MPQ    ��    h�  h                                                                                 ��B=��5^��k���ؠ�0ҹ�/�G�oۗ����/��E�t�Me�&�{�h�:h��j�kp��R�*4���Qߠ��%�h�8U��K���q\fo��I�B�<�k�枽��{gM?�;k��ã��o��K.�����}$Z�=��&1Ϯ�ߓ��8��K�?F),�!x�DC6�]�����Ax���e�暟g�e�Y)�s�=��R�*;5�h�@�BoI��>�E�:��D�gU <�9&����R�䒁j���Kn�7X�ɜ.�@-Ue�h���d�'ӣ����}�RO[�a�>����t4 ��0[D":��K�:���� ��'��g�>�g@�
�à����;�ڛ��.���6�{3���5=��� F����^����G�V� \�+�䩇��V��w��{��M!nl�ġ�-�2q�LQ�yJV7bBr\�Hfd�D8�s�c��I��� =X0]Z��|��穦�ѸB��63�n�>||�ү��_�7.�5�l����ͅ'F@�y0\��\'$���"�:=x�|�+�oU�>K �
��JX��(0�x2M������T����g��w�=y�h�L[� �7Yr�GƁD�:D���*=Q�v�m�j��"�/��@/T��Gn��#T��r���0'�N�P_
�ý5q�Y
�?h%�Bt*~DV�@�ʗ�=%f�!���D�ntWi���)���E�8�ԗZ{�+Yp�Jص,b���B���0JV�,��L�~�����1�֗@��w��v�VS�Ax���b����H���k���L(�E���sM{�
*�P�C ��]b��Y����<��V�":��R(�S�G��²m�	�����r��.j��i�cc������w���k�$%ئ�pVٻ���Sp#���v�c�КxH�E���t��5}�����Ȯ�0A��Ev{��[B��hn�
���cz6;��ڗh�+fBa��(5���3�~�[ű2�Eͥ	�\&G�Z��qr�"��!E�!c��s�ҪA���"�hдj|~��V��1XO�/gF���ޯj��el��o@e�>�|V�n��hyV�- ������kP4��B2�7+Jƈ̌IM�b��[�M����hP��@яB��sFL�8̠�B8vGʶޏMxo7y�E.uG �f:T����[i.�~a8e�}a/X$�
�Z�"��d�2W��J33:��`�J@
a%�������i�D�xi���1%�%�P�s�Ò�?�4���,��������9��QU����m��2���3Y�<m+�/��Q�}ZG��u���)�+Sԥ��3A��P����)�fT(���������Cƽ<���\��V���^� -=9��i�zJT�v��U�f�926�>𕣢��o1���},}��E�(�	���0>��� ��"sDK������]Ӑ4���>\���2����^�b��FB��y��]�ߵ����i
-���g�I�)��s��UϬ���i� |�~�E�t �潨K�����=v��Ŵ���s��j�z��Ϣ�8��l�Uj"f���!�^�˷���+ٵ�A��xL�z#{M-z�����<�Vq�@�D��U#z����N�秌�.��:f�M��R
S��w�D�x�B�@xZo�������/�k�D�2��x#�#P7q�R�C�-�9���i��.U��Ɵg(�R����dWo�&�XNdw���@>��q	5��T�K�,��m?2҄gt���g.�C2ݒAadP5z(\0�*������y �����AS�F`�a����/a�ˍ�<��:�1��{�I���e��� �Y��
=�FL���?��"�mjX��(��� �!�c���ӁQl�`���4�NvuZ`8�T嫌�d?N���J[�lb�F�i$�!��7=�/&�^*���!�⯵�$f��qҟBw) ��ؽ���2 ~�u/)DA�8�ra�0pN�ρ0y5����f��	����ТD�E7ƽ���]E�:�C�J�Q�(�*<~�;m��������@���ް���
�eH��r��yu�4�&k��f[�@���y9�4�M�^��L���,�4 ���I|0��z�A���{�Xp�;dP��T���ע�?8���=#�٧��ipUf@)���l��{3K[Ǐ��^g�˜����$�iv}���ťhPT%�BRi�j8���o3��xv{��<�����X`���bҷ��ñ�>2�b$_>T\�ր@��U����	g�26��mt����u�LN�_��%�g,"z*�GB˧s��Lbw��SQ���BzL`0ne8�M:��x��l�+���c�6p>��f�p����v�?Vm� �L 鷤�f�&]�UY��u1��'�����f�\㆞O6lD+�z���8R�v>#��6����ay�pl���gp����HA�'�Q������/R?$�C�|/V�؇�1���M+��3���H�����4��'�z����R؂�|����J��ra9��H}4Jƿo^]�� Øt�����k����s��T�k��\��	��Z%�ݭ�H�N����ʳ�y�q-������о*/�}�������!Yu�bR-� �07���6'��L�k�F��]Dɖ����)�;,	��苣�����q#�e�v���֢fZ���R+�x�j��,�������Ƙ�_ޚ��#M�~x���zTv/}m�|W����C�孟żan@^~�����h��|$����ը~�d�\�bp��z!!/�
�I �������4�)�Rp��r�8>%�^�� b�ߪ�Ns��Z��xVCu.�w5 �F�/Ʉ��x�@�^��x�����<�8�:8�0R今�(�[�"r�c��R�c�psLH�4�J	q���ƙv!��Y�&�&o�HX����Q�	O�8�\{4d��%6�zBi*�f��c9��Jh0*��wlN��_W�;�Zيڴ�H��� �#"1<�<��q�UD�I��r��*X�|��6j'-���+4Q���DhhQAQ~S]�k��(����w�ͼD|)�7�a����bY� tx��Q��`2e�g��Iz��X����n,|n�<0v=8�#������\�/�\d�J(�M����5�L �m�¿�u�\th����*�뛩7:����M��DWҘ� ��g!~w0�GL���^F�w0��{���D���M���D<V����'��������}����:�?O����t��I�ï��o�`�����v���E]�����2$�k�>Nq�o����SYt�ܞ�~9����)�����[���׆���Xt<]r�i��*���5gο�Vp��Tr����\�j��H�� 5���;���|��^��������UR+r�|��VԔ��ڬ쯓�ng�N�<k����>Ll�J���b���ж���es�H¤oH���XKdZp�"c�J������6.L�Ι+O��J�'�L_$m�.w�l���h�F;fy�6�+0$і"��:|ٶ/o��Kf�K�XX]m0bS2�N9�08��j5�F���J����hg�6�;��7Ԉg"�=D��|�)�R#Q��XmI1j�=c���v��tT7��G	�#Ofer�8�0�h�٢
(�w��DYEr�h����=�~�@I�X�X�B�����
�tt�"H��,�)A�`E��rԲ��Ҧ���%jz,�ZA*�A���oJ��Lt�m��c[⏂A�s�F1�@0�4��IQV�ݴ3?ʋ}.��K!Ķ�S-�qaL�����r��؄��/2ު�#.�8�,HE�RR��ο$"p¡��c�n���0Bm�Y]	ɸ���ۖm��.��6�$�c��z��ЎR���=oL$����o$�t��m��d��ަ+�S��܀�σk���k�6�и��w�K��wbmEQ���'��9#Gn6��Q��:�;߆��ㅾfKt�cZ��| �~ֻƱ�?s�`T�\A�Z��rv���Q맼�*�nu����Y�h0]Yj���̖��l����	+F���
 � �Kz�o���>� �|�ʫ�ev_V��ǉӚ��W�4�W\26�pJ�ˌ����w�[ʚ�����hD@|B�y�N���J��c&�q���9� x*9��`g�G�v��R'T�W��V�@.��a�Ƙ}��sH�
n�"ԩd��WF��3.'�=@�xi������#�i0�yx��,��pܘP<.í����y�ؚ,��O4��i�9"�OU�=�S��a���_<���/����R/Z����.^�Y^�&��l�A�tP�a���B�f���(V�!��6�r��Ƙ*�K)�\P�I����-�-�'������Q�iF������2�_�P���g�F��}���(^�d��g�>��K x�<s_���j�؞���ܘ�44Y��9���W��r,�y��E����.��2j�P�����/
���"}Ӡ {}�U��L�J� �~��E��ءCsK����j��v������j��e?��4����Yl6�}j��ǂ��ę�����k�i���EWx5_zz��?-U.�p�קXVlN��u���#1xSr��N��ҌL��䂘�f�T���})D�a�B�LFZJFJ�O��*.yk�����=x��PRE~RV����%°���.P@����E��s����W�&�Jd�H����N>�x�qd�c�L���|e[�2�!teg�m�C-E����P�(w��* ���+�y;Ǚ�q��<Q8�a�|`Oʐ�"/��Y���{< Au�̾WD�I#��e������{��T�
IIL��?$Dɢ�j�x(�F �w�����FQY� `J���/�vИ�8�^p��:Q��o��K�7l�BT�dNV!�#�=KĐ�yV��L���Tw$�����"�l�sBҽ� �#����1ڭ�Py)�H8+�F�+0�NG�d�#p�4�I��v���aZD6��Ƹ/v��/�I.�^�ܢ�h���?�v��= +�K���4صAU��7����e#���A�X�/.�&�Mr�D�5[����؆��ę��w%���я��� .|K>�zT�H��w��TB�֧Y��Ņ�'�#��8�Z��e��=��7���)�Jf;��LlG����3f�W�I�J^B፜'������vxה�n��`��T@�6R�H�j�¬:M��w��{��I�^�h�Ѡ`��bMUv�� '���x>O?�ۂƘ���g���6}��t��d� =N��Z�U���"!�,=N�*|�B�JB�(Kw ��SL �`��8��:=t���2�f�i����k��r)p���|�?�6��!L[�ͤi�&X�AYDoVu�zB�o��A��\�6O�r�+��z���8$2Y��5�Jžera�@�p`c�Y���H��ͻlnW!_<�
L�$y�|��)����1;��M����NF"�û����4�'��%�6�R3a7o软�4Sf���9
=�H�Aƺu^��Q ~	��)BR�x���]�����T3���W[	:�:%�ً�c�sm�ʎu@"���J@���l�*���h�U�*RA�<C�u��bhN� 1$���U6gm��ƹk���ذ���ԫ�d�,�]���@�?�y'����+b4�A��/����D��)��g6�����~i�L�M��G��9�Q�?v*E�D�Йs�C���@
�n[��"jx��w�:�O�f�c�3d�Q�b�1$z���E����%�����O���䖂p�rd�%ڱ��;)�z 0Nn۽�ܢ��3�����w�N"F�-Q�� ܝ L^�I�f�Z�U{�<��:�t�R�d4�c�:���dc��󲾲Kp.�KH���J�5�����𡨫�&���!A����lE�O(��{\���&?�6��?i���O��V���u*�lhl���_��;�z�5ԁH�F .0A"���� �q/F����]��rX�X��Qk�'���s�4��~����cdA��]Q�R�C��Z�6]xGD�/�7�/��C�b��� ���t5�۸]�B��I��X%Ȗ�ix�nI�b01t8�>�/����\�j��dP���dF���5[�Ĉ�c�:�i�7 ���]x9�떋�:;��;���_;z�S;�u�z!C��0n��͚F(N�{3��׿np��Oc�O�V<�n��8��\Zm���7"�"�����*+"�p�<ê���H�Х<���SHu]�[����U����9\�=�ଊ�S0�C�W2�~���=���Ֆ��4��P�&���t*��rH�����p�n�q������`��C���߂�0O5�L
�vK��^�TX��C��vo�+5g���p�V��y�3Z6�J�;nb�4��䧽���L���J
��b��ͤ�Z��z�}s�M,�����?�Xf��Z�T>*���z�xA�6)����A�H�B�0_��>.R�l1�	��zF6Ky�0���p}$�"
��:�~|b�o���K�����2X.0#J2C:Y吋U�� ���B��J���|h"��Vq'7O����D7�I�ĝ�%Q=M�m��X!#���SjTr~.G�U�#J-5rU߿0�uE�.
��x��_Y�I7hR��8x?~��h@���s-��cޯ��E�ot�L����)��(E>(:��8d�!�t� O,�G��K
���JJ�/����B�
0�N:�1>��@˗���<fV	0h��狘������j[��Zt=L^Y&��0kV��9h�JrT�9gl��3FV"��'B��H~"�j,��oC����z��m��j	ҸL��h0E. �%��&Rc�l����-�^�x��$7\��Վ.�qr����z��e��Y�Қ.�fܻA���ϫ���y�jR%�f�	����E,���a,�Ԥ�n��?�����;�]��^@�f�Tj���>��L~�;d������\\��Z���rQl~�9�ŧW�N�i`$�`v����hK
�jr� �������e�F�r�e���M7�o6|�>��|�0]� �=V��k�gӺ�uc4��}2���J|�Y����[�F>�7(�h���@8��B���)�l����)l����x�Z��{��G���^�T����p.���a�G^}�h���
��k"�`dM"�W�t�3)4Ă�/@���-"��ʹ��ik_=x�U��'�"�˳�P�أ�� ��<k��,@B>���@��9}��UAg;�2X��(
���=<�ql/2�����Z��ZB@�)I{�!^�Gg�AYs�PH����{4f
S�(`B�kc�����s8���\�T��a�s-������p=	�,Ek��M�o���z2���w;�.������}�$^O�(�v;��4>Q�� 3�:sz�`��j�f��Ӈ�4�ۗ�4�Ղ-�Ԕ��O���̪wͦ�&(���5���
���ݗ��;��i@FU�V��LJE ���~����	'�\�K�����va�Ӵ)��9?�`��Y�uݮ($lQG�j�����6�Ծ��T�ؓ���K��8xP�rz�>-0���R=n�r�Vg���P���V#L��킸Nd魌����L�f�{*��N�8�$Dk�Bxy`Z%����c��L�k����#~x�L�Pm9�R��u�`U�;
�.K��U c�ȶ<����W�Ӳ&o\�d�Ǽ>��>� q�#Y�ʾt���h�2���tH[,g>͌C(�����P��(�z�*�x9ݝ�=yv*���7ok���`
S�=�B/������<[�#�g��-�I~�&ed������OCy
��L��?��}�V,j8�(u� ��YQ{�`��Q�T`��1�*��v+�f8T����570֜&ѥ*l����_�j!E��=y�̔���Ǡ��e $�+�H���g��B-r$ oc<��*�(5�+��)�k�8��ö&�N�ng��΃Ó�\y������NFDєBƳ��:�����y�6�G����Q������B���+T��p"0�0�n� ��e�D����4�*o?&!�g���[�揷�惆����ԉ'S��0���a�|f�z�D��c8gԏ���q��ǜ��>L�z�]�ucO��}�=�B:��y��f6M���M�a��3��P��X^�?�b���Z�vsD����L�x�T[��R_��j�uJ	��{��ʹ 9����`ub���t��[/���#I>JB��6���7�&:�g�*6X�ct�k̫�Nߛ2�� [��Y�,X�f*��B���ciw��~SG�I���a`��$8��:���r����l��G�f�a���p=Rt�Ң�?L ?�2L�1����&S*jY�}�u�T]�Z��Bv�\Y�Ol��+�^z?5!8Ȉ�t�<�Vř��ap��u�ѽ�l\�H��w��U?�)!��e+$<�!|e��·�1��SMy ��i!�>���R�4WV�'%*&��R���t���l�꯳N��2�9E�7H��Ƶ��^l` 9��D���U��8��o!T�Ɖ�RL<	�ߚ%S��~����cP�i;�]T�������(�*�I6�#2��E��·��u�$#��~ �7?��ܯ6������k	�-�S=䖓�Pԟ��,?�H����u�4���:͊�9�����jwr׮m���F[D$��]XW���|�� �M�B'�����v%-�y+��TF�C�
��wDn�w��]"Q�ǯ�rj"���D��d�f<bf�Rzא꼀W��PV���ڪ�옟p7� r��%�$�vި���Ni$j�7������w+�pFaKi�#c�8!�^����~��z;<�ď:.R�-����͇X)Tc�wвq�p�?�H���J����b#��߆�F�G&�Zξ�
Ԁ����O�E\��\�����O6�D�i�㶅
��"��<G*e6ilĮ	_9�;�����:H;1 I�"'�V�� qjV
�,:�h	���pX:��l�0'#	C�N6�4ǫ9�R~�^�RA��]�N�^w��F8CBD�U7"d���b~� ��9�ݷ��V_b�S�I���X� e�d�n��)0��ܣY1K�����}����d����6�5�]ģ� µ���'(�hW둍;:�H���e�z?@Ҏ���P5�!~0	[���g*F�����b{N���:AX�\qE�H}<��`�����l��(�՜�k���V���p�e��	KåM�%��`��ᚪΰp]��[�h�Zs_�4��j*�g#�SK�����e~��xr�5���-�ɫ�F�A!tERdr�Fx��q�̫Y������M�]������4�z�5���ѱ���`^����X�`�1��+P�ڇr-V����n����Mn]Iw��}5�c_�L�TMJ���b�~��8��s�r��Z��L�2X�ҾZf��A�WJm���6$��O�T��k]�_8Q.-D]llu�Ğ|�F1�AyAKN���$��"�}.:·8|O-�o&��K���X�#0>R�2�Ee�k��:�|�~���Nj�h�_y�qdz7����eDr~��_�4CQ��{m���s�������$T�j�G?�0#EAr��H0X�L
xŽƄIY�@qh�`~�3*�~Uʓ@������3�6�ފs��^t(�n���)���E����פҜ�����3,U+` k��/�Jg(�����W�����)�K1y��@f�־�O7Vd�[��I���Q�A2��E�s���mL��Z��1^�';��eҲ��ʖ��z���s�������"&37��C���ʺ�m�m�5	?�{��c��.{��𚅿c�A��	�$�˝̳��$�'6���t�̐����L��˂�ƚ	d�����Ϲ�o��]��]�%Ƕ��ʒma�E������oFln�~��Ȕ.;UƗ��f�~p��
����~�۝�C^.��I�\w��Z��zr,A�tԧ�i+�dˏһ@n���hf��j�o��v���i�� ��F�:����+���"R�Uo�7>�6�|��ԛ�V�����Z�0��4~�2,� JW�x���3��[�᪒s�h���@S�Bu1��i������M�g�׶�x��s�9�G��:��qT=�,����.�DfaI�}�5x��c
d�k"�7d��W|n�3$a�q�"@;�Hi�>�͏}i�x:���"�ގ&��P��=��:�y��c,{
1�����Ϝ9��U��}�M}��V�Āk<EU/����N(ZX)����DY��-�"�A�QtP������fe��(���8f��hP��Nf��\��w�
�oT�-n?������%���:&�`�su2G�����I���<�t}�����h(�]j���?>��q �s�S��`�h�Ak��X4�-��/����*�^���D��;�d�R�/�a=�߆�:�f�
>?�Ș�S�V���U`۩�j� M�N~�����
���K��?�`*v<�R�d�6��I�[����_o�iyRll��j�H悥��������X�<�U�rݜxk�rz�>I-Fɍ~ �Y�Vb&*�QL��I�L#gԱh��N?9�����f��cm���D1��B���Z �ٜ�I��`�Mk���Cu�xT��P�M
RL����W���N�ֳ
.F��ư|����	�ۗWx��&J��d(����2>˨q�n��Q?��[�i2c��t��'g�L�C#ؒRx�P>.(�O7*��x�y�����l�2�z��
`����X}�/�K��\�C<�=F�JH6�I� e?���+���Qz
���LI*U?Z|��*�ji�`(0�� ڃ�Ԫt�;�Q���`���%7�v�u
8�ҫ���<�wZ�U�l3Pw�Z�!�V=�M̯A�B���@�$�P�B�b�B�Fw *����\ڣof�m	)�0.8aXٶ!�N�m�a�Q�jb����������eDll\Ʈ�c�nd�kQ���X������{��잜�s��W��A=�+#o�K⍲{��e��#�J��%Ј&|.�躩�[��f�M;�����{R�6ܞ
���E�H�.X|��BzJ�+�>����������5�5\a��<Ǌ[z(=���Xȝ�:�;f1A�O����3�G��?^�^�.✝����F#vn��$���/-Tv3�R�MHj�b���g���f�{~_8�X)�G�`�(�bC�w�K��W��3S�>Ee�֑g����A�)g�X63#Wt35��F5�Nډ�Ό���,s�*r�dB\�/����wV�qSBR��S�,`a�J82?�:3��� m��3�4�oaj�(8p������ ?�)vk�Lх���!&Ny�Y��rubN�x#�>��Y�\�D�O� +4z���8�U�1+���tcYa*�|p=� ����Hr�%��\������$wCw| ���7U1�9�M4��܄
�ڹS�7�4��.'�����R������I��*4�o�>9�3HN��ư�x^nq� �J7�_���n!��X��$Ti$\�M]Z	�{%1Դ�[?�iz��D!~������۽�*@�����`�`n��2�ur��ކ gk�䃎6Z��}I>k$�����c�n,���e,�z��ف��Ŋ��ڌ���!14�����9�Iw`���f� ��%���Bc�M}��C����x�v 57�2X�9�C�c��68nѴ���]S�W�m=ƹ�b�ٗ�dۛ�b��Mz�x@��:ɯ�ŋ�!p�\Y�Z�pR�rZC�%�����̜аkNd�撓�������w��F<��^\���A�^	(T�2��˘k<��:���Ru��ِ��{c�v�tO�p��0H�w�Jz���	�'�?���"&�$�YG�KK���O��A\,#��\�6�ٮi;_��B9=�Fyפ*@ zl��7_�\;}��rH�{� dTt"��x��)_q��;�d���G�(MtX��wˇe@'�9D�)v�4�H�� �Y�Ab>�]�-��y�y�P�A.�D-��7�*5���bj^� P����6��%s���I++AX[�K�_pHn�Ր0�A%�t��%��ά� �?�d��$��0�<$5��ľ4��0x6���?c����댯G:�"���Еcn�	���+�!�tJ0�~��T�F�FOaα{i��׵3̦7�7��ŷ<'��Ȉ��Ǫ��&2�\�9g�е���禘à�;���I��:��I98]fk�N���m��/���7��"�jSfi��M��~��ۼ��Ѐ��F��!���d�t`�re���_&��l��h�������~�������,���A5�^S��V��M=f^�����@���+ki{���Ve ������'�nX��M7��DL��J �rb�m��4�f���s��µ�@���X�9\Z�]�=թ�t���6
Ϊ����� x;�_��.��l�UI�9d�F,��y��\�H\�$"�T" ^|:�wB|�o�2CK���\x�X�/�0YzT29q]�F���@���N�����gh���یw�7E�{��D������Z}Q��mzE������[ �fT�v�G�\�#@�r��0�L5
��^�� Y�Wh�_O�.��~�۞@z�󳩵H��V�eV��At������)R*�E�����m�#���(,N����c�{��Jm�3���
� �ÕT1���@����V�4�dx�΍��j� ˎ����L��g�����	��6��R��/N���m���8�#3(ӿ�%"���>7���x��p<9mo�5	zd�����^8b.֝��U�c��ƿ��������;�$m��,��'ϱ�?���"�Ot��W��1 3�Th�a�G�i��[,��1���E�6��G6��
�n������O9�;0lz�T�f�Ȇ����M&U~Ǜs���͑�6\���Zw-�r6ִ������_V��+���9�h���jh j]�Yț�^F���� ˠQ��m�o,�>��B|B]�6_�V��4{����4'A�2��J2�'�5R�Ρ[�����ބh<h�@n�1B����	N��h�4��bcT�J)x[����GL�\��TxM3�'V�.��;a���}M"��t_
߸�"e.	dæ�W��3�ڂ�z@�Nc�X����j�ti�� x�>��6���IPm�����H�WR�>_�,��W� ���93�U�b�h�u�����x�<Y8�/hL���nZ��3�0�_�m�a����yA�O�P~R���M�f�ci(���S�����|�)�����\!޲�N��g-)4A��L�f�n�������$����2��!�����dt�ʷ�@}�L+��(/d񦭕�>�� ���s�/��HӞm!�I��4*�*�*0��h>��.2��]��0��-���rV�!���z�*
��j�S-J�q1ʢ_�U;���ª� ��~�4MV.�ҔkK8���]v""���;~,�V�5�%��$��l�7gj�ׂ���JK���z�������-مx�X{z`-�7���&ب��V]�m�g`�	�#�2��:Nkt��y��S5f�)Q��cK����DL�sBn2yZ��ٜ �����;k�L����xfP���R�a������9��q}�.A�H���>�����W�&%��dc�<�t�>�p�qu���@.�����2>�t�kWgt�C�N��jP�k~(�D�*����Sîy�P~�Bw--f�r�a`���s]�//��7P<��ܔ���
_�I4IgeڒG����E��
��L��g?�\9�\j���(�� �9�O$����Q
�!`g>� ��v�n8�;�����+���R�.G$�l���U��!�n=|B)�ʚ6ʽ����A$R��~��]f�B�:� �B��)�=��v��%)0�8�䆶0�NX������p��R�/�u7	��ѹDd.Ʃ�t�ɮ�&�H��C�=�/��{e�'����6�	
�Q��C�f����e�z�^���ӎ Q�&����uU�[F������L��J�Ho}��Ѡ���dc|��z��ߒ�	�ǧ2ƣ����8ް�)��5��֖�=�z�ٓ����8f,���]p��'�3�+z��Ŷ^Ӆt�������vi~��T�őT�ERU oj�d���/�HK�{y��o�9�i�`���b���r�-�џ��΢>@���	��A�\dog�S6{�tn�s���N՗v�f��S+�,���*��B7�N���w��\S=+��w`��8M��:���\���/��H\���37p�O��OV?BSQ��L�H�:��&I�nYU� uh7�t	����]2\���O�F�+	>ez��8>���S��t��O�aeNp�t����"��H-�׻�������W$���|�H6��y1L	oM�UGܟ�4\��t<J4�v'[YOݧ1RD�Kh�J�G��ԃ�Jr�9��8H�9ƫG�^ɖ� ��z�#�����4�_�TT�&�H�t	K`�%Ɍ>��.���$�'�Ӷ��_۸ J*� o����{,�­g�uMf�S8 �'��J�6x �8�&k?+��I�/�I��=,u9����Q��������BĊ�H֢ҵ�����䠢���������G���;���(MX��~t��"�v]]/ZC��K(C�����n������h0&�`F�Ք5�d���b\�z����=0����ߤ�`�%��jpm-�rՆ�%kj ����KA�N_���;Ԩde��Ww!�1F�I��u�n�Y^|�wH���?<#�:$��RPR����`�c|�>��M�p_�IH�x�J�B������bͨ|�U&����=���[󽩤O�1��6\g]���cZ6�� i�l��"�X{U���**�l:z_oI�;x�ҊF�
H��� �"�Fը��q�֠�������A����X��0ˢ'���'4=B����nT �A�:]��s씇���%)�8�Dh	7XX�|��b�^� �����L��ӞfIf�1X�1J�ZnZ�0b����!���V·�!d!���i��b5���ٍ«����'��I%4��:L+��l@�а�҄I��Q!�y0?�~��a�F9��{��z�0F̦:� c<���`*�"�K�鲜&&����#�������b�AH�Ûs����֖��U�8����]A#��������*F� e��ݴWS�Y#�Ȭ�~�N ��γkh����ay���t{�r�����m!�!�ȿBY������qD��H~�����m�5���'+z�蘤^�a���'��|�+�d�h��V@d������xnS]����H
L�l8J{��b�| �o���K�s�K�����X���Z\�3��x����I�V6L��)ېy�����_�z.��l�U7��k\F'�cy�ߪ��$=K�"{^�:���|�#�o\�`Ktl����XD`i0t��2��A�!\N�{��{��o���hS��ۧ�87�"E���D�(��w��QNm5������<��&lT#�jGu�#;Brf��0Ίv9>�
�C�|܎Y1�ah#~x�)�~�@5ZE�ĩ�xr�@���t^�u��`�)���Eo��v�Ғ���-,��e����v�J`�Z����{����1�O*@�VY���V�vً�B��7�|��2��>�L/YL��*Q�K�s����'���¤���@r��h�Ӻ�s"�#���J������*�mJ��	��\�ݖY�.1Ѳ���c0���(��|,�)�E$8�ƫ�ق-@�� =� )�����k��l����g���P������}��c�KE�����2��qn��8Pc��
y�;K����/�f�2��O/���r�~�{���i�L��\���Z��r�Jʴ�R��(��Z��q5��E�ph�Ѽj��8ֻ�X�-�6��F���v5ʠ�����o��>\�B|}#*���V�2@�x���F�4B$2"XJ�f�p#�i�p[�
{�Hj�h�^x@���Bk4���F�6E����]:����x�D�̋�G�(�7B�T�4��$.�hma���}/���
Z�"@E�d��(W��3 �'�@��~g@���Ek|i� xp���*����P(���ooH��/,������L�\9�{�Ur��'�����z��<�K#/�a�ʑZ$�sQ>�z�B���O�A
nDP8����'f_(BK��n��^mi�"|7�\�.��E%��-��0輺��ҽ/�2�0\B ���2����<�����2�X}sJ B�(ʊЦ��k>b� dV�s�+�Vȩ����܄M4�0(�%���â{^���1�7��q���"߼�P�ufa
�=s��d��4�� .UE���
� �sm~|���ؑ؍�FK0��V��v�A��{��P�QK�j
���z�l��/j���[ʟą��%�?���6�������x��z��-����a��C��VX~�������%#���^�N��_�8���&�f��>���i0DgFEB�wZ����;Xb��h�k��ƺ�wx�"�P��6RB9�tjǡܫ�g.<�"�fջ��-����Wn��& R�d�=��Kw>�X�q�y����@4�@QQ�2�ft�#�g��CQ��}�P��)(�Y�*B��.��y'Ȉݡ�(�-��`;��ӎ]�/�2����<��8U��I��Ge�5����Π
� �L��?�]��2j��(��� pʽ��8QE�?`���ռv<ґ8��E����:�-"p��li���P6�!V	�=7W$��F��8Ϧ���$���C�XۜB>O ��P�D��ڙD���P)kd8��̶p�N��0�ă����ip�P�b���AD�{�Ƥ�A�$J�`��ʅ����/�q�g�b���j@��DeL�ء���r��qn�e�E����v���&2�H�0!�[5P-��yΆ{ą�d��6� p���x�풻|�6Oz@����:��@E��B������!G������N��Q��=jF"��6b�p�f'�����s���c3�/��5M^����>`�+Z�vdKg���%�L��T��YR��!j���&��O�{to���fj���@`��b9*M{@�G�i>;9�G̔�� �w)}gu{6��-t��u�|�oN�������,�N*h�iBބ�w�@S8$9�	�B`��"8hU�:)�]�7|�R&�j��W�a��v�pn��#��?��E,=�LG�/�հ[&DwKY�h�uءs���G����\
c�O=��+��zP�*8�vůQ!T�*� a�)psf~�z�Ԇ}I�H�$����'I�vs$�^|6�j���81��,M�0�ܺNگ�a�Oa�47'� x�bsR���#F��)d
� �Н%B�9���H��Ʀ�Y^$�� j���9�de��-����T�?��Cߊ	�л%�-��!��_���L�������۳�*����T����
��(	�u(7�T?# �2p��1 6��@��L�kZ��ĢG�$!�P4�,l���hᬈV�e����ۊ�䢭ܮ���\��]�U���Θ;�8HHM3X&鹁�����v���NЅ~�C'X�,�#n��x���φcCB���_�O�Mdf�b�ӧzh�ܼ1a�P�,����ڻvR���*p���rP��%F=��'	���6�NZ�W�H��9D�e�w�H�F�d�Ԯ��	�8^��Α����A6�<>�:���R+H��O���),scw�ϲ*l�p�&H�4Jp�A�`~G��m.�*�&����̀���ص�O��eU\�����6�ci�௅;"�sr�ol*�S�lu~�_
V�;s:W���#Hlq ��G"���Ճ��qG:�P3h��H����;Xk�-˽߷'�����U�4x�c�#�O6HA	$]=O��?�F���c�D���7�w��b  ���.AW�����t�I�-�X��`�U�n�L?0����{����b��VXUd��:� G	a5GUy����&�3ڣ�ٯ[䳦�St:����'�����0ޅ�Yy!/��0������~F����]\{�!�׫xX��L�; i<]�Ǿ�X1�}y1Y�W�A`6�����H������Ö6�6�Б٨p�3�?�+]�u�ā,+á�%�c{�����S�i��C��~��Լ)���H����ɼ��rL�t��+r�2�q���\����iś��i��燨������5_�\�b���^�P�i�+�b+�딇�)V�>����ԒnNg�
��m�L�(�J��bd��à��A�s֡M�k��}>MX�g/Z����,�*���sh6� �`xN�40��?R_�X�.�r�lvY�o��F"��yRZ9���[$Xȹ"�~|:_�F| O�o�7VKZ���X���0�*32/(��6,��9��My��N/�_{Sh�<����7;�i	[D#�E�0�<�1FQ�z�m����Y���=�bW"T^��G�#6��r��c0�|dTg.
��t�W��Yl�h����$ �~f^U@��z�߽����D1s�t�2���=�)JE*���9u����l#C,�<!1��q��Jx��90� �q��%"���;1*Ȱ@7֮��HVu��ړ���;��ֺ��F��L�C	��h�o��l����>�%�����2��Y��ӵ��"7LX�~�����f9�m%oA	�vf�]�T��.�$"��a�c1���zM펙|�dd�$�J���J��ݫ���J[�;���E�h����ܧ>ϊa��{���ڸV�Ð��z���QE��`Ὂr�@�n��O�7����J;f�z�Jj�fd�㤊����߽~�{�T�7��.\���Zm�r��%#8�Ð�U�:��_y� /h��Ij^��H���V��F��{�ъ)�ǐ���;o"*�>7w�|�	��l�gV��ԉ�<�aҵ4]'U2���J��5��m��[�6r���h�u�@��sB��]����qAܠjxIX1� ��x�!S��d�G%��T�;��]�.�*�aZ�5}�[��܎
�'�"|�d9��WM3�ႂ��@l����v�,� M�iWx���U��7Q`P�#��4�=�����X,,#B�V����V9��U-��䞬~����U��<�~/�a����Ziь.���I �(���2�AE�ZP�=��ן�fv��(�.훉h��+b�߯�rW�\W�q��5���-��1�K.U�\��ҘhSm':�T����2X�����Ț��ʭ5�}N�8;�N(e�����>�7; �s�Gl��g��j^ܿp�4`❶ ���'$.�� �����s���*�=�W�?�p4
O���B����E�UV~U�)�8�� �~w
��5�H�eKK���>Dv�!��_qCz�L]<���ݚ+6l���jK�6���W}��X������Mw��0�x���z"�-�k��>0��RVSZI�b���zv#�N��HmN�l��s���Z�f�Wh�tPH�$�ID��^Bdk�Z�1J�v
�1!k�9�T)@x���P�I�R�0�OQ�L�Ȱ�p�.71y���و����,U�W��&���d�
���}>�`�q+�p���wO	V�ޠ2��t4�Rg���C$p�c�YPoG(��|*}��	s`yb�e�x�	#'ў(e0`���ө}b/V����<G�f��
v �I�9�eP���#�^�;=�
_>�L��I?+~U�f�jzEn(a�� +Ewi��hmQ��`Q^+�� v��u8@o��.`(!�+����"Bl���K U!��=�� Zʳ&��N$$��'�v��Sp�B��p [�
�_G���;��ʌ)�@82^���N,��Y������HO]�+A��:�D=��Ɵ������6��p�3��L۹���n�D"���Z���\儰��[���Rej0��`"�S��M&�o>���[P��x@��VX���L~@�����V���M2f|҄z��˒�{�{�����ѣ�8��Wp�f��ߊ�/J=E2e�	��h;f"2���M!3�SD����^��i�N�%��v_8R�5Mn�/T� �RK�`jZȳ�a��~tK{o'��%��x��`.��b�H(h��G�����>6�֢�蘷.x�Sg��6Ċt���ŘN�+��b��|�,�!*��B�X݄O"w'uS3=��d�`�$�8��:�̯�j~���B�ʁR�D�9�p)�J�>{y?8�օL�Bʤp�L&?&dY��u��s�v���p���\E"�O�s+��z�ZC8�[8�+~�S���<a���pxq�u%*��-�H��H��10��-�Q�$(c�|�!7���1Me+c�ՠ��*g��*��4Ca'�Y�=qR� ~����D���u� 2�91��HD�ơs�^A] %���7��C(����ՈXT:���>P�	a%?����4y��})�Ւ�I��Q�GۮX8*Qw(����£�7u(�K� 8���8�6.�4���Ckuݘ�?�����ԋKd,�(�ʗ���� ����[���^��#t�V@r�T����p�Uu�I���&�����MJF����X��v~�z�@�4CB���mnb+n�IC�$��^v�K>�
��d,��bRzC�"�l����:$�~���4ߘ�bOp�vr�m�%!0��bW1ЁLANU���쿨�,7��w#F�k�Uܤc0^����-\����<Y]P:��R�֔�]"��Ccr3����(pզ�H(��J��K�;r����c����&�B޾j���|�x���bO�C�@�c\�1e�-�E6�XxiLuX��A^���f*ѝl�;_��p;n�w��P\H'p ���"���^��qV��������j�9��X&�n���'����4�Xo��ȔJ��Asn]�)��0�������D�.�7�yr��b{�� �Z��I��B9j�I���X,Ï�P�n��0�eף�)������=AK�=dW ������5�
��F¡M��~[hw�bq�}Ք:����/��i�z8��P�!j��0u鮴ےF�(�շ{����&�p��8o�v��<���p��ؐ7� �\������a<��Qt��w�Ñn�T�L�j��5����W]����t��h� �����S�]S��믾�U~[t��d���q!�}Q�����-��t���ry�݊L��̗�>�x�뛭V�'������8�͂��5:��ѝ3���^�_��ī��^+���^��V����Z�S�Q�nI��^#-�O��L�JqR�b?�Ҥ�����s�F���):�8	X�.eZR�����C_�P6�λ����~_NT.��lX���
��F�uy���y��$se�"q�.::A|;��o��#K�_��mh�X�!@0��~2�����1z�񏷐薎�릺k�hɎ0��p7���D�wD^C������Q�Cm�y��߷A�x_=��T�[G���#1��r��0D�o�"

j�2�Y�]�hY��2�~�� @�s�����nT����|l��t��\��:v)c�E�]�T��҈ʔ�Guh,������l��JӅ���)�;���qsS���1e`k@�u�����VЫ���y���-ԡ��b��dwLeN�����ʨ�'�۬ђ=���y�Z�m}A��3FӰ�"��c�o�_�z���g�m m	+0S>o�O��.�1��@�cLZ{���ݎt�{̟({$>���	��8J��p�=�VKق�a��u�R��+�%�a��Z��X�����uےY��Es���d���Xn�S�,�ȀX;�qǗ�Ĭf?f*��� �lV~�����&�´�\�U�Z��r��B�`�^�΃P���'�R���1h�K�j�q�%�Ζ��ly+F�R$�, 頂����o�eb>"�|���hV�e�.�ܥ~j4xJ�2EJ�A���%���p[������hm� @��PBa���p�H��]U��SH3�[��x��%�^�G}A��y�T)c@��!�.��a��[}~����
P��"��pdt�W�u3U����@'�X���G��N�i�Q=x�����玒�P���Oc�e�7��,gk��1��9D��U��0�Q/�4��0 D<
�A/9Q|�kZĞ��"��٥�ڥ�5A�
�POck��xaf���(�2������T
gƺ]-��b\�/�����!�-Z� �f����Q�s���������n�2�U��!ȵ��(�m})��v �( 8����>�> ��s�3�L'�������4�����{�y���]]�!�'�;��N��M����$ǻk�
���Ȅ��� �ЫzU�.��s+B ��l~r��g���KfϾ�Lߏv��p�P�V�G�	� 5�U��l؏yj65�`��\�[ֲ����k��^�Yx�q�z�X�-wqm�y��y;PVNV��yF�5]�#�PT�HN�G��~��$�~f{Ι��f���<D�x�B�7YZl����慏��k{�����x@��P��R8H�*X����ٰB��.2�K����og�G�Wd�&��&d���ET>�� q���q��jsG�2�n�to�gE��C��cP*�L(�#*���z1y��W�W<�P���`���Ľ�/|�}���<��Y�n�����IE�eN��>���
:�+L5�?ƾ���j��(ߟ F��P��qRQ�ɗ`�	v���v�8�8ɫIa���h��ic�QZl����F�5!<�=�������.�⬭}$�O�#�N%�B��� ���zڏ���r��)��8�J �P�Ni�WM�ƃ�Vt��T�����ub�D�
�ƚ��M�W,Ȥ ����k��';\��K]�������L���fT����g�eE;��������&�o���[k6��&��1���������ѱ�P��]|���z6���ܽԶ��x�+�����I�Y�!#���w�G��= >x�D%w��@fW��n���Ζ3�E�+��^dJ̜�B��a�vZE�������N�T�/R��+j5*ᬜ���X{j�fʀ�+�3Q4`I��b/��u���8���Q(>11����|�r|���gk�
6�BEtBw̲ߙNƁO�w���U�,�*^�BȻL���]w���S.vŢ�DY`M�8��:��w��Ș*���bM�C��]�p��YAG?��&��L��Hv&:��Yf��uNu8�',��:c)�\�.Os:�+��!z4<8o`L��s����ha�{p����p���32�H^$������,Ǔ$cX�|l����7�1]7	M F'���ڥ!�4~�',��8+RU[w�q��_���vΝ�Ar9l��H���Ɯ9�^��L �M_���Z�׾����T��V�9�	\�%�_��hG�U�ʰ��������۩��*�R���S)��&����u�87�w �y���_b6����i�xk��gǺ�[��[��Ƃ�,F5<�ŉ<�bˢ��Z�"�C�OE�c�)䑂�׵�9���l������A�֚.�+M�[v�/�8��=v�x@����C�C]��"{�n=蓬����e(�Yɮ�q�\����dG�Rb�d2zX���^���y�k�q̘F��p��rF%�B6�������NPq����u��@�2\Kw��F��S�J�U�?@^�7���?֭�S�<t�$:��HR������9�_#Kcm����bp��,HC<Jfp���řlm�M��&�����yԀ7^��.^O
}b\�;�Ȩ�6�m^i�)������e��*�_l먹_@��;i�4�W0�H��� ��"�b��9��q��	�����~����X�4����O'�;B���n4�όY��E�A�S]����=�<�h�D�v7)�*m�ub� <ƥ�d���/�d��I�{Xǻ��K�7nkCn0�\��������o���d�c1�����U�5�8`�*YL�*a�Y��O^S1��xw:]o%��]�48��_���g�!�}�0;R��H#FJ��Mm{��ס=������j<������3�]���w4��oa�<���|x�]Ì�춿�@@�����5�O]�
�:�a��Pc1���vS��+�9G�~67�����<W�x��rBi�賈t�9�r���'Ws���W��)��p^ꂎ�y
̀S���}�85'��g��k�^��G��s�ةd+��·�ˣV�O�������nD�(��\�
~L)&J��obi�� 8��E�s���!������X#Z͂�`�ĩ~�X�MT6�g�w������S_�c�.t�l�:ĥB�FCy��4��$�"?"��:w�|vto-��K�����M�Xu�A0�Z�2%_w�L8�,9���>���|?h������71��u$D��<�f��Q_�Emf ���5���P�T���GF�M#,wrwe60����_
�����Y�� h����!~a�@f0��F��+M�ѱ���Wt/���W�)�[�E��=�o�����"�,:w�gg8�gw<J.m���G�V�y���0�p"1�Z@m5����RV+��P/0�:"稌f��*��'LL y��D�%�Q�ͅ��$��@�5y��K���ɕӫF"����*FX�+e��\��mۊ�	f	6�>ܖJ��.B+��A?�cg0]�p`��Ow+��$$�ষ�Yٓl�+>�qQ�;F��Pg���%���������̸���"����EN��3_��vNn���a@��;��;���@?f0�� �0���~���
[4�}߶\��wZc��rsIǴ�#*���C�K®҂l�vPxh�jT����R�	����F�(�އ��=��Bo�>���|.6ԢU�V���u���I�4���2��J����!W�:D[�Y�7h(�@��UBܨ��K�Q�療��ߺN�����xGż�w*G�}p�EeTd����P�.�+a�a}9�0�^
��"�Id�/aW�.\3"ق8l�@➹��'l���p�iͮyxA���	e���_�PY	]�j=��2��X,��������~9�bDU�������
�4��<EE�/���w�"Z�f����ˉ3�o�iX�A���P�9��q�f,A(sVۛ�-��xƕ+^�I�\�����&6e�-/�����RK�N:��/i-5d����2��m�h��x�ʣ>j}���a(��~��=�>sJ" �D�s�b������[�5�b4�����ԏu���6hْ������숇 ߍ��f֭
�M�?،��9b�K!#U�S\��� Tj�~m`��=ؾkpK��R�ǟ�v�����}��(�BI��{z���l��j�Aׂ����6䮷�s`��f���Sx�d�z��4-R��ɴ���D�VIr��~��c�#����kPN��B��j*�!�fvp�*�E����D�AjBZ$<ZG	����Տg�fkvT2�
�ax�)P��R����ް��.-��w��*�H�bs6W��&�gadO��S>��-q�－,R��x�Y"2��t�g��C
*��t�P��(4Y�*s+xݿ�Ry�����Fì��`l'����/��=����<����	��B�I���e�!�Yc��1z5
Lp|?a��.j0�(�=# aR�;J鵂��Q��`����2�vM�}8�"��d����־=3�Fl:!U�A�r!g��=hUn�6ʩi�,�$>i&���I��BOL с�ؕ�
t1�M�4)��8hW.���N�JO���8��>z;��ʏ��Ds��ƕ|�5BФ���)����N�ǟ�z�m��$v�d�����:ò�@�e fJM%Q�����&C���aDv[���n-���0�6�����s�������|�z�Mh��]�������Fu�$��d�ZX��H�=�i[�̿�Ae�f����5��Ú3#������^?!������evUr������}��T�~�RA
�j����m���{e����켈�3�`d�b�#�ޡ��� ��:!J>,��X�P�-���8Wg�t56z�tZv�MsN�P��'�?N ,��*٩\B�>,�ž-w]��S)����`�8���:�ix�ȥZ����;�[H�^�� up�ʎ�t'=?.9��g�L�
����&5�IY�s[u	����y�P>��\� �O!�+�e�za-8*�D���yŻ�aQ�pD���kI��V�H�ɻ)`�~����r$�mP|{����!1��'Mۀ���� �����4�7�'�7C�S�R�հT7U�z{6ꑖ��qG9��,HUI�Ɨ�^5l� �����z����r�Z^��K�,Tp��4��	��]%�;� ����^ʋ~r��;��|�ۤ0�*Nb腺5��d'��u�i� nM��˦m6��\�$�qk��5(X��7B��,�s����0����3�=ӓ��既>����*�P�\����f.\���k�\�����Mč��ji���Qv=�71ж��Cx�៝�n�鬿�Z�h�T<���ϻՀ�,db��bH�)z�ߟ���!�t�����p�m�r��8%�u(��S.з��NKz"�Y��Pt�M�wEF��̄�����g^�ڑ��r�<�i!:G�R��� ���N�chQ�;�[pKVH^�SJ�E�񹼙NK�荓&���� #���2&�)��O���[Q\S��c�6���i���l����໮*���l&nL_�;�;dڍ��/.H��} �^r"	�7��	q�W?�!Z��I����GX����H'@�p�&4)�-@��A)�"]n�n� (2�� Z�UDTۃ7�N�hJUb1�� �Q���E�8�|�?��IR��Xb�5�Fzn���0Ns-����������B�(d����X,�5x�y�E2�&j�4S��e���s9�:�p�X3n��n�p�ǅr��!���0��3���/F��d%{{�δ��E�~����
<.o��� ����4����Lβ6��Ǥ��F�Ç?<G9���Z��֪��]�Ba�u���2}�>��Z���W�S�YT����~�����\��s�����壗�t�<ro�X���1��[�����ݑƨ4y"�n����Ҥ5�:����TG�^��A�z跸��.+�؇T �V�3��T,�H�n?����śLD�Jgq}b��e�[�����Gs��=�|ီ�X#iZHm;���)ĸ�i.6L��q&i�e����_���.O��lΖ��@�EF�xyc�e���$���"g��:�&|��`oȯGK��4�#S�X0c�0�"�2�*升f�g�.�2��!W�p�uh?���7����ZaD�e�z�eFQ�,�m!����f�n��eT��G��#'wr��?0�����
 �ѽ��Y�3h�8����~w�@!t�0��d#ެ�"�Y�t��$�Ҕ<)8�E[^"Ԋ2S�~/C��x�,uD��)�b\J�t�L���q4��gn��KD�1��|@ ��a�V��R�*�UWU�#e��g���
uL��Pξ���C�֓��󪖿����9��*�Ӧ��"H�����ԸFp���$rm�ȋ	���_a�E�.��0��]�c�&g��C�*`���$t�ݦ���������N�����J��+���X��[�k���������#֐#�ԒO^�E)1M�ny���n�]~�t�����;������f��;u�T�O~�;Ʊe�b�8*�\z�Z�h�rN�{��Sq���p�F��ݞŐ1&hF�jϲd�йD��Ȣ��F�
��J���R��Jo�<�>�ץ|i|��=ctV�vz��U���5`4��K2�SJyM�\�ռ�[�z ����h�y@��BW�^�&�"�c�;��I�I���x��8��Gsڒ�1�T�ì.�_.�0�akQH}��IK�b
F�I"��dꡱW�3����@����/��ͱ�<i,�xܵ���H�P��Å7�[K��,�[(�'1n��9�DCU^������%���/<�ذ/o�rB�Zz�c_t`��Y��~BN�D��A�&VP� �Ȋ�f�=7(.������J'��p#�\(�D��T�ȹ-��鼜���p�)Ӻ��p@��E2iR��(Kt��	8��}�_��~�(6e����>�� P) s7\��B=�c���po�41�϶I@�/tJ�Q�L�ep�tb���\�(���a�T
`�����7���l�ƶwU��C��˭ �QL~h;`��y�[K�)��B��v^���h|B�C�=�8���+����l�cjume��uM�q�u��1����^l�ԣ�xxzv%�--�a�凜دlVD�e�s�U����#	�J-�Na��$wT�Z�fqN����U7pD�*\B�0kZ"��'����kq&��e��x�U�P*fqR.������װxM�.(�d��4��.�}2�WZ�r&lY�d�2��{�!>�8�q<W���a����=G�2���t�DSg{�C]��t6P���(O��*�c�ݚ��ya8�I�)��9=�`'�����/r���~�<�2����\�tI���e��t�{�H
�L�as?�����?j�(��J |���c�]�,Q1r�`"�����v��8q,]����V�֙1�nl�w#�<!��d=#���Q7�$�,�b� $y��[��D�B��j ��Pذ,�څn��(H�)Wp�8�Զ��N
���Y�;n߹�,������bkDƐ�����w�6z���l)��Z��Nb6�����z���Y؍���S�]/e�������lX���&�� ���[����S����5�q�zOj��_4�gf��~V9|#/Iz,���`�J�,v$ǮD��������l��ƍ�2�==ֵٺ����Tf;`�$���~�Z3>���!��^b���.�� BvP���F�H�8VT��R�\fj�Ml��o�O�;{`��6n��6�`e�b%����l�����$>'�/ֳe��w��}�ga],6U�t����t$N��,�-~���f�,O�*T݅B~�{� �qw�e~S$HB�uUp`ï8��:����>�����lC"��JĔpZ���-[?���`�L3ӤA_q&0�Yb�u����زQH\��O�'%+�?�z�F�8�� 1`tzŖ\�a��p�l�f��隣Hԣ��D'z�2���a$٢|�W-���Q1�eM���&W|ڛ��4�4�wh'bLĎ�Rp*��������l9��H��cƒ%m^�1L VL���P���5Y0��+�T���/c�	�>%p7�;.��K��f$��\x�"Y۟�p*bio�@A������zu���@0� 	AÞ��6? ����.k�X�ǰ����3��<Q(,|�l��̀��o�QtX�XL��V��d�gu��P���������z�R�w��$�?M������)��vB����q��C��|��n��o������a�O��'�Z�;*�d}z�b�u�zԇּ.!����ou��',Ƙ�\p�M�r<��%�Ȋ���RM NF���eb��(h�w�B�F^�Մ���u��^���>��-�<�F:���R�+F�;J����ccn��%p�CHy^�J\�3���������D&���{�[��'S�D&�O )�Z0\�`Ŵ�˫6���i]�R�'a�ߎ�[U*b;2laS�_v�2;_���O�HX�: ��"��b��F�qH���Q���4+�J+�XW@��)T'��	�K�.4dꊌ��";N�A��])(�`�2�5OaD��7_vc�0b�@/ ��������l֭yI���X���AX�n!�0	�N���������B	-d(���"�53�W�`+0�C����Ō�P.��n:����c�7���C�M�y!¯0F�����F 1���{�ח��Y�7�'U�<�S���xf��
E�T���̚�I���
����H��Â�=����}������+�]�����E��ˆL��'w����S�d�/N�~��f�r�|�n|��(+�^��t�r�(�ݒz�H�F�I����8�����_ׂs�<5˓��N0���B&^�Lx��6��N��+p)�ϔNV�7��V�"�kn:?[�o/���@�L_Y"J�0�bЦ��,��R� s��0�׶4�i=UX>D7Z�w�y����C�P��6?���\� [u��_w�.*�Hl	7���q�FY�y�����|$���"�@:˶|�;�ocK�1M�~x�X�3q0�
�2��h���R������R���+h�A%�.��7'���`.D'���bC�a)Q�*m��v�0�5��q�Z�TJ`�G|r�#"�'r-�	0u���K�
{o3��gvYX�:h*�o���~��C@�	:�KNP�:Qއ�]<�te=���Y)t4mE�
ԥ�L���l��*9,�1��p��]�J������"���&��1��@�6��T�V�B�Ji�p�g�]T�B��2�L6.nι����6X��"����-H_��Tӡ�"�-�ࠍոa���R�nm�&	�V$���@P\.�� 𷜰c�<��f�i��P5�$9����I�I���}����1o���ܓ;����t���i�>�Bx��>�m��͢E��ᩳ��16n��ɂȱ�U;Җݗ6��f�#_�vI���Ѱ~��D��9����\4<�ZYnr)�`���//V�A8�8I_���h#�OjJ�u��HC�=a�F�4G�= h����Suo�>���|��<�ؐV�W��?V��MA�4�s�2��JT��pU�[�&h�Rh�@~�B��a�ot�]r����DM/�lOSx��6�S	�G�V~=Tژ¬�P.�r�a��}�N�f-�
��>"��Id%4�W���3����@X��b<͌�iC�.xw��������P�nfàQ	֨*�`�d,�����ͤ�9UG�UU��
�� λ���o<���/
�m�%Z���Mc�J��5j���A1�<P �����f╭(��ٛ�����e��K'p^��\á�腞�KD-��ļ��G�H	���=Y�hc�T��{�2� z���C���ʙ�G}��'^�(�+V��Q�>)݉ .?sR��Ͻ%0�>�ܫY�4��%��\�x����lVH���ܪO���QN�Ú�\�
��ȵ����AlxU]�Z�$̱ �Y�~c6ex\F�4��K��ӧ��;v9���t.�M7�8���1e�݆.�l)�j�߂�0Ĭ�,�������_�x(�Xz��-C��*�3�J��V?
R�ΫͰf��#$l��N<�J�_�2��h�fl3h��C�	�D�3�BP]�Z�`�b,��kl���.xq�PEZ�R�N��,ȡ8�İ�F.#e��-cR��t���W�gu&Gkd�~�҈>��q�މ��Լ�q<�TT2`Et ��gJC ���ϸ�P[~�(j��*i���uR�yN�&��V�����O`���>/�#��Y��<3��?!���WIV�+e<)��Y@�'7�
�u�L���?�@��v�j�RB(M[ �1��8L"Ql�b`�̦�
vj�8,Vͫ�$M���tE����lp�I�7h!x=ޞi�l��ʟ�\�=�*$�}� =z�?�B�� G���c�� �W��)��8������Nz�~�ك']��4%ʮ����&�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�ڜ4�y^�*г�j���&|f~o,KN��xslЗH�S��ޣaQ(��OU8p��ӳ�ę^�|�ΡZ���%C�A�R�n�X���<���.���R��_@n^��g���+�¦���,t�_�_��t��T�(�gџ�l�0����G�KA�����tf,�8��'��J}����/rĞA�ɢ��`��F�qX�ߌ�����a����:��дd��-��q��!���7'c����~ZX�ox���\b� ���y�1Mfߖ�E2Gb.�S��^'��I�d�0�s�fz�={���|Y@�.����su@��_7ᢈ^.�)W�{p� �H�>��~νU��M�ز�����
�y�Q��]�����U�-j|@�'[vv&&�/&��΂|�S8G}(;�^f�&�<4�~]��X/�\�4�Iށέm�<�	�▴�����G������X͎0	��h�ٺ)��An�l�jǲz0��{Ո�᫶��S�� �� 9D�1A؋=��c�lR����U<��-�e�
��Im�g95K�^���(��jc��K����52�� n��e����z�1��8K|�j�|��;s|/�������`�D��K	�p+	�THˀ`�o�FRD+'��
8i��1V��05�Q��wExu��O��VGc�Y��leykD9|l��[���0^�mO��x���I�k�����T��ݺ|Eo�E0~���x�;H�WH
��i��������EC��
����v��(d�i������F�7$�z�$��Iy�,��;M=<� ;�$��qGU���n�L� �μ;,���ѧⰾ�]���t��[���1����>V`��y�J�^�}^�����e�kbt��'����ඟ>�u��>٤X^8%H
��ɭ����]�&�4�,Ԙ�r��p�$�:��$ˮ����r�� c}~9�Ǉ���c:2��|�Ll���[r˔�����٫،���,}܃�a�%"�5l�f9܃�&�%
���AO&�la	-�8��3�D�5�;;'�<���1<��rV )4���\H�i��y Z;І��ڽn���L�e�D�V;�H4]m����)�9˯բm�a����R�sd��J����p�\֢�h�E�r�A�Sނ���-F���">��_�A^vӀ���W��36���sM��H��~Cmh1)V��%��w�ɮ����Hqw�nۣ@m�7rVE0�;��h�zF�饋�U��Q���ѥ�(	�������.�.}@V�2{5��X��B4S��/
Q��T�}/B~4
O��NRjWף�ؤ{�
Yg�o}�?�����J�d#�	�r�KWܑ�\j*���4h1��D�^�d喂	�����	N�6��L=��C�1�3�vM	�XYg��X�ʖ�����ᩣ�w�г�s��\M�˹��GC�k����]���J��%�&�2��==�ժl�Q	hr��SZ������둷i������F@�r�st�%C��<�)#3j��������G����N5C�P=~�"lIZXM�|o�q�^�e8=u�&X��?�әI�t�0�k�f��*Ms��t��&���De#8!4VW�����H�!'�s$����~��v�O%lM{�Ǝ���ұ��%I�6��q^���gԻE�\Mk�*?���+6�'�!S���?-�?>2 �a����4�ǜU#>'��-,��y�n�=��0!���4����E�$3��#l]����'N?��F"/���9RGt�,N�ܪpE��s����朿8���(y�떦�u�`4�:-�W�Ƶ@�_�9�`���56zo��ĸ�B���#�G�ûDz=�ԇH�,���>��Z�@�B[4����T����G/���> ��k��UI��gl�˅� �&i���*=����hAr=y.gB)���wzW���i��6�4�	;&r�S�C�D������T�sLS�'3��P�ݞ���C7�"t���\T0�Uv��^f�P��}u�*��2A��>k���/�������_�2��f�|ex�q���(���P�� +[���}%��A�!��c0TI?c����"њ�L����y��F��w�hu���^�!�H�^�yc�2����"���O��'�d^6�*C�tp	я�j���Y�v˫h�e0���'���ە�{'�n;�` 2�z�nJ2���7R� �v�(�n�pJBT�W��V84i_~�e�,n*⪣w'd$r���l�;L���_j�dzб">�����9��e��T)l:h��d�H��������A�'�ۭ9�~�w%5���<�b	������Rq�%��6���w�� �H9�ػj
��Ơe�|�$����0��.1�0 p%qEw0���e���z�JQ[g��k����߿�4������n�H˩zMZb�� ��WG,+�+��b�����df-� ��v��X�Y��ųxb\���,�y?	2f�W9E=�.!��)�y�t���(s����~{2�|d��.���,@�0�_���I>�)]d{g� ��ͩ��I��U��ؖcL���O�����-y��j������,�U�<�5�'F�|&qY�/ѭ����1�(וGHI��h2��R�<�u]�8/.�e4�f�9l����D	��FE9<9e��ci2�;�E�s��A��A�<	�WNާf��Z�ް����*x���!{��X���;�|�)�P�>�Q㜑Eh<"�5%���1i�������d��?)��I��B�T�J,�[+�ؽ�����u���5��">�X_�Jt�d� M�\re�#V}��@�ŕ�Ηgcќ]-��l��(p�7q�2�(Ѥ�!I��P6]R(jr����_��1q/p�� �CC�]��a�KՖLa�3����&��_../��iX��y��_�K��R�Zܤ��\�$N%��f�X>��}�����I[ʲ����#H%x�3s�d˟�i��ƀF��/��)<eħ��c���1-�Vy���4��Q��������k����G��7���}(�Lfsw����S�4���5⫒�*N�G�N����f��Kl�xLK�AQ#���ca��߳�	8�u9lY.�R[o���0Κ�V��Z��N�RAN����@Ck4��0ʍ��;R�-�_�^K/g��褒�[^/��,M�J�Xt���>�g*�~lzT�#>�� �xA[�i��t�q�P�*�V���n�!/+�\A�] ��o$�x��	8e�i���W���A�K�(����h0��h�玀m7�X,����+��6��e(M�AM�Vx��[I�����c�����T=��O��Cp��"M4϶�Psk��P8���:�b�Z3�!ܼ�5�:��ϳɽ�0]o!�)!`�2��X�jP�7�v`c�U��na}�M���6��b��ǩ�r��!�{�x�vi|���߄���6N	�$Hw�~�6a���u�=x�ƅS��9�J>�[�- \�F����M rt�?�uh��	�Y�[����8��/z�l��m54L�v�/�he���D%�"�Y�e��.IJ��˛57�@� $Q��;�v+mp��m��n�'J,l��۷s�-)U	%=ې�\#���Ha_�,��.4� +�� �O��5.\�I���X!vқ"�s~�Jx.��y��s:���ù�2��T�v�f�[X�R��Ek��I�&;Zq����jH�z���dԳz�i����Д���1ipb̵C��C0*���x�T�b�VHo�Zn���w�\���O*���Bw:<��O�]��TJO���@wա�|�9��Ґ���Q����M�6E8)
I9��(�sz��-�?�1\Qm����#�VڢS�+��,K���rR�)��|p��T�8�
iهÒ+���$|�}':<L���fF��H84��]�!����)Qڒ��sz�U�?�%�*�:<O����߱�`��Ւ�a�����e��C����P�$��߾_䝖71���p�{x�k^z�H*�؞�NGr~|W�]r"F��;����'������
��R��J{�1��F}\�+)I�X��w[���IA�M��=x���l屡ΤT�m$]��^��C��ź�2o�$��-8�h�j՝m���2В�?24>�M,G#0��n��`6�_�_�KvI��T���u�fG�gL$�\�	.�آ�!9^A�?�uTUAQ��q�q����4~���R!hN�fox�ir��A����^���e����GR�ߥo��ө ;M�N �1=M�	I��թ�����w-'͓�h����y�b\�!C��e�L�I���|��ަ4G$�T�0}1�b<����<�t��e���-A�,Io��僴����@��5�v��J*C2���a'nbNoYv-�[���xwŒ���b��A�[�_��(/�c:)dN�X4H�����(UI�G`Hp�z�,4c�%���<��8��t��=�7�~i�p�� Y�&?axՙʿ����_=*�?ul1q!%�#?V����P;ʇ��/�5��es{�mJ$�DnE�7?�Q�Ji �.�s�|�#�鲄+#$4�ɻ�.���ϕ;@~���M��"��6�A�f��B�y�ˈ�*̄~7�qc*.���ǯ�( �`�yy�o��F�P�{�$"J�;��a�{����OF�j�6��~��2���E��wx�jo�[w���v-��0� �|2C:���rD�E��i�Ԍ�D�����/�W%"ѣ�,��AYA�KO�ʌK�Q1���"!|��v�yGFY(g�6�x+f�S���H3�14+p�)��
�:��cX%��@��M��3#i������D�6�7�N��"@��e@���g�1�:�ֿ{�5�6�����o����H�H(hH��n���D���@HAK�$��������<�/�9�I xU���`���k�Һ�4rņ#�9e���N��4��������Y�ē�(�(���l��Ag2N�ƪ3[��`�@/ϨZ��I�SO��<e �8�Jpr�N6u6ֶ�V�� �{�8��:�Z�ۄ��F��t�ub�T:�
�G��DF�NKO�Q����
��gM�V��~�\���}~8�Og�WTT	H�:Z��up)�ZU�3	\ʮV�$�͘U��.4�i�)�;n랕���z��yE���pǶ� �z������5A">�F�6RF���U���� ��]ٲ_���$���� �3��!�~�.�<��;�Բ\!i4�`����z�j�*"�8���W��n�Mw%6�����x��W��	��{����x_l��t΄&l�6h~�CH�ЂgH�R��k�1�:��D�ا��4ɜ�5ī]#q��q�P�������"f��F���>�;wo]�Չ"��/�� .�N�7
J�3�\��e%OD{��)
���#WD��e��R7�,�<�'�\I��SI�����7D���髝�քyO��~��wu�M�q'"�V�i��khb���뜻9��y�ӆփJ�����]�2A��Ǎ���������p��=��O�My��H�[DO��ݮ��� ����V�Ro�3<R\���W�L��ڣ������ ⫇R?���,�d�rh��Bͅ���X���oG5�[�0$��y��0:w�S�w��Qp>�>�2)b���Gg>Iy�u��~�#K��[�aqJS��nT��O�n��@7���7��`o�_>�`SO���h���@d�)�-ފ�n�C^`m+R�����TQ��f�r�����-Y%l�-����\�}-� �պ*��(�̄_[k�$=M۷5ҡ�2S[v�Y�G�dR��2�>�q��MD��bƦ��X��d�n~)�.���!�<&a�ӳ�f2~��-̼Y:Zn���S��d���ȟWa]Ȇ��iB`޻���@�1������uޕ�U��8o��l�����Z���3ĸ"�p��ꝕF��ZyUg��f���o�����Y"�:��M�4Z:���|(��_4o{��t�4]���� �~I�2
܋||v~9!I�a�]�P'v֩77ǉ@I�9}�����|�
Q�#��p$��ֽ�8�{hC�N�v�<�0��Ѷ�d#��.��su�847���Xʦ>[r�0�4�Ue-�k �!J���Q5k�����Z�&�Z�[�wHׯ�-X���Q����Ü�Z;����[
�pS�4����B�)���h5	�V�r�v,���]��vj�tUI{>E����X�����u�a���W�̋"�:�V��>A�#lM�PL!o<7�-�9�*��/��&���˜`�e>����춘���1��*ł��Я7��ӝ0�eq�w*��g7"�6�yd?���W�z'�W�j	�a*�Ʒ	M�������Dg�?HIq?U��Gӻ��DMm�~��g�"3l'��Ȩ�����.?����O�<�4	��U'A'v��,>�y_�������7��I�#4���������	����jR���]�IFYWb��hsR�XV����a��ߚs�3�U˛�o
��~��L#�`��-�M��~����M�p>�訃
�USzF5��{��B2(m#]��n�zt�}�_�������`j�վB�ŧ=�^TN��~s���	[���ďB��t���b( %e�i0A*t�o���Air.��O�w��U��W���i����kw�;=�(�JǯC��~Dhb��s���A���D'j�NP���8FC�8��PG�n��T��_�o,^S��P�Gu�_ ���AR���Յ��m�^8�]�>f�vT�A�S�Nx��1�}�6���S�G[1����%{����Ej�b�I��݈�񡆒=c�U��=r��N�u���^������l��W1�T���"�<�&0��ޑ�^�D�C|;=p`Ѫ���z��2�Y���?ҁ08w����	�?쯅r��ƥE��wq�q�yJ	������ ���z+��O�Jy��W�zcV/�H_U�4���yV�w���$����Sjl�B�ט�_�*�d1�B���e�U|�9O-�4�lQ.��U1�,"݅���|;d'��9~�~���L���3^H�J*�|ƀ�'���؍���� � �\���R��#���re5Ę$H'�.�.h\ �`&En�겒�
O��zl9�[��[�¶��#������J[�Ʋ�H�h�z��Q�vI����W+�H������e��;�R̷��X):�rUb��ܹy6��faikE�iN.���4�����B��s�������{	�K|�.��-q�@+�)_�6׈`<�)T%${�F� E�U�@�ˌ��U̓����u���r���1yuZ��_χ�>�U0��>�']HE&h(d/�[���-��VDG����*��>�<6B�]��/Q4��l�В��F��	Z|�}x<P� �ZF�8����c���X�	��N"s���Z����D3��5��7iV{-��8�_ǳ���gq9�H�o�sۚh��5������4���<����N������T��JJ�b|+��_��J�4/R�,���U�r�J+��w�K\�>��Z����`Ō�|�>b?�$�k(��Bq�u2�3��7�I6487!��~��_A��q�iɶW��C���X�K�c�L6��:pf��,���/�9�Xߛ2��t�Ke�������x\� %h��fOmOXU�h}�r�Μ�I�����Oc%[D���,�{�O�`/���A����������|�c=��%?0-��@��|��Q�
}��3��$��Z&˱�D(��	�}�Nf
��9��ً�P
h���.*E�y�%Ď���of�ԏK~ǂx�ݡ�xfS��[�a�1j����8�NOI���=^�=���!��$ӷ忔�RSñ��������S�Q�R-�4_3�^��g�W�[�W�8w�,��cˏ�It��]�5�g�%l16չ�"B�wN�A�C\��t�i�h� �L��E�"�/��?A+c�,�����k� �$	Α6Y��ex� FK���)(Q;��ѭ������m�kD,�G�� 6č�(d�M����ʍo����M2c \��EW;����Zd8�ĺύm�P*|��x:�@灔���3R����џ�1i�ϊ��4t!>��`h�U����j�ڿ܍��LQ�n8��M���6qXW�z�J����C�{����m���h�1�[Ss6�5	�O(H�g�g�5{���1z�Ã�n�)�	�.���w]8ML�&Qސ�ӵ��I"��M���w�M˰I�]��,"R0�/�`.�S�7��h��BdO����>pI��L�DSme��7���<�E�1+���e;E~ҡEOD�pc�����͵�^��L\���B.<"V��\�G��b�2f�1��Q�`��r���$m�����J�\c��<��G�p�+=�yd�i�]Cp���2������~!�%�RD��3�����5�+������柟 �r  �R�淡9�d4��'�'�B���z����#�� |�[�0��y��:,���tQek>k��9���͂g{��y��3�$K.��V��SkTT�>D܌��_���W�7B#Y`ıSR�F�|��e��))�5�wV��zS�w[��u�i\���Կ\',�Z�&����H�s!z�[{�=2ߌU��+mu�M����Yv�bm̾7�U�X�贡�*(b�5�Zy}�f��E��!.�(,�g���r=��Hsb���iN{0��|"U0.�pf��,@��_�2�Ǩ�)��{i* L�o�'93��2U���!=��mX��!à�My|���F��4�U�+��'Ģ�&��/��J��°⦌�G�~~��u�o�<�]'��/,�a4�B����$��2	Z�Ф<�Gjᡛ��96����J3��`	���N�ہJ�Z#o_��y#�����({�d1��)$�::�Χܑ��y�G�h���5���oF���:����\�D��܂�?��J�k�+�=���o&�O�쏛SK�s�+� 0u�#J�*��>��\pԁ��62�\9O���>�esB�=���w(���q��Z2_���^J*I6�k6[��(`6�e��_U�q-mh��onC���K���L���!U9�dV\]I�/eI�XF�+��K�7���"��o9\�5�%Zf��X�s}J����I�<�}f���{%m�Ij?����������e�����g	�ĥ\�c�ţ���-�O�hm��Q��1�����oٚ)�v4�:����}��f�Х� Lh�2C��>���*��ڳL��œf��_KESHxJ������-&�a�H���8�SV���Đ�:���d�XR��>��R?��cޓէ�/��PO�����&,|�+w�}���W�噰��:����L	}ٱH��b�H��R=�3� Y�i�V��5��^M�}��\�ܮ�cӰ'⥟�k���l-k��Gv{�7079�O�4�x(�k��kv�R�F�����|���E	ͥ��gx������
 �ig�ҏ���l�eEB
�|��޶�h�r�����7݂'��ރBu,�CyMv�Y�$�H-q�~��T/��%@��ǡ�,�Q����P�VL4���3�cD�-p��[�>O.�˒1JR���֕�ԓ�4�'��k���b��ݓT��5���LlӗY!X��D%�B��j&�����Vr�M4r	��ѝ�::�l�����t�r�dA|%4~r�.�����":�㐟5��LE'#�T���-�����2J��J�ٳ���̀as�p"�� �9��&�����8�Oߘ
a�+��1�3��M�n�};��<j����+�B &`���H�5�O;)�,�S���'�L����V	Q�HM��m�oIڂ�=9Df�������UE�lc��c���F���^�\p0�&�s�l�3�S�j�����Ț�{O���A�A��EU��0$ڊ,'��c3��;��I�em�֖VJ�G�w_Kɇ����3�ajt��w��?���)V��;�&h�"ʇ�H��n��Q'V]�*�3(�4��"�*��#�}ǘ�+���c&�U8�Bli�Zk�
������}�O�Bw��O��.N���W0"����
���o6;�`�B�ɨd<���L�W5Y7\�����<�eiF1^����)d���	ι����կ+�����!m1��<vF9�q�[��jB#�egQ,�a�ᣜ�Ќ����Sf֥� i�x�� �;]�3�y���� &�4D�C�="��ž_	�k�r=QS�2{���֥���&�? x�qNR@�y�r-"_���;��z#,>A��)?�G�,�^���9��z�P��"���MZQ
̕��qR��^�+�=��&񣭇�~j�"���x֘k��y�c)s#t���&U:k���8�G�W��Ͷe!`�$s}��.}��iI~�K�MT�<��y߀�(��^�7�5�q׻�� ]\��Y�M�'܋�-�d��'#�j�K���?����:K���"4QRUTϤ'�0j, ��yas�����	Yu��(4�/o�F�M�}�å�s��lt�����FKv���R@E6ۅ��#���|�s�p��װC�1�/����$�;����`���-��N��7��V;�2v�誳���z�mn�=��B4��#����z6hɇa����ŏD�=��B�N��T� C�@��������?��6|��d)� g*Si���*6�j���A�U.oD�����W��W9��i}��-7	;?C���4C_��D*����\��K�%�p',P���XC��Eț���p]�T��8O+^ʓPڃ8u'\A�q3A�	��2���G��p� ��x�G��ճ�ջxw���ybx�����[�JF���%���z���ܺ�I�<��G��s[���&��wL��ӖЊuI�^�i�|��Rs�:���"Im���<R��.�^�yC�{p�N��������Y����@�0������������y��g2�y9�ݳşJ��^�ZȨ����/���G��J;hW %1Vq��_����{1Gw�%$K���~�l	g���_d��d�ٱ�M���?9�2���?lS�hăt��"��GK��~�$':��9��~���NО�u��b���l�Ƃt��a����px ˎQ�ŋc�/��$e7'k$��E�	Z�.*�� �t�E�b]����Azn~J[ ���DD#��)����ϾU 7�H1�HD��z�>߸P��0��+�(���c���=!ǽqt�y��!XXRס�×bU�����yx��f㫞E���.�����M��M���s�.���{�k�|�9(.��Zoް@�Ғ_��b�b��)�c�{tM� Y��B��}�U�Cs�\�Ց���]%y7�F�a`�À��U�p� �'_�9&���/*&̰RHY��ɭG__�e���<8f]"��/�E�4pSځ�������	ܭJ�?ƨ<R���Δ���m<�eF���o�	s�
N�`�s(Z���$5�6'�9�9{o&b��m�uF��i;%�����-�h�I�5��n��R���ֹ�����������w�����J�?%+Q�ս������"�6�E�n8s�{l��X�J꼯��R\K�i�d�����)e���5�֏����()��q��2�3����I1&6�W�=��� m_��q�v��EC�<��K.�JL���<ղ���8<�/���X�M��JK����yݝ��R\C$%�zfm�XW�2}E�{�P��I�!������z%ݵ���j�}Ŋ��IY�<�X���u��R�E�Ĵ׫{
p��TJ���b���1���p�1���:z�0���,�~��~��C]��+F)6u�4X$�����<�-�8��
�xg��,�a��F�m+Y�Xږ�w�F�5>�A�a��m�#�P��.��XumT�����Рs&��`�Ƭ����n���/6hmA�E���-�!�5>�#+2i�Υ�bb���q�L"(2�A�Y���zӠ2-;m��f,�
����6XS�(x5BM�A���oi؂���c� :�Y�����O�n�ƭ�ϡP�?+������ߌ�� �3��D����ŋ�Ϟ{��{L�!R�`� ʩ�f�j�yܡ�؁���nL�"M@�6�6��d<��\��RYx{�I���|�b���6���#D�H���g������1��%���"f�>:�]L�}��;�']ȵ_�"i�Y_a��pc�D��]�%B"�A/�-.2X7��1���j�p�OM��Rs֛�DgGe2�27��<���E-P�\��1�5�D	]��4[R�-�c�N�V�`2�V۳P�ZVUĪ�[u�b>�m�E���c�� �S��bD�{zF�0��2Sr�0�p��=����V��q����?�Fjc)Ɋ�;���NRXO�3E����Ŋ�4}���&���4p( ��>R(�D�5"�dH�?�L��V
g��P�k��8(��U�0-߃y��:�����X<Q�ѿ>7������rgn�y�Ǿ��K���}�Sa�TL���.���iL�Ο7�|`�=��U�S��[�͚ĥ�d�KW-�n��`��Ʌ���QVzR�[�w���}-��_��.L��.����&kd��,��=k�<�̭��k�^��^5[��T�?M�Y|�m_�[s���;�(*y�-̖�@x6��T{ng��7�F�J�I&�`y�J�k2�T�(aʼ"�n��&S����Ԛ��Fk��@�i˻��Q�}@��+p+d��m_�O#ց���մr푬�Z+e�����"������o��ZeЮglOf_E�o�$�We�"o�ǇVҰ4�C��O�/|����&�o$`�t������ �BIUr
%U�|�p�!��rJ�m$֒6�7�e�I𖯎�њ�7���	�#Bbo$id֦k��=�w��w�0w��?%=#SD��+�uk�94@����Y�>���0E2�U����3!S)���)k�m��O�o�'���Σ���XfXV1�:?�{9�L��B?� ����" ���=�9�l&�/���C�<}�O���a�0-����3�u�L*;�@<�h��f��	�[ ����H��u�;Ǟ����j�E��L]�sB��Vg�3Hk	�mדU� 5�9��
�$�6���%�8��uC�Ux�$����D�p}A;�D���M���/�S5�����]�~�k��Z+mA�؀#4f�����g��=u��Y�粆m?��Vh��U<��%>��_S���٦��7����V��;��h-Y��@S!���!Qpf���_(�=U�@ ô���}�����r�����3P�B
}�����
pq��ͧ}��BկeO���Ni��W���{ʦ
��o�8��'-�dZ���`�W���\A`��Ȏ��C<1���d��d)	��B��gb�-%���^��1;��v�� ����z6�����c�`	�z�-�*������������:BӐ~�3]��v�F��@�&���K�=  ۪cF	?�#r[�vS��]�O*I�O�f��!�*a��\@�r�rKG׼�2��kJ#���	���%�����=ė$��ݙP�oK����Z� �̳��q0��^��Y=Lu&E���C��5w��JVk���A"s���t��&s�ۤ�8�f�W����f!>�MsN7��nŇf��0M����	��<��-1�q5+2��M��M���:zI��>B��'�Ş�������?�ft��gǋ\7*4)IGU2�8'��},^+yJT��nS�o��i��4�eq�$z���+��\��"�����_�Fy����HsR=R�#p܁Hy����s�'��uCK���)��~0��H�l��`v�-�]���ε��������ȣ�y�zf�ٛ^�BRX�#}�O�:&sz�JЇß����(��RB\ҧ];Tnͣ�O���iӽ��H��*�����t E��i$(�*����23�A��Q.�V���u-�W9�i����D;]+��jk�C���D�;$��#��������'��P
ޜ�6�@C.�������b=Tǈ_��&^s"P��7uD-��Ar!���uI����X:��^�}�T �ڻ��s]nx�hB����V��s<.[Q�k���%�t���:I����%O��Z�.�����]���n�u���^�,�����/���,"'MҫF��}=^�C��'p�����Ҹ��Y�ga�_ڹ0X����d�_�\������a!��yݑ��J)�ͩ�	�;�/���+J��W;�VOsT_u�����&Gw�V$$�Tu�sƕl'�$��|�_�dQPj�ـz�up@9o�$�8��lq.#�Y��?�rݥ?ƜK�'�968~ :3l�`�S�� ��7Ơ#Y���uح������ �x��R�&ɨeU�$hs ��.�8� ���E�2����}oըz���[�7����C��۾3γ��H�t�z�ߖ�ŌζG+e��,��	�[����A-��X6�Y�<�kb�N��8�>yV�
f�� E��.؞���U��%<�b@�ss���{)/W|;qE.�Me�@K5�_�舀<�)t)�{�U e�`Ќ�FU-dܖ�Fq�&�ŭ��p��Iy����)�^LrUPO�^��'}��&�l�/�#����9�ߦ�G��1�#4�*<V�C] J�/%�4΂����f5�	zʝt <p:�zʂ�2@���`���9���u	�^N5>7�:+�Z�f ��l��bY�W�{M�̨X�&���z��1��h���#�h�5�{"����"k��\,��/~�n<�p��+GJ�Rs+/�-	ӂ�,�T/��L���S/��J+;���b\�ֈ�z��� Ŭ�@�^
��4���#@~(�q'`2��ɤx-I��6T 6A�k���_a��q�A/�w�C�h��xVSK�K�L8"&�Z��H�ֆ�/�5�X�]���K��S�1���#&\!q`%��Dfo��Xu.�}#Z����pI27���C��oM%{|��h���������ډ�"�������Tc]MeE�-�d��u�sQ���(��DQ����/&�I����}���f*)��Y�z٫��*�e����*eO�El��Qf�K���xÕ�"����a�u���8�x#�A���]����y�D3�����R8;ɱ�vf�q���8I�RM��_S��^%:g�S�{�,�X�,Ĝf˯	�t�e��U|g!�7lQb,���~���A�{��R=t�)��p�N�-��%�M/A!�҆LD9�I��O�/n���tα&2��Yo� � ��V�(>QO���A�	�����m�{�,"΀���p6�)�(���M�Ժ�r8�����}'c@��e=�'Y��z���9ϭ5JPJH������`;����L3r]\��1��Q͌Ϫ�Q�!�!^hR`�H���j��,ܭ"�l�OnX�M̨�6��旚W̩��_�{����+���t�{6���H��gr��� 1��$��c�-@��)l����]X�l�F�	�3�j��м"��c4�����=�]o�"r�/a.�W77�u�����R,O���^V���Ds# e��7�=�<.O��Q[&��g=�0��YD����03�9o_��*Þl�����\�V���g�bʖa�Q�j�q�Ş�⨃ߘ��+�6���<�`�����OHp�J=�	e��|�}[�(��R���I�����Q�Rd��3Ѷ����,gڗs햲��@' 7l�R4jC���dT�GK$�bڃ͚��n#�Č��K�0�� y�	:LtD��t�Q�o�>��9Y,��ݻg��?y!�i�S}�K'N�v��S��T����������<7b�3`��S�LS�l	�Yc/����dkg�-{9n[:q`��Å1�;��Q��gK�A��-�z��V)��zg���2�6�U�����̹�kY%���?5�+G�X�yTY�٩���Z�g䌢F�14���1q�L�]�GM�ns����Vw�&6���V�2�+һ4����n��S����ݐ�,q"���FiW�&�][)@$M|ͷ�cQ'��������|��v�Z7`}��;�"��\"���{fZ�gx�f��Ro�^���"{�U��M4�0����|�띣�Vo0�RtA���ˤ� ��I%��
��#|��!^a~)J�-֞�7\y�I�%�	U5HP�wX0��@�Q=�У x(���x����A	}�������kq�BB���A�
@�$�#��}��&B��Oc5N��WW� س�G
HmoL�6���_�d�B����W��\y�� 5��{�"14�M�BdT
	�D��׌�E���;S(�;1s��v������|��#������vG���.�b'��"����!�r"����c]䪣�ێ��|@&TtX�u�=8�٪���	w��r�{�S�J"����Ls����USy�G�y@"ʾr������,���#���AH1�]�b�4����3V$��P-�����Z�����߾qh:�^ҭ�=�<L&G����Q3��kF��ys�s��t#��&�Ҝ8�:�W=i�#�=!v��sS~��ĥ�ſ�j��0M*;%�V�ԀA��td�e�qmH�V�!��[M���rE�z0�'�e8� �M�.9)?�H�d&���h4a3VUj�$'� �,�w�y����|��#k¡��4��\c\�S���2t�� H���T��F��d�5��RV�)�[�;ܹ����s�5��g���13���o�:jۤ+�`C��-���!����=�� np!�vz��ӝFB�~�#���r�Iz�ey��El��j��O�BJ:���T���"`��:��~���Ҳ�̊�
} }6�i\,�*��j%-A�/�.EN�Q���{�WON�iS�6��� ;��Ả\�C5�D�Z?��)V�#��MR'��PB@$�n��Cf�t�1t�� �T�u%��^�ՓP0:u=�r�Gs�A����-콋�΃�)�ME��&��������x����(~��;���u[�¦�9U%���P���r I.��]�Y�I�o�f�mR�S��?ǖ�Xuu�A�^	�4����(<-Fͣd7"_���~�6�6�^%C��p���,���d�Ya���0�����"���UL��.���d[��{���R[Jaҋ���{Aw��E���
JќZWV]tV��u_���;fѤzw���$!A�ë9l_�܍/�w_:ۖd��j����m�9�I��p�Fl��M�2��w����W��9'P�9nrE~8���5��i8�ao���ɸ��a������x� !�0�'�L9\�^@�e�rf$�������.��V �zSE�3������XzĿ.[6�3�{�M� �k����NH�[*z<N���rÌ��+>(l�>V���z�ǓQ5���e)�Xn*U�t��b����p~�y���f��EL�.�"��ۆ�#ҍ�s@sS�'�,{a7�|s�#.���"�@��b_Q�+���u)��/{J�S �ս͘�>�w�Ue����駈^�Э2���@yͅ��e�Öy�U�#O��+'�Jp&�u�/ T���0G��XG�i�[�h�@.�<��]8X/]�4r�(�.���	�LP��?b<����C��j�ҭ*¤��-�B�	I��Nm�l�r�Z4�������9����_q{�������,��������3�hK
�5z� ���Z�N��2�M��˂M8��c�J	�+g�ҽe-O� 7-��A���GX�Q^7g�+Jc�ǯ�2�\!�!���ͤM�a���B$�l��[f	(?�q_�20�i�O��IG��6���y֖���G_��Iqލ�����C�°�XK�ILpѐ��v������/6��X7n�28K��i�i~���qU\Y�y%�w�f�̗X�ؼ}[KP�&�IjV���I�����%����d�����,�Z��U�i����[`�V2c� �}9�-ƍ�?�qC�Q�p��Oe4�|5���A�g�y�Kb��ң}7�fbW�Ǒ����)Zb×�VV*�ꖳ}dJ�Q�f��%�0���5@���VS�|�呉���bY<�Z=�Qľ@l��r��׾�ʄ���#`B�ˇd�'���>������^Pֲ���3:Z1��u	�q2��^�aH=�q�&����hљ�)�X�ak��^�C��s�&�tmc�&5Hlݫ�8�MiW������!@�Ys]��/��I7���{M4�Ў�����>=�o�q�M���*}���*M�ֲ���D3�'½�J_~ڸ�u?�&�����,�4��6U4)'���,���yAE���Z�ސ���4}���&���]%�|�I�L{T��A���F�l�ӿ2*R _��ei��󝎘ʇs�zy���n����
���ۮ/�`��8-���!d��{��X��ь�_z�����wB�G#�B�|�z*�A�P���؏$���r�B�<	�_4)T��� �H�z�0���T�����D�w G��ifcY*-���FA��`.O�6���7R�W��i]0®� ;�ٺlًC?-�D
2��k��픲Y�'N�P�5�8L�CpJ0�{�1�P�6T�	�/i^���P��[uv��Q]�A��ƪ��x���������3�X�Z���.����xW�Ū_���+i	Ը�wֶ몐���S����Č���r���/{c�a�@|P�r�G��;�8d#a���X�7|�Nm)�)tO�P����뎑ZA��̅hpqB�u^���=�6E&�8��fs�h��k�X��SIs��t}8�&E�}�.8�ȴW��À�3!P@sm�l���Y�~��]�MDC.����ە�N�v�q�B����:��\�M�q2�
y��`T��'e��ZdI��f�?���*``��9�4���UD��'�y�,�fyQ���;�����5 4�lR�6[��m�i����\B������F����R0e�u<��(����]s�3
����!�f���y>۾9`��S-����d�	g��"������0~z�v
�-"�B$��#��õ�ez&� �Q�׆�?�4��גB�C�o:T��C�0�7������ӏ�'r�&���Tf W��iv~)*&�a�f�A��._�����Gy�W)��im[D�&�;/��|�jCO`�D�r�{!������'�wP�tK�Hm�C��;ȋ���`T�2w?�3^��P�01u�O�a�
A�֪��~��-b�X����6�hO�����T�xgJ��o�h9��Ō][����\�%�JN�jC��a�I��0�7Ͼ�c�n���R��֩oﭖ�2u9P�^�}ȿ���B���ң�#�"9x�������N^��PC�epү͏�~���u�Y������0�,>���ɼq�}����W��i�,ݣ��J{�1�J/��>a�w��7��J+v^W�a�Vat�_�&Z��\�kf�wА�$;ѻ�ͫl����	pv_T�od�Oe��r�����9�S��(vlC�f�>6��;��7���n��'*:�9���~�$�>ݢ�eYtR��w���ry1��Y���?�`9� ��K�`�Sל��0e'�$zu���J�.
 yavE��:��^��z^c7[,,�4%ݲ�(z��i��E{��8
�H4�Wz��xߨÎ� _-+�O��0�ըǭ:�i�����XH�h���UbEs�
Syhf�d3E��.�n��Ҡ|�=2<��ֺs����.�{{I|� t.��_!
@�s_���RW)���{d�8 �N�25֌�U�>�L�!��a���)��/y'z��Q���p��U����L'O�&��y/���Bߤ�>lG�q��u�@��y�<(��]��/w�4`���L��x��	���/E<Bb�W΄����7�U�
��bf	c7^Nǀ���Z���~�䓝�)�a{_	���[��e�{�YxƑz����f�h��*5��D��%V�t���R��'�遍�g��f�J�d�+AXν�Ăz$X�&�"�^��k�H��aJ�����;�\;�D��U���žԩ����ƶ���a(Iqy��2�>h�醛I!�6�c�T:�p[_s �q����	�bC�)�1K�xL�	��,����\�(`/���Xю����<K�� ��p����\3w�%ڃ�f\�XGS�}50�@f�I������K%�v��t���m�������,]���_ ���W��I�pHc���T-���Yz^�"&Q����):ٖ�P�T�naz�%޾�7�`}���f�|��ky�����:����*w�糗ձ�p��f�
�K��VxX��*/���:qa�8<�8R *�P4��C4���΃|���3��c�R��:�E����1���o�R߽�_%�c^7yMg^����3�G�j�~,��Al�t�1�g�\gs"l�\��������A$��'ut��E���9�������q/��As?��ފ���ӂ�����=΃X#� Ɔ�r�%�4Q(I���t
�?�PO2m�_B,4,���_6vTc(VZ�M�Cl�!�f�cR����a(���,�Lӑ�KB��`ZP�ݮ���r}p�+RF3l���*�c�t��K9ԙ([!0b�`�|ȩ!6�j9W}��S�~��n�8�M^"~6c���}3�X���pR�{�����x��ڲ@�k_6�Cx�yH@�bg��/��� 1��#�KW������{����"]��R�؃��v����"m1�w31��-��9�]U�"�7/��.�
7�!��c��O������6�kDE0�eЕ�7��B<���#����y��߅�S.JD�o����!֋*!�lP��>���h����Vs1F�9��b�!�룃��U��l�\�}!�ϙ%�����=���n�p��0=�E���
���:����$w~ǸE����=͗R6�g3�^c�b����[I���:������ �Y�R
��ӧ5d�Ȱٱ?�4֖ͬ�_#��V�9�=0�"gyl�!:�L^��_SQ���>�mt��w��Mg�oys܋����K��ʈS�,Tj.��r��)�+�z7��@`�@*e�zS�������\�d}��-e�n�hr`���CC�`kQt6M�9+ʛS�-�PA���c�b-��(�~��*��&���zv,6>�"�k�7��["5�*v9g]�?YZW��7���R�%���"咽�����CnEL���1���&ȵ��(��2�q��	i�@��nq�S�!(�H|�ٷ��7�ii������@���Na�u_�jt�֟^Zȳ���/=�Z�	���"�4����h�Z��IgJ�Kf��@o�9)�u�X"M����?n4�d��m��|c����2�o� t�mW��N ���Iw�
C�&|�_.!p���h�7Wr�pd���ݦ*�KW�koז�6��͏@P�_�:�]3��C��ƺ�L��DC"��bN�
�@.׉e��ҁ&1"Dl����{�1B��҆��߼R�޾~i��|ohutg�;z�����M�KiYl�ͬ�o���j�+���9�r�xq���۫&�6�����!#Ɇ���e'8�NOc\�*����A�v�"��v��xx��n�eN[�M3�q`*�7�ʧ��LwI>i���� ��E���{��u,�������mj��%�:;����\Wc��+uo0:a)G�BF�s�Owt�C ��
g��Rc�s�n!-�2�m:��� ���vx��U�>������#��C�G��UeA�06D�$Y�>��i#��PZ��o
�������� ���z����d_u@%���2�9oVu|�=�6���Se��ua�[k��\��j�n��«8 }J?�nh�eW	�wL[4��ܭzl4l6�75?�vh0�;�@]���+�Y�u��yVݣ���5BL���1Ng���������8�¹�D'�]���Bhsv� _�=����q�a���\�^�+m��o&��`8��j@�Й�v�׮���gs.�ػ���:����D�;ĿP�v�ߊ[7߈�=���ˉ��a�q�����H�1�6� �^)��t{���F��_���\d{bW�����*����_��bV�ko~��n�{ww;=��|�*E�#�튌<�����ۄB*���zw`�|r!R�v\=aQ�X&܀���)55�6��^^�x��?w;�Qx!񖅭#����~�/+��,6|��)ó�S������8�Ӣٲ�+'����}a]q<���DF=��8�a�]����pl)�$b�0�|s%l"�g�ʐ� �;��&p<�<��`�_��@�s�U��p�jC��0��#O���I:��1�p�삹v��z0���X1�yK~�s]] gFDR!���S��d��wYËӮ�
�] �G9��1F��+ԯ0X��wƻ��Z�A�ޓ����W<��y�����m/tڮ�V1������u2�����c�����2�m���2;�?���>G�/R�Y����D�_.7]VCʫ}��Tn�nucVG�=NLO�TW��M�!D��+�T ��-y-�HŢ��Bq��oXop!sѩf�\��.rG�g�pR6�r���"T�d���R����~h�&�K��فi��M��xفմ.�2b�Y-Rnu��^����b�q�Cv:�W饚Uq[�d�_����u�0h��b����v�,t���5E����W��lb����@~+P���+J�N��W�aaR �N�0�-�$�+��wpBΉ��άW�[�s,�S�0c
md9k�I��d�N(`��G��^po)@��c[�}��{,���t``;=��}~�D8p}Vl�.��]�ac���
�m�F�2=5 ��cf<�$���Z�����9P//�O�p{�$}ēE��H�l��iK.U��p�.v`��w$�-���JT�Σ��e�~FK�����-��6���1N�B����)y�o��~�-�c�:��ݻ����気y�*��L��P�^o��ܸ�Y�@h��x����z��j6AJ�i<2����H����`j�=sw��vX�:��m զ(2��h�Wg�D�xS��a8���� u{O��B�����/��YL������yf1��-�<������ѣ{G�z�Y3P3����+1N����3�&�4U���n˵���'���d@����x�3��øw�9��r3D�����Ni%@���e7�=���1����!;2{7��@���D���:����I*�ӯIh3���d���X9�K�*K'��K�M��
�hُ�c�9��x�/���K'��#��i�_�����e�YN͉`�Y z�����T���\��v��,�N٭W3�E`(���&Ш% �I���03 v���r����ou*�8�[9`��ے�c��:9���Ƥn�c�W;NumA:(]GbR�FsHOu�,���U�g�E�a+$��k\[�}�WMO��#T?��������2:)׬VꞤ4\���D����̓�@�8�+2��)�>�nVm��>[z��8�e+�|��,�ۛ�,E����?D�G��q���g����U��bN��@|���h�5 ٴ�b�Oj�	"K�k�
��ix���4���?��8@��j`�=�p��|����ڝQ������o�eJf	y��H A#�D�aR�̚���i��V�L5��X~Cz�����Z�X��c�n��!	k��l�7h��~�03��O���x$����kr0c���|:�|z^�ETz��1�x�ڞ��r
���i�JSҋ͒����Eл
$0.[���{�à��@����7Y����y��S,���M��U��$�+q��Q��� �!{��C<�,�;��\�R�ɝ$t�_���2������>˄EˎD�JΪ���*��Ⳇ#�[k�\ǘ�y�Y��˗�*�ӓ*�X��%�B��j������@�Iҷ�x�r����+:�NrY}ĭ��rN�kx��~��%��F��E:�[!��1ELA����*Y�)�T�>m�.�k�o�ٯuI �ao(�Y"�'�d�QPf!���'Q����S��T�nW��p�W�^r7h�3`���{�Sn��_�ϥ�_�d�*�-Y��na��`�Z����ʘQ��'�-���Ǆ>-Ԕ:�\���V>����x�L�[���������k_.�� (5m�4-��ѕ$YNv}���ʺ�L}��׹?�æ�(�M�n9��Ic��C�&<��¡2�O�zC!��Rne}�S���<�^�2l���Jiݍ����r@2�B�����X�^<N�%ȧ>�p�Z}�b���-"���X���Z���g>?xfq��oُ����"A\�hA�4Ք���I|W�?�)�<ov
tG�;���x 0,Ik�>
�B"|��!�P�&'�Ӂ�do�7��IBL+��1��������#�p�$�߿�xV绖������mIv0I��Q��#��1�LvZu=fo4R���r�>6*�0�U H�fnt!�x��*Pk��]�ND�o�ϕuZε�ת��X�Kt�@)I��C;Ԑ,�єVa7�/O�-�')E��hP�2���br�/��ؘ؉��veV,Uz�,> ���	�W���P樃�֋��|�?㌱S>���#���P�@(o.��@B96\��Zd���ݨ]��*��e��ȦȘ����2 *���+������Ӹ�Pe�p�*|�7]�:6j� ?����V���G1/WI��Ɗ�6uYLFB^m��.?Y]7D�e�h<N����6�����Lp�u�W��5v����чY�6V��J2�'�~�\��k�!(U��R��㗥�n�[�B�*�b(�0q��2�b����Ivt�6�)Rh1����_Hv�qm�<���CQ+��iIK�LL_���a��㤷����/��&X�u��3�sK�`�X����4\�G%O�f=X�	}�[%�5�IY.벽'�Vt%Bv�ꉛT�"3���k��!�DPز���*��奋c7v�=-0T��NQ2�;Q�}��r���ךiw�����z�-�,ũ}&?Xf1J6�@��r1��J�Pp*��賌�ݴ%�f�<uK�4x�끗?15�m�a��-�N8�$*�����t�$"�Θ�O�˭s�F��Rs�Ϸd���5��L�R�I�_ڮ�^�^DgSV��}y��?)b,�wm�V=�tk���8�gh�,lx���fF�~�A�-��=�t=i��h.�L�T�\�,��/���A�����%�ʨ�(�7v��θ薳�\l����I��(ž��L�C�����m�T	,	ȩ�i�6�9�(��Ms�&�8���0ɂ�m�c'�{�,����@Ơ;���sPq
������G#5����3��zd]��P��އ�.|!e��`o'쩖;GjN7�4�C��Ϲn��M��m6����-��T|�K�{����
�Ϗ����62����H�	�g����ө1��@Y�T�/�0�񔱉�]樞�ΐ�[��0�"bX��9K�׀�˷��]ʆ�"�T/���.%.y7u��� ��^O��3�%�p�K�D�ߑe%<�7�7�<U��X���BW��h��D���'�
ր�/����sk(��6>#�0V��9���8b1���>�no�ϸ���/���NdϮd��]��%s��Np2�
=��!�ɦ��D���˾�ٺ�s3���g��p�Rk�a3�;���)ӊ��0��"�Ki���h ^R;�/���d���\b�� ����TrO��6�}�0�	%y�c�:�<1�sR�Q��>�����&sg�[�y�B����K�½����SҮ?T��=&�f����7	�`k���Sv@؀�G��k dR��-���n(`i�ą��P�C4Q	x2�n�W�(�S-U����͉����}6y�͈|-��&T�6^̀�k ��I�*5N�..9�PWY����p�.�I�����u� �����n[dnz��Ϫ;��(?&݈���s2��b�{�����n���Sw02��e>���ȂRui��'��nS@?���γ�Js����ִ���h�3�3�Z~ʍ���"��0	�V�B�VZ��"g��8fR�o���
x."��(��]?4V=�ӂ��|s<�
3�oweth����� �I�qL
X�|rp!�9jŘw�̅�֥e�7Cw�I��v�/J}�Q����#�S�$#�ֹ�J����Jw�5�0
���2�4#����mJ�u~�"4�b��T��>�&70�xGU��.�g3�!�t���3tkY	����¢|}�V7�Ζ��׫�X	BK�M��������P;u���W�/7�0�0�q�NM�)�Oh�����r2_�䙼�٬�vfn�U�F>A)ޟK�����L��&ヌ+�qI��M��(>=�#�^PHb�o�c���9��T�4G����-�e:a�i	���������*�#�L���h��semt*_�7iO6Ka�?���w+s�W��~Q�����L[;m��?Z��D�Rk��͛�AW��e��|yaL1 ��]�8�w�٘g�L�0ĀT^^$y
��j���~'����0�>�H������q] i��k|$����x��E�ƍ�s�͏!lL ��%�E풊)\�B/WZ�=;JV�ͪ���D�U��o��(V��Z4�>���lvX�;x�&�U����g�k�U�<��8B�Ձ��fB7�K�8��YR]�F�-�%�����o��q�S���Ƣ�S�!���5�[��\�"��.�� �Db?]� h@=	0B�[J�O��EH�l��p5U�av޴�h���������Y��1�?<��}�5X���aZv��Aw��5�����O��'KO��_�s����5=\L��NN��a@&蠲�b�A?��a�������Ʈ�Wh��)�v����x}��W.�CN�Z��:e��Z.�ĕV vg�6[Y
��{*�W��Ї}�qd���o�H��Z̄vԴ򼝊o1���g�������bm%����*��i�Щ�ugb,��o?Qn��wQݣ�b�'*��O�C@E<o�۞%����Q�HS�wv3|H�ɳ����Q/:������F)��L3��4q���R?�ܲQ��9�[�o#*�5��Ga+�h`,�uު�\�	E����t�8?3R���+=p���Q}��R<Mk0�^F�F8��I]?G�ʆUp)����Y�s{�5V�fsכ�|�m�R��`��6��t3��l���(�C���$�����_��^��1���p�[n���z-��DI��?j~`x]38�F�d�]��t��Ml*�i>
~w�]d=��L�F^bg+*LX˖�w�D|�f��A(C�ޢ��[@���U��mE�x��U������;�^2' �|�z�I���kyKm �2;�?�ï>a
G�|��/rm�A/G_�t%l+��SmUT>�uq[	G�@`L�`��w=أIb!Z��‌�T�����g&�^~�š_���D!�%f�3`��,r��<�����HO����ݓ����h�����~�~0���H�曆����M�F�������%�$=D-�>Ě	:��O�b=j�C���m_R�+����2���ꯥ0>8�b����� t�V�>�S��ݭ�,�����6Y�8F@�"�����Jksz��W�a��wN.4-��/�z�w�/։���΂�[8i�کd{c  �d������(v�G��pU��Rcq���"�t�9�=��l~��p�,���s.a9� ʠ��O==K��`bҝtz,~����}^�h�Y/���܆�@{��$��EZ1���LB��i�֚�t�k�D���Ł$�1
�<�H�1'���~~�).�N���C��6�H��ǇWB&U��) _�E�K~B�c+�ǐ�M����I�| \y����b�%P�l�+��`!�%�#���r�e��jL���?b2tpx�ێ��Εj��Gw�v�2C�� ��}2$�e���D�,X㪘ӌB��v��e_��&ф���vYb.�W�����1A3D�������g��GG�YIpٞw��+����P3�a)4��]��G�9���!f��@d����
�3��ĸM�X�`5D�K�b�N?�@B~�e��Mҕ;�1��E����{�STV<
�$J���T�R\d���h	��O_��E�@�a�gRGu�'2����D]�~����#)��	���s1�y�ʜ#ב�L�2<Y���V`�^<�̮��a�a���dC��q�1y[����S��+�1��7p�*���Az<�~��z��y�~��K]i�;F�ʈ�����I0&����_�=
�e���ܔ(��FT^+��FXAh�w�D �\�A�ȓT?�ꆕ刊��m��_�,c��$���q2��Y���
�?�<�!��mv 2G�?��^>��G:E��eI��7�_:���>ݫ���T�/u'CG/LLbș�˚�Yj!�̓��T����9����r��סc��d�v!�dzf�a���qrS; �����~���w/��p{���t��k�	��W���eǧ�(�M�\���"�@ZQ>��^P-^~T�p���Tnb3C�9����l�aZ����k?¯S�0t�b��ǂx�t7�m�j��I��c�A�����W�@���Q(J��:��:�a^��N���-�K���Nw|\4�$c�θ$P[.��_��c��bdE���p<(��QG��p�c�L@�c�����:���~tl�=6�$~੽p	]��:[b��sao�fʖN�R~*=����V���0�/m����\��^r�/;;���d{��o$	c9E!n2�]x]i�2�*b�������$������U�~������6�~�ý��B��U˟2��{�8~ʀc�h��i������r��y�~c����P����H���<�������˯�h����Kej����u�2j$����X9j�\w��vd�f. ���2�#�cy�D2����&`�8);�,�����Nb�z�M;�}Y��ƻw����1�|�9B���]��]<^G�$.Y�;���+�Lf�ȸ�3�24"X������#�V�]���@Z�Y� �3:�`���i�V�mD��qZjNu�@8+�eC�����1쓡��7�{C���IV�P��������_�h?E-v��24�׸�K3���Ԙ�̻���`씖t9���x�U��e3v� �D�)�k�
�:�/e��NY�ٯe��4V=�y��,ڵ%�����8�Ne�>3�`�,)��Ĩ��-I�e��� ��/�!k�ţ�u�B��g�
�w:��o�4:�ڗ��	a( �c�u�4�:+1JG�|VF�O���v��g�?�����\�	}�2O~��TK�ˡ
� )c\v�EJ\!r�P��͏�����>�l)�3nbZ����z�B�\�B����~Q�Ҳyȁ3v� x�y�ױ}N�M����U]@n L�kT��>y'��5�V���)Pj��'K��"ݖ���uIv�����C/���8L��j��|8�|rn�(��f\�!FV�w�J�q�	�H�����R�5JĈe�i�sAV�65��m�n���P�o��dR�c[�y�-E(k%l���|`O�30��sO�[x���   �  �  �  )  p*  �5  @A  �L  6X  �c  �m  �t  �~  `�  ��  �  P�  ��  զ  N�  ��  '�  |�  ��  1�  x�  ��  �  L�  ��  e�  '�  �   K � (  �( 0 �6 /= pC �D  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr�	p>!��L�>P^�x�#\`yq�~�tD{���O(dG6â�ߘ<����F�N�B6��~�'.>I��]�(��d_�R>`��	&D��3$l��� ��'y��T"`/"�	�|az�H?X̴Y��ǘ^�B| �e �x�@�?	hlHG �*&���ɵ@�<A&��H�'�T)r��u����`��/T�i�'�S�č��F�P�+ 8x20��ĺ�y��Y8#N�P��1�P	�BL��'�)�s�Y�1~"AۇlX<�XAL<��8h�B��.z��s��N�@�}�'fvM$��E�d^� jSG�>l%��ρY7H03�,D�������b�]S�lZ�r�̹�'i��1�	��~=Xc@ѯMb����ėL��Մ��?�Ox��W���`�~�p�B��>eBV��H�Yw�^�]�*�x� �nN}��/!D�����^����b��WL����O�B���J�l�٧�QM�H�R�ϘB)&��$:��«z��u;!L��;-�Eaș!��5z�y���6G!���.Q��G{*��\�Ǭʓ��-W��S�ə�"O^���.ONA+F��6[� j���%|O0`� �B�v�ڍq�ڂ�x��i�ўʧ`.Z��y��V�k����=y����&j$�y���^9la��&^r�8Ql����)�O�yA�B��6-�Kd�+�j���yrj�8tE�Q���T�*�2����y� G�g�j)"q� �O>&ݚg��,�yb�D�#ˌa�E��^02}RgN���'|z#=%?�j�a�/>o��rw���b��}�S� D�DjF��$o�`t
�H��,�n��1�>��p<�R�� ��x�h�&RI�$��`�<)Ǡ]�S���C�g]wh(x�ԟ4*	�)�d�p篆%%Æa��*`��H��Es��:u��n+���ᑧ y���A�^89�`�<�0��%kwL1��9MV���&̟f��CƸǬ5�ȓ��q:��Ϭc����U�� ���԰�&]/+�d<sF��4�.��ȓ׀)��[�A���Ȕ!d�(U���Ҡ؄�P��3�ǶnO�B�I�'F!�6�@��$ZB*�!Q��B��7s���$�p��� !+ց?��B�IWL����C��sT� q� Եa�B�	�23���BK�8Uzuq1�S���C�)� j��Q/�9�1u�M�I��Xq4"O�����	_��K�	��7���"O��L kމ����-u��Z`�'A�p�<iڒA�Z��N@W���H�n�<�`kÌf(����B�"�j`�"��<Q왻Z���z�䛫b(h9`�@�v�<��4W�̅RQiQ2Ć�k��Ui�<yW!R#b�H%B�̟�`�.��M�<!@�s��@�B���$����L�<A�}��D���^F?�5�p�RK�<�3��-6�&�i&+��
��XGjAD�<��F�a�<:�B!|��aE��i�<��c]!ؼ,��&�06�ݱ��i�<10m���(C�I��8�	w/{�<�3n�'�$={a��;�\��3�	B�<a���zsҥ��F]5g��(i���v�<����~9zBd��W�.��!�o�<�擰a���N?W�t�e��f�<!4)��%9g��7iC���W�Z^�<Q7�'+�𛅏�6?:P��V�<Qt�t�T<Jb��Xd,�3"�k�<��a�?pY��Ht
�*T���Kt�Q�<Yv�H6�\xa P**�Hh#�n@T�<1�
ס�ΡS���)
ֆ�I�!�z�<AE���)4�1χ(U���p$_z�<iա@6��$�9V$0�q"�r�<Qt�]%L�4�2RF�]�jq�M�m�<�Se��\gX0���r�T$�6��p�<ɓ蝟Wp��2T�a��F�<ٖgE��(
@\��2G\�<ī�}ߖ�I�E�l�`�[PK�}�<�%��{�\t� ��>D��� w�<�c!H�Kھ|&�Up�!B�q%�C��CWx� �i���-���
�B�Lu�u�4�R�i��#Q.p�zB䉾^5k�)�T�p1�3L��>^B�	�U��a���=n(��3��i&B䉺k�����Īsx`y%o�'x��B䉦*I�ӁRZt��rD�<U5�B�I�Y�ș��#|�(
�� l�hB�	'���+ρ!AVy�N9}rhB�I5���۳Vm*�b�E~�B�I����U'Ѐh�^��-�B��_�Di:rcʸs�6DY�+T�O�C�ɩNQ$|2g��E��P�a�im�B�ɭQq����S�)���sE�9SzB�*�ع#́����;��â�NB�	&��
nLo��LXg�I2^B�	;����#�����e�KO�B�;i����55�R�Sd���xB�I�E+`�A��Z��h�'��C�I�q�Ґ����/~�Da#֬��0�rC�I-�H�(�ѾSJ�ҤJɂ$XrC�I	���w@�4�>0�BL�\�TC�ɚ@�B�� �� 1�I�K�)� B��T�@-�4OW?;7�ơCI�C䉄Bq�Abe"P�'&�	���	=fC�	3/&)9��]� (���Q�G�B�I;p�i�OӤ-�&��c��q�
C�I�4(��];y`�M`�/�8�B�I�o���3 �X�-"��G��C䉷s.`�B�S٦	9TΎ�8\B�Ie�θbu��:P0��'F7u�ZB䉃>Tb�"�ɏ%�P�āc6B�)� |��V'�4�H�P��-]�(U��"O^�3���h2j5�F��o�6hp"OL,�2��9<ct�AބM��A	�"O${)�+3�y��*��U�D8�"OJy���C�H�쨰1�
U��-��'���'�B�'��'���'���'���%u&q+G���'��Y0��'���'oB�'���'c"�'�"�'�z9Yq��*g�Hr�F�A�^�ʕ�'(��'WB�'�B�'h��'�2�'b��yQ�H.&�*`�`�I=�\��'���'!��'���'��'���'�>9Q�� ���g���l���'z��'��'���'���'�B�'t�H�r�P�7 ˔�G�VC
�a�',�'}�'�r�'B�'��'F��s���L
p���M�,\���'/��'�2�'���'��'���'Z��ql
�lr��D�":��I1��'���'-B�'�R�'a��'�b�'���a˖�c��X{����TJ:X���'I��'!��'���'b��'@"�'G�@u���\H93B�p?����'X��'8��'H��'�R�'5R�'V�H5�-r�,�C�$Xd0���'l��'��'x��'D��'RR�'b<$� '�<3�)�� H8mxv�'m��'��'��'���'B��'c���Č��Z�b䡈5'�iCu�'�2�'e"�'�b�'p�hӮ���O�x`E@�a��B@���EЀ��Gy��'w�)�3?�B�i�!�B#�g�̥�T���$����?��<��mA����4�B��m�����?5"���M[�O瓩�jH?�0��[��<`����B�^%�2"/�I̟ �'��>�"6��Q�
%�QI��/�T-Cr�Z<�MC�a̓��O
�6=���#J=Lkܽ@t��=�J|�@��Od�d�Pէ�O�1 w�i{��ܒبg��
`.U�p���[�h������=ͧ�?I��)X%8dyKT �Q�"i�<�-OR�O��m�N� b���W9�A��>e�x���'Q��T}�I�@�I�<��O�9#"�%%�|SG��j��Щ�����	�i�,�C�:�6i�R�Z��(BU�D(����/�l������ry"^� �)��<� ���u�"L�MZd"%ώ�<�S�i�ށ��O��n^�S�;eպ|H�bk��vR`%:� n�����|�ɾ���lm~2=��,�S�U�H9'!��jX�ђ6ƷVjڠk"�'�<TS�' �i>y�ڟ���֟��I�f8l|�Gꐝd���vL�$[|*5�'3�6��U�~���O��$�|����?)�ɐ��h�.)�T�ZG��#��IӟH��x�i>}�	��,��aó$.���4eЁ25�c�P>?4�hoZ^~�`�B�����?�����<�/O\1�R�@�c�  
R�̴yIrd�ҋ�O,�D�Oj�d�O ���<���i������'O���O%�Pȫ������ti��'Zr�|��'���ҟ���џ� ���`P��d�M���g�zF�lZ�<���_�p:`?��'����w�����E
&O�-�bM�:7����'\�'�b�'�2�'g�>���%Ƒ&��|*U�ߦ}k`�B�e�Ol�D�O~ow���͟��ܴ��)�$����d��Yk�f��f}+I>i���?�'{(�1�޴����2$Y�Fß7���h�2Tk�Sq���-o:����䓯���Oh���O���A�r�>�Y�S2� ���ӄr��9� ��"A\�mK�f%�3g���'���O:���c�t�eӎG�|��%���yB�'�:��?��O{���,Z�N�!�F��^����-e<H���ýjw���I�?�� �':(�I�[Ij扂�<�Y�K��7�&�[B&7W� t��͟�����d�i>u�I꟤�'O�6-����yHcG�^� ���}�(}*RI�<���?�,Ot��<��.:aK�l�>}kҠ{1��:�����?Y��#�M��'hNY}�Ԩ���Մ
5k�*�N��"�M	c���<Y���?���?���?�*��HRwm̆B�� [��Ú@��U��򦭉b�ڟp�I�%?�	�M�;:0��KNn�� ���	�4]#��?�I>�|r���MC�'<*���e.�(0��;AQ9�'\6 ��������|�Y��ȟ�YV�PT���IF���D}�U��؟���ߟx�	Cy�~Ӽez�M�O��O� b���C�i0Lu 9h�(�I���OZ����Gy��m�E�T*�FL"��&?ѰK�)Y7�AD�׊��\5���
�?�@��W��d�S"�$2μ�1�$���?���?���?!����O�]���Αf;�\�q��6)���r��Ov|lڭJU1��ԟ���4���y׉¡ ��"C�_�;���Q��_��y�'d��'׼i��i�iݱP���?5Z��o���À�0Il�������'M�I�(�	ӟ���ӟ��ɷ`<0�kZ�HK���%�wJ`�'�7� �8H����O���t�	�O:��>	8��0D�B4[ΚDZ�陸m�<��'���4���$�OR@��B�nl�A��hH)"�XP�h����6��<iA� )�����?�eW�<�*O�ۗ,��e9�i�EMZ4y@w��O4�D�O>�D�O�x `#�<�V�i(�28�>�Z�V�(����UFUh�U��'�d7�1�d�Ob��'���'2 ���z���@a,V!�U�-/.��i���O�5Т����s������ 5��;B@�8�㤍�o�,�'5O.��O���OV�$�O��?yS�'���&"��F�*�t)
t��������\h�4iÊ��'�?9��i�'��]c1iL4���[4�S�M>j��3�|2�'��O:J!s¼i��i�5b��
 	�P��^'?� ��k��0:����d�'8�Iٟt�IꟌ�Ɂ}:0ٹ&�Αo��h�2"O--F�D�I۟\�'�6-�6����O,��|z��}�Bh���k�kCM�z~b)�>i���?�O>�O
.|W��?�@nFe&� ���#qQ�MrĲ��4��X���`��O�A�1���Lc���$m�x�i���O8���O
���O1�:�EH�fLӸ�b,���6�j!zv!R���'M�`w�D� ��O��$׆l4�؞�|��U	�UYr�d�O�����c��Ӻ�6Z��U	�<� o�r�a1�d�)+�
	R��</O����O���O���O~˧b44IWc�G���u��'m�b��iq��h��'�2�'(��mz�a{ �K$9,�K儇K��8�m֟��I|�)擊�6]l�<� .J~?"a�i+�^D����<���&���D4����4��&�%���S3��a!��Nv�D�O���O|˓G����J9~��'7��.wTH��`�z`�
���O2Y�'���'r�'-��Z��@:7�8y@���Y"���O�9��Z:?�pD�%�:�?�%��OM��Er
�)��?~mB�OF�d�O�d�OJ�}z�ZG���S����(�&�y���=�6�޵>���'u�6-'�iށ����>"�xb�I�k�2�B��{�P��ߟ��I�c�LnZ|~B��L�R|��w���%�3�T`Q��688y��|�^�����p�	��	��\{OJ�18������Z��-��xy��t������O��D�Oj�?��KEk�,A� �V��
���%ȟ���OJ������	/HcJ`���R̔���ȟ�3�ԲףG�����'7Έs��Ο�Ӗ�|�[�l�h���`�<��e�ҟx�����	$���By�d��ԣ���O����o�<Yy�����ۘ@y��Od��O���|�)O����O���1u�:lJ�k��1Ϥ���#��@��kr�@�	ǟ, ���c�TU�4��Vy��Or��?�la�P+��[ڬ9U%Ǵ�y��'�r�'i��'����ǚz����b��tÌ\1u���P�p��?�i!<):�OO"|��OR��*�gx<(@+�L>)���$�O��+�x��ش��8T�|���P�y�Zˀd/�%CG�@��?1��(�Ġ<1��ɮ;3����K�Ha�5�ML+�O(�lZ8������	v�D�U)D�p�1]2<�Cċ���EB}B�'�b�|ʟ葑��:����W#�Ce>H��TzHP2E遯y*���|�a)�O�I>��i�`q�\+Q�P�k��I�`/���?���?���?�|j,O�oڂ$�9Ŏ�E,���cX��8dޟ�����M#�rd�>Y��M��3ꖙ�\lI򄅐L1ֈ���?q���M��O �:g悯�2I?I��Eށu��Bh?KH��#�k��'���'�2�'O��'�哢O�a�œ�]Yz��O�<��4m��)O �$��8F�O��d��]	
�lM�5�Қk����VNR}����쟤%��S��L�	��~�lZ�<����7s/�z�dH�C�*����<9�A |I���z��~y��'��"v|Xe�j��~����kN)k8r�'��'���M�q�?�?a���?�v�H
}ˎ�Іm��z	�ѣQoU���'����?�����z#$,XU�E��bx���4[�'�}���@�t�����~B�'�00�� �z�,FE�m�e Z�<���R:|! =��R(�< Cp�A�?���i���U�'
��n�z��]�D�f,��+H�62��UMב3�\����Iݟ���d�ɦ��'t~U�5��a��lݎJIjl��∞%��T�	�?QcK�<)O��������O����O��!`��9���G@�,�&pHv�<��i��՘�S���u���'�R�B�Hxt�U�_}�(���0y�I����P�i>��	 �Gh�7}��l*PA�+n��(@Т�U���o�[~� ��"iV���䓶�d$4����ʂ8d�*q��C�Ah$���O���O��4�,˓@����4���¨��ـ�@F�HoR�1r�xӞ⟘B�O��$�<��H�R�V IEG������V�3B�	Qܴ���[	P:�8:�'@���n�+��̲�L^�HN�I����2���+�OX�	���,I�2)�FȾ�(`(�Oz�D�O�Imڿ +�+\�Ɯ|"��.)p�I�A�U8����(J�'X����� }c�V��L��O�=oR�<���;9d��YPz�G�oV��4�D�<1��?����?9�-	��4!��_�>5����?�����D^֦A��Lğh��ğ��O���QA
�4�ҁ�ӌP�C��U��O���'���'�ɧ�I �%�R=c����0j����=D� ��-�7Wv8[S���ӹo��|�	�P��x7N��G�9��'սC�^��Iϟ�������)�FyR/m�������p��L���ِ|�0
��Q޼�$�O4mZ�aC�Iݟ ���Y�d��A3��֎#�;�ȟ��I�I��)lZZ~�#�#w��=�SJ�� <�*�+T;0���ZR4M�%��7O@˓�?���?i���?����)�)����f_0fn{6d7ElH@lZ#���I͟X��Z�͟h�������5?���:3-
TNd�SĎ�?�����Ş&�}�ش�yR#L	e�Ό(G�\�]��A0�Y��y�L�r��)��Z�'���֟���b�&HQ�/\v�J`8��;L���П���?�@D�'�6M/U$���O��䍤G�FqZ�OV`�����i���D�<���(����H�?q��Ҥnk���I)�}Q"! �<���HшѩF�<|3.O<���'�?	���O����|NT�ǯ�S�"�Ba�៼������	��G�t�'��`D��1O��}QE��V�ѹ�'�(7�"�n����4���ɝ�w���S��3C��(�?O\���O���;N��7M0?i�LV((��)C'�y��7RVJUrF�H$<$LT�H>i.O�)�Ov���O��$�O� ����
?�USɋ�uZ~�2a�<!ּi~���'Zr�'��O[�N͡I�F���iY�I�"��c��/)*���?���ŞM�zJ�}��ՙ��P�T�w^�M[�OB	"T ���~��|R_��Q$M*;�0Q5�@�~;0e�t�����I՟��ҟ�dyr�t��c�!�O*kP/�S!�t����R�@���O�$mZY�QG��ݟ$�'��-�j �C���`懀��`P$�+Ư��������}N��Px���eာ>� � �G�CB�2�`����ǟ��Ißd�	���2�f�9oI�`jD�g��;�Α����O}m�,�����0Qܴ��`�Ũ��-;d���f#�|�t1JN>����?�'#.i�4���3P1̈�EH	[\���ٺ)W�kU��(�~�|�V�����,��ПH*a����l	���@�Լb���d��Zy��n�6@Ԉ�<1����ɑ>��)HV����AwE
,/��I���D�O��<��?Ś�JĘZg�͓����r�����i�D���w��%ʥ<ͧC>��Y�?˘A��E�9b(Y�f��%��D�	����I˟��i>A�Iןh�'L6�"\m�pK2/��v���S"�wC0�����O`��Ȧ�$�������O�5�s���F<��@�]���Ps��O���@4/�07u� �Ie�x$9�ܟtʓ7����Ď�5I-N[F��(0#��Γ��D�Od���O��$�O0�d�|�g�H�D�T)YW�+�t�rV��;_���%�B�'���d�'�7=��� H��m�@"�	�K&���Od�D$��	��nR7�e��!èΥ8�<�᠏"""d*�g�T�s�	�!t��Ey�'M�� 7M�
w#`�K�!$Q��'���'{剏�MC2Ȃ��?���?����o"(�Q��`m<E������'U���?������̙�$��hoM�RV��'<@��D����Ȅ�~��'�5��Y$e|�1jҨ|�L���'�6�z�cC�
>��œrN�!�b�'q�6Mv�j���O�TlZ_�Ӽ��È�L�Z�ɂ*F?:A���	�<Q���?q�6��Xܴ���яn�uQ�O_�hŋ�4C̊�Yo�x� ��E�cyr��(P�X�Ba"���S�
��jy����,	������	_�'6-�w�	� tJHؤ�����	9�S���Ɵd$�b>u�ėNK��g(�5�e��n�b�lZ���S�WCa0�' �'��IupR��֜~��� �^���I�x��̟"eߦ
��L�'w�6�@;C�����3Yؔ�B��@{�:���-A��DZ����Icy��'g�듖?1*OP�iۣV�h�Z��(��ғM�`��7|���ɝPL�9���O���'v��wz|�x�f���4�L�e���6Dz���I��(��埤��П��:t�N j�91D�ǘ�(����?��?q#�i����ȟ��o�X�	�@�8��¹(w�H�e�Q3T�'����ş�S�J`oZQ~/Гl6�mZD)�-R<\
��(���"�g?�J>)O����O����O~�#��� Ls�ib�B�(��)e�O��d�<���'Uf`���?������xdTp�Hʀ�8P�Y�<i�ɤ����O���&��?���f�`)SC� |*��f��X8X!���2?���|�M�Oj���n/R�Γ]@�Ȑ,�HW|(C��_�o|��@��?��?��S�$U���?�M�G���(=��QҪ1�f�@���Q���*O>�$ �d�Orʓ�?y�-��X�P�ߡR��#�a��?���%Dm#�4�y��'S	����9O�Z�N�{f�!��fM S�$�v>O�d�O����Ob���OV���O@ʧ
ծT�f|6Be�� E�-�M�Ҹi�HJ�!�3�b�'���O�'J�wb0���P�\��s&��2,���'X���i>M�	��%���� W\U{���5R�)���B�̓f�8���O�@`N>�+O���O��+@	
.(����a \�T����`�O0���OP�$�<��i��X8�Z����1%ؘ�9��=z��]���J.<�?Q�Y�h���T&�sDQlW�x�d`+uh>,��!?���ȲlD�8@ڴ��OȊP���?!Ъ��Z!�4�ϪsK�l�%�=�?���?����?���I�O��r���GNU�� r^�HWM�ON�nڵ\�I�| ݴ���yG���H��	�м�!^2�y��'�"�'�vIPE�i*��4/G���ܟ� 2eab�D�:`�* _�`Uj�:�$�<����?	��?!��?!"��7/[ }���X�KyJ��i�0��D��M�q�F��P��ԟ�'?U�IB�R�q�*�7kHQ8f2�!R�O|���O��O1�bt1���W�(�&�ϗg�qP�K� Ak.� �!�<�J�J
�ĕ�����19 aJ`GX	,\^U���N�h��?Y���?ͧ���Yæ=A����p��K�h�p����0r�����+Y���޴��'v���?����?��n��xݞ͋�T� o�Ueh �r�L��4��D��\4�������P�s�痎Y�bD\�.]�髒7O|���O����O�$�O.�?1)��\Q�5AU��l��i����ӟ���џ��4�@yͧ�?ad�iv�'k�ઁ�QB%T��$+H6f��i:2�|"�'��O���$�i���+�j�A��U\r��(S5c�%J��$���6���<�'�?���?�����	>�$J�-G�2IZ$�[ �?����ę�əńןD��˟8�OA �@i_�v�ToZC(��y�O���'H�'�ɧ��@�C 4A�LY7bu TH4��~���&�N�x�us�����*�BLM@�h��h�'�*���Q���=�� ��͟��	��0�)�wy�%q��5� "d��]��$����IĘ��z�*؛���u}b�'6�PI�#bNT�r�(Y%Z����b�'=�.�������������<��e�� m��(A�z����i��<�(O����O��d�O����OH�'�2]�!u<!3 Ϡ5��
��'��dA��?Y��䧁?1���yǕ�v�x��@�6-��"��z���'ɧ�OV�y���i��F�vF2�I^�E���Z���X��t�̟xqB�|b^���؟hS���8-���a�GQ_Z;'D���	۟��JcyRO`�x�!�C���Ofayd�1Ht��aD�r�"��O
˓�?�+O����O��O�uA�LA��<SA��z���2O��$�1(zP$W:2$˓�Ba��O|���9�XĨ�G!�n<���ι6��dP��?���?����h���_�U@<@���d��=qbm t�������
S��d�I��M+��w������R�Dl�xQ�x$�s�'	��'C�=˛v���ݮl ��SLRQ�B�]�Xz PJ	�>�蒕|BZ�`�I��<�I��|�Ip�"�9k�(� �-�5x���sy��i� ayR/�O����O�����dV`���"]�H鰁��
m��\�'i��'Vɧ�O�b<�g�6��ġErR�iH�L��C�J��c]�@�$�64�Bf�g�wyN�xà=B@.��e`����EY7h��'�b�'�O��� �M{�n^��?	�L�_�N����81�7N��?�c�i�Od��'�r�'����$��} ���yC��z��0ۈ�(�i��ɦ#�l|�tٟ�����"��M�TW�9���ω�|�D�O���O��d�O��d3���[��Jtj݉(��i��@ϸ|�8��I៰�ɕ�M��*_�|2�s_���|"+[er����S�dQ���@!��'�V�؉�A�æ��'��=P6��:V�T��FD�Vy���K	;����	�Q�'���şl���x�ə����2�K;|%��#,Դ�����'� 6mCw���O����|�,حm�� u�2�	��ZI~R&�>���?�N>�O�@x�d��}�@����+�.���
O<�|���G��i>����'�&�x�Ŧ�.@^��$���G�B�S`�Пp�I؟@���b>ݕ'�7�M\�PA�p��`z������M}!�F��O���V��9�?��_���	�=�p�y�'=��� /�!l�����؟T��		ئ9�uw"<���/�syb�A;u�Ii����2�L��l���y_�x�����	�������O���+<���'Y"M�<LP�KjӚ5ӑ��O���O������Ħ�ݏE�:�rdȲ+b�av	F(��	�$'�b>e��Ǐ��y�:Ī��`کE�R ��J݄qߜ�Γ!
&��䫥��&�|�'���':a�%WY� ��D�_~� �`��'B�'=b^�H	�4\S�Q���?�Rf��@*��Tc�J�m޻��b���>����?YM>�f
��F&赛��"�
�Qp�e~��?�(�ّ� �E��O�,��A��I�	�N�`�q���!�$m����'l�]��ɟ���0�	E�Ӷ4��П �����H7�`��Hl�%N��J�4PV�Xp��?���?	-O�9�����@	���Y��Ԭb��jW4O��d�O��$E4�6�b�p��O��R��}2���3@��r
��"�Q�� :�$�<���?����?Y���?i����(�L�b���.��"�!���$�1�E"؟$�	ן�$?!��F��r@�=|�)�Qo�d�T��Oh�D�O��O1�qq1���wҩR��a��hiW�˪��	�&�<9��V�$�L�d�����S9_�,���)U��LM�4"�#pTv�D�O`�d�O��4�d�c˛Fd�*�h�T�D�S̷3����W���y��h�㟤[�O|���O���H
NT(f��4Iv@�)ʂ>EΑئ�iӲ�(�	 b2ʧ��;&K�'.�t��Cō1��K����<����?)��?	��?!�����X���?���K�%ſBEb�'�Os�
(�F8�$��ަ�'���K�d���c�	J�^`Vy���@�I����i>5��A��=�'�D�
� ~�($j
�k���RK,V�e�aՋ�~�|�Z�D��۟X�	�ɷAk�N��b�8REZE�T֟���LyB�|��u���<A�����yR���O�Tr� ��8t�I���O|�$,��?Y�W�c�����9*�ʬKȥ~�H�q��������t��o?1O>��h�bB�AaTAT*z��$1Ш��?)���?���?�|�.On@oڿ*�L��������l�;
J��!�Dܟ�	(�Mc���>�OF}Y�����p'�"Ob�����?!�́��M��ODe�J��O{�q��g��n�f�J��c#.�x�'R�'��5H6��'���'��O���7L�e>jֈL�Z����N`�V��l�O�D�OT�'�?Y���?ͻ9	,�+�̺ p��r�..6��<����?IJ>ͧ�?i��9ɐ���4�y2N�0�;���+w"���ɖ�y"��C�ȴ�����4����A ,;acɏ���c&�ۍ[����O���O��5���C�Xu��'�b���̩�aM�S4p����¦U�O�h�'I��'6�'32�҄��v�`Px�.3e����O^���fޜW��7-�^�S89��D�O♚���)LR����dR�i�^]T�I�����OB���Ox��?��b��<��%|�(�"�n�|d��Y	s�i�I;�MV)���d����'���i�55�Kw��ɰ�If6�)��|�����4�	�	lEn��<y�>��+6a�Rp��CO9o��,��%WO`L37oJ�����4�
�D�O����OV�d�
x�^� ��c�H�x$m��[�˓\��#�i �������mH�h�t���p��oW�?�������	}�)擷MO�����W�8]*�ݽRv�S���b��{�r욷��O�YM>�/OH��sD�/מ�
�MM�R�z�)�O ��On�D�O�)�<�S�iJ��'����{�<� C�R  ך!T�'��6�3������O.���O�� �f�x
�KEN2��H׳x`��ݴ���"�M�qџ�����nC�更�TJ�.9i�5�� ���d�O�id��O�$�O���O1�(H�jS�E���*m��T���O4��O�o�6.p�����X�	`�?dL�˵��(��Ȓu�N�{��H$���	Пd�	�W�h�lZ�<�����Jjܼ;8���#��/vF�!a�K�a���������9OۢQ���E&�h^8����MsE���?����?)�b���̄ |�,�U���7�`(枟\[�OB�$�OH�O�ӧ0P`"��2��m�ȏv	nyZ �;\P�n���4�����'�'DLɓ�n�b��kp'HA����'��'r���O)�I �M��X�2��tp�O�D��@A�^(9�����?᧴i/�Oz�'��I�9��y�T	V�5��(ʿF���'$��A�i�I&i޴
֟��9��`�ELJ%w�F=���	΢a��M�kЌ�g�פk��� !���< Z�NO/c������ҁ�QO '5��q�s D���,�dP�,�O�`-��!ǀV�rGÌ
������3��@D���ܢ=ظp�f�R�����Ak��b��]:C�cr�)��Χ�H�W�٨)��Y��U�����i�!}-�D���14"�1a�ău=�q�$�D �������`�8a
Qu���š��%r-���Íi���&�.O�4�΄3�tt �&��sZ�)	C߄/��5o�ß�������S���<�ӌ�'(5p�K
���4Bڑ֛�Vc��|2U>�?qR�^6xܶ��!�I9Y#pH�S̈T��'=2�'{6,X&�>�)O��d��XCMT%�*�x"l���Za91�1�Ɂ	{t%����ϟ��I5Q*�$I��Z��x 0�D28q �h�4�?��.
k��Ly��'�ɧ5(�5^ �Հa�.&��b�ʞ���ď)x��O����OR�d�<�"� ���Ԓ6�3]
�q��W *5��Zv]���'���|��'�"`˛+��$��Z/�dͳ���Z�2)�y�'�b�'��I�U7h�ИO
V���!��hi�y��J�8�4$��4����O��Of���O��$���ز*�)�h�A�=ʠ�)�Ⱦ>���?)���Ą:�̌�O��*�#0.��v��Z�+S*X�]��7��O(�Oh���Ot�3EI1�I�	�DL����-3$�c��6V�6M�O��D�<qG�:!��͟`���?��ˊ	S򢌪��(Gex�j%D�3�ē�?q�X ��x�����d�������[�8%R��G��	�M�)O�B��N����I̟�I�?��Ok�s�����׻v��vL4V�v�'|�o
�B�|b��[�9��ȋ���<#V��e웶�ċy5D7m�O��D�O���_h}R\�ٗ.�m4�H����'?�ER^hX�4j䤨�2���OFm��Jw�4P#�����5�E��-��ǟ ��_����O6ʓ�?1�'�xҗ�Y��rebG8i��8X�}R���'�2�'�I�n���Je���t�\)$0L=�6-�O<)9�n�B}�S�|�	P�i��{r��\��%@��N �>��U8�䓫?����?�-O�a�Ε.PX�L:���̩�D��y����'!����%��������s�]��12C,� X��E�3�H�:ł,$���	����Icy���7#-���>���;ƢY:In8���i��6��<y��䓖?q��:d�'G��ʥ�k�j�@4�ڰr��٘�O����O���<���l���̟���Ϡg����&�L�f �� ȗ�M���䓿?��M[���{
�  �{%��=d|��LB!���i���'��	�{Y��L|r���1#��11͖,Q%��@e��'���'R��'���yZw\^%�A��� ���U�[Cђ`*�4��d��nZ���i�Ov�)�a~��҇_Z|����QT�y�I���M�(O����OR�%>�%?7-�	�bTʁ,��J9 �#�=w�6� J��7M�O
�d�O��)r�i>�h�B� |!<���Ŷ4�@X�Q�-�M��?�����S��'��_�O��ˀ�B�&���$MV�7-�O��d�OF J��q�i>��Io?)�$� +
�T��,��G��u+������\�I-������Ia?��hՇ-\�{�č��@Q�ɂƦ���5:*���'4���'�>��U��j5J��"���$"�$�5b�1OP�$�<i��P*6�Z��V$8�j$�M�Z�@DϏ)���Ot�$9��Ο �7�p���`�Ud�H$��1p��o�1��c���I}y2�'4��՟2�&dٵK?�d��&B�$6F��վi�R�'P�O�$�<)"�Lަ��Gb7휘q� <Snm��<���O�ʓ�?��l�����Ox�ڐ��G��D�cW
p�V�kۦ��?����䈵�'��tq��55���P�^,+���4�?1���DEsj5%>]���?ט�U��]�c�O�j�T��0!Jf(O�˓�?�����<��>8��χ�\�f�q�<Ǆ4�'?���(�B�'�2�'��X���4?�NY��V]w��BdF�8_�6��O�˓L�:ExJ|�^uV�1д���đ�@�4k��ƌڢ��'�'4�d\��:V��tM ,26���L�,�;�]�\kFN:�S�'�?^0
��%O*d��,��mږK�>�nϟ��I֟,��,߽���|R���?��#
�I���3�"I��P�.�P����'s2Y�0ʯ��ʧ�?��'T��5��Wk��X��Z�h~�� �4�?�������A�����|����5k5j�H0��a���'��:f�=?A��?�����D�'QQ�ڄE5S?p��@��\�R8��a�	���j�IryZw��� ��ה%�ͳ�"�JdI�4�?�+O����O���<����X*�ə ~Q�QbZx��x�"DPi�������ןL�'�[>��I�(���c��ޔ�@�7#������O����O��?QWKV��i���Rt�C*aD���Uo�T���w�L� ��IyB����Q�Nဉܽi�� 	#-Ʉ��8n�����	QyB�ؤAO��'�?A���5dC�c�&tI���:n�xr��<I��	�t��ӟ��f
l�,'�D��
�rw$k�X��'�+�<�mnyb<Y�6�Of��O��)�P}Zw��f�ԋ'��uzu"�&I��4�?q��Z���ϓ��ϸO����7'ӂ-HiEa�{�R�[۴��`R��iZB�'���OR����đ?P�]�4���Ղ���!�r�m��*�I�Ж'�� �Dص?����Řd�4��G�ӪR��l�ݟ8��ƟxGi����ĸ<����~"`ұ7�lx�B*I|��c�̓��M3�����سt��?E�I�`��h��1��B�K
r��1h���o���X��BI��d�<����D�Ok�C�Ә|��Ժ7�1��+O"O �I�6$(�I��|�	ȟ��	ܟЗ'�4�rf�� a�t#sE���0$F&��gNN듯��O���?9��?�pC�e�����|dhQᛀL�͓���O��D�Oh�r\��S0����ڂ2,!��4
t��r�i\�	ȟ�']R�'!Ҫ�0�y�%(	A�u�3iX�(%<��n�-s�7m�OT���O��D�<����f���ޟ�7��}ͦ|	g�OD�t!� !�Mk���$�O*���O�X����sӤu����\)X�Mǂ|]�\ˤ�iLB�'��	���믟���O������%^�T�85�jJ0�X���Y}��'R��'�l,�'�U����0(8��ň.�:tq ��5�֩nZeyB�p�7��O:���O����u}Zw�X���'<}�!1��:\$|��۴�?��)%Q�}�s��}Jq"�%[�D�uKƞ:d"'+¦A�v���M����?A��R\�t�'q,��� �X8"b��d&���Et��0��2ON���<I��T�'>�%3���^�Hࢋ?5��Hq@dӞ���O^�dʋ1���'^�̟|��,m˄iP�3�TY��N�2 "Xl�cyr�'D��yʟ��D�O��ж�H<arm�I���CYl�LlZɟ̨!���$�<������Ok�/;i��q���[�@Tk��ɧ~����{y��'��'��5���^^u ��P�d��<1�	�Jvvu�'��Iʟ��'�2�'(�[�@4P|��`�o��I�
�dr:���'	�I���Iş �'@<�A��s>=�`,38��S�+'�HdR�sӜ��?!/O��$�OJ���2��Y4m�Y��*L/(�tͺ�A-@\Jn�`��㟴�	Iy�^�MR`�'�?����m��ĸt�vD#�bK�9Ϟ�mZ�Ԕ'Z��'�rJH��y�U>7������EY`g��[r�;i]���'O\�,��%�8��)�O��d�6ԪC,�H���Dh�f��i�� �P}��'Rb�'s2qٝ'��s����;�=@�"�#oo����a�J�2�l`y2�����6��O��O&�I�S}Zw�X����Hn��Pd�5w^�޴�?��0�����?/Oz�>� ��D��
� |�0�S�T�u b�izpR�}�@�$�O��D�����'���.:�(�!�ˆ0�VA��͞^��(b޴*b�͓�?�+O�?���ü�6�Z�kБ��W3}��H�ݴ�?����?i0+5��Imy��'y����/����Ӝ<��,S�"6z��f�'�"�'�*����	�O�d�O��� �]�vab�c�&G ݈y��k�馽�I�^���O���?�.O����N�Z�� #lDt8�LK$U?���RW�
��c����՟�������ky�.B��Y�<=*�(��f�`qp�>)O���<���?1��'�N��$�̛`O��`΋93&��Z�K�<.O���O�d�<1��ܩ1����
Â`�Q)�|r08`�@G Z���Q�d��Oy��'?��'�$�'�}�aNQ>P����W`�O���SQ�s�����OX���O��.�<�k�[?��I9E��z%aC4o�,���-q)9��4�?.Oj���O��$�R��$�|n�����xg�*~�FГ�EܷYnD7��O��d�<�������l���?=㳈U�*�ԑG"�
<Q��L	����O����Ov��A8O���<1�O}�̉�(�:"x`)p��3$�]k�4��$35�m���������S ����X!֌�!??pt{Q��g�:�ط�i���'b��'�r\���}B�ؗv�Rt@En�#�0�qA�ަia*�:�M���?�����Q�,�'����S�4��H��˯^�|� -x���
W4O����<�����'Z:M�g�,	5 ΤZ�r��'I��'�#��'v<�����O��	��yqG�[M#$�V�L]@6��O��$�O�p	�:O��ݟ���ٟ|�W%ʛ=ň���az-J2����Ms�����a\�@�'N�U�D�i���e�
"d^鰧�h�6���>Q����<����?����?	����Ċ6 �>�%K�,x�p��;Q�Z���^�Iן0��]�	ן4�I)y�@��%k��5���)A���Y�p	��$������Iڟ��'�z ˱Jt>e�$N�9�M��m�M�6KD��>a���?M>i��?� ���~f�%���'h��D-��K�������O��$�O��\z��0���4��2��])֬��KXP�ԭ��:�6m�O��Ov�D�O�]C�;O��'F�mB��̚B�-p�N�%M��#�4�?�������,%>M�	�?-B�#2ĨX�R,"��x�bK�ē�?��x �������4��!=�D]#&倥D��e�/��M;,O����Y��)A����d��n��'ĔKPb�5z�%�֏�p��!��4�?��q�Z(�����OP�����
0%F�ӥm}pqP�43���a�i�b�'b�O�*b���Qǐ�{�5s7���.�������M���W�<�J>َ�D�'�����N'�p�눣0�:��b�q�����Op��XS<=&���I��<��4���t�^ }_>
d\��-�ڦ�'�41��~��?A��?����K�0�ׁ�}!�6TP�6�'���4�#���O6�D"��ƪ b���{�tY����wLӨ���m\�<Q��?1O~��kO�on$D�Rć�e�@0xf�ɪG�\P8іx��'�b�|��'�B��T�F�X3 �<w���1c��[��Qڥ�' �I͟D����'KDm�e�~>q#&�G�}T���H�4*VT8	�c�>����?9J>���?Y����<��C�$>�V�!�훹+�f�����I3��ȟ���H�'��:�:�Ϭ	��y벦�5y����*7?��`l��'�l�����D�ß�O<��qEM�a6��gŀFq�l�B�i��'��IfG�@�J|r����1$��J�iBh8��R>��>�+Ob��6�i݁跨��v	��b���opr ��e���O�9���O(���O�蟔��á��L�N��.ϻ#DxAr�L�9��Iy2$�-�O�O����VB}�vH���jZҼ)�4�&DP��iw��'nb�O�����Z�q�Dh��i�S�$�{g��4�@�lZȟdE{��|��'���OԪ;ߞe�G���`C�!qӶ�D�O"��3C)�����O:�əw2��G懫i>,�fۚg�`Ҏ��d��ߟ��	����Ҝ������ک|6v�(Ea
��M���8~bX�-OP��OR�|"gG����BV�ϔt����k�*s\�O�`B���l�	ß��	ny��-[%`����Xt �;�jC�����m6���O����O����5K����X3�C�#�>�{p�!Yxc��������I˟@���f����0�|��pm�-ALQ��� �4��m��@���\$�D��qy� �'�M�@�'ҠLsG�0YV�
�&�X}�'���'h�	�ȕN|ڃ!ԃ����+�mS@�a��3����'��'g��'9�ˊ}�,1%^�C�%O?k�H�	�LA��M����?�/O�M����D�۟��5e �j��//`�
�+ي��݀J<���?�%N[C�'4��X�'H���0���Sd4�S���hO��T���Ŭ�0�MK�T?A�I�?�(�O2��,L�;:̨PD��q�8'�i�"�'s�����"�S'ㄵ�M�)�6� c끉/�p6m��	�V�m����	������?]Jl9�&$ Q0�+Z���ٴ5���Gx���O��1�,]�Ę2���^ː=i'������؟��	�S$P�L<9���?!�'��J�g�C\�M�7f�,z44��}�`���'�b�'1�+=� H=�H�.�p�+uMJQ T�i�r�\���c���	}�i��Kg�ħ(/�P��.6�(���>i�	�b��?���?/O�8�5��u�&�`�S�`��a�e�C
!3ް�>�����?��T.�]B�iL�M�$��a��vA�����\yܓ7�$���/v�k��	�5ڰT��i�p�4,�+Zh!��m��1c�2_�<�%$VqO����R(� L��@�P�i2d��`�I-
ǆI ģFF��C�^�+<Cp|PB������ 4{���G@	:*]��s�4m8G�&w����H-T��=8���4vF@Q[���1D�ڄ��j����'�X	v�0���-C�d���O��B,��2r-P� ����kP����zDV,��������O��C�x����%[P�����tS>�y)ǎy�X����;�����e7}r��R��q�	��7mZ�'N����A+G����s��"E�>�<�a� ��O��hem3}�BA��?���h���d̦0���Bq��2�$K��\
S~!�d�~�b�21��"$��ʀ⋸Mfax�)ғ�0�#��'c.���گ/�|y Q�D��ȟ S���(Ko����џ@�	����65�����W��!�
�U� �b�Ŗ~殍a�
�t!��v�g� s쨴L�HA��Y#LS�:�j�3%�zl�����q� �2�3�d@"/ yK�ȏ��p��M�.1�b�D6?!֩����`�'���҇T�MA��Y&!��m
����'���ز�Κ�hb��axp)��O��Gzʟ��ں}hVNءM���"2�!9(��+Kj�~Z���?���?aV��4�$�O��;E�y���Ӷ^����#Ԛn�E�W�S�>�7	�� Ta{��=���S�t���$�AY��p���N�ID�=lO�����Ŧ%*�1��t
t�c�+�+r�'�ў��?�&��,��I � �
�v�K$�^�<)q�Z�� �jÏo؜�w��C�}��	OyrČ�,� ��?��m�b�p!ԯ��B������?)�Nk����?Y�O2��G��9m�h#����q�0������O���� ?��x���*G�hqѳg�n{>�	�TҪ�e�,;���y�gI�l�j�񄀔�r�'��A����4��%c�+m��5hc���I0}>���_!���h3�S�BNC����M�6II/)�ty&��$���'fQ�<9*O��3�i���u������O���I�'D<�8�.�(E��[�Ék����'�B�ӧOV6�5���|�'P�Mx��S�2rl
�d�g��qO�Ы� D ��F8>���t�6pN���t�Z���A���.�)ŗ>�4��֟�I,�M�����O �X���:;!Fa;�$Q�6��'���֟ ����+�dE:a�R�S��ѱL<�1� �%c�x�i��7��O��mZʟ�{r- �-z�ԈV�O�4i����<�M���?��)�b�s�D �?A���?����DI�!!����B�Әc�Nh����8͘'���
ϓeJ�bff�F(��d�� F�4�=	��[x���ԅm��ݨ�O��ܩ@����L����)�3�	1VS���7��������H�!��TU�4'�Tʎ乇)̗E�����HO��(���{���pէ�+È��Ĉ�A��e�r���,}����O0�d�O�����?�����H�3d9�qȑ<��9J�g��9��EksD.��}BAߘM��hɓ���<Eɠ��`զ�JgO
��}Bo
U�|�	��u�P��V<)��Q���?y���?�*O&�$2��N�x���Ϸ�
��었�C�I4J4��Q�ޱ}��<Rf+�JFzb����O������CS��I
(�vՑ��<�T�Q�JY�8QZ��Iٟ��UCUٟ�	�|7���j[-`���0�$�A�l��X�t��� A���x2I!V&��LƗ����0F��Ç'B;	��rѮˬCrT���ߞ�2�'��I,$#2��''Ƚ�L9�@`
�I�c� ��	*Q �(٢�<r١�+�\�vC�ɕ�M�1i�0����B�^�:$ Z�M��<9*O��"�/�v}��'n��.:k���	>m���0��%7l�@`�β!�>���ɟ��`¯7*��*���&^�8$��S��\>��g�%Z�R�`�mN.J��	�<�'�r��oߐHu�]�B�|ۑ>��gH�;&b����NM0o��`�%1}e��?���h�X���=�pu�Q헓^v~���fN���C�I�eyV�ۣJC>JMp��.fSaxBM ғ2>��c/_-_���HCHv�n�!òiv�'_�E�(�:y(p�'���'�R�e�Q��ʖ����@�݉NdP����GE�m�H��	%	J��C>��2⎨~b�\`��8<O��K�F�6Y������G�M�ua=�����|�Њ	�^��7垏g)��Чe[��y
� << ��D�jK���,l��� 7��ؙ���ӮG�n�I��:V��{�dE�a����m5���	꟤��̟�A_w�R�'���:(�L��*I+!�)�0���0O&�sħD6
4HЦ�y|tа�ȧo!���6
]�1C�#B.�h@���
 n 3��'�B�|��'�����:=H^����V�V�IQ��I�Y!�d�
[%�1��.j��H+��"]1O@��'e��
��b�O�D�,��=3 �E���)I
ɄE���D�Oj�2��O��db>}JC�0T�F�H�.G�~⪍�F�h��r�&rjXด�د�p<!׬�A��P�A2U���҆8�
%R�ǹ\�3T�i �x�(��?����D��ҝ�Ć��1�JA�kݴXd1OF���R�KtN�8`Ӑ;�2Cv�T�*G!�d����I�C�0�0P�wjH%َ}�W�b��E{��)@�u8�x���\=�9�tk�")�!��0h�F̓���b�H�sDJ��zx!�d@�WĒ�qˈ�H�h�����5ht!��3z (�+�J&RuԴ��$�(_y!�ĐY�y��3V�:�E�Oj!򄈨;��0 ��g2�r�b�4*�!򤝀7�8� �d��q`K^�!��ņ	�.8��`Ӕ*t�Р4`X�3�!�Ě�-�ӗ��nj�0���T]!�dS18��m��_�s�@i����-	G!�dϩ7L���+��R�㗆A�B!��*u��t�k��zW�:!�D�*MC���� �b/��r����!��K�Y�rq7�o�,EbA��;y�!�]�}�dX˒l�0)��,8����!򄄁p�\ي�W�O��<b�$�!�dA�AV$i�I,EU��)_	_�!�[Ze�i�E�m�8{�V��!�
� ��aK�'Ez9�FiϔO�!��ٽ&�^e�b܉}T
�Q�+D�!��/���80���@�)�F�.q�!�"T��8J�IM�I)65˱@̷�!�۹]��i���Q�P|���d�U!�ܩu���f��<Q�(XP�I.x!�]�2}���̋�C�6�"��Y!�!L� �7�C(i�4�3.�Y!�dZ�lr���E?l�p�d�Z	E!�D̘z�;�޽oTp�i& T��!�䓣GN ��䊟5|�@B�R�!��1�|a)��Q-(�v�h�(:BO!�/�tų�aY�g���SH�9k!��N�8K ��[N�"p&� �!���3����NN�ut���増�=!�D�W!��J�ƣd҈+�L�-s�!���:U��5 �H�98g�X��(L
!!�� *=:��H�n��p��U|w!�$�P�̸��	+�y)T CbU!�dO$�*�[hZ-�,A��1'�!�Ăk�x�)�o�<֌�VPc�!��NPցXE�رE�z�mߐ�!�$�{����/ldp�o�F�!� �~���͖*Q\�0�!/�)�!�ʜu7���ŠM�\���.�	(�!�d
��9��G�2p �gٲ\!��,x�ʤ� nO�N������ȥ6Z!��.Vڒ`�Bgߵ#���a��A!�ӲnĦ�����$�h��5�!��P��h�ٍW��ړ�Y�F�!�M� �@B� ޓ��9An!�$*]�99��Y�q�VŅf!��=&<-B��&��̣�c��^P!�� H�! d�� w�hk��^Ej(��"O��Q-̾�$���-*�E��"O�y)��R:ʢ��#j��;"O�E�f�K�7]v(����C�� JT"O`a���أR	� ��U�<��ܨa"Ov����Н�h�*FHē�R��e"O�h��H�}5�л&�݁S����U"OZ!QU ə�d���K�/[�|��s"Oh�ab 30�x��w�ޤM�%�F"O�%HҩFt*��Й��Q"OΝ[W�W�L��(6j�'X.�C�"O��ɤ
��D�� z�	���`Ad"O�MA"+�A]��b�B�C�K�"OT�##-&#М����{���&�'��i{�収m���Y�j� ��]y��W�B��4^������]E��)��	�C�`��&C��>���^�&G�px���T�>a3�
N'V����V*������:��g"r��:s�܌@���4�Q��/Ĺ�ff��S���Y��Pp��g$�e�e
�7��B��λ_�z��ȓR���g�����ZB͝T7���O|�5��?�~dW�G�`,$��E�6TF'͡MZ����6���	t2��-��3\ԡ��C�$"��X
ci׀.88�M�z�dI f��E~���i4j��%+�1�b�:� �r�t���
]��Z3+�gi0���5+�FI�>@��8p��!XX��Y��v�աk����v8����o�Dr��(a�^�af8�)�>ѓMG/�*,sC�YL9���q0B.U�L��/��P
r��$,U6O��E��0H|���DH�,8���M���䞮&Wܐ��V<W�(  6.H���	�Q�l����B��@����$���~��;:�a���$���c��5y���D�^!1O���@�0��L�!/
_���Z�����'�ܭa��6#.����J�o����b�A�?G$�(�\�K�υ�a^�'�}��N�x��Kd���x����ϗMn����B��fX؋�����O�pC�_\���ϫ �6���D<s<d�PCc�?	�a�9̄�1�K-u�Fa2���K�'����ƈ�{rH�aŊM�/`�c��n쌙�����K�j�a��]�f����(�$MY`�R� n��">i�$@�@d��!̼��~�<ݘD� �%���C`�|��Z%gL*Z�� �@璮#��(�f� LLĻ3�d� �Ź7k�K�.�86a��2�1O( ��ML��Pa��>ga u��-�)bք�*3��8	��0:�B�
�-ڄP��+��b-� ��f*xt��ئE5?�(Ҋ�0=�0n�6m��v��_���e�n?c ��3|4��ROU�mKvh�D�V�'Tآ�7*�����:y����'�@ʖ�;�P�.p��e�(��D�{@�DxܓO�Z 8m�Fx�;F�@��T̼a���H�#W� �B%��I��A�,z��J�' �=�"#h$�c�<�&+,(��$`��W�.T}  !�I9w-��*�dM?R 4I���Ģ>1S�J�F���!AP�tll�DI\7��h���1�Jq{�.�i�������(o��D��i�Y���8LOfY��EK�-���2�N�:���@�OLo7�ꅩ7�?J�fX��M[�m}��0�J��h``���=H�S�J�S!�DR�",����ʙ���㠊�+�$d(�J��਽	�Z;
�1O���JJ"xͲf2�<�TK�:5��� �Wx�b��';�\��KA1����$�B,�6 *� ��\��<�<)�(��v�=7A�(�,5�6g@�1�k"&TZbh�bǒ�F�x�F}2���b�RĢQ(��k�,�i��q!�A�K>���Aŋq��93@�;B�t���S��T��gA}��� ��Cȕ���T��a�a���ZƦ?R.B)
Sm�L��TҁӪadJ�ce�dI9X�B�Bpns�R��gE>q!�{󄜈%=th�A�?:�Z�s�̘�L�ȈZ�K��Yt^��C�T>#�1O^��G�DcG�� 1�H�`�ß� �����:�����'qbb�h�;f�1b.�1G�n�;p)իMZ��<9t!ŋ�Z�c"E Fa2q��\̓A���(6�ܰ28i�lb�(|G}�'�&��X�8h�d+"H(}@'�qH�Se�4`�j +DK�t�Ji���u��Lb��4T���	{���� �=9�F�K����z牍Z����7dU�d����3;#����yKFc���dX�O:��tg_,�.P�\ �dH�P�:�"~F���P��AOM>Ĵ`�S��8`�t�ORH���Y�H�RI���9O��;?�X{����L��"�^��L�'�1�2�'�&m���&s����%��:ƜS� ���'�ƝQ�(�F�Hl0�g�a��S�:Id���D�TK�[����J��8��L{����L���Y����
p��3� e*2�7���Q`,&���2#�A�b�Z�s�;P���`B
.s"��T?��$�E�D���Qi�">��%q�s�������*�R�O�D�x��Q?��?!���$�.��������k�In���ڠ)d����	O$�Z�UI�5V����м]�E0%�� ���ɬG��CD��k]v(Q�F�L�">��@�3<��u�ۮC�j�ju����r@X�8(�����!�hxE�B�<A���c���RV* K�r�YP� �<9Bf]%%� ��"W�E�
qA����h��HJ�L�\��08 ��!'d�i#W"O ��C<S�l��5�S �(��#
i0�11�F;C:2u�B<��g���6,�G�_�
��|��,�L�\͆ȓj�QŏfA�B�� �3q�EѦ-����$���{�,�_�"!"b��rU�l�E�3�hO`!Ip��Hƈ��b�L5j�v`´�JB�X�YҸ�*�ѷiF��j��B�<���+��1�M��oX���6��Ħ�g��fB�H���ZYFp�$��OQ>ט!E�z��Ǎ�e�mˤ�#�$B�	�)�,aP���0c�䩁��3.5ܐ�v�&�?1�C�:8��<�V˽~J�E(�I�R[H�P�[9��0��=�����7E� 	Vb�W�L��`��3v�B�҇�E��zA�DL��<a%T��=�S�ѭ/��. �I������ܓ�`�
g��n|sf��0�0M�*#��͖���؂2�2����~�<!�"H�&���,�QaFm�Nr�� �d�OI"�n�f����)��y'n�4-`��ːoV�/��aW����y�Lȴ��t�h��;�(1˂&ʓ���5�hP`�]�g���ҩ�C⟠���<�1�a�<cLx%KV�/LO�2f�f<$)��]8n9�D�?�u���4H|����冣�4��tKI5>)H��DY�jHu�\��#�X"\I1O��'�H����D`q���A�Z~��DX�s���:2��Sg50X�Q�daKO�<��E�T��4c���]7r�1�i�.��!I3$_F�na�q+8w�Vy�bM�PˉOf2���w�h(�v�X`p��I�%����
�'�be���W�^4�ą�=W�&0�6!W
�>�9��T#�H�q�b.�bd���7^c�Xa�7&��`� =�:\:�<lO ���C���Ѡ{ր��G�	�lzV�Կ%��I�}\��Ѱ��d؞p�'��uh� S��	�H��H9�ɴ�XpK���L�O���R#�	_�$$�4K>���'�跖�1$�L��'�
qF(�[d��p	��OQI��3?��ӛCR:�Y�/��6�[���P�<��,$C�0�ԡ�(�ܑ+V$Fh�aq��!�:��1(�&����!;=��4��H�az򃈭z�X�A�ST?!6$��Ԡ2�M��ԡ3��^�<!���>C���x�&ͣL�L	c@$�A̓�( �(�3b��~%���p&քYذ�bQm�D�<9��Wy�$���<��LH�73�@s��0}�#������/_2�1�D[�~q�%i#L�&7��B�ɡw�D8{�׵Ey��P��B�y�C��B�\X��'��`ѫU�w� i�ՀU�B���ӓP��i�&V��hK~�s���,.8+��ξ��C��-a�x4�aE�n�|�ʍ3mrb�|�ƕ)S�����7Cj��adHKx�Y�3�ʜ7��C�	XXJ�F�Y�ʡ�R�[�6"����L��T?����F��O����9"��Y�S�{��ء�"O`Ȼ���4�2E����/gP�����;�<`J�&KDX�P� �Jg$���	0e��X�d,D�<Z��x�D3 �Q,%�J�F�)D�X�ˑ*)0:Т�Хd�z�qU�$D���Cl�T�Vĩ�s_��(U>D�x��@Z�q~HJ��O6G8|+�:D�h �
�(Wƽcb���d����3D�8�6͎1W<�{`K1�xxE3D�X����	&�8�r0�
0r���Pa$D��؅PWƶ���ʏ7����#D��B&N��y�}�pM�r�~(� =D��9gKO�z%��/G7\��c�O D�H�s(9x���beGk�J��5#D�hS�G�2q��A�=N�J�cL!D�� ��sB�^���yDU� '��s�"O(�,A��h�4��@�d@2"O�3+)u`�Pᣃ��Ҵ:""Onq��L�;RY����Y�"հs"O �6-�6u�Pp���_��:4��"OIcэ�6_�B�"�mɑClB-@"O����u&���vW7Ee�E�"O�(�V��h�@a0�x}ztp$"Od��$Ř�G�f('�\�YX�a9r"O~��Q+K�&�z�Yģ�)/G��e"OZ�Q���U!����@�3V�kA"O<(˶�Xx!��ă��*�t�"O<�.�4k=�`	P�Q0g`2*Of=Jf)�Y�vug)3T�U��'��*@��$?�T�Wj�R���q�'_�H�eD�<��ř4J��I{U��'񐕛u)�?���{d���O��Y��'�M�*��F¬��sa��^*�*�'+ u&����y�DV4��5�
�'��1��)иKj�"���>����	�'{T(Ar�:><�F�K9�Y��'Jia��B�z���:�/��$��'�<�X��S�NA�0�(U����'��d���G�[��E�2#OH�m��'�z5����?5��j�ŰA�r�Q�'M�P�N̪v���f$:��p�',�T�6`��3��!�v�:�͸�'U���,G��Y#�� 6�����'QZ!���D�4<�(����-K����'@��v��"z� fR-9�~�Y�'�jqj�G;L0�����"O���
�'&=��M�wzb��P����R
�'R$�6_Eb63��Fˢl�	�'��Hb"O(nlhzU�Q+�lI	�'�pe�v�IU� <D��ya���'��쩐r^��b�^����c�'�*%5JT���N&r����� &�yb��w�-Xq��h�D�1���yN��W�1�O��bZ%���ybJߨ����& �r4HIK&L[��y���^������bły�%�˱�yŗ�C$�,i�/��% �ÈA/�yr@�c;��I��&�"${#���y���sN�۷�J0tD�r @��y2邇�,k��+|m*�
���y⯍+|
�Bi��"�i�ѢG��y�'Ȩ�t`�@�r{İ�m���yRn2ŀ�a��Z2j�z%��(�y" �b96E �닼c3P��tǌ��y���&8���6�73�Z`($E*�yr�6U&�y�n��(��=+FŇ���>��OL �xC2Q�3ժ7N��蓨.D��PoFP�Jf��/!�pY�(D� �wM�3ˈ�0mʘy�d]`*$D�l('_�\���F���R�骁�#D��H��U������Zw��ӵb?D��ȰgO'���&�L�+���Q`<D�x�U���ITDX���n͢1�u�9D�8A�)� g�p�@
Ji����6D���D-}�|�)�k�F��De�2D�#F�Ϩ
l�5S�AR�2 (�5D�<���**
Z)c[�W�ؽ�`�>D�(Z`I�j�v�Ȧ*�?���2�:D��(A�v݂PZ7꟪!������6D�� � ��<|��%.�2C��\�"O��)Q
�l5��p�ź����F"O������JB]hS���ԬѴ"O�I�#BJ�d���9vYX$"OH	H���%� �����$&z��"O�J�J�[|DL���Y���"O4e:�+���Qz���(l�ly�"OxY	tn�A�a�1�T;di9b�"OXi�e����A�F	f���V"O�mqf��,�p6��
0RLyq�"O�-cE�?rf9pk��c?�@�"O>�At�	�4 �Y	£�28�nm)#"O�J�.��L�q�O��dX�H5"O� ��ƭo�0m�C�C"Rt�L�"Od؂�5{�a�d¦9n$��v"O2Y�!##�\)@�B�kU���p"O�$�Ζ8t.�i��ӁtCN�qA"O�a(�)�!=f�]�5�Op��k�"OJ�b�ˈ���7�4c$l;!"O�at�B�F��	��/\�OHZ�J�N���������E����/'#&�i���yR&H�+"�BeCL� x�B"ˁ�y�b�!T��욤�����Q[�Py"kĎG$���s��%5�{�Nz�<Y"���-�r%8��Z�u�h�ꤤnx� Dxb�00R���DG��e�"5�yr&ĿK:3`ݢRT�iC�c��y��G'[�j�j���L�ym�&�y��'�NL� +��A�<��'�0�y��O�+�Vl�k�Ks�9ar�M!�y�@��|��o�x�N��P�ִ�y��A�KN��� \��W��y�ؙ2(<S�"	fZ^<*'�֏�M��'�3`o��oQ�����+��m1�'�i{3���%d�
E�
����'~N�0qL�0A�!��@�'ln��	�'q�eY��W�*��dPq��W�`	�'��8���S�LR\0�D-V�.8�'Ѧe��3GP"�f�S�6ʺ�[�'��`�qɄ�R�F] �ě)q�|��'7,4	�HҫA��q��⇿ P(p�'e�����'>��L�a��8$>�\x�'T�3&Ǜ%�hhI��!��d��'���Q��N��'.��m��'����gJk\�a�/�z�P	�'�idh\�x�ĭȆ��@հ�'z�Q"@�H� X���e�B ��'�z]�!]H�	2��!V�̀��'�@ 0��E�F���釠b ����x��I�(�����YZ,�u����y"E��y+ܔê�5K��|h�����y�,~�����Z]�x������'�ў�O�����Lf��a
��P�b�4�P�'��(�ZM�����Bhc�'H�ظrJ˴|�	"��˸c�,qj��:O
��գ�:���$g3,�4j�"O|e��nKiʚ=�;I��� U"O�Q�@�V;&dxxY������'l��`��H�6&��1�/W	i	�DzB�'_�ܨ5�A�b�;4B��T�{���2��e��i� ��"���L��`"O���c�& ��P m�Kv�
�"O�8���." �8�E�>]k^Lt"ODa�ȃDy8�q1�X,Q:-i"O� �����M&~�NLR�)�,O2}	#*O�x�W��j�αP�!Up\I)�'٢`j��4�+T�O!Q���		�'u`1�Ck�8F�.�8Fl�D*�Z��6�S����j�\���߫T�t�Rӌ�
�yb	D�j��!F��S��r��ɬ�y���#�l���M�x}�ħߠ�y�F�{&�d�Gi[KAB���D��y�3h���'oA�J�<�bް�yR��"^��xǖ�G�ly��˽�y�NQ�:�p�ch�%=��ݻA�̤�y�/&-��`�`N�@��xpm���yB��0���!O�1����*��y�+��r�P�!����%��h����y2� d��T[R���$��DC ��yR	�#+��h �-�� *�i%┷�yo�x鸠�ri^�L4�G�.�y�f\t��F�9|N����AZ��y���MCt��Ȍ{�Ne!��R��y҄�|D����J�i���5�U8�y�O�\X%�b�17@�a��yB���L�)�f��2���	�y�H�o������6�)��P��y⡂ryXi&���4�d$��Y��y��JC�D�IfգyF�($IL-�yB���r��3�[>�$ЖN��y������ۢh��F��Qp�Ț/�y�DD�JITp�������y%�Ǘ�y2%<L�J)���I2b�'�y��ԣg���R��-)7� �����0?�*O���g��@R�H /=Qot�"OZ�Y�ҹ�����ɱY�`(!w"O�a�e�Qݕ��P�{��83&�G�<Y�dξ���� �X� ���[�͐E�<���	0)v����A,S�ċP-�j�<��?��PW��lܬ���GL�<�1	ߴ$.P�DO0hb|��*X_�<�����ZvD�Q3���.� �U�<��+K�iߎ�x�e �w��!�ɖE�<Y��ڒk��m{�oޟU��d��u�<!
��V���!�J�z�h�#��Y�<Qa �9&b���λ_�d���V�<鑋E�n�x�q�K�%���0��	R�<����o*��5�ȅKn8ѱMR�<�'nƉJ␩��|�b�)��r�<9��D�Z�KcBżFތ)���t�<��M�v	4�b�B�D�rQieMMv�<��M�=����nB�vu���Ee�r�<AdC�~�h\H�"�4��8��En�< )�$:�E�ĨWZPxK��B^�<!�3�Z���%{Y��2G*A�<QtD[��DT�N�h>�S�X|�<���X��6�ܘ4� �3#��{�<�jF�1��p��P9#�
_�<!���T�9A"�7Bz$� V��A�<���Flᮨk2N�f]�P0f��h�<)��5\�j {�S�fm2Q��fCf�<��ݸ<2�9��.D(.(��X�L�c�<���P�pxE�٫g�B�В�`�<�⫝��@ź�Kר-t"�!%�^g�<9큮!��Ja�էB�\)�`�<�J%1�0)rM��U?z�Іs�<15�s�q��'�X�
c�<��:~���j�UIj��uU[�<� ��@�����2�(�W����"Odѱ�l�4u��A"'E�E�¸G"Ox��DF�3d�0�£]<	 �xC"Of�y�c�:,Y����$�	i�T�be"O��X��4���â�(�(�
"Oڬ��ˋy�nl1�/�S�F�p"Oje�a,��U����JB���#"O>�bF��G��+�B�+aƼ1�"O�Q1�&AnZM��V�]�A"O�$JքؽP���a�@��s�&h��"O�E��KS�L���eo�-�D0C�"Oj	࢟�T��ʦD�/x�2"OB��T��7U�]�$�<x}�"O�� �X�W�D���t��'"On��O�pO�t�UI��%�[�V"Of0 �XO�"�G�K�0�F*O��q�逑z��X ���4Y���'<�4�!�%h�Z4;�L�<WَL�'e�QA�녋b͘�`�Y+S��ē�'R`LP��è%�V���f�=q
�'(����hL�zuv��V����`��	�'8�8�oM8n��tk��T69��
�'���z�H�4H&4h���K+)����'���B�f� ���i� \ĸs�'�����˄!Ξ���Z�$��
�'E�Qdq!Dh�G"
fdQ
�'k&IJ��ܢ+��<�d;��]s�' :�P�E��v�����@oM�5r�'��sD�#/pds#�/c+�	+�'��Q�m� cH���bE�$-���'R�*F��GR�����0d��'v6��0莥-���@"��w����'m*��O�=-�xA�A�h����'!`p�v�U((��%Hg Q178����'*�X8�Ƅ?a�`��F�/6�`(�	�'F2�c�͛7�*1Z�	����	�'HL-0�Nٙ]�Le�o�i4m�	�'�L��֪�4~�nu"r♐��r	�'8,��c��4{<�����A[	�'^@,�B�F�"����@����x*�'�����ĢPb^�٠f��h��1�'O�#R�2@{��k𡏳�*�P�'��U�fN� ����j=u:����'vz����p�P]��M�?x��c�'�I�&A�=�8�I��5��(�'wX�dl��n̜ Ǧ�}´��'�d1��`
�̌�F*݄p~�i�
�'u�r���)jdc�o�|F�	�'`��陾Db6��5��ml����'iV�R��ܚljpň�âW��I�'�$�;Alݴw4�G� b�9P�'Uzq�M_4)j��vG4i+����' ��TO�0B&Y�����e����'m�u�u.��_,��h�pَM��'���r�+�G-:�O��9�p���'ppQ�k�[b�	�MZ�r�'UȔRh��d�$M��b��v$��'%��g[�j�rIP K
����'f�[�_�G6��"7Ϧ(&���'�Xq��T�`���v-�--.p�'U��DN����3/�O_�i;�'�~�ض�yZ��I�c�22@�t�'�4���;u�h��+�!0nf�'�x��LܝL� �H��$�"�K��� �qY!��!.6��]%J��""O��)rF��8@h����Ϣ��� �"OX �����Yd���	�/��ѓ"On	C�su��U�7}m�"OҤ,וl�F�!���W�L��e"O�A�iX��[��R�Xk�}�<�1���EG(\���̓<�TE���U{�<	�(��e�ƴk�G�8j�p�F�t�<�#隿q�h���u���Ze@Np�<n�%^y���C�N*���AF�
B�<�Q/^&	� �Y��$�\U�Zv�<i�T�g ��:���#IoZ}�"K�p�<��iQ�=Y0���>��Q��Gp�<�A��j>�����Q42�Fa
 B�T�<�"�J<��{/B�U8��ׇS�<Q��0X=�S0+�*�+��N�<��l2[$�n�-"�B�Ka��M�<�cGУE۔$�TL�d�tHs��
H�<�v	��<��Ţ���O�6�� �G}�<���57,D��G�`V�mj"��|�<դצsm���AO�og�,*�D�q�<���&Zm��X�Á�>���+�A�R�<�d�72��u(��_e�e�P��P�<a���~�hڇ�@� 0�]#�I�<9�mZ1j6Q`��_�H��ʅ��@�<��bͪh�⭸� :càQ�Q��S�<QK#,/�� �B�55��D��	O�<YQ�C�VT��!dgX�XS���K�<IFˆ�@ۚY�p-8[�� I�<�ǏڂZ���i��Y�U��P�c^P�<�C/�&4���
�Vy2Uz�s�<���VZl8��_0���S�<Y5e�
&)B�.�5{9��\N�<�B���T]*�S���u�TB���s�<�c�۱a�p��&EV�[H�����u�<�U�_����
n�(S��E���Wu�<)Ef�?��5������ ��q�<��LX�\�V	d��
Plxs��x�<�qj�.I�D�,�2W��u �Gu�<!�m	2�X�1sk۰�2�+�WG�<�N#�F913��Yw ��w��y�<�r��oު�ґk\ P,mzծu�<Y��h>����Y�r}"�bKo�<�O_tA8�K1�߿a&�tҕO�A�<�f�9k��JǊ�"Y��Y���U�<�Ќ�;b�[&�.��T���l�<�E�	��|H���U�&�a�#�T�<��K8M$�h1mȗn� ��u�<�6���'�L$�1
)v��u*�o�<)3n�W��:ňM�A��k��s�<YV�BК�j &A����R$�n�<a��2&�%k� ٧���P�L�g�<iCl�,-sb���^%YjY�ï�}�<a�)�Onu"Vk]�UP��2hu�<a��K�|T�� Sֈ-�7%�m�<�e��!�h��Tۗ*Ɍi{#o�`�<�JQ�*=��@R�ks��jS�B�<��BŲBT�:���A�X��J�}�<3�C�.1�� iD'��E�w�<E,�G�@�wLJ$SĘx*#GJ�<iԩ[�t0ѹ�׹o��mr��[�<q�,�p���g�2.\�n]�<!͞	;I�|@T7%}��a��<�GK��)��y+��C�����R�<� :��榆�;�jHÀB�&��lI�"O���m�uz��"�"(��H�"O�h)1��G@ ���A©A�6�B"O]bb�,{l�	[���¹	�"O^��7��qB*9)�/�%(+�I�"O�M��ʊ�d\9��Pp�d��"O��$-Εi������H^��C"O�Ԑ%NQ��@�CeRL�j�"OB�8�/�Cpz�K����2�{�"O�@���&�X�r`f[�|�x�P�"Oz�1bi�Oo��ðĊ���e:�"O����]�|�҂�?�2�2#"Oft�P���Z�Q��Z<�(�b�"O�,
�j�|*@y��J�qg8q"O ��$�?�\��hMOt	7"O.�hHm��:�i�{C��"Oji��%ӞF��t�ӛ13���"O@!���?[2p��@��Jx�"O4P�c X+��;�٘d�̐�"O���B-^b��̓V&1\L�"O��c�ł�2��� `jmZ�̂�"O�q(���hS��s�	�n2Ir&"O�0Z�%
�z�jϐ�6O���W"O�� f�5�P��ş�(<P%X�"OP�SS&�4b]bѫcW�5<�dI�"O��p� �d ]�B!��p+Vmj'"O���錵|�8rb`&��c�"O���3��73���`M�33S�)YS�'�ў"~�e-=OUn5���9g��=�!#���D'�S�O�<����f��%!ƍΙ!��r���'����łA�fP����>9��)
�'e&�F�:Q��Q�$���h�	�'i��ˁ&Q!Ox�%�F*��kR�,A
�'��<��OU�f!��k�@�1��I��'�H� �&x�V�֗��L>I����> Z���K0�4LC���,�!��S(��95�x���k#N݅K!��\��h�������mÑ��O"i �*NC���YƎY�x�̭�G"O2H�Q�:���[g#ü[���0 "O>���7
�樘4�ώ�0���"O�Aё@N�l�Z��v-�J(-J�"Op��NU� Zn��"�_�<�`��"O�͡à�mˌ-xc�S�L��ɠ�'0!�ĝ�H�*�ŕ�L4j�-� q�'�ў�>�scS)��q´��%�i���,D���סI(,��{7�֙K j	˔,D�L�S"�6uL@��@ur@��-D��%�>x�q��Њ�<���`7��c��@hs��
M#�����	M�R+2#6��]���¢U�<@�0��/8.�A�/D�@�2���V{��?53�	�C�Od�=E��4Ojq��� ����ـ�*#��lX�"O��(�d?ތh�JxizW"O�c�H����Uj
وv���R"O����%	���p4�Ս3�ZH��Y��F{��IF l�<L�g"��:K�ܻW���da!��8�N��j�
6�8�F�](>!�ݺK�JՋD���*<$������]�z���$��B�`���>{��a�ڝ�y⭍ 
)�Qɓ�\��t���yr(� 0�v����B�7�y���l�P�c���Vi��
bF���yr��� �eFU�\AqKH��x� |ɉ5�I�ba�zI�6>���"O����'@�!,���'�l( &"O�A:wn�2I�*��0��$������!LO���Nڍ2M��7�(Nh�y�"O����蝆iP"��8dŢ�"O4��)X8�ZV�X)I
��Q�'�I�w3�1rԠ�P���FǄ�p�B�	\,�}X���<$�}���҈U�y�ɇebb��J�l��@��߅=eh�O��=�y�L݊6�J��1�*�>��G��yB���"̎� Bϊ>"FL�����yr £@%���v�oi< ��y.@P�Ȑc[5e�X5�f���yRLW#\���AP �Y����k��x�'An�H���Ϫ�`��0�؅h!�דc@ +3jB�y���pr(,,�!�GEQ�l*�"�F���42�!�$ƳpC��I󡔃n qd�M0F�!��N�d�:xe+����+�h�G�!�Na�����X�P�ʃ ĀY�!�DL t���#��4X��z� ��$���;O�zU��EL��g�2���Y&"O��c̔�e�ڬ�&L=,B�4�$�<YO>�˟v�b-< ��+4h�J_��C6"O�$���
+1��D�7��Vb��"O�)rŊ��-�8���G�h ��"O`u���g�*-0�HU�xfI�"O� G��$ꤔH�GZ$eP�1"O����n+V��zT�:X&]���	J�0、�zVE��%�"n�⼘5�8D��0g�3L��%�G�d��e��!��������F#(xa"h���'�P-0�f��q�kЧ8Qo���'�X���a�#6Tp�fTB�t	��x��'7&��qB�ѓp2|��Z �yLK�%6�|[�
L<kXZ�@�h��yb�рa8�����0�h�S�yR�>z�.i"i��u�|��C���y�I��AJ:pRr��Q���y掅7�NU��gQj�8<�^.�yRş�^ώ��@AE�f�<��(��y�,n9�����,Q����!���xBI�(���S5�@9i��� �N�'&�!��"N���D;���� NG�!�$_�l|����LZ�+c�=`��@��u�`��7E9B��Bֹ͚��ȓU�\�W�sC���c�m����'nd�[�'�rQ��쒎g�����'�!a�O0�|�c�G/[�9��"�'.�e�r ��t%��,��D�s���'@��&�Asq!�f��
2�	���?��*��.uX���O���"O8:g�܀� ���+��1�h�"O�U�7O��JܮLZW�B���"O�᧧I��qv��8�r� "O��ʁ���T��WiȍQ͎� ��0LO��:��k��!s��>M�j$c'"O��qK�����C�D�<{x���"O�����ػ8�H��އ%pX$r"O<��A�1�
1�l��XQ���"O6�J3/Iej�8��Қ#?��u"O����mΛ�)���� ��"O���R�O�@�6<����
>	�a�"O,xyAk�2��v��)!��}� "O� xɳ׮�͖ш0o	�F8�"O����
O��f��V.��lX�҃"O��BQa��HHb�,{��x;�"O��{Ӆ��wz�[��f[�D�"O(k��"òHC`�=����"O �r��(K���Q4Ꚓ!�N�Ӵ"ORM{�eҌ ��8'�D�X $��"O��:A�^�X�\9�߄aj�80e"O�j���D��a�ӦH�H�ޱR�"O�\!c蛂Aj��y�F�"�	�t"O���C!"����F �)�\"O��/3f�r@��΄��č��"O���hV�k�H�RX�v��� �|b�|r�7o�,�J%�ђL�-��Ȟ�BC�	�<��)�F�V�A��Pj�C�yY���4 \\|p !�@�!�B�1bsR��A�KMD�����n�B䉲���qR��h�L�=1(P���d�������=b6���V��ъ!,0|Otʓ�y�OӦ/F�:q�E�I-�Ȣ��&�y���}P��2R�
�A�4�04����y���(��H�AU�<�>�TE0�yBa6]��}PL�7Uu�O���y�MÖioT�5/;Q��yiJ8�yҀ��]C�i����7���*,O��y�J ����ߜn�q0�jд��3�S�O,�lނ��� ��v���'�b�AT3+È�aգ�����'�)�A��'`��B~�BA�
�'�(�C����)��p`�	�
�'�%!���.G�1`�K�b"��`�'���C�O1w$$�����8Y�*y`�'DB�aV��	�l�gϖ�>��99�'�B�{�ʟ{�D�&��5BCX� O>����iý,��æ[*9���#��.e!򄂯ń#sA�#�%b��!`�'+ў�>�! iD,k7���eM��cQA�@%4D����K�\�f�I�@�s;�C�$D����`�'^2��j@��s���"D��H�C�t�`�
�E��|�0XB��O��=E���E�Z��l��j�V'�u���:�!���.N�(�3��>���"0`��W�!�D�&r�� �J	)����sM��P�!�S3Jgz鐀&x�(�/U�1x!�d��Fؼ�Q�ߡI�*�����/{t!�dN�Cl��BD�$9~t�!�i-m!��*(�,�#f��Ja��C�_3:Y!�Ӄ+
H�A�BԿ!�D� ���WS!�\�+Zp2�l,v�z+�n�2$�!��$(�B�RSLΝs�Q7䁀��'�ў�>�8&/�2+�Liਖ਼3^�$u3��4D��[p&ٞn#ny��-�5T$u�f(D��#� E2�J��t���)�Y�(<D��V�[�ie�l�,R�AE2QJ�=D�TWiEff��zE�]�C�0��<�	d��k�ƟO�6S�ɝ�xK�![��9D�0���ɯh�#M����Ҫd�!��20�pgc��*C��$	�!�!�¤=��8 '
8l�13W��J!��?D�%#�oX	!$�82�Ζ<�!��,����$��Ya썡'S!���/C�,�'��'`I�'�иM#!�D/p�3 ��"3�j��tm��
!�o2��r�j${�6�D��u!�� =������!��@[��B���"LO���՚n2�lD�ҶXs�4� "O@{�@yrܥQ,ɺWkt)�"O�!#���8(BA�U
n��#��'_�d��Zy&�Y�(�P��dB��FS�!�dK�=�BP�'�@;_����*9S�!�D�+lT�"df��$xbń�!�W�	�T	J%J<"4x��,�k&!�$@�3�6H֏�� 2��`,#Vk!�ʃp;H�Pr�`S Z&�ջ5!�dH�H`�2��?4AP k&��3!�D�>���hׂv-.e�l�3!��'x���p���#z�jVAҎg`!�$�;1�R�����X��!p��M�9]ў��S3�2$)���Y�r]{1�$m~�B䉬~T(P��5L��`�FwhB��6?�~���ǾQЈ4#p�"�R�=9�'�d��C��,w�8S`�]�v�`M�ȓR����F�]NX�bVoߋ=y@u��y���B	Ӯ)�lt�F/PS�tX�ȓ�e %'�<tb��2�֊��Ą�,4ƭ��E��N�'iT
?BNԇ�>�����`R���h!m�Nz���?�zĭ�w��L�MU�^H���j Ys"�c0bѡf(ӕ"�؆�IH���́f��@9 G� ȓM�
��T�J��
A�ʛ�T0���s����R+�mD�
o��ȓ|��զ�!�h�G��z�5��3�&,�DJ�B@��� ���iO�	2L�S�,���cX�S�̇ȓrb"�T'a��\b��0#�~t��6<�(Qc�)G�j�I�k�� ��1���Kм	�q)�#;|��|%}�4�$̲a��ND�@���wp�y(�֊s���H
0���ȓ02�x�I��y�g�J_l�ȓK�`��ƀu�0���%$݇ȓGT��*JДI3iP3�`@��t_J�7�
�d�:�ǎ�{�bA�ȓ2��s4M��i�8eK�/���ȓ$�,��nW9 �����#�0���G{"�']JH���(��A��/"�&�)
�'�Ą8Bm#*p$-C��ճq2nb
�'��{狏W!��zD,jQ:r�'�vb,� b��4�V�c	���'lX�ȓ���P��3X䈰�'��p��b��(�q�ٛS�R���'h> "�>$��|��j�EP���'���`TfD�O	�A);	��'$D@���'�� ���7E�,r�'�f�Zh��7�����N�+*Nȝ��'����@��:�Dѓ�HYWδ1��'پh�(B�L���S�FwV���'T���'1Cc�0Y�IԞ)��F{��O ̹H�H�%fK�J�K:�P��'3����2`�d�lR�[�@Ap�'����7!���d*۹W��(�	�'5t���G%E{�a�@Ã:����'XB�;�C��`P���N�2�T���'=X{�BL�::�R3h2uz��
�'"���%"C̀ �����V�P�P
�'6�q0�d�JU��kD�� �v@a	�'��9�I�#}�>Dz�O�F{p8���� ^�1@�Q/w
@��7:9�6\4"O���AH�%;v�R�Y lێ�a6"O~�0i�	J�����f�2T�$�{q"OB�
�*�- �vP�(1�� I�"OT� �JҵZ!P(�B!ۻa��ٰ�"O�5��D�)*������!*�y
T�|��),6"�p��� .�q .�K�B��%Gc(���L� J��u�A+�6oÊC䉍d��������J⣖�vw�C�'�H�a)	�.���Z���h���=��PF]�"!+{H��۷GD��j��ȓiŲ�����K��H;*f䕅ȓ*�~�f��7;�@[e�j�ֱ��:h;�I�M�`[q-�h�}F{��'9V�q�dE7%"�"�)�?.T�H�'DP���̗n��(�5�C$�p9�':�ia̚�g��H�ݠ|+�Ku"O�����N0��B��<E3���'"O�T(e��3�f��*[�&D��"Ot����Hk���K�A��u�'�ў"~j��#jkʼg�S�T��ȡ�(��?9-O����g��j#�9�|,S�I�`����^��͢e�ĸ�F� ��ϕX��ȓeN�� %��, 8���܌��A��Q>��wK	w��U��dB��B��ȓ4�|۰+Zu��ݺP�åY��h�ʓ7�!�Ǫ�\�lQ �a];�@B�ɺU�L �ˑ7�2�a��5;'B���Y����&��`���᦯˚I��� D�2D�@.e���;R �?��)�6��	!�$�:ab�pW�6�]`Ձ�=m�!�]++��
C�Įn�<{&@ěo�!�d9=� D�&CM4)m���άg�!���@=Z���EU�A�F�t�!�$�	�Х(�!K�DOj�#�L�9�!�D�iPx͒�nթ1�	C��v�!��E�i���a�����YG�!�$KtN��V�O9#cfI��%��6�!�Č�o�:��%��78FJ\�é�!l�!���/3�	��_�T⭨�'��I !�B&k��	���2Y:�9gǞ!�D�q��Zw��'%�Z��e)V�!�D�7Q��À��'����EA�V�!�_�" ��)!JQ>S� %��F��/�!�F����U���R�kRN�!�ԛF��a勅�x?�U
��<�!�$	�J�;%���h���(X��ȓW��P�����-�*��cb�.�6��ȓp�IC��*&W\��ON�O��܄ȓ]��1�%�P#�x7bK8/6&X���R��Fġ�ihm�>4
�D{��O�mp3N2.�z�8'c|!�A	�'�HQ�6&8,ap�VCC�CfP���'��(���C� t"�h�;S�T��'Ħ�{�㉄Y|Ja{GC�Pw���'M��A䀨^/*13Ðys�eJ�'j��5�	347��;2J�5����'@"#��؈w��gJ,O,�p�'�]�S��>~���� ��XY���'���ɇl�?t$I��RJJ���'8�Ekf	�B�إCC?4o2���'݆�X�f�1��#5iC!+���
�'����n� |JI��苶�28�
�'M�*�&Ƕ�>ɑ3��0h���	��� �����_�In�����^)ON�R"O��`�N�5u�nE���J�0IZHAd"O��S�,�N<Y��C���04"O��������iӃč,%��9�"O4�ɗ��#6��K�bEY<�6�?D�D{���7 N��s�Re�Q�&�>D��*��5�I�oߝy�r���/D���D�'_�(�v�ް,�P���$,D�H��c� {�@<!��@�^�� ��>D�Th�ϖ0BZp�t��8 ����l)D�̡`i؈d�B�ײNhD��p�'D� K����@�z��H׹z%<9(5F$D�d�'.H�r�)3�U�1�i� D�0rd�1[w������M�f=D��Ge�Pr~��'�ĩGґ"ō/D��0��O/��a��-GB���� D��9#0e��c�nA�	$��/;D����L�:?� iV"8��Ex��8D�8�`N#2&�$[��I{�����4D�`��D�L)��@�C�NS��8f�8D�L�ᔂmz�l	V M�����;D��be$�����.F
d���1��;D��9v�S�+Dy`VK�!%z@�D�7�O`�.��q���P�I�$�@��Y|\)�w!w���J�cg&(�ȓ{6�<	3��`M�8K&`�,B������G��l��y2�	1u��Ȅ�mΰ�ϸv( ���+9�$��ȓb����� �%�x�x$ӤZ�f<�ȓN�� ��ͳ(^�Ю@�r��]��06"�@�.	��x�R�@��h�ȓc�f�!�*ߙi+��%�L#zP)�ȓ}+rX*��/)���H�'�d��ȓt>}����4����o�<rv���,0X���V��q�# <f����P���0n̍O����!޺9�0$�ȓ[?�LZcbT:WE|MsVF^�
5"%��9^��׃M6R7���p�h���a��q���_	D+��C��J=]����ȓb����OҊx�*dk׎=��E�_�,�|�H�9{�z�N(��x�F�N�<a��ͬ� ���ʮ>m(��Xt�<��\�>��!	 #�y�C�[�<��G�SވHkWił�쐺6��X�<I���<�=��cؾ�n3�`�S�<q*�m�~,3B�ٽ4�b�"\g�<Yd.G�G��+w�Y4
�\)H6Ϟax��GxaH;6����щ*/��u��,��y�%.m�<,ĉ��+P$�/@/�yroB"V��Ҧ��*�Z�����#�y�g4)?��Ʌ*�.)����0J��y
YTY�����8!4��g*��y�&��
�� �%7��a�F�D>�y����Up��o��{ޱ�s����>Q�Oj����Ʉ*����_dV���"OV`�%\G銌��/��Ye�B"O6�rwb�;�f8�(�S��d34"O����d�U������3c��iH�"O<lH��Xn�Q�,��-��9y'"O4<Y���9�U��_�b:����X}�<�a�B�������)Ų]�ŇƓR��0#`��Ӽ4@�@\(Q�*��'/�Ek�*e0�Yj��ˋBK����'4�Psd��<vX�G%�)@�~l���� hhSO�$��ЮM/
���"O���듅c�����ʁ�%"Oکע�<J��\*�����1Cv"Op5�6`]���C�� D�~�"O��Q�2�hI�A�e�F	 "O�`���B�d�sK�2|��y��"O��A�ʑr�q�$��	L*��"O�Xj�܀1���V=����"O�cS��%��|���&�x˧"OP,p���
�긪g�Z��~abC"O�y���e򐈠SLZ�3�:Р�"O
a�i�u���y�Ȏ���S"O>�A�_[4��S��=���T"O��;aH�h�|��eZ<��%"O��a�Nϥi� �3Q%�%D�D�)#"OD9Yq�':RAqVK�6��!`"O�e��K_ƄՓT)�*u�H�"O�s��I)�2�!J��^�(j�"O.M�R��/Q��հh�*~O,A{"O���p�@�K@�<��T�`��"O찠����6*��2���	7��)�"O� ���/��,.��E�!"O�8��ҼqN�	�r瀫:Il�1�"O���F
۶7,l�擽s70�"Ox�9�瘝' ak@f2'�)�2"Oڑ�U�%@�&�$5*4ݡ�"O y�SlӘx�N�S���P�"O�!�c�Ø9��"�l�,�|���"O<��6�m����JĨR�j�{#"Ot���[
O3�E�RDܛ-�F(Q�"O��LV+reH<H��Qخ�J�"O.	���
�`r��,VvR��"O� ��o4T�p�!ɺO��m� "OV�aUjHD��eF��$��$��"O8�"-�04��-��L�h��y��"O�k���q,`�U�H}
���"O�Հ�
��=Vj%�q		�
d~U�G"O�HБK�4�T��K�A�X@�3"O�A���˛@��e����/^��RD"O�d�����%�ebw#��Ĭ�b"Od�j%��KTذ����!H���ۄ"O@���"�@pV���S�4��|�R"O�$s�P���j�W����s "O\�:d��rȾx�1E@blLI؁"O|Bŧ��'��c�mQt�"OZM�&h�@<-2W�W�\BhiH#"Ol\�҉ƙ-��Ur��1�U�"O������x��1�c@�9Q(�\��"O��q�G�-x䐑H��<h�"O�5x�X"w��lS4�ֽj(�X�"Oh��o�%EU�I�&A�_�.lq�"Oذs��	ra�ǣ�>1v��6"O
I1�!��Y����a�� ,�4�x>��rM�P���A{�F���&.D�<B�H@M*$�D-��o}�)��.,D����=}���E�r���j�8D�̐�`Z�S�nt`C� �=dB$�QL5D���C�՞c��	0�ę�=4�y�%5D�##4G,X�h� "�mY� 4D��ʒD�R�<"��gb���/3D��pkT9/�D�2��k��9zF1D� �!eȿe�j%I��1Tku���.D�H17L�U^0�2B��0�4�㴧(D�L2#��$2��x���U�4�vB�)� �� h0@����A&�
AT���"O��Pf	ʏk.���  
0+944ɂ"OpK7*�sT�ѱq̐�.(�$��'!�ܐ��ݷPvh����<	f��U	%D�X��<��r`Y�]du���#D�\�lINz5���9��H�j"D�� �!�%�����!.$0���;D�p�E瓬/���:��X�"b���),D���lX�^��'�&#�&�:��5D��"�kɯ0&����#�8b>�Z�9<OD�$?�	n�Ȱ���S7�iC�(L,)�hC��sY��`�ʡk���0��
��B�I'4S�-�dg� T{\Z�̆8	<�B䉨t�<��f��y�1|2�C䉎p涰K���<}�A���A�C�C� t�H�����6At�p���^�C��,5gPhC�ϩ|�p5a�
.8��![E�=� 
/%d�3�Ԍ1k}�?Q
�
�N$��'ҍ[��)��A\��u��SO�`r7�	��fR�)P�0|���!�l�i�)���	��c�bą�C��膊�b(^hI4��]�ȓ(<�x�*A%�*`�HIi��y��-�QibE 
Ʃ	�
���Q�BѢ��4lZa
�#A���܅���L�T�,m����.�r��ȓk����S�385S�-:X/N��� -"�%��1e^i��%�f�* �ȓ<*( ��׎/W��(�Ɣ�2Pи�ȓ*�&0�	�s�x���G��t�8��2d.-�SW{�j�c턚WWj���f=`�@%T�[�>���VC'���Et��KB�za�H�h�4����ȓDqju�dNa�-4��\S&�ȓN�4q��
�w~�P�0퉓�l ��4�����'B�sd����ʊЄȓQ�h��B*���i�K�+T�Նȓq����U�Y�x)WNI�0.���ȓiB�X0����U��c�|�j|�ȓU�T�yp(Ҵ��l�"ɔzv��� ��신��1<�>��r�?�Z��ȓ.�,��dn�.��,y@�[.|͆ȓ�=��n��!�c��	�ȓJ�a�WY�rɁA,�S�6Y�ȓ$w������n����I�i�l�ȓ9Z�a��Iօ)\��BbfN�4����E�@��d�N.T:�}�E��$�^��ȓsv��I1��1Y��������ȓ,��m(s��.:��>��P��n��8��^,�4�rLޤb�ZB��t��9� V��x�Ɇ�n�B�2a¾YӔ��CY��ѢG$b�B�I�t� �C��W�ș�&H8=�HC�ɹ ФM�3�C+=���@�J�6��C�	�f��0v�ҏg�E�a���C�	=n �XR�똞]G�R�*N;�C�I'U�V!��CAY�D�
��L�hz�C�	 GS�LҰ�S�@���(p��0P6zC�I6F�fPB��2B��A1\$h�bC䉗�\�(�3}���E�)[�2C�ɾ�M����\��fH�)��Մ�g�x�@�[8w��E���
>f|�M��L���Q�&�)��1�-�>9'6݅ȓ/+�`�+����Hr��?� ���S�? 6m��Ç�^�H�R 	�k�Ҁ�d"O����<]q���qǈ�>�^��"O*	AԀ�4D�,Sл�����"O�]&��4����&d	�����"O�B��)H6��#��Цv�CC"O\��f���a�	����6"O�	P ע4z�𮊝)�}I"O`L;V�9{L�!�L�A0�"O�Hs Z10�� KULɏ7�ira"O�M��Ĭz���@ߴG"�p�"O"�铈ݟ��E�E[�k�@@�F"O6%bE*5R��ip
_��v�k"O�=����mw|(�(��^\���"O2��s�/t@B��?BE�1`�"O��hq�Bxu�#����~ pR"OiK�����:�e�L�F�S2"O8E�W�o(H%['�J�4oJ<��"Oz�A hG'��<#�%c��a�"O�4ˇ���*n�
�SJ�}:6"Ox5y��K9���QC�6P�	0�"O��*4$ZN"\�$ �b�	0�"OԈ���"�0��e\-Q0D�G"OD��O��T���"c]2W䶴�%"OԃK�$�\��!�>@��i/�y� ��LSB$84�����6�y"l�1�V�1�ɰ)���w�E��y�3iB<k��Ŭ)D�!ҵ((�yrς,\��y���� ��a5K���y��Ӎ9N�A FˈK<$��$	���yR��8V9��G�=�r����N��y���#QB��D�_�4�:P�-�yr  /�(��F L�3G~Xhb���y���fO�CR�^71�ʌ�$�$�y���
��Iq0��.�@ ��޵�yr �Nwl��G�)m��L�y�Z��T�7�O�(��C���yh�ȞT�غl~��A�ퟣ�y��ӱ=��@��=N8�t(UIH$�y�LG
�Zq��z��J����y2n�	o�Ŋ�����i����%�yB�ޒ98,y�kǰOݤ)"�%Ƥ�yr��v-�n߇`4\3Rm�*�y��	y�!r��^�!�ݢQ߸�yr]2}���T�Ķn4��@Q`�;�y�	O�"�����c}A�6�y��ߨsq��#�Y? d�1�M�y�)V�Dg��*�X� ���p�i�=�y���w_:8Q����u�B`�C���y2�q;����s-Xm�c���y�͖	���Jg喞:������Y�y�`�2J�.�*ƊV�,�\lI�&�y� CTTL��D��W%X:��Ά�y�披a����3�+K����գڪ�y�G-Q�x�ө�.?�\��W�y�H�	,&!єa 40�\���'��y�M�/{�0���A"8��˱���y��$w�ܸ�lP�P�N��O	��yA[誰�E�*E�P�!<�"C��-i�ȸ3�V i,Qo�"+��B�ɸ;�dp�͜��qsTF�+��B�I�g���A���0�����G�!�B�k�8	3�.Q�p���R��b�B�ɷ4����d/�EeN���&bB�	>Y�@3���B�>�'j��(B�)� rԩ����QsP���p�""O�!Y� K�c{`�U$�
�t��p"OJ$�R���Xt B ƽ�
e*f"O$Ejg�A��@9H��L(d)�4��"Oj�s�� '�F���ǁS��=@�"O,,�兊/�jI�@TTux�0"O��!th�a  0Q@�]Y]�"O"D:b$�lŦX �oR&WRD@"O0�P���z��0I�+NjH���"O.�a@h!�ܕ B�	e0`���"O�X�솤>J��W�ܠf:����"O����IW���8!p�Ϟ!-�9��"O�i�O�&
B� �'Y"����d"O.rc��!WÞ-���<1��j"OxDS��N���	GD���Z�q"O����j޿Q�$����=N�PY
�"Ot$2.Z�4��Az��;O�`AF"O`HqEoM�U�H亠�)!8T1�"O.�iJ�?�0�)sE�9 <�;�"O�`(ժˏ�T� &<� �S�"O�h�Q��	N�-U���;$�7�yrjڝ�6��Ȍl�8��l���y��a�ŋ�+��b킅��E��y��iM��*���G�DPQP��y�&ɘZ��z�L�*���ρ�y����^}[�慮W�"�H��yb�A7�*�:$k7S`$$`���#�yr!M�*:i&E�@����	-�y��P�_"�U�7��@����#��y��	N<�����5M���ŉ��y�V+Ჴb d�;/��H�BRG�<���J�G\:�cs L�t��P��^�<�B ��2�T�@+�ţ�'_2;�C�ɩ�ځz�m�
 Dy���۞.VlC�ɜyv2aH�i_4iG<mJ"��9Y�C�I�,��|q��%��R�"�8�/D��!r ӏZ�t����e2�k+D��H�E����̼*z�X$O&D��"����4���L�3G�*'%D�� �ҕN���Q�cݳ�r���>D�� D�FP!p��B1``i�>D�dI�e��.
J����%P����)D�d�T� �RJ��ア�2�����+D�,+B�@�%���T�W9^�<<��)D�`��˫x�(��dԗ��5q�()D�8X��L�_� ��EqA�dв(D�l��6M���Q�m������$D�4bB&��G���	�8��8�,$D�8H6aE�*,S�ș=�@�S�!D��b��B�kl���m��W���"G?D���5�ʞ-��MX%L� \:P���=D��S#bE�6
�� �%�� ��C�7D�4	EK�,ip�H9��Vi�pd�)D����'@:	q#��T�-q��Sw�(D���uF�-R-x�W�&��ts�'D��K�Ɏ�.tHզ�3�TI�m2T�Pq�AT�)�$��(G;C#���e"O��[���<N��ggH���̀"Oj�:����{��ग़�p�҂"O� ����T>��rař���{�"O���c�3UXn�w[*[)dEr�"OR<�C!O�3v-(4�Y7y|�)�"O0t9��M�K�NG:Q{�i"O�]Z��S�l�*�.�>�4�b"O� .����*��@ N�=K>��7"Ov�0r������^�1��"O�u[�J�G'���R�Ȧgs� �"O��3�Oѷ�~! f
T`�Es"O���s�(5���ֺ$��xr�"Ozx�բ@�HT9KU�F�D�"O����2!����/���X1"O"BC��r:}�P�Cd�|R"O���߃b��ɉ^�4�v�rs"O\�R(�"-���`նq��Q��"Ole�%��� �K��'&J�{7"Ojh�Pl�;-��%S -¯�`��"O(�@��<=��2�+�-E
u��"OX��i��"�C�̓#��H�"O`4�1���L�ʗ�[4X4@�3"O&}bj�5a p�#B�qɌ�� #!D�ȱ�Gz���I7t�4��D2D�\�G�<v,=8s�E9�
�Z1�1D�!��]�>s��Hv�e��$D� E�߷0�djLY�kڌ��e$D�@(Bh��X8�#�*����ad#D�,�a��*J]`�Hւ,Y���7�?D��S�On���c�Α]7腡�� D�lh��F���كN�=c���`"�#D���T�;W�\Q+�@fۤT���'D��@@+�'�^Y����#Dy�u;�9D�<�UCV�s�9`ү��N+�8@Ӡ,D�$ccG�'��`�SI�vК3,D��JK�#�(i�*K�~nV��@(D�hapϝ�D��µ	�+fN`��F�%D�x�`�^&v�Жj���Zk��"D�pR�h�
=|0���Y��a��=D��(�`}_�=H�'@(2 h��;D��۠?j��2b���%D�H�6ǂ	d�6��oB�Z#0U�W�%D�I5$�=>��<I3�_	ac��18D��h���)G�}���&k �5D�A�e �J��e�o��Q�� D��5�E*\��U+T�'. �)�=D���v�W�J��C`b��a�h=D��h�/
�t����)�Z���R֭<D�$��]�k�H��׍ߤ?���AE+9D�dI]rF�4��Y<d���O��!�D��Q|<���#W�bXi)VhͯH�!���&��9Y�!�Ա0˸o�!��ƄG��<����;:�E�I�T8!�k4� z���1B5��d&�o�!�!;'0�j@��5'�`Q�E�:B�!�dϯ#S���'�$>{�ݐb%2!z!��
��1H�FF�B`�,[&#� �!�ƨM����M��b�ys�S`!���i�:����#��j���!=I!�$Z-��d �w�\�����%�!�$�>S�%�C^��Ġ�!MP�K~!���S>�(��R���+"���#!�ă9!����� I�eeDY�7�!�d�j�K�g��(;���b�,�!��T�-�����_+��A	��!�$ݍ{�t��"厫aJ�Dł�9�!���&%�����_�|]l5��Lx�!�1A������S tH���N.�!�+|�hIH_�Op�hYv�n�!��ɲc��ݰ�Nވ.I�,�r!R�q!�$�n��Q�i\%�28�p#�=!�� hի4��7�x8Ã*=x"OT��e�>hتi�$Yx*�C�"O\��s�p�(���:�H(�"O��R�
�[��S��V�"O�PR�O��Lz�dh�	594$��"Or�c���,<H�E:w�۪$`a�"ONx��f��6lP`���()�|ف"O���(�;0�m1��	'<:��)"_�����<�2B-9���s����e���V�OX��O�����2:����eo_�T��2�"O��ી�I���s�X��tڦ�,\Ob|�t�T�)(�)���R"JDQ!�'ɱO�8rA�9H�����	Ϻ@�M"O�٢���o���x�h��*�<�b"O\}ؒ��l�Q��}���A"OP\��H�9.ѳ��H�C�| ��Ii�O��ed��[L\�M�@�x�	�'�8��wC��,�dE3DX�2'�Th
�'44׀A�>�(�n�A��0
�'��4��J��n�J�O�?�6�Y	�'�Z��AfZk��Xz�GL�Y����#OMA�n��ՙ���=�2�)�Z�X��I�80E��-��j�B��R����.lO��'��5"V���X��I]�V*4�
듍�����,T�A��+�L�"���|��1}J|�OT$ap �8��Ȑ�kD.X|�0Y��Iw���ɓ�~w�� ��^�x�f�h����M�����,�����!J�]مF	� ~�  �¥W����G{�x�l���[+R����s���-�X��=D���c��.�H����C���m���6F隍"G}��5�Aլ���)��:��-zE�-�p>�ܴ��dǪ\�L4���D
νȴ+�m��D�O���$� ?�ҝ������J�iX�qa|��|b��8���kP
­l��Z�o[(�y⫚�Z�=*�M	�8�r aZ-�y2�5K���xC�D��q1�
�y2�>/��	��Ɩ����ّ�yr��n��|��C&N*ƵZ"����?�" �OdU�C� �ɀ#⍍s7�9�"O.̚��N$.�b� ߪ'8A�&Z�|D{��i��!���V���CEC^4A�!�V8o��h��4��aR�a��:��d���=���ٟ- XI����c(6D�� N9T�!�d�.�%9d��!V�T�� �!���P���NآB\��E�j�axґ�$'���_�^�ha�i�<kk����j(D����'��� @��ϛ�6�����)D�l j�. P��#�m��(�R��(D���C8u�<@��eD< ����� 4���� a}*�hLW�6m  ����~�<����h#�q���[�eGt���C�S��i�0��h{*l{��{���8 �6�6"O�WN˔w��!CH�
�D�в��G���O���8�

'߮��CAؗ?�M�	�'��H� ��P� ��Fʚ+�Z	�'t}� ݼWw���ա�N���	�'j�8��U�K���˧�0`�@�'�T2� �E� ���n)C����L�R}�_��S�'~d4��\.Hq!V��!J�h�rs� "Ar�C�^C@���R�w2F���L�-���C؟̣�
X��6�e��<^��D�=LOV��$I'w�)�2�?T� <Q2�<Q�	p�'2�P�H�<.�l��c�.. l[�'�J%���j��Ӗ�O������� Xr��.C��{�bE�	��e�b�|�~zǥ~�����߭iY��'�ě /��;D�@���GEJ��&��n$#�8�	X?	���O��P1$���y��1*Z�����'�X����$�,�%��O/NY��'{$�Dy���S�w*��p�;Y��t�\��yRb�1��H�a�N��y�Sj���y2�\ 0�q5��d{�����	�8�1O�t��'i,-@��vt$�C �<?����\�$�8.\��aK@�3c���S�; x��^��$}J|�'N�dp0ۖ!���a��<rZI���HOډKtM}0�!�@X�Z� R!X�(���)�' ��9z�ƛW�Ti�	�i���z�r,:d�ЇW�0pjS7y�
����M#𧒟*�<#���,W��+4�TC�'�Q�$j��'v0�!��ҖmS����ʳ>34����D�O�#}2񏗙0�=�ē��H�1/����D#��?#<9E�Ѱe6��kL(|����Bk���'��Q� G �
�:e`D�`(Ru�dO��xr�6)뀵3$�M�t\�կ�%�0=�شj��'�P�N1`RHXE�ٰ �.W<D�4aѩQ$Bht�U��.?X��� 2LO(�(C���~�8�8Q&}��_�<Q��	!+v}{K�Is�M("�X̓�hO1�d��!���>y�3�\�⩺�"O<�A�i�f�Ң�l�0U� "O1B�m��;e$TZ �5_��T�"Ol����	�����_'q�q�"Ohx�À_�)Sɠ U�Bn"\)C"O4�;�]��0����>?���3 "O6�� &ʹ���3Ɲ�5NĈ"Olɒ5 �
���B�%�r4��JP"O��26�3\�b�.C�B$,���"O��pDO��	��Ś4��;n��Ɂ"OD�	AfO�h
�`�
���I�"O4�xA�ʔk�͚`ϗS�\��"O���J>Q������R*F��IS"O
��E�A�ay��Q�ϣd'�|d"O�ur�B���(�
5�@�1"Oܝ��n�ex�@+�bP5c<TA��"O^���ܼf�¤��A�" &�"O�\g�'D=ZQ��O�V�dH �[����ɸG�1R���< Y���g��}|>C䉳	d���
"w�
��7��C�	�<�r1 �O�_��y1�e�B�#<я��?�I��¹G��	�+�&_֕x0%3D�p���d��іǖ�B��L�X��I5�hO�>�ï�e}�U�bJ�i��()�@;�O��y�m}�]���5"GRX�cIP�y��* o���$j�m�Si ���<!���� (�r��L���sd!���^��d�e�۵V v}ӵe�ab!�D�9w^�4 �+7|!�FK��#1!򄀝#� �.��N����J
+��Ic��x�c(�)(<Txa	G.s�	P
3D�䩡�J�R4�ّ%_'K�b��@�1D�@�l��.H�C: �P`�C�9D��05ir
��� ��[���#D�k���xP*�� �M�eR�h��"D��a>{ڌ
�C
`�D�BD`!D��X�ɝ�u��$-�=�8��3D��*�*2���a�K�e��ٱi1D�03�)\02���o�%� 4S �.D�`Q�d�,���Kp��������!D�� f9���]�x�>x�"^!"MZ�Y""O�u@¯@�U	�j�lW?$��b�"OȍD��]�v����X7p�k�"O ����e���z8���"OԴu4w�z�A$A�Dl�0"v"O�������| 3F;@2=�#"O���i��_��a+q�5C�*t!��I����N4�yq��X4��Q��2y!���{�R���2^0c����!�7m�޼3f�	�:i�I�c!�$�!HW�D hH \��́g�̅L�!�DC�?/�����'.x��h�>�!�_�^��Ib�+���b��҃zz!��ՁAv�TAƆ;v��ӵ�6>�!�	��a7m"j~e��[�fT!�޲N�|QZuPF4`� ���K�!�Z��A�S  
T<H\���	u�!�Ų%�F���K�O<�e�`��8�!���L�� e�!-7Tq(v,�g�!򤍥lj�CK���08���z�!��]".צ��KZt����JY�!�Oj-�L2��3	/(�����A!�� r!,��w߾V�J'�< !�ē7�H�!T"}�"(ZE	%�!�dq+R��LS�LƐ$��Es!�ė�2Ӧ��C�����0mF�?e!�$�)�zx2�&�PQ��A�>{]!�$ߗ�T�r��\t�=c6ʑ�P*!��T9��� ߉~~�hr��2�!�d�S���(��gb�a��	^k!򄂆#��H ��V��88�E(@h!�d�.�X�� ���{¦M�eL!�D�/]�
q����9@�� G�L�n�!��^��\A�K��W�N1C�;�!��Ƃv���Ad��B�]Hu�Ѝx!��MY��6��+T9��ܐs^!���}>J�i�'n��u1��45@!�DS�|�R<1�ʆ�z��m�Q(!��4�r�ɵ�'j�4����.A!�_�8���YTD)J���a�;E'!��%�������i[�23���?�1O�J�kZ+8�V�"��XF&��F�'K����27�H;�̆�F!�$N�P�dD�d�D
��h)�D�!�d1+� Dk0*�|B�had�)�!�Dז��ʷ�X�0=�5SQ���|!�DʡTH�-�L[�n�lYы^�N`!�$1\�,l�`K;G� 1#��j�!�D^.(o�����V�#��}�&C� N!����~���6G�8��d����!���=�lJ&J��?u�h�d�K�;�!�$T�!D.]{�K�x(�9RM��!�Ï��Q��e�;gǲ��c� �!��+ai捻��ȞT�&]�ç�	
�!��(��m��G�6B� `�݅4�!���;,�F8��+����d�Y�!� �"x�u)��D�4�#��Ĺ�!�y�JI��&N+}���D�߇�!�ųjz (�,�u�٢��c!�N�\hD�B��.b�l�5�W� k!�dP	s;b��҉D�u���m߁SG!�$ټ7���Au��>���+� '!�D�0sdhz�D�B�rIy��Y#�!��ޑ4����V�Ð1��;�o�)|M!�ĕ1%k[�2T�l��V�ݠl�!�� �se��0�B� pJ�^����"OVH��)�"�X�c��_ �8}��"O�����b�f �g�0�"O�Y�'��0�s��1A��9��"O:,pEk�>b��X�4�U�.��"O���-��C��s�a�`��9�"O<m��h6.?����W�H* �%"OP����6R�$[bݦ
nʥ�r"Oh\��$��2 �nH�%G�� "O��Q1�K,h����clO�=D���"OZ� �` fI^��ЎR1orH,2r"O�@���'x�=���J�~z��ô"O�x��8>&�Y�j�Lo��"OV�X�`
����9�}!"OJ�1f�S�z�N|��
��K@iX�"O��@��Ѷ�׉S/KIX�yV"O�%��kHg�2h�h�XPҶ"O�p�䅧-�qI��H�Y�<5cu"OF��Q+O$z��`��{��P'"O�Pp�OC1���q+�,@�"O�U��BQ�JY�-XU�Ȋy��"Oj�"¼Ee ���I8\�H1 "OH�	V*
n�P����?gDT`�A"O@	�傅
�lIhp;QH�
""O����.�;�r�c���D(��"O$��	J�y��!�'e�	y$�EQ"O�	�*E�v���z����9��U"OJ�w�\�Va,�P�#�^f�5�"OxP����m���� /n��d"O���Ւ.	�C�`�0_�I�"O&��u�SS�����@�D�1�%"OJM�aR�p�\m��uaR%I5�%D�@��NԮI8�,I�N� �%D��� N<)9��9�VpI�d�<)� ʔ2@��S	ӓS��x���u�,;��N�a��e��ɝU�)�$jR�~�y��p�b]�U,ĤK3|a�Ovŉ[�#��x.�&C4
��,/Q�,٢��+g��b(�g�FjT���	d-�$B'p�U�ȓC5���$���G���;5O��!�\8t�	,K��*$�J�Q��)���F�_&8"~dr�/ܧA�,�a=D��;`
��4�1/)� ���⤟�`e�@��`y)t��]X�(�#X
�ā��+�`3�9�O�+� +a��;
5Ӱ�2R���3�.h��Џ^�tC�	aB��ᔬ�?6��dZ`"�T�.�<Y�	�gN���4L�>��O�j����шw��{���u�ԍ�'�"!ခ��o����d>d]1i,�QX}^��S��?�"�<���nΞV�*q��.�A�<A���3׮���F���EȡN}?�V�6}ش�%��<�®�"Bl�K���>]��C"OVX�@�'.R�H4�K$.��6G�*;�DͺG
�_�B�	�u���#kU���ԗ ��=Ib�ĝ��pȌ�iҗc�B�p�kf��A�#���B'!�dû'�l��f��J�Ti��i�r�Q��k��	l�>�X�M�)���h�d�y��h*�<�V⑒p����$V t��@�d]�K���13��Fq��I�Q�d�-���t&�$#����n�^���y$�D(`颅дb�CC�I�H�6xrŭ�UΥ��M��B^���.C'W�^Q@U�[�:��q�;�>lZ�m�D�I�?qbխB���M� R�"ljP�#��+�ax/��`qC�i ���ï�l�aE$�t��eJ����X&N��4B�TB��8�j�榵�'q���v��qj��֓4�$���$�U2��M �	�f\�h'	��7�@��d�-O ��E	t���P#�ȅ[N�n��m떝�$͜�(�	�@˥O���ܧj�Š����0=�"��;��R!�H�
ߠ8���V4-��I��M�~������.�hu��ʘ�	9�i]�m]Ma5k�R�$���ȏd���IN;,�THo$�OB��B!	=h��(�"?ڼ�����#dҌ��V�� &D�!�M
�OR-Bvm�<h��8��\���D�2i��q{�� �Q��-d�E�F�C�bMd:�ɟ��=��)ڐ/�=��*{^h�)�I��\ڲi���K�`CkܼQ�(�u-;Tl=��Z���$		�nӬ��"�)�	c,��"4mD�2�	󄪋�g��˓����L�(-o��;�d��>�U3�M��i�2��bfX�pI�ם�36�b*
�)v䄈����-�牬$������	*�x���9;�����)�n�@+�e���o��B��e���,�p]Ҡ�v~��)�O�b�8��g����ӬW�Z+���P��9u���`�`�U�x��DU.W�N@�ƇI�J&��7J�rĘX�����mp�̂❱{� q0g�	�9�ם������ś�%*&�C�.�B}�%��C�9��+��D�;���6`���'(�&1�%M5Y8xI��->�>�����'P�h�u�{��i>��ڭ����N<QQ�U�ʥu$��!�T9�b�ry���������H�T?�B�`ވh���5/#����%Տ>��r�a؞���>TJ͈���/���I�pɢ�)����>���#@�&d�$�O���'���H��Q&?��g@���c��^�aV`���"G0P�5�u��F�T`��X��<�U��m.�$��5]���'4bV���
�As�'	���[w]<��/�/��O�Z��@JO�>Q��	͸F��-(A�$A�p��c?����I^V��1aӢ�,J�\9��I+,��0�i����O�qr�"8uNduQ��N����W�0��ME2S.�#��>E��J<6J�*�&�/V��g/̾��D�54Y@��N=z`ayR��#�^#��ܦ|B��*۱Tp:�'�(�T�f���~B�Z�Up4��+��x(���<
߶#p��$N����I>Q��0DUGD�Ii���I�h��O@iYd�ĉ(,������<d�>āH̥E&�Jr~Jџ`�p�"4�%�@���Ї 鲉�"]_�X�2�	�y��Pê��v�5��
��<��$[�aB�h�?��)�'

�1[ %�8<Z$j�X�Ct�!��xT�Y1r�Y�����'�[ rċO>	�^Y%z��|�<y֌��Iܲ	��Y���u�v��{(<a�U�Q��i*��T�
Sry�L�,lF%�?���e�'-hF�9���,8�P�b!D�<Q��:P4|��K��R�$��!D�H���+άdO#f�v�1��-D��s��QB��h��]�ipH�5f(D� �u/�)N� I�B'e!Ftеd'D�̳�b��$�"1Q	[�X�*����0D����͑R�T��UiR�X�RL���/D��Bg�Q�
S�\*�e���:̚'�+D��{O��s�dda���39uؔц*<D�d(砏�i�Դco��;h�zV:D��Y�"L�|��L!FAX }i6��t"D�$A$@�6�D��$�8���dI%D���� �:�����Sߌ ���$D�옔�\�%o�0[�K�|��@�@A!D��ңaP�f� ��UH5[�xs>D�P����*pjx��/�l�+7?D��ҲlĽ&�H5��}�\ɸT�.D����n�,��4��EĦL����#,D��(�,^1`�h�AMI���"9D����b!���"@I��ِ�4D�4�U�&~���S��-����&D�(k��
8s-Xe�Ic�q�5�&D�h�Å7`��`E@75�Fu*1#vӺ�I�&8��>�b��J*���낹9jj$���B���U��46�A��O�|9t�P�A|�L�3LM�o] �)s"O�e��E�(�TB��f9����x�(�#�z)%��6MZ�D�Dgjam�O&��zI�$�q��'?�s��#V� Q�௛�/��@٥��e͔=z�*�O�!���H߸��C|�"^$(U.ػ��Ć>N�VΊzy��P� <�r!���c㠤���K�7��	�DJ�Vg)�Q��, 9㶼P��4O 0S�-�f��Y7G�!��"SN�Y7 G�9���S靲k�!�D�/8���Y�#/���ό-����GZ(�k^<t)�e�5=�Q>{��*^�x�K"�T�q���k 8D����0��pP�L�?�ukW�<U5��K��H�D��̢�#��r�ʓ��b�����N�~X^@�an�o)|���=�O����.� ��
� ��Vظ�f�A���vJ̯
�z�*ď?l�h��'H�T�c� b���Ň6[H����dNz�2T�U�E%�@q��^� ��\�U�~�f����	�A�r��(D����\
O0��s� ��S������<YO]+zZ�Z�N�-��	�Bӌ���{�n��~}D��ë�(�ɉ�"O*����T����0��˛`�j�ax�Z=)�ʛ�H��!&��s��OI1O��*/K�y�X��m�;h���;A�'e��s�X'Zi�A�`�e�hT�4K�8\o�Q�%��b��,F�N�az�a�0?�j�;3K�2I�D�����O�гE/-a4\��E��>�d  �O _����I&{F<�0�P�F4�B�I�[���nV�"X�#	L� _~�iF�7&S�Y��8�U z�ģ|B���/Wh}����Kx9;@C	C�<it�i��PJg���1V:0�Bl��C;���vl
$ut*�C��-�8��|�<��&Z)�T�q&�6~<1k��E(<a#-T�/&�:�[�=��A9���ur�r��¨@�u�S����=�F�q��]
G�K,(����K|8� �GI<,8��0��-�D�mZ�'߆9�$"^*vV4�8�ϑ=��B�	�c{�T0�i�pUv����j��O���U!=���F,��h�@�Y�����ĚS�2@O�hJ�"O24*�b��R���WhK�q"�(��G�##/�"M��AF�/�g~��P-bѐ��X�F��}�Pꚭ�y�)�8A>�����">
�{3�S��M+ �'0����K:w�̴��.A�	����dV4z�!�D����m�.��"�cB��!򤒋z�m+�j��D�����NJ!�D/j�PIr�ةc������p6!�4(np�q�B20U�5�w�D!��2�8�a�͎eM��!��z�!�D�8;r����(��a`B��!���-	������3�����B?b!�d˓I�`pJ�M�'�4ȒLܹ`f!�D�>=�͡���ktp������cu!�"��p����g �Pf �]�!�d��c��E����*�"��p�i�!�$�`y^��$
�s��#t�HZ�!��ȫg��ce_ݖpU�Ʈm!��hѲB#�,R�0x�3+�!�Ğ%���fHժT� ��BA�m�!��
?+h� 㪔�R6�6!H�!�$ϼA��w璅�lE0�a_�!�$Q�ir����R
H���#၅��!���|瞤( �DX7��G�+�!�¤>� ЗEW7_5.!
V�ۗT�!�$�2z��;��E���
HH�c�!�D!n&5R�'�i�g��!���r��
��G�n��y�À�!���c::���^�'�t�@��	|�!�d�/S�f����l�"�����(�!�Dz��XJ�d�8j��U��e��a�!��"'-�A��K���0V�U�*_!��)�����ŉ
.�$�3���!��K�dSB4�ӏ�w�&���b֧9!���V\�P+�)ŋRt�V��_%!�*x��5S�g�~K*%Rנh!�D��^>���:�$�� �$�!�ʔ��r��	:�B���� �!��I�e� ԑ��G�Xu�k�+�!�D���z}Zӫ��H�XA!��ҞnJ!�DO�'�5�DF�O���`@(0u\!�"[�2`�7^���a凁5&!��A�I}@�Z��*[�`<s`Ǉt&!�D�� ��p�/��]��ijd��4<�!�US�,�1�����遵�N�Mr!�� 3���&�q$�(�nCT
!�� ��1��Ύw�b��QFD5s�B���"O>Q���o�yqW�Ŀ�>l"O((�����˗OŜB��A��"OFe˒��*v�<�8,�.���g"Ot[�6Tj��e&Q�xɊP�0"O`|B���><��V5-D`��"O�p��A�2AA2����A6a��ۢ"O�� �`� O@�
D��;:�b��"Ot��,@�3kP���jZ��B"O��`��F��L  ��)~�;4"O�EꂉJ�M��&LA�!��#�"O�L�%�_wנ%����F��<"�"O��+�X!M���K��P�d���"ON]�e��4u2�q�G�ٰd��xY�"O&��׊L*C>�mA�(w��1R�"O���(݄}0�Ͳ�%M�/�v��"O0�{��T
T�$hU�.$�V�a�"O"�j�+I�8r�8Y����J�z�1�"O���e� 15����
�r"O���+\�\�(��Q2I��yz"O�8K�D�2f� q��J�D��"O���o�<���(��سB��""O��������΋�S�=K4"O^��7�}�]�E-Պ$*\�	q"O�!�3N��"4��C�J�!b�$b"O,X��#Iy��È�$mW�%CC"Od�B��Z��麴$A%J$ �c�"O��̔�M���Q�Mח/L0�P#"ODؙq&�D��D3��HM��!"Oġ��i��QG �ӅT9 *Y:2"OK������7k�X�`'��yB��8�r����D��`� ���yB��+�����ٔ
j���g��-�yRo��26~��FH�	�� b����yb�-V*8؉2+\������/�y�*��W������֭L聑 ��	�y���Evi� ��*
B�@ ���y�jɨ&�*h�C����+PGY1���H`T�� LOZI�l�\|	�c�P�9�|�;��'rT�h'J*#��� �f�f��T�h�:=v�+�`�Mh<9 �=�T�$���*�"_]�'.��	Pc׊:�@�4�	X�j��R�<>�j�z� ̕$~!�DA��HݲŢ���t�Wa��f���A�U/^&�u��+�wy���'�����¡[�F1�EHQ"�-r�'��c�ɇY�a��ǅ|�V�'<N�:@�	(82:�+��'�V�I�gdQ̤Z%C	vxHM[�$E��A����a\��(�//D��t�Y153�Q9�`��x"�[6C�,��4v��l���aZQ�$8��j��iz�Z�9 :�F!O$`����gI^979��ȓn�|���o\<+�$XT�O�3�<�L�l���s�˃GW�)����L��i]�pCD�����:D�\#G�)�n�S�Q6o�-(a���HQ$�\e��e�5(IX��a��J�R�J��H,{�괠UD �On�I�2��0{���98�\qp�����i���<��x�"�nf��s��ۮ�!A�˒��hO4��R�g�^"|��*ۃM欤	p��*ֶ���kb�<�G�	3։)��P ��\D�'e�#�X�O�"y�AQ�%TH��2������(O�X1�KK�=�nǼ2B�Xդ&Nn�8�HT�<!��WHBi�L>%>� 1��)���'/��d�������a�^� �C�	(�E�h��1��YccFE�~ވs4`��l�r��45aZh�G��8F
Q�f��N���?M�hZ��L���
:f\�2���  axrj��]Pr�!�i&A� ۤ�~�i�jp0�" ��#R��i��d���������'`���hu:� �Dʹv���r� ;8\|S�f��zy剁A��H��՛ ����\�1J� `�N�X�!@o(��� ��)�*W�-�墧��OPv���O�xa�>��i�
ӓ\� �ˆ1�f����#���᥉�x(+-_����\�V��1۟N������~�؂D�F��8A��2pzP� �h���֒E��!���w���c�V(� ���a��w�l� �nκ=�v�����*i\�!��V�u��˫OTAې��R��=	)��e� Y�v��@&�L����$>M��z�����HSMӼfE�]b���"G� �s����F6PI�-]85�

 �tҴ=ADS��QV�"U
��)�	�=�	@)۔M�l� U� �8&˓mV8)�����X��υk
H�E0&N=I���F]���lB:�[�F����j�N�6�^��>7�t�[)t�&���(������WI(�0+��у9�؄n�>V��c	e�0瓘T \U��O*�<S�@��;�ޘb�J�e�$���J1�"2o��4d���Č3�tU0c!@/��	�C�^�(�y�GȆ7L�RL02 ��U�y������A��L���M?)�~�C�����Q@���5����!����'tM:��Y���M�@
R�0<]P�D�"UA��S0Nݕ��i>�r��t�d M<��LX*����xȜ��&FyB#�9g��p�F[�T?)0S.F�1��!4�:4q�@C�d�X�F�B�����D,)�	�j�"L��	�I��1�Ѵ^6$��#����!�L�@ЇA�4j	$�'?A�ǁ����dn�'lJ���cE���q�A5y��\[R�\��eg�!���P�ҐuR[�, E(Q*b�	40�'A�D�\w�P�������O+�]����d 	�鑍Q�Z)R��ңzL�q 䈧�ħg�f��f��>��Hc�&@�E{v/V�o����c�52��)��L�WbҢX���#�XH�0B�ʵ<��6ea8��H9}��)�*o � '�R׋��S�`�ѫOʁ��C�1��B�'��ȪP� �dSv��M����I.}�L�2�x�kg���'�ܥ����az�;1���Ӟ�"u��0�����'���з��.�QY�%�$~3r��baԻI�@M����U�	T4���L+�'i���`!�B��&�E��F҇�LF~ �X�S ZS����?5�P\q5�ժ�^C�I��x��R� ����D x�˓Kc���!�ӧ(�p%P�ɑ/e�v�T��-@H�p"O0��rJڃp4��2�&�$�f&#���&
�.�0F��dA��`D!Tk��p���
x��q��;U����Sg�oԄU@�,��x2%�	h���jS�H$[K�%�b���y���/"��eːQ+�
3%Ɍ�y2 �/t�̻�AQJ��8@4M
)�y� 3�,�l��Fa�0XNX	�'�<!k�C��!�5�I  ��]��'2��ǀK�V��{&��7$���	�'(8y��E3 ��a�`[	
�u
�'���+3V�����&0tb�y �']:Đ!��=~��I@��k�� 
�'��z�������b 
pl��':�@*LZ@is���
�n��'���[�n�,LV|\QdE�vȸ��'�:@��bԭy���s�ƤXY( �'z����*�<d�&��C�Q+dP<P
�'�~X#�׌U�:��FF� e���	�'E0�sN�h���S�L�a�'dv�Itn�v��P����2�%
�'�H�xA��\�	�q%Bq�	�'�T=�s�]�e�<�a�(1��-�'�4�e��R>��M�-�|Z�'S�F��b��h�F&_A�� �'iF]r��{�"��UM^�'��<��'u�8Xs ��cP�͹�hޞ��)��'���{�� =W�L���&E% fV[�'����ƿ?6� �M��.̉�'g��[� �)}���8�:4P���'�r��\,��V��~xj���4�y�&��;p@i�C&.G��}�Q��y��M�s�j��<�����޾�y�/��jlxZ�T�,�`o�y��?f�]��!q�
	��V��y���4N`��B�.Z�rB,��܄�y
� PtH��ӈEZ:��l t�J*O��B�ټ.����Y������'�]R�h�I��	�������'��(��E[D�n���cV��T��'C��q��59bJh93��VIn���'rep��(��A%KI����Qb\���>��:=�6�k���P��ȩT�[I�<��i�5B�Vk4g
��"���/�E�kv�c#a'���v���8.<���H�)S�	8E"O 8� �s��j'�;(M����@�gb}p �>	@?�gy�H�I�FI���)~Z��k��y��ńW�2ų�,�X����M;c�X\H�n�>ƾ���uf`ɡC�)�����ƴ�뉻g<	�DcD:3/��(��Hw捋"�tLi#"4"!򄊆5���8�d۟kˎEѵ����qO����C�	K^:���iT�
��s�XG�vY���E�w�!�$Ѽll��b� 8A����*���F��"�U�T�|�'sn��T%�h'T(2UA�b�옣�'"�  �N}�#�Vd�,��aZXJ�!Ԇ�0>iw���_1���ɑ1mT�Y�G\��xb4��sQ>�7O�rg��R��a���p0n��"O�e�u* ����a��@����C���=����%6�bF
�+��ɻ�n�K3J��@�ȓJ|x0�D�͠��ț��t�B)��ǇHEqO�}���&�9�F�$S$��5��7��ȓ4�ެTI����cf"Q��}��&�L��տ^�9�BAO�mB&�ȓo�H8J��@?v2�r@FCx�PԇȓsHȍ	��0%��A��,�v�B)��t̠�E���~���M_0Xl�����8Ӏ�/-Z>�*�bW�⨇��0-8&n��V�0,�l�R�Q�ȓ.UB�(Y�O(��A)�Y�ȓE��y ���%H�\�*T��p��ȓ;�1���@>@v�B���Z<�ȓ�� ���S�|�b���69������F�.j��0*��(T:���P�0��"6���9���u�hM��i���t)�����Ղժ3!�4���2�*��
�H�yBB@� /�|��;K�ɪ���}�\�@!`����0~����L�A�l[�m�%s|��ȓlWb�S�A\�t�kFNݕ	����s��} �f6�[%/�	���ȓ�n�x KڢE�As7��uL���!�H���-z<~p4�ZѤd�ȓF��t��lǇ����<y:p)��2�l��U$Y�yzT���{8�H��1}(��y�f�����VY�Q�<�	 �QV�mh#gS�z�n,�w�{̓l�H��Ө�t�LH�s.ҳ �D��ȓa{�:��ǟC�H��(�65&���/o��в�ӂ�A�3E5�6ń�NaTt�T�udX9"5��H�R�<�v��<Oڮ��`��(�8���C�<�,[�
P�l��"º.�v����x�<��$�cܪ\����6%}F����L�=mK�"<�'��	�T2R�2q��7kפ��^h�@T.�>����5k���I"rq����B�ɟ��$�L��<)LԬGM���W��2Ph@�d㓌B��I��)�&_�S�O+�jS�K;wn]����;�\D*�O�زD�)§r/�����56H���pc��I�dH�P��<E���\M��;�/dw�Y�1�ʛ{*M��ө_k�l����d̂1ؕLE�b&֣<!vB=�b� 6�RU^�2�j'��Ѡ�$��(O�Op�<���Q��h�d��~3�xH>�y��3� ZE!��*o�i�FT�p4p" ��>I�O�Y�S�dl�(6�6mC�aXA)��X@@M��"��`y�hTaA&
M�ĂM���6��L�����|j7) m�N<�� c&Z0��LR}b���o�;��4g됢�@B�		��) ���O�� �͔�%������1���t`��<�	�'(�QQ�..'n,�e@LW�d��@�r��b�f���de
v>M��隍�U���7ETtL��䏱WҼp�v���,��C�$~���'�H��t("c43�2�����	Z��rZ���0.�#�qOQ>řB��06J����8� ����OL�s���ڸ���"0�.��Z
�xIF)�\J�(&B�?ᰝ�=��'E�ɳ'�0E����iCt�Y4��4!���?�'�NA�`G(B~<e�V��a�&�	�'�<\�@��'|̠$H�ٗ`Q x	�'�N\i�+�4�&�����R�� ��'��D�߻�<����{�=Z�'�X�14��.4�<YR�N0+r�A��'�h���L�.I��A���D�'�R���'k8р�G�/�8)����A[�'m��G*��R@�!��J-{�'�!�b�כg�h���ƋS�H�	�'�[ H��5�9y��	4&�|z	�'�P����#�\����
&�֥K	�'r>�J��N�:���A ���h�	�';j�@!,D&���:AoG�Z����'N���pi��4���O��U���'��h���Mf4�⤭�8bT�S�'�~䉳��1n.n��$�`�.-j�'�x�c?$��@�ӈ�,U�t(c�'t���8n�Na�#�P�EO���
�'%(�;�H8�����
b���
�'����ɱ#�cw�݌X:Q8
�'�ܵÑ`�#g�4yuC��s�q�
�'�P���<X��9�D
��<�	�'�����N�"�b���@ ���(�'S�X§0R�9(�k	 k�i��'[((�2�kn������W,����'邼�7A��@c𕰥�Q�DXָR�'�Ab�M4�L�z�8g28�
�'V��� O5' h����X,4�@�2�'�xU����5#2HJ�㌈Zj��'��i�F�Vږ�JW"2�8%P�'�@��ǃ9W��ɶ��h��|�
�'z�M�dH@�}=�x�%ُY����	�'������=����e�T��D 	�'hyk�NY�hlT�!�D�IJ���'��	��J�)� 8˲	�{�$�'�>0vL� Q�H�Bu�
�zf:p �'"�0��\���h�$pJ�Y�'������T1��;���7V�i��'����+�n����͌��y��'v$���T�����~`�E
�'9>L�P�.z�E�����BDٺ�yB��|μA�嬜�� ��,F�yb�%-2���aE֣N�;�H��yD�n4~����?9:ԫ���y�-��{��4�
m��-��y�㐡16ʁ�æ0�U�����yr�-@����z����(F��yRř�B{�r#��&L\d�V�3�yB�ޝ)A���u��-�QxsI*�y�B���ҹ� I�\�<%c�!D��y�j�8@���a���\��A`dĽ�y��T�	t��{�ЄUy���Ǥ8�y�%,O�����I��L�7��'�y�N�8�B�"U���8H� ��V"�y
� xh�g�Xi����Pc���"O
�d	5E[ e�ý!O2P��"Olٰ��Y}ŋ��L�,���"O��spI�c�(��fD��
�(�8B"O�`�����N3NECp�ō1�
,��"O�i�uO��]zJC'��"]d=�"O8�8�œ���I��C b�ʝ�!"O(5��+> I�b[�
�*�p�"O����H�-s�mT�Hs���"OD���ʟ"A@ٔ��i,�z"O�A���0���'2\�Dإ"O�M�P(S���C�W�?�>��"O��� ��c��y$�<@v� [�"OqW�5^͢����QZj!��"OJ�ȳb�?�x�BB0{E�"O
�I%���.����5X�8�"O���C.H��Z��1 ޚw��1��"O$�(%���C���)��d���
3"O�,�s& +����9U�ܖ(�y҅ҏk%�D�dNI�SSJ��0�ȱ�y"l�2	mڄ�V_d �� �y��I+��b���h@�wD��y��^	@p��ғ� ���7�y(�@�R�"Ӣ!vp@��fJ��y�$ђ'�4�c �WŤXzk�y"L�G0���)�:��i�����y�NԤ7�{�i��d����0�՝�yB��:zX�xA��Zהa�P�$�yr�܆��)q��JY{�I��m
��y�D!2�̤��N=z`C֯K��yr�Z��y鐉9[��kUEM$�ybI�[�����;4*.�E��0�y�#�hy��s׀U���`� -�y2B�83���P"k�J��$z��A��y��'	�lې���@�l�����y�lх&��S�̅�2�ڤa��y��(X��[Y�����O�m��s׆(��̘(`��q'�SX���ȓ8�԰���f���n4�8p�ȓA�
H�enk[�(�eoO�[�乆��d��P �=Rݸ�g)V  en���x�U�"��	#�q�*=b� �ȓ�D�`�(ٌk��X1NB;d�ņ�Wb��E/��?�n!B�*I5�$!��H�r�%U!�:��α�Pu�ȓ1�H괉S�v&�,��	*-JY�ȓ1-X5IF�ې�pJl��k V�<q �Cu�r�:f��+O����S�<��,I#�r'��*SP\��PP�<QVLS�B�D����Nؠ����r�<q��ߜ*&��R��
�'z\y�/g�<!��۵�4 2��n4�Bq��h�<�RUX'ܽ30i�VO��ҡ{�<����*DZ��3�&�6���C'�\�<IQ�ܕn1* hfL�cَ����r�<��ܕjXTQU�ۃx&t�jŀ^Y�<���j���*Z�(�2h^�<���-�:�:��Q=jt�RR�[�<i�FՃ%�X�tn�?YD��b�AM�<�À�9wc�j"�B�.,N�:���E�<i MP�'��t�ufK+GX쐂,�A�<�tEҡ �4$��l�}l\���G�<V�߻��]�CBN�V�%ip��@�<9D#�9M'�q��'}`��7 �z�<� H C%�W3?rF���Q�l|#f"Ot��H�4z�
�ɐ��42pf���"O>4�%�ȅk��4Qt	D*��D�"O����^��!*� �3L�%+s"O\��*��)��Q*qIQ<q"O0�Ѐ�g`�Z���YKn��S"Oz���
.cв��@�C$/�=P�"O�qBuI�<&�N�)���o��\�p"O
�F � �Db׉�&�����"Oʜ�QC�#P���V.K5b�l@��"Oĵ��EC�E���΅,1p&�"O�e�v��.s
��rPǀ,"Tj�Q5"O5�C^� ��q34��2io�չ�"O��D �/��i'���M{���@*Oƭ�-�*�&a
W�!<��k�'�8e0�(ձB� ��f��	���'�yae�[�1X��T�X�4��')"%IT�Y��;SK�C�'���q�B�0I<�bsF	1}��+�'�>�Ɇ�A'/���P �кv�R��'�&��bMe:iÚhxq�	�'o�9Ҳ+L;$)6����޷b&�%�	�'���Ä�L�:+�x���ĕ`���"�'�t���c��k���UZ�n8��'�8����B�uI�|	 iU)&�\���'B�Dcg�4%z3R��qT|��'*]�Ao��8�����h�3K��h��'�̉����YC���B��DLRE �'��`h1��7��x"A�̊C&�s�'�� y�
[+C&�������U��'��I�AeɭH���J���
�T��'����������烽�p��yz���C7:R��@��ɀ����T|���t�a#B^�PM¦�}�<I"%[%G�:5jԋ��}���jM�<��$�	>^��8�D�K�b��3��K�<��+E��� t��&pJiyB��~�<9�Ꮢ=�� ���# �|���͟N�<Q$"IH�	�J�1�D�#��@�<��(\�'��Q�"О9Ĭ�r`Fs�<9�J`�����d�ht@'Fs�<aU$P �v��s/�H� �ekf�<�K��1S��s�Ǝq��Y��Mj�<����s���r��%^>𰙇��h�<���:�&�0�	 w��q	&E�d�<�Í�fq�]�� �V�Z,�3�G�<ar���&����������!��7�yRd��d��%��5`��y�G��p�`P9V�S�<�����y2��L
)�fJF�FZ�L��Q��y�{�\�T�R�@(���%�Y��y�k�,P���bI�g	2d�-��y�$Xk]$� �܅XA���U�J��y�S��mB�+L�M:屵���y"��u���a�E�	G�����Ґ�y��ۦ
;�P��N� #K��y�Ʉ*<�f�"A/\)CV�]��y�թh]%�"|�V��ugP �yr�t���'��u��PiԷ�y�n�4x���i�
~S�ukd)@>�yr�ԗe.��oޥs��٘���yBM̭����N��8t�#6	O��y2��� C��2.t$������yr�W� ��"�dA%����@��y
� ��fi�N�N��r�<d�a�B"O��r���'���E��VN "O��#�X�Y�`�!E�?YM`"�"OR�z��]�2
T{U#92,ؐ�"O|0�aJ"\�^ )���"w��"O��; �(@�Ax�A�"��tr�"O���ȅ�"R2nYJ"O�%�@Fޔ[�x�����l�,t��"OXt�"Ƃ�F��Cw��G��w"O&��PK� A^0I�A�)^x��"O�=9�-�	���v��{	F�S�"O�T�0f��D�d��O�"^&<r�"O<��/@7�P��5�;�݃"O��G]W�����.9M��M"�"Ol���   ��     K  �    �*  �5  _A  OM  �X  2d  Bo  
{  �  ��  �  �  ��  0�  F�  ��  ��  �  [�  ��  �  ��  
�  ��    x � [ �   U& q- >4 �: YC �L XS X[ �c 	k Uq �w �} d~  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR��D�J���ӳ] �K��F/]$	����kϊB��.p2:d�a�,��������=QÓh�D}*���\�<�{ĥ��1	bq�� U&�2�A˼m2��v��$&����
rdk�A�)!��T��ΣT�8��re�q���W4O ��Z���+�'�δ+Rh��Zc�,��D ��2�S��f��zA�QW1�ɢ�݈�yB�S��n�A��M)3|��
I�v6�=E��ULD�S��"�l�B�C�tgZH�ȓp�(8�6̎��.��7�(1�І�_�%�l�-�w�K����ȓ{��4���`��n+h,�ȓd�Y9`X�^�zQ0QN�GU�ȓP~�����+���
u����5)�ذ���
T
���A�N+���F���c�H�h�>�Io:[�M�ȓ���G���,�+�T�g�0��ȓvU�M	���}0�P;�/a�f��ȓi����P�C*r���� T/jt��ȓ7��0�R�#!�X\�4�c*)�ȓ#���H��&l��:�"?r�����na��جT�0��j3R��܇�Z�ڜ�B ��w7��1��X2���ȓY���K�K<�fX�&�VL	�ȓe˜,�ӨN�Tu2tX��ĭ[NrP�ȓ�x�1m�(H��dϰ:�����4x�M*O�����,�\��>�8� 'ְ%?�8�3��t�$(�ȓy_��Q`&��fut�@d@Ϊ>�-��qXXգ�
�?Q�����'����Q�հ <A\ ��j��#o�0��Z����-�;�`��q��-/ y��g�&]6HK�Q �/I�����"D����@�,c�vh��F�<��"�g3D����l�Z3���^2CG0D���Р� 'Ava���ƴ�V�1��/D��A��� &C�5��gļTzJ�7l-D���rF�+%�(:��_�Tl��7D�`)���6 e��@����B����+D���a"ϑ"���b�C[t�$��s�*D�pڳ�& �*��e�لF]y�U�&D�d1�-q���/�rߖ �&D����oH�B����w��JAn`�.(D��:�`
q~��Kq�^>2\��!T�XCe]��H�Z�@5h���2"O�M��4l�d�
׃��8�ndñ"O�1b�b4��-	c�σc�4��"OH�y���ov�y���D�s�jU�"O0<"�*��0@p��-b�
��"O>`��7`��ܱ� ˅8:3"O��S��=ǰ�Y%-��N���"O� &��'��=y�~���L����2@"OT�	���Q'�Q0JI)RXIw"O��KD�5�F��(N;( R"O��#R��39���(ٯi�4A�"Or�PVꜴ-c��e�؞
�����'B�'}B�'��'o�'���'
&p�k��8�5i��3O�AP3�'�R�'U��'�"�'.��'E��'�Ќ
a��R�`A!�D�K�^���')��'�"�'���'�r�'���''�y3���o��@3����3��'��'�b�'�"�'�b�'�b�'Bh�CQ�S��)en���K�'A��'+R�'�B�'�b�'���'ONI�GXt�"�J%Cۓ�8���'o�')��'D��'�B�'���'aV [c�]�DJ�)�����bD�'���'�R�'���'2��'���'��$��D��ߠ��4*Ol!6�'Q"�'�B�'�B�'�R�'���'_�	��e�,y5���U������'���'�"�'*"�'�2�'r�'������ė/*��;�)��c�u���'r�'���'\�'<��'�'�3P�)-X(�q�fA�����'��'�B�'���'n��'��'Ԕ9y�HG�<�����dݷ6�bLH��'��'WR�'2�'���'�2�'�F���+��: 4��e�e�~ ���'���'$"�'[B�'�NvӮ���O��	U�wY����^�!�Ȭ��xyB�'h�)�3?�i^�ik��M-gYV���#M�+g�����"����ڦ��?��<q�zXU�C��W>�B�b�7A�����?yt`E��Mk�O��S��J?�7�7eD�G���^�,ٕ�-��ş(�'��>-�C���
�o؄p�!u��M;�A���O$L7=�28�jS�	Y�lN1fXp��r#�O��D{�ק�O���ºiE�����\#�Q�I>)�PdN x&�$m����E�=�'�? 
�(��e$(���׎��<!(O��O�@mZ�?�"c��9��]�bKB陁*$��`��X���I���I�<�O�`e���̞���Q��٩2&�,��O��K�rf@Q���?Y�b�OTx��ꖂ��#���(:�|�q�a�<Q*O~��s�,�wfP�<\��o Ԁ!R�c��ڴ�b��'��7�&�i>9��ƚ�L>j$���S�����l���I�d��!\�`oi~R5�da�Sk���P#C
5i�E���&n��ꢘ|�U��ʟ��	Пh���|��� =!nJP�VkW� t�ەIAyrA�O.���'��'V��y��;���x�`H�IW��+����_I��DX�v�x�*�$���?��SgT8��	�^u�#C`�H�IS.�����542���7�2	��f'�'!��0�ڵ��$N0KWxAx`JVU6����?I��?���|j,O�n�<vHR��I,
�<��*̫4��+0ρ�C,,��	�MC�2�>�#�iN 7M�Ŧ�+@LAzGX�5N�i@�����+F�l��<!m��u��8g ������z���������"d�4�Y�E�0�%� ��<I���?���?i���?����,߬��dJ �L{k�p�4F[�5���'���f��1�6�t�d٦�$�({%��,OE�����&O�8�3
2�䓈?���|�E+���M��O��]wx�b!N)˦�����=�F� �G�O�t�*O��n�iy�OC�'���(M)�]�2(��J�&q ���"�'�剂�M��e~	�I�$��P���O;d�&�b�̡���.6����Y}
l��m�"���|b�'f�j�q۝��,�$�^R��|ɗ�.ъ`��ML~~�}�y��'h�i�'�wH�z�(�W#E�	�h�Iրt���'��'���tR��ݴ!�H���"e���C�
KI����i��?Y���F�'�'oh��?��o�g�����Aպ'x��""<�?A��i;z��D�iC�c>}��f͆�����j稄�I�|��e ��^@:P�)�M#*O��$�Op���Ol���O˧n��ӐgF�fC�
'K�'���ĵiʂ����'�"�'��O�ҡr��2�{%,J���c��0�� Cv�'P�fi;���(�D}��;OzaׇG ��ٸ7K��I�A�P2Ov 0R���?��Ĺ<��i��i>�I�iH��x�M�QyP!�r��>�*��	��D�I���'G:6-��f�$�O���ƣw��t��)=N� CӉ4h�,+�O�qm�M+��x��
�\�x�h˞]�l�M����іͫA�����I"�u�I̟����'���$Bڭ9\���G���].����'<r�'R�'	�>�]�d�p�����?ZZ\z��U�s���I������*���OL,oO�Ӽ#SG\�B�`���8qx8Y�R�<)���?��i�x���i���=�,1C�O��ףJ@5�����^�1㐅Py��oӲ��|*��?)���?��#���d�[=��P[�-A�it\��*Or o�2Z�E��֟\��_��֟�#�ڋx��R��)'�.�@E�[/���O���j�i>=�	�?"�O��>DaG��mdQ+ԧ\82�����-?�F�E�{e���^���Z�՗'�H��W�V��4�3�K�dY��S��',R�'�B���S��c�46�F����-@"mx1�+k6�����8I�D���8ћ6�d�ty��'���ehӒ	D��.-�`�ǣ�F�[F�Y*)�7�r���ɥw�(ut�O%��H����� �!��a<{�4��DL������7O����O����O��d�O��?�r#�T����憭V/��ٟ��	���ߴ7~��O�67�>��S�*��𢁓b��,9ԏU��2�O�4m��M�'�
�`ٴ�y���n��$Z�BT�r�L�R�^�A�|�7�X&H�)�u�O:��'�r�'�r�'̜u�c��2k�\�sgϝlE�U���'Q�T��ܴZr���?����i �W���z�l��̕Cv��;6�	����O��D,��?I�g Y�VQP�	!$ �q�LТ"EX�{`���4�֦���ĀSA?	O>	`k�	2���̰,�����)�?I��?	���?�|Z+O��o#��|� W#l�j�)\���a�GmN������MӎҪ�>���nm��*3M�~�x��*�m����?q����M��O�LS����zI?I�ê�(.��82� M|�5��k���'�'���'%��'�S��4��2(МE�`�f��'ވY۴M+z���
ش�?9H~ΓM��w44ѵF��]n��w��*n}|����'+Җ|���e��EY�4Or%�F��5d��wm��0,��1O�p:S#�.�~�|�[�@���kFD�QlΉ�!��EӠY/�۟��I��8�IPyB*~ӒaBG�O����O�P���.�(0��'���xrO1�������O��d%������Đ&��#Qꩩ�(_�V��I�(�``����+K~��`�������l�GM^#St�+6bϡe��9�I������IT��yg�W	t�� �	Q84Ś�Ķ[���f�zH�5#�O�������?�;�����üT�x�ʳ���p�r��Nӛ��s�b�oڄFz^�l��<I�:���������'ϫ~"����*'����t�K�����4���D�O����O��W�)�fŊg�r$�B�!&˓Yb�*�P�'�����'�riS���5>��i�dh�
F���h�>���?�H>ͧ�?�����	j��q�pi�:�֘;��A
@�X�'v"�0����R�|2]�H������L�{�RR�܅�@��������I���@y2�~�R�:��O�)c��Ĉ/YB�@�c�&l���O��l���$���O��d�O����,Pg~4;�� ��
œ�v�Y1G�?��3O����B+�*��L���?i���a�5N�6/Bif�!�H����|����x�I퟈�IO���D���8Yk�E*ƍU1b���?��G��f�X���$\ڦ&�� &�Ns����mO
D�&����I�I����i>E���Xʦ%�'.���K�CM\萗���4���O�X�������4� �d�O�$�`�4\�@2*d�2g%�O��d�O,�u������_O������O�rH@��b�Vy�Ř�'���j�Oĥ�'HR�'�ɧ���'���au
51���(��m�e��ϝVȌ}���i�rʓ�.�:�	\�	��`��=]zPY����"��I�L�	���)�S}y�moӮ+D�-z��tCݡ8^�h�2�хp@�	��M��2�>y��#�dls�l�,O
.�h7�Ԗv��(9���?9v	��MK�O� +%�ׂ��O:�ٚ�G�
�b��b�'����'~��˟�Iڟl���(�	l�4jͦ�����*ʹ^�����̑%�r6-&*U�����T��y�ǜ4�$�˧����:�s��&�b�'Qɧ�D�'b�䊥.$�f4O|�C�I��c���m��#�2O6�JJ8�~�|U����Q
�=�ʙ�s�EX���9���������4��Xy�e�&�����O��D�O!�Sd����q�c�SJD��0�����d¦���4J�'m���1 ?:p�� J\+�>�ڟ'J� G	,���������Hh�V����ҷ2 �E��lT�KNMXBИ'tF���O,�d�On�D1�'�?q�(ю��Qc3��"� ���]�?�ÿi�6|�g�'�ңq����1*%>h (��S��U��^�u��.�M�P�il�7MS.9/�7�m�8�	q��z��O1>�3��ѿ�ֱjp�D�)C��}�Ey�O�r�'#�'���̆-�*�I�gW���a��cД@�	��M+����?��?�K~
�	8 j-[Y֨[DRsO&u��P���ڴuB��)�4������X��t($�"X"@�Zv���(�a�R���c�Kt[��D�IQyR΋�\�p v�ͶIߪ���m�s���'�'��O�剨�MCBω��?�m�>l&�P!C�V�+�D� 4�Z��?D�ib�O���'7B�'~��Ob����C�x�@h=1���0%�i��ɡ-�� �ҟ䒟��/YV��1���9#�� ��6��d�O��$�O[l�ܟ<�	}���0Lbfd�>`8h6�ņo\fLB���?Y��C��6�����'�t6�1���X��X�V���1�]� A�F|ܹ%�`�ش��F�Oa��{�i}�D�OƱQ��9�CLׁ<�}�oD�X�,(;��'�t$�<����'��'r2�iW�ٜ�T0�GUc8���'{"R����4w�v�����?�����IU2v=|�Sbn\�����¸d��	���Z���Y�4����)J�����!+�˂��|T���5�JT��h �j�3��i>�0�'l��%� AF�����U�����.]ܟ���ПH���b>��'47-ц:z�b�N�(t���˅�r٪1���x�ߴ��'��듪?��ic}Dr�����^	�� ����?�e�ܗ�M��O��!֣B<��π �Y0�@_9B�&`7�&F����R1O���?���?A���?A����I=F-p[Ч��@���t-��o��n6Y5����ן��	S�Sן������e��#�6����@?)8�U����%�?������|
��?�6I�5�M+�'W�X��$ɒ;����"Ot��j�'K�����Xi?�I>�(Ox�D�O����-HrIn���(�g�O��d�O\���<d�i�x�	��'b"�'k: �`RM�9Q�A��9���'�'��듵?	���$.4��"�al�颥n
�6����?��旮f��-�ڴ$C�I�?#4�O���u��9a!�����]+׎��2@����O����O��;�'�?����jh	Q�ʪP-�YC '�?���i2�QU�')��s�.��]�W_h���+�-�}��=9��	ʟ��	ǟ@�!��٦�uwW�9�ɐ-�h�%`��mrr!a%!�|���Oz��?���?a��?��P|�!�0��P���`�ת��",O�l� �T=�I�P�IE�s�P�rN�8+�!��-�*=�*U�߁���OV��"��ɔ�7�(1t�4h>�vfI�*��]�U�n��0�'H��D��m?)N>.O԰[K��[D��R�PMrY�L�OH���O��D�O�	�<�t�iJd�@��'l,u#b�TB������,@p���'7-(�ɗ����O����O8��X9ci�-p�/�J��� ��/{�7mc�x�	>U}�!xڟ>˓���W���X�,�e�bYx���>��?!��?y��?)���O����/�\GZ�	Wl��b}�=��P�8�ɡ�MK�*N�|��
��f�|�4��\�Rm�k��i%��3]+�'�"�����38�F���4	�4�R+K�kYR��E��+!��H%��c?�H>1(O"���OT���Oܐ��`�:�0F��$k�C�����O�˓<��o�0<r�'d�S>���L7O��YY'�Բ4�H:2�:?)�^�H����|'���CD���$�r*�!�V�bo�=D���Y����Mr.O����"�~r�|�/�$*�`eH���
޸�@/2&�2�'�B�'����T����4qsz�a�#M8����M�Nb�(�`���D��Q�?�\���I ����4��*gr���	֟�q������Γ����4�	�<q�g*6�hD�	8! kW��<A+Oz���Of�D�OD���O�˧%_�M���ʀf�x�M�/K�d@аi挤��'1��'M��yR|���#
L޸�ъˢM�b�_� h.���O��O1��(�+x�4扁o��")��m�a�F V-OA��*�"�҆�O��OJ˓�?i��sH�+ѡ�B��ʅ��<��� ��?1��?Y+O�<m��(�h�Iڟ��'lHI!E�'42��h�c��n0�?Y�P�H�	ǟ�$�����T\�ą���+��M�Մ&?3C��3r�s�4��Od���?�D�5����+H�H�pM�,,��d�OP�$�O��2ڧ�?��P�|�@���G�}��`���׊�?�]8��������4���ygo�:XRQc�v�kWL� �yR�'���'�S��i���O9���,�����	-�}"u��r��C��(	��'��i>�������џ�I���`�&IT�]���J�|�ĕ'ـ7��"bU���O��3��1Z>�b�K�O�N�ѷiӊ��P��O�xn��M1�x�Of���ON���̘V�(�Fi��6Lv���\;,Τ��O���o�9�?�0�İ<�A��bA�G�2ʚ-��F�?9��?����?ͧ��d�]�w��͟ p$0q�e!�By*fM������4�?�J>�V�d�ߴ	��&�yӸ|��� �e�B�H�#���:u.�MӚ'V���E���8��dퟲ�.�5G��|x�oR���(���'X��'1��'�2�'�����Ӭ,*(\ahN�r�0��c�O<���OjLm�<�b�#՛�|�L�4҈;j�8=��Cw�ѩa��O�Yo�-�M�'�vLߴ��$��i��5
�<6�Ph0v� "o�uP���?1�/%��<ͧ�?���?Q�7?T�K�&�;��0%ꗧ�?I��������b��Jy��'���?#=�U���6v��v��&,t2�9n��֟��IT�)� K�3z��a�����"<�m:c��
��<S��*\�l����-�ȟ��A�|���M�T��ERĽ���24L�'#��'���T�d(޴h5�	r�T�%&bh�U��7V	��K0n�`~2�p�T��*�OR�䝖
� M�b*T�ʤ����8��O��Gi�P��ӟ`�D��T���<��G�YE2@��oXi��(�1��<�-O��$�O��D�O,���O4ʧi��cmC7Y�r���OV�|��i⵳i� ��'��'���y�Jr��Q�F|z��lS.<
Y�K�m�����O �O���O��DZc��7�{����%�+*_�,��`�$x�����%g������[��,��<ͧ�?Q�gW7F�~�R�C���LR� ��?���?�����$���	Bg�e���۟���e�A��E`���q��a��s?��ܟ���E�x�D�bM
�RGFxVa�4�ŗ��)b����\nZq�'[6���ş�2T��[�tиC��6'���[�@U埴��H�����G���'K~<k�M�J�VU���O5p?*�t�'��7��]^���O0�l�g�Ӽ۳�m�tP�I_�@���*��E�<���iT:7W��! cn^Ϧ���?a�-�*~H��B�? �H�"b�7q�敊�+ �1��*���<ͧ�?���?9���?�U(�zr*�Å���۶��K��d�Ʀ�@�wy��'��O����58��@�r��i�E+�33L�
]�v��x�$���?�Ӿ���B.l��-�ǣػ8=�O� =��u3Bq�tG�OR��M>�,O�ȉ�ڻ���Q�k,:��i"�"�OZ���OJ�d�O�I�<1'�iӤ,K�7� V`�s��X���@��KC�'Z�6�;�I���D��A��4n��6���2TO��x�̙�&�ԑa��i��I3gj��¥�O�q�N�N	%��tp7M��i�� �F+��}��$�Od���O���O���+��	~J(�����F�ǧO�r �	��l����M��f��$�ͦ�&��rb+X ���������u��#Zm�֟��i>���fB�Y�u�-X>0�@ňC�./� ��ÁGf���O�O���?����?I��2Z�L�[6�m�&Am���?,O2-oڬN������h��w��\w�R��D�Ng�$X@��"���R]}B�'�|ʟ��"EŬ?�NY�Ѭ�^h��xg*.RȠ� �}�~5����&MD?!L>ID�"�����⇯+b��A���(�?9��?	���?�|(OTMlZ�U&��I�#�\Mp���8$ㆁ[Xy��y�8�hp�O���<5k&AST��i����E��{���D�O�B�Ma����K"WM]����P����KC&�Ze#B+.HԵ�7�y�`�'���'���'���'N�ӟl�<�#v�\�=XH��G"[�,#v�X�48������?!���O~�6=���c,C�W�ذ)rG��	�P4QU�O2��-��I8O��6�~���� t�T��>6�z�{�p������A��d6�Ĵ<���?Ѧ"H�r$��h@H�}F �ɰ�?���?����ݦ)��K�ԟ��	��@�N�?(�H�P$I� 6����`�T��q���� ��l�	P��uS-D07ߠ���2Q���	���s�-s��n������z���'12O��nH�s��(�Ց 땩\�r�'"�'������R�eՓxJ	��"Skd�qh��$�438XH��?���i�O�!L����F�+����f!�C������ش+����$u��F��H����}��$�ު<�Z�bB��R٩��>a��&�̕����']B�'3��'Ė�� E�i���%jH�N��P�_�\��4=�h�h��?����?��C�2=�`0��NJ��ݡ�g�C���	�M���i\�O1�Z`QA��K�&�Ԁ�	_^`��J5[jI�䜟����Y)mrəD�	Sy�/g���h�"DU�Tը��Q�0��'2�' �O��	 �M�W��?Q�>�|�����$~���L��?!q�i��O��'��6M�Φ�8ڴT�Nh�׈�u{��A@&eZ��f����Ms�O��;X�@��6�S�ߙi��I?Qn�y!����crL%�'�|����ҟd�I���	����B蜑-�Ȕ�U���X�T���G8�?���?�G�iN
�O\b�|��O���nͮO��`�j��9�E�v�9�d�O����OD�QpӾ�Id� .�+��<+� {a�h��
��)pj��~�|�_�D�I��	��<#�T�th����/X��m:'�۟���_y��v�hmh���O����O$�'?�D�� n�x:|�1M����'�>�]���%~�(�'��=\� Ţ+��XӔjDv~)�У��N�D]*�i~�O�����R��'7@���J�?�ΘV��> �� ��'���'�"���O��	�M#A@�����,K�B� �7��*��5���?�Ƹi��O9�'�<7-96�݂��
�y�ȍ�W�Y�)�ҕoڷ�M�v�Ĥ�M;�O��Z���
��O?	��Z�\} �}���s�z�H�'yB�'���'3R�'��S�J�&���S�x���o�3�~�:޴_S�p�-O��$=�	�OJ�mz����-(�Q�Ņ�i�Hlx��6�M��irPO���i�%4�6�x��`�k�;lE�!J©���в'"v����ۤ&�B�Am�Idy�ObKJ�xh�5ɂ�N�EB�L��ÃK�B�'��'(�Ʌ�M;�L�"�?a���?a�,ɼ@�D��W�"M>�� �J���'\듀?����'�Йtn��ѥ��$z9`�' H�c��M�r踋���������'��"0�P(e:����m�j49"�'�b�'�2�'��>����a?dA�����k�FA0�z8�I��MCvkW��?��h��6�4�B��u���2Hr���@��
�4O���O��Ĉ 8O�6�b�8��
'���E�O���w��"I?�8��yɸ��ӗ56�O���|���?����?���,�� Q+7�8���o��\�~� )OZ�n�&�&��IȟT��X��J���)��<��y�C�C6/X�0�[�������$�b>�qqN$���0a�%S�ju�@%�h��SQ)5?���@,,���S*����!X<Q��R�����#IG�}BV��O\���O�4���rs��j̧�y�&��f��&E�E_6MK� _��y�)v� �8��O����O��d
�C �p1i<ul�ĪG@�o�^I�i����ş��;��*0��'��T�w��p�wOܾ�R�rǜ�}����'��'O2�'���'���Q�KЄ=�IUd\�BE"�S"��,����Mˡ��\~�h�@�O�$)�HD1rƸ=��A	���#H+���O��d�O��pӐ���HI2�1� ���g�	��䁡#��~�c���~"�|W��ğ�	Ο,��'�2b"�5���|��Pu�����	}yRӴ��������H��N�0B$5
$i	�1d�h�����$XR}��'O��|ʟ,D�E9�r��r��!�f�s��B�md*�"7jlӪ��|��J���'���&�K5
D�Q�G�q#>	�֬П �Iџ����b>q�',7���X�1qVG]U7��3��x5K���\�ߴ��'����?��H�5H�m��	C}�`U�M��?��Sip ��4��d�K[ry����őY�
����wH�w-!�y2X�������� ��ٟ��O�N%���'�J��d��'���+W�~�|����O����O|��|j�{K��w��Hj��K�(�F����V�p��ȳ��n��ymZ����|Z�'��eH[��M#�'�8�HA�W�!ʺ���hՍ=&��ɝ'�~�b�K����s�|2]���)���`%[��I�O��0�@�ߟ��	��L�I]ybnӠD)��O����O��"J�6H쐖$� T�q�.�I���D����ٴA�'*��f�Q( A�PN]�,C�'��҂�̅���R3����3��czV�$�*=�'G6^�:Al��qՀ�D�OP���O�$-ڧ�?�t�69h��A��8p���zA����?���i;��7�'.�zӦ�杹h$��i,��I S�gh��9�M�°i*�6���u�p7l�@��1^*�a��Ob$�1�@�ePj҃/�h{�mC�nL}�IRy�OLR�'l��'�b�~�@�fF�\�T�5NZ�)R�	��M���,�?���?QK~��N�<�A�mL�^l�! �B�>�x^�<�ڴ;���5��i_� T(���)�F����
�����o	�[��I2�0eie�'�ڡ'�l�'�li0j��.��p�ǋ̕R�N-xG�'���'�����Y�8�ٴ7��;�'Kb9�솂GCpI�*ܥauA{�\Λ��ds}��'c��'�nl��[� )f")Ee
9)��H�4�F<O�$J!e����'?����?]�ݮKAN��1�Q�E�j�'�3TZ��	���	ҟ �	⟬��Q�'M�� �� 8� T���,��}����?�����F�M)����'#X7�#��]�V��C�)��1��� ��M&�`�4^M�f�O/\���i���O�E���`��	d��1K� ���8��E�r�O���|���?��88�SMns��C��
�����?I/O��o�A��������ID�4��:F{�H
��ae�!��C���D�r}�|��mڜ���|��'<�^d�4\0Sq� �;���	��V�m��qRS��o~B�OǺ���_+�'N�}!�ƵG�6d!�*� )@P���'a"�'���O��I�M[���RdD�He�W��D�[��1t�2���?���ii�O ��'Kf6͏�o�6H�f�B��T �@�U���d�J@n���J�l��<����سt�����'<z|���O�DZ�Lz���(/zn���'������	۟��	S�4E+e��1�4Q'S��;B�K�0��6�ӝ/�����O��6���O�ymz�}���&yVٲgN�1&�n��G�ߟP��l�i>��I��{��AǦa�|�x�qf��7"k�T����[O0@�f6�|��&�O��M>�*O���OPLde�$v袭��f� _Gu����O����O�D�<� �i���r��'�2�'Q<�Pc-�9q5δBs�	����D�Z}b�'U2�|���X��W,Bv�ɀcL��y��'v~�#���s���O����?	��O�aCf�T!z\6|*�I�;K�X�i���O�����I��P�Ix��yG���$81V�4n� b�(�?bX�	h��ݨ���O���i�?ͻOC���たTx�����6��Γ�?9���?��#޾�M��'�ReYy6\�S$�	X�S�8w�ID,$@�l� U�|r\�����	�����şh3J�2!��;`'�[���p��gyB�j�l�!G'�O6���O���4�$>kp0�2��.A�P�@�P0����'�7����5�I<ͧ���'>O� ��N�5���8����W����a��A����'��eBRR���Z�	ȟ�}�T��7���(X���� �1�:Y	T�Oh��%���6�N*?���Or�I	�{ƌ�<��
�0:��!dO�)=�PI21k�6�?��?���?9A�A��e���h���`�ӗ1PEK��2�����5�����Γ�?!���<>b�2(�������
�Z097B� ?{~��-��0����O����O���O��d�O�Ygb[)O0L[��Ԋw`�����Y�saM�3���P��	�O��dX��%��e|�|
��n>1'�0�����`jb�T���=�C_v� �џT����0�	�|�t�l��<y��r�R0Ì�W���
�^*���&�Ȩ2�X����䓔?�O��'n�%�A�p�HV*�h�ڱʤ��3�|=��0��E�3�4�Dd[A����'WR	i� �Θ�C6����?�:���'��|����b�$�����r�y>��O�R���\8��gGs�0C��),d�`���ΑɛF�����:A�$:�dԁ'�bI���\��q�A#WT�.���O����O��	�<W�i���k�K��(���fM�����s��G46�r�'�7M?��6��d�Ϧiچ��\�	�&]�fl8勆�M���i%��z�iA��]E�m2��O��'p�ao��{*u JY��Γ���O��Oh���Oj�D�|B�DN9~Ar�ш�>N]C�K�E�F �%^#��'�����'�z7=�1#�@�:/������-�\������@ߴGo���O?�5�&�i��� ��c��8q� m���E�D��!7O�B�ї�?��h$�$�<ͧ�?)7�C���q(٥)��]����?���?����$Ѧ%���r�����hP"BF���(�W>s|�`�AOF�3n�I��(��|�=Xe�FmϫB��pQD�B�P�	�\*��#m�fDm�V~B�O�����?i0��m8�\�p�Z�L��?���?���?�����Ov�R
�-6�H�3� ��໅J�O�lZ7$�tv�6�4�L�	�N�

���#'^�O�����9O��$�O��D�%7�6m3?ɗ$� "~���z��C�c#�xs$�+ M'�`�����'[�'��<��\�퉌�`���jE�+���2�[�h۴U�ZX͓�?�����<6�c�n���V8���@ᕿIa����@�	E�i>U�i#����m�~�[ �-Hv���$>w�H�G�iY�I�����C�O�Ob�&565z�F�\I�V�_�( <����?��?a��|�(O
]o;et�2mQ$̚elƯ��0GK_�=1�I��M���k�>	���?	�o*t �l	%�*,��r0@����M3�O��p3��
�(���Μ�b����?H��X�W+V���O���O&���O��� ��=#`�9%üזA��G$~�~��ܟ��I�MK���O~*g�&�O�}� �Z
"U�x��N/"6P���?���O ���O�Ia�g�f������Y`*��8z\5W�=�h����On�Ov��|���?��!D`��٢_���W� {Ȭ�
���?�,OjinZ3I��	�����?���C��I' ��s�T1Q�\2�R�H��Iן��IF�i>��+Nv(����1���� ��EMzm���rߠ�m�g~��OI�e����n��`1-��9�&(R��k�H�����?����?��S�'���֦!����D�8 ���'EO�i��f�P���b�����b}��'g�A�b�9m��ku�ц%�ʼt�'hb풇Z���3O���ļ@�^��O?�	�J��@*v�S1&.-ʆI�/��	ey��'o��'���'��S>q0���wf�`�č�� ��|p����M�s	�?)��?�H~2�&���w���cu���N�)#�E� $��8	Q�'�|�Ozr�'�}øiS��]�K�0!�t�٩i�@4���3O6!�w����~2�|\�H�I���!��B��ẵ�m�~LW��П������IOyfh�n���%�Ot�$�O�	��Ǚ�dO�[A�E	r� X<����$�O�7��I�	$��;��L���;PH��4��������E̘DpmI�!?���?���d���?������0j�t��T��<�?A��?���?���9�>���ʌ'*܈ʒJ� c������OH0o�3Pe��ߟ0sݴ���y7�ԩ.(fxx�GGt^��'坯�~�i:r6�E��	�%PѦ���?�ЪD�%�r��U[���סR%�Z̨���h�fl�M>�(O�I�O�$�O����O��P�y"α �����(C��<!�i��Q!w�'���'��O�2�ώ#Ġ��$�ܧ���a
���	�6z�0D%��S�?��S0U�P��*� }�zaƆ�+h,42F/�8K�6�bW�Y�Tl�O^mL>�,O	b ☴K{�uo��3����Ak�O|�D�O��$�O�)�<��i�ց��'��b��E<x&�q�LB�BA �'�\6�/��<��$٦��4M �fOнF[�h1�ED�p�.��y����6�i_�	�X���O'q����xa��ônH����Ӌ~y�{�<O>�D�O���O����O��?�a"׏B��C#�J�Լz�J\۟�����|�ڴot��ϧ�?��i�'BL+.�� d0i�n\�Xea$���{ݴ�"d�W�M��'��!�r:�@���R�<�]�aBP�]���QeB�ş��c�|2R��ٟ �I؟,���Y�3����&c��-/lQZ�Ɵ���|yr-g�H����O����O$�'�T�*5��;½z�@�)j��P�'Xr�
���Nu�Z$��b��wfS�}�!�բP7�A �;j��Q3@Yk~�O�V��	�V:�'8���L�{j���Ș�S�81���'���'����O��ɞ�M3��D�4x�l<U{赢%(O7�� (���?���i��OB�'��f� �/���"�׶y��T��L�S&6�RЦ9�+���'��d����?}��6@����s�b=�7Ι{��|��9O�ʓ�?!��?!��?������׀;�P��	�@��|�q����EmZ�Mw�=��۟���m��79��w��Y�#?\r$:�)_�#
#��{�"�m���S�'9	:y��4�y2`C�_��Y���U`\��&�y�J]�I�Z��I'��'��i>��I�s��G"��*4�cX ���	П���ɟȔ'@7m_%`J���O����
PT��$> ��`�����c��4!�O\nZ�M���x��!�Vy8��K�Z��8����9��$�1��Īԫv61�$�9��s6���G(G����c�Cw�8d�'�*���O����Ox�D!ڧ�?�� �1��h{0,��W�:���ɛ7�?)�i�����'~"jb�@������p�53PHQV�]���I��M���iZ�7Y�[�7m>?��̝;�i^ �6y9d/;�h%P 1��l8I>q.O��O���OZ���OD��`C�q���jc�7�2|+%��<!�i��@���'"�'��O	r���_}����C�1
��$�[�-TJ��?Q����Ş	 � �vh�"E�H}���3S����~��͖']�$���WT?�O>�+OFysR�ѾZ �|҄����}k �Od���O
���O�)�<1��i��	�'ζ�e*P)b�x�ćW�b!�'�7�,�ɫ���O���O�쩂��1E7d� '��̨�k�._�W��6�(?��nź(z��|��;"��S �#fLJ�(Sg�%|IB�̓�?���?���?�����Ox0IّCL�J����A��R&*\˝'<B�'Q�6M��Y���+�M�J>��	�~���
�/t�M�@������?���|z�ʇ�M3�O��qA�/M��))�m�oq�t��G(�����'b�'s�i>��Iʟ�����za�A
!�P�$i�<5��I��P�'KV6���{���d�O��$�|b�ǂ+6M@�ꔥw.�R⡟_~���>Q��?IH>�O�~�cG��('�\� ��SE������)v.D �Q���4�x�(����O⽋��L+h��yx �N�S�P��1��Oz�$�O��D�O�ɗ�*2����<�ջiI �C���H���*b��::uF�X�䘥�y��'hҗ|�Oo�I��[�F��!���K�R� �@��H͟�����m��<��iCε!ɖ(��9O�Hr/��"���f�Dta54O.˓�?9��?����?�����iA� ��)�3�F�x�v�蓆;��o�.��ϟX���?іO=r��yǤS0?X'�	�k�����j�*,r�'�I՟�џ ���
Ml��<yc͎��"j��د*�,$k#��<a���!V+��	[�ky�O<��ʶT��u�r�^7Cb���Em�*$2�'��'��	��M#��ѡ�?���?�U�R�+���)ԍ�5�,�ȓ��'���?)����:@A��*���#��^�J �'&lT' �8𽐉�t@ҟ��1�'��H���p���L���yٓ�'T�'���'��>���w�pw�����ȿ.�d4V��ӟ�ݴm$�'�7� �i�U:%G�v�@R���o�&� �m����ȟ����7�pMl�R~���	Bi�''��g�KC��@e�}ߌ�{J>Q-O�)�O���O|���O\��s(П^���oQ�8g���ν<	��i[�0C�'���'���X>���|��`�����.��C K�/��ѯO��D�OƒO��OT����wa��aJ�?ĺ�ړ(�8L8�9�D�s���8q�p{$�'즍%� �'����Pg[4�A����6����'r�'R����U�L�޴*](t���Z�����љSU0��N�;�:��� ����'��'P드?!��?	�	�==(I�Ao�:�04�aaG4UkƬ��4�y��'q,��V�S�?y��O��i��NՓ����@��0�
�rᘱ+�6O�$�O ���O���O��?-�a��F��1aG�E������K�h�IӟH�޴8�>}ͧ�?�@�iUW��%H�%�8s�n�}9�IQ�	����	ßT ��W⦩ϓ�?�K��8�
�X�B	�2D�`B��i�`���O ��I>)+O���O����O�y�ǌ�]��Wg��
���s��O~���<I�i��1k��'0��'H�x���Y�fH&"֒�����5u��eF��͟���^�i>����*���z��5$r��f��|�����/Y�	�r�oڒ����LI��'F�'\�xO�4�U���J<M
t�'���'n����OX�ɇ�Jd̟�7��5!/?������O	���������۴��'����?9��JnU
�'��f�G���?���J��E9�4����Ur�g�?��'����2�<QB$9���wW�Dk�'��	��t�I�0��ޟh��[��lӺQإ���H�.nz�B,'f��7m�z���O���8���O$�nz�	��O��{l�	��HJ���@Ɨ8�M�b�i��O1�6�q KvӘ�E%!`��f������<O��r���?1�-���<ͧ�?yeB���@�R�]� L;1�B��?���?i����d��h1��ß�����(KR�� e�1��
S���)AL�p��'��8�Mc�i�rO���:�VD�&�ѓh-�Q�v�����FЇVG�ܡP�6擀TM��ן��D4\TvBN&��9f'���������	��`F���'�VA�'��wP�Ac��cښ�ˤ�';6��-w>�$�O@�n�N�Ӽs��ܫG�u
��C���B���<y���?)��O6� ܴ����B�:���?����5o�Bupv�B�/w�}h��	M�IGyR�'���'Q��'y��ƿ|�ܡ�H��h�@!�����3�MCtG
�?���?AL~��	]:0u��j�HD
�b�\�	�U�T�I��'�b>����ۭ?`���W� ��Yib �sT��l����J�'ƙ��'l�'��z \�AT��e��b�4I�d�	����ğ��i>-�'Q�6��Z���� ��ɁA�C+j�w�R�[���dZަ9�?�W���	ş�ݏw�(Т�D�p��T�R�C��:7��U�'v�
 �F]�H~��;����d��}�F�qcU5�J�ϓ�?a���?����?1���O"����F�r�H�hIъ3YR@��'���'հ7�J��i�Oęn�t�I<0\0:�Ř"�p�3�)<	9��'�,�	��S�'$vml�R~Zwz\�h�ϫJ�H��B( )4�x�c�F��D-�d�<Y��)o�mё��܀��b�-�OЄoZ��M��֟t��K��@1l�r�b�����8rM�����Ox}r�'��|ʟ� h�N��K��(���p7��pLP�1�qG
c�v�����H{?9I>q�a�=@ l���
�b�8BmWx<i��i|�ʀȝ!5��`�$�-�d`�(�$����5�4��'I��?1w�M�sn����̀�l�@���4�?!�5l���ݴ����P�{���?�'c9��R=��T �?��c�'��It�� 
�I�}#��
��T	���M36���?���?��d`l��>r(U�g��K�����.SN@���Of�O1�j\��be�x�	�+EI�@�l	��E�� �0DB�'����P?YL>)/O˓LԼ��(a^�C��8����	/�MS��>�?	��?�U��?7ɖ<�D�	��9�t����'�J��?������Bc\�H%��7#�22���ABH~�o�VQ,����iR<���\b�'���c*pdk�&�Q�ntxL۬�y��Qo���;񂗦UB�h�T��Y�Rls�N-#���O��d��?�;V�p9�ǪU2�cG��PQΓ�?!���?�D��?�Ms�O�J�T�ov�)Ŋ�V ���T�Q7%RZ�%���'xџ؛�J�	�r����$�Q�6?��i�椛p�'���'���=Ѷg��uZ1��i�6�&�9
VS}��'[�|��$�B&8��xG˓#VFt컑��?kH-��i���}U Y"(���&��'{�X�4��&`jl4s�n��`�j)��UY��Gb�+>m��S��/t(�aV`D#�rCz��⟐��Oh���O��ƞ؜���(� Y@��ŝ#Dl`�j���v� ���?E'?��]''z^9`���<��iׇ:_~6��C��DQQ
�j���j���%/R�q�cB՟����Dc�4*�H�O��6�:�d�L�}�ą�7�,��E��o�p�O����O�)ˀ39Z7-6?��{��-�C�&kU�9�6H�{}|�C�����~��|]����ǟd�	����f`@�M�L�M�Y�|�¤T�d�ILy�'b�Z�"@�Ol�D�Oxʧ1�+$ωΑIw�\�*��4�'n�:��6�}��%��'$���WM���,(���E�ehr�]� ��zŌ~~�O!���|��'�\%(���+�܍�w`/,�1��'Yr�'e��OV�I+�M��`ȲE6�yJ�eW<���S��<(C���?1ұip�O*|�'G(7혙07x�ISgLz{J��Ea��i��m-�M���C�M3�ObّWG����M?�1wCkn��b�͝Y>���`�s�$�'v�'O��'^r�'B�� �V��f(֖M3�ԃp�H�[QRa���V������?������?1W��yG��9�3��j��]B������7��֦��M<�|ଞ��M��'� �I��Q�pwjp"�`����t��'lY	������|�V����H��U�c��Z&JX�3dX��J���������jy��u�>]�7��OX�D�O���k�,O.(pe � �l��)�Ɏ��d��� ش��'���[0��<}�A��P�i�����O�d[@oS�����C���?�C��O�#���*_
�ٔ-\+��"��O���O����Oآ}��"q��s/�z�6Y�1#�@���x����O��k4�'�6m&�iީk�����[g�W0$L�=�gc�p��47ꛖLiӜ��n�L�fJ����/���P[s#�g~<�6m�74 L=����4�<�D�O����Ov��8':tє ��NVy
F��3���%�6� �0���'���'��QD/�+�P�80�M�wjP}�6�>���i#�6M�j�)�O59�ʂL|��� m�ڹh�@���N�ڬ�����O��PH>�)O�M�#&�.'�bݘwO3�ڕ{f��O8���OV�$�O�<Ac�iu�H���'���FRZ���lʤO0� p�'�h6+��8���AԦa�ش��$��n{R`˗R8W�tAQO=���P��i��	<Mo`��O�q����8����-p������Y-\����O����O��d�O��� ��Hx~�d��$&�
PD	=ߚ��I��P�ɻ�M�&�|"��K�V�|2�R5	�]���9dp��዇�X�(�Ot��g��i�'>�6- ?�e)�����l�oF	+�I\������O>��N>�)O�I�O����O�����X�ti��K��<">�3�`�O��Ľ<��iB@ӂ�'���'�S6F,� �K	'T'd2�aA21�.�g��I�Mˣ�i=�O�ӂx;�9I��+o�����Vb�9��ht�&1�f!4?�'-�0�D@(��q,H��P�� $O>u�(�X0����?I���?�Ş���ߦiWNK%G\�8�풒��ܓ�քʶX��ɟT��4��'Fb�i'�f�R7C.V$�"�՞y�1ǬXf(7�Dʦu*&�ݦ1�'#R����
�?)��<�"��Zª\�o#�P��9O��?����?���?i���	�}�� ��a�	(������M�~�Tm��@_>`��ڟ��	Q�Sڟ�X����Ū��t�t賑iM&��� CU��rݴT���c3��	ݦT(7�c���#��/0�)���?�B���"m��A���R([��Dy�O�
	e�Υ�.�g���S�/���'���'��	��Mc�γ�?����?��#L�G�^�j�mĶs+��c����'.��w��֌{�ޥ$�� ��"�T#ԡ�K�$���CQ뗐9\�8V	$��;�����C��?���p�8sP"�C׈�ϟl�I���	���E�D�'�:�Ꮾ;�z���A
�(>I0�'XZ6'�8���OX}l�T�Ӽ�n�WI$���T��p��â�<y��i�6m���Uc�)�ަY�'&�1�a��?�"Y�f���p�2Uߐ�y��J>�.O�i�O$���ON�$�O����(X�/��ŚW�Bk9B�!�<a5�ir��!�'.��'��X��勯��H�@S*�T�1�k}�r��,l����Ş5���C��;J "�,ɥ+,,-���hd�p�'RX�X��K�T�T�|�^�0�능R�������72̞i��H ş`����	ß�cyR�f�Y5��O
��p�ۆ|Yp����4W�V�ۆ��OelZO��h�	��M[Ծi�7��!H����1�ɣ'a"�#�D�3��E�|�"�ͦ	�6H�@�>9���;uvɁr���F�'��lrϓ�?)���?q���?!����O���ԑY���lW��X�e�'���'��7͙�|����O�5l�b�"T���.�K���6Q^y0J>Y��Mϧ=S\���4��dp
��p�H�TA!� .�*5�6��c���?��1�D�<�'�?���?)���l.����-
0��2��.�?����\릡��o|��Iǟ��Ox"�`B�݁-���I@.FZ���x�O���'|��'ɧ��	�/ =S�Ǐ�V�в�lř�����F�J�7�>?ͧ	�:��B�	�1�$	���#3&�a���{�R��ğ��Iݟ��)�SKyr+f�n$h��ްT_�E�0-2�L���ַT*���M���>���Zщ	��UD�!ke.��6���H��?A�Κ7�M��O�@�
Q�O��]��!�%fz!YE�
��	�'�I�L����Iϟ����I]AD���ΠR�bD�w��U�p7�B=����O\�3�9O��oz޵Q�]$5�f�Qa�o��
!�T�D�IZ�)�ӛR3:1l��<Y�ϖ�L�̃�o8]~�����<�@ż:����h��\y�O�rM��NcD,h�/e���X�h�1D���'UB�'��I�M����<����?�d�;y
���/1�ؐ0�Hǚ��'���?������D����Q�l�&��J����'���ؒ�8�f����~2�'��U��]"��a�J�M�L%q	�'�bܑ��c ة�/�-��ڕ�'�|7�&JB��D�OF�l�p�ӼSlS#I�Р�[=wU�e��<���?���6� ڴ�����U�uC�?�"��;z4�	6B�w%|�I�Yy��� !�z��uc�2����{�X�D^��Nؑ�I�����s�' ��u@T�V3K���c���
	��\���	��X$�b>�CDΈ��aFU�dt�93�"la�0n�*��)_�e�'�'���;#�l��LP�tr���e,%��������{�!����ޫ9�W+�9Qb!�#'����	��M��r�>A��?ͻ�0���U��(pÉ�~Oz�"�+��Mc�O�=��JG���4��4�wU����.�#{�|�PlK2��,iu�'���'���'��'!"���Mx&ђ�'�̘��P�>�X�� ď�&���#�'	��'X6���Iw��O��� ��øvXЁ˒hʆC�$tr�lr�t�p*�Sv^�D�O��d�O�\�d#|�L��꟨�@�k�8�Ώ/�tiWi�]|h������%��)���?I�&jl�@V	U�#	be��BW�{V)67j�x���N�����S)������?��)�f�wM��
�F>'nnm�J�PjZ<x�'�66M�@�D�O��$S���i�|J���uC"Nאu�B�G�g(03LS���]��4������'��'a�S!�-x��9VǄ�9�L�$�'���'l���T�'�2S����4[i��C��ݒ'EV8�Sˎ�R�����<i���?�I>ͧ��D�O�� <.0)��͟�fL\u��K�O����H�d7�g��I.8\�Z��[@��'�(\ˀ�V7J��y��BǨ�ja��'N�	ʟh���(�I�����q�4�$! |	�`�(-�*��q�ʍ�7MMS���O<����ʧ�?!�Ӽ�v�\cH�� s@�;>EMU4�?1������O��Ol��԰fv(6mt�s#�H� �ȹCNY"�Rlg{���g�;��D+�$�<ͧ�?����ms���(Nc�x0�b���?����?I����[Ȧq�A���������*�Ä$��IZA��R�>ɉ�Wi�	՟��'R"�'_�֟p��b�G��m�5/��R�:)��4���Z�b������)�'I��,�(d�����\�c����o�0h�|I�cO �i���*�?�N�#M�;&�l@9G�D��� [�m�:|�,���J�E���(3,���)rf��/E��Hɱ^
CP��cj�)q�&,����o�u��� �.��ɲ���%Qʨ�Ї�S!8��,y��-S��3~�<���q����9���!d怨�䇳Q�*4n�8�88���<&���RB�|�YR$��_�L����)7�̊4g�SN�`Z�͛!���93 ȧ^_�����	�K#��R� mr�c���c,p�# �&]�Ā�E*b�ZQ���Ŧ��K�h[�}r�'�ɧ5����2�a�c�� ��l�e���d��771O��D�O��D�<eK�;.�h婵hՖ>RΘ��he�����x2�'JB�|"U���`(�/{�8��L!	w�K4��n��b�@��埄��Cy��
h��S�|����d�)
�i�i&Tꓥ?�������^-p�)� x���@7
4�課�ׯS�� P����ӟT��Dy�lҁ]���~=�g�K�3��]X�F����c��u��z�xy2`ә��'>tu���E]��[�l��&̫�4�?�����d��-�jT%>����?����B :]BcGS�Y���arN������0	-��L������ȯS�P�B/��{��npy"�Z�z	j6-Nh�d�'���&?)e���1[�`"��C6%��ɨ'�ئ��'2\����I'H��p��A�� �!�����fo�N��7��O
�$�O�)|�G�Lh��\54S�`�폪-���ҷi�:�ȗ�4�1O����: � %��&@ ���h��wDPm��������,���8�ē�?Y��~2�	6�,��	=b0Y��lX��'n�J�yB�'��'�p��)HD��"�X*W�`K�
b�0�D#j��'�t�����'���}��fb��j6���$0���x�@��<I��?A����L�_����J�o�=��[�>�PgL�Q��?�L>I.O> 9�͞�#�Up�K���!�����h�1O����O��D�<i����rH�i[�X��@�*_�i�0(��+�=!0��ڟL��f�Zy�����$�6���˕��HO�L��X�+����(�	��X�'qK��)�i��}@hC�r�~���_�P�6<n�\&�h�'*V���}rL�=���p%�����@B$̑�MS���?9���?��$���I�OF��q���E�v��YU�8Ã�5v�'z��''�Z����	�	�xR�l�&�.5r���Qr�&�'RCD�F���'��'=�$�'�Zc��j��50��	�%�VF�۴�?��0*a8!%w�S�'t4@�Kf��6�����Y*��-m�'?L�Iß4���\�ş0�Ir�do�7���/ �4��2Ӻ?�J�ξ�Gx����'?��Iū|-�l�rK���t�!��m����Oj�D]H$����i�O��	�Orݒ��E�(-�4)�!۝[$X-��d�T�Sǟ ���D��H�3)<P	���%���*6�ʀ�M�} �T��'�2�|Zc�\pEʶ���DH2C�C�OUe���O ���O�˓c��Ivd\�Uy�ř=~�p �& @� $��jy��'"�'���'���r�[�5�T�Ƞ*��ݺaK��4�bY���	ߟ,��ey� �*����<��Q��>?�XDPB��p|�7M�<����䓧?���5��1��'v��h��^sy�4�@�C6Q��O����O����<i%M��r�Sԟ�hQ.�)XѰ<����&�"@���Z��M;����?1�D�zd����	' O6%3�ӦE40�8��%r>6��O����<���]�S��S̟����?�-&I�0����xo*��6F�;��1$�P��� �-�Z����%�R �#E(R, n��憶�M�)O��Hc�O�=��Ο��I�?�ҭOk�3=v%���[�#�jI�6K��_S�v�'�2���O��>����q�0	�/)�|�3�i�p�Q�	����	�����?ڮO�˓mh��3��3\����
3(���x²i��<����/��ߟ|��/��G�l�u����vI��a�Ms���?9���(��Q�h�'���OѱB*@vfUp�/8�t��U�dF'Ux�O|���OB��
)Mͤ���O�.if,�Yq�>�ʴn�ԟ�s����<��������'G5X3�}��g���Yr%Ob}�b�7��'	��'�B]��'aP%v�aj��_��Ha`�Cauy�O8ʓ�?�K>���?�'��=a���!��Z�H@�W�f��bI>��?����D"aJ�'�ZY�GfN�~fJ��#�=��0�'qR�'B�	�����4�'�,D���E�yc��@���w����>���?����dϫdh��%>uqqb�8��LGG$7!4U{v-��M������4�z��?��_�~��P�b��(��p�U��+�M����?�)Ol��ӯ��S矸�s���'A�jT�k��DqcrU9uE�>�����O|�D%�9O�n~��([���h �p�7�&N$��_�,�G�C �M�ER?%���?��O�)H�iؤ ~�c�X$U� �iH��ӟ��I�ħ�����ES�����^�d�c�tӊ����I�L�I�?�ZN<ͧ.��x`&	�F4@��D-X&_��a�G�i~j�0�'��[�$?�f��q�O�q|�1��k�%!&�L鷹ib��'D���)��)�L���7��D���)LW�H����0��'|ƔP'0�ҟl��#Q��AH�Q�Qy�kדM\�m��h����ayB�~ڌb�@�{鮍�P��RE�&�G"B��(5�4g��H̓�?i.O��$�?�"9s΁69�ty���
w�]:�
�<��?a���'�����b�
}��A;n�\Dy@d�	Em	0�B��'!rP���	�E��'v�"q��n��x�"�FA�:�m���I��?��O2|'iBЦ��c�#�H�U��MP4:rJ&���Ojʓ�?9�j�,���O�T"�Xl$
���S	F4�!�ʦ�?���?A��0���'��Yv� 2`\�(y��<ID%Ђ�b�V���<A�8�B(�,�L���O���Ɩ(Óa�<n���j�
�,�n��%�x��'X�A�g�̑k�y��� r�HCݛg����i�=Nځ��i�剓!��tk�4b@��X�S���A�H�I[��P�Fu���7)�Y����k�ޟ4HI|M~n,u��� A?ͤyS����<6�Y�d�OD��O��	�<�O���T,�	�N��T��8k0$HZ�dcӸ�sd�k1O>5�ɶq@�i� ��*Z�����4f]�%�۴�?9���?A��pw�����'��d�9
�H3��;S�q�?_��F�'h�I�
�������O��d�OB(�1=b�9#���E�r�s$�ަ���*	|ց�I<ͧ�?O>�����'\v~xД�LmPD�'��e�"�'O�	��X��ǟ8�'>�(�m�}n2#U���*V��w�߲5O���On��<Y���?1`c^�	a"$�v+F�[���бK��G�����d�O����<���qF���a2��PBE�u�Y�Ug��M����?����'r 4�"��޴g��;T �T��T#���7��X'�T��Xy��'����V>��	�v�va��M�B,Y��M�ai-�MˊR�'X�ȍ�7M� I<鄬T77�a2)��_��"u+����Ο@�' ��A��+�i�O���Ƅ��e��� ק/���j��x�]��Z�c�럔$?9��]7"`��Z\杘�*�j���m@y�n߲U�6�X��'��D�/?�c�W�z+B�rTf E��Z�Hmoy��"5[�B*�	+��i(T�NӞd|b&8 ��CڴG�0hB��i�'�r�O@�O��-�����G�NQ^4��"[�sò�l�&;Z�A����`�'���y��'�Z�A��+iRLI� �
l��&e�6�D�O0�$�q5
�$��S���K1�# A��+ܮ���ʛdn�nП̗'�t�3c��~��?����?Q�$W��u"`ʅ�8����B�P�6����'\�Xs��6�4�8�D3����eY%��*�$FDҗ�v]�X� � ��x�'��'��Q���V��2�0�gh�O��XP�P�˝Y��͟��Ik�MyB�[�oe�0��eN0�a�F'�e1�T���'u�ݟ���ğЕ'lZ�[�n>-і�e"X��ᎠWw�9c��>9���?�K>1+OΡ����O�0`ǉ(y����GjPb9.�*��n}�'���'V剒3H�QK|b"jX���qT��6�r�"���w:���'��'��I�f��	^�����z]jXP�̕Q�Ù�\0��'SZ� �O_<��)�O�����[`���C��}�ǂ�=�H�HE}"�'���'����O�˓��TM&�Z {¨�v�}�%fU��M�+O��cW���Iݟ$�I�?���O�.M�CGJ!�o�i/<l9�ٟY��f�'���y�[���It�'j��P̭	��Dh"ϼ6��]nZ�By�Ȣݴ�?���?��'%��	^y��&K*8%C���-��?6�6-S���O ˓��O"�3u��y��,J��Q�働.��6M�O����O�8xօ�]}�\�h��]?���L,zJ����b��4�\ۦ���iyr�ߕ�yʟD�d�O���L�lv����bD�z�B9j�Tm��Fo�6��$�<	�����Ok�J�9�meA�R��h�0�١��If��Ɵ���ҟ��I�l�'34a�-�Iv�M��CS%�����-V&����D�Ojʓ�?y���?QU��%#,�+ �n����\�c�`�ϓ�?	���?)��?�-O�x��E�|��F� W�$�0!dR�uͦ9;�����'�\����ğ���	>�P�A'��!�E1\�"m��M[s���4�?����?����P*�fM�O�Zc�eP�U9bѐ����$��4�?�/O���Or�$D3�<}�<�LQ��E�n��S��ʋ�M���?a/O�@�f@�H�D�'�b�O�@�C\���X�"ġ]��t��a�>����?)��q������9O2�#^��ei�
��݀�@K��7M�<y2�B
=ٛ��'���'��$H�>��O�r�{F�W -KD�JVA'=~t]nΟ��I�G6����$4�ӵp�pr
��e� ��P��0�7��%fN4l������X��8����<�aY�S�EBY(/��3A`��Eʛ���/�y��''�	i�'�?��g��U@��B;I�})TՔw%�F�'@��'�(E�r��>A*O����������o%�7�
1����@�h�<���<����<�O�b�' ���R8t��%d��d��Q�F�'���a C�>Y-O2�d�<Q���$(�jTu�$�D)D�Z9"�g�v}+Ҭ�y��'z�'��'��I�"���/ƍNCXx{�֮B�d�ea���ĺ<�������Ot��O�lC��I6mF����Cf���3��+0t��O>���O����O�ʓF�~�y�:��}�gM�h9���C�����i��	ޟ�'��'y�b�(�y�	N�6:�B��lF��連`Nt6m�Oz���OR��<!B/UB ��џ�X�x� uQ�eYW�8���蔞Q�86��O�ʓ�?q���?�����<I,��nQ�P@`�ʎ19D,�Ĉ6�M3��?�)OB5°�]N�$�'��Ot ���G�w^�Q��~5�Q����>���?���lny���9O��Ӟ e~-�Q�W��Hk��]�Pt�6��<�T�G� �V�'lB�'�����>��n���ɐ.|Xt�@�Ep0��m�ԟ4��81����^��Kܧ9�v���ձ�.����K�Aa8\m��7���!޴�?����?��L���Wy2�O�����dYP�R�3�
h�6��c��d�O����O�Rh:� |�{Mݳ4�q �		���0q��i�"�'R�ߕ&֒ꓴ��O���5���t�ƍU���Ԏx��6m�<9��N\��S���'�R�'��`;Aߟ�����$�����f� ���>#�n��'��	񟐖'�Zc[Ԥ���{�-[�\�v�(��OZ��>Oh���O���O6��<I��<%�T�R�� Lq^��mt\N̓�Y�@�'�Z�D��П ��n���ɳ�d�f²E3�z�r�t� �'\R�''�P���c����TE^�>5�ȱ�J�/ ���@��"�M�)O��Ĥ<����?���`�~`̓}����9Ak������L}��'���'!�0=(V�詟R��J&n[x0��A�5����ܗ$�lZןė'�2�'\��[ �y^>7�Ғ���k��� /��#!�H�6o���'8�U�P��fI0����OJ���r�SS��=��Xc�/�"�Q[c)�[}��'`��'�Z{�'L�'Z�i9�hq�����<[����+(e��6W� P� _��M����?���J�[�֝=[2��)��l���V!?�7M�O:��ѡ'��$�O�ʓ��ONDՋ��B{�~	cBn˿j����4F�X�W�i�r�'E��O����Y<K2�`s ��e7�R�­P�`o�o$�	cy��'e��$�V�Hj�엘*0UrV�,��hoП��I某�!�V���'��O`��  �==�b�bqG�	���:�i�'�D��)�O|�D�O8�d�٪d ��/ng ���ƦA�I�K$ޑ�M<���?�M>�10�b1��)�I��I�%΂N
���'E2�k&�|B�'
��'p�I<Ay`�s�	I .�Ԙ�v%Z���!����'�2Q���	ß(���7��C�I�6��}�&.+�,�w"`���'���'��O�-�2
~>!�jR�e^�XS��ݳ&�̩�3H�>����?9O>���?�U��?I5i�;a���I%,@/鰙����d��	�@�	� �'阄��L=��ا!�f�	[8b'��21!�Y�w�ŦI��E��L�	�JUHu�I|��:*�!��D�"��*���3ܛV�'BT���r%/��'�?�'"�Ј�'���R�kB�( ��������Op���O|xR0O.�O��|��y�⍙i�x��D�X��@7��<1���$OǛF�~J��2C���q�E%:xHe��K�N
�k��rӜ�$�O�Y =OX�O|�>MX"���ڴZ���ᅔ(m77���-+�m���|��̟��S����?��oX��s�R9iuHS���S�m��t�]��h�Ix���?��)��8Y�%�̓R��a�b��Pk�f�'��'�����-��O"���xa�/��a���Z��m �L)��=A�\0'���������.��&���)��=���W>TfE��4�?�P̒�[p�'/"�'�ɧ5���K~8S��U�> 6)���D
���H1t�P���<���?����
3�&���g0F�yQ�:go��:C��m��?iO>1���?�UcQ*e�>yIS
ЂGd��$���n�B����d�O`�d�O���Zȡ;�La(�BU�hrR� d˺[v̙SZ�P�IП�&�T�	П���~��C�.ʔ��Cf@��*!�Yx�EN ����O����O �L��I�b��%�/l��$B%{Uv೔��2RT�7�?���D�O��'@r�i�֏!�E�#d�4gx��H޴�?y���䍥_9,9'>A���?�؇{0���@&��Դ�xfc��'g����a
���᠅�4�䠸"�i��I�����49��S�� ��$��k.hQa��LX�MJ$g�Cz�	Hyr�'��O�O֞X8��,hi
�$O8�l9�ݴ!�jqBR�i��'2�O�LO�I�!R�f�kT�Q�i�p���)^��'�����O$���ǜh:�L���K8r�]Ѷ�<7M�O����O���OR}�V�T�	[?qEF��L�ls���{�@1A3mЦ��Iҟ��I�&��)����?���q�f��p.X�&��2P%��X-��1��i��Z�������O���?��4R�9	aL��a4,�kb��u����'�6�ɚ'�B�'���'��s�l��j��:��4j�Z;��(qN�pQ�)��O�ʓ�?�.O����O ��>�8�C�ػ<n�c���!s 8O���?����'lA4s�<��Ȋ�܋����Ee�4"���C�iZ�I���'[��'�B��y��"�|M�W�֚8�b�{U@O�8qX��?����?�+O
��g�L���'�|mHd*�^�`�q�C�a�ȤQҠvӎ��<q��?1��7����?q��!�X��4��4r�͐�fڥgW�2�i���'��I4X���������O2����FAqC �F�N0	 �Z�:��'b�'�RF���yRP>�	b�#�ܲ9 �U�5\�a�i�ߦ��']~l�B�l�f���O
��򟘐էu'\-N��L;��S��}�C�'�M���?1����	eyB�'rq���(�YK��`h`���zr^��P�i�����Es�H���O8���Ne�'��/�`JU�ܪK`�����?t:޴td4Γ�?(O�?��	�T��i)�-
�(0��b 
P�4�$�Cݴ�?���?��狄��	fyB�'�DC6,r����^9q�blb�n	0R����'A�	*0�^�)���?i��,r6���**�P��̕0Aư���i�B��=
`�듾��O���?�1!80��b�
i�h�0gǌ�ZC�p�'� 4��'e��'b�'�B�'IBg)� ���K��	ކ����a��������Ĥ<������?��'�VX")%���vOw��t�ܴ~4���'"�'�R�?������|JQ��qv��t��n�ԓv���A��֟��I՟��?���~r�K�Qx؀a�k����'����$�OZ��Ob��O,P2�O����O���A W��kVcI �<��M�����u�I۟��'�Ƶ�N<���5u���s&iZ;�X�@զ=����H�I�$���K��T������I�?���O��'�k�l���@[��ē�?�)OF����i��j 
Z�X�b��� H4e�cj�B˓/f�ɕ�ih���?9�� ��ɞ�`4JvM�-]f�k�O'd�OQsG"$�I�?O4N����)ď��'�ƕ��i�H�p@�'���'�2�O�S�$l,e���:2�����;W�օ�6�fa�uGx����'��A��J�@C��`I�:%�����o�Z�D�O.���)�*��>a��~�� )��8��x�"����8��'��Mq�y�'�r�'� ���%J�1��G��0��sMeӠ�D�y7��>�����k��Nyʐ�)�
;E~�q�Q}b�:��'4b�'�[��iW�ȅ~�6l2wG�:�
��#�K�����O<	��?�O>���?����k!đb�HX:�4���U&��<���?����D9H���̧Q��9�
��WZP�gL�<h����?I����?A��\�'}Hm�0
�8>�ME�vi��ɫOD�$�On�D�<�G	̢��OZ"`S�eA�g��D
�,*Uf$K Kb�~��;�$�O|���O���Ձa'p�E^�G^�c��iR�'��	q|��J|2����e�#:��Z�&Mwj P�c�.��'���'������T?cg�؞(x�u`�o��UT"��� q�N˓W�h�%�i[맽?��'-���/2��"�M�������rk>7m�OR���2}�b?A8"%X"�d[��4^u��n��G$Ӧ!��ן ���?�xJ<Q��	�L=J2��L*X��	��Ai�q��iQ�!C���S�$��ЂK)�xA�O�"�MocD�M���?���yb���tV�x�'�"�O�����%s��"��S�v�ⲵi���'�����yʟt���O
���jQ�5��i�:�$��D�v d�oZ���2�LG+��D�<Q���d�OkL�v�.0&뗏<���g��':�	Ӡ���0�I����	H��'��ቇ*E.5㰘V���Ԋ��w�F�xPT꓎���O���?����?���S1��qP7hT*�JY�g�S	W�vU̓�?���?i���?/O�kE��|:F�_�T:%?��9c��0�n�}yb�'����������B`��k���>�B���d`���E��	�M���?)���?1)O
�1���r���5�b�"6�����J;<T $�M������O��d�O��X0O8�wD��{��L?B���"CK���ir�'��I�w �j��|���O���;pllm���3�4L`��X5MUD�'Q��'�R
��yB�'�ICJ���7"��$�6f�
P�bKզ��'
,�[��x����O��D��קu��"6
R]�	�({4������M[��?�%���<�M>��$�χG�H� �³l0�f�[��MkĈY)qc�V�'l�'E���>9+OH<��i60j�����0^�P���O�����f�L%� D�d������cF�)c}� 9уɒ2Д]@(:D�l��b����$�CF�>�X�� *$�OƄ�傊+ʈ�u�!���f��7Z�\ #p#��Q��i���ΡwT�C4J?�hy���l����=N��@��&��}�����N�T0��ѲZ:��� \x��5�Jif�Kd ��!5h` ��R'��p�ԸN������X
9��l˧��7f���)%kzEd�2��'���'�҅���'��i�@4��0`	�>Z:�m����Q�Q	U�mE�Q��.9j�$��h�N�'F�bH�(�4� �<����LT�
z�l���SIu�7-ժ3pACag�U>�#� �� r2�'�D��/$n��ʵE�A����I{�'@V�ӷ/�}��D05�Q+Z�x��'�����#D��G�	K�m��'�V꓾򤊆8����'#�R>]�t���:���Va��&ű&a׍H@�Iڟ��IC}�y��E�	�1�G��?�Od��i�Î�$��ɚ��۷HF�\i���v	h�� �Hy�v&7�i�����M� ����S�Er,�GyR�Һ�?�����O��!rw�P��)�hq:"(��<!	�_�zHb��jlxC�P�1�rx���-�ēJq��q��#N�d�!�ܪb��H���W���Ip�D��3&��'��-$�xS�]8F�� /7ɒl�a�,5~,A���	h}*�"b>��
4��9�@��<M�Lœ�(��[� ��HV�=��T҅�ا����O���T�� 8�0 2��.l\�Mh�dٽOU��D�OL�S�D�	),�AC��� �#YIY� B
�'���s�	Y4"�\M u.X3+��0���HO���cAX���J�s���BJ#S;�����(��D�@פ���@�����[w�r�'�h�8�oXP����A��?�Q��'� �	�	&>�d���\M8��   ��A�"x�X�$׾*�H�f �*�@�r�C�6h�92cD�9U���=W�.��L�v�
���.����	-{�ԁ��ޟ���t�'i"Z�H�vMZ��&Ee�;�4Z�":O��=��(�'%��P�]])�9`G�"��&�'^ɧ�)$�I�`�iSi��u�8� �92�tC�	�GJh�r�g��1OjRsGQ7zB�I�b�`u�#��[m4�Ȇo�+�C�	��|��	� V�N;V��^�B��6�-P����a�2�j#UqpB�	H>FU8�3��&L��HB�ɬY{��
qNZ�$��A���c�C�ɘ_����"�?U���e��9BʄC䉳^������K�ѫ��XkbtC䉝#Ę��vU�:�b\yl"!6LC�I�EOz�1����:�L�Y��a>C�I�ua�p��7G�h P!H2݅>D�`Q���J�A��K+�6@��&D��ɗ��
�&L�0��>  ر�*O�a(�M<*�v	��
���B"O���p+��2�q�D�_�m�� �"O�����O"
eniA@���xp�"O�I;�a�+y��z����$@c"O��s��ʕ$X �����d �iɡ"ON���i
7-f��:%�4J�$	�s"O�e�%.��A�b��K�`�B��"O�͋��L�,�r�	
T2%���"O��H�[�C��يQh	y�ui�"OX��8]��	6�KEp��"O��'�з?`�k7�	2[��h 
�'��U")�5�.�;s�ռ{1���'{.9CĄF�w�hA�]8�<,h�'�M����q�d� )C4L�N\K�'���l�%�j �[�n{��	�'펬�G�z��@g�d��`��'��p����=3��< ��C&Eq�y��'�(q�%(�N��X��r�����'/J�J�	<+^&!��E,R�|���'�QP�N$&Q0`0�n�45�L�h�'9@��gJ&\��d��Dۆ;��1�'��#&	��<�0D�S��:SV1��'��h����Jj��2C�,�D��'�<�[4߇���s��W$��`	�'�z��pM��+�rI��MY��>m��'����Ά�m5�S��3xԀ�'�A� ���h���"�@�'�F�2b 8W�<5�Q*����'���&F�akb0BΝ��y��'��[G!R�>�1�*�
q��I��'7,4{�G�
G��*)�#�LJ�<9
U�|hN�9��	*� ���+�|�<�U��T��������]���Sz�<�����w��P�ӥ3�-q���y�<ɣ��2�1��	��֥Rv�<Q6��4����TUNk�1x�ct�<��M'>o4Ș3%ڕb1����+@q�<	'F	�`^`	� �D��*Q�j�<��#ȏZ�F�wgA�dFDKg�<�g�I,IjY#�n >�� ǈ�W�<q���\o�� ��F,ܽ����U�<����%x�*�q��`�h�k�<iF��3k�9;B��B�`Kt �e�<����{e�x�wIL�C$����ώe�<!��ƳH8�i# 7���
��NH�<	˞�Yɰ�0���i9:�0L�G�<� �����

ufpS�ȡ	j=�!"O��{2,O*h��q����3�l|��"O:��
��Ox��!R� �v<rQ�"OҐ�B� ю�"D$��v�$�"O�h[A�ԥ*�FQ�Q�_�I
���"O��IU�@�#�f��V:-�p-
�"OH�(��{�H{0A�Ɍ���"O���"D89v�	8�j�	���R�"Op�ЅbZ6k9�+���������
Y �E��i�d8|�2�#V��%��`���y��E�
����T@L���(�5�~�憤�D�=E��oY�{��I���>Z`y����yH�$�Qiȶ>�.�Ȅ���ɒiu�}��'�4�� ��@RC��D@5x�TU���
>g{d�	bH!:*xкTI����B䉆D^������`Jv�׽&i�"?arJ��#n>��&OȊHW�`H2���5Q�+.D�����ۚ@�\�R��J� ~<��uf,D�h�C�G�T�����FhP�d7D�h��N�/�lS�c�=�J�Q�,1D�(�J��N��a1�UH��{�%<D���F�:�Bd��a?E���ps�4D�t�g��1E�:ใ,.HB�Q
��.D� J�:M�2؉5B�.v�tI8b��O؁���)�'r`}�&��*$d�yZ U�OH��a���$A�x�(�
Q��8aZ�Q�J9[�h����?I�	�/�|���*޵��O��S&e�8u�Z
���i �:EM�`�6�G�D�t)�y�M�d�kL�`q<��P@�Q��l c��77>�K��C]�V-2��N���z�M���Ѵ�6\�u��D|�=qdĆ+v�(���MWh��Ua!�_!����0�Y(K� DJ���T�7aϱT�\a�*,�2�)�Ջb6\��?,��)j��'�L�h�iҷ{5�������:�?���Q0~�P �2kF�QB�ER�jދ@%�'��d�$�Ծ��Ϙ'k��פl�"L�6��j��N��<��+�(k�3d�V����d�4'��;Ì�'aq����Z�a�$�e�[�7�H\R��'�4��a�K�wD�Ay����K:r\��b��e�P��b�7��ٸ�򄝏2b|�qb��a��I����2�NQ/,R�fK��fV�=�)�##̡QЃ�TE�ؤ�����&�;M,8�@��[6��x0���<�7l7�Tp��@ ���2�Է[�h<�E�' ��@�� n�H|����3D�?!���W�q�8��Q?5LH���l��'b�(А
 �Ϙ'�D�iV����3�K�d����F)���y���;7?T�I�@N�*�3�I*Um����	ʕ=��`Y��Dd\L|��@���|��,<O\\�a�P�M�}�cF�>�1:��C0ML,H�A�P�f�w�I�z��zA�B2ID<�j�����?TVR��ʎ�I���G{��)g�~9j���T����O?�V언�p��Ӽ��U�C!=?1�l�}0딇Cx>PT�ۦ\h�c�&D����pf��O�M�e�Ff�B�IbI+'�|����&?�����|3��� ���y"���J��u �ڼ�@(���	$bx�	}���*J�8t�N!��(OBP�+DD��B�L��h#��ˆ�'+����(� E?�Y���xA��Z&s�@BF�G�t�X��'n*�H��͚N1p< �#�
n�����$��$�er��C,\�q��ɰ'�ӉSE:L���N�\q�"O��EI�Qu]�#�-3���x%�'��]P����Z�r�0�O?QR0�K�I�X�x���Re`�*�
�V�<	���%9�XRmV�w��貣-_Qy�AI�]%޸�Þ��p<q� `�=��m
�q��E�4<a~�A��P�_��p�ƃT�`�"�HR��5�4� ����*��r�ra��R&j6��	A,�ѓ�� 24����FK)�����F!���e��a�1�X!/����U��������
\i�ᓡH�Й�NG4u3�/@sȖB��1')��`���5DΐU��,�6�tb�T��$�Ye�x����G��,1�#�+6XhB��U��x�薔�����F��}4�$(!(� H�*�e�I(<��@IAA����o�ڳ��B��'�'�qO� f�E^�
�(q�r� 1zn�%R�"O6$#Viś��e�c(��֙�<*Ð7h�qO>�3g엏S�n�q��.|��0��,/D�tiA/�V�Q��`�l�\�#.�	�,q\��'j������ +��R���Ѻ
�'ꢰ���^�J�@��S搨�(�+!��S
OV0����}(D�����{���!c
x)�ՏR��OA�9HAl�\b��J'��	�',5�t���ORV���N�
��A��i�NPE�8}r��Z�O��)���q����'�?u7�a�M�2��OD9`�a�`����A�Ih��g��hǯ�>q���X�'e���,b4p�$l��m�d�q��A�Y.>I�!�E�}済 *��k�X׌#K��%qm�#b�"��Va�=y����-sp��'
@^IhJģj�Y�4�
�p�셔��<{����m�p�'�y�)�3n�lT��#�3GӲ�1��y�1�
A��#4���R��v��x磈 4ʨ1�Bg��L�
�i�O��SB��7z�d�'%N`�1����вgL�B�lC�rE��� ��;��=뇪M@:�Ի���!�x�����hZ��Z�{�,�f��X�,J�k�&s�
��q%��Q̤X�l7�{��3J�E�ջ�U�h�R-`�cA�kĥXҍ@4?nT�W�a\8)�"O*���j�K�*��������ҽmV����[Kj�9���*\*6��<��>�.�/CȨ���� �����L)az�'���dL+er��r��I�N�z�cuj�@5� �ͱ[�9��_)v�^��]h�Z��4���`sㅏyВO.�I��Dy�����
]������ڲ֢�H~��i�1�j�Ӄ��:��J��K
?�zqZ�ψ�C�]��
(�8��E��E{�Ii5��%QY���ψB��\�aP�`�d�AT�V��hkʧN%IF�Ob�1�d]8���s�$Q:rJ��"N#V5�1m�-�f��,�11�r�� HRd{f���X�gj~�@�A��(��d� ۰
&F� 5�P�A�C^v��C� ��	SE]�p���8�m�8@[�"N0�9�D���
�n8)`u�#h���L��'+�t��6��UK�~�1A<I;P1����e� B�e�5Y�����Gc��hYD4�X�')��Q2������-��} �Iώ;�5Ä��w�"E�R�����O �k�)+�R�N4ɒIS�Fu�P���ABÏ(r~�ŊqgL'j���B�8d��� ��'`����N�49 �ղJ�zE�FA�Y����$M�1 ZL�t�W�d������).Z48��ĐWjeK��Yn��ªʧQjd .T�QЀ���'/@C��S�qT(G��'^Mn �wB`�H�K���j���8�``�R���V����݀FbF�	��C(W�a�pN�>7~,C��
U�%IhQu�ʑ)CK�,>��SQ�K�t��S��V|��ǀQ�	�hA<(Z��<i挤:(��+˭N%�(�/�~x��B+ʯJ-�Ӑ#��2��i�p���w�<��B�/x�� ��/J�9�G�1#���R����!L֘�:�C3	 � �<��b9�	���ܴV=��ZS�P%`6!�'!��.c���`��#�*��*�U`.C�	�:ˮI�T�ת��N�6t� C�I-Vi`���~�Ybť_�R�C䉗@����hۨ)��8��"ڕ7�C��'*���3�_m��)ɇ�
#�C�	�q�8��\�y��MӲ
#J*�C�	J��l� ��-M��r�!Kg�C�"���׌W긨{7��$[o�C�(0�p-�Q쏿��HfDѩ%~C�	3��|����'.����b��5�C�I�WxrM�s��=n�6�����8y�>B�	�6�h���<�R���-Z/�B䉟M�����1|(�d�h�C�ɣ1T�(�i��L L�P0�Ӷ��C�ɄQ
J!z��O@�§��?�B������+s��� ��*^*C䉢8Gh�(B�
�NB�Do"(�X��zLD-;ɇ�f�y��q%�=�ȓO���W�X/1F"�0f�\��DՇȓz-ā��U����M%I΄�ȓ�0;�͟7&ʝ�g��z���:9�H��^�=?�1���P�a<�<��9�%1�-%wrBU�ӮB<O~����N��@��鏬#la�[h���̑@�<� n��Pu֩�5���E)%
e"O��������Ԥ�)@��C0"O�,�C59|�6��e�p%��"O4B�D4Co�œ�!�E�pŃ�"O"��3Μ�V ���/�{ 4ɠB"O�Ȣ�˩Qcb�X�#	1r�0�"O����/ ]����$�ψtR �c3"O������Rڨ���K�	C(��"Ox@Y7c5rJ(Y�VN�<r$� d"O�)���$R�����X8C����"O� pɎ+e	M�eYE`IS�"Od�:wꋁ-R%z 瞣?&�Щ"O!s��*g�"d@G�¢-"�( `"OV�8�HL!�j��6K
�Q�@2�"OX�"�aP�~,f��v	U����Q�"O`���	��pF��5�2î�h�"O�� ��צIVh)E)�
{�$�S"O@��"
ؠ	SL���%D�(��ɰ"Oj�����<�u�E�X��\�s0"O�K[�9��kY=3���6!�C_����`U�q�Fia�*Xu!� � ؎h���8A�������!򤑲qȆ�Q�A��"o�.I�!��٫6~����84�`.P5Y�!��їx���0)C/��Yyƍղf�!��=4Ӳ����+5��m1�,կdS!�ď�SSi�+�J%Ae��"?!�D��+%X�mͯZ4� fY6�!�D�,p|��k�+�(vˈ�+���4�!��<.@�Fm�P����r��fm!��M�!_����/-5��]���#Xb!�� '��p�����qk1�B� `!�d�6�r�FN�;sh�]!�D�%/�`��6��C��u�&��G�!�dL�+e�T��?J�� &A�k�!������cA � |�л�ŻGT!�$�#!��B�W�Byr�&��6N!�$GJ<��֢ėI��qD���_!�$�c��%qr`�!P6�,HV#
 G!�D@�yr��� N4g|q,�;>!�D�K܆��LV�/f8�MM# !�dԵ��p��.��XL�FA\�!�D��i�ٛ�$�)W�\b�\;V�!�dϻ �� 
6�N��8ɔ̜<p�!�dj����d�>H��\8憰An!�����%�UD��2���H�#"7�!򤑕&J	�֎��.t2ܐPI�#!�� Ű���UT��)�g�^�!�d����EPQ
�HRr��s�Rb�!�ГY�ݢ�'�l= <�ׯQ/@
!�� �,7�� &kѐ+=�󮀥y�!�$ԲR϶��엇{�8�% �CB!�d1�0E����i�x����:1!�$�{M��·"�?���a��/5/!��	�fa¤X��b�X�0)!��,����cȚ5�NLJFcgIc�'����p�|��&�^��ԑ�'� ���Y�p��FT-]��s�'�D����6P\P|�oŅO�  q�'���e(4��tī��IN��
�',e���X%���*�tR6Hr�'* �I#����oЃ?�<H2�'�Ƶ*6�T�G���^q���D�6D���u�ٶwg�1���2"z�Ѹ`�3D�� r������Sg*
�o��B�"Oģp���(
�b�n�s�4�(�"Orl@C�^�K-R3�䟴jʲ��"O�5h�'���ٲ��.㎜�R"OH-1��0_�X� �w��%;�"O|h�bN�$/�IG�W�W�j0"O:�A��Φ4�n�Y��O	1¡��"O�e��W=�Z�cw��6Q���J�"O����
�+F,XP�E��A�P`0"OVX�7.�*���*�(J\��u@�"OJ� ƯG�G?��D�t�9r3�
w�<iP�K�r���K�,ph���p�<�&�Pj\�l�S��c,�l�<�Ue�7g�je���C.r�y1`�c�<�bj�e,�`���N�=���H�Ʌbh<��kY�my�$ݰX�(��G��;�y�N�p�Tm�Ï�!S�&`�����yrd�D���H���@��3U��y�#_�pԜ��A��3�XM:�)���y��U9�.�#� H�����y"�ݱn(�Ϳb�>P{����yb���0��d�F���Y掔`�G�y���'1�� tIA�U�-X+��y`�m���
ef�8G��:ŉ"�y®X$9����ǍגKy0�������y��آ���`�W�B�V@*��]��yK�d��s�!ـfRx�����yr��Cw: �P�+r� ����y�o׾k���
��P)q�ļ[�M֑�y�^5;���r�N�b�T���ʔ �y�H���Ȝ���R%e�~D����yr�����D��7^[< ���S��y2L��
�+�>cɒ���^�y���G+P\�B��6+��A����y2 \�gn�E ࣓>*i܄�3EU��y���z�!d�6 ��pK���3�y�i�$����m��d�H-9!�8�y¬�3[���E;_Ρ0R�>�yR�6x���1�^U�<������y���&J�}�U�[,a�BA� T%�y�i߷;��`�-�}�Z��ͅ�Ps�%2k_�<��X)���|N���=�bT[�h)m���k4E��=��@-���Od�а�!mE�pH�ȓ\z��س��#���Hd�F�]�n��ȓ �jp���;JҪ����n���R��驢"J#Dm\Ѫl ^���ȓ!0Ty��R&�<���� lꡇȓ� �/�Sղ��aK�!�`�<)ŌCM)�<"��Yݴ�9#k�[�<�ƢNh.MC$�^,U[�H3�Wb�<yu�]�8HpTNB+- (�Z�W[�<�M݇X���r����s�8�
�*�P�<9��H���vO�J�q�	�I�<�s�K���@�K¬|"9� �M�<���%u�s����#�U�y�J�Vք��O[�A0�`�M�-�y���!F~�)#N�*=�Qr�n�y�K9{T
�b��O/"מ�6�J��yR"��F���a`hÍ)���%ۍ�y­;��Y�AG�x,�ٛ���y���]֪p��Y1XH' )�yM�<U	�#uJ�0M~�̀7�D��y�(7+������M�P窚�y
� �)���a�N83shQ�kܖ�c"O�y	3M٨9F��2H^�����"OxȊ��.�P���ݮ_ʰq[u"O�����E;�~��6�1`Ĳ�`"O <)��πa�p��!��o���#E"O�2Ǉ�gO��v
Jm1 �c�"OHɘtJE.% j���"K�|����"Op�R f�;S
�E:bб(��<��"O�xgP�7CJYA��ӄ>���hb"Oh\A�.V0{�E��${�}�u"O~9��(d�Тv!�U\ }8�"O�p�&��bS��4JR$O�xQ)f"O���#^-5�����<A��)�"O����55�������O>� �4"O�؄��[�
�D�ӟ.�E�"OZ��a�S���Bɛ�E9F	�S"O�`�
�?��[�"�-ú9�"Oz�ɇ16��u+�!i��}��"O��@oJi���%I�+8K&"O��P�I��8�$Jt�\�H�u��"OA��a��;ndx��L�{�v���"O���S�ߴA�ɢ�B (���"O�,:��׫-0���� �bw0�h�"O����#ߤW�h���\�Sp�1�"O��X�'��,����@��(n�q9�"O��G��
,P������sg�ظ3�'Mў��L��m�u�W�f0f�h��1D���0�&2DI3(�_�\PRa.򓞨��i���GR���$x%�B"OtӁl��zp���R����"O�p�)Y0 ���9)B��`"ON�
e�In���Y��ݥ3�HT��"O\�Xq`�. lh$�(T:/$��{p"O6�9���BN,�9�撾><�}X�"O���D��([����@%N\u*"O�2�D�)*9f�Z+Ysٰ�Ґ"O�����	}(`��u��r�Z6"O���"��'f*�#��_�{�굑"O��F��f�`-�X�4rp�ط�Ii�O�����
]j��ꢇ�5�$h��Ğ$S�ƞ%/猙���	?�]��!�"�i��
$#�H h�'9n����e��| [" j���1��
v�ن�D���e"�8rI��c/�L���Z'��z��ڈ>P:�j�j 9\l؇��8e�ТO4n|�������pϘ��ȓY�˥�L��z�	9pt�T�ȓl*����
�U7p}
%�� �4ч�H�@�`��2��9
��ExHԅ�l�f Wc�cd�E׊X�����]�>�X��
:�͒��M�D0�ȓPC�ԛ�cnX��D�99��ȓ%00�VO!w8E���+�+<D��;�+�*^��SC�}R Y��	3D��PD0�����(�+x� ���+$D��6
r�1��
N�Y4�6D�ؚQ�0Ȱ����3\rQЅ@4D��̚V�|5ْc�]\���'�1D�a�
�n���k"��+����0D��z0Z�6t�U{�bب 񆕱�3D���gH6�
��Ժ �'@0D�<��썄~~�X��CV~|��WD+D�$�R�
Aɮ�R�k�J�%D�Li4�	�X�R\�'�v��h�%D�� �,�����p��걧��}]f�K�"O�嬘`E	0�GY�H?���"Oh��Q�,5�����kO/��ҧ"O�l�a�I�2�d*1kԨ-���"OL|1T�ss�X��D-f����"O�3"eİ;����d��R�Ƶ�"O���5.؈��Z䌈ie$�A�"ORi�$Oے'İ�a�D�L�ʐ8�"O(L�Ś�%o�p���K.>��cG"O�)˕��kQ^�*�L�"��r@"O�̑fe����bs�@��L3�"OTI���<[N��a�CV& �F,�"O:y�Woݔ%��c����q)V"O8��nT�}�t{��_��"O�Jч'}�ƁK��#/��x��"O�����Z;d���Ϋg�1�!"ON�$	�C=�,���ϖ�a
"O��7e��61ްA��k�B�KC"Ov��� �̥K�H΂���!4"O�<��"��4ކ5.)c��=k "O�@�H�E�L���M� 9�fD"Oz-�� ]ar9�D̀)s�Ib�"O�����L.���!�����
F"Oʁ�#�L�
��)�	֍<�xm�!"O��B��̛Y�<D���D�H� �"O2)ЗIBZ������Ŕf�$��"O\aa�Gk���-�4Xޤbt"O�<(֫�	q(�%8�-� U�-J�"On<P�f�,H�jË.##�1i"O��',޴k�Dm�C��1�$�"O�MZ !��|<�PIE#e��*5"O��(`�?z4�d12jX%Q���"O>uY0�$�%p4ϝ�-�f�Q�"O-[��_;Y�dC%[- ���c�"O p9Q�Ft�]:7��Wmbt��"O�"��pt�x�����P8�H�"O�y�@ �0rTcֈ=Ldٔ"O̴�f�	,>��6�^���@��"O.�X�^u��P���*�(ti"O�X����)5Vd�q��t��X"O�9��ar�iGaV�f�z5�a"O(y��K}@��"cR{� ��"O6�ر��?+��k���;�B�X�"O����Z�/��)"��|�2H�C"OR��͇Nv��@J�|(d�"O.pq�����\-����Xf�i	S"O����)�(�T�`%
�]�U9u"O}Q0@�Hn9��@�<�N�YS"O��B���yE�+��(F�X0"O.�+�jD)x)oC>�X`+�"O,	�B�֧z�d K�Η�f��W"Ol@�����B��0��K�	�Pq"Oఠ��\$ � �k�r��"Oe�� �<K��y�b�E�-슸�2"O�QI��B�;�h��OP�K�,"�"Oحj4!L�O�����('�ْe"O����*Ю%K�gF<�ơZ�"O�	����i.H������z�ٖ"O�ʃJ��y �h��ڇ5-���#"Oz��ժ�y�8���2$�x��"Ox�H��A�?���y��Z0Z �P�"O�t�B&+T����Z���[�"OҨ+"��p���t)��J�"O���`h��W>��8AM��r$��"O� rP����\�Z�̃Y����%"O�m{4�Q�T|����^��i�e"OV���(�B�"i"W�ħ �~��"O�MJ�g�[ZQ���^Gb��"O"�acDۭY4�Q�+��vc��JF"O��ǆω^��B5@��GI��"Oh��E�LS�-��^$ �����"Odِ�M��+�8��6#ǽ]*����"Oک��N��Z�(�"3%�8"O|�شO[r��ٹW�Еd��[�"O�R֧B'D���d��ȸ"O~lb�G8X��!b@�0�.)`�"O�`ؕN۫Z���X� �~�n,xa"O���C'L��ɣe��\���"O�Œ,
"��Q�� ,�B�
�"OrpK�AC�&*ze1��W�~�PtR�"O���R㏡���C0$�+]@��""O���,	�*�PQש0d@PB�"Oh�S*�U�,�R�K�ifzx��"Or8���O1%�(�Y��	F_|��P"O
M��M��X�X�CG��#NF��"O����U�I�(���%N\��"O̪f�Z�su*�8ÃϡonL� "O�Y�A�	9Z8T�#��S��-{1"O� �nM2jW`�"�
q�#v"O$�5�[2w�%�k����Z�"O
٠�[9�JT9�oW�J�J��"O(��W��8�d����)O�~SQ"O���"Σ>�=����#��09r"O`Ȩ�eE0\�PE�����F"O�-��+ �.¸��c��E���:"O���	C�2����l��aq��b"OT�ʓ�
�Q:M��L�	"�"O:��������C�MԾ/�2��s"O�LJ�NW-#� �r�G&���97"O 鲨��m��ܸ��?:v�$��"Oa���Ѱ[�f`8�Na�K�"Of�3g.�?�����N�L��E"O�!�,��������9h1P"O4�Q�ǯyζ�s�iԕn�j��"O�u!1nN;����ȕ�L�u�G"Ot�Pd\�^�8���':~2�ݑq"O:E�B�uӂ�c	&��إ"O*�X��\^�D �͖.e���"O�d�����_�L�@����w+n,�"Ob��5�Җ����7޸0'�=:!"O8jC$I��8�ɛ�N�~��U"O��"W�Z<X��H7%�^)��"O�|�B&�Iֽ@d'�5��`#�"O6<���ڀ�^�a�TtB`��"O�Hh��6��Q ��tiF 9�"O@�B�Ȁ+8�A��Ҽ{Z��ye"O�T�Sg�?)�6�#�#����[�"OjD:c��W���%$O͖�ڥ"OJ+���e�4,)&D�(C(4��"O�Yh"f�R�f��䘟(��"O��{�L��*V��b�ħ�R�23"O̡3!�ُB�2]0s�]Fn��u"O�PgHA6F����',F�E�u"O�e�7�q���b� C%Uj�!g"O�Pb`�I?I�t�0��7QlHI��"O�����ڷ1x�!E�BR<̻�"O��d�_�k�<m�'��/?*��c"O����P\ެX�"_�Y6B}(�"O� 6�g�qRD����+��@"Onř���Xˡ/�K�8��"O���b��e�~�A"�
�K ��7"O���?/�9b�N�P1�p��'d%����r���Z�k0}�JH��'v��Qږ&�T ;󊛭g��'>"926oR�M�z�s�ꈵ_錥��'N�q�~ �|cC�PM,����'�`x8��7G�h��HN%He��r���hO?��O2u�T�R��W��9EOQw�<�r+� 0W�����\�:�<Z�e�G�<� +�(@��A��ȊE�D� w/�A�<��c���܋C��8N��Bb�z�<�@[�J��I%��D���"�x�<QR�P=	Ԑ�^+�z��B!�uy2�'����S�L1O���if�)G��}��"O`-�� ւC�h	����|��	ZT"O��C����r�)Ң� w���a"Ot��rd��)O$8���X��Tȡ"Op�c�ܠI&����T ��Xp�'�1O�̋��P:Uz�Yo1R�d�S$"O�d�'I�2|m��M�,N�D:%�'�!��r��
��$P��,�b�0&�!�1ajxc��Ǐf�jp1�K�w<!�DM*�r����t�<��@��M�!�DM�S�u�3�J�0` ����p�!�d �2y�d�-2L�������!�$Ԗ��8jB�Ⱦ?�ၥ�@�-��d��Vvd+b��7�M�����B��>v} ��Μi�~=;v�V�B�I:I88�M�g�|ي�eE�l��C�I�p�Z����<�*���cC�S�C�	 &��u���� Q�`�SI M@�B�I8 �p!a4���)��B����)�hC�x��(�z਱�E/˒ՄȓhJ4��J&�2t�F�(RBj���U��bM�*?����#c��Є�w_ �1b��:Yߊ �&��~V*0��A�����L��\����Kך'��(�ȓ	�0��N�-<wn�*��@���ȓ-��0� �05E��ʕ�^�=��p�ȓnC��L��Y`�?s)V0�ȓ7, �VA�*p�<ȕ�4_����	Z�'�lpkDU|l��f�*^��x�'[�ق�%��;�-3$V���Z�'��v�_'ikm!/��K��Ah�'�xd٣��*R�R�r�엪B� ��
�'�&<��m�C0���%��<�
�'J�-���!��`c�R�4�������*�'3�0�� '.B�@����ρE삭�ȓ1"�}�#�G�tDXqgB6g�Y�ȓE�"剧lE�Xt����Gb,ф�*�Vx(7C011��`���SYR��ȓB%D��BkU����4��`��eDLʔ.���j9��հ,��(��
@T�� ��ac̏4&��G�'>M��
 C]ȱyP�CU�� �:D���S/�z{HXrD�7mh�X�D&D�x6��`�N� �e��[K�%��e!D�t�H��#)I)ΑZ(���*D��Pd#�7Aa0����R� r�i3T���T͂�s�4]x�EO�sN�T9�"O�Ѣf��g���c�D:j����'�1O���܈d|�!�`�ua ��"O� �<��i��@ zQ-G;[����"OֵS�Ŗa��c��Z�8�2� "O��j�@�n���8�"WO�U�"OP�����6��ձ"���� g"O�����ȴ4s�;��D�C���"OA�ᝧ/�4�P`)��3""OTPٰȈ�4"NY�g�w{D1�"O��0�Z-[U�����"�0�"O*��R�9�rݫ��̊[�ċ�"O��{�r��r��[Mt���"O$�	R��J*b�� LV�#Ր��7"O����=FFp��=1N�B`"Oԉ0 �K*`����Q�CH���1��0LOԄȳ�^,�R胶�ğczT��`"O��X�@�~��9:��3�ؔ��"On0�
˜�:�Q�I�0'��% �"OL9�#(��l�ڝ��g�fY2�"O��ī��t% `�V�5�Ա��"O���W���)�!{��ĉjaT�a�"OT��t������U)�E��$?LOxY��S|�he��gFޑ+Q�'7!����#Z��Α>��y5"[�!�d�=B
8�qҏպ|���S���<�!�d���<��&ô0>Yk ��O�!��Ŀ��]� �΍ZZ֬�1��!�D�~�4���$B���w-u�!�\�XV��P�ʹ9)R%��.BS��'2�'[�	O�'��$���J���x��P�x(����h��ə"�xy	�ͭK���т�TC�I#����ɀ,u���%G�\JrB�I�>1���t�
�&h����
@�B�	%x����L-�&`j��^'�B�ɥj	��Y�PF�Ɇ�xLC�I�]�4��c	�I�`� �X�e4t�=�-Ox�?9�$ˋ�vD����[&|:��j���U�<I�L���HX�/���%�>m�nB�ɢV|����c�m(IL��C�I)o��jl�-���D
{��C䉋A�f��2�F9��p����C���1{é��=z��q2'��W��C�I"f�i�Cg�g��ٓG�60Z�O�d�OJ���O�#|��eL6"�0�l�_� ���_f�<��ٔ8�Q�4m�Z��KP�Ni�<��&O$a�ƹhdZ�?�����bK�<�WJ�{c������}&p�b�}�<Y�g�2ev%�rAS�0����|�<�c��YH����ק1g���	�|�<)c��V�UGS�{|���@T�x���O�bH����/��(��.
3����	�'>>�&J��z�脪Sg: K�k	�'�fU��+|CjXP 	eߦ1|B�	�v����Ԯwm���q �#l�C䉒|��k�ȍl�ذ󃟒��C�+[Έ���R<v����%K_�(��/�S�Og����a�m1z`�3�#B��Xqg"O̭҂W��L��c�B{j�2q"O��y$(���=�d�^(@^2�Z�V�F{��)C�r�����-�`E���ً@�!��òb���R��Hp%F J�O���!�D�ZY>hY�hא<��B<��'$a|"�DP�
)(F.�	\BP����'�ў`�'���R B�zZj #wO	Y��l��'K�h�҉�(�����bD"N�؝#�'�h(&��b:%�Ə��E������� �s�?>�����̄����e"O,uIE#������ۉA����"Oġ�Gm�! QQ�?GId��c"O�U��>?�TY���*�"hkq�d1�	ߟ��'�PaC���O,��a�h�Dl�
�'�x|�L�$�&)��ā�zm�u��'�|aSG��S����a�1<���[*O8���O���VA�uRL���yI�?�!�DE�{�4�t�Y�;|w(Ɋ�!�䎲i}�T ���2D)r	�+/>!�� o���Ȋ�����~�!�X����CpZ�5�$��X"D�!��ob�=Q�	|���6J�!�$��qr$�A`*5�ej/A�!�Ε*	��hç��,�̡�4��V!�$ۤ|�J}�3(�:y�=B�ه^!�ĎѨ�,Vm�.�"�11�O��d-���r��fz8� g 5�H���'�ўb>�'׸�R�)
:���L��h'(
�'�\u�1+Ģ;@��OY�Z����\�,%�T�'�9C�䎛i�b��q��
P��4"Ofx�HJ���A���ഴh&"OP�1��-cd��p�],��Ђ�"O��;�%I�)>h)6jE4d��@*s"O6p�3��+�b}T/�gs��3GOz�a��N�XA���^�S���9�	=D���Wk�Kv�L�h[/ ���9��hO��I;R�k��ūn�b:1� d�C�_rn����"F�z9�EfK0^�C�I���]��m��6��M��'��R ~C�?>��eB�ѰjS��	3�'C�ɒ&dR܊3o@1Q�����C�n���O������;$����q@)3�윰k�!��cy��A�-�5�)��*]��!�d�Pt����$Uz!rA��¸R�!�dۮ[p2%dB���x�� �!�ɧ<�$u���	6X4&+@0{!��V'!E�)�A��7c4�	��J J!��5/�;�c�� %xA��O��Y6!���!QVp���<����K'!�$؞jE~�q�ʷs3 ���C�n!�Ͻ-+�\�Bc�{��`��y�!��]%@��%@>h�ڜ[���"�!�d\2:v��&�H.C+X�Va���!�$��8*�Z���9�{���h�!�ׁ�0�H2&�F���1W�!�dK!`��A�DK�uѪ�a�nO-0*!�I-Fp�W���d��q�bcǓCm!��y�.� !i׹6�,\��!P�MY!��9�YJ3��-��fG�M!��Q/_��u���
0�x���:j7!��_�[��*��1r���rml�'�b�'2������;'+ �i:�L�
I��v�|͊T	T8gu�IU*D���ȓm����X�bQl�3��ղ%�(D�P�7劏�1vؘ���w�1D��Xp��"��p*�R$~kp��/D��YS"H-xh�����E�4%c�'D��[�G�0O��M���܍%��l�R�'��G����]�ܨ���H�\Q��͙\'nB�I�%�4�C�*ܿ,ؘm�P�M f�(��0?��l�5k
�z�!�o��19� _�<�S	ֻC��tY�oB�VB�sR��Dy��'w���'ܫ(7T@#Y=f&��x��� �U8�AŹ.�����A����"O:,H�(ԅ9��!��D�	���D�'��'�r�'�ў(����/z|JI��킛G��R&f�y�<� �� v�!�.�1��(2	~�<����U��4z��M�`�֌p᠐z�<0A�)"��2`��%; �ЅLv�<��'Q Y�p�˚%I@0=�G�s�<���ۯws ѐׄ_�!�a{��l�<1�,ĳG�D�C�A�q��E� B�]�'FaxR
Z�+e���@NԲD��y���,�yR���D����f�-{~��dA���'laz�a����ڷ��1!��l�S�
��y"�S0q�;���3l�1�#W:�yRHO���B1�î/���`R��y��9�J]����~���KC)��yR��6{Ӕ�)0/�I�h�R���y��X�in��U*�9����[5�y�M�/{�K������yRR26n�'��4�B屧�Y��y�ß7N�0yP�S=p�4Ӈ��y�ÊV�H�B��D���
g����y���0��9�M��C0�ҡ���yR�V�KmP�����:4Dj�Pb#���yRB>co�u˂�R�&(�0񢡃��yf
��.I��
�FY��C�(��<��D��t�\��r'[�N�����A�!�F�
�j,�GD�E��s%��9!��/:Pxm���K�f � V�Y�!���4.��j#H�q��5���GLg!���=Ǒ���/L�ճƍN>�Pyr�L3p�V���m��Jw�$� �y���E;2����J�F��T� ��<A��d]�<႔*B�P�h�����!�W.6��q��/$�
��@G� �!�䗾t�hz��W��J1`<2�!�dF�FX�g�"h��%��Ӑw!�D�	jeQ��I��"Y�sEY�n!� ��i����X9â�}P!�Es�T���Y\�� �"+s!���Wg�鈔��S������1c!��&B~!{Q�óQ8�����<!��	w�D�c�͆�*rP�s!��`�~��`ҜC)�����x�!��)=n!ҴnG�wo�]����<<�!��q�b����Mbnʸ�``ҼJ�'5a|��ǆ{>�$�V F�B ���,�y�D���������>o��jO�-��?i��:JŉŠޡ�Z��EなDL^���'�5�4'^4��p��LI�'(��'�J|Ka�0�����Q6u$��
�'-\���E|Xx𛖀�{05z�'��XA���bI��!.r��+�'��ڵ��?�
��Ua;jh��+�'+ܘ�@LۏJ�,��ANf���	���'p�>�I�t���s���2������X;9X�C䉺
4 �Х@�!��Y5��1_LC��v~��pt2F":��¼:LB�I�\�>�u�ӸGT��Kf�V&ʓ�hOQ>A3���ҕ  
�c"ΑKA6��+�S�'l�V�z�n��L����A�,�މF{��O-p	{��C�t�]�ѥË>���#���2OH��� nnZ����;�"OB%X5��T_��(����I�r%"O�P����h������xyr"O� �(tNB�VJ<Ӂ�F$j3�=1�"O0%����LӔY�N}��q�����O���*�'~%: (�ܵ1�H�ڧ��7T��UD{��OÎ���	�%T�1aɄ���0�'_����E&zJ�i�A��]��h�'t.8j�I�\ry���5Q�^� �'� �
 ��8;�^mkЬM�Ih��Q�'�y��K,�XA�n_�4�@� �'3�M��lL L�"��p�>.'����'�J9��'�x�k�fUxlN�*-O8�=�O��	�{�씨���*X&������B�	�
D^��X�M���`��� ӸB�	4$�Q���6Y�$��3R�*�~B�I.A^�s��@�J[��B�O�X�jB�I��ʹ��OK�|���QHdB�ɩ�6Az�d�(8B9��HU7Z�C�I�~_L�G(����*w֋�n���O��6��?E�<y"L(,~Ёakׄ�e�g�<	�ˋy�j@��C]�F�|ʄ��b�<ٗ�O
wi2XZpM�����΍a�<�wоZ���z�W�l;-LEh<��k�#E�$p�� WhHA�mP-�y�h�q�@�#l�S���U,^�yR�� ẽ��'6M8� �wh׊��'�az�f�c�B��Fg;I0��1a$����<�J>E��-�;vpQ����FQ��ٖ�y�̰B%H��W$�P��������y���;�L%�ƥ�K��(!M����x҃)g5�g;}���`� �vX�O�q���u�΅�v��B<b�'�ў�G|R��DD��!B	{aĎ��xX �c	�'�N��h_�Aj���cͅn���I����D>��ӧ8����Ӟ@�Pi2Q��3"�@�ȓj�,���U[��Ń,A� �ȓ��f�#'�2$��BH1µ��IR��+ԃG5L���hAf��ȓz���#g��a锱�W��,G��%�H�	D���'��P���6.p)B.����i�
�'4T��D�!�6A�h�L�"�'�<񡣢��M<b%As�0*Xe �' �ԛ6�T1d���A�M(T.>�#�'J�L��P!"�e�d焳yk����'_naaAbډX�P]#$��7D�-A�'���q�M1||ڳ�Ք'V޵X�'��5�
S���$���iIP�'�l�S5�		B����𦑍5F0���?1a�Y(Sr��D��W�iN��y�j��TB<��A���'
7jbj�ȓx<P����(���dԽi�L��ȓ!wj�b �X�!�j\����]0Z�GbZ���|z�F�"(������̏|�X����p�<�hO
)��L`���p���/�B�<��X)B��u��jܻr�ԙa�AB����
}�Ji�fM<^�$�b�<'fч�6X��c�<_�݋v뙒o0�ȓI>��#�A!"w
8r.�la�ȓjkԠp��T"��������]����P�k��^?i"(��� %l�"��+D�`��J�+P��4L���p�&7D�d���܄;`\l��K���) 6�'D�\k��R�t <h�$'Pb�mvA&D�����ԙ(O`X5��$��!c7D�d��� ��p"�/һ3�*e*!D���Ƈ��K�q��32��Y���<I���3� �I�� 	&J%��s�ݟP.�ѫC"Op��	8�`]K�&��5}��J�"O~��� ��:�dX�%�+Lֹ�"O�Ih�+̪3��D[ě:8r���"O�kK-_ 	���u-���!"OD"
���\q����7^Q�b"O��(J��I�<�b≲A��hr"O���I*#N8@"��1�[��"O��*��� e��u��,K�Te*1"OD�c)]<	���K�\v�س"Of�C�� l�#0/^�9jr8�"O �����(�FH���Y�����"O⥐�(��z�$��Y�G�0a5"Oҍ���2HZEpvL�~�hya"O��0��d�T��d��|���!�Z�����<Ȑ���זK��4a��݅5�>��0?yv�ox"80w�N���ㅂ��<�7k�?R8`eM�g�8HHs�g�<���ޕ&�N!�Aؖp�fP�g�<�ĬJ9>�<�הG��p����k�<��h�&������րy`��j�<1�,�!H��ȋ��e��^�<)�çj�f�I���!��XZb��o�<���AO��8��FThV\��h�<9p*ԤXgj��g��2.ҡ�,e�<�Ta�,<(1� �n����Ϗj�<aǃ_5phLrD)QtӌP�Ԥe�<Ѵ��?���
3�s$\j7�]`�<��-��.���_�|��IЁw�<�6M J�E��.J7tD�Q`q�<���/i����e����)adX�<i�o�>X�DPF�
&����TU�<բ�>0,)�f�	(�F!&bWw�<�P�յMք��p�z~P�0SMAw�<�J_65�
ic�*T1x�� �w��o�<�Į	N���h�N��)�ڑ���i�	hy�X�lD�d,FP��] ���$\�=X�З�y�!S��: �C�RN�L8���4�y2�B=��
�#�>ʅi �R��y���3��$4q($��oC$�y�-�Pf1�B�-�p����y��^j̖�q�������A�y�#O�V��Xr6W�%@CQJ����?����e�4 )JgA-n���g��y��s�N4�E�l� @9��Ƃ�yb�Ѓp����@g
j�n��CD��yB� 6����s`��y�t��C!K��y"� 06��W)�q�؍����yRN�3�BkCѰ��eO<�y"B٪ H�#3Ɋ�e���P$�]�y���>ltM�-V���s�ߢ�y�O̢O���P�S��ϡ�yK�i��q�F�\56}���S��.�y��d �(�R$)St�R�R�y��T"�x������\��y�޻0��1�6�Q�Npa j'�yR`	i��ȁ,%b8i��_��y��0�v�H`lV� ��sCG���=y�y��Z%�X��'k[�qQBtS�d_��y©$E�J�sa���A�&��y2ć�;�h�.�|(zY0�Cѧ�yb	S�*eʭsw��y�T�a��
�yb�пb��YO��oTrd�a���y��܎N�b�h���=f%���a�Ӳ��'!az
� �(Qq��5���WE��R���'`1OQ�q�֏z|�`��IQ�����"O<��U,�G���q#/�F��l�"OP�g6w1ܴЎ��|� j�"O�	;��I8x��xe�G9f���"O0I��$E�i�����G��ʟTF���ܫj����@f.9FL@��ˈ�y"���U�Bꞣ����uc��y�"�zk
�R�-�v�� ��y��= %p0Q�CA�iX��S�6�y�
6 xb�]	Z�A�R���y�dJ�"���q��V�f�I3�Ρ�y U�|��1�D��#��-[��K,��O�#~*�c���P�3� ������W�<�dO ]�\�ׁ� w(�A�FQx�|�'��Yk᠂3/ǖ(y̆2/.�B�',p�eD�U��c�&Dv{�@��'��0�2Ù"E(<=A�Àp�*��
�'C"P;�ҥa�ک9�
��B�	�'�8d�PC�Gv�z�f��G��A��'��u3���M-:(r�a
:+88�'�^e3ǭ�/)52�pgIZ2g%�
�'|��b���$	|�	��7m�B��
�'�p������Q)iֆrH���	�'6H��p*C	7�(p[�A�:d�d]�	�'J���F�P�,���!�I�T%�i�'�T��/�� �b�ү9z b��O�<��3�Z�3(�b ���"O�
�c܊X1�Q$G �aP"O(Qb`�/s�&8�E��[5�U["Ox����^%�0�cg��Ib�"O����bġvmvx�lD �b{"O� �SF��$����P	�v0ZH&"OTA���(/��m��C�B{F�1�"O���f)B6��dj�,�8n(�@�"O| H�E�p
�c�+^�H ��1�"O� s�f��a,b�B�,.A�<��"O�%I�)��%j��@�%�2$@�"O",�`�O��x�̉>&ՊQ��"O�xч��H�>�k]�#�n�3�"O � �%¯ex!��ĚX��9R�[��D{��ID#���Ȁ��l2T+�X�!�DW4��C&�./��w*?.�!��L$Z4j��Z�İ
I�G�!�D'y��q�d,GzD1�VH���!���t%��T]���R!�#b�!�D�v���a��J\qqO��v�!򤓋;�Sb"�\�䐨`��!��۫%Q�-�s��r�>��M-�!�DA�8�V�I�vnQ��Ã!��
c�p�@F�qY�%Ⱜѻ`�!�D��'Q�����c3����BVQh�C�ɺgE�`��
)X���F� 	tB�	�GZ*�� *��<n^E!צ��'�B�!A	�4���~�k��
5K�C�I.24-J�A��Z��x(��'D�8S�XctҡI���جc� D��4)���NM�5�VF��4��2D�P��i��Pq��΀�OJ�W w!�ãFB�@�2�"8�:�i�@V&J!�B,!U��
�"F�\��a����S�!�L6����Y��RI�`��!�d��B�*��2h�w�\فO��7�!�Dd�0ؑ�������o�3�!�� ��!.��(�8�G�}4��E"O��1���G"�P��D��Kq"O�a��C	!�.����&a9���v"ON���/e�t\��[�N��"O�u�䌓+�h��a�I=��c�"O2�i �
�d~�#Da��
�Lm	W"O��)�+��0�y��I�j
г��'�ў"~ҥ��A2����F�*	�A�����yR�M1-���2b���N;Q����y��� >leSWB��K��d�alP�y���-i�$����,K��!B��yR'�Yb�{�>0�I�)A�y�K��Z�:`�2B�8W;�IY�%�yB,�?_`"Ԡ���|;d�A���y�����6�2
Q�|h�)�)�y�	�
��U�E�6����W8�y�R45<�j�_(Xf|#a���yG�T���b��L y��M�ej
�yR@
3Nҝ�רW� Фux��	2�hOn���O�܄� w%���t�X�-�,�[%��2LO|=#�n�� S��Q�.A�k�\��"O�Mٴ���S?��)#^9x\�S"O`�Z��
bb|0�D֩~��P"O��	�;xf�Tz��Rf���h�"OV	{�#I TB&5�U	�.�7"O� �pፙ?�J��� � d�4"OĈ�RJ°�;���<�����"OFu��R?���fhva\ 2�"O�R��ˑm2��8���9`L�r"O,y"���X�q+T��<o58z�"O� L�ǌe��g�!B��)3"O���UBێ�^��"�Ȟ)@�
�"O�wݨ^
6؛�)�A���8��'���C�i>y���@�a�TXCᑿ>yR�'N��y� �b��p��GnS 5�v���y��U���]��.��l�&�Av(Z�yҥ#1?x�`2	&p��:FhJ��y���	�N}���G Y��bR��y��|���1�ou$r(�y�d��?�F�9R��z�d��ܣ��$:�S�On�K��;��-�g���K�M��'�<A�E<\���"�W�\���'UNe0)�'y�!�2B�'^x�b	�'bB9���B�v/>E��H��X�\H#�'Rz���hH0pn|a�!���Ȩ�'t��S�\'�q:D-�#"���
�'Θ4S4	#}r�y���;F�����hO?)R�$�B�CB"U&A�K��B�<�t)�[�b���^'k����X|y2�)�'�nu�cmH'8ߞ�a4�F�T�V4��C���k��58P`�I�S�,�P�ȓPB�DM&y���7�B�Ĕ��Bah-R5�Y�ArJɊsM�����ȓx�5����#p쬠�D�)�j���^)]�D��
$� ��4,̤Q֎=�ȓYK��I)�N~��/
;2�8��ȓ0%v��e�R�?���ㄟ+�P]��bF�qW傭vݴ!�7č?$&%��A{4\q��ڻO�Rp)�g�i�����&>|��G C��(�,�W|�a�ȓ%䵱Q=	
�(DoAC����,�\S�OtL�i��Ė����E���Â@�=~�Ad&Ȇk"X}&� F{��t鉑65�)KVi�S�aAEH�4Bh`����?)�Ʃ�?9��?a��z��y� ���c"�[����aΖ4A����"O0(�ee��BE�$ K.D?P�2"O�Y���όD8��(C��m͚8�w"O�8��$�s�Z���ٻ��`Rb"O~-2�(�9�yDC� @w� "O�;�o̗���jC@�nfV�b��'fў�|B�'Em���獜�$�ԮE7�d��۟L����->�m�I^~*���0�~��tH��!N<1�#���̙�ȓd:p�d���x��l�sx(���̚��T�QD!�� �wԎ}��:�¡:�FI�.�q$�� o=�<�ȓIٮ��	������ȓ�|���X�B?�d؆�HhĦ���_y"�|�����`E2�΅V�h�)�IEojC�I5��Jb/<;�CC�NP��C�ɫR�p�!%��!M�<��o`�~C�=���1�a�d��8�q�ZA$C�ɷ&�d�Hq��c��qCG�4<� C�I�I�Wj~$�`�զ�),�C�I�+�ƌ;a�
Ib<H��;Tm�C��o沠 ��!��[tc��2rXC�6󰐳v�Փs���颊�&�|C�I�'�@x�B��5��9���Z�d�B�I�v��D���h.ɣ%�6VoxB�I�*"D1��K�6�$I�P&�)AjhB�	�L�(����ò`����2�3~=tC�I��T�囅P����a��0~~B��j3���^yƤZ���$���	�'QR��&d�"�X�q,��2YD=y�'-�F�W%0���D(�}��:�'��J�
�1��QtKތ]>�R�'}�ะ�\�m�^a�3�K:�(	�'`<,y��I5xC(��"OH-r:X���'Y�M벥и�j�$�ҨV�NI0�'p6�(��PKd PC& H�z	�'�� I(Q����kw)? l@+�'>�Tac��*|P|��3)�5DX0���'�T�2�hުb|�&��H�>1��'f$��ӎU�%B"T�F���BF��'x}��ʷS��|k]�;I\��'g"1�G-�:\���O H
�'����E��?Va��S=,�L��	�'v6DIS���
�� ����(zc	�'||d�2�նh��k�L͏!����	�'�>�pk�K����Hgc��
�'����6�J�j�r�A�!�3�T	
�'�ıa3F�9�:9ZS:3~4[�'��r���|�bZ��	�|��'��2!��J��B�Ë�{s� ��'^d�H��ě0�hܪ���y��!��'���aD���,U���j�.} �'SX\ad&P4&�3��F�eن`�
�'�B(Ѵ��� ����7iA[N m�
�'���1a���E�>a�g��" dLe�
�'$ą�/��S�B�"7�pL��yr�ґe1dCC�.r�Х$A��y�L\�e!
�	\88���E�ϛ�y�aY��(U�Wa�:Aq0��@Ŕ�y�,�X�P�����8�x5	ѪK	�y���Q( ��Uj
���I����y��S[�2b�&`�T�4	
��y�%*y��s"Z�E�N�D%@��y҉ �����Q?=��Q"5����y�CN:n|	�eĭ!�P$Y��2�y
� &����Wj
����D�VQ	�"O��*�ˆhU^����	uO�<��"O�Y��(� `�U�h��04����"O��j$愗q�`9��V�(2�1�"O����/�0{Q�<��!`�����"O�S�/�%�Q	���l��"Ox�`�I�����JPs{�ݓ&"O6}c�oE�rDxr�߾}�&��"O�4��*�{��e�S(;�jP5"O�d� .�@�Bi选�.y�|��"O%��Ts��=���6Yv���"OrAEA�P�m�V�@�9rr�T"OjQxfLލ� �%�N�sbD� �"O>��	�8��H�������d"O���w�B�Č�D`��.ы"OR} �ڽV� ��O8-V�K�"O��T�<;Բ���dG�"O؈�cI^CZByJP$��b�@*#"O��a�ŋ<Vjz��Py|$pG"OR��u X�8}�Y�Ո�b����"O i��)�����IAF�R�j�"O>-�$��?6����Ɂ�g�BУ�"O��4� ?W�a�.w}lY
"O()�'ՎW��۶L�Rcp�е"OFmr�@F.ST���e�%U�|��"O���(W锨Ie��R�N��"O䌚�o^#��(*�㚜z�L9!"OD��D�P�V��%J�MR/�ޙ3"Ov��f�Ƽ4,��3��I���"O���SK�,F�!����g�
�YU"O���؋8��\A����5WrM#�"Oj���P;i HPJ7 .̥�6"O�y;��<e^���"��QT� �"OZ�8���W��\)ЎN,xP"O��rbo6wL�x���ҩ�0�Q�"O�tbV��^�f�Pc���f�J�XS"O
}3sNG�j������\���c�"O�ڱ�N	&i�4��U�{ҁʢ"O�����7N�v1�\�US�x�"Ox]P��H!7����:<�#�"O`Y�R�S�isz��υ���2�"OrdK`P2k�(8���q���r�"O@�+�hͳT�ik�.N����"O�A�pjԁc��k1̘�|x0���"O8-��
�p�0�j)0`�4r"O2mxRc�:#��QهG�+?a+�"O���K&\�8ڷՁ_#6�0B"O��6
�pP�E�L��Ho"O������MtVM����}��	�"O`���D�$��EF	�.p�@�"O&�h=ˈ�b%`G�
jH4%"O�� ��9\��If�Q1��P"O,4K�j�$�x|ӆ�,qE2hi�"Oj�0�����h}�"FS9���e"O.����ħO�B�����/}zr�"Ot�ȧ�F,^G���FA�-�e"O,ܑVI��F���zL�	�  AA"O�i��bT-8�J�ӡ�'�d�t"OV�+Ю�wZJ%P�i��M&�Hp"O���F����TbU.h��%"OFTb$</���a�F8R�
���"Of��Q1�Ȫ��3K��ҧ"O�	a��ф6Q�i�5)�8���"O^�BuC2'5llfW1H��s"O� Ԡ���ښE����N�0-&�"OTШ��#ZP�UB�ͪ 1�w"O(�{���t���'K�"�5;r"O̡��bG�d2�A
�9J��,:"O��z��0
����aJ�6&讌R�"O:��ӇE,ۣ"��p��\��"O��[�$l5FTPtc�g�¸;�"O(� ��h�Upb�[cz�j�"O,�¦�G�v�fx��YFDX "O�9b��\* X�F���T�H�"O�Diu�B�s �!�"�f��r"O�eH2l�*oY0]���QkP�j�"Of���PV�� �-vSX{t"O�%j�JI�Y.D��b_m6p9�d"O��BB�2[q�}�!��sDP!"O
�#NO���@Ѱ��9"���"O���m��3i0���E�� ,��"O���
�d��M��%W
�h�aD"ON(�RNV	H�ޙ�v�7�8�"Op0!��39�]P�D�*;�	XQ"Oll��ДvAf��A�G��Y�"O��e- /K�蚀���u�d�%"O�-�W!�z#�d�p�g!��\�z��m�2���l��&�!�D�p�j�C3K�-8�ޕ"!C�4�!���HN����`�;N�ީ��o2u!��̓7:ъ4	���
����A�*�!�$�f�ص@C� �phj�(�n�!��L6�J4��:&�]��]o�!�D��-1���2`�y���9E˿xt!�ą�QB��S�����`Q� *�!��Y#r��i��A
2�����ϔl!�$��D	Z��s.џ|�&�S�d��Bf!�ǭ\bb ����'t$���X$i�!��#sXm��)M�$"��d�� &!�V�]=�ēV�M�?"����
!�X-B��{E"͞���4	T�!��U�`�J�fű]8l�i�)�!��[Ha�@�T:b�Z����l�!���,\�p �U=1zX��B�;!��%��9į�Y@�c�C�;,!�M97Z�(8��4  �6��=%!��ώsed�*e�́{�@�QA`��J�!�$Y	q�� �9����G�ӥj!�ĝ�&�Z9�� ?Z�$�s�mO�!�d�� T�PiҧI�|��U��d�!�	�#lz$"5$�W||{g��6�!��Ds�D�3յ{X�h𗂄0$�!���.#>��"��BPG8��0�U3�!�$	�U�����(,4� ��\�m�!�Ւ}��Q�I�7l&̈�7�
6/!���)LBUǭX�/-�x�GG�c0!�DH��p�a��˛���V��f~!��׃�>ԣ�nD>@��vN!��G,C6�(�'K9O��D�P	!��D&RE����&�p�Y��T�i!�d�|A��5fI�1��ɐf��d�!���k}���b�/W��}�Ԏ�'=��Dy��'�������+5�mȱȕ[�ޱX	�'(��2O}��3V�_�S�4<3	�'��X�RS)B*E(1(Ԡ d�Y{�'aXp �Mܬ�a��A/0N9�
�'J�MD�X>_C�T�H4߶ Q�'00��f��0/�d���R���#���>ʓ��� `��B��)^�̴`���e4(�P�"Oڡ��ҁ[��l��²��X�pGyBj&�')K� q'Z�S��ŌLcH���(���jR)�sT��9"�A�4��4�ȓ�0qi�#�`S��[��*T�ȓ_�����DRTFX��{��pD{��'Tt�8Wl�6�X[p`F/�4��'�݁Ҍ�}��������?��*�QS�B��S͚�끠շ)st��'�ў"|*R��$���I�2@� �'��t�<�hʧb�H���?H�4[��px�Ex��� ���eϕ'e�E(e�x�#A
E^�A+�N�G�J�b�;�C䉎׊|���S�:S�k$ɖAS�#=Y��T?]Q�д=�vq��+^�/��Z@;D�x`��G�U�nآ���4.Q���E-c�b���S�L<q��!��h��,�>�li�,ȓ\L���	B}�IRrd��e�K���<�!
�3�yH��L�:���.�v}���\���O��~�Պ��A�d!�&�ܺL4�5��J�\�<1�
W�� �J��uB�D�2�U}��|B�*�g}"��,���z���j���i�>�yc�%xpI�F�6.X�D�'�M�	�'(���v��+�<oܭ|����"O&�2ǂѰg��bP�21{�I)�"O���v䓰i/\0dV2�,�h��I~�Ie��x�-�4���J�H��V���>XRC�	>;�� �d�A�'�0�	s��h��� 3m˄[ �� �'��0S�'Q��:A
��HҎ��RQ`}P�`�p�����>���9����#Lq����g�q�{�^�L�Po��9tH��P� B�΀�sY
=��I}�'�"����޷j�:53g��G�����>�#}�!�K&xpj�:��$4��0�JY��B8����eH8+A Ɇ�8�ژ�E��,��4����O=���U���0�M��a��@K���6�!�Q�r22͒ �ޅ4�Z�b��E��p�Ն�ɛNf����e����ِ�+7�C�	2poH���9q��uS҈3Z�yE{��9O�9����7:&`�n"c!����l7D��ڶE�b�:�
Q��XLn�lt�@���2Y5��9gG� |��y�ȅ6�
���<�� I����RŔ-I��H���ě��B�I,_뒰X��Y\��4�fg�&p~�B��g�i�/��l���q@e$2B�I�F�qC�/1�|��%Ԑ]�b�d��P�'��:�F�9���D�v�2@"�4Z��	W�'�iD�4�	IS��AeQ8E0��,���y��'Aܖ=��@��2eg������Bܓ���m��:}��q ��2s�igѩl\��0?����r�E�#A[�2c B��)��O|�[ v��&c]��@�υ�Y����I'��d�>Y��@�@����%Y��u��o[S�'���=�'C����H�*mL9i��!,:x�=������F��w�,	 � &
��Uoݞo\�0��-�q3,��L�c��0� Ȑ�y�?��9��V�<w>I��*t@�Xu ğ]�C��4R�� -��f����wǆ7��n��hO���D3��p!�;_�x���, �V���He����CCc��^!94�%:p1�>�����W��\�+r� G[�4!�K�1��'��3�)��U;�E�`ɃV-t�I��	j�!�$�.9�v9kC�H8	%f�bUo٨m��O�D2�`�IX5��J߂?�q�M�?)��B�)� Υ�&��+��94I�@��Q��"O@�Fa]�s�X���R.��$��"OF����KȾ�+�&�"u��tӂ�'����;#�.%�|Iۦˆ�ՀǦ!D�P�c�N�j�aaP�fF����G�>a���S3|.��*�/�$Q�0I�[6�"?)���PcR�mЀb�\� ��k\H�O���D�k���h%�9zl}���C!�D�;�V�[cFm䎑y��)!�D�i��@�˅>�x���N,xQ�`���/~B���v�ĉOIjA"C��f_��P���ȟ&�0���U��9�W ���v�Y��'�!��T�l�+�(�Y��r��+��D2��z��~��S;W�n)���O!m�	�E�A�ybM�V���2�E�gG��0%���yR�6g�YF'�-,�"iS��ީ�yBI�\�P�e@5&2\��0�y�h��ٓ�K�!�XTB�ᆫ�y2(��'\���"!���dH�$���w���O���CpD�ds�8�R�5<� ��'Y��z�A�\	��cl�N� 9�{2�>\Oxc%�B�#u�9��X�7J��G
O�7�I�(<���E_-xN�D�5���a�az�D��X�B<���tE0`˃���!�U�ØmAF��oB��"�!���2y���ʊA<�y�"�J�\�!���H�h�QV6o�n�	s���8�!�$U�9��xZS'�i�8���[�(�� ��ɔ���Fk2-(s�ŏe�t#�"O�i�� �+6��Ħ�%��Q0"O
�"��+^�*$�3l���"O� ��ː< ���#e� c��S�O��j���zJ�]r�g�?6���&-d�܆�ɲA��ā�τ8�tS�G#����$l��b�8с �7�
t��!^;+�jkfm?D�lH4�3k�i��iZ�#V�Sv�>D�T��+���U��&Z7Bf=[�<D���$B�~�<�$���p�H}K� :���<9�R�x\�,�!�� S^	:�G]x�'�Q?=� �Ӑ�P:��Β+�8�{��8D�ؠA��+'
d)pҁ�Y�>@X��<���'1����&N!g�r,A׍�8'`A���:lOFm��%W�r �)�u턣UQ����
OF6��7+�"�ؒ͛�=s��e�A`�!��M��� ����7o&�"!�Y5=��x��	�)*Ƞjv�	���Ό$O�>c�����)�ӇVz<ਖoE}��a$���2��B䉺2�@�"Jj��A��M-��+cDB�S����(q��H�g@�Җ�¡nB䉢'��d+l ��"H�s�K3=4z"
O���I$l<����[-lf8��'�:Da�S��y6���}��dX�'���R�2D�p�䢖1:��1#� R��!+1򓿨�>��V�Kň}���9Ex��Z�>O>��U��8 ��*��W�*j��z��Ëp���aAÐ8�P�*���p0��O����Ԟ!�0���"�<-��m8���fh���C䴟����'	�Sj�aʄƐ*6)�tJ�Y��B�I<'V����r( �(Eo].F���$?�S�O���:�I� (� ��(��
����4"O 8�ƩU7�L�����d��8s�"Op=pvMؑ*T�-�"f%w>���"O���V���_vVy�CE�9 �M!�"O�5����V:�;����$�4�qV"O� p���l͹l��y �M9���9�"O<U�� <&t����T�j�"O������}�e§�/x��0B�"Ov ��"�.<��V�G!>qqw"O�-"��|�P�0 �2X��"ObX�2�OȒ�;����#��,�"O:�"��8D|4����3����"O}����]���"ЧM�+�bғ"OZ	���ο~�J)pW���.��"O�0�d��W���rC��rx^��v"Oƨ�g�/,C����薓-Z��I�"O�\y�YmT B�	fQ��÷"O���j��8c( Bvd��q+R4rP"O(J�`����碚�U����"O��pSƊ7L���V;N��5�@"O8u�g��KΝ#",�:��3"O��-9O|L�qIC�R��]���yi�	���cQ>=�HXs")N��y҉��2̌�ό2�� �'���y�HܶK�̸#"O�-���kG��y�䎐o����6독 �R4� c?�y���-w`�J�[�Dը�E� �y"�#-�vE���*u������y���1�z���Je�2 �qʄ;�yR^�d2��p�T�VѪ�Dd�0�y�M�����+�%�A���y�h�%�����Y� �¡���R��y2H���SRbj��Ɵ��y�i	������J:�P��EV��yRj��h4<������p3 �5�y����F�`u�4�	���F���yR� �,N�4o
��H�/���0?��$�e�X��E	y�����a�	��,N�<N���8\��>:KP5�g��p�<���4� ���*�@�RӉm�<c��1E�h š�&Dʀ͢��Jj�<�t.�%0P~=��#(��E"ǆ�k�<�A.�f@�cBã>��k#�MH�<�0�٬���.ܳ>���I�b�<9��1BN��$�J�T��	���U�<i�� +���6��`�cT)e�<���I�d$I�h�I���02�Uf�<Q�X�,����'�(C�� �(P~�<A�	��J�Tn��+�)�m�t�<Yh�	[����%!�~�h�Bw�<9��\�;������X'��͒R�Pr�<��"k�H��ЭV�w��i��Zi�<�����@��%���=cX����VM�<9��Y4�I	c��X�\@�q�<I"���Fqaa��8� ���Vj�<ѡ3`5�T��__7���u&`�<qg�*Z	��"i�_7��S-�^�<!Ǎ��9טqh M��4S�g�Z�<a�jJ�:�V�§H�Xj|hH�kZW�<٧c�L���*�r6�-BL�<I�j� a&)�o{�4�D�a�<�C	��h�c�� o��`ƨu�<i�� U
h�[Q�L�h#D��1C
l�<�wƗ,�P���L���j�Ai�<yg�MH���	ط=����f�<Q�eڢ7���h�D��%ǖ��%(\a�<q��{�y1�$Z�@Z�zrC�k�<q%K�2|ؤp��&}��!�c�<iЮ3E$Q�q�*E�
yh��RE�<� J�uHb"�Q�ti�:+���"O��Q6��uN{&�%�M[�"On��!T.L���#5΃vz�т�"O����9c@	����'r�pz�"OL��B�G$<���#E�vǶ�ku"O��`�a��3�$yb�J���Y"O<)�)"uHvEbG(Z�v���"O�z�˙2��c��?,�Nm3c"O�4�RO�.Z���D�Xξ��"O�%h��ϴ[5��	��ɷ�B��"O�$�Aи?J,p�m̞m�F"O`X��D��'���5+�,~�J@�c"O�h1�DҚu���%�14�H���"Op�C"�ϗT�
���f�D���� "O8�ZN5��� ��Ir�"O~�;ꙻZ/���K6��Q'"O��07⎞U$=k�ˑ�k/F�c"O�� �B�:d�p���@(��'�\�a���8�Go�?w_�uzd�ӹ~d���-(D�����QP�<�0ҕ:���7L5�I�h��{����:�	@ /)n
���M2C�I�V=���*�7<`���D�@�1u�QܓU'�>�!�&t:�#Ǿ��K¡=`����ȓ�L9�-��Fiԙs�n�U�o��D��I��'H���ĎJN��W`�]#��(�<�����<�#��4f�*���»-#jXң �`�<1`��NZL�[����blF�
F�P����ׁ ��y9�A��6ml ����!KТ���xc	������%S+�~�N��w�@��h��D�;�z���K�7��i���:C!��B�&Y#e
R."����,N�_�!�ƳHu���N�	Ǥ�*"J� (!�ÁV*�Ȳ������jjqI	�'��Qc2(Ǖ��EVe�:]��A!�';��3l�	J:.�B�QWx��B�'s��XtdJ��#���v)��'�c�AK�O���8�Ǣ's����'���`$�L�\�N�0�lƦ68",*E)�G ���I�{��H�T�6\��`��,H{,���1n�>d��3}bBM�U�T��T��9������y2i'L�*$K�B.��� �~@�!X��$!��E	P�~�e/�JG����tiIȭq
bT`V���q6��ȓL�E(�gM w�T �a�>,�$]��'��<y�E:�䫒����9O�Tx�
�R�wG����ę�02��q�E �\��� �V��D�}0t͢c)G+:���hY�bX�#V�>�x��+O~ �%��[��p��4mbH�)��3>�
�� 	u��"=9E�75.μf��[	Ri���~2�k�Nx ���V)�@I80��Q�$K����i+�H̇�Iæ��&a�]j"萦O�G�h���,�8h�����h*���%�yh/6pL��#���Id˟)_�!"�K���BB��$MR�+vɔ;)\�܃g<d��%P�b�@��1T��D�A����(oV�0ż���ϣ}���  "U�Kz)��-@8�@��L�62�3(��ez���tG�A=�L�B��0��ּi2 թ��O����Ro���q	�E�N�1R4F��1��pS�X�+��Fy"MP/B��FA�4�����*)��ɑ���AQ��e^<PdF��\�Ⱥ��� "dl �e�A��xzǧ�4��(x�.��Q	 x����CA���'��.D�(҇�|���O:�n�G�oZ=�
�CD�ڧ7�(�`�����DQ�i��H�L<��~���"�F�T��LЗ#�>橙(+plt��H�}9VЙ����?��Q��T�ǃ��4��w(D�`�bBUkr��%oX� #�3�Ȁ�+>���Q*|V�\��i2B��a�:a%F
%�~U��X�=�JiC���]t�X�4�?�'ۨn��\-6\0���dTa�\H�ф�}�F��DM��w�'���z�	[�+✂q��
(:�4�O�����J�bΨ����7�Xk�
�A�"@�F�9G��yi���6k�d<%��I<7Ɛ��֊�;qQ���	��LL���)j���7e�̟$��̅hچ6�v�,��D������r-�П�CЉ�$��@��j�)f�)Z�7O�
rAƪ�ēO���0F��+�PH��M��\��,�v�I�`1��	�k��鳕��l����=�g�? "��"�A97FҨ��O�lh�@�x���%�1O��q��;��=�|�xdk��q�vM��G��7㦘�s���F��I<=��y���|�;n�ִ���W�R'�1�3"ڻ�Px��6��h*A�\	I&������D>>I�qn��Ɲ��	dR}@
Z�aC�|X%�2;���$��j��ٓ�$����;t�5�& ��/&8Y���R
�'_��D'˥u�8��'�[-d��Y�L<ѣϔ6X�>)�N>�~*� Q.�
L���b���ʧ%�i�<��CT�P �s�
�Kj݋b+Թy=qO�M�5�<�3}roF� Fꍣ!dO�x*�Q��R�ybK��P�F7y�L�3�"�/�y���^�p�����kt����AW8�y����8ۖ�!ŌX;aMZX�G�&�y��2}�����3����ƌ��y�� n����0�5��$�a)�yRF4Rr��B��˾-H����y���t'ް93�K�=�L�p���y
S���0��"%�4���F-�y��@, C
��Y"lR� d �-�yR��.YSL�����,P�hRAmM �yB�,=�0��#�M� ��%pāٔ�y2�M24%n��k�I��]4�M)�yH�g�}a��X8�� �$���I�r�����(pF�E� �(c��8�I�9O!�D0��HJ���[Z`$c�H� `2��Ob,C��!b01�1Of��g@$8MP���gA�ȫ��')b�t��A��;v��i<�����xU�t�aR@�(�Р��bުn����e����Ox�r�^�|���;J|�"�ٴ%1y�G�n�x�#l�A�<��H�+��=�V��qn�ReMQEy�`�����G�W��S�O����a+U!M�D���ĳ#��e�ǓU�<} 2e>͎��O�gt�P�lݞjF����I�<͘(�GH
�� ~�)��NQ�3�	6~�h��@�S�~\rdHI�hv�;�ဴhPM����oѭr��K|2�m� \�����2N'��@�'�.Kx����S����"9NV}�a���/u �H�f�M���r�i�b'	1c20p�OL^e����+s.��O�Ll��0�v����b�r��c5�OT] ��&n�7�>��y��Έ=��;BF��t�$�Ӡi*�<��<���'v[��� �>᥎΃z|��ƻ%.��#�u�'��!��ʶ���Ђ�9�v�����"?�1z'�¨;tzDZ��_I���8ⓟ���C>���GB�o�h��U�	�6.��S�g�����$��/\&���Ś6^�hQ���K�d�
�&r<�:1��I����.��N�6z��h�'�
9��g[j�'��Y��J�a~~�y�K��^�]3��� �|IF�V5�0��U�P���6�:��uZ��y7o�#��D�"�N�DBZ�E!?���,�4�
�J+}J~B�]�[����#�J�>Ԍ� �f
M&�	�_�Dع5ER�n�R�!�)��܎�;��	�:S\��g�.�L�E����I��<II��@�d�z�'V;����ņ'�h�AT*Ǩq��d9u��!C��l3�ݗ-1̉`4��m�b��,�O�m���!.�b�Ѯ�F���$�	4�0��n��(1��/\H؈x�@�!-�j�!��� N��M|�Y	h���"���`i��`�''�i"�I���B��I^FF�}���_J~�]���A�t�y!���}$���D�4?<���Z�=8��'�����DZ� $،�"Lސ
@s.O�X�.K3L285�9�'u���I��O�}�,�:��I%��}�&UJ�`᧍�5g��1N�jx�Y����+)@X��F\�N3�]�5�� �Τz�R���i֟x@��8y����.;�6�]�R @�")�d˟%eAx��)�)p�챰��R��p>��ެO2�Up��^��cb%5�Fa��R�\�`�'`��)V���(��G��,��=����jR�]�P��k�>��:��Otj!�B/�h���4��#[�z�H�������:`h@�C9����ՙ?�0MY0)����E��O�(c(ʫ
��q�5���	�t�����Ʀ1��>E���"4$�K͸a��]���8]q�(RS�B B�Ĭ[F�4B�$��������.և ��,��뚭7�z��I>��6�~��� ����5�p��Q�4� �+�.m��7O+Lo�t���i�!���sp�ā>=��Å�u^�O����NK���<�H�|xb>%�,^�f4	sg�.Ahhz�'D�0����V	���l��t�*qED[��I���)�p�R��O?�I*U�vP��7Q����%~�i���� h���;ɢD���/)��P)wY��X6E�a'zAɖ�'��0�RQd����P�*��4��QTi���~:.Ł�εd��Z�h��&��d�ȓB�Y��`"+�J��D�
�50Pd�ȓd���,�?}vD��p����2��x���/u�����M�}��-D�����F�\T$�Z:sa���/9�T�a.Ĵ9ӌXwE������/fI���(;��@�D1d{���a1R�K�ñS�} t�h� �ȓ ��� "�E��M �@''H��ȓr����4Cܻj$V�j��$L�p�ȓ8��ѥ�יn��Jr���x��]��J[��5��{�2X��i�.�a�ȓ*���0n҄KM^�$��~-�Іȓ&��Cä`p�QӨ��QP����䃗��l#���G��� �� ����("E�K�vm�����k�轅�ܮK�ΎJ� � D�V�[`������
�Ké[58���H0>e�̇ȓ��!�
�%`�i���&w�ܩ��*�`���*K�@�8��# I�6�z(��V]��¥�׵z�@��GְM�N���>ނ��o��I�G�)_-$��4D��r�� ���؄�ߊ�<`�'?D�غ�	S�j�!M��8�d�9D�|	rnU�Z�x0��n���1��7D�`(��'O�}�J%,qp�4D�,��!S�w2����'�,�BQ�7D���b��B�
Ѯ�#��B�2D���Ɛ�v���CH
s�́�f,$D�0�����l떼���r�X �.D�$Z��]�'~�4Yrᏽ�z�8S�8D�,��T:��Eq��Lz�:� '#2D�`He�B8tL`]`d�
;p�xp-0D����\��� ���Nx��@��*D�X���ߙQ/& ���2}d��'�$D���d�1	�cFM��d~�}SC#D�d"�G��\h��iQ�W�\<�f�#D�l�1Nɛ�8Dh0�O3"�
$�'!D����푕m��@��C&���;�!D��)��I ��B%@�;w�5�A?D������U4�Ņ�Z2�I��<D�$c0�X /Ц��.ņ5ԞY�Q,8D�|��J_���*׫��Z�`7D�"�×''�4u&ث"t��"��2D�lcB�D���������s�3D�T�@���i�	P�N�&	�3�1D���G�H�c��Gj�PI4�A�-D��ҳ��I�,Y�g$
���[%'D��a�d	�^+��R�&y�C��6D��IL0H$~ �t����a�$4D�|��FC6Br�i�c��6X(���ti8D�����ψ�D�"m�,9S�9�3�:D���0I�ny�Ú�K4��c�9D�p�4LN�(�:����_�o��pR!C6D��;s@\�=��QEʖٶă�+D�ܙ�
Q l����O�^�cf4D�P�t�Z@;��E^�#��)6D�Dȅ�K�qW����0��x��4D�ı2�v��9�b!S��p�&3D�$*d/�$D �%-$�� �1D�L�匈hT���K��P�h,D��z��.!FL�F��5f�x�!D�� &���ǆjS �˶��<�n�  "Ob��u�Z �L���?�6	�R"OX���aZ2vn��Sn�@Ű`q�"O
�!Q[�l_�t�Ƌ�ȔP��"O�XP�_�i�%#�EW��ya�"Ol�ѫd�@-p��ϙY�0���"OB\[�O䬐խ1k�ҩ��"O�R <{ذxYt�A���U"O����/�"(Cd��a�G<I"�1CU"Od�C�I�F�H��B(Y�ƍ��'D�×m�<>� ��LS�F��Db%D�(�֫���X�82"L+k9�3E$D�4��*�*Ar(;#�K ���k�O?D�0����[To��3�b�J�#/D��_{ 8��D��<��-D�,r�KY34��ʣ#
��͙��<D�h�0�B�BO𤫖��2V�~� G;D��p^�`P�"�퍼8tQg9D�0{��;X�v�Iq�I�xѳ�7D�xB�AуP�L��U�D&} ���#6D���Ԩ۱�����c��Dh�Ӈ6D��Ӥ��eF�PX�}�&�ʗ!��)y��h
�"��!(�!nB�!��{�pR�L�M�X� .J*s�!�F�w���=4��i�C팈"!�V#:4HQ�[��T�U��4[!�D\�)����M_���e��h!�	�sX��2��ǻ#H�]�ЌN!��]��.��+
 4JQ��F�g�!���3ld8Ec֯]2V=d�ZTk�0�!�0z�8 W�ǀ(%z�E��<H�!�DO�4Z���e'����Y%IS};!��ƪ>��R�K�2k(H��Ñ#I!�@aL@ �D� �z���P!�\#����\�d��ٛw�!�J�B�8�"�O�HOޭ �k�!�$T�$�9�!�J3s60R�MU�_�!�D��:�n�a��44<AA�N�+V�!򄚟4�Ј�V�M7�ˁ�,c�!���;^P9v�<XH���4:
!�$";<��}�Eb$0$Oz�(\�	f�BD��3����/��͒�*ѬуV:BP��,V:=Ȫ��I�u��8q�l��>^��
� \
B,� �dn+�!��1�Ɖ��F>9�l��ǔ� �d��6���K�6?���H?�#��+ox�*���ݰyc@9+�!�?/�B�	2%�t��σ��C ���qBc�	g��HQʁ����`�'Ur��'���"#���y'�_5�������&$�����>��K�M��MAĄ/��!�ªR(p�E�%U�|IZ���n#��D�V��9Q!��p�Q� �S��+���yp%��,ި���<���iw�LQ������mV��?�n�e�@9_S�ICvC_:".�)��-֒_���e���0>8uC2� ��W)z�T�8��E. �|�cGd6Eh��ԍv�P��ޟd�q�'���hŮ��k��4j��MCd% �	��-Ar��q�<�Ԉ�x�}�Q�2 �Fh���M+N��I9��Z���S�[��%�^?!�DW
+���9�w�e��m(?��90�'����P��!𝃃�׺@,uyRƝ��� �F��~��	Qw��6-@&<���I#&�ъ2�85<�i�BF-v��a��U�H�*@��(O�"䎇.p��1E S�`�@j�?�k��D>�-��h"wϾ��gթt���D���4bߓ[p�Eq�*�<%�%�f(��.и%����皳m�v�P��Yr�I�?aԻi� Ĩ��Z}q����Kaj8�%:n����at��xQș�(��4%%�6;[�@������RnO�WQPi�s%g~��hq8O�[E�շ9]�,̻g���<WUru�,9�|���v���˥"لFq�De;^;�k!g�$�z�+&a��UZ ���4�?���z�*�v�
�u�|�?A���E0d�1�L��q��@~�'[�1J�%�#3�qC� �<u�'7Z�� ����ͦ(�ű2�]�@u��0p�84�L�"�Q(w���DT�K
������D�3F���y��X?Z�H���8bV�Q��ן��:�⅁g(��2�=����8_ b�"RD+X4���`���yҏ�?�>�i��)i	�9��J���Q��!�fZ���1��>t�	��k�n	@@�H�[4�C�ɭ<G0�9𩂺 �"@q�@D�����#D���	�%v����|bOh�h9!���q�l��Sm �Px����uѮ퉀M	�O`� ��#�X���[�ޜ؇��)\��h1�Sa���!xD��E�M'�����ܰ���S6t&`+L����5����X�!�d�$2��� E�E2�6�p�)�6FƉ'�}���S?l�ɧ�O�h��`
UF�����:&�
�'�5;����>��t����9���0B�0`�z��OV��@gQ#ڑ�Q@Q�~^�{6"O�{���qb �Q�σud��ʳ"O���f%�L�����<[t�R0"O�$Zb�Ԏ����0g�+W(�3�"O�M��؃]:V ���� �d ,�y���7J�"��D%�U,ҽ0�͛�y��Ȯ\k2��!B�._s��h���y���e[��J�Y��飇D�y��M
'9ؤkAi@D��(��ʫ�yR���F�d̜L�4�����yR�]>	�����8ARȊ���<�y�[�5��,{0�^<k4ʙ���I�yr'�+M9��y�Oזcj�c#ȵ�y�ON;-��ԡ���]�~ Qb�
��I3���P���	(|�� G�5c�t��Ƥ�4R�!�+HSȀ��Ww�re�X)=�r�O�R5"(?�1�1O H�p'�S
1Hw�5,�}�s�'\� g�<C,Jv	
�L�PDȮT���Sa��`؟l��#	�Xe��S��>I��)ؗ�/��%<n�!��OE� ��U�3�'(���`��U�"{����"O�d��l�Zm�!	%Ʋ�V\��C��C�(��֓>E�dD��v����eN0ލ�g�nX���ի3h�O�x����	2��� �� Q��!���&��;=���Vl�3�3X($�Ck�l)��`7�I�N`,�"�\�Ñ�JM��PF�Di�-���M܇U]�*��Ύ	O������o��u���(k�줋��Q�]���!�� 1@�↨.?q3׋e����vWD��451�;'��HT��-Z-�0�VJ��Y��i#��0D�Y![M,����Y�V���r�Xoߌ=�%���Su��!(U��'>>}���)(�ǐ<jȲ4���6���H$n��D��=�ʟZ��tM�m?�yJsh� ji��%�DI"o}����d��j�̄�SOwC-"��*Y�F˓{�p<3tY�-�j�
���ɵE�Ȕ���@$�{�F_/ܶi��̩��O
�P� ]�Fi�O@a(���`��[���Nh9�2�T���$��E��4� ��
4n���Pw�E�y�^8���$k�I�!�� �K�H��S��*׬!c�Qu�)�g,נr�N�Ѣ�ʿ6�^L8u�'�<:Rm���-@#âێ*�*)RM@#��l=�T�Ԩ�D+��O�n�ƨ�N���$�yo�8rWΒ�&\`	iB�Y�����$�"8~+��@k�C9H��!C�2uG�A���Qg�&��'>I pe�:�>����¸�v4�a�*��\�n����� �ɟ8�A�l�*3�nԑ� ��!��#�$
�#�+1���JMж�3W�^�㒌Pʕ|^��-y��3�;-P�qE�D�4M!ФmCud)UF�:,�$��4�@<�JنE�~P
c��xUj)K �1+��e�'V�I�e� ���ϸ'�~���+Q��2��˱bX��X��t�r�H�E�t,��i�ҦaإpW N�vQ �G�L��0?a�F˿9��[A'�seIk��NO�'���2��	4�?	rD��VH����V�Ze��E>D�@QÉq<�����͚h��5�6�??��a�7��K�M&}��i�*DX��D�	��T����Ub�!�D�6y}��"���1�샧M< h'�蓇�>q��'�l�eΞ�ư���
.^R*�X	��� �<`�*LO�n�xU+�?r����"O�	"�h�T�h�0IT4��k�"O4<9�n�'�ФE�:��e"O"�`�3�Ȉ�s�Խ-^r=��y��w�H])G��&�N�A���3�yr��9W`��<�����Fِ�y�U�>NP��Cڑ	`f�1���y���&L��� 
Z�{�p-X�$2�y�)�q�-@d	'q�<�!k��y��8іL��ʬj�j�� ���Py�l��`��eívFe����[�<���hYp��Q��.jpt����_�<QRC��e�"ɒ&%ϨaRD�j�#RX�<��jڲ(}Z�)�_/D0�*4��@�<�ï�+%�\|рO����-k�Vp�ȓ!^\��wa�o�`�0+¯i��y��{D�*���3r�9p5JR!	*��ȓ@��-���F0�Ha�c�:�v���b �� g��I��\�f�K=rM e�ȓ&@$�VN�;F��p"A�]�U�ȓ#|�Hr� ����P�+�\y�)�ȓ��X�#W?!���ĆC%c܅�ȓVLx��'d?���%W�4�\���%֜��%�F�}�X ��Z��: �ȓq6X豄���;��r�.�U�zQ�ȓn(@�)�|�CW��!�� ��o@��8E��/tyX��|�����\���`U��IՀ!��B�t^ZL�ȓc��Q:e���$�������C�I�p�d(���vÂ8 �ɐZ�lB�I�D����Qb��L�H��$���9 C�ɵcʴC5
2?~< ��X�M]�B�	,F3��Q͍!#L�� ^C�G��	3Ռ˶j�M���5��B�	;���0p����0�
C�i�HB�I_������[����*ߑr�C�I($!H0��"7ӄxtΜ3�C䉹w���"�O��J(X�-�~C�� p/�1
���p��5�
�qHC�ɛ����f-w~�Ń&�ǰb�&����2@��� ��OFz�ceHݍvq>��!B�t-!�d[�:tЅ�T �oz�p;��Ɣt!�����dQg�bvH!��j_�^!��/! p@
�HQ-`jx��(�q�!�K�Xo�Y�ؚmhr�[Շ�=�!�$��DŴ a�&�GV���GGÙQ�!�D��x�a�!��#S�0��7�H�/!�(\��-�-�� ۣ(J:?%!�$�x�&p30-Sz^E�ΗK~!�$������U�e��VH�G�a{��!�;y��1��# �qJ�>+"��ɉ�P��Sl# ��-�"t�����K��5R���&"��ذ㞢2��.P�uPFjد�Q�b�ߟ����=9��/��U8��%dnh<1�A	"��������b>eq�J7j7�<05���QJ*}rJ��,���=�g�I�7�!��%IZ��8�.�z��I��,M�?E��dWbF�南�^�T��f��jIt�80F$�)��M	��K䩋<6��a�I�u���҄��6��O���'o9� @�,�v���TH�]e�=o���'B{B�"��h�p֝�(丄A���\�P�!�S8/��݂R���U��)՛�?�B	8�l��!ɬ/(�;W	B:.��A1�ƫ8�����<�bh���a������Դ���� D$l��c��6x�=p��O%*qǞ������'G� �Ò'�)����d&U��x�<�N�d�L�':2����O�"��i!N�Ь �����̬�ڴC�<i*�)]�4ҧȟ� ���a��O��a���}D�`w�ٝLD��'�J���s�p�B����w���r�'� �b��0h*H�P�`Y�`f��`�'+�lI�*Z�k��p�lZ$�qC�'�!�	:8�a�J��,��'>&刕*�3:X!s�ώ�%`(i�'�N�R�'E�D���8�ե�h�!�'��!K��W\*J�x�c��| ��'�0���W�����A|J�`[�'J<ꃏ�4��!�&,ɍt{(x��'�����gL�j�t�Pa�>MZ���'
���E�0K���gHח;�@��	�'9>[$�!�z,��hߏ0d�@	�'�28���'aK.�k ��Tu�9
�'!�h��Rk�0`0ϝ=E���	�'�\�:P�*�<�����l)�\��'D���ց�Mk��0�R�1˰x��'�|hb�o5��� � v�Ј��'�~�{'�q �@�cK1D���	�'��S�hA�-�"E���3>Ǽ���'�j�r�"���\�4�ې4m$y;�'��(�� I3z~����h̜{bN	��'�^1��@���>� ��ȏoM�,��'͢�� 	]������C��m���'��ĚQ�ӷD�LШ��'���'_<Y����A�p��A+C/@��'��l�7Dޞ�\�Sѣ^7/ҭ��']t�O�$M�|ʑ̄!�b���'�V�Z'�4u��q`%��rTr	�'�4��?LN�uY���^8�
�'k:�	&����uc׮�r��(	�'d��t�]
S8@3wF��5�n8h�'���tK�=f���Ӿ&�`���'6J��&��C�Б{����*��[�'~Ő�i�<���Ҕ�ܼӸ�Z�'+�٫`�ih�ys��:V�ȓ}��;W��L��E�#�E>�T���m�|8a���
�>�(����챇ȓ.����u)�E�Z<�rLZ2V)���Jm$�˧�	?�|y �Էz���ȓ<n6�Q�&�q��x r��6���ȓ
��X��DeS�]���T0!�����&� O_������+�ܥ��]�4@���6N.t�P��%zl��@�Hp��	 Lb�sd�E�w� ��(`�hBW��X�p%�b�إPx�U�ȓd���[ЁՄO��MSŅ�f ���8�\�����J�[pC�: �х�3�j5Q@�0jj�z1/]�k_&t�ȓfK��h�)I�|�
���.[�xЄȓ(ZF�2��KrмR"��6���~����h�{i�z�L��Ψ�ȓV{<���(,ty�q �ȓT`b��\���#`n�=Z��U��e�B\q�� �Z�ⱦ�5h+���ȓ{�Ʊ���f;�@�� 
��ȓc0$m�[Z<^�[�M�h�@��8��k���10�v)�w�� m�X�ȓ_���O�4��4GԒC��ȓ�z��PI<Q�t���p�ȓ*�m�鏲o���B���K�Pu�ȓIݼ��cl��Oe&aQ�Pr���ȓ0\�� @�Јdf�0�VΒ\xԆȓq)>)� �V<j�L)��(�5?h8��S�? �9�T�j�L�6�\t�:"O�	hޖ#��$95�9�Qq"O��(ek��3��@qmGf���"OL,B`C��l��$j�-��l��|1!"O"�!�(F�(/��xЁ�aۄ}��"O����DJ�THF�G1��]`"OԐjf�Y7:6j��g�g�и�"O`}���#��kUǈ,�\�#�"O�h�KܹD-������9~��T�"O��1R$�!_K ��"1��"O&=+L����d{bVb�,	�"O���완!'�y�#��%-(Juj�"OV�8�� O�x�H�@1W�|s%"O�x�%�&���I4��-E(R�d"Oj�8f.�(�VM�Y���3"O��X�L�1V�ք2�	ul.�"O�� 0�X�\�}RP'�����N�!�dA�~�1�I�c�|��u�E�X�!��4'P�9�ʜ�J�{�E_*Y!�D�������-��hjB.!���/�t�Brk�R �9'���FN!�$����áF���l�,۬a�!�Q9��U[d!C#�V�Q�=�!�DO�zC���FX�"2����D &B�!�DX�:�rl1�� ".(Z'iU�*�!��ӷ^/��K��3"
� �7r�!��{�� ���$ �����p�!�D��o�=��Ef')�f��O!�N
J�jTҷ��(ƀ1���&d3!�d]�
�%�w��((�sfeݼ]�!�DШ(�2�v�4	�!8F���"�!�đ9e�@���/bɺ�h@��!�$���P$P�g�f�*a�F�?5b!�ҡ.8pԺ�l�R����p��gF!�D�+�zٸ���:&��d `A-+!���EI�u7DN#��i�O",!�$� Rl� K�|w���
Y�K!���3����ǼcH�w��2�!��J��s楉,~oD�G)��f�!��*ArnXSpc�5~^��e\d!���="�����ޖ
�h� &I-oG!��ƚQ�}�$@��d�$� �P��ȓH�NM�rH= �
�F�ĂQ'�A��{8����m:=\���b� �tć�D9��4�G����=Ay�d��P����OE�51� RN'H �ȓ>�^��p+�'Y�!� ��"j�9�ȓ㺭�`,��b4���P�I�ح��=��I�NDa�yä��	HX=���42$_6#��@�� ��(�ȓQ��ċϖD�
4H!O۸Q�2��\!0�ɅO|��3A�ϝ!w��ȓ�Ɛ2��#鞜;g�E�2��0�ȓe>�UcuHA]���sҗ'�DЅȓ7ꔜ��	�dI�1���͐�lD�ȓwc2�����-){��D�<�X<�ȓ9��S1��V	���6L�VZ�	��,�����!XH��"/�:�6ȅȓ~]T����B�0cj� ����Nk�8��KP�2�V!k�ʚ3^���ȓS��9��M1$6b@�b��H}�H��o.^�8�I,]��s�&�����ȓ_��ӈ_�`��rV��P�t��+`P�ۦi�%d$��r��W�A'�Q��S�? ���N��6`��C��9]O��[�"O��: %��,�?Zq	V"O*uB)�#cy`P�ci���ӗ"OJ�ҷ��+���c��8���"O�v//R6��'Ƚ�� �"Ob���D]	Ն�!'L�^vLI#"OJ��%E�2+@1.�+����y*7����ŏ%���y�͘��y�#[2i)7K��R4r�*�(ɚ�y�v�(Q!V�^	?h�3�gƛ�yZ��	�BA13��rC���)
�'���d�8X�
��g�B�4�H�j	�'H`ěT�A�N�,@�7���,��'��|2p�C���H`��( �)��'�`�{��~f�A�ϸ O�y�'yT�k(����0P�f������'���q�U�6T0�@�{=�,A�'PL ���>hX��v�������'��T�Є�Z���;��C2QxHq
�'�-��i���}"��ǈ~!P0	�'F������Bl��#�?rԵ��'.����#r�E'2s�a(
�'�^���n�?"����$%$0S�'��%��E^����B	��'���C�Z���UO^���c	�'B~�)j�V:`{��P;�x��'l���W�!RPkO6G���'����(�<q��� ��QHL��'�&�b�%\�x�*�it�x	�'2R X�J@'�h0AB�:{�h��'����ga��s���x���#yM±��'��02���qc�	X���?T�'(<ЁgØ$�x�@��n��#�'i�����-�!��J�5D�X�Qbϗc��Q��2W�pa�4D���׃̓���g"��P��e�0D�)W/V�H��1��O6j�[@d/D��A'M���lb(O%a��i���/D��'T�q��yH����i�-D������t�쀑 �'i���6�7D�T����y��+1aZ\ИSr 5D���a�So4q��WD����*4D�H�d�X�Z�<��%,T(��	�dG$D����#	��X�0��.,�`#$D��B%h�P��L�$ʷ�!D���9_�Z�Pd��<Tu�m2�� D��k��.D~A�Bn�8�c9D�Q��� ���s�Ю`5�ZA�*D�x1F�>"�Y[Q`�	-8d��";D� �$�ͺYC*�蔧��ỳ.D��z�ȁ$fhD�A�c|�F�7D�\�������勝Y���3��5D�A0�D�9�"(+@�E(hf��`C�3D�@Z��Z"?�d����?afYY��-D�$��d�.I����4:�Har��,D��8��V첀�`��u��p�w�?D�Ȉ�Q�T����nJ� �wI3D����O���z�� ;���Ң�$D��9���[s�ÕOT"<�l��#c6D�T���Z�U��
�E��N.���7D�,¤��
"sl@�`�S�S��*:D�(B���7�Zhh¥,/���@/9D��� f4aJ�ӕa�z�ڑiB�6D�`륦ռ�6��m^�3U�9є3D�� ZX�A$Z�TA�!Ş"�^��"Obu��`�+3n���	�=/�|�*�"O�)����&��4��fR�\Pm�"OL�aF�[_�(5�@ ��V�\�"O���3�߷-���R"�E�b����"O�D�    ��   �  c  
  a  U+  �6  �B  �M  �Y  Je  �p  �{  ��  ��  5�  6�  ۧ  %�  ��  ��  8�  ��  �  ��  #�  w�  ��  �  R�  ��  �    � � $ 4" , [3 F:  C �I QQ �W �] �b  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z��Yb�с�5|O�"EG�;֊�R"�O�~Q:�F�'VP���Œ�'蠢DO�	J厈���4D��@Q�Ђ:�|@��Tfs���(D��`D�J�=Np�A��׭7����Q,%D��z�oV5H�r��.Q�����$D��p�L���Uk��B�����F"D����`���2����{�& �E�<D��PL��j���H�G��:f;$��S���T����t��n�����^�D��� �F��9^	�F�=[`�͆�Im�)H''��*-���t�S:E��ن�	�H���
�e�pڶ�3<K�̆�;�؄�c��v�`����֭wXވ���t~� �6XvD�e �8�HP��E��y�D�9;�px����|	J�fƈ�HO����"��aA'ݥtǽ�!:w*7�!�p��`�:�4E�*ɠ����Gu��E{���\�B��8�d
5s�.,�(�8zE!�$ǈ`VaR�킍wz�q2T�
�-!��QI�V}z�f=n�����,a~�V���J^X+ָ{�儏v(p�R��5D��)��?1� Zg#��o�2���(D�p���%HА�(��� ��Ȁ�"lO4➼�eO\;xz\���%$��1
!D�p
`f	 CHA�0���-ƵH%�<D�pZ��CX��wf �B4F<D�<��"J!���#����.�aDO-D�qU"Ո0<�i3K��$��X��0D�� @��#aǵu0�IՊ[�zl�s�Of�'�6�NQ���I�k0L�F�_3��݃�!X8Xaa}��i�d	x�Ա$o��\�j�� ��Vhm&H�(#<E��4'u��D��* a�<x��S�RU���Ms�B��D��<3�Z�V��#YRy��,�OҜh�k��Z�:i��m�N[S�'����O�4�V� �ń���/( H�"O:mKw����b�GF	ڷ"O$��$L�GE��;A��t�V"O�p�##�&6yK83�� ��ݬ�~��'�̀�=E��' �R�yB&Ӽ!s�$�DH�:�y�DކE����B�
}x�^��'J�{�A�^]~|ӄԅ<(��B'	I�yb�����1q�E�-����ȗ.|�B≎;삔t�+I'�h[���8E��B� :��)2��a�,���	�3HԮB�	�s@�@���d�j����P�B�	Z�
�"�7d|�b�KD]�B�ɝIhZ�q����*�y�JO�jC�I�ynD4�7@ɫ	�8��B->0�>��}b�f�qiA�'-P�i&�G�C�z���DI^�<�sh�E$4���(�D7�)Z`?1�]��m�|yr�S�\Ӥ�#��J>�+"
E�V��C�I7B�F�v/��q̚���2j��tE{J?�����3>k-���I���A(6D��u@I(S"���n�#^�u#S�y���>9��'��	�E�l���4�\#�4����'|��R��-Mu��;�!a*�e��'��D��EY�3�F�4���Q'��+��D �S��퇺V�N�ر�	�<y�0��+Z�yAP2ez�=Hb��##�А
��~�ў"~�Tӂ���`�[�$��iD�Rԭ��a�$��΅�U)�%a��.P�l��\�.��hǾ �8:�a_� �����B̓'@�1�F�z�BQ�M����ȓVN^��ؽ���Qp§ ���n� �EE�0��Qtn
&V��_�<�ەi�#G�L�f�I� 	�ȓ=�r!f�,`� �2�1�t��=fPH�bd�3!��,�
!H����l����JƑ@��\��OC�f�4 �� ��Q���
� ����[�����-��l@�m�!_~����$��2M�ȓ^`�ђ �8z�Qb�1n�Z���.�C���J�~4aC.$@�ȓp�D�z��

�V1�S)־�ȓM��%L��	B�� �
S"���|/���%�3-Yt��N׋]�����.�ѕ�Q�F&~���̈,M�]��t�����^�U�FӅ.��S2���i�{�J���?N䉇�����fE�,Mq�(�,D��Ѕȓ	� �� ɠ�:��Ơ��j��-�ȓjJ&]!g�B�x���blV�k��U�ȓ{R"q�N�!r$0QR�&z�}��T��a��W(x�]���"^���(�ڢFC=�8@��j�g�pQ��G�"�BG"f��lљr�4�ȓ�M�P/W>o���x5�ŕ"��
�''�#r?B��K���a���
�'\�P��mɀ)%�;���
�'�����X�v\�[4	=oH`	�'�����U(���i˺	0����'4Z��[1����p �YL����� E�����Y0�)�J�iw�!q"O�q�ʇ�gs܁�˓�*I!�"O�Y�6���I	@�R�`M�"O���# R	
R��0K�B���t"O:�!ck�a��L`Æ�'��xi��'��'&B�'�R�'r2�'��'u��W)��C�5@��J�L��'��'*��'���'�r�'���'���L�1d���XC��qՊH���'���'���':��'�"�'p��']�e���nA(\�ƪ�u��Y��'�"�'���'|R�'���'��'�����M�	`���r��k��y:E�'��'j��'���''��'��'h���@0
����V�V)qJ ��']R�'���'m��'rr�'z��'MD� �^9D��8R/�)'M���g�'4B�'�B�'|b�'"�'���'Q�����Eg�j��4@�(��4�'���'���'u��'$��'���'�ژ��-���J�_���ze�'��'���'M��'J��'��'�\];���u�eナ�'-����c�'u"�'�B�'/B�'�r�'�2�'��+I��``I ��7Ȱ5�#�'}��'��'��':b�'R�'�ʱSA��,ol`�2oH�=�����'�'�r�'Y��'zr�'�B�'�J�-9	⬱B�W&S���A��'�B�'�'K�'���w�
���O��[�G���"�|�2�:��ay��'~�)�3?A��i�BU�e���Z0d8!`%֘ Bh��������?��<A�M�	S^`aCN�#s�RI ��/�?��:u�\��4��dz>���'���5!]ZA�0��~���mS�`bc���	ly�
ff�ZF��Jo����&44,�ߴ>�*e�<I���'i����!T�(�+6��q�'�4s�n���Ox�g}���M��3W�V<O
P��dٳ2w6�a ��>
t�-�5O�牛�?�@':��|"�Ql�,°a��A���Bq� 5t0͓��$%��F˦M���7�I�(��9��������ߦP����?�X�������������glJ�
0�H\�Ũ'ʗ"h���l���^"#Exb>m���'Dx��	�Lxf��+P�N��dr�h\�$�Jt�'L�	��"~Γ��Gf��F.�9��f?i:�ϓjR��偫��$�ϦQ�?ͧL�|hh��v��$��hb�FAϓ�?i���?ib+���Ms�OB��+���L�f��:�=R�Uj�dKFUO���|z���?���?����t�'��)O�X���g ��(Ob�o�t�,�	������?}$?岁	G#��`d��]iH���KĖ���C���ݴ:������O;�$/C�Ty�����Ս@�`Ԡ�ݗ|\�h �ih�˓2�u 󊦟�&���'�]���ȈW���c��:��8�'���'�"���\���41
<��_P��n��m��Qt�!+=��������x}��p����IԦ�"Ջ�9؜sW�Lu�Ը��L&�oN~r㊍3�N���6��O�fT�E:<�$�N3�N]�����y�'�b�'��'V"�i\�j�0���I;t�:��b����O��d�즵`�gl>��I+�M�����6�3Q�\0j�.�n�:WN�$�� ڴz뛦�O�Θ��i��d�OB�w���V�`��$�[8��$��lP�`h>LH�'��'�	����t�	�]�D��P�f
!���<I��	ȟ��'�6-t#H�D�O����|���}*dt:u��'eP$`t.~~RĮ>ac�i��6-�J�)Rт	����kb�]�g��,#To�-<a/�?�MqX��xm��9�D�&6"q���39��°		9.���O
���O���ɷ<���ij���lѧ�r�˱��?��Hq!
.,�b�'�7M1�����$v�~��'-�Q����Ty�T�@����ܴ<,D8޴���H'D�U��O/�	�R�>���LD6I�бʗ�M��	Oy��'B�'}��'|bW>���h�=0�j��-j�~��o���M�kM��?����?1K~���w$�Ҥ	Ͽ5�`R�H?��<YFfoӴ�mڳ��S�''���ش�yR��7�!be+6Np��p���ybA�V�@q�����d�O��әBIL����i�������)K����O�$ca �O��m؛��?|��'��*
>?�J��>dд���ٯ��S�������ē��9k�4�?�)O���F�GuhB�f��,v~ũ�:O��D�&?h�0���LF����?�y��'��9���v���kD�)��Q��6Z�8�	����	ݟ\��J�O���<Ab�41f���i�w�����$l�I�c�<���iM�O��3BS,�����a:��3�N�&5�dxӔ m���MK�`ͅ�M;�'%�wk4��'-oj��BՏir��H�ќt�NԛH>i/O$�d�O �$�OT���O��$_�NB��!L@��t;dϲ<q �iA�M1K����'*��֟���'���e��N�Z��'c�@D�i��>Q��i��6��Oܝ&>��Sߟ�PcŅ�l,���B�zv�IR.Z�<Ϝ4�V ?y�d�z��������dV3oU�HH�`�	x�ܩ:LT��$�$�OPa{��G>�4������q�;k�Ԍ���4�d���D	�0pG)�!'`�Q�9A���X}��'���}��2�iϜw�v���.� �81G�Z,8�P7�u�h�	3�a 5֟���*�{�? ���gcD6I�HHI�I�*!�F7OD�$�O��d�O����OZ���$'�n��D�%-�(�x�M |m,�u��Oj��Ʀ�@B�MBy�'��'k�TF�U���Ր2���B�a���7��6�q��	M{(,6�}�$x�fK�0���ô"�x�&��&B!���)M�M�0T��N��h�Kj��?9��?���t�}��ÍEO�����A��q���?)-OX�n�%�<5��蟸�I�?���-$p�1���a{5��62�����D�'aҴi�D6*�S7Z^�@��Ɋg��4�CDN�;��`���Մd��y�&?�f��h(#0�m��`��?ͻ��ו�-Z@OC$|��x�&��Ɵ����8�I͟L{� p>-�	iy�p�]x�o2>�,�qT�I]����h��t�ܟ�����\�������[��a�f� ���-�b�EIXw2li�`m�Ϧmsܴ6I2D;�4��ě�&�&� ����SR�h8B�cY���Fȁ-iLz=)�4����O���O|�D�O����|ڠ�ܲ��圳M>I�sh��9�X��ݴW��e`!O��?Q��2U��?�'�?�;.	4������sw��	F��(�:aⰰi�26]ݦ����O�`�v�i���}��2Um@�EP�$�v�����,X�H�h�d�Z�c��R���۟��wC:x���,��.�qA����|��럄�I]y�x���d�O����O�p���:����-@�K^��f�O�˓�?��O��$h�lody��Ee�(Q��5��y"�����j���� G�F_����u�FM��P���'^�\��I�,�\],B��D�tg˝�?���?����?�����'\2�ޱc~���"H�#����@�+CREz�� �g��O���O���<��Cs�Jw j�y2BU	To���aT?ٴ �v�mӪ}�d����ӟ�j����Ĥ�nzd8�Յ�Npt���bJ�r�\$�'9<7�<ͧ�?���?���?yW"Q(�u�Ҋ�|��\i�m�����榡��ʃ���̟|�OB�'���CDX�A����!��)�1@X�X�4	w���~�
����	�B����T����Kw��j'�tSAaA��u�@��\�ƣ-2R��Py��{�P�1q�Q�K�;r���`,Ǖ9=�H���?i���?�$�VA�6�)(O4�o�:f���S�J"�"q�߻#�6�a$@M�:|�ɽ�M[����O`��'���i#.7m�	���fY�=��[G��#5E� q��r�t���$xćH����-?���n'֍Z�LNbi~%t��l@�D�O����O���O��+��H7�LI+bOF&<��geahj|	E�H����Or�l�j�'���'=�	�8[��*	U���h&�@ `� <�۴��$|�!Dx��R�6m"?)���:�����ag�`Dj�?��m���O�q.OT�n�Uyʟ���A�3�g2�!�B��"<Y2�i��Q���'v��'m�2Q����D!��At��<���G��̟(�I���S�D@��u��,ФE=
gIG�Z�lG)����<ͧk8��	O�	(��%�V��=hv�iѕ��q*N�������ß��)�SGy��c���1�πF+���WKR�b}��"������O� nZt��L���Ŧ1�!d�!u������C���"��?YߴI��t��4���к�����$v�˓l�,hs J�mi,�y��g�P�͓����O��d�Oj��O����|�q����`)Z�(Ҟ_U�h!!��a��䐧E���'/ғ��'�7=�8<B��M1K�P)�� E�m�ń��=!�����|�����5�Ɍ�MØ'2�LS�1��`�㚘z�Y�'���J�˟��1�|�Z����ß<qKS�t��	!F��L�:���NX�� �	ԟ���^y��{���Rf�O����O����P�?BP��%�/�X�>�I ���O���1�d�hb؝��-��M��a㎛ a���O.�Z��+(�&	@Vj�<���O���DX)�?�4�67��2�"�4/���C�/ɟ�?���?i��?Q��I�O���#X�$F��b��d˗��Ot4lڥ\�����ܟ� �4���y���x����ABJ�,
V<{5���~��i?�6m�ʦ��p �榑��?A��ޫLD��)	<
쀡�t��'
����R#$p���J>�.O����O|�d�O��$�O���BO�r���:��]�tw:�Iϼ<��i�ɲ��'�2�'t��yR$w���GF�¤������(��Fl�F�&���?����6}d��.��v	��D�	;��b��H��59(O�HH�W+�~�|�[���q��3`,��'��cC∫�ƚ�4�	����I��Siy,~�zةq��O��%l@�$d:�+N1�Q2T��O�Ql�F�5����M�Q�i�7��=�] �%ڪ$Gة �G�a�B��q��"$J5�?e&?��]91@Z�jr��
�]g((X�9O"���O��$�O����OL�?�fG߆|��+7�� YVџT���@��4<$Χ�?��iS�'��pf�0�`4�dC�1*d��.��Ʀݚٴ���NB��M{�'�b�N47�Y�����pȬ[3,ڣ��5M�T?�I>�.Op���O\���O)�GV��L�@lD�\�eJ�O*���<�i��*�'	��'�Sy��j!E��|��`�7� ���	)�M�5�i�XO���$2˔?_qR��W&�f�x��H�H��eF�o�b�'C�d�q?AN>9��t}���e�m\`	���`<A��i�l���k7%k �1�a�>IV���J=���'��7(�I���d�O��� ̝4h<!c&���BA��O��m����m�w~�N4��%����� �Z�H�SsRl�@��h �(9O�ʓ�?Y���?Q���?��򉃳t�JH+%�7"@%�q�L(�f�oZ��f�'j���ܦ�ݛX�N�SQh�1����E	ן+L=�	Ɵ�K<ͧ�?��'�>aK�4�ykT�$T(�X��%��	�����yb��ue�l������O��D�^�ʹ�RE
��r<���%hn2�$�O����Oj�C؛�hq�Iş8�ֆ�0/.t�RR�//\حhDO�'�$c�O���O|}%��Z�LL9s	BY0�Q�N
a�e�������jBwQR��<��'_nJ�I��b�
0Pj�K3�ϛN'n��A� ß<�����I��PE�T�'�0a�&��W�H��I�0f�|��'�7ٺt6�����4� ����A��I��	��U�77O����O��l��A�~ o�g~Ҥ��u���'`�	!cJ<)��	)�KN4��TIL>!-O���O����O,�d�O�!�ǋ.c<A�T�Aú�Rb��<�e�i@�X��'��'��:��C��):�q���p�4�82��B}��'6��&�󩘖b�qs�B�f_Z�:��č_�����v�z`�'%n�S��_l?�H>�*O����%[z@Q���	N�.�:`m�O`�$�O����O�ɱ<'�i��p���'�!�L3C�5�%�
C[|�W�'��6�(�	���DP����4�6�	g
U
�d� E����S���o?&�ZѳiU�D�OX���MS���tP���S��	��L�O����C��N��y���I��	����p��W��,`2�AB�ǙGO�`�E���$�OJ�m��I)\��֟�*�4��l��y�C@��aj�m!e@�R�&��V�xB�`�ʽnz>H! �=�'݈���]8� �YƍE3?�I3b�S0�ҥ�������OZ�D�O��DT"��Tif�ށ@��4�U�Rl���O�˓A��fL�d{�'��Z>�X�N�Y�9�Ck	j�!5�"?)eX��+�4Tꛖ�$�4�l�I�-�<A��2�VɁ��>}1<�A䎞�z(r7��xy��O�����[I�	Z��ހ.��[S+C�n9+��?!(OB��<���i��t��ʊ!Q��A���T�;w)���r�'k�6�;�I����즍�b�P*D��`�pX��DG��M���i�豓Ѽix�d�O^%bA�۬��dR���G�8�* [�$�=3@T��kx�T�'�B�'�B�'�r�' ��`���	I��bR�K�>� ش��A��?9����'�?aw��yעܦ(B<X�F�P4"�$�� J-���c�.&���ZM���Ӥ�	�F�3��N �G�)+��?�P(�$�OܓO�ʓ�?q���\-�q횁0P�vH�Wv�m@��?����?�-O��o�
pM*%�	��.U����j�#��)Dǆ�a� ��?�&^������!L<�Ѐ˶p��@���ϙ�V ��~~b�	�3�e�i�����	��'�W�+�|��M�b�N4��%�S���'��'�����3
�� ��H��)g|�#7��ȟ,�ٴyt��?A��i�"�|�w�.l�C����q�̍�b�YC�'26��ܦz�4�\:�4�y��'��p)f��tv��t�d�e�C>v��R�H߅�����OV��OX�d�O��\�x]�m���
����d!���P����)$w���,&?�I&c��ч!Fu�؁9"��~hn�I(O���h�"�'����lJD�>h'.� �D=r�FA�u�ԸO�6m�wyb
Қ��m�����D�>D��$-l��ى��?B�|���O��$�O*�4���C@�V�ǷS��/�p�r���<U�N�bd�Ü�y�&s���0�-OJ��c�:�lڥw0�x�fO~�\܁��P5k�BC������'0����M�J~��� ���V�R�&&+2
]R����?9��?���?!���OW��Iq��*a�NŃe���.�A�'#R�'�6�B"�)�OxnZ~�I�:oJ�(M��)K:P`�����]�I��@�i>�r�Ϧ-�'>��(e�_���J�哶M�-�#��������D\�'��i>1��ݟ��I�7�칷'	$Z5�*���40��Ο�'�R6ǇI~���O����|j��'�i��L|�9�V(K~���<!��?H>�O���J ^����ѓ72hx���>
�`	H0.Z	F��i>ћ��'/E'��0��6IK �J��L����!�ٟx�I������擖6���Iy��f�R�aU#���p�0#�&dQ�
I	@4f�$�O��l�Ɵ$�����>Is�i���F�7f�d�q���l�p8��yӦ�$�� *�6�q����]ȚA�Q�O���`ƹ�U�\:Rq���d�.�]͓����O����O����OJ�$�|:3��%P��LbD#'�2��$��DIN�ݘ��'��O����'C�$p���_2L��1��	B�a�kS
�5o�> o��M����4��	�OV4k�y���ɹ���P��#7�F9)0"Φ*��<bR��O�lI>i*O�	�O��/�P�)N6"]��zV�W<2����O����O0�LV�&�G.Q��'^��>=�8�3�M=y� }A�'޺��O4A�'�2�'�Ot� ���m�9Y"잩��cԝ��s�@-eK�lZ���'Vɜ�	���q�h�_�*��V�4P��r���ҟ��	�����4E���'ߔq����8ެ�U������1�'9�7��"?�����Oz�oZM�Ӽ�Ҡg\�}3�D
�VA"}8q���<q��?y�is��¸iH�I+ �>�  ӟ� f�U���
[�ѴK�D�gA?��<����?���?���?��hʨW1d�QD����Â�H��d�ܦ�h�ן�	��$?�	�{�Y'�+/y��T&���PX��O�}m���?I<�|:�!�1�`dD l�ޡ	&IͦFv���	���d�$(���E�8�O
ʓe�J=�U��W�<h9�O�&G���{���?q���?y��|�,O�=o�	��=�I*~���çV�P �l�wT6V���	�M��b�>����?Yտi�t�z��N�T� �ň�;�؄�E!� tϛ����cSf�����:����p�wIßWR⽐��ҍ1l4Ɋ�'��'�"�'2�'���ec��������m��@Q*�Ѐ	�<������^���d�'��6� ��_+xb��
�C�<8�<}�2n4:���&���ڴћ�O����b�i��I�V"���"斃2��]�7C�VeX͘�#�;-f��+���<����?!���?Dm£S�6��ro��F�����R��?�����$�צ̀����<����O����&j�
�(���6���Oj��'K46-��IkN<�O� ��c���*�n�{cC�9�Y���<v=� �i;���| k���$����cܤ��W�P��L�3�ޟ,��˟�����b>��' �7��
t7*�HA�g~��Qu�N:�\��e#�Ob��Ԧ��?m�>q��i���{w��/ ��Pˉ�$bEz�l~�HTm�z2�x���U� ����?��'�T�ץ�>b�ظ�0$�*��8Q�'Y�Пl�����I��p��d�$@ڶ����|a�� ��8-�7�K�A��d�O�D!�9O�nz�� [=9B��	ufް	2�RAɁ�?��4�?�O�O���Q�i�dO0_*S#�R+Ov��� �<^���1>�f���D��Ol��|��%�:x�w'�3*�j���y
����?���?�.O�m5H����I����ɇOk�
?���r�ݑ}U�����j}B�'���=�d7+�J�*r��9"����f��X��OF��j�vRQ��`�<	�':'��$�?���X7F���a�5�\��,@)�?���?�����l"!L�j�fa�a$�%�l[�ԟ��46N�����?�%�i��O��<k"����I�>h|� (Ѭ|��$��1����M�r����M��Ox�jh���&�W�05v-sC��s�e[��ȾN,�O�˓�?����?i���?��
�j\0�T�*��\��;s����DO��y���xy��'P��|ꂈ]�o)td UC�K�t���oy��'|J~�5 �"G��r�*�b\40`�4+�T��q�;���ş'в$�e�^�O��Z�f$ӃbJ `���W�js�a����?I��?���|�*O��n����'	ش#�/�]cࡑ���:�0��'�7-,�ɼ��$C������M��#]B�&T
�΁Z���5K ���4��$�.�.����UD���0�.�:��1�`H ~5�A����-e��O����O����O���-�ӰxV2�R�h]90_N���җD�f��韸��4�M[����|*��A��|��Ǯn;�8:���1a��XHtKB�	xO�im��MK�'+���4�yr�'z�`�B�ʌ�↏+R ��sG��I�('�'�ɟ���۟h���
���ŋ�=R9�׎N3B����̟��'�d7틵[n���O��d�|�ˇw��т�'s����~~�+�>���i^27�y�)���˃X�D���M43�̚�k��)?=��NV��M#�R��t���,�d���RX�U��$�Q1
�"sK����OV���O��i�<a�i3�Q���v�~Y�PJ��T�qH>{�"�'L�6�9��+����OD '�ߜg��M2�a�)-��S�b�O��mZ���oZQ~b/Χ}�"���W�	S--�tI���?O�2T0t@4 �$�<���?���?i��?�+�캥
���|I�����mE�a��Z�	ß<$?��I9�Mϻ��,�5m$l�����z{J�� �'қ�-��O����O��$�6�i:���`8�(�B-)f2�8�������&):غ�1騒O<��|���}?:�a���V)��AUc�q_�����?����?�/O` m�&#�P�������iʸ�wF�n���Ɗ&͆��?��Q�������L<a�j���m��,Y��S����-)p�U�[���|�P�O�h��krݙ'�҄)D	�qhZs��+��?��?9����zxx�¸U��;nr���`�������юH�y���M���3�?���?����4��N��Q�&<��V	p�n �1H8w��d^Ӧ8�4�?�B �<�M��'U�X	A�ơ���r���t��}�P�T�M�;��%ƙ|]��S��P����,���@��� ��� �.�.NCǃnyR�n�䨠�Ǽ<����3_�?���.��ZV�9:~�,ڲȕ63o�$�)O��m�>�MK���h�R���*
�5��EI<yP�!��fP��3����#�� ��f@�	Cy��)�^ų/�:��ƭ^M�R�'��'w�*�O�剿�M;ū�&�?9�\r��0a�EVb!�ٓ���?���?).OL��>?���MK�uPځ;'���-&�5�ė7p|@� \��M3�'���hȦ��S���������u�Cm�0Ud�ɧ������O��D�O����O��D3���T�,��@�t3@�'V:���j���I<�M#g@'��dR���Iyy�	DFN��e� �D
G���rT��A�4:��O�\	%�iU���0� �E���].%�LP�B�<Dݞ�)����?���$���<ͧ�?Q���?�2�Z���(���Ew衸!L�'�?Q���?I�h��tZ�tHB�?���?ֳ��4��-������fS���r#)��${}r�'�BJ?�4���d�� 4����o>Z	i���0&_��+@��/_�6MMyy�O�z����Z���hh�
KV�:p둿A��#��?)���?��S�'��D��y����H@bրX�m�8ڇ���]������ߴ��'��#���m0a�� �h���b�.P�6ML��dMRܦ��'g��#��T:+OXu#�l�AE�K�)�a��D��9O���?����?A��?I����i)pG��]F8�SB\3��mrFzӐaX���O@���O�����I���3lJ�xz�nB7:�ި+�� kU���4?n��.��Ɏ�o�6�k���G���.����W@&GnH4�d�d���'	~1�� �Ĭ<)��?�q�%SkX�%��L�&F�B��?���?	����$Zצ��$�\qy��';��څb�$��PC��H�L�X����a}�@q�p5m����a7�1���9�B�&V�_�|�'v���G�<Nw��D1����~2�'��"Td�"�a+�ߞ?���a�'R��'"�'��>U�ɎnK�8��EqOF���b�$��	��M+eh�(�?���l����4��i�E�8t��c�I\� 1�Z0=O^��O��n�[�T�m�<���t�"�HR��t��A��7;5ąR�#
M��R%�D.�䓈�4�~�d�O��d�O��d�vC������/!=��
��{T�q��vW��'�B���'Sޔ1B�ҏOv@9E�7 ��A�˩>���y�x��tb�<����M�`��@��i�b���*F)�]����'��%���'��I{3L06�ꉹ$��[߆�{
�f����/'��FS�b�p��Fe^�Ie.�9l�b�<�p��OJ���O�lnZ%._D-R�a�3miu���!>4*숡�\Ҧ�'������V:L~��;q,V%��E���id%�l ̓��?�� �P݌�9s��(�	2"�!�?��?�#�i6��������%���W#�"	���Rk��^e�<3s��?������l��i9�6�#?���\&􌀹�Ɏ?9���b� ES�չRO���$�T�'7�O����J7�1X1�\��RY���!�MóF��?����?-�v�ZQH�D�]�6`���P,h`�����O�)l��M�ґxʟLl׃�n�,�X +� ݖX�eĆ=���z��%����I�f?L>	4n��	�~x�f�4'�5��U<qU�iw\� �WT���R��.�^�q����b�'��7�6�	���}�j��q��%֦��F��E?�8����ڴjL�%�ش���ДL֔���O%�ɖK��Dd�w ���P�@�o���qy��',hHCW�őA{��Z�/N�ƨH6@`ӊ�� ��O����OJ�?=����!hC�����Ř"<��E.^���Kt�4�%�b>��D�Φ��>��Ö���"b�Q��K�73d�Γn��Xp1����$���''��'��DO�"A�T=��,)�Fu�5�'�r�'��X��cڴ3�FL,O�$"�e��)M(><��n��54⟤9�O@`nZ*�M����d��&V)1���8-�(�n:?\��O΍c�I8�j�;�����S�q>��ܟ�i�E�@�6��G�P�r�(D
џT���X��ş�E�D�'�.)��D� l	�184��/����f�'fh7-�!�"�2��&�4�iSte�e���q�F���$Q�<O�|mZ��Mk��)\�Ѫ۴�����(a��IW��#π'[�0mj�\�X�
(���<ͧ�?	���?���?�t葓�(I��m�(*�>9Cb�&��dO��135�<��ȟx%?�	�R舩Bl��9-
�p�L���p�O��m�3�M+���O}�T�'�4ER�
RL�0�#�/p�3��::p= �O0�F�ȝ�?� d*��<	��V%U[ذ�c':x6,�z�� �?���?	��?�'������
�,�П KtHI,N�����r(,Ui��K��y2�w��⟄�OPnZ�M;�Q�����ΌXg��H2�K�l��+2���M;�O��л�b��d�wm�@Rq�ÛGd�yP��s�x̋�'���'�r�'q��'�p郷*"r����C�
�"��0��O����Oj�nZ:i;d��'�87M&�dB�&���F�*{�Y�n�&Zv&0'�X�I�p���C��oZ�<�����H
BWܨ=KČ�~�R����'Gt���3�䓥�$�O����O����J��pK�d8�26M�5TT��O�ʓVY�&ň.`TR�'�BX>9$�$�KEj��VXXJwC8jO�I����O���~�i>q�	�}-h��/ޏ2�`�j��I��I�w��B��*3�Lyy�O���I62��'NJE ����G��y#�%�l�4pv�'�b�'k���Ot�I��M�i���@%�iQ�hk+[�Z�J{��?�6�ih�Ob��'��7�� x�tC�OR5���z0k؈q��	��m��!�ߦ��'z�IÇ��?��X���Iq�|\�UgM�e@!�wDj���'�"�']��'"�'W�+{�ra86�R��-���kR����4��Q����?����'�?���y�nJ))2a���Ue��Y�(X32
��'ETO1�8d�o`�`�)� ��zW�@=w�P��1
� &/t��v5O
��%�W>�?I�b7���<�'�?�rE��:�$���ab�HpC�ϖ�?���?���������g/Mϟ ��ݟ B�
D�8�2U�����&��e�D
a��]��I���	<��(�вg�&pzi�h-z��!͓�?� '_@�"��4��?mzF�O��d�#^#�T	��P�i1��Ir�@)	��$�O��D�O��4�'�?i�II)h@�ͪ���j�P[ ď=�?�g�i�X�R �'��w����]!�
�`2�˔ �>�{�B�+'�牖�M��i��6M��Z6-*?�熟�rVF�H�Z�qfa��كL��J�X%$�̕'��'��'[�'�h�RY�](�!`A����)6�前�M�3�'T�LB��?��'U3�ub���?a1e�7l$�e	�m4	��0�f��ZW�I �M�s�'������O�����$\m�K�鄉9���I��� ����>��	'qLl���'��x&�h�'��:����`���l�5�BL��]���I����i>e�'��6�\1C^����GŲ�KPƃ� O��aBoRJJ����e�?��^�<��ԟ��ش`Cv�3���B������N5*8h$)�I��M��O������Ĝ�4�wR�}�6��<�)�f�t��p �'2��'xR�'KR�'�,)���J�eI`�g�U6)�P��B�O��$�O �o�{�R�'ic��|�hW�J��Yp�(M1v�ۃ�tO��l��MϧCq�](�4��$ѮW�BDõ�")$��6Łm�T�j� 4�~��|�S�h��ϟ,�I`�D����<��%��	�NZ�	[y҂f���	d��O��d�O�	��T�X�GF.n�F<���XŐ��&��s�O��D�O`�&�������dʛ�[�m"�F��6�P!���U&M�=X%�æY�-O6����~�|"��R�H��/��a'
��T�_�x��b�6(��E�3a��Q����H���aM�P^����O�lm�b�_z��2�M;�o�L�ED�<s�����)ڌs���M~Ӥ,�¬d���l�MUİ?Q�'�����R-\D�a��+J�:"͇�O� �bćO�(q A�5��Z��W'thP�b��:D��ς�[�h,�PɊ*(J��g$�8;
�l�w�	9���"bE�/vR:�cȍk��(�
�%6qhiB�5!9��X��v��S��qo�=d�\$�GA49�"e� k�Y펍�FN@�l8,�3r�U��N�1�m�3x�,�j�B>-�r����4?&� ���"L)��$�n������6ዲA��a��A�>v]@1��>7<�P'�z<�=7�N�H%��B�O<��pdj�,N
$���y���ON�d��`4�'=� ;��Dk��AzF( ��^��)شNRXy������OCB�UF��l!��Zs*�eΘ�f�"7��O����O��R�l�d}�]���	B?1W�J���������ئe'�,3�l�ħ�?���?�R�Y�ک�`�R�lxzq
�B�,]��6�'jD�a�>�-O�D&���h ���ԋojfZ6�(m�4�FT��i4/��\�'��'�bU��p�H ]���D�#��ɀc�l�&��O2��?�L>!���?y2�E��8u��!`A��h��ɷC�X�<����?!�������ΧYX�I+�F��}��(aa�A��n�{yr�'��'#b�'Ĝ �%�O�TD�H)R�2�h�B�%|�z��X�P������TyBcX�EZꧫ?Dm�<$��]�a���9���	4i���'�'7��'�������
�W�X���'��X����r�Q�x���'z[��Z !�����O��$���3��S>j;D�U��m��D%�r�	۟\�	���q�?)�O֘�i�+M���q�+K��Hڴ���Ȕya�Qmɟ��I�\�ӂ���ƪ������>�$hx%�S�V�6��v�i���'�h�ß'��'��>���@3J00qMc8��I����TL���M���?Y����P�t�'��a��a
�+������7�"@YQm|��-�QE2��F���?)0
0n��}���R�ȡaG� fٛ�'tR�'�L@@�>�+O��䤟���JO�bE� �-g2�,��%:��7�Th%��������I�*���cH�5��¦
��dj޴�?i�'�5��	gy��'Hɧ5��_,�$��ɑd8L9%M��dS���O
���OJ�D�<)��A�dR$�I��
�V��Q�ֆ�"5�U���'�"�|b�'���$c�T����&`d���J{�d�u�|��'��'��2]�q��O�.ə@�_?�h��Y����O����O|�O��x��h��,Ԭ�G.�	{`Ґb�E<,�1P���	ޟ��IHy���2�J��+)S*>�>�3��צQڶ�j����e�	G�cyB ���b�~�ֻ���)� \`�:$h������ԟ �'��p��=�I�O����Br���7a�Ј�b���z���x_�p�	���'?�i��ːJU�lA�(��!ļJ8y@�v�P˓ZTQ��i`맡?�����I�ru��;�"��XXP1C�Х'�27��<���?і������4-!6�:Պ\Lx)ʤ���%n�,w�Xy1۴�?����?��'[e����&=���u��TD�S��6��L����O�����<y��$�NP:6��<��-K����X״i���'"m���O�I�O �	%�h�c-^�bt%ҧ��	�@7�O�˓<�iq���䓔?��9�������A"�byX�!�vӔ�D �I��L���P��`M���FS�f�T4¤FD�K�MC�Y��z�ܙJ��c���IRy��'��� 6�Zg�u���G��&U"��@H�(��D�O���+�I֟p�I#%����c���hTxn�%}<��FR3@).b�p�IyB�' Ƒ�Pڟ�$����	)��9���N�|�J�i���'�Ov���O���a��G6�6��	`�@�����U��Hbcj����?-OL��Ư`���'�?	��Vf�p*�Ƕ\H.]��G�WK�����O��DHH֌�B��x�e�@��񐲧��"Oʱ�$���M[����O4m @�|���?��[��;8lN=�"�W�Y�M�K�I��,�I�J2����h2�~2��Ec_�� 7�wD(���n�Ŧ��'���*��}�"Y�O���OA��C�l}Y���4v\$x�f�Ϝ_d%l�m~���?�������4F|<���ϫ1� �@ōDy�b�oڥ�VPcݴ�?)��?��'����\cNpu[BĲg²��3gՏ#H����4O�1���?����?��'�� Zb.�29�PE���Y� ��К��ǁ�MC��?��.-�x'�x�O��O��q&�P(������V���8`�i�rR��H�GHʟ<'���IX?A�M��;�f4�?W	X0��ͦ��ɪ2T��'l�'��'3�{A��kȼ�F)�J��e�$�d��L��	ğ���ϟ,�'��Z��|�҅+4��U1���7O���O�Ĳ<!����Į�.]*� bԨzL�-ڇ�P	�M������O���O\ʓ�Bj�0��)��O\�[��c���J��!P���Iß\��Hy��'��ßt�n��*
ι�r�����KD$������O��d�O��~�x�cR?��ɒ*����ׅHmH}p�#N&Ei�$��4�?!(O0��O��d�����3}�Ï&┓�(NLGV�@ ɝ�M���?�)O��r�G�S��':��Oj����M��t�r��Uw��q��>1��?��R		�����Tg��	��lڀM��j��RŬ�?�M[(O���Dꦉ����h���?aS�O�.�4CW���ФZ�`�f�/�v�'��G��y��|b��uQt���M����䬝�盶oFY�T7M�O(�D�Of��Aj}�Y�H���I�T 0ĊU�� ����M�g��<�����.��ȟ��jQ�s*����
#U���J�R���O����O��E�_f}�V�<��{?Q�꜄}��]�$ĕ�aGȁa�mQ䦑��}y2���yʟ.���O��Ĝ<�|Q; +�<p
v]��ɐ:Q���o���4k���$�<�����Ok�D6&����F�J|��1�AU�&�'�2��'6��'u��'�rS������o��F�1ke)4a���O˓�?�.O���O`������%��(P�1�&�&K����8O�ʓ�?���?+OR�(6@��|J�$�%\}��BO1�F�� ��I�'S�L�	ڟ`�ɥgrr��%K�\ѠE�3�bYn�JuP����i@r�'���'s��`�����$�����U�"��SB+Z-Zf�oZ���'�"�'����yb�'0�$��x� �@	8���4(�ܛ��'W���%�?��)�O*�$�7@�3���r�սwD�����l}��'���'�V���'��s���'S�b|���u&�'M�<o�mnLy��ΩiQ�7�Ov���O��)�|}Zw���E��#{Zͨ�OԨ7���4�?	��y��9ϓw��s���}*���b�����D�'��A������hfi�*�M���?����rX���'��DX��@�����tp��@�@��v���y�|��	�O���dʝ�~�f��$(�H@���U�E������ ��I�X��Of��?)�O�L�����A�c��?�8���4�?A+O�X��6O���� ��ݟH�r)�-5 ek����8�K��M��H��4��P��'�R\���i���#�)3������%jN.8���c�h��&Y��<���?Y���d�s�\���� ��$Sc���B��e��Jh}�V���IQy��'\"�'��p	���;_T�u�Ԁs3/�:W�D��?����?���?�*O�DR�Έ�|R�Cڼ$�NԀu�_'�P��sk@��i�'��S�l��ɟt�	M���	�y8 �zO��@D��	G�T�n���B޴�?9��?������Ҹ��O�Zc�b�{5����m*f,i5Px�ش�?a+Oj���O�D�<(�1��F3�U�߀g:x	*�o�<�M#��?(Ođ9�[G���'���O$<�a��3n�,9Z3L�<pbY��l�>���?���(�͓��$�O���'+�Y�I�>�j��rK82�7m�<Q"�M1�v�'���'���N�>�;n���ò�>S!J� R�n���x�ɕ_���	����O8�>}:��P�hʪ�Y���|�u��~Ӷ�3M���-�	ݟp���?)��O��9��({g$�5J�0Y`��"<�H��D�i?&L����=�S�h3��ӟ36\��D"�"߽�M����?���1#��{�R�\�'��O`�s'ƞ�(1���EDE�l��)�Ծi�2U��+��a��'�?���?y'f�:{�B=I7(=��d̾-����'�F����>�*O�$�<���[b���8����h�F-Y#��Q}r-��yRZ�T�I��L�	iyB �$s�$	elr����F�ŘB.I�h�>a,OF��<i���?��.���T�����+�/ `�����<!��?���?!����E�1-�xϧ7f��@@�'�T�2� 2,�o�Ny��'�Ο��ҟ�z��a��8�9	| 9���/Q�h<��b���$�O���O��0�ּ�Z?e��9�� � jՄC.0*���dA6o�"d�t�i�2W�|�I�4�ɀ_����v��K�[�pi����cL���$͎��'�BP���� �����O~��Nŋ#bݑi��"o�����u}��'���'Dhųʟ0����+��;���Ղ��H�*���M�.O44Y�EWȦ��������?	�O뎚�T��Q�ĭ�/B��j�ៀ����'��τ�yB�'���'q��=��%��-3z,����'$��F�i�ph�3f�����O������'%��;-�����=��K���6����4|��`��?�.O��?�Ipƌ ���/k��e�P�[��� 2۴�?���?	U�\8e��oy�'c��C�3x�f�A�$� ��Qd�"CR���|�(�yʟ���O����Uڨy��8Uj�{1� Q@(m۟ B �J3���<I���$�Ok,=�i�Ѧ��A��h �#�-�	~���	؟���ߟx�	Ꞔ�':�t��(�2 �@��VS�E?*s�O&���OĒO$���O�42��T�v�y�SY4�m)�g�J�L�O��d�O�Ĩ<�U��+�	�	�z8�/�t��\�KW:z���� ��a���$��y�p��Zh*B�ο\��:���U'���'r��'��]�܈�����ħ�\D�F�{�B%sPf�	"t$��i\r�|��']���yR�>1�ґ^^<��Y�J2�hXb�����I؟$�'�R �Շ(�	�O2���IR�%3�D����|��BT�*�Ĩ$�p��蟸Q�D���$���'H�J-1V��6	����2Ryliy��� j�7M�G���'��$I;?!�G@"d�� ��&J����,ɦ�I؟�u�ߟ�'���}rW����CsI�#��(�����R'��M��?�����xr�'��,����%,����#Y(��Ox��(�%6��F�'�?yPO�uKl��c�8B� i�rb��)ћ��'R�'�b�Q�J:�	����]�z �`��P��&���%�0��>���Qa��?���?� X	?\�{��'f�@��Њ	�ݛ��'O�8�D�4��˟��'8Zc��h�	X;�x���? �-��OQ�#��Ob�$�Oʓa{n�"�Y29��`�7e��Ey���Ƌ�]!�'�2�'��'�"�'+�-�W��Sq���1�~u��+ˊ�y�P���I���ICy'�XS��R�Yz@�оp"�c%n�"SӒO"�d>���O ��*!����8<����㊪/��!�r#�}����'P2�'��]���'C߉��'n���pd�α �|ס?ހ�Ҹi��|"�'����u��>�1͛b`y�.�*�����m��ş��'Q�U�f�(�)�O�ə�'��EؠQ��)�:
�=	�i;��O��������;���?sAb�1���1��MG�P�ՠm�Jʓ>7ȼ`��i8���?i�':i�I�kE��g�+Do�m��">z�6��O.�dҾ0P�/��-�S���"�_�l�"��S�P;N7
6G�kS��oZ��I͟@�S����|��	b�=2��n�R���[���N]<a��'��)�'�?�"�ׇ� D!��°�B�I�7AN���'���'���ꦦ)�4���'O8h c�d�zdA�@ѝ�ҥi�4�?�)O�e�ЈFS��۟0�	ßl �+����	S��R����Ѩ.�M�%�\���x�OkQ�P�3%�1Tt9��D�g���0��>��
<�?q��?1��?�����d�?;�8�i	/us�U8b$D�8i9�cSs�	ޟtG{��' ^l��I��:���cG <�b�8�G<���'��'�"�'���	_A��O�|��AɅ*p"�u&Ǒ+�A��O���(ړ�?Y�-б�?釣ÃYX�TC��wu��"R�I�����ꟴ���`hU$S����	ʟ��B,Q���1��3&�pK����M������?���)��m�1��q�4mMR�p�O*">�XT�3y�J6M�O��Ģ<��ڶR*�S����	�?�Ig�<Z����C_�Q�*х���M���lR�5��On���^	��7��Q��ZF�f]���i���'��`�'���'k2�O��i�q�T��hU���L�(趭S�j�H���O�<��	
51O���y෫�(^�,u��ǟ�Z`���iM| E�'u��'4��O�B�',��]��P���������
���P��4d�N�:��O�S�O��߄մuQW�2.$�������6��O���OTM`��BB�i>)�	����F"�1d�#���v���GM����'J��y2�'��'�V|2GC�<7|��W��#T���lp����ԮH�N�f�����&���P�T�}�(Q��A�>K4���,����Dr�Yv����	�����qy��_l��(Bâ	����D�ڕ�� ��g)���O���-���O���I�I3p��f4N,5#fO5j������O��D�OT�4�
a�5:�������t�hD���&�%����ē�?�N>A��?�2�L}�,����S(.x�Uf���$�O�$�O�˓H�yJ��TF&%&��4���)�:Y�	��u�\7��O �O����O樨��đ�}��@���24�e�ݔ)����' �P�X�m���'�?���u�Q�� �0$���b��nR����x��'����O�$���Ϻ@-2��ӣK.	��7��<���M�g^�6;~����ѕ�� �� 3�T~��kQ�(>�%�F�ia��'c\�ʌ��)�2h�.x�5�F3P��#�^.��h��G�7��O����O����|�H�(���e+, �8�d��q$�q�i��-���d.�S؟���AM:/w$�4G�8!����u�&�Mk��?��a���S�D�O����^6�=צ��4/\����% $c�dCU�#��۟��	���pgi1oZ��Q�_0��m�j���M+� -���Q�$�OT�Ok�$[� ���,G5!4�8���&���S1�c���I֟���ayb��/~*��$ �u�؂ G�49ָ�7�"�D�O��d<�d�O��$�- )X�ýB)�&�8��ԫ����'���'""[�h#�OP����$,��p���kS���o2��d�O�d*�D�O�җc��I+.���
z�x�D\?O28��?9���?�)O�ԘQ��\���'.���G�(��k1��>,s���E/vӾ��<����?���;p��?��'`8&H	�+A��r&L,si�Cڴ�?������ſ�\ �O>�'��dm���7��"=V�$f;kB��?����?�efD@~RU���86:p�s$Ftb4�Ii͵�J�oGy����HԨ7��O(��O����u}Zw%�,0''¬�ҥ��#@�][hEp�4�?��[�:1̓
.�s���}*�-�=K\\�C'K�:����G*����T�K��Mc���?A��j'^�L�'��iNڝQ�ˇJ�!Ȃy���hӴ@g8OR�$�<��D�'���$��1z ��+�+���Ƅe���D�Ox�d�R�h��'1�ğ��ZZ����]PN��"h��% \�>���ZS��?1���?�g�ȦJ� �b�/����Eʵf��F�'d>i��>�)O
���<�������Qh��A^,2���E�CO}������O����O���<a�%�oն���C[���H�^�H�1a]���'�RS���	�����kL���)J�:dG�Ύ�Ь�g�$�	Ɵ�IߟX�	By���4è�.?^l�s�ٿR�}��B�4I(�6��<�����O��D�O�٠�:O`�h�F�,+JH�5K��Y��&Sj}��'UB�'��I8�d�í� �d>?���Ђ�N�$�"�`���">��n�ʟ��'�'*r'Ʃ�yrP>7-Mg��xR� z�0���`+(D��fU���)T��I�@,X�#�Tu����%z��ɬf5btH�� ��TC�I g���c J.�R���_$�˗�QV�X]���u�X�E�GȂ�_J�A���N��!��V�d�T�[䇗#8pX����.�|���A�Hܠ�#@ ˲�B�I�f�<n��d*���9�|�`��B^#'I�\��Ic�b��H'�����#����8 �7E�Q�pP�Q� 0�,YB�c��
Sd��O����Oɬ;/�<��FS���\����*y(���GI�����Θ-��x�ba����O�f�'��q� -�NRQX��Z��Hұ�/+� ���4�����9�.��3J�|�0 X��4�ݴr��B ��1W����B:����a~b,��?�'�hOR�㧣�-Q�|�q��.o@�8A"O����������,X]r��<���?і'�,�Z����,Y6�ې́�{-��6Lٙas&mʒ�'�B�'���`�a������'Mn�2ӊ��W�|er���p��+����X�Hvl>`9@9ϓ,��$�e��d0q��"Q��x�V�X?V xC�	`�+�[<VP��m~�cA��-Jq��)��̟���r�'��O�%`�,ι(Tܰ�B׸X�0hA"O���sM3%B6�{3B'N�F��e}�_�tB�	����$�O����4��Ei₄0'�mz���O����1X.j�D�O�擠 ����`)7�V�s�'82�Q�j��H|�� ��ݕs|���	Ǔa��U0���DwTu���O��I�Aj��0�#Rȴ]���'%�!���?A/O��6�� 8D��r���&�4����'|OTmˤ쑖�XJ��<5�L��eO��lڗ@@�l2�F�V'����F`R �`y¯Z B���?�(��Xy��O��� ł
Mx|��",ߝ3
i���O����;� aH cX#hX��O�a��i�#_�Ԓt��*��� C����	�V!L]�BdY H�ra�Gn��?Y8���Qp\T��I;z;����>}�K��?���h� ��&BJdf�N�GK���Ь�:)�!���(<�H�+�:f����e���axR�5ғO?��ې�~�dq R�V��.���[�����<A��ˡT<�-�I����I͟�ݓn�b����(T � �3Wy����O%�I�2DL�@�)�3�$���`:��(%$�RS�|��Hq�=3}@�!q� 1E������]��剶H\���#��E�Ä8�̡��q~R���?�'�hON%�MX�G"�x��3 1��"O>LrwD�Ce0@�F���h�F<ّ���{���?�'����u��3�2苰�D�����/��~�� 2c�'���'��y���	��d�'�"J����n$Jt�@�$_��N׹4�����Ј
�H�Dy^}�Q,�w�
)�$�� �`����`X@7iÞJ�[t+T%jx�Q�ɘğd��)� ��)��E�vo�!�$�'[��$e"O}��M0I8�r��;B^�b�dD�]�,+�i�B�'�R��`�~'V���O�t�z�B�'�m��A �'��H��|r$Q�?RB�*T�T�	Ɗ�����p<1G-]D�YR��(���9���Z,xv���S�x1��[�	���bG�T�K����D��JC�I*�@k�Iy{�����$3�2C����M�"Q+� �$m͐l����,���VW���i��'�哐88��	 /���1DG�z��M��`ӟ|R�)�	ǟ<��ԍfvE�$�����|�+�A[����L�����1��>���NA�ab`�v����'I3$�Hf��s��$��ؠT���'�P1i�ɘ��O=�QT�(���#�B��U����'��@%����C��y���Ó�X��Wm���v(�x��릋��M��?��S!T�q怯�?���?��Ӽ�-�[rlV�r������+0z�
P�;O���Ӻ	������|�O�H��:d�ñDЪ%
��*�x����z���̶lƠ骋�L>�2b
�c8̝���ŠN���c�$��'���S�g�I�#4�� T4)/$Tp�A��8B�	/p*�s7��;9�X]�6B���@����"|2 O:NF�;B�Y?y�Bx��`�9�Ys'�;�?q���?��M���OH��v>1��R�O+ - N߶j�.�PĬ���C��'xGXD�q��MN��6dH�L#l*�)�X�q�]�}Рq"�ˠ9,��&݋<���(�O��8���:.���@ړP�Z-s�"O��P1�EL��b4H�Z��0�q�Ni�(}�C�ivB�'�ֈB풴	�>P���R5K�x�@�'���ոlw��'��	Z�?b�|�e�.mB���%�NQhG��p<1��O��FB!;c�?cY�9�&�ӓB�@�㉍����9�Dİ?�<����J��M!�>]�!�D:{\Pc1�ϸA�F,*���6!�!���q��M�<D�x}��O!9P��N&�I&l���4�?����)�2����"A0���Ơ�2�P�s�P2�d�O�%���O�b��g~"�UJ��qR2�ʮ���$呐��m{�"<����kLLc�{��yY��T�DF6a�'��O��O�ư@��^�p/�\A�%Ä9gTH2�y��'k�y��I�z�JQ�X
��Ց!���0<�!��c��@q��A�F�)�$"�z�8޴�?Y���?9R/��cv�I���?����?�;un)!�o�7<,�[��֓!TB�Z�y�ۈ��<	�l�r\䀐F�[!^R�b�fܓ)��9�牔1@"`:�m>�x3��[�(�0��<	��[��>�O��t'�'*�05�� ë)����"O��9����U8�i�¨_76d������(���Ӕn9��Z�)³g��MgƒM����޹8m"�	ʟ��I՟�R_w�R�' �i�L���Ѷ���C����D'@FHGL����$M�{ r�
$�V'Y�jCk��]��"�ɦa���䉦aEn��� `�:��B�T-~��Ȉ2�'���'�B[��	y�s����&C�?ynv\�'g�4�<���e���@%L"h�{k�3k���<��T� �'Uf�#V�iӺ���O���*3i�Ջ�#P6���h#E�O���Fc9�$�O$�ӻ�A���
&�pa�'
1q3i�y��h�`D `8��z
�z>5;����"�e�%�O��K4`��$R@���;�-@T�'�z�h����	Fd]��a>��L0�>����(?
� ���|�ԡ��ϒ)oYn����W���,U�@�j h��)�'ǘ'��\p�	zӎ�$�O�ʧ1a�82�"��7��Q��y�R�J>HI�����?�UL���?��y*��	0\��5���,���#Q�ܫW���'\�b���	\���B2d�c�����>1��A�S��_�<� D���4-��_�2ͬ ��X�{�!.N^�B�I��l+>Y��	<�HOf�Z��\���RC�1HR��a��Q�	ܟ��ɅA,(,���O՟ ��Ɵ�i�{Em^DJ4�R@�L�P��D����a.M�q1�$���;��L>���>;Jxp��N�U���Ş�g���PE��A�4XYEEöc] ��}&����Bҙ&$�G�C�[������g�X����)�3���	S�ap�a�F/:�q�n�!�� �m�ʮ����7d�	�ɲ��02��4�4�O*�ǧ�W�����D��� �+&A8v�ˢ��O����O2��ݺ3��?1�O��h8BEܕ^6�tpa��`=�T"��x2�ю�����R@`Kօ��`yT9�'��Z�OY.|%j�e��5�;�I���?��SDV���Cr�je���P/����ȓ3�N��`ۼ!�XMbD#07�b��<���DU��(oZٟT�I+q��(�AȤ5�aI#�$zd��Ɵ���%�ԟd�I�|ʳ�e57M*����BL�rD]qyq��*R�&�xB�
��'��ms�lX�<��R��%�����b��h�Iz�ɮ(� "S�[�d_��P�-�-?
B�	�I��fI7�fX3�舲u��C�� �M�qb�-h�x���@H�@5#�v̓;ݞl +O����|�5$�6�?�q���5P�1�P�ũ@i�%�W����?Y�g� S��ԋj]V���kEN?�O��s�E2��H�Yi8�ѧ��<?"�'��C @�,M1����`�O@�<���Z!����U�<��2�.}'�?9V�i��"}��'2�$49��� �pțE*U�1�'M����ő�}�呫;ռ�s	ÓPq��H�� $X�P�:Ec� iX΀�)��M����?��,lSa�&�?����?A�i��T��и���	��ᓠ��Jc���P&*<O0�2LC ���E�n0¨9B���,.�yR�_��Y���O�5��JO�/$1O�%�������6pȒ@�9`�*����(RrT�� V�X����'�P�i�؍{�8��'�<"=E���W{�l.��S*�5^a���p@V1u~���'�"�'�a�i�I��̧z��y��U�\�n�W�N�'m��g�@F<A3�?>����gO�M�i@����m���=���3$CR�t9P�R4�I)x�X}�A ��P��	/��8��L]:��Y�ćК��C��f���BGU)"�x#7K �bc��؈}�
L$O?46M�O������F�X�����A�(|�n���Ox4���O���j>���O�OH5��a�d��Ñ�׵o{n0���'[L[�B�?e�<c1FQ��*	�c@�
�p<�`��ٟ�&�$��X��0� 4A���r�3D�|��"\9J�P�{UNۥ!3D #e�0��ܴ%4�Q�L�'A\={�M� ��<7�@L����'*�\>�sc�џ`�4��1��@�(��f��]c�!Kş8�	�x��	
Ŋ����S�d]>�����"Y����҉�4l&}"�/Hf��P�|��4��t�j�N�d/���iԶ��ɾ���Oj���O��?�����bd��XDa�?l�1�C$�I�����I�aͰ���F	^���
���[�p���@a�'Ͼ�Ru锋@��I�%焬B>��(��{�$���OH��)�.4�J�O�D�O��4�L	����,�1s�� k6��#��4�	�QU(I
��'���&�?@I��1�L�"8� �{�ߑ))J͆�	�O�(�Z��NmaV��"U���IG~��3�?�}�I�����+�\Â�
�<qqd�/�>y��/�4;�HM�i����5e��H7�,�����D�O��<�r))�U��
�!��|蚈�4�'5���ת��as!��DkҵA���6���9���+�!�$+��DB��+�L�b��	~�!�D�?\|J��2�Th�B�ʢr�!�dJ�Iܱ�!
�����C�۳!��R	GN�$�R��6��@%��7r!��'ef�X�hj�j��K�ei!�d�q�T��oҠeV�{�˵sM!�D�K 2�B�����R%��,;!�d� A�Bd*C���W�,�+��Q�/!��J�xe��j��ǋ�\�Ze�BY!�(X��%aѓT���	�j�-�!�ܦb��t����&2`�z4$�{�!���tB�A�(�h���3����P�!��>6P��:��'9���Y� �<�!��̭;���+��[���a `�9u�!��  �+��/|	b�#��:����"O�h�Ă%LJ䫅��q�z��""O�IcT>S�hYu$����U+ "O�iS�#�����8S�T:v���"O ����:?��e� �O��8��"OLxq�K�+s�b�x#_���� c"O>��FC���ءe�W�P�\� �"OD<yū̾��83c�S I��3"Of�QdK<u��jS0l��7�3D��S�i�q�n̓w-X�t��X�n1D�� `$ݘRG�����5Ya��`Gi+D����Z}R%�4�ȕ^�ț�>D��e�ћI��0b��&Y�^��b�>D�@ E�=����V%�J�dd�ѧ'D��I��9ØL���_�-Lr�1�!;D�,ڳ��7`!ND�c+߂-�>0� �$D���,a�.�{���*�P���4D��k��C�D�씻��D��b��1D�����*u&�q!����n9�Ђ0B1D�8�c�,~�Ti�4KQ�`J�9˳l0D�h�·z�>t`��0�v�(�2D�ԣ�lıx���M�
��P�'<��.�&iR����.=e��T��kK �I����}�|�'̔kJ�� �i�@�'�w�T\�A
�(9�]��';����"C^�۱#_Z i����:3���w""�'/1�0�6E�A^r��^:0��ȓ5!0��u��>SRȹ�/�9.{\�X�X/�sU�|���'FL\�	��Wl6ɩ���/t��p�
�'t�)��˅Z�"�x�
L=��R�'W>�ڔ�ƩRha{bM͞Rr����K+$ȗ�7�p> ^�C�Ty۴S%V	����a( �A�ѷP�v�ȓm�\}�O
�P�
E���k�b�Fz�c״a�.}Ï��J�����/g��M��( �!�d�5a��`�R�ܤ#�T�����!�Z�A��ip2H�Edl����l�!�D�/.J�iTӸ_O�|ѧ�N"c}!�����aZ3u���s�IT�o!�d��$�A�(�����Ƣ�)>u!�ĿN/ұj+�%|����&:k!��	B���(_������-9P!�A"P� ٪ h�R����#jG9!�$"�YX&�=�~Ah�`�7?2l�O�ștC C���H?��P���U��uk��� q��Y:d!#�Oy� kC?�:M�b�I�����	�3��K@��: ����~�����$	�����ڇf�ҭG}bg�;�Zm� �P�]�O���íP�b%�dr�˗�}T���'/\�VH�cL�)�ҡ@�8��'R��X�NC�%JF�Gr>�3@�^�n��IX^2 �3	3D��Q��7(�y6��'z�:,���"��ɱ},��Ua@j��g���y��)� ^|B���+8bU��	�\�ZxRܘ@����b�-4�*�͒ 5h<(J䯚*)�~��ǒp��`��Dy�n4;�� ��y�&3� d�� @�L`Sc%'�y�`5kq�M��?-�r\��f���y�(F�EQ��e�P��=!���?�y"HТbi��HC�+F J�ˤ��/�y"Bʋ	�8����X�o���2U!���y�+	`@ݰkɞl��r�ߕ�yR�[_F%�č`�(���M�y2�����@RhɌD,B1��V�yr��5M@�� ��=5~pɐ�`��p<yp��t���!KR�	���jqE�
����f�6�\���)B�zBڠ��'��C�oB��w� Q�Qz���>)��C��q�f�L� �%ėB�ȓ�� J��
)���Nϼo+�|���^j�<� ��� � 1s�"�+ ������y2π
r��Ђ� )���r��	��Ɂ7,A�p���p��XҐ��/^���Ă�L����+vL6�;���&=�5�"��n�R �lۏ~Lmїi�>��"x�I3���J�4�2�s�����S��@��6�|�`4�	(e�����K�q9�A�k��`��
��^�4�*�A�'"�[S�&m,�ȩ�M�韰�u*R�u��x�i�r̒ ���J	LTb�l�0�"�$y�>�{G%��*L��'d��(�R�(pс q�D��v�١$ɒV�V��,gJ�At�4��0��/Mڼ��$H%w�,�1aJW>�,�#РŻ?Ts5Ί7���2��~���1�t�3���VX��H�� ؚq�ל!��|X"�B����1o�O�����C�����!H7j�8��>&��哇ƚ:��v��>Y &�x���Cc��{u^�g�j�����'�!s���:%�%I��W�~�*я{�R1U�p��;$���j�!Q2m��Q����2cbW�G,�}�4�C$2�u�c�G8w�fd{�
�%�8eC&�H7}Fz�3gjG�����q��7>����M�j}N��1��9��q���=0����>�8�r��~=���E�*�N��'�M��l�v4z\���(�قuȈ�N�] ǣ�'n�a}���	����!�
F�D:#bX���q��d�j]r�a��H�jeH�=��	�Ϣ�7 S2.�̚R��92��AjeT
���qo�m����J��\�XggR�7/�| @�#z�v	
��J #��0R��A9��m�p?it-��^���
&�	�,{�Xw-��F�B���z�v!��cF�+2�$Q�T�~i����O�Z��ۃ�B�y�>�HY�2Ez4{��¯H���/��$:���H�=�ņ�/x���T�C��@���4ر�I
��OȤ��T�O��0�
I�;(�娤�\�|P���r�	=#h����C�jJH���D�W�2�Y�{�����e�⌨}Ҭ�� �"J��s�J�!���G����>	��Uąy���yr��`���o��Vi��&O N=c(�?��H?9���hh۷�Awϔy�"F��Yt<|1e(|OD9�A��7q�iر�Y	z�Șk�*����*����Y(��-]$L�@����R&Z�Ia+�x���B!�R��B�tLɡ]�jȰik��
��O�\�s��7\(���E!�`���'�|�Îu���y�F��$1À")���u����2(�9FLH��iך k�#=Q�l�0H��U�I�l�$U��<O�� �ix�<����j��q���O��Q�Y�,^$T
Z���Q/��4�h��C;��	d�^u��I��6��|�D�E�>���`��J�LJ�����4�Z��c����iɴ4*��*�L;�I���;���rUO]�]m92u�,�,7�O`����;��k5̄(%�Ƹ*3L]4\�:����v������9ʤ�sQn��d�h��q@K/m�+W�ɞ[�>�����P�T����h����ė�����µ}�F���l�J`qǢ2`ȭ��$�j|����Oj!r��**�"A�¯�1A�`s��	�OQR8�K�&xԔi5m�T,��
��+�b�$F)X�c�!Z�@��}��Z̓h�QB@��;@*�  ��1(�	�n	D���"�O�!���P�� CMU[��*	�>��)mI�I��eQ�;��|�2����Υj��![6�J?C�d)�"O�T��.]/5�|��)�dm�I�R�L�'���O%m��P7�W-2�H�O�2iߒ&6d�r�5ȮpY�ܵS�,kfK6�̕����%+��\�ι~j��O? @����ǀ�05��IԎNw��A���;�io�Fq0��Q1��Gz��<�)��m�<	��q�w�]1�PM!��)X�ȑp�=���,�1O����콲�a�;K�T9�(N�����	_��Gz2�+*�D/�m?�"��;gh��jCHG&z�p@�C��iR(�q�'�1O������',����w��-��̇�tA�r�3E�2b�yr�_2`��r����b�fNEa"
%k����� ��h��	W(ڰԈ���3���|R��i����v!ƖB�|pBG�P_�̴(7��,/�bm+��4���)O��A}��AJ�	8>��aש
L�0�i�:I�3	�G8���pO���	��V� ��Qɨ<��4�n�c;6�є-ô31*h2�C��_zȷ�ծ�0=ѥM�J=���bG�,����c%[�FK��I�^��QT-Wn�Iʟ��'�l$�g�y;NA�9�Y�l�1%i� E	��}!kޱ:!1O�| %cΑz�Q�)�N�d ��R��̓A�T˄�H0袤��M�H�'��������M"�o F2�1��d۶��M��CYzx��d�5v�l�4g��0%�����	��|�'s�(9�`5j��$j� V0��N��sVQ�B�^��p>)c��� paϏ3{v}"#�Uy��i>��'��٢�����Pa�ўqҎ����-3az�`�)�h����Y�0��ᄒL8&�(���(��a��U9�<9U�=oШ���݋2L�Qp��{���E��,��e�H<c�1O�a�X#0���'j�d�H>���9CT�ӷ�-0�@%bFg���p@$`Bo�B�ܓ7LU=���=1@�������W�A���8C8Q�����t*��-(`c���a8�`@�fԌ`�lQxRA�X� -���&t�F�
b�'5
WaH�(
�d�%AS*
�֝aO>�!IC
��<	#˜�%��̀`�AS��1��&S��p=q��D�/��˨On�p��]t)���C�D(It(a��'����G�T	�)c��F/�� hUsa癘y���F�]�r���'�y��T�8�� K@��+{���Q��ۯ9̅0����17d��O>1����q�d���D�<U������LhܓN�2)��"buGj98��<	Cb	C���0!�� ����$*Fg�~]�t"R/V1nz٘���mbhH���Xbub�B���IaX���
N\2��C��
��"�I�I�����c�<��t���oB�y��8w�
P)V 5� ��G�Ɂ !��J-p߶h���6wHf4��HI5y{�y��7�f5��@Y9��� ���i����b/�%��eh��b�az���2c2�ks��)��L���1&�bY9��ۼ} ⫁���=�"棑�|�a&��y���=��
P���'��>�Q/Pp� N�� H�������xy �&�����ɾf�^� �c��U-�oy��i�E+r_:�3
�S.�����7%��D�����'�J%*D��&^�@�c������S�'b��@��ނ��Dpae�S�ć�0 MCUBÍ�D=�����1�J�'��4�z�@��h��y̧h��'re�ւ��z< ykCK-&>L��'�rd�f�6�h���@�Z�N@�#�%�mQU�(O�tآq�}rz1��I!\�^��@��4o~z�8D�^�n�t����%2ܤx�׃�w�t�� �/� ��Չ0G }�t�Оaޜ���A�Px�ϙ !����9o�x��A��dW3�ޕ1􄋣l,�8�dI ����Z�6���� M�TE�<+��Y�y"F�;H?L�s'Ó7O̺�J�Н+ⴼ����7�<x����$0ܻ��ԝxB����ܵbv��2�xa�ȇ�yRɍ�X�ȱ�V�[�I[vl���y�%��r�f�8!ȗDJ�5:���4�ybfW(L�-���7@������\��yRG��aN�`k �Qan�k��P��y�c)iL>X�gǎ>,��"�IH0�y�N�<�uZ��͚"<�W��	�yҪ��WX��3`�`Ț���y���Br�T+ËL�6ʣD���y��ݶkd��9�m^.c�$P#jG��y���L�,%y����pbc���y��-�T�&�)r	9�Dʻ�y�H:��@A� Rܰ�Ԧ���yR`"KtJ|�N�,!��D ���Py"�P4v�z\˴MԌCM����t�<qg(;M�����-�}���)��Sp�<���I	/oJ����	P����J�j�<فC��	�|�
��ẔjJ^�<�E�U|��9Z'�W�!g���"�GX�<y��G�n|c�I0A��<#unFZ�<�E4�ƀI���25}�X�f$�L�<��֔<�+��G$[pă0�	A�<����i��ԩJ�Y$Yۂ�r�<1U$�@�8�����
�.�y�<A��^g���E�Ջ?��}��'�N�<����L5�P��2_��0�jFH�<����R��
��
R�ޕ���]y�<��N�/y��Ȉ˄e��p �Xr�<i�!�3Z�d<c�a��(8%Ęj�<1�.�����f�C)��y+F�g�<�����p�3�Lu��ۤc�d�<���:M��}@�
�fC��b��d�<���F�@�&��Pxl� �X�<��d�ЭPu��c�ڌ���<��$���S�Hc�Ԩ%Ør�<�w�BR��tp¢GUTv�X5h�t�<�&��:�H��ED$R�U�3�j�<�S�/o���"$n� `]���b��f�<1S��6#��]�b��������N`�<��ܺ�6ݡDؾv�����\�<���1� JPO��e[|Ų�BIr�<I)<D|�M�r�Hv��ы,l�<�T
{L�edlԾy{�J�g�<� �#�,Po�|A�Ȟ&XިE�a"Ox���)G�%PGIׂlI�"OF�xf��'|��`0� �8;��Yk�"OԠ��	�ao��� %A�pM �"ONQ�V��Rb^��� S�ް-�"O�H�f
AwH0��$���*݉W"O��ٷ)�血���48����g"OLh�A˴z^�P���R� ~@<��"O�܀�&�.�D����R8STu��"OB�ȠJ, '*S�؜�I"O�����RY'XA�#�����"O8X�5j؋R������Wj��CU"O�m�R������ԤANn1s6"O�Ͳ2J� ��	G�õ��Bf"Oh��p�2l�T<yU`ƀd���e"O��{����z��/ȥ �-��"O"��u�N#�>���\�H �,�@"Ov��2c�=�ĥ��$LI�"OL�2"���~g�	� �V�٘�"O�8ʃ��`Bf��2/��2��%"O 0�Cy���A"N�,���"O��S�u�r��Pi�OU�˴"O:��U��wk�m ��7MB�)c�"O �R�eψp|b��g�s����"O��� Ũ~n �����V�4e2"O�qq�P�>/��A L�*i�U"Oh[��F-Nx���嘸A��ec�"O6I�a�6J�< rE�6�|�G"Od�����x羼`��K,v����"O8���l�7��0��L4�ࢄ"O�h@󋌓-�,���
���aY�"O�4�FiV$�骇c�G �hp"O6�i�+T�zU�Y¦Ȇ��ι�"O.��%��(N�*�*2H��y3"O���T)�%y*��v�8+��=p�"O��x!cC0h��3�ŋ�W��!��"O�0�q�H"$6x0��I������"O\��ċ�.�`bI�^�h"O`-�
F�5� 5�V��8��"O$�K��<I����cŒ�t0�"O�	i�̀�z��ݣr�E�@�(�"O6U�GZ�r<P�E-F���()�"O�y V��y3Ȅ1�L��q�@}�%"O�,y�mO_Wƕ�f+|��!"O���m�<�HYБ�� ��)Z�"O(تe��$PWt\B���8�0X0��'��'���h��Ö
��p��N�	^@@�'��8�A�F0�aT!�0 �����dԷk�����g��-[�?W�!�Ą1)���qEȖ%sDePeJ� �!��ӽh2��:��	7Y*|��	2�!��P	)8���X�J�
��%�9N!�O 8�>ڲɛ+m�\��AL��!�D�<2��`���_��h���D�!�D��O7j���D�,�P��2EX=�!�_�T�����C�`xR�ɸ�!��&lB̈w��4�J�ƭ�!��	�y�F䂕D�5$���0�ͻo!�E�n(�����K�����-]�6O!��.�BD�[1Et�TA���r>!��8kɒ�*���0n��Tؠ�!��%)4.T
��S#nW�t`&l��F`!򤝔:4 P���An���Л>9!�K� "���	k
�!S�-!�� 
�I%CI�
�yQB�=|*��"O�-�Ql̨*6D	�n�\^�R"O(1�3ǊC�ʁk+--���R"Ot](���+��ᑯ
6�8a�x"�'��	H���D�R@���q�
�'���FN19��P��9m�%��'���@���(8�҂�@-�İ	�'�
�@!��qM%b�  l�A�'��B���<P��*⮌�'}�b�'��BaD�j*$�@�IJ0m��=�
�'��LJ�O��{�/
_���j�',�@A@AJ΅���ۋJ[��;
�'�P�(�O�S|:��m_�FΊ���'�p&cЎ>��%�g͐I��'dzu�A�8|��Dg� a����'�v��#&�yK�_�K�.��ȓ3Q��pR�r�q+b*�-Նȓb5\h8E�!>���#��Ϥ	~����EȬ���2Z��Eb�o�LM�1�ȓt���Yg�9Fj������@��ȓӆPX�똏_qYIc�Cr'�ݤO�=�J���;q�,;�8�7�T�<qw��0zP�y��+J���y z�<q�c�W�b���'�?OB��Zv�\�<i�'�;f��	�#�T'Z[�x)5eTV�<Y��*r0̄�F���"l�r$Q�<���4<0��5lޅ#=(��aZO�<���_%f�x�e$��N�ػ �Nb�<ys�̼D��x���ۓ �y�C�S^�<�C��:zl��r���1�0˄�[�<�h^.�"��""�:ڎM(�F|�<y�MY���ۀ��K	��A�'�a�<�ҠY8�����.G	U��!����d�<�pG�R��8&�ZR��j1(�U�<1f&�?@�D�E�H���VF�R�<�w�J4��,�d��<	}(�`"$K�<�V��'%����[.SP0j�o��<I�G(z���ʥ�Ȕtt|�q��u�<!���.,�l"�!�%�_>-{�B�I�}�h=B�GѨa�R�Z�읓*U�B䉅LT����#1���්[[�B�	 q��p�Ƈ�5G�c�V��F{J?+��
4D^(*�<�D"&�!D�x���8m�m3�+U P�fT;�o�R"<���O����EU�e��IjęA1�|Q"O��Cʂ!K	z�x���&1�)��'ݛ..�O4�R�+�<���C���@��3"O0T�C&J-!x�)å�ۚq�E ��,�S��ɔ;��H�D��=%�T5����Zg!���c����ݠ$d��+eX3wd!��"a�ݣ�`��d�!4ʏ�C&!�D�=�z��D�=x�j$�4j�Oԣ=%>٘Ө�J��@�%ΑV��J�a?D�Phgɏ+1N]�Q�wF4}��!1D��0�@c�v剷�S�3�H#g0D�����6;����	>�Ȉ��*�>Q��'A�S� dպX�s��`�f��'4��{3�W�`8L P�кZ$ʰs�'���G!Ⱦ`AmCR&!P������D!�f��ĉ3�;^O�� GR����ȓ�j1���(�6ܐ -�$N~�H�<ы��	S���۔�!����X�!�!M>� e���
o���q'��fd1O~��C^<����A��jd���lJ!�� n�� ˔_O�miB�-�P�t"O4=�#k��hx<�c��8`���"O$E�%o(:¨ɡ� *�@i�"O^]I�J��O�/�&j)�"Oؙ�"k�qmj=��u�����'��	J�
풠�R�|t@ɢ��<��B�I�L��r�$�4ӆ BZ+Y"����7�Ʉm�.��I[#{�L��I�B�I�4�~%�bk�z��ۣ%��"?ٌ�)��$�4C3�D('�����!�Ą,�����"��~3���'��Kx�'_�i����'��41M�&3�F��	�24��
�'�6lC!�ǂ�6X"�D>/��
�'���a*��(�L@�c��+E�2ۓ޸'M�X���]|�H2C�F'$p~ i�'B"��ġ�pT�i��/��*��'����6|�Za�֩
�H���'��a#�\}���LM!	�n���'�ў"~
ceب �ֈ��D��KQ���a!�q�<ٗlwt��"�Hx83Wϔj�<b�W�!2��`7�ir�tK�a�g�<Q�'�"-Vmp��O�XƖ���eZ}�<���y������*Q��XF%Gx�<��� 0�( S���$7�:��5��s�<a�mB�+��a�kJ 
I��@�I�<�D��"K�=��͕CJ�xǧE�<A�h..�ŉrߛ�B�K���V�<9P���a.ap��TH\���dT�<y�H�r��Č`P�b� I�<1�-2-\}�ˋ�8Lؘ!�
G�<�
#y��dc�G���O^�<�ҍ�xvP]��e�M�,���%�W�<	�&�<b��U ���
c��@Rrk�z�<��+[�~j̃�K�-#U�����q�<�3�նj�5��N�P�v$��ny�<)��L�J,���ْ=������u�<r#Թ}�$(�7�B2�E�"Y�<Q0B4\��I�V�@�VF����.�o�<	�ڿ~��,�p�S_?~u�e��<q�7W�40�LZdFF�a!n�T�<i�F���7����RTq�u�<1���-�� ��Z#'�!�&q�<qү�9	U|$�g�J	gr!!MUi�<�Gj²�b�����T�8tNO�<!�FčG'`�2�I���]��$R�<�G,9N�h1��f�z�]��o�i�<�ΟZ�aҕ��g�n��R�h�<Q�`��Z��{j�M8�cWa�<	��	 �!�% �<�z�z�e�U�<Q@ϊF���p�c��͐ۀ$y�<ɡ�&jp.�A�!F @���7aK�<C��=�h�RA¤D��`�O�J�<���&$���	�7��mP,�F�<a�,�(Zh� �s�~�-�u��K�<�$A"kAF�0f� �,�:�S�IA�<	�O�W��U���k[�u��b	y�<r(��#`d��W,��f>�I��w�<)�� <^���K/2&7��/�yr� �̸�I��Z�����h�	�y�OT�xԫ#lZ�r��&�Ӷ�y2�M2>�V4#�T,8�(��J:�yҩ
�
�ii���2G��[A�D��yr#3.f&�#���r���I�y���j��mb�߀"��CW!�5�y
� �%�чI�W��e���K!���q"O��B��!��cQ�G�,q�"Of��b�?$���m܆��d�"OqR��S+g�Y�v�N��<�7"O6�x���"�xi�!�ī|
ɉ�"Oj݀C��7p��ʕ�*g� ��"O��
@Jβ50V5�e��TY��	 "O�< �<I����O�T�L�"O
r�V10�0}�E&I����"O$\�q��M��5cV�D+0���"O:X�d���������H�rh8%"OB	���0P;ȍAW���D��JW"OT�aM���xh�O�%�Y�a"O�riT5@ ��
w��w�nA�1"O}ǀ8!>R��#��,�4UBe"O�4:�O[v�p�J��H#dYl`�"O�e�7ɝ\�>�Sb	#���"O��ڴ,��fp��@�aP
gxQ��"O��`���	$<�E0�lJ6ɚ�"O��Ҥ��J�%Y��R�S)��2�"O1���4� ��d烟C�RE�"O�a�O�: R��(ӚQ�4�"O���L ��5?��h�c"O��[��V�Tc��s���	��i��"O.� 'oǒK�LPaȈl8�, �"O�}��:y�:�� :�0�"O�\���n�p��u�^>aa6"O���e��Y��,�M�5�܁ "O2�y�����.�[���i�"O����z�<��G�	� m�ى�"Ol����	J��C�O� i�ɚ3"OzU����1��r�+�C?`��"O��S��Gu(�35l��m1F<h""O��	�a��t�\��5d�8��r"OD �-\���B�Z
��ٱ"O�d�w���f����M��5�"OZ�$��&4l0EU'���"O�`iԁV5J/2=Cc\?x�
�"Ox�z�����.W��6��"Op]����8)4�3�O���>�s�"O��C��
��@��o.Iq`,ل"O:l:+Ng�5B�B�2�β�!��F#z� ���h�R�ȩ��	�Q�!�D��J�d�H%_�1s 1<.!�dq��y9qd��t�5�^�
)!���P��	� ���T���bm-!�:3����b�)\Q�Pm	!��Q��a��`V>H28��ˆQ�!�DM�Mt�đ4l@
�L  ��P7�!��i
 ���ܯD���� �#$7!�9o��Z¤ϸ~�~�:2���$.!�$ � �v�@��@�@��4��*!�� �N��e��Z
��3)�6	!��[�x���sk�]T�A�j��J!�D�8$�|Sv���I �$s C�
F!���C��e�*�!�z�Z"�
n9!��&<��x�`�S�S����i !�D�\I����� ޖ�Z�I:!��9/�
pIe	��T_���i�O!�d�9M���Z�cF(9�|m`�Z*!�D�7	`��� T��JP�]6!����e�7 ײS�"�<Y��C��n�f���^�>�`
ŤQ�C�I4��h��7�n0�Eŝ<��C�)� ���v��2��� �	G�P]�`"O�)Wg�&0�����%Ǆ>��,a�"O��r ���V!�Tb���ê�y�"O�e�u�́NU�	cmK�~��]��"Op�I
R=d4���-a�xAt"Ox�C��-vD�hE+%�"O� ��P���\�&��an`�"O�\Ó���8@�$K�XL�"O>!��<�b� �J7�(ux�"O
�SwB:7��M*U�Y�a�`�y"O4Y��Ag�k�AL'|u� �"O<aY��.T��d@��J75h�i�%"O,���./t��0@V:Y����"OL��g^�>>|��ӅVu7��K"O�JC���5���Yc �쑂"O�S���I�$���F�D ���"O4ͪ��R�r�%�V��]wT�#'"O�	�匄� (jթT�Μ.�`1�"OȔ8%}�1��Z�l�ڶ@�!��RA4�B0�)G4r�q"OB��`�܀e�<��%��R�"O�+@ �k�dys#���:�s�"O���񌘙 ,	����y��Ԁ�"OB�z�#�j�@ӧ�d�fx��"O���"K���<�j5(��T�`��"O�y�f��BUu
2*հdM���"O��â��(��D���)]����U"O�0�P�ոWN�]�`�[��~8"O�Z��FOx�ófHZI�%"Od�ӓ��&[�!�� Z/LIj"O:�k���:�ѐ���	<9{�"OL�+%I�<.[x����ǋ%�M�b"O�MZ��ԏbhf��e�#~��c"OнbP��ij���-2�0ZS"OpT�3���`��\:|PJ���"Oz<�Ve �><�mϡgEr�"O��j'�̑Df̠3@+�&Q*�� "O�J��Y�<�	%�w�"|Sa"O��q ��M�p��Q�
�u��#%"O8q�Խv�Τ1uhN�1��A�"O��i�*rA�@:ҦN)ar�h:�"O>=�����X�XRA�K��(�"O.S�FiR��U�j���"Oԩ�dO��[`#��:y���"Of�8v�3Id8��t<*�xA"O8��'�en �`�B73:}�"O���M��}&�A�$ߠ�h	t"OzѢ��W�V��Qj�����"O.t�q,X�����S�B�,�"O�vY|� �H$j�����4"OxE:�ϛ�Z���F���ad"Ox`k5 F�#��b5��r�p9
�"O.��1#D�X��=sf>Q�r�K�"O��k��A�2�<2��:�0�"ORUj��9:>�P�@�9S��d"OH�+$��y��y&�=>\��"O���U��bvtpQ�AY����'�B:OX\�e�Z(P�yPU��nk\���'"�T��(AKؐ��eI�~g܅���3D��b�N�?pˈ�;�낗EX����0D�P:@�'Q[6�Y�*!%h%;��,D��2An�(?8��!დ�My;7+��i��P�P�>䞝a�m�0�0�ҕ�+D��C�ϔ2D�����(>] I���(�O��)� ��K��;g���i���?d|J�3GT�F{R�'�1O��R3�wl��0]�K%"OBQ�`��$F24���6xUB(b"O��㵀��"��ԁQ���"�b�C'"Op�0ᇏTx���)ݟ5��0ئ�|B�'y~8yc�z62�1��D+,�C�'�b)�B�֧ ��qX�-#D�<es
�'���b��\|hxȇA�'I[��	ϓ�Ol�
��H�E��NK23�i"Ob,3F���i���E��t^�Ц"Oh� T��*���flZ6Z��"O����H�]¬�����2$A��:�Y�����)X()R������f`|!�B�Ib�K��0A`��� ��IG�C�	*9��݁(�J
���)��d�O�����BT~i����i���׬ΏP�!�Z1��0r宐�,�� ����\�!�߼Qۢ�1%:�Č�p�TX�!�dT�0і%�6[�`��
��r<O֔hse�[��lJãG$�z�"O(�۵�/�lQS����?���"O ��"	1!R���W�R�33>���"O� �1	��P��D2�F�I �p"O\q�Qj�q�N���d�F��P�""O�(�'�?�H��`톹S���7"O4�{�j�>f��a�R ;��b3"Ob��qL0(�8 �)3=�l�g"O*a2׉q��E�)��
�"D"O(Lx�N�6i+T��ǉ;aRL�T��3LO�����$��٢�DC�<����[�|�Iٟ��IIy�T��O?N*s�������J�T��'2�h��\�	p예4�Gxt�'WPEj$oU�NK����雙>ր��'"��G.W̤��&@7 5�'x.!�a�?c�b����W0 ļ;�'�������+x�h� LM�j��`���.OQ˵�	6LD�i�� �f!d���'��'��)�-
�k7��7/�� %�5xH��'�����L9_X�퀶A���
�'"R�R��'*� 1�2�L�db�0�
�'��\��ڲ]lmт3_��Q@�'1F@��Ez:P�Q�[_0�-O����O����_	c�8�* �T5M�IK�,Ȏ2�ўP��:0f�h9q%��Cĉ	� S:r�O�ʓ�0|b OUt�tl�sY+!{�`X�K�<Y���6+蝡E�V]m�\ؖfAI�<9&�M�IKh�w��/=�]�P$AG�<e�h�{�L��)���&F��<1�d	�r��]�ǢE>\�$���Ŗ~��b�ȠG��V-~Ȉ%�S;vᱬ*D��J0�"k�nu�̊-?�B0ð'*D����K�x� �r>��[p�&D��D��	�n�`�O�O�
��#d"D�0J T�q��y	�f��-+���l=D�tّ�YW`UӰMM�c�8�g7D��R�%�7���Qn��|?�x�6�O��DHsun�ѷ!O>m(�m���4o0�B�ɥW�(�#���D��A�,�j[�B�I�8u�dhSgԝ!(R��S'Z�>ئC�I�-f �P�ZiނZ�C�>V�C�I�&9ؠ��#��q_�q�V'!,�lC��B�%�V�L��v��e�0a��㟀F{J?��ж*>�Z�i
��5DG=�O0��$��i��l��r7��t�� ��S�? n�˴��&Cq �)Ȟƈ-i�"Ox�1�A0H�P�AI�s��iY�"O�i�ф�'UJ z�*3H���"O<͢v�:���i#y��!��"O��:��P~ڈ���A�o�ʥ�0�|2W�h��S�@��t
s��AhP{cϚ�z��B�	 O�9�3G��;Ц1Q��\7!�B䉻E X\IFG�R�.y���ع;)j�d*��r���]�(x���Q�CS*uj�,!D��R�ÔN���2caM8X�p%%D���O�=i��)&b��0ъdR �6D�p�$��;VM�S�̜']��J@7D��)d��2y����@��x��6�5D�T���$9���E*���+a3D��8��~�R�Y��
�&?�`bC�/D�lQ�H�����:h���) D� ���h@�ص,��%�"�!%=D�T�u�\<L�=�R�>"�
��9D���G�@"w��۔@;o�2��sB"D�D0%Mݑt�m���
�iE�w�?D�xZBN�$a4 ��U���g*OfM���e���3n�7N�D\`���z�O�����R /r��f�ȳb"|A�'ZLs4��e�2x�a* ��'�"H�+(y4�2�Q�RL�@��'t 3��Z����3�O�,��
�'�ܹ��f��E��2��-���'rtu����u�pK������,O:��dR�*��g��$,��hW�Qq`!���t\� b�l���fb� P!�$�v�� ��o�
3���bȬ,6!�ĝL�ɒd�j(s��;!�D��)Mօ(&#"���gH�eў��ቶ3��-�Zr�ݡAF��3����@_����I���{��J�zl�q�uI'U����O��$*�OPuBPEF@�D�s�i�~� 	��"OB�����z���7(�}��@Sb"Od��Y{n ���-L����"OH�`U�$1B�8�kڝu��O4T%�'8�Qaƈ�1*��&M<D���bΖZؑ�a,GTD�g�<D���cH��mAv���"Cz��@%�9��3�Ohܲ#�-�|=�UF�2gi
��B"O
���|S�Yb���UST��"O��В-;_� Q�c֮A�ГU"O�X"�����`!���9>2�� "Ol1���s�qA�N���ˀ,̊�?�O>!,O1��?V�B�Z*�����L�������<	U��yH0�1�)ѡ$`Z���C�<a�S�ɔ��e	N ~�v���$��<���%I�������|���q�<a7kU�S��\`�2�lt�w.�j�<e��,�T�p;W�L$�*MR�<Q���5b��s�V+�
T�ΑPy2�'�����BL�����ھ�k	�'{H��׸y'���� l҅b�'y�pAɈ83�L�*$ES!D<�
�'��Ax���6��<���ѡA���
�'9��E��h\ʭկĠ&�P�Q
�'/F�Jpc��Aj�����e�c��y��Y�~��W&��<�R%1VB���?����sS� ��jԾs|ءef�->�d�ȓnr!���<���G��D�ȓ%@�zU.��^�v����2d��̇�S�? B ړm�'�0y��:l�v���"Od@������eȉ+��Bp"O��!b*�a�8���V��}�D"O�e�g
$1G� S�Hڣ0$4��"O2]Q�Nٌ!�ޭHp
��$�K�"OT%���P�I���QU�,s�T(d"O�H�Tg�.�6!JJD&|lZ$��"OX�0b��#oӰiJ�揄KX�|�p"O�d�f�8<�D(�A-$W�9�"O*�ެ&�d��["9��w"O�RWDE6\$ܭà&ۡXW�) `"O�����Ӏ��0��d�'p|��1�'LO YcdH;O��t*�N/��2e"O���%.�S�D찆n[+k*�bQ"Ō������N�Sė�J?��re"O��a��3h����!�IK!N��2"O�Z�B M*MFiЕ-����"O�dKe���D]�ȋ� PLd@@��W>���
{�������D#�$7D��Cg��a�rZ6�A6kJ�y�U6D���4	٘B��[F͊�z���'M'�Ic�����m�줻��?����:D�����J�T�8�bd��C�Y�0a:D�$�C��Pl0�3��\_�	JbF>D�l�#Ù�s�p�G�:�<=A��<��0|��*]7J�us"�R�l���"PN~�'��Y���n���({��UY�x0�
ƣ�y"�� 2�C�g/�Sn���yR�B�v�����Ic\.���ކ�yb(�5Q��(0ħ˴r��bWH�8�y.�M�H<�g"��T�~�2�E��y�h�MA�Ib����c�f��v��?1�R��&C~rr"I�!�"���,ٲ���	� �'�Ш���B#�\
o]H@s�;Ҧ�B�%/D���&�լ��!�[��<Ɋg�-D�@S��ɄM�	#rJM3$����*D�lI1�\��`��U��I�(D�� �N��=.���L^�2��"D%D�L��A��6�@�4I��j�.�8t$!�Iʟ\D��'�lX�4��&0������������?����	A�g�dM/!�F�dc('��H�+ރP�!�����S�����xB�N�\�!���YB �)�,*�&�[Gޮ�!򤛙H����׍��J��!F313!��]����2/V�F]r�Oʅ!��]�J��̺���Y�ٳ�Nܢk�r�|]�"~�$$0w�4��/��{�b����y��>W�x���H8au�����yb+|<��AT���
R��b̓��yR��'����G$U� �l8��y���6�HB��U k1"���=�y���?V�X���wҀ��Ee_��yB��L$�-"�*>uʚ��w
��?�����t�t����Q�+���q��-_9�@�ȓ6+�M���9��R����vxȇȓ��A�m@mp�-����'Ŋ�ȓF�p�A�F\5΄��9#�@l�� ��|�����Y=4���6p�b��ȓAZ�K`�70��`��*EB�@���P��0��H� 9��i�!z�0���)]����J��|;��o:�,��fD����G�E��2�c�>O�̈́��x!R'X��@�r�O�i�(8����0u`I�z�: ;�E�4t�M��S�? �YpQ�kך!��H k(D�P�"O�i�L��-�ntBJO�P�7"OjU�&M8&� 03���*n?4�T"O����FIo����I��1( ��"O4�2'jC,.T �Rh3M/���"O:\�RaΨp?H!�Y�n��Y��'bў"~���Y+Ji �.S%(<�����[��y�n1��E��C])����"��y2DX$f��Q+��X�ZY������yr+^� ة�7l8\8\��ꄣ�yb�<U��l@rJ�X�v��,X�yrH��h?��HH�]�: �v���y�*6��л�Y�=I��6h�=�?���������8�C�_:6�R]c�lN&�85a��,D�P�"�:F� �q��{\l��A@+D� 6`�"<<*�
�j(��7D���4�F�*j�2�c�=i��A1�4D��k��x �$��8<m���-2D�����K����� �Юz�x��+D��ʴ�W�7�����n͊b˴�i��(ړ�0<�H�.6D�Jр����Jp�Kr�<s�.W�k���,�&����H�<�a��
�rѪ�/��yz5�SF�<�Nט��:�$�&,$�0�F�<�a�@+1��ј%JB	m+܅*�MC�<���Ųf����3��r���q��~�<�ȕ��q�G�=Ų=���x�<m�\NlR� 7X�r9���w�<9Fō<F���3�އ_�$A0��w�<)t�[�;�p��U�܀bX��2/�X�<�e�|.�B��^�4���Qz�<��؊���p�ŵ�Y�0�u�<)���F��)«�.A��`�U��e�<�Ӥ��oiV���˒T�zE�7nBy�<�䄋,�>tq�OF���}iӦ�z�<��ܡ}�f`���1�ZyId��`�<���$4,����v�r�a"�Z�<��(�\��ِA��  ����V�<Ia/�p+(\h���=��Q���T�<�� ��$b�����J�,�#���h�<�!�

F�xDs����80r��~�<!�	M,k��2��������Gv�<1@�Mm�.U
�&���m���Ug�<Y2L�Hw�L�&뛧�a�Ǟa�<�BlL�5x4��a�ڠͬI����h�<i!���5u��To�3ٜ����g�<�0&�Rߖ3g!�u�ѓ�I�<��)+��M0o����.;�C�I��)��l�%Nb<ْ$�(Wf�B�ɖN�L��5jJ:p�h�R�U��B�I�c�+%�Yd<�s��� �lC�ɜHܱ�a헤��i��j��B�I'g��P`0���4-�E�D
�� C�	�Z�A�U��5w��Ź0$�6C�	�aZT�֪I+[�mhp 65B�6�����P� ˠ�y��qd�C�ɻ=�4$�J9�Lqq�Հc��C䉬#@�W��4l��1Z`�-k�C��&
#xiI����7���w�F$K�B䉤2jv�I�MT��zո���$�<B�ɗK��+�>&
d%�Ձ��a
�C�:,�̌��!��FI��c��
��C�IU\���t�'8��U�P�Ň�6C�	 �d4�6$��h,� ��.]�C�)� �K�O�9a���`��Y�"O�l��Ϭ<df��0#�9�&�2"OV}{sŋ�4�B]�`H�%V��%"O�`�fԹY,��[�hϝ�� F"O����0��ehM�@i��{�"O�p���R0��ѩ'�u *!Z1"Oĥf	S�Sfk�L�9KJ�U"O��yP�B�+�R`��	52�ȃ"O��3
�#}�PӪ��5�E �"OPq�)�M��U��o˘mטy@s"O��'�UNZ�q����`�S�"O*`�TرU��(Y��2�6##"O�u�S�(!�SF��<���a�"O"�&Ǐ?�`���@ƽ8D"O �+����G�Z1�%lS�[��ؐ�"O.!rĈ��<�P�qa�C�1d�('"O�i�3�?=��adN�G�}�"O����憕SdN�zbN�[��t:e"Oj6�9$$3vF��6ps��<LO�H�秒�K�@��B�Ga���"O�Q��$
� �����gU4�+�"OL���pd5r M��1K��%R����	��p9��\���E:8B�B�2M�&�)І�g3.�h��&�B�8d�Ĺ��&[����ԂO�4)nB�I�:��eY�H�G�U"��w<B�� �r��P�Zj��ZE��w�B�	�zL�$��`
�>��D��޾�B䉼b=��G���%���ؐ`�=!:$C䉽V�<��6�	~�]��P�HC䉴I�%��П)�VT31��%GD�B�gh�]����0<�a�
�\�B�	)E����&"����f���|B�I3eB�Tb$��+�
���Q-83\B�I�"|�TGĹp0p���)@B�	:N��`����.>֕�4�O"_�C��	�r��6�ֈ!POM��B�	�X� ���0��,#" �8��B�Ƀs�аy'�Ƀ�@�̯8t�B䉩t��bf	R���X�"I{��C��)xv���Ū�?�@�ȇ�eB�C�	% �|� V���J�bd �)&��C�	��44�R�S��(H��F�]�fC�I�h^�|I�^�(
n��n�:g�*C��6j�V���@� b�ݽi
j��ȓa�Xؓ�.�(=i�͚���,��ąȓ�و&������ݶ9����)���"�M#;|�`����O���g�5[���i�A��#11�5�ȓV�p`�
�4�nUS�#[6b��X�ȓ9��3 A�aH4�u�D�=� ���B�z|��L�V��K�'?�Ąȓ�H�q��
,I4Z�r�P+{���ȓT�\0vnǙ)3�t�̇;ڤ��x�x�{`�BdT��k����+�p��ȓ	�l�Jfɋ�q L�S�z�����[��YK�
�XJB�X���9�����$�$�+V/_.v�`��"�:fHK2D�$I�fو9�thz��	������<D�\��ܻ9N�A�d���z�TW�8D�غ�ĩ$"ԌĄ»a���I1D����ǟ8jBfT:��@�%����3D����,B�BE�"!��}��P���5D���pf[�p6*�x��B�h�Ҋ/D�� .��&�B	n���"!(�6��"OZ �1O	�Wv���eo��G�Ȣ"O�%�4D��rP<(8e	ѣOҖ�h�"OLyp�[5P���N#t�ڤ�s"O����6+�~=ʡa,K�&��"O"�S%�,��h�`U�s����T"Oڭ�D&@�*�إ��7ҵr�"OR�(a�e�R0YĚ����$"O�`���C��h�#�Ɂ2�*	�"O�8:�'H���Ug٤	H*-�"O�q��)G�	�hy� �1%:� �"O����*�'?���V�L#6j��R�"Op}�$A�/W�h�Z�F[snL�"Oĸ����<}c��P��A8dC`T��"O��)��N/|�ݑ��n�ZH�'"O��3ALR&=�ȕ�pĘ�Q�hm4"O���r�Ф(i��9�c��i�`�*�"O��Ra�� ��u�P��� 0��4���O ���Ћp��2�KP�����'�0-�!�[�R���RЉ�"̲� b�È/!��Z*c^d�7��b)Ʌ.ͅH�!��,ޝ��	K	u��9@�#�36�!�dW-'�||{�E!_��UZdcD�W�!�J���������1�~�!�d��vl]�uj�������Ð���O2���0�Z�����O����T� �!��?R�8����I��@BB�uT!���#T6��3+Q�R0 컧���q�!�$�&ry~���
!.�`��H��5�!�D��<0��(A�&�ZéL��!��Ӫ*{N����wLx(Ƃ�{�!�$��j�-�Da	�e�\ =	��O����`$��pFN>G�6�7瘤u�!�$���Z+���9[����U��!�ěo�:M�a�V-$��#!H��!�$��W��1�'�@�S�d�$�!�ж[�ZMa�7L��@��#�!��ܗd��nM6R��8`v����!��N�(|��e,�(�EƜZt!�dͤe��H�mK���TD
`!�˴b�H4N� ͈ir�Ғd!򄑢3�<q����'#�"Q���.;(!�d�)��"Bj�(?4u�X�:s!�$?!�By�
Ϟ[0���럮x{!򄚖	�&���*�e�j� �
��n!�DB�n�@�E�W���H���u`!��[.~p����� I��� �T�S3!�Ė4��=k�AU���E*mR�{�!����JQi?!�q�MP�!�ݟe�F� �Y�<2����l ��!�Q;.d�!m��2��(ԫ;)�!���B��p[v��E���P�I�a�!�$�{�� D�B�tvfP�D�!�d�bL�pI�L�H&��!��S�n�1@F�+X˾q8pD
�F�!��ߥ~��9�B�{��S��͜l�!��\l
�K%��(u��h�Ə̩�!�K�B���P�e-�����H�!p!�$O�u��X&�V-[�(9#Ǯ�Y!��R�mEb2�f��|+8鴍�:=�!��G�V���r�k&�IeB��E�!�$$r)��Q��?Dd�e�7�!��J�v�N9�b��']$�5�U��I�!�0�� rThD�	(պWcP�B!�� �<��惥XS ��GŇ*(��"OR�P����bD3��8~x� �"O��X'�ܹJ^�
d��y�����"O>\�#�Y.g
�$۳�żH'v���"O�9#HJ�z�lYIA��q�"O�lUK�i�`9,	��9� C�yb��1x�ҕV��6sb�H�t
щ�y�� Ԩs�#W!iR�Ak��@�yR$a��{4�>]������
��y�d�d�)�f�Z'@�ҩ�T�� �yrj�Y�u��@�97FB�Dm_��y��Z5qL� `�֠���a6���y�㛊_`���B� FHH��ք)�yҢ�3m+�<a�@D��H��h�
�y�("t��)
�CP�4^���Ua��y��"fɼ����0��������y2�3h�E����)2H̑R�ڽ�yRk\�-`|�#gT+N�Ċ��/�yr*�Vn�:�ƙ���y�le�\�G�^|�*Ǡ�y�������[!z]�������yRBR�G(~��*��h68A����y�
tq��P*[�cS:�����y����.�����D*�rM�"�y�o�'D4ӠM�==H5
�$�y2��:���ۆK��
�Z�٪�y�	ьI:x!�G�U)q��A*v`���y�"Ь���g[�8�$L��y"N�E�:�s��6c=��4AS+�y�j�;j4x�c�`�ne�Fo��y��A/T����UJ�[9&y;�i��y��Q9$=��8U���W�JÕ]3�y2H߸�zl0�톭P�6�+����y��8-C��H	54�����jC䉅d#h ���
KB
]�񩂉?LC�I�C8����C�x��0Rm�]�FC�+=/n4ӔkC|��((��3��B�	�P[4L�G>�t����&n*�B�6]"���قl� <����Z�|C䉻d�%���ct�}�G��+HlC�	 }$8�b"�X��q9�G� LhC�I"/�� ��^���Ui�
ݍ�4C�ɯ+��1�В���i�Jۖj�C�I�*��(�!�?���C�3��B�	�A܄�I��X���. ��B�	V����L�GqN���㛂�B�ɪ����)�6uZ{0JZ�h;�C�ɵ�Rxb�� �qJl�R׀Y5ZVHC䉯�L0�0
Fj�`��@/�?t]C䉥=ʼ�N˔;�<)k��#I��B��3"�I�%,9�6{�'UB�	.M��5ۥ���'WNxT*3Z�6B�E>>�y��}�2������M,B�)S����U)	������KAO�C�I�U��J�J45N��G�,)8�B�	�<��Г3���8�@��x�BB�ɤ�P
mX�b����*-�nB�I���q�7H���FK�&�|C��.X��
>I�Ჴ��'
�\C�I� t�ic)ݣl��MQ�Ǡ��B䉎~dv��
�0>���7�ʽ|��B��%e�pI���n�&�H��	�N!xB�I�l%���@dB&X����a�2K�jB䉈N��B7@�ƶh�0�Y-zc�B�)� ���@AX�����cY�gz��A"O��q����|`�D� ���"Oڐ���:]X�#!�� pa��"Or-R"L��r����Օ��"OjP���"	��p�e�3G��J�"O4����ŢZ�X�� V�]!pekp"OT-Q6΃k��P� .S�v%ɳ"O��C ���3�:h""�V�Fk ���"O (�KN������hjA�3"O�t9���M��% �K�DU��E"O�uZ!$�$����*J�W>|q�"O�L���$h�N$�D/�"08*�Z�"O^1��H�4m.*���Ώ(v%8��"O�t��_z`;�mW� n5Ca"O��@Ӄ��+�j<��~:J��$�&��0|���A(p��ͱ��]�@e�}�<9!)T�5�M)S. ��&��f��A�<����:x�X�㰠�6e���cP�YS�<i�@D;t��lÝ߄�˅+�Y�<����oų$_�mz�D;�oAS�<	"R&f�z�㍰
ưk1 �M�<����M�*,آH+8�� �
K�<9�˟<h� � �+
�@M. �G�<��)Χ��4�%<k�!�%��E�<!rjP�Tf~�r��G��`aNZi�<іoηV����h��[��9���c�<)u��/+ �Cj������^�<�����*V����[.C�`�� �`�<�d`à1�ay����ы� Hq�<��ѽR��D�-�v�v���^Q�<с��OS��A�a�.=�q��W�<�r��1N��:C��nX��b�ƆS�<��!�0?�MyA��H���g��R�<�R)L5t�{b�W�an ��U	 N�<�g�����@��[�H���JV��_�<I�ρ3�(ٶIH+Fz����GC�<I�g[4IT,�u�٩W��8թY~�<�7+¼y�:��dBQ"J�:��B�<�s�i`|���Q�SV4�A �I|�<� ��:5�*�!R�7����A��x�<A��\D<T�4ǂ9?~:LyG%]q�<��*�9o�@�C��G0�h��g�<y6E��<�2����9��#�~�<��"�7Q�bܓ�Y�6|Q�+�N�<4B�_R�U�H�� _��"�I�<��ϟ;1=��i���H�����]�<�\�8h�2n�0�CUB�<�&�����Ɖ�yڑ�c�@~�<i�LǼUф��$';#FI�G%�b�<�Q'��z�x� ��F�rrX�:�
Z]�<�� ۗeq0���'T���^�<���K/%�b11�!Yh6�"��\�<�AV�]K J��"����1��_�<��G1��Qd��"}b��r�U�<�s�$��UR.��%�vm{�o�R�<�Fǿvf�t�J�!#H����XN�<1!�k����T��1/�]�g�Of�<y�hƟ%�lA��i@�"�vи�(VL�<�i�#�$@3c��,�F(�tD�N�<����Z<L�XǞ�O(|��c�<��ʛu]�
�䄽O�Μ�b��W�<`�OL��R��W5d���G�l�<��My�n�sEV�"<�x2�AC�<��=p0��#�0
L0T�<� �2��fW�Q��Ė|U�0I�"O$�
�J�a����uJ*Ѻ�"O�)�f"�E>��%��K9D���"O��#�V�_� ��!ێ�\ݻ�"Oj�-[�O��F�ב �p���"O�P�V(�M�Eڳ=E�J�94"Or���mC�)���7��=Hή�Ha"O`Y��E�3A�TNܲa�z�A0"OB�1�F��؋���U��:�"O���� �DtC��ƙ�B�"O��yS�}m��0�F����0;U"O�\`�[���[�M�P�B�"O����]Kߔ�@�D�ں�i!"O��3ϓU^����ү3ª�"O��"�GԔ�ce�%�a�"O޴)U���>�s�A���m�6"O�i�5+!TTq��Y`�d��!"O�����΅3#�=��C2�B�`"O^����3ʖ��6�J*�>H�t"O����Q�lH�1��܍W��I;"O�LR"C�v�z1[a	B�f�p"O,J�,V�#!�d��+���X���"O>듦 ?6M ���kU�C�����"OP��ą�2F��E�l��dՆ�P"OX��]�	��p����i�t5;Q"O��Iu�I�6�"Q(�KS���Ȋ�"ORe�4���x�H1k��Ez"O���H�7&�����#ޛZ���"O��׭Y�T�D���I�qmT�"O��6jF�"����.f氢�"Ol�e�P.�d!k�CϽ{]���"O��Ӕ�Ԑw/&X)�c�>)$�0b"OlH:q)הoR��D�S�4�rݸ%"O�5�!�I�+#�hi�֨R��H!�"O��a���-�= 6�28M��"O1��oS�P�.�"w�	�:�4�T"O
|2T`��I|�!�5J��6�+�"O$�;q�Ɩ(�����;����"O��R�N��n�؃q'��^�&tH�"O����Q��A(��Y/1��Y2"O�	i &+���߫>��ố"O\���l��M�XU8*��! �"O��)�*X�T��:]���`"ORq��l��=,0��Ŏb�z���"O@����"{�N��� W rH���"Ob9�r��^=6()�Bֹ&$	Ȓ"O4D��є$����+�
��H �"O�e��n	�K��:��3TLF� �"O�eq���=�K��̢heB�a�"O|a�3DQ�d�,9��#�� q���"O>(J��*IVĒ"Ɉ"p&8x�"O�=�EL��*�ʀ �k׼hܺD"O�5Yf�G$`N�p� A�v��l B"O����c��j/��X�/�1u�څ*&"O��qЭ/C��d�oĤv�A�p"O��y����v��5��YsJ�sb"O^@�/s���y1���<lĀ�"O�Ѹ0��&9�i���0�0\�e"O� �r�[�e�zY8s�̇����"Oa2�肨b�b���o�F(@�"Ofa���ߺ�����U>H/��a�"O��@/�y���@���66jq�S"O������V������5<�ᩃ"O��d�\9V��M��,Z)�h"O� n���Z
o�T؊ċ�/���"O(p!����)r�X.c��̐�"O�(��H�gDL1�I�%,��5�1"OL̊2� �DgԘDH�;`ą�"O�U@'��g�Y��T}�����"O`t�� =W��sqeP�[�$�h�"O^q�"��'U�0�*a�5��@P"O���5��)%cS![3,�d|B�"OfĂ�E��Ah�c���c%l)�"O}@�'M<��H�!oHO���P�"OTٲ�ϝ�I�0ٰC�Q�6D��"O�$���	�{eH$_��@!�"O�%	)�;?�p�ZR�S?lH��"O�	��	7������-I�-�f"O��H��UF��@�-M7X]�"O:y�b�@)~����C*7Ԕ �"O�q� `_"��ir��T��zɁ�"O�R�Z��t*�đ�@T&�"O&�Q!�D(0�N}C�c�u��U��"O0Q�O�6!_b@ʶ�̣	���$"O����Z �0}�G�Җv��P�"Oʌ���fU���Dgu�9X�"O8����U�MM�I��W�X���"O�|��쒶"evl�f� ��TQ#"O��CG��hs8H��%��<�0$P"O:a��gM���/�y���q"O�����G״����K4�P@�"O�}B�Z�RI!8E��R���5"O�ԲgO�	~]���(Xn����T"O��ZE�L	<
�`b�Y޵F"OH �FCߪ4�2e
dlP�C�"O��'�m��BLE�]16lV"O���cn�����5�}Ҁhu"O�e9�k�I`�
3@%P��y�"O|9�ꃏCb E�W`�4:򼵓"O`t`�IU�i$n[�tb�"Oġ�$n��=���J��Rp"O\����*��Y����p�@R�"O��
��~�2����P'���'8n���o6��@��?����'X,�!Ũ^�H��-�f�ɵ8VR�@�';t�`�y�^1c6N�.�l���'����qF��4��aV�̽0�pX�'�,�8cΞ�}c2)�V�%�f���'��h��h�Y:�������Hq�'Q�ɪ�d��{gJ��,��]���!
�'��Q���m��	j"��`�61�'�TEIR���E4X��'�W�F��'�ڠ�sB��3zIصč1K~Ց�'_��0
�/Z�vثŁ�4F��'��r!EQ&s��m�0��y��(	�'�h�hV+E�AD�]C e�*t���{�'�q�&F �D�GeB�eW���'(r��ŋ�|���S����`�j	��'�R���.H�4�b���I�U��j�'F�Ԋ��Ə)�Թp'I�LC�U��'?�tp���d[<����LÖ�8
�'���K�,L�y
q�L;r�l��	�'��l�l��FxHd��
)V]z��
�'��qH�̪Kxv�R��6b��"
�'�r1��f
pF�!kS��gf��
�'�~�Wn��w\��㮓*a�L���'$�8�����n�r��!,���'..�3KM+;���J�,�2f6���� �x�$I�@-���1CA�m�ID"O\���3���%� �:
օ`�"O ��ݿI"�i%��3	�(��"OBx)գN������NL'w�t�6"O$Z�99���J<V���"O~��B��Y�x�;Ak�T�4-�""On�/zY�f�V�r�R��G��$C!���]N��&�ǽ}w��q2��:�!�$�=,r$,�eǑ3V��H2nοx�!���m�4���Q��Qb�Z0"!��ŏ:����n���b�I!�	�!�\T���Ά�N<#k�)[ !��!i+�@����7��X0��K�% !��k��<+��A�W�������k�!��A&�uQ8�`�� hM�nG!�$d���4�
|�6�x"�I�!�ğ>-�u�S)��{�T�8*Ў9�!�$�A���ׄ˞<?<9��jW�!�D�j"$M�!(��e�,�*����!��ڝT�x�(��Bk��ǭ՞*!�d��8��%�ri^����E4!���Qǚ�{b���������;J�!�DѤE���wdٟ$�9y��Ff!�d_./��Aȁ,��M��� !�dN.zh2,(7���
A0K�:-�!��Հ|��M�gC����J���#|�!��P��x ��?�E1��0e!�ۭ�6dh�"��p�,Y�'�?N!���*wH����U�9����j3!�D�o4 ���>2���菀`�!�B�R��u�ܻ	C�Z�k�!��*f��4ab ź�
����Іd�!�d#!����Ɇ�`��̠'-�iX!��ȍ�"e;��u-�UZ@b8'!����"'M�0T�&$H��lv!���v�4�u˓|�`��B��l��Ox�=�������z�~��$
	0C���	D"O ٺ�O�t\��Z3q �!"Oؠ��ə�wEA����"\ܥ��"O���غM�J��b�X#t��"O�<cdA<4lM�gƇ&i�m
�'�����N0y�,S܄r���	�'�ĩy��Mb�9i�m�nҼZ�'��9&�ޜqH6�b*2�a��'����F�430�򂐋*@�i����6�o�	�e�H�0Ձ��j�N܉�"�(��>����,-D�L�t�~�Q�dН{�Op8�͈GNV1
7%�
M��u��O��X��R5'�ʖ�J�Q��y�n�,��'�ў�b�,'N_eY׌�m�h��C�'o2Q�&�/o
��X��9~x3�'��10H�،�u�,h9*�'�lL#&�%m" t�) Q��'��-q5��f�ry�Bi�6I}����'(֙����}�8B3O�C�e��'rҬC/;�Q˛	B>�9��[8�y�o_��`���aϬi��;)��O*�;��#}j �V�V�lZtl0/�N5��J�A�>�S�'FF�01$��2�Ԃ�A*	����/O�O?7�,�΁��[��,��W�U�����ޠ�F�ܫS7��sw'�"Ɣ�'�ўtGxrJ�O�^ܠ'��l���2�l[��y�Ի����h��\҅�ٸ'*ў������@1t�eS�7	|9p���.�S�� ъ�!<�p�kWJ�a��P"O� a��̵,�4��%�^I�� #�x�C�����Ҧ�Z;��
�g�����:$�Ȱ4ĕ/W�.DI����$.X��$�Q,\Ur��'�'o�)�s�x��NL��`�@��Z�7ݒIsA0�`bz�}bugK�a:d����G���jQ��f̓�hO1���h�hO�Z��u�3�H^�z�� �x�eB��Xe�=�~� �6��:F�M-�F�Z�'��y�K"C,�طI)+�:�2�ҙ�p<Y���
%�N�{�jQ�.�حIcE�L�p���'�J�d��iצ�
��<X
�'-nD����6��Ȋ!4����	�'��yXA'L�Őh !&�r��1	�'���p�$�~��0l�>�%%~̓�hO1�T� �o�����F9V���I"O�-�!�Cp]s���33˖�(S�Iox�p����6[�&H3��]ohѹ�o&<\���Q$�$L��O�YG|�q�"k1���Ӡ`+ ��'MZi��߫v�` ��	�<!���˛(���ɧ*Ϻ-�x�E�&)!�dM�z=��AU옃7�p!�#��g�'�ў�>���n	�N0D��ڠI��� L"D�t�$V78ܦ�`r!XN�(��!D�$k��ԏ|���>[P�0�:D�,��[+/h�M�E��7FΥR�	<LOz��J��%C�n\��˦5��Ҥ�V?�!��Q�� �̒)�Ji��*ξM�!�dؙ.�`m�F&L� ���ڡ�A1P�a~2�Ol�c��������3qx`�:2�
f�<C\�b<�(�%�2�$ �cm�m�<)��<Ȝ��2��;*�@��i�<��՟*'�Ii�b�B�I^�'��&��h��\��:���>{���b-D����E��w� !-8��y4
�i�O ��)�x��&%5�n)�Ə�|�bYq�'ғ������3���8v�|G�����-�#=i���O�,��L�G)2��d�D��4�'��OԢ}�A<%q�	��@�A�9\���ɕY��݅��a�f0H�� 48'���fڋo�C�Ʉ,c��(��8��3C�юC�I�Z>}Hf�s+�j!�R�D�.C䉴U�b1u�P�l�9׌C��C�	lL�`�
}tlzҀ@0q>�"�S�O&�!�"\�h��ke��Pq��'�qOn���i�HJ1ʵ�
�m����"O� i�)@6M�Ib0iL]�nԣA"O�!�	͘;�&�!'���S�2(bD�D �S�)B!G���g�i�����X�X��D{��v�!���:(fN0����*̪��{����>deh"�&9e5\yp��v��=E�ܴ�x���,̱L�����(c�rԆȓU��,hE��.�4x��/��DІ�(�$�1��e�(됎X*���)���;G(H�@2� �^R�8Ub#$��
���&x�"�D�Lc���C�#�~�'��)�Cۃ,�HX�R� "/�����(On���B 2��T���N,s<mH�"O���]�w��]�s�]/W#����'3!��_�7=t8AoB�>���`��H�!�D�$_��xmʠ3��y��l˿)q�}�������
�9���@�U�<�؜!�-D��a�%�|����+�n������7D������^L�(3䎁�z�Xa7D���
�R�$��kY�>GZ�;2 4D�� �BΜ7
ոu�FNJ�\�yP�"O6t
s&G�X��	Q4-X%S���P"O��[p���B��� Q���V�OH��D]2z���H�<Vre�e/	�!��ʦBo4qҷ��'����FB7{qO�����
n�:�#]�-�v(�SQ�!򤆪xIriYց��(�DXH�a����^x�������w���G�[@B�e8OPJ��dI�i�d��H�]p���\J�!��\�'����� �	��m��m�1O,�=�|⡁A�U����1��i<���'�I8��$���.ƅ;�,�ЦE�f&���#D��K��7
�y�s�a�0�F�!D��8�l�/
ր�W�K�b�&)A�	?D�Xr�
������$T�B�E����<��'�qO�2
��Q��ν:�>���Ġf���$1���  Q��q��r��i�@�R�9֬����<��OdU�'/@<��t�hPR��<��"O2�0@ I�+1�xcDHQ�:�P*a"O��!��ABtH��,**���!�'��'w�K�j�@��"���JA
�'P2ԑʙ' ����b���m 
�'a�A��E��S��s�hTBH8�
�'�0ɘed���h�'n�3��B�IX	�m�� z�:98RF��Ƥ�����	�Z����Ǖ�{����?q�E�IY�!���7g&�����D��&�����ʁl2��y��ڢ ��u�e;D��Xv�Q
_�|Z��F�QJ�y9ņ�>�I���O���$խ0�ġ�	u� �XPB@�r�!��[�n؎����O��t��#	+9v��:�O�ܨ�$H4}�4x�)ڃL0��� "O 9Q,��r*����&!S��c8��hR�9�vE��Ѻ/��K��!4�����& ,�c�"�e=~�r����x� �R�nQ�q��D��k�h���<a���$"L��1@�4+d�ȳ�ӹO�!��	4јP��B9oI�4����'�:�IR̓i���5�.Y����8d�0�ȓDIB�[�BV"+'n�H�	'V�j�IDO9k1F�,^<2i��KY�B7�4p�"Oր�6��0�R �b�S�����"Ob �M
�5��\HQL3R��U $"OH�0e��btF(��(Y: ��|�c"O��h�+�0/�Ѐ��%8Y�`]�"O�M��jƠ7�Z�S@��.��%A0"ObES�$ۖ O��БL��/�U� "O(�Kd�:R�#$L���,��s"Oʬ���C[���,]���@�"OR,P0)y5nU K�!=Խ�C"Op!S�(�Q��UA���~�#A"OdMh&fZ�$�8Ep��9��Ѻ�"O�}iѧ߽f�0� ��1N��ZD"O�a�7�Z�x���{�lM9�Y�"O<�Bu���"��|�P+X�4��1��"O�-˶���,(��#K�8"s.u�P"O��YG�D-T`J�j?*r����"OzI���ߦBwR���Hęo.���"Oxt�A��%HX�!0����Ya&��"O�r��΍0֒���@�s1�<0b"O�L�/ݶD�tY���^�@B"O�mqP`ŕ�~�	� �Lv�yP"O"Y��iʜ@�FJ�X�0�T"O  �&xY��߶�X}:�"O� ��U	�&1X`˗ǒ#M�v �"O88IS+��v>"�0�fI��,U0�"O�9"V��N��u)$Gº8�F$�V"OF 9�d�<v���@[:7�FY�"O 4*�+�1�2���ԕc_�4�"O�5 ��#?�:	��B�S*�Xq"O�%P�	�?`��(��A.�`۷"OZy)� �g�<�p��)`����!"O��J�D�.	��`A��5n[�="u"O���GU'xPV �B�W��"O�U"p��Rz8�H oRD��2�"Ol8��K
�A.��IQ�:r��A��"O��(����5S��D�t��|�"O�9)$A��0�b'I�p���{�"O0ђ�̐�M�<�l]�p�0"O��P��U�M�����+�����"O^�Ԩ�3<�hY�$(���Z�"OX�82%V��T�q�C�(���(D"O��G�5�%I�ȊY�v# "O�t�$�O�4�l��NI}��#"OFa�TO�@��DIc�+ `���"O�Z�  ��iU�b޶� f&�	\!�S�)r�� ���%�����>}!�d�2cA�T�%.�
C�B$�a�?!��Hm٦Lxp�<`�F�{���!�ד'"�PsH�Wݜ��b監Z�!�D��Ag� *  ������ �j !�$�y�tz�N8��Yo@š�1l�A��Ӹo8��(�n��y⡉9Y�y7YW�mѣ�yB�]B�L
�C��e�� �=�y"c12"h���0,,���e��y2a:7��ȹD��'9������y���m�8���-������yb&˽�jM5M�<1:��f���yb뉽^4��H]
,S.������y��7]��4��D�1^�Bh�P%�y�ET>-l,PȖÅQFI�g�G5�yro֪Z>����'I�z��ŉ�3�yr�ޣ.���l�%�� BE�E�y��.5lP�Ƈ��$�,��7�,QJ:�B�F����h��ߨ|��92�k� &�,�C�O�!�$K	F
�:lD�8����zH�ݴF���-�E�r��	$��ze`�!�`�	�f+JE�z�8r��J%�ƭ�~��Ԣ��F�(KalH��y�#����jg.�B�2��B2˸'��3�a�l�f铯6�`���oZ
]��$��bA�7��B�I�[��B �I�GD�h�!"6��څ��#ʒ k,O���Y�@��mµjI>��bd��%�&C)D�8�e��E�@q�ʧwFT�� �Y�D5 �D���hj�^�H�A��>�����¯*춱��*9�l��0+�h�r�oڻ������M'	�����z.�s�<��j�v���N���+���Kܓ{L���t��$Q���`���`�`r��1et��˦�T��!�d%+�4����&< :ʓi�]�L��� 9K�i�'er1G�,O����ƌ"�R�JЯS�����"O����H��fQ�14���P`���Q�i�9���J!��Q��I��(��Si�B��a�g@W�i���d��zp���&|�c������#"/�>i�)��O&D�,C�~��K%�Q�@�N��dj$D�� D�Ρ]Y���N�<���O�ʵeZ* �&�O?ա� �9E�����* �t�>Ա�O�h�<Q0d�#E�2l��>#><=H��l}�![�r��١�Bx���"��9���%�"����@.:�O���V+�8k>��� ���r�.W�j���O��R�8䀑�LlH<� !4���3�EIےiD�Xn�'ւ���@�#1�������(��L� � LQbhiWI�>�!��ȲHx�R1[�7<t�󓆗�;q�$��"��*���yy���'(MX�@E�+�,[@/kKX�<�j�`���DWN'(	��N?�ՠ�5!��LZ�H̰<A��44�峳�N�,5��� �HE8�܀b��$ȱ�S��%v��2��v��@�4�Y�ē�nDb��ݗ):��
!���m��EyB!���zl2�\�+8��M�,AU�آ�Y<|Xl1�"O�\1�R�[p��Cs���]R,��I,?�+��<E���)� $���4���5*��v�Ʌ�T���@c�[�Z�d���"���'�6Ųv˗�:`D���	?v]�H�e�5I3.�Bs�C���������s��m�`�ե֬U�N� ���Cf�C�	s�� �$�تښ9�� 8�C�I~��(P��}���вq�x�)܌�	�n���R�x��צ�F�ء��I�{j�B$\�غ�IV478�.U/aDN�Z�%D��Kg#G�rtP��(���9Ԧ �ɾ>��<���:z2�M3̟�v�)��.ɪ�t�^42���P*^X�H���$t~4�R�Y�bt~��6b@<��Qb�{r0�$���I��H�R��kM6�~bÒ[�Hl���[�"ʒ��l��y�e��Q����/��&tLx�ǠS<�?e�
+�n�Xg�6|6�[����?��O&vHp�瀳~z���
?��d��I�Au�͉�E�\��9�& M>���-�,��ÅT�"�x�R�|����N���� �o��4k$���>x����U��3�.'���K��P�l���E7$�`��h{��U(/8�5�t�Wyu�9�h 7}哌_I���̜����H1��^����X��؅�ahڎT�h���]�*��!��3D3b���C�m�<������Ǽn�2����.���A�B;jĻ�ꂘl�>東<^���%N�{��1°k^0F���Dކ1E�/Z�jQ"!�N�P���x#�U�l���S�@�$��8[EJ[�7�P��fOʺApQ:Q�'���(S�T�j�{�0��ʁ�H!`92M)���;庄����>�z�2ٌIY�(ДG:)��� S6�	�����H
��v��8��
i 1��O�-PW@[��6!���|�=�@]�	�����L�8U<������䦭{�z[��rg
F�7��T�� 8���ge�)��Iү�T���C��11���jZ1D��
g#�>N;�q!c��B����D�03,��J@(
���#/��a�sc�H��*M�P��6�Hza6���z ���`�O $�~�F�l}���t�S�Y2���u���p>YV+�$P㾈A���#j�
�)��x�\=i$�	;Jh�f���A��L��(�D�@������Ğ�UI�K"e���te��DM@1���J�J�4i��(O@Q&�� @GV�"�!N�F�*d��fS�<`�`î.Ghj'�w�����֖g2�o��,�u�F$4>�8A`I������#Xpxl#�����4��,n��(�U��$5?�Ͽ+�C�/����ҕD2flKAB�m�<Q�(Ʋs%��)��<0I�MK�N&�h<#W�Zp��[S�#�"H�'�HO��(7+[�z᳠(�38�2z�'��4� ��&x5��r�jȴ{�2�Hqj�4|ր�Gg\�!��d�����a}�6r
Kŗ%��d�C,hаEy�fr ���Д#��@�v��i�S I�����
a�ݪ"V�h��B䉊F�0�Y��Z�B�te�&�A�Z�֨`�h��ay4,�ik��
�h����5dA�s����P,jݸ�k�)�y��)y����'g6�؀Wꐃ4+j����ɑ1��aJ�}�p����@�q#�& t���,Ta���*B,+�OPA�$ؗk4~�8VH�#^�����C~��q��P��M�#DK�5�}�ș*gQD�1�Y +֐�T�+�hON,R�j��r�Xvh�4&5 �'W�����ݑJ����&ɜϒe��y|!��'�� �(5�$�_�B	�I"{� P*Mw�U�Qm�@�O�b�:0�!&���2I	�;�<�"w"O���/�)eڄ�;"h	=�H2�l
��~2�]�@p�X�!�R����� e�t쑁��?��J�ы.wl����@ɬ���������&)$	W蹹c(��/������6T�ܣM�
�hH���ax≚�m�T�=IP��;���Cޢ��}k���B�<�&h���t�Y��ܚ�r��J}�<ِ��e����T��:��8��+Tl�<A�k�Iy���b��!Mt����L�i�<� >DЂ�̤?=�@8����~�U"O�A��O���+��p<t1�AE�l�����Ox<rc��R�R� �҃yu�y3T"O"E���I�Ro�(+�*A��H�2�>O��	�&ϳp����B	z�z��� �U��d�E&)�{�,X�}"��ɦ�#A��Ayz�r %U�z�J�
,#D�``P�O!0q$���
 ,�$�!���G�4�`�Ϟ@b�>	Y@�I�I� �҆���Gf#���` ��i��@'ȭya��(�hA֍�x��Y�ݙB��O8�}�exz�i�F\")�d�E�Wc` x�G�TnqO�}��_ՠ����Z:Hq*ĩȯk�Ե���{<���e��&@�a{R��(TT�X`H�,��D��,�	�?Ye Č �>��8�����|Ӥ	���+ra���"F�W0�h��'fj����g}2�X
0�,��D���"��@������'2� �/G�fQD�$M�pZ���ń�/'�����!K���'Q8Lq��Zj�OVhYݥ!���Ao��W��+A%�V��E�1b=}B��PS/?�Zu`l��F�	�Ξ�6���È{B���MK3ym�EW�� t�fE��k�0����s�.	��I�e�H�P�R#62������Vn�	�.=�቗E��2`3O��u 
Q9��ƍA!�*1"O�IH�Bܙo-���"M�r�
��"O��h��4r)zU��E6��"O������P�9���P%ڭ�"Oh�adM�n�,k�KI�q3"Ot�k��2QT���U=.		P�"O�����Q�N��G�([�m8�"O:��虸Fш��ǂ�'����P"O�t�7EԾn����\"�� j�'@�����ff�Ɇe�j$��H�'*�t�1A]�l�^�)��?S����'0J���L�2��HF�e�����o�~�I<)���;g�	9 �iȘ:D�]�<�U �G<��$UlXb��XF�m] Zä8�)��\� P��aP?z0A��[	A�B�I�)�T�c�֪�0�sK�2���䍘Y>�S8,AD�Ǧ�:�����97��d1TvGζH�m`0$�;��ycf#�dp����Ťg��L�`��{�(����a�az�L?
f�O�e��g�^��"���jS�4ڠ"O�l�^�G���E
?G����DT�<@���{���'�k�f�Y2&E�$�i��յ�ycP#g�a����%&%��˞�}2�Ћ��<aUa�#S��3��5�{Pw�<y�i�)v\i��M�:K�V�p Z�<��c�VX�)�5T4���T�<vNf�A�ɰn8:qtcP�<�'nTL�Q؂	��v�Z��e$�Q�<�hΒ8F�D���	~B�XJu��W�<a��8|�0�8��w�:�BV M�<�FI�B��aB��tC�Uja�a�<���K�>��u�q*�)l��Ka��Z�<��n��a�P���)|]؜�e��M�<i���E>D<�2l�?��m�/]f�<�f��m���PT'W=9��*��k�<�" ����㦊F"28k�z�<��Ή"l(Z]Z���t��b�w�<���ɬj�J3�9ݐ=�4GH�<��j1>�=("�K�lp�KG�<9�n��H̰�O���kf$�A�<����/z�����1+e����}�<�	Y*�6�����6�5I�V�<�3	��Cp�(�Qۿ/���(�Sk�<���X�U��@�YW<��rN�~�<!�AM]wx��	ĨT
2`�R�<� ��Rqe¶��CN���@"O�0���1x &J��ڱ��"O�=X�`_�$H�+P��8�"O@iKw	D+;�4x�@
</�(YIp"O�A�C�9-�� 8!���
�+"Ob�aT@;ϐ9�s���P����"O��ʧBI+<DCU�MO$��b"O�q2�o��jH6 ۝`j�*�"O�z���7$��LcD��\	�V"O�!�!C t���⑳b$��"O&�y��#P�9���4���T"Oʄ��Q� Hs�Q&#�Ll"O�ؒb�]/P��h&1�B��"O��ɀ�j$l����A�Z�t"O"�9���/�M���F�c�$ٗ"O���0�!;I��3uJ�?]����"O���,��iX~���)8�Б"O��вj�R�(!⇇9H�3 "Oڌ�D��_�
��Vƅ��V<�7"Op�j�(I�!}�*%�B$l&�T��"O�����������l yط"O�xv- �m�ff�"'ŲW"O�$P����{F� ��Ä!�X�`"OdBv������^, r8f"O.L	��T��~�."Vv�XPS"O�X���2I�z�C7	b�|*�"OJ�X�dZ,b�:	ԍ� F�ѩ�"Ozi����^��iSmG�	���"O�ԙuj��V�t a��_&��3�"O�-��%:~�bq�T1<6f�"O�!��wY�Ͱ%'K�Zq�hK"O���A ��_���FT ��<��"O�Pj���.|R9�ৌӲ��`"O�AKv揯
����V#�VQ8a[r"Of����
�3�蹐���qW�<(�"Oڄ�F�msX����N���"O8E��O�\4R��,N����"Oj9�E�V��$�����<a�"OJ�J��}�	�0-�=˰�
f"O89�!��"3�]��T1cĜ�"O@�!��2G��H�6�\�$�:|��"O��1��ʑ<J�b�G�mf��@"O>L���DJP�5O̹\t� "O44��j՛X��1��eS�+L���"O����У2�)�r��3i����C
5:C�|����#Eȶ�b��ķH�l(0�$D�����*2�$����>~��9�RDl��trf�x:��ߓFu�u����:����۔Z�\��I,~0p��FEֵR�m�м3���rx����0��B�ɉPF�Т�努W��}��I�$��XI��y�Z�r��U�O�Z�O��Zae�S�^�C�'�P�C�1a�.is�i
~~i�S�D#?��8+���<���/�gy2$M$sn4E�D�0J�����#�5�yꄃ_�|�\�}�����Դn�J,��!40���J/lO� �"2!-��B�t�|����'�4�Ӑ�(� e"�i�E@�D�<���R�Ϗ�xthQ��'P����Uqm�4�]8dR�h�{®�6#v���`�=u��>Us�T�y�@i�$�'���	sm/D��y�.;|�� G�8����Am��̬��I� ��5�(���n`���AbĄp���0�W��dC�ɺR�p%�B�Km$�@�/P�*�6��*�D� )��=9��ȹ{�`|r����en��a�c�u��LH�f�W;�]�E��;�̐;T� 4�����4��Q�҄��"m�3&��й��S�? 1xu/4SNA�S.�
J8T2�'F��R���;�ɧ�����5(]��Hh2��21x:`�a9D�� �
�*Or]P҃ϓf<�%�G�>��k�y� �!1<O]i!��8x�ޠ�`�=�!���'c�3���DPVܠ�OW'b>43�N_�h���x�FU{�!�D�2klj� �/� a�=�Q��qM0	aD*���z�' ���&�[�yԚI�eN��c�v���*%�\��!�1,�%��[�:�P�rb�=�(� ��3N��)�������|O ��oE -��f%D���/�y�|�xD�G�z��奟����Š-0�Up�˟~X�����M���1#΅�anH3��5�ON���M�Q<���' L�HEUP3�����dM-&A��'��E�M�./���ꓨ��u1��X`��m�#�,,��b?��e�K�.Z$l2��Ϡ?���ӌ(D� �# �'�Y�L�޸Ã��< X�I⁎���2(O?�d�$^�ZH���=/h؅¯+A�!�d�ML�����3[DR�F������r��3i6�y2A�+"��L���<(M����W#��>����#u��*"�ώ&;����!��3%���y�݁<PA�JO�:�`D��y�D�}��A����To(Q5�ז�yrO�z����� e�P�e��y�I�o }�����d�+u�;�y"nI;K���*e"	��,�ٔl��Px��� ,n���;)D�Z����F�Fi⢆�Z����R�'A�"D[�e��}KD_N8�DXÓ ��9�o�"`��d����%
EU*�X��j�nc1s��*D�C�D	kT$8���-t*��5+,-B��ΟJ{pp�#IX'K��#������V���Ի1<�#׫�	=Aڕ��0>�Q��/F�(�i3J��i��]0� pp� �T*Y�Ne��_�������X����շk���g�~�hHtmG�U����F��$X�A�OtM�͌'I(����o�����p�����IJ�z,�b�a�T��RеG�<��F�ʓL*�p���)�����ʾtȅ)T#
#>YkAn��0� �ʅX�R���t���Oȴh�E�U $(a3ю����N�c=Z�⥈\H��:��8���34U���@L(����-�:�|;Nߑ�8u�2k^�K��3ǳ#��%�@,�ǟܐdm;�d kb�_�|2fNI�.��pqGˈ~�4[GUV�'_�\�cmE)%���Q^��+e��?ݪ}��"T9/�tʦ�I<Rm�S�[.ҢΦhP�qѤ#T=��3�	.Hzh�iH����@VF5˓ �DL(P��Zx� ���$Pz2H���)��,NthB�� 8��|@��C�7�dq�q�S�w�ȹ�HK�V<��D�i�����VS�� �jݠfqn�ѶHσk�~�`*Kf��=:f7��ؖHQ��(iV
\#�~R����*a-^�M>������?	m��^գ�K�$���	��O��je;GmԿY�>9s��s���j0LV6r�D˓sfȥ�c�A0X���(y�����K2N#����i��s���?��"-t�,�G�'{����f�^�}ڰ�2(�o��E�PE�4 s��R�M�A(<� ѭI�Z
�KM(hJ\Q1c�Ojy"hD/6��5A�́?�|	Xd+��W�F��~���:.7�����B�����.�Y�<�����P1K�N:b2n�䈂���b0f��U�g�v�
��JG�	�X��ԡ�� ��D��F���W���r����tm��u)*�XBh�,x�jC�	2R���c�m�#�-{'&S6�C�ɭ7�P���G:]��A����8n�C�2fĥ)v��;;jN���K!r԰B�	0,d 8 F%ܫc����6��1bZTB�	(W*�ѐ�B�P݌�7k�*d��C�I.yJ�A� �JPE���ğIcC䉐-�*X(�g@�%�6U��4��B��?��Ѣ�����R�^	��B�	%m4p�)���>c�ؑq�݁�LC��(K����!9?,�ZH��SdC�	1J��1+�1jw�\R�o���hC�	 �x���"�I��
�L�!��B�	�Z��2Gm�aF<4���=J�$B�I�c~X܃�Lz�B�b�
�W'6B�I�o=9᥎��t�K�
G���C�)� 6<iP��w|C鈷T5��i�"O���r�\7�6p8!)[=s86�Q%"O�áN�*,�T�ƏYC��"O�|+��R�RwH�QZ�C��c�"O\I	bR�&�6%���04�11"O"�b0��P��X�kǂB�]��)�)*�����O�]��j@v��Тi�!?��e��"O���Z�,�j	@�b��w��p�0O����V($���Z*�HػP%��PLjR&D�1��{bA��%bL�(3���8�i�<2�(�W��0u�Ҹ��g%D�����0f䮡`�����p� �ɗ@>90�,s��Ɂ?1^-��K"8�$�Q�N�j�!�ě�EBm��˾(S��Fb�:?��D�Յ(Z��Oz�}����X�`��r~�0u�I	O��ȓ,�f�{ЦاK�9x���d��I;j�M�tAXE�a{�lS�z�P-c�ρ���d�` ����=�`o�	
��P�,sӔ��U��U��ÕB?M�q�V"O��`�f#~}�3=�2��`�dY�0�A	�H��s0$	�bĥ�e���N�І"O>�
�HG?PN]�&b�y����C��z�P��U�$6�g?�5k�����Z����A�2x��Ke�<YINX�hbƭ��-�����<���ϧd����
�i�P��r( Z��X����*shh���>�ı�1O�!"�F��������R"Oz|� �V2Gw��1fɎ~�4� "O:\�C�O�d���5�[���`��"O>m���\�̚�(�Ă�1�9 S"Ofqha?[p4��"�{7dRR"OFMSEiӌ+��Țt��1A=��;�"O�����^3-��p�p@�+�0��F"O^���f��"q����Mѧ�y*�"O~�*Z
Ep� eW&H��"OF$ꃆ��06`�� �:_�& h�"Oʹ�ѡܳ]��8�.,[L��#"Ov��?�D�1e�<&1�q�"O C��B.�s���%_ͬ��"O�A�"n�.��i��54�V�I�"O�T��>�nܰSLGL �"O:ѓ�)P�i^Q��ɍ�9�v*�"O�`{S[�16��bF?����"O��8�J�6LH���	 �Ȁ:2"O��@�E6���g�݃/�jl��"O`Ĩ!��114������}��,h�"O���RP�*��)�!u�L�t"O�m�F̎0n<�uf�{kZ �"OvŻc�V6�\{f�����2W"O���M�>q�Y�b�ђ!�<��a"O(Xf�J9h��5�:�,3"O�5�u�	j�V)���)&:P%"O��`pfıE4dx���kϖ��&"O���dA�7���2�]0(�\�1w"O��v�h��Ѓ'#U��ҕ� "O�E��I�<{�)"U/-�TLs`"OP {���j��  `��Fp�9�"O,=�ׂϘ9�8xiW�@Bur���"O�d'��	ؖ�rP?Hij�b6"O�i�ᡃkW���2Ͷ��G"O�P	�N��N�t�q�W�I��h`"Of R��	�&z�	3��F�{�
��"O�aV�ɢ��PH� ���K�"O�E2CJW�>�xm���.Gw��"O����Fބ/���UIֲ1s\i��"O \ʔ	
^�n�CRj�j1"O�L��C"|��L��C�3Rnu�1"O� ,��i�=u�Z��B�=xZ*}H�"Ov���L��58ș�ƇoO>=�2"O��3T�Ќ5>J�#�)/%<���"O��aj��	�Ti�ǈȖN��<�"Od	b7�L,p"��ѧ�ܕtz �W"O�yђM�����c���+j�X�"O�����^&�`c��x0N�q@"O�5��B��Q< �Z&�ӅM"d�Z"O����+��\ǨtzV��/'*ijs"O��J�T�2'����^�!�xz1"O���̊�	�h�q���/P6Y�"O6aS1�Nm�&qw
ߑA\ђc"O2���:FܱahD�L0��"OMR��=k�܊6�J�j�v@�"O8M��,�p�5��E��"ɸ�"O�H���D�Ei�JG�.�be+Q"O���A�oi��e�N��`�
6"O�D��Ò��8I�C� eT	��"O�e����4��PbDl�sEnYbv"O�u�	O0Cz�|�%��'J�	(V"OH���[�m;��h�%L�Y8lЪ�"O�,!e��\����Ć/GZɹ"O�܈2��F�t�R�#;.��a�"O���!I��u�8���ßg/����"O��9� �\�L��O�)+,a "O� �p�p)H7I�m �:�"Ol2�GG�^2�Є�G���HC"O�lJ��I�8¬43���i����&�&$~���
�s~�$��(���Ӗ-&��8�]�䬐��ϱ:��i�r��c;���-O�<�O|"47O���Ov��D拪+�&|+td
>�&��AOe���')� �D�?��Ģ��Xv�k�c��)r�����ZA�u���s>	S'�D<5@����=d�nuѶK3}2iC#{ɠ��Mצ��H����Q3@�4�����B��@�O����G��T�>%?�'B$�F0f�1q�%D>?�$�b�4D��� �⌵&o���/O�?��R�A;��u��ػ^��<���/+d��`
����L&�)"ҧ`��M2Ԍ��+$ ��P-�;T�ulZ9I��$�O�����O��sӘ�6��(�VA��d���B��i�Y���(�TO�?�R��<�H�if��4j�B��J�+��I�s�$�ĕU>��QlY�G�- �G�����I��Ĕc�ā�i*�Zȹ��Nܪòh;H�x��V���5�p$��A�Z>FL��Ș���� <`���]�a��䜶n�#�H�a�+�kq�Qf"�"�4�HDK���y_�e'�(�Ak�D���çU�4�7.Ջ~�@U�擄jF�Xe 	3~�P���* m�)�' �~���Z��n�{���;
{L���ǘo��a�Y��9��OlZ��ԃ�u�x8�S��r�Y��'����d #y�{�&�
k��m �'�
q���[�Oʨ=a�� �f!j��
�'�F�j%�-�h���IQ�Q���y�'�" Z&�[?x@C�g�'z)�s�'�,���U�7�|\�L]/R�y�'y�4�"kCo6z�;�NM����'/���W����dAfE�0,��'jvP�,�0s�0qq��N�e8^H8�'�R��0}�~��g�ۼJ�p��'�: �%f�58<�a�O�T���r�'�����Ί�U�=Y�D�����'>��.�`�h�ɽ>��4Z	�'��ٙ��9��13��	8;���'�^0 �@�#����࡜8-��U*�'E�bH.)WΠ1�	�8M>��'gx�	Gn̶$V�i������Y�'�&t���͞E���dIΠ��A��'�,���ZFU:X��!̄����
�'On j$*!%4չ�N�LPҼ��� �� ��� _��*P�9{����"OP��3��Y�Z��f�U	z�� 0"OzM�4D��?8<�\T��*�"O��k6��`�MBc�ͅPJ�D�"OJq)��;=���/;p,�X�"O�!��7~hi3�n �yH�"Or�C� I����S.D�i�l��"O��Cfj�9_,ez��j�>���"O�jE��o�V�C�
K>�zS"O�ሃdȆ?��8�䘍Q��-i!"OBD���ߤP1��aj�-,~�HÓ"O޹�t�D>g����:zk�(0"O �2�Һ�&�P�oMV4|��"O�PD'ؒo�`@	�n��80�Z"O��B��Zm|x�!��#Н�"ORE�U�ћ1�ތ��J̲�6���"O"���h��k���:�L 5R���"O�A���w�A*�o=�0��"Odl�4`I}
��
��y(Z0��"O�1ˆ��`�����B	h22�z "OD�cu�ځ-��4 0aґJ<`�"OnY�D�/�V��בr
:D�`"O��X��\�	�ҁ���(p   �"O�-[`�݅a��2�J氨s"O���6��*c_��p5J�)���P"O����9�l q0jv]P�"O�5A��$JO�Iqc�!dZ���0"O�1¶Ҷbg�,��A�$\I�\ˤ"OD0�A�S��� ���]5��z�"O"ic�I�1 �Y�,�,�m�B"O���X�M��i��i�3av�4xf"O
����;@ob���G /l\ր��"O� *�d�Y��F���<��mQS"O��V$Z*��B���v@J�"O��!�Oӗr��������l3va� "O����Kb� @�ŉ�%yJ�� "O�,�PI����HՉ�EbXQ��"Oĭ�f/�6{��5s�Yd)N;�"O�|s�RI�R�P0A"��"OJ�9�&��P��4"Q�+ x3G"O�}k`�R�RU*�!�;���#Q"O�=�dC	_PT	S%;4����"O�$���١l
�%2�̿A&U��"O*d¶�Q3Ҕ�"`�>&�=IP"O�I{G�3�q��;! ��r�"Or��GHV:��B�Ǻ'��A�"O��5I8e�Z�3��~�,\�"Ol�� ���
\z���9���	�"O��!�ǹs�>�9w�H^J�Ū'"O��@ĳo#ؼ@�
^C�$��"O��b0�W;��p��w}.(�D"O@��"�ɒr��!��3_Z�M�C"O�`Y0�%[{����$o���Q@.D�p1��СM�|�a�C��b3����/D����A� Űg�B�I��{%c9D����ə!H/`��pg
$�DYa��8D�\ڳLE^
�|�tF�"E��
�*"D�d�2���7��$� )U����("D��Q�]?j!�WD"j�%x�.D���cc��h���Ui����d+��,D���gC�+y�4SA�v�[$,D� 0%ɟYApD���٭Bt2}�s/=D���5*�qy�Ī��53���*Ӂ(D�x�5��lp�MyЇ0M �ZW�8D�� ʥj���Eo.�s�%J�8<�"O<x���1"�aA�
��9��qpq"Oa�C˝�o�FD+�AR�"ܣ�"O��3�.N�Qp��� 6.$Ч"O>��lO�@���6 H��)�"O}6�Ia
��!��/�JA��"O�\�kɡkG��2ӦɴCKb�{s"O2]V���L���$UK��I "O�Ƅ�F������;e��}D"O��1�M5�*�Ǥ[m*]��"O>�h�ص?�X�9���!-x��h�"Of,I��@h����#-\L\��"O$��`�%E�@;��уpH�D�!"On,�UhZ�kC��H�ƕ�n6��"O�Hq ��;s,���E��k$�j�"O��[dC�ݠ,!�@\��r�"O�2$��eI���p�T�$��QCC"O��ҳ��*�͚wɔ�d4�<j�"O,�ZN*ea^a�����=��Q�"O�t�S�vyf��牖�{�V�C"OPPЇ��H���R/�v��"O�z���^�)�w�ǀf'��
"O�
�H*���c�b	z2��@"O�u!$��!g<���G��t��e"O��(T ^�t����o͉1��h�"O ̣��,�8$N׭&�H��t"O~��$E�-+��K��_�?�	��"O"�8�)�)8a�b7�΃p:�Q""O*�C�A�=�48�D�;B� �"Ox�J�B�2
�N����t��YC"OƐ�W?(@>\Z�ޤ�l��y�F�h�!�ԋYC:84
@�y���4?������W�MCS悫�yr	C�$��˴c����]��윸�y��'�d(���^��uz�ꇝ!�D�P��i�W��]Z~�(�	�!�$߂ �����D�##Q@��)_!�G�,U�]"t�D��l��EJ��T!�Q!���`ĩ��L�Ԥ�b.9�!�dڈ&)Hsҏ-I���;�&{�!�ː֘0r f�n&�%#�OD�!�$S$+��P��V�F|�5P�Ͽ8�!�$ƬJu��k���Q[��pD��9m�!�$�-�p] �HDZ��!��bH~P۳f�P1��8P  pg!��= 8ᓆ!�2� �R�"k!�$Z�f�%�N�g����Q��@	!�$���Ȅ�FªP�\�s&��76#!�$F�4�\[�ז����ԇS�!�$A�gL	�Iܩ/������G�{�!�ė
o&��s,h{��)b��!�d��S�F�b��`���d!�K����#jO���\�� �>y�!�Ě�O4�m�$u��hT
Ǭ$�!�H;Z�(�:�eA�-k���ܞ-�!���o���@T�oL�k� 
xq!��"Y��	�#��7����,f!�D5��q��D�H6�%�GW�N[!���5Wx�
�J1?lH�e�V!�V�'fڕ�,�=sPt��n�,�!�ǼD9,�AnR�7���g�>�!�Dڅ8-A
�Y�B��%��x�!�$�?j��I+���L�$�� �ݘfp!��ҺH>���C/z��ɕ�_k!�� ����ՆOJH�A���<OL �"OXZ�؍+�5�&T�#(���"O��z�`
�~#D�#�$�`¬�z "O�L�a��Ǣ<�g��d�ޙ
%"Oĵ�G����P�9�00��q��"O�hc6/�?1����J�Y�҅2�"Op]��/�0���#c)˶ELt�s"O8����ԉ|{b `��V�9S��Z�'�R���F��T�:Q1'L��$e(�
�'Y��z�/V!p�NT��hZ�!���'�DEbwV�4�H0��♺D�RD��'�����\�s�L���H� Dz�'��bQ,ע��1Q���x���x�'�h��(B���F�C��h0�'�6��REf���g/�k>��'��Ŋ϶D�� ���ҁw��@	�'���Ԃ	גYQ��Y/��T��'���Q�+=a��X�.W�+n��
�'Z�|sDf��s��hß.r*�	
�'�~��#ڸ57Fp��#� dR�X��'�%�&#�:27��S��_S�-��'O���n]��@j�!Ef)�"O>͋G�Dm�i��dM!p����'"OFL@�b�=B�`��f�� ~^�&"OLuHP�0���$Y�\�k�'r
����փ
�����(�	�'H�ܨ��E�#g8(Q�Mc�����'���-ـ_�Ѻc$mӪ��"O���ӥT6����D�{��("O�X��-Y�I����E�W� �H"O���a��C�4,ӃN�a��(u"O�(�@*�C'��z�L�HW�H��"O:�p�(U;nJzQ�֯�14Z�=�T"O�P����43�p:��/X����"OH�OH?CF�@9��O�VT. PS"O��s`�>U�ԣf�\�B�� �"O,�Su��=+̪�@�S��3!"OX���4p�T�Au 8Z͈�"O��aLQ�V�tYqM�=��R"OJ��K)�6Y!q��|�
1@�"O �I�P0H ,8;�Ӑ:S:M�"Oν0EN������^T�8��"O���A�'&!����i�9m`U"O�,�Ge�vH�����^�PȆ"O��Rg㗭����x�$�u"Oɱ֢�'H�4A�c�����"O"�A� �5 �*AH�ݖO���A�"O�I��͛hNx���K?���6"On]c�	   ��     K  �    +  �6  �B  N  ^Z  -f  �q  4}  e�  O�  ��  �  ׵  x�  ��  ��  !�  q�  ��  ��  ;�  ��  <�  �  : � ; � "! s' �- 4 ; �A H sR <\ b �k �t | B� �� S�  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O��jg�=Pz�Aa`�#�h��!\��̇��#=B8#���fB8%pS��H�����fȉ'�$!q!c�	^+F b�ǂ!3�v|��'��EK%�ݵXF|ԲBER�/�f�ٌ��#�
ّ���5�`��'c�6vH��C$"Ox}e��N&}A�A�3Z`X�"OJi1�Hճ,U��I�	� 4Ft��"O�D�tkI:��͠�(A�Iddi��eOuH<YS@҂+2��p�T�w޵����h��\�>y���BdlcL
�g?x<����d�<7�5�)�늁yD	�`��J�<�"]2����ܿf:����G�q�<I&��d�ɓq�:Ρ����X�<񥮀�8TΩ���y\^P3�N_�<	BdJcV�����P2.�"�J�,�v�<i��1i��#P��,+=hR ]q�<���	4M\���#���:�����o�<i���3ZJ���5Y�%ԞU��g	h�<i�-
�Z����&��U@�ɱF�DM�<����+�|�h�O��i�ʤY�h�K�<����u�
� R?
Kv ça�<���.-���4��*��ZVŀY�<��ꈍ[����Se��e:��Q�<�%��$f��F�S�r��TeXX�<��(g��K�GįDlz�iU��P�<�w(]�>c�r!�*8`9K�"O���T�W���!G�Q�R-�"OHXB�X( �i#B��)^i"O"5K!h�5��В��+B
p�Ia"O��Y�Xr�-���,�ِQ"O���j�"�U��-�~��"O&���Ǚ7�l��t,�V (�"O�a 2]`��:G���ya]�&"O2K��ƹEέ�F�� F��QS"O�%�⋖�s�J�y"nԵ'��ۣ"O�Yk��z��i�`�@�p��"ODY�̙<RE��NK�l/2!��"OJ�jv�۽;�P;"�̼#j�P"O\I�/���Y�	I����q"O�D�$j�4F  �H1e��N@b�"O� ��
�/q:��W� �!��Ժ"O깚��
=%dU�f��3���7"Oba�6� "j0]H"�sΑJ�"O촁LTf�䍐ANL�r�4 T"O�LU�]�FP���2�xX�!"Ou���]�9��]ao��)��"O
�H3 ��Y��Qo�)I����"O�u�wƓ-r��@�7c��_���"Oz9T�ȧ&u�h�IK��< D"O��!�5�6���\�f�"�"O��k�eK-fCu����:���ar"O� >��sc���5S��	�C"O���I�8-��4�nO�G���"O��X �].8pw�R�u|�#"Ob�[h>S`�b��C"4]��!"O"-���[T�]!u�v%���Ĉ�?����?!��?����?1���?����?�C��J$d�bbT*v B��?���?���?��?���?y���?ٱ@�&i��(^@i���ز�?���?9��?���?��?����?i�f�	2J�x+�QEr�5����?���?���?���?���?���?���)rev\IQo�Z��=��2�?���?y���?y��?���?���?�� A�7{��9��+X,�ᑓ�?���?y��?����?���?I���?�jȍaBN��3�N����S��?����?���?Q���?����?����?��BL�`\��ߑ�v +p.���?���?Y��?���?)��?y���?��ᖚ͜�C�\�mHP�$�?���?��?����?Q���?y��?�U΋�@�Bi@rdݭn�����A��?���?1���?���?y���?����?���<��� ���m�BE�CG��?1���?���?����?����?����?AR ��d ʽ��  T�6��'f�+�?���?����?Y���?)��?���?�֋Z.1P�u�#PR��a���?����?����?���?��dQ�6�'
RgE/\\PC񋄇6\v�{�eN"�Tʓ�?�)O1�����M����]xb�� B�av@ ��ŕ�P8%�'2�6m&�i>�I��q���S� @p�f5�T���K�����	3�Pm�[~?�ڱ�S}��[�#�d�b��-�,��`�1O.�D�<���IĆz#B-��N�:%��y�D��b�&�lZU'�c������y�ǔ���1��D	7�����J ?2�'I�Ĭ>�|B�E���M#�']
��s�R�F�>e�㣕�m���'�����6�i>q�	�9k& �`��a�����+t�J�IByғ|��w�|�kv��n�����Nd18��U&���p��O���O6�|"�Z6D��ؠ�TU�#����Ot�����G�1�t���G�J�$�(w��x� $�<{�v=j���� ����O?��6fH�ً���y\�a����Z�牱�M�&��u~��yӎ��Ӱe�p,�'e�Np����42���ҟ���� Ӣ�
����'��i��?-��"M�SD�K�D�2T��h��?3*�'�i>)��ڟ<��ٟ��	G�9c��*H6��A�F�]��P�'�\7�g4����O��D4�9O�)��L�e�=�"�Hqǀ�<����?�ش2r��T�O!�t�ϸ!.�
�A�:_�:ӎ�) ��R��By�l�3��� AC�8/�Ɵx�!dʓ2�r��M�v�"$�O(
�����?���?���|�)OFqm�)z�r��	!��s�=|�j
�NC D�J��?�M����>9��i�7��O�uʒ V��q��o��5@�iM4x7�v�l�CԦ\8E��$A.�i�	�?Mj �S���nϨ{���h�A]�n���H��d����ȟ���˟ �I���Jg�̊&\�c��NF��5JE)��?A��?��i1���^���۴��S��2��	�0"cnL�c��b�yB�i�,6-�O���eӐ������ך���b�	B�+��@b��)r".ͱ��'� Ȕ'��7��<���?q���?��M��A�}p��Q�:�.L�֪���?	������ l�ȟ��IޟH�OpA������,ѢJ�j��ON<�'In7����%���?�8�h&�,5�N$yn�`C��3�I��N�?hl�'}�֝����dy��wa~����Co��!J�@ ̀��'?b�'���O��	��M#`o�S�k �%a�AXa��j*�+-O|�oZJ�g��	�MK�/M�vK6��T��:}#�< �B�I����'.��Y��iK�$�O�-	 ��1���@�<!��8]jV�����;��=@pE����[���	ğ��	�d��ϟ�Oz`%
C��t�<�:�"V�l|J��q�8����O^��O����|�4��w�����:V�\E�6	]�OS&�z"�O�6m<���I�O��6Mb��jP�sG4�"�J�d��#���I?��X#�'N��'P�6M�<a���?q1�����PCP�����K��?1��?������F�J��O�|���|*�I�q���kH-��2dK�C��$��	���o�L�ɞW���Ԧz�\8Zӈ$���I�h�7�Ŋ(.��AB�ULy��~�͐��'�X��I�F7d]1`H�U����T�G�=�e��Ɵ �	���Ic�O�R �OOz$��jS*�3��I�:��Z�Wo�I=�M��wLz���
(a7z�:�E��@J��'T���g���U6�c����q�"x1�O��̉�l�AP���tL�&N9FE�&l
Ny�s�:˓�?��?!���?��?*�6�o�Ā���ܫMr�)Oܙn;�\e��̟<�	w�s��kT���W[�����K��� �������ĝ䦅iٴ���|r�'�?Y _�(��G�;�dܡ��D�+���Ӈ!Q��򤖺_u��k�Fy��X뛖T���r΂;`��t�M0�݉�E[����ܟ��	ϟ�|yb�k��5K���OBl�&i��/�6	�/�9'� 0t6O�Qn�f����I �M���i*��⠴IQ�$���0��,ɶ8�q�im��ݜ�`�����B��e���MA[N�� �s� m��0⡈S)~v�h��4Ox�D�O����O����O�?]�it,��M�	�E�WcT՟����l�ش�Ĉ�*O��l�E�I|��@ o��Y.f���XZ���%��[ٴ@���Om3E�i��)L|��Scg�L �0��7	;\Y��j�0L��i�ЛÂ�'���'@"�'J��'�@e���R�fR�y��#R��S��'�Q��j�4�d����?9������C$�r��#|6݉ jH�W����'���w��v�a�T�O�"^�������T�k��C$
9�U��1�@}h���oyb�w�}��'����y��Y�><4
TD�[D��	�'���'B�'�bc�<����<�'��Zj��Mz<��'�[�7AYʅ�;]^�ʓ;�6�'��'�r�䛶�ͣ��D9��/'N�`�,̯e+�6��O�p��`ӎ�H\L�xd��r,OHx�#�F��Y #�������K�צ	�'�'h��'�2�'	哵u}B��j�.T�P$	���3����4_\����?���:.��A٦��:pz��%o\�;M���7�ˑu$�q����M+�yJ~R�"�M�',h�ٕ�-`��9  ��$#*���'��FPޟ�H"V���4��d�O���ۓ¼�����&�A�h�8���O���O4˓Z��G�����'��$� Y��L�I9���C�]Vk��|Bͽ<����M�I>�7��p&�d��I�����u�x~bMS�B|2����H)R�剷�u�E�ݟ�"�'F�ԁ߳~��HsǗ (`�4�'^"�'4"�'Z�>�]�q�Q�w�5Y ���Ь��5�����M�U�
��$Q����	m�i�iA,�J�2D ��;�4q@�H��tnڐ�M���q��ܴ�y�'q����c��?u˔-W<lN%d�݃x�\q��Ԇ��	6�M�+O2���O6���O���O
�3r�U-��9���L�q��L��B�<��i&����'F2�'���y���;x��s'��g�9g�@�wz*˓�?��4�����'�?���$�"�s���SV(�N=�V4 ��.��Dѻj��;��H���B�vP�3cƠV�j-!��:��b׀���'�R�'k�O��	��M[1�
�?	�F�CX�(ŅVyH0����<ѣ�i�R�|��<����M+�SS܄+�`Ʃ~n�^ x���R	�9�M�'��,B�{������S���1�u'�w�r�8Aj\G��hs���0�
��'�r�'K"�'���'��e���#=<� �g�^�R/D���.�O����O�MoڤJA�-�'�7��O$�*܌�wJ��tOT��ˊU=��aH>	C�ijj6=�@1"��t���*2��D% H�q�k�o�d�{�`��]W*������$¦��'N�'��'̒�Ӑ`@4T���C�m���P"�'6�W�Hr�4K�m��?i����	݈)��黦D	f2kMPX��Ot)�'�p6�̦�'����?�	&�@��)��
� �L�;�NQ� ���R��#a�"��	=2�����q�\�����k�A�A�XiS��E?v�>q *��?a���?���?�|�.O��l��8x��������ѓc,���3?��iI�OLL�'�6m(	�q�4��Q�Lsf_(Z�n�|ʑm�ݦ�̓�?	���!�V���Y~2���rD�۲�M>R�0�d��6m�<����?����?Y���?�+� ѐ�K?/��p@1�fK����/�¦� %�s�L��� &?牍�M�;d��ͨ�IȌb��6k��@��i547�9�4�N���O��@�goӊ�	$��SP�Z�&�(2"�9a*��I������',���'�6��<�'�?�����4��%���B	V��?���?A���d�5j��2?�����:A�x\�8�e�%��Mj��k�>9%�iq6�)�d��6�2�H�U�6��(ՙ=;��O6�r�ƈ@�����,B_wD$�ɞ?rb޹h�t�ȴ@�ԆhcՅǨ2��'B�'`r�ȟ؀��D5x¡��\������ϟ��ݴ&e�5�'Ƥ7�7�i�u�P��^m	��M�eki��㶟�n�M[�GV\�s�4�y��'���t/��?i⠥��2��	��� /T����JRS[�I��M�*O�i�O����O:���O.b��V�G7]R'f�!i��C��<���i��A�'���'���y�K����M߮{6@}ځj��FJ0�M��fgt�F�O�I�����= ����e��#`p�A����8@*E�s��k�I�M%��$�'�0��'z47�<��2&L�\#�K7.xޜ�ũ��?��?��?�'��D�Ѧ���i���`)�&2��d����32�>f��1�4��'���'`�6�|����$	��P⑬�.6@��1`N'NuN�0/f��:�˔�I�4�~"ù���NYIe�	��S%.��yj���OF���Ob�d�O���5���vx(�E�^�~��,�bϛ�#�������I?�MӦ��}~�����Ob�YP�X(MT����B�S����UO'���ŦѪ۴�?Y�n��M[�'�b�"h�d	ԈX%M�4R�nWZX�!��Nԟh��^�<1޴��4�����O��䚂6��h��' l���kQj��kG��$�Ox�YT��J��y��'��X>u ��V2*��}���_�V�E@%?�q}��tӺ�l�p�i>���y�*�ce�� [ K0hW�:�0���o�^Q�E�*?�"���|���T�˓��[�"�9ʂ�I �qeb�*⧟?�?i��?���?�|r.Ot\l�
�;�MO~��A�s��bD�Aqy� lӨ���OdhnZ�5o`�cWl�,FD�O�"�~Y��4P���f6O|�	#\�J�(�"�վw"��$��� �-�cg�^ۜy�gA��hĴit栗'+��'�b�'�R�'h�'@�N�eT�ٵꋄp.x4q�48Yٹ���?������<7��y�
�����D@'v�Za����6�ԦXK<�'�"�' 8zy"ܴ�y�˞(*h$�Ө�r��t�6(ъ�yҢF(:�`e�� k��I�Ms-O����O��2�
�A�ЍA�(�+�K�OR���Od�d�<�d�i��0��'
b�'@BM��`5���.V���2��'!�'y�˓�?�޴r�'�Sǀ�p�^yhw"_+pY<屚'2镍wRܨ5��	W��.�u'gM���p�'��ez��:jn 9*�g�N8��z5�'[�'\r�'��>��2[���,��'�ܭQcȖ�I��	&�M�ܻ��d�ɦM�?ͻ<T�%�,E�4XN����Vg�&`�̛��k��oZ6:�\�lZs~�ݧ'�.q�S�D��G�8W�X�cꍸi�R`DU�jٴ���O���O���O���:�
��	�qNV8���
"�VʓLe�6��L>��'	���'ʄ0��Z)�!B�������<9���Mc��|J~Q��!��A��fR�H���` �
#�(��i��$�ph����~Th˓�vS�����@�8k����_K��Z�kZџ�����������Dy)p��IZ'�O�!	�ϭA�����J�t�U�F;O�n_��8��I�M+ŵi˒6�C�<�����b�ZX�4@V"IPry�akh���ΟJ�Kʸ:����Gby�
q���Q�`�R�V�5Þ�P���!0��I柤�Iȟ(�	۟��I^��XF��IX���`�ƒQ�m����?y�؛���7-���4�MI>�w�>W���S ��!y&�L�zV�'�R6M����� $čl�g~��
#�T� �8����!�Z"�t䪴��֟0�C_����4���Of���O����'0���b��.3h(A�EI�&����O<ʓ=כV
 ����'8�T>��Æ�&�)��Fؼ7֞L!V�:?��]�8�	ݦ�hJ>���?�gQ��xW�]((~�H�"�p��X��^�wKV��'f��]'2ReKyb�w����D�E��@+"��E4n��4�'���'�b�O����Mk�B�)CP6��ߊ$H>��'ϩr�Ҝ",Oj)m�_��"H�I�Ic#�\+*�T�Q� W�����8�M�T�iJkG�i��D�OBUq�"ɫ����<Q��$-	�
�5�<��RE���R����ݟ���ٟT�Iٟ<�O
F��&��N� yȀ��C!6I���cӜ|��9O���O���$Z��]�$�mޓu������UX�41A�FD=��J�"6�w��#$���r�l8����-x����$�|��+g�)K1��	K��hy�O�� H�6�-Q�9�"(��A��?���?Q)O��n���	ʟ(��#?QL���O& <I�F�q�)�?1^� �ݴ\��i;�D� �`���E1�X�:�Fį+�I1$6�q�6��_
�b>���'����<!X��A���f��!b�G�]�����П���H�Ip��y�E,B�Vb�#�H�v���D٧QW��rӐ�p���B�4�?IN>�;|�0H��E	�i��$JS�ۇP���kX�6�r�b�mڜ<ln��<���2ty`��.Hಌ�'M�0m1t�מ��	�BJ��䓙�4����O����O6��, �M�'�yuJ�sE�s��L����2���'�����'1rD�2n�7���z����`	�S����4f�f�7�4�6���:��A�.D�xqA�ƴ�X1t
 b`�����<a`��)3��� �����G��%K����N�A$�
Ae���O`�D�O��4�d˓UM�fŞ,2=2 �Z���ڭ5�&h)��	��yr�q�|�`�O�HlZ2�M��i��|�q� ..�H���χ�4��a,�/R��1O���^" a���^\$����;S]�L(`C抍SU@к3����?���?��?����O1���<*�����L�^�ej7�'��'��6픔T�b�8�֚|ҍ��"��X��Ӑ]Qܸ��OB�q��O"�m��MK�'OZAQ۴�y��'��*b��;q�8�&�c�\�!�6p~>��ɒ&�'x��ɟ���˟���3<�0����( _�؂� 6�����T�'26�(C`���Op��|��H���zh���ukr�kCm�l~�J�<���M��|�'��S���/��i�`Rtڵ:#�ɢ�.ycq'��S	<0q/OB���?���4�D�w�Zr̓1Id=@i��8z����O��D�O���	�<���i V��$A�a�x,��i�1��|�^&^K�ə�Mۏri�>��iB�3 ��+v
�!Ǐ�2/�d�� t�r	mZ#N��Qn��<��rBH]Ac�y�-O��x&��G��i� �U�>y��as4O���?��?���?������O�48���L:�MZ�&���m�h�@1�Iȟx��u�s�������JS�6� v�
�͂Q�������`ӄU$��S�?i���#yv�o�<�I�o�0����4��
�<�VNн2��dL�������OT���ET�xՁ^�<n�@'kގE-&���O��d�O�˓+8�6���B�'��l���'^��=K5�;�Of��'�6-Y¦͛O<�ਘ1gR���񎉄*�4JϤI̓�?��p��2􌙕��u3�iV>�� �1N����A4��`@2���Or���OJ��'ڧ�?I��I�	.��� �R�@���H��?!�iJr�2@Q��H�4���y'狇[3��Ek��t�)�nJ��y2j�� lګ�M�TИ�M��'T�.�(ά���ۀ �ၧm��]� ��ٳ�ᐵ�1�d�<a��?9��?����?Ѳ.�:�xi�BȴR�.��� ���Ħ��@ܟ���̟�$?��4'4P:��:[��A��	�+0�r�P�OT�n��MS5�x�O��D�O�>�J�i�
g�0�r����b�����9���P[�x��"�1i��BQ|��py®]bV0�DlұUN�)��ĝ ���'��'m�OM�I��M���J�?��L�1��Q"TeĢ;k��!҇A�<�i��O���'W�6�Lަ�Q޴<_fAS��f��5��[�5a�	�1HO��M��'2B%̧Z���S���?����4!9�leYU��9������Пt��֟��Y���6�x�mE�8����2F�1K۾�k��?��4]����q�I �MsK>�p�#L�%PrM9Z��"g!Ѱŉ'46M�Ŧu��(2pt�l�<!����1�@���H��b�����\���H$GT�$9����d�OV��Oh��GwB����11�B$�DǞ��L���O�ʓc@�栕;���'-2_>E@g%v����Fό4��(���O�p�'�*6-N��ipO<ͧ�
�А"���&�Gh�k�I���:1`Ơon��*O��C��?	p�"�D��|2�a�@lOd�<J�$4����O��D�O`��<�i����N�ʔ�qW� 
̼�q�'�<!M�I�M{��Π>с�i����Έ�V�B *��"$쬰�ha�Zm0p���l��<���tD(��&��	p+O�ӓ��t�v$�5��+���3O���?Q��?����?����iX�4�DjQ���IJ ��ei��?��Ml�,%h<�I��\�	r�s������37�͝C$���
�B�5���33��v�`Ӌ#��ɞ4u�7q�7nJ�-,p��"F�%��3�
w��b��'Nb�	my��'���
��8:]����7�]�Z������?���?I-O��m�/x%�������bTN�Y��r�N��)L7{���?iA_�$@�42�6#�=BR�@�h�*qRmB`�!n��OI`�~1آ��<i��jXp�D���?�Gd���������4����?���?���?э�	�O&0���^���Q�gS����Kg��O��o�v��d�'�6�8�iޙ�VD[w1���r?�J�n��Rߴ ����|Ӧ��եj�<��.<x�$���hc���"@��1&M� �Byq�O�䓡��O����O�$�O���T�,��ъ�c(�2��0d��uh�	*��G�!�'���$�'_�� �R�7]�Y���H�����<)���M{%�|J~����N��j^�BL�9�l!���p�ʗ:��гU� H��S���O,ʓ#�����j-i%�Ò:h��?����?9��|R,Od�nډa-64��5Nl���� ��@R�D�"��I��MC���>���i�B6���q��8��T:G6h� ��CpmZO~2D�#���ӿ<%�Og��>��� g�Ӷmo*�0���y��'("�'=��'���)�-����p���I� C�3��D�O��$Ԧ��BFvy�v�ΓO�<(�×1���B�*	�MR��:caJC�I��M��i���~���>O��ʃ:tE["��P��L0SQ�yQ䴩B�4�?!�i#���<����?����?�kSS�]��GԊr�\uZ@MT��?Y���D����(�#O�t�I��8�O��@g��$�!�B��]�v���Ov4�'�t7���*K<ͧ���J�4�n��&K>�x�����a�3Ǜ�Tk�ԁ+O>�I��?�Rg'���O0�r&E�&�[� ��5(��$�ON�d�O����<�c�i&�̈�M�2��]�%ON]=�<��"h���MÉ�O�>qҽiV�ܠ�E>N�e��I�&� �9g�m�t�lZ�^BL�oB~"�E4O�Y�S&��ɣa�J`8���~d��1�ȧqTX��Fy"�'�r�'6��'�r\>���eųzD�� I�70�|8�f��M�ń��?���?�I~�?=��w���&��Z�{ .�*��i`�zӚ�nZ-���|B���j�͊��MK�'��97ɖ!Gj�(piڪ=La�'���	rϟ��3�|BV�����ĉ��)aFЉb0�\.&
��*�ɟ �I��\��Zy����d��O��D�O����?ݺ��̈�m�v����;��2��X�����4!��'�����mx�X&��gmP���O� Z��R�.�*��:��^��?����O `!��'���ʓ]���1���Ol�d�O��d�O��}λ��p	�͍)�12�"�S�B)K��k�6
��F��I=�M����Ӽ��/K���afK�kwB����<�q�i��6mݦ���M�����?�F'� O�����e�u����;���p� �|~�-�K>�(O���O����O����O�YZq��y���5EEaX8���<�g�iR�E���'���'���R>�,A���9S%^(w3rP�P)�E�R�O�o=�Mc��x��4��/mdZE�QCZ�2���$+�'U��*��Փ?t剮l�PmK��'Q��$�|�'�t��e'G+\;�eLR-x�|X!��'b��'�����R��bݴSV���A����E/[N( j�\.k�\�"���'��'���ӛf�|��o��{Ϟ�y��^�T��lr ֟SD���HC�����?�qjƾH���������l��?pa�Ɲ?M 9��	BS��$�Ot�d�O����O���5�S�h� 3`��iz{�ƙ=��}�����ɿ�M�6!����ʦ�'�r�׈9X��"��	�is*�z#C� ��0כ�imӚ�)�t�7a��I '�z� 8��TC&��D(���^���aRcG>�?���&��<����?��?q���{��	�&�/2�%zȝ�?!����ėǦC����	ڟ8�O�m"��%'|���A��<���r�O���'װ7m����M<�'��7G\-OgJ����Z�'_0�)�șYs*����/C��u{(Oh�	߇�?���)�䓯K����,<N��D���(k����OF�D�O���i�<q�i+V�z��;��K
: j̘ӳ��>w	�I�M��K�>��i�p���Ö:m܄���D���-X�cg���nZ`�>�lZ�<��:%pҦ��ص�.OJ؆�O��i$S<#<T��0O�ʓ�?����?I���?A����<*��sF�ֻd�D��$p�j4o�=F�K�OB���O���$�Ȧ�]?1�����7C��[�FU�u���	۴����0�4�*���܈Io�,���hL�WA�#$�r�C@��(j=��I�xb�Zr�'��'���'��'���U
��H1�4� G������'�2�'�2Y���ٴYY�PΓ�?!��E�L!��ϳ<���y�Onx y���>���i� 7��o≉;{�٢D��$|�@�D7���蟬@�N�Cn�sè#?a�'Q�$�dP��?�@�&Q����\n9��0s��8�?Y���?���?���9�����R�0T20�qC��R!�\33M�OX�mZ�Ssl��'~�6�4�i��bC~��E1O�;�.Y�r�p��4,&���nӜԺ��~�l�Iğ<���m��B޹N�4m!�fE�o2
l)`�K $��&�x�'�2�'#b�'���'�V s�ҝ>W|��g�ڒ'��Q�]���4w��8͓�?q�����<iDgE�_Cn�	��E o>L �g�H�>v�I �M��i��O1�t�I��
�b^�����4�sDO
<_�1S���8h�pRL�r��Uy�ДR+��C�&�wmɁ�$u���'q��'��O�ɟ�Mk ���<1��")���q���'(��	A�I�<Yſi��O���'�ҳi� 7m�>"�=��T X��Sa��&*�&� ��o�\�I��@��xu��L-?a�'���ݱ_���#�ė�47~�07�S�<���?���?���?����؄v�-�3��>�`@�^��yR�'���v�@�J���L��4��Y'� �oZ�,�*���C��$��e�xb!g�B�n��?��������?�u�F����`�4;&h8*'e�2���p/�OM�K>1(O��O����OV��ۿ-���PC��$�f��G�O>�d�<d�iJB5��O��D�|�h،B�)Ď0�r)j�E@~RI�<���Ms4�|�'�.Ll}:w�
H��r1�_!Șm�FC�'l8,y��i�p~��O�rx�	�a/�'S��(�*�Z��U2�I�A����P�'���'�B���O���M��V7
܈��)TQ��qyC�����a+O�n�Z�W��I �M˳䚡G_8�bCt�a��7J�F�k� ݱ4 l�8�I֟$�b�����my�!�/>z���$����q+C!��y�Q����֟��	ԟ��	韼�O16�;���V.h0�q�
'M�i�t�|`Њ�O��$�Od��������W�����$_.��&��)iv�@X��M�ě|�'����j�Z�xٴ�y�b�(V�Uk c��^������y���(���I�'�IƟ�I�fN��i�薏.�N��a/Q�P��	֟��	˟��'i�7���R&^ʓ�?ѣD��f�j``���E��h0Ц��'��V���x��'�\صfV6�H�jT�B�V���Y�y2�'���0�ܱweddtU����q�@�ş��!�7Tk�!)´q� �#ҏR�?���?Y��?��)�O`�)F��2�U4!ݏ+��9���O�o�=d�$��'@�6�;�i޽���߷dþJ�C�z����"l�|B޴t���~����r�d�t��🬻��M6o*���M�b�9/ٶ�a2ؽ'x�l$�x�'�'�R�'��'*��"���.j�M��
*Z�.�#Q�ly�4Z�0����?q�����<i��ߚ�$���Ǽ�ܠ
����nN���MK�iC4O�i��(�	K0q,eb5M����`9f��V{f��Ґ)�%��$�{V���V���OZ˓)�%��՘-4֭#��P�bx�J���?!��?���|*/O^�o�`�\E���_`�Qf��ԁ`��,)y�I��M�n�<i���M#ӻika�k�t�",P��1\�P[����=��:OH���'��4���N�˓�j��_�����E�}o<1:d���bo�D��?��?���?Y����O�<�@a�P-Qʱc4m	r�4� ��'���'��6I���˓P�&�|��G�?i`�(B�S�}�ëܯa�zO�n�+�M�'0_bQy�4�y��'�~<�3���yAp,�F�D���p�'Xi�����A"�'���ȟ0�IΟ ��,��)��EĂ)�E gN��jy��ǟ$�'�J6�-^�8���O:�d�|B��Á��u�P��1N��0c"Tn~r�<)��MKa�|�'�j @K�	֩�v/ǵk�9��H$-��c�^
/�@L�,O���-�?�1�:��O�=���*���yANH!����O�$�O���<q2�i�[��I:������B4?-ȱ34�4Eo�I��M[��<��4�B��5"��L��&�A�x�A��i�B6͒�[m�6�$?�b��O�������^u�`�4&p�Q0�E�_`�d�<����?���?���?�)��9(���+H�L��6v-捋�̦}BvL�������L'?�ɀ�M�;'�Եт�HO��9���%{��r��i�6Me�)擝Aڜho��<� ��*5`�7M��c���t�4�8O�xk�HJ:�?���$�Ī<9��?Qª� 7p�ke�/��vO�?���?����d�˦�sr�ܟ�	֟ s���x;G�F#+Qqi��Kr���O��l���MKD�x�c�A V�X��Nu|L@RI��y�'_A`��7�	Q�W�d��4��Eϟ�6m�KJ]�ס�UQ���W���	����I۟�G���'Dq��ʬ��jǌ
�a�2�I��'��6͏t�˓y����4��Ha��؜MH)��gQe�&���O�6�R¦Y۴d�r���4�yB�'������?U`¢ޣ;�~aţP�0�t��dAP�vm�'��	۟��ȟ\�I ���LP���t�G�Axʨ�a��ה��'�z7M�$#j ���O^��5�9Op	{b�W�|��̹v%�=�l5$	pyr�''�&�9��O��t�O�l�qSf]=ta��"���$�	��r�ֱcR���V#��U.R�X�y�hF�_�daS4�'���т�H>9���'=r�'F�O�剩�M����?Q��ۘ�:,���S��h�U�<9ָi��On<�'7��ܦ9kߴO��]2�eI%E����R�X|�0I�M]��M��'f�&�J����J���?u�]J�P���j��`;�-C�)��}���	ʟ��	����՟��I_��ܚ�{�n�{�d�1��	TU�}p)O��d�զ��U�#: �i��'�Фs��
���s���!̰���i-����1���|�r���M��O"���D�*C��a�K�Rd��֩_y|�R��Ox��?a��?���DR�}�-L,4�t���*�xlř���?�)ORm�_�����̟��	D���Xb,д1FIDT�Խ"AL�����H}B"v�>o���S����3����g
VZu�`�BOFJ�2��зMZ`���T���A���C�oD�`	$��F��	��N2Q;"!�	ğ0�	۟�)�SHy2.|Ӵ�U⋉���P�M��)��G΂s$��d�O�	m�|�@����M��eǅ�l���'r\���@[�fu�6-���o���ퟠ@A�%#�ĮXxy���H�����}�
Bt����y�\���I��X�	埸�����OÒA�k�:E�V���Cj��9"�~�T�b���O���O��?i������,��E`�u���mт�)0Mϛ�fl�T�$��S�?����E(pn�<Ir�ׅq tCF.]-�f	���<!7 7j���D�0�����O ��u��1�J�;S:��	�+F�V���OX���O��[B�ƫ ���Iß� '� ��y���ƹvŎ ��Z��x��	��M�c�i��OH����$��0�QBZ%ei6���8O@���$����!��������O~$+�o Q�BaD�jH]ef�*!�Xr��?���?a���h�*�d�%���{�K Zn�@ #�~���i'�My2�oӊ��]8X/8�Dc&R"�d��	����8�M{r�i�7m�u��6{����=A������O68��I�*f60��cг� AH�&@Q�IsyB�'���'�B�'�N�-A*��6Cɝ3��s�L�j�� �MC�.ֳ�?q���?�I~Γt���� T<hNP�/$%�4���\����4>�&�=�4���i����S�eP�B"�	i�<���V�]^�>��d��<Qv#�y`�������Ł\�f���FR�}��`��ZS��$�O@�$�OL�4���|�f�9).���*���p�*ަX�
�j�Q/�y"m�^�R�O\l��M�Ŷim�̚B:QyTY��
N 5�1e�|��f>Ob�d�27�x��'{�pʓ�r��Sxx�@`ƾrV����E9%���̓�?i��?��?����OL�9&	H�-&]�U��f(,�S�T� ����M��B��/r�h��<��JN(+��IU�E7}�`�GV=)��'��6��ަ��?���lZ�<a�/�����e�!N���xND&Ѣ�!_8�$ލ�䓚���O����O���@�y2�EX�MM3H>��H����:wd���O����&%	����'y�S>�ka�ٱ1�=3��L��O'?�!V����4i)�6,�4�f��=xW���X�M�/C�^$ʳ"=lU`<ʡ-ѴN��ʓ�����O��H>���W��E ��\+q�,�[�͊��?����?���?�|J-O��mZl*Ip�@Q:o�u���֫kP c�Dy�b�R�� �$�E}Rnl���1��d|��ԇ3d�֡jV���MK�4	����ڴ�yb�'�R�0��?Y��Z�䛒�K'35����,A<���p
p�x�'��'�r�'���'��z��:1�'i��Rq����hQ޴U� 8����?������<a���yG�̲E@�B�>'tfa��%�9~D�6���i�L<�'�J�'tq���4�y".�n���h��^%��|��)�y�.^��i�I�<~�'��ߟ�	J����R�k�(�zQ��#{u�Iǟ�����8�',�6�J���O��䎽" �S�_��Z����5_i��"��u}�xӸ�mZ���(�E��/ϡ$XL��P�N'b�ܕ̓�?��Ł�`�J42�^�����R�waB����$1R�̖($V�z��O�^���D�OR�d�O���'ڧ�?���3(r��@(�A؎0�녶�?�b�i9x�X X�޴���y�(4y��p�aj�~ڒI��d ��y��o� n"�M;��5�M��'&bM��No���3yU<�#/�Vʴ<C$)�8K^8�W�|Y�P�	��,���L�������J@�Q���P+"h���pyRBiӒ����O��D�O:���$��n� I��VT�h�PhI��!�'��6�Ǧ=�J<�'���'12z\� ��G����I&��Y����bʘ���6:41��.�O�
L>�/O�=@aL�4E�VDD�ְBdV8���OJ�D�OB�D�O�<�Կi�F<���'"T�
��ȋB<a��*]=4��ۙ'1�6�&�I���$E���Y�4�?����5�����P #��i�2	ʍTU�T�ܴ���$N6m��'��O�>�،#@�I�g��;v�=�!�
� �H��ԟ��I���Iڟ�	M��
\�����{P��$ڒE�t	����?���Ư6�a��M;M>�����4��&�a��@6���y�Z��(�4tW��Oe�A��i�ɵ�j�b_�*����"�^�(g�,#"`�\�Ily�O-"�'�b����qh�m�@�r<�#��CO��'�剂�M�2���?1��?�)���#&�A�k��K'N�fi~�ps��0�O��lZ��M;`�xʟ�hfhܭH� 81������e%O�j����3N��]|��|j7��O�u�K>��d 5\��D�����Y:����?��?	���?�|�+O��m���:P�.��4��k�4K��+�iycr�����O�l�k�0�:�G�8�d �5/�/$�|���4q囦��.�V3Ol�$U9M<~���'{q��{��u�@�+z�IwJ��.En-����O��d�O����O���|r$b�R��
�뀱iVT��tЁ_�V��9U���rS��y�S �<	�� S�����J{�27��Ǧ��K<�'����-$����4�yb�Hn�����܁T����2��y2��Jx���.)��'~�I�4�I�yva�׎��*�I���rK�M���d�Iޟ�'�7-X"�����O��D	)IL���m[*6|�y���-R]�⟴��O�m�>�M{r�x2�L�nO*�#Q%�e^$!�+�9��$J2Mˤ5 ѠBqlҒ��98��slD�D@�n�;�O9?[�!ʕ��. �0�$�O����OX��*�'�?A!O|*$0�0��R���?A�iV� h!V�`�ߴ���y�"��oLd=�gQ7�F8Q4���~2�'���*d��i�ҍp�6�V!�)�@ �}��K�;[�����
%g�P� '���'���'���'/�'ŘM!Ž1|l��Ǝ1�P�BY�� �4�L�	��?���j+��<]䚙`�f V��ф� O��'�7m�˦�SM<�'�J�'y��K1nԳS\P����y�I��O�B�L-j/O��"���?��4���<0G��/�@T�Ձ��1�����?����?��?ͧ��d��q�(��t���5ڽ�*�#cE�m�C�h��K�4�?yL>9�R�<޴m��%~��!�V�ۖ�D��ЁÏz&��t�i��6�w�H��t�h[@�O:���']���wS��9E�'L낌�@�
J�t�'���'"��'ER�'���:FB�1���d�F��$�3e��O����On�O��'��6��Oʓd�z=���P�n�����5\��xh�x��q�n�o�?��6��㦝��?y�K��@�so�E�>Pz�a����0�g�OԙYN>-O����On�D�OЬ;��ƿMt�6Қ!
"�� ��O�d�<E�i?��e�'o��'��S�(�y�t��c�����D_rd�p��I��M�#�i�,O���R	�?;�܉����f�YP�jȠ�d�*�-��2z˓���+�O�T�O>14�ֹ1^�����3�L���K֤�?���?����?�|j*On5nڶ2X�P���.
=�=D��٨�j�@^@y2Cp�|�d4�d`}2�a�̤� `Qc!2C��!b��{�l������4a:H�*�4�yb�'�,Tj��?usTZ����F�'b�a��U�41@���
t� �'<r�'2�'D��'��S�(z��q�5*��C��!����4)U�x`���?Y����<���yl�_�8GA�:;�8�W���7��A�I<�|Z��@.�M�'����@�/ >�y�A�m��2�'�P!��C؟4�֘|�U�0��쟸#���7,?t5��@V�X�x���@ퟸ��՟���Wy��l�,��2��O��$�O�42����B�CĀ[�F�0�.������զ��4�'����s��
R�Ju{v홮<m��1�'����*gl:m*�mXq��	�?-�t�'h�E�	;Aҥdm�0X%��H��:� ������ܟ`��J�OwaR�'6��Ԡ��l�	p��#;2�d�ʕJ���<	�i:�O�Nդkl��I�J&�p��e� vq�ݦ�ܴ@2��CB$��2O��D��d�x��B�БuUIs�č�(^�Zϟ���OV˓�?����?����?��l��0�mJ�)W��{ŋ�� ��/OĤmڧ	�U�I��<�	V�s��q�Hͮ3�|!�3%	10�P�S"��'��Mܦ�۴uH���T�O����C�5�1���M�����B�lEY�^%J��2,
���'�(u'��'�l=s�lH>�����O����'�"�'����^�8	�4/P����x�����'Z*lCf��w�!���}�����_}��z�F!lZ��M�Md�f��pF�IQn@S������۴�y2�'SJ��4���?���U�T��ߥ��T�&��a��E�;鲐��r���I؟���4��⟘�Zk�3R�Ҽ�'�� �E̚��?���?!�iHXڳ\� ݴ��s,D��
�O
�8��Y���L�|��'���O͂�J��iJ�I8Ubi# "�'E䌱�`,x
� ]�,��X{�I~y��'*�'�ҡ�SՎ��v���wS �£N	�?9r�'g��6�M�ӧΩ�?���?y/�6�h@�{��y6mvK�������*�O��n��M#E�xʟ� Ne:��˱)��]Ȳ� P��JV,T&8/��@U�� ���|Z���O�|�H>�k��3��w(Ld��#�,)�,���O���OL��<��i�fQ��9A����q��0cS�K���*��ɲ�Mˊ��>a�iQ�t��b�8`��-!�*F�+�"���n�Pm��3h�El�D~�"`��1��+��%k�0�1$�Ҏ�t��,H+ ��Zy�'��'Y"�'��R>�{�'�&p��s��,
蒰���?�&�hyb�'��O}�b����F�@�E�dx@�0�Z���Qm�M��x����Ǉ@i��<O����2@F�8�]�2�ꈳP5O>-��ǋ�?�s�&���<����?!@���Z]Z N_%xb�:�Y��?a��?�������p���ޟ��Iğ����Q�|#���J7
"	�#�Q[�yu�I�Mc�i�BO�H���˼B�T���}B������8�4

�w5�Iӂ�C��u9B��ӟ�#Wc[Yx� K ͅ�k��a��F��L������ݟ�G��wk�����[-?�� Ӑ ��6G\�p�'�7�#G���O6io�F�ӼkS��#�������@M,dY4JF�<��i��7-�Ӧe:����-�'��8�R��?�x�m�VZ�֬� ��ԁc�U-T��'��I矜�	�����㟰�ɹ0ˮ1������љ��<&\���'�N6�ɇkG����O��0�9O��� �A+[Y�$��Á/DxՊ��Uk}�Na�\�n-���|j���R"��$/q�-����.d�X�a
wehP�����Y)����wO��O���H`�СEDQ�x� jUo7XlP���?����?1��|Z)O(pn��mj4���.N
�����P-���_2*��7�M���>!ƹiIB6m��5Z7�/L��K!0%�͑6Q�кi��D�O�92�fһ��a*�<9��ǿs����f�L�T���/8t���?����?���?y���O�F=�<$��TC?B?��3t�'!��'L6�^&X�h�j��F�|���fN�!0�1j5�9�b�K�2�O��oZ��M��d6eh�4�yb�'=��bȂ���Qs�j�7_-���2G�,�$H�I3��'����p��˟��	^c�c��8����m�)]4vd�Iܟ��'�7-\�'���O���|�4�����Er%e
�J�}0��WG~��>1��iu�6u�)"�)M/`���3�Ɛ2Nn^u�엩1�z��Ƃ�j9����ǟrԙ|�dX!q�h��N�9V>��ǭ��r�'3b�'����Q����4E*Z)�'+�&AD&�c�+�;n��al�"����y�?�[��*޴1��!YS �s�'��!Ό��is$6���&6�/?�#!\�	����DȊm�8*�\
&�,k����d�<i���?���?���?�.����Rf���-S�4��N��:�E��L��ş(�RG��y7�����x��S/Wh�ي� �*�Dj�Hu&���t:E�z���	c|���(z�F�s��E�&�.�;l� A�'�'�\`'�H�'���'��D1u/�*@��������I��'�B�'�_�:�4R��TZ��?)��q(�(��"b�H�"U�PwXi!���<i���MSВx�Ǹ_��t�CF6�ʅLT����^̓φ(|��f��������'	�qv*��`8:���A����OF�D�O���/ڧ�?����e<hi)��T�u�q8�ˁ�?�'�iMD���^�,��4���yJ��%5Z%z�� c #;�yRG|���n �M��E�M{�O��րE5������P�5��!>᪜ �o��G�|rU���	ȟP��ğ��I��L�QG����0#�ćIq�E��Cy� k�n���N�O�D�Oz���$���څ��L�z�t0 �� +�B��'F�7M¦�L<�|��	� d�=@�o�>��7kG/ T�G�����ެx�0��wKҒO��5�l��Q 2}*AX%l�-������?����?	��|.O�oZ�@,^)�I�Y��xH��/g�4�!7�Q(5�X牸�Mˍ"!�>��i��6m�O��"g�p�N��R.\qJ�胉�g66�>?i�#V&4#��)9�Ӗ�5@Z9 ���`�	Cx��N��y"�'���'���'���	�!�b�����?V�$L`q�t���O�$D˦��b�ryB��F�O��
Ѩ\�pn�Y ���0�`D��{��'T�6����Z��Dl^~MU;F_�Y��o�8�I!��mMt���������|�V��S៤��ʟ�0F��&ٰ�����1&z�	ş`�	Eyc|ӈ��I�O,�d�O�'%If-*���:K���%�-"�i�'f&�2���i��$��'bu��¤� ��q���O-FxJ}Vg.XW� 9�����4�.Q��vt�OD@�d"�n�~��O�o�r�KG��O��$�OR���O1�˓	���i��lt
�h��غy+\h��&�E� �fW�\cٴ��''\�Qg�vML`��KSL�!<���1�O/?w�6�֦��$�����'b� Bc.��?��1Z�d@5'�0��q@j�0|$��zQ�o���'���'?R�'�r�'��;]�p͚$�*��xц��-��t#ܴ�
�H���?������<9���yW�B�<���7�#QQ ���mu$6-M����H<�|2��Ҏ�M��'h�)���'9�J��ǥGP}��'�j�����ٟ$qt�|�]�X��˟	���.1�B�(���R��nٟ�������tyaӜ ��O�O���O��%�\�k�>��� I�@�*�P�h.�I������k�4&���� 6�2�ٵlԸ�p @3	[�����h�	���P�q��V�ӏ�⏌Ɵ��V(Y�q8T���� -�t�	"������	ҟl��ԟ�D���'혅�$�,~���)f%A(�%�OBxo�2)�Q�'�7m$�iޕcEۊ=<b�Y���96���ȧ������Y��4s�ʡq�4������ �'-��X7��\�>�C�M9xu��Q%C(��<��?���?)��?񥡚�	��uAkҽ�%� �P
��$�㦭���Dy��'�x�ӂ
^���)GN߹&.Ѕ*��W}bAm�t�o���Şv�
I��"��Ү9���J�9����+�_/0�Z*O^���_��?	 J!��<�,��ZH$fu�j �7���?)���?����?�'����=ۓ-ȟD��ˋK��Y��݊c`�Bob���4��'6,�5Û��hӪamZ�NF(�c�n?� ��qP
���m�Ϧ!�'ĝ `ɓ�?b@���w� ���.h���'�Y�w��eȟ'�r�'�b�'���'��fmX�g��9�xA��Y'q�8�I�.�O���O�n� ��͖'L$7�?�$�&����TKK�&	���3��j�%����4^x��Ox���E�iM�ɭ;;1�'HғE��%���,~�)�	ъz�"�B��Ky��'���'7b�ȫy���c��*s�B	�͌D�'Y�	8�M�4�<�?���?�.���C���'�8$��́�}�X�[đ��[�OؼoZ��M�%�xʟ���nE�51��(͇��@g@ϬJ��l���3U�R��|z�%�Of-CK>a�lΖS6\����z$�0���?����?����?�|
/Oz�o�33I�13�+FP#VN�S�rs��sy��xӘ�`#�O5l�-ot����œ�1�l�+��@����޴3s��AJ>4�F������S50����{y�Q�ɀ�r�j���yA�,Ұ�y�\�\�I៌����`�	���OZ���CnB�|�3^��U��͂�5��pM�I�|�IW�s������cvl��o��I�A� �l��:věրm�x$�b>�i�C���Γ~���#�?v�>�	 ��`�ϓZ:*�#���OI>	.O��O �PA�֔�v�h�!E3.&���tL�O��$�O���<Qֶi}؄ј'\��'J&I��A�q5P�#g�В����r}�w�*lZ��}�D��7mK;z�Q���(P \�'�`��l�qr@���dNܟ4���'��NO�i��#�
r�`�'�B�'�B�'��>��?���Qq�ͳ�nZ�:�(�	�M��G�b~2�oӖ��ݨr�и�'���&�AW�&��牳�M�V�i�6-�>9��6�%?���@.$Lr��A`� �6��$R�!����-
PL>�.O���O ���O@�d�O����	b ��%�̲8���2��<	�i�,u��'A��'���y�IN�[9��R�f�wy��+�dl��di���|�
�'�b>�z�	X`et4 �]�D �aD�F\����/?�"R<=������䓿�D�� R*�H悆Bj��Д�[R�t��O���O��4��˓V�v���y�EC�r��yђK�;'�b��n�8�y@x�z���O��lZ��M���i�v`�ͷY�� �/N�^�ꍺ"'�9�v���w�J1P������h�I�0 �\���8%��)�&3O����Od���O����O��dI�ZV�9�<��A���.UfDE���#:ҥ�K�Of���O�mZ��tA�'R&6�-�D!%o�a���$.�NxZb钄@��&���4z���O��◺i����O���&[:0�a�	�&E��l��
'~ ��+��d�V�O���?!���?��8<�,��(ɟNN�Q,�$Qs���?�`:L0B�,�
w�(�,O�����瓰j�2A[�CP
�b�T�S$*Y~�t�I��MB�i�RO����@��.�<2YP���Rd9p�kge&�@9�d5Y��˓��դ�Onq�L>!S`�C���B+�#[?��x���S<���i����@ο:��u�vF�%	���+�$����&�Mˍ�F�>i �i�^А	�>?k
�ض��	e�0��eӒ�l�.�x�n��<I��O:���c��D�x)ODi��M������T!ztv5ʠ>O\ʓ��=�,���$�k#LK14:ZI9��K�$���ɀ�qo��ʟ������y�⌓jt�H��*gV�9���ZL�6�ѦM�N<�'�b��E�d��4�yb�Y�8��$rVLR����kRFǸ�y�/�g�"y�	�&.�'���Ky�̌q�,D`ê�#� 4WǕ5�0<���i,l�� [��	�a�:���d�(+b��&��?QFQ����4yQ�fl(�$_�NV�EIu��4^����	;m�$�O�)��e�'D�.���d�<���9��D��?�a@R�6�f=4�\^��d:��Wg�<)� �1)�>ɪ� P\�n�{�-���?1ÿi���b�[��{ش���y���{0��P`O�%P��y�D��yR"c���m��M�4�[�P#;OJ�Ċ6~�^����7���8�%��s/aK5���*�|��!�D�<I����*�,�:�*��(I )6%��	=�M[)G���D�O��?)k!�:���+���'�N�#������O�6m�I�韴����x"� z�%@۰d�@5I$��y8���c�<!�d��6q����䓵��>�H�92�z�AB��a|r�w� �H���O(u�� �Q�`}�Gl�0Zk����;O�IlZm����4�MCտi�>6� B���h2̊b�Xa����
N� ��7�k���		X�Z�"��O�2L�' �t�wrl:��l���cgɏ�&��(�'A�2��/�-+01t*P��Vɇ@�����x�ش2�^ �O�6m#�d� �]�S�*i�Mi.��Ro¹'�Hm���M���q&l��4�y�'��m����"m�����%J�gH �b��:p�5�I/�'v�IE�.�1��NW�]�$S7*C�$}Exr�rӸ�X׬�<1�����T ��M �HY�"��!X"
��ra�������O 6M\D����i�<�V��%�
A<q@�)�6Jx�c5��	7�Q��<���o$���D���U�N����ܸ~�DdsA�r�x���M�˱�p�3�L�g/��Zp:
�C Q�L��4��'#����Vl�/~H��(?v2��J0�:�6M	���
5N���5�'N���I��?�J�Q����F-�~ݐ��Z��srk�̖'=�{��_��ѥ�O��'Ţy��7�G;�p��?���$Be��>@Tc7n�.*DD�b$^	V�@�m(�MK��x���f֑ �6;O�ܒ��K,[��@0��h�4O���K��?)Ӡ7��<����?aB�A�}�z�{�.G-O���C���?����?�����礪���ty��'�(њ��

���� �Q�p����f�Mw}�/j�fo��ē6?Ԍ)_��pq��N�����;?���M�1Dl�(B�X&��"A�mZ�Ll���H�D��7BM�)��DZ,SJ���'0��'���S�$��֕��@	C!^v���П���4<p`�'��6�,�i�)�����RxBu�}�����l�Hj�4/��v�d���a'}�t� 'R���|ם ?M��3�@�5L�����&]j C|�R���͟���Ο��I֟r�ɄS�ܔ��E�u9Ī�hyBai��]��8OJ�D�ON�����Cԍa@�Z.]�����
M9Aθ�'�v7MP���!O<�|*�,;�r�"�Y�"gVA�&y6`���i~B�L�n��IRB�'��	�*�� ����x" ���ϟ#�`t�I���I��\�i>y�'��6m�~1󄌌&�2�B�l
��`8� 'W�H=��U�?�`[�4��尿��4ev"Ń��G4i��2���<�U���M��OxR��ܝ������wt�x�$Nٔo'zd�#�3��1��'�B�'�']�'�(�Lڄb
Ak���m/|�y�1O����OTm���>�:қV�|2d�a�@�ځe�Z6"�� BI�Ht�O$�$i�󩎪7|7>?!��0:c��{�� ,3`$Bk_>d�l��"��O�	�J>�*O���O����O����\h�� ��L�;7��x�n�O��D�<ц�i0@�'W2�'��S�?�RoB!u�:=����$
l�:�����M׷iȄO�SG�h���1�H����1r�Y`0!�j߮�<?�'xԮ�����J�0J@���NF�:"�G"����?����?��S�'��ݦ��$�~�t!�D������Ǐ)fc��A�&�D�A}b�y�Dp�wbFj��)��I*e�ftʢGT�� �4��2�4���@��i�����SԐ�f�9,x���c�6��Yy��'��'A��'
�P>�Cc�CǮL���Z"��ܘ�@�1�M��&��?����?�O~���c��w��:'��/}ء V�T�v�����z�D�nZ���Ş.o���ڴ�y��ƴN�pAH�+U�R���6B���y�	T�Z���mb�'���؟��	�rUĜR���"-�V���}\v�����,��럐�'�(6m¶^�Z�$�O���R>M؜���(T|~��P�ԥ�:�X��OܼmZ��M�A�x"�="d#j��i��d �hU?����:u�P�d��*rΤ��h	���~�&�-5����R"&5"F�J"*"���O��$�O��D3ڧ�?qc�>-`H|z�o	�[���;0m�
�?	�i7 4�A[�x�ܴ���y�n	4}�Ҽ#�+��X�\2�d@��yҥm�xtl�M�����M��O� yt�ʁ�J��֣0c��X��B�tX|�� :n��O\ʓ�?q��?a��?��I4i!3,E�^R���C��[@�-O�lڦh4&x�	�	n�s��s��>3֐j���?j6��v	����X���47Љ��OCF�"g�8,���;e��!g�DPs N�w�&���_����`:12�Co�IFybh�ZA\�ۥ	D=%p*h������'�B�''�O�I��M{�<�A`Ժʌ�Z�N�C�82�i��<a��iI�Ox(�'��6͈��(�4-���81M �	�%��ܤm�DZ�, �M��Ol����/�j����w�-���3��C+���a��<	��?Y���?i��?���� T	\:b�M�KW�	��X��y��'�"Fz�Bl�!�����4��1HZ4�$&3\3��s�#_�� I��x� g�<�oz>%���զ��'e��a���'�l�,� df�%���eRX�	�`��'T�)�s�H��J�(�xq򰢁2?���� �!�j%�&�X+W�񟀗OP�������T�br Y o����L}Kx� po���S���^�"$2`H �[��d
DgS�&=�=8am߄i���[��3|�b^|�䈸�������P��8B�ɕ�M��f��3� �*Cj�|�0Y���U7_�f)+O`o�v�z���'�M� ����	F���]�pb��U�Ϧu�ݴu����4��$�DF(�+�'rbDʓOb�0�I�0�0T�v,ڑ�z�Γ���OV���O���O���|�Q�=f�^h�ɍ����7�B�:��D�O���&�9O>�nz��3��?B��RqטrH4������?	�4�yb^����PXŁ���	�_y6ċ�k��^4p}����d���I�hq����'1*,$�������'Q�ES�%�`�R��$�:60����'L�'U�V��9�4������?)��8�Q�G�>&�P��1Hi=�%/�I����O`7�s�8�'�����k���r@G�*�q�O�ӵ��3��TТ�Ɏ2�?���On8����|���E%�M��� �O����O����Oޢ}��j��I��f��T	f�M�z~l���GP�6E *��		�MK��w)�ht,����8R
������'�J6��Ԧ����t� hoZr~�
�� ��ӃF��1 ��3{����8z��+��|T���P�I՟P�	����g.	�EID��7����U��ny�{� �'�Ot��O�����F
h���"G�E� ��ȉ�<Ҏ��'�7���!��H����P�?��U�5�6���Ǉ�%u��仢��
ǣ�-v��-d@ԣ�N����[�GQ"t×(څO|A+�V-趥�����[�"�$Q�a!�Ӆ`Gr�Y�JۥCG*!�Q/>���5���C�l�4%�9(�r-�2��h�cj���T�T&f�B�ѓ+K 2�.��m��I�@qRf/8��0P��h�Ը;$� k�z���Iң֢��e��Ԑ[�U�|�m*!��7$AnA� �c<��jtL߹,�r��Qc��'h$p���X�H�ܑ1F̔�2&΁�ƈ�,�R���`u�d9�#c�c�@�ҡ��/^��D�خD赎�6"����q�6�G�\"E�(v����5��^}��'v�|��'w�J^�$��!Q�Z1��S�h@L��%ài�6M�O��d�O6��O��`kC�O�������c� ./�̩�3� �0L5�'	k����>�d�O��H�RV���x ��]�Ȼɉ����%��MK���?9���?y��	$�?���?�����ͷDrr�!vl�#0�R疭6�'G��'���8f����������c��)G��8W��Сp�Z�X��f�'�c��:*��'��I�?������0��y����eR��4�67��O��D�[i���f��I͖+8@�f�<|�����8z����N�cr�'�	�?���џh�'p�Y�b6�u����e�,Tk�{�ˆ�B�n��y����O�=��T	�Ԙ���A�r2��J!�˦e��[y�_�)���Zy��'��D�U����SHD�}:�5ae�ͼb�*��<y��?��'�?���?QE,�Oꂝ���@+�ԋ�2;���'?$a�R��q����'�ē�?�I��+k�@�f-E:t1�'��.�^�H�O����O2��<ɦ"�\�H��B��FpR�*c��$ ؉�cX� �'�2�|B�'���ݪ,Y@ Vh��֠0ǁ�&�|��':��'��	~���K�O .U·�4jT��Hrb��b�x��4���O��O����Oz�9#����p��+$U4�ЄR�2�j�B�>)���?����^J]�O$�	�-BY1`K�>���� c�ws�6��O�O����O���>�I�@��ȡ՟$�
1-�@� 7��Oz�d�<)��ZT�����H�I�?��v�l���J�/�ưH׋߱�ē�?i���N���Bܟ�8�G��0���U� �2��i���
t
�L�޴�?���?��m��i���w�C(Ɉ�+G2h���J�z�,�D�ORd�,5�	nܧ X�@�$�9#`�hƠC0Tۮ oZfd\Zٴ�?���?���/(�	Gy6GJZ`��?VQtu�Ҧ+�T7M�e��$>�$)���h���e��lTB£cR8A��ʝ�M����?q�<��]��[�h�'���O�R�ς�m$��qC��saf�`��i��'K(b@L/���O����OV���Rg���b��B76�4u�$�TצE�ɸ�|q�OF��?�O>��+�R�cm(=���l�&Z���':`����'��IƟ0�	� �'�H���9 ����0��,x��Jq�ī�x�����Ob�O����O�p)UFͮR^e[F�"C�%��΃=_ВO��d�O��$�<�'�N�I�bڭ`�(ÖYtA�E�x��\���Ig�Iӟ��I1����4LX{����� �C���r��O����O0��<Aɏv��\{sdX�m��ܸ��Ǣ8m�Y��-ǂ�MC����?I�}A�Xq�{r [��"|�ũ����"�� �M���?y+O��R���K����s���M�xjq��a޲E��qÊ=��<���L��?1I~z�O�z��bE��*��D�p�L��޴���6;*�oڐ��i�O��x~��5��}pS��.%�v�����M�)O��`Ť�Oܠ&>�&?7�[1. ��8Ō�%y@�x[i�<nZ76zx޴�?q���?���v̉���@�}\� A!OZM��q)G�t 7�ҷd`��$�O,˓���<	��$S�1H���N��J$ȒD@2����i`��'���q�PO�	�O~�ɕ���Di���H��։cF���4�?I*O��p�J�}��'5�'!`�����#ϩX��x��^�v��7��OJ\P�L\�i>��IY�i݉ rG�h�r���Eʎ5���9�#�>3@��?M>i���$�O�i����2�i�e5�t�dj�-1�ʓ�?����'^��'e:5��N6Hdx0���Y;V�i4�GHf�x�y��'H�IʟLHƃ�X� �8�&Υ*5������hйi=r�'�O����O���CF�;ϛ�
�5	�N���������?.O.�D�^�r�'�?	X�ډjɂ$�����)R���nk��?i�d�:T���q�I�w��ժW�	�Vy�h��ұ��6�O*��?�E���i�OZ�D��klC�=K&8�%��wcN��aJ:7�'�R[���.6�Ӻ3'`�p1���� wx)�L}��'�I���'��'���O��i��Aw/���uy�7�0d~���D�<� Jz���'L ��a�Yj�|� c�	HL$�mڹ���	�	�<�S}yʟ��iqD[ 0�Ƭ�CΗ�H����\}J��O1�h�dP (�:	zr��=�T��b	��l�꟔��ӟLQ�dٛ���|���~�F��2��A�`M�>=�6�j���.�M[����$�S6(���y��'Y��'�ʄ��+0 IX#/�:+�4pf�vӰ���?j4h$��ڟd$��݈Z`|��	�x�lq��F�x�F����$�O����O��e�()wJ�X��	�O��&� �ےk����'L��'�'M�	)*��5s�@�	b-��P�B�XJ��d�Z��0�'"�'��P�0�������d�ƕCa.�#��,;� ���
�byr�'���|b_��2����9�%���lyF	<7ص*T�����$�OV�d�O>ʓ�,�Ж�A�5�Ι�$H�Ex���P�L�u�$6m�O�O ˓RV�в���(h�d*P���#@n��sǉ`$6��O��$�<���L@I�Ou"��5F-����0{g�۹d�&�QHR����O�˓}`��B����'���욿g���mݕ/:b�AGU�����O��HC�O.���O���⟶�Ӻ3u$�Y��&�=J�P\�)G���'Y��-u��y��Gӊ	�u�4�W?v^��;PL��Mg[!�?���?����
/O���	O�D�"�%bk�E(p�S3ga,|�ݴZyܝA���N�S�OW_��xJ���$uԅ��I�:|T7��Ob���O�����<�O��p�&!B4��+܈����f#(`���Hg'֝&>�	؟���$DLڸ�ЍC�N���#�#:���ܴ�?y���	dщ����'��QZA�O i����p�0Y��$�eL�j}b�]#QRT�������	Qyb��!z2$PE�V��B�ÀS�nY"I#�$�O��$2��<���9� 03�FΗHF`��B]�B��?Y)O����O�D�<i��+��	A�AF��C�H0 ��@�J֩*��I� ��J�	by"�hy��H`�Z�I#���)�����N8듅?����?q(O�ѹ#e��d�'�Z( �Ŗ�g�"�����cV�hV�e�p�Ĺ<���?���~�d\ϓ�?1�'���c�l��Lg�*:�XU�ߴ�?����֔i�^U�OZ��'�t�R�a� ��I4���Ef�����?y���yҊ�m��^��'"N�T�C��q�ܸ4
Ncu��l�_y��3Q�d6��O����O���DL}Zw�[!�� ���H�&(i�ش�?i�dK~H͓�?.OB�>ʂ���)����HB�M�Ԩ` a��08$e��������I�?�ʯO|�P�^���GĎ\�|0d �B�y9P�i�
�a�'��'��z����dQ���S�Ūbi���֊#���o����I�ԫ6D�����<����~BL�~<`����T:n���g_1�M���?���x�~5�S��'�r�'}�E�3�?�>��!�� �H��j��dS70���'����$�'�Zc�,1�O	�_�2]�b�[PK<t��O�`�e;O����O����OH�$�<��·RY2���g�,B�a�o�IF�x�U�D�'��T�@�I�����-4Ad8H�b��t�9�<�I�4�Iܟ��'|J��u�x>qh@a#p)�NT.���.v�8ʓ�?�)O:��O���U���
jx���(͘}�r����;rՔ��'���'f�\�PX&J^���i�Oz��6�H�p�<4#�Dj;����䦑�ICy"�'1R�'�^���'��7��4��N֏N�t}����F9D�m؟t��ny2D�D���?y���2�H,%�޴u'�-XUNGJ�"lu��������8§�q����ly�ݟ8!"�
�9���#��� q��2��i��	F�y�۴�?q��?!�'3q�i��#k߬� @掍	���ȓg�b���O���t3O��d�<9��$�W"���#�ɑ7�L	��k�MCCj5���'���'�����>.Ob1x��/
HUaQ���h�������R)h����џ,��B�'�?B� �Fn�֮X�i�&a���}I���'�"�'y��(5@�>�.O0����[E�Y3C�e ��
4��]�!�fӘ�D�OL�D��OM�?���ΟT�I1g�&��#�*��ϒ0P2��ش�?��.�A��Ly��'���̟�(3G(�a�ǚ����@�]�uD�`cb���?1��?I��?	*O>�b�OѵBע�bkROx�PrX��!��>�,OB�$�<���?����|Xg��%��`Ȱ �P�a�# V�<i*O0��O����<�C!ZL�i�| 섹��W�f���wJ�W�_����|y�'v��';��!�O���V%BXTE _�(�b����M���?��?�*O�����\����5��
�H`,����/�ހ�sBO��M����$�O���Of����?�q`d��j�w���`!]z�m�ş���Ay��Z8�4�'�?A���� ��k�(�-����4��28^8V�h�	䟐�	[��T���'���
�G�-KSe�&	�,܀w$Ρ`���X� �#�F�M����?A��JvT��ݪn�B�# '�}�\)�AH�d7��O���M�\��,�$7�Ӑ[t���d�*��DlF�7T7����.�nП0�	ğ��ӛ����<a��>C�� Y�%�4����h�t@�6$0�y��'@�Ia���?ae˄N�>�"�H�C��������P5�&�'Lb�'m�y1�Ŧ>!*O�D����GL�+=��Y�D
�n� �Bp�>�/O&�2����ݟ��	���]20�e1�N�#��L� l��MC��p�l�YUT���'��[���i�u��AU�RPBa����#k&�x�&�>���M�<q���?���?Y����d� zS"�q(�<U��Uȓ�ԫ>��dj%%�[}B^����^yR�'�"�'�q�� uZ0�X�gA�b7|]�E���y"U���	��TybĂ�Y��,P��5��(G��Έ�l� CE7M�<!���d�O���O<�(�:OL����:�����R�
1���Uܦ��Iܟ�������'���Q�G�~2��C�*�/XtUUC�'oI\ɱ�զ��Ijy��'���'Q�:�'�s�#��R|�T��)��O�&�i�B�'��M�α鮟6���O6���70��a�
eq�lҁ�Y,j̕�'Z��'�B�� ���<)�OҠ��� �i�m�3��&{
�*ش���BK���o������O|���}~`M�~˘�9se��4sJ�S���/�Mc���?�����<�M>َ��ۿQ��!���,7e�!� -��M����.��6�'���'��T�>�ɾQ�4�#@%�ts2���HRC��ٴ��͓����O�⌀�_k��wA�i�'�?L�l6��O,��O�R��BM��?1�'���$�)fB��LӄD�F�Aٴ��M��M�S���'���'�>!R��EN��店$:PI�ԙ��d�����<v�b)�>a�������7X�����>'��i9b�C}2͇�A�_��I���y¨��
��U�S��\p���Z��EQ�0�D�O���*�d�O���Q�/�ҁ:�EO
)��@�B�M�WpSU�O�ʓ�?����?�+OH�����|:OP!�&r�"��	� ����l�	��$�H�I���y��f�*cŚ���9�%�� ��b#b���$�O<���O�ʓ[�l x&�������y��E��~H�%,�
)��7��O��O>���O�uJ�c�O��'v$�$�5=v�1Q�&E��=�4�?9����$��4&>q�I�?��MܵZ ��(]tڸ������?!��&Ix�����䓂����
9N�X�E�G-s(�`��!ǻ�MS)O��	���Ŧ9���.�d���Q�'�� W GhBGÑ�1�}�ڴ�?��*h�����OH��"� Q�/���
�?)����42n�$��i�r�'0B�O�b��"��I%L�<4��G�&�EQa�-�M�%��?�L>����'�0�R���
u� ��h� Q<V�r�Is�����O��S�}/�d&� �I�����]՜�Q!�>tv�Ab��2aB&@ns�	;/����sy��'���5�Ԉs)3�Ё/*�l+�ğ��M;�r/�Ǖx"�'��|Zc,����.t^�1ՠ�7R�h=�O�E�3��O���?���?�.OR��ǂIx� ��H�$�`����6Z-H��>)���䓘?!�� �ڨ��d��S3�-b¢�eҵ�.�<-O|��OP�$�<��L$��3,��J��/'ԍ�uF��r1�	��xD{��'��@{�''X�"d@�W� ×�O��1�cӆ���O���O`ʓ5�6勵��d�)J��0 �ص�<$���1M�6M7ړ�?᧡L��?Q���~ªJ(vH1���(<��lʠ�M����?	+OLh�G%IB�ß��s���# 1N�
#���$�1׌=�I��l���Rǟd��ly��np�u�2<&X�S�L(�|pz��i���'����'��'z��O2��5&I߇[�Υ�@(�:d��H[��
��M���?A&�F�Ԏ��<�~Rg"O�8����Q��UD:���W�����X��M���?����J@�x�OG2096GJ�t�b�{�c�v�Dx�t&x�Jh��	>�	�?c����)�J����� '�Y#�ʰ8%z��ݴ�?	���?Y�#�?!����I�O��ɦJ��`�fʆp���G��*?ԐQ�yB'<;�*�`��O��D�`t�IA���RAP�ǅ�La�en��T�V���'t2�|Zc
��K�'�f\�Q�G�g,.�A�O.l���d�O����O"�S`�q�!M	y��m@�JTVn�� ��ē�?����?�dpaKe8_�,D�D���>�`��q��?q��?���?�o����œ �p�pg�*'ZL$�L��M[*O��d(�$�O���	U,��i����W�ˊ�����+�$�8�ЯO(���O���<�2��4�Op��E�5JH�1�@�����c!�}�H�d�O⟘�g�2�ӄ�liH���A�JT�F��(>	�7��O����O*���/˧���&��#��!0�0�BwNKZ�bQ��U��柰��t����i �~BAD�k3P�A��:����@Ц�'`*DZ�i�꧔?��i<���#ў ���ą���n�:7�O\�Ĕ�"9� �}bq��"��]	"d9'�R�Z�����c�զ)�	ʟ�	�?�J<1��r�� >���c[-0)C0 + �A��iv����ğL��D�='��r�}@�p�F���M����?q�~�,S����Or�	(O��gi�n	�!���H�b��5�9�Iҟl���d#���UzL$`��0jת8{��7�M���B�Q�q�x��'H��|Zc�z��q� ���Cq��>�A��O
����O2���OJʓ<�Љ��d��4MfͲC�įNc�`$�FN��_y��'���ߟp�	��;�I��� )��焗 -�QPEBo�@���|�I��	���'�hU�P�{>)Q�3t0�e� H&�t��+z��˓�?�)O��D�O|�DH@���I)K45y��A#��[f/U{}r�'�2�'��I?@lfȪ�F�K�%ij���Y�w|�ٳi�	^٨�m��l�'�R�'��K��yr�>y���80�vi+rj�y���T��ܦ������'�7�x��'L��Of��Sp(	�Nࠤ?e�:,����>1���?A��`��	̓�?I*O6�/���i�䍪sF�1��ÖaѾ7;<���%�V�'���'�4�>�;-�ʼ�e�ȁIӾY�#�V>Zt�1oٟ��,/�#<��d���}��Ayr*�7fJ*��U.�M�5�]�RL�V�'���'���>1,O��K�G%��uQ��A�>Y
o����St�4�'3��)�OLP2!�Z�� ��i���[ڦq���X��0���P�O˓�?��'e��Z��A��Mq!A�!?@<�2ڴ�?�*O<p�4O�ǟ,�	y���$�>�����1N��s�R�e�ɻoKPq�'�"�'�?yH>���I?H��nA(w��+3����I�fUbc�h�����	ٟ���9Q&���#
~�V` @���A�Ly2�'S��'#�'R��'G6p���w�ҼBBC�/"`�P!gJ�N�\��O<���O����<c��
MP���6 Yĭ��-�:ot|�!��&L=�f�'���'��D].<��ɭ,c�
�a�'���@�Q���?y��?���?�fFH��?a���?�
0�8� �02���i���C���'�'�P�lr"A1�$W.#�Xȣ����$ш��!��k��~"�ֽ)����%�4
�ƫ�y2�%@\&��m�{���! �X5tp�M2�e��M���w�KQV�G�#MG�{�l�j��Q�R?`X��r���DMle�k׭wdD�{�(�LvB|��CY9D̞���Q�z�i$�� p%���mܻ[<��t- �X^ܠF�[�5x�%��W�`7@�s~�`�aA#>�ʑC��Cư,�aӪ]6�$�OJ��Ov��;;6�0�؛67 �1S�̘	�Ę��fW�10R @�
�\������Oe�'Ő�ҶL�x76�+2�I;��Ҧ�U I��\ɔ�:`֠S�]�I�x=��+�|�E�%K���݉W���2⦋�W���G/!�U�Ie~b�^>�?�'�hOYPv��:)���s�㗶U��p�"Ob��V?M�(I+�!����|�����i���?�'�\5'��xה�W�C/-؜�f$��S�
��w�'�r�'Vr'p�Y�	㟜ͧi����N�~�#���~����`D���\8�V�R����ϓ&�l����ڇ'�`٪��$utt�# m���I��4
B��;
ϓn��(�����8���?�(țt(������o�'��Ol髧K� n�6YYg�
^QQ@"Oq�����Ii& Q�1˂��M}BY���������O��cegK�?D�fN�l	�7��O��D !��D�O��S֬Sb�|K�j��5�
T�OgF�8&'N�����b,6O�!���(V��u,�*l#����#>.i��C߳.��i7��>�p<���Ɵ�Ity�Yr�j�!��*�4ੵ*B#Ϙ'��{���O� �	mj�\9j	�xb	r��Px�Bǻl���嬂��xtC$8OD�B>��ڴ�?y����݌?�����gW���V��L�+�)��P&��Or��P/B�l�v@�7�~�[>��OG�l*׋^�+�:���;2�O�P����S[����L�~ŞU��ڼS�ҹa��?�ɱ'�.(�tj�퐈aN�A	(}��ۡ�?y��i�\6��O(�?90%�
&}Yd,a�T82h���p�H�'B�^��g�S���Th�OvP�鐄Z�;""��<Ɉy2�iv�6M�OV�lZ�4R��@ ѩ��ª3yD1AaT��M����?���cF6�FC��?����?���ҿ!�B!]L����V�x����N
'Dh ۶縟��׍� v�$?c�Z'׆z4����K@/�y�GչD�m�T\�s���s�̒Q[��>5 a�<ɖ��x��#ՌX�_dT��$�^��?��i�r��*���,O����5V�\iBA$	8W��i�.Z�����>y@�D9��ɒ5G\m`��c��B��q�X�m�]��h�DP� ȲB�0G��G�� )���� D��Ћ��u����f(�ZMD�>D��2tdѦd/�=k���%8V�"�7D�,�v�A1��t
&��2M|���:D�(q� K	i(���JJE�AKk9D��;EJ��N�$ܩ&����Y�c�6D�� $�WB����#��<�D���"O�i�M�
�!�`ԌE�~��"O$˃��L�ddO�mrx$"O��.CҶ��Ʈ* �����"O�1s  �&����N˨<˄��E"O�XQЌ�^)ld��k
;Pj2-;1"O䍨C��BI9��U�-N�T�D"O& "��_�9r�"�'"I�}*�"O��щϺCd
1��=v+�ѡ�"O �J�m�#Z�|���	]�vA��"O$��H�<P�P���nH>�X��"O�J���T�f�
Q�e����"OH�!b��kj�lZ�
���@r"O�-�q`�3�L�
��a�h�i�"O����]c�>�; �T�X~z%+�"O
I�G@���@��@�s�%��"OF]�0��=�(���A�"`[d1�"O�Z�GL�?�(��`�:n^2P�"OP�p�̓.hNt)���
��ґ�"O�ْ�5�u�MP���"�"O<(J&)�6N��Y�V��yS�"O|m(�"�'o�*�Ɔ���"O|EC���+�f5�Re&k�}CA"O<�i�>/Vt!�qi҈N�^�y"OR�Qd.��Hb��kt�<�dղ�"O.C�I�\���:���,�<9kS"O�4Y!G�.y%�Ī���-sBdؤ"O\�p�ۂ/�Q@�n�3Wp|�A"O�)��#r��! �ѫ"�f4� "O�=�R"�w����KƝl�\��"OP��Nٛdv`��Ȣ��#�"O��7��פ���F&$�J(kA"O�����#&��A�"�����c"O�A@��r��B���̌�R�"O�Y�%�5R2��넏C�<��"O�0a�_9G����G�#|<��\��s�j2�S�OU��+���H0̴��Ȑ�zR,���'�D ���F�/:�W*(-]>�I>Q�**�0=�գ%���kC�V8;�A�!��M����U��Un���ŉ�
TȽ�����n8��&u�u���Ca� ��v���u�ER��i>s�'�>׶<�p���y�6��� 9D���v�C�g���O�A�>!����<�Go>���(�xIT(�<W�
Y�R���y�$"O j�jӷ?B�R��E)r�n��2�|B�D+v�az���/W4j�S'�V�lh7�{����9�n�bc*�0���\�j�L�A�<Q�"5X���#��.Q�	Y7���'�pub6�S,u$.=���޴%�hI�N3�C�ɱ��@*�Fɠ"4<	�A̘
v<�!�����i=Q�p��F�K�%n�0�7f��x�!���pf�Q+I�,�f ��PXq�'�v � �'S�Y��(�x��&į�~I��'[�0����`y��,�.i�b@�ˎ�y2�"L�ű�l�rvl\�F�G�y����2^������,� f ��y�,[�x��q䝰ZL������y��t�~����C!? �A@Ȓ�y�H�(�B�k���\r�g�H��y�e�$N��	4��� ��H���y"Y�D�y�%Q
hݢ��Ѕ[!�y�+E�<l*=c�e|��A��R�y&/wU�t�AÝV}��'�R!��'�txjL<��T0�.�fY�W�O+.7��{WJ 	����S"O� ��qG�*$:E��i��\�tԁ1@���!�0���(���)^�6�yr�Z H�����h�DB䉱T�<,��F2V�0�O�}85�'d�'+����!���R7C�&X��Ub�4=<��C�;|Ofh�C�>եJ��M����UZ| u-PU�$�1��a}R�J'<'b!��i��\�j$a#���')|��L<e&������� �|ՠ)�J(Y	`"O�̱����u^|��.��R��Eo���' ��P3��H���]5��u@ӂ��c���hQ-\�"��C�I]6�iE�<F;��h���$�打R<������6ZX����Z�'񾠻冈�i}!�$O#R)� �@�7��-B��$~X!��[=��t;�V�yL�(�A*�!�$�(K}:="�%N@f	�e�N[�!��$s\�}������|℅�/�!�$ܽP�\s�JE��U����T�!�D���t�6��%�s���X�!򄊫U� ��V��c0J!�D -i�to��V��a�O�<<!�dO�e�5k�i��,��l'��6!�ϗD�:ibpE.2�<5!�e�72#!�P�;�`���20�B1�J����y��P 1O�a����RJF;E��)��"O ����k�x`�IO���z��>� ���X��x��$��y����ӳDLd����yr���qB��Q#��G�NP���0gxQY�<�r�����'?� c�Ο#�Z "��|�J]Q�� �O�!`���Z��A�Մ;�l�%"�:��3̓- �Lڵ�'и"A�=�aې�/9�"�{��� i�n�s�öd��bE��|:P�B�B����59�Փ��x�<�{/�Q+��7�����uyB�X&\��Q��3��B̮~���`��3"��(�.!W�&��UmN��!�D�k�3���(	���u�(K ���V#L<�n��~z^�Z�e;��ON�c�O֨)���1D�z�x�oז^D$�QOV�*�̇%-(�:�h��`rJ�e��V �Ԏ��J6�	 �D�y���8ŨO�)xH�7kIzQh��Pb1h�;��'�<XT�[�XE"�G��M���P�X<BH�'R�<�x�Sᗴ�?�E#�B��l�V_8�2KY�_a��b�o)?�Ei��twRɢ��ǢM
��F��}�f	Kq+-�d�J>i�dI �LG�HxZ`*H�y¤@(ּ̉���?��1Ҥ�̚z����g�Ӭ����7�-�N���4�iR���'<�!��,��X��T2[LD����u<� �[\p�A*�P+���`�X2	VRL��	ߎxd����W�K�$�d�i~(�����G�	����
`NI�S��X�ax�C�035 qCuF��n>���+��,��K��ِJ�yA�fޤt{��;u�/$�Ař?4RjdA�@J�����-4?Ʉ@��j��p �)B� �(9�NZ���O��9��b�m.���c 6e܄8�'Wf<�� m��prF�"G��(ui�YH��	��)Yb�P#req��'R��Xr�M�[8t�P��9��- M�'C��i�a*��~�d��r^:EI��s#L ��,�G^�J`�P�,ыz��zҮ��T�!tK�����΢���/9`2p8�{�.TѨ=(�ȭ�����ݶOR�tK���-�@�b⃏,�!�$�wo&�+�
u�jЩu��%��'�z����ERs�n��~҃O�_50�z���Qn9��p�4�F���5��I�~� ��3��,���ELi7��	���Z�A��J�/.���I�9~@"|
����?�Al�9n*�!�W&Q�7��C��Q�c1�4��"'NV�_�J�b�F��)ݸ1 �cG;"d��A��f���	:�ʐD{kH�>>A�w9����*�0=������A��Ò��m��[����R��cL�sì�<X_�����i��8��ɴ+/�M���R�2b Y�*\=8�O X�"Lx�M��jj��r�E9q����o��ih-�@m;�8y�  ��{�!�D��τkEx-�6���d��\Q�K߂Δ<+�x,�2���$�|K4?�OҮ�˙w���(��&F0��E��D��	�'���Tݒ(�@��&�ݤ8WTH�0�dB�k��x�D��h�E��Tm�'�T\�,]0F����a$9o�p��ۓ<��� �% �|��2� ��a�l�'u̦�bT _'<��!P)�;&IFxP�d�
��t�ī�{X���'�N�vr̈s%��'D�So/��)rT�ٗ�4z���3'ƅ�s�FO\��C��� Mc�eg�V�؇�`H<QSF�??�@�`$��-R�`1U��=u�����+��P�&�6UޓO駻y���.�Vز�oA�7�&��怽�y�o��
N��`��[�	Z��F[|&)%���NK6���L�*v���ɕ�5��d=��p�)n��D��F�|-���,�1 �cA#|IzY�4��+[D����Ȍy��3E����
��AO XH�͚HM_x��s��dY8���8�l���H8Y��#�'k#K��1�
��<���}�T\�/�,K�u��"@>g%F�a�'c�hǈ�jxB��`��c0�*1��6h��/�J�> ;kـR��)���E�#нp�8W�>�l�r1"O4=Jd��=�҅�wa�RuBUFÃt�&�KK�tj������i�4a��t�תX�L����ҏҧ-N�tf0�O�u� ܀NpZ�i]N��[��?<��{� M�t�@cˑE����	(\O��ʲ�J"Z��������1@�� L@d�T-X�L@Z.r��M<h|B�BF�#"��a #A��N]�ȓ4���b�J�W�����؜h|J���lF��{�b�!k��̋¯ľtv����94�-�"��$2햰#A�e��?�"��#8`�?mB��YP��2��0'������͔%^хE�
S)�q�9���'!#�O�� �
7�4�j����
�^��1�A���b��E��̬}��|��H�����0��	������9�x��X�0: )lOD
�KT�ì�w�T�J� �sp�'�TU���+�DD�1TT���[>Xe�D�9?T%��)+�Q�A)�Zg�;P�[1jU�@��I��5�.OD�8���h�P��խL�_UܽCcP�@��͎.�J��b�*V<;��'ҧs��#�H�	!�5�U���*4�?�pV�b�?�.%��0Z��X�4:y{"�ڟ	�~VG��,S:]
�<�U�ߤ��g�*�2x�d��:*���I^�d����+����'��>���#�7��H�ܮu�ޠ��C]u1�l�t���G��'�(7a{�*��}�19g�ؗW�쌳��D��y�i�w��#<!��O�/��Y�!�t�L�m�{���ST�
s�8�jSM�PټB�	�?���,��C64�:s�jM����׭<w��qf�S�|4L{�c]�b"��:��\T,C�	�i��@ ����6͘�bZ���6^f0��CFY�)��<c	]�Br�	�B�����U Y�<�v��-�!1r�L�<Szeʀ	]V�<I4�p��@�A�U3Ut�D��J�<!���  ���!Z.��|�T��A�<9�kA9g�J�s��(2@=ʣ��z�<)��?a�pX9 ��*U��!B[�<�v�A�<8��ZSG�.�ʘ����V�<�bE�#T�j���O�806L0���^R�<����`C�ţ�
�5�̠ä�B�<)�"��k�P�9�E��-�mpF@�<���X�N��� &ׄ�@(��Xb�<	�*&c���e&xP� �G�<� O[]+L�Bf V 8��3U��Z�<9���!������O��t�aZ~�<!�*�7h�4�g��dǲ��NA�<	Pi�j	LCe�YQ�%�H�@�<ArER�0t�ܡ�!@�.�m��z�<������nx�i�>�jTq��\t�<�R�2eC*�{�/�R=��X��n�<�'��WLy��=+
�1r "T��	BKɫe{�)���f�P{`�;D���F�fR��Ef9#��@�S�&D�����ۼ^��tqD��4V1A�2D��q�D]�Pyd˵$�+�B�:D�+D���!�@:��0��HT�0�H(D�P�c��P�N�*�Η�C��Qw�2D��J�#��rtQ�b�+OD�<a�:D�@2�D�C��#��G���B�,:D�@y#`��t>mh�gN�|���*ǎ9D�Ԩ6��!�4��JM���`�f9D�� �5�����QZ/݄DZ���"Opt�#�35��	w.ɔT-H r"O(�"$��	lL�$�[#H50$"O�	��W
7u@�3�kD�@�T"O2���"FS� ���@�dXQE"O !oU�D�'�Ⱦs��X* "OT�:Ff���ȉd����"O8T9@�� �ġa�"���"O����&��}���@�S�s�Z�s�"O1����.�q��E�F)J�"O&e��	�Z
�Q[£Ǐ?��1"Or����=$H�#����F�`%�t"OBeS��ӫ��8V�	�C�n�"O(Qh�1�~aS�+�$d�x���"Of	ɕ�̺h�dH��%f��"O�@ȁ����֨��CW+�L�"O�aG(T7n �K��àl��B "O��a -��8��q//r�V"O�l�c垞!zR�3�M�aՐ�"O�!� C��k�(�A�Q�&D�D"O��^ �j���^Yڰ�"O�!'B����Ȅ-S�K��A"O"�aaXU:���m��>��e"OD�bC��
���I��;_��"O�kg�
5&DP�I�8i�"O��J�f� "E:S������Y0"O��A�	�RW,�맩�1-�`�"O�`�FX2o�����gS�)��!�G"O�x�t�J1q��"��X�d���'��%��+�R�`QI���0�'x�"�ڥ4O�1,Ҿ>
ZE��'�.eZ�j&WnJ�9��/>�J���'yHl�#�L9b����Ŕ;<z��+�'�N��.VS�^��G�#9�V�I
�'�~���h7m��|q́�>�,�1�'��w�Qei�I���%1v����'-T���n;FKX<P�Z�R�Z�'# 10S(_*j�kWeW4NL���'.H�F�!h�pegn�?l`��'G
���I�m�F[Fl�*'��#�'Wb�%�߇S�T�dH
�i�"E:	�'kZ@rw�%��@D�C�s#����'���УO\�.�lx�Β9p��$��'d���.��	(x�`�G�=�
Ւ�'�\LQA��l��4"D�/:4�8��'^�@i'�N�/��%"��܇5�
@�'������Xb
})#N�3,��q�'R�bI�1XHi��]�.>�Ɉ�'��h�FH��?0���\�����'s~tQF�
&wiB	��m�$P�������*��)*m�o]*��p�P&.�!�D[�c����o�+G|�2#�5.�!���dHl��j��\��a�k̑IK!��&ytֵE�S�_�a�TDT$�!�DA��9��އ9k޹�q"�?&!��#�J�$��:HUX��b��V!�DL<�.������/�����i!��f��{7��@�de#'��5K�!��2D7�}�EC�&<�Z���E��~�!��<H��en�7��m�U�m!�ď&e�Qq�B�<T#�X��
�e!��HJ���F;zr�x�cP��!�$U5'�1� Jjo��ҩĭ)@!�$?[E�8��g��y�����N͝F!!�� 4�ʖ�
>m1
�x�J�,� �I�"O���j��J� �3�G�>�D�§"O�iҗ�X����G
1�`����Iu���	��&
�����W��ECb�V'!�d���Zx��dC�R����g(�!�d�
�4\s��M�4���fN/L�!�$بs�`�,�6�@Ec4�P�]�!�d��O��h& X�G��E���8/�!���ʪ0(0,��r���J��Ҥ�!�����'�
�V�z1`i�!5�!��s.����O%Y�F@���U�	�!�߻��x��ށz͜Yxa�R1k�!���B��h��ޯ,X���9k!�	4r��3G.�5j��	��!2{!���a��8c*��:YR q�
"Fl!��o>XT�T :��!+��W ^!� ,r쵚@�N�@��1dˏ_!��@&�`��n��1(ZA��h�=6X!�V aw(qc�,ԅ3q'��!�Ps��S���T���oZ	�!�d�Z�f'��!��aSU@�[�!�$�2>�P0�0�/N��A1ae!��O�E��B4̘,i� ^7(:����"O6������O�ب!�Yi,�$��"OL�!hG�k�n�yŨ̬w�D�:�"O���a�W�*HE��҄%"O Q{ӌى\�,$C�M9~�>ŘV"OrQ;W��*H~|��q�.-�-H"O"�1�&7O�PjU��%�6L�"O�Hy�%՟z��4	Rˊpڦ��"O�I�v�ڬA�&9��J^���"Ox�6��o�~e�b������F"O�9� b��F$0�U�2��\��"O4X"%E�lԮ�3.Ǝ�2�i�"O8ŋ��NG���GB4���"Ov�J'f�qnD�F����I�"O�z��´��`R=6����"O��0�;�|P9�[)",X��0"Om����tm��Ԭ�;��U+v"O�% "�˅��m�	��l�"OHM�懌(��j��FG�bF!��y!���w�l��7�=�a|��|�#yUD9�B�?q��-�`H�y"�бad�  k�,3�|]9ceˮ�y�ś%�p� ���(U��(�A%�y2��M�V� Aj��k��Uң���y�Ʈ��!%' i~��뒋6�y2�]nAi����c�N��b�U��yR��Y ��T̀?/��Xy��
+�y��M)&8�X��O4s�̈�y� �*;[|�0�U�n`bwo��yB�O�AȾ����T�
3Hy��+3�y2e_&i��8z`m\�{��)c���yb.�8]��Me��f�2�
SG���yR�\<}6�@��?6�y ��%�y��3����)��t  B��yBA�b�j�Cu*�4�S��N��y���[p�9�&��fP[�N���y�ǘ����(�a�H��:!��yr�Ɨv��� �;=8�}���V;�y��3��� �i�#,���˥+݁�ybA'=X��5@�=�8���G��yrj�	l&��&L+}s�y���yrui��w8��*V(���p?q�O� ���Z"kY��Y��дY��9�"OV�ڦ�͛?|Պ�C�
* ��"O.I���J�V�%C�#�>\��A�"O���k�,"�x� �$
X�+W"O�\�Ǣ\�3��tC���*ɜ}3a"OJ�;f��XJ���2D�ih��Q"OXq��f���p�A!r��Y�"O
T����"�N��$E�5a���"OT��P���z:(�I��QU�h��1"O8�`$��=i��\4u���"OL���艥L������^ ,�a;�"O>��p�L�\g�i����@�)�"O�	�g��Q�X�36�h�!p�"O� #^�ZG��3 y�b��"O����(Q!�`M`q�E�ش�`"O�$�'!�A���"�!~�y�"O��Xv˝Tb�`�p!�P��9#2"O�I�� �:>�,�!�	h��x��"O|H�*?B�p��b V�2�"O�Qs��!���V��!��Y "OQ�2��'�쭁 ��,_�� g"O��`�ǅ�0����A��&дx3Q"OĤ$�ׂ?�Lz�LQ�*����a"Ob� ��x��Tp���X;���"O<AY'�T3hX�dx$���f1�P3�"O�M�OM#��� �'��+ hi�&"O��!�FYF��;�E�.5ٖ"OT� �C�-����&W\��"O�CEj��T��j!/��@�D�3"O<qb��#LŦ�"�nC�v`��"O�h��^�N��B�]��� s"O�z�$�&GS&�Y�KށE��2�"OR 2󋈾`��d럊,}3�"Ov}�0K� En�x���{�xyYA"O��IwE�=D�,="�����E�!"O��iS�s%�� ��^,z�(�"O�3 h 0i�Д7cO���e�"O�ع@C)#0TŪUG��p��!"OP�٠�ы�HJ`F7n���;�"O��� ܛ$��$�T�Hx��!�"O�ݻ�C
,{��I��.�"i��m+�"O.)�t�s��(1G�?X�2��"O$��ɒhI��r�K �8� �p"O*lhe�͊Z��eH�o�
@�9��"O<��N9L���j6ُ@+&$�&"Oz�pl��n�Њ%�¹}6��"OX�2���Y ֌
siѰf����S"O�$
�Aڒ{��|0`"���"Oā�P\8j�	��ሏ�h0�d"O\�������n��$�s3"O�����D��\Y��NI��s"O¥��E���:��_�%���"OXDY�%�(:��-soO 9�T*4"O�5cK�H�Ҍ ����(�m3"O�嘕��?�^�tOګCfH5��"Oh���IC
W�1��@"d��"O�p5�T�/	l�:Ө�� �"O�Xf I}�<4	�g�O�2Yrd"O���DaB���z����C���!U"O�B�!'&�c��$z|1(B"O�l ���	ca�)r̊���T"O�I#W��9W�R�ӄ텃����"OF�1�l�T�n�%�����"Oj`IE���̼�X�BԨYz��"O� ������3z`�H�qcC	���"O.�aw�ʡ(�+���_� ��"O��FBL_��QP+ɰG��a��"O
 	�B?�ĐuiD�c�XI�"O4l�6�@�.Mx]X@/�=VI�@"O8�x2�P�F��!QM��Y� 5�"O�(���A���땟%̌Ej"O�0��<�9��,��ȯ�yD˄�`���MD�Y�h��I�#�y��I�E�~X�#�T��prД�y2��|q���T�4u9�t !�D��y�-L)Y&���e�7��m��W �y���Hk�uB^{���$	 �y�X:c`Бh�A-		6=q�F%�y�h�m՘<�R���-��l
d��y�"I��BU��9}\��*C��7�y�J���tEJ�(t�D#�I!�y�Nn��@ '�'rO:4�r
���y�3`
�L��Ϊf$s2
��yb��*;,��J �`"(B�i[��y�KA�J���V�b�����I�;�yrlҖ(�x|��ȋ9X봴����y2*6K|:���BM�?����,��yr��"{~(ەl=m�\�r*��y"+�,2 6� ���%c��QAG�y��A�:d�9��_�f!Ӂ����y«A ,(���*ǺP�ȴ:�a��y�CH;/��ق�Ԭ(`q��j��y�ǝ���Xw��#�XH[�����y��ϛar�����{ؼ���F��Py��Kԉ�W)դk�H��[�<i3�ч3�� e�J���E��S�<�eo�) �n	���L�T�@a?T�4�G�O"��8��)A��A��#!D�<�u�Z�疝pʅAФ�#!D��H&)FK�P��P V��"*D�*2���\U�$9PiΑiX�Cj)D����րd��� �o#7��Bֆ(D��(�6q����
�_��IQ�8D��B�� �f5 c>v�����i3D�h(�Rl�TP�ڪ	�8L�R$D�Hsg+&��$�e��1 ah�
G"D�`�����;�%�R 
Su�%k��?D��c#��6�����L�y��>D��swI ITZ�Mިa���i��&D��rŃ��Lp�Ы/A�5�`ш��$D�zD��K�Ⱥ�(�=:ƈ�;e -D�,��o�3, �H5��C~Z1��9D�(��h�%3�޵���<�4Qx��2D���rm�6����'kY;>i�/D���#�.&�HjS�-	Z���(D���SE_�X��dI�f V$�m�+4D�h`!�ߍ%�����2T+�ءF�3D�D�($�%�+ɺ?X�̸p5D��	���
�����Z-|��rU*3D�$��#��'�<%��D�.�D���n0D�$ke�ȽR�Fp�0��G����k.D���E�PTX �G���b����6�-D��A 	�?K0\ �(J�ts����c,D��	݊r���8��U?S)�m+b)D���B�^�:>��Ժ��	2�'D�����/5���k�0?cz�kF%D��T
T�<DM�VMʒjA8�3��8D��Ça�o~��1��A:�L�q�:D�� Z�� �_�i=ԁ�"!|T�Y�"O\	��?"�z25"]�fE
m�3"O�0p�&E�A}�1P��Ύ+�01"O�*R�M}0�j�!\�}� ��"OTdf�5AP@mR�ÈW�D=:�"O ����4�d�K%�<� b"O�`��Kґ!�$e���T$��x��"O��3*��H�h�A�	�H��Q�3"O��"��^-n���YOF-+�"O�,�bBW�N`񠮆�wK܈��"O6HksB��D���G�nCH�6"O���,�:<���l�*1U"O��v�K��J1�&�H��\��"O�ГaB3����I�%f6I�t"O�)0K�V(@�!���m�x01�"O�5;��R?�q�07��1�"OH��5N�'`V���;fj�,X
�'�� x��Bm��,9E؉+���
�'\h`�G�9Q^Y��c�3 � ��'�`��$D|U��(�C�J�'�<9�E�':F��+g�,��`�'�pؒF��-U�+�%�"#t0<��'#$QS��[&[�.)F�k�t�k�'8�E�U�U�tƊK�y���'&|��m�aI���X't�B���'v"$b�搭}~�Xv��v��	�']�ĻBn�	�¡�U���bVؑ��'::��AS�, jI%T&D�r�',ƭ�V��l-�Xu�N
PO����'Ր��#Ͼ�3b³O��<z	�'��m!�j9�
d��˳?�8�	�'^��[g�F�oF4l(wgҜv�~݆ȓp�P5C�%xB��#1���A��l��zh
]pl��lJF-���X��Ň�C�&�@AZ+�����.ɖk��B剤�n�F��4NSr=��m�.p�C�ɕy.��� gK�C,p����gP�C��!gjt�`A�&|heE��lC�I<<9���n�;�>�7�_�d�B䉓iP9xw�!��P0SG]d�B�	�+P�}�%�U�R�,�b��B�	�pԥ7,�96�\��V�e�B�+k��a�2���ep ������NB�I�U�.���P<Ҵ�H�f��+�$B�	����]�S��Uzd	�c6B�� 7��xc��^B�~�"Ƀ�cG�C���@��ym0�!G"_܂C䉇!~��oTv�Uf�ZH�C�I$C�J�;���@J���D�١5O�B�	�Ilp�g�2���e-�#;/
C�	�#��h���"*)���.�8�B䉭L��9���"_3`�ċR��B�	)��#�'ڬ%q2��Sa�)��B䉷�Ԉᷫ�*{��tHJQ+��B�	b�m�W��8��4�	ۯb�C�I.F9h�h���9��q�D��N��C��>x��$� -��*A�q�	�#s��C�I��(}[ī�]���T$�![(rC�	�(f,��|����/��wdB�I�t��ڡ(s��2Ӗ{��C�I,V�����8��Xp�O�J��C�	�^d�)U�#��"�� ]���0?фo�-פ���M���a�s��t�<���҈G�|�҅ܓ�0`�"�p�<� ��I$�ߚyw�4�D�&"22:�"O�%��ՠؐh�b
]�0"O��)���w�^�)f�\� Ӥ�8T"O��T�	�^T�9��"��{f�	�O���e�	#�였��ޠSf ���'�
��gS=X�(��`ьJ7�{�'7Ĝ�ӧ�(���i*+B)��'�4���9�x��)�$"�9	�'���3�۔H��!N_/	��p�	�'<&,ۓ�� �b�f%R��5��'^�U�aã.EbP�G3BXTq{�'E�T�JA1@�9 ���6��q�'�ΔȁHԭS Q�#�n[�'7dI���^hxs���P	�'�.�r� ɁXHT�+H��(L�h�'$�qYƬۢp�"�z��%���@�<�QG�	��<����j��Ԡ"�c�<��!$|��0�
�z�f�p7�]�<y��R�S�� 4��N�<���d\�<ËU�V`�#D@4Md nY�<Y��D���!��l{�] ��HX�<F�בt�����51�X�dQ�<���6x�M�uH)l�d��7��x�<�%J��>����ċ�;3�C
l�<���Y4z��Dn
�K���bD�Q��y"���%�z=��J��ɘM3t���y2%�:8��B o�s�UXI̐�yr�aBE��ā��4X�.��y�d�p��Y>�Y��W"F�=�ȓ&{� G�/dC�0S�lK)&�f���e�2��_��n��7m�
�p��,b�,٧N��f:�� NW�bX\��	ϟ�����C�}R�n��i���rrB_{��O��=�}��cw�p��Kp����!^|�<Y��0d�D�!��6H����I w�<��͕$�ڝږEK�G�By0p�[�<��N(f�>R�N#O��S��]~�<ٕ�ՐO�A+pKC�b�\�cWR�<!0�I�M�:��1���|�R͡a%��T��\����+?��I!)��Y�¥B�i��$�Ŭ�N�'a���94�˴&��w��8ǌ/�yBѽ'o<����A,ı*�,�9�y"%�O��(#��:ݺȁ�*�y2KN*\�~���%�*���p��yb���\���&���ġ*@'��x1x3>�9�늕	T,�҄�R[�0��*n��e�c"M�%��C������d5�S�O���05O��c����4M�7"O�����;}�4�0��6s���sF"O�� �#�?.H诏B0d
���U�<� �4$4Ѩ��7�Xr�,Gj�<)��Bl�*�!����D��`\p���hO�'ca\E�f�:n),1�ƩɸS��ؖ'o��'/��$+��a�.%���v(�:��zR��A�<�'�:A�@�9e�[#@�y���A�<1�b�<&lj�
#7���i�<��B��1�Nh���R
��%�d�<��O�� �B�Ύ�|0ش�%a�<�� �P��©��"�\�ro�^�'�?)YC�ŪTJ�<Qw�H,c�
hz��,�d�O���<�����k����J?i�1Qj9"��1;�D%D�0롂U�v��(��Y�e&�`�"D�t�aG�<4��h1j�w$Q�
<D�`Yh[�RDIQ��
!H���m%D�� @�����g�V�3t�Q>.� �"O4�:�oN�[D�I*!�XC���b��|��'�t���l@&1:�kIe���1�'����%��3K�2H�nFX��J
�'��9���S�n웅g�K�"�{�'T�H9�ƠK�d��%F��6��}A�'�Fј��>zƬh;U�9.���"�'D�<�rB��?SDT��G���Ti!
�'M��s�͏?������6ظpH�'5�k4��h��(��.ۋpA�P		�'O萲����ڪ�2�@�<i$��'t���E����2Cۚ1ܭ
�'"�����0 9TXA�+"����'R���sfЬrܱK'U���`i�'	2@�Pϝ=�B"a_!D�ȡ��'5�-����N+�̬f
�}�	�'��37�*x&��#�^4	��в	�'
|��f5X�"�xCX�z��'.�	���:Z���b��Cjt���'M4!I&cäu�DyҌ�=5���	�'cq(�*�0��P��у/�T���'jD�� �p���j:*G���'e4����:H�\��t��7%��`�/O�=q���z����H�}�ȺN�w�h0{�/D�8�B��izr5���KK\\��N-|O�c���D���+!vXٔ��=c%d��*D�h��k��j��B��3s&����)D��X�`�'!:0("�����Q)&D�SħS�S[��[4�N��!Yҏ6D���D�;<a� ��E�|#�=���OT�=����,7��'f�*P�:��th�Ȗ�L��l�*!���p���F�_.�0Q�!��!��5n�mbfK	��Hyr
��o�!�d F� �£�@$l�0�kb*V8Jk!��S�F�J������\�1p���ZZ!�Ƕ[���"�M�7s�b�@�ʊ8Z!���2�6�;kJ�V�ڴ��O��i���'�
uY��ɝhϠ��W��9����'z!�Ğ�W,�B�ˏ$/x����8!��0va"�J�ԇ]p8��+B�H!���.��U���>2��a���|5!�$ێ� ���_mҦ����O�!�� %�:�k��>�D�sr!�ב?���Jr�7�(��K!mM��P:!����7X�����^�WP��0?���׿d+@���A|
��6�Ay"�)�'E���R4+�	q%L��ES�:C��`��:�C&?�V��遌xc`T�ȓRsT� H!x͘���l�Z��D��IIZ�:G��jC�����F�DrN���e��=�5A�C�u��.K/�����.	Yש�3��0�%��:��(�'�ў�Fx�&c��ҡ�
�����K��yR�1���A@�<3B��v&���y���g����-
��Zf�
��y�-N�[l�;'/֛nG�)��'��y�`�F:N; A�<�p(+��-�yR��,70�j�W�;g��(�.ɿ�y���;U�ȍ���(. ɤ���y�>A��Ƀ��4�&���g��y"%�)I��37nH�1%��+��#�yR�¾�R@�5�W9S����'���y2S�0�ؕ��X$E����"���y��[�h<\U�$aX9>�x1K��y
� ��	�mW�Ex�Az X�
rZ��B�|�'az����`D㊛O܍���@��y�_�0�b6�$|��I҆���hOq�
(	Ƭ�%/T��O����=�"O@ݛ�'6�H�p��Lp~��"O�E{t�]�_��tҕ��-B](�r�"O2ap!Â-V�K3�VN$�+""O��X7A�lӀ��YB�-���|b�'���#5J���O�9����6͐��!�CoI fFw�`@�Q�߼ y��I��(�L�Q�/�(D���p"�y�"Op����_ ���JˑEW8̐�"O\Dk�iU�qz0<a&I8r���*�"O5�Ί�P@����ҁb���'�:����{�&�ZG�2]�B)C�'�2���N�Ԝ�f��7V����/O��=E�䀪�f\��MU.1F�P����?���?��<�š�&EvL\�p�F&'j�{i�Z�<A���iX<��FOА)��I��K�<�Ӛ34�J��V�fPb���E�<�D��$-\��D��xU��"�Ln���?��o\XGJm\�pV��1N��5��ئ�C�mצW��X��,+�PA�ȓW��	�茳3�% VD�Gt���ȓOT�!��*B�JaL���VNm^؄ȓ)'�P�sB�r�H����KѺ��K}T�Z(���Eg��~�21��Ӓ'*�<�x�J�+[%O�2t���O�=E���/U8L#��7D���'�өQ5�'ў�>}8p
�=l�!Э[b:H4�L7D�x���KB�Z8T-E,hFLs66D��DJQE<b�ȠJ�C�Zh��2D�`��e[&�p�d�U�^�)�,3D��!B�.tY���F��$A,D�p
�呠n���i��Yʨ��$��O|�O����O��=yd�P$O�B��4L^"��}h#���?i���'p��`��ǲ�̜�`�L"]�ȓe�n��#�,hkn4diE;1��ȅȓs�D�qp���L�.�{��S6���ȓ�|\�ĤٝZ�x\suK�1{ؑ��9�.�A�g;�<u�G�ǖW1>��P<��'��"֖}k2쐎n_>�ȓ�������B�Q�"�(�H��'*�':�\"��O�1�&����hR�'��Y�t^�0�4�#���"�
�'�P�0N��_(�٣�N��y��Az�i��t���F!!�y�Gb��å��
w���K���y��H:\Y�)R��'p_��TbL1�ynH�t;e�Y�dlL��!f���y"
P��YeÖ,XZ`�Å��y��!
�h�x1��Wդ�3B*ׯ�y�	W1�s� '^�^0�1E��y�@
tH�DلbU�XO<`Q�+�yb`���lp�G�D�U�`�����y"�ʭ%H��[�K�29G�9��F�7�y�l�f�N=�E�]?,�	q���y��'c\�8j��B�bF�S!=�y҈
fi�x���tI.(á�R�yr�˨@C�9u�<j��Z�"V�y�A].����2FJ�`�@1���yb셍c��P:�(��-6��HK��yr+�1�R�`����$*~�"L��y��D!2�]a!+�$0LHM"QJ�y
� ��I֏
��3G\� ~h�0��'��3)J�9���P��8�e��g��B��%k<(�14���壌7"�C�I���ۀ"A�a�
��d��7g�B�I�wj�J�<MµJ1,�7@�B�;�*�y��(@�U	D�)c�C䉵D�@��h`�!�ʈk���H��	�j�2����Bw�B�T�J� ��B�I�'�����bv�9x7K�,���ȓaF$��B��<r�S&��t��8���pQ�F�D�����'�ń�	;��+b�8g!�ӫ7/*U�ʓ*�‡G�F�8�ird�<D�jB�ɑ*R� � W�&+8�0��1�VB�	)o�U�!)]3K���	1GđQ�����O�a0��ׯ$ʆ)W'��X6 D��%/�*B���aL�;'Ф�;D�,I��Ʃy��"�F\o���b�i$D�a�N� s�����3W\ Z�K'D�(Zq��+R�` �B�6"#X��� D��%�3/"<�p7-��S��	)D��"�a��W�@1/I	����%�O��D�O���F�1/d���T�G6`n~���&!D�����$=Ob�hA��99�n���,?D�\˓B�M�� Q)��m$X4�w9D�,Q���T��]���V^F0�D�!D���o�`�v\�ec3r��*6� D� 	a#`���� Q)Y5p�`�D4D��P���"N����iХ9X���?�O��d�Z��	Y��^l�|+@(����C�	g��\�!_�0l.i���?P�C�ɤ��H�4��\���%��v��C�	�~�h��5,Y�A�ؘ�bB�+_�^B�ɑ�y�
��M~���j�*G	*B��$>�FMa2a��M�t�B6�*$*B�7L���O�U�&����
W����z�`;�!�(�h5k���+J��	�$=��K���T�'b�QV:qM���Ê�{5ja�u"OT=��݄>�Z4y�@�$t�:�"O����4gp"��n�E�H�"O<�*@�֨�ȑ	5M/.�6(��"OL� H�h�8��%�˃�ע$H!�$�T���7m��R�*H!�I��d�!�s���	�E,q��˦EL�N��Oz�=�+O4�jU�(�| +���80K�hs�@�OrC�		���P� ٣6kbБ�FǛb�.C�7@^6Lr!/�_�Z|�����C���̘���S�S�p�1G�Ήv�B�	�O�Lzi@:2*�8Y��L6HC�so>E����?�p�Ŋw�*C�ɥ�̔Q�G��l��T3A��=�H>����J9""��ۅ`�Z���8������$�Op��'gǚWB]q�u��C"O8�k ��g(M�sI�!j�|@�"O�I���Z�zU��)�Iy�@"Oƹ�BO�����лd
>��'Բ�s���:��L����v�1R
�'�0��Ņ�\FeP��\�h ����*��p�΄�N'2�a �@�z��'w!�d�DZ.�( I�q�9��]6W�!���9�����ƘV<��	C}!� �ᤅ[����S�^�Y���]m!�DS�L�zd��܎H���aţ o!�ʳ`�b=���'`4޸XPb�t^!�� F�J�l�]6���VO^2��9��IH>y��6L����D�Z���bv-:D�����r�ԭ��>c�ĩ�Q#;D�@3fðzD�h��K�Ab1*:D��� N�}��"�疓b좥�e�+|O��<?�4�/!(�'� ����'i�i�<a�J5�h�f"_�Nn�|�<I�ϋ"dڅ*R͟1�D��a'v�<Id�(S`��)E.��v�.}@R*�J���hO�-��̘��Ņ��YD(� ��ȓvH\m
���w�r;��QRч�Ej��y�i��֝:Ao�;Lr�1���v~b���n���G�NH@�1W��1�y��Z7f��Tb�?w>�`&.��yrO>s+j��昤8a4݋e�;�yR ��	�nX�F�ڠ[�����?���0|"�$֣z�tQh�" �@��5`�I�<Y�l���x�Z`JA�(:�M���Q�<ђ�29*F�[`eڜP��x#Du�<q�J \�\�yA OH��IS�z�<�#���D0.�HU��3A���f�u�<E�Ń>�	��%4��rA�^����?9���O��2S�8"��Y�H��y�J!�DL�@! D�|}̘�rmU}8!�$RSG�Yd�r
x<��L��x�!򤀉f!01� Eי#M�r��<(�!�D/�dH2MD&=��lS���Rv!�Q�2����J�*
,"�FО1S!�-}>�`K���u&
�Ge!��Iy�ԉ�� �M�BdΟ6!�d��zU��wD�ٔ��:�!�_I����ŕ���h� ٶX[!�$�+�p�	��Att0��
�8^!򄜚R�(=�Q��xT8��f���!�d�F��)�cO/-�� ��Zk�!��úq�>@a�	�	[�`:��*m����#?(��G��="��D��\f�B�ɉj�v�Z��[�sVD�T�,�B�ɟ\&}��.ٔT��Ce[V��$Åa�M!��)�¨�!fĀ:(�'vў�>y+�&Q&eF`k�ɚ�`�R8y�a#D��5D�Xb��T+��u���qN.D���C
Ō6�Z):F��&~�����L+D��+�]��D"�RYpƁ1�.D�����N�8o���ǐ�G>Hr��+D��H���5Zz,Z�jN�~wE��3D������s$e��J�@��q %��9�S�'A�荛aa\2R!8l�5H�2�̵��~8��(�(T��X]:R	�6B�ȓ�h�uʉ��n�(���*$fŇ�S��p׭�N�������7�ɇȓ.�⁹7�G�!�D�
��(��`��c��İg�F�.�t��˷Mg���ȓ;*i$����԰�C5'#'���IS�Sܧ=|��J�g�.����l��ȓU���0���+k�D�4��TqBh�ȓ	F��+/�<p���4"4~5�ȓ%�ؐ�g,�;^�$H҄%M%�����;1"���Z������T$\��h�ȓ;�Ȩ��KX��X�▥״st������Cɸz�@��!E��q29&��$�@��m�O�,;%��2�TAy��ջX_,��'0�1ѕ�C���3-9ϐm��'S`�i��S������!<ޖ�B
��� ����A�|����bT�
�3"O��A�ӤI>~���V�O�%�"O*X���3M���Q�^�Y4q�"O���6.��"rؔ�Cb]i�l��u��m�'���9g	߯@ޤ��C�����0��"OYx옲v��(X������q "O��Z�AA�h% -��쎜G�V ��"O��k�?,(��C�ۜl|�z�"OHa򧤃�t숍+���zV��"O���"�$�p(��+
/EH�Y�d"O�	9�i565�8�aɳvA:�@���S�'u�D�I�܉g��3 \���LoRO�`�ec�urqɔ���:S"O���4�����I��]�p�	q"O�A:P�ل�F%��I_�k���2�'�ў�I�<&�T��J�y��l��M�ul�-{`�Og�<	����(�� ����"^X�<Qo˿w��� 5a�!g�Q�<��i��}��Bh�c�\*6AhB�	�K�x}0Ī�)����P�%XBB�I�/��7GB�X���Uh_�3 |B�I��m�2-ۈz`H��Aʎg�0��d�<�O��e�D���Ub��"Ӫ�q"OB�˶*?� �['����i�"O�r#Q蜄�1�_�9���"O�"C�L8��`�8���y"OZ5*t��
�h3��?ﲔ�C"O x��K/΄I䀀>Z:��9"O2Up ���x|r�+K'rf� �E�|R�'.b�'��O���<J��湊6�*����B�4P�	�'�:x���1wO�p��ʊ!ON��C	�'*�"3��n���[�OF�K��p	�'�pD�)>�<E�CP�(L��'ָTx���$���*M��d�r�'("`M&qb���g��nL�'le�A�ʅ0e�؇�ܞx��S��?Y����OJ�S�'��x��!�4A�^xa�!��E)��	�'ڲ���쓊5t]�S�C�EI�'Vf��Ej	#}Lh�n��?V�@B�'�̝��ؼ��a�*=�2H@�'@��i��χ#���%���5�$���'�T��ԍ�w��M�+K�3��"Ov�Q%*  �xP�7B>Vn�H��D&�S�I�=�֌����5o��h�ԩ3�!���!Op(�Mx%.�&ɋ�B�!�dHR |�G 
6$����Y?3�!�$�7f݆a���U���"H�^!򤝖o�h�2'��[����i.cA!�u�mi��JN��\��
cC!�$�O���QW�wh�pZ�@Ɲt5ўX���e��<	t˒�D�h��'K_>�|B�I�,#hH�7�Ù,��U"��DB�I�Rw8�#�|r�_)O:4B�	J�0�;BbJ)�P�v ���2B�I*��u��C#�)�\>(�4C�I�{V���	W�r����L#9,C�I9H���V$�K��(I��O�d|6�?щ�IS+: z��O?D��H&f�j�!�D��5k���(��eƕ"�!�E�H8p`A���aŠJ�H9�C�;y��׭��_ ��
�BC�%aG�#�-G�f���#��-�fC�ɦ"�H<���[�� TC�I6o�p�UG�
�D��w�I�T�?��� ��W%B:A h�3��ݱyL�YAD"O�1�č,�V������3D��"OЅ`��ЕM�F-��@M=!����"Opl�C��ڲw>�!���7D�k�B9g���+��b��7D����gGK�[��l��P��7D�L�Df�(�J�٥�H�@E�x�v3D�tKפ��:�SB�k�t�"	6D�<db��A��݉Uk����(��g!D��b�K���|aJ�q�r���"D��Yj��GL�%A��B�!D����=jv��a'���l�`�S�2D����]<}�⸂�dƤFJ�g�-D��cPGC =� �0���.cd \��9D���C��9�����Y9���c �8D�`���+W���&B_���ɲi5D���P���ZyI�
ԇ{��1!�@>�Ȉ�n����VWz<܂s����u�0"Ox�?Cv-��Q�L��Q���y)˘��	0�
�	����gN�#�y�HV-;�r庥��Ut�e[��O�y"j��N��W���i�y�W!-�yB��`��Ly@FU!S�q�'��y�	�\"��EL>~�ά�6b�9��'���O
��D#Ҙb��8'���BP����yRjjcuyq��&fld�qЊ��yBh�>T�<����]f�!�d����y"���v8�9ӎA�Z)���g΢�y�.�UH9cS6{8�LK�F7�yb�Sd( ���y����Dm��yr[��pe���m~�Dh�&����?)���dL܄M��J�h߼[��K���?Y�'����U�)`�ɹ���.��-*�'0B�@�fAg�C��
���'nf ��V���1AdÇ �t��'ֲ�s�4g��	�3�C%O��Q��'2D	0DŖW 40A#����Y��'ͨ���Y	M!ތ��ˏS���+H>����?açQg�	��A���fȨ���E�L���I~"d�)9�\)c�%ʁ_J:m�C�D��y���'L�:���=Y�`i��$���yҧҸk �� s
��`d�!H&C���y�C��v�R�H�`���`���y��. !,���I��/�8qеJ���yboϣh�zA+�-�D4�u� ��d ��|b�y��L*�1���\�}1�yb�;)^M��`^]l(�x�����yB�I�X�S���bM��+=�y��� ��X7�f��TQ&���y���a�$P%g۫g��x2v#P��y��r�i#$Ğp�[FJqI�ȓɔT2��C�y�f��O�D����}�$d��)Ȧn�5
 �>�
��9�ecK�%oYp���J�8aC,|�ȓv��bs � I��]�d��"4��ȓqe�%����8wT8Q!�"B=FeP�ȓ���"��Y2R	!��t�]�ȓ@
��F�RKF���%R�m�h�ȓwD��{�^'8�� [V%��6r-��Y �y�ʴ��#rE {f��ȓ���e���A�4��Տ��̄�I�֩ڵ 5��9Bd�\�0��	�ȓNӂك��:V?�hZ�ϕ�DT��[�|��#Q*�i�MǘQ�*���S�? ��"�'D�@���BL�X�a"O�����6zW�Ȫ��޼D�N���"O6���ε%�u��kQ��N�!�"O�Qi ƕ5@�� �EQ$+��ٙ�"O���ÍH&qA(�U'�B�`pq�"O&9�$��w6c��F+��'"Old�%e "�9Q�qS"Op���g����$� �5�"O a��H���3�T�P$bq"OB���M�R��M
GZ�|�b `�"O��	�����,As�D�I5�"O���N+��#T�_�e��<��"Ov�{F�2"l6�;B)C�k�*m�T"O޴Ƞ�J�>ȕ@B*��D��#s"O��CP]:� 	��(�I�HI�"ON`!�ߊS��*���=�H��R"O��ŏ�;z��I$@��XӺ�
"O������/ +���0�$����"O�%���T7y�����fRfn~4��"O>�ʠEO��
�BƳC! a"O�8#'QbN9�jܡ!Ŵ��"O&�t����V��ɳ�"O:3�b=9��(��.B(vy�Ԫ��	ϟt�'�1��tF�q���c��BQjPHCt"Oĸ�'�/l��EDH���"O�QsS�
 ��eÃY�D���"O�P��2z��usT��B�j�"O��� ��E7@���3� 5��"O\���
$Gc�xb�Ԧ�
�P"OT�q��$��0� ]�
��ȵ�'���+�Տe2����	��1d�%9��$�O���B���IP�$S���$4W B�I�tW�1�'6�j�'F�
B�"B9'�
���7�[�O7�C�I�R��ĉg�/T~�%A�AFxXC�I�9��dZUf�'��1�����>��C�ɹ*����t�\�=10����Q�zB�	WR��ضM�N%"�i���#H�B��Dl�l������YWϠe[~�K3�'D�pQ���p9���L=}NL	f%:<O�"<q ����'�=g��MR�� [�<�B&��{��q!b�_���r�j�U�<��nY
��0CAM���@���y��V	,������4��T�"3�?����h����%��B�R/_�b�j&$�?4�}����a,��#�\��d�N"���C/D�$j�*�?�} �o
.�m8��2D�k�`�^�̨+YD��)Ƅ#D�h���֜ua4�Z��pI��;D��F�0x.^m����YY�U�d�8D���/_mj8&�	%��q��<YH>Q���O$��D�b (�'�An|����'R�I :���I"O�aG�m2EA�2EC�ɺ@x��������v� 2�?a����#;�H}Qg&$�i����I�!�䞨w��*'�<y�,L�Ҋ�q!�D�t��$�fc�9��ثA@�y4!��0��n�u��<���Μf�"�'/�'+�>���l�����W2r�\��@O�t�0B��Eh��5��I�)���:�*B�	�K��b� � 9�"${r.
�btz��8�I��G{2@ѓ.D��G�h�(�ZW�B:!�D�VG�,�G��$���� �-!�d��Q�����,xpnH3Chȅ�!�� �e��L�FҤ	�+�� Ja"O`�@��C�$���r���}�$i0#"O�qya��MR24k삠�(���'z��'N�ɱp�b����H߇T�#��',axb-��W�}�D�]�V�x���Z��y�����e;���P,d��g�ǭ�y���z^d��� ٿOZ����	D��y�lQ�!��b�K��5�j�a4��!�y2��[9�3�W��PTsc�+�y�Ѿ�s'�Q
�Ε�!����2�O���bQ�t�f�0��<(��Sc"O�C�i�!�h `Uм`�>�4"O��X�f�=�
$�0���	r�!HE"O���J�v�4rd�kLԺ%"O2�9��?�"͓"��Se�T�"Oxe'ǋ^�n���S/XyA�"OJi��&��T�f�t
��K"l@�X�D��	�8��B����x���qs�A�4�C�h|��� g���x�Ã�$C䉼qI�P����喍��CƶG|�B���YcGIP
�fq�5A��B�	"h���Em_�3�(�Z/�)�C�Y-���f��:8 c��-�vC�	2�(݂f*X5/�Ӆ��n�2B�ɎZ�h!c�:Mb�$+b�2"B�I ���+��ݾ��ISu�d�B�I�{IZ$1�&o]��{����C�%9���V�F��e�`"� \�zC�|�X Ggj�N5��۫+�PC�ɒP��C&��5�2M��Y��B�I���Y*�Ʌ�欣�?A�<B䉆c[x�e-���s6�¤	<B��6����G����C�E��tJC�	�#Gi'jbx�KEᐐ!e.C��	)V�XFX�Q��i�Ȑ�`,C��^�h@q�I!;�¬#W!ٴ}�C�I�>Nl	�`�4����LH��yb��#�.=A�$%{r�,��Cގ�y2���v��*m�>���ز�yr��WZ�A�b��3��(�0O�9�y�ŏ1-8j܊QȀ�Ɛ�5�א�yr%�T���K�h�՘d�Ϝ�y"�G�H� ���`+2�z�M�'�y�#��P[���F������"D����,PK4��q�qU�y��	�0(��h�-�&lxQ�N;�yRd�	#�9!�F.1RDp��5�y�II����j�n�'�e�p�˙�y�\�i�q�Ug֯z��X`�A��y�
�3{�iq�H�<	v�QcN���y��O��z)#>Tx]�rL�6�yB�Ha��݁5
�N����
��ybl~�8|�䌝�?C��	ՀE1�y�T�X\FՋc�PE�4�d����y���\G�@yu�?DL]����y�Jt��� ��.1�������ybnZ ]C�l;�Ӫ�΅:�.9�y��ΠQ��yw)�}�&���yraܙ%����c5���F��0�y"�ʌv�B�Kq����^i��ۍ�y�LQ����+Z�W�j=#�n+�y�B'OP"���m� WP�p5H-�y�B�q���E�pTX0��y"΋:Yj�D�Pl�(<����*��y
� �lz���/䀢�ŉ�T*"O�12�C&o�`��`c� w��YBT"O�4R�T�Z��uxw�ތth��&"O�x��]=Ib����֐����e�<����	5�a�e���Y(����y�<9��)+6�xa0%��k
J���c�l�<�F"(h��5� ���x5v���$i�<�@d��H��ܑF'�"�#։�M�<�[+0�4PBခƀpsEƖH�<�P`Ls�����ʢ�l�{ �D�<A��G)�%�AB��F��"�A�<Ѡ-C8U@y�q�ɾO�r !hM{�<���1��pa&Ȁ�1Й굋m�<�v�O*GV�;q��0r�
 ��M�<��?t0-����K��m�+W�<q��.- d��hȩ9��@��B�<!�A�>3���KA��jn��zpk��<�`�a5���W�ݧ"~�ҦD�|�<�Z$~:.���s&YBծ|�<Q��4�xe-N�
�|͢eLC�<�a@2�u�$ꍀg�,TzwB}�<��oB�:��Qi%-k�pb�Ey�<��U5!�d���S�{��i�C|�<��B� b9��Ν�At��F�^�<�4�@2V\��"Ӝa!Lh� g�E�<Ih2����G=�!6��D�<�5�R�A8��{���<N���PP��B�<��EB�A�7aҴY�^U�<�%�(%@��Hs.A63�>�H5�CP�<��>8'�� ��&t{ �H�L�<��a�NkH��h�"u�>�s��OE�<�Q��'vb���l�"	2ܓ��e�<)�� �?q���(A�րYa�[�<�`l��(ؾ5\4\Bth�Y�<1��K���RB�T�>�+���A�<�E��v��Qa.S5h�@H���]@�<I���1岬k�n5!
�|b4��~�<A5k�>nE�e��R1f��(:�~�<��-m�����F��-l�c�%u�<d@���r�C��TB�r��l�<q	�-oR:�A�酿c����@�e�<q�)�xFJ4R�� ��������`�<9Ԉ���	`P��F&��ֈ�E�<!#��$Q＄�c)��<� �h	@�<�rD��&#����;Ș���a�<q�A�L60PS⍞8��1��M�T�<�.�	�9 B/�;�ݫ�)�i�<��B�1�� � ��%"�+d�J�<�'c����2 �P,E��Y� ��]�<�V��(�e9 �ϼY��r�<���݃U攠#�KK�\��b���w�<qv��3^�\a�T��>�v� c��<)2O[�{�
abFďtr2��`Lt�<I��T/D�|��F�D�
�@�&�Y�<���"���H!k��U"�遅W�<�T�L ���ll��EלYlA�ȓ%ff�0�ߡ#��uq&�ʢh{�����(it��y�ެ:�ܵQ���ȓho慡"�"��� ��/?�����N�d�X���"����!�\���I����ւK��mK"�#VX�ȓPR����.��{��k��٠R�5�ȓ%���J��$%R��
�L�`�ȓW^(p�ѿel�ч���xP��S�? �@�iWrE���Ҝ1���`"O���O�4�xqC��L�HX"OV�����\x̹#Q�ܧ3�E��"O���f�#Z,�Р%�'�>�0q"OFB"/�5^�d�h�F�!z��E�""O����A8Jt�X��%�)|���x�"Oz����vZ,jQ�������"O����$J�2< ���V��"O�C"j�@�vQ���J0\a`"Oz�q��5}��!q��BA4Dc"O�0�(����i�ЍN�2F�s�"O�X�El���5fJ�'<�0"O
�8��H�^r�y�B�s)��'"O.�P�惙_���z�а��W"O���L(>p �B�%�|Ը�"O҄��/˘u2El1�䤀�"O �:�D+jԬ���d�� @�"O6I	�Ș]t\��$�łe�����"O��؄�Ѐb⦠K�CF;����"Oz�3D�D�)������"�x��t"O|��g���j�.�CU!T�`�"O�L)aAԸq��)�B_��(h"Oh`s��	*ot�09�O���Q��"OȀ8����1�fDa[�E�l�n"D�0��矄&��L:2A�`n�ͨ��8D�x��
Q�)��e��E䪕�D�5D�	Q�� �p�;p��	���x5O D�B�a;(�(�c�I$}JX�u�#D���E�(|D�c���C;2l�!D��ʗ��;9=d�@lA-P8P��>D� S�H۴_:�:�+��Uv���B-;D�Ȑ�N��L,�&��><��dm-T�����:$h�r�,O#2�dp4"OR�X�UF+ @���[�*B�Q؀"Oʴ����%gj��,A>���*O*aࢃ�ot�<[CG1n�%i
�'NJ��EOw�颓��\j�d
�'qb�{�������G��
�'�N�H�ʞ���X�BI:���Q�'�����i[�9��膋ƫV�Ex�'����!���s���2��#I h9	�'�:`HsbHɀ(	 nԕ?:����'*"�b���:s�h��º;vQJ�'`��X�,��2q�I�%ۈ��'�}�F+��C@\�k�@Z5#<�x�'�����mA��-�g�K�J�<x�'�2����������g˙L�Z�'��A �=\+D�Pf&�&	�Zx@�'������Gt\9v�	�|����'n1K eh~ĸ%1r	:�"�'�n�h� ϛn��H���k�4��''���tC_ 6���p� ܾgI�DS�'��as�C=:زlP�@	L\��
�'}椋Q-]��v@!�e��L�}�'(d@�.��t�ҡ!�d��K��}�'�BU��O�QmX����A�1	(ِ�'���Y���]�$��]��'�V�Ӯ�v�h� ��^4��e\���<����*H��� ���L���i�&G��}���������@��A��I+^ك�7D�HCD�\9kT�T&иul"I�i3}R�)��9v�LIq� �qWH��f��c�؄�I\�����q�ӥE�F�����a?)��P1��1�D
iC�W]�<� ��E�?W��R'��\0�!t�'>ў4�n3Wтl��N$5 ���!D�<��E�=z�t���b��I��"D��j�&B��ܨA�%%fN�x�G>�OP˓���1��_i���!��Q."(�'>R�'�x�(���*R����P���;���y�>�`�3$ -�D��?�y"퉲Dr��ᗉ	�(y�@��.���OD#~s��	#*�ؑ��,"�����D�<��eV#F�Q4g��f�+ph�}�<af�U fB�<۵�C"]�n�EX� �O>��Q�
o�Q�whۗ��݈[���� S�2e�����HP��I2���5���<�;�(�2u�$�I�e�`��&�-q85���:D�$"a��[\�E�a	�6@�8�9"�"D���@[�5��1��Y�\�ڡ��H D���gNY^����?�~T���3D�ԨQƁ#`����ޱ@�L|���0D���*W)H��)��
ۗ# ` �7
,D���ƙ.
�zE ��\��'+)D�\s�n�1g���t�V�
��*�"'D�����C� �l3C*�2 �:ykP�$��hO�S]�:�k1e�\-�8�ƊP�kb������`��J��\v�6� A-C|C"�n�ş(�?E��4q����7/�)a�����?�LFz��~�b�;mQ�Di�D�<H�
ف6�[?!P�O:��dOC��n�Ix��[E(5P��r��1O\��?���JA��P�%br��⤗pH<I$LV2?,(	�mB>� !J>.��	h��,��+����x��.&�S�A6LO�⟬z&�D�K���pL�Ȝ�S�N�>)�>ъ��wn�q� ���2[Q~���[j��&%^Ni�!�@���s��p�>�ۓ�����+��s��9K���,[�B�I'R�6�!4���{�\Q ���6Y�C�	?/����bED���$��eɘ�DUz���I$�I�n��E���4(�$��"^3�bB�I,$��I��ȞZ�K'��ŰS���4�L	Qr,@.��c�Ƚ8;f8��N?I���ϙU���� E�a��-�&�)���<)�d��NْC�L�I�.L� �d�''@8Fy�Q���F4�D$�7"�6����bO>��xB�. ]��ᇌ�S%��VA�$D��o�P��h��q����T
�+4D
=b� ��'�qO�"�O>�"�'��fȅ�t"O�Pc�	ͬ|׌ԁd�)~d���&�>ъ��)�	<����s#�'.��{���fF!�D�A5��5�Ȁuwe�592���)���`vn�*T`JD�L�~�p0/9D��`��_H��;��ؙ|�@���!x� �?1�ט'Z�S4K�:���@&�Z��ML2#���m�H&��ib�́53Xg��h#��!�v�8	1H�S�O����SnS%,��rO0uf.��'k<C�Ϲ��P� U,q�ZTA�'����Ȅ�V�Jm#�B�<��1�'�s��6�P)��A�
#|uy�'�����	 0uL
q�-o�{�����&eT-Oc4x�f	r ��#��y2荿~_nT�#%[oD���&����<�OR�Ђ�*I�����m�3.8D�(��	D���	K�1[��'�+�6ذvCN\$!�����+�C���� �0bA�1�k��ħ��I�"xRa`ff�;_�썀3'��Ɠ5*r�j� fPfru��Vٖ��	�<�5�)�~�H?��S�? h�ℏǣ\ŠMC7�C���S�'��̧>iCH�h��$�T�R� ћ�l�[y�'�Jy���'��5*膤XJ`�CU@�)b|����D#��?��ɷ1�rϒ`�$��S@�; )�U��!8���s�Ж*a\X���y��C� I�#N�E��ܐRLL���M�g�Z5���?NIt�Y�!Ewar�O�q�g���̦��Q��j���'ԛ���{���U`ި Y�yA�g�,sK�B�I"1��tS�&�)a�z8 ����G���<E��B2	 @L��ѱ`EN�T��y2�>x��sLŖ_��I`�lÌ��'�$܅�I<#�n}�fi�'	L%��e�5|ߐC�-)�H|ˇ���`�`���^%A�NC��uV�}'��9iE�� �Z�RC䉃B�ja��۝'��*v#�
yvC��3k�^tz�T+D��x2�LK���⟬E{J?����o�B�+k��^�(���:D�� d�!"�jLAS�R�J�X�{Q#7D�������J*`t ���t�v�	�A6D���U���x�TykR*�oF�tm(D�04E~�U����9XM�%D��@�e��Fpd3�eݣ{��l���"D�T��E#p��� �'r����,�$��1z�%�$��}0�Y�A�=H���p?!��܄mD��[�F%Rݓ�
y�<AA ��`� ��2k_R`��I�<9I��h�݃��	�@��(*���o�<�g 'i��xjgk�
{\z��Jk�<����(>��SSÔ��ZÔ@�<	Ď̂qp�أLN��X��c����?����:%T�a;��E�}}��3�O�X�<a�B�'6�L��gG<l����`̓ט'�0�|�JH�f�PdIp懸F��]9�/IY<��85�a�Q�p܀3cPD���'�ў"|*��-,AD��KF�΍0E��v��D{��� o������:�KebK���'���$�&
I\x��BMD�9�&O�GR!�4���2�*G*>�	i�M��!o!��ڶI7l��%�+g�RD��ƛ5���gy��'� �ca!���\��BL�4�
�'��d�`�ͪ�t|Yʈ)t�p�b��$<�S��b���&��Htb8 �jɛ�y"��]�@����%,�q���mZ�Q�Q�"~n�$2. I��ژ!�4���H�P��B�I*�v�jA�Z�rrE/��.�B�!�T��N��&��YS��h���	v؟�k�%�;9B�]��-��kM��#5D���1w��үO�=9�'�J�<��.�
"�9��K^j	.��#ꓢ蟂�3�@�$v����$9�(;�"O�l؅���.%.(z�OD�+�aЇ"ORT��oÞS;�uZP��fQ�"O� �[�v�`��P�Åh�au"Ox�Z�)ǈ{��K�%*�@}J"O���P��	4�H*����^`A�"O��GLΟAJa�s	; �h�"O�ț'30PTH%ŏy�nppE"O �qf �z,Ȅ��m_�N� �;�"O`\#�#X\4(P�ވ(b���"OR���������wϞ-T��"O�P�T�*8��i���8�<���"O�1Ɂ�7k�vd�qDH#h6bUc�"O�T�q,V���-�Y�
� �"O� �Q����4X�HJt��"3r0���"O0�pqBD�D2E�sѱII\�
�"O�L GlL�Y��M����RJ7"O��`�śH��Г�+�:^$��"O����Z�0�٠�, �2�"O��s���d� 0���(�n��"OmS�Z�&z:Uб��\~�\R�"OL���ώ�k�6	�ݳjl8��"O`�x5Ș'd��"dH�N��s�"O� K�G��d�"�� �k�V\@�"Oh��AN^��y8)^-1�<i��"O�A�a
�$��
"G��\�\H�"O�Y�W���]L	���U��P�"O�Q�EW|�P���!8,Y±"Ol:s��2_��d��I�%}���"O�Hb%*�>����e,z�x��"O�օ�Aײ�� ["l��p�"O�<���7Lr�m�`�,	�"�`�"O�	A	������Ώ�ʆ��`"Ot����DZf��\1���"O���uk�m�F���<d�p��4"O�E{�%F�Y�e��.C�f�(Ɂ"O H�#R�_u�d���ƉC�V`3�"O
���A'+���Y3$^H0��"O���gJ. ����~��Y�"O�L�"e�X��Q��F�-5bΔH�"Ozm��)VT�bd�3�W�Z	�p�"O ��Aǋ��4X�m��E�  *!"O�ya�/5$�p��6%��i����"O�=�`H�6ލ��ж�`�"O�I!`��5yC0$���Z�2���"O��b�S�)F=��I����9�"Ozi����S�ڕ*0j��A��Ը7"O� R¯ײU0��ɧI�E��tV"O��	001@�0���"2�X�"O>���Y�+�2� ��=g�T�"O�]���T6~l䱁�ѕ*{~(��"O� DȢ3fA Ӎ��`��!�"O4���D<Hf�a̙{�rܙ�"O8I�!͈�c�f���i��t�$)I�"O���c��_�����G�2p��"O&�s�B$_��=A��:X�ƕ0�"O�l�1"A�RXÀKL�[��|qu"O�4��I 4E2z��'I�����"Ot9Xc�T�s�,�y��6$�*���"O����/I�z�Icg��$���0""O���Ǚ�3 ���Gm!3*5D��;��l#��3W��v2��t�Nm�<�"M�A�"�QQ"PM����c�w�<��J"f��e�Ň�"4��x2�	Y�<�`C�8�J��U�E8�| "�c�V�<I��R�qf��IG?Pxyn_P�<�ևp�Lڦ�;?�B@[��N�<Yw.&bǘ��G��81'�L� j�R�<1�eD�GcX��%I0M)x�����A�<1((�~�S蛲�Z���&C�<9�$DOǠ*5aγ+�~a�''{�<鐏ߗa5nА��)�H��g��J�<Y�H�|,Lp$`�{�2�Q��\n�<u̖�3yl��т��T�1�G�<!��DNl�i�R��\|�<Ac�2|C�E%�	�ڨIIwL�}�<a�i �E��r�]�	i�U��";T�����Ԟ�&�q0k%c�ˤ�u��I1,B�qO?� t�9�aH:�d('��
޶��P"O�q�H�;l֌@��lJ�Q��X �Q�\#B%3+BY��Ʉg<p9@�գh�Q���P��N��$!@ȁ��,��!A��"7�s�Ԋ0���u
�'�mq�)_�y���k�͇8<�J�+���_�u�����Խ��OvĔ�K	"����s��3�����'O������9���F�� "U,���4:��B����lӧ�����UDX�z�	u�D����p<qQj]'��'#Mi$iJ�7�f�h5��\=X�OީI�ㄨ/����
ϓg�Dj�˂D�i�ᇏ�z�'�����CO�S��c��r��h�������n���x�"�=n��7H@h<��	L�q�����Y.�( !�B�W̓�<,q�b��ؘx�k�*��IN���۴H!�Qr�dH�hݤd����D<���x����ϨEMv�"w���Y�����iO�:$�:t��/��I^��M�p+ҭ���rƯ'�xy:ed������}�qO���/VU\�!���C.���c_�����4 R��'"e:�ΈO���AM��~ (�Ofe)PfÛ鸧�	ڎ|9[p�S�RO��`�*�2Mӄ�9��ʄBoRT �'&j��� O�������'j��0D�P㡎 N����5
Qt*P��p�g}�O�fI@�ƅQ-r�8cC�Lp�˓	�R��!fB�D+"�\"��$�۸D�� �R��RJ�ϓN���kĨ-�)�'$��YS �
Z�4l�J�qM���Oa�b�U��D{��;�c����#�����p�O$�3R��,�0=����T�upR�Դ!�����O&g�yiP�x�B$�;�q��N�L3������#_Z���-a����$�Ԋ�Px�@\��` �H� �X���n��<��i� �(!Ҝ|��@��8�=�S$FFykD�$���KEI�7����-+��7���2��_�ZT�Q!��5�L�#�N�.��)�θ�!�����S�O�Z�"rQ�`p�8Q���-In"�
I��YҬ
]��t�eB�k�OZ�]�W�C�p��܂�m˝Bd{L���u%9��8Ǔ2B��H5��E�
��SM�K=�lx�dڋV���5GT<٨2��l(�g}BaLn.�J�	��80�$ՁH^���됯%^���ɯ$	N1���s�0��4g��X�G`���t�䓻�ē�Mki֑K�6��D��z}���5{�B�+_2\��a����L2�p��	�e�h�Do�(��DO"S�@��%l�|����!e��O�1Mo�\¦��(5!v�	A"Ц�~RF�7`9\�Y���	���c�4q �W���S�ȁ�g~�O��C��	e|�	f�}YK�;&����&!a�:yh��	+D�a�D�I:I�e�IOw�����I�y��h�Hp2�S��ɪ��};�옮�P 2�)L?s�c�\�{q(�'23��Qt*�7{ڀc�����N�P!��C�+�8L�h]����(�)�F�"a�:��t,Vu���1Ï#y[L�S��M�N��,��쎳9��%Թ&Uƈ���H�<���q�!|QX�3�N�����|0��38�@fF�)RK��H��'	�``r�Z1 �(1���`͚���B�,�%S��S�v�Tc�L�/>(��%�� x���eʐȂC���TmD���x�A� �J(u��'���O�BEƎ�X �$��r�E3!�X���0�%�M
xs��ڑE��m��o�>!p@ۂNў�tl���$�n�,�����$�.Y�h��<���ޑ~�|I2�"PH�2��Kƥ(���O�q�!ݝ@N���/_ *�>���Oil��1� ;�a~���!��!��;����U��;_s��A��0�F�5�>=8�[?%��Ϟ8����O.�X��"MT�A�hD�[N�p�C�'�*�hr旇A�:��raĹl��X�pe(Tk.H��v��2�E�=�P�5���+]�E��k�Q�2�[�|yaxboZ�kZ<@Ҧ�v ޟ]�6�Q>?�B����@>Z�YV+Z��yRJޡRm&i$ğ;��e0p��1��$Ȉ>tZ=�P@�
f�R�k$
Md�O2\4���]s���9����r�� �'(�Q�%���]�������a��lyע�']� �㵨���1�Jȗ��g�O�<�aᏠ����'ʨ2����I g�:��Ab�V� �Щe0mXQ	̖�p�ɕU=�� �SF؞hR�M�Z."�Q��׿kNɻG�;�ش����F�t�f�~��yBYw6��t��9bJ�`����7���+�'�h�؀��B!8e �.�*�Y��'ٸm
DB��b`��Z�f���;ҧ'*Q(���Q�H��e�e��N���bÂH�� �?-\���O� )3$�رd�(3͠s�j���D��f)QԊܓL���'�N�:��}2�?8�Z�!V  2sh+2oG���kp��+B�<y��4!�,`��TH����7���� �x�}0AK�}ў�)AB�15H�� ��u�\��˃�'�� 4ږ#�"�"��'׽�<+QL�cH<9��� _>}B�x�2}�l���E�%.�����d�v��E�U(U#�;��Q�R��c���=�!M<+L���'�b�[քD؞$����AH�iZ�iC�E�� ".yX�h�����_�V*��'Dh��.[~�P� � �
H�������w|�����"�Rap�"�ZuH#J/D�܊F N4.϶I�Ն��i���Õċ�n�dۢ�[Xf���/��^O��҆��6��	>����S>Y�x ��� M՞�y��I��hO�%�ďV��R�$�7#l��BbX�L�z�h��.]HQ�&M0YI"�#҃Zd�<ɂ%D�k�0�'ʰ#}���rb昪� �r&>��CG&]��D){\%a��T2`@�5 �-qh�`�q%1��$�'탕{���m=Q���������@ݽn��j�'˴@�$��O�y�
�7 ��2���K��AȔa_71��T���΃��Ƀ?meZU��� Y�u���bMV�����-\U�T0� NIa~B��&�	+R�ɼ4�6�1�&��Y�����C������A"lY��05�pɽ6�4�I�h�OE0u�4gX-~����8v����$�Mw����MQ0o7���Pg�~�s�Y&K�ɠA�Y+co"�S�+�?e�� $Ҕ��O?���|Ν�����,�R��1��-<��Č/��q9�"�Xd�Q�#%��� C�!�, �%ʀ�A�v%h����}9��чnp��$�E�i�e�fm���R��-*�epA��4cCg���fA�L|Γ)n٪©�EBy��G��Yeq�3b�a*�m"�O@q��g-d�`�r�|r�`���+?F���R�Ȇ�M����n�?9�lN�3�^�{�	_\������_�r":}�
�֙��G�OF|�v`�*u�d���ʲ��4���{�(j `�8�8�1���p>��D�*޽�$iT�%��񃦚�'�@=	�GC�t�2M
��I"b��?�� ���Hs��!�n'N��4�b"Oj�YD�� �`2�
�R �!�'vD�H���$7��P.� Hz�yd�����Â�V'Ҝ��[?��\�ȓ$�p�F)�2W�tm���ָ�v�4j��)[�ֵ�~�S!̗a���I0h@\7���y�@��ƚ64�8�F��q�S�'j��D�䌛�Tͮ@+���h���"bJ����Q��J5q�T����,�0>��3Ŏ��F���f��L ,e�`#�kV�p�Np��ƙ�?a�p�W�.�� �O�t}[�dY�@�A��5=t��Rߓ(Dq�3��>����� :���0H�I��f����j�ቢv����*�,f20���j�O��X!`��.���c�@G�օ���;8�%���ɀx*��@a�Լ5���g�M	#� t��b��N�� ~�ؐ �^>�Gx%U������o��Xs GWF	j��.�Ic�O�a@T�U�n �3�ϳ?�@9SGH�R�\X�@8B��(ӓH�s8�P����3A"yҢ�V�Dn��d��OL�	c��&��8�H�C��On�XT��9���&8���t�M��|CH3]!a|��C��l���jJ:f�{5��,&�؉��E� �G�`�!g�����#-�^H��yB��$�>;V�ٟ?����S@0X��MC�b$�0�>�wt�n��`	�Q�7��S}�y��#��LhuO���%��7U
�0Ђ��oe,��׭���ft[�-� (@��Ų'������k<���I/%��IF���.���o�$$��g�=@�]�Df�6&C�	�s����Ce��XX�MJF�E�0|�,���Q8�ЬKv�^�O���5�ѕ�jQ�Ю�0V:l0
�'� u�W�߈r���GL���|�a����� qG�<��'�gy2��[x�{����ju!jq��y��J�b��y0M3:��P�\�h���	��O�\#�#lO��A!�ԱX�z��Ƭ�<���'$�)��gξ!����i-ҽ:P���
�L��b�.*�����'���P�b�{���җ��,/�ő�{B(֖��T�GDċ��>]IGh�/Ip:��%Dq|��w�-D���$A� D�1r�K�8�pH���N�Q@ Z��l���DɩIG�M�r�H�i@:03�P��!������j]:�Q:ǧ�6b��
)!�����'3�X���޳f���뀈Þc���b�'�P�aG%G%3�Se�!	]М��'��A�A�j�5�Tm�rؖI#�'w� ��s`�Sd��#cj�'l�@�0�����A��0E#
�'�(FY%G��=+2�
�|���Q
�'�`�I���}M`�J�M�z�1)&D�� b`��ȉ(p�V����ߎ�h42�"O �����n�qo�H��y`@"O�DB�fǧ�T�)�.WA�Xis"O ���U��Jݓ��
~DI�"O^��:��лC�08���"ONb���10�r��5n���ab"O��y��!g�nd����z�
q"O<�)��X��L�W�G"r����"OT��g>#1&�{W�Fd�1�"O�I��nE�i�������=�A`�"O���@�W����3\���Qs"O��Bc�1n��0��
x�2�"Op�d�Y'/�p��N�*>�����"Od+��c#ߡCϨ�q�j]!�](4�`��pF��2� =���W]!��'Q�ȣkC-{��H�"D�!��M�,
|| ��O>�e���7�!�d��-�d�$HԛB!b�צX��!���^CJ��u+U4
�-�t�.Q�!�P7JD������a�ٌ^�!�d�r�I1�ح&���r�� 0)�!�$S�6ư��P�
(`��ip!�ޡ!�ټE~�!���	~ö��EG�`]!�䙺HwB�;%�M��ơ҈&k'!�dтV�b<h'$6y���� k!��ޯ��Yb��%s�M�K\�	�!��
.C�B�k�(��01B2�D9!��X�&-��!�������,�=?.!�D�>>��xᤈ$~����+P�t
!��>�k��X�S$ԂT̗�!�$	�"��\y`��s0J-���8$!���A�pH+1·$)�d	Q�X �!�M�0,���EnA�5a��MV�!�$��F$�I@Jj��CVfLz�!�Ā7�^E8F�|i�1��Le!�$R�#t��C�"����ac���q�!��JqZ����:�%�M#�!�DN��J��s��+s�f�s�,$~p!�䃂8���0r�q��5iJ�`f!��}���s3k9D0��8ǊT�!���F����vK)>�rt��&�!�D��<��<a� O��0	�LBT�!��2I�yg�<5��yh d�.|�!�E�JO�Uh��� i�V�[�!�D�n�"pCp�6qdV��q�b�!�
8� ��.�C���'(d�!�DR>Mcp��dk@�[:2$��g*�!򤅘Q�dMHC�z��0�+Q=:{��������$͙�Fr�Y��	���A0-2���8u�1H�V�&�P��u�!S֭ـ8M���ʀ`�@���QP����v$�􂇸{�����\��D�R6�A��,�(��ȓ>�@R8 |%�T��Q�$q��cg�M�4��� ;�)� CR���Ɇ�锡`�H�"�4W�[|X��"J�Z`A�0+%�R�i[+����ȓYi� �	@��ԎL�<�,��ȓ^Ԑ횇�͠�5��@G7Ype���ԝ�VjR��qk�!E�"nЅ�U����,R:x�2�ô�Ɔ"Q�M��4��-�U!�$.EV��O(����pI�F�Ͼ�(A�(I-���ȓ��Pa&)�$Y�!䄊*e�FH��S�? �E�*���i��էP���{�"O�r�b^�I���s���=T�4�;�"O���CS�����e��}�n�q�"O@�7؆���j�P�jhAz4O�e�1�L-Ƹ�������A��zy���V>P::!"Od;�V�+�6%�&-S*A����^������5N�T ��ɓ85B����� �f���E
���2 0@rƨk�zM*4�1L-��H�$���'��9�"���=��m� 7H�0��D��h�EA���O�4�Z�n7b���#"ƓyֈD��'( ��MM�8�X��,]Pn�xشbж�I�ǖ�?g�ӧ����dۆV�����2��YQ���y"$��Y�,�Z��A5a��s����d�#U�5[���
��<1VnG9�����A,�
�r�vX�xE�U<j���Ṅ29����E^jtEԇ�!Z�񄔚b�<��.o��c�*L�,���l!5
L2kv���	3t��Q����A���rS�L�V�!�$�)��xP/S5D��R�O�wɛF�W �U����@��s� ��P$�?�>��HɀG�,8D"O⍚7�T��͊�g^�V�t��W���l�&;�����'�f��᫁8cS@(��L��!7�H�	�Adp���V�u8�1Q��]�A�>-H� %:L`PQ3�>$���a!�$������ɝ,+�,����f�Yb�x�ɏl�q"�S�)��:��ɘ��A�tT,__^��DE�3�ɫPi�(����^���[����R Iy7�d�+����{�����(�蔊��Ȉu�~ŠQ�"M$����1C �G�B8���I<jZ���$E�X��R Q�!�$�dr<��@R�B��Ö́"⦩;!�GsyB�?1���}&�,�$h�!1mL4�T*�vz��V"9�`:D� �R�3��X4��� ���ZȄ�h��9V\�M��ɠ�H��� �
	8��A�Mƒ��$T�\�@@J�`�`2�
_J�
3$�	G�i�̈́H�q�' I��	T�S�O<�Rv�	Ad̬�PP�=�
��I��q���.w�%�u�G�O��{�C����&�
7Rj�qN<4�k����p��1j��F�()\�z@(��-�LQ�꟢d�剡*T���E��I?�.�N�[���왁BW�r4�9�#��� y��>�O�Qp@�Q�f�hA�ߏl5�[���� �D �.�W�O6m95Dxɧ�[@��I�
��t��)��q�p�c��ҷx4�r7�'�p�@�ě$m�ld�.0�-�"и�aFؘQRF��QK° ��9��(l��)U���&�	oR� s,�hⓅy������V�V3c�FZ �OT#C��X"��A�IU)�10nx��!ł��M�� �#z��H�<�4���
�5��y���A�  b2���'f� C~���q�B�6%�(O�	CR'����i�4d��<�kH~���<Ĉxp�\ g*�l5��Bm����ʂ��-H��/�O<H�b�P,C,����H%iN��K�&+��"AdB�9M�L�FĞ� �<@���.I8��	�oF��wZ�Ċv	XL�L�����wxQ�0_�����֗����W%��R_,Mx	�*cvUA��Z�z_tm)Ӈa����'�N��ҋ�(-��O�~]�W�_	2�aфG�R݆����|/Ќ$��+pP]K�fK��u��q� �@�E�C�. �d��9� �O�%��'��$>c��Xrc�6ˠ4(�A�\�9���<�F�P�
8�K�g՘#��0�-��Ij��g�I�`�u���y��`��P |���AQMV_��T�5�.J�@���j��r�h��GP]y\���O�3���4���O�D�Ҡ���p��~
��#�� %Ǻ9Y���ob���	{���Գ,�)IP�Q�dQ��F<"�B)۱Xr�X�)kqO.�N|rD���Ua0��+!�*���:O<�S%�=@����D��.n��lZ�%�,�y���8A2�OB�6��C�8R9���s�8<9/�w�0�'��yhRD޼"�Q2���E�>����1H����&s�ԉs�O4D����˜�N�t$�m�s�P���>��u���#��L��~R	O (���C�D�t&��q�g��y�)U1\&�'\�m��u�7��?ё���*}�]�&�<lO"��B��0.;&����but ��'�x9j��*W*�lZ�z�1#��;h�6��P �m|�B䉈}X6	1� )��ƯڔpBV�P�B����x"�S�Z�l35b����qb��C�)� N	q�V'.�~�QqJ�7{�.5VȔ�"ba�"�'��s��c&a��<��E(ϒ�G�\ ���$D�x��.��$�ӏ�7j"�ٶ��p��dI���q#.<O��z�EM�$+4hg������'j8���~�8��Hҵ`���L�G[��O���R�1&�&�2W�F�V�ЈO����d�#�(�"��Dc^0n���80�ذ
���� ����@c�.��
ۓn�p�v���*"���q	|�i�6O�A��eȔ�x	<}J|�@�$m��z���3��݈�Qg4�R��nB!�� �@p�`���?`����[5��*|����-a�` �e�N�~�'�f� ���GE�	?k����2ֈ���ٌnKV��:���	�Jv��)S�+Լ��1�ȜU��IA�>y���O��:�m�Ê�
��� ��AE��:Y��
��3Q"q�(p��aǬ(�|�I�J�O��r��ObQFkN1Pxh�ӓ�xA�e��K���@DHŠ�`a̓[C䌂ꋏG�Pҧ����~��E���\RV����a1�� �L `�L�0"Oj��+�l��)N�\�M�%�>yӏ��3 �t�p�ί_Nf���B#}Q?Ys�MT�W=dl(�E	8������"D� �f�/�����%A:�,B���zd�؂���J�Zҧ���ǺY��$9���P�uP�.
<�y�B� >��`��n��_>�p����~bFt���aǓf��K��=~Ozh3� ��	��t�R�;�O�����c��������Q���YE��'��EQ!m�<�3o�R�P8�m��X��I1P�/<�ri;�'�21����T�'��P�x����3)�
�J! W[>'�a~�m��H�@�+w��O��\X����H���0�"J�C��E���n\<��I�|�$��q��.45.!�"���w��=9����
�rB�+�I��H��F���to�W� ��F^D8�(3����y��
+��h8r�^2E�
��ף��?�Bʊ�&=�c�y5>Pq!K
�h�����Z7��!��p��M ��%D���vB��}�,ъ� �6d@��DF�:n+�P�G�R,K�X#�D�@a:�'�O����ݳ6m��X�;x~l�U�'|fѕ� (?�v\R!$ěh,�D����U�
�q>*�(�b�7&�S�aKH��Wȇ�R:(��J�hG{����%�QL������ӆ/��	�_&lP����b+^��h���!����^(��<sD\����6h��l*��s��D5z��AӶ͑���>-�#a���RR��n>�S"�Z�<q�g�V�X���W;]�XHkСtz�[U�U,a�v��5Hŵ�O����dMjzH���G!V" a O-�O� ��'i���8�XL "a���x���12 i�	E��p>����-hj���0�2U.�:Q�W�'ZВ�f�ϟ48s�ҮT�ӅJ�F9Ж��A7�I�gΎ�HvB�	���04
�uj�� ^5��{��A
�}E�d��<f��m�F�p�j� 7��
�y2 ?�0�����?e��!� �I��a�Sk
���>�p�d�`�W�NBt@��i�b�∇�q��l�����UaA�U��	g̎��>5ـk�a{r$R�>8$��'Ĥ}r�r��W��p=q��Y�HD�զא�M�VCD��	��s'F0��
f�<I -B��f��
f�Yx��N�2�"��2�F�Fr}����<"����J1sa���_r�!�$D=EY$�"���(�ҳ���V�+T��-G��'ft@F�,O$,��
.rb Iu�3'���#"O`���mZ�A���VlW�v��	�3�)޲U{�/�n�|��ɗG�|c�KY�,L8�XӅ[/l���dM5�\�v�$[7��U8-ƬXͦ�z�j��5wjB�	�[� ���ZNZ=�R��w�*�@9�@�@�Z E�W�O"T�si��{�������@��% �'�\�.4:��)�b��hP�5��j��^�xP�s�>a��>qB�}�H��CbO�x���E�m�<q�Ԁv�lD���7;�2�)C��x���.��}���)L�d�� �\�,�BL)���W�NC�IE7)�vk�i�*��㇨O~>C�ID��������T���i��G.(kC�)� ��JS�W)�PQK�Y�"O\yEC 2�<����@�[B"OZě�f��OT(NO�;��l(�"O�R����v�8�㵣��D�B��"O�x�@� M�B*����bD@��"O�� .�A	�!��{���!�*OlТ"�\<w��}Z���h�����'0�%�D�	G�D�04cBd! T2�'�DYp��
/F�d�+PȢ�)�'}p�;�o�6`#�|Cm�]���P�'������L�=i2�""�6�F9	�'�ɪ�"�YɄ�p,s�z��'|-X�
://�ѱ��Ĝ>cpez�'����I�5�����I��*S�4��'��1"A�,T
���1�G%]j�8�'X�)e�1����𭅇^_֝q�'hR�����<�`!��W�DM��'e����Cp�\�{�R�LU4��';t�j䫅�!�`�t�����'���9 e�K����ƛU8�'?�����شW�~p�UI!w�d;�'z8e��c��|��e��/;^t���'����e[�.H�e�SF�:ި	��'kJ��Q B�z��񭒄 ��,�'̒�4b�D�t����z��	�'K`m��Ϟ�V%��hG6"�<�'��q��� \�n���l�S����'�
��M&>��%���]�Ț
�'f#�ԧ&i8��"V�p����	�')<|+�#��b�@AL<$r"���7BB�*B��zO���F�9q[�X�ȓ,{��+��_�is��F�-m� ��bYJ���"Y7@Pj@ lG���ȓh��)	ʃo�ݓ��ttx}���̱�q�ͅE�IK�����ȓ]� �r��-~�d�w�Θ1V:���m�D�+Ui��.L���f�C�R��ȓk����eT�/ޖ�k� �4�:��ȓ!(ȂD��O�N�A�_#A�*���_���$�O�֬	�HR�(M��+:���'�0*���;eń����aN��B�7+7"���(L�?"n%�@J���ا�O��2�]7�v̛���c����'逼A�C�,-&ɧ��L���(u�)��
��r9�<)��>;����%�Pe9G'���X�((Ů���z\�S��-l�5 �R툜�O,܄ᓴxޢX#�"H#�0tzO�+\�DL���u��W�^��}rN|�K�)Hm&\�A)Y	t�j]T�A�	�t�hY	D�R��M0���M�K(�9[@��H�,;�f�.
�`�� ��@b F��6�tX���R
��W�G�R8ap��0�����p$xШ�œ6H�	 	{>�9�FM�^�����M�){��\���H#h� ���ݖ���M��<E�D�J��:U��
�$̞�)��
5�pq�좄B��OFT��Ӊ)3�HP��L6jR0�A�1j�Ƙ�"#τU��ʓ.Ū}�'G�ά�D���țg���7'ytΌZy2O�!~{ܘ S��4_?�1��@��%��y<0��#ƘO���OzdPG#&�)�SU(�i��m�r vă��Igw��o"����G'L'����T�:j�X)�^�!�d�<�PL�"A-�hKf�P��!���N�>����Z��0U'ݿ4l!�dޓu	VyfD+�4 pƟ�%h!��޺!����n C���P:R!���@���IaO�M0�����+8R!�D�653�M`�%�$~-p�`��~;!�$řu����o�� - p{�N+!�B�=C���n�|�������#"+!�� �`
)NM��M��H�%�Na�"Op9���U��}��[$`x��6"O.�3eAؗ>K�%Ju���zG�� "O��	؞����e�4n;�q"O$���Y
U��r�� ,��Yh�"O
�{��H���Q�M��V�"OH�r�/ '$��ɴi�6Y@�v"O�<锠� sPb=���o����"ON�c��$Sx�-�A"Q9���qa"O����Ċ�4��(Q O�y?���"Oz� %e�";��Ѳ�78 Q�"O�L�oa�̀i=�L#6b$\�!���0�6���H�(�y �]M�!�d��u��;$/A!F PD�<+�!�d��~�+��� 	����Dw@!�X�;Z墳��IPu��Ǚ�%!�D��Bܠ� �*�n��sl�A!�D Ft��kݐkB�A�&˂��!�d\�4\X2l�.`��3C�<s�!��+f��u��#�~�(��D�!�d^=Ƽ3f���B���#�^�/�!�dα��+���sâuq�I+�!�$��`z,����[�^��=Y!��)�!�����2+0�Ь��^�7S!�ďL͢iR����܁NI!�$�I��m,b���Ҩ�=	=!�Đ�k`P� �o�X�Ah�#M!�D�9(�����\�Xy��@X�M!��[�M "����\$4l�U�􅖒*1!�$G ��	��OȯBk��P�;$!�$ʷF\��*�K��#fqx��=!�d�Q�4c��.{Z�%afn�=$!��g�z�cq�E��|���͆�2!�D�4U�0yIUH=�H)�uc=r�!�d�0e�P���n�">�ҍ�hP;F�!��P�h�%F�G����eh\�Gq��$ʷW�茒����M�`O�6�y� N�?��$Ӈ�3D��!�ehO��yR��k<V4IRDǣ":�3u���y��B�,y+@�Ps
�P���!�g��VB�T���c�}!�d�1>�,���D�Y�� �Eˮ@!��Čt�I��	!�d���%�;!�䈐V���3IF�$|$��#Ε!�P�s�l��gY�*f9K ��7!�$�:���q�N�~��r�-�K�!�
K�MB�FR3q�N)�e,xd!��	cܸ�S`�2Z��(ru�οc!�DY.��x*c@�5!� �Y�,C0)K!��B<F%���"�ʙ�U���JE!�\�,��p��"9��4C���:y5!��ư�U��M_��D��a���Py 48"0hQ�LZ�~m`�T�yҨ�/u��I���OFx����yboD�?�F���H�&=�v�;PI��y"�E�I�l���"G:�LQ�����y2�H����Z5�?9���؅ �3�yb9
�8�)&DӬHL�a�C���y��ήW��M3� A�<��mM>�y�ўD�P�Ь45f<a1�]��y+0"���$�	�3mt9���8�y�'�n�!�9_+l耵�8�y$ڎ�xp:*
M� �ڤN��yb�PV?��kD� C�ڠ��	��y
� �q�&�8,T-qpl� R{����"O8q2�I�Z{�l��n��ɫ�"O`�hI��@�,�2艛w�"��"O��Rq��^
�t��D�Kk (`�"O�0�fd|(�)�I̢F���"On�Cщ�.���r�=fy�h�"O~H��h��b5$߄[e��i�"On�e ��I\�-��(	�,�F"O��r�%-RT�!��~D�q҄"O~�2�f_�?A����G҈Z�7"O.d�Ή'�\I�p�ϦN�A �"O�i����-��"�H��)LH��e"Ol-aw�P6_	�Yh�F *~Sr]��"O" �V�Z�p��T2 &9`�"On��삛t�����D�MuLMBq"O�`)𪅬]Q���/��L_�A "OT�X���Ze8�W�@�w�XX�"Oa!�gG�L�@9�� Y�(!�"O���*ʈr��C��L*�F��p"O�q������Ү����d"O�Y���n9jí�`Y�"O��J�C�*(��!�":ڎ��E"O`����R� ��p/ɐH�&��"O
��2��F¢�U��;�Ҕ�f"O�L*�
��g0��M�M���"O�����#c����c��b�5"O�� R	���&0����!����"O��:r�;p���1Q왉z�d�Q�"O���0�Ɠ.v��I�#��;U"O��3g�?�VA:"��.3����4"O\�UC��5-��cV�Z�ƨ�"O�S�✎U��P�مo�0��"OX)��'�86j0�"���9�d��"O���/])S���P�@��r$��"O�Hr�(�@����m�?KL�!"Ozq[6n���@Aw*��)и�!"OZV�Y�Z�� �B����"O:� ǋȡQR�Y ��X��"O��q��J�O0�@y�d���Y<�yR�v� �Td��{�Vy�5���y�F�3<��`ȎF������yB�u9���s��8�ir�g�0�y����?�M�͖4�ʩ 4G���y2"��YĒ�:�(O&)����T�ט�y�˥p��CB����~u�f`�9�y2��[��D��+ O��y��;�ybH��Ux&�S��n�x4���y�L���j�����0����(��yR'��Q�]ѣ�đ~yp1��gא�yb�Q"7��"鎤	�
Qx3����y���g��9�!"H .���Ac�y�"%>��q���1ɒpɡ�� �y2G�4;�%�dK݌(��k�:�y"@O=$<*ŋ%L�4�e,���yr�6	<��	���+0�8�#��;�yrMՈ,�u]/#��X-B9�y"%L�yv���Ch_�d٤͟�y��L7o8R`�!Cбe�z�4k���y,�N�|� ��>e�x�yC.�yr���c������g�I�C/\��yb�ǡN�rM�4'�R���5��(�y��N�����FFE��i�d���y�M@�
$	��d��Cv�E�T6�yR��(Xp��]*?h����+�y
� �˃*�&�e��(Q	Y��h "O�}�B��<{Ҫ�*�'	7�p�Z5"O"��o�1~���� HkʬC"O�]��ݝ\�"M{S�R�t]�� "Ot����j?xM�ʕ.3A|Q��"O��&j�"K��©[�K9�x��"O&EH��P?S��4H�B�&�^]�W"O,��m�5Pr"�
3AQ�\�F`!6"O�$�ƩsӠ��Ǡħ]f��	'"O|��T/3FƁ�C@�1&c���"O�a��ͧA	�ȶ&E����"Oj���H�(}�b��BRR�؂�"O����j6>z����Q.�v886"OĥE�9[����Z������"OB�!P�C�\�t̓����"�[g"O��
7�U�@⮨bP�L;l� +�"O9���ݳO����1�߄im,�u"O�����qڸr��
0l`�@�"O���`�ۚo^��J-ɛ �H���"O�|{��/����Vk��J���[V"O����僮�pA+�lh ��"O� ��菈GԸ��dʁ��F3�"O96�7RN�Z�	�E��|��"OFD�s�ιXݘ����H6�dP�"O�A�(��Jg|�JB��'늬{d"O5��	`����%���p`S�"O6ͺ�O73����l�}�B�X�"O$t��#�* �Q���!w���C"O&) �al@b G)u�P$z�"Ob��$,��N��Z�nS�\�D-t"Od�ć$!b��R�K4���"OL�����,M�"-
�h����"Op���Jߘ\7�k��ɴYZ@��"O@5Y�)�b�B [��*�j��"O��ʂ�ޞ[��pU�y�`:B"O�s�'�'��� �����@�"O<��t�\�0��\˕+L�
� �@�"Oj\*Wo��r��#@�?H�"O�5���`v>������`M���&"Oؘ��mǱS�$i�OD	Fn�v"O��ҮJ�2(5�.�)-"�Xe"O�ԑ��RA�JPx$��.��&"Ojar���q"C"��`0��b�"Ou�sF%���n�"5C��p"O��K���PzQ[Ƿ�N<x�
h�<y��.b�Z�y�,۶���S#�c�<R�O$R@DЀaM�ܰK���K�<��Ɔ�R��9:r�K�^�C�.�l�<��`��B>Y���M�6iTh�I�i�<䉖<@X�k�oPL�H�8��e�<�΅;_>&){筛�_x�`�K�d�<����E�ҐH�̈́89jUh6�
Y�<��S�&?�T@R.U����Cn�S�<	I��H��0! P�4�����e�<�-�0٣����ܳ���J�<�-�5>'0<���5xV���,m�<�B�]C���b-E�l�|ԓbC�<�D���ؚ�^V���HW�<1! �u$f����I&XB�#r��U�<���V$ @  �P   �	  >  �  R   �&  2/  t5  �;  B  TH  �N  �T  3[  ya  �g  �m  ?t  �z  ��   `� u�	����Zv)C�'ll\�0�Ez+�D:�Dl��F>O$���'h4�l��n�p�2���cZ��
J<�v'�l�6�H��́M ���n�SA��?�/��?��A�d=��pD͜�-��;`Z�"оI5HN/`z� �Pf��S�c.�#�uBի*����'4t� ᢇ�X�~�i����ε�fߗG�����-�OD����I�������$��۟p��ҟ�������S$Q�#�h�ч�$�!Ď����	� �Ly�4���O����D�D�Or�@�/�U��c �	�8=t�ca��O�ܣ"�<�������u�u�	�<���\#*�3aE��!��b2��.��p��yR�ϥX%��[��C� ��U(q�����>��~R��j��p�O(\�[�F@f
�V���܈T)���?Q���?���?����?i/�D�]�a��Ms6+��_�z9a�c\�oF�����%rٴb�6��>i��i5�f,�Mkr����?�#$՛*�򩂦I�kx��м-g���f��"�Mз%G%4V�8�C	X�t�(2HD�}�p6�IͦY�4�Z������'��	�n���04)��k�v/��ԛ��Z3�:�kRn�(A����� ����7$b�-�� �2z�\8�ʆ*+A\��O>����#%B�X��'�i���$G8џH�	ܟ\�|Z�
L2=V@��j��i���Ouy�)§n��)b���y�~(*P�I�dS-;���hOF�d�[��o�s����� ��5��#���{b��;�?�)O����O���5���1�E��8�^���OX���Q��xȦ��7<�n��*O��%�/M�t-u�9U#��D�H��<��G����k2�l]�	�5M�	韠-O�$����!p����"	Z9(T�'n2�'��O1�:�I">����nY�EL2Ijq�J5oJ��E{�O� 7m׹mҰ���C�G��Ԛ�H0ey�o�Z�zH�؊��O[^�5��W��13��%>2FUق"O$���dT�j���C
ҷ~�|A'"OΡ2hO��p��W�F�(����"O6$�sMJ�)�MjnRXDJI�R"O��s-S3��i�G+�0�aU"OD�z�gF�y� ��j+*��԰%�'���a���S��V�c��(Z��6��'���ȓ#�T�D�5Ȏ��ËE�E*�M�ȓ\�t��ħS�t��msUi�!����ȓ-�`�8�
�;;{z�BP䗂�P��ȓ>wEcfA	�8���B�������ȓDe������;��ԹY���'u�i��d��� �ۘJ݌}Q��(G`фȓ�H��Ž}���5�M�P]4|�ȓo|LJ�ǎq-��ɓ�d�r9�ȓ+Z�[vO�&@�`Ap���7���iRlЗM�t�
� 2JL�8Y�͇�7'#̘`�4��D۾#3��(�
��2����\��"R���Iϟ�ϧ]VY��H�UᲈB$�?��E,�|i��L�<y���p�d���0<���Q��}�7!ʹ����A`�A�䘚 z�����S�AR���%��$�Of-n�ϟ�Qb�V?9�� Y�|��YP)Qy��'��OQ>�I��B�X��$��e c� �N%��۟�D�MkӔ5Y����]f�qR��(#z�ؤ-Ҧ�$��:QH۳[�H��?��'[hJ�qV��L�Z�QLƷ��8��'���4/
z7�(i�_�b�\��'Hh��� J#��� %�nI��8�'�M��퇫|�M0�埂e���+�'�ZP #�!�(�xBĆ�[:�h�'%�z4l��Gjʩ5E�X��ײi��'�ޤ s�O���'��X�<
��[�=�<S�!V&Eؼ!�A)>0)b�K�/M�`2��+�f`�O������1"h�jcR�hؙTkF�j�s1f�6VB&I&A@i�jc>�5��Y��$�8� ��� Ȃ"����� �l� 6͒ByB-��?q�����?��c�`�`�V>xq�m81J�-\�)��u�O��Q�>Z@Bx�*ܘ v���'_��gӊ�oZ]�i>��SSyᛑ_�N�x�$� �X��f���x{��dӌ���H�a�a3�X"D-��ҥ(�IZja)sO�R��U"����|�$Y���ގ\�!�DU$r�`��o���cא^�Bv�'�LB�	�*.��%�e>޽R"I,~x!��C1DZ}bR �:~�"ꛢh�'ŀ74��	�7�o�j~ҥ�e�6�����_ ��)tD�?�.Od���O`�d��wJ�"�����J��z�� xC��t����l��~�X��'�� �Db3T;�aJ��3�y"�ΠZ{� a4�A^	VHH��0<��I��`@ش�?��Xl#���#�I�bm�y 0�����?���?���䧥�'i\�s�#�O�<�8%٢w��Q���q���K�
H� \F�fj�S��?�-O�͡��Ӧ�F��i��$Ƃ��(Q�� ��	OP��ɲwa�"<E�Tċ�"����˳(�͈�����W�QE�"|*��H�B���}�ڐYr���s���
�ڭ�I���S�O��"!��	�Z$0��'+$�b�'K|݋���5Ш��2� ,0|���A�OCn���i�1DȰ��Gʤ|�dā�i6�'S"����O9��' "T��04�ȥ@y��0��֊ysL��3Ʉ�����OR��p��Yg�F"��+=�,�rn��~��'N�3������*�6m6Z�"@�e��?"�D�ੁ ,4�%�"�ݮl��m�8�ć0dY���*�<a�h�h�eEO$`�.䃰�նd�T}��D#��?�u� �P	���ת� ��(�3�?Y�� R�	ey�X>��	zyB� 0F&�A���rl�R&�P�N!d��r�����O���<�+�F�D�(R�S�Ζ^X����?%�LRk<U����ɬb�z���L"p ��i�͖>�ٸ'�M��K�ǔ#���	x)�.ݚs'�@Ȣ�ښ&��xC��O��m���'��	�yE��:�`(\~��:v̆�R(��D6���O*��(c�$�%�ܟ%[Q�`�D<?� ��㢱<Q�l��'�ɿ$@{ش�?a�'�&�iB��3ߪxȐJ�7�0pHÓ!9DDxB*�B4��G,���}�r���0<AR	e�'��i�-ś|N���*����l-�4��7��F2�2HZ�o�e����d�t��c��� �RkjXc�K�2P��Ɋ�?��K� pBVdٱ��iҤ9���l�ɛr*v۴������O��1��RWx|�愗5%��=�W��O���E#_ ��O���%�S<Ф��+�l��FX�yPv��'��@c&�*9�rTQ��K�d�>��C�M� �(��a"��8p��X�g%?u��˟�ٴ��:�If>�	���?s�!(f�A�r��(�$<O~���O.�x���i�E75X�Mbr-�52p�E{"�'�����df>�؆L�@"MQ���?.5(��6�̦���Ay�K�3�t�'��'��F���!�H7ʨ+��12dH�O����J^TQ� $c�'7�����#j&fH�g��r������+�P��5�h�����h�DZ1�1Of��D.�9� ����$B�f�#�'R6m�O�i�D(�O�b>��?�7�I?WR����ʆ@�@������hO|�=q���&]���/L���Bv��-oX6<��?9�U�|�'��O��I y��G�	FC���]�>��U�u.P#�M���?)���D&�ɒ:E����Ƹ	�(@#Wii�e��$�^;���I+mNL��e��'C�1%���f6���J�nԼ᪇"Ii��l�˓ݨ�"C�� Iؽˀ��$z��3L����Ƀ�M����$�O.��c6�]6 V�����0n5x�iu&�ןF{2�'���V�x���1�P�pIH�2ԠN.\����ڪO@ʓT������i�5O���`��]7*)6|H'�'@����П@aDT$\�!KE�ƙ;v��JQ(��9�G��KJ|P�n��0<� /C�:R�Y�FϢ@:�L�T�i��)��.������RE�l��ej�uȤ��	<�M����?����]aW��F ��E�?a���?��?�J~Ҍy��;iK�㱇�/ݞ$*o���'�ў�+�?BG�	�hlpv�ƒn�X�/���$�<��D
?|�F���4�6m�O4��E��3���
T��!Z!	�O��D�ZCP<A��T���,��f�O��?�+�"\"u����&�R��"u�3�S~�I׼P��rA9Ŵ(g;ҧ"d�#�Qv��IĻ|u��'8��`�� ���C`Ӿ�d#�'H���c�#�R�����A+9�ԩ$���I៰D{�O3�<��AA�y�Z�t�$�d��D�OX l��ML>i����5>�a��L�yp��`�9�B)X�3��O��Q/��H��[���`�腝E[PB䉦ev� �
ή���;�.#@��B�7p�`�����N)���s,3Y�B�I�t:�Q`DGT�@Ӥ�kn�]$B�	�Wy.52W�$]���sI�4�C�I�w>]��>u��d��״˓MC)��*`���iW.�:s$���Q�0B��C�)� �8 f�܁$�~(���-<�E�B"O��7-@�L��Cg���!8� &"O���A�zx4P��#W0֋h�<�� Mz��Q�W���kQF�gx� �������@��+� J@	V��zk2D��pU��o�ƕ�e�xS�5�P�#T�`C@E]�P����>���9�"O��)�EߥVD&9X�ŉf#x4H�"O
��䉊hcry�g�	'����"Oh$�����=�,��*�|ݼ�!�I�e�ƣ~ʃ�ߟ|���b�-,A5JQ{���I�<����:%&^ՐrC�+� )��BA�<q7�
�'x�شř�1��̚��s�<a�� 5]���*	
@��r��p�<Y�FWd�|#P�аg3��A�.�W�<q H�{[*�١c1%:$b$��|CXH#<E��B�y�*lqU��w�������.�!���6Ő��Ua�*M��9�炘/f!�	�X �Y#�mƭ%'@��id!��3Eƨ� �Ƥ��2�䝈ib!�D�[f��3F���:y!u���j1!�D�R�2�,��q�(mpQ��j��	[�8��$��1H��L`�x!Cf%Z^�!�d	4�
���w{�A3���t!�$Y՛⋞	I������q!��ؗ7W��a�"��]b���m��N�!�D�.u��L�bꚭkTI�t+�$��}��R��~�C:�d$S^,qv �%�S��y�-O ~����b$�
:!|�2o�0�y�Η�I��q��	5�J�Z!M��y�� �Bhx�b�+/��`�O�#�y� �?9�z�aŎ�>$|���庐��'��`Q��'ڬ��B�C�S������G�F�Q?%�$*���h� �?F9*�b'5D�0� ��K�	!�+&t� BD2D��3�Q~��a��O�8��jT"2D��K�.�+�6$�l�&~ฐ`�=D���gl��R��x�֮7�@�M-D��#��\��mr��D7`���e)�O��12�)�'P����b*�/o�H$��
Na5�	�'����􂒵<u@�,T��d	��y∖�0d-R*_�_6�U��	���y�[�h���]�R��tS���=�y2	��Q2	��Պ �`��X �y���`�i�%��J��I[E+ˤ��I�9;�|2k]�8�@�9I0+%Dd3e��9�y���D���2H��� ���>�yr���Jy��`	���V�p�@S��y�@]�C^1+�MU�|�p�Q����y��yj�q��f��w�؍����,��>Y1+ S?��	L�Y0
��@�/ՒMl�!��'����@¹�Z�W.��L��	z�'�z�ڳGßK�X�	��Fb���
�'XI�� W9p6�0�c��ge<=#	�'�d(��FB:��@[�
�'�d���A�-r��Ha�g�=��i��D��f�Q?��Gg����u)� J.Bt��Rt�(D�L�1	�,/�x�2Eʉ�Yu�Xb"D�T��תX3�$�
�"�Z\2�4D����FЎ@A4���NY�CU�P'�6D�t{��R|�.uã��H��U��9D�`�򢔗Z��[aX�]<�l����O��R�)�Rn�8B�^�t������ "�'���׮�wV,ts�n͠d������� NР��!P�,�16Ɵ�w� �0"Ol�I� w/ء�P��Z���2�"O<ɫԋ&y�ƁHӣM�DSW"Ov����C+Ήc�ސmw6�7Y����a:�O2��.��p���+�!~S��*�"O�!���>���$Ĝ:8()��"O��'���<���C�\��@��"O��ːm�a%�5��֮qM`���"O���6�3s���d�&Gİ�$�'�:M(�'|Lۂ�ݥ@:n�
����M�c"O��PTbJ40t��a)�:����"O^��U!@ZL��F�:�,3�"O�9�Ŕ,mS���$؈<
�<:�"O��Ѩ �S�έ��DU�C�� �w"O�����Ɖ��C!�� ���I���~"SٴF����p�]t�t5:���c�<�P���e�xK���>��cmF�<�r&�v����A�0�2X��.w�<�Vg_UL:Y3E(����h��s�<i[�Y|L��,E	Az������m�<� ��,="r� ��Q�w�p��Q��0)��8�S�O�V<��Eޤ#�����A� H��a"O��* IY�ĄF��4��\"O)q��X� P�$�/*ي��2"O�Q#ë�I_@	r�o
�$����"O`)�d��r�� ad���؇"O���D�\�v�Ce*��^c�D�V� f�*�O�9��S�BШ��c(�`c"O21��y����#@K8��ep�"Ov���@:<�a1�]3�X�P"O(� ��)�Dkt�=��q��"O&�����P�	��%K��u���'@8�P�'��8�d�.+8L�BeVX0�T9�'�J�9n̠v���-y����	�'���ZB�4��
�ˎ�k�=1
�'Ҥ&�>[E �IM4v\��'��v-&^J�%�w�����)��'5L4"�.bZH�Zl�R�@Ȉ�Ĝ�lrQ?]B���B �GQ��$��$6D���5DC0Ie��U>��b)D� R����G�lE��L���(�&D�X�#��� =��
��I�ʗi%D��bւo��ٳ!�Tl0��E>D�\�%l�Qo
�x�V�1n0�p���OȤ��)�M٪yKS���a��W�@eXX2�'��er!��~������:؂�'~� �g�&5�(�Lތ�r�P�'��(�5gĜ@��=�t z
�q�'C���F� ���4�En[�@�'̕���R-k,�T�0��"xǾ-A*ORL��'	���V�C9��(��K�h`ʀ9	�'g0�� P�9*����cq�ɐ�'��Q��H�T�P�'��_:Z�'����Q�O\�@��i	1M{�	��'#��TmP�wJ�p��֑G��i��8Z���u=�����PA`��(L�o4pC��,D`��7	�����Βt�B䉗)"N�0#��n�6ʢ˺=�B�ɯh�A�ӏ��X���R�)
)
B䉇����(�����s�
-�C�ər��c(��_Ɣ"	T�Ab��=Q�I�M�O|�\�f�[�~	��抱yբ}H	�'Rdd�w �[��j��]t<�M��'GfD�tC��1��L	�N�T�\�s��� B@���ҦK�~��gFO�(�I5"O��I�'ֶI� Sq啍0غ8"O�C$"��f�!�ڳ0"4�S��'�|�����~��T�0���2Kb-BDɃ�aV�ȓ�*UD��T�d8�UA/��M��-"�`��|��l��çx��ȓx��Aaӆ���]xt˕,�$l������BB9X�X�	� ��,�\9aS�L/|�C���YP&��'B��
�	#Z`ʆ�ߠrT�� F(&��-���� �D�߾Z$ 	�J�/�6\�ȓ���!cM�"�x�d�M�.(��W5D��?�� h3�K����ȓ'�d�f�D\%��KF���Y̐���I&3n�	3 �*��c�-{�8���y�jB�ɱv7�#B��($7,qUg� O8B�ɼݺU17&���� �F̩@@*B�Ƀ��b�Y��5�޾+4C�G�XT�@'D�O�F�1����fB��=OZU� Aϼ$��qԉ׹M�V�=�� Lz�Ow~��u��	;�l+���|�	@�'��视OiqC���	2$\��'��D���߮U�h�s�=P"O H�&9+��`��	n�R��"O�`tj��^� Ts�Bл��a"OĽx ��5����KIq�����'m0�����M�0�	B�5�@�0M����vx\���DM�� Q�є �ȓaw6l+ӂՍb���%Ι�QM��ȓb8=x�j-^� "� W��Y��2��`Xb��j˲i�R'�&Y��Ɠ�6���M �_�8���_9Z����#�����'6 q�'���z������>��"ʲ�p�H�Ck\�3l�4#��i�'�FQӡ�նJ��|�r��
���s�'��hi�l��J�6(��Ł��d@�'��PY�l�E���1�Z���r�'� )��^�$`�7ό%	=.��
�'x<J�ëHε�'Ó ��9���
,�O�'�$D0�'�%7��s�,�m�$L������m�yB���e��fLͅ���Eu@�?z�gl�8���ȓ\Z���&��/����R�F�J�V��ȓ�
�����8`-�h��.W�B��M�ȓ:�v�2! L�"��[�5,�MP��(��h���� '���aH�&�>��qe���!�$�~����%I�~�d���c�2_u!�;H��A�$&�u�vxX� ߹\l!�R9|�����I�RUXp�_fP!�ɮ��0�iT
h�´2aد1!���v�0����*��U����v+B�X��p?���ـmWL�jCO�XV��!	�R�<�����rg����6kb������!�NpyOF%ld�UReJ\�~�!�D�n�R�H�'ڱ@0K5I �K�!�7 |J\��[-G�
���Kps�{�@O��W�4D��JΟB�E�da@
n��B�0%�X`v"H�po�p�A #3�^C�I4dL��	�2jl���J�X+�C�	G>�8�"�;Va�=' �2E��C�ɭ/��L
��M$���C���L#VB�I*�6��%�1��i� ��<⟜��%�S��3zy�iB'^�S��@P�L�8'	!��T4to��:t^A���F�b&!���' ���[E��rбF,�*C!�� �]8�5�D��G����Y�"O��0�.Y�BXxx�OK����"O\�+��[�،bvȁ�	d4�Q%Z�OT�}�Qk����ʞ�tGXB���#xf���/ṯ���L ȍ�`�,��ȓ&hh��bNzL���b�6�<��1�����;'J�xf	/��0��B����A.׾Q��h�L�[Ly��`NN�x��A�o9<��"�CH�)��7Xt���D)���RB����A2�/ԭ%�!�]4n� i	7> �X"FNǯ6!�d^)u|KY0'm������!�\h
�'�,�����<TA���C�f��	�'v`��兘{M��B��+�(,�ʓh�$1[j�'O�j� WM��\��5�ȓUoIs�k�#QҚ�� ��k4�x�ȓ8`6%;�c�*(�T���7�^u��ז�S`$Z�-~PU��`� �2�ȓE(��7��Q�H��: �>Մ�ۮ�P5��V �kI:_�b�'6�'�ɧ�$�	
�{F�I&�ŭ$ݚ��޵o�!�䗩_P� �H�_հ�;ť�%��O�6�8�Dү��'HPIu��>3Ĺµ!�#�� U�i��g�8��S`]��'@���'D�$Π#mN�3CA�drN��@�V���/GӦ���lB���I�<)2��znz�	�ȟk�\����Rm)0�ZT'&Y�YA��?������yr��.���O����O���!Y���ۄ�C;���mx�F��K�Ob�D�l���$t���*�?7����O��Aэڰ	U�� HN�2z���ڪM�Iҟ*�G������O����z�DB&A�	0��VY2P��	3%���	������O�p��O�扞RX��s��H��`	�Thv�v�KT�ã��	�[�,�Iğ�:t�9���?�'c/pp��ZY<����Ɛ�x����d���y��8�?���vK���O`�	E���s�¨�SX�Z�Z���՚�؝�剺8Ԍ��e��1 �O��X?\����l�ɾ|S�UY@gL$.dd)C�Kn^��ߴ)	� ��'N`�r��?A���?A�'Ӣ,�O���gDX�f�����b�'bɪ���iˆ4���'�	���)�>�e�<TxȠE��3m	+��yJX�!'��r7��@�q�π$�M����?+O.��O~˓���lH��I��D�
�����e� �w�i�X��	���)�O�˧�?I���*_&�"P@��d��  �[՛�Z����Wyr���U��2�N�'
jDC�	s�����3�yb��-w�4m�w��VR�Y��EM$��$;�Oh�a�O�6��PIC�z�6��f"O.!���8�������&A�X��"Ol$!E���,&vI��Bq�Ι�`"OЄ�@�x"�1�
��5��"O�y�4��H�l�v�F�&��$��"Oz��3손3gMrA��%�n9�"O���6��u�m1�`
-���@�"ON�`�H����73, d"O*��ei2�����S/M�b]�"O,򥃇D �l�r��r�����Ԯ15�@"dk��(���b�p4f���B#L�N���&Y�lTlի#�1@��;o;�82�˱N�~횢�wYb�N��#�i#�bV�^Ӯ����8�ٚ2�ޓ�\ �鑦x�};C̨Bp��I�@� \�&*`��0�`�.zH��/]�L}*�O���F�8WPV]�X)��	��{�<q��A���)�J�=��ԙ孟S�<��#v��؂3�Q�#�h�(��M�<!0*ə�tb��
*� 3�YJ�<�ƈ܇f�@��E��11�����|�<YA-�#k�L��&�peLU�Xp�ȓ���:I�X��Sw�N�(v�i��K�(�z�Ĝ+?|4*Ӫ�W����ȓ5�8���!�i5��q0�E�:�d��)|�I�ʋ�U!���G4�씆�4f�X�%�4�]�2���v��ȓk�\K����T4�L�0L�/�Hم�~�C`�4��s�H�!xI��S�? �X(F�ߘa��£R�~W��*�"O���@ P39fx�`\PV�Y�"O\aJ�b���>Y�2�Ӄw3�E��'�̪�`B�:��y�H������'ξ�����j��Ԧ
�wHY��'g�X:��G9Ihp����7jq(�@�'۲HFf4Kz6�)��ڤ
(�j�'�*p�FU/s�<�"(�#+Hle��'N��X�o�\|�"��</
���'�Lxi��U�w�~U����??({�'�,�L�8�x���u��-3�'�1z�$F;i H�HK3?�"(!�'�B�c��F�X|�(`���7���'�h��gЕ�&Mѣ�N� �'���B��d�s	A���
�'xi�!�Q����j�l�:f����'>���gn²&��m�LM�-��y	�'����-Ę<� �c )�9T{(��	�'�Z�ˠ�è]�.���f��Hjz��	�'��4"��K %<@S��ϚN���[�'nة �#G�8���H)H���'+j�Y� ֡_���R�o
�h����'�J|/L�\+&eE2*ZXq��	��y�#�*]NFq�1됣(����&���y��m1�d��A��JL��E�F,�yr����g�,
h<y6�χ�y��U��^��ࣈ� �$}#6���y"��e�Z��֮��,�jB	�2�y��c�L@!&�U�
 �)+RD� �y�!>�F��-����(q�I��yR�*><N��#Լ(t� 셏�y���i�Fd���)sP�{Èɀ�y��T�<c��D�ow@�3�H��y��т"[2�6��8KV(A#H
�y�"S�JL����Q ,��j��y"�
�<���9Tbu'έ�Q��y�FTA�����O�?l��]�1"ݼ�y�Fɺi�(�ƌ�jg���7�y�j̀}PĤ�"K�^uN�a�_��yb�J_c�d�T��	Y�l��ЁS$�yR�}�n����ݜXw���ׂ�ye̎e����s	�C�\�1�һ�y�Dܫ8%Ԑl�P/z�v&�y",��xT�����O�̄ v� +�y"�R#�l��e��Pmx١e�@��y@_��*�!�՟t��{����yB`W�L5d��ƇŪq,¨�pA��y�C7xX�i�fTi5�U8`�[�yb�C6]I�]�
�j����gI��yc�R7RhVaO�]�F�����y��ܚ�B�sk
�[�~��c�yZ���sm\z�.����.1�C�	j���� )�b��칱�͕
ݒC�ɽ}��zd�K(NQ����̑�&C�	&#r��'�C�'�2	
�@C�	�'X~ੵlE�wвu
$�7~8�B�I3tE.-��ϱ
L���C���B�!W�\�1I�?���S��	Wq�B�	5C���K0�1l��AF�U��nB�I�C첩!v�ׄ\��R���B�&��d��\59�j�#���.:�B䉒u `�'�S8ǘu�9�B�ɅW��{IL<h��B��X�B�*`�HZ�5f�"(j�͗|{�B�)� ���C�
��q� �΅�3"O�|��.��"��	A��H�p���'l�}{ J��Mg�\z��7����
�'P*��+��iؑnY�r!:�'�
uy��,�T ;d*�P@�
�'��*�J�[����bC؃L�Vu#	�'����P��2-�Ds"�I
sI�A��'���	p��!eЁ$Ob��Qq�'�2�3�8b�+�ONWa�@
�'u\�!�Nċ.�d9�r�J
�'��Z��]�R�# !�6�*5�	�'� AAP�_ X~��ƽ(>�Հ�'��1��ټV$dA��N�)�'�6�ȵ�Z�A��ȇ�!k�'�[����TM����B%�	�'�А�dA�S
@C�� �Թ�	�'q�Y{Wc_%�vXB�͑l���',�U*�f�'pl��� �`�5��'W0�9'B��1�aH�!��Qj~9�'^r�	��]�$���3�%ŧR��Й�'��(���e���;��جH{��H�'�ē��$T�U���;���
�'{�)���%�褈S`��/~�i�'>t31�^&��@#���'�vp�'r8%�Ҿa����ҋ�)p��`(�'��(b� .%<�����p�Μ
�'�A%�	� %ty����<w�p���'��XᥡŐ ���-M�|IX���'Ȃ��j0d��%�h�$Bqr��'O�y#�F��$��B��#���8�'�b!x���; �T3��{� }��'��9#��*߀�gD�p�
��'��"��9Vv�6,ˊa�>1i�'�,� B�W�("��B�D0S&�C�'��1��&x���S�#Jzi��'"
p�[�*�@�B��-Hxf4��'F��!扂�T �|22��);4db�'�Vu�Cʀ�DrY@��2U�����'���d)�H�<%y��NL���'?�X����;>d P��Jd
���'�`���c@�*��ղ"�G�D��h��' �
#��#A���aD�L#��Z	�'ߎ��g
r�p����>�x�	�'��-�Uj^F��	�)^aG� r�'q>�2teط���3[�}��'4���ʋO.��G�ښN�x((�'�Z��]�#�%�"��*;�u"�'t�h�B��6;(�j��/&����'���,"c��q'@�T�̼8�'	��W�ȗtHH�HG�Z�Jj�e�	�'���;��X�$^Ĝ)��E�1����'����VlD����GEʀ/�|�B�'�XW��Gh��*%��;�\���'^6�@H�����;F�d��'v��Z�� .������P�i�'��Ҕ^�4���R/��A�zԁ�'�&��g�.�c��ԠNf�1�';ɢ�k���z�	�aO�5F���'�`kB���y�v�ǘ�D\�'��6��4��AZ���m�:a)�'�~d�r���Z���w-�l�H���'�����Kv�p�o�8�����'��A��\�i���h���Zڑk�'��1	fǇ4W�txj�aBUKRй	��� ��A�9T� ��JG<Au��0"O2��FϘ;}tj��R�u�h�J�"O�9#�-,f:4��%ڨ#��t��"O��2�ʈ~�Z�{ 䒆P���"O���)p'�9zD"����R"O����X,O�Ψ����,{z���"OU�V�F�"����&-�&Y�"O������q%h("�ۅ�HY("O���r
O�/���!PkJ1�@��"O���(Y����ʃ�ek d� "Ob`�?Ϝu�bΓ!9�iʇ"O�����Q #&l@+!-�
{+N}:"O�t	��V�H%��!�)A�Xm#"O�!�n�2�n�@%*�1�0X�"O�}3S�����ac��.�y��q�<���!76H��kץ^�hdmKf�<a��߶@t�Q�
ß�l� E�i�<A$*ʢ$��y����2�T�k�`Bb�<��٦8��B���8�VQ��l�]�<a�[=<�RɈ���
�d�o�<�s��|�+��6^�!�I T�<Y��7�p�z'�I"3؂8�C��d�<�き�N=F���E_�N��H�OEb�<��.ȢX��0���2u���)U�<a#�ΆF�A��
S��$����H�<����z
��Ǫ����qfa�j�<9���-eG���4�
��`y���r�<!q'N��j�"$eO�(B���4	s�<�o�o�hj���2PGr�Q�%Wh�<Q$mK)�<�+�!ZN�У�HTc�<��*�{�nUh�n�
�z,�Eg�^�<A K ���{g���jXx����B�<��FE�='���	�\s�!PC�F�<����>u���0ץQ0`��pTd�@�<�'�_�2 
�)6���!�v�<��F��a�TQ�u�����1ۀm@~�<�tR�dn��L��`�JTs$nM{�<I�FS�2� ��ͭ{l�u���SK�<Y����X��d�ɧ'��4��`q�<��-����2�mrT�EL��'�d�[��ۑs`�:Ӣ�*Q@���'̼]p#��n���y��C�6��	�'M�Ȼ`�Y��q�����2aX�'�LI���L��1��)�����'�F�;�뙫9��+ "Кh� �Z�'�DAHfIә�@�J�iF�Y�bt{�'x"tb%�߁��X �E�S�p�
�'L��Z�(�
C'hdz���L�v��	�'=�A�EE���@���ML�	�'�09f�շ2�0 �M�{�|u�	�']JL�1j�e>��(r�}IY�L�}�<�o8Vݔi;�f�P���M{�<��F:Ru�$�4"�Jx� �y�<�ECؙ1�Y{b���MB4+��M�<�Ck
�q5�#g.�:F �*$MI�<����0%YTQb#� �foF�<9�`Ɯ$�2���IՐf�.�0"�[B�`W��)�&sf$H�eŭl�4&�@ł$X��ce 'U�����yr�V�n����JO|�	F�L�y�'N7�60�3%�M�zŲV����y�F^9|�^ �$��F@$��5�\��yBMG(#���'ޏv9�h���͸�y�]�������P��T�ڪ�y2�E�=��ݨ�b4T��y
� ,����]�5L<,3�#���k�"O��nǪ?��Q("�К�ґr�"O6��R��)}$ (w! a6"���"O9���]K7Ƙʥ��44��jG"O�<aI�:LT)kg�($"$��p"O5���
4��i�d��4�z�"Oܹ!��ƫAB������z����"O�tô���U�r���y8�xQ�"O|�cSC^�>B��+ �2|p��"O�]�`	��p2�X�pJ��_~Z�`5"O�M˱,� �a�NR23�]ғ"O�h1� �v+<)��MƝs
><�f"O�Tx��ʺj"��R�P�7 �}s�"O¹��H@�`+�)���:W,��c"O��!�e*����戉�-�8�T"O��2��+4x��Z �B�a�(E�"O�҅\�	�( �&I?{�rq�Q"OFl�� �!%�@�:��� �|��"O��#5���"P�B�� `O�0 "O�TI#�TG�leP�	:j��1a�"O4P��%2���9gjķa�Vt�D"O֍h&�S0
EX&�E��qf"O���p�I�*�E1R+���1z"O����>�:1����%���5"O��@f���Zo�9�"	܌C��
�"O^�A��W�RYk�o� �,�0G"Ot��=N��S�L�0-n�0Ip"O ���ZtxQ��
bH©[7"O�xa$ڲ'
&`���8�V�Pg"O��	C�^�\J�	3 �-��K�"O~A�*ٍ'����G٤ ��ѩ�"O͐��Z9K����S�0��"O2͋"�&t�|#��b��y!"OZ�a�<}�.�Y��VNbz'"O\T�VƜ�b�A'���p��"OƱ��e��B�f.�4��S"O�IءfZ!I�^p��E횥�"O�Uصw�$��̝�;��4ZC"O�+��0����2t�0�ha"O"yy�㜲��I�$��x�:�"O�8RÑ4s��8�M�0o�HkB"Op�����^.<���
��y�"Ov���M�1Xp� )p0��"OZ����-:�R���Y�Q�V��"O�Y�#�_r����п|��A!"O��BoRm6,��c���\ڒ*�"O&��g	5� A�h��]�.��5"O`!��̓7ϴ�J��q�
=��"O�슃��`��de��
��ua$"O����#��Ds�O�0���*4"O�*U��!��ʣ@�	`B�8C"OnTK��֪0p���!I�l�B"OI��D�F�x,���&�>ecs"OP�i�n� �Ҹ)B톹e8$:"O��cي'~�{�cͮ>3h�"OA���!Q$����I�T|H��"OVx``̾54Bp��E�3j�`�"O�az��"R��dĚNd8�u"O���)�8��k��ܝ�"O�m�f�\�� jej"z�rȰc"O�= JP�H�(S�1���R�"O�lۀAC73B8���;�r�;�"O���s/�q�,]K��$9��"O��#�#ǻe�9��^W�is"O� v�X��>Y�N4p3E7��dJ�"O:M*V흦x�� ��/��샰"O���$�@L)�/�"2z{�"O�l=1l@kW �H���s"O�l�t��eM�eXA"cx����"O:]Q�eˠgRR[Ǭ�L���{�"O�H��l�Dt�
ׁX��e��"O�xbB��`P�T�ã�,p�"Oz1 �f�����a()i���{�"Od18p��-gx5Z���o�1�u"O�9�7��	�0HA-A�MU���%"O�x˄&M�4�R���*�D��"O�EC@`�$@���F�m�v�+�"O���ʁ�}������2Ǥ�8�"O�lk߱r���f�]�c�DY#p"O `A5� H�k�l���%"O�P&*Ȏ/��2�)Q�^ �U!�"O��ӄk��\PňY*wq��{�"OF���J�]p��W�ѭqb|�K�"O�d���'�*@1��W*A�X�y4"O=�ѳ_�ZE#�Bĸg�Z� �"OT����35����!ڰq�|�� "Oq��H�d�r�+�@V*!���"Oz�tiJ+X��r�g	j����"O�$���<*T0峵�M�A�(�:$"O�U��GX7���z��lE��p�"O��4�J</�����87��tkS"OLUѡHdO<����Be&9�ȓ'�0\��� �r���n�ly��)X�XG)þ2*�����E�KH2��ȓAψp#�C�0�a�ac����|��Mx�b0��k�]!��n�ȓ1zx��J��a�a�&�
�/�Ԩ�ȓ",HC�;XrEH�L�D]���@pX �(��`?<�b�߃1�.Ї�TG\i����#��`D�x�Ňȓj�����G"O���I�+U�X����\\ �'��%�� ަ���s�+F%A	'�DE	�
���ȓ)=6L�d�+|l��F"�p��ȓI���c˟��}����;.�D��$+8����V�["�ۓ
2N�U��+c�nC��j��A�Ů��ٲ�'��1��<F�2!��O)�H��'��=X���<}��Ibp͙�FQ��
�'��$"gj�V����N�Ez�4��'j��	烇��q@�`�+I[ ���'?P�Q�=��¢�Q?I����'�@��2�,>�Ep��Q.~G�P��'��h���� uضʒ�$��'����@T[PH獇*29��P�'�0� -�(,@�t���
�Zo�ܸ�'9�;��_�XСׁSWGb� 
�'	��kE!�j<��f��x)�1��'��aC4�
��>)����p�H��'h�J��^�\�:8��HнC��x�'��:�D�yT�:�d�>?���
�'�tq8B _&��+0�X-�,��'���D����s�ݺ�,<I
�'S<5��4CT��2C�ٝ
��h�'L*��$�S�D����ŠQ#v\��'�(12BNP�8bB)�4,�<QWBDq�'zA�B�N/&�0r�lP�`� \p�'�l1	�~(�X7mŜ��C��� ���f#Y�_NJ�s�n�s*���"O��[�'���`x؅�Hv�^XY7"O�`ғ�зO��h�a$�+S
<��U"O�)ɤ�X e�~!3�!� ~�g"O���"䊞h��=�p�Э(gb"O\��D�"A҅��1d���"OЁQ�J�M ��Ŕ�	_F��"O�IbE��]�81BA�B���"Oҁ�"'�	z���2��.`2h<B�"O>{ �2]�t�a�(��"O�HPjf�|9���!fڼ��"O�H�ϚR�V�9@�Y��ћ�"O|�Q�E�Uc�i�
d���"O.��c�ܚ�(�U)۳wBD��"O�\�A��C���q�&0�ԝ�f"O0�Hp��%
��K���}����"O�ع�BAPeT����~�j�"O>]6gܯ,�51�^�	���:!"O���D��i�fh��X�d�1"O �Bס	�.5)щ���< r"O�S�i8��(�hV�v�5"O6q�4M\�{|f�PRN��"O�m`ej�3l��]�R/�*7��Ԫ�"O��W��#S�X�oP�/o�l��"O���GC,;���%ό!]`Ĕ�"O�q�D�,8�\+Q��"�,�0"O�L��-�%��5�l���y�"O�4�v�N0����l)uֈ��"O,H�Rl\%7�:9�g�L�s2P�[a"Oy���X(�`]��A�.��H�"O�p��.�75L�a���L.5�I��"OѢ��ʾ�~�q&�S=GȎ� �"O��"j6� 5�1hM/	3�}*"O̅rE#��g��H�q�
�j"O<@Q7F�U�����J	)�x�R�"O�$"&�G�up��I�(Ϝp�l�"O��V�Ϡxr1[0�-J��i�t�<)��V�z�t �T��#֖Pb���p�<)V!Q3x6��9kK�g>�(`�H�<1�țߊ9o'�`�:����u!�ނ%#f���`�=�th�r ��'!�$۰#��^]���N�o�E1�"Ot0��2C����Pm��0�� ��"O��
�'��4^���6mS�Ut���"O����E�~�	Ŧ�\�H�"O�H@��0L�Ωa$%ĠS����P"OZ�
W��WA��1k@'�\|�$"O$�Kcgy�YYu�ݟ2���;�"O�X�2c��L V�Y��X@�C"O���4�-(��'GN��d˵"O^��i��.��hե�)}��hڴ"Ofq1�		 ��$��bX�	���1"OjA�"�-���/�"��+0"O�<���C�C�%�b�ɽE~�J�"O���f-%�T`��Q�?L�9B�"Oq�gnW�hO��߬��""O�)�/�9�hkΛG~��"O쌰`�?8 ���n�43���q4"OԔAn��N�>���o�P�D,��"Ol�r��ޏ+�H�7NK$����"O�-����,l.�҇�8j� ����yPvx��kɌ5�``q��.D4�'�� R�Dթ6f���M+s�EA�'Քa0������S�o�:�`���'�RYa�R�3�����Н4+8P)��� ��y�N���B���1_�*�"O=!R� �t��%���L@, ���"O�C��7Q�̐U*��@�R��e"OF����%7��8�"��hl\y
"O��8#�,Ŭ�s�ےC�~�E"OH�y�ɦb�b���J�=2�JU9G"Op�d&Ւ8Df��D��8��E��"O(5{B
����l���/�}�"O��s��L�
�R�@6Ĕt؎�h�"O@�1%�������S7z�`��Q"O��"�+B�L���&��'� I��"O��s���~5V���#�?��P�7"O�w�@D��ЁC8z4,c�"O4T�#.U�k���ҵ�vF̀u"O�u��2xA�0�P�<2њ"O��rbQ"0L�[r�ȐU����e"O�iW� %0RP�d�(��� "ODԻs�5U� ���������"O�m�1C3v���a�:4�F"O�4BG�$��d�s��p�h(��"O� ���P��܀��Z�d��<��"O����6� s� �3?&�v"O������
M󨡢d���?)l��"O 8[���*]7��k���*�,;�"OBy��@�;�n��b⛰k3�С"O�LB��L	7*�[R�E�$�<�١"O4\z��\t�6�"��� ��"Or!;g&y����K�yypA�"Obx�"�3w�E;�J
lZ`�1�"O�Q
S�V�&!�t�@�&�ڹ �"O��8J�.yJXĚSgS#�=Y�"O�{�,^8�آЅ��P&�'"O�I�,�6M�ŀ�D��
���"O�FB��PO�;��C����F"O<�u�Z�x��	�m� lA��"O��RS�
�Y�&lr��ֽ	�@Y9S"O"�a��XZ R�j����"7"O�a���["YĈ��R�m ��"O��A�[ _�qc��+�D/�!��-[*�:�`�A�B����
�]k!�d��$,R�����bP���j_�Q!��
8|�q��Io������Z=6!�/U1�8�CK׳l皕�tgɥ!�UY��Z0v0�%�Iu!������z/ |+vFĲ&D�,�"O����#0Ť<SQE�~-\��V"O�PQ��^�Ƥ��O;.�2�"OI��cE-b���C�(�Q�2"O`\!F�{�`���B��7 �9�"O��;�N�:urm�(�X�Fp;"O�0 ւ��t$���Y�7ɴmQ`"Ov[�k�:hXpy�N[Ol�'"O�4*�O�)+5X$��*ց#�8�"O<q�+��|01�A	��1^q�D"On��5�Y�&*$�n�P�f�A�"O¤Q�ɾpQ$�ȦMԶ|��8T"O���d��QEʁ��M
hyڤ"O��fEO�m�|��`�Teb"��"O�\H�Y"^��11�M+2Q���"O�e
��B�Wm��Ռ�-A��"O態	
>��)��˙�V��\�q"OD�3N�t�����lH�c�"Ot$A`�ťScĀ*Q�Q/j{ C�"OԈp1(3l�.�0�&S�s��b""O� ܥR)�5}��٦��q���h@"O�u�V̌�9��u�#�V2i��I�C"O��6��Pin�!L�.�Z�'"Or�(r�8dG�U�r-�3���{�"O��a̝�a=n�(�&˕t<8P �"O.�z���*u�ܒm�(�(7��l�<Q�
̱qC�%�w��G�h��C�Ok�<�$	^�A��U�L��ԡ�Pr�<��#�(X�h��H���)�Fo�<1�#R9N�Q#����W� (�)�p�<)�E�	@��l��.�!Wm��Vȝn�<A��'R*�C�MI!%��A��f�<qЅ'�"�yC��b4 �^�<qB�i�Bt��*[=1t0#D_]�<Qg�6:|@]�$!�w$f����d�<q��0琥%U�c�D��o_�<Y�O�z��LB$K���d�D��W�<���/_��<#�[,=�m	��w�<yA��4��)�ٻu}(��3�{�<q�Θ�-�N����ޫC��� �p�<���ۤ5���Z4+N(E��]�'ELQ�<Is�Ȥq'f���JÛn�0X2�Þq�<��'��fV�U��MZ�Y�r̐��5T��� (D�P�0� J��Z��bc1D��˒@��q~���������L#D�`$�ÜPy(��ec�92� �%6D�$�Um����H;�!�71ZQ��O3D�D����)|��ЀI�J�����1D�� A/�%7R��c�j�W���	�H*D�t�4� -��
ȥv:45�g;D��ҩK&�P�D���\�h#�;D�h�ub�%�@��LV���R��8D�4�@
$q:�xjl�ex �Hvc+D�|ɠA6f@X#J�6Ĺц,D��r�A�1E;�4���Zw�� �>D�4��kZ�kS��R#OچVhҹ�À.D����l҄iIf�Iq�ęu�V4��-D��ЅO��"�`죰�&���dg)D��*âVSך�Xr"�yrTO)D��h�B!B�T�ꡎӈ	?>]���%D��q������2��.�Xh࣪%D�|F�I�.5���$��*B8���#D�4��c�+�"T�ҩ'9�� �i7D��C����M�^����G#�P#C2D���ց��S���j�$T0%bA@�B1D��*thݔo�\)�-�7I;8i(qi/D���t�*�PG!�?�8�ۂ�.D��z��M$]y���w� �B��-D��p���.M����=�G!)D��C�Ҁ1,d�i�AN= ���$!"D��#�ϵC� 87�&�P��!�=D�|��"��*��A��Ϩy`�x��:D��Ӓ���P#.
�[��[��9O6"=Y �S,

5!�$)TU����r�<Aa"M)B}�a��'ҍ�,A���LT�<���M�&6���Ѐ�\0R$SO�<���@{�>HY0�<ƪ�1Ꮑq�<��`Ԅd*�%�i�d�!"��b�<�4둴`��$�b�?��DĎX�<�B���fj��i�i��7b\�R�<igb�?P訋P��e1�,�R"P�<	ԣS�Dء%�ێ�VԨC�P�<A� 6G�"u���U�&Uؔ�@�<��C1
0�9PUÎ-=������u�<� l�c���e� 2`�40X�E"O�8p�
�&Q��	���
[�x$R�"ON������│C�v�u�0"OBq!Q�p����A��=!"O�@�C	�(7tq8�N�"t�"O��Х�7H�蒒��3(��s"O����.dh<<QĥG�	�M2d"O4H[���ԫ�A�
�@q"O(!�DO�3r�������P(�"O�� �C�I`���4���X�Jd"Ob�I'�\Ŋ�c�R���""O�x� )F�i�ᐍ�0�
d��"O���0F�Gh� u��'�p�"O�4 �gQW$%�
+I�����"O�)���|�Q����,�^�Q"O4!���9���#1��=,f�"O<����v쌘��f�Q^��v"O8����_hڽY��!zߠ���"O�}J��\H�t����E�~=*b*O�M�!cf���E�	�"P�	�'�z�g�*i���*DM̦m\x#	�'i��"�KLӨ�Ѓ�.v�D�#�'P�@r��T����à��3gA�'�X�ؐB\�!T ��V3^�����'\4�Idh�O�n{wM �V�e��'BJ�V��1Q���2gD�&�̰�	�'QT�3��C(݀��#���%!�UI
�'M�|j��I�d�`s�ƿ����
�'�\� �]+�B]��O#�*(��'���kA�_�?O@L葎��"���'�� j�B[�g�8\�V�N	(�֜�'�����e�#J��Qf�ͺ!yx���'�2X�,ܳ��0�%�ݕF���
�'.<�۷���<�f`h���1;�d�`�'K�A�v��,�l��Ǡ�8:�0c
�'�������I$Q*�P$�	�'׆@��DN�U֘�� Һ�a	�'�чŁ�>r�2�d024��'(����ף�E{$�D<n>��'�h���_���Q��� y+@���'!��)�"�t��(�fC6Dj����'�L� ����}m��xG��1>kXy�'O\�6��+o����W�3�q��'Af��A&r�����-�c�~0�'a<1"V(��4������X�`�	�'�b1�u��D�!�'+T��)�
�'��EQ� �TY�UM�2;�81��'P�I��2�KmN�/�6� �'<Hm��K���Ĉ{���o���H�'�<L!�㜀 ~�DN>kD�ܘ�''�����19��ϙ�U<(K�'���k��k:���#I0L_M��'�d�
���7�j86�\Ib�@X�'���Kd�A�oߵu�d9	�'ݒ�(���4Mv����gPoK�-	�'0�!�2L�Z�Z0PD���V8� !�'����o�ؐItFGQ	>�*�'�R<�PB��hC
�`�ҥHIh��'U � �k�:S{�J�Gя	�����'�| ���'�Yc	�uyj���'�:�#Ё��Bh��,Vh^�ѫ	�'�D(�ɜ8Z�p�*��ŕf�:�z	�'�rpB��91Ny9գÅ/��h��'�|=˗���8 .�it�HV��չ��� � �-ɍ $*Tb��!��@"O�(g(��f����91p�iR�"O�|P@bJ^�b��sK�;we��z�"O�\�c��E��5@�珮KG����"Oh���X8/�);"��=><x�A"Ojmң$�o����瞒7��0%"Ot�pĉ�!dv2�X�J�.TZW"Oe�I��S0,J�ǔ��r���"O�u�#)S���Ʀ+N	P"O�h9AD̩�qNɵZ"���f"O��Ԁ��#�Ȝ��P�Z@�"O&�Q�K�3b�����&��$˓"O�MۦL�A3���wj3�0c#"OHqv�B�H��
!�:8��"OPp@��V��=T�:�@ :!�Ra��3� _�`�XMA�& w�!�dģ;����p$ѠBR$+�O8�PyRnF;2�"� 'BB0��ѵ�yR�B%EdU*r��P-n�XSf��y���6�\H�W�լC2���3�^��y��.
A����D�b8IC�%�y��,5S�9�0j�n��=zF`��yA��&t����%de�5H�4�y�!"JebY&�X4a�Z��!�y� �\ E��n6.	���Ӡ�"�y2n�)]��8�ɕ.�z�Z�����y�ڳ[9b%Ib�D�(�x*��N�y�͙m7�L�T��"��X��Ԝ�y⇑�KnZ�Ps[��p
 ���y2 _��<��!@��0t	��y2�H=tK�Ö�����l͒�y���$���Cߛ���1�V��yr�Q�Ц�{C�Ýq)Px�@�<��A����ԁ��b�P}˂EPK�<iīM�{���*�%�?u㦔����Q�<��)WcB��
��z���Y�<�G���Q�,!r�	H=+��^j�<�L.1H��gd��y�֥C#Di�<1��(��y{5c����If�d�<a0F��d8�L��h�N���fG�<��K�5�y���!UȔ8�4ǅ@�<�3/�����(�|XHAC5r�<q��˙|<.��WND�~҄I��je�<�2��9;��)� ��kr��3�Q_�<Y�ǚ<i�L���R)\�����*�W�<���;� AP&6:֕Qק�y�<���]>����J� 0�D��R��j�<i@Oƾ4�nhi�^��H���h�<�ƈ%%���3qKK��-�R`Ae�<��`��`�xXb��&�(qf��I�<q*MTL�	�'��</h��FI�I�<��!T�J�#r��rA�$��m�<Q�fM��z�)��=u����Dg�<1F%�aRx�S��ʵx�Ċ�c�f�<˗�J�"����/qE¹Z��^�<yҀ�;v��8�$F�kn�ъ�$@�<��NةY���q���35��p�D�<qD儂
\��T����5q�M�u�<u����drqo3E�`AMs�<Q��<�Xm�v�ՑH�~1�s�<ɥ��zK���O��(�83mJr�<Q�IU(�( sD����R�4��y�<1�I�-XFzԀ���k9��b�x�<y �Z�L���A�L��f��b׀w�<� �	wG�H�
���;��	1"O��[�jX1QT̨�c��a��!2"O�0�MS+u����&�6Z�� 
�'.I��f��ahB�y�\���'Y�y��͐C�C'��l�Ё��'��$)���Z�ظ:�O�9_^���'q�H�B�`�V��SJW�l��'��I¢N�l����%V�U�F���'K.p	$Ĕ/2�Df��V���H�'Mf;$^��������l=��'$�M��#�s��26*�(
�E 
�'8pGJ�3�}b�����@
�'���!nޠ��c�^~�֘b	�'*��s�1a�:�ÂS� HTPr�'@�٠���8��%a���	t�1��'���Ģ�!]5��QDN��HS�'^��rb�3�V@[Q��)4����'��$3�͓%dPՙCiR�C+�j�'��Õ�/MФa�F�5��y�'A��1RnM@̪y�b��|���'3"\�0�I�!���0'A:y/�UI�'���b`�E�Zi `�6qB�9z�'�܅�!��(|���l5��9�'�Z����ڕ�㛒�b�#�!�Z�*b:t�4��_�N�1��H�!�D["ȤUZ�G���"9��)̄-a!�X�"�Ê�3�ܠgh�G@!�[�t:���%�1[��͉G�˗a$!�V:(�tab�M^���s�O�:+h!�l�Ai�%T��lA�oEYx!�DY�r��]at_���M�K�� ;�"O���iB%jz�!�"ȵm�4�J�"O���s�
F�b���3#h��"OX��@
'\���z��*\�C�"O�E�-�N�L��7�Y1V8�z"OQxan?+����`R�M�nPi"O�q���
Ә0Ӥ��h|l$��"O.�w��U��Pm�(]0=�"OԌB�*��?=��Q���1=���"O*M@���_f�����ԥw�ب�S"O�i�h��l�!�)�
r��E3"O�MW��nF�yT�T��Y�2"O2�	�I{0`<��գ1Ӟ�6"OR��bɃ"mm*pbpDݹ/h�y!"Od���Ǟ O�ލs�c��q�nLї"O��)��/ ���z�� ^���pV"O����|q|���`�5�|��"On��3��$��1��۩>��x�"O�t���0<���v�6"]���"O0���
F���[�.	RZ,�!�"O�]Z�nY/k���� �ų@$��"O���@��l�Th��K۵n "O%Q$�ŕz_d8@#
AX�B�"Od�7�Ԁn@XX�ʌ13����"O&��Rm��q��1Qr�?j�����"O�I�U"ŕHz��cb��N����@"O�
�n.uj�@��<>�$9��"OҀx�G�!9("���� "R1J�P�"O�MrC�$�ى��Z�J��T"O� �@'ʈ?HqY�߃0�"�P"O�lba�Һc�4�At�ɔ�H`#"O8usV�y��u�d"�"~X���,D��C��T?#3&$�CL�;�l��3/7D��bS��KB���S���SC�X�t�5D�� �%�M�$A��Б�K^�7�����"Ol$ 0��~!Fd�e	�F�Р�"Ob@qP�C�v�{�gF�~ݘ)!�' ��U��%��`�cm
"fEl\	�'+�h	���=r�����թ3[���'��E�� M�8 '�ŧ)?�4�	�'4��H�%Ӧ*���Ƨ��>���'nfɐ�G��G�T�f�B֐�
�'9����=,b�P���ݓ
�')����k�.[%� ֤�5�H;�'���"@y�����M�-�
�'j���g�Q�Ϊtc;H��	�'|���5݌YK�"^�9���'Ѡ�:e��w<E9��ͣ%��X��'��X7o�8M*vC؝� �`
�'U,Q�`�7��3���=��T��'��i@L�:Q6HDȓ˙
�l�'���b�Orv |s T7|�r�
�'������^�H�C��h`l�	�'�fi���
��`���M>0�3	�'����M���H�㓚,�lH�' �i��*�X%��h�#r���B�'���0W���f�H�p��=�08��'��!I���j9�ȣR�5.C� �'kJ�I�X1rQ�,!���3%�~�'����P�M�4`�bA��>q��'R|�kG�
,_&`@�	��,�Y
�'����NX�;�<y��Ά�D�~��
�'1�A���5p�Њ6�a	�'�ֵ
�N�xê�N .<tMK�'�F�9WHŢtҤ�SGA�5���y�'�����cI�]7���6o��y����'Q�	�(F)�ƌKq�q��x*�'v�9�H$!U0���Hk=���'Z����Z�s���� �+j�ʝ�'����"@�䴘��H�aD�y�
�'m⤑@bجz*�T	�˛�V����
�'�`���KY(���g]�I�^|(	�'l�|c@�	>��LJ1JC�)�����'�V�
�J
�"*��I0 Y��:L��'�rp�MˑH$��0c�)A�i�
�'?��r�K7�l�0�]�Vn-��'Et�"�J�I��Ipj]:_ެ�I
�'�p1�GʍL��*#DUl�=Y	�'�ʘ��@O�
c.u¢��Ȱj�'g��i�<ǚ�ue��]x�B�'���c�@/n����"R�
4�Q�'i��U��~2�FO��b��'$�y�qo�e����kQ9}|�@�'�  P��%^tz��"�s�$�'��X@�Kܟ&��-��L�zȈ���'���2���\0D]1b �"qҔy��'z��"��d� ��4O7�<q	�'��!V�C����3�5�F�X�'�����6朢Ԣ�.�n���'�.�@�^Ehy�T�Y�v9��'��Lj�U�'d� �� _p,�
�'�V<�v�׹/X���&�ĊT͔,[�'��4��^�@~X�s� Y�Pt��'�H��M�	�~d9���c�����'�l%��&��!Ѻ�.%` X��
�'R�$ V52�@!��Kl6Q��'=�e���$PƐ�$"CG����'j}�� ɼ1"1�v��<Q�%��� ��Τ,�d�1�®�y��"OD!�D�59��@�R�J 8��X�"O4�k)�8oK\��@\'�<Taw"OTը)����b0�ɸa�z9�S"O�u�E,˨G��f �	k������lCq��W����'l��T?����MTt;�f@�^i"�K���cG^����?��|#���%�[�rt�����\��D`>�^�6!B]�i���%�.��}pa�
�h��Y��	�W|�0 ���v`��`�2l�'�I�<Q��p�e�*�`�0в��O�oڗ�M����i�tکbb��H���DҦ+G6��`�S��?�,"��߸�r��@�M����I�M�ֲiʛ&*H�l����s=��	ׂ��~�c�I����'U�W>ų7��ПH�IȦi;q*Qo*Ձsh�h���5��6�j�X6���6���/V�nm޸��?ŕO��t��reJ�@�b<����G	(;�$M{A�iOZ����(��6��9S]"���U:�xd(rÂN����D�p�Y�2��T�@I1h��	�2�i�=���0��z� ��+��Ż�͈�bB�H�+˲#��������bX�p��ƑB�n�+�"J�l8v��ҁ8ʓW>�-w��O���ݭ�&*�:L �9�HA�6RQ�f�
�?�����< �P����?��?	�S?Qm$p]1C픀<��DQ���p�#d���v�� � *J>������:c�:qM$����dT����B�����̮8�d�fV�%j:��ˁq�$�ƞê��P�zy2��
z(����@*�B�(��Scr�ӿ�t��Φ��uZ?˓�?ɬOR�h1KD'����s�5bP�|�"O�0�ȗ�i�2�дc��5������L��MC �i1�'���OJ�I9mhH��(Ή`ʊȳ��S&�l��@�J]���I����� �%Nȟ���蟬�Bx``!�̀�[u聊��T/R{���i=���@P�/�Q�Q��)_��̓"�+:��	 f�H�Vļ����=�蔺S��V�d�kU���+�R��c�@3�qO��V�'��&JǗ}��5�7l��{-p�C<,��<%�<�ɀxD��?�;���b?6��H�l�.y�����y�@֯v~p)h煁 ��WC��~�%f�Zum�Ny���Hr6-�O��$�~�'�);q.�*'�H�Y���ӌ ,	.D���'���'ܐ�Q�FN��xK���b�F`2@k��|��D`'h���c#`i�CAc�'Y�q ��8$R8a�-�9�F� ����u�]�\�����<���&��E�<���$I"2�'>��,7m�!@���C�C ,n򍉷LNl&q��T�S���� �z��#%ѽZ�BT
<U�|"�sӰW�9�M3�i��W�,�R�Z+{�{��Q?�&\2h؛��'�bZ>�r���ݟ��I���CĮ��1(�1dmӚ#^�aT�L�8$����S�����U�|w��7h�?�O�����LmJ��XB�;�h��6LBQF�i����n�'D���X�$��}��8���*3�x��l�H���V��73��¦%[�����i#��(�+ۛ��~�d�D.�禭ء��;�v|���温��`?i��?�����d�Oc?���ȓ�"��D�^��lR��/ʓ*B�iO�'���Z�eJ��ME��Yd(�
H�<�K>�ۓEa8I�  @�?  �쬙��ۜy	��z��L�<!���7�@ĐP��$4#��ra,�@�<��e�4R�"]�e�e�bd@�x�<����x�� SGY|��@���z�<ѧ�R�d�\q#@B^�P�§�x�<A�	^��	�K�/a����[�<y� BN�)�%��xFR`��P�<9h�*fah��p�	!��p:#�H�<��ݏ6�� ��>ON��Q�/]l�<	 �3i��Y�n�Ao�$� �g�<�vĭn�r�a��9L���a�G�<� BU�ybN���;GzYY��Jo�<��O�8n$�җ��4��'��S�<�B�\�&Z@H�,_�O��{D�L�<��_�%{��W��#�4���E�<y��Wz5f)�&�%\]T�X��X�<�ӯ/J��#���
��Ӌ�y�<����8{� �wD	�0��Jq�<i�e�F���Q�)O���\����l�<�&��� �j�i sw����h�<��J�쒄�笗=��9"�k�<�� �9_h$<�֨��$b�|q`ʙj�<�a!A8{��9���o�-�L�<� ��9���4<�@���� 1b�ys"O�(��M��G�xi��+<?rA""OD�Zѧ���4�@$�\�2�"Oj����<Vib�3F��R*�s�"O�iа"	g�Ȭi�"Y"\�Ub�"O�|�mF[椴�爃P�\�qs"O����Wz�9�0�"�څ�"Ot;A�J��DA*X$�|�"OJ���O�.µ��l� �f�R�"O�=Pĭ��^�Jm���-	��"O��x#�C�=A�T��Γ,a�ཱ�"O�x" b*�h�9e�V���z�"Oԥ���?iL`Yf�A�7霅XS"Or=��� V���z%KǢ�~� 6"O�u�V Y��*9��)��g��"O�HD��B����A��{�`���"OLĉ�*�?	��*��E"hڮ��W"O ,5�0�6
9~��0�u W�y�̇$e��<�`�� x�(����_��y�+��h�K�酯v�䓦 ��y��6�콡#��_�,����yRN�,���BNӮV��-�V	8�yr�:%���I���ܜ�e��y�I�4�F�d�2�!tCؿ�y�Y�i�
m�&�	2�FU�U1�y��BfV�zR�{�e��GE��y�e׆q�ΩCd
�l�c�I"�y҉A6t����
4g+Ta�&珟�y���*$��Z���9(�l�ʠ�ԡ�y��ڮ9���1Խt }� �ڎ�y��0�j��îW�r4�)3Q V�y�OQ�nDDW�M�eb�����P�yB�A�B�\�Q��aM�1�G�J��y� ��r��h� 'VU)Zq3�"[h�!x�m��To���)ٔ.)@���O�7mI�l����b�e����!G�|���X⁃�]�xuB1-�M�$�3�,�5��^���O%k,S���|��W�<8��W9fD��^�TG�|B �R\ ܴvl�ܫ�jɐhI��C#�|�12ӐĢaG-Y� l
��3FN�l�X4����Ħa��4�?9���i�t	ᠪ^�ZH3�뛡c��e��'��Q�����}��#S�M3�49r���b"=��4q��V�|�R?*�$��2hdE��ȉ'D�t�'`���?��)F�h�KT��?A���?��B��.�OJ7��=P�e��1f�Iуb;`��a:�@V�g=
qKFE�(F%
%ʒ�?a5�*P;�O�pj�nF�d���q`A��7�n%�1�'5�@�Ǌ�Y>%I�h����S'a�б/��w�����Nq0#�I�/�>��!4N2��'�(x����?�1�x�'�R��+@�!/�HQ��?�������I��%��}�� ^?� �� �g�E��<6��ۦ5$���?��'b>	�3 _�m�2 �����ɡ��%P8�چ�'���'��B�m�R�'���V�f��8���	N� ���E�!� i���ԽRb���������j˞aZ��S�\��VPz��͍9��h;flH9y��q�BcE�y��`�+��s�XH��ˑ�)QV ğ|��<�?��(��TC��F
1�&$H�Ȅ�:z:�ӿiBV�`�	ӟ��	Z�'�H�B)�R"�e��>I	콅�W:d��i޻rS�B#��<7k
���F��S׶i�I51��h"��O���~��Z�>�,\R�Q�6.��H&�q����'L��'qԍ�G�����)�9 V���#����s$j��n��"�ƀ5;�Aa T%�Q���1*��~��0��a� Vܥ�R�ؓ���ņ�_�ɨ�"X�+1|�Q0nY
���WP�	�
�DЦ��۴�?9���⏙ݥ��Ţ��Kǲ-���'B�O1��O�KS��j�n��������%�'�"6����o��C�h���
�9�ְ�2C�c����#��|q�O��d�|BDo;�?����M�vC�� �h �[i��x�I�3EF����K�*�&2���E���jgD��N��P�r.Ch���O'k�MqT�eGF0�h5���"Z��ŀ�3جt9�a7��]�V�0.&�	�+�`I���\>�ظiܼ��&���vz��M#-�6�۷8�R�u��lןp�O���MÇ*ݍ7�εbN�CUR��f��i?Q�Ű>��gU9�hI��5�x%�g�'��7m��&�0�O���ǈ˷,K�e�q��`�~Ђ�m�O��߁�z(�Qj�O���O���F���i����,ޔ0^xt 4��]��ڀ�M�/�2�as�D�M.6m��hn�)�< nD�CO.�� s��nES�L�5,����$�̹��� [�&�^$�L_9F��ӞZ�F�h�W�,��|ɤ�a�h[��*�(n/����'��1P�'i�A�,O��d�>�	*�b<�ᮂ+P�bR�m�c�°=��hU�!���F%�)Bg� �u(�
Hw|7�B�A%�|Z�j�?�$�讱\(� @�?�D?f<)�2���'l&B�ɈZ�P�[�F����Q�(^�o�B�	#����dU\������ZG��B�/ L��⓫*Kn�(ÆX���B��(l,.�[GHĆ�@e�5KY�GR�B�=B�qi�\+��b@�3	��B�D>�0�&c	(��F�us�B�	� ��)Ӯ=����1c/A��C�	�@K�A꒫X���i�A-��dxxB�If��<⡎܏y.���E�1Zm@b��D{��$��>�r�b&�Ug��4�Ӓ��<���$]PMr�Jǖg����4瓹x!����M�sLL����#[bn��T"O�d�q�>I�����8"��L	�"O�|jM�8@ƌxpAQ���)pO\i{i��2��=ɠ����`��9D��r��ԔM��5��Àe��}��7D����; � ��<L��w�3D�4���;XVi��E���VyD�0D�ɱ�OUd�pʷ��M�j��v�.D���$� ����@i[BCU�B�9D�{p���x��ݨR�:)x�"D��JqO��X�h��Ů�x���C&j5D�X����'[  �� �N�Ƹ�wO2D� �$.Y�Q�Fd1�⍫8l4¶.D����ߔ\3~dy5%O�z�2L���&D�6�V�/Jl��Wj�!.�LC��#D��)Ve��pU�����i%D��	5�X$gJ8�8dɅa>&D�=D�$��7	��"���x�� ��M:D��s��lI����,� ��W�+D� {W	�.5�Y�RJO�6�9��*4D���t�o��i[�b�*&P���3D����a@�Zx��tHT�e��(�&1D��F��:�$T����%M��� �/.D�0�c)��p��|��hת6ϖ$� �*D�8�G)���&л5�)$����!=D��X!V
I����;c�t�	%O?D���ġ���Ir�睸``����0D�$�6l�N�Zɰ���R��P"�0D�,��L��<��ԅe��1��.D�(b�'j��C�Ӌ��2��0D����(٤3�p0Ԯ���q���.D�PJPJȉH� �.�30�Ҍ�Tc!D�p�B���n�Ђ�Z~�d�� D�|끋�#����#o�=B�%PW�:D���t/�7	����eZ�
����f$D���Q��b~m9���_&ڙ�3�6D�P���J,,U
ÊV�H^�@�3D���1 !+���5e��%+Ntإf3D�,�Ɖ3"�<���A�!�<XyuD=D���r�=i��*�`O�s1����<D���7#?�$�c��|\�����:D�h�Mt���˙D���0F�6D���hn2�`����[w����'D���m�Y��A�$�Ҽ����qh3D��#�B����B�6���F1D�\e��9����~.�1p��0D��gԪh�ZS"b"��ˡg-D��2Q�wp>����1.,5!d6D�� 
��3IF���,�.jRPˠ"O� q *�=��(q#�L�9gv��"O.1Ĥ��s��H@*]�5QU8�"OQ�6nH�$�`E �	ڙ(��i�"O�t���ճ%)�b3:����"O��K�i�/�M��T<"P�x�"O��X&kI�zd���!X�.
`���"O`I�Ɉ��P�Ή!J��Q�w"Oܽyɉ DP��g-H'�@��@"O�I�Cn dժ��q4"��"Or�2Ώ��x0��o-<:D"O���/r�왂���=M.I �"Oj���H���4PD�B7h�t"T"O�Q�#��^��c�g��{�"O�t*�Z/wv&d���̀:�,�a"O�m)�'ֻk7���Ϭn�ި�e"O�@+��N�\�4�(�ڡOʮ!�"Od�:��]1d�1a�'��:-s"O�4�0�I�Fg����у[wƠ��"O�4�$�2U����@v�F�!"O�Bp�j�ƍ��*�Bw"O��[�G�Mx�Մ�9���F"O�`P���YE��1��e#�a�""OT��
�<�Z�X��
��A"O,�^�����,ˆ}�,ݳ`hX�<E
�(ز���#W�J��Kp�T�<i�HȽr/��V��1���[��O�<-mNR�0�U�ܬH�G	\#Q�HB�	�}��j�M�u`���V��
jB��:)s|�0A# q�hLB���B䉖1ЖHu ���6�Z�*�:5~�C��	mFx8VN��p)"�Q�K�MȖC�	)}�R�ڶ��"��Y�h�b�rC�%u0��F���{�$��R���XC�B�	T!:�kJ�A�V��j[�B䉍?�v�z!5��a)D�a�B�	�F/v��(*�5*���yb�C�IMo�����T�����}W�C䉵Uwjuڐ዗x�����]�.�C�ə&�$�pGJ��|�f�!TC��G��U��O$��0y���1�B䉊'�F5�#���<0��yU`�-q6hB�ɦpwh��Vh��)u�5 �Jϒ-��B�I�e�����ߊ9bpQ�",�o��B�	?i�A�L�%0hy�B��q��C� n<4Yɢ�Έf��AR�#�c¸C�ɫz��}3l�%<Y9I
{`�B䉛j
�Lk��^�(g��hN�<	��B�	�x���C���Lΰ��τ^��B�I1�]r$��*0ÊIm4�C�I�}��,� ݔP������9ky�B�ɨ^'^L"�K<B{�-��&��Z��B�I��YR�Ę/p���bF�*��C�I2c���h�R,yFi�EdP
!��C�I4&�d#�M�y ��B�K.�C䉵�@i`�ݴ\���zQ���Q�C�ɻ=^�ĳaB8R	��9Q�,C��C�	w�NM �i�.��锩8b�!�D�G��`�5�	�MW��	3�!򄊳Ϭ��ql��Mՠ�	ť�0
!���$��䕘m�-2e�30�!��X$#��4KV@�[��(h��@K�!�$�6���v��>�&�� (�� �!�ԊO�,1".қR���s�&��J�!�� *�Z��({�ܚ���3_��"O���w�<f��;���*�u��"O��ibݱ;�f���
09�2�Xu"OȠ�7�TY-���Z�D��dC7"O�|9��
,�eð��:fd��"O����Cܛd�h���c��pp"O�d���F;$D�S�ڜP���"O�͚�a
�/���2U��V�R�!"O�h����018�s0AD�`þyi"O��ag%��Ox���c�u�&"O���]�`~`Ij��K�ErԘ�e"O�L`���:`��e�B\{����"O��!��z������zp�$��"Of��`�� w��0���v���B"O(�c�E�x=&U���!N��� �"Of���+�zr����(����"O�IɥA�1L���H6y�LS "O���-��f~�I0g�+�����"O�u�g��hh���Gn9��"O�Y���c�������js6�ن"O� K#k\�p3��zu#b�m��"O<d�uCͶ2`}�s��*-�ix�"O.=�G] BW�d�@�A�u7����"O�K�6i6�aD ��lA��*�"Ol��T�B%'H���E T�#��-��"O��CH8l���B���qP��p"O(�V�Lr��M8!#�14l�hB�"O:�0��y��FaX�� "O����'�!�*�Y��˝*~1�"OJ��5J��hT	�	~0 �*w"OiҶG��&�P�H�1<��s"O�]����t� 1SsE�~&�ԡv"O��!�#R�����%FRN��"O�٩!"��
Ԝ`��N�`a��"O"4�hG78&9cU !=�P[�"ON$���:��I #��I�#"O��z��� �T�+�!T���b"O���J��2�q����|���`"O���N΂|��A�t������#"O���#��6Myp�bּ}� ���"OY"G��8�[�kQ�VW�Aq�"OPi��O���IJ&a^�T����"OTDR� =R��rt�ɖ^��Lcs"On�"�h6�ㅮ�F��w"Or!���3�Ԁ�p�K�Etnd�a"O�9���Y�ޠ���z��|��"O��� �[0Aj4Cv��$YH�L1�"O		�HZ���
cKܡ}bu�"O�-b�	I1W^ld���4'�fi�"O�����2>x X"��d�H�"O��� cǒl3���3	�����"O�z%D�;Z�(��
��4�lȻ�"OP)�'l�#���C��Y�?�|XE"O�p�caؚ@K\��QH�&y
��C"Oz<��AL=9�(z���{��|�r"O� 1%���W*�T�#HI�K}0]
@"OP�c�ME�^�����3(����"O���F����4b� u�L)AQ"O��V(B�D�q1��at�"O���wkV�Qo.U�B@S�Df.��"O�#fI��C�jPRiʃ@P&��"OD=Q���#\�0d�2gX�m�P�"O�5qb��m-�5��hӾrώ�A@"ORи�b�-�>�#ԧ��A���5"O� d$hHMcs�g����Mc�"O�Ib���5�X�ɴ���t��"OB����-v�$d�GAtv�Q�"OJ|
v�A=��\���h���"O��r�BΚ�<]ȴ�_cd�Գ�"O�y���iLHa���I=E Tz"O�x:���=Y��0�N9@���#�"O�`h��*��x��K�B�X	��"O��ҩj^���WŐ�M�=p!"O\P��T���U��%y��y"k�`��Z�܎b!�%�d田�y�U� ���`�d3*ǲ(C�
��y"`�.)��G�+$B��:�� ��y��Z��t0�&�+<UaN�y��Ki|)���ɪzǲ��g꟟�yb�S-fR�#�;=�v��V��ybiPgd:�2H֜HX��-�>�y"�ޛzp�H�բ��v��EI�j3�yBÛ�2�R�Js��%xhD��D �y�A8,��@O�r3j��(F��y�O ����bX+h��H�0�^��y���>e�Y���ҜX�xUc0��,�y��X���<�&�G1
�uB`��y�B�%G|� �����D���I�#�y2�C�f@J�� uC���l�<r��\�v�[��:T���3�CED�<��Ś	L���T�ڙ��}�<��G+%RhR�D�35�� L`�<��\� B��8u�/ �V����]�<!5?�@��-Ԥ[i�m��[�<����Ahx���Wi��He��[�<�2fY�Ov�hP�͏V��x���O�<	�lK_n����T(�% VK�U�<	��0/V੐vG�F���k���U�<�vk�51nn���ꐂ��LäTV�<���ެ�d"7�ʾx:�#m�U�<�Ѓd6V� eޔ^���F)D�@뷎��WFz���ߜ<��㑢(D����M�BA��fd k-А�%g:D�l:p�]�tk�I���ن�y5�:D��B�k��E�vU��F��[j�"��:D�sX�44 a��XV��T�S�&D��3���g��`B��9N�hx�V�:D��QeȾ/�I�U҆s�:H� :D��9��`�jIz���\���=D�xc/��mV���N�,�/D��3���u-����ʆmD<���/D�8�B5y��@�s� ����Fm;D�\)2@3T&���@�81�#f�#D��+b��t���D!��[p�� b!D�L�7$Z�;Dݪ$��k��hC�  D��QόR8PAf 	X_�P��`>D�H�%I�&zm��mK�D�h٤�;D��a�A�9�`@K�ꊇ:�T���.D�ܐ����	���w%\�V�T���g-D�T��m�!t�9�cސ|�<����)D�$���9�z=)��Χ|�89��B'D�����lڕ롆���Z8{bB#D�`�bGO�žܘ�`��C��*pl&D�{ �ߠQn,�K�gL�{?@��uF D����-Z�y�3�
������+D�D+b�P����iW`�zBA�צ%D��3ᄋ7��sdꖆ�v��'  D��cQ�W�)��=R�FǸw�B=J�K2D�� �4r��T/�1#�
G��8P"O|�eA������'ۦA����"O:�`�<�*��Õz,����"O~L��O�l���	���?t(L#"O�l��V�&��b�ͲHPH�	�"O�}6a�[��IP��!0Vb�i�"O`}�Cڊ]�AH���|Ip) "O:aa�#��N���%�G�=�����"O2��Ӈ��X���#��;@�"���"Ot!8�ޝ)�\*�
�����"OJ����)j+N̑3*W�]��|p"O�!�Gk��s� ����Ww����"O�H9�cգ ���1Ս�xZ�9w"OxX��y�.�(Э�	 SB�(�"OLY�`��^Ct,@1OC`�d"O��Ch�P��DyGK�~?n���"O&\�%�6_`�E�(G;j�۶"O�ͨ3/�����1���(,Ѫr"O��A��Z�YHt��gЇ8����"O�q���;�{af�N:|�[�"O�8&��VCAZ�eL�R/���"O���@c�+}&�y&D��mBD ;�"Ob|��MI�a�Y�e��}I��1"O44�5��p:���\6S6I��"O�,�舆=O԰7F\�ˊ�r�"O�0��_ŞH�v�гy�|ͳ�"ORUHQd��8��Y�r@Z�D�2�"Ox�{b��4Ɉ�� �йqv��3"O��R��0`>,����O7Ut�|��"O���D��^l� �*pLQ#"O��C�Џ�4	��Mȑt���g"OTc��	1��jqOӽPߤ��3"OL��@��C~���p �=#̩�s"O�b�X�!9V����Yy�*�"Otɫ�@��uVt�QH�&���p�"O�1Z���$�,����e�U��"Oh��Tnǣs���(�� ��l �"OB��#X�x~���ⓧ8&AAe*O�	t'W�?�Zsrʌ��x#�'׈0�u�$`�(aKRf� C�xj	�'`����0�|#S�]I�P���'�xl�P� )K2xԁ2O'SK����'�2�p�ĵ/��r J�;9�Y��'�y�e��(���9ʒ~4D��'=J��̜.c���+&τh�'���XƄK����*�0t���' lQCEu6�����*�D��'��Uz�ߧ1d�|klSr�\��'����K�;�^E�S��%�T�J>�����$4�L��k�97���'�_)�!򤔷~�bT�Ɗz�C@I�3Wa�8�'�f�+v�F2\�nehG��"#y�'��UЋ�qK�@S���:���'s��z�-T
 -�`�N�x��U��'�z��#��^L T�GI&�`�'k�B3��#�n�f#C�<^T͓J>a���II(f��PK�c�δir���ZQ!��H�@M8��GW/n���1fk��0G!�W�g��q�RM���q�6L!��ώ?Z�*��W�L���P�QT!��Z�,����@21�\Puo_�N�!��-Wt  uh.]��p�����6�!��^�:�N40d�ɿn}��� 6�'ў�G~��7k�Pp�v��,5Vx1*�dG2�y
� �����D�T@zP�G�
�����"O���`� �d Z���V�L�0"O��YuF2Ìa�����M�T��q"Oܴ���� �z�c���8j�nID"O�x
��;��ѳp��,Q��f"O�dF�ѮadѕG�8aĮ���|��)��tI�X���;;��̒S�W�DC��;������J�R�l@P'g��z8<C�I�g8$lj�·�eKP������C�I s�n�𲏜J�^�A�/�%DC䉯rU����o�rU❜o��B�	%;��BE�I�]
Db���o��B�~|#a�ɇ��e*J/U��O>�=�}��$q��p���!�¹����P�<����(^�
fD��\)EE
L�<�QM��y6qi�Nš9�X��C��E�<�l·$�x��c�X��h��D@�<Q��B�����Ĭߚ!W��R�IW|�<�@ �Zphg��+2��Q�6(�_�<��n��Gq�J2m*E�h ��K\�:z�H�?�}�sa��.��8�uvp
�D�W`�<qte̢∀��f_�b-�QP4��U�<Q�.����֜<; 8լ�x�<!��ƥJ�F�*eC�"9H��C[�<iE+خ+�T HSeK�$U.(�ׅB�<IC�2KL����>K�7G�U�<�	�n�+�S77>��*p-��o�'K���i0#����D�mJ9�%Fԓo3!�"h������ۈ�R$�]��!�D�?���ٓ%�
n�� �B�T-k!�d�>F��H%B+���C���
!��u���&L@�SrvP�GB�S!�$�E& ���%՟8���
���(!�$��,�����A����T4C�'0ў�>y��GzP��ّ�ہ ���g�,D�$�kل</��Qc+���*)�gc8D����(�"ש;��a�#7D��
��P?uj� �bS�aLހ(�4D��HA F���T:�gP�"4�hCe8D���S��&7�����B�wEv �­4D���늗2b���0�N���%-��(��|z�O���U�á	F���fA q�Pd"O��ȁ��$S��;�j�rԬ�C%"O��Af��<bi�����"O{@�%�x1i5�����6"OHS�DY?)ġ[�M��U̘p��"O8)1te��gq
��g@c�p
�"O���b���}�j���H&!�j))��|��'��Oq������3�4I��ڍ_�XiYu"O*��$2A����:tص"O�L"fiƢK>%�rą`�x��U"O^�����.�d%�0P�N��"OZ-zу��F��1oQ-u�*�#�"O��Ӷ�q$��0΅:==~�c"O��h�$��H�<�cc��u����"O�mbE�1T��s�炔-M�w"O�[r�@�kc�=����r�ƝXT"O"X�2d:i1���� yy��Y@"OZ��m%?QVa�u����"O(I��.ՂS��Mxt@-�޼jP"O�|z4.�Hb4ps$/( ��ܚ�"O���ci
z'(�pu��
����7"O�3`\�M��[�m�G�ę��"O�%� �8
BHݩ�2l���"O� ��R�(��;H ����^(d����A"O�`��
���nq�`	@�J���"O�9`�NM#�\� ���,Eǚ��@"O�<�A��y�L9��O�~��\��"O:�k�P����Ya���"OB]�#L�A�p��C�.(N��(�"OLԻ`�To���&��*�r�"Od
�IՇ��{6e�u�e�v"OP��iT�e-v��u�F7L�J�*O���@d�-�a�����X{�'&�(�˝�IP�����>�9��Y��@�Uċ��س㇘6�������p$#��[�m��>{��ȓ$e�W��bm�Xõl\;J�@"O�L�7�$��̫�@���"O���2;�v� c�-/+82#"O��Fm:r�^�Ԁ��"fx��"O��sbM�)�B��w/�q����"O0�e	|-���׮�(��a��"O�%�,���z��.��_�d��"O��Â�x"����ǡ^��"O�֨I����A挑�f%RW"O�}�!�e�$�G�6J���!"O����� 7�T<�� �{�:�0�"O�xHA'�9`���E�k�(��"O��&i�eJ��@��Z&&V� �"OX��f�A���cH�_��h�"O��s�H��_�� #,O�
�1ae"O2�@'��NM,u�תЂ:nh�"O�0�!�(5V�؅L�$�8��g"O���)���x��˄.r�$�1"O��p ��II�,�w��V7PX�t�<)#��h=�c��7L�bE�$�BQ�<�7�PIEC,v�p"B�
*���X��Eْ���pp�c-��]��Q��
?��x˱L����!��'���u6ݳ�`�g@(X�Y*Q�����1�4(PsM%M&dM�
8tM��T̀�b,a��ν4��Y�ȓzyb���Ȕ�V9v)i��='z���1_�a��HH�y�
Ք���ȓ!��3�%��'uP�qG�,2|�ȓi��c�,%EFѠ���,�\�ȓh��7�R�$R��(%����'�<�`f�8�8�B��7*�(�'u�h�C�[���chL�~��LY�'�TY��-�@����*�p��'}`!i@�f|��e	�1�B!r�'�<!�D �:?M2ݡď�&@���'R���Q��&p�*H��ǆ�*��(2�'�^<�V�^8`@2�<-�R
�'=�1K6�]�l�>�)���J���'/2��2�A�1�]���ޮ|;�'��8ՆWB���sr	�~r�J�'v�:p�Y�_!�1R1I�n��'��Q�ǫȰfԌ1��pl�Y�'=v������sY@p�@LM2o�d�
�'FjAs�F�4=RL�-O�/�8��'٠�J���(m��zBj�*0�r	�'�"\ �\�x��X�V�׺Qv�i�'�")#��]��hQ�j�*R3�#�'�^���(L����{ �W�KE�,��'���;d�=%* �3�\%
	�'�0����i{x�P��®I�	��� �=�Z�yײ�KT�֜
�0$"O�5�2�
�g����`��Y�"��4"O���蛥#���x��D45��!�"O���2%A9a�1Ǝ����|��"OT��f��h��q'�F>n<lb�"O�E1HF�*d�A��aGQP�|�W"O����nƼ-Q���E�j��d"Oh8�U�4���a�7j܍*�"O�Q@��F�@�T $/
8fXN�{�"O�{�hƢ.�@���D�[��,�a"O���CmS��Q�T�5��T�"O����I�s�a��P��A�"O<���#�3k��E��ޢ���"O|=�ulR=��P�u��"�"O�!2d(ًF`�`f͓�
$Qa�"O��87j��l0F��3�Y' T�"O(�Qݔc��u{rm�S�@m� "OP�P���
.�`�b&��ud�9"OK_9)����'�LA:�L@=�y��!A���W僔<v���O�y"�S~�|�`uE�T� Ӄ�:�y�h�l�����$Ο�`�c$ƒ�䓼hO� ?YB��:| �H��J�p*Z��DΘj�<���Ơ%vB�ʀ��IwL�3 �c�<9a�ʲ-q���Ӥш8i�E"$��_�<�'�R��hiv���p����E�b�<�0�[����*s��f	��PnRW�<rH�I��=�V�D-(�`�"L�<a'�V8bd��b�ED3��l�s�<����:ZT8a���M�̢7�q�<�@jߕ.��	a��N=K~Ax�ĕk�<���!����EčyʤTpe)Yl�<)����(�ެ�U���`y6�#S��e�<ٰn�<LZ��u�9h0@u�Kl�<�2K�<5�b��0�F?y��Y��@k�<qW�Ut��AP�ܲsg0���+�e�<9��,R�ʦ�+V��Mi0e�X�<I�.��T�A�ɥ.��ؠ��z�<	��Ź���H�K_D�鶁s�<a䨐90Ԛk�f��?������]F�<A�X�qv<̳��#[*@�u
�]�<���7i%�<�鋩=��ՙH�S�<AF��Lmn9
Ba> !�4�CřR�<���N�i��Ц���&OLm˔d�P�<�NF g�!��ƷBS�l�E �K�<��ď�Vs��bS6d�J3d��C�<����1B��)'�'>0��F �C�<� �����#���#�h��$"i�<q!ٹJ��#6"�"J?��!C�{�<���@98ʘ|�􀔞%��j��z�I���?�}��,Zb��a�T��6�4Srʟ\�<��쉯7��`��A\u(u����Y�<�1���.���	��;���fHY�<�G��3�qc0+N�bh���k�<i��ޮ)�z�RW� ,ppYT�\�<	6@J,6���5B޶;��I�	Hs�<!�E��iYS#�ip�h�lGo�<Ae��
�if��9���("�G@�<����	d��C���vX@����~�<Q�
W��%�DL²�M#V��5�y��ֶy��Hh�A��a��}B� ���y,J�<��0dQ=0�85��y���?��ࡂ��"�� ^�y�b���P�F��~e����Kɕ�y
� � Re��+2�(!�e��4�F$��*O�(�B)��v��`��rVH��'��i��Y<������p��r�'����bg+<h8b�Pe�-�'�`��-(Ğ���LH/
t���'��hZn��x�M�`Ą$k�B�:	�'29d��p��%����:,���'��ZqoQQ�f��H�)[�
ti�'��]	��ڐ8�̘ҦHҬ]/:��'(z
���=��&E]	����'����UٔB�l�+�aU�[�X�'%Ԁ P��X{��:�hUL\�́�'e��@�vc�hKǃ8�~��'`���M���|sf��zy|P�L>i���i�i�p��@IE�y�潲��]�!�Ks5숀�b[�@�F�1��q�!�Ě� `(�O�:�Jp����tm!�:���i�� ��<K4�8"k!�DR����PC�3C�0�IbB�O0!�dКV��Y�҉c~&�IQ���?'!��P�,I:�n�,)�B	�a�X�(�O�˓�����i��Ֆ6@Z�g��E=�B��'�!��
!>�tа��L4u2�h#�L�!��H	�+֥R���R��W�A!�dT�7�\�f�Đ-�4 �W��2,[!��Y/�Hr`��%j+N��L$>!�D�O��@�͚$^ ����f�!��W� 3��E�O��x��	!�䙓�zYG�Gm��ӣC,{!�T\�νh2'��>�F �#	�)1p!�$ͼ5�~�����
G"))�̼m!�|ÎD�7��O�Mq��!�d�@u�L�8"�i���Rx�Ć�`���p�ǥ�0˷��X9��_��Y8gC�3UN5��S� �b��Ddma��D�HT��ŗ�	�݇�	F�(u�ߏ(�δKHҁ���ȓ(8�P�g��iW �ېeǶg�B���-�~�aOF�.1���%O3i�J<��d�>�Y�
K� F�����_԰�ȓr� Pb�H�"���s�R��.0�ȓ�	)a�I�N�����g��$��C�����Qf��ă���JU�ȓ]��X�ь�^;tI�C坻9�\]��6�����x���3#�+~Ψ��T�d]��NQ�j���j̐����ȓJ�p5��u0�-C�]�]�ȓP��p�4�[�|<h�h��v������P�9g��?0�iX���2]� ��vQ��J���0y�  � !�H$�TF{r�'���Ӗ_���{��O�}=�-a'-@6.�BC�I�
�Jt#�U2ʄ%�@%�:�C��?�:�,��D��.QxjBB>D����K�-%<����
M!����<D�X�t�M|�ޱ�CZ�B��Ò�:D��a"×f��e % �)]�5��9D����JYs�$x�d�&S��,�b8�:�r���]�ORޔ�!�*$������B:@�ܱ
�'�	Z"!��,m��@�c�>���'A��00Y*n�R���26�|i�'���qL֪0�Д���z��
�'��s%�֜Ｔz�F�ӆXz	�'����%��	�1��	?f�Q	�'ˀ%*B�L>wb�����V�y�T���� � �� r�j��d�Z83b�x�"O�E[�*�xI	��[����Z"O4��R�C+Ɉl"h�2r��+�"O��/���e3� �?&j��(7"O(d�M�5�\s`�EMN���"OJ=(Â�7k�T���aN�=7Fe8d"OĹ�� #��Ւ@�6G���p"Oz�j�'\�0�b���/�[ʠ���"O� ��+�(UG�	�D�C���`�"OhਐG�(=ƑbūA0"��"O�B�D�p���SM� a�.�Y�"O�����33�v�Č�h�V$��"O��iЊ�	t.q��T2X�T��`"O�UH��^o&����X���RQ"O�hb�
�}��q�؊0�``2�"O�=0n�<�2f.iܶeK�"O�l	W'_�-$��)�'T *ؠ�sv"O�ⶢ�&���
�:�8�,�!���8lĜe�eo#7���$셢1�!���r�@=hF&Q�_/d��d�k!��u!D@�"�! �$�3�X5!�d�W�B�JcJ;+r��lMQ�!�ā�H�l��օ�,h:4(��y�!�K�7���7���24� �� {!�D��$�:)X�AΥm������Ũ`!�䊰LtHyy� �N�<�� ;Z!�d^�*?p�U����
�a�-K��!�d��ZC��AHK8F�ȹX�C�!�d
�J���ڳ��<���P1�� �!�H)��h���"N��qkX�F�!�D42�z\�2ŗtx!z�˱=~!�;a >mʳ�� �x��)״r{!�D��D(
v��r�����f!�)>�X�T��1�,��ӄA�n�!�D�+ ��[Q�]� °� �CC�z�!�$��J�I��@֑F���YPb	�1�!�d߃4��yP��~�P�HV`_�4�!�Ċ.�Ȱ��K̆O���w�ܶJ�!�D	�m��p69oƴ@x 邪:�!�>3�na��e]�\�����i�9!�!�X<(��<Q6�+2P�@�t�L��!�$1<�]ru��g;l���� )�!��=��D Ы�%���q�EV��!��&fR�ӆ&б"R 5h�dʊk�!�d�'��1#b,U��ԉG+Y�!��<V�Hw��?J�4Ԗ �!�$�=^�t��b��{I8�(�O�F�!�J(o�J�y҂^�*R �(P��&�!��z�lҗ�E�%DNuP"O4���2m�V�sVa�*E���p"O���� �����!ޙ-3F9B�"O���V ʭU2T	����&@d=i�"Od+���9(NrHb5ꀀ���"O�*Aj���8�DiY� ��$J3"O�$�"��T���x��Ք%yu�d"O`���J��V��0�� '<(}��"Ob�+���E"���U��$Nq�4"O�T!���% l�}�7�� ���"O�R�a�88�<�sh�:#�f� �"OΨbR��)��!#�&J�B'�Y6"O$�G"ѵ#30�ҥ�Цxn�x�"O��XD��op���3d��6"O\i�B�B<c{����(�t� 2"OD#�L�}�Q�1�H-|�La "O� �E0�a��qK8q��>�ȩ)�"O��8i�7c��آ��1U3�M��"O~Xb��i�TL
6�Ҳv����"O"�2"	�!��!�fJ�gq��"O�(�a�Ҭpr�p"��NT���R"O��	 �G"h�X�q��0=�X�"OD���C,��!�AD�}!�Ps�"O���i�&7��@E� tf�Z�"OL����ȫ$<�\s!Ǜ���+"O8���X+�i��XH��܉t"O��r#�� k��]��CU���;�"O �� �IV�!�ˇ5^��c"Oh���#&�x[K֘q2D�t"OB�Zg��N�,
T��.�`{�"O�E�CY�����ڥI�> �"Od9bÃ�#.D�f��!g�`��b"O~� R��8"1�$з;�<�W"OR(U@у;��t��W
o|"��Q"O�Q�P�2�y�m�m��e"Ovݠ���{`�拆o��0��"OBؙ�i_4~�&9����;=�z]ۂ"O츫��T�dp�O܉7���BG"O2}���C4zq��`$�����"O��;d!]��.�Ӵ
�Lndi2�"O��8�؀$ԑ�	^	p_���"ONx�eM0�؋ 	��l_T8z5"O��ڵ��]��8C�F Z|@�V"O�p(�kZ�H�8=p1fLO&��"O<��4� S��c �{Mv@ C"O:�P�(W�%�H�6aP-�%�0"OBU��MZ�xs�m�#͘x�V"O���PU��A����5Iw"OhT#҇�Ca�B�
�?�rM��"O���@�D�m��`�l��`�J�"O��
�ۊ��*ϵ	�N�	�"O��2Q� ����x�I������"O0mI�,��Q#BP����u"O��I�j	a�q.AT��DPW"OV�'�c�@��'��N$�pD"O�B-=xG��)Ū��	�"OP��_x1H]�3*۲JҔ��"O���"V�_^zԡ��ˀ ��1c"Od5�/X�Ak0���� �4��"O�e�f�*TT�*����^���"O5��L�+����J�)Ndjlk�"O��r��ۅ!w����ʦp]$9�"O`8x�m�x��%�x��40�"O@(K�)��H2B���JАtba��"O�E� )[�12��w ��]��"OL�6���laa���i�\�js"OD]�4$�kE����R�@�c�"O ��@!P�B�H��n��p��"O�5�s���\dR�n}Dl;�"O<ɪv�54U�:�#�(ۨ�D"O�9��J'��k��A�V��U�	�'�"���L՞~��8{�!��_d^�'��𔎓��T�8�F�]� ���'�h8pP��
ٶ���e͔�F�'`�'태q�4(a�)�����'ot4���1)���a*����'A.�� ����4�1�\�~et���'1H��GM6P��(!�8{�F���''t�YG��#3	8�#"��~aVj�'e�0������N�R���(��@���� ֜���G8����-0`j��E"O��pE/�&8n2ؑ��U2f0ҁ�"O�z5�8B��1��<3Vq�"O�=0E���Ey��(Aa�|6�M;"O�����;�x`���$�u�!"O�4� Hɸ)�F��pNBV��;�"Oܙ2��ӂ%�xY���K`r�!��"O���"[3�єMАr�f�G"O��G`V ;�.��FQ������"Oȹe�<F.���"�y���B�"O.D��A�>\��٩6aG�F�ڃa'D��z�ȃ$U��zQ�\�e4�����%D����@.^t��D��~ 8J��&D��K���M���(Uu�I�J#D�,��M�XWV�!ը@,fix�{ƅ D�����6/<@"#k�8�����>D��Qt�D0�X�R�[f6�yb�j7D����Ξf�
$Q�)
TA��(5D���n���)k�;,.�pj1D��ٳ�V�o�6��5�X;sؤ�.D�@ �6=TT��!ɼG�Ơ��:D�L	u��!6��� #�9¾ ��E8D��[!��,�K7�@� V��*U,5D�0���}׾y�Dm)	��pPO/D�T�� �SE��PYk!|���,D�|b��E�>�z�餩˧oPJ��3�(D�ȡ0�ݐR��#�E=d�FTh�L(D�$0F̊BC�q��k"K�� &D��w���=Tx�ā52�HC("D��0MC�����4;D�$qP��g�0�w-�.��Q��9D��9S`�,aagn�L����j$D���2��~J��D7�0`�Q�=D��s����3�T9�ĩ�@�8`  ;D���M_��,��c�=% T�!�%D�|��&v�.Q���N�*�J	�p�.D�$B�ƚ8h����k@���g,D�4K1-̧G���R���'2YT$�1D,D���T�G�nM��qs�S�8l���'D�DsЏ��-|��h!��H���'D��B�,�1�f�{F
�}ID��'!D���C၀GN�L�v��[]r � D� �U�*D�ΐ�μ��{�*O���œ�r�b�1U��6=���˰"O�y#j��cS\q!F�#q �"O�%�p�M8I�jhI���� �"O��e L�:�I
��쁥"O��� �
�6�v��2ω0y�F��"O�1"���b/���ˉ�����@"O����Oڗ7�,����2�byP�"O�!�`̥%ٶ��f�ƾp���!�"O�8ِ#��\z�C�ПZ����"O��g@�!e���W
ͬS�V-"E"OJt�S�ڼ"jB���Z�R�t ��"O��#+�mo^��H@e����5"O&�U����0�i��/�ʭcC"O.S�ٝq|t��GgW"��hR"OJe!�B�C�y;6��I� �д"O�m*�`�8Z�\t"�M�K�	�"O�S���]�4��G/#�l��"O`�* �S���XV�Έ`�H@�E"O �[�A
5!�s���ɒak�"O�,�Q�G*i�0���ʤ!�
�U"O��c��^�C�j�ذG���%��"O� �U�͇}�p�&�p����E"OT���JU�10 �h��%0Id"OP<W��!PL���O8Te�`�"O���  {a��%*ѱ|N4؀"OF4�T/^0e�*iShR�
zZ���"O���GY�,�u1�ӧAu|��"O�(�P.F aK��S��[R_
���"O�!�3e��	P��H�.���"O(��C�]c�(� �JǼ�˰"Oft��R�
|	�i����"O�QeZ 5���P�h���4���"O4`�f���~vF��$�L'	����"O|i����kѼ0����b�3�"ObQ��	9L0DA��+c*y�b"O�uS�l�1p�ҍ�S&M�&W�Y�"OX��RnB�2 P�0�2CH�+a"O.Hp6�ѳ3ީ��f
S9:�� "O� +�-�"�Ι[�l�;s�p�f"Of�)%MI�@��T���Ql�t��"O�]�Q,+��d�2���`���Q"ONE�W�ʻG���Q��B�8!8"O���	�5S5�ՉVdš/����"OD��$�3�~��A�L��N��P"O.�:G� H�H1��g����q"O�i�_�uʸ52f��$]�B=�"O4��p� -#�BE�qo2�Vak�"O����#��~3eA��X)i�$U�"O��х`�.�`��%h^�T ��u"O8�`f�1\��I
L`I��"O��E�YTb|p  Ι0B�<0�'}�`���� b�q�v��c{�!�
�'<ѓ�)Q,n����B�T�*�	�'!j��Rl4Z��@Wd�D��(�'	H|���D=������80`��'��P���*��a�>,,@��'_rP�-V#@�s��(�(��'y4��Sg�Yö�ȅʔ.v1+�'�p`��!˖e>�@��0I�JP��'(D#��.��7�����'7n��#�1RN��W�	&�hc�'�$H���]i�hK�,K&,��h
�'S�=)��Yi����ڛ̀U
�'b^I(��8��|#mOh۴ݚ	�'�f��gI�(<��誃�s�L���'C�LBV$+�PhkS�"s�RD��'��IF�Z0]n�<@�(�"��|!�'� �Àl�0�aÔR�4���X�<��D�=��I�,
�/N(���IY�<���M0A��r`׽-f��ҋU�<!�KX7*�J(`�D; ��x�6��y�<1v�'PH�(���A�v�@	p��s�<a�� )d��r�ʲP�8$A�Oq�<�ց��X�B��)v�b�c&�i�<qĐ���҆�B#-!2���K�g�<�'���:P��
�-Ǻ�(��Rc�<��m�9O5���E��&�`�F\I�<I	�/FA����A�)r�D`bnJn�<y7�˾��8x�cN	Q�Pڶ�GS�<q�iJ�7��h����1k���yQ͉R�<i ��0�JI3Bj�&>�r���Fx�<�hYU��u)��N"����j�y�<�ˈ�>�zF@.�9�A��{�<���p��m�"�ϖ<��`��l�t�<!�D�T���#F��p�AăUx�<� �-���K�8�yBi�^Ut!Rc"O6���j��ja���I�E��!��"O��#֦
"�,�ʳgW�g)�UR`"O�4�T`�1yʝ��EїI�u��"O�`�`�F=z��ṅ�"a���#"O�S6#��n�v`Z6&]�Y]PLJ�"O��qA�"*`�kw�P�)g��i�"O�Eb%�ŁH���r矅3e| )0"O0���eE>/851��L4V��a"O�d�a'(v sGE	�1��=�e"Ob��@%D�#eb��儹R�J5y "O(0��%�"e�rx�C�ΏMz�@�"On�Q�ED�>�0E�7�L�P�i��"ORx���G-m��I;v*9��A"O�4��#�<q�B�z�K�@b��U"O�st�z��)��%��/�y��)\"�[��2W�4i;Ҩ���yB%�9Z��0�̖3T�H�D��y�H�Dh(�dY0H]�����D��y"I���AÖB;F-���jس�yb@�=6����D%?�<�"#fL��y2,߱~β�����>�09藯��yR��X��0��IU,>�̡'����y��YR�t���/M(X3��<�yRK,�`9hѥ�8ZP�a�<�y2\'7䖔���	�*ũg霱�y��9i ��iAl��p7H� �y�HŔ/�l�)6B
�yj�P0V��y��̰L.���� v�*�p�
��y�����J �C�����"Ǥ�y�
B&I �K�:)d4,�ѩ�yb� dfԺ��A5'�.�s��y2�J�� �A�lA�oa�a���y�nܙ����d�^ m��8ZcL_?�y��8֮�[�i��a�D�CC�M��yB���[�J�rHZ�\~�J����yRJ9L�,lp �L,G�y��NR��y�lV�E�l�ZW��Aϐ���h?�y��ٴ0��b3�9L:l��`4�y�B�\|�8���$~�^A���Y��y�ν%�9���Au>J�BM�7�y�)�?~���ɗa�ޢ1�Ԧ�y�mE$���ɣM��?�A���y��]J1��`d1~�\�"&O]��y2!ޯ!e&	��f�m�H�ۢ� �yb��}��$�g��ը"O����^(�|��dƳYK���r"O�DSEC3����p/��K@vA:W"O�����\�AFR(�h,=&H�)GOL�H�$٬rw��{�k�4IRp�W�C+9!��Z�Qrn4�G�K80�H	���Z�!��Ybo�@��վ0��`EI�k�!��զ>�������$���i�!��ϫx��e�X�[�d��`2#�!�$�-pP�rsE�c�4�YCo\�(i!�$����V:���䃭Rc!�ΑyT�4����2$��LR䢟3e!�$зy�0�Jq�I,J��8��O�N^!��I�Tw��§)ު��	@�/U�V!��'vRt��/����L餯�>v�1O��Dƞ?�2Q��M�*ŀE:�� �;�!�O�P���g����-�3"�x��O ��Kkx��B隺~�~��po�J]ax2�I��.]��
�,��-��/�����D2�)� HۓG@�@���J��J	w��2"O&�Ԃޮ9cJt �J��V�tDpA"O�`�:���EI��gv��;��'�ў"~���
KЬ��W-�De�d������'U�{B��,(@�9���6;�������y�A�<I���kE�67��H�8�y҃T Z�l�)d�1G-*��s�^.�M��'붡Fybh;��kVy�a�H�(�I7`�;fe����<iփQ3C\��"���f~�k7�CP?�F2�S�O�JD��7A|-`A��|K�5*��D"�R�⤆	7u�8X��ѿ2���"O␚,�!�iXP��<֒����'�ў"~
΋<,p���ψ.~Q�ܩ�G�+�Px��
Ⱦ�I7�#/���C�
O�}�tYmZh~�9O"�i>q�n�I�jU[���:������ֹ���Y �Od�B�vT|���l UbE��"ON��qk	�~Q
!�e��kUTu�w�>��>�S�'h&�h�4� M���z6��D$�͓���@���!���PK�Ę�S�Hk�-!�I'eAazB�9��]�I_���1�8��x��0/D�EsA�X�=�j�3Ai>���=Aד}�=K ��:��=+!͌vs�ik�H��+%�<��b/2:d���J�N�Y�G�6@dI����Q%�?!��qyr˟���K��I'X$t�0P���'��z�'�`@=R�I��I�n�p�0�HO��/U��Y��œ�J�$�J��A=�C䉽�����b�!.
�v�ӱ/�4O���h�%Uq��y`�hM �R1ꁧ��m����V"O����L�%V����d�v@W"O�yp`���0�(i	���9g�nt�"O\s��S�tkXe�w�4v|iI�"O�p��$��+J�Zw��M�<m+�"O"Tئ�ٍ0svQ����3	w����"O�"��Gl��9�żk�ј�"O��*'f]"U��l��+ھe/�+d"O|`�b�OJNl���"-|�A�"O8�4l��6g�}葌�	<���"O>�Wl� f�"��=AvB��'�!���#A��t1�Ũe����a�!H!��*�t�$DFۜ �ů�ya}�߯?�B�@�r�K�-��y��o�;'���p?ɤ�ۘ-��9��
�b���1�f|�<�`G*A�(�[E��4��%نL�!��'?ô�S��\%W����Ԫц,la{���-ge�I2����Ffju��J�Od�U��<ˑo�"%��Gg�S�2��*D�4�!�W@���e�Ȑ���@$D�L���
�Q�C�D�A 𴨂�#D��*��ԒZ5z4��>z}�p�A
"���➔��I�(E��Ì�rX��$V�*�M��Z�4��5.�'6˨ ��ᅎ�����8���@e��nƂ� ���kr)���?1g�9�4LC���q�L01��R�<�I_1\���`�DC�o��Ƞ�	�f�<����1h��G/kaT����]d~rV��F{ʟЀ`�NU�P��ib��gp2���"O~�RJ[.<GH�{mj���"O�q���} 1��' ��\�C���u}R�S<|�r��4�6��ō�A�'C��F8�T��*�s�tJ��؏)C��StH0ʓ�hO�S?�R��q�F�T�	q�gŮ4�>B�I�Z����&�Z0�5k�N8Syb�O����G���IÁ	�h�����\ar��ߟ� |��n�?�5RqӓV�4��?O.���LW���``�V�p0�9�6�P;<�!�$�o�T=��Q�&����MS��D:�O�7�r�$��̜֠O?0�ӡ�'����q��0b�G��`����\�!�Ûh������i���xҀܟP ��&���jA�@A�����瑙�,]�ȓ=~��J�I��x���t�r4�(�'a"=E���Y��"�۔ 
P�
�JBF +�0<A�<�O��p���h�<����!j������=D��Gkƒ"@��K� [0(Ĉ0@�7�OL�IqB�(�B`%����H�fC�I"+��#�X��)��0m\c�̳�)�\�;*����'=X��rf���[I!��] #tRH���f��:q�D�`|��U�	%yHax¯�'=�n��碁D�T��e�Ԯ�yRa��C,�W�A�A ���X��HO����٘.�8�9��[P���{� �!�Ď6%��R�M��-2�c�)>�!��Ķl�0�z6EY�J��<��d@�[���0F���Z�W8�iUȓ�l,�];�$�2�y��G�ה�@'G+z�.�	����y2mF�m��AЃ��wE()��.\���>����~��Ŧp�D r���-pa|]yg����y(�4C�޸!ag�Q���j�`��y���I������M9bѣ��#�y�@�&-�LɉG��E�P[� QeYў���i��4GE�n���Y��ЍV�ZX[B�"��ȟ�i���/�|PH�DU�#"���"O�$�Խ$A���/uh�s�Of��&�� ]�T����*٘DpTO[}r�';�x,L�g?@Db��,�Ҭ�
�':I���h��Q���ƴ 	ۓ��'��Rw��e�)���_����ۍy��)�S_Dt �Q��?c�ƈK4�A=	*B�I�w��u�+�!EH�|�CG�."x*B�I��F���ߊ$�:��F�r!��hO>�rf�Ҏ�����#9"@�Tg"�$�>�˓;�c�f�s����`@�5�Nl��>�p��F��!SbP����1�JA��1jB䐔��.C�eZ�c��+̪��O�'�L q��U�:p�pe�d��ǡ/LO"�  FG�*M)X�qF�)K��-D����O�#vh]���H­Qj,D�;�Ե}t�`�F&J^�p�&D�l�#���H�q�Ȥ	�8����2D�p+�#=;�l�ŋ�T�ʴ���$D�0�u�ކwJ��5�EkE��e�#D�LX��M	`s&�_<5���"D��ʥ�._D��QE�B5?A03cH D�0(��E�v�����TJ0���3D��Z1ᗺz���G��]H��6D�ʓK"rD6q��\��!u�0D� #�Y�(��m���Y,&�`t�3D��
eOW&E��X�
$*��D���0D�X8��ǂr��EK�<C��d�2�1D��˷nY�ߺ��`�W3O�p)���=D�8y78B�J�b �3�|)U�<D� W�] �B�{�%��U����;D�tˀq洑���Sr"��#l9D�@r�Ā-H{�h���I82��V�5D���aG�~j�|��\J�B&D�!���<"��X�%�c�<$��$D��l�Q��@���b�h豔	"D�� $e��,�
h���J9z, H*�"O&0%I��.���`��$^�ð"O��	�J�q��88�C�8�!;e"O�e�P��i�L�rg�T/$�k%"O�)���{9�}9��-DK@cs"O�����Ի>�����b�����d"O U1u@�/;�$�q�9	�4�C"Ol�a��� ,���yt`�~��y*#"O�m�AƉ=9���k��Uk�P���"O��P�Z�1�H1IR�֨J�`��u"O�LxG��
ˌ��r.C��pLp#"O� 1��A�5ȖH�0�Gq_�=�b"OD���/D�L���s �%~��	��"OPա���:]��9�UNݏ���B�"O\<RT,;=MtxڀK�45���s�"Ox��#A��"��5*¤�Hk�1�U"O�M��I�$u譣�W�&`���e"Of=���$C��hPrH�5sF��K�?O�uJ4jI�"��aK���>�x�e��?�"P�v��1?������gE�C�%HVm����� I�D�87�B�I�$�&�eH���������^C�I�#!�xk�E�|G�( Bᜭ!��C�I�l�P�Θl(�ăw	��+z�C�ɢ)�P	a�%�*7�P�Å'�2
�C�I$?2�t���Q�]�Fm��Á0 2C�/lZ����1EVu:AAPx�|B䉅|���i#�G�O��]*૏*(�B�ɋΈ4�%�_9*O���' Eq�C�	�^P��Z��×W����&�)�B�ɔJ �	��"�4^����'$�h�B�ɪE��e;� �!=z�|1w��9h|�B�	#]1.�J�'���xs�GH�lB��DXb�K0L�ܑ�C�I�B�I�\� ��ީ+9�����%�(B䉟r��p�GM�_�Xp1��כM	TB�	OUA�Rw�}��W�uv�B�	(ݬxs�Ɋ� ڥ�0I�/��B�	!�&��7,ýb��ձ�)B��fB䉋0U���� &n��,bWlߩ�l��;,�\�'��Dd�����װ(2e�V���shC≦)4�t-.I�"�1q�uF�=�逊L� Q���5��O�8�y�`U���E���@�"�x�R�'֘$A¨�7=����A�;���4$Je���9QWx(��B��"~nZ�T��AE)�*?�HH�ą��B�	&u�z����/͐� ��V<iZ��:���ز쉏��8A5��?�=q���IKFpq�&Ԅt"0
��`��HXbáS&�,2!��	�� q�U��*���_+ZA6�����V�a�䀺��3�
=K.������'���t�A%��W�Qh�xR�<��N�."9
t:�)	Hp�"Q(@��y�j�$9�a$��LM~�`�X��Y�� P�C��I�T����ٙM?��I-�1��':�"fl���@c��'��'���@+c/0��p ٭m� �(���%�C>���H�	$Wre�A�_ M-6�G}�;E��H�C �+���������HOz�,�#Ag��9 dUcz|�cƁ�1����, � �D�!�M
'�%����"j�� 2$�y!t� �%�	g�r����Ⱦ �*���F r� y�H�*���3r|�f`Gl�b�h��b/	�%�$��7]?���A*�A6��l�cb��9�剘Jx ���p��S�O�� c�#N����i�R�&�Ss�9�@D
	��)������$YP\�4o�(]��ɳ��8��#A�أ���'L�1�AZ� 	0��Hg�$�O|n��>;*��^��֐a2����d��Z��Q��י%4�e�� �L-D��P!�t�IR�dȺ\gkLߨu�2��6?��֨ bT�bw���B2��@��bU��?U�py�G�X��r�,@(W�>���
��G�ra�T��;6�j$���W�[���a���H7~�k�[��*�GѯXP6���N�/K���h%'�-��=�@�E*Fe&���jV3UyX츢�ہ#N�:��î	�~=CU��/��5訟�n��k�J�@���&�n�*��05��f��Ab���W�cO�~r�S�S�D�r7$���`�TR�#�,DTJX���]�t 8y���"?���E�m��i
�O RjPcʯB[Pl�&��'r9� ��b����0��mP6!�~к`�gmL/e=���gB康-ʄ���z�á<�K�,�I3c��[�& ���v>�`/Ĵ,���k0���Re	��b`LK�]�&<�vC� �A��i�uiv���e�T��MW�kC�M]ފ`�F��+��9�TU�p3V`$�,r&dR��0:s$V5g
J�)�A�2&�ؠS��5IĽ�rÔ4�X c���&>@Dݩ/1D�P�υ�&�ր�@�%3E�7MF)����D�l��� }K�8H�E��8q�pXtkV^���g��P_�Ry�X�뗝Y	��ɗ���wILx���R�I��
t-:	 ,Q��R�
�
T��݆|
��Y��w$��`��D�E��@�ڼ��	�[��-qEАu�A�����,���E�`]-Y�[�l*��'[��51�}�}�6"@�)��3t� �K*F���Z6�	B�t���Ġ)�B�1%�8f*�`䯁���G�
斉�w�=TYj �t	L�q���F5ڗ�դf�p�� �AJy��#~Je��׍qx�aDT��P�7��& ��Iu��j8�Bd�	o0� ��YP@D���#?&��2;��Ȗ���ZA�\��F�b��$�3��/Z��v�9>�:��[s��,���iKZ��:H�R$��2>��XٷD����ꄐ����w'z�#����>y���k�2�t�G�3^��q��)�h ��M N#r�;��L��ϿK oG S0�}���]yÈ�B�C��d,@�Cޅ���g��2(}.x�'R3�a�0��Β8����<�.W�)���A$χ+>���qJ�N�tY��ˋ�D�v����^�����O]�,��4)8����*KI�je1��$���.���G�36!��N��� �R�@�y�,����S�ql1O.���Ó#po�0��[�2�N�2��~�,p@F�#�?!S΄����e�K�=*�N�A�b��3���0_}
̓R�C#L�����πQ�@�i$Oж@V(�D���'�"Y(&�[W�OqLX�[�������_�uA4!G�$K6�8���s�u3�D yBx�ģ���������?1�wF�E	�b�*�X��p�H�9q
�'�TY�]�s� �j@e�5�ѸF�ԧ/|ԝQ'L.U��
��[m�VQ�B��p�.�*�_.3����V���S��5e�4�3+K�B0���Ɇ1	�Њ��Ek.p���+	a:�C`L�)�n5(0Ǖ4no����F�8�������xHm���K)l� �?Ѯ��M��k4���9�ɶj0������L����#J��]����N�-J����	�|�$�ސE�1�w��:eJ��� ���N��	��	$D6�b�GN�0��p��e�{�ja
�c��Cu��H��W�\�WM&G>�:4'��M��#����λ6���E�� �F|!4e�#�V1��^,�� F����@T.���U�I�l�X�-�		�Z���j�^.��@�&P ���0씍-�����ib��h���6t$�2 BI�ly��Q	�;J@$5;���P�dǂ)t�M]$���e���+$�"��V�F��a��X�d]؂� � `!rD�I�mȎ�\�� b�8g[Nc�(R��:bPTa�6�3R��� �J�&+¨K6��kŔ�B���hMXY�M��g�$%��*^of�)1FJ6�q�l��RD�	x�����WZ��b��eǪi�2� �)�`a��D_(X|c�웕+�$��WH��բĵcͺu��@�*�r59��<T�(�A���:b����	�(۸'��ٴT-w�"t�Ϊg���T,�MZB��'Y �:��&6٦k�
��`L����.T iz�
�C�p	9 ��X �E�$3Ӵ,S�V�jx�%�iK�((։A0T7pjG	;n���{���`�k%�G u���f��8N�$8ƹ�R��q(��&�-��A;��{������AfJU"#KG6��3����V��8ժ��T[A��9P��lDy��Ĩ)b�X�	�<f�!Il�cF�Ұ"D��	�3��v�2Fĩ)f�@�	ܢ;k�9�L�?U(/]�T8�Mi�Fӎ_ �CDʘ�7n (笤J���*5�z�B�, 3GLڸ��n�G:q��E��}8X1(a	A-u �����}T�h��#��:��Q�@	>}�w�m�� ����E($��MHIP`G&]���s��B�G0��a�x�MV�plK���+&Ș����pUHǶu%Ɓ*�  *O�j��PfU�a@A�e�I�w��I<
dXUrp�T�]�rG�ګL�dٓ�%bDI�E�I+u�����<�ᧀ9<}���v]F���Ar�0�R{�d\ �%D�
�9�G�; ,]��뇇tTV�� JJq�q�]%Y�S�@�>����D�6����	1F�dã�0YIBe���d���5�qhĸwԘɱ@� !$��J���L���̘� ��-������;~İ��iCH���t{>d"T�K�O�2)�r뙩rQ|�I�#�CG� E{"��?OB���
��}���Hї{>��qF��"���a�@0�d�Waҫi.�zbj	�/�1	t��{:�ڱ��&��҂AZ�E<�L�ס�G ���5��0h9t8��B��OvZ�H@�� �`�aa�� d�b�(p+ĵ	��K�p�4��d�	v&�PC�1մm��i�nYX!�$�?!6Z�i� ]8e��%�Dr�y����� ���N3�j���,�WC|�A��KE����G).�h�h5���� �4D��	�~��⌇ӿ�am>E����o�3vh����|լ��8=��3'��а<�H�M���S�N��C��˦�N,��l�3������G��dҁm�O�����ٙH��o�L8�� �I�."��P�PN�C��e��a\v���A��E�fa�p
��B".��/�\@�� ©Qf�%��?Cā�b�E0�"Fݳ���C�\()�Bx� �O�13 ͐�:Oҩ��-E.!��#H�^���T�ϩJ��O���EO(M��rh��=�
D�5�Z�NR�����_�#��˥n�@Ξ-���[�S�[�bH9�M;(X3e2x�	"x�\i7\�F��){f��w�T���g[&Jvt���C	2	V��h�^�q�U¤ָM:�0��ϏV��3���'N~d����	3V��̻&}JE��L7@<�h���L�A�ix�'ԕ�$PCD��>M���$��y��;���}_��	��O����GL�;p����'ŝ���q�ALx����=yQ��m����d�<�P����]H�t���.U��{�$�'>���j%�?�`\�򁋤Vʀ�&̝73���F�-�L*P�Lo�ʱ8sc0�nL���K$V̌�F�\�24��(cL��.����ƪsGi�f����R��7鉾H���iQ�ո"��|��ّ�b�<b�����
�7_@`�3�#���{�JN�+�(	z�eĶ8�4j��=f��誒� 6]�$�
c}r�U.
+�M�v�U'&�!�E���?��b[�m�X}�I�����7
�@���Ų@�F�A1ǂ+\�5`r˗�Z�&!��`���$�v�����sv�I����m��%H��� �� (�&L2�B&P)9<�����'��Tx�D�f���s��)
ֺ�*�'O:�rV�(:9����-�-�J��풠Z��\Ȁ�'�Ai�I�	2�&�u�'�>0×)ʏh��Q�q�2��ЍU�ɋde4IĤР�(�������}�bc&gYn�J$� 
�t�19_���ٳ9��H�	h����A�%��R2�b�`ŌY�2v���T�st�a F�TĈ�у��c\��1�V�v�5,X�:x���T<td����'����.Œ1a9E^(������.
����A.Đ5MQ���&�� hΟ\X8˕��7�|��U
�$:z���eD�Xt�!0��9]��e�`��TJ�U�'X�%{�O
k8P}RD�{��|��ᛳC����&C��qJ����%\�5c��
n3JI:���M��µ:@J	%TS � �d�x�����E�T�*Q�P�ֽ�w��#�%ӣ)�5]�|�Su�y��а�bX1?��A�l=T�΍����'�!�c	�7Y�n��;E��]����* ��V�4D��ȅ�	4cҮjf��!Gմ����>I�TX����hr���L�+N�dE4����`���ج҂��O�Nt�poYm|��!�M�P���)o����Ҁ�
N\P���6�K=����ǒUӶɻw��1���D�^����S蔢*rX��,�*d����"��:�P	Rb�'Ǫ�"�i�,7!�<�èU��hO>0���,�%�*�$QH|I�$��c����H�aR%�֗JO(X�L�+��T�ѧTBli���e� �+c,K�I/���v�X/n>���A�<6μ���8�O� ��Z25�hq��̫76�	�F�"
�;�)��PuƸz#��h� �02�haU�(0"�I!6��)���c��@C�EX��'�2�.�z���'A75N����Y'0�`!b�uzDa�'�p�qg�u���@��V�
r�Fp�V�)��$�0d����M>~%�؋"��o�Q�(�v�4l���p�?}"��ˢ��k�r!0#�Y)Hk&-�Qi�:"��#o�'x������R�s�b�;4�i���+ͨO쭸C�I�A�(}�v��?wFY��ƞ�:��0(dn�k����T_f�����H B�&]����}Pm�5�_�?�>�%GӬ7��}c&J�!	of�PpECQp0�F}�HY7g��&�3Q�>�~)��	q�8�I2G���S��$f�ܡ�G�iȔ4[��P�;�t�fI�t� �hޥF�ݡߚ�s��*gx�x�$
)}� E�U���	TR��"�2�Z�*�ur�ѕ��	E� �K�g�|�R��]�`�h�H1�&��K�+b��5��@�4� I���NdlH��� (n4蓯H� *�Y�d�<���O?  ��h7��Q8dz�G��c�`��p(��$H Ȕ�� �'����ᕜN�Tx�L؝ۦ�-*`����jg�'r< �ʅ|�X��ůƽH�9�JͼlϢ@�I�Y�j���D1k����VLK�y�B��Uχ?M�%��*�?j´h��鑎]��a��#Ph��R���!Q���J���OZ%�PIG�ؘ-�%%���)�y��@�D[���:��ˊ&�|4�׎
RD����+��H��G#~�� ������J� ��nV�p����5E�P�`��-Z��ɗ-�5*j�3�x�:��H��nZ�j��tGR��fU�@E.)��O�	�
p)��^�vcP�9T$R�(�@M�����u��1JGFH8�B��Dq�#�?I�L�"a#\A�
Kse����%��D0:�U�(��F
�[V��ͧa VYڂjJ�wh�����[��J:5j�}�JP���G��0�2F�V�Np���E�[�(d $�ъQafU�_�㞠(��Պ*��	bGl�(.��9�wc*/��b)��p�B���"~3���"�'��ZG��)+���C��#��`�i�!tR��5l�1 ��v��	\ӄ�Y��#"�<扞X��,s�a"o���x`!@�L\��UGؖS��e*cƁ(\2.���j�oz�U)%�ܤ6l
����ӎ�����Y�T��Ir�F@*Y;:ՠ���kr�u��!5�A���,��Feד*Q��_�l��ɷ,��|ɂ��,���m�O��X��۟�ܐ�[3�Ȝ{�HX=֜Q9剙4��������#-�S�rO۲�ƄS��9߈yiu�X�6��7-B9.p
8%曥.nP��H�=B6��b��Qg�y�r�Ę ���#��?��MR4(�4 �/�	'�Q��b��].	�)Q�8�\���k�;/.���A��o����?����B��_ c���"۩[7�A��敼i|81��C"2��,"bC�`Nճ&�ǒ �. b#H��'<�y�q��hp<`M¢2��0R��d��Ba�U�XPE�"t����G�)�%NI��'�"פ8,��	�C�7*8�e�P�V�x�:a��[�ip�T��$��Rp�؇�Rf�!�V�I+L��a5�{�>Y���Z0lz�t��D�Rt�З.C"!
t$�g)���°���^��ɥqFl;���=r�ڠ�HC�m2�g�4+�H�+�0��A�p����kͯ\��
"���B�
�Y��Y���؂a�/#�4ɕO�v�B�KǗ7�� λa��O��"�b!���d_2 2FAA�~j�M�dj�#�%����b|�c��!a�Ck7T ���-ǇFF�I� 2�N�y�o�b\(�ў`A� Sk���Oh� ���yY�y�JO!SƎU����m�����7A�� ���O�����J�xZ�I(fͶlR mM�PH��+;NZN�K�J$����^�Q��˙�L^H�C��]:W�$aܴnw�E�P�8j&��6��2����7"����Ƣ�<hft��)O�\��c[
t����1g�5@��Q��?���$���&�͠z��`��6��V�rBj޺d��:��8�Pɏ�nT-��͍�'��]�bd�ć
�6��y�Ʀ����/&�� �)ƋJ���,�*3i��r����Pb�XeVX�yS�W�U=a��)?s����	J� ��P!ά��	MR�q��sb�Ќ��V*Q_<��E��#x�@-c���`h�-O�U�,�&��1$>c��Y�X4��2ost�AbÃ���RN�F���UGր3?�(�a���L(����`�_w`	��I2~�Bg����0�N��)�>��Dܩ/f(؋yB ؍%�2�k�Aҙ3rV�;��O��y�M�
U´+��/��[3 (�y�č	پL2��@%KC��B��y�i^����,'(��%=�y
� �}��Ǵcقq��ᒗ~ҁ�b"O��x�\:P\6x�7`@6a����"O�1�C�)eؤY�/BXdM+�"O� ���)C�`1��4�p"O����A&Gm��v*ƤFP�3�"OzD�%��-�,�"�+��b�@�Sv"O��W��$��;ŬS{���cT"OL԰PG�6���ⵄ�0��1�"O��Ca�N�s?z�)�霕:*�}#�"O&9�S-��^�8��J;Dz���f"O��4�.?�0�bH��2;�"O�p�	�_004b�i�!� ��"O�lK0JA�*/,�a����{6��`"O>���ť�(��%�U.Q@��%"O��kү�9<l��̒?F&xw"O�9Х�L�6���
ӫXG���"OTT:��;$_�EЗ�S�NK.u"�"O �q�A�Spe�p'�nv!�S"O��'��:9lܼ!��%�X+�"OP][ ��[�t�7έd�6�""O|p(�A�_�@��ȹb�P��5"O�	i��U�8�R��܅�8�B�"O�|�#�$DȀ��f�P�~�2"Ormˑ��> 8Q���&��%"O�����),� ����2F5$�5"O����H��qk7H�ht� ��"O��*�Nk�ݰe)܀}cNE�"O,�˓J�j���B��EY޵P"OZppPDJ{����;(g� JP"Ora�di��G���B�n1!!"O�4��nȣ1;vx2"�&Z0q�"O`H;Q�S�4RrREX7�pj"O��� ��'{�Ѣ�B�b	TI8P"Oh�p��|�X�k� ���uR�"O�k#��~������EJʭk"O���&)�\������|;T�R"O��Ӏ�۽D���`l'��	#�"O&ء��;)f�*�� ���"O�ҳ-��12Y�dD�M�xI��"Oʥ�u��/gyD�b�-̈]Ȯ}�"OX� eF�({�Hsn�6M|��W"O��Y@�P;1�X�0��w�PA�"O���ҧʮv+��M+y���V�'����˟_;�ݢ(�&i�~�S0�Ȁ/�b%�O�-
ėX��PA%D�^��Ѓ�I�h���UgּF2PT�|��+��s5�e!����Sb��h�n�<!��G�v}{�/�;�e��fצ�XB� m���1'ݵ���s�̡I��	/od	���%{W��6"OhYu�e/.Ea��[);7�ӷ��埤A�b%.����:h�퉇Y���PT��A���{�Pc������3BK��ScaצcN��b_�>�*�ǫs<t��e���<*�����	���� aW�P0�	Y��Q��0� �6=:I�'A��F�j���~��*�z�Ҧ� '?�s�O�e�<W�[�a$4 ����hV B�pv�MY��8�mpq(K�b"���fT�@�Q����'�� ��׬��I�aMbJ�M�
�bH�A�r�ϒ)� i�#D�=�t�R�c��'�z�@RNR�f=D���c2��Ɗ'�"E}�Ǎd
�薞@F��qK�3�HO��`�C3	 �e@TkO "�����h�`0pCr��G��R����|2�)�"�ʑY$i-ғIj!��/�I;���iZJ�T�4cN2F���+0�ِc��9��DJ4O1�,{�+[9��)yɛB�@o�~�* $�5��
#�N\����Hn˓(�L"A�«*-nҧ(��� �@	�u����UǦ;��ȍp��G�J�H(Z�`��"��I�[�uq�� `��+����dJ�H��" 6����<)始��&L�G���4.4`����#z!�آ���m�dA�+��Q'�H�K��`�����p@I��4־��Q(&�ɵ.on �q#yƮ1��mS� Tr�:�X$�,Ш7lڳ|��	1M�y���7b�M�C�
�B��0@�y��o9� ���#U9ub���$2k�9[7n]0>8T�[f�. MXL�'���`N��t�� Ya�LZ����8%d��QUM�7M�
�"�Րm~X�k�fؙS�Q�dM� `\��GU�&c��i5�ѶL���3P ()��y��B�e��s��U�<��h��8"`T6�2u�P�8��>�Q���|Ƅ���
d>Q
�h �S�rA�S�Gz`!�犉� �4�@ѫ�(�3TW |���R�"�.�>Awp��JI$"�(�r΀+��1N6�.��m�!(!��	�v�D���OѴ=�BB�@y2�B�MD(i�&h�<3R�`�W�;2��p&�i���a����f6@�y mU�<�~��E`\.%qlt#���Ц��G��l�w]�_��Mc7�J'��ƅ�,�[��˓U�Ҥ�R�;=�t)˶�����*�\�����)C������.�@��"+�َ���
k��@�"�ğ/�@髀-(G�ൈV+�Ħ���5���؈��P��Ab+<�x�e�΅��J	�% `H��dY`8�)��<�T��M�L�d� ���2��KV���!N�H�L(���و��M�X�䌁���z`A_ͼ�Si*q�H���+b���
�Ř��?-�.m�*�B�
J�4]�ՐK>I��ʪ0T������(rH��U�	�}I�������<53 �:]������ (^�5JA�1wX��-OzQ���N��1(Nͣ2��I��S�8L$� '��p��(
C�>�dEr�� R�,�.�&ɳ��cxF@X�� 4�L���!ȰX���h�c�Vc�iY����/����:?��j��W:8q��_�Nxb>e��@�\5>HH7mW,t`�ԙ�e�+�0��CBr�l��N�-R�T�B�	�Y=.��m�n��7���C3;\�9�K�p�"1�r�A�Kh<0��e�"L�11G��+v���O�s��
�D8��2�lD;%M����ɳ3!�p �c�N�R��\B��F?��j��#@��54O~l"b �mN���+��5F��b�V�lc�%V�Z�޹�V{ܓz��I��\���(�M�"��S�	�f��f��>L�"�{���;	��
fon����"�Io����mB;:�nU�Cf���a�%�A�Y���� զ�	��S�7>��%���?�| "��[R�0����6x���a�P-{2��A�-���n}�����Z���I��iY!�8��A|��yW� 	W�9�M�d��x1GʛqhB5��e�%� �y&��{��i��	U��ɬK�<��&O�fc$a�E^�xN!�$�J�1�P�Id5 ��Y1=x���,U0�J�d���5�c F�B�Aa�(Aph
���~��2j�%X�
�S����bQ��p=��k dap�Ԫ^8ð�z��~L*Ф�0:Bh8��.3#�=���N��!���t��*�?���p%�0`��ЛA���BR@��<�a@�*AZR͋p�K,^�%S��O>	j�jT�T<	����h3oĸ3p��6z���ƿX�(��K���>�B˩j�3�L�j����i�=J"���v�P;�t@��*��x��B��o�c1�i�B�#ϓ��yG@�-Mʄ�v古lc��Z�E��y2��,_�d*%a�8g54U�*�۞���&Q�Kf��:�l0�0���/W�HB��O:b=:I�s*F�ъ6�ע[�l���sPDr��O?�azb��� 6��"��~��:em��p�6e�1A�q� >״(
 A��e[8}@Ӥ�;`-��M
#f"=	�
�ʠ�ThL�P�n�X1IVV̓Q�d��)F��� ѬM��0aՊ��tMQ���(��L[+Rn��͘b`�������
� �,�����)4j��.��h�TDZ�e�P��Mɧq��(0#�@5LM��1���ݞ`Z7M�4�d�4D[`�h�A�Ȥt��< 3I�4HD��ID�F9g����ڋ��k&{�t�9Ѧ��;6�5{g�t�Zh�P�3l��S�Y��@SSA�;ذ���}�r�╩̷2��c @O����)֪Y��\�9
Ę�M�x�h���4]�@�c�V�&�(�x��3,3���%�� >�b�@,B
%i(�B�O�_�F�[w$���"i�e,J�8�x�+ȁ���y�O��>ƅ�!j��\�!��%��c]�`p�q�����UDybI� z���jr�ނ\$��uJ-*���W�X,'S�5�ɐY��в��!{���rR��[)�(Ʌj�?�[C�Dv��	����еi��5+$� �'��*�2�<��C�����5i��1#4�@4&W {�z��cFN!}]�i����+!nt	�w����K�(��d�ͮ��[w}�˂��=/�TY��@�(�V�O/�f��4�؁h�l�$��"G������%U�&u�����-w��5k�m\�U@�RMB�2�`�c/�cSNe �'�.D��j�:���f%�by@�j$��$1�j��SOMbQLmƇ�G�ҡ�;yБ;�ܽT��m;f�Z�G,(�Sg:f���u���f�jt��8|؉��ݿP��q!��5v�Y�壀#[�9^�9f��x3D���E�?0�E�#�b�pe�g��}\�#=��H��LHs1 �+~�"5�3�ђ}������D�	0���j��?�%�'�.�Z|���)z�$%nZ#$�@�5Z�{
9��j��~{NI �Ƈ%|V�@���Z�ў�B JߜV����i�S2
�YイR��C1�P��R�s���O7(HJ�M�?�O���xp�d�¤S��<#ѣр�^�;`�	�zt���j�uXЉ�*��D."o8�'R<z�ɝ�B�j���̀0 =�7D�R��	d��?����_5rȼ�B���3sXH�J���M�VNY�VF���	�
X	�IT<o�eS5�
m�0�&�IW�W�_4�\S≏?��R��Ýr�`��7 ��`�C!Y+5�6�a'�֡Y9�h3B��?���� ҆xȐc�J�*�0��/XL>Xr���	5�1ɴ��2�z��I
zt@��iEH�z&�^%�LAt�F�i�R�)�!��g��i"�ԧG{xT�F)�V�j&�~Ө��(�
�������o���Q�țB4p�v�'���!�əF<@��'��]fv ��8a��@g��;?<X	 �&�w+֭ۑFwㄵ���Հ3op%xW]�h".:;5L%`3f� s-D\Xw`Q����5Ǖ��v1�|"�U��z	��rիቊ?XvP��A�A]LH`��E#�t��Z�`��I�f(^�7h^8n�n��D� ��Oͫ��͉C40�&)��c��9a�^"@,��͎�&*�4��#�b$@�W��I��M;���Q"B"�PU͏%,�<�3�o�A{�ςl�(,!2�L3Y}�`H���4V��0���&��$���'�Vر�G�3�Jl�3
Z&6Ү���(ŝK|� #�E�?��Yj��z�Pԡ�'�0�ZH�Ê{ӢM�'Gn9[��Ld$h2��^��\z�&���+$t@`!s���C��M��'Vאd�� H~�4`�߄;|`7��L���-���@Ǐ,)�)���	��u�r� �y#���I^:��2_�,��< a�I	"̶�뷣�%.1�����N�g�LH� �1\0Ѣ��$�ǆHF
�pS�Ձ-�D)���{o�lp��·�:��>1�aЈq�u��,Q�|,��bٟ�7�ܗ���O6
�4qX<�F���8a�ƦuzRμ\V������I�jM�$����5%ɾ(:���@���xZ�I�'����M�+�l4��Oѓ�\���B�R	F!~����T�$���	�-ď)�b(�����ZEQ�JX2dMR�)]� ����e�&&9{!fХ������9ʡ�t�,7�I	�K�!7v�£��On��a�6�T:�,8ƽ�ԡ�5�M9�K�:�n�0o �$)�:>,�i]�|"�Τw|@`V,ۉ6ot��s�_�(H�(Ѡ�ް{�旿:�J���
�d�9jQH92elٓ��
[�"D���!�̘+��Eg�0�!�ÂN��`�BЧո�Gyr�ۺF`�ɡ�J��e"Q�Ҵ�CD��ڒtr�B>*�-s��Kb��,cP�H'<>���3C���A�m�0ӆXx���^�}��H��I	$N͒���a������,�&��h�t�*n�mh�_~��D�I��K����faƦ���$�|ybQFL�04�YC�ԫ_�:u�a���`�<��	^ U��*ъb%P�C���!�>��Ţ��,��x���84�8��[,a�2J�`#@�Ӄ�%�*�![��GJȌW�, �	�-G:��$�!L�Eaa�+n��Z�o0O�&p{����
���.�(D�����7 Z!;q@�.嬹T]�I�0X;� T1��J`��O�n�X�
��ؗ(�}���	6.{��ū�N� ��^2)^�Y�bGۢ]���;%�PT�ᄧ�=�9���>T��X�aDKt�����v��s���@�'�P5�⊹{��y؁�̻f:��{�nM(����N��ܜ;��<q�D�T��8x��U�Q(�c2��+�K?"�Z$�R"lؕ�p��3ªZ�M� �o�Fx��Q�f"j���3A�'j��g�N�0`���)��9�m��A�~�Cf] h����X�m�8���o��+b��=~��L��9BGh�C,�O�BfDh�=aw(�4��p�3H�+�"�J��ŋ<Q*Y����@���p�`�v�^y�3�҅]t�(!�k��sP�GNtB��ݐ=�|���=ʓ 9֙KІCFTz�ݒ9�l�X ��c�y"��C*m/��1զ�� �"=��X�G�*��V���Va�A@�꒲b�Yjt��%9��L-z�lc���Z�V���Ҝw`���SK�%ٰU�e��^�<�9�F�	?�L+B��&^�@ٸŊ�rd�A�,�<ig��R5n����*�u�v�G}b&ۑ@�"Q'��A�M|�< iń�v�,��`�@i�<�W�BPA>�q'lӒ��)�Ly�6Q�Ût�&�q`m��
��ɸ��YI�� '�PX�'}�B� M"���!?��XH"�G-A�����H�}Vp��C��$ݪ�;1���G����'嗫;��	rM�:�A4�ɼx_d��-!����<��f���X@���<4P�NN���$�gN4(؀��;8(�1&��!,Je F��
F��s X�M�!sW
�Y�܉y�mI�g��)�4��3s�D��E�ܚ3؜�i�*9�V˒e���1F��<���X`H}@V�HR,�[4l̢{H��ȇ��b���qu��3C���7���}eF]�I	�T'�,ct(���x�w��l��pHF��9T�����w�' �%�V��5x�p�����G���1�Ef�X� ��i� i�,ъ�l�\ԾD���2z�l�&N�,Yɐ��UmK�Z����Gm�4��;U3>-AfΏ6��!K�G�^]�!�'p�ye�;8�Ԫ������v�inP�KΟP���$���l`��VfA���;.���0�X�ĸ�嗦J'B����vT�/\pu���9*������"�l��ꆛ0F��j�"�2���@BX�j�c�\/S$HKc9��`����5N��z�b��0���"�"�.%�����	�JQ��[��ͺH�T�2��5=�������!1ʌ�į,!���l���x2YR�E+.|f|�aG@./'D�+w���cTБڂGF6rԊ��źt&Mj��\*+rtT�g��)+Z�[׀�$g
=r��Zi&�!�@��q�I�Q�cҠA�FB?��!b׮a�����~P#'�pֆ�e���1c�1 �5rb&��q���UJ��I���1 �\Y+k��@�d�4j�%P-�7vj6��1c:t�,��%G P�|�G���$->�B�@=�4��e;w\]�#��B 8l�'-��)���G�	>dD�"B��Y!�J֢�d�PC��7'$1D�_՟4���
8nT)�"S G��}a��#�M��L�?Y�2��� <���34�\�O�t�%��I�0$��[�E����O~\bD�z��=��.W�`��YH��]�
J�[r�;"�x�	e�s�] �8#�"�sb�W yp�!��'
$iX�!��j
%� ��*T�������5�6�IP�Q�	g�Z�̍4���Rd� �A*W�����#H�6�>�1B1��H�/��"����W��I�-���q�2�k8�	8x�ɵ�E�^WX�Pr�A$uj��g�����$���J ��PQ�"~��Eb���(m�D���Z�oߦ�� ��5N��HQ��"��A�&i�k�����Mכ~	F�GFy�7_jB�)$�X�E2D��(z}�H�U�E�CF�˧��3�Z�X����W�ہ)"u���^#<����)_=~�5`��҆�S�x��Y�F�ĊI�n¸;��E�Q��)���C�I�T�,���
���8�*�.P;��,He."���>�0`ENB�:�rI{�AL�'\d��Ŝ)�V�1��W�u��H��A$� *�F�q ״w�"<��C(XF�%�z|hڕ�P� �j��e�+aRm���$Y�R����)[@��'9 ź�hPF��X�bjOvk�� ���Y
��ӡL�XY�f��q��#=Q��N,^6��
I�xw�L�RP�-��/�p�Z�mޜ11جc��>���yq��H�.Ua
��k�\�l�E��������<^
�`�ݱm\��Ҏ�D��xO��% ��u���Ο��h"$ָV:H aV,�?fƞ�Q'�ɍ'@d�s��g�$�{V�ɝu�Q?����G�� �rL�C���a�B�B��$�jdp
�L�IT�ç�>�V��$}Q�K7וa��]ҩO&훢�:q��5��N�'��(���L2)ƚH�Џվ"��q���By2�?T���Z�!/��D�zf��h��]RZ�X�'�4;�� J�{e��"Ə�+.�D�d�ę*E�Ԑ����!`�̆�ɮH�x�˰Lȁb5���eMD&L�����2 �Ѡ�y
� �9�FN�+��ݰi��J#�=�"O��
�.�	�bl2��ëE�Z	�"O�� E�Q�]��B� M���"O�=J��è-z�d{�i�e,<١"O)�P �,�`�8f��8�z9!"O��s5n\� ��E����;8s��"Ov��E@�$�0$��ol�B�"O���@�f�b�C��ڗ��Aq'"OzaS� D�N�̉Ҷ�D����s�"O�h8 C]�p�ϖ%��Ay�"Of���B�A������EpD�JB"Ov���yAt0�4I�6ih�P"O���eڠnX��z��#]"%Ѓ"O^A$K�0xr��5�pӞ�b"O�q�-Juݦi0���y�>%�'"Oa�!c�����Ԫ�]��� �"On)�"+�M�԰p��9�(�"O>���3�h�0�e�K> ��a"O4�2biٻ)�@��<xr�Ȗ"O��(�NW�+��̓7�֏*	F]��"O���,�W�Xy27� *-`l��"O�	p�Go��=�@�>m�j�"O�q9Q�D����#���9�"O��p�j����) C��.|����"O�$�����*L@@h	��0����"O���bI#��
��Ȝ`-����1O��I�+*7���q&�[������I);*&J��:ڠ�+� �
�����BR d�bT��-J;B�
d�0�?��U�ρ�&yiG��@0�p�5��a� �6p��ٴf���i��F�l-X�*�$�:�)q��~R�a��u��MZش3$Q�o*��8�g!X�M�f$ ��Ɉ0^2)@��k�`є�i�=�����2�<�[F��:)Rތ� 3F�T)۴�ا���$Ι���:a\0d��T(-���'�H��1O���7��0|*�iU��z�2e��r�^!�L�E�D��[侹J��iD&OK@�K0i�;>d*@�ib�DI2��Q ԠS �I#��4�0����#6�2s��B�Hk@/S!)z�}8r���3VL�O�O���ưi���X i`�D���(�4
�y �C,�
y�e���<E�$Ĝ�]�>�t���I�@Y�@C@�Cέ�u������ 8 a�t��t��"5-/�I��*ϐ�I�Z_�-���!a��K��/E{�n�'Q ̛$����;i�Z@� O��<�ٴ��>�3ĬE�J2Xh��E�Wg��1��OXТT�fXZ0�>E��KӞ\8j����Z ����?�p��#_�OQ?=z2�B^>������/|����#'�*0̓j/����'Q�g~�-�� �� 7�����׽3R���M P{�'f��)��@�6�k��E����pQh�>1$�OrU`O�t�j��Q^�I�4X,y�Ttr���<镮��̋L<E�$��)X) P�P��=��p�!��0l�n�nZ�J1Oa�D̂�0���v��@�Di��l�.� �y��O�?�A2!ʡCx�m�U��8|�� .�I(�?�� �<����=�"��L;���BB�N��<O����.%�)ҧ{�-���Ȫ!��]!E���nz~� &���Kn��
��)B�BJ3cV��#��\6���m�I12O؂T���'�T,.(�ȓT?r��թ�!Oٶ��gT�d%�9��a��i�dN¢2�2(H���UBNх�PY<z aV!2�DTrS#��&���$5�Eb��T�+vN�bcJ���%�ȓl�4ʕD���k����Vm�(��9<0�h�
`��h#��5PB���giƊŭ~8 [�\`��H��oD�h�d�=,�"�
�xD�ȓ/P�����=���aEQ����ȓ�P:M�y�L|�f�1B��݆ȓ��#�D6z�tI٢F$���ȓ�@i��D+N.Q�cCI�&�Y��S�? �����:_o���j��+���:�"O@L��e�(sՔ�C +j����"O8`�Q�L��H��oF�/N�k�"OD��"�8�L*S��;N=�-�"O@�17j��w�.t:�- 9H��S�"OҔ"qjH[B�t��l�&uEa�'"O����Cт`e(�8�ꘈ#AL�[1"O�yǋZ�h$ѳ�� 
,����'�
�B3_	}�L�EW�b�
#	�'�����x�(	q�憈`����'�*(����n���I%b�c:h��'RX� ����H�r$�3���<���'�>L�P�j��P���uB�	,�-���L� ���_�h��C�ɀw�I�go�7�$*1�\1K�B�	�(��X�SE	c���� ۂ�B�	�0@�0�vnҔl��#%K�B��= O| 2�Z%k��E圳M&C�I>k�)�pb�g���̐�5�B�I�l� �[S��.8O�hz5ț�Q��C��#�P��T���a � C�nC�ɤ+�ԋ�[)qֲ�f�֝FLDC�IsG�h��O	l`L����QC�I��$!�(���Fl�b�D�&C��R�)A�"Dʩ�4@P8t��C�	~�"@D�*D���"�:��C䉶K�FՓ%-��v Ѣ,�I|C䉭%���`�ĞP�t�1��^g�C�	^3��Q�KG�*�ɚf4xC�#B��9S���`i����?JS.B�	�V��� �&
�9�Nu��n�	),<C�I�<�ЇĎ��0�o��s|B�I.;<ı��+�.Q�u�R�4�bB�I&Pl8u;�L�>w�2]j0�Ζm,0B�IX����v菿	=Rc.X79B�	�wC^lq��@�l�����f�VB�I �����N�����F:B��\F��t�E�Y�(��� ��T��B�ɿ �hj4��;79>Ԣ��4p}�B�*̭q֏�v(�P��ԀwbB��!�R��+I�#��x�KS�*8B�I� ����oU���������5q�B䉌'�
�-y��țS����B�I�g�8�CC/u� 8Ee�I��B�I	h¡Q�)� ���'	c(C�ɒ��h�kEd0��U�}e����']��� �o�d�8��� P|���'�Z�Q¡_uT��cZ1*K
9��'J$(Bb�G�����N�U���8�'��fn��,Ϧ%��j���p��'���	1��M:	�W�-q�x�'Y	�j�D��q���S� 8��'���p��`��� �`��Mж�H�'�.��v�KQ����X�Ibd��
�'������I~�� �틌E��Y�'��A���� [.����I��P�R��ȓ'�&�$�J�K����q^@�-�ȓ���2+H�,{n���!A�rd�ȓ)n|�1Wĝ��P󋁰@��M��{}�:��΄��!��)(>,��g;�yС�2Y8"��VP��.0LI�3LD�#T��+���,�ȓ4�@EU�U�� ��$>�ĭ��5d��@�X��ܒ#��
,����S�? �I��nE�_�t��	U2S���5"O��+V�җT�4�!�{ת�!"O�<�枙{¦���]�QՒ���"O���h
OQ������}�"O����ɟVK�$z B�0d@a��"O���5��:ᰔ�� GrF�)�"O��C�@];��#��H�J�jC"O�@��a��@��E8|��,�$"O��jC�Ŝ]pp�q枫d��-�"O�śB�.��0b+��b�d8!""O갡�A����@�;��сE"O��y�㆟L���s�2����f�<����&q"��[���7vT�)kVm�<���pr�w�xJ�q�l�h�<��Bƛh:���@�2W}���DVd�<�ǌ�/J*��T-Kl�t�z�<ID� jQxVe$Ð)P�j�s�<1֯�r��Тu���1m��S�gl�<y B�	7,��Zf�	�g���@w��s�<��ģ�JX
��G�N(�Hfg�n�<�u�Xx-���� �8��H���`�<�6�I9�
Hh�iA	U���棙Q�<�ca�)q$Z, ��T'�$�$�M�<0i��<vʬʑ�� �ĉ+��M�<J��g�b�_�@S� QA�<�#e�'
ޘm��Y+�ݑ���y2��>�h��	�W_���Ca��yr/�1H��d���MhC�oY��y�cLZU�`���	��܋�B[��yB#V�na��2C�r|�9B����Py�d�; R�� c�.*�8y8�VS�<!��_�~h��I^,\y�E��ȖW�<�@���(�)�`�s�:�SV�HU�<ф$&~����@�'�H�;UOj�<��nPzH!�I��xVд�`j�A�<"
O��LФ�̢�A�M�{�<1��E�0��qWϟ�/���i �Tl�<YceʽU ���ʮo�
�	�i�i�<a�(TP�~��M�\a��q���k�<��.B�A�Ry�S勦%� }�QLNk�<�c��Y����N&�p��J�[�<���ǗZ�2�+R��#SX|r6��X�<q�F�<�A@�`b�NZ�<�P��P	J�j
EO�$�T-Y�<Q�e� 2�¼{a�W�.>ȍ�ģ[O�<� �̚Q*��Ԃ5�Qqt�S�<`a3EȠ̘B�B0ʹ�AP�<���j�.%�$�2�n0��FO�<ِ"F;�0���O>k� Q�c��K�<q��R�~Μ8�!��dq0h�mXI�<�4��>�@�Ҁ%ӏ/ ���EC�<1Tj�"���G�h��Q$~�<��O�'4��M�WgDt�0-/Q��B�I�İ���r����.-a�B�	�5jr8���Y$^�!�g�.c��B�	�>P��;�Ǔ9]���ӍK:`hFB�	��`��0�Y	b�6B�?H��C�I9<r��և�/0p�U�G/�,��C�	, ��t���c4��$�ʘ�XB�	�&Ʀ% �H[N�T�#�%\PB�ɂCʪE�Tg4\��cďI�pVB�ɽ$�ܥ tÛ!0��a��m:X��C�	!n�ų��& �f�	�'�2R��C䉊+�Q`4��ZO ��I�zVC�)� `H���!T�� M�9���"O� �5㈆of�E��kʭG-��{�"O<Z���$~�9�W�9$)е��"Of�2�F_ �Ba�C�X�<¶"O��r�Z�a��5�=�x�{R"O��f��4[{ڀ�p�
a6��e"O ���&�c �ے> 8��"O�����#2f�!D&S0u��"O����@�1��  	�19e"Oz�8��]�����Ř)�(4�U"O������V� St��9�"O�t)�Ƙ�Lt9�&�P�J�:�ѡ"Ox�rgD8q\hܩ&��y:x%0g"OV�XbL�rN��ҵ�St����q"O�ԫu-�P$R���F]�R��$"O�a� ̚oKX�JĮ�>d���pg"O��z$l���F�`�N��ZZE"O �R(C�x���(M���I�"OX��V�&/h����>!"���"O����y{rD���
 ��Z"O�ȲFoĪn$��@U��>F�0,��"O^@�i��~2p֋qgB	��"O�5�bcáGbB
�,��j0@)8�"On�rD+Zt�(�4i^`}�%�"O�@JԄ�2��k��1m�T��"O<HSI�@@ě��d��5"O2lB%`>qP���A�abȳ�"O��Ѩ���T�Q�٦�4Y1W"O>æ��k�ꭡ1o���<��"O�AK�̎�t�4�NH�F�#�"O�@��R�0Vl��cC�$��	�"O�LR���*{zbr��sf�iZ"O��H��TEq��U�_fx��R"O�)"$��}����Iߚf�r�"O����kpa�Rƀ�(p�p�B"O���6��BBj��ń#
Ii�"O�e@-$z���2 &�Lm��"O��[�?̈Q���72�($��"OzA���̽�bݲð���"O��b�˥]�e�3'۷�"���"O.�[�FȠA'6�x0&;L�"Kp"O��V��'$e�1K[)K��	��"Ot�
�o�V��U�0�V�9�j�YC"OFy�DG9wS�t� cU������"O<[�JX=i�h�f�w�P+ *O9�c��+O�HXacHT9DG���'�bY!S��	�b��h��`q��'��M� qsE7n��Y�'�p����Z��5����(r��Z�'s̑PD#աZ��$f�����'I�)3d
�&s�t*F��\���2�'���k�J�& KNU�Ek�Y1���'F��x�B�3�n�e�!eV��'�a�5LM�%�F�juϙ�i�Lu�'��&�.�D=��� ;
���0	�'�Q   ��P   �
  �  9  �!  �(  �1  -8  o>  �D  �J  HR  Y  __  �e  �k  +r  ux  �~  �   `� u�	����Zv)C�'ll\�0"Ez+�'M�Dl�Dpw:O�1"�'"d�?Y|��̛'"����E�;Bc�T�`��>DK���(R�9O %r�%e�i��#�?U2���?���%�f�:0������R�#���(:�\٥�HC��h#B$9ؘ��ǖ��u���!����'�M��	q����rj�7y`�1ud�$L�jq����O��h�ϐ�,���9�@I���
���(����<�����k��P�Q�C�Wp�i��"Y��@����h���fyB�'z�q��O���'S�Pi&�ؗ~�0)��I�#���@��'���'-bY�L�I$C����h�����|@j9K� or�){��!��)��	�<ywIɏ({�upd�˶w��y�rJCA}"?O��O|�	�.�>�u�?���+�2��@0AJ�"�j\� ��O����O���OR���O��$�|�wG����I6z��XWAG� ����1Gb)bt�'��i[T�iR&wݙYÏ��u�#Gs?�6����q0�m´b媵�`M5����iU�
��>��1�@��is5H
1G�b<8�-�!r����kۋS���8�+Oæe+ܴ[o���O1�	"n���c܊{���`�-H%Ct+W oI�7-ҏ�j�Q�O�"a��]R�-T3�r������t,n�)�MK��i�n���#�#ɞ�Ps��������R2���527m	㦝q�4.u1��ĚkDJؘEמQvĠC�_KؐsFBH>TI�u0C�=�����9w���q�i��7m���h���!U�񱴌�##<��+��i�܀�Э˞���9B`��I�OF8b�gc�ܪdR�`���O���HC�-cV9;�Gh�n�������?���?�rO��؛F�?����:ؾ@��� �J��q��OB��?a�����C�������������U�i����@d��abJi�i><��;��'P����p�y�G��u�¯ڬ-�8��2�B�K9N��!+X;�0<1�	���8�I,��DO^輁cv�����j�a�	s��'����io�ē'TG��mBh�[F$K.�O�o�6��pH%dA�8�z9�c�8��lY�4��$a��ulZ)Jo��	X��MR�3W�$�ʸв��w���.x} �-�9L�'�|-���'��	�\���kH��ن�D�Uy��jbÔ�$?���.\h��K1G ��B(ħ�h��u��%�!�%#�
�Y�R����RF��O��n����O��4?�̔�tH��|砽*cl��nb��#�'���'%�I��~E�傃{�@�� Y;80F�=�� .�	Wy�?��b2`H�t�iy&��67!.=t�'�x����D��Q��I���N�h��8�$�#1�.D��'K&^�'�@f��;��(D��1�"�--��I{1*-RO����l(D��#!H��fY�,َ<t�k��9D���c��z[(ـ���4Ր9y�k6D�p�����k�#eĬ#E�<Y�CF\8�QB�DU�l{Vb��)T�0��7D� [扉:5ø�5��{NVT`�)D� ��dJd��J�n�x�|"q�%D�LY���$f�*��'��F���)D��*��&�p��)��UKL�)(<O<[!�����I�����k-t��,c��&g4�Y����۟��ɦK�@]��Ɵ8�I-R���Y���ң/ח0�7��,#P"�H�x�����	�0<���	%���sU�إi�N�P��Ɇ�|��sJ_�!��2%�;@�����S�V�$�OL nϟ��a�kJક�қ9��+�Sy��'L�OQ>���#@>i��g��i8�}aF#&��T}B��2�M���[���!JY��@5
��(�6�|k�7Q��;����X5�V�Rb�ks�ڦxˆH�q�"D�@i�*H6���1��)�"���L<D�,X�HS=?<��p��I˦����6D�$��hD��>Ո3"]9sL�B�3D�Db���Q��1q��ߴ(k��k�/D��0''�[<��p��t��)�4 ɦ&���A���?�vӈ��O�˓@Vh��`�-}�,J�G]H��hp�z�Vis��5����IZʧ}��O�q�⠉�m�Dx���+�ԁ�2d*k�0�%�ʿX?��R1�]%%1��t[B	�~�A�yhB̀u��/�z��2Ő�H�H�<��D����|�I����I452�Qc�p�R����͙|���&��'Kf��G�K}�F�0�ˑ�#��)O
�nZ*�M#J>ͧ��+O�t;��A[4H!�6��=X�,2w�@� ��({B#�O�$�O*�� ٺ+��?	�OVDDR�~�F!ѷ蔺y�Mʕͅ'�(@�dk�O���'���wƗ���go�7�b�(�* 9��xBώ�B����'��p����2�R��ь�:k��aF%�?���?��2��KNԺ"$�&@3�X�C�=�]�5@�:ivtB���hA
�O��m�H�'d���l�~��Q	<���v^�]��	�4y�q���?!B��5�?�����/[��sʍ
��u�_��� �ؑI�-W֦�s��:1h�%�ALP�'��i�ū<���h@���P�B<���Յ7�-J�ǟ%[}�5s"c�2C��#?��l�8��M~���!)F�;�K��W�tcblG����0>i�b[�^(TUڗ,*;�H�r�\M��(����!:�.��s�����>4�Ivy��I�6�8�I�|
��D|��A	��x&�[�N!���Q���?	��L�6:����jӂeb����������O$7�����΀�Z! ��6��,�tڎ���K*9�#~�cE�$L���+�8�V���N�e~��W��?��]���&?ΓB���!Ors�1Cwf -UlT��ٟx�I������-�2Y 5��6��!�i�Ui�?1��S!wx.k|�5{�mV#R~^,���L妩��͟����K�]"��ڟ�����8��ʿ��.�Q�q
%/&
pC/�V̓I����ɒxw^���N�?<}�E���_�d���٠F4��	n�rIh6-*�3�	qZ����#�E�����.T- {8�%�ܹ���Ohb>c��H�T�y���W���aYR��Q$&D�@R��)
�,c�g̅4@.�F�O|�$M���$�|"
��9��xY��'r������!��کE��'�"�'���]�0���|*�B�)4�L���Y�u��L�w�X+0&v�#��ЪO�OQ��p=���/���Glƺ&�e���_'k��+�O���TE0\Oh�
�����
ѓs�ё	6��i���;gB�p�J9n�L��Y���Ȫ#o�Сj��))�Ѻf"OfȘ5��"kk��ϝ�Ub	���|��>�)O>�aG'Ħy��Οxz��)�vu��H�Wn��2��K �I�|�t��꟤ͧ
��	G�[�$�y�� �6.TtX��"$,��	�JjX#<a�B�p��=��� �Q��A
a���7/�O8I$��`�W�H��լag���f2D��Tf��$i24�0hӲe���Kql1�O�8�I0:���HRhֆf"qi���p���O���YǦ��	��H�O�$Y�u�'�؋�OZ�|}���R��D���@�'��fT[�l�I[�L��br��r���j`�ʊ82N �!'?�'E�/���d��L������ [��9�q�D�M���@��#sV�	�,���٦����D�OO�)Ι?�&]��EF�pI��� �8Y�y�'�b��8RmA{{���VaP5\P���8��?�gX��'��I���e0d���Sb�QQ�k@�7��O&���ON�� i�\6����O���O�(tK|��^1:��|��1C7`�6~�>�nfz-p3D�]��8�	�G��v��6��UkW,��g�x\0r�Y&V�Z���k��v��p�+�%E�0�^ˈ��fk����5�=��}�ɡ�M���Z��a�������$�O�Ȃ���Ij���2��o�,Xr$��hOT���f׆D�Vإ�$@_"���$�O���'��	Z���'�剰(.����R�P��;v���: \0�B�0�,��	���	���
^wn�'��,	�u�8�ZccR�>���C$	�(���
�'N�EY���1%����$F�/'Z�@�5~��y`@�mڤh�l�}p���(��7�:?3�4�`R�x�'��<~��Sˌ�V\�\��s���' 6�O���?���`��`^��Q@O��qpV�n�B�	՟�Ig̓3��8����C�Qy�ᕰ��'k�
jӆ�d�<q�4UQ���'~�$%>11��)���L��
�:�R�4�	� �	i�r�{�g�:"�z4�A��<q�ֆc�P�"3NNO�T
�i[�P����a6(8 �^�y�扺vCм��L�Yu�4��,R�[�����
r�i� ���O�dpW����[�]8h@��XF!�Op���O����OΒ��c�D9�.8_��P��k[/P*�{��&�O�����&��`�����Ԥ��2���<a5�Jz���'I�]>uB��Qş���
,�\�1΅�+`��u�PßD�IE��d�dV����O�ʧ��	Zd�8y�Ϫ;g6���Ʌ!`R�u�bvkW�v�|�i��S=YYB`Ifa"��o�D#��!�&-x�	�@���C+Bu��=�M#��i{��S; �`�+�4D�̴e��=V�ГO����Oܣ=��=_��_2mUP�f G>:�*D�~��xo�A�ɇ9x��0� �.|jTfK�%<D��s\���?A�g�'�
2`/k#�}�DȊ�{P���'��'���z�$�'���'��sю�<f<�3��vș�'M�P�DЭ2w�y#��7���a�'p%6D��"����#	<k��B�'�� �W)4�^1�ߐDC��9sP�\�e.�O-����;{L���C)�@��"O� ��Ʀݏ0�b��J�a�"O��C���+*u	«D�51�"Op�P���%�ʍ0 �.V��i�"O��A��-H.�|!�Q8X�]�5�'�*�'�D�"�I�K�$�q6�=g�N�	�'��@��S � ���BUg0`�	�'��E�v@ ��c��c����	�'�0����2	��xeΞN?l48	�'�H�gh_�D���@jC�ȡ
�'I|�Ӥm�j>�1:
-��P����� Q?e�f&�=X�-Q��\�q[&��3�.D�����7[��[�j]��p D��1��A�tuB�X�ҍ���+D�THf��?��e��`T�]h �+D�LRG�>�H8j��W�[n�	 C�'D��"�iӕo,"}`Dm�oX9�D`�OȠ1�)�MRT���S6j �h��AG�H�DE��'�E��Gр
X��*�c��6�D ��'���@��`�"i��� ",,��'��a�B:.jj�U�7�\��'��x� �[����m��s�Z�Z�'�좐�M�
V)�篛+}�8	�(Oԥ�R�'��l1�ᎫN3��.�G����'���Wa�ed��'�J#Pc|�`�'�����o�.'n(�V�� GT&��
�'��@
�d�q��2ê"H 
�'�l�qb�F58gt53�&��ڑ�	�q$l��:��H0РUSQ���1K~�NM�ȓ~y̴ u�۷P+T���y����ȓC�^1B!�D�9HȔ�ی@}� �ȓ
L!92Hp�L�卓�g�8 �ȓD�ԄxDK�Hk�(�T�X0Z��x�ȓ��*4�uLE�ҡO�~P�)G{R�
������`K�(�ؘ� o(G��TS�"Ol�5�P5OY��q4�֞XvjMJ�"O赡�Q�q��ȣ���*D��m D�8��W�w��)Hd"׳U�,�:6 D��؅b�v�
icv�-��X�k#D��Q&��qcP�'H�[��4��n�O� ���)�'_�)�nʵ4Xb +&�26Қ��'���
��R9xn	C�N�3�|T��'�p���d�R����'�!�`T��'fB�r�%�rGNm@BͧO}����'�,��ɡfT��;�Õ�Y�:�'�­��
 o��}[V%�V��/OB��'� ��b�pf���PD��|S�s�'沄����>)MZ �׼r�̑x�'�h�/S&������r�z�b�'	49"S�^� <yu���c� h1�'�*A3�
�;cx���-Q\�؉C�#a&t��1�DSg��8x`"i{���+x��5�ȓ\�����\�s��Gߤl��_x1�%��&n�q��$ǖ^�޸��#��k0��F�N�4�i��ѣ�'KD�� �ѭeC�4zLeɱ��u�<�fY�/Cr]� ��_����u�')~T�����5w������n��(#�m��u�!򄖻6���A�$ �3A��+A�}�!�$�z�(� .֩U0YB����!�M�P��� G+OPUjPː�E�!��Ր�T� G"�܅k�i��|t!�B1��UC-?�� !đZ�$�:�O?��@0BRn����0Cq� ��@�<1�OΞ�2 �T)|#��Д$�x�<� "�V���0���h�3�*M��"OJ��㇋3n݀]I�,W`~xxj0"Oɘ!h��o��� ��L*IvZX��"Onp�wI��:0�U(�bN�d�@B�V�<k�N'�O
�S�t���p"I
�F��"Oc�:dhXQ'�)RKz "O�"Ѭ��H����LC�e1E"O�*�^<k��98�}�Ƨ��/�!�D� 0�@��%��Z5�̑��Өln�}Bh�~+�f�阖�Zr,���S��y��پ5�aX�jZ	0D�Ój���yˍ�6@�e�a�݌+]����ĳ�yn�1 �nt�1�+Yג�z�X��yrG��nhr�[d
��P�.\�E���y�	�{y�)�u��=pĈ�G�ذ�hO�������d踪�h\�L�04Z���{�.B�I�f-L9���Y�w���q(	+N�!򤘾@�����i߭)R͡&'	kd!�D�"�j(���C�r)z��Ńz!�$J�����^y���J��$!�ާh�P=*���]lN!���L%|���
�O?�Bi���a����Q'ؘ� C�b�<����`��iƧƕ+������h�<�M��l�p�ȍ4/�1`\`�<�� ڟ�	裌O�l%��L@]�<Q�l
.	 ahtD( < ,�A�<I���Y����3�N6C�9HTBAy2���p>�kψ3�Z�`.־*�.<����F�<��a{J�˴n_�-	�a��M}�<a��;���%��#��Lq���S�<!�Q��`�a-Ȥ;7�0��h�<����X*�QӠ'�*eP���dx���H��X�TE1 ����0
�6ΰ�/D��xT��;+�%��g@(�����-D��R@O�=�v �3���M5@Հ�8D�����["9(l���[]�""+D�0[�A�9/(�d����u#(�')'D�T�`��'�J��1��%q��v�$ړl�ʥF���:�YxB#��w�E{"C��y�ד
+4<��nS�c���q�ԙ�y��(In��QL�n��BBꖜ�y2��i�$��FC��T$at����y��qK �:N�(u�S욑�y"��<J�nq�΅�L�豚sJZ��?Ys�x����(i[��$:��m@�[��u�'D�tKwgӺ���`P�hy����M2D����V�#������^�wS��Y��;D��b�%E	7�1�s��>~ٲ�"�4D�,鰡ޙ/���-��LM�=��0D���q@�9��G� ��6�WM�<q���~8�D�uIߧf��p���$ S�J,D� �W-2m.}YP �	<���=T�l�VM�D���V�3g� c�"O~ٛtNV�q\�Ԫb'�3?~N� 0"O<͸тI�l� �[QL	.Le�X`�'�h���'��ı�,�d�8��3#�JD 
�'M�2�aP3�N5�6H�jLtt�	�'��(�+H��<���S�a�^p�	�'��8�-�B��X���ދk�\=��''E�e��^Blu8sņ�3`���'��	��1|�05����;2I�`�����F�Q?e�F� �^���u�J1	qx�R��/D����H4��ۥbT�0�,=sT",D��v�ha�
=��)zP�ƩY=�B�)� >Z�5/*�x�l�*LNܣ�"O�h� �3o_:�(���"�Hk�"O6��
�?<�$QG��0 ��'R��
���S�c �).��%��t���G2c�:d�ȓph �$� !��-B#j� פ��'���#D�*��<Z�܎-C����I�����I6"ȕb�� !B[Լ�ȓR=29+�c(�~�҄G+�͇ȓDܬjaMمN�4��Uk
=P0�0�'���(�~en<�4�¶z,����D<4���dWJqB��41|Dx���?�H��ϴI32�K�| �ӂ�(�`��l6�9�ۇ[u|�s�K!%f�%��E�s��
If$�C�#�X�T���	�'w��I>Z�BIz�"�,I��!WfߚV(B��b>\Q�K"�|d�tB\���B�	�ﰐ#!��=;��9Ұ�Y8ߘB䉠e#��h"L%>nfI!��9<�@B��h�c�+
(��@
��ԇ�nB�	1k�������!����;�L�=ɶ#ET�O������MP����g�����'[��DfI �R�	r��]�*)��'�*�G��>�8y�!�X4�!�'�:�8�&Q�`��p�`B�;�B�)�'�8�b�,N:^��<��ߟ5�l���')�Kd�	!�!�AIS�vz����;)bFx��)�n����)��_�T�KbN�&רB�
?J��3���I� `�G�/NxB�	�WJ���E�3���O��#{xB�d�䍈K}�|0��J�jB䉎4�j �i�ZH�p���UwRB�Ile\�2��@Jޠ���;nY�\��^��8F�I�����r����Pɦ	�g"x�W��*Ѭu��D[\�0����Jh8��I����,1�|�g�W51� ��&B߉n���� � ��)��`�\����g�(~T��\�(O�A
7�B�a	�I�`I�*'jP��M^$z>ڥ3P�ĥ}�"�1S�?C`����!�(OBC�'�&6��\�<�:��տA�T����,�˓�0?��,�-���w�i�}C�b�mx���(O�Yz#h%}��i���@l��Z���!�^㟨���#w���ƌ���ϝ�NXPa�J5D����V2)����\�D� g#5D��Z��Q�d�J)�2ͅI���v�/D��;fK�H��VAB+g��pt�/D�f'�Y�d��@J��ˀ .D�@�e�E�`��c��B�)ѰB��K��tE��'�	3� $H`�6��8(m�}�	�'D����"!;Hބ���:.����	�'˾�YD�>`��T
oD���'�P\�t�02 �~s>%�'y8u�V���M�x�gf_w����'?@�'P�O� �'��>g%�eQ� ��؄�	�C�Pc3FR����b"�HC�s����ݣg؊=Jd!�z:C䉟p�*����
�^ۺ$�o$�B�	�R�LCW�;���ڊm��B�I��V�( ��	rE��dVo�,����5��*���ҥ�H<=��<
�AJ%!X�i�ȓ$�D������u�X���{&o-D��i%cI��i�k(����ro*D��k�JlHVt�2�@�P�����+D���Ǡ�2�p���5<Ϯ���'D� ���%E���))�5�Ƽ#rc'�	'��#<���X��_�y�Ŭ�Tj�:�"Oj9b+߰Zel��ϭm�.ug"O�ՠ`�.] РXR.9�`�B�"O� ��h�JF�~r*$ �*�o{u8u"O"��dX���9���=�� Au"ON=�dN�$B:�rBA���(2��OX�}��6:!�0�����w��-U���ȓ��t�g�ɪ>���6ɘ+*
!�ȓA,,���nӘN��g-�$l�ȓth�%���"\�����$U�1��}��-r��9	�*�jd�LJ����A�h	(ԥV�$b@��Q��I?=����D�29����Wh�1Rh�sE�9,�!�dƙ	��90b��x$�%rE*^3!�H/�Π�tc͛
B}:q�Ю[!��H���h1	��0������7!���'B���c@�I�'ezA��	џ0˶�M�M3��?�O���iG�"Ӏ�R�^���^�.�����?i��v�]����M{d��",7�}>�9vZr���NL`�s"<�� �S!���b�q��Ct��S*eH0�rc*k�l��'Do��#>�Q��П��ɥ�M����dCϨ%��j�E_�%QV�A����?Y�������X��D�
I��Q�W`��X���(�;?��O�c��'�F`j�)�ԃ��8(�/��b�
 �<��@"���䧚?��O�ܺ�ͩ�䔋���h� @c4�	<�h���RH�>��S���
�^�0��Ջ!�'�V��Ij���ɇ{k4�i� �9� D&0��$l?YT�O�T>�*mO��Ӷ�"N����K��s�8�q��]~%}�'�>��	9��'O�5�i�@�.��' h ~=A� }r��E��'ByIu�  ��kl� Dc��􉉒�I-H���'ox�'u'��(v��E� =b�C���,)��a��'&�]R����E(Bp�TO�k��!�탚#���H
�1��/-�ݥO
�m_�^����˹q:���`�5H\�*���O��G�4�ХS������[�B!�����{��ӧ�9Oh
���j���6-�v�2G�J�X���S�0�e�'V0){�'g���i�O�|PA�]�2Z��S���r��K�UU�	aPE��D�s�x�C��@�B��3"�Xu/�{hx��2+�O@���``�#%F��-x4 ���L���ȓ9ٶ����)zRU;�*Ѿ}4moZ��L�Ioy��'�rU�<��5�e;7�.\s�-Νa����C.M"�Ms������O@y�O�2V>��	<7.��0,�9:�ڹs���F��d�I<y���$�I�<1a@����b�>�x�7ȏ32!�J+f���Q��*{���&$!�X�ao0-F�İ����\�k�!�$S	N��� ҒN�*�f#˯~�!�d5��RW)C�D�rYbבG!�D�%�`�(�м���G��"F!���:��� DȮo���� ��8C4!���Eȸɨd��<�n�����t!�1�t�@a��1+�
q"Ýp!�d
L��U)↟�6��ŀq�S1e��ۋ��?͙H��R�&Y��/�'-�uX�n+D�<`wc� 9�(�˚�/�����(�	,�"1	�`�Y��b@�U�cȘd��.�0u���IBK��q�������u����a��#
�\���i� ���$�P��M��M�NXa@��A�X8��cA'Ew4���,?�d�B��^N$�4Ɓ ��1H�
#��a6�J�ufȱ��F�kr� �c�6���f���N��'��Y�,�:cb�=�IHj@�� W�t(�M>�O���	-���� 7zHP����o��O�D����k�*Q��!$܉U��=�Ԑ�ƪ�$�j�i� Wc���\7�`���S�I8nb�����4�?Ɏ��,�U
ihE��3�uA'�����'�"�'���P��߃A�أ'�ݓV�Tш
� �Q�p�s��=׊���EޖjBy���_�6�0�����?���p�����?1���?���2�0M� !�K���GZ�o���ADE��<w���'H���Ű��� T�M���Di3?�p�J+i⒱���L��n�k��5:�f|�6�T#I�Ү�9�|ՂJİ[�t�'0���;V;��G$�'�L��S;N�P,�䪚7�M;F�iVB��:���,OH7�L)t���6��B�c�'v��\��?F0��	3T4�a"4�ŤOV�Ez�W>��'|1'�X�)$a�֋p�ޥы��<�'4���f��힭��a�7V�dE���hO�>� ��k�'N$t@�P3�����R�"O�ea�ـq��M�V�j��+"O��æ�'M"�RI-mD�컧"O`|���D�9tr$y6�ʀ3�PU��"O�H
�`$'%i��������"OBq�A�5%�� �M�7���"O��RSg7~�r�J�FT�y� �"O ic@,o,A(���\�	�"O��w(�����*�;��m��"OB�Ձ��T�	�(@�P�����"O|�#A�	,����!'�X�
�� "O�"���ܕUM�
�j\j�KRi�<y��Bt����V�z{�aQ�eOo�<��⛉3Fj�{e�*X��Ey��Rj�<I��H�{BJ]�S�.w��(rHDd�<Dc��6+�(� 5 ��ؘH�E�<I⓴;�&i�둆B�WGCA�<�cL�;��88ڼq���Jn���ȓ8�p=��b<)V����m׃@X���P��	��/��i@��Y<<���ȓ�J ba��=�X�bN�@���S"*Uڧ+X�2�x�d�^�6\�ȓ  �!j��8!@q×L�Kܠl�ȓU�
0 ��3�|:��Բja$���F��k�?k��DOҮUʊ��ȓgdd.L�bbAD"7�ɒ�BHT�<i�� �+� U��[�%�$Da�JO�<�� ]�<�:��=1޼��tF[p�<���*>�0�7Ms����'�m�<Q`�T8T���i)'�h)Y��D�<i15~Ƭ���]&c��Q�צ�w�<�����
�*YS��;кC�IXU�\9��ń\V�iW�G #�zC�	<r���(Bw�<�R�B��NC䉸B����O �/�"M"  �	`C�<-��-
c�M,�ȫ���<��C�	�H�������x���AQ=�C��pvŸ��­��ѳ#]�[nC�	.�$mH"�G"��at��+&cZC��<3oz"���[�aAf<>��C�	�P��hh���a�dea�҄��C�I� {P�����D�`�t�&Z4�C��g~�c���_b Q5��F�vC�I���ղbׯ�LX8���!�C�IrT�����#QLx��J<hC��&$�X���NʞtPp��͔+unbC䉬/�6Z��_8}2����ӵzs�B�	�7�1H�K�r��ȗ�ѝbi�C��$	��E�r��2�8�i�'�@C�I4J�4\�`oU�N`�lȖf�A��C�&?�`I�4��J�dt
&�y�B䉞)zdb��!f�:h��'�cC:B䉴0�Tc$�	b��7�Y'3�vB�IY �Pi�� ��7bٓo�C�I�v2�ᗈ��z��}�p�� ��B�ɨ{����'��MG�qpg��B�	�K�u;GG�5I[`�s����B�ɯR����3)J<�!\�B�ɱF�B��D��+D�a�@ 	 
��B�I�C�n) �H�*��yJ�oȎN�xB�ɳ�� :w�##����U�4e�RB��!O����*	�В=)��%�BB�	�]h|asȦR�<ѳ�"	�l�4B�ɐ&�ei!�]� �J��)&J��C�)� �8 �U�5�R݈������c7"O>��w��c��\S�����H�"O��f�L,)\���D��_���"O����=p,A�UW���P"O�TI��]/xwI������F#�ye��c0�SP��<��34K��y�
�bx�A�_�0��x�r��y��#�~��B`ՙ!�L)Ab��y"�E�O��ecD���d}��.��y�e��z��5�@JMs�1�Nţ�y�͵�<-�D�Q�R��M��y�J�05xtq��H*��eP�y2��B�,w��3��Q�~�&i"�';�3bj]3p��GFQ�J�fU�	�'A�`R�����8ه�A�3Y
��	�'�DH�FU�x(��΂*يm�	�'�:<��KR�H�@p�A�8�L)�	�'��Xw�e�JL����8W���'^��x7��)'q.pQC��iִ{�'>���j�#'��	2 ����;�'E@u�`��$~o�%ʗb��~h�L�'�8u4P�L�`�'�#u�u��'.:�HuBѽ\�p�q�	ؼ!綍��' ]ʥc�'2��ݪ��� %��'�x��
�	T�ua5��A�'dܣ�c���i�lM�|"���'�� J�fH���x0c�J�#><݊�'����Qi�|�|���KMp���'j���*3'�uh�.CK��A�'0(مd��>R	�5=e�q��'
��1�a�/ߴ����B;���[
�'�4X�L�Y�����04P��
�'�l�B�ݼXr&���L�7;P	�'�${���������a�8�p	�'�l�ǖr�9��$N'X9�'�d�i����.T���بJ�#�'��Xr�
%[�`�l\�F�$)�'�IQ��'�0���00�(M�'q�QK''),J��.�>��Q�
�'f�q�^�2��̹"i�Z���'~�jV��+2� $��a2�@x
�'LVA�RN^&7�|�S'�`d��
�'r���c"/~�8�r��#Q�FX�	�'[�Dc&��ZR�x�!Z<A}���'�����M `f�pcҗ5l��[�'��iʕ$��.jhZ��=@��ph
�'���zs�L`Y� A�?���	�'ZH���¡
?�3WKC�8N���'~��h���N�D�CL�5�|Qz�'U�73\��H"���;[�d5�"O�
2#Ԯ+�� ����\։��"O$U"Ѡ�K�<@d�Nd�9"Ol���xq��a@�䅋
 A!���:?.�m�a�Ēn��e�$�ѐ�!����ט)�&Ɉe!��B� �#!�$��Y������7>�D���Ȃf�!���fVXYc7暴'��y��l�!��P Ě�bAA	�@��(>+|!���h��:�D���h�C�B�!�$��Z\ʧ�$Bs�y)GOS�D1!��g�ބ�$FL���Yj�(/x!�dY3v4�s�F������rHI7t!�t�r,��o<�T	����e�!���(���7 ��C����t�Q�b!�� $�򤘱5Ֆ�)%%D�QH���"O4m!�͒,.�T�xFꎚ6���g"OJ��|��:G/Z�F	���'k
��m��X�K���QV�M`�'`j�ʦ�
J�H����4F�x��	�'!A�S�턭�BB¥'�b��'�<\ W�I�Z�d� ��-6�*
�'՞�ۃH\ )�F�(P��5C*���
�'?�AbB�(EU�T���8ݨaH�'Q���B��&t����WaI3j
�K�'�ȭ���̲SzH=B�nD�'�3�'%Ҝ��g�0^9z�nB�b8� �'�����Q@�$BW(ײ/��8�'�t���(D��Fd��5��p�'ި��Gc^�eQ�La�(������'�y(���Z3��
Ʀ4yXh(�
�'K�i���:gE�<1T� ?^}	�'��{s�[x���s
ݭ:4u[�'�z�"�'̱������)��'l
�	�N�W��֪�s@Us�'�F銲HB�D�v��թ��h��]��'AbQ����3LP��k��e�")��'�>��R((2�is��A�F�Tm��'��hJf�%$~c�L J�.<Z�'�	�	Q8O]N(90�ѸC�:��'�N<����8� �5;�jE��'�|�Qqc����BD�M@�2� �'� ��diC�9�P�k�o΅9P�h�
�'%$E�vK� ߂���3ۤ�R
�'���rƂ9��	;Q"@�(�^�Y	�'U�Lx�J+_h�Рs���*r�+�'q�XjBa	1�����/��0fQ��'��8�aH?U�(�����"C�Lz�'
�@s�n�(pP��w�Ó4�|��
�'�n�[��!N�>m��U�Y����
�'Q4
b�ܛ ]
'ɚ5T�j
�'�n��s�[���Zf��7(�c	�'���h#.�~�#cF�$(�ܚ�'���S,ͺn�ҰZbL�$�$\��'o��#Q��~�����.Hy�'���c��[�2�HPK�/S��P�	�'��,k!-�g� ��*K��ĵi	�'�ب� �86������E@���'/�j��.L�R��4KT��Mi�'(�
�nj����۝� ��'�������l�zlK��Z {�D%z�'*N5ag!��f1��� }VB�'OL���X;�L�g��ӏI�<��dB3!GČ*R'�0(<��φl�<р�����@S<H-ఓc�Uj�<�
�>Fᐶ��-@Ș�C�ψf�<�E��h�хc��T��!��|�<q��J�M4�,)��5��s���{�<��m�/P��(a�� �+B�E�עu�<ْC��xǈ�@��|&<01�j�r�<Aq��L&>@z���P�jQl�J�<!�d�N��t� �;h��Ԇ_�<Iތv�Z�9�lϏw�8l�qA��<��Aq���T��3t��آC��<y����~��\���/3��$y�lR�<�����~(P��U����h�ŀr�<9bGT�� p�Ä�F4R�x�'�p�<�FE�>NC@��s��+�!�U��k�<�D��?l	p�eK�:H8�+2	�c�<� \A��\2mqHI�G%A�"�> ��"O� �'/GA�8�5�@$DՎ�j�"OX���!�p�hW.A���A"Or��V�TzʈD#�(&-�"f"Oz$d�ɛ9��'F�%O>
P�/4�<��H[�w�<�D�̓xR΍���+D�h���>�0��;}��ˤ,*D�D���E�\�:%�	:u,����+D�����U� q@�	j.
�H7C'D�d�D#�% ��Բ�-��X{ 4rCo%D��R*ɾ�̊eg��i������#D�\��I�b�^�͌[�8
sn=D�̰`��
<Y2h
��*�:�o9D��
�@!zR����$U�4:$D����� ��-Rub��IH꤉v!D�LaTa�,��pr"�Z��P���$D�<�B/ �M-~�ˑ�ڽz�TcP�=D��(��O�'Ǭ<�sa�u���:D���4����蕡1���n�Ƅ17$:D���JR�w��,�P�������#'D���E��4u��hÞ1��+�) D���S��ߒ
�Ó&Hs����/D���$׃<�|@[��R�gؔ۔F9D�p �T5(�'Ւ
��T��'D�ʢ쐧@�lUP��66���C �$D��;�&j�������?i �D7D��+�(Ӻ/�A�[)_����
6D��q�� xf$ ��>vx`���5D�4 `k�)�ͺș�eBt؂��/D��@�L�Z���ʵoʏS'l��2D�<ҷ�M!@QJ���1�@��i1D��J���
ZU���� o�"�Q��)D�XZ#�JE�d��wH�;�H�7D�x�N	���IK�Ʊ��j�H5D��r�Ţ�b�`�J��:oѨ�!9D�#�h�"'
����*Ùc�����8D����,��n,x��U�W���2G&D�|C�]��� ���D�&�BD"D��yq�ӱLx�d�"��򽐦�;D�|1�KS:��!�6-��{|��*8D�(2Չ�"��լD:=N��B+*D�(��(ۘI�����B�.!�O6D�r�Q�
<�s�U3{+��DA5D��id��?,0��k�H&x��sP�'D��)0N�]4L��@nH�O-���'l%D��;��	[[�m�I��ي��/%D�����<U�M1taљ|�b͸��(D��[�H�4�ИA�_�a42�;D�DӀM
,-,A;�/x �Wd,D��P��<�h�����vn�	 ec+D��r5���+Kd�9�B(7��}��&D���I��&U�P�aK��E��}@g�8D��K6����
L�8][`J�S0C䉫(��L ��E��
M�Q
:(C��,�&���+ Q��m���	9W��C䉂ae�E�ڱ7�P���嗇�C�	
/�:��r��xZj�r��A0�`B�I)9�f1��"���� ��� D(NB�	`ԑ#i϶?3,uxd�ΰQ�B�Ɏ9� ���E*?�F	�(H@�<a�h�8�Vi�$!�F�ik��f�<1M
�Z�`�1�O [L-��Uf�<yad_�q6�1`�_�n�$B��e�<I��'f �����L�c�~�pm�V�<� �7(�6;��Ð��ƼX2s"O �"@'�?�Y�B*A��PջE"ON�g��D�Z=)b���vQ�("O���TIT�"�La9&�@�LG2�z�"O� 
�	��<�l��rbա\�jt��"O`�j�]�-�ꀡ`hX�f��0��"OD�C�D�p<N���G*��"gA|�<9�_�HR�I2S�S"T�z
U�Yu�<�!�U�~�Xw˻MT�c�/�z�<Y!%�M��]q#��"R�c!�x�<)���/�$�0I��u?ʽ˄hz�<��C�,\R��a��8Z̔k�)@�<�W�ߔ0�j���G%`�X���	e�<!���	������7�4%;��W}�<a��G7.�1�7H�(����Œx�<)��	?�P�;�参=T%��'L�<��
 !JP��S��S L���+D�<��F�|��<��%�5��5#��_�<!v�Q[+�u��� }�rX�'+\r�<ywAL�������#�e�<���u*L!3$v�]K�j�<��`��l:p@�
[�r}<��	�{�<�G���J�`�ҁ��.x=�����_�<�f2C-j�ȥ]�u�:=Y5�BY�<����D��p�� O�^\~�j0�q�<Pg���Z�J		WL�P�_s�<���	�@3Ȥ����Kn�+�fSv�<yU���5�1�� *��=�T�Xs�<!�H� A�����l���Q��q�<9r��Lh�i��"��rc�J�<a��ӃxBh0�倒	A���O�D�<��H��q� S3�܇	��i(�C�<��˰�☻�N�B+z��e΋@�<Q��E'���g�}����G�`�<��'A6{��$A	�Yi���p�a�<�bJX�����N�
tz�Aԅ�a�<Y�GN6%��H7B�}�Jh	�n�`�<����fx`����a~\1� �C�<y`K!FC�Y��CƓ%`"=�� �H�<�d�8F�t}�EȒR������Y�<�t͉KFL�+S�K4�y�D�X�<!sFM����iJ�{�����X�<Q4O*e����դ-�8=��hSZ�'�R(���>�' �l�̄�Xpb��L�2��(X���훁U�t�����jmԨ�;]�Z�C(I߉���Te��.��ԝC�A3;~�%�f"O�[bM��g��<P�A�	���+�[�<���"O�N!�&L9�0<����@M��9��R�E�$�z���@X�H��(	�AՒp s�A�G��)	e�O�/����5E;��{�'e�a;an�0���b,] f�P�����
P�Y�r�̂!��8��HZ����ɶ�Q�9�dH�H؆N�xB�I�e�N|��)�>:(�H�_2Z4Y���{R��ש�O�����t��yҢ�
0+j���ٯgR4��N���y�+T�(h�l��EΌB1��_=B�H�J��NK�)[��� T���g�'o\4�!�G2lx=Q��H-Tպ�	����@Q��Y�\5�u�[/4�ܹaꇜQ�v�ps�U�"'��F+�}��|zAeF�l�@YSbߣu�°�v-,�I�p,�\	���YE� aE�)<�6�?ѐ��g\
����H:�Ƽ�.*D���VcR*6���ˠ!A9��0X�-��/�&�`��L����!��MG��%h��0H�u�$H���ͬl�2�0A�(D�X�O�s��6��B�$���E��M�w�0B��R@��⸮�X�����U�`tu�0 �w/^����4lO�"����>����|����W"�4Q~~�j���/(�%�S�N=?�bI���FJ"��T	ˆwϐq��1!mRc��AgDX��(��fBl��<A����3� ^}suo�.d���"���J�z'"O���D��-h��%��LQ��^=ZDND�܀�L�XO���ŃEd�>-�X0��6�R�TB���=l�rՄ�L��M�+�=G��ʑ���p��UÐ�	1��q�Aш\��
�&M�?�>Q!�V�e*�x�&���%���I���K�'�L��U#X!�$ő���QLa1�6S(��EB<ٰ?qW��^���+��V�^���@�'%~��a!���*�i!���)��2��q���9zhpQ��#�y��A.�^Y��]�%�H��t��~��ʟ@m�-B������S�m��ࠁ��$`qΙ�PJ\�U�C�	�;�Ҽj�G��r�:�^�?� �-�0�jqF��2 ��	)	fظ�U'U�Jf6��V䍶y����dN=$$�cG�� �遠%ߘy��M���-pDlp�	5F��Z9*n� ��U2�ȰD|2�֨ �])C�)K�a�T��$@\H"R�X"lQ6&E!�Đ%U�BCV�C�(��M
����	�b��E�?E��kQ����'hH`��y�R�y�O�IԴP2nԒ,| 4��Ɓ#�yr�M�3*�uq�����.�0�Ć�X��2P+�bt��ȓ�J䱆ȓF$D��b�^:Y��آ"31���ȓ1rP�@�D7o�8�2�Y����q��!��9�:���џ7�2�ȓg�]�2���)\F躖̓y�*y�ȓ���R��~����Eɓm�愇�iK�0+��.t�6]Jm�/T�Є�P;�EAQf��-�"U�5#S�A0�p��Y���E�gt�)B�W�b�v�ȓ;�с�G]�M� Ő��>� D��D~�C�BΩX�ʼP�,̣&h]��.r�L��n����3Żt�܇ȓd\��ԋÍ�\2��cX���h���d$Ĩzi��+1�	���*�x[�.Y�(�ǉ8���ȓN�h]:�χf�Ic�Д)u���ȓt�j�ў&Ǯ�!&%�4c,ԅȓ=V`$�b�ֱ`���;f��fz��ȓ#(e��?a�j\���̑R�(��ȓi�ȅr��If�cg��eE�P�ȓl�n��H�'FtԨ�1��h�%�ȓ3���蜗`�N\P�v0rY��>��C�IR�aE
�+qr䘆ȓ,�bD���ڱ �ȩ	E�ťW�Q�ȓe��� ��Q�~Ѓ�I���fa��J96)�"��3��{�eD�,�E�ȓb��-�D������/b>���tr`�RpgN;r�\)+rZ�pWPȄȓG�X���-�>)�������bzF�ȓ�r���-5�>)��([�&іE�ȓ3b�
��ӄ<~t`�3��<��D�tw���p1+�!Ѱ����-D�ر��ˠe�<�(�D��j�8�t)D���3�V���*�)̦F�8��v6D��p�K	�|����8lYaS@3D��bė	#L��Q�!�@��s�3D��K�-�0kF\ÄF/��c�>D���u���A`�=h}蕁d�!D��s�+�'�&x���%C��)vl.D�Pi���7��x�&�X�*�u��*D��
�]����%EpH�}*�(D�챁�̽i�<��4�=��-� 5D�h	��
$}"���K?�i��� D�� �#�FX���6��d� D�쒇�ҾK�bU)4O���M��)D�� ��h�Z	�����"���Xc"O�PI��@u��zVd�17� ��"Oh<���R��KFJ8��$"O��z6Ę$!�x5:E�~�V5!A"OFt
��\C)�д
�.s�4�2a"O`�P�U��8U2����*�"O�|�DY�$�~�St��8+���D"O�����)V�jZFOVg�f��"O�9" mN���)�DܐMRP1h44� K������M١;R$�!):D���!��1$�Y��רJ �Z5�9D��*�*�R͖��V�k��%!�e=D�H!Ǎ�3Mu�A��
�:�>��An9D�t0�c��UqrH���BH5D�4��Tb�RC#�5nn ����2D��Bv�5n'�A$B�2B%��1@;D����S��e2+�)�q"��9D������,!�8���BI�����j4D�tPD�5��b!�+��4S�%D�䊁�5�,���nϔ�	��%D�Pk�,�}5V��̆�UE��q	%D�0��K�r�� (���_�,�r�#D�8Ñ�9k�)�d�ߟT(<�p�%D�4��j�=��	�@�%~�����E'D�蓑�.EX�e:ag�5R��ǁ%D�����W�� <CP)ٵ#㎬PD�#D��q��H��M�vf��79Z8�s�Bh�<��(ϐ<�.`�@S�f�<��1��a�<�G��JCr�
����D0ke�]�<���3$�,}"q��vlt���C�<AVHQڼ���c�8/�8sC��t�<��.�W�0 k�;�؇�Z�<	�%ӝUal!�B\;;��X���n�<�rD5-��c�M��f�� t,�_�<)
J7TT�Y�PY�1BA�T$^D�<	�M�0F�t�C�2C)����Y�<abBߎ}���e���edtk�+�a�<y�'P�p�P4%�4�%s�,O`�<I"M�	4A1�Р0a�jA����c�<����Q�f������.�xU���e�<6�M�/��P���K��x)"*�u�<1�苰7�:D�ڲ>���� J�f�<q��Ϟ#�y��G�PC�� ,�I�<���<I�p,���1�d�
�,�|�<�Vf��e����!e��F~�!��	�z�<�E�N�3y��@e��u�-pqņ\�<�,N/ x�ThV�`<������f!�dڰ�h�gŦI�J��I)KS!��
���N�%[���1���1T!��-6�����Q�#�\�gn�Gd!�:hV���ǫ4f�dD���Y6.�!��t�!�eDى ۚ���ƩcO!�$۫�,%��a�8�p�&A�'B!�_y��AY7x6�s�E-+2!�B8p<�l����$z��1!%�B!�d�H�l��,}�ՒE�^4j!��Ȟ,�b�b[�פ��"��h!�H��.mRB��V�(Ļ�ߵ�!��2ra�Xb�@�!p��k� = I!�Ѳ'�l��&-ȧ?����R���1 !�D�
�l񷍗-v�Ҩ��[!��?c�fd�`�ְ5|����H�b'!��-
n����A c�f�J�M&!��A��ݺ�n@5���d)�%!�� d��Tb���鈲�}l��"O���� P�P��jTź�"O�L8��%:��A2���r6v�K"Or\�5 E9��-��*�UDJ���"O��r�ʔLAV]@%K�~���"O��e�%����Q�^�c1�[t"O�1pÎwh �6*7,�
5"Oސ��&J�1�D���K>�)qt"O�b�o;������..����`"O��3&WQ��Ī���'�	�"O0	ZR�� jx�����l��x�C"O�q�lֱ��q���ּF��(HF"O�
b�� }�9+t��C��/�yB��,<޸ӕ���bq�%�4a��yb�πZA�𲦯��Դ�r��!�y"�����iF�����E��E^��y�K���P��c��T����f�I��y��I���ߩu�<�cAI��y*�1�rc �'_�`��Ή�y�X�;q�j h<n�9��&�y2�1X���5nU�X|0���G��yR0�q��0L��B���y�,V�?���S��A�����!���y�G6-�����W�<��p�0F��y�As����ҞG~`��t퐃�yR�R|3�5���./�"d�5�y�(�+9{�a0��L*�4)�0�Ց�y�'�e�=j���;�1�0�A��y&Uh$|��#�S�8N��y"/��"r��;�]�Eoٹ�y�bϾ
��P�1��n,�ԅ��yǅ�N@l��׉����GB7�yr�ŁϞap��:|h�0�&̇�yBŒ�=���
GHPy���tD
��y�C�=�};�$�8@S�a$��yR��dVFdАb��>=,��mϠ�yB�/���q���F�)`�n��yBL�3��R3��s! ���%\��y�"��0�.���B�q?��[2LT��B~\Q{�GUQ&%�b��*��ȓ?�na�pb����z��!�l݄ȓv��0�$J��bZ�]�d�9T ]��g�lEjRI�8%�tO�y���ȓ	��8� �0(�ũ� �\�bŅ�?V�%D��0���g�
�pȆ�,Kt���I�sc����)?_|`8���R��@E"g`D��
�fe���R�^��D��
��d0���j_:ņȓY]�IA7���vwޘ+�+�L��X��V��[�h�kw�}�W�=H�z��ȓ4�m����|<S��Q;L6ч�{@�%K')�:Z���޲�&Շȓ`xp�`7o�<(Z}�#"p�p��ȓF~�Y#��.����V�bnل�}�V���Z�3bāS�+A2Bƨh��?��Has�˧6�@!B��f8p��O���偌�g�����.Tq�`��ȓA�`Y�#�3{�.)1!�Ia� ��ȓO�`l����D�9��L���-�ȓ!����P��ިKb��i��ȓ[��Qg�.G�L�c`���q���T���]��[���>nݴ=��;��ͨ��&-,E�E.�9蠆�!D�SA���B�"�)��*j�Ԅ��S�? �딮E>&�MIT�ڶ��Q�c"O(�`aG�@H� PF�M�NxT�FO*��ºX�N���$VL�p
��ѣ^!�dtV8��-��-̨0�kC)�!�D��I� I�#U�"="0yGk�0�!��ƹZ�T	�$ �[@� �F*�3F�!򄚻�&h:`HΚ3'LT�	�<�!�d��U�łGBZ�lj�E��Aí�Py� �U�����iIx_he�%���yr�̿a�VX9eH��<8v-�yr4S�0���!؆	<���j�y"��U� 2ƀ���,�U�_��y"_.@�����!���b��)�	�'�h� �G/#��C�ŋ+B.,b	�'/p=�F雃7�, �Fǌۢ���'V<����R"�X2KH2$�;�'�Ld�C4%3���v�U�#�� i�'� L��	��z(R�k�-)��L��'�H�b�Ε��m�� F?�~)��'��0�B��Z�u��+�~�l���'�n  ���&B;<��%Kԅ{ntp�	�'j6��pA�*����B�"�T�	�'�AӷFûa J��E�!N�q��'M<4C�A&�}RT�ٛ1|���'Y
��:�r<q�FQ6�`���'q��B[�k�Ęq�-ƥnt3�'���n.K���k�o�0rKص*�'X��FH�=xH,Ȣ�(7�L���'�ٺtfց&tθjgG.'-,�'��9A �Ys�c4���g�=��'n��3���(rh���b!Z����'{F�Q-�'Pc "(H�J���'s:E��Mx0&� OZ��"�'3,�`&�� ��؇"r��#�'�����%Q`��)d$U���P�'� [v�l�H�L�"LF��'KH�ZC�6T�D����9q�B��
�'<��F�ܯ\$`�2�Vx��y
�'�(Uॄ�M}2�X�% �H?:�`�'Mb�Scl��GY�a�U�Ў:�ȥ�
�'X�h�	��=u��+Ԯ�4D
�'ފ!��"�^pH3V.8i�e1	�'�h����؇&��LK�(�*���C�'�X�30��~�)��(��DR�'h���A�>2$���0�ċ Xp���'}"1p���j�T��0O��fO�yr�'#��{����d�A�N�e�8щ�'0�偕��
?p�5�мK,DZ�'IZ<��C��r���!ߌy�88�'���#P�[-4��wM�Hޒ��'��!&���2�60XgdC=����'��"�#ޏ Ŧ�v+�)Đ`��'��$&G2W�dsvH�(�ⴚ�'���i�����Q��H�8W*y��'	n	!�5g�:$����8F���	�'0Lx���.pn���M�Q��M�'��q�U��F���&�L��D��'�\)�	J�Z��u"�%z9��'ۺ��R�<E!�#��M���Y�'m�ԡc@4n6dXD?}b$��'%@��F3wSl�R4/LIɾ�3�'l*�������L�� >��ݚ�'�x��t< {s��'K2��
�'8H�P�ęh��|*�
�.؁
��� Ҡ:O�P$q)��	�3J��A"O���!,�c����˅?�4���"ON)���7=��X9sD2��d"OXm)V	��*6<� aΚJ��i�"O2T�� _3�)@/�g��]�!"Oj8�i6r���·��$ :%"O�Qa'ÈJ|��� KkZ�Փ�"O�P�ȇ)zY��EB���Q"O��8Ҫԟld�UA�-�]*uc�"O.� Da��*��(�1�N�N�i��"O�9���8�1�E����� "On��rm�8��
���<x�Hd��"O��ׂ,��]�r"̠[���9"O��D띂M9��S)2�����"O|(���1XtH���
�  ����"OZܰ�!H:"6�����Z�%�4
�"O>�C��"G^�)��6;w� S�"Of�P�	��±Z O5R\�'"O�I��T����:[�@��"OF�-����C�L<\v��"O�(� ���.^�,X���"OX$�j�>���J@-��e<�)�R"OB�@G�&�,�`��0:���"OZ)���+Z��d`Q�
n)�"Ob���F��,�Rܐ��X$�*�b"OF��G����j�j\-���[%"O�	��!��	�\z�j	�0�e�"O��c@��n��!jд��X�"O
�Ҡ	�pX$؃�h]:(��}�2"O�<����0m|Qc�l�LB�q3�"O6`餭��GF�E�IӗP7��i�"O`%s$�R�qz�����?�@� "O�U٥�Ю���0�E�Xm�x�"O|E2�#@$9.��-��]y�sE"O��)qE��f��I��F0��4�"O���v苋f��8�e�pbN�"O���tB�_pt��td]>k�=��"Of�*U&�V� GdG6\����2"O ��GI�p��1����T��"O,@��g]�<�>X�E!-"���a"O�	`��� R"��1�o\*9uPQ0"O�a�C�U,�u���Z��}`"OTA
g�&_e�QAX�@�r�X�"O��k"ˇM�Q�ԗe����"O��['ءm�$���	Vd~��"O��tR;z̚�Z���	U����T"O�@9�X/I�xC �6Ir���"O�QSC�Z��֍�2=�(9�"O��!��t6�%���E�w�D�3R"O\Ypb� �A!Ǆ�A�: "O��B�=mXijkݷ9Ŷ�B"O�E3�E�g7:����5I��Du"O,�te�3E̸��&^=��	"O��@MQf�4I�M9!�\CD"OIj��1��P�&�m�j,�"O�1�v*�+�Hŏ�U����"O�)�`��*Xv}�s�ʂ\�p�2�"O��"�dQ% �6�Hj�(��r�"O�L"eEM�H�F��V�9�HT�b"O��N� #��(���R�\�N���"O ȓ�C�9�R8z�(-j��"Oh|�q����)J!k��Q��q�"O�$�$I?���%�NP���b�"O�������J��8�$�/rt\���"O� �X �c�/CK�˒�3RH��"O�Q��7΂�0%�� :6q:�"OJ��aOS�Ul�X0Č�'w�.�`C"OdPU�¿Y
�i��c>�b"O�@�f	E.d��(�&��\}|8�E"OF����W{"�IӅP1�$�"O�T��(��%Q�x�rN�/x���"O��Q��C\��P�1p~:��"O������gI ��kU����"O��4mM�~}�IP���B� ��"O~����ѭ~��i��+Q�.!�9Be"O(����@2� �G?6���"O�y���\���u�ň�;��� 4"O$�pr(Gz�,|��!C���"O�A+�	����33��ye�1D�\!Bo�\Z�x��� {�(��.D�|P���/(�tt�p�U�k����B�-D�\�c��
3>�d���2R�h���6D�X�JԨo���p��w�����b6D�\���^���Z$kDRy �.!D��T�!Y"&,����cQZ�	5.4D����k_,*���nʇ��̚T@2D�X��J{��<�R�	�<��R0/D���Ӗw��҃�63���@Ə(D��c���p��ЇX8K��cU@<D���C�+6��]�$�9dF��A$9D��Ch��I���z���*`��͢��$D���U�O�JY�Ŧ�,R��!�d/D�0#dQ�G$j��^4U��� l(D��A�Ì2+MPH9w㜏+E�		��1D�pbЇ	z���Pl�]�n�s@*D�dJc`>�놆C+LdQ�@�'D��Ywb�=�ܩg�Ժ;�$c1�$D��"R��;fD�c*��?׼�� �$D� �3�++:�����A�����<D����h�,!Ɲԫߩ6��� O0D��{�e���X� T�\�I�Ԓi8D����h�aAb�
�8*�IRH*D�����
IV���Ǐ+��O58!�$�>=R­․+Y4��s/�:�!��u�쭩#�0g1`����&B�!���.�4e
��Ϸh�0k��J��!�d� 0��Xjb�ֈ^�Y�'�b!��5P���NŲV��d�[!��۸e�fX�e�ύ8.�4i^�!�DM0����0���r��M�E!��
0t6FE�էwP%re+B!򤞴c�,Ay6e�&a�-S����]!�$ثS-H���ӑV��)�ˁ�D!�D��#v5�'HD�lv]�䄑c!�''�ƴ�!է�,,�L1�!�d�_�|���[�px�5 eb�<�!�dV5|<,X%K;ɨ("vA>���l��(��}��?5���ԋ^�Q
�� "OXP�i�r zB��U�8��#"O�����m�2`�#�v�F)"O,�D���&�|,)��T	W�VmR0"O���� pʁh�;!�H��`"Ol�cT.��FP�������x�"O���S*�6�u��&?�ƀ��"Ol۔��^��E�?��<O!���8\�d��>uT��f�YW�!�䗎����j[.9�I	ah�?��z��dGK$|·֣+�}��"f�!�� ��r�S3_� ��!K�aĶU�1"O�P%���|�9�t�B���Iҵ"OV<sD/�h��XQ���b���BS"O�kBbH?3���!�φ+_����"O�
�B�/�}��B����:"O�H�­ԟ|"����o�zY�&"O,YJ����,۲��F2Zw&�1"OVLP�n�����H1)��ZL��"O�����	�����N5Y:���E"O�J�cɹR.�T��!a/¢�y�	E��I4f
�W��� F���yR���τ9a��R xD(���yB!_�2���`�Q��YJIȤ�y¦STf@�T�/*u��!�y�E��MH�BmLQ��'�y�%P)@�!Ѣ �3���Ҩ��y�ꂇ3�.������w�n0��%�0�y��UJ8=���]�?�p��-�y�K�e�9��M"�=�2�	��y���*�`5��M�9�^a�G����y��H�6yR�ʀ��8�Ջ���y�N+lbn�c"m�tٰHq�i��y�C�C�Jp���l�D���R�y�.Y '�$hpg��l��=Cé];�y�(!��C��9T&.���Gߕ�y�̊?��M�wM�w�4�!΀ �yR�߸Y��#�cHp�f���a�*�yrȗ�6M���ǻeXf�2%���yb
��~XM��L mL�=B�à�y��׶��4A�
^��;DC���yr"U;���i�$�òq�����y�'�^�p��7)R��,9g���y��6q%��"�Á>�JI��%�ycW�!`}PV��)s�+V��y��R�[�L�����0W��`��
�'r�Ѩ�Ԑ!�*B  ݼ�@p��'r	zA���]� �����,6L��'�J� �C&b�V�SK�<k�f(D�<�W�Ι`B��s��;) �X��%D��F�6� 9�e�+/C��2�.?D�,�
� f�|[P�%D���H�:D��X�&Ku(��A� 鳁8D��PA��K^�;�#�z%����N7D�dV���LdcW@ 'v���*D��e�u���sЪ�o�<���-D�@�Q��2LՂ	�Ǯ[�`�kCD,D��c���V��<eI0\,�s�I6D���D�(t�ܩzJ�?u��}���5D�0�D�̰C�h�W#�+i1�E#Cg5D��P.F#tt�K�ő1B���$')D��*T�ƚq~ T�m��1O@�!�&D�h������ i�ɄM�1E6D�$���ȃc:9�D��Y.��` �6D���"AR�%y&HWe�(��2�/D��HV��b͸W�̋�̄j�" D�@Q�j�1?h�X��k'4�تF�8D���F�1$Æ���Ζw�(i�*6D�Iw D��&-z��
:X���9�' ty8pN�= o�l��'l��19�'��T�z.��ER�}���a/�A�<��&F��ػJ�*�"���v�<�� ��P���'5"���!5cCp�<	V�6#`��ů&>��enj�<�k��a�M�䅊(<�Y����^�<� ���,	� !۷"M�~~�Ļ�"OP��P81�$�V�:`t Y��"O01�E9$�z2�S\d��V"O�c �I�Y�.���jT�	Bjs"Or��蛍;w0��El�V��p�B"Ol<���N�E�X��wk��$wL���"Oj谢kO!t���p��E;a��T��"O�ql�n:ƕ��N(.�6��.D�L`Pa[1_�\��ՀZe�X�&A.D��3�TK5(t���¢,��p�Wc,D�pj���8a�P��(K���3%�5D�$� F�1 W�y�eF�0do���O(D�D	󡐂('p�2��M�F~.ʔ3D���G)�)Y�j �"��� &�1D����cE�4�5#��F�d��0D��b�K	Q4���G!�}0�)0D�P�fL�0pO�}BB E����a�m���$S�1���iayK�7��uӥΆ�D��5�'�L5�L8pPn�<V�l���iP�Pk蟔q�����@Y$/Y! :���5��V��0��t�G�M�jt��~R���nGF�{��~b�X�X�JMTb1�P��X���D		u���dN��1�[?˓)͛�^� r���؈ЛaFҠd `ҡ�2D�$h2��1h$��e��q$�]��-\YD��eӤ�O����^�^Ǯ�1��͉1kԤ#�-ѐh����UL��wkR�@���?I��?�T��	�?���?�e�Υy1v)r�A'�����|���@���2/�F0�1.��|��ݸT�i��+��$"d1��e���b킵{u�Ջ��
� �vEA<[�`9�Fd�d�HુM!S#�p��l��\4��mr��D�gȘ�@Dc�O�(	 ��̡4  ����K�Iڟh��u�S�t`P(��l�c�K�o�Ւ�I��y�.�8�f<�!�g�.�����~��eӒ��<�V� `$���'��P?���H�]Юhwj�S�&���j٫O~E����?1�5�H�c��p���J��=ꐬ��(&�-�S����1�UO�}��c��TI�'L�y��59�Z��Vm�I��J��Z�	`,�[޳D�MQ�I���� �v �%D<�Br�|R" ��?��n����'��S|uT�����p��JF�0���V�����u���O� �ߠ:�@���чx�11�e�g��TX�4[Λֹi��P���RU�xy:��Y2j�.㰩���dW*K��%��ԟ����?�aD�X�I�A��]�s"����_�y*�e � ��K������z�'ϲyc���H�IK�}�)�B�	h�m���'���l	�S"Ġ @~�D�H��#A�j�hr(*w���ug��7G��S��Ԓ&����[�R:{����A�I� �G�H6-:{�R�a��lZџD�O���M�	5O�J�Њ5mҶ�
��_L?!��°>���O:Y1����%^�j2��E�'�6���]$���ƺs�aW�m]�(IS��:�0��7��W�R�'}��E��b�'=�'� ��lnZ�z�N$2�ðw�5�v�@�;�����D?���W,��U����A+��+G�L1'�Y4'ѝ!d0�Ch�� �v<�uE��M�ˇJj��5���O7�T�P.�# ��<�v�O���NRW��*�&�&���ߟ 0e�Yɟ�y�4F~��gy�'��ɔ7XX�R���(R��1��q��L��'S�9�������@�I�p�|Qcݴ�M3[Xu�J>!.����@�gD��*x�b�'[B +%
՚8����?����?iv����?Q���?!ձ^茝ч�4m�^�$h��4SĲg���5}�D�����I�3��	F�	P�2P 1NҳG�9`cA46�^Xj5j��n:"1��c�6y�����5a�f͒E%R�j\ �%�ĚE��O��a��ك�4l	��Ȼ,ϒ�!ҋ�(29��lZƟ�'9"�'/��	-iQ�0�DY�W�
��7FRO!��[�cj
8b-���	�d�,4�d/��-l}�	>�u��'y�'|q�� ��$   Q
  �  ^  �   %  `+  �1  �1   Ĵ���	����Zv)���P���>��'���qe���Ox�q��P�3J|�t"�+��aX6"OL9f���H�G�N|y���EfJ�h�Qjr6$�!E��WMvt�f拍��Ё��f,���Bzr��X�j��wv��jR�ts@Z����;�^iۤ��Q�0��F�{t(#o��[.P�/D��
���a7,�ybN�/ekȕ�eOx�1���f��!�7�ӧ|�H�h�}'f���?���?�Q?��@�_�U&y�u�Y
ȭxd៉���"w,�)8��?LO�"���Z�h� �'̦D����ƃ�9!<΅�fo��ti�PRK?y_�&lN e�/_�I��I`+ �ǨE0/��3`��lf�6�O� �E�O6�m����Y�P�	X?���5T=�-�A��]�����f�<��I�%�^9ZeD�7/
}���E٦�����J�*�\���<�Ӧϰ#L~��S`Ƒ ��Ĭ7+�A���.�?Y���?��pa���O���`>�%X
o�tQ#��I�$�iY��r�N���Z;*\�B�P�(�\Q���ܨ~�*\82D  }%~��-Q.R��U(��\�,�Dp�tC�5O���:��"::U�Aϊ<}D��O8Q���'���E���A�!*mA&����{�x�oǟ\�'o��T?����ͫg0���J^#Jn"����8D�HYH�ha�}��׌kWFY�c�>�S�H�'+"�TefӤ�d�O �� 4z��cd�!�R��B���JX6-�lu����O*���w	:��Gc�7Cd`!+4C��q�'
�.u��;]��m2�n�7=d�D{�f,?��U��,٬@�$1ڣ���+D���c��v�Z=R!�S?7����B��ў4p���Ox����m�IC��%��* ͂+J(z��Р��٦e�Id��|���pv5��@A-��BA��R6��O��!�)�V_�0��N�"/�$!��n��U�!``�ˮ���
0
:�qlZ��(���$���I�������)1۾0�b�߉	��2�K��M3CV��?1)O@���|�>1֣_�Qiޜ鲅S�.`��������bv�Ä2����V�V��E�TO�<_��96�D�d��!CS's ��ߙ�?�w�iT��S���O}���r�	��غ*$x�3����(YF~"�'�r���5�+��N11N�1Y$/��c\�O���h}B^�H�Ok4��f�F���;s-� Zό�+4Nw�x�D�O��(��V����D�O�$�O��;�?��NZ�!�0�2�4�d��[�E�|h��'x����	G��Eq�Y>�<���5p|����N��(wX<���ȸv�����~�:�qeH*/%F��(OҴQ����RTN#>��d�I���9	���'r���?ݫ2�V�$�� �E@����T8��&D�(R�hV:J	��sp�v��$��0Ez�OZ���#^ YЕp�/�DH�����Sa`f	�%]͟��	�����uG�'1B;�$=86 VdJ�m;��M<6B|���X��@�R�ھ*�
�p0ryTE~2�
V�*ձ6�N���u�u�-��A�K�zĪ����
m�ꌑ��"�]A���h�vL��E�	9G��g�.)�ݴ�hO֢>�v��[jr5E��5��ma�<ɖ�V?�,yI��^2Ė���^}�&t���D�<I5D�;0���័�'5�4�֋�&���C�F*V_In�:%z���ݟT�ɤ`	�"���~�h@�����h�4��ʇB��pY��
��=)q�΁�4���cX�/��"@K�H�� S�������	�����ZҦQ"��D$�=��<��̍��)Hu�ȕ��$�O�����5�t2�0�Z��B+<�a}Bm,?��DST�a�%)!dN6a*��q}���p� 7�O��$�|�⇓�?Q�}y�ͣ����&*�bԢ�$;�XU0��i��R0�'�1O�3�I{r]���W"0�$�Y�����Ix�K ��_v���fi ��\Z����D3?H��QÜe=����n�H�����S�Oڞ�[�ɸr����E��2	["OR�!Ɖ T��ջ�Ƥ\Eh��$�O��Dz�O�8ɄkM8��!�Ċ�!��PY�(s�����O�]u'�Q��D�O���O����?���Lz��@�D�h�6�ЌM�^X�'
���	�6L��Q�D�]m�p@��E�'5��p�i9��$�ߛ}Q�M�ë ]��'h�EI�H�az�����F��̓R)˔�y�i�d�ن�q~qE�*�M���i>�%��s�I�.�i��V!d�2e�I�j'pac�'Of�Q@���5��-Z�wh���'�����+�k*�%	8b7l��'D\����>p�X�ǫ�	x�y�';��r�����Vy��諤 Dy�<����R���r])�Tx�0�
/ z!�$��Xyce�ՐH�ǁ6w!��ʐ"b�X�)В�>Q�GM�!�� AQ���!#��a#o�v@�7"O!S׋�7Q#�!;�NԱ{�%�'"OV���.G5��퓱�ϠNӃ"O��*֧|p�9�G����ň�"Oܰ���gz�M��	�DD�=1�"O�&���v��U�p�5+�NL�"O���gLK�9�:9#QE�>��h0"O�-�ɚ�t�O��Z��"O@���@__±!�Ǖ�$����"O��H1���y6��7f�~u�$P�"OX�;7���᳢EďK�p@"O�CĜ�Y��K���23��a7"O����V,.��q����1Q�"O ��d�;2�v����8�V�zE"O��i�f��t� "U�{��9��"O칑`,G�Q��j y�ȚB"OZ�k�a�L�^���C�%?�� 5"O�	@fӯ-�I1�V">��@t"O$(��ا���q���c1��ڃ"OA�ee�5&�R 3t!])��7"O^�z���,�PC [7<�Y�"O��ȁhٮyg��`d��K����"O@�؄�K������r�~i0�"OdU�q�� ���k��8\��� w"O^���gWoL�=���K�a�NP�"O��G����%0���9�D؊$"Obx�0�"	FLh�^�b�FLC1"OV�����( � ��c�%/���d"Oj�3���?$"d�c@M��3�"OZ ��*j{�BE��C�yL���'.�4�� ��@IOW��	�'m|-pOۀ��)%�Ϙ!�$a*�'KZ����_NF@A#kX�ܴ�	�'��yY% �#�
ԏ^�Z�x�0
�'0����/!�"�PdխR�P+
�'��#Q.�v�Nu�a�L�U��'C�x���9���V��1W���'�rE�0(G4�x� �2�.�@�'�8uO�T��0OY�[�rq�
�'ȄU�qd�"=�Z�PB�Z~����'/�d{4.˴b����R�H� �*q�'u�-z��լ0�bq�O($�l �	�'�8	��O隰9��1Ѩ`j	�'��`	Ȗ� ����0m���';`�I��&&�l�S-��"~���y��9�� ~����*�zĆ�NҦ�pNI�qzU��˙��伆ȓ`N���ET�c�l���.�.+�ȓY�>�w���!\4՚�Z)Qqd��ȓL�&�Ak�$Ɲ
��P"z^|��ȓMN�y���yh��S�3Cl�ȓ^��Ī5  ��,��Ȅ0tфȓut��4ڢyI�㟊:�b���]z�"�CGg���bŭa��%��J�Q0)*v�kPe�)HZ��nT})��ҫj����犾b~ ��%6���I� LFI7��"x��d��O�}�%��,�«<p�4��ȓ=��9��,�&Q[�aj�A#C���ȓ~��Ѹ@��}Ƹ�8Sk��6�ȓI��0R4�$kEƕ�PkŞ�f�ȓy���C�T�D=H7��k�r%�ȓ1ڎi�D텔�x�1�.��#5����be �p����w:&��T�[��Ą�S�? b��G�S�����:/^�D+�"O��2�-O B,.ِ1�C�?R2��"O
��a�ӑ@�BtR�5�J|q�"O轚��L@8�-�@�0"����4"O��$�,YU�Q��"C�@��aH�"O���Q�׃K�RሴNk�PJp"Oty&�
�x�u!񍚮�nHW"O��Ra��{Ԛ�aQ�7RB����"O����C�s�	�q��O��y�W"OĽK$ }�H���ъ�A"O�@2΋��t���A�,�:�"O�8�E	�jSh���J������"O�!0q���.�&����`���C"O�䁲���8��ь��JŚ��"OV!�%.J�@v�Ecb�Q�š�"O�57�]��vj���aczhp�"O�p+���?OT����,bz���"O�t٧�LMn��6光GRf���"O��·G�c1`��^�)04�a"O�,e5�s�KX Xy^	�·�y"E\�[ظ1���?����4���yR��I�6IF��?A ph ��H(�y��jv���h�>�"�L�CrC�I p�Ќ���9]�b9�vb�N��B�	���	���<�b- �k��VݢB�>"��"e�ĸ+�����V?[�B�I�N	(��TGG�L`���O;Z�B��>]��8yu��
�*q�K�P�PC䉲(����s8 �0@a�dC��C�| ��o�
أ����	�C䉒7<y����_ۘ ��D��u���P�����^����E1'�n[����b	�"O|�"u��E�K�E	:-|�=��W�80YH<y�E;�gy� E�l��FD�;+G~$�fO���x� �Z$���$�)iX\ �J 4r�A�J� ̲���5|O�<c�Ɲ���k���H\��'�'�i���7��	�#h�O�)I��>z�v�[��kW�q�6"O�� ENYe�hѲkT�Q���>Ѧm�>z(8���o��V �h�&�S%@�A����Z��1C���r�TC�I7&�"%n�kʸ��c��6$�ua��[b��h��i�t�ю�^�g�b������<T����z9�C��:"��X�KG
�2b��Dh�5,\�E>t���%Qc6 �EG4LO�U����_z���vf��ҁ�a�'���Ї,��s��t:��/#m*]��Ń9�HD��fA:[ʀ�����5�yR�ʸ'�n	�G��Xuzhb����d&�`��%��2HVթ6�ٝ�������5�e��g�$�p���1�y�,�<�h�Ҡ�Į����D��H�qE�VM*N�l�ap�	�����I$�D�B�T�p���l@ 3�޵_D�BL�#���!x2�9�T�Qa�M5�m`~(�/þPL��+<O���'MZ˖m�S$Ίͼ�z��I�t�h,Y��^�x�j5�6♻>z���B�-N���kd�^�gF������x��E��V�����2иq��횹��^�sK`A��ޗ+f��y�ЃU����TQ�)V�9@ɽiޥKT�y"��|-)����U.�kR��#RHy��ꀢ��Z���fE��3N~Z�y��^_lpR�K��
�����$�x��N0]�����¥a�%�ׇm��`�9`.]��J�:�X��
�\/��X���;Gq�LH�/��ª����*�~2)Y�`�	��
�+{>��%A�u�޴����a�����"O�0P��C�_+Č�X�5�4{��d��DM��I�HŧO�~�|�b*�mh;�N6$HT`ۓ"�x�<YФE���@�J]�7,��� ��E�Z�ke�+t/�	�H���
9�8� "�
Ú<JUxB��< �}0�c#,Y�)�1�F<&V����'�&0���r��(���+W��A�Q���xE�p�?lOJ����(����S�? x��N�/_�H�����h�"O��j�N�zD�DKf���L�1��T�!�̍���$�'H�0�G�n�@I�Įʍ��ȆȓW�`Ҳ�W�:o�Q�a�[�)��IxAA��h�����	i���B�уS�!�dL
�(!���D0G>XK���N�!�߫ko�2bD��w �u��b[!�!�dB�s�t9��ɀ"F�L��� R�l�!�$�D�fp-���������!�DH
$)��d۶��3�
 �!��� �6��B'n�Z���/�!��-�>p#�T�S	��u�� �!�*k�:��T�j`�R�#�l!�q��8a��� M��b\�d|!�Ԉ2OX��$���I؜��0aHa!�$E�$x*h�n�d�h=���@�.!��r��Ոqh�=�4e[1'GPp!�K�>�\���_&ZXf��7eg!���4FQ �E�k8ba�u�ʍ_6!�*�{�I�/�
X��E�(�!���Y�d�I�L��&9�b�]�S.!�D]��
Ź�oT%=�.��U�I%�!�K)j�4�!�B�=(E�5噠O!��.g)���b�ܕ\�Y�3��3?�!�D%g�!���R�}�Ω�p�թI�!�䀈qbNȱ�����y�i�? �!�$F�v�d���د����э_2!��1>�@��65�d��q��!�!�#T"��R��9���Lh�<!�����"�ɣ`&T5cW��j�<��%Qо9Ӕ�P)�W�RZf�ȓ=_l��f���B�"\+Aˊ.\D�,�ȓ���j DF5C��'��E�Ն�C�j$���Q�=�ը�bBOhĘ�ȓ"#�i�+Z-*�xi��v6vq�ȓ]ǄxD��:�Rg��+/+\P��w�4Y�QN�(Hq��P�H&��o�h�������ˬ5	�݇��̑geE$.l��*�3��X��,W𰠕a�
T+\��w/�H�<͇�v<L03��!�����N�+(����ȓI�,��jF�>'��Z��&\هȓ>��+��� ��ʶ��&y��H��y���S�*�/K|ت�&��uuI�ȓ`d8�gό5L�4!��_�����jH22,9`��i����� <�P�ȓb�u���@��i��'*@p]�ȓ�|%��rl���]����ȓ[$0�R�с(?�)E$߽*��ȓ�M���0~��@��v�P��ȓ!6B��d���K��`��⅊!̈́ȓq��msQ��"1�6yFiX����@TAp3�U#�0�*�-��Kz̅�"iҀ�	)`L��J."�����DUZ��V-G�
<��
+m �ȓ������B�Ze���&�.���?�zA��[�E���c�%T�,@���b��ǰO��dY�$#M6 �ȓ*b�`�fרA�$Xaʧ@u�̅��l�jd!��U轻6��-G�����	\XX��G�()��=Z���N��\����y�,��v�´0%��?lf�Y�/��yBȍ?Imx$�do�<4 ���N��y©Θa���@C΅z�.�z�֥�y
� V��m��wl�R�8!"O�I)�M�2���@N�E=��+p"O^U奜�b���ԇ��0�9#�"O�$
��N	(��q�3'U�2X�"OrD��$�9�4�`E�<3O�,��"O����E^����X�� "O@���+o��{��J�\ZT��"O���Uߤy�fiCbYY�ly0"O$蚂"��a%zh����-�T��"O�4��6�f�P�	
J�f�A"O6��PMG�GOjiPHU=�&���"O�PH��D�p��FS?&�ݠ"O�ѭ��_e�����-{vVأ�"O�P!u�[�F)8d#��)�jpx�"Oj11a�
�V�	 ��Js\��0�"O� �e	��qc�KvH���"OX=�B�#
��E���ٯE��i�"O漈�	E�*Vx�32�fy�"O^)1�"sXՃr&%Px���"Oz�ˡ˃�)Md�R���->^���"O�	����p������N#6���"O� ��n=h�Qb4�ܻ-�$;6"O��t�y*�o�,S ���"O&qu��V�2��`��� ��K�<�#��4b%2u�c�Q6n�A@M�E�<ir��8\eԌ��gG�	vV�H�O�A�<хcĺT 4[N��s�ND��|�<aȗc���2�M?����j[n�<��ǘa��#t(4`s���tɃ~�<�SM�_d��N��[y�A�f͚P�<9��Ç%�t� .S�v�,�
�%M�<��">^(q0�k�0�` R�<��/_-O�F|G�`d`ip�f�F�<Avhت<�^�`QB u��!��@@�<��Gޥ!L|+�T5W�ąI��UR�<i�	Q�4���H
p����,L�<)g��6:Iԩ`!��G:ȕ���J�<�qF��@��$L�|>RD��RF�<!��Y�mh��bL� t:ָi4(GD�<٣�� ���)�EW5�R�頮W[�<a��ܦc#VЩpg�9.�� �sJMo�<�����c�y�e4-�p�d�Ng�<��2k�d�;t�W1_+�dR'�H}�<��;(�u;�hI#"	�s��d�<�V���w�d�2�&y�L�)"Hh�<I�l�9�Pe�6�ی?oF%" �`�<����)'�%+r�Y-�5S�TT�<	��6S��PфH�@��Ѫ�)FG�<ѐH�+m��HO,Sr��R�z�<!�C�0c�����+`ߔ���L�<��)L���|�&K�x<��z`�J�<q��M�B�}���D�+,�I��WI�<��A�_�\�K�,�_5R�!�C�<	&�<�v��BT�N�(���L�<��.��\YG���v�r&Äz�<�"�?M���p��ݑ&�$c�'�n�<ql]�
�^��6P.�RQ��e�<�����$$@;��!��Ŧ�`�<�c�Q�G��!iR�X9m%J4� H�H�<���<���*R�t.��p@'�G�<�G&X�%�j���ǎK�*��tGLC�<�SȎ��eB���\:�����B�<A�A�#��`�>M4��h���<����qc�QEGZ1E�X�����x�<� $�{�	�dy��v+F.UD���"O�� kJ�l<��Q��*0G��"O�� V���z�H�?����"O�h�I��is���R��50��a�"OⰑ��R�yਘ��-�z樈�D"O� �,��
��  @�{ǒ���"O�4bv�F�[�z\�4.�B� �R0"OD�tl��_[���R�="n
C�"O�T��BS�T�I�t!�!~�]
6"O&]�a"��<�jÆ`кCp|	k�"O��S&���D^N�)!�� =���"O&�B�/�b�H�nۼ*� �� "O�h�^%x'p}T@�C
y�q"Oj��2!ޠP�
��2��7�zu�2"O�}�bC+4d�B�ʧN����"ONi1���=�.�g�ۊX��as"O��s!�@,c�Ty
Y�8��Ԉ��y�-��>0T����u�@�8g�N��y�lK�#��X&��o|<�;�i�y�a1N$M�YbB�P)�N͝�yRE??THrƀ�.^I��v��&�yG�fqkl��I���F�"�y#�;o�8AaD׳Q������y��
;77��(b��C��Ͳ%m�y�#ܴnDb�Cf��1;����yRd��_� �R�hc���B�e���yR�b2ء*ͼCp,%(W�'�y2�[2A�D��ˈ-6����+4�yBȵe�|�sd�!�F�����yB��O��Yd��ô���L֐�yR��76���	�i�%�|�1���y��1]MЌ#.�h�x(T�"�y��SA��A#��|Υ#`�4�y�%���K� g�����X"<�x��OSr �ҩ�yz�u(b�^?1(�ȓ\m&�F�?=��L�%H:D�"���D��L��+͊6Ґ!p��-�l�J���s���`Ԣ_�=@� �D��69D�x�, ~5����#.�ǆ6D��XFa�4��%�E�����ѧ3D���lZ'D�LpA4NZT�5)��<D�0�4��>�>Ȱ����"� ���7D� �q�_�"Z�X8$C֝
��)$b"D��c�i� &m2i��NT� ��	0�L!D�H5l2<Xıg`�ܦ���#D�0*��@/C���Q*�n��Y��>D�����)x��0�Ƒ|B�w��R�'�Q?���M�:�>� �!W?{u�)�&D�0[U���4�G+փ��Y�'1ғ�hO�ӹ;�p}:f9FQ-ad�Z	1B�B�	Ov�P�`f��ͨ���U<Ǣ6�!�S��M{a�N�5�@Ҍ�73���AN�<ٷ*��Fs�x�G�X���	�"GU?AP�'-v�B�+�S��0��3�
듋���D�7##�E�z�B�I�p�����[U�E����1:H��<A`�|�g��3B������ Iz�Rl�<��E48V>��'Iδ"4�yShf�<��/^�mN,q�7�O/	<&���^�<F�>4�mP���/�Խjf�t�<q"��
����עV3*�h���J�<AP
��v��M����#����A�<���5J�4H��;x�9�'(�b�<��_ �`߂e�@s�<� ��6)}�zu)��P�j "O�u)W�Xu֩Aǭϸm�pI "O�@��Ȑ?5}j��g��2Wf�"OT��
6o:i��K�1MލP"O� �0���n<\ @nپ(*.H��"OxQQ��������,]�,�X:�"O�	�U	0uG*�I�AD3�Q�"O�٘�b� [�A�ኄ�G^�s"ODeI0�/=��!�UQ�qS�"O�L�WƖ.1�p�1b�СX,��!�"O���� ��`,���J ��j�"O�i`�*\3&���uJ�K��,�T"O��Y ��<.���R�A�.t�"O}i���rߜD���I��l��"Oԁ�!��m��;��ܵm�H��W"O��z0`ƶdzX����+먠3s"OP S��掁��&�-��)�`"O@�P��4Z���f ��j�"O������p�Q��E�V����"OZ\85H؀D�9�t$���"O��8�菕�>Xz7㓈r�H��"O:mvN�ti�����o�%h�"O0�.�2��b�+�/60����"O�Z!ϟ�N ��u��'D�I�"O��hW	It�����A/m�7"O�l���W��b�1����kB!�D]���j�e��0�P+�!u !��	�^<Tâ�5^�Q��K�"!�D� [A��{���aE�p�$�B!��^��9�5�F�$�<�ط⎎>!��	ِ�ҠM����rcPV!򄌔"��eA��.� �!`�Ƌ:!�d�k">��`P�>-�
�� o�!��ކ�J�bk]6x1��cm�0A!��$}��Q�W��{.�]��MTGK!�\$b�z� 0��C-�=3�m\t�!�^q�������:R� b⋘��!�D�&RH9@E�;[�ĭY����1�!�$Ź�ڨ��Zsb��%K�j�!��2;\�� AE�h� 8Tj��/�!�dX0P7��ss�^{g� `$/;�!�D�"��|PV�H�g��`P�Ļ3�!������ ȍ�g3�}��f�0{�!�d�
���:d�d|�D�!!!�	S���@�I���&��W!��^[�i�����.��d���:�!�DԌ�h�5�ɩG�XfY�R�!��
 ��
):-<U!��`!�D�
�z2�C�X58ajUL�!�G/�yT���AB�q��[�!��B^�"(�O��r�P�֌K;)�!��s��@�C[��TصK�8J�!��ڏ�(��W��k��9kq��j�!�ŲUCP1��dW�$X�r&�	O!�D�&�ʼ�G@�Tu>��p��9T!�D;[#���a
'u4ybԤB��!��Mڀ|��n�3fl6�8�d ��!��Y�X,,�C�8U|bU���WyH!��Ѵ(�Uzs!N�:�`�1C�E=!�Dθd�X��+D/��iA��,%!򤀕x�6��&l��}�BI(�N	8->!���-m��@h�$Y�X6T��
*;!�N�E��� �ˈ@���4�ӝ2!�dȤp <�@��7�&��Q�*<�!�����! :  T   �
  �  *  �!  �(  �1  �9  ;@  }F  �M  !V  ^  hd  �j  �p  .w  p}  ǃ  �  �   `� u�	����Zv)C�'ll\�0"Ez+�'H�Dl�|��00O�1"�'"dWJ�� �ެ`H���exV�O v�ll�6hFf����u�w�%1Q�^�?Y"�CP�?�3u�?ꅬ(��LqQmH4�P�WT��Ɂ�f��� �/IDם�W��)����$(#��.�t��ÝI��1�Af��U�z��O�?� �<H�X5�A��N��V	�8D'B�'��'��bO�:S�DSS�G�h��* bv��'Ղ926bx����?�����?Y�Ɲ������U����j��?9���?Q���?ad���?y�[ߟ͓�*�0CiB�P�A�G��z�c�&��?њ'�寏͎Ј��̤vJ{eF�>)��D��l�rc�	���\)l��4j�!`�0�7*OrH�D�O����O��d�O0���O��'�yW�A5�@�1*�+v��KB���?i�i�t7mئ��ݴ�?ap�i�0,0�m�l�i��O�X
c7���`1�ݬ/��i�%�l�'�d�9�(�[�OF�� 0����̢�,L�H�tT�%��~�zD�����!?�P��iN`7�V�����?ŘP���~��piE�YBd@*ũ��|� �JD��M����<�4�Q�7jJ��ӊ|��� ��Rq0�fam��lZ�bOą2��*f�D!`4L�_A�t��e\��}��o��M�i��6-�8u���7
�c4�!�,��\;pƙ?/x�ҫ�%-.lA��dS�g܁���-�Z�n���M�iN �qA �^�y�E\�'���u��4��#t��t��< )�)7a�xj�`LW^��n��u�R�$QId�=�W��)A��0�C��\��D+�	џ��IP۪@�ٴ��iE�F_��e�Z��0�$�iJ�T�`�IП�̧)����I�|�xQe�M�B�� aڐ ���޴U�ݰ�C��0<ɔG/��E�o���Ll�/)�)KvM�4Z����vB�3~�Ԅ�I�j��$�O��'IR�
�b�18BP�#"ɞ��f�(���?�����O-�dT�]��a����,<!h�o{��NwӢ��4U�vI�qt8���q	�Ц�'/�@�"�n��r���O4�'1��]��'|t����JǞQ3$��� ?&�E��?�f_4�?i*O��d�|�O|l�t�ԖV-���0G	)YnP�A��`zb�+;t�e����G�4l���)� ��Q��YR�����i��U��,&���?��'bv|աW蔿k^�ᑧ� K����Iퟔ�	R~"+Լv�NI�n˧3�v����Î�hO��D�_}bV��'d��ф�R;Vd�4�Jȹ[D�I�2����?��g�'�18�G����j�-�Ez���'6���HWD���p�Ы�2�+�'���� A���Q&�u���
�'ƴrN�W�`Yq�
�l��
�'�Z��G��'����0�C�<^.T��'6(h�fQ���r��:L�2�*+O����'iN%����.娤Z�́2���
�'��]���*xع��@�-+j<��
�'?�e�oC��ٛ%G�&���(
�'�zT{���R)���&W�%�(��
�'ؼ١�o��gG��j�#���)ϓt��u#�i0�'��y�3�Э���!�""$��E�'����9��'�"*�$���頶iU���K���ej4�?R�%0�Ɯ&"4�QJQ�7O|-k��8&����BJ�����#��*.#45�2���*�kE�ax�����?���9#���'%�P�6��zV6���J�ڵ5Y�0��c�S�O��� K�eeY�D��}��`�yRU�$F�d�yӘ!K� 8OZ�X�g䔎d4��g�M�=&���$v �?y��$���vK7�V��TJۉ^�Y�
�'gh,�1F�*���0��8�<r�'h�Yٴi��QP R��H��A��'�R��7�C�.͔ՙ���1��'�DX�C��i�չ5O��Sj�)�'l������F���·O*��i�'p�q�O
"�'t�Q�h���]2 ip���?Rbp���Ʉ_�ĽI޴:���](hjh�1S>mp�r$��
����@�p����D$/gꈁ�/ӂ���W�N.e��0�T��V�
��QA`���3�8�����+�`Dݴ;F�I�D^��?��OF�d�ON���ȉP;��i@n;Q�:���%"<O`��?�w��-'��%Z7��G��	Z�`@yb�~�&$nZ`�i>��Sny�җ+n�E��g���be�����O���銙HzR�'R�'f��]ܟ<�	�|B��� q��@�`�O)�Dٵ'��.��I�U���
�	F�C)�=��EKB1��C���m\j�C�E3�Oı��	�7 T
E+%ш+�2\�eϟ*aD��2�O���
�<NY��E���\~L��q"Ov��q̄�+iJ-a�vu�|�#w��OFD�����'1��I��/"��{Ц�4_�b���D�O~�D�O�����/��4)b˛),i��)� �y�a�WO�3��I�&���ZA�'Hp9KQ�\�l���`[��y�K_su����;x�� ��0<鐨�ןL�۴�?��q�:�����d�L@A���+
(
����?���?���䧯�'��po��*���)�J�p� 	��oq�$52&���-1#�4� ���?�/OdL��Ħ=��ɟX�OBq��'`�)$H/+���x���
 �b�����D�Ud�ן��<���	�)(����տTBȃ�苉.D��\��Ex����,$B��Џ���
R��=���!<��M�)�'���:���HR�C�=���ȓ;t�Lx�������� �]҉F�*ڧD
:�A+[D��@�֒-C��B�4�� o�Q���?i��?�(OE8�Дe�����1]8Fd9��M�g$��� t�Pr��ȏ�b>c�X2L��Y�J�#9^���҈����(r�p3�'I	
v�c>c�Аt啲J#XE�Um<l���JBͦ���럼���Z����nyR�'���'�졊i&�f�Z0 �tȲ��#"OFQ�`L������,�����W�L��������Jy�˛C�B�s�˕�@0��	��1uDa�d�߲1��'�R�'�@�ǟT���|��>�H$#(]tQxM6Mʺ�`�h�+2� ]hg�Q�ay�#��dVh���'_Q�i@QG2��I� �R
[~�CY�$L��DF�&��$��m�;`*
��ܥ>%�#B�'�Z6��O��$�O4���O�D�O^�LNX�`����l�pP��K:v���d���(AJ��S�p�[�ƄC���&�Lx�OV�Q4�1�P�i��'��·o�5Vpt�rBϏ�5�"��	۟��pH������|�e�ҟ��<�⧖�?(��z�lZ$J
f|�@~��82�9�9$<�a恂�YPnE�/��ć�	1�dF�I�¨H���'��Lr�d|�C��y5:}��JP;B�В��	P���$��lb6g2u�@Aס�1jpԠ�E$�D��M`�l�˟(�I`� א,.�B^:A�8�p�C�ia��he�'e�x B�'0�Iȟ����Br�i{��Ԙ}�B8�G�&;n���bI��B�w ,�bm���h���v>S��h6��
%����Ѭ�O�nZ���OK��4�X���-F�H,�rE�5�v���'_��'���1~@����5`�ԬB�d/|<�=i��oI��Zy�2���&($�tsC�8)eޝ �j����O$��)$�� ��Ov���O��db���BBN�.k�I2�Y�L�Ã�,l.��!�Q��)s�d��G@☕O�$� c�Cb~�UXg��6��� ��ʩF������OV�=iJߖr�jb>�PPM2?�Ne �|�� �+G� �3F D�pSݴ�?)�h$�?ى�,OF��D�.@�Xk��M�a�]�+��hO��=i��@������!���A6t���9��?�eT���'����T�'q($h��.AS�t�%%LM�R!���?)���?A�%��n�O��d�O4y a�įJZ��s�ћu�bm��c�8x�M���&G�98T�ox�H��&45yB�H5�խmVMI�KΗ170�Z� �mc�Y{ef���.� 0>�^
��bD.5��y0��եTZ�͛'/D⟼��?�M�������O�㟼����v�IQ%L!W����7kꟐE{B�'E��Ę�F,��ZU���s��9m�;E��	�xh�4�?�/O�嘖��m���<y@n��n�,-2�gǿCW�P� ���L�'�R�'�2�ѷ{� h�B�ԇ4�d�C>OR�9%a�1�ز�-�6%C�S��'PL���R�]�$�q�1�y�/B�Z2-��I�k:�Y���0<��i�����4�?Q��X4�r�j�� �X��$ߴw�^�����?����?i���'��'�
ȹG,��
�ح��ɧl�6����=��	�+�HM:b(+-�v�v���?).OV}��k���9�IğH�O��eB�'Z����Ќb��kUd͇i�`}z��'��F�o"��t��>q�����|r�'B/Jm`����[2S�����]���D�)Dx�( Bء*�����/ 70Ӳ�j���灢o�x�ҷ��&��Y9��:��$S��*mӔ�mZ���G�DFA(l#�QY�ޔ�B�JS��5�䓘?	��hO�I�*r]0��pJS/@��q�W�D�=dџ�zܴ����|2�ġIL&|`�F�v,x�)O8L7"��Y�O���	X�L�K��&P���P�,5|B���pH��ŒC��U�P��v�B�	,"�PX����&ZfS�͋�ϒB�	�t��@h'��<�`t��$�K�B�I�b����m�����H�k�B�	%#�i�3��).z���Y�e*�ʓA�ZE��r=rpr�W��Ӈ&�"\�fB�)� �mzV�W� ���۱�N�"YX͊b"Ob�ŧS;�|���C����"O�1����x����O1!���2"O�8�p��*5��5��G֦��t�')X|3�'/v0f`�4Fq ��5��0�'!�-�.]AuD��0I@�dA�0�'E� ��
]�Y�<h )C	%�uc�'^�
%�U;���h��K�z�	�'��!A��'L����R�Vu����'�tQp��ɸJ����"��{���ɋ��Л"�Q?���Ĥo���)���S�D���.D�k�A���șh��ɔ��I*�@!D���f'Uy1M�!����c�*D��iB�K�$�}p��y�P��<D�����ߦFd��e�:)t���;D�Ģ���Y�ֵs�Ƒ+@�Ě��O��b��)�'C��4"�]d;r�YC�
2u����'4^5b�eV0u2��i�HK�Cຼ��'�=�C"[2�H�6�W3e���s�'�p�1�N# �`��d��'�pD�FOP��#E��\��M	�'��<�p�_�L2H@ ��O�T��M�-O�4���'�\��я	�+��L�bƎ�H#�(*�'}$��K� �t�"r�V�Q�X�)�'������X��t̡V�Mad����'�4�ň��8G�a� fP�S���C�'j6�t�E"i�(�� +A�>���>>�L��.1A�.D.�Áh��h��$�ȓY��2Ĉț0bj�3@�.@��8��ɪ�s�ld!b$k���bfR���9�*yÅ�)�`p����?��ȓՎY���5/s�*�%�/fצ��ȓ\�������W�1�E��(��E{�Ȉ�����q�EY^��ᗣ̕4fh�"O �p�}�4=����6 �mz3"O�`�FO��{� �1a`S�l~��a"O�	k�iȩfWT��ėdc�[V"Oj��5E߸���� �$�ԑV"O^e�����i�Ɇ&�-D����'ԤT����ӊs"䫢�N�Q�T�1���ΐ�ȓud�(��ϯlR����ݰ���ȓk�b���B�r�Ѫ�AҮL욄��.3���`'\�(�\�²ɪ,���2��Sg��Cb�4BwC��T5p��F#0�"3�ηN�P`�˟����' �DP�5�JA��M�=T���+���-!�
�ȓ��4��GM�,+����C���+N1S%��9i����(��>�ܨ�ȓn8r���iΜFh s�$5*�ȓ.��i����}���ƫM�J�z݅��5R��	��|���7:9vIے�0PԺB�!M���%��D�j�I��ƌrTzB�	Ff��(Tყm�>�Y$WH@B��	���QL�w����B�(p�C�ɯt�
|�6a���1+'E�q�C�y�䬢���?S$��*�/�7ej�=iԮAT�O#ԍr�kM,Ru�$�A$Ιldj@��'j�m"�Z"k{@)9a�Q�d� B
�'�����RUm����L��T��P��'�4@V)�0%�X�1�F�T*�� �'��f�ʖf�H�jBn��yR���'��,i��"������ِr�dH��Y�MGx�����<��1y�,]�fYr���f��B�ɏ\P\ɥ�Vc�xXi�{��B�)� Hu矂BC�<���Iqr�"O>y:��!R�"��O�.@<�3"O��4L��ZĈ�U��RT"O�p�\SPfd�!�IV,���X��bff$�OԬ��5���	�#�����"O�P�@������
p��U;4��"O�)��`� &����` F�6�h�s�"ON${���<u^�)��.Џ�<�Ku"O31�	Ūm�u��w�p��'a����'M(	Rb�YmH�����2=�m�'�dU@��٧���s�����T{�'^ΙZ�K$7���a2D@~�h<+�'@��g×�T�T�Ȕ�Z!pn���'�*�:t�1�61!N�1�	��'�NQV�Թ$ἅ�f�7b�vU`��dR,�Q?��� ��懙#VI���-D������ܦ�ӵ�Z"t�T��!0D�@I�T$�&�aB���M�p��9D�Z�d�8G��r/Җ=�H���5D���&��y�y��O�EA�5D�<�W΀�\�xi(�L�n���SD��O��2��)�'Pҭ�6ꐦ4��IʔN˵F��A�'KYSE��"8�}���	rzJ=��'�h����v�����:z��'��1��G�8}#T�#Ы@:&6$��'��}��Fq���C��2Ȁ�{�'�.4�K�
А��+� �-Oֽ�E�'(B}Y�JоA���(L�
��
�'�f2�ꂽwo�H�u�_\�Y�']���Ax�>ͩHٛi`-{�'6 PC*F�7x�S��
�񼙃�'?�q��ͤ�ꈲ��X�
�L!�u�f���j��	���'\�v�a ��\,&(�ȓ>�f܃ƫM�g�n���f�l���\oN�{1.�d�[� �0j\5�ȓt�(d�v+:i�u�s�W�n�҅��8`By��#g����׈u��)�ȓ:4���ϮBE���܄��yD{NѲ���ܥ��%�Y��t���g��m)�"O������$n�� �g W��8�:�"O0Hs5��6b�V����]	I�,$ˇ"O.A+�i��y��m��-��ֹ�"OX9
uL�bڮ�!F�	�q�>��7"O�8kF�
rx�1L�;H�bt�%�'��UZ����(PȐzɀ�6�Ԑ"����b�l>D�h��o��St𓴋�/&Hp�ar�0D�\[�&��}a���V�]+|�v*D�P��X�S�X-�F���9]8�7*D�l�Tf�AUV�N L��a%D����81�D;V����@K�ϸ<���z8�pH��
�M`��� ,޵�(<D�$�%����6���_6`�)�Q�:D�Ty��$=b��xAL[�zu"�,,D�TpB%7i��4"�,)��l��i+D�hFa_(!��\��B�V��g	=�O�mB��O�A��H�P���ˀ���h���H3"OF�%�F>t�H3+�50���k�"ORA)5�@/Q�|�@E��a�D��"O�y�"Z�Y
�Q3ys\Lj�"OLuCtD�m�VA��&["	^��"O�QAV����YAFG�:�~�X��I��n�~J���{�����і'J� qU��]�<��JӢ0���я��g�y[�I�Y�<��H+\����D�ާ3�
�"5ŚS�<� ��P��Ar�8�� �|��Qy"O^�
P�Ϡh���(A}����G"OƵ
��E�b^���R�����\���'Ǧ�щ���<�Bh�'lE)v۬�z��F�|.��ȓCF �a(�s�h#���}xޔ��?s��"P���,w����
Xq�n9�ȓ^�ݙT�H"V�~��Ŏ#G��@��s/R��2�_4*��s�&_R���A�������8�d#����'�����yJ"`p"є,�L!Ǚ� �P̄�v$BI�����(A	1�	�'f�P�ȓňT�(w��	����7Q��ȓV$��Qh�v�̍�����U��F}����D=:|3$I7H�p̄���7&��	�81�x�cD��dp�� `M.�B�I���@5���%MC1Q,�q�"O��c`N�wZҥXg F4K 0��"OD��(8-dys�.�h��qC2"O�<z�,B�h�H�;&E�$��4�"O��B"Ϛ60r�!�aҿJ���˃�ɩN@n�~�D�W�Zẅӣ�ǂ��=�7�I�<I!aÚ"��yaD��9k�*5�!�n�<a&�؎7?rtP� �6X�|�����o�<q�g� kT��ѯZ9LubՂ�Hh�<9����f[��+�J2J4���Ą~�<y�.%0͚Sv�M*������!�S�O^pX(E�j��U��� z���"O��E)�#�N`���#��|x�"O4�*���<�� ��;��K�"O��a˟��BثE�݃E�H��%"O��!pmD)I�����+;㢰��O�=`�ĩ916T��J-W�h\��*�O��'P"� �&m�Gb���R��]ß��6���c�a��e���
FF��s�X|��S���I�H��5�r�H�hD�V�npk�@ �3_\�A���v�*A@��$O��dM��MT��Q����й}0μ�Fm�&���뤊�:�2�:��^#`���f�q�L}Yϔ7T�Q�d[��O �mZ5��'z��I[r�S`�L�m�$�9�'sa~�"�b�
0��f$wl1�����>�s\�8�G W6sqnq�`���&q�i���'�ɈM���?��g?�����}` �Atn�"���D\Y�<����PeJ��1	�2�(h��$�T�<�� �"<&�c�`�o�!!��YO�<�b��=鮴��Vx�X��Q�U�<�b;3��-�[��`p��w�B��ȓ!Fp�7�M�E$���'�.(V���5�;�h��D�EOMQT�+_@⭒U�
4
�!򄝟2X^T��aJ�y7b�P�����!�	���R�c)��b��$�!��L�����p�T�X�o^�mY!�d
Z�ⵡWnƤ1��8UN^�eP!򤋷R�X��o�PQx�C=P4"�V:�p?ɡ.VhF��KF^�x2��H�JD�<9�M�J̈��/P�f��)����<���A�b����e�$R��k%HS�<�B����\RF\�8�0yveV�<	���&1��Q����2����aBT��и��0}r�Iu� G��a�"�QV� ��y�H�+8��9Yt��1�.�k�<�)�?d7J�����Ts~h�#��<��X�T�HVJK�1�* �5��}�<�v
��\2H����*ܦ��a��n�<y�쓣&2�b$��R�"��Gb�P���qExJ?�t,����h��'��1[�%D�h{�K��j�ׄ4����9D��i'��9��Ԣb��ݑ(7D�� $�ц�ܛG��Xy��޳��(��"O���Y�7���K�7bc0�I�"O���ax�F%!���|v���H��O�}�@�^)StG��O��)z��W*c�Y�ȓ<wP|r�B���Ԩ�2� /�D��
�Q��D�f$�]�'� LBP�ȓ7��j� 'b����M"#~P��a��l����Ut��PeO�Xx.a�ȓJ��I䈌�[�uB� ם �����#;q6��dӏzj�C3c�%�	QQl4j!�D^|�r��r!�j$���ڥ{d!���==�(�b+O,�Z�je�=D�!�D[�����D?f�>�3��8!�Td�aJ5�_���i��wџ�����M����?Q�O�.9s5�כ]��p��9b~h�:�+C�����?!��K����1��oЦD[r��>�'5�Ҝ+@�V�R���c4.���B�E|�B]�AtQ�3��M��(�1�gۆq\�:"��5����ɤ4&����K��4
Ԍ!��R	+&��[�!'[Įф�PЄ��B#�b$��*:t�'ўʧ+���6��:d�ڹ_��m�+��$,��?�����|�����ҕ 날*�џ��9a����8џ�����*�¨� �
�#��%�Cv��O�|�1�x�χȟL�O����7�@V9���g��p���2�Op|�t��T�O�s�����ex��� ��#T�*\���'B�'|<�J��H|ʄ��Xwn�g�� � �ifl��Nh��'��	\��y�"ȳ����p
V�KAtX�B/8@f�8�N��xN��z��=}��~��)� Snrd@�B/b~��KI����8}r�֒��P:"��K�}A�DA<v(v\�P��Od�$�>� �>�fAm�����y�'�:$<��',^�Q���Q�ͧ<!4K_O�$�E�O}�G�[k-.5z��9V2�в!���l3aI.}*��]�7��	�g3<0� D�:���.�*dpI&ÃCy�o�;q���'
ؤD�D᏿7�8x`c�4r����RK��?i�����Oܟ�&?���]�|���~mxr�&�����:�D��?�sg�?
6d	B��m~D��D+�b�<A�`��P� ��3H�}GC�/
Ԧ�I埸�'T��'��C�\cf��� �N�d�<���%�\����4�?9(Oh��V���'���Ґ������
҆(��9�4�X��M�,O4�İ<AL~,O�p��գ��Hz�$Q�q$�S�<�`��lW�1{���Drؑ�qkP�<���̫A`$��7=.]	��g�<f�ِ?�%SC��7�D�ŉ�Z�<	$�M*�r��  J�`n�Y�Q�Z�<�d��ZS�Y�)��<�[煊K�<��&�k�� 3� 'Nڕ��"�}�<�����8aŅ�!�`����|�<�'�P #L:r�[�l��}#x�ȓ#��x@Ъ�;d����%�@?$�Gx�O�G=��H���M-Fj*��0���]��Q'���^�!�$�3G�9!�<3k�AZ��@!e��O��+`ș�#��8W'���a7����y�ri�kFܴbk,2���b��3U��ӧFO.�>��3�N�$�R�2V�$G#�m6g0(��-i�61�$@B�N�Lјe���:\ִ���B��؊�MS�0\H�r��q��Ʊa��U����	 �4g\u��v�i]��q��Ŏd*�0p�4%D@sե�O��d5����aFh�|��"Y���& �f!	��Y8ԢԘxb�_ )�<�)FKܝ1�R��G���J�!�2̃c�ȅ���'i+E{����	��O�x��'3�7-�ɦ9��`�'-;�x)�T*5��!9��ٗD�$��=�����<q��=kfHx�^#E��ÕM�s8��c��D���Z��@���&=y2��H >Mp�����ß��K޲pZ�������	��lx������Ȉ����3�����'{1��R�ɔ�J��j�'!���Łv̧q�ɂU<���1)[�5	޽A��Tʘ�1�e�(�p�(����j�)����fHN$^>%;�����ygd�c^vx��ֹ"����;}F։oڸ�M��)d����S�gy�i����
.w� P��ǈ:��u�G`,$�x ��R�,Ϧ�@l���H%<}�n'ғ��>�ׇՉ!�v��U���s�P�`�!U7~�Ρ8  I[���':b�'`rם�D��֟P�U�[<�㥎�t��k��:1�~u��,�^z@dO�%��<��� ��&�1�Љ��
*5�����ʮN ƜZQ��{�F { �9^�DLG|�)@;`(*�a�K	,��q��U�������?���iLrP��	h�N���0%ʃ"-����]�ح���hO����O�OrI��*��l`S ,��ud��R&�Dyb�'](6��O��<p��r�i��i���ԫ�/`N��6Ȗ����ɨ�?)���Tm����?q���R�������i��P#�J�5pvdbr���T7��Q��'��TQ���jݼ��fM]^�I��Y&f�5`t��#T0���1,O� k �'@f6��@?���L�v���2�X�����E�b�d�On��$�;*�hy�����L9iбkH����I�t�'Iў擖UŞ��� �l�;����}��ߟЖ'�yvaTdB���?y��7�<��4}kre0�#�95���ħ]X˃>�?���"����&����Λv*���'�u(��O�B�ոv�ɐ(Z��'��R
�qj�r�Gں8l�aD��LX;]��H�A���e�b��!ʨ�ē6�N���؟�G�t�i���į-,ԥ��b�$�8A�+1$��i��]�����G^�A��	;��&O�Ey�M7aꂤI ӎ"gHX��FTZ�poП�	П�Q�!ȱ[?�A������	ܟ��ܹ&��%�č޹*`�"�ЭVʎ%Z����	ڲ��}�yF�y�'Jq�I!n��#��e�R���,̷zu�e�r�B�� 9s	 j����!0��'��]3y7,�PW+���#oܚQ���	A~r'�8�?�'�HOB�a3���l@
U��b��\�0ke"O�Z�`���V)��B�k�u3>���i>��	c}��V�̉��	�,e�2� �`�9���S�$���OF���Oލ���?�����ԁ�l���B�B�@m(��*Q� ������T�3/`�k��{��$#f��
Q��#�L�����&�Q;�t���%b�<P�'G����oD�W��嘐�A�4.H��eA9�?��i�7�-��9�O�h����W!;F
Jp��B�t��'����[b��8Ӌ��-���P�{��>i�yR�~��� 6膕��#ת;����օ�ZyB�)�'W4LaR���k�XD:�B5$)�O��d�4d�HQц�U�0ih�)�:#!򤓸k7��+�JYh���!��5!�$>�h��<i `���3-�!��TXH:���,�p<؀�Z%m!�dێ9�E+� �2[N6%9we�ng!�dɮz����ϟ�f5~a��Mq[!�dїVa�q�P�Ѩ$$\��7�I�!��=\Ɖ:�é�@��Ā&�!�DT"�lh�s�PL�0� �E�Q�!�\�`����c�
v�t0RWB��!��ΩR����'G�~>M�F���!��*/���Y�tډɴ�/&�!򄇉,|���l�0bh-+��Ê:�!���G�ҭP�)ۼN"�Lks픜,�!�ܩK &% pJ"_�4��b	�!�d� c8�� C�u�n���*�!�D�Z��ڣ�Z�5?lL��
��U�!��	"(��$$��b+ 	�4��r!��,S$��{E��^ɚ$�)Z��!��*9`haS��e�nx3�%Gi�!�D& ���(�%��i��݌xe!�D_�n����S >���P��\(���$.�L��M�?.���`%���yBNB�`�y�aݨ:�(0�M�5�y�l�Iy.��c	J�7,�pkËY��y�����Xq����(v��	���yR^��Aa�b�	���y��MR8�u�"a�.����H\�ybbCh@����G1�t۵�B1�yKK�o��Q�/S�[:�!����y�em��I�TZ�[����h���y��Ѥ}�P��&̒�^9"�����=�y"�ǒC�d��� Ir�t��I\&�yRƏ.hA�T�GD�G�x�s ��PyB@Y̊��" ӵUx}����N�<� ��x$�J%�P���!��w(�H��"O�T��))�U�s�A&r��Q"OT	b��#c!�\�;D��!e"O�:���qP��p`R�0�6"O�E��lݬbn��'ŏ@���"Oju2�����㩃-�mx�*O�D�f��'pj�Ĥ��B1����'f^|B`�6���3Si3�$tz�'�����`�2`ZCL^�' (���'@�� �$ܶj@�㈅6!*�3�')B��;m�^�!Y!��S*!T�,[bZ�'[H�&fE$u��6	Lh�<���,}����f�9*���N�f�<��甉~�V�#D�� ~4"GDM�<�0)��0ʙ�0�Z�*��P����F�<IWb�&���d�ق~l� ��Z�<�G@:8�<����
��	R�<I�/q5u�5Bսw\�,#�g�L�<q�I5Q���qϜ�5B�c�.J�<�C��:I�d��.?e���r�WK�<i�&���M"��5%�غ�CJ�<a�J�91z���
� V�*9��a�<�s�4kB��p7	����$�Y�<�s��M�4�?,D��W�<���<q*�D���[�|�2¢�O�<�k���6Q���tm�	Q�o�a�<q�I	�]	1	_r�4ˤN�T�<�$ǃ�,AZб�d]"�h�k@/�G�<	�(ǯ�ک�V������	C�}�<��.Z6札DL�p�6i�6	�Q�<Ɇ�E����ң�1UH��a��v�<Ae�6�ȹ)%FRj�Hr!�]�<�%J8lP���M5]N�q{�%_N�<�cc�b��q7#֯t���٣g�G�<iChK&��24I�-�R��M�<���)=�{1h]�N_{��R�<�!F� �f��fݤZ��u㥖L�<ċ�W.��rO�$%�ޝ���B�<�uA�Ɲ��B�!Ύ݉F�U�<�2��;6]@1H���E ��U��T�<a���$H���è�)n���mP�<���S4;�N�a�k�rR�)iNL�<�DL80�:u��MN�
���2��D�<���\�#� �`�R�.�,�!aO�v�<�C[^��sB��}N�|�ӣ�z�<I�g'e�>���I�����7lu�<����3D�L:3�S�N��#��n�<A�k�
��8�'�	:G�	W�Zg�<Adʔ�HF����ƍ��� ���H�<�2�Ҧ@�V(<�:�[�jExR�B�ɧ2��J�KR�}�`��Q��U��B�	��M��+�I�~�7��B䉉tdI'�� ը�@�܋=��B䉵-�,��2�[I�P��d ε8��B�I51g,ՑS�Ѽ>�XC��s߾B�I 6����0$8Z�����C䉨��D��L�5y��� �\!��C�	%"�X���)Ҡ`T.���"�5$��C�	":���`�Ǝ>]��� բ�C�IK1��@D�$;��
����� �'��u	�� �h�f���/,�6�
�'�`#6��[��|�`�)&x���'�<�)����/zLjp ϩ4�<��'�$�)�' 5�@�*M<y02�B��� 2���( �p7:	5�V���`�"O��gf�h֤&�)-kT��"Otr�1~P�,���Hf�h�"O�=Z�l��Svp,���X洙Q�"O��ɲ��#xA�ij�a� �ĤXv"O��`#֒)T2�p� �V�����"OX$V�x�0dIb ��4�n�3�"O�M��*�]9��S�.T�[TN "O�����U�K|�]�t�1Q"�qf"O�Q�c�@�P�9�gn�8-H�"OVPp��2��@Cag�?o+4$��"OF٥
�w���M?)����"OD\Y�A��y���j2��Sn>|�`"O����>35�j"�G�f�drW"O����`O0'�ذ��D�2ND� �0"O�{�@ӄVJzD����LH�̈�"O��8�K�<Ĭ�'	İFd�1"O��Gn�'x����&�V,���%"O����	F'#?�y8�NA�lv�쩷"Of;nI�uC0�8���c\��3�"O&��@+ؕZ�
{���$?aR"O��F��X��ϩv�(��"O����͗�7��8C��X���*O:t�׋�&�ZQ�%� �|�J���''
�i�b�#����]%"�����'0$�����J.�(4� �K���'[~�����TP:6��7E,N!��'�@ ��'��1&��7y�#�'=�d���B`!�t��G��1�����'�,ɳ��"{pE���E-r��0��'�5�0Lܪn���G@3����'�2}"aʕ6ke�"�6m2IC�'.�x���������C3Y ��'�`!H�A����2��L�֍�
�'�< ��$Όa	�Ȅ�LP�-��'�P�XfE�:9��$��B�@�<]b�'A°���ϭF�)��͹k�r��	�'	�0�Ӣ?K���1EOQ��\��'@�����DPs@g��L���x�'i�PH�$�E�
��Cd�A8�'Ӥ8j@������AW�(s^���'�ܨs��p"�}��N�N�nT�'�h�,Q6�����6Z��D��'����*�6(�^]X$�W7". �'"vT1)�/�d9i��E=u06�
�'�0L24 ]�r����� i����'
�MJ����zZ���ȯd�^�K�'!ZM9�j��H|��B٪Z��'J���$,�s�8� �h��=`�'��Ti1"F4�\i �A�%|�, �ȓn�Vd2s�����GD(�~X�ȓٌ)0��  o�N��/��1�ņȓ^���#4F��I爁��M%,�歆�cX��7I΍j���`(Y�T�>���`v���
��?<�{Al��6�-�ȓ��}S �7r������#<z@��`�&$(�ù*B蠅��[�ڡ��%A�c�/H���� V�n>\��.�b�K��Y>n]I�,��0E��
�衑	�:OH�ͣR��}����	@�!;�*�S���{���v[���ȓ@���S��{-��Ha���r)�����M��F ���(��=�l��"��@W�m�N�FZ�|-Х��S�? �X�E�A8@�D� 1*.�-k�"OҔq�H�X�-���*^���7"O��e]n
�Ma$��Ұ�Q"O�5��Y�$��J�M4۪h�"O�4 ��p�~%9�j@�
��\bP"O��C��:H������lJ�I�"O��2���t�y���$I@�#"O�P�EO� >I
��؍7�PK�"OF�"a$����ul�<"�"�x�"OV8�b���F��A��)Ðe�"Ob)r`�U�H�d�'	G�A
B��"O8��@�8abGFٮ9G"O�c�"�
Yf�XW�T�8ӞhA"O�蝖1�@JpE�nβd#A"O���oH	b�}j(/�ٚ�"OXxQ��ݪ���Wi_b$�3a"O
�B�bǌ%ђ�̞��!cG"O�	���r�� *ƥZ{�t��"O4�զX+E}|���iA�����"O<X���؁Ji.uv��Z�m��"O�L��N�b������\�"O�\[���E�L�)#�%E�t\��"O���!j=QH|�$�]�C����&"O�������y"h��!�K.V��� "O��x�G��RM؅-�L�)"O�A��.����T�`iP��"O,qȣ��#@��� p�I+[Xvt��"O���/K1!��u��eE�TBbq{"O��"`W)s��g��7>1�p"O�91���'�ⵂ���U&�v"O:�(࡜�d�(S����e�u"OFh� �ɌH�
�k4+C�ʕ��"OֽI%+���fq�@��f�`D���'�:�a��98�hiZ�"�<Vk�-hr���,�L!H�h��M�ȓ}�l-A��=^u��j���-�ƹ�ȓ�d��B�|2�1��K,�|�ȓt��� �Q���6�(6%d���7��E���E��.iHg��A,��2�hyy�T�
_��#MU�#��ȓ;�L鰥W�J�����ۃV�9��i;J��fmR��)v�ǋ/�	��-q���$� A{�g�3N~���z��4KҦ\�(yF({6��8r{�D�ȓ��lRF�Ɗ~�ڵ�7�U��͇ȓV_���" �>�:زlا=��9��ane������(+ѧ�!O�>݆ȓ�4R�[Z�fLz�o�?W !��3����q��2l����ޱ:��ȓ6���h4qp1ba��	�Е��"�>������z�Je��eP4q��|����YN���(�dC�W|�� �8�܅�z��ڑ�@�<܁��ׯ��E{r� "����X1/7�y��/(�M���}oŲP)-J ���4Y�b�B�Gg"`��@G�Ӡ�(��ؖ��$
�8J��{2	"�
m��*�g'���)��%-��0$�[ :S���a�u��B�	 |Ʊ�!#`��%[W�^7J�� ��d;>r�hڥD����D�YC��$�ɾu�-E�c��m��L�y����D�Y�R�Z� ~�I�FF�(9c�e��!�� �%d�$q-�4+���c����A�Lv��ʙ�3��+��*�ĉ�s����B�(_���f�I8O��:Q�b����/�N}b�'��v�^�X�ǜW���Us���n���f�//��@�Q��*	�4ϙOn��T�I;$��7�~���[��n�(<ݣT͗e)������!�d�(�RuiB�:@��ѥ�?\�Xv.M�F$|Т(+>j��׉��A�RtkF�=z�b�� y��c�.��#Jyb$`��'��`�� �7b*䋓�E3at�q�FO�Nll��
�Ik*��!�LG+tt�����0��ߓCےP2@I_�jp�T��g��;��O�ի�%�2#�,
t`KjF��*R	F�
�r,0tcْ ��T`��Z��B��
�0�����y��IJ�Y1�	,^���Au��7J�%�0��0����W-4���{��Aj��y>�Cq���y�l V�N�HkϕP�   b���0?1�D՟�(t�
#����3C׋K�ta����"W*11V���Y�t��O�+��+p�C����rk�^�$���0�N	�,��On����kӨ!yB���$�aѽqR���S@��e��hxBA�VRfvn�E�Y����Đ���I"�ܔAq��)�$��DH��0��	��I�!A*|d��-,3�J�9�}��a#��_8���! jak���h���:!�]t�!��B����)ο'�NH�C�
�1X]#�"Yob�z�휴X�,qY��b�ʧS����aU��p3Eq#MM�G8�4��i�<a�[�}P��K�.�	�F���+V�0��i�mb�"�h�8;9��c�K�=���I�r$ʥ�Vo Pt���a����<�Rg �ؖ�M<�:��u�h�b��� 1��y���)�X���:J���׍��=��)�6�� $����m�'�9J�ϓ)n[�#4$��x��t�`��D;���i	�?5�FJ��8�)��  �Z�DS�M"D�a�"J8;+\��X"���)�1F�����JɥX��A#.F�QXr`�&Bh�It��Ð7�,���\�yt�u�
�l��t��
O�AC��W905���1T��1&�
 ��4�E[㦝8�� �DX ��ՏF��T-8�I�M
&$W<&о	��A�N�
G$��q�A�"�'��9*B(��	T�dR��A�!W0�)����O��%I$��	[��q�'�4yS�OT.3(�Ћ�A�1u��s�Or�Ce�N�8�B���4W��yR�K\>hLЊ�I�5f�n�� �p�MFy��M3Si[ve8l�"O4A���BI���)`gތL���p�JcӸ\�"M�El͘�E�/tN�h�2����ޜY��C��e�!��e%ﶅC�H]�1�ȫ'O.�O�!��mGZ����aA@N�M��L:��t�!�l��0A�� pl�ٓ�τ���0�ъ*O��sbG�S6^O���AA�y����_����"OD���(<J`��!�t�h��'�|�)�42�Oq��(�� \g���2��a��su"O:hP�ނC7h!`1�H�-����2"ON8 ���=Y}����c[�����"O��:�WP��2���3,�(��G"O��B�(�o�|%"���3Pv$\b"Of����݇m��!��f�&x��"O�|*��ׄ	���l���"O{b�
Xs��	t��K̔LY"O,Lj�f\�-$�M�'�+t=��"O�Xr��M����)�����Ze"O,�qm/5��X�Wfw�j��'D� Jc%ۺq�t*O�'x�`B9D�L�E@Z���l ��_�v98�D=D��$H. X!��	�LY��.D���c�&��1@���))�6��k8D�0�E,[�l�,��Oٞb��=br�)D�� Q75���P�F:c��Xɰ�3D���ėo���Y�U����
0D�DY��$o<���U�t e�*D�TZ�"K&C3N	�EGދ7F���G�*T�X�4�\�+���3��׭��X1�"O��R�&P4u,�K�n��u@�"O�1��dV!����P�@Un��C"O����Z=4O>��d��"SR<{"O�IP�
�C�(+���%y�L��"O* �BNTA"�i&_� W"O�<��G�%��l1�� .!x�P�"O�U�ml�tr %��p�<$�6"O�H�AñZ<v�0��Ѥ
\q�f"O(˶�
R��t�T��!Q���"Oz4+d�/�Z0ɀ+�>�j\�"O���܌"�,�G��if���"Op�Rŧ�@{иX�D%zTL�%"O� "����/�T´�͸W�̙�u"O"��B9b�lآ���5K= <��"O��
gF�_XƸ�p����Z����o��H0�I�f-�
"����ل�zi����T�@*��A0Խ�ȓgp<QB�A1��p䇋�A��F~��2Z�Q>q+����Sf���\ A��M0!�2D�T)R���g�
�{���!��i0q�<{2����$�"~:T�)�؈8�aԳx�e�u�Y|�<)r�B(JOl�!��<���+n�y~BSI���S.�v8�����,|p�����'h��4�Ч<�O tk0�_9� �����"&2
!�&��B9�qJ�.y�:)��X$ A�'�;m*��s��A�M�8tFx�! �0HA�vG�7ZT�������F��a��/���tz�b��y�%*$)UH)Ms��b@�h��PऊP����0�_F�X7�s��S���U6y�T�ò7g��h��+D�\ $�L�"U����k3~}����% B�Ð!B5� (�2��'~?����-��
�Y��|x��J�z���ݧW�|�@��?j��Ц��H�T�{4o͞v�xfȉ/-ھ1���'5КpI�S5�B���Ɉ}�Ն�2�rDc�Y�NXZ� ���'^�0Y��"�*�:Yq&�Yi`���rE8�$-��78p`S ��m��� S��R2h{�EP��r��H���ΓCۜieĤ[�=��ĜE̔�ȓ �|!���։aX����:bt�iXz�85ہ4{�q��IW�u�!�eE"�k� �|L�iQ���~5����mj���ѧ��?K�E�CB�G*�	��^7�e;���/q��0y�*���0?Y"K�TL9��AѫL�b@~�A���g�l9R2��&/:mn:�S铯O٦ aD_ ��)��z�<����(�H���/,9Ϊĩ���
����u�D�mB���Z�j����
�<1V,AN��$�|ڦaA�L�t�<�b��>[0gg��D�f��w�@�j�(���1���H b։9��;��Ot�"���.�*Y�&�� ���'��PEH��u�&k���tlC�{mR�{�Hƅe����D���p?�R�U;zk�ZQ'Z��5Ju�g��)��E:��XU/J�D��O�г�
��?���$�ʣ+��!I	�'F�a
5��J�V�*�9+�֡��'��UȲ�P�)�X��V��}B�#�*\V:YQ�ӶP�V�Q`A�[�<�J��c��h p�ؐO��i'LR����D�a��	�F����3�I"ii��3w,	7 g(ÊD�~��dU�!?HIG,L�|B!�	S�D� ��,-��5�#O.L�q��_�� ���%xGb}�3��4ZG���Q!O!�O�2Q�'�_�v�=P�A�J��Q�'�Mb���lc�K���'@�����fjɧ�����k�X�T P�Τm�F���"O� �D��m�w$Q�}��\(Øx��X�X{�zb�ݭg������-M��5�F�yR/݃ �8U8�bҰ6U���E�^
�y�K�'?� �Q�44�ix����y"$��y�e�"Ӻ4u�D���ݬ�y���x�B4R��V%�8)����y���H��؀t�ΪYA�} ��X��y�Ȁ7E�y��@;K�z�MK�y2E^�dM�}��-�@��$�P��y�����B��(�5�>Ph�Q��y�o�<A9��D�m�aca���yd�"N�� ��\|���k]��yB#V�/�b�2$M�*U��ª��y"�A�[��9���X6LH���)�y��,K(�a��\�I��H;�˵�yb.U������Ģ8�����cDG�<���	�T�H%�f��1�`�<qC��%-�8$��Gk�P'oM|�<)C��4�$�AL��hz�"��{�<�G� ��E�D��G��0�T�Ct�<�  yʠ텠\(�̣f+U�\�"�"O&�8 "U�6�,��S*��k�bG"O��"f�A?�mqUF�9�4�"O�1q�!#R`�E�Ʊ7�E�"O �3M�4�6��G�M	Y}]"�"O���Mإ1�|����?-m}�!"O���eLA�Z��)L��T���S�"O��"U��@npa�ĥ�@��"O��@�ǁ#.�$(�s����u��"O��փ`�ҹ8B���6�s#"O^�a�)1������ikv B"O8�jg;���`�p�BD�v"O�$8�BI�I����ȋ;��I�&"O�(z��Ԡ8?���I#i����"Of�9�m�}�P"�C�6b� ��"O�LH�%H�J��,��S1����'"O�	 �A�j����'�F��l�h�"O����%On��s��>�Y "OX��#噍}�0IS��͔C9L��"O�*��]B����a)��d"On)��䂢�|l�c�C�x8h9"O��2f�%_�`ە�ھX؀H@"OPj�/�gz�X����^'|5`�"O�Dz*G�0!�/��#���f"O����'��>|�EN��e�H�"O���K�nY��oU$8�u"O:}��g��tT(b,��S���3"O�YX���^5�H"�	��d��Ua�"O�Y�T㔮f���B���e��"O@�QA��%z�+	��ʥ"OҠ8vg  ,z}3q����@Q�"O�d��J,�pɊTʅ�1��L��*Ou�h�L���Y$Ŋ�Gv&YJ	�'Yv�s���b��
��]3o��u[�'@�5
���;j9�u{��ͼl�v��'y|P8�f��ߜ��F*[�z�H�	�'ܼ���/��Z��LJ4&����דv7x ��A-@1�p�T�>vL��QY�/-,m:�^��B䉲 �H�g,�4Z�Ԭ�lG� B�C�ITo�Z��D���bF��!��B�	�m����`��,B�p�p��8��B��"_�"��p+����ql�:��B�I�m�d8��Z&� �W�۾vL
B�		8"�xPdL"r�`f蝋�"OX��1��#y�d�"�hՌ_M�	��"O�D1�G"Â4Pf�/LG����"O����ᗞ�,�:S<4�ˠ"O����#,Sv�|p+�8��H�C"O�y��ƦAW��S��4� P�"O�|Т��0i�.�a���0*�v��"O�]����c�(9& �>{��j"OjY�t �8@��s%b�'Sh��hd"O$���-��J,|�a�;����'"OT�p`� �j���R ������Q"Or`2�
~U\LP����!"Opm�AȚq�|̑ďE-]X��6"O@�S�l�9��C�J�KP*�"O����ͬCpyB��4�Ty�"O��q��S�l����P�3Zd�"O*�tfL0mTB�w��$`�"O�Q�d'ߠ �	�4��'L�r�QF"O<`��'�5J��O�a��#�"O��(6#���d���O-#�}�`"O��@�i[)DIa&f��ʔ{
!�� ����k��p��$R�j� ̄�x$"O����m���s1���	yQ"O��I�4PZ=��
��+�PA�e"O�}R��۽!��<!�H�|�Lpg"O�H��/f�U�$��h�髄"O`x�À+K��-���WY���U"O�,���Y� �L<���;'h���G"Or��&%ĕu�q���-I �0"OK�*A-ĥ�B�u�5*5'"�yrJ�X���0���=�̉a�
��y/C=n�D�����|�0LB��R#�y�,�2Sh��`Y�r{L9�\�y�b̷
����Qp9ri��y�J$D�VL��$�Z�Q�[��yr�����B &u(K��N��yRF�h iq���H�`��P����y2�@9j�H�%H������Q-�y�A�2^n��g@�0RUp��&�y�(�|��ݻ���!�xrwNߟ�y��'3r�ݰ�'���e�0�yB!׆0c<��g�2,�Ԥ�$�yB��8��8ӄE�9(�ȁ�����y�,FgY���)b�H#�$�Kr!�ē�4���P��K�p4$SgW!�䀹;ۀ��EE%M\fN��"O��b�,��M�t07�/l4fac7"O�@��N�<Q�r:%�ѷf�Yv"O������ ~��� ���h1�"O�-s�i^�ZO�%(/��ly����"O(�Q���PyG+`x< &"O�x��e��gtk$K
2D�1�"O�:�@*�0�HیC��M�1"O����5cĵ�w��.z���C"O8d��,a�\+���9$]���"O��:%o�DJ�g�={X,���"O(����y���#�]qE���q"O�8���dTntBC�Q,��A�"O��m\�8Hq�����!	&"Ox�Jf�*+2 �!���.�ҤQ�"Ot$y�-9F�ҠpR��<p��i"O�DI��(�Ta�Q�	_
I�f"O�}� Ò6E�T���	D �yd"O�=1����'wnU��'(?�e�f"Oup���+�2|��M�n�)��"Of5�Ce #M���H�E8RI""O�Tk�dWY�`��
�q9P6 "D���u�܀�HZ�*rp�'�?D�h�&��~b���$)�UF(����'D�\Gʌh/��4���6_P�C'O+D�tе�[�.$yC��Ԯ6&i��(D���HK�t^���sQ�^wN���#D�h���������A0���,T�4���3v\=�a��*[b��"O(W�[]��4:� G=>\1��"O\���i�]:f�@F�G�ج�E"OR�1�L�K~���s*Q�V|P�7"Ol��(Η*���ˀ"0��h*2"O&�zE�3UN@s�L�+��`�p"O����s�:Y�%>m���1D"O����|4��"��Na�9ؤ"O6٪�J=��t�Vaܑ1Z,��"O��ǈ�*�P���oK��@��s"O2���
�b��XO�
��ܻf"O�@�Ğ��P���mϪ!�4�"O� �0kW՞}Z�x�ČP-d��Ԫ�"O��?npi̑5�v5A�"Ox�I�bS�0�4���j���d�T"O�����/;�\�%�U�W�X�SR"O�xK �L/D������tB޹��"Ol�
@˶=�&�YcB[ ZɄ�x�"O2`"�f��/&�i;!a��!Ҿ���"Ob�Fd�-|z�ꣀ��l��Y�"O.S"K"��Z���u�J�g"O�Ր�X�[�	{�O��Y���n6D�[p�J���y�th�_E�%Ic�4D���1-��E��qb�Ϗ^b�u�#1D���W�Xg^Us�+V��(��$D���@�l�P��˅%d=�8 �#D��j5@N�q,&� e� *I۴��� D���� ����%�^(B���%�$D�L����N�z0�)M䪉Ѓ&6D�pa!-˿
�P8��#�!/��%q�2D�T+p L:&���-��Z���[�-D�����9i���S���'��1Bf�5D��zvo�"�~X�n��JȚ���d6D�� !��V��2�&F�k�(�x4�2D�|�P�ɹ|%����jG�+M��Ae�0D�HBDH\#��rA��{�t�c�/D�l�wƊ�t�`���\���M9D�l0��HN��l���f�N���e8?ъ�ᓸS��� �V?+�n�(A��z�B��=]�������JT8�A���R4B�<;M����]�pD.Q�!no�bC�I�\?:����,+��Ĺ3&�&�RC�I,C�e!NZ�S��\�fa�9��C�I�d����_)RE�� ���3�C�I.3�f-rD��F���� ��5�bB�	�w�p	;�O�;�% ��i�*B��*9.���DTE��@�1�6C�ɧL��`���*HK�p !�qibC�^�qƅΩn�h�g�6�\C�i��2��Ŕ}C�QP�HיVuLC䉼to�hC��͵C���a�TpC䉡h�6����ՎM頽�T��;_8B��IlE!km&����J�`B䉥#!ԑ�`޷PC�"����(	�'	:87o+>�������2[�Y��'�dl(C�[<�9ӁM�a0�u�
�'����E��a�`��R�W+|�Q
�'PD���@p�H{��ֆ%�|���'-�0��#٣HZ�⠙?)Y`�"�'d��9��A�uŸ ��>M��i��'�XĈ����(�lu�g��!rd�D)�'�.3$/����ъS�f�zȊ�'��P���lB H�E�l&(���'�nݡ�+�)]��I��^w�v�!	�'�R��� L�L�j��Bd�����'�&N�<m�<���FR���'�JL���eZz��d���h% a��'�lQ�%�K\0�3�J�5c�x�I�'��%�'��,#�Qi��(��
�'hмz�I,�<��d;)���"ON$SW�%%*�8��EF7R�`���"O�l:�G$_𮈑�%�f&A��"O�l#��V�XCFY�eMR���t"O$I��,<����qeE/A��	�"O�I��H�s��I{�b�8'!$x�"O�P�`���U=�� �=����"O� ��K+D7y�F1JaG�c��"�"O���E��'�P�s'^/v$�4J�"O$;AkxU�)����(�D��"O(���
�'uv��ő_ ��"O���!}������!'�=c`"OA�Gυ% r�x*���`q�"O$0˓bP�,��C����"OV��&"ƦT�(8� S�X�XJ�"Ol\#c��8���ѯ�� Xd)8�"O� Q��iq~APWlK7M=r-��"Oz@;G
G�R��:CH0F8ra��"O$�[�䖄c<����jغ/���	�'m6��&��nLz�{�J!{� ��'.^`aW+��K"��s�\��vy�'\48��3[���A���4P�'�(�ES�X�
r�&0Xj���'�%�7/�:"v�(��-~��J�'Kx�:�GT	�b�sL�s	�d1	�'���"jɵ=��k�c�{�5	�'n��T���D
�oYtbX�
�'OZ�cu!�MF4��C�72���' ���H_3l���[��Г6�8i!�'B i�i��G&���͗�ݤ���'px�	Q�� j��Bxs�2	�'�4i@����H���ȗs����'�ny�%n?���q�^��L�@�'�j�s��>Zqa\B�II���b�<J�2V�x0����9&ZZ`�A	�\�<��OQ����چ��,OC���C~�<��Au[ة%'˟F�v�<acB��(���+��#FlX\Sqe�w�<iR��.Mf$q�p+@|౫Äw�<yG��|�\��w���>�dzG�j�<	"n΍V$AwF�>��dp��e�<Ip�٪>ݨYД�юk��M��c�<����y�
���Hщe���d�YU�<1�j��l��L�NG��pH�G�M�<!� ��|���Qc+S�g q��čM�<1���@�7n�j\�eb÷�y���"9P2-��}����
�y⤑�@�L�#G1yZ��`5 ���Py"���zT@��5=r��)���W�<�eɲ%E$UR��7{��1(�
�y�<����g�� 0���}�n-�`NIa�<a� �{�PCwcˑP���a��r�<a��O]V\9�4*�C��Q�S�<1�bg�FݳQ늀cU�(v����y"�ܟ� \`L\�TK@��IK��y��G�"=Ψ��]�8�(�(�Z��yR��A�
�+��8R뵇��y�l�,d�v�B��mW�	Z��^��y�	�*�� ���&_ЊlJ��A��y�b�:�ؓD)��Y��!��ύ�y�댍 ��z��9j��ᶁK)�y��ăD�������+�H5��IJ��y�N[��+U�D�u���y� �-J�1��)[{��P���$�y�ް"��9��
�J1H�@�샥�yb�
�V�[�D�G1�y��R��y�٥(�(A3�(Z�8 ��rC�"�y!V�|\���c�2Rs� �y"�Ya�����t�d���y��;��Q��-Tl�`G��yR�W"^�%iU�\��e��
P��y
� X�2w �D�|���F� }�"O@m)���k��X�6��Y@"O0�����s�v���R�{.@)5"O̔j+֌"ݰ1A��$lp,��"ON����Z8��O9Qr`s�"O���+� �r�r@%6Ob�%�"O�}K�]�V��uyk�TV���"OF]���ޞC>�k!��X@���"O��(�_�$��,q��92g"On��jH�lv �lيMm2ĩ�"Ox����A���iT�O�|X��"O�� �F�4+$����9E�0�v"O�8��
��:c�҇��.\��5�w"OΌ�Ί�l��Yq�g�H���d"O
(A��ؿ4�엄Dj����D��y�sD�񳂉ND
��A�N�;�y"D��r�e`�¤B|2A�RJ���yR%Z�dF(P`P�:F�CB$՚�yb\q�C���+�Z�����y�.���y�	N�v/�A����yr�X�+��d�%�nb6��!�H��y2!ѳ@K�	��c��]�T�)1j��y֡`��ҢT G�����KQ�y�o�%_$:��PʼC'^�p����y�g�<��c�d`����G��y��CLH2�;�i�_)�lw��!�y2.�g��i �oD�[r~���j��yR��#;.TkPc˅Um̤( ����yBN�#L�l�ڒ�ӡw���w��;�y��/I��0p�X�IG��/�y��<'�H ����$4d�$D'Ɯ�yr.I,H�@��V�W�_�h�Ϛ��y2V}�nL���0����͊�y"fX
n����OˮU��ix���y��_mhy��\��`�#"f��y�ē�e$4s� Yrx@��ю��yB���zd��Վm�ts�	��Py�׀~�T�Qt₩j�Nͪ�%�s�<��%�� �yk�ͧNV�R��f�<Q�b�Z8`I�1*V$ �f;��X�<��߫ ����Y�[��\�j�M�<��O�QX�Pږ��u�n9P'�^M�<���0��D���Y�?��2�UG�<Q�MںC�j�I&b�X�['��K�<ѳ&�"�
Q�L�>�(i�ce�H�<���F7f���+�lu-%��A�<�0}ȶ�T&Y�H�Є�Ц�b�<�g<i�(�2F�>Т 1�^�<��/\�
��i�s$P7}�ny� �\�<Qp���hay�DY6����U�<��˷FИI� ��8P�!�fF�e�<Y�!h�������3K��谪Xc�<)�h����A��4[)���]H�<���3H��ɺ�e�?�r1�#D��t��cd"(�5�<�JAp��%D�0)��E�7D�*ݕw*� �"D��rq�6W���ӤE5w��@��b!D�@���Dh�����Cװ%oބ��4D���.� S�(��	������I4D�|��\��<�q#�X��0�Pf5D�t[��L� ��W)Ɗ��jՏ1D�h١�'=���Aʅ�f�=r�/D����F����@��cd�� a.D��p�A6Q�6�0(���1�a�8D�� M�u���)��%���sو�ل"O�� ��
	�J�������mÄ"O(	�ŮÁCҦ��aB3�����"O✁s��nڨ����*7�Q�f"O�ة�� ��~�`ʣ?x��"O�[Tj��-p��vm�?V.�	�"O����L	0�+�E�H�X�"O�Y.�jl�6i�l|R!"O�1�JI$��e�6jR%;Tdu��"O�i�ּL*@��c�\0��"OVYCQ��#��U�Ӣv�hp0"Oؼ����Svb��6���ps�"O&u��h�Bp��Zr�m ���"O����FQB
�dzF�؀`U&�"O��0��"+C�l�L�!9.H��"O��	S��>d��#��L,V4�"O���Q?��Tp��ػ��"O�@Y���[|��9�i�������|��'���"��1w\#$隖n�A�	�'�H9�q#�r��	;0a�)b�na��'�0ٛ�%@�jE��kv�X�*	<���'�8	S�<��x%f vH�'����
��m��äÁ��H��'�j�3J[A%���Sa�	 ��'X�Q��f_�jR$���M�2���j�'�r%"Z
�!3�/J~���!�N�<y��	 C��-�
:P�0��P�<���O.s��4hN�i���@�J��hO�O�X���z�2�Ȥc�,�R�Z�'b��4BӌC��x
��!��<@�'�&�{aD`gbŘ���q���'�����).�|� o���A{�'���D�ӊZ	h�)�����'��7M��&g̨;t,ב^���a�
H�!��9�q�a��m���5�Ǵ!��x�	�V7
���	��h�q(
�<�dC�I>p,Fxy���#f����&�^�.�y���"|�E�,9���`�H68{va뀃�b�<�����f�=3�x��q.[G�<A��G�(P ��M�@�h� ��{�<�FEN'�Eh���3Vaz����r�<9�!**(�%��/6v�ǔU�<��M�!x�=�gGSn�0�f[L�<7 Y�or������������]�<	!̌P��,�u�o�����c�<�'@�]j���M����` v�<)�iK�_2.m�d�T�w&���k�<A��\�G8�b ��Q�8f�[P�<Y��]&@NlpfH�6�h�E�
e�<�e�d�^hˑ`�38���ZяUU�<��L�~�H��2�R���];�
�Z�<	M�/�:	ۖ��3��E����T�<A� 2d����ȭ4��z��S�<�U�\�H+�5��`�,8
�,�Ҁ�Q�<Y�&԰-���I�*PCYP�	�L�<9�F�����M'R6VY;`��I�<�"�S�8�)�1��p�iqCJ�K�<AG��1n�����Cԝ_@ȡ8���E�<���Vbm|uڳ��hX�F�<1���>6Zt�0o͕N�:�MJ�<�6�̎Lt7�����
���y�R1$<�U���ld�]E�Q>�y�m��]�����_ҩ�SOU��y���)N��T��+��@��.Ӳ�y
� ���$d��$e���G6	\�{T"O4�����a���B��,���pV"O�}�֊�$>�}�BA�a�VT�2"O0L!CFP-R��G`Q�+δ�F"O��H�l�� $�h��i�&�x�4"O�p�΅�$��5��j�s��³"O� ��ɾ]V���C�V�]V q"O$@�6�́VQ�p2�K��5��DkC"O��x���g�Nl�1K��(�]��"O�P�*�1�nM��d�g����"O��YfIJ�a��1*�C@�E��<�"O���g�r�(�3ԡ�J��h1"Ot*4FݥZ�j�V<%¶a��"O���ģ�#�4`�Ï3�ԩ�"O*��Ʃ�+_���*w��(d"O���+	bt|��ࠃ�G}N��"O�M:�R)��a'π���,��"O���%��o����$�F
����"O���$/�6�)�Z�B7ڽ�S"O �U��>�n �&�]+*�k6"O�-ip	A�s�b���eT=h%0���"O$�K�@ɨ]���"F��	J�"O�vm���l�BEN��[y ��&"Oڄ�1$7��P��엲6qX�!�"OH��$��0��{��T5~{�d�4"OjA�T�T�K-� $E��zoF���"O��C�Va^!�A#S(x�"O���U�L���W�5�<*"Oܼc���1`�AՌ14 ��W"O�=��bV�q��t��j��1�w"O\�؁#0��I�,�3{�0 �"O6�B��C%dE:-�VJL�)�D�J�"O��,y��h��E��YRf�(D��
�y­N�cώP8�G�)��i�$C��y����5+�-�R#ϐ�fQ��3�y��?�V��F�߯@�V �H���y"B��CX��X�BJ2!FN,�E��	�yB�X�~�K��WFd��7#&�D��v�؈��+D�k46�h���3|$<��-2�Xh�M[L���(C*�1bs�Ňȓ�&���˗Z�LX�(b��ȓHz
HX�KшߞؑDH'T� ��F`�|s$g�{��x0��Ӣ[����ȓT�hP�4��JJ$!��)���p�ȓ{lzx�ҏ
00�b�wG��r	.h��	���C@� '05<<q��J�6ޒ�
Ӣ� {�X|{t����?���?1��?��=y��?���{���]�� ��Y�n%����!	�YÌLؓ��*'D5y��$|NT;�*E_�'��pHP��P��A'w>�5ke�}����d�C�V���;�%�(de-�d���N����|B����?!ٴq� 9�Ё�0}�vt*r�һ3�ʰ�s�8�d�<QT�8���u�6������5z�}y���$L��cT�X�0ʦ*�d�d���C�I��q����?A��L�tq���':�6MV?9':X�;�?���?���k@��\���]����j_�����?��u����e�R%&-dL��(�
!�.Z�P6(��@Mg��I������!��LS�'�潈��0`Hd� ۢ���^�iԀ�q��|���a�?Qx� Si����X��|BI���?9��i�`6m�O��'tHN�Q��}�@ 8s�(��A�t`N7>�	��H�R�
n �dkG�g��� �eY��p>1�i��7�j�\tڀ
��$re2p˒�a
�OƉ�͑æ%�	ʟ��O�p �d�'ҿi�B�H��V"bڎ���HT��*L���MT��#���4OǎkRM�*��=9�#�U���'��]cf��{�Ӑ30�w��=�R��ٴQ&$�3�dB��ab��ӦIX�)�?v*�t� C��G?�s�]swB�<5%��8�jBa��Œt�g�JL�w�'�X7M��i��~��MT%JE!z0��9�0H�@�GM?�����&,O��2-+nf������~QA�I����ڴ�䓻�I�{�V�(S�ژ$& c�Ч6(�H��ݟ� ��JK9
U�����ϟ#^w���i���i�&͕S��P�!�T,.��ʃՁV��.O$>O���EU�
���	f����|
� Tt�C�
hFu�#�),��`�GK'�DDXg`�4}�̠R�G~�!4�x �pb�	 <<��P0B. � ��!E	<�P�'������?)&�x"�']�� !d��8���B�_MXd�c@����	ҟ$��}Z�#�9��i�d�DرD�U3\7���I&���?��'�fuBe#�9+}F�� 	�k����i��ű2�'E��'�2�Q"+����ݴN�vx"N�F�	��	�y���;4
��1�B�!O�MF�P
��R�x������z�'�^d
���,^5�PX�]��:���(ҮT���B��]ˇNgi�x�Y*P��!k��
)��Q��5�	?D蜅(P���:/����n�sd���Y��M�����Ox���O�b?����X>+Bd\`F͎�� �!v�B�	�%mf���%����b��z��7B�(-�4��J�b0�1��'��U?M
v!_ i�(��gG��lϒ��� ԤE����?���L��kCbN���9;$AǬk��)�٤6,ܰ �W�#�4� "�ƹ'�F 	AϗP�'���������p	!Ŋ�׮� B��H��ͫ��փ}n2|�4�ŵ6c��:��H�z�=@ԑ|��H'�?�i�6m�OP�'9���� G�&�A8�!�g��sx������'��\�"�Q�Ǽ0�W���? �"	�E����v��6�;d�����6��5���L()Q��$�D�>!"_2   �=�x�1�I>H�fak���0����)26ۘB�I?t� �  ��L�p/d,@�'4D�P�4K�s%Ic+�:4�|�62D��l��$x���*��+fV0��lJh�<��-�:���
7f��xq1M {�<�v�X��X��>w��ز&�v�<���4�8)9�,/'���׍^I�<��
��0�$)N�t{&&n�<7b��6e["���i?�hq�N�m�<)1��,�&��9���E�D�<i *�#2\-�WfE��u1eCQF�<� ��E��L�aIS�:�ar��|�<aT�W�f'����O*Yl��+�B^�<	�� ���ٱH˥6
4L�W�@F�<�唄>��H	�%ΣJ�����NC�<���֊y��)�G�� r�!4�X~�<�f�q�a#\@-90	NT�<S�\Y,h� ����N2�h�2��Q�<�'�ֺgK�d��+0&T   �
  p  �  �!  �(  �1  �9  @  SF  �L  �R  �Z  a  ]g  �m  �s  +z  ��  ��  ��   `� u�	����Zv)C�'ll\�0"Ez+�'H�Dl�N��:O�1"�'"d7�R�)R�ĞH{b����L)<H�yi[i?zhЦ�� �7C~ݵo�?�ѧ�?1Hw

�mR{VA� t3hň4��IЌ�'�Z�*������.l�C&g����?��I+e�.}2���7X!���d&lŢB l"đ+��o��z�-�U�n�91�i:�M���'t�'d�'��$��	�$2$D�	`Ν���'�r���>/vMkR�T��v���Sȟ��	7�2̑���x�Rl��M zL,��Iğ���Ɵ���ar�]�	���$m����9�p� �$
=7d��v�иK&�����<Q�&~oDZ�	�:�H���@BB}��If?�&U���U����A���\s,���Għ�1���(�	��8��؟$�	��,�OH��<_�qk���฻C�GK�Br�`o���M��R� �ܴ�4���i+΍���'��ڐ�C�\���ks�G�t�å!(ғ@i��<ҧt�M���UWl�<���Fj�Ъ�gܺq�^��R#v��y�4&כ6*|���	�(	(��@9�V`�T�HFJ��2F,��P�KD'AƦ�(�hI�k��EJ�j�脳��^+���"ԌX�M�E�i	`6-�9>�1b%�
*�6��@�^�5 @���_�^H2�h������4\^��ݮYw�i�ˆ���/Ў&Ve�󃌯�؉��6Kw�Dzի�$?�Ѫ�O*q&7��Ӧ`ٴ_R�8���85c�]�įӫ�>7�,��8�
8A�}8SŔ�W£As�F���3��-r%�S�;B��E6*�"F�N�{v,����
�8�� �	柜���F���ܴ��	�6�8��kT�j^p���"�0~�Y�8��˟|̧,%�H{��$'6890���MS��١s�Ը*���2�z�G��0<�����g���nك/�z����I��`�`�h̼��A���wR���	�{���O⤗'GP����ھM4N����x]P(X���?A�����Oc�dDT�U���5k�tc�N�k�BIg�(�����g��l�U�Z�pMҡ�3-�ϦU�'
�e nu�nR��O�ʧh$M+��Tr��� ���K+�
u�x�ǬEß��I�,Zh��wy��'��3}Rˌ� ��i�fX�lj`�&F������p0����,&n*�X�#ڧ3vT�p���.+|�1�p�B	i �u�'S����fћ֢2�S�?�'e��+���v9�-A�-{P(D��Iڟ ��~��I�5[��6
��$$��hO��ęm}RQ���'`�J��h!e)����8�f��I?u�M�?�g�'��A�5oQ�VP����л5�\@�'�L�t.�"�4��A-G 7J�(b�'�)BF�<""�zpj�81�}
�'�.��f�]�����U��Q��'y�1����+$��DE�ұ��' f�ȰC�I�&%�@K\= ���a)O؄ac�'2 ��cQ�L*��##�[b$�܅����3f�HB,��3@�P;mC���z���j��(�����w����fU@�*`fǒoR�D��O�e�ȓ*��40��>j%<�Z��&���I�9���ڴ�?9����n΀K�`EyG�A�\����?9��H��?q��?�D�CP:
���48�=33!��r1!`�H(-��(!Gj��h{ޖ�0<)ଅ�	,�%�񎗄 "0��&b��W���0p�+X�f�aC�V1c,���	c��d�O8o�ȟԨk�8Z�̭����>a4���ZyR�'U�OQ>!���˾-���A�!u�����  �IY}R퓾�M�!z�X�!4:J�{��\�0ܛ6�|b��\�F������¤���!�<�0�
�+��	Ǆ5D���b��_d� �$oH� s2=�c5D�L�@Tt�P����%�F�!��; ��u�# �A܁-��`!�"O��t&Z6Hnd�w"�*�Y�"O����\�]�fR���Ŏ���}�L�O���@E��`�D�O~���<�IZ�Y<Yh G�::�zfK�*H�@!�6�ib*6�Ό�vy���|b �D
�.PJ5	F�נG��}��O�a�� �Q��	Ps���׈Ё�����T;�a�'����*�!�&�Q4+��q�1�@7�hykơ�?y�����?��.��9@��+ ���s�7w%��	ϓK$�Of � �i~x���ڋo�xٻY�ݴXӛF�|�O_��\�h���?�����ɒ�D�J@k� |{H ={��X��(�I���ɍ�u��'@?����7���'Č���H�?��M�� lcH���'c�E)�K�x�\ �\Ȫ��W���zp�_�����΢>|H�0�@T�r���I�̟���#�l��b�Y�NF��c���D ��e��Q	B�^+r ,��Eɓ���@&�9ڴ��s�(`2b�id�	8��[�K�#N�i4��2-��ĸ<)���?!�k��yc�NB�d��rrj��y
� ��肂Y0,Ni���Y�^��i���'��PL��'�`Gh4�y���J�����&~l�s�W�0<IŇϟ��4�?a��H�`pس�=�=H��ۏa�|9k��?���?	����'��'l���.(�S�$���	��f�Beܐ0�L1��Ê5�0��&oW��?�/O> ��	���E�I˟�O(�0��'kҡ�`'ƨO�B9��%P��f��4�'R�\�m9��T>�'c�Y�M+qrЋW�������OlX�T�)§^��Cn�. �f�+�,�Qڞ9�'GK���`�M>E�\�Q�P�9T���R3r�ҌQ�'I��*uf��	NP����Lo�P�H��Df�O�~Aau���_��q�aM�;D"�ֽi�2�'{b�'� �r�'���'��=�ܒ' �>`mv�e �7q��D2���,G�az��'d��2E-4j���$��ol�HCA�U3d�RS�{�D����y"ʏ�-��� 7,�hD5�� ��S��'L5���ǘϘ'K"Lꡢ��<\p�DF�j����'�4��ae�^A��R�&�d?T�̓�?��i>�'��iׇ�0���9Ҭ"�FE���ً)/~qVe۟���ϟ��I�u�'��5� 0i�%2
%����,��hɣ� ������0_C>��Kǌ�� ��=dҨprG�X�f���PU@�>�:`r%O�G^��dϷ��a;�&{?��>&0�$�'�@6��æ��?Y���G#kl���-z��h0H6!��	�*n��c" ��Y��Ǟ*�'N8���D��	t� lZ����Im1����3w��B$�'�4���ɟ8�h�T���|�1������<��	�>w��9r���!H��A��~���I=u�d���;�h4��BPh�����Im����@i��%un���f̗}fB 1��M5$�C��%UdRъ!d�)l�r� V��$���dڟ�d��E��b��5	����9��Z�I`�lZ����H�d�T�,�2-�4F�R�񹄏X�y|ţ��''B�P�|��W����}�L�̐� ��h
�R����2�l���8?�W��%[S��x��\�	��؋��)S�}��`�ңz��$Fj���$F����̦Z���O��)B�d_"�h�*A$'� 9ZPb
#��yb�'�▟I�/�[w^�A0ۆ\,X��=��?1C[�d�'��K�X�XJ$�V�T��}����5V`�6m�O����O�PÆn����OV���OV�]9m��B$��r>f̀��L�v��f�U�-�TlZ,0]�)3��j�C.�	�lj����RΠ��%ӂ��Q��k��U���L^0�b�4�*��>3�����P�D���$�!2�&�����M���t�Ļ������Oddq�K�}	���!�|-����-��hO����Q�A�ŊC�F��S�γh� ���O���'t�s�$�'�	�`U\l@� N�l��Q� �F�؈S�E�m���	ӟ�����@SYwj�'�.ۍ�^a��L ��5�
N,����m�l�r��VdM�n-���D�V߈"��ɦtI��B��(�T���`�<pq{B�6D��(��	�s�X��٦뒹��'RT�Vl�O��$��1��Cy�'1�O����b�bGa߂<k�����O��=����?��ybe����r`��
��M�6�����O�um����'�j��kӮ��q�4ag��lڠ��"�Ǽ;����C#�O���?����?���.[��~�'[�4h��'� �YN�?������hw���
�Y�>�g�ɴL��ڰH�<�
�J��
��-o���zn[�\�� �O&|o�쟸�	y�&�25m�+r��@!E&[+X���⟄���l�	B��j�MHH0@��_vX�$I�+ �Y��I��?��E>�PС%��,w��0+Xퟨ�'��: Gb�l���O�ʧ����z/��:�� �$��Ş�.�8���?���ŎI=��!�_��IE��U>�b�T=1�d���G���BY~	G7|ZB��!��S
1�䀗,G�B0�}��`��XU�����'���p�ȈW~���?)Ƽi$v7�OF#|�q��d�fx	!#�s2	 U�X�ן���Y�����E%dV����K<Z�T�����Onmڰ�M�M>�� �X>>�H�X[~��j[�?y6��'����d��h������ 4K���xG�#L�!��T�H��l�UcM�A�P!D��!��D�$��T2�K�=kȺ���W�!��F)_1�����0�t	K�%`�!�$�/8������?8�q�"D�u�!� �lYJ��RET*��Y2'#��s�剪.�V���QHrX�0�g>Rl;���!�� �0I���?�\)&�U�{ άæ"O=�I���z���F�?2��ʃ"Ol4��(����f�LT=6"O@�+��� Κ�D�۶�q3�'$H��'�إ��;~]UXq%j��'NT��4��`�\A��!b�9	�'7Pz������7��-\��M��'�y���.<ѐi�M�V���'[0��� �7����Έ�E��@
�'m~]�'XG��$�0�
������$ �Q?YْMǤDY�t��FT�h�H�*��%D�X��@(|WxlRp��B��r&�(D�����ػsw^�ʀ��[ ��	(D��CO�>B'<ٻ%`�4h��a(D��z�EӺ#$�=3C/� D��鲂 3D� �!�<o^8�[��:e�|!# ��O�5�)�~�i)�(U2?��]9w�ԿHk*T��'�fx��K�q[B��bZ�Hh[�'y\AC�+�}���F�?�Q�'��9CA������]�z6� ��'�:�A@f�,.q�yV�A�o�62�������עU	F茱�7�<��πt8�L0�^k!�� 5,Qp���&D��85��>+���x1�P%5�"l�#D��H `IPA΄��O��a��iP3D� C��J?X~T��"�9��MJ�2D�t���1
��B��y��5ȅ�"�O&�3r�Op��a�٫v�P�$悤|���A"ON�� ��h�Q�����rli"O��E���k!d�"]�h+"O"i�VG�$x�4@5c��<� ���"O�ԡ!���Mٌ�S@ˑ+C���"Ob�w���.�i����
8p�����I(g��~ZD�J2y�`i��'L���i�S�<鶥�tm2�R$-_l�>�i�)�N�<�VA�#G�����%��QD�K�<��Ҹ6xF��!���@%ɑ��A�<)�F�~��x�ٷb�F�Т+\A�<aP-�v�
mC��ٽ}o��g�Oş���A/�S�O_L�#T�5� �;���6e�2h{�"OX����Ӽ$&< b��N�����"O��Y��QA�DY�`�\��V �A"O
���C�l�2L� �O�s4,�"O(�˶��*͌5�rD��`SQ"O~�c�~h���b�1w(�_��[��4�Op�b��Y_#ƕƢ"X[���3"O�p�@ãLW��j�LBUIlAs"O` �@[�!ît�֊�؊!U�r�<�nϻŀ)Q���$ a�]`��l�<��F¬��d�r���b��I8UlPjx��â����J?P~�r�Δ�K9&�"t/3D��(����!{�DYg,��!��<D�`��jp���W�rX�Ԫ�`0D�,h��R(ӊ���7
�T�dc8D�q�4F�� ��'��T(�8D��"dF\$4��yC�j���ٶ�8�H�dF��N<M>�p�i֢4�T���K��y���kH� ����-Z�VI �yra+R��X��j��%��b� 0�yR��?-؄������ ��F�!����rEdCbr	��哩k�!��
$n��be�cd��SkE�-��W��O?��6���*�T ��N�2�z�nI�<��AW�!e���1�����P�g��\�<� �I���]�hl&y�pG- {Ҁqp"O.Ɂ�Â�z��fքy� �Q�"O�hiԊ$o��$��a�8�*"O�8Z��[��<�� �G�O�()RR��	��<�O�	z��ר$�LC�'�!K�4�"O��s��Af�Mp(�*O��}y�"O���hʆJ��צ^(����"O
�s��T<�`�5n�t+q%��yB�ܧeY�D� CE�`��4���V*��>ywe�U?I�ȏ�M��=�c�!'f�	����U�<I���j8��sd�C�T�H5��m�N�<��#�tW�8�5	���RԱ#d
N�<���Z�5�(P�EQ�t����`�<�f,�!7@.u{2��7��XK��A�<	��K%�\�d�&w�i$/u�'+���iP�6�U����#1��gE$�!򄂦��(f�9"�t��B�!򤜊
T^ɫ��{R�q&D	�!�۸@��`�̙U�0�d�'�!��+�;��Q�hEX`C���!�ʋ@������!?)Qf�U�1�򅆾�O?����.m���1�D��@��W�<�	��v����cO�Q�VDP4�h�<1���,~���Q᠋
~�pA��fh�<�v��;�X			Ra
��d�<Yw�q*�
@�6z�A ��^�<1�&�3<��}+B���8I���E�O]yB��p>��Y" f��� ��$ A��Єn�<�&F��*�Еၣj8̑���h�<��Ü$�j��&j�&BE$)f�<�$�|*�93�We��(#'�^�<�煃�Mv^5B�o�B4t(��mQ\x��s5����� �5Jhs�M�;�"�[s�-D���B�Q:{~L��� 5��XC��*D�0�/*xOU� N$}p�ܙ�*D�\ccd��c��I��:z�Sƅ*D�TYvJ�SWR�0�X�i�6A
�
*D��w�L);���@7NR�f�RK3ړ2�< F��/��Gs�BpC�NWL�@ ���y�nɾ�m��e�H�fPA��yRiZ��G֫/��I�$�̶�yr�ߒ-�p����� ��� ����y"=_܈���"�V�X�eٷ�y���'�~��@��Nh��&��?���C�������lp58��u�֚f���P�&D�D�6'L���x�@*ԏ#
�"(?D��ڇ�N�)E�}c����o{|���:D�䁢�C�a0v$C��1AL���$D�|�AB �_���<�*�)$D�HzƈF/"�eKV�V�K�KJ��6���d�L�9�1��t�!�n�L�!��A*�\H�2 �;&��.Usu!�dB.�:9����"qӼ%�-�s!�$b�>i��U�-1����k��hp!���
�9)A�>Z"@A�t��9iA�}�S��~
�tv�¡�R-�^Hs��Ҍ�y�������P��Zq�ꎂ�yC�K��d��˰�ژ�1���yₙ�rfm�} .�a��y¤�;H��mB�-c��k�C·�y"�Y���T�����*tz15@���hO u�a��/7vpy��b�?$���У����B�I36����ǂ+������f�B�	|	x��b��Bƕ�ʃ!_�B�)� � S��΃ �l��J=G�,��"OD�suI�yz��Pl\�y�hc�"O�<{�dK7$�� &Ԙ��1���'�H������`�� �+m�� (D� N>͇ȓL32��#BL�3�~L�N�����>���I߆c�h�b��4kn�a�ȓO	̣�d�f~Z<�fY1l���9�����˃,l�0Y��1)\68��I�,��e�C��%�4ܤx�'�����$��բC-��2���kP�ɅȓQQ����a�NX�$q�N���M�ȓ{��@E���v�de�bn[�J
�ȓEƾ��Q�]q�,u@�o6I����ȓx|HZ�ȏ�E��Ԇ�r�,ɇ��0��I	G[U{�酄Q��� �y+�C�I
D�ڄ+�OWC�ʥa0��-%��C䉑¥���/[�lysU�׵P}�C��9Z MZ�_�(��A�|5�C�I,0��b��I6���ԭP7L��C�	�c�2���tM�YpTʎ5W�ģ=�� �Z�O�@�`e��&�""סX�">Z1�	�'��\��f��d��z'�~(<�
�'�FY�U��;u�Z�r��Ý�8�
�'2�IJ��A�P��a�� �`Mp�'q��YgB.�CDΊ��L���'نB��5)ܘr3��gn��`��;�t�Gx��	хLQ0%IsA]�th�<cR.i`�B�	¨T
�	С.���h���f�C�I+�-'I��
��
K�B�I1�� ����<��
�=H�B��#HNB}1�'}t�����(C㉨" �H��a��{��f�$`�le��K�YZ}2�L7�,i�ߴ!nXZ��b���O�� ��iG�T)։Ք�?�!^�?���?��Ї/<e��&[+8Թ�Ϙ�5�)r��FbEs �ʿ�<4b���"n �Dy��r��c�N.<������? �Lɧ�-�M��גz~�;�� �*��)DyB	���?)��i����t�! �Z$s��i��v�n-�2R�����+)d�����01��]��+Q�r����Ď_y2D�d턙�4	P�U`��3�9��'�X}� ������u���a�!�0�2��s�i)!�Фa�<}��%2 ��F$�h$!�䒬�&�H��\7���
T�4!�ѢU���(��%&�B��ƨZ!�9'�4�(��K%&�b�.R^�!�$_�S6���J�	��(�m��C�����D.�g?�7%��V<�1��T����2�m�<i��=\H`	 ��=��Jg�<AF��+]���/BQּc5F__�<Y�--~m��Ϝ (jA{b�Va�<!�($��U���
q���cN]�<�4���s���˄;?�A��F�䟤 �2�O�m c�תp�X�R�Y�.-:T"O�\����"4�5�@e����ݩ"O��BB��>����L;�DE{U"O�����n��QS \;z��!�"O�P�4J�K�(�@�87Ǹ�[��'��}�L��8����\�"�Ycg\�}� !*�!#D��(�EPD�8�W�[���'�?D���!
�:w�̌���'@}j�3�C=D���g�Q8;�P�"T�I0G�L���I<D���u␊)�� ��~xP4�/D��a	��}ILi���"@�%(��7<Fz"<���!iN�2 ���?w�,��$"O�E�#O��M�HYɴI@2���˧"Oz<�!��+��)"�\�=v-.!�� V!�rP�v�p��"��!-ZPe1�"O:��Aڄ�h<��EŜe#V���"O��H�V6}��
�aF�Z�i�!�O¢}�6{~�ÂO�:8x,��)> �Ņ�QdVUQ!�͕)Mxl�7"�:G����}�d=�(��4�Re�ƾf�R��YV�yqƒvv Db��R�hO� �ȓqжt�2 �yXn5��n�$�h�ȓFCĸ�q����9NyNV�I�aN��d
xa�I��Ŏ
G��x"eيL*!�!V:Xy��̃/7��"�خ �!��+`*� Q���.0ظKF̓�1y!�d�����CP�����ܦ/M!�$�)J�C�`ׂs(�<��ʃ!�џ`ʥg� �M��?y�OQf�q@��7`c����O�{�8{�{�}[���?���o�<��嘧��
�:<j �'#���,��-��O�]0��Ǒp��@��Q�z�'0�Bqp$�3@U�E��uib�F|rFW(�?��ɉ���	"���U0��[�
�6+�!���Te*��͜ ����,E�d��'�ў�����ƩO��p[�lP�xE>a�m\�eU�����s�i>��w~�ř�5�{�N�3Ƭ#b��?a��9��K��
� <P��� I���"�DF��?1Ο� � 	ތQ����`���.����t1�'�,�IL���<)�%Y9I�3���yv�ՓӬ}{@�I�O褥OB
��>q����/�d��YҤ χZ���c�!�J���Ot!��h����p�x��� c%�59'�<��E���	��..��'R��'?��-H��*� ��l�:$W(���W��'O�TB��i�,k�:M V�0g�X2�ۏ
��Dӆb����i%�`�Ot�lZ�D7�1hb69be���E/4�ʓh�樧O�DG�TM�q+�Y+d���O�V1-�9���	�6܊ӧ�9O8Q[u�����ʃ9'z����$L��커)Ɔ�<��'�*�*"�'Qn@�O��-��<O���
jG�,s�Nu��	�'T��IM�s��CbD�����.[|��/ƯsX�ۢ��O��Y
�����.Ԋ�8 �F�A78�(��*���'	�k�d�v��W�6,m��0��Iy��'��T�L��5�#�7*��y#HG>`~��#�R+�Mk���d�O)�On�^>Y��7I�����s# )�ŋ�)3�X5#�4��d�O��������0q�	���U�{�6m�!� /Q}╄ȓi݄ѫcы׈A�g�Ô;��؇ȓ	u�%*B�]�H���[t�ȇȓt�����FH�8�����h�ȓ9��I�jJ�P�����U4�q��q�����u2�`uGқg�<��+͊��2,$��E}��ȓ:2
hPӭ���:��7l�
'�^��ȓ- �ta�G>	�,����mOҭ�ȓWp��E�:���Xb�EB�Gx���_���Y��	�-n]h�
 �}�y��_:!�!���cTm�bXw�\d���&��O���*ɦ(���2gV���H�a���@c��r5�Ʃ
���F������U�g��A@���ru|8���+����E�>|K�A��2�R�Q�X�|}r���y� �SH��ds����Ң}�&xǏR�6� �a��SI��ctjM�J�н���ӓSdx :U�i�Z�ؑ��+҅��Ćr�d4�6�OL�$�(P��)WLJ_�|���4*W㛵r�ҭ�reݯ�A�x�a��mr敺��?P����I!%3H�vf�*@���S+b�,��_|�H�nݎJ�O�����'� 7�[æ���m�'58�S�FY��ۧ�]�x=�=�����<I�	����d�P�<ޠ|�wcIN8���򤂘t�p����R@��e��"���A'�N֟T�IԟxkB�ª��@�	֟�����I'A9RQ���,��D�@�#��}�� 
6Q�;�Bqr��N�"-� ��IBy�'C�	�Vl,���/���*%�A
� P(����*[��*��:)��DG�^�e�8#�X>��P��yǃ�j��<iD�������G.�6|<@l���M��)p����S�gyb�i�L�
�V�V��a1L��v�<9s�"$��ӎ�Cf�Qq�ȕ4��Я.}�/���i�<�A��^6L��%���S�*X�3�ϟI�$`�P
��?1���?�;4��O����O"1�s@��;#r��f&��^��}�@���:f�"&Ƞj.퉦�Nx��	� T���T�^����K�<��p�cE�+߬���K�*Ȣ`��LLV�DF|R�۞H܂�aT0_.q(�Q�m|��	��?��iG]����Q�@����?�䱓&(V�����hO����O�O> 0��M��Je%Q�_".)Q��CBy��'"�6m�O��1�\�S1�iFB�i�ȉ1t#Wr���v/'��	0/�OR�$Κ�Z�d�O@�dׅF`,���<	�4d>�I�Ů-b�Qд��.�P�剧mB"�23��<3"!�

")fr0۷ �~t",i��T>��a�˓#��|�I�M��O����	>�BP
�K�|[��>i��ʰ=Q�B'f�Dp��㟐���r�A?Ug2�'r�II�����'c8.Y����8�pW��3��'�剞w�j]ޟd��O���ݓ�j6���0B��z�"�-fB�����N�h��I�ZR`�E��ۗ��" .f�B�S�tY?%b4O˚R<$��IN�[[�!ڔ�:��Y�i�n�BE�Ͻ`�$��l+ʧ{g�x+c�-ظ��d��L�l%�l����OB��*�'�M����K�|�� ��p��|���(�!�D��&��x�@)��f�i���0r�x�=ʓfh�pKQ����P��(C�tn�a��oӈ�D�O��G�5̀]���O��d�OP��w����vMA";5���u/��9�jгT.��{�ތ0��m�p��Î�&|��b>)��O����?k6��#IB�Z��ѫ�
�eb�ͦ
�̰����*ӱ����'^f|��^�֤�Ӎ����e�O��"'$H�i>Fz�*ɜ~CF����-��q�Q��1�yb��%��u0�-!�eR�!���HO��O�dPn]@Bg[����+>;�@�$A�%萉 �'�R�'\�G{ݱ�����'-&l�#��֝[�t�2�`��V�`�{4�%D5*a���yv��d��G�Je&i��Gr���;'Wj]��)Y�q�zIJ��p=qfg��a�n�@�ߋ
+V��#�YzV|����MkF�i/�O�Q�}�`%Ue��P�1�I���Itn�a�<a��
�2��r��v�h���^���Ip̓���x��1�G�Q�b����7
K�����hOQ>� ��')��qJu�݌=x��bTC1}��'�^��+ԨJ$J�С��N���'FƜq��%p}���qA�5����'4�-;�0��h�`�
���'sL���cԁh�}�J�'Y��;2�ad��"{
8��b �y�G.2B�E��&� �~�B��yR�̵}��Iw"]�/y����mO��yR ڻW'�	�6ʉ�%��!#C"K��y���ĕ5d�|�$�IC��,�C�		l�.�*L]�i��dY�CR9<C�	�2�9�"#�HX��:��� <�B�I%�쨛b	�3��t���(`�B�I�N�����E�T�#�T#+GrB�ɬ��x�`G'6@\�gӺ^eRB�I$ClE:�E��N��tP!AĬN�XB�Q�X0;��'lx�ԅCW���ȓNT�����/wߊm����IN�\�ȓ@��x��H�:lR�#�n_4k�p���""�mJF`ٛĴ�WJ��
�Vm�ȓTW̔C�+H�?CQxa�ʧ>�Ɇ����q���쎩�b��#[����ȓ(7����B�K�T8R𧆛���ȓ? �����Z%;ixt��XҪl�ȓu����Gg�
���㰩�p��؇ȓ�(YE�ޛx?�A�Z0)ȇȓt��jvg�����R��&�x��K�|����)���R�M)G�)�ȓu��ɳBЎh!�j�@=d���ȓ^ZB��AZ�L���Ҡ��Zja�ȓ0�*�'�×>����)4~��ȓ[����e,#YzГ ���\`�U��H~��Iu(�%;0�33.I�f��ͅȓZe��cԫʲA��˧*�9���ȓkgF@zE�Y�����=Ob^X��@�����!ʳqH��!V�b━��S�? ֤�&����5�0��$+0���"Of���Fߐq$i�p�B� ��G"O��P�}��s��p�!0"O�<Ad�Jbh2�!q-_�$�x��"O��bDL7eR�Æ�@���2"O�:QIE	C��c�������T"O\��A�L�R�>5�3�%5ӊ|"O�LI �V�?��*��H% �.%
"O���vEv�P���	
o�<
�"O�� ╰;~�M��M����9�"O��õ+Z*�`���D����"O���ŀ�E�^U���Q�lE��S�"O�� �X>$%ʍH��8oі�1"O���.��(��p����
�@1�"O���n��`�ݐ��B��D�R"O6��#I�,R�*<[���	GD`u"O��ԃY�)t�;c��1�V��"O����N��%�0&�^q��"OfXr-ƃ;��1 Yv� ��"O4(�J�{����OX��"O�k0*۴l>��G���>�H�"OlAH"J��|����ϠX��"O��!���0�6����
�P�J�`"Ox"ǁ��V<���FЃ/�fh�`"O�p��aV8x��\I$�'��e"O&ix�F�m�l��"����l�&"ONh�⦝a���\1G���"O�yc��ֵA�8`� ��Y�x��"O��9�B.@���/,���j@"OfQr1Έ-U9N�S��ąI��T�"O�e�a�A�'	J�Jq,+�^�xS"OP����t������LJ�r�"O2\���{�ذ�ր��Y��̫"ORԢ��ɴޮ�8Ď\{q���s"Oʝі�ؔ�n�¦.ă5��,��"Oܸi�`�%Wj�Ah��,�
�K "O*�!�a��-k&�2y����"O����,����J�o�/a�)�"O�U����8:�����.�@��"O��xk�?U�LY��qFZ��"O�4@#*��aJ�pJ�JU)�ZR"O�@�#cTU]��CԈ�4G�4xW"O��Jv��	��H�0}1���"O"�9V>6	�2��%P���"O�� �ױQ)ĥ�G�P6R�ZL�Q"O��2����4&��梓F	|M"4"O�����1 ?�XE����	hv"O��w�Jmd�PlE_5B)W"OJ���(��&��u�@�"OU ��>b6�]XӀ�:'(�c�"O�i��E�]�|�j��]l�و�"O��ёnK G�H40w��,�"O��ŀǋ�^��B	5��R"O�����
s@�+AG�"a>���"O�qI�-�,��fT(QNN�Y%"O45��\%YG�IKwe8[1��"O��BB'S�P!³��;p��4"O�����
 4���eB�	,D�S"Oj�'Vad�#Gɻd���	�"OX���A*
G*����[0��b�"ON��м&�t���O���p;'"Ol���l�eL?xR��3"O��i4��J�D�:�D�df��p�"O|Ĩ�̐n�2 ��^3x�d2b"O� �dڣ#I�/gA QC� 5�аH�"O�	b�B�&}�"�M�R�D�J�"O�m##A��`��n vLp��"O ���&�Q�	���Ϯ4_�ɻS"OfL�PBי9��Sf��#*J� 4"Od���;��l�l�q���0"Oؙ�#Ľg=�0��`S�-��
5"O�ɸ�=S��I��!
ވb"O��h'IP$*��pM�*[��y9�"O��Y�k1�i	��W
iIީh�"OhhXN��n�ڙ��#F�ن"O�{R����=�pkW~*,ȓ"O�����9U
tѦ�0w8���"O���D�!%��! b�<L��QB�"O��/�
}��9��G�\��`�0"O�L�p���3����!�xxP"OF����s<P��R�Y#c�t1q�"O(q�o�u*\I��D����"Od�@�l�zx���mQ�)�[�"O�}ڲ`ǝ*=RE���O���!Q"OС�� �NuM!��!p����"O��v.V8��m�'��u�X�s�"O�0�Gl���MR�dKT�� R�"O4�)t�Je�͸�F�"�<�@6"O`���7+}��A��:t�a�"O2-��j��f�uiJ�` �&"OR��׎].+`ȅ0�M�b3����"O�ɚ���$Z�
83���1,���"O�L(�d#�� ��d�l�k�"O��0�FחQtZ���M2N�"� �"O ��lL-=�^ePe,șFA8yH�"O��0�E�5Tp��JX��	"O�!	�+�8�����GO51�h��"O�r#Y�Ԩe�ɢ6�:�xV"O~%��.:`�Q&�2�̀Y�"O.���X.7�>-kE�D���3"O����#�����dؕ�`a"O&�rS[�e] ��2����g"O�T҆J�:Q"��ͯj �D�"O]���ɂh] ��B+VD�"O��cj���9�,҆#�[-�!�dLl��EB-����g��!�W�$^X�E�[�2U`� �T��!�d?^M���Gُ?�PpA/�^�!��H�gqz
pLܚ1�8 ��l@�)�!�d�%C� �SIL,c~��ԫ��!�I�>���$��y>b0*W �.�!� 2Hy�薝@9���m�*i�!��	������wL�0d,О�!�˪&|��5�G,a���`k�_;!�V&$�l@���3�0-1�j�!�" �PY*��Ü��z���&c(!�d�M�=#A ��}58<C�)�,U !򄈾Wݦ� Q$r���@%$�!�]�� ̢��(�i
�g�i�!��7Z�Nd@�!���ـ��_�!��E�0��U�cK�<\����m��E�!�d��F0T��`�H�I��'s!�$U"
��IH���b�m�C%޳N�!�DP�"�B��`a�u��=[��<
!��Dp9p��Y�k��k��S�T!������R��D�H�z��Eq!�$:v`mb�_-3��|����97l!��\�2��b��%p��A@��	�kH!�� h�	L�e�@���Q)���"O*U��C��@$p(�ܘ?H��`u"O�&aB��Z�4O�y_0���"O��`�C��/�p9ɥk��:^b�!q"O�$B��xA����(R���"O���KɟC�Xe�ƐV�ظ�"OٻP,�%���PiN)^�"̃�"Ob�����-U��s��SK�^��"O|� OV }[Ta�OÚY"�0"O`s�/Q[b��B�f�:���J!D��KN��p�I��O�D���cl D�Pۡ�F=
��I���̭%�,ZC�0D����&��P����+y����(2D�x� cϱX�ҩ 2�:z���0W�2D��
Q`ȋD�Lܓ��Е��UX��/D�����&7��Qd�\.y�i���8D�Xv�j)����)wy��L�!��%�╺P�ðp�F�2AL�<:�!���&�1�voP�^�ryEF*0!��$
F̣�D�q��u��HY�g�!��tl5a�ɑ(�ꍛ�GV7�!��R�_��ӡ�{����2��f�!��8fݠ m_"Yn��ҧ��!�dC�7�)W���?E�����w�!�D~�,��F�W. ��x�����!�Đ&uJڜ���x��x0AFB��Py�-$"��rC33J,��C�'�y�`�Z�@��SFAz�|��#���y"(���j�bE�
d��c .�!�yr�gl��AB��`���wfY)�y��Ѭl넝���Q-W��<h�L�>�yR���T�'$Ȟw�~��A�Ӂ�y�-��:ޑ�"5'�&@a���p=IEɁ�)���Ej��,�jbu��\��A�/��t�|�z�I,D��1	P?#Yd�xq�ۧ_$�z�$8D�S1,}�(���I�8lƲLA��$D�XB�@�W=34dCS���@ê$D��RH��g���6�1��(D�l���Ѳd�~] 7�-vl�$���*D�q+�4鰨I�W��*~���@	�'��s��O�Lg6��5�,unRi	�':r4E��{ ���q�4���'є�7�P�ܼi�a�n��p�'�de�I	. ���ń^�a�.ū�'9
-���,[xp"�
�g>h�1�'+�5�-�
v���S�j>V03�'�lLP���!�,�%_�����'5>E��,\-w�@��B��v��'0>|��	�ph*�"��Śs���	�'�"��U�D6Y_�X��8���	�'R\����:4�� &Ӿ	��p	�'��7�J�P�H�"�I�:�02�'T�Ӥ�� �m��.M4"pt��'�t��$�(u>a���ևJ����'�t���hB�g�����i���,��'8:4[�Ե%~���U5`h:�'p"ȋ�iI'���P���98,:Y0�'s��,B<I{�\��h�0XT{�'�|�r��q�@a+��#���)	�'<�ٚi9Sg4\�0$$�ĕ

�'z�qT`C�Xn�Y��'L&��X�'s h�HU�jq�ǹ)�����'D��K��4)X��* '�=_4����'�"M#�ED�5����oA�^N�]���� H ���ĎI�ri0�8L�l���"O6�H�C �N��e��6".$�P�"OR� ��� Q��L鶀Y4�4h"O*�0�Z8 �Du�a�5UH ���"O
��Ϫ{(4��@�HX	%"O�%)tk��8��ѷ&֘�EC�"O����dֺz
�:�@',Z�"O|p��/X�^�a㇟=�jr"O0�)�j�(:ᖌpb��c6�KU"O>-���1>](1� <
��"O蔫���9q�~��F-%rT�p�"O^�KɄ�@�x,9�aX�\�$08�"OԈ (z�2�"Çڛp9��"O\l�1�LxvP����%q��iKG"O���@�		�Q��Ō��`Ɋ�"O
�R��5c�&�����$�r��"O t1�Kŝ �<\���Wt�U*&"O.-�B�Pc���ŭY�G���"O,l��DLNvĵQSj�v�lL`"O��#̭B�Q�pƑ+S�6`s"OB83����Ш�٥��
�tUi�"O�a"wϓwg��y��ܯ$84��u"O.@q�<eC������|��"Oz@�r����&����Y~'"O�����N��LH�G+s�4��"O��٣l��S�(�@R�ԺK��E��"O����,4��)E��l5�S"O�C�	��p��i� |��w"Od؀�㖓rl6̙G�*@��"Oᑣ�Er�����У-��*�"O\ԈÇ� a�H)8F'��D����"O>�`�%�)qG�4�%�%"O�Œ񉝷�Di�����Y�u"O�)�'�UdF���΃�UT.��"O�ɳ_������*2IJ���"O:E nB
��I��ΑJ���84"O8��G�K7܄	�@n^/f��{�"O $:5��)34�d)s�D���p�"O\���BQ�8�j���j���B"OFi��G�Z�Ƞ�-_
{��i�"O�ez���@�4��c��x�Q"O`�b@��ʔH��OΔJu����"Oԍ�c+�,$�Kw��sV+���y�b��af�q0 �=h�̨cDά�y�"ÓA���B��h]�Q���]��y��6}?N� $�8J���i�͞�y�M[ d�T��8{�ʁ ��_��y���@n�y4�@��a+��yR�U���ă��rN\h3���9�ybh�O�ZX�A�(���R@[��y2*JZd̳���ɰ�XR���y��?l��P�T"�� ��p�զ��y�� aI��0Qj<K�m3��y�(Xz4�2�-�:0N}J����y��܉.C^ə�"+����Ȍ��yR��$O�� ��#}x��F	��y�e��K��)��D�e�hLȳ+O�y��]��H�DLS�0��D1�yR��^4B� ��!Hڰr3"Ǎ�yb'RTzE6ʜ%B�n��ݒ�ybm��ĸ���D5~�Q��mT�y�H�#i&Lis�"Je�quH���yrnY�e��ݛwF��dAP<�$)���y��	uCX�Z&��``؅�Ɵ��y
� z����M:l�.�K�$�7?[FqHe"O��ʕ(�
+6���@�E�V�Yw"O ��ƋpM���C�3c���#"O�e��FU�&:��gE��Y�8� Q"O�0*�K�g*���$jI�|�^!�7"O4�6h�_�"YK�i.O�� h�"O<�x���0׸�UJ�-3b�aW"O {�뀁o�`�(�)TL+�(�]�|) +U��اH�>�x�Ř;��ȓS��P'�5��"O�5�0V�u li3p�ϡ���a�����b���8�C�@N�@��A�R�z�$��;Ќ��I<M��1�U,=�@Q(��h��,ܟM�ɻS�£�xB��*~)R��pM�W|�^��HO���Pi�T�LX��.�Ķf`����[B�FU����$f{��ȓ�
E���$R�=���O H�\)K]~"Ȃ�Q2iO�P�/ �MG��'����G�$d��n�pîx��M�̰��	H�`���`�߼�p�iV��0a���닗����dS��� D�9e��1�㜠��{rIX?#��H�fC1Vu������ä��%� 'dY�	oHQ��I�~�I%ߩj�0�!r)هO���?�T�<��h�"Z�U�`�G�BR���/X��ؕ��$f����`7�!�q��a쏎=R:���'ǂ6���o�)]F���'�C�J�r-n:ҧv`��<T^ DZ�4~�Z� $ �a�!�td*!�[O~؂FD�o*�oZ$ �x��!�/P�iX��}ݡ!���T����)��Â�n�ڔ!�X=a{��̭2E��W��p�y�LW��8�$��)o�R)21e�wItTy%�#�O 4p�"tᓨ�)D�hb���Z�O �D�&@���
Y�$�b�z�Ο��ZU�G5bՄ峳��"pDQ�"O�`x��ĴGfD��*	a�RA��GxNMy�hV�y>p��nȦ#}RE6O^\����s�����GBRT���"O���RI�{���Hfʄf�y��EY
)e���3���$&Lyb�ā	��N:�.���A�e�h����h�t���l��0��A�V���;36o�����ʵ�bt�Q���s�@`�"�<�O���b��Q#<,¶n(������}?�f���<-��fH�
P�Y+C  [���aU֌3��B�I?���u'Ʋt��5��n���I�{�����퟈I��q��h�f
ץ�.N��(��&=����Q"O<�i�!	5v5��NnQv���3?iR	�Z\��')$����JD�t�Ղ'�2���X��0?y$U�xD�UhGOկ)F(�2 ^�eZ�;u(�6tT���9�苣�E+
����;?�,�D}�+��x�Z���&:�Sv��*3�ED�d�u�ڭ3�C�ɘ{�Z!��$K�pM���K��I�Ur�M���t�)�'%��D�gʆ16HXqEG�X�̕��@dR�K�B�>�(2���R�&7�'��� ?��۴gJ�B6�,�B��[|B�IM�e'(Ki�DrN��|Y>B��Rސ���D� ��l�Pj�d�B�	d�M0V�d5��h�T��B�	�0���Ue��<2jmR�#
&�B�	"w)0�seT�Lx�mb��V77I�C�ɡn���J��K2{���˷H�<"pB�ɷF7�9�D2��qB$/A8^B�ɓKf������%WL�i�$l��@�TB��U�"!�p	_�t��q�'�Ʃ}^$B�I�=b�K�c� )5@`��C�9"B�	�8�*al��\��@oCB�i)� ��AO�\
�)
	���hf"O��cC���A �����Έ��"O<$�ՁB�i�H�q��<�9"�"O�Ik���F�p�õ# $�`�"OFաҍK/Z�,�ʱ�Ɋ5�C"O�9��A�\��	�X��i�"O���$e(>�&�{��S�B��"O� &5Q�HI2)�|]�2*,�Le��"O =�Δ74����ЮWVT#�"O쉓@��U�4����[��C�"O�u�%��&H;�x���,�$d"O%�A��Q�B���\�(�q�"O��:fmÐYt�p�H�&Ey�!"O��sRG>	��K���'��y�"O�pˣ��5	�\��ϗ,~f�["O��������ڡ�e���"O���JڎN���еgH]⤠("OX`1���~�Ch��tm��g"O�����c.|��`L�~T�a`"ORHè�W��, `�݀$٨��"O��`E�)g�l�'D��*�|��W*O؀r�`��\ ��R`G3;<LK�'�
��T,���5(�\��D�	�'��1�� �e�ՠk!`�	�'S�L�`��7dY�@��R�a"�8�	�'���y��[2\[�9�6��"��5i	�'�ֱ��B�^����VYo"�	�'�zm�'�����Յ�&BH,��'��ua�L�\}����eL7�6t{	�'ӲA�Ĕ��8q� ��	����'*�Cp��;A2��&�(=pP���'7��%��(I	�M�?"9 ���'dt9�P`�a�t��Ed�]���':ܢD��-���w���(N���'��xb�wi"��\�z�� |�<�6�V?��!s7b���U"&�Uv�<	f �mH��& J,Rd��r�<��iͻ=�$�;7A��`-��s0G�W�<�q+�YN�l��F@!S"Dh�g�N�<�j��R88�\�?�� �F�<颋��~vt�B�X�������@�<�/L�m8la�$�Q�4(�#��Y�<1�U ,D��!�TDo.�D�
X�<�t��!�p�� iIejZ؁� �[��H[C��66 8	�b�-JƠ峦`ޮNJ$͹�"�0J�F�8�"O��ӊ�FT��fe���;�"O&���٦3�fq1<$x��v"O����{�����N�@
��"O����Ԡ;��*bM�5Z6p8"O��W��f������(.�xv"ON0(� 
D���m�	"�R�"OHcb��_E�y�B+@�	��"O
�z�L. |�Q*�J�1R��x��"O�Z��J�mđ9uoG0:���"OP�7��N0ȩX0��C��X�"O�<*�gU+D�1P���/9��H+�"Ol1[��?[�)��C�7��C�"O�BE\1�dD1��(H�te؁"O*(�$	�)D�Z��pK�%w]�=�F"O0�y�lO�k=t���
�'JԽ��"O�497J��`�݃���4g0��ۦ"O�81�m�!)#g�)-�h�"O�3P�T�V9����gG�2��y"Ob�Я�-���bh�/�\��"O�q�T�	W,���g���j�"O��f�SJ���[��7A^��q1"O*8ؓB�,k�����T3�p+s"ON�����O�8e� B�0 V"O�%R∛7I$XE�'cD"%�mS$"O��%f�Ud"=��]��{�"Oh��b�7xK�k�*?�<�"�"O� &�� �A�Ġ��/ժQ��p"O�LZuk��5^V`�&O��t��MҰ"O~���S����@�\�u��Ṥ"O�ٺ'hί|U����kɻN0�"O��X%�N�&{�(���Ƅm�t�+�"O���D,�? �$��V�Д=� |Q�"O��6� �&����R0u�#7"O.|�L���1C��F����"O2����#f� lʶ#����"O�q%=�q u#_����7"Ox��dG���ԛ`BA2z�d�9V*O�`�ň8W4���(>A��Y�'nrX�f;Z����Ç_�Ġ�8�'<�=���/H�ؑ��R2���'/�A���;>�m��BI�~�N(
�'���W+;cQ�����pv�a�	�'�6ܱW�)Q��DT�J�8
B���'9Y'͔�Y��dIv�%!��;�',6%�'� Lb��R��o[���'�P�1�B?<����M�t�\-��']�	�8�3���z\�*�'�D�1T��y8��!�Le�����'���;ԢO�Y��x���$���'�(�l� l��Y/6��a�'a���E!C��Hɹ�B�&(����'8�5� %�i�Е��"��L霑��'��q���$v����dۥ<t�� �'��XQ���4m<����$e�:�'~u��/܊#����ZD��'�Z�S�L����cէ�'�v,��'K��������15怖/�i��'�B��5���c�����K,l�`�'���Ѫ�.UG�[�j��~��k�'h\h8��G`�X�"�K�q����'��}"�ߢlx�$��ě�k~�(�'l-є�L$F�d����f��y	�'���IԌJnu�(iQ�ZY�4az�'^d�I��tk�P�%e��b�ij	�'1V�sNF l�xAvū,�H=y�'�4L�]Xp���T_V���2C���y���e��ݢ�XP����	���y���S�RA��JB.E�lI�����yBj�=_At��E�D;�u�L��y�J#dq4�@��Չ0�ݨ��ϑ�y��av�9�%�":0����
7�y��S��ı�)N��L��ƃ��ydQ� �,%��$S,��f[�х�3�&��A�W8wR�)���e�
Ѕ�!�v���3a�(�)�H(�ҭ���`�⤃�,j�`�e� 
�ୄ�?�x���6N-�	X��_�D׊0��Vtݒ�A]3>W�Q�P'֞Kp�q��`>���vo�
_Z��@ �F���@#�����G�D)����ȓZ��(��l·M�zeg�D0"���y��4�U��	V0���R�� =�����{BI�K֭?Q�M���鼙��1j�����w���񦆗T�H��6&0B�c^hJ51cΏz��H�ȓYv](��3w��!�'�;$��b�4��T���\V�%a䂭m}ę��4L�;B~�$10#�=Cڅ�ȓ �b�Y���4�Lв��
0��ȓ2ņ��qg
e��I(&�
3@�̄�S�? ���c�0X9`�a���T$� �"OP�K��
�L�$��K�8	��cp"OX���F3|'r<a���1,����"O*���b�'�fx�)����C"O&��L?/���2T�ή!>0��"OJ��O�6��x��a��Z\��"OܽR��%V�����B݈?�h��"O��k� چju���'
.,��"O�d�c�
tx���T7R&�M��"O��e$Wo�l��jݕ5����"O��h�/Q.8���'��Lx�iS"Oȕ�JM�~8����?"���"O��PG��A`'� �˲(k�"O� ��� k|�qI�S`�"R"O��d"��^��ͩ��7K>�0�"O�L	cۍ,�������l6� �"O�lҰ�'8|ٙ$e�9]5 �:�"O"t��f6l�q� �N�h�"O80@���e��ؼR	ȉ!�"O@8 �_lhx*�l��}��(��"O�eS�͙_60ѤS�w7Q�"O� R�A�h��:�C�b6���B"O�8!�j}����C66�T�[B"On��@�[o,�2����8p�"O�y)bJ�����э�57y�Չ�"OP�(��7Q�nuk �ݡ�&T �"O���pM��;t�S��х?����"OƝ�7��2�H���,�h@���?|Oft����,5�X�x�J˅̸���"O���3A��R��"���.a��z�"O�1�&D����C�ӵ)2X|1u"O�mh�I�.uoH(CH�	$Xt�"ON	��L��]�pHqt�M�T�UQ"O��+ ��,DFXX4 ��	��ݪ�"ONx��L	r�Z�/֪gJx�p"Oa���\�1*� ycDCQj����"O(��eI%��-����Z��X"O�8k����&���E�"�U�s"O�sF&�x�bA����u��%��"OD�X��0\�� �!�T�6�S"O`d۵�6I�$���A[;�ԩ�&"O�\R�i�w(@�� -It�m��"O�����v�H|JQ�I&ld%�R"O����n]���[���*�:�1P"O24@�H��2�T��h^��i�"O �zG�\Xh�r��=8�n�:&"O�y�#� +Z}[ul��6�u"O�1z�bW�X4�r��-���"O�u��
)Τ����4�.�"�"O$�22 �+Wx��	�1v�R)�"O^W�=bИ7��=J�F<kv)�\�<A�",NR��n_�����Z�<AR/N*R髢�k�|���T�<�!ިlI���Qf�9����P�<!�*�ҍ2A��P{h(��E�<IfXfˢ��Ofl�	�#�X�<3�s��|�uJ� RB(؃KQ�<��N�kw��@Ί	d��!�UP�<ٕ�D6k��8g�H�VÒ��F�<��#կ(*�1k����)� �[v�M�<�RA-�T�A$�//97j�}�<q4H��zJ�a�����@)�@�<����1}��ك�
ƭC�6�2���x�<qGJJ>m�Z�H�+����q�<� !,]7@j��"���x��"O~�S�HR?͐ur���rF���"OT02d�D�*JL�Qϕ�%"�Q"O�� 
�A�>���7����"O���F�:& �%��f�=��x3E"O�Pd�����Ӣ��#_q�Hj�"O��{��Q�@Қ����9KƄ��"O쌣�7bH����.�#m�A�r"O�}�D�)X,�����
'0����G"O�� P
Я5��X�J�lq���"O��yL�A;*�3p�4lM�c"O.ؚ#m�Es�TɦEӱ5S�1x�"O�� ��_��X8kt%��>�, �"O4��6��^�<�#1_�A���(�"O*�I�oJ&.|�YS4���@f"O���V��j� � s�(x"�ۤ"O^̩�hY�8���'��m:��"O���ČֆK��5�M�&b$k�"O��2G$�$YI�ʁ�,y�QF"O���"iR/��10��	]oh*S"O�ظ�
���H�2Z��Сu"O��� �O���ܻVdطW� ���"Ot)��"Cqu����nq��b"OfU��&�,
���u�7Rb�r�"Ol���Ȉ8�`Be����`�"O���aJ4t`5�#�	\�`	r�"O���kķ������̑^�6���"O:-���]!IW��8��L�^��"OV0
��?M"�	g��W��$A�"O �ʖn]�L�|���J��.qf;�"O:�I`kH;[l@i1�޶@^�p3�"O��R��F�f�P�d��:Ct��"O$�c��½xn��k���g)�X��"OXԘ���*�@�����r��0Q"O��`T�WnjU8T�X "hqr"Oȡ�@�ֹp���ےE@9�.��"O0��4J�;jY(ȳ��A���s"O4�b�ǔ)~a�11)D�U��a[�"O�%�@��Zh(��w��/N���w"O:iG�148��ӭZ�i����"O���q�� vMD;7C�	3NQ�"O�XKD��W
J��@�B7L���p"O��	T	[��	K�D�Mshd�w"Oh��C�#yJ�5ٗ�L�npܼ�E"O��'k�;(�̄�O��dA8}�"O��)kƢ.��!P�_ ;�T`�"OƩ1'��>c������d+!�Nk}�}��f���N���ݽ!�!�?��qo�@�>E���!,{!�d�1X2PL;��L���! �kδiP!�DС,�!�#g��7΄=�țp�!�dV0 �L�T
�Q� aF�O�a�!����z�����L�\�hS�9	�!�$�`�n-�trO�J ��Mx!��=r�:�j��UH�l�+Y4vr!�]�[�r�ޕw�Nѫ!Dԧ1^!�$N*W�bL��=|s��뇂�[S!��1��|��G+l�&AS���G!��p�hf�>*��D�Do\5F!�$�<LQ��*�>)����6���=�!�C�:���" ̑	#�\9�l��C�!�5^t��lX�N���J|!�D�~��Q�V&f�@P9�&�?�!�D��*k�
K�B$�4��E�0�m��S�? j)A1ۢM�(�93J)2D�Q�"O��8�J-�L��3&�(P#jx��"Ox*ŏ�k�tŨceGPz��"OB��E�DD���cC�R��P�"OV������/��\ �aP�0H�|
�"ObDp#f�3,^��CR 2��s�"O�� pʅE=�hC�(���`�G"O-���uL��9���QÌ��"O�)aW \�wΆx�D��<��P3t"O�H�6���RC\�����"OF�� �E}B8�B��7
z(A5"O�)�P��
oT^��Ĭ�H�"O�Aˣ+��^��@���
�سw"O�V�+o�Xci	���5xu(�K�<!wb, ,�![�o҂h�,ɣ���D�<���>I�����N�pR&�����<q�
���� ��6]�DQ��n{�<!��>������ꦝ�U��m�<����,6�*������<��l	`�<�a
�sf�}�g�H�pݲ����U�<�����0/4������o��S��G�<q5�I6��E�נ#d�)�7l�E�<�Ddڼ�8Bd
 YP��+�$�G�<���
.b�K��әO����!b�D�<	�N�I�s�*P�e�
u'�C�<�B�1y��U;��'Ѕ���}�<q��PIj����V�&C~m��Ha�<QѪ	����z�O�!q����CZ�<���+.���CƋàs��reB�^�<1�����q���, =H��M_�<a��#sN����pl�4��Ie�<�F`̱S��dΙ�z�(@dHBb�<��&S ��Ɇ��1.��pF_�<��r��x�7��a)���Z�<���
ay��P��,������j�<ɵŚ�E��!��qJ�:!l�j�<!")O�U���p�e�I��"��j�<a����� FOD��ǁ�c�<ɳe�)<��I	f��=�htJFe`�<Yf��5o���)4d͹[}*\�C��Z�<Q֢T�1�b H�o��=���3b�N�<�sD��j�85$C�H'��x��I�<Y��T��朹w��F{5s�NH�<�g��HH�m��ȡQ�`�ԢL�<��,��O�6�Ho[����H�`�<C؟n��h+d���$��i�\�<qQ�/wY�d�v˙4�W)N�<��P'B��X���ʘK�8��@�d�<1�gW G �
��ϕr�v����a�<����$b� �Į�T-ΥQ�FB_�<y�HN�2��0�#�65z5�u�[�<��K(��"D�˺�a�Y�<o�T�,�7,A,upY�
Y�<��ȟ-C�Biާs� Q��Q�<a&�-���7�#%��� XK�<!�,��-4�)���6��q(s�E�<�gQ>L[����a�9c]@��D�<)���I�0aFË7Zsn��ရX�<�R�q�:d��K�4{\d�t�DS�<�B�H����u�2L؍c��\M�<a�k���ʙ�ȣ���!1�_�<ɠo���0�Lx��qi�k�[�<y��Qm:d�� _�=܌�C�DT�<� 
�D~�d힦�	'��L�<� ���u�;h���	ޘq>B�!�"O���ďkN�I��M�Fנ�r"O�����X��Bg,B:8�Ȱؒ"O=@-�%mwN�� ΜF�\a�"O0=��H�vkx	x�`�tTf��`"O|ɺa�ׇ_��!���C9Ψ�"Oj$���M�/,`����1��JS"ODx���>x4���[���1"O,�!��!%���B4	�m���'HPɓ��_Kh. ��z����'��}�(B� D(��ƫJ�ADl�'Z��{������ɲzqD|!�'�^��0Aܒ��}W��oH�(�'+�����+�>Q��fZHA	�'
�����;/���6�ҴY{�i��'B$+$Kթ(t�9�Ea^}��8�	�'���џ@��}��΂�B8k	�'�����ׯ\����Ӛ}1�d�M>��O��a��\���.�:@��ȓ�>�k�c��jrܭ�2��YP��ȓ92|p�'��6p�<P���/$�܅ȓ��#  ��j	pU��*k[�̅ȓD/dlч�Ƿia�+�)j�х�U���C�M�Ly>P�B�O�\V��vlv�C6mK=l(8��-���Ʀ �GHH�$�3�a�"�"X��>�* h1�E��}�}�ZA��P@���A��c�V���C�a����=�����Tm�u2�����$b4@����y"j�/����&JF� �*�Pc���yeݭ-hd,B���(�Α��y��דa��Ê�S�L|����yR�W��n`A��7Z��jw��x��xӺ��׏-?q�Q�f�A� m�"Oܑ�U�C�d�*\ڐ$W�9@�8��'đ���@I$S7B�J��ŕ[i0i@�7D����@�/���b���� L4?��)�'X������+F�J0�l�s\���ȓ
tй�C��z]�m�MWJ�4�ȓt%n A��mb$�χ�"���:ъi9�'��Mf�G�
���ȓt	0��ACڰ�X̢Cʇ?M�$��<Q����(�<Ek܌��f �c>��ȓ/A��2���nXh�(���i�V�ȓ4�20�H�O.��(�j�/�q�ȓ`2�@2�-`�MhQ�P�m!�T�ȓ	A`<T/�5,��<���Ǡ31��ȓxfIE���p��B	� Y�0����Z�Jw)��T���PG2d���I�}�����.0s��Q.V.T`��<M\��B/^;Ԙq��e^&	%�ȓr�\��)Y�x=���� W�J��ȓ_� 1�nB ebyx�I�+s�m�ȓ�́ ��m@x�SuEJ
*Ϛ�
�'1����e�e�mڵH�4�]��'$T各N1Y(L �/� �8Z�'�fx��8��lD5.�P�'���
�-��N��{s�܋3_�;�'W�ݡP�S�adH�*��\�,�\B�'$<���FW6و�ӬW��p�k�'�ĉB0�J��r�����x�'��9���9o��]$�:cT<p�'�@����D1j����ׁ3����
�'�а%d�,xn������#n>}�
��� |���".��ԥ��D>:��S"O��IF-	�[�䈁�˞k,0d��"O(Ѡ΋(*D(��]�F�$�"O0\�tl�R���R���ar�"O��%�-CGv�a��RI��"O�p�&�'�<#R[�!��,�&"O��xga�fN�����o :4�&"O��q�"]�dd�ٚ�lL]���B"O��0`�ǹ{�\X�F��d��[�"O��Љ��7@d�B��,��x2 "Od5;B�y��}��ͩR��
"OxesQ�Ǖcj�Ыd� Md��!"O�@��(�*^��Ĉ�����trT"O�aD)���b�ڥ�(x��S"O�ȑ,�?g���!Ï7ZtIPU"OR�
6N��c0�#:<򭱲"O�y�bǗY��Uڅ�~-I`"OP�7��h����ˆ�6�ey�"Ox��� 7M�i�H���)�@"O>d��#u20�cD��/�$)i�"O^�J�bW�#�]�aՏ����"O����j�t��P  �}Ң��""O>�C�� aB-�$i�2D"�#'"O�Cl��$��i9 c͎���"O0Ѥ*��1�쐣���3\J K�"Od,�0�N�"�����OӶ%8�r"O�����756`+��6=Pq"O�q)��؝U�Ѐ۔O�3�b��$"O`ui���6���U���-�<e�t"O5jң۪f��c���8hֱ"Oh��&K�"��)�UN4���3"O���mM�
+@PA`�<i@�s"O���ȓOH���΁$>H���"O¬s�Z2Xy�͋��Q�� ��$"O\�r�
M�4��
Y{�ʀ1�"Ox���EȤgܖd3@ǈx����"O
�ha��Y���
[h��W"O8��'�A���X���w>^,SB"O~�)��˸F}>Lð@E�E8��Y3"O���B��^�x1�oV/hR�e��"O��B�(��j��Pbf�Z�v"O�i���:"u��*��_11�$4��"O���G�-d�p��d'̄�!P"O��ۃ��r`y�4MӰIf�ap"O�ҁJ'e�J�[�L82
ҷ�'`�`P.ZgB�@�Y8%�X`˷M��h�'1�����O���O���O>���O�5t���l�t�S�����P�F�� 9 &��䥀=F��;ËE<]�����y0Q���&V�D�:"L�%Jtp�ϋih JU��)��x���=�v�	�AK;m��Mc��@{�ɻm����J�[c-@�.=��ݜe�%������M�����D�%B����|⡁�	EX���-�N2���@G~�'cay��̣F�xT˗���b��h�q_�"���Żs��]n���`��4��`�q������O��w�D�ӂ��.]�Q��Ċ���K�)Q�����O���N�(=c�.O	<*Q�����#�t��ѳf�()����[�dZ$I�?��LQ剧!������5>��sw/�?���:鞈:���`�D�4:5x$�M����&��&��i�O�nZ��M�����ɍ,D��y[�A/K�t�X�E��MZ�hB�4��'�"}��=TĞ)#�H8�a�R-��A���T����ڴ�M���߇6��h8�e�Z�uX���O?�7�9$���'*T>�(Q��ğL�IƦ�ҩ�=D���q�ޜr�^C�� !�eJǪ�&B�� n��#��S!o�=~�4��)�R�ih��*tM�ՐT0�J�?�F�p��a������g����ᗸ#��F�.R��:��D7Z���5�#**Z����"a)ԑ�$h��MSUEKݟY�4�J�ğtF�ܴm�zсf�_6.�J�#���Y��?�)O����\�M3A��9�Ec�:8 q���dl��lu�l�T��cH �iW-_�N�����)-�.��O���O���D�O����OT٭��?�޴}��!Ї�� �� r���+\<Ր�OG�D��Hͳ�ʸ��%]�}����	�(��jJ>� R�j�@	>��!�%�T�^�����"(u	\59�HV7T�2�ە�U�"N�
q�R�uO2V����>��9#�o�Z�j���-�(@->�'���
��?�R�xR�'��T�ܻS��J*9��P�h���Ӧ废|�I͟h'��}"q��,r@����C�R�|�1�l.�7M��)'����?�'H�$9�� �N��Ԓ��@h��aG�͝l�P��'<�'��EߟN��'PR�Z,*1�7MF��8Ek`ʞ��@��,gnh�ui]�4jD��,�1�m���d�"��yS<%�@`��Zn$��`Fy8<h3a	�a:xȅJ[����c`p�O�����'8t@���ς2�X�V�_��0�p���l�6-�O���?	���?y��d恩qJ�{�#kb�ز�e�3�y��G'Zl\Iƃ�afȬ��ɞ��~�U85�6��<!�	Y����Iȟ��O�� 9���b����A��#;h��/��Y����O�����@���i�H�Y���E�A�#O�rԯ�(H|D�B@תhjr�bB�"g�+a�I%)I�ԃ��ۢR�rQ"! �;rDI�'�|y��*_���?X��@�$UX(��*;�$F�$l2D{�Z�l���O���O Q��!�/zT�K�¦��?q���O��I����u0��#ƃ$�y���'�46M���mZ�x���(���Gxz�rƊT��<�N>�}2��v <  �   d   Ĵ���	��Z�tI�/ʜ�cd�<��k٥���qe�H�4M��\70<����z@�v*ɾE P4%�M�R]M�Q� �6��Ϧy۴8��$ �Ibybl� \�!����V��XS%�,8@ɲ0�PK9�=a�#?t�7M�dn8,��W*¹
�c�.2���&�ʠ�"��RG�I�Us �j3͔;���<2Jڽ��%W� 9�P&�92���Ej�6*;�v�tTx��/0�H5�V%�?)�'�������%g� $�r���9F�(�fbSA}��{��c˧~f���'�(� >0�kÁ��<�cH�y�p�I֍�I���C�+UC?�� )�Ƹ��Dy�+�	�0����Xg7�	�q:\	j��W�8����J�6��#�ߢi�~�@���δ�O�y��?l�ڠ�ጔ\^8E˳��X�'���Dx��A}���	���ɲ G=r�`��+����ɱz��;��$�/��*�:Fu12�V�+��j�K�'�@�Exbb�2G@�`�+cx���13�� �}��LT�'�pd�'�ر�BD�]Y��H�!� Qhh�k(O�d������'/�� 7�,h5R���#@�u�N<�-�t�'��Fx��˟L@c�ýV���6���@ܙ��/>�I���쉂�xr���%�6�J@�=7"�-�~B��}�'�i%����'��U[���CK8eS�էRub����v�I4���	��iݩ��rD����y+pm���1-Ƹ��%S���'�\%FxҎST���n��N�(Sb�!H�AB�P8�Iv=�x�1�I>H�fak���0����)26ۘB�I?t� �  �a�U�<��	v��p���wv�T�B�U�<� ��RǭJ1I�13"%S�D�v�D"O�Y²΅�"�`��G���V���"OP�4d�+YȞx[�S@ڴ�@"O��"��U�@n��:�g��-Z��q"O��A.͒Z�b�X�ɠPR�|*g"OL�i��	�pcDM�H��¶"O�l��_��y{B�R-V=:���"OT%����d��`��@�Rȴ1�6"OD�j��>x�
mN�a��lZV"O�Y��?Nq@)����G�p�1"O��q�E	����m@�.�B(Z�J�ON�{`���M�O?�ɥ\�긻��מ6͈y�e�˶	 ]¥ã=:騀��k���#&�8h�6�>I���H��/��LL&�+��V�nJ1�g�i8����A�Rm��0f�n��T   �
  w    �!  �(  �1  �9  @  SF  qM  �U  �]  <d  ~j  �p  w  H}  ��  ǋ  Ď   `� u�	����Zv)C�'ll\�0"Ez+�'H�Dl�N��:O�1"�'"d7�R�)R�ĞH{b����L)<H�yi[i?zhЦ�� �7C~ݵo�?�ѧ�?1Hw

�mR{VA� t3hň4��IЌ�'�Z�*������.l�C&g����?��I+e�.}2���7X!���d&lŢB l"đ+��o��z�-�U�n�91�i:�M���'t�'d�'��$��	�$2$D�	`Ν���'�r���>/vMkR�T��;l����ȟ��ɰZG�8���+�
$�C� �~p��	۟��	⟸�I%���	�b3���`���CP�cf��*-�Y���7z����I�<	��*s�Ƥ��RE��{ƧBs}r�j?1ҡY56$�'d7p�ISK<"��|��oL� �P���ПT��ßp���$���ĔO����d����Z�"JPju�'�b$e�R8o�
�M��V��	�4��1`�i�DIyr�'�T�P5�E9]���X�^J�H�B	!ғJ	\��Ղ<�'ɊxC�jEt�x�؃-��@Z�|����t�T�K��W(]� 	ܴ�fC}���)�T��0�3CD|�ˆ"���H��-ݻzEF�g���e��#~��%�r�Ȥ?�L=��	E�P���zu[(�M[�ig�6�7.�<Hzq�ײ
��Bb�~aC�k��S�T���l�n��7-B�U(�4?�pX��J 72<�Kզ�.����fg�Q�Xy1���!�1���;�܁p��������i�7�Y����Q�ʥ*{n\�ٗ?�4�R�i���Q��ڊS����� �G�V�k��<Y�����X?�.z!K����������'j��Aҁ�`��t8�}t�uj��'��O8���O���4�Ŧ��O���2�A�{�� ���4)q�$*�����O���d>1	Vn�|C��0�IƇ���o�1@���Pb%_�~�� �!F2��M��I��
I�DE��5E��
���z��ե	N^lca(B�ByN,�'@#O&EpR�'ª�<5&�,�0!���'.m� *Nڟ���֟,�?�|
�'/P�-Y� ݌���+�7�a��#6��I��q �cq+�>p�E[��/:�7m�<��+�(t^�dNa[bY>a�����?�"h��Qo����.7V�حj���柼�	�F�����jy��'6�3}�(D�l�&���.��m�,�hѭ����/N�֑c�$%+P\�!q�5�'>ռy	f�T|(u�!�W�ƙ�'�V8���r?�f�1�S�?��'{NPh
5���K��,ɱ�
�R���I�� ��X~��
eN���%��f	� U��hO2��Fl}�Q�`�'��å�I&6��\`�J�9{�Ta�I�#�b9�?1�g�'W��X��U"nF��`!R�glp���'`h�u&�Lܮ�P��*X�`TR�'���I���?un�lA��Z�6��
�'��;�!Q�@��� G�~�%�	�'�D!���`�j�ёD��Li��x	�'+��z�bY�ep��`!�6|*�$�)Oh<j�'�"�b2�Q�0&N<9��!m%L��	�'Z�����<�x��i
�4>�I	�';2	K�(��jb�)�EK/7�"�K�'00\r�֜h���w�D�(���Z�'����f�|��l!`d����APϓo(��h�i<�w��h�o�9G��K�5��ˀ�'�2�����'���]"pĞ�1�i'V�����ߵJBπ�O�V���CO�!�&�xE�0O �C��<��/
2Bꈝ�d �?> ��ơ�A4���Kax"��7�?���p���'8��KǕ<<8�q$#F�4X� �S���ID�S�O���s�.B�t>|Q�Q9Mz��yBY��D��u��Qj�c�EԜbA,8X�2��WjD䦑&� �T77����?�'f�HP0�Z?�i;�L�
�.؂�'��<J���{�XA)��l����'lp��P�cJ��!Ə��d�:9��'����2�J�kz@�cV!�=M�B���'�X`�
�O_b[�^�y��T�
�'m�x9!J��~�<q��\�{a��AQ�i!�'�,� ��O7��'�\�� ��H?�( 1F�/!�>e;4���P�VH�ڴ�����9�ޙ��R>1�#D./��I2$�D�TŠ�	ǯ	�>�D��Ҽp���JE
��t�4ۈ�DH�G�����*L5����<����?\�h��4��	�w��$5��O����O��� 8oT4�:�P�/]���g&(<O���?�dA�rypV��"Ж����fy.z��mZy�i>U�Swy���
3vT�U�;vm�OC�q}��`��8O�b�'���'~�]��p���|��揆��dI֯�a�
�K,4|zmO����u[㔡˗Ė��fa@/
W�d��5�O�t��� �����<��ec�, C��1�O�9��,Ҽu����#��*��؀"O$���O E!+��F�	(���|REy�R�O�ⷆ���'�\��������K\:/� ����$�O.���O81�'��|��qR��ΐ&��)� �[��\�"H&tPT��("�z�B��'�R�pQ�G�iEօ�%�	�y⧛�x	���!�é</J�P4���0<Y�L՟tsٴ�?���z4���`�?hNȪ�̀;������?9���?����'��'t��sN��D.�lW��T�+�OD��	�wZ��KW.	6 ����ş�0Q����<���_{��f�'��P>8a)�џ�F�l�2�8e	 ��E�"'Yȟ��	p����	D�S�L��C���H��Ds�H-8<eh��#?�(�[����l��W�֌�`��7�dP�0���9#�Ob�$�"|���r�@� b�����R4-h�<�!� .7ͬh"���C7$���	�f�'G"�}j�L6^��)�K�	B�\DP�Ĝ
�M����?�Pv�U��Ş�?i��?���y��!b��)�uN�%�2DI�-Z&��'���h�nz�y%�L��� �����	@�f�G�L���S�YPa�RX�g�2�����d�,��d��xr��AK>٦dAşP�|�<�p!'aX�G/�;F5�\kaA�R�<G"C�=����g��4g[�lP�F͟��ɲ�HO�i:�$��r���**媢l�}�N��S��2�X�d�O����O`��;�?1���T�ýoG�PPՌV+m��sI�Wׂl˰��b�(��u�R���!bDգ<���V-^�p�+��:qr���JS�|�:a3�'�,�ڤ'����x����[�\�Z�E��?y��i��7m6�ɾ��O��*�/P�wR�u�5��م�y���Gy>�`B�I�/-l�5���P���qy���2��7m�O��d�?��!0Qk�"6�U��n_������O��g��O��p>=I���O�c��X��~Ȋ�1.�T�ށh�N-O�H"�	!$n�lXǯK�o�8T����<�j����;~[B�(��$�u�8;*�ʔ��U!�D�5)��4@ȚD-ZxCg�� e���O�$���=I����BQ�@��(��|b�Wt��6��O���|2����?�#����SU��n��z��]	�?��\�J9������Ot�g�Č���а��C+�)1Uo�)��	;����ңp=|a�F�O5U���W�x�z����֙'�t�O��B�'H6M�q��ڞO8ĵ�2." ���ᑪ��z���ϓ�?�����O�v�H��r@vm���O� ^ў�I�����<9�OǦ! ТKļ���֭��`Q�i�"�'��J9=�l� ��'R�'�r>��8�u��I�*TBtaS�t�c�逓~r���Nn�* �D�f��'A�ON�瘂_���
��M�,/f�#�	�2:9L��VN@�0i���⢛&�1�\x`a��d�����HV��d� *i�����O�IoZ<P5-͟��|�'�Ҁ˜:_p�Ё!Hl�� 5#T�I�ў�F{�'^�0�`�6�<찐oW�O�"��'�B#�>Y.O��'�?�-O�P� �4Ax�Z��_<1��§
Vv��d�O��d�O
�dº����?�����ܸ�� ���R��YP+�l*�BE
$@�2�]��@aq��'e�غ�Ŗ�=P��&j݅'�~�h�͔�;0���a۔H�>�9�h	t��9���D�5z��sv�C0V"�8��l�ܰYS�'�"�a�F�$�<����'���e��3/H��e��o�R�h��',ў���˟0�<a�l�
1�ȁ�`�,x��l���HAy�'M6M�O��u�h�`�i�B0O�	5�M	O�l�q`�7;�I���'���Ɵ@�I�����>([��uiB<p�"yΓ>�`���M�O��f-j��I�w�@��`Q>W���)��{�p�I)2��Icp
��l�N%QJ�54D��Z�S52 iӦ��O��k�X�P;2H�Ye����-�Oh�$�Ox���O~��Jc�$���)
�g�t{� C�J_"G����Oۻ����$��a�ʶ:�z��D�'x��!bJ\jٴ�?a����_7+����ܸh[ "͍|��إ�ĉR�����O���Tg�Mۺ�'��W>��O���a� ~��ҤP6-��hT�� �"���_z��B.I7Y]��"��8##q��L�bM��Q��k%�W�h*4Rԑ�0�׊�O�an��M������|!0�7���ҍ�e8�1rF�|�'"�?%B6IWMc�`��H.�h��:��"��`Ӫ�OH��7h���FU"b�W�yb廴@�O�����;���?�<EE[bʨ�{�ĝ'/�� I�^�<q�cŠ�ÅE�V;ҩ(�]�<�/�\���Q��`�a&EX�<)��
,����d�n�@\��GQ�<���G�tpJ�AP7v�%+��L�<Q���<���j�r��dJ~y2��p>1d�0pVBEP�h�5G�lH2�.�O�<� ��H��ϕ*5�\�J0-ځ��"Od�K�@��k �����\�E$����"O�)��$^�M7F!Q��Z�E!"OM�v �6\jH��A�`zN�F�'����'1�]�b	^4gY�ĸ��@|*���'���H�-�`e�dgI>v�Hc�'RZ�	��!�d|�t��A�^�I�'�tmQ��)[���2�]��'�`3��!x��Q�@J�:7j�{�'�d�rpn����y �Q�G���8����&NQ?�rwuH�mq@%C�O+�\C�8D��X��:~l�q ca$.cIQ7	4D�4���P�C�nA���O����餉4D���ra>�I@A.�7����3D��%Z%@	f���.m�^�;Ǫ<D������/@�2$W�<F�M��.�Or���)�'cFy��j֣+�8�UP^�f���'��I(o�!�4�T�V�QY2��	�'��1f��#C&��
�&ً{�Nг	�'��h�j.M�*Tصg�.m����'��.>�HC�HãVd�)��'� �S1a�4�!�Ĕ<E上(O.����'C����3'��1��@ 0��+	�'����՟j��i!�ǫra�ih	�'�ne�0��K�TQj3ŕ*q��Ac�'KA�0鋼���T�h� ��
�'��p���?t�&mR�%B�R2��;�-�H ��*m�L��^5��@�	�mF���8��C��J"����45"Be�ȓiN �Cɞ�C�,�AJ^� �Շ�x���I_�`�`
�ό�(8���ȓ]�5�p�U�]N���oT22�4��ȓC ��/U�*$�%��)vj�E{"�����x%�C� ����|5��"O�آ��ю+�EQ6�ěr���0"O	���`�&h���OB�p��"ON�TNG�_l��(��	e,�A"O���UNU�剢��,4�"O0��'�J8��
��k�$AYf�'��ɏ���&3�Y1G)נa
B��'P$��Ї�����.��tkԍ2E��(��E�ȓpL�$ c#�7����,�3Rb��sNyIA�_�B�dY���) �=��L���u�H��U�%Q�܆�;7�ec1#ˏ �`�@�	� vv��'�|�y
��j�ZG�� ����ӣ������ȓ�$�B�XXB�p��D�~
�x�ȓV�n3�ӎ?��&��x.�Ň�}˔QpF&��k��u��'A�]�Նȓ�� �E';Y�Ȳ��~z|8��I����	�-d�)�m�;��%:v�vB��?Z��)daYA��I8a�*I�dB��$�����^�Eg֡pT�^.^8B�I��ґ����1b�Zx��]�gԸC䉤	�rU �dO"0|�	�	��h$�C�ɻJj�K�e��N���X�D[�_�j�=QA�{�O&�E�1��jkr���	�1g�j�3�'��`'���2M�l����m"����'�b��*ؐ�>�aA�e1�U;�'5��V�y���ȥDZB�y��'�I u*QU����5U0 1r�'�>�R+lmHǪH�Mk�:����MFx��IY@��胄���20�ϫp��B�I2����J�;O_r)��� ~�B�)� � �Vb�9,$&
Z|��"OM��ͻ,i���djGk#�$9�"O���¥�;X��j�B(���"O8�
��C-Jh��`��kZ�H�Vj!�O��;�	)eF0� �
u�V��"O��2��L�V*&���^&3�lK�"O�03����U2��4�0�"Ox����WW�~	���΄(�Ry�R"O�Y��)¡L����"����2�U�'[�� �'��iҢ!��S���M!NO��y
�'<��Riְ)�K����E!]
�'p�`eǃ��H���tL� 	�'�HI��+9�P�čQ�br*���'��M����&%����a�4���'�������D_��H��O(�F�2��$ˉ�Q?}p,K�N$� �B�3biN�}!��S	}��P`Tl�$��RI�:{!�&\��UrD���8��rgGQ�%a!�]�H=�� �'ť�X`�`qN!�$V�\�{�b�3U�!C�dId?!򄍯W|<I�O_2rN��q��/	/,�O?=`��ɞ,L���&����@'͟w�<AR�ɿ���Q=I {�`�t�<QmH�7A�݋I�|�Nl��Ǌo�<�'� �1�j Sm�;|V�J�&c�<i&�S8�"�5z�(��B
]�<��a�]���A�neZ�����by2�آ�p>��yr��+7Κ)SG���u��T�<	�K0=_����'j/lI�u&�H�<Ag�	�-�2�LX�n�B�JD�<�A��8B����M�와��X�<�sgR����P�_�b
.��@hLWx�\�������1KJ�<�0�D%(��yC�(D�P!$h� %LU���ǻZ=�0!�j:D��3�@�j�h���C=BYp���&D�d���P/mN9*f*B�^R�8��#D��@w�r��e�\�^��7�D��y�Ѕ6�Ȥ�����T[7,��hO��˃��)*�= � W+pW�,˄����B�I6=��uMA���	3��>Di�B�Ɂ]����gꍛa#�eAP-�>�bB�;)��H�l�&Z<B�Z6l ZB��:p�2$񑨎�z�
3'@� ��C�ɁƪI0E@)J��tHZ�x��D/{��"~��Ń01Z��E���D��d[F�;�y�FDa��p�0�9��Xg�\-�yB�����!�.*�p�EID�y�Ȓ�R�N�s4���&���e���y�Ǟ.{�n��dG��x$;���y�R�F�p�������E|L)�.O"	��'�	c��8Gy谁��NDxU��'����Ջ}�4a��Ωd�	�')��[�/�>]�ژ9�䐴X��L��'�!�=s�0��ԉ��S�ܭ 	�'wV����!��
��XEӎT��:,p���N#�`�%�:�n�Yg	%�6�����ɨ� ,���9&HGh$h���Q���� L}=��So�?ɜA���>A)p��検�%�À��P��/N��#F9}�p<i3��71H��}�����_0.�FC�uIr�D{"�����ɒ7�Ѽ+��w��-N�(9*�"O�-�f	A?bQ��[���+�"O�`:��\�S6tk7�O�g�Y�"O� 0JvD��N�n�B��Y�:C^�!�"O�8c���u�~1���WR���w"O���E�/�hip�*���>Y�R�'������St�t���8)����|a���X��P)�+��v_^Րulݪe�Ն�^�~l��b�9<�m@�KD*;�e��Xo*ua ����L� l��e/ ��#��>X,���_^�}��n~�#��e���X��Y%v�j�'{h 0	�5N*T��@�`S&��`E#��5��d�4���Lʏj
�ҀkO�=iΔ��d��9v(1�M�2搕�ȓo*�����^
h�2=��ǩpv-�ȓ9h��Yр:w��iBB���B��� qx����c��U��G�0���`$D6NC�IV�tU Aʶ,�L��4xg�C��-���:ʒ�@�Ι@d�����C�*aJ�`��O� ��e'I�3|C�I�u;� ��nN�N��ՙc���{(TC�ɰbI�T2BH�:䈭J�z�B�=��C�m�O��(�6E1'�!��M�{d�z�'���ð�ۧO���e�p�L���'%�\�e�*%� �´Ȓ0tH�س�'
L=x��9c���SKY?nn�D��'�d�ð�;X���S3��`t�e9�'��ه�\b�����8z!���6�Fx��i_r���@��톀eÀ5g%<C䉍 ��A*���B�,� �܄w�C�	�bx�P� �w1j�[�"��C�	�P}�5����,+8��-�,C�I6;�Ĩ�C�S�k 4kt���:�*C�I�O�ę`��:_p<L�Q�UB\����v�dWT}Bm\$Hʈ��4vÈ������F+\�rܛ��\�rJ���ђ�?� ��=�?����?m��<�T]c��@&(�H�˜����)sB̏S(���d&H1e�v��'�NDEy�AL	gG|� ̠_��`"�aC�$+���V�-D%������ [�f�QadK��iGy����?a��i�b��\Mh�@?_b����
�6D��R�X��ɱP2�cp��x���Q������@{y򈃻�
���dO72��e1���6��'���*a�����E'!2���s��8Nd�ҠNI�!��\k�L�W+�J;�$�r�3�!�dU?r��emï4&�iGK� ]�!��M\��EĜi%0�Y�)�|�!�	P��ʒ�6 7��+�g��!�$ʠb�T�ۃ����l��]v�\�щ�"�g?�A� H��zAJ]�k��4�1e�h�<�4j�o�|�Cl�	 $Q��|�<i��@3�f,ZVG��k�pp��IQ|�<)�^�T���ÊƵwE�'�w�<	ҧ��o�4q�J�ri�-�x�<���٢q
P�$��H'�����%�O
�`���@������~&�qD"O)(�bΓM��dj0�/_���"O����%Fa\��tË�`6��S�"O� �!�%��%��*-�L+�"O����ʏ9H$^��U��4v�*��'ʤ��L��c��@>=*�0_� k3�0D�� ��$��H%�Ĉ �T�"`!D�@bV��
�ر�v�����B%!D�(��ȺI`Tۥl\�rVq�(#D� ��b�/A���
�h\�,�Z�;g@"D��[1�	; %�3�T'0�@�?�əl�"<��0��� Tx!YRk�,��"O����Y��]Jq�E61���z�"O,��g���`9!J�f��G~���"O� 5��ɭyҴ�B�EW�J��p"O���ǝ=?�z`�PoS+iH�w"OeӠf�s �QA��"3���b�I���O΢}��0�0Z�CA��]S��ۨM�@��ȓ_��&>KP�� �3tZ�ȓv�1��	C2:8NEy�^�`h�T��o\%ar�W "U�7F�(pHx��ȓAT8<RA�Аv<F�ڰEX�E�͇�jS��Qȉs�$�W�֜�\����azb����䥒&
_4��Yʧ��n;!�D�eB
����J�/xd]p�Z�l!!��@���A 7H�H�ݵM�!���<�&�� IٛZ�d��`��x�!��I~���tiɻA醱1�
˱E�џ<�Wc�'�M��?	�O&���"���^G��L�����?!�ɀ��?!���?9���?�y�O5"��
��{�樱@id�E"��D�?)yV)�D��q���k�|�
F)� m�D� #�(m#��Om�'^���y��Z�a�χ��3� ÷ ����"O:dq`LD�n������X�,����|��i>	I/O��3T'�:l'D3��U(N����X���	���&�������'�z�$'t�ҕ�G���!�"�y��$P\�O��hH%��2z�B��%GË0Ø�?Q&�L�8��?m2�j@�=z����lh�Rp+�h9?!��O@t#�>��y�,ө+֐C�Y1&(�2�Öo�2M Q��D�N�tAC�3}��9��d�q"�*�& q:��� ōS�>ɀ�O��}Γ5��!B�Z�C�Z�{���.g'�!�!�`��M�Ĉ�j����S�,��D�U��E+z!r ٙRX�$��XZ�0/��D�Te�<~$�d1��L1 ��њ���/%L2����	��I26�~�'�>6m�:(B�bCZ<<���I񯞹#D�	l��'��#��̌z`��*%N&�ЉC�Ê
)#�D����S��'�lK�Ov�����GÀ�Q.R1?����BaY�ʓI������?I`5ҧl�����%����S��8A���	:����:��$"�9O�5z%�OX�����]����kYh���Z��'�l��I(T3����6A�]"+��M��B�	G|�D�%X.$N�{��Uwp6M�O��D�<����?�*O�����۱D�h���O@�6�s0.�˦y�	[yB�'�\�'�?A+���ر��4��.�Vx6
�9�V�lqy��'5�	u��Ly2�؁v�QĄ�_$�1a#��l.>B�	6X���0�#u<���Oϝ3B�	���Ň�j�g��PB�ɯ}�d��̇v%䰣� �H��B�I�:�2<�2��C�(ZF�E6U�C�Ipfp� ��01N�8$�[��B�2u����%�6�Ƹ�τ�k�C�	�eL!so�X�ޕ��ʗ��!�$"U3 a)����̪��%�!�DV�_H�T�5�5����ظb&#<��K�?d���D�$��L�REb�S!RO�y�A$��yR�ш��xq	��;"t�� �
���'*H�B�E+`"#eܧs���H�'�! H�=�\����(P�d �������bOI�d�V����Hzk��؂-���|d���2&8f��t���'�Z9[�ID�P� �K�^ G��!z�"G#}�d�!��]�i����->ZD �Z���J�B
u�LQ;d�9K����ŋ��X�B�/24S��
�U�q2@A�?!�-Kv�zv��7qɧ��~:HB0�\a��F�M�����@�	bR� )	6�Bř�D��[p��D
b��0Ps�Oք�����S�Y�F�`O<�7&����4-��6�'���Q07�& �j���6-Fu����O���dܙje2(�CQ(n�,eH�O�\�xR1�u-��j�_-	�����:c>89�#K�6e��'<�B?u��]i��'r��'~BK��"�8��M�=�L��]0�䠃�ޒ#�`ؓ)!S K���1����'�rY(�"�
Cb�����|@8��ڜ{) 9W����P7囌۾�Y�DBV�D�^K:��0�,TS��&0����F�R$��Ѻi��6-�O.|�Q��Oq���Ц���S��IGQe�"a"����x2�F�T(>M �.�
4#6`X�O͵���HOBʧ���HN�$e(���^̔{4N՘�����Ț!�<�	����H;[wO��'$P8���c+���=@��M<�4@��ܔ���a2�ט`R��$M�? h���юq���vAY,��U�
��i!6��PcRU���gr�AD|b!Ё�^�+5��![*���%`%3��H���?���i��V����S�+�.`0��w6��ǧ<�x���hO����O�Od؁e�<*Jtic�5*/��L�]y��')V7-�O�A[��	��i$��i���%�S*�-��L��!K6�j�O���$Μ���OD�dI�gD���<ݴR[^-(� j�2���.�t�剏7�ֵ�R%ˠ"2�yƬ�8��'�!֬,��.]
�P�˓@�a�I �M�b�O� z��$�X�b�ٮ[����>�Ѱ=qBˇ�NU��yѮ��o�sЭ�'���'��Ia��� ��n���B �EU�����KsVU��'�剛'^��QU՟��d�O��i� �:7�\�gM\H��R�7dRm�c�ͻC6���̟��q`���
g�U9W!�p9�S��^?���D]�5Ⱥ�1��Ξ<�rq�c%��ͅU�E��wZ�S�5�'-�B� w`	�,\1�k�2Cj�$�D�b��O���7�'�M#a�˽R���If	�S�H�R�T	T!�H�}X9�&��1�4��ܚw�x'$�p�vx��\�a�x
D�\�W�	��Hg�8���O���]�8��X���O����O���wMhM�t�{��4����؃�F[-XEJ�䪓�{'�`@�B&/Mjc>i�O зj-#:�y����*&"��Y�pZ�*�+k�Co��e$I���T )?I�h�03��x���6K��|'��D�◟����O�"�|��Yit�1����Ujd�ȓz5��'*�����Ǎw���O�Dz�O��_��cu�%�
�U	ޔK!p�ɥfL<X�Z�X���?����?��!����O���>)rr�{>�-끭GP[z���ϵ�����W�����6�'��@���i>�Ra۷IH��`�6X�i��W<#V݆�ɗe���Ғ��U�e��g��6^��2��O��m��M{��;=R�z�G�`���-�	[��C��
� ���6\�\0!�/4���˯O�b����5�pi��:ڲ���8j>��]�lG{��	�\�l���O�Z��P��V��ذ>ץ�!0:�B�4K{�)�V́u�<����P��Z�mޖLI�Ty��o�<�B腟$���f
&ފ���#@�<�/V%F����C��''SbtSm|�<a�P-�@��3Jz��L�r��L�<�QC��	|xݫ�HR�h�>�
pKK�<A2��=n扒'-��Pwz�����`�<ɂ���(X�/Yy&��UhC_�<9�ڦ^2����E�&llH�H�Y�<ْ�ҥ!�m�x��}�OR�<a��B�o�|,a���e���tFX�<QW��$${���%���>9�`(CdW�<��I�#CEf��3�Ґ[t9P4�RP�<t��������j�j�;"g�H�<�G�ʔ���V]��ђ�k�B�<)Abݣ/w81B�.��6�P<�CYY�<��^Dy1�B�Gd`�����S�<�gMħ=�ʄ�T���u������F�<�q(�&9�A	�?^��%�SNB�<q�ّ]Ʈ�ŇշEs4�I�g�<�����'�C4?�<y�'�b�<� ���U�T2v%�.	N��d�U�<�V��O<���D�q�.����R�<�7DR�YX���HV!(�~����XM�<��`�
lB��sŃ�G�|��hJ�<)� _icF�zg�oO��h''�G�<Qd����0���u㎕q@ "D��7�B(i}�XH��	M�L�a�-D��:�Ӿ\/BCw�2�<��D&.D�t�3I�\%%G2�.��p�'D�ls���oV���Ŏ�(� �D1D�PI���M~�1�rɽ2���cS�0D��(�E�A;�������P�I.D��[�J���lx����RF�@ rO,D�����0�d@(�(�5M��4p�A/D�� ��+R��,�1�U.Mh)D"O>(7bA�5\��@d�+"\��h&"O质I�;�`��1
�Vۑ"O�e�%���p!r�֣e~(U#T"O�@ۀ��%a�B��g�/dD1�"O�i�c� Si,ŁG振!dx��"O�u#���y��1��/�-y��,�"OLLI�I�f�H�7��oq0x�"O�h��>5t�2$/��^�B�"O���M�$��� Q  "X>��f"O
t��c�W&�[�/�< ��� "O�y+K,-����0�1|#f r�"O&���L3S�s�� <
h��E"O�T���0�$�#���4t��8�Q"O�
��=>���ҏ�����3�"OFt#�� {���n����"Ot�P���16 1Ь �Tp�])V"O�2$�;m���P�
�`�q��"O�z"*5:Iʍs���
9_�!0�"O�:t��B�NH�2�
�JB�1�v"O�Y��̝"�jY�8Y)a"O�s�YS��,8e�c�Z�"O -�S퍥��p�F��,H�0��"O(����K���pj�hh��0"O����l0vw�u3 ˅�8��3�"O$�1w*F��|����r�X���"O�L�WVE�$	5��X�"O=���^�>�4�A��g�Z��"O����E�D]B���޲c�(�"O�h��R%K����߽_<�d�`"O�p��o�`$�b�N�s8�C"Ol04F߽�Q3�C��Z �4[a"O��W=�Z���lј	-��#d"ORY��m](v�XI[e�] ;%���"O�I e� p�N�s�i7D�I�"O.9����� h�����w"Od����(� ��Fጢ*�<QȠ"Oμ�h�8`�jw�������"O����K;UV��Y�����	�"OL�rfo��3đ[�Nov��"OrqS��~DF	Z��dT���"O���꜍#�:HW"N:p2"�"O��yA�K�r��+� �^��6"O��v�Z&TKH� ҆'h�tY�"O0�H��ܔ\��<3�jؼ
�蝙�"ONl(��ބA��{7ꄈV�xMW"O�P������䑖HH�90s"Ou���I�8�.Z4`���D���"Od�sE?��⴯��z]<{*O�}h�K�w|X\gL�&�Vy
�'��8��
X�}Ɗ�1S�	G�	`
�'�RH2�o�%8u���>��8 �'n lx��w�j�HޭM����'"8X���ϹY�ڹ`���4UD���'3؈���B�h�l�+!�U��]��'��p��\,+ę�_�;�RM8�'�A7/�W����셤.2~���'��@�I�cO~%Jʀ�/?�P��'�^�SeI<����4a��Y_�̀�'	^)I� [-��TDE�
QQ4!��'_]�� �(@���9��&3�X�I�'���Hp�P����p�S���t�
�'!��I�m2JH!���$
:���'d������u�^��HڜLȖ\���� �����BE��j���>e�J��"O�x��� ����7i��H�B"O� 撲#w   ζBuf���"O���Бx���Z�� fj���"O���aH��M"��{7fKVb�X�"Of���O1��䥄�nR&\�"O�mz���EUx�!P놗?klLS"Oxhh�ʒ4G�� �a
�]u�Y	�"O�
W,�l���HO�mTr"#"Ovɉ��p�"l�S�#sRCw"O�镦���t�Ei�7 �����'O���GO��f¸[d�½Rw�}�
�'���G*��?M� �f�!xDy�'��xsF�"A(8J�C�z�h�	�'\P#�ǝ
��%#�*~�:|�
�'a}[ F�#jtB@�ī�uȄ�0	�'�xAC�*�Oz��A1�ɐ��P��'jayg�+t(��� ��Fav��	�'�����j�����87<�T	�'7�����;vi�I����$(m Չ�'3��@4���͙v �
"�ri�"O��T�V�\J�d�G�}�ku��u�<	�!V��Ν�q5^OyK�r�<��̆MM,S ňiZ���$	q�<�4Ȅrf�����Z."��J7Ml�<!�;a2�M��' ��`\l�<�4jٯAF|�&.��w��]WMOj�<1e-�:~�����fL�S��A�<�e�
��=�͇*U"�p�`�a�<qs��(��<s��\�%"K�U�B�	�e�T)zÄ��R��q�w��|vxB�I�2Na�u�
�@�<�,��EC  $D�\�c�Z�Rv�B��"�x�;��$D��J",��C|�JS��	�( ��N7D�`��BN�=��mk1iS(,�ʔ�9D��0@�I�V��Ш��,e����8D�0 G60�p�1�N:���tj8D�T��ީ@I��CU�g��$i1D�����!wQ5��=S)|���9D��С�N.q��H$�;FN�s�"D�$S!�̣5����u̞[(2�D?D����Fb6l|�"��tj�%ȗ!D����ܻ vB�G��m��}p�:D��HF��.x�l,z�)\20w��8#N7D�����d�X�(�:xm�K)D�����s�,9Ra��
Yd�!C�,D��
�`� 4�L�&���]^Jc@�+D�\�O�hM��Yẹ(�\�G(D��ɇ�*�Дr`Ǌ�|KT�3j&D��C5		ev�z1e��kQ ��d�#D�DY�����6J�6�"X���?D�D�Tc��PV��3�OQ~ZP�e?D���A�؝x�!{Q$Bj�.�91G>D�h0�H��6f���Z��s��B�<q�܏�0���@�(T� ���C{�<Ag��#�H�@$M;er��a�	u�<�c�ߌ)�����6K�>x�!��m�<ѧ���Ra�E�3�:�"�`�<�	�}3��HBG�2��T�%��a�<��*���Y�G�K�2?�`��/Iu�<�#��:`�:�)�E?A�N�X��s�<Q _6O���ã�7� U�s$�C�<��C�,T^t�0�J�VzI�� E|�<Y�9���*�;-Ȱ"F~�<� �Z2'J7]��
�`�()��D��"O�(��E�g+�Q��[�"Ȱ��%"O.���i�@؈DI��#I��R"O*�	����8�# N� {x��E"OFA�$΀"
�
\���F�m�4H�"O�dˤ�Ϗbk���ݣ[���"O�%�A$I�=�Q�Qd͂An`ۃ"O�	��l�&�Z``%%�X�C�"O4���ך-�p8!�y��1e"O���b�$TjP��F�\ �"O�aWcӵW�+W��5R�<�i�"O��sЊ��i�k�Ab	×"O<�
�#D?~�J%+'��
����"Ov����7O�D�T�R5[�t�c�"O^I7iܢ<�Th {�W�c�!��/��p���-KSZ�i�n!�$��!bfn�BP̸��ƅ�O^!�D��09��0�B�lR�@�V!򤎊\R񂳀��]���Iᮋ�(C!�%�����I;wlrZDM�'w�!�$�=�ՙ�F)bwl�JT�B;t!�$��2�������ZY|s4�:-;!�dȩ>4J���ǋ/<Vi£a�
3!�N>5=�u��լ-��@ �2$!�~`<T	1h�mY���iT"�!�.qf��f%�W�T��HV�w�!��(�!Ct+Ӊ,A��#�f�e�!�dD#��I�'��/!N =��C�g�!�Ӑl���-�2.@�FFS�].!�dSr��|	��׬@�Ȁ��d!�D܀Q��z�:w��tpC�D�C!�$�U �pkT��ӊ=ʳ�L�E!��J#v[lq�Q �Y�`(Y��ސd�z�i&8
���5 ���Xm(�		�#"J����G�g(�1��X�<�T��0&�Z�@��2D�����o�<���[}X0ҭ@~��A6h�R�<y0*�B�ڑ7@jO�iɱ�!T��$#��W�̐B�,�N,j��5�"D��Ŕ�-�<d�#!ӣ�B ��)!D����I��:�,��DR"L�zU�s, D��u(ԅ*V��s�*-��l�W:D��ՠ�<^��Q�f�!F�x�K+D��h�dB�MNP�#iƣWb0Pk�	.D�|�V
�
�:��郐Z��Egc*D��y��� Z@H��-#�d�P�g,D��+C&��F�bXk��%%.��P�+D�$���-U�f)YT�ņ+���Cf*D�$��
�E�L0�"�B�4�Z��=D�d����:m�>�qȏ.�	�ҁ!D��#��Q����c	Q*IF��ir�-D�0 g��,Y�8Q���Ӭ)hʤ�$*D��p�*#����<,��%[&+D�$8�!B�2t�Y{��%j�&\J�"*ړI�m���Z��:F�r鹖�m���G�<�Ĉ� �s,`���BC��y2J۶<������d�Dd��%��?ɡNA
�j�@tJL&hR�7N��#}ʣ��2�D�����#&��"��C��y��ۯ�`�q㥑{dtiD��)]8���Φ5��e���41�_>���Bh9D��` �B�<�R�r6�Q&��>q4�Y6UĦ�B��D˦ 0�'$j��0a���f8��I�h�"�,qC��'/�-@P9+H5�C+���!N>�G#�1�?�f�!���� �\���h���җ~Z�Ո�h	=*�jwa�O�!�(w%�s��P%&5[��CGv
�pW��*g�Uc HQ�%���sb��8�M��l�Tˁ����C���u�����SC�r<��K���xIHէX2�L�9�BW?�0]{����4�
T#c�̊k���
ۥWxHJѯH%���� ���tn�4qq8H� H�z���'S���$��0� ��c*2N���"��	�B:^�vc_;ٸ���=R�0)���.Jwv���+��Y��������M�H�� �O6X;�-�,M"�C`��*k7�q��e��s"��-Zd��D�.n�r�v�J�P��� B��y��[}s  9K�?yb<D�K+<[�d�3�s�4��%�� >����S]3�Ik>= @�[�y$2R����M��A��-��(���0?Y�@Nן��4�V�,�����
�m�t���I��,�$��W��1�H߯HؔY�0�F�l!����N��]\��@w�Q�m��	�����O�Hҵ�{���{mK<�:90��+)z�-Z��D, q�ճ ��"����hղ%��Q-+ �a��I8�и���ºx^4ih����d���	�*P�	��A�� ����II`eU� o����X�B���(5� �2A�N�n%J���ŝ��!��B�A#v,�7��]ca�n�x�K$�"G�iq�+�v>�����$˧4WX��˼{`N��l�e8vLY;o�2�j�_b�<���e|���'�F��j�� ���Z�K�8�B�c&��F* �  ���%����Z	�PQ��S��ڹ ��M7��<��C�]ڸ"�]]@.��2+Λ1;���)?6a�Ю+�b��g�y`z���'0�a��4l,Td���d&�ēM"2�*cI�8`��&=vli�".��RV����a���ًyX���7����R"O����+K�e���m��b�P͠�Lh8��[T�o���+��<z���/#�T$�Y��.\|`���cٹu�,��.oY���@F(���2z��+��аRd\��`�ʁ\��)n�"e�T���:X�Q8��O�*�`���^�-�3�\�	��(���7�'�z�I��ߴ�?���~���pT�":��]Y%Ń6~42ăc��]�)�q�Յu�h�E�'|<ܚGᗐ"	Kf㔄x�p*�O�e�AH['$��ܴr<�ܛE埀,]�	Jd眔XZzpo��°�a�Ҡ%�ܔBA�:i���#"O|�	�I�k�~��*�v�lg�g�8�u��?���b�m!������IE�Qlf��d��sq��0K���s��L� �� �O�qu�͡�1���P0@�kĩ��6���y��T�e��k�@���g(�q�2�"O>�{�j%S�O��!G�B2X����^����0"O�:��LqzMAG�M�c�y҅�|B�]�#/�Oq�.�#@�Y@���k���|����"Or�І-̠@	���7i�ƽ*1"OP�qu��Y6-JblYU���R"O���r/NT�&��#��g���pa"OH��c�l��@��kϴJ�ܽ�"Ort�	@�N�;�ޠ���@"O�$��E�b���!���3��̂"O\E���0g��	�bדM,��Z�"O��M.kܺ� �G�`uR9��"O��p+�$g��e����2��<�"O���&؋
�Xbf���2�n�1"O��a���"m�S@��)Puj4"O,���Q����'E;`i��ȥ"O�$�r(�EW(Z$hP"OB�YB؁4kF-�������g"O�Ac�o��6�*�p�� ���"O�0A���>`�4�r3��=Y@�9�"O����"� b&�Yb񪖂�T���"OTA��H�F�*�YGCD�t�����"OZT��R2G���
'��W B-z�"O��s�R�>�d�`���%���y�\�.a�ӈع&͜(x��'�y���'�:7/��_-P�횄�y�)�'j�V����߸U��a�g�ȏ�y�AT�q��s#�T�P��!d��y���)�������\��
$L˩�yb!ؑ)��ݨb
�P��5���,�y�̴^�"E�բ�Vf�R�%$�y§RT*pA��*U��{`��&�y���83;���(P�\�aK0�y��^ j��3��KO��p�Ɠ5�y2�ÅT���ӄ�
F�숓���3�yr%�D�piCF
�z�H�[�����y
� Đ�!�T�e�ŋu�*T�̸*�"O���D�}�f��R�v��0��"Oث��T��.�(��!?�1�"O� �ꍺ@W�1��.78�ܖ��y�N�-.�)BA��n�´���[?�y2��XaH!�&K����*�劎��O��G1ʧ:�n����	x �X�+Ӎ^|���J�|�  e��c�%����L� ��U�A:��S�O�̣S��z��ə�ΥF3���'���+#��*L&D"7J:?O�@��O�M�@f�4��݃Ǔ:����V���i�N� HR9;F8����2�v�.	��PEIg���d�+a�<���L�@ՔՆ��Zʨ���9_,����o܊p`�Gx�
154�SIK2>X��3���1�)���$=N)����y��M�M��(@��E�~I^��T�1K�u� ǜ"/\���՘E`6�s����%R�utH�Pq�=@��5��b5D��bk �T��ݑ�Z*�}b䖡j��I1'�=0������V�n����kՊ���J_�1��8��+ե#�h��Ĝ39?R\8f���+U��8"z��y��
 c�(Ҭ©3�2 ��'���!��6_�<xr��ӓ}�r8ш}�l��\�4m�B�38[|����Y���e7����
���ר�8E8��ȓosDt���!K� �b���*�8�2OT��^� Vk����H��9ϓs����j����$�V �1�ȓ5P�b�`�k,��� -6 �EY�ilm`u�%uŢ���uw %�M#lpHsm�%.��|�FIA$D���I�/Q((�����"F��4�K�[��ܐ�mmcrI��ǉӺ��C�-�0?)4hX?|���U@�2Ax��׋�r�$a��`����!}���GCD!	K�o:³�J�d�m
`eH0 \���-�Y�<�Ɇ.U�Pb�\)����3Al�PU-5a��ʚ�h̛����<q2E�6Ö]��ي!�DE�a�V�<Y�/�0C��@p3��)A�Ҩ��UyR1��$w���,P�n����ԨO�mX��)d5�Z�N�`��$�'j$�"�I2�lZ�ȉ���	�lT
:�LKf�Ѷ6A�Y�%'̼�p?�&*�)WY��ǅM3H�&��"* P�t��$�	���Í](�Ob����l�q��9��'v�4<��'^��Y�)�?
��� CKr�~���'q�P�Qd90���S��}� ��6i!���w
әU�8$��e�t�<���[�U�q'�V1F�Y9��]���D�"�T�v
U���3��	xa���t�B)�Tٙ��^R���I�L�	Ǎ)�$� ��8��L���(%�p��O(�.t�T[u�ʛ�lP;�/�]Q���sb[�������4�>9V����1o�������y�)�6��qe�ݲ#$&0m���y���,9F�|��)Q��	;�DN���T� ��>�!�$rᵎ�;n=�(�"U,�΀�xR�U�v��zBF.�����m��w�j�W!��y���#N=a���C>\���M��yb֟'��P����~�
q���\0�yRCi��}��ω	$6�����y��=Z��Q�`HFu(��V
(�yRG P�攸W��j��`e��y2�ϏGH����Ĭh�d�4�º�y��]�7�!a�����f��yb˯[��P��`zi��r�U�y�Ɂb��c�P�y�xh�%����y$�2tִMKpKZl1���y�NQ3�,E��&^c L���ʍ�yB��4�6A�,����s/8�yҤ��.�fH���T	0�2��R��y�I�`��T�#�� s�d�'���yB�]�R�� �K~�R�jdÓ$�y
��*�d)�0#�'ֿ�>��ȓ�����Q�Y�[`�F�$&	��:��j��I ��NX�8��S�? �@�ӭ+�ʗi�$ol1�"O"��gc>X���*��
o��{"O�<�"���E��q(*1��"O΁��NL�R�:�zBH)��a��"O5c�hۂ�,����T�d�D��2"O�4�a�:X��E+q�I�
Ԥ݋&"Of�R�f�`FV��Ff�2V϶("F"O�JBƍ1U��[V��j譋%"O�@v)мC�|��% �_V�(�"Oֈra�+JX��(D!Zg��4"Oz �d�x�����K/z�)�F"OL���O%n�� �K��ON�Ă�"O$�� �5k����-ǳXݢXJ"On� /Ξ��!S��N�`�T�r�"O�ܐ�jͥa̸��t��b��YY�"O��Hc]�Tk��
Uͬ! ���"O��X�@0�L�Z`L�&5���w"O��ա0���B1�^�y$��r�'1*�R	R)��ձs-���s
�'РT(qf:w,�T9c�J���0	�'����W���K:5;�ڴK�4(�'CJ���S%9P$���� U�0t��'X���j�*�,���K�R��'�D�a�X&/�>�A���	r���
�'Ga��3d�d0Z�f�eT$��'ULq��7me��zb`���\5��'(�آt�������%��1=F��	�'�%'�>R/�]k�̗g�$A��(΂�CF)˦:�S���(04��ȓl�8�a5�B 24ܐ#hY���ȓl(���u��U�<�N�%h����,���Z�����b� Sen���^��H��U�X���d@3�a�ȓJ�^=�%�0t��넶aB�����ec# U�]暭��K۝Q n�ȓ}a<��vl�6�(�1݁V#��ȓt4\� D|Ȁ}Rǚ�e����	"@�TŰ$mQ�\�Ry�r�h�p�����,����+�
`�!�۱�  �)*8}��ڴ�S�@�!�DR�T5d�3���c���@�
��!�D�\���I��4N���d�U�@�!�ā�U#�H�`Ԓ�n ���0�PyҠN�-��Y� �R�/�.h�-P�y2�*	�̈"k� (?�UA7����y��C'����u�ßx���N��y��G�2���nC���H�/C!�yR#:s�(�� 3NAae�D��y���6�h���i2�6�`� ��y�	-�Lј�G�N�r�]2�yc^�{���b/[M,�q �R6�y¢�=\���f���25�ͽ�yB�@-M���s)Y�f�ػD���y�(�S*��)3
���1;t��y'\6 �� P��^�-��г�� ��ybK{�$�0�o�*v�L���Q�y���"V�.P i
,i�~���炠�y"���g�6�������׊��y�J��WgfUh�C�E��%菭�y���<|�F�{Cb���Pm�Yp��'�b����R�t��@��! ]�Xa	�'�X2t,V�~�,�2� �����'a����
3��������x�'�t4���E�D�J��բT�b����'���5�#����i�
V�d!z��� nP"�`�=��8��A6���""O�H2� ;O���A��6R��hU"O�)�#�Q�/�܌S�I�'��1"O���	A��x�(,Y�{�"O܈jB�@]iJ����W�P��"O.U�Q'ė�Pȃ�eZ�=hM�"O�\��C �T)�O�X�2"O��yr�X����(G�eX��"O��ՈW�, ��E��@U��� "Ojxy�g���igB(WY�l�3"O@���(i�Tp��`H
#N����"OZ���#��#rdU�7o�	?��c"O����S�b=�<:�Ύ<1�0��"O`=�U�
,��x��H-.�1��"OL����=We����h��K�ɉ�"OT�3ԇM�'��ZS���(�,�(4"Ob5tF�N�"����],e�VLcu"O}q�č�C.x�tـu����"O�����N/v��D+�)�YC�"Oj��):%,%	���d�>@�"O,]
2 6�XaVE�z�d̐�"O�P����`��yQ���N��h�0"OIpp�S#Bҍ:��R�V��c�"O4ݨ�g��I!4�Q������3r"O�fn��M���Br��@Ie"O����ʚd�t�PgW�N�V���"O(��ч�]r�d����]2t;"Oل���[d���~�<��0"OxQ��¢aVmI�IM%h��U�t"O������e熸�'�[]�>�2�"OD�1�G�*zľ��g猇��B�"O �ؓ�W�n�*�	6F�+B
���"O8J�	3��!�E�*a)4�:"O�]X�Ʃ57���C�>��T9"O��#�lArX�AÇ%PG���"O*I��.�7�����'ځg4��"O�0Z&��6]�vh��FY�R�6�u"O�y�Dh�!X�q��_�"���[�"O(��N�jC�x�D�N����"O�	��l�xO@,R�B��޽6"O�U��HD�%�%a ��2I��S"Ot�Ókx�����*v�`��"O�ܱ3@Lb8!*�)+�6��"O`H8l
x=3�_?o�� ��"O�J`eѝ�F�a�˯q���˄"Ov�8F�M4 "x��%.S�t�p�@"OB��2�R���uC�M/c���'"OP�@��N.$5JE��e��J����"O:c'�Nw;���b
.v�e� "O��XaA� wzV���
5��+7"Ot�G�G�VŊ�,�!�1h�"O
$��gY%cn�mb��=Ji�"O��1���&�x��@�W�h8��p�"Ov��;<��'N�^!(�4"O�� F��q��pրր�ju�"O\�D�N�	��B��Ӗ7�J��"O��*��&W���rh�,X^0��"Op�*@m�TF��(��MO&���"O�)Zd�ޫ;#R� �>Yڤ�"Oޙ� �َ�,|`���BS��9"OT��H�%�$Yz�IP'b=^��"O�ԙ1C5I���I�
� d"On-�3��F���ʑ�،�yS"Oⴃ`K]!l�����M^�a��!�� M�����X^8c�,�-T��"O��xF�)S1��J�&�c�ʼRW"O�����(Y����O�8.�hB"O��rb�=L��qa���n*8�	�"Or���i
7`��k�<]**�Q"O�dqO6x|$X�
�' ��yY�"O`d ��(L�d����A�nm0�"O��Rc�G4!=��� �ػ�<��R"O
\�$O�3�X$cP��e����"O�qX6��I@�`����A��"O���AlA(I�6�P7���:�zH[�"O�x+%,�!_縙��쎌\er�"OB�{��B�B��D�n�0IZ��*�"O�Q�WBЯs� ���D�&�Pݲ�"Oj]	#�\�u�\�z��


��A��'s:sw�^�~!r�IG�>%6���'9t� 䘜V�H���O��9�'�z�X��$ �N�rV� �[����'�"-k��iij4#�D�_�d��'��щ��w|���Ej�X^�5�'�h���ВV��Q ���5g���'tR ��ҖQ#�eyE��'�laR
�'ߒd"ߜ4�.}�TOK����	�'C<Q�ϛ�
r4��#)�	�B	�'Tj��P�Xވb�	�X����';��3̝�JI���u@��Vf���'���C��C l�.m� ŋ�`�D1K�'��8b�I+o���Ǫ�Y�-h�y��'WF	J��d��c�@7N��$Z�'�J��C@�%*z]��Ȑ>��8�'\Lx��d�(nέ��Z<�\؈�'D��Q��K��\�S��,~��'�2��r�͉	�:��JM'ȸq��'kR�SqK��Z��$�
���'��r�7�����lۓ�ܕR�'Lx�8�.J|l���EZ�[�r(��'���E_ r��J��*LVx��'�^�H��}R>�����"Ot���w�V4�C�M{�t	�"ODm��H�6U��ȸ��4`�db�"ON��0/P'�^�y��]57r\d�W"On�Q��:r��Kv��9Bm����"O�`�tB�Q{V1��U�a\�u0!"O�)�t� T�,���OJ�I�"O��;$ )a�ΙǠ¹s&����"O�}��j�y�"ɳ��:*#�P#"O@q�,�p	���o�S�ڤ3!�dAV�!�CC�P"Rua�h6!�����C��Șn8E�3�j!�d�fKfq����K��DIcĕ�NV!�R=T�P����TEؘ��C�V��!��5N���A��8����J!�䃮#0��+Dᐌ,B�2gL�"v�!�d�:Z��m1�'ܸe0Rl���ȉW�!�$W����F0(0��S�D;�!�dC�H�ތy'\�Z!��i% �/z!���,}=&��2#�,g��:5BU)h!��c�v�:c�=8K�D`��/�!�D�>�Hq�&��=������tc!�d�Jl:-�?9�H��E�!�ݝm�r�9@n�
dkfE�����z�!���ܘj`J�fn��&b	�Fv!��O�⩸A��p}:��Ί�7�!�4V������#1�X�i͌�d_!�� ��*&G�Tԋg*ۦ$fƄ�w"O$lBs�%�<M)2T3!]p$�c"O�0��!7S�U���5%�p��"O�t�pѢ)˔d�E$P	P>��Ӵ"O���������R��[�k�d"R"O���.ZhB��F)B'f��I�"O�9�� �*� ��(鬹31"Oj!��*�9	���a�4m��]*U"O*��cf\.{j�����0:�����"O:�Ȗ�:=:^�:���+��""O�|Xc�W�d�#OY/_��˅"O"(�0�� +?4���ŗjo���"Ol��T�=׈l�m/R��i��"O|�եY�TN�I3a� �܌;�"O EZ��ɦ.䆤I��Z�����"O~8�A@T�Xll� |֬��"O��9��FE�:�"���^!�"OF��"�?<�e"��I��[a"O�Q�!F�����T��ֽq�!�$
#h �S��Է3B*@����!�D�'z��p�d|+�	Тc�!��/o��s�.E54|��dbW(1�!��<�P��f�Q�=I�d�Ǡ�W�!�T���ёW�Ĕ+,��Æ��<�!��+C�~5�w혭5'��Q�W+/!���XXxp�!F���#�NU!��
��x��援�� (��#MP!��ũ(�h�ŕ��4��ڒ;!�ʉ=@����+-� ]!k�wJ!�d�!1P3�C�R����׃C�!����$R#+߈�E��*�--�!��	�3��[�n��	�8���>H!�D��~�[� �Se�ܚG��@D!��E���i%O�d|lI#�G';6!��C�j��$�9Z`�����l!�DRhs`H���T-_�	����Z�!�D�L����À�"2Z}��'�!�X�)~5��$�m�C�=!�!�^�
��%�0C�`�ӫE+!�$U#$(��hI�l[z}�c��d�!��
�(<ۗ�ZP ��Cd��?�!�3iq���f�]O4$��Bǳz!��_6x� �Pt�Z�8M:�D�[a!�$�3PT�Cׇ��}@���-ܐ�!��[�v9�c�K�7�b�.�bK!�mt�fD�-?�nU����
7>!�O�=袅�+�^��d��F!�ʡ\?@�c��<W��U�E㍘X�!��@�.�ɰv��;��]��Q�<!�ەR�"�Rc��Q�ݸD��5!�Č�l���Q$K8pp�2�#�4s!�$��;s��[7�ȍc����	- !�$�� x
�!ͧIV��H��Dc!�DQ*w�
ث�߄9M�ѯ� �!�����P�Jŏ?;N�
B�׭]�!�WP�R���"D��D��-�!��,-?,�!OE�%���k�C��~�!��R��M��՝c#:,�6�G�d�!�$�+�M��-�@�~|��×J:!�1��!���K9D�N5ء��#2!��G�\�rDs�dȈ�a��G@	]!�$_�(� ���:�z�����a!���7�t �� AwB@r��S�'!�䆴!P@�#�^9,a�6K�s:!�� ��Hv�A��\)��ͻ2���d"O�����93���v��Q�0��"O$��ф�>p&�a��o眄K"O��c1��
�d� 2��C�LNm�<Y���57OB1�eBлꞌF��Q�<s�
�a�HdbH9&���v��L�<��o�I����tgҲ.}z�H�L�<�d��#Q:��f�ȱ"��<b�+Bm�<�#�Ҡ(�(���%P�c�THs�<�f�S�b���+<���*l�<�gf�3�Rd�P!�H�ZQ����g�<)�a+
���ї D����Y�<	�h[�{�.�xU�:u�N�
���~�<�tO^�#I�@�$g9&�N��Ĭ�@�<���S;tx�A�;X����G�{�<���L?VȜ��,�(h��LB�<�Fil[��RARs���I I�<�q��-$��	����U����OPn�<	Daթ���D�#&�D��qN	j�<4����e�^�dy�	O}�<���@+1�p�c��%�%0^�C�	�Z�ۥ�ś+���B��^�B�	�\��A�Яt�`+q Ǘ>iB�-�N}��N�y��@���H�/
B�-Pd��6i��M{�] �`F���C�	I�ԉY��.'|^(�%�ɰ0�C�ɝc�� ����`�@���B�,C�	�kC(d	�=>衁�;)�B�I9��v�։*>|����u��B����e��%�G�*1p�,C�C�I�RX���%��I]�x�KQ:9,�C�I�Q�p� @�(O���#;4�C�ɀ^��lI�DR�q�1j��F�~�vC�	b@����I�&����OXܬC䉺|M&���d��yl�i��Tg�B�	�A@�uC��E����`�Z�B�ɂm�V��/@��Ҽ����RB�I�:��Z�+ ���$h�q2B�ɄE�N]�D�ˍU{�@�[��<C�I=!�6pJ�&��f��uXC�X�6:C�I�5($��FAl~�(R���h@nB�Ɏ\�0p�P�vv ! �W6i�C��6\N�8��	(d�x�[�6D�H��̋Iy���VɌ_v��Q�l"D���"E�d)�	�C�%1y�!p D�����L {��%�Gև ��S�*D�,M�<�~1����t�����h*D� ��酪t1��ᘓS
�����&D�̰���|3�EyEĘ�M8� �T�/D�(񨗺�<�!CIگ\�̀�ƌ,D�\���ؗR��A�ٞ���Z�)D�H
�B�u��VJY��l+�h&D�0;��T/	p|��sBX�wb�|�1	&D�lE5��\��A:_w�Œ%/1D�1PM۰u��x��S
h��`�+D�P���Re�	;���6/�~��#)D�l[fƙ��z�Q�̙VMt�s�(D�x15�ڠkېd��&�� ��`{��'D��*ō�.d����J�|�n;tj3D����K���Ш�K�\.�Ғ-2D��@Ť��AV��H\bg�Q���,D����m`�0'��T��E@�0D� �]� ܔM��/544���,D�\��d�PO
��a�+t~"|[��*D�� �xY���5U�Ɖ�!mJR ��"O<�r���C�h<�Ì�&(�ii�"O����Y6��$8���1}��"O��j��*��M�b�FxQ.LK"OTt
�h̪l�Pl	7oĲQ#n0aA"O<@(3퇟T�"q�7�"�"O�����$����ī�����"O8|��%\0e7^�Q�@�:-��D@c"O�pZa�%
�
4S�nɓi�m�"O���2��IL��V�<h�z�	�"O*Y�'�<fd,�`�"&2�>=*�"O� @7�G2fh��ٗ"O��R�`�	�\��a�$.g��{�"O�2E(�� �)���<Z-PE"O��eL�� �Ju�����"OI�2gH�3~Q���W�A
"Oju���|��Y�a	�Pd�4"O,�pd��|r��ځ��ݠ�)��|��'�:����N84;�`�65�&�
�'0d��t�X=`�b��A�)%���B�'}:��b`]Mo4a���!&�
�Z�'-������x�P/G�h�H�
�'Q4Ep���$�h�p	�VnЈ�'0�|+0扫2:�|�W�/&��=r�'U�}��Q�?Ђm �%-����'zܐ*�jB>�|���[4?,�	�'E��B��OYd���`֤5`)	�'��� #D����%H&�<{��)��M�jx�͊�3c��qBn���!�$گ+��g
@P8Cw"@�D�!�X�v���,Ni��D'�4F�!���>&,`y��е��\�S
G�%�!�dۖ,� y)5E��*�Z �3*�.>X!�TȦe�p#G 
�a94��{���G+D�0�Q���~�q���v9.��P�(O #=�U�W5\'"LQ�g�K]���E�w�<q�B�92X�|C��(�,�I
�r~B�.�S�O��@q��)]��;���4(:h2	�'A�P�ɽ��́���#/��9P	�'Kh $��
� ���'��5;�'�ce����Q�l](�F�Y�'�5�aU��Th0'�Y�e젢�'�NL�"�C�)�O�_�����|�<Qpe=Ϛ�1#k�>UKH�4��^�<9H_	�n�z��O�64(|�\�<鴂_A�fm�o5uK4�;�EW�<� hX�rZ=P��TQB��Q�g��B�ɚ0W$X�ba�����K���s�B䉍H80`d�=a�d��(�>��C�ɥ ^]�6���f8��Q�9�\B�I���=��J��^�<����ܮ�B�ɫ80���<��r�oϢ1	XB�	�a9���>q��r@M'[4B�ɕxk�,���Sd*�t�MGb]6B�	;A<�iTđT�~$��#Z
�"B�I�b��m9㈐8AD���NB*X�FC�ɫ
c2T���9Up�!ՄD�.C�I�Ю�B
�R�(���{yC�I�E���]�+���vO���B�	$��yjr.�y]�\hb�S�}��B�I((�`��!�,6Gx4�TGR�P�pB��l����ICiâqЧ��U��C�I"��<��Č6�����+X�b�B�I�+l����JE���� ���� >����[.}�m�%�62�`�"O���|
r�x���j-B4Q�"O� #Vi�
bf�̈�D#i|tx�"ODD8���e{�$Y�Uz@�3"Om�!��/J��7AH��vE	�"OL�#���8f|��r�����W"O���/�`���A��I�v�J�"O��IS:ڨM  �O�[t��;�"O��;�,X�����a�~��24"OB0j��-@�4h�Jt~�l�s"O��ť��=P�����36|�;�"O,5)1#�<Q\M��"<%x��I�"O�u��G�Y^�4!���Z"O�M�S#^o�!�D�кd�j�R6"O���W�O�/zp�a7㊆d��YБ"O��z%��!�x@O�?�D���"O�9Ҁ�I4ݩ�@ùà0��"O:x���Q�c�����N��m�"OP��C��.v� ƃ30��͈�"O��Y�P�>�Jq��B4V���	�"ODpAtŎ7d��b-	U�!٣"O���b�9=TM�����}�"O���^(�T�'�րc7Ե��"O��c@�ئu��Q�� ",xYRV"O怺�͚f�ΰ�q�G�')͓�"O2i���>;���%���rp*x��"O����I]� R Uk�*_bNp�"O(у�S�]W$����Cp|$!�"O2�ru�1
"��(F`�1?
�84"O�i0�H��Q�Z� �L�
�-�"Ofm�R�@]/��!kJ����"O�@s�_�(h�0#�ċ~�DPS�"O�i�mB$y~Hqw�Z�z�V��A"O:�[��W�<
�苏]��MJ�"ODE��m���N��� ��"O*]�RÜ%>��\��b!�~]H�"O�\pp^������ƅ[��MP�"O�l�㊷s�S��N����s�"O�����;s阐�%�?�Xc5"O�����?^t<veM!=�Px�2"O.HCV�_,_���P��OZ~��s"O����`R�������Dd�U��"O�X�g٧��-��lZ�Hm��"O&�*B��2dC�Z�ǋMZ8���"O xŊ��n�-���T By����'�b��8Ca�b����F.�u�r!ʯUi\q�9/��$�O���Oa:���O��$�O^Acc�r��i�a_�T�ԕagJ�)p���Bgo�uZe*� C��s4m��C�Q��/�e¹+wa�:���
�� R^���݉k��#Ӥ���
��#%�9�MɅ� c�9���^�
 f�,�ȸP6�ɪH5���հ�M����$ӼR����]�|��fƇt���Y��ٽo5 E2f�`�'aayR�N�r>�c���f�T�T�ܪ4e����6Iܘ�lɟ!��r�`L��u��'�"�S���;bR��U΅�f���	0%\u(����'�2�'BX�����O�MۦɅ�v�<$�!Bk���@/#�T�s�F9E1|@���@�h�<i��J63��i�r�1sT���&�v��|s!	�< ul�h��,2�֕�B�әM��+Sg���L�1����MC�i��V?i Q0S��ِ�±!�\���e����DY��?��$�"z�x��r�t��Lk O�H8����4_盦�i��$� ��@L+^%c.T8�U��sQ���M+��?�+���8PI�Or�dӖ5(c�A5+m�x�mӒu�a��e�t�В��P5ߦ�P�֭^~�Q��A�R�O��Ա����CE�(��Ȼp����T�iM��GCP�Yo�u�a�.�Ms$!�p|� oL6|w����A�V����C� ^+p"�Aґ�˦��c�O��o���M�������L�:�fU��M��V���b�D��~�'��mX�p���+@�9C �����01��/��M+Ӹi��'��S-��q8��F"_
5��HAT$�����?��P�*~�@���?9���?ه����r�|�k�Ny�����=��X���$%�,�q�j�YJ�[���u�|��S�P�F�іg)�� ����U�c3�P!�H�����C -��1�'#C��X  �ºc|��$.�@s�C0���z�Ƭ��%Ҵe�LA��5*�'������?1�x��'<"U�DJ�G�j-�1ѳA��y@�!R鵟|�Iܟ�'��}*�*Ǳ)?Xj$�|��A�ժ��7�ɦ	%���?��'�8i1a*Ʊ�`�Z�BG�$HX�s�H.;,Y���'l��'[Bϛ���'�d���bu�b���n��1*�W�H~B=�A��2.T����bں}#��X8,���dZ1\�!h�l����S��I�='����K�7-��nZ�2_H4�p �2������#�@�OŢ��'�D��A�.��i�w}\ܓ����>)�7��Or˓�?!��?������������^�{Ș�ygi���yr,-A��k��^n���Ǝ��~"eC)A��7�<Q�N"������O�B���ɒI�U����P)�)s���d�Oz�$؝=��TO3&�	�B��Ri�S���D��0��EH)�D��a�Ș=�t;��#H�t���D!=��	�rCƘ4Ul�+ԉ�g&H��O��R���>�b�`B�8l$��j�@�O�alZ��MS����i�:e-��8��Q�vl�$�bSdˆ]Sߴ��'��#}��Z�٪1�U>>��Lar�1����d���ߴ�M;5���6��&�_�;�~�
�Jq�'��' �O"i��  �   d   Ĵ���	��Z�tI�/ʜ�cd�<��k٥���qe�H�4M��\70<����z@�v*ɾE P4%�M�R]M�Q� �6��Ϧy۴8��$ �Ibybl� \�!����V��XS%�,8@ɲ0�PK9�=a�#?t�7M�dn8,��W*¹
�c�.2���&�ʠ�"��RG�I�Us �j3͔;���<2Jڽ��%W� 9�P&�92���Ej�6*;�v�tTx��/0�H5�V%�?)�'�������%g� $�r���9F�(�fbSA}��{��c˧~f���'�(� >0�kÁ��<�cH�y�p�I֍�I���C�+UC?�� )�Ƹ��Dy�+�	�0����Xg7�	�q:\	j��W�8����J�6��#�ߢi�~�@���δ�O�y��?l�ڠ�ጔ\^8E˳��X�'���Dx��A}���	���ɲ G=r�`��+����ɱz��;��$�/��*�:Fu12�V�+��j�K�'�@�Exbb�2G@�`�+cx���13�� �}��LT�'�pd�'�ر�BD�]Y��H�!� Qhh�k(O�d������'/�� 7�,h5R���#@�u�N<�-�t�'��Fx��˟L@c�ýV���6���@ܙ��/>�I���쉂�xr���%�6�J@�=7"�-�~B��}�'�i%����'��U[���CK8eS�էRub����v�I4���	��iݩ��rD����y+pm���1-Ƹ��%S���'�\%FxҎST���n��N�(Sb�!H�AB�P8�Iv=�x�1�I>H�fak���0����)26ۘB�I?t� �  �7j<C���Ci8,|�)h�E&}r{�'.��=1UI�jR�IJ�!v�V�"2��ʦ݊�ቮ[N�dхĉ� �����I4]q��P��8
$b�TS�I�j��I�5�A� ��܅0�cL�*��� |�#<�`0�	�O�TaAFS���bK�#���t�Ɉ`�X��'�bh	w�N�[�:}X�G��>(ybHJW�'��&�t1�f՗,�<�1�� <dXm�������	(S'�'�����h��OB l,����b���xy��Z@?!�l]?��	��� \w��H�A�
h��'i w�)����;�O���H��b#��KF���Q�6�tD͢>�� �4�"<���5D�ThF�H�_2���A�<)@�� 2  ����C���q�.D�l�#�    �	       m!  �'  .  >3   Ĵ���	����Zv)���P���>��'���qe���OT|#�j�9]ֈ���
�*U��r"O1�4ŋ�/^LPi���0HEfIqJ�O_�����+�\#��i�,IP4�4>z�Qv��:\m6�1�I�Sg�-e��4MD`ri�i�rA���o�B���I�^p8���O�f�Q櫁�d��k�}�"�Xu��s���*_V0d�2#ښ!=���$�89�]ەNL&M^q�&GD���	��	ßభ�:������q�de�1a�v���l\y�)ߍO��q�2�'ˆV:)4��a%t(ՙ�oR.�:m�QE\[08q�ۜ���'F�Ƞ� 	Z���"�����Z���񖂍�)Ŗo�ğ8�A�ڟйܴ)��<����~��W�1���IhV4�vM"�ɳ�y�O�qmV� iT'ޜ�2� �M��qsV���FyL�O�}(W�+C3��C���`;��yռ�����?����?�`��`�d�O��%�z8�[��>Ղԣ�0�� �i�-M����S�߶x=�b����O��k�Fd�|�{!��TB h�@��0k�-;%���@�B Go�bs�3b�jz1h!��B3b��-A$C�6b_� Þ�%�Z6m�æ���yR�')�O��W/X\���It��P�� Y�0B�	�3I��	f�m��)զ؁��(��	zy"���B��7��OB�d�?���/ם^<�4�� >����r�}�6!	��O|�d�Oj�f��P���!mK�w�l�m��F�:%�I�@��:tP�X2�m�'��x�Ah�`t��2/� T~����I`Ս]9N���)	BTH̥ ��	�s��D�OJ�o�꟨��$ �Q+��9s"��p�n� �v����9�i>uGyF?)���r�]1/���
q��M���?y�ʟ�x�'5�p�D�Ɋ�R�bĨ�Y�pYg(�>A�	J9B����'��'��D+G:Yb�'t�� �C�cQ��S�L��-��mj��)a���O���?A/��O2��`��n2x���ؗn��y���'�"4yed�-{�Z��E�ѝ=��?��S,ڕ1#�9���7P����ȅ�H3��OZqo9��T>�Ss�t勳[:��SQ�T�,�����ww����I؟H�}�qjSu��J�r��)3��W��?QZ� �'S�> ������8/:�@����<:-�Ȓڴ�?)�?4p[�����?i���?q��}u�n�O@�F�T�MRRp:s��2L��Ѓ�ڈ^�����3�&���F-�`	��(OD�ٷAԭSv����X2x��`Ps��J|��%XsP��d+	�6�3�]Ĥ�wȌtC� s��~�t�'i�y��?����'�	׫x���q䫎 F܂�����l[!�Ē�tYP �3�Da�hPGm�+7Q�f�4��|���������a�	%Y��`���=D���Rcɒq����O����O�����?����į��DN�ĺ'o�-/��\�����~�P��6�׍Yv���@�Oqxȣ��(�yцh�S��T�y�u%�iK41���D�O� ɤJ۞l"�T��]�p��`"���Od��%�)g�%±fUL�bZ��Ʀ�G{��ɅS\�8q��:zA慹'��m��C�Ix��ztB%/��B�s������'��3��p��J�D�?�Zŀ�F��P���� [�XHvCo�B���H�O��d�ON���	��hI�A�A-h�ԟ�R@C@=_�����A��S�ؙA�ɕZ��`qS-��'4���d��� B��Bi�
���<@�Ņ�hO�=�@�'n�6M�@�'="�	p��'h�9g�ھ0����'�R�'��%ӵ�>R ��+�It���
�Dm�ɟlS&a��iD�k���i�eϥp�j�lc�\B"G�;���V�G�	Ӱ�GzB���=ת�K5B���HjaE*�y��U�֝��A�|-�Tۅד�yBRb9S�B%&��vgͦ�yr#ψ`:���wH@�T�Е�yR�'�	�n�P��)�(��y�b�#�L1v	T">+�e˵ᒱ�y���B)IGa�h4B��	�y"/(5�bh
��O�C�K4E��y2FZ{FhKB([�;��� �"�y"Ƙ�V�B���fP`�H��Tb@�yrI�0�ޕ�JݘNF¨xdh���y"��<B�E��b		^�T ��]"�yb�D<%쾕I�m�:���MC
�Py��8j"�z�F�-*�`��u�<���c�����0b�n�8�]N�<�Ь	$���:�a�&s�h�j�F�<� ��j�H切�0�6Y`�ďC�<ɤo��w5��0�ߵ/Ң𳤘_�<Y�*���9J�À�x�`��B\@�<� �\0#�/dhlh �>SgE��-�3p��C$�Ζ&b��2w�i?>#|J]�<�$�V1��%��L�@�X4
��1D�
rI�14H R���k#$yӮ�2�f�)� ��ɆP-$*�	�]�H�Ђ#Z�̹�"a�qm,�����J�\d��ၨ���cGΎ� ��P ��\)J���x�-�lh�� U؟P�󃅯3�y�Mۼ5�m���3�ɬ?"m���5��;Q��'�47��d�L*Q���ABG(a  UŧJ�y�AE�Q�&��T�]%#�@y�D�BG\�tWi
�o�\T1t���M���?�sS���?Q��O\m�.A'����cYv%��'�v$��Ŷa�l� �7V"U�΂�L�� !�i  �ĮK�j�RYQ�M���Q���H '��%��&�;m����Ì�O�Q�����X gh�$��.�+M�j�	�Ǆ�o�s�
��Ri��0P�X�2�
S-X��@Y+�BS@؟��" ���с�ޟmW���Ic�@��(�~������B#y��i�	L8
@r��W���s���o�� n�p7*[L.�Uq�a D��@�
ߡF�@�h�"��=��<����pkFܸv�2y��f�����O$@�j�*��}-�=��O��Z�)P
Q�&q�6|����'��HP��9���7_��s�ütL�	���ɾ68 xr�����J�`��z��j��7��Onh�@Y�@wP�l\�O8=��$ՇBrK��@J2��
�� ��|+��0,w�����1��BnC�@�S�4>���-(�O(L�#�!@.�=����+�@�����2 �U�':���g�H�PP�"�Oc�ܔz�����6m�Q�4��& "!�'�R7-��:5++D�0@u���������w"#t�@C6��/X�Pm���������x��&t�4u�3B�>�ǅ_1-� ��ȷr���2�]\8�0���� 6��p�SdȽO�~��@dD�g���z ��*)��� �G�/��zĮ��'����o�]�'+F�q֫إz@�1[�B�}R���d?'=�\�l
�5�tpY�#�^k��pT���Î0�Q�J+gC\�h�MPkU��Y3� �O��v-\��#�BRa�<O���q�^q�n�"�(�`�L�t=|�h!�]�S�X�*q[t,Q�Tk�I�4x>B�Ix���׫Oz\t�>`�3"����׫N�hA�Y	pc�S�ft��.i��1*�O���P��M�f��q
B
�4ب��')4٪�M^�N%R�`�\^"ؑH3O2g뾽��*ͺAVJ��'���p$r���+(�R�F~� ��n�L����1H�@uUhЄ�HO&MQ��\�?�w��cຈ+6l�$%Ltj�F�ސ�ʝ"G[PL�wA��vX�t���'�V�J ���iɒ��w"��{W�� cU�D�|X���'gȸu��!�ִK"ğ�I����t��w`�`Ĭ�W���Ö�u M��'�:D�c��
k
��rvDCC�K\F Y����1J9��(ݴH(��� 0+��2D-�����T�H�G�]�q��](�a�.��!��'�O�q{�9�$�mywF��� � "tR`�V�w��6��8����"��tSb�^�W�J`���dSZ̩�e�]?*M䘒�Lӷ/#�h��mԆ^4�Q���G(y-I�p��rDL����#!�d֎z��,�� &T�~4F
�7�V'�%�`�|���i��a���v���
tdU5&��y��'�8�afO݉~]�p�o��\�2r�O��1�/|O\u�ELI�#3��r���)�0��"O���e@�c�@�W�`��"O挻�&M)C�8�!ᇟ<)U�ā"O�,�ǂº6���� �%d���y"��nP��m��.z��������yr�B�d��Q���+!��aѡ쑓�yB`��L�L���,L�e}z%	���yRd��H�ѩ�,<�`����y��_W�X��ƀח���eCG:Y�!�M�[x� gΈ)5W*Җ�@�H�!�d�xLʑ����Lg�@[��� [�!�D�>@�Qp#�U�d��*��!��8��H��V ���f���{�!�$�<��q N�_��A�L�v�!��S%o�S�G��0� *�hS��!��e{
D���Z�S���BC/�!��2t����Vl�m�J���қ6!��L=�T�E!�f��@'� r"!�䔌9�ȴau(Snڠ���T�A!�ǚ<V�P��ˎ.fL���'R#Mh!����\�U��)QM�x�u��G]!�� j�8eX�*9�l�p��$#V.��&"OV�$J�$YU�<�q��4y�P�"O��7��aN���X�j�c0"O��bg�0�p��l?#պ���"O��e`��y�F\+eͮb6vy3S"O�	s�d��ԉ?+"d��"Oz�����]�u�%k�7���آ"O Tb��E�t�`r6*ע	�>��"O�eC�ɒ�z�r�Jw��'REA�"O����&�'y�@K�HԡW&B��"O�q:�mЇI��%P"�Ëf& ���"O%��f
�!�H���>'
)�"O8�ъ=��`DKJ;E�q�"OV :���a���'�}��"O�u:≚6�ލɅ�p�(� 6"OR���_�rqCFћ'Ot@@""O���VjTw����n�
 A���"O��c�� n($|��\�BxQ]6��O*�}�>d�,�UGI�Rx�m1�J�{��t�ȓ{ �Zp,Z��i�Ui�]hL(�EG����'�Ja��f&�Q���[4CA�ד3����@����VANb�l�J[�)�"�%�B�I�#��Q�C
J����*���O�����
Zy�u9Fd�J�O���� o
Ta"�2dEr�	�'�Eâ�#I(�9�鏁\Ӣ0S�BAp��<��j�O��1%���� �D"��T�Ln2�;��߇/�����P�;�J)� �O�P7:����L U н����KR��	q�'�{�²�O���a�p�@�����U��D*�[��Աf���b�C]�2�m���[�y?�B�I9(3�!y����g<b< �-؝Q|�Ox�zD&K�{���(mdo<9F�dg����Rf�H*%�B�0�:�y�.�tg��*Z� �qĉ��mBqHsnQ� ��a�?h��L~�y&�����3F���HY�pR%L��?! .��B���a�@��Y�@�9�.Ep��Y]F> ��J� ��w�'��,u��0��|z�Iul2�b��$ĽB��݀��=�԰ˠ��~�B��CcK����T�ވ���Y1=)L��� 8&� ��yS���h�:
V9�'��L[�R�j(9Z��	pIs�t��WcLI��"��Jt��3�D<��O�
�
���x�����l����� ���`����"jӐl�F+�?��~8�'X�� 7�P�+?�`�	�4���M؀��A;mQ���'�Q�W�,eu��yo��-O9�Dz�B�g�y"�N�p����êb��•L'��Oz��3c[�O+�|�w��r��נ�/a�T�r@�v	R��4��.�TB�ɄlM�1卑����ـ|
�9���a+
�A������ |&�0D��@�h�l�2�uۘM����/�y�$�J�@����:h���S�A�a�P�JX���)���|�<�0��<T�H�ɰ[P:Y��OW�<�D#C^,��Tj��J�����ȃ֦�a`��%4J��P��v���k���AvfM�daI)lOέ§��l�`!�Ӽi�(��q�I�`mjAhe��W�T z�'��-�$A߃_ �A &�e[�{�A��,��f	�h���G@�Z0��H?��u"O���Br�q!�S�dp�d��o8��"�xr�<�g}��ەk���Q�L�c��H�rݮ�y��S�a�.x³�D=3�D����:4B�|{N��d�=yd	�ŎV�V)­q%�-o;�{�*�:Q��I
�)� 62Q�h�4�C�	�;����Ŋ�܁��լ?�$C䉯#�H��ea.	��Hsa�<S/$C�I�- ��7�F�vw�䐶��,i�B�	3��d�Ɔ:K�T���T$)�B�I�6Jvɑ��Iw�d��7|�B�IX�>�B�1@p�3���Ii�B�ɤjD�(�g�:T'&�ޜ.�B�)� �q�s�QO"Ց��^�7 �p�"O`�Bc�U	rʈ�ABg��Qe6i1�"O�s�(�N<ԡF(׶!���+p"O�*�`�	.�����(J>�Bݳ�"O�m�Q��%T� �&� ?�(��"O�\1��%Lx����b38�lR"O�]�f���l��#LU�*M�P"OLē��}#�܀`L\HܺB"O><B�Bч����!@�+kB0!"O�pC�C�,�4�ɑ/�'�<�r%"O�L�b�Q�$� A1daP�R���"Op�0C��M����(3���"O�l��Q�eI��2eG���0"O�*Ó,9!���c�;_B©�p"O �"��43���D'�z����"O:��5�E�j�ti���ӑ$�zh��"O�
��T�Y�|�Rs^M�.�:�"Oʰ�G���ږ��8j� P9�"Ol�0��F�.e���	��qP�"Oq`�FRo�<i6)�?��y�6"Ob��3I�������;����LW�q �[|z  �1O��܆ȓ7�� !'Q#M*�Hu�^
#�I��G3��tn�%"���sSf��1�<�ȓF��i��g�~Ũ��{���ȓ�ެ���Ů2i>�KV�ٚń�]:���-a�x��`DV�pp�� h�h�A�-6��#�h@�S�]���A�U9�rY�7�("��ȓ4�>=I�kI"�dx4	+xǶd��D �أ3�G)y6 0@PO�I����cf���!蓉,�ΐ	s�׭``L���h�8���W�:��R#�^�R�؆ȓn�hؐ��o �Ś�EM�dl�(�ȓ}  �P6C�?���&��#
�6a��ӢP&ݣGR:�iҦV�^� �ȓ?���0�G[�/�����z�숆ȓ<p���5eH:/w�Ys�̉� ��ĆȓC�\H$�0#�r}���/����ȓ�F��aFE�OP��ecʲ3)�@�ȓFo0!�WmFm�x�2L4E~5��wz���#O��0 .[�{�܅�sUB�b�T}"�GJ(2
��g���c`�U�LsƝ�	�N�t���9L�dI��wU
�P���	;�2�ȓ
K�����z������� ���tz�)�%[�W�>E�En�_�Q�ȓ[9��eM��rH v�Ƨ;����ZU@x��dy~-�%�	GHN��'�X���l�<Q��8Cp��
`�tb��ě6=�,EH"�@�(06��aDP�!�Ĕ+ZV��ĭQ�b��Т��Ԛ_}!�	�M�:��$���!����L�e!�$�>����'�I�RQz殈�U%!�DQ� �	�0Jn��y�-ն!�N=�8���6����uk�(N�!��Դ��i8F,֞%��ꃠ�y�!�D�d`)�'�O�$!B\�P�!�A�2�4ړ�	�|1�4��W3!��ƛL�>�tK�&6�*xB*ė%G!�Ċb�8���S�tySW��&-!��*�BQ��/B�qۥ��(!���ՠ��!�Mcr�!�p���4!�ٻ^Y���L�4d�0,V�g�!�L�pLh&J
ZQ������P�!�� �(s�.B蠕��a�lT�!"O�Di!BR�0w��hB➂sT0�1"O*5�F�ژB!VHӔ�F�|fnMb "O��	����@<hs�W LW��J�"On𒖯��hԖ{4aT�s��PV"O�,��cV7
�+�J�<x�<��"OV���. �pp��j@j.+\T��6"O�8F�j��0+!#�8	�& �&"OB���^h�\�â�HV"O��XC$�7�eyE� x���ib"O���ID*@�n��bͧj���"O�����	��� ��D��qI�"O\��a�!il�Y���=�:���"O��2TMJ�|3n�h��ݨ��g"O���G��k��-�ciZ%��tK�"O��C2�ڗqa��)WSʐ��"O4��"�u�f�V�Ѡ)�vӒ"O�`� �c�2��)UXwDɣU"O��ȑ��G����Ygr�#a"O�\�C���Z�� H @|��.�!�DRt?bM#aJ,1��Lx��M�!�$�
t�<K"�S5f�9�FE�?�!�DU�~��r���+8�� ���#=2!��<1�n�P�ŶP�c�E4_7!�D������Z'����!\�!���J��a�fLJ|�>�1U���!�D��f>(�&�� ���q�!���pH�"#���#ӿyO�ȓ%E�`��oJ�����\�[����@���
�lG�g�q[�-W�`z�E�ȓ �Ax�%�Bb};ƧU94_>��ȓnM��jC�2,�ITG�~Zhl�ȓM{�=�PӉ<2���S�1v�ȓl'Xh�U��_�z��ӌ�D�и��J�呥D>b.h;��W=T��̅ȓi̍���I�$�4c�ʷ�B剭9HK	; 2<��M&�Z�f"O"�/�L�Ul x��'@�l�C�Ɂt_8C�l'^زa!1O«FٚC�ɉP��Ѩ��u�!*���f/JC�	98�U{�mU�x�n9rg�+�C��2H�Đ����:V9��%ч��B�I>W(t����f�$��f� �B�	�d�.0��1?^i��
�K4B�	\�^4��)[*e�J!R��(;�C�IV�Bǀ-i3>���NEY�B�nj�A�ʻ#\�x"� �TC䉅iT��%�<� ��r��yNC��\Qn�{�K:E��\����N�B�Ɂ �����\�0�|�g�^�u޸B�	�>�*�h+'�`�B�_�^��B�ɹ��9��h�>f�P�b%k\�&��C�I1<��e���Z�Ia�rE		�HB��,j��uZ��^�?�Ԣ�"�eFB�I5?cD��)U!"*�<�9�nB�I8tJ��ʖ�U�C�T�җe��
�BB�ɗ,�(��E;l.􂄂�j�B�	�^`��!���L��B,?T�C�I"l�bA��m�����QBD�]��C䉱�6�����V#�ZcK]k��B�ɌrZ�P8�@���u�$��|B�		'���i�L��e�`9�vi�(��C�	�w#)�P�:հV	Ç^KB�(��f\r���$�.��C�)� �<�'��!8��9ňA5��#f"OF��pC��4G�M:���f�Y�4"O���P��5|Pܩ�AP�s�� �"OdP�#�Q;Sr$ŨS-WR�@#�"OD�C�����[#��X��mK�"O0�5DF7�Z�r��	�(�����"O~�`"��1L���˧Z9�D��"O@L�F$�61F�Шg�-#<P�b"OV��Q�3����속Q"��'"O��9���SX� !.Z����"O�='��Xe �̋<~h8e"O�E1�)�*f�IR)��~V�D�"O�Z@�\�sx<���fB��s�"O��A��6*��qg��8e9�PXd"O��&��q���1W.Ʊ4z�`�"OfdXC��x<I��=gr���"O���֬ў3��H�2g�W�D�"O��[��+�JU�0'�8E�P� "O�m�RJ�h�!�Խin�j�"O�x:E�:;��sV�ޕk�]��"Ol��ѿn7�@z$��.s���"O&��b��Y�%�T�A�@M*�b"O4�v(Խ#��(�d��?�e"OZ4:�#7!��2-Lip�"O�� �Q$f��T�_�/,F�0��'��'�t�Hg�LP��}�E+L�9~}��'g�}��d�'���	��ʉ�f]��'�l\��L�aZX�QC����	�'��Q�Iy��Kb�Յ;�=#	�'��=(���)����!�_�GJ��'T�͛�dR7W$�<�D�W�;H�'������?C(	��b� ^#���'�H��ѨA��eP��& ~U`�'
����K�x��QMނh���*
�'��=��΋J��F��n����	�'���jց�#S�EaU��t���$��%�OXq:��N vY���E� \����P"O�t���Œ_��h��=F��"O������NHl8+qC��tL^4��"OT�K��G3g�����U�d�F"Oz���]?�P�r��(a�m���	�HO�6p>�H�`�7F8�|�çM%?#�B�I0LQ��JGeS�d��JB.��I��6�%�S��M��AK�a�t�[U�Z�)�����N�<�c�M��Ie�ĩ�"���	K?�F�'��|8��H*N1!�1��9	�'kx0��K>,(�!p�ń-à��ʓ+��� A�9���1f[�QLP��ȓl�"xq��(M$d�P��C�B��X�ȓmw�!`��"���5��5=�,ԆȓE��x�% ���$x��*�-�&��ȓM����$�U��hk7@6	�h�ȓc��=�cH�-Xt$Hm(�ȓ\�`�P�M��pċ�Ӿ��l��/\>�s�0M����e�ws� ��%��1��]�İ��
P)9:Έ�ȓ`�V=:b!�w�Tm:ǐ!nC@���y+j��0⏂z=�8jX�0��5�ȓ�>\�7���&�i�Ɲ�t�@\�ȓ9��B�n�P72����	*��݅���m*'E��2��@S �,�Ԥ��a'6E1wG�=1�E����(\F���74��3�K�1(� }j�F�"J��ȓo����AV|W�Z�d�U52\��S�? �!ʂ�̉;��,SwaA Aj.q�"O(y
��Dg����v	�!5"O�H��Ԭd�iq�"Q��a0"O�=�L!q��`���P�$�0���"O���DV���H`�����;�"O|�!UcZL;ƌ�%#ݝa���"O81kEV:�x�AtAˤ=�x�"�"O�!e�ϝX�$*4�_�f�&�1�"OJ��5苖)�x,9`-�"x��QJ�"O2�b�HC���F �#h����"O���3h۸H���R�J�>R<xv"Op�sq�>J�Z|	��Q#9Q�И@"O>1�J6!�M�4g�K3T�K�"O��(%A�0+�Z�����||ʅ"O씪��T+ M�9r��q�,
�"O��0��^�h#�F�!��"OZY+�Z�	>4Q&�O�a"��"OhAW+P�b�М2iT4e����t"O��d��%2��R���r�	�"OU�҉8!;|qIWgS����"Ol\�g/�"r���+sd�	0Q�"O^�٣b]3~�=!�C�LV��d"Oz,��O�d_&x�(��bKz1�"Ob��rj�8�%D��+�"Oz��4ჍP��A�᪃.,�6��%"ONĂ���k4���O
y�6d�r"Ox���ⓝT���#_=��!��"O6t(2��\萕��	�+!�~��"O��r�)4���i��ޑ_)��2"Orm���KB�U�Q��	B�A��"O����-#�j�z�@�"?2({e"OE!E)�*%�ȍ�յxZE��"O����#4�X32�Ěv]�ɉG"O(b�нJ�rt�r�&O6�*U"O�:�@�U�`���L�=d�T@�"O�܁��Y**�����N3�Ĩ�"O��s%�#������0(Z��D"O<��b+G�VEb���}p�m��"O��K!BJ��$xR��C�E�0"O�Q$�]-Mz����� #�8q �"O�	'H�bL�r�P�n�j�"Ov%h��-�-��o:��6�3D��3!K�3.�^��t��B���d�3D��:ևM�(I8R�ɺa�� ��=D���4�݀��U��+}��h�!:D��
`C\�A�1����=CSg7D�DI�Ւ�م�}�ʹR��0D�p�� A/~�R]A��;_��5�0�*D�p�bj ���y�e�D�y��8��$'D��"�d�;����#GΦ�ʣ($D�@zVM�eR�t3@4u�u� A"D�T Ԃ�)^~t��K�8�Ni5�2D�H���;u���1�
�*=xC�F%D��   �   j   Ĵ���	��Z�tI�.ʜ�cd�<��k٥���qe�H�4M��\70<i���:G�&�����0E�5��y��cA�6-Ħ�q�4x��$"�	}yr��2�p�Y`f�lٖ�&�H�܋'왭e�a�=��,)�=`6�ĺ)Π9Q�$�x��)xׯ;w<�ɋI�q�ǩ�{���(�8YvN �q�	 ��U	"�$q�Pa�� �`����[$��͔9,�%�	�Q��`�d�?q��'�0�%ڱ��E�*ߓU���p/�EdUI��A�����d	*3�i��! @9OT��U.
e,�ɏ]�����b�&�FŉrP�G����d�����Au���t�nY�t�P(H����OF�����BTƕ+u�ҸuG=kՀY�[H�a"@\�Ƹ'0�Gxrk7�YP"F�]�CF�p�p��	�*���a�Z��h�����ڔ�290�x;�6}B&V�'C�X�=�SDZ��`�W�\&0��bb���b�ቮ^���%dV����!�c�(��Z	L�Bc����A(��NFM8�%=o��*E�)v� �'�B"<�d!���2,<��-F�+U�"���*>"4(ቻ��s'�'즥���Gb:}���HW|I��y��y�'�~�'�xa�ժ�r�ϼ@�(@T� <�~���k�'��M$��s�'���Be�1]�X$��*�/F���C�+h�ɄU��	��i�M��Kp�dņ�I�ɠfQ���s�O���'��Fx�
b�DN� n<�2�� C6��d,�I�@��`���I��0���E�W)��a���	dQlC��5>�� �  �&4D��ic�OZ&�g�{K���"�3D��2�g�*�~|���'�Xyw�.D�|Hb�	;_��dy3c��W�@��4,D���n�����[	T�9`���ybO�5V�y L�1&��;T+�(�y�B�2�`�F�_�.H� �#�y� C7)��q'�\�(ke���y�l´uB�5I����X�H�HMJ�y�MZ�E%R�RþP���¦R��J�'������=�\I"�iĞ���Y�'�|�T�K&��I�Q�� ���Z
�'�N�E� �� [�@�H��)	�'��C��W�l,��瑄\�����'U�5A���o�C�F]�i�8py
�'j"��`��%:p(Yǋކw��$��'H:)��ω?��j6���i�4��'ðĠ��M�F�Q�Ի�    �	     (  �!  �'  .  W3   Ĵ���	����Zv)���P���>��'���qe���OT|#�j�9]ֈ���
�*U��r"O1�4ŋ�/^LPi���0HEfIqJ�O_�����+�\#��i�,IP4�4>z�Qv��:\m6�1�I�Sg�-e��4MD`ri�i�rA���o�B���I�^p8���O�f�Q櫁�d��k�}�"�Xu��s���*_V0d�2#ښ!=���$�89�]ەNL&M^q�&GD���	��	ßభ�:������q�de�1a�v���l\y�)ߍO��q�2�'ˆV:)4��a%t(ՙ�oR.�:m�QE\[08q�ۜ���'F�Ƞ� 	Z���"�����Z���񖂍�)Ŗo�ğ8�A�ڟйܴ)��<����~��W�1���IhV4�vM"�ɳ�y�O�qmV� iT'ޜ�2� �M��qsV���FyL�O�}(W�+C3��C���`;��yռ�����?����?�`��`�d�O��%�z8�[��>Ղԣ�0�� �i�-M����S�߶x=�b����O��k�Fd�|�{!��TB h�@��0k�-;%���@�B Go�bs�3b�jz1h!��B3b��-A$C�6b_� Þ�%�Z6m�æ���yR�')�O��W/X\���It��P�� Y�0B�	�3I��	f�m��)զ؁��(��	zy"���B��7��OB�d�?���/ם^<�4�� >����r�}�6!	��O|�d�Oj�f��P���!mK�w�l�m��F�:%�I�@��:tP�X2�m�'��x�Ah�`t��2/� T~����I`Ս]9N���)	BTH̥ ��	�s��D�OJ�o�꟨��$ �Q+��9s"��p�n� �v����9�i>uGyF?)���r�]1/���
q��M���?y�ʟ�x�'5�p�D�Ɋ�R�bĨ�Y�pYg(�>A�	J9B����'��'��D+G:Yb�'t�� �C�cQ��S�L��-��mj��)a���O���?A/��O2��`��n2x���ؗn��y���'�"4yed�-{�Z��E�ѝ=��?��S,ڕ1#�9���7P����ȅ�H3��OZqo9��T>�Ss�t勳[:��SQ�T�,�����ww����I؟H�}�qjSu��J�r��)3��W��?QZ� �'S�> ������8/:�@����<:-�Ȓڴ�?)�?4p[�����?i���?q��}u�n�O@�F�T�MRRp:s��2L��Ѓ�ڈ^�����3�&���F-�`	��(OD�ٷAԭSv����X2x��`Ps��J|��%XsP��d+	�6�3�]Ĥ�wȌtC� s��~�t�'i�y��?����'�	׫x���q䫎 F܂�����l[!�Ē�tYP �3�Da�hPGm�+7Q�f�4��|���������a�	%Y��`���=D���Rcɒq����O����O�����?����į��DN�ĺ'o�-/��\�����~�P��6�׍Yv���@�Oqxȣ��(�yцh�S��T�y�u%�iK41���D�O� ɤJ۞l"�T��]�p��`"���Od��%�)g�%±fUL�bZ��Ʀ�G{��ɅS\�8q��:zA慹'��m��C�Ix��ztB%/��B�s������'��3��p��J�D�?�Zŀ�F��P���� [�XHvCo�B���H�O��d�ON���	��hI�A�A-h�ԟ�R@C@=_�����A��S�ؙA�ɕZ��`qS-��'4���d��� B��Bi�
���<@�Ņ�hO�=�@�'n�6M�@�'="�	p��'h�9g�ھ0����'�R�'��%ӵ�>R ��+�It���
�Dm�ɟlS&a��iD�k���i�eϥp�j�lc�\B"G�;���V�G�	Ӱ�GzB���=ת�K5B���HjaE*�y��U�֝��A�|-�Tۅד�yBRb9S�B%&��vgͦ�yr#ψ`:���wH@�T�Е�yR�'�	�n�P��)�(��y�b�#�L1v	T">+�e˵ᒱ�y���B)IGa�h4B��	�y"/(5�bh
��O�C�K4E��y2FZ{FhKB([�;��� �"�y"Ƙ�V�B���fP`�H��Tb@�yrI�0�ޕ�JݘNF¨xdh���y"��<B�E��b		^�T ��]"�yb�D<%쾕I�m�:���MC
�Py��8j"�z�F�-*�`��u�<���c�����0b�n�8�]N�<�Ь	$���:�a�&s�h�j�F�<� ��j�H切�0�6Y`�ďC�<ɤo��w5��0�ߵ/Ң𳤘_�<Y�*���9J�À�x�`��B\@�<� �\0#�/dhlh �>SgE��-�3p��C$�Ζ&b��2w�i?>#|J]�<�$�V1��%��L�@�X4
��1D�
rI�14H R���k#$yӮ�2�f�)� ��ɆP-$*�	�]�H�Ђ#Z�̹�"a�qm,�����J�\d��ၨ���cGΎ� ��P ��\)J���x�-�lh�� U؟P�󃅯3�y�Mۼ5�m���3�ɬ?"m���5��;Q��'�47��d�L*Q���ABG(a  UŧJ�y�AE�Q�&��T�]%#�@y�D�BG\�tWi
�o�\T1t���M���?�sS���?Q��O\m�.A'����cYv%��'�v$��Ŷa�l� �7V"U�΂�L�� !�i  �ĮK�j�RYQ�M���Q���H '��%��&�;m����Ì�O�Q�����X gh�$��.�+M�j�	�Ǆ�o�s�
��Ri��0P�X�2�
S-X��@Y+�BS@؟��" ���с�ޟmW���Ic�@��(�~������B#y��i�	L8
@r��W���s���o�� n�p7*[L.�Uq�a D��@�
ߡF�@�h�"��=��<����pkFܸv�2y��f�����O$@�j�*��}-�=��O��Z�)P
Q�&q�6|����'��HP��9���7_��s�ütL�	���ɾ68 xr�����J�`��z��j��7��Onh�@Y�@wP�l\�O8=��$ՇBrK��@J2��
�� ��|+��0,w�����1��BnC�@�S�4>���-(�O(L�#�!@.�=����+�@�����2 �U�':���g�H�PP�"�Oc�ܔz�����6m�Q�4��& "!�'�R7-��:5++D�0@u���������w"#t�@C6��/X�Pm���������x��&t�4u�3B�>�ǅ_1-� ��ȷr���2�]\8�0���� 6��p�SdȽO�~��@dD�g���z ��*)��� �G�/��zĮ��'����o�]�'+F�q֫إz@�1[�B�}R���d?'=�\�l
�5�tpY�#�^k��pT���Î0�Q�J+gC\�h�MPkU��Y3� �O��v-\��#�BRa�<O���q�^q�n�"�(�`�L�t=|�h!�]�S�X�*q[t,Q�Tk�I�4x>B�Ix���׫Oz\t�>`�3"����׫N�hA�Y	pc�S�ft��.i��1*�O���P��M�f��q
B
�4ب��')4٪�M^�N%R�`�\^"ؑH3O2g뾽��*ͺAVJ��'���p$r���+(�R�F~� ��n�L����1H�@uUhЄ�HO&MQ��\�?�w��cຈ+6l�$%Ltj�F�ސ�ʝ"G[PL�wA��vX�t���'�V�J ���iɒ��w"��{W�� cU�D�|X���'gȸu��!�ִK"ğ�I����t��w`�`Ĭ�W���Ö�u M��'�:D�c��
k
��rvDCC�K\F Y����1J9��(ݴH(��� 0+��2D-�����T�H�G�]�q��](�a�.��!��'�O�q{�9�$�mywF��� � "tR`�V�w��6��8����"��tSb�^�W�J`���dSZ̩�e�]?*M䘒�Lӷ/#�h��mԆ^4�Q���G(y-I�p��rDL����#!�d֎z��,�� &T�~4F
�7�V'�%�`�|���i��a���v���
tdU5&��y��'�8�afO݉~]�p�o��\�2r�O��1�/|O\u�ELI�#3��r���)�0��"O���e@�c�@�W�`��"O挻�&M)C�8�!ᇟ<)U�ā"O�,�ǂº6���� �%d���y"��nP��m��.z��������yr�B�d��Q���+!��aѡ쑓�yB`��L�L���,L�e}z%	���yRd��H�ѩ�,<�`����y��_W�X��ƀח���eCG:Y�!�M�[x� gΈ)5W*Җ�@�H�!�d�xLʑ����Lg�@[��� [�!�D�>@�Qp#�U�d��*��!��8��H��V ���f���{�!�$�<��q N�_��A�L�v�!��S%o�S�G��0� *�hS��!��e{
D���Z�S���BC/�!��2t����Vl�m�J���қ6!��L=�T�E!�f��@'� r"!�䔌9�ȴau(Snڠ���T�A!�ǚ<V�P��ˎ.fL���'R#Mh!����\�U��)QM�x�u��G]!�� j�8eX�*9�l�p��$#V.��&"OV�$J�$YU�<�q��4y�P�"O��7��aN���X�j�c0"O��bg�0�p��l?#պ���"O��e`��y�F\+eͮb6vy3S"O�	s�d��ԉ?+"d��"Oz�����]�u�%k�7���آ"O Tb��E�t�`r6*ע	�>��"O�eC�ɒ�z�r�Jw��'REA�"O����&�'y�@K�HԡW&B��"O�q:�mЇI��%P"�Ëf& ���"O%��f
�!�H���>'
)�"O8�ъ=��`DKJ;E�q�"OV :���a���'�}��"O�u:≚6�ލɅ�p�(� 6"OR���_�rqCFћ'Ot@@"��.H�$���J#s�Yi4�G�uaN�25M�@�!�$��pD��Q���N/��z4
�J9	Cl�|�	�
�Q>�4���",S90�F� sAN�hͅ�Ax�H�Z�j�v-F�o������DH�dcԥH���&�U��\5���B$'�H����>\O�)��Y�"���'�Hh��VW�	)��&`�$��'�����j�x7�E���Ex��+N�$��e$D�]�S45WT�G��q�p=0CdP��� _�y�g�������mI�k~�x��닝�F�h��Z��$��=��;��L>၎�ͮ@��+�26r~�`�Da<ᅆ�6���8"'� {�1�dpԴ���c�r��o1ɶ��������G B��<)&��J�ax�-M� ��@�Y�pi�T@�o�'��4����D-��{I*Pj�'�քsaI�f�6�E��r)�V�<ic�0�:}"�
"kօqiY�����KjZ5 *�
#JԵ�PQ�v"O�9&"���i��#�tmV �w�α#����%���{<�MB�n0<��O�1O���f�=Qy�$�,����!�'r����|{���v,
+c�����9�q³/��,G��0"*1����D�Y��ؤq:� ���Y�k�џx��j�0������'�`�2J��kǀ��+��zA�M	rGX�pϦ�
�'�2*R�W���ݲ %ִg�Tm�,O2 s��S��P�m��L�U����Of���CӔ��C�-Y�k� �'��0��H������ĉ-s�<u�� :䰛5�_˦9�aƋ�n��OT��O"�)gÂ�C���ڐ�To�YS��'�"�+cˍ�J���Y0E�6i�:b�
K5�	�@b_�E�i�%�����D�,,���&�� TI �&PџX�sdD+,dQ�&
@A�A�&��b�ltX��}�xyC@�E9x����b}�Q��JV	h�S$	�8,:���',Ѫ�@�1�t͑C�j1�Q����
LH�Pg M'>�f �/��(�!��N�q�&�*�c\�Q�M�b�<+p��g�b���1/�T?����y�-����};#��t�I�#@Ƹ�y��ő;w�|I�.�)3��[����M;v�^�o�֤:aN�p=� ƄOO��PA�:FҨ�Ӧ_]؞�zG�X:U����7I|��)E�I�r�8�ض��u�dE;"OR�"R&<��	2&́Z7p c��P�[��3�j1F�>�	@$�3$�TڧME(�,da�l1D����	N�3�@.�<�\sB!ºX�8�1�Rd���^�*���F&�8�xI�q�Z��!��Y�#Ü��D�Q���"�GR:�:6ę������	�3�,���O=�%���Mz:���JJ���_�v|{F�Êr��T9�CCbp��O�P��p���S��e�e�٫l:�����╂D�-XU~ز�a��`�ȓy?�DSFܖZ�Z�*X�p���N�$�[�&ژ ,���)��q��@� �U��?0�x| �㏡^��!�ȓ�bE�k��LQ0g��*���ȓr��0�GB&58�¬��%��S�? cT'�J��X�'C��E#"OR�j�CY&rp|�6����B� �"O���RmK�L�\����'M9�8z�"Obء%`�}��ga��pQ�"O�����09���!swu�"O�yy���JЈ�;D*L=	L�w"O�A���o%�H��+߅l(ԣ�"OJi���m�hd�>�}S�"O4���I�(�DL8�O�.Фݳ@"O8h��N]�0$�16`��|�PU"O|�Ā 7"�iKD�Ć+�Ny�'"O� ��<Y��}aqc�+L�⭩�"O�BǠ�h��1Z��ˈY$:�i1"O}��%�Պt� �,}f�YB"Obe��1\�,)�l��n�⨰"O��jg�R�IZ%���8�f��"O�٨�E Ȝ}y��zR���"O(�@�6b�д���pR�y"O�i�j�X|bF`ե@�0�y@"O`�&��/P&��SM��(m*A��"O�ERí��N��p�0f��N^����"Oڡ���6���'��7d�q"OA�'JI�ڌ��Z�<+<�y�"O�0j���I�vP��,t�,p�"OpZ�%��SW9!�_�JdVyA�"OpYFG�7jhN�j��		8~��B�"O��&FY�,<�qY5��53���0�"O�t�ġ��H̬U:t�W(�r	+�"O L�jA1s�ţa�(�΍��"OV�؅!\�HN08�CQ����V"O�Ăs��r��2 	���891"On����2;� y��K�>[��g"O(	B�K!a�fi���#j�Tx0"O2 J&l���֐�DO7yc`��"O�|���,X'�TX��+.���"O��S&��k�6��0ߝq(�� "Opx���V"'jM��O}"����"O2Ac����#l�P�֥}���8�"O4L����A�b��6a 8�*���"O0`C�U~�]2 ��4���""O��S�蜉&�J��4	ɷa�V�e"OZDH��E�3SިC�*�t� I(�"O�A�pE��w�&�b$I�3����"O���ݾG:��[�iF"z�n�xT"O� ��A�F���� �Fq��"O���F:��Tա8_��!"OR$���ťx����d�:���"O��a��d���z ����1�"O|�1FP�_b�zģG�g`�9�U��[��3>}R<A�ő~j�!�.�Ph��������Y#n(�D�ȓ.��&ۍR�����_+�)�ȓy�� �Wi
dmy�l��A�p�ȓr����Z�GA��Xb�û!ÊՆȓ>u��H�B5=���p�\�;N���0�Mb����[n�P�L�8B�N ��5�бQ@m��c��eAR�¬�ȓ:�F i��[�r���ڒ ӿQ��`�ȓ;jHiB �\>S��pRfl_�@�z8��vR`��W:��ꦪ�11��9��j� !d#P꽙��ԫ��Ԇ�OyP]���B�U\l)x�ʋ�7�t��ȓcN�Ae'#h�Xͣ�ߝ7��X��U�<8��ĸ1�б�琴5����ȓ^=��g��:>vUIv:):���S�? �y0�l�
l\}��d�����"O�$��#�_�D�X� ��o��C "O���d�>A�4��L���Ⴃ"O��X��Ȓ����MWy��I�"O��c`BF�/�6�C�,N�B��(7"Of�[(��\�����T3�ă�"O�01�J�����S���"Oq@�51�sAL��+x��"O�Ȓ!qi������O�֐�p"OV�B��#dr���Q<[���A�"O���Ӌ*o��Z��A-Ra�h0"O����K^�s@���?'w#A"O��IڣD5"踖BR)=ϒ��D"O�| ���ZO ��V'_Pĩ�7"O$��ɉ!bJʐ��ŝM^`�*c"O�u�掅$VŐ��F��ʅ"O�hp����y{�������u**da�"O�1����(t��5���\|�"ODC�*P>�~I2"��K��E:"OʤQ� �c׈XY�j޲'���kT"O\!h�J]L6]J�)�#w��)9�"O�|3�*�c��"�">/m���"Op}�bi\���UƠ�i�"O��K'���C��6m�@�"O&��s��@$��c&�ٖ�`JQ"O8+$���YHv(�!����ؓ"Oތ�F/U2@�J��tcϗ~$Mk�"Oظ	�]����b�Ѐ;J��3F"O(a��M��yv�_�2g��b�"O���7g�69��d���ԝTdp�+ "O��J�D�K(���CkT_E�$�P"ODQɣ��-3��{
��
�5�"O�!���A�zQT������?�\�0"O��w�_�?.<m���\Td�b"O~��C�D�"�����^��B�b"Oz]���kFb����$9��4"O�s�'5x@a󂥘�s+&�"&"O��(����D�T��dB،n�4�%"O,)�vaOHZ���CB��:� �"O0ĩE̓�I���c�=j� (Bg"O�T�6#ެz�4��L�9�|�J6"O�eC��4 ]���+w���3"O�1��D�-�$��5`?[Ui�"O8��-G�r}cs-�$��"OJ�f
� �L�(�ՠ�8�(T"O"�h� �n�NT*���/��,�P"O$�3 U(6S�Ar�Ė,��1 "O�@Y��Z0j�\�X�$g��0�"OĔ���M�%&bY��ڧfZ�!�"O��X���.u(,@� #K�a:b"O�E�`4T=XP8�?.*�q�"O�XY0�ӦaДr�Ò�JT�W"O�Q#ahS/(RzXb�E��TYF"O���˃:��`�`Btcb"O
}A�� n�ܰ��ʃ�.���"Ov)�5 BO�5�R ;t�P"O�J5ɞ�'����.ٜ8k��x"O��J�� +����.u8��c"O�9k �2N�Պ�a�RW��F"O�5P��P�MZT����N4�Qp"O�:�(%'t% �@����"Oʍ{@�L�
 }*@�J&f���"O"xP���Io����ϞL��y�"O�pp�92��Y��Ǿ�
��V"O� ��"��/r#�Q`6���d�@�KQ"O��{�ϔ|%J媧�P�ymei�"OȅK����S���Klj��"O�u���B{W�DP���4l:t@�"O$���&G�b�y���`��"R"O�Th��\�`��|s�b��1Z=ر"O��T�)�TŨ�[,d�Q�"O�+'��]�!�Se�0����"O�d����r��]�f
�?Ld�a"O�X8���"Z�V	S����0�"Of!��*;�1t�Q�z�,9��"O�d:��
6�y���ϳJ�����"O`�2uN	�&k�j�	��9zs"O�\k�b��"��� ���!"Oxt�EI9z�6��؎2��u*S"O��X1g�i�r��4a�0}QS"O��I�+@�c|�mX�� vvT�@"O���WF3F|��n	�p(	�"O�M���D ���V��bSpu�c"OvH�AЗyX�;�c�2���"OjHxg�&�� %��n.��3C"O~	��K¨g�1%M�1X K�"O��aN�8�dp���#.4�"O��D�&i���+rD�=e+h�S&"O*�'�;��j���(T2NQؗ�'��'�4u ��H�(<ja���~p	�'zB8�pjA��A�g�Q�$p�'�b]�Wc��4ѷ��PIf8[�':.�f@��H�V�;�d �HL��B�ay�惊kv^�+�a$'h�ȓl���ro:B�|�c���;$�D0�ȓD�P�����dj�Q��b��M�x��^5z��F+)k�tY��k��20� ��=S^]�qމFԋUa%�H��ȓyT(�!V�&w�̋��#�xć�@�4�bU$L?�����n�����x��'�6yG��[��\�VӌKQ:�h	�'�,h�gȣU%��Q���mF�$��'�t$�7�Ԥs�*9(���e��$��'wtay�I9w8��.�HA�'���/Ң:9ƌr����-�B����Dq����C�8�����6[J� D�3 �!�d�*]������X�\��@��6�)��=����N�8��_S��"#�!D�t����`�ġsa�a���#�����ziΜy�&�;z^�@h !^;{�
m��r�  x��>�^�`a��#9���ʓ}��(IEI
���5P4&��q�|B�ɍW �腵U��9
H�.D�zB��!q�D�g(�$~��Uk7G¿`�:C��<����RG�,�R�Q&6'K�B�VM���
)j&
�0-�8$rC䉘XFZ\y�c[�C�:e(޼g���ȓ�<�b�ȷ?(�1� �Tt���G�t|ai>�1:��W�+-�<�ȓ�hʰb�m�R�������5��?T�zrk 2���ƍ�=)�]�ȓ$&��a I^-t"��w#>\��r���Sn[(zxq�b�TK�V���F��<��ɉ*:V!Ѳ�Cc)�@����%K6d�/����vͅl�29�ȓ5��c� GTU�Ŏ��]��9��Z��Ed
ITU#f�ȓ��$9q�Q�_o���I2���S�? ����)D�H����<��s�"O�HVAǼΆ$b�	�<I*���"O�	G�M�TՆ�(=��:f"O��8B��$/w6\P�D�=~9�$"O�+�8nW����bտ"p�Q"On���-��W�q1Q��4��q�b"O�� *���qe�6��Q"O�X[@����ic� l��M@R"O��"�j�=IA�2eͺn�.�XT"O��ؒg�P<i� Cѐu���G"O��!�ʆ	E�HJ�!��U�`�6"ON�0D�&��9`���~��U�#"O�8���M:y�6�g`��n<3�"O��P�K�ͰL��/\�?19a"O���F��-_��P0�7hj9*"O|�+��$^UL!�D�Q53��H�"O����Z�$+LıW�][���"O�P� 7B:a��/ V��(r�"O$��a�n�8a�����Kn����"O�� %n�W��������m��"O�,ɢj���=IE��˪��S"O�(���©r2�e�]a�"O��ٵ��>�t�����.)�8�*!"O�� LB! �B�;�E�Q�R�"ON@���;YB\��b� V�h��r"O4�0m�ZK��hT��w�����"O�h���{��� �*˴-Nh��p"O�-�O�(��@��.l���v"O�,yCN�V@�H�g���9ΨQ�"O���&�֐��y��fC#�t��"O�J2%5�.� Pe[,�� "OHD9�B�(;H��ƭW���8:�"OV�h$IO?|�Ĕ��Jڸ^��t $"O�5��W/ET���(]R4m[$"O�a��Ԕ&�V�XW��A:nmA&"O�T�-��C�US�`Ϋ<����"O�Ű�*�a�����קF|A��"O�����
�(r�V�3��(w"Obx��J�O�81���~7��[E"Ox�S1G��J��Ƀh�l|��"Oh@�bZ�x���̏h]�9cd"O�\��kĥ~��WkC6`�pق"O�sE�"'?�%�f�ˉe%����"Oĭp�霝A��-����6 "Od�9�H�0:�,�H��k�<�!�d�uTD�j�坊�[r��a%!򄓖J���:ɶ)Dk��+ !�ئ5��*$58�Ƚ���	m�!�dJ q��uZ��_�t� }8w��Q!�$�6Ǩ�1�&����|P��ϫqC!��A>�2U�b [	o�F z.ڭ�!�(D�Rt��a����S�80!��>A.� u'��.�v9�яR06,!�dU�Hg h  �   n   Ĵ���	��Z�Zv�J�(ʜ�cd�<������qe�H�4��S66<��ʄxG�f�َ%� �8�MαmF���򄒻�7����۴ub��=�	Xy�dݰ|N6��#f�%~rN �E^+Wa�:��]9ap	�=���3�l�&6�	o6MhP ��=�r	���G1���Æ��C읏8A�		9�[�H�y�If������`kP��%m�<&���ťR�Y��MN-c�0E��$S��Lj%˱?�I�'�X�06*S�!RHHh�A'$-�$��O1��2r��By��G�FO,�0Fk�O��ϓ&}�|�E���y"�ƭR�#���;>+�!2A �"�~"h0�N����	��I6�ꄹ���5Jv�g\�a�DW��۶O����K&�\�b�H�iu�;�X[�h�a�͊c%���Ϗ�[��y ����O�����^����
^n��U�
�~L>;B�!L��'�f#<Y�D �I�h<ٓ"�� �`i�g�߹�6M���O\���D��
a&%�1 e���RD�ڈ\J`�s����O�!�O���T�	+`�p&��X�����^�����I=vO�O`�E2�.ɰ �I~�U��6�O��;��DI0�?yC�\==���RRHKS�TkDP̓zS#<�T�5��O 4P���\_�A��뛳-�d8�Oʭ�H<��-Z�MK�G��H5�d c�S-pi�ԚG��ßp{�u��
��S��?�2�>���~��d �j/�X��O�UL,�q�d�?�OJ H�x˵˞9���5���*	��μ>ѱ`9}:�#<9���;9�+��ʴw�e)Eȑw�<�qN� 2  ��*�Of��e@�&+�1sN�9U��)��'�� 3w^�yվ�+�h�O�U�#�(-���v�C"�H��"O��S�Vu�tx�e������P�|b���NA��Tm�xun�}�6��_z�{��ѥw|B��@m�J�<�p��D䘲�
�� *V��X*KzIpI�	;.�6M�*W�BI��L>)�f��.6
1tDD����E(<I���5r�Qf�M1(xY�A$���X'O�<�V�������z
� ������9�q%3��I��'�@�b��Q�ka��]
&`�l�҆"M�$:��N�{��������yB�3hv�!s�o����0�����*_Rp3�i�C�y`�$�>EQ-`�D��ț�Iq(9�!?D��QPїo�6�sVcԫwa�岅�9E�|�2`'���&��60<&?�xI>���eC0�"��3�~D{� J�������v��-RB!I�QJH�D��;� jCB�e�������T˴��\>���łvi\-Sl@�#��G�G�;T�ڤs�l\�A��!����h~:�y7I�f��xH��=IvD�34��:Ө]����N6[e$���͢<iBb�zYl���K8�5h�����?š��uZP���-�2Iw��Z!g4D�H�����kV��+Bpx�7���!8� �柞&E�vM.oyfU&?QaH>�Ү$�F��7�[�q�P�b�jI����֦�!��@�_>H���, � ��Y L4�tr�+��!8Ʉ�(>�f�xC��s��I$gDI����;2��)��^y��I�rH�3�	�/V�k��6%�5���2�"O`P���w���L�4Vy�%*����d?�!"	#4�(Q��b�O�i��`�B��A���	�"ܬ8��'N�3�E���؃f�_� 2l{R�D�ys^�8�C�]y��9�g}��Qܴ!�`�A�Q�1;�`ȯ�y��S0.��y`��X�M!���M��5p�����\؞���"�W����"P�[+����H+\O��
P�ƪ(+z5�&�'��8��!��3�����+Z�i*�' ���wΕ!�n͊�L�B-H�}��������/�[G���An���SH� D��<��p(��S�(Q�+\��N&b갠��u�'j��E�,O.�ô-��q�:�X�N�6nP�"Oy��_0:WZ Tp���]ßp�G�l������#�p��^0{�vI��m=D��&aQ/.��Вc_�+���z�d(D��B�]�,�j�Y�B=�)�-:D�ܩ���N���HK�i���q4�<D�`��	;��}s� r��P2�;D�P�5�_#c�컇 σ>�����;D�`8�<^ ̩���RC�T�e�8D���u���aD<Jdʖv���YE'D� A�N�h.�F�._aZ�S�f$D�� Q�ׯŨt�R+'�Q>D�0�¬�h����!��r	'D�����I�,���Ǐ�L�4� D�<�T�E>9:0(q��P�0�ԝ��.D�ɥo:X�u:�c6T_�R&,D����n�3.F���A6Y����G)D�xk�K�>�V @V�4}����*D�@�G�G����R5<5b��<D��B(ױD��)s6��1[Z^%J� D�\�d��,� y��-�Q�q��O#D�k�b�=&����'��g�RL�D?D�����J?}�:؁�B�=ju�I'D��-�S��]Xf�0"�A%D�p��a�k)���͛-%��%�)7D�hc��ȐG��A���&'�3�3D��SlI 7��J'�	�� !b��0D�\��2�u��\�k��q��'��4� k�6�<�F��l[����'$��S0�FRlqq6AO.7	:0	�'�`m�㍎�
����Z�4jm�	�']�)�!F�;������2��Dc
�'����#�S�7�h���+[�	�'��!�E��$�H�" e����U��'I�a!w�	3�8,�*�T��A�'Az��5�ˈ/� ��t�>&<�
�'���!���aMz%����"��+
�'r�"�N
�-)�ԩ��Ñk��:��� �EkU�3A��e���L�;���a"O^h�Gf�5.ڜ����"�A"O�X5,����e�b�D�l�Ω��"O���G�cfj0�L؞(��\�2"O��"g��g�`Ӂ��r�<�)�"O"%� ���S/f�s�IBy��ᢢ"Oz�C��l�N�p��l�P���"Or$��D�-ZԥS�-� ��<2�"O�4i!�<�ty�0�Q�/����"O�QyF�؟}�r!�%k�7KR�r"O�\�����@A
��|0�#"O���T�_G�X۰�֕Q���r"ODE�&Ŝ=�`��B�1E�lu��"OX�pQ�|z^�Џ@�s�,���"OA+D��+)$%Jg��>�����"O�ݱ`�
,�\��6���tq��"Oz���}�T���l�S���4"O��ƌ^�:���@<�@���"Oz=+q)�vMX�5�@(�D *&"O|��3��z��bJ�Ӻ�� �	�9@���!�0�ԩ~�6�O�,[�t���GL����Z�O�!�$X�(���G��:J
��	ݽ#�!��ƩD�Zdxa���tfT����@9!��-C>AX��� l�PHaՃ�^-!򤘠'�h�WM��|�e��cװ*5!򄞺%��A�D	'z(�z4�%*'!��s�,㧫�2!ǊL��o1!�DF<E���O*y�"\h�-Y�,�!���:CӾt����`�L��7�D��!�$h异�*e�V�R��$��=�ȓH]�aBB� )t��Yj��'�5��}㔅*A�&7���!F�R N[^���ii��AΈ��ޅс���w��X�ȓcC��ꀋ\�V�!)Ё��s��M��	S0H�&1���r%�������4�2+ۭ)ڀ4a���o<�(�ȓbYDA:C	X�#��(��b��U��9��G�ȳ`V�~��M��S�t�y�ȓ.�1&�^�4i�g��q=1�ȓo��MPG�	@�
h��]�쑄�ʒ�Ѓ:W�]ДE	 /H�ȓe6$%��D�*1s����#d�ɇ��J�V�$ ��JF�8b{�n�9p���2ʎ�J�k��'Ț���jI���#�b6%'B�ȓj!����'V�J����U�Hs��ȓ$��e���[�h|��B�>\�(��7��Ec�g@�aƔ���J
"��a��]@����d����pW�Ý�����c�x�[��U���*k�>4�\��Sq����LI�f(��ʑ�C9c2`��VM$]Ar�K�A�tZ2�+F���b�\�@$���"��& 
gݦ�ȓV<v�x��]p��Qb���ȓ	�-����K�Р��I�)��8���bO�l߶<�u$��md�ȓAhΘ����4s���Ň�Q'�!�ȓ(t\�8e�ڑ>o@��+2<L�l��[x�A��D�L�mӣ��豆ȓ��� t,��zf������̅�C�9�FfK	�����|0%��u	a��m/|%�q�0P�̅���$���J�`Ĥ}`&l'��T�ȓ/R��1!'I�Ah]X��>���S�? �	��ڊ��a���*I�T+�"Od8�M�����`��H�]�F"Of��0��n��U9�7���(�"O��1�ύ H��{��խ(�`aR`"OH�{�E�N�{�l`��"O����������ͅ/+�(q��"O��g%���j�eW"J�^��r"O��rC�h�dP���`�8�6"O��r���:�RH	-����pq�"O|Yh�BFK"|��"�ӄg��t��"O>��D�tx~Yٴ��R{�	�"O.��CE��,�u�a̓�qg� 
�"O�c�ϑ�@��]JDL�qKn� "O����!9[�eb`
H�7�� q"O�LRd'BT8QZ��	n��V"O��zWJ�|V��*�.-^����"O��7�ñGq�����Y�H�Q"O�� D�<' ���o�)|��t��"OM(T\ xL�1!t���,�vmQ"O��S�&��4jb� 5}���3�"OX]"�坺AO���gܐB���:�"O0q#��ɂ_����� _�����"O$���B���|���h�|H�"O�A��`͸;=�2�ł�<Y�iC�"O�� �,N�,���d� )J��5"O��C!ȳLw���d��g���#"O(�9֮Th���@��:|i�"Of����z_�)s�*��̱�"O���P�h肩�A�ʾ$�H��"Ob�Y��M�Q���2�H�?�6U��"O��z��ei�p�,�*}¼�ȡ"O��"���3��
�Y]҄Yp"O��)��E��(��L���\6"O@A���� y(А1�ŹG�z9""Ot���%�/��+�h��p�Z,6"O��8Ҍ�rN�(�
�>s���"On��'˅
���`5�P�����"O�;R	�2�1#�A�F�^8!A"O�B "��P��Ћ~H��@"OXus�J�}�<K3�	[񈰻�"O�d9���u�B�`�+#!���k$"OМ�@�(���K��
�܅3#"O��S"� a愒UKՆN����"O��c�k�f
�]�pJֱ,���b�"O^A�`�J��=Fd�(�<k""O�aD����@�^�@|p��"OBq5 ّnt���Kߥtq�iy�"O�2io�� ͒=�mbâ]!�y2�ɍa} Ф33`��j��>�yBɇ.M>x2��H7�P9`�eӼ�yB%H�Lc�`�����3��� ��y��A��Pq�%���4L�;ǈ���y2�Lx�I`�ceʰ2����y�
%,	�I37�×o=�A��&�yr`�"~�*1'Q�b�(��JK��y�.�Z>
����T�D�r9�S��yB�9�<��^�7���tΆ�y�$�1D{,�	/�43�)*&�'�y��	#.��5d�A��;n?�yR-�!���AuHZH'�`�B�
�yB�k$i�0�V�DD@3"˖�y"�'���kT��Nkڀ��4!�$X2	�'j.M��]��������'�����U
�(�h�LO��X����� ����V겡ᲁ�jnt"O^����S���IB��x"OT( ��d[��@Bf�&$��"ObA��ل��b%*T`���"O��l�NdR �2FM<*xr���"OvY���5c8���T�q�,y��"OL$%�|"u�!߳���s6S�F{����.G<r�8��B+m���%`α4!������I6 X�a�Ԯ�0k!!�N�>{e�PMؾz	,�Vn��~.!�G�>jƩ
�j�9���:p!�$�tԜu��c�2Mr2��4MQ�o`!�D��-D���KXI���m҃TU!���3#Y$z	ٴ�R�"6�_�=!�^)V��ɲV��#=�	sk�b!�"�@�Rc!�TFȠ�1ʚ�!�>%��" ��1�Hl�2�'��A;�IM�j���Pc�̖8��A@	�'�T��fٰ	n��>18J�3�'I�4C%Q(}�>�k��-W����']�Xը6W�d��W�M�	�'�Ƒ�J��)y���.�����'��!cO�A��$PE \8 ����{�� ZXI�P(��B��y���(~a��1�
S�L&���@���yr��8;f�#�Q�Dh.q� �^��yR��t���[ ʣi����4R�'�P����Q,2v=
�՗i�����'������X���BǩБqS���'�H�5��*V��p`�[lĪ�'�p4I4��.$%��K���V��T�<��	:�(0	�C�02��i �m�<���A�/����ņ��f;(-����E�<���_ �
�iaiY(#�UJ�
B�<�p��<W�(��`O�!���y�B�@�<�0]S�4���ؚ4�n䩒D�H�<Qs��,8Մ!�@�G ����Y�<A�f�FM�w-�:ך��"S�<IU�ӦZ�T$�Ō��L3����M�<��A��v��Ek!��&�5q3(E�<��ׁ0��	���e�4����C�<q5Ϙx_��w���3��hf�<����:*����`Ez2q�&A�E�<�2N�/p���t�F�Jp��[�@�<��եb�Xd᳧��H��;�)`�<��M�����U BSȊ�r�k�v�<��HK1����� s�"�� Z�<I�ρ�i�h����8c����gT�<b�J F�>�� 	�LX�At�<Ƀ�хpR)B�"F�J�)	�cLr�<I��4�-@b�	��yр�Bv�<��n�����F,B.d��Gv�<�Cnٔ7~�`j�`�%_�<�!0�p�<�ҍ^:r��V�$=�:����n�<i֋E YT¡��J	 �2ك�jf�<��<t�8:�+N���1�%�^�<a��w�`�I��,te��Lq�<�BK�򬽒s+ͤs�N��o�<Q����t�g��2h�]����l�<�rГ7=āZN��.AF�Q�h�<aF�X��$@R��F�D�i�n�h�<A�eS9%Ld���:VH�"��Y�<)�(= �t�"#�p���g�W�<��DCI0aH�!ͺ(��Z�o�Q�<� ��T��$j�hs�+ܒ1�"� �"Oq��*
6S@��R+�!"��6"Oh\x�U3����O�e�4��"Od1�#.Oe!P�ȋ"kX$��"Od"�J�J���!��~�a"OX�S`��1��DJSE��p���"O*p8��P�#-����ۢ6���0"O�� Fj�;���y�-E�x�����"O�]BP��1N�ƌ�	~���"OV񻐄�P4X���@a"� 	�'rȡ�J��ls��4�B�"�̊�'9R��;Pv�ySbS��N�`�'p D�D����y*#ʇ�P<��'u.:��L&},f(���@1"ۊ�
�'�xd��KJ(.��1�0G\��	�'�2�9�Iʙ=�.!���%J˂�a
�'��� k�k#~pg,��v�`
�'Sr�UfE�k.�CFK�tx t�
�'�fdhc>du8�0��ǖW):���'
�aHV)HIA�;SHH�����'>�#�%�-B��`�ץ<S��ʓAzThz!JC�$> %1`LϞ�ȓZ�����%�`���ź%���D;8��ꐝ.��)W�?]�r9�ȓy�t� � @�?   j   Ĵ���	��Z�tI
)ʜ�cd�<��k٥���qe�H�4��6]22<i�ʄI}�F�>A�,]��#��r��A�7-�M+3'��y"���<!�BA=&鸜:W�&��P�3H۔e��[�A�)r�������Z�FÆ z���r��*�4܁%�7��$\
46v�# EJ>��Չ'�� $ߓ��
�7T>�z�e�#`&��[��ׄ
-�#����/�'g�8�5�ZXP���U-ѯy�H���ގ` ���=��A-O�!�ɒy���H&ƾ��A�'�`%���~EJSh$$1�OX%N*��`�%�~�+��YM���RG���D�	k��b��
�}d�+�ՠǙfR6� �1K(\=
��B���(x�e&G��h���D���d.7cN�K�cM�O�����Ċ1��Ć�#,� ��!`{��"*4{�<�#<I��'�	�/���f ��9�#F(Q�X��7-^�O@ų��d(�Xh��F�.\@�)� ś�v0X�Ĝ�O��K�O�) �ϔ/c�l���K��8�r�W�p*C�	(N��Oj�aj�2-�����Rr��I��Cٞ�O�)#���ɰ�?�I��L(��$x"TB`t�[x�#<�c�0�$�
�����,F�r��K�)łl���ʵ�O^PAI<�G"G⟰�GN�1X���T%<#)����O�t:O��kRO�ܟL����M��SQ?�2��ec�G�v�p�P �G�]g�2�I
�ċ��>IRa�m�L�@C، �v��D^}"oBx�'E�Gx�e�i�-�W`ԕ�}#Ei"�y"�Um d  �y"�ݬ:&MS�b�87�D�CI���y"J��q �4
I�M�R�-�y���_^�H�/Z�'"q�g��'�y�o�"f�´HU�Ң.�537�P�yr�;���H�G$	�Å��y2 ҋB�8�����&f�����ybX?y�v��呄�8����y�O6eL�!�"�~BP:�Kέ�y��z������ds�͈�y���Bt,��a��`���@��R��y�k̢Kh��C��3X��#�+��yBlE�_q�X�+�
K\I")� �y��N�[�^@��G�1DFMB�o�2�y2HD'`��<{�dҷ,�B��2�T�y2W�]u6�с$�#�]�0� �y�WD>HɣG�ϴ����yNE;Nv��C�
�
�RC�V��yBF�� �LzdF�W��B��yB-��[� ����|�D9jҋ�y�O+p3�42C^� q*q�R!�yr��j���a�2X��p �4�y"O+��@b!�0��(�����y���<Ѥq �F_9i�&$��e���y"k j��l)f�Fc��MC�K�-�y��&P򩺴gH%[��YA�j�y2EǚInQzᩝgB^t�6Ɣ�y�gJ�F��ьv�f`��]��yre��F�H�"ŤM'$�NYҵ�@��y�B�8I�<����Fi�5�G#�y�i׹I8,%#qC���d:%	�y��F9K� -j%$�fd�!ʺ�y
� �x�k��E^&{p@�=F(�X'"O>�#�h�JC����)
zh�|��"O�,+o[�D��Ѹ�.Q;ZSZ�[p"O�|�O�1A�� �홨L?���%"O^�!�-�y]� Aި%���+1"O8�8t���su�Հ"�Q�j�pV"O�(�p�݋�sd�X@�$%8�"O$	;E�()4̤	��@8��P�"O��*�1��Q����Tn�X*G"O"�[��ԛz��y`N!J�%��"OFt[B֊~ܸ�A!�#���"On���]4s�ASB	W�\�18c"O�iV'�
^�ܸ���O�t��"Or�ɴn����51D.��AFu��"Of	9Ń]�2l�X�Ы�!W@$��"O��z�nU�YKl��o�kT�:G"O0�u�ƛd�Va�4��?d���"Oҙ��G¤_U���nPQ��s�"O,�9�B\;~i���.ŎW5���"O&�IW��:����L�0F.��:f"O0�"�(�'|�E���P�0�g"O�!�3*Y T+*�  ��7n��Tb�"O͡p�9%�\9�>(P�3�\|�<���J�"���kW�ԅ)�te��ds�<�uc[# *  �   M   Ĵ���	��Z cwIJ(ʜ�cd�<��k٥���qe�H�4��6_?><y�ʄd�V�k�,h"�l�A���օ�0267���հش=�D8�IBy2 ��E�@F�4mBԁ@�ϻU�,u���:$c �=�G�"�o�6�"eZ�p��7O�|�	3��
;2���<&f�J$a؏U�Ɂk*���Ȏ;q�I U Bd����:~�(��(�,{� .��O|p$)
�=��'�D��*ʟ?#�PȓNUoO���$DlPN�o�Z��ΓC���͡<q�O�e�P˩('ąm��6$>ax��L���p,O��*��J�)7�jC�䙲��Y�y!_3"���Ƈ,5PVN��yb"�w�'�L8Fx"c�J����f�q����w����#<�)T���%sp�����T2����&�W��O�)ێ��J���'�L��I�=f࢙R3#���:ͩ�461�"<���9�@�&9;��Ȕft��CV<�����O�H�� "<A!?A�͝] ��pON6$��s2�Ly�B�'����?9���JU�tȃ\��~t����2ܒ"<��a$�L4���H1*
�i��G�9kp��l\= �1O��	����1�ē:,�"vɉd
�yY� �%G, ��4NJ#<ف&6�[?Q�L��v<�k��o�z��%���\��P�l��O*Րg)"��'H*ם�f��`eύ$�R��Ʈp8��=	W�(�S��'�$�ޟ�B�kB���<���O �Ȋ�� �O����
��~�z0j�	Z�iR"O0�p�  �x�"OfY��IE1{�%���L.P]Z7"O�Y�D�1 ���)e��H��"On@S���9Y���s�ıS��T�#"O�$Ѐ#�Հs�a�Y[�ъ6"O�d��J�:�I1�E�$fИ w"O�)�9R�� pХ�\�հ�"OHu{�̓Dm�1h�d
<q�z�{�"OLx��Eƾ( ��uW���qȒ"O�8�"��V�9�2k� 3�ڑ�D"O��xs�Պ ��0Ѣ��/�u!w"O�D������� E�5F6x�'"O�1��/V�F8��Q3E	 "���S"O�li6�z0n� �_�N�P}�"O�QP��s��k����	�4�y#"O���c��0=v"�'�+���X�"O��ۦi6��yXtf��l�h�(�"O0�AE�(X2�9�c�D�.����"O
�X��Z�h�xQ�)*�����"O�}rd`S�tC19F�5uk���	�'<6�c���#�XI�@]	E�| [�'��Ĩ�� >1��bc�+,lII��}�65���1)���
���x�D�1�x���K�Q��(��|iL���E�'%��a����$p!�}��{�Z�@�J�8GR`����#����ȓ^ځ@��<����R	�Z��ȓ2�J�x�d�[m 0�M��M���v�����L@�+�b�{�Hs�⑄�N]�99��K|���g�ѱc�*���AfLZ���4�*Y���Js�@�ȓV�b|9���>3��c��+�D�ȓ8{�I�D���:
��` ����nC�O]�H��jR*�>G�B8��[ݬ��JB�8!���Jӌ��L����ٕ~�lHI�g��gl�%�ȓ	�^���)"�>P��I�TI�T��*�4{���1���iE-SL�&��ȓnf��jWdǠ<��v���ڝ��y���v@�H�̩��f�yҲ���^�5��.�!����з=����Dr��bR�Y������0��ȓL~zP�g� ����Q�܅3�>e�ȓ&"���oH�w�L�R�SC6Y�ȓS-$�K�ʈ�x�P<�3 \ �"���f�`T(�� tX����"�h=����k��EAd)E�m#"퍟D8���!̪d��<Ԯ�btGA�Mآ�ȓ!���Pe&���f/¬	�"h�ȓz��iҡI[���Y�͒#e�Դ���R��ī=;VX��oWH�@l�ȓ.�|i�2o��R���a�&97�хȓq��з	7_�u9;Et���'���wnƕ����V1B@�ȓc�8Eǘ�<N�� �$ձ\�~8��L)�I��)�f4�ɐ��*|l��ȓf<�mԤH
da�p�j�t�&)��� S�LEB��'�8�L �-�
4���� %J��X�'�\��¦�v�:ɬ�'q�Hs�.�4���[e"��H�(���� ,�� y*zX �"O� \m2�-�5��\�Aˍp��Ȼ �U��,�a3*H���)��<��*�?`�����W �6��l�E�<!�͊6 �t�� ��.��)�����<yC�M�Dy�­=\O�����9�
�`vm�y��	��'�����O;3�ra�E YjN��'�K�f�^0��y�"@�lQXt���T���`�!�4�O8��f℃\Ӭ����)�3d��c
�w��Hq! ҠZ!��77L��r�8k3�I� �*X <@�C՚*�`��N�"~Γ^
T�
�W/7:��yqJ�i�Q��9������Ϙ ThY�p t��I�y|��i�'B��$��F����
�J��ez���a|��
#Ḑ�e�ӣD�d��k�d�5	�F2p�a��'׮���AQ�W��-��������䟁?��u������(�8PI�Z7 �h g�]�>m(q9"O2h*B�\�^��m0F��7o�@Г& �Ĺ�uH^���)��<�Q O/OK���8*����\p�<�B�Sx}� ��]l��t����l?�3`E�-��h�e���G�EU��� Wb����	��"1��'��r��>FP"��'��P�<��'�l���%�	N��Cw�I*���'��mV�B8'����JJ?���S	�'�d�"J�"h���8V癈Bh��'�~(�����<�P�됞w+bɲ���^;�>9(��W����S��0d�]�oK�!�$��P_x�T]�d��!�n2p�]��A'O���hQF�S�R('��O����6Kv��(.�~��7"OD�8�P��%��x H���@@��9�s��Y[JT�'�T/{��I�^�Ԉ��;M�� "pD�8l�
��d��E��9�m (���Q�F��"O��`c��)c�Ԥ�sB�`���'�ea��JSB���AMGG�ȓ�}��2 ���K�e��( D���79�O��b3�_��$�k��D�2Vz͙	�'�L�
�͂0Jz�p��@�(^��ao�+�<(�$癀�A�����7
�,�I.�\�șw��К���P+Rh�Ј5q�X	�']�L��;�7��i�����!ʗK3N�p§<D'�u��-L�T�d��'~2�k$�ݗ��	=l���Sႆ$"�KfD��4�4��d��9s2���}��!�L�$S� �i��%����T�\�1Кt ��H��B�J�K�I��q
�'�M��`\��� .� |���B�y2N��~�����7h�4��h�-��wȏ)7�e��[�I�a�$O��CBڇ#�Y��'/���P!�z�b���J*�0R��Έ�T�'O~�ҙ�AB�#-�����|�l���j�(� z�w����5F�h}� �G�ۡ�i	�'����Ռɍc��X"w�Y~��e����Q�0��H&t��e��j�_x��H�,�a��pz�
�y��M��O$��%HBaJ��׌Ϝp�D�	�v�<1��]�\;rAS�B���%C�+'H1I£�.C���b�ه^4�͂"�$>��bĬ�+S֔u��	�;�6|b�˔1n"ɚ�����RjȘل+וO
�eKpi��L�r���J�nu������� �ѱH�y[c���N��AcJ�sH��'�� c�؏wZ"�&#���s��06Z�� w�D�@mօA"�9��(+EtP:�Ɲ% �䑛wo�U�A�'X-(���V0$�~�K��5j�}���C; ��q�РxP`1R�M�^�$�c�A�@�1��E�"6����O�r�(Ѿ,��'��)��Y*6�����[�:��э��d��2s�O�iC�hj�DV+pB |{
V�t��4��2;�:æ��6v�b˓>���`,;,O��[��LUߊ=9!�E,����V�t���W��+�nK�#��1��ն`LL�>i��'�M^�0���i��(D���Ñ\��	1��t�M;�-�H7�������s'N5 �l����c7�>���I�F*B+�? ��K�*P<�3$]�|���H!� "ZM ��UJ�<T����w�^	W 4�����X���۰<�D(�2zz���g��n#s!�J8����j��x�2h�L�A)8���@-?���`5B��7�е� �"O�5�6
Ͻr��m �B��$� �Ap��S�I��h n��Py�#}�k `t ��������
B�<	D �8i��xK�i��;��ġíѡE���v+w��b�����H���G3�Y$F;Yy!��H���j ��n'���f�F�W��	���,���Vb)|Oi�DꄖVy�\��3a[�j�'n�2�ٕ �V)��i����NS�R�~dpG�(�6��	��� "�zv!���Ԉ"�O�rU41����)�Tҷ�Ա�h"}���0@|��70x�y�@Q�<A�jTXP@�`��3$g�`ƬZ7�RE��EU�dC�I�k4Q>˓��8;��8�����[�&����ȓS0R|����l�F�rQ�R� K^�l��u�rm[�T+n����O�]C�:�d��qmH�y�{r�֝۞T��g��������TO �ք�`l��+D���
W>Z�^-qg7p&��@�+�I$V�Y��蔯~��>E�	��}��KH8RP@d"�L)D�����P�����K�_&n Q4-�;}_�"����	N��~Bi�)H�M�1�[�nɚ�dņ�y�k��(JDO�Y�X�"P%ƍ�ybI�#F�=���'eĂ��-
�� Ϗq��x�?L�9��q�$��P7Qф0�W-�7=� 9��-D��p3̝���,��/[� ̼s'�&D�$����r��8�X?�)��"D��:�,�
1�����?zٔ@
C�>D��Hǝ3^μa�`�fN�ɛd�>D��h4(W�s�� �Q�Jt����+D����$f|��f!M:L�6'D�l� �$kVӃ��.��ܙ���� I��eta|Riؕx30q	AK D<�u.�0>)�`�.A�xa��L\�{��4S)����ۢR�\Ʉȓ=�B��� zg^9�4���`�|������	�g�O6�#i�|�ӌ�i�:���k���y ���G$!B]B�nSL��3+-i��5��Q�FĮ8Ѷ���=�Ъ�ZL��~�� �u�+@�؊��U�U��K$U�.�H�㉒V�R�3s,�Uܶ�sPJ�<�h̀6m3~`p�A�V�W��X�!�'��`#��`���I�$�N1�
�+���@�+���W$��W ��V.��+0^�' \i��8|�B=K�N۔Q~�H��^= �7��!��]G0-��&R�}��ɂP�ڠ(ƴt�DҁXa6��G��-@����X@:%��O�"�+���M7g�q�r�U(:� �  �J�5�az�j�A�X̓^j��h�DηE/���d�Q�0�~iI�״SC�|;��N
�`�ח�?)uϵF+����!����'���t�է,��"�h�Z���L>)��CX������@RU�2'ت�2ԐթK���	�'��<��Q���l� j��G6�?��l��$4q�FI�G��y2�9��xV��j�Yv�J�T&%Ё�ì�1U�L�1�H��b�'2b���<���iÌ  �tR�R�z�rP��	\�2K��j6$C�ɽT�.� �GD�wdA:\XK��ζi~<����dB������r��d�V!��? Pp��z?1Ǉ��=�9X$�O�(�x2�݆Y�=�`"$,O^�0��S��<kܴ
i��T\- 	� �0��K����^}��ѳx	,e��Oqy��W
A����Lr�I�0a*W������5�8Od=ڥK��`e8�4E���˷��G�b��� M 'X�]�I�(��H��1��dQ��K�:�Gr���
�FY����آ;� |�b�A�\Y��E�Ơ���K�O����N�R3d$���S�|�Hَ\N@ �vb����?�Px���o�2�90��4��"�+1hn��iқ���.�,��f�n�>�) �n�D��|�n�7\�
��Q�R0[�4XE%FjX� �c�$c�
�y�Z���
Z*:���.�-��)��Dl�^Q{�4q�ص�M�"~nڮ/,� {Ce	,���@�
x�O��!���z���	Wed #�UNJ��#KY'��I�l��lj��\X��y���K��ģ���en�(X�ě6k-���=a�u�'UN�u���?K�`c�Θ	9�<���9D\�%��'�MԋόO�����,L��C����h�~����]�tY�� E�%n��!�CA"�!��ŗd�`T!wj�( �sR�A$D�!����`�pP�
�����NS!�#�ڝ��I�O�
�����%!� w�y�$�.Oٔ"t�)P!�dӃZZBa*QkRC����c X�m	!���+z1�(I&r��d�q�@�K!�$�φ�H$h�03�� ��34�!���~�0��6.ǁj��\��n�>}�!��
Y�XXcCY�f���@�^�!��O5��e��H��S�Ʌ�e�!��Q�Pd�O� t�,�!�� �P�c�P4"i�Տ�mX	�"O�%8�mR�#���0D�٣[�T�4"O����BOS$�q@!4��"Ot���B�*�3R��K�Q��"O<�����H?��� ��Z"O���K�#b��S`�C�p�L*"O,}ᔯ�N"&���Y0X�hٵ"O6���(��:�c7cP�P�XP�"O` r�F�M��2�m��~��4"O�i�ӌY4̖�a6>�%lO��y��ا[�����Je��f�A��y҉&0���0�(�NW�����'�yBL�=�f��̩~e���b$*�yr'S�I�v�C ��8`�ĝ��y҇G-"B�D�E� v��yF����y��{��er��}b���(:�y�Cԛ3ʘ����t�i;�H�y�䞁,<���˜�\�*�:!�R"�yB	�t���Q�"��U�>i�`���y�%�u	<k�њ������D��y2�/'N�,rC Ս�&��Rh ��y��I6O��2���3}�e:3���y���7ܮ%���
5��(٢ �:�yҀ�j^��CP� ����=�y��`��aϾ�����&5D�p���70��d�68��-3@l5D�hj�藇:�%�Y�^��c7E<D�p�bF��\v���f�U3��L=D�L{b,ښ,h�
�'F}�)ju�=D�8f�66t�k� �[�4�91F;D���2��y�ұ� �U>4��#6D�Ъv]�K��Spd_�jt�27D�D�2�Ջ@(�1�?�ѐV�3D�x�1)�h�EJ�C�	��a�#:D�����6W��+"ݍi����%<D��3�IǢK1�\8�iO/� ��(9D���ᄝ�nM�A� �>�ꠘB�4D�ԋ�^W�����	Z����S�2D�3�N
h�N��`�K?v����2E3D�8��4�>���"ǖ{r-
�#1D��(��&Tg��9��ѿ7��(��.D����dE�xAK��6�zܠa*D��!!��DX�X3���8�T�r��5D�8sB�'A�$T�C�^�^sD3D�����ɣP��l�q��.���Z��1D�أ�hK�WX.3��D=D�� 	T�"D���a�v���y��^?Q��QBn5D��	�Kфej����Oe����$D���M�\�x`�R�(�j)�c#D�h����nn���e�!^��1Po2D�Tf�alHU{��+*.=��3D��I��3s(�ّ�E;7P	��.D���𤘋+	Rܱ�dB�y4F����.D�$1��Þ*��ذ��/�:��d�1D��{w@�C���� 1T�e!�5D��qnO�e��&� �Xc�'D���N�9Ʊ�P�S�<^�`���0D��١�.�R���]�~zu�WC*D�8����&OC�i�O۪|i@�o+D��x6��	"Q<�i���6�HA��c&D��&$%=T��Y����0��Q�3D���A�G�7k���*
2����!2D�`�І�F��XЂi_+���ڤ�'D��h��߅>����%�ڷ-{�)׏(D�� �I�F�"�S�]�xK�0��'��)@ �$*CI�&g�H�@��������rd"D�h[5鍽{�ޔ1f��<Fl�\���"�K� |sei=�H�(���n1(��q���$�ʅ��"O��� 6��Irp��H����oذ}g|Y����)��<�qN�xd-��/� w;��T�Mx�<��%A0��k5\6����U�<q���)���a�%3\O����#ˬE����F<�)�C�'�,���X/�L����fA�A�*W ~e 		�	� �y����:ij�l�6l4� ��OM�@����&�(��Ă$	B
d�^�13��0A��S�"OY��� ��!�f��()��Z�Qf��`�H_#��)��<� ��1��E�$�~5"(��G�<iW�^�x�<��w���e�����`��<�g,CzXr�`&J=\Op�z���i�C�?	X��q��' �U�r���!�� �C��"�����m0Bԓq-��y"BʒY�H
�k��b}�q����Oꤢ�� /����$Xk�@iU�4#2p�R �Y�!�X	�����L$T���ψ1(����Ѐ��*ږ��L�"~�|�����U P�j,$�@�ye�]�ȓ_Q��X3�ʀH��L˲(H2f�h�ITP7��Ű=�`���&����!ȝd���
ҥFX���5��	B�E&,���L1hQ��,�$�y��؟z3�]����3�����ą�y��,ݔ���'Q9#,��C��y"fɨQb�:ƂAA���p�dѥ�y�Nʊ��6�M6.P�@�K� �yԀ)��MΫ_�`�Wƌ�y�EM��J�ΑLHμ���A���'Iʴ���R�S�'9
�*�̜<?6�H�HD~�Є�"�R�ʔjR.��cA����FQ�o�m�ɱ�LE��Oq)�%ά0���Ɖp�IjdO�t�&B�ry�s�,�6d�!�#�Jg,���_���>�0@'6Z����i�NR��rA��wX����RM����R�h�Ԣ�=E 49�a�0u�i%�-D���ǤK
��[�	ξW!�PL*�S~!� "�Aؕ�M��B4�c?����t|�9Q�B�#x0X(��+D��dM>Q����F���~�᥎I���+۾Bjn諁H�[�vb?%�Odhk�a�0c��x�5
'd�HO^tЖ�&]�򙛣LA0m�SÁ�n�tQ���߸8�P q��<0l��I�� �ʀ�ߒW�(|`j�"F!��D�>&�lm�� ��D�J$1c��$/�=��"�Pn���Ԑ� |��\s<�󌅠>�f�34��k�(T	�%8�\ ��-����Y�L��:U�ܴ��D���%8t�	���%	��n_�T�t��-�S�r��B��!�D߄V��;�lK�(ؽȥ��/��!y�� �θ��`�	YTX���o��% � e^@U9�NE/,�^p��O�������y�<H�E�-�H��I[wZ�)��]�r�hR�̣i&t��Ռ�iq2��$�'3r��C��^����v��	aO�eb�'�;1)���2/����:�i��Ǻ:R��.8L��M���h��ǉ``�(��ďi߈i��.�|�h�o^��ZQ��N�-e�bL�a`֩
�ꥨ�'St: ����UA���d����V������^eo��za�W{Sv@�O=��]Y�F��|���w�N�x@Ư~a&މ|"�=���h�@�@$F�d�b}	�'�Y�]�և��QKz�+��gv��eˑE�I�fr���%�1��S�~����e
/���[q��*=�џ(��"�/��aҖ/�2|�������@cœj�>�����$�h5���|��]$�l1��I3+������<r:0�E囚g�\˓C��`L�j`��#u��j�|#}�K�P��u`�"^-vl41y�<q�H^4{H�r�)R=Fp�	��E���yy�G�)6�"�sTg_�)Xȭ'?�ԛb��)zc$���lڨ�`c�)7�Ћ")�kh�IW�#3��U��ʝ��=��!Vv� $S�e��P97#Q�F���	Y@��ݰ�O.OA���fw�3cF��y2�g>�3ǓQ�F���A	��y/�q�^u$_*1Ķ�X7-Y8��'�n��6l|�G��됇@��8�Ԧ�4,�Y)6��5�y���-b���y�m�.[�`�V+H�+B�B6l�����:PQ>�S�? 4i���2u�Y���S(~��M��"OHI넀�) <)��,P8.�>4�4L|�R	� ��ă�|��qArخ��r�z�"ܷ.q�C��c�X]�� ւA4���	��y�ꝌG�P���/?k@�ywa���'"����N�P�t$��Ӿɪ񙗨�f`�8P �I�C�I-+�.���O+Q�paF�5N��͊m�X����*O:�K��Y�TA5b¨]�s�Eܹ[� ��!/D�Ќ׀TZ]A���1�lӘ�2��@(,$��J!�'���5S!`Z@ڥ�9$���
ߓ\_T�S��^-(�
6�M�cOZl+f�4t	���� X�Be!�d�t[�����P�S��[ i�O�m; aL(�R����0�`�F�uY�2��2o!�ċ�ٰ��jVH��C뙉'�̋��J�b��OL�}��9�xd��M�હ���,�� ��$B�䓼r��K�F�MB��ϓ|B6����>��=�B�CJ��yI���N%fmb���C8����Ʌ�F�d]��Z���n�=Є�G��,2�!��=w�A��@��!Su�ǅj�!����ad�@�G�T��b���!�Ę�}`^��ŝ�D�{G�~�!��L�cU8a��O㪬�T@D��!�""�I2bo�7٪L�m��\�!�F!L|ꅩJT�i�aPSU#|�!�DN�!].@V������Y�K�>X����VP�0��\��@Ӗ]3�0�$stم�0o�*����̟��gJl��%냯K�l���Ǐ,D�P��/����$q�M���4��O q)`�ϒ�~�eϡR����G��A�O�B�QG�j�)�)��n<Q��"OHi�dI�0�$0�%gG�e0��7�O�@i@sJ�Yw~�Q�'Q��Pb��h��Sq�{�+
�TXђ�,ON�����`�*z��05	�`�E�5,�M
pj�aB�$	 �&�?I�Y��N�)v�/lO~ęU�(d�#��	/s��a[��r@��\�����ȍ=���0�����)�Ŏ^3j���[wb����s�,"�
4v(h�'۸��@k��`pC��P6z\6AX��
�.���F�U]}��eaנ��+C�|J��y[8Yp�w?ęz�^!6F)ф�v�p�(ӓ��`R�*f���A�U1~�~m�b�Q;��QwkI(�q��ו)n��î�p�����'{�nu�Bf�
>���<a�c��98������i���Aov�h���/Q��P���N;O�!�֌@
�Q3���*Bl]���J27زP�s�^+-`M���x��8K���$?��]�
�8�hy5�?ZA�b%��pf�8�S��M��ȂX�<Q N�Gx��r�����
R��h�g/>k��,<�y��E��CL^�1�
O�%��HD�RV� J��J:�L� o�m�T�J��ȠO��{A��#���ʖ�ĬQT���z?�o��A(~K��M��8:�F8��l��F.,O��IԨ��v6��48�]�ʲ�����[��0�$k�K�S!�K�I��= Q�Mcy2�E�+�8�� �a�~����V03�@���oFwVO���e	�<����4k��=�e,��R�:�q��t��}q��n��
���S5Z�j�@��S�\��e���I$�'^:h*��A� \t��#�Kuh�� �B'`i��@�z=�ԉ4�W��h�0�ӼYa�ѻjP�6��m��_��ć1�A�fAV5���u�B-v�ب�E�$b4Pc|��b@g�z[I+���V4��'���S�*�t�@SN��*]3u.�9@Z���:-I�Jܶ��V=9l �$�Kc���!!M1Λf�G�	��� Hg�ӧ������o#�#d�����R�@������z����0|J��ǺC�l����}�̭+���^}r���7����4.Qx����S�}��9"�)��;�M0��P�{�qO$�p��@	���S���\J�@�{� %��i�`�B�	't�`	T���qKʘbC����">)��N-�ȣ|T�<(��S&/��?hpP�,RP�<����7 ���)��w������E�<�e1)�2�+�$S�R�١�%�}�<�a��F��KvC�K2�a2��}�<��JC����j��MG�%��a�b�<���Y�FE6��dɚP�P�
Z�<��k�$��$C�ޛ0��@e�P�<��8y��@�<��UX�+Q�<� �10W�'%jl����ш,Z�`�"O�"�S2�|�2�S�6� �i�"Oޠ���n0��a�T/��Aiu"O�����ОMU�-�BgM �X	�C"O���nV�>�y�#HA�,��"OpP��İ*:�X��S�1�65!!"O�#AF�1vq��"�����"O��J�DL�ð��ʆ��I��"O�\Ba���B`Bn �?�luӴ*Od�Kg�[��=���27�8�	�'��]�df�/;Y �*F�%�"��	�'�EG�D�i����/,l��@�'Ǟ)Q�(���L��ō"e�f�#
�'mx /�fz.��@�>^�0�p�'�
�p/4
��p�G\!y>�8	�'��i��W�� ��g���49ڽ��'0f�	.$r)L��e>Y����'�(���fϨ��i�Dȣ;���'��ar@Z�,� ���5ː`��'�t�����]�T(�A�.[w�Mp	�'��,	��R-Zwba1�W_����'�j%0�ƈ�3R@� O�W����'à����/�8�d�E)�)��'u�x��"ε��*P
M�:"��'m$�Z�Yuj�R��F�2�6���'����cH�,���fX2%$ٺ�'�6T37Jͦi4"Թ��(:f�'�~-���$(�F��$C U�&���':a[�$��n���\ �����'�~i�e�֓M���1허)����'��k��>E|�a�`���_�4��'@ �*�͂c��tBӥ֟C]��a�'����`��7���z��;�8I�'�L�鷈:w�ā��$֪S���
�'4���V�^<�%� �I3��˲#)i:��Ë�1-����|Oȝҁ@�Up,M����<u?�]��e'
�y�헰+�����������L���fɊ�ohy��,�D5��ȓ<�p0C7HY�{@�T�Hr@�ȓP��%��^� ���F�e����M�����G3V%�-�"NQ��b|�ȓ*T�ƭP���ӧ�	����<�ÇGI���O���J�)V�@Er�Dd��
&��'�`7��؍�'���B^w� �3?�')�d�$�4J�f<���V\���kFA��E�,OrE���O=L��W%]�,(�hT�g�B1B��T�|T�	U���(1��	�fǓ0��	�M�d�8 ���@}rh�6i@!�֡@���	Ll�OE�Ub�H��%v�u��h^B�HSd�V���Rr�7��%���O�?�yPƋ4%�А�œN�	�1Ad�L[�@I�A\8�'���	ׂl}@��"l�,xԜY�)�ZQr)��'�,Ô���Mx^Ԃ
ç)�R��G��jѨw,S�R�x��Ż�~B�=c�P����+����O� J��p��cyp%%�����8=|E�X^M%�����۞r��d9�����d��K�UD��!7(�<a�kFy��IZ�a�J����w
L����تΦ����,��	�'�8<'?-8I~�6#�20eb� �q�$�6"
�h2И�0#�V�m�;a"��}n:�+	�{Q��B���=�4��/O�V������������|xX���S�{��@�b�*wU�  BF� @�h���OV��'@�2S�W�?����j�|_�<еJ�xg(%�@K}"��.U[��3S	I%���Z �\ �+ZGjX 5l�	C�D�$�����x�f�E�~�>q(7���>sPF]JY�@��`��S�p�^3�ݠ��Tb�ѩ��\:�!�$-]��J�O 7.5ry@p��
%�!��/1�X��AӑL��(c�'�;e�!� 
g"�9��L�S�Z���O�i�!�d�>.(*yJR(�8φ(K#��2!�� ��S0��?iT���J��p��E��"O�)pE�ڸ��q
���7����"O��!���o�T�ZB���8k"O>�`%o��%���($���mrX��"O�I��ŨN�@"q��M���ɐ"O�h��K��P���	��=A���"O�;��Έ@r�� ���0/2F"O�%�`����	�b�:"W�c�!�ٳBl⸒7/��>i�	�v�ͧN�!�_�S��`��-4hf��nE	2�!��4d!�Հ�m���P�L�!�FY�<=�;U6����"�!���I#���'��I�pxQ�B�[�!�P�R��A{U@V�H�P�����&&�!�dUz�>�o"Z�&H� ��!�DX%=��b��&Z܈c�.Sk�!��-_$*w[�byI��"!�=~�,���@e>NEZ$��'p!�^�@�Z�0��L����-z!��2�`�"�F�SH�!#g�<r!��3WO��j���a>��B#&�:gp!��w`�t%R=r{7JB-S!�*W�|{���-�T���F!�%)�����_�m{�@�fA�$)!���{���;rT$d ����>Yj!򤌆@�T�3b����E���]K!��[�R��!S o�w���(r��y�!��-?���J>|���T%�?F�!�d�.���g#R�tx�U	��aK!�D��_a(��ԁ̏P�ĹQ)B�#F!�כ[� �k��(��	1����m�!�D����4#P ��0Z� T�A"[�!�W�y��q����O�@�	㉈�!�L:o�.Q�q��6�D9� ND �!��0-PZ���ʅ
����Т�!�ĕ�GjLfB�Ut��qɅ�!�$=xޑ�a�: �r��6)���!�d�&@E��
Ԣ�F*h��P탄b�!�D�>|�t��$�Ux��<�!�d�F������'���ǂ���!�$)3��c��-Y4Re)G�N�/�!�]%o����ʰ*w6h`�R�y�!�$�?����ӛjZl}��`	J�!��͒Lŋ�̃{���@" ��8.!��LJV�P�b*��e��rr�̇%!�DÁZBJݲ�	�r���3��|�!�o���`$Z�t�0#� �!��4E@0�#���4#�aD�!�
'��4��([c`��+VN�a!򄛙R�&�3&�8nC�11�lS6rP!��VG;Pp��M�P*Z}��J1%�!��Ǟx	�B�3��*�jѵF�!�D[>Y��ģ���0FըQ��O�!�dNcs�HA`��� ���*�!�d %-���1&a  �0�RW��*U�!�Z�4�& ��LSX���g�<q�!�d:9<�5q��4v��y��Z?\�!�č��b{�M��	�R��фW%�!���}P� �`߇�4M(���G!򄀃=F$`%FP�d�8����ZIV!�A��� Ʈw�y �\%SS!�$������-�-a��7L����R�5�r�!mڹ�lI��y��֬P��D�!��}ɦ�9&ڗ�y
� �D�g�ʁgF` ���!j.�#�"O����Z�<M��$�UW��Y�"O�a����"'K� �C�<o6pI��"Of8{�C�>�j&�<`%pE�7"Oj��b�Ēx{�HE�]�5�Ekc"O�)���\&0�@8����2�`"Oz���ߋ�2��v��	� �r"O:����
)��|Z�#	Q�ؘU"O��q��#ҭ��E%Җh�2"O,���/�`����#�+)$ʬ�C"O���D� �TK���d`p�"O�)sW)��Z��#\K�l�"Oʴ�P�&�>�I��k�`���"OΉ+��ԇX���X�^]�~@BW"O��D�ϯU�����KW3v�� ¡"O����n7����٢#��	b&"Or`z _�
�xE�s��r��a"O���&-L���A��_1R%09"Ob<�'gq�0&j�1��I��"O5�$�B�E]�e*ѹK�}��"O&�xD
N�0i5d�xS��i�"Op�P"i_�1��0��P�'<L�5"OJ��t�V�H�� �%[��§"O�|ђi�"rHhׇ��pҐX�"Oа��C�$���ǔ$��u�0"O<���gÈP����2&�-�x�W"O����
�HO�Ar��W
)��iB"O*���ܧ|X��{��Ü)�X��"O��R%́�#��cg-��#�V�iD"O��qv��B�Ѻ�픛"�d�S"O
d�d&�6��X�M�d.�qW"O5rc�7>l5!���Ѵ(�"OH Z� ˕)��`+2%��[�t�"O��`��8��ph�a�z�Q
d"O������(���OR����"O*��uAH8^�~9��d	�\�R�"ON�"(�;��	t)�._�,5�"Oެ���3�j��'y�.�C3"O|��n�r~���`��;m`Z�@�"OB�+pD�>ڌh9�k^�r�z�""OD�[�N�7'��y��a�t�"O��*���k���U�/b	I6"OȰ!�f�,J�COQ_���V"ONI�S�ޟSs ����g��%"O8���K�{�������|�� �"O0TZ��H�sm����K����"O�%���()���F� 9�(d	P"Or(���f��]��Z�7�P�q"ON`��c�d�YC�k���*V"O]���H$"#j$��l�E�z"O8���ӎ{���I!0�d�a1"O�l�kȗcGb����kYr�qC"O֥�U"���Ait�X?�ũ�"O��{��ѯ2�@,	��̵P�0�"O�;���a�U�� ԛ=A� A@"O$XV�v�� 7�1|���	�"O�`�ǟvg�t�U �V��e1�"O������4C�,��(Ȱ	5�u��"O���#�X�{�����@�&y�D��"Oy#畑 ���'�D� \{ "O.Q�C�Q3
�� �wE�]1֕��"O�9 D_�"����]5x����"On\�g���p�L��N
��"O�FI
�phQ���
Ҥ��4"O� l!pa��	�d ����/��9�"O>�"�[:J�0�"��s��A�"Ox 4
�:|��1uDFb"O8�1�˞I���&��d�)�"O�n�*��Dh3I�����OժD�!��Ƞ@:ݙ�l�j���0��!��Je4���J55�Bu��D�!�ć�?Qr,�g��*�	`d�!�D��V�@кA��"*�j��D�!�dD���1,�!�F��UÁ�_�!�{G��6AN�/^Xj�!�H�!����@�Bd"\�f)`���4�!��V�j��M��-��`p�E/�!�$�L�Pq��C���=;�D�F�!�d��Y� ���
-'��I���P'Oޡ�d�$5�
�p��:}J�`Z�A��y��� i��S��O�]k��i Lӊ�y�Cݽ|#�K�,C�H�ɛ��V0�y(C�nhct䔤R�tH!d��)�y��]1�̀a�ڟ���
����y�%����9�ԥu����D �yb��r�ŋ�'o(D�5��-�y"'S���p�sJ|H���d7�yB�NFP��e�)<m��(�	�yRlZ�r�B6E���!�ϵ��4��'���@eD�1=�A+&Ɛ+lX���'�4��̗�xO޸be'�	r���'�^�J�V�9�rk�/�+�:Uq�'���QmѢG] �td�3
z��'�*B�@"�@�3JC%����'w���fȀP2<�B�+U��(�r�'t�����W�������Y��)q
�'^u;fE�9}�0�K"A�����'��	�n�?w����B��<C,�J�'����a�Т�F�5����'3���@�1��`"6��,&e4p��'��ԁ�Ɍh U��X3�Xx1�'ǾMA&���S�X!*����h
�'֌����+U8Ȑ�tO(u \0
�'�����.Km�D0�	^<t�X�	�'Bh%7��w�pT��9 �D��'p"����X&���#]&Q�;	�':�`E��q�<P6��C�
�
�'Ѹu`Qfխ	e�l��4�\�	�'a�})΄1l��A���W���\�	�'ox9��j�T|ma�\�_���'�x,���	
 W���b�� Pm��'J���e杹��,bả�f��i�'$�����6^����C&'���R�'{�E�biB�{�0��#���P�
�'�B\��c�%#� ujG�H4���@
�'�Ι*�@Z+L%�D!��-#�JiB	�'�xe����b�~l��-ƍ!�P��'"����L�e�h��2l�
eI�':Z��aش"*���e��j	�'l�idA�O���A�0$�i��'��4�P�	��+�F�#@*�@�'�D���Kj�^�"��Dh5��a�'JhH����L�Re[W⑴p����'Lb�"�	qF�]����#��Gy�<aw�'\��UrU'\-p���AFPt�<� ]�L��@��E���m�<�4��0�6i��[0ޘ��#�	f�<�2�����dE��)Nq��hM�<�+w�   �   �  ,  �  �  ,*  u1  	8  "?  eE  �K  �Q  /X  r^  �d  k  _q  �w  ~  W�  ��  ې  �  c�  ��  �  '�  ��  /�  ��  [�  �  J�  ��  A�  ��  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C�>����鞿6�!d��x�^��I��~�!��
�l����v���:�9a��:uZ!�L�,Ƞ�#g��UԀ�e��t�!��v.qc�ʁA�P{U�C-h�!�DD�x>B��cG;c�lK�,��"�ayR�	� Q2���F��u�t��� �/��C�I�Ld֘8����D��T�U�#�fO��=�~bh(e������M?��m���Tg�<� �������T�����R�g��dR"O���ѣi�A	�͖<|l��"O�ȁ�N��SO��µ'�#{u�L�"Oҕ�sGY�>u�0@�'B>]ԕ�b�'I�O 5j����)ɲV�л�"O"}��J]�P#JLa�׊R�Q�֓|��S���O��Ḡ/��l"�88�n�:!�D�	�'X���P��u�҅� D�l7�<��'{���6f-虡4��	.�<�R�'L�Q8�C d� ��욯zA��'a�l�3�F!C����4},0|ϓ�O�4 6g�'���z�h�!�P�R�"O�$Kue��Vrl��MΈӲX�S"O�!X$�ZD��z%��B����C"O:0���b�V�a@���VĪH��I8�\��׆pT����Y)i3	=D�$�&���;�#!a��9��H7D�|��BP���x� 脖~g�T�#5D�H��
�Kh��Fo�Z�s#�'D��)F�^��$H�/ǐ'��(#D�8�\�.V>���bYO�9�4m%D��3"�Pq�f�2P.p���(B��$K
~%x�b1Fb�la�CN�.��C䉮T��[#A�$I����(��AC�C��H�XtN)qH�!!��A��C�IHh,����s�6C K�R�jB�	����#塕��Z����}�B�ɥ~�� 2
?<�[�"��nZ�B�I)&�ĝ[uj	�%��a��;�hC�	�f�-� ���=��d�E۸a� B��;}�܉�e�1(��1��ġ=JB�I�!�\3�oԾ�p��C2h�C�	FxXz�g��dp�Հ	c�C䉇>�6���a9yVa�W�vdlC�	�!2,ҧ�?U�*�����5�0C� XwZp''�q�1c̀�ThfB�I(wM��+����k�I�@�ӽ	LB䉆���F^�=*Q�@GB�	�4�ܵ�!�� (Yv	`s��7�B�	?s�r��d����hj��I(8�C�	�g��d,�(M>�h�h��q��C�	�TTx�5��<�� ��&��C䉿[.� �� �a�P��/ԌV�tC�	3F�!wFY�b �'NV��C�	>=F�m�FǵxZ8U�ց�	tLC�ɦ:�p�n[�u�ҴY�!ӣd�BC�+;���U&�<b��T�@�����C�	<+A����Ǜ �R�I�.ݻs�C䉂Ԫc��T/T.nL���ܴS�B�	->�N�9�N��T]@xËZ�a��B�I�E�Ĭ1� ̮j��� A��'�B�I8[�2�r ͫ���TP�]`tB�$�0C$�!O�偷ƛpuNB��]EdP�o�4'��m
D�ُ9.2B�4$�t(*d�8X�}cRd�+DB䉷L�T���k�2n�i�CE�[SB�ISQji��6��{@��/'�C�	�sϴ�;u
�?�X�:b
��~/�C�I�F!*t��N�:�0�h�-	NzB��<�C��3}"%���CW@B��&`H�ܸ�Ζ)��p��+� .fC�	'�n�x�$t���2�I8�^C䉟2�F�@�╧Nt��q�ŪXtB�I15D�"� 0h},�H���yA�B�)� ��aF�H=�`z�aN�'b��v*O��xc���2�~�0����}��'���� 0����
Wl��*
�'��ԁH>pxcG�o�����'\za�2mF�3��H��ˀ%o�����?)��?����?���?���?Q�=�q���-xpB�ѧ�B�j��9��?i���?���?9��?a���?i�vD�U����;�Pĥ��?P����?A���?���?���?���?q��S�x�+��� &�h	���#OVlI���?���?���?���?���?��j�$X�գ���l�o�d����?a���?���?����?A���?��(b���[tu��+�B�h�J�2��?���?����?���?����?a�I$>�K�m�����Bl����?��?	��?���?i��?��,�lyGm�1��x����n��,���?��?���?���?����?��g�x˷EǂP�C���'�
�C��?����?I���?���?���?�7ⴹW)>��
A�������?	��?����?i��?����?��s��A�N &)*�n_�a ��0��?��?1���?I���?����?a����*��)[�|��� ��r�J��?Y��?���?���?y���?Q�z�(��P��
^CB�ve��A�Z)[��?	���?1��?)��?�c�iC��'�:�i�ƩQ+x��r-dԙt��<A�����0�4)�f����s�P�p��&�:�S�C{~��nӘ��s����9��S�Z�A�u�_�ƚ-��՟�R�(����'Z�	P�?�����uc2&MD+0�ѯs�du�����Of��h�d�Uk�19�A�v�R�q�2�a�����#1!#��L�'Ad��w1���G�[	7��%�ECN��xM9�'$�?O��S�')����4�yR���B�@T@��)T����pM��y�9O�����ў�ş�%�dȌ��#QV5���%`�L�'�'67��-�1O�0�vg��k��Lץ
�ؑ��/�����d�O���u���'|��Gw��Ȃu B�}{�O4�DK�1
>	���I.�?��H�O\�p�n߲iM�:Q�F�Bc�m ��<Y(O���s���$ޑ6��$ѳMyE��uOv�`�ٴX�t-�'f�7-+�i>�ꖉ Q2�8��Q�'�a���o� ��ß@�	�ED�n�q~�=�,��&c�<hJ��~KL,�&ş)���#�|V����p��џ�	џ�Rp�N
W,
��IV�LH*3��oy�u�mIB��Ot���O̓��d^��%D�8Gr��i���Hb�Ʃ<����M��'L�>���O�;5($s �� �h��MM�Kx�S� �>��@jhy`�ьO�ؖ'c(`�C� ��,��D�	H��'/��'�����S��ݴ`� 	�@F��	�/􁻂�D3`.d	�Z�����g}r�i� 	l��tK#�^�p� �G7Y~���D�Uo��m�^~�닥�ܠ��w�'ojk�3=� !e��!'2<)�+�T���O����O���O��$9��b�.Iy�$:?F ���>/�(���՟���9�M�$)Y���dNߦ�'����M��d�di6�ώBb�(CUFN:�ēM���Fu��	]YD�6�7?!g����(� 
����s���?�Jx�$��E�F�$������4���$�OX�$R)�e�5ᛧaU�l�FnUd�$�O�˓Z>��.M�\��'erZ>�05#�+$�����LDA�=�l)?�_���4 ��v
&�?]SGKE!F�:�tB��@¸��4u T0h�I3���|��`�ONd9L>9����IF��Q.2�Ψg�ކ�?a���?����?�|"*O�$o��Zm�U��h�r����L_!h��I�������I��Mc��B�<�4w���E픧��=9� S{$��sǿi��7mC0H+�7�??Ae힧����3��[�j�x���,Ү��qe\
�y�P�L��ܟ���˟(����ܕOΰ5���m��eg��$��XXmq�(x��-�O��d�O����dD٦睈B]�a���q#~-�
ӈh%ډ�	��
O<�|z��0�Ms�'�ص 7���NcHLp���A#��؟'��)�4Ǆş�$�|rW��S��k���FTn��"��6%�Rw�\�������	hy2�{�T�*�OF���O��.���P�C��Ii�r�Э8�����D�O�7��]�'e�:D�P�1R���i�d�	ǟ$#����2U#B|~��O2P��	�x���0'��(e�(ј	h4&ז�"�' �'E�����"�!�3����^�qo6`x3�C���4.G~�S.OBl�l�Ӽ#����Is�y	V�A<e�L��E�]�<���?��i0�a�ia�$�O���WJ���!*�v'z���n�4���2#�F�RUp�O���|����?����?����>4��D�5����LN2,.� )O�o��+�m��ȟ���X�Sȟ��G/�-?�н�d��Y�b�*�(C����I妹��4Sg�����O���H�3U8�UY�� Q�YggI*Ly EY��d�*\�n����*h��Of�(2��2�K�4�X�d��蚘���?	���?���|�+OzUm�
INL�ɺ/?� IRa�8:x(�cC+��H��	6�M#�2$�>��?׵i�\��R�*1ՎQ�G�N��Q3#7��:O`�d>Bf�Z��Vb�	�?��=� vmS��A%1TCV:l5t0s�4O���O6�D�O$���OZ�?ᘡ�.n�Ȉ�ɇ8�Z�#"��Ny��'_F6��+5�)�Or nW�	&P(vă����j�*@M<	���?�'hҰaش��d(<	��E�ϢiR�|
��G{J�#�C*�?�&�,�d�<ͧ�?a��?�U�O�"ߘ8{V�5i���Y�	�?!����������ٟ��I�� �Oh�I���.�J�*��6�&��Oܘ�'R�i��O�S'Y��YA`�<1B,�!!���t�Dy�eo�()ں�s�:?ͧZP��DH���bd��q!�M��1��ɮ�	���?i��?y�Ş��d�ͦ5q���$u��j���v_����+^5A�X��'��7�>�	���pӄ�b��;L��6ʍ[=���EOH��P�4*;r�4��$��X;~���'��5��]�5ɂC�5{��W"���Iuy��'�R�'���'��[>uP�Ɠ�e���QBOϫ�j���gۀ�M�Q�?a���?�H~j�v}��w�"𠱩�
,��(�EC�g�ԵSv�b�v�l��<ɪO1�0�1�}��ɡv�j����W�Jq�偄�qUd�	�js~q��'6H�&�����')n���J�X�����V.TEK��'��'m�Q��"�4h`Bs��?���'�N BT�O9z�*q��@V���i�B&�>Au�i��7�WC�ɤi��9:R�II!b��2
F���*�#ϟ�t�D�|�c��O�D��0��#�d@(5�pBvI�(]�
�c��?1��?���h���$Λ<�f��S�[�8s�Ao҉H���Ϧ�P�B��D��:�Mk��w�t�d��3[˸p�WlI��`�'F�6m�צ5�4}��`�ܴ��Y L�6 ��z�v-c���m��!�@�~���cB7�Ľ<ͧ�?a���?9��?���1]lM)eeA�S3���r�U���dW��M"q�ןX�	ڟ�&?�I2de<��4�E_@�y���إ
��IY.O~�Dr�>]$���[�Ş_4�ځ��o�(M�wӄ#��!���\����B��f�	cy�
�nH����K$t��Y@��f���'zR�'��OL�ɪ�?AE����@g�ż'�� Y��'g�@H  ϟ�a�4��'����?���fk�QθZ�K[vhrYyA-V�2�h��iH��e�X����O�q�d�N�& S�b�ײ�0�����Z>��O&�d�O����OP�d1��R�L0B��7�^	���->t2��'$�ix������?�j�4��7����N�.6�6�`F���\0�x��'��O �Ҥ�i��I	T�{��&L&�`��ǌo�� �p�ؿvn2"Lf�	y�Ob�'�Ɍ�J�4�A()8[P�ԗ���')�ɮ�M{����?A��?9-���(��Ģ|.��S�D�	���8ѐ���/Ot�$g�\$&�ʧ�"�c�X�n-�HA��:G�2�#��D�$�N���"}~�OT��I#z(�'���3V��VT�[r�ϊsjV��V�'sR�'�����O��	��M�1%KmȾ� #Z/��
�!��zF���.OT�l�`��/�Iݟ�w��	[��ٛ!ǆ�}�\E
\🸠�43�pڴ����H��Ÿ����+Z>�$��2�r�U�1�D�	my2�'���'���'��X>�WDF3Ӕ$��,%s@]A����MK����?���?�K~�F!��w�h9c�[	T�V��W!�_wZ����'�2)%��)��+��6k�� ���M�p�!�'аC��б�$r�����#|B�H]�\y�O��Dؼ�p���f��سQ�Y�4��'���'3剸�M���I��?���?�sd��l<dK�C��L�2`C�����'��ꓬ?I��H��'V�Hq*��Z�,ʳ��)+:(	(�O4�ٖ��(J P:`�IN��?`��OF)x$$�3���Ԥ�<�l�`&��O����O*�D�O6�}:��4&Te*��4k�t��0FS!{GR�(��K��f�ɸB�'�J6m3�i޵����u;����$þ���i�j��������;ش�R1޴����(oȤ�'|�8��6?��H���9$i��*v�7���<ͧ�?���?���?���=|&�u�aE�L��%9uFY����Ӧ�1
	�,�	���'?牝T�d-��!V1b(�3���>�P�S�O:�mZ1�M��x��t���k�$	׆��l?�0Y%ˀ��T�aH����Q0�����!"ؒO��.Ɋpk�@��#J�����|���H���?����?��|�/O�oq@v|�I�E
j�!�J�� �VA��ɺ�M3���>����?���i'H����?U�zh!π�(�S2aWd������lA�S!������ld�Beǡ�썣+��H�B4Ot���Op���O�d�O��?���E�`�8����U�3
d��b�Gϟl�I�d�ٴfy ��'�?��i[�'&黳��-������
�i2O�W웦�q��\|6�+?q�ȆD�ШB���3#7�#�윀r���H�O�9;J>�-O��O��d�OĽ `�����)��� ��E�g��OJ�ĩ<�'�i���<��柠�Oz��(�	�H�Ĥ� d�zX��O���'k|6MS��i�S��du�|B�I�Z��"�F6Q��	V'uSB�RS_!��4�P����ָ'?2�h��M�8�h�A�.x��	�'�^Dt�/ƺڂ� ?tI�	�S�~�-Дh"q�A��Q=�P
�e��5<��@�쟃�С��B�ncn���@NR�iX@���HvgĐd<��6错;� Q3�O�R�\� ��e��oP�yh�͹pT<"�̟E�V�Q�'��0��̛���4/���H�B ��A!"��*��Ap�,�8���f��[���,o��kf"O��g�F8�(0_XeX��S���pT&I�c��'v��f�7��ݫd�L�y �E8F�F��q�Ȳ ��k�� ��D�F�[�|��`�`�����N"r��4���Ŭ<a>�F��e�A�!��F|-�FDN&aI?:<z8H!E�bXlaH���-H(5*��.$���%"�K$�� �c�O\uP��� >�6q"D�K�9C6�9Å�O��d�O�,�@:Jy�nW���y[�IG��������X��#E�k���Jg��)�(O�<s��*�� �	�Y�"+$�r���T<E ���9P��a�'Ot�'r�D����?�O~����t�z�c^���´c�:��$K�����?E��'��	�-��`8��`��,�>`����'�'�����
Roâ:�&����O���D��P䊦o�m�R Y`+'4!��թ	<��!�1Bz<�ꡨǽ4!�C&��A��;W Q�pHߋz�!�$�2��|�Df��| ��J�AH�Z�!�d9�Z=K���bg��%��br!�$g��e��m�� L�9�4BƃXh!�$Y�f�T-�5���B�XZt�@�y�!��i���`1�Q�T��
C���,y!�T�{V��%/���P]PP��H!�D�7Ul�@���h����Lև!!�䕘6��B��Q�چс�AJ�r�!��4 Vl�$J(P�x;6�)=�!�ě�a�H�8P�%�9��$�x?!�d�/&�b�F���l��S7@�!��+ێ�(�NA�+"*Q�� �2r�!�d�Q��"U#H�a:(PoZ:9!�$D6~=�UJE�N% Q��՟;!�6NS*���	� �'�n�!�$T�r�p�ra@A���u�<&!�DQ�.o
��'�Z#'���׉�2�!��� �@��A
B9��-Q��|�!�$D<��y	d"F�b�^1"�m՘x�!򤃪q54����YXX��l��r!�ĝ�[�6��GBY��{�K b!�DZ%�X��_�8�x@�%��uK!���*N����(����cӶ28!�"z��Lyˎ��jd��O�_L!��?-h�D� [5G���V!�䃠��(z�SN
}S�f)R!�ď�{��S�'߳7J���Q�T M!�&>�$����
n*�U��O[d!��s�<�)��?t�l�ir��RL!�){z���n�;u�>��Z~�!�$M�17[Q��E��yұ�л�!��g�A��{��I�V�z 衇ȓL��air�O�E���Ƃ�4`�괆ȓJ=�!�*w�x)�JB�d��"O��bR!JZ��݁B%��g}t�KT"Ov����&��)���)���z�"Oh�wM�0�p!��u���(r"OL!	R@>R��a��f١��R�"OvL�7K�e0�����ߘXՊ�s�"O��%� =hV��U�nӪ�2�"O�}x���ј�cW�W�N�V��$"OR�ă��3`ٰ��W�N]�a"O�Ps��ϻT
�#
6`��m�V"O:ԃ0-� &���cJ���[�"Obm��a������#��BGJ�k4!�D��N;��h���)eF��b�>!�d�#"^ �B�B�B �͠���EG!�l���k��W�H̢I�'d�>?!�D��Ji`��Q\�,�QB�?.�!��C7'�8.)v`m�7IM6 ������ i!C$µu�p�n�30���"O��A�a[�F,,l�-C&�nyx"OB�0d��2HL�x3���eې�"O&M f�G0
8���.I�bl�q"O�xcGE�X$A��+�|�"O�ѣ�FG����Q�N-SC�q�"O�B"��@=�H!W#�+vEp"O~���X61���g_�"l��T"O�8I2�й_Z ���'˥����"O��Zu�h�挠��� LN-J"O:��чѧD�9�4i�#7�t��g"O>��C	}_26'Y�<%R�94"O��B��������ܪR��A�"OL���"�=p',ac�Ϗw.c�"O��!��8M�H��/#����"OR,ٗ�qIr��:E~0U��"O�+��"���bg�'5{�LJ�"O����n�S��qq�JE�MD��T"O��
'� 
�Xx)C%'�UI�"O�p���*3`�9Վ��.�Pl��"OD8���܇pI�`9�&��T��*�"O��Y�,���N��e/�g"O�yg"�/v�$�H�#]�*,d��"O|��p�Z�1!i�R��A>�y�"O(	榓�]3&�+rb82�"O��sVk� j�M��K^�K�j��u"O��!��r'��:3Ii����"O���Ǘz�A��s�^(�"O����o"*469 G�HXŪ��C"Oĭj�DI+!����'+�=�S"O���0��zڂ�Y��Y`�y"O�!���>^��)UD�_\]P�"Ob]��HV�+�\y�RC�]�։)"O
�fE$ }B�Ŧe���"�"O���5�V�?�,����Xئ�	 "O��2��������#��9��"O$)ht+�0Vs!���'=���A"OVy@oϦb$ ����A���"O�E�N�`� BfݿK�zE �"OP�A�'8Z�����	�$;PLB�"Oބ2��ԌPW�p8������"O��� �]�%�X�* (V!�@��D"OLb׹�V�ز@��*_�P��t�<A%���}{�ms����"i�4�]G�<9�/�2q���K_=b)x �fQo�<1�4a����ڒ!|�4��Q�<�LT�P,h�!bU�P�:�[��q�<	�	.XP�S��ňb�y�"��q�<a��ݒr�&)X��
�d��f�[l�<�I�7 :fa�k�8���ʑA�<���6N��Q�g��V}�`�+�{}�Rx��	���)a��FF�_�����%8�O������<�N�LѤ0�&mj+1�o�<qS�D�;	�-�DI�D@h(0�KZC�'�rHi�0�k�uc2�1*=
��� �2���O�����G��d$}�ek�.����N�i��O?�ɝDB%�� I(�:X�R�2"�JC�r�($K����
�2#/�0J�$��I�D;�@��$��#��lx��b�ߣRt�Ň�&v<�p���A	��$�\4 ���O���b�(@)*�!�92A�Ѹ'�J�D>�Hr�'IH��'��Ip�/Y!*��E��Oƃ��<ȶC �@=��D\��yr˔;1l`5��D�zH���jS�W7L��&�ņR/>�ZmE#)�M-F��é��9�����S�? ���Q��
/3j80�(�7 rg�i�JX�mV-ǰ>���(�$ً��:O���x�@K؞�Q�aǵR/p ��$��z����Dd~)b����w/v���S����c
�(�b��iH8EDx�	׃H&�����T�9�lyU �4;Sn�b��E�T!�䄑(�� ���L�H��+�l�N��b�/ �' �>���8�pv��~��(�c��*Z�zB�ɜ+~J���Ϩ]�]�Q��(BP6�_�`zZ��R�lCP`\2H�8���I@��%q�$?lO"1K ��d���~h}�1��0��q����7�^��ȓ�$�s��JzX)� -2B���?�AN�Z��H��I֜4�ԑ7'Z�M��L!�Cě�!�d�%/ND�,�$�l��C������թH��b�"~nZ��ҴB6��a�
	+�n�vC�	��`��=%^� ��j�L�@��+��'��xb��U6W�B�`��IM��u1�D\�d0OD���64����*5���r"O�-��/�;l�����!4�)��	�dm���):>@\�a�܄0��IBᏑOb!���u�<�&��?A���z��׬]�����p�=E��4�p�C�\H�I:��N:;�&��s/�x�ph	�K�E�G@]�#�U�'��[D!��=�0�ӗ:=zr�- ;���c�JX������u��6m�p�\��E.k~X��K��^�!��,&I<tXf뚾H��@�d�Iq��H�Ee�D��>���!��Rq�TKc��D�e�*D�<�U�76���ӵ�!.l�`a��tӪ���
LK�S��MKCE�4cBᲖ�l��)Q�Cg�<��Ы-�E #�^�^	�`�g�WN}r$(a6���d��U2QТM�8X@=z���)~4a}��3<��I.���e�Q� ����G;6B�<3ꜰ0&EG	:�i{�Oq�"=�!L�)�?�"�D�.@1C[�t֒��<D��I��J�5�<��Z�G�8T�C�d�4\����w�S��Ms�F	����B�_.Q�Xm���[�<I���-Sr��{ �. ��f�Uy2��p>yA�\�V<��KթH'9bA`D�PN�<iDh�c���#��L0lJ�UN�<A�nX�����*	(�}���J�<yG���'Lx�D�E|�lp@�_E�<�5bz����!b��{�����[�<����m�V)*hj(�S��S�<�Qn��6����'ԦN��Kf��L�<y�Ē�7��r�*�96�飰��l�<�`�ƨ!��I�愜��A�Ġi�<Ap���/�:���J\��xp��l�<�ҦȂ[F����	-[<�ي1̇e�<��f�l͚l8c���j¦?�B�	�nw���#�Y4U�2aCj�i��B�I3&�I$,
�-P���_�`&�C��8c2R��E��x���T!�C��0,-��ȿ4i�ZV�Y0`zC�Aih�@�G��BU���=@C�ɑ*`(�j>>Lr��?��B�I� p���+9�d�x�N�a�B�I��h�;��E<� ��&L��Y�6C�ɷ������( �I�C�	*n͸���e�	^&3C䉁?�b�r�o<!���� 7)לC�	�Yޚy�FK3e�l�h��`��B�I�i8��W�5=���;��B�I�U��Y�v�?A���HԤ��L�\B��`���JgIka4�Ǒ_!X"/$D��� �ϠVbR�gL@%Yܼ���/D��  ��nR5W$V�b��b.Љ��"O���a17U4 �0́�S%�	��"OPi��jY�W�<�d,�?~ZI�Q"O�`�-Ϟ �R��g+�5�@��"Ob4z�,I�U��4
�)Z�3@"OXM�1��X%Z��6� K�l�s�"O��ƒ3>�
���a��I�:��'"Ov$ ��2j���f(s���R�"O��Y�,ʙ�
,1�%�YkX�F"O ��'/̀���CϩR~i�#"O�Yڄ�ޘ\&�\Ygτ' ��sP"O&ܰ�
5Y]\��c"0�&@J*O�S������sV�1�`S�'��񩠄�3�1U���K��XJ�'A��0�*W<@� ���ِ@ 4�
�'ۆ�RO�1`����OH;᎘r
�'BYʴ���V������I,8�ƝS�'�^գr�[�k��Ea��ڢ&@��'�ڙ�D�2<���ϳ~2�!��'����F֟N�,�AY���K�'�R�!B��YD�k�i8~�V�C�'5�y���΂2��ᓢ�Vs1z���'[zDZ*��z49��4l��@P�'چ��g�#+VX�q�[�d����'m
�A�#�~Y�P��,1��`�'W���OA�J|h"��<�x��'͒�R�f 6'Yb��`Ç ���'%��IEOQ������V&��'Ȣ��g �4b8�	�	��}Q<���'8�����'�� J� ��@��X�'#�]s���|��Q�eEm�X=k�'�h̹!a�ڎ�C$�� TT�':���ʃ��,z�i�)i&���'�8��w	�>lܴ�C���̴��'�P\�e-JBg&�h�]:!����
�'�z%�S-S�H����s�ܸ
�'�2�Fn��'�&9�v� .�ab�'-�)S�N�Q�;A��-l�έ��'-´Ҷ�N.@�q`#�ؘ\��\3�'�q+���S�9+��T"?3\���'+n��iNb����8��(C�')�xpi_H�\�h�JP�/a ec�'
,� gV3A{&����(�$�Q�'5���˖8�vDQe�-ml��Y�'�8���"L�``Q�
�����'��2&�Y�2��{B�]�;p��'o���@�6!iQ����*���y	�'���b�# ,M�I0�����I	�'4Zy�AOP*L!z�C��N+9æ��'<�:6�TE u�&��
i�	�':�(g�B! ���R)�]!Ԣ	�'�"I����첢k�,�F���'ў��f�46A�[�&���j
�'A�8*gC�Vݦu
�ψ4#�<z
�',)��	(%)�(���t�9�	�'��XC��O�>	zU�O�X�`S�'$��23H�x��q�����v�����'�xY �#�+�"itO�$�@	��'V�]3�EE���������'���{��& �������"�A:�'�v�9r�
c`�0K����;�' p�AAǌM$��06G�=Z�'����`�pE��b�ŋ�'���	�'$e˓�S�i��%*�iZ���}���� I�F��&v�"�R�P#
�[�"Oj��nC��X�Q-D,u6Mp�"O��V�&���;����"O��R�l�b� ���#h����P"OԚTm�)=�@��bQ������"OP\��&�	]������L�$�D"OV="u��BRx��qC� �����"O ���aֵ���K!�Y�?��Ԛ�"O�@� �ʍRQ��yCAʎ�ĸ�"O�5Xp��_���Q͕�K��ՙ2"O�8��&ڋ��	P���cܤ`��"OJ���gUHD��p��Ы}��X��"O\���])X��-��c�F*a$"O����7
NLm* �_�/�(p1�"O:�!�'vH���l�(V,�4"O,���ۈ	5�pr�˅Mv,��B"O6�K�ʚ20[�l�-ɚG^�l:"O
@1�LD
J��h�U�R�ոd"O�9B��O��KӬ�&8Jص"O�=���L6D�B�"�N5����"Oܘ�@ ��P�N�"F�S"O�l�0N�"��9����I�1��"O$�s�@9jEBT�@�r!^���"OD�r%(T!Cv`u��hs����"O���H�r���P&�V1'�fi�&"O�a�Q��!zZLD��ǈ�A߾��"O|$��K8=�d���۔a���"O�	�#F�h׋�iqL��G"O���piX�R2�I�kÂ>il�0�"O$)Iq���!�/�CGt�JV"O�%#ծM�mBdXc��Qb����"OFk��N�WP� I`�/O�̊�"O��;p'�r�0(ʣ�
 ?@�p�"O��@L�"Q2�[�14��p"O�;3L��(�����:@�y�!"O(x�b��!%��l��0�y�r"O@�5圐i�<���L�;:VFA�P"O"��Sn��`((m	;<h, �"O���af�g�Эj��J�Y"l�"�"O�hT�\10Ą�ɂ��+#"O�l��0W$I�E��P2�"O��t��@�R�3���(��J"O���jLo-������74�,C�"OF(�UGaJX�!Ƣ�C�]r"O��YR�F6�
�i��B(�fd��"OB���cT4(��e9��9æ�w"O�Y.�1%��b"%D�N�Ľv"O���Ǝe�����CM'��H;P"O�i@��Ff��$BɳC�����"ON��ો�V��a2���T�Bh@�"Ot؄��W�yC������"OB�[�d�0 ;�92 �D�g�%��"O�2ri�I��i���oؔ�""O�i
�_��+��@� �|�jW"O
�{&�P1����V��
�0��"O�M	6#�*�N`0��2;�,�!"OtQ�Z/�6����
�Ŗ� �"O&�`1"��.i�gh6�fe) "ON��e�F'U�.�7�¨B��P�6"O������X͊5
C*Řw�40xP"Om9��+�Ui0�_�R�8��s"Of9SV(���-�!� |�"O��*d���P����qm�r��s"O�����4Pz,�r�oΌ��"O� �H���[�^��R�ΎF�!3W"O��Ѧ�;&�
�ٳ�(�����"O�́���P�����b�$�i4"OZd  ���&�9�����F"O��Z5t� ��۵62���"O~���'�uN�� Ê2M0�)�t�'��D��(��h�$ �O�r�=�ȓ;�$	aTd�V�4�PR�6��	��y�Z!�ܬ#R��R��?4"�}�ȓA�ָ-9 a���]�H����aJ4D��u%;\E:��CA]��-c�*O A�T���X�n���n�{���D"O��#6A�JNԥ�$`	�Iѐ��r"O��@���1��(q"�;V'��ا"Oj�:" �>e"͐�A�u
� ��"O�l�r#ʴ<�L1b�<_�	�"Oh	�I:6<f-i㠎�;��u�"O�-�T�Oo�i�f�Y����S"O|ܢ�ˌ5�~��u�ژf�e""O
pA���T�p ���6"O�����K�AA���dR�0g"O�����.���#�N]��r0�W"OFU���&�~�K�B�~Э��"O`T� �B�q �C�CK�"O�T+3)��|�U"M8[��-Y�"ON����.EcDq�
B��d��"O�0儋�R�TÁe�p�ޭS�"O� ;���f�$� ���c���X�"O$H�C��A��U�BM��/N�T�"OJ91$ܤ	��X�ۿD8�x�"O4P9'k�G�������MJN�`"O�IiFg�;D��d�`G�}��"O��@��Ne�%"ǡU
M�*D�Q"O����B����a�����w"O��" = L�Kp/E20��"OVԓ�I�|P�=�)_�Q��"O����Ίd�� TB
:fni�"Oֵ����@�^̸g�@��h"O���CBT�M� �����"O�!�MX-P�fPr�^]�k�"O���D-2rc�V��T��"O��k\/���
�k �5Kd"O��a$��>ܡ���%T��"O�q��b�b�nm�w�[B�4��"ODmQ
������� Q
�I�"Oڬ��@V.`���
T�9�I�@"O��9��\[&@��R�T�D"O^�y�]�+@��A�;Y�0�B"O($�#շqæt���܇��y��"O2aԩ9� 8��BÑ �~���"O���a��Da:�h�n~���D"OxB2��!@������"nl,y�"O� ��n'A|&�BP��P_\�rS"O��>y�bG_>S"��"O*@q"I�l3���#��?I�#"O���R���`��	�m�F��"O��	��̑�nА�핳M5*$�"O����ڦR@m��˕Y n��"O8��`I/M����*��jT@$"O�1�E��d	�
4�J,W�H�+3"Op�P�ˬ�ܘh&��&>�(��"OP�Zq	�Sb;�抣e6&�U"On��g�K�j�BE�P��7��J"O&��螂(�J@/���p���"O� �s���v�F��4�i�<�cD"O�I�$�!0��Q�#G݄}�&�#"OQP#֑��y;�^��:�h"O��[���d}Ԕ��>,$��5"OB):_2L�!��_!:>�0i�]��yr�4͈U����(�l�w�Z?�y��@ld��0拷�쩓VjP�y`����Ҽo��정��$3��	�ȓ"B���R�%"�H���L���ȓ,{r`�3����t`X��_8��ȓ��@cA� �X�w��;�l��ȓdx]p%�C�uH 8�I�b�х� ߆0;AGQ�t�:t҂*R�B����5Z'AV�&d����K7Ji�ȓ˰!�IW��l�Qj7�^Ɇ�b�D�l�!((�֤\
��ȓc��U@�G�t����T�$���m�(!��$C �L��%��(�9�ȓ.�T������`)������ȓ��S�gU9��H�&��[�x�ȓ6̨�cង���Q7-�k}4���POZW�6)F ���F)xp"O���D)BtH��aID�� �q�"O����k�Z	��u)�#j稬82"OR�y�F%S����t� ���"O��p�=c1���ǈ�^����"O޼��-*�� ҡ���\���"OZ���ָU�^�� �ȟ(��͊�"O䰊$j@.K� �ׅ�$�|��"OD�Dm��U��d�#�0�w"O\�`'L��{H�Y�գ�?�Q�"On�Q��؂Y$<�h���;:mA�"Oq�3����}��- �"O~�	@����Lb G�*e~l��3"O���rd�D �{@�P�� P"O*A��OȥoX:�"Q3���C�"O�J�r�X�2�O�����"O$$c��_9>T@��:��4��"O�=��qk������ 8/L�Z"OF��Q�.~�6�!WԌ9(ܼ:a"O&%!����|M"lJD�ۦ$P�T"OjĩE$.A���ظL��|�@"OT|��9MR�b"c��E=L�+�"O�H�񮓯6��H��E;̹B"O�@1�ޚ(��9@,�S'N5��"O���e�9F�ܤS�JX"^�ٻa*O�Y1T	�Kba
���}��y)	�'w�Tѣ�D?8]ڭ�S��<�ޑ��'f"�Ig/њtb-1$E�np\m�
�'&��s ��#w(�f�S�_���	�'d���cԋA��j60T7	C	�'.�C֕B٢������FrB		�'����.�2�r�dK.>���Q�'����6Nͮw�x���S%v��2�'b �����)A��a�NIG�)��'ly�%�ͅs줼S�n�	b�8�'����*)����+�$K	z@��'���H�+�.��8 TI��B6!q�'��@�+<7\��-%A(,E{�'���q�œ?BG����8����'���#��ݵ{�H=+p�X�B���x�'���@�u)���@΃DJ�q�'�j�!C�yG�a[�셞B�ȩ��'���@�ɢL�QcQ\B���S��� �E�$D�yj`�Bc��(xx��{T"OX��a��=3>�)��R!No(��"O@�x��2������MW�@��"O��[�Cѡ}@Uk�$n>T�"O�l@�O��P�����vak "OH��V�c,�c��h��y�"O�CP��c��4�;#���`�"OD���R9"nB��w떈Y|:8�&"O�b�������Z` x�e"O�a2���Y�T�CҨ�!ET��3"O����\����-h1��b�"O�d��	�.�dd�m�
�*p"O�`����tۤ-&�C
�����"O�}���8<pAx ��F�D�6"O440��]3C� GD��3�|�5"O�����DIP��`��d"O��YW��l�a�T�.�xYې"O�����T	�e�3��&\Tlp¥"O4��ꃪn��@�B�F����"O�-�r�W�4������K	1^��z�"O|(�fm��V�6AW�0%4�%"O�R3������!ǰxӈE�c"O������
�z�ՠ�&�F�#"Oj�bs� U�x��o�~��x��"O,�"���>@�$����� ~~e+"O�9�^:(�b�Va3zY��#�"Ob 3eτ�	� a�t�<K$(qQ"O���p K7Z��H�5C��2DT"O��� �E�_R���X6{���X4"OP�+�j]3X*
�`��3��4��"Oh�i]�M���WFP�q�d��"O��B*�)�\�H�l�hH�"O��fhϮ*>,p� <am�5p�"OʱӅ�V'i��J�O�_V�T �"O����2Z|�K � �[�@ �""O2�SƬ�I��`��O�O����7"OfL�UB�%Q�:@1�b@�+����s"O�	*�MVj�q��׋j�޴�@"O�=�e� b��1���_����"O�=��,�%�
�C͂�_��1c"Ot�@`�H���Dk�
�Y""O!12��{����I�y�8��"Or�b�F'uK��qۓh s4��ȓk�����7x���9dN�r
&$�ȓ@)��pm�;���%�г.;~��ȓjhm9�HU�D��Ap�/T��8��ȓr<���ä��F��Y�`e�zهȓ/0��sa�Ia�Qn;ꅇ�&4��(7&M@�	qe�M2*$ҽ��|��}�G��&�z)���O�*��ȓ����9-�)�RŖ=E�r�ȓi�J����o�й�A� �g$��ȓ<$��b��3?`ģ���2#EDՄȓN�B�[��+"��}SU�׬��ȓCe�[G�:]]6�9�_�c\|����BcO�>etT9j���!UVh��#3UA�#�63^<4�H��ȓj��<��@7/8��i��Zk�����a����1LB�m�#$��-f�`������2���`k�9����Ĥ��z"���.а*u���AB������W�L�z�MĆ\ڂ))�-P<Gt��ȓ�����Ȝ�7D�u���� ��@rL3�O	�)�,����Z�D����S�? �4�El^%��1�5�K�
���e"Ojt�7A�3W�<��!�;z�Ѳ"OJ��'B\��i11*�2K��"&"O6�k(^��lC�iY�wH��y��E�D���K�V�"�1D�·�y2N_�B�L(�í[G�,ȓ�'�yR�0�p���DU.	|d&A���yR���P�z�z&�S"}�r�b堆�y".�v��Hۧ�ֺa�]sD@G]�<�al2�ꈚ���.)�]ҥ�}�<�h̰/A��/��p׊��W��a�<���U��h�G�	�t���5��t�<�j�=~J\,�A�Ğ�j4�Wlp�<�d瞽"��#R�v`���p�<�Uf�.>0�B�6^܉�NS�<)`L���z`�Γ[(L�+�Q�<a��	��lɷ%�n0���`NO�<y3�M�i��h塌����eEO�<!�Ay��8���?M�;a!s�<!S!eȆ3���2u�EH�<q#�'LCT�PSU�|�l9��N@�<�VO��ZTȄc�~8Șb��u�<�E�j�����z��0t��t�<᳉S�W��D���]�B=���m�<PB�']Vii�eƉ)�d��c�<Q%1Z����^�t�����A	E�<�w� )�x�	���`*�H�d��e�<�&S2��8ɐkK��4hRi^�<��@��N�t�Cϖ�f4(A�$S�<yeK�Jn6e�o��a�N5��*�t�<�sg�=c�`�'��c�=a�o�<�%�3y�*-�Dτ�6����#��l�<��-C�>Q�JX�n��]�3 �s�<�ӌ�#�P� ��I�tlj�kHU�<a�Ӽp�ذ+��@�1�萫Ӂ�M�<A���O���DD^�v���e�o�<��i%~.�`�ǋ�4{bPk���g�<�v�G8ze:�b���h_^�(�_I�<I���8Z!�ѤX�`+n8xdF�<�P�Q��2����M/��1��-VI�<�nƌ&����큈G� @�Z}�<�7���`9��ˡfQ0+ʰS%B�{�<�1o�D�U�s���P9�9{�k�v�<A�I��8hZh�$��X̮���)WX�<1RK��l���Z2�K�̈���Q�<�⋕{����U��c�:9���U�<y҄�=th�!j�fW��F�`4D�O�<�W�P$b$ք^����aV�^I�<�7�G�*�<0a)�)pnY�BO�D�<��I�6j8t��3J�2�����@�<�3�Bj�zͲ����*M��Dh�~�<)6�" �V��"-ON�!�À|�<YSN�>�V��	ؐ`5>�q�kSz�<��(X�Kyl��ve�"�F�+��vx���'LD+1B���a2U��i��d%O���u�~R�"�ܞ����"O ���A[>��X`�DK�{�La��"O�A7C��}�D���D	U�� ��"Ol��� o|����B�R�|T@�"OВ���3ZJ�h���7x�x��"O&��m��c&Nb�� �"O� 8��� (j�|Ç䒽pC�d(�"O�P)�l\��J��7ߠf���8S"O�,���!���a��3 �LI�"O� ��*w`з,�Ā:�D}�
���"O����Nɼl�������E��S0"O��b OԿ4���a��܆&��9��"O��p� �w[�`��fҼS��=��"O����I��$	h%�랖D~���%"O|�X� ΰZ�� �C
jN؂7"O�9�
S=k����d*�Ch�|P�"On�y���3B�P�Hu��}(��"O~���)œx�.q[�	E�m�"OY8��	,J��PfߋX�e��"O�u��H�(��a�ܳ��("O(�!�&�6�3$�0i�؀��"O����$\���t���;�"O8�ã�+|�L�*���g�2�
�"O@a�vHc|�dC3��|�h�S "O���6![�g삡�$�&���"O���'D_� �WD0A!��z�"OD8�1�Q�!,�TB�$<�L��"O,��^�K��L8�&O�B�09"O~i0D�"�ZX�ͬ%��$�w"Oj�R�k_�
]y��X�U��0�"O��R��9x�t���mI!I���U"ONA[%iEo��t����F�0e�t"O��4��uD��	8*�Ќ+�"O8xp�G�^��uږ�\#�*�J�"O�<kQ�ǒ&����A.^����"O��@4�Z41F��p@R P ]� "O�0J�$��f*T�ϓ.Cab�S"Oz�P��� wΪ��mΝ����"O����ʰ;2�ē��I�߼�1�"O
0��D�5��������c0`��"O���g�dNԴ	0��F'D|�"O��C'��su"�B�Ȑ>E�}���D(LO�YQ#@�	R`���OL�~��pI2"O����\3$I�yXh�f"O>�86��L��xKfΔ�_Z ��"O��p��||<���9iC~�S�"O4��I��"$��l�>O*��� "O21�P(8�rt�LҰ5z�A"O��A"�Y�T��@ ��-qX@Qw"O����홻%�Α)�(�̄$#"O�	� � �BZ�g��d%
�"O�Y�
�8b`XR�o����!��"Oꉺ���BC:IN���uH��|�!�$���`u����={B�h:���!��ğ��q�.T".�=��'_vz�y��'�1O��p�� /�U�5�?pQ���"O,�**��l# �85�I�(J�k'"O�d�D�m7p�����O=D�)g"ODLi��ЗA��UJ�8_�ԡ �"O􈈆!�@�V�����y��"O�LS��J]b���f�lp��I�"O�Jq	�.i�r�`��n=�I矰�	çrwR�Z�!�i[���G"Ht�ȓ]T���\�"�T%#�E]�^h��*�~%��H1DD�q�Ӌ���ȓ?���TJ(
�.�Ag��+�ʐ�ȓI&���C+|���x�$ɉ�p��ȓC@`R��}�"�
 �̯J`��ȓIW��7�LY-��{SL�@�0��NNl�j��2G��	q!I �t��Wԍ���?ٴ4`�%��!��ȓt��k�cUv���OU0�z���}oj�"�拍��S��Lc/Ć�S�? l��5�\?�!J`HYgܽ�"O>% �b|���  IN��"O.���п7҄�SL[8 />�q&"Ox%A�#κ'e�]��N.X&�m�"O0GD�.�t}hւ,X�+�"O< �s�W)�جw��k`b��'"Ou2�o[�\�D)�gU
\U�� "O�Hx�ϋ!V�N�B2G^�{��v"O� R�c��{��P��&U4��"OƝ٠"U,I@ �PB1n+���s"O�����	/6�;�B	_"|��"O��U��,�	إ��9�T�0"O`�S �Bs8���DJA(�"O�e���B�m��|��@�y�n��w"O:�����
.����!J�ē5"O�TA���$�|�*BׄAН�"O��ub�R0�};�@C'�b��"Ov`"�,C�h���@���Je��T"O�<If���%0$X,W�`�)�"O�y{�/�Nr��A<y��t��"OTH���=�l�ʦ8���z`"O�����%�Z� >9ҒU�g"O>�Z�Ǝ�W��@���:�B�2B"O�q�5�[
~�l�o��a�i�"O�P�ii�J��-�t��I��"O2�b��]t��X���M�W"O�6�P�k���z� � h�~���"O�d(	??aDٳ�P>Y�>a��"O��X���(�lh��،s����"O&�vI`; ���"ĥy>�m�"O\����[��<��!ޮN/0��%"Ot�4�/}t�z�� W�HI�4"Ota�s@͔=R�	Ǭ˨#�$�j�"O:�q�횋P�E�ԋO�S5V���"O�t�����Q8�%`*O b���"O��kM��0���2S��0la�|��"O�9J	޷T�
���ac�i��"O
��e��G�ةq���2va\T�"O�Lx�N%t�D0#�֚"�(�"O�,�C�0����b�,I���"O<�āU�A'0�:Adçy�`��p"O2�aɂ�^��[f۷NYf�i�"OȰ��$O�<ĔAS���-��u�g"O�,�B�)�2R#�.��hiw"O�������)�7�U5-��Å\�T�IK�S�O��\@� dB��qgX@+.%`�'���`��оRi�8Х,�=�2uK�'6�=b Nؒh�E��O@��;�'C��bBN�T����\i�'����,�Z����#M��6ܢ�'5����A�.7ɰycE h�|8�'�RAGӏނ	�2�ŚtQ��Z/O@��)�)ʧ�B���ΧYT�\���]1�\��`�L�¢
*(�)��#!�\����Ar&K>C�f0Ɂ��8a��ȓ2�(9w�D3mvI�]�UxL��ȓ7��X�e�.����3O�J�d��ȓ 醨��))}�� b�#4�ȓ|d
2�ġ:L\d�t#�$t��a�����1Vz�@ �I�g;�|�� ���j����Z�.�#���)���0��I�5C�T�S���i�l���.�X@�򇉅n�N��e��%je"T��\����:�� ��"byj%��S�? �y0��]�N���Y��3jq����"O��p��p��pJTA)k@����"Oa�	[�L����t�� \949`'"O%�C21Ը�Ue�8s���"O昀� �i�`h���!H
�"O��i6!)ekL�F�Ն)��
�"O$}�512��C�X�x�"O0	g�<~n���`������'o^��Rl	�<�݈��Z�ER$�'Ђ�Z2�� %��T���U';Ҭ|�
�'�t�ä���P@^�9�
��g�2�:�'�6�P��W������oM�S���'5j\: '�6[\��q@�$��Q
�'8��*EC�#��ps�,��t�U0
�'d�esv#�R*
�1/��a����	�'� 0�	�<Q��a�0h:	{
�'Gb��U����|%i�	ۦg�e�	�'X��+X�jy)��C�k���G��`�<�q&��|�d��̄/ar��w�`�<��0��@��,EK�q��I�Y�<&B��6EtM:3��#u�X}�֭�O�<ɗ��8V��BL��}*ZQ �g�<I4˕�>�`� V�V9�eA�^�<�e-td�(�7��^R~$��+b�<!�9�J���R/k����/�u�<q�gȣg��Z��7��{�TG�<!$M� )J��7�LZ8�q�Jh�<Y��m���郞��u��m�< dY
.���՛v��"���`�<���T�k��xVd�C=h�z���[�<Q5�
6-~B�&����dB5�DP�<	�L���p���_@��r'&
u�<Y"O��'�p��ǖ@�䙥��i�<q���VQ��C!7�v�Y�UJ�<��U�j��J���b�(؋#@I�<���P]�ڔ*��ܲEQh\e�Nx��'?,�(A0�P����L�t��	�'�:(!�*1�^]���L�3 ^H*�'d��j�%�	-�d��p �~���'� ����\�ntc��_6�L�
�'�@�!�d��	�4�i'�F8.�F���'t��%�A!~�J�f*�= >��	�'{���,Y�?�P��2m����t�	���'q�}��-U�{�Z� �jQ��:	�'e<	����%>��������'���R�ѺH�r٣R���߂���'$�+���"K���pO�#un`��'��쁣��
K�2Q����!V����'p�y��B�3d�-��%�* "�xi�'�%Y'h�(@���kR����бr����F&L���qf˚M@l�b	�I�!�d�>w/.�㔦J�tD6�"�d�L�!�@e�Y���8�1��
�g�!�d�Q �%������g�&_[!�$[�9t���_8i�V	��b� 1!�qt�4:TW�U}^�
�AG,# !�<, Q%@�@l�����F�]k!�A!��	�a��wX�m$ �`!�d�SH��3�o�)BFpcc�݌Q!�d0g�QX��@�E�Y��o�?H�!�$�#"�2�ISbB�u�,8�h�%T�!�W�A/�=��مg�j��:&�!�i�jYZ�D�� ����B5�!��Օwa6��2�C�V�z䇔�5�!�� �᳗b��5ߒ0!��	�HQb�"O�-�C��;J^Y��	�6uԴ��|��'`az2݋v,�(j`L#S)p��"`��yr�Q�:���H���`�1�F���ybg�L��Q`��]��0�@�yB�."q�[��A-���k�i��y�ᗃz�%D��y��Q�:�y�ʂ8621��J�=qo�)������OT"~b2���K���"e�,v7LP8RC�K���0=�di�:Pڈ	�"פO�HX�g�G�<q���^4�� ��"���P�B�<�!I�P�8���5x����z�<����r�`�u�H�H�@Tq�<�M˕R1�9C�냒QK��v�R�<q�,:(l�h� �3��0p��IJ��?�	�'6��ɰ��B 56\�^�VA�u�ȓ��h)�EX�k���k��H:l����Q��ab&g�HR<�9@@�l{PU��z�P��J�W�8��c�<@�z���J%`������(����|���ȓA2ĉQ�>&�pR��2�:9��a̓2�B��n��^`�Y�Bl��s���G"�S

��4�֛�Nu��!0ԨC��4A��bG<k?}S��Ò;��C�Ʉ����hU�`�1�6�O��JB��<U���Zf#��)JDK E��
�FB�I�zx�} ��(5v�hn	�c�0B�ɸP�$i���@4A@�j3�\W�ȣ?q��)Zݶ5`��� xr��v&�"�ў\��	�h��@��"��e��Y��H�C�I �ιc�E�K&�� �K7 TLC�I/�␙EH 7L��U�E,N91 C�I8g�ʀ�+n8�%JᏜ�C��2A����w+��G<��iwꎲL$C�I <>�� ��ɿ]R��gE�����d*�)wHh #(��#�8}�"���4B��H !&�����4#�@'��F{���G��U�
e�DBG�������yr��L%��j�W�y�t`���ybAA�.���9C,6�x���OX7�y"�@0\$4������&FB�Q��y�&@j������JG�$B��S��yRf]�l��j��F�@# 9䎏��y�)F-(E�Wh�9d�RC˝0�y2��m`�i��s��1�@ŜpI!����Х2��P�V�����I1!�Ğ0L���A��޼>��qR��#00!��&:b�Kdș�l�8,r�&ײ*!���]U�u���� 
u2L���; q!򤟦j�F)�4k	�+c��g#I�:�!��P�pi�a!�*U^�ab�*�!�DǑP��(qb��o:������~x!�$ԭA�R�z���@1��ի�rh!�D
�\�D�!��*�Ä�
]!�d��aͨ9�����F�I�Ĥ�(p!�d�=�vթ��d' ���eD!�D��=���#���rg�}�g�!�$�'s�ࠃ-H8v�%���!�
*&�4��k��a�@�;!�$#p��0hС,w\���b�5�!�$؈��D[R)��|S��^!�D�^FҥJ�Ê*"T��.� .�!�$X�t�L���iǷR"dU��ݖ{!��DRm �h��jb�\R�� t�!�� F��eG�]��+r�P�BߺQ1�|r�)��;9C|eb����}Ė1B�N�=Pq�B䉡;L~�Kw�Ʌ$����&U�b�rC䉍>�4ɑ�b�h�A�D�h8>C�.6ta@�8W(��2.TD�JB䉳OW0a��O۩b�I��b��H}�C䉬,�%���_ݞ��Ev�C�	�
�n��%#%W��sD����B�	�>�~ɓT���,����H*B�	;��4��1QɢȰaKD�2�bC�	�@|d8b���M�dI� ��B�I���Ű��@�i�((�%!��_HC��> ��`c`�v�(|��e�?@�dC�Ɉ>2|�A���-W�8S��G,Z C�	�1W�0$퍫]]D�d�<;hC�I�_��8UK'Z9\!�w쑝Q��B䉒,M:����O�Y-D�d�B��� ɝ���E(�p�!�"O ܓ2��,Nɮ�	�f���Ca"O������6�L�#��o�ʵ�T"O�:� L�s���9Ab��v�"O`���e(Ǣ ���Y�#%���"O*�����p<x Y���!��`"O��CM�R�.mbBBW~826"O�Up�(��
1 ų�(zYj�٧"O��!��q������qQ��'"O�#��J(lb�j�)?=x@"Oj��GhO����J�wN�Y�"O�d ���+��ݪ���vM��h3"O�%hf���5�6D��M_�>���Kf"O�YKV�-4�Z|a@ύ(%���`#"O�Z�Æ5�pq �����L��y�N�&n��hs�Y�5@00���!�yR%o�U����.��h�Ȕ��yb F���P�X/Q�*�RC���yR�O�ѣߵ7m���n	�?��ȓj�l�۶�?z��}k&ÒGP��ȓ�|��$��5V�I��N�P-�܅ȓ7�*��(�i��튑˓3+¸��ȓsن8��׆G����E΃-�<5�ȓ�|�)�#�R�"!д�]�f�4��ȓ4��3�-�B�}1�ȜHVDH���t���A],�$=c�ѠS�Ņȓ#��Y���I�NRTc����fQN-�ȓ^�b�	�lQ%<�"��p��E�d�ȓE ��
��XP'V�q2� 9x5�����l_&=a�t�ӱn�0ͅȓn{����C��$C�
!���ȓ�T{�瑒2�l��.60\�ȓjt|�gP5
�����pS�p�ȓ)��P����]3�@nRY�ȓ��@���;J�0;#��/hB��ȓ4ƜeK����/�4��Ƣڭf}!�d�20:�k�F�[����E��/!�B�kq"5*����(�@yZ�KM�!򄈱�$�JP�ݯhu�al�	!�d�9mԖ;oO��eHG*	16�!���.-�m�L�$& ��)_�*�!���=,qn�����{|��G�ڟi!�$ܫ,u8�:b�Ѿ���P"�,-!�ǌ�
I�7��<|�4��Вtm!�,:�*qm٧/�|��ʞc!�ɇ;�ҕ+"� B�8Hҩ�<a!��(V�BŨS��X��C��!�� �Ũ�kɚ+b���6�Ӡ8M<MYW"O@-�Eh��GKv9�rG�2נ���"O��i�A�~H�po�����U"O�	���U�� [�+��<��#"OJ���B�x���j�
v�,a3"O�@�D@؎h��p��RchP�@�"O��w�Eb�xDk�K��;^raH�"O9�S��TՖus�HB�~'�u;s"O��kpH�(<8�ၰ�]�I!�I�&"O8-�嬅d_&I"�e��8���Q"O�,[%	� �!�V���H�x�"ON�c�	�vt�aI�0F�p�4"Or�#v�ӸVa�h��4-��P"O��ÀFO7j�qJa��C"`��6"O�\��I�5�~�� H#C�d �"OD5)�(C#a�J�Z�'��{IV1a"O(Y�Ƣ�5b"�e(� `���"OZ�SKX�Z�L�a��Wۖ"O��Վ��!.�"v��=~��Y#"O���G���X*w�3n7\��T"O��B���72h�]��)��J��k"O��ӲSt�&	��(
�cb"O �Y����L�"I�3�^�S�d�QQ"OBM�Ph���)r�ֳ%-|�P$"O���Q��r0Ec��� �|@"O��p�o�!F��Q��["d��"O��sda��%5~�`U,iV��z�"O:	�Ɗ�8�dI�#f����("O
�	���PW
�2a�2��$"OH�J��
3����hI7O����"O�m��LtP�Q�Ι�Ol,�&"O*@� *��@��y��5�"O&�#���u��Y��?�:��"OސZ�I�8=�ԐR1S�c��I�"OJ-r�䇓HV��S�(����[�"OL9�J	�<���sG�$�0x�"OV�@�d��4p�#���hն��D"OPq֬B�G
��T��I-�	Y�"OF�"� �5r�b���fܬӷ"OĴ+$F�f�*B�T�M��z�"OzyX�遛b��+u�����"O�T{�O� ����G1Wt0�"OzH(`�'xl)��_�n>��#"Od��!�3�0�� g��u*��[S"OhI"� #D�p91���h�1ZW"On���V�r�d��hȝ(�vT�"O�]�4��X�,���fٝ~�Dܘ�"O��y��ٿ#.t|ʧˊ;*T:�:"OL�C��,�LT�mְgO��"O��4d���M��,Ǻ2O\Y��"O����W ,D��
C�s���+�"O� ��,DE\d���JT����"O���dE� p ��V��3r5��'U����H�\"8�W焊G.�"�'��;զ� qu.��Z�j�6a��']�E�#�I�h�<qc�� ?\M��'�v�wr��[�a�-B��e��'�V�)�咇�L�iT8<*�Ը�'$f�A򨃤y׬EA��1-��L��'H*�k�j�2Cl8�ʐl��+����'����P N!�00�*Y�[	�'!��8��
/`��2�� :M���'匕�. ����-"R.��"O¨r�'8b@�y��Ǒ
o)�e"O�  �8���a��m�fm��&Er���"O����e�z���8>jZR"O�P��k��t��cf׉G�x��"O$ �g,E5/N���E� ax�"O�Ay"�B�gߞ�sd��RE�@A"O����J��<�h�JtC0JC�Hk "O�T�`E�S�4�b��S>H3a"O�}�� T�D��騐����M���"D��C�`2K������`���3D��ƏZ��H���G�����*3D��4AŏJ�"P�H��K
�Qx4�2D�����/�
Q������B��/D�|����P��e�Z-@g��h �/D��e.ڵh��LcF�� G�4i�f�-D�(y�OZ8<�zq�U#�$��1D���� 12�\�k�`Q(���e,D�$���8z���a�S
����(D���l�|3fK��l[�Hj��!D�����R^¶���%> �����#D���qkA�ل�C�(M1�$����7D�@�#�8q��,
7��:M�����/9D� �5���]���pǆah��9�j7D������%"�̹7�Q]xHqAIb�<�C��4KO����	ژh��嘥�IX�<�dK��d,��tǜQT�MТ�K�<��"Q�l��8fbN�{ɂ��cŖI�<Ag��������ܾ!O�aA1dC�<��fJ9����*��I� !@�A�<���3�xx���]��]� ��t�<��KM�=n	(��X4�셁D��m�<���A?p���8�������`�FA�<��)N�V�nY( ��;H�`Q	�A|�<��סFDv��@!�Y�||q�)t�<���#$WH�PԎZ7w"�9�t��m�<�1d��[z��33��3 ��1��Z_�<i"�Ȗx�bݢ�hX�'>� ��^�<	4N�n.���[�0�3��Z�<y�[58�p0��_�:��SG�Z�<釉*k��ɓH��8\AYcG�X�<1�@~,ze{�Q�Dw �j5�X�<���ԪNS�0� ��&,��i*p�RQ�<���9Ąl��`	";2���b�<���-�*ɂ��8�(��Da�<���V:v�N"���\���`�r�<Q��U�=@!�R/�G1T<��cIo�<�SfX1_�t��$�!��aE-Hl�<yA��2"�h]�Sh���ܙз�A�<A($E�JT�6���9>�Ҩ�t�<9�!�0Ĭ���}%�蔌Ae�<p$�(taPo�WR�YHԯ�c�<q�j��?]d�!@��8�#��Ut�<QuCM/xn�:����B׸ZrBنȓ4A�¯T�$E��Gɝ���ц�=�����m����F�%*��݇�i��A��HE����b�j}��S�������HT�֖�<�ȓ�X}ÄK�.��V�ۑ ����ȓa�B���i	�z��ro��\&���ȓ��\@�ΐK��岷�P����ȓ@�~-��%P��Ja�R%�"���J+ � �\�6��cI 3x ń�L����L�#�&� ֹb�&�ȓm���Q(�7y��<�Ңa!2kKG�<!���ް���ܸa�rQ
��<� L�3��\�N�6�0���
@�*���"O�\	��T!'wv=�6�S�-甬��"O���T<B���$I;ֲ��"O�qQ����.�4 �Ï�K�=C"O��S a]�`}�QJ������"O�}�qg��H��t�#m^5k�F�Q"Oh�86C+%B��*BϳYE<0��"O`hHa�F+M��G��� >rX"O��y�,rI�.�'6,�B�"OPu��G&��{�C����"O�8R��< ���C /��&�T�`""O��JtL�QJ���sC�i�B��"O���F!DV��1)�!A3i��
�"O\�`5䔉S��d�b��A�t�Z"O`D�s�  �<�#Qg*��"O�}���C�OϞ���AF
\T�aP�"O�:iƲi��˳.[�L��\Z�"O,����
U_�di D,�άZ0"O41{7��=h��\�v��+M�����"O����'ބX*:l�R@7nLMB�"O���P�#"�pCD.O�@�az�"Ok�*�T ���,�(`� �"O�0S�쀑*���l�)!��3F"O@}:�����(�j�"�X��"OZ�{n
'?�D��3�:���z"On��T�X�M��<�2�H*�ZA� "O\T(&��OA��îP�sr��8""O��	P�Ln"J\���> ~�L�!"O��j�WfT4 �/�Cw���"O��	h�d�d��\q@��"Ov�{�l��б��o´e"O���)X�G,d��&�ΟCC�i	�"O� :RO�@_,q�Ǌ)d#*�Ї"Ojh��Ę��M�G�;��ӕ"O��r��l6��@O,�� �"O
LP��e�<D@��O�I:6�"O45Ѕ,g�	�1@\! ��� "O�@yU&
=�H�6	C%-�ŉ�"O�P�M�8 (�k��L�G����yB 	�{��k&n�>i�ⳇ���yL:Q�V�X�M)`�@����8�y��\+%�\���]A�q9Gj΍�y�/���>4`#.�V�����n�'�y�aĘx�����B�K^b}���y�MG<l��ٺ����7 ���ì�yB.S�"`~m�2�A�'^h(B��y�c�Jp �V�ܣ@�)�w`Q�y�˓X�|�`*i囶D\�y2+����`kC�HfB(�	?�y�cͷSF���$B�\�������y"hZs��86G�4Qh�$(6��y���2%1ܵYV��Q��p���y�D�PY��1q�F:r0���ǋ ��yr��pv�`�G�ΘcH�j���y�n�+����_�	�V�CF�Ȱ�y��4y\!��/�t 􀸶�ِ�y��V!+,���M(�j�UHO��yR�2�ޙ����M��0(O��yr�ɥn0�2 �ģ%6 �CJ�y�I��P�yO��V�@�P��y�ؖ6�je����V�V�IQ��?�yr�S%{�x���Fz̈��C��8�y"F'F<�d��	ۛx��+�Ɛ��yBoW��ָj ��s��Њ��[��y
� �9A���lm(�"R�75�V"O���b�
\�e!���/2���"O P�2��3������y0 ��D"O�J��U>/N���2,T��c"OB0"|P�8�I�$�����"O.�#%L9y쑢�a�x�� p�"O"u�"	�W��qb�5f���""O �Y)P</�\���}`U�B"OT�p$Ӯ$T���Hp]�I�7"OB�2U(�/3	t�1g(��L�j"OĄp�GN%���7�˟i�(�"O�dQ�\�D�P$8���&DX�0"ON`���ȈR�l%���q��� "Oੁ���%'���jg-��z~�s"O�{Ť�.+bR���KN	�\�
�"O���`�ܠ���{Ɗ��z�|�;g"O��C��;a���ĩT��8�"O��ZNV�IE�u�%�{{4�@"O����!��K���7@Y�0��"Ot��gM���9cK�J����"Or�#��V$��8;q�V�}��0�"O��&�Ӫ}5��@C����"O�qɢ+��f��t��*x�Q�"O:ɚ��W*o&�!8!�Nr^� "O&��1���&�����4�>��"Ot�A���BA"�3�6A�P�"O�嫓A�[�������s�T�a!"O�$v`P�Fm�`.������"ONi��j˧y�Vŉ0(�Q��p�"OҔ�1?hd��'H�&v�>��"Oր�F��Z�z�S�蝰0���C�"O�)���eu��*��|�bT"O^��1�[>Z�X���*P���Ec`"O�`���JL�� 8n��L a"O�<�F���F���j�3�(�!"O���AG^�Wc�ˡIǊ6�h	�2"O&AP��
.mP�9 k^�t�5��"O�%�����[;~490����z-�g"O��cqA�p$�8'`�=,����P"O��`�T�=~~�#�nWC�DP�"Ox"�Ƴ&�RkI� ��U�7"O|H��	�	:�t�8SJ<~|yb�"O�p��4,Y(,@�	���is�"O^��6�I-�b��k�}��	� "ObyQ-S2�$M�$
S,���0"OD����u�Р 	� Y����"O�@Q�NݮQ�ҡ��D�B��<�"O$��ڸ|}�Y	Ą�	c�p
�"Ovc�Z�l~�	w�E�Z��"O��fa׺n\��P� 
4O�a��"Ob!K�����\4�y$y��"O>��W�(6P-0�ȊA#x�f"O��z5O��[�����Q�D+S"O��b��w�y1�/� �@���"OH� э~��Y�Go�?^@���"O�!Aō�O↼��]�r��"O"{��&�`���];(7�՘�"O�A�@��s�j� �_A�yj�"O���򥗦#��Q�DH�[2�]+�"OΨ`A��!%��1BÒ�*x��5"O�!���#J�	�C�
����"OV)FL�0��8CU���V^�:�"O8�Yp-߰� ���r��P�"O�-�T�:���m��b����5"O� �HqQ(�9k0�qZ��	:�i�"O0���MW�t>�JCM�c��MXV"O�T�b��(7>�k1�,	�h���"Oҵ��ӅFO�(
�㕋\�} "OjD�r���h7��եL�"�@u�a"O"i�'(�6ڪ��n[3qў���"OV}sv��;Nn�ڱ��:�0�{ "O�,�iب%\�x �g�?,���"OD��iG�$`kw��W�PH�E"O�9�B�^�&!A�A�n�Ka"O�� �@C�$���o�RO��"O�i����0Ce����hs�h�+2"O2��(R�~�Aᐭ�7ۜ`h�"O�A�� �Q��{b���(��"OT:�ё'���b�k�;y�0��"OP	D�Gˎ�h7J��pLu��"Oz��fI�B�L����Q �}��"O�I���c�� �bIV�:�Y�"O>\[Q��`�~1�*G�V��tڤ"O���҉DN��3�*K`aZ	��"O4ub��ǡH&�E�C�ܿ(�
y�"O.��5/ ,:��S�³T�|�zU"O�ɲ �T�]��K3Q��"O,� ���BG�:UdM��㛝M�!��Q�e�)��2<r����!����,bqgI�V"�9�UA@�)�!�@�z�����."�<�QV�\�fF!�"sr0	WE�e��A���&,!򤜎T�,$k��#LlZM�$D�h!�DTi�ɻҨ-u0t@�c	�o!�d���F%�G�!~�(p-�u�!�:��I㋚�$��ݘ
�!��A6x4,�td��tm����2U�!�DK(\1���1�����	J�!�ė*U 	��ᕗ^Ķ8���e�!�D�&�2- '�C�0f%��i��=�!�$��UL!Pc�{�|��)���PyR(�2hX�Ls���oVZt[b��y�K�-Ҥ8���� ^����� ��yҌ�/KW��Ӂ�#Y1Q�R���yBۭ�jԙ1#���^yyb����y�o�(x�F�TjW0��bsB�y	�=P���&��7b�R�U>�y�BϏ3�>Գ��.�@�����3�y��G�^�����J�z1�ᐅ�y�N0
0ir�Q�t�0�
�����y¥A-G_�e�Ǔ�@jU"����yR���Mn]�蕊����m�y�	�n�nDj��T�xϪt�&����y�D,K n0��_��iㅅ���C�ɳ;6+o]J"����=М��'����,��;Q(pk0���a<�-��'~�y���[= ( R�l�V9�
�'V�=J�a���5c�
QǬ8��'��i���0�����J�n{�'�:��@4I�5�ț1�3
�'�̜ia ʔa�j�3%A>�L83	�'�� �/3����`K?Nꈫ�'�j�b�ǚ�a"� ���=X���
�'X��j�>��P)�$��|h����'� �çh(}�|���ʿ��9�'��X�Gc�"<� �@Ջ,%@��6�\,0��
v{R�{WFMx�t���A�S.Ze������
9Tԅ�S�? ��� P03�V�Y�ʥ~ȢD"O�]Y�>Cf�="ֆ�,��9q"O�U�d�'4Z����W��aI�"O~�fiH�A�����?4V$�aG"O|qiT��~l�Y�D��)@v�&"O�(�F�2*��lY���
GL
��*O�Е��h�\�2!�����
�' t�Ϙ�Bb�R�G���{�'�F5���TG+���Wn�D��EH�'@h�ȝ2�}�PKM�oԎu��'�㍐�j���V���a�L@�'t��S���0�^/X�ੇ�=�z܉A��_�� 9�)̓\8���ȓe�ĳ��ݑl�<J7�&k}� ��H��} Ǭ�?+�.4HS��1$���JO�(ɥE�a���a! �B�)��{�kƎ��@��F(��v� �ȓ:7I�D)?Ρ�lV�3���N���9�+� +�6\ G�
ݜ���7}���O	�AA,�Ud!��@$��H��|�ׯ�*���`�ް�B�É�h-@�={��ȓz�� ��2N��ȓ4�K�7,�i�ȓ'>�X��&�.��P�7�(I�ȓ/�,�:6ףg���#w,ӈD��H��#;�8�V�ɲA�sá�WFE�ȓ$���FB��>~l�ȓ%�RE�wk��t����@&ي4 F�ȓ#\ �#/T�� ��ʚ�=�޸��M��Sv�- #���Eك&�0��ȓ2�b����]�Hf@�k�ޣ:'t-��TT��2���@�"mN�ϪلȓdN��'e�6)D��B`��n�<�ȓV�Py2�@%њ��Z�&X�ȓV���H䀅'��⡦Bv�&��ȓ@&��e�
�E��D�ԅ�i�b̈́ȓ���[��U�vפy+D��a��M��wܱ����	x�����	�lhD-�ȓ6��zRh�i&P�
)���ȓ����ȉ�>�d�'AZ�!��l�ȓq������7�PAx�aF �q�ȓo���qM�4i`�mȥU�VT�ȓs�FH�ŬC�[��҃�|�p��PU�U����%�ԉ�K�(�ȓ{EN��Bo�%����b�ԅ<�@�ȓ?��p��/�aB
09!� �:����z^e���pNl�(G�P�V��ȓq�0 #Տע4�����]�@���$����
�$�3�mQ�6�����7,.�P gC�:� � �f	�Wo���:Z�x;�� "
�@1@��ދJ��I��t��a%�{�8 `�/e���ȓK��1����>�\ccL�S����,�Ry����9j\�����[X�L��x����#��<1ؔ�#B�ftZy��g6��glD�&�����iiL��ȓL��-��I$;�2��ӧ�1H�8<�ȓ8��,�&m]9Y��{7鋖Tr�<�ȓ�|#��=R~�!��̝'��)��&x��&kϛ�n	i���7��ņ�jb(W�q��_`���ȓD�\�����	KO��	�J��XXY�ȓ|A�X�&
(	r�
DK�+TH��g���c��d���"�)NC�)� H�Cdin���ʇ@ƚa"���"OxM�E&Z���ŠL y�]�"O�|�7��.z�`�`�C���"O�4� \�s��Rn���"O�M���źdp*����>/YĒ"O(L@�o%r*TYc��.K��j"O���w)w� �	��ݕvWʬS�"O��	��6z�Ljn,(3Rp��"O��4�_0}yJ�X�M�]�"Op��ԨV�7�6 ��
���K�"Oxx���ʤ��"C�<d��d�v"O�XS� /;r��t�RHan�b�"O��0�zD@����8b�����"Oha�7ʀr��Q��c�5�Ї"O��3p)�	>��V��	v6�2A"O�y豍ƓEk"���HT�kKr<k"O
��玨~Z2&� K,�%�"O:\ZB��	={$��"&�D� "O̫�Gk1P���n�"1l��'"Ov� Í�}2���  y�^��"O
E�I\�p�|�R�"�2p��"O�0�@D���u�P�z|B�"Od�����#���`�\�
���1"O������%ML���-�f�D�0"O�����\�f`C�e
�Ph}3v"O��a�!�5[�$5�%���d�K"O���E�B�\8:�8�ҮO�!��� �zQT�V�mN�ř��%$�!��6i�5`%ɔ*Lڑ�"��M!�dC-!6h`�2�*���nĊP�!�$Y�5�x���VϜ|㴇��^$!���(<"���`�8
�E��G�T!�H*o�j� Ì^�;��<��Ǖ�b!�7O�h��bV��zi�A�p"!�D��]�p!�H����$�s!�d�#=��;EF��U�8�p��K8	!��?%J�ɷ&��tg���虄n�!򤁯7-��!c�X���>�!�D�hC��#���4 �y/Z�(�!�$�	��k���s�t�I�!򄍧.0�Ei�A�cj�� ��^�!�$�2]��C�MV2HR��s�σ1�!�� �aN"��$GW?�퓐CE��!�dI�H��!��ܣqB�I�#�g�!򤅧\��тӮ0W��%¡��+8�!�dMH&�2'�
�Z2U� L�n~!��֋	xt�b�C�ww��(p�$2w!�dC����PWIi�X� �H�,w!�$I�"�z�x�	 R�X-�al!���Ȥl��#����'[H!�䝬=��q�m72�P�0�O��x-!�$��j3���B�� B��j�<��N��k�ŉ�f�:��.���ȓu�������r1��+~�*�ȓ%[.C��(�D�"� *-�`���th8�J�˘�f:�*��@?9C���A��=+�F�9ڎ���7T�B5��@�R�����Vd$�+pV����dUf0���9�0L����N�ܥ��-�d�t�ӇWv��ۤ@X��2-�� �@@�gI�L�J�I*�LV��ȓ ~J��R7U^�9䞼����a�L1�`�-���r�ݠe�\��
��j �øG���j�"^��Ȇ�S�? �=���� w��\��:��(�"Ol� ��;gj��#Oэ�&�P�"O�"UA���r�C��|���"OPD���� 6)2���U�4�A2�"OD��@/]"<�"��6�ˏ1 �ʴ"OH�yA�L�$��f#��B2 !�"Ol96(}�2���#M�� 
�"OZqɠeF�9��[�,ܪ#�jK�"O��d����h7&^9!U�
�"O��"���ifB������K`�rS"O2�$K^'1����}B^��"O���G&@=����±)b !�"Oz�
r��x<��q��f	l`��"O�bk@�^�na����,*��9�#"O��ؑ��d)�B����t��f"Of��5�Y��`���#*yXa���?D�h�@A�$*�h�3i�.-� K*D�\���5�p'ҝ)�6��'�&D��R��EN=���c�ì�(��!D� �Ѕ�g���BGhB5����!�>D��:gA�OLT�DdV�U���
P�;D� ��	�&gP�C�O<B�\M���9D��Z�/�ѸT;� �<�~�h@�8D�:��ߣP�^�q"��*v�p��G<D� ��IC�s��$("����<���$D��+�AE� t��(ǥh��z�f8D��s���S���s�:Fx�p�#<D����L�S5AH�o��&����9D�<2'$�D��D�����b%D��i2�H^%���G� �ɤ���7D�H3R����V ��L� px]�0�4D�ء�ر�6m�#I�>f9�w�0D�P��G k 0�	F������;D�����y]�ah�1V���$.D���Ȃ�Nd:|��aA>�d[!� D���C�� k�@q�dA�ckhQ$T��r@�Ymmh�9�-Q��8�a�"O�]��m�C�*�@&�E<�0���"O�<�o�&L�B�KS%˹8c,��'�(]"�b�-V��a#�P'iL �����!����-�4>htER�H !�!�D�3/�DC��|G0A26#�1�!��V�^&Д[�͟mMLu �i�){!�G�����z$vx�&�H�!�1 ɡbә�4��!�DK0~9N��A�ث6-��A����!�D��
,+wl�,SPa����9�!���k�"urF�	�L	�d��6*!��XlN�SQ!c�h(i��W!��6庵�d!F�p�^�z��Y,d�!�dS
��[rW<���H�H�+�!�䚥N�z�'$?G|$�A�Q�!�D�?C��C�,Ɲ!�����a��!�d�-#:����-(ʮd��C�:+�!��$An�ȃ [1{�����Q/Za!��W�/B00n m����!nİv�!����=D*�"��7(�����!���z��9yu���������5�!�$FzN�M2q�I.W4%y�ϑ�
L!�ė-'�.)����AD!��	�'�����ԬM"�p�"a��R �3�'�����"v��e�"k�U5����'pԁG:=���AG�ZM$�ϓ<��ag�V��D&y���$	�e'��Q
�qs!�d�?0�����=s�ء�j_�1��'x�\���?	`��� ¤��.�b��tp�f�{�2�Yr"Oڸ�j�((4�
��t��SPbͺ)�B�,�(�9�`$�3��ۗ{2QU�?MH��A��T�E�!���y��2�PR�x�yeÉ�A|Z�:˚� �5�XX��(")�4�HX��G!F��ط�(�l�ttᥓ�A]�)��jb7Ÿ;��@�0�2. }x�!p�<9Dh4`h`����`�sy�ᙇwPh�#'���i\
���(���sM�x��9�!��8yg�`X�kA801�EC��(u� ���
���3#޵Wq
�:�Y>�<�Q���ű@��+��Lkc�UHX����F�0F�ɓ	�6�]%
֣�x�Z�I[���0[@y9E�Vc8�:F��� �n{��!��Q�$�q`P�3|4��Q`D*it�=�Q ����ƅ�m�}��K�+�aҴ�y�X��z5:Ƨ�
���!3���I�"`{T�	1	Q=Lxu r�l��ygA�h�(y��צ�~Ma�.�yb�Fo���*�e�}����BX+�|���kX*AP��W��2$��Z��o���Fy�D_P��\k K�pǾM9ҀS���=GL�'.�7$��U�:A����v2Z��Р�bt���]ݮMr ��a8�	�g��ed���tn�uK�����;�I�Rq�U{�F�����3	�j��0;5G�?�°"�m�:I��ƑP�qҮ<D�4J ��p���I�MK!>�ٳAi\����bg�C֪(��iѾ��-j ������@ߙHY䵰"�=4$Q�4�w�<!�.Ҫ�q�#j׉(���g�֮$�6����P>�h�����-{�r�"�Nҫ|��<YքR-xh y&��z�Z�*���i��L�QC�������M�P|+��c@��'�Q�]�p���4U�"\s���:�p>��	7�8�RM��-:2�ã�b�ũaϐ�H��6	U�o�"X�a��I�qQV0I���6y�W���!�$�1\���C�e�,�p�E�H��<�%�^�SU|��2�M�qU�U��0��O�*��;�Z�����8����ɞ:
8D�ȓ|���Y��Cf�\�RaB:q�,1�7)I��* �)�.0�K��ӡ|���aP�"ʓj� qK��ͥYIH�yb��9b+�!���j�|��.��c���JTMA0m~�����<C�(h��
f� �vN�-ւ!��"\X���6nA:�I����	�=�h��K�<�r�F�v�m3� N���謟FAY�R$���@g�6#���D"Opzt�})�!�0+O8�a��v�|  �'��)��D�0@�P�J'§�V��MXa�c�#d�n�(p���6L^C��-�h=�#$��$�nM��4��l�R��=E�s�5-�֘`n�ٺ���N�.:V����#'	P��ӟ��{� ��wj2�9�M�,9��D.� !=�A��@��.A��c��,A�	
�� l ���(��Aѩǒ8Kh	Ex2�-#�hɑ"����Xgh�����ah��oOЄ�B"OH��&j�>���Q��V�{OF�T��)m�2��͍���S��?tR�5�Y[G�\�VM���Kv�<�R��98�N� �EXr��f�p�<9�*ÈJ��X��A��\1AM�q�<3�ސ[�����QQ�t�E�n�<��k=\��)�i�?�`��RC�o�<IM]���yqh���e�A%�d�<��+7~��W&�*8���Dz�<y�	;m��*%a��e�E��`�v�<i����j��+V�!xvB�P��]l�<��Y$n�: a2M�"X��U�� �D�<1ǌ�'ǘ��T	�=��9�	_A�<A�L��:�F�R��W��ܼ�F�B�<S�ױt!��0r ��4�L��M�{�<�Ģ��d�!�Αei>�C7/JL�<�CG�*F1��޽r�4"� O�<q���6eFua����%˕@�l�<��\5?���WI���T[���T�<9�+��d�0�`ې'��H����<9@�ǈg�(�b�ě�88E  ��m�<ѵ$��t�)�:F��DX#��j�<	3���Nu���7�B0MZ ��De�<	�f��$���� �,.�n��i�D�<� �LsE��L����_$~E�T�"O�(Bp�ߡ}��;uF�"x>��HT"O�,)����r�`[�f;7��@��"OS�%�7임 �ޯ*����"O�ڲ�!H�<٧ٕ(�� !�"O.�f�A`�
A��#�R��Pq"Ol�b��9:�c����SV��"OB���N�3�hX�!\�.F����"O�Yє�P�_r�Y:�[�i� �"O�EZeH�3~� U²�4@G��92"O�@��·W���B��A����"Op�ۢ͑(`�,U��ѓ\���"O4|�r��$?,�1׫�3d����"Od�I2j��c�RA�F�D���U�G"OT$��
k皔 @�PZ�0Y��"OLU��ɉ1�$�YBW.(`ڒ"O2�[G�܁`�H�(�s���e"Onњ���b�CF�ߠ��D�U"O�U�����ؚE�<1����"O�$3�ț����yb�5�mk@"O�P�ԯ�'���!�G��d4�@� "O2,���8�}k�� �"��"O�Rab�,C"���1�
��F"OX��Ī$:>D��d�=gPI��"O|l�w���Lu�����ˉqH��;�"O���M�:5�Z�{� Y8O�ܰR"O������>Yu����τ�s4d��"O��yc�A�[(1*M��f?��T"OԠ��9K����퐮z� "O�<��"]3\�j�P5LK.�IY�"ORLr�Z��Y��k�#1^`���"Oh���"3hȹ�)!p>zź "O,Mkp��.%�V��F9Ctp��"OJ�R� �v�����G�ok��3"Oƅ�.7DQ���Z=�0xg"O ����?10�V�J�L"�["O�t ���[�$���&חV���"O�TYюW2*h6YJL[��"O~���Ht����#*�=	�:��F��'w٪�ڍ�	�Kd�)c	;D��1�HٲJ!�d�=j�����˵ l*p��ԁ24@ѻ��I?��gl�|�'�$!Ă�V�`˅EA]3���'@tB�eV�X_��4�I:W���b2j�E\n5��刡LA����	�`���!�9yYDT�%�խZ���d�*r񺜀D� *Y��ۖ L�.�![��P�4���0�l��*���!��ېI$
���F��f�'�$�G��	<"ђG��3t4�F��)Pu��h�+��nO<�Ò��1�yBh�X�vq�F*��t��1�&�U�x��8�厗�n�t�CG���i6P����L>��n�Mc��i�%�v5D"�(<i��n�|P��B�p�9g���Sa���&��pҘ�`T·�q%���G1�������!,�!��Φ/�axR�ߦ<� �(�mX�z~$])��a� �`�T��h���� �̵!�Orh6Ι	\͜-JT眄wU¬�Ɲ�<C�N8澨9��H��!���s���xAAaKG�]0��IH�~x`݆ȓu�HCu@Ŋ-�b�&�Qq�A:7K�7R@�ಯ֟[k��(�G�f�'��.Gf���EW$B\F5y���KV��.Dn���*݌?�n1�`�S�6���X�����C� =(5QC	��<���(D�`��ƥC�u`tp�Bs�$�F�6*��kC#��w*��ʳ'��w�u�%�]�
�ڡ��-��\�Ɠi�0�#f�\��%���R4cS���'���cDMZ�m;D!�m^]dΜ ���L�`��� ������	4�!�$�T���x��`�
t��(q�dG�Q��!��0LƠXLC1�ĒO�`��iP�l(��u�$=�0
O4]�$"��v��9�J'�%��^�8
�c�N���0=� �PB0��=`��ls ��6��@���'���
�A9��T�sF-����4�Aa!�;{V\[�H�I�<��g��&�h�Rp�7
-$��M�ɃoR\v%[�}����$^m�Ojd�d攈c���6L:f�����'�(9�Ĩ	��`��Mv�6*ҒEJ�b������ � ���ē� ��슰(�@�"^sBh�Ɠ�*y��	��.u���ՐEi�y���R�yԒ0
щ��
�Z��䒠pL��/�I%z3v�zr�z�#�	�Y����<�g+R�X��<AR� ~HiR!��Z�<� 
:>��T ���,��g@J��@�c!�v��d�!(�B\8��^�y��.�>�I�)Cy�~5`��ѻ_y���ȓw�@��"{���×0*k\ ��_��c�"�$h�"��%l��<�ȓR5B�+�)n�+-"n�`�Q�"O��rA�I&��óLs˜u:&"O�ѡ��՗r�`Q豮[�w����"O����D�?C�Z�;6�]<��m�T"O(��q�Uk8�R%�
2����"O�)�'f��lF��&*B�*�,1�d"O2p� �(�X��P���w�1�P"O��%�47�`1C�,B
M
2,��"O�tt�2T����A��q�	
v"O �Y&k�<������&h�Q"O�)3a�)Q6`	aC/�zeb=��"O4%����302�{�,�#zEΉ�q"OdS�l�s$r)c녂G���kG"O�p�����*zpu�j�8st��[ "O�}Y7Q��R��d�Ot֥�W"O�̓���o0~e�`�!P�D���"Or�C�ʁ)M��l�� ��p�Cp"O�q1�
�z᎜c�H� dy�xr"O��8hB�о����/fb��"O�a��SC�F�pǫۏXfN<��"Oΰ��a�;%���bQD���� ��"O����C�h�:T+vĞ�[�z%�V"O��r�N�0��X�	Q�a��8�F"O,��r`�#k����ȗ~���f"O�u�VC�;pF���7a^}��"O 9���t�Q��V	)g�ċ�"O2|�2%�Z�8k�)��at����"O�EPT�D�MZ�И�'6P�{�"O*�s#�V�O�u��ѯd����"O�,Z�M�:\�,p�Z8iT^Lq "Oԉ�c�����r�.��N_Z4��"OvuZq� wƴ�'��%ʐF"O��!ਛ/n6\X��ſP �q�"O�]�Q �4	N�� �M�[���4"O|�
GEU�lf�8�ϳy |T"O���I�W���J�&ů\QFy
A"Oh���zҥ�g�[=*�b�"OP)CD�B�iu�\�a/y*�$��"O�cg���>���J�oT
P��"O���P�Φ0��уM�7
�4��"O JN҉�6�Q��D��.�"O^�8�V�Z( @8t��ag���g"Of�7`�*�`�)���W���4*O6����ܱv���
�V�s��1�'e���C�	���cϝ	�f�S�'E��1A`ʐy;Z��1fye����'�Lِ�cwJ��PPѱ$���z�'�81j��p��m G�A;���'��cƊ	#JR�0:'@";�$�H�'|~�DI*%R2��fG?�h4I	��� R�Jt*R�|.DT0&�,)c!y7"O�)�k��v=5��C�?ri�t��'<=��׿��	%I�.IC1�O	6xձ��� C�I=7 ��R_"�8M42[�O@�ib��jg�t��Ef*�0�g��p�y�o��g?�B䉺�Tͩ�)�?H<|9� iU�(}��Cq.U\~�a�+W�T�}&��W(��'���"�1g�h`��+����Ø+}N�H4�>H�Z��a&y�h����GE���K��Eʂ]$t�վ��b�&�w�@Ah"�Ō��]�J�q
g��V���o�J�E���W�<Av��8sD�!�w��*��d�Jgy����dL���"�>,�����	�;|:%q�Ƃ+H4�`�C�f�!�����[d���o=�с��D�I�t=apAڸD��p����{�Z��]>�<aa-��u��Y��)V�8;�Xh�KsX�H��D�5d(�y���G@�F!�g̍.k��s#,-X�`xxU�|��`��	� F���+�e���p�.֊YJ�<١%T�&J�ۥ�c���(T�����O��	�@�&�����6VX���'���w��9\���-�8ĩ(��x�ց[���1%vd�q�I��E��w�rd[G�hW����Z[(�B�'��lĄP��* ��/��u�h�BI��A �#I��R˟4���o�'�Fi��#Z@���j\�t_TX��n��Y
W%D�n�PE�+�!l����@a��q��i��d��%j��^�I���P����&�]�Ipu�fb�f���D�l3�v�c���8^�:܂��51�l�SSY�@�C�^�(�V�%\}�PC�I$	��`��b�K�耺t�F !<U�`om�"A�F&S{^a¢���.Y���4�sޅb0�U�Z�b����u�j�#'=D��hB�+�G�4���$LV�a[^�8ⴍ�t#�/�J�z�cF&G���0��J8 �Kt�X%�@����5���d�9,Wfܢ���6 H6��t���c��y��̒�{�Թ�L7nH��Cv��5Y�$!��I"c�(��F�Q��q�%W�DB㞰����'�-���j?L�j�L�)���0�O*��R�Y�8Ć��k�?T��yC�'�8�"4��mA�XId�<P�zlƩҪDL ��$�B��kE���a�0��~��x���T��sƞ��vg��F�D�b �,D���-̸v�]����(0��A%i�t���;'�i��\Ӳ��Q�����9r�Q���'�~<�
f�XC��b�7\O�	A�%r�����D�thVH� g�iؤ�8��^)d�,�AFĦy��-�K8���q�_�jQr!���U�Sjmke�#�	(����`�f��}�����dȨ�k�t�]�E����ȋ���@a�
�yҬǙZ��BF��Fw.`['*5p�t���.��`͸5P'��v�:M;���k���-�!��
$qiJ��nD�M�!��G�E-D��3�%Ji�A#A+E�3�v�S���<�@L����5�Z����D|�EA�JZ�#%AC�Q���rPEX���=	U͟/S�����AKx�Y�͔.J�x�t���WZ���	�N��	a@v@;��Qfѣ�I�+id�#<i�;.ƈ��F�Sy�O��Q��{�>4��f�!FX�];�'��!q҄٩dH"���Y'7�F��qO]&O��Z�Rz�)�矼
��%�����_�q��\��$D��+��<,��9GK�h�
ݛQ�"D�P!���s�v��@�eF�89�� D����&Ǽ_v@��n"tMR)� ?D�\#�FݏB,�u�p�q$}�cd?D���E��:�\-�fC�S���ڷI1D�xB�ٰJ�=�[��40��L�!�$�PMz�Q�Lϔg�MjA����!�dJ�Oc�)(e�ǝ	�����x�!�dӪ}G
8�D�=*Y>ݐ���*De!򄏛[ǆ�p����x@���&�#?a!�$2�	����7DT��(�84U!򄜫YP�@! 6�������:G!�ĝ3��Q�m��<����-�I!�$<vpƱ�5J�7)R}�흽P�!�YGB�뵁9?�@�\%�!�H�Bx�A��� f���oB��!�^X�u
�@�N�>՛�?V�!�� H�8#�Ϩ.�������H��"O<�YS���@6`�2��<���"OHU�A��_`��,*	�}S!"O��#L*RL����!��n���[u"O�YA.��U���ˁ,전�"Ovyc��ppSS�I49��"O�x�/�t:�h��%/�Y��"O�AbU��eD��
Ts��,e"O�)�V��/)�(b�j�3��J'"O�aCP�2�2H1		��!S"O��0�ǻ�P(r�h3�a�R"O�3 (D�/,
9�ѧ�M��@JB"Ore���L�D0 -8�������"O0DR�����|�*�G��w����"O�����$��xYW&A�T����"O&)�e��x���%�����"O���ូ�Q�O��g�d�q"O�<�P.�DX��J!a����"O4��B��}*8y-ȈD�����"O��FYp���B�M�)
@}Y�"O�i3��$+,PP�6&�p�\}��"O�u�b�ށBl��)��J�
��!�"Oz(c�_�}P�Z�gU�_StJ�"OĘ8@��T$��D��@���*W"O>�s�cI�1R��PD�rQ�X�"O��P*8&�,��Gʞ		@�qA4"O����ZTX��2G*���"O�T8ң��/�QF���]�D"O�,)��		~Z�$SV�F��rA��"Oĉ�J��^��c��X�A�p�&"OR��R�!Z���Ыk� �I�"O��"�ŽT�^�:dM�/r�6(ʒ"O�	bu�R��J�.N_UR�h5"O���Vc#����l��s312"O\m#�L�6m|<(ؔs#f r��>D���,�w�	j�&Gu� ��"�:D�X �/���Ƭ8��?
y��ɶ�?D�8� ��#~[1�2>K���(D�䛃�[�^(��y�R�F�����) D�9d*��/,���BM/~HD��s�;D� �a�Z�H��5���)L�f�2�9D�xa`��b��[@\5B|<i��:D��ۖ�nz�8	d�� i.H؋b?D��I�eĜi� [��W!FdLB�N/D��b�ؽL�V��'l�lE*D����.F��Za!�d��F�z��&D�hI� I�6�J�k�*L�
�����$D�x�����T���3rf̂,D��3EߏN����K�B���� D�$�A��2-��zW���8��<D�xs1 鶴�5&ݝD�
����6D�4ĂT�-�-�]��0��8B�	�z��L�k:@�J e۶)FB�I���p�W�eB� x�W�$:B�s��$q&���8�p@��9SB�	�H�vE�C �Q`�����Q&C�I�� I�bذ�d�b`f��C�	1ne�zs�é�����`�=�B�I�q�D�1l�96eHAk��A�O܀C䉩��L3S͜L�N5�C��m�~C��f��LD��~���&�6QMjC�zZT
�3M%���o��bgvC䉟s��3�-^3k�U�@�	/~W�C�/?L�H�c:&�X�с�8�<C�)� ���T´C�uC�m̊��l�C"Op��3�;v�;Cl�{��љ�"O��Bu�ҏ_o� �,�p���S�"O�]��MތH/tS�!n�x"O�����,
�Y;7l�a/�ę1"O��hW��(F��Cu���[!"O\���C.v�I�'*<���"O��#�P����"�$6.�2�"OI'$D�z�x�x5!D�h����"O8k�@<DZ�$����<k�"Oz�J��;|C��r��{G�!"O~)	��F9k��|���SJՋ�"O<)��G���6a����aZJ	Y�"O��B2�;1�A�a��"���
�"O��{`@�)�\��/iwԜ��"OVؚ�+�b# %P� ���2"O :D�4K�tض���9kBi��"O��jo�������4m\2�ڇ"O,ܰ`Ʌ��89�����9ؔ�"O!���?^�ҁr�(�Z��<3"O`@�C��6}�l��B"5���@"OF���2 ���K"�A�!���j�"O��ѱ*�+g(8��oB��� �P"O�}��͈���bcy�"O�0ʷ�3�:�b,	#(_\�HA"O@-y!O	a�)4="D�[�"O4X���}�RHt��'�]ʢ"O������Lɘ��ۋ�I��"O��Y�A�|�*�8D�� #��Mb�"O�\:U��+��m��'�(�� 4"O�]����`�ҥt�ɉ�X��4"O^�Kd`�,��m!0e�F�V���"O��"񥆉|��,P��FPt�xA"O��' �:�Zm��E%29���"O��A!IQ�����4]-r90"O��V��'�\����w0�{"OVɋb�-���c*�j�$*�"Oh9�Ř>*�����
�z�����"O�ZÐS����rE~�\��"OL�y��Q
��ue ]�`�D"O��4͵EO��aD
 0��k�"O&�$R1=t.��֗S5��� "O$Y�a��6xA���1<�
�"O�E9���$(�9�nO$_>.<h�"O��8g���M����a*ļGJ���"O�E���Lrb�8��U;D� Y��"O�x6�ҜX��a㗢��� �2O2���ٵy&$��1���$�1 ��ɫ*ϒ����,@�X�$�V�f0B�I�.�BMjs�_&?�����('3ZB�o�n�x��=*}�����L�h�C�	��� o\��Z-)��Ȗ����(?q��U�~}�5��M��`�<1ԌˊX��-q��UQ�H�1U�
w�<�a�¢��@` "�k���S&)�l�<�*j.g�=�.Ԫ��_e�<ɶ疼KpxH2'UM�ܐ��J\�<�rُNHcƝ=S$pZ�bRX�<�g,֢?%v���G WE�	��nJj�<���7h�� ��DP��	d��b�<rDث��E�2�r�,^j���E{�G(�����"	�2��x����u��<q�����'v���yU�C�2LP<����&WQ��9�V�4I��ا(��$A�أx�}z��Z��76O�9�'
1��?y�>0nԐK: ���E��E�f^��D	�����?� ���Ԉ;?.�Ivcէm���Z���H�'
v��i�'`��p�A�&��Ua�.��Oڹ��i>��\�`y��S�/ت�����!pz��%�P{7��o�S�.PX�g�ݺ>��S���'�%�'���a���ӟcԘ����! �x|S`�ٿZ�>����(O?1�WDϺd�	�	��ł�"ac�<��?3mZ��kMe�2]
4*^�<Ys�  ���'eV
K��,jEq�<�%[�M̆���d��#u�� ��v�<Q�O q���A(��(�6��G�u�<��d��*��=�t�zA�^p�<U�K�N�0��q�5JӁ�v�<���%(�p�ڇ�w�p�³#�r�<A�čA�Mh/	s$��+��s�<�0�\�P�2��@�߂��!BIW�<�� Й-�0�c��,+5�CQ�<�AI b��e�,j�x��&h�<�r�S��Hf
�*�T�#ĬNb�<�p�O��t���n�"t�ƽ����C�<!4�TPj�!]:�����=T��J�M׊GP�[��(1`��,D�$��h�4���CF�0_?��;�+D����n�?U��P�a��t)�	��(D�v�i�ê���j,�+^Rܘ��'c�0�����8�ʹ匊+j��x��'�\	/Cd'���Tˉ8_(rt��'[D��@�1~t��3����2��'��Ĳ7�ù^�003��%Py�i��'z`a�� ����oV�xXҁ"O�Q��R��m2���e{�"O~���
Ւg|��f�OV�8m��"O��{�jP%H���S�|x�0`b"O��"��t[r:�o#O�\"OT��c�޼G�D����G��};"O<� "Q�Ԁb�G�K��9��"OF,KՇU>�\tq��2\{�"O�Dį��@�y�i�6)�NܢT"O�3�Z�i�D�V��D�aW"Oz��S�L� �q�����p<�"O*Ⱥg�?}�x�Zu%VT�\y�"Ox�Z �I3"\���� ,:̪w"O�$U*.�:�c�@�#m���@Ot�<���4\ܦ�S��R �e �iF�<�0�<QLxPc��X���t�C�<i���q4�rD�O�S$BY��|�<���W|�qhEF�	(�\��NJp�<��-�8vA\�����f3�4��YV�<IuaN��{&b�*�n!s��\h�<���:H
fLЙ�4���Ίm�<��@'NO�E�D
H<�!�:�	���S?�b��v�C�!�d�;�Ԑ˄HG�a�Tat(��=�!�d�)U:,hF���p����>�!���f�p}�$+̀{�d�<D�!��;�p��C�� n��i�cܓn!�1y�J�" ��J�����4x!���+�ΐˑiBS����T�'
!�B�=^�yжK��+�>i	��I�X!���(}���#T�2]*6�1a͌!�σ.2 ��ߒy���cj<'!���x5f�s�)^�+׊ZD�C�{�!�$�|O
͡P#�M�E���	>�!���
�3qO��e���1%�ՐF�!�� �,��l�0���!"�M�!�� �4�se˥H�N�s�)��aQ*��"O�ɘg�ωS��E�O�{1Δ�@"O<4BfIE!g��0���DЀ#�"ObT8��Mӄ�x��>�@��"O~��@��Jy����(��+�"O�ܱP�GC�0��0[ɪ1�"O.��"i�&E��ð�>�.�k�"O@з��&/6��j��LĲ�"OX�C�jB
8��i�>��9;@"O�ҥ�%HcV�۰g��i�DQ "O��`Q��6Yd��(��[�B�Q�"O�lySǅ\��j����\���p7"O&��`�M:����83��ɉr"O¬�0�)[�X��W �F"F1��"O̙��A�"_ܲ��ɪ��/E�yrN)
Ll�����	�~�� ��yG�L<b��d�BVI�`������y�
ڀe�$Qum+c�<ēE%Ԍ�y�X"�YG�C-^Ȇ�B%O*�y«��l���b%l�;f���8 +@�ybM�2<�LAbq�-
^�,��
�y�i�d���r�9|�´3G`�?�yr�7|���8�h�KB�K:�4�ȓ_nq�1�ѷ	N$萦�+O���ȓh0�"�����['Z�9[�̈́�~s��b��!�r,a$EB�2�:Ʉ�,,x2V
����i����%�0نȓ �%8�mX*���V�R�5����!!g	7~u�����ޒ
��-��{��T�&̂��ʔ�We�)-�l���$�.y�p�֨Czm�f)�r�L��t�RI !��+;�4�F��ni�݆�7V�m�"��Q�F��e�%���|g�� 瞹+�A�SI��j �i�ȓ?�*	A%r�lx�Ğ�_v�����s�K�����E���i�`���-��1 !��R��72)h͇ȓP�Ј��ŕpf�u�i�	hE���(yy�B��WQ�|�'���8�ȓj�"�Y��XZ�P�(�*n깄�~�*����	�y���TBD<XSd�ȓ*q^��m��h!<0�&��k���ȓ���1���{��)��ί>M(X�ȓf��" Z�h�b�[�wX���G����׋E�7���$Ҽ~�怇ȓx\t�h`-��7P$�s6"\"h��@�.��b��	=�|�U&�5��}�ȓ7b� �I��T}��	WKP�r�J�����QCːx8�6�3A��9��b�� ϞY�at���捅ȓyŎX�s�R�q�X�x��A�5����^�bd�d�@ ��bBi��<�F���elv��S,�gꌨ*��� �Ą�a7�$
���T�,l�րB�4���qr|˂̀[w��!����y�ȓ	>ژ:�I�es���.�(Y���ȓ_nD���M�8�%�P�ը�2�����cGGD�J�, �Rl�ka*M�ȓNX�z��߁	_$��jӔR�\���0���g�TE�4��c%��sC��ȓ_=4�RDwfe��KW+E���ȓVs�T[��?/����R/T��0��G�r�J�
aĐe��@�7rp��;��Y!	�01�A���S4de��S�? ���O�>+�TMc��	3LY"O~��#cP�Qy�tP�h�
N4Y2�"OJY���N� ��8�i@�dhm�"O�e#�AYN	��&ޮh슑�#"O0�a�k4m�~�c(ҳ
s�}��"O,2��D1,a3L�:;�Q� "O�u�L�� D��e�"Qƭ��"Oޭ[��/�>�D��RW
̊A"OX| f��&q�8r�M|<\�P�"Ol%�r�-%�uʢ�!4-"�z"O��pʍ1m��M�D�A � C"Oބ�IJ�,a��Cm޲|z��"O>�+�(Ē_d���'LJFRF49g"O�8�FJ�{A���*�<1�=�u*O<e�#���KO�M���f���
�'=�Q��#�o���D�r�ؕK�'*|H���M�5vјU!�>�&P��'��%� �!z$t�����G��k�'��G��%�����a��P_�eq�'�����	Ю6u�� ���I�H�0�'���Bl�=���1� ҕx^��z�'njQ�#�!=�TE�F(H�;�xd�	�'�0�ڲ R�,\�+#��?3���A�'��[�l�;ޔt钣%1�XZ�'}d=q�OT(+l.������(Bd���'H60���̅
�;�!V7%:&���'�jh�C���&<0Hpd��(��k�'&F�;�Ζ�5������$���#�'8
0��j�c�m��5p����'�,	#���d
d}8��ye�a��'�ӄA �"G>���mϚ{��IB�' �����C��V8��d	@�G[@�<�&�t����7P��A��x�<�b������(�i��8��ae/F~�<a�fG�`Ɇʧ��
7�N��ZA�<ԅ:S�6}��A�npj���g�s�<A�o1p�u�0
8�l$au�Pl�<��N1Rm켁`!�%V�p��	B�<Yq�D�06U�a)N�q�v�#*ST�<�E
�
A�]hP�L+"pP���P�<��ŋW���	��I�x���+�g�q�<7b�'Z���he H��b��Øm�<9ԅ��K�\T�F�ucd�`��!�yI.~�8�I�G_
���
��y"�,7Cz���^?B� tH�hܒ�y��7C�\����F�"ȑ�V��y�%SA.���J2Bi� � �D��y��b�)��CR�:����ǆ2�y��D+v�^���AL;�ptYrb��y���	�@ب��S�d��ac�B�y"	��j�Bd�T�^�`J�J񫑈�yRf�.j�1F�G�j2 ��֪�y"Ɏ�=�e���K%��M�u���y�fD=���S�H*O˒���I��y��$����hKS��� �0�y���[����$Ets�ّ����yR/�=��Ҥ�O.W2�4�_��yRf�D�n}��K�op �	��y�j�)5�n��FJa8��K�AR��y�Ȁ/I<�0eŔ�{�`��P�y����f1� ��M�k�hI��ˋ�y�oA'!>������dq��T�
��yR��zGJ�B��n��1����yb�?%�R �7.������y
� ���ЂE�'�X�+�.;��2"O0z'�T�[��U�K���6�"�"O�dxV��	�^A��*ɡe��I�"O�A�VgV�m��u��	�$DB$� "O�=��E�#���
--�\ �T"O���biQ4j��-�t� V�z�1�"Oaa�bU*�RP;6�� ��٦"O��X��ǆe=@
�k�=� P��"O�I��6l� A�0�
, �JQ�"O
a�� �Z����g�'g� AI�"OĀ�f:M�T-3�
�[�\�"O�����Ǫ?��^�D���4"O��x�
   ��     �  d  �  �+  �6  aB  wM  vW  �_  l  lv  �|  �  m�  ��  �  3�  v�  ��  ��  E�  ��  ��  '�  k�  ��  ��  ��  ��  ��  ��  { � �  �/ j9 @ [F �L �M  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�	�� R��g� �t��B��1�s�Ee� "<E��'�����?l�i�|����y2�6�Şw}��̞�� `�d�ǁ���a����dE�D��p�i^�;>��S��%+�|�L3}2jN,m��+�lRu��iT�y���>�����Q�g�عQ� ��Mˌ��%��|ph�9IV��1�!�;qu��UA؞X$�>�XR��V�ԎPԜa�g��:]&���d(8a�МA��řcYx�h�G��%ڧ\�ƠB�!3]��`��G�44��^�Ȅ�-J�S�d�Ӱ%�'
<�'Bў��$��Fa�,ʕ0�i�9j.!�$�!i�;��@�f�I�Iſ+� �牰D�-�Dk�;�Q���c�C�	;<�4Qd �
����'�4��'��Bm_�K;�HاA�H5���|�����Hȸ-&�tbr�Žp#��v�/�yb(Ͱ6��9�L��o�(��^��~�!�S�Oaƙ�gh�[8|`c��e��e�'% �;?ʡ��� J���
�'��s0i�3y�Bd˖��Vy~9�	�'�F��A�^_8@�D_�M}F��'����7�[�Y��:C��JF���'�*ex��N�d�B��9;� b�''��SѪԮ4	�#"K��7cL�8�'����d �el�0J�g#����'�HS��Q��*�р�	����'a�|@0l�9�0�p�A|�`<��'/x2���93�]���:%���`�'W��P��҈4�����)뎨2�'R2K����y(J�0�D�Z"m��'�~���j�$)ԡIg�0����G��O����^�E�� �9rdx05$?��{rɚ��I�m#��Q��Lm��$*Ǹu��ʉyr�'q�x��H��t��ѯ���r�H0ND$��=�3U����"��M�霂���.�69���ȓAR�L��/�B��ǭ��-����=���?Q��Ӟ6 ʝ)��^�%x"T�&��~�<Y���7?=f` ���4~D|9qM{�<����J�Fa@o�`Ѡ�sS�Q�<�[y|�d[� r:���`n�EB�`�'F�|�ڮe��)҅��F��b�O���	^���O(���b�>�bI����O��p�	�'eF�Js��#y��L�Ǆ�U�
yK�}�x�鉷4��9{�ɐkL����N4Z�rB�IlZ6�+l�	<�ؽ���Pdֵ����'] �cV�`����jG�%��9�'jX-���_�"�ba던�Da	�'�bY��R&��l�� ���$��˓�(O��5,��N�R$�7/T�j�~�J#"O�BS�]9af�K��G�Y;b�s���=lO�A��ydVEk��ה:0��"Oȑd<$�X���$Υ|����"O���t.R9ǎM�1���S
nj`"O�:AJ���,������eh�ha�"O\�!��שn=Ҍ��$�	'�<Y
�"O��#@E�U��C��W�9���"O�؀�J��}:5��k
:�P��"O�D�G@فE5ZA�Cj`D����7O���df��	Y0i؀}�~��)I�5,�,���'���ɉi����AE\���z�&I����5�I�|9������?& �S &�T|�B�	���0p#� ��� �<}��B�I�Jz��5B�% dY��T�A�6�F������ ��A��ƛRTV�BpH�>���6"OL�ke�I�Z t�A��V)(��2dU�p���h��Q#w��
T�� s!�F�H�ZC�I,A:� Iv�CQ��2�iħX+`B�8P��(��_�!�l�s�H�3
R>B�I�T=dX�!��N�ZAz���._B�	,$��rVk[	l��-q-�)
B�I�e|Lru���Z%��� $��>r�C�	0����ThW]jP��-B�6Z��#��c%O�>�ȉ0�F.`�����4�O��$�QԅƪuJ�AK����>���0ƈ3D���� 	F��AƂ�5�a �M2扃5���?�|b���b�c��$��iIGhd�<�0�� T�4+	I����a�`�'O�yB	Q�$�� ��>;L@�cc/_1�y��%&�&aYF.đ-�E �Ј�y�C���v�Pg:��P�7J<�y�n 'Ǻӑ%�0�؍qbC��y�ώ?~�Pt,(t������	�?����v\8���,�H�Pu��!i|���ȓ@��-Ӥ@+n�P�Sd݃B�v,	��O�����!3��q9�(��D���fcҖ^����)"?��,�;�2%��۷�����(�f�<���H��z�eZ�j�
1I�<��l����v����¡К3^lm��	�!n��M{�O��e�k�!�"��"bN؜�"O$Iǣ�W�$�����w���S��D�O��s�{����P=j��1���{�|x{V�D˟̄U24�K4�ҔT�X��CDP�(��:g(I�&�ݱ*�������>�rԇ�,�*I�K�J��f�3��!�ȓ%�M�adT/J�������n4�ȓ�Jt�0o�zB]��j�b���^=�P������[Ôpc���ȓSܐ�bɇ,�����ODN�ȓ&��MJ�� m=j�%)F@�م� �]Y�Fѫp'T�C��J�[@�ȓ?�,�B&@�����1FTl��b3�Y��N��z�	d�.n�B�ȓ9����[��䪧(Ų!xPl�ȓI�@��Q�(]�r�I�Z<��O6�dұk������@�]�(��׈��H $��<1ѧԗk����n�hU�ݢh"69YŨ�<�\�ȓ[�p�Q��L�r��a��_p&ȇȓq_Mb�o˗%�@$�+�# �����<_p�+3
�h�F@�3$����@ua���7���9�'A.S�\�ȓ:����<%�.��P)��(����|��6�Ѯ#���ޠg��=�ȓ-�E�� '��ߓ4�� �ȓ"cr�@�0!{�	�fΈ�
@�T�ȓu+�,J�$��P	�)+vN6Utz��0܅�P/ٮr�\��v!�h��x�ȓ^��`�$5)x,�N8�f�ȓz� 8��O�]1l�RT"�39���ȓ{/������-��$~(�ȓi<ش!ĭ�_<"c/ק!а�ȓi�Y�&T�w�^��n�%4P��ȓ*�f�K�JB�$
��R�ĩ�ȓx?�W� ❩3 �.��\��`�Y Th.���)˯vD�ȓM��R��+�:v�Փ"6E�ȓz #U�$ut�A��7-�4q��S�? ���*E��t��Ś���(&"O�"&H�8��U��e)���u"OnQ�A��r<x�D+^�@:8�W"O�h��&Y���k��N+/���"Ob�p����U ro[�[Ά�[��'��'��'��'&R�'�R�'Ӡ���J<OT���ʗ/p�4���'���'t��'�"�'A"�'�"�'�4�Q*J�$BLc񧆈aR��!��'�"�'HR�'��'42�' b�'���D��'�� �1�u�3�'��'���'���'���'���'h�v��k��<"#��>2\�E�$�'���'���'vB�'R�'E��'�Dm٣��"D*����Y�r<�f�'���'���'>r�'���'��'&����
���`}�&�ȐF.Jp��'/��'���'e�'1��'��'"�����5`�P� �R�F�RC�'Z��'{B�'>��'ub�'�r�'@����k5c@�A�*�-5������'���'�r�'e��'or�'���'��)�ը���e��Ȓ?'�=�F�'�B�'�2�'#B�'7��'���'_dQWhV gg�0S�M��˂�'���'%��'��'Q��'"�'���AЂ��t��!�,�W�'{��'�B�'���'���'+��'u�� coK==�vlz���f�R�*s�'���'��'���'R�a�����O�Ձ��	{����rrgjm(*O��D�<�|�'*7�Z�-	�&z����g�8�Y8W����4�����'���]hXE�5'�E�~q���Z�;2�'�T��Ƽi����|�U�O��_�̜ڐJ4�pLp̑�� H�<y���D#�'*81pG:/�Pxz�	ҕw8T�3�i��$K�y2��A��ݪK�ISLK���hjp�D�+�P����0Γ���I��e=�6�z��4b��S�>�BsjI�6$�q!$d��Γ4�rCB\���t�'�k�R,4V2���kǡm���'��Io�ɱ�M3�j�d�Wx쁊��H�m� � ���hJ��{�2�>����?��'��	�H[v-��[:0<S�ޢ���?���F���|��O��K�?��B�萚�.�00?�,�MyRZ��)��<a�-D!g~*�[���=�>����<)��i[6�J�O\,ma��|:t�ˊ>=��r�*��+��ȉ!���<���?��O��4���i>����.+�� ǂ!&�t��d�I�a�I�l(�ĩ<ͧ�?!���?i���?�a�%hY`��ҕ#�r��Z/���Φ]8�ԟ�	���&?�	�Y(���F��
Sq̤2�'])2Dh9
�OT�nZ
�Mu�x�O����O�%��E�Nђ�á�|��e���]�\Y����^._�Et�Ioy�MK� a� Qr�>M�.E�0>���iM�H��' �̉�Lԇ��yf�Ѕ`��u@"�'!`6�!��0��Ąভ�4 M��jO� ���G��a1�H{¦��e�FUɢ�i��OnTДП����<��'UzkLA��1�%�0���I�	â**��O0�d�OB���Ob��,�I�OF��� �14�t�Y'c�:%y��ó,�O����7�J�����C�������d%�� ��\6���g�q��7�[��Mc�V����4|��F�O�>�"�i���O~qq�M� �N��tl%g D�BK8&6�4��DǄ�O���|����?!�G���0%�*�r0��u�0�I��?�+O@�nZ�o!b��	ܟ����?%�;nSԁY�p�����"$9�'b"��X�	���Qߴ)��O���'�.;tM[�F�R�A	�˃,@�0##һK����O��	C��?q3o*��	wj�2V�6*A��Q��.n>���O�D�O���<!3�i�T��L�<����1%�&��Q��P�	��M;�b�>���i<�RW�O��D�u��oe�0�Nc�moZ�p�½l�<a��\�pR&���4|#)O�<���$��@
�4=��`;O�˓�?���?i���?���)Ϻ.V��l�K���k�"���fpoZU�����ݟ4��^�s��@���3��!C-!`(�&<���%��#J�f�a� &����?���)�o�<�Q�ڧS�o��h����bX�<0E8q����
����d�O*��"6Ζ�j0��(O|9�k�a�����Oh���O���F�ٱ>���'���Y"Tn�hC�<?f��d�׌}R�|Bʥ>�7�i�"6mL�	�Xܺ!`�׵��\q�P�lt��	H!h�.*���QT�h�S�,%BgG���"�oL�r�9l��D��qJ�A9D��
�㛔H�p[ë�Y�tf���h��4>�$Q`���?i2�i�O�.�#�@��%�0 �P kƃ��Dզ�0޴=����Fћ�=O��D�"?�6,��'p#>�K॔/Xk�ȷN��sE8��pK*��<���?���?���?��j�-Qr�P��-J2���$��iS�L�ڟ����$���?��Iޟȓ��]*d>�tb���<��.xyr$rӐ�l��M7����O���H� GK�=�փ�@����t�N7-c�x�Z$���Y�UX�0:��G x�O��W���*2^�(�-���)C6<��	��M�'���?A�S�=_����B��J�&YKd;�?�Լi��O�|�'u�7-�Ȧ!�47��]���	a0j��v東&܎@Kr"Y��M;�'�B��iFL-����	�?�]� v9��NW4ID���AL$�V��t;Ov����(�[7��:V��@P4%�,��?I"�i���̟��m�S�5V3`�Zt$�"�F��D��U{M<a�i0$6��F	�E�}Ӹ����|cF-Ӣ�I�)�>���T+�Y��'�R�&�\�'���'3��'|��Aυ^�����.@�n`p��'~�Q��شO�b�����?����%	9r��q
*+rT|)��ײm$������󦑚ܴ��t�O���W$�p��qĈ x~tM���Z�q�M�5"Л8��I�?�s��'q�4&� ���[�u��؊oK*X�4hc+�ϟx�I⟤��ҟ�S�X�	Jy��l�`I�� �f��(���e�l�5��i$���OF��+���OL�D6��D���a�V�	�"0��O�'i�\7����2�$��-�t�����������I�?���w�T��N-C��y���@��6�+���O���OF���O��D�|RhBt4c���G��q��p���-f���'4��'��7=0D�<:۪�����1)�4)�@c�馉�ߴ(����O�53Ǳi��DX����s�˫C�A��J	�$ػ/���B�k�,�O�ʓ�?1�/��Y ��I�`��T�E�h�p!���?����?�,OԤmZ�d�T����D�I=�p	Pt�:CR�Fh��+e�dn}"�qӞ�m��y�鹳��
9D���d�b����?!�Cf���h�)�����e���;����J�a�Ӡ�Ǌ2M�&�ʙQ/��D�O>�d�O���-ڧ�?��*�%W��zB	Bp����� ���?�i��%�!^����4�?yO>�;�.�.@�VLt�cJX!��@̓(�6i�b�nhO�m�<i��;���S��AÄ,G�T
4��7<�T��s���䓾�D/�m<0�!�թ(��@��,YxB��'v6���u�b��?���tT��(MSG��8a�>`�K��+%d�'��c�r%%���?���%Bp�dS��61�$�#{м��E�}�)O	H���)F�A
q��h���q"N��!��{ڨ	Ζ5�n�з,�|'Z��&�7��<�SnEsךQj7#Jj�ѐÌ���4*�@_��!��͛'D��(��i!�$�j�BU4	P|����A�"�x6m�$]�R��VˍTN	���R7Q"r��Ƭe	��h7���]���+0G�4U��S�oC�`��(z�*^�o� ��C&#�ބ�����i�
Uj�A�-4�RhN�T� �7b�,�L%򔇀4�,�1��n��a�IW%Ae ��L_ DPdxUd�성���.'٨H�le���HrcZ.Z:�y�N�=��+�IGE�	şT'���Işh�pi�>A�?G(��2+���"s&�V}��'���'@�	�4d��H|r�#�~x�1�!�-P���W���'=bS���	� 
��!�/<���W��NVl%���M�����4�?Y���zA �'>��I�?ט?���b��<Q�����9.~7ͧ<9���?��EJ̧�?a��M����8�n�4.],sʞm뤉r�X˓(����üi�(�'�?I�'N����ȅ2���/�p�/�/�$7��O���m���|J���&�$BP#Q�s־Y)GG��1y6�ڥ�n��;f��q�	ޟ$���?��N<�'��x ��m�f��;x�ܴ@��iU�P��Q���Iʟ��3����@�Fֆb��� �� �!q㓍�M����?��H��x�&�x�O���'6�	pA�.J�F�)F";.�SÀ�>���?iEh@Y��?	��?)ËC	7���Bf��ȅ#��0��ij��B�7y:O�	�O���<yC-�=��M!3ZЈ���_.ɛ��'��k�y�'���'�剸v���Dd8�����X"-3�\��ē�?Q���?I*O<�d�OH��οL@lJAɕ[R��*W�+M�1O����On�$�<���d���"u�a�)��e"��\����ϟL��ៈ�'?"�'�i���Z	���ڭj�6YrI��%�y��W���Iݟ�	Fy\"�(��1ɕ�1�~H�u�_�Y�E����ƦA�	O�	Ay��T���O\�I�ō!+�@��V�T���Hش�?������;�)$>��	�?�����ʗr���Pw��NJ(jܴ��$�O"��M$F1�&��&�)<�p3��p�,Cs���MK*OrE���ڦ�۫�~�$�
��';��q7�_�/�J�����Uʽ�4�?�{b�I+O���?O���c�71q�\�ԭ�9��z�i��d�&LnӀ�D�OX��T�%��SwLL#�d�:-�@(�U�&8�4��Z/O����O����O��q�M�B'0�iT�շH����!Aަ��IƟ��	:�:��K<ͧ�?�m�����_�V!A��1(䕺V�����<��2��៬��p?y��T)4�*�;��Wq�|0@+�����Ip��'r�'��Ď8��u�1F԰>�I���W8^}�	�9�@	���5?���?�,Oz���
J!'�ǿ�򼸕(�9{"n�����<���?����'�rf�
AHJ;/rm���� �(� ����D�O���<q�.�l�@�O�(R�,�'�%Zĩ]-e1��ڴ�?���?)���'6x-���>�M��HX+�N�i1��B�X�FdK}��'��V��ɽ$ĖO��ŤtB%RDbQ�0w���Xʛ��'��O�䎼D~�ꅟx�略g8���%�&ҕ+ӵ�Ms���$�O�)��|����?��'C) m�4�0*E$���*T�հ�$�Oҝ�f��<1O���?dRd���=Kz(T�r �y��?��I�?����?����*O�� @5H�R$�$X%��A=�`P�X���	3?�����<�)�ӈ��ڵe�2Bi�X�AH0G7헡q�8�$�O,�D�O����<�'�?���TmK��C�!�"~�:E���<3����5Xw�Y��y��I�O:-�j���l��@Y�W%|�s2�S�=��ߟ0���=$4�����'���O��FO�!O�= q���[Gމ!th�~�ht��ك����'���O2�Pa���z�WG�b�I���i/r)R|������������=����{��]�������#ɓ���mX�lAQ~�'rr^�\�ɣ��D�዗��x|��Cʞ �NhA�pyb�'��'��O��dZ���u��x�j�m\U,�� �E�!��I�`�IBy��'3�xjQ՟���
!�=��i_<�x�å�i��'�"���O�*u�H�|9�&e�+i�XH*a�T�@s2�@��O�����O��<q�	�6�b*������:���놁zqx5)��66�,��lx�f��8���r�C�$Oz�YqIF�vO���LH�~$ºi}r\�D�	/u	���O�b�'���R�A� dۄFR�w]�l��[�9�Dc���',ޙ ����	k��ok���̚ m~ �X�|�	�UT�0�I��������SWyZw 8�������i��R.5�N<A�O�#�|`GxJ|Z���`�B��_)@h�a�#LK�-*�����L����t���?-�����'xͳԨ�,�`���ǋBn�yc�l�>)��C���O�2�;�z�#�',�Āa�ü��6-�O��D�O�sE�<�'�?9��~�(�4+��h�A��4^���ܻ[p�c��Sf���'�?9��~�Ɗ�Ϡe"�K�W�z��F���@�IN��@�'�r�'�$A*sșb�LU��9`�18V��9�S�3?I��?�/O��Č�;���y5�:4�0��O�$��!Q�i�<����?A����'��.���Zǌ��:.f�)7K�� ^�	�cD����OL�D�<y��rv�O�8ࣆAцR��`�⌵@`r�M���?����'x"�Z�ԅӇ�M�H�5��dƅ�-�I�v/�u}b�' "_��I�@�μ�O`r$�&.I�	c�ȺU}�̒2����7�Op⟤��v�*	bĤ5�$�nc�<B�했v��8��A�!��f�'��៰��dMw�d�'���O��`�q/8Y˚�BR��'!�|�)�	���
�b��/3���ї P���6�:Tu���'���� !R�'���'��tP��2ws�ɂV�(P�6���ƙK+���?�FfٯK12��<�~�p�O$-ښ���l̅o#�CǘĦ%�5Jܟ��	ן<�I�?����t�'P"%K�*�,!��q�+�&�L�#B�e� �C��C�1O>��I�`K���g�/����k�0<u����4�?i���?��#ȕ��4���D�O~�	�Qa&�zTI
�;$�5�\	CPe
W̓Y�������'�2�OR���B*E��d�c�@��3�i6�CT,Q�Iݟ���֟�=�e�S�c~μ�f�T�r�"A�E}��^8�Y�Od���O˓�?�B�d��x���vͪŉb�	5���.O��d�O��9�	ҟ,��� FT���EJ�m6|�7�OM����j&?����?�)O
��C g}@�S����ѧ�#o:-2RDPxr7M�O��$�O����ɓ-��2��~�浀��k��r��[�I��"�Y���i�7��<���+9��z*�����ӊjA�ԏ����k��; �iL����O6��0m���'e��e���A!З+v��ߴ�?a+O���X�(~��'�?�����6�9 '�Lؖ�8����A��"3�Ot��L��~aS��T?��a-ƋJg�LI�?y�墄��*����OL"aN�O����O������ӺC&Jk �C#��"_݊�B�_}�'�iQ��ϫ����O���:`��1*^@���̰8�|��۴���#��?Q���?�����4�v�DӁz��a�T'%�`�TB=/"8�mZ	cblSK)�)�'�?��XB��2�\�~B�B��H��'Z��<y0l�����'��O�!�ۿ(�TA�ND�]���B�^�,)�����'`R�Ox��Pb�oEB5�'+��k�8p1�i�?f���ɟ|��ן��=��mA�$������<��;d� |}Jۮ!`^��OH��Odʓ�?Y�ga�*1i�����`�-�Q���.O$�D�O��D8���4��ζz	l�pdF��,�u��O," �P`/9?���?�+O���Y�g�b��b��ȑk�(0v�ڡ��H6��O|�$�O4�@�	�Jij��6Ig�N�c��ʷP�\�S�B��&���L�Ity��'qji�T>�I
t\T��ĄʷNd�=���$��T��4�?y���'�� o���@��Y�VO՛B�(�b��Oi�6�o���'|�J�6R��SGyr�O�,���G���0�D����P��)���0vfЋ`Ҝc��f��m��-����㰅�:�B!�' b�Y�-���'�B�'���Z��ݘP�pUI�DF��y�sN��w�jꓧ?1t��0@�<�~�en�
��L*�H�mr��K!���{SD�/�M����?���:2Y���'S����I)��,��I%l<�qH�ai�*݊��D�'�?��D@~� zF�
NeH]�$nʇ@�v�'���'A�	�Po�>y.O@�ļ�� �ͲW�.C�:H�v�@$?m6A�q�i�rX��� h���?)��?�W��d�>� $��tG���t�C�D뛆�'T}���>	,Oj�D�<�����!b�J<�i�MJiz�^}r��8�y"�'��' ��'��	�Yx�����N�@=�"��4Ţ���"�����<Y������O��D�O�Ւ�F^*0c�+�&ց_(T\9#�W1O&���O���<�$�N�48�\&b�T�kƫu����WϚc��\�(�Izy��'X��'�PJ�'�ԹY��;MIz�[�톰x�`���|����O���O�˓|�L)�AS?�I`?� Yq��6X�u�pA_{�t�޴�?�)O���OP������W?���	�Qt���� �ry	����I��T�'~��c�~���?q�'/ 1�oƂb{�5zb��o䮤�Y���ӟx���%����?m"A�JN�T�(UH�e��%z�Et�J�f,k��i|��'���O���ӺKψ�%���ė�El���W,_���֟l8ala�ė'��ɑ�s��QP�U�vP� o�9m���48��7��O"�d�O|��G}}�Q�|�ToO1#��� D?���F�/�M�<�I>1��T�'㌸��>_Z���%�d�Z��p�f�����O���X���'_��՟p�Q"���Z�6wEBQ��THv�l�d�����)���?���M�R3Pt�Z�и5d6���e���Ѓp�PnZٟt�	����	.��I���(�oĩHp�XS�¶ ��s&�>!K�<���?��?����D��6�V��	0`j�󠭋9_��\��i
n}�S���	Py��'\�2Od��@m�I�D	���®=��@�A�"�y�_�����T�	~y��Nl���cE,�(и0��� a:}�&�gӚʓ�?I)O����O|������%*2Ԡ��*G,����5i�"�l�ڟ�	��|�	Dy�֣꧍?�10jA; ϕ�EEVX�)O,g��<l����'x2�'���D�y�>��ӝ(�*YUm��H�O����	��d�'[��ZT��~���?Y��Fw(��R@�G�@r�K�?��Y��W����ß�����h��M�	Fb� �6Z��HS���O�JtӀ�[�a�'��9�V�{����O����:tקuw/���f��3��LIbt�U*���MS���?�����<�M>����V'�RA��ꇽ,G���G��M�p!�O����'n��'��t�>1+OJ�h�%Րf�.��T��W.��ɈΦq`�u����@y����O�1�B_}>Lqv�W)��4�Q'�����ş��� \g�$C�O>��?��'���#g�6ddi�hoxR���4�?y+O@���:O�؟��ğēF�

�jH(�E
`_T��G ��MS�a0̀6\�@�'�2\�D�i�u�d.�����u��
���0ų>��
�<Q���?���?	�����rt����T�J�J0Ap
�5�L�0GXx}�R���Ity��')��'~��D(����͋��<ESz+�����O����ON�d�<���Qw��`��IcF��x1���KѪi��\�@��ky��'��'P䢜�5%A .���n3 ���$���M���?���?�)O�	�%��@�t�5�/���c��a�$�D���M������O����O�ݨ6O�'��-(�l�?�8 #��1B��H�ش�?�����d�H�ƙ�O�r�'����/*��%�6k (c�-0C�Q��?���?���H�<�M>��O��DDЏM �bt��1M��)
�4��DG.3�<dn��(��ϟ���9����2�����&=��xi"D5Y�6��`�i���' �Qj�'��<q����[)��Ԩ�#5X���"U��M��d�KV�V�'k��'c�䦪>+OH���ʨ��@F��4l�bF�㦁h@d��'�\�����b�����*m�y�sĚ_s��b1�i�"�'}��H�^Ԡ�����O��ɻ'T��E�&R�j軀%4J�V7�O��.��S���'Tr�'&T�p���7��!`2ğ3x�$�Ѐs�v�dN�,Mv��'@�ğ��'AZcFI2���W:z�z� V�R۴�?Y�cC�<����?Y��?Y���D�4Qo>��&용"��/u�Ba@�<7gJꓽ���O���?A��?9�!�.>�i#��4���Pm+3J���?Q���?���?i.O@u0���|r�H͖E����@�յ��=�P|�I�'�D�	�԰w!p��٢o̢��eS��Kd�8�T�J<����O��D�O�˓��|I�����l=p���!XnP�t�c|��7��O�Ol���O4e���d��3BK%�T>��b��E#~����'��Z��cmZ>��'�?��� 3d�gE��0b���c��L�\��Ԙx2�'�R!�*�2�|ٟ*�r��õ}�Ĉ#��ѿw�vH�s�i�I�r����4"'�����3����
7j�Z�CșG�@�H�V�'
��H��yғ|��鎋2�Љ�Z�'|�ĊcEÍb�
F�Q��7��O��$�O �IJz�	����	�^S����'C;7��X���(�Mۦ	P�<AO>�/��˓�?�+ݙq�l�#S� ~F�H��C�@,���'e��'�h@a��%�	��g#���4O�f����q�4���>�0�L��?����?)�ʌʞ4x��Ԫz<��IT�^�}���'�S��'�$�O���#��Ɩ�+" S�f%��{�� e���bQ��OZk��П����,�'5�Y1w��tS��ˆA-lJ�[u��s�c�X��C�	ş\���� ��u7�n���B'Y��P�NY�<q+O��$�O����ի�BL�|�lI'P-�Y(5J��S݄H�eAv}��'k"�|��'j�̆�y�����f09�h�vn6�k�@gÄ��?����?.O�U���F�Ӹ��x���!*t! ��|�P޴�?�L>��?9��J��?�I���Q/ĮT�l��tK�+4 ;VhwӖ���Ol˓y]��� ��T�'��T.����s�KN�+����l��: Od���O�`��3�I@"��>I�xf[��Po�ۦ�'��-�bj}�x��Or�O^�����Qs�L:s@�]�̙�-h�m�ߟ�����l�Il�Sܧw�bq	�8}BuQ��%��m�3b��{޴�?9��?��'	̉����t�!�(0K���°([�6��.JU����O��S�O��A�Т&JJepCW�H��6M�OR��OM�Pb�<-�����2�W��019	fڴ9�T>�	�Tلc���I����	�^>�����T6�	3	�P�x�ݴ�?�!NԦ�?���B���֟�%���m�\��arB�V�^t��{�́���×(�D	Y���0��ӟ��~y�,[5�n���'�$a#�iϝC��Xs��>)���?��?	�"�G:;T���X�Ot���P�eeZ%�Ҝ|��'6��'�R�'�DiSv֟
e���"�<�Ū'Cd��ҿi'2�'��|"�'����>��1�4�։3�Ys�I�C\n���'QB�'!r�'�cM�9�����5G5CD��5EY���Lʠ�M�����?���I�]���f�I�S�� sHA&�8 1��> �7m�O|�İ<I��)8����I�?�"��9������@�@�ި�M����\x��O@���.��T�+�@� @-ɜG\֙$�i��'e&����'�B�'��O����5.�1zԍ�	�]�|Ո��M3��?�7��&e�`�<�~���#� BvK�-W����"L��5!�b�ԟ���Ry��OA�)b����D���gě$:���abM&�VdF"9	r��y��I�O�q;@���t7�x˒C�o/0P�`KȦ���۟L�	�-��}�'��Ę�{�ZU�vm��;5�����%-�O,,��'J��'bo��+�b�GM9$Z�ڱK�'n��6M�O�ӕ�K�������x�i�E×���6u2D:0�ČVq@!{�K�>��oW��?��?�+OMʄ�WA�BH�Ҁ��r�-���$c鎨%��	�P%� �I�Xy��mR�Z�&�+7�) C�ơ:<(c����t�	韴���l�I�雕i��$������Y�4�?Y���?�J>Q��?�6dE}�%Dq� �RA�7$`���bG����dSNɸ  �"(HXPR��I��E�d  Nv��"��#b��"P�yb<�p�%�P6,�<e�٪�~B�����yId��,f���1�(���TO��TD��w��	�RD4;ۺt�(���r��e0�5�,I"j��1!A+�={� �E�T.�J���Z���	�IhU�q)��@����P�W,��am�,dk"�t�Y�,�2#���/!kХSf��m��L�'�O����Or|��-��,�F����ҩ&�S�/�4K��H�I9B��U���I4��O�Ԑ��C&ܘ;G�ǻ����HO�;������ɩJ٢t�����U�St�ٳe�L�L��q��/AN\�85�'z�6m�y������+	��:�,^�:
xmr�B.�y��'��}"�͏_d ���ͮ[vU2��ߩ�O� Dz�Oc��T����emH�k7+��Ĩ	���?	�-x��*���?����?A7��h�$�O<2O�>��H�Z�H��$��`ڟ�:S�D/X�v=�5,��8	��I�:��@CC'�2fi	�_�lP�m��jEQ�fR�s�bQ�#�?�=!�O3�U�1� �$]rSa�Q?i���ğ���V�'\�]�t유?b
l��.͐l��B�I8�=��@[S[����&y��{���?Q�'/�I�~ӆ܉ŭ6T��iF�O?,��ðe�OD���O��d��w[��D�O��S��t$
��E�H��I�T��i2�!��C�r=�����м{,�U�牚EIPa��`]�kdD�[�n�'UtH	1��-|�D�@����J���I�}����O�1�J5��u��� �q!�7ړ��O©ʗ`ހ%L�C�B&nu�u"O�"�%ƒo,����̥(�Y�1O���'~�	�/Ţ,��OD�D�|�K�bDD�)��X骕R�`C�!�^s��?��m\�dQQ+X9 d9�˞_�*��b"��[��[2�Н �Z�S�	�b�	ja��K��E:�&� Ԙ)JVa� C�%��bT�p�5�A�?
���Z�I,$`��$�O��?�!�g IV4Hp̑Q���ci���	sD0�#��/&R�P:�oV oxx��dV�I@�d !���*��Ūë��<A��I([���˟�O��hR�'}��'2�	6I�/Ԟ1��-W>�4[�!�Z����+�:�l;%�O�Su��d�d� z %��G��e��:Q岡yq(�
���e����t1u�����#|�-���OɓOK,hIc�R��x�JA�L����	Z~J~�J>�e#��>P�Q��.{8¥m�K�<� �%ɀ��(T�0��Q�E�32቟�HO��	�tʣ���̈r�O�B�	����pf��/�8��˟��	ʟ�r]w_��'ڰ�3���U�\�������'�}��B8�A��<OH�y`ʂ+f�� po(j�mч�O����Ë�kd�91��f8���F�]�p�׉(:���q',���R�K�O$��)ړ��dƬr�j]�������,9��=?!򤓯J9�aU��>�����>5�Ezʟb˓����iG����E;TWZ��$�"T�8��'x2�']B�мBR�'s����7m�O�P����%����T�F�FC���A�'���Y�(�C�Y0�Yu��I ��hqO>�O&�h��'~�6M��w��b�HC���� ��G�%�mn���X�')"��?��F��Xv*�	1K��AD�WB9D�<�f]�j@�(R�W�S8��i kw��S�O�ʓL�����i?r�'S哽kT6t�qÅ
k<��X�D9J7jCğh��ȟp�Wi�=B����<�O	j�H��P�B��P!��
��¹���D��{p�@����f�h*eNB�:�p�G�t�>�<I��S��`!ݴ�f�'�S��X՛^������5Z�`i�a��ߟD�?E��'1F���X)(If� 2-�?R츀���'.Hy�BK���u��	�8�+@�<�C�M����'�2P>�HVF�����ӟ�����
8����G�N�� �
Y�>�Yڴ�����	%�R-kQME�f�$��kľ*ά�I˘*�������	
3�d8�o�}v9w���0Y��0��'�����#����� 0G�N=�ف#%ȕ�bg��Igx� Ȱb�.(��e�p,X3d	��F�&�-���'>Z�2���*ת!
�h]�$9+��?��/l8t9���?1��?A������OPt�AH��e�8���o��p��G�O����g@I��{2�3$�)KV�T-rk�DL��~"��)9��-�ߓ^�&2/�#RO^A!2B8~��%��@�<��?1�S�'�RR����Y�%���ښh�b5cU*4D��ce�%��4Z$b�z��$2�HO\�A2��O�?��!��n�²��%��p�KY�2�c��O���O��$\-:h�D�O��Ӌr �ѳ��!�	�*���b��%=&p`��c0�OpP���Oa���1	eZ�B���"6ʚ�Q���p>y6bƟP�ܴ��:QCގ:�i�c�+��H�&�i/�R����x�S�t(��3�"Ś��*��г�&��y"�5W"�`�ի�/��h��.K��y�.�>1)O�iZR������� �O%���g�ͫ,����^��9P���yZ�'@��5d���B��>N ��d��6!�'�����<W�<�jO��\���Gy"F %��$�ŭ�`�<qە)�k��S�&�8��k1�$5+7�\ģ<��A�X���2�4�?Q(�@AY�G�U\H�HC�E!l=��O��"~�$.^x�3LD8����L�E�@��ɐ�ēG�$=! i�"��$�'��9%�����wN�(E&I����	��S�m���������U�lM2���s�n`�ƈ��[�91�/���
d(D�F�]��& �	b���.������œ�vx.ŉem�����i���a<��j��m����)��Vy6���ߩv��6B]��;&��L��3&d|��CO��B�e`B���O?��&i(e�g�ax�܋`�,!�d�{ҮI"��B'4t��*��T>+�`1��4�D��݈�n������`����=oQ����Obag*v���O��$�O�d���?)��;|y���3 �X��NS26}����j�|������ǰ=1�풦�^��N�(FXD�2,N?a��F�G����	ۓx������K1:$	��X�>$�)���'�������6�d��Y���ny"��37�(�x�o	�/��D:Un��yHS�'mِ�,�*�^Y��ެ7�"=�,�d˓Ĩ�A��i�T��WH��}f��KR�Y�["2lj��'�2�'E"]�6���'#��l#5a��i��+�?T� 9P#���N�2�'|�T3�%�>���Y�?�%{4`G#�m8�.���p>��Xٟ\s�4GȈ�R"��b/�(��h�Kw�x2��iB]�<�	U�S�T�Z�a�F5��� ��mâ!K�yrH�)(28 �IV�p#��Kr)���yRμ>-O�50��y}2�'�哭�jg&����.8l�ˣɋ�0������0����b��ݧR	�y�q��?�Ou
x���C����w�#��������3J�ه�u��ᴎŐ�n���OY�����K�*ɺ���mx=I��d�d��vX�~�JM$�9�`U2>��ɳf˅�<����>a�ظ>�\P�-G*�;���B���H<� ��9!ʂ&t/��a��*w5��>Oxh�@�Φe�I����OR���'���':^�Z���`�4H���¬Q�4�O55�В�lνh�,H�FB#%C�X�'јϿK�D� ^긍S��)0�z�8�@ϟ4���f�,a��!#Љˎm�pP�ۘo��)b�JX�	����m��^�T�ީ����)o(4�kF��&Z�<���O:��?�G���g�6���G�:!�8� d҈^gt��?i���P�E��t�v�Z.E5J@ExRG9ғ��I�6Er.9��e����A*W�,4f��O�p�Ƌ�	U2���O����O�E���?Q����O�,m6X{����؀��^�*� P'ֻ%Ҧd��I
tbwiΛI@���䐰+��I(|�9qd�+�`��$Z�hW�H� @T.FP�%�w���8��D�$:���!y�t�'�V�����@�O4��M��^',���?D�L;b�X4$68�a��5���'
�HO��'��ӼK,���~|苕\�
�Px�<IVg����CKߎK��"�u�<��i�+�-@�k��ɠ��Cr�<i��U �\�3s&ǒH��`4F�g�<٣I�wj��lF��@�5G`�<� ��09FL�'qF �#aB�V�<Y'�O,���N���C�h�i�<����.}���I$c͗|���v��h�<�EEJ�tLr2��L���$T��s�O?,Ra���aAj���7D�L��H\;[1��J� 	���L:��4D���_r��xP��	�~���2D��-�18S��r��F�0����1D���j� ���jG�r"j��A-;D��С ���2� ��	i���-D�p��ꜳ��"�-C-,����b D�D��M��sD�ȗ�I�1�
!D�|:�@/H�f/�bBl��->D�|���f������%ArL�E<D��c�JO?������ u`�`;D��"֋��x�䥹��)T�4��g8D��ۆ��`�a��Up�f9D�L���Z)y��(*�KYi�9��8D��iY�/\qwo�`bUZ�G6D�T��"~�tU�6�;ŋ��5D�l:��#|� �p↺C�����b'D�$�0E��B�IvF�=\�Z���:D�#i�="Ѹ��ŮoT�`Q�5D��ȅ3A���EĠ'C>*�2D�|��1��#�vv����"#D� 3��!�ש$�xh{'!D��k���o̰I�'�я$g\�R�%$D�x�7͙�)�-�R	У�z�0e� D�|�:qQ.9���m�4�IWd D�DА@��p���"$��J�S6�2D����m��
5t��G�@/z�޹!�N+^_�	�TKW�?��$��OtܼqGB�輓��\B�*���.O�l)jT��md<���L�F��Z�)n��8�2 Y1yY�]�OȈs�mP�"r���Ԡ�K��"��� >����F;���#��yax�hW���4صE?YXDl�� �+���е^ =\ܘ�jZ Fu�$.��4��խ+�{���8����	�����ӹ���S�O��؃�!Y�7ٲy�e+�U��D�?<�u8-��$0p�+N�� Q���Ke��+�"O�U;�E��0�RCG
�B ���oJ�'ѤkQq���h�0O�T9�M�|�ƪ  te*��;0b�]L�:�J]1��ƓX1��p�\P`����[�æU� i�Q�_�<�p��q ma��Y=�d�	��Ow��b%V� ݁F�	;"fH2��0<��~��`R5K��T�-��""x��&@f���"�$K-qG� c���%��c	��=Y�b�����h�\82����D~r���Q0`E��McD�4�8��X�'�x����O�2aKpO�8z �<3uΙ#�!)	�'�;��
.�!�����OJH�THڐS�����
��蘻4���~*�6�s�aS)i�n�*(���R�'��[~���AY��D�~�����̘��#?���	;d��Rm�xuZS���~�����Fc?���ø&lT�yaΎ=r
Lp!�֟�i�NU�Wf��=� v�!��چ:���2�C1/#�肂e�>��O�l��g�k�<�6J�h�f�a��K�l]|��k�`�RUJ�5l�35F�$�S��O��#Q��C8Qg��~ʟ��&$Ї z<��)�m��[���x:#Bt[���wS�%��H��782�7e����G0b�L�TMU	1x��!H�dW~!��ؔ
UT���ڑ�~��9O��)B�q�=ID�.��$��LA�"U��ʳ4�qO���B��Ũ��F7���b��#5� �̓Z� �#�K��h�L=P� "�,��jcO��4@Z`�F3y��,��h�Ē�&rX�[��3�i>Q� 	U��M�waWY|�R�o�.g��k�"X�9�v�>��W5~v��v�ȝF����]�BW*�ceF��L<;��I�b���FxR�'��tGʭ�<9�Oz��(p�Қ���r�gD
/����r�+Z���'���U�48%��0���J�{�'LJ��!s�È>�����/�Z\�6�.����O���	ef�;�iT?:J����>ٱfj��'I6$(0Ѭ]k�{d�ƞ_���>�{�'!2(ps�A<�=G	��^R���'W��͑40y��-U]�'!2)r/���m��܏u�t�`�E���I��HO�i���޴Y�v�rR��Jo���Fb�A�0�!c'�gn����	-�������'؅9���
�0晻A��J�Xs���<�>���'�X��K���r�Ũ�6lx�*?**�ϔ�Q��I*>�T*�E�	?#@��ɦM/R➌X䠚�6S�%�j�2�: H&A=��_0%���p�R�Y�iu�s�L�����O��H *F�o�45Kw ��VD�))�$�D"�DC�4���Ob5���ɏ2����`*6/v��j1��w����O&B@��oߌR�N!{3�'�Q��B�3�Y�q˄
8��)r� �q,5;Gg����$8§Yۄ%y°KP���MԺ�#�B?:}���	��p?�]	N���-ʞ�J#�ʱ �'�<3�NT��yB)�0^א�������LJhx:��6�q�2/D�t��f'O\�B��x��x#f��w�<���-F�o�>�+��-�hr�c�5��䂹fp�@$��*���'7E�ämF#��Ufx�d�5S!n����35`ܥOB� e��g�j����W���b��I:O�a(D&Y�Z�����JǇe[�����!b+*t}Z
�|�,��).ˣ(P�=���m��  ��"�͍71�贯�xxb��?c��R��,#T-�UDZ6,�N�ڠV
O\a��M1`B�Ud̵���+w�h@��'W2U�?)6�'�ؔ��w6�q�k�68q �8pN.
��+
����S�Цz.l9�tS E���#(�6G�\�T�i�n`�'�69���'6�I��!�����`�S�d�H�8a(S M�0d]ȳC�ENў8�����B�"�&���҃j��	���U�/��<�`�¬�{6���a�7=rps�K&oLjX#˓Gl�h"� ]2'����
7� ��'�N)S�'�U�@��8Ĝ���'I �s-�x�ӂH
D�B��d��	6�qe"Oܝ���ʖL�4���|i"���9X�m�`�Y����6r^\b>]�$ɇ��N��Rv�D�k���A�D�r���';� P0BP�1hn�sT�]n ���2e��	0����@�;�3�	�\��}�RHH�l�
A�%E�o�1�a��l��2� 4Ҵah��)�'y���t����hf딓=�� �D��;S��\�#��9�-�~�(3
T�5����Jv>����wF�(�� [bQ:W�ާ��Tb�#ʱC4)���ɡCe��`���������>x���d^������r_R��T����\���c���p�U��A��~��<�w��;i~`�F�G+DȮa�ԑ�J���'����$�e D�á�Έ4���	�&��'X(KJ@�2�K���I?m����B��##��Q8�	�#T:��Ҕ�V�oD�<1���X #�T-Y��E{¤5)�~y�蒣#��u���W�^�ZQ��%[>xvcL�<)~��'h~x����c?�t���O�>��Q����	[�v(��N#r�ؖl
-k0�"�T�
�P=��#oÄSFLX!�	�r�+Q�<��mզQڐ��d%0����!k˔<��M[�	�m�b1ϻv�a��"Wi�TM�0��K�����ɤAW�y�5�V~ʠe��J�:�"�S�U5#��x"S&4��/)E�U�3�Пa���>z>"�Q�E\���z*C4H�4�QVēn�"s��82:^�ل&.�{�Ż'��%wT0dbfnJ0�t�ΓJ�y���[?�Ɉ���$~M��q3��Q���?K����0_��d(c��/4��㟰2��� M��A��(`�Ip�,c�,(�4�i���Æ��$wO� k�@��;h�����ر��K:N8����pQ�5��% lX	C�-1gZX�u�'3��#3fV ��s�)n)Iڎ�Yo�ϓZҘ������������Ir��w��u����zR�xr��>v<��a�tg�����f*l@�?6f�%�A(׸{ �В�j]`6
��9����U1��?�卆k��U�ΰq��(cs��6HQ�p@3�O�y��#<�0���%�AB�˧)�)�nH�<2� 6tD�<�T�P�g�Ltx䊂�s���=qAI�ٟ�!V�цb�<qc��C��'W2�k ��w	�ً�I^�2q�mCw-C����9��\�h���y��������T���w��X���@$i����쓩h�n�󵡝�M_E��	�yI>����V�џ����o�z�`Ȝ	]��a���-۾�I�N��P�;"�8�ɗ7=��q@<#!�ᣃ盘+s��·
C�\����牸k󸙀7
B�X��� ֑���͝7�q1�	<�`���n/��9W���V���sF�?���8mƱ��A>4��-A2$օ+�|@Ä��(O����P<0���$ׇ/�|Aǌ�|��#27C���e��1��p����!1�ߛ>^=��%�,��pG��]���t���E	J4�$��*�n�`���
j�X��T�bl����,?8�D��w0��3��!lP``Ѧ�No��{���q�:�	$R�������џDradEM;L �%D-f[q�BOW�Vuа��$P�B�`�A1G���S��&F��`��(>r@SAi[ed�@�0�_0�y�g)��<�4�	&��xͻQ֦X��b�W��0*��A8|_��ae��9��]s��b*���ۏU޶x�7b�W,�1(N~��gٶ�f���E�$o�
�{(Uu�'o��b�ߒ-�&���	U��[�dM_7B詠E�T�D'��ig���&V�tѥ��(�X�p�ɼ6ƈ�j��ɨ<C@-�iq�&�%�pU;�lP��Q�
�6�\ DG�cL�PE�D=O(���H֛s� #& �(Ѐ�5�©d�;c&� ��
(�(�?���� ��0�j�t<����H^�9�j�f!c*F�I�+ٯX�D���~ʟrҗaϥn@����'N����&N>T����6T�.l^����xyPt �����s���7�,!;C�;O�Qj�j[7��y�Ƣ�x�t�B�[�S��p����t��G�ӏ7ʡi2��)����0�ӫ%B�b���b��n�F�*���$4�]�B��P���R��YBh8N���2W���V&Lq)�Q�aƠ� �3�yia�Qy��Е�84�w��)u��s���\;��S�97��P�������ɾ����ɪ8J� !5(K�JP�V'_;*A�����2��� m��.��Er�Q+;�z�(�/
�wkX��"E��"7����z�1y����k��h)^w-��Ɏ� ^ř���
K�(�1kF�"tI
��@|8�,C��֎]��!��G1Ĝ����_��TH�	�,!0�K����/̨A�a������J���'u'�)㠩��`ؖԉ�L�8MX��d=��#o8#���:�@�/�Ib4<�����~��w�3C�T@����y���'6��D��?����90N�I�<�U$���'y$���S,��������o�<Q��*ؿ}Er��}"�u�i�2m���;^$�����?��ő"#�H���A���{��a5�H|�$�fn�x� CņݎN�]b"�W�)�f��C���̪)��~Z�?q���"��DT��Adn �L�>��ǦQ��
�m�z����NĜD/�E�5��E�&P�b'�QKP�;��_v�2�:�g���X��Ϲe�a�i�)���ij	2�
D4z��I�ǀƆt��1�}�)ͧ|���BTY�Ĉ#�#Z��U)tX�Dں)�T�T1"��AZ�J�u�dK�"��䁘O��IY3ҵJ^�'�D����[�lC�Lʫo��#)]6J�� ���� @�����!��OH��韢qzW?��|�B��GSF��s�ԮW�pd��7l$�z0mD�|'ay�aK3C�"�PAJV6�R��%%
�b��53@ �,Q,tDQ�%T	Z���f�`�+���?і]��i�G�Qp^� ��� iEc�&��y��'A/!kAk��T����!Vr̼��ϑ,XRB��4��<1��2`H��'��ҧ�s�|�(p�Ya�${"�
�YXs��]�8�֝�f��'�<�C����K?�ʆ'DwG�( ȓ��R�@�$�[���%��sӎaS(�W���'��=�o��8l,�P0'�{�M��!ȃ|p�I���/E󒉲��$����ԟ^���D�e��Ө\�QM^�\��0�B��e����	��R8w�ĩ����a#pU�Q).�30�N���Ï9X���S�,O��'���%&�q��0�D���%Δsb�i��H���ǲF��8�][�Ș�G鏹:J5'��~Ű�'�̌�ԩ }��<%?7�T58��s�D0mlD���H	2dB�ɿ'���`]���,9~�
B�	�؅��TY�"�R4)�/ly�C�I/'S�|�$LT�1+�!��r�C�ɐ,gj�[�c�5S��X�Ȏ�BdB�'fc��姟x1��SI
IBB�ɺD}�QY�d	� u�WAS4�B�	�XM%�K��T��%�xY�C�ɻ!���
Q� ݰ1�����q�HC�Iv�T"ch�,=�����%"xC�	���v������ �B��'I�6P�w	A�:ʰ�,S,?�C䉀j"�](
K.	6Ό�G'
A�C�	1�P�F@+t�����Gʛl�C�Iɒ��7ES�A����M 98�C�Ɋv-�����M�/�HHq&&��b�C�I'x�@�T��e'>h��l� +�JB��<_NUۤ��:1�:p��J�i/�B䉘~�r	���C�9�ޡ����P*8B�I�)rX�����~�U��i�,��C�	>^�Q׉{*��%/K�g��m��S�? 2i�" 3:KN$C�>LL�;�"O\ c�b�V��"�ؔB�h�"O�8����\���j����"�6��s"Oh0¦�=��q�n�D�"��P"O(p��D°rx�p�.��-h�RU"O����*�J�DA��$	��b"O��h���Kw��ؐ"�@��z�"O� ��H��@[��WM!����"O.�A/�Z�f�ۃ�	9`�(�K6"O6x�#N�5�l(�S/à-�ѕ"Of䘅���f�2��WG��*�b�s"O�:�l�M΀hdkC�H��P"O��rcE�V��H;ǇIX��"O�=�n��6�U�q�^�K@�Q�"OT�� f�_��E6�׌[Ų�R"O�T@�+^�7�Ԁ�h^.t���""OʅbV'K�F춘�h�<:����F"O�@�-|�D=8M�B�~U��"O�}�P���I���"��<�jM��"O\a���l�y�ҊD� �^�*�"O�m�LT ش���3V<a"Ov Y��ՐBk䕢�,��8`���C"OrX; %� S�܈��k�R��R"O`�qA`��r&X�k�֝>5<]�g"O6H�W-�$@Qڙ<"�A�"O���ä�uX`��i�qٻ"OƤk��J�D�P���(�*c��"O�hc��5k֢��ԶZ|`���"O�T�5"ٽi�,�9�/�7Ax��:�"O�ز0J�������ɯxB&@b�"O�t[�ԩUA������)a�"O��1� �'�Y��F�O�l�R"O���c�O�&r~(&�Ǚz���B@"O\�����1,Pa[�Jײ ���p�"O�$IЀB�/���T*�5�
�Bq"OtH���D��1Y�
�&�j��'"O�x�H�dB�R�����@B�"Ol���Y�?�@�� ,�$@{�"O0d��i�6 vD���jR�0��"O\`��#o8��!-ѧH�<�w"OޜK�S/�w%P4-�>��V"O�D{C�֯\xH����%��A�"OD9x�O���8rg��oo�d�c"O��@��0����hF�8ZE"OrU����ܸ�׍ɐiE�Y�"O���lmkX�u��#8ˆ,+�"O@�bH�6 `�l؄��?�^�"O`��`�Z�$R�񵅎�(���$"O�x����}�Jq����K?vA)�"Oz@����cH�U�Ҟ72R�*t"O�$XpH[G�x�� ��0��Hd"OL!k&�F�&f�0��!���
"O�#Iμj��M�"�ߟ_�Re@@"O��9�o�Pr���$kԎ6� 5��"O̩[��K�+bش������AG"O�)k���8]4���	�ul�l��"O4=����s*�h凈����#�"ON�Ia�kؤ����,b��x"O����΄�nW�D�L�"{����"O�Y**"Zf�Kw�(m"� �"O2y����<���"�Ǆ�ԍsE"O�Di�.�c�\(��N�@���"O��@�aR�^��bBŇ�:;<���"O����)<9  �v%�/�2Ui"O� <�Z2!Go�]�&Ҵ��9�"O���#�2e�L�B��&	���X�"O�X��
3(��IAo�\��ܙ�"O�e��FچK�&H"U��&L����"O~��@�Ž^A�,+᥁�h6ܤh�"O���j��>@���_1e/���""Op�r5�a��Jr����0JP"OB#���)u�J�*����]�:���"OryP�
1$�2��t�K9q����"O`�;�܉&�@�
��	Y�s"O^�0		h6D�F@� a���Ir�D�PC$6���D��5P��;$�0�PAӧ@N��@3� "%6�*0�E��y�I0r[��s��@��F��)�y��S��$Yw�Ɛ�rq�dϏ�yԆW2xl1��۩cr��ԊA���'ўb>m�1&�x��Az��u�2�a�<D��X�e TLvpa�$��#$L<D����ī-�4�7��-������4D���չiH.��?RR�P�D�3D���R�@#��U� ʋ�d���X*=D���Uc=;� �j䃉*yI�A���:�If���'z�:��D!�%��1w�lU+9D��c%Ϙy��a{a�Uj�����$D�p2�ǈ�$bly�GR#W�RM`��"D�@��,	�fO���"(�/<Ն5��!D�����V�$���n�6I��V�C�	�kD���<S,�Ca�*-�C�ɞI�� z����r^��dM�
DVC䉬CR8P�E��NMdA���;Qt��d�>�PJ,4����p�F9���G�<�FGܖp	�����q{$p;LEB��~�f�O�A��c�&\�넨�Vi��'���A�`@;�^�h�� ���)��<a�dEh���YEO�J��,�� �r�<A�b��H-xe�eE4���f�_k�<f�Ɲc����C��wĤ�)�e؟��[��a���E 4;�#����h�ȓp���S
��M�2��b&X����ȓf�$��M$'��4s�lVr��Y�ȓ$$�sw(%�Pqzu�֋!�A�ȓ?��k�`�G�Bu aD �b��Wa\S j�Zz�bD)�2J�
$�ȓ2�̋�E,[6�dJb�/^.X��l˴H��ݸtLVd*g��+t�d�ȓ<�H�i���:*I4p��-c���oAl�� �
6-�P*rZ!v �ȓ�r���I:n��])ak=J�Նȓ��D���P���e�@;?�`���I�<A�O��C\��Z�NW�eS�]���Gf���=��ZRN�(M˦2�X��b IW�<�d��#�1��	����Re��\�<A�jV6N��8�U�@��]*'Rt�<�p�=T�U��)^�<44��Xl�<yDR���5�'���\*n5)F%�L�<���}`^8���z?hI�Ua�<��޿[l*��E�g7�Hg-�e�<y��DP=�! Պ��&<�P��c�<�"�ݛ >v<Z&�)%���*G_�<��/����h^
�F��0KVQ�<�e���)�L\ɒ$
�AU͋A+v�<�S�)�nU*�ȋ�����#��r�<Q�덛P�b ��P7$N�ZR	s�<9�V �T*P}ҒA����V�<�  � KB�92�q�7��2"O��.�TX�<����1=��xca"O���I��A�<x�"a�n�5�g"O,i�g�Hv��oH	t�Y*C"O$qU�{u���7�JcVQ8G"O�ը���N��EF�n��ihR"O��+�+�=A�ҁS���1�v,��"O,���i���<�b ��B�"O���i��R�8� �Gև1�\�s"O��S��>MH&`zFF*i�6(k������	41� μM*f�!2
ۋ!R���$���c��}2\V��1.�ƍ�.D���5���},+������<�B+'D��ɣZ*: t�f���{��0D���Ѣ
� ��G֫T���em"D���@�4)��8cU��h�"$cD$D�Y�Ñ|���!M?a��sj<D�����9�Ç�a�ཡ�/D�,b�G�y���ĥG2�3#2D��JR��58�t
�lä��#0D��)s%��-���Pa�s¸��G+)D�x#�A�'-��`a����eif$D��JS�" ��L��n�ʁˣ�yR���g�Eq$ T�n���Y#̇��y�?�*!`@FN�`W>a�nՀ�y�����RXQ���Z�6���b���Oڢ:P�/�"�`�i�)%ڌh��G�D�<�u$����I��͙G;0T��X�<a���y�Zu�6  lzh�!��n�<I�oîA:$zl>�ai�ek�<!3��+�X�7.���!��VR�<�҇�!&i"t)VD�irX�Y��Cz�<�4��z\ƙy�.��4�JABF}�<I�D�itLi�I��f��"��O�<y�O��C��a����e�����D�<����]-.H��L�	ݮ�j�˗B�<q1av(�C�$/Th��%�����xR�3���h%e����+1����'��z"�	�6��%	-Ͳ}JJ,['�T��y�� �y���`��Ͱj��M����y2琕_�|}�`�L>j��I #�ya�3겤æș�iܘтK�����hOq����лX@����N�%�LqZ�"O�q�����؊�nD?���Ȑ"O"�R���z�!� Ά�rʵ�W"O��� �9|"�͹F�Ҹ=G�Q "O�i���B($j`댄C�X`�"OJt1�^W=HQ�i5;����C"Od�� �;����p$D9Sb"OZ�3��0�>�p�^�G9���"O���D�
E���O�1+.�u"O�0���=�HIJV��1T'`5:�"O4�r&��J�AaOI?(����f"O�!�ƤL�N>��d˖�W�6M8�"O4��i�C��Vk��L��Q`"O"-�����QCP��i ,JTH���"O ���jQ��L���#_�<΀�"O�Lj�FA2T6���@9F�r4"O5`�&��,	���o�3�Lд"OPZ0J
�R����D,�+E4]�s"O���P�H�27[��m�B"Oua�\�l�hkv�e�X;�"O��ɗc�!����ůN�R���"O��Ԧ^_vh�֊C{us�"O� jI�@�X�j�Tl(��OϖA�"O��҆���J41���Q�ڹ�B"O��┈`���˒˃%C��e"O|$3�C�(�43*إ}�8m*�"Of%�"c�*{��|���zؤ% �"O�����Q&���:��_�	�F��s*O�ɡ+�.n����R!�Mx| ��'��b@�f�"1�͏�O�d!��'���vJ)'�A��C��A8l@�	�'v,QA���q�p�R�F�%;�~l��'GHH2�	@xn�A�@�5�ء��'�����5C؜ ��+&����{��a�>#X�S�l\��&<�ȓx�
 C�ag�����Ϯ~�XɅȓsP=�W�ȯz&9+ �ƧA�0�ȓB��hd"]8a����ٞ}"��ȓm�~���٦`����Hn\�ȓ&HR�ic	�w~QA��	Zf ��ȓ��&m7:4ɐ5(� �
	����������	��d
�iQN���
u
�Y�m\�Z$�1���ip��ȓBaf�  ��O�zU0ၔ*{�X�ȓT~�����s֌���-��mw&D���^���i�Dɒ�{%k�I�؇�T�,`�,N�>l4�;R�(��E�ȓA� c�߱T���!i՟E��0�ȓ"�|�0�Ϳg�9X�N��?��,�ȓdD�87EH�_ppi��%�����C~�aԨRd�d4y��.z̜���X����پU��X׊G#8�ȓ�ps�Ξ.IX�h�D����ȓ-�4�m�%
�,��N��%`%���Ԥ�f���E/�m�XM
4�f�<���bf\���-��	��хA�X�<IHҼ('>����0x�4���X�<	��71Z��V�_1��l�"�S�<���ҠL���M�艱fQ�<�1A<8�`�l�6a�py�jK�<���	T�ܙ���[�K)�QfEDJ�<����P�����ުE԰hJ'�D�<A���`�[���>]n��C�g�<	R�T�}��Xc]�O���
U^�<Q79Tw��0��ȱ*�����<g�[�Gx�܀��	*`/F�R��b�<�M�l�S�^�,�5:�I�<	�E^�(�h��U�L7�6yA3�QH�<I�+��, f�/:I*х$�Y�<���U/�I9�hK'uվ0�3�X�<�䁋:�&�(���>Vֆ�ʁh�K�<�P%ݞ/�F��S�E=Lr9���B�<���#*\|@DJ;f��12֯�C�<��?�e��"�7
���a/�C�<��D��4��
�Ǵh?���GJ@�<���1�ƨ{�̆�$�|��|�<�@Ȍ�4��9�M��̂�H0�|�<��>1e@`/�	[�0��"Yu�<Qw������p��0��Bt�<y�E*T�^M��		h	D��U�<9��H�p�cgŃT��2��B㉣'���&mغ15L`� �W�P�C�I�\x8C�/UT���Sg�Ò'��B�I &("�*c�@#A��)�(?o�B�I�fN���A�B���{f#�-�B�	�6? �tՇ��� �(�+h�B�)� XА�O�J��d��0� i��"OD=�g�'L(P�' �6���""O�p��&l�vd���#I�!2"OBaRÊ�7u�,cb)�X��"OąH&*�01�y�qnJ7,�m�"O�aa��ه#�4� mW�o���c�"O�ZWF�6R����F�˺0��"O��듫5}� 
v�<r���;�"O a�@JuN��Ď@�C��-��"O�9uJ'�تӂ� }�0�"Oz�B�ߚG(Ju�R�C�`o�p�"O����j]m�ඤO?-k�"O��t�b���z墛-8���*0"OL)�PL��f��*��ʇ&M
�c5"O<`���>4]*1� �Z�h�p�"O�9��I�8ǆ����"2�����"O�AA!�ko�m�wL��P���!Q"O�]���C�0��+U��X�"O��i"�U�L���'�U�SǄ|y�"O&��v`M�D��kȗ
�FI�"O�	#�i@��mW3K�Ȃ#�
x�<���>4�8��f�+wb�ɫ#�Xq�<)#�"��l˽&H�5il�<i7��)I �L;|���)��S�<�5O��eo [�nzK��0dDIP�<���L��2��,E�ᘓK�T�<��&�0x�)����*&��U΅S�<	��	%|	T�(�N�%fKJ%�f�z�<)DĜ�n�J�9��VȕXp�u�<���+>���2�lN�;:�{�@�u�<R�ͱ�Z��#�T+S�
0P�mr�<�`�Ӯ1'��(VꉐyW��d�V�<�e�!G��E+� [m����m�V�<�ׯ�3x #��sK
l{��k�<	����\k��Pm$����Gj�<Y�ۉ������k�����i�<a�ܸ
+��)j�6@)��Mh�<Q�`�aܺT
��.�P���`�<�6�ʽ=r<��[�lc���aw�<ɠ��,q�qBW�#u��G�Jv�<qЂG�8N��e�	/�,�1��h�<�  p�Ρ���ɫC3�yB�"Td�<ypE�5"���T�ȫ=F�h"�Lw�<1��E��f%�V��qE^���Lp�<�C�ˣ>8�rGeH�T�촨֤�m�<��9b���A�
�I
�����N�<�h�+��C0¯.M��c�d�F�<�i�6[="�x3m���\Y�'aOw�<����#D�����ؤ<����c
t�<��J� @�H@���#N�D�)%�p�<��L� %�,�"o�͒���'Ej�<qvř.��j�j�N�0�F�Ac�<)afN;;3&���튝��X��G_�<	�ʃ�
�je�¤�4+����[�<)q�N,dz���&1`�e�T�<�3�],0��	��E;Z��	(A�t�<1�1c��0hB. ��[���G�<��%�8V
������bP�-��lF�<�ӫ]�ab���6hO�d��h�<i���S�`s3	�.FXȐ�JE`�<郧U�V�s�G�V�mc`�<1d��1\P�ĂtB%zd�c��Z�<�×�8~��� �(�B�9��V�<����!1�=�a�i�Q5�U�<� ,dQe�_-I�	��ₖ#m$	�"Of�I@ �;0kNT�UB� M\|Thb"O�l;���7���k�A3pM�}�g"O��Ҁ��A�QJ'Aؒg96���"OPx��
=,��1/�2/#�� A"O����W_6��E��:?w|s�"O
\b�*��e#v��5l|mb#"Opx!��,a�DA���&K���"Oطw��A�~��6���2x�:F"O�H�G@_E�,��0'�!O*dE��"O���P�J.sږq���� &$��cR"OUCW�Q�B�pQ1��D;H�C"Oj�i�'9�~�SA#Ɯ]�;�"O� ��	�%>�h�ȱ��w60I"O~ ;ǉ����JM�O��k�"OzpcE�$=���)O���
b&��y��P�7���2Gx���+�D��y�C͔Ea�8Z�#�k�r5C�E�y�d\3d�,��@T��X3��5�y�d�.�K��F�J�H�aE���yb�Ъ-���c�bA�3���g���y���z�@��e�4&:�&���y8mrz�@����	{J�D!�(E����b�֗	A��#$��~�!��^�O��`��¿q2V9
�i��F�!�IsM�B�U�l,0�*5G�Z�!�˝�N�hf�D. �H���Ĳ_�!��9�x�`�*���\�!�$�����N��9JA���-�!򄌆~��e�Tci����ߙm�!򤊐y@Š�˓�K*ъ��X\(!�H'H�(�W ��S,�\�)ɮb7!�dJ�8ؖ�QC�Y�N���ұ)�	O�!�ǹ3T$�9���T��K��D�M�!�:\��(��+M�Vub8
'��53!��$=����nƟOg�L��Nޮ[�!�Ym�riX���/Yn�aϳ}�!�$/#�h�9WMX&RQ6`��Z�b�!�D���	Á�2A����=|�!�L�|5��/4�&�;hO!���x`p�@�
��\(P �)2!�74W�t.)$F�Ņ��%�j�'�j8ã(	�* 8��#k�ܭ��'ڶ,c����ε%Ŗ�q��P��'�rhe�=����E��eu�4��'}�����;��;���Z�����'��,�Ū�gb �KS��YΚ�Y�'54�@+�{�ve�b��"R���'���E�~��DQrJ�v�qb
�'o(�g ؟s�������l>�	�'����'A�'jU��@�X(�	�'�^��Ёˆj6.���*x��b	�'A W����!�rh�2l>@A�'���qoE����(_�Xi`�c�'``�Q�gG�N6�u#�!A2���'��@��c|bq��D�4�FU��'M�L�TF�4P��:��6wt1�
�'C��3VoȦU"��pcQ++.��
�'� 
���
����ţB�{�-H	�'�v)�"b��k&��T	D=#
�'��ࢷ���[�/�9J�\*	�'��R�ɓCTPۣ�@�DL��	�'�����	M3c-.��g�Oq����'3BM�@�<M��p����sJj����� �a��m� ty%\h�8!v"O�h3��J��<��'��׎y��"O���霆k���;��ʟx�D��c"O��S�&nt"��0�ҿ�L��"O�9�� �|( ����n�@�Zq"O��" JW�e�ɐ�	.����"O ȸ$$����,���(Ŭ	KA"O�ܘ��N�	hv0����Mju"O�r`�R2U$������Z�vq��"O�01eօw��iR�ҫ	�q�C"O��Ӫgb�x�*��"NE�"Of�-߽g����wiD�L�𑨂"O��j��|h>�	�G�0/"�*�"OT1�J�n���F�.U�q��"O ����s��\��b�`�\���"O��;��zc����@�L�"O8%��aԀ7|Թ�$�-��]�3"O�fb�nq��r��
��H��"OH�J�G�v��ʶ��.�����"O�cMO-f��"rꖏ���z�"O�p� E֚<���R娖�ou`	24"O��O���9���2>���"OL��vV�q�� 3(C4�-P�"O؄+v'����� ��4�0{�"OB���Eb�<䣱�D,�D�au"Oౠ��3�&H`R���Q�v�1�"O��"B�M:��q��Xɨ'"OBM��	�2a����$4����%"O���a�4�� ��H�2$8�"OR��3o_O\�\��'T<��݊%"O`����bjʰ�u�2��͊E"O�u�T)��s=<�P�]�S" K�"O: ZF���Z�4\&�,i�i�P"O��G���Ha�ER)8�`�4"O�} B͟��Y���F�
��"O��P�@ 9�e�R�]�k��j"O����+�U�z�z��W6*(%�"O�9$F*�E2�%������"O�a0p.F��@Q� `�"OLt��⎚3���CGL93:a3�"O�Ij���=O�tP�ЄO�!�Ԡ�"OЎ�Pwޕ�&�Gj�i�"OMi0X�JCx[ӣ��5a��B�"O$i�ȋ�:��1�Q:x\�u3�"Op���ޡ������W� ��"O=�A�Yd��&M[ 7Ll؃�"OR�s%�hَ8c��ga�]l0D�y`㚬B�.1�(ȡ�¬;5!�F�?��S#R--L�p�����* !�D�)u�Q'ʑ0=v)��S% �!���4x��:�.H�&U��ȁ,L�!�d�%���cC�E
��L!�!�DQ�{ (�@R���#Zvlr��	$!�ēx
�D��Bܠ�F#n�!�$J ��Z�F�~���ڳ!3�!��/R|����z�:u���	�!�$�16�θ9+�"k��9"���?s{!��ۗu+�� "W2h�t9��J��(�!���EϚx0�E(�Ѕ	Q����!��F�PZ��@�ȐT���ņ�#E�!��S4Ђh8�L�W&��s#ֽt�!�dL�8�xQ�Q��NJ�A(2LM��!�DF�.

QId�\�-��A`��/�!��;*��aI�N[	�b�㫀�r!�� n����
/]Z浠�,�$Y�V��"O�����M����H���<n�<h[�"O����Ȅ'#�~)���S�~�hK�"O�A��*լ\�h�!6/О~�5��"O�P�K(i�Dy�L���Z]�"O�U+�!��?&�%zd�:i�,��#"OP���↛r0�A�Â Qܬ��v"O��RGD^�O%��16�ǽ%�P�I"Ob$�`�y��k����<��""O"$��HR	@e�UN��a�" �6"OX�p�ǅ7hz��UR膬�"Ox�)��J�c�U!��
0���sQ"O|=J�Y�a>��箓M�Ԡ�"O�-[��E%k�v0�`&H���:E"O48怘u��U e�ڵc�А�D"ONd�')�qS �6�6��"O��u兯V�p1��TSIJ]��"OP�V���6�����4)�J2"O�H��!�.iX`�9�� \5(Q#"OL�f��gZd��`��D�	�"OQ�B�Vi�B�AnG�i,`g"O`@is��m��h���1Y|	�w"O�)�S�;N���2Ķ/�c�"O"t�,R�0��5��-��"O8��$���h@Y�����لT��"O�a���	h�>i��j�V�3�"Ot��W�
@�)�B�DYڷ"O�1c��q��źg�F�^x��p"O~�A6+ƞG9p�A��r�s�"O�m� fV6Etv��d-��� �c"O��@vc��e��D(��]X^�"OL��׬�4f��E���6�� "O��S�	&7��D5ʙ�X��|:C"Opy�Di�z�!"�H\3s��\9�"O�����6�����V�;p�]�s"O^���Q26I4$3� ��Gft�K�"O�P%dv٪���.� q0��"O��)A�|�	s��>*T�)U"O��X �z���c��D�)���Q"OH�� �\�o������ւE��B�"O|��s�IqL����j6�qh�"O�ӡ��Y�(�k��]Q��!{�"O��r�'�n)�h(�'�~x0i4"Oʜ��#ʷI0�����56�L�y�"OPq��M�[��ʔÐ�*kb�*�"O"���'31���Ǣ����"OJs�NK��^��C��9+}����"O�� �É�H� *w	O�6֒e��"ONp3d�)+�$�9�h�Z2� �"O%�@��������1pq�a"O ͡�*̹AZ���>*แ"O�4���z��}h��%���V"O��KH̳"�t|�D���y�F�#�"OP�;�`�yb�\����,>��U�a"OИ	�a/����
�#�|��"Oڥ*f�X0|�|��"M'9nq�@"O������ECjG�k��) �"O\#�A�������~%> "O�,���W�2����q�Ң$0!�&"O��j��:
���%A֞z	���"O��P" �6uI&@C"�Xi"O�M����G��9�r���@.Ec�"OP����Zu1V!ҧ�O�loz��"O�0$b*������B}��"O� 5��͊�l�舻r�K�Jl�XY�"O�$y�M�=B�Ud�Ej���W"Ol��◙z���
�±S�J���"O�5��I���u*�� �f�ejU"O̝���j���-�5"3�"O �Z�CW�HM��� ��0��"u"O�Ѹr�6C����1�Z�@w�I��"O����抂|G�2���dl
`Sc"Ox�P ��.؄T3  ]��0�"O��k�B�<�� �u�� ��  0"OZ�I�"[�*H�3�a�qo�h�"O���tcǌlB����0���3"Oΐ�2�	F�ޭrV��
%��K�"O<�VS$(�Zun��m��h
'"OD�*�E�*W��YrN��w�-K"O�pKw,&��ʲKK-wđ��"O�t��AQS5|YJ�=N���V"O�!�"!ͦ$�=��
�("b\�"Or ���>{�4��ל?F�p�5"O��3W%�]�Ț�)��.W��ҵ"O�x����=�.����7:�)@�"O���EM�M��CW�v����"O�hxsfW;%��3p#�<{�"��B"O=Y6`��0���;U���V���҆"Oi&�H��ƎėmP�['"O�� ��Q���@1��1oY�(��"OpQ���(i.x�����/6��"O.�jQ�Ȃ;���㇚wN�["O(�7�J�R¯
`��G��yr-\g��C�l\��<	��yR�r��$���0Ϟ@@Ǝ�
�yB/٘VЙ��ϟ�zT��Fe�y�X'	Yʼ�Ո�&~KP9��œ!�yb��;�i(DM��"G|�`�F���y�_a��uZ�"� ���,о�y��-$�|���ܘ)D���D���y����f�����=RR��
1���:�!��[�T{�,1⍂�=N�C&n�8!��]5WDEْ㕉,���,���!�D�"銁�s$ ,@֬�+j�!���Mk�Tj�MZ�QyT��7�!��=Nؽ��� mגIb6��;�!��7}��0sMQ�g�D�M�,zx!��04Q�<�դ�bA�l�cfO�hd!��\W?�8�œ�\�b,�Kť,!�7e�|}K+��\>J�s!�F�n��Q�b�Z;P& JPi�-�!�R%]�d�����:�!#T*}�!�(�x(� ��/1��9V�1'	!�D��<���lV�K'�(`#G�"!�dE�-�B��� �ftdr��).�!���#3ۘike�� �  8 ��V�!�$DrSFR�$ʴ��e���`�!�fa"�W�g�� �
ۓ*���"O����[��$����(X"l,CF"O\(�l��~d�}�cO�n�@�	�"O��`��9n�D�G�˯�-�b"O�L���c�d�� ���1�r"OQ�mI, P��d��e�T�b"O:��v��5��t�Ff�J�P�"�"O>�W�S���\����7^�8X�"Op1���u��R/-Z|H�Bq"O(%p�̌�;mf]۠�CyP�zC"O��J���P�Ҭ^���"O� ����G\C���:�hM2%�hIf"O�Dc��wuN�9a��i~6�B#"O����Gƫ:��Y���W�8�|��"O�e�HɆ{!8� �CW5q�(xc"O�=�w�ټK��i�1E�a[b��"O$|�Gd�< q|�y�ҐGNzp��"O4��NS�r��C�Qd*,�"O��%kH�j ÂǫRFN-��'� A���s��0qQ�"]r�'*��t��`� ��3�4��'B6�Yf���XI*@��	�����'��p���	yB��E�<{����'N^��J��i��z�LA-*�"b�'%� E'3Q�p�ʃ�S�9D��' j���/��U-:!{ӤB�^,b�8
�'�D�$L�--��]A#+I'WgV��	�'����֎L:lV�����5����'��d�G�5cGd�cD��7��<��'�v8Z����-�~!��@�T��8�'���3�Д<v��SͅH�}��'̘�0��@���2#��Dz�;�'wD�h�*�%�rȣG�הOvQB
�'���Շ��e�vxR��=GV��
�'��B$/]���8�*��K�H	�'~9�h��9���F@>�i�'�b��`��)H؍(�	����!a�'.��z��~a��MV\t�zp�V��y���Ec��X���^㢘y����yO�$m�`�5$ȈPs��2�݇�y����y �r@��EU!	[��y�#�7I�(y�$�P.����l��y�.�	Qci#�_8v�Z���X,�y�%�*$�2a*��[�o�e�%@��yBă�\�>�Z��KdW�a�0���y��V,�8m��@��)XySQ�Q�yBL�8w�R�҂gڦNPZ����ͣ�yb@Ϫw�RD�RT����]��y�Qin�(�d!��ZMzH��O�yr�X�Z�	��ԢP׺�Ȥf�yr�_=&4|� E,GK��m�D�y2��!
(9EN%�4���!F��yb�<m��DzB��%w_b<��F��y2�Y&)�r�S�v\�1j� �y��Y	��)�@��6���Y�f���xB��=y!y񦙌`R�!�!hG����)�<��4��ꟳ52�%���6?�4�@�'6�b��Z�d���`ǜ5���	�'bF�!�Q(1�fF֑zH0���'���`*P�h���ŭ��� �'¼�1C^� �@`o�:||�ͺ�'kLYae�	�
���J'!�v|�	�'��5�X�H�q���8f,��	�'d0ar�;d���Ĩ ,���'��� �48���[���({4�'���ժ�W�b�S��5x�\y�'�^-�'BJ�7��9VI���,5��'�dk��8-�x�b`� �>;�E��'qh��܇E�q�P��>6rn�
�'Cd4��Q�̠���е+�XH0�'�T�)�:��$��Μ4xٻ
�'����Bƣ?Y��xg���<x���'��h5B�4'�s6
]�}��M
�'x���,�.��b��hg���';,�*e�N?~��	����=
@"��	��� X�@ס\p��E��-4	Ҽ��"OXyq'
�r\��j���k���E"OP�`"��'ۘHb5��,�(�"OtYIFǉ�
���y�(��!�"O`���E�k��|	�'�7c�,��c"OP��3BI
5���F�#K��$��"O"I2 \#1�!�.�(��Đ'"OR�c'�K*�A	w��C�N��OR�겨M, ���{uj�e�O"B�	�22z�;���1K�l=K&�؁"Z�C��">hP"(
 .��1�qlVތC�	27pU;2�N.���6��	�JB�I�DѲ�кbA��D�QP�lB䉘پ��Q�ڨ;�`�Do�&!o.B�ɥ>I�Hc�f�2Ӏ��QE �+��C䉔B��%(�/�d*�@?$B䉌O��0d�
�Z�ᠠ��@�ZB�ɬ%`���%C-sM�,��C�:B��9|�����V����22]1MA�B�		3�R�O8�S��V��C�	F�|)��O�2v��h�A�*r}nC�I�����:S�\�hL-MLC��#�na�d�̀���G�}9|C䉥H��9%*@�'���9r�ħ cC��!ج�֨�3r��VjÚo�B�I�s&��Db�=g�	��AU S�"B䉬3"���2/��#"��qM�	F��B��=)��9r5�	�p�j�
bC�	?/��*割=��9!g�J��&C�I��"i"ׂjmz�Sփ�<"�B�I�(����v��4p0x��爌zټB�	�D��-�d�֞	�X��W��P�B�;S�YIVo�!�8�q���3lB�I85�劅ˇ�a�L�Ƀ+�%�<B�I�)9P��刈�r�H����%*B��%Vh3��1d]���5�JC�	*R���:���I���r���:|lb��ȓk{vً����
@�V��3�X���s������-'h	���V�|X�ȓFɈ �gdJ�d�>2���J�	�ȓC�BȺ�e�,%,�M
g�7#�(���8(A�΅p��ʔ�6jCt���E�*98����; L��钱��؆�J��ek�P�4��0{ІP.}�D9�	Wy��'>ў�O��5�򃘖j��%� !�}��'�0u(��*Yx�爄�9
�'�=P���#&�d�p���# ~Q�	�'�00���r��4咻%sh�p	�'U���B5�m�w(���l��'k�h�烞��dd�X��c�'d� A�W$k��ː+�G�Ե��'XtS�eO7f���W�T�8-4ur�'.�4����D�HAj�-3f�M�'��K��:s��(��9]��'�PI��$%��D��k�?�A��'BH��u��/y6���O��k�'0�+GF�j��(q$f��~N��'xh�{��]�X9'G]rc(�
�'(�|j� �'�41P�q�>a�
�'s��+�����*Vg�ڰS	�'J��0ƥ՚@�,@8P/��^���'�~]S�h�M-fu��çc;,-��'���K�ϝa���	�*'p�'�!�0c�q����s�Ҥ���� ���a׌i�,�)�E@�Z��"Ot����'W���c�J# �� �""OJA��Ƙ�~�`��f�� �dU"`"O�UwDԼy�FĘ0���"O�X���[���j�Ì�v��u*V"O�h0&��<�x���C�m�~��#"O�	� �� ���
�*�=G�ZxP�"O(�G��EP�A��ۺ�fi"�"O���Qɛ̘]���E G�l+�|bV�0�:��y�mU?��9����/7�$�����yBiևUd���4מ�Q�D��y��ВwG$L#�%�)�]��%���y��=�x�!��7aȀv �6�y�o�$Bnʈ����m|�cm���y�G��-�w���]������W2�y�E�r:��ӵ��X�(9�"���yb���]���R錮L+���@���y�
ǋF�ܙ�֬�:Ez����mX�yR�i$J���)Ui8H��]��yr��8	Ƭ��G�u��t��/�y�lϠ|�l�i�&8f��5L���y��
ug"lFm�kx�(d�_ �y2�9	��x�#H]�ϴ����U��yb����J�I��%C9$���$�	�y�!v)�Ȋ,rKĜɖă,K����^�#!NZ2Q�BT��M�$W~ć�-"��&�]��T��u"Ѐd��لȓ��}����A"2B h߄-��d�X��d�3=�>4R�NڻOzx��3p5�0ʮ+{���[9+��ȓt{N�c5 *d��I�V.=����4�V�[�W�=�(zUb�'p�L�ȓ)M$�
C�U�\(�af� RQ�]��B͜�:�h߀I���>���ȓ+3Z��wa�*A��|����L�܆�¾�BӅٺ]��q�OV�a�8�ȓ{�l�9�HY<@S�
�8��ȓ7�n��`��;C�ꀸpJ�{�ȓ2�ĭ�ٳHa��f⃳;l���ȓ!�aU@� .ֈk%	�kV��ȓ_B|2���I�u������ȓ6p�DI��j���]�Y�ȓBJĈ�#��:UP8��A���=�ȓ`��i#�=J\
�2,��7N"�ȓ7�v���rj: ��� ��|������/M08�������T��%��L%b��4���x(�ȓY�ʤdR�X��6��i���ȓ}����ðJojI�vg@�L�m�ȓ
%���AĝqZ$��lU�B�d �ȓ[���*u�T�.C(q�޻?ZR9�ȓX��XP!�5BKz��"ϔ"X��ȓ]��IC�
��E����"UР��ȓa0�5�E
�D`����c�#�>��ȓ	��kTfI&/���7IM��B͆�$H��0�g�7(3ܥ���Z�&�V��cl�!�M�_ڌ�"_�O	��O.���&�˶%�e��a�=ځ��Ӗ���M�>v�`c�$֖l���ȓY��q����4QHL�h���`��x��)x��7� ?�dMP'O�5%XȄ��V )-�飂.\�N�LL�ȓ >�0A�>۸�S�E�4sI��t00	e(B�6��dS3�t�l���S�? ���6��� �^�A$�J`� ` "O���@� � ��5��9C>�
b"O�� ��YŞ�j���85ZUK�"O��tVrײ�wJʻ����"O$�`�@n�@u*��/%)`��"Or���:)���@����g
x�§"OA�d�r�8+& э=�29�5"O����1Zj�!ڧ�"��� A"O�IB��V��+[1Z`r�"O�;qhS�|S����G¦Yc� ��"O�u��#�Zje��:V��t"O��D� �̵�ghγ["�[�"O�!��e?BD8�9�&� �� "O���UEh��ӑ��r��x"O���O	-OGzȃ4k]�.�5ke"O�q#�,QIg��ެ�"O�lj�@�j��\�1	��W����e"Od�B���7TF���Ȅ�V�&ђ"O��a�Erf#"�o�B�J"O�=�ނ^׎MB�.��z���J "O �0�R#r�e�'Ίz�,��"OA;u�93�H��dc�!�bY��"O�y�B��Ca�X:4#��n;�j�"O:�r��M���T�X:'8*�R�"O|8��L1�h��t�	@P��� "O~������g;�h�<b0d�Q"O���NE�9FX8�������"O*lpc� ��Ч�PY����u"Oh�"�Q ('$�)�~� Q"O:}����H���g���H �A�D"O�0��΀,J9�e��A@�_�Bи�"O
�B��1ڼ�a&`/� �"O������8,<)��8x��	�"Oبb�N�$O~��b�˞iܱH�"OF���D�J;�J���"e���"O���IYJ�`TL��Z	�"O%s�Cm$��#z��F"OV�irǌ�	�>8c�b�lq�3"O�������W	�%��f"�Q�"OY ���=(��l(V��=a��"O(T��GH���А�5P�h�"Ob%�p�\�[��D�7uh|�4"O&8�lҭ7��pC��2?�d(�"Od� �L�]�H"�J�*6])"O&�����%�� d�/xj��K�"O.lc��Z?#~�X�H�1Y��7"O0����JH���V��l@b�"�"OD�gN3md�0`��)�dB&"O	�U+�n��p�O7[.�)�"OV��c�)v[��"�
q�A�"O���DF
-G��ٰ���}��"O�@e�$ ¤�dńu�2�rV"O�"S(�u$���l�45��6"O\��4#&n�6;fa�Ȑ]�&"O(s!��Ԭy��I�4uW"$ �"O\� ��Q"d�|���XN�"Od+�j5?NU@-�*��"O����"P�db�,��CR&:�p�BE"OЭ*d"�v�C`C�*X�^�(@"OR���n�bt��G 
2�&�"O0��
p&�8�S��rD9��"OҦKl��azV�Ļx���"O��c��9D<w�G�|mK&"O@�	�͐u�,�BcN�T����"O� �� %�_�9[��A������"O�LG�6r�F���0��s�"O�,�R�ՠF��ĻT㚺��)��"O������tm��bq�оv ԑ`q"O�<8�,�9p��=���<&�Sq"O:�{�;*,���P.z-(<2"O���1G@���@J&ڱbN�p�"O ��ږe����G�P��a�"O���@4����l��{�"O� 	�$FV�qI�\%��"O` {5��)�l�x�(�T)��"O�k���,p���C��P�Y"O]#���sw*�#��20��U�W"O�8�W��vX̪%l(l�@h��"O^��fгh�$ @��}�*١"O.�����b��<�"��{�||i"O���/�r�|p�@O
�`)�"O��t �.�����g��f"O
��%v��2 ��v��˃"O� �'��y��/^d*��v"O2)eG�	N.��#�u���@"O8����G���beK�e
�XD"O�T�P�֔
�>�HA@�K�ЕI�"O��i,چ*X|-x`O��^�F1�"O�\���O��Q�.X'3o���"Omy!�D.DQ<!�F-۞v��i�"O�YY �݁��qR���+'��X1�"OHB�H�~V�.��1y&�1t"O؈AfÈ�#��X�Ȓ'Ef�Ј"O4����'q��t�Ӿ^�|���"O�Z����;�%�>��\C�"O ���-�H|d@2�Ğ0/�*s�"Oh�*@O=T0pm�V�ą+��[""O���1GR�5Xr�Hw/!<r�RP"O�<"�F2LS
 �d�� s�d9%"O��¨�8�r�r���*>P�r�"O����ȃk�T��`�aOHKw"O�X�uCސm������V#EEt-Pe"O���$��j���B�í~A�"Orq�4ě2�BС!�ύ&���"O�8�6O+\4�q��Y%zRq"O�ͱQ�Ȫf�f��F"O��
���j`��ޙh(!�"OD��bڥuL���$�jԪ0�V"OXD����3Z�|����&l ��q"O&�i�fY�yօBơC:B]4�A�"O�	���$eU�� a�"SO�ш�"O�y����i�@Z�2>isr"OA�u��� `��pb
�t�u�1"O�HF ]�XRp��G�3g���q"Obw�?6��2�ɔS���:"O���@̋��ZTe�y�0t"Od#�j
(��}چ	��"^���"O�i"��C ��.!T�Q�V"O���,�5��5��g�nS��8�"O�1�7�\3o�j�#�{\ΌQ�"O �"G���A���^�MiH��"OTxB�j5d{��;���+28�Q�"Of�K��ĭ0ר�t�I)8��]�"O�<��(04䉧J�!���h0"O���%F�+����(�+�8�K"Of��o��} �����Q�)��lр"O�L���E�)E�${�Z4&z�]��"O��s��L*\{��d�=I:1D"O� )��D�([xB�J�ߜK�Ԛe"O����c ��1�X%&���3"O��K���s�`���*�9'��y�u"OQ�6��E��m �X.�&M�"OVm�$�½ 8Z�R��)�����"ON0���#m�L4��nͶ��T"O�UA���xI8��PMc"O�ڠE7,�B��F>$�l��"O��Hq�P�=^���W���@X"OءҧH=<~<��o �`�"O���,�Bx0a�#��Vغ�Rg"Oqp��ߒ��da�D��9���"O��`(@<�:I��c�#M��ip�"O�S4nUp���*e#
�2�޽"@"O�Ct�ӟ/(
�ǂ(�� s�"Ot��� �sM����Ůzx�� �"Ox���<�*�X��[D��)6"OL�c�*5~�Ps.�)PX�x�q"O����t���P$.N?(a��"O�5�bC^�.K��g�
 v 8��"O
 Xao�f)H[�W1bo2-#"O %C��)	�A
�F�^Y� �!"O� 8�ԯb�Nl����/K��"O�u�&��j�v}�Rd� Y>��"O,��如?�U"��M%26�!.�!��o���F	In�ӷX�^�!���f�JhTl�;y\��@�cF�[�!��)�j2$Է@-h�ف圷H�!���>�0a�,�@�C��!�$Q���bJ�-��jv	\�!�����p#a��qR�}�"�n�!�$@�~u��Ã(Ge�`�Q�X�j�!�֮â��v%Y,T�F�ʕ�Z-5!�$�  �f��(�L�c��V�+w!��&�$9P�%Ė~Ȳ�	���"i!�D<�r�A�L�(�2�{�Px!�$�&{J��q��7���ǌ��Ri!�D�.\f�詄�Ȭ{�~�Kw�ނ@g!��9DT��z�fܛzS.ԚjU��!�����1R�bmr����[-#S!�$U!6���k��u��iS�FZ�?!��Bb26�P�!#8Z ��+�OB!򤟯gˊ|[���"nˎ�` J�>^!�䍁Mw��E,˴`�^���jX�f!��&?[�m�棙;�Z�� �^?+D!��4l��9�vK���	[�i�W5!��4J����ڕ)tfM��
M)!�d�?,W2�#G	�^�0�7,ъ5!��C5}�́�,�F,����%c�!��#����ʾ44�0��N�k!��`f^iprŜ- +.t[��C$V2!�d���赻/G�-2�t�$�ҳ[!�$�4�>�Qu�:�"�3ۚi!�d�9\��#��%��q@�hS�V�!�E�j&tU ��]4 ����'�/|�!�D5~ >�A&�B�F���I�g�S�!�dUl�,!�SA@�C���r���*�!�D؀J ���g���|#"!ku���!�dU&et<��k�E� ��&K�D�!��!j:�	�DV�h��
T�4�!�	�T=���X(4�C�*[�mw!�d܎�R5�5�	�'�(�&�#is!��Ph2�Jr���4ܘ��D3wY!�$ЫCIl[�&A������X �!�� �Ⱥ&����=`�!ĭG��"O�鐶D2!z�1�N^!(�""Oҡq�gƍ.2�!�U��4@��"Od���DH�����䓗h���"OfM�d+�%&e<H���hfI�'"O�ݚR�ӦWtiR���.I�B��"OU�G�dufm1 k�-3�`E��"O4�a��^.n�9�d]+_�<+�"Od���i�+6���CRā�E�0�{�"O�L�f�3�8�T%�"SP���"O`���*��H؃nOAGTh�e"O.1�q�?�:ԛDUc���"O�3scd�LD����F��[`"ON�1�A1� 
���;~��=;�"Ov`I��ͫ-�P��=!yZE�"Ox@�3H��%ɴ��%oȻrl�`�"ODt�l��}�ЀP�3dN����"O�0� ��\���� �� S"O�0R�k	-	��-Q1(�.�b"OZ骅(�V�� �B+��R-�|B�"O���(W�A��D�&B�f�A�D�P�<��MC]3���b#%o༈��%�J�<Ae��mu�Q��ƛ]���UG�<	6�ùp �PB�!=�Bm2$A�<��AZ՜�Jf�P�1I�!Я�e�<���XIz��D�k�,iu��^�<���4dZ=1���M�T�� e�E�<��P`�ܱI�d�5;�FDIj�<Qr�T�7�~u��g�4�,�j��Uf�<�t��#7Q��FL�W�1�Ėj�<����88�+[b���.��o��B�I!)����Ld�}�k�Qn�C��N#�pRcE�APHH@0!َ�vC�ɭw�*Urƃێ-�]�$���3�XC�I(&:13Ed��nh�ԉt�"C�I`J氐�H�]f(��@+nQ�B��4y*���b�c�><c��U�= �B�	6pd��e�G jv�y�>C䉐"K`�SѨH�1]@Q��ڮDTB��Fn̹�R@O8+��bC���hC�	�=r]
�O�4A��8�NĒ7�ZC�2�%����L,���O� <DC��	Df�����;et�`h�Z�a�ZB�	�G�a�7f��v���bG�0fHVB�I�C�F�{À��!P��E��
PTB��*w��@�w��M,8I��bs"B�ɶQ8dX��C�$����/�7��B�,�L<hP��1t�`ҋ��&��C�əh�HR�(��b?f$�Tj�
y�6B�	�jR��$A�%�$|��>y<�C�I�q�d���۲oj 0B1B8GAB䉜>A���i8A�0���]�7�C�	1( ,�5��2q7�q3b�ڋq��C�i�fQi��-.��e�D�	}ԾC�IS�>��iO�;��:�ꕖk�PB�ɕFg�HHrȖO���So�7Z�6B��&� ��O�L��'��+��C�.��0��E��#�(�ڒU�8tC�I'Av�s.w�Q:�6 �8C�	� l�[�۴K��`j���nB�	�))�J`��P5~�2a�ďw�BB�I�-�\���	��*��1�G�;�B�� mM�U:�g�H��Px���3�B�Iw\fDs�!8v|��0C& 7D�� hM�a��8�yY1�եU�t"O =�E�>Dښ����0�4�q"OL�c-@��`XuH�(�؍��'�,�Y!f�6�:Pq��5�>��'��(yWO���2���N�l`�'���G����0�U�vĨ8��'��q���JRe��iU������'#����'B��;���ƒm{�O�!b���]f1�'�  �7�]�&����-�s'W�d�xX�n�,N��I��H�P(����y�2h����00ę��K���rɀ�n�*5�W��1W���ȓN]Vp�	�aYrt��F�`��T��� ��-K�u�D(�cR�&pF��ȓGYddZc�b�ĩ����,�hQ�ȓ[|Е+6���q��1�* 'b �ȓN��l�fF��Nt� oF
�$��]����eF�Hm��W����,��IC�'��pR�n��� r ���p<�a�'j(\�U�V]�Ȝ�d��i���ϓ�O��Z�C]�0�|�j��ԠR��a�"OB����j8u�QL�#Қ(C��!|O��U��� �vt��n��'���9��Ix��+��I!0D�����;�F1�g�*D�t"a�[�6�����	ȮD�Z P��6�O���Dh�N�"�~�����],���Iw�'��1��vO<��������-1D��#��7!�}��ZP��J!)3D�dJ��W�-7zeQ(ԪN�ڀ*p�5��b}���t�x�4�p
V`�{VV�ڑ�z�jC�ɋE�`��P�a�:�R���?8B�F���OR~�~#�PeӃAt�i�
�t��-�ȓj��Sa��Q�\�qT��X���'Ma~��Hq2$�Pc��;/U�|�WBW��>�O��uȂi�%��W���"O$�ˇ�T�IO ��4զҚAb�>���?�'.Q3�HZ
g�(B
=}�f��6Op�'��zBC�R��9���2�X@��Ķĸ'4,<R�5��$�'g���bR78Vy��k�L!�	0�<�%9���f*#��If�O���]��� ��SG2N%�0�i8�`��	�*����, �ض��$T�dDC䉞q��[������&���O`�Ɋ{"�4���:!O�06�����at�B� x�c�n�.����l˷�B�I2L�Xe1��m	���%��lB�ɷu6��P1m3N9L���L<zF�ćW��uW�I5N�P�be,�(Eap �2��A���D�\�<ܤ��b����p��� [�@!��_���S�H<*f��gHBut�eF~��ӜҠyg��T�I�#c�-5y��H���<�pG�!&T�#�)cŶ��eNu�<9�j!���s�Ȋ)N6u�B^q�<�6/�$Hٲ �2 �"W����B@�k�<�`�QpPd��lJ�b<��j�e�<��O��\�6Xp��C�LdJ0#�U�<��kV+qy�x��h5���9c�}�<3l�8E��i9�_-x��q��w�<����c��Da���"���#rev�<1��
�My0���hI���n�<���;"
�gI	rLd�`^s���hO�'N�8aA�`�(k�p�
� �y����ȓ"v��Gfԯe�z��)�"%�Υ��W$��e��q��pC�֞x��o� C���iy2�8��� f(QO��|�PXٶa�+x��!q"O��2qI8T˲l@p@RR�V!k�"O�0����h� |Y6�I9]�] s"OX��!A��d,�r$ǑW&���ɿ�hO�I�=��e��!�-L.���V"C�w�!��%3QAB�-�LothY�#�T�!��e��x�鄽C�eB��D�:�!�D����g�(c������8�!�d�n��xɃEV�\� ��ňX�	ޟ���$/ʓ ��A��A��b�H�h�"1A<z��ȓZ��AK���)l���D`��~�Dx��):t -i�x�3ƚ�%���i��L�<�.�*(H�9�vmQ�<���e��F�<�� �:U�u�g�>,���w��l�'2�?��� \�8X��4�[�����ko������4P��b�N�8���I�	����B䉭b�l\󋓒Vz��+gO��P��B�ɲk%D-3q�R�q'���c
�'��l}r�x�P�$���1g��"!�������#��/z�C�/%� ���Sl�-/G;����O���%i� ��7�,�k�,l�џXE��HɹI���[&�^°m�f���y��C�9njhd�Pʶ���ɮ��DG��/}��I� raY����t��Vu�!�C�FTxTS��G�)�0�� �C^���E{ʟ����~��i���$K<)c"O�|"&��-�6�#�.'gԀ�[��G{��I ��A!5�U<8���פG "�!�kE� �'"����Ph��*��*<O�tiv�U�m�!�h0R�'Y��	�<I�����>�����=N��B�I�w�0)H�O(1�
����1(��61}���UyJ|�<i�=	��D�v�W��l�<�����c.�	�dǄ;7�>�pu@�jy��)�'x6�!5��1KB���	 �K/^\�ȓ?n�Av�'ZԠ{�WQDn0������`�H��^ژ��ʙ
�HOO�,A����C{r����ID[cb-�ſ�y'Ҭ.�b����O"�<�:i�,��=i�{��N������8�C��y��)j�xqg��(	��XM�y"��D�lA�����S^�p���R�y�g�?h��p�(�W�4�"W��ē�p>��P�D*�	� ǩcM�A3�.�O�<Y4L�3R��9�@��+�=+$��N�<!��]|w`P��c��23dK�̦m�	Y�S��M#�þ>���s���_���r2^H�<a#͙(h
�����h"ڜ
b��F�<9aJ�$�vh�D�;:V��Q�ȎN��$�d��%έ<Β	�A�F�AL�څ
%?�Q�*�O�;�a�;L�`bF�&M>�R�>Y
�l��A`&�:s�U�w#ݐS�=�ȓF�x֊�ce�U����=�<�&���'kɧ�O�8�E/̓rtp"�a��@��	�'�Խ�"b�V�+k�J���2	�'�Ja�q&@�>|x!RAD�Bh���D9O�Pj�� @L�g%�9Lp�tӱl&4�4��HքZ@~!)��M�W���pP%"D�h��*� )���cPG �H��s�$����/U�-H"Ӝj��%�����e��#?��O6c?qc"䅅r����\�)焤!�/D��c.{�4�@IV�qVx#�-D��e��*"䭒Gi.,nTy"�0��G�'�IgV���c�9&%*q���}��B�)� � S�Å�9"Hy@4ŀm#�Qˆ�kx�H+'��n�L(��/_8��3D�`�#F�l�,	�W%��Մ2D����WlĉC��;-Nĥr�
/D��X͚ܬ����'?�h 2�)D��	�	0H�p*e��.hf�x�&)D��c�!W��d(#kQ�$�n��1
<D�����(��䳄��|�N�iP�;D�Dy�J�0�@�ѧ�P 2���+D�p醇D��0�Z��!���.(D��`���RbB��!k]4�x��'D�̠��KN���&� {DBw D�$��٠fFu+��PD�C�=D�9%k�J�Aa�P!J24�Jq�=D���FH?u�"�8����N��T�`�:D�$:f��2�v�ciI�j>��3�9D�ܚšL{$���i;&���sp�7D�|���ڠfH��b�X���i�fJ7D�t+#�ؐAu�؀��T���RJ6D�4�p���KW�<G��5:D��b�h_"~�v�A.T�����Ǥ-D�d����� �B�*�Q�w��R�,D��;$A�/W�	A�h�'Ȫd���+D�����  � Aaj�3�Bm[��+D���Q�U7-Y8f)L�QAű�I&D�0�D�e�<�r$��9\@lB�$D� �q� [r� ��*l+�$5D��(��
wFfE��	��.8<A#5D����H�7�5b3��<�,����5D��"Q`T@.��)�MK�}r"e D����)O�l8��ሠa�b��c�*D��DAG�贌�F�w7���((D�,s�:j�&��^ZL4�4�"D��dO�0x����ĀC�<��L�!?D�xK�k� ��mǥ$��Ĩ��?D����m&AϞQ�t�5~�P�i?D��{�샡e;0�J#F�D��\��7D��9�ZMy^�:�FB����16D�+c�R'9�J�����L�6�9��2D��#� ��E�_�u��qc$@��0?I�@�n�,``�(�@,� �.E\	��]�<���V?(�0P�&ű7kX�C�L�<���?��!��K$P�V�҃!@N�<ن�N��8mzd̠a��x�R�FS�<�Ѣ Z?<�	i�H�@�y�O�<���˛q}���-�:^��c��I�<	��
p����D�)~4�]�+�D�< m�P>, �I�+����v��Z�<i�k�3:	sԍ�o��ʵ(P]�<��iU
<
x�""��@`�8�&�\�<aW�̝��������H�e�<ф����zQ��T�!���Cc�<��B� �P�0�������X�<�V*҄ 5���p H�^=&�J@��y�iT&e��Ă3$	�;�<�"�y��լZ� �uJЕ=���D�,�y��կg�Mq��(%����#O��y��]y8$��u��KS�+@�T+�y�M�p�}�����9�N�9�y����j��5hϐd0:�� �y⁧"(.�Ff�){�٪ӉQ�y2!O�21�Έ[�j���a��~��� wD��2E�|���C% z�uH2�<�\���H;!��Ԣ��y��
�`$��6��	)n��8�O�U0���)� �(qsiH64�� ����8ڮ���'p�Q�EK��'k$��R���@�0A\U�m�g;+6hń�	��R-���"������`d��<fF�\1�rF�? ���O|
A@�."x�jT��>�iZ��A{�<����oܐDJ�r(<jBn-}���ȶH� �M!QG�"'����'W����cՅa�*�qd2Q����'�F�d�>@��2o.��=K�*Ğ!@��sD�*�2��"�2�����V�-���˂�]�]��噼,Q� ��B]�[��D�8Y��B��&2Xp5N�f��Pd�\@���5i�S����	��{�V��S�����p�8�����8.-���֛��֠�ځR�C�b0��q�ZY�tƗ64�X��F�U�\���.D�iD!��/0;��1J|ҩ�L�� ���*�#8�&<�D\9h���\?��AX�<��as�@?�2+ǃiA|}ဎ�[�T���sܓZ�v�֭9�S*\źmS���UX H��]���"Q�EU�i
��ʟ>-8ґDK�,� ���� u��&���@p�wA��~�~�ڥ�;j�^1yI>ɕ+��i�N9��6yp��+-Y�L��֏T�
]B�a�H�;�bY(���4"��\�P儜G��O����Hх:r�ժp�1��F�꫃o[."p�a@E?N2����>�-��֞P�ᣄ���V��#/Ҫ��AU�;	|�)�دF�)��D�_�^X�`�x%�Ǭټ&|����:��P����1��=&�ִ ���%hT��ɇMB�v��L�r��)�x�44a1h�?#�ƨ �쉥hRt��A��<K�瘓G�F ـ���p�����<����Ȅ;���S"��%$�8��PU����n��&�� s�i�0a\a��O�@�B�K˳$��;���W����nD/%���I�bH)uA�6V� �`��I:L�fl�B#��A3���D���'bPTX��U�
1 �"Y��X4�E�t�F��*	?cr �w�ը.4��ml�����G�y�T����� /��ʉ=j`鷈T**8���u��OY}��*�jDvt��E�!.�툅'�7����$F;]�n����Իe������y�"٢\�&����A. ���Q�N�W(�7m]�;1$�����.�݁��|� ǆ���dB��08�X��rHƱ��J����� L_�F����p���hq�i��^C�瓋p���xQȉ��ذ�v@�	!ch�#42Dй�Eǘ'P���{�
�s�f;���XS�K�r�PS2�9��$��,�,���YԮ�-�ص@�Y0�#q�r~����G1�$p{��b�Xƍ��S��j]	��]�*q�M�D�ݺ}q� p3/I�IH�;�Hnʱ�'�<)uOH�bW4�Iw��4��CJ~���5G����`瘿~be{��ƛO�fI3�hޟ
}�Ջp'�75
f�ɔ)�t}���<����s���G.�,)Ҽrg�Ƀ_F���×�|�h��"aL)r�� Х ˟"~��5b�-��2]"7" -����p!Z!B՜t8�j�q$���^��r�ȅ�$iJ�@�(��λ*�m�ь��cD��F��3�����g/���2V2����7扲W<��5,��Ƭ��f��e��`����� ���i������1�o@d�����1}�a��d=J���hBA�P^�T
S��\��P�0	�f�]��L��i���PUYE�Χ5�(1���͖
�DJ!臆DX��B��w�8PBĆ]�p|h���l�I�-#�Ѐ��[����}2a�^�>���� Y�a�Y�����a�B�IC�HX0 ���R�	_�&����Z�s�%�S/�#w����E �m=�p	�"�O 5bG�O0:_ ��N�"~
$���������*�>�qkH�G/@us��n7z�
0�S���0�'������(�(5���C?	0ŗ2&.�H�9;6��h�!�b��Ѷrth��}Zww`���CA��ꢤK8k�R#"��k����A��,B��۶�D3'*���v�ޟ�8�r$J{�'��pqlE�� �@&Eո\��b�{�*�.F|
-�_&���bނž�B7��EF��k0��]�>4�B
����=CGjM)u'����N�#�p?�VJߖ1x\E��� �� ���h��MY�T<
<� KI#&5P���4)i�Ҳ'��v	4	�y��=G�8���W�t q�m��yB�̐1��\BCl+r1�X��@���0a�I&5���2#�_DA��3��x�,N)v9�p��Ł$��ݵ#�����J�$jW���g#S��0=A�/@R��!��x�=I����\����@��H���C_S�I�I]�	����ո_6��	U�_��hOd,��@��� �Fe�6v�N��$�$\�t�^����!
t�I�� l^�A+gԪLhr� `ʪ6�h]��I("�~���F�P���:��J�����I�R�"p�A�8:�,�"_��{Պ���"�A�#G�����I<Q�6<�i@�,9zČ�"^��]	A^X��,F�g\3�n�TB䉭�.�A��	s�Lb�h�)^��zaN��2�N�0�/ S�n��%��-� ����u�X4Z���+[� �ٴU������ch�<[�/.'�>�P��p��2�FO3E���zB��
U����5}���l��~�@���ƳF��E��<)�XC��=h5{4�[8�$��8b�(��"�̓\�'�1XD�3� �!?��3oQE�} 㠁�
�����I�=��1����;��ɓOA�4���H����!�$%�|kRN ��N��8ғP���@��u��!w�jWx�rI
�H�Fȃ��@�`��`�F�)��x����La�hN�lUtl��	��Ї�@�.���m
�9���R��;.�)��\:K>1&N��+��@#[���K�k焙s��J�:�Ȝ���+KE8�b%)X�B�����iP����/V���)�I�{����Q�T+JF>�JEɘA����G�˝`D��ܴPr��0�
�	�"�*�dؐ!��H��Ϲ	ۺ��P*C�vN�A��ЏTu���
)�(����"��G�:h��P`ELڵ����Au���/�S̴AqH�C=a�'�	k��p �򄎇L,4h1a�<ouh��a�y�vD�4������G	�4��'�O*<DY�)?ixr����~�rt��g>�9��䞔6ղQp�B�w�lH�c�:N�Aa��ޔ4Ӣu %�
|�@&��@�? XA�2�҈����F4~�kuʕ(�<�8�O�	Xrt3��O"D�iE�CN��P�	�ȕze*�M��͐�KM���P���S���K<�p!O�@��8�`�!����Q˵yzޡ���B HU@��� ��B�6�*nZ 
G�ѣ���Td9p��E.�,���O?8<T8�)Ŗf��ߏ`v��ƀх�d���ң���Pц�9m iP/�4H'>¡,^�g|��V���@����"���h�f�u-F��0팩d��B"+\���g"չ�ذ�MQ�%��MKQ*,�q%�Eb�m_G!&���Nǡ�X�r")٦4���X�bÚ~��ɧc��X��B��
`���i�F1�Tlҙh��1C���#���P����L|�٣˓_D$��1N@����_is̴Y׌H�x4���t�@	(�)���vΈ���ϚKV�ؠA�"�l�`��+~:������8�I�j׏pĘ��e�����Y�êM���0Qǰ�$���q��e��IAA��T/5�Ї���VdH��ٗ��@� ND`�؛OK/9y�m�5JV�	�6��z��q�U��(�^���@����G�^�\w1Oh	a�E�B��q���5l3������bP�PK���ɊD�fΊ?fxQ�勷F��],CG�A��Ĝ5�����}Q�����K�6�yQ�8M�%��e\>����4�S��<�ǋ�$%	0��#/��5 ��B4�	�@��EB�@��9�0�zc��B��l�;�.��3/R�5$�
�A��Qr���hH^����	+h�!���5�0=�V���6X��HS�\#�F�a?P�%J��W�\:��Q�i� ��x�
�.�)~6P�3�@���-Sူ*P҃�ʄp�D�R��p��M��$�p�O/w��l���׆9o�Җ�	<�e��EI*|i���)jfHt�_U�T�@5c�af\|�@f�����'�nXCP�͉J܈�F�J>2�ƥ���dH{_�9�B+��U-xd�,����%_*��eja��WAd��Kк��
,v�ZIp� U�G��:B�"�9�Ahf�=0ꐓ"'�L*��1�X�d�1 ��#%���	�`.<,�v����C�b5ff�{D� ��:��S@�L�]�'D R^��K�(�3 ��o�N�F�J���9����Ni*H��/T-�p=��
Sa8��e ?8��`n��,��Dx�� {Ur$��	/�����M�<��%F >;��*0/��PP���"�y�#�S�(���7Kͦ8���R���>����$D:�E�?U�b��oN�h\I��ə� �\�#�)��o��ثV`�%;��i:�(E�P�t1�6�<iXE��i&�y��HL��@���/4�K��Ȑ�HO����B�$Df��U�@��	�\� P���U'�@��7���`�|��E��
Q��A�D�^�l����\�*#>�2��S:f=��m�-O���RL,2�|���,ڨ���쎒-Ȝ8�B#͗R8n)�RMK/J��<��H�/;�X�s��6}�~��B#C�{U�8)C�<�hM�wjG��>�e�L2T��X����)V4z�(BG
�Y���.�%?P�bU�� u���k�3P��d�p��)V:`�`�'K�e�9/&D��ԠNdp]�lm�p2�KR�d|e�Za
�Q@�N.İ�&:9�|̱�$ ��m����1ǧ�?��8��Á�4�x��M�uw�����ß��6O�#�8��3eN���*�G'_���@�-_A�]�!-y�p��:<�D����l
0՚Q��6]�<{�T>�D�F���^D��N��T�3���j.�=i�K��iaVAiU1�G٩g�E� |I4fЗVu��2vKQ��)��Gd }q%��`�m��� C�^�	�D��L�a�S )��(pN����>	Q&�)`�`%����_F�0OB�h�r��W��j���Ŕ� J����* !�.8��2� ���y7�U-e茓�cͼAHƨ����0>Q�E�B����4��1� �C�%�'�\���[{��!Sk@�EX�y����]������4�����"�@��
�
��I��Z3����W�\\܈C�әM���Ex�i_�7�t8q�,3�0���$6��a{�Fa�fE1nK0�R��D�3>Vy���7�tQ�/z@p����ruc����!OplãF�`D�i�0I2T����Ǵ8`0HY�$��[�e�ܣL|x��F�eI�]��OE�m�0�o>�XD��2e�a�R���X��}�(��ի�>���姝� ށ����Z�<�3�J�X�Uz�`�x�0��U����1�E���ҝ�;6���Be�8y�Z�U�̡%�����	�3����#f�bw�x0"E.�e@V)�vb�=Z�M�.J�ѰB_e���@Wf�!A[�l2@�&�M�	��ug��'�Hr�B� &u����@A�.=��RR�!�	�D)9��Ҫ�$�S�6�U����W4���@����S�����[!M�`XQ @�=��q�٘MŰ�*&� }zvČ�v#
L#�ϕ;a��$jd 'fD�j'� ��V�SvI̠C�\
���r)T�/U�b�����%cL�`�ᅒ�����%fԈ�&P(+7:����d�i�I:1捙m�˓8|�$�"�F�FN�aQ�ج6 Y�s��0-_r�
��!��A�=w����(DH�yaX�2u̻%��t"#)J�pv���5�J��0��'4��iv��(R��&	g�OI<=�4f�;��4����]�敢� �4n�!��
�"Lَ�I�.69a�&�=���$��2[���b �S?
�4�,!H�#D(\by��*-E�L�X3�OF�2�(��Q)x�I�����5�&@BU�"U,P��V�ytR���ឪG��J���8�n���g���*�M�+f�b�[A�6�ɷY�\���aǱ�duRȇ
k{"	�7�V�/b4�O��w�~��6G�x�t���O�n]��ƈh~.-��MW�)v�1��+���b��0n���	ˬl�򭉢+H/7qO�H�u�ɕ�F�!�\4L[da���FY��@-]o�;& �?r��%�2
�bX�%fQ>ej����ϹBQ�%��-Yg�v �:{�{�e�0\@�<�T� ').q�Q���X�ƨ�'>�p���dX�����]�!uI
 S
�0�8F՟r	����N�m[4��
B�'&+!��ՙ��6D�4���ԑzfD�z�\J�E�juT5��F�)%���m)s��f�W�:}�3e��7���g�mdf@Qu)S8]X)ɠ#�?m+CC
�L�$���
	Y\u��%�%�fqp�-S�:���7���_�H!��c�&�˃��}��YPe�!�li�<`�K%�
uCu��2C��qg��L@��5S��s��H�p2 ��ĈCU%��2B��2ac�	Q���B�^E�Poـ !�s�H�ؕ�	��́�H� 1O���p�	�+�L`��_z� �X,��	�Ԫ@)q�h8�&N�|^��R�3K��Zg���m�����/���$j�*w�Xh 掀|X���I�r�? �9��E'A����^���Q_�����Y��؂��U	x�Yc��Iv���L�|R�9����A�
dQx���G�){Jx���/xx��EƫyGdT�b��9����!
eRp��䇇*~Bt㱳it2�Y��פKʠ�����4������Ә�|Y�$L�-�\�#��ګ]v�S4^5��:����T��p�B|���a�-)V�2�Áky| �w�-L�""T�5
�6��}���=�Sc��Kn���ܰB��i�Ђ<\0d��.d�3�ٷ%��K1�B�jh��Rf�B��u�b޾Z>|��+a T T�R�n��`(���]I��F��F�"�ɖ�.�	�Iw�����)p-q�c�  1����R�\�Y�ߍ1T�B`bX l����şDS��C�- �%���oݙ+agP�z0�@He[>5�g��`��a3b��m� ���C3}rnD�ض2�A�&&��T�l0j�V�Э� ��I��[�M�A�D# �<BUĪw�dj�E5#@ �g �WsJ��Ag)�'�y׏F;~@�P7����0#3���<�j6�(��p �fmj���t�2��aٛweȕ�����uy����!G����h��{�au�b�0"�A:������U橚�!N7�V\J�E�g A��O��i�R�(�~� K?�I�S2�1���T��rs$çH>@a�6(�41(E�6D6t�ۓ����f98R	k��1z��\��)�Ό�C�1g:"�Ö�c�бg; ����U�S)b�֩	��S%���d��`�"?�.M���<ad燥��:.{JXk҂ʼdS�H���P]JB�ɋ�Z���LW(���(Ƹ ��ʓ3GX��,ʢ�ҧ(��|����9�l��―����"O�P!�++�n��G�T�+���9����H��yÓFhdx��#D�[��x�@�?b��ȓY<�a�C� ��A�# ��7��ȓO�B�ȶ�NR��z��?
����ȓ�4Xꀥ6, �`b�/Jb�,��3K��������`��,��s�8��]�Q��Z�+�&��g ܈"@��ȓ;�)yeE�(n� ���C �=��<{��!��s�|�P�i�1y����ȓ9�xa�@R �H��*��!��2�^���bQ)f(�ɷ�X&yX|���T�`��Я�|Q !Ѵ�"�4|�ȓz�nɰ�$&e�阁��!=╅ȓE���Q��̦,�T4��ƃ# ���z2�u	4�W]!�X �$Y�c����ȓ<�պ3������K�I^q�<��.����r	�3a�)ㅋ�|�f��,`x8��
 k����Q�v|�l��1��]��o��}S�Wi�<�(���6h��+�(M�gz������~�D���YF�4��)�.pkx :�
T`d�Ն�R�s �L�lǸ�r�W�-�����v���+v�C�4��L�`�;fT��
�XM3F,;hlm�'b�a)�8�ȓe�8�Ɛ
a����n̍{��-� ǎ~vM`aK >��-�ȓAQ ���,ainI90S A��(�ȓJ?�ѡ��/�������x�v	��<�Q�se$�2ԋ�$r���:V,�	�[�=��=���$T1�ȓk\�󖩖)N�xԣ0\� 1���l��f]Z-�q!&/�< ��ȅȓBm��At-K��~�pAŻ����ȓ[r��a�6M֨q-[8 �D��&Tz��&��o(z��WE�ai4�ȓ!��q)B��"�z�RR!L6}�ȓKVL ��B�lvL�u�\� ����76D�b
�y\d%��8���ȓ]nP�!�h��pR����*H ���ȓJ��"BgM��ֵk�Gj�Ćȓi��,�d剅k�򸋴 S�t�ȓ��x�p�J.k�lc4MQݴ �ȓ�z�8ckīO6�0�F�	B����k��@�m��:}�t�ti����7�a)�Ew��,ڼmnF�@!��c�<�b�Қ4)i�
�{��iJ���e�<� l[$�Oڤ�P��k�`�"O��P�-oǆd ���DZt�"��On}+d����O�>��vlY���� ��@���Ǥ/D��2&� `���w��'*�\�hw�<�7��C���jA�]-�0<��!$D?a+!���O��(hR��\X��A�$;72����J.7����+�z�p LL=58��bs�'ؘ Ԫ��y Th�K�	l:��X��4Ҁ�J\
Dp�k/��5N���J�a��$j0��}!�O(k�!;��GwvȂ`� xT���F�ٳ�hd1G`F-�x�)��t��o:B�eRk��H��/D��!�GM*�8��[�'�h[�FQC|԰��KA�a�}(B�W�An�3�`I�T�I��A�D�>j�.PF}2l��eiB�͓$KN���çfɌ-�2P�V�"Y����M^>��!�*:-C2�O�#s��*��h�&V�w^�h�'�Nѹ�NPwnf�mZ���A�F�=Y�)BQn-5��9+� ��%�\��p�
W	�6�Nq�ȓH�l�P��{��DJ���d��H '�P��J#O����Nv�t$K�Q��(r��Uu�$G/N]:8��&�\c�m '�%&�qO����R���O����D�]��<��Bec�X�v�H�x��4y���Q��LӘ(!�#%��[�G �w���0`C�M��)��� <��A��l 0h��I9�DF�n>H�tI��i��@���rГ�`�Ib}9��IpHx�Q�k��[� ו n���?�2��:�8� �f�#���%p�1ď�%LpLH�'�/7\�\r��J�P
R&~��b��I$d����Υ!Kz\X�ן���&(Z��� ĵ'-$Q:�`�aK��M0$�%QQiR��S
�',@B0e�Mj�D�s��C8� �"D�R��|�v�8�&Pٳ���|U�n�P��<�(�"d��V�.�Ї�eW�T�"�B=�\�Q5�Q?��%Z�*���g"����'_�lp�^6�4q`2I'p@ndZ�ռns@��� ^9>�xd'��&D�T��F�T?
���&pAj`Ztս�y��^9=�j@JףI?_�M�R�ƙzB�ٷ�˛<7�г%�݅,$�I�.j��h�oW�q���!��P~��Ң��!�f��e̞Z;��� �^�{ـ��)�9C]���������MXޟ�+��^1�����_�x܆�i�q	#Ll�b]Hs��/Z�g��,�0�^*8�Q����@�#�4,�(�O5����ʟ�.�Ĝ�!�J�)Ix�C��"���m30',l1�e�-�-��C���4FD�)��8��y��λY��ѹ���Z�؂�U'z�@����z�x<��@�*�F]��D�|���G�^�,�r�$}�Z��UmdۊI�΋C��ţ�%=Vn��o��
���iQh]>{����7jL:y�,�剧)���J#�_�h�8̻r��!&��k�í7����V��>(b
&���d?,k<2��K�b�4�b�/=m@2�Ӓ�-D��K�!C�S�P%0��ZM.�:�:'4\�'�l!�4�E�k�P��)�U��O7
���#�1���[��><2�Ce� ==600L]< t���3��>W0�۫O�	���ߞ��;E�diF����pVkO�k��zpi��+�H߂d�����S��yb��O�ؽ��f�{xȌ��O\6�	����Oo�ف_=g��k�%��?�{��R�|��I�f�=tY��] w�f�9�EP�a��Iy� �<���I1-��CVM˱l��9��1n��Ye��8[��i�C	��q,P �Ύ�]fxuSu�:��(Z�A��Й�V5Q`�A�Ù>��,h��0�'�c�T4���_�9��ٙ�;&���(�k%扻'���xv�0,R��Ӊ�<FāR(��g�B�H!!T }�!M����g�f�@N+��'���("!F"S*q	����n�������.7�h��,O�5O�|��Oގy�t���	�m���SD�h���g��,3�d���y�&��#!�$��	�尅إ)�?12���)�lJp.;}���+=�e��L����P)�/�^�Z`Z.ִ	�)��F݂�I䟴m�A"���혀���	��D��Ml��Xt��]�Љ����p��3���A�7�iݥ#����fi�BE��3� �G�mKa�5/�4<X�D�7_���$�5)zm�2��DIQ���e	ng։�3A�*Z(yac�!��,���� �?+c\\Sc�UWN�����g���b���Mn����:8�re�&��W�ܱ�A֫�p?�Da��35n�1��_�)-$ա��Hfy��Ǜw!���r�����ܴ#m|�`�N��V\@�CC�?�y���(�U�J�'���P�y�ɕA�� 0$�X���#�V�U�BeiDi�B�䡑e��8t�!Չ��C��$`���P�幃��S����>2�z�ZDfW��:�a�*̈�0=)��ʌl��1�&�,p'�y4B��D��$��B-���@1@,��z�ŊHt�8qd��Y�4;�ϭ�hO�`A1�	./���v��K����,L <�%�L�ٌ��BLL�m=
�1䁐Z��T)�MؚX(��G	�	4�yi2ٱ7���Ձ}��D��I��A0�,H%0� ��pnƓB�>�	�!ڇe��t:��@�
�pi�+R�qX&�I&6���Ά�C�0睄t?0�� cɁ�<9��� 7PC�	�H�E"RO�k~r�$D�
�}�ĠX�$�z�����MJL��iPH�er��֚muf$�t���I�ܴK0�\���Q+AqplcS��=ڤ\�$�J�m?�4GG�6T��k�
K1�� 9=�����hX�|���$Ö�pAPV��]KF+w���X�lH�X��Y7a��Uwh��!ό8���ڤY�N1����?bI��gcJ��E���T�{�\�;�d{0�p�&\�F)��̄=fG�,���a�%��/Y�� ڷ'O�=X�L�C�Sʔ����"~~�Gz��.U,ԣqH̨gOn��7H�.��4�F�2{�uZ,^�(��]�$KC�L@n|#gޥ ��q�B�\��M�E�ɏhm����D�<+U��Fi����a��)Q$h`�a�6�'%ll�V�_�1�%������2BƇl���Q#ٓ�4%��˄N�Y�W�I�R�p��h�dD�L�ᙕ	��Y놬\�6�&Z,l��,�= I������E��6� hDP��Ŀ6m��*�`B�T���&�Gq�\�+S&��&6�{���i}xX`��D?7i����B:V� ���Ƅt��,0���k�v7��%���Q�	�jJ���mZ/6�2tj���!��Da���y�'oHر�@ģ:�ت���+nh{�۞@<��� .^w ��@G5Q��Ł� !?���UG@�P%	z�h�"�9x���L�8���!,�8 �썠3!�aZʢ<�̮<�����:&�����!�=��Ls�1,�f�2pm��I�6)�����12d4�ү֬�x�I:��l3c��*�d�m��M�&5��+ѲN���8R�ߋ@�<e��K7`��'��m�TK^h͚2i��J��+�(Z%J��U���#g���g@�3=^ bc/M3Ӗh D �Ms`FF�@j�qVZ2�tC�Not� ��~>)3�������I&4��]�`&�j����IS9��X*C�ܖi����+�:��q�	'7��u�F�8n���b	��p+�b���!��&Z1��P���7p*������ `�ˁ�� $;j|G}�9"�����[b����.ݯ'g��spb����p&��<�F 
3�r؂6�Y+s�d6-��2��HA&��)��1v�	
*l:���NO3>ayr��\�\�!�'jjk�?K\���c�5+0�]�Wl
J�\��Z�E2�q��#]{ʢ���žI^��i4C�O�I��,�L�F��D��Y�6u�DE.k��Y�S��1'V~O`���G
5gD�Ԋ��W������V�/u�Xsf$�.?�|Er`Y"|_�\����:>�fI�!�����K3Z�H�h;�� U`C1B�|�@���'����,��8\R7B�b�t�CLރ:��X��B'q+
�	���$8��ȃ쎔�.l
�b�`�h��;>�H9�7'޵L2�@�Z[�B�#/�~z�q����`����~%~��Q�D�l�F}�5�H����bǍ�N8�N�XռY�Kʪ.#|��1K��o�VU�E�{�fM!�E=�����+p�X	� '��!�0�'z��T���S�`��hF�w��h��ڣO �+4)��J�*y���K�V��)R��R�C�|��D?O��x�Jb?�ԃ��y�,}��eE�k/p!X�T(�"�_:��<�=��o݂Bc}+!K@(=Ъ�Ra��	��- T�Q5�X���*� C���l`���M�M��x�+�6l(;��Ƌ4˔i�=�n݆}~>x�F UbExrHْ��y�� DFb�@%'��!�������@�nH�Ea	!dK���YL
p[1k�V9�� q �LŊ�$@6�|IA�cL�$hI��'���8w��aA�(��Z#q|1�O�+��3`cI�f�|��	��M�@��qz!�̟r����MŇj���(B��5���	�%�'n$������f{����+�vm�������HgDE(�GX�O��6��^�!S�ɍ�����)W�3��x˥�Q�w��.�����BC�L��Xs��+��}b�T�	�Td���#�d��3�ڌaT�X�b�N�;�K5�b<(ckMDc���Կ (�H@#���1�؈qdf�a��D�t��,����#3�����.ޑ�t���IT�D��P]
h}�c�B�n�t����*;���B#�5,q" 2�+e����s.��*2�P�r�"$��j�
�(��Op%�uG�h��Q�I�J�(S
�]t�|�f���:�l�w�A�4�`9�E	j��qC�{B� �WX}@(zT�B�,-KU���$m��H CM�H��2�O��Q֥W'	��Qa����;T杞`Wja���ڛ#���!<Ca��i����	��Aay��c�6�D�I�L+Yp�Taޡz�=���'�
�[��P70(��
6*�9|�n�#U�%�L�$̄?=�*���f���d B�N����G&v����8H8�4I�zwT� �gJ\���[�����9z��d��67ؤ��i��,���AՍO{�8�j"�]za��0KL����'U�Țqȶ��&�,��K�
pH	Q@�o.�aF{⎄2x�v����̉#�L̓��8L`w�ٽW�`]
�F�X���	�/��r.����W'"mX(��
�a�`p�"X�M�Uy�n��obp{��R�ul(@�ؗc��5��6����O�!N��ru�7j���#�Y�l��t,ިTsPh���X:2u��oZ�E���c���	i�h1�w��la�8N=������=���	�<����@��yh�c���G���n�y7��QG+Re�|��!Dy�T��J�r�<�0V��J�8�n�'{4���K��?��LU�R�Ҽ0k�i���$RH�'�"T:1�(1�h�!�,פ8�L=8�i�>��r�'-"��)�.��8d��#�bM�҂����ȳ��#��]	�����O453eϒ9U�L�F�<%#��Sn�3Q�"���9dn�k��	4�&ҸW�\�K���� )�ɺ<�Z-���&_�Hx$K	�B���	ՃH#(��$	�����!&5��;S\�C����Ъ�:n��!�Oн2FȅXtiȯ����F��3��s���@��<1H�sN��Pё�C���|R��~$RP��O�Ҍˠ�*k�^i���I#|���ό�
촢��յ�(�QG3L�ސ��a�o�JA�!.	�t�I*�(��Q��'0���
0~Ѩ�{����l@�)�x�2�I&�\�>t�a�G\��q ���=Y�Li�q�s�RM�60����)B��k4��=,=،�D��jJ��s� �i��U��}E٫�jP�s�4ȓ*��iQ�p:_��}+�H�:z �U�U�)Y8�T��P������DY92dQ��� 7�7��y�D����ÖM -("��{|�9���7e6� �-�?L!p�3J]:w^��3 ��d����BW!<�ءC�e��4
�,��N>H(d1�;'�`j狗ku~A�Ugۇf��͕'���UE�n�U�ǁI�OH8��	L.�������t"�=I�eL0	���*�k�9���B� T��0I������Sm@+r)�`e�q?�cy	�앯G��[F�W?qP~D�I�	l��2����r#c>es�*�!���P�);$��-�-���RFJّA��,���@v��(���j�
�N������f��	���<�ɸ{F��{'*�;'�Đ�a�QT?|${6�[�z���#�Iͨ��yu��0`,���O�θ����W:p ;�bZ�|���/��,O8)1͐7�Ȱ`�T	�����S"�qO�py�)Hm����g@�q�H<�GL~�<R+Ӂf�jl��doa�n@�y�K�+R�`�tX�`�N<v���w���%�"=(ƩǄJ��[G.���4[�f �.����d�	"bFU���}}r�V�8�\<y�
�a��Z��G�`e���0��I���E��'SK��隦`�(O��	�79}4e�4HX�i	��$n��a�SgҔO���� ЫI��IaOQ��ы�N	q���1/1Z���m �M(氉0狈�*��_^��9X@�ȧ)ٮ���v��&� �$�@���s��.^C�a�e��׬m!@��<�ɪ�d�Y�� � ��V̓X����M��:�@� o������,�ժ �R	pH�����MD~Ű���>�PG��m���]�Y;���.��U�Ek_VR��7�˾/"�a�,&X��E�1E�o̓X��]��D�zh�ȻB���A�UKM<)~���]TRԹ����"Z����Ba��Y,�u�E\:x.t �%��=*h!�u"��R^�����G�X������=u�ɑ���8%,D���O�2��Ʉ~8�5!�B�w��i��9��`�#�*�`�W?�i5OL�&P�U�I�	�Hq��$U�态��æZ�����A@��hUb5l��M� X�e	�
�x!k�W���k�8lGR)i�d�/gN�`���=����FD�B����խ�X�ӛ?Is��L�^��rG��s�V��5* a���1��K�m��i�v�T]�lQ���50�@�Ə��n�\����V�n�l�*Ǔ:+y~ܘ���L�<�['*�&L~<���G�J����8s�x\�dӻ)|r�����/N�"�sG�F'L"���6C��Ĉ �?1iTS@M��@{���
�:c�<�s#B1L�ΰY`ÍhU:yb�M�&�8��Kԃ"���i�.��5�>]���҃�Ō��R���S���ۚ����ە�@�W���s���|���!�x����=v���e�z�$�z��A�K<u��	da��w�v��!��V��pXAd&D�M�ΥP��B.ޡIQ��GaL\�.��~&��Ҁ�Z�O��.�?�N��$�>bN�e"��Tcѐ�o��c���׌�I������OH� 6=��+D�	(�t��V�&7���d���C�����G�j0�|R�N?L#��I�$}�f��j'P��ǡ�4P�D�j,��\#�b>
���bU�~Γ|�a[��d)�	,t�	��AZ�{ʑb�t>L��r�0��=����(]�C1�7H�P����H '����a�*5��P���e�
U
=C�m%?e�����m\:L�����N:�|0�5o�j��i�O?e8fh�h;ԘzR Z���{# %D�ܲS�P備6_��.���@�<Fn�}�t�#'}��)_/0D�D�\�f�p, %>-!򄘱 ��	!L�=�X�a�NòBxqO´@�!��0<Q�d�[3� �Po
*&פeC�c�<)УN8;�D��m�XH�m�b��_�<A�e�5 ,���UcQ#n�Y�r�Z�<i����
�f������	>�B��S�&� G��9&��Q!�l^�?a&B�ɩ"��@�wB��7{x��5!�`�4B�ɠ-��Z�E�?C��)GH "!LC�	�!�(A��E'a�ƥ��O��y�RC�ɔ,"�Ї�]:>~��00oJ�	�B��'h�6#�&~R�!#��R�C�IN��H�gK���{fcռ��"O��@�z���"�HK�E`���"Od���᝚r�`x!���gZ�ep�"O8}�X�H2R���1| �"O�9RW/�@"��2��	fXxe{1"O�ceD�x��S���R�~Y��"O�����,r:x�p��);�|i� "OMQ$AL��0]!g��R�"O` ��g� PJ>�8�_����"O�99�� �
!)aC�%=�4 x"Ot-( ��D4�LD *�����"O$�j�FD�J���=)�"O\)���&i@���KP�s���r"O�a���#���X���J�����"O���@
�0JQ�ҍ�5�T���'|�؋��U�He����\)�T�e��� ô[�{B� a[��W
[%o�Z�Bq�:�2{	zw� 9� Z��ݿN=r,��G� wƛ6GX�D���ǉN>�h���5(*�*�L�Zp�i ��E
fh��&%RD��C+N��T���?�V�!N?8�PX��
�Kb��N 1���O�$��>Î5��.�4$Ud�U�H[����#�c��f�n#<%>��f��)*M�j��e�l��&;�D���(O���t`҉�+��A8�?���Q]�X	��)�';u��3J%N���ʑ���F]o��RQ�"�� ��֐�w-Ӫ-S��1#�,�I!JM���	��0|��d�R}J��K�J� i���N�N L@�'M�$ҶO�0��S�m�z�CD��|��j�n�0�f@-�y"�':�dU�=�~�1��2���QUB��lX�$n��A�?c|ج"1a�G~��I��T�j� Rb��[� 5"�ģp�6�C�V�"$�G�ʣ|n�?�@dY"pH4(T�؞\M���E�!��M��� 	�Y���)�	C<4�|q���c�����ƒf��O�e���9��Af�R5���!	��x���|�I!�z�I4aG.qD�� ʨ�O��7�� ���Y��	�"�O&��'KfO��]��&}t4ҡoO�k&�e�!N�' ��b��O�X;I<E�d/��#�
�8�kO�_�j���yPJ�$���a��ʑx�l\���%�`�8$�۔1��O�ŐٴnR�b�b>��pɭ	:P�He�`���$?�d/vӖ	`�y��)���q���U8
=�5*�dP�5�_矀����	�`�`N�%V X4QP�' �(ܐ�����y
ç��$bI4�Y�t�`�ր���Oɺ�'6Z��O%x��5�'If����?�T/��+-6d���I84��C��g�<�è��D?FA�e��5Ԥ1�g�<СN#8�����9o���BăEc�<i�#��.)Hw]V�B���C�a�<aB��;_�A��l����p�Sa�<���ݛMC� � ����Ёs�<�����hH���*��0�En�<!c�F�7A��A��(x�p���(Zm�<�7j˻k��# +ʋ~(�%��+j�<igoP�����d(ʃ����}�<	���R��5&R�L�~t� �
z�<����:hO�x;vL�}S�b1c�s�<�@�}�V�sS�����g�Z�<��O�zaT%���Њ
�fu:�MUY�<�Ƃ��vp�I�����l,�)�k�<i��0YX���Ŕ��&\�'d�<�"⟗`�����b��}��I�<A��ٴfU�:��l�z� j�K�<r	œ8���\�y0P�D��E�<Y��("بIg�Z,h�)�F�L�<�b�;��"'+�9���ٖf�_�<�#��);�k��64��OC�<��L=UU��QC�Є�m�Y�<Y%��`U^���<XXРQ
l�<��C�q]\m�O�#��8J@nf�<�ue�D{��v	ۄ3��ⷠ�h�<!�.2��U��9�t��a�h�<�'�?]�i�BL&3����E�S}�<��
*V�����'Ф=/YBEN�<��.O Z� 11aKߤ^��q���s�<q���&xs�=�����I�-���En�<a���D�p���/ք�2��g�<�@V�n� �k$��kC��pB��\�<ٲ�	�)���I�LA�s�$� ��C\�<�7��={,`x�S�b���0��|�<�$͌F>BsfD� D�ig��B�<y&�@K��!S�aǢ=���|�<��JQ1���D-D 2�
pە��w�<��.Ce^�"PD�'�i�5��s�<A펂
������y��aGaw�<��3Z���1#O7!.�h7�t�<A�g�?2=��ډoiX� ��u�<`@�;Q2L�0k�?ELif�k�<��HNwL��b�)O0U0�p8�-R�<)q�[�%,|i�CS�$��P�.S|�<9Ê�8��(i�錟p}�)�I�p�<q�O�PP����)�XH���p�<��ߛlF\���7vμ@��X�<�D��Ax�@���%g�Beh��W�<9 %Їh*����*�`q8��l�<A!&z/6\X�F�"7u�P�$�s�<��j���!�"y��H"�F�<A�텠;�a�M\	v���dFD�<��۾uh�-�u�̂(à첗��}�<�aҚY�-�V`�M��}
ƥZv�<a�@�Mr��2��W�A�p�v�<� &�vi�%��!G���7�^-�G"O�1�+pc&ժA��:Tb�"OPh�f�+R�J�Ƴ
����`"O�Z�N"%J��pe
>�.�	�"OXT��%8{<
�CM*?Aa3�"O�|���X'\7*�(d�[�N.�!s�"O��ǌ=K֌ HP"ιE0��"O�Q��#Kx�AM�0�B�I�"O@�r���(�le�s�,f�Ըp"O��Y�-D<�8�3p@Ɓ%B��t"O�kQ΍F���nؾK'���"OF�0s,=�6��s��M �1p"O�J�
�'��3��=T�2�8�"O���U��5RE��@�ʖzH�S`"O����D������Y�}ul�j�"O.x+��S,M�~��bE�ztX\	�"O\@�F�W ���"�W�&F�H5"O�8����7U��8Ս����Iq�"O�5
Z�Z�@D��Q$$���9P"O�A�4��$�D���QY�
��g"O\ݡ$�^3m�x��e�<�)1"O��L�A?`�0Gf�!�t��t"O�ɉr@� &e~��&�h�����"O�2�G�a<��$�
l9(��T"O��N�4|��C�'"7�AG"O���S�^�{E�#P4%zB"O)m=d�X�(�,�d|�3��3D��u�ҥz)���R�K1�čU�0D����OL�i��j��ͺ=ѩ�,-D���S��5Wʆ�1�	�,@a5D��#Ĉ^_�B���B2B��A�$�4D��ħY�.�0�pa�L���aApl(D�xb������х�_������'D�,8 �N
�(E�,#��0�D0D�PaS�894�@����2��m�w�/D���nD�َ��č7��y�2�/D�t�+@�jdr`N��V����h:D�H D��%I�`���-D�H��IG�l���Z���-RHV�Q'�6D�:��݀d^������&�4E8T�4D��@��X3�Gg��AU�DL1D�8��#�5u��ɒb	�bd�|ڀ�-D����m
�yy	HP�D��\��Ռ+D�����ۉ!��p���`���/D��h�O�	�
��o^L4�YK�-D��Z�.�7mg�1g^�su�X�	9D�X��l�C@����@|��"6D��rBŷ%�\�r�Sn���/D�XI�D�QsB��Ǡ��0�@�p�1D���g��Y���Q��G��Q/D��Vc[�/�)&�ߩ}&̉S��,D�h�s���r� �Ԥ� ��!p�**D���-�=��3��=P�4D�2D�����4�L�@�Et��eO$D��&�ԳL�i`�.��o�p �<D���!�[�y;����inH��-D����E�1�R�	,ֿQ��e�sd)D��y�N�*;R @Q)_�4$�mZ k9D��
����0] ��`.ۙz���I �:D�@���sòL3eۆYX����9D��j�΃�gz���G��mS�u˗�,D�(G�G�E�^�x�(S�m�dG}�<	C�u�a!�
�R	��&�N�<q��&%��F
kt%�R���<� t �g��604聐��*uul� 0"O2y�@�.2L5k�͎�p���"O�)� �DJ����)t�n�h�"Of@5$�VyԨ�F���6�@�"ON��@G��I)R�����XP��"OT���͍̢��oT=sq��)�"O�� �49\�]ᵭ)'hVH"O�H���R�(���:�(��e"OH�%��a�ت�%��O���C�"O43a@��jx�#X�;�>d�"O�%�q��t;�y�BA�S"O��҅HFyҘP�����9�"O0�ȑ/w�L�s$ �*D�Hԡ�"O�IP
NU���jC�ē 8�IE"O� �ab΅Ɣh�E��$0��2"O @ji;�lp$.R�@v���"ON�8b+�'?8�Q��&�t@�{E"O�U�טX�|ͫ0 N+\�8��"O�i�0�G�4�wn)|j�L"O��LN�'rb)bw�?n@�Ж"O�Uc�$.:M:��6=``ة"O����Љ.JX�Ȃ ��4Y �
�"O�D�	p�����L�)Rt\AG"O�a�gX�R���G��6$�,@D"O
A���{�N]ђ��2g}HEP"O���rf\6^B\�P�I�u�}��"O@Lh�L�;�,\��dĄSh�!&"O��@�b��BJ !�&d��kW����"O^���A�?E���� tL�Yh�"O6$�WЉ�(�S!2���p5"O�@;V� �>)��-�7.
��"O.v�+���BZ��d/T�a��U�ȓ6� ����ջj����"�I8��ć�C������;".�qveڳz���ȓBp ���\	gSVJ��/v\ u�ȓ-t�c��ohF1Kf���x�I�ȓ �<�igI�%�A8���&T3��ȓx�n�J�搵^rD�GA�!@j�Y��_Т��FC/M�H<���X4�ȓ �1ԏ�2+�Y ���9*����ȓ4��0"�Ŵ#�F@�GV�6�B�ȓCX��D앏�|Q���^5v%p}�ȓx�,xq��s+vIyԫ�k6M�ȓau�i��Kͩ}&H��cZt����l�)ц�(~�RX��$��7��5�ȓpO�xy���İ�(QV�n���e�Xy��փ?Ȁ�;�,7��ȓ�pIb!���*���$�.��`��5��E�p�H^���A�J7��I���@ӨT�X��*�憂w��ȓ\����	��Lb2��t��<��X?�q�Q��9zf8����D�ȓl�d���C�[@��cj�z{b�ȓ_�`{ ���.'F��\��z!�ȓ,8^����G�:ƴ��և��^/�I��@z��s⅐�t*=��"�	5����$c�Ð:jzxa�U�ݕ	+R��ȓ5MH$@p`­O���гG�zĦX�ȓrWXp�2���n�`�ѧϜ9����!O:���Z� �峲�ښ8�]��m˔[c��ew
`�g+
`��h�ȓfI�gY�"�D�B��MJ�%�ȓQ��D��؈hdK���/m�z���$p��B%(��Q���ہm�5��S�? �a*W��>�t��v��4Vd��E"O�ܩ �	�3G��a�_�{7���P"O��� #�4g���a�"V�V�ޙV"O�ݐ���6{�>���Q8O��Шv"O���B��su��B�/^��yc�"O�Ei�N�*{����qa���Dy��"O\Ppf��*!�d��E$.��yS "O\����V�V��D�b�xb"O^��X#8��e��*��{\&���"O��ʴaG���	�iK�&qr)B"Of,����PC�ՈqH�m�
�"O\h���
�BA�T�V�� Hg^,�7"OH�/�d�[F ��Y��B̾w�!�d 	� �  ��   )  �  ?  �   +  �6  �A  �I  `U  ya  �g  n  kt  �z  �  3�  v�  ��  ��  >�  ��  Ĭ  �  I�  ��  ��  a�  �  ��  ��  ��  ;�  �
 � �$ x, �2 �8 s<  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��Y�1/l	aCڷUClM��%ɘ��n8UZ�&]�KR�P��,%T��<A����!Ez��F��\���i�L�/Bl!�S�t�3�a[��~��	9"O��"��IvH�	��EL6j�"�"O�aY���VAv,84jٟ.��"Or�{��+Q���A	L}>q�e����D,��ʆJ��t(T��43 �B%�!��/@��*e��-�tF�Q���hO񟶙��$ڸj7�7�B�Z�X�,D�|�7�g�Z���\� �~���|\�S����M�o�|P�L�"��uȨ�Z�'�L �r�ϓR�<H��Q/_��e���$*<O249��G�/{@ыR�%2��Se�'F�,���s��P5�!�s��5E~���b��ex���*x��ᐦO��HO�����`h%���a���
T�V"O��X"�@57�R�6#�^vʸ��"O0d�7@ 4i�8![���Z[�݊�"OaZ��R�,�"�;��T�xD�9X�"O�#�EMd@R�+F
]�� *��'Z�̈́	�dlqi۹&�ͻ���z���$=�����"	t1�.r��'�a}�c'
�ǓE�T�8c��Ұ<)W�>�O�����mF���& q��I!���F{���(aDQ�p�"Ǵ���-�2�1O��̓�4@�2�3�  ��B�G�ecʜ�R�.���"Od���/Ƽ2�K�Ȗ6nƲ��3�O�=E�TV*�\�b�Z,�T�k �N��y�J�v 
8��&�b��,��y2�
/B�R�x�k��1����jD���>��O~l��M�Vk��8ċ�4$��1�"O����B�)G�"8ȡ*�8U(Aӵ"O�l�E+Y�U>�48�Jӡ/�����"O�-r@�C�\ ����$z�t�R1"O�����'6��]?Y��R"O��³C�&���	¨|����"O^�{��G�
�d{�"hh *O�M�5g¤%�-ۃʗ1)}2�H�'��Xp-�� �\t��m�kJ���'ڴ���"F�<�b��$����'Hٲt�S#����!�
k�ܒ�8.*�6ڰJ獀�6vP9I4e�'@���m�|yZC�%x]��N�����Dz��~���IX�Չ��^k0NXǎUd�<���F'W1�%I O��՛"�Ҧ?�"=E��D��I���5yb �`%U;S�؝��B�z;�Hņc�6�����d�,T�'_a~���T_���+��X�<�j��L��?a����8������(c��BS�9+q�|��]fI�����ht4tZ$
v�X0�'�a~���[K� �	��C����᠂��y�A �f�\�iS�n�*����y��K"��0ՙj2�䫓bR��hO%��)��8�4={�I	
kƞ�v`[:*�!��·|&�!B��� "�� �ռ7�!�J�`�����<�R����t�!�A�_�t,��-�'!��;���|�!�dӗg"%pEhތ�2���jȓ�!�ɲDEz���$��o�ӉĔ=r��x�㉳	xR���7`�bAj�O��
��dh����i˹2s
��)���&#D�`X0�Db�����ᗘm-z�j��?D���"*��Ae̍�C׺r�0�鱤(D�\E�Ґ +��)i����㤟�D{���H%��1� @Yh&�A� =!�$^�yUVxi�V9eǒ�Sr/ފ6�Ѱ>�a!�[}���U����k��A����'g���r�Np��d�{�l�X�'���:�/��{()q�R�v����v��E{�'99�\B���T�]h� ��z}
���9�TPh��/f��PL.s?6ɒ��9$�t[D��
K�,���(�X�Т�#LO\�@�"J�O	<�PSe$*^���a5D���Q$_%&|غ�)�5.�;�G4D�d�Ǝ�D�Ea��k�d�)�O1D���$ޠ�����H<P8�H�ƭ<�$�:�S�O8*���~'L6��*��i�"O�$�LUaa�q�ƦN8eLy��$^�<Y�~�R�� �-I��{Ώ�"`���	J�	l�@b�j%N�

��n@�8#�'k��4	ҏu8Ԥ�TCֶ6�L��˓�(O��#�1d�����BS`!1"O��@���.�HU�1GR�eEޙ��>��)>�S�'~|mc��ǃ>@>m1��@�]Td�ȓs�\��Eő�2��Ɇ���̇ȓDz�8`�Z�(�8=���B7�0�ȓw�.��!�U$��Z4E�}DD܄�`�0��2Þ0�쉁ōT�(�ȓ' @����	$Vd�T��	�v���S�? B!(d�ʑ�xǁ��W<�D�xb(/���%��1��[&H�8a�"N>4�F���i?�p�ҒR7�m`�
VUԵ�EK�<���+���p.C[qK+���D_�Q��7�eq���H�)�ȓR@Q0���*���� 6D���ȓN��U�@�ƈu[Q1��ο"�:%��@��Ϟ�D�fq�(�or�ȓL 0�	AS�8�DI�F~��ȓ;����g�ӱM��0�i��;�m��}�|��GMQ5
�-X���&T�(��n�Z��@U�]d=���д��\�ȓ_��e���΅S��!��.'n�@��	c}���.A	��0�!P���z@
��M����s���C��5!�m���	 h	�"OjiBCN��l��B�]�!�f�)�R�̅�	,��"�j
�>Q�P�����~V2B�IKO�
�F^�%v��%ƅ�>SDB�ɞ|��D�g���d`�h��+B�I6
P�S5�(��!h���\��B��ӟ��'L��$(J���-܅+/��P /*ʓǰ<�� �Tx@�1c�D�+ƭk�'g�I�h��h��Ͷ	F�B���(�MD"O�}��%�, ���U����{I�<I����b׌ѓ�"ڰatz��[��C�	5�]I ��D��=� ��;�V�=yÓR����G��<��M�`,(�����?7E	2(�V�ì{��=��Y�<�A�We��}�֪��5��=(�ZT�<aWob��r�LN�3����FS�<yfɝ7�*�:��Ͷt �h$Rt�<���؜9�Q��	�5��9b)�o�<1A+U�����F��!шP��j�n�<�U!�2���boӱuH�]a׭	g�<��n�9���I��-����/_�<		�7.�����f5�dx# Yv�<�w�
�������*� 8G�o�<I�i	#�Y�^�,R(YQ�"�E�<�t��!Dk��X%����t����y�<Y3&H|�6p��i�D�0@��r�<QT	�Z��r��+�0%!!Ak�<��&G�k����� ��'�	h�<i��$`�zH��b"x6�Qc�k�<�a�]T�t�tMU4R0�a��Ap�<��E�&F�����
8`���u�<i�I҅D�����e�!21,�Q5��n�<�GN<����F��_��#��a�<a�c�(��q)��\1JM�Qx��^^�<�E�|����挭.�&�P�Ht�<9�%9\����$G���q�p�<�r��1��u����R5�ea�<Q�щh���Z%K��2��MD-TZ�<)F��~��Tc�#�m	�}��V�<�W
�w^콂 ���d́'EIN�<i��ع"zB��@�cs�:��H�<�WMӟk`"-�S��j��
�Z�<�V��(gDT��@�=u�B}��b�W�<��΢<˜�����`2Q��}�<13埦ZN`��N/D޸�p�O{�<闇_�F��,�o�vG��R��B�<��2u��8#�E�_K���"E�D�<�Wʄ���-I�ਂ�&G�(B��1"&~H'\�W9��!���QBC�!Kz�$��,L��,!'d˰ �C�)� �����E\�k!��$SH�"OtM��imƴ"@N7 OV��v"O�٪��`�;r�[93�@�"Oܔ
5#ԙg���W%O/\��@"O� �tl@�~r XפM>$�$���'�2�'r��'2��'KB�'6�'�@�A�E(uYT�+���(22 �!�'�B�'���'pB�'�'8"�'�H�"�Ȃ�V ղp	�A�\�r��'���'���'��'	r���isB�	ߌ5j���F����o����O���OJ��O�$�O��$�O^����Oq	aP㚂��!CcA��$���O����O��D�O���O��$�O�d�s-J(�w ߲���+	"��D�O��$�O>���O$�D�O���O�dJi�\q2P��)������{�V���O����O����OD��O��D�OB���<~�ܻ��� iԙ� �7���O,���Ol�$�O���O����O��m�Z�[K\"� � ��8dZ����Or�$�O���O��D�O����O��_�Q��8l��5�i���@�����O����O���O����O����O��d_��8���M8�����'ɘ�d�O��d�OD�d�OL�D�O����O�����܉��U</b��k�;8����Ob��O����O��D�O��D�O���0+��e8��
 ��s'�A�����MK���?Q��?���?�׿i���'Z����Cʗp�~S���;�K����������$[����	1 0
�Ěs?='D0Y�-)?�3�i��O�9O�$�(XFaz0GL6�xb��������O�4"m� ���$$��O��(c&ķ�`4H�gO������y��'���Y�O~�2���"������C Ǩ!���t�Vm�F�� �ӻ�Mϻ<���7i+4��`b)�1Nx�|���?�'��)�S�"�n�<�1g���#�mC OB>,��	��<ə'�4��ò�hO���O��i��K�U�0]���(q�B��7O����"l�L���'����L�0ghŹG�R�qs��j}�'�29OT�Zx��Sr��nW�xC�F(�0�'��&ѩA9�)������,�B�'�P�J�>S��\�q���8G�)�r^��'F��9ObH7G�X�Ν�E�P!=w"��q3OF l�3h�
���&�4�f���B�ŀ���-aD @�4O���O��$�=	
7�6?9�O���
+�y"Ɓ��F�ND@� BGvh��喺[n���HI�A
�ᄑ!IF��$$�3k��$�"GS$&�yS�4C���`�%�9@��%�}I�*��l��`q�g�?%�ݲ�oL�_��k���LF���'NҖ��d)U��M�U'��xE�l�(CD1��٘XM�!oVUҀX��n5��)��ҟ�>��d��*WlF�A�ܖDGt�Iˊ1,�f��b���0(�%Ŋz�T�b��X��@���\Ej��͇' �֕ ���
�`�h'��f�$(��D&���y�AZTh�`+R�J 9�;�HR ib��������)�I��\���?y��One���0�B4�����!�Ru��iU�'�1S��'��'{b�OF�'Hc���S�k���cפH�.��m�H��4�?!��?��'t4���T�\=K�tt;ӠW�=Q�q�$��m�7�L���P�<��۟L�3��џ��qH��r/�U{c���������M3��?A����q�@�x�Of"�'�ʡy4.��SSΩ���\�!����`��>���?1Ң�B��?���?��Έ�@<BĢ	��P�7a��s��f�'�)��l<�4����9����x5"�.&!�T!�픵�g[�|
�6�	�d��ß4�'��HeP�(����,ڢj�v�
EM�	$� O*���Ot�$�<���?y&�ԱF�"�C�\�C�%��B�T�J�<����?�����䅱t�Χo8�����Cpi�%�C[?i�$��?���?�(O6��O�ȋ�_?�C��J��%[Ё�����pF/�>q���?�����Bg
�$>�kG�λb=�v�:�����O�#�Ms���?Y/O���O<�g��эr�3'��>��m)M�5W����'��Q�P���F��'�?!����B̽W�qH�P.Wwn��ō�Ħ��'�b�'I�ܘ���⟛F-�d� ���%`ݜ�!%�Ɗ�M�*O�������UX����������'D~�ʆ.��9� ���c�4�?Q�����*O��?OVt����:��Iש)+����i��j4.g�Z�d�O~����$��_����ucկ��ؙ1/(b���M����1��$�O~�$��1O,��/{��0Q��]e<����@:e�f�o�˟���Ɵ\��і���|����?y��RP��l�@&,�%�a�����Ɵ��	43.b� �	����I�T�*,A�@ u!�tڀ�@)�v�S�4�?�D�Ě:����'w�S�(As`��?�Dq�5$C�Oy�(� �Y9�M���FV��<����?y�����@�C�F�#d�I�,��P�cJ�!K m�i�|��՟D�I�0�'V�' uSʇ�D>�<s1FF�!v���.ٳ��'[��'��؟p��KxrcD7������/�Je�*妩��՟��Im���?� G&{k�<oڌ5�t8��b���x�s$���듃?Q�����O -��|Z��J:�U��+E��+b>�b��Mכ&�'+�Of�D�'Cc�uוxb"��`���׻.6ͺ�'ڐ�Ms����D�Oj|�a�|2���?i�'u���&MP$��h�foR6w� �(����OpC��G�>�1O�3� � �e�n�2O��[|⡘$Q�,�I85`���I⟴�	�d��yZw���.��,���h������O��d՞��#����aR���WG�~�|HW�LԛFD�Y�2�'���'���]���Ɵ����۰g�P�iC� fNp��˙�Ms���D�V�<E���'��8�`λ'N�����g1� "%~�.���O��$A�i���|���?��'�.�W�"L��|�Wf�4H,� �-�I++z�E�N|����?y�'�-*"e_)I��;f��?N|���4�?i������O���O��0s���7T�P偕�x�Iۑ��>�YB���R�!?���?�/O0�䔫!L����R�Mw"���KܷlZ��Ф�<����?I����'hb x�|�8���(�U�GD�o(��%$�1��D�ON�D�<I�66Dys�O7h,	��m3(ڀ	���Y`���9�	����Ip���?1%�Ԯ8p�-o�� Cҝi����,�����?����O2�)!��|"�'xD��פB��1��)��sJ��
�4�?��'l~�P4o���K��TC�+ Sh�$"�J!8_�Xm�ӟĔ'WR�1@e��֟@�I�?ѩ�o�!� �I�O�6���D�S���'�"�@�zxx�y��J���/�̈!#���=n� �"V�|��8M��P��۟���՟��SQyZw� U��Ԩ+��)����|1s�OD�DR�Y����O!2������G-�J����W"Z�6 Pc��'���'+�$W��S�(�wN��uq��p�Y�d�\!�����M�gfΏ\���<E��'N���7@ �Pp2��#�P�6�g��x�����O��2RM�<�'�?Q��~�յ{��I�R�4YG����2B�"<�����'^�OB1H0m�85���G+!�v QR�i"
æ���П �����=Y���	bV,�Hq� k�b��g"�z�ɔ)���?y�����O�����O
C�@�p��6�
T��Rt;���?1���?��b�OZ�90j^�o�d}@�L q��PP��i��0��O��D�O�˓�?Q�cG���T.����ՙG	� H^�e�R��M���?����'crĒ�O�`hp޴+���VȈ#-�u��#���'j"�'K��ҟx�  }��'B�iY��.�`U�0�"X�f�c���D7�Iޟ�擆	?�O�0f.>Q�A�13W��h1Եiy�T���I�R�	�O3r�'��4%L%-$��i�;:��9쉟WJc� �	�*�>Hk�(�~��H�c��y���k�"$�e�a}�'����'��T�\��FyZw�\��¿V�4ܳ��.1(�p�O��d��\���r���	0%�&�Q-V[���T� ���c0<B�'�"�'��Q��П���͋��P���B���[��Mk3HьU��m�<E���'^^hɇ��H9�D6�C5�~� !�n�D��O��$U*0!F��|���?��'����:��a���T�:8�a���'&V$��C2���O�d��|u��]s��d�C�/LbG"f��d�:�N˓�?1��?��{2��7�*��A�` L��aղ��C'C��������	Ο0�'��,Ϸx�� 8���?�zt��ƙ]O�0�g]� �	쟸��q���?Ã�(�r�z��.&$�0!��T�=���r�ÈS~��'W�^�4�	�����'&2�	%̋!�bm@`ɕ-M��l���p�	����?���<o2E0�lV�A�3��N�� c�^�0���>���?Y,O��ă!i#bʧ�?ׅ��d��¦�ֵ}�4����N���'��O>�����d)s�x�C� ,ϮL;� ��xE:��`� �Mc����$�O)C�b�|2-O��I����&�Z�$y��Y,. �>a�jXp���Me�S�$���`'�Q�q,W=Ȇ$�hɋ����O���$��O���<�������8ժ^0S:��XDB�)R���p`[���I�~��m9P";�)�S�IH�!7�=*�Ȅ�n�;2`7�7����O��$�O�i�<ͧ�?9C"ɑ`�V�+t�	!�z�a�튔F��Bz�Ś�y��)�O0�BT,�V�`{���x�,A�p�ᦍ�I�`���dEL������'��O�]-�T��s�X����fx@�y��X�E��R���O����I\1 �%\�.�x������b7��O��3��<����?9�ĸ'w�5����,�1"֡3�噬O�LybaWoN��蟠�I}y��'�@�z&ۺ2}榔-U��[BE;g���ٟ�I埌�?��Q�������;y���%Lѕ2VL�������'J��'w���4sEGD����
�ذAǈ�'���p������	ٟ��	T��?��;�In3�Is�;(��yGΞ����?Q���D�O^|��|����<�Ԃ3+PFm4B���ـ��i�b���O �D��~��'Y���D!�X:�<���M7fbJ۴�?A+O���@�xp�'�?���J�i�b?��r͛ �S�/Y>�O���Ϗ4t k��T?H0��+�Z�ga<����>��~$���?Q���?�������(a@l�
�u�o֞0�"(��R���ɓD��x��6�)���Gh�{��!��a(1��07T6�Q�P���Ot���O��)�<ͧ�?	A��!n�ԫ�E�j��aV�T?��&��s�>L�y��i�O�5� �� ��>p��s-%|if�i9R�'}b�-��i>���ɟ�v���:,Jn�1t#T�k�>Q�P��/���$>������I�Qs�=���Vq�%e�^4�L��4�?��n�*R��	Fy�'��IƟ֘�s���q��;z���S��TV�p��q��?A������?i)O����M���a�啻%\��� D't�D,�'��IПĔ'�2�'@�T�)i���cD,w+��A�ʩuTT�r�'N��'tPa�p�';�T�r�������B���[p�X��ؑ�M�)O �D�<���?	��u���4����	Y�`��=��+��?�p}�irr 	���'_�bb`ѭ���d�7j�٫�,�Y��J�-@�*�(o�(�' ��'�R)���y2P>7��^K [�ą� ����6�Y�����':T�0З�S��	�O����Z-9"K֐��A!�)b�:͚�B�a}2�'��'�F�)�'��s�D��a�6}2v�Y��X����6�m�fy�癁w�7m�O$���OZ��b}Zw}�5���_�4e^`q��;Jx���4�?a�r�H����$K��m�}��&�c�`\Q�i�,q�`���):�M���?����pU�4�'I��C��|����e'<����nӮ�t4O��D�<y����'쉳�\��(*0�����ͭB��&�'"�'*�����>q(O��ĭ�t�G,�tz@ �6���m�b�i�oӀ�Ob�3�8O��� ��˟ˠ���ر�ӯ�(��9��I��M��> V�$U���'2Y���i����hȹm�`����)���Zz��!�FyB�'$��'�I/2��F��(^Vظ�jwU@��F���ħ<�������O
��O�M���ǅ�`Y'��#��P"��S���O^�$�O(���O�ʓU�4���;�|���NG��I#�/0�дi�����0�'���'�c�����W�{�љ��,v���Vf[�9W����I�ȕ'�r�E��~��{bT�7�٥�N����B76�8i�&�i��Q���	��\�I[���Z��4z�f�ۦy�AW�C�Tbڴ�?�����QQ��O���'��4�Ȧn���Jץ��"���kZ���?��?�]K��|:B������q���j�Q�ά�SS!�Ms(O��Sf�ަ	������I�?�ɫO�N)��©F���I�f��]r���'Wi���y�K�~���O���l�.�>L&
��tX�4N>ir�i�r�'B�O����򤊸l���Y&�>=X�˳@�
���m�R4~�۟�I&C&����'mV�q�_*O-��MI�qP�A�i&b�'�2+�##����D�O��ɇ<��tK�J
N����%��6c�7-�OP�/���S�D�'�'��#&蝁A9�󫚝zd�eV@}��d�7}�X�'�ʟP�'Zc�>��f��Cgܤ�S@�g�$0�O쨋w7O����O
���Op�D�<�C^�Ztԉ�E� 9��VD�irW�\�'��U�X�I��0�Ic�u� Bs���J�L�&��)p(|�4���X�E�˟H�	Sy���"�擲"Њͱ B͓1)�av*�f�0��?A���䓐?I��+����iŲ�a�Eo�j)[�""}$���X�l��柀��Oyb�r]�pI|�a%�V �3�lы2o������ro���'��'���'����A�'��K���ѡ!�%+��L��p�.�D�O��9��4�a��4�':�4��8�z�(3揑<X�B�e@�l�Oz�D�O���A�OȒO���97�R���L..<�rI?�r6��<�� ���/�~�����%���1S#� /=l���f�
%��A�`�h���O��ХE�OF�O��>)�#�Ȕ^��՛��_�~'е ����o�����ğ��$��'V�p+�Ǝ�f=s	R�y�i��y��qp��O,�O��?1�	�0��Ӡ��F����H�Ꮈ�ݴ�?����?)Rē��'�B�'�X�Jΐ۱�ʶHI4�#�[i��|���3��.���O����=jH䓑nA�/A$$��읉t�oZɟ�s�:��'��_���i�E)��!�DaEںP�C3M�>g*��?�(O^��O>�$�<I�Ɂ(�P��,��,� �Yu�݌�@���x��'z"�|��'{"�Џ0sl�xE'�{{����\�f�c �'w�Iϟ���ҟؕ'��� 1v>����.(Xj�ђ��.\K�M)� �>���?�J>����?�&���?󩃼mJŢ���q��#���+���ܟ$��џX�'���[��'mƽ�N�o�u`�D�S���D�iy�|��'x2�R% b�>	�ې;�<d۱�<� ɡ������Ο�'�"�y(���OD�	ِX:0r��U%��+�oN�"���%�\��ܟ��``b��&��'8��1����eQ��[RD���mty�& "̀6��[��'#�Dc(?���M2�5���3,�4IEm�֦��I��0Jr�Aڟ%���}z��Ǭ����hV%ۤ)a1��Цm+��^��M����?!�����x�O
f���S�a �*A��&�L$�`�s�x!1M�Oj�d�O�uF��':q�΀��
�I�M�</-$���pӪ��O���W�/Rn&����эU'y�ħ=�bY�Ʌ,"u�֙|��/Q{������O��D�	L|>r��J�ہ� +��m�ǟ`
��T���|ʎ���#A !�#%�#��`5`êb�6�'�"���'��	� ��ʟ\�'Rh� �Es�cH1��
׬N�;�F4#8�'b��韰�P��=����gnۃw%��� �.yƴ���}y"�'�b�'���'Pp�۟ ���!7\�9�c�ة!�(c1�i��	şd$���Iş���$�4�6-\�]�f��1�2\�2]�pj+�������	ß\�'W��Z%�~��[�R���ܫ$P�(&�>b����V�i��'��O%ڠ��ڠ��@�ЦZ7�uHDhX%JQ�f�'qB�'�R�H A5�Sly��O'��6l�VR>y����Fk�̲l&��O���47�x0�"�T?��gA��@ �	�
l�\��w���d�O�Q�M�O����<��'�?�����
��b��$���t�XT���Y�	̟�� �45?b�b?]��95`	��ɸ0����"ii�j���R���	�x�I�?u1�O˧n�$��k�& ��(�H\�]�G�i*(7�D򟂒O���/e^J8!�oˀ\�h�ڑ��=����O����OH�h�<�*���䡟�Z7�L�:�c"��8M��١h���'�:L�Q�:�i�O���O����k��=u
4)c��-*�H��@��ʦ�I�,3n�'�T�'�?�L>�.D]�lt�ʜ�
`�',9v�	�"	�Aг������4�Icy"-/y�́P���./Zœ0����禼>����?a���?��Ț�?m��30�O7k�DU�P(�+f$rY�A�|��'��'�b�'���kf�'e�� �W*�ZP�d�/�����x��˓�?�I>���?iB��!@9�mmZ�U��90W��I
�2����%�l˓���M�Xx4:çKT��w�[����!���c*���ȓBN)��NL�#��{Q.��Z����JcV��v� �*&��"/����w�e���ǉ��t.6�RC�M�G��"AA؎V���C`ƋK��ؤ�^%$x\]�6o�#:�L�
@�{�0���Fאb�L� ˑg�X�&��$*���7"Tp�y��%^>ap��F^<�@2!Z%Oh�d�Ab�
��Ⅾ:��f�O����O��9TBS#qC�HCd�"�>�80mKtQ�c4\�$	45)q+ΐ�dH�O�1��gG1'n�ݐ脩d]`��¦<wy֨�q�W)�"��3)��k��ɭR��pn
2V.����9a����%����c�IP���䙓��	�X��'��+����FX� @	d��<)@0�ȓ[n��P�E�U��Y�Ě�k�Fx�"=�S���#��9�
�vQ9QNנ��'��1�U��"�'��'�v���H���g�ԑ��h	o�^$@���R��PB��C�4���g) �P���?�=ٓ�S�Iy�0��(_?}��-��
^�B��.u��=J�@i�g�'��qKҁB<X���xf�E�t�0K�'��B��?Y����<�Q�	''��zg�/v�����	�Z�<1���
��`�[*l�D���㙓|������$�< �o�J����"5XX�/G�uY~����t�	ğ4{���Ο��I�|�1�	)@�>T���Y5g�"m�@ł�V����,�VT�z�_���<a&�K1/8|K��7�$YWIv�7��>)�t����-?N0��	�)����O�@�'xcB��D��"��`�7ړ��O� y�Ȥi�0���$ V͙�"O<4�� <5 h1��޺�Y�9O�=�'�I�55��s�4�?������8�
|�7�ԙ���;-c,H��-�O��D�OP��!�z������S0~���|*h{~MK3͂(~�� �W�'b�CnCC~mb ����9)dN�ﰴq��-��i��݀K���C!\R�'�%��Z��gl�"�D�|�$�KW���C��ͷF��02��?1���9O�iP�ۉ&�ڵ҂K�8Ln����'�O�\��G�kf���)����K�6O�rv�Φ���⟰�O$�D�'�b�'HT����g?����l��F:����XJ"�xd5�T>��|�IS*�M�vA:9���gƍ�BV$��dP�X��D�J>E���x���õꂵ+".(� ��	�rԋ�	��?����?������Ҋ]�{�UP NK  ���Pҡ��y�'��}���9k_"�b�Ǽ0�d)�/��O�Dz�^>��B�$�i  �x�����ß��K/��������Iݟ��	'�u��'4҈�v	r`�B(�b]������~�f�u������ɝcFB���	>v����ʐ>$���ńpw��I��&H���K�@<���ˁl�꤂q�N�N�ָ���ƃ$��Ռ;w��mӪ9l�V��a�S,,�楙q#ŀHRj��`h��izC䉥u�H��� �|H��3V������Ē}�Q��6��'�M� ���	:���� �Sn��Ā��?���?��t��8���?)�O=6x9�,�>�͙4��.��(��ҍ'�6��(X�~��X���'�����UIӰ|y�"Ğ3?$�#N�oTDB�.ֆK�$H EB�	������dJ�AiR�'����E,K�b��ѹ1� ��'K�O�}Γ3k�sʟ����K�ŕ?tTQ�ȓ�$KgC�<X��ӤK�>�L�����qy#U�N�7��O@��|RgOF��+f��89��[���	F�5@���?���=�`}�c������ �|Z����HA�@̕=�}�S�	6y |J$ڧD}li�B�n��a��c�<#�R�Dyr�Չ�?ɋ��@�s����Ƨ �h�0�g�13�!�!_
���:��('۔�a|��;�R���X�ģ	�M�xDJ��T��H�p�TnΟ���k�T�ؘE0"�'��
�	G� ��R��7�4��w��+`��Hi���'�ia��M9H1LqK5ͭ~"���;*����@��:���GEеUTn���9/c���Ŏ�I#��փ���>��'��tم��<M\���,�Cϐ|�Ai�O���"?�[��?��Ժ3P�Eʢ(˕'�^H�3#��<y����>1w��tF��;GH�z jR��A�'��#=ͧ�?�Cއx���:��Јn�@�Q�&@&�?���J	�\i���?I���?)��j���Hy������M:AfQ]d�ré�����*�"�4yaE��p<��b��*��sD�ɦ�\JaY]?!R�?@o��fg^
t��x����B:�j�#��Z#�� `�: *�Ð�Fx��'n����O��arX{�/L��YA>���ȓr7$� f�``$$
R�N'O7V�Ҁ��}�$[��P�o\:�M��	�6�xep�f�3[����#Ā��?q��?1���������?��O�Jh��O����ƚ�}^�� �Ɨ�Z&E�EXY v�ٖ`��0<I o�7$�:t3���('*��@N�d\�����$Pl
=ˢރDjP��	�-&���֦���E�/���`�,��D�"$��M˻�M���/3��<A�He�t�a��"���#��HP�<����?tH��Q�i>|�cr���<���i0[�(Q����M����?�*���#$�K�>Iq�%�p،�2�±9���D�O�����$*�|�&�7n`��eם$���ٷ�r�'(���ӳ8���d/��k슁H��)0�T�<!�N���IF�S�pƧ>sx���0%W4ef��T������?E��'�`|���%|�5�[g�R1��^#�'��d�gڤ(�A5�������'!^���{�����OF�'0�R�����?���p(��ڤ)R��t��u_�1!
�o6��'�>{h��Ȧ�'���?	dl@�t�)!BldQx|ˑ�_�@�� y��U	�:5�E�",U"%G���r ���\��qyg.4F�|�1��?yC�i���'(�O���',�A�D䠱��U� *sF�ֲJ"�'a�}b�S(�4��'�Q=K��U�uŒ��OP�Ezr��>I�MF[�ji�f
K#CؼY�BNݗ��xB�=9�d�)D�i���펛�yb��2r����Ψ`&�� "+͡�y�l9BvyB��U^���E*�yr��W�Z���@�	
򭨑��y��m���d�C' �N�pj'�y��*����F(�0Dڄ� @��yB�� 	�)b�k��R�t�1"���y�#T8a�� #P�4N��b�
&�yb�ϠW�̪F&��x��T�G��?�ybjS�\gj�5.��l�֠���ʄ�yb��fR��3�	�f���+���y��?g4��A"O�Y/���K��yB�_�#-dtZ��@�Q�l��bO��yb��.8e$U)���V�D��"K��y�g�]�.����	\0)���yr��8�&8�'J�$�s���y��@t�D+���%r/<��1���yBbM,i�Ldǎ�9l�Ұ
���y2G'w�,8�F�_k�8�P��y2 �g�*�BrbH�h�RYć���y��>��S �[8]��ICc)��y��F^R���*�9`>����@�y�a��.,F�p��6\\ޱar��4�y"��]��Xs��T1V�ٱ�o�ybh�
�R��2�$ Įţ����yr�	�w	�m]1
*P '�y2�1H���x�cB��,S'�ͱ�yb�%ź	h��M" gF��D���y� @l��#��w�� ��y�J�#J%���Vn"�9��>�y
� ��[S�ݴe�psj�g�\ls"ON�P�ʚ�
)n,����\�$�A�"OZB�[ E���	�K�fc "O�0��,��z�N8p��A�t��"Ofa�h"�������#�,� F�>QGAW+kǦX(��`�"~�#����1)��Ց�l�Q�*G�,���Ol�S�"W�?����r^K��x��˚8z�@�.M�mc��H�C�s�<��U�8l2�»d�T�2K|*�eĥ7I��長u��JE�H:l�(��#��HAP,�℈�4�����z2�Љղ�O�KGo�E�H [֌_D�60��%.&F�RP��xCrb#n���`dj��� ZԈWd�60$�����״"�Ʊ1��X3�(@D��?+oQ�L��$�-���<Aʐ*��'�"����6�>���A��D!��!�>n� iq�*y�h�5F$�|B63轢9�AB2V0��v�=����8
F�7B����фQ��IG�e�e^���eI𮼢!"ضn���ɨZ.PAф��)^��L�Zw��x�7��+�4��v�>��IC���S.܃}94M8g
���3�c	��?ٓO˴n`�%>�y�/��-���"�[�T�(E�'�[Qyjm􂓷N�\#��C�9����Ɩ �8x���UP�'��e�O)A�ltKGO�c�Z`�ۯ?H`�Qb�^�4�xb6*�Ev�ܸG9a��T
�K�"#�ɏ�`�Sv��p�8j���0�ƨ�V
"o��IF}���&ؠIeb��e�!�p�'�ּ�@dN�*�!�ς�l)4��`݉M����%j0jx<Y��jq���Dl^�]�� �O��睭I���AJ�p��PХ�ơt;|�T!|��G��#)���3���h�F-A���^��]�`K�:��a�Dk��<�E��7�����A
<�Ub�jP8�mc|�'��!�<[J��;�c�h���Z�� ������'�ƨ�����ħ;G��)]-s�j<�P�U��y �T,�(��(C4$!Z�-��G�~�C�ʜ".	2EA���Y�5��S��	Ued(zZ��$(0����(�区�<��I�B#�'r�=����)��u9g!�8Yr(����	�1�<�6�,���#�Z,ml�%�K>�?A#b^�*�]Y��;y�*%y�-Ou�.���{�F�?嫂NԜ@纀д�Vc����cKְ�=�L�H�ˎ�!��8y��D7P��ϐ�l�rʆ�g��iI�c�n����1�6�����#���=���1�uw��-_^�a�1.ʆ3��>�<qvRc�H���.>��1�o�#� Ton�y3��/z�L��̩?� �y�DR\���Qc�!Wszx9A��8;�@5"���Y�p1���S$H���I�NvX�Z�A#>s0-�'�x��4�`���EZ��o�%�b��?Eb�� �T6ݸ�lA9,���Xq�_ư=)��U����1n�b�� �A~�0�֩��|����(֙q9�]y�,�e�O ��O,Z��XI!s��;1��bs�͏ɘ(� �	3e� ��F7�u��P�_����L8!%��W�R�P��P=B�T�#�Ĕ3�~���o������቟~vŉ���n�9[�a�,M8���shG�(��
����Ѐ뺟�����AkL	�K�F^r�23��yYph�΄ 1<�~�a�-g�&���l�}@�jA"�&���p�'; ��"D+R��1�O���杻��X+����E�
|s�&U�*"��䋳v)zU��ͯ?̾�[�� �~�|Dk3��s�$U���K�Ez�!g�H�O���"҇��(�&�%?����\�d��1ۑ�N3�aإ	*ʓ�����L�$�0ٕ�^R��`��?�˅Hv7�z"읬+���!!�4����gB��x�jZ]���g�'�
�ZG,݄0o����B0{I�y�JX�H
����5D����ְYҸ�+Qm�yü�h��
Z�n�!�ۚRU����"_�qK��'=�n�r�f	�Uo (���D��ʓe V��O8�q+�+vK�wF@��͉70�*�k�ḿ2�2���'�.���%��a��QfC*9<����ҭ��ɦ�y`%��O��S5$J�w
�$9Щ�h%�I���V6D���'㠔z�/7'�Y��O�<�"ŕ�8۶�	���!<	C� �m�\�͓ �n iʃd�����O���Ȟ���Q"ak.j�����$�@��oW\���~�g?��# �~��e�B�b�̅#�NE����C�L��~R��P���a�(F0s=<�s�ȴ5��	�S���T߱bS�Γ?��,��l����](�B�9rY��@�C���S��:�\*���PU���@%`�\��"��"��	�e	E�K
Ur�E`�I�Ou��/D�M��x�t��!�E
Z++4\��$�1o�; �HAia��\qB9e �u{��}�Iz�+��^��������G,���?ёH>i��L4S�h8���k�q��X~R#@��-᠍/q풕�bB
-'5�g}Z9n���#��r���㉖1&��Qc��\x��z�⛋66b&jÐ0x& a��ߎ'���jg+1 "6	�o0&��ֽ<��py2�؈k,��HT�=�y8�՜1
�CC�'���J`%֠N�� Kޣy��0�g�+�b�h�<a�ˈyh��K:�<���|��w�R�����HӖ�뱆�'�0<��֮r�Va�2LO�q�.����ۂ�����b�@ƿ�<�p���y� �d|u=��W�d��:̔���W%hy&�'��(�/��X�mR��ۣ4�t"T�O���� %�$a��
SL	6(�I�uH��7� ���O�J���� b8q�@�5H��qHyT*���-�1s9���ŪYG�C�b9s�P�u�H�	X19�:��T5��Y��!Cx�|���p�h�O�X��	�q�p�s��J0Э�!Ǘ.V��HPw��x	c�A�~��h��܁��P9o�,�K>*�.1,���.Cet*6lY�$H9��PdȒ�y�-�%7����᠝�M��� E:Y�E1�`�S&ph�`�I�~��<"�G@4�f`9a
�O���'��ܩ�J�_X��J�ƿ{L��0�ڽz-��N��p��g�ŭ���WB�%�y��D�] <e�BFm&�\���A4�B�M O<Kw��Ș�M�5I����.��v�0�(��PDX�M�"l�O��$��#8�D�ƻ�` T��'/4N W͡,N  sÓQy�u
ؘ*�ds��@ ���Ow��$qB���pr�ăV�U�;�t�0�f^0c�:K��^(�^�G/�hOv�bW�N35���0��Ī-WP�%��̓ebQ�ۮ��CƎl*�k�N�>].�1��e5t��4S%@qCKF�094�(��7���2Q
T1w4dE���+b�TmҕB�o"���!L�o*.� RF��d���(;L�T�&��	&mDL��O�A���U��.?q/�*�.f��e�����4�!�$1���[��܃Laq����QC~�D�q6�X��T}r�6`��e�ѠB&�����߈��D��pN�]#�H�d�%��*TiLax��
��%�� &!�Ia&LUg\FI��*\�7$ �����C�m
Gm��K'�D;�
A�;&�[5�'���H����fn��͔�FB����O�e1�-�E�	���WI�Փ��\G�����MC�n��.Ġh(���i���xBaJ
F��\J�@�Ow�Q��-u���"��م$ U��G���D���鞜sj��!6�<Ս��n�`Id��lS�c�O<��X�h�QD �02��T��K��C��y��A����L�$�+p��	`D���'��K����wˎܘ7�ƽ� ��ÓL�����מ���"�_$��[H� 6�̥z����&�{A��U�`�L�K�|C�aR���<YA�3��0F�T2ig�$��XA~b���$Zލ�*ƓF����e.K��y"�ܺd�r)�'B�(д;�F�ʄ�Χl�<�ȓ�jM�5-��VJhѢ��M,�N]����&S��j�
��Ń2�Շ���<�6���S3�ܶ��ԉ� ��m`L�$%\c<Q7�̖?7������q�D��dfH�q�0D��M�.��sú�9�):Oڭ��+D%D���N� :D<�@��j�'vX (�2��cf�Q'r��A�u�����8D��!Y2��eZ�>� [6���y'H�D�;#�+x����v���D
p��(V����`�|�<�����n�`���CD�a���x�t,vS!�"�����Vq��O虚5�^lh0Q�B�ۃ`��A�����tÂ�O�<:��5��O�:mQ7��?Fhh*`�4�y&��65h�a����b��M�3��pԧy�K�R
8�RA��]8���)ڼ��~9�P�B�=%n�$?qHg�C�9-��N�B�P�LK1��`˧J�Vz���$/eJ���"�<*�c���O��zc"�/���ŷ'&H�NɈs�RA�'G\�h/���L˧x��sŪ��y�ݳN6YU�εv�*Uhe��$��	�+m"T���X�	.��y�a2�O�T8`CO?.aĩ�rfƚp�r�����>�ԣ�F�8*o�$�E�X=�%��tj�P{7k]"��L��5q�X!(m��Ze̓�J���Gi���{"�yӐ4�VNΈN,8� ��	�4G���'IbpȒO�$z�h�Kg�:Nh�C=O��o�2t0Z���%7�����W���ݴ;}0w�}�$�g�40Z�穠|��iw:�D��U���CE%{��rs�Si8�<���ݟ�pA�*v����dg]F�l��F(+S�D� S�Hv�cPŗ�(���
�HO2�c7�yH1��C��7�RE�0�D�;)"M�i�ihq��̶a�Mr��ԬW� r��;���&cr0Q�W=O��	�S�l0"%;Uԭ S�x��Z }X$ B�#�0�I ���t��҃Mt�剄���}�  w+�Q�����?�R"��f ��C IցEa����J\�E��Ծ2� �8� �sP���Ƀ6M��sCK�!�x�%��7E*<j��y�ρ��\ JЁ�����?���U�󮏳%�� �d�C�;�Ȅ1%�O)�9Y�Ny� ΄~ͤU�� ��Ń�
D��U@���x�M�5	C+��B�f]%$��Q��6Z� �����<8�
��y����|�&M�.s�p8�&����'p9�"��4c�	z��9O�VJUh^��@�Ɗ���B4k�D��f%�H	���(VZ����Z<Fi ��Hq�dޘpe���� P3>���J�lΫ6��SZ*�ʓy/�ɬ�<�R(Azl��0d�i*�o=���N1w�dTK���M����3�:�+⦌�*�@�RǓ3��`̓�9�T� �!�*HL�8:�a�KV�	�t+ 0��P>�����^�N+$@G�S)�H���㏹n��D��%\� �F�f� ����~�c��WJ�i�`+�,1@I�u�F|$󤬞�H6�Ē!n�y)���h��!Ēxm�y*���'��x(���$|�i���O�YPA��Z�j�ㆀ;��[��Ɋ>S,�$G��D4�uK�}���4"�X�p�o��t*�I�j@J'
>��Y�B���'�$ݹ��Kv
8�O"~�Jc��;Avt�ï�&�����i��x#��_����,ˡ9��xRf�/D�N�*@aL>kVI
��oeV�@ �����"i�d `��Rޟx�3�)� �P*v�]V�``�Y)r6DA��FEH<q���_h�ix�CЛj@�Y8��V�<i� nC�\+BD�0�nq��A�M�<�5'��v�Y�#(T�CVf=3GM�d�<�ao
}ۘ��r�Z/\f�`��h�D�<�BA�4hJ�����4<ۦ����}�<񓮇� �ʔJE��}�H@�Qo�<9�;]����p�9�pU���e�<���C��Yxq�Θf�}���j�<�r�Z�>���W<xz���� �g�<��@��Mh�C׫�5-�h���`�<�q�ˉ8�0���5BxH�!q^�<�g傗K�Lz��޲so��I5(X�<Y���(jc�pp����=��9�5�PU�<�R�v�y@֥%+�XI�O�<��	]���F`)%�tb��c�<ٖ�ˀA��y��[�v�V}���Ew�<��	
1�^��Q�J���0�
�s�<i�2a��ꗁӇZ�$�!s�<�� �
r�� ���Q��,�Q�Ap�<�&�u�l�!+��Zx=I!�Xk�<�A(��p?�A���H�� �Ae�<�&k��j����P�oA\�R�^�<9�I�(_�l�:d$�&;�
�ŝ]�<���&x��	�Pg�gk$BT	Xq�<y%cO?&U�ժ��x�Ybab�j�<qu�+��I��ޅ|��5�\e�<���Ӄ_���e��"eq���b�<q�S6!��	K�¿�qn`�<9�.ȞV�$�
>�����_�<�n܀ZJ8:ak�.z��MI �UZ�<��lT�c����Y�]Kz	Q�A�n�<A��7[���Ă.7�t	�'��P�<�g�Q�'N|�2UGS�2$T��d�R�<��B�>�㤩�&0��)j&,L�<)%�/#B��'o֢2T�Q��F�<Qgj�S=�����ŊEv�ق�B�<���\�:���2WjUA�j_�<$j�zk�@���\�MjHI�� b�<�g&��H�D�<Z���Ї�`�<q"Ś/f�E(�.V��X܈do\t�<�/��}Ψ�´ǎ<LN��Xp$�I�<�qɎIRz�C���8���0��H�<QS ���!�D �,����E�<�R�%&���҆�%h+���g��B�<� Ӭ��VK� z�nq�(�h�<i�B͟S�LUz4j��BXۗMj�<�!-ӻ:f��� A�����f�<��脾s,�He�ɧ-���vl�e�<A�Ί�C� h0��$�J�w�F�<���1uF��6�ߝm3�H1�o�w�<q!"���܍�tiqkxP�CH��<��AM](���J�S���Tdt�<�3%PPpF�{šDؖ&)���s�<���֍�������p�T��,�r�<��El�����><�]���p�<��v�b7��� ��q�
y4PC�I�dڈ�p�/	/Q�ܝQvd�>$�C�ɛ"�J�Yc��5{��9в��6!��G>p�l	��H�P��@ku��
e�!�ě�a�ȫ�@�/*��`3�ZT�!�d=TX�uh��pd��k��!��'KF�C�ʒ�yf��*-Ɔ��ȓq�T��Cm�YJt\��`�U*����S�? ��$i0�83�i��w��p�F"OT�A�K�9s&��+���Y�"ON �C�ϰ8, ܈�+���1�"O���'��t��|𒥌%�J�1`"O&���D!y:^a)%/�0�����"O2L㑁��7F�|��P2R*f�B"O$��٩7W��A���B�^���"Opy�`��g/�A�կY���A"On�h媃.w�T��D��rc��"Ob!�7@�^^T���i��x�8TA�"O��s!�"}Fұh�i�3��`"O�$���'`�ȵcb��_���r"Oڬ␇ַ0s�\c����z��8��"O����X�m�Mq��]�ت�"O0��)�:<M���(�b�s"O� 룍��(ơ�㉈�N`i�$"O�$���A�lV�akW���a:��'*Oh�;�`'�j�{B���,���'�����L�d���Ҷ	�|Q`�'O��"�*6ɪ]����:��
�'^n���1i6.\�@C8t��c
�'t�ݸ5˗9f�Y�f�C�*b0
�'5���S�UrB�Bu+����	�'���ZW)M��e�O/�2r	�'��8R"וk�V|�t�_V�r�':�k�@m��	�J-wbQ�"O����9I}hPegP6_N|`�"O�a���ևH���kί^X� "O���"���8���ӊ�)*�J���|��)DҠ'��]q"	��	B��C�Iu���X�.K�/R���4`
��C䉾:9<��셤e�XD	TC�;P�C�I?_���;�i�/qyp[E�s�\C��+u�~�)V�L'l��5�Gi�"'��C��,R�بS�69���s��H��C��/��5�9Zgd����د~�VC�I��n��f/K�2�NYH��'G�B�I;q�b鋔oWf��TI�� *�B�	�&>|�S@�*\����5��a��Oj�=�}Ҵ�[%`&np��O
@��*XY�<ّ��Wx�Ӭ��_;�(h���U�<��lHN�Z�H�:T8�SWF�T�<Q1O.c����K:O:�k��TO�<Q��*��<��!"&�$"��N�<�k%-��+�MΤ*���1�  F�<QS�[�k������+t���AlTB�<	�ȖcH�t��o�f6,��1(\F�<i��A�����'J�}.L�<�����=�G�*-Wza�㋟E�<��pB i�䥃D��AQ�SW�<)�,[�x�F|{r@�."�2@F�T�<�7i�G��a��O�&2	�r#M�<YcX�>N��+U#fT�eR�FH<��ǵGs�[p��?o8��U��1!�L�M��!
�g��d�E��O5@d!�S>�ʔ��:=�`�b�#C!�d�0`j(����$<��V�H!��
?j��C�i�!�h���*ռn6!�R4`�r��g���m�6%�S$��J�!�$���[�,� ��T*�c�U�!�D�������L��}�U��7!�dS50BН����_��	3�E3!�$����rb"�8*��dp%"�
�!򄘺eq�a�������[3 �!�� >�����Bp��E�#0zH"�"OԘ;�+՛:����ӫV0XJP�
�"OD������4�;��C�sܖ��"O��vN�5�J\��nل���� "O�5oV!}=Ɲ�r.�4��Y�g�'h�I;v
� 7�<j���#��:`B��,M��yz�'G2�΍��K8NG�C�I2����4�E>i�e9��_c B�I�A4Up�j�=]~�z�ğ�`����0?9��X�S��av	ʩ�^p��eTL�<YM��7ft9jw�Dp�eTJ�<v�̲:E�(
q+C�$k�n�IV���O8�y�Ȍ{�	�0�4Y���{
�'Ⲙ9�T"NQ.z�K�.|j��
�'��$�Egݱ@Uha�a(��	=���	�'�����B�jK�}\hE+�'v��W�u�@�0%��?oа����'T��rI�	O�f,)�Fޘmg��8�'Nj�c�j�(��8 ��b�:� �'z�̳�c��n]ҹ ��a��i�'j�"�U�~7�X���[x���'�|���
�5�r�H���i��]��'�JH�2AWA��y�@��b�����'�@]��ݑh�8���(���tp��'�R���b�0Ext�*���?6Q���'L��bD�Ih� Dj�5- ��'$�I8Gh��<S��u⋛b�r��'���/��'����ϽB�d��'D&i
�n�3��(b�߶&�VM�
�'�Zț���3[�Pɑ�I�%�����'ou�j�&+D�g���p"K\�<��Ǎ�40��"S�لL��eȂC�s�<�S�U!5�B�9!��FW�� �G[�<a���P���	%(U�<���QS�<Y�@��	5���%�RB{�<���!{��b�C�s��ʵ��b�<�R��|Lҝ�5L
# >�@�ZZ�<��!��Y���N a�%���m�<�Ӌ�W���#�@S�����-�j�<�4-��2�����-1��ȳS!�P�d3�O9��"�(6T2a(��-}� U�'Z�]�-���#�
ND�m)� � 5!�ē�=K�8�$G IԊ=����2.!�D�V��I�0M�d�z��ac�,#!���TL�Z�"H�\Y�X9����?!�� "�L��t��AG�i�훗M�!򄛬��-;IE�8�X�+R���S0!򄈖@�� �EK���0h�q�Z?H!�r���\���5��-�����'4�|[��F=0�+��F��08��'sF���'J�l�)�E�)EHP���'�~Eړ�F2�6���F� A!`L��'�`{t��yE�pS�bY:)��H�'�b�ɗl��G�
p�s�Zs�:��
�'�ވK5b_�A�^��u,�,i�2	��'bd�
 h�'�+��ēe�0K
�'������20n!�c��+~���	�'�N0�t&J)=t���B��:����'�88U
9t�xc恧8.v\��'�����	CZ1��M1NA+�'��Y����+�>E2ଡ଼�[�|�����X�L�, �f�P�Pe�k�!�!�dK�*�D��iɇk������:���Gy"�@r��5\{@�:�) .�6)��"D�� p��`�|��B���!:��z�"O��D#\�m�X�����F�(���"Ov�����}DtE�%�  *<"Ds�"O�A�'˧J�,@,�Y��!RT"O*A��e�,HF��k�dѐ�"OH<{�F�S=`\B�e�o�u2�"O�Q�t��#g�}��.��p��"O�냇P& O�<2$��< fy1"O�y@`L/������F&0��"O�A��GY�^c�A�\=(���"O��ի�.L[��a��*5S���F"O�l����'v"VxӇb��"(�"O�AC%ԇu,�t�O[m32��"O�\�pE��&�(��D�{H�M� "O�\��MWse��ѐn* �"O�T��jY�P2<|�m��	$�S�"O^���G�K>v��3��K��1�p"O�!��H�;V=pˁ�Z�2�[�"O|�i֢�7ٜe�����֔��"O�%#R �L� ��"/�%q���"O.���J�-Z�h���4Ih��"O�<a�N���36m[S	Α2�"Oֽ)�'##�D�{��S�O:�qE"OtYv(�5e�\�'oL�b�\��"O�8Q٤z1�s5�'4j�t"O~�H�Μ�s��@��U�4"O~U�2�ʜ;�^q�����^��#"Oj̠�Yr�0b�)ڎ��"O.��w��m��)��N!�ZuA�"Oht�-�\��9ڴ��%�>hا"Ot��3
�2�C0N�:���C"O:U��MO>�1`�BB/#�8���"O �5�Š#��CL	�f�N�9�"O|xp���HuS���r�.���"O,ar�$4C��a����i��WT�<�#c�-3�Aۦ`T#zrH�7�e�<Y����m騙�u����B�&��y�a��3��l�@�_B4�9�$H$�y�e��vŮ	�R� �0]�  t���yBjo}�5��lK�q�Ty�E���ybd��Z�|��HC���h�뇓�yRj�W��Q1)�4?��qy�H�9�y��E �J�h�L�ijФ�S�y�Ø�8�n4��q������K��yB'ܥ{p�Y�Ѡ��a~�!F��&�yr��*.*�"��	�X��9��
��y�D�_�T	�ҬMX�F18��y�j���slΈhZU�B�%�yb�DWv̛ %W�k2��)����yҮH�Z��l���.1��y�bB'�ybnK��]�3nݒ/��T٦	ѩ�yb�@~�<�'H� ?@y�Ȓ�y��R?J��HC��ܬ8�6�rt���y�WQ��()��5M�9A���,�y2�@.��8+�+�8B�`��3�=�y��0Zp�����q`�%�����yr*�X�~ ���Z�4H��`ܓ�y� _�p0P! D��]q�逹�y�ȝKp^My�ǅHpf)�g�Z�y�P;x��:#��9����I���y"��v+�%�DHþGό=��\��yO�G���ed@������4�yrm��a��[6�:6¾$����y��(y����'��SU����y
� ֘ڗ�М�`�ش� �(��"O�T�$�����u�S�^�hI�"O`(��B߉X��Mv�B �p���"OF����#�"Z	0H A��_�<q�ٗ1c�1 ��IPD�2���`�<�B$�,��HXd��;Rt2`o�c�<�ƮX" p��̧	*�)��b�<��拖#����9 �\`@�L]�<�'a��R�`@�[7CN��
S�<����W3��Qr�0SgH��TO�<a�gԂ3��@��#��A2# 	M�<ё'�L�|D�B�
f\H@���`�<a�M�zU��R���gYq�<!��F>:"�i���(
jT��/�n�<�bFG]=��/�0b<����T�<Ѷ��I��b���cw�8k�o�U�<��蔖x�L#Ɔ Hj"���)�l�<	Ă@
&�9;��ٌ1Ƹ�ϟr�<���UM���K����`]�J�k�<�� YH"���ٽ�(Y�Zi�<y��1E"�viG�����c�f�<�4K�c|�-#��՚g�hH�4c�<Aq��Ii� 2��>l�ډ�pE�[�<駤H)Hp8ySi�#UV�-�Ԇ�r�<ɲ�3\�����cW(k�b�[p��e�<�V�P�
rD��E�,>3���CLF�<1i �
���qъ�+7xۄ'Jg�<���� ��M1O�>�鵬�X�<Q�Ӎ`�|"�mʃ;2Rm�DB@`�<	bMO?6�J�P�ƿgg:�rgj�Z�<Ap����(Lb��6g4�%��~�<��#ݚSj�Q�rJK�pr$��1�P{�<!�S�X\~��C�K��P(z�̂N�<A���AF�H�abZ r@�^q�<1�*��l-�!��	CO����[n�<)�jP�P����Y��Ѝف��A�<���
<��0�w�ʜ �$@}�<��A�:h��9ՋY�U�\�$B|�<����� �D�B�^�J0��F�Py���%Xu8�:Fe�q|^ur�e��y�d��u�h��,ӉS�n%#��y��L5!�f��G�I��x	�GA5�yb؈��v��"u�� �ˏ,�y���7h9d�ȼmO@�1!���y(5pZ1����OLC#GV��y�A
���,i3F�`��Bo���y"���O�FL��K!Pqؑ��y�gH��b��a(���9�"#�&�y�HJc?0���]�qzHQ�\��yR�Ƌ4���9GO������ߪ�y��X�}4p$�j�0k&�#�o���y�C+֩q���%/~�MIs����y�
W�k(����ϯu9�i2�oʽ�y!F]z6a7��6 :�C(��ybd�:x�tJ�kP#*P9�����y��#AL�±-
�w�8��`D�y�b��e�,�*1�6f���K1�R��y��ݚn�Xw�>Z��(��yB'�-G�$�c����8
���y�J] F�l�#���
Cݜ$0��K��y2EH24�"�0��Q�H)8da���yB�&X;���5'��V$����T�yb�Pl��,9�kXLH&�y���yrK��o�pʒ��SѲ�v�_�y
� �*�,��"G6��G��Oł��`"O*����X����
\cZPW"O�9iEա*
�M	Q����x�<�耹(~ ���HQ'u�^I!�B~�<9�,R�6� g�U�d�P@�Ey�<Y!� 7a`A�3 ��h{6�%�^�<qf�ܻrz��O4U��ɷ"G@�<�ႌ�
�E` ݅d~�U�[{�<���H�y�b���<2�<��r�<�_/Z���A��'�y!n�B�<�՟[��<� \�����|�<�V��/> ا�ݷ[�8hdJDA�<9�f[	Ha��L������C�y�<'-G�C�ּ��-$B����}�<q5Α#�D�3�m�.r�lȐ��_�<�r��_�Z�c!��2�.@T��Y�<I���I�B��q䈿gM[��Y�<Y�cD0#,E�@J=7�.�r���}�<Q.о'���Ea�1�*�*3�T@�<�w�,x�|Ҕ��#8~4��|�<���480R��	�}�����y�<I7jG3 cnEC@��4��Z���s�<�"nY:L�ƨ��L��|l#��q�<1*�9H��MP����b��_n�<�Ϛ�S!�}j7n��?}��z�+�j�<���ǁO�PEY�H0$���uA�^�<Y���\4�Y3 �3I�Ƙy��F�<Y㩕y�,�	�ǅ\�"��@�<��=vzٺ����&� ��A�	w�<	������p��U撨�F��u�<��F��ѨMK���0y\i0�̈́l�<�f(�2�(,y�Q!s����%[l�<��2Pe�Q�­\���� f�<IaMP�r�n���B����(Kf�K�<QEJA�;������ܢKA"f�l�<���>vŊ��Q4 ϴ�b7�p�<��i�N�&��`BJ%v���E�c�<q��X�P��
�Ȅ3�,���o�^�<�ů����&BO�Z�4h'K�X�<ɲ���Nu�H�e�L�H�#2!T}�<QS&C.�&J5��Y����S�<A��a2$�d�IlH8�D�[�<y�@cI�<��>�d�1��JX�<�ѡÒw��=$L�\ t�qC�[W�<٥'ΕF�$0	�GM
D�IJfG�T�<����ߎ��d���l'D�4O�P�<	�Ɂm'H��"�
�h4z�
f�<�w��cZx��L�gcܨ�V�R_�<�P�Ӱ=���X���<|���uU]�<�1-��%%��уh˶LV�rj[U�<��K��5I�؄��9,�a"$i�H�<��%ݼs���H�,��hኍ"���E�<�G�O�"?�[�Ȅ�)��܁ao��<���� �>��\�ac[e�<��a��*�x�fػC4�% �_�<�t�K�>����ܲ��0�Š]�<�v@7:����'&!X؝�g[p�<�B@;�p�cn��$���䇝k�<W}, e�F�	�C0�Ph�<1Do�(Ì���U�3�!xE��m�<�� ;Q5,|㯊�>�~U�!MMR�<IP�	/6�м�1nPR�*�� ÑJ�<A�N�R��a0M�A��(ΗB�<	C�
�U�T#F��Ӷ��U�<�  ��ަ�l����+�V0Cf"O �gg\�b�<��`�%'8��p"O���%kE&1Y��WÇ����!�"OD�@�틃>m:��#�w��\��"O�y�Ɗ�n���!"�}��13"Ox���A���MZbA��qx��R�"OV��b<7$�H!" ���a��"O����H�� !��U�J��"O�(�����,TT ޠ4w2��6"O0��#�Ǭ'��}xu�Wk��"O4�*�[�
�x��M\1Qa0F"O:ujc����U����B^����"O��ٷ��n�0�`�ݭ>��1�c"O6�jU)W(�X���G�<8���hp"O�9�ăD-tl�4g�~|Ψ�Q"Ol�ydo��M�He
�#�����"OxWI�:�H�!�r�(��"O9(��^� a����6n*�8"O���hQzOف,V��r7"OL�;ŏPf�)X��V3I0���g"ON�9��Dz�����A͝��c"O��e�&3>��°�4!	����"O�)gK� d
�,C��3���Q"ObD0��1fz^�J�o��h��"O�Mrr��&C�Z�;��w�@�"�"O��a���Te���7�*#�@��`"Ov�;��G�6���p5.����"O���0�`��B�ML�"Oj8�rj�4z*�YA�bP�^�����"Oh��6�A3 �a��%RU�=� "O���@�vrfMȱb��3�l�4"O��%',���7!��W^�홐"O2���+c�2=R���{ft�"Ob����2W�� � DƘ��"O�q��◇K�y
�o��;�V�j�"OҨ�"��*j@�Ԋ�F=\|���t"O�l�d�ߐb �i0o�ǮLQD"O�YQ�
�u �+�p�l3�"O��1�O^l�y��_4��!�T"OF�H�k�*�25�,�@u�s"O"\A��-��,z�&��:�yb8Ǝd �GN��Ҁ$^�yҁP�Fa�I�)A�q����P��yB�M�Z
�*�+H�"�
����yb��fv.@s�
U�>���G/G5�yRCK�A�:��S�
#o�4];��ȓwa���r��Z����`�ѳ&��Ň�5\��_�6�$��Z�� �ȓsc��Yw�^�K��X�ǉ5!�
4�ȓ������=F �t(�� HF��ȓG��DI$֫\�tXw(ݓ�0�ȓ%��ꕄ�U�VP��U�z`bć�b80<�0�>bu��[���D����ȓ	yTQ��E��]�!ÕW�|��j9Td�V#�.I�{�����݆ȓ^<���ъ:�*mJ$�"rxe��bpT�t�UJM�d�;j��I�ȓv�4]�e��w^�D��7$�l)�ȓgnH�� N�xl
E��N^*U�����9�k
G��U$�|Rل�3}Z5�T"��g*�#C��w�b@�ȓF�@�C�ÍX�~pc���1n�݄�A ��%%޷-�|h�䣟�2 Ԅȓ�`1�6O�4zt�!�ǧER����S�? "dy��Ѐs�v� ˗$! ;�"O�T��'��h��)��2$PPr"OT��W��(N�,�lB�0�
 "OZI��(+b���+����K*0��"O��Qe�ˉ�����Q+j^��"O�ۖ���$�0�!ي:jR4��"O�5���W+d\����rR�:d"OfT�$���%<d\A��P�]�"Of��!^W���C(ك
Q�8�`"O��u.(����F�EV�1�"O��۱�LI�Ā���]�8>�T��"O D���Ҟ ��eQ�IO14@x�"O�m`G�Z%G�� ��73�UY�"O�!nFWsvd���8J02Q�C"O��:��ݽ6�^� �mD=&}�2"O��C��0�d0��JZ0j�5��"O ���	�19���@�гR>�b�"ON���'��2����H�)
!�dS
V�B=�����L�d�$t�!�P�c	�|�h���$K���!򤞷?a���)6�Nyz�J��!�$H>4Z����	6.d0D��!�D^��� ��J^;6��%�J/!�dX,=� M1�NU&( M���7 !�$�("���R	�b)�����|!��<p�H3����d<�5�5	�!�$�35�v=��B����h��.#*!�#��ŦT�~A��h�>�V�t"O͓���;#n�DQs-��Q��"O�0�R��+��B���%d�B�!�"O|)���Z"���qǔN��TBe"O�A��B���ʌ�� �~�bI�"O����h�G{�i�W�Д]��H$"OU�p٠W �Yb �"o�r�:�"O,IH���:�8am�!X��`3t"O|�
���>x��<)���a@^YZ&"O�r�Dɓ�>51��܀��05"O,�P��z�\��,��0]\�CP"OШ�n�9��3n�1&�R��"Of\zhE0d0��&��:8�8��"O�[�"I5Xċe���A0����"O΅�U�N����χ~*X9��"O���woC*r�6Ɗ,7�D��"OTe:����Z$� ;׈ʉ	�A��"O�R&�އ.� �a(��#(���"O�A��	\D��%s�	�w
�š2"O,���J�<��@�O�pũV"O��L*T��)��H�N���t"O��:�,�Q�l%� 쏛qVĔ��"O��2G+��[�H1�3kS�D@n�J�"Or�(E�12`5qvJ�X3�t� "O�\뵉Z_���I#{���a"O�9��)P��abj�2 ��s�"O�׏֪s`Jh�t.ė �X�Y�"O�4v�?,�p��e�$�P�i*O"��5j�%!�(
",�Yz�'#��9d���% �F˖�$I�'Ͱ�@��в'�
=  L�Hm��'e�\�0��]�j
� ɬ�z
�'� ���eѬ|��YSC%M!���	�'������rv��A���9%�@�'I@�nϓ!� `�R��.��h�'8�ш��3C ��6�U�x}
!��'JjH�t-�1b�iW����� h$r -I4'�(
�産*��}��"O����W<ws�	:�ŕ�V��"Oj�{Q�؄}�Z@�;[h����"O�|��Y'zm�է^MHF=s�"O*��
�}���s��I��y��"O�5�E�)�<��F,�� ��8�"Ot�� o( i���(l�E{�"OJ�b��ע3�Ɛ(�%[c����"O���MT$���C% p鎸qP"O�$:���e��A3�܈*���"O�9I�R.R��F�gu��9�"O��p��)rǠ����\M�XR"O����I,%��+��`e�=��"O�Y3�C�,�(5���9Z��"Ov�{�Q�R�:�k�"�*�
=@�"O��8�"P�,�(oO��]>H�B"Om[�Ò�i��@ փ8�m�D"O�a��
m��y�W���3�^��d"O�0s`f�R��XZ�ٙ �8(kp"O���Lɒ&�ɉ�L'��H"O���_	U��A�e�E=A9�"O����+>�MH`�&V,x�t"O�1�W��ND����ɩ�@T�v"O
��j��vόX���.��\��y�Dz�x	I�Dk�p�T�-�y���:}h$����?ؒP0#��yB�=v<&��6��/ٸ48b#�yr�ŋ=� y	B��/��걩
?�y2��K��;��߳f�J�Pv%R�y")��f�D e�z����y�B�Z�PԱ4o�-RQ��+���y"�)Du��%������jH��y�� Q�:9�3FU*Lϸq)u��y���H��(_�3�����y2č�>�j�_Z\ȴ�"ː�y�GUj�*%��E_�M1���d��yRI$S�2�!�؍O�nE�6��PyBΛ���PF�	vRR�a'�\�<�gH�e��݋��%�B<���|�<�"o��s��D�
'qt>y���o�<9�ٗCW�1��T!K�
=CT��O�<�T�Gf�GEՠ���V��_�<!��F���������B�l�Y�<y��?Ǝ���u�abei�R�<���V;:X�4*�i�*@�sD�<'燝U�����1frFp�r	@�<iW$�
2����#�J�z`:�(}�<�aLN�e�HE���D &�ER�fWu�<J�L����FB�.�0B�o�<�$�íf�*�r�ºA�����@Hi�<���[�$n�q����y�T���]f�<���*7�E��f��n�p�b�&�`�<9")�$	<0`I�ςtP���l�Z�<��F�3<��Is��=T��y�m�V�<	p��K�$%��
()	0�pE�R�<�`eM�!���2�%+��-�D�M�<���qd�u�&A�)6�IJ ��n�<E�^�H��}�,@%Si����Mr�<�q�$Q4f}x�)� Ɋ| GGr�<�G�ծ�Lcu�@ ��Ԁ�y�<��A(��3%
^Tg����+�|�<Qd�{]�(��G��y���@d�<	b�ؙh�kP�@� A�S�]�<q! /O�HPK!�,�qQJ]�<� �����D
Xe�s��tLҼ��"O��馆4E��0�1�P�b��i��"Ox���D(�l��ڭL���� "O��ȡ���	I�P��b��3��*�"O��B���9� ����M��]��"Ot�8�^�	��j�J�i�ĉ�"OҌul�l{ pM��*�jMh�"O((�EjV%D� Q �F;_�dqt"OVXd$�t���{��;��Q�d"OJ�0��6Q�X�d�w�ެ�C"O��&fۦW��h*��4|�|�[�"O��& �1�F�k2��#0�2�"O�X��Θ-�0��A��x\A�"O��i����XW��3�aD�B��Yʴ"Obu�WB��L���q�t��"OV��0��'"F��q�6Xl��Ku"O>�PB(�A�0�`b$g.bU�"OHuSBD3%�L:sޒ�Ś�"Oڜ�u-�?jc~(����`6-2D�0�2
�u��M��"֥W� A&i.D�h!ʳ.� ���oI4w_&��&�1D�dp啑>�4��r�9@	�P��$0D��V��aղ�3ׄI"�|Ċg�,D���q�H����UH�1�8-s#=D����
5
�:R&��Y'���:D���ul@%b�z��4�j�e
7D�|:�c����3M,�$ �2D���*m����.Qخ���/D��W��z���ZՃ�_�`	�G�.D�L�1g�2Vx�3a׻7r>�h$�'D��a�ؑ8�N�JpmV+����D'D� ��K�,A��|J%�S�x�>i9T�$D��BS+j�
Ur��R)[���j&�!D�`#�L�|�����>����!D�,(T`ڰ;�yW�Ut,���=D����I�es*��Vm 1�0��P�1D��ȗ�K)����C�v����q�-D�H���2�,���M�pڕ3w"*D�@���!C>��ƸD��MR!-$D�P�FAW����c�"�Vf����N,D�p���*]4)2��?mi|��L*D�����p�r��" R�M�*XB� ;D�H�@���xvN�B�Eʍ$��D�p�9D��T@Ɩu�l!�ƴ!�hyf�7D��x�
#*�q(�,_]VxiE6D��AC�	�lR��d �4t��4D�Lz�`���x���)D�2�p@)1D�4:�K,��h�e,.H{N�v@$D�dJp�W6r���p҇1�r��)"D�����E3!q�e��C�d�:@!��?D�@���2�Nt�5��X�R%)�j<D�Rs�
=/��l���,c����5D�,ɂ����5Y��9F24�k��1D�0�eG�0~�,���
8�Vt��+D�D�6�Ѿ�1�Q��6~cnx+&�.D�8	#��J�򱳦��Gފ���E7D�ذ��ȳ`��t@�Ҙ<@Z89��)D��rר�E���o�7fDP�06�#D��zDh��:E�a@�0
��I��6D��Rw�^�P����2)W�.+�M�5�6D�, ��#<�I[%l_47�\� ��*D�����,Dx��ް=��xjB�'D�<��/�50ݨ��F��,�����`&D� ���?,<H!�*~�ܪ��)D�� `��
;P��ꔌ�#M��r"O���q�%G����2K�76�Zd"OB T&��Qf�9���=z*�X��"OV�G�N��N$Y���2��s"O�QYӊՏ��@B�[-?�|�@5"O��I%�(<�0p���
CT�)�"O���eY�r������	�"3h@�#"O��	��&P01� �X��)b"O�h�/,\`�Aք@|�YC"O: ��E,W���0$�K�$��"O8�"�H22��irEY�W\��3"O����\�b.�U1"��"3����z�![�eHs�`��ôk�Y�ȓlV
9��U8g�V�1j95SH�� 4�l��*�$|���hf��*-ܜ@��XHx���P�P,��FX�ȓ8I�����M�x�Tx��H��W\<���,�r n2xI0��۲B%�]�ȓ!�,����؀v|�P�r���z�4ͅ�&���?���Wŝ�I����ȓ8�X�p QgdlC�@�$|@:��Cz	B��ζK�Ή���D���ȓ��})����2A{�݂2"����4�tsd��XU����3]���ȓ�p�i1+H;�0��  D`z��ȓ,ѤX3w!,eªQi�d�6R�h��̨Q�s��PoF��M�;F���8k��j�D,��X8d�NX�lE�ȓ	��1ѧ��o��Y���� ���ȓi@��Ĥ�D����#	�PS���� er�p���ͺIXpG٩u�RC剓Ci �ir��&n�M����J'�B��;U`xmY��e�Z�!S�Z�B�	t x$���;q��)�d.ϯX��B�Ʌr>6��	� �P���K�&ׄB�	�Z����Ġ�4��%I�Jx�B�	�]��kt�s!���*�~���%D���V	[�>�*���iP9y�B��".D��(6�؟y�]���3n���O,D�D(�� 6c� I�f�!����D+D���sH!J~ 4MK,v��ѠB)D�P�ᅂu�H�"�G�\�NZ$�;D�@�V�����1q�b.eu0��5�9D�|��B,-b69("��.,Y�07�5D��2��Pu�*�B�G�{���go&D�� 5
Y�I4��5W���0D�)�ɍ6�$�0����X�@�j)D��R�O850K$�L�ʶy(c�(D�T(�
�z��΄�z����Ш&D��)��%l��� �_�Ԑ���"D�(��O�:34hRr�T�����6D���`/�g�L��r�H۵�9D���U�J�V:��C�W�3)��0B�;D��!��eD����т48�	1�:D��� ��I8"�SĎ4:9��R�9D�,� ���zb���4�߀%��Yj4
4D�����Ps���9*��#p�8�T�-D�$�E(��iW��B�O�\G��cF�,D�tY!LVm���\+�:�sV�%D�p�`Uh���q�l��z���׫?D�x�b�5�|0�E0��U0%�<D�X�aR4��rs�lv�!3�#=D��2EHI)p�
P)�`Ď}�f�2Sj9D���RM�s���Y�(F�e�Z2@�2D�� *鰵��+���`B�<(�Ȩ�"O��S��F1C�e×3&�"#"O�`�4o�3B���I�.P�&�D!#"O. 9Q�K ��ͳp�ϡQ��{�"OZ��&�H�6�4��k��[
�P�G"O"� �3r`80�)L�6H!"O����\�w� 4�v�ƙO�1��"O�@��)Ҽ|�W�כ2�b"O��{�#8�>�c�i_y�|�Z�"O Qbf3���U	K�'�@�R"O��ɇc�0��=����{Ղ�X�"O��F��a�޽�Fg^!�Ђ"O�yY!��6Q�^�AF�*	��)�"Op�S���=v��mR�>I$|T�6"O�$;���P��):Qwh8@"O���%J�3��X�B��au�8ȅ"Oj�Y㇈�2D��i��R	��e*�"O�y���ѣ#�=r�?? ��"O�"�d�Z��d T0J�8��"Or� 1W ���8
�j�"O8��H�5Q~�pA�����k�"O��#�}ʥ��M�=,���u"O�(Ⰵ�)
���� O;�-
s"Or�֪�8�8�R��m	w"O�`��"ڿ�XQ��&�
�X�"O6}�w �;��κ<?�$��"O
�"��?\	�VŃ�C\�X#"O�M0�i_�1~�qR&%�v�R�"O�@C�F�M�M�"%�<mP�D8�"O��&_\H���T��H�"Oµ�FLЇ"x i@���*<��"O|�����4T?�� �+KcQ"O~Y�G�[-t��e��Ն5���g"O.�0�Ր]��Q�Ї�.e�d(�&"O�-�4-�n|�l*�	-B� 4e"OD��	���� ���P�r�[�"Oݑ� ��(,�ʐ"@�h�T8�b"O�pᥣ�6�HQڣ��}���F"O������b�
�[`̐v�Ш��"Oȥ`aK�������1?��"O
q����6E���y�C��x�F�R"Od�S"Jb�V��CT?����R"O�4I�1N�85B�b��mh�i�G"O��3A^�Z�LP���^�aT���@"O��bP�2`�Q��G�!;ju��"O��f�ha����f֧	�Qh"O��#��Z�.5zƧ�5|^ d��"O�la��D65����B�7LDy�"OF��k��diA�Ģ9�u@"O.؃�MV�N*ء�	<$���"O����E�0Y�~�p��O�/&У"O�a)�A�)|д2�Q\ȼ	�C"O�M1�j�6Y��L�+5��I{5"O,IZ0hȧHN�����1!��۳"O�U��	l��a+�� Z�r�s0"O��ŤN�'��1�U�>��QP�"O\� ���ݨ��X�g�8�$"O�(��׋�jh���S�f��`�"O$���+t� �G$f�l�S"O�q�ț#�f�2`"�$.h(li"O�9!d k�Xs W0!�����"O&4{���o�n�qT��0g~�P�"O��eǁ�4�P���g|ĭ��"O8caD�?F��T�5��5M�� 7"O� *��&j��`��T��M�=M��A�g"O�вs�X0h$���L�;Ό9�7"O�����}��8�cl�����"OV}�`C�b��Ċ�đ�o���z"O"!��.�/&���h��ڠ(�+��O�<9��ʬ�Iق�Ȼ+�����G�<��B�;w��ъ$슻j��}	V��]�<9U��(5V R��:4����E��\�<a���# p�3���Q(��Z�<��DL4��%`Įn�jyഀ�K�<)��r��4���̤O�	�FƋF�<)����hlI�$/C�z����Þ\�<��n(k�TI��(S�q\bEX��Gp�<y �Oc����$M�6�Y ��h�<��Ѷ �:h�gD�p~P�5��N�<qGf�<g F�A�X�:�`�X��L�<�`�� K��aDc�<( ��G�<	��A�mHa;�癣d��p@���C�<	4�@�Kh��D��~\��F�S�<�b��
�HаQMpu�牌L�<	2�^�'E8����)�ư��`�H�<i�'�A�v8�F�;���k�n{�<�E,��4���$&��%5, �"�y�<2�ȄQ-�bE`U�L�,��E�_]�<aSj��5�d�Ł�i]>�uG�q�<1'��� ��U��`1ፂB�<�p�_�K�BQ[֠�e�9��FG�<��B�%]Zd��C©D�ޅ �`�A�<Y3��p�����.[�MJ �,_��C�I���hSj\O�x����0.8�C�	5��J ��-pfY���7.�B�	2!��]:R�^��$��d�)2f�C�ɴy�v����%I���!)�7i!dC�	B+J���Ɣn�@�1�a-&C�I8"PaP.�#.X��$
=*�^B�	�j��1�"bڶjW���ʄR�XB䉯��U����X����]�DB�	��@���Br�((5O�,��C��*_�n�R��`� �����[ZB� gf2T@WKΐ[��T8�́�.�dC��9U�"��0#¼z���MA�h�C�3K��\��q�>���ޞ�$C�=�j�#��*�E���v~ZB�I������BRY����.dC*B䉰:�����O�U��х����.B��+�H�zs!а3.�5���)��C�	�$b�]����(\��袩��y_�C�ɛo����H�uv�s�@�++�.C�I�k.��0"�٤fw��c�靨/�B�.SiB��Ϸv�Ф��h<CA�B䉧!#� 8f�<IE��(���'E�B�	 ��@̀8w���T�R��B�	����'�K F �����jǚB��'<���Н,�0���IҾ'r�B�	�[��V���`u�1�΄lGVB�	3	|%����7P\�0C��<H�.B�I�j.�8g�-<�f5+ǌ#:��C�	Ur��c�2A@>q�'J�v�C�I+G�}�,��y�2٢�(]��C�ɾo�p��AK?X�0튅,�&"[ B�I5]�yТ��Q����! 'k�B�ɰZ'�� 
��d�xx1,R {�bB�I;�\1��	�M����am-K�>B�	�Ь�Bg��/l]��@w&ڗbw
B�)� �%hDL�20�l-�p�Y�*�R:1"Ox��6���D&]1�� �j	HE"O�q4���H��L��*R�3�(i�A"O2u�O"�drJ��]�22�"OfUy
�+4G�M��&�&HȆ��"O�t��j		+� Pa%Y*��͋"O�iq�!C�L,�rPE�
��R�"Or �'�^�<-KW%�2� S�"O�eYpi:��[F��^�څa�"O�l���� ;�uz��"Od=��B�oږ`r�
D#:WH��yr�^7$��iĕO��Ġ�eȬ�yR���Is�� � _�U��͖�y�ᅥP3>ТE�E�(%�-���V��yrT,�X�����7/DĀ�k�y��0.�@D��R&/N��$�$�y��D��"Qk�
�0��@jU%Q�y�K��h�z#	�'\���������y�k�2,�`�@:�l9x4Ş��y���e�T�∬q�x��>�y���7:2ht�ԥ�%e( �2��.D�da��Y6e�H� �I aE�9�R'D��)B�ǧX�F	KF,�,�h�PE�!D�P����MN@���ʄ5g�����F<D� �C�h�H����Q�
V�6D���#+�~��T��Č�j�1��4D��T�ȝe�j��A�Sc*�;t�3D���G�^_zd2�)]"X6�S�5D��!!��(_P��9x�y*�4D�4I��	8>̅�rm�~���J0D��K�#*�~�@���"�~x�%,D��*��r�~xp蝭$�F�O?D�(�c�N>T��gG��a�$��4�=D�ܢ`	KdAP�fC�3�Nd� �6D�<p��O�!���u�@�;��)�6D�tӴ�5~ĻF�Ea~b"+3D����;d.�ʃ\�l܀�"2D���B��7%\�xt�5*-!��*D�t
�K&	Ά%)B��9��H
��5D��9�a�'<ڐA�װP �AzF�(D��� Ϙ��|��b԰;��Q��4D�l���.Z�(0� �,$E�}�'2D��#�*ǽf�v���O��Z�K��:D�ȃe�(�	�L�n�4{�*#D�4*�➀B�J�c ��pa�U#!D��R!�D<}ך	�׏�� �DY�p
;D��:�k�1�D��d�X9�Py��4D��vH��D����X/Y�����3D��B�jĶ(,��GדJ��	���0D��閭� {�0	*�$<��$�,D�؃3��(�(q"D���I�l��&h%D�\��)V�`,9�@N$P�B2�8D�kFe��'�䉲�Qa`W�!�d4O�"g�U�Oe\(jV%�|�!�$�k���ؗI��X>��ʤ%!�D&'h� *W�4ѧE�;!��,���ۗ�/>�4x�DdV�i�!��mF��Ҏ�so��{עB�*�!��D�tY"V*��F�D���5�!򄐐
�v` ��),$$�D�8&�!�4)q�`2�ۗ� #�,�,W�!��w'���	��8y�]�!���N��QB�$�L0��߫v�!�d�;H��5	{L��@�.}Q!�� � �aK� ~�˶����b"O�����/1�EA0\�* @�"O0h��]�$�ʣ�VYd�Y�"O9��@�`�<���lF��Q"Ođ�&�ձ)� �J�'X$/���U"Ovq��E���a��C����x3"Oj,����B.꼺��ԏM��D �"O�(B4�Gܖ\!ϙ��p�ٱ"O�eK%��>1`��-��c*�2�"O4H���W'
�&��e�΃pp�Y�"Ox�r+�bn��GG�7�Fx	�"Ov$O��@Q�8��G �ܱ�`"O�"���c
0���J<�2"OƔ�Ʃ_�J}�#BZ�*�ً�"O�c7K�������ٗ^��1��"O0|�$��;���
%��VЮpha"O��qU'��Y�L�E�F�M��80"O�d���/6�����:6�*�� "O���п:��X��"�/8��P��"O�� ��^�d�	�̍_ ���"OQr���0���Ə(u��	�v"Oz��P�EJ�u�p�	VWPi��"O�bF�LP6��O���-B�"Or����$��tC�F�Z�)R"O1����<h���"�Q�A�PB�"O�l���(m�h���^9���C�"O��I&�����$2�߽��X9�"Ol!�U*$�@�aռ4�.��"O
|#j=<� JC��I��ɧ"O����%�)Q̸Qr� ;sU��QR"O|U�gͺC<\Y�dO�p���@""O��y�"��-`��x�G�3;(�(�"O���3�¼���I���(RC4H�'"O M g��3>3�b�.ٷ�.�k#"O���  R�E��<�G�Y'8�^�%"OhL����]� -�q��2�|�"O�����w�h��#ޒk�,�(T"O^���;=rc�1���c�"Oԣc�yI��S� ���P��՚�y�
W�D�|b�狞t�T,s�BJ'�y�E(2� ����t9x0u�X��y��
D:ܜ�
Qh���4�<�y�˒�v8Yʷ��Vy�1z�c��y2F�yjX#@��cȖ	��L��y��U��*��-λr�(ɘbO	�y�늴AJ��b����	S͌��y�C96H��e��2zP:�92O�y�����A�r��%	�y7@֬�ya�
�]� _�G�4&h��yr��8s�.�	���CF<�(�,��y� �� g�-�R��<!
}@�mA'�yB�U�o�P�@!�0��h��C�
�yr��3x���� 3-����t�W��y��	�$/r�2!h�+2����V��y���:v�� �`��$��i�����y�o����C ��:!@kd�ԑ�yB,�,�x�teH�zn�S���yB�9�ZA���:��Urc�%�y��<�ލI�F�S���Р�"�y��T�M�ir eJ/���G����y2�\�{�.M���ǰ
~�Ё�	�y,5�F�aլ?z h�I�C�y��EC�N	y�c���E�ЀƑ�y�&Ȣp�X��S�[�*,Y���y
� �ѫ#�5A��
���.`Eh�"ǪA����3B�(#-]k�Y��"Oh�����u��H%���!Ӯp81"O*��b��쵠��J�P�"Oތ�7�7fP��̉6�\�!q"O���`�µP��Aq���-/N�Y@"OE��ʷM���ˑ�G�8��E
7"Oإ��Bܮt��(#�ޑ�"O�x)�IJ;ș�a���8�5"O�D{��pJ��a�*O��,+1"OT��"ƕ�`f�t��b@#*M��"O��Vf6B��-
d�.���"O��QsiY�xخd0�d��T�ڃ"O�Ś`Ɔ�9�aJu��8@ `�"O���f�ݛ�#P�&��(�"O�2E�M�4�d� �OW(d"O�,����k�(�K���H��H&"O|=��-ه[��Ap���z�>`�"Oܔ�$��bmtiG	ɸ�M`u"O���W�J�Ѹ �Ùa�Ʌ"OT �B�>���(L�)��Y�"O\dv�Q�<&�b�_v�X+w"O$����rϜ���gY�.��W"O���(�C�p´$�8-����G"O|�r�#�3s�鱀$�%r���S�"O��ͥ;.$�K��P<w�Z�#�"O���@�$D���!�J�U��3"O�t+dG��� ����EtDj�"O�T�P��`Dj�0�$x���q�"O�h:�(�1o�.p!f*�#D��$�w"O.����73널��OȻ�F��q"OXmxE�Z!oO��³�9�lyҖ"Oʤ�$k��e#���!zf���"O���4�.J�� �c��<M�T�"O�D9t�ʪ:d�!��("�Z6"O�11ǎI�ix�p.��a� �"O2���O�8d�
���rpx�"O@M�&���{�D9�,��$��pH6"O�x+'�ɵrQ�@B�D6N�D	A�"O�ykW���n��R�S(zƾ|��"O�M��#u�����,w�<Q"O�p��'��-�9*���"�"O0�1AÚ��i�* 3-@��r"O�D*W&��!
�	@ɝ�pw��ۅ"O�(�6�IXdY�g��\��!"OA[$ ٘��ԣ��N�E�h4h5"O�i�F����3w*�s�h(3�"O�����E�<�E����L��*"Oҩs��� S� z��I��z b"O֝k�,]�H�����,�7�PЉ"OވЕ�!t8�)���ȗK����"OX��`K�i���r��y��t�"O�|"�C<'0�<�d�V<Q�Ne�"O`q�r�
 ���q��@��B"O��r�cԚ
J���\�4b]�"O�5+�,F�<����hS�H��"O�����.FR�I� �o�ޕ��"O��3�i�d����@n�C�2 2�"O꓃M��R���E���"O��YG 	
;�`{楝�Z�0"O���P�m:DX�7P��  S"O��B��Q�'CB>g�@�s"O��H"��	{R@#@TF��"Op��ѠʭZ[�툥/O���H�"O� X��@����$���/0,�	�V"O�p�UG�!y���6�Xh"Ot-��]�%��Q��
�u\���"O��8�c��?J��)D��*��1�$"Ot��b�_�x��@B��A�a "O*�Y�K	��,a�T�3�U(�"Ox�� #9!����{Vnm��"OX;�*gрj,�F`dZ2"OĉHB뇔$SjI�H�O�����"O��b��RY�*�5E��/�LY�"Op�"���d���p3�T2�nȚC"OT�R���e�*D"���(*�*E"O�'$�w���C(W켌"6"Oz��r����@bT�Y�b�A�"O�����CQ��h�)D��1�"OlLy�AܷfV�(37!�<B�"x��"Ol��0
U�u��O]a�0���"O���R���B��1� ƃ]�N�"O��i�-2�� �m��<1��"O������&nɌ`����-k�XE	�"O��9�KI�"dġ�)��A�9b"O@rPh����!�ʥDuF��"Oz�i��]�3�,����ԐOw��0 "O*����ѬP|����!eؐ�V"O6���K[%Kvt�Fn��z|�k0"O��9EΕ�,xpal[���q"O�Y�s���0��8�FB˭	��r"O��H�� $:�H�(U�Eq.�)"�"O����d��P� ��1,3( zQ���s���	�[>�ɢ��'��)�q�J�-�O�<
 ��8! �P �&���"Od���5z����s�)��9rO��d�l�C� �"{&�P�KT�,�!� 4z8T`��5 Y�vҫ	�8݆�U�ʽJ�T������M�މ�ȓa�P�&"^�I(��Ă�Ŗ�ȓ�@��@����B���-1���'��5�$���~$���_���a������	�Z�X#K(6 j�	Cnŵt��B�	%ST�sУÈJiXA�֪H~C䉢* Qr)N2�B�����29��(*	�',H-�QhY�ž���$Յ{�eX
�'��!�l׼Q�p���O�0r�ΐc	�'�p�ӈ�%Ai,mY0� �5]a	�'f�Ye.�q ��w$�"v�I��'n�P�ug�2)�]FM�u���C�'b���=m��6_��p���O2˓�~��$F�T�y�d��ԁA#9����3�ɩ�y�o�?+�ܭ��U4s���N]>��'��' >ի��5�=K��1a��� *LOH�'L�$�O�:�B�� �qw^$i��84��܄㉼XN
�X��A�ZIڴbi͢yW2�>���Iب`���X Kэ^RZИF�+!�䝤-�nd;�I5q���1%�<6��$.}��>%>O ��&������f��9G���'1�	7f���2��&���P�����6mw�y	�������>r(�ug��{�����@�S��`��W��|�DcF�%w����*� �Q�t��P�ȷSl`+��������d��x1���Ҕ=�����!�$O�|3����&β���R�!�d��O.��B���ɂ��y!�R�e@��x�&��z��J��<j!�d�+g=���%�K��5qg��"gi!�� ��e�H�{r1�a�9!d4�"O�qAC���7*���Wc7��Y�"OF�!��H�q�a���0I4��"O�HP��P�g���7��@A2� �"O\a@�c�cD9s���zEh��"O�qh�nI��,�y�ދy9\Zw"O ��!B�*�����/v�@"O^(�w�$k��ě�i�J��1O
�=E��cæN � :�&_3K��SѪ���y,N�,1Ԭ1ը^�+.NuA ���yJ��S��!��E���H�g��>�<���D�1Att����&J��1�f���Kb!�ߦ2�>�CZ9��Y ��_��|��i����gG��s~0 �%C�V!X��I��X�Iܟ,�E^	1z&����ӥ#���s� '����{B�)�	g����CI5���k4c�7>�!�d���#�I0�֝�"G-R�!򤖨7E -�D��(�LDsfB.N�!�سa�bu�*�.�ZQOU�!��_X�� ���{�"t�B��\�!�@1 ��S��E�;�@��O�$;G!��	3�R���EƝ�ԉ���TB�I����;LO���C�S�z��lح8�PiV"Or��Dœ���-��-E�"�R3"O �C^	�(�ċK�M�� K�D����Ӛq������8^�["�ݰ4�>B䉴j��!*��l+�МV�B�I rtI��N����r!�J:��c��D{J|JG��q	2�*b��#H@i1rc8�~��'�FM�0+�u	�l�b��$����'	 	J҈ϗ5��UkR�Jjbz�'Wb&O�qY2)����&T���͋�֘'$r�$!��B(]0��#I�1$L��K#�!���{'��cc�0w�qz��΃�!��R]������hj U���˓X�!�������Cmצ\|ZE2E�ݝLC�J�����7te�1D�B��vB�ɡ'� � �H��_-?�:B�	�B;$��!�@�p�ȄB��G�H?b�d���`����UCN8V�8��Eۚx��C�I=uB%8��|l�d��V<ܪC�I3i@�E�Ւx�v�F� h��C�k>쨨Dd_#|yv0�ᑲ9�C䉀 �H2��L�x!R��M�)�ƨ�`�)��<їd��p4���#��xSh�	�H�y�<Y�N<�ht"ga�P�AB�s~��'N]��?-�̭�ҀѪOJ4I�'��,+eA��Jd�P�)��X\�	�'�ṭ�U�V���;AΘ~�f̫듸�=>=Z4�N$$�2(("+�%�C�ɩob|h[�)E(a� t�&E>�|C�	9Fv���L<U�q�V��C�>������B�==Pp{���?gZ؄F{���ʓ�~"�'�v�hN�iNp�@Ϟ]�Ε�rO�ubr��uy�!��j��,���
���;�S�Iٖ/�8����fn�-JъE�a~�^�(��B5W!L��� xO�� �1ғ�p<�!�ۺ.�|<q�ʙB���6	�U�<����*Q�I��ᙙ (UCW�B˦Yz�,�(�����3NcX���
�46�����'��)F��-3J��#j_�YŮX`�	5$�T�uCC�2�j�T/ǔb��¤�.�R�R�񄇓��@bE�O�})q�lɊ0j!��]�Bk0q��
�9�^��Q+"p!�� �`� 3k҄��G_�����"O�|P׋٫B����c%\'io��;'"O���)9r�#��D5?n��{�Z����T�'�Xq2Ԍ5*��$��18h���'T�l;�d]�`f��ZE�W&.^�y�O��=E�TnM�G+t��$[��0�!����'�~ ���������Y�O�3S���+B���y��Or�"~b�(R�	ì)K�m���!0t�WG�<�d���8���an��;���F��<�ϓ� �p�U�^���*йNO����	�<��(y̜#F�ӥ'�r�BT鐰��x"�־f�q�B@�BtBkt͍���On���iԘ	��С�cI�N��Qy��ܟT�1Oh�=�O����A���A�*?�j��E^��!��b� t9���^�m�C&��2�!��"L˞|�#��5wP��Ґ���(�� Y�8*7�1o$���W(��il��'���iy|�^��C"�:}����Dk�);�L,D�L�m�7pexE�E��>t+��)D�ܚw爢 %���!i24d;%�3D��Y�JL;g�uhq�ug|�F��<��5�ڤi����4i!�;Nz���s�'�����H
�j��As�#�����'/v`��*+Ql���e/����'�����G����D�)d��'h���E��6�ͪW@ۆ%@�š�"O���fμn]fq�Aώ1P�d��"O�ԙ���D����2-c$1J�"O��H"���WY�/]�:sz ��"O��*E�<g{��I��ӿnm�b%"Op�Ǜ�XP��u��2rT�@��"OB�hMU
����J˕e_(U��"O��³�
�c��,xf(R�Ub3�"OF-�H:h�8)�@�L?8Ha�"O��ŏʰ#�dŚ�B��1�,��3"O� +�c:]�� 5]�"��\��"O(<i4�F��f@��@�V�<pc"O�ZA�-`��d*IfSjԺE"O,����5�L!W���Z8 �!�d�D0t�Y�D�hp���W<)�!�[�q(R��C��'Hc����#C�!��w�p��)I�7��I� _�w�!��_4n�l� `\�p��Tk��c�!��ٓ0n���焠K���D�7*�!�D�g�(�F �"6i4��gfܶP!�$Jx@t�� O5\b@���J�!k!�$ tm����(^� �<1q��?Oj!�䇴G'�u�$LR�i�B*a�Cy!�D�
�pLR���@�$�+��ξdv!���7Cr��Zv�R�#���8���8Y!�$^�+��1�F��e�`1��"�:�!��j��𡋊�Sj�`3q'C�>7!�$��(���M�m?H�2Q�Q0{ !�Εs).5��&F�I&�J�k_�q�!��͚1V��_�};�h;��1D�!�D�iȼ$�)ׅ$
��QkE%F�!�ִ ��d�򏋫V�nP�֧ø!�!�U�6�ŠCY)_�u�'�%�!�B=�Zm!χ�O������fy!�DB�#�0��qI�>�������J^!��0� ��]�	�s��AE!��L�\d�hj���X�Dd��.�fP�X��H%Qa~2��
�ׇ,���z�E��y��Da����CN�&�֌Z�� �y
� �m�fjԻ[�H�6i֒3�*�z�"O�E2%,H,z�d�x�q�F���"O �4Ԣ{������V)�.e�"O�kBi[Kh���.[>W^� �7"Onq�D	5�`�0s̀<P6�M�"OZ��b�.v1�� ��E�j��3�"O
����Y�?�\̓U�vVL%Y#"O�[��%ԦγmLF}�Ԉ0D������<�#� �r��a/D�D�e%Ә*��p��ř��y �%1D�����f�D�w�V�>ﶉ��.D��+�a1:�!�"�U�X�U�6N-D�D�o�7hp��Ff�
\ق)ؔ�+T�H:��\X_ư��m�x��Q��"O���+�ТB؜�B�[�"O�ȈQ&�����ЛIW��B"O��R���|C^��տY@.}1�"O��9'�&o~ BtfߛGjl��"Olu@R
�V���(������V��^��y#�'	��zCh�ZN5X��D)`�bq��@��6�D��	�F�rv�ә=��b7%Q?�Rlp��ˡ��	����O���)g�;(���'�蝈������Yg/W����"��~�L��gbʐF"T�Ū?��$�a	��^It╠\�"�J�����`@oՐE&�	h�'/�D��	E�e�h�)&��	�qF{҉K$�>yZa�*i���;f��ɄB�x�ʗcجXc���k\�B$d��}8�Dإ_��� ��L>1���;�J!PR��!	�pQRP[���h�c�O��Da,N�@s��(�\�XWAQ%G�P,����:=,�P��	'u2�� z�����Yb�ȁ�	�w��Ș��4�t	c1WܔDPw)L��y#h�|±M�v����!@�4�n);�Q���"6\�z$
�jR*R-lO����)I��!��@�.�h(pG[�	�t�t��K���A��� {��p� &J��%�$i1h���Ol�D�>�TBO"'��u�P1j�L��`�P;!�2-bR��A�	; �81"���_>5��hս��+bHS�?���A��v�1���b�Rx��%��o�iР Gߟ49�Ʌ�oQH�ӄp�)��Ǔb��e|� ��e��n{bK�%0��Y�ǌ�zV�4�񡇳#��% �CYa{�,������0iŌ����q����0�B�)�S�b��-�<�t2A�ï���D�bH���$Iż5�*Ih���}����cS�&�N��/��T-��o]J9"y��)��mD �l�//�8Y� �F� A�����Y����B��e?�N*sJ�w���49��i�:XS6Y`l��	!�pGH�[��`���^1̀�����s�t����ʔ_�1���(�0'�G���TϘ�eGBLсJ�?.��$���F�(|��)�����ҩ�Ry҅�&7Sp�zS'@b�@��$XdhR��OPv�F��)�Ш������%�oN��b! �XS���,Pt �DK��1B`�4���w�p$�E�2wք�ۇ�¸I|�ثQnBW&+�->x4�����z4�e�2vԀ�ӗ��Ky�̃��C�`T�5)Ȓ�2) �1SpHu���F�[��Qp��%~9s��ն[�l�dɑ�*p�bV1Rq哴6�`4R�kL;o�$%�5�Q�6h`y3Ǣv�ʠ��k ]= 3f55�n(n�v�t}"4�¢ l�Ъ��݌JD�)�"��e�V�����;L����ٳ. �
��x�acՌKE�s�Hh��D�Q;>5,֎�|����2 y�F/�3o&|� x�0$@�4m����"���L�wk3#i��I2l't�x�˗�L\6�U�A!+�Ji;%߁.f5�%8R`�'�T��D�K�Z�9�H�-WМe�' ��d�a��1tF��T�U�"��p�e��
& ;��^NHFQy��J5\\x�1�C�rK��$��ֺ�bM�O| �p֋M&��dC�L�@CSE/�Ms���%1�`���Țmc�L�u!P-�Pzɇ�?����KX�:aaH�0�ʐ�ei�0=)�X%G59�k���]�R��B\T]jx�SA�����U2;"�%u�����T�QNc��Qd��85Т/ |i�d�GsT: � -�8��G�Hh��	��@$  �����~
U�d*"o"v�yqE��R�p�	�6��=�B�OVQjp߂U�� 3J�b��O��8s��lH����>���`���`:p\h�`U� �.����[� |�:�#G�d
B�1�
B?���X Ǜ#e6f|8@���tl��
���W�<_y8�k���L�z��0���&b9�A� ͜�!����I_)�P2 L�!�8P뷏]�4�*fĔ Ŕ�92+ô~�ҝ+��Q/gKV�Y���$�"`�Ϝ�:�z�'A�̓D�֔�8	���+f���1D&�>A�)�wrR%�'� 0
�Q��+��R���0ׇ�2fu�4B# �榱��E
��Ի��&Afi��!�{�F���h˾��Pr� �6\ �-���iуZ�vu�'v��P��XH^(uKC*�+jxx�A�@[�ɜ=�4%S�2�R�¶�W�r��a,X�LT<Y�j�)mvd�)W�ۍ1��ec���"~�V�j�-F�L׌�)K>a�m� MԊ�9c);ғK۶%�����T���2sC_6*���4Ȍ�+���*39�u��k�+I���P�HV����^�,�����荂,�|� k���Ũ��� ��q!IF����E~��<1�q�N	L8,p��M��Z솔2AU�D?^�KY&�u&��qCN���j��+Ƶp�Đ XaH�"G�(
�<8B<�\<
 �PbL��Pb�g���(˵�߇T�0ii�	C$��ǲ]��] �%]f�Fm�C��u:����&N\�qHF씧8A Xx' �	��y�nѭN�ı�&�4i�0���) ��M��)T:s���Ɇm�3<	u("Z�P�s7��hтiS!��Q��%��)�V�4�0�R��ޑ& �E�!�� >�j�"����c;�DU�Ҏ��	��9*��\�"?���nՄ-�:���J]�#���)�c̼ �TIВ>�!�D�U���b |I��Z �'K��zp�5��أ�D�0/��2�a�3x0�EK�?�N���	�-�&aj1._�B��7�(�2">	��ڥN(��/Z�F���X(~�6�b-����!*�&E�^
�R�j��[�����O��������Or���A�v�b��@'-8^� �'A���ԫ|<e���ǹ8bpA1��N9N��|���)������@'u�$HZ�G9?:��'��A��n��Ϙ'8�5a�̑xm���Ø�,m#փ�5����J-Cz4��!j����A<��1�i�tHK�"��yqB���+�����Pg`C;E��G�D�>��{B�yq�IA�n���t�L$�Bq(���W�
� `�6"�*|y�T� 
�Uq��P���2[��3�u��X�ZH(�(�.R�W���E1��On-��B�L=N��#�U��Qq����Du�K�S�"��cI#0���1��P似E
��8��$:�n?1�eE�Q�D��Q����	�I�����G�>�t��N'��D��:T�	0�|}.ٻ$� &B�H�qC[<ܑGǓ?ND" �% ��I��F�?Y�8�5_���I��'mP���Eȡ_i��:Ȝ� ���̚��$Q<\01V�"y����m_.\�eJ��f�������ٲ��إS9V$�̣z���XA�^�]�����8(68A��t�~�@�ܺ*j:$���C�0=�SΝ1��X���BN�Yr"I��M��Np��xd$\� -�L�H�{���(WI��AH��];0n����0�]B���3H�;Wjl�熊��'hd�3���	� ���Idb\(9����	Z!B�zr�Ũ4N�0F��.A~�J-�N�r��_�e;JȲ��cR�����M�������h/�l"ٴ����*�ViI!��,^F��̌6M��FA�D@/ZHl=�o��8��*0jTK�.3��ܣG�I
LG��!����/�r�cQ"$���Ȅ�YA*8��G</t%)"/ڈHO��L>!2oZ�IL����fL/v�ů� H�j�t���f����Z�T�Z0����N��� �M,q�9CE��I�z)��a�)c�([����Or0�M�2#�m���W�b���D'����ɯa�aE	�D4�uh6���L�x�*&��p��EA�'c�*١Qb�
��4m���&�T��83H��aT�"���S�*�N�뮎��x8%�H�p�\�Rդ_�mnB��d/�X�rl���dӘ��m	1�����V�I�t���
	>2�Иx3�_^?�G��-QE���#ޖ �<�����(AGXXz��ȻX2�EYp	�ڄ2$d�����C�*MpB�T����4B^�?hQ�
�5е ~qR�P����%ȕ ���M��n�E12!a0��Q#c�9{�2�ґD�!���;e(@�R��&�!#f6M�tn\�V���4|a�t$'*�ĝ��*0?��hA�Œ�w�L��!��!@���M$Ru��C�����m�������T
%G	�S����A��"tѠ�ͧT~��k�-M�
�-!���+D
�ig�
&6���������}�b�0?	�CÚ$)N����#6��d�d���s7.�!��Ը+nVWi,d�b�L%5D��bݖ0�\q�f"W�+i�\Js�K�[.�AY�Եi-�&�'1N�0���|�(������a���#j����k�2"�yp�J� ���J?�	��ә��A´�N#k����S�i=.h�v���dU��a����wa4��Ї�38EF��ቘ4=3|AwƓ���'c���@(Op��`���§�!��@`#�5tnDy �f��/{@�h2ឌ;|+O��H�䂼|<�v���N�7a��n$������h3B<��lD�{�xR��p���`�G�JŢR*H1|Xup�Ñ9��88q�U�/�� ���4H<�۴! �µeU `〉 ��%yRMY@���@" s=j�ґ�Ĩ��u ��6E�a�!�F�n�c�UA��d�\8"� �/@��۳��HA
p1K^  �2��8=<<٤����`�?���CLH%�'�>L�qߠG�@ �</3��p���O�%�䏶p쳲C^��,d�Yvyx"�ڀ��t��@6��r��9e��׈VgzT:���*���F��j3r�`e�ǥB�����	(��@�e����-肇^\��ի�"ۊ"T|0�(r�Y��X�+��P�eF0��	�g~���Ҁ">��� �¤�.Ų %G�e��|2������I�lX��Ӭ��xx�#�-[�7m�����88ʸQ�GG�Ш9Q��O�o]����%|q�kqm4h��8"������ҔF�|-R�٫0ܬ�0B��oܓnTb	'&�l��$Jd+�U�J���EG�qbv�i�Ӕ(V�ِ���F�:�ATF[�w�<A�r%�XUit��O��a�O�҈��b��,2����;tBR�~6d�����	�@��M:�Oƍǖ�s"�=G�-,01���`�
�9�-�!v�֝ɺ�u�H ���8T��78Lu%YЀ$)��M�AR�����R��@�U��|2t�ʘ
22X05k���!ci�KϺ���n�Y�"P4����D�ʣ)^�-ѶN@�5'�9CI������ؓo�yS�1�襉�gT�d�wT�Th��ۚk}�xů֡|�p��E�Bٶ����!�	!l��X�� T0��m��IߛT��d)`FҊx�Zy�-�$O��)��� b(���ʔ6��}�ԩ_�Q��XA���~�&��A898�����e����a�b��#��D{r�&gG�tc�&'n��Ĉ�ܞ1� d@�U�QL(���+R=Fl��Ysȃ#�L�iE�SN�0�3d�~�Vʏ+#��|�ٟ�*�A���8YP�R=$�����P�IS8(��d�Z�T`ܺ1,qh��@e�+I9�!�'|`����ø+X�p �ō)�|a��[-t&��R�XАr�m������/J*(�"���m���!� ���`F9 G �8���gOS/T0�qQ��uh�[��	�|�&զ��0��G��u�Kן2=���U�_�GXu�@冏K�n�a	^�����Yx���KV�hO2d ���o��U����%z�X�Ă�g����7-��a`�F�BF8pXF�l��]���݅ r�a�R��ۆy��_�<�V/�!��"�&C6�d#>9�D�E�䙨CDS�S!��P�Զ�x�8E惈K~���Ό|TMa��Vl"��$[�����O�D�Rc!��?���h7F�?��YC��ܓՖ�����n;��CG�|��A�o9��k�ܴn�1�0m�>�p�&[�<q�FN"�=X�(�2����B�c���yRoрQ��� �.�,�H��Ξ!�)HՈ3ɸ���胏g���m�-	����C�x��ؠ�O�E����� ϩ;��W��	���,�.�Q��}�������F�⥉2���D��LзCB9gͼ!�g��ul�oZ��b``g�5A�� {g.L�w���� ��� t�q!�I�dCZX��m�P��}RA�[�����I�9Ԓ�x,ݧ~�u)O�|k�c����b3� .���)v�P�6���4E����X��O�b�b<H�#G3Ƞe�UHT�-�0vͅ��Mj4�L�@���a�1�X��a�$@���c$� >J�=�Q=��yrtO�<@��t�2�V��1�AU.s�@�5 T%�'#O���� �� �8�P�#pdԃH�6������!��t���GcB8t�������ysT���.�#{=4�;��xa駇*�(<���C;q���ࠖ{v^���N��y8��ۄCp�$��+%'����Đ5ڪa����L�V�Z��:DaP�M�HPʄ�D)!+�͠��1ӸA�j�Z�1�%�=6�)X�K�/��͛e�͑2ZV��1�� A����"*��[�b�Ġr�?_���w�ȾW�P!Q�������ޏyG��{��#u �k���(������I=P�H	2��?����x�� �Rɚ?ҙ�vJ�3���0/����p󤍰.��ɋ���
o��]�࣏=�����-�K���P�J��n��E��К ΋�1���`���|��q����<+��U�V��G�OjM�W�!/i,�<�`;r���P&��ɚ
����C��+@�?���pd��xF�P�1,ȇclT��3��@n��lܵ7������ײk��L�57�V`��R{x%(OQ>�ᰲ�(z�E�kK�y�#űN�D01� sRxݺ��Y�c5L<�����t(	B��,iN�%1vC�2H�n��g�ƅ{����j=hZA�A�]BpqN��
\)��"���'����J1g��R��S5��IXtaJ.T���|J��nځ@��
%�R��4��/���(��r�IH�{Ϯ!��*B+"��ePᬐ���'(�
uRd��q0�ԆSM����y�y���	�1���@1.Xn s���Lq�CZ�)�8�F3E?xE��^0*�V� Ë�HR�|�iؼ�y2�1��)��E����7n�1(�R���IW�\A`�?x��%���D.Jl`���z �GD�j���PĂ$�O:��֠�-t�7���s�4������i
�t�0G�;w�$�����l �$��F	pp.�cW����.�Rf6����Z�ko�}0*��3�a~���X��j��׸-dD9J���/�I�G�Q�`��b�աc�Ȱ�.Z|pu�@�V:)lH-b�L .�����Ă�oïE(\���` ?���@4�X�y�5(�:��8�cG;X�Χ-�`��B�2�F��!�8PV���ƍ<%�pa�(E��Se`T꺋���-m�$��%�Z' !8@*��������-+�4!HAS�_z�I ��6�4����8ˀ�Įk�M�፝�Q0,3��/\h��BJQ��e	�\Ip��D���fPy�ő�,�D�h?)��*.�hL�E)�/'0PyJ���W9�����F]��]�eP�9�f�VN���©ŀ���D mϪs��C�� �Dْ���z�+�%�0�����+M�q`/.u�&mY�oC����>����	[�oV�c��{��l�?q,U?XF�ݺF�9��сf8-�R���H�{FI�1w9`�4W��qÛt�>�zf�?�=a��@�o����ǉ�l�Ғ�J���t��{�OCy���q�%ǂcW��"e�0�j9�e�,` &%N��p?iR�؃������]'n�I(�._�'~����@�.w� H�)[�S�VX!��ǥ8�`R� 7[��B�I8�H�����o�y1b��=����*(�`p���!b�ի駈�Hq��/S/7@(�bP��<I�%*3D�T���qߐ`�G�ڵJ]>Q�auy�a�%h� a�倆���	�)lrXH� W��@I��G�h������z��ѱ�Xs�,���85(�g�N:9�(��'��a+�NϠk4l��s�����ƭaD<9���įݨp����n!�*���@��y��W�N�x�Ț:r=�D��� �yB$P�u�^����it���N�6�yB��b����%
oAHt�N��y�K���TzǬ;e�b��e���y��0�P�$ΐ	YI�MA�Ζ�y�%{bV��R��&̪̔&��y2���TV�i�&��*�WJ˳�y"߰fU��_[�8Ƭ�
�y�=+E�]0�߬[D���	��y/޿Q��(���J�m��D��y��M7|���JA�FI��#v/6�y�E�E=��3.J�6v�B6�Q��y���;r�=@+�|�8�
 /�5�yREI��̰9�ʏ?g�8ݒ��3�yR�::�T�"��*^����$ �ye���6*��Ie8y�D����y�`�-(&t����A��)����;�yBfQ!1q�KƭD�q�>���@��y�B&EV�a&�S��#�K�y���A؀�p%�-C}
�ȇ.W��y�I�L��$8,@)<h���E��y*�4]a�t�wl�X�^� ����yBr��ѧO\Դ�6�y
� P�3�7kZ4�z��U1$zP���"O�8G��2tc�9`��� ^h��"O:�3�<zn$A��+aKb���"O�Uà\���YД/��Z>^i)t"O	s�gҡ� �"VLܥ3?|q�"O���KD1z��;�L
;Ij�S"O�}���-mV�sa-��x���e"OZ�X�쟶W�j�6�ڪ.�"��U"O��˷C��H[��G%ؘ�e�"O�G���'�\]2"�ŰoA�<x3"O��`�ҒvIR�+�Jܑ?���"O�Œ�J�����ɄS�p���"OF-��DW(O��� iP#ir:�T"OX͋�S�@4�
b	ٽK��#P"O$�[VA��`�:Q"\�(�ԤB�"O96�ʁr�V�7��g͢�xw"O�q�%fd��� ����v]�U��"O0���R�;�������w���j"O�B�n�m��c}��D��"O��#�Փ,�hL�"�weT��"OȲ�h,w<���K]���P�"O<�� ��O.f�Y�m�N}�%Ҷ"OP�x��	8h$��0��;ή(����f�j
ç�j13CZ�^��c���h��	A��326�����\�؅ǘ�	�N�cڟp��`9����>�fY�O��E�EJ������'�J1Js��,)�[5�[,`�� Y�%I�|;�h�6:LhT]!!�0-��W-xJd3@�D@�K�mz���'�6�Ilܧ)t�z'�R�WB��c]�	[p�D{�"� ��ţ$bՑl���pG�].�)U�.HB�
q�НjX	K(\y+��0!5��D(Q�@@z��L>���X K�	�2g(3a+�9�6�ؠJ��b�)0f�䐡g o^�F���X! W�y����0����j�C~FA1噥o3\�0���p��Q���(L��W����B�Ȕp�* ��rӂ��Q��,0�X瓁)J��`�m����*C�U؟t�_dM���q#F�!�݁k.�O��#��=�ؗW�&B\� M� 9SZ]��-;!b]B�BE'����T\2,���▤+����8R�'K)�(��6+/pl��ރL�R,+a&Q�s�n�OP$1�Q	w�zE�rFK��	�*3e�i�)9^�K�*䰴��'.IܬZ1�D?v�z�D��*'�Q�B4�\�[ǎG+簰�J�4  \|ě6˖7[%�b��ANpHb�F?l�~Y��/�^$9d@�E���ug��$J���P�پ%�t���@�e�_���S2`�
&�P�<:�ω��'h��	�������cb�`궎��U��1��)�)X60Y`�oWc�O�|%�v�i�����7^����L$�QГ P���@�vbP��o"��i�´���އ8��@e�=(�4p��EE��a�kF5]�.���k5teVyt�i�p|�eB�.�&\SG�D���Z.E�M�5oT![2��`H� �#ª �Y�V5�E������+ �v��WnM<8ڇH��mɆ�
�I�����w�M\.�1���ڗ�,YSv�H�}̨�Ebق�u�1,��a����7'�Y%��q���&}���pQ���<5.TyA��]�`��E(ɗg:��S�T�L}�W�[��`I�Ú�5,PqQ�\�j���i�p�@��8�\5a1��@�6�1�mN�Qaك���^�Cdm�7��p�=�D��:B�2��O>dJ7��W#�,(q��/pJ�*�c�'v6H�[ebJ n(�R�$ޡ38xrGCd݉�R ������M� ���KR.��1W�!��C-����%> ��5�]�0����P��C*��J.t�h`ѢH;wW�`)C���&'T:1�A�8�F��#%˖3�R���$�0���8]�DQ��D�?Q*i1:�H��c��6�ƥ�0Lˢp�*�Y�M�>��a���ɤ0"��<��%�t"08��(�:
mP|��|y�%����ZbՈ^_�9H�H�P,�#��̯$�T��]$�9 �,�0G�i�H��Zwd	��{.-S�ʌ�(﮴��X3�M�7�i�X�QFE��(S+���<J�L�dY�})��0'�t8ð!a�N%xS��7/�Ɣ��aЍQ���I')� 2�.U���ͻ�0uIq�� (��+��GD=Tq�F�d���F��Gh�h��YѲ��ӟ��Q��~���f��/��If)B>L݈����l��e�rېd�(�K�쁾J�V�1㉆�c�����r����?�dC�0R�b`"T��f�3?)D���g��Zg�����E������q\�b���.-"t TH��y\�(qGE+s	���R�F����agĈyH�j���>�m���ܣU.�������Y�È���5��I:D`���ϡ@{����F��s�t��'�?	�iJ�皯_k��׬�;{L<���k�%v�тU&ټu�`���$S=����,��H&���`Ȍ���H��	Ez-�YxK焳b���[�M wݒ �ش,]V<6 �֑��A
3�rE�b�d
�i�Q`��-��8Mty�釁so�\�b�4��t"G#<����"�����jL��M{���QD�k B�^5F�1s�ŌCr6`��87(��U#T�5�\�P���Bh��PŃ�DJ��5�N�4�2�OH����/5�6I#���V�@Wp؁�'�=��	���z9�rh,��	C�8���W�D_`ġ��7��q�B�k�5O�@A��:@ ��O#(=Jl@��K��p=�㨊�� �©ՕC
�$�ХZ@L�)���F@aAT�Ͳ_�]���3�"EX��TG�0��e��CK�='�� �HqQ�N�E��	�S�ܞod�I���6|��`�G�!D���1�70߮�Q��J�`�%ÂnѢz �*�.�����9�H�.�9�w��+ 늄ȡ�'ޞ�x�ޡ.��9�*ݧ
;���4M�T��7�J����!3�1Q����B_*89C��:Np:S�[�Nhg��c�i!�䃀m��۳"O@5��!i�4��K�U�-��oԣi�P
�f,i���%Y3Z�D=�����!k�$��J�]�1��?�,qЊQ�4{�����;S>qqW�'R:}Q����I�Al�$^�-�G��Ỉ*��ǂL��	�E�t����<>Ȇ��NR�H[b#>)���L�-��gY�A�0)�,#����I"m�
Ȓ�G�W����ͅ�?���L���7��� �PjP�����~{3�C;c����>�~��ī �Cd`��4.h���W�˘OX4���7F�c_�3�r�+��c�䆾Wdb��g����l�@���KhHٲ�E������:X�~ex�,+Z�}I�����*X�7�5�`%�h[�$vls��^?GDȨs(3S���``B'|Op9+�h[�	��D�7/�'ZK�����L�_B����ȵ��d��$ܾN��̓�E�(
��P���;�/*1����)���9*%J��`�L/}"��E��ईhb�77q�����iB����E�)9�Ex��M�6������,_\���t��p"C�Y��T���'�&�Cņ�z�P�ҟ����#m�����>�$��V�y�O�K=�!����"2��$ZwHN�3����#_ [�bO q�,�7*��CJl4ң*�e�z @!�|�����#?�,P�놂 �$�'*=ғ2*<�$d>5OBh�U&H���z3!1KI�3C���\j�#�H+0 ,�t�Q�7JHh�%&	� ���C1 *�xJ�`�*��	y��@+YI��XbB% ����'�T8	!œ	C�<�g�[�bR�F�ůdC6�p���uݨ-P�f�klL�
��C�D�,�#M���{! ���M[ڴE�&�0!�:y�2dj��1;,�`�d#�$�1:(�h�'����wjB%@3J(ۃa�0B,�X�(	�^,4F���3��5r�2J9Z&��J4�:�Xtg�W�d�����*��- �)R�n7M�)`+-Ѵወ  B�d@�m|����i�0h)�D��$��QMNU�L02r�IN�bb�����q�,;	p��&h�~F��G��7�n���A׿m�t �w�Dzn�m����~��N>���v�Ib�X{�q1�D�n4�M�-��#�Bm�E'\�>X��F�^݂�9�o_s�YP��8o?�eQA�"�@E*g�6-1��lì��9��B��tL�r@ѳ��� L�<8�e��d��q�e��6&>^��NC�9����m���X@v�P=ii��oڼ;Z�I��B��L���:zz(��#�Z�((뮂2��e�Ξ�J�� ���A9gxU����k�6B 3Z4�
g�n�� ��+'
(�E �*v8���o��mQ���(WBmKP����x�d�@� �
�P���yA(�6]Fr�q�� *QI�V  =(ő&ˉ5���	�FwAMK�=̀���,2j5+'��м�s�L要���.a�����'s8�a�ʐ�[c2�rfHO�]"eɕE6��E��	�/18h�ՂД_\�ioZ�)��(Q���N�R�⛟dI��K�	�|�x�E(�9�A#L��� ��-S��x�2ϐ�m�	��d�)
h��J5�+�5���X�L���@FˬQ��`�2o*d��� ��2oM��ۢ�I��j�@	��I�?d*EL��ֽ36�sSz,�s��SĠ��b9������ʍ�
`����&J�=����lK�>�J+b��#�OȤ��D�?O �p�+^`�����l����,���r� Q���~Cx��ɬZ�0� a��Wp���$�m���ݴ"`�sr-�=$h �j�C�j��M �Y; �t�î"3h��Ξv����]�Ȩ���{�	�B��ŀ����!bg���.�,�y��َL���i1�Y#s�8��k�C��F�)Xpŗ�8�$9#�$��e]����`�/&�t@��	�O(HA�E+O���q�"�X��Ŏ>+��H�T�_�juh�b_�n��ē �H�˵�ֆu/��-SzHAA�Q*w�����<�8��Ӓf9��:G�S^�lMEC5#<R�!�dP���%0���3Q�G�$�|(2LƔD"RyX�R��{J�m��1�5���1� [�E�A���L�@%XuH�'R	��C�j����DP$+9��1C�K�W���Cw�\�r�I��c	6�8(�.]=p��IgK&.2��aӀ� U����s�Y�#ٱ<W�XSf��Z�H7�V�c�=�刄0g�P��`ʹq�n�2�V/���A
 ��r�C�ޢ-P��*k
|q� �8*8$����V.��fA��A>���b����+%���|��J�o��Qn�4�O�}8��)�d�?�Z)jP	H"N�𰕠��8����!�	҈8��j��_���K�91�؀�#M���5�Ϙ<����q#I���*8Ƣh� `�J�8����Շ7�f��q��C~��� f�K��pdI��(�*��G�\a�h���S���0��;-��Yqv� �:1h��:����g�j�˟ԉ��]_٪0�u��x����7NCȝ� EG/]YȜJ�i��Xؖ�H81����
�U�d�p)M�l������\���)�����B��#'V5]Â��Ɇ%>�dL�/<whE�U�On@�q`�CÎ�5\���#�i�$�DS�/�bd5%^:��V�Y�*�����T$Eҥ#Y�h ���ϓ�.��$A��_9��f Y�8��2I6r.j�	���)T.fq. �Z��7q*f�1�'�(W)hmڴ��F�u��$�uξ�KQ)G(��c����ӈ����I��l���Ѻ!�I��m��;�4�1IG���K��5Ӗȸ7S?��-��:��uA�,ـ:��1�Lʳ>��e�s��W�']<�`�"|��R��7z�8�`�AЩ\��a%��;U��+�aC��%��Q���k�%ܾg$�'Pw��§m��+����L;������[��	 r)X%Gj�'�0"�!N5J0����JM_��%@�i!A`����ze�y"Ý�e��PiĆ�P������";ʹFI��El��%��=������OP�:�-�*b����-�ta���Pb���'o 6��]�B�]\�(uF
x�|0�.�ri���� ��W�-V���a�(9zj�Z�l�W�RHS4N��[���s/@�`�EHķC�Ҁ��ŉ��hOL$����L��D�RM�#��=h�$��-g����)�|�	2��1AF0�r�8O��L���&���'0:����+Ϋd�I���9�j��Q�[X��Rf�I#H|���DG�,w4bt�qK\�$��%A3��SꙈ��G�l���bIߐ5s�8{%���>``4��)�~���Y��F�q�#7J��	�tg��-�Dy�$ɺ((Z��c�r�()^��5�3Hr,\����E���B	^8z�	%�� "I����e}"uP0�W`;�����(�6�V�rI8��Z-*Q�+�d~(m���f0�����RŦ����%tN��X3�\�qt����S��@z���4���S�AF�l�H� �(M$wF����]8rt��ƎD�T��4*���7��P�����h`�Ł��uF��Ɯ��AЏJq� ���[e�O
=��ȉ*�2���dC�J� �a������B̟,!텋^h��ψ	����*VPh�OZdi�C��%x��3�ӻ1@��oݕ?i�Yx "�+��'�(00�+UZ�ЭI�N�|��i3O�j
4����[�$4�&_��8ٰ��Ӽ58���j��i��r>ᛰ !X�"4����7�,Ř֠ܞ+�i����murըE&�#�剘��ɉգ�l�LK� E\z�m�78�f�j����i��t)� S�y �2�4\r��X�y�/�w8IQlB�`U6��%� U�
i��0�>HZ�e�Z6�G�v�p��Q�
L�Iw��p�n�2��_`��Dېv�tTg�/p�f���E�#D�Q��ǔt�|�rG�˰>�܀W�&��S6LE:x���+A�y&�pB�>a�@��K�?���<!'˱;�Ԝ+RJ+2>��  N�r��Ke�̺ ��Y�"����;��^�T��K��^,="��� =q�����:'�^���i�*x����.ڕW�n͑��D?[���׍1�	?Z���w퐌O�i�I��L ^�E闝a0~,� ȃ6R�"�RF�/&�r�6C��*\K�M�)%b>�J��`1r ��H4W�>�Jƣ���ǘ�a�l�qM!�2���ʭ�~Bˍ3o�pGIY8Zp!���2|�д	��P�s��e��e��;���Go,j<�q��S*�p4�Cf�5{������f�4�:0�;gY��(��9��kQ}�!���YS8I�j�0>� ]����#@���еe��1���SKP�~��!*�*Ɏ]Y.-!c:�l퐒�@��H c6a&~"�V���m�J�8t�5�s�� $F�/Xd��	3=�<���G�$��EC�R�W�d)�'=�8i�i�.�J%i�8�*���eǟ&���I����@j³y��9���E�E�̭#�ß��$��k%A��b��� ��-�̽7(���5�0XN;0ƿ���j�A��  ��D�Xz��n-u�HI��=h�M��"��+*PKء�2�I$h/�(�qÆ7��=Z�(¿n�A���O),D(��"�(� fصL{rDӸ`�8;�̖�O��E��;��?I���8.�j�լE�]^��·� M$��/��_�P��Ee�/x1��r��+�z%��̅>XV��gc���P� �p�r9ځ�Q�0^���MB���c��A.��b�B�0j���!�$j.]�E���*T(�#�c��{"��FҴ\d��¥C�5`���aSH*�'��Mٴ�8�����O;pQ����Y�+���J��A 4����	�.K�)bN�`�4oFVb�u8u�L�Om �dIH�t�1�晅Ulܐ��>)�Dǁ��TX�Kc7\�:��B?1w&B�]��8�a�W|HJ?I)6ů�pP䆂Z��X��W7+$�e�+?�Ɖ�� �mz��D��p��}��m�7m���a�D=0�,g�O��<ej@O�5
�ҵR&a��sQȤ�c�F$��H�;&�u� �S�`�r�S(>����bD���Gԓ+�� ����� ���WyJ%��*I�:�5��NM�1���q�甒)���}ΓQ	&xU�T�z��xEg��4\�GB��-Rj콊g�U]�S-)���0�ڗf����G	�d0�����i"TӲ,U=���wF{£U�VXޤY�<$	�y�Ԩ��I�yJ��"�ԟ��X �T��ޝ�%,�(+r@ r�vcđ�7V�[ʼ��'�O$� �M��b�P�C��(�d0�퉮H6�t�o�3�툇��4� h�#)T���3w-�y�*��/.�0P�, �f�C�,�?�¢��<j���18���)�/i�yJ� ڀtAʥIGŅ
(@:(*�'���b���
j�a�FNߔ���C�X��J�	[�VXT�GO1Fx��A�x�D�P����e8VX�gi\�p?7�Q���%���-%j�� W9p������N��C��${��,�aj�9Bz�Z�	��6MF�?	�h�,��b?�r�.\����J�9Y���3�4T����D�D�֔�[�}ބ��"O$p�,t9�`7�	X$��"O��"��ʙ��!G�eM��A�"O���f'���!BE��A"��"O���ҧZ�h��l���!6
�C�"O��RS,O�&8Q����*DQR"O��Q&�[�Ew�����3$ �!�'�����)3>A��IK(2X��'�����+�;p^8���A�n�,@�'2 ]₋�D�@B��Ρ�2i��'��������@eH^&	�>��'�u顧G�ZE��6�di�'�~�q��<e㞙s�NΥ C�|��'Y�-��&Q�+�>��ҋw[ q��'��,���ūGr=p��A�78� r�'_ �(�E[�`��ds���\��I��'�N�2��Q2	�N�� ���`�|2�'�	rs �����H�ilPQ��'�v�iB�a��9#�׼_/��R��� F٠u�X7�X(����@1"OE���,�nak�E��q~�#�"O�h�!R�
~��PVc�PP�8�"O�y�Phέv+�呀25M��"O�����Ux������6P{"O5�����X�T�L�z��p�g� �Q�1�ɵID�@��؍�~r��,�A����nJa�0!K�0��7�!�d�,����	6L����R��$ ��Q󏍎#SO\	Z��_��M�ᓸr�C,M!
�<e��S����4�*8���f�pOQ>%�l�]@<�ḟ�G��"(�䘏�(O���Xd'�����B�֤ۆMq�\��`����h�q�|�-8Ց �A�{<�R�e
��M���E':����Sⓔ�e�;b�R���C�C�lM8���=�z}�I
�����+{���ç ���[W��,B4��D֕@fH�"I>�y2d�Jb�Ij>["? �䐤&�:��8��S��b�Ik��C9>���$>���ǘoox�rD��gN`�`'cX0�~���G��?q�$��v3�х�Ӫ\���!M�q�w�EE������j?:��Z�y\YK1�ؕ�`��_��m1��(�����=?�r$Y�/Q* �%C/��41�X#Z3J�;�� ,�5r��OՒA⟹o��h���}��LR�0�\)��Գ#�ȩ�%C:Z�&Q#�UBXH93�'3���Z�[>Y���c�0c㖰^�d,��ڥ-8�J317l�uk�"OI���	�[��[��7%Mh%�L��L���9��J;u�x[¤�����۟Q�֝8�*��a+ <(��s��,@.��'�T"�'/���	��1.��겠@��z�3N�5/��~2G�H�)�'O��I E�`t�I�*��=2�	�~�+�V�i�@��Sp��X"ŉ�
���|��A��i�:�A6?��'e~Z`�FF<mpD�@+�%R]��n�t���'�Jq���O_��gE(8������S�F뼥�免q~���'\����7��ɴN�ڴ0�'LK�3�����O��ض�Y��M3s�J���>�"#��eVT��V2l~� BoS�ovHl��f�R\Q`�˹vӦ�8�ď#@�X���Є�S؊H�ve�pO\Q_B<�ȓL]� `Ջ�::�h,8�J�x�b���:U>P��o��|��ȡ�u��@�ȓ5 ��ׂ��+N�ԃ���K���� ���iV�γe���!V-׸����ȓu
�L���$Dr�@�a�R�"I�܇ȓ�ܬ��/�'\��\*��7wj8��/@)�vG�R\�8��l�1������a$��3rx�v.D>����ȓr��;s��0]:�D�7��zdt���Zb�tۄ�ʺK(Ke�,ZlC�dQpͪc�EP�d������s"O��!K�f���J����f�1�"O�$�٪KԔ�Q���#�Jh��"OtآE��	�dtX�ζSyl�"Oh�P�׀@���y�+U�~�+�"O�=�P�ۄqK�m#�ݿ[���D"O|��uA� ɮ�9`�4.���$"O�t�҂R6Q���eة
�9#7"O4��΅�.Z��B
�M""O`A+���o>,1IDa�Q���W"On\p��)(L,4��	��1���"O<Y0�.#RX��j)Ht ���"O����M�T�B%Ѕ/��*��|#�"O0�`�	I���c:)�	�>Xspm���0d�ղTy�|JG��e��-��MJX���s�ǨE��q�,^�yb��.=�RyKb�^9+�$��K+�y��J=w.8����%J,@ڰ"ŏ�y�F�;-�n�ʐ'�M$�e�Z�yr�J`H�@���|��bý�yb��20���Llk��P5�	��y��O$���2Kb$����3�y
� ��iT�D@�럨=���"OzXCda�.aƔ8d)�Ezl�@"OV��wE�����È�am��"O�#���>��k�슩+E��s1"O���m��2�n��s�K�!�p"O�ࢱDMQ�����AK�1���z�"O�q�+؏X�V Җ&L!`�2lJw"O�0�sOaq��q�0rBE�"O�����Q��ځ�#�|f�ɕ"Oz�W��'#����*;I �s�"O�p�"f�~	�i�uյJVl��"Oqp2�7akj��I��m�x�c�"O�ib�$)bK�2�B�Q�0�`�"O���<� Ā�w��H0"O
�Б!��O��(�r�$%� �!�"OJQ����#���@���1�R�R�"O*#� �W�D +�C�|���2"OFI� 9^�x5Ʉ�	veN��1"O��`ͅwz�١ǚ�,[�0"OF囔�0���С�_�I<�0D"O�uؐ �%`�V�#���!'N�!"O��$��(���s�H18t�CU"O2��$��Xe�L����*!R�k�"O`��ٞ��mc%�^���"Oh���I�(4b"�fU�L�R�"Oʭ��&�eBT����h=40y�"O��!�'���A�#%����"Of���K��҄�WE.�8��"O��J�e^�@���7�.���!"O ��i�X�A�$�	\��z�"OZ��B��C�xH�bDT�X�@�X�"O��K�2H��PgË52{���t"O�`����*GuL�H�+�zy��"O�Z�N��D��(GH�xi�L� "O�)���ŧ`��`�eL>yU��{W"O��+D�u��R#���#�UkC"O5���M�~,�� �O�x R�"Od�R��l�*��#��}��d"O�@C`k§'�I�桀��r۴"O�THe`Ј,1������C�T�[�"ObT�@˞-,gR�x���Di�"OL�`b+��2�MZ'c�-^�B��C"O�tm=VD��L�	���"O����q�l�@K�:H�p(;�"Ob��J٘
�J%5,���R"O|�[��m�$����Z�"Y"O�9�	�G"8�֦\���"O�Q	g�A*e<����2�vu0"Oک���ʸP��uA���N����"O�)c"G�l���a�=xu�X�"O�,8rM�����%��D��"O!T��0D{0\�%G{�N�15"OT����Љ�6�K����J�"O(�jn�!��y��IڒQX#"Ox�n
Xi���AbZŚ�Ip"O���M��c_fTi��J�R���j�"O0<	�L��:��M��i��e�lLx"Ov�B�@�#�A!����T� "O���E�܃>6���	�� s"On)�B�p�<�
�(Ђ���"O|�9��8H�H&�4� ���"O� ߫�(%$G�_�d�B���N!�J))Һ`����"�&�"�OE�[7!�Dɻ��c�"��VÕN�j!!�� ���E��;��0��]�D��I��"OnD�O�0t�|����ؘ(#"Ov|*��[(��\Ñ�+�n��"O9H�n�B�Н�և
,A(�!�"O�ɪ��I���;ֆ̔5,ȑ�R"O,\1Wȅ�~�4x)uEޯq�IG"O~ #�
�yhИZ�.äU��I�ȓf�� 5��J~�S&��VTH���Yޮ(kp��iG01i��LU: ��:�v����.4ː��bc�*)�ʀ��|�)��O�R5PdQQ��#Ofe��:��P���h�1���!K[���ȓjϲY%�A�g�$� �,$� i�ȓ8cJ���Hҟ�j`Eᆔ?��`��}�Z�e��W�u��ᛑ+�%��5z����I^�2T��#��M�Fۆ�ȓ{�<i@eX,p؀�)b)�G|����c�L���e�o�e�"��?wxp�ȓ�����S�=g��l�P��H:"O*)�!ɉ2h���+O2�p���"O�JQ�)�k��-��i�5"Ofu[@��.T~e���m��x�2"OdMKC-B�P��1�Č�*S�h��"O��c� �a�l�3�Οp#l�Z�"O(l��͆,-�P�ڑ�\�\4#S"O���dJ����ST��`�(��"OvMP���2=�
,ȥ̅c���"O2]��gڽ~%X��(�+*��R"O�a�"�	�U�w�eN-��"O�%(��J�e��<�̍C]N�{�"ON(i�����p��K�!�0��"O�Ը�f��(R4b�
�;]��:w"O��K�K9�h�P�H.��|��"OFt ��ZRJ������*�<4"�"Ovi:QD
�3�ܴ)�CЯȠ�Y�"Ot}��^;�P�Iu�<T��|K�"O��LX*��E��I�e�l}P�"O�-���0s*�J��4y�<xY"O����/�M ��	v��F� �XU"O�w�OO���YQ���:�h�"O�kUoєrN�K'�Dg�]�"On���?�*ɀ�i��ShK�<Y��WK���@!5� I��KC�<Y1��>�r\e��a� 9�fD~�<iGZ?6W���U��h��k��y�<�AeB�:M�sb�=l<�c�x�<�ShG��B�$X�;Aw�<)����/��eB��΃����Tp�<y۝s��̊ zG�Xa��B�<AE䎂k�e�fCQ�����&�B�<S�A�U�$Ҧ��HzHz��w�<ylE39��)w钵�	RS��I�<&��8R'�x1U�bD�ia�H�<���Z�8���b�%� <^�Y�BA�Y�<�%"���r�Ȣf\�{�(L��G�Q�<q7HP�FI�p3UMO�K���d�<YqM�	�^Lkj�'Z�xK'�x�<�fNR�O#����)��Et�$C0��r�<��+k@�H���O�:kؙ ��Zl�<A�,��W����.��B�`��j�<aF��4>�PRecĚvμ��ц]c�<A�-v8d���\=��ș%�Pk�<)�N[�m�،	"�W�]�&��a-f�<9EI�%gP(�ɍ��yD+�J�<� ~��d�E�y+7�ȟ=T��x�"Ox�Z ��1�n(#S�MR@�"O�9�3D��#��@`�i
��K""O�m���պq�Z�
�mȗ}�i��"O$��UP�[� d9R'��-�|yH�"Ol�s�*ٚ~���f�!�i�4"O�����X�Q�I�$
�"O�<p�n��pni"1jG�O��]�@"Ol0�ǀ+&��=0b�T��ed���y"��F8(4�3��59�,u����y
_
t�@���8�� :a*Ź�y2&��]���b� y㤄�sE�y2➂m8e�X7`!C��
�y��ƽ��`�D�	"b��	c��yb��$��Yô��l��!Ó�� �y�I�=G�H�c��^��̀����y"J��'��(�fآ\V�<B���y�j�0a4�uJB�}z4iQ�̱�y�7j��\� ��w��������y�ǎp2h�`�#P"r"5�¡N��y"	U8�Ra녓6R�l�r,��y�o[=L;¬y�$YZ�pܡ�bX��y�
�4LD<�C��5Y���cn�H�<I���!�"H9�.�y+>iz�	^w�<���W�T�C���%5`�e�J�<yF�O�W��� ��"A?0)�0BAC�<�Γ�=N�!�2�B�؋FlIE�<��D��t��eGK�t9iP��v�<���D�_)���%K�b����)�s�<y&*� m�!�D�Y8�rYs�<y��U�0g�|��x���R�G�y�<��_�N\�T�%BS�{��(�!B�r�<�IL9W��D[����B��f�<aG�É?�N�w얺psjy���_�<�P�
�B�J����ó�����]�<Q�`   ��     �  d  �  �+  �6  nB  �M  �W  `  l  �v  �|  .�  ��    �  G�  ��  ˨  �  U�  ��  ��  8�  {�  ��   �  ��  ��  �  ��  � � �  �/ l9 @ \F �L �M  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�	�� R��g� �t��B��1�s�Ee� "<E��'�����?l�i�|����y2�6�Şw}��̞�� `�d�ǁ���a����dE�D��p�i^�;>��S��%+�|�L3}2jN,m��+�lRu��iT�y���>�����Q�g�عQ� ��Mˌ��%��|ph�9IV��1�!�;qu��UA؞X$�>�XR��V�ԎPԜa�g��:]&���d(8a�МA��řcYx�h�G��%ڧ\�ƠB�!3]��`��G�44��^�Ȅ�-J�S�d�Ӱ%�'
<�'Bў��$��Fa�,ʕ0�i�9j.!�$�!i�;��@�f�I�Iſ+� �牰D�-�Dk�;�Q���c�C�	;<�4Qd �
����'�4��'��Bm_�K;�HاA�H5���|�����Hȸ-&�tbr�Žp#��v�/�yb(Ͱ6��9�L��o�(��^��~�!�S�Oaƙ�gh�[8|`c��e��e�'% �;?ʡ��� J���
�'��s0i�3y�Bd˖��Vy~9�	�'�F��A�^_8@�D_�M}F��'����7�[�Y��:C��JF���'�*ex��N�d�B��9;� b�''��SѪԮ4	�#"K��7cL�8�'����d �el�0J�g#����'�HS��Q��*�р�	����'a�|@0l�9�0�p�A|�`<��'/x2���93�]���:%���`�'W��P��҈4�����)뎨2�'R2K����y(J�0�D�Z"m��'�~���j�$)ԡIg�0����G��O����^�E�� �9rdx05$?��{rɚ��I�m#��Q��Lm��$*Ǹu��ʉyr�'q�x��H��t��ѯ���r�H0ND$��=�3U����"��M�霂���.�69���ȓAR�L��/�B��ǭ��-����=���?Q��Ӟ6 ʝ)��^�%x"T�&��~�<Y���7?=f` ���4~D|9qM{�<����J�Fa@o�`Ѡ�sS�Q�<�[y|�d[� r:���`n�EB�`�'F�|�ڮe��)҅��F��b�O���	^���O(���b�>�bI����O��p�	�'eF�Js��#y��L�Ǆ�U�
yK�}�x�鉷4��9{�ɐkL����N4Z�rB�IlZ6�+l�	<�ؽ���Pdֵ����'] �cV�`����jG�%��9�'jX-���_�"�ba던�Da	�'�bY��R&��l�� ���$��˓�(O��5,��N�R$�7/T�j�~�J#"O�BS�]9af�K��G�Y;b�s���=lO�A��ydVEk��ה:0��"Oȑd<$�X���$Υ|����"O���t.R9ǎM�1���S
nj`"O�:AJ���,������eh�ha�"O\�!��שn=Ҍ��$�	'�<Y
�"O��#@E�U��C��W�9���"O�؀�J��}:5��k
:�P��"O�D�G@فE5ZA�Cj`D����7O���df��	Y0i؀}�~��)I�5,�,���'���ɉi����AE\���z�&I����5�I�|9������?& �S &�T|�B�	���0p#� ��� �<}��B�I�Jz��5B�% dY��T�A�6�F������ ��A��ƛRTV�BpH�>���6"OL�ke�I�Z t�A��V)(��2dU�p���h��Q#w��
T�� s!�F�H�ZC�I,A:� Iv�CQ��2�iħX+`B�8P��(��_�!�l�s�H�3
R>B�I�T=dX�!��N�ZAz���._B�	,$��rVk[	l��-q-�)
B�I�e|Lru���Z%��� $��>r�C�	0����ThW]jP��-B�6Z��#��c%O�>�ȉ0�F.`�����4�O��$�QԅƪuJ�AK����>���0ƈ3D���� 	F��AƂ�5�a �M2扃5���?�|b���b�c��$��iIGhd�<�0�� T�4+	I����a�`�'O�yB	Q�$�� ��>;L@�cc/_1�y��%&�&aYF.đ-�E �Ј�y�C���v�Pg:��P�7J<�y�n 'Ǻӑ%�0�؍qbC��y�ώ?~�Pt,(t������	�?����v\8���,�H�Pu��!i|���ȓ@��-Ӥ@+n�P�Sd݃B�v,	��O�����!3��q9�(��D���fcҖ^����)"?��,�;�2%��۷�����(�f�<���H��z�eZ�j�
1I�<��l����v����¡К3^lm��	�!n��M{�O��e�k�!�"��"bN؜�"O$Iǣ�W�$�����w���S��D�O��s�{����P=j��1���{�|x{V�D˟̄U24�K4�ҔT�X��CDP�(��:g(I�&�ݱ*�������>�rԇ�,�*I�K�J��f�3��!�ȓ%�M�adT/J�������n4�ȓ�Jt�0o�zB]��j�b���^=�P������[Ôpc���ȓSܐ�bɇ,�����ODN�ȓ&��MJ�� m=j�%)F@�م� �]Y�Fѫp'T�C��J�[@�ȓ?�,�B&@�����1FTl��b3�Y��N��z�	d�.n�B�ȓ9����[��䪧(Ų!xPl�ȓI�@��Q�(]�r�I�Z<��O6�dұk������@�]�(��׈��H $��<1ѧԗk����n�hU�ݢh"69YŨ�<�\�ȓ[�p�Q��L�r��a��_p&ȇȓq_Mb�o˗%�@$�+�# �����<_p�+3
�h�F@�3$����@ua���7���9�'A.S�\�ȓ:����<%�.��P)��(����|��6�Ѯ#���ޠg��=�ȓ-�E�� '��ߓ4�� �ȓ"cr�@�0!{�	�fΈ�
@�T�ȓu+�,J�$��P	�)+vN6Utz��0܅�P/ٮr�\��v!�h��x�ȓ^��`�$5)x,�N8�f�ȓz� 8��O�]1l�RT"�39���ȓ{/������-��$~(�ȓi<ش!ĭ�_<"c/ק!а�ȓi�Y�&T�w�^��n�%4P��ȓ*�f�K�JB�$
��R�ĩ�ȓx?�W� ❩3 �.��\��`�Y Th.���)˯vD�ȓM��R��+�:v�Փ"6E�ȓz #U�$ut�A��7-�4q��S�? ���*E��t��Ś���(&"O�"&H�8��U��e)���u"OnQ�A��r<x�D+^�@:8�W"O�h��&Y���k��N+/���"Ob�p����U ro[�[Ά�[��'��'��'��'&R�'�R�'Ӡ���J<OT���ʗ/p�4���'���'t��'�"�'A"�'�"�'�4�Q*J�$BLc񧆈aR��!��'�"�'HR�'��'42�' b�'���D��'�� �1�u�3�'��'���'���'���'���'h�v��k��<"#��>2\�E�$�'���'���'vB�'R�'E��'�Dm٣��"D*����Y�r<�f�'���'���'>r�'���'��'&����
���`}�&�ȐF.Jp��'/��'���'e�'1��'��'"�����5`�P� �R�F�RC�'Z��'{B�'>��'ub�'�r�'@����k5c@�A�*�-5������'���'�r�'e��'or�'���'��)�ը���e��Ȓ?'�=�F�'�B�'�2�'#B�'7��'���'_dQWhV gg�0S�M��˂�'���'%��'��'Q��'"�'���AЂ��t��!�,�W�'{��'�B�'���'���'+��'u�� coK==�vlz���f�R�*s�'���'��'���'R�a�����O�Ձ��	{����rrgjm(*O��D�<�|�'*7�Z�-	�&z����g�8�Y8W��D9�4�����'�	�"�� 5_OՒ8S�	|���'��U;f�i��I�|��OO�A�&�ۧ�U=��d�aM�?�6i�<�����D?ڧ��;"n��d��PE�,T�+�i����y��i�ʦ��4uu�i�����Kt)۱��
}gJM���Γ���I�k�\6Mm����&���@Ad�p�t��q�q�PΓE�Hx�����'���`��\�#�l%@��Y�F>rU�'��	n�$�M� HKZ�2�i�Ǭ�?�B �B��}*�2�>��M����y�R���V��ctK�����0�GH>?A��Ǩ�I�PO̧ƪ��P��?�gM�i�J���ì��q{�D�+OP��?E��'l�����R�\$�U�g���Dl�c�'�D7��7C��ɽ�M���O몬��.�j��m)'N��-�'���'�R+�>�f���ϧb���"�#e�ɴj�:"��
�.��^�z�%������'��'�r�' ��;����"�cg&�"{T�i�Q��3�44�ݳ*O�d7���O8"�)�f��dAb
1VH�U���D}B�kӠo�1���|�'�ZT��CY|١��C�~0��/�J�9ї%$��ҿp*<y���t�Oʓh��مϋ�!�x�b�H���񉒎M�����?aPB�9S?�-ၩ�3H�0�5�?���i9�OV��''�6�_��50�4���Y'� wh� �gjފ�^��Ğ
�M��'�b�Ӝ *$������?�\c��|;��� y�ڈ�Ai���`ј']b�'�"�'�B�'��OKra�	�
����G4�l�-�Q��'��nӀ�2:����O��O=*R�O?'�ে�8�8�i����O�xlڶ�M��'L�xݴ�yb�'�͸����w0Z|�F�b�uq��øG��z'�E�m�rP���i����?����?yCP? ��K�/G&⌈uI�!�?����?���_�ၣ?�?1��?��i(�TM�q״��I�o �f�)�yr�T.��|·6O���b�0m�;m���|���U� ���Mdld"��,PVX؈Tɞ�4F�TP�U~��O@���+��'�d��\K��u8��V�ʩ��'�B�'�����O�剠�M{� �c}�M*GB�9T;�U�ڄ?`+��?���i��OH��'��6�� /���DY)l�`�#���+T�l��M5c��M��'���$�@]��&<D�	Y<P��q	�2oN��$"�,���	oy��'4"�'�B�'��R>1ZuK����T,�2-��$zSˎ1�M�$�Ӛ�?y���?QL~r�	���w	
M`��G#T�� fJ�0�h�,p���l���|Z�������M�;g��M1RL�(6�����$S�u���'��r�
�O�[M>y*OT�$�O��21f�W0��T	̙t�-#�D�O(�D�O����<�i�1�T�'�b�'g���vHژ2ȠD��r*�2�'��'��֛&�`Ӡ}'���A�'Y:k������Rmz���ɠFi*5�A6+�8��'������T� �'� �W�݀g)�����T��j�'�D�eZ�Fa���� š�O<�oZ�\1<%�I,j޴���y'�U2j�r�@�ؚ[R�j�ѿ�y2�w�o��MWo��Mۘ'D�A��W����5j`�p�5�Q.p���O�T�
@�ג|�Y�����d�	�l�Iş�Jpm=Z�FM��aW$����@k{y��|�xz���O����O�ʧ�?A��)���#��yJA�ͅ.���殮�ش��9�I矼����+��p�Mb�F�2�)х����R��x!�	�u�u���'�B�%�d�'�h��6�I�>���;e�PVd�4#�N��FL޸b��߱2�A"ᦂ�E�h���FbBJj����(�O��l�M�i��a!Q�{�|����0��A3�(XYr��3OR���=F�Y��3�0˓�bU���  %!��G8*mhl�cd�4sn�J8OzB��6#��8�5��i:�i���O�3�|ʓ�?�Բi��M�ΟJme�	�ƅ��Q�vx�Tb����I<�#�i��7-��Pq��g�������$\IZ��Q+J�/N\��,�z����4�'��0&���'���'4B�'\`�[#��#���Ѡ# b�����'��^��
ߴ_^Z����?�����	A9L[���6�ۤ.l�YiӤձK��������	�4x����O�� X�� �.@���1�����I�$��ӓ傓?P���?Y �'P�@$�8 F�C�Έ��'X�l��m��EA��Iǟ��	ן�����	yyB�f��Yk�����;�뚙+��2�n��d��$�O��0�d�O�˓e����9.Bܣޝ[�f������qv�6�Ȧ����QΓ e�q! "�|���	�?�S�o�H8�nO�(�f�QH�d�7-Y�����O��d�O\�d�O��D�|��p��$�%U%���)Dd�@��igL����'gB�'��Of2!q��J�0<p�[dҎ}-~ 
DU�M:`to��M���x���Đ/�V?O��	�g�Pn���5A��[!D�v3O&	AĦި�?I]��'�����T�	=_'�1��Q�l��UA�fDll��'���'qrS��[�4g����+Ov�$�*Q�qFo�'V��Q�T+<?\��ЩOm�*�MF�xB�ց�H��dK�c�J�j��y��'�� 6F�
� �QU�<�S�>b�Fşp���_mQт��[�d�"�K'DϟL�I�<���D���'~�U�C�W:�pj��8��'7T6��<<oD�$�O�n�ϟ�&��(msh)�^��*�#T�P�X�:�M�@�i��6m]<rհ7mo�d��*3F�#��Omh�S4�L,5� \8�F�QE
�!Jl�Cy��ѬxÛ�:�͈-�B�� B��j9,����<�� ɉ�r�%�A��gn 9��=D��&�MsöiD�O�����IǬk��-����~4���A �73�t�#�ԢNR˓[xĨ��o�ֱ��&�	Δ�qR#J5 ����k���Fݜd?:���G�����*�2e@���6"@�BeP�1O�G�Z���ІPW�K��H)�|0�T,�(ކx�3ɉ�jÀD���Y�,�9�O��3���r�-K��M;�_�:�����QîY�a�;�J��\q��PR2 �q�u:�̍��tx��M./(<�,R�	���Z�ʊ��\0��E����C˂�/����aK4�,0)q��D9`��#N4*���J�S�x�T�Տ5&�Ā�eO'ސ�(b� v\���E�	?Y��kڴ	E�Ю�pg�����|�B�JC�M�	ş�&�H�Iş���!�>Q$�
;M�(h(d>)���]o}"�'���'��I�$o mM|����(p�q תډT��P�q��2G���'��Z�<�IğLq�� ��8��ݙS�2^2��B+�'k�ߴ�?1���DΠE�>�%>u���?�؏k�V|s���i����/	�7�<A���?����ş�?Y��ae���4A�US��K'&	��u��_,�E�i�P�'�?1��%��� �nU�4�3���e�B7��O��DZ27p��|���&� � �߽�&�	I�bX�=��ArӀ9�����I֟`�	�?!�L<ͧ,�>]���R�KK�`�S86Ҵp���igt]�gY����ş@�3�	ϟ����ng�*�Xڱc�]3�p�۴�?���?�,�Z}����'�b�[*T����S"	�]\@�j�!����?������<���?a��U�X �뙎`h� ��SY��s��i�2.���6O�I�O��Ĵ<	��Ka�x��ꖓ=	����CUt��6�'���x�y��'�R�'R�:ߢ��4چ4�>��&[�wT�����?9��?�(OV���O���w��M�yy���q���!NT2^1O����O��<b��8%�󉁀[7fT�#��$z�
3c�-!���ݟ$��؟�'v��'6������)�/�B|����k�i �\���I�d�Iyyr��/w��i���4��%��E@)S%v��l����	q�Fyb����O&,ҲHG�*�pu��,ك`�Q�ݴ�?�����ܲ5�d%>-���?�أ
��T���
�8S��D-p7�<���?A��^�'�?y��e���4	F����Z�����&yӼ˓O���i=�맢?9�'eR�I�W�S��;��p�F��6m�OP�N,�S���ē@0�PϘ:�@ L��N+�1m��Xz�I�4�?Y���?��'Gꉧ�4��!�Izm-W~����,E�6]&@L���?9����<q���Ω�tʜ�X?JMP���eȚ���?���?���T鉧�$�'*��Ԯfޒ1�BȘ37P��.����?���&��a�<����?��'��eX�`ҹO�8�Y�M H^q��O�Y��<���?1����'Ɔ����|h���m�z:���Ob�����d���\��ty��')tDk�lQ�k>N�e���Q��̛
#���ן��	�8�?	���z�@�����-C�K�t$,ixi��d�'���'�I��#j�s���qTJɠ6i�(1P5��ܦ���蟨�	a���?���$�x	nڊvW��Y2�ŦgΠ�1F\����?a������O�y�,�|���)�j��B¢G_�4���@P�d9�p�iW����O�$:s. �|��'��[$K�{�tu����$�
�۴�?i)O��$ڦ$���'�?����ڷ�E$3��%��3�����Ί�D�>���x����c�M�S�Ĵ<�@���t�4Ś����'I��T3)���'���'+�$X��=� �)@5� ���eŘ+
�ڑB�Q� �	6Բ�!a+�)�n�v]���D�J۔L{�j�$��7M�%5��d�ON�$�O��i�<�'�?���P[�]��n9D�����+1՛��ڕo�&وy����O�mq���'-��*��H	:r	h�o������|yd�5|��i>�	ȟ���m�t�Pn�& ��ip�O_$�`Y a󤓟rꞤ'>U�I����rȠ����R���r�H�dIo����8##�ty��'�B�'�qO0L3�m�,�2��F�Od0�]���NY�j�,��?�����$�O�db���	"4�2�k�$���d��.<����?��?1�R�'e���DG�\2PZ�d�v@5�R,ֻY���OX�$�O,��?�f.W��d�߃)����HM!S�:�X�KD!�M3���?!����'����!z�d�4ZFP9Cĩܱf��Q��Ԛ	9,��'���'��I꟔�	�B���'��- ��{6����&N�yBv���nm�R��$�	꟔*�ǝ%G�O*����M����%���B�tb���'��	��\ j�w���'�r�O�zͰиKB��SEȠ*�v���*�	ly���O��isLY���U8-> �LC%ZZ�	ޟ�[�B@ڟ`������	�?ᕧu7ɺr���f��*�̹p�"���ķ<�#�y��ħO<Xc��=Db�1�J �7���l��'����I��,��ݟH��Yy�O2���~���P%^��=ð�E�Nv,�Ox�Ex����'�~,+P�V��L!c����� �s���D�O|������|���?	�'7L�3˂=66�A�4�Ӄ,+�	<Hp(L|Z��?A�'Θ��#+n;�a��cHI��@��O@�0�/�<����?	����'��0k@0z�D�!K�>��	�O�!i�M�&��������Vy2�'L*�K�D��?q� )s�����)�J*]������4�?q�r��hc�Ϥ�@��D%/�M���
I)A�'qr�'��Iҟx��JLR"�J>+�
��p�GGp�tZ e��u����p�	[���?A�L�.tj�lZ,δ�A��Mk����đ.J��?)���d�O"���I�|:�'!�a���EԖ�Y��C�?�~<�ܴ�?1�B�'�N �W�V1��]c�p+u�O��0C��B�~ H�m�ߟ(�'���91E�ӟD���?Q᦮A�b�J�e�̶a�*�!����'u�IV6�t4ъy���$*eT�Fb���˟�X�Z�
'Y�0��+���������	�X��{yZw����"��+t�ur+��ҫO*�]Iz��;��i��^�B��b����0QFFS�����Zd�'�R�'��TW����D����_,��[!C�j�z1�����M`O�� Ԛ��<E�d�'�~�P�*�X�P�����l_��7�h���$�O����#y���|���?��'�n`@�K\�� T�pæ9�ɱ8��8I|����?9�'�U ���J�I26o�)Y$� ܴ�?�X��,OH���O��d2�I�&
-��C�&�d@F�@&\��;�ti7��M~��'B�Z�P���>��P��N�<��8q���s�T�Є�Nqyr�'J��'��O����zp��1C�"Ԩ���ᎷG^�8�aF�l��	֟d�I]yR�'�LHk�ҟN���Nh^��5! q�T�t�i�B�'�"���O�u$b2,C����>+	8�sS�z|�h��#���D�O���<���:�0��)���d�z� �x��7!\8(��y&	mZ؟��?�bR>�W��Q�If�����;1���`� 0j6M�OF��?q6'K���	�<��';���	K�,�,C�K>B������O���Wˁ�S�1O��9�`aS%WC�����f��3���?I@Ö��?���?����B)O�n�*zb.q�5��
��	;�~��	�,�G�� j>c�b?IkU�� <���"D�dIV-��{Ӵ���O���O�D矨��|��-�|)"F���Bua�1C�����i2����M������$��QH���G�P⺑Y�\7_,,oݟ��	��@٤�EEy�O��'����-oT�k5Ø$/L2��F��<OD��<ɦ.8C��Oq��'���"H�I�'�U�Tb��2F�"g��	����'��'q��D�&:�ۢ��N�|�R�N[���I�> ��l*?���?�)O����W��˰���#v�<�		��ȵ��(�<����?)����'�bL�6}楪j�/�� ògX
��j ������O �ĺ<���U��X�OpI@�hE���ۂ�#"���2޴�?!���?�"�',ht�%ǣ�M��Q�	�>��GNό)�� ҃�l}�'(�Z�0�ɓ���O=R(�}()r��ȭ&$luG�@�%*<7m�O����I��lK"�#�d0�4�@�ǉQ����,T蛶�'V��ޟp�*�L���'~B�O"�1y�����-h��޼7�F� ��<�I韤HC,5T��c��']�����43�l�*���U���'�2�?���'K��'��t[���$w�����}����$/Ui8��?���ڮV��<�~���R�}��u��՟
��p�sN���q@�
�M;���?����Q�t�'�� �Zؼ6%ޗe���Aר�5�6��]����Z����櫛�A.&�bՁoL|���i���'@rL�oɒ�����O��)� <��de�2yR�B�J
眑��i�2_��B��v��?	��?�dŎ�uP��g��?245)԰>6�f�'#�u�c��>�+O����<���[AB#hc��J�1M@���Q}bKG��yr�'2�'��'&剶��2��,M��؀@�ܙ۾lI���yk�����O�ʓ�?����?A���5<m�a�Fx�ڴ�$Y�-&��<����?����dRL8ʹ̧q�:���Q\6z���~�L�lZay��'|�	����ޟđa~���Ƃt��hC1
�@n�p�T��MK���?9��?�,O�t��`���'ҽ���W6fV�����c8J92�t�����<���?��bJl�' �$�K���f��2ZF9�gH�F6���'�rQ� O�4����O�����T,�!Ck�F�u��H��X*��t}"�'�"�'��c�Oh˓�����b|X���/'w�y�C���Mk.Ol�1σȦ=�I�\���?��O��I�@K��3S�:
����C����'gB���y2P����Dܧ~��ըW���+���l��A�m� �h��޴�?���?��'���ny�F.Yʲ�A#*�1
�.8�W��]w~6͑�-�=�$9��ӟ���Ǘ'��
�9&�+���M{��?9��`�vS� �'I��O0���MV7faL�Z'O�1��-+ķiq�'l�ڟ��I�O��$�O�|S��.�D�u�W6X��]�b�ۦ���<!���4�?���?��*���R?Ʌ�J1s��qڱo	/"a	c�UR}r�V��y��'���'3��'��9x�J �0BD=Zº���b,���.��ı<Q������O4�d}�X�`$2�Pxrj	�t2R��#Ρ&i��<i��?����򄘆"02�'^�J�ɆjȳI�Bu���2#�,<mZky�'4�	��I���Lt��⣮�e>P��ģ�r��Ie�V�M����?����?a+O:�A��y�t��5�cM�o��g(4k�Z u��=�M����D�O��$�ON���9O
�'j���t!�d�#v
��C֌�r۴�?)���ǖO�`�O�r�'��Tj�((YnȲ����#�i8P�h��?���?��D�<�O>	�Oz��h`	�I!�qaV��9f���4��Z>:^��m����Iҟ�� ���� 0���'���tB�
j^�E�A�i�2�'�`Tə'3�'�q��P놀�"|8�2��sn�l�T�iTz�Pt�b�����O ���~T�'��I9L@HhۣZ�4`@p0-2X�޴Rfb�ϓ�?.O&�?��Iͦa��	3��mX�ED����i���'j�e��d�>1+Or���`0Sힰ�H�[D��i}��s~Ӯ��<)�O�<�O-�'�B�ޢq-����?8��-�u��,,�7��O�us��x}�Q�0��My��5��~��,�#ƅ�g�eP��?����#h���O����O����O>ʓ/�V|���L��l̘ n�"j2}hM��#�	Fy��'T�IƟ�I��[�h�,�H�Q�	e~�GM�h���?���?�����$��k�I�'�\$tI�C���ܿ&|l�Iy��'���ɟ,��۟ a#Ag���?%_�e�@$O	$iݒ���/y|6��OF���Op��<QńN�@��ğ�� �����)#H�!��M�K�N��?a/O~��O �$��* �d'}/��m48�����!X�5ӽ�f�'�R^�x@
�����O����Lm�pe�->@�M	�,Ա+��V
�g��I��Iڟ ;��a�'�0��.f���+�'I��J���aZ�o�Ly��U'^6-�Ot��O��K}Zw �U
A�ٳU�"	�U/X(eV���4�?q��WԂd�V��s��}j�-;cr�=Yc��-i����gB���wl��M{���?�����T�@�'�ؙ��a?.���@�i ���$1sld���
67O<�O>�?��I�YE�-��KV4VP��)�7�8�4�?���?y��o�Ity��'��D��U5 ء�&

�i�IF���'��I���)j���?��U58�A�$Ej4��a!�<+T�P��i3���0�*���d�O�˓�?�1�J�iV�O?4�15��6��ml�ޟP"��m��I��p�I��L�IayRIK}��j�^-A�X�"�K�9�`��±>�(O��d�<����?a�P���A�¦�4"�"�SI��c����<Y��?��?�����@�@�5ͧ!��� �Y�[�Fkd
�b�%��IP���	�:��	xb���B�5f�P��8���OX���ON�d�<I3jŒt��O��@R!T$fu�`�7a�nl{@�~�H��&���OJ�D�L�O�=rv��v.Va��כ�i�W�i�R�'��ɏ.�� J|.�M��'oGh�@f�e��K��}`q
�x��'�B�Z	���|ڟ��,�.Tc�I�!��)6�i��I*+�drش}�֟$�S�����$��X3�Hl���^�a{�iI��'y�H��'J�'�q��uBM�K��Q!闆Qkеˇ�i�8�[CB}���D�O���䟸�'����j��2�K��`,�q(M�%��)�4F�������I�<y�z�<�QwHWa�p�Dn�&�:���i���'���@)vb�0�	N?������	1 ISPE�q�T!f��<����?��� #�`�K3|c�m�HR��ŵih��.bO��$�O�Okl��0,lY�e�Ճ}��k���"S�	P�'����П��	KyAY�ܓ��ݰ/����@mO�6�:����!�����%�T�����p� �Mq��N�&�PQYtkSm"�:��H�<a*O����O,���,�2���|�a�T`�@ ㊊D��ѡ�F}��'5�|��'4R
�yR��>�Zq�Y9$���+%��q,ꓠ?���?I(On�H��[�St|��j싈C�0=:*�
߆l ش�?�I>���?��߹�?!K���qaJkLXj�ኩ3p ؁Q�a�R�D�O2ʓ1�n�����'s�t`�?f#����BQ�p�tjp	�3Q��O����O�L$��a��HkS.4�#�ɪ���5L�:�M�*O�<�@�Qӭ������ ��'mzIV&�;�Ν�A�X@{��ش�?��S�N������O����B��:w[��31���>�P�b�4�Ԕ�Ҿi�2�'���O��O�Cx,����=����G�q��oZ�:g2����l�����䜑f���g�=��/i� �ӗ({Ӯ��O���B�6���O��'�?A�'k���0�܇��b�)	����%��#;
b�0��ß@��#R(nBQ:V�g�V�I�Kٴ�?�S�٪��dXJ��'��'K�<z�H��(9���R�8M�$�`�C�>᥌�%�:��'���'k�X�ؒP��,�[u��g�j	��K!� ��O����O
�d�O��4���-0�xl�iA�j���a��{.4�&���I֟d�����	�%�� �I.0�X��
zp`
5�+>�"d�޴�?����?�M>���?Q�cS&�LoZ5���9��x�!�NH"Z��?����?��?I���?��?1p`��E��	+��H[��8���H����'��'���'��x���ēx\�	�#��}@��.!,Vx��x���O�˓5��1&V?��I˟L���0d4��h����D���0qݴ��'��������k���W�� ��zk4�r�ɯ(����'B�S���'�"�'���]��-x�&�6��L�풐\�$��7��Od�dDn7,}d��ɘn�^	�悅�:���Q�ĶC���%U�a��'1��'����'0�O�,Y�'�U�fp@���-M3�X�r�Ql�qw1O>q�	$V1���c�F8a8�(�$-	 ���4�?���?�oȴ~��O������
�I�]�LU(�,�D]�p�/�ɤwǌb���	��I�&���tn�	tL^I��e��ش�?��g�+щ'$r�'9ɧ5�+��&Y�����`����Ьͷ���D�H1O����OB�$�<��́�BG���h�:JUp8�v�.[ ���C�x��'��|��'��&9�*��C$��.��q�GRg^��q�yb�'B�'E��'A�)x�՟��B�,�E��hwC�7����Ƴi���'�җ|��'�R��$��D5NG��;�U9+�Aj�mF�^�I=O�2͉�
UJ�0C�e��K���b��b�b	��t<�fPS,!�Ͼk)�D�tiڱy�
ي��� ;����JІ٣&��Z��0�qg��T�9
D�:d�T��[��{/}R�̈��!��*�μX�ءrg�ŗ>��S$iӿ|� *�1A*r,IS�;K��kw�Ūt�h���g:A�y��e�a��&k@8:cn����::HX���]��`r�d	�4/���Ȃ;,��'xb���Xff{/F)(����e͊��@]�&a����\끍�<�O�1��Z�K�&�q�ʐ!2�@`m�%t�4q�'j��'�*�p�%�<E��9!�0���L�s�(@-ژ�#b	��?�U�iB��?�G���B�VEJí��sڎ��5�M.,�}ϓ�?!�kl�hj�l��f���R��*̡ExҌ=��|��P�T�Rf	R),p ٪MH���?q�cJ�j�Z���?���?9p��4�d�Obe�3�H�K�<iEk2[��Ѓ�������ދa�����ɀ�x_����8X�-I�^i�$�
)U��I���z�)���%iX)�Ac�?�=A��K�1�����#Xr���/f?qE�N��	K�'*�ɱ=/,M��G"j,I��g˖|v&C�I�Q�LݑTg��W�Zpjf��3����?��'�9 �kd��x��Az�.,�s([���Tg�Oz��O�$�4u����O���:/0U0P��YR$!4�3
�z9�fb��e���	t�欆�	�:�<�r�Sd��X�1��/D���g�1w�t�б���)�T ��ɰv�4���O0YK��'t����@�"��y��#5���O�!�5υ5pء�"�F�"�8�Y�"O��dka��i�D�E`i�1O��'w�m�~9�OV���|zC��_��Q�@�	"��`�U�g�Ƒr��?!���U0��!`ʜ0��ƍ%�*����B��e6E"��N�U��)���u.Ri�A��-��Cv'��U��E0��Qr(�fՔTf~ИPb��x�,�Z��)$�2�D�O�?���e���"e��*��ayzI��@w����g�$]�q �%�� S�S	�n��$�g�I���;��7G/�[d%�.!�I�M�Pms�O,�$�|�[=�?!���?���\�	�&�=!��d�U�>0qf��&�(G	��:���kB*��c>�DHh[`T��ֵB@Z4��U�D��"��Ⱦ�*� �8vj�ZE�ċ[/�"|��0�Q�)F*46t�&�Y}�1#n�l��[~J~�J>�W�+O�)p��L�|�G)T�� �؂ӫ
0�;@D�1r�I��HO��@̂�`#�H3�P���`���N���ßD��@�0����ş�I🀺_w�r�'��<I��f��03��ӻ9�1R�'(���@�:��i�b�=O6�Q�/*�n�� �űB^����O���-(AB���d�\8�\zu�Yk���h����o�b|y4���DD�O�d-ړ��DٛWuh�Av�B�o*�d��U�#P!��B�&���j�����ЙFzʟ�ʓ(p���i�����+�+:�bU�۠s���i0�'���'�2g��r�'�)�;C�7��O��g)�%L��� �'8�����'>FdI�U� C�	Z�)f8��W�ޝD�0Py�"�O-�p�'4R6��k�}Cq�
Y�`4�f�@��lZ���'����?Iْ�E�JJ�	qn���}8��+D�p`��,s����VW$հTEv�;�O����)�f�i#��'�d���1Q��+ˌ�3V�	����Wd�ޟT�	ៀ�	̈́M*bx�<�O=�2
IC@���4^/MD�6�I�����8�'&��Br�]#0ƴ0Bp�D=5QGyB���?Qd�i��7-�O@�'k�����L��r�Q���8i�d��������$�>q�ar����#u�]�' �a|B5�dT�!HZ�Rag
�Z$�C���1�d��|5��m�@��c����4-�r�'�B� �D�� Rq4���m��&��,i�bb��g�';P����D�:�Dȩ4�1X�r�s�c��k���"~�I�L��9jЅ�dN:ܹe�%�Fф,�Ɵ���W~�'����@$'� P�YN|ڴ�	�yr�'"�}���0k�r7�Քu����׾�OEzʟЀ*���f�N1���8`u��,�Od��]�y��1$��O����O���C�����?a�N�v�t�V�X/%]���1�T?�qa��r�����ɝ~�fZPhӨ}��2�^�97���u��mCe�.|O�i�˂�����c<�2���O ��J�O���O�Y�l�	ky�c	:=y����`��Ph�Q81����y"�E�|�E� �P��qZ0B�Q͠#=Y��J>�?A*O�,�N�˺�AcErx�!)ak�/bv����X$�?Y��?��z�bD���?A�O4���,�%Q�6��D{����F�mS�p��d��p>�����k:~,��40IT��Å>@�n=�ND�I�l��I��<��Ҧ����M�9���JG�Z�R ��S�K��M�����$�O~��'|�>�Q�NV�0T;Ǡ��d�ȓR�]8$��WLu�pJ�k���%��Igy�Sp�7��O��d�|���/,�#�JD�
���F��%f������?���bW���@��&ul�2�M�u>\R�W?c	 ���1�q��EN*=�$ʓN��bP.9%�$�Sr��q=��s����Ol��Hܷ	LY)G�	r4����ߦ�޴�?-�8�jg��=0���ǘ�S,��4�O��"~�S��8�E.��������/->4��I��ēz�� ��Fۿf�\選y����'Q(|�d�+<b�'�"�O�0�b�'/R�'6M�DcO�xq:��c�Z������]0����:C�@�C��ق�^_�����>��X���W�r���J�ݬW���c@�lo<�P���-f�ih^2�&ܘV��A�pIӶX>��
I�����l�\$�i�>�l���I)�S��?9��J�e��Ё4W�?נ��7j�]�<I�!%Q|p���l�$-�'!�b�' �#=�'�?���3�L=��#��p`Ze��͑!�?9��:wuHiK�?���?)��ta��O����	o:X��F�7j��%2��8|h��t���=lO\5��I�G�(VV�=v�� ��O<��ѩL9z����@���&=?�5��f�|H����?q`n���Ӧ��t�'tRT�t�WD�<nB��pǮnt��d/&D�,9�	��q���a�_�9�<�(�� -�HO��'������oګX�B�Cq"��z��!�4�#� ��	���	���� �����|�R�im�T��4^��ĉSw��Ci��? p��ɴ$��l��Φ�I�S��ZH���-ŵY��)6�O�5��'��6���~�]��j˻6�5�s�c�*l���<�'r��?�{��AưaR�߃-�P��*.D��agkNm9� �@h.��(���k��+�Opʓs&h�FR���	A��g�^�LxQ�E]�ɂP�L*d����'���'L��`M3m:T����4Q.�T>��5�ZT�h��
�	S��ӣ�1�����"Vpa ����3S(9B���?Q�AMKh ά��Z$����!`+���I��M����R�X�v��s��	1/S�]F��O����/2�<����<�l4Afx	a|�L6�� nX�U@��Pǐ���H ��n�P�>Ot�!1̦�Iğ��O��<s��'Tr�'�!#��2�R��3kLin<S�C����"ط�� ���3hF��'�ϿSC�V�s�:H�1��u�PH1��15״�ZԨG�/���R��#�J�/B�:�rX*���fV"EO`Pq6�ד$Jpl�bF ��?��O����O�8` �<D�ų���?]L,t��:Ot�$3�O���\)������O<0lж��9�HOʧkRD���GŐ���ڏt���2���?���+RN� ��?����?�ƻ�����O�p�@�WN+|���
������O����GvN%	f�']�L*�+�^2Ҙ����9��3�'�F=� A�~L�ϓ\b�J&��04��;W�ʷ<4�`���a�����et�V�f��Y�@�I_y�� ��� ���"}���Hӌ�y�nΟakT\�`�/K<�B�*�#=�/��O�.;6��@�O�\V�8[��І!򄜡g�~�K�
�� �F�hS*s	�
�'u �� *@ +2�Q��1��=�	�'���۳��)* 5�͚w�ba"
�'�x��D�� ̔e�@�Сk��a�'�0���Ц&_j���$@�ykP��'��LAh�#<���X�o���'�z�:�EzN~����)e�$��'�>x"�AU��HdN0ML����'�H�Xti�V�-Z3��/=)�|��'�|�¢@�J�dP��@��1c}K�'M��r��s����s|��	�'l8%��d�\������B-zȸS�'��pU���Lͤ��`�
w��"�'�N`7b��~y���8�X���'�� �Q��D��T+��`2�'�tY1��,D� D�6fȠp�X��'$^�W˄*th�$�g�X9Ԏ9��'7�)��tb�g����	�'At��`�Ћu'���SkZ�x0�'#�����fÊ���M/NGP�2�'��	���G- T��B�ބH�>a��'��l��aG+Z��ǢPG�T�
�'K�aE]�0Z��%�=Et0��
�'$쌢�H�j�ܙ�D��&��R
�']~��&μKZ:��&%�t��Y��'�d���F�P�qv	W�Y	*u��'�� ��Ը��$A5�T�{6:�:�'������ "�q e/�ׂٳ�'7P�H6 xp y��\�|��e��'�J��Qa�;�T�S痖��<!�'�b*҃\�Z���PwD�R  ���'t�m!W�X�s�Ե�f�K��x�'܄(�¶tE�a�f�� 9��(��'$R9�U�_M2Hآ�D>1 �	X	�'��)� ŔB>���ҹe@�d���R�RM+��?`�ɧ�S�3K�!+20��y�U��_�Ҹ+�H�}؂Us�O�x�Q�H;f\E�7��K��06"�,
d�dXedT����gϜ�(}fq�?)��C�azX��JG
p�5E�m����J�%ւ9P�+V�i�l��:X$.űGo���0����6�N��A�B<;tf�X�l��0JB��:~J��"�O�(���Vk>?��M�*�X8hg������P�_�<����rVj�a�'>����7����d�j�8"�ȇȓH��sE��;���B�/ϸ<���L*�a�@�$Th͓~�q)�z�%��jG���; �%��a�tEP�fުB�!���O�V�i�B	�?/.U���@�Oפ�n;O���s�S�^����E�Y�F�+gJ�{�>�\Ѳd�EP'�A++[�ĪE�.O��B#$�e�JX�&,G~��I6��4X~�� i[&/�٘v���m�a�@�J�d���*|Ov-J6��֕�#C/v�\�����)�O� ��}�viA�=QG�ƘV�t�ɵk�6���:O���@�φ�JOx�hZ�=��B�	�WHxkČÜU�<��v�`��Qx��wÄӾ9,ű��d����|���A*�ͻ\�2��+��B��(v��	�0Y��,�gt@����$G��d�Y�+�V�✡�i��;���qGם1����;��P���|2����F�6��K�H�ؘț�� BT��"�n����=��%��-T%ΨO�q�2H�!�.Ӈ�K"]Rt�`�ȇH��=�Ν"=��1򷍟FԞ]�@�̑jb�(з��O�xc@�ɅL���"��~ʟ�i�o�"OFu;�hĖv;a0㕟��r���mmv!�d�m������؊*���Vf���i>RA|+��ês�6�ڤ�ݥIF�!їb�<�8�b���~���O�a ��3T���0�
9Dw�ۂ�&��<A1�Z*ø��i6��	$~r�9V �P���ZÅ�.>?��ɹ#�2B��q������	\�rع�jJ�?���!��-`;�8Z�)}�K=@vms��4��@U��צ)"�K�y4dT��(ܠU��M���b.Q���CKV�x�XA�Ʉi����OTrphF��F��M02-]$�"<a�2��ĠP�O�L�'����@-W�B�V)G1m�|�2�AF�"Z���a*x$�
v�SQ*��=�Ә*}��O�w�h����Q$.�(��{��;�'"�d\�J>��/͛4~��I�x�D �!�p(Q	�/�䜡��	�����Re�c��=���h��6(<�y�#�Yt>��I�vojL�F��5xb�dC#��>NC��ˤi�F�%B��H�D�`�%<}2B4�S��@�t�"7-W�lF�xP��=S,���*zNrɊ���AE���7�B�>���w�*�[Ն��:´��@1�0�E�$���y��ߨ2�,��:�?��'�JvV���
SͺU+Di�6v3���6f	O~R�¨-lfE��e�2^?b�I���'/p:�O�C\�����Җ�y��y��6���ɳ�?9�G�ܦ����¶��>�c,Q�km�m�dY8NmڼP �=zF�͓h����H>����V�'V� ��)#?��b��
<6pD+�'�z�0v��R ���dWT8�L �c֠�|��%�64��i��$�f�eŗ;������@�l˺+�I_������\kd�)��R=����w�se�SI�|l1V�x��B�x2j�D���ɳe�<P*��~�˖7RG����CT�C�<�b�X=A�򼲢*G=�0<1��@���5����%�ׁ<T �#�مx~l�sF�Ɣ@x)�>j�}�g�x��*@��5�ǟ�6NH٦OL�NM�r�r���9IB���>A�h]7l󒅐���@���CN��%gN|��+X�d9�}#�I-j�Z	�;��I���"�Р�%O<���.����m)�P���2V�i5�����mB�%*�FJx"/O��y�$ث-f@��&ƋQ���2�A̛\˂��aX0�ʈ	M��;A\"���M�q/�I$1��OԜ�	�+�睔j��(��ҧn�����H�.m���B��-�V%�y�.P1c$ˋ羉15���Q�йo�
&剹Y$<���!���3��ժ3_ę�A�>�������� �ҳ7{H�ٔ Y{�'m�<�uM�b�2	����>R�6$BҦƣ{׾9Ce��)�`�#�0n��;5�����'�� �r��N[X�\�B�^�9�T��1?��9��,:?q����#��q��I��h]��'�A?�e��S��*�H%��x��%S��Xp�W"�y���7o#.�@l[;��<BtŒ�?N}�2��I6��1O��������,���w����ႌ �Xz>��N��!�D](@b��kgk�d�ru1CL��]TT�"
�<����vP�|�<!0*��--�aE���lm�=�b	3#M��J:���Ҏʣl��1E�DlL�i~F�"W䕟.��B ��x���z�k�2�����ާ�Qn�grN8V��yU���$�\�Pe�is"#��0�S-�82�i�G2�(y���Y2�f���gb�&d�֙� *X�T�:Q��$A�Hс/s��0�Ƅb�Q+��1���
�>A"�R)H�d�H���,pȘHaF�SDb���B@��@������O0�/%nn@��n�?Fy�A/\��O�)����݂0��?������ic�C�C&h��D�גJ��87gƈf�:`��8+d�,�"�H����kg�S@�'�h �G�6+>�$�Ϟ�Gr0�����<8@�fK]tq��8 ���yB�k��%�ǎ����������9��(u�R)��ȂF<(�Aդ��7���Qq�'���@��W>>��S�B}"iX ��/�yb�y�~�cP/��A`x�C��w~���U�)&�2I�wm���c�Ej,Cs�+u��-q�c�X�!So��r�^�;d�=/^�%��jҏx��m� BI��f����S"9���E�܆(`��o޼$��b¯8t�l�JY�GHf�C��Z,���A�J�J�u�L�'5�� �\��|�.ɗV��-ʟ'�P�)�2����#N�{�,ZB%ږe��˓x)Z��	�(ۖD��\�i���?i��	�/�YR����T[U�ԆZ�1�V�q�01u�O��LlΓo��XP�	�U�U���AA�o)f�tb�@�"\X�a��� 4t��pg�_&�)��	�_`�S���!8��:3#�0/`�P��{�<�g��7;�(��Ư�(���O^��觿kc� -�������v���x�	�x�����	HH֔s�	��==;�ġA�֤3�A�Gޘ��Pc��P�.��xbH��)��o��=���T�Z���h��M��ݒ���8�!��	D�b�I"��s \��/�O�"�ɛ`zp��IL:R �<٣�
k�Dy1�5�7"���Ӈ�Ґ %��>MՐ��<�Ѕ��Ew�"��U��xƭY�N��)�G�0�a@O�'\�D̓�� �
�8���ߕq`ǟ�&�l�BF�%.sJ1ө]9G��8k���$��P�6���Ҧ,��4|p�+�z�������!pv�]�E��<���;]\=B�o�w?��k2 !4�@�m�^�1��aۇI`��	J-��<��i˧h��I�Jo�? �}�ARF�ԁ8r�:�v���΅E��D�cW�I��:i�B�?Y�GaW?j`�]ZP���Y�9"�E�OR�}�� ���@�t	�/-��3�(�&3��D� �T�d�6iM�@�-����C����06�a�R�6;R2��EI]D�(���i�<Yn�UV�s�)J�X6���aV�[�i�W��r��Р%sʹZ��9�>����$�T؅*��]Fd�S��S� ��pH&�^� b���L>�?YUcV2R��TM,mKf�NɆ�f$!��݁UD�вl.za�m�'�?�O|�	�0�׎ �l],3YD kA/%�8��#d�.Y@�yB'EF8���w XiR���Wp-��'�;dZm���o��sq�'�ҽ!D��}HIu��Sp,������$�&	�e&ЙL��hЦ�O ��ɂL��\�s<�a�|�d�O$f�*La�g�%Ia�-N>
&�E ��6R�fyp�,<P��E��_�|��A>=�L� �LQ�15pD��7+����7�D- JWW�aأ}b�'(��HcÁ�G	~4(��&|D�a��J�t��y�V�6��LP�O>�џ �F�3&�,h��ޤF8�����)T�0a����?��Lh��P�8�>�u?�Oa���h�bO��pH�Q����"KC�(�K��	/G�xB�M�.��$&m޹��̓\$������=Y @8V���m^<�A�O���	ґ"]�L�f�,^�ISF�.���D28�Z�J�j��%@^ұOp��ϕJ���Tbу�(���'�d"+ ���gS�D�p��'�)��� V��8^ $��;^8���I�<ɡI�so�\rC�':��8R��\��2�n���|��u ��F���OU�N�{��a�9Se���Q�źc�A��6��4M@���?A�-ީD���0R�ޅ8b�U��-G[�,2�l+r�R<q^*�⒫p���S��SP��B�gźl6]�`��0~t��m$��xrE��6K�d���i��e��J<r����3q�k��R��~B?O��i�hH�="˓b zʟ. ���� i��hъL�n�`)�h����'��4�e)ҕB�H��T	v1�82��~b#��>Už|b�t,��p"�"v���Q�OXU��D�+��T��1��B�'��9J�j����,6��ʅ`�#~`��P�I5<� �Ú���]3��I����O�'�_�	-Q&� ����*�p���o{��(e��yA�8�ÓU[N�S�A?!�.͈��ԙ5��yZ��DE��Q��îL�\���O��'J:}ڑa��7c��rV:� 2nL�r��}R�JJ�}"�$T����� �y� �Z���3�U�y.�YAg������i/��q��
xc�A
���b>���`F�2�����=[r�a��0۱O�%�"�Ք]m�����KPld���=�4�de�z�/O� �"���عQ.� ]�ώ��*m>�x�'_�`"�$���-L�Y��_�f�rȂ��ՁcI�U�չ��t*�%��^b>Uj�Zs�C�'�����B6�� 7i��R~8Ey���?Z��aQ��Q-2v���I�L���KD�(Ց�`�+:�d�@��`�C?����V� {����}��&V &H<`�	[�ѹ2��`��IA�Y������=2t�I���j��9˅�P��$Ɋ{��H��$Ο��O���M�CNí%�>%ZeW�M�M���V��Op�p��M7�]��`Y��6�	0'���8<|��h`+�
.�m�CS��;}"/��J��i��ȣ�ۊ[�}@ 3D@9z0�k�	Z�Y X�4 ��sS��4���e�gy�O�xQa��v��L���Ƹj�<��5��d�=D��T	��,O�見Ic`l�F�R�>�"(��$^�n:��0�+�.��U��gyI�>	����Xyn��V��R��l�����P���@�&���dO���;B�εYd�S�K�	¼!�2.^?!7�0��cT�)��i��-� Ew>�p�$��H��%"O�U���Z�$,9Y���S��%�p"O�8p�
ʂ6�� �SBO+.�f@�""OE�!�� +Dc���5mѠw"Oh�Q!KF�D��f�[WH1��"OX]���G�9��Y��.��&[r��"O�0��O�l��P4K��+M̠��"O~0#&���(��P�Xl-��"O�X'ͮ/�(�ZT��:t�6"O<<����Q� � e�G�"d(؁�"O��#���Y�L�r&��tcnq�""O�� *B��9��I]�/_8P�"O�`�ӣ��<����H_�EI�� �"O�xfgH=8ْ�		��H�K?D����"�3�8��j�\隭�/?D��A!O8f�V8�H	�zf*��A�'D��y`*	�7s��K�����D��	'D�8�G�
��Ͳ�`�#��A
ǌ&D��P�߰6W.��.]7f��)p�%D���F�^K�@��Y<rP@��	#D��
p����t��!�J�Xp��&D�� ���jO�gbHUr!�H.(�dj�"O%R�ñkz�U1'n܉
��	W"O�	P��F&�p �$¨�W"O��V ��bj򅑲���2�"OPQ"6�W�������#�� �p"O���w*��R=
4`A�A�$�x�"O"��bc�`a�P�X�(p�"O,ss�
m�@}StA�'i�A�"Oxt�3�]C���T�ܦ9M�	�U"O�4P�0'����R�խ#�Hp��"O�ԫ�,�3U����Ǟ�&Z�l3�"O6�t��$s�0��fNV�^�b&"ORX����'��j�A��Jm)�"O�*d��8��Z���L}� �&"Oa�B����!j��Mo(�`�"Oveq�iԴ��M���S&L�2�"OgÆ�ِ��F$ c4"O�D��ĒY-�iSR�V0i'J(B"O $�)j2ZQ� �ȕ
���""O���0�%[5n���!,zd�J"Ob�s���S�v��4Ć/8�V�'"O�����,̰m��"�t�� Z�"OȜⶬI8C0Q�����2��u�g"Ot=˓�ϖ6�hi �fɓ	��L��"O��R��NZ\,CF:�t(2�"ObyѲ��q(��坒*�PY�"OJ1$�^�\��q�B�xup��"OxA�p�=!��5q'�&>f`x��"O�LiRǌ@���*rDU1oj�ds�"O0С�̃k�ܓ��.�ٸ�"O49��L>��jĨE6@�mɢ"OPme�3 $�k���!�<��"O�����A��tH��z�Is"Oqjc��(KU�,�t�·m�z�3"O��9��ܻjD�
�Ϳ$�D�F"O 0	`D�:*���&h���ޕ�"O
��b�:y��#'�_�����"O��!��X9")�B��,B��"Oz��VK�#iN��W�A@@�"Ov�����%>�U	"F�k��Y��"O.!���Y�cˬ!�r�߻!p	�2"O��{@cH�`���Q�@I�:fH,05"Od�`%
:�C�O��P��"OT;�Ę�l��D�c�U�p	R"O�����,PD"v��#�U�"OT� ̙X��=`a^w�p�"Ox-�����;}n�@��C�UZ�"OD1��R m��h��R�   "O����D
aN�E2vf�l�M"O�����$ô�J#H�1O����"Oh����7�X� b'_�)�浺�"Ob�c��?$Lh;���P(��1�"O�,[�'�4�fQ��%Miv�Z�"O��P���@��qK!cӋ �E�Q"O�,#�I[��e��b( ,���"O�����>d#B(��gQ/�Y��"O�t�GI�,e\3e�s�x�x�"O ��T!nI���)y�@�J%"O"AZ.��Hp> c�����` ��"O�h�(�,Z4b��'��-���`"O�Pà*�Z,J��ch�#X�>iX�"O�d	TT�I="5T�k�R��u"ONY @C�(ȱ'� [���q�"O�eH@��a�`9�2��.'�$�aR"O� �xy厉1nBڵ3f���Z��bD"O�ux"dԥO�hub'��7S���f"O����	фL3\)�6��*�f�h�"O�q�e�e'��v�	-�u"OT�j�)[:f����ѡH:\���K�"OH�s���!��-�+K�H؁�"O�DA�.�B���J݊:��*"O0$�W*��j�Y���'u&ժ�"O�����S�G�\��X9I��"O�XsQ�!w8�#c)�
Ֆ��"O�5�M�a���d�@5�v�	l��!%EҶL8DI�d��?O���5�3$���DI���� E7=��L��B�,�yƳ1�=Q�C�2KL�c�Y8�yR
� �
d��P+�&h��$Ø�yBk�e��*j��q�lt�H�9�'�ўb>�h��E}�\�R #(� ��#�;D���QI+�ycC��?R��T�k9D�8c�-�I7\��%EЩU4�ԉ�k8D�x�6ˇ����r��)=�"#��4D��PF�$_����F�F��Ĥ2D��X��K�W3��	s�H2WM
���/�Iq���u� ��@l�&��*g�MI�|��9�~�8EX�b��)�ƀ֖l+�P��Q��y�@�F���s!��2&�}�ȓ7�vdp6K��|RU��j��o�"%�ȓM��Up���:���N�>@X��%:�0��Qa~�p�\�"�J؅�U��b��S2L��&@��f�ȓ�ttȕc��1pVusb�Ǆbꔩ���g}���0��Y��F<hx�`"Ucύ�y�G��-6��ҳ	I�/?X�:�) ���'��$�����<��E<v\��R�]�}����"O�Tؗ`�=D�S�v�@�8�"�S��y��j_f�Z���jD��"���yK_�g�TI!�Խ{�(�����y�"ڂh��9Jq�F�nn���aMA��?i�'\��r�3e�����5��' <�(r��y0��l�ij���'Y����CA8W��+0�˥�pɲ
�'�.lb�� b�53b���!��k	�'V�\Bs��8V,F�r��vl4��'��,hD��[�~0@1�>n�Z,{�'�z��$ȍ
0X�pl7>�+�'��]yT�*�@�
q.6ꮙ�
�'�" ��K�ipa�(�OP�B�'�h܋f#��Q�:�i�j^S����	�'�������.s9T��mD�NV����'1d�ąJ WP�x6� �xH�0��y�iڄ1���s#��-�������'��{�B� jY����"�fl�B%	�y�/[�3�L��\��8��Ɨ�y�ꆄ8��و��©[�����Җ�y��@M� �ьX�"<�d��y��)�j����,�l�w/Ǆ�yRjBr��e剴�|��8�y2�L�.PT�j��]�k���GC"�y�e���ju���R���I
*�y"I�"�I2�υ.¬�&^��y��&f�����o�|P�h�=�y��![$*q #��j��Հw���y	S'9^��{�H.y/�MK���yO�V�ƍ�1�Z�]�Љ�!�
�y��N��`�!0�@�!ﰼ0��
7�y
� �ZDg��LyF��F�pE��"O�U���qx�sD��-�$̚�"O h�!��kn�`0c�?U.>Qӑ"O��*F�M���T�� <A!ca"O��c��(������C7�Jh�"O�D��& 9���!��A����"O�cAl×��xd	�� ����"OzT�!
Y ����ũC���"O@�!�\�j�"(��n:b��hy4*O�eې�B?��v�K� ��O������l
ve�2�J�<���sh��!�O8 �H�Y�|�; ,��6w��"O9+5�&a4�z�	�Pԁe"OB����X�1UPT�B�H�o�n]�'"O��/[9z{�u
3/L�^U�*O�3c��Z,�F��'ڼd��'6�H#���$W���ɡ�ɱ�:U�'z|"� �D߾њf(_i,\��'b���k�#Uʘ(� �^�P��0�'�,ɡS�T�t\a�E ��ڽ��'_}�Ƨ�@���N���)��'��� 'C��h֣�/K����'Z�cGK9��jt� ���"�'�"y��U&|���0��"�'U�Th߈9�8K���<�2"OnIs�7)�����Q������q�O��]�G��D8���l�:R� !��'���8�iX�~w��P����A��'W
�(v�Gb���Ƽ��'\:� AK�-)���aՉE2=��'�y��ũ�2Ai�6Ob~��'��Qz�/O;jMBѪ�JƝ2�����'�Ɲ0��u��p�Ů�/$��Y��'��m�aӞ�>��N=#)B� �'�b�bȐ�i`D�IG.nlɪ�'���ru���>��ŒƧ\�j�x�9�'�ڵcD�x܄�IQ�a$�Y�Op4Z�C�*3~h�#0K�! ��}z4�d.\O����;����!��"g"O���M�9d}!�L.,�xa�%"O(el�m@*����O7!朱q"Oj0�4�G�l��R�m(�॑|b�)�Ӝ=$��q���7���'�4	�B�	u��4J�葃h.\��&@�Z+�C�	��rL�� �`k*Yhpd�� �C�?&�p�����0b�����-rC�I�aH������5g�\`3��3�\C�əvmXD����4*��8�$�Q
^��C�	'C�`x�G�g��M�2Ώh�C��2RB������+6L"���J��B�	�51FA��P	>��P��E98�B�2Qj ����H���RT���B�	���	� G/�y2��V�V�fB䉫L���rɇ>FѲ�)�J|F^B�	�6K�)�W��D~��Ga :Q��B�I8��x�2��\$P�����x�B�	�E��-P���J� ���P�B9�B����A���ҟrʶ �Em�5��C�,/�Ȱc�+m��XR�^�9|�C�	�-����çP!��0��� BB�I$/D��5K�(j�✩��B�	<<(6��d��.8u.�![#Ay�B�	<@���:BHа>r�{��b��B䉰&Fh���`���J\�:+�B�)� x��ƫ�%�ڑ	 唗AՎ�ے"O����&?�R��'�A[�q�G"O.��E�ڧYm���°a[jaH"O����8vN���M�u5�<��"O�!�A�%}2��JQ/1н��"O���腯M�d���	� ��"O0 x��C�i�Q��M��@���0�"O�e���;��i`�N�Bܠ�##"O����N1!�ִh4@	!�6X
�"O�q�pcȫ6�h����.�X[C"O��������ꆏ�z׮ȳs"O���䁍F\H8�H�!�
�+W"O\���CO��*��ȯX���P"OD<*�mB!Ͼ5�P��#�8|��"OL��m�o�Ԥ˵�� cǢ�*�"O�E���.D�L�  "��,`1"OҘ�/̑A��YK�Z�e>A�g"O<Zr�	? "<Z���>^��zb"O�T� &�.ː���6Or�C"Or���#>_"���)Ȁ�B93"O����s��asÕ26��=�D"O�ѳ@�ϔ/~40
q#ƮBFT�+�"O��YO�]����0-��	:�D�!"O�K��e3�X��w3����"Oj�����Z�cƮU�$!���p"Oph!"K�d��������֜²"O�
G�)|!�Ƒ�F,��"O0U� ,���dP��!@��P�"O*Hi�L�[�r��p��b��B�"O��	!)�5}?��b�J�"/��x�A"O�ܓ�A[31Y�B"I�Va�E"O�0���M�=s�U���(�"O����
+��Ѡ�̈��"P"O�@����4�h�[�O�B��u"O
��M(_/Xp���(X"O���ꙊxӾ)�#�;=�l�rW"O\�#U�ā�j�)�H9C�C'"O�t�b�?H,�JVkI	9��m�"O`h�e�w��@٥K[7Tnv�S"O��1uIP1-�h'M*alt�hs"O�M����I�\���޿W.�x�"O���ӗ)�)?��Xq'ۦwG!���i��BL���*@���/[�!��E��-"��X1�,x��Fp!�D�+�\9�̳5����6lO�V!���#�nвP,�-�B��3j^,�!�ڜ.H�XbF�|m���S�F�W�!�D�Hذч� C�p9���đy�!�Ă�EA�D3�cW�w�8�t��g�!��+J��4��;QDr���nЙa!�,��0⬛#d��0�pT!��G���TY�˴U^*�H��a!�Dª���#�ė�iPx)�5Ξ�GT!�$�	*����N]�AA��3�͇$X!�D_:װ9��)��j��b����8�!�$�L��l��kG���H슂
4!�D��ߦp���8f�l�%�"t"!�W�
^Nm�蟩o�pM�kց!!�$C�����P+P'WK:T:B >j\!�D��9�6����"d��W��7>!�$އ6R�%���(<X���+�1>!�D��A�۪�PF_��k�ϸ
'!�$�_i�� W��x(x���D�-!�$<	�<�iG/�g�tQba��!�� ���V�ق"J��3������T"OX�je��jr�رpGݨ$؂���'t.QK��8$켉����M�]��'
f���$m�s�C�:	�X��'n(X��K- �vD�s�ȏ �*�d�<��")F�z=P���j>ms��N�<1�M��L����u�O�L)�� e�<���X5��Z�[
e+����@Z�<�D�3g
԰��_�Fm���O[�<Qt�2UP�@R���%t�A�`�M�<�w�oO���Q�I[TMB2hAD�<��͓�'�I���� ��S�W}�<�G��+fD�xvn±P��x��j	b�<!$i�
i�I�#�x砐�@��C��5*n���ՏoT���d��E*C�I"U"�|P��\�T�j`�1�ŁB��B�ɬh�8�
'�&"�r�r�O�$#"B�	2�.���J ��j����+u�<B�X��������)�T!��C�qj|C��<���b����`t��(mx$C�ɦ_|��C��P-3�4L�W��O��B�I"<�q;U
>�RHSIU
Kk�B�� b ����c�6\I�ťr?�B��;zd]��	W.���Dxq�B�I��|����YL���M�?�rB�	:w����@��N�(���j-\B䉥}��j�O$�"'
Q �,B�>'s�L��$x0D$�[ �B��=v�*�q�`�:[(� w�Y�q�C�O������(r�d ��\��B�I> �XA(��&1�;�m l��B�IXk(4��ۦ<�mj��Ԛ@�nB�9?O�$�b��`�NQ�.H�m�B�I:Ov=�� >���7��=tǀB��0N*y�/�eM���"� 2�vB��"d��!��
�tQ�b��f?$B�	�p��5`Ə�\��*��K�u �C䉩:����=���@�Յw�C�	���<��EF8{����0$S>w�C�I�	�5)q.ה3L�:6�Զ��B��6}�j��fI�٪�Q��2T�C�	���1rbG�N�v-r!��?LC�C��2ri��s�����*���.�pC䉆v1fa�h^(Y�<=Å&�u�<C�I���4���DO�.���H�	q%C�I�Mt"X����Y���!���B�	3\��Dh�	�m�5�ad Y��B�I�v8p�"�(
=&/X�C�
;��B�iif��\/�)y'��5���R"Oإ�u�6�bQj�F�OPn-y"O�$����+Rvx����!��y��"O�D��	B�|�.H�NL�w�,�"O��Q��
j`�� 4Lt�W"O���*2?�)Sc��V��t��"O:�` ��+C��8w*��R�"O@C���*VTXi�C�����KA�<�G���S�D13�Klh���@S�<�K'[�<|�v���^`N���#KM�<!@�[o/r�u�=4�R9�˅G�<��.E�$�F;�%Ϡi�x�)�B�<i��Z�Ct�� ��]��u���@�<1��=~a\�ڐg
-xV�a�k{�<qu�L6m>��P)] `��M�<Ĥ����wLW��(+1��O�<� ~]Y@N����P��C��P
"O��s��0�(Г'H��k�|YB"O�"�#�>*���Fl��SA"O��A��Ƃ��%�����R"OA" FU"
.�1dɍ�?��i�B"O��;���R�$�+SIQ�5�\pc@"O\0�A,V��|��h�1eE���"O@t�C���&��V�Z�r�"O����h�� i �жٚFў�p�"Ol]��� �Fe���Q*��p"O �3DtZL��B��K�4 "O 	;vχm��\��'W�(�H�"O�Ir�4]�Iu�ށ%Ƶ� "O����6~���ȵ�P������"O2X���P�;�vA!�M�>�\y "OZxAbaJ/��y�U�&��i�"O\��"<N����b�?AGv�b�"O�1��@��z��A`��@.��"Or�f�d`z��d.�>F��5"OjH0WI�+�j�┬��w!�e;�"O�E9R�ǆe�(!B�yf�s�"O�8�ƢA�Nрeȡp�*���"O���L�*�X��C�B�]��c`"O�<�M����l`G�� ���!�"Oj��d咜*�2t;C��6�(�v"O��fA���0�	��ŕ�6���"O�\[���:b|�`��L�!%��L��"O.���Β�P����E=s(8�"ON pÄ1E-*�Eɱ_�B���"O<�
����T+u�+��H�"O��#�XO��)I�̥>�
4`F"O\���j5`�2���#�o�P�"Oˤ��MT���"�3���� "O©�bᝆ/ �b�׻�dXQ!"O�" #Ļ>hR�f�
"�(D�r"O�`HÍ�0o�~��Q��*߼5!�"O��C0/S�w���ڔn�v��"O�s2K��y��l���A�A>�D�R"O��C�54���q��"$,fQ�Q"O|�����?��(D��T ��"O�@9֌>a��U��IP�hŀ"Oj���/Y�����RX��`"OVU�e	S-p��;�愗6'��"OJh�n�#tP�KP�O�8X�3�"OX�ѫ��e�� G�ebN�yB"O�yg��%Y��US�&P�Z�
=��"O�m#�bBn~y:��κ`�ԉr"O����#�t��Q��*�:G�x���"O*�a�űa��c�gH���#�"O�lxe�;�p����07�mC"O�|Y��#ӰI�Qe��\J���"O����:'PFhRFٟH�X��2"O���E�u��aJ�C�1`p� u"O�#�E�+�h�V�ӃQ2�X�"Op�s d�q��ӣ��	��y"O��8THC;E�J)Cd,H�M��6"O��p�a��H�q��� ��"O6��슨q�0	�h+O����"OHi�A�0Q�ĭ`a�V)xT#!"O�y�fH�>qt��x�G҇�|� "OtIR�@�2���ɱ%��X)�q"O��R�ѹ]f���� �"O�還��<��#֡Z7����"O���5D�1Qe�&.0��W"O� B�
��[�b����ղn�+�"OJ�35��&M���S B�g��p6"O
� �B['R�E�b�
�OU>�0	�'�0��%/�� h@P�3Z( ��'�DHb��4j�8@�g��a 	�'c<-P�UD�����+B S��Y:�'B���!�)a>� ��3C	p��'�*(�e��T
LӳE҉z4���'B�a*��G<M�u�W�9H6Y��'��u�ͫp)��Y'my[p�z�'�$·��>C��1���+ *��8�'��1H�m��5�|��Vo�7�a��'�hi����� �RY[��@5e`��A�'����Ge^�i&�)pHǤ+�}
�'������E�M!�T�e���+5v��	�'z�k����~覨0$��vI*�'M��[��%QKl;3O&$�<�
�'�=Zai�	 pB�I����(�
�'��@�J4]�~\�a��ݦ��	�'4�\0Q	,q�4�KQ��=t���'*2$�d aU�*�H8����'��T	˖�4]�uÉe��I��'���Q'�
�`W
���ȟa�dՊ�')" 6o	�gO�<As�J;Rb��'��Y�R_�0�(������'���š¡���r �n̨K�'$�tIt-ȟ+~P��-B.^/0��'�t%�0LJ*D�8�hV�J����'+�]q0B	�Z��D�(<J�X��'p<
���1�1����D-Ɯ�'J����k�`�^�?��a �'9r���T&bP�V��6�z}��'�(�aG��N}��9���7N
�8�'o��&��E���+�mϥ2'����'K�<�%I��e��{�C�.���'l��Y��:o�٫c�\��	�'OZd+"�<M`�ۗ�TE���'Y,a��J�4q�x*7IN&�~��'|��Q���9W�>�{���..����'٢�����V�E �
�8	�P 
�'�t	�I\"&��qG?p6��	�'d��^�~5�� *<����p�<q�Р�R�fM��*Ӯ�0-5D����E���h��t��3��q*�#2D��k-�O=��	 %Ρ,4��V�/D�0�H�^�M����!>�Z��1D�@��g�#t犱B�	KL��'�3D�d���Ԣ�i#&M�OF� ��2D�D���$ܜ��l	-��b��1D�`���~x(�����/U����@f1D��Q7 ��8 ���X����2�-D����M�����pV�p�D3��*D��ⰋD�S�  	���؜"�I%D�R�A�b���MНd�=�w�5D�Ȁb�F$Q�,�$H�>04��C��/D�H��(��I��u3&��x�4�+"D�\�FOK�7<�aN'��x ��<D���f�S(Ᾱ���
=��P�>D�T�U,S3_��A��2��%iю=D��:D�Ӝ$��@%Aț�e��b8D�P/�L(�%c��>%�l ��٠"fC�	���T"���d�$Q����TC��
�\���f�-��l4�Вwp�C䉏=�h�2(I��0��Z�&��C�)� @�Ȃ) ɐт��	�4`�0p�"O$�%C	 ��}�P�G���)R"O|������@�h#���N��""O�t�dG�aOb������ɣ"O�0S�N�c��hr�M5@��Cg"Od}ʐM*o��$is�T0ԅi�"O��7H3�T�:�jq����"Ot���(=�����T�\� y�A"O�l2e�a0摢�GМ/�ꌂ�"O"��)JA���QU斪%�驤"O��k#9k,t�eЅd9�Mx"Or��	�.m�q�����m8�١"O�ZA-6������N#�q1g"O�	IF �
Q��	"M� �d��"OVfD���#1kA;rB�3�"OX�d�$R�]ұ� H��"O�J�B	�l04��'�/AK�	�"O8
� 2;�a�ŭ��6Ke�"O�����+�d:E-Ц}��]�#"O��!&�ۇzX�y�,�
��"O��`ЦS(B�AbeÄ�H�c�"O��	��v�Ve��cÑLƦ�"O�h!�!�X�%�B������"O8��4h�)�<Ի@ѻ3��"O���C�����A"a �h�9�"OJ�8�Sak"L��ƴk�|͋"Ob%�.�\�����0x�ɛT"O��yPᕓ ��)�Q/J���S�"O��5�߹n�.	yt��9��9Ce"O�BDL�%�
����R�vN����"O�����>x�"k=$�
�"O�t�"�Hݞ�2�J�, (HHPE"O~u��@A0*ڔS�邥cu�ك"O���֤9�^�)G��?���S�"O�cv%�}���ӷf��ё�"Oa�wm/0�z!�-2��a��"O� b�lۻDֽ��%
�P�p�q"Or詵(N+-@��Ǥ�7�f��"O^Ё�K�<~���%2)�Z�"O�1ҡ�\&0̼�[�d����x�"O�ejU���\�fՁ1F=�(lhS"O�p�@�X�lp���b��`�  ��"Ov �@:^$l Ă�(0�$��"O:hX�	
�\؞t{�G+|ؐ0�e"O��S5i��x� ;%�
�V��l��"O��P�J�)�|����ۍ-�%a"O.pX@�#�pܘ��B�<ʤ)�"O@2"+�a��@��K�_��Ѻ�"O�����ᆹ4a�p�<!6"O�Jኋ��:yң%�'S�<�
�"O�D��<�c��D�gPذZ�"O��آ�Z7v(��"�d$��"O���a��#m���#a^�l�bg"O:԰3�w=&��.��
�޾�ybI�y#����K�?Ǥ��6��$�yB)�;4~�ň�hU�/�B�4�y�	�����ᇶp(�i[0���yBmO7<�t
!
�z��x7����y�������h�����)��yr��"K���V��B����4�y��L�?��IhT�0�E�u�އ�yB�ڛ���%ÁiW�x��1�y��C+�ZEQ��_c ������yB�Swyl���#�P� ]�%d�y
� p�V�v�5�	H���"O�+F�p喝Zק�V{>d2"O��"ō����H0�O�2oy0m0�"OTH�E��:f�1���K�5�Q"O(�9��14<D,A����y�n�sW"O����@�:u�B��ѩj�}X�"OZ�$']	,��q0ᗽ_r����"O�e�V�� E�b@^�7"O ��%^;q>�(FFGb�E(�"O����fWoX�\�w*X�"ΑpV"O��1��t�>01��P#(p�a�"O��{�d��+6��$E���"O�-�#5V�<Lcĩ
�Q�zM�"O0�EB֤	f�@9GH~�$4A�"O&H{��C�PO\|*�GH3�
���"O�a(�Þ�x�&�&�o���"O��S�Ťd��`$�R4�|Ȕ"OJ��F��y�&lcգM
*1p$ c"O,c4�PdH��fE˵l�N��1"O��pb.R��=a�dT8T��8�U"O@a���^D:eAm�(1I`"OR�(��dQ���A�����yr�M�@�F|��gۅ&]�؀���y"��)I���H��C� ���� ��/�y���]�P�&G�� �����ybe�����p-�x$JЎҴp!�d*�HAPD$d�0����:S!� �n,�"爤���r���B"O������,����(��nu�u"O<���T�Qzn��,T�e����"O\���ÍM�0L#���=�t 2"O�()�)��I��1ԇ\5S�"OD�A2+J�7��S�N�p�T"O�0�F�={lX��@�+���r"Op��еK|��j�EǺi 
�y�"O����<D��⢊�F�LE�"O��{th�E����A���X"On$�r��43��d#��9"�M�V"O��g�С��4�7n���<2`"OV�z������R��R�(fiB�"O�u��)OZ�ĥa��4NU�yӁ"O�hX Er��I*��@�G�>q٣"O^�i4c̄V�xȻ�J 2t���"O���$ئCi�M�D�\���"Ob�p!��;נI8�*�4�i�D"Oh�9V+_�'��{�D�"+�f�	"O���5�;,5�0��T�@�E"O��Z���2E��j�:4�ʕ(C"OF���m�,)�4�tj4�Ä"OF���(R�i@��a��E2d"OF(�B׮8 K"O'jhC&%"�y�� 
-n��6��=p�Ҵ1f�Q�y���W�0��i�#l���"�E8�yRDگe��H�k�^9L�)�[�y�)ǧo���p��?��A7���y�X0}�x}�䏙�K�(@��y2�
�U"8��� H+`�2u�V�y��%W0E@WE�P����?�y�hI,?��j��\����4�yb+t� Eq�B�>O$4��LV?�y���A��AthG�|���+DB���yB���$�>I��]7},���c��y!��F7�E���q��Tjc�]��y�������"�A�W�F¥��y
� �90���"�9DjH�
K0�)�"O̜�%hJ?����5^8�3"Oh��L��΂\��\�ri�F"O\�S�!X�3�rx����*�<���"O�����4%�}�wh��Q�\�"O�aH�N�Ԡ�A�DV%�h	d"O�A(�C)`6r]iʓ!J�I%"O^ ���) ��4dhŹ`�C"ONp[��=fV�l�'�����&"O�!�I* 5�+q%�<R�h9�"Ox�r� F�,� ���N'N��P"O�,xp`�XD�ۂ�Gn�x�Yg"O&<��Y�<�v��R�������"O�M"�b�צ�"��mHX��"O����-
e�P[��/; 	yu"Oj,X�����t���c 0lp[E"O �Q��)��zAB��{�5%"O�ez�L�u疽3d_8��4B�"O�H��ᔍ�8[�b�fu�h6"O�JBG�1��\��
K�ib��B�"O�%��	�rB�{��޹@��(y�"OXB��߿#WXT�6�c��Y�"O�ib��MgN��#�AHv�:`"O�qUG���db��
pV� �"Oв� �BtA'��Â�C�G!��!s1�͏m���" 
֒�!�Յx�\�*�G)hb�yʰ��<[�!�D��E�h��C�Ui`�xa��p�!�� �84癹r^Pp��ED�0k!��Ax�t� ��B�ƌS�C�
�!�d�?Frʑ��N�	4�j�ۀ-m!�¦1�%A�o�'>���AE�Wi!�d�.3�(���[c,��S���F�!���t*B���%N~�|���V�h�!�$Wd�lQv�U�v,,Q�É�!�E:�n:W�Mb�x�u�30�!�6P�dX6�)><`̪�A�,M�!���;�Ph�E�֕G�����<m�!�$A����"���k��R�L�C�	�.rb�x�iZ.N �Bb�K>T^�B�	.h��Ԣk�"yf����mH�
��B�	84�&C&��,�n��kȕ,Z|C�I�Fkv	BWI��z�:)�F�ŧ|&B�ɕh�N�CG��0,��RiC$�C�I"��e��T�60�S̈́6���IP����l����[{r(�b�iS�`���A�5D��P�#w�xx�f�Q9Iʠ1` 5D��"�b&P�h��O�(Qb����3D�йF�!i\�t���L�HNLy�*O@��Ej�Iuҕ{U��)�] "O���V��$~���B�,`Z��"O�I��@$�0m��D�x0ؼ�q"O��0MR;&��݊��={M�D�3"OvL��O݋AE\E2A�<v�P�"b"O2\���À_���SkX��|� "Ont"�kS'�ʽ�r/G�t�ȹ`v"O���ǀD��Zh���T��E��"Onlb�(Y�6�A��؀n��"O؈���?I>��2�ds���"O�pяY/ZF�����O���1"O|�� ��tt��#!ΝM�4�"O�!� �,Q���JG�^>p��Pp"OZ5p�@�OE����"�:�	"O����2H�&����[7"�4Q¤"O� ���F-M�8��I�8v�y�%"O@
�gL'������D�n[�l�"O�I�/��A�Z�Y,i���r�"Op��28�3��|�nX�p"O�u� �G	νY!�T�M�rHSP"O^A�V�˘u0zY��,��rY�@n"O�}�"hɃfsv�{�!C�#�<��w"Oh��� ȉ(a�R���"s.܅k�O� *F(��\q�s�+]BL�J��O*B��=>����_�Cx����,�B�ɸNo�X�$�E�@v(Rơ��|��B�I�}� �W(-j0�$�ƈRcpB�	�c�����%s孲W�9c\�	�'��C&HB� �$�ևD�T~�-��'F����N>d�\h�փ�Y��!�'a��� ��=97�� ��^��~�S�'�D�� G[�gEL}�e+�$J����'�X�C�+�7k�Z}�u��;yO��;�'���17�.~6^�,�u�:�2
�'�N����S>���F�-q΢t�'W�x� (}k��Z&fb� ��'�ũ�ȃ���<1e���a�<��'���*&F�3<\ �k�W�Q
�'6N��g^�l�/�N���b�'`���#O�;Wh�����B!:zf<�
�'�F4R1�.�d��r��7m�x:
�'&m�$��J��P�G�S�&�H(k
�'&!+�.�������vux	�'Ͷ����׎{��Ѹ7�X�t����'�E���[�$BǁJ1I��!��'�6(�7�<��VIG�1�'�������2�͊a���2�'����\R��M�'��']�l��'����V�A�`��x·�"	L��	�'�"d
3ȃ�;KP�bW5DX s	�'B��VE $Fռ����@	z��l��'WA
�\ 3�f��#;`M܈@D"O(�ȗ,
�|@d-��$@*�w"O葲����L���bɢO>�C5"ONH��C�;��� $ζ#.8h"O<]�n�
?���v�U��̘�"O�At�X�k�4h ��)-�n��7"O���O�2FA�䓷��%{t�"O�)�R
�/d��Tj��es�uzG�' ��ȟ�G{J?�[�nV�q3�(Y1"�C����&b=D�<��hW�A7�|x��3*{D}Ba�5D��u<�vea,�/2���5D�T��*���1f#4aU6�c�'D�ظG�H>w�"���♼y���ǀ0D���bh�>(2�4:�eE�8�H�@"-D�(���LO�r��b-*�zh�	 D��ڢJJ/�ra�~���f��y���*'��L�t���jK�1����y�f�/%��U����Pi 1��F��y��D���A��M�>�pt��y���7%P�iц��Bw�r���y�,o�����ڨ7�"hH$�y�$S�s��X�-�pY�����yb�.�UQfe�3!��a��`���y�阚Q�f}#��� �舳��W��y"d�p�%흗z>i0`
��yB��?)zƕ`�b��6�p{F��y�
Z�����	Yt.)�._��y"-�NH I�Pā�'E"l�%���y
� �Qf�	�]����2�HIr "O�}ȱ��"~���XWE��Sڌ�҇"O����Y]{�Ր���;����"O���%ѭ����F�׊h�h�w"Oԍ���I� ������Af@�R "O �@��*��F/@	;j���"O2���f�Ѳ�o��_�պ""O�t��[��d��c� 6P�h"O���O�B�X�bD�F'$P���|��i>h�ʍ֟�&ě$c���AVb��z+��ʅm�s�<�瀼/fn�[��!�.�z�+�n�<��!Z=)����1N�"EE@J`)�s�<���*�p0���I'��F�o�<��m�.7��Q�G%һT�hiD�e�<�q���\Ҭ��n:}��q�A{�<�)ұx��"V�E6��hƬ�x��~���O���3q�SX�plC���U�Z�'�$�(	"���%�Y:����'2�{�`�%}�j�J�L�9�
�'��ysE�Y(���cD
�DBЀ��'16��w%��A�#Iwh�Bf	r�<QǪC�Z�@�M�5n��s/[S�<��,6;H���Ԇ[�\���F]I�<Q'�Ėb*�!�F�G��B�m�<q7K���Բ��τ���a��e�<��Y�[M�`RbF�:�qᨆd�<�3GQj��a;ѭS�"iY�E�<!�+�+����	
�����W�<�Ө[�2�:Hs�c�k0��Pŋ}�<���D�I����塈�i���iK}�<a�i�~�T���#� x�T`�Rn�<A�厄ka��ZF)J�LȖu
B�l�<��
,&]8hCĥZ��ȹ�s�a�<�rN��BK�)��	��$N�p�u�ȓg#�qAD�;���{�iR�x-�U��#�!�V��DE�y;������$Z2���� ��c��χT^� �ȓb�%��ꔣVB|cd��* "��ȓ:  K�:*�jDcD�%+���ȓ~�X�a`��� { ꀍV��T�ȓ8B��a���#��-����S��E�ȓY�B� ��FjJ��ǃ�/�:=�ȓX
�("c��&�n(���ٺi�V�ȓ,r�ѳ�EP���!_9K��!�ȓ=�*�;��������4�� �ȓjM`@�S�N�c�e�\�!�ȓ7��5R���<��ĭ�-n*~U��D��.�=��$�G�V,RT.ф�utp���N�;��A���! !�$B x?ƴR��w6����'?!�'Iei�Ҁo2}4#U5!�Իh�@�b@À�t�1��f3!�L�S��s�$�Y&�E�-!�DLW�m�E��� ����&Z0�!�$B�~�p�(ą��2?H#e$��H�!�Ȟ<�Lٲm�7�*5�7c�5g�!�҉>���B�mF���:�B���Py2�U�H���Ǌ�=�:T�!��y"Ń�Ī#��2vD��QR��y����J���ra�s�БV�J��yH��3�Ƽ����y)�8!�
�yb,E8<�X,�ŭ�bF����y�j�>
����	š##�]������yR�Ġ""��&C�
R:�@h4�N��y
� �D��� ?|�+��Ӑg�z���"O~��AW	\M���"X��Ř"O�yW�@-p��E�G��h3�"O\h  �6eW>X���V[���"OlY��
�"�e�_(*C��$"Of�A�]�i���K�3?l���"O�)��Bˍ+Ƹ�0��	2<-��"O��ce
(�;�D��%�U�1"Ox�B�р[]�È)c����"O	p�H��$�p莾-�b$k�"Od�cA��# :�1V�
h��	"OF��C��%*=3�e������@"O�ա� �x]��DKi�xY�"O��8r��)|��r�̗2�Pc"Oz��LA�D"v⛤�P`�"Op�����Q1��b�@L9�(�CG"O�D02�ߨm�N�`��Czv8r"O���s)��A�ub�:��,Z5"O:@@;����� <kf���"OT�:��H'~6����iS?f�@��"O$�3���:�.tS��q~�(��"O�E��!�I�M0ˑ�'��mS�"O�;�Ȏ(>�A���=��ɺ"O�,6A�����S��M,ֈ-��"Oy����(vg"��س.`l;�"O�e�Ι*3�<0�	�!\���"O��`��B6b.b}�ӈ�z�\�ѐ"O쑁�	>2op�h�ᗅ5��#"O�0iWB�d�!3O�Xq�r"ON�J4�ێ@����!�G g�4"OHp"�Z"���K��ɿO���i"O�L!bBJ>~���Uΐ�j���
�"O�xr���^t�h��O4]�c"O�ɲ���=�����጗5xf�yE"OFD�R1J��`?�9�%"O6"�L�=e�(3m�%> �ۅ"O��)K�)r<cu��$*��"O6q�F�!��,��3pH�"O��Est(��L�
���"O�q�C����J K�H��;�"Od���A9q��@����;�>��"O�;s�1z��(�ЊJVXJ�"O�Ƀ�N]m�j��V�[*�
G"O��z!��<<�-ST#T���f"O&���hʴ
v�������C"O$��&��%*Ȃ ��l��]�f���"O	��m²Ll�*Є����"O���e�͏f���TI���L�R"O^��!��!&���$�#��		�"ONac�g�$u�˵K�h���"O��@�Ǝv���#祓I L�s"O^�P�N]�\�͓sE=(.�uxg"O���`+��7E^��E�X8����"O6hP�$~��� �z�V�y�"O
yam�N���$_�\s���"O���� ��L����E�d\x0��"O�hrOGq�}��-[*^?f��"O��AE ++����clN�?L�b"O,)���B�x�@�%�[4��"O~IHf�ÝpR����7%x
2"Oj��5�6;��ӂ��<$�م"OXu�-��`��iB����+�)��"O�X{�%��3!Z���gD^����"O�LCE� 4�;�F�T{���S�? �a�A��F]�y3�&A��a6"O6�0%˕5+@ȓ���(4!�!W"OvE�C�3��l*��˂I	�d�"O|[�"�=.�&�Z�[$	�L��"Oj�V��2!� �飦�%v���"OD
�J�#��\�����%�q"Ov��3"�(q�]`�S��4"OrذRM�U�ΝR�H��@^9�"Of�{A����xq���A�B=Rj!�S�3�X(���J�Ydf܍iU!��O2N����)���)Vf-S-!�D�N�L��G��f�{e��0!�ğ�6�l�2�&<��<��j�>^|!��K	0B�bA��q����<)N!��%	�ի����z#�eh��M<!��T)
/|�Ps�J$
P@�5��V(!�$<YxyK�Ub��yFf�.1!��4n*�:����Jh����߬
!�$�d�puA��P!����ĢE�!��X6ez��-��(Y�C/�@!򤐉4����W�f�s��ӺH!�
�D�H��6I������л�!�K����ڱ��8��E�cόr!�$�x��h:a R�c�f����	�+!��B"CIt�{ED�$�����m(l�!��ܥq��i�RJ
k���JVl->�!��]e"�S�T7g��-�w�ۭ4�!�d[�s��QA#F����]q�I�!��2D��0rD@ �<�F����DP!�So-�QuH�"i0�!D�?!��K%�Q�,J�{p�K D��%�!�7g_��{w�T>f�s�b�	�!��8loޖ
03�r`"ˊ|9���'5�Q[c��>N�܁@��|f� ��'y��6n�[5���H�r�t] �'?��Ҷ$�-�jT���X�r��PJ�'�P�I� 
�䬐����x5��'[�X�1i�g7���̈́M�L��'��m��卶n�
 � d�
@ʂ�`�'/�4P5&�aDy����4�>� �';.\ ��9`>�9���ٵ.��I�'�.0z�������fS�W� qs�'��&"/HŰ�$P�8�
��'���n$V�0�Ι8A/����'/����n�(d͜�RJ�";�Rp
�'�μsT�%��0�a�Η`?ܸ��'ytYv&׌3��I)A(�k�|��'��q���+M��x�p�4y��1�'���R�-P3T���I��L�n;�,��'J-)���
�]𷃍k�1�'Q�=*$��xnU���j�+6D����/F�H�����m�Xq"8D�`�j6P�b�IC�L�Q2pM#D��c)ϡ6	���M��@Y��� D�l8�hO�bo�pH�33
���&?D���҅B
��8�S�H2_�P�A)(D�ģ��ͣj��\��.E,ss4ġ&D�8gHP"<��hR���3D���0D��j%�״z��=S�[-4����J.D����C<k4D���ivP[�k D���-�i�&�·�٘R�l�#4�"D�XI#GJRN.�yw�����a�a�>D��r�kCT|ذ�ˬ@;�5���7D��*V��p�8ApB��2���!D�� ��� o�6l�䘣�G	},��"O�L
2�ػ�l��H�&�\�W"O�LZS�[�k0�\	6�A�,i!�"OX�6��R�^�va�"+$dab"O&��狒!.��qQ�� 	�,�pt"O�]�'��F7D�j��3(�(���"O
��R�3�4���1l��x0$"OP���B�P�,����2]O|C2"O��#
�&}�$�S�6֠Uzw"O<M�Q�p��Z�#Y�x&��"O܅��f�u���jrW�r��dZC"O�8z�/��gt���C�@6��uA"OBSi9%�Ȅ"�<9}Jt��"O��
0�߈������@�"O��BF�V�M�h􇇗^���*O.͘ e��� r�`d��'��X�ǚ�c$��k�F��i�L�
�'ص�ؤ_�nӥ�U�fp��	�'9X-`�E%&:t��%ռ`�J�"�'��D��+Յ]�R�����9&	LyQ�'� 	���-q��}����	g
�0�' �� �MQ9(bn<{$蒺+��R�'��Zf�H�v�͚��\&m��,B�'�d|;�0|:ܨ�S�R<1�L�
�'�N,[A��-P^���F7H,��'��b�<��83�"�t��')�UR Ǖ�v�^������Q�'��q�qR�tR�t�=�J�h	�'�t�`��
|2��R����0�j�'�@u���p���ݠy66 ��'R����R* �&�q��'�
�z��Q�;����4�޹�'A\��G%#��+q�Ȝ
h�S�'[d��A(Y�C����q��8��
�'��x��3N��}�F⎜hƩ�'m ��Pl%u�#V�\-Tyq��'ߖͣj�}�X���M�6<5�ɲ�'���(�(�'#�6@��ߴGN�,{�'8U��h�<�7�h}(�r�'Ő|j�-ʙ3� ��閝����'S�����[+X�DԺAMI2�=�
�'�|��w�[+V��䂵s@Ȉ
�'��*���8;br���/wP���'�,��tL�4��!�l�l���		�'������+4��#P���'h��F���ta�B\i�	�'}�P�-S�8�� ��DF��8�'�L��,�*'�8�hpB�IK�$��'c�4B��όD�!! ���t���'GLL�G#��P�1ǉی
0�i�'6
D�t��A�V͠U�3Vup���'��t��#Ҍ�0q��ѩK����'�Ν� e
�wR$���EWc�-Y�'�pMajD�:��Bh�7nR���'�)'�:h���s��&,����'��y�Á�?��d��Y��q�'�HV��l�	��D��=�D���*D��H��
(����H��[~��GG+D�0��ǌ[�\�1dE��)��j<D�|���@&R3DQ��b�n�zV)/D�,`2fޕ/c�h���]�|+6%%�,D�X�Ɖd�*|�@�+9���!�I/D�t�v�R���w�X,,9|�hq#/D����[A��z��:c�zQ���8D�� ���q1G�p�a��#�ȹ��"O�k�j�-O�LIf�è�����"O>�r��a�a �(�+eR֔��"O���E&\�V&LzA��Ok��&"O
�JuQ�z�����l8l8"O����Q������ ~ �I!"O��7�+S�<q3��R:8/�6"O��R��(�Z8�C	�U-R�I'"O�'Fw>� ���CrH"OJy��f�\z��RS�_Ȱ8�"O�M�婔�"!8�qЙf"O�h��+e]~�rGo]� #�l�S"O��m��\U�;��̯y0!*"O&��F���$-|��(j�"OJd���x50��*�7��uR�"O��r��@��TR�HF%0�2���"O��s�oo�R���)���9""O����D�� HI* ���yS"O �7$^K.�,P����"��(y"O��� )@�|~���WC.|H�"Ot���V"c_"��oܡ:,ti�"Ox����	/>�*8C����/�4�P"O�����U�9 �`&��#/�Lj"O�uH��(�VPY���>)��U�"O���͖p���R�6�8��D"OH2Fo99�䅻7k�.�jl�7"O�M�#�4�TX�'�X3$5f݋�"Od������9,xp�
-���#"OB$�M�>>�Z	��``dt}�"O~  �V�b��m٣Ҿ��d�c"O�Yǎ+� ���L�GgH�"O���j�)��|RG/S(g�v��s"Oz���9�J����FD��#"OZ�k�:Uy�h��n�9*-���P"O~�@�`�^�x�P��0�ѹ�"O|�!D��M�~i�3�o���XW"Otl�5�A�]��}��ϛ�u���7"O�Mjw��k`XD!ʮug`@�`"Ot�kĹA�d����Jq����"O*`)!�M�f�:P��?��%A1"O�����t��Q9�9����"O�l("c˒~J����U�?��U�$"OF!�g�U3Tc��C��L�`�"O�Q;����~Y���Y��D�"O�0ё��/x�Lu�T T�l�BQkr"O^!�I^>w=�-�V�Qz;\!`U"OH���Q3AV�U�%�U�n0����"O�9�õ�Dq	��א.f�S"O�x��-�U�y G^1�l]��'�.䩵+@�C�dhd-"�ڹ3�'jҝ�@g�w6,�D�ܓ�|ɹ�'�v�3���0�Đ�ΐ�h��R�'�6��Ή�d)l0#��dl ��'��c�.8v��!�=_]�h�'e�Y��K�C���XB
c�.���'��@r
ُ@�-bV�B�S�h��'����󧊿3��Bu�M��A��B�<	@l�%3 ��(�L��b��0�D�@�<)bQ'�$�x����;��E���Yd�<��.�	D��q �����ċ�f�<Y��D�#E  *���ogL�6/Em�<qF瞈�|l����ZO�AF��q�<���{���c@dΝ]4��ûw�<�&K�.�D$;#՘BS�9A�L�<� �	��g�=hvҁ�
�`*�U�R"O�pp�M�6����S��bL�"O$P1�����Ç��3�,BB"O��K��>q�e�Ԁ#%CN��0"O�$�X� ��}��@@k��i�'"ONYP��OR��q!a]7�h]�2"Oz��6 6���+dKS�L�Ll�D"O� b5`�!rmƘ�j[�bU�9��D0��)�'S�X)���]C���4���ȓqO��ѧ@S�-�<��L�@@X��%�tec*�`6�d�[y*Z}��v��5�o��`4��+q�S:b��=�ȓI2�\34�B�c�DI��f�x+�y�ȓHQ�����A򈆄���ȓ,+ �6%H�Pb�[�������ȓ]:T� g�0�L
e�#*��ȓ����hR~F$��]�
����Y�.ay��"{� �B�9,`Ї��G�'�L��fP�a D��i��a(�'n��k�w���Fh�2����O�x$Ў"��)1�P������"Oz�Q,�+w�(]0��V��@!��D#|O��KD��8�ȓ���f�08���]x��k@�4�ڨ����.,PD�*D��@��+�Vj\*/PI-$���$0?�-ٖ(��IǪ^�oX�(*V�c��E{bM���c�
�� i!qKW��y�b$4�e��(�tyP���y®���̐�or� <�J�-��'0�	r�O��ɩLE',80!V��l'���fh֣�yB!�l,� �k�9x�,P�@���y��)��-����h�eJ�
o��<I�,D�	�!�OFq���Ŋk�����%���f��L*�`�3]:iSe���B��H��&6�O��j��)# !	�.B���bhU�$O�L�� ��ؘp ш(��dH#*��G�* �OV�Dz�Oo�Ie&�'�S{�h[�'�?D6�͓��	p���q�=2@A$"�U@d�9SO-�I: �Z��$�!��8�`+àR����@� ���$�_�x��W� �J�n}كl �ഊ��9}��Y��4�0Ǖ�P �����<���Ĝ�O`�q*C1dsbd��� 2�$``"O$e؀���M����0`���Ւx�BLl��(��5�$MP�F��F�p�0`�"O�)p��1:�M	�G�vU2���"O
�ta߆���jd��6�,���"O��a���4�l�� �e��AQ�'3b�=���(OX!8��E�Z�%#���0XF���u�'��c���< ��@�@�!��Y�"	�'7!�dN#"Լ�֠��N��x��	�����D�De�.Z"�O�vmA�-�y��.,O���"ۗwJ^L���@3��=xr"Oze�bf�{(�=0��Ԟ80�*OЅJ�+_5���k���=���	�'�rLY��Y�&���oOe�	�'`QG.S 3{�$��ÖV�F���'8�11�����h��Ğ��ı�'��p@��a�"M)�J�7���I�'J�žp��@�a��'� )�ķiLfu����-�q�'1��5�����q�J� OA����B�)�4��D��"�(~6u2De�#�y�cH�M��D�O�o����b �)�ybaͳ[�U0�kQ 1[d�qL,�Mcu+�0�?	/O��G��t�? d�J*P<  ��Z�=?| "Oh20h]#
l�;&��*#�d��"O�M`�ᐤV�	�R�ޓu��T[�"O$b��J�T��@�Ǉ�@�����hO���3W|С9��Y�Eab�`GF�=5�!�$�`�Y�P��|h�/�=H?!���:��e �F�,��4�g�;�!��-_�$ �č-BL��%��!��5H,t(S���[��Ay�mS+y���⟠Җ�D1ʓ������Z�g.6�!��Z&��ȓ��ɧ.B��jLiV��{�̕Ex��)B��N�V��hB�W0��Ls�+�X�<RB�4_X ���=�( [�N�<Q�n�"&��!��O%2�f�ga�'�?��b哶*��ȶ��6����m�ԇ�	�oSdU���VL��� �P�T6�C�In�z� �>n�ǮN�x�DC�	:@�@XZӇ�*)@� "��oV~��{}Ҙx�Y�4$��ݖ������H�$aj�b�[�C�	�s�3���MqLɣ6�η\����`؟ܸ�eA%=sK[zv"e�3�H>OBџ�D����4e���w��7- �f�h�J	�'�}�m�b3"�F�"�X�O�z-O�ҧH�M��˧uD��3f @�"O��Z��̞P\�@䄓�{3��3��B���I�9��wFط[���vOұ;!�D3<lD@6m��l�P�(O��=E����V}pp��7�0Q3%���y�BǇ!�TU���-?��������y��|2�'�*� q�#�^����U0<|  ���Mh�d�ju�!��h�HH�T�w�!��	=��+���$Ep(Te��֒>Y��<%>c��ْ�2S�U��"�|��s�>D���b@5D��H�+\�H;�,B��<ɏ��&u�V����ٛpv��H̟8�nC�I8�djs.� (k��!ň"AL7-[���?Y��8P4n@�GIѕE��X�5��c�'C�'�r��|�D ,5
���m7 ��yD�b�<�s�
(�t9ⶌ�1�V(zU��_؞`�=��b˶>H*�X@�z�����/�[�<1�i�p�@�x��� (��`a	W�<��!
�HA�9���P�P܂L #�M�<Y�� d��,��-D	5bJ(�"MVJ�	]8� ȅ����.XHFj����9A��#D��͖C�
D��
��o�����!D���h�D��`��A����r�s����0�)��]y4I�d2Vu+��@�N��"��1D���&��C4��#��Y0kkp,���+D�8�7�ؼl�
��2�C&�TH�2�+�OԒO�D�"�����r�Źd~��E���b�'U�����7:p�c�&��x�h(I����	"w��9be�Q�_�T�h�l �v��C�	������
?���Y4�\���O�˓��S����Bӎz���@�ېc:����u�0���7J�D���
[�b���h��t��)�tK��#�Ǝxhj)FzR�' ��j2�\�+�>�2C�\�߲�YCO�x:7��;Jεz��*���:1"OF�r�HϦV1�;�ޛeN�\�O��Y\H<��bˁ�:,,T�B�Id����'���� �GBG�$aP� EGD|r`"O�ܪ�[�VQ��5 D�a��"O�p��n�Q��p���aJF Q �D,���$�	+�`��Z�g�i�c�ƛ&&!�� Ԙ���C�찹�&W��]���	ix���2�E�7hy��(@3i���B;D�|�e�շ%��M����qM��Z�3D��Ӄ�V�2!F�Z��R0����0D�Hs$gԑqzLj ��Y\�Ha�.D�h��-��U4h4fL7	������/D��J�ܘ$b���J�rT�R�a;D�pi���p��yꁇ��./\(���5D�8مl� t�@��&��i����&D��`܍f�]k�b�8O���SE(D��3s��J���f��rz9{Џ:D��v�Xot��&� (�PpRa&D��AT�r�J��&N��ZMyB@9D�l
QC�r_D��p�ͨ�V5���5D��D�*�Z�����8�$݉�#0D�h	�K�!|bحh#��.�$Aj�I8D�Dɂ���8t�U��&=HB�/5D�xc�e�v�Z�Чf�$)���+4�4D�H�R��h����%&�R21D��0e*-+n�K���/�R+�O+D��)��P�~eʧ���1֐����'D���uP�:�t�w�	/FŲ�s�e*D���aI��a��(0%�L�ؔ�=D��£@�8�&d�5eF~�Y��n<D�\sWNQ�Qæ���C�:XZu�R�;D�#��ȼg����ݞJ�\b�o:D�H�ˎ�S���@GK�\f�聃�"D���f�4sp���[�Zkʐ�%�?D�|!��#%v6����Y�<��H���>D�4�GD�L�����
�Բ��8D��DB�v�BM���6�����;D��Ȣ�ճ7|��DÚ'/�*�3$ ;D�X�2�QG�q[0ᗈmW��g7D��	'nT7��8(�J֢v��� ��3D�)��)��$6`�6��@���<D���QFG�ZN� ���F�U�7D���ӥ�@�����MX>�8�0�"9D�����!�r�h��
4  �"�+D��ʧb��U#�eK���[..D�L�%��&��A
�IK�erB'�O,=AQ���f�@$`�X�&L�u�-��:�"O��E��?b�#"G��h�s0"O�	rPF��	��Pb�_�i�z�"Ox��F���DJ�@K>t�^b"O�1a�ѥW�j0C��J��J�"O� v���,=�n۹E���Y#"O���U��AbЬ�͆���]�!"O�����@13,^i����j�"O��#IV�� $��x���2�"O��1i	-%��P`������"O�Z�	םkA���Dھ.�0��"O� xG��F*� BdO�k���9E"O�=!g��-+�\H�t$ �o��c"Oꌠ���F ����h�^� B"O�e�b��}c�P���"�\X�"O��vOs� � R@�<��uj�"O�p�r N�(�e�&$þ AʝkS"O�	�c��e�F�Q�ؕDMnśD"O��#IS�;�( t�ԩ
q�0"O�U�Gʚ;�Ĳ���	�@��R"O�Y��I� f�Hj�b������"O����d	=���0E���%-���|cz���%+���,���C�V�O��U��8	hB�əe�\�ƪ8��al��vR,���̪��0H��A��S�? &����@�4ja,ъP��� �'�,�U��%B��L���G?mY �/�
I��xJ|����4��ZR�H�b��x��7
�<Y�ǀ������ �1��$�Ɂ�\�zEy��5nxz�7E�?�!�D����Η�T���H���Q9��O�U�l�E�E�<�)��0�6���|o�H�ěv����`>D�(F'�����!��U�P���߁cu�e	AI��|6�`I}���3�ur��sY9L����@L6zS ����b�X(��4O�h�W�j���I�/Z)8��RU�ǵrm�xТ�
|ܶ�� ݮ�p?� �Q;+&�|/i�܄s'�acB��{��'�͸�M̌�	�
�۲���d�!�<j7٥Dd�8�iC'g�v;����y�C
>mV!{�`E=f���_7r>���S&T1  D�#���+K��y#���5y�^�c�NE�珻����	%�~�Y�mлn��ڣ�.�	�A�^��q�)P�U|z��#�n�2 .����F�+H)@��(O���a�ߒT��I	ՉD�v��fh#?�aP�̇-oǪi��S�4�"	�%�_�C�z��V�:����A�t��֌��-M6�Z�M�X��bt�F�k�X����A���� H��mk�aψ6���?�:=�M�%	���\Iɒ�R�dx:!,/���{aU��8�zEJG&1��r�ٽHaJ��ӭV�nh*џ���I�n9A閌Yی� Bg�#3���H�K�nnA`���0|�Ǝ�.\���
W8��y�*	m���(�"+���PE�IR���̧\��XQ3��9�I�l���"���Q3�؀��Z5*���ŗ�.����e�Ȓс̯+�Zl.�+�1���a��=z����F�K�?����'�Ħ+���Hn�m6�l���>x5Dp��+�U����V����/_�<��+rr�@`��dJJXK�aU7���Y0I�$4
��p�$5��$�?�� pv#��ހ}p�� uw\�c�̓c?���BƐ'�l�d��A{�����,A(`Q�l
C������O��2�b����D�_tz�u7H��B4\���3EPn�am���p1���7*;����E��l�.�d�#æf�����y��E�<�@HD'�0_O�	AT�F��X6�G���sF��;'���@��|�#Av�r!W��<-束%������:tnF�;����*���	+�r��ջe�<)��{>�ʠh�8qb\�CL�*���Bx������7���H�7M���\݊Q�ؚ|�a(�I�?>�(O��������"@��V�=��*!���<]ܙ�� G�up��ci!�$ǐp~���)��h7��r� �C,Ru6��#��7R�"ػr��z��ݻf�(8�nYEH}yb�ڴ �������� b���!�&ryvT�QhB4�<��fh��DyGƷ�0c�i���������HJ�j\;��cbK�C���yg�@w�
isBď�&�,��l^�r��Ig(��?E��';��c3��`J��2�K��ʔa�ãI?2[*}`�dX�P��H#a�%>:��ScB��Z%��6��A�w�4@%f�>Qc�83�� Kfl��'9�*#Ę�M hrU̓N* (҃Bj��2����y��(��4�؜Y�c�f��G(�g8x���̛6��Q��`���6f4[��^ C4���3(4p�s!�³#��#� ��'��(�c�:!z��CF?�<k����&<�%�SeߚpePk��̷M.�Y�%Z�O\�!fE1�����K��`H:���D���R<�3�>sɲlkSυ�+
`D�9�X�S'lJ43�J`�A��D���<p̴h���s�B-��g��0qJr�HF.�ϟ��B.؜p���>E���+<���QΔ, �u����-*�r#ɹ�T�" �Y1�lx �O=���.���Y�ec��~��ϭ7�npQEF�t}��2a�A-��ɮ#��)u����%��^D���X�k�F��2�&���b�S��I�v���*��}@lޚ&�	p	Y��Oh�r�ǹ(��ہk�Wn���D+3hma1C��O4�q���Z�,�Z��V�?`p�DI̟zH�!���/a{����V%��ܑ�d�B���j�U��I������0��/uINU)�ۓAz�0�q�[;t�n��+�}c(O;rAW ̼�Q ]�9cL�i��[�Va�C"��J�<Q�/0z�� �۝}c���rS�,<����!���'�Ȋ-y��Q��C�y�<���ڟyj����gI��?qF�V
D���r���|F�H�˂Z���c��<�Z��a�1~�B��'�K�~utE�@A��l��öh�{�L��gVFP��N�h����*Qў��K����T� kA:�� �C(�Ɏ;�� ��/��裁m�����c��<\�0�R�J�<�V���[�Q��!��
5r񤹚�JD)*�������s&AUn纝���U�����	�`L��[8[�z+��ظ�����h묵�+F2U��;VzР�O�*�@�b�WK�مȓ�h$�O�iv�`�N�u��|�@J�;�e��Ǎ���HW
��b8��/Єo`� q-��q��H鐺i�\����N�j�2���<TH82���j�����V��5<P@ 2�~�dK�U���Q�](R@#���v�����~Aq�Áo��	1��pϮ�S���f�&,���&$���	4=�&��q�K>aWRH���ߞ?�vL�3H�F��FE*���n��8�2��$��e_Np�2�=�bd��HS7`ʐ����&�L��g�<&.@kvlX	���x���FK"����ށ�!f��_}� 9䎎8]�L��`�΁q��=�LE����ŎL�8P�I�#]~��(�u����AH�"iC�+O-th�w���(`Rx�1,7]XN�OPp�q���^_@MȤ�7y��ѣB���\i�Ņ��O/p�^�*�i��W��e('ϒ�UcF�R�'�Xa��u��y�ɐ�b�"�Y�N�T��iw���}oZ�J��A�rK�D��i�5��
t���*�)��d	$)�4^�-y@�FI��M�B�F��}�e@�	rذ�Z)�F���# �|*�$k�W8]Y$���E;5x��"�e	h��EÊ*�V�Gy�.'+�0�F�_�X��B��:3�b�M!�v��5j��z5	'��(��#%d�
��P���xp�I
0R�xaA��	>ށ��⚈Wo�	�V�N6�Ո��		:ҡ�G��Rc�9���O��� v�������P�ORF��t�D,����$z�IJR�>E�Oڰ Q�NSr��7I"t{�`b��
sv��s�IK�3���$����!�H<ɇ�PNJ	+�a�y�&]�����y��$�T1`��g�Z��8ajܴI}���S�ρ��YXQ�i$N��&i�|r`�a �R8"إ���9k����g�� .��=լ�p�e]�P)BU���w�����-ۍ0P�:��!RO�l3_�����ǚ-� 8@*�(&o��t/i�f`E]�pњ�X��ͅ4#�%	U#]�mY�-� ��D`ےQ7�%D}�E�L��i�GG	�Β�k�6.�H���&{q�0J�̩<�¥&r���i"H�3$�6�[�yT�l�4�ʜ�.���K3�p�Ƒ
/�ay�K^�e0t�&��R�q����� �:4���cA���XK���A΃�G��͈�N�2�������;�"�Jĭ��[��
^D����.C�A�xq�7��~�����(K�p�nOV9Ss�QR���Z��-�R�C��3xM!�Ο,B����/;��q�f,�G����� M��F��M���(O��pMNK���!��6m�j��<� g��h��&(�|��"�X�!f� ���L���)�L��p��e��8�
$-�l��RM�8	X�!Q*�1r���D�(���PQ��)CwJ�D^lٱ�	^x�,de��mS
�~.0 q��CRP����7r� �هC�`q6q(�O�Y[j��?��BQZ���D%Hb����C���m;�&�k��D�����W��5+Sc$-$�a 38CE�"�tA��G"�
�.�
2�F�P2�F��?�!OX 0許sK�� �z,E�F���9i���-M:h�'�ֆK|�!�$c"�%?�x�Q�ȡ}߀E)��>h�0P��l�'�8�M��J,�'�ϏXr�Q[.hJTm	�y21':D����.�p��ܟ�qO|]y+ҺmW����OP�4��D�W�v�.����� �IS�̄!�~Y�;H�M���þB~��#a�<]R��*Ǟ�O���i��4|ST���.A�fx�I�4��d?�M�'e��	�0��I�c��}�E,��28��)e�*'���b�L���)�B��ðl�6�V	��ؘ:��UKu6o��j@a�LF5
��S���,h��,�p=��"�63	^�����l���M]�OTDX�s��"w��aV�
����4�At*)��ď76�!���~�����#-N�ҺoD�Y(tE��q�@��g��P��}�'Q�.��&DS�G��$���>H3R�P���{*]D�L�04�t�U�'���@�B���0Ó�J0P�H�iH�x �Dݽ`dTq�� g ,�Ѓ8���h�n���	H?�����΅`�����p�jᧄ#:�^min=g���kǭvZ��h���3殜�r�~�*���;K�Ls0�ɯ/�Ā�.K�3u,���ʀ5Ē��2O����X��úI� DS`,�-+�ШCq�1p"��T���91�Y��$B�`K��
�ѓ��.�x��D�4Gcn�xʏ6^�c�abNx+��Ѫ� ��8Gn�(�@D�Dd~�0�Mˌ7^�$A��g�.	o�6�qq��h9�]�t ��ha|�%>����b�T k�C��t � �r^���E0v>7m�",nҐ��m,�Pf�F X��Bע��i���O Lqe^7~IZ�
0�U�"%��	$%=L Є��?k���� ��Vm�DH'��!ƁӇih�)aLV�Q�(=X�.��d$I�F���|�K/ C�V�q!D�'�J̐�/�}u⨋� ק���+`̄�Z�e����9Nf]����8�^��Oڅ~}�����z���S���_��A�i�Dp@5��
HE��8c�؆T��MX$�'�X�
x��䣓#��2�2@@ѩ@�v��ā��?>Z�3���hbߴ9���Ǉk�M� 2��k�i ����lN967�i'�'q̥�ả�W�ށ��X�q��#\�
l�v�C�I�,�ŇݑTQ8�����k� ��$A]t�5����_�x����O҆�6v�|�d�K� Bp��@�Y%�O�9��L�h�l�j`���H��z��N����.� f�j�)v��p�t�c J�@�>16M��dM�AKLF�?�TK�+`��lh�	b"�x��O�?�����玆WIJ�`�"
�<�`Ż��ݾ*t�H(�䔈`'�X�3�V=9����(!��ՙ�!^�L�{&	G�2�sg��*��ڤ�'~�0 ��� j��D�$$��S&�Ac�
�N!�f��OB��#%�3t� X ��"m��p��dʹW.�y�w�d��*��f�V|�t�P�(`
�Cof<���H�8�-�2f�q�%۶c�7*�L�hŁ)l�!Jg�Ѳm9�H��+ċu�B4�R�� r��#�5.�F�P�Oƭ#B�!5L�I��愝���.q�qO����e�waJ|�&ɳJ�ʼ�Ө�
Pd��Ƅ�,�BU9w��)X����o��jn`��B*U�w�.���̌4�-��&6�/�V	Y�!�D���	�#�r�ɳ	W�!��
=pl�lzbh��9�d)r��X�%�H�3�F�& �f��c���$ʘ�Sf�����}���Ĭ6�v���׼d�Q��������B�J�,ZyR��l���k5�A��s�+�y�`����8P0�0���V��8J�獗i�Ґ[e���
�� Cu�!�y�nȯ��͚@N��.VB�g!�I��a���q딕@�N(ҧv@t��CC�;��!��B�QyM�g�ڿ<9B=(��� �ig��|ܠ���#U6��yq
Tse��-����g�	i�!%�X�=�X�k!�W�|�����'�����\	]���M4���r����
�΅�_���"b
��Y����K	����qED��𠕯	/5,��H/�RN ��*����'2�"����~�"H�7Vx��-Y2Z^L�'h�*$�Ay#%�%}ь��d>�*�HQ3_l�'-�VF`駈]>k̩x��+"�$ꗽ.�����܋ٴL�=i3NE�hS�tq! �'U��y�ׇ߇7��s@��">�+�	�%~��1��P����π3u�ڗ�����_�Tѭ�e� ��\��0���^�D����"U�\ 1� �aD�\��O���	��r9{B��X�~Uh��ѫj+��h ��?��K��|��B���ii����m�p�W��+T�N���&A�G ��f�x�����Uja ���$Ëe�d��47��&*V�:�Z��ɗ�,w���A��b�f��*�o�`���ǈ]%+�U�BD����>L���`E��#�2	��X!�~�K���6��$2�O�z��mI���8`2<<*
 '�>��y"JJ�$�*#����M欙���1	n��'�ͲV�`�W�����	s Wz��$c)@�O����!Iۺ����!3�Fq Y�WXJ�s���	����Q 7��1!%�վu^�c�49ue�<qT�QS1@^+K[X��YW�4�"C"�p�Hel��AI�(PI�!�ݱ4��
'�, qD<��Ч��Ke`� ZB�� x4pvcì_�%�Gn��6�eʖ^��� ��>vrh%�q-�7v8,�1AW�	��k7������>��<!q�_�c��x׍��n#L�ѳ+�I�r�`�r�\���D>��09A�ߩb��H�mT�m&D��ûie�������� '�
'N�P�&O(Ҏ��) (~�(�pŉ g��U�|"�E�F���e˵��t�M�.�Zs�*VL�l�`��$��rA �#1mX�:e��4��l�=9��C��2���k{@@ǥV�X�M�,Q�p(��gD�wTA�ˀ����jGkzBhEхT� Xᭀ/T�`���&�A�~M�5�P	��#N�9KdL%9T�7�IRJ��eɖ�FԂF�⨃�nS#)���C`�WԾ��G	�/jϘ� ��>�`ae��8�t�l�*�ם8QLq�B.����$$�R=��o��.X�x�DD�/�v�'\����H�g]X钴Dҫc��ApaE
k���h.�$�!�'Z|xT�C-�Aiu� y�Y����B7����W4&#}��wZ�h�4
�j���P���R�H�o�D�`�d�T���zu7�� �U0V��eF�{��,M3�ă7�ܥ^z��BF��v�8��d�=z��I��Gn>#>����Dj���"���
�0�2��&
���@ߤL`����:��y�H¯F
y���H6bH �-ǜWx\�1��P(Y��LxPCFs�p���`а�\&�� P��Վ�������%b[�������5B�3@��D-�)c��t���Az�V�cv�Ǿ��OL+���	���?��%U�w�r���{m�u���ޣ�yB+9���� �K�C$��MY!��/69������)�'\N�ѷ-[#l��5j�QBć�798PK�O�+TB4
�)Ӭ$���=ф)֒Y����$#B��	�	N(><����8�!�
I|��2�=ut%�q�=z�!�ď�>��a��M�#���;��֐�!�Һj��թd��Y�*��W�A�3�!�$H�'/�P��NԊ/��VT-R����ȓr��e�A�D�D�V�� n�21�츆�oN��R���NND�:�G�2ߒ��ȓ$�(5��F��U�,Hwg֧| ��ȓX�P5��b]<hMP�S�8SD݄�=�����U�U�r�ӵ��-�����Ԡ�>@u e3�Я "쁄ȓ/%0�h#�F�!��Ĳri�*8���I��"d,B%K���FǕ�P�*p�ȓ!fn�0��0�4�0�W����H�|��cX.'�<�H&�_������>US��K�\����R�K����H�=�$l�)���`F�M�U3��ȓ0L�'�>A���W�D�T�2��ȓAF�QCi[�v(������ņ�[4p8Q�ڈH�xh� !Q.�:��ȓ�*T8�͌�H�4X�!� b-��5o�8ӫ�X�]�U�51&H��	�|���=C�L�pGΔ	bڠ�ȓs��8��'��`�Z"�DI�]�ȓ��}C�ܼ| N`����E���ȓnF �J��,9�LP QGR�p�����v�J��ʄ�y����p� ��TW���5�b��2v�/K�R�@�"O�lc�[�H�MҥOE�J�̼�`"O�)�d��$I�ҙ�a�٭8`z�U"O���fEC�$E:A-E:>�4!�w"O��vG�rD���J�*R���f"OZ1 G+ZaJ�K��C(?X�+7"O�%�A�,��X+Gg"7U��b1"O�Y�V�.;@^ ��f�02�Jdɤ"OV���lC]e��1��X�u�,�q"O���bCD?_$�p�WJ��C��(��"Ox��fʞ�.;b)�V�Y!*���"O�m�$�ƖK�6XZ1H�"���!�"O�� ��J!A�&�qŇA-=�� ��"OŠ�щs�h���e?[�b��"O�)hSl;K�9a�a�[�<��G"O4��R�"ǼL�Bϗ�>��"O@�!AfB�d�n���,k�jl{7"O����JC6J�^�ǁ�9�E�""O� P��nGP'|��2��_�6�D"O���#'T�%�� ��dXs�O=�Bm	�!���O�>(E�
$C�����Ě7;�(��3D�xfK�h�����x����<Y2�Wp�U��0<i������e^�8��I�ƕpX����ͪc(����,z0p,k��2
Lb��Ų�'M@�!���H[��`g&�B�ȍ�	]IJ��m[�K]��@G!��_�-�$��H� � ��C�4S�!�䊕c�� ��	������UA�'��P!�k�!<�y	`
]�Z�9�)�矨KX����ӂ�n���q*z|!��2�V�҅�P�h�8�K�@��1)J�-_mUY�����`0�<���b�@�-%�m�C�@Vci)�e1��2�B���+3����hՉ �����Ȁ�.�m�f/�/���2Ŏ(+��
��v�Xhw��8�ddb�bZ}�V��ɅwŌ���.�&(�����]�, � N�w9���@Et�da�#=C @t���g�~�;T���!�]�d�ޭ���L�Р��`�>h��Yaf�\�I�d��(��rTj�4���S�.�8j�ʒP���	�l���X��@�zz֡:#�XM�㞘�rl	�f����{�i�{�҉`��5b�(�٧�Q��������M�f�S�;�`�cBuɺd����"<	S��j�����\�J�Q�'A$F�����Z�N+ȓO���c Z�J#��Q �$}PRt-�=8�հ$�F�Sw��iT&Ɨn(BMx$��.C�~D%��[��� [�-�V��H?y���w.|h������AL�'	z0 Qٸ
g�����t2�˄�ފ����B|��8��y��F2��)a�N�U|t5�t�M��~�		s����k��!l���ӌi�"�I�I��A�K2dȈf`�+0E�d�t�@�9Nܙt#f>�:��I4M�4��aH6fĈv��-2Lh�a��E05��>GJ�z���$�1h	>, ~�-xn-��?I��ˁ~���e h.}k��ͺOO��e���"N��F�g�ڠۤd�![�&tIpb�m"}c���:LH��%N�qf�51<��ӂB�d���P��z(8dBc�.-\	�)O���	6������ow>T"G�����(/7Wݲ�r����6i`��ɥA<`c�m�����̓�'ʘ���6T٠�"QmТ�&qH�<O��7p��A@6;��aKN�&K8��30' �NP��虴`�d��4x�@��� mu�Ο�nM�IF���W�N�`������PnZ� 5�Œ	�.���'���$��\�65���V�ND�; @�kmXM�\�z�� �	��7ӎрt
�� Mbh�p]�|z#͘I�D��D�� �%C�� 92��!�R�ȿ����g�R��	oZ�GW.���?V+���JU;dl�cTU������(P抅���n �Y�՝/�@Dj���5J���ٶ`�X�5K���& �`H��ҩD%�`H����h h�s�E�V|�����ąu�6�E��9�J�P��_jy�CT�Q_�Xs�#Ԝ{�n�*a��'޺y7R@���Z��y)��M�Uq乫��&( >I�(��Q}�@hu�;���x$r��T�?�]��mÇĘ!L��Q��^47"^��A!7xA�1�D�����A�)��<�â	0뀴�Co�;A�-[��M"=+� !�	8;�"�+$��3$�0��'芨����G����1dmΨ��C7O���B�a�\?yCƍ�o�Y��ǖP�b�P��'�	\�<��E��o�����iR0!��oZ�9A�@m�1�*ejf��2|�tؓ�J g�Q�O6X���Iɤ9��A�5���Y�,~&㔣޼��Éy�Þ=�
����#-��Q�B'�2K5�����dz�b^�4A�GB�z�<�0���C(���o3��ŃE�Z,�+ߧ)�J�>��R���Z幱�1R�Ҽ�A�?,�"#��Tw4s�N�(~Kʕt��hdj��9��2��y��ѻЮ�$��|ƒ�b�@N��?!!�jKt��G9}���D&Y, q��W�k^�b��T<G�PQ�!�#�`��^�j��U>C�J��&�t��v��FP�+��Of�0��
_	�Sf�*\��YRw�>��LT�c�֝V���$�U�K�A��n��d�&��@ HK����<�"f,ӏ�4��K�|�u�C���j~�bC�� �p:	ށdv�㞘�4o 38ˊAhs#י�d, V��M�8�c,��324]�c ӊc����P밬�p-R;:�(�ؔ�˅�J
xJ����\)Ҏ��M��Xค�g���e֡j�	/�M�7k�
�Bq�M9R"���wp�5�����] �E"b���'O��H6�N�Yu��W�fԩ)5��c��̉e'�d"����UO��`F��\����&
l��A��'VqY�H�p;�)�AΝ�)�	�@ð���݀��ʠ]5�eq�� ��B��K)-�����Z�L(��.�,A����r逝Y<�I��D��`)~M�GJv�L�+�K�8�1OH���=�ެS6�5r��)7�?��x�s)�:f$��c�N^Vq����_$a���2f�>3���IU'
IX������Rs٨c��A��hQ%썎z���C�Ǒ9��YD(Q�����ɟ<T|��Ӏ�E��lAumޥ" �'.��x#���d��H %+&D�""#��w��Yed

i�¸B'�@#%<X�wlћU@�����+u^*rÔ�r��1�$�j�̘���M� �4?�ii@��]� 9ksЅ�jA����D�х�36Q�0[?1�U�,@�����Z��р���0xPY���v�0�2b��<=@G�':a�q9���$[R��A`��HOB�{ƨڠ3Dfxc��3�!��A9g��	2cF�7��=�0!� _V�#f(Z�0@p\##�0�5�%E�c��d �.��h	LQ��q��!�b
�v�V��Ơ�u�'��ya�F�9^��ka%�sㆀ�0��Vڴ�%ѰZ�x���`$Q��Y %�ů�_��4D.��)#K�b��=�p�ܑ1�TX �^.5@�ZAG�]��y9Ę|RE_��WŢ"���g��^�a�ץj[=B!8,D��U�]���T�a�P&!p���d�^�����/O��Uj2�ƛ,F��J�=��@�Q�"b��r�� ��S��Pm��x�#VQ�0�0*]?e�&�%<8r�!�oB���cрДl��l�S�V�S�<� Jܽ8���-t���3bB�6�dX��n^�'�=!"�t�@N�q	4�Ȇ�5�l
�XEi�l��Tb "�~1��(�S��i����"I*�5H�V���x�	ڴh�1����Ob	�0hA�T�&��ND1H���J� o�^mi7�R�2�N�t(=�I���
 `�i�FA	�Ɠ�4℁k���[&��u̘���T(Q�����%�/XÀ)SQm�� ̎�U8�E�X���th�Y�Ĭ�0%h��~�^�CG+Z�0}����x��5i�I$�����o	r�|i��G��L!J��1��СC�<X�L�C�,_'�m��4;j��gkX)<�t���kĹIv��!��{����>X�D�I7� ��c*38TA�!��1�eè<<���Xs�@1��`#Z2���
��64|	���8��.�"pt�x&��� 
�2�Q�W+�;���Ч��J��1#��>��YҘ���KF����͕-���YP�ɘn�t,��_��bֆ �#i��⑤G?:f���R�����ݱ�`H��&�Kd,�r�ӧİ<��	͏9��tpUJ��I�Ε[f \"0�0DP̒<=w<��!nͼy�)��BB�8�3��ȋ��#1�*|(��'q6����?~�B�))j�P�BزF}�X��D�d��'��d���Z����s����@L,��.�������Q(`@t�zx���L�sd��V@]�MS��,w����	�x���PH_���J'ϙX̓�T#��'2����r�F=  K77�fIB�ʂ$:<�rǪ� �D���%7�� XB��q�H!��~)V��ਚ
R�F4��+°7�h��Ǣ�	���x�NE�n�$��I/��Ę� �%3
6Y��f�$I���Ɍ	6���$�J3�����Yȇ�F� ��,�M������`��\�v3��Ueσ/�ɐ�.AN��Ժ�gaA��qj ��12�Դ��ݱy�m� �ŷO�T$;�N�*�	�G���^@�4�а�`�O0a���ڥR"��i�.QPf]��_��Q�0�I�} qO*|��D�?Ld�Ғ�Ì�f���8NV�`d��*�4s���Y�����%,RL8��@j���'�L!Ѡ�*�����<D,qO�d�R �}SdI�&l>=he�6/ �p���6F��h���S�Wu�`�� Yf<8��Q�"�l�����ݼc�G?�A�z�Y��Y�e����C�4�9dʇU�MJ��/O����LP-o200���B��_�|��a�=�@��{�NYx�����C��0O^(�h��� �3]�8� ��U�M7��:��
�8��a������0��˞������rH�e�a��S���!�iT�8�v�H�k3<p6ʑ? ��G��n����wzL�m_�R�\��fb.XƖɱ	�XĒũ�灅--&��ǨS�U�Ɛ�CʰW�\Y!�Ӊy�*
��9?7�Kաɔ%4���� Q�ʄ�cJ0V�Da�'"^���"��4d���>~���{��$^���E{��O��W�=hl�1���9e \[P@�h\���1d>�cfA�D�@�ƴs��9&ႁ:b|G|�"�`�n��c+��fV�� ͖�!)�iN�:��TQ!T��vJ�]a�j��+͖cB��pm�##.�EXV*R�z�TlYlM2)�4�8��)�6�7�ŗ4��}�ô'b�0ȡe��4�� j�# `+��K�_�m��mS���Tab5$j�����(ɋ�*�7�yg�ۋs�Y�$̎�Zd���OQ�0>�kL|��(`d�D�~$t�v��ڥ� �kXrt���h$���A���c�ʍ)�Z����*\�c�a��>ޤȀB�'^��C��ęH9��`�N:���Ey(
(V��5��M3��R��O�������[�WA<Y��.��T/ ��hVL�I_쑣!l�	&�1J���N$����y�'���%�	{8LX��F@��~��Y���WcŦod���M�w�ؐumшx0Xt�&恘	�j4i.H\��e���!WNU�e#��ܰ��C(�4�^�	R�'V!q�C�-]B�lSU��?PMȢ�Б7&���D��P���!U-^ ش\�����J@z ��05��X`R�V<(� �b&i�l��c�'y�tSLV�%s6AT�(dv|Uc�&x�^)3�M� �BVg��uQ�e�ɔ�Ԋp��*a}fa���{�X=0�RGA�hT$H��� �������O^}Ѣ�π!ڰd�g�'H��ˁ�T�+
�8`bM\�O�ꅐ��BELt!*��4I����M:�DD֣v�pm�4@ݎI���zƯ�m�|T�6�ȝ1,T���@�f� �v��'lٞ�Y�B�:i��:�O�o�rt�7'@�dP����(Z^؈�\�haj`yv%�?����	*V��Isf
�` ��+2� ���i�c�K�m>��rIR�|�¤�6��X��c�$�L�5���Y�U~�@�� �$Gw���3�'�����	~n� �*z�~����A�Opt<2�`�d��G��	���A	,A�^�ˇ��Y��CQ���dr��(*�%��Ÿ_b�\'� �I$F(�� �&/�@9�@gȷq9���$Ӻ\�e����!İ�&��\�����9x^Z�Z�A��l?6���M �.*�G}��.:��5���+�c���C!��
�?��q!��ua���đ>���q��*� [��	N�
_�qx��,��A`��@�q1�!�L���BiJ�"�,O�y�ԁZVmʔ�&Z�-����YM��&�+*c���2IH��U�d�Rk���F�/��,Kq>�j�!a�W�ƜQ�Ɣ��ͪ�S��
C�APmy������-9!�}�͝C����h^� ��[̄�gs��9KJ!x��C���`�F\B��E��8�Gȟ��
�f�O���O�n���q��gr�,3�L������r��%��f�+�����^��@��^�?a���w�΋R�z�al\2a��
�ɖ8倠`�놞U���k�^���K�pEZ��E�j��|��#�̏OW��ʂL�nׄ���')�Ԩ�e�./M���M�{^@�!2��ٚ�MjЎՠ�'$%����E>oJPq��m=����ߧ6P�;�D�u~➘PS�@>5>\��/��4�8���	5ߌ� � �8N:,���O�Y5̚�I�5b9�#!\������@�x֜VZ X��0�?=<l���"+�ti��̾�qq�͔�qb|�KE*�>�-K�j���{3��(VHq߄ݲ,�&�Y������0I\HBb�C���!%�I�^��*�D@�%'�p T���SӐh�%O�(sLx�"�G���q�M$X����`�ఒ��­ F����i���@W��)=�&�Pd��/���k��r���� !	�D)��4Y�v���生�� B�ǥ�	+�h����W���K|_v���!K� \�1�Kأ=�V �GH̓<�\<�E"P����F�$_�
�dԷr�^r���+;m�A�U ^�gEXA[�� U����s�Z&]��P����Ԥ9�
Q�C�D'8��`CWwo�M��<,D`���$�>*TD�C��3�`�YǦ��<�U�7J�<�%��&Œ��:�0�c��J2L��`S�
{Ҹ���?R��!aD��>�Ҡ:�:�K�h�ݒux����%I:�j�F��%�8qRIձ?���`�l�*�	�A�!�V-#`��~B�Գ:K�uO81�W��]�0XT����\gD� z?L�`E��F��ّ0��tL0%�'cX�<p$�i�L��֎[[�M`�"��Fd^!�,��o�����A$LDT�D��?	�VȲ�M�A���*��QEb�'�/l�ąQ�se�0� ~��͐rfA�EV��GQ�Fh�=��Hʆ!:hA�@M J쑭�`����FP�X� xS��za��Y�j�c5��I6�x,�7fg����F	U�LȒMV8x�
��$�ܙK���;�]�)�v��7-����'��A+��qb&��t�`�U/_�4=��y��uL���EN�;��YS��v��@�˨[������u���&&�-�rʖy���D'e�09pF��0`|`��U$["��I/`�����ȶEY�����R$���B���-���'8#�$�e�d�p���!@�x���#Xa�q��3��	*4�W��H�V�	'��)��E�?OR1q���xڴ��;p��(#���yӱ����q��
�"S��Ph Ӎ�9rȓ-a/0��q�A:�Ȁ�L!�6�3�(�S��J�}�p�I��DБ��{?A�o�h��h�&�"��'����-L�,�3�*wZ����$k-N��q���2�D<a�%<lO�=I�	$f �;5�*|<QSd�`Xe��;Q���jH>��;P���b����EW�O� 8�0���mK�8���4F��ڼ9�#`��fF�V��`	[4��r҉L�;��8��&o*���ø7/⠒j�0��і'�ڴ��*�(|2��OQ>��p�^dW(,��ĨC��}Q�B2D�+�M� 	,h҆�l|Yp�1�ɀ6�(���'�!��8l	�qҠd��^���
�'�����O p���0�^U����'(*���E��K�-��LA8O����'�xt�c�׏ (���Ǒl�z �
�'Ja1��8>k.]ؖ���ۢ�X
�'ivQxc-��̛`FV�n0�	�'��Jr��i¨˹LZ�L7�yR�^a���;���|Ұ�Y��yRh��^�r�6+
\7t�!�-в�y�I��B�b�@�Q/�)�@EF��y�*��+�)��M0E]��)�e���y2�
�O�T��u��0���l¶�y���6k`���0:����y"ͅ�L���d�P�-�j�����ȓ��m���Ʌ肤i�D°:_���:���!'T�&4h)�N*)z�8��s�� �ǜ��#���WH�����){����}B�����'p��`�ȓq�X��C��<��C�ov���s�����F�71#��s�Iğ�4���o�N� �e+p��#���{����=\�	���ԜL�]�Ð~K@�ȓ#{6�ʑ�M�:>@�C�g�����0H�<��	� (h����덄zN�u�ȓk�H�a'd�<f��N�!�>���	P�a۵��8��m�Hw�NY�׍�������`��ĵ �O��@��#���'P�����Ab8F���[�`{ �P��ʦ��h�C�x#�O����6��o�8�P1��;x�n��LI�����T�+�r��<�a�4�sը�z�GD1bC��A�X�xt9G�
+7�'�a����`����3�I�Y�V���_� ���v�>1�4�O�O�j�	w%�7|�4Y���c����J<�0�?�S�'j�j���K�J�R�wl*{�'c�PFy��iHj�*H���l&L�3CK�k.�VE��ȟ,ȡp�O)I�2��.�L��x���
�����3}��!� �I�`��˒[����}�p��%�D0���<�(��9Za��.Њ
�Z���٪�Ƅ�|� ���k�X�P��-:lqO��V�[f�+���vE�=+I��un�=`Ĺ� ���oV��S�O4�� �(�P8����M��0EQS�I�B�0Y	���d���s��i%��ٷ��(�>�`�#Iy�eX��p��m��,t ��/��O�'%ɢ5,MxP�m ���Y�}" �`~a���+� [��R�5����&��S�1��6OR�Z�.2�g�? �	��FS7w>BT�T�u�*��O���'m�O�Su�8]��ie�
3�$��(�/�����OV��M<E�D�D��xV.٢/W�TH��B7�y��A�$nha�4�S1M����b��$w���D7^2:O�<�4�zc�b>M�"#A�u�|1���!/��"R�5?id+d��p�y��)�:0���a���6r#ʹs�mT�7���Mޟh+'��S.O2�I�h1#0�L�ƙ�B$V�����˓�y
çzĬ���C��F�C1B2DC��W�O?� ��$��?]�d͟��)�?�DǮi����� �x��1{��0�!�D�3e>z�YЯѧx���I�/M�!�$�!p��!,������!�ɮ��0����I�n!�(�i!򄎫A
��9'�T������$!��إpM��"�/ ��B�"|!�F3>\^�i���#F�0yTC\,�!�$س"<�+�Kܕ̦xR�L	�0�!�$��r9R,x��ܪ&� �b�m�8q�!��zfr�b�G�<A��x0lV�!�dZJ,���.���%ք/!�dW�eQ��+��e ������Z�!��FF�vC�;[��Ac�3mx!�D������2�"S�ӵ�D�-�!�D�-��Ԓ-@2j����K�mQ!�d̏+�Δ���D�o�Fia�n�-OO!�ޮp�ȉ�̉=��d� MK�Q!�$ �	S���f!!�F�Wf�Qz!�D	�k5�S�Ԃi~@i�U�ͫq!�$H7!a�<�AŞ�L�Q�nU<xc!��9�\*@���qP���A�!�ĉ%,��d$M�	���6<�!�O�H6��A�/J�L6C�σ=~h!�d��O�bL��!�n�K�v��t��'w�5�AL�zxt�'gB���	�'��r�ƦQ3V�Ń;k��)��'�q�pJ�}/y�3d��l�$��'($����	�i|>)���ٶMd�U��'�lP���b$�(n�BF���'�1� �+TѸ�� h��|���'��H�s�C�df*�@��^��t��
�'C��� �H�EJrG'U� n�)�
�'N|RF(��~���F���'�ֱ�'��,�Q
)}H�V�Uht���
�'Rt���K�H�H�Ћ[~�Q��'
����Y,J���ӌ� N2����'�`�'�#x��9:�+% b��	�'�LI#uLR'e��L��)�%���	�'�"����8�V�&S$���:�'��KW7W,`,���u�]"�'�ȴ��GIBjVG��PV�Y��'�0D����$ JH���GܜIB�'��m�#bZ	s̺A�t��(�f�+�'�v�0��>[P�9��#:��)�'��U{Q�X�~0��;��ݰHn\P��'H�(�`�@�Q]\��lV(@ZR���'���s�H�8��92�O�8*ϒl��'��(��î\�P8#@d҆�"����U�MO�k�L�G�Y70����?D�h; Šw�a�6�(L,T$>D���TʛV�j9�T�՛=�,�Vd=D�h���H�$� )֕-,����d/D���'��I6F�;T!�e&-p�n/D����E�,�a@�(_�TP$��% D�����ߦe����e�;ܕ��?D�� �2N��0���FO�����>D�� ��c7C2=^2����g���
�"O�UyrC�qx8!��F^��e��"O49"�$����OW�x��"O��2#��!`��ဘ�Hy��9�"Om��̘&d?L����w$���"O��Sc�
9��@ӧ���S�"O0�b$��J��a�V���5p� ��"O����?Ttss��&8謀6"O��r4� �d�$Ч���M�I��"OJD�գyL~4�v'��.:" @�"O����,[V"���ĎD^�S"O�P[7�S�cR �g�<x��T"O2����׸x��Z3U$���"O*��# 5P`( ㍐3�=��"Ob�H7J_�WDx���@k�H�<Ap�ܢ\��YA2`
kP�xI�&D�<��A�_��O�L��$N_y�<avAC�cEĐ���W>7��4 �ŏq�<�s�Y4�6A��eV�]�EqB��n�<�F@CS�̡�ViՁf�bYYuiKr�<��*ǣ,ь��̏�3vx���o�<�����wo���4kM��}b���l�<�ŉS)~!Pʶ��\��8�Ch�s�<��aѥo����D��:�,=�w��x�<eeW�Q�t���Ju�"M O�h�<�Eb~VՑ�� PF x@"KY�<��bHm�~���һ�HtH� �N�<	 @L�Bf�X"���
T\�æ�C�<ƤH
h��H��l̄N)p��!D��PG@4r6�\�U��F�~��@!D�tQR +c�����^�D4c � D���u/��$�S�	�r$�:�4D����È,�JD2cʅ'�I��-D��#�K�8^R��k�IǇ���2�G(D�����@u�*$�Qr�%�e$D�d �f� ^�10�aQ,g~n�	Y�!�ۘD�T��#K�OF��g�M!!��ā
�|�����|O������3!�d�c�1�����iH��XU �RF!�DJ����0�C[��9��.��^A!�!>�.Es�eƱ![��@�mJ�q�!��� DH���˔AO�r���!�ݱD�V��'DQ��Y�Lĵ�!��]*NI��5/�̢��5=�!�ē5hZP�4O���faވ�!�dϋ)Ը�77�I"�#P!��=z����BL�3V��R��!�D �X���J��!5~�b2�)Ai!�d�y~�e�A
N��q���ʿV�!�$X�_>�8��F�����T.�!�D	"j��Po@�B����f��!�ąaK>1&� g^�:D�#�!�č7-��]{0��R\�5h����!�dC��&�y�����%�)���!�D�;SD!����c��8���B{�!��;r�����&��k����A>N!����K�7vP3Waֽ:E!��,U���s���0r�&^�O2!��-\�|z���0{�r��Ug�� *!��5z�P��A2~�R<�0@)P!��@�CE���EN�	I�(�j1m�B!�d�J���3i��\�Y1,M�G!�d�t�v(p篎�uݸ�r��&,�!�A�7A��f� ���ȗG !��  ��fo�^UH���\j'"Oк�c��Sܤ�s)A��4܀�"O"\�BBד^�bQZ�h	�\ך�i�"O\��dMD8����H3o�xQ!"O�)�hHu,�"�Ƚf�$%2S"O����H�v��bÅ"g�x�r�"O�< e��c@�P�Ď�t����d"O��b'�&Q
�ԃ�oӘ6�0p"O�<Z�iY]��ه���h'�L��"Oxd�B%ϩ@���B�'%��c�"O<S7�<�"=C��E�r�,4q"O �����"_���*pb-1��y�"O8Z'IS{6�!��x�J�s�"Oހ �!�h��xs�/ǬǾ���"O�Ti4��X���4P�x%�7"O0��U$B
X�� &Ώ}0P��b"OzDU� �cxP���u"�(�"O�1 $S� �M���S�`Az"O��W�ܻh��ҋ׵H�H�"O��q�C;�~-����$t�Z(�"O�L�r�ˌ\?Ld�C釈����v"O�l{FV$k ���͉�T��	��"O�4��AD�0쨡�4������B"OZ� E�8H�@�Ѫ�W�HEa7"Oh��# �/�V���jCU�}aq"O�D�5c^[r
|�Jˊv��@�"OxI�w�P2{�б@���cV9��"O�4C�L�m>h�X㧟%&W���d"O�����C�eTXx�G�(��y�p"O�����X�?��)�t��1O�J���x����*���P�1I����ȓeDf]SB-^e�d���q'^H�ȓX�Ґ�VF�%y�z���E�'v���HJ���e�G��,�D�_�~B���^\cf��x`�A��%Cr��ȓV7tH1��YL�ZY��%@��-�ȓ"��!�D�T�4j��J&MR =�B�ȓ:��q�e�u`mJ�/��o��5�:�+e���*����D}+tm����3���]�>} 3�N��4��>b~��e�ٱ)�P�����M�`D�ȓx�f���lsP��cž@�0���|�@��V�ߊZi�j���D�xĆ�w(��5Lׇ;���k�f٩38^ �ȓKJH��`��ʦ䚗m��-2��ȓ
�+��
�. I�!��z�"O湛T��/0��-z��,7���"O��h�.��e��][�hM>�Qse"O4��!H��n3Z4��f�� ��Չt"O�2���kf���dR;M�d�У"O�}�KM�!�D��۫`����"O���PIW*J��I�hȳ9l����"O ��f�	�����/e�a+�"OVyK���9�ܵ�B�Km�~�H"O6��/
�,\L���E0'�`5�6"OMS�DV)�ʸ[goF�*�xhr�"O6��XB4L��H�tᐌ�(N#�yB�2zR="�肄#��uz�L�9�y�L��E2VKޥ0�� {���2�yh�WĪL����2,*�sBK �y�h��h���B�</`&<���!�ykW�.U��L& �F��5F�%�yr�6���B
�h�<�r)��y!�C� ��(X��C�ɵ�y
� ��Wk_!�
ҊR�:�� #"O*0˶�ơ,=ZIJ3J�A. �"O�@
�Ǹ*6��a$dZ.U��;�"O�)��9!���2hT�8dPV"O�|���F��Jh𑧀#2�0��"OV�i�i�(W�%�D�ׇB�@Q"OƵC���"$��|� �?���7"OQ�Q�Ӛ)��Uz���7���J�"On����ӊ,��a3A�	 }�,P�"O���d�T�IgH=�sD�(׼���"O�!����`s"��#�X(Y	�"O�r�.F:d�
L1�\2SW����"O^L�wL�t�x0�T}R�Q"OR�   ��   )  �  ?  �  �*  �6  �A  �I  ]U  sa  �g  n  bt  �z  �  *�  m�  ��  ��  7�  z�  ��   �  C�  ��  ��  V�  �  ��  ��  ��  3�  �
 � �$ m, �2 �8 i<  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��Y�1/l	aCڷUClM��%ɘ��n8UZ�&]�KR�P��,%T��<A����!Ez��F��\���i�L�/Bl!�S�t�3�a[��~��	9"O��"��IvH�	��EL6j�"�"O�aY���VAv,84jٟ.��"Or�{��+Q���A	L}>q�e����D,��ʆJ��t(T��43 �B%�!��/@��*e��-�tF�Q���hO񟶙��$ڸj7�7�B�Z�X�,D�|�7�g�Z���\� �~���|\�S����M�o�|P�L�"��uȨ�Z�'�L �r�ϓR�<H��Q/_��e���$*<O249��G�/{@ыR�%2��Se�'F�,���s��P5�!�s��5E~���b��ex���*x��ᐦO��HO�����`h%���a���
T�V"O��X"�@57�R�6#�^vʸ��"O0d�7@ 4i�8![���Z[�݊�"OaZ��R�,�"�;��T�xD�9X�"O�#�EMd@R�+F
]�� *��'Z�̈́	�dlqi۹&�ͻ���z���$=�����"	t1�.r��'�a}�c'
�ǓE�T�8c��Ұ<)W�>�O�����mF���& q��I!���F{���(aDQ�p�"Ǵ���-�2�1O��̓�4@�2�3�  ��B�G�ecʜ�R�.���"Od���/Ƽ2�K�Ȗ6nƲ��3�O�=E�TV*�\�b�Z,�T�k �N��y�J�v 
8��&�b��,��y2�
/B�R�x�k��1����jD���>��O~l��M�Vk��8ċ�4$��1�"O����B�)G�"8ȡ*�8U(Aӵ"O�l�E+Y�U>�48�Jӡ/�����"O�-r@�C�\ ����$z�t�R1"O�����'6��]?Y��R"O��³C�&���	¨|����"O^�{��G�
�d{�"hh *O�M�5g¤%�-ۃʗ1)}2�H�'��Xp-�� �\t��m�kJ���'ڴ���"F�<�b��$����'Hٲt�S#����!�
k�ܒ�8.*�6ڰJ獀�6vP9I4e�'@���m�|yZC�%x]��N�����Dz��~���IX�Չ��^k0NXǎUd�<���F'W1�%I O��՛"�Ҧ?�"=E��D��I���5yb �`%U;S�؝��B�z;�Hņc�6�����d�,T�'_a~���T_���+��X�<�j��L��?a����8������(c��BS�9+q�|��]fI�����ht4tZ$
v�X0�'�a~���[K� �	��C����᠂��y�A �f�\�iS�n�*����y��K"��0ՙj2�䫓bR��hO%��)��8�4={�I	
kƞ�v`[:*�!��·|&�!B��� "�� �ռ7�!�J�`�����<�R����t�!�A�_�t,��-�'!��;���|�!�dӗg"%pEhތ�2���jȓ�!�ɲDEz���$��o�ӉĔ=r��x�㉳	xR���7`�bAj�O��
��dh����i˹2s
��)���&#D�`X0�Db�����ᗘm-z�j��?D���"*��Ae̍�C׺r�0�鱤(D�\E�Ґ +��)i����㤟�D{���H%��1� @Yh&�A� =!�$^�yUVxi�V9eǒ�Sr/ފ6�Ѱ>�a!�[}���U����k��A����'g���r�Np��d�{�l�X�'���:�/��{()q�R�v����v��E{�'99�\B���T�]h� ��z}
���9�TPh��/f��PL.s?6ɒ��9$�t[D��
K�,���(�X�Т�#LO\�@�"J�O	<�PSe$*^���a5D���Q$_%&|غ�)�5.�;�G4D�d�Ǝ�D�Ea��k�d�)�O1D���$ޠ�����H<P8�H�ƭ<�$�:�S�O8*���~'L6��*��i�"O�$�LUaa�q�ƦN8eLy��$^�<Y�~�R�� �-I��{Ώ�"`���	J�	l�@b�j%N�

��n@�8#�'k��4	ҏu8Ԥ�TCֶ6�L��˓�(O��#�1d�����BS`!1"O��@���.�HU�1GR�eEޙ��>��)>�S�'~|mc��ǃ>@>m1��@�]Td�ȓs�\��Eő�2��Ɇ���̇ȓDz�8`�Z�(�8=���B7�0�ȓw�.��!�U$��Z4E�}DD܄�`�0��2Þ0�쉁ōT�(�ȓ' @����	$Vd�T��	�v���S�? B!(d�ʑ�xǁ��W<�D�xb(/���%��1��[&H�8a�"N>4�F���i?�p�ҒR7�m`�
VUԵ�EK�<���+���p.C[qK+���D_�Q��7�eq���H�)�ȓR@Q0���*���� 6D���ȓN��U�@�ƈu[Q1��ο"�:%��@��Ϟ�D�fq�(�or�ȓL 0�	AS�8�DI�F~��ȓ;����g�ӱM��0�i��;�m��}�|��GMQ5
�-X���&T�(��n�Z��@U�]d=���д��\�ȓ_��e���΅S��!��.'n�@��	c}���.A	��0�!P���z@
��M����s���C��5!�m���	 h	�"OjiBCN��l��B�]�!�f�)�R�̅�	,��"�j
�>Q�P�����~V2B�IKO�
�F^�%v��%ƅ�>SDB�ɞ|��D�g���d`�h��+B�I6
P�S5�(��!h���\��B��ӟ��'L��$(J���-܅+/��P /*ʓǰ<�� �Tx@�1c�D�+ƭk�'g�I�h��h��Ͷ	F�B���(�MD"O�}��%�, ���U����{I�<I����b׌ѓ�"ڰatz��[��C�	5�]I ��D��=� ��;�V�=yÓR����G��<��M�`,(�����?7E	2(�V�ì{��=��Y�<�A�We��}�֪��5��=(�ZT�<aWob��r�LN�3����FS�<yfɝ7�*�:��Ͷt �h$Rt�<���؜9�Q��	�5��9b)�o�<1A+U�����F��!шP��j�n�<�U!�2���boӱuH�]a׭	g�<��n�9���I��-����/_�<		�7.�����f5�dx# Yv�<�w�
�������*� 8G�o�<I�i	#�Y�^�,R(YQ�"�E�<�t��!Dk��X%����t����y�<Y3&H|�6p��i�D�0@��r�<QT	�Z��r��+�0%!!Ak�<��&G�k����� ��'�	h�<i��$`�zH��b"x6�Qc�k�<�a�]T�t�tMU4R0�a��Ap�<��E�&F�����
8`���u�<i�I҅D�����e�!21,�Q5��n�<�GN<����F��_��#��a�<a�c�(��q)��\1JM�Qx��^^�<�E�|����挭.�&�P�Ht�<9�%9\����$G���q�p�<�r��1��u����R5�ea�<Q�щh���Z%K��2��MD-TZ�<)F��~��Tc�#�m	�}��V�<�W
�w^콂 ���d́'EIN�<i��ع"zB��@�cs�:��H�<�WMӟk`"-�S��j��
�Z�<�V��(gDT��@�=u�B}��b�W�<��΢<˜�����`2Q��}�<13埦ZN`��N/D޸�p�O{�<闇_�F��,�o�vG��R��B�<��2u��8#�E�_K���"E�D�<�Wʄ���-I�ਂ�&G�(B��1"&~H'\�W9��!���QBC�!Kz�$��,L��,!'d˰ �C�)� �����E\�k!��$SH�"OtM��imƴ"@N7 OV��v"O�٪��`�;r�[93�@�"Oܔ
5#ԙg���W%O/\��@"O� �tl@�~r XפM>$�$���'�2�'r��'2��'KB�'6�'�@�A�E(uYT�+���(22 �!�'�B�'���'pB�'�'8"�'�H�"�Ȃ�V ղp	�A�\�r��'���'���'��'	r���isB�	ߌ5j���F����o����O���OJ��O�$�O��$�O^����Oq	aP㚂��!CcA��$���O����O��D�O���O��$�O�d�s-J(�w ߲���+	"��D�O��$�O>���O$�D�O���O�dJi�\q2P��)������{�V���O����O����OD��O��D�OB���<~�ܻ��� iԙ� �7���O,���Ol�$�O���O����O��m�Z�[K\"� � ��8dZ����Or�$�O���O��D�O����O��_�Q��8l��5�i���@�����O����O���O����O����O��d_��8���M8�����'ɘ�d�O��d�OD�d�OL�D�O����O�����܉��U</b��k�;8����Ob��O����O��D�O��D�O���0+��e8��
 ��s'�A�����MK���?Q��?���?�׿i���'Z����Cʗp�~S���;�K����������$[��qA�	1 0
�Ěs?='D0Y�-)?�E�i��O�9O�D߇o�V��� �a��8Rt# -t���O^)ا
o�����Td���O�"�cӬؘ~τ55��7*�mc�y"�'+�	s�O�6L3��4'g���'��+xI��N`� �#��>��1�MϻI���u��<O�ܸ�Jt� ����?Y�'��)擽0y��o��<iΈ�R��U�p&įN����A��<I�'f@��hO��O�i�FU3�
�a��ȱ+$��#�;OV���XԛV�۞ט'��=�R��;QɁ���<0����	f}R�'�;O4�9�$��D�25pyp�	�	��d�' �h�>00]����H���X�4�'H�� R)��T745a�Kڒw�x�T�ؔ'���9O�Yʓg��9���[�DU a�:�Ӗ<O0-o1%������4�L�:ńL�v�^��d�;���#=OH���O��dÀk�b7�1?Q�O���eF޴�D��:	%�Ā$C�2ah���CC�r�l곤C�}&�|�F��T$4K�+ĭ$R�9�A�8u@�8+�@D8t2��镤��*#������d3(����D�d=�x���%u�����-@Z$��� �a:�
"ݓy	ZI��i��hf+��S����U�b��{DТ;����V)&sŹ�OK�y\,}��ݥ9�E�sDV����14�f�����jj4�� ��}���H�OVriK�O>bb
ȸ�,���$���^2�TCg%��Q���YqJ�[n��d��
�h����O�s��@22�	OgTu1ì�'2<�Rg@�|���'g�'��`8?)�+��x��uyw�F�g4��2!V٦a�	��ԅ�����	ßH���?����]�D�G�zT��ڒ�b����u�i����jӊ���Ox�D��fQ%���,
1e�����F���	��� 1�4%Q�4v�(�z*O�d�O���d�O�H���U")�J�����.Ly�I��ܦ)�	�X���(!�՚K<ͧ�?���E��}s��U�n�E:��N�����V�p�I�@"�?�I� ���<i�
����K��5�$�r���MK��uz����x�O�ғ|Zwi����� b�&���A΁M ��O�A���O,���O�R)�i ɝ-}^���M�_�P�ڀ쐚r1�'���'��U����֟H�Sk��7�.�h�6���'J�\66c�p���(��ay�"��YDt�S* �����H��p�G��>n��?	��?�)O
��O���'P?�Ȏ$:jSFإ)VX��u�>���?a���d��e+'>�C阌;Q���ȇVֆ�i$���M���?�(O�D�ON=��I�"';DI�0��;@ubw����f�',�Q�h�$G�)�ħ�?��� A�kn��Y�+]U<*��q
ئm�'�B�'x[��Iꟛd�l]��G�(�b""� �M)O�D�P��Ӧ��������*1�'��ՠ�+�/:�&I�m� ��4�?Y�j\��(O�S�?Oҭ�4E�0(�jj��Z9β��P�i�hf�w��$�O(������&��ӭ)�ƌI�lԀq�B�$�ǡ�<���40��=(O�$�O����On$���q`)Q��$="�0Xq \���I�h�	�# PN<ͧ�?Q��~����K�7I�	C4")\�zl(2\�L���|���.�����ğl�����R*�� �G?4`���4�?AsB%�����'
�_�H�#��6h�ف/�]�r@�Mk��r۠�<!���?Q�����~x��a�PA��c�ٌen��!\W���������'�r�'*\ !���4*���\0�r��Ø'q��'�����K��Y`Z��~>�P%-���l�{ҫ@��	� ��I���?Y��#}>��l�2��܁�`��,ˎ���f�+K���?�������OB���E�|�'a�M1��F�FƊu@U� �ډC�4�?ɋ2�'p:a3%�ējI¹y'��+E�r�	G�lZ����'��($���ڟ,�I�?�s3��V�V���*�A�K²��'�� ]/s�X��y��� @ePլLU�5�F瓈媜h"V�����x�F���՟��I�H�[yZw(�p���}!�yX���i3V��O��Q� 5��`F�����n� ɘDh�W.^f�O%Uۛ��,� ��?Q��?�����4�V�d�y�F$3���'-,��7i�0[s�o��� �Sj:�)�'�?ɐ�	2R�m �@�9���ŇT7����'B�'�&E��W��ܟ���[?9£%�f�[dF�K�feV
WL1O�}���k�S��0�IV?�p��#�
u�c��H�ĉU�@�]�If�\�'��',r��K>dӸ�/��V�)�!��*��ɥF۲�K�.?9���?q/O��� 9_69R�/�'B�\���!�&p��8�E�<9���?Q���'�E 8c*��ZC�\�e949�U@H5O�<�qT���d�O����<���.�@}�O����cד��,�ՠ)�I��4�?a��?����'�>�֦��M�%�S�A�����Σ~��Ԯ�}}�'R�\�|�ɽQJԕO�©	v�)ygl�?!��i���n7��O��|�I�h�x#�H"��%��%��)z�!ZT,F�6��F�'��⟨�S��G���'�"�O©���N�uƌ�+�AF8f��I0�&2�I�����#��E(b��'	�0l0��˓�1��f�.l��'_���62�'���?��:���P�LiNQ+���Z�b�>���X��Hm�S�'HVP}�c�$G"�A��)s��m�G���� �'��D]�����r)%E���¢C�!��lS��M�p "��5�<E���'�ݲ`��Y��@J�H�GN��bb�l���O�䑝zx��|z��?a�'���{�#O�_�d�� *֡��R%d7,U�O�'i��ُ;��bf�� 1.��� ƔJQ�6�'N-4W�p��ݟ���Xܓ'���5j*�J1)�+&��Q&�h��E(?��?Q+O��ė�:�)�j� ~r��J�D�D���<���?����'���S�c6�Z��t,�V�L�*j������d�O*���<�:�$���O�ͨtN�l=��	�
�}\����4�?���?����'���h���M[��b&dc�*ݚT�,�S�Qi}r�'�T�p��.�\��O�BaGA�<��QG΁=Ԙ�;�i�)S� 7��O��0��gl����;�$�/^J���r��;o�6�m����f�'d��П(�B�Wo�t]��+%�Be����G�zi˓�H�^E�d`�}��'�85e�1՘��)�.C,RQIaĔ`\�i��
���	ʟi���՟���㟬���?��u7b���y`�K�(Z��B�IC(����ON��s�ʭ1�1O��XUr�F�*s�m�R`#E�U���СU�2�'e��' ��\��ʟ�Y#
�I>�D�"`Ԙ������M��Hh}��<E���' &��G��2w@-)��6y�v��OzӜ���O8�D�z����|����?��'�8@[�BZ�ge�QYB@�	7��I�e<��5,=�1�M|����?��'꾹�1n\�	R��Q��I��HS�O"�;���<Q���?�����'Srȣ��ޯk�<l�@i�i��x�O��:V�D�5l�	�����Yy��'��(�!��]��Q� �BE��)���#��������?Y��K�ˊ�������A�DDh#��`@4�W& ?���?Y.O��$�����5a�*�I֢Q�%�X����=�*6-�O\�$�O\� �I�9�TP��g��)k����ّ&J��r�0e��P���	埌�'���ɥ;���$J7�I<F( �L�sH��!�U��M����'1��ЗL+0�jM<YU`N8y�j'ǚ'�HQ�S�����NyR�'Jx# W>}�����Әp�L�9�Ŕ'hn���b�~��}��'�$�S�������	��!��zۮA���T-��	��Q *�ҟp��Ɵ���?m��u�L�4.���fIԴeXD�z������O�I�V��;�1O��F�[��.PRF��6+B��0鰴i^�ӕ�'���'B�O��i>q�I)x����"�|ik���~	05��4/�)9�+NP�S�O�r��W=p;���7߆���;V6��Oj��Ob��p�<�'�?����~�bR��]��l�$|�ܠ��F.o��b�Р�)����'�?���~R��5c0\	��H�} I
G����M��=o:-O����O6�6�I�cr��K�
�Y4�2o�N���#�p�0U�In~��'t�^�����UW�ZRJ+6I=˷��(��c&��eyb�'���'��O���s3l(���mv�����Z<K�豪E&Y�1N�	����Ify�'@�cVߟ�1ݹ�E����h9�����M{��?Y���'��$�t���ܴ��m� �8�Q�l�o���'���'��I����T@�`���'�6�����)Y���SG�U�A!�~�p��:�IΟD�d�آOĪO��oB.o2�zE�ï8A��鲾i��V����6�~i�O�R�'��,8~{]+ed��&�r,��H$"��b�|��$�8��B+�~j��L42�s��H��`�"��G}����9PJ��'��'���U��ݖS�5R��Dh ��%�t�<��?�ħ֠#�]�<�~*�홨}	Bd۲&�>2`���˦�j��ğ4�	ğ��I�?�����'�D�R��U3x�<9yB�ݖzC��{Fdӎ0�$�@�X�1O>1��+׀ �8��%x� l!��M�$X�=�&�iz��'b�(Y'g��i>��	��h�H},I�b�q+�@3� �9nq<a��F0扬(�@�0H|R���?���K�dd8��2&.�u�	\Nh�z�iF��,N:�����ORʓ�?�1]A%���x�ā�Qcֵ=/�5�'&uZ�'���'2��'�[��0�L�N��3���R'�$"�k��Ȅ�O�ʓ�?�-O���O��D,)���x!�\h�Ԃt� x :��<O��D�O��y���O&��<Q����:$�iO�G�"�2U�L�Yh�'M�Ni�FX����GyR�'���'�l���'�Y
U'����,�f�l���A3�`����&Z$d��O$˓(�֕ppY?i���` ����Ņ�Ш���۝dTn�8ݴ�?�)O����O �D�z��|nZq�aQ'�������	�>Hy
6M�O��d�<!�̅L����|��?��F莚Z�PH�m���U��L�TyR�'B�'L���'�s�@��8�q#Ji$ y��k"�oZgy�l ,��6M�O*�$j��I]}Zw7�=k]T�c�MҊ=.��'���9��ꟸ��A`�X����,�R"2����А�iF"�X �*I�7m�5ӂ�mZ������<�S���$�<Ѷ�K�XH�ɖ8Z���(���6D�1�y��'���N���?Y���!x��x�&-J�0rt%K V
�&�'��5O  D%�>y/O��䨟T�T��8y7�t��D�IT��"�'���7Gf��?i��?!G��	^�+��;Q\|R(ں\�61OHp���>�-O��$�<���+wo�$v*���F�	�`A[%�Uj}���yb[�H��ȟ��my�(F���bmU�E��uB
�F31n�>�-O���<���?Y��N)��3��?y�ޝP�	�-'��r��<����?	���?y���d˱n�tΧqW*�Wɖ?X(�W�۰���m�gy��'����$�	ӟ�j���~�iH9JZ>�y�M$���2`�U[}b�''b�'���p����N�DH�w���`�sմ�v�ݱ"3��n�����'�2�'��J��y�^>7M�DXaRU$U=.\�9�g돮r��&�'��U��RW� �����O���0	 ���!�Z�C��8E
5ʥ\}��'FB�'��Қ'$��9Fj���-��lHVM��g{��@
Q���m�[y�Bտ�V6m�O��d~��)J}Zw�PU!��j�� 䇹�X���4�?��K�
E�}��s���}�$�G�>����˩<��M����h`:�M���?�����pX��'�q�1�j�襹��*9%��Z$�s�й�8OH���OZ�� ���?-�m�8A�9�$���k�&�����M���?Y�'P��FX�8�']�O�h�IG-!p`㊟���AָiJ�U��y�/l���?���?a�iJ3s�Q:B��3pG�H�Ʉ�t��v>O&�p���>	/OL�d�<����ˎ(�L�����!��@�1)b}�d��yR�'["�'R�'t�	�mgJ��)�?[��Ċ�#�<u|<D���Ĕ��D�<����d�O��$�Oހ d�˪�F�'��	0rJ���:2��d�O��K�^�6��OT�E{t}��>�Ҕ�r,�*�m��ረ�V�"^�<�����$�8�����σ՟L9�lɑ,�n�H4���`-z�������O����O�ʓxw��cF��D$�0��\r"�[Z����4a�6��On�Op���O����j�Oz�'�8��c�D�t�6H��*���sߴ�?	����$A��&>Y�I�?M�E���);4i!1N�a�1�4�ē�?���l�Z��������H'r�Xj�\�t`�PZ>�M�,O�,�#ZǦ�b��$���Rx�'�XLJ͒"(�4�!1�S��,���4�?Y�upd1������O4h(�Y�yYZ���\fp2ݴgی=�i���'���OZ�c�x(!��$ܥFY
l^�Rd׳i��5nڡHT�-�I`��d���?�����T��� �%k�H��a铍R뛦�'�"�'��`��=���O�����|ёM�>�,8��? �x�fӸ�O�pg�M�S۟����`�I�YsvU[��_">P씙��/�M����&������O���?�1@h��,ʂI.���ᯋ{��'P捺��'^�	��	ɟ|�'V2�qD��)��8�B�*H����G�VO^�$�O��O\��O�p��;�6 HG�S�T"�a�����l��<���?q�����6k��qͧHa��SJ�P�}4�@5�:��'���'�'���'�Z����'c��k$Kс>J�;�,R�X����J�>a��?Y����D�4L�@H&>�RT�16�DM
V�J�;�� zR&Y=�M+����?!�/�z�������&��闍9~�{�J�to6�Oz��<�')Lx��O���O݊7�@qE ��B�\*i�2E �$�O��� ���(�T?���%Q`�!Aj��K��h�pӒ˓I��Y*c�i�맪?��Nu�	��ܺr�#?��Yb்*+�67��O���[,���0��0�'/Բ��@�+
d@Y���	�W$�7-	��EnZПl�Iɟ������|��&SǮ��@L�%A����U$O��?��Aʛ�?9���?1��)�O2��FҜ=�|��bH$:���f�����ҟ�I�q�L�N<�'��I,I�ؼ�c�Ű�x1�ǀ7�t7�:�I��&>��	��T��8612�%�(�lx�ħX�� h��4�?����[����t�ɀD�p�m2��y�@D�%�l7M�O.0���Obʓ�?9��?�)OV�� 4XsA�>)� �xb�D:�Ig��5cw�'���I꟰���˄l�,�ۤ���TH��A�3'�6��ly��'���'��'�,���'B���^sU� �^H�����rӊ�$�O0�+��O2��E�&��Ǹi�j��׏c�hX`׎�&z��AZ�O`���O�$�<���\�������D5����I�uvZ�B槉�M����?��������O"Tu� X>2�6��U��9\7�\��4�?���?9�k����?Q���?���&���Z�'iPAb7��LD�D�x��'����\$\�0�y�����!	BD���gܝnF����'��-;��'=��'���Q��X'xn������4 <Es4&� 7��Ox�d���8ك���U�*�`(3t
A`�T�2�J�o��ŅesH7-�O����O��i�i}"U>��kT�"MriqDm �f�n�	��ݻ�M�Ď����'���|b�'�$���N+"O.��V��T��y"i���D�O���F��f���O��'�?�'.������;��d �k�>.˔�&�I�d7�AK|����?q��v�t�z�/�9C��]aR����m���i�b��*+^��'��꧳?qJ>q��_6�<	�'h�ay��n�/F�|z"5��8�I����py�hH���"�?}���jA�V��쉤Ǩ>���?���?	�����o�.�A@�<E��$�V�:hvX�t�|"�'R��'R�'\���֟��3�?f,��&�Ȍ���1"�ir��'�r�|��'�R1����4i���r��>uڦ��#�"V��9�'�.�R逩.����O(Ω{��m�`���:8t���'�����,U+.6D�e�
�1��p�'�Xyh��h^���&��Q�ұ������j�$[�KA�{���f۾�����D�����cd���lY�Jܢ�B�J�1�����ǼR�NEʇ���&����3���W<"|KtiR�|�d�C)F3�HD0׭��R�ʁ2�nǚz�Rd
O��@����m���2%�^E����O���;d� U	"�V�,~�a�h �I ��:�*��r�]h�������$:9 ��'ۘϿ+gb��"�b%\���y�fԡrv����ϧa�PT��oĝ@	F�3\fV\���2Cf�,/�G�M�<3�l�2$ $3�l�rҬ�$5TҘ�C�'q�����x�O����Y+�"�����-/t�"O���D���Y�$�\�֝ۡ�	�HO��@�����,Yͪ	[4��b'�i�I͟��s��NNa�Iʟx�	�[Xw���'G����&I���p��:h��,��b�O�3��g 딍�
����č!-Yl�PrH� �>m���#9t�9�#C� i���?�=Y�)c�@�pƾd^ք�u�K?a5JUɟ���c�'�剣'�tXF@�.��9S�%C�rdB�	#K�Y�#�#l�q��+ )-�^�I���?ŕ'�(��b�:9!�"��o��ᰱ�S�C*q�Ѣ�O����O��6e-8��O��Stf��"�@
"g(u���0��
ܱ/Zj�!?=@|����%y���Ó&-0����
0����É�;]���x4�5��	�P���O6����Y.S�
	��.�	���5E%ړ��O���:,V��RD�V�z����"O\� F��h�v�b�fو��6O2��'��I�ndDPݴ�?a���ن��9��� jVr�:��.Z�ˆ)�O2�$�O���E٣|� ���O8\?ne��|:Р��W��H�D�Bo}����J�'3ni��Ϋk��h�W/Xޠ��V�cl,ꓪS�z+|�ᬓ���5V(�B�'� )���)�֌y�N�D�|2с�%s�Xದ��L�${錳�?q���9O�`9���5R��Sꞯ/�`�p1�'�OT<����C��Ĺe���� D:OМ�4O
ܦ��ǟ��O!� 1��'3��'�Hpd��9�2��S�OU4Y�.�v$`�k��/�T>E�|�	$�V ��UIU�pkq���=�R�P,��,�U�O>E��pr|�Q��=cEF��� u�6�7�Ǚ�?a���?Y�����'wJ�X�m_�B�B�� �y��'��}�*�-,�� 5n�sbT�1�	<�OX�Fz"T>	�'	v�8%���']�T���Ȍß��	L᨝�`@�ʟ��	џ`�ɥ�ug�'5r�V!T�$I{��MC��9sK��~,V�* ��j�"J�m��x��	�4и�R�Ҳ�Dx�aɦ{�~��k�H]�t�O��Ybu�'k�Ua�*F1ug&`� �Z<���'6��3�Z՛�-l��� ��f`��LQ�>��D�2��0 )�"Oni볥ֶ۰�`Ҁ� �fII�'�����M't�~mo�OF\D{6��+�lĈB�G�d��I�������E�ϟ����|��Ό�&5$A�g�L,/Ҽ̂RIV�"Mc0cܔL6�|�q�E���<�%�zZ���r��1"��&@X�)
�[!�X����5V`�Ѧ^d�'�&D+��?	�e��v�5Q��;@��5hՒ�?ɏR�s����
*��:�X�&�����$D�|�e恢D2��m�z(2mh�x��)�O$�)��T�s�iLB�'&�R�8 B�j�#m�f��'�Q�JEd�� �����П��0
 ���<�π "�"8�q㛴|zl�v剫V[����(ڧu�P���=4{
M�"/�LC�<FyB�ˣ�?q��)����[��Ջ2�����Ty!��0(D���vÍjwԝS���ZTa|R#���13=���H]�d� D� S�Q�$*$�±oş��	G�$�W`R�'Fb#ʇ><j��OB9f~d�)�b׳&&&��p%��%��s�XY��"��~���;xU��'Zt�`Q��Ǽ\�t؀waN4h�����b�|Hz&-ɗO;�>�n^�s�,	�$�C+Z~@tMO�x$�(���O�$$?��d��?9�ع3����ߘ�)� ��<y���>i���/�V�H���:+1�`�w�@D�'	�"=�'�?�ER�	@����H'.�� ��C��?���r>�c����?����?��*���ܟ�A�6M6�(�DЫkؚ؉�｟$[C�I�6Ѱ�R��ί�p<q��4�Nu���#��8��Zp?��LN;5�F���BUW��x�E��X�Aj�e�6�*���	]r�]�2�'�����O���l%�(��a����+�����ȓ4U��p�*I���/��j	�YR��d�|�*O��ɂ�զaX���:c�>� �T�?c�%#�Vş���ƟD�I�g+he�	���' FYu�ҝV��ع%��xH=�$R<�~�H4�k?��8�F�Z����lK�?�����`�C�Ig!�U%�A�Äݕ%��b��D`X����&�үd��"�lÈN�*����Ֆ-^L#aJ�Q�?�C�s��U���D��4N���)��f0D�ta��ҹ,5�Ɍ�hp�6jn�`��4�?�+O�r��)�Iԟ�O�|ܰQ�P	]������Œ�d��O0���'��	��y��T>�`#�4_�r, Ҽ@���z�H:�v�D���&�F�Z�K�z~�"7N�0�Q��S��OX��(���O�\(7�O�
� &ߧ\A �TD�O��"~�8�4T�)F��mq5A�-n���I�ēUDZl������k��Շ{�4�r�Y0�i��'��Ӓv�܁���,��#(��Iї�ưu��+f#��(��}P�N鴐Zf�!P��遾��I8��O޼C�˿S㾕���˔|� � �/>�vd:�(W�<�Z�Ȇ�?�Q?��Hb�����U���ck�,׎L)���O��m�X�IS��T�IҟS��%�z,��.R�BM�JL�@��Yx��� L@�����0����*}�Ǫ(���|C�O^ls�"��@�W�Y2y~�u��b74��92톊ܦ6�P���9f`WP�<���2:}8A��R|dq�q�<�%%�,�������B�BIg�<yd��-L�z����(_V����O�<�խ4O<0	TO��x�]I�<a�MH  ��A�˖J��+�� T���d�[נY�TD�?�ȵ�si6D�<24��{Ah���� 'G+NO��y�ƈ{�p1��Z�dfp �Va��y���k;̩���Y�r]�%�B�yR�J:nN���A#]:�xţB��y�NN�w��$�ÒV&ne��i��'�n���͘ %x�\��5C{zq[�',���kz�*5HR�V�<{DhP�'|��K4��Z�k73��R�'�d(����L��!餤�22?%��'�N�����޺���-��3��u��'&� �E�ۡa\�,�JN7+b����'�Ji���
��jx�)�#h*�I�'�Yfm�'3 x��@�=JYVl1�';:�C$�P�h\��X%'O�G��h�'d� (%�ԛD����50���'hN��E*BvT��$�;���'e�A��X�2�6piPÎ�[l�[�'��e���M�x��t+�� 
�I	�']x� 
Ӊ,BJ���?y�h���'S"ՠ�]�D��!�'%�r��'��q�tb7:ώ��q�ֺ԰��']J��W;}�QD(6bD��c�'�BY�uD����0��5+b�5���� .u"g ���P{v�5
=�;3"O�{�M��z�ys�7
,��"O\�$�-;�"=I�m?'d�[�"O��;6���v��s", )�lV"O
T������X������4 ՞>����gX32-�U����<�
p���&R�}:�8R�̱�|� Z����@ 7*�c&�ȇ�ē��1�@���Z ӕh�ȴy��nt�PH�=I6�sƈ\{�S+$��m���O�z�a.K~�tc�!��)%�����P�9����/Z6�bؚV�ɩy�
�G}Ƒ>k`�DefM�"�L�7k�k���^4�V�(��3���ri\� �dbE����5k/�@W����Tj�f4����'V�
�s���
*eFl"�XJ�|aӦ�O�QkB�E0Cq��ABaA<#�(��q�	�f$^1O�<d��16��k�S�4�r�]ґ���Qa�;3�R/r8"���/?yqjV�:,`e����+�2p����nj@�ۻZ;�Q�@���C�`ϓ|���5
�	����,y�1��*gz�B2}�GG$䅹'�ԪW�&u)1N�"�t�rBNF���cJ�r+��N|Z��״
mF	Y�Ş<vb��F/;L h��g��zb���%ǚ.|b�� ���9Fha�#.�*�O����.X��Q3��'�z�.��`@��<�6�R5��G:����%& ��샧e��; ���<A��<|R��;勄!H�4(+�@�:dl �c���O��"G��f´�J�O�6B�6�Dߔ_	�T(��^��
����L�( "i�����$���̓� �P �����ɼ;3`
V(��3#ƚ�W�v}��DH~bJ�Co�����p��Mb��	*�5��c��@;�c��(�dْ�'3&!Y���w1v�&Egݩ��,¬	��p��Ml���;������<~�Pq���Œo��0���աh:��K�-�`���':n����K�J�'��K�d\�0C\!�:ષ�^�{��a�C�5L��t��:�脹����o��x�o��7��C�.��| Hۄ����&zQeSh�X��$�dC/�ug�x�)�!Ej��kb�R��.��GBD}R��A|��#p$]�l/y��',tL��O1 �R,� �A:8
�3�{�(&\�qO4I�'0�X��a���:���n�+�65� ��?��U��li6(Y �����@��Xg��zI������Y�^��I�ܥ�SÏ=Gz2 ��{�ώ}��nǫ;c0�q����j�'����e2��!6ləx+ڜ����N@�X"�'C������9�	�՟��<���w��P'��N����(E�;h�(r���!5�N0���L`R��䂖O+�3��۵*�D8���'�.i��
X �M�R�(3�O�>�S��9+ ��"��]�.e�l	!�CZ؞�	ѭ��m�$ט=0�2���L��
"Ȕ�)��mH ����	�<h��'���H���`�O$ C�����=9�,"7��*��$B�(I��'�FPyv�I&���O�ظX �P1����]�rcv�J���k?�uE��OnZ���Gz���$�F���U��z��1��DQ<:�r��dL��̡�c��H�ġ�O���ɋ.[��j��'3!�0�G�dϐ��-���p?����D���� Tgp X��Qn�ȑ��(��8��*Dzӧ��O���2!�M1��4+�=�$A�8a|��Ij�Ń�h��4`*��\���I!l��{utK �R���� 9w����O�����{����F�#�h� p�U`�Hܑ]�X����I�;�F�!�`�8@��Tb�@̱X��@���\�y�`ȐJ^��8���:\��`�����˪#?�3�Q�*1Q��:���1D�ĊK��p�<1@�Ԫ4�qq�3��g~�(�����Z4a�hR(�P�$B��u����}b�f:m�Ϡ,�0����
/[FhAc��æ.��Ik<l�'�d����?ͻWnI� ���j�buR�-�i/r��/ZQ�t��3:�Hx@��8;�>i�6�U���1��|���'n�rbH�:I��O<Y�H��6�*XX'��1|�.�����u�di�4F�x��s�����?E��@Ip��%'�(!�Q�X	��	�D��Zv
��P��g�')��� ,)�%Q`�lj<(��OR)I6��|Y�yR�-5���$`��б-�tJ�)N�p�[�y9�fD��p?�g,~,P��b
S��0�ɏ�N�f��,OLDJ&��.:�?Kn��������$�����7�޽  ��m���wO�%��.�,����FI�L���A�n�*B���NP���0F-��OT��?Q�Q��J�QI�.�8�q(C� O*��B-��$��P���B�fՃҮ����K�5{M�0~"���O�=*v(�>���O��(*���1x�*a"��'��´�0���Z�J$��a]?b��;�B$P����	�0�;A@pF��fʕZD��&��[ff�Wx��!��2Y:~�#��� ~�`L	�e�<�P-���BX��sִ0ږ׽<��`y��U�v��΅�AvP�:C.\��j/��?I�#\S&� 1��*Vq�HKgD��a��2a*2��1A���n� o�����\!"7J�LTH�is'��;0y��	��&A��J]���D���-.���N�Ge|�J��+`���0��<yP�W�t� � �C�Ax���n�1��T.ш<�$�A��'?��L�U�h�"-uȬ�������/�$x(��7����1l
�k������H?Q��e���� H9��,w��adk�Rβ!����eF��0��]=6�$�Y�H8��7���i�'N� ��0�,|ZQ�M�2-�DH�E4�H�O,}XU�D�S��3�b�q���*�)�X�xu�
3#��X��,.��0$�U��1q4j�5���O��V��q��qYR'�#A*R��՘>ᶬ^�T� S�a��'&j���8�@T4=
,j�Hvf�݉�mE$�굑g��� f�bcNʽZVE�d�N;9�����v�`��W�Y��3�j`���b����ě��<G��`@�ˍ,2uAS��g�b>mJp�޺Zq�$3���W��E���F��lJtÎ}�N-�W�V|�ڨ0�jG1��ɐ���0y�z����}��P�*?*�'UFP슥E]z����K�I�K0,�YW��J�p�H0.L�!��ɸf�Dʟ\���1!��%�%�ׁ$Z��bᖤ5�l0S2�[��`�Q0i]z(�tC�:0��(��%0�V)\���� K� Ic�֓v�%�'��i���gm&I�"�+����h�4d���8Vf�`$B7-95H�$�N*�L��DԮs("�Q��P!1�a~�F�X<X��fa�;�|I �� ���a^,ZQ���*F�4��ŀ|ٓ0-����I`pb4�t흵�ƙ��̆vj��:$O���p�L�X@x s��Hp�$�W�-��tȅ�4ϐA�'7�L�p�R`�<�;[��8T�O8���Ը-����nX�?�<�A�'$�l��� 6C��#��(*M�4! [�"���àI �:�Ύ�]�a�&��.-�ӊo�y�c��v����D�%8`\��f���$��`�����&C2v��u��Q��*0����4Ji�l`֥ݳB���F-qL�u��'UZ@�R�ʔ)���{��L\*�Jѭ&h��M���Y�W�ܴ��Oq��x�+�C�8����Xh�xo��h�VH�,E�!���2�=�r?|��S�֓[�f9�Eر,/ P�q�O��H3�Q�lB�d{��[>H�+G�|"@jp����39��� ����X-.��8;*��@Ex�����
��((�G�΅g&���W,H�K.p��$��;��]zb*;<O(uєA��a�@�h��;jm�3���:�(��3\�8��n2��5$i��yC��7�`扬V�(]�Fo00Ĕ�2NM�B�B�	�f�����"-6ܐ����n:,�x�Ι���!�		H9�0�&�O�s�0�"�c�Ճ4�C�#�bqE���<o!�ԁ0�Ӿ58"lۆ(��H%)'�?-��#ôi���I��h�t�'t��UI O;*��Pg�=+����I'�
� x�ՁM�~�x�`� ��?��"u�N�� �� i�ܡ��i 0�(�� )ܠ��a� ��c�V����E j��9�ZJ~A��@��i�w��T  �quT>c�Pʄ�� "w���E,M�Ԑ r�&1�	2.�%��A��ѓ��H����'�$oƆGD��:�K\8>\1�DJ���U����?F�oܓ�xb>�R.O3=Z�*#��6�B�q�,%`�5ѧ�K�r���c'"�<7HQ��#i�qr� n�0��
�69^O\  �C�b������G�r�̧.U��U���W3 ��S��8p�V�9��HX{1�}�����?i& ��{c������Y�"�9j�����䜱MD2,��	bQ�β3Fr�]5 ���[��^���Ê���'���p'�5;�45k�����>A��^	��qr��L${a†V&�U�p-�#_��S��0姚�+	��fh�N����O��5hݘN�p�
�ڤI���+�7O֌�p '�Ɉ�M�� F�t�l�0a��B���1�+Jz��)���j{)X�G�/JL1O(Z�O��p<������'!G�-_h��0CNQ}� w�b4�r�ǛL��5���=L(�#)W���I�)��B�"�i�Y�TIP��  X�j�S� aS��`;��{��z��!(j!,4K2ˈ�����s�>P2��S�|z���&rS�Ic�]�N���4lB����X2)��6��֯8�s�l���S-�<J���@L�tKS^�|�pU"͡@���<�!�/���� �LOܙ����<V���unKB����ɍ�(�X��gm�<i�Ǻϓxޖ����0 P�?�B,TL�0嫄:%}r� �̦����_&|�R��_�B�����IC>II�Y(!|Q� Z�):K�a��Γ����%�6Y�:@��&!��	ܢ(Y��
�wH9��!��k���f��5_����S8�����5.V|Tx���ß��@��4y+e�=r����@ 2�2��(\�R���d�� w�H�@����ˆ�Q"�y��4�"S�
�5U��lyס�6ؘ'7�m{ө����JW�9OP��%��j�dȁ�ˊD����\�:@��K���	)G8�t�ҥ�.}�bX� RC�䚐-z, 񃬊�G����L�3߮ۦ�2H��r�}��<����	�=ᑆMe�S	�v��ɪ���4
�9J%F�MC��O5Rq�B	Gi���Ǔ6��1k���I�J�cTE�G"��k7��v��I5)����V>����D��v C�A�Rb4�k�H���8c�1�H�� ��b]ve��t�7.�c�ā����x��AW1=c��[5�K<h��T��
/�y'�;D��#V�Щ\�F�m����'jF �e��GB��A���O-�ˉ�>(" �Q�Ƅ_aA��	���LW?T����uk�O���P������D~� H�y��a�8�䚸]���'���;.��w����O�V�9��Hf^��-I)M�X����i������ux�$+��+[Y�x��G�g�nX�0a�
/�6ТoY�d|Ex��5�&��bjq��I�ٟ�y�3�)� ~� �)�#'���E�AT�����mH<1�1��u ��@�T)�Û�y�cS<+��`�#O]a��0�!�(�yB��4)�� �b�:\��kW$֮�y�C��'\�\ԡ�ce~�sQNE��y-�<?���M�EMd�pֈC��y"�6�DA�n�DV�դœ�y�e�;f��i�V�.g7� ���P��y�'X3;/�![cU�fW��B�B�<�agD�^��	$o�IQL	Y�u�<�ԀR�'<$lQ1c�-RR�I�p�<Q�Ii�p���+<@ u�7��`�<�����y��nH����0 ]s�<��F�+�����~�>����<T�P��eK�w1���HG�`o�L�� D��r焮�B\�c�6"ߎ@��;D��C�N�(Hֵ;d��1#�r�F#D��i~m}
����^=\,�e�!D�� �ӺI������$�:L�� D�L*U�1
�J��O�`<z�vN>D��!��G�z8򯃶Ail�{�f0D������7`"T)�h�=�p��p�/D�āFʟq���E�YX�#WO;D����!�"L(X�t����`0��O:D�$ˑa��~v
�Q	[��1Wi7D�@�HٳA��L�A�2&�zq�T�/D���ŀװ���@1@��0��+D���#)I}Q�Pr�D�  ��ɶo*D����˻ }�a�r�]1��)i�*D��"�� g{��$�!޼�1`A;D��JD���k-p���B*}g�4sO9D��ke�G�E�.,�c�M���B�e8D��0!@�-a�����ބG��Pwo6D�X�t��;^P�uc�`����3D������S=&e"'χ�*|]P6�.D�P���8N� $	�=�Ti�Uf"D�H
4�^#mK@\E��2x�B��e"D�J��ۺ$bRp��D*0�E0�"D��0�ϣ���Y��_����?D��dG�'6M�V 0(�%���>D��k��E��liP`d^�/��e�"k7D��2$��,�RȚek��s�j�B��3D��j���FX���gJ�L&^�A�1D��o�<(vV������P�n�C�<yGK,NT�J�G�#�4��� �}�<aE� =��� ��^�����^z�<�n�>�����⍠��*�s�<q�i�ZBV)�A�j!#^y�<ɵ�U!Zx}��U�]�����_�<i%��w<f�s��%s����]�<a�a�O�fՂCV��HE��`�<�w)	_2�5�.�\���Я^�<9���p�(8�e/؈]���!��r�<�g�/Y"t�9����d�7n�v�<t�U�%�z�� �q��@c��s�<�"OE1+$x��Ŕ+�bų�h�<)�G)��8�b�Zx>����c�<QH���=[�S�XJ�e�	�y�<4�	��<Xq��ѵp.�e��s�<	���œ�*3^ v��EV�<Y#쒅[t�e0~hTTC��Bl�<�B�F�G����V*.�����L�_�<�� H�	l(4s���֌���^�<�"��i$m#�C�(f�dA�Y�<� ��$d
;Z@ك�R4
UD��"O��!���Yf]�c,�;G�Y�"Oz�ۢ�����,֓G|�3"O�륬ۄ��e�RK��.�b"O>(����E���� �ә	���a"O��a�b�3ъ`���˽K�V�@"O.}2�ቚa�^�Z�A]nN܁"O�=�	޿{f�a@�~�8��"Oz]���Z�*	l[1(UW�ཻd"O���H� �pT`07cs�u�%"Op�c"�"3 ��2��#u��"O�<����-Dj��#Lǿ4t�k�"O�C
�~�pLJ����?� `��"O�i�Hր2�
�7+��g�8���"O�Ȳ��P1y��M��ꎞ�<���"O��BGx4`�G7w��$�"OJ���V5pX:��fJ7���a�"O��N�40��!��a�,ˡ"O�D��r�����%&{��t"Oj`x-�S�b�[��B�,]̘��"O�hU�=ok��HgN� ��,�"O��C&
MGA��K�Lk�r�xc"O��k!�۱x�i���EQL!1�"O�Y����r�H�6FO��01&"O�M3GМ���{t�F�)�*��@O8�%aB�-��Lj�`Ǉ*}JIH�f5D�Hct��'�p�֪ʦ[j*�J�L7D�p�%C�&q�( �&��Z��T��5D��� LB�i� 9�d��u �S�� ��5�Sܧ
+2pi�o�P2��3�K93��u��
�0�{��z��@B"ܷ$%^ ��H&�ha��ږ��TP�ʐ(U�֥�ȓ^�:@�����,0��`"Te���ȓpU�*��9`����/K)	�ڜ��8w$�`)V4ʚ�RAb�9 �ȓ|�V��1�կeRĄzr�����ȓL$~��A	�$����cO�W����Mr���d_2$���NʄPn2��ȓtv$vE�
y��8�ҷ��y%��E{����P�~Ix��E	��e�J%#�B��y���l�"@��N�ꬁ����y�戙hy$Y����V�YPK�y���>u,� G��(�.��g��y�(P>T�|��d`[%):(m��yb��1sRu�T	6�޸Y����y��v���F�+
��݊ ���y"H�;�6 �!�3�ީ�w/P��yB�]�!�d��H['qE��H��y2�'p!�`���� &c�����#�yb,�'3~���l�8���[P�Dk�<i�R.��|C�]�?Q�=K�mDt�<iUE3{f|ݣD��U��jq�o�<��c��o��!j� |N�{cpH<��	���a��y��W$�< !��2�PTȱ��\�*���[�!�d4�
�A� �Y�̈�"�!򤗠k�L�[��~L�
f�	�=á��Y/.�J�@����C��؅�yB�*��i@雜U�v�r�e��y��J"f(��ZCFΓ]0<T����y�,�7C�L@E
�Z� Z�D��y��q�dc�%�&M[!D ��y"�S�%<�Y�t�ڔn�}A񨂅�yr/Q�`pug�$�
B������ Hxq0�7�e���.I�F#u"OƐ� ��q2�G75ڌ�2�"O����^�o�,��IV"�f��"O I�D�5�J�N�����'"O�����I��z$� -�N�F��!�'���-{���#5NZ�XT ۅ��?�TC��?1��P��NFr8Ȣ�8H��C�ɡ4���7��{�0Ȇ���B�	�P�n��Pg�4��m[� ��q���0?1�(Y�~�:l�長{�8+3�E�<a$�:4~��я5L� t�d�f�<I��{�|,�W�Ȱ&F�y��`��m���O4�<��E���A䈷!ؼe��'���:6� L�ll8�,�p���i�'ND��W��=~��d!�&L�`4��c�'���2q�S�,x��ͣP>�M�
�'9��ro@�&4��L�K<�ۓɸ'0ܰ��T1o�����J���K�'_|%�Ҡ����I�r'�7JH�Q�'/v���H�E�<�Z���,L��	�'�j	�"*��p��ҥM_�9n,�z�'���!�.��Q�|���э1x҈�'`\�:b��}ښ ����>�P���'�>C��U)z�0�:�'@�dS�m��'���v� �+H��c�E�]��k�';���d@E�o�8�cO�ln��K�'�
1iK> @'�^#f#�c�'�xX�g(=v���C>Z���j�'��Y���G�8�nH�K�u��'s��k��.X֖͙T�Ůp5����'ct�C����3�0��AbS�h�Nuh�'���h�V�H�L�eB����'���Cb'�4=>�(�o8�B��'���X�L�a�\e��Ó�iFP@�'ab���N�7�,�
A��"x �'=6�Z门ep@�p���%j�%3�'=�ؒs���M2�R��%	�t��'#�\�W��+��!3�նI�:���'��X�Sg�X�,�Yr��A*�P�'T�Mɡ�и\Je�a!�>�Ĺ�K�|���=XH�S�#'�����D;����f�`��c_ <�p����~N��8�$D�,��	D9!~���e��)r:�k�� D�PZ�`O=;vxk�`Y�!�J�S�=D���F�0<��q�i�-ll
]��:D��Q(�c�X(�cjW�p�.�ڒ�3D�pE�F�C����!�(���2D�\S��-4��8s,S&\3�9��.D���`�Z�'����D�� �ه*+D��+�O�hT��;4	Ζ}��h��)D��J���6�`�r$i<a��%3b'D���ю���S挤Sx�iKc*O�AX%���t_@´�Z�,�=K�"O �b��(@�L8vˎ�!$"Ota!��O���#t��!ńp9"OH�$I	�O��|�7�9j��
�"O��z��O�VŃ�E��8���i�"Of���+͕sHܼ�R�0n �{�"O@���@ݦO�<\r�c��F4Z���"O��;���/Բ�����0 "��P"OZ p��I:m����6���I�Tٱ��'���$#v9��K��vǐ���D�/UTB�ɵR#�!(�A�D��q�G.u�N\ˎ�*�g?�CMJ��)���%y$ܐ`��SM�<� �\` /�CbH̐�'T!,Dx�"O�U[�&�h"���H�-s%n��w"O0yѮ��[w�Ȧ	��-�"O�H���C8E��bq�K�p:X���"OH�� '�=d�Ld��4D����"O�I`��/��c���6H�.��V"Oz4�D���#t��;|v%�"Oͺ��A��ԓw�%f���!"O��%A
�ib*ŽAlX���"O4��w��@$��[�H̠Z\|�V"O(�{Fh�0�N�kW@W��Т"O��&��9t���0 ��V;`t�"OJ��coܞ���X�o$����"Oi@���""Q i��nCV�#"O�@��aIg��M.�$3A"ORh�툎a�*\QaK�^(ʑB�"O�t�!��:2j�m�&�7l�Jѹg"Ob��'�
�=> ��o�D���2�"O����O�D��hI��ܨ0I�B"O`�Cbk���%�g�E&VՒ�"O�� Vω�zh-PQ�݅ b�A�"O���E%@g\��B��I�hm�"OB������UJ֊J�l��"O(�I�z{��J
�4�2!�0"OJỲ��;;
mQ��Y2d��x"O �f��<�D]��Nz�f�0!"O�uI�[�:$@�!�)ψ.�L�i6"OE�����&��P��1W�t
#"O��S-K�/�)9�%;�"�ۡ"O�ً�Ο�R���5� �M0BD�"O���ڞA_��)P�\�.��)�"O^�b���~
��c��Êj0��G"O"35Ā:,��ꌐ?�}��"O�݈�E�7y�@ I�
 �y[�H�"O��E,C+Z���#I�M�Xi�"O�����(&A��xBry�R"OL��U�W۲������(�����"O���w�#X�8��$�X��u"O*љ���O��ЋԺ�,��$"O�#Q&��NUc���i��K "O�i+����4��JS�̱�BU"�"O��`��%*�����@�B�x<�"O���� (�(����[�i�0%�"ObL��IQ�J�I�g��4n^� "O�Q#,�%GtaB��=�b �"O.�Ae�Ib�^m��D�~�cb"O��$�T����V�G�wނq�"O�����7H"�RSU'O%ZX:A"O�Ld�S&h�	�t��y{<��"O��2�]���	R��
3x���"O$���Ɂ�;%�Ac�ZBb����"Oޙ�M>y
� ���:��G"OHi�&!C�}N�]P��J�;�`X��"Ohu�A펕mT��C䆹Q,�\��"O� [�\X-���3���&�S�"Op�ꇎ�mƈ4zqg�1/�43W"O�q�C��D�>�K2�B*7�.��"OtԠ�΄!,D��[7�"O�ݱ���"�-K��^�2�J�j�"O@�:�f͌�@���5}i`0�"O�P���ϲu1��o�6X2x��"O `#�$�����[�D��(Ir!P�"O0Z�،ـ ��	�p0�b"O��A�{G���E6%'�I��"O� `�Hq��Z:)с\;���"O�ڎ[i���� �4)#��0T"O����^�
4���iuN��"O��vbـD�Ă�Ζ�Un\�@"O�l¥hG|vV+�nT�LŮl%"OpB���ԺI� �O�p�R�"O�M����|�=��Ĕ��`��"O�*5�Ɗ8r�e�ήu�fI �"O�iP��<d}���d��43�"O��S!Y�ܡ��,ީ�r�*@"On���\�L4�`�l�/9�ָ5"O��!�o��+����}"l|J�"O�
b��x��}9&k��"���"O�*׉j3��"i�6漃�"O�H�a��E�|1Ag���#�"Oz	�kTo{�
�&��(����*O��s�DJ
F�@���:` 	�'������!��dI�	��h"���'�����M�F�~�8t�^7�X�
�'V�k��9H̹�f�3Y�"��
�'n��ə=�"� J�M�F]
�'`R����i{�a@�/�|����	�'�l�y�H�:�-4z�i�
�'n��2t�-a�HuG���x�H��
�'�89wh��X
��Pf��3q�|�	�' ��W�}�D�B	��[�l�Z
�'��4r�_{�Fm!�N
&x��	�'Ҏ�Iu���^30�Rq �1 ��d@�'\-� ��)څx����NuP<H�'�$PiӉ�?7����$bR2Gr�,�
�'��T���_�'�( �c�K�M�*<�	�'���Qw��9����	Iv)�'�X���X� @���P�k
�'�B�Q�M؇s��]����N���	�'� ظPk��u4J��A�� `���'d��#C�s�����NEP�r�'��P�鈏{������I1��'���cu���s4�ZQk���6U+�'������� EZ&�#���
�'�aSA&�y"�:V� >���'� � 4T�\�Nݘ!�y��I*u��<���Z[y��H)�y�I�/rBޝ��	C�O�4�!�+@7�y����lyys��xX����@��y��q�",�CݻZu��K��y�o]�[IT�T#\	~��Ie�R��yrJ�*R�ʌ���H���q���yb�Q��v����ݑ~��@Á�
�yB�2(��
�$�=`7�X�a����y�
��4��QT��E:��z���6�y� �o��i �ȳ;��"C���y��Z�]��p���+_�������y2��uR0Y`�bU>
���$J��Py"�]��ܑ����)6���x���X�<�f$��3����B$PK`�H��HW�<���6]��ձuOT�~��,�l�R�<���*U��Ic�ᑗFߪ�0�)H�<i5�^:y�*u��f@���|� M^h�<�B�O6 i�r�ND;fl�i�l�\�<`A�V�`��.X/F{����GTY�<�+B�r�%�fݴ@Q���X�<I ��]�2u�0a��{�Ah�̒~�<�p��=��\JG���\2��[�.�t�<�QC�~1\paю0
�m����s�<� \���L�$m��3�߄O��8t"O��(ӳ���v��?�Z�"O.ố�!/ܜ�v�ԝRG�=!W"O��B�(��{c��(h)��g"Op8��5�
��̚�04rACu"O:�Sjy	�\��@~5�uH�"O��1�!�D��0��o��y2�Q�E"Ol��*N0(�r�@M��"z�(�g"OP�5O������G�Cb�9�v"OFA`�OZ�*�� r)0cAtQ�P"OR�BA�?B��"��*ŮY(�"Ozm����jH.\RgN�q���"ON�qA7h*�jS ���P�S"O|��7bD:R-�����(��qD"O�a(BK���2g�F8	.TJ�"O����	PQ6���e@2�� �"O^e�"Ƒ�!�2�G$]�n���"O*9A���Tu�IsF�J�\�݈�"OT)A���s��Ԙ"P�p
�,�""ODTq���6z!�r��.[���#"O6�آ�H�5>M�q/I5��h"O(̩f�
�s�x6L��.��&"O���œ>uQ^����p��5�"O0 � ���xŘ�<��[#"O��ȅ�W�9�@�҉��7���h�"O�xˢ���j{0�9I��P ��;�'���p�%�%d�A��Fε|Kh(�'��-	+�0a�|��6��+)$D�x	�'d蝨3�غY��!7g;)�:�@	�'�l�`����'N]���D��'ڄP�G�ˍ��	z'I1�mp�'�R�0��C'\LI��!p~���'$�UB��V�%�lQ�I�:fz���'�~�k�J�T�j5yaI	]��;
�'�$D�A�ɒX� ��W�zeP	�'_�=;T��!�|����Z T�(I	�'Yz� @��9�v�,����'���P1e�[�ݱ�hנ"����'��V[\$� u�.�k�'L�Pԁϧ=�% ��f��3�'E�D�Iެ�:̱��g�@�c�'6
x6��-f��IU�ѥX�`q�'���I	3����k��Y@�}��'6�X�����R�k A	�R�2��'��Mʂ�����5��$��)p	�'O $c�ğ�[2n�Q��I��p��'��3��I�u�jG�� HM�mI�'B��u�B��DJ���i�|h��'��MY4���$d�H�(��e��!��'���3e+y?�����2K:AZ�':�]�P���r&N1{�nۥ5M�J�'�U;��n�����͛&�ޠ:�'��� @���C"��;	�'�h����L�y�E�&H�
8�Y�'v�}�6�	�}'2�0F��d�ҵ��'i��!!�ˉVR�eC��R%Lt���'�,|�da�z�hxG��M߶9Y�'NU;��#4d��8Wj[/tK2�'>\pI6F�k������	p�4 �'�8�Z�l�qb� �(ҖURH��'��= ��
e���&�������'e\�
Q'$ ��ᝧ�h���'P�0���W�l����Iԩ y��#�'i�a��D���-P	�{���S��� ��8�m��?Ϛ��H��d���"O���gHyX|���T� �"O\�pD��)�%�f�q��M�U"O@��ZސTzr늏���"O���aߐ��|����
o��Q�"Ovx��C\�rH ��W��-}�Y"OJ%����m�hT��뛘d�  T"Ol�@ -Q�081�I�8���!q"O��9��;�Z�����640�e"Oֈ@�@�^�¤r�C�6��!"O�
u���a�����
&�lИ"O^�y���9�@�'%����"OF�#�`���݂��H�h}Q�"O��k���:��g�]�`��b"O�D��#_�H��\�����_�V�z�"O�4*
/� Qe�1@`�2s"O@!��g/#X	�N�2�0{�"O0�+� �X�FA�����\��a"O����cW*>{�e	 *߇"�|9S�"O<��6M�,bϮ� �D�p�:��"OT\{��=/�,�sl�"9x��R�"O����Ťw\��2à'h�J@��"O��PD���;L�S�_)gK� 0#"OƀA� E" 0����#��Y-�9��"O4�I��@�zZ���^�աC"Ob�Gᓲ;���� d�ޭ�q"O��ƞ⾜������"O�q�-X�+�0H�'i�&.��l�"O��`eK�w�*�+��Ǫ0Bq(�"O.u����DF,�ЅΥ8&��9&"O޸CS�E�&f�A��[*׃B�<����X �XRG�fdT��q�E�<9���aj>\D>A	N)�#�}�<���4m(�`� 	8.A�DЖC}�<)d���O��1c �\�pnڨ����q�<9�j�:*�i�+�m��E�iVS�<)¦�k��i�˜���L[�YJ�<!3����<a�,]#BNɲe@�<��D#0�$�#	:ySP���a�y�<�1WOF��R-!'@��Q��^�<��*̽P�q@��+kT:A��b�F�<awkZ8�-h6�/�^]�l�i�<y"A��O�|%qu#��@OPi�<�G᎜�=RQ�ȊgtDcE�Xg�<YP:	la��μ\->�fe `�<���ڿ=��I'ݰn�&= ��B�<)"���B`B��K�1� ����f�<9�៭k{�U���	H�؛�hi�<) ��#F`t��i���Z)�!�$�e����
�".��C�L�#�!�$1\q�p �d�#�5{Q.5v�!��Љ|�#�ы^H��vKd !��H��၅���x�%�r�!��3��M�2`=�0���!��Z�`�J��F�D%��+�f�M	!�d�4~�T�Gn��n�b�$�/�!�M�u$��A��+��	���
�!�d�$�*�"��,"�p25a5p�!򤓗c����H�3rhx �	;7�!��&q2P��k�h��2�>h�!򤆊8�~�8V�h~����J%b�!�D��a|����X.p�����M�!�䐴[�6iӱG�_�����C�!�d��e������ɻ(� �5d�oz!�� *�s'�I���r�;G;%"OT��0N��4��)�kP�,#��B"O�a`�N�E��9�s��
h��%�w"Oz��CM��ZG�5i�D��q"OheS�a�h�;��ѝO����3"O&��vL]�S���]���	�'�Lt�Ucɫ�͠�⃶�$�
�'0}X�l_'�<A� KI=39�A[�'��IƪW�yh�:�.ڲ-"�'k�H�3NS�3j�Ip��',>l�'X��٠��As�xZ���/%�:I)�'���G�>(�pK�O�T���'Wxdf�@�ÆJ�
v��'��5���"/��h��X���x��'w�͂���&*y�|A�BN���x�'�
i�8cƤ�4$�x�X�#�'S�|+$B۷e~�@C#Dv�"���' ҝ�n�$0ļ���
VbWf���'Z����*B�6iF)a���^t\�z�'G81r��;F�z8���'�x9��'�>� �(C�V���Q���3�a��'����5��L�FaZ�-����
�'�V�Xc�m�l��g����
�'� �b�5DG�O��ʴ��'�Qaw�:�0�R6-Y�B�ص{�'C�Ic���N(D�RT��5K�he�
�'猹b"M�Z�mZ�a�Ffjx��'��X���|��xbA�%;��q��'a>l3#,��t6j������8�|��'�&b%��$0N ��J>G'p
�'�us Lʌ3�t�2 [�,����	�'�ZpHS��H�Dp'��/�,�

�'������[�(�+��� �Nt	�'�f	y&�O>mi�	R!O�-�0�	�'U^�X�8��$֦�#�A	�'Ƙsc�	�v_r��e/y^<y�'��dK�cц�ps�m�4j	�'b�-mD�Iv���sd�%R��2	�'E��[w��)��ᗍчl\���'�$]�Ώ,4�6�aP���٩�'^� :�IP�R�\H�V/J�o���`�' �K@��'���q�^{�P�9
�'�6pr��'����9l�%�	�',4 )3!C�*�8WM�1uK�1��'�P�8�f�6+��$�3kŞfTH��'y&HZb#�]80��i*coL�i�'�.���ŕy+h�0���.Vj��'� �9E���vԑ�"h,�>�:�'P�}�"�Q3������x��!
�'����)Rn��1�IQ�> p�'�8��j@'VYM�%�/	�r���'��QxW�\�4��aq�̞o�hy�'x�x��lU�p�r%���E�/�#�'&�(��5۬h�%F�)m��T��'"�l�� �=�J P\�$!�'���U�I���5#'���
�'�2�{�MCb�e Ux]+	�'
�s�	�6r�2�4� �⥋�'���C�R="�^%���U^�	�'L���J/s�nY�#dD����'�>X�s��j:`�#�&/(�� �
�'��A�(Θi�4I��_ L,H���'�lXxV�N�_~��+�QI���	�'�rp�$IH`�����!B�TM�	��� �x���[@Ru���0�N�`�"Ov�Ң� �q���C/�>����"OZ��#Jw�� �(�/�X郓"On�×'ʪz�V�b��LmPAp&"OV%z�M��:�T��P+����"ON:C~I a䉛)-���"O�吅$�;]APؘ�'�����"OL�cbC�g.��K���'P����"O�0�n�}ԞЉ�m�c��|�"Or��S����$���M�<��9�v"O��(�[�|Pɢ��u��!8�"O�P���G
�,��*�<��@"O���5�V�(���jU{���3�"O<��"ȉ_��D�f A j6���"O��p֪?9�}0U��<,c���g"O���C퉩�,R�LN5f܍�5"O�d�&�ΗG^h�FKByv���"O8�1$�xu����t�7"O0�k��V�lPd((/q�hcU"O���آ ">A���>���� "O>���$ؕ��YfgÞY�*5s"O�4��K�:�c�"q-�Pi�"O"�6�Qrv�b�g�(s�Ҕ"O���faR1��(1AY�!�6�8g"O�Y3Dk٤4jl<"��)R�t� "O���S�C8�4�1$NyL58�"O�Q�R�ٯ�S��v�<K�"O��)'���4�	��9L�th��"O�]�!�Ej��EH�|}��"OfѤӭ��q`��wPh0�"O����T:�|���m^�Si.m�S"O4�E��x����̋�_J�0"OX�RU��(C�jg+�;G��4"O����Nå!����f��t.�j5"O&X�O��eM>	PqC�=jT�%"OpU�c��;�����>%2j�"OD ��E2ZU`C"܋ �a��"O�<Hӭ�$t |�[ ���ȸ�"OB�Q@(O��0�H��O5�QA�"O�����G�{�]@�K�!0e"O�t#A��}�Vh��h�%$�*��"Ob[ ��?"� ��%*F!*C�M۴"O�9	tc�\&-yg��6Ӯ@r�"O��	�eݸG�0�c�H%c�8�"O�X�\��� Pa��+�>Y�R"O>]��*�:ԩ���G�4����q"O�FжJ"�	7����"O�h�"KH(�<����r�&q�7"O�$:a�4�H���@+`��Ac"O(ɩ�U��ݳ�
�?��Ԣ'"O`�j��NvL8�bI.�L���"O���c����Ua�� �����"OB��ć�vN�A�R8x� ��"O0DR�ҤM-X<�3�	�/$�{w"O0�@�摴8׬�� �]�,��d"O�:Q��N
Q*�_�yjv"O4�*�H�)0����:_��L�"O�9B6�;B@5��rV��4"OĜضIU }�2�3�pm�%�"OJ��D�
bP�)�K޼5S�U�b"OvŻV��8�
�	�݆q2j�SB"Od����ʤA..�*G�`%�()�"OzA(B���0̲К$@[�(vpR�"Or|��b��B0��*q�Om���"O� \�C��k���:cQ�7iD9��"O��A�E�
�)�o�l���"OPQY��ǵQvμ�c$��b���"O`!��uI4��6�.H�:�"O�h����Z7��w�ņ~��̈"O�0#"��G�n��W�-\�h�"O\d����!{>nQ`İ�"�(+�!�Mm�r��� x�^�����M�!�C�rʼX2�
2?Դ@��"r!�ċ@܄�p5oI$g5T2�%��Q�!�$�JZh�㶧[.(}P#��3�!����\:��S�ŚH����7.�!�$_$dj�Y�OW)i@����\��!�$OW�x|9eb}��i��3�!��!��h���D^�Kp�
%�!�Ď���d�U�܄fMyҥ�!�D2*p�aH�@?W84y��ݪV&!�d�4���Pb�q:�!��ٱi{!��dNX}�Eb�(IRPcw��
!򤕫j�KVE��a
2,���&!�$;Ԝr�k��T�Q��Z0Q�!�\�25���Jha����P�!�P�*~-Bv�O�}S�\ QK��w`!��X�Rq�N�`2PY��Q�9!�$/NPl��W�K�^��03c]�wu!�DǷ/���d,�O�"����/m!�$�e��u!3I��K�rL:e�T�d!򤂎#�QCׂC#�Vѩ� �`!�d�+h;�B$�Ԣ����v`�@�!�Y9*A�Ң��=�^A��)�!�[$3�n�JG&%&��,�a̅3�!��Wd�(�%��\��m��T�[�!�$ѽO��=���٣a�@ēb+̋B�!�B4#_:���/0�����K�{p!��@���� w�+�5F���jc!�Z���m�8��A�o�!��'Z����ŝ(H���%�K1g�!��r��iZ&�[=Y�~���
;�!�D��.:�p� �ՌL3�KU�@�!�]"�0��[�R�f<��L��C�!�$Cy@�drD�N�H����,��>z!�&lg�b�@��r��P��j�$ie!���9n���1�ď^��i�Dɑ�o�!�DA.*��0ϔ`P(��55�!�=�}�+�u4����1�!���-f�6lq��	�\-J=���Ɂ$B!�d"��i��H��NF��cf�*2�!��.����,
 .Y�Ñ�M�+�!��]�&�`E�RuK���C�B=�!�'
�t�ĤaG$�����!��܉_�ޑP�-^2߈����T�u}!�d̼rڰ�h�Viـ�Q'Ȫ_W!�d�?5 "!��ˈB��@���ch!�$��J�h�`@��[�R1����/@4!�'��}"�	z����2��^�<�cF-�B	���l�����X\�<�ԭZ�=`1�/�8Fln!��U�<�D�f4𥳥�7_9��/�S�<�˂H�J�pG�����D�P�<�'XL�����PK|�RV�R�<��3[�qz�&]�E꓎�F�<�r��;/hIȦD D�pY�qnC�<飧�9B��"+�#�����N]v�<1�,O�jXp�̉-D�=5a�n�<� Dc3L�b���Sv��!�E"O.���I�+��[ԭ��"��"Oqct��$.fH�Xc�ۡ�xE�"OR�[�d��j���sĥ�
F���%"O���A��	4�4�dS�,��y��"O�4�f���@Aμ!ЩZ&!~ڸ�b"O	za�2$�r��Ǎ
���C�"ORqJS��(���T��c���""O��a��s�R���/8��-��"O(i9�fӯ	4(�0E$�$ �N�A�"O�d�Ң�1b�r8���6,���"O��&���fo:�s
��P�4��T"O����gIO:^�z����a����"O �C�_�Oy���$�[�*8`H
 "O��c�j�ł6	^0/3���"O֤ F�(&װH���m-p �"O����eP�K	��ӄ^�z��D�B"O���wC��tMXyid��Bf��[R"O�J��K��$��E�lc�dqW"O�Q�f��KZhh���0c�iPc"OX�cWgܩ<�{e�F}����`"O2��2JQ�	�
D�PH,C�r���"OE�O�N�0�*P�T��̻"Oޔ����!�fR(9	�a*�����y��Oexȇ��-4�N��O���yb̯g��-� U��A)"�R;�y"�4�l�7*T6�~`)����y�CA�D�c��(���տ�yB�X���X���"K������y��K��iX�́Dz�X�AK��yB@ �v%yV	 �:2Ir�";�y�lͬ_Ϭ9#AŁ�0v�,{p�@��y���=���넭!>�F��L��yB���u�����AP
4-t4��,φ�y2N�7u;n-q�c��+.��!�F���yB�D�K˰Mڃ@�*%`�qcH��y�c�-()�b�9�2�A��y��O�V��X�A��	��22l�<�y҆@�<P�bH �A���ξ�y�ȑ�Q�L�KQh�3�ҹQN3�y��ڙ%&Q�q�Z�)`@�&튤�y���1��eGͭ�5I��
�y��Y�H+����P�.�8تgk���y�i�',.j��V��R>Ap���y� �D�E�D(*�0�	@��y��X9��I5/��?�@�C��:�y���g�����
�L��H���Py���v�9����*� ��I�<I���KA���7�/P���A��<�B�
A0��J�|Dk���~�<Q5�ۧ>� �X6ˎ�]���&�Sz�<���K�jZ��iƌ��%�EHx�<Y��1eZъ��ސ|Oؼ�0�q�<������(`���N!���T�<�닔~v����I)�Pq�j�<�$-W9#�P`�A
G���ҋPc�<9q&�:Jd�cQ�_pC(D����b�<�d�M`�8� +A��*��'�^�<q��h?�Hc.��IW���3FR�<�w�Fi��mq6�[�*�:ّ6�z�<y�^�Y�-(2� �qDg�w�<�'Ԋs$6�r3D[�:�ʤ�e��w�<�敞TXJe�g퀵c�.@I�<a#��~B%P@�5�0��\]�<� ��A��$��Ԫ���'�����"OF�� 훍b�z�����C9�y�p"O�<�Î�2c�L��C��M
<8V"O�$��mӋF5�P t$Q ['JE�"Ol�aD&ʵjL)㣢t��1c"O���b�8Dr�HB�kʹS�"i�F"O :�@��&�x�U�L{̤s�"Oޘ��*�vA��Dп
0��4"O�1�`�M�jq�	0�<��"OH ����V]	�@,W�H��"Oި���T�q�R-"@&C><�
y��"ON��@܇ �p�dEY�"��9K�"O�M����/�H�X���{t�Rq"O��ʂ��-l�|�0Š�$,�Fp*�"OLM3'� ��8�/�<~�բF"O�����5m$n�2D�jrPQ�"O��1�G0e�`�D�1>S�T9�"OPe���Z<E�Y����!L|�b3"O�IUR�!�K�+@0�-�"OF�*v��8O7��;@�A�yOx��"O�;$EZN	<�㓫�=v�P�"O��T'�H���[aʘ'>�Ij'"Op��!���q�@#�3h� �"O��b"#7y��!���3,<�"O�(�LD@�2d̒�f�q+�"O�#Gӯ
N�u&��l�t8ذ"O8Z��Y�6A�;���f
yd"OvP��ńr�pE:2h�+Z�&("O�QJ��Ov�$����T;$�Z<٣"O��kW�,C0��7'HW�8;!"Op�EG�=�nA���Ԅn'P��"O���6�3
���ط��}����"O�(Q@aU:-i(�Qֶ5�:�%"O��b[7h��"�Ɖv`��(@"Oшs���ز���PQ���"O,Yy�ㄔ��ܢl�5-�x"O��c�nC=�$��s,٣1B��)A"O���C�We�0��*��W)n��"OL���� 1(Ȥ�A% Y�pj LJ�"O�œE!!$Nё6�QaG���E"Oh�"e�G4	?z���M~]�"O�-XԊ	�)�D���W�1ʰ"ORE�V�خG]���!K�����V"O�Ÿ�bѐH� 	 *��o���S�"O
a� ǦU�$���Pd��#"OFm;gi��)�%��Ѩ]�ĵ
""O�@'���D������"�"Od��5�d�P��.�`���"Oz�y�i��SQ���R_*`)�Y��"O�}9�\�j��#��}x�Z"O��4�̆�~��)ԔY���"O�Qم!�
�� (�<�2,�"O�I!n��:��89ņ
�v��"O^��eр8P&m���3C
���"O�y2E�I1E�KP�ע6<(S"O�U�Ү�Gh���E� G2�8��"Oʵ#��Gn���/R�f)\Y3"O�r7mI�;W$xH�'N�|��Cb"O�Y	A �s�e�C��	���3S"O���7�}|�y����̑y�"O�9�r�%7qR� �DÎ��@�v"O����8XY
��%��U�}�"O���`�˂*bؕKԤY2H(�;�"O�@ۑg
�= P\�I_�Z#�\�"O� ��B7*�,@z�������4y1"OȚf�B1!Ǹ�����a �e�"O�{%˒"�M��sW�[6"O$4��F���ɰ��_�`9�V"O�ؤB��N�\����@�o D�+s"OXqZ�,~�:�ja,E�d�YP"O�\���T���GaS,0l��Y�"O�� BH�;>e%!A,$�!��"OpY[��r:����Ņ<wr�i�"O4�C�++c�� ��-�u�$��"O�$@��O>h�>��"LTxs�"O<�&�	��K+�*b$@"OЙ!DE��q��e�s�=r\(#R"OL0�S�N2md�s,ai~�`"O2�!t��5)��R���yW��KD"Op�Ԡ�M��`�M�F�a�"O��)��}���F܌HR2���yRLS #j� r��G�@�J������y�͎���yz©�� P� �Ѡ�y"#
�0�.}�t�#�r�
����y��Z? ��Ui�d�$1w��d�D��yB���(�pM�cg�/p&�*��X��y�_,4Q�HG����#(!�y�?6||ztW���h�c�%�yB�Zz�&�A@R�o!,�Ї ��y��T7N��ܸ%�>S:f�;��P��yC7f\�h�ˉ� j00�eH��y��U�3�P�RDf��!���y�>Z[R��7�Z�I�l�@���yr�I'y
:|!A\�I,�shE�y"@�4!|�D0���Fl)��]�y��ҕrN�	t T9M�Dz.�:�yB�ۼd\� �c%��
�mpKқ�yB�,P����˗Y���%*���yb��(9�&(����K^�h�uo��yB��$�� �r JT&R�!D�G��yR�P)n�b��R���F��yb�B-��`CƴAczp�&��y��I:+�`2�%[�H�� ��
��yr @�6���k(LC�ԡf�J�y�ĲF��$y�#�����z�� ^�<�v�@�. �a��uB"�P�<��ՙETd����!�)��)P�<1 ��F�	�@�8�����K�<�7l�:{|$y*AK�HY�u��E�<���.y���IV,�C��J �}�<Q��,y8��!ߣL^��*f D�<U!ɽB��aC�ҚNST�B���[�<�gƘ�O]/,lh��R�~�$�ȓ&���c�L�&5�Lq����꜅��|��H`�Ĺ�t����[3W�(X�ȓ�2�j� �D1� �A,o%��VDJRg�&���`�#ߥ/�湄ȓC6lܪ�푸(_8���B#up@e��&\���q �5�� �AJ��ln����k�L\�VFW9FZ�U�6���n�耆ȓO�
�*�m(�L ����*�<��ȓ;{R-:�M�]4�0��H�,��ȓQ`x����|޼����g]ȑ�ȓL
�2�+ͷ /P����O)#�I�ȓ5�V���(2�Ρ0'$^C]H\��,H�1��B��vܙ���-K ��ȓ.ȩ�b�X�H1p�J֖/Y�9��Ig4q���T�nLR�K�B۔9�� ��S�? ���'`�4Ri&���A��Bf"O��S��ք	��1�n��(�"O�i�nI$	a�d{�A M�"902"O��(��L3c�X�a�N�VL�Xh�"O^<	��N�Y �%:�L��Y<P�A�"O�t1��Nت|����,c'�x�7"O�-���D�d�Ҥ���m���;�"O����W&_���0K[�o���1G"O�,zL^�J�F93P�)7Bi�"O�h�'d�1|�TR7	�T�� E"O�q2� �J�y�hG�v���@"O�ِ��;H���K���\�F��"O����e߯pne�d�O�z��L�"O�\"g
�Br242E�w��5z!�ݿCI:���+
m7��Zc�ŝ
�!�$����B�4N� q{�c�!�D�V!U�o�4 w4�{�"G&}
!�-2����w�ә]dq� đ�V�!�$Z"!T�Sg�gJ����m��C#!��#ӠՊQ�_$� rLX�\0!�$&
x �x��AF`<҂J�bA!�dJ�j@�8� �HtL�=���Dv�!�DԳ &\͠7hH�q74��C�Sg�!�Ā��(� ��X'4#�q��$(�!��K�����M�'D��1�VƆ�E�!�Ā�l ��Z�J۝9�\��3!�D/&��҂��2,���	�c�oW!��R	! ���Ռޥ@�1WLW�-F!�d��_����J�O��*P2VB!�d�61|����3��R2#�Q>!�DZ���@ U�+������^�!�D�46Dt��B9��yk�� �!�䇥K���G-0	�tI㫊�P�!��tD��-i�<�c�Om2!�w´㤎N��*�*v!�d
�;r�<i��G���3��T9d!���?�Խ�bj̄��ۢM�(p,!�ɺo"@� �	���0AC#P0`!���:O|,�����5U��9�Vh�\�!�~�sD��?���uA[�5�!�d 3�^���08��/���!��L#-��%:2�R;	(>)�l9:�!�D߃z�J���bK)Lj��sd���!�D�"��� t", �\ɳc�mP!�d~H��AI�<��p�)��J!�D�9i�wEٔ����2a/!�$�
h��I	���Q�04��֢C�!�Ē1*�*0k A�!�d�$g�<l%!���%8� H
f$�+�!�BH�!�dKm�`�+��7`��%2���[�!�	���W��"U�$q
1GD 	�!�D'C�u�#.w�����}�!�dQ��8�AO�z�6�)w�&5�!���lD2�ç��ab�0Af!�$�ޥ���3�J�o�3ޞ�Y�'�&!�,�:��"!2�p�
�'x$1�ᮕ>>#d�PFW�D� p;
�'G�2��Ų��y@nԱg��[�'B����ǲM����7G�h���x�'�V(�eK��l'6aӦfV�NbhA��'y�����-Z(�P��Ţ=m�Q��'��{P瑮y'jQ��鏸2�Z�x�'��a��Ǟ�K���f�+2��(1�'/dM
�P�a����/��R
��� �5�/�$�,�s��Y	ZZ�Y��"O�0x�'
;?T� ���4�L�5"OtA����QumӏK��F"OD���ȭV��bl��O`PA��"O�	3� ղ��釛mo8�"O�Lb�g�:X��A1
�643T��F"O�⑫F�J���ah�/�젒"O�!��&
xJ��@�{%�D("O�˔�<���PsF��
�:7"O�,�&�,h�A��
�ͺp�b"O<u�'�5��1P���r��4��"OT�%�8Kl)�ÁW� ��8�d"O ,a]"$���A���j7"O��ȡи�`���(���c"O�)4F�0D�����)Q�L��A"O�Dy1.]40�~�)A+ �R���"O����΍!k�ػ`�� d� "O�p!d� $��P�\�;Y���""O`a�SJ��Tc��bHFY�"O�Ijp��lh���T>V��%��"Oh�^	�4R2�Ë ހ 	S�<y6�Ae8� 9��x�h����y�<)���k�t�� �مPM�lҠv�<�B@�6���&�RY�Z���@Z�<9V�-1SFIa�&��{-��QcE�X�<�S�6���g��U��}q��T�<i���7M�61��A�� ���BM�<��D4�x`��1���Pg�<��`�i���_�`�/I@�<���t<`�� ��E�r�����y�<	1�17����B�傄�s�<�4B\��>��x�̝��P��pC�;1�VɁ&N�����kK1�JC䉹G<�
�昏'�@{��˯M�C�	�[��\#�Pj��C�l��v[�B�	#F<,���@(S�����G\ �B�I
>�)EeW.=�`��ˇ��B�I���A����I��t��L��C䉂~#<�J�a��I���f����C�I!d&Phc�2�p;�ܿP��C�	�Q#8���e�\V��Hr�=f�C�	23% I� �:G�����X��C�I�v����f�4^�	07��j.�C��#�0����JcN� �B�$�B�	�ke�� F&�lv)����v��B��6m+�\�Ƈ^�,y: �q)dC�	�E�!���ѱA����Z9>��C�I0^��3���:���C���"s|C�	$](и"'Y�5.X�a��O,[P C�.�\m0�#� ?t�BuIےZ�(B䉨)�H4�s��
F$a8燕)1&B�I�8]�� �̌��8*Q�֑N�\C䉺B���)���l༰��Q.3u`B䉰Jk��3�A�(W;r��d9?�B�I7jd�[��Ȟe@Q���m��B�	�de�\C�h ��dŘA��Q��B䉴Pޔ�#gė�0A�����(hzB�I�HdV@af)��4�,�9��ڷo>>B�IZ>�1�I�eU]���X.�jB�I&�48rP��z��<��׭<ȊB�	�-�4x�4��X���r2��a�tB䉬*�IH�K@�Q�℩�R�'VXB�ɰ�6�ӗ"�7��dK�N5!�DB�I�q&�`�"FT�?v��Y��D3(�ZB�)� Э[�j* ����(�dA�T"O�ш�b0�q�Уԑ5��i[�"OƘ��ΌA�j@R	�٠а"O�<q6,�����R�H�E����"O��h"�+;��1��
!�l��t"O����ۜ$����4c���3`"ON�`A]�[W0�!X_������b�<	�O�*F�8@a�5��ڳ'�f�<%œ�{	�UA���=^�Ų��\n�<I4EJ�}�9ѣOA���j§Ph�<Qt��vf����ō~��M��d�<��O\*4_h�Yr/���<aĘX�<��,�< ���ȼ��&F�P�<1FOW=|��Ԩ�'��/�Z��)�K�<Q�)�-�����V-�N�z1�O�<	��[_��U�%�M�Ȉ%�J�<A��;=WD!�unZ'�B�d�^l�<yC�@�NLr��!���pĉ�i�<��Cyʎ�Q�� @���8kJ`�<�Հ��l��,�l q�������R�<!V�;|Ɔ��C�tU�y�U�R�<��Ⱥ!�h�`��W3+���2��s�<���b��!���zxB����p�<��IR���N�<+N�K	�R�<�G��SP���$H�u#��S�!Ht�<�2O����F��
~n^)�f�q�<I@�]e�Q"FZ��U�Aj�d�<����,.�V��%We4�ҁ3D� ��
0~��Q����ö�-D�l�௔s I��)Y+4CF}c�6D��j�@
<�H�r�� ��S�C5D�PQ6���^m�C�oV-v���Z��5D��9ANG�X|�+���� O�X��,3D�T�������B	ݮDKWd2D��
׋�`mR���8��ʖC/D��YDъF�d@y��K�`9�1��d,D�d�h�";L(`�%�O�r18�>D��s��L�(`@T��˔z�&�2�!D������`�:̀ࣔ�W���5#D�tiw,��RS�!�n�&#���K D����ǉ1������Qi��B 0D��¤��@;Xʇ�O�9s���#D�D�I҄"�ʥ�uQ�f����H!D�  ?�vU����p��,a�(!D��wgԜ��; A[�I�F}�I3T�D�0*C�Y(��.$'6z�"O��R��"�����
F
M:"O�\�gKT�i��?U#�|!"O`HtfƏU(���0��%<.x���';챙f�J
$jp�fL��@�h�'PJ��WB1Ld�e�J$ ����'!�Z����hp�1+�{^���'��(S`i��
S�`��m���*	�'�`�{�#� ��A��N�k!����'R��BbAA0\(���e9(}��'� 3�Y'!
��V��
\��ē�'�9SPE�:����H�6$/(e��'�05'��k.Ԓ�o�_ބ��'i\�8��)pB�n%��A��'[dg�T�� ��'!��`�'�P*��R���4�`��6z�9�
�']\x� �B�՚P1ao�YzV�{
�'F���cb^�Vc�+�O�O
8�	�'
�K%o�828L�WeF�v����	��� [4� $�5�s��1"�c�"Or���ə"X��e�c-S75�d�1�"O�����y������c�p��"OF�K�d�4��ɘ�D�V�h��G"O�CI ,�4r�Cնd}��r1"Ot�)���MJG�Q:0n���"O�a[��9oR�;1a�3O��S"O�Pp���	ĄX����WG�DB%"OƩ;�b������=%�
�z&"O� 0���x~��	��=_�:�2"O��s���j2r�bA$)|
A��"O��Cc'�BeT�!3LɾI	؜y�"OHH2&�~���sWKO2�����"OlX��F�
�HH�QJN�v�by��"OF����/!x��g���&ЩA"O�r��4B�:�F	|l�ͳ1"Ol�����qV��Vlm��"O�4[�A��^�lȨ�Î�"jn��"O葂�R�&7ؼ!���N,�sU"O��ʑ�l���	���2L��=G"O�#�E�p , {�U�^zR�˶"OHy��l�8Ƈ�`C�<�Q"O�@�%R�[�hU��G6�q"O������=V� Ug��)[���"O<)SPb�gtm�2g�X��g"O
7�;J��KGWr�H��%"Oh�Y���>/���Bv�@�K�~Tx@"O���A�!L�qU䑊{����"O�M2e'�<�R=��e��� 3%��|���	�C�x�d �8[<;u
)���)�O ����6	���:feG4@�6�Qp"O���P �&fA��Ë�x{�O^��HMo~�  &�tܒL0�'*Z!�D՛<֎1Z���#=ZȲ����/�@��ȓa�� ���V&��8�G�!�~���7 t*1�H�w�r�$� G-�l�ȓ�4��e�T1�hYWO��<,�8��~�AN�R��a�SjԉRSh���	�Gz�	�bײ���+G̜�A�  }��B�ɚGg��A���.�H6�%,P�B��-��c�j,�Vl��@��lP	�'P"��!KØ=� L�b�9#�'R�qRDE,f�y��K�Y���
�'���j�Κ�g^L����S{�u��'����W3H�#2o�P����'������2
�*�@<JLP�'���;m>��÷FUv���O˓�~��ƟLF�4`���[@(^Ě�S����yb���
F�`�q�ǷO�9�S!���'M�'7>9�B*�#E�J��d��{��I
�,LO �'t�d�f��x��.�h�@;T�>I������0�0�8�g�O�5J��Y :أ>i���է+9���6'М2�.���H><�!�$��a=2 �6� 
m�DM&�J�v��+}��>%>O���!�xİX�P�,:�Y��'I�I�^�q��ǃ4Rv�A�mW�c�T7ms�X��>9�$q�%�T���ֆ7k�Ї�	M��\n(p2��}nu�4%��:t�����rFH�.�� �so�(�$��������󤋵.	0�B��nT��oP�=�!�$βq��@��͇�h�aV$?U!�$�8��"5�#a�T�#ω��!��=`t4���E��uڌ�oY�I9!��H�q�Dц�΀��բϝ<}!�� �l�'a�#O��1��Ӡ=�l=j`"O"l���G�:0� ���	H�>-Kv"OQ9���h�����*Tuب��"Ovh[���H��Ƙ�g�`"Oڅq��Cz�^�8PF�$:X�e� "O��§ �����fW�K�H	;�"O>�q�2<X�0�Bc�?nԮ�S"O$�*�-$�꒢֐(���>O��=E��o��C��	������7�y� ͪy������ƀy�&�ɦ���yr�;fc��+��Y �"��F�C3��<q��9^P2���^<R@��(��D�!�P@pت"/!,��pDݐjV!��9HbPBB��#�%0�O�ay2�'.��'��-�e��� �eK�:��)������G{J~�H�%*�N9��%��<jDl���U�<iVC��9�r��#NS�n2(�4oUP�<�G&��%��dr��� �ʍ�f��J�<�ACX2X�0U�D<xB��H�<i���F�@P�DN��,pR*�O�<�p� �}K�a���;��-��fI�<1f�4V`x"���qlb��V�TAy�>I�~S�@�r��3��K3`�7�8ȇȓ,�8yK`�j��D���4DVЅȓ|��X1�ּ+��Iץ�����>��'^a��!F�E�����X$;j���h���y�Ӳ.�"{�퉾f��	6bW4�yR`��oQ��Ŝ0^���d͚���'�ў�����}��:UO('�4Ī�b�� ��ɩΐ�C�V1��)!F#P��$B�	�vFh����>Gܹ���XO��C�������_���9D�E�JݚgN-�I��4�?�N~u^3����G5PE�D�Z�<��O�"��)-�k(��Ӥ��R�<!@M�R�@i1�@7DU�i�� CP�<�g*�� �L5r �F��B]K@[��xr��N[�I*���X00IB���
	�'���Xq/�"�Pɠ�אLj&hC�'�Mۗ��?m�y��ͣ�ź�y2�'�Raؑ��Qb����?W���'�r	bJ��A.����I�`,B�'����p!�m�d��`�D�$la�'<��wA �UWȴ��N@�\q��'���� ���������QS/WPg��<E��'�"��wd9/���w�9S<R�'yj�"��P�:eI�-R��y�O6��$�.0�y�Эf��=5Ě�w�!�D�&0Z�G��(4�x�#�H<!��8Y�f�PA^g�RM�F �I�a}��>�5f�Uu��9 0`PE���x�<��J�{�|�sd�4v���A���y�<A��&\0c�j��K�l�ԧ�t�<�uѮ	�U�fa>R�$�G`׭�hO�gy"�O��$�/�$�
�I�d��*1#ʽ��C�	0q>�%{ՂJqar��FR"p�HG{J|�(H	Ul4q��%�a�`��B$�O˓t�NU�׹GU� ��)Q6v Ez��'B��5�ѨM'������H��
�'X:HpE&�.7�^��dJTNdP�4(����%~^>т�	BV�D��|*!��6"OL���g�s�6�JlH�h01��qމh@Y,��c�Y/@�D!DxR*^`8�tI��;$��e��|E���1E D���f�S51¼=�bkk�)���3D��  �*E�np�	�H �U�BP*""O�P㫝}5�9	����$���"O�2�-ʻ_:¤�7� Jèe�dY���A��o�'O��a��/{�z�ВPTR@y:	�'�ؕ�V���F�xmq�(8I^� ��O
�=E�tI?��0!��	0N���Т��'k�`V����A2���V���K�<���cџ�yR�O��"~Z,�2��#O\�9s�yi� ^z�<Y�@BR��Y������hO���<��nX�A�X' �Bh|�������<9�;������Z�pLxtf�;��x�_�"G��%_V���I�+��O2 h��IGh�BՊ�*� W��APLP�p�1O~�=�O��$�=�$�E �'�>)P�l�9�!�d�$<��� �"�`y:`I��l�!��@�]�T軂#ި �����(�<�!��+x�;�L�{���WW&:��IEy�\��$��'�� ��χ���y�� ?�E��'S�T�2MF�+�����R+L����';��3"�@���5����݌pi�'%|�q��]� \����|P|��-O���Xm�4ب�X1w%�T��@�%�ay��	�L>�sF�%,�@,��J# �C�0M	��H"/�SZ���@� w=�B䉸[���E�({Ȕ���mK�T�tC�ɂ9���D\��v�P,˴�B�	3�t�
�@��$n�h��Ό .B䉀~��a���F�S�Jp��c��L�B�u������yx�VnХ*~�B�I[]HԘ1mɏm�R�!6���aoTB�	..Ez聵%� G�õ�%�8B�I&`؝
p�K���A���hB�	45�*,�qoB� ������`Y�C��U�xK*�=88�[r	̻1�|C��#3d�r�`]�p��Ș���}�,B�	�G�Zy#�
�
3 �754C�Ibw~��
*��6��]�@B��'g��=R1Mȅq�:9�DU$M6B�I�56=Xk��U��*uh�0D�4B�	rN���1e�4�B�c�*̛7�C�4v��<Ѡ'�'[<���/�~�C�I�AL-�R��38%#˂9�C�IC0�����,7L8��`�f/�B�	�-zL���!�R�Aa�L�jC�	�H��६�D=N��'��s�B��������[H��(��B�Ɉ������oa�P��M��fтB�5�jL���©$��#�`�34�C�	�<��xHV)�<~�@�P�*:B�I=Ptp���ظ`��<z'��}�XC�	�q8s-֋$3@�0��H�o�VC�ɪ6�ʥ���S#f���A ǅ\oHC�	.Z4@s��!���K�!�C�	�i��B��>���[����.�B�II���R��N�nmp���f�B�Iiؚ��Ed9N�R���D+:�B�ɲrNN�";�(��t�6wbC�	,<�� ���شU���� �B�	<Y�*��䂗�@��Q�(�0w�B䉦s��Y f���\����J�B�	�Z.�� �{�h
E#��t�8B��y��jnO$�lHb5히;!��釫�)a�����L���,�=�,�Q0f�?|���
�'�0u�v4�ě�@��s�\ �
��� ��1MX�h,�IFW�Z�fy9�"O��3uoҤzwb0��.��	�p)�F"O�4�	R�\�dpj�䍉*^LZd"OP���aS�)��+e�D4h�$!�"O&��T�ɴW�⥲b"�r}l�!�"O޵�P�@8�Ԙ� ­6N��S�"O�h����9u� ��OF�/NN�i�"O~���↼5��,2�5]BTH�"O����js!R��el6+�0
�"OR�2&�`�j�a���$��II"Oҡ��L��{�����˪:�H)�"O���C��=�Z�����&Q�J�sB"O<8ac��lX��e
f1z�"O*��
��xv��1H��%z�"OLi�"��n|���c%�A�b}��"On���,�j}:��re��l#PH+b"O�p��h�QL&l;GAˎ|�e�2"On���֍S�s�n	���Ahw"Ovx�t���*�iڄ�X�%�"8h7���c���'9܌�z��O��(���L1?�Tm��툭Fs$��	�sG2H@��+�@Q��+`�l Gd���I;W>��OgZ@5�B6Q�X��'�����7J�6��N�o�҉��t�.ճ�X?��B��V9':�ʷ��;a������O�ff9�s�ê~�p�;&JL?��Iܧ&閝K� ڍ\���1����E{��:d�,�F�ע@!v��)g@�IԽ2�IF�g���v�/u�J�ˀ�S�P���5B�v����L>�� Լ,���:B��: �=
WN˦���%�\�J\�7���C�کZQk���(����L4v8a[����胈#��d��46<X���9��,�t���wҭ�䏙�Ryˣi� M�&\b ��I�����v��	��1g"ӼacJ}`dM�Oy��l�8���W�]j٢��'�p�	���ąѱl	�ip��	
H4����'�J\���Yab���Ø:|pv����l�I�L2���O?1�0�h-�В�%�w�:��g�:qT؂ƒ|r��vD��fBO/=TFMGR�|� ��1�O�Q���2�����k����dA�Kw$�8��'����Ȼ���炍3�����@��:k�حۀ/�m.>���nă1�|�������z|�v�
o�Xx��ֻi���?��;u��Q鞟\s l� -J�b�Z�!��c��ɑ����
ը� Fɕ1��d֞ @'?�[!Ϝ�^�D	'Oŧ<Ht3QC�;���z��Ζu�NH���5>>#|�b�&p*��$
�,$ 4��z^���F�I��ؒ�O�}ȳO)'3<�$>7m�>��� bS��K��!�d���
�F����=q��ű��+�����*	��+7�[�(�|���?i� ^�Nʘ@�w.�"yp�r��= �|���2�W�T����2'S�S�	����+v��y��+=���#�
�2�� ԯ	�����<��T��LA����� ��=�� ���K&6��(ďZ��?���I�F��ƨ���Q�O[U͜�T�ԉn��\���6h��u	u�H K�@����O��U�6��WȖ�4��9E����5)ѴB�x��r�w툄k�)X� e��ǉ-/�i1�.�8�?���зD�l��BB�T�D�-^^xq4b�����5C"�x���eWD&��2��Z=��x"
֬]Y��H7P"|%�kƲ@Fɂ�+�4߅�j�5�\�i��!p#׶\i@���^����f^�<fM��y�G�<{��ص��H \7��q�(�
�b;{�YC�s`� aw�B,%%���7�I$@8�&�s� ���Z�y�yф�(7��h'��kp� p��٣[�%那�sZ�ܢ&W�\8�$K�9?�I��뛟 ��;v(ք�~b��P`�@�w��^YY$J�#��y��M�x���8���aI��k.�Pc�t�7I���xu�d �R2�9*A��8p�*FL@Ȧ�3w���J�Y
�g��YϚ)0Ac��2D@&u�,=�c�@�g����]�z���a��^�d�K�b.'���'��8^h �U�F?D,���jA
~���FX�|�b��%���"lF�e�N��C!bح\!H���.R�ࠐ��;,��5��j
\�R�����#���,_&F ����m��DK ?�y�QV(�f�� �Q��?��#ܖ�r]��LG	�3?��,G���R�٧9�0��?5P��,��,��mʃ�����U�/�J��"�&?�4�#���;?F��l�*,����"��wC�B�ɗb<Qbٙz#b�KwD�a����,ЋO���8��ȓX���C���F�0�o�
l� -h�h�6QD�adA@��f���ˑ�c��)�%�C�X�Gi�0V(��ڠ���-��1�
;H̼��ǃ����-S�UJ�:��z%C��	}�����&b�z��S��+P=��Ɛ 8>�H��kݼC,����}`9�C���K4�ۂ* �/O6����	l�d8�T?Kd?@c>8q���"t��1eC��C��]�t������z8�D
�Ck,!���>L�a�3gE) fGs���s�ʊ�8��P�0��J��>��`�P�HO��EI8C� ���ѣ ���v�A�\Q���JQ<,�b�H jSl�%��F�
���oѡ%��$���4XY��#Dd@"n��9���p-j�o<HF)���XԔ�����z �ij��	�Mǐe!$aR����hQ�ҥ^"����B �z�kΎ� I��B(H͂Et�����X�xbڨ��T�矜Oj9���ؤ�HO.k���Fh���cO�$����&̒�1�@M��@�'#,|�0�HL��,�x��ӛ	�m�bG�!�ΰ�1���<as�n|����AN�K"�]֦mʁ @�+���� {M����Φ��Ri@�����$�;-o�h�����/��6	���8I,���S�? h䒱��<ULLp���:*�0$���ƮJ^�S��A�옄�2-�l삑�<TIPHѮ�8.� 8�8�����V">Dl��A"�~��C�'�x����1oH�5�Q�@Wqzy�s�Ҹ+�.�������I�D�|�p�-��c�����m�([u�">!�h��K���6Tu��E��3���2&�|OH���OX]�1�a�S`�I4��rs��i>n���H!�Y$Sv�#�eG�:��
`�$ŀ�c�-8T!�l߷l�t��l��O>����5KZpABb���qS�� @��D(Z0�-�����X��LRUQ2n9�]`d�[�ة�+��W`1�փZF08|�u���#Z�G2:6��8�ri�7B�98�Z%�w��\՘%�A��'|&���c�5|O�t�'B���t�d%M��w
�;$��k�ͦ#OxH����/z�ޡ; �;��`�DG��ިv����Pٺ�@�/wJ�c��Y�?ດ��I�x��1h�@�c]�
�4P���(�ZQZGC��1�1r�(�E�,I���U�v0xS�i��e�h�J�'�,��1��H�1{۟ظK�>]4a���$��ۤY����ӟ4�Y$�_$HeH��#eԝ+� �!�.�A�a��9W�|�%�^�=Ӯh"�#��wmL5�e�_����
& ?|�0w�աET�t�5�>ғV�4M����^��E3b�7D�hY8��&n����k[�$��A;ԩT�>]�V+�=\��E�5A�vaX�mR&AG�}Xt�_ ���p���eEI�^A/�8��'��0b��C�z����RU�Q���V/:��꧈j�zq�E���z��CA�/}����n�Ӻs6)�5�M��4|�!	��G.B(�1c���4\�<AaJ(���4]�8Ei�'�x�b� sPy�k� ��a!OƍV
�l��>��0�Вcwf� �I'iJ,,�B��(i�`�(%�i�"�`@�C>n�5�N���V��0*pY����`>�}H����.��4J������;f$d�p��mN���j�!�r��f�7"zq��A��(�(
�,ϐM��ܴ$~\h�#���Ѣ�٦;J�y#b��E��$�|+B�F�D���ƭ8[3������-w#bM��Pi���˥��i���r'bVR���-�;_=���N�r+veh��k�,t�ď�.b���ʃMyQ�CJ�*]��AVp��ׇ)��Y��%-cIQ�IO")xe�2ɟ&�Q���,*J�8��"?7� h} ��U�ɟ�b\�Ć�I�%�vg�?�u���<p8�Ah�v�i��"ǆ����ӀB�AԾi�V�� �֣�YZ��@�k���B�l	"�h��`STn��l �Z��h��U&K4�T��m�(5H�a`Z,]g�TKq�?H��:q�i�P���͔n!���G)�D�.�"	|���Źkȡ�&�x��@�9-�\�oں����4Ü�8M�XE��u�4�c��M?��:7ʐ7@�͡�6����e���w|�$IS$YܦŐ��p�B(���%h��1.�r��L)B0}� χ8� ("�䚵>�^���R��b����!3O�M�s�Q<}� �G�
�:*�$�6;�R�0��5��K�n�#�\�A#�"�H�[�E>V��4"𙟔���Kx���9ԠR)3/rh����"� �W�\�y�����샹HR��0���X��4��I��l�(����ɍ������{�𕊦�OT��p`*P?^���	�cZ��*ģ�����["p�j5#n��d#�DX6��j{h�*E�3(Dn9�A�bJb��FG�/�MkfE��Z�����!yJ&t*Q�ɵz` �KN8�7����x�7A ���
�Z�:�]��H6-� E:\�ɕ=&E���҉a�!4��4K�R�3�$���2�Pf�>��$I�BqJ񌚣u�ҙ���l��}�0��?�*�ag���x["��H��� g�.p�r�T&
%��=!qf��1��D�5'�Gn�x:�aP1(þi���2�H�L�	�"�)oʅ����?%�U U:�6��7g� \$�5Y�N#'h�u��A)r%�Ep/O�F�+��B����0W1a�EW�4�ʣ�}#��C��g]z=i�ϙ#9p|��g�߯�j��7��1�+O��P�ᆛ�T�+����k��c�EK�'~��Aʔ�ո��戚05^�� raG��D��j>{åK
!X��6�S�V��lX�R�9z���n�05q�iJU�*!��� ��p<��E7%^�P��� 9y�C<VhcrAD�'n)����t�@�����������<�)X?�9�c�L<�����FE�N��䃞k�z�
׍sv�!��땯L�je�>La�#�۳�PݚpD�"P�@�ۑ ��=p�9��K�	E�8"�딼Fi�'���b��/3��3�P�NE�*���'�&tyEH�� �r�� �U�d� ��
�V��p����HB"�!J�pE[��z(�@�Ǎ�$0V�D/��$ɐן&���{��!�GB���uG(@?v��\�T��=KD02#���M���I�����I	Cj��� ��{�ZY���:1��H$&��u��>d��ōO����7���
��0���k�Z����ڈ|��H�4:l��;����w�2�� ��'�4H�m��V38%(��;���P �B��0�#ӃR����H���2@�'V1<)0��ށ:�����C:��Q�}P�E�W��Y��lk��3@��g�ٕ{28�EhQ 0���{�� ���H�I"'������_�3a�<"�"ҁ�f�" �� �<a��{2 � %��!�_ �C��9:�HS�'Oꄈ�g�nM`0 c��W�:�X��.ړ:%.ЉĚ�����!L�t�� �L,X�R�qJ	��PN������Ȕ;���  O@����D�ڡu�
��Tj�2R����΍VK�p��L���O�x�Ӭ6��x�e���X(�4?��aa��?�J�ů;V,y�c�3G�t0�`�+1�F�����5=��(s���	�ʜ��+����f�X!Z1U�d6�h%��gP0a̸�E�1^y�adV�Or�H�&̚l^��H�aT�Ix9��'0�&ªM2��"���2Y�zqV Y�1Ut\��1\V$���Ɠa�yJ��&X<ys%D0\�n4E{'	i���K�(Κ�De��GK�
~���o�=1���1���'ys�,�@��n���c�h��VM��W?m���$�A�Ē�
Ť���F���e���Д��O�PJ5|�.� �`�;OT���K=z�����_,�h�A�m��!��㆛�j9�%�4u�S$7��kȯs��� N6S�l��C��+"�X'�ݗ�"q'��P�]�(e�m8'��: bӈs�Y��8O`��1���~͑sB��C��9��2_\a��֞=*@�t�ٓм�QEԄ�z��BՋF�����0T�F�l6R��e�}ƠA���=�4����{^P��,�66j�1cр��>(���sv͚:�hT��4k�@A �/	B�0`b�ƒX�>��޴n+���A�F�� �2����!���E ���G`X�2��4��=;c>���#
x	�mS��"�����=.1���wP����O�	��i�r�? �DZ�"��)�$�Y+"敳�Í'$vY��Arܓ�*�����r�J5����i6	8�HU�R��s��m�Xi �P�E��a��*��v���8���k�!Вm�X0!����^�5F��4��uY���c����Ô0��$�?�A2��ӌWȆ��EL�}X�7m��N�x���ٰ4�(�Y 
=lgƕ�H��i�^��EQ	���Ff�8/�`���*�"76P`!ՠ>i`̝�2(�,k�T :��E�S���7o
��Ø5[�����-�z4#��2�I��
��E�4�!Hǂ1d�J�Y7_���SD��/�hh@^�B.f��	��I\P�g
�I�"F}��պ�!�9{2�`! ޅC-`b��xq��G?�QV(��q�F����fPe��`��u'�N��� �U6}5�aR�v�^��t��e�#ۧa��u�G�]3֢@���>>�Gk]5zc�%{A�Dݵ{f�+�K�N|b٫ @u��A�g�͑w
^- �KK�L�p�îm@�a� հ���Do��6��F�wXk��ʞN�`�0�O��Cd.�3�%���D�:L`�e�s?y�	'/.���J�e؆j��ś��l�`��.��j����w9DD�#�3<�ұ�CwJ��i�_9�1������T�$�)0�t�S�O��p�@ ��R)B
?1���#C,E{�Yx�a�4�"���ɉV5&�r��Z�ZQ��<9��H��KF�ҟ+��)�JE P.<��,��e(�'�T`b���ʘ�yr�٫I�:|��D���(���P�z�%ƶ@�P��^��
Ӧi��E��P�
X�j�Ox$H6j�%�!C���4x�A�D��e���X��L�C�1*V��� m�X���Lt�e�5�����`c��� ,�����^�<�#a�ʹ@4��[@�۩8�dE���a�la�a��V/��!D��y"�Ɛ�J�q�`��c�h�SW*��A�����"���%5]P!�P-��T�IH�E)t]�IJ�%5�O�A� oY�&���c�F�|I��ە	���K��9?F�I�L��u��ؼ"�����K�H;��49A�.�f��2b�<( =Ss�'���	��Hv*�ȅ���q���� � �y��ͨ"�F�k���xt#@O�VzԬb"�8��a�П���
��@�C q�:�0"oAbj#>QA Bz\X��YC�!���|��Ϙ)H��1FK�Lih����}����t�e�L�$כo�@!���O��y�B�^w��+�e�(_S x�s�O�����_�*+T٢bA[�Bf��O_@��E�5?����#�zM��%`'��ࢋ]�TI �p?!��R��`hb�ʄ@a�H ��
�(Q��sU "ӆB�t�T�x��C
b?.<i���3o*�P�e�Y`��](��8��� Ԝ3"
!�OF)���]��.�A0�Z4L
&T�@D��K ��1-&�m�t�6N4�2�D ?�$�Y�:�s������*�4���ۿ^��h3��<��=����O�o�x�d�ݐ� �RLĢ/v��
q�1�Mҁ�C_�� 4�O<_)��3ړ`RB���	�j�.%S�H��9���O^YZ�Bъ۸����֝[J�!ò�\�>!Jva݆��@��=
�u�%O�e�~B�\:s����B=S�I��hOp��.��)I&��0O���'6k|)�.�c�88��*�ŭ2D�\���N�2Bxl*3���Q� �b���O��1c$G'1T��2�lЯ�~���Nwf�����jdj܂"��$P��C�I�\]`T���6wv�C�,f�a�'w�����F�'��18ϟ�PK@K��!�l�R�ðUhT��w�7�O���uM��()��bF&�%gx�%�A$��W�`�ۯ�x��E�M���^���]��V4��OLQ�
'��OX�	3S)�Y�^��v�@�D���P�'�D����r�\��U�a� � �'�(|��hP�4gB�,��	��I1�'~��#�=\�@%�di���'�C�,�1|ΐl���݋f���'"�XCK��dCd$�K�X\��'hV89����Z)q�9�t�'����G^�S�!s��� |"�j�'?nl#���?=�Ț�$y�H���'� �УF�K����!DؑD{�(Q�'j��8qM�ۚ����i�̙�
�'�R�����}Hd`yL�d�d�	�'ɌU�b��s������^Ȕla�'� �[��٨t���
 %��M�*`��'�KG � `|����ٌ
g���'�
M�%�ޞ-֚M���O� j|(:�'rD�f�5����b�����'�f*6f؍TΘ:�
G5h� p��'PNl�cl��j��)�I٩?��mk�'}�� �a����MR0�XpB�'w��ȕၼ}ގ�t��;*	`���'��\Q�G!o�ԩ�th�m	�'�Z�"� �@iy&��ynR�a�'��LG��ˮ�B�,��e���� ��ԥ# j�q�aK]����"O<`A&���S~�%;�Ƒu����"OLu�c�uE�@�$��&ꈭ"O�����ܱ���)�1�t"O���`�%Dlf�:�d��M��%��"O��0��W4ڡZ�b:�I��"O��Bc�و��D���&�0e�w"O8u
V�=~,�(SG Q0�\4Ip"O��9���_Z)r��T�$�i�"Od�'jA�'�<����!8�N�"O��h�O��R*i C�\�X����7"OxS!k]8W~��c�B'z���"O(����5l8|Hg�*�z�!�"O���!�#DN���r�K�4�x��"O"\y#�Q3I��X$O٭$�<�bC"O�h��ޫ8p��C휭s�x<�u"O<k�.�1P<���įs��p��"O���¢PJ�L���·�(�( �"O�����V3/Ԅ4{g�S'����"Ov�{u�5�;�L�E�mp�"O���-�(-�\X[�-��4�@p�"O���h�;���[��L�B��� �"Odm%$,B~��I�Kԕ~�$�A���
?g��$��'��� �)�\�� �b���>��1��A�Є��	IR����5<C����Ȗ.����dE����-^$ �O���Rl�%D�<|�'g���}"���v,O�I��ܢ��4�l�)�j�5�,��!��F���@�
($�Duqn�+}y���˪�jrϔ6��	cܧ&*�auƒ�	��Y���ūVu�D{�	�)F^�����uQ (J�*��A �)�����`�
!s0�� *K�Y@̵���]��D_�Q]x�:��L>�[1ǔD�R�X����Ԩ^���X�
S �p"Q�r�
�o�<BXG�D��0R^��c'I[�b���4ŏ0:΄��<r���/�\����kp|��Z�A��5J���� ̚f���XK��#��� ���S-jvp�%�>G��5"p����(�$�D~n=�a΄7��H�!�O�|r&��<){��,7ָs'��P�q��������s�ѡ�坵.r�	��`/:�+QQ�'\x8�cw��@IS3��#��=ғO��� �9����'Q��pi��K�`x�I�N�\5�b�7*��-W������͔z"R���-�b=�8�^=�'�6*��J����^�|�����H��IY`�N�>5��h���/���IY����S��O�'�uOׅ7��S%E�V�<`ɗ��Wmducˏ9SY�!a�.C~,��`�V�`ѷ�;��'p�1�&����̴�+�	�
�ig���n�
h8A��z�d��A��[�O����i��-Z#�
'
\!��~'��0�J�0�Ċ)Y�d��MP�s�`)���4ML-;`Ѡ<H%i!�F�b�R�fHH�a�)�� ��~�(v3k��hH�iQ#:Z1���`�P�S�I���l��(��c�9]���$M�G�v�1 NҽQ>�	�p�%��gA�O�R٘T+�%w"U;G��?�A �P�w>�%��3�p=�� �z� g�]��4�Q�Z��I g�t4���H��r)���ߍ���Cv΁�Bg�	3�a�f��H�ܘxć�/~t ��[a����O��Cwʉ�RGF�0�u��ƚ����s��6j�
�䅋\Z�0q��bn7	�B�H��E-�䡊u����?���T� #H�r�
_h�$�
�g�d sW���z!6 �c߰e���Qm�3u�� �B�u8�KF	�d�j��)������xɌU�B���iA�T��� 'E	�z2�\�xI�f$���?A����#9�A��&��9O��PgEG�_��%Y�.�.W��@���"}�uAn�=J��b�H}�j0�7�����.��P�L��"|�a)��J��:�
�2qpq�,\$�(e� ��#@�^s�ֆ3��˓K��R,�[�,gg��K�(ȗ'q��:��/4a���I��6�r�gJ(d���RF^?�`dQp..Rv��:6(ڬ5e��べ�����-��9�GB�1U	���1hG�x��x��t�J�(�r<��6P�-�z��	`�dIc�m��k@+"�X����S>8P�:�ģ �i�Oҥ-�"ɣ #T�F�F8 !͒`�*I��'1D�Z�O��A�o�?�℣<]�q��v;&p:d��O�8a@�-�)#C�@�ъT�
*y��B��r38LZ�+�B@ߥ_b�o�M�~��"�M$/��i�U����?لlW�-��l��M�$^`�3?��$_a���EƎ�~;��Q�?y���u"�Xl���GcѸ{T᳇IK�P!Z�еf��{3���}���Y�bĈXc��Q��B�RF��B�z �I�'aR:H`�O8��p���e�e�p�3����&A��s��=���Zq�8���
k�\j��\��J���G1	�����
&v���p�O�AhDn�\�h�r��5�U)���C�'m 7F�,qX�E���s͸<�����M3Ư��m�T��2a�BR�k �^f��e��T�,V	R$��>r�1�' �`xu�х�ı�O��RP�� �u3K#vѪhS�4P	�Ḣ��6Hm|�:d.��n":C��,H�u��F��B�}���R�mr�>�� Y�p�>�)�B9�٤q�8�1�Y���O���P��OȔ9r��E�t(������(q�4�#cV�q���+��Ѝ҄MϘ-2Afs%� ��4PCg�����EC��R'�p ���u�^Pד6J�+@!\"Qh]�!��5j�A2b_�����-�݌I�&[�%'�勡oJ,R�~uȡ-�7o�yB�~�)� "���^�2��ebYQ��p��5)@@@�Oʆ��
�,F(o{�I�BAĆB�:��կ��h��#��L�xÏ���*�/R�}����4<O:��p�� �� HGKȞ+���׵i*��rdT�|-��T�>��x�Ł�(BR���V�<TF)�CϋY,�J�F��"I�."��a�(D��c+�D�����G�2��i)G�;���Z��/\�v�zS�ޔqvh�CkL+D����eJG�6��Iw�f��@a.�_���	amģN��*�`#�O�2��Ï����^{���'��>W�D�W�À/h����O \�ZbA�})h�����M���G|�I@�_N&<��ōx��I1w���e�E%D�ԉ�m��A��@!q�^�8�r!�)���Y�Q�aI��:����dQ ����J���д'��0�$,P�.Ѩ�ݝqr1��$;3�ܾi=�xh�-Ԉ_jVLؕ	�2��	��Ҡ��K3�3�I��j����*rL���iȡ	a\`��
�		ฉrG�.{���@f%��/y��n��/4T�bҬS=?�F$����)6�9Qw@Ȓ$�0��.b��(Y��S�R!b�4=��и���u�J0˴cR%�T�#i�(g�$bO�2N? �yA�<��Ԭ;:�����O�N�G"�yj����џp(0�߈8�鑴�w~dl���1���Se��3m�0�G�$z�[�
ɸT$,=�&�â��i�G���~B�6R�+����=��P%�1(B�ABs��:��[.�	S��s�T�NXy��e�<qe�� ;�^����ŗ��$fn�[+DmJ3I��[Oƽz1#ʪk�N܈�b�Oa����)9���V��Z*D#=��O�&T�8*bi(E����'g��lEu�$�L�*�ˎ{}di��'V�2	2��F���������fABs��O&X`�'$jht	 hͻ1ky��BE7]paz���6����ƛ� ��T��M}Ш�q�ڍyk���a
��O�:Y�T'�8>�ɠ�ƚ��쭻H�<�۴�M��ft��Pǖ�"��PQDȯ<��O�T	q�/�ybg� }xiA�J��"1Cڐ
{�y��l^�*�x�p�ϽA�ȉ0�%
��m��nK$��#�	ܦ��T�xӤ��b	Ç=�5�'�0�.6��5oL�(r�a��FD�]Wiδwj�P�ִi�0�U�I�m�4���̛mӂ|94�V���󶮓m�°�F͈/Cކ9JD(X��qa�)s��:-�wB�����I�0)��
�Gֈ-jO>��G��FՀY	�`JJ2�؉�$D4L� }��U�7����Ȟ}BRx�D,R�=X}ys�KM:���wD��M�0U��AT6�xa����`�tc0�C
X����R`"�K6��	�+�B(��.b
HixQkP�bXFX�R�ăw����fB�&a:@���JF�nڗs�B�����k��C��
P�JYqwm�L-�n��Bq���B�9RT�A��&D��R���K�$H4RV�x�ڌ���r>v�ڄ�ǣE����)	h.N�H7��l?���KdP(i�!�)`��)���"0�t������2X�ћ�J	b@2H��
�&�Y!yTN	���K��I%5knp����S��{�ឞX��p�FN�d�+u.^�����Im���Iԯ���c'��<?�h��ƌ5N�i�b��/X�i+���}�<�#��U�%(��m�2l��q��Q�}|�ڣ��(@�N_���(%�@	 �����Kp���BU���!X��V:�|1�]�s)@}1O[�Ft5�ӏ֣.y�={W����=h�Ė�lYf!�#�ؖ{�u#�ՐbaJ�����<`��!�ʀ"C�
/Cs�0��ϝ7kjt�"�ͫ4֪��Ī/�^`�,�4l��x�TM�mZ��R��{˼}_�P�ĭ��hH����埮Y���ȤI�^�̓�H��5�è�~���O�)[q�� +�[�(�걬�?Y���ҵ[��\䛅����t���)Zr�G�\(����⍾3*� �@G�,�HͲ�!��s#
0}�������ፎ��O;Z Ա�-O,@�C��	J��� ΋�W,�d(���:���� ��<嶐Ubd(L�K�hY1*��	�.L��gV�5W�A-_PR
D	�v˥E�s�І�ɨ*싅�V�[�}i�Q1���0%-H,>c�)#��s�9#QKۍRԎ��SFa���2.�e"jeӑJ�^p��#怩�q�ܖ&�đ�A�X����+f�'�~�����;+@. ٳe2��="Wϖ�J-Լ��cM�&K���|%�P�VGw2Ұi2ᐱu
0�BΗn~�0W�'�����~"�t��W��bed��*�J�/�=~�r� `MĨWC�q�˓,����.���H�*�6�8�z�O��|P��UN��9���+X^��y���"o�N��Iߘ7�ԥ��%Ȝ��-�f�T�>��x��Ɠr�f��WC��5t��3H�hYf$�.:z8��H���8��`���Fs�h��W�K2f��C8O��		 <���48V��BE��p>I����N�V���� JBωڶ�����1��qI�
�#'-䰘q͊�Kb��)3�����8b�B�Ҥ��T�I3��i��y.ꈀU �/DZE'.I2.@&����.�I!��K1�ĭ$`arj�:tC�YI�a��qT�` D!`D �P���)�����U�WD
F$���Г��'Z����?Ad�`�q��
g�Aٔ��$p�4������f�~��X��@v�l��c��Rߔ��i�	 O�PW��0<�S�h�i�;D�nu%ƒmf`�5�8m��{tkV6Rf&}���F����&q#��|ڦ �_���a���Wo@�(��0d���5&����	�)w� �1b�A@j�k3�]/�±
wO���� T�V>4%��� )��r���\J|H`D䕼VĈ�*�������$�DBP�S%l-�����?�Ɉ{�����/�+�������'�PT0�f
�w����1阽CPu��1n�9��Y+������"�PhXc��~��ߋu����!��6?i�s2Ê/W��`WJۛ�hO~�Q%������R�Էy"ґ@�����"mGl��t���F G@�#�����W�I/B��0H�~��е&��A*�ҟ�@ �םmj�� �{����P��z���R��Hl�����V�d�O�.�I�'�~�$�A��pu��Qt��`mVdC@Pd���S�D�
�Gݒ���`��F*���T�>�����%�2fߓ,��a"��q�N��)�0/j�!�k�#�`�i�Ś��-�����s�
4>y �.b ���*��ي�!�  �D����~2�R��.~d!@�픘�hO��Y��Z�0��OŤ[�}@�d���Q����E%^�Q0d$p�h���ŉ#)�@hnx�4�G�M�z��Vn�dx��⃘�RHbP���i�r#>9�l� uVrk0�I�k�,��уZ��*��9s��R�ǒ+���eJ����S��-)j�OTf� ��9Iz� ��I�z�d䱃
ǲ2��<C�%\�X�@yf�|�ܽY�PQ6��9�v �O�1!T����A��<��� �����܈
�Ä�@w�}R�oY�i�X��`�̫9@�1dG�'"��f�T�	�֐J �E�F|�YB/�ɦE���*CՄ��F��<(v�]�"YB�
4��0)%`8�Q��f��Y:�%T+@ݐ4۲�G � 6�&%UXi�����* =!5�:������[��E��&#�T� � ���X����Q+�O������2��U���ٓ<)��X��">�`Bs�֟ �#��Re�)�#n�"���N
l;@���Oj�E�Vo�Hٴ�x�ˌ3|R��;�n�>�������'~lҦņ_a�����\3Dw�d���ȕ��c��Ƶc��IFbN$c�T�q
��wcph���؛c-� ��h>��f4b��!��ρ#o�H�Q�ʮ}&z�÷#�uz>	JD�� ��I�����(ɖ��+ދZ���l��?�jacYz]d�SA�#���zTNA�O��U�3Qiݎ*�o*D� l��
�9�Q��m  �εjD��M��A�c��k؄7�>8�Լ�G(&b�	�GM�mΊ�ۣx��}��P!O� ��X�>���h��g���$��iƘ�Co	�n�buq�-�/Gx���#G�0����
֗��j��	y6f�Y���o�dy�<Q[����
��)�2�HQ��Ja"�s!�L�Ύ��(�	�F����=�d*�LX�/�(�8�ͅ�Lj0�K1�쟌���W�6�eY�F4r&�s	�<
�j�)Îٗ7�nb��9�.�3�xpK�B�"7���z��
�F�Ze���>�p(p��!K�hp$����n �$�tO
G�Vi� h�;�l(�j��<���F��D���Z�Y�t��U��~���oѢ�zt��-Eu���c��Q$��f,C�f�z4�ϼ>���` �{c
p0� ˕B�F��B��	@�'�@�H4͔.z"0M��(���WƅC�`\0�%Y/y�`X�ᬚ<vhJ0x�#Y���g釧ˢ�[�愃@�j\��Y�}�vl.�yGm��jA%��SwZ2@�2��]��̧O�l�L�Q�1��$�S�����ML�{�8(�@�
Tj�p��I1[����'L�>Y�f�5�M��ˍ�}� =HF �Pm�`�6T��S��L=u��9k4��*��DSB�o���[�$��B!ۿb������ߙm@������[�� `�:D0 #�\F1����1EM�*֬=�]�U`Ւ{ڊ[���q����Po]�HxTgCK%J����Ɲ�Qdw<�t�t��r������KrHQ��
�M�b�P7�	�;�4�ҮB��+P!�&a▴�@؟��FPݥ�$���@����xxShůGN(I�A��p���`�2�L�T�����7ON��.L$+�P������<q�ǳi�a~҃��ri0q�%�2'��C� �d���LX�|YH s"i@>#^�Cπe��E�#��k��ĉe��	��l�^�	S0�!�.gQV���N<�-��A� i$�⵬
�[ڍ�'l� �1�	�
�Bl��	І;���f	Pq���`iE�O�A���@���dG�(*�B0g[�/�(x�a�$���ւ;��8!E�	U,��"��"���h�A%tk��)�XPƀ��q���G���"-�����	�L\J��:$Tb$�0H�/�л���e?�2C�C��iq5�^t.:�!��/;�](�o�V��]G��u���T�X�R!��Iط�����=�&9����VS�I��KZ�~sv���(I�[��[e�68����g�+M�����k;WQ��>�2_%B�Z�J�*�t��m�<Y�?�+و*2�����#��P�h[ީ����d8(x�F�[A��޴��I ,��
��T��(�?�=9��V��F����%:餅��c�U;Jv�M�{�O��ꁊ��P����Ǌ�n'��@��#����$�m	�3��7�p?��H*�! �U/	T@��I[��Ōʪ#�D�s Ъ\��v���ڔnHش��E 0z�07"O�1c�Z�u�t����+ZD��;��'���x� ��]~V��u��{?E��Ur[8-{�gϨ}`����U�Zz!�d�}���rI ��O�-mT˓'E�5)d��>�����Oz����� )�@�ꆶ_������'��=񵢞7y[�}��Ԃr�|�2�a���^9���G<��L�o�`$4(ب)�$�
���a�'s�Œ�@�`�'3p�lp��N-+�
�~�=��aVtCBތFg*�rq��_*(5�ȓ��!���AU� 5I��(�t�ȓ50�]�w!�D��c�J�IU��ȓ-l�q�RӵcpF���+���
��ȓo ��k�m��ȷ�+�VU�ȓF�L��A#�5z��)x���s��,�ʓyp,J0�����{W�;	)�B�I�Ba"�ش��3rYw�ݒ)�B��R��=���R�[Un��V�\��$G{��U���v��É�y�!�d�u�Iq�W72��%�c���!��Ǥ#PĶ��I_uV�H���?�!�A�JP*A�Yw�)ࡈF!�!�)n����u�@�Hb�� �J�w�!��G�r�E��8P�.�3�Z�z�!�dǞu�>�C���np����	�!�䇆I9ve[�ԅ#�ʜ��nõ�!�DV�dc0:�"@ _���c����\r!�Ău����g��?ᜑ!@�R�:!�� �!���ջo�(���'�<5���;�"O��K5f؟h�^%	�fƑm��!�"OX�!�A�{qX�ct�["T�fu+0"O$���ہ0���0�N֚��"O.�u��0��d��p���"O�X�#�G:m5��P�hJ�s*F�b�N�;}`����	�%���3�B���~�䁿i��0��4(��r���$J6�?��E8:7���� z�$]��.QaT볣OF�O���G�M��k�JY#$���d CgS���Hfvt��!lӠOQ>�KV"ȚeEP�#E�j4]Z"�,�d���(O��B�r�
�*�9�ք�S��ij�W��P�韞McҞ|�&c^�"���)U�z�ť^*�M�C��Z%��l�S�=T_�u����z�' ,��QґA� [i.��I/���A��Xh�'Va���CoY�v�f*��:��j���y�O�!r��m>1��c��j��t:t��h� ��Hӟ���I'CF�I�`��$>	2 �9wS8�JVʟM&@�0�ĂQ��{'�C/�?�t"�3{B(�����]2�+Z�&�pĊD�@?�5�a���c�ܴ��J�G�J�c?�l��&  �bt��(	�A!��q�&?�@�`�@��%�"�`� х�9�؍������0���OR�1�N�<V託���}bVAKMѺq�'��]�$yt,	�f����[�|�؝'Ɛd��&X>1d�ةcx������8ibZ�U�@7��2��N�O�M��� uxR���	(_��9��O�_�f=-�J�t�I�_��1��_�d9	��A���i��K2n�F����H�X����v�K~��~b�+�z01��y���a��
:ʼ�Q�S����'u�}%��|R�, +�B��T��*y�P�m���:�'�T�#��֝5#>�1֌ �{�VyY���#p�Έ�w�C�c�
6͘�/���0|B��Ѣe��xP�����q�e�Ħ9R��W~"��=a��ΑA#�l1�b����j|���'�,Z�iq���)�%A$		���@��T��1��d /�J��4I1�; �S<D~� q���9��ܐ$ �<e���H�t�<� ��'2���lѱ#28R /NY�<9&�=Nne�FFF1?�9����S�<��섶���R�n*6��C���W�<	u���n��d&�*/���v�]j�<AT�[�,�z�)1�, ����Ac�<a�N?9�<xb�\.+�i���D�<QЇ�2Z�qb�B�( mjL۴)�i�<1�U�y�NԘ�Eݠvx��7�Aj�<����&f8���c��q��u�h�<���1���.X.{g��Sa[H�<���L� ���@^fњG�@�<��K����6n�Ⴊ��9�!���D�~HP ��m�9�f�Q�!�ضB:Z�hr��ag�1!s�O�v�!��Կ.� �0&��\��3ƣ��OO!��w�� �kE >n��A�ݻ\!�Ę�i��ڔA_�p#Ե�� �	r0!�֛zݘ�R�LB�Q��B��ќR�!���^0��Q[�}���ʁ/*�!�D�Ukl2F��	� ���ϓ)!�DH"OH��H�냀�	cT6!�X�0q���L�-|p�q�b�"D!�͘D�~!AeɊXe��;�!�S�!��	t|2谐�G:j���hv.��'�!�߸.�t0s��;~���(sM�<'�!�͔DФu� B5��xIe,�7P!�W�%�X�`�J�Z��1 CL_7`!�d��X�e�-���k��0K!��)J�>H�a��^$�*�i_�A�!�d���!s5o�h�S����!��6!��z�e�saZ��ǧ?H�!�d�/�,="���C\xS7�Իo�!�DEq��X�&�Q'jL��` �l�!��� S�6x�)bHVH��P��!�� �@
!e �(��ㆵi3���v"O�|{ׁ]  ��!Yp@@9,�s"O�Ѓ6�a�L!�/��_��]�7"O�Y:��7^�&�iP.F'v� HJ�"O�[�C�<:|ِP͎�&�R��"O����P�Ph*7DW�Y��Ir�1D�xq����__:u
`�SI��k�-D���f�*H�VI��S�=�EKj+D� zb$X�m���(����Dt\=I�-+D����݊k4� ��Vx�`m#G�6D�
wc�E��"�eՋv��DB��5D�8� ��gs�3C�*U=P���)D����j�"?�`� p	3+�*�"Vj'D�dA�&ݩ><P[ .U��!�U+%D����E�tG6xR�z���dn0D���1%O"*]�؛���3�)���1D���E � :�(un��d�$��g@.D�Tz� �0R�2��U��LA�+)D�,�q�S��+\�ZL$�hC��X�<�w�P�`��@�c	���k�Z�<��&F ;�`��N~�<=�Qe�K�<���&88
�������#n�R�<qG��4"�"S���Nd���c�<�6K��4)�D�����=�L���Rd�<1$B�&耉��Ԫg.`,B�N�^�<���.�9bKmX�=S!�A�<1�b >J<��"�_p��rD˗}�<1���>P�t倥���8����q�<�͘�D\mHA-	\ptrW�@g�<) ���M��d	��G��` Aa�<�_�(�|���P���\1�%Rt�<�$�_!Q0#�D	�&NzD�	e�<q�^�Pn4�
���^�a��b�<)��ߠ)2��C
��v�8T��G�<1��Ƭ
������1(�^8�r�FF�<�r��/4��T@�.'
.v!����~�<�����i�S�s���aa�|�<y���!l����Lb5�`BLa�<	b��:�h��/
9?��)�d�XR�<��@� |�b$�,�E��d����P�<�qC��9�^��̒)"'���RE�<� X&��i� �j+� HD�^V�<aEE[	�a`��{ضQ�G�WT�<��d�4>�4@�jE7Ҷ�g�
F�<	b��`���t������b(h�<iW�E��D�"�"ӊ�� �d�<�G��l�d�i�N͈M�0Eg�^�<A�d��lZ�D� ��xA��,^�<i5iߎ]������6k"H��D~�<a��
*yN���2]�0%��N�O�<A�K{�\ԉ�͝$��YꑈAw�<�4O�)Lt�ɺu�,y�x���J�t�<��� KMٿX�J��FFk�<��K��4���!ֻ�60���Je�<��V����P��X�|T�'�_�<�G��4���x \� �SU�<��ǂr;�阣���=�]y�%�R�<�����9�1��+N[����bO�<I�A9S������R��`���f�<�R�N, {=3�f���unk�<�tFѦ8�ĳa��F�����~�<�W�n/�̰���/�ll	#�\Q�<Y��"m���f#I_G
|�e�T�<i#��&f��s/��(�0u3�`EO�<� \���⟉d�
�J���P�0I�"O�5���rO2=0U
ݓk���h"Oq���L[����?#��!�&*O ��E#�+���i#B��H���'HC����p	 �ꓳ�v�h�'U��ZW�A`�.Y�b�R�yH���'���b!��,JڑI�d��H�T��'� xcd.� $�Vuh��3t� �'��Q��έ7����*x ]�'W�h� ��� \7A�8>FH
�'�b��CD[줵����fUB
�'ҒXx㣘�;r3 i�3{���'�9��A�5�h�2柵q���h�'t�s��O&G�zm����#S����'o�������)��Pv�M�T8��'+b!�)KC��ҵL�I���'�@�cB�� [�J�zh�Fs�P��'xT�����	��RtIK�0A䘇�n�&<F��:skh��tO�,*[~��#IX�!"�y���fR�5a�ȓI��#�|��q�T��� \V`�ȓ8C<d��R?+ L��Ţf�$]���~y�vd@8�ȁ�	� G�:��ȓG54�uD	0�t03�x���ȓ�Ȑ;͔v>�lPF��9d���X���	�D��_n^�+�bN1
� ����t@�4��FLb��P��8M�bчȓx�� K��΍U ����/�1<��%�ȓ9zL(r��tztm�nB� �̈́ȓvG�E�r!�]f
�3f���"�n���q>�J��Z�p��5[�Ҫ,v"�ȓD�ң :e5<��wj'Q�`���P�"0�
֗:�.h�.̉,�a�ȓ�����N��T�t�  Cڅ ]��ȓ5'�"��?��jd�ê�p��ȓlU�C��_�@p���3��.h��e ��`6.��Q!�;�iÍn: �ȓ\㔼�	y��,q�5&�Z���5�uZA��?����f�0cr����qQrpYW	�*3ڼ�8��˫[��ȓ�^�h�]�z�d����&'_����,_L8�V�
v��I����W����>|T� �����h�O����̆ȓ|�F�{e(F�Y���9���A�\��ȓ.L�=�wJ^�ZБtLR�G�z��Ί4�l��6�w��?4�����fL���j�!\�堊�y	�e�ȓ[/��`�#wBФ8VKˎ*n�0��bޚ\P��;{���;�hǠ��b��=
  �	�0L��C0�%�ȓU�yAo���[w�Y>hʈ�ȓx��!��_v�1�'�"9T��CE�u1� J��P�umK�;�hІ� ���Vd��Ɣ*�jׁm�v`�ȓe�e��H̶R��]�O�T�ȓ��0"&�^�bo�}���R�-�l��%o�YA��{���[f�\�>�ƕ��|��܁_���H��-�0\䝆�&�:���E��=
�kC�
�A�%�ȓ:�������	���Q�􆘄ȓ4�%� FS�r ��_b@�\��-$�4�s`T�Z�b ����`���}�FI��#��r��9�UN�2����{�4���¾!`|x�&�2-��S�? ��bWk�8ע������UqA"OV��瞪;vDYrfˋj�lrc"O�� ���7d���T�)`��"OJ,꓇_�n	T�cGő5EE�Ĩ�"OV]ReW�?޶��RD*>A�@��"O��9����Ë�U�n�� "OF���OUs�d"ƢŤ-�j<{�"Of�㑅]98�����!D� X"O�eҁd�"E�8ɂd�@�Xx@"O�]"E߬c�$�Q䁍���"O�T�B�|��c��;�b�+�"OF�#��J�D������H-D���1"O���J�T!(�cƩ�	P��� "O�%ڑ�דg�y#�?^e� y!"O��S����d��� �NG����"O�qB7����@y�1,F?FP�`"O�QK��#;r����k�4�0h"O�aV�ŭz=fk1��<��W"O^8A���*)sV��s M�+�@�"OHZN��D�&�������6"Ot(V�O�]a�йE��2��@K�"Op��F�+d���� dY�'�����"O&�KC�X�X���ŅnoX�S"O���T���@X*��2���{�'c�Ȫ#�Cp��DꋴCb
���'b��!B�.C'�� �l�GTr,��'^�)�-ėyU�i��\�Ff�c�'Nu�$t3���F=�-��'��2�hB�ct�CP
:9�,`�'��4 �-FT������ni�'������p�	3�����q�'��%Iq�V뼔)�j�O�(�'�T	���>��1A\9�fX:�(2D���0�E�BDݡ�Ғ�b|q&D��p�B׿��9��N��U3Q�"D�S��   �xԡ/e{�k��.��Z��J�Ś�r��9�AO"["T�ŎP�pV��a�JF�AbE�4Z��R���s��	���!^*X���i]��P�̟sj�,8�Gň.�SeQ8��'�
 $tF����5_�G�� ��gl�$�A�.^�H��(%/��s�K4)V��e߀@a4�2B�M�4-�t���+/]�	�=�R�,fҙ��Kij�a��	D2�h�&��䉆���.�@�R�#`ލ�N�ik���"�5B<�h��\��.=*Ӈ�,�����MK����Q�S!6uv���/8�	�0��#��7/"* r2lG�K��/�&����)L�g�0�&�(�vaQ�K:>�ƠsV,��?f���"ov���N�4�C�X>$�߂j.UR0�̉��\�V�/}�  y���П`�N� �LҼyQb���	!ό��G0u^h}WJ�oR�ҡHM�|{�er����%9ҧ�yGT�H_�db���(j�ZH1%E�'�B7͋�N��P�щ-�Ƚ��t�S�TLj�wR6��p�������;���V0�#�χ>���(�9~�x��ψO(u����$�W#� ���AR�N��d�ǐ �0�Q6��s�$QrX#m.}�4H��hH�Pr�o5Vѻ�A1R���P���=i�A+BԘ�zw�����ɺ.��"���3fX+tq���<�D+us��	���p|'?m�&bƽe�0pa#��`�*��'D;�1�= �&��RCM?��`D��;1�	@��4
��9D�(�у��{���r�S�G��9���<��&�N�5��4}���ړK���#@�N1!69�a(�-f�!�D�^��G ��U&$��g���H)qO��#c�
$�0<!��ɻ`eNU�b�ïH�zpyçDK�<�RHJ!5�XPkW*�'?i����Iz�<��B_�l ����>��FZv�<1��3m~=��*�X����p��m�<����|����	Ϛ% p͛a�<aˈ���b���R��݃�-�W�<ძW�T=�-���d*٘$VP�<�"*^�1ȉWc�H�����P�<ٷ��=\ X�k��9� ��2"F�<���\�x �#χc�B]8t�<��ǁn�-�V'Ղ?g�e �`�w�<��\�@��(y�ϑ�k�8�'ŉD�<��C��L���V���Ӄ*�{�<�V�)^�i	��6&=��K���H�<�J�\��)[��F7k�ٚRf�N�<iQR8"�Ћa$�����b� �M�<A1�M�+��1J����4 �D/�P�<�	R�s5� (�'H�<H���IR�<�ML!iF�#
7~mNܻP��[�<힜6�2!�g�SyBp[�)o�<1i٣Q�TtA��"�ORp�<q��O@��IՋ5&k��@�<�D��UZ^��5�d�RQԩ�x�<�$�9����B�=!&6n� �y#�8�|&�v�x9bL��y�(ƚP�o\=�6]��̮�y"�$-{@|�w%�.pY 	h���$�y�
îW�x�tT[���0���y�m�����E^���	`�y�̀k�4p�ʊ�J< Q�wnʯ�y�-Z5e9���a�?5'ʘ�&Ë �y�� ?�8�[b!��,���[��yB�]��>�R`�]��a+�y""SR}pI��i��I����y�틮V��# H���b��A����y"eƣ8�Z����
F !
�A��y�*��:J�Av$?>���ćW��y����!�
La�i@��h�X�b��y�M�070�$���&t�|�2�4�y"�D�J4h0��	_4�ZRc&�y��:l8؝�C�0$gH�́�y2��m��ȗ�W!���Am��y��]�4��4��7�:	jqIJ��y��R+�6ܲ�T�
��۰�V��ybo�i��� ���f�ݡ�φ��y
� �uS��=V������anA{�"O���,��s�P{·nb�����O����Z+i��O�>�Z�#
�u-�m�a���PҒ�+D��i�f��/�� �%%E\�L	�<	�(W�a�}�e�$�0<y�A�p�
@��'L����HA�RfX�X���$N*�$ 3)�(|^���g�фW�l���ڛN�����'��Q��&ΪaP6��t

4(� ��D��o��I۴�+bV<��T**�I͔��� ���^}���+v�!�d��~�Ā�Élk�Q*`�	��F��7i�\�,��6ۤ2�H�)�矌��fE�DB��`��K*?�r�:!'5D��X`'�8٤ع �F�H\�ߎw�Ř��J��x����78��3�Q	k�Jڰ	�dՃr%� G�`%D}�`�W��	ϓ(T�0O���i���<"P��'�Ճ*��ٻ'J^�
�:�spb�{���2㞷9	2Zwi�ϔ�5��O�q��@� t���B�4B���r���i~PP��^
��{��3("5*E"'Μ�Y9ֽ(�'��҂i��F�Ɛ�1,��Z?` ���@�.�<�K��ʼ���#���iУYgB�0F�M,2��	�-���c��X,n�@UG�2	➤�)����L*3��Q.V,[�ύ� �\D��L�/l���f��M{4��
����'%L�r�����[�'\��{Èã|�p���հ%���2��F>0��aOG�+
B2,�waN�i�PC.�.�<���d�!{0Y !��;H�D�M,��F�ԪԲ���Xs�ԡ�ښY%�m��u�X�S:+Q��=#��i��![�[�mkE��2 ��;��n������6W4Y���w�T���/�2t$�Ҡ� m��,��'��A���j
|��$YE>�C0N��B��9ѧ(�;������;�,�	�.��}�D��A[>m����C���H����ˆ�;� h�@�%��顕��,6��yu�N�>��-u�j�7�Ωq6}��?���1>�(�$������6L֫a˶��K�*C̵��	�:h�`�:�K�O���R`D�	����l�+b̾̓Ḓ�@)��l1&ɚ�<]дP���+�8��q��c���+O����nF�Yɐi����6.Х,STxep�C��`�J$S�ۄ%���Y��B�2���*�25-�Yp��7� �:C�'�D<sc�Z �O)�yZw��liN��3C�Ɍ�*g ��[g���h��ѾV��(�"Ɓ�e��L\�d��'J�Y��w��Q��MB0�`:#�"t�e.~���b"�+L� ����Mϧ\RB$! �����v�Y�/]�V~R �!���:��ş�x����5��)�j�/P	j��W{\ K�mݢ���:���X����꒠3E�1�rK��iL*Y끦w�FAT�H4g_d���l0�ܪW�Ԥ����"���x��V����	�%n�@j�,�1��a�ʘ�<�$�O�A�*�88�0(
B�&ˊ��������s�7m�0r�O�Z�b%(��dfDD{q�ʢ5�PʓF��Q���,����� ��':>*��楍�W;X�6��:�:��,hW�4#@�nښ�{qÑ99$��'�}�,��?��63�Ԥ9@��-$��a F��"5��h#퍛�z�b�ۇb��)�)��<�0��b\@��DOE2J�����d\�hV�E�L�P8���8J�t����c_Jܙ�/�L���D��ʼ�s��5�ة�@�St���a(YA?���&b��3dA�b���c�D���3����z\Ƅ6�t�Х[)7ڰ�a�Ƈ%hXXCP�@�U��R�C���j�'�XK� G�68F��$�2~
ݹb���.�����&ےO�(%�<����K�>���.�Xѻ¨؊d�����0_	��B%��D�FD<R"�`	�)�%�@ D��� X4h�$�^ܧ-Jn|��,�o�0CW�?&��ҒDFZ�6�֮�q�Z��*ɢ+FvL�U�Þj�(kgϴ?睁h_������	�~�^���N�O����Y�z�BK�"~�fM��0���0c��N;"���$\8<�`S�K�4� ]ؤ�9Bҡ��'0�����K14ݨsD�z?�)U6!)�H��ھ/�"��ePR�$ѵ|]fAJ�}Zw^nUb�+� W8��.W-{Z$a�n]�v��i��G��l-�BDS��U9�J_*\jd���VB�'�İ��ǹ9/�P%J���{�Ȩ �� Vf��h�̴�f�2~��j!bfoB�HuK�T�V����A.ti¤
'�AQ��a)%�O��q�O܁����j�w#�j�B�C��=�H�+�`�炁-!#�7-:'KR%��u�D��$e���wʘ�{�k$�5p�*(�0�T��Py��H!�*̋�R8A&�+��A/QԐ�i�hC<9�,���=0�r�m�"�8�ۣ�S<H2�{A� ��?q�A�39��V�N>u���S$��P��|�5矸k��JuM�	���% �>�ݪ6�Q$���ӣ���Z�ы�Hѯi�-biX�9~$��@�}�'6ntkd(�e3l����7��\h�y��A�4��p �C��C���iF×RT1c�͇C=t@o�.�ĕ ֣m�i��7�`��H���d9��	����qc�"P -���mP�:Q*=;R�P�� DPl`��)���Ӂ��![	H��l^��Edx�� ��zy�c���<�B�	�8�.�!Ō�|�~�;���Zv ��COS�T�6Q�7	������A8� �qu,җz�j���
_}Ȑ�4��`�3Cڷ5T}C6�M�X>:�+PK�:1�uS� U�dR����ヾ�������bF^��1���4������=��P�P- n��@#PK��0�C��'	ٚ4�֊�6��ᐈ�$ǐ'�vPIW^(_62(q���h!tq�jGtw�./��k��¶3�9�Cʻ8�P��q��9�4T[�R����P�ڥ-���JZ � DH�
�A���=ғ�~�`uKs�
��D�@U�D\�e��=+�&ڽH��8Z�jU�I9��@���26d����ɠB�JYo;�f;̵֦y�HQ��ըh��v��I ���Lqi`yH>��,�sone"�
��j����d L�H�J�(���& ����>J��!�%ϐC��I0&g�z�����c[�4Y��e}H��	�K����OA��YVg��6� 쬐b���> ��d���LcD��-޸�����K��H��7A����"�
?$��4H � H{t�N�(�Ⴅٻ/@^��pf	�?�`��iQ.^���r$�c���#�*���%8ʓ\h@Hd!�0
&X%�s�ӧ\��+�'�BB ːB�9x$I��j�;#wfXh�AE2/D��g�O�;gF�Erm9�틐d,�;�'J�z�ʹ�%�P޴�a�"ʓe$�{eg��|�ҕ镏�V�f=C���UF,��&�r
�@.V0s��2e � Mhny8'@a�8;���QX��Vp�Q�.�1p>�2%�7���`2%C;#���C�x�
uN�1��&��QO�h�0��D�H ��3:j�iXUdK�a�ޔZQ�Z&��1h�^�1 �4S*Tt�#�D�1 ���+�4Ɏ�a5B�>�N擾>� ���v�^%+ŕ,A�l�X��A8n�M�1t^F�z�nG� f�p���s�P1���D�z�bfA1z���
9�lAyp��8�"��@�%Y�J����W��t���/S�Q��J�'�z�(Ѥ�!C���
��1G���ff͋H4
�κd�.�3!B��h��:햅�0�l�PQ#�f�	#�����b����Ħ����YX������}�ч�6Bt�6D�*���r+�9	��� @F�*E2`�r�X�,�𼳀�
b�B�*�����
���p���2,I&@��]%:ې}��^�zL�,y $G<�����ar Ɍ}*v���'��J���ЯH� �İW�ֺN~��02)ߧ/�l�@@Ê#v�~�0�	Φ����	l��/}V��ē�JW~�ء�&�I�	\<#�ޝt��|;DΚ�ڐ�D7���)��5@��)�A!
T( ��_q��T�>it\�)��i�	Bg�a	hI U�Ӆn'I�f�$}REp&��T�0Q��$)Α�`%��k|�u�ؐ6�S�b�	Vvu����[Q�(�0/̅� �W�hl��Ex�b��8�(�ː�
i�TJG* �:f(!��'E.�E �9� 1h�#_P`LabÅ!,�$�2% 8�� {�e�&0R���,R���c8Ox\qrE`?	��͝@U���B
m|�$XPn4Z\�1�O�n�v��=���7{�PI��g@�w����Y�n{�x����?s� �X3h߸1�/�����+��ԯ�Mc6�x2�H�Q�*���6lO8��=�PBĹtN�Qh�G*��Q��''@�{�$�%}ش�iZ-T}�@���1)�6�n\�eU��4$�L�!ck��)�P�c�G `%*ES�NT�0��m�"H�0�xF�'��\�R��/h���пC�<�"�O|y`3 �f��5�g��F^�]���M��l>C�:�2�5+��;��P�AkcΪR�4`a(��������$\�#���O���r�H��$vU�ƏO�����o\��pA�4
���9DC[����ѯ#M.���-_A1��;|v��8��G�W��!ٲ��8`@���I�9bF��W���)>��d�ʹ0�Q���B"c�����A��G��\aC���$<
��+8��[O41�]-v�Ih�Fx�B��*j���c���=��"=�EG5A&�Q��j�7G�ą�PeFYu6H#\��tZ��[ I�z!����k��-�`#�%�(�Xn�I��-� "�T��$�-/~�!S�f���R,�T���M4����G_3fixа+D�J�ع�#O�-}�)s���
�F��,�O1���BG�&p&p�c�01�`D���٣�0AJ�� 59$��ϵ oˢ����r����hSR��0.Z����.&�p4h�N4#h0�R���������U)L�����6;�d!�k]�9�a|�g^���aU�#+Ya�I^�kŖ�5�M��N���Bѕ&��7�Xg�T������Q�@�rDR�+ݘ)��zL�0�K�O����\��(x���8:���2቗5Rj�;��,��`HԿtx:T	��v����CD���P�#��͉'� �ɲ�T;M��M�>GtƬ(2��*7\����@Y�'g��ё�:qAH���U�|��=RT&Ț�4�{�$E�7�H���k��Cl����l��rI\�zk��y��*�I��z��bP)9��	YPoI�h�l�rƨ..��S�'�г�⋰V���h�H��qaʾ-!�<K�AD�.x��6��;���ڴf% �c�t����U��y犏�߸�!�K"d���U�[��0>1���6��9g�<!C�l����&F½(u-Yet�� B$Ȗ+�]cB�UފI(�'�$I�D�iP7#Lҡ E��a~��H�X}��Q���+l��ȕ�$T�(Fx���F���c䂢]ʠ11KR�M�HaT+O;9Ֆ��jܮ ��qcˎB�����2���Z��ʒ?��h�@�<݂%�������QW�ʱ'���X6N�deB��M�qo�4+��f���&���y'�K3"��� ��>X�X��YBiY<.TY�D��"v���*<�O�ё��3(+�9���n����o-c��r#�x���i������FI�-)�1���>j����?�� �sKL&*!4�C�KM�b�S��'@0��u��4����b�R�o:z p�gY"�ұJD�[�/�6љ�F&z�b���*F��]�2O�l=t 8'ؠ�ܥr�X��9�i��b��;��Kk^Uz��Ӹ'�(5�S&̨NN�[e��V�x[pʓ18lи��A�Kv�<�d��G\�jQܖ9W����!5@>��ޫb�a�c�ɪN|>E9���b��h#d��BA���!��R>�LI&͏4GH�b�ČX.}I%��d��XS�D�FK�����V8�9s�	��G1�K�ŪW5���w�Y3ƨObPaT�^:&_Z�buC�<���K4v�d1�3/����0���Tתl��W0>����j�3K�J��qm�6s�t)�OP��(�D��ؼ�b�4p���έ~���ClNOy�o�:��a�R�L�;>�D�Do�?j��9�*"N&\�"oEiB��`-� �b�ℂ$/�$$f���Qr��'E<hʒ/�@`K�����ƴބM#�I�K�֍QV�_BMb@+�'P�H��n����)�mŶ9������*L� �� :�I�r��q�%�
�RCJYq�o�#1��x�K�^��S�$�,-:�A�v��O�t0RB�,T_�mؐǕ#H$�0�?�t1Ue[	qR-����7�:�;�	��|�����O6�c̓��lP�e�w��2���5D��15�<r��[ ��8��X�{����h�yR�+M셻��_9�z����
�i@�Ck a7��1gݸ~��hӆ��6��5X�c�qҕ�7��mH�,H�k��c6�-���;{����`.K�hW������7��)�Uȱ>�B. ���)t.ȮF�r| �ET5)bp�j2oI����Ã8.f�#�.s`)q�	�4��eC���;�"� �ᗒF���_ݨ- �q�z��pK�Iž���-�#���d�gA����tT�"�nH4A2�BFD��*t�XkGAū�0!�OI�3��%B� ���#`� ��:��4e-�#��D"'�<�	�T҄QF�?d�Z :b�Ͱ%���zu-Xu̓$���:�-����țG��+���^���}�1�
�}�v���"���	�̞���ȋ�I}* �� {P �Ɇ�\�y9�3w~г�86!|L��.Q�V��)S��T��y�g�?N�K#B��Y� }Q��σ zT��j�=(��x��B�be�(���F�ÒO6�4Ha�f�%uH�y��>-��d�M``�h॒ mN) SϚ;KFj1�M_L}bx��}b��؊i�h$����#�����' ����O����W��M�~���U�0kX)��#˾|������F�>�L�Ysԑ>����R�L�z��Sj�3lT=ᰃ��qs�O��D��B�0޶8�b�i�X�Q�T�n+��H3͊v!�y�O�B�a&[��N�˶B� ��FˉÍs7o�	"�`�&AX%3�f���[�r���pbaʴh�M�M6�	��.WI�~^�@7�W7a�ؼ��̀=��E���� v�|y;f�L9!�8����|[�x7��b���K�b�>��y��Ձ ����2v�>�cB��H5X��޿>��$�>���O�?��i�D�	x>bu  �Kjn�J�CDo����BU�x��t���@?N鶉��Y+T��JIohȮ;J�E2��W> �'vJ���Ē�� �m��GYO(I�G�"����.Ƀ��©TO�й殈c��H\��0�R`�#	�<3G�ף6���QQ�ê&<��`2pQr1r��ۼ�����M�&i�D�:_�L�SU|.��	�!ʈ�Gt=����O�ĜP55�Ƥ����xp I#��0�&��*zQ)��G6�Bs���;z����kF$ jF7Q(ԩ1����V���Z�`��ܐ�HО~Γ�-s��jD"���W�X}���S�^����B�ڏnx����'BLY�!�.;
����1��(��&�W�.��c�;*L�%���#�*N�	Ӌ�2��' ����6"E���D�-�plD~�''uѼ�L�%C��<$���J-�����a®^c��ȓR�ab���V���D�5�0`�'�^�J�k���̦OQ>I[�BE�G欸�)՟v4]�''D�ܓ1�߮kW������{�R؂wM"�=P+hɳ6�'�L�Z��J�f�ʭ�D�O�sb"l��'�h�u)�N�|T#4�
,�j��'�>	v���@��Q��Z"~����'t1�WaWBR~�D�L}���)
�'U�HPN��@���0��D3k�j�R�'<��Z�Ӝ.H��@��Qe�i��'˂�H���h��58�a�Ar� �'V*�!
,v/����&	%0Sha�'�RyX�!
�$��`�G���*���:�'�X(��.�K�]�6i%+l�P 
�'J�|d(z����%.S
1�	�'W: K�f(H"���=:�K	�'���j�D4*x��j �-)Ґ��'�J�ɐ��g��0c��# ���[�'��i�ш�<Q��S�zd�{�'SZ�	V���BN�` �6P��'� �D-[�J
n���
Kw�%�
�'�l�0�u�l kR$�9vT�	�'i�P�aMԍN0/��aP<�	�'�T��Aރ�B$rI�*$�(z	�'ΐ�S�2>���"+ޡ+�Ƥ�'��۳� �C�rU@3�޽
��@��'H��8`��+@��4�C�� }ʭ��'"���#�ծp��lS@�jg�-Q
�'i|�ꦃ��
�� W�=��	�d���0c��[Qΰ� D�;
|l�1Y�:�L �=����P'قb��!��U����<W4�C-�4ys l�0���Ik��{�a��M�6ON dTy#I-��Xڣ�ڎ]�X,S��	9��aB��%�Mӡ�Yc���'��9M����
w�p�2c�%<��
̤W@��x�(W�3���'�����U�V"L����F?Ȩl81��1K\b5�$}b�i��ܤ��N6Q@��"�iA1wd���xRȓB���O2LlGI��[/rD�ƨ
Z"�s�O��r��铌m� ��5�	-��<�7`΄u��6-X��(O�?�x�̚� �@�l��o���j &�'ͮ]HA/ K�$V>pScQ�S����	61р�bi[�74!3�+���y-X� �������M��z�� +=L�0�j6j�*|q���<�ӄ��#�d�b?����;Mv�dy$���HEH�#}Q|��t�G#�m��BUc����ڵ�0Mƚe�h����fx�@�=?��?��� ���z�FR�XAܡ��l�6"&4�)��<�ݴt1�i��f�D�Y��O$d�����ЬB��I1*��yK���ʴq����RKڼZFa_�0va�>�'�
8fAm��!���k�π L� A�T#)h��8��ͨ=
� ���OM�'��O��[��)O:��Q�Y�I0=�Ai�L�"�j��O0H�I<E�� "�0��dB��ġ�N��y,�Q�$ݐ�a��a��d���v��)5�z�e��%c�Ox�
�4^��c�b>]2D��!�H��3�Q�1�i,?	Gv�Dp�y�����	�,��rd�� x�Z
Y[���,���>T ͈�-;��� ϯ�N�����y
�'Y+n4�a�T%�U��#ۛ�����S?!�z��h��?�8�AC�T��ͭ?�C>J0vDoX#|�
-�Sf��!�DD��6 BD&D0k�\	�*M1/�!򤝺w*DcB�e����*]�`S!�$��_�L����o�0]1���(D!�5<�:� 7 �U.f���/z�!�dƨz�:�B��'�E�b��w�!�D�;��I��"��\WJ� ��@+K�!��-S*;�NX.[��b��[�j�!��ϡ
�<-a�ϐ<|�8IF��'�!�d��E��P��Q���H8�)��R�!��)
����aVظ��� ��!�$��:�4P�O���z��] B�!���,s�`お��8�DǐS�!��l��Hr����{3�=!��qM�)0�L�Bl���eP!���)|�"��#��^-��b@�!���H�2dрc]o'(�x��،�!�䄘W��hڈT����蚊f�!�D�\�Ps�(�h��2(�\�!�D�Qv�(U�������ڍW�!�I"� �����W�<�)��C�!����D�􆅽�zQJ��15�!�d<��M�f�nhə�kY�*'!򤄂:��y�%�#e�M��k]�o+!�$� �H�C�i@99Sfy3�
V�!�D�O�.�2�蓬>�<��Qb	!���Lq��b�;j� �ҩ��;!� � �TH�0]���&(��#�!���̆e	rk��F�~�hBFQ#�!�d�(r#8�3�D�Z��x�d��!�����E;�`�����!�H�A�֒%��d�á�L�!�K;�Ι��OǴR��l��N�!�@�j�
�j���=���(��D'V�!�ׅ_z$+��
,�t�C+��'�!�Z�����S+�hHҹB�鏨)�!�$ߢ$v��y�-1lH�6nĔ9�!�d_�rc*:&
r1�
�`�!򤇽*����
/%�1�`��!�$�, L�	�DNE�7:�ˇ��K�!��j�Hʔ)ƕ^c�����̬&H��3�\�	��T<Utqw�Ĥ!� �ȓC�쁪�ކkx����&���*,�ȓz�*�jF(A$x j�F�l ��LH4��6懯ǘ)JQD�>�X�ȓKl��'ټ�%�Y�|��}2�,*D����Kď�v�r���)k���HSg3D��Y�i,#��5�ֆ�	�T�K#G.D�D�+\$T ��`��aP4u1�b>D���j7 �a֊Ȕ��=�"�:D�$�ҏNR�����,=|r1xt
8D�����o�b)2��G	]�F}BwB7D��YЮϕ#u���Ç�P���"7D�4y,��f �y�*�he�H�� D�(����.>���3|�PKE�?D���GJ�2,���{�����K;D�� $�v�Ҧ3��;f#�`0��R"OdXb�]>/s�]ڢG�C�y�"O�q�`�׻|�<�H h�M��С"O��`BȈ�;�<;�h�hoBP2`"O��!W�C,9L�`�0(Mvn�U"�"O����4�1cf��(=PF���"O����뉘) b����;$.�j�"OF���0H���Ǯ��B��6"O���p-�kh��b+�2c��`�"O�xBƏ��j2xx96�O	\uBw"O,�H"e	�ՓA
��l����"O�Tj�*¾.��eN�i�,xҒ"O��K�$V mvP}[VC�-�t�!1"Oz��˙#Gj�w(�~r�	jS"OD����8̍�¥B U���*6"O������ �Q7�ݏ$���"O���������h�#��N�^� "O ���ǟX�iЁ��`�R�0�"O��kȠ<ZYY�@��q>=��"Or��.�2n���9v��4\����"Of���(�u�Ob��0"O��t�]�;��8R��Ї{�  H�"O�0���@�D�>T� o\�y�X]�f"O���B�!���b��0>�D��t"Or�x�HJO�x�cC�:;5Dr�"O�s�W5!*!�'�G&��2"O!c�"�"����aU�+�9!"O�A���I�Ԁ+RK��o���"O��b䈲KԂt('
�"%m���"Od�S�K01�� ��K��2�T�E"OƸX�*&o�0�0T V6h��y��"O���ܴ"Ū��z�jH{�"O"Y;N�+ ��j����p��h�W"Oj\����v����$�|xu"O�p
��_~4�#���ցK"O>U!bgB�\r�W7a�X��"O�@���bA��٬��|��"O�q��D:yG<�{�-�.x�8<15"Or��a�&j��9�B�ƽjٮ-�&"OHPj$��%���4=ɠ0jc"OH�����$�L�$[����w"O���P�G�!gF�J��'t�J���"O���W�<�����ܭIݒ}i�"O� �I�#R0���A�z���"�"O 	e�V�B2���'^?s�XE��"O��#��	�a��X���G !X���"O i!��p{L8�T�O"Ey2"Ond�6$Y�O
�@z��L>0���"Oތb�F�#h�8�0�%(j�;"O������*b��Eʕ[[`�Y�"OJM�`��.V}��{��P��$�pc"ON�!��\v���P�KT�S 1��"O�C �P���B��#JD��"O�H�s@G�%���zv�J"C�s�"Ohp��ʫKrX��čO\� jB"Or��#mF�7{�I3�E֍f~�cF"O����MLZ).��S�̩[cP�"O�����;J��僖*}Q��"O̠����K��A`+>h���y"�.uT|��G�5]-�+2@��ybNA�s��%�BD|B(�� ��y�kH7�5;Ug�7�4�P��
��y�m�uqf��rc��y����Ê�yRcT:,DQ��	y�V�H�ˁ��y
� ��SWFϫj� ��h��zbPA�"O4�����]:ڑ9wL
CF>��2"O�\#�%��.��&*o%�AP"Od������ZEb#�Y����"Op��`^�)���B���%��"O� �7�2.K`ődϻs��m[�"OJ��r���F�_-
����0"O�P	�Ԓt� ]В��f��"O��J�(z%� �C�=C����'"O�|{��
)q�Y�%�T�?��!CP"O�*R�H3g���C��7z:`�t"O���� ���#Q�˅%L\�""O�ؑ7k�a`�� F��:%X��"O�ay櫎?h���T�9��J"O�	�5k�z1(DzBh��%��"O�T�ԋ�
�T983��=|�H!"O���a���n�|02�NB
F���f"OVm���#~��07��#z$z�bc"O���� '�~)�P�P9P�����"O`([��ڋC�Z��� ��P_��`"O�4qC&C�$�V��4�C�Hfr��"O\)4��1 ��\�Ə0K5"ؑ"O��GF܁aɄ}h�M ~�M�5"O�juJ�'�\�!#��6h�"O��a倉�;��$�K�Kx F"O�Q�e��Mb��� E^�K�"OV����"F%�Q�Q��~ Xl��"O�|�d-6k���P��$@��1"OJ����#:��D�)
6��kb"O����b��oH�P"���1'��M "O�Q�CB��и4a͟F��j"O��V���i�fy�.�2�~�"O8(h�$�`�@�
6��3p��5"OL,���U�v��J�M�ef�|�U"O"�p�cֶ{	�H˗J}�@9H�"Oj,���:����oɹ;�F!R"O�*si?5q4	6'�9�Y�"O�=�afE�J��(1'��.H �"O�����f���cLES��*�"O.���Aa�J�EKH1�&`�w"O`���$�I��آ�W`��٠"O��P%Ĭg�H���Y��D=0�"Oh�0���e�FH�QW<��UD"OX8��C�`=��s&�B���"O���߮x� �G#J}���23"Ojm[g�I�R	�2��|fd��"O
 ��%!irP�ǌ^�~N��"OX$)6΋��
� f�3~	��r"OT`�f#;%��DE�=���q�"O 
2�[6q�.\8��"l�d�B�"O�lAD#gs�ŚSᚽ}�"M`р+D� !�E�����Iچ(��P��A>D��1��C$4F`�WI˓~��0� C=D�t�BI>^xT� ce�R�`xq�m6D�4jN�1��� (�s�T(� D����ю8����M�������++D��0@�PN-аH��O����(=D��{g���4�r"˂04����-9D�\2p��!3n����%�|ܺ�&;D���	�mQBTZsi?.-tDQm9D��ׯP���2��GTp0��f8D��8R��#9������]22 e0�8D�t��b�7=��ʠ�Z�zO����5D�|ZI	Yy���AX1%ly'h3D�� R����H����ҫƽ	�$��"O��B��-��Q!&G�f���S"OB|+d�����=�1�`��T:�"O$<J��п&7��kPL)t�P�R"Ol�I���%��p2���= Uc�"Ob�qT��(A���#O�:+Xy�"O<�9P,�vmX(˶��,v��"O<x3#�B�����-A���E"O¨�&�{k���:5��ɓ�"OR�h6�	zQ>��i�:���2"O��{S^�fV�3���2��A�g"O�`��`�&Mx�2� �RzPh�"O$�`�G�$F�J���OI��\js"O���   �>�M�"O���   ��4��y�>}5nӥ>Rl:���,2d!�ȓju�՘��U��� J� �>�^чȓ:�:�y��P4�fX{� ��q�ȓ+�eze�E:C���*�K��E�ȓ?�6����M�|h�E��Q�<���KU�E�� �h,��M&Ԟh��_`�Xy�É5=�����%��ȓ\A� �P��z��	rg�<1-�Y��(����I'U���g`W7G t��=,$��R�@�|%.�it��,K�F}��
s� CBN�=A����%�-u���ȓS����Ҧ �.	3��ê9V��=��!Շ�~�2��	��(����^&�((����T�!��S� %�!�ʯ��˵83�8QpaҲ#�����Ol�xX�+q��@J��Zj�#tO����#R^���9�!xĀ�x@ W�,9(��hO1�و�@|M��	�s��UH�D7u��u��I'M�Ʊ+'�U���!��M����{���U;ܼaB��̖��`@6D�\k�ȥ80	�Ȁ�|F��R��<��"�eXE�K�"�ԡ Bi.ҧd���B�A�5�e����#��Ą�S�? ���FΈ="Kf5[Vϝ�b=Nu�@���o���䖳e����T%	.�'f�qO�x	v�/]��A�6��y�h��'Ѯœ�N^�(�@ ��X���H��ĉ:�3eLF=��e�A�BT�����Q�f��$�%V?����2�W�L0$�'�6�g���&�PB���+s��h�я��z�,0�%W?*@��R�V���ʂ%J|	F"O�\���;3g�"��4�6�	���z'F̸A��SG���I�p�ۨwd�u&�k�w���h�C�X	n%wJN$bbЍȶn��g�4Ѐ�{�����1�H-��'ױ~���T��--�S��U xsn�G�M}���rl��3�D1ڗ痰z��8yOm��g��@���;RD|I��5+k� ���pN>��?n�(b��عQBvQ bĘ>0�J��`
��$18E�$3�����:t��#�h�P�E�?)0J�!
Ll|iG�u�R	�E�
%�b�cs� ::�py䑟���FHD}`X�bȂ�cf�l�Z/g��Q�F*�6�fK�|^Z�y��_<Gr@��%�9g���"���0W��Â���>1�,�e� %���_&W��:��P�jV�0?��YU�@*3�f�q�ԭ��	S�TF���;��<i� X-������0���M�݀B��-}]�D@�bi��`0��Y�f�矬i�bj��U�n�jT	�&�%�L��6(��$����@4dnd�Q�o��a`@�hB-Ys��&�X�ə��!{P�;�H�!!c n�R�yP�ܳ,��k��՚6t�'����ıPdX�XPe[�ldSg�O�`�13��O:N+u����4SF�۲1�����~�I����3d�M�;L"]Kp�[�
� Kf��-u�*���1����2wU��3���x����ݗ<���(ոT�l��_+:����Cd��C�B�!��Q���gU�p	4�
�20.��42�T�C�+��h�w&f��iыr@�M9�w��&
�9]N�`3Gu�F1��n��������3zT�!�Ε��������\* 4>��1�J�V��,�C��
lG\��$,�,U��KJ�#96���+y������ s�X���ކ��'RʁZE��1"�"�^�%�&59��ϢpK��I��(g��Ahrn���J��[�=<�Zv�_�#�"99��O!vH��I�Z�m�t9K�I�P���Jve���FF%��녪82�I�H�d��@/��耂&�j<�IYU�C�3R0Q�HP�d_��iJ��Q�4cE�4��V�c��@QU���3S$a���>Q5GJ)|f�Y�捝	<��m��n�:sE�<���6.:����͗n��Q���Ne�b#��򩎾a���2C�S�~5hDT�uB��sV�L?$4�A��!L@mHW�<e���#c��z9@bD�pO��֭S�0%��@��>��Uag�� i�|�z��S3̼�*�uW|���6�ӕwRt�ƍ-Q��A�eDUj��H�4?)�-�p�$XC�ui��D�dm�3b؁˲iµ�[�Rg�YD�>٤��E����N_�����O�""RU� 䝝2
�镋��Kl��bB�	C��1�N�[������%/@q���'9̬� 	*B[�� m
AZQ#����bą�lRO6a�(K�ܮ��M!I)l�9�K�?5�nIB���*�vMѶ�R�R�C��i�L��%Y,,���;��{d���D�6jY���M�6�x��g��*�"�c���(��r�\6���,��B��61�H���vhN�i��4
Hw<  n�	�T��`��=�� Y�� ���l��HDy�	��JI� r4�'	�P���`ڃ�y'^V��h3�]i�@��&T�0�Ah�{
�F�O��.=
�|��%lA"!��U	�,͘1����Z�,	�b��]�.��q�ز p�إ,@�$.�$ʍ{�P(-l�(A���;ꄝ�f`����O��b����.��i0�0�l�*�l��`	�*����#���]�f-��*V�K���"*��<P��ɓ*|d�h$Gb=��K�@�]��ɣ<��Q�^j�Ū���8�d r!#o���m�2Y�)��g$�5;�h�GmF���V�"C�	�~P�r��t�6X��E9;@��@G�,B��P8��B'�Z��3�Q�y\�R��u�<DHR��;>I睾)����!��0|�cT\������.R��i�ć֟7���?Ƞ ��	���d�I�/�Ѧ]���3,A��c.:e�{�"�t�q%�Ԙ���>̺E��<Hm6)P�2��*z��՝cи|Rt
�%5�����G����8��P�N1D((	<g�D '��Gр�#U�'���[�� tX���ƆD,D ��X lOIY
�*#�h��ZT@�� ��H�T�Q*1���f�E�A
�`�,N�OV�J��ɮijB�z����mM�$kM�!R	�g�J.ǐxRiE� �@��$(���+6胥�X�	���0
��p.Y��	+�L&д�g��bu.]��2G:��;P/����Ù�^Z��. (*��'�xpy%�����c(�d*z�`���W�� �A�L��J� >H�`�_�t�"�����f�!��E��y��ӫ]�"��6D��^r�8O�Qk��G�G������0�j1���5'Y||h�/\!?�Z� s��/��YK�EGC��1�#(��3�|��k^6#P�lS��֐�����."#��{�	�&�|%��	I�I�,�b�|�'n�*�$[��j˥*�L�K��Z<t�|�g�Q�M��D�¯T�b����q�O�~
͋��
�,�H�S޴~1�ع����u�DБK�x�3��]9F,��[�w�'��}���H�v��*��E+��{���6mM�i[EB��;�\��&��<-.�!�3��U"��s��o�L���"�9��U+�8�^��)�=.)�=�c߷W'�����&�H��RhR�A���A�'=�yY�9*�6�Zt�[��+����"�X���/@�����8S:H!%`�7* �Ԭ�=�L���"P��)c"1H�������X�B5:e N�6.	�T�<��'N� �(���=Jl�񯂯`�XX�.�5f��Ė�6�zViĦM�� �#��?@z��aoC�f�D��=p.\��ֿz7��S�Ô(�й�C��)�f��ؼ�8�<A�/C�,�ĕ-2g�bh�m���r�K۪w��:�*`��yɦ
O�!���*��qh�
�8O��
bKڨp���"�F+c�Xpq�$HŚ�+v`��\�2���P�U+��"�Nd��!c�c�+I1)"�(+R��/ 2�B%r֩���D�.X��oۃ2ś֌�@;���eK���7m��t���C>��' 
F��h��W���g� ^$�P޴P�0P
�:8��X�D���8���� �0����OH�d���U�d[dv��q�K6yÐ-˷D� x�ሯ�I�$�ѾhS�O��J�W�p��ܫ�h�{n(T#�j�ZW�H��H��ᧇ�u�L�$�"J�f���)"�H`�� BD��&J�$���C"(O�S\�������,b��Q��'��\�˒�(UҴ�Gj�0�68�3d�� �T*��9y�451ӯ9C��H���'f����
Ӓ3�>$�D΋��P�z� �!f�Z6q�0Xi���|t�n:�p���:J�1eC[4(L0���3�X�:P�5D� ,s�'>��!�T/ �"Q;t+@�9��C�]=����h�~-06d� K ,h��3���h� F�)8F��c @��z���-�Of����:{�)�*N��P��F�-0V��� ��h��Mn�	4��2w3�a��U��."p�ΞCQ��ݖr�J!	Al�#���$�;�k��h ��ړ/FJ��T�qԐY�hNS��-�"��zcFEk��o��@Heڒ,G@��g�Դu܄u�F�ipr�p�dͯ>� �yc-��m9*h���tI����2��S+�;H`|Q�b Q82/�a���ɶ$��4账֗+�KÂ�˒xc"�
Loly��'#�i�l��hb#K�Nj!Ka.}2��sգ����>����2�>����J:R5f	�w`�Ml�I�Y &`�J]�vm��0��ؕ ��M�x �J��jw$�_خ<�4��!�ao�*^�6��ɦS��H�'�z1����$�@!�rI͡x�j�K��ף~��!�I��+������580j�G��q¾�����G��T�C@�!vT�
l�;=�
�X�I59��DA"{*���B�T���Ŀ��y����<��M�
�*ӎ�#s:ٻ��ޔU����_Vl�%P ύM�Te�L?8d��[����� �%Q�����&�p=���.�(�Ʌ
�
�.dJ��4.}��J@ʓY�� �OB�5*B@ےGޯ�&��J�
�&pb��.y��b���tq�@r6 �q�1@m�$��x�ˋ%~���m�lܜI�!	ධP��I߸��&͈�0��@��
'p���m�iׄ4����㴴@"�O�|>X�:�)U>�J4 `\;8�aybL��6yP�@P���s{���'�e,�9�ۏD�R(���1�Q��$5��P�m� �$�1/�f)�1	҃[G�Bb�Zf⌞Ql�8eE�)����0}b`
�$^��w�� F�T���j/ ��X1��>|�f=r�śE6,�q��R"DG�H�備8e��Ab4c��D�>�D��^+��[ϓ)�����>}b�;T\;`��!�B`ϓx��ػ�AW�G ʵ+6���-�0�w��<yl�{�"}yۥ.�v��3���3D�[D쟠B#���	T~���#�M�+TP�1P��d�"��m�n邥T��P1Y|~H�q�	6|��L��*�]}��8���L�'���.�VD�N��g�l}���a��r��'�)��˂�"�8�GљX!��!���RBX-3w	˽G?��{5�Oy��q�D��u���$�̼R>АT'��QG^9�I�>A0�'�@{�(��]�|=�N�ci0M�O��R�'�i��T��F_lE zeK�c���,�$n�Y�V�J�:�`�s���'Dh�%����/i��3�׺r2�H$晣9[L���iK(�լ\D=�t��#|0du�f��\�ҁ��1KW0���V�l@�E��	�FiKG�hԲ`�03 �m2v!J*��q�D�B%��I�2%���W�Vm���v&9qجSffN�+TlR��ʪlt�m�cg�:dg���%ףRd����Gڤ?|�=*Qb��v$΁wM�a�AϜ�9<��Ѡ�-O�C����၁��e�@[��	L��usTO֊Q2t��gIj��OX�A���8�MY&EmHa;��H��e[$O��1O2�$#�A�(�z1+ņ_� laƓ�T���	�|i�b��%�t ʀhS�\(h��k�(�bPp"	G�( R�,A:t}\��7�#�&�ڢb�3{��{�g�
{�,����r#4��@�ٱq� ؃��}��k�Bҝ3�=[��-�p��G���w(,����w�4�۲���{��#7B�U��IЩ%x\���Nb��D�M$�Sv�YD�i�u��h����=d�M)�a]�_�>��f��O(�{&a��G�q�J¬l���¼f�L���dϧc� {�	L���(��mN�t*�- ��<�F���Dt��FG#H��M�@	�*4ǋ�9D���4�	���Ғ A0Ct���äثH.�$���٠/
 Gxr#��[`� �N͸w�zh�d��1�~҇��ui��s�c�:�ՁeZ/5w�G�]�C5 P��!�^��b�����J�KZ�{� yR��Ǟs�
ma	�(&���>��m��gp���P���X���K4����HϠ~�:!���o�3�ۈM?������x�(	�� ����#J)������¼ ���&�,ժ�- 4$⧯Nu�D��Łf��4K�I�u�;���f@(J���5}e2�M�[8��;�AE a

h�w�'SZޔ����>gF(B� �7xQZuE�;]5���_T��e
/8G�@A\��x��E�+P�кd�~2���`���h��) X˳oH�Lh� �r��0��uN��>���dF��.�te���	\�t�/��Jc�$��������X	�4K��(�m�0T!3@C)e�l�s�'7,�=Aab>�:&iW4:�E��>d��L��e� �^��N�hD9�m^�MM�̸B�ΑI)�!�&�$��X�Cˢk��MZ�eвHT01�rmG���X3�9s]=��eR�*�V(�K�0�ԥ[E��KS8��mՁC�����;w[9�4Kі/�>q#a�E�� O�p����{�G	9\���:dE
�J�Faq��58|��ӕȜ,DZ�����2Q�1����z9>�Y0$I;6��S� ��	�Ԫ���C��[#˘�S �%�@H �0.�a�dh�=@�fP�4Q��g���VȊ����e�#�|�ƴa��-J�b x��P?5S��S�_/hY��� �2��t9���9C��uIF�)(��k��ؘB�\ r��C Yȅ��e�+��)rw�J�3@O���1
�$!�zA�!K+L�p��K_��q�V]���D�7���qJ�$&�da�qEK*A�\��+ݩ���A0J=�DR�!�?&mbE�$ 0�t���0��⑧W�1O�<���ХR��l� �2/�~ݳ�bH�PΤ�W(�T�q�RM<I"�p%aM�}��ܩ���)�z٣BH�S°���[�A�ҍ׽���`��AO �A�#T2F��P��#V7HŹ�+����l1Ĥ�"�#���(� W4k��"��9��x�2�
~Y�fʀ*�ȸ�@kH$-j��I��6n�
��"��
��p�����#q�-p��[�O	T�t�"B\��ł�'�a���XE� /(�yI��/w��KΟF��b���[b�h��K����sa�I�7E� �@W�Q��l�@��?`��1���$f�H����k1F)��8- �yu�Ɯ8��3#\*+�����Sxv̙�A�9Q2Ʃ��O�Y%gF:���(���F�X�^�(Vi�s(�S+�V�~��E�D�f��`g��<��U�>�dO-c�P����i�?  �#sČZ�-A?t�ĭJ!���~�a��+��k)\�P(�@�%yΘBѽ��eB7*���:Ի�N�69��k#.��]� ���ί�O��eO]�lq9�&j���a�[����F�k�<A�ʘ�gؐc BՌ#	b��'����F܂�japKT���sEl?��.����Z �͢�U6f4��'v� �%`�즹ڦ`L'g�Ĳ���g����t��9Rtq��FU�^BP8��Ċ0-2�3p�W�mj\��5$�boD� ���'M���eEW4d�4�IEg@�~�d��jO�\QxU[�OV���9O>a*�.��ʼ;�@�w�:��S�O�G�Td�P�L;r2�i'��j�����-ͶG.Y����v��
�D
?O��|S� RN�v�A'-�$O�r�QM�AL������%�Rǔ �L��LF����$�h��=
�H�*���`��CM��`��|4
��qFSq�<����f��\�Ћ�_(�l�$�Qs�m��9r6g�A�Z#}�����[������NF�ح���n�<���%
�0��ƍ8:S�
�_!�U�� �@�S��?Y�e�6r\zM�#!I��e���c�<��$(G���b�C�1�����T�<����
>PX�돹C`����z�<ɀcM 8�P�0vQ�5���Y��i�<�������d�5W�h���m�<Y�[�8�t!��ϓ�j��XAJ]�<q� ��uu��[1끰 ˞�2 �q�<��B�0>��aQl�/4��c��l�<A/́>�DБċȧ������n�<�������VA�
YĮ`p�L�f�<��������CdH�	ؒ�z�<�0�
Wp���#X�� ���C�<�mD����x����x�7J�z�<1���P4	�s���I�T�s��L�<a�LO9`�Q�ጇt��9��J�b�<!�Ӗ~r
�C�`��r��(BG%�b�<9$&\	Q^��p�kظ38R�@3��^�<y�i֢HZ�#�H��	�&ѳe	�w�<��(G+~| ��C�1qIz���Fo�<�F�^�V򀓴�����f�<A��H8�덿<JX�����J�<	j�R���r'�Hx(�qE��@�<�p�	i�"�Ѐ��a�\�j�b
B�<y�)L���)Cщ\�O��e�SK�~�<�GnٖV�N����}M�,
��a�<y���s�B��Hj�"����C_�<a���4#��}��U&0�$Q�6�V�<1��&h��t	��ԉS��x����[�<a�˜=�qF�ބ+�Nqb�Ci�<��H
���m���QE����B�<�C����"!9�K;Q�.��W�Yy�<��N�0g dq���� @t�<�ub�T� 5 ���)�9C"�p�<�5�!i>���u�K'R�
A{�$�p�<�V��� ���E)	��*怇o�<	�OKe`�F�B7
�x���a�<��-ʳ ܞ�r��;t봈r��3T���@��%W60�q���!�"y�f!#D�TX��<vV��vcM,l�Rq� D�l �j(��0��FF]6q�U�>D�l�4�_�(l�Db�N�M���A1�>D�1C�����*p�!j�e��a=D��R+ǦH��+�f�247Lɛ�L,D�d�C'DI���P��"Gw~��!D�ܲ��ŏS?uA��P@n� @�>D��uǞ�W�n�S�;II�h(D���O
R �J��R�f�\�׬-3}*�{��m�OX����]X���Qa�6*�
���>��	0���0�Y󣗫[��+���Q��'�jm[���>�NK�zp�d��Q��r�j�uH<���HUdLŨa�>�u����\���yf�"���C9|O� �#A�S26�I��(?nF � �'�$԰w��"O��1���}��BL�b/������4\�0�a���y�C�F`R,`HQ�Ka�%��3����OPd���h�J�OtZ(Tϝ\��0p�g����

�'yvY[uc����4�c�*![��y2'�P>�E`�+�=G�:�eʘ��Ϙ'��@��W�S=��C��&���{�3���;ҡi�|�Si�'7��D���Z���b��+P�Y:�H',l:9��펬7^�z�� �������G;�� ����G9��kY�4|�7��1Td8y!� ~r	�fO;�X�"��()��͂ ֥"V"O��
��Q4.�L!2�*��<(�@��E�+�M��Ԣ�±�s�L6mR��J�O�4��	oq�V�k�e� 5c�RE���z��`�1$I�	�4Y#�5�)�'p�n� �W�����<(�8�۔�����	����W��z�Ḧ��Ֆ9�����DJ�ت�k4�O5�~�7*Ĵe��
>G���I�h�i���'L�Z�ԑ:qY�)�t|k��"{ �LK$��:Z���S�j��bB�ҷ��Aۊ����+�	w�a���qƀT�d��Y���S�E�v$�!A�D	�����FX"H�t��X�~L��p�5!��9�kI ����m6w2"h*�-f!W�i�qOz����	�TQZI�va���ʐ�O�"�Vic%Y
b�L��)ͫT���O�W���H�̄�ڌ*U��|��LE0`.��؜w�h� ����up�D�'vh��J�u@>����~�#?U5l�CrIՍ���OP٘QC#Z;Z4�� [� ���+$��V�. ��D�M �m"P�ʼC@�Z�¡_6@V��i�س���Q�R��
�4�4CF/_�\��M�1k� �@�SK;vܢE�D(��+O(������X �O(�.��4�F5w+�h ��$��)�#Ϙ�qlD[��ȇ�b�[R�3;����AgF5t,��ֺ'��˓OY�x|\s��X�D���2��<�D`PiȽ2Ռ�v�z0@�� &'��|sf����M�.�c$<��������d	 ��DI޺k<�!���].$�q��ЎL��7�ǳG�X����1����|b���x1z�ݏ;7
1�E�̜lH&5�#iD�г�\!����`u�����ħ'��\3�M«uhj$���Vt���\H�T���A���!��צM�Kɞk�P�ص��:7���RǑ_��I"b��vJ=�!4!��Ale^k�Nu��/���	AO>�P��4�> ��/(*��+S�ըBo����E��	��$!���Q��u�&Y�*VrM����6���
-O�T�U��)#H���#*���D�/����pj8�ʬ���(����%u\��E��S]����Ö�rBqzr�>�L]��� ��[AC*ȸ�$�GMF.S�	Ӑ��a�H*EUtQ)FmHw�O�j5 ����q�Ab 	��g �Z�	�T�Y '��%�B��@P)V�~`�a��p�$i�d �2�wnr�	V��n���dKg�*�!e&c�XU+�'Y�(�%	k�gy�FWc�6TвN�y��Q��ciʬ�4nC�/�n��ghߧ3��fL[M�"d�B����q�H�@�@%D� /Ʊ�B�I�{	����� T�JP9��ܚ+�ث���)���W�̒UX%
��"jܫ�H%U4Pr3�F����&�|�Ly��e�4�`��!�xҡLl��Xq��<{���	�8bD�5Cף�ȉ��ƛ{��.F$��[�C2=�q�'�m�r��"�>�0����Cp�LV�ԋ]%��k��קW��8��1��W�V�� ��Q��ȟ���#
��h2ř!/JG�L�A�.8���Q�� �҄�����S�Y���4K�/HB�l@Q1�bEI��>c"�)�?f���`��qO��a��in�ɪ�7p�3��ʤP*�%����p��  �9 ڼlrEB�	�01G�^�?`�S"-��V&qOD���`���NB�%�Be�V�	I.���N��s�0H3∕$m^��T�U�G�R�qjT&bވ��ć��L�9�IĘQ�PMb�-�p=�@�2|h����BW�g"���#�h?Q��G���SqDX%(`�ؽ2�b�l�b)����胩�(���ڂ��� ��J��!��g�<����'��	��S%W���GN;-q>U"`��Q$i
�~���GR�����%�T�̨�.O�����4.�!E�G!K9�� ���z�����3�ΈK`�įp��;�m��&��1Cj��J�2�4{���@g$Հ6`X)s'���[/��
����-xW�τ�UP@�:Z�t��r�I�Q��{w��w�`7�U/P:PUl��k�>�������ʰ��0Vz %�֫:��O�yp_JZ��$�A�r`*�mء>�����·�!y�d�&`ږ5����I�l�2�'C�D�jLzFm�:����$N�-$s0`)�I�6���2�-k����2No"l��K��ᰤ�;k�LXCAڧ=_$��T�	
A�ˆŶ0�a�󅒿M��0D��k�FDK�!�$;R2��;m{��(A�m����.�=2x�'�!cp��I���eh�h4H�pa`�r�TF@.A��h��V����O�I��W�͏�l]�j�#���qQ�٭=������6��	"p��F�O����)ŤN��؊�"T��X����\=m�TD�I
-(/Bq�A�Ũ{-�����&J����B�Ԧ�N��"�>i�򐈃�2P�@�D���jf8q *�;@�S��ջF~钦S�'1�40E�Ĝ"{v�����t�|i�,�J�^ H���:Id� B�G�`�����ꅁVvn�ÔFO�r�xq�4V�@�@ꎍv��0���R�1�|�0���jo
��$�JS�'s�8ɳ-�-2�r��b�9ih��tG�=�P,��3\]�� �e����FE�l�zh���~ �HA��
�VfH�VM��0^U����f���*�ƅ�n�4h�g
`�n��%U-%���'~ �06��Y�@���ʣ(8$t"�gd�~��enխ$��Rョcy�}�˟G�m�D�'��S��7~��)�:J@�9���;7,�i�׫�F�q��D$���+d#����c�mG|b@�V�S���K2<�Vė� �pK��g$���oMj-"���U���J�y� y	e��7L=�v"6;���7l�rV8��cԲk%P�<�f��7?��Ӈl7Ya��r�R0`%�MB�OS�G�4L��&�9+d*=s�b��� �3$�ô]l�	�g*�m�R8A�6P��ڦ.	�݂�Q=tx�k��K���T�4�S��t� WΝ<7ȁ�0BߧJ�,A!� ���d�?DN� �����xҨ��nOx�ñ��˦�P��L9j�	�|<��2�fL,-�Y��4��XP� ����ʆ	����-iRh��Z#��8E�.5	 �^�#@44� b�,18@�S4ґ	��b$�#�����#;�J�D%�UZPD	���y��<��D�KQ>�eD�n����l>���C�#=P���4�q�&ƙ0>��E_;d_8�Ac�rfv�a)O�E��$ǏhK���E��M{w�O#R�s H��WP!��,qL����pX��Zb�0]��qt�s�<ac� jZy����� 8��6%� �V��O��<P�!Ɂr�2eCrk��jWE��� hW嘍H���a�Jh�v&K�HOx`�",ƌ �jI����>tsE�$.�xĀ�iW�U)��3f �!1f�M�V醄,�x�k�]�c �F�L<.�&ـ�z�\���lA9Ei�죢�R�|�ǨS�	��L��+�8���� ݼ�?� �K%k�2�ʳ�]���CH�:
��l�˂�:��5�A@�?;�(��@&�>�����bް5�yɡ��.Xg���h,�#�P�!\��F�>��O��Qe�6!���@���?�,QKIP��|3R�_�UR8q𰃋0����(��"���hUES9�S�	٦��$۶'2��7�
'i�]��lI�y[b3LO���7&�X���V�Kq0R"�W[��S��;TbE��g�#%��Y允�<�HܩS�w� 9r��~b�N�),����U~�c�	�t��ی�MJ`e��>\� �g��L/�ؔ��"VQ$�1"+�a@kq�>8z� j%eB�#��6��h�ɔf��rR�X�R�R�y��O�ġ�LՎBX�	���Y(���$T�h�f/QEj�82�ӑ6p�9[���Vh��X,���T�y�N	�,̦/M܁a��@�~0�h�$�p��d���]w���G���JF �ܟ�OJ�Jqa9����B�r�hD�����'�������(Z!>`'!�?SZ,��̦�3K)�r棍~�"y�E�ِU�D�2j�`<����J'Ye�zR�Q�-��v���)!T�3f���@Ł6�8��ccQ�'��\j޴G;�( ���q~|��$�IȐ�{ԃ�:�`�0�.��W�.ՉD�t�����l�� �0��qj�'T3Oh��J��=p
��	C
�avR�D�دFf�3� _�3��Y2&GձK`��R�V�ql��� ߣ)ĸ�#���B���)�GQ�a��Q��r=S�,L�p�쳖#�n�x$��b�d��+��m2�V��5�@�av@�}��c�o�t8Hc���g�d�4�(E�
��N {��Q���E�XC���7�@*�r!"��ڡ\V��I�,p� i��Q��z��e��;��y�D�K��V�Zoʤ�a
Yx�@
�G/\��E�Y�/��K3��9 � Db��Y���тn��6~�aB�c��B%N��5iY*��+��46�q�aF(U�X���nW!A08��[���a��F�> h�E��bJ p�!��~�	����Z�0
����MK�ON�xD��k��È P�®!��`3P'�n "��\�y(d8xw�*M��e��I�������8vSFAj�l��_;��3����u뢢�(0�kE?<���@�]7(#�p@B�c\����Aȟ
��U�b�I��Ml� �,đ��U���D�z�"*��k��ø!����	 ����`2��8@� �32�,/��2	��/�}a�M�t/��"�H�.�x���4;�<�bY+��<��дnEq�AJ[�[�Tb�� y��D�5��!��)A� ��|B@��hNU���Z�-Ȅ��HV�f���x4H�
%�	7�Ρ灇�p��R��{H�T�B�ȴT�� B&n2��Q��)��TK��"!g(�6cHJ�\�∉6S�� B�S�h9�0����*��q�I�^�ލ�C�	n12��	�H����g.U�iT\�	DH� ��Vǎ�2�h����ÿ!#�����h{��CS/�
l� �c�"O�^Ԁ����=0�b��m�|̓>z`Ea���l�b�3��&2UĘ�'��Ո
LIn��aGGέ,�n��M��y������K�up���2�Q�~U�h� U���Hq��bx��#��$�HhňK�����b�n�a�"&-ֹ��#��Qh��=r�"Rb�l�)AҌ^�g�v�C�!  &�6m�%��y �M	�ڑ�S�F��$�Ҍٰ`���$��C���� Ȇ`\�y��eh(Pq�<a�T`\4JQR����'���+��cZ�a��l!DYH�N�c�����(�f��4mR�=��������.���`p��1��}�����`�@S&L$L�� ��,��D�V"�7dq�6�^܁ �S�m�P� �M3B�h;��$ƿ)��)�jK�8��@�-V����	TX��q���a�n��g�a�5e�qa0�9�+�*}6�maPi�D��k�jS6in�"�'�r��)Tn�:e�0mG}r�F)P��I�C �д�I�����]f���4k�!u&��4��(E4v`����H��8'���OΒ�B$c�7Xl���d+��yW��Mі05�N<U��(t�!��'�*�tb\�u��9A*�]�'(TR)��6���xwN5	}�X��e0-\�3�؈t�L���*WT%��ž2����.��p�l̻M�H%W��~,��� ^���H��t�!�q!�3or�D$�ӷ9y�P0�%B��Uitɝ�F��������< q��F��D�	�R�iQ�Ȁ�P|1��1C���� 5�	*IҔ-H"Y|��"��U�4��ܴ�L���N�_,���VP����|�����tuhUi��n�b����Q�:�����-��`���G�&�<!�Oy,*�ъ{�a����
�&Ӹ����P�]��豤����1�Gh!%�E�M�ORDP2su�Ƃ0Y�����%��qGl)1�iO�X�JЫ�i�&k�P��E����h��B׽zr�����_NV2Q�0Z'*+p�ۧg,{'؁UǯMkp����!4z-��zcV�4�fp�P���pk1�O.=|ir��
��(���I��;%J]��X�sĄ�f�P=a���7Q��=Z�o<AF�MA�LD��mU���B�j�"Lߨ�R%NБ:��*��yT��hp�.x-�C!�,1}r�ş�"�J��V�9��rcgF�}\��XH<��d
&s�>�)6k�#Jdq����oK�LZ7�Cd�:<cDצ/>"t��
'r�"�Q�+C�"J`E�r���uIY���zT�������2s1����K�B.���Hٹ"< �<���Y�&(S�cY�
�"��&��-��7�}�p�N�d|+���
~x�3�Z'	n�D���!jj�hq��5�Eʰ�td)F�o�=�oT�d;e� &��fb�`�@�֥
�r<����z�@A{6C�lti���n�PM��'�[g� R���v�͈�zy8ɠ�Y�$�$�b�g[�O�Jy�W��2���{Z��%ۿ� z 0�/_�1P��'��#R�!�� ��Z�%��,]R�_�76`4hr/�)3S��'5er�p��8@�Z@�j	�,A~�0�,}"�[o� ��`�B$� ����A�8A�Rh��I�.Bx�H<⧗/hu����j�==!Z\���M%tb���H�-�2��C"MY�h��/iv����ʃ�?'T\ɴ��٣�q���
���U,Aw��$&���@7.��4q:�	��S�w2`@j�}¤]�� ʇ��5���[Ԣ�2x�ɋ6/L�jm9�?F%�뗁Y�m���D�V����sdb�1}�ś^w�&��5�-}��З�/�.]3A�*� 镌SM�'��y��O�	\�Y�V"J?@h!bkX����I�/���m3�d[2��E���R#��D	%ߘi�5�J���犉ɲ������\^�CSa�% �M�'ٟ��E�U�4��D�?+S��q�%!Z��n:�/R�>�2�������F� \�X��i��1����]l����+EM�g̓wh�t0�'�%�b8����
'�
�H�FNGr�jrOS?�e�%��<I�烷PGZ����[�r�����^�VtE�E� �8��eJG�.��zbcS\�&5@��7:q��X�(��e64����Ңàd�S�J��¤l�C�
�e� Rv�'����AM�gt�18���eӖ�IE؞4(��n��)�࠘�.� Q�a�˺2� ��!�Z����'0U�d�_�g���'��b���To8=�d��H��҂ J �l�;�� 5"Oι�Am�l5�0�揊-,��c��+��y�F���O
��bO	5|��f�	��`��"OT��F���q O
��%V"O�dk��Am��!i@ Ѝ\S
�yP"O��d�ԓv�p�/Ȼd�t�rC"O@Q�ɍ�
�6�y�G>s[���R"O�J��"6�Y��.MF����"OV��v�Na�e�5g�k�F��!"O��$���6�ҩ�E��;O��4`e"O`I3�
F5����m)Y��I�3"O6 )���J��B�l�rL�٠"O���䅀#���J%O��Yj0"Ol�5/�̨��0Ǒ"tŪ�"O��b�hд'��ۗG1Nf,U�u"O�򷢝*J��� V�E'DLb���"O1��쁺?�>}qn%a���"O&\���ۮe��Ŋ$��#
j�i�`"O^%âN�,F�B1e�ݦ	�%c!"O��J��B�ad%+@�C�|��"O��#�'F�)����%�H� #��@c"Oa��lQ�N]zb�ʄ[�\dK "O���� ��@&��Q�剫`�r�;�"O�1a$���1��35Ò�~�,�Y6"OB�P`��"X)����[�E��zq"O��c@�; ܖ�����l���"O���K
�cV^-��f�&+(�"O�E��g0v�Ve�f
V�&t���	�.�k�O�i�b��A���ҳ4ܳ@Ø���ЙQ"9#�a�� 6���Ȧ2#�O��ӂ��C"�	�$�/&	���:,834b�Цar�%��"@a��E<uK~�Ya���U6���.]V�[�ėڦU�G���^V��S�O�ij�l9>S]�ڞ�)�w���i*�G�#k��S>�@H�"=?��TkCf)���&I\ʦmY��G��y��0�&�G��e �TkL4���:a^��7KJ�E��C��d������z����OU����,�$H:���_3��9G5O��ʠj�$#m"����4��{���|���C�u�ʵX�#@=7<��.��?1�Y��|�����&���3����f�Φ}����}W�=�p��?�.�)�x%��g�}P|�;`U}x�@2~�|��<'�N�=�O�HH۶dY����v�(1R�TJ6��Q��B�Qc�0�ǧ	�f,���X�NDإ�wNUk��)���0q*��<s��\�h�B�: *R�K>��P0Rf i�.� Q���C�N��I�<��I��uG�7<�%�qZ))���򁍑o���y��v�6%�7^?�5:��O�������FiK�h�&"���z��oݛ&B��m���T��_��'Q�J|���L�"IB�UMT5n���ó�M�@	 ���B���x#���w�@����-F�J狄�Ni����J$m�J��rD�<�7bl>��!�*Y�x��$-
	Z��HD�1(���0<y��"��`3G֨UҸ��`bS�jVZ$�`��tss�&dԮ�@D�6�nx�֌���)��CR�k>�H�?O���w*ڂ(=&q����"~"4A��$���ɚU;ĩ���ȾB��X�j�j��]�0|� ^��#�߱G��e�Hò�r���8s�sԑ�`���!�pk�F+3�x�J3&B���!A7fX�IfM�4bW�#�3�	�����/�i�l��PH�<�`C�	�\p��$��<5SlLbE�2�"C�	^&6�:��O"i�:,�E�B�F�
C�I�2A��@�.5m?֜C�\�3ϠC�	w�%� H�+|���x�A�4M�(C�I�r^=��J��<�|�#� ��DC�	X��R>H|����Ռo�C�	�8�q;4�'I�ts��3Z��C��&.0�0U��;[f��SK��s��B��^��`ӁJ�T�*���P!M��B�	�f-�����],�����"��OƜB䉍g����AN��)�V�����L�pB�I���� �T;2�h����3�hB�I"8	������Y#N}!2K�%@B�	9�ء0w-և.�����
~�B��E���r�f��xm��&�� ��B�IqX�2V�� �4���q��C䉈T� �������f�`�՛��C�	�K�rԱ���7�Vu����7VC��4<!�I����X��5f%�%,�TC�*,����N�� ]�$a�.�bN>C�#�h��9`��<B!bE��C�]�����A�s)���%��I��B��?:^y*"@�!5bT ��^\��B��
f]�H���9Q~���Q�SC�	${n��%�L)Jѡ�a��l�C�I����SU�<i�*YZ�MΝ9s�B�	C�p��� ��pk��(~P�C�Im�n���"�i�0��p C�ɔ��l�D��HI� G�Jn��B�I�L�I�� Q��)@��*H�B�	[W\e��-��D@��Cc).�B�	�?�HX��P�'���aaJ�k��B�I�¦�j�-_���@];n�B�	� �d�4�U��B(�0�ضtbB�� o:��SG*L�.���iWG�^B��),�}h�C<ye���'C>B�I4�����CÀE��q��l�>D�B�="�:9�u-ڥQ��q�d�]'eD�C�zɂ�ۣ�ۣ-���U,�*-BXB䉜&ł S�&I:y��kwHPc�pB�	;`��l0*��H�\@D,<}�6B�	4+U��0c�? �Ȑ��*?5B�ɊQrV� ���(����/[6��B�	�P�8�:�7RzCKi�rC�ɨ?��D�H6/2�ܺ"�U�D��C��'.��!�j�'��B,$|��C��CM@0XꟖS���QvMN�V!hB�I� ���N�gu���v��Y�rB�b��ZtG��=]�yS�Զ+h�C�I�*��Uk &A9	�<�#å����C�	��Y��,��^��c��N7�C�ɭ
�Y� M�t�`�KK?=�B�*Y��A�Ø�Jx&I���ʑ��B��$"𤱩֎��y/�C@T=w��B��6tx�n�i�(qӕ�S88QlC�	�y�^@����Y$=�U/�z�.C�"��h��e���P�~�C�I�+�8���O<i�XI���/\�B�Ɏw`�ī K�(��,X��<�vB�	�+�tE[�N1������jB��&\���W�#h�@$+�$ݘoB�)� ؝�2�ɹ/e�*e!���|�a�"O�|���rf�DAt���j'"O�Y�խ�A��r��*�截"O���gL�6�
$af�1�M""O�Y�F>,&��׊A+E�G"O�8;��ڬ`�*$�`)m�"O����m��<�@N1�fL!g"O�l�G�L6[ǦHʥ,�5��-��"O�,�`�9�v�!�U?W��ع"O�DRRkL.J|Э�"�i<2�"O*)y�lׯ_�"m��]t0#B"O�C�ꊋ,�.�#�R�x���"O�Swf٦_;���"Ǟ ,A*�*�"O���AF�����u�(~Ύ���"O���V-8��-��V���2"O���
�N�����*׈^�B=+6"Ob�!O�$Ѯm� C_�i�7"OuC��:E���"YK�9�"O�@P�͐�)��ዠ#�N��XP"O��҈����h�+C��08�"O���B@�B�R�� EG�#/��h�"O�����?�0ю�� @�j�"O��2Uo�ĺ|@�׬  zG"O)p�U�]`��G��m��=��"O�i;PcŎ/s8�iWfX�E8D"O��:�j�P�x���EJ�+1�a�1"OƩ�t�_Hx�����d�d8�"O.`"a$Z<;�RXP�H� 0�)�"O�ثr�Ł''�A3s�X�/��E"O@��gX8�,]%ԕ��"O�I7���4�:!�V��}�p$��"O�@t��#f�6�b�A�%�*���"O�uy�k�'%$��ɖ�
�`�vS�"O���F�F"I�&yⴊ	 J �r�"O�]�E�ź-���r��PB�(y�"Op}�eě� J��"C�?1@T�r"O�������ا"_�M��肕"O��/�RZ�+�l�0ep�q�"OF2�bN�w�I�*�+)g<�"O�!v"�k���{�NE45@���"Op92���E�,¢�˴HI��"O���Fv��X��;G�p0"Ox�FHC�nL褨�"\����b"O&)��"�-L'hG�4z>u�1"O<b !S�{D� �Q
�1�mJ�"O����I��<��4h�II5p��s"O����+d��iŹ2 Z|Cb"Oxm 3N�3�����!*G�-�q"O&��&���/#�dRt�E1�Q��"O{qф*ix  tM�"vb�"O`�B n@&r/����S!S>���a"On0B0MF:�<�B�ҟbM�1"O��!�C�?��5�%���HE"O�:���R2�z�MћTNY�"O�]Y����,w
!�pL�i���r"OIB��?��1t��>����#"ORP�E�ŋ5��S�*Қ�%�!"O\M���6�=r����]��"O�L17(�G��$1'	��XM�p"O���IA�#�!��|�X��C"Od��bΎus�P3��E`�Rф"O"�y�Hw��ao�(�&p�2"O`�0��dȪd����l�Z))V"O�-i�A�����_�B#�"O� �l����;�8!w�:��A�"O\jf��D'z%qC�Hy�~�B"O0�p��HA�ތ�#�ƉL���"OdȢ�"w�����6J'4���"O��yR��}u��Y�-ΰ8<�"Oҡ20��
�4홒c� 8�B"O��f��Tw0�Y6cO�`�P��"O��a䄙+B��%1f$\�P�h�"O�5k�Π�Hz���9�z���"O�
FĿj�z����	t��ܰ�"O���D�{C0��1��	��� "O�� �@H.iWjMy�h�Bs"O�I�$/��8��Yҕ�l	xƎG��yr���	�p�P��_�Z�#�(؟�yR�!vhTz�CēQՐ\;���y�n�* p���L�R�KA��yb�.7,�b#g
@K��8���yb���	J�it+��p��'n��y2h�"#��kW�U/|l�+�솆�y�Lt:e�5�z#��;E�1�y��ɴ8�������k԰i$�"�y
����ũWK��c�%Q���y2%K&t����膶-�T)� a��y��գlq�%j� .����b;�y�
�f���p��
�����ǎ��y���h8��E�H�&.�gh#�y��p;�h#�N�$��11���y�O�#������	o�N�1Ό��yr� �߄�P��M�9�P���%ܮ�y��i��ѣ�2~�z���,��y"�9*Y��paj.�I�`���y�A**��a��ؕ��s�D��y�C�0u��;�e� #�}��Q��y#߃o�lH+$�!|�V�{t�΀�y�LL����C�J#af�bdeO4�y2j@�dbL�%��YFF`����3�y� �5*y�ӭK*TMX��qG.�yR�׷u7�ȳA��9�2]�`�M��y"hO:^�d�k�O8ľ��P
?�y��63�l9$!O74#X�YЩ�6�y�n��~�(0;�K���P!	��y�d��<�T�����#�a6�y2�	&�@�� �{.�˦�ט�y����D���J�|Q~�9'�P��y2�>a�I�Ћ�? �(�%�^#�yB��l�k�ɋҡ�G���y��֕vӾY�0��"����'$&�yR��2d a���S6; `G*���y���~e���O�X������yR)�5)sԃ��@�"��#N�4�yr$_�t�"��v��>E��t��yr̓rԼtb�h�n&�|�SO���y�m+*Bݘ�)c��u�c.J��y��{-�a+`�\��x�-��yBLO�X��Dy���b�)8����yl� tbE- q��	�����y⣆($��8w!Urmʝ�'Bʀ�y2c)T�~  ��)t���R����y��ى�@]���L5r������y"��Q��=��+�'�����K��yR���r
�T"���%PT�c��Ǌ�y�={����Bg£;`�R".]��y�O��Ri�A�V芐C �Q�T/�yB�y�P9 f� ��)SA�ζ�y
� �|��cY �& �N�:G:�I"O�]yp�E�EV�(g��[�,��"OHp��K>0�n�SEM��b�>�k�"O�U��*@���52��тc�<�S�"O
L
� H��N��l�
<?:e
A"O���a�
?W�6�R3ˌ�3�6��"O�xkؘE+��SFϑY���s�)D�@�g�    �P   �
  �  K  �!  �(  )1  l7  �=  D  GJ  �Q  ZX  �^  �d  9k  |q  �w  ~  ��   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dl���2<O�1"�'"d�p&$�#f�<b�FX �~���$P�0�ȡS5�ʸ?8V�媜.�u� G�~�dM�r�Th o,�DS�F�"`���d�%�]pv���ZFZ-���[!k��ם�y����џ��.��:e����@������h�^!I�
R�?���kư�{��-K��6mB.D4B�'e2�'��c�c��Sw
B�y�=z`/Z#,��'���c�Dx��	��*G@^�?����0҅�Y�R{�1�0�C#H�Z�Ƈ�����ן0�	ݟ�)r F����N�OX�I�?����6j䬃��-������Tu��\ϓ5��@�`F���^yɤ�Țn���'��+�$���{� ]*��?3��  ���;QfZ�� k�N����O����O����O����Oʧ�y���h1��0��V M�6d��?��i� 7���ᩪO �l�+���xش�$1��� ��!`�	��#׀�Aa��q��R�����������Q���<;�� �$�>2)�`3���Q��]��#�THb�o�-�M�e�i����O��I�J�D>H]I��'1T���������t��-��#�5p��H"V�(�(�J>�j��ɦ%��4]��V�X�~�n���fι�Qs�Ow��3�ߌG/~|XV;�MC�i��6m�?�X��D�h��at��(S��|�B����pATN65�����b@.�*�� H�6A�D�oZ�Mۅ�i5$O�'r��qբS���Am�l�h�R�#�]�p������G�(�P��!�F�m��6d�r�9�IZ+������L?@�*�/&N�y�	_��?��InѪղi����\,r�P��P���RK�#.���<����?��O{BU��)�?}ɲ�±}����y+�<e�L����a�Ti�S�'�x)Ң�)s�܂�L{�� �,���鑧ľ`�b��#���0<�ħ�ٟ`��=��Dj���ɰa�k�,��eǜ�R���'R��)q�X�0��B4��d)�1=��u�.�O=lZ�m�4x� ��Q �j�ΆO*�5�޴��$�	_�tn�ʭ��H��DB�t����²M�R�;��T�[�	 ���Xr"�'H�1Ɇ�'Y����(���	�f�B��DA�%!�0��3��j-D�K�@%Z����	ѳ�h����@�"�\)���Dx|�q���J���OX�l�5��O��?���Z�
�|un��ņ"P�S��'>R�'i�I�.||Sa��h6|��k!  ��=��` ��Oy":��`#��)n�6���▤���g�'\�e��d��Q�`�`D$�ڠ��DZ�JU� �;D�d9����!�0č;.�baA��9D�L� ��c@F�'�,QXv�3D����6j�x���	3,���R�3D�,r� G��Pr1���O5�H�4D�tPD�D�%F=��j�QJ�<���o8�S���JI���&-V&u��`U�$D�<��L�:}�4ų�J�#�8����"D��sC�\�p�f��$�|hI��>D� @�76�q$OɒP���Į;D��PL�mE$��A�Gp6`S��:<Ohrt%�Ǧa���4XR���d�ѣH�S���B�h�I2Qʊ$�ID��<�R��H�Ϧ�B��
_,#�L��\z�e��q�	�'BP��0<	VܛUl遰�]'&�rh���+�����ȏ\P��B �-)�2<��ɜ?G����O�hm����Z�Uǚ�¡��9l�|�`H�FyR�'��OQ>�F��XV�\�fϙmԱx�I>��Z}r���MsקD|l�P�n�e ��g�_�x�v�|B�θ
iӵ������P�F�up)P S�9zf��X�y"K
;yGFQӔ���]{�bS��y�,��|e��������A��˽�yr�{���xc�]�wn��J#j��y" Ώz�樃�K�9p:�Ec��U��yH^�!����j��?�Rj ̠	��V�|R�N�F�4�'��'���NH�#�d92��Q0�B�N�� (�#�&�M[4�iU�S�޷ �S9��'��p�mB�#��'�X�0m�T=i��`��@�q�h�,����O����VM?�@)��C� \����)uFPI����M��X�@�3��Ob>�d�O^�$��N�H*�bA�{^����
/¨��dYt�m���K��L�����#B���'�7����1&���?і'\lU��`�n0i�V���b��{���t�����'+R�'�B@l�A��ɟ�̧ج�uK.��� �'?����+��k�4�ѱKضQ#�x@	�B�� Pw/�&V�
��FZ��Lh��e�C��S���1q v��ϓ@��{��
�7U�̡Tc^;9Jn��Ɂßh�	՟��?	���T*?p�H���!V��lr&��~ !���,�m���S�	9�5�'&�$_��'�R6m�Ob˓ �u8��ih�S�kc��a��G�h�NI���JmQd��<Q���?���7%����$�!f� ౑`֏�y
� ����nW;2�����2w�ʴ8��'�\��	[�v�-�H2�y�䊋i�&��O�-DH����Ə�0<&iN���8�4�?Y��k��\*�;_YR�����5Tn�H��?9��?Q��䧵�'�� b�ǝT�V\�1��5�D��#j�,ȧ#n�j&+ p40�Qd®�?�.O��aGզI�I؟`�O�|��%�'W0�#�N?-DI!�T��R1�'��C^8h��p��)6&��	K��(S� *����cV,k��-��܊ �S	9f�24�����52��EW~��R�o~<�O���ɒ$P�8����a\�=���O��;��'#�7�Un�O��)��N�.��� �e��6#��	�'�2A* ��Ԭ��/�J��TЏ�D_G�OB"zs��#
�Vϕ���m�2�in��'�R�A&z��	��'"�'�"5�v��!��	W�m꣡���p��۷=ǲ���aU=zTX�771�1OX\�# ��)������	�4s�E�-w���3e�\��@���(751�1O �4+^�$ʌ�*�R�0@�л��'%��%�~��'�ў�2���s���3ǉ=U��+�^�<)�>��E�׬7$(ɰ�!�Sy�� ��|����$I&x�Ո�区
��(x�L>?2��!C]��$�OJ�$�OѬ��?����$DC7p�&qi�	�<Af8ԡEƣ�����'���H0e��z���x� �0!#}�g*�MS�8���d+��bA�'T�8�t'�~"�a�!i�<.NZ6Ĉ;�?9��'6��PG��+6fB<�P�%Xr��ߓ��'|��)�G��$�f�A !ðUo�T�K>���i��'��-!��}�N���O�ĻCiҜS��p�0Eˑ�X�	�d�O�drS��$�O��$Rg���<Y�w戍ӣ�=j�.�b"��G�y�
ÓX4��T&�C�̡{뎌�?�GkJ4=����/�*�c�m[V��YdG�Otum7��d�y1 X��#˕V)�p�LO�{ �	ޟ��G��i�1i�d��㝖RԘ��͟0�'ў�S�?)a/l�6��� 7;�X�5)�蟨�'�658��>I��?��'�Ȥ{�X��������(���3(?��{��?���.1���c�8E�<����%���ST���c�8qэ��v���c5]D�ɝ%vf}�PG�(P�B���
͒W�Eq�G��s�������?i���5Ez:)ٳ�,��"��&?Y�g�8+�4.�F�'�>a��K��{u�x:GgۺXk���q�&���O����O�˓�?�Ο��r5`�i`�S��l�Py�V�	?�M��i��' �h1qA��[C�9s�š�X�#6�h�,�D�O>�dV�$Φ�ieB�Ov���OF�d��, s�
ɨ�Zg��]肥IJ�"�Z���u2�p˕S�j̺N<9�ϐ�UC`��-�q,�9/�Q�`�I�U}�1�XS�b��08ʧ*��ԪflLҼ�»�8��$�/ }L��!�T�M+��i�2+ S���Y�$��2m%V8P&��y��J�Ψ'ȑ�Iß��'�r��>�Ǔ �
Ms�DΨO>�u2��sy¢n�@nf�	|��^���'�!�J���H�2G�ԥr���/E������ߟ��	矸�ɣ�u��'��?���Cd�̼g��x��V�y>�}�1�L�.f��$4�����fW�'���!AA��(O��۴�	�#�LA�	<�封�>ob��H �B�8���֔!NpY�eA���(OJt9�ל`�\�u��!��Ƀ�K`�X�Gz��5B�l�C.�ڝ(4	]*.B��i�-�4��ɏنXR�|�/pӰ�D�<i��^�x����\�iS=�0�[��@&*ܛs�����	�0�����|�'�؅p���s�H���X#Y��]0#��
b+��1U��h��i�
�||iE�'ʓ~+�<H��[�P�f�$3⤀$h�)}eT�dK���\�-��z�DI���8�J	�u�	��M�*�P;��!��$B���R�ۮ-��&�@��	�y�Ց��̺N�2��B������Y��8a\���!��sئ���Ol⟈ID�$§�y%�4df�qi���R-ĭ!�d5�y"ꗷּYpd��9J���0�F��y��!�H��r.��5q&��\��ȓ9r�(��$(	p�+"��wQ̤�ȓ0B��b�R�+%ȸ"���2v�l4��4F�@2Sc^1=���R$�,4�B��ɛL�"<E��灦HQX����ɬaDp:wk�}�<y�I�-�T�@��>�*<U�}�<'���M72���+�����.�n�<	��(���y��&i�&��#��<f"K"Α3b-SY�D��![|�<A�=L�\�����~�ʌ1�-DOyi�'�p>I�`Ba��%���ҌȀ���]r�<� nX��Z�#Ǻ�H���9��$A4"OڥKR%S�t4�A W�ڍe�<�q"OR4z$Iv:���ٝy��U�"O�B��݄HbXQү;T�ـE�'j�${�'�8�A1!�-R2�q �.a,8��'TX���^!lg>y!�c�.��di�'@�@a`�8(��Q�3NT1:�$A2�'�6�A�ڳpX��`F�X*:���
�'  ��k{��A֯�q�TA9
�'|
�[v���:
�!�N�;l�:� ���� =	Q?��5�V7X��`0�lظe��� `k!D����U3'�s��ќ{����P*>D����@	U�,����pl�ȃ@"D�ܙ��Z�IFT�S0�L�b3(t�"D��U%�w�4�A���Y.�# �"D�L��(�:��aId�#!RQ��L�O�mS��)�`b ����:�H���G��K}����'�*�8t�:��Ӷ��>7��h�'{���Ϗ�#�\��vC��*s�\��'�$�Y7�8v�>ђF���<k�'���� 	�,q�����(8F�@�'����/��%՘����˥?�+.Oh��A�'R V*ÙqN���"���(�
�'��=s��*R|��$��r=LE�	�'%�i�� @�ڙ���9t���	�'&u��CD(-�
hz3LU�e���	�'�0ݣ$��'xsZ�m#.��M���'8�@�'G�rr.�/���BkJ�aۖ|z�'%¡��bƛeh<0�(S�Kǜ0x�'���B��F({9h��`� wņX�'R"s�*�(�V}A�G�)9�註�'�.�`�H�#4�I"�3|T��'Lغ�b�D�����q���k��DF�lIQ?5�(�Rx��Ë�+X��c�4D����I&�zux�l�.*%r���E.D�8[fG%�, B�z���Q�,D�(Q���VT�4A�Q��mrA�8D���عt �S&)�q^�Y��2D�d
��5���"ͰI�<���O�Ă��)�'P:�a�����hV��gOS&/��@�'`���H�� H�E��'Lh��'E"<� ����x�FD���l<k�'#RX���ւ��XZ���r�^Es�'�8�4%O#En<t���f<��k�'�p�����cq�"��Ԇ	���K,Or8���'_�=+g�CJ��l{��Ȁ{�f8�'Z���S�J�1� B��r��p��'�P����3��A�&�N �ܐ
�'vY2�bN�"T�ͺ�jA}���
�'c~��a"";(t��!]��Y�"s�t�#�5�c�O�/�,@��Ш:�v��ȓji�T95��WK��p�*_�����<�u0�*Q.�����ND�-�>��ȓ`-,,B�JVU�Qx�b��K�⹄ȓxpz��7/�&.LL(��@7����2�`݂�B��v=���/��S�L�E{"hӘ������g�B3#�ꥑG�		lʀ�"O^{��W�#-:ղ�ȐF�b�Z%"O��S�,ݰ>^�ݨ��!Cx�ē�"O�$HB��d���RG�h`��"O��sV#,4����PL�z��Y6"O�q����j~��Ɇ��ifUC3�'S�\Q������)��L"0u 0�c^!`�D��ȓ#���L9f�ֈ{�"�'SH-��S�? .��.�>Ax�N/A�쪆"O�Z��ڏyH�fT?j �W"O��A��5]��X����,b��[#"O��X���=�<8����lha٧_��	O1�ON���o�.J]�����|�0��"O����#�!G��)&�F7#�B�P�"O�E�AV
A�	'�˸pF�PR"OZ�C�O9gZݭ ���A�^=�y��>%��$`�&D/�Љ@�ɞ��>q�ha?	d�s�J0!'ß~j Xs�Sb�<�1�S%?�Bi���
B4�5�e�]�<ٕ�l��DZte^7��`�"&QX�<������`�׫@�c�`�Kl�R�<�A�7YA��cD	�.V2�˵.�Q�<Y5`ƾ{�`��
9 6q6�O�'���c�����}�J���&�y��p�����!�$g�
��&#�b������3I�!���_� 	
4�V���*a�<�!��� fU^̙P�$,y�9bAU�!�HI��\�f��
[r4��u� t�!��5#-4A�-��Krb�)��!!�"�̫�O?��%]�R�X̀ǄK3L�t`�*�v�<iSi�V���F@^�
�H����]�<��NKH�)�q(�'.��q�l�c�<��ɔ4t
A��eL�Y�$��d�<��h�}��QI'�Ra`3b�\�<I*Au���:e�J�G
I�B�YyBK��p>�3�)'�F�B�r��%X7'�W�<	���T�:B�Y*d'n��1�R�<1��F����c�=��̂%n�P�<A��,(��BR�֕V�zLk���J�<�0���GށC5&ҝx���:���Ix�d�p`������C��V�TK
7 �Bŀ��5D�T��?lsbɹ�j�U$���4D�lac��D�^�c�OKЭ+T5D�� �I_�:EKv�
3����J.D�$锊Z*��脥Y�\4�9�0D�@s�cD\%��Oݰ~)>)hb�-ړI/�D�䧏�� ��!�vUl�G��y�[�3X�e��
i� ى��6�yb'I"���1�)]SX �1	���y�	�<'�8��l�m;*-Pq��y2(��a��,k��J%dy\1�-�,�y"��%�����&�1`S"��?�� a����:k�j�h�4`խ[[u���d=D��i'���8H�}�G��M��8@�<D�`����K�V�*V�siYW�=D��S0c���Ġ6���G���gc>D�٣�ͺp� �`1FQ:0�r	�A�9D�Xv�ţ�p�KkS���Љ���<92��S8����m�:��f��", bhJ�+T�l�d�4R:���B��H��U6"O����>7p���b��xy�p"OL����;(�H]Z�ؿi�C�"ON��f�/i\�`f���Tc�,� �'�P�H�'�Td��&�6#�� e�C*ɲ(`�'�䜀w����L�fE\�1by�ȓK=x%���\&Zkx�ë���݇ȓ",ZdA�f\V��be��F�ȓ<4�L^�0!D����t�ȓ�.(s�U1I~���"��E?R�F{�DY���f|�A�Rz��JN �Z�0�"O�;�J��3O�h)��օ��0"O��%b��K��9C�X8�
�ID"O� N��H��o�� �3�v��"O��	&U&z��/ˠ=͆�"7"O�}�b%�
<� �Ҡ�-Q��j��'�|U;���~��4�Dȥo�<���DLHN�ȓ�rEB�
��8H�H��2,f}�ȓ4�@͉QH��k�.| ���23��a�ȓ:��d��
�~�]X��9F]0���9S"4�`(*8��)HP��9]�
ć�-���K�_I�f�Q6�ŵdu�ٗ'���`�'�t1j��8���v��ҩ�ȓ
�pc7�� A�bi�&�M*1ZH��J�X@��ȤV����j�]��1�ȓ *j@�wlD �*���iW0OT�i��P�"�-��{��`}R�gPx���v����BցN�ՙ$"]�|a���o%D���P̗150dY H!q鮄��"D� �J�=Z���(�y�rx�.D��P��؎B����Y�z�z!:��0D�|JGI�3�� )]Z"H�H�N3D� �uȔ����˙�?]����.��e/�''�ԝ(6!��{|�ҠSw����UQ�L;D��r`���^t��ȓ�8Y�!��7�@B�
�F�N��ȓY��(��@Ah�"���Ů��'���*� ��P�P�&NT*	a����Q" <�!��2"��Y0c	C�J��=�	�gM�#<E��䇘)c�� �Q�6$x�3�`��B"Ol!�0b �{>�׀\G	�@�D"O
U����Rha���D�f�`��q"Od����5��`Cf�	1M����"O�m��(_|��!�R #d��TQWO��F싱;�r@���۝�����OF�'��	��'�r̋@)FԦ�@B��?��S�]ƴ����1{��Zc�P f�P�Ƀr#�4��ퟄ�I�u�\�Q��ʈ[;���V˒E�'(������H�L��h��G[4X���E|@��$q�/�w{(����KB`��3Z�l����-b� u�"�f�'��I����|�s!�<�r��DC�0U�pR&�hyr�'��Rĩ����z�ƺe�JTq�a剬+�dH�W�D?1�Nc�ȗQ[f� �օ�x�����Wbh�թP�e�v�׭~�<��Z��t�R˒7b�V ℊK�< ��6����Gh�m�QC&ZOrP��W(�uhY�,�v��L V� B�	M�A��K_�'�\%蒡
w��B�I�g�\1`�1j��dx��1f� ȁ��{��~"b	� E�u�ͣ@Х
P����y�A
%���+W��8�U�"ߊ�y�B**��x��J�';{�-�����y�o[�@H�@yA��J��P���y�J$0��C���,J��� s�R��y"��ce� Ӯ�k=��P���?��)�M���q�G&U�n��({x>A@@;D�y1�8p�b�W*�30��+��-D�����=yV$y��e83�DaSD�5D�C�H�b�8S�Ϳ*�>-�n5D�9�ǀE�4����<��5��.|O2�2��>AB���0u;�g0d�~D����d�<aD�8&2��5i�>b,hأ c�<	�ǓjY6p��(;D~�`����J�<�r��ih8���J71����R�SC�<)T�LiH�qڅ`˴g��D:bH@�<ɔc\&�M�$O7YȊ�#� ��'{�i���~��F�E+2��6N]�1� |i@�h�<�5AמN �0uabZD��	�d�<!���u�F0+�V�_%	�Ea�<� p9����1�0� EA�*[@��
�"O�������B'g~�	�'��}ztiĠc�4��H��o�&��ƤX�'"�>�	 �@8����=
$P�fBB�	�u��{U��[���vi��rrB�I���d� �NL�l-�$��c��C�6_��t��@�H�F-��\��C��k��q8�g�2;p	 d�)1�C�I�r?`�H��}��Dj�.�+���1k��~�ɥz	�т�g�e�� ���yB�ݠ_ֽ��j�i�f�PI�	�y�O�I�@�HP�*+�ԩ�G)�y2Q&sS��㎝%q�*� �-�yb�O��<���j�ع��c˘��O�L�֋�Φy�Iǟ��'00�JI��'��	k���4���yӐd2���O��D�OJ��B��Oxc�擫s����O=HG>��%��v.>">I�(�F�Ow6�3����,��1�'G!aЈXQ��n� �I���Ox��i�iO+-a�lp�[�RN Ly�'������5G�9����PJ���k��I7 ��oيA=�i���=EN���?�����|�����YZ@7�ǆ4��9MZdџ0p���<`����2S�2,��K�BF�Ot	��x������O7�0�4��RI�U�G�ڼO�����O��K��\�O�s�̨!d�&v/:� "�H���U��$T��'��'p޽K�\YI| f�=Y`����0 1��ab�'e���S��y���$�F�)S�ìMI�p#'H�\d�%�M�ԫI��*�F3}rD�~��-T*~�V�;���^��U���K���:}�k֗��RM��h�	i�H�dn�Rɺ ��Ox��F�>ѥ�>q��RF�DS��!Sq�V��(l����E���@�<��RQ�D�\�OJ���e�
-N��]��b��䴟D�u-}*���B�]�	,9��x1"57�XE@ࣃ;#A��C��Hy2�����'$DD��,�MM"yt��;M��zV��?�4D��p25dP��|'?�;}����I�lD��� ��iC\�c8��d����?��m�r��@ӷ.�N�X$��\�<1Aɜ
{b�X�p�݀0�<�Z�K�����Iџ�'/��'A�	f�\c����$��.9��,q�;c6���4�?�-O@��F�4�'F���$�\�Y+,�2������PQP&��ē�?q��OH�MJ�5Q�A�G_n���B���ȓ-�x<�B�W1�0�A�b
�}�(�ȓ6#���A�M��})BM>Gz���ȓ^��[!H�K��9%�V0v"�M��c�Ddq���6r���_+?3����SF D�e�K	�����H&>lpt�ȓh����B���J�VE��B-lf���X(����r�|\#�+ا-�1��L����h�n(�)ǝ�|�1�ȓ%Դ!�⎔/"��֍I�/�|Fx2"4�S���~E�4'�3rGpDp&+إ�y"�W{���d��m�����9��'�v5�2��]�)C@��]�=�7�U�'���:a�G�x�[��.o���a��&f�EŻ���/�%��!!�kȨL���4[��#���
�Z���/&<�)�@ޢ	�����o]9b��#Cќx�]z�K	<5���0A� F�`��R�'�l8�0�З2,QjشF�܌J�C�+k��}��`Hx9��hT�'_"��zmLT��E2�T>��O*8X�������xZ�\Qi��J<�v�!.�,8��	���c�Uxx�$J"� �<��i9QH]*@. ��KQ�F7X�'8`��b��ot�(��"�>�$��F�	�b�b)��{|T��IzX�����	^��;��.X��!,%OޅFy��4V�����R�!!L��|Ia��O��ą:$�Q&OZ�X	�x��#Q��G�j�0(�r��]6��(j���y��+g6.�Z��J_D��G�yB.�  ���9D$�
SV-1!惝�y�ȃ�z9�	T��:0ژk0�%�yb�D;)i��yAT�"��t0��	��y�K��>~x�(d������x�쁫�y
� �(iw��B�b���A.Gn�l`�"O�p�dS���U�U/ĵnsN�c�"O(0x��ׯc1�p"���p�Lx'"O�1Eγ!)��Q�L�.�j-��"Oz���O/ZR٤��+:��)�"O�}��EK�1�����A�W�bp�S"Or�)��1�9�/
	S��`�*O���G�	�徐��D�dnd�'1�Q!7��.W�Ь�11S�%��'��3�lŊs�J��b��(�h��'B��bdX%~� 'Ă�:�!�'`(��C�y�"튕&�8�Ł�'y��� ��l¼R����~�;
�'W��: JJ�4	���*4�tJ�'�0Tx�ڢaZ�� �dQ*�Hp��'���Q�T�{�2�3�j��'@���A�3LnX Y�뇉d����'y��Q�F:n����DL�o�B�'���ņ���-�c������'��X ao�ʵ�Á]�ft���'�$IC��ݗ[���§o�]�� 
�'cj��S�K`q2�\;(�B�'OX);R�̂U� )2���>QO���
�'�lu�}JM����S�1
�'|�yoś���q��Lk��	�'�����'��?�!cA�]�?��A�	�'\���"c[�̪І�4?v ܹ�'W��q�%N-
>�xs�5��a�'2y���:�P��h�0`ʰ��'�-*3h/;��i�s�7u�6��'�\��v/�!`���AU�5~�y�'�.0c�ĺT��rMG,�����'�&�'a���ڡ[��^�%��y�-U.o���E�)f���Ĕ�yb�Y�89��.�� I0d�ҽ�y�h�>y���ÃV^A� ү�y���n��`*BA��za�`	M�y�@T9eAjM!����x�ઋ1�yRO&"W��R��˭4PS��'�yb�߳ckа�V��,~<t��U���y���E���8� �q��ze&�!�y�mI.�ޡ{��h����I[�ye�\L�d`K����5�yrl�" ����*ՁQ�:0���V�y��B=9xd@�mE�G��-��A��yI0na2���F	*p�vB	�yB��2'M��!&�V1Q�ʩh�����y��LN����'ʙ+`ڍ�R'U9�yb�S�{�RP�3����z�ZB�M�y�B�2[��Ht�������aH��y���4O"�%��׋8��I8a��y��r*t��ǫ2�,��ԅ�y�aI�O�8H�.ɶ"��]��W!�yrF]"g��Ź�j��F�*@�آ�y�H֔s���3ɛ+1����O��y���O[��X�jI��@�qN��y���F����/�Z���H� �yr%��V�Bi1�]��lp�A��<�y¦A�^�z�pdi�/�D:����y��)Gzvʰj��[D�� �,�y����ԸAJ	[Q��������y��RPޥ��7S��L�`�L<�y뀖xܠ-��j�35�b)���\��y��`^�@���(}.婴aT��y
� ޝ �`��;������M�vES"O�!�Qƹ)�X�k���{
(P0�"O�h��hD:N���H���2gY\���"O؁���?\h|y'�)XL�%�*OJ�Z�I�q��J���i%�	�'VF�y2h� ȵCW��Y��'[�Ɉ�C#o!L1Ў-{m�8�'$�	�L�J�����vx�8�	�'�z�z D'�}u+V"͐Ĳ�'HB�EI�<q�%9Ta�,��2�'&����l��,i�`
�n��'q�eA��*�asej��T)hu��'�t$"#��6dj�B݌w����'G����54ۧ�@	{sh���'7^:�ƍ	��<	f훉L�pc�',���HJ�v��8�e�H}�̄b�'DD�Qd�(R��5c�+�,�#�'��IѰi�:|�Ɛ���3u�M��'
^t;�Z�5H��d�_;Z��{�'��̰#EĂq�Np�$D@*U�!!�'x��j��}G�3D��{��A�'	�,��E�d�`S���*E���'|X|�0Y<�+��>rƢ�i�'v�  �ljy4dU�p�b��'��xu�[2V���@�?oZ�'4d@2�c����P���'c`�
�'��1!��6�
�`�RI��Dq
�'uj-�5j� ;5��c h׵H�b h
�'�vx��m��c��|�wcO<^�Z
�'":��o��.q�u����;4��'v*��%�	I>�%���3��u��'����`ӟInj��L;W����'��p�!��t�<A��Ʈ8���'�1Q�%��T��C-e����'��ice�(^����/�7bn��	�'%� 9R"6D���@f�J� ���'P�P�3/ˬ
�2��R1>���'�8(ɤ�''��c��Y:4�����'uxX��<j�0�Aܓ2i�t*�'�J��S��2Xi��
�L�&A2ı�'��KW�Ʌ9��YF� ��i�',�}a�/+b�F�AQ��C�l̡�'�P;��E"&���AK�4+����'� �B���DE�1aa�H21Ne8�'���)b��' ��݋0���' N)��'68����"�B��
�%SĹ �'���OĴ~|��A�'L�:�'���w(P�t���j��G'(�z�'ԨKD$�֤1b ��0t��'AP�aң�=fX��W�7	�����'	�u�p�
�Hj�� ?$� �'��ҫ�kj�9�K>s�D�@
�'�x%Kq�15�� ��eZl2
�'����ea=�l���
�'݊�S��V!dPv�B�ִ}>u��+^�9��*�g��\�2�ѻ]�L��ȓ6�vP"'%ڙPs�Hю;D-��'yʽ('
 S�<pc4U}���ȓx|(h�5] ��wl2I<��ȓ  �c��v����O�B�2l�ȓE��,m�$@B�ª	JBm��8D�0B��Ӈ,�P�1�,�f�)v()D��"ǫA�!t�٨�MżKW���%D�@���)����+d���RJ#D�� �ؙ��E����塆&l��P�u"O�������$(�!��[n !�a"ODE�+2kf�� �V�m~�I�0"O ��n�T;�u��¾Co��s"OT�k�F y��� �F�J[J��"O�+P��
������i.h@�q"O��ac�:~JtP#�Is'2��"O��0jD�H�8�@�o�� #F9��"OH`�"�:"50s��.D(\�"O�)[b�:160k��U�-�� E"O�a��D��Yӕ(
����D"O����Ӥ�Ј���R�~T�5"O����$o��m�Q/ћl�&�jc"Ol9�î��H��C�#G��82�"O"h)�����*oU�O5(�T"O��E��4(B��@��C%֕��"O>8{���<tXP��Q-�`"O,MZ��1�lMB�L�T&��o�<��$S�
fr��W��y���8m�<I���/����#	,#������R�<ID���*�8���"̪2�>9��De�<�գH*L��i��w��m 0�x�<i�N�^�sk_4�`h0R��^�<�aA�� _�QQ�ɧT�<틡ǉu�<y�͚�l�DI�צ<5�}��_p�<��V��XZ$�g�~��F�LC�<a�)K�d+��_�9N���@!�e�<I6�8S�2Т�	T�S�6)p��Y�<iMN�&>j����,�@��fF�a�<��B�a^�EsP+H3tA��;,Qe�<���;Y���k �m��TC��[�<A��.��dHB(8{Ȅ��I�o�<A���WH�h�ɢ_�xi!���m�<q��
vTe��N~R�T��j�<��C�e�A7e��^F�@%�M�<�qn�V�zP�7�
�;�*s�B�I�<��@U���- c��``i��_�<�&�/͖m�FJ�ɺ�6]�<)��ݩmݮ��$�61D�\Y1ZV�<Q��S)f�X%&#۴7�F<��fDj�<��h��h����b��G�b49v�i�<a�U�:�(�ɅAW/`��ŉ�a�<�&I���d;�Q �0�"LI�<�ĕ9v�\P:�B�f�<�G�F�<q��Q!�Z ����j�0�q!NB�<�&Ct�����eO���	�|�<�ᕤWňq�X?�R�E�^y�<wm����sH˷%V5�vf�I�<a��Ps� ]���IK��w�
M�<a0c�C�P%����V9脀 J�<I���l�N�ao� Zs 5��N�<���R`=�1�t�_�f����r�M�<��	C�n�VE�.��7l���_B�<��kO&I���c  K[��S�d�<	��ڣЬ��2@R��,��V �^�<���@#�f� ��+���:�[�<!���'H���A���|�D("&#�T�<!��]�0R$0	����;"�Uz��Q�<鳧կN�>� ���:���&d�I�<9�H��L�������f�`D��'D�<��=K+ ���[��y�;T���ӤU(Wk�P����]S��?D��@�����k �`��Ah	d�x,�h���	���nx�|Z@�32|�Y�.V�VR4j֩5D�� � �AO��DT�SoF7łS"O~@�w
���	��W�p�Y�T"O�,�𯆛]F�}�f �^gX�Y"Ov�Su��dhց�-͵Z��R%"O�]*�A$��L�LQ(>�ΐ9 "O8\�4�-���hӂ��d&�rD"O>�s�)04�sA��4j�D"OF�iF��Nh20�E��#Iz%ʤ"O���!��4�|	ZC �˒�B�"OH��'�^dJ("�կU8Vr�"O�LI�� alF=�g�-;�p��"OH�A�c&-(ue�f����"O�в"^��p$��U!�"O����ˌ�E��e�T�?��Y%"O����قPD�0G�I6{��]��"O� bC��	CDH�+���p���"Ozi	�:8j�aq��0?4�c#"O���6�V�
ܢԤ+M*l��"O��0�˞. �����x�X��c"O��1da�&�f�sS`�� V�*�"Ol��5B�d�"Y��G#q
���"O�x�T'=`� �{�Q�
O�`hP"O� bF-rH�$Hٴ|K�=��"O�y��
��B �X�&���R"O�`�S������ؔ��	? �e�E"ONǇ͎pa�j��(o_|��"OR[�D�(�>�"�A�UD�X@"O��*'j\;]��E�<����"O�}�W�SXn2�+��J�~�t��"O�4�n�F�]2�+��(t\�"Odi�
 E���"�!Z��b�"O���P�_���B�ML(F$�:A"OX8���hԮ([F.T�^`&�RT"O|`�'�2R��BCֺNX���"O��D�ںX R}ӷC�yW�Y�c"O�Ⴐb�[3�q��/J��k"Op�7�*��XIb+֠�>�R"Oځ0��u�����k��%/�d� "O~�(��
l�1T�@�Ay���"O0a��Z'u:�	a�>Kw|�I6"Oz��BáwΝ��]�R4l�"O(��gڃ?!���7�< �P�Q$"O ���!u(PD��)�b"1"O���׈6�,a�H��J*	��"O�	�F6�Qɧo��\�H"Ot	"`��#����n̈́�`�3"O��rM�y�y��j���9F"OZ`��J6^H�#I�͈M��"Oh05��L�E��-޴?[@\z�"OzM�K,E�& �0o��k�6p�C"O�A�Qj��%��!Ju��=q��0YR"Oj%b��Q	� ��e�!O���"O�`-W���lR�|�f��C!��Y�	���#�OՓ���'�[ +u!��I.5[f|�`�S�������"bl!��My-��O��Z��QQ*C�>l!�N,
��a[���'l-;�]F8!�DCl��Y&(W�ʉ#��#Nd&��ȓb����&,]�)8dI����(\��1�$@�f	U��bӣ��>��Ѕ�4�� 	�c�M*���&42���S���y�L�b�j��N[,�lх�#A�5:��*��鈷�!*F4�ȓhRtM�5錫4屮����@_���S�? ��;��Y��}B#Ҥ"�ui5"O@R��J�s��D��I�/�b"O����`Y��  I.A v���"O�:�����Pb�'̳t���d"O�`E�/�� !G	`|���a"O*��P�F9�v�""F�-=c�P�%"O��Z��5!d�����~��"O��`��%��#1
�<t`��"O �۵�����G�� (0"O �B"�ٶ>߶Q��\�Vޘ��"O(�����*a!�J[{�m �"Oj��&&K r'Լ�s#Ǟ>	�W�f�<a�*~���p����¡�dO{�<)B���8��}ʘ�tB��0[B�<ɳ��Quh�qW$ل]p��Gn
[�<)�)�%${T�u'�:Y$Ѓ��T�<��(��FtA��L0{$V��$�HV�<)dD�*W0�����t�����(�T�<�0��L��:��2I~�]�W�	R�<cJ�pQ�b�GT�x�ʀom�<	�ٟ
��-(F��w��6��R�<q�K��,6��IF�hj�J�P�<��BQ�4� $Y����W�R��ōj�<��.B� �!8%@Z�R:�m���De�<Y1	ȧ*�h��
z�4��<I�! ";�(��e���p�`�x�<Y���N\��K�蘋nSݑS�C@�<�����1��$�A�W�/����$�F^�<�u�M4.�li��ǰ0�k�W�<�)v��f^�/�.y��_~��(��{�u�E��lT�{� L�v]��M0������=�8�r���E����f�<):2@���l-2��K;T�v�����M؋,�����
��=��"O�͂%X\�p��@�4$���"O�q��� ����'���`��"Od!��F�+B^�`%M�L
ٰ�'���@	M�9s��k6H)�8�p�șD��B�YZ͐���c �����0��">�%cR�Yr��a����k �=�W�(�4�;�.��yRb���؆b(l�d�%I:6�U�2�ȦZ�(m�\�"~n�-X:�I8V�M:Nu��h��� CtRC�Ɂ���M��]�Tz֢
P�B�(��V=P��	Ǔi.V��G�/Ll�1f���j��	�qd}2S��W�R<CC`˵'`�4#�-z'
t�bm�t��]���(�dOФGt^��s��	=<v"<9��׮m�2)0����	��I~��.��\��A�(J�N���NL�<I5$E�i�4lC�BI�6b���(���R��R@�$���8d+֘+�	G��'�r h�n�-~Ɉ���F��z\�	�'�r|�Pk�s:���fFWv�ѥ!׷I5��2�+ڪ(��cpm�:�F}�!�9+�]HtnL=Sb&8£��=��=�cB�$�4��#+S�3ִ�c#د��J��[AD(�G[�|������F=X�	�.��e�A,
��Y�>q�8�r�hd r�0*����6+�mq�a<��E�ҏ`"xC�^Ƹ����]� jj�s+P�	4>�a�:Z��d��F�y7�D�3�'�~RiX$gMVzv�	�D<�q/��y�HO/[�M���>-@)d��5	�U�ɴ+^.��
԰�(Y�]w�Q�Y�a��8@Rm� ��DcH�b#4lO����`	#�l���Ӫa㖏�	^��Tj�'�-[%��مh .yx��$..�&���N�(3�	8 �Y�}�Oi�cO�T8�A� ��Y#�� �0��K$_#@ۀ�_�"�1��A.�y(�����rQmɱ
�H��}Ҩd �WU�����d:`Ћ��O�d�Þ���p�E�L#b�$��Q"O���˂o)�}��d�5g����Y�> ���5e�8�L�F}
� �$pG �?.�a+���qo6�Q!�'�DK��D�����H����O�d� �#�DDI���Qj�6c:�|��"܇^�m�/�Y%�l1��
��|&?��$`��k9X�L� ���)D��0���G}�! �hS�UR�ṟ<��)@�@E�N<E�Su$�Z�p_�y���x�<)�R,-�R8� &ʔxq��A��X�D\�iq�Y��o8�pyԋЉd4+��ҍ��-�.�O�t��ۃ���_#/$9WɌ�M�b�� 4�$���'oF�՛ՋK(r>��r�9�8x1��	��d�v�ZN��!
َW-!��;���"��ҧS2�!sȈ�K�!�W���Ii��O�S{2d�g(I>%!�Ğ(��u��G�.urqc�܍m�!򤗹d����ھcj\iRa읚Q�!�ʓiu(D�7nU7~i�4:����!�$A$.#\��ǝ>[����^�!�D	�<�D�{��.@"�u(́h[!��(I����`�d��5Iկ�3!�DF�b�=���m�\��� �D!�$����<�b`�n���p
�9!�Ċi�*��JK	�ycqM�R�!�	�!�Tq���+�*��d��,!�ϟ�mDZC��~�:�����t�!���&ˆ!UA��Xl#t�	��!���������s���,	.!��K��╅�5OfB��a�F[!�$G!L�x�1U�Q{Sĝ0cɁ=�!�d��_A���V/�
��MB��88~!��8�x]������ �T�+{!�$
&<]T��>Mb��2�*ߋCb!�BFc`��^�aCz츐꛰}c!�D��4��q��EK�+�����*\)w�!��	�4�:Wm��T�"��6@�(�!�dע�t���M�_x�x���j�!�$E�n��,0�KYm�6	�ȑX�!�dm�ޭ��nU�l�t���+J�!� }�`ݨ��ߺ,3��@'��2u�!�D֎>@DX�hֳ3%^��,>m�!�]�&���Y��� ���,Ǔ{�!��=��@]4h�$8p�F)5�!��|n ��cE�����a�^��P�ȓ(�ΩPw�H�7�V��5��&#A���ȓC�(%BP���" "|T��J�-���V�s��+wgޗ:|�=��f<�#挎(GVI���K�\�q��2��X��8K��AD�&4g�Ȅ�:)\�Rs��fo|p����%/T�ȓx�@����84�p	$�/����l!p����Y�p�"�N�\����ȓ}�Jq��eN�YX�-�wI�4uC  �ȓQ�&!�u�Zx��UΔ�
KT5��K&�Qt.F/eS��B�M�9I�I��^mn�xw��<=4&A��4q�e�ȓW�X�B�;6)~��AH�2��0�ȓ\m�Uc���9�pr�̇p��i�ȓe?���T�Ҋy�6<�#��2C��Մ�r��H�\�)oXLR�U�LG������u����I�]��M��!/��ȓb�����Hs쒔"E�@�%D�dZ���0j�x����	`N���/$D� �mD�x�`����P�-�`���D D�B�'̽�����D$��if�!D���ݓ]�i�����g.<��.D�� ^E��"-"�j��$� �"O
p*�)>w��r��rP-�"O��Pc���:#�T+��%٦�F��٩1&@��pAX�i"<O.,��/��d�e��+ �氱�"O):���8\��q
��=D��53"O��z�+��D�	��,B�"O>�[N�����(ǒ����"OX�SfB;X���uE-mGL� E"O���"MK�L?r)00n:G�0�"O��p�ڃZLh�凙�ez���"OB\	C(I:b�X8�f�'bx�9@�"O�-Jv��2���뒃ؼV��1��"O���ŵ`�F(�bмhh] 4"O��k�h͘�؂�S xO�l��"OV����%^�(�Pm�M����"OX�"(Ԗ>���C��2$մ�	a*OX|
�AD%Y
S��Q�f&V��'�V���H�6��@���X��I�'$�����(M5�tR�G��$M4!h�'��Y�jɌa(i���?
�V��'�dXLB/��`� �ؽ���;�'&���@U9x����^M80k�'9���樔a	
vJ��x�n5�
�'�耢�&�;����UNZc$X�	�'{�D2�zyYO��+�`�	�'��l�h�!�D@(7ɲ� ���'�4Q��O�6�.�!N�˲ 8�',�ܣr�����3��J6A��R�'��DO��rIH��Mu��E��'�й��4�x�{Q�X#����'�|����_/z��ɲ��	�P��'z���b]<��i�ӒH�(��'3j�Z'��T��d��KR;#~QQ�'�TY���Q ��efM
/.����'V2D8�K��<��(�d/ݗ!�~L3�'�aC�)m��{�늀q�`���'ޤ`1�K�4���V�׸_t0�H�'�$�I�K	)Bb��V[�"1��c�' &Ya4WkuP����<��
�'nT��щ�YF2�q�H�9�p��
�'�]�uʛ+c����Γ��D\�
�'�&�23	��w[
a�@B�f�P��
�'����m���Q�+W�dȉ	�'lVe��F�80H�ɧM�x�")K
�'Ў���C�7�.!F�ЉB�J�S
�'��D��ߦ�Z��Y*4���
�'�B���D;�%p5��4����	�'�Q9��M�:e�5"%�]�`��x
�'¢	�c*�0Ox��c�i�p�X	�'-�����e�'M��	w<��'�H��"bܼpÚ�R� R�	����'���D��2s8Y��j�}F�80�'�b��)bબa�݂^���
�'w%�ph9*�T��K�XÀ}Y�'O��ET2)e�)�+@8&����'/j@��	HT�� �㋘t�����'�p�T�Ϸ3H���`�\7vdA	�'�\��ᜆmB���P�u|4$
�'���&N�>��!���U�ql�y��'�d����@�Q�	�d���'��P���=�>�״�3a���y���n�z��!b��j�T�����y�*�J�\�3CI^�s� HAՉ���y��V�q�|h�ƀ�q��H��hM��y
� �P#�f۩Yqֱ10�؄�d)�"OHL3p��K�Hk���zz�,�"O�ɓ��Kj�r}�v/�,n�<�D"O8����+o���W.D�MVT�`"OjE���R'j��:nM�
dD� c"OTҤ)�	�̅B�&�5cڥY"O`��&���:��rfМXj �H$"OH�pD�$Kv�gK'[ 8aF"OT8���DS9���_uE��q "Oh0�� �b��WDT�N%B�("Ot�蟛+/ܨBƃ��a��"O��B�l޴��D�w��1K��0�w"O�hG��M�pCg���1"O��;���To����I��Phv"OZdH�,^���Q��ɰ�Q"Oba�vF�Nz>,HG@�3�.�y�"OF5���Y�?��q!ϋS*�A"O~9��+�V\E�>#n��0"O.e���4�����e�+��س�"Ǫ�we;�NA1���.��(d"O��HCDTW���Ԏ	*��Q�"O��*fDǐI����҉D�MjA"Oh���i	�n�sQ����J"O�`$��<-:�hx�,�����V"O�!b�\/�,,Ac̍ ���"O6P�A�/4����$_R]�2"O6dr���x�`8�7�ĝn�:I�6"Oĉ#�ł)�1���F
aں�@�"O�)���H�L)QC���F8�"O<����4s�< �q�Ť���"O�$�G�.�Z(�ȋ/7x��"O�����B� Qp�j�0'�,�"OPU{��Ӷt@$��H�%\{�"O*e��ʯS��=l�9B�"OT��Q&�5>�	���E�om����"O��F�ڻh���@�ܨ	[V�#�"O�:�'�		����uG�q/N�a"O�(җ�Sl���� ;�M"ON�R�k��0�~�8����h��"O��S�J)�l�JWC'a�\�8"O��o�.>���*��H�%��xI�"OR墦�)7׆�0� ѥ3�$t�"O����´5�PQcuA�K�i�"O�ѕh[Qkb�ץv����"OJ�酦��Op5K$��.:h�bt"OJ�@�/�?p����6ʘ6$��[�"O�IX?L��<IDo�Y��{dO�Z�<�tC���B�͉j%�f)Z�<�Ư�@���+֕X�~E���GU�<��.q(�)'CG`�,I��U�<�����/7�Hv�(N��=�'��R�<a����P���ص���bPW��v�<��/Z9�*,�v�������1��x�<���>���PEy�F�y�<�f�Syd���9�z�y��t�<�㊜�}��ġ���ze��Q�m�<Q���\s��J0�B�H{�p1!JYl�<�E-ʞT�b�S�V/�& �	H}�<���#"�0�Bb흊�T��@d�<�lB�c�vH �A�(��X��'f�<@�V�#I����Ѕn�ZT���a���=iv�ë0��8�M��pI	�j�Z�<�"�	Q�j�ѥB�-B۰q8�	OS�<ف�͗B�ҡ���Ѩd�e��\I�<� ��򮜊��1�0����"Ov]q%C���`��ʉ|��� �"O~�$$�h����p`F����""O.���晳�l�����tQg"O�dڕ�A�+��̫�C��:�CA"O��I1/��G� �z�)�"x�6(��"OJl�r�E	On��$腃 ����5"O ��k8;�ub%GW08�F�:5"O^1�����Ўt���$颬�"O ��1�� g�R��eD�65��ɖ"O�)a�R����³dP� ���t"O���E,�Nl#�Z1 "O0�g���t��_i��9��p�<1����h|a��Y0�����n�<���F`�恙���;	��us���B�<yah� 	s�J#�/6��]�f�CE�<��&�{I�Q�U�K��Mk�"�V�<��T�r�Ԩe\A�����KP�<�c��k�nJ�`�ڌ �N�<�p�B�"�dt"քǝ`zeX5�SH�<i�vj�چ�CB�(�A���i�<a�A��*|�}(�
%�h�C��f�<Yw�֧0�r5"�,G~ �B�~�<ن��3����"�r�3m�y�<b�J��a�Qb]�KRh��.l�<����+M�"HR ޯ�,���	c�<�e��0���S���PD`�2ծ�\�<!�@ԍ�RlS���tX�Q�+n�<��C��bդ�
��������m�<�R?uX<A�Po��4�I����k�<ن/��]L�H�`�.\k�%��V_�<ɇd����� ,[�"��$�Z�<A���1\��B'.��t����A�n�<1�Kيo���0�cAY�B��Og�<��dN�kh�;jP�R���&.�{�<�Sg�zZr����B���w�Fv�<���4i�3�K��'�e���Q\�<q�J��y���hA��(�XR��[�<�0Ď9Gd�;�C]����S��|�<q��2"�`��i�Q j��ԩPO�<�E�G9 ��@c�Gi���¥�O�<����30ZD�GX���@b��OR�<�5��^���1'�P��F�Q�"��ȓz*��¨�&]b� bn_�{|�a�ȓG�Լ���8��� ����)���I�y��ۼN���)����x��u��29����m�+�2TYWk�)K$�ȓu��u�
Y�8T04m�06�ȓw�y�c_��i�¡��.X�!��tQB0�7��w�>x�	+l6�!��B����d+"�B)�@O%4�����L�ۖ��;t6�
U�ȓD����w�ы7�z`�%��4b�`�ȓXJ�r%*EW%�-���*�]��H+�L� ��&-CBY ��W(#ц��LăG�Oo���1ЇZ"Vu��ȓR��������4G�S���\��ȓ0'N�r��� �(ٔ' �H���.P��`1�N�n6�=#� M*J�n����q Bk�	�
��ЀR�l�L�ȓ4�݋�_"5q�T�B�H�FL�� ����C�n��90D�]��ȓS�N� ÿ�r-���"a�M{�"O�s%`Q/hLӐխY���"O� ��BS&�Q����#?@Q�5"Ob ���?b��G�@5[����"O�Ӥ(�S����O Q���&"O��u�@�rW�@��Dܷ~%@���"O�5�\�,�T�����1�]�F"O��jWc��$DH6C�*u��"OR��!Q�	&�	�N�"a+A"O��@��Z�C��!��N&N�9�"O�*��P�N� f�؜K~NAKP"O �D��\���PՕwl�]+E"O��K��	R.��`oR^&)��"O���!.R�O�E�Հ{�����"Od�A�h� E�`
!n�	4$���"Oʠ������"S��*a�`V"OvE���@�{;J9vV�"��X�"O�)H�H���X�K��H���;�"O8�q�E�Ur<��I�,d��k�"O^�@۶y�.A��o�3|�> �"O�YT��.2������9�����"O�e����X��(�à�S�D�C�"Ovpr���)�*
oP3�LE��"Oj��r�[Z���T.�G�j��s"O<E��^F���
G�M+gnV-��"Od�)�HWr� +�OI4f��j3"O�c.�q�4ib0��[��7�1D���c/��[(�Xi�Ι�CVB�c1D��z&I
�5���2�*Iu�UB�K-D�4�fz)A���
b ��M�5�!�DV�b�n�"�(?@�Ѕ��,�J�!��Z w��a�@��&��ezqJ'6!�Q����7 �p嘕ʑ�a�!�DV�S\9j݁n�\���If�!�$R�^S�TS�E�%htmY��ܽI)!�dǂ��@A���Q�B�:�F�+6�!��=ӰK�@� l�6%ɺ6�!�d�*�|(Q�$�����WY��!��ٙ@��p'(�9���P�匕n!��V!�]��ْ(�4	jd-V�!����!�*шx�E#$E<�!�dM�d�
�b3��rP��JҤq�!�	x��۰j*<E����Ȍ;p�!��4 �N�;�l׮e��q��� x�!��ٓ�T�(&㛆(*���	>!�A�aS��U����)�G^^Q!��h�D����JB��
5���^b!�d��#�R��$�H�7aP-	�R!A$!��^�n���4�Jf�1:���<'�!�$�=�v�Ic�'Vlt�*��~!��2+F�=���k�-�4��Wu!�$��)�=3rJ]t?d��L�-�!��4c��`B��q@*h��S5vX!��6_Y�������1��/uA!�Rhv%(�oC:o R��u!���f�&3�͓�s⚙8E$�x�!��ȃs��X;@�Y�/͘���_�	�!�䗏1ڌ	d/L
O���8�f��G�!�$I ښ5K�H��Z,��'L��!�ą �$��d�
~d�m�����!�$_%X�)C�B-Ny��ϔ�{�!�d��U�p�ݡL^�5�VNCl�!��A�&�,�dAJ	M1XYZW&X0�!�ВOXp�zEc�M L�IucM<Qb!�DB=c.�T��H Xn�Q񦡟;0e!�D>l��H d�>9b��4�E�1I!�� ̔۠�E+@^��@1i�R��Ht"O�%a�b�%[}�W��wv) "O q ��թ`�� �U�'T^d�h�"O�]if�W�N��4b�8vz��v"O�hH�� 
���'�K�m_�=Y�"O��vnӝgZO
y�5f��,!�䚀g>͓V�]�#=�y׎F�Z !�$1g��i�66x��h��!�$��s'�}	!�R�D� %"�9<!�D�<Q�\Y��M��^��c�D�i�!�$�9��8�2fƀgQ���`��!�9	`~ՉE�ҌmI��%�ǯx�!�D<x�$-����j-YP�ڂ�!�DƟ}wԉ�ƥ�� ��uJ��-�!�DPcGrq���R%#���W�O�!�䘃b)bĨr@�{�fH�$M;M�!�F5�Lآ��"C�F�qv��jL!��^1Db<�[0�ĺ@u��Q��HI!�d&M-��`A׳$�t���H�%�!�5 ;���̚��:�6'�K�!�Dڧ~���1��l)�֌��Is!��]�����M�p��f+�	 X!�D��0�R7�[�d��!�sD�7|;!�D��7��xC�m~6���� <�!�Ę�|S~	���y`ɩ�ʇ�!���Bąp�e��p�&J%�!�D�b� u #צua<�����+l!�� M���E�L�W��-�S� z
�'<�t��`Q/\������ E�HB�'�F�#��P�!��]��옰D��P�
�'7���V�G*V�)�䗱HP���'�� ��VbƍA7랏��	�	�'����ϛ�4�ъޣU]���'��˓`��B��"���E�^3�yR�K>2��*F[E���d��
�y�d��M2��C�%:�5q���y��|�*�3����ʙ�����y���:��E ��<Vt��H��y2�Uk�i7�D�ȬXFަ�y¨����F.��}x��w`ō�y��W�9�Uz�%2oˬDpVѮ�yB�5u�Y�ʘ�c-i���y�ֻK��t�fA�C1���d�R��y���$b��"9^��X4W��y�nB�G`��E,h����y"�5���F�ܝ$Ց�D��yBo �1ըܹ�)��+ !�5��O�"~Z0�E�!�4���mMH��1:D�E[�<	rH$T��0�sPfb��SET�<�F�>S#��P��j�֝�"*�S�<��(\�h3�]����=�̭`��Q�<icK�>̠�p����)�Rh(DJ�b�<�@D�3�@\�g?=bB��t�<�C޿r���E bx�ЫdQY�<�VF�� em�Qc��pf9���S�<���\0/�j���8C��xy��JN�<��I7�؉	���6:x�Q1�B�<�q-O�M�`A� &Wq��l!� i�<Y���.���BȄN��99�)b�<I/I  �Fm꓂·?���#QaQB�<1���Kg�a{2c�v.����@�<��.��4����Ĥp���%O�~�<13-^cjD��8O��lFS�<!C��&��8p�*��;7��I�<� p�¦	'O0��iBh1(J�C�"O�""üi ��`���`͘�RA"O� D��N����@�ŴX]����"O�q��<5�Q�&Ÿ'B��sB"O�=��Ț=e���I	 TL�{�"OE��Ϡ;���8d@A�qM0��"Ov��H6�`�Do\�I�6Չ`"O����L"S�z����Y�I��(� "O��J�i�'��d.B�6�nt�5"O���&���&��� �#�J��$3D�`0c���T�	�M˶2^n��� /D�a�*�E�M� ʰ8�&��
,D���F5+:���C���a<i��&D��pB^1J�x�q��/P��=���(D�$P�)S#��P�1N�:/��˰�#D����N�|��h�  	wE���E"D�{���-V|@/�Mx(���?D��adDҴ
�^c��S���T`=D�����	)I����]�j4�M�j-D�Ա���7bt���F��[�xcċ)D��b�,��0���UJ.@vԊ'3D��	!A��W��p��n̨F� �rfa0D��x@��x�ܴ�� &�����e)D��@Eȕ�9n^����ï� �p�<D��:%�6Q���7���lO���`?D�h�T��.>#�� L��*	�����)D��V*�	�2�۴S�"��0lZP�<�&�u��(������a& g
!�$U�N�`��k�6E���`��t�!���s����M�i���dԢ�!��X߾}��N+��8�ƅ�v�!�6c�l���D�%�v=i�eZ�S�!�DΊSU2��A�>pۚMk�EP��!��h<��X��q�V$��^&t!��'�ZP�X/'OB!E�];Ig!��
}p^�*Ɨ#	gx���ر?X!��[�F��0�A�^�EV��P��W0!�Ǵh���q��P�HQE^�yE!�	�4�Hr��eSP�qw� E@!�D�����c�Q%H9��Ή�H>!�D�#����j�9h�	�6	!��Ŗ+�@!��N�";U*8��iN!�dǹD�H0����:L*�K���!��Vt]ɴg��*P�5a��!�$��&��Q�nX� �L�ʂ�ѝf�!�D�Pv0��� V�R�.������w�!��G,���Y0JV�S`�x�T.�,Fk!�D-mHL<:�C��u<0�ڗOÞ8!�$K�t��-�� 	@*:�a��N"�!���8w@>�������y0�ԛ^K!�^��}���ܓbx���C�a�!�FY��ɘ���*)`�pGW�b!�D�0p��ʴWE�%�t�^�YO!�������Ǒ$D8� i$�E=IH!�$CW� �po�8ҝ���	*]\!��i1������HhŲ�pt"O���nO'#���`��B�F�c"O�l2$DP��/̥W�0	30"O�EYr�ҏ~mR�1r+��Mu�`��"O�*�M,p������-a����"O��;�(׎2�C��I�?����"O�(:��:R��i@�U�0����@"OPu�b,̬��@��*{.1��"O\�� �s*�S��
�8	"O� 4�!��ފ^�D(�%̜��h%h�"OJ��$���q��,�Մ� �B$r%"O$�j�)T#m�t�8'M�f�@Q"O���v��3=��9A�Z�x�D�"O]	�c��	�����o�*�Z�"ON� g�
�8 +�$�q��Q
"OViRAI@^,�p�4-�ya�"ONt ���> �|�V�[�)8�"O�]��@�"LP*0�aCW�I���Q�"O$A�����d��A�)�t�["O����a�_��}��+m�T�ᑆ�O��e�\��Mc�O?��<F��	"�1A��)�P�j���k���FL2�h�U)݋��¡r���>Q���@�(p�8���͖y~D�`�iM���e��l����$��H8�ʋPvpH8��R~�s��(���9\����L�%[ՒI�wӒ�;��'�"jz�V��-�禵r�.}!��z�"D,7��$��ȶ����͟d��	�9�ȥ�Ô�q��S�.µ05�<��iU�7M?��ܺc�K���W,[-���w��)v�', �ˡ��?	b�'���'���]���l�	1h��%E�c��(C���d.��[czz��v���J��%D�����a�Q�`�'�샖�M�"�=��9&�!1v�#h�t��,[�h���`"�JV�U�X\	�#�)�Z�+�'�9c2̒
gY�(P��/I���H$��O<�x���O~qn>���<��'���D�
5�mz� �	#l�j���!��Ģx�lu�A��@� ���8SmL�1޴(!�v�|��O�t^������|�^<S�Շr^�1��b٫Rw@4z��Esx�4��+r�4��H�Gv�;�n�!X�����$�b
	�.#h�ڍ����$x%��$� N3DY��J4�_�=�}(��!���H���B��=�ڴ���
C�$�HEy�n�'��%�H�	�WP��B�
 ������� U��=�񌁱�M{�����Ŧ��?ydџD@��/Ŕ�5 C�-/@�ٙv"O�a�bv6�ӧ��/M&~0)��O��oګ�M.O��aºޛ��'�BW?iP-A"*�x�r�F}A:���-���%���?��u�����hS�<��1�� �] �L"Ժ��D�K�L����ᮞ�|>�I9�.��Q�d)sHƀ\�n,��FMT�H�)]�3�vDѧ�դ,���{��A� 52P�T�-��kqnԧ`�
D��O�dAg�':7������1	у�9k�����(�5<��ـ���?a����'�(9j���t��-�T
څo�k
�4�v�'����|4�@�*^E'$�)f#� �~��΍`��6�O<��|�0`Ή�?9��Mkq��O 83�����g�6p���th��"l�1`,|h��B�Ó'����'��Yc�}
���"�^�Xp��-5��̐ߴg�P8ǣ�*+P-�����*�n�c'/	wo���RF����Ba����-i�"|���UY#׽iR:8���:m���M����~�s�<]b���xـ@���H�v9I�OH��"���'����ŗ!G�@ݐ���\Iv�K��$V���4�?��i�"��^I���Mqd%Pj�͠�)Կa^��I���d�aiB�������	˟��_w�r�i (�#"D�%܌u�o�9IBf���d_""6��2k4߶���Jo *�i���N��|�˄/������"=bqP�GA$Ap6m�):f�C��" ���A�p�ăʌH�nt�G�Q7���Q�~����a�1S\1�(�e��.0���		�MC� �~�'�[��[���/A޼����u_\a2Dc���x��#�Uң����<"�.G�M�4-���|�^>Y�>�i7 >  ��PDxªM�c�= �%G'($
U8�C�0>!U�ҹ,ײY!Ӫ@<p+���a�3;�MR�gT�U�Ќ�T��QN�y0�'x���	Π
�b0���7B�h���-�s�
�%�:�#�A�k��re	�GP�\ҥc4J���y"/XW�V�i�"O a��7���U�b���;� J�P��d �4���i�g��W�A�`�5	�1���>J|g��{0 �7�
|�!��V�@��9+�-GtE�fg�(z��HD�����tHN4�V��;��8)�	-I�1OT `�k�fg�@0��݉1�A�&�'nN�z3�M���A�:[� B�� ��!A�.��`6�
 P8�A� �0=�S�Ј|��I`る�>80��C{�'FZxj��Ƒq9��:���5w��]0ଔ�rr�=Z��ۻc X`��kّ���IcL���y��¹N��!�?���{sM�]h,��B%��{º��e��WtИ�ûJ�(����w~�K7★(���ŋɰ22�A�'�4Q��J�A#"�i�_�M�t�E�]$T�Y�.[�Rp��2@����B�㢥j�y2�&*�l� bT���3rA�0>��叱k��a�fO�aƎB�Z!<�CEb׉אi����8���B?P,f���ɏ>�tKS��:2����@"#<I���_�4�3����*N~�a�N��$�^�_0��#b%Iu̓[8��c���)_�=��vI�<H�`�ߏk��D�'��Wd���L<&1���s����O�5Qv�c���'t���Ƭ����'��+���2c��S$Q
TBۋy�����lWߟ|2�I� ������-/��F���,�8��J�:&����Oם:����!�*,OLQyae��{�d�ѣ>ti1 �3^Q�6M!eU���k1��<�he9��x��	~���l�̌� K��Oda+5�c���W�9YX`���@BEH^!����6���������>�|��ʑq��!����=�=�UkVA��� 	��n��/O?�I��!Cp)ɒp0���U�zGJ�k�}�ߓ���I�P�0DP��L�~�*�� ^S�I$:ʅ��?�
���!���N�e$(8K�㙒X~��Q���.��<q���e1�5{�OV���q$A�*x��oX >��� 4ثO<� t�:㌒+Lj����>s5�!1!�	2S�t�8焂K�O�8p��"��Ds������y򠑭��b�b>�Dˁ�,��G
�_;N����'D���'�Н]ͶPr��\�d<���-��'G��1�𙟸�������rE��6+N`j�4D��KE��`in�P�� �8'.P8�钽P\X<A���XW�Ҟf��t:�B��&t���I�{T*=(I<��J��M�5J�&C���IBY�<9�F�|�x�� �bI��a�X�<a��P�U��	��(, ����P�<��8i�$)���ѻfh�dB�	�	K��С��6�*��d�VB�	��&@2��=|�	�2��f^<B䉯��i��H
R���'ғ,���D��@�t�q*Gb�.q��f!�"O����R�&Ɠ�Es��3�"O�xx����oژi#��X9G~$� "Oz�E�#<��}·�r�]B$"O`x� �0/u�y �$Օ:@"�8�"O����:{����bQ,�*���"O�!����#@(�AŁ�Vg�YKg"O��f�Y/M���A.��hM`��"O��P�1+��=�D�Kۜ�(�"O���ȘV�1���o��	�"O ����ϙs�V�c'�ԕ"�*h�%���
GN�k��|�\�^K��ӄԨ���q��(�O����Od<�qK�?nh:��#o��"OLM����7�Z��U��{�N����9�!F���=~C�Ũ�S�f���ƕ��0=��^�^�#cJG�<Qw�ο@��肤�/���c��<��DK������,S��^�9�h�A�gߒZ�n�H�dސ^�~��K�01�?防W��"�x��@.�����)6?Qq,����=$���~���yu����R�q
�?E������__~r�����	 8���Ӳ$�y�b�@1݅=C�ɐQ��q���|I4! �#R�-Y�A�c���D"�O��H�[w<z����
!�`t�W�'�F��
��e8���'l���(�u�\�;�j�X����'�=l���S���Ӈ�3 �蒌y�1$��҄oہ���:�B�H�.L&��ROIe<x�0"O�Q� ]5,�N�?r3N�t����S������1�g~�"Fa�4��ˇ$r��P�@C��y	�O����#N�WS�H��x(˄˥s�nm��'�i�`
��O�@S2`�`�#x��:2�!LO d����;^F=�U0Oxy�6��,	�b�"�.�<U�\B"O�}�U�==��� �@�16D��A�5>T�B��ٕX]?�k���0Z�ۆ�"�"R��?D���S�P���\ 1��>tx�<��^8M��`n-?9�-����F��ڽ��f�;N��s���W�zdۑ�܉k`a~bjťy�tā�L��!��p�F|�GOF<äЁ��4�<�{��0c����}k3+�� k@l��?D�0FB�=3�!E� $��a��>�	  ��!u�?�"8 +�ZP��(�v��0"Oxl�#'�YQz���:��|��Ƥ>z1O�\[�3?�QkЦW�z���F g�=q���K�<� F�L�� ѵ@7&���Y��p��(
P��|3&_*p���KB�d=X�J�	"LO�C���$��-���acX)J�f��� �&B�I�R�V�)���w�>E�mF:���?�Bڎp���<�}���1@x9�g�J�� RN>D�K�Z&ad����3 ��4�����@��c��p�'�g~Rᙍ�H3f�# **8a��yRb�_�L�	c�4&�ᡇ�v-��5���0?1���t^B	���@�zۀ�k��~��H1� G�i�������fΛm�0����C60=���S�? n@s�B��k48���^�sX�*�"O��G��
�X�cT���5�
�q�"OP�j�?�V=����=r��"O��Pk\�2� �YD�[*_NU�B�q����'\��ꂅ1�3�R#>�@�W��i��"PǞ-�!��*FD�D
3P��M3��S���"��K�4�[P�'� �2!�/WŠ4��^�A	�Z��a)+>�>t�'��`�+ �i��iu#
J9<�I�'��0�$+דm"��d�^�2tЊL<9S�U�@m(���iU�O�0QB-ʅ������VL(h�'vr��3 ��u���B�-
',�L���'V>��JPĹ0���xS[��# �V�pJ� �.G��x��W0��0�'i��c~��`F@�Y��$���!}��z�2m�U�G��>{��u�P"��I�y�����$<
�"�*�5H\1n,rl#GF�m��ȓ��(+3f��y;��I�oѻn7��%�XS�ޠs�~<K�#2�$E�YPs_�b�jeف���`Ԓ��ȓ7:
`�CC�x������^��ą�0���Y�H��=�L8�Ǘ/�d��ȓF3�8
��g���J#ْX���ȓ���઀�f�@�Ā��W�Ƙ�ȓ?+�<Q2,ܡMv�M�5�� |>��ȓ=�&q 򨉺݀%㣋޻�4ɇȓbπ1���]ސ�҃�H�Pćȓ	� ��M�4w���k'�9B^��ȓ>��L�e��fB�6`dq�5�ȓ�(�:UAֲ.���2�<V��ȓi�Q����~�p����r� �ȓ5%��� �Q�4[& �2�J���>����Ci��VM���AO_���X�ȓQ}.D��G�c\�2#��Bx���ȓX/��/5C�$���UO�dh�ģ&D�����Ɔ6W�<�dB��$��2�)D��т�_)d��7�6)el{��&D�����)&��٢B)<,8"U�%D���"�X,)�((���-)���#�"D���#k���1;�@H�x�l1�f D�L)��.}��j�E
&l$UHԫ=D�Ce!#.Z�#���ɑ�I:D���GK�f� ��S�]�4l��	�,D�(��i��[e$a��o`��`�5,+D�TA�J_R���"�\�6����b)D��*V��i�d`I��Y���D�܆�yR]� ~�ӀK�Q�^D�F���y2����8���^�Q�ڕ�B��y�5'F4�(��=����D�
�yb��%(��Q*P�/�>�qCL��y2-�3�Z�����'�B��%�_��yrj�9Q��0G*ϼÄ�j�㏋�y��
f�Ҩbp�ջsHL򃏘��y�(�(y+րp�e-*�h�
� �y"E 8�Tb�ռo��m�
�
�yrAJ�+vX����a-
1�E��y��#�����d�Wd��ť�y��*(�8:6C
9E�h�$��y���\-���ԈX�'����@W��yR��� N�����\����z/ �yB��B��<��cJ'M@��q�
��y���Y�����>U��t��;�ybj��N��q���ĔG�"x(`& ��yb��0��pk�A8>H�y���&�y��-H� 9Q�n�C�q eC��y�=A�������j�X� ��ybD �mJd�H��Y�W���a@D*�y
� ���Ѥʀ
�q3E�	{�{�"O^��N�?vGt�Sa'4}D\�W"ObUyV�@�RKv��Vȑ�
$�)2"OLr�'�9��̋���z���0&"Od��O�jf�BO�+lJ�"O�Qbd�������.b�2%"OΨ�WNO>*'�,T�9v�����"O��3��D8� ��$.	q0�B�"Ol��ǀ43�e�4c0H �"O��B�^2d�U��\�f�~�X4"O8�
�G��Z���T�U�T`8q"O�`�Ѫ�V����e+B�{eйY�"O� ��d��)Ĝ��3醍W+�5�U"O�P� �[�xI�d�˧,*��ذ"O�1(�d�B T�x#�Q�R!�YF"OK���Wy ܣg�)336(Ҧ"Ou�bi��:�D�M.���"O\�t&�X{�� ��5+^��Q"O��	B, J���,g,8�'"O*�`�eG�J��}�d�,�d�C�"O��s�iR#,`X�ZF�Is����'"O�來�TOB��
I�Ѭ��g!�],v���������̍Q�!�@1>qM��I�[����FjO�q0!�M?;���{�O<q�T�	��!�M�X H��ԉ�0f�ƀ!6��*�!��ݚv�@�p���%�zAaԦ��<�!�dĄ�����Jw-�� ��éx!���2�:et��&H�ԡD��1�!��X2��o^)L�,hH��2!�J� �x�Z�5Ѐ)iG�1'!�DB�}�H�� Ƈ4�pU{͛
!�D�ch�k� Y�S��{0�/�!�Ā�	g$���g�.��-��Q#!�$)=R,aP�-̀P������!���1���r���l�HiQ���!�$��R��%y�ʍ,-���*Gk�>$�!�dA;�2�QS���l9У�M�z�!�d�	��Q�c�8݈�P'�Q��!򄐌6���'eT5'2t��혜^�!�$Z�/��9�G��ZsReӑm֑F0!�B��\���蚦)Z�d��ŕ&3!�d��%���)a !��U��Ŏ2J!�d�A�<YK��-�f�fG��T�!�	 ^�0#B[��9"5$�/|X!�䙊B�f1��j��]}%�fA�I!�F. �@0cT v�у�A�[/!��N�r�A b�i�8��l݆-!�d�(xu�׮Ov���-X�!�J�?��]*��\�r�gT!Ux!�$Բ|���`�=w�<,(�e�*�!���Tꆍ�TC��n��� e=\!򤘿G�ŋ��_�VK�x� o��O!�_6���ꄊ��U:���c.F�
�!򄏫"1�B!�/r�<=��,��4X!� H�P��Ah�pn���K�&nW!�D�@ 怪�wXhZFT]k!��	K��1Qwaȫp�� B�67N!���Msp�S6U�����*~�!�ĉ�H_��`c��%�N%�R��=4�!���Tl�y`�B�}�.a��}!��#�@�����x��lh���B`!��S:QWba�����McU�=hK!�"`��[��7X�HA�W��'>!�� ܭ1��Z#AV@@
�9C$��g"O.x��̓/;A�
�HA>y,,p�"O���� jI���ӜV]��"O�D��cS'8d4����ݻ53��D"O(!�O�7-�C�C'y+\�ْ"O*��
XM��M���X8p�#�"O�}�%�FLiv �w�;���"OV%�B��	QA+#���{&mP"Ov ��ִp p�M6'�会7"O��sff�jP�����1c��"O����P�>w����-��Jh�!�"OF���֦+߬��7��1 9ry8�"OZ���I�t�.Ua�,ʵs�4��0"O����䛍G0\����/@.F�#�"O�Ɋ��X.Tb�}��e�X�x� F"OX��Ċ�t|n�Q��%)ϮY7�'Oў ��h��eF�CQ�N;\Lv�h�J4D���K��<�H!B�R��DI[G	1D��*0 +{Ԇ�{�%Oi��y�@*D�<Qk;(�<��%�5����B/-��p<y iKv4M���K!y�80�&\W�<YF�=��pA�	�c>X@�V��H�<�q��j��C٣����+[`�<Y�������!֣O���G/u�<�U�R���+	�qC��¤�Rw�<A�Ί+
�$%��̄�8qZ��t�<��[�����zn>�+��u�<��F!%�Ҍ�w�M�D`����y�<97c�$�2�ja�;Ev��CI�|�<�b�G�rM �� b.�ⵘe��z�<Q��1^>V����Z�VC`�8�Ɣ]�<a�k�U��y�>=D�S��	B�'7ў�'Wʖ���%8��ˡ
�<o|���ȓC�>�S��X.4l񄅻T~Э��;���y�I�<��ā�.iŅ�Ic�%5�(�%G�-{��3�I�(3��E��R�1��޸�l��b�I�L>���ȓ0V��ړNH�e�����W0>	��-�0��ΎQjK�lZ�/	(��'������" Q�x{�͂��\��L����LQ� ��m���5:�X��ȓ�&m�nSQ:N���AB�i���ȓa@ب ���}�V�1�U5.��A��($0�C��ͤ_�Da���d$���j�r�82��|�4tp&ӣb����8"Ds���u�)�(������&��8A+�.q�b���͚N�lM�ȓi|�y��^���"`і:"��ȓ����KJ'_j��p����5���u�������'tЄ�M����$�ڸ	�^1-��5@�g�1����q�����M��W/�)o�q��z��"E�T.]��G�(�
�ȓq*�eH͏7xD�s�� ^Q��ȓ[�8Mi"�3){��SV�;C<���+�����8tr�	�clO˂#�[��hO1��Q��o4pur��ŤN��� �"OT�A���l6*���h�,��a"O6M3�kޢ]�*� 1G��X\�"O$�p�(k�"�¤�8���!p"OB�T�ح�క�+�P�	R"O�(�#n�1;�T��Jݛ>�6���"Ob�i"m�8��s�E�p"O��#S7\� �L!�6I)�"O� 8Y�6�Űh�֌r�%W)4�¶"O�e�"U&������^1;�$��"O�0"�,���x��M� b�P�S$"O&yBU'�/eP�8�˛�M}<5s�"Oti�̐	vs�\�d��/�x��"O�%s�Z?u�&�qedˁ5��Q�"O�b�^�MÏ�X���"Oz�t�LG�@e ��]�(+��2@"O*QK�h�_���;� Ӽ)&�q"OR���7 �]�ab�1dh\�"O@� N��.����M�,8�"On��B�37\���#�<{����"O��
Um]�j���!�����Br"O�h�l���6K�T;�!��"On�K��^ 9��� 4��/���0"OzW��5!3j�	���1#\�3"O&͚ �P=$�%i�mL�Hڭy�"O��0D��- ����	��ȁ"OFĹ���rK�LP@K��f�u "O��xPK�+X�F�T�C10�5�"O ԫ�>lԩA�̎Kv	
�"O��ȁٓ&�j0�b��
#; =��"O�}��%�)���)��O� x�@�"O��%�W�D����$��(�	���'o����� �Q�|8�A�!��U(�B�I$O�B	�B�z���HwFɢlJ�B�ɸd<i �f��C���jQM�1�B�	�D��m�,�p�{�%��?TlB�	�UT���Fe	%+��A��[&�6B�I�RSh�{ׁ�5P���S兜�6Q:B�	1V���gЕ2x"�!Y�j��B�	<)m��%I�6vp<�3d�+Z4�B�ɬ?�j�KC� �ib�15nC�	>Ұh�e#/5�t���>4~LC�	h�NňF�>���K��+�DC�	7L���f H�Kc�HȄ-�;pC�	�	�|�*�6E�|@�a�p�B�1]|h)w�B�*��!
�5BʰB�ɪYg� �7�pm����S����`��<����fur�E�?\ub��ȓ1z�}�Vl
=	# ��!L8h&�-�ȓ`��-�C��	%��L�t�M)5�Q�ȓd ����Y�b�j
02�Y�ȓf��Չ3n��fB����	��e�0��ȓz����)H.* ΍!S�W�i�����رj�#��>���Q5CT�ȓh1"	h�I�b' �&�ڳ%N�U�ȓfn�p!�H�r���(Wb �cL����D{��Œ!�]iD2/-�-����He	BN���Q'�ij���ȓXiN���T/z�ltS�φ�R�~��ȓE~x �K�B<x�� �W>n͸����|�Gׁ9M��j��C�`Lh�ȓO��ŲGL�*p�r�J�b Q�	������'�Ę>$��RB��G`P��� �"�@�%%@ܜ�p�H�~����ȓ58Ƹ��\�1�ƭr�&�Q���&�P�i�ibH�:��G/��I�ȓ���k�(��I�~ȡv��T���ȓB����P2�>����f_�͇ȓZ��J2#N3T4p���ͩ6�D�ȓ��h0�̛2]R*�c[�k�Є��d4�`-�0 {~i�� .1]��$cr����H=c)b��D.�m0܇�S�? *��.�Y�	��`'\�Z���"O���B�:h
,k���@D��"O*��`�\(#��j&o��@��"O&�:c��2qb5� @6�t�"OH�  L���D*GÞ/N$�5��"O
50��ʑt ���, �M��� "O�={��ZCb�Dr�,��H�̕P"O Ii��"a����Y�nDyW"OV<! ��R��樌	�&��"O��c�̀ �4T����0W����"O����`�5 � !lH�)�JQyG�8D� ��3iE���$��[:E9��5D���G��3u}��Pw��3>X.Ma5D�Hc��A�8/��q
֊Xg��4D��[�KM#I4\II�ԫ`#�e�EH0D�`���L:��0#���+G`	:�-D�l�1o޺6s����Ϙ�&�||���)D��A�&�9|�{��C&';DXpR�<D���$�"����R��<d&2T"9D��U�UđbǊ\V�U��$7D� ;s�>V���q��m�g�5D����Ҕs7�x���X+|-���3D��RE��AB�Dsa�	3H�,�W�=D�P�$���ty"���F(N��� D6D��B-�:%��P��ŽkrҴʧ7D�p郇�$@6P�5�4����+7D����j��ִ��ر^��9ӠH"D�``�"��-�r�y�$��H��-�-D�dB�/�3�6�kH*df���C>D�X���5B�p$�!F�~���=D����eɐH�]�B��Rv��<D�Գ�@�e**q bb����Q�b:D�$ ���@���+����y�Z�Z �"D�09"kԢFC�T�wg�'�\�꣮5D��a+�&x�4������[0���M4D�4ca�P�L��,c񁅚S�K2�6D���S-�'�N�����"o��\:Bn!D�$���[v��P6J%{UҰ�S�=D�
��X�E0�sD�]�`�ڶ&D��"e�J�ME�Z�-֏o�b�p��"D���f̌Z��Q�s���T�@��!D��/	?�0Q@s�\<UD�$?D��A	U<��ds�-�aVB���n*D�(��c���t�7��;]6�³c5D�����P ?��E 3��8�hI�K D���D�&R�<�f��?Y)B�[��>D�8�1i�-s�(Q�wǫyw���?D�L�"�շ~|e{���,�
�H��<D��h��0T�x�G A( ��t@�'9D�,���g�V(�f�C�W�>4iC�!D�$��/��hPR���Tn,�`I2D��*��G�-����kug:D�l3�G�O���Q�[�0Z�8�%4D�d0�b��w�9�*Ү��V#3D�l{Ԯ� E5�BC�L�4�S�I%D��1��L=��xRw�۱y�N-[��-D���$%,_�j��G{9TTr �6D���(^�;�Ƞ��ڨo�2�@�c6D��c�_�O��s)�3&���F,3D���dҭJ/PQj51Tu�
4�$D��+�̖M� !�A��'��8�.$D�X�i�<����"G^�:j�\��#0D�8x���^�h�ia*iܤ<��!D�"ҏדo&��! ܕ	�b��wf+D�� h�5�Вjqd���ζP"B*�"Ov,q��@�{�Q�d���>,y� "O��#R��Hl��FJ'$�A�"O�Y8�+Sprxhٳ��V�%V"O��{b�V^�
و�g�Ic8�"O����9Ii�A�FT�%xx���"O�|�̗�#�n}�҅M3)eD@" "Ob�Q�D�4W�0x���]^^���"Of9M2��A��/�n�V6n?D� ��GD�I��B�O$�u�� =D�Ш�W8S����̓'3`��':D�8#E`��d�k�'�W�AQ��+D�P���ߎa/P�S��;�@���6D�t[�̔��Y�F��"Uܱ0��8D������TZ���D�?3��u�q�:D��hC���D���F�K�;�Tc��>D��زDzB�#��G,rN�A��<D����(q�H[�BF�����ń:D���/C�}?��0�B�pD,E.4D�sQ�*V�x}p��߲<m�ab"4D��Z&��$Qmx���/V���%�3D�@)�M�8��=�B�%:�vX���6D�0��)��N$���.�3^�`��b4D����.}�d1@�%�"�k��1D�Tѥ`�:?0�Fj>X�V��3D�<�h\���\k�
A9vk`A��A/D�B!I�a������s	�.L!�dV��"�!'�\afH ;!��C$=f- ��۩ D�6g�}�!��9J�`s� �6R'\Ȣ0÷m�!��;f���`l�\PŪޔ"�!�$�	l*�q�,� "�H��e	J�K�!����� �)*-^�iI�!�Ĕ�5*$���zh�ѓJ��!�C�L(Ӭ-/J��r���H !���hb���w�
�p�����i�!�æI���+5h �2��s�����!�$�4Z�l�)�i�� <#!�T�l`ZB��g2΁��@�!�D]8G�3i�:M~��"��3q�!�+	b���C?eV9��OJ�!�䍑T�kA��a"�����E�!�$��(k�PY."���.9�!����ꕁVh:t�b�֣�8B�!�$A� �h���3#�ģ�%� Vl!�E&/�H�&̤0�<��$�V�RO!�d�7w8��$hJ�A��YB�զ2!򄟋(���!f�IY���p�O62�!�$4RG����G��j�xv�٧[M!���Z�nICF�S Xr�b�5:�!�Ĉ�7c�Jv-ܘ����R!��n�X���:�p�v͡o!��]�T�T�P&K�I��D�o!�$[y͂�����c�V�Kq��R�!���[?����,�~�v
�k�5&�!�d	=B���bƊz�n�#���H�!�DU�LmT��"iU1B�^�)��ͷ) !��$?�ޡӓJFh��G»V�!�DK��]8��э	n�Jc��7!�ձ[Mz}ڷC�(V�h�7�7D!�$πCZ����Q�>R�]Iv�##2!�dQU2 P0j	</A����
"!�9k=�e
A�]�-H�R�.��Y !�DN�,�`Ycmޠ|�M*�#�1T!�� v����?X��+ʘ-v�$"O��ڐ���U�.��#+��:����"O|�
����~���&)�1#�~`�4"Ov-��#��
�*��D��½#�"OҬ�E-
#K�� �T�-�~
�"Ol�ӧ�m@"Q�a$������"O�]@���$��J��T(�D�Z#"O@����T8:h���Н�.�a"OT��WF�6M|���b�$����"O|%���[��0����ݮB�:��q"OP񩖇'c&��G��5t�@9b"OD�!u���)e4��O�PIyw"O$�3��!w�z���*�V䩠"OR�0�Ɲ�tU�=Ф#�dA	5"O\��}Kd�BQ�	:�<��"O�4��D�O\�Õ��.���C"O��cIV�����`B�p�Ҭ� "OT�&��gnT�@̑?�b�"O��Z�@0�F��RV"�bT�<1���#d���n��]�yCǙg�<a�`�r��@�t��s3�M1���e�<����f=x�J'!��-Li#�M�<a��V�p�X�qC"�G�\DIb��E�<)�a��
�p� AL0�XW�<Q��C0 0 �A�u��QeE�S�<A��A�S���`@�ϋ�r��N�<1�M7-�>�y�&C�~gHaj�h�d�<Yl�0=D �W��8�L�@�΋a�<Q'B�i��=�2�+<�r%N�f�<�&��>@mR�#�&]��i� �h�<�a""���EE!<�u�"B�k�<� ��Z8qf�ğJ~,��!�b�<Q����b������@C&�[�<Y���s,.)�#�_�<`̥A��q�<U�I�O{|YR�C'g��U�n�<�%�7�\�B�!¤y�����)Gh�<��fO�W��!���)h
��7��e�<��
3=��s͉�F�ၧ��L�<��o�8
1h�p Ļs[�0S��P�<��d�?Y�|�P������L�<�fCQ��3��9)����f�D�<��kA%T+��c�lۏFr ���~�<�` ;|�iȀ+ր���R�|�<����e9����GQ�:(�pb��u�<��40 ���*X�Q��X�䭇u�<ѥ�� 0H�1�T�6��|a�o�<����n��Qц�UWr@	�˜m�<!���X��
��|0��HR�<� M{)��|	@��ao)#�~B�I�1:�@�N�5���e#A%&�bB�I�?��X@��@�_��C�ɧ|��I���onX�ZE�BE�C䉌2G2 �wNH�,T��N��&4`C�	,G�uk�"c04��BIP�6ÄB��/ R�փr��U�fL?j~\B�	���C։@�d$��Js�,	�"B�I��&4ۂe=Qx���AQ�T��C�	S�4p0V狔]j��)PNLM�C�Is�B|0�(Q,"3�̑Sk d���?��?����$$@F�ϬR�M�D(�
�y��.�j�'A�O3䨨n�6�yrm�U�②�d�/�B��v!��y�6 h�yj5%��R�+&����y2�N"X�f��E)�\��Z�0�y
� ԝ��&��@��f�˳i�8���"O`yaDE�^�p��7�^�j=�t�A�ILyR���X)��g��$�PbC�Ke!��O0o' Y8U�I� � �*g�ǀ~T!�dS	���Њ�<!�8Q��GC!��	�[ލ��ϖ�h�����,'!��#���¬N�\ϲp1'KX�!�dX+dA�xb��Q�y�d��jP�r!��Ӗ8.Xy�ri^�*�"���FAQџ$������|�B6�T�{P����D:pM�P�<i�C� ��I��M���Ź���J�<i# ��W��Dr���B���S3�G�<IP�I�4�:���ƃ�4����ĨJo�<	RF�2�6@+��D�0�;Ьu�<�SJ�6t�����c0�	��@�m�<B�+ .p���ܢI�2��b��l�<���R8���Is�US4jEs��'T��
Ս΍kf���1A8s#`٫U2D��+U�}R.ðj���8k�J0D�|�e��4�j��^�q��Q��/D�p���u�ƨ�p	��YC�]��/D����-j����4�וhx)�4�,D��q�[U4$:��Ŷh�4*D�6��B��k���V�X�b��NL�<a�DRCR�ڲ��9u�x�9 ��D�<�Rg�<�:x9��R�����VE��<94C�x��
'Hҽ+�D���V^��%k1D����h����G�#iI�=�D%D��yg�Q9\�.(@��ً��-)�A"D��� �@)�J ؿ
���*Q�!D� :���{X@��A%���A�	-D�h�j�q�����D��l�8�)D��rV���~����kK�hsׄ�<�+O����#��)�A��&��c$.��q�!�ĉ�FA��㳧��#�0��G�#�!�dѾ>�FaʳxhXl�#��wt!�ڿOzRd�!�(� TsD��
b!�D�>\4a�����A�f�ZsU!�D�o¼�K �C��!�~H!�r{F�!����h�d�ʸk!������rr�ʑԐЄ.l_!�d�[�I� �L�Ftb�ퟋ,�!��Dm@��! ,	�*"Ԡ����W�!��X�ıb�R"	���p/F�E�!�4c`�(�jӬ	��xQ�ěOg!�d��a&�!ye���^b���.�.D�!�D\���[�I�|��bpm�)|D!�䐿f�@�0��)��(�k�|�!�� S�z(���WkUd24EܒQ!���r���(+7�r��Tj�$C!���	A���ED�<��3t�)!�$ľA�\�A��R nJ5Q�Iў,��I,9lK�.�0u�0�TJ�3�B��e��p`0zībkK�,���'�S�OR�e���+phf�R�[�	>4�+#"O�2���*fm�I�G,lPJ�"Ov����{����P B�]`��"O�P�������J0"�&��"O�,��fX	Fl�h��"9�L4k�"O���ʓy��V��-����d�|�)�G�"Q1��"e���Af)@6���?�S�O���S�Ɔ�|���:�c�
)�F��1"O��pa����`���Eu����q"OB]�PC�*L�u��)\#��Q�"O� �!�(=��(S�^��<M9�"O"	��Ɏ�Vk�d�C�Y�)OL�X$�|��'���>����0HI$��d%��{ c�<	w���p��y��H0z��M�c
�4��|��|��D��
´;��+�H�b�m�<2�!��5��d�(�����pOF�s�!�ϱei�D�c�Aw{`4�$�"!�d��� gM�Ye��"��L
�!�$E�������� D��!���'�|����3WW"I�U,�8���Ȳ�4�vC�	*Q#*�˃̒����z��U:���d�C7�"~��bC�����'����k9�܄ȓET�ຄ�,^$��B��Tk�E�ȓw��C
ٿuo0e���%�Vd�ȓ1�0��e�U �Ar*̞W����ȓv�2��W`C�ΜMQ�l��l7:��?����~b�%[9(��j��
�`�`���YB���hO�'
8�9�DA�.q�HU��'o�6�[wl����<E��'�0i
�(��?��=[0B�\�b10�'�Xܳѥ|��GH4M�>���'�yxЯ��n�"�����?�4P��'sDt�Q�ݘ8���C�31�t��
�'�l�@��ؙ@e���@	��W��1���hO?!Cg��b���4`}��5�h�<	c˂�Mhek�ծ=((�BT!�⟐F{��ɚ;;���2
F�M!lUcD��)FB�I�'^fܒ�%E�c����C� t$B�	�?/���m��P;�]�Sn����C� S&��\ %K���C řS�^B��dM�$�Y��a�jX�˚���;?y&%�rh=33��K6t��ey�<y&I
<��qӁo��e���&�Q��`E{��)�h(i9u�P�n���jX�4�|C��-$)E�R�)���� .�.x�C�I=!��q��/͗ Z�M��C�7��x�a�<$��Y�GB���C�I�E���w'�*ފ�CIڔrӲ����O��ɮ;���y7*
����B���0�zC�Ɇp (��Yn8�@�V��.,�T��/�S�O��Ic#I�tډrCL����v"OL����Ӓa��u�4��+H�:�;�"O0�Pr�M2d�,�R�� 8DV*e"O���q��)F=�HDn�$��W�'���"G��$��J?T��w!�?qbHC��<	��z`n�T��`��-�#�nC�&�*���ؐk�h|�Q��1˞��Oj��{�'�v x�@�YI��Aqc�g+�'�f�؄��7Y�dq�	��� ��',5��D��4aES{.�L��'2�0�ԂXH�AP\�o� y�'���+�g#$�\ P�,P`��8��OP� f@D��Y'��r��"OL�:�e�]&V�Q��&x���#�')ў"~����)
0d��L4Z�đ��P��y��H�>��£OB-Pm��9t���y�)+G���c��	<I&��/I��y�A4�z���K�lp@���K֕�yBd�F�ڒ�!e�����%�y
��Nm,���X3gG&!q&B7�y�hC�<~�c��\��BA��y�A�|��ԤV�\� :���yBd@�Xc�|(�B�Lx� q�ė��y��?>X,�`K�G���U�Z(�y�h��
hIрǭG�"\p�I[��y
� h�c�"�.��)���c�J�{%�	\�'8�hCF��v��:��
�`�+V�'�ў"~"��W'7��k��O�y*ѳÜ��y��>.�	��_ o�
�R�H��y��=C��z��e��X���y��ٟV�^l����[ P�1
��y�cܐyҔ `���L4$��)_ �y"i�'.��(�"U�w�|!!M���O,��?a���T�UB�P�������$P����yR-�V}H%Q�ʊV�|�nS(�yb�
�7��iy�D��N�\17`�<�yBHݲ4��5��,G��5	4�Q�yRUd(P9RӤP�:;@�s&��y���?.T�i��o�<1�M��g �y���38�]��#4y��t0�����O���.§4�d����L�s:��d�א8%聇ȓ���� b��MU����&��v�z��*�.�D�Y,��f.��[�TD�ȓi�A@$å��8ۅ5"��1�ȓJ� i1�@@�~S�bƯ'^�����@�ۍ7j�D&^"�6��ȓK%��q��T(Rٺ�@,�,�F{2�'W?��/�3¨H���:@s֙x�N4D� �Ao�5!���4R�Sg��2f�,D���D,��A�������A�%D��j���8Ch��z�$0D�� 2'�h�TԢ�,R�1%���7�8D����δ;g��� #���8U.8D�,��	J�~�z��O��v� �<D�X��ȬTDZjpKLI�J4���:D�p:��Q�]0�PA�--$��ah9D� @�nÅu�bXɞ�3�ꝑ�<D�@��E]�IX�0��m��bd��b	:T�02fF��4��cQ*u��`�W"O0X Џ��"J�:C�
��-C�"OP|ۀ担q�N����J�n��Tc "O~-+�^��p RT�U�]u*�d"O���j��|j0��/8y���"O��À�M�E���FN���F�y�"O:5�W�g~�5���ϙZ��YA�"O��0��5�~��2Iމ;�%��"O�8�` ȡ^^��g�"���2"O��J�gV�oh�:UȂ|�@��"O�C����M�ȍ�1�S�K��l+�"ODi�D�0�"��䝩5�x���"O����>l��*��C�Dn��hF"O`���F"^�A���3GLL���"O&��j�V���[����d�0@"O���%&9^�F䡤oM�[�d��"O�<�hu*,m*g�A�4��"Ob����F1	}�H��Q�&���k"O^��C�����H)f��E�x��F"O��c��#�LxP�NRV����f"ON�@3ژ1�H�$�;z��r"O�%b��3D�M�#/�N�����"O~�)�+8(Ҩ#�.��'���6��Y�ȳ��i��}�����nPS�+�D�O^��� "Y]D��ކ4��3d"l'!�Ĝ�JT��|����#�
e!�	V�T�3�N {^X���aW�%�!�$�0?/hC���z8|� ��
4�!��лz�|�Q�똨%&��z�V�1W!�;c�nd �Fk�8�"\;�!�$%�Ԥ�v�4A��ҁNC������Iz��� ^�J��E#p5f��$��2ȂuYW"O� ���;��a���W,���	g"O0�+�5-�B����MB�X%�"O�z�
S6�hL`�Iʜ�Di"�"O���f26z��5N�%TD��"O
��F��5f��r�,_Op�"O�Y q��+X�5,���	H%	E�m��Q�H�S��I�{a~@� ܋K��� �ϝY@�C䉋A8���СZdJ`�4�K�1/�C�I A������3��١'ʕ�(C�ɹScT(����!p�!ܕX�FB�	��H	��ϙ/�ڹH! �6tB䉺b��2'd��<h�xP��;:$:B�	�L$re��G9�,l�c��	v��C�#Q_����L2Yn4؁@iԉ�jC�I�_�F̱�J�����w(Q"�dC�	�k�&H��FS�	[ȉ��,	��4C�I�Gz҉���Wy����"!(�C�� Ӗ��W�V.|�k��Z�Y1�B�I*����`D� f�6K�%c��B�&3�J��2�ۓ-��@�ǓNFB��o�ٛ!�	9L���d�+Q�C�	����G"A� ���ƍ�Da�C�I/���!"-ҋ[��*��L�Q��C�("*�����	��8à�
�uaxC�I!<Š�R���b�\��cE��pC�IVT�(���hGv��򤈡z�t��>��|���
�jw�u`��]lGƙ e��8�!�� y��y
Q�Z Q8��wc�8H!�dџW��Y���%wN��RGiM+!�Dч�Hy�$���K2.�)�I��!�U/0�3��_�z��Xy��R�!��ؠ|��Ĉ��;�l��%��<�!�dEP�!�E�$A��vH0�џ�IO�O�B4!��Q�N����A�D��'�Ĥd
�Q���Q�:	�
���{�J����`K�+��u�!�d�&<�&���d\>V��ѤjαXD!�J������\�EE~Ux@i�N!��ؘ�����M�f��E�ah
��!�D����f��%7i�Y�ӆ��'aa|�
9¶�ӄ��`B���y"��(̜� A"�����2�ۗ�y�Dޛ"�0�Kd��b�D�B�Y��yn�8�����j��T��\�y�����#�9ic�k�cF��yr��$e�-iv�(u&za,��y®��\��5!�2jʪ���g���'aў�Ov�
� �1-Ju*��ڤG����'�d]�
^��J��S2"A��	�'��ӷ'�
�a`�#t}��'n��Q�M4$H�����	�z���'��=PP��(p��3�k�#�<��'R�l��L?~씋&
ӡd�V��	�'e"ećX@���EW)Y�X�A���?����������K�� 0V
ŀ�K��һ B��m��$�*F�7i@�f�.�C�ɨ+�0l�sD���	H�Ş�k�C�IT� E����8Rj��OپC�3	Y����C��	�̀	dٮC�	{E�m1 "�̨�d�W�B�	�3�ni��� ~�t��A	����E{�O��d��TT�(A��f*��B^	_3�)�'*
&�
���-h�@��Y�\��LX	��� >h�4E�"6���ffI�II"Ox���bE�E����Dȴl��њ"O޴�ƣ�(4�zfe�(��=�"O�I9�Ja�b�"A.��.���"ODW�h|H���Xj�����P�I���OC�� ��aqD�%@_)K����,O �D1��p�'� �c=&�(e���ݴI�$��'�n䢥��WHTh�"l��Cs|L!�'	ɘ3��uVH��ʞ�?���3
�'�nѐ��C+|���e��>hZ� 
�'��ӧ��� -���5�K�2>�h��'(Y�h�jؠ& (�̂��D*�`�I��B;� ���R����'�ў"~r��Ϳ4�v����(Cff$x��yRH�j"��Y�`K:wz<P�Î�?���S5X�|��͓~}fe�Q�Y�^�B���a�8ѸrG�) zN(�D-�J��ȓ&z̅ I��S���(w�U<z1L���F0��Pq��F���S��R7Zj^��Io�IVy���G�(&�p��+[��E2�n�(��C�ɸ9��UK@�ΏU��Y�a��e�B�ɖ
W��dd���	aFA]�wp�B�g�(�rC�ɒA�H�h�ۏ ǸB��5JN��¤�V  m����^#�B�Iie�)*��Nh�TiiA�A4��B�I(#�����!M��y��ԏh�|ʓ��$��)w����MA38$e*a�"�R��A%D� ��S�(���1�dةF" D��kp�Z-_�T̛v#�"�h��ad?�Il����	 Pp��#i�2Eֆ��adV�LvB�I�fH<�g㍊)����a��#�dB�I�M�����K^d�Ԏ��38B�Iuʘ�zv�0*�L�/�:C�I3_zpuHs��wmn�ɉ23�B�ɝGw��rE-�fi���H
��B�	�K�IH3Ɛ��P=.")����?	����S�O ���rAX��Jq�RaNd��'��*@��#�R0/�=X�&�P�'zv@� �R���'E%A�*m �'��	GI��V��9�3���8���)�t�������'�59��x����䓺0>�5��	
��\)s��V��v�<�`G3F𱒇� {����b��y���hO�'��,!̟F@n\��VD�ȓb]�qG(F.8�az�J���LɆȓ��d�3*D�����e�)Br<�ȓ,�Z���)�*�
q����1:�2��?Y���?	��IL�c�
Ա���� �sp�,(V!��4	�!�e�߹&�j�al�  Q!��(W�[ԉ�(z&a`5���Iğ��IS�)ʧl[���%Z$&{p�Q� �N����c�� �S�NUjM���X5:D�ȓʖ)k2Ϙ�EP$iQI��y��1�ȓ8��"�G6�j����(�G{B�O��1��i;I���Ë�f�ՂM>y���?�t���?�b�ձ��Os��H��<J�Ju���Z�B�H
�'�0:4�
>z�mX���.>�^I�'Nv$2�I��ܽ��� "=e>�I�'����8\�Z8�J�9#&��'<�ɣW���kN��# ��>'�zY@�'�&���́	�dç�ėLR�9�'Q�aÐ�@�C����W+�t���S�<dExb�'���xp`ۀm���#Aٚ�y��G�}�(i�6,o��\�@���y
� �0+��L�s�� Q�^�~�|�c"O8Mj�'�i����C�09��i��"OR%��m��T�f�h�m�"V<:02"O�tу�'���C�TY��T�'�'�O^��!?�);���ᢘ?{@f�E��P�<1f��6N���J�	�:Zl3���h�<a�$ό�@�!L�cDݺ��{�<i��X�lRX��	��z�e�\�<Ѱ�{�0ZB�f���u
FX�<�QÕ�=��PL�|�9p��V�<a@�K0�ҴB��Jz�(]` �V���hO�R^&�a5�$�Q�cLn��x�ȓH.���J��U�F8�-�Zo���	_~B됪W�J�R3`ʴY�h(�t�^��yrf� h��[��Y�"��GE��y�'ՠjƔ�Q䜛W�� a�)�y�[�M��9��P\"�fٵ�y2�ΫN��@2��[M6�kl߅�yRn��3U�T�'S�E�ȹ@5%C5�y�N�5gs CI�P�h��DGۆ�yrd�2ڢ�(�ʜBt�X�êT�y�Hٍyr���@ϻ?�Q�")��yB�лz��Q��F�<�t	{�$���y2IK#M�A�#M!6��U�a�X5�yҬ�df�#�
)3��	X��y�Ƃ�v:���ֳ1�$�Q��*�yҢѨR����������B��.�yBL��z�2�A���a��oE��y��L�!>9Ġ�*>�Q����y��έ%��S�I9N�QF虑�y⢅)Gtz9��#�4�ڴ���yR�؀EX���%ɕ@r�����y�!ߓU�ܠ���t���aumM��y��)P��Cr��>���t�P��y��[w�D��46�&�s����䓒hOq�n5��0��)�F�i`���p"O�)��"��\q�n��r��"O��j�b��QrT�Ĉ�"O��1��E��Z踄J�?��p�"O��(��\8"�Ĕ�E�PN���B�"O���a�R�`  	f���_ƶ�QU"O$eB0�F�q��oS�f����&���O
��&�Q]~G�FS�D�F�Z��	 	9#��Q���5aC9A����K���Q*		N���b��o^9�Ɠg3�"Q��6om�c�oT�KҮ0�'���v�K����Β�<5J���'\�ppU# X(�Aē�/�ȹC(O�$/�O,��M�
�z�j�G&EL5�5"OZ�r&�O�����:5t�"O�(9��_5�
]k��?Q�=z�"O��� ܕ0���񁯄4D��iy�"OJ���h�
^$��R��U�:�(��'R�|��اdע �� �4��9sdF>D���&V� ��ȡ�G<<	����I!D��� �_�p�p��--�n�H��,D�l0�
3R�`�ǫ�s�`��4�,D�X!'��7;��A��=U���H�*D���'�ْ�ĵ2Q�Z�	,%��(D�p�!j�$�NE	ŮĴj�V�{u"�<�I>���O��k��i ����ƙ40�tB""O��Z���U��\r#��z���1"O@����L��
Ɓ�AR�3"O�`��C�&!n�� �;H����"O� D�`��W*ty�$��&]��ku"O�4iVhJ�*�z�#��̑VV6��"O�\``E��U8D�B:!Gd��a�'��|"�)q�ƿQY�]����6�x�B�5D�����i�z���D .e�f��$�1D����  �Uӳ�\��N�K��/��B�����c�n�SS���.�}+VD1�C��	f� �@/θ!wzy��Mr�tC�I�A���� �.ٞ���+L;H�~B��xON�x�n�[ll���G,:B�%BĺI���Ww7ZD��K��+А�	H<�'$�k�P�h�b���|k����<AQ����g����#��� �q�`��J֦㟔�	>!sU�'qd����~{�~-���5D����@�� �۔k�`���!D��
���Uy���]�\�2�C��;D� �����]�$X��nێ5޼ᨦ�8D�8:#�X����*""M~ VPS��O���8�O~Xg��O_�	#R��*o&����'!��$.�Р��˹C� ���aéL���r��`b1�+:AL�͏�_ɬԅȓ5�@��h�8���i��z���m��c�9�Lиb�\F��E�ȓf��Tҵkɐ����ǗU�Ṙ�Yq�\Q&���
A�,y�$`�'�a~�n��`M�H�NLي%HS4�y2A�M�89Q��w��52���
���hOq���x�6�
i��	8�����"O �0ǃ�����P̏ ^f��A�"O6��cË29��"�=6=5j!"O2	;���>d'�KP��o?�MZ�"O�<����\�HФ
� Cx�3"O��)�G	$M�V�P$�ۮ%�n�(�"O$� ᄆ-x����f��X���q"O����c�#��41�U�]P$"O�e�� (-��8cJ�1U��c"O�i!b���}�w� w�,�"O ��a�4��	�#(R!Mn��w"O@� �� �Bݨ@�ӌ9 �(�"OZ��d�8=��J�>a"0PB�"Ot�hN
`D x$�_$%��d��"On��r��!4���dH�e�1;�"O6� teπT� ��Ħ��D��"O�̙¢�:����H�'Ά�{�"O�:�@U�+Ɣ��N�&g��1	D"OX`���4+Cv�k0�_��΅�w"O�tk�N�>e�*�Fѽ��c�_� ��g�S�O.-��	�z��Ր@�+���'����:"�ڹP�ˠym2�C�'�,,ɲ&Q�����A3�,("OJ��Qn�6L�P-�ƯӚ$L�)��"O��� V-%v�Ń%�I�FMd��"ON-�S��R#Z�(wMĂC�(�;�"O�=���(���ap,�v��FV�xG{��酴^��H���G���B��~T!��A%-u�y .���0y@`�S!�d�?BZP�) B:z��$��[�!�N!p�؅�� ÄZR�W��1N�!��>mܪD�%N��$Y�)@W�!�݊J��E��)�;o�:�'+֕k�!���K��E�ʹ
�XسhY?c�!��HZ{�Y �p��uS�4u�!�$-/�u�aϙ8���IW���S!�D��*ފ8p ���ꨲri��%�!�� �c�Αg��t�Eg�8%
]0e"O��Y��7ZT3G��2��Z "O
!�*Әg���Ae�U� � �"O�,�"J�iX�	@ �N�B�b�ʰ"O��0d�#F��l�s���fc ��$"O�D�AE؀F�81#Q�\pd�0"O(��"�X��tR"��r��	�""O�5��E	=�ޡ�� ��y�6,"OhQK�%����G�*��A"O(<0���Д�T�I�N�p�{�"O��{�瓥%� Ba�F���"O�H2�ȊdP #�.�=)^�D	�"O�2b`
YL��! ؒW�"Or w�Фw��I�P�Z�l���"O����ѕ?�|�ޒ"�u��"O�a �"A+Qתm�UHT�
�P`yA"Ob{ǚ�-�f�RF M�.� V"O��@��4b�Rb��}�$��"O�0�Zi͆�r�A�=��G"O��4�l����L~q
�"O�qB��f@�:%�=#X*d��"O���pc��2B��Ʌ�V3#U���Q"O� 
�gO#� ��ᐚR8�U�"Ol�Itg�e���J��/l�U�"O�ei�Âg�<�5莝����"O��9׀�`�,��጖�pw�(��"O�,��l�6IY�I{Em��|�c�"O�X�h[�M����l_� ��A�"O�!��9R�\|�6ҹc�j�z&"O�Y;���CrE��
�"�B"O�$�f�5g� 9xK<jp�)p�"O��*&k��a��U@qj�o~�-�p"OĀB%O�.FP����!z�%x�"OP�XP
�O��QE�\֞�S4"O� Iw��:*}pXk�N�+a:H�@"O*)9���Y����`�Q�l��C�"OTM�R�
����v(U0n�x�h
�'������*�LLq�6Nq�
�'?�E��Q�l� `�*Cz8(!�'C�A�
�!	���0�W�@�fi2
�'o\�+GBU#R1 ���`�	�'*`��EʣLf���GF�t��'a.@�똚�R�B��T79��Uz�'���	�/�*%�%��$578`�'�R�
��9 � ��C1R1�' \y�G��0C���*�T�Y	�'�d���%�Cp��Z�F�+´l��'3<����D)W����V6X��qx�'Vt���b�$2|S�#ҞI.�h�'�pᠴ�ʌ���[whG�P�e��'clh��`	�I�q��?W�z���'�Ԭ�&怫t�@0�ը�?z����'�
�a�S&�5�HO�k�\���' ���7H��uޤ �,�h�(���'����.�Fȱ:�� *h�=��',xA;�ϥ}�j���SR&	�yIS,�HrQ@j�};�k
<�yr�Ċ�d�+h��f��HX��ȅ�y�a�6�2�j����h���tGܼ�yF�N�J��W��]�� ��NZ��y"e��A��툱c���i%�Ü�y29�ر��`^Wx�sSeٛ�y�N�h�f���AI&#����R�S?�yX�;�s��L
���
r�*�y
� �h)c�W�"
�y��Pn$�e�!"OpĢ�B�nc� Wcm ��&"O捩F$K�`��P�mO�0R,�Z�"O�!���V�V�:u��_��x�"O��	�&g8Hx�3.�	e|2� "O���c�<��1�l�-n�F"OVB�a 0&���1Vl�r���"O�/��[��s���df����!D�Ԁ�M.7W0�qbD��oj� �=D���G�.SXY�1A�O�����!=D�p���>_�(��u���w։���/D��K L��2)��-P�D,D��0u`_(#^a�a�KV���rr'D�ܻf�N�`R�QC@�ǒA��y�&D�r'ew֥[�ؑIp�sB�$D� �IYjoJi�����V�@�g>D�l����v�$dQ��B��
�7D���Ҏ��g��ٹ�L�*�@��ŋ D�(�@j�8�1��B)hTF���<D��H�d��d mJ���-#̥B�:D�D[�F,M�L��N^���	�:D��J�W?H.*���o�SY�6�4D� �t�	 mq1C\�)u�4D��c!ξa͆Dy�@ 0�A9Ѡ'D��c�o�x�2���
Q��$�g�:D��p��]l��j֫S"r �H�6D�p����F�X�	c��O[*��4�2D�,Pa���<`�g.�0��|��%D�(��tFΌ�꘬b�T��-D�h�%�ۺV�ɐ�B�Ls�|��	.D�H�n�-|��+%�Q�'f��2P')D��
pȀB���ۓK
 *�����%D�0� ��5yl���e	�8B�a�!D�Ț0+��XP��
v/�(a6~\s�N>D�$Y�O�*Z*��bt$1M�����<D�4�\�#*!⒩���z�"M D� S��t�:���/aO,���3D��u��<�{�,�5
�m�C1D�HY�'�, ���+�̍�.C,�.;D��	G�b�r�bŊ]�
�@�7D�Ġ���L��=�0`ɔ�YZ�!D�@�U��>A>%��-_� =��<D�P�f$P:Z&Jȹv��Z(�Pd�<D� �b�<4�I� �	����g�/D�|���d{HA9��0��0"�I1T��If��yn����ˇ�k7!�4"OhEBs�6F��㇊�-Mh���"O�0i�#�9+/İJ���	Y9*X��"O"��-~��ڢ�߳Z4��w"O�!8W�E!�zq����7�x�%"O�YG#�1wh�2S��1� �"O����
2"������"!Ҁ"O<< qKZ�JT"wV;E�Đc�"O0LhO*6H��2���;\d[�"O�� l�4T��b�CBSG���"O$=��d�YgX�cĉN����yb�>M����sfD��<Yچc� �y��k��}C�A�y�80ƧC��y�ܓg��sՌ�-��0�բ��yr+	���LS�rh�%���y�F�Kl~���膗k
$���ᚶ�yr+T�3��웄�NZ.�Ce!ߍ�y��1!`D0�� \�6��TrQh���y��7f(8�k�� �X��f�]!�y
� 4u��%D�^�$���IY7���"OhYrh�%M�&9��̎���"O"q)Îԁpl3Qf$��k6"Op����/b�0|���&"� 1"O�d`�f��o�*�H6Mܫ9� ""O�9�"b�-z�Ġ-Ʊopv09"Op��.�;a�<����54T�y��"On�s��
}�N�a�ٟG�e0�"O�T�D�،OV`BQ&Øb=����"O�H6�ѣ�M�7eL3}04"O�\9��62kg�Cev�[q"Ob�&#&:��!e�<Z{^��S"O��`�i� �6Ku��k��B#"OfD��E3!$��d!ւa�.t�S"O*K.��;L\`@�C߆�y"O��3caF�gqR<xP@�r����q"OMxT�5_,�M)`	о{�"1�g"O�5� �"N.d`�F�W昐;�"O4�@��~���s�%��9"O��HE�-`!���	k�>�3�'�Pl�p$��:���ч<u�l{�'$�жcR�\ AKW�dI�	�'u�İa���V�H�p�j�}f�*	�'��4KlXazu�ǅj٠|��'䲌`𥗥  �뤈��dq���
�'�ʰ�4��+	 r��dH�c�@@	�'d��sf�| ������_6����'�	��`ۆF�`@��Q%�z���'�Y��b�-,��@fE�4#Α��'ښ	��Ā$����G�&�y��'|��QjH Kz�ɷdB)S�e��'�>��V*HA�������0�=j�'Ҳ"���.(zK7@������'V6ra���豙����U
L��'tv+���}�HE���R�	q����'%�2E@ѧeW�tF�{[^aP	�'�u0���7�U��O�8s��t��'��a���g��avi7q���'�p����4@���z`*	�'�=W% �5��2ix(��!D�: b8p�i��!���a;D���Ƌ_����bI$���)9D�0�C�ߍ#�ڬIe G6d>��[e8D���R�.���G��D�5���5D���NxI�#�,!
�@aa@?D� s��R8T��@�RE(qi�i�C?D��8Q*A"#YhaI��";uxhɷ�)D��Y7���8b�Q3�m�\@>���&D�tKU�!")H�pB���4�g�"D��sv�M�1����5�@�`�٨��5D�ȓvĜ���b��K�l̾)C��2D��s�I�{
^ �,��Z=V�ra�/D��B M�j�zl!��@��hP�2D�������4�F�O��h��*2�O<}�O��S����K���gj��~��̋A�2D�|�5lF�K%���?g F�2D����G�d�8�'቙H� E��O>D�T��'�+u�aX��=@�(Z�#>D��	'kN�e�� �&E�j�d?D�l�Ƣ&\�
���G�Q�XX*��9D�p�̏�/�$Hjbf"k\��M7D�pҕM�.��@#b#���j�0��*D���Bg׷sfN`�p�P�te.��T�(D���Vh�1g���mK�a|ހ�si%D�� `��#Źd�� 	���rM$S�3O����]�Ԍ�ĂW�#�蹱#dS�n>!�$�2�ji����;$�ݳDҡ�v����X�r���efF��@�o,��hO���+���ڂe�m�a8���y�x">��I@�<SܙB@�%����n 1!�ǘRG��r��۽Q�����)!�dЎ
dȜ�whU:Ǻ)����F��O����5b�B���w�ΰ�f�2��7�O��#�)O1�*�R�����}�"O�X
cj��o4���eȯV��	��'��D�t�>Q�4��z����I�tn��*��DRn��yrI�o��q�+�@^�鲤)L	�0=y���W:5fHhAgKٶj�bĬԮ�(Oi�� ڹ�voW���p��hV�vn�%��E{��T!�
B�$z�߄���KU��y�`�!��Ѻ%��ީ9����'?az����T�؉�W!6�^���'J��p>i�>q1B�5��Pj\��i RƎßLΓ�~r�'b?��O�N4+�
�>��f%Yۦq;��ɧ#ĢZ�#��!U�	%��W��{��n�<��!CI�$�����&dS�ٕX!��Ey��)�OvXrf�ɞvW4���E��9��Q2U�@��	p�p1�W��;r���y���Ysh�	�a~2	�G�t1��p�a������>���<��d�Hx��Q.��YGXix��	D}��'�icfg�N�[�,�R�1�'A¸# ��6�p,Yf�J!H���'��M3�ǵ5�d���H�@-v�.ON�=Ys�Ę�.�@w�7��]�QmR73��	a���;��DC��	���/��q�%�7�r�L+5�O�`崽��)!����(6D��y��;=�HHS�+ {b���#�uӈ��m̓e�Q?!���ȍ"L|�ad̚Ίɑ`O>D�(2S&7� sSO?dXEԥ<D�ܸT皣J�fM��K�4%8�$:D�h��Ȇ�n�P�[��	n���o7D�pRb`�Tl��@#�C؅Af5D�,�pFۿ-Z���hHH̚%C5�1D���a�
�/�R �¢�(4d=��;D��pb�W�%���|rdX4�%D�h8��$��
��Q��H�T�#D� Y �"3,�i)�`�' �@g�5�O�II�F��T!r֪}	1��+?"�B��HM&E��Z�[,@�F��0��B��)�L�K"K�*�@� 蕭-E���$�/U���<ad*J!h,�"q(�{��}�؞D!�Q�`jqJ�G�e��I� ƀq'!�P�/R� ��i	*�d��c�!�D��7�VL����a�B��S�HD���D��,T#Ԧm`G�H�\�����!10!����B��E26.���P����9+!�#0�@ԲLG\8��C�ߗp!�$׳xsT��Ś� u\h��b��P!�$��x����C�)6���8���)�OpHP�{�����&�Qwo�1IGh�!BL�:ǒC�Ʉ2X�ar�B�&V<���g�mfC�Iڟ���G�F6er�AE�Z(��
��2D���1�]�/�
[d�C�X��;f`%D��ȡlB+'@�5b��η��d"��"D�4��ߋT%�T�G?V�N�6͟jy��)�'I?���!ʗ�8��T�����K�jчȓ'�
pH7�� ,��@���Z~��� D1A2�]�%<z`#���BD��'2��z�S�π ��[��a��䭟7M�R�"�i���o8�Djs�Ϧsf��Y�'6h1�2�(}�)�ӫU`P�A 2^p���һߖC�	%m.t�f�\��z�#�Q5#%���&������?8|���Av���(lO�Lyb�'oX�%K����!Y0����	�'4Xt	�B������2fp{�'L"�I�`l8��,B>UX�bO&�y2/�W�B�*��F�Ѭ��1c���=��y�X?x�`L��BK&I���!��N��y�L�{
C�	J�"�qAk܌���;��&�'a���0�ǉv���`��Q�;�L�ȓQ���!��6h�L؄�Ѽw��<Fz�g2O^���'�#[��8ũ̻b �%J�በD��Ix����Hȕ@g��P��A9E�p��"O P�G�B�enp`��^0X�QA��'f1O�PL��6�Xc��W$V�bհR"O���Q�D�a�����F����W��;��)�'M��2�C���([�"�M�rl�ēR�J�P���
� a��Y�"�8��>I�`+�OH�wj��p���C�ɋB0H��"Ov�eH���R�P��V����xb�'B�0rA�I�{g�"&48��x{�'�h$�7�
��>U�� �(��p)�'�LEӕ���8LXǈL�I"ы}��)񩇘N����kFƄ�ZAMA�2�!�d�;w��5`#"��`�0E���["=�!�$�O���Eɐ�̚Ē�K�ay��'[qO8��4��%W�A��툐A��ȥ"O��a�FгA�9�r�P-N^��"O��� �ϟ2�����q�.���"O�����,� ���3>B�0:���3�(O�c>�j�&�
�� ��%X8H�����$?�S�S�k�u�s�W@� ��b�tB�	n���bR0Ն�q�C�;�^��d�<a��+W4Aq�JE"(��+�W|!�E:6)r�҇a�'o�PH�-�/o!�c ��x���;��S�?$o��XF�d�K:SR�ܘm��4 P���D/�S�Of�!@֏�y��0�S	�2#�TT	�'�hI1*�7k��p�+p�h�'G`�A�#�3Z1�8��%?����B�)��<�hT9�, "t���Z��&F����'�a}�J4x�4ȗ(��~8
YzBJ�y�� &~�XƦ�eGɹt� :��?A�'����G�Q�m1&�_a��
��'�>E0�iq]��c'#�2;[�����5���2��3�޾4$p
	�T�(Їȓt�<Q�G%O��!1@� �d�dH�ȓ4O,|&��6q�z̐��&*M�)��x�.���.�� 2̤���l�D�������9��m�2J�ݚl��{���*'��L���bko�D�ȓA莌H�郭iR6H*w�g���ȓn��4[�L��,.�`Z���[R���ȓC��@[��ˣU�|˕�A
xt���'4���AC�h�8DB��d��B��a�r'�8lET�qҭ�i��Y��
L�)�B�Y=!A���[T���W���؁Ŏ�D�ũ�FA�u���ȓ]�*�䚔Jæ$z���c�V]�ȓ}c��G���Ň�7)���"O�U�G�(I��!�\x����ʡ�y���*$�����)�g,Ξ�y
� ^l���TPґ�jL�+L���@"O��� D�<:N�TKR��j,ne)�"Oz����5�̨��T�(�T��"O���`�Qܰ�Yu��n�ف&"O2ܺ�O���
V��?R+x3f"Oh�k5σ�:H�|���˖u�v�9G"O�-�f#��5������K��� �"O��ң�k��2�"�f��EJ�"O����G�\�&�BV�N��j�@�"O�a� % ���E�3m��3֔p�"O���Uj4sy�L�k��'��"OJ=� Z���ēd���3j`���"Olt��%�@�iႦʂ h��2""O�P����8 vdR��R�n3h !*O������p#�רc6x�"�':�!��Z%o�VT ��<
�:���'����&�&I��� 3��i��'����B	�{�y���ܒ^~���'۰a0VKD�j�
 ����L���q�'���ZTk7$5|4@Ņ�6TR0��'����$G]��9�U�^�'�>4�'X���cf�\�2Tݞ	����'oL��K]#�D��&C���)�&�2��	j��U<k=9�$�Ш@��=�d��h �92͆ȓUD��F(J1=��u�f��E?�؆�2��|pCV�J��0J�^�V�r��,���杸>ݪŉUD�8XNv��ȓ\���6�ǄBN ��m��r|��ȓe�TY��~Pec�*DZXx��tq� Y1�T�W��b�*�0���\�x�҄O�
z?��z�̉�X6� �ȓ<Xข1��0��7C!.�椆�k�(�I�BF(m	����5���ȓo�T`Icm C7�0��]�5�>d��2d�H���!��`a�JM�M�"���H1�̀���#��I��ވL�d�ȓZ�s(�U�Y���" �P���;%�� 2�U�|0�a����񢕄ȓo��% ֨M��� ��bZ�a���ȓJ[L ��(�$q�(Y3�^�*��m�ȓ0�x�J֣�a����t�>`����Z�>�;b��6�N�bd���p ��ȓYU>)��U�04;T�ҲQQ���9,����|B��.\v:W#\O��e ��\���
��T
�o �db�,�)T=��ȓ�Ni� )�,YP����?^�'�����׎>X��1��f�O�(͈B�v���A���z�0���'LԥA!�Io�t{Q@�1O�6А���v�с��O�q��!�u�g�	�?TU�I�Yf�l� z�B�������\�`7+J	v���`�/c�$��Et�����r�p5�T��:���F��U9b�?��h�9,��h+P�O5nX����|�)�g�2d�<�J��2?��pF�0D��� A�+(*�1����	����f��DYq�Q��&l�w��7z�l�pE���(��4J�h�Q ��ހ@Uzd�u"O&e:��I�&A!qL �%o �"���$u�� ��Q�4r�Q)W�&a2ׯ�&I9�{�C�3�����9(�(��'�0��<����)�$��G�1=�${��@'n,q�h!RhZ|��U�X�"Q�y�"0��Eg��Lj"왑A�3C�T��.�3�*<�@)Q=�I�7*U9HN�)�#�6dl�rE����9KN�=kA�k������J�z܊��Yy�'���&Ko�O8�ч���vu�CM��B���)�a�,��Pk;�MY�n^�g,����J���!r��ϻ"Z䘉��\�HM�F�I�;�%NYʽᐞ>!����u'f#]��V�,^���ŉ.�bB���1K!f=�ℍ
W�䰢��"U�9�t����'��\�� �*���ř0 N�d��4Z����5�0N�(8��.Gb D1�I? ,B��
�S�(�C�5�F�Aʓj�0X%�Q�g3`��<��Oƈ*E�ĨL]�=
� �ǀ ��ys̏5Xu��+5�[c������P)��5��Q`-^�2h����ϖu�PT�����)[wR&<�%K:®����E%K���[%BP�ʓ�$�f/���]�!�t�_��B�'�԰��N� .�T<ZF�V2')�0¨�o�5��jĠdp+�&���S/�����D�߹X1���d#��.,�@J��5��õ#�<L0��I�U�tM�'n9Y2���D�Yy��9~�����wN��X���-#, �Z�o�U��L1wDڎ!3\�Z"��/`�xE(MsE��0bc�/''��'�޴x�g�;x���R�$E<`\��4r���ǭ�%MtTJ�S�����?5� ��iP�Q��33����;D班UQ\�2Ǭ�^����Gr��J��q���еX����s�4X����]Opz�:�lI�}{�t;a�f�����-VԐ	�ƭ<y�f]�2��L�6g�h_�c�����Y,SҘ�O��<5#�i��k�GW�/O����΁T;\ ��a�'yv�D���Xݴ�>��JK��ͼ� �մ㨰����?��8Ѣ�I�	}He�A.��)�S�M�*ւ�� ���矙$R���A�*kǒPاE�Hh����M[��R���l�~]^`��FJ�Kٲ�K���
��t�EĔMa����]��ល7l8	��&ݕHD�ܙ�̂ �#�#(g�}�N:�<� ���3f.=�"��OK���Ӭ�"�3&R�>Y�`AM�
|Ҝ��b޹Rxc�#�����`̻*���'_:` ���5�~�����T�0 �RA��{�'�*GԌQ7 ��dE9Vx�����sj}�ǠA�RC��#gY	/MĨ�@֖{ t ���&�r&O�"�&)�6H�m��	�@�Q�m�	ݒ��C�%P���X��$�˧s��T{��T3���(�l�0b��@��1sZ�qc�މ��%6k�w��HK����|:��_1f�����aB�B�P8�����) �(��0i]�'.8�ß�"���:�H"�S�}�Fi4AFH��9"�ě#1֐0���уI�`%��B��bN�-B��H����1]#�zFdڠ7ۆ�7�x��t?D��Ò�p���I�z2��i���:=$U*���B����M+`�N�|Q�R+2�v�sF+p��RA��FD������!Q�P��GY.�(d;Ԅ�*Y�8b�`+��X�X�>��'}��W�;rEP�C$L�'161
m�	x����:E�,lj�C��uڬ�����tHF��� <,R�mJ�z�� �;4Lqa'�ǝO8���I�EܓI�����"��<z2��g�>C�@�<�&)F � !�@����s/�a�:B͇�J�l@!>�*i�0��Y���ہ%Ev 
��P��̩��'r���7ǎl@t�B�"͡5E�e�#��6GJ�)����/�4�D�>o�D3Ԥ0oGz�P��"3N���8�P�h��p�C��<y���F�2�B ]��
�;L,��G�]h�6�P��46�4��6g$N����>V��`[jR)i�h�t��K�������mv���DA�sV2L�2A��D�O�my�eB�(� � ��h{���A�p^ d��-@����FD"�U��J��tF�����Y�BB�	�vT ��ω3�|� �q$��G�+������9� ��M;�D4l��A5"�l�;XȬ�P�I��e��4!e��?�i���
qܺ��mG�;L�a勇Wo�����g��Z�#D [�D 5�/��AHo"0X(�K�Sf���J<i'+/"�Ic�H�}u�(�����'�b���d�o�Y""Ofd=�.׊Z� ���@ՙv̡Aaˌ�d�.��Ы*N��@���p`��2,O�3��u!��˦"�����Oa���U�GȬD��	W��8֭O��@�T�
�(��� E�g�����XT�(�܇R����R
�*�E}�e�c|�u8����^�(���Z�,i��_���+E"շ,$����4��=*1. 8V(RE��B��3�^#��%"��'<��XJk�����#4.��S`�"�t�|Cv��6�E|	꼻�˻".*��'D��~>��`˺'%:ĺ�&RVÆ�㡌��8�x�dm��j$�!��	>�(��!�%KѦ�� &��Tƈȳ,�.�ēp�ݻ'N�V��,��S6�!�-�<y�2�JU
��>�4	A���p�͋WN+R�� �㋓�0�%i'͑�$�����R�V�f��c�˓�KMZsf���鞩O����E�
�(O����/ǑYth0�2�
�3h�c���M+X{%P�/�����1&nԍۤ �4P1��H5f��'���h@�@T��s�FFQ@d�5��%6�ƐB��N�'�����GBYPD����'2�֌r���>�4�� ��y0p���6�8���'R�] 8\�w�Bk�m;a���Hp4��Š�z>d�K���2���G�+\����H»w:����LM�:��ӂ�i8YP�Nv��y��tP䰫��Іr�` q7��q�(���8|=A�T���S�9+��1��A�Ms(tHq@X�5�b���2*�L�dG� ��{co�x�I�"�꽋��X�=V�0K���G��q��_9��	�#��UZ��	d�M�&�����)ز?_�5��@�����.{����j�"vQ�U���r����Z�����\�J"=)g�΋T��a�So���t #��R���;���F���	ǳT�P*\�Ul(�@�Ę�r0oZ��F����A�DL�(SC��t ��Y��O �9"B5'`4#=��;Y��1$�
 ��(s�!4��{�U1 �x�rl	?+{,��F�X��B=C2L�( ����炩i
�}kphT3%�p�2�,�=-p8��& �6��$̏�.�Fm1·�3}�1q�3:y��%�)n*��x��� C81��NUС���]4o�8[bd�<)W��Pg��Ӵ)�3'ln8�N�_��x�L�!3b��E���OЈO��Zv�MK����k�����ʨc,� i�ߝ_3�A���>"���"�b̐O�����Xm���[��
)c(���gl�f�f�PF�W�L>8!���y�X�y��'�lX2���GLW�&6&x���*������PpjaybCB.v|��iʛg5�qg� 4&|m�yX<EIc��O���r���5�D��zŉ�ӅO�D0@��DQ�7�J����[..�D�3�F�
K�q���pc���+
�'�|�t �HT\ȡ�8��l��bL�O�$����dكkK�!�p�OI��zp���v	h��٬>�d3�'f����Wی����L5v��Z F��zH��-=�Lc�.�.b8�q��1?i�M��+݋|�Zl[Q�S�F*�&ܥm���ꄴ�0�y��ɗ���"����H�3�ӈ*��MI ɚ)�����$:54��,ߕ���B�
���\�c�
-��a����.��Y�I����� �'|/�i�@* ?�a{��Ż,@]�tC�I�&���dU�Y�0�� ��M>�}�4�ӹ[IX��eHS�p<���c�N��fK)�SdZ��� ���gD'37�Д�	�h:H�������X��}$b� h ��A����+�AA�,���c�F�5�|�2 �ő0wϺ�6HK�;2���7�C_{��k>�ئ� ����� �n��<��$�\@�R�Q� ���O�^�I�'��d�:.�
4v�X9�!3��Yq*D�a�ҭXS'L�cdm(��X��F,FN�?])��J�HeP=�� �	d��"��
6����D�>�c%f��L���Q�P邙#|�f�ŚIU�P
#Os=�IZ<xL�q���
���ć
�2��ѫ�
�zRn��Y���V(��	�l��t)!a�kJ	��E�� {�t�΍�Aˆ���R"+�'I�o��h��Ӧ(����N�<:�h�qNK���x�i
0�U��ޓe�ް �ߌKX8��I6p?�	!֭�����d�ýX˄H��^g�ʜh�I�NP6��5L�6r�"�
�*��f��*��1N�Q��Xpb�e�)K�	�� N��8r]%��ik��!\���!N�Bq��j�5 ? )�EGɲ*=�d(U��yC���#Yu�'�V���B�8K9�l
e�S�/����H�X�T
@�Wb5K'�]qx@�B�)ƔN�
t��%�uҁ���1ᤘh6�6B��Trs�A4C��"�.�c��Ms�
̤5D����&_�Lpf��%4��E@اG�t1RE�Bj�5�㏫^�QT�A�#R�x(�f�� ?�� ��F�@I�e3k�:U�Q���b�vɻD�3�E�'�M����P4�}�tƍC�lܫrnѫR�Dk��7Jb��0���=)����%6P0�Y����F�z���NЩ�E��*!� �3���!jĹ�bő�p�
̇�	�=1 � �n\�-�~��� _�Gԉ�A
� OnA�� YxT���Z�-rD�i��ٱ�F�O3����ꑡJ`a�v�^�	YiT�ʒbB 4�	jw���.��k (Stn[�P�eÀ+�UTLxh ���C���@E�7�ƌ:0A4^�Q�G�o3�Qwg��!!C�ܗ{��U�V�߅��<a@%\;s���Ϊd������ Y؁k� ͌_b�����	8H6�"�E�u���uFO�`�����R�Qʽt�C�*�(����[�Z�88�r�ϯ��?DÈ#w>���gMYB���)�-c�TIR�B}֬�e���:�"�M�#v:�0�\K��HQ�/f�DQz⧂7 &	K�LY�v�X�`mݨ/����	�g�8�{Tb�1m�RYIDl���Mx3��qutY	�*�ZDZM��z�$g�D�*����H4�i8C&�spzyY�"�9~"iA� S�&\���a�R�G��'O�Py�ߧF��sW�%) 
@jW�
�p1�Ej$�	9u)�`� ��I��� D�� ����/�1("U�t�Y�Bqb�2l=\O�{���+^D�	��!f�\��^;4M̉���#��="j"q��3D /TR�aB��#c�^2����c�Թ&^@!���R&.5�!��~�'���!U��W�O��yKc&�&���"vf�[��
�(�52k�1qB�	�eg]��,�!P�zas���$����f�_��,ReHW�6c��)��Q�-M����[K�@R�dIR�y��$j�ҧ��P$j����$�%Q@��yu��+n@ʈs�.[,`p�H@J
�N����V��s���`�W���\VHEk�&9�(O�5k���9O�: piJ�B^`m�:OΕ�D� �� 9�e&?��;Fb��K�($p�I�GTrq�S�ݲb&����08DH��x����X����V���G��L�q�7�C�����g�-R��U3p�� Wٺ�A�)ΟG�P��$�@�?J�
�"���)��KyܫáA�Uܴ�"��A�D��t��?>r��6fg��l"<Zne��( ��'T��Ki��83AX`�dg�����BFnI�t�j�$�al���P�պb�μ��.ǩuK��b&�����;`�ޔ�dΆ�sA��λ 6���FR=�¥!����c�e*0C�j0��g��Z6�o�����?�@�"߳:�,1�aG^N��ts�CS11���07�ܐVF�DJ4r2"-cCkȎp[�!�dK��XW�34���$����L��P��d$	�#���!��8|�T e`݃NJ�pRA��F��wL�V��$��!���d9~�@m24	�3���i�tXL�rf�N�Fφ�rY`��i�;.�|�P�� �W��mۣ��1"mz�s�Q8l�=W����0BUҠI���E������9ch03t���u
�mH�,N9]�%�&G�B&Q3��̘��8
�bY�4��UzCB0�� 5��u*��Ѷu�ܬa��
#1-�ps�$5 Y;��wm:A3Q��'= *�/7$z8�)w��6F�}ړa���\t[�grd.U;$�%9<����yw ��{/<EU��f�(�����(�H�Gb�VaR��=.t��� �$x)4I�O��a�F o8ɛܒ��P��B'){h���f�?N���IQ�ը�?��&�Hb<ͻ�n��D����P�yo�'�H�14MP�uO�9��nW�}V�4B&�ŜG�qS'䚱N�d��7�	�g�@�4-4sF���NW�z[�<Jh��G��%g$�_����
6v6X�uʝvJ����K	=0�|KW�!�		<4�`�� 'Y��H�fՔB��r�  �0�2�
F�_kPY��\.sdSC���g*��զ�@��z����2�*�J��ÌZa@E1t��7Nd�8ӵA޷g�N�����I��D@��A%��Qb��/�!;Պ�c�`b0oۧX�F5�ȲP^l��I%�p�����m�� Sq�$E2�|RM�8\�P��PB����"�O(,����9�R�\9O������'%P,t��k3+!��=}�uJR%B%��Ò�]�L��'>�ϻLr�q��Z_�^&>&�H�)�=�.� Ȓ/-�4}�"ދq�Fd�S���>����S��ēM���M�H�L �W�N�,9q��a��y ���ʄ�yq�lۢ���|���M-J�F0�7�N6-;e� ��61N�Y���1M�Xl�օ��b0^1(�ㅚ�T=����4o[�D;��D��i�f�z`fG�5�6Hj�C
Hl�X���|��q)gå2v��q d��gZ�(��Ä'3_�3qkO�PǶ�ǁR�L����3��4R�;�Z�h��pÌ��[�_����46Z���۹m��P��K�x�؁oD�����L ?��X*�<�W�71��b")�z���/k�O>��J*�h���I>M��y�{�D����{p)Q,XE�ԧ�1^�D�ڣj�ZN�[1g��j~.�%*�+<��eo��y)� �f��|b�սy����E�Z�93�)�Vţ���X�^h��'�AE��O�0�O�6+�b8ʵ�W-X�,�b�B�`h�B�]�|ц� 憊'I(��'F�k�:7�И��D�t�>������J
!'a^�`����]!��=�`IF?*��s�~�  c`�\̈��e�"u����T"O�  �X�dG%PѤ�@�oK�fq�PkD�I5F&�P���(:JU� �*m��� ��ˉl�.B�ɚ*v�0l��&�u��KU��tB䉈?ph�p����Y~N}����7'�`B��.524����+&��+�*�	!
�C�əI#n�"CE�$���P�L�C�	�,/� �,�2*�,r�l��:<FB�I.��Ũ�M��Q�����K�yBB�I�M$Ԥ�G��26�Q3�ˈx �B�	x ٣M� ���U��L'*B�,��h�l�
�0A��H>Y�B��%#ê�YG���Kn�K"S
�C�.l�ؓ�A�ђ<r׫�7[�C��2��)��!r@�[1��n �C�I��2 ��Kn쐒�'łB�	��y��LW�:�L�D�ȟ-7�C�	�Cr�!bw�l�$hb�H� mSbC�I5/����	g)�hH#�$�.B��8<�(�,��:Z��i���q�B䉌j�n�3�Z�n"�1��P\��C�?��ĹU�Q�g�h�� �Ca�C��X���ª��c�^I��L��C�	�ḫ�PN̂	uDBQ�Q�"�C�<
��y���*2��3/�B�	o*%��eͿv��xak�/qRC�	�d�PHy�M���#+��B�	�p�!�B�W��KeG�<��C䉽����!"�;Zz<��̂�i�tC䉻	Q�1�7M	((} �5A�2xۼC���ЗCP�n�:��r� 'b�B䉜"��a��*@Etbu��c�xB䉧!Fu���	*![��ѱ��>�DB�I�:���0"��a1��I®�!
.B�	"n(x��Y+��#D��zd�B�	8���r�ߢ�|�x$üe�C䉜`q�̀�a9�.��4%�2BC�I�7����"A"NJ�[7�
&(�B�	�iG4y�t�0,�^�Ҩ�,��B�I4V�=�Q�
�ewʀQjĥ_�TC�ɲ*��cT
��K��b�C�� �B�l7~+&@��xln�[֯ndB�I7qF�,ɳڌ
��"g��K�C�I�<j��d��<Hį-5l�C�ɺ`Z�K�G���5���	 '
�C䉣a���	�n���#�mNB�I�sA(�vΙ!;G��5@V*^��C�ɦV���XC�Ҕf�N5ӆ"�(ƸC�I dXz ,_ �\=���F&Jΰ��$C(Vͺx����>Aa�[̸豒 	$#j��1IUO�<YDH�(� �A�G�#��)���8�O)��/A�C| 2�a4��Е�bG�L�@���������ȓ 4.�A�L�!G�rm�R��r���#C��6�z�'�ܙ�4�>�3��H�X�c`�B(AN�]�vm�<���d�$z�,P0�cL&J�x ᨏ�[D����l��P>�x�DO��������?��H,�?z���jCnD�x�B	�7a�l���ǩ	&�yſi#̘Bģ�)@DWG%}�T$��'��\�W����ř�A��"�p�Or��cc��sO�%���h�ˏ�i�	O������� L48��c�K!�d�V�LE"r+>#b1����w%.) ɕ�&���0֣k�,i �bS V�HM*b;�1O����c��E�B]��ˆ�xxF�'�FU��F6zl�^tXs!P����Q� ÞDyFn��0Q��]^5�'�t1�%.�2C����e���RE�L<Y���j"f��)�&��Is�US�2��Bרl���r��P�!�@���e�	��RR�X]�Q�p�e��3!�?�
j�I��xs�ՆWd��aM�,S�|@�$
	�12TM ��]3�p�Z��GĦ�'Wf���f�� \�S)Ct4�[��r���k��Ŏ:�4Ygc�p�$#���]�7W"\iSk�8bx�5"�fU�m\X(���7�V�;��أBk\m���D�4P2|)�kT9a|��c1i� v��-�Jmqp��Ea�$��S3�JY��.}H'd	���GZXyv�QP̅%>/�D��ؘ{��<�&�&-�L��&m�����h�n��m�>�ț�s���ZP	.���0Q��U`��Uh�:^��u8�l0?9#P��ܺ�)���0��c�Ѱq�R�� �١$����e^L4��H&�@�:��C�w��K��Sy��:w�U;0oXId ����w��-ʂ\�z~���n��l��u����)P�������M���FJ_I��=Ң%�~ZힷQ��T��^= ��A8a��92fe1y��uCQ�U��3v�X��?�7@�_?�%Ɂ�`��=2.Oz�0���)"�Q��A��{�	!�� *{t�j�X�F���g���x���G+$��e�Q!D�{y��+ )||�D��v~�r�҈][� j��f7FB7��)R�2��%%�!T��˓Z�B��$B�*�F�26'��M`	�%C�^���L}�"�Z�mR���Q*䏕o������-f�(y�!�$C�Z7�C?�lm�eL�'	18u�d��@�b�������1�'R�p�Q"XE @L:���&��ϧ!�M��E���)��ݲ|ـe�G���cG��� ���KQ-
�\��y�Z<uw�(��ݾכ�aK�|����I��]B�xh�H�.[�@�c�0+���I ��R��I�o4-�B�;�3?�c��b$��0A��rr�T47�N=� ҟB6��N)$�NU[�K�j6�A����E��R*O4��D�C˾�9 �NW�Qb��҃7PL�al�����Y5I0�DJ��	���'0�>8ce�Dƴ��aŋ>]z��V�"�-��S����be+��`��k�>h��ɕx8��:���8�qc!���|���6���P��4X��UC�>?a�*m��m�VNH?
�.�x�F3ޙ��o���@h�s����V.�Jr ��"����;�O� 4�E5	.�߈�f�w��u}����Բhf}#��G~�WG߃O�R#0��7 +v0�t�2ovUC02�`���.I�h�T �ՅGmv�I�=�(��O,4r��̫����D�<���Â8b���UD/i��A�=?+��c�F��YN0��&��8'��"[�o�Ԉ��xRg��m�|��w%P�7�^�,K�@��7 �7H;DٓR�]�۸'��]d�L/R6�0���CЁ��>&�	�I�{˔l�D
�h.ȨP!�S�vÆ4�l�K���<�7,�H���Ƣ�>)����r}�1�V�B~2��G��hy�mF�X فt��U��\"f`�5Y�v�����J`��yE
̧f`Y��o۠^T�oY�1a����,\��4�ç1/2Q�3o�%AҰu��lٲ+�yI3��?�nmj��Z5̌��Ж7%"M�/���}��̙�(�Yͻ[�
�xf�̠Q���H���C4�����f]�c�� �<����[4��Rq�B�A8.�mp2i�	^�r���	�dp(f�^"�h�����)f���r�D�����өE-Q��z�i��*/Xj�ə�*�:bF*`�ܙ	�@�6H��It��**�bh���\�T`D�7�۝@�Ҥ�B�'��ћt�Dj�x��)b3�z�'�Ԁ�1�Ǎ2�Z�b��ڢr����̻Ld�8��E+g:�JG�޽H�NdB�1T�"D!@h�$�O��Òm�#��<pW��:r��=(�&�`�΁pJ�<���G	(C��oB�a�nH�$,�p�i�5��Q7,)p`YU�^=Fu��)�O>H�𤐂��ɀ�

�mtn��҂�,n�8�YÝ+�����G�(#䪖jә!;���"
�ns`أr�n�ɜ;D=���@_sf$ �R�|�#>���G�C��(�3�O� �J@J���?�b�J��֮ND��q��\�ց� ��P|Ŋ��	1A���U�]	
cay�Ϛ�!�a�|�Z9��Ƙ�y�!X�r�,��T�	�n�v�[��BG��y�@� ��f��ը!A
r��x#��Y�t��@)�)³_P�>)w�7#��=Z����S� <�A�
s�P�r ����A�vn͏^�nD�D�խ����]�j������ƕM�L����:��U��NL[�xl��+u�+M�?��`��RrZT!����� �V��˒j�놝���_ Zr�he9������X+l0�,��GX/b�|��h�$�����-�2K}��bv��<I���2�ɈKր�d��`�l�D��\�I�p �bt1:+]y3"���arP��,D$�	��B�7%<�#!��s(�Z���3? Qq3BS���E�'�3/�$!*$��kl�`{�D�Fs��b��FK<��vFO�s�F8`��D�Gw��MR��X�O@��(4��dmd`aO
�'��h �(ЌB�n$qֆF7���0"�IF��ȱ18���G�N˂j�=+�zӑm�W: ���K�'9���l�?/�j(�m�S2�#���:�|퐕!J�lm�K��F+��BV���[���f3R|��i�"K.e|��U�J8oj�c�ڙD.��j�Z� �q$J)n��
!Sْ�n_0�M�Q�
�m��Z�Lқ42��[��
�O������+�8�9�c?cg�4�A�@GТ"��a�%:��V=Ga�AD�ʠpu�@�Y�X����L?��M!dn�! ��'�l��ϓ��tJ�˻/�N �FK�~�*��@��$2\����LE m�L�wϒ8�ljJ9*�\�֡
�<�ЮY>��e�H��)8��ɑ��� `�[ӊ<�D�=�c� �P�	�s�����!�&	�0E
#M�䝈��~�u��J�$7�^��d/_�+���A��e�曫���s�#�?�,P��;3�ޘ���-�d�;�A$�!�h��n�`b��8$WP?�5���[�H�� C=t�:Y�S�߈a�h�$ ��6X�3���%8B���AT��`Å<p�.u��Ğ�e�b�	�O7��{��X�U�8�H�Cٸ��٘�i�|s3*�%js�׿��Cw�V32���F���-�-Otyc@��]��agEv"�aq.��4���v&x�����BaC@1�9�h��P!5�t��癷@x�� �N�c�=*��>@{�MCD�N
4�6�Q 5�`�S$g�5Gv��P�N��H��Ź��4� Ŝ���9@�a��zUZ����9H+	3@B y+%�ڭH���Ã�;�v�A��RC���I
70���m��GM;%�z�,MqFƖ9~Ҹ ��
6�����' �GD�q���,w�ўX�A�40`�Y ��n��1B�$<�,#�Gu¤�R`�XMP1�!�!f�|Pa�[���y�����I�wĴ��k�H˂H�m>U�v�@;s�v��[H!��(J<L[T��9q?t��e��i�����4a Ё3�Ǟ_N1��(>IQ@|{6 ]�"����A��[L(`GJ�S�.���O(���%�|��p�B�#��#>� �)A�yvJ��"BT�`�2ԓ�2m���''
*#D�8�B?\z1Æ)��zrN��b�
b�"�ӵ��O����f�u��G��3^i
��^kmN�Aۓ ���s#m��]��$���U*�5�H�Vڬ0�0�O*I�H�c�a��[!�(y��ʳ	T���ܴ|��'�"\�s,�n�HM���H!��	hfڡ��O��2M� �pkG �i��V�[4LjNx��Q_��3��#��A�ܴO]�!��T�#��"��I۴��'.���u�
� }�)Bz>�jaD�8�\fA�?G21�#8���{�pJT�ưҘO|�tRtG2V%ܜ`D%��P�e����$L�FI:!�B3DRRl�1���	,.A�d
T$1*<SE�?a���d�b.�[�O'�����g�M�ҥ16�>)����ݘf:��F&���m�"6�"�s̀-
���Y���0r1�l�p��Dj*ղ��ڜ'o�GC�zb(	����d�PH4ˑ)�8M�ŠpJ��ҵ�O* ���ФA�&A�dT@�g]&y��b�)�N�q��Ƅ_)D�BDɞ:~��}j�
M -�ēQ��ي��G5{Bޭ��ѣB<�+6��{lz\���]�=�j$�N0dH�����5xG΅�3� G6�Ę,zh(��W� ���I*��{��'�2H�X�A��,��p��)���ã�Ⱦb$�9��0x�IJ�H98R�ػ���v�~!Ч�%���Ӄe�?j6�iO>�f ��^=ll�d�L�T^2�"7
Q`��Z���Dh�n�D��� F�(���顪�Q�T	R䭁���2D�4����X9p��c�@�@�>i�l�v���'Yz%�p���l���.B�r|��3�֐�����+�6(��9Qn	��	^�|7�\�2���'�.&rp�1��=t6��フ[�hx 'e'�Ot|�Qg�2(*��w���TT��SX�K� �b�+{!��` �*9���
��3++�����P@���K�M�����1.@�Q�c��R��2
�')�ax"�ͫ�`�0@b�W�*i��k���*�pfd
q ��!Q�5I< s�bN:�x��/�
��p�>�H6R�r(�<�|�"_�+Dܐ�㨜%Œ�s��X:�����M�A7F�2s�N�+�ɘUw�����ph*=7C^��*��V����4��]A�`&l[�$E�:�LZhq�%�;<O4!��ꑫ^
%�F#�DQ����R�n���@��h9��!%]?H�$	�vJ�(T��#ۛB\���ĬSj��Be$��vU�80� ]%9O�*6�:�O�jdKF��{����V�T`�t@�6'cuɤ��w�LI�ŖN@Ts�fPJJ��g̀�R�@L�� �4#ee���(4X�q��ֱe��%r��y�axҪ�"��	#wo)2��k�-�w�]Cb74y��`UNH�Yk�A��' �|SSg�P�H�%F��~~�A{w�mX�И' "�c�_%l�~ɋ�JI't�	N��W�U;"�^Ȑ���ap\����-}�D�SB��8�hz�G�2��%�R	$���c���p����/�zU�񈉯�p=�7��uNd��SM�|%t0
�)�"{4$<j��*9B�t��BF!&��$�����pDv��y.` ����y2k��zݤ���B�,}x�����v�ўp+$�޷)�>������"�Ѕ/��)���D[�g���ӻI"n��,ʀ��-�Ve�ywv����?K¶<P�ߑh]�e�WG�|��5a�FK�:2AU�ޫm?pq��H��'i���3}�����C�P�⡚fC��y���Z1�ܶf�r�i \#oN8���G)�U#��t�)�f�R(�j�2�!�c�Q��e��/����V�1,����)��<	�eR��`p��J�[���(����VV29a�G�'"�����
t��C��H,v̳���?DE���M�=��TbF������	��Uء�NE��``�P�KC�U�QW	 \P��e� � u�d�^d�h�ĝZl�LYMHK�yȁ��%T^��U�� �e��%w|zD�D��?C����.���̉$�O����	ҿ?0��Ճ=�Tm�#	k�4�;A9�B	�s(Ն>7ޕ�ƨ�>:<��ӈT�;�JY��c�m���3�r�H�ӽiuڤ��(��(�1	��A�.��'͊�M�4;�jh�OoT�9�K��fy����G[�J:����f� ������4z���d�)d�-!�(4&d#ڞO1�ͩ&��'R��S��=�hP���5��{e��8��������j��>dZ����-M=�n 0(M# <��Kv�_�=��b��K�gH*q��/�@�V�#��ϫc���;��{�ޑ����}�X "g�^"btN��=ak,M+�F��;�>��4O�?�D�3vF7%c̸�̂;H���s�E<bj(yK2��>�,���X!;�F�+��vypB �0i�[���$�֜ˌy2��0'�¬��+�>"�����1G s���8M�*��)3L�u���:��`���]�ְjs���n�h���m5�j4�O�+6I�a�v�>��x��gޑ+�D_�Q9�:s�|��E81@�Q����&�.�+OǮi*F�k�ߒR�ӹx=rE#�b�'�h b�딚M;̬��(�U��8EgǡP�F�ᤣ�Oޕu��	Uy`4Z5��H1ތ����y��Zg�����?l.�l�h�یP����Z�ɳfB�l�z���-Xc��a%��k$�d��V�َX��A�P���R�F 8������0���E�=+�t0�)�j^t��yihYd�Iî
<X���d�/Y"�L��=-@��+c���!L��ʵ�:|ɨ��˘<1���3���,^ ���wl���C��	�%K��;�BC�~������D1C�pW��X�X>��k7BB7}������5^˒-�5#�:q.2�)#���l㖕2É/lU2Ȣ M�0�\��0�>Њ�eB��X�I��̶h圙2�ɂ/mT0̲0�����wD�I��*ע��ga@pCJ�y�`L&�6�j!͚�{�p�DE��%>	̻<U,�p���� d�; ��܃ÅS(N�e��Q)D�K�N�<T(�@��~��P�xAN0�����yi���"GP��ÀGIQ����i�& b4%J�|zuL ��Jĉ�.��FR���`�ș2���*k|	��C�$xp��h�/�_��i�2Ɩ�x:L@���d	I��x���߸��dyAȄ��d!vc�D���!���^�ypHΔf?
�X�Z��p���@u�(��G#T��ĸ���
WF����ДUEB|�HZ�M�%z����,qh�T)��G�m{"a[Ր&�Av�2`�u[� ���T)��<I��n�8�%Ėj��	Z�LXd�O��X�'�I��@�"aю0 p-h�{�G��Hg�>�nDF���7Lϖ ����ap�%��!Co��A�0�MKLN8%�4�>�O�d���4&q��äUk�Y��'l6\SB��<M��Z��(���G�? ���)�n��3$�(Uf��g%9q�0%yq�ֺ?B���$غx{�qBR�hOb�eR:D0�/9LM@!HSm��#��z�aD=<$����kJ�AXT���&�>��=���m���Ad�|-(q,B��yc��Q/y#~�1"O؍C�(״aA(-�Q�Ɓ`d�c�	�:t܅K��z��r-Ҍ8*�|#�B�=`�C�ɟQ��I��X&��凒<X��C�If���S��W*���uÑ7}�C䉩x��a�)͛;��x;�g	
�C�D��0a�]@zd�`�D8&��B�4!k��y�*�--��#A��U��B�ɊQ�TP7��+-���E.��wN�C�I<k;�����V8L�@A��	3�6B�V��;ei�.ņ��$���=�C�	U������J�d��|T���'|�B�I
���3�)S�}ٸ����(o�LB��5ZF��q�M#}�TP��"�<F��B��2�f�_'|��P'/ֲV��B�ɰM�n�#�/SK���O�1K�jB�	&[�Z��u�٥.o�h:�Jؐ
όB�I�8�e1�OO@I���򮝹j?�B�]o�2�d���5�T#A�~B䉆J8�1�\�H�p�Z��
C�I�F� �b��1�R��GB�^^XC�I
kT"����ór�b�K����C�I�.���b���-�xX�G§\��B�ɾz���cab��^�EJs�W`pRB�ɒ0�t��S0����#0�VB�ɢ]D��w�	K�!�HN�`B���ܤ����FiР+� FhB�I�}J�# j�ؼ���#.�^��W����Ha�gb�>���ŚzD� 'U�(Q@D*˧[MR�r���8�tZ-Ol1A1��0|�R�!�@DZFBJ�%B�! ��R(M��I�)��!��&K�Q?��K�Y]�jɄ�0��!��n�T���H'��q�,�l�)�'F��ak6��"s'4�)E �:�6ec�	]6fRh):gb3���:�~2��߈R~���THg]���˗�SY�'ϸH��s���h�e���h�K��y-�EO6�$��Nľ�b>��!N�X�$QJ��u\���7}�ȵH����y��^�JZ��s@%�!z�ȩ�Ҡ��<i���ȓ!Tf�j�VF	������d��g_���d��2�-"�M�e4�݇�J^�a"hL�bU�C�[^�(�ȓ=�8q�e��i��i�7/��;��U��`XP��cNƏ&}�-� �Z5(
�Ԇȓ設S ���.4a�-E����ȓ5�F��+�:��q&�Χ?�\�ȓD톄0�G�p�sF)F!q"����1��Ɉ�ɘ�Y�лi�8�x��E��ˢ-N;P/p)�e��=^6��ȓyN���D"�2:�dA���=x�h���g�L��ՅN'��5���*�1�ȓrXz� �A�J-@i`�*_�,`��_�");���Nئ\����:�8X�ȓI��:R�F�P<�䋑��#k��ąȓ^6%	M�?a�%��A��)��cd����ۃQ�@X���Y9�2��ȓn��K%���
����(*x�ȓY.\��$R�%y��ʀ���xPb��
ޝ
��}kj�
}�I��{�M��K�JL�R����Z���v�%��.�81B4��J̤oY�D�ȓg;z��� 7f&�J�I���Ї�s�����L�s�����W��݄�Ll`;E	�-�����Wb�U��S�? 6��f�5W�Z�{� Z+4(4ؙ "ODq����24�-t�W�K���H�"O�(��_�&��X0�´`����q"Op�K����P����a�����"O��(���k�8`�� h����@"O����2��q�f�ȝ)����"O2�K�G�D�9���έJs<P""O�|R#�ܬO�F-�.8e\m�3"O"���$��B��4���"O�� W�m�6 pn
�TЂ�"OP�2��>0�|�d _o}2Uɐ"O
zDХBi�� ő�4c��"O-#2�'e�Z8���	�yct��"O�q��AW�cU�� �o@PKV�С"OҠ3h��'�`���$]�d/܀��"O��J���&�h�s䂌x�X#3"O@�u�� [@I����>��U��"O�suoL���$�橗g��yU"O�s7aA�Z'R�A4K��3���p"O4]�.�/w�+I��7n�10�"OR�3F��1&IP�b��@�[WY�w"O��Q���0W�qpG�^"!���b�"OT�q�@ԙf�0�kkZ��"O,+P�ڝS 
��4-%&6]Q"O\�2�Q5H�P�Q"x0�"O�԰��G�R#.��fL�_ܪ��"O��B@-K�/���q��'3��9"O�A��J7O>.�Z��J=��u+V"O }0⥙2<cd<���Wm�diu"O%�fZ�K5P�t�̍b�����"O$�@�B0[R4�q��/h�>��"O��BU�дkY�@�E�ٙ8Ҹ$!�"O.���dՒIj��a
�D"O��vF��.�1�c%tq�$:0"ONĲ�	�L"���b�1J7�h�"O��ۑB)�ژr�a�( ,`�"O = ��D�!9p��d���8R͐R"O�y
 n�2&�{��X�f�qAS"Or(�$ѪY��`1A"��z!�M��"O��X�ț�M�\�$�
/lh"O4�s!I+	:��!�AH�0��{�"O�$(��_ >��݊�S'�X�r%"ONY�d�&c���k��oF�2�"O�8��)�1t�\x�5%H�M^�W"O�ք(��rǦT�`!0k%"Ov�S%�p�M���4#h��"O$���^�)���P�A��"O}{��m�z���ؾv�P5	7"O
���E9j���&�) n�p"O �s�Qd�f��P$D	�	!"O�]Sv�9�������-Ԑ�Y�"OD���VM V��q�C4�n�I4"O-0DIF�n�����=,���{�"O"����0	0v'<@�Hr"O4{e���t��=bW���@��j�"On0�PLθ!٤�X�'�/zr�+"OP�@�ؠ"f��TH�Z��"O�p8#�ٛ3�  ��o"�`I2B"O�9��vC&�{��E
#��ٚ "O�Lq����M��`���9|�[�"O�Z��?Jx���O�����`�h�{��N#G�����E��
�H��my����1z������$%�Ć�|�*�p�	��,t��f�]q" ��S�? ���<}&59���1�xHi�"Oz!��ܤK�v���m�?�B$�V"OXu��b���b�+R�U_�q1d"O��Xb)סr��pza��
vE\@��"O,� (T>u$t�A�bI��9"O(�� H�m�P=0�A�946d3�"O6y۳�G�}�@����v(�D��"O���@�d���Kb��#��"O�d�����<P�pvK�D��2"Oh�h��\:/���W�?�}��"Ot����:7t����B /ٸ��"O�ݪ!������*� k@͙@"OH�YR�:"_��5ώ�G
�4#"O:�#@�=�H��0�C)g�eXG"O�@��*m�]c��(��H�"O�d@��������dB������"O�����8�xH�'�E�JK���"O�!"�m�4LS�4�wl��"G�4Kb"O謁s&H�?]"���76J��T"O����Q)Y�Rhk���G2���F"OT�˧,ӴX�� #�X q0��K&"O\X�*�A%�X9��!l�y2"OZi�j�!&���kЄP�^�t&"O�I��N��d�S$Ӽk���"O���A�?_�2H#��ػ�*�2�"OD�3�I���Y���-_pr<��"O"и��éQv�E�E�Ik$a1"OphY�G_�w�J�+��� Xr��h�"O��k2�8��laS�""^�aI"O�㑈�""B��豊 YBRmS�"O�����	]`�E��,�"OR�X��b>~	;��C=Ny�ar"O��$�Na���� �  !T�]��"O4�1$M�޼x�a�-V:	�G"OH��u�Ue�^�8Fc^�L�ʦ"O0(����4(sD��8>;T��"O2��q"�'�����f��7�$�"O���6l.@��1�$�1/ -Qq"OyX�.ޓq��t�P�G�	zI��"OJ,�g�.%��QV
�%�"Oh;��ɳ]���F�Q�0�0�"O�(����s�8��� }�d9�"OPD��mX�c ���ƈ?�v���"Oz��j�%0���*�����%"OVSDؿrP<e:�Z%q�"O֐!4m�9Y��xb&bK"�.��"ON��go+T�4�6`����&"O��J̞n��`��!�06�~!�"O��AP&�ua3��,%�V"O"�p7�@���΃4q�p���"O6�j�GT1tĨ7�+D���p"Oht��M9T<n�XW�8{]d�"O���"��R��U�D0Z>�D"O6���g��]bZMr�"؅EG�i�"O~�VJ�����ͪJՄ��"O�� ����@�9Ҁūe���!"O�Zb�Y�~�8�CF�����v"OxA�5�ϦM�`�W[?~�
s"Ol]���=qJ�I���p��q�"OTU��сr��5�e�,|�8s"O~h�փ��s������N$�R"ONl{҃��}Q�N���1��"O���4+M0y� M�O�{ꄁ"On�H3bå_�@5�Fg�&�zI�s"O� ���a T>�(]F�F-Lg�DЂ"O�mucR�N3���dD�3ZL@"OR��.ӑ,���B��/�Nt��"O0���,@ ���k<��	V"OZ��T]�2(J1�°I��b�"Ot���N�I]̠�"��/��4P"O�Ya�䝡%�p+���
Ni�YQ"O��T�I#@�q2�6dd�)F"O]0%*̑A�9�aE�B��8(2"O.�{5�Z��T��fĠY�4�:g"O�|1�jv�[�&^�P��u+s"O&��E
��'"��`��&_���r"O��k&'BO�v�$���e"O*�h �R�E��q��!%��,U"O�5��Ϛ3�VL�� d�����"O�囒�Fv�@Sj����"O���4bٺ1��@_'��B"O�H��Ppy�`bC&2�ڠ-�y� �d��š��م!�s�n�r�'}�+ƎS����5�̠�(��'�ȸ)'%��Z�����M��i��,#�'��9� �&Sະ{�N4a��Q{�'�"yǥ	2����C�\����']]����V�����%� V���R�'�� ���ѲQ�� �C�:~���'۸x'��<�L�ccE�/Jn���'���!m�v���N�(��s�'��U�(��FpVE�R�Ѷv*N �
�'Qb�9��|t�"�ى���
�'��D3��Üxld�u┨d:Z�S�'t(8W��2ڴ$�3rN,��'զ�G��KgBd;/�!*�pA �'^�ؕOE[5���cܭ!�ؕ��'(DB��[c�hZfB�/M�<`��'�ʝ"�̋�E(j���P�����'�@$�!L�!&4���w��3	��2�':���$��?(zL������R�'AH
 ӤMS �9f$��|���'�zF��lt�0�Ą��t�����'Ɋ�C��1'Q�9�D��l]6e�'�4�s���=~J�C��$HZ�'~(�)s��%ErP[c���`��c�'x2�Q� �"�I�O�<[�����'p�Pd�5-�T��u#�(M��U!�'�$eكK�} ���᧐�p�u��'�"�J�)�WˎU��D��HX��'ְ���n�/2�.��"�W>/���'9l�S�@���)U�Ђ�L���'~�P�R��\uڥ�Ɖ��6�@�'���B�dI0s���;w䙽�(��'������B*D���E+O��q��'��0����<�����Aiz�"�'贡�H�j�����8&�$�	�'J21��]�.e� �s�W�.0��	�'>��J�A�Ug䀊 	Љ �>���'�{ע�z���;�O�nY��'jv`HSI������`�T���'iph���Ք5B68s׍��U��89�'f���Eߍ @0�Ɔ��9��Y�'�� ��Ǭ\��p���ҐG�:Y
�'��i�  ���   �  �  �  '  j*  �5  0A  �L  "X  hc  �m  6t  '  ��  ֍  2�  t�  ��  ��  t�  �  T�  ��  �  V�  ��  ��  )�  l�  ��  ��  =�  �  �	 F : ]! ^)  1 n7 �= �C �D  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr�	p>!��L�>P^�x�#\`yq�~�tD{���O(dG6â�ߘ<����F�N�B6��~�'.>I��]�(��d_�R>`��	&D��3$l��� ��'y��T"`/"�	�|az�H?X̴Y��ǘ^�B| �e �x�@�?	hlHG �*&���ɵ@�<A&��H�'�T)r��u����`��/T�i�'�S�č��F�P�+ 8x20��ĺ�y��Y8#N�P��1�P	�BL��'�)�s�Y�1~"AۇlX<�XAL<��8h�B��.z��s��N�@�}�'fvM$��E�d^� jSG�>l%��ρY7H03�,D�������b�]S�lZ�r�̹�'i��1�	��~=Xc@ѯMb����ėL��Մ��?�Ox��W���`�~�p�B��>eBV��H�Yw�^�]�*�x� �nN}��/!D�����^����b��WL����O�B���J�l�٧�QM�H�R�ϘB)&��$:��«z��u;!L��;-�Eaș!��5z�y���6G!���.Q��G{*��\�Ǭʓ��-W��S�ə�"O^���.ONA+F��6[� j���%|O0`� �B�v�ڍq�ڂ�x��i�ўʧ`.Z��y��V�k����=y����&j$�y���^9la��&^r�8Ql����)�O�yA�B��6-�Kd�+�j���yrj�8tE�Q���T�*�2����y� G�g�j)"q� �O>&ݚg��,�yb�D�#ˌa�E��^02}RgN���'|z#=%?�j�a�/>o��rw���b��}�S� D�DjF��$o�`t
�H��,�n��1�>��p<�R�� ��x�h�&RI�$��`�<)Ǡ]�S���C�g]wh(x�ԟ4*	�)�d�p篆%%Æa��*`��H��Es��:u��n+���ᑧ y���A�^89�`�<�0��%kwL1��9MV���&̟f��CƸǬ5�ȓ��q:��Ϭc����U�� ���԰�&]/+�d<sF��4�.��ȓ׀)��[�A���Ȕ!d�(U���Ҡ؄�P��3�ǶnO�B�I�'F!�6�@��$ZB*�!Q��B��7s���$�p��� !+ց?��B�IWL����C��sT� q� Եa�B�	�23���BK�8Uzuq1�S���C�)� j��Q/�9�1u�M�I��Xq4"O�����	_��K�	��7���"O��L kމ����-u��Z`�'A�p�<iڒA�Z��N@W���H�n�<�`kÌf(����B�"�j`�"��<Q왻Z���z�䛫b(h9`�@�v�<��4W�̅RQiQ2Ć�k��Ui�<yW!R#b�H%B�̟�`�.��M�<!@�s��@�B���$����L�<A�}��D���^F?�5�p�RK�<�3��-6�&�i&+��
��XGjAD�<��F�a�<:�B!|��aE��i�<��c]!ؼ,��&�06�ݱ��i�<10m���(C�I��8�	w/{�<�3n�'�$={a��;�\��3�	B�<a���zsҥ��F]5g��(i���v�<����~9zBd��W�.��!�o�<�擰a���N?W�t�e��f�<!4)��%9g��7iC���W�Z^�<Q7�'+�𛅏�6?:P��V�<Qt�t�T<Jb��Xd,�3"�k�<��a�?pY��Ht
�*T���Kt�Q�<Yv�H6�\xa P**�Hh#�n@T�<1�
ס�ΡS���)
ֆ�I�!�z�<AE���)4�1χ(U���p$_z�<iա@6��$�9V$0�q"�r�<Qt�]%L�4�2RF�]�jq�M�m�<�Se��\gX0���r�T$�6��p�<ɓ蝟Wp��2T�a��F�<ٖgE��(
@\��2G\�<ī�}ߖ�I�E�l�`�[PK�}�<�%��{�\t� ��>D��� w�<�c!H�Kھ|&�Up�!B�q%�C��CWx� �i���-���
�B�Lu�u�4�R�i��#Q.p�zB䉾^5k�)�T�p1�3L��>^B�	�U��a���=n(��3��i&B䉺k�����Īsx`y%o�'x��B䉦*I�ӁRZt��rD�<U5�B�I�Y�ș��#|�(
�� l�hB�	'���+ρ!AVy�N9}rhB�I5���۳Vm*�b�E~�B�I����U'Ѐh�^��-�B��_�Di:rcʸs�6DY�+T�O�C�ɩNQ$|2g��E��P�a�im�B�ɭQq����S�)���sE�9SzB�*�ع#́����;��â�NB�	&��
nLo��LXg�I2^B�	;����#�����e�KO�B�;i����55�R�Sd���xB�I�E+`�A��Z��h�'��C�I�q�Ґ����/~�Da#֬��0�rC�I-�H�(�ѾSJ�ҤJɂ$XrC�I	���w@�4�>0�BL�\�TC�ɚ@�B�� �� 1�I�K�)� B��T�@-�4OW?;7�ơCI�C䉄Bq�Abe"P�'&�	���	=fC�	3/&)9��]� (���Q�G�B�I;p�i�OӤ-�&��c��q�
C�I�4(��];y`�M`�/�8�B�I�o���3 �X�-"��G��C䉷s.`�B�S٦	9TΎ�8\B�Ie�θbu��:P0��'F7u�ZB䉃>Tb�"�ɏ%�P�āc6B�)� |��V'�4�H�P��-]�(U��"O^�3���h2j5�F��o�6hp"OL,�2��9<ct�AބM��A	�"O${)�+3�y��*��U�D8�"OJy���C�H�쨰1�
U��-��'���'�B�'��'���'���'�~�����|���ZW��tZ �'�R�'�R�'���'���'���'�jp�5*��I�x!�b�7<��'���'��'��'���'=B�'�xt �j	Amtp��@ИS8���'���'[��'��'3��'|��'���Eb֖_�x�b��ڠ-�b-Y�'[r�'TR�'���'��'���'UZ��)���pi�f�0,���'���'��'���'���'��'�\���A�SJ
hbB��,l��U�#�']��'�"�'���'b�'�2�'(�����{�f��D�;��'��'I��'��'���' ��'1�����^�p�l-X���}�Ty��'�"�' R�'fB�'y��'���'����F��
�1RN͏@�"+3�'pr�'���'TR�'2�'���'~&Y������ֿ�K"d'�'�b�'��'��'���'-��Y2c@6����P�y��tkS;5��'�b�'�"�'Z��'���'?�<�\-qD�ѕoSb�"&M3<W"�'���'��'���'�`6M�O,�J+"�I�F�]��9��L�I�*��'��T�b>�z����5H2�9+0�˩g%���R���J����O|0oy��|Γ�?)�&�$�<!ⱉíURȕ��Җ�?���{j���4��$j>a������<�N�IV၆"r-Q��F�.]�b�(�	ry��	p���w$̳+OH�����(3�@`�4^�,��<)��4�k��Ƒ:�.����®���Pg�ҡQh����O��I}���!�0��V<O� Y���>�<�2�%��B�� �5O��I��?!T@:��|J�{%> ��G(ƅZ3ƐC������D-����z!4扨-yx���'�[�p�h@�H�x�̍�?q�_����ޟ����D�2�T��#�	+!gZ���a��O^���!H����O9�?��g�O��È�^�	�#(��@t�pç�<Y,Ov��s����I�.|RL�<N��tb"Er���ݴGc(��'�b7�.�i>]�w�3iy��$jݵ=�����~�8�����	$vv�]o�D~�<�"!���_ۤ0 ��ʍ%.�aXW� O��8���'�T!��'6�i>��ǟ�����\�	�<�B�IԿ	����&З;��A�'�~6�F����$�OR�d�|���?9�B�,��òm,-h��VD�7M-�	Ɵ���w�i>��	��\8vƛ(J,p8�g�.�@���9��oZe~b�W5,"�h���?!6*��<	)O��*��{_�i�I��O�����O���O����O��D�<���i�V���'��鱓*	�{�N��':���kq�'��6�<���OD%�'�r�'�2�����f�:�f��Cd�_؉�B�i��O��M���s����߹K�S>�y��ʷYA�q���t�t�I����ԟ��ğ����Ń6A�䄃�eH�P݈I�UF��?9���?��i� ���_�,�ڴ��56��b�*ԴZ�I���0
w��AK>���?ͧ�(�ߴ������g$W�o��i��#g�1X$挞sD|�	�����O����O���^�L-��3��-t���� �O�V�1#E�l5�ʓN��ƈ@:��T�'���O�'��E��0��H	�hqDq@1	J�y��'��ꓙ?���OUR�Q#'�i2B��B���2�0Z�L�pFS#]���?1	f�'�t��I�4�	YW�MkoP#J="yx��m���h�	ßL�i>����8�'<7-.����	O�lu�EZ�{=���H�<����?),O��d�<)�Z�@��V"R� (��jW�N�����?�ԩ���M��'�����M���d	zo`��%śg.(�䭆KD�Ķ<��?Q���?���?a)��="#CU���D����\�T�C��I3��ߟ4��ɟ'?�I��Mϻd��ԩC�7v��Yxc�3[U<�J���?!O>�|*6Γ<�M��'o$�j4	E���(�pFV�tb-ڝ'�P�Q.�ӟ��P�|^��Sܟd8�nȉ@K����,ִ�,ږ�ß���ݟ4�	fyҠu���+�O8���O:d1�׿��Qb���	]��y*Ç"�������O����@���x����FBњ#l;?�4 �f���7瘝��'d��D��?1fO\�$�^���B��\H�c���?����?!��?َ�Ix>1C�
��7��}0��4C)V�J@+�O�n�}S�����<�4���y7d 7|-R��6oL�S���E�ɺ�y��'��'H��豰iU�i���	�?YÇK���HS�Ř|<��&�C��'x�	����I��t�I˟T��;4.X���']�:� W�ʳ":�'�,7���BT��$�O����b���<�'hԔ3<�"����Gla@�-��	�|�?�'�?���$z�M�m��U:FP�2�[�)M�Q���Dڜ�/O�4�dL��?Y6O�ON� !?O��M�R��m�4ga�x�3Naj����?���?���9q�=K*O<o�-y�d�S��� /N<'��}�B�eQ����M�O>���3��ן��	ߟ�!C%�L�� ]<>��� �e�	�el��<	�� ��JS�*��' �t��� ���g�#<Q(L3���=z�s8O|�D�O �d�O���O`�?Q�䬉�{D^Qk�f�8�R�9�䟤�I��|C�4���'�?y&�i��']�H����=?T:�	p�N�HR�|r�'��OQ��c�i��i�!�GI�!,⍹$@q������I�K�'��d����l���P]��07.ZU��uq��@�	ȟD�'C�7uD���O"���|27Cz5�8������@&&�T~¯�>A��?�O>�O�b�I�ˈ06�LRr�G5�İr�)�D~��p�@���4��89��I�L�Oz=����>���C�J�?P8��@��Ol�$�O����O1��˓D��v��m��QҦ���Ti����"�F��y�F�'���y�T⟐	�O���\��FTۥ�X�q�U��(��n��$�O�5�4�q�F�Ӻ�%����(�<ᷥK�
ͫ��A�]� ��FM�<�)Ot���O����O����O��'V�t�d��"�=�p��M�"ೡ�i��X;f�'b�'�Enzީ�uMS%'��Tcϯz��ɀ"�ڟT�	b�)�Ӣv_~�m�<�'��+cW�� d� N�ջD%�<9ve�
A>��P=�䓉�4���$��.���H�zc aQ������D�O����O���E.Q6:��8�I����8R� ؗ���K*�����	"��=�?�T����ߟ�$��x�g^1K�*���Y�r,"'�>)3�&VǞY F�x̧RƖ�D�8�?�!�����q%d��r�KlϦy���� ������D�O9ǂ�U95�5�;���2���\}�`uӦ�Yq��Od�DMƦ5�?�;���qJ��B�ͱVϗ ����?)��?q��1�M{�O��S���1�*"fҋX���P���8�$��f��)�$�O,��|���?	��?!�6�� 2� I��ƈS��6�\�*O~(n�Fmj���֟4�	@��.A>�a�c�����"�@́��80�T�d�	i��|����?)4�X�{ծG��>W���SFC 1pz|0UM����O�����k���O�ʓN�^8D!�, >��H��1p��?����?����|�.O*�n��u�d�I�y��@TM�z��9��J�7d���ܟD��sy��',��ӟ��iޡ��)"��5ȱ@��E����Yf@�B�iM��O����������<��'��R'pdF�&��|0t9���<	���?)���?����?�����V�P�pta˴V#t	��%�T�2�'2�r�$���:����զ]$������0��U9���f��7�4�	����'ߜ�e�iY����z����t~D�s�g���կ&���V�oy����#�Fpr��_2�ܭ�-N�u����4\�$(:��?���i[�=J0z�C�@Ж$���:��� ���O6��$��?A9��
?p������+N�a���#����0a�3\6�����Jş�h��|rE��-B��`B�%H��4đ�)��'oR�'Y���[��1۴?�N����3;R�Â�W.O��!��N�?���'�����
n}r�'Q�is+��t��ܸV�ŧP�,��'�ҏ;Y`�Ɛ��ʣ'�12�T�~
eY�zl�S�Y� ������<�/Od���O�$�O��d�Ot˧��X)��N�&��E�W�L-wٲ�(`�i}6�ۂV���	�?��HK۟���)�M�;Bs8$��ۃH��X��͑!v`L ��?�L>�'�?I�i����4�yb�32�9��Ȝ�@�<X�b����y������������O����3"P4Q�hĶ����B>�T�d�O\��O ʓa��b�b��'!M�^ަ���V"H��5/&��O�y�'^��'@�'f�f� [�� z�`��D!��O�q��E�{	6M/��	j����O4)x��\�V�TX�A�3R �"OTa�爑SBQ�PK3�zM@ ��O��	�0Ժ���Ob]o�\�Ӽ@�S�S��d#ׇ0	��q[���<9��?���#�� �4��$�2]��)��O�����iV�=��%C�Q<tJB�'d��y\�����?]�	���	��;�b\�h,M�0�ڏ`�&q�5�nyrBg�~a�&)�<�����I�Op��Y	�.g#�;�x�x���crʓ�?������|B��?�,ǵk��m[��#T�]��P%1�h9q�4���W�U����'*�'m�	
I�JQ�E���o��\@CҊ/�����Ɵ���џ��i>	�'r�6E�gAX��M�$	ri�T*�8[�^19G�T^��$U����?��]���IYy2� (} Y�r`�
RT*i�-,U�!��i��I��$)P�OS�<%?�]K������nb��i�:7"4�	^��  �g�63NQ�w�2y�V�;A�M����	Ɵ����'�����|BhW�M:���Óed�Ԋ��/6��'����4(ş}��v����h�w?��s2�&+�|��AY��x��O�O��?���?i��L�>�ʣ͔:bZ�av ҃G��1��?�)Ov)n��@A�	͟ �	b��5\	ئ�.+�>A�t�5��$x}r�'��|ʟX���Q�b�N��gT(Y����u�E����:wi߸}��i>�%�'�6�&����{� ��Sa�-\"��,W�t�I͟���b>m�'հ6��o�
10w�X2=HI��a�V�\c���O��$SǦ��?$Q���ɧ�M��CK�Z��,#���//� ���şpV&���'���҉��?���� �=)��A�72��#�O�����G8Oʓ�?���?��?�����	I?$=&����	/�MS���)��DoڣPF�a�'U����'C�6=��g
+/ 0Q"��2ު!薇�O0�D ��IލU��6�z�x g�+m5H��C�zV�9c��i������O����a�Qyb�'��]������~������>HFr�'���%���0�M�������?!��
{���%�?�|����?�/O���Y}r�'�O����� .�����3fϲ�1s<O6����V�F�ԌQ�Z���S<Y bFM���!宊�x%���E�ڵ��;��^Οp��ɟ����E���'��[��/�.5�aیr�AR�'uF7��+|�4�Y����4�h� +{�!BK�q�x�1OR���O��$?O�6�#?���Z;��)�� 
LH(V�M�A���b�J�,!�H�H>y-O���O8���O��D�O�����e`n]�q�]:�H���'�<��i�f��t�'d��'��Oerb�Y���҅K��O�<h�o�2<X��?�����ŞF�h�r���+�� �R�>!�Z������MS�O����^��~r�|_��re�N<�.py������N�����ӟ�	��Hy2�d�`�Ѵ��O,��gbQ�_zxh�γ1}H�aŢ�O6�n�M�@��	���'e��PR�ڗbȴ�bP�8� ���A0=�Ƙ�@ ,ϛo ��%�J���-��CJ�pb�����L<Se9[X�	ş(������Iğ���y��6�x6#ǯ�j$�@�˙�N��(O,����M�g>9����M{I>iR!�&y�
J�d��!޵�䓫?��|�Q�,�M#�O�T��玺�
��0gK� #�L�Q��D���#�'Z�'x�i>M�	�L�I���0PC�K� ��3d�y�a�	ǟ �'B����-�	ڟЕO� ���h�R]�����Б:�O� �'���'�ɧ���(w�2���F�.?����𯑷5�^�r����!$B7�Bgy�OU����P@Ԁ��/*c�i���'{��y��?����?��|���?�)O(�m�K��3/&u>��*f,Ђ
8���gf�ٟD����MH>��Y��	����)O?__�T���L3�ʌˤ�ٟ,���S�@o�<Q��>�	�?��'^~ V�Y;����q#I��9�'��͟��Iџ��I�	���Z{�a	�;I��(��']�7m;)1$���Ol�-�9O@�oz���n�f0�@�����x��k�ޟp��d�)�)%n��l��<�P��fcЅ��/1�[6��<q6FV�ZK���@8����d�O^�$���|�����^a"Q��,
�R�$��OX���O��^��)K<0���'b5S��� z_���E莕;b�O>��'c��'W�'	t2�%�^H�7�p8�]������ !7�|�rc>�	r�O�D�5-_$�3bo�,�:�z1�F�z!��ڠ<��X��ݰ@���+ɾDb����ş��7��O������?ͻ#�X����'?�xU�äz,�Γ�?���?1�cC-�M��OB�2)���d�<C���>V���AK֚B/�'��K�'R�ɋՂ� $\e��`�a��O �I�� ��OB�D$�ӝ�^h���Z�<��*ۭɶ���O~���Oj�O1��m��e��G��J��V�(�ޠ�0Јs��7�ky�ŕi�D�������$Ī���F���t��t-��@�`���O�d�Ond�3�r|�ʓ��i^�^%��>j���/��p��[��[1^b�m���D�<���Lg����0�'Ed8���Z�9ve�9J��(�7È$��f;O��$����X��<$����)���IF�s.�x%O�Q�r`��?I��?a��?a���O����F5["99s�ʇd	$�B�'���'��D߼��)��$��ѩO�c���8�d�W�Xɣ%��@�	�H�i>1�0��ѦY�' lt���B����O�c����d��g*���䓲�d�O��D�O��$J��������y!�G�=F ����OZ�Sڛ�Tl���'�rY>�Յݾ�©��֤b��)X*?��W�(�IΟ�'��  �|9�ӽ{�(�����dǂ� �ė�.�����A~�O,I�	��b���yR��M�=ZjI=vA.]��Z
96��'��'�ʟ��R0��<�"�i�M�EJ t,�Z(O΀���]��"�M;N>��'y�	Ο�Ò��p:pq��̊ �L���������Iw�vm��<a��|�Xt��?��'�j\���o�����Ə`���'��I����P�I��$��P����$1̵��� �����!2�7�� |Q�#���O��D�����O2��J��wΔz6O֖#���$ˊy��	��'sқ|�O��'h�P�5�i�����\�p�荒+x���PN��x��E
�� ���֓O���?��.��#�퍻O�=��D� A��?Y���?�,O0�oڈC����'Djȝ2 �����!�BT[�M �"��O�5�'@��'��'�Ʊ{���A�����K�O"���!�7�Ta�S�	F���O��FL�84��,��2��굉�O.�D�O�d�O��}���^dT�t�5���j֧�8!Y셊�W���\�Z��'��6�4�iޥ ���傑J +2h����q� �I����;M>nZt~2Ȋ<�i�g�? ��cr���.�� Jti�/$A� ��2�D�<����?����?���?�Ef֮:޾8y��%>V\I��\	��d즱���J۟��	ޟ0'?��I�w�`��EV+$@�`��
�,�O����O��O1��$;`�0/F�9�'�>��b�/F�Q�̈Q#h�<���>�H�� �䓒�䛣4�VD:�Ԭit��l�p{���?����?�'��D�릭R�J���c��E2���ʞ{`qP�e��0 ܴ��'듍?���?ٰh_1�hJ�C�	#-����eJ�um Q�ش��dK�>i((�	����:o"��*��ݳ�zX2w5O��D�O��D�O���O��?)"!� lt9��t+��; 'Kџ ��՟p �4^x`ͧ�?1��i�'ČuI��5j�y�V��
((|R�'��O�����iu�I1cs�9�͵J=��r�N�auJ8�a�ɠAc��6�$�<ͧ�?���?qQ�ڸ0�x�r�)M�9�6���?����$����agH�ԟ���\�O�h��$H���j����a�����ӭOn�D�O�O���yNp�@�_(bj�Q��^�DA��䄞mTU#� 3?ͧ5
��� &��e��ث��� $m���T�
�Ii�<����?����?)�Ş��ğ��q��$��"��ӑɌ��y�D�8 -�'�$6)�������OX�!��
2?Rx[f�S�l} ��ъ�OT��ƌ$f6:?Y��ďߞ�ryB�\q����܇#��۔u��d�<q���?���?Q���?�)�xM*�"���*�H� 5`���g�����$�埀�	۟�&?��ɞ�M�;P���a���QN�A�@��8~:���?9M>�|�5IE��M�'��m`F�8gL���
E�q�'ƈ�r����hQd�|�P��Ꟁ��"�j�f���B	I�:�Б��۟�����jC\Xy2,��`�aA���D�O�̐V䈅���o�`Z�W*�O���?	c\�����%�d��MȊ��x�g^����@Je���ɓ'%�jE ލ
�E�'M�������:��'v�!(���	�#�n	 ;�4A��'4�'�R�'c�>��I�p�NI`�C �x_T�14hRሐ��
�McQA�*��D�����?�;���?j}rd�7WI��̓�?q��?1f&��M��O�7]K��� =A�@<[S�	n���Xpkx�n�XN>Q(O��D�O��d�O��d�O]��lԵq������#��6�<1��id�\���'���'��O�үB+s�Ir%\RI�v��|�4��?I����Ş5<Dej��� rRPh�ca���x��f�8z�(�`-O
�2���?��<�d�<�(�3K�เ�E�͌ ��Ş��?���?���?�'���F���Qh�����D���r��C��|�Ta34N�̟`cش��'���?���?i��(2�!��i	���2M�>��)��4���������Ol�O��Fܷcr��礂�9���ӳ#A�y2�'|��'	��'A���U�y���ea̸��Ē���w�T���O��$O��h�Iv>9�	�M�K>)tEϵ:):�P�H��%~M��ia̓�?�*O��Z�yӮ�BW�\c�T�LX�B��.���l
�4D@�$լ�����O����O��d�)2� �E�I��<�f���*�����O�ʓF�v������'lBR>�h>z����b([4˪}D<?�wU�|�I��'������S�A<S��@�#IE�n��Y�q�+@�B��F�H/��4�*=3��&��Ox4uh��G�\Mi�̗�P��e9W.�OH�d�O�d�O1�F����ڪW�DqT�Z(0�(�s�ɭnl�s��'�Ҩ`ӄ�XR�OB�$�K�|@gK�pFN@Q��V�R���O�`��GkӦ�Ӻ�e��7��Ͽ<�$A��Mè��w�܄��u����<�,Ot�d�OH�d�O����O�˧>b�J���6x��:V�\� �iyj�ˀ�'V�')�OUr�q���<i�z��P�U�,�(�T��u�j���O\�O1�Dٺ�}��扨'9� ���ߐ),����ꖵ�l�I��Y���O>�O���?Y�0g��(��Q+\�J�V�����?	��?)OplZ}{|��ɟ���C��r�/PJ �b�)��.�ȴ�?i#U���	ʟ�&���F�4U�āѷ��q¨��B<?�/�`}���"G���'j��œ�?�3D�n��18�@	�J��S����?a��?q���?aI~�B[�|���$Z���'B����#�a>2M��Vg���T�>��'tb�'��I���7�ְ�AeX F���QI^0Di�	㟸�	��\����ϓ���L^5En�mM-+^! M4��U#���y*2�'�P�'�b�'=��'w2�'�b��\>zZ�j��QXT�KR��1�4=ތ����?����'�?!q��;Vn �R�;!?�)�v�ˏh������t�)�[Ov�p��� g%��*�[&kL�q�gP+7�"(�'C��0чޟ,�0�|�W��c�a!RO��B枥�������	������hyrhg�.��f�O~�dĜ9P.�Um�&f�*9�&7O�o�g��v�����T��ퟐ�r�XJ0����6d���{VnL3+�^%nZM~�ٲ1+�PF��w^\=�#μ3�Ԙ����JkBlj������(�	���	ğ���덺q�|�
���5�	ӱh)�?1���?��i�a(�O���h� �O���A�3;Iƌ������<(���*���O��4��Q�7&y�j�+��P� ��v���aWhUb��N�A�lp�͊��~ҟ|RU���	П���؟�*�&]	:C���3Ö�p�� �g��H��Ly�z�8��.�<�����^m�hjW��m���rW&Ǟq�ɸ��$�O���/��?��%搟b������iu/J�ZL��v �	��FA?	M>g/ �(�QDY�R�D|C��
��?���?q��?�|j,O�io�(c������4D�����BJ<�┥ΟH�I8�M���o�>���a$6��	��D����6�
H��?����M��Ond�Ǉ¼��O>�Y3���aT� �˟�V�
�'�������ܟ�IƟ�����ӽS|��oD6�Z�P��2J��4$j� ��?	����i�Ol�D�O�n�7�6C��5|�L�*rM�[A��d�O
�O�i�O��d�"R��7�}���# �2 ���C���(u�j�
b-g�,����$���6��<�'�?A"aG���%���ͣ|���A���?��?������������T��ٟ�"f M.h��W���J̾��j�o�\�I��	J��I�I+r�$�:�O
�n�j�V�I
U#S�M�d��4�Fg?�����<ː�\�����p\�	r���?����?��?�O5b�9E�'�K�2*v���q+��,�����z��$��yچ�<��iB�'(�w&&��dd@�D�0	�&ڳ�@j�'�R�'Y���]���3Ox�M�}	���'r�"44�H�ʩA�CX%v(ͣ�"���<ͧ�?y���?���?��̸E;� ��Dʆ١b��z����M;�eH�����O�"|�$�*M�0I �D�c��L�����D�O��i�ɧ�O1�9�BO'}��y�%i~���� �2}�\��O��(���?�t%2���<�Ջ"-�	�%H�i��\�(A��?q��?q���?ͧ��DW�+�V�@8`��"PN@��P@�}+2.�ğtz�4��'�@��?����?�"���;֦PQmB'?F�`,�:!��}8޴�����M��؟Ғ�����]�5{�-6�����!s���O4}����OH���O����O1�p����	 b� *p�T�S��MY�(�O����O.Uo92^I��П��Id�I/i���r�ߐTd��F�F�v��&���	������+C5o��<��^�8I9T�ڂY�r��C8��\xs,R�F��d:�����9O8�X&���[D4��c-��?u�M��ɿ�?��kП`�I��4�O$6 �U�� 4Flc6�ʞ8��O^��'wB�'7ɧ��UV�r�в�T�_�)p�Z# N^�`)Ίc46�Wly�O`T���k�܀��U�EF��UeF���EX��?����?Y�Ş��d���� E�r��jT�P$����%f8!�D���J�4��'�L��?y��4�����u���a.��?��X�F�!ڴ��dưPC<��Ot�	9�<Lb��ʬ+6�T�⡒=bz�,��L>턼Z�BJ %
iCg��/0��#�Ϧ?̴2c��3~BČ�SN�{��fC�x����4�z�@sA��v�$�ė<�P1Ѣ�A#:�#>i�O�5�P�a�h�"| 8�%ɏ:.M�X���8�~xbW��(J��xC�狊!� P!j�,`9p��ʈ0:e���G���G��iC����`�£Lh���T���8;��� Jr�jťːS)�)¢���\��ũX@�\a�b&dS�M�!zF0����T�j%�Ħ��ɟ���?՛�OD��Vc�	M�Zy`��F�:z�@�i<2�(`�'��'�3?��	�TH���@��]H��A�@պi�R�'��`\���d�O��	�\H���Ǣh%eHDJ�� ��}b��',I�')��'w�'Z�z�3�1-WK--��y�i��*[�-��ꓣ��Ox�Ok��lV� dED�l]t�)�@��	��3`t�l'���I����	qy"J�} &���	��$������m��M؇�>(O��d9���O��$�#ٖ��U/OZ؀��T<R� �[���O����O��ǂ�'>�^��h��M�Bu��c��$��(1C�i��柨%�h��柠��A�Y?�0��b �p'��yTtc�BG}�'JR�'�	
�f�#��"��-����-G|}��@&�	g8��n�ßh$����ß��$�R�	��a �T�a�,x��i���n�Ɵ���Ey��p��꧉?���bS�g�D�^�n9^IG [W���3�x�'��`E3{���|bן��hrI��W䩳gOƀ("�([�iL�`Wh
ٴ�?A��?1�')"�i��f��|&e�[�t�&��@eӮ�D�O�l
0�OȒO&�>�V�*X�AP�#T���(a�d�:�k6�����	���I�?Ѡ�O
�R������.�8�Qb	�+R ��i�x`z6�D(���Hh��>����ͅ�; ���'hٌ�M���?Y��c��)��]��'F��O���e�9���Ӆ=��ar�d���P�O����Ol�Ė�X�rh o��D���� ��{���mΟl��N����<�������p@߅T�nH�T
�pt�U���G}hʠCT�'�R�'uR]�	GZ��3K�7p�=��g%|6`��O�ʓ�?�O>q��?)"g� ��`�+�<Y,Ih��>�B�H>����?�����x��u�'"XK�=)�P���l�61-�~����?�H>����?�B� B}�A�C@�ِT��-�"q�p�ø����O���O��G�`���R?��I�CJ��;^�(�H0*�%�
�U�۴�?�J>���?1N�ĸ�� qe�T�d��K70�6@jǷi��'��ɹȈ�K|�����N��>����NЮQS��%�,�'\��'}��yZw$dYb��ĒC�ܸ 0���d��|۴���D�>4�(o���I�O��ITr~R%Ï|~$�CbL\$i���(�M�)O����Oa%>m%?7��Lz���Ŝ7v��0�*3��F�ü��6m�ON���O���NV�i>�`2MC|��8�"��U� ��P=�M����?�����S��'�b�7f��ш5��@�H����DE�6��O����O,���_�i>Y��k?q4D'2<�s�ؙT펙��iSڦ-�	F�ɭ�������a?Y��D=���Z;�]��$�ڦ}���{�T]�'��꧉�'�0�b�%b�@�㇛�p�p]�m'�$Ј$1Op�$�<��S�hm�SbN�e����c+״@:½���ɶ��$�O
��+�	�p���Z#팅y��l���T02�@lZ�'�Zb�l��Cy"�'*a��֟б��ǐ�	�(��"Ϛ��!�b�iir�'�O,�d�<a�����q�s�0w�dx���%�<�"�D�O���?y�����i�OZؙ!o�=�5�Ŋ��hJ������Ħi�?�����dP��'�Nx���(,`L`�v�1epvt�ش�?�����䚒u&lt&>���?��:'��1�ߦq���`���J�rO�˓�?1����<��*�������TRd�c҆!U���'�r+ܚ�R�'���'G�4Z��	��EKS$��y�|�Qb�5bY*6��O��oDR�DxJ|�s̖2gR�P�l�˨�z�,������,��ӟ����?՗��閲~���q��:yt��k�HE�3�x�'�(4X���I�On��7���<�>	�ã�Y�,����������8��t\�CO<�'�?���2θչ�"�=p�Z�Br�ƼT%d�k��i��'I�I ��)�|����~� �A�>�,Li�R%��۴�?IP,�����X�������ЊJwYD}3��ȁc$x�'�t�� ?)���?����䑎?��ݓ��^�/�j�c��:x���
}�	����H�IqyZw&^�BO7tC�-c��Ԇlm@�4�?�/O2���O���<��hD���i�#�`����> ����H�Q���韄�	����'�V>5�ɚK����U���dvb�#g���XUF�j�O~���O���?y�Q�����O�����V��8y�oڸi�Z�Qǫ
Ȧe�?����U�'���z���3!ײ��a�Ι�8��4�?�����kĈ��O�b�'��땧PX��UM��X�t@I��Ĩv���?	���?aa��<�N>��OVBB�޷ ����a՗�>�ڴ��ţ=���lZ� ������Ӂ����i* ��G�̸��D'�0ꢽi��'�ڔQ�'^�'�q���q@H ,�r$zJ�-�����i�X�
��q�d�d�O����0�'[�B��M��ۧa���Ǩ~!F��M��(��<�����:��ߟhE�����v�!x�$�A!��M+��?)��x�����X�ȕ'���O�8�1*�> n�(+O�m�`���i?�W�<peeo��'�?!����4`D�� T�r$�VpD�`�g�3�M���6�<�Y�Z��'�Y�S�w��a隭CW�J )�:e\	�'*@�'���'8B�'��X�dS���D�R��/;n4�R�G�l�  �Oh��?�(Oj���O���
�%��P�b��*,��N��)=��xw>O���?q���?�+O�S��E�|jUÄ�l�@Jք�`�d�'G����'��V����ԟ��ɰ����
e��������7,�� �ҍ�ߴ�?����?����ެc�X��O*"�Ǵ)1��ZFXҵ��^�d$�7�O�ʓ�?)���?-�����ܴ?��(���-O�(�l�;�oןL��By�&��b�v꧁?���C3m����GÆ�C�@�[�IƟ<�I��PZ�)s�x�Icy�Пle�V÷v�)��Iϝ��r�i���5#��Z�4�?���?y��"�i�U��"E�Dv�P��_C\H �d�R���O�2f<O����yb����J�@�C�/�5z��{���,s�F�K>z��7��O��$�O��	~}�T�����.d� Cݒ5�\�a���3�M{pJ��<a�����-����`�� )9�,H0e��;1���R��6�M#��?y����Z�H�'e�O$ͫ�@�#��℃ Q���i}�I͟D�%�~��'�?9���?��OȺ}�� v���6X�HӒ�B�^��F�'|^�9Vi�>�-O:�İ<����"�5��4��ˊ��T!���U[}"䗃�y�Z���ݟ���kyB����Ba��j�0��C������>Y(OX�D�<Q��?i�����f^ry�pk��z���Ҥ��</O����O<�$�<i!S�]N��ƀ)��-aP��8v�n$��	�yI��U�4�	Dy��'��'x8�R�'Y<A*
�7M!�qPr�P(W���r�{�B��O����OL˓|_�,yUX?��i��r���n��Hb�ju�
�Ѧ`tӸ��<����?���4͓��i�dQ�0��2)����ߗ7� ���4�?�����$K�_��]�Og��'��D���kj>��V�X\��yW��Hc�>!���?���
C����9O����o� ���ɃLa��QЬDn7�<��'�2~��'���';�ĩ�>��;�T�[�H�5`�h1�CϛV2�m�����u�l�	矤�'rq�� �A;�@��
��gG�CfD�
1�ifLͨG�pӄ���O@������'���/�f�e��0K]^�c8&�a�ܴo�&�ϓ�?/O�?��	�XF\� �^���K�-H�C* 8��4�?����?��bNz�	Ny��'%��̗�:(�L]�R��Т�*ߍPX��'���'~$�������Ot���O0�k�'�(s�n��U�J��KЦA���6��mɨO�ʓ�?A*O�������*�*�h��@���h��R�0��B}���	ܟ�	���Nyb���@X
.�C�><���BB�qg�>�,O����<���?)��k]{M(s��`%.�3n'��"��<)/O���Ov���<!����U����&<�(��cA�h���a�*��FQ����lyR�'��'a  ��'x$�R��E�����92$���`Ӯ���O��D�O�k zu �Z?��5$��	�+q�
Q�m3**��4�?�-O���O����_��$�|n�?r 8�F3h>*�Zw#Ly��6�O���<��L�M��͟��	�?�� ��7f��xE["�D�pB��)����O�$�Or=8�<OT��<!�O�`�Q�\�<!f9�gZtW��X�4���U�7�ޭoZ����	�\������t�w�����P�� �'�L`���i�B�'�R=c�'>�_���}�Ul�f��Փ�/Y�{$�A�R̦�X���M����?����zV_�ȗ'�01a	\<��%;E,�U��*a�!#W5O��ĥ<���t�'����+82L,��T<M��mr���p�D�O��DBa/F��'2��ܟ���j���H�+y��E�O�:P mnZ� �	���㒨l��'�?I��?)��k!ܽ��0k�.�ApDPk��v�'�I ��>�.OR���<����l�we�ݣ$,��P����a}BcW��y��'���'c"�'���(E��� M:��c� ����&� ��ē�?9�����?1�Kd@5�.)&�S$�V�3}< ("Y@��?����?�*O^}Y����|�d�uR)ISP�c�����n}��'�2�|��'�B�1u�D\>��͈�hܖ`F8a���-��	������'YX�Ғ�(�	��
��@3tPg%��~���irӘ�D$�d�O���F�i���5}�j�6��q	��S#kϔhP"���MK���?a,OT��[�ǟ��6L���,ĥ_9Vy�U�lw�II<����?ylN�<�L>��Ocbp8g��	V�9k�.�9��ش��d��^Ȍ�m������OV���\~A�,JD����L�>��p�[�M���?1獄�?AH>A���Ɯl���rLlR��C���M󵯚�OP���'���'�tf*�ɝlR���)o��}�&]�N#|���4F�Șϓ����O��@=�h��Q��'[��%`@D�=��6m�OH���O�q:�gY�I���\?)vM�/�H�(e�(Ʀha�.[Ҧ�$��X��x��?���?�1�I!Za��
���_��͸U�#u3��'�Ęp�4��O���*���Fp���06V�@aL�6���k�Q�X���g���'s��'�O�̥��C�*��ƈ��)"$@_5N�D�H<y��?�H>q���?�V剁ri�A��ܦ745�w� -}P �����O*���OT�����7���b̑ (�0 ��Ɉc(���W�T���X'�P���h��w�� �']��]!�����6�Z=��L�'P��'��U�|+���ħ�V�)�˜�t.u!J�_@�a�i��|��'��J0v!қ>��(շ��5H_�s]Z�ٴL��M����?)O)��(w�Sٟ�s�� eI�=0��D�AB�c0]0d�3��Fy��'��O뮜#6bAᘳ]< �0�	
��v�')"k�6��'B��'��DR���{���ӗ)�jl~ِ��|<:7��O0�K��DxJ|�%d[KFT���u�hbƞ�=9T@	8�M���?����BQU�(�O�z0Q���-!���ɓ�K��H�Gq���d7��䓺?�BK�#Y���zd̆�K�rtK4�P!��v�'��I:JѸ@�'��	� �<��ak��I�+�m���U:�I�ħ�?����?9�-� Ҡ��ě!I�N%�1- �{K�V�'��):X��[��6�2�$&Ύ��so��05���䇜,/b�'���f&0?���?������B�)[��b��-C��a ��)H-j�ӣ�Wn��T�I��?���k ,|��d@�d���1��I���<�<9��?	��?A�O
6pH�O3��ϸ�	��ҧ6i�[۴�?	��?yL>�����%f���L�o&E�T�CW�(�R�Y	��$�Od���OH�>jM|��oN�B��Α,|��<
3jZ?U��F�'Q�'�R�'ɾ-��}Rܔ$\��ZR��,axn�Y1Z��MC���?��O"��K)��O��iH#��e0oׄ8��HR�	�&��Iӟ����>���FU	Qߐ���b�lޙ7N��M#�O"1pG%|�е�O6��O���O��Ӆ��� ��c���] ޔm�������G�\#<���'IJ�Ur�B˳J�X���?р�߉�M����?������x�' (�3����xq1�
A.*����+hӚt;q�)�'�?	�A�#wMX�bq�A3��E*3����F�'-R�'E���1���OH����x���h*�DAb�X�M���o$�I�|�c�X�����I΀ ��T*�9R��'��&�hp��i�2�[�~�c���IG�i���=����Qm��:�u���>!�aWP̓�?����?��O��h�n<�<�Cv�Y�3�h�K]6�c�`�IA��ğd�I4}�l�ڧ�?
�}ӵ�W���%xf�8�I^���b�˚#F^�E�to���Xs1�^�()��"(ͱ�y�`�>S�&%H � �@�k�����'���S��ێ[汪����wW&( Ek�>������.͎$H�	��'�(�8�
@9l��mJ��ȹ����	!�a�DX%:�^�	2����i�S|Q�%BkGkH���wq(����'dc0�gV�m�A�Wй=��25i��=�m(S���P�e�3E�_��Z��7H��Ct�
 K6��rWʉ- ������?1d��C�@XrÌ	?&z�k���wYJ�S@���ۘLl"L�ԥKۈ�*�����	<|�d��V��'���شr>`�V��^���`��uĆ�l���P%1�>q���'��iIs�'h2��џ,Q�7r���!�
ʐNN袃 5D�����"�D��c��)m7 "3.O��FzB�n3DAb!jôOB<܃3��?���'E��'yb$8B-N��"�'~���y7�M�&�cuʚIhDc�T 3-�X��IN�bYn���/|y��3"�|�o�y�*}��2�y�q*�3y��l��ޜ���dR�#������L>ņ�x֢Kb�	O>L�'b��?�Or� ���4퉖=J���;8�AR�_>�\B�ɼ#�J� L��4"��4GJ�%đ��'����0��j��M�,
�d�Ʈ.Ey<Q+��+H�����OF���O��;�?!����DH��(��t����)F���pfʹ]����1F?>�\�k'�'lOF}I�/D�YgM��`�,jf4d��꒔,������܌?m:I��I>������jZ����*�$��O|�d9ړ��'�N !�,2{��`<S�<��	�'/��fͯ7���f��0��y��>�)O��
��]}��'[�А�πRZ��Q& R�	��!��'j"�!e��'a�	�h+N�S��^#/����F �h2�쉯GA2(�2�ý+����I&�̹��.F%�l,j�'@�9��F�C� ��kZ�n����Ǔ2Q���t�'��1n�� w�LP�D�$6UZ�ҋy��'
$�˳�d�fxa�0�*��'��7�K�u1 ���OSS堬�"�>V�$�<I�M��A5���'��\>�R��
ԟ�*���13G�p��o��z�ퟜ�I�  �9��4������#��WՂ�s"�͏��)�N!}� ��(y ��A�-]��s�-�D �e�J~��&mY��P��2�Y��B��Իecb�'�7m�O&�?$k�+�c���/1����kd��'��V����C�p8��M�'��9*�����p����޴�?���i��k[4<�óC_�?���у ��듌?q�IR ���?����?�׿k����5tV����E�直Q��S�A�>�5��

��1�|&�|�l�nຐ"t�^�:����,"���X���#���W�q��'�$���c�VY�E�R��p�U�'"�ɭq�N�4�,�=їm� �T���N;b� ���m�<�F�E�?�i@W`[�$��\hQ �h~rA?�S�$V��3U&X�K��AX�G�	/����i0���j`��ǟ��I��@�	:�u'�'0�;���2���6KK��k	_�GT:�jC+��U� �FB5�O�L�5��^���m�?#$-Â*ƠKq����&'�O���7Q!e��T�͕+��q�Vt�"�'���'��I����?B����\���F鼹P!nO�<�"�_!]ߘ5�e��
x�X@���P̓��uy'G�:ꓥ?a��\�a�b�1�}H$ʴ�?A�Z�9����?��O^�|�&��*W�I���>A�mZ#4�G')$ l�S�#O�1q7���l�\�h�u?QѭʳTS�����s�[�N�I8�P9���Ob�$�<�c��bъ��'(�����p~̓��=��HS�}�v��a盺u�����	v<�i��`���48�H�����3YT��*�'��	,ƞY�O����|"�I��?IgH^��8�-ڈ@(���-�?��y�dE!� �.�S���*���'y��Ce�_)І�_�ft�@�O���S�\�^�$����I�#}�ꎗN�xs�m]3W�(1CQc��f��'��>U�	�h�
	��	�~�R�ԧ���0�Ɠ�% ��E`�Q!�T������HO� 1�����Y%W�V5�)�ĦU���<�I�kgbAUm��I����	��u��*
Lر*O�7t]Y�S1O��8��'��,*G, ZF�T�S 4��{�-����<���XO$��e-�C[�����<ܘ'\����S�g�'����AI� ���\��C�)� P���C�ܠP�l��������Z����n}P�&�N����8���x-�$8��?v�h�Iݟ�IƟ�^wV��'"�H�gG�x(Wܢ���R	C�̂#OD��4�Q�J�t��TC�u�� V�	�0!�тJ�:��hۑC,�40g� ���y:��'&�';��'*�O�a�.	-��q���s�B�"O�@+W.H ��Ӂ�Ra�P`D�d�x}��i>y;�ϩ!�B J���7�VqZd/:D����Y��5ؑ�ӑH~l {�6D��x�@V�S<d�K��̄1�^�(1g:D��Y�	+
�]k�I�*@ST,9D�4c�oV$ @���C�h�ay��8D��0`�_(v~<5pA�6lܙ�s 6D�Hڔ	Z�4��0aߑ
��A��6D����,`<��I] `��!��(D������>g	 I�)��t��IU 'D�ț���4����Y�d�($D�\���G����9��\�����"D�\"��1$Iu2uDC"lD��b�l%D��!��M��Xi�'p�Y@V� D� 0Eb�>s 51#�*�$Y�d�9D�@a����#�|���T�l�H-���)D�p`��>�`�; m�U���[��2D�X�U�C�Dp�Q��M�f��͐��2D��ᄅƷ|�>��D�K� ]��Zrh6D�4 ��N�}�2	�H2��H�3D� *��h�Xd{���1Ί9u*2D�� ���;Z�Y����~U���0D��1��L�g�@] �IŤgXI�4�"D��ꅨI�M QTK�.Dm�Պ�"4D�l�sdōjnBa���o|,��k0D�,BQ�
r*��(���-����,D�|��
�/o4����`��� e*D�HK�)�T ]sF�R��إ�)D��t�Q�v�ֈA��D6.��e��&D� ����r��P�G����Ub�2D���IN[Ґ)�sJ�\�8`/D�(�0��E��#'�F���,x�(D��iӭ�=��3s��i~�4�4D����C1`($aE)"l�|Xx�#3D�(�do��B/����^.��3p�$D����N�;py�-��a��h��ms!�!D���u��!n����O� z��)SQ	 D�`
��V��a�p�!m"��;1E>D�D���Ä.jRģVc�'`v�ӧ=D����bB�4S��q�EL.1n��$?D����Yp�x��y���i�e
$�y' 7�yp��Q:p�����`C��y"�ӊ1�x�9����U��D��S?�y7 Q4�� �O�n�QR`��yB���N�n��S%�Tx<%����yR��#㮉*3�ղҽ32�U��yR��6Gnޭ���v6^���C��y2`̝W2�p�U�@"Œ� 啱�ybl<,!�,B�ۊk� �˵n�"�yB�E	1cx�� ��c���2&"ʅ�yBgQ�4�(�`�&ۑ\�]ؕ'K;�yҠ�.FJ|Z�M�O�\U	_��y(M�?l�t"���@�ɹ�(G��y�(Y&��9be��Ѝ$+��yr�R5 :��FA�C���x��G�y�b�&T�{�DĮ?dP�Wϣ�yb��o��aI��	�I�&e�!��;�yN$F�3�U#F� �R��y
� ���3�O�g�<k��G12@��"O~E:d$FZ���K�O� ��H�"O��Iah�����w�@41�HD��"O�(H�A�D!"��e��O��tQ`"O�X�W/�./$=����k�t��t"O��)�P5>�$T�O�7���q"O�1Ru�W(��!�md|e�"O����#�!��,�TcvPA�"O��(�J�U[XQ��D�z@��[�>A"l�D��Ho9��i�?��rv�<#�L�|�T���ϊuj�����-����s�OM�L����|h�b�\��4AԌۄ	�N�"~nZ*�D4@C'�p� 5��3��>1�HE�<$@1��4Ě�S��B�jU��:��)����+yrߓI�dX�K0P��� ��Y��`��[���Z�+��S��$�a�G�-�Y·���L��l(]"��yǬ=D�xK����p����@����zRF;}�@�L=2]qu��/�v5�FP����~�����
T�<���8�H�h��ҵ*ߑCXa�s�ص$�ک��-���U�ֈ�}/�|	f��_��,O��z�-(�s����V�\PU*¬V�r������	�f�(��Sb=:����A�E�A�=�X��Bم+r�X��ÊŗPJ.]�D�S8�xkR�
e�t5��-�;��{�A��&��aSrGGc?�OԱ�?��t��k��4jj��C�J&C R!����frh�������O J�$�#+˘ȣ%>�Zu��Ò	��5��Z����\�~����H3A�V���Sސ�g�$-�}�%�
?p�2�i[`�� kPcO���'h�!iTk_�J������S�4�S�O�8c%��j<�qe��Ǝ��F��!r�Ȍ��g'���:��QCn~+8�1�`-#��D��=��y#'k ��1�#�_$��g22�Ce� ��9��FB�0V�lt`d_ 	��H1]w �	:!��F1�2'�W5��h�'����a3m�RHrQ��V��8���U 2 "F�Ƅ)'T����1l$���)Ψ���)B�Ȱ+ L�H���VD�>Do6�8�H�h@ "�Ȏ<!ń�A�n#ړM��!!J%PH)�;<x|�f�J�+�F@;���?&���O�Af.D���C�p��c
A�g?�5�>|�z�#☗rH1jQ�i�$0Q�3�ɦ)u$1 U���}��x�%��V�.�C�� �Fϖ}@���H�(r�f�I��<,tlؕL̴�#�OX�ڴ#�t��hCb�,��C�'m v+��8,͉�Eɕv�ny���! 7���Ǌ��xޔ]kK<Q��Y�<)���=�~r`��F��k�'r��4��c��~rHM!xY����A�^��	9�J@���4�:�7&��2��C�Oֶ�	�E2>�NO,m�
ЛD<Н��@:�{�p�d-4�p��3��6�teH��VBA�
֝9k��<�ƽy��iAG漫n�';}� Y�$!�9Yp(T�
��y�I>Yr,\H�OK��I�������&��a#\!a�.,:�yb+L!.-8` �*�`@�`�И'�v	�f��&�L!�� -Εp�4!���ێ}2C�gl��ja�-h��i�t���';�MH��IC��(à��}Y�P�rظT,�52�g�Lz ۓmU��p7G�7J�	Ӗ@��?�t�JrF��pp�@��@B��;��G�sR��'��hI����<k4٩��%qaj0ZT#E��yb��'jgX�B�A�&����rE�%,6�|�r�E	$���!�+��'��#�k�\��w&�y�Vhγp�L����а5X�q��7���c�
�B5(�V"oX9��a�~��c�8��i�'>��*P�B hd"��%扶o�acA�� ��L3w��"'`,�>�B�
Rl�B� �3�,p΂�/��T���	,�v�V�(���ӧO(:����a�^p`�V�,LO�"׭��F3D�1Ea���;�']�9+�K?�v�*ufK�sM� ӭ���D�3A��_7Uj ���)��X���@���-d!��C�8�A�)#z��ʣe���na2@��:T�P�r"�ά8R1OP�p&�ތx�&yx�4�):��[+����X� �P��'�D��"��,�@���X�\�:�٤'�X�x��<٠/�5Ux��tT�j͎t�q��̓>ER-2��>A�|�wfA5U⼄D|үY�A�vԙ#�̵/{�-��B��P���Xd	��TҒ1�࣋{y�i;!jݕt�XI!%	#I��鳓/���?I�������x��) ��9�>hI$��s}���b� Vxx��'瓶2�@9��O��C�|̓�޹j�mY�/@@�ɖ��G��q���fX�T�?E���D5�H���@Q�2rHIVC�A�NUAE��)��)��i>咖���e�杞dG<{���.O1���C-Q|���[;<�B���� H����c��d���T�'�hi
�*6�'44�p��Dh�j-K�$"<�AS>�DU�8�h��Cl(�zT�a�?�T����D�Q�C��8LЎ���-҈��i� X����hD�0�GefI!��!L$����9`����̧^�� �L�0�L��V�{H�}��?��?�����Q��=`�g�n̪��DdD��@ 6ҼD��@y���1��� Ԕ}KR�{�� �7_i���<@b@L��)� �,I�dC&w�v�a�A��,�5@D�ɴe��m����0鑗��F�M�����6�U���csÂ�ÈB䉲F��ɰ��Y#L�0X`D��z�d��-vL`@��R�(�)#KI�)rd�}Zt�R�t�0t�g��Y�$I�v��}�<9���|Zd ����r�lX��ώ�1ʣM����H��		���fhSp�n��D��J���T�C.J�"��-�.Ȉ���v�h�H�D�O�f��6ᒬH��9c��Fi��t�e�5S�rlZ�/_4f2�ʀ� �\����6犉#�6�ۓ':s�Td��:X��]cTe���	�)d~��"O�aL;8�:ɘs�ўD6F8�`�i���b۠��s�/��Q�(�Af�(�k�\�����	lD�x�"��N!�5B�DEI�mҶTO��K��Li�
X!pGD��lI�,��4Ε�BT?��2�d;����G��҈Z���(�z��קt"0���Yl�Z�,N�tP��̊Z��#�.C�u��P��L^'%�έ�ߓF�q�ś0�^��
L�8���<��\�?��ݹe�
�}pP�7�P��O����J�/P�9sU��]@8XS�'6�d��%c�\p�uc��S�si�6�X0R���ȈL�����)�<���ǡ�)\T9��l�<3��4�s"O��6GU8[;@��t�3 � )�PG�9m{D��1ݙW�8T�L���2OE��㟼���S���qT�J�3���C�*LO�9�u-ù�⍣D�M�g]\�)#ɦmm�����[#n�+�����M�R.�<:7���ɺr�Hag��j[^�#%�b��+\��X%�ݠT��)���,.�p�� ȸ�u���=\tw��6!D�124%�+�y��G��X�%� [L������P�r�M_�5�I�͔�n�,�B�C䒟<�Z�w[�`6F��
�x�)a� �1��'?�dB�/�+�Bt��˛�/��"pI7�9�!%���͘%���<���Ѝ\A���ԓWo9�$�@��$!��ͫg�N1�'���	��W%+@Z ��������'f2 ����K>:���#ɂ9z���y�/Ѳx����a*@�OU�(�̈́_J˖C,���A�'t4�&��}��7M	/ Z�� PM^1���O4���3?i��]�J9.$Ar,؏d�� 0��v�<ၤ9f������ʀ̊�Ѧ~��� �`A�i>.���I�j��g���)�KX(eF�ի�n>&�P,� C���Z/�!���:"�����6B�5H�`�!�ս!�^=B�Ɣ3 Kb�<A�ʍD��Y���0v�E�	�.m��C�0B�B�	�,'1I#��.Ű�cr�EI�8����	�Tr�fR�PG��OPK`gԷG8�����E�,)�5�Q"O,䊒F��
o���+R�\+T�[Q�Z�H�t٩��U�p>ѳ������V����#C�j���k'�0.�~��vS����l�3jv�d�>W�!�S"O,ݳv�D���<0U!M!2�av�$U6A�bp�����&��a�B9Otҥ2���?R	��"O6Ti����v��'�
�s�:<(�g[�&�h%�<+��<�R�Άv�X\ '�O(P_�1�TFe�<�hQ�T�� ��K�!SU�5���i�<qp搼�yq�@�
%��w(Bi�<)B&[OP��O��$^<B�J�I�<)�N�S� "Ąu
(3e�z�<aeI�4��q�E߂=�0��*�o�<�5�ώ	�VM3�CQ�6)PX�g�\i�<��(P����B�:a��jš P�<�6*J�t@<��%�H�0�atv�<ٖ@!�29����1T���c	o�<�$�Y�9���c�,1%�q���`�<��#cI�1)�D�'=�r���)XY�<��Γ$�n��ώ�4���K&�S`�<ar�P��vd�� [�
�� 4�B�<	�M� kO��(��H�
�svc�@�<ѣ�P($�b��"aғD ���{�<9E�̑
�px�-Г6`�	!�,T^�<9��s~�/Y�:!��̈́��B䉝V����Ч)>�l��H�a��B�)� ��#`���Q��9�� @/%輪W"OF�S!@�FnJ�f�Ɔl��"O����e-�K�'�]��"Ob�2A�Y�]6z�
h��S���t"O����G^�C�,�tǍ wXR��`"O�@zj
j���¤8C�T��"O��Ұٟ2�Ƚ��C�;=�"O��!C�Wm6aR3C[<= ����"OdQ��-�'���qL��7/b�b�"O��Ђ�]�6,���E��bs
�J�"O�H����hQ2(Sԅ�䖪)�f"O�zҌԉ'����+-v�6��D"OB�S�$@�nH4��+�Z[��;#"O�����;n\%jĈQ�uf���"O`�D� ��ɣ�0K~|��`"O�R��09zBe8�G�S�*xj�"O���O&}�%�FeX()R���"O�����>T? ք�,
�v\�t"O��A��6��a"%�$����"OR�c�Se�,I��T�V�ll��"Oxp�kQ?^��Pp]}ڼ�y�"Or ;��U�e�%�߬|�\tP�"O"D0��eP��2��YƠ�S"Oݳe����<��o���z���"O�QC����
�x���D$f{�!�t"O|�5&��\W�!p#d��;��Ua"O��[�#n�~����:��lCe"O�P�J�d��P�R�_�\ �"O*�xX���*R<y&~ �"O�����W�쩃�hD�m>
��"O4�p�P2>]��3�}��I�"OR�!�lY�$۬�6��:�� �"O��񅫎�6~�i�!�D�6>q@B"OF��ń]�J���ɤ�J�&�܅��"O�hA���r_*��@ Px�� F"ORD�G/�<P>��� hZɛ�"OXHy� дHaO�4F�h�"O<�p %�$%ʹȑ�d\F�-��"O 偅���D�95��-�Up�'�!9�Q�W��!V�e�\x�'��\+��V�\І�VY	0���'7�5��FZ`�_.Tj|@
�'Q����e=3�H{PN�\�C
�'1L��5��r~�H`FB�[�����'N]P$た\�
0Ii�P��b�'��Ñ�F2|1gН1<�|�+O6���J�!�:�`��<dKUꛐR�!�A_��Ԉ�.�.������6,�!�$]�ty88��N;|����ʧ�!�d�4wYhIaD[7?>����3�!���L�d��4�C( �H�ek�]�!�dB�M� �
S<�Ы�* !���I��	�J��)+�(p�I�F=!��<R��u� H�l�=(3h�J!����q�6+#m�� ؠ䙏x!�$F"*�D�b����N�\i���Y2�!��bI8�IeL��N�l�Z�� �!��9��@0C)F�:� o�!�$��:�@�P"�_~5" ���O�!򤑂J�b��&+	�q�nP��Щ�!��R���!e�c�88JdGQ!M!���G@^M������(�H�*g�!�DD�E"��	�nzLtP�(�Y'!�D�P��5��ŉ�bg�Ⱥ��L!�� 0�ui�"z !��Ε�{>EI�"O�P�0���;3&H3V��.xul���"O�Ds��M�4�Z٨�N��ogT|��"OȘ��.H��|���,Ua:���"OLy����k01�`���DU�q��"O,-��"F<c��܈�d�>'�J�R"O����
)�1�c-R�9� H�@"O�]�k��i�~�ƍ��W�����"O�XQ���������R����"O8����J8t��
X�xz��D"O`��bO	S�t@U'"rfV�R"O��S�aL� 2�E�.xF�e�"O0`�Ǐ�.q]�rC
SH`=B�"O�\#0 ��:�*����E�>4���L���X�ue��jp&#��H����!�!�䗱8ɪ�c�.\p���1 	9!�$
�B&9���N�R�� �0e)!��;N=}���8@n2%R��O5U!�$O@y���(Z-_�arUa�8^��φ �|��ߩ~S�K��1�B��>ctY�흊4��M��"ȩ'Y�B䉒_>�[��P5%���@s(�q	�B�	%Q���F��	H�-��%-/�B䉣P��LEa��Kל%sՊ�q+dB�3;V�S4&��*LA$��PaC�ɳ$R��? �н�V�R�	��B�&P,K`�ťM(�!kŔ�x�B�	�c%`b%�=`z��rER�Qk�B�I�D�b0�@�T�2tȲ�L�{��B�	�
��xQ�l��"�
��J���HB�I5h�n����2r�AZ��_,r�C�ɻ�B��w��>,K�qQA�&�B�	�#���q�Ħo!���v�T6	�fB�4i��}0e�N7/�NI2��p1C�IMF� t/�W@:��4��,�B䉒(���C@ͨj��0z�_5w<>C�	�j���0~�Ĩ���mp�C�i�j"�C�B���a����"Ї�O�&�3Ɗ;}�@���"�'}�ȓ�LBT�ڽ\��c�(��(fLB�ɏ<��U"�o��{���b!Ϗ�!-lB�I9GN̬8td]�h�	é41��B䉨�f���Y�+�1q@�B$GT�=�
Ó&�m��nПK̸t
�ʌ�vR0�ȓE_p��4�d	�*%�C�	�g� �r+��n��T��nl��8�I ep���ԽbW����#7��B�d��b�K�"m���P-7`.B䉲����w�ɝ>��"�� �Pa���E{J?�C�m�w��*4�]���%3��&D�8���G�mʠ�'�6y�)Q�M%D�,h���(��E@pJ׌:1~MV�&D�@�U* ������2!�09�+�>.O"�=%>�bc%���)I�酴J�8��Ĥ �O��|�,e��[�m���H��L l4��9oT5�W�1c��Z�U"u4݅�2���tI�q-�8(ק��( 9�ȓF���{��+���i_�h��чȓ�x-AAH��YK���.U�s�z-��U}֘)"��?@��Af��%y����H� 	 �,�-9}L�k&*��	F8��s������a��\s �./
���	I��!0�
={��58 !��X�C�ɺ$Ӣ�r�D�|Ҭ<��n��!�� �l��K!uG�T(�+эZ�l-��"O�j扂�qZ���L�_�2�K'"Oh�a�ʨpP�)�K��_Z1yf"O �p���%b`�,0*R��ku"O�@��ŕW�laz�!�0(ЈC"O֌��ѓ^퀍K�Fղ"� �"O��Xq�# w���ħ�Ȕh"O�)!�.��0��`PC#�� �"O�`��h�J@��
#-��w�L���"OV,�v���|1�L��&!a6"O�1`"���Mf�H P,��9���۰"O�0K�N�9`�v����!p�X�x�"O
�)�`�Ahi@lB>5��S"Oz�p&9��tJ%�YS���X"OL1���/ I�%Y��Y�B���"O�A�g�m0<���dt�|��"O��* MЂ�>�!@� 9쥢�"O�hXS�D1rO���S��a�x�b"O�
P؛��c#��T����"O��٠�"̬Y����R�F��'_^���`;&Uh�L �xҪ��
�'�����ϗ5��� ��2~�p��
�'�0��e@ MP-����tj��	�'��ɹ�A#�`���h9����':�%*�!�g.�:�@�6�q�O����T����j�	q����C��h!�3�TE#'LH4	���a�;ng!��_�/|���.ې<��]�&��:0!�Dӡp}[a��NHtay��L4K!�T=LMYԏ��<H�	kE�O�!�^�0�8e#K,N<�M2d���!�$�:�����k�H�0�07�B�K�!�d�<됉p0I4���R��ĸ��yR�]� ��r�C�}��%��ğl�<�v �	��ɐ��?.��a)�H�`�<)�C]M6�Z0'�$Jy�Q���N_�<��!l��V샫c���0Q)_Z�<��ș#T��q�b�}`b��]U�<!W�t�ZAAg��&e��|ȅ��V�<�%�\�m�"M�@�K�g^���'�U�<qs��#k��#(G�W�&5b��]�<�RK��"�^A�QB�n�V$jD�[�<�5��q�X��5���?�X��M�<F�J�!4 �G�H St0a�GEH�<Q� 7��@�wc��T��Q o�@�<�7�$���ǙQ����a@�hF�C䉸K�����W�>�v(R�S��y��+&���M(l��(�y���K3�(���J�XI��c�.�y���������$�=R�4��	=�y� �0#�
�as�ة����T��y�K[�YL�"�<L�谦)Y�y��b��ܪ����U0F���y�gZ&�=�惚�D���c/�y&�-j��z��z�L8!��В�yR�аh�Z�������^2�y"��LR��ǎ��<���c�V��y.�9Q�7K�:.�^�[F�ҹ�y2�������a���"�Ҹ��G��y"�Ľ&�H��$lC��zE2aHS�y�f��/H�`���M�ژ ġ.�y�I�/FZ �w�N$\ږ%Rd"�y�	�l��S��_f�֌C�y�L\��"���WZ*�+�$N/�y
� rPaա�=X���z�
?�Ҁ"�"Oҭ�4,ƞ8����C�l�.�"O(-��Z�l��+6��G+�XiC"O�h#��~�:V�S�<x�`�"O�Y�qmQ�,=B@�IY�fe|U�"O��!@+�2.�)�I�ad�{u"OP�(g�]!P1`u*C@&<8=Ȕ"OT� !��S�p� s"ȵNr�("Ob��+ۋ&٨E��+�$]騬��"O| ��BCw��@�N2	����"O��Qi�)�h;���y;>���"OΩX�P�;�8R�M0�U��"O�u�BQ7a�u�K"U�*b"O��B�[��}�R �-Z Z�"Ovu)�K��E�j@a�m!(l�у"O&��f"��L�LH�ČNx��"�"OL���,� Z]<�1�lG�E�5"O|1�ۆv��R�$����"O��&c�>%��s�_�p�(F"O`H8�ʖ]j1��D^�J�� "Oz-h���u�ISf�IR����"O���f�+[6�x��n���9C�"O�B��E8^��<x��r"OLH	�DN/R�&��ӂ�G��@�"OT1h��"�0) �݅�^�x"O�TRp��j�3�I��2iCs"O��+gh^8���f� k���s�"Ob	(��Ce�\I��\/ v �"OU�CN�W�^� ��/v��}�@"O��dhS�4?��h��F<�|��"O\���Zt`,rWв;�F��"O,�a�g��D�����p�dc�"OT��ǚ1&7��p �Ńtq��"O.�#��+�6��"�9{s��"ObH#`��!��x�!�ƢD�6 ��"OPb�
"9��p�������"O����i%��!��hԣ ���R"O|Ջj�0�aG˓~ �Z�"O�,��j	!Hx� �E�!{��\٧"O~��� ��0=�P��	)p���s"O.9�W��?�H��Ղбi U�$"O�db���+S��Yu�ȋa��Q�"O�L��GZ�O���R���MG�`��"OJ�v�U�!����#"K�U�j�"O���V��;1�[B"�2TLݚc"O ��$��8��|k4�$0J�y{�"O���Ԭ̋4v|P����uF�5P"O�Q�FM�5
h�m$!9���"OTY�:3r�#�
�k�D�0f"Oج�f��;��Q�Z	G�lq0"O*Q�rdW�dT*��@w���"O
��!�[���䆗*,j���"O���j�l��I5#�6U^\��"O�d�W�[�k��H1p���X|� Cg"O����g��B�0`ӏQOez���"O�h�$bJ8`��y ���-^�4b"O$���l&`��l]�Ma��{D"O���ŀi��tx6ldS`���"O���� UC	~j5��;4��R'"OZ�K!J	y_�dQ�I�T��I[v"OpĚɋ=^�j��%���~����"O@�"�Z��lr͜�c��%[�"O� 3��ޒ\`�E� l^]��9p�"OE� ��5X !�Qʒ�6�z�R@"O� T]�a�k�^-��&\�8���V"O�X�h�$S朒5�?�\��"OL�[ǀ7in��ac�Oh�k�"OtT��˝�|o|��U�U� ��"O:���Pr�&B�X�&��v"OZ�XΒ�?f�*�+s����"Ol�{eρ�)˺�sF�ϔS�2!��"O���Z�p�d�؁oWX�>x��"Opi�F#�|�\x�dP�F�T�s�"O|(JdaV+Y��0��)g||��"O�Y�R��JUp']�4ZZ|K�"O`:We@�b�ec�-d3r�u"O|�j�W�QR(]�R�f0YP�"O.���c�;Ld�9�d�O�]���"O�`�̿^I��hD-�p��Ȋ�"O� �W�5a�"}c�*ۭ�*$�v"O$b@�ڨb[��q���U����t"OP$�c&O</X1�'W�${�d#�"O\��t!W� ߄)i5,�4&מ��G"O �#J�we�����
�#$=z�"Ob�����3t�|Bi��@��D �"O�x��\0"e���+���"O�|J���$zҔћҡF<i<D"Od$�7 ʴE�rx�^pR2l"Oz��΄F�]zv/�@���� "O�D{0�87[>8CT���p�0��"O� ���ߢzN��P�W1P��"O�P3�Ο>oB)�E�ʺ@�@<P"O�0fh�5�JC��P��>�b"OTeK�Z���)����jt`�"O]��ݒ�fr�-ɪM�Y��"O���a��?�6�X�L�J�>��s"Ovmh�OC�SV��U�Z�A��%�y�լ9�±��hģN�X�Q�߬�y�\�+΅�C(N�|�n2e��'��i�r��%�<��O�#Y"j��
�'���9���+x�@D#�*@��Ѩ�'���ݓeS���Z?+Hԉ�'i�U�c�ܢZ���
�h�;\,���'���VE	�S���E`��8O� @�'�*h��� 6�����5*^ѐ�'f�M"��������w/M�XR��i�'3,���-�2~
LhDŐ]I���'���BQ�����H.QY���I�'0�e��I!y L�S�\�O��'H��V
ގ���@Ǟ�u�0���'ݠXC�$O;:5Ps!ȋ�8��e��' �����UʆdS4fЫY�|(9�'|���b�Ows�,��Y�M���q
�'�R�BE	�)�TJ!L��m�1S
�'0�Cc�%Q�ع@)V��M �'������G��ቀ/O�NYX���'$~y����k8�s��A��ih�'�d����r�hx��3>�}��'�FTCd�/ZV�jG�M(-n���'�<`J���i�>xA+�*z
�!�'<LQ���?{:�Ѩ����$wL��'����%�/�0�
�H!�hm��'�:h��L6\���ɡ�Q�?��� �'����ٶ71�b��<�T�
�'�B*�@aX���7� ��
�'o
p�E(��|�5OT8'���	�'K� #4NL $�l|���-�F]��'n� A�Ӊd��ݛ�%?_�l����� 𙡂�0��Da��R�r@q�"O��;�䇁��� �#���vDk6"O�t���g�@ �ԃ�!��a�e"O�`#E�$̙3���;���"OLa��Ie��� � �3k�4�ٴ"O.���^�MJKQ:j�XbE�4�yλ��#�� ]���)��� �y����m�G�D�N���%�؊�y��,O�t�bg	�L���,�2�y���g1�0	�ȑ�7���1CM�;�y§�=|���SJ�3{O��ӣOſ�y���T�d�U���W�i�ᐲ�y"��p�TX���%q-�)kfZ/�yQ%Vv8�1��N�dZ|a;����y"�%_ ��R��k����vfF��y�,�$��VJj.� V�Y�y���2bz�VgH\�)UFץ�y�� �q���`��hBDoŷ�y��_�u,F�@��G�Y/���
1�y�lU�2����0U$Ԁ�	��y"�;wq�����S8E�`�9�G�-�y�_
2�ր��댁l�D��!���hO\��3Q��@���8����F:џ�F���0R\Z����R��� �����hOq�ܘs�b��S#�d��[F �j�"Ola�W*|�=HE��)g�6I��"O.P&K�-�$��Ą˙s�j���"O�Ġ�m!�^��EiOYpTi�"Ot�@C�7U�:U[(�ak�y�U�'��Ⱥ����[nx��Ve	�ܬ��p�)D�x"@���6@+㣈�)u�б�-D��0�b�NdNi�Ҫ�'��xk�)ړ�0<!J���d�������!z�R�<1P �;*:���E L���qd�P�<��LȊV�����l8�9��P�<d��i����UM�I�fe�t�I�<�-8tC.0Q0Bԁ+����G�<1 �K�j��9A���;sL�+�j�p�'�ax��.OoD��Ƀ$o�8!:�#����<���G�>R��� ��6��0�ΚZ!����V0xbK�8� -�v����!��$:AD�� �h:�k�"�!m!�䗴v ��jSoB�s��!��X�Z��'�ў�>��1pw�x�H\9`��@�Q#9��7�SܧhL ��ԧ�l56ZF���g�H#��͟d��5Q�ϛ%��=E{��OȂy� �;e32�ڞ��y0M>�,c��`�Ӎ-��-�gO�V~Іȓ`X��'6��}���"?~!�ȓF�r��%�"jO� S��ڟj�
D��S��xĸP,��6��D2�k����C��$��y��;j�B�j����x��C�I#n���Y����|v̈1����?����) ?��+b[�KED���I�<����;��Y�4�{r�mS��K�<Y`O��X `�YЦ$SPnũQ�F�<�2��{KNA����0I  �m�~�<OխC�*���[�K׀�#3��}�<��UvF��$�^ AmH;C��A��0=A`� �JlB�9# _�O/���U�V{�<��q��x�l�9jv��P��z�����O0�$��N���
�nU�����'���S�%�g�p���<�(��' RYl��;<��B�Ԟ.k�%���� <��b׎ }(�(�Ý�F��q�S������|�&��CO��P+|��"A�-6�C�IN)&��P��6"��5�t�O��x����x�'�d�D��l�Q�S+�x ���x�
��z�u �R9 5r"F
�y��Ăr��9�M��*����'���y��]�wRIaf!�r�0DF2�y�i-�`jDjq�e�R��y�ƅ;Y�|������ 3��8��'Gaz� 	y��%���4 ��KAn��y�A�� :�&Ʈ) y��!9�y$�"���5���'Bz�#P썋�y2m@�B*J�C�3{x��4��yr-C T�Xӱ�Ψ�����y�g��)����e�_>o�0pbC���y�J:�0�3��LQ����T����0>1nR38���ѣݥ?N��R-]d�Ik�'����<aD��Isuj�!A8���[a�<�V��v������on`AkA�x�<�T�1|�
8�T�:K�R\�C��?J\�YB$��Q����E՟B]�C����b3C�:Dp�eC��Q� �C��/pu���!��*�q�^1Tn૎"�)��lN֎�"���#WX^B&�Y��y򏀰<�j�S�lQ#Kn<U���D0�y⏇=}�
����Ќ>� �����%�y�E��ZĴ�#me� ��װ�y���eH��t �"U}��hQ*���hOr���@+[���kakŭ(��TK�
��x~!�U,v���%	/+��hC�nF�)�!��I#�J����@����#��2O{!�DǕp	�£K�El�}�`�MI!��kH����٘Kh��Ӕ�Z!a�!�ċ'@�<}R$J3�,������!��_z��Tb�
|8�:3*���!��W�b����I�p|-Q�
��!��\C,�|yvN�U���cB�7��O����xg*Uh��:E���O�${!�đa[J�;��@�%#TJ���S!��@6��tI.��[p|:��"C�!�64�jL[��I�h�1ɖ�!���)�`Pg�_�"9H�'O�!��5I��x���v�8�c��r�'Vў�>��>Y�a��6UʚT�§8�$*�S�'�Ƒ��L��^A �Θ�o �t��	b~R�.���.��җ\ @�J��
�'��#G�� p��f0��	�'k��ImQ�=�aS��D�2<��x	�'E���/Xǂ,s��#�����'�`�0����У H#ZBQ�I>������1?v�k� K�vXF@Ƃ��+2!�G+x��z���
{AȘ�C A�,!�D�!z$�5�ƤKV���<L�!�J!�����%��DK���A�
|q!��U`�d��@j�?\B�P���!�Đ7v^T�WJ՘!Br�h�/G�!�I�Qi�焦j�lhq歁$.!����4@���V��)YWBƍ<!��L��1��Ց:{䍑�Ւh�!�C�0���t/X�Wu ��Y�!�DĚN���nmb�SO	�!�$	�gy���g��`�`���z!��Ta $��OE�p�N�BUI@��!�$Q�e�p1�g�����a�`)ȣXo!�� "�ʎM`h��lDj��@�"O��Y�LN90#Z(Ɂ,�)���Is"OZ����IUR�È�;?�d �b"O��Z�fQ�3�j�����k����B"O�
6���1����0�W8�T�p�"O\��3C/w�dʄ-·v�>�1�"O����.��P��A��'��'��6B׆��􆛜_��@�ȪB�!�Ĉ�G]�rdB�
����흄*�!��)g��I��D�������&�.�!�� �)f`�i�m�>w��mC�LO�!�G3� L�g��J����i�N�!�K2F���-�0�Rq�o��T�'�a|�E�'�<���'X92 �j�P��?�(OL���P� ��`i�iA�X
��6d�o!򄘔V3��hs���y
F��6B��3|!��D_�\J��Fz^�����Mx!�d��Y��u�vJJ�
����!��SPnm�En�0��-�6P:�!��j�$D����6�r R�횎b�џ�F��M��2��p-�<O��v�B:�y"��>��ip�+��E$4k%@՘�y'ԹBo���g��<�P�)�
ŷ�yB-Ln�R�C��A-k��TnK��y2#����!c(  ��<�'
��y"f�2-|����$�Pˆo���y�e���҉�1�Ѽ"�As����y�	ՇjR��#�#=�ƍ��ɨ��<���D4�\@���#�V�X��ǚ*F!�DV*L��0��RF�0S��,[+�y��	� JmX�&�WHf��*]*"B�I4�e�����iX(H���+'B�C��6q��qm�c����va~C��1R@��A�����p��OE��h�=��'���eZ�u|�[��Zܰ�ȓYa�S��>�h�c�FIa�Zȅȓt�>9su�B�m���5� �r�4���鶨��F�A]]��,��F��ȓ_ЮL��	\t0ؖ��'𮹆ȓc�l��3,����[@�A�Ky�!�ȓ7=��IE	j���EdF�%�0}�ȓ��-�rd�(�X��s��=�DX�ȓ���h�G����cs�<i�x����T�f�F�T�����6<N��d&^���#�����*s����ȓaP���2��9���7����qզt���c �#6NM�Q`v���$����m��镎�3����ȓT%��`�8r2s��W��%$��G{���M�v"8�;�\�>-��b�X�y���V���<x��T���y"F�T��z�㌮~�t	�$�E��y�&S�#( ���B���tɇ)�y�j]���
��;����AG(j�)��#%|LR#�϶5n��&K��j�|��ȓ!������Ի)�: ��q,XY�<�ǌ�0���@P��y�ҋ�T�<1��S�F ^�䁛�FsМ3b��w�<���߄mP��1�.F������p�I}���Oܚ���ɗ?��´�:�pQ
�'<z���Ƃ�Ϯ�Aw�^���$�
�'��5R��8.+���(� �ک�	�'|` ҖGр�,֯.�d�I>y�z^�I�V žDz��RfEI:l�p���S�? ���
 9�FPk��l3����"O�������#]t=�w�]"D!}��"O��&֞�(���Μ6n�ű�"O��Ђ���v��(����c\D�""O�Qc
$T^|X)w ��E�x���"O& Z�/߹')SRA�"6T�p�"OU��+L�oB�(���Q��"O�ɓ�%��(���!�0|����G�'����ʱ�iY�}����Y7T\B�ɵG�J�(���4����[	2B��7
�`��E�$O�q�%n�����0?��Iו6�z�pUbY1|�:�*����<a@KZ!�&���
.O�Z��v��~�<�Uo��B�(t�"��	��[cN�}�<"'V3{Ĕ�J�/=M�Лg�a�<�5�& ��l:�l͹}�l����`�<��Ŗ��!��H=�2��І�R�<9G[0)���ql�UmyfKAP�<�Ч��@r���	�B@��NZK�<!�@���䀐��	Yj�@D%�]�<!G�	y'���BgQ:�F!�*�n�<QBF,�.�el����C &�l�<AA*�,�j�`�/c�l�K2�l�<�aF#����G�"{�.���͈k�<a���@��"6���+�0����j�<��ܤ[P�J@����D��e�<�#L��M�����DЬ7�� ���`�<�BE!l���#Q�Lޒ����Y�<a���3h��c�G�-Z郔'�Y�<y��3M�!�c� OA����U�<���*��p���oV���N�<��˝9_C�ة�X�nI�y9%�M�<i�@�s�^�I�*��9$�MG�<�o[�r�,�@d�d�T@Q�Hn�<9�.��E���i0 Ô~V}	$�Rm�<��F]�S��H�sĜ;E ��*&̚k��hO�':�!J���;l��g�eI�ȓ�M`Ʀ�)�(@T��!�r	��K��|��k�h�I��Ɇ�D ؠ�ȓDI�E�J�ʅJ
��!��|�<�V�ι\�p���7�ؔYâv�<�w#�;Jz1��.4ROd�I�]r�<�+ۊ`"�=化�Rg�:3I�F�<I0b�8.�1!���N�����E�<���Ő՘��D���:p��DC�	�F��-b��ڢ,v�UkEOW�(L�B䉘?������i<����V;,e*C��	h�P�7��D~UkQđ�N@ C�'��哳���/*�T8���2:w���d$?��-^�	E�l��}��	���t�<�K�
vŎ�cal@���Pƨq�<�&��?>w�t�삁W��`�)o�<���M�w�l��Ũ(?�J֮]A�<��K�z���xg" 9JV� R�<a���v�He�!
9ȼi⧛K�<1؛x���᪛!X��a���k�<�m���(	 ���!�Fi�<) �¿�\���--�xi��Ky�<��0pkH	�*D���bNL@�<iEK�� 6<8��R#p��J�I�d�<�R�P�V�~�4�� 8_��R-a�<)ck�X}h(�6�0��X
VT�<��a20�mb��:�
�.�S�<90�3eD���U5t�����Ux�`Fx
� �)�W�ϓ{?D��`�݅)ٸHW"Oj���L6_&� WC��*�vtI"Obe���y�� ����q��jC"O�Y����Аj�D~�t���.�S�)�b�6{�Ԯ8���G[�{=!��-v'��i�� ���1%��5O!�dߟH�
�A����[fEL2!�$� �$0�ƃ�:�t��d�!��Ob�=���ukƢڨQ�>Ts"��4_\V<�"O,=k-�T��d!	A�W�!k3"O��C�B��E�g�;@�~���"O�����H����MJ�"�SC"O�)%���W��|�7FE#��RD"O��D��[��� ���k��@�F�z>)��`R�r�
P�r�_�i'����Ĺ<�+O ��7�&�J�bOC L@a��p�8��"O`1ƃJ�E��x°�U�<n�b"OJ���DD$���&�/Hk�,��"O����
��\�-����f��KG"OBI
�7v �M�񯙿
c�mb�"OTP%��
�����JK�h1"O� qwjİ&r�Vj_��
�����Oأ=�'X�x�0ԉʌb��Ԛ%H�6d�L��Pa~U��J�?��zχ2M���ȓ%��e��'��Y��P�߮3f8؆�?�\��bʄhGN'G�D�ȓ\~��$$:�y�Q�D>\`�ȓu�@P�"h	�{���3�J���l�ȓ�T�a�׏S�TY�んu. �ȓ��M+3 �-/��MC�ꀕ;���ȓ/�2��������sEm�i�✄ȓM�e�T朅1D,AS �%v����ȓ4�4�����0q�+��!=X�لȓՂW\�!��=�� �<O�x�P"OLa@ ������`ƅS? D��"O$�@�HZ�0+��-(��"O�qb�/$�vD�&����D8�"OX��U	��E�.���
�����"O&�KtC��u��(q���z>��E"O`�{�����ʅk��g�P�"O1��M�c�N����7-hL<�'"O)@r%LY��p2 'ϖM]���q"Ov���C��O�D�[��P+LS�dI2"O�|�!� ]s��y"*�%�>��"OJ�Y�S~�X�`@#G]��0��'��	�6�����Q+bp�$L�4C�	:�v�bi[�W������FdC�I4_��@����)hX��.O�DB�	1#_�ѩ����J� �B?H�8B��*.��eR�b�r����f��(�"B�	+Xk q���ڷo!�B�ɚ}o`ȊW��(�İ�$�\RivB�	A<z����	 '��d,��O�C�	O�8����՛D[�FF�`��C���%���{%�8�|��"O��O��a@FXaB�P��p= �"O:�r�Г:8�z�M�;��ʲ"OL���k���Z���S�;�HH t"O`�cb,U{JQ1��h~@QQ�"O�� 4ĝ[�q�L�k��c"O�mj�̕
N�ՠ�JH�,�J�Jd"O6��s�]�|�:��ށ�tt`�"O�@�TH�02�IuGK�N�z�"OT@hb!�4'��M*�-�Qj�H�"O�  �r@�P=�|��5Ɯ�S{��a�"OH��古P�,�4@]�A�da"O>�HD�c�u��Wx����"O�iX&@��	�غ%,C�Bd�'"O��(�Œ.�@����1+���Z�"O`P闇 ��/�/�TY�"O��X���E��̈:�.Q�"Oȵ�0C�7�6AF��l.��(C"O��!g(�M�6��!h��H�1"O8QѓҒy�L ���Һe�Җ0�y�ŝ�b�B82gb�	@hZ������y2�I�o��EI�ď.Mdc���y�%Od�}Ycˈ%��DQ0���y"E��5�0=hu#�O	�tSd$���y�۴>w�M�F�E�vh�S.״�y��?w'�4:�i��:��8��)^�yB�,{�`	�$̎�1��$��f��yRG�#��L��$�te�ä�����!�OL�H�%��T�Z�:�`G2pq^���"O����K:�$�QW�Ę`"%p1"OB���u��X:�-E�NL�$��"O~\h@�4F�t��FT� V5�"O"�@��%%T�Eo
�U��'|�cF�D�[ ��k�	�R����'5d``��uQ� ǂЌF��)�'v��JU����&Ը���'�R��
�' <��SF���(֫P�1B�
�'.��7�(O~T�ȥ��*+�L8)	�'���*pȉ�.��Aش`� p�h�	�'? [��,I�f��qX�� @	�'�l�эNL����AĠt���'�He��C@q�3Kքp�R���'�H�3�/�-,�}�[�lY�-y
�'�X�h� ø�����Nxr	p��y�@��<ҕ�C�=*���[aDI��?��'���F����,���Ƙ
L�0��'�Z����K�_~�XYQ���|Q0b�'S��)Y�?��e��,=�NA�'�p8�I14������*�T���'qx�Q�Um��H@�E��� u0�':���eV�Xࠨ�b	�(1��'(f�2��FĂ5zu��*R|f44"O�����;tV�z�HL�I��"OH��!IK0��	S�N0.<:�I�"O�(Y	ͭO\�3��G�rz���"O�|���ÆcZV<2�D%\�H���"O�y��@M?u�]�t�+}.�˂"O�2��R�"�X��vbI�s��Z�"O���5�������DBk��R���D6�O �;�Eu;B\�g��G��a�1"O��y�HW�dU�e�4%�����'�p�e*W*��B�D�V�9�'^~d���<�=�1FN�B�y�L�edPi�A�;�ވ:��P
�y�	T�M�
����N�:c���Q&�y��?��!�i��+��I"�4��'Jaz�(P�}� ��eω#�xs����y���Z�B�D�i��lZ�(G+�yr.�.p�v #W$װY�R�3c�O��y� Ҥ1��q�P�Ь(ب�r�c6�yB�S�efACǉ�P�l(����y���B��4Q�HH�H�ƭK��ݫ�yjkh�� ^u�x�0J�y�U;��%�2g��ӇF���y
� �U)��-wy���T����"O\
E�6*���I�*�>[e�U��"O�X!6LЁJ�&������{"Ov	�Fg~F����A;;�����"O"�[��?S����&I�]'��"O�hI�R����bfF�l� Bd"OP�C�\�&q�h�#U�z�Q"O�5z�/�0{f���fc�<-�ꍂ"Op�
�G% nd�#T85[��4"Or(��ʓ@� ,٠a@I����r"O����#�;Q��x�31-����S"O(��Aa�q��mT����o"O���#סK�^`�&cD9%�� $"O\�(wI�2J�xl���O�b�C"O��B"-u#J�
u�L�L���1W"OL�[�O9�lڒA�C��0��"O���.L1SنB ��y�D�Ä"O�E+���.n�T �a^��b@#"O���M��z$�����8q�D���"O�!�DL�}���R�-
�>���˦"O�@1VeE�7(j�����/;��"O>���l�Τ�����$<h7"OM�ӊ��25��:�U5��D��"OH	�rlF+g�x���?Qڌ��""O"p�Eꑍo�P%��aײX]d���"O�V���/�Ea��@X�B�"O��R㩋� � 8�).,-��5"O� �d��0r 1�Ph�$^$L�"O��p�I�&�v$�I��`��E��"O��*1�\�
���*y�z�cU"O��fF�i9�ybP���2����"O�����e�4�+�^����c�"O� 1�Ō
<�P��DUx��+"O��bV�DrB�1��)�9y҂ �"O�̪uk���I���&#f�dp"OL(��nS<j@+d'�4����"O2�93��o���p�����5;�"OnT �L�d���W#���W��_�<�HS�"�9<�E �-�S�<��=>҈4���܃DЮ9Xc'Q�<9�n�$w�$@�T�CV`3�^d�<YS�bj��1��.:��T��G_�<)��X+[�ro�)-����!�B�<���+�e{�ʋ#}�KUHOi�<�`�?30Kd�
�xt��(i�<yf�Q<`�ѧ�P(~7td��K�<g#�?b�H������ � �-�]x�8�'���"c��5�
1�`׳[�|��
�'ۮ��D�'L��r@M�6F1
��	�'s�p���Y75��h�į@�8z�z
�'M��D`�+c,�aHܧ4h
�'6R亳e0$����\t����';>�$S�Y��A��.<u�BP��'|<)�e'J5g�n�2�Q�j[b 

�'�*������֠��D���&��
�'��*�c����K���c%Д3
�'����g�,-�QfGA7' *
�'2�!pV<H��9���	v;	�'\�9k�A�6�.y{5�W&����'���A�?&�$49�ۚ���'�(��������;���'���	eU�f������-��"O��3F�V$dn�ȦCΫ\n�#q"OZx��'�z"�?\�@�"O� �x��S�Mt�R(��j��D2"O����Ι.w;Z	���(~V4�W"OB)r�gM}�FQY��S� VR�X�"Ob�xŇ��b�����D�Dd@*�O`�T��G�6A1U��,^�:�xT��OPB���&��PփRA��m^�C��4x2%RP_�'�����2�JC�IQO*xQ��:����d�~4ZB�I�k�(��o"$i�AӦ!��R�<B��&E�|pb��T�m�&a2A�+ �&B�ɋw����^� 
%�U�$-0B�I�~�RA�P��%Rl.��ՊJ��<�&�D{���+�����g�Z�1��,�C���yo�����j�"�p�3�Q)�y��?nb�hEc�#h���B�W��y�삽R�� &B�;a�~�9�bݘ�y���ff��W���*�x��T�1�y"!͔S� )�G6kE��Th���y�	 G�T0R��j^�i�5.��y�'�:m쨱�h�N�KD���y�J�Z��U��@����)3ɘ�y"Ϛ+B*,�bT���%�r,
��y"�X�q;������� ť�y��V�c~����Q1l�(BPKC��yU@�*y�1G�Z�x�����y���H�����d�e����5�y�l�(bX`9�'V4��('#�-�y��8B�0�K�R���B��y��3�0-����*\��	��y���gk�E����k��g<�y���2K��x�'ò�f� �AǼ�y���D?hqG�U\�,H��G2�yB�@�+9 �cd��a�تvBօ�y�WM�ޜɴ��_�xI!q���y��ŎI��˷h�?DCN�Y�j��y���S�t vd�$�b��+�y�����$-��~�#��^��y��͚��c�>	&�C"KW)�y��H� ���FQ�hR	0"�̉�y�j]�6J�x°�X6���y����y���1]�o�$�t� ��	#�y2��;^��}�Fď3<�6D����y��;�.9�e?.6huP0	�y�!	BnF6�0aEH����Yi�!��\h�=��l�[)�]�"�	b�!��>g�v�d/3.�Xa��&�'|!���e���x2���n�`�"�p!�Ǳņ��J�W���	v��Wb!���f��iЕ�N]S�b�a:wU!�D x��8jV� J�1c�`[�H!���7�F�;V�G=jE��)s��:�!�d�t���z����  n��F�W5�!�$A�\5�=�pƻN���m�js!򤁲0K�� !��c�#j�	=�!�����`��DM�N�Rw��	!��.�p�EY�z��8w*B�	�:E�9���"Df�� ��:L�B�	$@ P�I�<}�l)��1�C�I�b�0b#�+�8��A��F�C�>'Bi�a�@)%t|S�$'z!��D�F�BMCDS�	3�A�����&�!� s�\���(��1���®+�!�D�g��bV�!l �.��O:!��'6�J�hքS2*B�a��.H�!�� �d��.0w�\�{�Ù[$Hã"O��[�Nߝ2��`З�W�A$�'"Oe��.��K�"e��Ce� )�"O�p��ߔf~@$���֨K��}��"O�"�k�qRΥb���O����"O�!�1�X-N�ȡ�4k�(�"O�R�`ڪY��m�q�F%�"Oz�z_)n�KBb�H�r�+��t�<aPa�3r~j��1�3d}V��[�<	v�ɓ��e�%"�1�`I����<i3�����2fB�!��d��Jq�<�&@N�~sfQ�#� ~�J���/�C�<@�R�l�Sw땢U��9�uz�<�S\����ǝ���Ш_�<�"惲8D���h�p2\����Ea�<1sL\&J@�B`/D �!�/�s�<Q�֖dz$13'�'3����.Ll�<�+�4�4Pb�c҉cAE�#Ym�<iw-�2��͠3+[�`b�#2�~�<�d�;'D�D"܀W���Ox�<�� ���q��LQ| �"�MHt�<��@M�d"}� _y81�VCBo�<��G�{�N(AC� �D0���i�<���[��d]	n"tBE�l�<a��Zx�1!���w��l�eÆs�<Y� :R�ְbE�/c�Ƞ� �q�<I�C	��1 �%�?;�����DMo�<�A톽nh{T��#|���
�g�<	Q.�<b'�)�	�&TD�y��	d�<�UfL�A��	���C#��@U�<���Ӏ,3p0�A�ӥ#��հ4N�R�<97��f�:T�֋ӇG����f(�Q�<���|�<Qѡē�t}f�%�S�<IEɃ/9V�02b�0u:�z��R�<A�iD�НX��Q(K� �@CTE�<I�o�O���;�&P ㎜H#�w�<	d��@G:l���E�l�Cchv�<�#V�4&&�22�R"�"�"!��q�<!�(��%��\A��/m �)�b��l�<�t["6��њ �@)Z �]�4�\M�<I���Ӿ���K�	/�+C%�J�<�BMM:>�tA���"������]�<�W�#��j0�&^|r9Z`O�X�<9��Q"
�VD`Q��$G�F��o�L�<a���@��h�U���QP� F�<QVe�-���#�Q F:�P�A�<afk��,��:�AB�U�v鐵`�y�<)��ȍG߾�;Mɶ<U�]���q�<�� -	��R�F\��J`�U$Jq�<9\N���c����`ĂF��!�$�2c_Lx�$�����у*�!��Ro��	���+�-х���p�!�DG�F�(�dS�8	�}1�=�!���N�Mj��90��i ���!�D�sN^$yB�Z4Z~e#D�:�!��W�jp�"�(O���+��Z�>~!�$�;<�Bȥ.��"g豢T�N/A�!��?d��j C[�d�颴"�V�!��ϋ���r'�`F*t�c���!�=
.�1b98�ؘ����lu!�DO'p�� ��mߝF�E��Q�pg!�d��h%�Ԙ=a ���AO!��R�
������xARX)�/!��ث_:$9��a�;0X��ĕ�j!�� L5;�cW/|�C���>0�P"O0R���-aӦ)��e:�:"O��@T,��e�J	Xp&��d�RQڠ"O�����VÒ�S�n÷�"r$"O��� �����l��,�*�"O��ԥônL�A{�m�	f��H�"O��7�p �ݸ��_�Ph�:�"O�SF��bąH� ��[I��8�"O6�b$�:]� Y�͂�$2����"O85 ���%��h�`L_4_,���"O��	D��fHW�IjJ�)�*O.�I�k]���eO��)�'.�hǆ�7����
���B�'~��t"-?0��B�H$
2�Q�'2B�@1'��B�:���d$��
�'frY�v�G�$d�X$';Vg��A�'�68H��KK.���]�H���
�'��BǂӌP���Ίt�؅R
�'6(X�#��-T�a�#Ѵo���
�'��ՑtmOr��ˀ,Ѓ\��H
�'��tZ�h�R�Cp��"(
.<b	�'>0��d߅$Y�t;!�~t���'ͤ�Ӳ(����Yj#��͛�'�\<rEL�? Yk���@xd�'��azЎ^�d��,X"_�� �'Kp�A`�E�8��ɸĒ�
�'�0Y�d
G!������ݳo��k�'_ Ax�B��t� �&�Ǥ7/�m3�';H�����;W���o�_�9z�'|=���A�F�
�8�=�	�'�R-Jt�5�
ȹ��p@�:�'�^����6O���)�Z���'1��{���-�`�SR��!R!��'ᄄ
��Dmnv���dS�'h�8�'������% K�6d	2�0��'�!PA�Π;���,��r-~dY�'��y��&M�2!D�[ŧ�=v9����'h�x#7��(<�|h�΋#n2z�*	�'���rSN�'�������e ���'z��"���k���(��ʊd����'���Z�)܂V��<���6c�jA��'eB`��)�Z�|�r��֊�x�'䔽j�NR�M�z�3��/���y�'���hQ.Y@�Ӳ�͑,�8�'��@p�������+Y1V���i
�'��5�⬜S��5֍P:b	��'�P1�\l��[�,W�Eb��',��V�S�wM�LJ�bǝD��I��'�6��cZ�s"��NΥ<�q*�'����%a��psL%���G�=ޚAQ�'* ڇޣgz(p���B&3����'�݀�B]�:V\��4�@�0P�0�'�@`���6Y�&�"[f����'��$��K�c�Z�Y3��)T^�$C�'C�b��� >ڍ�bV?,����'�x��#��Q+��+b�&0�j���'լ��b�IS��x�Vi�#� $��'B�(\u�:@I��٪"�hi��'N8�R2��]X(���$F�`�'ȡ���.��w˓ HT:�'��1�Ǌn��!k��N:z��q��'
��gIL2%������@�"a$%��'9N\�RBV.q���g��p�'O�`h�S�M�hp�v� e��b��� 	�g)�&���N/��q�"O�5J�b�%#���E�D/m�J���"O8�� #EM�~�kT��8O�N�۷"Oh4�GrrcŪ�1�|C�"O��3��pbԩ 1�L�]�X�H�"O
`�C�&J��6�5�8���"O�ݨ`�s�T˷�ݥQW�Mr"O�Țp��;���3,`�@�"O�y� '?�h�щ��R&ى�"O-��� �8���@Q(_5�^��"Oĸ��a߿x){��]-H}�"O�PQ����;�
���Y =����"O:	i�j��x��!���RR�v�P&"O`hHܪM@��r��h�"OL$8�æ}L��2�@�_�m�#"O֝���I."(��E�A8sY.��"O�,{@/��ձE��
V��z�"O0u�R�-BC�aI�� 9Q�e"Oց;`#W.����%W��;B"O�����s�ԕX�H�B<d �"O֩���� )����M<*�p�G"O�Yɰ膩 �@���G�$Dыp"O��eGۂDĐ������>\���"O�if��f�z4���w�`�"Ojx�B	%(I���h�
 g"O˶&>d��[����E)I�y� Ͽ
���[5��Y,F�h����y�T,<]l�sg�7F�(Ŕ/�y"�	�)�	�	T� �g햩�y�m�#x::��(�`��c�O\��yA�_F��@����T�ʭb�Ɂ�y2c�	�N���!��\�CfFP&�y*�=�� ����?~��pɅAƼ�y�IUr�0C�m�Ic���܏�y⃂ �Bd���u�`$�`��y���!��d���q�ؘ0�.���Py�� �|p�D�X�~~R�;�EK\�<�E�T�H�p�cVs7�ȈY�<�F̛�3�,�#�J��2C!�\�<AK��V�H\@�H��o�RA�@��[�<��I��2���.K'\G��c'�Zl�<��C��(�ʌ��CO$Bye�q�<�ь�6I�!ie$,���y��B�<p�Q��R�D�I^֝��E͹!�!��>��"k�,u.���'�^$<�!�䍖?��Q�ɜs!"��"�P1!�� �̉`�B&�8���!�4c�!�dD�Y��1���̫����*�#>O!�d\#X�$(��v�X/�	0!�P�-��L	TC#V�M�!��P@!�$ޙiY܉i�7 Fv�bw)s!�$.?D��2Ŕ!4
x`����!��2.<�w�S�@��1��A<�!�$��hb�����N�lά��C'�!�$��5U7ʃ�s,ۂk:�!��J�o+���6!Ƨt�q�#ߢ�!�d��K��Uj�Ybl��@�8x!��,1YG��p'��'�N!�$�0B�dDq��3�ts@j��^�!�G	����&3r[�(T,!򤜀Y��#PHV�Jyn�8�s!��ݜab�4����m�^` ��S!��0%D����"$Up!�R��H!��>�(���C�+���b��>]!�� �	�G��R/���3jX�;(N�9e"O�\3�(�TlC�� ���(��i+ў"~n�	:"]
�g�=�Ȝ� K��?_F�OP����(b�lJp�[�$k�d2�,¯���^�� )0#C0�X@�I9uD�8��5�.�S�'T;�L��h�!�P�u� gBԅ�e�L5H䩞�6ǜQS�+t��Q�On���ˇK����93�\��"O�2��ec(c��ƨX0��`"O�q/�R�J�W��	?(֍k��'��	6 �"D���
-|����YqB�I�&>Lб�^�*�(+�O�g�BC䉔� |�DL�b%���'杗V��B�	�eP3 ��	���!�+?
�dB�I�)-^���)��drs�KR��G{J?%�2c�/�@%�ͼ+yH��g�j�=E�ܴ��@��S/(p�qw��X���D{��'3�ؓdO��QAn
?/�a+�O�����X"��mݹ`H=����	W+�	�<�J�ЦOq�j��"
�2 Ҩ9@�.��J��7�'i�!��؇dl<��{@�V$�D�MH�	Ex��)T�r�R���� ���P�DY�=�a}>iC�C�Q�p�ްf'��(Ɇs�g��rD�C[���iƲ����f���'h֐G�tcv��yu�P4���L��!�p�A�4D� *H#	�Z̲���-}$�P���T;�4��SF{@�;fIؑxR ۟<f�|*�c ��y��{��ѹ��U
j 
��3���y"�'=0A �O$PcPd2�I8*4p%q�'mڌ�R�*��k���*�����'m�(�P��=\�&��f�O�"�li��'>%���N+�!�ך.6�)P�'���a�/�<ƙ��O�z���L<�r�"|OU)� d`�L ����DH���Q�O�U"�c;S_�	�e�]-u�  	�'B���g� x�B�L5����O���D�4D)�6����	!#<!+A�C��y�"$�z��G�$l��D��yB"�3�����gdv��Ə��x��'�IZ�N�2-�&��Lʂޜ���'�a��ȩm�)���.춨���N��y2iLO�2h8@���<MA����yb��/�� c��	"��wI���y�nΥ#����FT�O;&�/W���'�az�n��`J�9�, BV+�N���<��k�*#��<C�Ӱ�*l�$��@
�B�ɣ.Ԥ,Z�hf�=5st�@!LO�X�>`�Wr���Z��Y�q�� 3',��<���&"˪EksLP`�jYZ4��y�<�U���(���a���Ф�V��t�<���2f�(����4H�9	ap�<��c[�C�,��W��0������k̓�MKS��>IO|J˟�m�!�����D#��?���q2������'cʽѥO��D)fx0��2Z9P�6&2�S��?�&j��c�! �N]D��"'ȅX�<�(ΕkT�E9��؃�|yz�	�?���'���`cT�Y�uNU�͟�L��� � 9��ۋR!����F�"���ȓyl��2�J0Q��Tj��ٰ�B����O�'�Z`3�K\����j1�$Xz�N��3��'����E
�i��\`U%I�O�K�t�Ik�����>�6�ϡU^VP)�'Q�:�ّ��o�<�!�4�0!*���<��ᱠ�7؈OH����(D��ɲ��ԕ5@`'%M1!�� p}z�C:*��p� ٦sH���%"O&i��U�I*(-c�\kB�����Oe���i�Of���@Cn� � ի߰w%ȥx��x�We�����̅Q��Ӑ�|��Z��-� �=���'o�S��?K&"U���Ucb��@h?+.�C�	���r�G5^��)�-�% �P�,�S<��}�pd
�M՘@��D��Z�xQ����Q�<9%��I[�x�HȦIx�����c�<YU��*k���AɞyM"I���J̓J̑��'�H� ��R�B���l�"ap�q�+"�Dܖ�0<a���MVB=��� eߑ��J�͙�<�L>!*O?%���1����BK�_-�x᳥=D�����.Z4���bLK��J��0?��O�Ósl$rG�M$r��"�ߑR��p�ȓ*����G!4Q�4C��H�<�;�4s��oDC����q�:�M��y��X�]��!�#&�8:�R����e��D�>��!1���fV������az��=	\\��?)V��d̮F�!��1�g��z/�9��$ma��"O��Чm��*�R��R0̔�"O���
®�@�{��V�t�5He"O�u��HGWwd�qw&^(g ��6"O,��[M<���� w�(��"O`�t�r�:Q�r��vO���0"O��b2�-e�pm�*]>�H�"O0(��H��L�&	���	~=0P�"O��r�;�8���E
�:-4�"O�Y��1FL�<I+E0E���"O���B�Ƹ4�b� H�`����"OFU�A�V���dȚ(���P�"Op,��. �q�$��1	�L�c�"O0�2
G�z(`��0�����"Ox����m�`4���  �^E�!"OD Ys�ԗF��5:�A,Z�ne�7"O���� J�;��4����*�z��'Nў"~ZЏ�y�ɢ��

k�O-�y�Y�">�b��S!_lTS��@�ybDPn>�+���eϚ���"���0>iM>�dn��-J��q6��/i��H��^�<1���?)d@`Ri�)`���@֨K��hO�1E{��Y*T�kbg��k�Z1��+����m6Uis��5!���W���{� ���$;�O:�PCg]DRڅc�,̏e�t�(�O���&_^����f�3e;d�"D���,�R��R$�t�S`�!D���W���!Y� �wj��/�ȱ2	�''�܁��� C��!���$�C��hO?���5v��S#��5@\� ��<��ضT�<�t�O�,�	��NV{�<y�UC��<1�BJ$��u��5T�X��ث٢a��-&�|���:D�`���{�������Tlf��i&D�����\(2�`

Z�t���8D��S� �@߼�I��l�BV�:D����A�;pZ��dȉ�C������7D���%�N����wd޹rD�4D���q�G�b#~���N߹}��1��M(D�`� nO�`�d��-�{�l�� '&D�̐�!<e.hb"V
U�h��4�6D��1�"�:b3�AT�y��\*g�(D�l`�`ӧ��|eb�m�R,S�*O�]I��0y����Ǒ�Ȣ@�"Ob��RL��NVi�էK�1�\@YP"O� Z�2޴bz������o�^鈲�'��/���9�G҅@Y8�$ �27N��ȓn������ ��5�C!��l�$�ȓfy���rJ#"��F�$|MB%�ȓM��`W�;4��kš�
��1\L)zr�\+J~�y��!E�cȶQ�ȓN9.Qq�Ƶ�d�W �#|(X�ȓx�蕸���3�2����$4t�t�ȓu�x|�'Ý n?�h`w$7�i��yGj<3���.vH��v	ʞ?+�ԇȓF�F�SݺV®u�� +�1���T��u@�(r�͕�[�]�ȓL���@��s�I˓��
j��ŇȓC�Z�J@a[*�J��� Uin4��l��Au�$<�-�@F�{�rU�ȓ	���@U4O���%G3�ȓ0��pQ��2y��U��l۾�m��F���(Q"��(��=��l+�h��p��|��)Eh��:�l[$��@��v�d�##���X0�D*��Ԣ3}Ω��V.8 NJ�������Q�i�ȓ9�.D�s�FZ�4�F!��jk`������ʦ�Ė{8�A�D/[�4U���Y���g�n�Vcؠd:\9�ȓY�Ju��cٓ-���B�����b�(0����!A�H�p��1�K�<D��9�F���K�/�$��C��J�<�T�>Vf��ad�*�<�k�A�`�<�&,8'����.	��ࠀ��^�<A���%*2�#r�� �)X�V�jąȓ������KL*�!���L1�`�ȓ%�ֽp���$Nvyat%�,{�*�ȓ:�D���d� �Q�mơ�ȓN,�KE�H�<�0�"*�|�ȓ�α&ߟh�t�p�@ԟ!8Ҡ�鉷M�~��
�fNH�n#�Z]�i?Pn8C6ဗj�FC�	�xT
��􏛑<�D�X �ŗ,kC���`6�V�I(�C����B�Id�Z�`�#d ��^���C�I	�!B)�6&&أ��<<2B�	1$�T�����\��̂�e��C䉕/��iuH_� $�1��>	�C�I9Pv�:�U�I(x����0DzC�I�=�"Vܪbep�K֣�a�B�I��T��X[��2fiԅ:��C�	��F��M�>E��:�cH�'��C�	��lX$H� �)$�ʬj�zB�ɐ z�hp���=Ghd���F
nDB��-�&"`F��l0�3��+ �ZB�0�$��H��p�����i�n|C�ɹ.w������0p>��Q��V�8[NC�I�h�Ѣ�=Y<��!AmT�UZZC�3=�5��F?�F���s�6C�	�!���[�g�8���[Q�Ԥ	�C�	�&u��*�E�H���x����b#�B��1�A�0�V9X��d�%e]=x�B�	�]V=J��ѕ�p �M،L��B�	!Pu�yP���f�ba`t��U�pB�I{��� +�M�z9�U�̞$;<B�"���g�P	�2AK1o7�C�	+.�3�nD�>Q*�@��8��C�	#txص��=%'��Xr��
]'�C�� ��YH%N�8,r��C��C�I�v�^I:���bU�]p�	y74B�)�  {�!J/)B|�!�XTR�0w"O�XTG͋#7d�HR�+]^�G"OhAP�.�7 uz�H!� ���%"O.��
Q��e�1) Y�f�z�"O&��7��0a�9xC��ɪ��c"Oij�D @��[�!�'I�8P�"O6�(�K�!?�ě��]-���5"O�����6%&�����i�P+�"O��oͮ2��q���K�GX0�F"O���<w����Ɓ	*p^b�QW"O"\Pw(ͦJ�Q�� �Qd�S�"OؽFk�4�恊��W�'F A��"O\�"�f�2��I���$$��"O�!a5��$k{�$��Z�O�Qz"O$����*"h��qԎW����I�"O@ XG�Ø�0���+����"O�P����ݶe*d�Ӧp��h�"Oz�C�.M��;Q��('0HI��"O�h�� Z�:bb�Q���X� �u"OJ��/��h�`��E����E�"O&-�4���0��4����.i�>�sQ"OBTx�c_�>8PZ��ګxd�Q�"OHd�u�ܗc�4��Ao�B�� �6"Op��Q�۸1O
���N�1��}ʔ"O�*�N���r�{��ʬ�Z��'"O �����]�H�cю�}�<ms"ONX����h͚��*L$�!��I�8|���%��TT-9��]�oq҇�X�[U�|���<��U��JȕD%ƥ0�6'�B䉦#W ��-~8:�f�+z�On�x��`�(4A��d�#f&����K�i�x	�G��<F�|2�_4{)��H�!5���`�;9�v�H�b�on� B�[�J���	��䨲�qD@@xP��).V�<A�������rM�pGFL``�
���i��]����F�ή�˵N� !�d#o��!I��K���@�왿�9�&��"f�X�t�f̖��	��o�Q>�����II�邬Y��Eʆ�E�Lf!�1(ƮI�ж�YzT�#LВHp,X�aӦx@�#L�A��T�Ʌ������'����b�.`���#3h�@�r=*
�i�5(�5z���+]k����$u���h�-�-C�ܩ�V�]�O�xͅ�	�E�z95,C�um~y�0�Z.?h�<�C�@�n)i���venY�Nڟ,;n�R\ws�D� -�_@ĩ�Mnf�M��'WNcB��� �zWʌ����wń2 �ӑ耮t������|PB(S8���$�!U�P @t��6J50)�"O�%�3N»>��<C�+f�-RT���9�4�Ӄ�"r4��R&�� @>��vd��=9掐�H�<2�A���"mx���6bۭa�Yc��P�]�<�DLW���*ƮY�B�ջU.I�I,� -Wz�z���qh��tnκ-�,� Ř���O���+��vx��A�,Ϊ	[B���K���@�:f�\���aR}t���Iu~d�s����Js��h���wI|y �j<bb`<�'���c�˂�Sg�-cÃا=ML `��{�'e@��V�։I�8PR��C�2��'�J\��f����zB�B*F�l C�W!O��1�faH� :6�:���1�r	�d�߲m�,rb�ª���P'r��y�����FLU�Y��z�ʊ�9��D(j���?y�ثk��8�q.�3�5Iv��>��Iq���%B��[�`�>�c�MP�!�8����}�'{��� �0H�O� ��Wj�g��(���ɇC�dj�H�=W8�ӕ�Q��Q���#j_���"�9%V��#��ĸ-�v%��)}�sB�<��Z�r*�Tx��.扯_�T	X6/�<KK��A���Qʓ]� �G�1MlR0��/S���e��dr����zם�t�,��Ã��z4H5{��ѽi���ɟj�ہ��W�az�ě1@������I Zj�Z#pD�9;4�J6�,�� ��2+�h!D�C����-�V�!�9#ن	�c�3���B*�������t��@;�#����]�q�Bpo;2c�P����]�uA��(��s����z8j ��L�q
�r�O����CA/b�N=��]�T�#2E	5�d���ɤtJFu:��	�'�f��E��	P�(P����$09������1m̥��Bo�mJ#�I*}Ҁ1�V��P�,RCF��&�(�"�p�ɓ(�R|)��3A{`ʓUKDQ�� �������r�4Z��Vl�	1Dsl8�Yw�51��lB(V�d�a��<��I�'�z}h����<� |!r�V'&n���F.AV؄mא#lqA�F�J�d�����K�r"���$	ƮG�S�<qt��0t�T�[���n?�� ��%F�~b)Q c�L�LU�0y6��s&B �۠nϞ��0�BPy2��U�V*�D��|[�lZ;]��a�?kT����M�Y�џ4,36�����ͫ�ħ_�l8���I�|�����
�'���%/�$�����M��?�`�f�cG�s���ə'^�����)����Q�*�<i�/�<���1}��)�'S�j�Þ�(�I�gD_*d��Эu0��A~A���剷J,�:��W|x���N�pq�L���2Ǧ+���&?���G�sKZ&
��q&���y:�0H��,�Չ�[��|��V|Nm�ǃC(x���bG�X;e�U'x�'F�H��%	r,���)_�Zv�+��J0�AsaE1v-џ�	�	�\�>q�p����;?�|���*��C�M%�M{��׎!0�Lh�^~���isf�1 �)Z�ؠ93b��0h�)Olq[#f�;X�H��|�2"��$;P�%iG-Wk.%�0�r~2�X��LZp�'s�1�1惭8>U�`�\��@Bc'=}�aܸ)�5�����O`j'���:0��Y#V�}*��X8�p�
�/�6!`�g��l���͉4��a9�cC�Hr����� �OV�Xd��`D�<���&Y,�t��ɭFm�邤�R��O�b�i0�V?��4�&��{$�	�'��ZA"G�G\�[���>����O�$��lY+O~�O>�+A%ȵa��Uc�ԁ,.F�g(D����u��(W��9l�ᓤ�&�I6b��A�Q�'�*�p�&�GL\�9�͞>	΀�	�'@Zt)!eѶO$����bD�� �'{�Ǭ�v�L0���?��M�'bP��,F9
.4���V�e��d�'a�1�0o_2�s�KW�X����'����
.H�@�d�78Ɗ��	�'-���E�P"D�.�af+1欀�	�'���h"��\��@�s�$ �"O�8��R*���`�,P��"O�m���6R��˄�ƥqֺ��"O���A�8VXT ���!<S|�Y�"O*�:u�Z)%L��T�Āy3"O���7��+D�\� `�-P���"OF=�)D��H��V�9�>H��"O��kP��MC��� c�8چ��#"OX ���,Bp�"�".�R1G"O�D��H04f6a��)qs��@�"ON):2#�3@n<���݌SP�d�"O�u�6��*a��5{�-ٯp^p�"O����oA�1'F��@^*D�P!P"O>�H��^�S,H=����>Ա�4"O~$����/~"��fƂ�E�< �"O��SaI�K,°ڄX�I��(ܾ�6��i��Y�\c�H�6�� �P�H���	4�-D�k�OַV�k�F.��5��ͱ7�bqsH�g��|��]�tʷ�GI����V��<	�/O;�d-1e��!����>s�r7�i����'�~�!��D�X��QٕzI�]Ys�Y/C��)��(��F 2\���('�ߵ�H���H��Q�0�z�Z�E)oj�<�"O��!���u6�e�I,gL��1�Q���{'����j��A9�q��'J*��%�@�
��%�"#@�+�d	p�'K.���R<=3��fE�����a"K��"ٓ�C�mA\��1+�h��|*�*��R7��Qǆ7H��`E�>O���-�>?�i"'��*)�6[� Ǆ'��[e�=�x"3PwE!򤖏I0�R.\�T'P)3 \��	�q^X�xńM�qwf]�e����G�$O�)8�� "qO�f����W��y��
�}�&��è��A0S����gOC9:�B@���[�"mI~��y"��c"���@�Ӗ�>��FG��?�^'`>$L��Q�o�,�p
 �6�`6��FAɀ��A	ӓ/0��7�E�Cs��A��3Wj�G§ށ���"��a�t��Ċ|j5Ȥ*Q'L�Q��Al(�Z�"O8��Sb҂
�fx��$���<��^�p���ړx�\��ʸ������g�π ��a
�>DΖ=q�$�h��Tx�"O����J��߬l�5��N�ĳ�
މ�0��m�'Y#��`>.��O"1OB�I1AWb�ۄ![v����'{F�aQ�Y-�����ȍ+y�Ȱ��C!dy����J�=�Ș�)̻i<az2i�&��}�r�7|˒D���-�0<Ivo�� ߬�V�˽#`�����g�,���I��2LD�һw�I���`��#͆�+�u#ӏ2P+H��'V��f�`�N�0A Uz��D��l��7�~�K!���ty��D��y҃U9f�P��!�){fV���?
5L����$+ �D�RK�ᓈ�L>)���j�����ʹ)f���H�F(<�ō��p�i��J��=����Pg�|�	��[��=�D�P`GL��w��?r��K�OCX��j��}��5r�(�����+��b eJ�ju2Y�*ݾ�y� u�"EA�=>���D� ��'<:���$��
DD�dD��r�	."\R�-_��y��V'[s�P�Cl������Dt�%���\ܓ:Α>�^�`��2���q�:�ӱ�\�|z ��\w����͇F����c,�:_�L��ȓN\���2 ԋ��5�ɘ}����m�T٪��؞cAq�h��������!I��эlǮܰgj�}5
���ڜ��w���]�6T �J�<�j��ȓM������M�=pL�&��݆�XH8!s�#�$-h�(��A$) ��\8��0�&L�}�)emU� ����IN�{!GG=#��Y�HI�3HB����bգ�!�%�����: ����)�9�� Ͼ82��7C�h��V^he�U��1	P�Q"r�W��Xd�ȓ!��	��G��!$'L%iż9�ȓ� ��Y�;��6�T�OV2\��'V�=�`)�54�j���i3C�J�X�'a<� ʎ���
 �
���'���3�X��u�
����!�'I�\�Ձ]�MC``4\+��[�'�c��Ho����	j��
	�'f\e�X����̎xe����'�,{s�U
K5	a��вogQ�	�'��!2ֿ1�~�c�lۨc�.���'��tjP ��X�.�!3�ޫ^��8@�'�v���M�*ffNt�CN�Snd��'�B��e�>Ev�sl����I�'Q|p��4$k`9���X�F5����'�ruq�`[
�h�Q�.��7j�y��'\��i�ρz�^8s#V))U*�'���s��]<,� j'�·$g�Ԣ�'�� �d��>����6��WC���'��q���Iv��LiX�'S�@Ys�!y!�U#]"D� 4
�'.V��,�氱�4l��Nk����'��҉��L���H�6�Th�'#���dזj�R�J���7��U��'�v�ʇ�Km`|S�iH�g�`�'� @F�1�d
�(�Mk �a�'�t���ֶwn��@�ν,��p�'�8���H�'D�@g��v�#
�'YlE{0��>. 0d��3
!�`
�'@p��
�H�T��4a�� �8��'�4Q�0%T�k�Аrԋ[.�Z9��'���DN�-F.�+VfU�J�'Ԛ� 	�Am΁��k9�	`�'��nJ;���C0�J�<��ݘ�'���Ǭ;�Pp[C��2����'�r<s��j��`�"��2�
��� �A�
�qIZ��G
��'AL���"O�����MR\5�P;
Nh��"O<�����/MƬոdF�J)d�h"O�t[bgʀ I"��`�-+�x�"OX-xP) � _�X�@dU�7@�w"O��	�2�yh��W;�@��"Oޘ��e�>&��c��F+*��`�F"O��)g�3�ne��%�Hc^�8�"O���E�*����'��9q"O�5 _iW��q����P��jP~�<a��˦cX�$�2��mqo�t�<� �	/%U���g����#�_q�<)�
�5/�;Ą�f��)P�/G�<�G�I�\y�́a�4�cA�<Y�Ɖ#2��I &䝴0:Q:��|�<iA"̫}�A���7��l�΀x�<�'�čn���z`/�@S��	e�|�<���RK�,:(��� �D�<����T�\[�H?�\� �B�<Y�*@�sI����ǻjr� p��U�<!B�ObA�֨_�F���h��L�<y�!	Р�hх��l�v�<7��0�,�J,ax�3�n�<I0��*�|lsnD_���{#Dr�<9c�"����+/hRT��L@n�<��O��?v8 �4d-ǀ[��So�<���\1F�Ll�k��x�ıå�HA�<��X�u�gd�*u�D ӑF�C�<�&W�V�87&mv�c�&�S�<!̉�pT�H��n��2�l���J�<y$�Ϧzr&�����N0�ݠ�Z|�<I'��`����C9�t)�� ����ppH��9J:�$�"~F�6鬉a����X����=�yr�y*��Z$�*?Z4��L����T�"�^MЁ"A���<�1' 	d�����l+#�U2�o�t8���	>^�`�9bC)H��ɱ�MȘdta��H�1�2��ēAd�YC2��*O}�9���"�b�Fy��En�q��+M��vd9s٫5s2�8��#x��C�"O�DMԌ ��`�7DZ���Jġ�c�P�h�O�zD�-����2�W&t��M�r�I"LvxvmI�y�a��z(8*�Ń�r����P�~ba��+��PP#�.�ayѦA���0�$�%fC���#_'�p>a��H�z��u ��*�]bUdL�T��ԯ4l~��	�'H}��ϛ]�pp1�A)1o>a���M@U�AΙ^�tb?ɐ!�ھ���C
��`b��3D�tiS]�E�- �\ �C��<M�u� R�T�
*O?�d������Д=�T�H�l	�Z !���N��d@���z���+~9�O�-��4�j���` *W�h�ɠ�`Ϳ:�@ܳd�'�DԣDM��K�4�H���(�L	X���z�<Ћ�"Oh�������{4n��mK�Qk �'�H����37�V����$x�T.�
ynD�I�;B�XX���5��k���`��U����,*��F|�&qYC�&�(��O���ia�	_�BըeL�Q�r�ON��D
,a����$�r��Ac`�T�h���H���]5�{��F�,��!�h��s��O��	��D覽��#�8�x`� ��c�G,��ڳ��"w�J�҆��E�\K�"���<J�JĪo�~�j�@�A"�x�񮊡p�Z���4���f�9Z��D/2Z\���?%B6i��Ǵƣ?aQ��H���p�E.� @xKv�	3CL�"������ �
�{6GQ�3;��pbI��y�Dp��8�C�j��c�ЂŔ�mMr��PE�>�{��<ف�Bt��pk4�ݾ. �HQ����$TGk�@���� kݑC�T��b���8��������Ҡ��c�d�Y��'7X:��Y0�#���8D��A�"�E��]q�#��`Z�3d-,;@,���?�ݠl�,`鱂P�($Z�8��Z�0� �5�[i��
*#N�T�.X?h37
�'�S�g Dn���×�s�P�(BAO9fzZ)84�K�^;`WZ�4�4Js�7� f�@��4�I)�!��$|@�W�	��d���*H��A��(Z?�m�2�o����<Ǌ�1
�(G���F�ќTE���W\�L��6T��B�>�%-��2f' I�`�w�ބ<˓`(I�ߟxZ6��D�x�3�l���E�O�%
`����6)�҉O�:�2<���*���6O� �c� mS.�b��!<O4��DE,�<JR�ݐM7E��%���"1�A�%V�����J_(��l��.���u�Ij��넭G�nk�-�S�E,/4p#�lF>�p?��o����MYw�O0h�|m���@k�$@Y�tG���X�d� $A�bU�!����#�ħBʲ�#s5D�@#�F M�u���U�'�V!�X>�&>*wi�pW]q�gA'z\��"�N�!p�Rc��Q0q`��O�	\�AU��Qȟ�d�>��y�AƝN�~��L�6.��uH(}�Մ�2��S�O7� �C�_�,�J}h����pX2�'��-���U���� H',O���.�Ew٩���7faR��k��C5h
���`/��4m֝�;AF�1�柄d+X�q�z|�Y�b/2j�����}����+T�D^xQh�&'���1�S�,�N�[L>��/�Z�dE���O��a5�
<�H�Cf{e��e�'�WƎ��c��2a���<1�e�O��p��g�#q'B��ig������u�Ds�O?7R�<�ʽ9�+�>i���Gg�?��I/n+�f�KH�S�O��!׾�E(��1�Z����g~B �.g`�p�'.NPPn�8i��ı�K%_<�1��$}BmǖO�`����O�Ģ�� ��S��"CPv	��Q�]dZ(�
��+�1���D$\rDȱd��.$T��[d�Q�'2\d�e$�O�9Y �V��A�!eT�1jB2��� Z`�EXw)ƕP�O�d�,0�P��U�V��tMi�'u��1��+<���*��:7pX�O����v&l�O>հ J)`�҉�J��gr�d�;D��p)F9S�&a��)Ȱ7  ��+7�Mȅ�'��y���Pw:)��� ��p�'�Vt���5��L $qZ�l��'dv���KT%?H0Bѣ�_�hQ(�'�J�;P)
c�|l��GD�~�P�'���� ���1|���Dƭ�%%�W�<��
�(X�}iSL#0��iS$��y�<A�^�>4c4,����a�I�x�<��섚\\��YS�Ԗj���Jh�<6"�H|��a!��in�E8���N�<���:�,�����<�D��`A�<)Qըh����`���.��D�B�<1��ܫ/|�9�!�5oSfx�q�x�<�F��LZ��E�D/�6��AL�{�<�WξA����Ɨy�f���"�}�<)���C ��K���E��{@�y�<!�C9E�xr��[u���f�r�<��($�:Y�_�EZ�j{�<��;,� ��;"4%J���X�<1�O�>������A�:4H1"�	Y�<I�� 
r����l�z`=Z�gNW�<�&F�rd��h��:y�b�Q,�S�<1�i	�F�Se��4}�����@O�<�t'J�:]x�ǰd�DuɄ�P�<At���fN�+��׭Dp�l�ƫ�k�<Ib��B�(���+31p����x�<�&bH���"ή:��MB&�B�<y��_3v`n�t��.iL��z�H[x�<f�#y"&�B!L9��|�<���ޭX�%3����l4z�y�<Q�%]�Ɣ v)R���\����v�<Q�]>ob��GG�x�.�ǃ
q�<A��J�z�3����N����7kXi�<��ٶ�����$2��(A��i�<Q� �[����Z�j� _r�<��'��ҹi��!#P1����m�<�F�3ڹ�6�հvA4XK��d�<0/44��`3�
p�z��A��f�<���4�b ��&�vD����J�<� ��
G��!ip Y�s8�'e���N�KX�h�b씎!���0�L��;�d��F�$lO���%�ԭp�*��#k�dḊR{�=��@V�$�NB�����sI�
8���	�#T���� �A�_�h��V�o[<� �L3�4x5��1J�C�-��D��-�39Fx� 瓝𚨀R�M6j�6�'�-E�,O�P��1H��U�䃁�wt��0"OȌj���j:Ȝ�g�ѭC���C�L(tx�|�f��}�a|"!��c��M��+>k�0��T�G��p=�/�6
�*=؁�x�9t#F&x�N�B@�Yu�Z�� a%D�T{��Z�5<~��х�X�ٱG-��ܸc��F�?�#2�U5Q��8!�u��� 4g.D�@��+�ʂ�����2�x���6
��y�l(}b�B���`:z� 0DX�v`x�B�Q	S�!��z!Y�P鱴��9���A�_b��U��JZa|�̜�K�l��L��Uʳ���=)�)�4H|޵�'Q���5hKz1dL��g�"�¥�	�'��a���-�%��-O�^�q���\+7, �G�d���'\���bƖ4�|3!��!�y�H�������* �M�y�*߅H�!��A�v��Bc�L�<ٰ
�4=������O��qI���}�<����+9�R���,G�S��а�]z�<�D��!"�\��L�[��0Ɔr�<a��>l�	j��ޥ5[��P�)�s�<ycOZ�[	�e����)?��p���g�<�TmG�~���CρAɮ|HN�k�<)��&v,�AV�@�G�j�c&�	{�<a�JR>lTU2i(Φ)��oPq�<�R�
�V=�bGDROĔ���g�<���`�j0Q' �#"R��t`�E�<i��D����J& �D]��NAA�<I�	�l��-y`��&�����d�x�<	"�X9*1A� :Z8�Q+Ʃ�o�<Q嬘�/LdY�alL5~yڭ��N�h�<IW�`op4����7���D�R�<A�&	~�
�`G-�0 ���T,�u�<y�s���;��Ev�s�<�A`_�v�B�i0�P:(��Ӧ&
`�<qď�5G�j�q4��8N6np�`.�G�<���O5�B�PA��ED�פA�<9ue�9�@d�ҫ�4��ax��U�<�u�$�j���*���"�Q��4!0��G�L�f�-T">I���6i�	�k�W�  ׄ'D�T�!��x\�uc@ꐳ9)���Dg)D��i�!:��	[���/�-"sH#D�أ��˷%�
��c�x]F���g4D��A�F�(g.���d�(iZBIS!.5D�B��=�V��5�V�Q�EY�5D���D���;�p��%o�`���>q@��W��H�<EcC�T�M��hBg��X�,��imJ���R��@(O���T��DI�W��7m�(h
���'%U�]�M����z6����oӦ�"�����ԧ���	-vm"u�AF���q��e{r瑦R�"~*2��I۴����R�@:6휖"B\�Ey��	ƻ"���AI�1�@��_�zTQ�P�W�O���3!$��B<���gQ�7^-X�{��[���'C�b�'���b�!��U.1�O��ڋ��i>a>V4��g�)|l�u2'�����5�hOq�����r$|��E��t�A��1U�b�>�O'dc>a0 ����)���=}O8A*��4?�CO#{��t�D�/}�𩈣s.Y`g�ϟ'���hL:5��f�������$P: ��)�p���8t�\&c<�y0��S�L�G�^C&�a:6�s��8u�{>U��O��~4�۱�̥mE�3Q�X�&��W3O�X�F������	[�@���mI-1^z)�o��s߲a��hJh���kY�������� |�bR���Q���]�Ƶ�3�'Čĉ�.�_�S�O]�\�ə|���1���,!(N�����5>���|���.u�`m�<Z��hC����(����{���Ipa�DL?,�ر`�`O'h|�z�̉���i~�r��)�)k�.��R'�L9@�)`D�9�PB�I\M�x�!GB X`�l��FCBB�ɫ8^�:)��pW�m��^�lB�	=�P�B~�������b)B�I�aqrk�G�>[N|��T/�)P��C�	!�F���l��0�'��_G�C�I�e�$�¨�<����É5JjB�	�C�Ҕc�g�>��t`�R�B�	}���'ŏ)��5�ņ��c`B�	�{ǘ�ٵ.J%B��1���\~*B�I:m���W��O�h���_,PC�I�%֨ɐ��D�<@(s#'�3/"C�	kB`��H;,�$��	cUC�	~<���r�E
?�P�aQA�|N�B�I%N�<\@C�O=p�zm���=e0xB�	:p� 5SgNӥ/��<�q�Z'{�0C�_��}Ad
iF��w�Y�?8*C�ɣ*H����*�J�8�&>@5�C�I�_TQ`Gȓ�Z���Rӂg��B�	T���e���,���,]�OtC�I9~���h��C����T0DC��zJԉWΑ�H���b�;J�@C�I>#D���H[��"Se��e�RC��T!<�5K�^����vՆB�?{�9�� �4r0��*U��B�	��0�"c�|��A'J�&VrB䉒F�I3K�I�j�jpe@0sddB�	���躅	3~�L�q���}S�B䉫wY�Hr*߉k�6d�m�1ѴB�I"g��K���"u��{b�Z:6<hC�I����n"��]�1�vfC��t{���W�ʎ$`�QqE��,4C䉯F�P�Q���pi�p��?�LC��&-�` �Mϊ1�4٘���y�.C䉟^-6�@�įq;u #��dIC�ɍY(��0�9O� J�ˋ��B䉪]_T�p�� Wm���q�(B�	�H�S!��[��a�4o�(B�	� �x	���	i�0 ��6q��C�	�0�<�+�J��7��� 1j0fB�0�t� ��5R{�ݫ��P.}MC�-"�B�)[�ta��b&.��B䉺4Q��Z>1�R���[�|N�B�	�@=�@+���1XH%����?wj�B�	3�ޑ��N�J����/��B�I�\�B0�<P����g��B�	%�l���ɾ �n<����1O��B�RE��A��T�mJh�4�̬w�bB䉘E��e���_�6�"tÅ@L�C��2\��Aq��>Zjf�o�|C�I�L
"�jq#8���)c̪	KFC��''BF,IǠͼ'�z!��\g-C�<G��9�$Q�v.��� \��B䉸*�����X5� P��M[�_q�C�	�H�T1�H�@�� xT���d��B�ɪJ����%e;aoL�rW. �y`B�I�ӡIW  ��P��X|�C�	�d�0��c� �g�`���ͣM{B��sHI;�J1�T�*���qi B�	2a�^���/�!7H* �u�yC�)� �yR0�/d�ܥÂ�m �!�V"O��R"_j�&���'Șz�%؂"O�P����S�"���f��.e)A"O����g41t�I�rE�h�nTAp"O T$JӦ9�2���#��X��"O���H>u2� N�T�T�[�"O:��d�^�!X:�Yf�ɀ9�P� �"O ١����%2�����r-R�r�"O�yB����N��#hԴ^����G"O��Sm&`:�b����H�"OXMW�E",�sg̉�U��@��"O6%�%e�(^,��`
K�H���%"OV�IPB��@�4lkd��1����"Ox���K(2�`�ڕ��JV�`�g"O���󈄫#r��gk],n��5"O��#�in<X˂���*���H�"O�I��_=<��aJ��G>@���"O�LYrI[�#޸�qe��71��98�"O�<��%�[�D��eЖ? z�"On�#r�F�hH�Y��^34<��"O(к�lZ]�Xq���Ĉ�6��s"OԬ`W��0 tH�BE�J�F"O�8����%<�z���12jļ�q"O@À�ƤiU�.�1,2� �"O����ѯ%m�BV5I�y��"O�	��c�/f_����8A��z�"O�H����*"+�9P�"���t �"O.�����E
�9bF"I� Y�V"O���*@�LƖ��!��zW(�{�"O��x��c~�����0c�l5�"O ����v����C�X,�1"O���Q�)I8�X��-5�4Ń@"O���5G�o�ųe�u�j�"ONXv�״_K��;��D�:h��Y�"OB8�6 ȷ)s��"�(�iN�j"OV�Y�S�I")e�̉o\mC�"O��� �0\���T���:8�/�!��B� vЁ#��(����!��a�tp��O�0�ά����8�!�T��:,˂L��	R�I�!�$���<���@%h�HDФ(װz�!��*��)��̐Z��cQ�ё@'!��Ê|��L*Ā�7b֌�Q����/!���)~�ˀ�Q�0k�>!!�x�����C�I�RA"P/F!�zKnl"�}$ъ6����!�$�14#��X�!'8b	ru�P/C!�$=
T�x;j�6Q0|��ߩB�!�߱��90��.}��|A�4�Py�E���x1�N��=z�z@Ԝ�y҃
9\����ǎ�1Ҧ}�m��yr� 3J���fލ&�%����*�y�+,� \�%�$�:q؅�
�yRQ��	�L1~Ezu ��yb+ػ�2��T@�p��4�I�y2�P1m�P*�G�r�YBT���y�I ,?����8Yu�@�C+�y"�@ �U�"�$XZE����Py"��,lF�#�E�Y�������S�<�d�N#!BH�EK�5��e��@�M�<9���]��β��X��K�<Ɇ���W�Fux�l@+6����O�~�<�DNY.`��ő�f	�K�z��I�y�<gH�B��9�,:j��YrH�L�<� �����((°b���#Z7�I6"O>=h��
Y�!3WjY 1>�x�"O���E��:�4�G�!Z'$e5"O���φa�&E���!�m	�*OF|�n�T��%)���K�\X�'A�ʧJ�%)8Ȱ�Ƒ&4~��'�����W�`|������Q�'��x;�@�l����g'�	
��d�	�'�l��ЃZ�V��4'�6���S�'bh�!�ț`x�I6+Q�0�����'�q�+Ee�� z]V(;�'����J'5���lo	���'�`%��X�ڔ��Ya�����'����`j������
T��� �'< yk���:	#DD"�K�0��
�'0�u��$�K�H��B�M(�o@M�<�wb�	Z�dd!��6]�*��T��H�<�4��B)��g�	;Zk5�Ec�|�<��B�T��P�s�C8�Z���Q�<��$KA:�Ȓ֊~�X\	���N�<����p�=*�Q���|� *VL�<�7ˉ�9`�S���Q�O�<a%)�'r�
�aٛa�r�E�<a�搐)x�1J^�%V�II7̀Z�<)�I�k4>`3%�Tp��� d��R�<A"�M��x'��R]B@iqiBY�<�p��9W��a#���|&�}�s�U�<�c�AD�%�b
�+�� �MT�<A"��*��#���#9�l�k �.T��K(k��X�ժЛ_G�Aڶ�(D��p������ӑ˜p�]I��%D��Z�`E�~ia;��=R����Q�#D��ZcfY���;�!�	v���s�"D��S�* <K����JM2�hj�#D�hy�g�u8xͰ��	+u��e�?D�����."�&��B$ǔ�y2�=D��!g@G�Eon!�׻2�PH&����yrG�0��D(f�ը~������yB��c����'
�R�)��X��y��˟��� ���L�}aa���y�`T�b�*$sR�Ĥ"yִ
1���y��4:��h+���I��I��J��ybnH�¥
�;E��ݪGƑ��y�#Q0�S

�{@p���0�yc0%ṑL8_����i��y��uE4*ޔ�s����y� �*`��d��-HLQ$%�.�yRk_wk��S2b�̄�ق���yB�:�xd���򈫂�y"#�i�`$��O9|����&R��ybܺ6�Ќ����,��X��喷�yRi��R�p��8n5L��r���yR�I�q,�$��Q3p�@��J��y��8x��dyV�ȝ<(��Ф��y��Ʉb �BRiH�58������y"i�����k��0�q�/A��y�G>�͐��[(�5���E�y�ㄧs�:I�v��Od���ʟ�y2��-�D��@��I���(�*��y��"^b����؁luĠ�	��yg�D���C�ǘa��!:�	T:�y�f&|�@A�F�Mz�ލ�y��+eR�m�.� $y"dT�y�%�|��Õ8Q؄�q�!�y
� ���/�F�b�2�ʃ�O�a"Oj�Bb�!M��$��k.pֱc�"O���,�%F�`1�� �Rk��"O��N6al��S'�Rbj����"Or���B+K%H��BFU:�j#"O\`QA�3k@q���!oҔ�"O�m"���p/�]iZ5V�!"OX�j"C����E7H�
���"O�b�	   ��     �  �  <  ,+  r7  �B  FN  �Y  �a  �k  ~v  �|  �  ^�  ��  ��  3�  ��  �  K�  ��  �  $�  m�  ��  ��  =�  ��  ��  &�  @�  9 � `! 1 �: CB �H �N /Q  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;���ē]�.�X%���tM��aF��m���d"O>P(DǄ�.���w�G�AB�"O��UjGOV.mI%�]8Z�y�"O$X�Q��L�"c��=�� �"Oe	���0%�^���a  )�6E�c"O������r�ꑺ��O����e"O�%+�CdeM��1O.̩G&�eh<�E�ߒu��P�L��SF��h�]���	@X� 4d�N�F<�bi��E�Uzo+,OpR�O��dW�e(�EGߎxB��ݢqĊ��ȓE����E&6zn��8$$$��A�<�<O&�s��E�π �Y�P���.i���x�ЪF"O�)��B,]�X�S�b	|9I�O�=E���7` 
`Ʉ�F/e@^��G� /�y����`1�G�A?]���A7"���y"'�XPq�'T �W"���>!�O6�zee�82q��[�2f(-�3"O�a�b_b����E�Ie6|��"O(Q���r�F�A�E:<�|�
�'T�9A5f�cG.���ZS�bU�'�^�Ӕ����v!�'O��Y��'�����$r�LI`f/ˬB�ڡ��'���vOSNxX��d� 7�(���'�S#�$]墭�t��>#��e�'Z4݁R!$(\���gA	l��K�']b�qH{�t��gӣi⸋�'J� ��-�J�Jw.��H6Ű
�'F��	&E�J�K�e��y,�9
�'5 ��uoV��P�
# RA�:��'��-;C�P ��hY���3zR���������9��3� H�8�Gh/D��aO@�k���4������Ĩ,D�`T+��QB�"[Jh�����+D�X*t��(^�R���F),�%a��Ot�=E��C�#���IU���] �E�.G!�d��q�ɂ�!�'�~��Лg0�f����G�U����9����$D���S��&��d&��ɕh#D�,)��Q�4�(�1.�BG6̪�@ �SK�#"G�_�F�zY�#��+L:���IC�<9���@Z�(� bU�x��!�K�w�<fET[n��#��B8�����r�<�p�B A_����Lԃ4J�e�w�<i��gM�L���;?��P!���o�<!2�L�.a�3���EQ�P)�ğo�<���S i���X-/l�����h�<ѡeˌP}�K�o�(Ejt�����Y�<2mX7#�B�G���&�h%s�'XS�<QB"�v�J���"E�RV�L�A�VN�<i��J�J��� �M�:y�)X�Ǆs�<9���"h9��̀$(���s��p�<)į	�� i`g,���N!��_l�<U��Xۮyp�(?1���%$F`�<��d��*�����!��b�~�K'A`�<a�D�E������8���C�PZ��{��y�Q�KHtʂ��&g9�%@���x"G�����͌�z���mO�rO.t�ē-��ɒ�G1=��Z�D�9o�l%���w��`���T#�1��ܰG�N�]7��ȓ�TH�Jð\~����S�*<��ȓ3Z�]Z���-]JZ����T��Ʉ���1;�d	f���Т���'p�Dy��[� ��5�J |t:���'�1�!�d���.�˵�M1k��8�Ķ"�1O��Γ�p<�p)%e��8!ă�y�̹I#.�q؞�&�pBL?! �0�M 0&ϔH� ��y2�SD�Yb	+v�C�#� ư<Ɏ�� pbJ\�F(�S��zD�x!�װ1� v@ѹ:d�e
�BZ�"�p�<��D�� D�1�bE]	5���H҇�U�<Y¬ʤul�mĎ:w<a���e�<��\?�R]����oa�|�Go{�<)�B�P��	�<�$X�� r�<�	�=~�X�ʂ,��k�BlAa�IH�<QdV7h4aS`�1���@l�k�<� ,h7���?�XH��^��B��'�x�"7���\z<���(~�ˆk�0r�����R?�wK#,�$ �H��Yu��z�<�����$:Tk��t	�Q*�H�p���2�{���}�R�36B�&^��T ��ybk֙:~pA�iX�)��á���y��ʛF����j��Y/�l���ݯ�yR�F�AX�[��P�R�2�&��y�A]D
����S|���ptH��y��ɍ#�\5ȎJ�����H�y�ǞqК8��
-3H��3(D��y2Ù�E��E�5 �9O��)D�T��yG�nBlPr��3\N˳MA)�p?A�OL�����4|*��2/^�r�:!�q"O�ȹe��=(� Dct��2�2�4"O|� 5���
%X��	,=H��"�"O�t3��=�09� #˸7B��Y6"Oa2�C�0���Pp"U/�6H�W"O>�(��Ň6���#� 
�+{�i7"O"��� ��|w����5���sEOf�d�(�R�!$.ԓ{�t���*r�!�ټcnm�w��v3��X��I ����'lH�}r���7��(`B�Uxy�p1 ��j�<��a�avj��)�&e2	��%���+�S�O5���7��'�|
��ں0��;�'�@��"���Tb��"��Ѫ&�h�s��D=O�K�Gϣf���c��K,��ɪ�O���J��@t�j�NR��UH�
�!�d�?䔴�SJ]=n��9J��� J�!��T�!�4ѣ^����bu�c�!�䐍0q��ʕ,7�8�1�_s`!�M�*)I�2k�#N�<XS�O�G!�Dģ �p�A�N�������̣=!�d���)���-fzIL3*5!�d�qy��2"/�"O]B}�^�w!�Č�!^ HQ	�f23�˪!�D�(I� h��H��!��[4!��7�Vqċ:��I���Β`�!�d#u����"�$�0����B +!�A�cK�$��G�v�.$�&�ƲV�!���{֔��g�7#�F1�2��tv!�U�/ �q�㠟[���*�Ȕ�}i!�D�Af�5���N�e"��T�śY!�$֚d�X�aP��n0�!p�S!�$��m�t!(j-.�9e%�q�!��<	U:(RW�N�~��1`�#Y%!��t�yF%�/֊i2���!��[--j� )�C,TlЌ�F!򄆝M�P�s�OѸ?�x���" !�O�m XXAkN��Rµ�� U	!��Ԋ����;��D�#���!�ě* ���&�F�E�,�@���50k!��B�e2�k����_��ÅC��S!�$� v�]����%ܦ���̈́�!�$M�W� �Ief����!ՌQ�!��FK���eƴgR}��*���!�]$ �f�
��	���Q	�7!���H��|����+a�`
WE7B)!�D��? �pصf�.tVԺV��!
!��8�����5k.*`R��͘;�!�	鰜	w�� 3o�t"�η,!���S�ٻ�@3o@��	@�J r"!�Dި�U��^ WG���4�� C�!���35����˛+M)s�'��a�!�� ����8;,R4o3k�h�s"OΝHw�W�~�P�օ*~���W"OH8�D	�  ^�����[[�d"O�Pp��qԤ�9��D�4-$���"O���!�ɖw+�D0FHR�l@��k�'!��'��'2�'2�'vr�'>" ������K�P�i�'�'���'�R�'%B�'���'Z��'�>�� ��7��ű!��m�@��a�'�b�'���'I�'�2�'�B�'����y�Y)&�Ҁ3��I��'��'���'^�'^�'���'
�(���w�\@��5�|Ա��'l��'���'yr�'�B�'�"�'G`���U6!U�!<7�nܳU�'sB�'�R�'���'�'�r�'jč��	�DǮ�h�i�2����0�'���'���'�r�'���'���'�P��Ⓖ:�X}B�KH�>޸Cu�',�'��'���'���'���'}h�v:u9�n	'c������'���' ��'xB�'���'�R�'���R��,À�"�Ȭ>n���#�':��'	��'��'�B�'d��'4�����ӊ _��S�.3zKf��W�'�"�'���'�R�'i��'A��'� �:` W��J�YA΃cQNh��'r�'�B�'\��'�"�'[�'�A jV�r��QХE�c"���'���'&r�'���'�"�e�����O>h�!�1C�Դ��$�~)ƥb��fy��'��)�3?�i�^�����5�|U�p*�u=�T���N�����ަ��?��<a�O�$Ͱ���-�Ti��׶T<�|����?�J��Ms�O��;��M?���� +j-Y��M�ܰE8T�6��՟@�'��>�
��҆�b(�_?�P�W�/�M�r�l���O(`7=�*|�II*@D��g�P�c'z����O��f�֧�O���ӿi���V��!��<e��	EܐD�����P£=ͧ�?A��Uq���J&�Q��E�#��</OD�O�5nZ"U��b�4�A��NT$hL�C��(c��F��	şT�	�<I�O�x�d�!j��PGD:8��������	x�ؓ�<擉x����leL�@ʹ�� �M��<��n�fy2W�8�)��<)��Ge0 {�I�L%�Y�ON�<�ķiO��k�Oکle��|�J$&S����/�"�0�6�H�<a��?Y��Ϩ�۴���|>�0����U��	�<N%4Th�����c�;�$�<ͧ�?9��?���?���E	"	�Pe�%���dL ��� Ӧ)#S��gyb�'�tӢ�ͰSU*�=eQh��(�Cyr�'�&3O�N���O�L��H, ����B��(�8U�T��B���p���H5� y�Nyr�
�^OƠ�� ���}[֫�b�'#��'��O��,�M�"����j D�&�(mJ�m�&~4��j� �ش��'Țʓ�?�۴V.�&��
m���őO�pt�@c�������i��I�x �d�O��%'?��\c�9��"웥�� p��0��'��'VR�'>"�'/�d��W�<]� ���*����D��d����MK�,}�iz���O���s-ҟ��c�����m!f�ݟ��'� 6ME֦��b�\mS~b�/k��2�(� �|B��N�S��P{�L@韄��|�\���	̟(����T�䔴%ɾ�s��,"�E	́�����Ty�c�䙚`��O����O��'o�nQ�-i��� W�t���'Z ���#u�4H'��'{��
�@k(ܨs��rsR���/U�1,X0�F���4����
B�OT���&��! =*%#""RAV�O��D�O�����e;5�?����?��Ywr|Y���ӸLz���У;8��eJ��	����?!fX���۴U
|��pϽYoZ-S�� l6��i\�6M��5�n7m`���I*��R��O�섔'c��k����+g��E��d�iP�']�I��d��ߟL��ޟ,��B�T%�����vI� m\�H�͒�fO`7���"�*���O��*�9O�ozޡ;�C�:%Θ�ĩ�%�h#3��MSr�i�$7��J}��%��&6O�P$֩-WHMc�j]q�`�3�0Ot��G��7�?�
.�$�<����?Y���K�T���!�<�l�S��?�?���?�����D��ٺ�'p����ߟp�u���>z��)�-�/���se�E�y#��'�M�"�i,�'��a�b��:-���"���y�hӚ'��
/�����F�m���?J�xӴ�`�tm���Ć/�@QAB�ƒ������?����?����h���ĕ30�Lq��4~= I֕J F�d�Ҧu�Ĥ&?1��i]|�w����^O��0֩��9o,���'H�7�����	�&�޼oZ�<y��B�p�9"�ú+�EVdT��$BBӐ����%R�O���?����?���?��>�ޕ��S*�A����O��8z*O�TlڍvyD�9+�ҟ4���?���_y陕1 �\���'e�Y祐�1���4��VOaӢn�n�O���b`��/qW�T"�JR=V�,S疳-l��dQ��b�&�]���U�IWy����2��a�S�B��C�W�(*��'���'��O��I�?�	�ğ��Ӈ��9B�dZwe�����"v��ȟ���4���?Q2W��Pش	���n��uI��?fb�m
�͖fY-��f>7�b�L�I�e%<P���O��H�'����k�� i9�%ӫm�J �2[�p�={�:O0���O����O8�$�Od�?�;6',S����CNlt��c�����Iꟈ	�4#L���/OZ�l�X�I	Q�¨��)�dj���5�U.U�P�̓���I�A{ݴ�?y%	�MÝ'��B0	�L�r��g�zE^F����NƟ�{�|�S���x�Iܟ�4'ԔD$��b�2e�
�pd�]��d�	Wyr�rӢ}�j�O����OTʧy��!��lZ
.��xc� rȪ��'���R͛6�w�>��_��?�
�l%P���;�.�#>X���c��t0�ŘC�8���!j�O�qpL>�1�$���+�`rQhA�[��?����?i��fFXy��[���'5��By�sa��&>�usum����x��哙t��Qo���dEO}bl}�2�I��?(��kؽSF����"�ݦ���4Ô�cܴ��d�?eL�b�'BF��uQ�i��O߭2���
���*�&E����O����O��d�O��d�|���J�~o��ȟx�4#߉bg�U~?���?��'��9Oҁoz�����m@.��G��WڤTa�b��M���i���ĵ>ͧ���M��(�4�y�m]6,� �sIIFJ������y��
9�����O��'��I䟈�� 䚠â� A�a��ܖ�vt�	��T�Iޟ8�'΂6��~��'�*?׊p�bΛ+����-\�Z�O���'W�6MUܦ�2���dK�����-L�`��Cd�92��	ZXTy���>sG��%?���'d�i�	"v�1�"��E�I+�N�1������	���g�O�B��/����H���R�&_^��n�4�SO�0)�4���y���$?z��!f\�M�jd��D��y�mj��oZ2�MӷI���M[�'���F/y���S,?~4iz2"�#F�" z5$�*�������O0�$�Op�d�O����H��Չ��2�L�۶�J:8`��O�؇�P��~b�'�r�f��s�� �@�x7FT�@%!�ܱQ��+���ZǦY3�4>5r����O@��("h A�R�X;9�(��"�H%*�b����ɏ#Uh���'P�&�`�'944��i	�Sj���"��<R��'��'mb���]�܁�4G�2u���(�J�#3bӂ$TuA�������pq���H}��c�ƬoZ��M+�O&K�X���њv"h����?S4�޴�y"�'���gJ��?q�@Y�����ߡR��6f^��TЎUV�Pi#G|�d�I͟D�	ğ�I�l�2a�ۏb���R4�f���8�?9���?���i��e
gR�Lk�4��>X>c��͂"��@�5��/�25˳�x��bӀqoZ�?�7nĦ���?���0�$uc��NV���񕌟�Ć��Q��O�taO>�)O��D�O\���O���2�ګxz�؂��;a�	ccj�O&���<���iSb�Y����r���I� qZc�Q9�F���hW����w}��w���m����|
�'Z21�l�m�&I�Q���s~��$#Et�J�a�щ�yRA��O2I�O�O&��I�֘�e -h5ǈ
o4��KH�m��l��ȟ,�Iӟ��)��YyB�|Ӭ}�Y�Q��%��OQ�H$���Ɩ1Ϝ�����Pq}b�x��qæ��1�ܕp�-��}���������)B۴%t&p��4�y"�'��(��D�?���S��ٗ,G$ 2R=��'	�r%�d�i�L�'%��'[r�''�'��P\`&.��il`����5S�`��4_�v��,O��*���MϻNn��藁�*��0;�O�If�Ӷi46
j�i>��?�cc�����o��i��d��
GcR�/��	͓���y��O��H>Q/O<�$�O(�.I>6�!4D'A�
�Ȥ��O��OJ�ģ<� �i`B�rR�|���N]q�L m8���j�Ƞ""�I�����ɦ��4N���>��ʮ{�$j��'��-@���<��@~�XU�ӞR<�)O�iP��?����O ��r�Y���A�ޠPr��T�O��d�O��D�Ol��`���h�O�.�8JP�j���0(���H%]NR���U������0�M����4��.'� ��ǆC=!��PWoӷG"�ڦ�ߴ69�VB�f�������-i��e,}ܐ��#9;8Y�\�pjd�$��'%��'���'h��'ej��4�O�b;F���܇n�|4k�S����4IT�p��?�����<IB��]�5��'�OG �0��ژ`v�ɶ�M��i�ɧ�O=��z�B��Ht4���o�=�s�+ˊLq��"G_�$0Ъ��.' 7M�����ʞ?���ձ`�,��wۖk�,���O ���O��4�Z˓g��FI�5dWb	ɳj��D�+G�M�-p�^�y�b�p��"�O�$o��M��F��S �[��e���Б �E8�N%�M�Or�X �W9�����(|���E	�]U8"��ދ<��	�`�d�����ʟ �Iǟ���MLY�1x��
6k,�5���?i���?YV�i�$d�4Z�R�4��)�����iO�~���pO�R����'�����M3c�ia��Hz���=O��d��]u�����1|��1Ej�>4h ]C�fZ�?Q��?�D�<ͧ�?a��?�B�p�	�c��1�.��GK#�?!����\릩[7͊�p��۟��OR$��J���`��>c�"u��O��'�*7-L˦�Γ��'�r�˛�2���'�|�ҁ�O�Z�$����ž.�8��'��$�ɟК�|�N6a�h2�&J�ł�1�A��s���''��'H���X��[�4 ��qKu���J�y�ٹ�ްÕ�P���d���Y�?U��i�4A�ZH@���3A�l�Cb�3+�*	��i�|7-Qg^6mw��7B)_���v�OŜ]��?� ��KFF����Yf�2İ�*Ĳi��'��'y��'�b�'��ӎ`{2�t�MvxQ�'bب[p��޴ [l�Y4�ݐ�?�������D���]�'l�8����9e�PX�P�w�,eZ�4g���yӮק�4�O����:PP�6>O��K�қ%�LK�K֨��� �1O6�Ad�ȷ�?��6��<����?�2���*����8��ѯ¾�?����?!�n����ꦭ�A&��?��ݟp���J��
���f����Ri�ƟԔ'�2D�<����M��iB�\��'�4�&�� �R����	��8A�:��a
AWyR�OIJ��	.��B./��L��N��
�=a6S*y���'��'�R��^�����	�N)����צ��S�>Y�iq�O��-��m��h�6h7�!�'A�2�Ʀ��޴@˛���z�v;O���ٲ@$���<�:�ۘT��j��
t+ħ-���<a��?A���?���?��K�1[tp�E�	��l@*�E����U����O&���On����F�(t��5m�T�eÌX�@��'6�7��A����H�Z��n��@�F���i� &��q6fA�x�I�M�<	ǁ�J�$P7�䓜�$��*l�pK%��:ǾqI�X`m���OV���O��4�DʓFE�vdQ,6#�B0���hG�1\�> ���0�y�@e���«O@il6�M;�ia���&X-$�(�e�Ԃ:?����'g���3O���̿.7�ܱ��UH*��*��ƈ8KCY�	?�M27�N2U�-sd3O���O��$�O����O��?m1�(+�2x��iˬ[�>͹�BX�L�����ӟ�rݴy������?�A�i��'�$�����8 X�)0�	U*Lg���ub�T��'�Z7�Cצ���"P�o��<9��y��������:��#CR�Z%�ݮyf2��ߪ������O����Oj�D�o�\��`�?;U��p�O'��?I����Y��M�ڟ���ԟЕO��p8���"2��(�)�#Lf�pb�O���'��6� ۦ����'�.=4u�VDJ!)$xWKf�V s�mS#H��<�<?A�']�2�$�9��4�Jx�(�(@;��B�S�B�x��?��?i�S�'��D���Š����7��p$��$\�����P�{](Q�'
�7m>�� ��$����2�] 4t�ਁ@�u-.0�n��M��k��M�'+R����8h�;D�	|L�ڶ�"`�Ĕ!VQ�~���ayB�'��'��''Y>A�E��f\���w����§�r*�io�.]���	�����t�s��	���K�h�,=�.�K3$Ԣ���Q!��t����p���	f}�O?���'�Z%�p�i=󤛏�jU�p��:��m�A)�;xa�W�k6"����
� �O(��|:��HA��,N�2��ȉH`D����?��>�ta-O4mZ�F2y��韄�	T��S��)���y�č( �f�%���	������=��45-�^>�R0"�%�
C�L�)���h�w��	=�ˊC�i�BYzy��Oj\�Ie��.¡`sr�� M0X�N�H�Ϙ/X���'gR�'��S����HO!�`�A�U�7�<\�����	�4*�d��'g�6m/�i�a(�G�3?؊�K !��j�vЂ%~�<��4.���'#&\�w�i��d�O�T���-g��.��+*���Ь��sKȹY/^�'*N>Q.O����O����O��D�O,�qD�F��ݠ��̱~6�t��<��i�����'��'���yBG�7Z���k�_�=#�t��9K�`�g��6j�Z��L��?����F�RuP�eϤ9� X0��lM��00*�%t�2�i�  �O�8�L>�(O���J�}EMYBВ���]0��'�B�'j�O�7�M����?iw��:+���d��ҩU6^R�xy�f��J}BpӘhm���kB�ħO���U.����0�"]>pS�oZ�<��3�ơ����H�'n�D�i���R���Rx�����z���Iߟ��	ٟ���۟���I����(B�\��&!+7F\0�?���?�q�i�D��U�4�ٴ��\���Y�bFqh�;R�[/i]�P�'*��1�M[��i�R X����9O��V&[g@�0��F�0p��ߝ�Ee,�`��2�O$��|���?Q�`{��s�	��*m����,~R]���?!(O�l�e��I�����~�dfQ�+�\����2܈@�TL	���}}R�x�L5nZq�)b��5Gάu�7���s���7��;\�k��>c��:+O��
�O���m�y�ɇ">���j�:QnX6#V�������	럄�)�eyR b�*��GOV�8T2��e�l�"s�̽��	��M����>)@�i\uAֺI4D��f�H ~e�q�P�n|}P9l�<��Ӣ�B��S8��.RHy��,8ؐu��
<p0���B�dЄx�0�[�8��G��D� GΎ:��ձqu� G�T	+��Sc���6J��Í�kM��!c�߆U�Z9`B]K*��X%
8C�����^,0&�� )�ѩ�E*��&l�x@��-��y��	���!Z�1[f��M�p�x� `J��(�S$�'���a
����G��c�I�mR. ����Qe�(m�!�r'�{���I\:y�=����3K��QfoW$4��C�f�&q7����%�b�1A&ND��z`��X0XpYUG]�;�V�'B�'{��H<�$�O4�ٱ�P�� ��D�����BE���-��ßh���� �	�?$?����P�8|k�J�.0���� ��|W:Y�ߴ�?����?�Ab'������'=�D�	&PZ��w��7	�UC�����}yB�B���'D��'�
�A�v�(`�\�Ԝ)߭_K�7m�OܕᆋGZ�i>���ϟ��'�v�E[�P�P��)VR$5��|Ӧ�$˳>R1O��$�O��d�<Iw� �i�w␇C�t����<B�&�г�ц
$�'���'�'��1RSL5��]�v�RP	I+@&�yŧ0�៰����h�'�x�$�u>af�Y�y���6Y��8E�>���?�J>�+O\$zu^����M��A��Ypah��8 b�>����?�����
��'>i���T�����8]L���a��M���?�+O
��O\����Y;��
�m5gd��B�ր_���'��\�����'�?������Y�Pȣa��B��43`�M}��'��	�sf|#|��O����EO,7B�!!�b��W�P��ش��D[�2:��n���	�OD�I�k~�\SD�N5���T��M*O������禕(Ѥ�qE8X

� ^�$q���qӾ�'.�Ǧ}��������?��H<�'3�@��6�W%���#Gd�s|:ybV�i�v	R���I�\�3��������X� -Ӧ ��
)�e喊�M���?��yk4��x�O��'sb]�fI�:��QkG�F�%�e��>����?ypcTu��?���?�����)���R�dʩ>Vx�xW�I�4���'�&}0U�*�4�$��2�D
;ņ�1-�=?7y�d@����'6xъy��'��'�ɾTxdM��F��,@PWM�'3��Cc�>���?1���?�*O:���O���ʛ*/P*-ptB�3��z�A�:�1O����O���<Q�gT��ōkfD�g, .n\����_�a����t�����'���'���iX�m���C!$�cXHc�S��I����	vy��'"����R>���4H`��j�z}��2Mݵ-�69��4�?q�2�'�:�%ۋ��v
BI0�혤]�*���#�;eԾ,oZ�L�'�gJ���ǟ8�	�?Œ�hT�XRe q�C�^>Y���!��'��H%`2����y��r�Q��=RNe��Ž��QeT�$�	�E}�Y�	�I�����AyZw�����Ո4�.�	R��"AT��OD�$T�=����U��)�� ,p6oO�<����ޙ}Ǜ�kؔ.�2�'���'��X�����a��L<AY e2@��0U�؁�Qi���MCoL/3�VM�<E��'�k���y�u��F�J���'�v����O���S����|r���?�'�Nx�`Y�<��@�G�@'p��ZB;�	���M|���?��'T�hC��T
N@$����$l}��4�?ijC����O����O�H/�dS�3��e�nB��>aq�ւJi6��'���'��Ɵ��ϰ&��9ց�^ �+�솜z��H�'z��'"�D�OJ�Y�zd*u�)��a����(�<��Z�����ڟp�'0B�S2G(�	ؔRu>���͸7��a��� b���'5��'�O���w��u���iMT\�t��8w�بDN�'e��-K�O����O|��?�rI����I�O<H�@(��=� ����:Ax�צ��IS���?Q�� ���%�pQe��e�@H��;_�	�gj����<)�,���*�P���O`��Ȇ6��2�¢PZ�A7iM�
Fu�>Q�&'�=���o�S�T�[njI�w)@(���#�����d�Ol �6��O���O,��럨�ӺC�%�W��`��M4�x�A�MKw}��'az�5l�����Oc��j4j��b�����#�'5S,iX�4M���?���?��'��4�6�dR�?��`��	w�xu@ɔi9�o�!u0��V1�)§�?q�S;
�Ҡ�ף��e�ڬ"�ѕz�F�'���'��h�B^���4�	}?�䏆Z0$Ѐ�	�-��11O�
��	}�֟���_?�W?f�u:�Q�>0�ǭ����ɫЙ�'��'�b��۠T�p�e��K����ZSԉ'h �!�O���O�ʓ�?	5B�6U��c��Qu��Wm�	|&�i�(O����O2�� �	f?9V�זk�p4��˖���Z�j�٦	!�B%?Q��?�+O���F������ �а!+L�� ��&��6��O`�d�O��(�'+8u�ݴG�\M�v�= ��Y�jL�f�T��'���'W��� ��" v�4�O�9��5 B�Ó� �e�ſi�����O\�`�肰0	�'�4еBsBPr�N)s��]��4�?)(OJ�dM$@�'�?���ꠋ�=4���S�*"> yN�L�O���S�_9
-�#�T?}�2cН��esn�<ex��0j�>���c�������?����?y�������D�S>|�@ĂA��j�h��_���I�pz��A�<�)��*
!�����@����EIJ�v��7�@02`��D�O:��O��	�<�'�?y�W�+o�����X`TF�b�6m��Xm�|��y��I�O޼�!k�e���FASE�ZŹF������I�H�Ib��������'��O�)A�Z8mQ��q�g8t&��%�Qn̓g��msҟ��'�B�Ob�R��κ���3�\X��iHbl9���̟,�����=�6/� *����RY�I�%��i}B�Hߦh1�O���O�˓�?I�
ɃZ<"e�ȸ{���k�O6;�:8 -O��D�O.��6��ş��!״!\uJs���v��qq6��U?�P�-*?���?q+OV���[�R��:�\3@ �((�`�Ag"٧Fwl6-�O���Ol�p��$@Qv!JFa|�Rph�!��qފ�{��1�de�SR�4������'L�e�p��Sݟ�� ����\�pY�ăV6�:�;u�i����O�T�%m̰%&�'��H�P�\�` ��j�ۻuMV�:�4�?9(O��ӷgu�˧�����A��i�LH z���R&H30��S��?QqE�92����<�O�|P� �&?�. %$ɴ8 \\a�O4���H8�$�O,�d�O���<�;HLpq�ŌU�;m�J
��>.��'���f_BQ�y������5ZE�M�.+V�j��َ�Mk�=�?���?����J.O�I�O� P��_�.�
�s�N��	C�!��e�����W-�>q"b�"|��R-� ��G�O=FX�$�*��:��i|b�'�£ҁ]6�i>A�Iן���M��yu�ΏD,�94!�O��#��${*h$>��	� ��t���rN���)���֛��l�HkWD�gyR�'�2�'�qO��4��-\> ��IJm*I��_�`���2'�$��?�����$�OLX8�Fv�h�#1�ߔSU�Q�%n�)mf˓�?Q��?�2�'JJ�Q�Cпi6$�ăE�I��U� �G�.�� `�O��D�O˓�?��@����]'X�\4Z�(Y����F'���M���?�����'}�.�	+(H��48��J�@Ӏ&N$+�H��i��'�2�'�I��Hڄ�	B���'N��@#�'�  ���P��|ٲ�tӪ��3�	՟`��L��(��O�d���2G�a!�0pR� �i�RS�\�I��	�Om�'Y�4�t����R��v��*э�xlc�p��
5j�M0�5�~rT�X(t^��Sq�y�4��_}��'��̓C�'l�\�|�S}yZwX�����ĩY�$L��Ϫ@��͕'��-�7T�`q�y��!�3g���3%ͻ&��8��ɇ�M˲��?����$�V��|��p��1���7�&���E66�T���i��9	�;����j��	�-�8��1��	�T@����-��oҟ8�I˟X�a�ry�O+r�'����=�4�s�Ept-X2�
k.��<����щO�2�'p��+!oZ����E�Ic�Y�酏�v�''Ԍ!&X�@��П��d�5:���֢Mҵ
����\;ޠ�'�L`aA������O`���O�ʓb���A7�\�O�Y4D
	@�|1����P�	`y��'�I�����H�t��
ºL#)R�6~���B_���	��@�	ԟ��ԟD�'A��Ыw>��C�Y�F�R�`Ũ�p�R�y�X��?�.OZ���O��Ę�o�ĳT�L�X�^xY`%�K
a�� o�4yw.���4��Sy�J�+PT*�'�?)�#�CJ���.B�I"��F��'��Iɟ�Iԟ��q���I����	V�<}K7f��T��Ӵf�g�T�	�,�'�$�q��~���?���h+�5��	O�d+����Q(9����R� ��ş��	�|�L��r��'\�If�z��u��.��x��װ��\�4'f �Ms���?����b�V��2 ��]B���%d9C��y��7M�Ov����y��v��'q��#���Ȑ8��mS���p�i5����sӈ�D�O0���l�'��	h�2�L�u.2�S���76|�(�4u�U��?)�o�U8����O�̕ih�8��t[��1��$��z�D�$�O��dו�.M�'������j���b��O�g�0��q��X�P)o����'=�m��)�O�D�O���j�x��|�q�L�N�P���I��z=�tҩOhʓ�?q,Oj��ƪ��"��FS4�dW8K�>��Y��*��f�H�'k��'�2Y���%� #H�P8U�,|���N�Й�Op��?9+Or���O���<#���s���=8�n@�&&���z��5>O0��?y��?�,O�u�Я��|z��H5
�${��ݐ@l�
qkz�ʓ�?�(O����O�dNd��I���ْ6��4��a�bɐC�� o�������<��_yR-Zg6ꧺ?��T?��R�L[�p��yQB���s$�An�Ο$�'�R�':�k���Y��S�0F��{dˊ�f��b�n��d�Onʓ_ЍiAR?��I៼�S��� 32��J,TQ ߃Sbf��O����O���y7�Ĩ|���D�X3]�|���J��@�*�"Y	�Mc.O�q�J�ᦵ�	��	�?�+�O��#,�9@
څA�$�x�LD�W��f�'B�Ì�yr��~��:��OR~�{5���fe ��ӎƳ`�.E۴t�*���i"r�'��O�����+,(Y�5぀*�xq�/8]�mZ�z:��ܟP�'������N3<ă���d���&@�>Zذl�ϟ0�	��(SBc����<Y���~�Ӻp�2��tj�?�r%��Η��M���?� �a;*��S�T�O�R�'��!�%�� >�p� G~thJCa`Ӧ��-��'��şd�'Zc��z�D�e�������=y�0�O�}Bt=O�D�O�$�O��İ<�D
B�ք�����Ҙ;��ȓ3�,P9V]��'B]�������\��p�-J^(pS����	zT�s����������\��ly�	�uj�8'r<�pP5[� ���C4}��R�X�IJy��'�r�'�h�'%r�@�FG+s<nY�E��B��iH�&a�����TE ���O�ʓuKB�e���FG�i_��٦��,�B-�sc	%6��Ot�O4���O��B��Oh�'�x}RdlǱe�����Iޣt
��yܴ�?����$�l��$&>9�I�?=R�"A����r�j�:5�!k���D�OB���OB��P�Oh�O��S�r�)nB�I��P ��W-T��6��<A�C� ����~*������� �D+�e��-�R��f�@�d��@{��i���'�J���'(�'�q����M~9B͛��l裇�ioR�A�BgӠ�D�O���䟦�$����UK�n̎��qH'��>�B��4���������O)i��2����Q.^V��N�V�p6��O@���Ol�����N쓫?��'D@<��刭?v�+��$ `����4��Bi*�#u����'�r�'��Aj�~>�y��d�,'���@��p����N6th�'����ş�&���%Sx�%	�卥�ܥ ���W$��{a�M�������O����O(�t��pFEx� �x��B�*5mQ�D	W�O��<q��?Q�'�Y���ů�nq�A�ѐ5Ú��&d��?q(O��d�O���<ه��A�	,v#H�g��2[�����k�\�I��\��H�	��X������ɻ�t�)7�DHV�[5�ޡ+��#�O�$�O~��<�����Oc�	�A��v��PC"I%WAf���$z�*��1���O(�$@.-eD�d(}��!����wIȘΔu�AfO�Ms���?+O�:�P������!�2ihR$��*�>�b�$V�G��9N<q��?Y���?YN>��Or�	�	ϸ|�ԵA 
��3����4��dߘDi,�m�����O���Y~"�_�02識��Zy:�8[����M#��?d�Q�<�K>�~�L�.�J&д@X�B$�G��:u�V/�M����?����*r�x��'`*� �D�?X�\�`ǂ<�z���!r���FB�O�O��?��IA��c7-E�3�\���Zݸ\��4�?��?q�Z�?{�����>��NK-�bQ��o-��5�SЦ}���|���?�f�
J|B���?Q��d�(�4�� ?���!�bRgvRX���i��N��XI<ͧ�(O q:�-�3-)�mh�
w����U�x��d�̟`�'�b�'�]��w��6<��� �I�W!ް`�iǘ�H��K<i��hOF�d.O��a��m�%!��Mbv-�=�2�X���O˓�?I���?,O"u��.N�|��M��-���Zr�Q�y�0��¯�@}��'�ў<��g�p5�	1Rn�1ҨJ�M��`���>g�0��O����O����O��$	�rc4�'�~�ʜ�q~t$�f�^�,�� Bi��M{�����?q��p/�|g*�e�	�Z�Q��&7���cA�8W�6��O2�Ħ<ie�	�/��Sȟh�I�?]
A��fҀ��da�J4�d�HH��M{�r��������i�l�� n߼r�F���:�
D�޴�?��o:�};��?�+O<���<��Z�v����82dMy��R� 6!o����>Ye,���;�)��#c����G@ΰj��lj Ŏ9��7-Y�h�4�$�O�ʓ�B��?�*O��i�`T�!�4˖�C�[��2����N�'&�c�"|
�_e���7k.�ڬj�aH�M$��v�i���'a2�H<V듮�i�O~��֬j`0���WUҸ�C��1���>IVM����?���?ɰ+V�P��I�8ʶ��G��0mś�'^$��0V�x+��~�d.�d�g�f�2%Ƽ��-3�Хkx���'B��S��'��D�O����O
�D�O&���D;��U/�)R?�(�b�ұH��˓�?���?qO>����yAQ?
��]�g�
 ��I� '���2Zggz~��' �'��	�=�D˝O�MÑ��_�dcæO�5[�$�ٴ�?y���?���'�!�O�M�A`M�nޒE�敔"c��eS�P����8�I���I�N����	џ���`l����]�G�8X��אKB)mZ��'���	�42��޸T�NO�(:�X���#�\8���ׁ�=?v@��f�d,�g?9��W�W? D �J��� �T�<s�P=r�%Z@��gk���0��W �  ��D	��\�b�P���ӻ�]�@�K�vO�u�׍$�Rm��!E�֤���7_ͪXI�*�K����B̠�R*��b��}d�;q���!s�8�'(�_�@`s�[���=q���^��(䱝s�^���T����'DZ����gH�9�?i��?!��p�nM�_���a�[~�Ѝ�a�|,
,�l&!�f��*'jT���@-��<��	!��	:�'�`�H)s�D�fzj����ָ4259��X��f��F��86�>ţ+��x��E��y��Y>�����P�VC�P���2&��O�	'ړ0C��R�Q�C�0��K�|^�ф�W�f����ޚuf����b �1���'2#=�Oz�	�`��b)rxTX@A���h��[)"k �Iɟ�����^wyR�'���QV�jxSOL�LO������}g� `vI,����"Ǩ	v��"� �B&D(|�~�'���Q x���U�
8�K^�Nc
t �	x���#O��f�� 9ڭ`�Y����	G�'�O,i�&�G� �4 T���1"O�i R�I�8FX��/��8�6�ʋ{b��>�/O"�Nk}b�'�>u  ��=yp1���j��Y�"�'���׾^���'��D��U���N�4��Ӛ�頫^9e��KR43
Ȁ��'�J���D�G"��3�S���.ͩ(d<9�H u3,� vB�p<�`�L��IEy"���%+�u����
0THb#����'	�{��ʿ+�n�h� �G�$��Ȁ�xbu���I1Ë�F4\�2hO/�9a�3O��|����i���'"�Ӻ_�|��)� �ĺ�.#Ӛ!0w�Q�:��3�H�O����C������ c�n@������'�򉖂Fu����TH��X'i^)&���"���l�"`L"E[�èB�J;1�"-���'h��z���%0(���#g� �OT���' �7͇Ʀ��	\�'����$Y�{-����I��t�<����<�V���dER\3Lڒ!�ZW��B��Ѝ�,ĩ@F�V�i3 x�sI�(*"�n������֟�j�d�8G�������	�h��6����b	9eY�k���"��!J>���4�|&�T��R'l�D�H\��J9�5�@��-����6�(�3��ԙo�̘("�Y	��\)��^�!1���O��d�b�j��Y�����9��*���U��}*䦓�+z���b�B�!e�F�?�Bi{sM�~FI�'�@"=q+��
u�H�aܡ`����q����ͫ��Z�H�4b���?���?	�����O��S/Z?�@�� _!�iQG(��a��#�;����tӎL��z�B�@`��a��Z�e�񅚻(2��sǀA�Qp`�ֆV\��,xP�E!oh��;tM�JJ%W-��Z�$E��A�ܴ��'2c?�P"�0��/��9݆�7D�8k'��?���+b(C" ƶEP�	5����<ɴ�?�����4y�ߘd_N��v�_�N��g�ޟ��ɓ?n���ßh�'M<��� �ۻ}5&��4��Md�w;f� C��"�jY@�Kf8�����[�Th��鍸���kg��7\���A� iP�����pߤC�B$�Q4h��	󟐕'͡&�2"�	�q���D��y�'��yb@�*�ȅpE��=���#Y��x���"��!/Ks�<I�#�ߵI����w5O
b��֧���ӌX�� ��ܫ[Ѕ�+��S:!�d���>��Ae�-N�Ђ'�o4!�[�W"�� r�E���4�!򤔴k�Bdᗇ��-ȩ��,p�!��K3{2�Q�D[�M��칔�ˁG�!�$ݪi�1ˇ��>�ލ�p��EV!��ŌuU�a���;�f%1��^mj!�䒼 nv\��A�4yh�)�(^!�˥e>T�J6k؀&=%9ШIeZ!�dT��H�a .Dp�GJ�:D!�d� 
�, cҋ�f1l�co�l�!򤄳"V}򫆛O���C�Հ*!��U��2ɱ��ϩ�zlQA�Q  ?!�d��d1���$u�ݱQd	�j�!�_"�(��BV��2��Wcҿ.}!��*Wʒ�s3'I�ϰu`Uiּ(�!�L/�R�ѱX�x� �(��K�!���&P�ЗgJ&|�p*�'ԩoj!�dѪ[.����I�'���f��H!��<��*���G�B��#��/9!�d�v�L�(1���l[C/��6�!�MU��`@2�J�Kb8}0�듏I�!��@h������;
h���0kЄN!�߲"4L�H%��@d�M�Cڒ"P!�@!h�d�iFB_"m\�!W	��S!��M�5FN@�P!VF-�T�0�!��3^t��Dý1#<է�*�!��6?l!�a@Q2.�V��̏N�!�d͈_�����0��k~}!�G./������L.E��d�D��1[�!�	6���TlX��zΛ6P�!��&S�Xuѳ�~���)4��n!��ܒhKS`�2V�-0q��1;W!�d�8H��S�a2A�ω+�!�$I�2)0{é\(���ғV��|2L�
�Z`H��T:~�Zyꑆ/zgpx�	żM��ࡥ�G<!ĩ���&x[�)�����S��F�'����F�C%q��L�K(+��O���1i.a4\�"Щ6`ȑ�'�4�٣ʑ���mx�G>4�F8��E��]j8+Eög���@�񧈟�>B���(�4�,�H���!��GK����VF܆�����׿7R���@9�TLK�-RJ���x%�'�S�? ,�db�:�XѴ,�p�py��'y�A��9�u1W��3XjxB�ǐ�4�I(1�Ƚd5��:��O��i�MC�mM��Q�+�h�P[�"� a�B%��@�<�x��I=A:�s0\�a�I�)a������gb�q
J%s���2�V,��뎎y.��8�P��6��x�bο�����87J�p�'ʨ�f��ף��|� �p��'!����i�bԠ�FQOe�(s!IpU yZ��_bU���5���dò"��E�4�V_�M��N�@6��F,��1"si�4\+��
b?��e�=Bl>-�k�PI��		b��QEg]�j���o�^�&��dԼC��A2�D~�jCCۚv�z'IB�6��叜V����9M��0z6���(w����Ӫ*:�M� I��(6�9鑎���"<A֌�5������a��}pN~:Zr ����7g��Պ���Q;�=�=.��C�������xBa�Xƺ`9�C�d�*� T�P9(ԖA�c��31�EJС�> UBa�F�a;�S���9�\�Q��]�M*�R��ޡ~p���"Oh`����>`�B�����0��O*���N;$h���dG13A󩂪^��A����h�v�
���y�"���b�r��׮S����?{�<!'�Z[�<��{���'H!��K������O�p����>4����;��*��40��Vx;���Xx4 ��)>v:��զ�����	@����W�Ӌ��pH͍BĘZt�Z�9e>���əfbB��	q�t<����= ���R"��z`��;�j�9�D\c�\�"%�b��O��<Jp��(n�h:!Cc��
�'��˧�ԁ>=R�M�P��&��<�J���� �~��M̧�ʱj(ObpR�Τ~N��3�ś/�L���ObrV'�0.�q��
��E��5 �H,o��	!�*7m,P�X�OA2���B /��{E$���ƌN#����O �,���	�L�fu�߿>*p
aI̝b�AX��c�����Z�AH�����%P�H��ɠ9��֤�,n�D��G�'h�\��j7��(^�N�0/^V�5�S�ӭ��P 0oZ3>��1��.�,B�1a���RDڹ�� 
il�C[�a�@rd���H�d�Ʌ,F� �[�J!#6m<E������1|�4��%��#�"ٲ ��sjS
i6�A&�K?B��,	4cq'6��b��<$���E��V�C�  �H��y
���WƁ��0?)��]6bx�4'��]��`��@Y>��Oįg�p@q�[|���j!���0F�Z�lb D|b�_�<�P��%�Ŵ[F�O�ZD@b�L�p�RD0� S -�*���' T� ���5"(��eM�� =��'�X!��R�q�օ��T�"~��� �aaK��m=zAx�.�@�<I����6�YG���;�td��U`?����z�V�S�+�^(����F�ԻBI��KLA7�a|rHH� ���Kc�D�8�;7!J�n�,�:� ���H��fO����'7��UӤ�ΦF� �U�	 <��0�ݕ�,8��F#�6�5k�+Z����l�<�@�c"��âA�Q��m�T���Q�4�9"Jl��H)O?��*A�����!=��X��إ ���I*+C8=���=3P��3���-6�tX���H~Ɣ�1Z;#z��`�E��I����cD�?�o�&5�/Of4��/��D0YqmT�^���b�'#�0�-0����O�HhP��a�`����*���㑤F%��<g���?�O����CZ;f����ҋW��j����F-�:��!&��6LrP���hʧ$�d��ƫY�Z\��Æm�8��M�������5��Qsp�_7��r��Q�H+��S�G��t�%G^g�$��
9�缻u�S=1�Q�ӞS�i@B���<Q�K'��>��a�j��Iص�ʺN6��yf��.��o�I3�tS��uG�-�OUўX ���	����%/�30���G�"�O���e�<18bh�j{��q�ɋ�*��j�MB��m�2O�>���d@�3�x\�d՜#���������eHâ.������؈}�V�م��y�D	!�H@:ѩE��9JE��$�yr���?a��3�
VqđY�ѡ0W������pEp�G�q� w�s�Z��<u�v���^�N��Do7�O9����h�iʳS��0�5�_�Ō=ؓ�OE�=9ql��TY��ف9��4�OGў�
P��1s�l��|�K�8+��Q��dղqj`�Fƈ���D	�Z�F['W�.�NL��� aO�h���B*%�t����6	y�,�:�O6 �s�W�8Ӻ}��N�\�� �k�~G~�7�˧=nd��"a<&���V�<۪]�cF���9ﶀ��B:j%V=; �� ����"O�����4KD�I��ΐOJRZG-�.Q��l�Ĭ��~c(�$$�5T������H��ƀ0�R�9�hQ��� p�l��&� �Dt��')ْ!��(V4(�� n���>��D2�Đ� ��B�������\7D�J��- 8n�5�3����K܋6
��CJͦT�̠Dx��9T�L8ˇ�W�l�����!^��ƕ�7���-މIB������+F�
�O�.V� �'~���VO�v��X��J0}J0���(���i�F��N,T ѣӑ@�����^�2b�y�DB�O��w��� "[�o��0�`��$�0��'��h���A�WG��q�\�a�N�ZHi�b�@�SO�$���]�e�^��Ouyql_�Y��b��!�yG�E� }d�*0F�c��!�����0>y#`)@�D��Q*M2Hl��A�>7�j�@P��8^�r��D�'d��1��W*@�έ�!#�+������R�dGz��`!�4]1H���J)~�P+���HA����S�):b���t�q�شp=�L͊DW���tOp��d�U	�-HԭJ�r3�pj�)Q)h{���	�wD)3+�"���2/�-q���t�Q�<i�!A	(�����?�"!�� ǜ"e��P�-*!\�B䉹�ƍB��J�_���`�!]Ab��%cl����͞���F�Sb��/vl����B���WK�m�#/M��ꔫB&V�J7a|R�L5r9Ru�u#�a��j�f�'*��32)+ol���'�x�)�c���.�	���h��)��9C�׎S㌉�6�	�m~�8C��:���!����]'��O�H�2��~�L�i��ҽaf�<2���9Y��$��U#��!�i����0&D�4�"Y1��<6�,c�#Y+#��4���#�a�0B1�Y:��4��F��-�J�<}��	ˡ�@�xai���!d��Cf�P���ss)��~��[�C�Ot����ޟ��C%�7����A�����5��� �n��"��ϔK0NL��+�O�Y�uj�0�d�i�	�=}X���!�)8�
A�U@j��$TNyL���4�
@�QH8*0��ѳh�'l̪�����\��AJ�7��@��ҜX�T�# ^�����y�M�'���=2��@�*P���'3�B�"@�UY�y �&@0���!�y�F�q\�	��Q
s���Ȳ��-Z�Dl�m� =��2����l����Y�f���㜊ij@t˄�M�`)F��Q�[h��¤U�8�u�jD-_E�4���'Ӡ�xX�,����)u��\�עǇ�?-�,�&�Ը�K�C%xB5�	J�G�ܬ��]�,�*��ef��|i�}� ��U�wk����΂�8��F-_� �P�j��y�A
�{P�ĩŐ���\�Dh
@�
X�͍%�xY+0M��P|�wH?"1(���IJ>v�%� �ad̮eF�RE) �&΀1v+�^F��X2i��*��:'7�םq�'����P�� b���a��o~}(�y�i��/�qO��l��+�\j�
�I�D"��D��D՞Y;Y��Zb��}��	9�7l�:���.ѭ�`J�@~�0�v@<}X�@��B(:i���D�T睋?�nq(2�ԡ�ҵK�aP�@�P��$���)��-
��,�Z��@�l���q3mߦ�M���c�=�e��z�����K4~� �>m��n2�ae�	&'�
��-U�j{6G|�E�a,�8��,I#^�O'�-�ƮB�~�̰	⎐a~�E[v�Ȣ-l*��c��T��)[b/M��u���*qΠp��'ͰFa�M�~:�	Z���5i1��%���9O��0�^%j�`oZ9>T�ujE��<D�<V��WP�U�5$�~��a�Ҕi���v���un�����K�ڀ��'�*���OI�p�
���O9�,�9���鑧E��.I��QJ�0�'��	�o]�|�8����E�mz���X�"G.=�I�\`NE�"o�x���*v�<@8����鱟��ǀ9��W�B80Ӗ��#�8�A���%�`p�P
K~�'#[(i��\*��C:9���f*�8����r�ڇ%.��'e�:*.r�����OL�c�@��bP!��ޙ{��!�8O�X*b	0�ꜻ#%�<���&�Q����k��=�w%L�Z}<ʤ)�5j�����c��\�NSI�r�¦KC1d��%�Q@�Ey��ME��a4t�0!�|�@V!�y�FU�Hؐ�Gj<A���h"���0?��<t*����E]�7ފ)y3�̐ d$��/F�<y祈�w��FNB+A|b4��MMA��~�ʎ7U�|���%��z��>q��#>yaϋ

�~�8���u����Tk�L��fGW`̘�S�H��NT�"�Dp�vUs�|��G}�]Q�2�	�
���pKF*�~��^0}�1�=�O�  ����t���'�U�Yx���a��%_��Ã薍WXT���K؟(S�Ɂ�B,J�[I��$VBy�4�;D��Y��3��B��9s�leY�%D�8�l��=�3A
+:mD9��#D�T�@�07��D�@��4A�ls�l6D��/4�X�ݭv@\���>#�*C�I�L�0`z���${���i�5TC�	�QTܑ*������X$g �M-�B䉾	κ�鶆�/v_|UH�ߧCTC�I���`��'@�C�ˊ��\B�F$zy��o�KWx��7\VB�)� �К7�M,
��eJ�T�3%<aض"O2���"Af@�S1�@�M�g�'D���3(��Q�l�Ku!�$`~�[!�!D��BF�^ļ��G�v$\�ɳ<D������3w�P�_�`N(X���:D��F��8&T�{�<O��4F,D���᥁� X����G�=`��//D�Л�)V�.��G!�z��@25�+D��2#�Ø5j(
�X6�6i��#D���,�2XM� ��i�2����v�6D�Ld�ɀRW�I�O0eȊ�yB�1D�<Ca�O������G4z��hó�3D�qP�R�.�\���G:_���"�n2D�L��N� M�TH&��+l���b4D����ƈ�>a���\�@5�3#4D�0 �$ۺK,��TCŬ ��;��7D��Qfɪ@�`E�A5��Dr��6D��Ys.��,�Z)"���G^�8k8D�Y��@���س�\�(Q\�`��5D��c����J6+�,.���6�7D�А���gV��W��G��9Մ4D����ݟ,nŨ�/�!Y�`�1D��� L��%䄕x�N�+l���<D���U,�+ج3��7d�:��A�8D��� n��Cf��7o+o��ċ�1D��;4�<akl�.�qlx���.D��!v�E�s�$ё!ݵl�Ec'.D��bE$P*A�y��C��$=���.D�d��K�2"p!�O�1Fd[@�*D�0��8�<�cGB�x�ۥn(D����!�+m��;qi�Z�Zt`��'D��7��IzH�څC�",��1C%D��2�D�~���"E�J����#D�0���L��p�
]'t8�٥�!D� +2I �ZӔp��]+y� ��І%D��JAf��T�,Djc̛�Q,T����9D�k���+JXR�i'��+hԎ�8D������
�AHah�%o��"ƍ6D��!��S�Zj.�����?$b�:aj1D�p�6d�c`�{���#1����!D��WkD�>�(�c��[#�Pyf$D�P��IE�Q.XRgӥfb�T�ǁ/D���d��k�����-(j���.D��r��̈Tc� /l��:&��B�I)�����M�Eu�}�`ĕ�F��B�ɂ,\�x�Ċzfd���
j��B�	�}M
��A	ڐ-ш��,���C�I�%�|�27+�b!��E�#TlC�I�f��Z����)|\��V�A�
&�C�	�]��5��WS�x�+��4B�I7��A��`�.ir2Iɦ�D�iV�C�ɀ<\�
e%?-vp��l�Y�C��Z�K6c� �q)��R:ZC�4�Qx���4��a2s�Ҏ	C�	*�R��#�$
�`D��8@�B�&��E����
u�h(��B�6Jl!���)	+�u�%ʼ.8B�I5O5�����5$Ǟi��H0;��C�	�tq��fs�<�j��O&s�H��|���v�8��$�x\��ȓv���g���\���+0Mո;=fi�ȓo��|3�d�#"Y85�g�8IK�9�ȓjD��T��93�ɪ����.i��ȓ}f��Ʌg���rI:�vr���S�? �A�U�
	����;[����"O�e��^eE���'V�|&|�u"O� ��O��Q�$�B�O\�N}k�"O�xʄ��.��iS��(�T�W"Ox4����6�Z���GG�6�P�{�"O���ŉ�1'��2�埄���"O�e2��f pL�"%D�b�X�A�"Or���>N*��e��M��Q"O�`�w��Z�6��-W2�����"Oԑ#r�ڜ��[S�=�fȢ0"O��j�� �<���@��Ws4�b�"O�H��(�!<�pCs�
	\�Xr"O�� ��]�/D�i�o�U���"O���G�Ђ,�д�e.K(zV a"O�g��~FM��O�-�`�YR"O�� `��J�+	{2�b�"O>8�T�%��89���Ghر� "Ol�cHF��P�4�<4Y��p�"O�̳�`��4�ȁR�S�-$��C�"O��z7�7 �<����{-j�"O8�1���i+�d�g�H���"O��[�٪�ʵ�P��TR�"O8�;'��7o�1RPi�6J*�y��"O��3�O�2v�������9� j'"O������N8 �@�fZ�P�b]�"OFY��lʼ-����ܑN���S�"O歘B��#"�0�y���k�lQ[�"O�`�e���&��TjV1�����'��I�[E�J��Q-�Ҙj�$�05`XB�ɹ;r]�5DR�������?Q��C䉚E\2Y"U�v�IzU+]�UZ�C�Wz�ul�@���
Za��B�	GS,u�v��+sXJ5�lӝW.�B䉝#z�I��/ämAn9Y�
P|��C䉠Pa�(�DC��T�2�'/Y1{��B�ɼ��y����Iaj���d؟:C䉮&��m�v��C��49�B��1`�	#�aǊI}�0q�&T�JXVB�	�k�n)��O�Xe$ꃭN!c̀C�	��ĝJ�!�L��-J��N�SjC�I�-'��覃���1X�*H��:C�R��Ej�7S���¤7D�rB�I�=�4��	ˤl�t��Ζ'`��C䉖v�ܡӁ���μyf��g�jC��h���U'/��`{�@�D>C�ɼ/�M� ,R�"
X�)t@��C䉔�.�CƍJ�����*��	W�C�I6�����Q�~h��##�.̈́C�� ��q���<s3�)Db��{/�B��0gϠe󇭏M�jQ��
��B��8[�	�b/�	H�~Q�gLUo�xB�	:A6����Z��\�Ja�NB�;l��\�p B' �`�EȬ�"B�	?9�h�P�L�O.��C�S�S$B�	�?ͼ�P��Qzrj)�jS9��B�ɔB�d	#w��#�P����Q *6�C��5 � �D��%$P"�hr,O�'P�B�	�0���d��s�O]�`B�	!dJ��v�3:yaE��4GT�<�˓X����#E�����Nјj��ȓo��4�]�h��2" �`M�ȓ6,6)�PbI�S�Y�d�]UE�`'�\F{���"P�MH�j1g�D�U�'e 7�y���:9�E��Ū

�L�+���y
� DD)��0^
�����j8�i�"Ot,[VK]�5l"�3)�`/�qt"OFa����11���	��< J�
Q"O���dP$(��mC�]�]Tr7"O,y �'�*W�V�/צ@22�"O������#)���	�oC�f%b�z�"OP\�E�V�2��m�%P�l����"O�*�"�SH:��Q���Z�"O��(aN�>U�Q+@��Q�"OL4(�P�9�D@�L
w��e(�"O����[�a�Y�`��<b��m�"O�E{�*�  ����X��=	"O�̋6+DCH�YPN�� �.�CG"O��iGᔝ���1W��f���"O��Y��zI�	� �q8�V��y�m�%GH�=���#�īfk��y�D�%`�`U"�ʪL� �jf"��yb,��dnz1�p�M3W��p���yB��,7�8�B4k�S\D]ؔ��=�yB�`������F�r�z�%*�y��H8��p#�D�7�Bm�oȗ�y��D�RS�=X�e��*�< ���B��y�J�7`dY��E U�t��!��>�y����P`&�=#����)���yb�߫r�B2�17�Ψ�p�M��y��[#ur6�X��R���|C'E_��y��%~9r$N�+6���V���yRn�1FnDe%j�>#=����	��y�h��@�08�V����@w�V/��'ў��ք2�F��B��i��Ů<��-��9�����=�IѤ �5x �D{r�'6Lh�H_=Tj��K�`�2x�a��'ź��_8we�i�eU�y�t�'Y&��FI��>8�jP~:	�
�'��@a#\�;�x8c6�>"1���
�'�@��w�7llc%$��u"Ua
�'��Ti��C����� �"[Mx�'�>��ƀ�[0>����p'�]��'^ �)j��PeG�(a���@�'D$a�ݨ3�^ݡd�׈B�����'��xC`��Ct��kkp�K�'� I t_!������0ߊ�*�'{zQ����I�T�rЋ["#�6�`�'�&���HA�i'�@@w�Sa�'Py�6a�S�|�s����
�'��a�L�'v��)�g�!	�	�	�'Ԭ��4A@}E�š�ߴ��R�'�<D�Ԋ
_��V ��u� L��')x�[��Ӫ>X-	�솓n���'72��Z���#p*ʘhvṭ�'�v�t%^7��x4��/_l��9�'q�M���A>6���f�""m��C����H��}�V䃞7[�	qԥ[�R3q��"O�t���C�L%�H���{6JM�"ON��� �m�D�3G�Ө8��Z@"O��C�*"t�bQ	W�_<rH×"Olmz��ԕ
Ie��g�+a 4�u"O$�2fO�'��e�憂��H��p"O(l�p��4U�R����ݨ)H��z1"Oj�ɖ'A��Z���B07�-@""O�HQ�\���ƪȩ6lYr"O
`�'i�2㆙+"��&g8�)@�"O�<:�O;�$]�?����"O*H���lYTj��r4��2"O� �`i�k�Z����Y�mH<�#�"O����H6;�j@*TN@ =9�I��"Oȁ�$�$d ��-ʞ&:Tk�"O���2�ݏ/������I�%�"OL���?�)h"�t%�9s"O�t�H�"u�
�Η�E,v���"O���GZ:K\"E,�p9N�0�"O�-�ai�6k��2��%U�E*�"O,�%��;	%��b�+7���"O��s��4 �䠅�J�F�d䱖"O$�83Ȉ��	V�٦:���Af"Oj(��/Y��MCԅӫt7p��"Ot��A��F}��K�D��'�pC5"O�l���Z�l"�!���U	*���)�"O�`1�B^� [�Df��q;�eA�"O~����]�h�@l`p��'O��l�E"O�Q���0<l[�/Q��ę��"O��K�E�s"���O�s�ܝ`"O )��DL0U,a� MR��t��"Oh��o��=\�;捄�z�Ni�"O���b����z,`s���e&d�R"O�(X��S�+u:T)&G>|� ��"O�� B-6���«�>b؅�"Orɕ��l�@����]+ �=��"O���!mG�o?|(x�)P9]+R�p�"O�)��.#�<�3I"%���S"O������a$oI�8�+�"OF��S? W�x�Ĕ�7�� ��"O˖#�.9��A��W:-��0Z�'9��aS�WKn����% �ȓFr܉7˛&a�)	��Zzhh	�ȓ��MP`�H�`�����M�֝�ȓnkN���)��L���YG��ȓ�.�K�ĝ�H�4I3���'@	�ȓ��pĘ4p� ��ĮM�h׼U��,�f�h�%֗��}�l@�
�������H$�Ɋ�JDJ���%KQ���ȓ�P�k&%�A5���"�-bؖ4�ȓ^"�X�㗈hGx �S+B+$�ȓ	rK�?{ ��� �p{�d5D�D��c
�N��S-�3vp�*7�1D���g�_	#(l�(�Ȓ̉e	+D�H�e �?R�v�#��Ĵf�z��")D�H����s����B,��Eh�*O-3�i�,g��ߥ.%>��"O�m�"F��Tk� ���9�f�Ҷ"O��ðFRN�T$)�8U��a�"O֔� 
�2X�z$-?P���r"O�t�c�	XXc�� ���B"O��5ɛ;�|HJ�:<�u8�"OD���In�F�ʆ(V����'"O�${�eV�$`v�@$��)44��@"O���T��&Ju��@��Ս1~�\��"OF���K:�tQ��,����ð"O��2���/��˒"E����"O�XUK�2�y*�@̗x��H�"OԊ���G��ti W�S�I"O؍2K�;B8`d@�!I��!�q"OR��W'_f�	0��4b��Q"Ou��>"��IsJ�H��(��"O�,ҐE� �P������F˜�u"O^Eh�LPG�lً�o�7U!]:U"O����J���ԩPD�F��$[T"O|5�!FG�0���Յ��X��"O� �Dc`.ɆW�8�hP��#h�AT"OP�k��8L+ hZ�_�H]qp"O�u�5Æ!z��钴��r�,X��"O �2VkE�	�2Fb�	֌�bv"O�8Ce�2�����A�<yʐ�8 "O� f����d���_-)y�r"OT5K@,�u�dl���E�p�y��"OR)Z���)Q�@�(W�冝��"O��#N̊G[�]�"�ة	#"O�)`P�lmt��aA<��"O� �l����؃b��ٳ�"O��3򄔭I<�H��B���r"O�u�QB�8�E��ak�*��1"O���z٠x��Bv}�da"O��҃�Qph�oZӎ�1�"O�y���˖,@��9Q`��9k6"O�}�$HB@�Ҍ(#�	e�8��"O�C`�05��Ek���?da�I�"O X*���2 }���q��9�"O Ѓ�o�'�Z\"��5nt0�5"O��j3IU�\�
5�+��ib�i�!"O(�ؗ �B����0Z�=J�"O��󒫒J�nh�������g"O���e�[Z�0�CA?( �"OZ���dG=b�id%�@���"O��kR#ā8��Qjf�Έ��1e"O�)�W�	�#B�42qB7GkN}[�"O���6+ۀ>C,��D a^�x0e"O�%�CJF�\����ŀƻ*�2"O���&�߾F0�&@a�q��"O���F�
t��Lx@� V��#"O��b㌽\����NV�>(�s"O̡c�B�E �EH�:jD�u"Oʱ��C�j@�{��S�i�H��A"O(�F�Y#��0����F�Y�"O����N��ђ�D�7Z���s�"O�\"�ϴ^��5��G-�xc"O�������T��lьi��<�E"O��e�_:G~]B �K�FN�LC�"O�1s�b�%/|�H�,�9:���a"O ���ʈGp�C�%�AX��Ӱ"OX9�g��Q���嚥R�<��"O���aI0��`R�!�$/7��q�"O�䃧hŉIa*P3$ մ)�^���"O:QH�b��u�@2����FŪ�"O�mB�MJ���vlCs�ܝxW"O`�AuW�u4X�K#�h�#"O^�s!�T�RX>Es�I�˞ٛ'"O��Q�HëT�V$��H�v&����yb-�����ԆR�CC��`K��yBc��O�ESB��6gt�e �Μ�y�!�i~���'_��`��BQ��y�X�4
N�3'�'"T��V���yB�r%�끨�iF����&f�C��"t�ܨ7�~O,���Ӻ(��B�ɔ[b���g�;L�=x�h�C�'��$�D�8X}�9��)Y�+�C�	���kRI�>�pd@Fn�?*�@B�	�|O@ṐGD�`�c���2B�ɷnG��:"aA�e�zXBUN�"P	B�I?/� �[& D ����L��B�I#@KTPU�I���( �C��]LC�9a#�8�B`�2++l])t��|FC�I�N
��ڢv�nI�2�N�,C�)� 8���D�<B��i��ٵ
�]RP"O�<���s�򝙆i,��-�"O��&N�j��\'�T�<���2�"OH9A\O h�7dI0�d�	�"O�ܺ�^8/U4�I��F�i�hȃ�"Oh̓�IW ��`�COX�� �2"O�P�aG��U�$����?;c��ۓ"OD��c��#(��d��ibZ��Q"O�a�ׇJ��<�0#˒$R�x�"O�D�$��)6u�5ɷ��;¥"2"O�رƤ�.<Q|��	�,��"O̕*�-W!$����& VI��|Z2"O��Y�	M��L���T7"��Q�"On��3��B2��a�͙r����W"O�cU)E e��j�����䂱"O��03a-����g'oL5��"Odͫ�j��v�D]
癧dXf<�p"O�����M�H�Ӕ%!eU�ũ�"O���'�)!2��!d�~E�$�"O�3m��K4�p�fH���K�"Opt�ǚ+ �.;g�. �p��"OL��vo �!p�S�� �1x%�"O����I�@V�@�� \��"O|`h�E$X���GȌJ���&"O0�)�Ow�1��F��~����"O�#�"C��p ��3����"OZ�X�5;H\� ���"O"�
 N�hVh��!�S��Ј�e"O���O2�ڐS��={"O�}����~"`��P,�3wE"}��"O�@ÅoV�g��9�s�N4�D��"O|�R$	ٱ9���A�T'?JJ*�"O@��#��Y� T�hS�9K�Q�"OL-��$�Ve� �%�zN��3%"O��!���zBt��:ҜjG"OtUP H�s�ޘ�)���"OL�xOM�
���A�� �U"O���' Q|�k�gk�(�"O�	2�fD���ؗ-�a��](�"O�!�w��m���IA
� Z�M�"O�DR�!���]R/C�2E"Or	ec�&'B*���-Ʋ#���A6"O́�#(?�|����,P���["O�)`���l�T����'�H�"O�i���0|h�͙�#uv���3"O^�BP��>p~Зh�]2�i *O��[(?�Rɱ��ӐS����'�Д�����x��ȃ�vvh2�' ����ŗ� �4�26hW�sɐEy�'��TCb�¢a��򋒶7Y~�H�'��131m��vx ��%�.,W�0��'�\�Y�U�H�={�c�9ψA�'Ô�a��ԁ>���릀�M�$H)
�'v	p��=(���.�z�� ߓ�?��O4Z��C� �:D�	�O�¥۰"OL8au�èT� �� �!vߪ1�"O�Ti��ߒ��	�e�7�:�*T"OԤ��>� ñ�G�7�aг"O*�R�mԽ�@D�cC7��Z"Oj���
�r	�$�[;�t!B"O"px�a�S�(�aA�3�\���'
�'��T>�Ex��Ogt1��_��dT4.ܷ�yb�ƴY_�ı�H�$Q4�I@.�4�y��F5pJ`���+G�d���(�y
� 2D�v��e��{#._ +Gļ��"O(ts�ʖ^�>���\(�I@"O�Ay�e�`���PB�zy1�"O"� ���'�P��4%�y�v�'D�|B��8�)Y$,���3��I
�;D�8�s��<Ĝ�rc�A�:g�d���<�W��\V�MɖI՘'����R�`0��o�?1��pQ'�[��\�ȓe*�������x��ئ/C�R8�ȓB8����o#����M�jC��ȓejĭ���a�f�`�	�h��u� $0���
�x��%�ȓVy���D޴�(0��
Uf���CS�\�� �U�d̼"\f��TB�s��Ȉ�hCРآ`L��*tN���G�sKB�ե׵(����u �$��L�;�>0�qǜCyx0�ȓNt>� ��̃� a��Ë́G�<Ň�	T�']���BfA�t�6h��d� ͒�1��y�,}H�-94�ؠ8�hWC�y2`X��м�r�Kfw�q�G�R��yB��Rҩ�1VX�j0�u���y�8C.Ԥ�oW^%dmh%� �y"��|C�H@B�S�=@�f���y�@V� ���W+֚ILh�Ċ�y�Ƈ#?��"�ױuA�|���E��yb�D�]}b3�Ҟ{�Tѳ���)�yR�D=m���� �#d-��� �y��_�=�݋#!�� La#��y�k�GY�R#@�A���y�*ؖj&T�@�K�t��l���y�Y�1p���$iV��f����y��-#�L��c�]���#四���hOq�����]�&�n�x��\'R��1"O��`,��]VB\X!�M�@�	��"O���5�k �P�)ԟ0B��"O+)���@9(ھeY� D+�v�<���	\'��)N�u�rsǑN�<�1�ҩg�J��S$�ʡi%�Lh<9Ƭ�Zl�a�C+ ڸe �hš�䓧0>�uKE0AپȑG��o�J��@KID�<�O_		�����h�H��4���B�<i�C�\�*���E��yL��(���@�<������x�bQ�U�9Q���E�<�4]����Z���n�$�p@f�<�$��������~�p����^�IA���O/��K�e
P S,D�h�Ԩ*O�=E�dES:,�a��/�ZX`q#
.�y�`
��l��u� ��Ш A$�y�e�<a���*Р 	���!c�(�y"���j���U#�BiC���yb���:Ա��}�t-�!���y�B٪0B\��[�yMZ��F���y���2��#S��� �5�%hU��y�E��z�F��@@��L������-�yr!\/ia�St�C+4�H�aD�y�AE�X\�U�Dn�)\���yR�]�c�&�2�띆'��9���&�yr�;D�h�d���ԉ(D�?�y�O0*p,TI_?>����ƌ��y�B����x�I 8��A�����y���/ %��I�b� ����yr$
 E�.Uq�P%_�L�P@iV��y�FC�t��91��N�^�ĭX�$і�y
� ��cga�01���!�
�6^6��"Or�����,8x���ҡW��Q�"Oh�!�h�5>]^�pV�I�V�����"O�@ydaޠ|�`	���.�j��5"O�h`��U=5V���,��[[d�"OX��v���r�d��ӭIW�ʀ"O��x�B�mU�D�DE˗(S��`"O���bFJ�\�%k̀B:���"Ob延M۶�)@��><&ք"w"O�T
�%,��D���N(��"ORUP�i��X���*T�@�%�"O����|�$��m ޸��G"O&Q��ރt��QdB�qPP D"O�	��i�}&�heO%fph"O�`�#�Ũ=���	q�F�yc�!��"O��5���[T��LN�)�"O�uq0NKJ��n+^�\�L���"O�Xص��K��݂�鏮G25�	�'h��Ӧ�3X���3mF�}AJ�;�'#�p��L��ƄM[��FMh&��'O0K����|��\�z���"
�'q��(I�+�L�&��
��j
�'z I!e-�E�� k�W�}�Zq*
�'1����vt��W,��I�'T�-�qJ]�A�j8��MzLa	�'�*|���^�:���i��Q�ň�'�!
�^�r���	 ��� (���'�3�u�"DS�C�;{�5"�'�h�R�*X�a� 	�*���'�̱�A�[�+y��Itڢ�]z�'G~�k햨]�T|`T'
�)�j� �'�,q��M�2
d���m�/�ı	�'l�]ࡪ����$�B'r���'��i�&؝Q��M�C��>T�x��'�*o�	��h3'���:	�'�Vm�g ĲuDZ��nߩ��m:�'�n(C��}/x�����#G��!��'%��۳���G�\|{3+78�B���'�N}If!G�/�P�؃��*e�^5��'��%��fa�Ը҉@�7
���'���� �U�R�H��V�~c&Ժ�'��e��Mɓ0�bDR�u����'P�D"��Q^
H
��@z��H�'r�E��m����A�A"|,䵑�'�@�2̅	���s��4s���'��8C�E����KשE*kf�M �'~�X�L�U��
�C��n���+�'��i2֠��H�+GèlH�d��'c~4�D%@/m�x̘�f��bo,�
�'���!+ư�Ѕ�uI�W��1�	�'vA8��AtD�âM�9P��e��'���{��^'��rS��|X�p���-���b�B��D(3%ۮkÌ�"O��E⃿?`�uł�m�t!��"O⥸Ї͉��,k�c���X��"O�-�F؍��1�� �x��'"Ox	p��@�F���֪�^���"O���2Ո2t��6	0U���!�"O"|�D���XJ�g�K]HS�'a1O�Qu+!5d�8�ɶm�vhQw"Ot�f$_�P���K%���h���
"O�p�@ ٮ��
`�>K��m�"O�x7�"w-&����� �qD"O�A��c�JT��hH��z���"O� D�y� x�m�f�MȬ=�"O1��]#@�Y���Υc����'w����;����}"f�8W���^���r�,D�8�6�Փ�6�BE�ɺP~��d�/D��s�n^$)�Y�t�

e�h�%,D��#� ��v1��Y���Bm\1ZJ*D�����j0!������(ÔK"D���E����#-C�9�&�֣$D���%L
#���h�A_�
Dr@�.���?	����0�)�FN]e�:���DR/_$�'�L5 WiR�W6$�"�,	%���'�l 2P�H�s�x��J�
�J�Q�'��U�C�\>kƔa�싺� ��'ֺ��.]���A�M9>V�h�'ʦ�RE�� `F��Ĉ�N�(���'%��1���F�
t��&~�d�Rϓ�?���dDx@¥��˧tk�P��o�l*�OT�h�$�`�.���"O&��l���2HS�V�Q����"O������LwH��c�_6I&��(r"O��" ���f�{�#S:\�{W"OL R��?k����&�3J2V�`�"O��y��ۯH�����4�:������	۟\�Oά��e.��C��1C����K���b�'��\R�֏<Pl}`veާPO
qA�'�(A��- l��9�  �l����'c�|j�	SְM�2C�'�ި��'.�+��zl����D�rל�H�'Q�U"���v�iೊ�fF9��'�v��.��8V��N�ĕ�ߓ�'qj蘓�%V���)�D�;�V�c�'V�5�t�Z�L"��qdo�+7�6���'�9�t��'l,ă��4����
�'호��� �������%=���
�'����aٷ~<��`B/�1�(�+�'[�E��k�*0n��n
�"4�X��'���0@E_i���[6��F�}p�'�^D�2	Y� G�#����B-	�y��j\�AÏŨU��l2M�
�yb�tr�s��*<��!�5�yR툝i�@��D�5:^¹�����y"a���I�r�֞D�<ȚK�.�y���)���G��gdL����!�yb�Ӷl��$�C��;e��E��mH�y���D�=s��5�����m��y�
�*7H�CB��0>�,+n��y�"���T�y���60�F�y���y�\�G��3�8���ኣ�y�'X
K�X9���L�*�.<Z�C��y���40�ؠz�,Z+ZT,�1����yB#�o���#��޴��d쌹�y��^1�Bs�Nþh����D��yR+�#D��w��,F�!#�)��y"鐎2�.x�N(�PP*�y���v2�*R*pX�Cd+��yR ��%�ީТO(�q�琵�yb�	�N�AB�N�L;4h��y��5
c>}22�I��@IsmC�y-�m�  `uR�@��Ds�˚2�y҃=�ʴ���(;�"(@iJ��yB(��Pw����R�9լ����X��y�Z�s�D��QjX�-�v�i�Q=�yҬC�!����]�\�Y����yR斏�&��a�ˁ]m�A�vn��y
� IH��AesZ�Ӡ^8(�d�;�"O���eeS+�F�S� R��1Z�"OR���sk��K�O�-Q񲭣�"O�Xڷo=�~��@�*$�h"O�lkf/�S��!����%J䬻"O4i�A�^	vy
՚G�M3C|�Sw"O��@
8\��P�H!l���"O�E�C,X�`Ԉ19")8�.�Pd"Ot]�7���N�p`�Z*Z���"O�x��+R8Ab�qck�*�$<@w"O
<�E&H�9�T���,_t�e�	�'%0���l�䚕�#iJ�3�B ��'iHq:�5�h�҈ΐ,p;�'`�����6+tA+�kC
?"u+�'+&�i���0<%gLY�7/��)�'6\� �>�<<"Q��(; ��b�'�jɣd"%l͘pY�G߃-���I�'#�R�m�9��H*������1�'�ʠ��
_�� lړ��!)+�� 
�'R2 @��H9v���f�#K�j��'�4� E��{�p��%R$G��q�'IVŘ@�H���CJ+���B�'�Z�����H��q �A�%G��"�'=V�s�@�v
����O��,��	�'��K�C.,�ܡ�h'/���'C�\{�Y74	6p�SJ�F�2;
�'A�ݒĆ)�e�$�<`��+
�'�^AY�.�SN)!@>=�6E��'4���FP�(J�HF%EyV���'$I��
ۯl瀅#��\�j%�
�'|�K�X*��hI��Vi��r�'i��!B�X�B��2��a�v���'�T��Bm��@�*l���֣BW��	�'�`eK��9X� ���>��$�
�'`��GU3|A�H��*Zz��	�'�Lu8uIS�9���� � �&�a)O���On��$7X28Q��E-�H���I !�d�)BH�g�LT�P��'!�E�!��'L ����,G=K�����o�!�ā7*�� ��8Ǧ�JEI
J�!�<�}�C�
�(}+��M�:�!�W��(q!��<F��E���Gu!��
�~�åA
xi�`#�d�<D�I۟l���+dP �S���`���ŹYNB�	%2��"��PL��F��E��C��,&Ip��ū�L���d �0~��B�I�,� H�7y��#�b�lzB�I�4�眎��ݒ�i2��C䉳L���Q!���è�XE�YqNC䉧$�&�(3	X�<N�����.a�����>!᨟�E�>�0]��qAǢ\�y�F�NT�ð�H��(�+�yB�/�m�G50@�ꊦ�y�+��iJQnQ 2 ����yBC� ��mI��!2��u-�&�y"�G�?<���gi�/���C�����y�ŶF)0(	 Ł-=�a ԅ
�y��0zcx�C�N�?(���^(�yb��O�"�I�C�:��@���y�M�-���d�Ѫ���S�R�y���#0���S	��~̙֒Q��y��&� e��'B2r"�	@&g ��y"��>L{.m�D/�f�P��� ��yRf�7���v�Z���S����y
� ��[�߂S,�@��%�ʼh�"O|�S��G�P�K#$�(�H�S"Or��g�؁$Q��z區`B5*`"O
 �%ԵB�j���P�BJl]�""ODhBW�Ӑz�53vL	6�F"O��s���z�΁��3d��ҡ"O�t���̩hY����+m�:�� "O
��U�V�PL�i@�AJ�ܙW"O@������=_8,�%`ԉ�15"O���vkޙ#�l�3�A3I�����"O��NH���mH�I��*"O��cD���;6�:cmҿ,��D��"O���t
:"�\д��Vټx�w"O�������D�"��*L�L00t"O tHb*@�>R����#;�d���"O�V�2(�<*7$�L��"��FQ�<�G�D=q��I&��-���̇L�<�pG�\���5mW+}P�:A#�p�<ɣ���1�T�I��W���1cŀU�<yu��]�~�cr.JoL!*E!P�<�Ԋ0C}��X�cN�,ۮ����W�<�a	-?�,JqȺK���Q���P�<���Az]*��:I�����J�<!%L5�f�K�c�/F�,Hړ)KE�<لG�;?�����/���i�B�<Y��'Y<VZ1�@'Q�vm	0FB�<y�Ŋ�|�;�j)�����<9t���"���"F�Ց X�����Qc�<駇ق�����Cx�Q�V��W�<�K٩bހ܉B�K�,t�� �j�<iIı!��@ڒ!�(���g�<�RW�@��$JU��j���%aAh�<��G�E� �J�%ߔ: �4�h�<��G�_=<�+��s�>��U�_f�<9�G�lͰ�*�(�4I�f���$[x�<)G��K������w��U��ot�<�b�A ��:���[(����Y�<�6Ί�

���B�|(�i"�Sn�<AՏ9}���A��~�xW�k�<Y7+�;:��A�sE��~
(��d�<y��U3K��0�Dþ����]�<ᭀ�@�5�D?D���J�[�<��,I1>¬�(4ȑ�$�0j�G\[�<1խ\6����"M>�ҩ�� X�<y�% �+GcL��LAâ� U�<ighWg����Ɗ /����C�I�<�&kڵW�dh��/��S����ZO�<�D��j=h-��Ը!�|�G�KW�<�1�Ξ؃E��|���D��}�<!��j㜁ZV��;ļųf�A~�<y4�=C�6�0U.�,P��$Y��}�<i���	!%F�A���\(�GYA�<!`���l�����_�)�m@0�?D���7�۩5b�R�����A>D�<�bC��h@*���lS~"��3�0D��I�F6E	��'E�������$.D����{�=����!i�<���-D��J��Ğ��C�꜌q~�%��!D��qF"QG�AG�G�_�dI�"J!D�9���!p%y���e^��N D��2c��6h�tM�U�C;�q)��#D�\��FҫJ���b������!D���@(:3$���j�'0Ӑ�x4b-D���R�=<�*�:��ܰ��j�J*D��  �a�Ƒ�e@U��\1�|Pz�*O4�yw�N+K��C�%ȳ�����'e4HYB�].v�F�(�N�/��s�'N��&�؜n"�ʲ��T 	�'))
A��� y>Xaņ�"��ِ
�'e��A��5z�<�ʚ8c�t�!
�'�48�c���-P��k�%LZJ���'(�h��H$x�R��E�E�B�'I�4���ͯl҈xre�?EIޔQ�'� ��l�<]q��Z�MѬ5t�0y�'��!��
�H��,PZ�v�;��/D�p#劏�L�����(�THAR�,D�Xi� �-� #.��$��U��?D�(�w�� t̋J��ղ�7D������&�$�#���-lCH%	1@4D����mZ�j7��a� 
�$I���?D��ZQH�*�,C�([�TO�u�b�?D��w��9?�Ľ��X���`!�=D�,�&��,%9���C#v<�a+Ph<D��������A?��*��8D��Ia�_�a��*5���F�����#D�t����?!o�A��H� I���Ah3D��u��3�p	 �[1	�l!�PD0D����A��^F�5�v f\*��--D� �1�R)Q@ؔ2��-#I�B�l/D���U���6� �Eo�:)Cת-D��������
t��b��Gkp3!,D�\�BN�&M��I��rQ����5D�l��1;k�Il��cJ"�2q�2D����̈5k�5�P���"���/D�赦ЂB���
_�D�*��.D����[��Œ��.|�J��/,D��*�����~�������Ǥ)D����DE??H�q��쌬pS�@j��1D�:$�Y<n{�=��얀H|�qF<D����S8p�8л�`3�>��P�/D�@�B)B;C������	�hI{Wh1D�H����5`�y�a˾v"�:��:D�	� �H; �㬕9:��Yp0G8D��a@ʆ 
�(��K���@Q*D�p[J��y8����g\��J}@rN#D�0S�c�3����`�l��6�&D������ �e�rn�*[�FYX#"9D�L⧁�4,����aV�$%p6g7D�̂�`��`�$���ٮ�.}f�'D�LI�(ȼf����3�f���+D�\��s��)����A�\ٺ*<D����h�xH�3�Z�n2!j(D�H�ާR�T�j�o�a<xRh0D��rQ�Ce�ř F�]c8J�j(D� �!L�I�ؔ����nY�|;c")D�٠���[����ui9xhY�&D�PY��*��
��@Q�İ��9D��S5A�56�!�U�eӠ���#D���S�V�z@���A"��ub!D���1:H��� �^y��E�+D����ګ@�X`�� &HQb�/6D��1%�7Z�� �)h�B+5D�t����)�f�C9�	I�-4D�dاkT>S��9[b�?�k��4D���u�ۭ7�4�`�� �����-D����̑sN�� 4�;=�R|	��*D�<��֤w���� f�� �J�Ba)D�TԪ�X��I�Q��4�T�Q�'D�� \L�叴H�.�����	,&T"O�4ASD
*���Ünx̤@�"O��;���,=! %� rW4��r"ONP����"ذ�J7�C�2K����"O�9F�ҨU>@SG�3s���V"O��V`�4̀&�.���{a"O�Q�&/�_H�N?"�����"OR��`'ʝk7,��ㅒ7u858G"O��q�-Ӆ�����a�4[���6"O����ԡk#ti4���u��"Ohm۴a�m���@��]��H��"O��ĢA]�Ɣ�g�[�@q��"OX-��
%>-*���; jȘr"OJ
����O�`����>l4Y� "O�t[#��g�j �@�E�f��s"O���GˋgX�	Se	د,�\D�`"O�<Phll��u�� :�Ta1"OP@f��5�*��ň�p��u"OMHP��z�=�G�| �"O,5�IĨm��)�eќ3 �!;�"O0����Z��)�3dŜ�ݰ�"O�9Hs�ٛ��9���(�( �G"O�	+�E'Z��q3��֚	\�U�"Ov��/U�	xb�Kg�y���S�"Ob�a �ָZ��l�'=��[�>D���a Ǧq`:�s���ƺ	��<D������4᱓cZ�*P�m��=��0<���, y��HբD�7�n�zP�Y�<����*R�@�x���C�nm��UV�<1�E��q�}�1E��;��<�u	L�<qv�]�_�.���b��0h����a�<ɠgƜ��Kt��W��aE�G�<��I��",����-�9	�`U ��\@�<���Z�
 P�CB�!s�A p��{�<�c!ՓP1C�N;�0 ���a�<�t��7"� ��rT6���sD��C�<�l�N�hM�B!Z�'����+U~�<�t΅ML�"�J�� i�[FKy�<9&��7�tDi�@ȧAH�a7f�[�<	`Ǒ:���R�!�%+q�2!O�<�`I�(x�M�׊�%�ƙ���I�<��J�-�� �M!j��t�TF�<���A�J���{y@3�LE�<A�؍r���IP�Ԕ�V�ʳ-WL�<1G�F9Dup��S�:R��LVK�<)��;dv5�I�'���M�m�<Q��YI����ǔv�l�n_�<M����AL,)L��u�Z�<9�6�
� ���
%`��ӟ8���,O�H;�ʋ0��B7�(�,�ȓDi����G�;|�f-�6�E�hX��P��k���-%�&�cs��|T�̄��<����/ò��3�� ¨���9�`�# SX��pm\	xD4]��j�Ty��f^+,v�d2e��5P���ȓj�@3G4u�u� Q�<m��ȓ@���&���L�&�	�j�$24���b���R�`E�+R����-!V�rЇ�] p@��ʔ8܅q��=`��ȓrG��q�M!T[�=	�-��;U���?�*���4-��dI��_4^��ȓS�v�{E�"�<q�1�D��#3N��2��:�Д:���	P^��ȓKr��!�Ț�h�r�#�v�u��S�? N�cd��6�,����̓�=��"O�l����6�:��p��K�(x*�"O�5�@���t�WO*x\��!"Ot��E@Ur�ܲV�V�#�&H{�"Ox��3f�k����W�����"Op���+Ǖc���	�2�<%�2"OVMp�h#DԢ4�$�ԋ\�P���"Oup���s���P�I��4�x�"Op�d�N�n�\@��(�A�"�x�"O��I6ON;h�i���Oe���s�"O8�x���;�(�7�E�Z�cC"OJb��P-���_f����"O�e{phC�*�P=�VIE$zo��2"O��� �ŚcQ�Y��5>�A�g"OJ\1$��.�ƅ:��	<1t�"O����S��m����>*T]�"O�M��%�Jظ�3�D�,V��"O� SըE��F�ȓX	v��"�"O ��Vh�(K 4��Ù|�>\���'�ў"~�&�ظcvTI(/����һ�y���n�*2�dٸ��1���D�yR��q�t�$�<��i!�V.�y��N>P�.T�D�U�1�>�Z��ղ�yrc�'n �X�4�R�"#����� �y���7�0�3ț�e�=Y�Ϝ�y­O�Q�p| bI�f��k F��y��-o��d�F� ��*�s�h���yrI  -I���	~y��S���y�'K�!g�E��0z������׃�yr�Z�&��<���1��wç�y�b��1����e�bɂ��yb�H ���hƠl�bd��y�ʚ�q����ԥЕuG�0[�gB
�yB�4
y�P�2&R3i��-)��J��y"��\�rt�J��]�Čʁ�yr��72^��W�84J�l����y��Ĭ�dy�5�
3[�|h{�AG��y�됬l���(�f�5<�2Ls�A͙�y�^�hڸ�� �:��m��<�y��vV\�[���H��}�G'�ybjT	����cl��D�v�Ӂ���y�̚e%��vM:�h��GV3�y�
T0̂���-7�|�3 S��yҍ[.O��F9�� �E۟�y�KC�[�\CA����>p��.��yR��m��H%J�]E"!k�����yb��z����C�O�x1��\�y�ER�P0�SK�W+8	�rlZ�yBH�	lR���H',j`�7�[��y��ײ*@�B Ϛ�ZD;����y�m�" E(��I�v*(�
��y����%�&�ˑ�Ќt����e���y�!R�j���A��7J����y�`ر/�pu��O�.J���Z�yr��~n����2+Uf`�F�ئ�y"N[+	E����*V�/@2T�T��=�y�-Q�`�3�� 3	�SԢ*�y�kG2aѣ��.u�hy�",���y���;� ��T�P�Z�Ec�L �yb)<BȨ�aF�Y�|�Ђ�'�y�EU��6yAEǮR�b�s#e^�y�fS<��W�)CS��K� �?�y�!Te�q��A�V0uK��@�y�f�-,�سB�ѩ2u~�{AOU�y
� ���-�.7�԰�ߓ�vl�"OV�(FAA9�N�Q���0�*�y�"Ol����VvȺ�`L��fi��"Oa�����	i T2"��@�g"O�<6aU(��0%ؖn�e�a"O"ܸ&f�'�ppq��U�E~нB�"O�`��ݐ�Xh�A[(&x��"O&�����(�����*,����"Oz a⡋+e��m��ʋ))�}��"O�|����*	Ti�!�F�B�V!S&"OR˵h�,E��TM�Al"OV�;q�@�W�*�x���(i�Z`"O<8C�יon4���m���7"O�尗�)5�Zl�dP�[�"O�E�#)*W�X١��&:.��s"O����*Lq��¢L�<,�z"OH�T%�|��A��6%@��u"O���0��\`���tV|��"Ozh��(�<���y f[�(�,X*$"O1"g`׋
Y�u���S$��$ g"O�Ճ%B�T:� I0�ϻr��}ҵ"O�,�v�֘-�Pp����=I�,:�"O���&J�����ʡ��%��ɐ"O4�pU �#�����Xw\�P�V"OnA24dO?*0��W���IB�9 "ORu�ϝq:�����8xN"��"O��B�eŁG�MPRM*�v܈F"O�4��!\�">"D!U��n�d�3"O@8
fJ�"����y����q+.D��5���X��M��ul��w�-D� ���0~T$��.F�X�s6D�ԛ��	� ��� W(� 6��E�B D����-\V�nؘP���a�?D�8�C҃A�h��b��С!�(D��@3��`f� �,կ$۞�X'D����&F�UK��3���4��Q�%D��� 	o� ��"Y+s�� E�$D��A`��_(�)W�>vVE���$D�8ZS)Ǒ"-��)�F,Pm D�$�#��! "��b�m��86p=���=D�@)�D�/Ŋ]�b�@AZA��e:D�P)��S�rd� y7KL�bD�%i"D��u��UR^���<��A���?D�`U I��<��h����-�1$(D�ġ��cC��SQ��	s���0�3D���@M)��������Y1D�J���m�܅��f��!?�%ҷ�.D�(���G�rx�8���'m�����9D���b�׶�*��HְLeZ�`wb9D��*��H�E�`͙�O1>mf����5D�Tk�Α�%�`��$X��	�@5D�hPu�P�[�q��K�AKd��%l3D���qJ�0P\!���{J	��g2D�(�"����n�;C@��+�ڨ���/D�L�ď ~KB��gN�=D|��k,D�����Ǒ4M�!�gW;++($��/,D��ّ(
6Ϡ�{W�	L�DLq� ?D����	U�N�5h��� ET� W`=D�@%��<@9����Bu�4�(U�9D�hc�M�y�v��s�"[w�8D����o���,�!5�35��4��5D���%\1E���'�N��P5*4D�H����Ae2uH��_,Z���!(D��z�� ��}1G�,w�v|��!9D�� d]r�m���4�V*� k "ODQ�E-��4X8e��O��r!<�*�"O�X�TV2�"�0�.�"=���["OV��@kP7cb�UI�k/�=�%"O4��8@ p���Pq�ix"O4�����,XaAQ)O�	m�z5"O:؈̳S<�`�C��,XJ�d"Op�q0i��I�h���1���i�"On�%��e�fm3�xj�Dr�"O��Y@kZ!!��%.XM��1"O���1�Ž��s�^)t! 4"O��p&0J�6�a�@&;H�s"Oވ�d^6j���,����"O�dAccQ,�b7E40�NI�c"O����V���ʷ)lO���"O�#�P�H�éS2<@��aC"OR���F�q��@InP�M$"O�Ĩ���o��h
 �OKD��"Oyꇯ��6��[@E@<F�H��"ORm"@D�=
 �0�re�0;Db��"Oʱ(1�F� R�+T�Y_=��+�"O<l�F  ��ף�5=R���"OX�K��ɀ4ǔ������$a"OLJd(AG�t�q猕A��#�"OVt�� U�$n��j�l�8�B"ON��vC̟PtZ�����Q385�`"OZ�)wcǑ2�t!�WP�b+x8��"OD�ِ��/9���"�"D2~yr�"O��
�ɵ}��"O5<�E!r"O�� vR�F����r`��fW�Ii�"O�p@F�Ǽ5��sF ^�a�.�z�"O�}�@ �R�Ӕi_�'�L�"O��w�Y1�ՙ5KЂ���G"Oz�@��Y�Oc:�Dh�|�U��"O�9���� ��b��T�{�� `"O�!��8��2#� ��`�"O�La�aD:^!ꑱ���)D�� 
�"O$\��M�UZ�<�t���Y�<��`"O0d��BMm�B�%B;��P��"Od��Gm�5k�� h4��=8��!)�"O̻���LF�8���"N���"O.`���T�3AǮy�F��h��y�JW7P�drr�l; X��� �y�[Kt4h�,��>H�W��y¯Ħ|9��q�Z��(Ru�;�yR
�=����H���d��yƱm<�h����d�I��yr��(+3��HBS�}���j��� �y���[��)`��
4% �؈�C��y�u N���F�A�U�F#��y��P�f��p.��=��jaI �y�
��ft ��읤���Z��X �y� � #>u`Lĺ�B|�w&]��y2-��H�a������Sg)޵�ybH�xF�̉7N�3GT@�G��y"��<o�YCF'�&}����%�y��A�+k�4�7�P�N�T�7��ȇȓ'd��#��^>*]҆N��+���ȓ����-~���ڃ����8K�-���UҹQUE׆�B剹4ՎYI�@��hu�sb�c�ZB�ɬ`���C���0hDPՎ_^�^C�I+m���zg�׶y'
�C�G_0;�NC䉰$�����Kٞ���$�0>�LC�)� n C���!2^���˜W�M�T"O�(af�O�"� d
�4� f"OvȚ�nWM̠�׀y���1S"O��栒���{�(>t��Y� "Ob�#RmJ�����@�ЊmZ4��f"O����͐�4�pQ�GR� N��B�"O�I��z��	��>2��p"O����B�MR�Y�_*F ���"Oʝ��mY mG����ӕ �`���"O�a�$"��1�A�X�t��Ly�"O�m���&���j�k�<xT"O�����Aй〪��F�`��G"O�$��,r�8��hǡ
�2��4"O�[�*�!��(�F�<IGl��S"OX!R#Ҽry4��5�Ȧv=�I�f"O:	`�m��_�d0�,*e9�Y��"OPM�A&>T� �
�J'@�"O.���R�a�D A1��&��yUO��Ĉ�i�|�)fĎ�
�!3Q͆�V�	A���B��V*o�3�-�3���I"O84���W�
�����ʻJ����"O�р��
vJ��0��I? @M5�S��y��
8d�
��q@F�R�@����M����sӀ ���G+\�h� bțstBp�"O��y�%8���3J9l�p9�"O�Q+��a�a�Ƈ�-] e "O��+�MH
#����a4N,�d��"O�T �ͅ/v�6	�7�V1JX����dN�°<�\�l�A�j��3>��h��O�,$ C�ɿG�H��I�D����c!L2&��Iq��h�8�A"	\�M�D��A��G8h�Y6"ONUw��k�@9�Aj0�!"O�5a�M� 	�qB�,�=^ٙ�"O�ͻ��Y��.=0�ZcZ���"OI���̮\5"yro	=Gd�ѳA"O"!��o�>6>��C�hM�����'�U?��
�t$� a�7��������(�O�PSc��fô��4���r��=q��'��D��j���*䏄�?����XP�������gƾNC����f��O�Q�&?�H�T�IQ��u7�G?�B����#;D���+�y"Z�`���KM"!�e�5���!(C�I�.�p�2�/�7 d\��CȨ!�"=�O�d����Ȟg�p;3GJ�O�aᶈ�x�<�T�̓\�)gl��,1�Rx}�;Oh�����,O���i��1K�`x6�)E�\��"O���h��b��%��å3]<a�%�� ��ɟ/�8�4��,5��pb�o��{���$�O㟄M֚�LD#�EO;-�5���'D�@*e�վgr^L@���G�ą�0%D�<SF�*D��/L��9�'�+�B�I-|0<�¡�\�������LϤB�I`EX���x�^h��h/M��B�I�y���S�H�v談��3tI�C�IY�z1I�hY�fUh��E�3"p�C�	�|�œe.�:K�P�ic��E�\C�8u\�x�MȞ[�ޔt�N��LC�I+
ch��'ܯAql��
�.B���m��� �0$�Ma�j
�[ �C��y�t��A,v�Ȩ����~K�C�I9X>Τ��Ç)9׶4Kf/M�/;���d;�����m��Gɩ=�Z���ɔ
`C�	+9� Q��[�6�۶�%h�bB�ɏ;�t�+7JD�#A�fg��H��B�)� ����f��Ũ��5)�<;ST����Nmft�a�� �K$��1�PB�	6u��\Ɇ����z�c�@ HB䉡H+��ʵ�
?^P�Ʉ���g�D����'�r�' BO�~&���'!�QWlL�7(���a�BTD��'�R1����`���+�&*G�a�'��k�"�~.hő �E$" �@��'�.aH1f-~x�.L�f���9�'�6P���vrT�!���?Y��Mj�'2��I�F춀y� :� ��'ܔJb�_�ePvaq��)��L�H>'[�ԅ�ӂH$��*B(��u���Eޟ�C�%<�N����SXF	Q� E�C�-{~�R�oս;�E��]�)���i�(����uO�5`� /�������W�<�B�C�?d�a@��T|(���KJ�<��*7����f!��&�H��K�D؟���j��k������&�V\v���~���S�?h(���U+T*�2��p�C䉓1�̬"�A^\ |�t\ڊC�IJ�J�9���6����9Hf�?��S�O�r�'��ْ���+~2e����tV��'& �����XwB�$��
�'" �ө��{��ʥIɯA�b� 
�'#�����UB�=0�A�*1�d�B�'�ў"~r�'����r̍�7��qC-b�<� h8W���Q���&�X�)�A^�<Ar�\)N���X��q!�RA�'�ў�'?��H�e� ��o�r`هȓP
ġ�w"�	�^E��AQ�y��̇ȓd��0	u%w� Ճ��ܦ>
`��ȓh^�ꐫP�${�i`N��q�ȓ5��p�['p#�����-,�t�ቑ;�Q�L+t�Yh� ��F�-�`=���9D����Bڿ`�8����;�����H:��N���O8��
R������Z<+`E��'`�Y�o��*��m�g��lI"�'�IȆ�>3Jڨ�vhT�v�����'K��{��4]�z���M)`jL�}"�'�q�� �$��(��%�_���b�'�b��p�Ҷ+�.m;@iU?%��	��'���" ޟ{��xW�12�2-�Ó�hO��R 営B;|�{���5�p����O�i�.O���~Fzr�<�"�Z���1	H5�����?��'�*ċC(B�\X�C�9N�N�[�'�RM�W�(�8
1jE1���	�����HE{Zw��ah�1 � ���:'�D��'f"���fF�*A�#�KYPlS�O&XDz��i�/dɺm�g��:��
q���)�d��#����L݁�]�^�@=@�'�ў�}��
�Y9T*B=<d��6�s�'F��F�4�2b�X(��4x�5��*�?�y��UXB���D�5��(����y,�_�HmːF(	2� �R�I��y���t��Ma�FE�>z��FkF�y���;Bs�x9�!Z� ,6@1& �?Ø'yQ�4�}�c�ʅH��=B&
ϾP�
��qoGY�<a��(.���V B<K��H��-R��&���1�߲U?��T\�<4HPpI!�O�)�eCF��~$��	�Хh����4������O?YL�l�R�L��(�PQ�nC���a5D� �0��7:��
@���>��3&�2�I�<����)�2��s�F � �[p,	
�!��U�c^T���F�(z�`��Y(H��"��@��~
� ��k[�EۦCr��B���I�"Ó�p�%��Ph�*��6��&�iZ����Igy�ݳhL����B"S�~�����HO���$̛x7,cQ@N� �^TC3A��x�!���d�0�ӗp+T�$ @��'Siy͝�8�U�GS#��:�y��):�80@+�eP�T�RD1D�]����䓆�<a%J�1�Q�֦ȒQ� 1�㯋{�<���� � `��(Q��Z��Xl�<���.^Q��ߠ9��P��Fe��n���O�*؃cG�7li�󀂸pP⭫
�'5�H��/Y4�t��ɓ"|�ӪO>��D\���� ՠ!/_<����M%�!��J�<�KmU��M)яϑV�!�$S�lhF�:g�T*4���s�Ѽ.�!�dʻ��M��T Z� /�>I�!�D��%4���Kܪ	ZYY�..,!�䅹~2�T����#���P@�~!�/L���S�W��0���r!��23�ё2�P�W����E2m!�$��]����&�@�;�A�D��/�!�DS
h�l�9զ��Rn�v�%!�䅘^~hk���`@*$)�F�G�!��1	�=�T��(�t�- 0�!�D>M���ς?wj�P�YLG!���\u4��$N���cS�r�!�8@+�/T�t}qfOPO�!�E|Ðu��\�L��/��@*!�D�2v����,u���CU-�r!��ĘCR��D!��֤q�0"NU!�D�U�8�g͒�"Ū���.!��՘e�+s�W�*���N��~r!�Dԧ[�^Q�s�$R=j�ʇ�W�K!�^��fM �m�9^%vq���J�k�����{83@��
�Xچ�9�yB&��.i�Y�*I��b������y�%ޡ=�J�2�N�!���ag�+�y2$�(YX�+���H��R`�^��y2���W!��XSA�i��gÓ��y2
l��2v��4�A�4	ǩ�y�m�#ft��@v$�6x��0�T!�y���xg�! O�3tu�ï���y /:R �l���j�D�y��=�|쓗�T$M����T�y�l8��T�@�;���i���y2mF<�9�qa��-}��Ҥ��2�y�H�j�4�L�v�$��D��*�y(�o�����o�h}!�%̬�y�⁃Kt��g�;���D��yR��V���Z���\e �#W��y�+,|p�!
�d��RQf��
�;��'^x�p2�L��������!F�R�yr���r@��V働9!6�`!�U��y��8`�Xq����.:�\�P��y�k>��A�ł&�Ή��)�q�<�6C
,(�5�Sj�"#P��b��q�<�竇�l	��"a��79��("�i�<�� � �a)'��/��0i��e�<�se�!�`�����*[x@[���\�<� ��*��"�iэf���#�F�<yd Ÿ9��P���J�@�<i��P�! s��\�<���}�<00Py�$��
Tȁ��Gy�<�3&�
���(������M�QO�q�<1��L5;ztI�* '{֌��g�i�<� j�H��$230�"�!)Ht���4"O���f��R��=j�`���VT�"OJy cT�fz��CA�z~��"OjxP L�zE�����ߕ"�Ƹ�t"Oؤ�F1.jv�Q�g�/g�(��E"O��$̈́%1��`E�($�N�B"O�)H#g�*���%%�dK�A��"Oe�� �<�и��8Dop�C��'��lZ��ڂ;NP�9��_�x�	��H�p4��/����sn(�)ڧY��F����,t�Pe��v�iG{�-�>A��ݹA.�z�'O���4C�$�^��E��O���'|�$b
הD :=�剈/5T[�+O5�#5�NG��B��Wz���;Sr����c�'9z`��.&�*�Q���p��Ocz�u�7±�x������.7ߞ�s�,O����e�PwD�´M�$���dm^>]r�08���Nߒ�C�'���Χ$�^� wO0��x����"b����I�aH�� ��G� mk$ԩ=2I���_�����N"60P9��"= ��e�8y8��0�'�" E���t�p�VW�sƴ���(�z"l٧O�aC�e�'$�J����[�8۾��n��t^�O �I*���S��;�ʂ8"}:<
�'zL�%��F�8�c�âq џ0��I��"tä�@: `x6!e��� KC�I��#bfG�c��c>�b�2g��JF�+|o� 1�A�l�T�Ġ7-��A�p�=Q��%�S)~nhBV.�����	�C5\�Z�1��'`�ց���ܟ6�e�%��1�"TRv�\���a0�����	��B�?AG�
�|��̋fFwx�H�d�D��<9b``W�>����|{��Xp�A�Cx���ӗ|���O��1�D�XQ��-JQx�'���mc��Ջ��}���{����H���-��'�"$�c�XZe~8�ԕ>PV�;b�����*~����b��k�~���ˍ�!/ּ���

�� &N$06�ǾY����@�1�r�i�`�෋V�5@s�#�!FB�x�F��$3�ͻ4d I	�G]�R/�hXR��5^
42���Up�)IE�̄ 0��C%`��T7��ݩ5],*�F�F2��r��׳wr%8���1X�Rl 4�حq�l#����~��Z���o�s��(���
�R�F��}�ڽQ.	)2��@f�\�g�����b�`���Z�f�~���Y��M/
���";�.pSL�%%�Uji�p�N(�J 3̐p��$D����'�Q����2	�TŻ+�A���BAO��D\�!�
�`#�i���� L��-�@m��A��YQo�	�BT�Qʐ�X[t�� `�i���/A��b4�J1T��4"�>�`,T"\��2G�I���8a��"�B=
`�تw݈p
!�L����%(O�̥���J����IX
�´/��_xf��`�F���E�M��ƪR�ӱd�X��q�7�S� v����f	!R����uI�|� �kЇ��l�
5�[�Z��a�w
��~������!U��T�fch�S��QBp�� ��\:z$m8vF���Eh�G]���'���b"�%�pH�|�7��%(I��@.I;��'1i��*à�8�����+<�Q�����tB�	��r���3�d��Q�KM�*RI�H�.�g��8V�`��E*#�����IS
v���[�k�h~��S���Mc7
VT�����);(���.B?	��ś�a��y蘠B#]�$�� ��>_R)��.�)9 ��u.C�������zJ�[�j�C�&O�,�d�3"��gG|��M��XG$̂2ɀ���Џ}�����%�wN�PS̉�7�����I�\^�б&C��J��鏊.�̹��Ԏf(� ���i�����I]D��q�'�\9�I�	z$��!�λi|�	k� `��@-J0���v�֚�Z(@&�ܲ�@3K��ml�i��D�j�ʀ��4����0mM#sL����[al0�3���� ��� ���'Uh�F��< ��.��Y�`�tN�L@]�0k�,�>��vIL�M�Ȭi �U�
�l����<o��LⴎLBVq��+�*�8��&Im��KC*J�]�R�K�C.O��@P���M��KS�zOv����A2
(����@��bܹ�
,]�Xy���9���1�G3����k���Y�GϹ>����u�X���P�IȟPtഛc
\{�ш��ڍyB�d2I��T�q��$[�!¼�?��`�����$nR�,����#5zX�)��hA��E/IN��d��
\o&��GHyZ�ꤡU�O�x��ef��?�T�G��M�'>�\�w��-Ly���-�5��O�w���ɔ�A>z�]��۳���*��XJu�Ǚ.
��`��*t����8v��͵cjI��H�9��͋�&��U�x�`&�)�1O�|�@f����'Yh�Xs�� �0��r�^�)!%�	3D@�/A*��!7)T_f�`��-Pb���;�.���2���1``Ų#޺֒pZ�*GAOkH<�ņ=�.D��
����ȍ,e�F@��	�7{��%���\���bF�8�:h�'J^� ��hͭg�L���7+!�Ġ����V�j3�]
 ~ayr#[/$��u&O�G��FeD���5�5�+��p���ʋl^���W���]q�@?Wp���B���.]��;����(p`���!�Ҵk1�U�;�8ON�Q��֪�Qzp���p����v,f�bQ��'�Y��nƒp�jU�f��8�1�w�I�b$��'`�Yё��Ҕ	��Йr��ab�]�O��`� ���S��/�g��a��� W0�V1�%F�g�D h
�'��Q���1�D��DD��bF8�V^���E2��ĪJE�;�!n��]��	<?)f�c�u���!��9ˠ%�*wVN ����A8v���ɕ����1�<�0�׬RP�ݲ���m��2b@ѡ&%,��0�:H�!�:Ozb2��٢K��'Yi�r"1*�J�~Qvm�?I�o
���eI�Q��"PJbՇV����0�O�lp�P"��[C���`F�|�v�@�� h}�u$����d �g?ч��G�@+��D�0J}�/_8|k��I��͵q�Bx8�D�Z�w�_qwi�}�w�>-"r"�=D�L�h��Z�WN�0A�4EFH���^�+E���)<O� ک���Uڹq��ũw�H$p��8[z�1`��c�N�27��]ޭ�%ǟ Rʙ!&/D*������8����H�8w�qr�
�NJp�Q�'E�̉����~����Y���gQ�e`l$��ń'ˆ���!I�ix%vfF�^B`B��"�ڟBʄ����^ +%�<;�ɂ?Z�����4|�i�}��C\g��c0�٥�
@av˓8Bg.��ufY���s�U�uf�<�4���E�*��&�mB�(�fM NOPqj�;OpP�&!�wb�(�d�&D�(O�m���L3$��r�hHvA$��!M�� +�Y�!��`����E��n2'��B��ȄuF*Ɂ�]�I脭{����2�R��gi��lJ�R@X:vLVx��D������$Ax�'N�r`����Gk��#�2�k�
$Ȧ�(����z��]R��3v�P��,�
����ߧ!�&���˦ͤ�8���Φ��w�$�x@i�*�P�m��%��z��O�L�`���J*�#j�-!�P�IP�]���M&(1N��®�=7����W�xB�R�/�pD��cډPh� �G� �u��K�S��,"��zq@*[x��m��ZX	��F�
����^�"���@@�*d��`/�Y��Qp����LhQP�G��$�E��'���8 FQ�Y��y*F���;�|��u�T�Wjك5*��a<U��M׼]�L�Q�&�?]��UJ��Ҵ?�v�'�X�cb3/�уZE��a�g%U听�V�|���)�oZ%sDt:��Hʦ�8���6��Q��D��O��1	��N�g��+v���\�Jbȍ3��\ <f���+��&���x�\)p+\J���&��H:����B7��� �!>:4����R(^2�!3�[/b.	C�Z&��e�B�5
��R�S�������2E�&��T��d��J��㞟��gI�����ܤ-�v �������0��q���d%�o�8usa휬	^F\i�K�@NЛ6�ҵ���� ��c��I$@����M�w�<Lq�4Z�4*r�6G��t R�^�bD UH�`Ïn���K$��	I�D� :谦��`(/`A
A`�`j�͈���%����&a\�'�4�V��Ԙ|W��mމ��1m���Q�'Ԍ��A�	+��֐�[[wY<mS���<a��5�wh�h�(F��6T�[�lڰ��4����[��
�-=B��ts�N �-�����E��r�bPEθJ���3OS�<�!o��V※T +}�#�/X��Y�Ɂ�]u�UBb���>Jř�S�&�ɰ%J�ow��x��ԝj�4M@�؏^;���&�p>H��R.�ݨ5C�nw��Hw��lp �i��I�Z����cJ=�Tp�O�H�F`��@hO�<`��bCʶWbx������i�9(T���lٸ��RA���8����8Ɗ��񀞩���,�*D��#̘;��'����$ͯI��U
W��Ғ��uMѯE����l_'s�l$kQ��\� ����O��A:��Ƴ֐��ݴZ<���@j0�QP��4�,�TŎ�6-�V�A�L��	�8�b��E� Yҳ�2Ȅ$A�A
1#6��d)S'8ј C���B��A�2q�#�ɰ̌	1��%=�$i�R�!��w{8Q��Ծ3�����iv���s	�$]����&��%�Z�q`�$E+�*�g#@�5��f��MBT�٠q{P9
$n��YkN�)�*�&@"��Gu>=���D�ds�%V�@-xg�7��9�6���J��=rf��#�mo������թ���3g��E��(��!3��a��=���C�ؒ��:���s6�,�sJϽUÎ�� 5%+t��1��u	��P��Uep>��0@_���,[�� �$)p��!���-�WB5;�L�`m�
f�@0ٱe\%������7K��]q+�[�Y:�H�nm�x�ԊZ�?5ё%�eܓY"��B�㌐=�V�P����md��o/<��s����i���#i���r�C̑>�\�h1��im�9��/�O�8ygM�7@͜xC�P��̉�#E�v�t��6W��	�y��	4R��!�I�+7J	�� u�򕩐�۸�N%���D H�P �Lޛ���K�KTjNL� L�r�衱��[y�t�'`.�Co����J�,hMT	����Z	�'LP���E�[����N��n��vDT1I	P�����.Ł׫Y�X.Z�����CR����R�z��᫵bE�YO�� DEI�)�(ա�+��Y/�Ӕ&���$G/S�r/�r�A�B�e��xqeX�%�v�J�`_78L8�6+	T�-2�/ǭq�I�'ZL��.�\���u��<]F��R�
X!&�v��!�O���5�,a��5��/rhr���zy�y2ϛ�l�|y�˘6�y�Uͩ���c�F��c?��y�!_�X�ʰ����֝6o ���+X�U?�Q�7�\�p䣧� G���y�
��:��UMƼ~��$:D
ٙ%��#=Y�mݜ�j��f�$HM:�`�Θ<W���Z�Ƅ1x[�`�Td�
u��3��^�ElV<�E$HO ��^?%R�"�>)e:ibci�z�B�W?|��pt����hO�P�WL� ��8�U��6 �8� �&x�h{��U����׈�+� �� �SgJ�ȑ��3�>A�� ��A]@Ɣ	����F ��*5���i3.sL����q�T��'�>�S���D�Ȕ#PJC�ҀaG;"YP�t�8 s�pa�팛bw:�"#d���ɖ$�7_ʤAz�'S�3B��P�@�kD<M��['`p*�B�_����N>)FꌚC<��S.�\�����M�`�Ĵy���=�0U��*\��TJ̛A8��3nS[�����o�6g�ԜI���|���Z�iQ$tMrQΐ4Qp�T�7��/� m"1'�%�Q�Xja��Pt�@YZN9`i��T�Nu���98D6M؃#(�aR
�+
P��p�'"٘P�������<6Z�&���r�(���8C
*�8�)��;&�#�"G�s� �q�Ò�r�@�Al�)ddp�N��&R�uS�	:a\�<�f�R��A�E�"�����k�t@Q�݄#X�E3ڴs˨x)��-�4�à�
2m��h`�IE��%b�* �nL��$׸HH2 �����($�~P��D�9KM$�$"7H�ǧ*Aj����#6Fr �7����-�Gl#�V,8���"{�`��0�Q�x��jĀ7B~ڷ���	�1�ǜx")���L��m�&.lT9*w��x ��M$ۛ6E�F刹8áS�!<ܽ�T�ۥL^ڔ�nو4(�Xr�]��%x2GԾUF�i2BMQ�;�l	�%)Z�"x^�3դ�� �-�=y���k���i�k��Lj��W���[$H;�b��WQ:����x*�P!%�4`-ޅ�e��Nc�������]����VP4���ƌ�|TL�B��L�wc�5���Q�AV"�u�4�	�@R(��U*Q���柱,��DeB ]R@��� i���Q���92�X�<PB7��N�mRu(K&���E�§p
Y�D@^�U���yRI�X�8XZ�ѷ}�f(�g�	4d�|�Q��5�y�l� |=�<!�$$EsN��|�b$���2i�H����6�i�7,Ƃnb8B�έ,����?t�ᙁ�ơ �����ٞylL�Q���?=J�AN-,��O>�&�-�� ���?M>���!g��ʐ
L���s��e�Q�H���(� Kɼ@$��`A�`�В���vP}h�B�p��p�Ϧq��A�lѓ�׎\1Oݳa(׌Ytܑ���4.�Z�"�!��SL�z� �M��0ꅮU��� �D-F���d�@��L�jU��>RL�jĀ�K��cЪ,ր jdI'&�P�&9�V�_.w4���1��.u1��ȑ�ro8h!k���Rg#��bpq�FY��Y�����Dc �Ʃ\}��O��o:�y��'5J�
��~�8y�O��b���g�;S��y��B�#�Pb���D| �k���y�&"Ql�M{'�I����B#H�ͻ"=���^+8tt�%�G�)n6 ���c��s�
�����J�]�#ȲV�4@�a���X���![�-0�0S%�]��Ь�	O�i��cI�S�&`�E�@����'JZ*ot��R�Tږ���'�n��-��Y!a9>�T!�G��6U�@�Is�t�b%
 e}��xk�j45.�y7lW!_� �'
6T���}��neV���q�vPp����'�pDHFM�2���ֆU��*�	wLg>�YS���k��X	��7f�����C b�p�	��&n]#V�Ϩx4��D��K��� � R�-� ��K�'�-ꄎ�7 2=�B�o�ԠY��,��'��M�R�h#��-1`X���Ҹ�|�B�36I�à� � 0��*j��`�JP�lWj���7�����e�庆e�:Ҵ9�ъ/a��pJѮi]x��S`̙6��'c氐���վ��!-"ِM��$\O@�/�tE�����m1`�;8�6�S�e�*<�����5���3.B�_�Y��N�-�|3@+��{r��40閁�V���g��AlY���'r�� �����i�LTu��
����T	�+˪����V�r� �#���N�@��aLۍZT~� wM"\OhMK��8�XR0 ��$\ikb��5jz�c ���?�"���H([A$J#hDFł��i��4۷��-���A Zk�Շ�C�I[D�1�i�1�n��	�ɴDV��� �6�E�J[J�UcT�~���vC"�i���T:W�D=;�z}�'.��"�/��M�g�a�$�e����ޤxg(�7Wp�ч@\�\�pKM�v�bEW��c?O-�ߙ2~��ë���h�Of�:V�ы*�%�4��?|�*ѹU��ac���nY�HER��ۓ'q]�0�S	R���s�X�\����		Q���/��_���i�i�0���)�\�p��><����',*��W�ܶ����m��Y�$��y�-M�\�0��"¨{��>���k�d8�pNN�|j�`$D�<�EE� ��a��R�>���Qb��[W�@��1}���E���$A(	;�hA��4� Pq҆ſ6�!� ':��*��	U>�8 2��A��CʭL����;��HCևF�6�*d�%[<C�I�-?�(�CH�+��
C��Br�B��)5TT<B��̋V�Z�a�+֗v��B䉐{&xM���J(Z�>���;0�B�1O��AP.��4��Ԁ�;.�\B�I�ҁ��խ_ 9�p.�#N
hB䉟��Q�e�]�R�����FŞB�ɐ"���sP��+��}�Q'�$.%XB�I>y]�A��"�9uW����޴`�VB�1hՀ��d�� ��Q��<@!B��&����*��v$����!�j��C䉺^f�Q0�	��φ��6_�C䉅�H�3P'�t`R�M�l��C䉰']������#��(: ��4i��B�u�q��P�2���
�̰B�	:,���O����r5`��r�B�ɂ6������X�8�����e��B�I
m�2��p��)A���4e�5)�4C䉞%7�R@H7p��tˢ�ʛo�<C��=�f�H��т3t� �����C䉭H|���Z#D(I��֡*�C�ɴi`pYy��U�(r�Jվ`DC�;�(�Dϑ� [N0s�V>9C䉍,p��K��H�T0�Ei��<1�B�8����� �:lB/�C�I7
=Jq�Ƌ)98�es���7BC�	;k�0Tw�5s�9P�fB�g�^C�ə����qb؄q�j-c��=hRC�2l��`ҕO^������:�tC�	;��@{
�	�-�ţ\1\ZC�	�P ����*)ät��A�x� C�[rX)���4 [�0"H��/zB�	�`�n�����Wܸ!�"�,"��C�	:Xdi1u�G�h{���F���:��C�)� ����S.n�dH�G�,Vh�s�"Oa��E=� �q���=OX+$"O�ي#dG�AC�tѐ&�7���Ȅ"Or�x����W-�س&��I�$��F"O܉�P#
�8n��!�Z�!�洲"Ox�����.a#��9㌇^^�09�"Of�`�Sڌ�(��,'iz��f"O��VO�8d�����M�}U,��Q"O����������-JiK���"O�����Y>S����	��0Ry3"O�487)�[ �r4o�;��8`"O�aЮ�.#D53���x7�'�ڦE ;P
�]���a j.W1�A�� ���;减�Q�qO�>1���^���7����j1�E$���� +y�c?���*Ս��t�P
ro�8��'�<��i��UGα�Ì>,OPH�Wd��tܐ(�q�ڮF}ƥH�D4~G �`���3c��b�4��b?1��E�%-��ↄ)QA(U�U7,�����*2(mL����QVx���f@5lJ���+j�*Q�Cŗ:k hI��;i�n��F�%<Pv���� 6lF���'�,�ͧ���/�@���*��?%b��	 "��	Zq.myD�x6 �2���Q�)y(ؓ���b|�ىuJί3�r���
H؄8�'px�D���l�౉.Ӈ%���pʌ�{�ƴ�OP8�A��.�A�R>3;�A����s�O*�R��gFR�Ņ��/�Eb��'���S$�<^V���X%G*џHB6�Ew�b���-�0!
`�a�A�&`�T�9�KW�=�`,3����%�b>	�@�!�x��DU`z��g���8j��
��7�daE�|\�=)�$�Wav��S�X�p���2_Є��SJ�
=��A��<������?����s�X�Z�p�#)Z��*X�?�(�
ݥ(Ty4�E:��tDv�X��!F�XL���>���$�����#�7:���B�b�8^�NQ@A `���f�vղ%��B�A�	m����\�?�O���	��"�~4�,y�,l9�.]b� �(�'n�R��e##?�1��/K�Α8����4G�L2�fx��3��K>w�3�!�kN�	C�Y$s��o�7`�0d��m��g�2�d.A�l#JF?����q�s�6ʌ�i����#H3�.P�%Mr���̈́l����c	2�<x��]>�cr˛�u���%Z�"�(�
۽���y5�`�t(K�[�Ψ��a*�S�n*^�~�4x8\�����4i�z�zQ+�_o��E	2���C8v���o�,1�bT��Em����[��B�hǇ-�L��֠A<r����[D�@:�i�ym��E�ٙT�\	�e�H%P�`�wN2[���A�O(��D B�6{�����+@��r$H8E�b�u�۲{`��
@6��6-�a�]���[zD	�f⑑r��(��7d��8��G�h.9i�Q�FIz ��C��xr��)w�Fbƨa�O�̳�eL;�TZ��M�':�}�qO�<8_̜��iģ0a�&8`��ed��O8�X9%�NI�tr#8_B^����LP5�T�T��&$0v�����
N8�L��Op�H��F9]ADt�AD����"C9-�e�3AE;H��AQ,*4�Ò��:N`��!D���b"�/�Y��9��K�+�������M�W��$�]�7�詢0��+	ڜ���L'��+S+_�����y��-^66���ɛX�&�+.O"\���O�]��"�@��]k+�t�����|/��q��^��ft,@Z�3��,�|e�r�91.��s���Afj�jn�)��;ӂ;?��@ܭV(37������*��8����W�ŧ��e��f��J����Y~ITp*@h^me��� �:����'�ĥ��m�fFZ!J���kXcq ��#	D0�W n!@�+�>i2=�D��w\?5R��D{ ȱ�"E?aw4���#t��U3�4,~�qBD=L�B2'�۷6bju�R'�-N��tiĢu��m{3�'t�q���I�R��Am2Dj���*g�Q$O�
���'���"D���6(: Ǆ�� !K-O��nâ t�����P�>���c�]�u���t�2���S�]<��	�l@���I_�i�^�����C�s�浹ơ��U�A�	3p�(a��n�$� !&;�{��u���hu\��F�&�ʍϻz���K��H2`�]�"I�e��o�t� 0�L�HT,EС�'������P2 ��`�"�P�{q ؼ�~bh� �p��\������K�*��yP2(c$Ѕp�_�;��H�@Q��b��Ђ`�ɉ��'2D.�#�
 ��k֕jdh�"^gr���H��(~6�ҠE�!!�A!F���:����r'B/	RfAIR�U�	/P`MQbb��Dٱ��M��Ph�d1R�lOr���&H d�V�r�C�*?�^��@aVj�0`Ɗ�/%3@�
��ćPr�к��P�7���^�$�ZXXu�M�:�1OX\HU�,��'�TT������;!�(����D�6:����N?1,�R�(
K�ZH�q#����s�R)�����w0�u�fAϕ'Ժœ�/����'���jD�.&P�p�も7�lH��!ЫG?*����2*$pS�|�Z�#R�#
F�8p�5�d\ᇁ��,���M9s)\��
W�N���c1,OP,��k,<�� #	��GW���ϋ�_JH�����Xrm�VF˜|����ę�Z͓�@w���G��.q�$�"´Y��\�|Q`��O/����~W@�wON�O8�12l۵8R����A6{�� ʔA�4+���EEQ3(`8U� �gsdA��
*ܰ?�T��/��dy��ֿU�B$��c˩N� �ʂ늖}�_D�?�'aǭ�8x�.��v#�.z#:M9�'���Zv�V<2�kV� 0pːh1i��f�b��sc��g�L	���z&6?6yݕ����`D�Σ+�6���.H�K���뉯L�t�"�R0$f�����hx��%�7n��P6bBl��V�׈;RDq��9O$��1�z��K��g�? �@���:��y���φfD�̳���H�x����Z�w���Ba�ȂD�WmA�?a:��G��N��$mQ,	Yf��ϊ&2�t@ !J��L�˓�h���O�aXqÕ�Xv
i�7����X����0PU�gP��p�s�+�e�}ҝw���S�!��LRc��o�h�4@v�pBR$�JlQ���!<Oh r�ay�"�@�<�PW���Y �C^'M���$�P��0���T<�e�$N�?J���G�:�;��Z�����EH^�9�-Г�{���Î:i��)q�ըof Y�ۀ!E��7B�b��y��&ѷU��-X�d�!z'�E�Z
e�.Ԡi�8Q�h��%�֡�E�Pm���4�@ru��	�J�S4 ?��?S�-�)R�g��У�Զo*r�so��<�	�	�Ӟ�H�;��_�j�X���j_�~B���l�=5���̓|��m�����B�í���߼�"t��RC�I[��M���[��ʪG���r�d�7 a��� �ɹլ�
$K�/QD�]s�&�����k��K�h	���pNW:p���ף�b�Z�����`��G
�5�1&�	�c�^����i�t��E��
4�@m���N#I��A��.ZM&�(�L'��(-��V�d��UDC1�^]�!	�I��I�i�&4Aw�S�`c���4D��P̊�	�S�YS6M`��L�+��6��k�RAH���Bʩi�e]�x���h&KR�9A,-i�=w]ة��o�a�0�����w���[_w���#梘.Mj�$� �&y��Q1N��p|F�@��T�����Ś���a����T��a�Î�iI��B�ݝJ �+��T�p6�H�f�^/u�ݩPH�:mnB���~�f�Ч�ȃ� Æ&(0�����};�(����idT�J�!��}��q�t}�k_[���¨A<�D���ז.��m��	:'��YDc
��dY��4�0}I�а �fH�ЏQ�/Ws��\�$ |cH�hĺ��"��16��Yb@C%	0�����H~�@�Hj8y'�ؕRt �&�3�d��=7�P� g]-7����ÞM���c��ŏr���RS�_<4�?3�F�p�۟�ؐ�Oͥ>����\�K)B�U�z��� �T�"P"�+w�օ�t���Xڑ#Ʌ)%v�n97������}:-F�@����Ō�+LȈ��S"Z`�l �R��	���R��si��2W6-۩[��r$ͫ�E�
�V�Z���#D?D,ѣH�!3��X3��++B(jD�E�:��$Z�iJ6T�P�����A6Z���� 2�����gI�|mb����Q3[P��Øp��7�*h
��%�O2��@G�yfz��f�0?����=�ӥ�3�$� �F�J$�B�\�8_0�AHS	wc�X�T�C �)����&� �&	K>�� �0=V�����{w����8�LȂb9Oz��G�� K����I��hON�E���Q���__69�-��Du�u�QAy��	"W� �HP\/�vL�#��?����@�>�	W�F�9X�ݳ7Ȝ�m���Пs�0�#Ҩ�:�V,��o� ��O.x0$�ٔ�<�Y�_�~I�'��DؐQ�Pm��BW��i�K�ą\?pBIk��_0:H~�#��v�q,�����؜'���3i��u�k��jܓrD �!�\�r��l#��8;wh�S�����x�K7g�����vC��'r��tsv*;9vd�o��"��a�50*:�˕�[�y��T��(�RTL+�S>]���䑢<�yvD%y���)�0�\�a�Y�a@.�!��K�r%�KA�y
&�"pШtI2�x��D%dJ@�*�A=]�Nu��+̷D�(-��'���z��
�Ym���i�" �~��0�@
9�TQ��0I��x�f�y�������D�d��7o�=�����<�|!�ıH�)\{����ƭZ�!��J�N�F�*q��'�@��i��%��A,Y�9��J�K�R�Xq��
�t�ڻR_Z0&��.;�* ��nX?t���3�ŀ`�6�S˂��0=e�GN8�6%�]%����-U.�M� $D"kT����"�#gl�"%��EL<�;$ur� 2h��]�B�xG��E�PXK/҈T�ij¨�V�X�Rm�5%� ��Q��'��Ec��O�RP["��U�hD�ŻK�/o���c�h1V�u$]�j��)?2��9�pa�TC�ѓV��m���#sH_�F�C��i4>�)�$�?Z�ؐ�B�ZcF�:w�CJt��͹!/�c����k�8#*�E�e�T�u;"�Q���1D��xB	$E4vi��h֬4�l�	%"��h�� a�X(�6mʳB��prR?�I�jU�B�ED�L�ؙ���`2Lz#EO~�a4@b%ϾZP���j�:WDh�@6��5W��{���@Q��4�/FGb��D�F
YhUT�B� �R�ֈHAf�����5AU��;�Bo��B�X�
Iy�Ι�w]�(��Z���|S�@1r���s�eK|�� ��4c$	wY�sU��gNZ:���X���B��FIz���D�d�RŨ���%]�H��|�H `f*T�~7�x�ug�&EAj<�7��'�@|����	(<9���!p'�̠�섖+���`B�Rf� z�"���t�uRR
MC�F��a˙�*X
�&	L)�F��HG�~��sՉ�d��>�R�������3ғlㆡ�DH��IzJ���
A\BM8Ej%z�%�s�E="�� D�W�<Xr��0=|N��"K�G^�?����
�	�b�K�Gx�ȑB���{�j����<@����򮐜 z����._| �{��R�k����4��	�%F�=-w,]�Q/(u,t{ ��_l4��ҥb�����?�
s	��>�4�@sA��h�����M@�;X�!�2���~b�o������"Xf�� ��[Y�ՀV -�x	ⅆ�
kIS�I� �J�ꡨ@'k�YT�M7b��r̔��P��A��CO�@{�Ȯ&�T����%��k �G%�`�~!21'	P2��� }^��c�V q��Pe8n
��ge�:b�jJY+.(t�����v�#� װ>���Dg�.�qC�-_�W j9��9K~V%ɂ�\w�'	�}S�M_2U��d��X@��VEl��}(��i��s1˃Qٺ����4	̂%q���%A�~U��2`Jހ^�:�pQ;Ѣ"#�����V��㟰`�*�<3v���B�&ANPQg�O��p�c�G�<��Q� KZ/1D�:'#F8"�X���K�����d�(u:~�KB	��9��7�׶:Tv�P5FrC>��g� >k#K)%�l�����o��q0b�04�Ήj��^�ٶlN�(.8+��+�?�5n�i��4YP��	6�X��M#gb��"�O?���� b�{��Q0?3�YQv�^�]ϐX8���(Qf
%�cU�I�b!\	I$�VI��/(h V��gBV�m�fc����	�\�R�,�+:��(����+�a&P�y �
DY�����n�PXH����D� 4%؟'@��E���'�@����P5�`��ѕvL���N��tL�P6�N6S3Ui�D ��$K�@��`.�\{��rA�����J�X���P2Q	�% ����<�J�SSb؅�|U�<Ys��n}R�n3$=�3�U�7&�U��h�$$�|5y���(T��2(0���֐P!lС��D�L<�R��d`~)A��G�y�89S��D3*0���Q"��8�JK�@���zc�%}ȥJV��7���i��1[�h�����f5��(�ꋚD�����J'yƹz�̏2�� (��Q!�6Rָ�႗{'�x�B� As��M
~(p�Wb�.2�D6PԼ��"�D�b��ǡ�O� 2�������FxFi���Oܕ�'�`��g�T'I�4c��z����AZ�o�4�bb��#��-ه�-I���_^I��d�'�t��<�5�<$�`���iT72���)�LT��f&��]�tSP�#|��)�d�og����oV� m�qB�IR��vf[9_�l!#��џ&v�e[$.J'?�T�Ca-V�{�`}1f�;�	�z�jaq���4C�@���9�ry��M�c��usT.������bv��ra�z[nр[�?�y�0�Of��B�H�E۞��I��':/������J�ظQ攨-��I�c�H�i$�5��@K�l^��Rk��{�C[
d�>�R_d	��w�`pH��3����G�2U��ٴ�5�c�0�)�禭�����=~��TmӟZ>�H1�E~t��s��2H�6��� ӈ�^���'ǋ8u�<��-R�_*�AE�|vl˧��).m�0�w(P�$��1*�>LO�d(��q�!��oZ<A4rɂ��8,!(<����c�tXt��/���"�/l��y�nB�bղ�����>Af���\�4�"��wn�YCU{̓vd��h�bK�ըC9"瘅ig0�T�k�@ 1�PUH�j��U
n�1�� �N\�K��f�� ��Na{2�C�C̈�yQ��"!�iKm�h+(,`��V	Bb^�UѠ��^w %��SN���mT6, ��� �Р'��T*q�Q������+#XC��I��)S�`��o�L�26���}<l؁tKX3 �����D�d}�'��L��!  �j�\�v�Q�|>n�ӻ[��aA��ĖG|�� ��Q�]����.F�0oG�f)�w����n��b@�Ce��j��]�6�P�"0�G�(�%!dF�,5t�E8c�4��{b��4�ðo�>0DV)���G��'��Lѷ�O�p���ᐠ]F��r��)GK��8o�E��f�v����q�4��#��cUIg ?\O2}� V� ��S��+Ѥ�z�BӶsj���m������|��'÷
��|��M�,����\�Mf�@���
��hH��B�I*68���rI�$s�\|�b�X-v�6�H�.��A"�&+��:�Ҩ20���R�i�&�����
A!8-�f��*u2�j	�p>�ĉ��$1��	)rO�Sf%,��h�KY�k� �rWdM3a��A���'��%�f
1�3�dD$�L�	��@�X��eAC���d�&rƴ��G�
1�*�kg�33B�IB�L�;r$�(�/����=���>@�ոChƯ,�ܠ���Bx�Шs膮/�Ҽ)�da��&	̢"r���A��M��]8BM���y���)J=�2	��9hn*�OG��'ij 
��q^hU���ӨJV�l��bW�M��p�P��S��C�ɝZ��LY#K��N� �!I�M��ѱ�i�4���'���G�,O��)���V���p�FS�iB ³"O��Q2m�D�<�s�Nߢf����'�D Q4��{X����֦Tx(#�X�}��8ەA4D�h�t��Q ,\ˢmٱH�L�g�>D�pK���[��q*�J�]���1D��ہ�Y���,I�h�"� �.D�8K�T�5wZ}h"G]F7�j`O*D��a�쒌��Ȓ���  �����(D��1��"1`m*BM��V�~9b$k'D��𡔅�j`��Ǔ2�TUt�9D��{0͐�
�P3pjN�S�\��/4D���ԁǺ.�t��Qf/�
���@7D�D���G�݈��ˁwKX�i�i7D��YC��m*���ߴS�@$#A2D��16�#��	Y��X�@ �0
3D�੆BT�u��M�9Z+^T��0D�H�`G"N�}pЈ��F����.D�T�Ŕ'�D`	�C��Ql,D����Y���C��Z�Ĥ��f*D�H��oK�t��,�f�����B�4D��Cp��0f�*�v����M��4D���d�h���C��K(IF��*7N3D����#K����a���S�n0q��%D��JUh�
BZib��!��A��4D��	Q,T�f�.\!&��'[�D�y��4D���Ro��x�j��Qˀ9�@�c�0D�d�e�;s�P��f	Iv�=�(�ɎNy��@(T��K�T�6a�b� �戏b�4 �CG��,�bQ��.4}b�ΒX�����=���8b������tD���
p���H�W����0bM�)�'Vp��ծ�^w��ʅcçDH>��w%�.\�H$�e�)���/����u(V)Q�����$҅:w�5󢉞�^�`���?yN�Fǎx>�rp�@�!4���I�mK�����ڭ��b ����M�V�PX��3� ��BӏǆG�nQ���@I^�s��4�zhp�OnB⢈�0|c�2N3�u�c]�y֌���S�1w���ȉ��F�$�P����!�"L�=J�ٷ�C�75�$ɗav��A�>]8�%��?��v��*_���kFFD,	�ɤ������j1�$jI<E�$�՚`�܅k��W�C�ly��%\rZ���8Hz !���"��	(�m �Wo���MǧBʜ�*������d��0|���+@�Z�:��޿B��U��@��
D�E-s���3 D�^4�����ӶP��&Ծeo��j� ˚z}�u�!MKxn@�S��)�?��'?������yOP����%�\��5��	k\Bd��$���HX"��	^�a���RQ�&���M�X֭���n�,uKҘ[�� ��@��a�j��ç�ȹ"wd��b"~p"�ūr�� �1�|{F�� 6�G�~R֟�8�a�IU
��4�x���D�"c�VQ萐x�ɄE�a�䬑�`.T؈".:����ۂaω'u@���#J6�a�d�$)�1MЍ�
<X�E	LN��'6j�"�@�%92O�OO������*`m+!������4MҲ��a�O*\�oM/�~
ç��в���Ʈt�`�w�čϓ-��M�p̪��35n<���4�ܯ#,���-\��-YsnY�@���2�'��q�S>�Y����$)�F֧����`!e=�	��~�����<�Oe��c�f=I�d�#r�pU�s��� v!��ِb���RL�k� Q���	�6I!�$ڤ�P�F�4i�ڤ�ͮH�!��'t�^�8�K�,Nڈ�7�:z!�D(1���h�O5PAPm�3F�?o!�J.@�)O9H�|�f��'kc!�d�<���y!NX���p83�R�_�!�DC<���2��3
�,9[t�L�u3!�$�<q��A�/��=ߨ�����5K2!�D�*��bbET:��PΐG�!�d��1�F4�P�@�%�B<�s�K72�!��ZP�@C�e8x�!H�&��#�!�d�s�HD
�mK*e��[qf�'�!򄞻_f��L�?+YQ�״"!� e�2�(��6���c�N!�E�P<)�c�D�@�^��Ǟ:!�_�cbų�M��:�T�@�!���!���Y=��Q��&az\H�G)
�!�DѮ{�����z.��.��c\!�d�Bv�P ߀i����Ԃ N!�Ė72�"D�u��,~qA�H)�!�䚼O�,aɐ��
wb����	'j!�T�j���'%j���c0.�O!��E���mΜf�����hU�C�:B�ɫp��!s6-���W��hB�I9D�40���s�H ����TB�I�M�����Z$f�x���"�rB�I8p� �]j<e��*ɕ3�jB�	3�$�[�'�'���шF!	�(C�	�?X���Eҧ^�c��5V�B��)V�48�� ��L�a�*��B�I�Q�>u�H��HV�̳ma�B�	L~���F�x|�&Kw6�B�	�NĐ��%�1H�X �%ƛ-\:C䉋'�!ȖG�W���� -���tC�ɸ!��D��+f��r3 B�8k��E��ĘY�u�-Ha��C�	�F%	jdm@%��Q�  �;y��C䉋qi�02v����Z�V�xB�	X�v� �C�5Mp����WRB�I��I	�A�'<<�C���$��B�I,h3�4������=��J����B�	�Q��q+`˗�f������ 2 C�I�B?�������Y�����tC�I�}�l�0�ƃI*h�� Ɖ~��C�	�z$YS	[%I#�{@ L" @�C�)� ��!5t���>a�8�"O�][�iwv�x�΋�PU���"O�<��"�?l(��]�GF�(ad"O���Q��t��]��K�1F��H"O�0��&Ӄz�8���ʏ�I�@���"O~Q!�b�E�P1CD�`�$��"O8�rԈ�x�N�+bjD��S"O�0�=[ ��L�xƠ�"Ot!󀌪y�f����̹!ݢ��v"O8ݒt,�0`9�p�A�M[�.�9�"O�9�s"� (��5Q�НD��-I�"O2] #��#��������f��"O�s6�<���sf�ԭv��xp�"O���A�E�tZHD
\�4���"OV��ġɔ#�$��MP�c~�|��"O�EpЌ��mHtA� LĄ x��3"O�T���6�j�YB,�S�.�1G"Ot����K�U|�P�*<i<�Q��"O04ۤ�ƟA��(�oHGT� ""O�II��^�K2Bm�N?D��"O�p�G��`���IW�Ky-|8�"ON�s�BC�e4ҥ��Ù�"F| "O���G�ޏ6)��IA�=�8q�"On�[c��&IUH�Co�'2a90"OT� ��;V�X�q!��m�1a�"O��E�I$ބ`'N@76 &"O��3��=Hs���wLαy�L�2B"O�L3WL�2E����Iu޸��"O����!��c�M`cH��9w6��`"Ol5��$�7�-cr̎� N	ړ"O0�Y��߳J'lZ/R ]��"OT�5�<6�;S�/e�M�!"O�	Y��A�$k�j�)U�L�F"Oxu���5,��)93��;S< ""O�Y���M�i�FE�'��;EX؈"O�<�cF�o�`E��&A'E�XA"O�8H��J�!��t���65$ތ��"OD40�%
?x3�)��I��(� "O��s���:�C���г�"O�ȸ7��xzൊ D�)]�FH
F"O����E�h�n I�c_�0��B"O0���jROy�Y���� �%�r"O��@×p^b����E�@��e"OrUj��Ԓ,j�-a���"~�0�B3"O�x&�Q�aX9͹J�bT�G"O���C��~�
`��o)o�ٚ�"O�4IB�;LB��P�%.qZ�{P"O8�
D��tUtx ��V7"Cʌ�4"O���v��n\���&���_���!G"OT�@d
��X�"��Y�k:T"f"Ob@���œ2���:a��#���"OX���]5;��0+��X�]\��P�"O� �d�p-��Q/���3A"O�����եuLp����sԔ�s5"O�L���S�H����恅|�ܨ90"O�d�w��Ff�3� �<�!"Ov�`īN <\8�B�P���	�&"O��j��ۅ=���Ibb�1$g����"O܅����o^���0��fPD1�"O�%xB!�.,�(�2dR�.Bn�a"O��c0�v�L �J�wN@�"O�͛��Y
%�R⨈3l�bX��"O�E�s+�)a.��1h���S"O,9���>>��ɴK)s����"O� �]IA�գp�~��q�{��9��"O(x���n$���E	/?�BM0�"O�`��Í_���r�dF2|uj"O }� ��N~��Zv�B={�	"O��HG�H�uN�<Bs�g����"O��EV�y�d0"�N�/i��7"OH�Ӗ�*;��;�F"2X)"Oह�&VW@ 9
w������+D�D�4��-R��qzr�μ��� 4D����̄�ZQ~5�2�߻- ���)%D��0��֙{Ȥ@��A�1R�L�"a!D��9ul��`gV�j�'�P��9��"D��y�T�".��(ۤ#n�q��?D�@��ȃ� Wn}���/�����(D��b�CL<�2�ە�
�?�q�(D�t���ǯ-�~��Q
3K�Yk�1D��3����jyl�؅�F�v$�i*��-D�dCqK��q�hI��~��@ D�4S�I*_���d�}�p�2�?D�h�E�A-|����C�	ez$���0D��X�B>���Z�lB& z|�B�+D���F�ԥ�����Z�(@pP
t	7D��	7�8L�x�b���34��c6D�P)�k�"�p��W�D,j�� D���d�˥?zP�iR+h><�9p� D��Ӗ!�_= 8���3N$���<D�\9��.,�>t�MP<zb�{#�;D�,�� W�Z�Qֈ�J�>�b�%D�h�!<ޖ�G
�+A ܛ��"D��1UF�[�>Er� X�p:�i���;D��Xd۬(C�� 1�Ȋ���,D��Nʮ	v�P�e�C�Xm���8D��0���S��P 5�UE݊:� 1D�x3�a��f��*�ҹ!�6�7d4D�`P�L�TX ��N�3�� �"-D�h[q^k�N�$-�N�����7D��C���	w�j1Z�B�w��d96$;D���c# p��xS��9Q���ul#D�,I �	"�(1W+OF���C�<D�x6O�>?e�����H���
�7D��i�C�K��9�WB�7_X�!�E5D����D��H�4e�b�4���G1D�����)	%�=�0 T�r�8(Pl$D�|���ˉE�����O�(�W� D��9ry�d@1��=P���@+,D��z����ؤ��Q'���ұ�&D���5f�f�ĊS�ц.�,ee?D�h 4I=]�6��a�N�"��`)�#=D�؊5�кp�^X�T)�&?l�� �<D��
 0�`��	!D�P��2�=D�p;"�`m�5gO�E:D�T�&J�<�:=��T
-����+D�<[G�D�9Ÿ�82MH�O�ze8Qk-D��R%H\�(.f��F�p�zi���+D�Ȋ!�S7{�>�bũI�p<(���<D��ZC�!���k��1��C�*<D��zD���+ﺜ8�.����(�7D�Tc�g��)9�V�m�X�{�5D��Q:XsH�A�-j�8�{u�5D�<3֤�X��hyAAӃ�(���j1D�� R�Y0mGd���{��	��A.D�4a� �;Ԕ	j�؝E�v��E-D���R� �
�������f�Y��,D����c�+$n�Bf�߄|Bɢ2�)D�� �Q	ui��F�P<I5���b��ak"O�2��������n0|��"O��1��a� ��@
 nYH�"O�@2��5Ɏm�%'Y2�x��"O�	P�Qr�v���	��Lzy "O������nx��c)[����%�Py�NΕ]n��k��Wp|����X��yr"P2\�$��@n�la�аa�I!�y��N k.�O�	fBz�Y�̠�y���/0w��b���H�J�fJк�y2*J$y�V)5)�Fu�(�MJ��y"�B�w����'�n��(���ynڱa`�1*�.�<2���E����y����(�&�Y�9>�yDf݃�yR�X>	b������0��D�R��y�ƅ2e6�uA7��h*���c���y�(/:H>\K��ٰb3`q�q"��y��HƝIB.�^�~QRԆE�y"���U�D��(V�f�i�-�ybF���x��n�a�@�*7�L6�y)F�
�ʅA�f�3$��������y�Q�Z�\{��ėQ�҉�p����y�J�
h��L������yA����Ex5�[O�:��gG�y2�I2 @  ��     �  d  �  �+  �6  �B  �M  �W  /`  l  rv  �|  �  m�  ��  �  4�  t�  ��  ��  E�  ��  ��  (�  j�  ��  ��  ��  ��  ��  ��  � � &! �/ �9 X@ �F �L /N  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�	�� R��g� �t��B��1�s�Ee� "<E��'�����?l�i�|����y2�6�Şw}��̞�� `�d�ǁ���a����dE�D��p�i^�;>��S��%+�|�L3}2jN,m��+�lRu��iT�y���>�����Q�g�عQ� ��Mˌ��%��|ph�9IV��1�!�;qu��UA؞X$�>�XR��V�ԎPԜa�g��:]&���d(8a�МA��řcYx�h�G��%ڧ\�ƠB�!3]��`��G�44��^�Ȅ�-J�S�d�Ӱ%�'
<�'Bў��$��Fa�,ʕ0�i�9j.!�$�!i�;��@�f�I�Iſ+� �牰D�-�Dk�;�Q���c�C�	;<�4Qd �
����'�4��'��Bm_�K;�HاA�H5���|�����Hȸ-&�tbr�Žp#��v�/�yb(Ͱ6��9�L��o�(��^��~�!�S�Oaƙ�gh�[8|`c��e��e�'% �;?ʡ��� J���
�'��s0i�3y�Bd˖��Vy~9�	�'�F��A�^_8@�D_�M}F��'����7�[�Y��:C��JF���'�*ex��N�d�B��9;� b�''��SѪԮ4	�#"K��7cL�8�'����d �el�0J�g#����'�HS��Q��*�р�	����'a�|@0l�9�0�p�A|�`<��'/x2���93�]���:%���`�'W��P��҈4�����)뎨2�'R2K����y(J�0�D�Z"m��'�~���j�$)ԡIg�0����G��O����^�E�� �9rdx05$?��{rɚ��I�m#��Q��Lm��$*Ǹu��ʉyr�'q�x��H��t��ѯ���r�H0ND$��=�3U����"��M�霂���.�69���ȓAR�L��/�B��ǭ��-����=���?Q��Ӟ6 ʝ)��^�%x"T�&��~�<Y���7?=f` ���4~D|9qM{�<����J�Fa@o�`Ѡ�sS�Q�<�[y|�d[� r:���`n�EB�`�'F�|�ڮe��)҅��F��b�O���	^���O(���b�>�bI����O��p�	�'eF�Js��#y��L�Ǆ�U�
yK�}�x�鉷4��9{�ɐkL����N4Z�rB�IlZ6�+l�	<�ؽ���Pdֵ����'] �cV�`����jG�%��9�'jX-���_�"�ba던�Da	�'�bY��R&��l�� ���$��˓�(O��5,��N�R$�7/T�j�~�J#"O�BS�]9af�K��G�Y;b�s���=lO�A��ydVEk��ה:0��"Oȑd<$�X���$Υ|����"O���t.R9ǎM�1���S
nj`"O�:AJ���,������eh�ha�"O\�!��שn=Ҍ��$�	'�<Y
�"O��#@E�U��C��W�9���"O�؀�J��}:5��k
:�P��"O�D�G@فE5ZA�Cj`D����7O���df��	Y0i؀}�~��)I�5,�,���'���ɉi����AE\���z�&I����5�I�|9������?& �S &�T|�B�	���0p#� ��� �<}��B�I�Jz��5B�% dY��T�A�6�F������ ��A��ƛRTV�BpH�>���6"OL�ke�I�Z t�A��V)(��2dU�p���h��Q#w��
T�� s!�F�H�ZC�I,A:� Iv�CQ��2�iħX+`B�8P��(��_�!�l�s�H�3
R>B�I�T=dX�!��N�ZAz���._B�	,$��rVk[	l��-q-�)
B�I�e|Lru���Z%��� $��>r�C�	0����ThW]jP��-B�6Z��#��c%O�>�ȉ0�F.`�����4�O��$�QԅƪuJ�AK����>���0ƈ3D���� 	F��AƂ�5�a �M2扃5���?�|b���b�c��$��iIGhd�<�0�� T�4+	I����a�`�'O�yB	Q�$�� ��>;L@�cc/_1�y��%&�&aYF.đ-�E �Ј�y�C���v�Pg:��P�7J<�y�n 'Ǻӑ%�0�؍qbC��y�ώ?~�Pt,(t������	�?����v\8���,�H�Pu��!i|���ȓ@��-Ӥ@+n�P�Sd݃B�v,	��O�����!3��q9�(��D���fcҖ^����)"?��,�;�2%��۷�����(�f�<���H��z�eZ�j�
1I�<��l����v����¡К3^lm��	�!n��M{�O��e�k�!�"��"bN؜�"O$Iǣ�W�$�����w���S��D�O��s�{����P=j��1���{�|x{V�D˟̄U24�K4�ҔT�X��CDP�(��:g(I�&�ݱ*�������>�rԇ�,�*I�K�J��f�3��!�ȓ%�M�adT/J�������n4�ȓ�Jt�0o�zB]��j�b���^=�P������[Ôpc���ȓSܐ�bɇ,�����ODN�ȓ&��MJ�� m=j�%)F@�م� �]Y�Fѫp'T�C��J�[@�ȓ?�,�B&@�����1FTl��b3�Y��N��z�	d�.n�B�ȓ9����[��䪧(Ų!xPl�ȓI�@��Q�(]�r�I�Z<��O6�dұk������@�]�(��׈��H $��<1ѧԗk����n�hU�ݢh"69YŨ�<�\�ȓ[�p�Q��L�r��a��_p&ȇȓq_Mb�o˗%�@$�+�# �����<_p�+3
�h�F@�3$����@ua���7���9�'A.S�\�ȓ:����<%�.��P)��(����|��6�Ѯ#���ޠg��=�ȓ-�E�� '��ߓ4�� �ȓ"cr�@�0!{�	�fΈ�
@�T�ȓu+�,J�$��P	�)+vN6Utz��0܅�P/ٮr�\��v!�h��x�ȓ^��`�$5)x,�N8�f�ȓz� 8��O�]1l�RT"�39���ȓ{/������-��$~(�ȓi<ش!ĭ�_<"c/ק!а�ȓi�Y�&T�w�^��n�%4P��ȓ*�f�K�JB�$
��R�ĩ�ȓx?�W� ❩3 �.��\��`�Y Th.���)˯vD�ȓM��R��+�:v�Փ"6E�ȓz #U�$ut�A��7-�4q��S�? ���*E��t��Ś���(&"O�"&H�8��U��e)���u"OnQ�A��r<x�D+^�@:8�W"O�h��&Y���k��N+/���"Ob�p����U ro[�[Ά�[��'��'��'��'&R�'�R�'Ӡ���J<OT���ʗ/p�4���'���'t��'�"�'A"�'�"�'�4�Q*J�$BLc񧆈aR��!��'�"�'HR�'��'42�' b�'���D��'�� �1�u�3�'��'���'���'���'���'h�v��k��<"#��>2\�E�$�'���'���'vB�'R�'E��'�Dm٣��"D*����Y�r<�f�'���'���'>r�'���'��'&����
���`}�&�ȐF.Jp��'/��'���'e�'1��'��'"�����5`�P� �R�F�RC�'Z��'{B�'>��'ub�'�r�'@����k5c@�A�*�-5������'���'�r�'e��'or�'���'��)�ը���e��Ȓ?'�=�F�'�B�'�2�'#B�'7��'���'_dQWhV gg�0S�M��˂�'���'%��'��'Q��'"�'���AЂ��t��!�,�W�'{��'�B�'���'���'+��'u�� coK==�vlz���f�R�*s�'���'��'���'R�a�����O�Ձ��	{����rrgjm(*O��D�<�|�'dv7��%{�l�ƀ�M�hX6�	W�~����d�ܴ�����'���FnM2]i���5�T���*G;��'�:���i5�	�|*��O��>et@2`�h6�IC��s@��<A���$)�'~K\�9���[Uz�	6iǃfc���&�iW6�J�y��	����]2T����l <Px�G[�s�$�I���ϓ���i��6�d�����	P^j�p��?6���S�lc��̓"I�~�����'����J*�h��q�
�#�Z���'~�q򉗤Mw��N�	�|��(_-��h�c>����>���?��'M�I�F'Uc�M�7h�X��E�ԢQe���?��۰Y�Ȝ�|���Oʜ`�z�:��/F	������G�&Ѫ/O˓�?E��'�bi��	Us�ZȊ�#�O�xi�'�b7m��r�I �M���O�P�Î�3x��Ǭ�Gঁۛ'�"�'��$
��v��T�'h���O?Z��B�{��	B1"��;e��'����$�'z"�'���'N4��� B�U�ȑa@)?�9IW����4e���)O�� �	�O��R��T�Ttʓ�̽6}60 ��M}�*s���oڇ���|��'��2o�S�]QsF�Z$"5i" �6 #�հ@OS��� H�Θ �B=֒O�� r5�E6��#'mF�:f���	��M�ЄV0�?�$Ѡw5 ��6��&�"���I�!�?y�i��O���'�7�_�i��4r��(H#��aU��*��Y�4ǔ���b���MS�'�"㘥8���S>p���?��_cpv����P�����%�z�����'M��'��'7��'��O��1;�'�0X��f5V��].3��=��'��Af�˖�3��I�T�	Uy�AѠ)�8�J�,�1��B�#7Xg}¦|ӎDl��?�x��Gɦ%��?���^h�P󐥂�Z��U�ԡ3P�wn	�Y�������O�n�?���ߟ4�� ):0 C��up�1��]�N+�heN��Ok��ɤ\�"4�CM )UC8���џl�	�M#��&<,��X;(G�s�`V�y0��ϓ4���_��yB�'"�f��	Q��]k���OP�i��W�Q��s�i L����f�G`,�xW�8��d쟒x*�D0�O��R�K�J���prCT��2uc�D�O���O��D�O1�
�l��J�l>��#�/Y��ԑ��A�/������'���o�,�R�O2XoZ%�t"���-���Kŉ��SX�)r�4P���MS�IN�f7O��$�!0T(%��'A6�I�<D�3=Ƥ��plԅGfJ}���D�OZ���O���O`�$�|�̏�Tl�x0��ڿD�⑑�É-^Л�dT�d��'>r����'�X7=��P��ǇK֩CEOۢ�f�Bh���شw鉧���O��Ԭ��s���>O�	��-���T��Ân�bpw7O�Щ�-	4�?,.��<����?a�兎l%*ёP��'��i3wl��?���?�����Ϧ�*��S��t��ƟL��(M�h΢�3gCQKG� �����'����O�ToZ�MKR�xr,�'Y��(v�$^����Υ�y��'�N��0�(\l�$:eX�h��r��!�i�bҦ��c�_6N�X[�J0D���'"I9 �Xa6/۞RTD�(�e���$��4�a����?9R�i��O�N�xC�!��ك���?4��\��۴U��v��s���2O�D^=&iX�3�'wC������.���.iW�`(r�&�d�<����?y��?a��?aD
\���	0��.{��d��?��$����FMЂ*���	�?���PyB�� RL��s)˨Y�h��[�d]��5�M��i`�7�K���?��S�n��0�'�%m�TC�'�/:���ք����N>dvčA�y��O�˓l��L�ER��tnV.j�ƈ��I.�M�ej�?1��@�a!Є���Z}L�����?C�i�O���'U�6��H�4x�r;���,x8b�N(V@����'�MÞ'�2�
�7�>��S Y����?��\� R�;��x1dn�	6��B�6OZ��$��(=���цܭDϠ�#�)
c��d�O��D���e�� J"�i��'��ęf�ŧ
d*�A�	�7H�D�G�*�̦��4��g�M�'��ʈhBF�2E�x� 4(�lA�=*���&�����|V���	�����ҟCcٗ^����r�=:�ؼ�㈚����	xy�,m����O���O�˧k��5��$��lА��k�z��'���[��v�p��&���?�g�X�L�h�c�	$1t��Sg�qΌyZ#�V�tE�'\���Mǟd��|b�= 4m�06�$ ZIO�?�b���O.�D�Oz�4������I_B�S��ր�lZ��e�ײFٶ���D�o�8!ȆU�(�IB����$�'-07�B!v�
�t��[S���Ѧ�	%�nڰ�M�&�E��M;�'�
�37�N�_���H��'"����ύ>):��DmM=��lb ��d������ϟ���^�4�t����6�ش�����3`�ܙ��i&d���'7��'P�O6��~��.��Jpn�W� e��J�ɏ�7q�yo�5�M���x��$��5qƛ�1O�D*�&�2.�j�ЯՈL��%(�0O-�S�-�?9t�2�Ģ<����?Y�a��wʄW�:3GD��c�?Y���?����d]��eR�/PyB�'Ъ���[�SgƌB�F�; �a�����Y}҆{��mZ���[��4��ԖP&�\��lG�^�`p��?�d"I5sYt�1�΅����q���n����j�Z�c�`Vb�@��Ѕ��H����O$�D�O���(ڧ�?aTk�"Gǖ�2*�0*_\�:��?�?y�i���f�'�d�\�;�4��@�b	6�`3�Ԇ��x�<OVpoZ�MS��iw�͡��iE���OXa���&���K�;��хe��k�c�0�O�˓��O��� �8|R�Ȼ���1��D�P��`Y�4X	:8����?����OZ��@c�_3k T�K&iHC-���w�>��i2�6ͅR�i>����?	Ǫ�����='j���/D;��b ��Myb���	K�=9�͎o�Q���b���ܖ��A��sdyk���5N��1��8j�X��L�4m�#e�Y��<�&��__��*G��&>	�f�&*}�)5�^�}N�<iu �a�Y��.Ò/�����Y
-��R�=P��B����ɒ+B"c��t�_/It�0���S��}s�a�3�`�7�L��h�Z4/�2-
Ψ�S���r��$��
���j�2ag�Ѱ	K��C�#��x�)u�aF&�dh��2��. ��i�5pH
9����"/򽢀�ty�ǃ$���R�F�*�����J��x��#��t�!��r�d��O&��<��O$�$�#]���J}8����pc��r_��T��>����?Q����,�y'>��@��X���i�(e����r%X�Ms��?-OX���O��� �,W�.48��Z��VӳϏ,!$��oZʟ���jy���>d����D�k��Y���B�	�^�1��G�6[�4�	Ο�P�h)�Ο4�s�N�3�"�PH�E%h��A�iy�ɰ_o*�I�4��S����!��D@�en. �C�1�Icq�J�@u���'s2���x-�i>��	�?O�<	��ܥEYl�H��M�Z<�E�i+\ŲTEk��d�Oj�d��ze%�擪%FznmC��M�MGz�R���M��JS3��D�O*���1O~��W�8}F(�v��zO&	�T��)5$ml�ß����*d�����|2��?q��y_�,j�
�;}k�� ��
;�	����ɰ@�Nb�D���0�ɼ/^�I� �,�����.����#�4�?�֫
R�����'�S�Ln��]���z�Ǎ�q��
�K��M���=����<����?����D�N��9q�E�"Ih�M{e�ۄi��J��ES�����	˟l�'�r�'qH�	���*U����0�P1dT,��'���'�BU�(i�mD*��4��1\@p�s��^a2 �������OB�D�O^��?��Y���O��-j��̤@�N�3O�D�n�Y�Or��Ot��<�@Ɠ	��O�ژV�2R�*�u�әZ�ޘ`6�gӊ�d>�D�<��s�'���K���5��&�ӖFČ�lZꟜ�Izy�&�G��0����k�G�+"���A8ig~�wD��G�&P�L�����I�2���4�s�� �q���J5 ��qF��Z� �i7�&A����޴%���h������<T�U ǯ�+GdB��e�Y���'�ҁP
5"�)b�g�	�kk.�
�fީO/b�d-	<R�6-��u ��o�ޟ\�Iԟ�����|ri܅��u"G
Ʀ�2�~h���??@��ٟ��I�?c�\�I�}$�ՋD
�^(����.r�P��۴�?)���?��Y�v�����'	"*��;�8�S�պ9-�X{b͛���?y��F���<���?��'�ڡK�&�j��h1�Zut�Pش�?���З���O��$�O��ܺ
;~&p����8�Q��>y�JF/?{�=�'���'j�I˟�*���{��f��-8H��і�i��t�'���'����O]R�s�j��1e�ac�k&��А�����ԗ'I�М_��IJ�`�X)Ec)W��lK�K�e����'���'9�O��DU2HSj�ie�i)^YQ�ǐk옼+Ђ��U.JT�O��d�Olʓ�?�hR���O��Y`jY�^���I� xѰ��%oݦ���O���?���]�.��$��@AÔ�u����t�^�^d���v���D�<)�;�B��)�|�d�O<����'��	H�oʃyS�x`,S�?����>��[r2��ώA�S�T%�-"����dV6ũ �����D�O2����O��$�O�$�J�Ӻ� T�c�� |��ː)Y*a�#P��I�b��5y��<�)��3
6Mr2(�)m1���Q�'��7���IO��$�O���O����<�'�?!��C6!]\|9��B����s���:��(کآ�s�y��)�O
tRGFO�����"Xy���%�æY�	؟4�����`�����'��O��F��s9�J��~��@Zwe�n̓M��u����t�'��O(��t`�(+C�ub��*��p�r�i�b��"P�՟x��� �=�eج�� �R��i6]+U$B[}"J)n�����O����OZ��?�n3n�Ti�B�Т]A�H�G+V�5k.Od���O���;��۟x��薍I��l���p�����Á�u��%c��7?��?y/O��č0 ���Rע1�����W8hp�"L�Q�7��O�$�O|�`�I�2�����Nk�pa�DJ����]���8a%^����ş��'�a�;V�S�@"��R�<����Dߕ����5�M#����'%�N��E����O<����2&��!Q��@�4�Ȥ�Ʀ-�Iry��'Ɋ ��]>9�'i��L��S���@)ȵ�(��&X�R���<i��x��u'�:@_���)���T�`����$�O4Ha��O��$�O��D���Ӻ����uQ�	¨}N�{%�Tx}�^�`Q �/�S��>Y�=�WnbqF��Ge��s�7��J�z���O�ʓ�b-O��O�3�㍶�f �����2lQ`�l�q}����O1��$�6$j�MS1��)\'l��6-E�R��n�����'A ��V���͟��	\?!�k�"3�"5#�M �8����MD1O�]�-�]�S˟��IS?Qr���Jp�FP��(;�J����I�(r�L�'3��',2���E�.mZ��&T���(2F�`�I��R]Y 9?!���?+O��dP1	"p�� �+�h�����m%p�0 �<���?����'X��Ͷ��4�5	H�RK���3�5V�� d������O��Į<Q��m#��Oc�� C�:D��cL��)�۴�?a���?��'����W�'�M��C-"$T0Q3�b�3�U]}R�'@RX�|��� j��O�¡V
|�pL)R+�/2�(��P�Q�6M�OJ㟌���n�dYW�=�d/h`5`�@���S�� ��F�'5�ݟ�з#�W���'��ONШ���V�K�(�᪂??@���=��ϟ,���G�%��b��}�Z� h��i��G\2�R �'j�g��>���'$��'���[���Ky��D6A��X0��\�B�tꓷ?�v�F�y���<�~�U7Р#'�Yb��袀��Ǧ��F՟<��ן��I�?�����'<�bt�X
	�F�y��=I��aӆ5:G��E�1O>���
b��`��(W��ܴ��6v)�|��4�?����?�ˊ��4���$�O<�ɴi���@!��)�`�h���*��`�y��*�~���O����mJ� 
���y%�G�m6��OR1x�C�<!��?A���'p�kӬǚN�P FK� eҝҨOL"1�G�%��I�H�I^yb�'���*����:#f�'u5ʁS)/B��Iޟ��	����?���<��h���U�no��kgC�p�F�y҅�=D��H�'���'��	����7j�S��IŖ�j�04'��<"�KA�	ۦ��	쟀�I@���?� "� X���m��"	Dͺ�m�_>xa���n��?	�����O���«|R�'��h��H�6t~6�ڠ�ZhcLd�ݴ�?Y���'�Ȍ��\�����hօ��"%�w���`�H1o���'l�$R�[��柼���?=k��̊��gB�-�=CR�α��'�B�2�̅��y���A�i\�p4��a�� 4��Gp}��'��$�'sP����@yZwF�P@@]+=�`��ٵB�HS�OX�$��W�P�a����I*&&� ;��V��3��&x���f�`���'{"�'�T[��S���1QH�K$�aQw�o)��6	�/�Mk��N�S�`�<E��'.5BD͇
QpT�Ά3gyL�a�jӈ��O��$۞\;���|r��?��'Hl ��H/r3�A3�ɽ�`�t+9扼6,� K|���?��'a��a�H9B�P�6�����4�?A�,Z����O\�$�O����;Q�����\�4�j�	gH�>�Q�+�Y�'���'��� [rD@3GF��[�]!uI�䳕���vGp�'���'���D�O<2��G�`���g�]�1-	:!٦M�������ԟ�'5�@�iH�iץ.����%q���c���&zțF�'�2�'��O��	
W�� ��iW����\�w�b{�CT�7E�� �O��d�O&ʓ�?i!�,���O�L6GߓV�㓊�\zƱyq(JΦm��N��?)g�Ů��&��P��[�(�S� K1]Tr��S!c���İ<���P�Ȭ )��$�O��)F�]E��c��H�Ƣ�'I>v��>!�7�f�����p�S��!��|;v���dɣu�p|��N����O�}Y���O��d�Op�D����Ӻ#�/�2�쑪���3}xrU�O}r�'��`�/L����O��uiӏ-&,vu�i�H�"��4����i�B�'�B�O�����L]n��0���<.����Ҝ}��$mZn2\#<q����'�H�K#hF��V�%.� �F!��Af�R���O��$������'��	���S�? ©G�x:$TX��0����i�_�T��@f��?���?G�٬ǆx;�G�"/Aޙ �� ���'OX�QdJ�>�(O\���<�����h��|a��E[�:�H�}����y��'���'o��'��Ɏd�䐀T�d�����0<D|I`j���D�<�����d�O��D�O�d%,ܡ
pR<���V]��E)�b۵�1O����O���<�H����J4'̺�H8>�9 $��0ěS�t��dy�'���'��D
�'6N41�o��T�v�� �>�@ [Emx����OX�d�O�˓Lj��7Y?u�I�A��̺tN�b����
Vz���4�?Y-OV���O���D��[?1�㘨	�&����
>����¦��I͟\�'�����"�~����?���k�6��$�y_��2��m�.O���O6�����IXyRݟVt���Y0��Pp*?�bR�i���{�V�R޴�?����?��'#��i��A�L��dXIU��P�XREzӚ���O���d<Ox��?1���U?t�xE�G
���@ɵ�V�Mc�cR�/����'X��'��t*�>�*O����'J�'��T�]0�
)R����U�Bl��'�H����;U>X�B�ۥa���k�ɧL��ݛ�iz��',�0{�$����O���2'��80$NI|7&�b��=��6�6�䄖2K�?9�������-0w�����wL�=C���WN�A��4�?��cϰ��v�'&2�'yrb�~��'\b\R���)rT���'vR�O6I��;O���O����O���<�	�2�0JOR���<��d�0z%���S�L�'��\�H�I֟PΓ]~�}�B����~]`�mB;w�aQ� u�h�'���'^�U��;�����EL�pm��'�2}d����M�.OR�Ĳ<����?A��-���n᚝#�4b$�x%	у���U�ia��'�2�'��	']�p���~��Ɛ�sg�L�S'�I�4�	�i�zu�w�i�B[�H����8�ɑ)Z�Iu��<`	�!�`��F^��+@���AG�&�'T�X�ȳ,
����O�D���%��(Ggr�I����'r&��Ћ�u}b�'�"�'�RQ��'��'7��2pڬQ9�Q"�lջQ�3>��^�����=�M����?1���zP_����ZM(p �!�Xs��	�:7�O�dœ`��>� �S5G���Qd!�F	D(XGMS�P�(7M+)��ioZȟp�	��H�S�����<��'^Nk��J�-��?��(҅�yB�'��N���?�ॏ&p���ш�	U�!�kC�L���'9��'�а��>�)O��D���#��O�r48����
�S�6�Oj�Kbr��S�T�'���'k��Y2ɑ�-{��A����囕T�&�'S@IW��>	)Od�Ĩ<��{`�D�q���Y��R�V!�@Y���T}�K��yB�'.��'�2�'E�I���e`(0��˶@�#X d��۷��$�<�����O�$�O��e�X+yH��!_�^ä��SHL��������Iӟ��Iiy��B�,�5
,Zp�N-lHaR���
�Z7��<i����O����O�t�2OkV�>5Xf`�?K�&8C@�&/��V�'���'��U�t��˟�����Ok,�	��]Z�N�It���b���)��6�'��	՟H��؟t��+g�@�O�%k4���s���p�kƕ!2���"�i�b�'o�ɉQ�����D�O��ӴL~�ċ��ڥC���@�lP4p�'���'ҁ��y"�|�џ6�+vn�@��)z׌Sl���
 �i��'�h޴�?a��?���|��i�UP�#�������?=�T`�t�r�$�Ol�Yb7O\���y��	B��X�8ք�Qz� a�
6E��Ĉ?d�6M�OV�d�O���SS}R�`xgAʟ?��X�$n(l����/�M['�<�K>��t�'6�TRU�B�X�0�J��R�w�r-���n���D�O�������'��	���������`׭	S����N���QnZ�'���ٟ��i�O����O�q��7�ы���4N�]�AȦ��	�Ʋ���O
ʓ�?i)O���8���N_N��˃-A�w�}E�iI���y��'���'��'(剗&�@p�ݩojfxaf�I8��-PP���Ī<Q�����O��d�O���*§xnD�gh��0!��NY��D�O"���OF���OV�@Ԅ��d4���&�E /�6L��:.^�+7�xb�'e�'_r�'�.���'�d��sĖ�Q�`�9W(߂ h$8��>)���?�����)���'>���n��(	�6rT� K"�8�Mk�����?a�B*A�>9�脍$�+ �.2D�j�a��ʟt�'vLA��&���O��醍V~Z�i�m��b��Ÿvn�\&����˟���˟�&���'op������\�Ҝq����ml�PyB)�C�6��F���'��K/?1�ŝ6P�*jǖW���;Aj ٦��Iʟh¤��$���}��&�`�@A�ã�io� 4Cͦ�fꒄ�M{���?1��R�x2�'��<����J{�i��3l���2�M;��<yM>i*�V˓�?�p��,�rdr�CE�R�u:�#yٛ��'��'��	k�@;����l�"���Ŋ�0x�h!�F����>	֫|��?Q���?�2�Ɍ�V�G�`N��r�b����'�����)��O��$%����0� K1b	�e!�c�Q��\�q]��xdŏq�IƟ��	����'�b}�c��%0$q��c;�(�pcZ=?N�b�@��W���D��ǀ Vl�p!ȑ��R)�t�fuSQ+P�<!(OX�$�O������M��|�S�T' `�'MΞ	�7�TB}"�'B�|2�'�H��yB�s�0s�L��E�}�b��;0	�OH���O��d�<ѥ�נ[\�O�\�b����3�-	$	R<Z*`�"�$#�$�O �$Q�Aټ�d!}�՛=۠�3�36�9�D��M����?q.Od����^�۟(�ӟ=����A[��Yk�(+z��J<����?���^���'k�	T�hz� �4+�:�}��Kh�]����̓��MK�V?Y���?���OD�)G�@�	��v<�~�K��?��`�������OӪ�#�[�$�ҷ)�#M\rEi�4g�pu�i���'S��O�:O���=���ƁV�cL�-�
֤jŴ�l�˴��I�Ė��*��_�$�4y�dl=3�"F<M���l����	��d�c�����h���'���U�pH���f�.e���s��U��Oxa��d�O���O����G���0%��d#� R��A}��A�(k�	zy��'{�'?j��4��`b�IՁ�>`�
9pű>	�/q���'�2�'��X�#�_�	��X�e�0P�2�;����.���C�O����Ot���Of��
�Ƿh��u��IH7H����ri	 +$@'����ԟ��	��p��6���I�h�J�""E�+v�"XD����h	aڴ����O�O\���Oe���,ڛ�˯S��|ru�W%lKls׬(����On���OB���O�P����O����Ov�zSf�ɀ�ֱF�pY�M���d�Iڟ���.B-�!G �$��I*�,�7eP�>�bu���ԛ�'��W��c�Ϟ����O$���f��'��~����!�%7۪Uz�����?qRl�"��'��\c���!�`Ͳx���S���F�ZQ�ie��'������'�'�b�O��i��2��
l��!"C����/yӄ���O��z7�C�<1O�����M+f�d(��A�ibr����'�R�'5"�Oo��4��n�\Q�!G-{Ŵ���Ɉ1l��6�F�8�S�������r%A\8�J�ʅ�'�0�r�V��M���?��"K��Je���Or�I,��$��	 J8p _(oc���+0��ݟ���ӟ��ȇ�u�$�˱f�'�¤�C�_1�M��Y��h1S�xr�'�R�|Zc��)�#�0a�mqP��l�F] �O
�R���O����O&�)M��r )�#+�D�p rr�	�I({��'?�'��'>�'��80����Q� r�k��0ܐK����'N��'�R�'��H*D��	�� c2U�E%Ǜq�2]z�h�(���'�"�'��'�2�'4��:�O�E�`鏭b٢����/>;�P��:��K)u�N� cn��<��e�g�+���4+v�W4ct��thR�7��C"O��b�[8jJ�p��d�
]
��O�@c���@X� ��hiw, �Ӭ�>2Rh�D�p�n��E '�X��;f�I2O;m��P�c�0Dn ���9i��@2��85O>�"'�%*@�s�I!Y�t032f�&h"���b�H�(l�5�G�-c	��ˍ �����RDĀ4��%� |B(���ų(�HC��'sR�'��H �c�2SȔ��;P�N}�ǝ@J����nQ=���S����'���gMT{NTW��I�@D3�A�O�d�ж��)GJ$�S��?)�L�6��6�s9�wfћr���G������ڴb����"|��WL��4��o����s�@��̇��5.v�iW/ƅr��pA��1#<���i>]�ɀ{;ލ`4�V4
�(�!�,Db:a��ٟl2P�XY7B$�	ʟ����!YwX��'u(�f��a�1��)[�% �	+�a�O�ܹ�G��]�~�1�Ө����$��*ot��S*0ehep����Н�?yq!��l��@�����3ړUN�ҍ��JC�Q�����D��|�m�d���˟�F{�[�t���M#�Z2,!��q���%D�4p�Ԍ8"��uf:~ԝB�	���HO��Ny�\7mD	��KabN�5���2���ef���O����Oh���@�O:��d>�K���6)-���?2T�A��G"}4�цL�@��t����Dx����k܁w�Z�2
54��Ё7�C%e�p|�!�AZHj�"PO�Dx�`�!��O���Y\6��@�.~��m B���-:(�=���3U24����0f����^�;!�$̧v��sw"H�t(��Lƚ;��@}�Y�lB�
���O
ʧ1�ม ۟d��k��άGc$@fN�?����?�4�9U��a@��^�.�����i��L4�X�̇�R��4�4�˙�(O ��#�t��+f�,4�' 9&:Ţ#��R�`=ză�3Xt�Ѣ�(O�,#�'����Ł+��hl^*'n�ԲC���I���Q���
3a�_d�C �Ⱥ\�6�3p
=�O(%� ���Q)Z��U�WK�zt���y�P@�J�����O�˧:�da)���?��^���դ��,kv|�"�>j$U�`�4k"ع�`õ��E���	+��O���k�b�NL�A"܇!��4��	�TZ�I
l�yQ��
@�:@�Pl%���q���I8�=���¦KK�۲��x����Iߟ���'��h�V�	�hJ�|h��@lH�2|x��S�? �4b�%\J�Hd!ߟ~���I�ቭ�HO�8�t���˛�u�l(�F�%T^v���2��¥d�>�	�� ���<�Zw���'��H�5�P�@�􁰍=g+.�R�'֜�k6fZj�R�o;O։�q��^d<�ӔcQ"���%�OXI�p���(x�Yv8��H���emܟ>gJ��E�����=g�r�'TўH�'B�h���M�'�F�;BA)�nu��'�d�2T�%;|ΰ��L�� gX"f�)�S�TV��{"	��MSu�Rи�"����p�P���?���?���b��Px��?��O�`�bu�i�B�A7?�Tk��L����F�L/�p>y�!W��dΰ@��)���פ_ݳ���%A�|b�
'�?9$�i�:H5!�yC�l�2��6������s�"��<	�������'u|���b+�IQZ��
�!���;n�a��)>~1*�0 �̕1Z���I}�Q� ɂB�M����?1*�X���;� �F�K(8X`�J4+8���Oz�DCPOZ�ڒ?�|���-r�n�����
?iRe���Yb�'�F�c�E��h��500�*H.��Kbb�6�������:��J��b�4�?�*�:L�ӎ�6(�!��a-�]H���O �"~Γt-�tåw0eXg*�D�,��	���X�s�����l�i7%�R�� ��+!�i���'	�%xNʀ�	��͓O�f )0&�>���`�L@�Dy�.)�6m?�|Fx�,B�L���sg)�� %���I'yϤԳG�2�)�矼�D�ta��eM�#����B-«_C�Y�	ǟ�*���'���6jͲ��4k��E�8a�౟'���'� � �h �x*b*va���Q�����:~PD���ڂx�(��ߕ>����O:Iɂ�
4B��$�O����O,�;�?!�!��P1��̨G���"a�I.G>P��� 	��e �T����sdU�P���z�(((� Y��FJ�#a�����?𾤁�R F��h�'�*�B�$˚xq����O��ԟ�	�<�'�:MGJ�g��A ���
�����';�y��<��A�I�4��B#�瀅	���dͤXf������Pu#��?��i8��4ܚ����?����?I�b�-�?A�����4I6ܻ��i�м@���cm<�p�UR�����vO�=�횫�M��B$oj�	1���MnVU���{8��QU��O`�lڷg.�F+��QḆ�a`���� �4�?1(OL�� �)��M�M�@es���x8X+��j�<I�	���Q��Ȕ"�Bآ��<A�Q��'`�A"Oc�R���O2�'j[�$j� �5���@���`z��!�V��?1���?����z����D���ݮu�І�<_�S�\����@ 6����>zv:�<��^͢#��$���gQ6f�(i�O��di5`�� �#wY�@����$��Qs�%m�T	n͟�OL�0JAdΜt�� �3M�,	��'i�O?��i��)��aI�Z*���E%'cP���O�I�sf�LX���(-�4���E�=�2�I:�D��RN���L��H��4!���t�I����1a���R�����f�&ų�B�"F��(�)�3Z1�hQ��&:��i+���0т��5�rxy㕙%��4<���s��uVz�����2=,L۰/�<-����EE�*�*���)!J,wި���:e1l)�猒A��qDx���'�j�s�G�qu�cI�)��%s�'05	�$6I�áN+��b����F�����'�l�6fF��`�v�BG^0��'BrO�cO a"��'�2�'��"l����� c��׎����]�=i�,:S㥟��O=�Zx���&�ȓפ� wV�t.�OA���/?X���n|؞X�6Wt�3�O�Ƅ ��V���$�=3�t�'�r^�x��I�LZ8�)�*�~\��%�+D����J�0X�4y�IX7Ű�H�Ȓ�HOT�'�򄝆+Yx}o�%N����9y�e0"��V��<�	���Ip�����I�|" aU<B���4le�)��CւW���
�Q*t`����*}���0
����5���v���Q� U*�:�OP���'
n7m�B��`�Qhӳ1�J\9UF=cƵmߟ<�':��?��Њ��>���dF��ER�JbO$D��94�i�H��!Ϛ,#����a��j�O�˓����R���	}���H�!�y������A�$�jb�'#��'��˳���7�b��?0���T>mhq�!��a(WQ�`�e�=�x� �iX��(�7+L�3atX��c���離&`v��3�W��2M���H��Q�8Ѐ,�O��m���O�`t���>e��T�K!vl���'��'��a����g+��AD�N�qz���-���� ځȓ%�7M��u�$���}118O�m��o���	��O#6eH��'���'�<tr��>FD�A�+@_��#�	�w���y�b�b�0�ņ֐�������Ͽr#Ͽ'5!�EEn�%��M?]����iDW��� �Q��������X0q��4�Ͽ+�S>���ںx�(Z��D�2���s���?Y�O�$��O��ð�F2h�`����Eh��9O|�$(�O�Ұ@�0.�W�H8&�	��HO˧}.My򧜓vJ�@��D\	dtR��?�GI�&�*���?y��?�Ĵ��d�O�|h�,	e!<Mz���?yl�3��O��O_�$�,�@�'|:1���K hKU�AjW�}X�x�'܈*!n�B�hR	��:���$$̥ ��@F�REZ��H:��I��~��Y�L�	by^#z��=c!�c;(�b& /�y�iR�+P�l`��-]4���6���3`�"=),���O�N̲���ã��2�ЊU�W�u!�$,�JaY�D�/��Y�ċ�'��Ј�ݭz����@�L>�	�'r�ՠ�d�'�$Cv�,HX����'9�[��ۻ7tҴ��A¦�r�'t�R�Gٿ'�����ɪ��L��'�HL�#��X�R�8c�_yZT%"�'��,豧L�p�4$S�b@z��#�'˪��u���!�s3.@�EM�9�'@ͻ�Cǃ{�j�s�W��HE��'�2�h�*z��r��	_��i"�'y�*Ǭq+��
��^z"I�'eL4ä�yy�L�ыТV�����'$�4(%�L2�)�F��i;�'@ް�g!H�~'
��9<6���'ʰP)�$���,�'��/�Ƹ��'ib�ˡO��v\ 7���/Ɗ���'f�=5jSpK
���V#��L��'���X�+$$ykF�0��d��':F�ir�S�$�H(%�ʏ�de�
�'���a N�:7�����"� R��
�'�<p��IŜp���;�
��B�ډ
�'}�P`Q�1����'� 8��	�'��pz�OYP��7��,ZN %��'��b�U>5�6�E�Pr}c�'T�!贩��@H��3V��Nш�'�b)��V��E� Jb��'��P�Ǎ�@���a�ȭy�p���'��:lˊ&�(	�1k@
�,R�'�YeZ�Q>�A�ں�H!��'�Be����LA$�À��qO��h�'sL��CC�+)v�0�>
yR�'R����L�;H��w�3/����'�֝!��۲U�4���oOK��*�'쌡��a$k9�D�1���K��	�'g�u�e�1o�=
6���mR\$v�C����*�� �"�E�@�6�~*4o�$W��ݛ-ʺ�b6�E3u�T=��Cɯ�B�ɻmJ:������h[�Aa��	�wi�ۯx��ic�X�r��E�G�p�
��b�"l���D>_T�6`�%g��b4g BKax"�ʔaˬ88b`�y�`YD.�a�|Q���A*
hʜ�EH1}<�A�5Y����܉>��{B˾;6MJIH45�ҝ˕i����(꺄x'�N xA��lߖ	��B�392,�������rR@<�"咱��;��  �"O�!�!�1+�yr+�:NiQ� �*f�BZ�n��c?�mࣰi�$XG(Sj��g=A/���wl�B"�/Sv\A	U� 5�TA
�'�l�@E��58L�����-���6H�(�?�A@�('ΘӴ��-ԭ����\���u�d�+d�y:s�S&%�p!`���Maxr�é[U��S�3?���k��*v�����oK5l6$�!DI�X�$�y"�ܭyu�u��nSZ��{���5�f$1�GPT����4��(��䟀@h*�eQ-5��pA��®`��)H"I�2��A.�"mԍR�%@����I�����*�"O �1JL�����Ɋp���x��|cD�i��A�{�(A���3&!�5B�|�&�P�޹λj.�b����*���c�5+�����x��R�^{�X{����+lCD���ڿ��GT
�݃GK]9x(��S�ӎ9��d�$��<<Ĥ��x�:�D]����K\
=p� "��T� -�n��F��:oTɻv)���O����N)4꬀�J��W���ԫ��^�KQĝF��Tp�&�
k��h�Q��P�@�k�@�O2������Z����~ʟ�y�f!'@���jM�L��r&���;�"�>kX�� �@NO�e�� ��%����FNd$�ӭi�bZF��M:N��GB�W�^ݘ�'ց%�X�ڠ딿8���s�D�R�עE��=K����<z��dI$JU�,Y2#ƃT�.� �Q��c�|ҖO?}����u�uI�
8V���`G �y2�KD���
OfpF}� ��Xb`��I>'�2F�\�B$���M��!��\TQ2b���R�J��>ͧ!�-���i�|`#4��(ZPi��6y�0Q#�V�'��i��M�6=�`��b�k�@pg��S7
�(���Z�\��"<i����lá�O�)̧ �esn�>@���3���<6`�	p��J����9��U�`۵"�����0�%��8��O6����G�4�����d�� q�'�I1�J��$	�[��b�D�����g>}r'����G�V�
	�U:#�¡i��+1���b�}Z�O���B(��y���) ����R��O4 �6c�+�ܼ FCO��O���j��?V !{�J��zY�i顉��
��Su���'V�:T[��i�N����@��>�[#-Κu���p��H�'��)�ÞuR�[�񧿫THW�t^��筙^����e�'p
�ϓF����s�Ox`�I�!��Бd��w��鷧�|�p���n� ��$y��r���"� 3��|}���=y��%�T��H�(�NY
$j�YIz�IH����'����2O�*ap E�2',I���vh_ g:����_�Xd� V:/�批N���&�p��/-�l��׼\o���RCYZfe�+�p̉q�H9k�0e��m&O�-@�h��(�ޜ�E��S!*���"$�ى��ݩT�	F�O� 5��fp��:sBϪgޱ�P�R����fb��s��~�;}R(�q	�ML��jǚh+P0L<!/ĮuQ�D[+>�g?Y���i�|�jφ�\<��#H7;�l Yp�YH�:�ꑄ]����cآ+LB��cK�
U�F|cq�	(8XQP������5?���I<Q����/�n9�JJ��'[�5�͂9#���%�����J����C�+t�@T��m�>�X2�h4�	>GSv�#�i��3hjhF��X�l�B�:���6 �,1�!�'�����#�����D�yشS���p���3!�}І��o�P,���<�$.�	YWʤ���G�
L�z�R>
b"B�I�D����ɝ�$,�d#�G^�m��I "H ��?��'��$�K��5U��;�*��I���\'ga}��ۙ��ᣢBO�pW�h{%H�/J�T��b�y�������:a�u��B�0yޔy���5}���P^��"�vqx�j�K��hO�%@c$�7E㰄��M< Z�Ђ�O8�(	/b�e�+i�t�8����p�1�)֐I�ƽ��A�hX��y��*9b@d�2�J4*��M/?ɰm��N�hUr���uO��C!Oh�T>�Y�f�K9l5j�Nɣl��Cc,D���eY"���#��,L��|�p�V�hٖ�#v��+x�x�䧘Oش���Nͼ��	]Ė,r��Yn�����[J�<&�(%V���+�"0��NN!�P�-O����@�y�1�1O&E� `L%|�F���A�r�
��mR�M��U�CdD+���"#�_?M���,h���sL�1<�^|"�)[b\Hˆ�~G$��	S"�j���"2�\����H5E*a�5-��V��, ��9�U�T�"�&����,Ox�	���	UW\�x'Q�#�kS�'	�\e�H�J<��W#Z�RZ��p`��=��a`�G����'��A 47O�t)��;J����&����W�'픰��G�e��z��,Ą������p��(c���PK<���$F�m���~��s�%$@�L��E��<%���G�A @h�4|�D8��J�?>���E{��2LHl	���L
��� A�i��!"G�մ��� �
x�e��'�Hm���+�����O������0�1h1�׫c;�h��+��&�,�/�OJ�C�A�xn��W�3>��s �T����:l�d��C8�ɭ|
��qp睫R�`�7O�
𼋵f��:���M�u�4 P�D�Dҩ[�Bڧ:��a{���:|
�y� +��a��H�Po�,϶0Y�G�/�d�7�Q̱;�(�"_AL�Y‏8?@�"<��2|'��#�@�A���0���<��*��&oT4�L�g�;V�|X�L�O�=Hs�'x�ћ�읪܀�a�dJ�HN��2(2�l�iA�H�D˦����)2 ����̎�I�4O��6 Hsl�kE�O'!�u!� X���)d;�aے'�;_�R@Zj���@��'�"#�<�P:��˺
K�����yr��g3���0����~bLI~�����`�0� D�Q%�|��s',?�O���2��9eqP:�d�	j6�Q6A1�^���T'�&����O������^���DQT&���ˆ8�����j܎Q�<eK�(Z>{s�D�cg�/u ��	��ĚY+xȒ`a���O�-B�-	y�Dri�:a��8��E�O�m��� :.YIʷ,�|�#�V�V��%�$��J�@��3�e�+�� ��JY+2�4	���<�R��X��%��ZQ?�4GV%� ��Ӏx�Ĉ�9elAq`hELBX�;4�'X�W�t�'dA��,T�:�F$�vɏ
�<��I��y2jU0)��x���ہ�~�_}�'��@p �M=�4�K�)B�Z����$G�y�! &\J��"�&À D<�C�#v�������Y�pE�y��Y�p����'�(q Dξ?a��G��N�T�áU*\��=b�Aѳ1���R8@��P H�P��;D���cr ڱ%E��!RZƊ����Ǿpx����A:�"���ٙ�h�i�/_L�����<�vL�xJPQ@�F��e�@D�4#�-GT삣%$�tHZ�T���ي�9�
���_�d�'�X�^����x�H�������: �
�?� ��3~BX�a�V�Z�v�a�B_��X8�/��X6l��!e��]�*�ϧ�?�O3|tcKP��a�׆�p|��X�N��*d��a��>��y�F��j��ҝw%�9��%6s�CBگNN�S���\�Ra1�'������d;-��q%4w�A��dƘ� ܪv-ш=bt%���O@��0���<A�Q�J�Q���H 
�|�B�.C(�(�v`�2��5X�� ���p ʛ.�6(�$N�EɈF��P���` �B5��Qc']/�H{A��y��(P��<u��T� ��W.�}��'ʔ��0�ԃ�#��8E(Z1�LY�M#H<z�I�8uz���NJџ c�&�o��XFN̙F�д�Vi�0��f[�%dĝk�I�(K��]z?�O+$s��T�dvn��΄;i����s��;gl�Ke�!jn�xB�ߩ��&e�咀EL�Q.��G��_����(^I�����O��P��� qbi���W�,p����/�i��X��k�Qq��P��;ѱO4U�%�^��
}`��B��Fă�J3��J�5����m��)�B�ծ�4m���Z'���OR6�ؖ&��*Hъ�<Q4䆣3����U�n�9�� �2�n98��	@ZD�2ȏ^��,E��O �Ka'S�%���j�	ְP�À
R�T�2dY��[�6`	�G�L( �?��d��`H���9���s���#/͖	����j̰0����G��<���~��$�p���MzI�T/K$	T��{��]%9i>��C�l4q��爠2�k �(VK@��b�4Iq����B���n�H�G�/p��'ڌ�"�?�� ��9'���Ks�!+^@��t*�AȱO<�@d�?o��xg'ܫ�yu�#�T޶%���5,�`���A��e�lY&��4���D��	�*Cr,��Ot�I'�$�B��-���f$�dgr%rIX�k�z� Ti�:.�r=Br&'�U?���йV�ՙp���ӣ�$����+^����1<<�FR;`k���dI�F��9rV"��oy��Iǀ�9��uh���#�rI�O�0����Ӻ�I	��H�� 1���A(T�D��2ʝ@�UX��U�b���$@�.���3Q�I)@�x���/,y�����6}���I����#��d��'̴��\"E��秘O0������e�k���4<�ڕ�jCV�6%|����%F�� ���Ȕ2R�EhK?ٛ�j�H-���d��3�p9�㗝)/��'��"v��|����V�t{J>au���:�0���WA	 1Xq�,w:��B9�l�S �U����|��O�T��&x!C���lb�x e�?%T��e�4؎�"��' �&�����sU���h5A�#Fxv��g��b�e��� �O�T� n��	��DpMJ�qt��D�
(��-�B�4��f
)��%�:Y�L�*!1�ё�S�6C�������I>��4H�
�?��>���&,�E����#�"�^`I�k��4:~c��X�!��@H@3lZ�0�Iy�-�N��{���1�� )f�EB�(�M���D<�s�@���	���'ڞ��կ� *�dApH�>f���噎}:��C@��eK����ԟd��D�%8����Ї9v��A�
��ɧ~��ʵk�l8������O�TI�p��|q��M�_��� D��H�����<����]}"��=� Y��ɄSw$�3�w��̇�ɉ{���������%kL�;oNV�Tx��
��~Bϑ8�r�'�.�S�s�((����U����S�ǎI�Tj�F9D��+���<Gi�Ea"ǐ�hC�@9'�$D��2����#s�! ����֭"D��J�a _Vn8
'���;�Z�3�H!D�D��́� [�hB�G�&�PTzfI)D����� �|��aÓO�$y���3�H3D�D���W=}��ء�*�m���{�!6D�8H�*�dT�I�B�� d���5D�$���f �i�1�6>"U��B3D��zb-���G$ֽk5D����=D�\1DB�7A��0���֨k��S��8D���p!M %f0%�U!p�$+�+6D�� eD�i���sl"^,
yP�.D��29HB8X�h��
���q��*D�\a�Ȟ�~�"�����L��f�>D��Ö,��h|��b��R������;D�0Ic�Ǖ�@JD�Ҹ\�<����'D�T�2>�Z��+�d�"�ԋ'D�0��@��>�X�!�3 T%P�%D�h�ĕ� �� �eM�[oм�G�=D�`��0h�4��A
2粄J�A;D�� FU&�QZ�\��eɋtW��"�"O�Y���X�y�*ɒ�FҰ�q�T"O|���![�=����6E>~� ""OlD9"E�|8�+�#�p��Փ�"OΡ� ڙH��%�爖3
���#"O���n�*U�ąsM��y���"O�L�uK��.��-�j�d��R�"O�$�n��	�H�l�4�"O��K5n�T����kP���<�"O<�iU*$&��!���F�y.d��c"Ob|S5�������ؠ/#Rl�t"O*!TE�)+}bl� �x��c"O�`��F]�f��c�O�Mt�t��"O�H8qaB�xG �a�?!tl��5"O�tg�	Cl��Q���2Uz�"OZa��!�L��@�ћW�r��d"O$�bs� �����vyZ$�"O4��B�I

��:�EC5�u0d"O���5͜�k.p{�B�[���"OFIٶ�]�V&J�2Q�ֻ�(@h "O�-�@�0��բ�8��#C"O�9�(Dp�
�ip��4YmʀY�"O��h7�u��Ta��ݐ;g�qV"O
��'˪P�$8���Ī&`�� "OX���c�\�~U�	ԥk�ȡ�"O�Xhh���P��ʵ
�t���"O2	��d@�,��BP�I�;� *�"O�Р��̆ � ��c�3/((�T"O�h ��;7~���K�8:�0V"O(,���)#n<����u�'"O�1��A#N����KJ���4"O8�e熞�܉��n�<E���s"O&,"���]N@C���ВE��"O�X$M�?H$���:�3%"O�@��.�Tj��_�J��q��"O�\��A�A�Z�'h��p�d"O0j�	�#+��f(v���K�"O~���mD�\���SA'p�h��V"O�8��-��4�����F�	� с"Op�p� �\ �h``U{n"`�U"OB��ɦs�.TC�ɂ�V����"O���I:rqV�Z`�T�87��ҕ"O.�ɑ��~Ѫq�I,$��%"O�H��H:�| �kP�v^p�"O���Zd�و��t!���E"Ol�s���9
9~h���+i�T�S"O����˖����q�D�U�b�q"O��[pG�7��}���[����"O�E��׶..0�$�D�X���"O����A@Z����4 X�ӊ T�@ ��G�����F��	:f��psB(D�Ȃb�_�U(����`,�*��2D��a�BÄ)�V�b/��ee^]��%D���� U?x����ԍm� �*O�����.]���QR(#�^l��"O�xy4N�B~��!0���x'"O}�ra�e4���`��xV�,�Q"ObIZ��s��t�X�j���@q"OJ�1��F�����ԥiyN��Q"O��Zc�lC���hH�DL�D"O�p꓈�50y�Vǔ�:��s�"O6��3�&TJv��� �"O�q�d��;M�0ՙ�$B+7&|�(�"O�Z�`�?P�B�b �?��� "O� v=������>���� ���{�"O6ȸ� L*�f�Jw-'��@�"O歐�iP;2�h'�:^R��"O4,�!N�mQv�ad�<�X�"O.x�� ,�6�D#��@"O������b����[�.�:�h�"O Pa�Щv<�h�A�;���"O��4�6�`a�����e2b"O��� #�%NuxXYe㐨��la�"O䩢b�]b-\��wO݂D$�Q��"O�p`��J���H��I6L�3�	y��$x�2�y6���W�Y�f9$���0���{�D ��T{�ڶJM�y�E�6����(�
Gֆ�MC-�y�";���I܏M��L�%��6�y�$�=|v%�1BʟKT�`%�G"��',ўb>mcB��j��8BUm(W���� D� � G*��0�K��4���F D�tˣk֭"�����o�gȔ<pwL?D�H��
j���z��|fpRР!D� Q�IB���0����y{8 ��=D��(�b���I@$�Qur�#&<�Ir���'zA"�ᗄ�
�\�3���f��\��y��0g��Q�`��F��i\ ��y	*h;qG�<d�e�Pț�@�ȓaƆ��Eϋ�^aV�*P�"l�|��s��M�gg6NeP�����Nu�i��~�whN%L7*A���DsE��������Q�)M�I�t'�<����H���R���`�A��A�������b}���,hjn����Q<h|%��o��y"�ģ������
�x�B�@���'���ډ�����s̍�#xr�(��O�oE�iv"Op})V &�cr* 6���z�b8�S��y"��_���C��Y��#I�&�yr	��0�\M�%�Ʋ���IB���yb�[h����JJ7#\ɒȏ��?1�'4�ږGC�Y�ސ� o5N�>x�'�Z�Js@�;�b��WkT 7�Z	��'��%2$�\. �廣iJ-EGN\�	�'M�Ab�Eڸ�P0��ʦG�T�q
�'2M2҉�&$Bp���6:C�4��'�(���OG
� QʤE�4��,��'p��&�(Mj~Bs�-,:�T1�'��5��WDm�x�'�S?+���"�'ԑrDJ/ ����V�Ȏxc�;�'٬���-!�v�*���0C���
�'��-�Vn)/��h�E/.}N���'��1Rh[%P�^\�`� =4P����yb�D�K�|�	D���w�8�S�b[���'��{rFڐ�d�,��i�ZQ�@
,�y�H*�D�AJIgY�]���� �y�F�"+�]�fc��Q��ŀ��g�<�͊��0:�X=D��̈b�N�<��&U�L���dƼ�U��h�p�<i�i�&"�����V�{^&�ZG�p�<)f�5m �*���}���[�%h�<�p��p����7Cn��@n@Z�<�a�M���,�} ���4MZn�<Q$�ĜNc@���� `��A�f�<a�V�{�+b�N�fX��A��a�<��/]�N@|Zү12N(�Dn�^�<���F�'L)��Ӱ|[�����@W�<�RX������Y0B��M�dh�i�<� ~�e
�(�:a��Y�}D����"O|�5k�� �\��H��U�}S�"O(h���.�4��F��6պu�"OT0ÔZ�	�@�+�l�l� �"O�x����;n]T�8W��8h���'"O�Qr�@�]&x�P�;� �`"O��:��[����[�I��k��`�"O���E�4��Ti���S��E�"O�x���#_ےu#5oQ�4���"Ox9Ʌ�Mb�����JM$��2�����ɫc�:�����iŤ��3�ED����-��ñ��Q#_��b8�W+B�<L!�$K�j� k�^�(?��PCː
w!�dI^JraQP!�"U& \[ظ~]B�ɻ>,$� �
;��� �'g��C䉛)��is��	 ��Ur$�M.@�C䉴;)�]�A�0)H֩��aF3+!�C�ɓ M��)>^X3�k��9��C�:>h��Ơ�9! 4�"�o�bo�C�	�:�m	X� ��r���`ש#D�Dq�i��ʌ�tO�[l�"�e7D��SS�Kf�ɻ��
+Zb��Ӄi!D�w�:B���S�1Vn��a=D�T��^;a1�e�r'Q2}q�҈&D�`��k�>X�40�a ЄRR:���%D�|�բĔ��i2P���E������/⓷蟊08�JP?EЅ�s�RqF"O����?F�̑Q�I��.�ɶ"O����o��dH����-Z�"O\���ו: Z���@�hձ�"O�h�F�O�c/&d(��t{[���'H�k@
45�D���!�-�H�[
�'V�=S!�>3)�aRuc#T�I��'�.�Y6�$|��X�sJ���i�'Q����*O�.I�����Gh8�'�\�pd/�:8�2��# :�{�';����x�,8YU��Hy0��O�eҲ� V �Yu�L�Q.��"�:\O���SkW�>��K�	վH!B(1"OJ�ZVD[ .�"e�c#ƥ"4|I6"OD�k�nA�.L��hEn�F*OF¢n�,*����M�|�pp0L>����߹a4�R���Dv�@�f�Tf!�D�	��H�ªN"yp�؃I@�"g!�D��-Dx"f�/+�ndـ�<\!��$���]�{�hp���vG!�DC4�A���	{�*��'>6�!��!j�=c�\�f�>]yCa"~�!���H=�ɘ6���"��i�%R�A�!�� RF(�r��<JP�8���h�!���>G�.�i�M^��S���^.!�D��p��Y�����V$�#J�6
!�L�_�0m����y�����&^�!�$�+�`)�A�6m�A��
	�!��L;$�d���I�W��j7� !�D/��m�G��E���<!�$�#4b��H� n�L�N�/.!�D�(v��1*�%$X�a١�R%+p!�D;r��� ��A�c��	��Q�fY!�dP� ^�8��L"R�� ��� pT!�):�m#�F%nǾD���ɑBT!�$%ր�%�Ѕ.6DI�o��V�!�D, �L A!ď8��A�7^�!򤉶_7^�J�ɣ$�Db��7!�� T��C��<I�L�Fo]S0hܐw"O>@;��Q��έ��˴,�-q1"O@hs���|�����%�=@洼q3"O�X ��� ��#����\�)�"O�[��[�"V���
��e��"ON�HU�Y)��THЅ���V��"O�@���6&��:�D����"O�� Đ ���kC�;5<��e"O�ěe��L��A�k�5>� "O�Ƀ��V6(Y�p2� �~0Z�"O�CH��ڹ[���5��A�"O��a��0yy��2��%�d\�"O�5@TlV�MJ	�4�
����"Ol0Y�`˥|{zL���4e��;2"O6�UA@$p���V.Y1O���"OF��2ɘ7,nPl�<3���"Oҙ��J߻цS��J�'}��"O�2�s��1'I�c9��"Op�A�QA+��%ܞ!L>��"Op������I������`�V�y�"O�� �!"M^��R'UɊ�P�"O�	+�U
*�I����![%���G"O
����"VD��Z1Nȿ|�T��"O���p�C& Ѣ!z�m_bl��"O z6-��> ��B�R
)8@��"O8hQU�޹f���;Ao!Q ��0'"O��gk�$w9�-+B�D�欥�G"O,IX��<�h����N�r0"O��#G"ԧ��Űb�T;޸��"O؍��cFj$�ъ��I�ꀓ�"O\A����3S�f����ơ)����"Ox,�UiX � ��֮-%l��"Or���O.���*U¶Em�"O�9H�F�h9F�c P�H�FxY�"O$M� ��	��ur�@���c�"O�0��'źP*�8���8E�,2"O�$�4�̒A�jD[�@������r"O�ر��}n��2E ԍA����"O�}�ޒWe���& V>0��S�"O����K�faT	�j~,���"O`�ĥY�X� ����-OO��"O�h��+R��ft���t�B��"O�u���{��@�7���~���A�"O�l0�ˎ5�Qa@�1jg���b"O� �� �!Զ�S0��)X^=Õ"OvyꉐG.����A.T`�E"O%�q!,K]>���C@�w�.�W"O<P��$�m���Ӣ�U�x�d"O������hb���z�X��"O
!3�'Bh� H�(��a�"O�`�ѕhv�Q ��Z�d��X�"O�X!���`���(�D�#[w��R�"O"�@�.��ݶ��ʺys0�:�"O2Y��#ح�bPyg�D���d��"O��	"��dy0���	~�C"O��Q�q����d�E??p���P"O��#��%gP�<�!"ڸV��!�"O<`#&M�Y*Z�X�+���ԑї"Oج�7�3���ь˖k\�!�"O�!��п[沈)��H8v��"O�d�T��JԸ-h-kaB�[ P;!���ge��Xu��9�8P#ÖE!�D��qpv���\=O�����"�P�!�]��:ġR,o�ĠT�#�!�� �@�`ڬ|'�$Ё��I�n���"O����ޘM!
��0L�>z�Fؙ!"O��g�� '�T�DB�
�
h��"O@���I�O;T��i!Kk��""O�����B�cȄ��Ađ���"O��� ���|���@�.4���"O:�zE̜#�*l�S�F|���"O��	tiO:%�p�cn:�d(�"Ob�����D��U�$AF�b"O��rӌ�b�h���,^mZ�\��"O�`r�63��U��63> ��2"OT��r}3jq�j\�i���c"O�ixtNG���J�Iɣ'��I�f"O�=�F�9_�(1Ί1rz�+�"O�Ѩw�ǩ2Ϣ��NA
0��@g"O�5�3�w�����G����"Oȝː`�|�hĊs��ܘt8"O&uA�%f��x�NJ/RqĬ��"O�\�sMÃ�dB%΋�m���"O��׬�0%A�l�jpF���"O�sr��lc~X�P� EdN�"O=;I�)/,�����,# �Y*"O�(j��O�l�+���	�'��P ֠B�a��!�gD�k�����'��m����B'�����	jX���'*�$X��V�h{ (�7�8\��	�'BZh�Ǆ�!|�"I����[����'�ʹ��` �!:�`v��M�����'Dh$iԎ�^�^�U� �[ ��`�'�f�
�l̑>��U�T!%d]�X��'�v9�(ͯe��0\��!AF��y2BP�"yY��PBV�L�S%�1�y�[�,�*�g�7P�p�9DD�1�y�E���&�t)�Ӟ��Cd��y�PE5��������� ���y
��Ԙ��i����pUL�y��T�x<�����wRz|ՁӅ�y��	e��肓�]�޶�H��_��yBbT�k�,PK����E"�t#�"*�yҩ�d��l�26~��A���y��K&e����k�>4�V�
�E��y�-�
���B�ɀ�)���a��y�Nڣ��E[�S�q����yr�K��	#�E^�����׋��yR֞$��Ó�"h� K.�ybkR;E$ʉ��	�9SZ4`#`ś��y�l�$,U��1�mȍG�3rO���y��Y�	�4*���;
*������y���$Tl�`�D�06��z�B�6�y�Z�r��c�)6qn��4�K��y���/6b�#���Y���sM�y2���jd|��ςIqf9��)?�yR�WW�	�veQ�*��3!�6�y�i�&c�)a$pEXgʕ;�yR�S�	ɫ2B��7I���,�y�E�"�@�JF�4�uk��y���kR!�*̾ 
,�KӉ݉�yr%%T{z-�r� t9�(do�(�y"���
S25���'؂u������*�3b���j&��thH4�8P��3xYbn[0kv:Ѣ�ojh�T��3�hř�L�t| �AAA�B�d��ȓ�tQ��$)�pk�T5:ҝ�ȓ,�XyS��B�8��5)1���S�? �H[�#��,�m�C�T�(��
$"O��)�N�n��X��âH�|��a"O|UY�#�)=5�̒a-ǡrK��� "O��ZwÆ#OJ9[�␇W�db"OР�׎ِ6�0��s��&U
�"O8��C)ۤ��E�a�턘��"O\���NK\�Nak���ky�,��"O*Bq�{�pȢ��5j�!��"Oꉲ֮�#-t`�XZU���P"O�l�0�N(P���K�D�A;̡�e"O�ahe֞�8��%J�p'����"Oaу�<>vL�Eb����"O`�kM�M�
�̍g$� �p"O�	i��ݙi#qҦDC�u0B�h�"Ofy
�N Hy��F.�ry����"O��@�˛\���a���#:P
�"O��3�^G��\@Q,C/+�r��"O&<��υ|�N8Y�k��T��`"O�d�gD��>z��4쀷A���aQ"O�s6�S�
��AZ�4*CNt��"OF�I�+�.S|D��wD$>�W"O����J�\0#Û�"S�)R�"O��b��Јy�lҪ7��L���2D������e���P1a��C��4X'�1D�A@0.�ɊP��b�r���:D��)�$ҞA��$���6f�+g7D�$���T�CĔP*P�K�_J,0	`4D���Ă��c��P�aD�P�$�8'�6D� ��1S6BT8�N�>D�2`n5D��� �B�W� ���$��hqh.D��{G*��1zc�Ҧ�$��T..D�� �)=T~�xC�N�O$�M0D�d8�$��{9~Bf�t�c�a-D�h��ʛ�w������G�Ҭ���5D�0�W�J�n�$���:��rW>D�D����#8L���# �`�C�D=D��L�-Y�� �Q@!G0*\�r�>D�Ћq�&o=>0��ˎ�)�^`pu	=D� �����LI�KN/h��0c��7D���G�q#~�����{��0W7D��q�Թ=ϼ��D�K%t[� 3�c5D�8�QZ�H�ᣡʛC
�t���'D�����7b����͚�	n��`�%D�Dj�'�VH �
ܝ,p�` �k(D��ڐ��B=�Ex���=Nr���h!T��S��,�v�*���}XN堡"O��r�`��N�Z6MHN�cc"O�hH�(��LQ�F�Q��"O��E	�?���
D�	
/6x$h�"Ot3�+�i2�qK�N�1 (���"O�xɒF����#m��F���G"O()��l"���W�\�U��"O\�W捰�s�*��講�"O$|��ab�<���1���%"O��;r+^~�D�bX1q�v83s"O Y�qo�H��p# ��"O���`*R+c,F$���K+=^a[�"O���f�"M����I,�i��"OP,���W�l)��� �]�xb�jF"O��ҥdʽKX��b�4o���b�"O�ꖅ˷"S�i�0��K���;f"OM*��*1D�#�!J�q*1B�"O�"E�=���c�*�/�iC"O�c� �9���P7bfuy"O� xm�R�ϽN�!��#��e>@u"O��sEьMܤԨR>I(��"O1����0"d'���"O�UqnW�x����6sF\3�"O�Ti'�%L��{C�7c��l1"O�a )D�_m.<pGÇfʹ�1�"OT5�
�	FA(2h�M!�AW"O�8�-Eb��uJ���g!�9�yR (O~(C�_z	�)?A ��Y�pp肎]�d�Ӈ�'�q�ȓHXL�3c �<T��k!��:M����ȓ(���J��t`��  /�Ф�ȓ,�=aƏ��J�q��=�bp�ȓhti0��L9�ڄh`�@NV0��j���8e��&i�������:)�I�ȓQs*$	�i��jn��,�
6nN���9��)��R�*L�q ���1��e��9����2'�H�L�y�`�k0��>��XH��{Vj+U��6�h�ȓ`�`$��_va#gL�<��ȓd��y@BC�XM��r�~���en4����[|�����id��g$<��#�'B�h0A٬ ���ȓZuD)ذCZ�غl�ƥ#Z��ȓ]�1[sDW�jC��)$C�si��ȓHW��n�0��5��-+xE���ȓb�2��Z�6I�󮑪0\⠆ȓ{��=�$ڞ`c���j�%^��0��^Z�jD �j�T�Ɯl���ȓ"�Aiɠpq:��R�%��q�ȓ�������`�T��� &��ȓP*i��/<&��w��$c+8D���FѺ
y��P��F٨���'D����g�%����ϓ�#v%�s)$D� �be �+R"��e�V0^E8�(D��BPC� 	��|�7��\Q� k9D�(;G@�f읻�'X�Gx@]C7�8D�P��7q����&.B>L�t��e*D�����@SHn�a_�N�~Isub#D�
�ǟ+g]l%P2�GL���D"D��e��;*�L|��+�}6K#H D�� ��T6-u�htQ��3�2B�	%3�a�a2[$�X&���j�hB�	���rV���Z���`tKA�2zDB�I�j��E��q܌+���s B�	��x�j�N�C��hU�U%C��C�/HV�P0j�6c�PÂ�7w�C�	-6��!f�WrR&�"�gM1i�C�	� ��i��MuZP��Ǌ�Rr!�䕯F��p�g�5)>`XÁ�K5F	!��*j`6��wΒ��´;6�Y>!��
�	Wʽ#��N;[�d���J�d�!�ی�#�M��D\�'�I�!��n~������q��p��!G�!�LRα�vG�/�ȍ�w�^�#x!�dT�j|23+±#�m��EE#a!�Ę�?��ت� ��Z�C2�� 4!�$'+����eJջy�n�`DR�!�#
$�=P�Cة ��@��+T�!�(TNp�نG��=�Iw �2v!�D�?e�-�E�^!$��%�ńʢn!�K2�4�0�פ/��$K�D�MW!�d�ZWLI����+\�c��&et!�L1�>��̮<��4���*a!�� ܠ[qi�M$x뉵6���"Or|��C�UU(9�R�Q(HPIU"Or�i�-H��ٵ�^�D�����"O���W��x�z�E!�(��p"O���b,�R������ݠ "O�u��O�%@��J��,b��}�"Oj��w��;l|ށA�mC&�x5"@"O��0}H�\��� pu��"O ۇ�1yz����Pm�H��%"O������mi�<;�!*�|�R�"O�``/ɇy���C&`��-v@9:�"O>x����,�%z�n��Hp蘀""O�ʖ��vh#��cP,�f"O��r��(T*�sg�M�b�qh�"O���gH�1n`az�C�2G�R| �"O.h`�@J�*�XAl� 4���'"OЈÒk �%�Z��e�P�xf��	%"O&�J�+B$Lk��	�hd>��!"O����F�#�j�P5*[=f�`C"Ol4�P+=<^��Qd�"}�^U��"O��z��,s�4��"\�z�8R�"Omk�7�TuA��4A��	Bq"O�ٙ��R�|������O[>1�"O��@�K �l )T@�6=2Ԕ+�"O��ƭ��S�<�Q'&D=Bb�"O(�0G6zE�X�� eJ!��"OB�tz�LDQk �Ax�� �"O��X"�J�%4�U��*�kaE �"O�|�p��s�Ω�I1Q�	�"O�1���Yh�H��j3��*w"O������U"@�X���h.�=z"O��Ȥ� 29��y�M���"O�{�@Z d�x��ƤA��"B"Ot� &��z��#�AB�#0~d�"O�P�ui[@��6��3��D��"O2 P!��Q�՘��?`�8�c"O��K6�Y_ր=+��+~��]�P"Ot����ҰC�W'�@T4�D"O<e*TD�X�t�%�#�eX�"O@���LM�j��ݠ!�4�"O��H�/���;� �>�B:�"O �����2-QP�O c@L�#�"O5�f䕑C��A1A�W$���p"Oh\��L�e�l�L�(��+$"OH1�6`����r,ċ-1^��C"O��#���(/����g,�r>�Be"O��	��K4*���ؔ+!e���#"OZp���%�nP�Q*�*j��B"O�9���p,�%�Z�p�2��"O�����gH���A��
@(�"O�9���H�V0g��
�`��"Ol���HA�Dd����U:#�́��"O��)��/+����[f��e� "O,m	H��6��x!�"^�{�����"O,DB�C�0B���RH�!'}�"OJ�a�J�u	:2$��?�%�"O�I���<��J�]�6��"O��'mM#BT� 2���8���p@"O4ɠ�6�*qq �҂G��T�4"O���$@ &7V��h�+%��"O�]���j�I2�'ӕ\$xy�"OtHx2��;l��s)&�,xG"O��R���↺t2�p5,��y��hB��Ȓq�LA�D ҄�y
� D(
��R�U��@���J>(���p"O||�	۬M��!
W>�)��"OZ������b%I���/ ���"O�\���	�8�&\:�Jǜ �ه"O� �V��(h64ԀE��FwP�"O��
#��\�⸻��#A2`zf"Oa�F��+�Y��J4X\
L�"O̽rІ��-~Ԉ��B�'U�]QC"O t����#	�TH`���T=�q�"Ol��#+X�vgnx�u�́5C���"O���"C-���Շ��|B�"Oeb�bԼc�#�ʓ%��Ke"OD$ v�R�Q��:�-ˍTTA0"Oz��&�r���cf�Z([V��@"Oe,��EJt�1��Z�lX�Hc"O����L�Q?聴f��t?|<�d"O��	�*+�=��F�{<l\B�"OT��	���P0z%��D��1"O�|�v�D�b��	���9;�Qۅ"OjeѲ��p���k�#V�L'	Ya"O
\��%T�%���P�L�'LL�"O�9A"Ì�1N�C�t�d��"O��Em½;������I��R�"O�p��L�3'�)7 ���"O���`�&��d�& Y;4B<Ҧ"O�ȓ�ψ-#�N�Ғ�Y�T �г"OT(�7��h�e)���c*>��b"O(�p"��1#�a�N�:#��@�"ONq�6���
D�4,�0Ph4Лu"O���R��:!8��pJ\-&R���"O�� +S��F $>� *1"O<�8�R
	� ��Ś�`F�Y�"O��Z�I޴Y@V��$.!�����"OZx�RFѠrt�N,7D�t"ON�uBшy@2��B�0IH���"OP52���1���� �~�hhy��I�<Yce�	_S�:B��t��� �G�<�ƈ�;Z8<p O@�Vj�a�m�<���K�M`�S�Jܟ#�6+��_b�<�+o*�Lم�B�YI�5h3��a�<�2gU+<=��`�c�l�S���D�<	'��RG��x�BP�).44�A�<YQ�U �BUPp�q6����Ji�<y��ܹ88�sIP2�cejLd�<A�I�9�"��g�X][���/�u�<��)�	_
]�4kH�	�l��`SI�<�&�&B<\!��LBvH*���J�<����3GD���f�-ЈA2���^�<�ǡ�<XZ�Y���O�B,r�ŔE�<���%�L,~��#��K; B�ɡ	ZR Y�+(��iEm�740C�I#u��0�e�,;�����j�RC�I�j��T'L=qP���CD�#T�C�ɿ9���+RG�� UH��F#"s�TB�ɚU��m`��G��0|"b�!�hC䉽S����w��?FJI��T�
B�I.�h� �n��+f�YuEߵ^x�C�I�D�50R��r	�`a��$�`C�ɟ`��)3�H*"s�-ha�\�ZpC䉇ac�ۄF�n�he�H�JC��zT6�Ȓ��EL� �W3�8C��?�0���7!�ʗ6	�B�	"NP��$f�� pR	5ttB�	�k��9����[* �� ܦ�4B�)� ����ʖ1���C ����hV"Oh�@�NۆF�ɐ�$��%�* 0!"OP��䇚�c"�2��ShЌm��"O⠐��-0�}#�(/���Q"Ol��eM1��2&��3F�*���"OЩ�QG:4�l% 1�?d�F�	U"Or�U�^�ҝ��LU�Y��D�g"OP�QT=P8� ���1�ֵ��"O��MŧD��4C�jM�K�x��"O��g�^TF2MzSCK�}�x|kU"O6�UL��d�0�	�k�X�B�"O8U�p�	8�:��NV\�["O�Y���fw�[-A:kh"��B"O�\qGP#9]]{��'gD��v"O�}��D0A�,6��;Y<F1�"O,�a����X�!�F �~Y��"O�}� �X�ب�Sd�0%���`"O��	��<?Kv�Ȯq~���E"O���F�	�W$Q�҂��0D� �"O�H�6.��cιz�B\e��HF"Oh}���Ex�S*
lbR�h6"Ox=cĀL�Q����V\p����"Oީ#���oꮜ���Zp�]�'"Om�R�/T���g�#=���8�"Oxh��Ps4��/�^q @"R"O�(476��$c5��,s��`�"Ot��)o@t��-��|xeZ7"O�MaRL�~���٩(\���r"OZ��0�ՠ*���Рb�>���8�"ORx���eJ)ো!@fB{D"O(q ��@�Cܼp@���#+�)S"O�:g�I�0�@�����,�8�"O0�{C�	���HFCϗ�<�PF"O���"@4{�t=Q�O0jϰ +�"O4͑@�ikTZ�$Q�=�t��"O~x�W��u6��:�\Q�ޑ+�"O�c1L�_o��qEB	:4�"O���4���8u��	g�j}	"Opٲ��W?K�r���ו@����F"O����b�6B�N4�iĄey4�Aw"OЕ��X5q����W��k��k�"Or��AG��_�����> ���"O�@2��ڪ;,���ϊN��ib""O������v�Zl#�M�Cά`c�O��@���C���!�Z:`5x��O��=E��h^�^��RW
�?6��Щ 嘠r!�D��^�D���B��;��l:Vĝ.&�!�$�I)�p0q#�d���%��`�!�	��<3�'I�q���	�3:CrC�IpL��!G�	"\gz4B�'ϦbrPC�	.|�af�vǞ`K��
�P[VB�I�O�� ��9vo�`�dȚc@B䉺L�9H�G�8X�α�*H�@��C�I�jRm��L2Ҿ-ZT���} �B�I�	l8�GiN+, ��) eO�ۤB䉄3�*�0Ō�vl�AsB�L��FB�	�o8�x��}q�-Z�˖EB�I;#%�h wgP�y�\3���:1�B�ɤN���el̥U����GI�`�jB䉻D>��ir�E�2��i� ��d�zB�	�D�r��Q�mB�(B� C��&���(@�M�F!�i�,y�B�	6p���M�	�Ţp�ǒA��C�ɷ,TІ�Y�R%Hh�QjC�>-~C�)� 8$��-A8��})$�<W��h1"O�a�� \O<ģ��IoQ yK�"O���פ�F���bK�%��˶"O��1�[2k�P����s^�(��"O�U�Z$^��J�&y�IQ"O�A��d�2��Q%1l4dI�"OHᩳ�_�\�� ��3n0�	��"O0%`�*��B���+$b�O��zS�D���L���n�z0�OC�ɦKцDLC2S�, ��3�C�	�$x$Bf�,�t����s0�C�Ix�̸�J+&�m�u`ݟevHB�
���ڧ��^+�0C�nΟQ��C����mc�O*h�����?R8�C�(P_x��IB�6��H;�bݳ3PC䉝47"9j���S�Z(����"fC�I�)'ڑ[�d�#h�:�c��[(q�"B�q��`�/Kb<dL:` �B�	>vXv�P�	AX<��d&�2,~B䉊u�|,bS� 6W/��i%Kg�C�;[a�92�piة;%�@0.�C��<e�$����-j?���Ff]�B䉜QQ���	c��M��I`ŮB�	]#D����ހ�8��D/�B�ɒ�T�nĢa�*d�p#�=s�C�əF��,��!�⬅���L���B�	�C	R�A5������F#��C�ɼ/�6�st�O/t*�e�G.�-O��C��,�@zeň�8qn��v)���C�	"M؊a�@a֌?�2%2#N�:g�C�I.���7ɖ�\�u�䑥V��C�-kyI�NȦz)�`��	�*iG�B�?�69H�
�[�@�Ѓ�F��B�	��H�a���
���v�H�0רB�	{���§g��w��)�AELg�C�I��8e���6�q��&P�Ou�C�ɇw��Wd*d���ǁ��:���"Onq[�(����k1&I`|��JE"OV�7�/s� tb%Ċl^�Q�"O�癎hh���Tg�*Uء(�"O����,��Gz�Ձ����2`��`"O�xA�/׉]r���LY���6"O�0�Aq �)q�a��{G�Y*"O�ݠ'/�>:�T���H�~6*��'w�	ß�F{J?�i����n� ��j�,��cg�!D�T�� f�:6��8Z;���3>D��e�4fL����uz�z�;D�l�0�Ӹ@���W���Cp�f ,D�4��EA����-e�J	JAl*D�p��"�7x�#�IL0%� j*D���B�-�<�ءa˝`�%ID�(D����,�(s����
�V
�Őv�'D�,��]#p#�48����7���i D����+*�A� E3i�@0Щ!D���d	+�`x�+j�Fp�£2D�8hB�:�Z�{ !G[/��K��6D��ju��q�(!�D c���Y�6D�x�`F� n��8��A�T�f��M2D������B8����A�4�H�E 5D��x����~�CF)C0L�f��e�5D�\ꓮ[�[u�0��+-�e�ҧ0D�����T�UF�A���&7H����k0D�hp���uOȵy��G�#��a1D�L�:D8��`9i$.�e!;D�� �@;��X~�ђa!x���"OΌ��/\ _��`�Gv1X�"O�����(k�L���/T=��"ODȻ��\�y J�Q�A��0AB�"O���
�M��D"
3,{�4rS"O�ĉ#�M����*Ƌ��
��X�<��%A~&�i�r�� T���)y�<�`�@�z#R\y#e�'.x�!��E\x�<V$(X j�:$��[ʀ�BN�������FJ🜖�(OFX:(�I�΁iA/Y���u��"O�9鱢�6:g�����Gq���"OJ-U�T4B���#Nu�!b"O�e�̗��`ș�'WҠ2"O��H�NY?�8Ě�CJ�b�� �u"O�� F�e��Z2���w@�8!�"O��XBV�&���S-�9Ƥ�u"O
E�6�z�B6Cƍa�R��T"Oj�v���~nZ�Aw���H�t"O�i��X��ۓ��#R�l��"OZĂwč�1_�E M�uO4m*�"O ��r8��%/>�d�U"O~�@tǖ�OKJsUY�@m�)��"O�M���( ކ��lB6$V.5z�"O6Y�6ֺxn���@�ڎ��!h�"OB5���" �hm:�*��#�bh2#"OZ}��	�Bt�cu�(M �[�"OL9��

7rD�8%j]�7H�8�"O��fF�1�HQX�J��I@Հ�"O4�E�(�N�0��T>f1$H��"O������ZNe+ �±6&�غ�"O|�Y���.g�شz�K��Xi�"O"��"eT������%0u'�2	�'G$P���6V����쟒;P)J�'e|p�e���pBd��tS�'�jYr�O<>�< �s'�'H� B�'X�"�J�(r��K�%ح=�j��'�����ڋH�ru��m��4�e�	�'�`}��6 �����:H��t�ȓY`^���O׿���q��M�[ ��ȓJ�ڈ�0E8L_P����Gh<�ȓH]�U��<I��-h"��*掅��O�Ԅ$�5��q���X
����xh(����!R�m�0>�ćȓOq�`�Έ�S$(局)S�^vPل�e��m��/+q6Ĺ��޶>�2!�ȓ!���q�l�6c�2�괣Up�L��m,8誄�:"n��R��0���ȓ� �;����0͂���(Q�a�ȓ"�*=�eHVx|���S�$$�@��ȓ���Ñi�'��P��X���`��-h0��ʗ�� ����ȓ�Ȫp�W��$�'a�F�z����걡��̀��E`G��#�y�� x�����D6'��@�_=�y2�CTpQ�Є>56�yG*��yr��F�x@)CÁ�zFD�2F�܍�y���im&9��A�:��4�"D*�y��0l4�T�(٤���x@ʱ�y��6�\4`p)����rl��y��S�%5~Q3"�آ�ؠ�fGG��y�OU�6jb
ط}�l��ڄ�y��=f
�i�H��}�v»�y"���852�*J,�- а	�-�yr'��*���ie��v�2!��ɉ�y
� ~�J�fF�rդ\*f�E� (m�p"O i#�j�9i:��s�Ԁ	l�k�"OH���fJ�B`�Q8�fյo�a
�"O��9��ÂD���i�T��!�U"O(e�g��;�.5��cһD���k�"OE�2I@A���α@����"OXQ*#��޺��B��<yq"O�F(�Ll��D���
"O�Tۦ���De�|�&�Ȓ��$"O�l��GJ69�L�3k!?�Z@�b"O` rs_-6`������6��CG"OQy���_�NpPs�՜Y����"O<My�ↅ6:tH�6�ķi@�d�V"O��3��W�5���tOl��"O����ۜV��yR$�\��`�"O4�Y4��Yhb"b &���"O�x+ n�W���Wf }t�)*�"O��ړ,[�:v��pdօ=frp��"O$EO_�'��R�J`�t�`"OV%�e��T8��K4HPb1h�"O���%�8u����+Z �<���"O���o�����@J�m���E"O<���<Q���w���,��|��"O�\3�O
?/�)0��G�@|�t"O��%T���3F�R�wA�4"O�	�P"秃�0	�����17!���<rH�Z���m��	q5ρB�!��[,e����?U�b�#��g�!��uO�z����y���W�N�`�!���^Q61��I�y
)@1�R�6�!򄏓S����a�M� �q�9 �!�ִ]a"iJ�X">ʍ��F�v�!��S��Ҝ��h����K��!��{�|���J&m�
�d�8J�!�Œ_����' � J�ޤb0#D�Ar!�D�hX�H���  ��0f��MC!�@�X`&k�,� �{s�U*s?!�7[ ���M�R�$��a�;!�d@���0	Y�WL�(����%V!��ٳrt���U��"q����47!�I����7l�?1����5w!�D�y-����
��)h&�Zlh!�DL�]˴(�b/�2�ƅ��B�&"Oƴ� kC�JH�@z\$<�u"O��(�Q�d��`�� �`�"O��C6�B�ݐ��=�$]�@"O��@2"K�/5*���K����J�"O�%�fm�4{����k�d���r�"O:a�	��@b�[���c��2�"Oz�3��z������C��${u"OB�Ѓ�]�8�Z *M���C&"O��)u�ݷFd�YIR���=�!"Oh����))��+&h�)�0���"O�\ȇm��W���hdɿ��YJ�"O���I�?^&^,����R��3�"O H�V��;K��|�t��"O��X��F1e�pe3�'ݜ;�Xir&"OҌS���/!>%�0F5_�� ��"O>�2�=�r���BZ�K��)!�"O$ ��ϕw����0 ��?�<�I�"O�륅_�t8�,H�n]2t���E"O�If�~��!W��y�:\1�"O�y��bK�@�����A1q��|
�"O(�+�i2C�\��"A��$�
�32"O� ��� ��G�Τ��"J�Q!*�x�"O��[��!M!h<����c4��P"O�a���g�t�$�'%�P)�"O�-��C^�`���Ġw۞�8�"O���1��j����N�	��Y�"Or a���N�X�ʢ͍�_OҜ�R"O��� ��|�@���.FV|4��"O,�����z2�@�>a27��A!��Ў����d�/e�0�øm !�$N
}����!�� ���箞?2�!�P*y��(��ȏ�o��!u��J�!�$��e����K;j����J^�j!�D�!{�����.ʹbb}��hEA�!�ޞL�T��1"�W�lbN�T�!���9Z�4��՞X�`�`&�7|!���7������sm�����,Fa!�Du�dGS1[\���KR�$a!�dN%h�0;V��)3s���֠�?;D!�$�)i�޼�SM�|y.9�4���j&!�$��t��DƀM���@G��!�d۟.N�y�ň�.`��)� C�3!�䊉��T��ڸU8X@ѯA�V-!��"��Eڲ�[)b����
	y�!�� yByy�i��);R��6�._�!�ĉ�ac�	BF����Z��T�!�43�
qA��B� ���!���!�DV�;	$��o�6��|Q R�!�1�h���&]���yJ�L
�%�!�@�sjt�y�a��+�6����!��W�&�±�K�Z4 ��M'3�!�$ _xpx�j��i���y��߭'�!�E�PPa��W�Z�`5���8'�!��ö_�<P	��):~V�R-ڸ`�!�
w���PsE �zt����Lխo�!��ٜg��E�e��;]u���ťP�!�$�3`�9F�C�8��Axe c�!��ք"�04걤���x(�!�$�)q�ac �h�(�c�����!���"��	��	�)S ����[n�!�^*NTtZ�@ �>�����N�!�U����7�M1��PJ�8T�!�$S2���se��A���(T(W=I�!�DŇ5|x�qwM�.��t �f̽q!򄅲\��ڤPol��&�'qY!����Z!����pT|�p�d��+��� "V,�d.� x��dNO��y�)d_֝P���`�\刡`ҳ�y�O\n��
�_�<i�5�y����!�t��&/A !v��IE$�&�y2 	[��e���Ɠ�������yb��12-�b�N�q0!�HA�y"�Ä?�jyݴ2%�u��*!�d�:���� *ܰ����"�!�$�n"��<wѤ���f!TO!�d�)5Ka:�b�<}�0a"�U�E!���� ���U9IȁH�$Q�Q�!��h�aqpbR�pD�92��e�!��N��ؤJ̰�H�fGp!� �+�$�XÆ��޸pt ąXU!�$����2�P�*�µ���¨>!�D�8�ys�g��9eL��HK�l�!�$A%ٮ���Y(X�Y��G"M!�䊌'`ÕS������Q�!�"��1q��1A�a�r�B�!�� �X�*��4Ӭ������n�\��"O>��`�N<f��t�-������"O�@k�*�q�2�8�,��6��A T"OX��ჴdS 1˞�Gd�Ӥ"O���D$�TYhRj�I5r� r"Oj���`׫X���؀)]K80�$"Op����-�����M2&��"O�u(�dS1djTD���ͭu!���W"O�u@OC���J�R�j8hb"O���ƀC�y�,IbBnN�vr��%"OJep$�0S�"!m�-VX� ӷ"O�,0s�ĶU�@#q�ȰL9�E[�"O~EU�@z���q�ɛ87*F0�"O���C�L� �f!
G�N14��E"O���2��l�
���W�-�LR�"O��{��͵/�
�(&#�$�ъE"ON��n\����Dc�E�<�w"O�ejN =��Q((t0���"Oj=qf�@@�(˵�-6"��X�"Oҥ�&�N)&+�À�������"O��p&',���� F]�c��u8�"O�`�����1� �=�L���"O��H�	����F-R�8�q7"Ol7!�U
�t@!KR8;�pS�"O^�0��("�5� ��5-6RC�"O���u&��/f�M[ǩ�9�H\14"O�:��R9S��&�ܓ/�x�u"O��p�쟑k�z)���
�7@Es�"O*�r�2�6,AbI�9|Q&Ep�"O�Ԑ��0MV�PA+�<1�`$��"OD	i�䌣	V����?�p�8�"O@!U��2A3B��A�λoq���F"Oʭ: ?��mR��˕hmD�"O�X�넪q>���q�A�U�#"O����N�0_�$̑��I�ҕ�c"O��5�W>���#gLP/V�� "O�x�@i��Z `R� �9ZG@uR!"O��6d w��8�7o� t�tY�1"O�AoL�.P���㈜�m˴���"O�I��"�bcgՑ�Ft�"O�ix���
Z��7�E�4� e0b"O�֎ �#�L�Y$F�Z��ñ"Of����+��8��E-���&"O��W�P��:q\���Z�"OLa��a$��1��b�%�"O��X5/[l��8C��-w��-��"O�/��a��L4/�:��S���!�I [d�r���X�:�-Z�V�!��,D�dE�J� oJ�Cv	i�!�Ćt����əgk.��_�!�DΗU�8iS"��'F�J͘Ӏ��K'!�d������I��_?-C S�'!�$?�F��Ǎ��aO
�'�V>U!��ɁX����g6�:����9�!��+�(�aU�ǾL�'�ͬ0�!�ĖW�!Q�i�>}��8q��,�!�����t��g��T��M�bÅ�{4!�d]
���.F%�����"6C!���
fcI��ڸv�u����M=!�D�t�x��3�Y�.����5!!�u�� @V:���,Ay;<��"On�p��K����]�@�J$�_��yr�ˊ%���``�L���8��b��y��FB4.<�`FRj�������y
� �<�r��{vbT�&�7�z�"ON2V�֐U�֨Bb`̏��SP"O�]��B_i�v�bp.Q�i�x""O�Y�a�>3n�����<&N�YP�"OB�۲�T�+�`dz&		��<P� "O:蹲L�}_�飀� X"l0�"O:�	�J��0#��y�f¥#����"O��dL!H&
�E�F�(]9�"OƱ���
��Hu��V(#��{�"O�Չ��P3Hp<��@�n��ؘ�"O�hDCز~v�<bjӓ^��d��"O��s�a̮KiP�RI�$k�b�H�"O�h�GR���]��	�b"OZ}���S��(s�J�"��i "O�Eᓈ[*�ʘX4(ޟ}�(��P"O������3�bm(�g�����"Ol��N�M���V�̍r��"O^���j 1�x afS+QT�}�v"O�uq ��b���#����x&�0p�"O\�9R.�3'D��j��$=i�"Oz�*��*M ��3j�4t@ܸ�D"O"���GI�">�ćX�v�2$��"O<]���g�.�6G[�r2a��"O��r m�>B�+�g�+Y�h�"O
<���ǨGJR<���'E�|Y�"O*�P��[\�`���^���A�"OP�k��L�p��y��Y���r�"O�apD���xiN��떦_�z�P5"O���a�¯xЬ�鏼�U�E"O��Hk�m��I�@Gԓf�ԥ:�"O��b�֟-������$��"O��"/�=x/v5�o�5o�����"O�S�"�(��qh���)Ȧ� "OV��&o�k6������}����d"O�I�H�<F����U!���"O��h��ա+w���dK׫�v���"O�Q�q%бr�H�%+�P��trQ"O�e�tj��.��@D�S6m��BQ"O�p"���+*^<�bh�Mΐ��F"O������vN�)&hޔ@�.%*�"O@�b +�8Sd���"�2�C "O��5I
$\�Ha��/[V��i�"Oݓ4��-�X�9�CZ�X�~���"O�d�@��z��U(�Dy��ye"O�}�^<6 ��B���gpp���"O�J��20���ir�4iY�����~��s��F�&&�9�E
Tp�!��Dkm�+P-L�n�Q7	�H�І�}�Y�V%�|�R�ǧ>U�A�ȓ)�ڕ��,c�ar�/�4لȓ0�D�D��+*�X�y�FЍ0X݄�>V����:��퐄*�%@W�<��3�\�z���O�J�!� �%��qҠ�MˉPlI��L�'�ȓ0��1UP*!��A!�?/:���%��	��*���8&+����h��B`.����G���1)�y�����&�j�% ��ՙ��5R2�p�ȓZԎ%�g�!�y�5*/ \U��v��z����B2��b��;_F��ȓl_���+�+f����")�Q�ȓF�JH����T�v��#�>�@L���<�cAbJ�i�z���m֮fK(8�ȓx|}���L=l�d)]`� ��S�? �t���Q�vtIѶd�I�I��"O��� L�꼃".���p�"O�8ȁhيD<�U�d�D�j�TP�"Oh�rhW�#R� �'�=qL�t��"O a��rcNU��H.���"OX(aA�� ��0���S�0~���"OhVJ��(P���!`F%����4"O�L����u����������Ԝ�@*T�)�'C��A��ǁ$6�����n�1i���ȓ"�^�چ�R9j+�8s�b��H��|�ȓ{��Y5�&db����kș����ȓ:����!��&X��B�)X����%;T@>��B�\�F�ȓm��ܨ��
��ȫ�݁"	"q�ȓ4K\d2%^|Ȥ+c�OA
���l����Q&2Ga���D�� �ȓ�5ꒂH"A�S��R�`�$��}C�����3{�ĩ�7@�(����r�'u�ֆ.B��|2uH^�wcv!�'��2f��	��f)1y��j��O6��'VAZ�� ��*} D"O:��V�ðO�y	���H�nM����?|O��Kf��
>���Ь,T�T2��IFx��8w.���da�Bi/+Ӳ|�`c-D��%��)^��C$�Q�!��ajSE.�O��5���`M��Df0���ϝ�D��u���J�';|u�e�H :|���$ߕc��
�'�����Je8	�)`@�E�	�'PYꕉQ+;ܜ�9���&\70��}B^��F��c��^��y�c��r���0���6X����'�@a֎�=*�t���=^�@|3�'�ў�>	�g8O\�Cr��|y($8�$E_�R��&"O��ˤb��بƣ�%WF��W������WL��`����>Y~�� �K���$?!��V����J�D�0�n�S,E�<��M�%x�4D�AF�1b��]
��K�Ą]���t���3���.n��Ƨ���t��C�<�I�����vQ4]�a	GG|q򥊓&a�4�"a!<O: �����xK�-K�US��3
O~��R��!Z�,�w�S�bn����.]��O�'�Q>�TC��٦5�qZ-N`��Va1O�eӌ�#Z�>��QJX.��4�t�%+K!�( fXa�d喵,���"�^4VF�'b>��=	��I�(E��L���"-# �q�,Y�E!�W�D�VIq�D�jJ<q��]	�!���c����&��ָ��T0"�!��3.�t1����J�B���KܶO"�&�Ӻ���s�dp���B�G����+
&a{B�<�I�R��B`B%�4�0r)��%#B�I<0�H��a��h>��T�<s�"?��	ٻWg6��(A+n&��\�@��4O�c�Є�xy^}'AMU��!�`��\4JC� F�q��W�Z`����U�pC�I�:�tB�=�J�L�3Q�B�I�Y=��"�X�������=��B�� �V]"a�]K�xX"��$�B����m�q�;]�̚�Ӣr+C�I��9AN4#^�y&����<C�	f��SN�-*V ��� �2C�ɨD���o��"�
�H�C�I�� p��³D<Ri��A'@��⟠E{J?��� 00(�AWMS&
��bgC6D��I4+g�$�0:ّ��xg�������Sg��{
r��r�I6i�*�n�8=��IVy�L7��� ���sɘ'~O��gnH� �0�"O���G5�4x�Ǜ%2�R��Q"O�A���ɽn�)��4��i�"O|���(��b�v+d�B�+"�Ɇ�hO��C�sd���4����oY;�!���3#Cr=�u�Qfet|YQO��vl!��S�;���R,1eZ辉Pq"O����� �`q�TQ�ե(Ŧ���"Ob蓧d/}�	�`��-Y�R�:eQ�|�	�qO��<9�hJ�
�d ሒ-|��8CX�<)oBzN�s��+�<�ÁS�'Nў��Z�i��L'1�~� w��=<��Ԅȓl��%�fd�W��8uo�:���ȓE�pP#�iQ `�:���nN9"��F|��ӛI����Qm�K�^�j���i{��IT��P���ػh�ԘP�b�6f@̨ 6D��˕#��wD� �U惣V����5D�$K� &ɒ=�D��}��s��h�4�'��' �	H�i���Y5$��X�!��$���c��"D��{�d�>'vT���M�I�$�֥�������E�fE���&s*^�У�#���?a��IL+[��j�	ɐ����R!�$iO.D�q�V+��7��8����c���l��kZ)� KV>�~�i&��!� C�I�W�Bh���F�&�fX�]��4"<ɍ��?Ej�`ǯ4PJ2tB��78�5�%4D��	Y�oF���F*S@N�� �)�<��哛!f80S
A%���#[��B�(G��h��ز$T�|���� v���Y�IVx�l+�I-3�m�$M�??�8����+�O�r��P�v
X���q`���N��ȓO2���"E�/$���G'�Q�^�mE�������yR-L�#�<��W��=w�eAa�yrON�{R,\X��JG�vd+4'Ђ��D"�S��ͪ�\9?�f�a�m\x� Y�"O�@j���p/���5̐?P��=��i�P���IG�� �S�̴���lH�r�F"=YN<���-��Y�h�@�o.xL�PbW/��Z�*B�$�ͳЪǗ	���z�c�=1����?�	�B��y"���"�� ��	i�B�(Z��B�J�9f~p03��^��B��15�,���
4'��H�>��B�I:J	�a�nCV��R�*G�02�Ol��$��'+�u����22�%	B(�t�!�Նh�^��l��Y�ظ�IFR�!�x����ؘL��80�hKA����'��O?7	>-m�R��^6���&�M�V�!�Ϯ�������{yPyJƦ�*�!�dʡD�y�t���<��S�ʎMa|R�|�h�2W~��Ȍ�;�
��cO������p>)%ۭaJ|AD)�THr�j���1�OV���gQ;<ul,���2{�c�"O^y���=y�9��E�V�Z�E�xbS�$'�b?��n�_�P��,A�]�0m�6$D�l¦��&Gd�`��+L8I���"D�I�AB�;��K7!ʩ_����%h2��p<�AJ�3-�m�G
��Z�.����x��P�)w��JLjE�C�
�y��
��Ļ2�@˪���熛�x��'�$	S�
�78{̸���H(G@��B����>A��$̘41�j�:� ��Z%����y�l?�|�����%�0�x�N�yr�9�h4���?�T���א��'�ўD�'S@�B��ߒV���Cl�5~0h
��� �<��f(/�9&'�
����G�Iox�d7@#��xC�@�Bf���c'D��Q��T�<̈́�h��_y�e�$�#D�X�a)�9>$r]ru�IoP�)���5D�L�@̣,4^�a�LF�+m�ca3D��3���	-h� [u�E
ʐ-��l1D���g/A).�����'z�����.D�0zQd�'=� ���@�8>�����1D��tk�o.HcĬ8thf���A.D���D�I�XVC�"��)��o+D�(jFJʗ!�D���͖�f�d�)D���!�Y,p+\�W͒�$��k)D����Ѣl+�@����J�{DM(D�,H�n�@����˺.�%���&D�"-�� ?Z@�Wh�c��pH��1D�l�M��h��6sɫ$@#D��[G
Y�b,�h�r���^޼�tk>D�,
�g�;yX)��OJQ����1D�@�+�Ġ#��҇��
�0D�t%�H�6��\���3C̩c#D�,@�hֵd�|��֎]�pp�eHE?D��cPoի2={d���@ Lm	�(*D��а%V�d�*5�a�p�I;�/+D��j&jOl�r�J�,��g�(D���g�W.0U�����3��@���1D�\СNðr�ޠ��Vek�|!�k/D�D���^��ʵ�E�̼�'�?D�8��F�*Q8�k��M{XS� <D��)��H�N/9�ʓP��)�U�:D�8!������IqP�Ǘ|Ct��W�8D���/�g�p���8m��@Q�8D�(���o�z`X��C%4|��9!7D�l����ma�1���
M���n5D�\���8
�QѦb��nйwL!D�蛃N��l2!���Q��8Sg�4D�D����`�N�B$�Ͻ?���z�L7D��H�
�`��E�E�Y�wҜR�!"D������q��<Z��Z|x��"D����$��]�p�m��`�Z��u(+D���) �
P�#��D�5�qL-�O��@V��#I$iyHQk�4<c�*/_z�sq"O�) �A8?q$��3�ݞVz�I"O�p�f8X:��FH�"v"O�X��l���JH�I=��	��"O A��KT�{qP�Q��;|a�z�"O��REbP7'�� �a\Ba�4�1"O�ݢ�C	\9��"�Nto(���"O@\ ��B)�h�c4���6U���"ON�ѥ�7-�|D2P(D�Jn�1�"O�[��ݪt���a�A��;8�y[�"OjS�M�MHaP� W�-�x��"O����p_?8$H)�G�
pν�ȓ�P	j�ĉ�fF)ۢe�%M�nȇȓ`����"޲(��XCt�Ŝ"�Y�ȓ,OI��&�/=|��r�M�3A~�ȓ�}�æ+S��� b�3i�=�ȓS�x�1�L�1������*<�L��e4��ө7b��i�I�N�4��Ku�A�S)3	���k>���wL�R�J�-R,�� �lW��`h��1BZ�6}�hD����~��Q��&��I3��3Q1�L`�Ȥ]�q��E�����&B���S�O�	C`��.J녁оFT4�p�'w��Xf�Ǵb Y5@�8��5�-OTp�1�(x�;�H6O� �1xP+	#����ǌ"C��6�'D�X1���
`�AW�I��rN�;��c��v��t��I-2�Q����n"�}ᓀ� -S �<�e@�/ <�i�Dl&�u�K|
���,��3��N,? H�x&�t�<��,e�H+i
%f��|���1/#��b�̀�V��p"�JφȎG��'��I ׆	�/�D����B��&��'	���*Q�I	�8R�+wSj�0� H;������!@D��"��׊a	��G}�`T�C���b�E�5���BP�+ڨODA)�H��(gX�CsJ�)���E UFS>���UH�:��A=y|ȕ�ZMX���I�Xb�`���2	�,@$��=�4�VWS��2�`H" @����C�zSx��%[�7�8`�?���B$1�|h��e%��unU}�<��☨P���a�n�~80�BA�4o,��Ju)���w��.��U�O��h��D��z�8�O�(+`�R)e�,�Y%�N����b��h�a��6��'_D�d�%�ـy�te�`LѮ�uz��)Y���������z ��&�~t��;_\��h��p��<�CX�f�(�$�.:�`��
J�1�'�f�)�
K�{9�)ZFIDHf��M��w���B�X�.���g�bU�5���,���R�?�I�^[�CgJ�'(�����E�Rf�&%+��;2�;����F޴+`�I�>'K��c�^�%c�u��&$ !��/@����y(�" V�)�#4Z-y�*Q�~����Nt�����W��D���D���y�h��/e&�;�d�\��y�Jʚ@�l1�r�ED���k>�a���1+o0�c$D_��YYt��AĜ�B"LYD|Q�i�M��8t��`�b"K�I3ȕ(r��`���-�,�`���>�A6���J%�G铟f�d�XT�,au��j,Ց{�&�9��F`�fg�+�T��)�<a$Ƒ�c|���r�� ����#��e���.Mj(x�L����Ϡ���q dUȈS���Q��ŭ+Ed<�!ۊ#�����3]e��� �)C��(�
�IT�-�FX:�?9��{љ�ń&-���C}�֝�����m��иU�\&�<��SÒHE-���Ϗ^]�� ��Қ>��4�D��o��ذ͟�N�'=����Z�H����)�%l԰yn�s_Phs��y,ݩ����TN�iD.IJ�O�?��]ϻpc4)�ȄHĦ���Lwl,uK���Ҟt��,�N���1���|:���Lξ���h�pl0IK��A#Pt�y��ek���!�|$��nZ.0�qЖ�P80eJs/��_N���^�����ͿId�r+�"[6yS�'�^��Qm�+�,��S6auFP���о��!jR�%W.MC�'E_
��1mK��"�IR�(��U���i���Gh�'� �hX7Nl%�'�R ���� d���Z�|��1cID�KE�4����0�1
ԯu_�����o$���HkڰZ5\�ŇI8 �X�P��w�ܟ H��&b����>-l
��L��WJ�r��>k�@�R��N��u"1%��"a4��fi�?/h$?�ݻszI�XY���ҒU���P��34��ԑ��]�R�$1�%��?C��]R�-yeK�]���
`ĔD�-7Ct��eI3 �m�P��B���R��X��(30��?:�GV�%�r��$G��dx�&�A� �0��А�:�0�Ů*��I�=	 -�7�J��b�E��l����%��3�ҕ�#��O����r�[�]�`�gX�<�Mⴊ�,s���e�6u����-��H�������U�P���Y�9������M��%�􈗁6W�,Р$Z�y��A´j:�d�4�������5E��"����L�!���k�[�@��
¿� ��t�[+K���ňU>6�6�ې�C-Jݢ��T���]�T�Cê?���weL��OE7zӆ4��i����(�Px��AL�DA	kdN���)ʥQ�N)����?P� !4��h�ir%���
�f�+��P�A��qʶ��L!��.G>T�	I�i[&m��\�'����OZ;{���pa����6w�x�"�i�u!QaB����'d�N��|���#n�Dbv�.*����$'�	bL�`�J��,K�H�Q�L!!D�=b����ʃemI(�A&7�,��P�ʈ"�̑���^. [3CH�8
8��x��I48qpB�$�Rұ��#Lf��4#��p?�R`�=�� �'��	c�LL�͆,����"��h�H���rаڴXqx�Y�o1���"cZ�y�͘�QbfX�p/ۭY�v�8]@0���[r��"쑃=��E#�HKN"]����/�1���شR����d![z�����8��ecU�
K4i��p>�����0��Ί�"1�Q��I�n�ǥC�:����H��#�C�w���,F_t����	�28(.T��g�E�t���͏L�%G{�K�`��!�4'�?�֠��.��'�д���̬"��YV�#Ktb���(L=����Qf��x���]�tS��� M Q	A�%|��ak�,�O����I�@�X�G	
��"@��:L�@j�Ġ~��tK��6V3����d$G�@ ��)�� H3�3�B�;r�y���P��U!`���1�"O���˔�n#��읜L����oI(Y�L��F��m���$������u�<k.�5��\N��1��Q�%��)^�`�UL��H�ԙ�Bn]5Y�~��%�K�YǠ-��l�9)��U�����FM�`��mq7���S:�kc��.4��� MN ?�����13N2�"��
��(�c��p�8�D�m�'#���a������ˋ_V��"�)�l��
،ؼ�ȥ!�>)�)�����A-�	[\��_�-�L�AÂ�;<�|� ��``J���lŚ1&�`��/�~�`()�2�L�A�I�8u!aݾE�e`ح_����A
U8��-[�Y����A܎K�lZ8ͪ]�&�A�Y�(��Q�Ɂ{>qȑn��*���H�iH⬴)I>A�	�J䢨���Б���6�؜�DnJy<yؑ,�$L5��*]�{)XTJ��޹��u�q��8����w�ĦB�𭛀l� F-����y-^Db�韻��7M�0J��\�d犟}���$Eخ0=)�J�7N~�ؙ�/�)NW��z#CP1I��T�$G����T��.1>�T��}q�!�e		A�j14�A
=�H4��g^\��0T�BK���hĂyy�<��'��kZ��ab�\��80RE�9ZS�D��U)JM��΀%X������aL���TZ����Z:[_�|{P�#d8�Ԡ0��x��9nJ�-:qᆂI��<�� �1
�
��b	;hA�Z�� ��#Sώ6�J���B">�ۇ�=5��L����Z�|Q34b��[��4�T5��+״@$.��
<6��(��I�Ҩ��ꐇ>�v݂Ēx�O��ub���)D�#_ �
� �0�F1� ��^�VtyR��,[��Xr"�E[ у�Q��\ɪݴJP�q�ˤ{sf9�5B\*]�J�;1����S�]!��	:j���C$T��x� 	̷xOn�ˆ���8KXu�q �$	��Xۇ9o�����6�P���̷zFz�N�L-��-�0\��ધ�5n4��t˕0(� ��+�/xI�P��f�Y�'�Zi�b��k~�J�3k1��+��)H�����"�j�|
�H�B��|���z���qÀ+di��iʤ�$:CP^R`Y2��'>�-x���"'���꤄�h_()a(��f�� 1$���{x�8р�W�^�*)��Gj�a�@��L5I%ĩa���D�6sl�P! �R�P$P0ؐ"r�E��ΎLL"�bA/0�����d�e�ߢ �)K�1�p��1��Y$�b�`��x�P5��%��!�j4[�ś�Qի���貭@�m4��(h��V
X+��v�9�	*j,f��ҨW���;���=ҁ�Fb)�be���8p�������i*n��R��'��sghX�>��N
C2����ٱ_f)BC��b����P$+< �1�`W 7�����r;ʝ��&� JO\吰ף��	���i�1�tD�
[jbA`r>�����"NEJ��شA-D#�G8a�H�[
��
��'-��h���IQPɻ�)�6b�9��B݉.�}��Qc�1 ��#���r)P�[��IQ�sx�̓(�y�u�O�3��ŉSDd�T���6^��ԅ�	�@4J��@nqON(
�)N!4\`�9P�E�-��E�$��"P��zc%G��ə�!ڂ/��L �ჷ9��3�l}�2H'�8�N�vu�y��`�,qO`�1� X#jN�}��%�&exvl�7#�"�)��d�|Z�hR�GG&}0b୻`��)I�!7�����I�̼�w��ZcrX���]�1���%P}�~��e�Ǵ\�		�(Y�S ���<��:�bX2Ҍ!���yV2���ՠv�������	��yӀ ��xT6�!`�*Y�:)�E�:TGfH0(����%���p=�$�C��f�tbB6����eb|�A�� -2@��Ȁ<_�7m.b7&����Dl>��c�1��&Â�]�B�8ز��a�������a�)��}�!O�(�&���͊?V�a��C?�α���.���`T2�"X�/��{�N�2��:N�1�=�̵��mD/��A�W����D�K�b��58��:yّ������*{eFP�t�3i� �����=m����,E&�V�9rc�=X�8�c���g�T�0rjD 1Nգ�o�9BtNA��E	��O��;F�@=A�P�{��=��Yy��O�bG�#4��?�Q�Iܖaf��v��=C�^�3��9��MQ�=gN���b�o��l�D'O0J���S$�%�����-�OJH��L��	� ;��O�7|hu�VŇK�=���35g��j�7mAZPؤLP� +���(1wz]��4�%,Ž!�h�j�f��cc���'�hf{�l����,d������F����a�&�rs,��[.6-��gH(�A�l��S`��kRo���a!V$C�1�fe5F�O��bো�&jX+P�K�A��)hV�ɺ��De�N�d;Z�����a�p�Pl�U	��"�A��d򕫂�)�
%��J�z(n�yM$Z�2����X���ׂF\�'�!:3mJ�]�6�Kl
Լ�2�`Z#0۲X��B<�� �mJ�%�c
6^�"�#���ܨ�J@� 5(ݨ2"�8=��mj�G����I�v!�/+��˓�'�����_�1�*��Կr����$)�x��Q3��4H�7(��N�����4Ko�Q�qfêz�	C9�8��,� 6�
]J�Nq�fuV�' ~�3���2TC�TV���F���`1hE�G�NST� ̈́
3��$a�Wvr
���E���\�`��c4nQ!W�H^�h�%4�L�JUmߓPFfd�FGո�O�2�)�Ncz� %꛼#���`�Ϩu�}�􆁯6�XLh��1��#2lU���3h��0uN1cѨγ'�Fuip� �0��PyU���ؙ�'�3r�v�d&O�V�d%p�	�,t�cnֳKl�t9%
�����R���t�b�	(U�8E��ѻW56`�5�
7̞Q�e�)D�kE�'SR�ѝE��ɒ�3X�aC�� �%�
�9��/ar�!Å5#Y @��ПB����FV�7P�y{�w�NRF����aH�� +'Lə	�L���E�7��}��b��~�PP Co����5ƴ[ �I���U*ĩf�XJtd땂\}��t �@k�����O"�Jb -jxU�4oL,2v�(x� �iܓ;m�` i��bEàK��}kr��sf@��\❏-�����<y��yȔ̆�B'�٨PY	Y���7j�O�j@"��$��n�{� Y! ��R��Z'5h>��Ӎ�6��2��wn�Q#���<�r�s �"��j�fZ%0c$��c��5��}:���jB\�:���)�҄�o\g�'.Ѐvd-apP�bZ�8�A�Z1�Z� ��W�y@⣌ ��%���Z��A%݄#<����۳�V���R�YB�m��I�/�s 
5���2!N�"�<!�$�8Ƙ 5L��%u"}����-(?�1�F'
�r�q��]�5lj4�"#�"r�`h�������cf,5�zǮǥ�h�)1��1dd�	�' ��)��:��8R�mH5l(ȀBb���~r���nD�A�6��"�ǟOJ����6gDan�l�Z$a�"�N=��	�$>g�I���b%
���T&U�#&_�hڱOKR?
֤�*�'Qc�M1a��hAh��O�Wv�p�]��T�Ѷd>t��ӏa�qq�JE�kHx�s!��R~%�+Ť_ܶa��)�&�Pzd�3b�^X��-[f�\,&ϥM�1I�#"�\bt(3c�X��4C��xb| k"b�`�� �
�J:"��G�N�rT�٢,,@����	6��qi�E�����/p<���)B�|���㆙�0�ʀp񅝀��D^�5�l�鄦�*� �$a�>s���Y�lW�JgB��	E�Iy0H�
�^mr�C�#�ܖ-{��h�$��x�*��N�Jj����E@@p�w�S�p�,�4�@-��l�[�|��'ꆕ]X̴�A(̿pKN�*W�{�hH��E����{gd�?�5
/)m�� Ħ�:&��rUK@�WH���Ϛ4dX�fÏ�6y��@E?j��e���ԣm<��03�QB��<!���[X��?V�)�+Avj�B�pG��Z珂�E�������GE>Hp���(u�<L	�
.Et�;	�	�ªܽ��qSMC1nIqẻ�jhX�Ia�_�@�$�H!�6�	4A�(� �×�R̎x�����a[$G:��xr�Ƅ/�6��MO�}z�����ud\�B��S����qA�����@&�,�&�!эxp��� 0�k0�ˇWR�U`E�f ��5P����
P�"S��Y-��!(`�B)
��b0� �R�� "Ā���� @�*0�E*H�@8�dr M:|f�0Hj��_��DhT#ʧ"���K A�"$�5ʈ�C=�h2�i��э@�r�4���!ɥy/�U9D`�� �	�8|�h���F�Ӧt�<<�T�D>/��&�e��,���ىt�r�{�m��1Sh�y�#Y���(�n;3� ,A����d��4�=��#M�^KVt �BՅ�n��6�Ug@�RRd�P(^M`p�o+L��$A) MZ`����l���b��eF�RB��U�ʍ��gۡ=c�M�"�@��x��]:+v�	�[�b���hsV�\�@b�;�J�*'n�=;Q�P g�FU����N�..I>�ۣ7wb�qtň��������9R��}K|uaB
»8��Ӧˢ�t�5�l$�2(�� �F�'j��P���C�Ҥ�ٕ}�zm��ُ`\ɘ)������\�z�X���V�`s����n���GJՈ9d�I�V�V��#}�w��9��96[�D",�:b���+�Kq�Pt��I���,��M�~*fi���y��I�P�����ߙN����K�H>�l�!��i����`�]� ��ψO�q �m�4c��4cV�[�����q���ٳ؄Ƞ�̟���s��a�Y�t��y���=h�)F�� N��q�`�*m~،�����=Y��3r���O;�@���P'>��P֏�+���{�/$��V�*���s�ı~)
q&?�م��b��낦Ѭ.�Q���(���+�G�6�`}�O?!Р�0��v��$9�~��C'D��0�>d��Ha�6�3�j�<�I�P�
���,}��	�4'��ؐJ�K0����@	Dr!�d�q�>h�5B0��tÖ�I�qO�e[�d�
�0<Y��T�C.���'
��S& Rp�<q�n��c��E�6���?��L#R*�r�<��/Gvs6����y�)�J�m�<���ՅdAV�����6$.8+D��d�<90
�q�LВb��:�E�f�c�<�-O�T��.��=/2���#t�<�B`�!��	EA�VF�+�#p�<��h��!���p��S�))(�vG]m�<yS��3J�|��eS�FE�T �@�S�<pL�eF*0�+2G~
��㧅I�<���	�EP8���T�]�LACE �J�<醇=2"~�0�)��P�a;���^�<)TK�-O�v��$Ϊe�����Y�<y�50��ȩ�铩\��&b�P�<�Wj�h��<����'1$�����g�<Q���NRbi��4ɂ�Q�a�T�<��ձ.�-[Tc�|ih)qPK�I�<���,#�̰`%ώn_�bd��@�<CO��Gz��W�ӉY��@�1�F�<�de@(?�`��!��_֕	�C�A�<ArkI�*YH��r�K0II� '�t�<1��Y�yvE�����T��~�<AB+�k�~p�!�>�RL)�L�s�<٠�A���Y0��2O�ݳw͝h�<�'�ZqX@�!/��L����gMk�<��Z@,�
f����2 �x�<�'�V<I
p�RR�V�j��T#�O�u�<�$�W��r���F@��Y��v�<y3��;M$�[�LF�}Vty��Bn�<y�%9g��	�$�*3vP�L�<Ar�E�(��U��J���X�I�<�â2��4!pf��V��t��k�@�<I0�C�/�̉᧨����)FB�U�<)�R%i�݈a�	���{&?D��"`�p���s)�6@�X�4�<D�����L={�>��3̈��lD�B�8D��a
Rr�h��7j$,�� �6D���	�xxD� t��?���2�2D�t��j�@\9V`��J���huM:D���A`X�;d5��+J�f��܋T";D���$Gj��1X�a��Q#�KRG$D�3!��-w4(jҫ��-}8q��+"D�<ÂB]�74�00�F*��e�7D����V�D��r� TT!,�9�&5D�J"�>���R�ԗ�{�A6D�� 4`Z�'��%H>w\���"OΈ�eI[�u���R'�	Jn�x��O��ˤ�: Nr�O�>����<����"՟m�V�b�)'D��Q#i
*�fp����G>|�2®<��!ʶOK�(�	K��0<��' y��P�@�i�b1�/cX��r 
�D:i�k�s��d(���5�r�"'Dӻ%���+�';�9BG�J
k���>G����ߟo?�2�9L s��;��ra�J�7;��c�L��Cg!�ěM����!e�yPf��7mȼAɔ�Z-Z69Їe׾Z��򧈟�� h"��q%a�):���tD�?�y�\��K�0/����HH'{���`$�~(��BO�)��\�G���|F|�B0GL]���,1��XB��*��O( c�����y��$7������C�B�64�Bb��`ࢱ�X�#3���OB�)!0���oXt9�� +ClL���G�D��ŗ����F��M[S#^	;�<���BP3\�İ4�3b��Z�M��p��͞����I�!�yBI�u����%����Bá�� V��b�ΊX^ɘQ� �5�5��N�����lp��p����ㆫ��}ȃ,W5
�$�"#�ɚD� ��)��G8L|0I��F�ΤrgÖ�4Ḵ�� ǧD�Qc�4T�j̊f�P�А��I�i���Ex"m�?3��X�Ƚ<5�<�%g�V�5�!��Dӎ�'�<�alY @۞��#�΢Zp�V�M���H�!l�x5�M��39"����W-O_(�P��VBڢm�?!b([5ObxPZe'�/��)/�N�Y�%Q�k����\�\����O�qQ͸ F؟o��ٕ��(+�Z�	'e�
l���џ�O�k�����6S���LZ��V�|����-L	m�h�
�'EЖ��7-� r��}1�CJ�c�$�Z$�~��0"��q0��b��|��!v��QQw�g�,�B$-I�#�����%�Bh�ЄɈ�<���b
�z?Qs�ON,řE%����'�8-��'�RK^ag�֡{c�I`�R/h���o��x�b	��Q�$�فbֻ8�����KV�{b�IR�y��{�p-����> �����V%
��	�pg^/E%��C"o	a��Ix��`�H?#t�A��B�qC2й���1����paD�I�lɒ�J�i���`��F��$l֭�d�ƇJ�����	M�z��@j �jz��i�Q�Ė0U�"���+�yC�]9bLC� KjkhS�~���ʷ��"ěd	�`�I
7��_��s��0�*�qҢ���I]�Y�,�GK���M� �Z5X$��k�b�j7=��A�BJ�v.h�S�l��y'EO�2��x��Q�!���"*X�)Pb���MbB!N�*�����O��l9@�P$'三�*,Z�k�P5&`EQ�F��'�2A w��M���,(�丂��$���#/٠i<J�w�2����?b���`5 �,�>Qb�	�U%�K@4R��rH>A5�E�Q��"���%�Dye�1V^\c��\�x� ��^�%�H�0�4�`�2@�t��9�(O~����A�=�M�wlÈ'�>���c��zΎ-	ŉ_�5˴����	��x��Wl�V��q��H��[�[���Do�d[��w��x6Hp�"XkLH�|z�o_ e��EQ�k÷R�~��4�������[����%�]>o�̤�f�0<��ŉE��
Y�����(��ksT=��/�����U�ܼj�֐򶧕28���ɣ ���05���n�8���ɶh���D�k�BU3G�N4+K�I��yb��(C�y�D��]F�IY"�N��Bq�eN&p� �`�D[� �����^�@@B�ÎeJ�iJ�����]�̚d�b�J�M$tY��ʌ	��10׮�h��������j��В�@���@���w�R��F��I�d ���v�������CH�a���
Q�x�Lΐ
�>E"�<8q�dl����Y_$0`�I&�j}�Dg&y�N%�E�� 熬0�,�N~|\�lԢ_T0 Ү�����w49Ku�A9Q�> �֮�e�����T%���o��ҧ��R]+F� ),l���7F����̜6d\ �q"Å:���r3d��\����� -&p�s͍.2K���%�O�����X�:�Q�뒯Xf���>��W%^� b��}{�*��͎�0�<
f�:Ov&�1N�W(dk��
#g�����'��@��!C�cT�$j��I�!6�p ���6R���"ޏ>���c!oU����A�N�ƈ�A�׿�n�a�E���F�:�NR!jb�^�r�h����7GF���	�  :w �?4�Ź�װ_�bM�P�w�A��#^{f9���W��MԎ�)uzȻ#AN/a�ɺ�wD�ɰ�)ʴ/�d�S�ٙe��+�'{�=�sjK� 6�8S��Nb	�vg =��\PK34K�E���2j{�-�j
�<�#$��Kv%���'��z�77�,��b�,rw��BӓQ@pqEO׻=�f���Ա=��IsJ�-ӛu�X;b���AҸ$gX��"�Z:K��&��s,�SR퉂t�T-#�i�?W3���%��3�Db���Aŋ�6�^ 	԰a�H�3�#,X�cE r�N}(��o�ִ@�I�E��L �f�����͋��>�u	��bX���$��Bg��`c�P_�،QV�YIx�i��
1N��	�dU�%DFo��hCD�߼���G���D���A ;�H��X�<!�
1�V�3f���& ا �%_���
�9cJ��h�|�P)%�	5�@0����,<�kA#R���*l+�@� ������#K��Җ 
	�b�B��������)��T:5�G��,N��k�Z,�����a�a1����#���
�)мWg.�P� �e�r�R�	�.��Gz)�$ٲ��%
��iV��X�I�6I:���^�fԂFŐ/|.����$L,�}+�+U_ݰ$�u/D1�0��st�M9g�OQ~ȋ�Ϟ;?Y�Z�g�y��4�I�(<��Ҽu{�d䎏�.%�q!��ٲa�0i�ǎ�7k�T$adB�ք�7~�T�n�@(�e9شc̎A���l�ȥP�D�/ X=!&D:Stf%:U ^�-�$��В|B`��/�(���b�aE(�5��Q ���B�B�	.\91d�ɲ�� �]���Co�
2��� L�?"��!��;7���@3A�ʺ��p"����#�؈6��m:� ��Y�G�9h�d���ȼT� T�A��at��N�����{�oC&W�i�'�i�n�@H�=V�,P�!dx6+$'ȄS���F�H"b�¨ �JðDy�lx�Icp�<F+��:k�')�Fx2,+�	�%H�`&�1xLIx��14�0�1�AEqn�-�!�f <4iҝ!T� ���OPqhv�3������p�"���M,z�>�;��@��
��c�Q��#V)�$dt�[7��2aTx��ͽy��;3+ ������T(���.��6��E �
.l1�>~��<KëY�!����f�P ��Ӈ�� '�T�G�ɴ	:8����$�ēh~lx���,O��{4�X ��ٖ!FE]*�ڔ�K�BFz�+��͏zz~��b]�S�ԈĎ�����/�F�sA
\���ъ�*����R1?���A�OᡄI�/+���b�lߨ�,P�M���*ab,'N�f�KL�����."��z"�iڨ���w��݉�J��~,`T��@�Ff~�S�
��K��bǧX]xt�8�£>�Djޭz��i���-�zS��%������ta����^�,�7�1Fa����/J;Ǜ�g	�j�36Kȑ^�f	�BcC`�i8�H!��<6%F� ɖ���PD_r%Ybk�&"��U;
�ldB䧈
��=���C_Τ�� ƦC|��0�\�'8����'�fxD'ɍ������H���z%�<5�,�Hs'R0H'�'k�Ib���e�Z�S��4�*�ϕ�6�>��S�K"��ɔ��H�2p�� �-ұ�V�7YAynڇ�PA��O��V+��J�LI�P�ɀ'Zb���R��O5ޅ���{�ܠ�!$Ũ,퐡��c\�%��Wk͈LL��2�x9�an��E �ۥƅ�".,0z�j��vȗ aElZ0������h�j!X��'R�y�($h4�L���� w�̵� ˋ('�Q�fK~��)27	܊����q�_�j1�P�׌�"r�¡l�W<J��d�D��9�G_=<�����e�4������$�۱C��'��OPF����B;~�$��п)E���$���G�� k�MRD���'P�h�����t��!�X��@�A��$.ކ$(r�҈��'B�`�D
K��rt�"y�D�
�B�� �-{�J8j��^��rQ�#�|����7�i�~O�-Z�^5��B�)ܸ'n�� � O�tBf-��UH�ˊ �MȄ�G�f��hSeA�1o��]�}4i��Y4;�\MX l�����Ɠm̢��2b�%C���:�h,�
�-'�U:���! _���dRɒ�rK	77���R�H�I�ZN��A%���]�dx�é�?�Ŵi�����	Jry8����ebF�1\vL4
'I��i�0��kf��L /Ś0Nn��*�;G����7e1�����,�!���K��_�yR�6Ɠ}��A�>v���Sq��!c0y��G�ywm��f֤�AL��4>�v����>	V�Q�=�@�Z��!LM�����R��:@!/!�&(�T�ɋ�,I��m� �<�"���IA���Aj�8Xa����y���#������!���z���HO�]X�G�A�B���Qvw|���u~�q��J.y��T� ��`��9h��\g����ˊ_f8毙�r��9@��Kl�'ef0�fL�L��\Z3�K �>�HTFր2k���d�
$6k�4
�O��Amh(�&LN��x
��
"�4�`$f6���r���nx<���h�"��z�/c� ����'af9P�E��,H�զA#`Xu���W T�mؑ���\mL(B��ij%h@%�&@��f �&iLY��w8D��ًctT\S��P�� Gx����6y�D 
3 ]pb�̪Gdb`�$��J��iMȩeH͏j�^d*���j0h�p�]W����V	')�b�+��P立 u`��V�"�O�}ki�8]> c����$X'�_5@�\`��� ��C�U�XͲ��.k�.ts!�C�:�J���J�_��$�F胶>�=9DL@�qp؝2�h�-u"�s��ĢB�XX�眪���
����B�Vb�L�ssҁr@��s/�34N�E�p��&��^h.`J��	)yv�zehA�?`�!��F¦��>qAf׉4��Âɟx�ڈb�L�&ih�8�ʀ�*��б�)fɠa2���ʦ��%��=�f�L���y���L�x�"���#������0>�u��\�n�"4 �<�θz&-J�Rg�./�fe�Ï�+f׬�ɀ�Q�r?XԊZ,͉���o\�L uhл%zY����ܟd��&�J4���#��a��,1,Y�=���8<2�D�'�MD�2��#N�иև�O��H�gǼYh.�ґc�fs&���J�0qf����-1F�Qv�Q�'��T�F	X�V��*�L�c*,:��Ll���;*\�w��z6b@�F��H�&�8U��1B�a������xg����ȝ$ϒd�G9ndܺ'�}�a~�O�90���$��3/�p��q��/���C�!�
L���B.����Q�"/��5ର��0)�dԐ��'�yw/�-g\��d�#�|�aaV8�p>��i�[�>��+�|yB|@c�5�V��HK�S�^�g��!:P�q΄����pE��<~L`xrc�7�B,��苊��D�O����h�uF�����0,6]�=I�%ؖ�$l�d�D�F�����6 T�Y� 郥Nܐl��c۬b�f�'�=���ɴ;0��z6�{��)I�ِ��O�D�C^�$�p�����i"�dω$��Y�
8\\X�V���J���ߒ#�`��u 5j%�J�Ď
"��9i�L�s����"��=T)���`#�l��D}�J�;/W��k�	�7��)x�0��A�7H�L��Ė�2��� nHۄ!H&+�FX��jS�}����6I�@�����$睨k����%Ƃf�r�Sr�ľ^#�˓	��1�	 �p�h�:�'PԚ��g�Ux~�*�����I��h�}��a�'�2}��1q��y�*���nߛSuh�rs'̜��a�W�����0�v��u7��c���7�2Ty����q%�ؚ��ͧxmp���J�P_��IQ� �S���	�5
��q�b��,f�Zl�WJ���@�����(�2����{��Y@	Lt�/GD:�-Q>L��ݳ�!�3F��J�F�	5 ͓�*ٿ~=Ctj �!R~8��3����a���B��R%��9�Ӵ*ɕ�� :$�)AuDݲ�d��@��H!"B��DptF�%jX9�ʗ�&��< �D�G�6�5O�GZ @8�#Lv��9kR^�FA*d��%l8ʴ�˞�&��O�CR0`xrR�N|��a�ӎZ�>Hc���oG2��q�E=����Opq�I� ��1ň��L��@A�6!������?u�`-�c��9�(��9�4TҔጓ$F<XP6�@�c�4�3/�N�4!��Cg��i&( :� x�DAM�!N2Lx޴
,�q��#�-�p�����}5D��`bڶ9t��_�2����Ux¡@�D�F�
t�L<��}8q�:� `L��Vt��T��#S�?�ܺWc�Y�f� 'k�'>5&a���.~?th�e�O�<~t��H��`�q��n,Lb7�8^My�-�%~�99��@$q�p�c���e� q�'��-�]0�Nd��5#���qV��2������-Z��|XR+b-�U1��ܞ`+�qas�M<;�xĊ�(�&��ɩ�%ӇIzU�Rf�q6ع�%/ZV*MX��+mv�Zc*Z�Y���Ffm����t>ԥ�E��S ]�VdP������!^�c�TXr��A}�ߖ�J9k��J�@3bh�E[�M���Գ`/*=�Ot�"��Xg��h6��#8��X�EѮw� �������UH��.۴]a��D�!f�1�#��Y�2���G���%тp���tn�=g��I%-*U5(�!��I�2좓�R�����?I����32���Y�#�!���k$� �A�Ɨ;��X�!]0@����2|X�H^P'�1�%aCT���`mE8h�-�o�/f��;de���[1��z ��� ��6�e�e���%��`>m��A3O^<Zd#�Λ1	D��p�^�Ș@OISp1�ई�T+2�i�}�c�NV׍��L�d�1	E��p�lM4#�Yd Jh���{SOR�1��d�`�јD�ЈF/
�5�*�X�,m݅ �fpɓa���	Ѳb�L�C�jG$)��ǟ)��	֊DJ��O?R%B��f�h���͉&&8���O�Y��1t���D_&�KT.�$L^�T)S��/M�iQ�!1E�>!�;�Ȣg"~�R�/I-�Flxp�i�ȭx#�N#P ��eSɦc?!��)DƼ�У�k�ʷ � V��/�>>Y����[�$B5���"�(��g�'�����!ZW@�P�A��J�aY��~""�;,
8�� �C�9O<`������W�P'��2k��ȒF�F�%�U?Ua{"+۹f�.��v �p���"�L0f.�@�e/h ��1��M�I�h��!���-`� ;H~�d�+]u|@ NN�BU��j�h�'�\劣@C�sw����~�7+�
"�I*ċ�i��r��	A�<1�$�3M�GQ
b�1C�ty"�_�D*��B�Ll��S�z�1��C=(	�9R�kÓV��B�	�L7�e�H�Ղ�`\�r1��DIn�9Xax��ٕ|P0G��U�
��7�G��y�e�8ohmP�ήJQ�ZրY6�yb� 3:��� �=s���9�$���y�-�5.5��7^��jb-Z��y���
��h�#�!X�М��`F�y2ㆄP��I1E�G����'��-�y��M��m �G\�;�x�X�ǒ��y,Z�g���!��Z��в�-��y��0?� �V&eޔu#�,���y�d��	WR��'��X!��(����y�f��o(��*rOW�P��T�$���y�O!M�\�A2f��8�l���	1�y2�<'��h��T2��u�A��y"8�s2�2'��	d�΂�yR��k��h��+̠�À��yr��7��B�W�t4� ���ȝ�y2A�-���3��=�,��pNM��y�NʅK�n��_�8H��� ��y2��8���qw��	�L�k�/A�y���[����doؓ�j}�C-�&�yRDȯb |��m �p[��#Æ��yr)�"MB�a�^#{�h�s��#�y��A Z�P���d܇&y�!{ C���yB�͖b~0��-'蕃�I�y�H_	f�s����X�2I��0?�T�C��t���&A��2����{��R�GܓR[-�Q��w��1R-�1Uq��ٰ�
�	�� .G�a��$J� ��ı�4A��  �D�����$N���т������h

�H�4%R�c"5��Pm!�d�A����:T��KȚ+S�8a�NV�8�Љ#}Ҫ=�%��蝔1���3�*T�@�p�������'��&�)�IƗ2�qe��M���t*ܞ]��'$�LGy��d�B�y�TA3D�T
n�H�t"'��$ڡ�(O�>͢!�ԀLO�D��o�h�����bӦ������J�%+��,	�e�>sR@���^)lP�*��>�v�O�$�k!��U�2�I%��..���@�k�9��USs������0|��DB5�n���)B�5Ub	y�!�{O&�X�8O �RC�����Op>0�֌]]�� E��Q���C#h����ŪQ�P�)�'R�H�P�耮qP�%���E��4(�����O8�a����d��.h��Tz�DΗ>���2�,�zw슖;O�6�R[G�KE�~֧�S�P����KD"��
SDC�A��`�>��@���0|�$���u����~I���bN�~H����'N����3� Z��Ȏ!#r}�3��+Q����O��'�FO��a�S2Lf�����+:��T�T�C�%�t�OZչL<E�4g�%l;Də7f4��Չ��y��v��S�|�a���$}�"5���H������Ҟe.�OpE�ߴKz�c�b>� �$�KJ���h�pe;b�3?�)qӢ�ʍy��)�<k@�ӱ!�K���@�ƾX��$�������56����d]`Þ�$'�>O,R�xL���y
�'��0���2p.���N��: (��
JS?yQ-w��	��?UH�LY���C��?��W$ N��a���y?�)��?,�!�y?J�X�܀ܑ�*D|!�DI+u.�:�	CJ'��*���!�d0s���c��~�x".ϊ�!��F��@ڴ��[�(�B�g!򄍯|�1����
��@��(��W�!� I�>$�V��|��e(Ua���!�D��9:`q���ɯkm�]2� ��^�!�®9����h 26.Ec��BC�!��R�v����,d�f8#��Y� �!�d��>"�Y� $1&V�C��Ճ5�!򤜯
*X۳��#K����Sn^��!���%B�t+��>�Й��l��g�!��S�7�z�ݝF�P=�U�ѩq�!�D>d���	(Ԅ�*&�499!�d�ti�eKɹu�&���YK+!��[,Q�d�g�2@������<m{!�d	,J����#�`�(�,Uo!��'��ňE�_�qe*�������!�d�:M*��T<	�T<0 � �l�!�$>}�	�C��*g�a`#ň�`�!�d�/&��Yba�5w�j(�)H8!!���-��QX�!Q;)��A1� ad!�$Ö`z���j�3���v�Ʊg_!�D�:l
��U�0Gl����^aN!��u�jʖ�R�cX��P O�Ge!���#"�f�����HF$Mz�����!�$ �AG ���S�:�\���3t�!�� �J�`b�ϯ1�.u�Kߓ�!�R�rW`��6 W�{2P@�ˈ�L�!�6K]�V�z<��K
�!��w:��R�DU�W�\(([Q!��	EG�E���	Cܔ�
�A��!��$:���Aճk����c�"!��8Bք\��T�`&/!Y!�D��2��D�c�ZN�� xU�I%�!�$GiC���&��u#��;�"K�8�!�D	�T+,�` ��d�����x!�&4��p�#�	G�`d��nžl�!� *� 
Q	�(<H�%�՛'�!�Dطt[\\(��(K-�������l�!��9���!�ʎLy���ܡ@!�D�'N�0$�?Ll�A
��_)!��y�� ��?*�y8�ǃ0a!�d�"&�ڦJ��\B���C'}�!�d�5ta�gM`*��(C"�hz!�d�6:�´�ׅى�(|��N>�!�$A�V~�,B�JϗO��	���w�!��3vf�8�A��yvp	P���0c�!�����S1M�)F���B�aW�l!��F:k��(1e�P�4�"4[!�M�pM!�$���IP�F	}�\)Ҁ�C�!��b���i�l�(L�~���g�>�!��#F���I0�	�4Y��2(�"V�!�D��z���eoݡ��Vd�'�!�dE��tJ�b)���!eb2*�!�� Xlu�>B��s��B �i"O�e��BQ�|�h5T�ͅZ�`�"O�:���=/��r�B?P_�-�a"O(��íW�d9d�#5���ib"O�8��Lj��*0������"O���f[	��I�7�TbZ򤺂"O,CT��g
@(�#[="	�"O����cP�o�(���%J$#�� �"Ofu�b�X3V"�`QS*Up���"O���/�8dr�5�U��+� *�"O�t�b�йtPB5�T�+	�mI"O�M��C�d<f�+�4�8X�q"O�L(`,�(f��KN�}�JՃq"O��zb^�o�pP[�*�$P����"OV�۲Nʏ��  �)�Q� ��"Of�rĝ0A�0�r�°�^l�w"O��H�E�xA�i=.R���"O� :�l�6��x�i�1�റu"O�HV+C��00��QE�� 3"O^ah�E�yU8u�'��`?z��0"O� 93��kh&�8�F��)�<ؔ"O�M�WBM�W$2(��/E��蠤"O���%(�e��k�n8��Yٴ"O6]3"֎�N�sH3㔡h�"O�%�sCõ+]��`�(�^� F"O Pbș^έ�`��[Į|Q�"OPzs��k�A(�M�AS�"ON`P.�;8)�f��Y�V��"Ov��S�X�"U,	;��8�t `�"O4���.Ο3|����"�(�"O�{F��ry��+��ȞK��XB�"Ob5g�	�L[��X�6�
�#g"OFpA5��eʤ�g4�����"O ��4'�(j���Xæ�K��a�d"Obu�c�� ����gڶ^�z��*O2YЖ�Ӛ<)�E���+]1ޅ��'������"m>���	K
@�6!�
�'��A��`]q���D��7�% �'߬s�M�֘�(݈;�r� �'H���ƍ��%�E	 b���'�؈b�\'W2	#��� .t=��'A8a�!g<Kb�Di�r�	�'2�@`��v��	`ǝ�#��!#	�'	���6��3[CD�;�L- +�I��bN�Ű�a�a ��άH9XI�"O�����5R����d��֝"O������J�R�Xc_�Y,a9�"O�C���P�J��!I2"�ʄ��"O�-H��
:	�.��f��h>h��r"O8-�u&Y�O�x,0r`�����c"O��zWG"��a �bx���4"OJ���>C��	Z�E7QA^؀�"O$$�3K[P�AF΁	�A01"O��0Q)�M�J��r�R?vSz�Ӡ"OX���P肝���	L5���"O ��&�{��H�F�X)5X��"O ����9.���z�c1PP�i "OF)3u/� J�(@�oR,J0["O��)`*G�����-02�٫"Op��(PL[F0�-:��4(�"O\D@�E�9x%�kl�T츍J�"OJ����6?�$�	(�FX�5"Of��B�W���æ��t�N�"OT�r�]1�|�c�dV�v]�	�"O� .�j2Ȃ"�z�`b�>�՚�"O��#Ӆ��l��U+��!Hx��"O��q���2(���@�>5/����"O��+�������%o[� .��g"O��S�O;lY�8b�=_����"OX���BRv�n$�k�+*(-�"O������8H��e�B낈�L��"OL��EĘ�H=�	�'��e	&�E"O��B��],N�\9h��$h�t@h7"OHՁ��r�܁`�T�A�>�Hc"OXA
�$�=����c(��A� �)�"O2ث#��7/(0ِ�2��z�"Otq�h� *�L�U�@h'�La�"O)X�+���qRN،���q"OpUP�.ҝ9���Ҳ,\�r�(���"O4剂nΏN�~�I6)R��:��"Od����ޭ%����(M:D��,�&"O,L�̝=�������\��K�"O�
#���V!�"���"O�x:Cj��a��낄V�B�� ��"O:�[G��Q@��0*@bX݉�"OLpR��d��8��H-_7̘�4"O�8S� �&�#���r$ftA�"Od�X!	C����A3�ۡ!$:�H"O:@�6@C"�}a6ƞ���"Oވk�/	�GkB ���7w��B�"O�����@�	�x`�T鏟?$q`t"O6���gV~;ɚEc!�LE�"O�,��˺�<m��\�*�L@�"Oބ���R���D1g��<�B�qv"O*if�B�pVx@��cF�4�sB"O����B(�c���|q��"Ol1*�(�m��m(��� ��h�G"O�ٻN!4��[�dG9�� r"O��6eӊ?����)�� ��Xф"O��WGV�(OD���a���aY�"O��jբ9 Z�ʀǋ;�$d�'"OH�(wc�"���FG�O�(�'"O���3�\1a5Rac���SC�Yb"O�e�u荗L΀@S�^%V:�Z"O��P�#��v���c�F2*�H)�"O�-A��ʈT�:��G�t� ��"OB�cb�k@�D��y��+"O���=V��Eȶ坦#;X��S"O��戲�
�	c*tѱm��P�!���1\�`� )���Ye�-~!�Ğ���:V*-+��
��ـD!�ā/������B�f�r����%�!��O�x���a�b�Z�S�^�%�!�$Q19G��(`!��@�~�ɕ�J7�!�d�*B!�\�!M�lP��G�ǃ'!�d :<��Y12N�F��*��}$!�D߭�����(�R@�p&�<`!��!t���gH=q��pѥ�28�!�̙-�	W���
a��K�8�!�6-(��]�T9�!��$˪,�!�D�8,i��)Ӡ�X/⁸R�@�*!�F$���󠪎���0��Ⓓ[!�d��@@G_�O��9�U�f�!��̚s���ذ���5�@��'��!���0~
���V�R#w�,���A=L�!�#a�Ћ�bP�S�X�nU��!���f������F����k�(!s!�ę�d�6�AE�K?-R� E,��5Y!�� �1!FFI-<`Lm��çPϖ��"O�lj��ϊy!�
X<,��0p�"Ol����M�ڐY�J�3�^��4"O���+X�_j� g�Z�Y�<���"O�1y�l!:f���CB@�1�"OhTrB����L��aT�j��@��"Or\rU�ˑGp����N��ز�"OT��pn�J�4�+dDű:@D�R2"O��r��.��ys��!V2@iʐ"O���Q��o��ܡ2"��*����"O4��.)|&&�E1�� "O�(��T�ҸMc�HB�Xa�A"O0���`� Ґ�qЍ�2V�2"O��2   ��   �  F  �  �  �*  �6  fB  M  0U  >\  �b  �h  o  Uu  �{  ہ  2�  ��  I�  ��  ̡  �  Q�  ��  ٺ  �  e�  ��  �  ��  ��  ��  �  �  V O	 � �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R��I^>�Z�l�)N�HI��S�6�CJ.D�Lh!Nġ ٳ�fݒ!�҉��,��T�I̓L��@|� ]	r"O<��w�R9{&m�7 �)Aj��P䘟�F{��i.[�����N�&�6��Х�}�!��U��0C�/��10.�`��s����<��-�|����G�� 3�iC�ą�IH��?�������O�3: � � D�<�%L���.�����%*4�U����h���� ��#��]C��5'�.��"O�у1mF�1�dIU��'i艂��O>�=E��܆5�>=��ҡtN�pH���y�mX�~�vu�g��G491ŮK��yR"�0A��٧�K�E9(ʡCI��yb��!G��p�$��i�^����P�y�eɯ0�<Y�(LO0P�3��P�y2,ئ ȷ�ɼE.x9u�yB�G�6�vy�*˰Q����	٨�y���TN>aJ�������"�!�y2+�e��[����,�ű�hV&�Py��G3h  i"��yD�RAXv�<AU��{1��s�-�P(�A�t�<�4 �xA�!A���O�hH�V �n�<�6J_�\~������Q�W��t�<1@�]�)p�bI؈k�FE�F+r�<Y�[.i�T�9Q%@+||����.�U�<�1��i4�T-�dym����v�<�`b�� �����*�K�y�<0��7qz��ekM y�p�#�N�K�<��:g�����+J#^��)�a.[F�<���ׁR��!�jI�\H4!x�<Qb�ݟ]z��۠�ۙ	H�P��w�<���f[�%!j�?���cl�<����E��iH�
�(fU��Ti�<	�!]�hRU����, ;�N
J�<��ÿ[�F�:a�#u.�G�D�<Y�l�&w��J"ٝL�H���A�~�<��M��(P�\�*�1&����/ZT�<)�����L
!*5c��q��N�<�S�]9�Xt��+F�yFiSH�<��E��y�t�׆*	Y(L�É�M�<1RB�VrȲ�.]�L,�`��N�<�Iƽ2����C�#�^Q�H�M�<��jr�, ش��uX|<�)�]�<��#,�<��嬌�roܵ�u%�Z�<Y��V�-5�i��Z�Ҳl	BœV�<q��2 �d�k���T���[��O�<	�+��>e#f	ڽ��z�L�<\�"C�|�AE��5�F�n�<Q0�|���`��T�*�����@h�<9�.K$.0�hV �BW�1ؔ�m�<��L�*������Y(i��j�<�A�s�"ء�ɐodA0��d�<� ��*c� m����T��+�I�j�<��m6$�4���6�F(�vȔM�<Ʉ�ɃRԀ��DO�����j�p�<�U�ǣ0����Y\!T�����b�<�6E�)b��m��$��H�#_x�<!�Ə/Y��j��@2`f��2D�v�<�F���PD'�-?��dX�
w�<	���%&TKw�Z2G5�Y���s�<y�Ņ;ra�i���­-,�*Ԍ�E�<� ���vcV*w�Mkf�G�<:eY "OXU�B����4\�ǭ�M 
}��"O�T;UaN�I��q� �R�D�B��r"Ox,BKW��X��
M(����"O�쒅D������!�����"O�YAd%ϥ^ jY;IGJt: K"OlDx�Ҍ[�<�8e�M�@\# "O� ���@*`���I�?UM��8�"O�E+��	7z�y��K�>M�A2"O�ڠ��>t5>l�4FȲY1
dx�"OVT���H�p���#� �I���"O�!�"�~��)[U$����C�"O0���Р0��ϟ
��:E"OF-�c��p\�娥�=R��(��"OH85�N�n"���&�Lk>�A�"OlmP�j��i@�d��*d^�j6"O����(G��@����.R��2�"O�qKeđ,����n4��`�"O8dbElًf��0���N	0�Ā�"O�ubQA�7��}؇˔�_/X]�!"O�쳲��@�D�/)�4�*"-��yR�ùF-,x@@�!7�,������y������1Q*a{��4�y�MS��H����V�~Ё�1�y�i��+<!��\��|q�/P�y҆� V��(�r����ƙ��ѽ�yR��q;���B�܄��͉AѴ�y�珳Y�H�Ҁ-E
�B-xQ�7�yb���p��U��\�9&�{���!�y�O��r�:vj˕ 1"!��j��yr���P��F�F�yA�-�gV �y�#S=V��a[��9r@:��g%�$�y"���!�֔��ϫ6����	�>�y���k���״0����K-�y2	]���`Ɗ]�T�2�A�m��yB��4�4�;�ǊNhy��8�y���>^}��8�[B��ųt���y�l	S��ئ�McꚀ$���yBb���8��۪W�؊t���yBʇ]h<e��K�0@9��+E�W�y��
<��=���C'_�yB�֡3��ȗ6��T�CQ�yBB]�=İ��ܢK�^������y�I*OM�$����H��-P��J��y�4R4P;c��1��}�a�5�y��=������|E}I��V��y¨�X�U06D�iEr-�Q��y�)Й3��|x�K�6g���p�I�9�y�k͗)q���qgU.1�F� ����y���Ȁ�"�R>7*&y��%/�yrCƆ}'`��M�,v������y"�L�jd��C��;!�q��a�<�yrLͯL������BQ0��0'�3�yR��zPY��Ҕ@=z]٠JԀ�y�*�/j*p�+#5�jP�[�y2Ȝ'��Y�.P�(�TI�F��y�aQD"`<*��7LF�̢����y�Et 2�lU�D\�Z���y�'��d�,����]�@9]+ʍ�yrD��~��Ň�:$"�֍���y2"܈e^��Rߍ9j
��Vg�y�/����s��1"pP����yb��;Sr��CA�$Ѷ}�$�ś�yB���1F�.1Ȁ�x�*YI����S�? ��r�/�;.�8m���
��lZ"Oj����e@�9B����X��v"O��ȶ�J�DVb�x���ABx�zP"Oư�e%��2�T�O��J;�dC�"O�ð��%'
�:�A]=#���T�'���ş���ܟ��I��h�Iʟ��	,#6��B��gb�9��n@$�����8��ݟ��Iܟ��I����	؟��	>,D:����8�;�N8>Am���,�I����	ן��	П`����D�	� ���0j��F9
X8Q��	 ���	��Iß���П��	� ���8��,@��Pb�OG�Y�&U��`ƌyf��������۟���ޟ�����h��ߟ0��9��S�e�(���)2MO�+�44�����	ʟd������ퟔ��՟�I-j�J�C��)��p�b%%� ��ߟ<��韔�����	џ���ڟ(�I�d�ڐ�S�I���J@"=ؐ-��Ο��	�0�	ӟ���˟������I�egpa����knA� b�X�N����H��ʟ����I����I؟��I*]��)�T`�Q�U�s�[h�ځ�I����ß ���@������џ��ɦB;�QAέq���JE�@<�Nx�Iן(�I㟀�IƟ`�I�� ��۟P�ɔR�*x�E�8r���j��_80����I���������	����������3,X0�;s�, �0�G�M�{�2x���<���P�I֟�	ß�ߴ�?���"������Y�_(��7��'/�W�jy��'��)�3?aG�ii:�����x��Qi�+2���Q�Ǉ�������?��<���U��X��ڎ3x>�KTe�%�2�Y��?���W��M#�O$����L?� v��5P@���f6���ä*��ҟ�'�>Q�g@�8வ��-m�Xke���M�%�u̓��O�L7=��<#7�f<Ѐ�1J@iٵ
�O���b�ק�O�xC�iW��֯$=�hĔT��\Z 	�<|��$j�LI���=ͧ�?�q�x���*Ō�3����M��<�/O6�OnuoZ�7�c��� �C�p�|�q�7�<���Cl��l�I韜�I�<��O��Y!�N���9U�������	(O�34�5��(N"�U⟔Z%'HjpB��ҜJ�"�X��iy�[���)��<�u�:�pP�'��h�bb���<Qұi����O>�m�R��|:ѪR'B���#�;ym�4�+�<q���?9�N
���ٴ��d}>��'JI���Ti��p�	ӎ�$��Pӄ/���<ͧ�?a���?I���?�wi�\�u#��J����A���Ħ�jp��I���&?��I�GٶPJK����5� �r@!�O8Hn�2�Mk��iQ
#}bDL��E�nˠa�U�~���]I�p��4/�~bc
W@F����'7p`�O���-O�q�pd�?�(8[�-��3���O���O ���O�i�<1V�i� pA�'휤qU�IK4Z�:�O3�X���'�6�$�I���OT6mӦ!�b/T6X,̤��%� rø��PM�_w�9o�f~������3h�O����7��&#��w��ʃuez��T�	ݟ��	ߟ���]��U��Q8��&Rw���ȑK���x��?I��i���D_��T�'��6�:�ĒI���kEK*F=!4cL�i(E��}}2(iӆ\mz>m��
��Y�'�$8�N�
up��EW/
�)�PH�X�.����~�'��Iş��	���I0Pɴ�s����}��a�6P�P�I��'�7,U[*�d�O���|���
svT��h]�N6�P���z~⊰>�¼i��7�\ݟ�~��&:h�����=� I�8i�h��jC%`P�Y2*O�˪�?�gi!���"o�� h���k�
��A�v���O��$�O���i�<QҺi¾5;7��x=ĔУ���@�L�%�+s���'��6�4��-��DV�=�E@A�SN�Q�H�3U����;�M�@�i���h�iw��RWJXq��OK��'�X`���`Y���/C>��ə'����(�	����	П<��I����]�J�{�bH9G�h��h���6m�K�P�d�O��<�	�OH�nz�5H� ���D�v6"�	*E@��M��i����>�|���M�'���P��m5ԉ"���B<��'�z�����8(4�|�Q���󟘫�"X���A�ɛ6��=a�����Id��UyR�b��|���O��D�Ob�0FϼBT,ɘ4-G�Z��i�6��)�����ٺٴV�V�T�qh�#�Np�5� ���aVd/?���1	8ʼ:�lˡ��=����!�?�3�19�*�S4�͸Xb�㱩��?q��?���?i����O8��τ�B[@ԁx禁P ��Or�lZ�>� �����Đߴ���y'�\&0舰��� f�J�P��H��y�Bh�:n��0 � ���q�'�J�r'�H�,Ǌ��	R�L�U:'
�(v�<K'���#��T�ܕ����'��'���'ZHL10	U�
�ԀG��/ Dn��T�h�4>7~1���?��"�'�?)�4n&�Q�!�h���T�����SDV����4<���"t��E�d����j"�[<v8��hf钸A�0o�X3�I�KE<����'�b�%���'�)��!< ��T��I�
�n=���'��'�����S��+�4x�@C��#�d��F�1Z�]IC��+k*Y2�yj����[X}�Jh�,�m�П�#�L[�!�`�3����q��˸tN�5l�o~b�	�,�
e�E%BBܧp�k� ��#O[1����J�1YV�-�R3O����OV���O��d�O��?�6ޢ/�L��j wA���B� ���I�4qZ��̧�?qd�iB�'® �J��4

��Իh!R�� ��O��l���e���_:`>�6�+?Qv틹f�ˊ.�Z����әr���%���Z
���{�Iyy��'C�'���97/����D��F�� ������'h�	��M���қ�?Y���?�/�Jl�P�օ=tZ�q�Ö	 d�Ǖ� ثO yoZ)�M��'x���L��;B@�����
2o�@@e�4��DK�C&*��i>]������v�|��(�ԅ1�,�*T�!��	1(�"�'���'s��4]���4R���s��E+U�L�[1�ݏP�8@�FG�?�?��;śf�'��i>��Ox�mR�d:��k�ą3�Q= j���4K��&o@
Y{���t*u�m��ԦmyRm̀b��9�7`-nb���"��y�_����Ο��������ݟ8�Ob^�;���U�`PӇG;IX4�*@a�`���
�O���OԒ����N���:$�(9!��D�f��!s�CQ"Y�	�4gM��8O�S�']{n�Rݴ�y�(�9�=���WA�w�6�t�|���TAɶq��x�kQ�	vy�O�2��� (���m2ت��Q�B�'�b�'m剠�M��ʂ6�?a��?��J�-}����F�5Zwڼ8Q@���'
�]{�m�b�IC}rl�('@��V��^,���Q���Y�q�*��٫F�1�P� V!y��2��;ڔ�1�b�;ADBŲ�'��p=̉.�M+��?����?�J~����?���h��B!%�7b�x5s�ɓP5*��5u��+L/f,��'��6�-�4��n��R�|i��
,���ӸI�$L֦�h�4-��v ��&֛&��D��-w������1p�-��l����}�����'f��Oyz�4���T�I�\�I:7�Qc!�	Q( ��I�!Rq�=�'a:6�1�
���O��埀��=���I�fB� k�j�.���jl\'���'���i�6��p�OȾ�۳��8�Vl�A;F7<� 5��C�>�iDX���p��\&�q�wyKK�L���ʱ9d���C����'���'��O?剃�Mӗ@��?0�}+Vű��Z�y����+D=�?��i��O��'sd7D�	�ش�6��/HT�9%
�.�X�E˱�M�O���.���r��*�i��s���4�F��J�=P� UC�h��<A���?���?i���?	���'E���B o����GV�dl2�'-�%k�V��<����AʦM%��+�ܫ6���vDF1�~MX�W<�?a+O���e���
+Gw�6�9?�W��83��Q���CE	�2o�.�,c2+�Ol(SN>q*O����Or��Od�O��%s�lw�؜LB>�V���O��vћv�
(�"�'��Z>��Ъ˲^R����4��2Ģ+?q�Q���42��L�O>b?z&_�V�lx�2f�Y��#ܣw<����1O�����JПDі�|2+�*H�!F��4�0$�
�2�'+��'Q���[��3�4$ؤ��@^U�@m �NH@]ޙ�����?I�r�f�$�{}B�aӨ	Zp��j��9�cn	WT*��q���9#ڴ]nv�
�4���D��)��'XT��O�F�,U��ݫ�[���Y*�`�\�'8b�'�r�'���'�哎^��%ô��-m˂A�[J-���ܴT������?����OT>7=�Р���!�2Q�P)�)ւX���ۦ]�ڴMW�Q�b>��ŖڦQ̓`�ұ�BK��+��c��N��<�+� �3H�O�đM>�+Of��O�Ż���x��肤q6�=�ׇ�O���OL��<AҲig��[D�'�B�'y��`�&:�P!ӢL(�����TC}��a�&�m���M;�P����挲c:��d/�	Fҝ(��:?�C)��u��[P����'b���$��?)ţ9Y1���jB�`�ԝCO]�?����?)���?	��I�OTHq@�r��pi 1Mw�*���O�0m�1{|,��ן��4���y��`e����	ۢl2�j�Ʉ��~��'ݛCo�Z-�%k~�z�z⽹%����e�>F�V �KJ�p���H>	-O>��OF���O��d�On�)�œ�l�\a2FJ\Q�2�+dŲ<A��in:3��'�2�'��O��Ƈ�*(藁I�r�D	pw�Ł#@j�LH���t�j��	M�OT��0q���6Q��)����P97l��)�0��Q��C%	\:S�")T��zyB"��{D0@C�m�NdYcȐ	��'��'��Oi���M��C�?Q����6*rC*.ǈ�k�ჾ�?���iD�Ox��'<�7��Ǧ�jߴ?�Q��P�J�1R�9z�ī�ǐ�M��Ot�1���J��=����[q�_Ҏu`�H�oF8ȫ&�F�<Y��?����?y���?A��>|C��U ʄ0���í	%R�'Bjo�J8�&1����֦�&�HC@��1�. �U̕*?�P����?�ODEmZ��M�'L����4�yB�'��yg��f!dKu*]�&C�+v��/p�ĉ�I�T��'��������쟄���oL(��e ��{2*l��ʛ6U���០��P}��j��g/*	��ʟ���$�M�'H�
�+BI�$���b6M_�@]�|�'e˓�?�ݴ#������Oy�fKY�/J`���͒�(1�$D@�l��!��g��Uv��?ISf�'XV�$�RW��,C*�Ȗ�RpE�e����ퟐ��şD�Iߟb>Ŕ'��7��<iVƑ:��!EWn�2��	*']���u��O�����?�Z�t0�4��A�{���X"����yV�i��7m	#t"�6M`��@o��nT�|�'�O����?� ���ũR?xr�#��XY���g�i�2]�' �'`b�'�'e��%���9#@[�n�E��IIOHYb�4?v�l���?����'�?�Q��yg��='K��6���&�:A�a��95&&6m���E8���4�0�iꟜXs��v�,�3���%x9x�r��;Nh�	/1,��w�' ZT$���'�'1�)�`�P]�!a��[,F�Ne�@�'$��'��\����4P�V4"��?��	;
,zPJ�1
(u 2k�9�hͣ��E�>y�i�66M���'�:P�`'öٸ�o�2���c�O�mSS�"Fq@M��8�I�#�?io�O���.O 8�Z��F�*h�m�CG�O��$�O����O��}���d����*!,i) ��[�Z�!�f��A�-B�'��7�&�i�1��+�0FCPQ2�Ŭ�� �V�j�A�4
"��b��+� o�Z�\�eA�m�JEA�$��	��P�4KʡH$u��IX������O|�D�O|���O���R:�����Ȍ�(�z�j1:Vl����Ζ<�'�r��$�'_ܹ�7�
�TTb1dE$H�� ��>���i�\6��韐G�d��s��4�#�I�?�q�P�^�	n��gϴG��I�z�"A��'��&��'@F�C��6XҰA�s�5|�pU���'�r�'�����4\����49�lq#�~�t�#G���	�uX\���-y����\y��']��/`ӄiy��^� ��`vmB�?'�7M"?����u^��	�;��'`[k�e3~�{�`�`�8�����^���O��$�O����O"��<���쓔@NDUisfI�
�I���I�M�%H�|�����6�|��]�H��`�\4��t9u
����İ>�Q�iG� �'g5��4��$ԻD��p�'0D�X��U�b�$TD`N��?�$�(�$�<)���?����?��䘊F�ތ���i�L-Z���<�?������ަYBjE�P����0�O](8#���<nv�	(��*��D!�O���'Q�6�Ħe;���O	�[�+'mv�p�M�#X�s��$,��Be�	Y��i>��`�'9da'�P���#�(21�ԕM�D4 �mGٟ��	��	ʟb>��'�7��?j��8��3j���h�U;�����O��DKϦe�?�cS����4|:.)�����8���A')uPM��i�7�P�=�7-,?��,��iB'��d^y�T�� H��W`
Gc��r���<���?����?���?i,�F՛��ܶI�12%F�%3j��$�����X^���	Ο�&?��	��M�;N�f�͙�&��p� �p�t��e�i��7mAɟ ԧ�O�~��iC�^5)�!	���o%r����H9U�D�~ڤ���B�O�˓�?���L�8:���Ϯ4�� ^I�,!����?a���?�-O�,m5`4��I����kTu9&τyr��`5l-a�F��?ɔ\��ܴy�����O��a��9�1��G5�CEХSd���'�j� �(�P������4���|�$�'�a����qr�9���S�Y��'���'���'��>��	e�BT�Rƚ=8�ʽB��#r�D��%�Mf��?y����6�4�P8���Q�uL��m�>����A�O`��jӂ�l�\��Tl�]~�rFv��s�y�*BW|:d�1�\4i�X�Su��	����d�O ���O����O�dnQҵb�_^\�EO�}�V��PU�d@شu����?1����Ou�آ�n�004�)�U�-��ڀ%�>���i5�7���@E�D�G�W}6ԁ֊B�0�\��U�7��R0d���I?H��J��'uX�&��'�B�Qb@&2���@B N�{�l����',��'+�����P���ڴf&����vԄG�Tw ��dЂ8M@�s�`����A}"�h�"%m��MCa�̝�l}����.�Э��I4gD��Aٴ��Dъ	� �J�'T���Tܮ1)ASt��-  ��2N��u̓�?���?a��?�����O���[��Q͞�fc@b������'N�'|H6�]���O�m\�1�dT�A*j>bx(esv����������|j�X�Mk�O���H q�0�T��;ȑ �o���`��GeғO���?����?��?(^q ��E�u�P�s)M�&D�����?I.O�m�:T�����R�N'QZ��'�^�pM�X�ɲ����y��'v��E�O�c?���'D�� ��&+ǵn���`�N F�"��n��m��������*f�|d	�6:�eR�a�?M���qb��\Tb�'	b�'z���\�`۴N���2��b�����I�T�`�D�?!�-T�V���W}��w�4E�.	�n�(X���9R�X7I֦1��5�oZ~~S�O(.-Q�	�V����D�̑����aB2�/�:.��<����?����?���?�)�ح"�Js��p�FBYk>�y�pI㦉�F)ӟ,�������W��y�_�X��Hȕc��6J.)��T.�7�զ�����	��6�j� ��n͔AD�Cw�[-qIDePf�}�x$��2u�r�FF�ry�O#�{�����ǡ+���%� t���'���'5�&�MS�ϐ��?���?a%�4d: SQ�G_�~j#���'@R�``��,x�b�oZ��D�4F��9P`�Vh�<ZP.O6��	�#�D"a�T�r2l'?�B!�'l2l�	<o�p(A�K���4GF��GT�l��Ο8������u�O�R��*<=H��FL�BJR5B��I(8�g`Ӡ)	Q��O���ߦ��?ͻuO�A( �1�Q�1�G1p�n�̓A��6�b�z n�5hT�nZ^~RИc���S� �Pxr`	��ܬ�A�çA�X��#���<����?I��?Y��?a����7Ht1� �3`���EP��� ˦x���ퟠ��Ɵ�¢�M,M��q����A�:�����M㴼i�D�8ҧ8\>`��.($,dċ��n��h!D�I��q�-O������?���?���<9�M�9�ఔC�-F��QF�?����?���?ͧ��¦I������l@vE;${0�(V�^�֤����Ɵ0�4��'��H����v�0,oZ�
��P�O�G�DA�q��f<��`ئ�'6D��� �?����tD`�1��@.cU�=��,�0�n���p���I؟���矬��埠��aA�6\��Rv��c�a���}���?9�*D�V�U#����'�7�*��կL=�<�D��8t6<� �X#W�^���Cy��'���O�>�*��i��I�_�~#� ./�����dOY��]���` R��N�{y��'~�'��bV�Ҝ)���7���WVR�'�剁�M���O��?a���?Q*����*@��2#%\�A9И���O�m���M��'���v�P�H�56*-UE� ���ZsaV�ؤ��ۢ^����|2���OF��M>�&�Ԥ����S&/���2�듾�?q��?I���?�|Z+O.n�|��%JT�\j|����7_��K��x�ɯ�M��"I�>!��iĝ���?8( ЭQ��iJ��|�2Pl���rӖ���� ���ݘ*O<��Ш@�_����go��> ű�8O��?	���?���?������)f92�z�昽6P��� Q�q�nZTL��	��IA���r�����a��Z�q`B�Gx�T�জ=�L���I^}���N^��:O\-3F��*i�z�r�B�]����>O
�rD����?)���O^˓���Or��P�e��	�į�t�Z��v)P�`�Z�d�O��D�O\˓Z���R�n���'�g{Qr-���/s�ԉ� _�N|�'�bm�>���in*6���]��O�-I�#՝&}$c�l�":�d�×�d
�ʙ�&:(���n�S� .r�����+�+PU�A��j\BónO���� �	��8G�$�'���Ï�E�9�׎��F��<@��'p�6��6�����O�Eo^�ӼC�N&BSB����Lp�h�A���<!e�i�^6M\ꦙ�s�O����'�R�����?��܉#�\	WeQ�k;������]�'9�	ן��IߟT�I̟��ɨR���rD拻�;���o��=�'�X6��5lǘ��Of��<�i�O,i����3���06�Ҕ5���)�lWT}ed�jYmږ�?����<�|�/ȸ{����`;w��Qȱ��n ʓ=�d9���O� J>�.O~T��m_� Q�i	��O��XH�L�O��d�O��d�O�ɺ<�`�iK2(Z��'��tj�+�[��yBi��tOnxS��'��6�+�ɬ����립��4O}�F���1�.P��x� �C���0Rq�iZ�	��0���OaL�&?��[c�~q+��,;֑x�k��z�֨)�'hR�'���'�b�'��%�ENݏ@T���eR�X���<9��+�*�.����'�7'���GT�3a/H���!���T^p�I~}BbhӪ<nz>IYp��Ц��'%>H{`��(���o�C�p0��Ǆ�3��y�I�x��'��	쟰��ԟ��ɾh��Ae����hR��ðK]nL�	ҟ��'�`7mC�d���$�O.�$�|Ba���4����: ����t~m�>�Խi��6������~�F,ae.�1���6��ԠB�En�ɂ�h;.��+O�Iâ�?�sl&���� �s��; �<)ĉ0�����O@�d�O��I�<�1�i����f��~�P!��C����&#K"@mr�'��6�3�	4��D^צ��b�!�Lp blU�e��<�B��M��i�Ҝx��i���� �H� ��O���'���[�SXi��$+�!�'��	��h�	�0��Ο���@�Tဟ���E�̢8�H�Ra�GS@6���@�D�OV��#�i�O�mz�=Xen�j���*W�����2Ѓ�?��4Z�BR���д��"���	/*�ة�q��*�R@�*�扈+XU��'+ P�IoyB]�T�����Ćȡ7O�z��:-��u�S#�՟���� ��ly�i��5��A�Oj���OpU��(�&Z�@Y*.~���5��3��$G禽��4���l�>Q�.Nb}�0i WpBⶪf~Ra�Ӣ��h�42��O��@�I32�RB~a�0A�o�{�ఄ�\�(	��'�"�'���Sȟ���8P�+�㐖>^ժ��:�4\�����?AG�i��O�m��Q�fo�-l��J��I40*�Ħy�4*��������f��p�UI��jn�DLQ�]�:�z�Ȼ1�� ��	�Am�&���'�2�'�R�'�B�'=&�:X�F[�,�t�(��RAG����Šu'�ԟ\�I��0&?Q���F=p� �O��)	J� �����(l3�O|Ym��M���'��>B��B)"ka��#Q�CT���"��#R'Uyb�o�V\�ɚ8�'�剢+��\r�哪ZQ����V
�ڑ�	����� �i>�'A�6���U��$U�Z+h�r�.�Rq�x ��t�T��R�Q�?�%[���ش^���nӢ����:L�٣�E\W��$��hςe�6�<?1��Q�|����P���i�k���[srebPK� [4���鎋aQ��O��d�O����O.�d?�S3� s&҇�Ɯ�blSa�j$�	ɟH��(�M��,M�$Cb�B�Ob!�J2��VBA&]{��hAa�� �'�87mΦ�#:���nZv~���� ��( �Mu���*r�e���\;���`ܓ���'/��Pʘ�?�dH�#!B�k���B5�}A��h�<����79`�W�1F\��>),1Q#@��2vf�q�$T��t2�#ԒbIB1��!Ө�KPB�!P��G��)0��
X�.��SJ_H�7��YIT `�k��x�Fb�{�"�qU�l����AsέP��9smVLkUFL�~]�q�:p��$B�b��o,@Y�"�/%��T�dDܴD�6��OT���O|�IO������ߴ'��a�@ě@N�	'����ȟ�(�
ԟ�'����sQ! �JȻ/�ȅa�iP�4�U�ش���_�`�x�mZ��i�O��HZ~�.H����! G�68r����ġ�Mc��?�/?�?	L>q��Tf��<�rtS��=?�p2�
�#�MӠfHa��'���'z��F,�Ɇ<2F�ф-�@f^	��ݔeR<(�4l}0Ő)O��D�OΒ�����O�h�@ɟ��й����~Ǟ`0��䦁�������;C㚀����O�Ӈ
�JHɡg���N���MP�S�yR�ͲQ������O���^	u$&Ac����is��qO�_��`�'U>���'�U���	�$h����ѢǞS��@ZVo�up���O��q���	˟��	ܟ��	ٟt��dвc�Aʇ�»
$b����W�Ce�I䟬���P�Ir��T��YV]����a0l�cb9�\�����Q2��?����?	��?��ы�?Is �q��c�g>:�=؆k��s[���'R�'��'B�'�,z���!�M+��.T�>�PA�̹d�j��w}b�'sB�'|�ɍb-�0"O|2�+�O����36�������ݛ��'�' ��'X̙��}R��	ш��c�^�����!�M���?���?��
����O������c�v����n�%�6��3���&�����0���1<��c��F,j!��q0���'n�nZß����8�r���Ɵ �'����'Zc.���<Z-@`e��+J���ܴ�?���������M�S�*���C��2�`@�cP��6 n�(vD�	ǟ�'��4�'"X�$ねL�h�|��4�"]r�q��^��MsBڴDg�l�<E��'����#�	�B��ű#�Q%M�Jy���'<��'3��'(��c���	m?qtJ�:�3�(��B�y����p}��'<R��%#H��ǟ���Ο��{�nAh0H�Ũ<)������n�Yy"E�|�)�[�a��N�D�p�h�F�.�"Lj�Y�x�pM���$��?a��?�*O8�cKN�S��Tg��prx�6% �4y'���I�d&��'7n��S'�"`�`X*��b�E�ͱ��'��E������ݺ<?���#�8½�d@��y�)��U}Zh�e@�J��C�$��'9ީyƠL����⊬����2e��m!!�n]-n|�WaH�M$\���E'�Vl���R$q	�d�������ò��Bҵ��gE�%5Լb�J9&����_>*��Ȓ��e)��)7d<0�S��)�@P���Ԝ��r$ϭ�"@��.��EAN5p��
� �2��z;��;4 �k�d|���ĜS�������?1v.Jkc�LI���=FTA:��Z���i�Df�@q��R �$#��"��V%��Ɍx4ĝ�F�^�Zy 0�R.����S@҈F娅�Oހ��暧7�"��.1`LJ�X b�O"�lZ�H�6�)���X�iG1A(����Vl*�B�	�r��c�χ+�FxcE+UJd����g�'��xsR [���b�o�-��rej���O����?���I��O��D�O���WԺ�FfǜorT9� ���bfHY �	]6�E��>��3�h���L>��J�(���QjQ&�t�A3K��p�a�/�&�9�J�ȴ�}r##�Ty�f-��Ȑ�v�0�Pe�+�x%�	{~Z`L��S����	���cA��7-�jJ�(��i�ȸ��~h<�q��-T��h����,&n�Q҆�a~҈4ғ��	�<�ń �m�vѫhh�t-y��E��dT�	��?���?��h����O ��p>}�.S�c�mR��r�*}�"���<R����?U��l�>|R���w�I�m���,�zȆ(���^�iE��)P�X��&����æa�6�D,w��b��T#���K>q���(�Y1����]I�F�B���#�M�Q�iTBV�D��F��[�$���)�����cH ��U��U�B�ؗa<A����B��K���<�#M���$���N|*G�>u����\)/2�|3��O�<	f&05��d+�(N�GLār$��K�<�I�2�8$@	�X[�u�Bc�~�<9�-������.π`�Pف' R}�<��F�>���Z��˔<͒�)�kB�<a�%�NJ�I'MD�ka��C��|�<�5oثrĸ]����(�8(jU�|�<���U�3b��� Ȍ��pLB7l�u�<i�$��M��&Ԅ��T�%�y�d�	h}L�J�΀,2�r��W;�yB��)z�R|�1�2Ft|��0N��y�B�X%v�����J`^U����y
� ��Y_�gt����T,��}r'"O�L�òA'00ZA&ؔ0��}"Ov�����f!�Ef�(8�%�"O:89&@�`��=Hv���7� �V"Opr�a�j;8����ۏ$��"O@D�@+�P�t�0��~b� b"OT��dN9Y�	{u�1��"O�q���8�H3@ڍ3�^qq"O,��āB�aXX����ȞHN�"O,`h��*����#��)��"OJx��;%Ŭ����8N�x�"Op�#��ըB�Z�B���	k>��f"O���Nk��8rp�\��
u�"OB�2/�
�XSAҍXK5H"OL z0"A�&(A���:K�0"Om�`̈�D
2q��@ۨSH���"O�=0o��:���SVo=���t"O�� �+qެ�G��)B�S�"O��"��:�~��Q�Jlȣ"O�������g̈́�z��"Oh�P���<�X鳔V�e��"O��1��e��  KA��zI[�"O�񺰋�<���I� � gܞp��"OVh
���d�I�@n�	:ܤPq "O�8ڃ,Ĝh2�m�����k���"Oj�B7��3�n��6�1|^m��"O$ ��U�\M��R`�f�4��"O�SeD��	��D+t�X�t�1"O��@��^�(t��@^��"O��R�18' ���dK�WI,��Q"O<���Q+�d�Be�HdfAyf"O����&�D���cR'pVXHf"O\$
��XR���dF�h�p�r"OL��!Ȑ4�ĩE&�zaF��"O�,�U57@&�"2�R�)�LM��O��2�$�Oԍk�%M�4zɻ`��q��L�7�'�ƨ07����	$v��c��-N��P"�?D����Z#SĒ����+{�%"�+�^q���)+�ar n�t�	�a�U�Rg�C�	�~[*�b��	t���J��Ҵy��0鳭B	v�1Oģ}�4��	2Fl0Z6�q¢I;
zZ5��)��Y���d�fi�s�A:��)K<ў't��W.U5v�Xڄ��L�|�J��1e�'"������<�,U���b�����|I,��ԋL�XpG ��v�Y�7F
C��Pː��!7��I�d���=�����/j�đ�h�;C��×�4r��'����2G����		ָ1H����Wnp�i�� k}�%V%��DB䉔�ʴ1#���	��LK"/�I���\;Q��h�xN�%�'�Z��O|�`�Q�A���/0NHP�Cѭ{ vĻ�N?D�X 7��8rz�X3�@ X���kD�%�?�!�_����A����4
�����j�P�M�sɎGY�ѱ�+�o�
8��Iz�p�C�%M!'>��+��+2�!���8MdV��5��:`?-��.C9B�̌�Bj�^���h�#��t����tb刐 7�	��"%����t���a`�?�7-_�dy�5�_&A~�h��ʟ5<���钑�!��<���ę .�����F&�\��1O+L��*\n��Uc2��%�0Q���yW+kpP�[Ӫ�WD�( L��y��8;�����MN��81����l��ADR?^-^���#�3�<�+^w`��҃O�w�qO�8�Q���`D��(� B=JTh
��'�A�Ca�*vXsV�@0Z͔�z���
o,X�{5�eK`��D��G�ب���݈7��zR��l(�A������G�ֻ��'>�Ъ��O90�hJ�D������:/~��'۞z�=�t-Ŧo��yx�%<}�C剹|��bI7�JY�`�U3OI����g�v�r7���j�4����=��aM~�<���z',U#m\���
kPR��'��@K�c
�:?�1j�G_9 5��U�����@.��	p�a�r3l�S����
�1b�0�8"1�>�I��-q�P�VY��� Ԉ�<	F�X�M��,s�	;~V[������ �0��H<,\9TL,7������)���q�ʅ� E��q�.�8��O�G�<��`�Uu�=l�4����K�gp� ����G�I�3�I�䁀�@W�t��}�iɾ@�2�"O� H��݃t�"ق�͆��\$��/�$<�6�F��O�a�%# W���ͻb�(A�fmǓj��5b֧j�jl���0�f|���ֆ"H(@0�L�=`����'bN.}X��G[�	�<���ïv���"���>@b���q��W �l�%靲#Y^���7��+RW �`��޵u. ��`C�%ǲ�?��%cC�J��+�`�},B��co4D��B'���@V^ ���ʢ�&"��4��	`�"l	�-xtf� �����C%F�-^�b�zFE2UȨk@��r�<�V�H;z{"Ay�c�3-�~Њ���4(��	�W�68�����M�S:�"�<�,,h$�ϙ72��%( ��R��ô$Q!=��
�R�<q8����%���(��Cm�f��/�{�\��	�*eh@4h{�ʠ��"؆ȓ ���[_-����A,P`��ȓ�@+Qa��w	Z��t��?^Pq��w�&ؒdE^����[��6$��	�h���*=J� KN�"0��ȓS5N$'ϙ9|�8�6�@/`M$!�ȓ0UF���ŎH��@�/w\�@�ȓ�����Ûpil���U>U���ȓ.���{0��<���i��<	L ���h#s�ƺ6���©��{��ȓ\d:8 ��˥hc��!Ū�	ܩ��{���xӁ�+BvD`"���Ze��ȓC�\�K�e(PtǁE|���mUԙb�E�Q����Df�+rjՄȓx5�Y8!���/r���*�
8ھ݅�vA��Dg\�e}�M�P��xd����	`d���dڲ[�F�Zr�74x��{�|e�gg۴��yr��ع3�깅ȓk0*�K��]�>�:Ub�a��q�ȓ �-� ���c���6�Ӊ"�����T����<BGRi�&��+�l���k�|��	�%}��J������C|VL�G��	^���q��əE,<������7�Ƈy)�� k؞��-��-������N��܁Q (��)��s����S�DliQ�Q�gaɆȓ4�2�![d��@WL��j��@�ȓD< �S%6%�p���//����ȓ#|PWʆ�|U<���S.|�Q�ȓz\M��m�*-��P� �F,�J��ȓy� �'둑B�e�w)
)t7Щ�ȓ��Qփ2/�n#u�D�/���� �&����Y�'V>�B [� ���ȓO�����HE Hi����P�ڰ�ȓ7���qN��VN�I{�iH*p����U���&��D�(ň��G:�0�ȓV���2,�:�^����\$1K֭�ȓU�[ê�N�قI�$�� �ȓ��˵	EgB���ˡ6�9�ȓzL4Ng{2���$^!�t���P��rF�&vb\���kѪ��ȓFpZ1����*ܮ��򬜴!x~�ȓz��	�`̎X�q�0�D�A��S�|����ͥ"2%rW�̌t�걅ȓ�n��p��3H!e��	�����9�$���J��o�xء�H�>9C�͆�`r��'�M�R4�4��7\��͆�D��PPG��c� #E��)vU�ȓF���R4�Y�V,
�YF$)��
\�0aiI�H�(A���T�̅ȓZ����Q�h�RE�ʑL^�A��S�? ����MR6��j`�9B^�"O|͸mRyW�YHEIV��r%"O�@��NZ�DRh�!��'@,|Ԩ"Oƌɷd[{�j)���F�T��%"O���茬F��E!�L�HU{"O��˴c�s$���B����xh�"Oj�b�G�0��M�U��G�A['"O��ٲ��ej�I��!S�άd"O�������ʃgݎj�\�ɥ"O ��Ao[�hh}�f�/� P��"O���rD��S��s�#H�#�fc�"O��+6-�>X ��@M�8=F2��Q"O���[���JD̊M�J��$"O8���-З߰1�
&@���V"O�#�\~��R��/l���A�"OJQJ����f	D1'(�G}��!"O|E�2����JxSǦ�rn�ٕ"O�\��B9�d��M��hc"O�KQ��59��0ze�Ֆ!4i��"O��`f��=�踨f�M�a%"O�Tk�l��X8����[�]J�K"O�P���K�o�2%P��XR,�%"O�L��O�R��m�JǇ:W. �"O���Aʶ,ʬ�hjOtdhQH�"O4x�u&
�=���yԨ��n\u�"OpX���#�*�Ӷ���n��X 6"O\5)p��#G���p����qe"O�	�a	kQ8�)G�H-~�y��"O�#�
2S�"�r�(P�R�"O����A�/:+ʈ!�^$!�\Ah"O�ٹ�gǸ',��ñ�ѣw��AH"Oh�*h�q��P��(t�@"O �ơ�D��t��kB 	�~�('"Olhy��6:`J�HU�J�t�"k�"OP1a��c�t�Rj!��"O``�&g�{\Հu��C�b�"Oy@䂥u�쁨f�_U�t��"O�M�-���*�p�GV$CF��"O�:2�%��PP�_�i&
]�"O �0��\'R���
_">hh�U"O�qS��Q�(�Wi��L(�"O������s)t$xPHW�_��I��"O�|���(_��d���S삜��"O��sV$O�}ƒ��"�&|� ��"O�h��
��zd마v�r��""O����i^�f��L��A��X�"O�����D[6Nс=��={#"O��D���8K���������Ye"O��{Z�K�.��.B.	�c"O>����G��葶��$>H�"Od$C�IEq����!�6$����"O��k���h⬄�fKV�R��3"O���PK�8 ޥA�
떵�"O�`�I�Lh`5��R���+�"OP��7@�)�dEK��Ė�l��"O��B+�-2�l�a/R�6�8p"O0aկK�����B�<�T�G"ORl��Ҁd�
�͘$j��EXu"O�H@��,my�@��NRSF�8 �"O��ce� �,��D.�j��HU"OHE���\9���kY)y���U"O	��&��a��!X��FN�X�*�"O�t����7�`,�h�C�:g�!�$Ԗ3�̒`��;Q7�偒i'�!�� ��رE��\�3��7{Pu��"Op+W��uI�u��%��$U&$"T"O�p��k���z�E�$C88T:�"O<�c�) �p@���O<�M�T"O�:�
W;j��FD3j�@��"O���«�#X��"�c�#h�(a�"O�]s�Q.B:t�ѡb�Gߞ�JA"OP�jG'�;)]�H0 "]�K����!"O�`PeB_�C٘51��_�x(x@"O��jGAZO�>�S&\�H��"O�1i�
��� P%޹	)��b�"O�]a��X%(��|a��I�8Jp�"O܈j�É�4MK�>KL�e��y�\�"7�m��ΏI���uh���y��"ꈒ�"°�f1�䄗)�yi0����
Y�x"�mD	�y�%ˁ2Q�l
4F��Y޲��S�Q/�y�ہh�N�+t/YQFnqV���yr���9�,7JLKm�L�5eI��y��S�]�Xe0� �2�~-Y4mJ��y��̗G(����H��%�ӫε�y�mG-)� Q��t�
d�c�ŭ�yB�-l�\e!��pG�x2�ⓝ�y�"v%@`wǗ�9X��;⍈��y2dR�$������+���;T@�y��L�\��� ��q�{f�Y��yB*K�n�6�r�����!�ܘ�yrH��|������ԛ&��p2`��y�Fl�䬸�d�~\|�sF����y2CH�$�@ju�ɳ@!�8�թ��yb'�o�Le�+��2��UFP�y������Eлz�Z�G@K5�yb���7�=Ӷ��q�
 ��B��yb��i58 f� :>H�%)��y���J����]�,xN鉵���yR�#hv�x��� 3������M�yBG!�.�J�$(��=��ۉ�y��M����+�)V6��� ���y҄8v�4��`�T�X<s5��y���u��!i�}
D͛�cD>�ybZ�V�KBIzl�*C��y"��
T^��PCa��	�ԔY�f�	�y��WXfL�
�����k���y��&:]�d %�9y�x��4BȔ�yEϢZ�zĀ�u���˱�э�yR��7��������,� M#�yB�X kx�8�%�\?v�6���I��y�j�9<.�Kf�­?��űe�˘�y�EX>��ڒfʿ��䱳���y"��N 22���
�����W�yR��
���Aj�64 I�)���y2�R�QY^�[�̑G`�RT���yB��&�u����=f��4�c�K��yr
Ӷ�4qva��YH"�1@����y��ȃ|�uكf�z��[@�Ӹ�y���+;*�ၣ�?	�`Iٗh��y����Ab�������|�,� �C%�y�G���yq�EJ|���1w���y��[2>D��P��&l6�G(�y�`˭X���4	ıS�fl�v戛�~��)ڧnU��[�LߦUj0���կ�8P�ȓ�搃F�N�k�L�
�)Ozy��iІI ����h���%�TY��me��Ӣ�?�f�#��D�mu|���S�? ��yTA�+C��H�L�C���zיx�.�D���O?�Tq�(" ���puk�2Oj�͘�'|~�;4l�av��	ÑF|��a�'���zsϒ�-#�$�@m��E��TB�'���,�,��( 픥I>*X��'�콱wƋ�LX��-<X^���'pd�B�s��0)�@S�~$B��'��l� 3x3:�
�R�x�pZ�'���@AԀ
��]��@�
G�q�
�'f�pC�;j�V�e�͡C��uk�'Į��Vo��]d��Iը6��1r�'�!cg����L!̩2�p�9�'.i�nA�B���K(tyԩ�'#��s%�/jqԴ��aA�����'��9ҩS7P���P�R�xY�	�'5� h�A��#y��&�ׅ.����'a@����*�~�x��/}n�U��'d��Z�@���]�?���k�'�X,Y�E h`Z',Ėf+<�'g�l�c"ڧQ\���A�,�f�+�'؄,�rLՠ,�lz��
{C�d{�'�B̪w
O�I=:��#�ĩcqŸ�'���y,P$<"E�SmĪn���'0~A7%��ze|tɢ@�Q��'U�{��=tK���QbI�"A+�'���Ae��P�X�y�n
	H��'W��(��ϚB�� �%G�3]:I��'0���!�a2 i��^�(~P��'��x!EϯY��\@���.Nt�
�'��T�Aӳ=��4�Q��Q�ث
�'ZB<�U�$bྉ�	Br���'����-N�'�F�h@韾P~B�B
�'�Rm��E\�H�h�P�a��I$��r	�'�$�`���n�tK����d�	�'� z#AI�Ma��I��B6$��E��'F�$���^<Y\���̽+|���'ִa��+p�](��I�!��R�'�A�5�*3�=s�Wy� B�'?d1j�<��=I��K���'QD��+",��ű�+I)jچ���'	2H�o�m���!U9\�m��'@�s��:�}��e@�K�'�ԼBB�W�Z9��~��1)�'U�8Y��%�ɜ	x2���'-����ٳ*�Ő�c��Z!�'�\�R	ۙG�Nq(%���jx!�'��ڋ8'&�3�f  D�	�'L읭(U�ְ �K�&� ̫�6D�z�� j@X��(��!73D��a�ń:>N��C�/�6H��a�1E2D�,�Ec�V���.�>��|�%�3D��	!�ye�S�ܸf0Hz�a1D��y��ߘ:�Y0�BN�$p@��<D�4����
T�@��T�+Aʹ�R�'D�y��JT��)�O-q��-i� 1D��Q`,�4��1A"����0D�0��Ɛ���E�v̵1�k.D�pa�XÖc&�*����-D������Y6�lڔmϊZN��A?D�� �eX�Z�D��cLVjIC�=D�|��)�*B��P�Yx���?D�0ir1��=Q��"�p�C�#D��s�aH�tY�1d��4V,���<D� 5�
�CHv�CA+B�F�Ց��'D�� ���2@
j�dTR3���xqp�)�"O��P�'
lƢ�S���h�"�"O� ��"aiQrB 0#;���"O�!+A�Q���Q��S�c"D��&"OJY#�Ƈ1I���O»U��R�"O���+V6**��2�$ab"OdܫPh��h>t��d��E��h�"O�4r��S�����I��T���"OQi2ȉ�n2�	Ua�j�t<�"O��s�L͙j"�Ep��ˠ:���`@"O^���K�@�P�@�M���U"O�������y�j���M�y�� �"OLu��n�;�4���
�ra��T"O����R6k��PBgJ�wx��� "O��g.[�{���c@�ur�`�"O�xj�0�Z���3P�9�"O���dK����j�/O��"O}A��/5�p {� ���4�;u"O�3��1k��@�-K~�u�s"O<�yN�x�77��EZe��c8!��Zo߾Ĳ �M,( h4-�1
!��Y8}T��G��m�@��,
C�!�$Y�|�x�jT&Xy�����!�dZ�\��i1��O�-,��ˊR�!��˜n"M��ѼY>��fh��e^!��&8ZW�ɝG�H�Q��TS!�ă�?1Xc3�C�4�&�B��S�.J!��D"��M[��I�ld�fB/
=!�Đ�%ļY��jLq@G�!��z��M�B��h�>\{�ċ�Qd!�䑡^�@�@� ��P�a�!��r
�c"Y�;���x��M� �!�]�k�H,dI#�n83��?G�!�DD�t����+d�dM[P�V�ny!�UC���k�5fܢ��({^!򤒶"�~�$EWyxl�y��;%6!�D�7F�p�ۢ*3�<����_q/!��4zu�x�&�U�u�ܐ`�煶p�!�dUj�Nա�i�4Uܬ%�Sg��?�!�$�-F�� � Ή���RťS�-�!�$!��q���J;f���S��r�'V�����y�2���Gŀg��C�'�xAA�ňKI���©�<[#�T;�'�T��!��bHJ�Rg�\�XJ
�'
r�@��ԬX�b,b�!S4Ym�lr	�'��@	�T��CG
U�tl��'�6,I� �1buI$h�2_=�p�'�@I
���)Ed�QaT�B"�N�1�'�6�g��;?��[�oF	�jm��'�8�����8�\�1ő�φ��'ި��`f �K���+R�H,��'*�{נO��f��P����k�'�&��p��6ļt#�e�w� �j�'�l�37�FD��0w��F��%@	�'�l���"1VͰ�����6E��#	�'޶}�MkS�L��e�9r 2�'���C�T$NN�Bɑ�.V�z�'���H.AN���C�Z~)�'��T���W�t�T���G^R��e��'V���Cl�^�nh�#�s": ��' ����v��*����h����'P�푥l5!i�|���T�M�8D��'��-)�EY#$����A�xx"T�
�' :Y�'Ԟx����
kk
Ph
��� - abZL�%��c�=2���c"Ot`1�dư	'�͗)Y/��Ȇ"Oj��&��+Tɫ�k�WD\Q��"Ok ��"ř�ʁ
4b-�5"O&̘�FH� ����C�TX�b"O�9��n 8PX8I�"#'�p  "O�y9!NB���ć��5���H�"O���띊E���zw��<8^��s"ON�"ĆP�"��#��!B/X��"OBl3oܔ%�dⶁ�e����%"O�]��I�&��I���~4��"Op�����&P�6U�WA�x��,;�"Oཱི�A!F��qcM^��Ve��"O��b��Z{��˽&��k'"O� s����R��S �
1�$"O���5�A�Q`����Ò"F��Pj"O���].T�XM�BH������"OP���h5�ٓ2-�%w(�k7"O��q�aC�Vd@\@�!u}�
Յ�@�<D+7�<��!�� 4h�"�O�~�<a�ÄZ�� ң�&�B��!K�}�<q�553�q%�<E3,�s˒e�<!��ϊw��W��R A����G�<)šW4O��mؕ˔ u���2�OB�<у��E�ZM� o!��s͂d�<�ѩQ{؆��DX"$� �c�<ЕIt����0fб�%�^�<��匝+4�g��h��}c�&�q�<�v.���<5'�
?��9�Kx�<��"xP�3"$�L��F��z�<��/p_ԙB��zơQW��v�<��j�J���Q�lԞp�&�D�[h�<	b��c\>q�h�6��{%�|�<1a�W�,".y��Ά����t�y�<�פ�.x r�I�L��!�VP�<1��+Q��"�
4��У6EYJ�<�dG5_Lx\3�#�G�i#��Qb�<�'P�=d�SC`�g(����c�<�W� 8�i�;2��T ��a�<�t ��$`x 	<"��!�g�<�׌�"~@b]4��:)�x�i�!Ba�<���,nR�1���(��!2W�M^�<I��=!�9��Js�� jE�VP�<�1aK�Nc��q�X�E�ܨ�#.O�<���Օ)A���N��9�LK�<��hO�yr�dmێ#*�ق��q�<�0&�!_��X��0z��x�̕y�<I-��{aѣU�,<�5P���r�<	'@��x��ţۦ�:�C"\m�<�bј(��
�&Z�<'r@�1hm�<A6d+�=�a��<]�!P�ă@�<�fL��N���f�8H p�lh�<���"@<4�S��57��<yU)�]�<I�a��\L];EŖ-2�H\k��D�<aRm�3 ��R��+Gd��R�%A�<�t�1l�j"�F+Tm���F'�@�<	�lL
?��u�VJ_'Xp��𶣞{�<�W��1
��R�_V�$$������:\� ����&�H !�+�Xg�l�ȓ/8F=�Ae_4����BeݷF�4�ȓ\Š����Ӝ&T�ċA�ɵKR��ȓ�|%�U@�otX�Ԭ��
ْd��2����.;l)P� K%Z���U����$ˋ&TZ��!�8�~$��S�? ~|�B`�7�Y@4��:F�y�"O�	yk g��	�7��)�.tڇ"OL�r�g�oЦ�����%��DB�"Op��@���s�M���:�"O����AR>Q�(���摼R(�)�"Olث��K�&Ʉ�5��5{[4(a"O�X"Q�
=咠Rp��&h�����"OL� 0_v����<X�B��"O��h`��Č�� 
� ���9�"O����hN!2������'�΍�%"O���j֡|���
e������7"Oơ�RoAV�Vp�NWu���@"O�tIթ�tҥQ��Sj�Ъ"O�@�m+uX:eHsc�)gl9�R"O"EI���ډB���u�rq�e"O���ǓX  @�C�%�fbw"O�A���w���6�(��4v"O�h���Z*.TȦ�		eX"O�{RL�3�|If�6Nʼ��"O�E�F:("6<cӀD/r8h!"O캃iL$?�y�5������"O�e���)��刀eM� �|���"O"�A
U�)-��r��D'�d-��"O�Ӷ�m�"��!bN*K�p��"O~h�Qg�+��c�ʟ��~ ��"O ���E$Ay`�G��9�MA"O��i�Ϝ)bb��R�-VH"�J""O����D��o��(���.5�p��P"O�M��;��KV!G9��y��"O^�[%�Ԛ~�&���!My�Q��"O�a�g��ل��P�@9pV1�"Ov����K7+\t��,�''�(`�T"O���#fC�^�����%��/��1"O���� ;�KĪ����rE"O�l��i��i"�����z��)�"On!h��yMP���^a��U"Oj��) �/	�"#(�9?,� �"O��k4��)~:�𶦃�-vc�"O�� s�Y;-2 �4喃RD��"O�m1eKP�c4�B�51��P"O�<�6f��LW��&�%lV(A�"Od�Z�ї`�!C/��:�a"O�t��o�}f�1��ğ�j� Ёu"O�i�Þ #\�TÃ�F�H� �"OX���9��Z��PN�+�!�D�@k����d�� �rH�C&�!�dIv�M�����}��d,[;P�!�$Ե	�����p �E�y!���
����F�R�A��bI7J!��D
Qê���	C���!�ۤ�!�D�$`f����+>h���^t!���6��"N�GGl<r'��^!�˘f�`(q��_)X�)�VcZ?!��<6m��p��/�j���Ò4�!���P�Ag��t��	�!F�=�!�ʶ<�0�!J����� Ł�m�!�Űu!�	h�gZ�~c��CO!�䙵<h�Q
�f�i����܆�!�d�$?���!���cTl�(N�!��N 
�h$8P�Ɋz�UX�M\�;�!�䃆*��أ @ྐ4&��>K!�4@>u�d�hk��@r���!�U"j�U��$�L��
"	L�!���.N�`���X�L���\�{�!�� �`��Hk@�x���[�Z�"O����-�q׈�:gJ�-�Ԅ�S"O^�v�̂&5�R��ͩ-���"O�\RR�OXRQ��ܧh���Kg"O>%]�?���3A�Q�/��U`�"Ob-�4��XT�y�	ڢ6�0	 "Oz��G�0"Qh6O�39ߺ�$"O���B�͛T�����n�&͎uBu"Oz������y�:ّ��'	�T�kp"OV���ͥvb�C���f�����"O�]�tZPy� ��%W!�)����$ړ����_1����{R�Ц�o��'|a|�BA�(��كE�+2�@e���y���k촄Ig�l`���B��yr��.\�*�:D��)^Jp("���;�y��/a�:� 3��Y鰄�O��y"��̐��ȀR/����H��y�.����-J@�I�?56p���S�y�b�	o�J}b��S=B?l�t���?��'�Q�g	X�`9 �l	�4���c�'� <�f�:N�҄���
'��1�'v�3��'v)��XC|I1��_�<AAIȲ6!<${%/C�9�|,[t�v�<9��11j���[�� �hS�^�<d㍘?��<+�]5�: �G�u�<�ҥ��(��E�U�ӠXr.œ��A]��0=a�FO�;�t<� ���p�˒E^�<	F*�-O�. ��� ����X�<�0#�.�������H� <ӳ�H�<I�%2z���PcgU#1�����A�<� %�(���b�c�e�n�p4"�B�<��!��/���W�b���05M~�<�u�� _ ��)��V�{ ��3�eHQ�<���'�p��c
\N�#�K�<IA��0)����&�!�1��_�<I�o$���3�V�6[ʉ^�<��oW 5�*]��_|<���@P�<���^] ,tX �Ur�6�J�RQ�<ACLQ/l�.�gD	U�����L�<Qq떷���� JQhj���f�Q�<	u���3dIat	V�Z>ʨ�`�[K�<���B4o{\;�
 �F����FA�_�<	EV�$8�����xk��]`�<q �V?�̽##f�>I���˲�f�<�@K#3��	�W!��v|@Ѳ��G�<��Κ?|~�y��óP`��hpc@�<iWBȼfXa�U�줰�^���'&a|�H�	�Ԭ�3%�wp���)�y��N�$��a _�@��Y��
��y�S"&��E�ʹ~�X�.�%�y�솴1	B
(�l��P���y"��l
�t�MO�+���7  �y­ϖr�H+��XF�{O_��y2M�	'�\���W06�{a���y��� �b�0�]�G碹�!V�y�O��U��4*x�(�w�E�y�9���7�БKr���/��yrM��M��EU�-���JY#�y�nK%ZCD���I�9BV���Mڲ�yR/ߘa�Ԁ3�l\IŲ�9��y�$6��"6%8I��U�u���y����v��X�8�"�φ:�y��3f��I�f)B�����K�y�`��{�P,��D_�C)�I[�͐�y
� $����/]dՁ!��J�I�7"O�������s�F�$=����"O�ez��B_�1����$ui��'C!�ªEA����y�JhQs)�)c�!�D�.sZ�A�B'G6lc�T��W�g�!��T�Hɱ��X�-D�H�'0�!�d�B�e� F�)����f�Q�!򄆭��q�%@�ycT�
W��9:�!�䓿)�$�0Q�[<;��%.K!�D��k��C HO"&G�9;BƊ�-i�O����$�`σ]dГaC�2A����
�'�|l�"�.c""�˰NV4(�d��
�'�lpc�^�@��D���&/Z�	�'�6�����^���Kc5��M��'7�\@ ��6�E��2�:��'�P���,_�1 i����S~��'h�#��ײ(2b1K�mҗaj���'F�<`��El�R�y�O�*���#�'Yܰw�Y6/�ꌳ&kB�'�&�
�'(遥��T(<bVBG��&U�	�'����^.v�zI���ܝ=0��2	�'���a&� :z���6֐��'�젩�ʗ"��<B#�^+;���a
�'��\p1���h��Mӳ3o�=�	�'�4�p��ck��p�L&Y(&$i	�'�jɨ�''�xaV5X
�+	�'�.%�^A��)�J��E&�5�	�'�riq/F:.�
���X�R��e�	�'(���wb��Ii�02���G�8 ��'g��*��}@��ݫC� � �'�qpc޶-�
��R�J�0l*�3��x�ѹ[����I:� y�=�y�Y0^	T��pOG���&��y�P��9��P!T�P`E(���y���jٸe�qc��{\�	ɔ���y��W(5h��r�bR0{�"�����yҤD�n:�<��:w����W,���$.����'��p@����	W� =�6A��'�z}�g	~��\3�K�'9����
�'^m#���Ńb`�2 ��!
�'��-3���l�n�HY�)�(m��'	���ʌWn�|��8;��)�'������5�[�0���iR
�'��b!˚�򀴀0�WX�Ԩ	�'��tc�'@�c�jLn��H��	�'�T�"�A>(�t�XW#�{n�Y�'�@���,�?eS*�����|�r
�'���pM�uY�f�J �d�	�'s�13,44� � B[<��'�<4�2!(#E�sB�q32�'��ʦ�O>e=(y����iCZu؎��9OvM�%�������!P̼%jW�D�Od�D�O.�$�O��'<�N$�Z�^�9�&���e"O��H5+�$�Ne�f��9�� "O��IC�4>�d�+���U)v� �"O��1��<9v����;\���"OXhx�#�tD��j�
�pz�"O&�@��ǋatPUŉ 7^����"O�lӡ�» �Xy�g�G?$u��P����ڟ��	ğ��I�\�IG����=1������F07�d�����y�.�1*<n˓爉c�h�����yB�T�w��鰆�b> x���yr� mZT����lߜ�s��+�y�mqUD�O�.b	d�C���y
� L��bX��>�`�K��rU��qq"O�=�M�<l�AK�2%�u�7�|r�'b�'�"�'�?�7#�(B�yz�kU0]Y$4kG�%D�\�d� T�h� ���B�R�$D��󰁌4�����@:g<�QE�7D��F��_��M�R�\�"�4D�p�'�֬x�T`�N�	F�֭(Ҋ7D����ߚ=9��gˆ;T�U@D)"D�t����e|�1�B'�.�ЂL ���Ox���OR���Op��4�D��Q.�dk���9�h2,��<��Ð.|�xx�k�wդ��0��p�<Q�K�`���p�N�@Y����GXj�<��"
}8FjZ��n��v	AN�<i��#�A��^: �9x�b�F�<�'Zx,�(w�܊R`*ы �	yh<y��� [�,ar���7p�
7�_����?����?	��?�����)�5�F4�5HH�B��Q�ѡQ�!���}	@���J�@���ƪI5�!�ɥ�nݸQ��2$�q�K�,V�!�d�;>gz-��d%��(��&l��'q���bF{Z\(C�K��w�p���'��*��eR��ql^�i�p���'��T���U�s��2��$B����L>����?���?9���?1ΟxQ��S9HO�u�pǞ�_�ٙ&"O�����D�K�e��c����"O���4�X�� JE�><�J��"O
5cFN֙%��8��	�.�X�!6"O��E���zP���0!��	v"OH��gB����:!M=P(B|�P"O�eQ�/~�]3�䄋$�|�'Tr�'�b�'��?	���B�|��V*K;Y�졊0�#D� �0���*~��	���?���a��!D�|��-�~�@8���9*�\%9l!D�����U�/��e��n�s��ץ�y")B*J|z���pg�M���y���M�L4�T�� �N��#@Ҩ�y����v	�,ׁq�p��թ�y�V��f�/q�pt�u�X�<�`$�#�젲CZ+g��ڠ�[A�<)t���X<p( ����/q�$��j�\z5ϊ.kX�e�eS �:4�ȓN�v #q���V���$$C���T 0�Z��4���G'$�Ԅ�F��CJ֧Bdn��g)�%��0�ȓ<&�10!�9,hI�艕B��m��-�>��S��?���ʤ"���q�ȓN�M
צT<QD�K���6s�`��R���0S �f�R ��hʎr,Єȓb����u�ݒ<����h��<�n���o_B�6ȝ�!.�!�O�o���'�џ��<�W��$��p��M����wn�ٟ������w�[1����M�^b��ȓUa�j�G��yBG(�����*R��?` �����p"Odi�"�^�b�Nu�d��dB�X�"O �r��8%��p�eK�7(�`��"O.II�"�?	2U�L=?!XD��"O6)�V��;K>�k
^�{��-+C"Oj(�K�� yEC��0�> 
"OT�[�IC.,ɐ�Y��A5[b�}Q�"O��)�΋�0a��(��utJe3�"O�aC��ܲa�A����"Ch^3�"Oℛ���G������<���{�"O>��f�-�<�&�N�f	��:"O� �B$w�� '�=(�dH� "O�8�-:�N�a��S��T"O�@��'���~�kq�9U�D` v"OHM�Ly����2K�����"O��r$��<H�xٳPn�����"O$!�a,��ED
�0���c�L��"O41��']Y>������w�\�!�"Oֹ"6��s�씫��<��B�"O�Śh
>�x]a`��tL��"O�yq�% s��:�OF�!��dp0"O�|���D�r�D�CR�ޝC)0��"ON<�$�@�j���إ0����"O�I�Fl^s�f���./uT�F"ORT���ЀQ���Y�s ��"OJ|9V��-±�glQƺ �W"O�QRq&~��p
�ʐ�g���4"Oz��E��M ,�8�ʞ/
��I!"OP�ۄ�N(���� k����"O���Q�;$qI����$���X�"Of�`�͇$g��r�:��yI�"O�C����w�\I
P"K2v,���"O�Tr�I�ZqfUϕ�L\(R�"Oč(��^-T�P
E�\SM,t��"O�8�qk8[}l BnU6=��"O*dBu��4x_�P+�R�tdS�"OU��(��rZ��0���H8�"OxT*�ŕ�K>P��'�J�O����"O©A���2#R�x����(�"�"O��P7u��Ö[�Fovha�"OX�26�	�`#p�P�LF�,A�x[B"O�����	 �\A�W�Т:��h�"O�hy��V�S4�C4�Ƌ}<�[&"Oڝ���@�`b��8x)��"O�]��!bN�Y��9r��y�a"Ob)�2���Z��K��m�l-��"O�!ie��K7<$�5�j�5y�"O��r�[)Bw�٢���4�2"O�(h���4%�H���r��,��"OƝ��L���YqN� /�n8��"ODE�$�E�O��c.�(Y��UA�"O�Y��~\�-�4A0�P�"O�M��$(T.h@!�P�
��a�p"O���!�I���;3�� MD
���"O���!�
��Ttd�B�� c"O� W��J�X��W䎽T7���"O��X�@C�w�l��Ë�<�pUz�"O"�q���)5G�2&�("��t؃"Ot)��ӊ$�NP¦�\26��4K�"O�� ֮��]�\�@��B.̄��w"O�A�4�����(8Y�v�s"O�L�@�(@�����<�R�0�"O�	�,ȿZ���J�)f��}"O��$F�8a5hѨi�,Er��"OJ�3��֒dt�����?��(�"O\P���'^5�UIc1@����"O��i�`Y<�s╶q����"O4 X$H]�\�0�K��˒ko�d�"O^֠ �-˰�x�bЯ;Y���"OPu�;Eh���|F�A#"O�%[���ǎ�@6�!I�"OVɱ ��$��2'�?%�	z�"OB��%6dB@�:<��@�"O��Y��2G�Z(�1�6����"Oj�B������F��&<R�sc"O� \T`�HS.>X҄�Va77x�V"O� b��v�@J8.+Ra`t"O:}��/?��pcB��".��F"OD8sn�3E�p�)<�:ѯW�<ђΚB����*�-ext9�Mm�<yf X�s9S���B�,�2 Q_�<I�(E�A�x��ʩj^<�H4��W�<����<� jSiN�2~����o�<)V#�p^\0o�9E"�-����a�<I���#��}�*
5 /�i3��v�<q!��T�NQc���/'�Ӵ��yr�O`d�s��áYۂ;�"�y"���|�F-#�j�=O�pS��H��y��C�|����)P�E�}i��/�yZؕ���ɄB�lڳj
9d^��	�'��A,Q�Dʲ�ѶK��e�	�'�@��!ͨ��E��'vBܓ
�'Z�zӁö^s �3VEC�ͫ"OlI)����R&���r�ޅg@z�bR"O�#l��rYqr��5:�"O������9!$�9�d�2p!"O*�qEY.r�8a�b�J*�ن"O�Y0ԧ	���#SA�)v�eH�"O:]�2Mk -�5�J	��(w"O�t3�ο)Yt�;&&3zLN��"O@���"N�/�"��R8j�9`�"O�ժC�&o���B��H��"O ��S��+~>�ys��1��̳�"O�!��t���H�OZ�nm�p"Of��.#-2iz����9����R"O�UY� ��-p�qq��,�\��"O�Px�M��SV�jԨ��&�1Q"Ob��%��V<DY�m�
u���I�"O<QHY?]C����DXNx��"O���K&Lzm��A�S�"O��v��;Ո�ô��kX�"O����(��'Q�h��kas� ��"O��"�ϙ�.tIҪC�6_�QD"ON��b&��Lx������+%t�23"O<QH�fy�Q�A[�AW&���e���y��+R��)b+H+0��y��W�y�%�%5̦1�)@0"Ӥ�	���y���M��s��ڬ�g��y�Yz��h���� �I�'�џ�y2(��pM@����Ȟ�������yB!�!�T�Z�'B��#����y����HŻ�pL�" ����yb�*�@%��T6�(�Р�Έ�ybbʎv \��ֵ~r������y�L'P��eY�lW$��>���ї"O�5(rKS'd_,�
S�	�=�(!�"O��#��	-Fȳ��S�K�����"Ob�[�D�-�A����\zB���"Ox�����k�<;�VY���kB"O�(�s��:s��K���O㖅��"ORy(t��>\�PD�c��	�8�*�"O8�cn��(�XЫBN�2kԨ�p"On �gG�hK���#@�Q`��X�"O!�#�\�[]�廗C��=�L��"O��R�j�O����ռ�͙"O��uNKK��YS@��q�R-��"O�U4�&YUȑ &OԴp�H�0�"O�E�'	�wH<���Y��(Ja"O ċ��
�o��YXvL��ݘ"O� ��q��628��rRk5@�j#"O���aG�>�ΌB�*� ���� "O�1Q��~�����(�}�"Oe�V�Ɉ��1�M�O��w"O����72�ԩC���B�p���"O� dd�b�|1��x�xA��'.�੡f��9��Q�U�O����'�D�s�jIwC���ț�C(*���'^0�@A_�QJ�m�#ى>�q��'8���T�s��`���"Lh�C�'v��; �T>g���捻����'Tj�bR"ǽ���肢M=S"�(�'4x��"��13��9�'��D���'ܒ���N4�f��Ү�,�X��'��!�l)��}T��	�'�^��s@׿��P����1G�I�
�'��9��?u(0�DR1��'jp��1I_:���$c�x1L���'-� 0�	� ����&/U�pp��Y�'���Q���#�!���1#N���"O��b�gO%l��� F��/��3�"O��P��T��=��g �},�!"O���Q��&p�`x2r�R;Q�i��"O�Mc�	�Usn=0o߉6�P�`S"O�d�T�[Ot��d��4��ڳ"O��p!��2o8��
A悪!�4P�"Oܰ;q�B�l{6aq�E^�T�c�"Oh��HJ�}�J4�&�לM�Hِ"O4=kË?�$%�'��5�:�5"O�0�)[�4�<�&Lɐ{=Z��%"OT!@����u:lJr��w6&�YP"O�(R��<G�=��$/���F"Ovx*�#�/c��`p+M�2n�"ON�[��%�*(�Ϗ�;���ۖ"O �P�"^�D�酥B��D�t"Ov������(��2��aE��V"O@�ٱ
P:k�YY�*D;�l8Q"O��#�eI[t])3�Ȧo�vMzD"O�L�0(Ԡ�z��	IX��2"Opi�Qf�.W`�m�� Ut����"O>�+����	���#�a�"O�9$����h��D�eX�]3�"O����(�,p$у�¿QKFtcd"O�`G锗&�I˵M�ZIp!˒"O0�H�Ұ!Yr�� �
�=4n�F"O��I�BL'm*f9 bKW��T"O�9����Uy�q����&
�x�"Oz��� _�zg�<�BoЩc���k�"On �V�<���ӳgP��tq��"O�蹔h# i��'��X�$�(#"O���(VGjV`�oԐ �hD��"O9#�r���P�n�nU�ib�"O�=��d���DB��֙L�rs"O��P�T��)���+,*�)r"O��qP��*b��@@v�H�T��`��"O愰'EE�06f,QĮ'��`�"OB�Iw�)5��B@�H;@�^��"Of1I��P�'�P���v�|i8�"O�r�L��|��x����:crn��6"O�h��ʄ5�01���:I_�y�"O�L����<��P�BLA�XG���"O�m��Q�����%�653��y1"O�M��ݏS,�T��0A!��"On�����rGD krn�>u�� �"O� $qC�I��}���ږo r>|�2"O��aI�T{�hҒ��K�&�#"OtmY�U4�<��ؒ9���y�"O��$��y� d�7�
�^� ���"O^�٦`�1%:@���JߦȚ�"ONܠ�O�v6����S?K�Dq�"O������(����U�{���8 "O�QK��1�n]q����D��"On!�E��@m����B=�"O��q*�'"8f%8J�
J��
 "O�Pc㪙-*S���$��#)�F"O���`
Sd��XP�R�,�Lĳ"O�ħ؏c'�y�@��>}B*�+T"O��G��F��%,1iHX�眬�y2���J�8�&o�n<:��Q"�y�I�_��[g�!l��ջ���y��)Tq��E:�V��A��y��H�~9��"��",��`�JV��y"+�>�P��T�*g�X�@�^��y���5T���c�J""��(wiB��y�/�|G�y�B�K��-Z<�y2,�
#)	��?��1�VDǛ�y�À5��Q��ؠG�|u:S�д�y�R�N�*hkc�	�I�
i���yB�?h�@�!È�@T{�	D5�y��R�	�ց)��V�f�z�S&�D�y�kB`���\�/��2Ɲ,�y�h�2�!3�g� z"�)��W.�y"���n�x���.s�,��q%��y2�%l��v���m����P���ybF�Md�L E-׮[)�ف��y�*�CT�#Q��aĜ�
1jɸ�y�/M�Ru�Y�W���`��ya�(��1h�z�>3������^�z0�؆�%���I@W]8Zs̆�b��<��[��@#�,]d!���:N�\��ȓO�tX�$��J���b�d�4['���ȓS���D"E�F����Vc�+$P����~� MU�+A�5�,��-Ĵ���qd�I���H�
+��SC�ݪd�ʝ��)�������(�:ܓ���Y�^M��x]RP�R�_`d�3��[=�Ѕȓ���g�՟Y-$��`	?VO܀�ȓfx *$,��$(��� 8᪁��1�^R��V-��0[%m��rȆȓ���IBޯ~�P�%�R|���ȓt���)G�^��� 8S��,|�f�ȓc���eLŴ)���r��Q.L���#����e�W_ްqE^�@X��<T�-�%W�*,�Q�	�'0߶i�ȓyJ<IG'C"N�����8�ȓ.�0ׁ�5W'~豬�d�L�ȓpȈ���ݮO�0��$ ڔ.TlՇȓW�^8#��;�I*��	p�>��ȓp�E(Wcň"o�!�bG�t������
a��� y���9�K�w�R��ȓ*���I��W���A�{�f�9D���!O�	L�-ˆJ�y.��06D��kUk�%*�ٓ��"MR�r�3D�s�nYJ��0زI7h�Wo%D��s���UF�h�E��ґ�-D�[ʋ�`�fĊը��Ӝ�P��9D��Q�ƃ�n9L9���1`Ә� �8D��������y3�, �e�aD*D�� ��r���+Y�8�0�� -�p�js"Ox�����)t�̕�d�Us׶XD"OB�
͢u�6�1�^�d"b"O	����OH���Y�Ă�"O�*�n9N��P��U��|�R"O,�b���5��uj�A��S� �"O�4zbk
�&]�T�`����"Opj�.�O��X*U��4�~@��"O 2�'��]O��9�iƎy��X�""O}4&��DP�$"4c�!%b�9"O�����)h[� ���Ň$��"O1�%�\9�vݪ��;?�@�v"O9(6�MuR�������&"O��8��&|����CE �6�꤀�"O� ��NV�j�H�CR�Ytb�q�"O����\��t���A��aY "Ot��em�	^�)0���H	Z�"O�ͳ�B��v욇b�>:R9yp"O��J�&G?\\�{� @ 21��"O����؉$��F��Q4nš1"OV�a��1�R�Z3��#O~xs"O�����(���#F�/7~h0"Oꠘ�ǿ!��S��3y4H��"O"��!�ǜ`(}Z��?b�@y��"O�(8�
J�
�����T�Pĥ�"O��#s��s�"\)��	�d��"O�p�Т�bk|9"(�H��h "O4�ѱ�ι*w��#wg�>7�	R�"O�}��狫1r�hh�K�� ��"O0�LA��n���_�:�jV"O m�2��;�ܡ�&
�9\�=a�"O���l�"�4�dϽO�va �"OZ�0�٦6Hj�ru�]�7�V%YT"O
�b�:�"!�@�X<f���0"O��[v��J���9�0-��"O\Q���	�d\Ȃk�:_�F�(G"O����՞��|��G�t���"O����bϪ7�F��J�$&����A"Oz���*�Ti�`��0B0�)W"O\D�ᯜ�#L��)�1c����"ON��"�^���0#���0Xt�AG"Or�y&�j�PZԡ�_��"Op���AƏO@�q׉�%:��e�'"OD`5d�j)2���$K�p$"O�p(�t�E�$�=��p"O�)�b��	0��×"Ԫ	z�P�"O̩�D�
6-�sSaWb".���"O��`��ٿM��5y�O�Dr��r"O�h��I���\)֡o����"O��r������V�G%UR����"O�l��X�
đ"��$7����"OX5*��֦v����g�;%�}�"Oh���.B�`�\)���J�E|�� "Ob!��E.l1�K�Ay�!��"Od����WWv��Y�h0�(%"O�)��M�p%*A�7�ɩ��;""O��yE�I4{�h@a��]�jpg"O���A��H	da��<s�j��t"On� W�
�U4��Zu����t��"O��1�D���y�7��_���3"O��V���=��M�&�2P����"O�ȣ�
���T@`��q<�F"O�� @���I�&l#k2y�""O�4�2�� >�<LI�J�4)a�EC�"O� ������`LD:4��`�IP"O��vN��D0�w�O��X�
C"O���Vl],�&����T�bդ)�D"O4D����ܙ�ӧ��x@�"OP�d$�%¤qA�B=z.%(�"Opm���C,h�����dM6z�hrp"O\`9C��'O<�;fC"���qD"OP��!�F��8t�7`G	roe*p"Ob�K���p��a�s��ɼ=õ"O�p�F��v!3⇒O�z=�R"O6�Z׊�m舼5a2&yz4��"OZ���j�y
�X�Ѩ����"O4�����Xq�c��m��A`�"O��a���p���CU�"VA� "O~� ���Y[�P�¢Y)A���"6"O`k%�6�\�r�^�A|Ƹ�""O�dK�fغ��=ӡ�!M�Y�B"O�!hqĕ&��£`҅1� ��"OH�q��;���ӎL�e���kd"Oh����	�P�`�<L��@�"Oj@�CM߅D}�w�ȁ+��4"OPa� @=9"Na{�ΐ��ѹ5"O�e�S���V��(�P�.� a��"OR�Sa���vQ&�ۗ兩C+�1z1"OzEY�LX�E�����A�����"ON�:`�Y�5��ջV�F�"O���EޥM�x[�-G����b"O�xcq�ˏ8ِt[ cΒP�lы�"O����g�''7N$bBƠH� 4#g"O�Px4có$dh��f�|��`�"O�|�ag� ��\�1�\�S�"O 3�∳/�l=X�
ӵeF%�$"O���u$��5��si�5UHa�D"OX�i��!"z�U0�,6�$�� "O4�����3l{^	�s
��E�9Җ"OΤ۲l_�`��#	A�Ro����"O�I�.�'��j�蜆�� �"OrJ��"��
3H�.QZ�"O��%�xT8IE�,Z�e!�"O��C��	3b��D��jҢ$q
���"O���"�,'4@QƩ¿Z]@�"O8�Sa�BD�l��.�?Y��4K�"O�e����8s����+�(C����"OȐ�G�''�F�7��?��9�`"O"1�FP�nh��b�F�B�"Oz8a�L*�n�" b��L�jW"O����`F\�i[b��O{�Y:d"OLiaR������}pl��"Od�aÇ-Y,�x&�::ilQh�"OJ *� �;H"�)����#TBP��"O쵈%DC�_��a!�Q,@�NX*C"OҘ���4����(Z�^BD "O�4ь�<`�0�g��L.��"O��Iaę�{d~�05&K�%��ڇ"O�i�$�-s��A����/|Г"Oе��k��|B�Y �P�Y u�"ONP�R�T�)�BՁB5*��:�"O��BR��$�:\CS�	����"O�Pj�X�%=`��Aߥ�NY�"O>1�s�D�
F�x�e �#{|��w"Oΐ�#Ulġ`���'`�%��"Oz  V E<L����6O�0KU���"Ou`��P#H��:����X=@�W"O�u�NX�=X|��P�D�$nXs�"O� J����V��hY�4��1"O@�g�[�@�vh2�ē+��;1"O��0O�̑S��=͎�"O��9R+�-R����e��@�F���"O�a�҈<U�)Q����)�"O�I8����I[t8�0�䍲v"OB��g�3$_"�:Ƣ�9W�L�"O��zw�ΊPˮb˟���x��"O�q����/�V���X(5�pQ�$"OR�P�� �a�r�b�v��"O6����@�^(����[X�1Z1"OI �'G4�V��|F�h"O����IH"8�TL�Ag�wP��!�"O����NЫ6� ��&�3]f��"OR��A���`����_�z��4�"O�4���ߨA�R�pw$
+�¬ d"O.�hC@�VƲȨ2ɇ;��6"Oؙ31�L<Wt��I�MY�X���"Oꨱ��L4�*=a7zؔ��E"O(D�B�G��Uf�u��0�"O�h�w�[����� �I:䬸G"O�����tK��s��+\3tQr�"O*%��+�1(D�JP�D{���"O���o�"��l�aE��&"O����/�5$�D�#l�P$�L "O�|��P�j��q+%	�D
��'"O��H�+=�!�bK�`�*p"Ol��u�ѱzPDժ̛=i���"O���"��#Ħl2�jC�5��xI�"O�pP���q���hK�|JL��"O"�B���P�
��#��j�l���"O�� ��װHWv��"��H�&�y�"OZ��T�(g��ĳ�d�<�h��"O�XRd��>�0�s�;Ȅ�["O�q�r���0f�̚��H�QerȂ"O���E�X�W��8�柃[
$J "O9P�_J�@�Z���,@�-�"O�Y���'p�iZ�,��g�.;�!�d�Ms��;S���6J���e�C�Yu!��'@PIfCY�6����2FO�5i!�ֆ�qbV�1��� Ug�Y !��V#x��-����~���E�b�!��E�09���-vF����ɑ!��R�}ʝ3��Z[��0��H!���X��e����gp��)���P�!�$Zy�9@g�P� �,�"/K�{�!�';�8l���56�t����!�DS�a�F��ޞc؊9�����Lr!�)S���aI-s��,r"oӎF�!�䌃$+��CУ߱E�B)�T�U"�!���O�>��E,{T��9��X%�!�$�A��{'�'YH.��!
�B�!�$�({�r���.H0Һ��p%��!���;#��Kv�E���p��-!�$D{��$Q�ǀ4	Ÿ��a� !�!�D��]�Qp�G�[����bG0S!�U=&�Nkׂ��y� �!DD!�$�i���qR�+N�8	�@�a$!�DN�g9
��Vi��jq��'�!�dh*�����z�D,a%/��c�!��R��\�̉0 "��d�k�!�$�f�X�P���5c5�|�T��%�!�7!{�!ɯ'44�V��7�!�]	~�|ى1n�<x@~�)#B��!�� z\����s�S>D����"O����,�w�d�
wn�(����"O����C`F
�렇%��P9�"O��2����]h� ƹ�Ф�"O���@
=x���C�
�^g^��B"O�(Z�̟>K�v{bD-r�\�f"O��i�5\����͇b�\�xq"O' �,T�tT��6��5j$"O~9�� @�
z��S�"�xA"O���
�ii�r���-����&"OH*uGR���<%�9i��s"O<h S�SV�H,�¨	�� q�"O����"o��=��I�(��tqG"O���H��LQveR�JU�`wNU�"O���3n��#>�P��[�o:�	�"O�D��C *B��[VĜR:���d"O��K���&�	ғ"^�Y5@�13"O%��(ğw�E���)����"O���F�?���� Z0}���F"OȄ�Y�fU��S��AKg"O��Q5@\�A�ܜ8�$�r�\��"O�]
GI��8��`�*�;B�"O>|Z���/F��9ei�7~Ӥ��"Op}S��]ULH�r�^'[&��A"Oʕ��B� ˂	�"�$�&"OD��gk�v�ީ3sV��48{%"O���'�;R�Y�A��\�04K�"O6l�1DB!��1��E��'��I�6"O�P ���R�8�q$	�2x�"O����0�M��D@ {�Ҩ��"O4,Aw�ӿA>L
�ep��s�"O̐x0'��Z%��q$�<�@١"O����2MX��7B>$���"OĘ�C)��q]���¨�\B"Oj���nt�<���JHXh�"O(�Tٲu����AV�&:���"O���$`\]{��CO� �u)2"O�܀����Uъ|���pu���"O�k ��dx5���j�5b"O�3r��9o �]xB�W,��b"O�0K�l�1do�(Ksᑩu	Π��"OH܁cb[�
b�y�`��L��)��"O,��@�n�>h3g���(���"O�$����^��ȡ�m�8B�ܽ��"O��#��	#���C��
0"i�F"O�q��*,@8<ZQ�#�D��"O*̉w��)�H-�J���"O$J���1Q���5"�E�Fu�x"[���<�~:��=����  �L������f�<�RB�z m�1�ֱ/��M+$g�_�<�U*� "��僑�����)V�<I�a��.lL��ǉ+��d+��U�<����*�da׋�0�"��4��T�<i'@�3]Z���Mv>�Ä�=T��i6��[5qՉ�c�v�a_<!���6P�U����*|�.��R��\#!��ԧu���
t�E����vAW"U!��_5g��AwH�=zL;��?!��'z��h[��/v���Wk�!��F��	ےEX���;v���!�䂂;�<Q�AGت�~x�IPA�!�$�4k�����ȱn�NE��GV�s�!�$�4h����I�F��`8����!��Q��%/�,ovT�s�&0�l���� ��2D��T��=�e)D(H�J}(C�'���>z�1�� �)���@��W�X0		�'�d��_?�~0)��$VP
xˋ{��O
�}��hl� 3FY�pGLtZ�耠*� ��P}.�YыP�KZH �Q!�3��9�ȓYz&ؐpJX�x�%�`k�+Jޔ��Vmb1��nä!�p�҃J�T�ȓ���ڑ	�M�s�ܮ"�X���`�&� �	+d�I��͒�@�ȓ��d��a�z��uB�5Kb.]��	\�$� ^�2e���.�ahQ,ãJ1!�D��$��r�/����7��}-!�d��z^���3�[8L���B�N�}Ҝ��%�S)pTL���#�Ch!C�#%D�h*F�[�~tp�'m�`���%D�T���68��2&Ԁ�VQ���a��Cተ|	�Eb�^�*���KmҪwTB�I5I��L�6�/.nڵY@��8�C䉪CT�P��͡L�f��D��/N"C�	�r<� ��4wL	6��<D��B䉏!BB퉆��~��y`ELWMU�6M'�S��M�AKJ*W�B�b���S^L�2�
XQ�<9\�J�R+	�4)�$2���N�<���o�����ƍ6_�f��fMJ�<�u�v�� 1�P5�
�@�G�<Q��M\�[�"�u��Y�Oj�<��,�
�T���^�̤0/M��D�<	 o�q\ƕi& Q�Z
��T�ğ �!��Z����y�k��3ؼ͢S��~�|b��L��Θ�>m���YQ�TY�L>�yB��8ZT\J���;���hc�.�y�
4^XA�  �2�6 ����y�ă�	6�M�0 ���d�8�y�LE&rB�h5�W�(�Aw��y2툀x�:�
���J{ m�G
��y" <uh�aqf�F1�%�v@���y���`�<�F��'0t8���;�y�N �9�&���Φ3�� ���D�yǘcѶ9���Y:[}�5	pgݖ�y�N�L�\��C܇W�j�Sp�Y��yB
�,��a�‴M���Ԍ��yR�@��`�`E�(1WI��ʜ��y�E��8�T��2���<8
��#���y�D�5n5ڸ`�&԰�����	�y"���<�PĒ7S�>�˲�?�yҠ�1$FƄ���H�Qаn��yB�Y�L�}:��&)�[� ���y��"ytPU�ui��4���N��y�Ŝ?{c���ce����צ_��yrG:A���"�K��~����F�V�yCs�Z�2@,��I�M+�ʖ�y2
�(�X4`��2tT8�'��y��ϡ�����$1��*�@���yr�b�JuX�!1�6�*Ѡ�#�y��]92��b4����q�W�y������
0� �J4�u���y¨	�r٦9*��J�fW,"r��ybE��]K��;Y{hi�A��7�ybG�O�䀀�H}� �����yB��{�� S�����BN��yb�H�&x.Y�S��p
�)K����yR��O�4��bM�l��Iz��H�y���9"�p�6`��+�%���y�c��A^��i��F�nT��;U�8�y
� ���5,�9j�k�̧I��a��"O ��f�5�� �S�����y�*O��Thö��t#�悅/�����'=8�*q�R?UUD�rN_%�H�'�jy�g)���䂫!���a�'�Z�[uJ�)� #�-��=�x �'.��q�*�: �%�^)~�����'���@#�ܦk^��^4^y�UI�'�Z�Rf.�8U&�)�����	��m�,)S��F,'Mb��"%�]<h���&�P��=F�A���۴D�]�ȓ`�Ī���9���+�Ă:E�5�ȓ��l�7�Ĉ~J2 [���m�؁�ȓ.�L� F$*h��I**���l��xp���`��@[�K�#���ȓ��u�
3Ԃ�ʴ��#N:؇ȓ.�d��2��?3�lIu��*I70��ȓC�t��Q�K�8t�*��.t��)��L�d��$N��أ���(y�r��ȓQp�+v��,k(L�b@
��{jV��ȓA=:d���-	b�N��T�Q�ȓQB��Xw��O0B\ф�O"$a�ȓV9�Aɓ��

��m�Q>B���(�P�:�.�F��Ԓ6	�F�Ą�t��a`���0xAf�츄ȓO�����Z5y4��q|,��ȓ����0/�IkJ�pȞ�9�n���s|e���<$�M��@�/���ȓ &q��ۣo^zc��.P9�ȓrX<�R̟�~`���	�7��]�D0�Νx��]b�FF.^#����*@��"�)�hJ��֬8K���ȓ,f~Y[#�J�洁�Ș�8�PU��ZY P����9c��7��i�ȓ2,����[%(h��f�`����ȓ���H��oa")76�LH�ň�b�<y�E6]�\���6 J���5�Y�<)�N��!R��7��봁�y�<�7�� C�6�X  V�L3e�&�<�2J��U0�+E��0^�R2I�d�<q"�	�N��,Ђ.Uе��x�<���A*��	ֵ�k=l*�)P�<�d�L
~��S�3t�z�)4��g�<预>N�	��C��$)LYdI�o�<��'V�!���"�b�)#\����j�<A��ڭ-Q�`����N0�!�a���<ag��;zv�3�49�xG�J�<A�D�2{[�y��؎'Ȥ��Bi�w�<�v��w�`��a5�IS���N�<�DQl D%�B8D��P�`n�M�<93���!��4d�ƈ����m�<	f����Y�)S�y �K��f�<�u��� I�����+:?j��ˍx�<����
���0E��n��Wn��<A�X8h*� iOs�a�T��|�<� Q�uq2JU=f^zc�A�<)�`�Q��Uqv���V� �/�s�<9�X�-S�4���*9
�90oMr�<Aҹr�y�&�X�X0ţ�7B�!�ʌ*�q�b�U�d�^в��<�!�$��p�N��@���Nۈ@�W�-:�!�$	.]�x�φ���AA��S��!� *w�d�R�OM>Ӏ�y�AL��!�Ԡ��=��
�^z��GK�!�� n䈱n��HX��ޙ+m��S�"O��Y'J�)]*���
�3�.	��"O�0���Xl�����B84P���"O�)ɣ�ML��w�:Tm:�"O򬹣c�_�3�˛�~���"O((�"�FK�f��l��g� B3"O$L�3G\��y�-ͷj؎=ʗ"O�\��I?&���*V�T�U�� �"O���"���J��8&U�"O6��6ͣ�FL��it��"O*a2�R-(o|u�R�H 3��833"Of�N�/\�QG��
����"Ot�xv�H�ue��`@ǟ�%n*虧"Oj�����%jlX���W��,�f"O�-9r�=<���Aɐ�L�ݻT"O�ᯔ�s��Mh�ِ7A8]5�'�8�;s�	'�����]�xk�8��BӋ5Z
�P���O�8Ei�'���s�E�
����u\d
�'�vmHEoɈl�Xq8GFZ�ZP
�'~�)U�oCb���!�]�I��'I�%2��A� �~�R�3Qǒ(J�'L*b�P1���ɂL	J�����'i���E��Z�B�G:9��ݹ�'s\��� /=����-V�>��%��'���7�z��{��ܲ�����'�ʍ�pk�m������ $�z�H�'p,�Cr���]s�Y�q$�
�"O���P�bӆ0�懘
�m� "O$ݒ���V�z�h�f��5���´"O��KC���]�M!'\�*M���"OH )#$�
e ����E��(�>M��"OH��ʅ�_�*��v$�2t�R�"O�����ˈ{�ڰ�W��3]�H@:1"O6!�eF�1����@�ʽO��6. D�����R= <��"n	��HU+�$<D�d�4��wPb�	�P�K�=��;D��y҃�@���`
L�V�@�B7D����1^���d��(c�x��j#D������:'��11��7/�F�{�!D�8�Ba�z��Ĉd8s=Ne�r� D��A��8)tx����~���/=D�t��B���81��.T�}��@(�f>D�lY�ĄlʴuC/!TɈ��"J!D���t`�5a8UDK�MT��p�(D���E��,����j�a�h0� 3D���G��pڑ�B,�%C��g/D���F�Xr���([�EveI%A!D���!�D��H9bd� ׌�V�>D�4:j�px��@1�[$ y
�!� =D��vN��$�P����E,u�2 �� ;D���	F�"Y@�8���7&��c
8D���Gɿ�	h�e,V���SI*D�H�� ٬:� Y�8B ��jp�/D�ؚ�e��^2n�����&M]��3%,D���#b\0��Ĺ�"ڱlC��d� D���&BؖS�Y;�/č%yHA8�a3D��sH[0|��C�j��}�:�Qr�7D���iϽ|�J�����1)<��Ǫ3D�@��B[�a���&S*RT�$2D��t�@�:\�k����qz�Ƞ�1D�(k�C&�<4h1嗌f���'."���d����j�v�b�eBި�ڵ�J��,�<ѕ�ʈ��].q��K�?aI ͘�^8��J��� i8��V䌿�ƹ���Mm(<I��B�<W�IfᕸH0��$o\9v*�����Q���Ȧ{���kP��(��<��j���d����� 2��A>����!�Z#/T0lpO�)k���H9cG��m[n4�L�f��=rѬ�25|����F�m�Z�C��Ӟ�b&�Oڲ�X�O��%K�"ӪtC��� K$����'G�M�&J��@t�	�3�t� E���]��1h�*��By8 �Ҡ�W��`�u�i^y��N�EY�����",N� 9�yh'��k�h XrM�,8�OX�xd�_~����0�M��N�ם���!��B�R� 5$\�-��"Ц��l��
uӀ��*O���WcM�U�f�
���ѨZ�Vx�'�T�(l��a%*rK���)�OHѳ2A�*Yr�RG�Q(X�BH�爕=*d��aE��M�1La���B&Ɩ4�ȳ�k���P��&ʈ,`j|i �I<z�t��$�S؀��򩊐izd�#��S�?��	9u�I�)���W<w�:)�C���M�1�Ҕ"����7�'Ev,q[2
Z��꤉r�-	�4X��	���T��`X�ز@L_�P�R4�'��ɒl�H%6��*�{5���c�A1;˛6iE�WB���5}L90v�ػ�Np`Yw�|ɛ���P	���NC�W���P��JC��3���Sհ�%�Xs7��
<��us��'�m*3�4u2��S67�u��'�����OzW���3�R�~5nD���+���w%^(:�"����G���"!��'7���1%X�RLb�W:33"����~�"I�؍y����?݈2I�,B+,�4�ܚ����X(� �E���D�y�!ӭ�rt���Y��ad)�U4Ն�	=^����N�� m33�!5!F���<��	�{��y��_�b��yH�B��W������Q�&��V�R�;����d��wU�a�W��%',C�I�0���f�_�et��z/ѫQ���Z��^�or��CG�s��ju���5��&��jWҼ�Wc؊{�A�E�M�p��q ���w�<�u�ʹ[H���t!{�0���Z/[봼�E$�I����O�����e���XO���$aK������"
Q�F��c�+���	�So����E=�~d34�	e���U�E p�<���-g� �@O,ZkD(R�+S;���$�&1,�Y`o�n����
aj�e����d��vX|0#��S���G��5H�ص9�%�20�8�iA�S1�܈ ��Q��M;��|�ayZ�p��͋f�O8sAbʹOQ"�)k�8#�.�ŭԁt+�d����� ����3Y�V9��̷IU*�1��<�t��S܅pcmS�Q����?|L~�Pb�U�.ߺO���$�*S[�}��U����oIH.��۷
$��"˝7i.,xᓣF(�,M"U��3.��I��BB8;f6-^%K��0fֺl�Dh�b��	Q�'�<+��r4CÎ8ɼ�b�@�`X�S 5; ��L�(S�4�H�t> ��i�A+EJ�f�l�ƯO�K9:%*ED�cV���lb����4�R QBNA F�'���9��P�	�D�C�	M��H�#��%��)��4��hɔ�	&};��mڢd6�aF�-�j��O��>.�&�
(o�)c0L��j,��a]��<A��(I*�pʡC�O�D9#�39j���.�v ��ze��8�8pc�F��M���D�[�x��2���nnؠ�'�Nԛ5J��*t�Y�f ͈����8���Z��H<�@�_���HV�?)���-|"��'of�!��A�aH�U#3`͠>�h
E�߂X6|�s 	�52���!�?�E�G>��I M�?�l
�{R,�^�2)�F��&�nݸ���3�"d���'�!�׏=}ưkSl��]�*�� ��uWcΞ3�^c���	tC_?�V,dV�(d�mP��A4���S��@Cd��� 3�����߾|�)��ɭA�|1#�
I���;Q�Q�'Ӑ�:�� �6��l>!�js[�X���F2O�xfH�YFr��pÉ�QخE���'Gv�� c��P��䛀2��.�=Y{R�Y!��.	&� �Ё�(������B�0��T 1GX�|�f��.,Ѹ�bfh29Hg�f̓fj61XG�<�d��6���M�&s��!�2ĸ#*�*C�yz������[�P!�VI�4�ڒ�:z}L�E���%h^���~r�B��U%�@�0fȢ5mM�*a!���P|�ᒒ!��P�)��؎-S!�G=@U��HS,��;<e*���23!�$�I��h teňo�$m�G�|9!��_9�y����/*�(�AE�'!���k��%R��u��s3DT	o!��@�Z���� �0I"����!�Y�α+�������ɲTp!��3W�R�R2nL�#d�@X��	_h!�
k*H豴�Ք8L;r���!�DKH�D���{j�yr*[p!��""*� ����4X�{�jE *�!�D+F'��s�O�� �n�k2)V#!��
0���7�T�p�~"C���<�!�$�#^��
B��
���BӢ��!�D�FV��2�*D=M0�,�g�v6!��:Jv���-?ZXV�gr!���-!�
Hi����2���3"O�]pf��34���R���2�"Ov�rʋdѺ�x	y�l��"O6e�%~4B��_,+$I"O��1��U��i{��e�Ð"O� VȂU���U����*['`~�d��"O�D�u�7|�TY� _�FSFq�"O�P���\�� {%�3?E<e�a"O��X�IT-�����^2����"O,,�q��I&�LzdK��\��"OP���!Y�3�V�B#�$B��q;�"O�h��	**���G�9�"OT����V-s�hu�eO�  Ny��"O�
Mn�B4cđ��QSS/D;m!�6R;E�aGK�n��pS1��"r!�d�
���sӴ�,��m!��֏|Ӽ�X ��K�j4���3�!��Q�~Y8�v �d�"̺��6-j!�R0|-�$�R&�?�@�IvÀ�MI!��?�����I�E#�ɹ��H�B�!���Cl��C�g,
`Y��S�!򄛥fqH��]:)�5�h �!�Da�>�AECޛhͰ��!�!��P2)��h�oΥ�t�?y�!�
�I�a1�Ŋ�^<|ò��(�!�$H�{���`�܀1����ߑZ�!�+R���T��,5n��Bo�v�!��U<9�X��934��3��)�!�D�#��HH���W� uar��/�!��H�z���S�X5�����!�D��:nH�f��	r`���
{�!�ߕ�A�.�?�Z����M�!����.�����ȋ-}�!�G�/��@�`�ɨo�葹�i"�!�?^�B��̈)Ƙ�XRS�|�!��o�:H���L�=/���>+!�ڟa�1��EԪ,�QTo!�!��G3p�~�!��1X�5т�9@c!� �����6_������-x!�dL�+�)�O���w#C�$X!��8&Y��0$��-���V���!�"&(r����S
zM��^~'!�DY�qF��c�˅$����!� !��WsA��
�*��m t��P!B��!�D "H9j�Łub��s�� �!�]�RC�8�ₓ�n�f̓���Z�!�d�.�M�%Aڎ\�5�SC[ t�!�,8�ғÀ!�
�g�
�!�D� ���;P�:/��2A`��L�!�d��yE� ��j�[���+5Y*G�!��n�`i0���Rժ��KV�R�!�X=S�M��M1?�-�6KB={�!�$E�y&꨸��O���h�2�PyB�TL"=C� >BV�ƙ:�y"�|����ƥ��GPr�Bӭƻ�yrH̅c�AK[E�0�놋&#�B�I#iL a#��T@�V	x�A�n�B��e�v���i�8�>}��KzB�5+�paAɛ��ԔC3	��@� B�RƜ�B@Z;~��S�`L8,�DC䉴n�����.��AI4` @�M�-j^C�ɱ:1*s'H�l�v�'�K�
$C�Ɉ7zʼ��ɛ�|�8l@C�8��c�HȮuC��`�呲BZC�ɡX���9u�
1H:HL��o��C䉯0�v|���J:�9��׵)�*B�� &8�<�'ꖌ= �9G�Q�ErB�IFb��r3�N���WHȑ/�JB�ɝզ�A� #��9�A�?�
B�)� ����@Ur%���̴<����0"O@0�bM��$�
�s��� ���"OX$���S\��(!�>*��R"O�� O�H�))6m�Bjl3d"OP�X %�C���c��r&؄�`"O؝ŉ�%+���,
�^�^t�"ODp"S
��&�%�*�L��A"O^���Ĝ�)��`i^4K�)�*O�DYEl��9H�4��A�#�'�pp��j,u��s�e�B%�
�'͔��iƜTJ��K<XLj�
�'�:<B��]�\�H���#�^9�m�	�'�X3g	?�B- v Q���	�'�vM[�/Ir�|u��O�U�x)3�'a�勱�� ?²УጘO,�[�'�J	�炱@�D��2��>;���'�}3�aƱj�zX��>+*�z�'�܉��,TMJT���P�]��'���eZ'8"I�MŪP<\K
�'����� ��l��૛?O- �a
�'q}1&��{zH��Èx�@0�'����quN@���w� !�'�=���ݼyk�,�2 \�[���'@~���^�h�D� ��Ӑ���'�\�����m�n sb�i�T�R
�'Ԙ@ �V�&w��ZscO f4�@	�'s��h0�
*q|y겈@Q<lAA	�'�n=WdC�jFP���H�4J�Jq��'=��y����Z�,�.C�0�0	�'�m��'��(r`�Z4(>4���'D�-�Ӣ�a3\)@��ҀY���h�'�0�����m�Ri�!.��_A01��'J������P�:��1ꃢQ��x+�'8x}��J�'�<a@�D�Kh�@	�'/�i�9��]��ܘ~l�iZ�+&D�Pa�"��/TY�P�4Q�Y���$D�xp!(�s�|���Y�f�HL�e.D�pz�̔4"�	Y�│+� Kw�0D���A�RFz4�;V�1Z!�$D�h�R	����:tדC�hU��n/D���&��]�9�Vi�;e�^��� +D�h��Ǒ�#��L{��F�{	<��u�&D��a\&8�U�uH��ux���'D� ذ�޾_�D�8s���4��D���"D�|$FDH��
Q"Z��<0�i#D�`�Ƕ��;��qqn���'4D��3$E�jf%+r��7iC�2D�$�M��X�`\Hd�?�aðG-D�0r�@�yۮ e��nUu+��+D����$Q ?˦	�@	M�X!�,QÄ:D�\�4�F��<)��	F:�<���8D�8��S<\G҉���a�O6D�THF���*�Ĺk$ R.PB<X3��+D�dY�_+yy�LX/ 7Ԣ�6A4D������<� ��#��"~NH��.5D�����Cl~�x�9^�p�9�7D�h
'�/;���%N�8BryW�5D�xi�)�=]�t�)@(�4YJp12D�8x��E#F��!5(�*C��@1�<D���1H� ���j׸C3�ŊL8D�|H$Wz�@�A�&׈��d�*D�T8!
]��r��L�*K��W�>D�|i�ІPt�(��<a5!{e?D�8���_H�8钖��(���"6�+D�� ����=iSLD�3a��"��H$�|"!�#�����	96H|sV�0Z�Fʔ�"c�4J�J�
��	9F
T�؟.M�pgF|1b��U�i�MQ�ƫ��)��1���q*�2�n���� 4�� ��î���(d���ٟZ|�(� �j�B�Bv�O}����� �����!hF�-{ȃ�qP� !O�1�qI5dGT0����#w�9r�>#�H{6d2h$jyr2�� 0r���iӂ�p��OF���Ol�A3ճ^5��Ȃf�OM�!*��'�b��1EL4p��L�	�:n�}��A�r��T�ǭ"`2v|�%A�^d�
׼i��	��ǍJ�,�ቐ��kd&͙=�f��`)	4`*Oٸ�ASn�@ �c�Ys�Q�[(��2�,��,L��!$W.G"�U��W2$Ѫ���@v���1n�
	l�xxs� 6�",���П��fʆ�0�`{���1o�,iӎ��o�|h[s��6�<�ݻG�H	��f��`u~�.M���C≵P�}s���;�n����  <�9� [4Q�zd�#��#}�>s����!ڨI?��Q�'M�-` 	L3ݦ�p��#�J�؄�[%
��Tx�l�mX����	�Orщ��'慃��81�Q��X��l$��"C�H��f�4�t�bXG�ZpHvI��tj�Aa��I�L&@�8�-]:\m���۸.!O� ��6r[H,����s�KP���	Ģ>�F�*�ʋ	H���E�HC�q�����P����A�n\���	)L���J�it�Y3�烊�R��ᴟL�o�?T���O���c� �8�)�#AZ.�n��,���&�rTc��!򄓕8>�MBd*r�" @�]x8Q�ã_���Dсx��вsi���	"�n������Q%/����ݡ7�^�w}cw"O0!�d�Y/_~�Qv�\P�i�
��M����%�>��5�gyrE �*�����H�{8�Yz����yr�1'96�#�5i���rژI�[���jX��W~�|�1
��#�p�P	��Q扄�I�$� |R�m��{ �$�-e�0)-Q�Ul���m۞q�!���;u�(��2�ĝ&W ���
A��Cg����DI/\H0"�G];��	\�� ���Э��K�9%H���E��-=����%�'I��C�,<��Dռ\�F�+��N-�ѨA��3�IE�G��r�fh!3�� �L���?���L@<@�}z�Y)Z<�����$�$�3P�v\	!�	�?ᡧ�=L(�-e��R��e*ف�>�yG �q��q��"���X0O��r
�AWj�q�@�K�f`������*��h(W큦��Ot\��"	^I4��V �Y��,;�Ň� F7m	�u��2'���@u,�;��	1��98B�I�!Ȯ,a��ڈ��q��� }�j�K Q����rc��yr'�"pɛ$J7�2�i><J�kt�Y�#@��VMQ�N�>���ՀJh!���'��a�玘�6�����c߾�pM)"�DQC'T22|n���2���i�N�����p���QA^�<!"��X%�)� D*Βh��� r�V9���iB�fF2�9 p��c�Һ�0��98,�^1ܖ$k�lG�H��i0V�W���-ɲg�t��$ <����S�l� ��H���c��O���VI�-k���Ƞ+�����ؓ�ؙn��[!#16��;w�NTKE�ʳw�>T����J(�����~�{��B�:��G!��t`c闺D���)D�`�qPK��5�t�C�4>�dq�7
n�Q쩈P���Y�Gl�'pf���$�r�&���@���XW�1;���C�D���͆� �Jţ5%_�d(D��:�`�B�'Y����^��ѻ�cתc~�X��y�#W�b|�\�'l`<kg��O�2�2T�  �'W�w��iڵN���Ӊ��Px�"����ٸ�%Ҿ̴�S@���O3u�@�~��!���tܺ�5�ƕ17�SB�<y���/(u@�e@�5�$O�Q�<��+�5BXkG��(Cd�C��A�<�V�׶���O_�>���d�d�<��G?J���fJ�p�s7cFI�<��H�>?�|���
��I�؜ʐ@�E�< �ڞ=��C7��-��;�)^�<vNÞmuj`[���HR� ��K�_�<�V@E��R9`u	X#l�h�)��C}�<�F囗^.��Y`i���	�B�A�<���M&.iZUAӛ&#,5p*�V�<�F��07��r ��(�| ЦIV�<��"�	X�$%��J�>hj��B�V�<!���S#�<�`��-\���A�F�<�/�>�V���*o5��*g~�<ɡQB�I�f^+4���iԦ�u�<��a�4>PvܻэF"~Ǩ����v�<���RI�DA1.���(6�
r�<� �􀓥��^Pqˁ&��(g"O~�;p
(�x�k7j	j2�L�E"Oܼ��J�'���B+�S�@�"Od�I��މ��CT%�3���p"Of ������c�4C�"O��9w��'�е��̀Ƣ�á"Or�d)�!�I
��ڹVB��S1"OxAbe�+xlT�pо�Le�"O^P�t�� ]dN�n��ȸ�)P"Od�����@��	WB�$p��e��"O�X1R��:p�Bg����L8�"OxN�eO>|��H��,���"OFT��
ˢv���C��=W�Z��&"Ot�#�
^�i�zq��%�Vm� "O`�+��M3z%�y#�R��pyU"OV�2�)�83Jy������u�4"O����H�/i�����ԺE�e�7"O�u�-̙n���Y�V�
e*"Oġ�ÑF��d���ա*��lQ2"O�AB���$/^����]pCw"O�xC�,�_�@�y ��Q��"O�4+6HK;jf�tLp����B"Ov@2T�^4Ddqm�0�����"OĘ���0Pj�e�`-	��P�5"O��X����ry�=H
�[��,�"OdM:��ߓ.!�mȑ�ȝGr8��"OJ��D��4�l�� - v`��"OX����<A(ٱ�o�4|,z"O�XIm��	b�Ы�(�gT��"O�Q���	
6)�6�V1>@I�"Om�� �X[R%A�Ȅ*.tS�"O��!F�`m ���g�4�Ɲ�!"OJ���l�B{�X
�݌7N����"O��P����ъz�(Wa�`�K�"OlYÓM�)}b���d��ݒ�� "O���QZ�%�H衷��E���1"O��{��@�Q��\�X�b"O>�`�m�E�Rm#E)�,�i�"OЕ;��A-!�`$��5����P"O��s����"��`s ��"Ox���
�a��5��"�>x��ɻ�"O���2�MR�}�PC�-mĚ�S�"O��pwAE2*��jw�ǭ*�����"O����m��W�� �B����"O�AK�X+ ���K(b�0��V"OX�r֠F�uk�d��@��
�|��"O���6n��z��p�Uۍ^��R�"O�@"Ec�/\R\���Q��(�"Oj8�1�IIi�`�WK^�r4iy�"O�Y�/�-_}�eDX�M��� �'�4	�eҐ� ��((2M�'�T�[���1A�<�J�@Q#D�L�c�'�f��&�F(�U`ajзl���'� :棕q��ܰP�ׄYP�Y��'�D����˫;<t�a�K1HC�Ip�n-Ӏ(+�2�c�lC:�BC�����\#n	2Y'�$�B�ۤ�Z�-�/*|1�m��`.C�ɇO���� ��*��4@څQ��C�	@�@Iz���3���Z���n��C����|*dI7;��t(�cY{��C�8B�@P��7$w��[��5��C�	w�"� �.3[�th�F
R��C䉣V��2kI�w�m�F��}�C�)� F �dV�a��H��L�z^�!k�"O��"*C�O������?51ڤ"Oj���E^�
4�|����=��:�"O!��1xU�� ��rZ.%"*O� ��ᅛ&�tZ�)W�J:���'+*Dc��^%k
�h���/B.���'�@� PKU��$d��Y<���'jrc��Þ|�J0�F�)"y��'���3(�
���h!%�ZE.���'r�h+D���;1V� 5��r ��
�'���SՈ�f�"�"��
iFA�'���zP�Q2X�m���AP�Q�'�ܫS��B��i�D^�I_>���'��
�ˏ�|P�J���S>����',�գDJϠu�(���!LAx	��'�U�@-S�VĵP��$;�XiK�'���p���\�b8��l ܬ��'Yt<�"	ډ7���օ �w5��*�':�dr'�z��(VL�)y$*�p�'�B	"�(
�\}�h˝瞑�
�'W6ѹ����@y���ӡ���B	�'���	)��b�����/{Kv)k	�'-�p�B�l��Y"����iE���'GlaGM�C-(�U�i��U��T(�1�7L�4�C��ҥ~���K`�	K������4� @����<�$C�73:�y@A��c�d]�������ԹM�4eS��Ύx��y�>���g��ħ=H\�P5��LrU[#�	jN�'�ࢦf.���|rre�S��$y��6����j�P�ʩb4�dl��L��%�ܪFR^UH��O��-���ԤV Y��J�T`ʳ院�NI"q�@U�bt��蟈�įK�	�咦��j�����L��0� ��i�����0|ZV@�C��h�sc��_7���q��e�-9�+�f?�,�{nd��)V X������vH����%S�F�`nZ���]��.	���`B¨8�LȲ�g��9ᶂ-t��x���� ,*��yF�ߓn*��JW;Oa�t��YA^*�ňD�\ � G�8h�%��%?Ia�q�a��ח;��4�g���|u�gƎ��yDU�)g�@���U��<(��ڮ�y�O�r �Qزc(h���#��y�DB�-T�$��ι
�^�����y��<rT�!�܏x�~��!����y�C��F8��8E�6��+����9�S�O����@I@23d!@:[_|���'3���i��B�$�$�G��
q��'�4	�)�@[@@
�,+�BJ�'Fl�)T��p����eG����0�'=��𧩌�e����C�3�!��'k�q"$a�Q��a1'�!�5�'�f�����%�	� �
�2��Q�'�&e��n^2hĨ�:U�'��y�'����υM$ƈ�G���r�'��x�L͛-t�]�1O�%<i�'��	����11^:`)��Z� ]���'�v=���633fq�dK��'��� ��'����7o �PBR��	�'�,��*�t�zw�W�0��	�'�Ȁ#��7Tf@�SmL)1�΁�	�'��t�4�K�P!m��툩q�����'9����a6�2�11�ɐV�Z���'��A1�J`y^ ����T�V���'��i!4o$tzJ�0 	F؎���'��v��$;��U�'�ѧDo��P�'|d] ���6+� �C�+����'��I3��cIf\`u+�3�X)�
�'�vup��2.�R�2������  �!ਈ�/3艻�c�]DF%k"O�,Ҕ�J����QC� 53����"O< �HǂlX���Ѡը[)��`�"OX�ѣ�k*xx����yY�"O�d9'�ܚw�"�B�,A���"O��U͞[�<1뀱5����1"ONE�5� �xT	ny�I
F"O����a�v�PH$ȅ%=��ȃ�"OY�bN�-M;�511��&S�H,�"OH��˒�d+��`��\���D*"O���s*V$9ܼ��D�I�X�ʉ`"O�Xyӆ@�yJ���B?�N�J�"On ���#r������r�6�Y"O�Ɂ��sNN(@�H�ݰ��7"O��3-�3@��#��I�y��\��"Oj�r	F��q/� h��`�&"Of�H��ʑ33���.�=X{m�4"O�p�'/]�]^�m�R��J B"O�]"��� ��A��l�8yg2;�"O����?�V����6L93"ObD�c�� vµ���ֵ@�] "O6"��Y�{B�e��AI�qr|w"Oz�hlZRȢ!�e@-k��k�"O$=@�.#�8r��  "�Y"O�z`��{�贫�̀�g�J���"O��ѣ.��3gf@����"OhJe!Z$tr��c��!�hq�"Oؕ���#5�IL�!���"O��y���8XY(P�P��2����"ON�9'�K�V��,`R&�<N�=�"O� ����gr��j�'m��k��!��~�����nhQ���ѦtN��ȓ[��yA傆0���S!�&�����_�����"�����S��p��A0��%'_:P�ER���#���`�Zg቉V���Q�i��p�x��A2����J+V�v聳I�K.0���gl�ٰ��%g>�cg̔GI���h�:�Έ�G�VA�b���I��w���e�*fId1"§�:&U�5��N�n�3� �&a�2ɢ���[����Q��b�Q���I�o�<y�ȓ]=�� ȗBa�	q�$V�9����ȓJ��;�&��N����^�@��]�ep��a�Ȁ�]�j��a��FVH�%(�>`�X8�64�n,�ȓ|B)b�K�&�<�IU��X�D5��W�f�A.N�f�)�6?�4Y����L�x.Ե���0n��ȇ�b���Sn�?Ch�ԈW�cy�]�ȓP�;3��&�h9j�֧)A^L�ȓf��P��F�a��t��5�T�ȓXzx�h�J+���a(U������!X�Ur�d�u����~�L��8<`#uċh�*j۴
�j���\����6$ρg4M�$%�J�ꁆȓVSh r"U� �V���N�V�8��ȓnRj�KrEٺ�8���Z �ȓo�,Y�s��9ǒ�ˁ��>n�H���]���֢H�j�����lɽP�ڼ�ȓ?�e���g��)�ֳ\��T�ȓQT��!�J�n���S�^P��K�t(�pEͷW��1 �!H�$E�x�ȓRc��(�N�;$`���^�jх�S�? ���gdkw�2�P�tTD͙�"O>�I#��YpwG|8L0��"O�p��#�xtk0���{1ҁa�"O�hTNM���hD�SN`s"O��a��Ϡ#����C�=��e��"Ont�0 �D8� "ƒD����5"O��[4n��"�F�P�H�4u &"Ott�K�/F����ʛ�h,˦"O�����[:^n*�	M�@�=��"O�M�ᇛ�A��|3���
�^�� "O�!��C1V[�X�H�/g�ݸB"Ohy;Rc�h@L���FQ� af��"O�H4�I�_�F*�N�=`.A"Of�ڣ��Rb.k��@lG.i�%"OX;�N0��- ӄY��B"O�]�2(]��Тd֣A�4�
�"O��˱�N,���!����,��7"O�Y�Q��֤�b%�$�L��"O�����Q�9�ҡ�� �X��"O��1Pc̦.�lkAT%7iNA��"OZ ��ݸ0�����'RKf�xV"O���jU11����T/��A0�x�"O�h�p�02�&L�#ɖ$<8�&"O:uP��o�m�.	�x�(�"O�;f
 �/��]�c�Go�rt"�"Oޭ�`LM7}�lC�JE?��m 5"Oeڐ!_	dzi�`i��B�x�w"Oj�:R(W&k�f�H�(G�AhV�!d"OFYzE�-t�d�g�;DQ��G"O���r�F=zh�"lG#=ܫV"OX�� ��*\cP�5� C|I"O���GN�$���u(�|�8"O��J��H(j �c�οs��%��"O��i���+v�XE�N���AW"O��gä6K��ڠ,;�.�#"OHXs�h]=^:���#iۿ��xR"O4L�a��(���Ć\�F�s�"O^�)�/�#$�,U��/�2B��ؑ�"OJI�1�B6^INܑ�m=!��;C"OD�j�e��s�f|{�L�G|�$�"OL�R5n��0� ��3|��bW"O�԰�8l$ ��B!a�.��"O<�C�+Ux�a����<F�D�z$"O����T>� �ҥ˕�yo�,+�"Od *��R�6A��´PnA9�"O��a�����8�R��٩qV�E��"OV�
��q�^��3h��Z���q"O$� ���c��G�y��x3�"O��U�ĵb,^�U��(2�T�s�"O�cjɼ|8l���՗W�dhv"O�8��V,g��I5�Otq�s�"Oq'F�6Mh�1���C�r���"O�@ 5��:p`��ц&P��X�"O�,*�B�792��1��بF.��#'"O��{��Jzs(K�n��yplAq`"O�A�CJͯ �;�nZ3FF���"OZ�a�E��9n\���deZA
�"OX��gM�He�	 �=n��"O���w�Q,�Yғ)�\� �#Q"O�0
&�<=�X�UiH�X�t�p"Oju�C�n����HD;?#F��"O�)��H�+2���ȼk 
��"Ohj[�.|����3)���"O>���].5��2�.40튑"O� �ŉ���1yw�� #O(j�"O�@��@؜M"(��.H�'0i)U"O���6b�~,��r ��.v�kW"O.dR���R-;u/Ph�T"O2��7/B&U�1�t�\9r���jF"O쁣`�
�L9�E���
oz���"OP�W��0����4o��Td�ՠ�"O�t���͍0�A�dl&+QraZ""O⽉���mT �t̂�=B��D"O���EA}>��&��	{��܆�_w8��uj�=�q����<A���ȓM<�0à'�k}f��Ө@�>y�ȓ5��p��� g�*|�uI��N�ȓa�6u��n¶Ƕ�3���F�,�ȓU�8t�d�-,^�K��E��^���6qЭ�򄗷<�p��a�6�&�����L�#� #�mc����/�i�ʓH� G@�%`��� ���+dC�ɗk���FN�+J�����U^\C�I�@�& BJ��D��q���#r�XC�	�V(�ck�x��m����U��C�I�DeD	e�#YI�ips@ScY�C�Ih\�X��^�X�ဲLQ.�jB�9d��(�SFR% ��iT�.)��C�,vO�,�V�
�fS�)�7r&B��??l8uG�#q��U��AX��DC�	>�L��N� �U�!��u�TC�&;dB-������e����p�C�		Q��٪���V�<Es�k�� C�IAv��L��I�:Q�bc �B�	$<h��#T�
�Om`ѹ6eY�-�B�	�[c�U��׆]�$E��?�B� DD�c��D��-�
M�K�"O���C�w���S,�7��� "O���	ί3ΰU��ζd���"O8��D�B�#*�Es�KR$*���S"O`��$��T!�UpD
��<�&��"OR4cc��y�´sg'̤i�p���"O���wH��n�n5A%J�O���3$"O4%!��O�l9� ��A�3d��1i�"O�:�.�z��:��_/��h0 "O��KZ�x4�Өs7*��"O�|3�=�,��!���m;�"OP�"���:7>qpH]�����"O>�X�D3p��$*7	϶f�,���"O1ɡ熖y|R��P�b����"O(����̂9&��a�$���"O$���˙�FV���e��5>�M�2"Od��pĎ���$��K� ����"O�ͫ��+�hI��� e��"O$q+%g�$Ƽ�^-��mk5"Oz ��NYs�@�h��"J�;F"O$l��,/^��[*�S"O��S   ��     �  d  �  �+  �6  eB  ~M  �W  `  �k  Qv  �|  ��  N�  ��  ҕ  �  Y�  ��  ܮ  %�  s�  ��  �  J�  ��  ��  ��  m�  ��  ��  � � ! �/ �9 6@ xF �L N  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�	�� R��g� �t��B��1�s�Ee� "<E��'�����?l�i�|����y2�6�Şw}��̞�� `�d�ǁ���a����dE�D��p�i^�;>��S��%+�|�L3}2jN,m��+�lRu��iT�y���>�����Q�g�عQ� ��Mˌ��%��|ph�9IV��1�!�;qu��UA؞X$�>�XR��V�ԎPԜa�g��:]&���d(8a�МA��řcYx�h�G��%ڧ\�ƠB�!3]��`��G�44��^�Ȅ�-J�S�d�Ӱ%�'
<�'Bў��$��Fa�,ʕ0�i�9j.!�$�!i�;��@�f�I�Iſ+� �牰D�-�Dk�;�Q���c�C�	;<�4Qd �
����'�4��'��Bm_�K;�HاA�H5���|�����Hȸ-&�tbr�Žp#��v�/�yb(Ͱ6��9�L��o�(��^��~�!�S�Oaƙ�gh�[8|`c��e��e�'% �;?ʡ��� J���
�'��s0i�3y�Bd˖��Vy~9�	�'�F��A�^_8@�D_�M}F��'����7�[�Y��:C��JF���'�*ex��N�d�B��9;� b�''��SѪԮ4	�#"K��7cL�8�'����d �el�0J�g#����'�HS��Q��*�р�	����'a�|@0l�9�0�p�A|�`<��'/x2���93�]���:%���`�'W��P��҈4�����)뎨2�'R2K����y(J�0�D�Z"m��'�~���j�$)ԡIg�0����G��O����^�E�� �9rdx05$?��{rɚ��I�m#��Q��Lm��$*Ǹu��ʉyr�'q�x��H��t��ѯ���r�H0ND$��=�3U����"��M�霂���.�69���ȓAR�L��/�B��ǭ��-����=���?Q��Ӟ6 ʝ)��^�%x"T�&��~�<Y���7?=f` ���4~D|9qM{�<����J�Fa@o�`Ѡ�sS�Q�<�[y|�d[� r:���`n�EB�`�'F�|�ڮe��)҅��F��b�O���	^���O(���b�>�bI����O��p�	�'eF�Js��#y��L�Ǆ�U�
yK�}�x�鉷4��9{�ɐkL����N4Z�rB�IlZ6�+l�	<�ؽ���Pdֵ����'] �cV�`����jG�%��9�'jX-���_�"�ba던�Da	�'�bY��R&��l�� ���$��˓�(O��5,��N�R$�7/T�j�~�J#"O�BS�]9af�K��G�Y;b�s���=lO�A��ydVEk��ה:0��"Oȑd<$�X���$Υ|����"O���t.R9ǎM�1���S
nj`"O�:AJ���,������eh�ha�"O\�!��שn=Ҍ��$�	'�<Y
�"O��#@E�U��C��W�9���"O�؀�J��}:5��k
:�P��"O�D�G@فE5ZA�Cj`D����7O���df��	Y0i؀}�~��)I�5,�,���'���ɉi����AE\���z�&I����5�I�|9������?& �S &�T|�B�	���0p#� ��� �<}��B�I�Jz��5B�% dY��T�A�6�F������ ��A��ƛRTV�BpH�>���6"OL�ke�I�Z t�A��V)(��2dU�p���h��Q#w��
T�� s!�F�H�ZC�I,A:� Iv�CQ��2�iħX+`B�8P��(��_�!�l�s�H�3
R>B�I�T=dX�!��N�ZAz���._B�	,$��rVk[	l��-q-�)
B�I�e|Lru���Z%��� $��>r�C�	0����ThW]jP��-B�6Z��#��c%O�>�ȉ0�F.`�����4�O��$�QԅƪuJ�AK����>���0ƈ3D���� 	F��AƂ�5�a �M2扃5���?�|b���b�c��$��iIGhd�<�0�� T�4+	I����a�`�'O�yB	Q�$�� ��>;L@�cc/_1�y��%&�&aYF.đ-�E �Ј�y�C���v�Pg:��P�7J<�y�n 'Ǻӑ%�0�؍qbC��y�ώ?~�Pt,(t������	�?����v\8���,�H�Pu��!i|���ȓ@��-Ӥ@+n�P�Sd݃B�v,	��O�����!3��q9�(��D���fcҖ^����)"?��,�;�2%��۷�����(�f�<���H��z�eZ�j�
1I�<��l����v����¡К3^lm��	�!n��M{�O��e�k�!�"��"bN؜�"O$Iǣ�W�$�����w���S��D�O��s�{����P=j��1���{�|x{V�D˟̄U24�K4�ҔT�X��CDP�(��:g(I�&�ݱ*�������>�rԇ�,�*I�K�J��f�3��!�ȓ%�M�adT/J�������n4�ȓ�Jt�0o�zB]��j�b���^=�P������[Ôpc���ȓSܐ�bɇ,�����ODN�ȓ&��MJ�� m=j�%)F@�م� �]Y�Fѫp'T�C��J�[@�ȓ?�,�B&@�����1FTl��b3�Y��N��z�	d�.n�B�ȓ9����[��䪧(Ų!xPl�ȓI�@��Q�(]�r�I�Z<��O6�dұk������@�]�(��׈��H $��<1ѧԗk����n�hU�ݢh"69YŨ�<�\�ȓ[�p�Q��L�r��a��_p&ȇȓq_Mb�o˗%�@$�+�# �����<_p�+3
�h�F@�3$����@ua���7���9�'A.S�\�ȓ:����<%�.��P)��(����|��6�Ѯ#���ޠg��=�ȓ-�E�� '��ߓ4�� �ȓ"cr�@�0!{�	�fΈ�
@�T�ȓu+�,J�$��P	�)+vN6Utz��0܅�P/ٮr�\��v!�h��x�ȓ^��`�$5)x,�N8�f�ȓz� 8��O�]1l�RT"�39���ȓ{/������-��$~(�ȓi<ش!ĭ�_<"c/ק!а�ȓi�Y�&T�w�^��n�%4P��ȓ*�f�K�JB�$
��R�ĩ�ȓx?�W� ❩3 �.��\��`�Y Th.���)˯vD�ȓM��R��+�:v�Փ"6E�ȓz #U�$ut�A��7-�4q��S�? ���*E��t��Ś���(&"O�"&H�8��U��e)���u"OnQ�A��r<x�D+^�@:8�W"O�h��&Y���k��N+/���"Ob�p����U ro[�[Ά�[��'��'��'��'&R�'�R�'Ӡ���J<OT���ʗ/p�4���'���'t��'�"�'A"�'�"�'�4�Q*J�$BLc񧆈aR��!��'�"�'HR�'��'42�' b�'���D��'�� �1�u�3�'��'���'���'���'���'h�v��k��<"#��>2\�E�$�'���'���'vB�'R�'E��'�Dm٣��"D*����Y�r<�f�'���'���'>r�'���'��'&����
���`}�&�ȐF.Jp��'/��'���'e�'1��'��'"�����5`�P� �R�F�RC�'Z��'{B�'>��'ub�'�r�'@����k5c@�A�*�-5������'���'�r�'e��'or�'���'��)�ը���e��Ȓ?'�=�F�'�B�'�2�'#B�'7��'���'_dQWhV gg�0S�M��˂�'���'%��'��'Q��'"�'���AЂ��t��!�,�W�'{��'�B�'���'���'+��'u�� coK==�vlz���f�R�*s�'���'��'���'R�a�����O�Ձ��	{����rrgjm(*O��D�<�|�'dv7��%{�l�ƀ�M�hX6�	W�~������ܴ�����'�B�3:*Ps��0vN�y`�*T��'����i;���|�6�O�'
,�=
p��m��#�ن.
��<)��� ڧL�`��.MZ�^�6�H�APP�iΞ�`�y"�I���[{�T�&Z�g���Y��ʢ���O*��~��ק�O2؜�%�ik�DB������0〉*!�
�q�K����=ͧ�?�S�*2C��F�6[~PR0�<)+On�O�hm��CX�c�`y�h=/7*��c�ޠ70>L{�aLV�A��	ퟀ���<��OP� ����.�y�&e#�����D�O��	b`�Kz1����KzR�d�7o��0Jϓ�܉ɥ���xN�˓���O?��.ht����'RUd���r�	8>��٦2կ,?Y�i��O�I[�f�Q�&R,RPX��K0 @��O����O����xӄ���$,����
"&�7Ȍ���Um��QPA�4����4��$�O����O����X��Q��I��b�)��\#��w���K8N[�	ҟ$?M�ɮZ��r�͌�\�$a֬$V�L�{�O��nZ2�M���x�O���OfЍ8\�i{ �	!�)~�(i8�g��{��M#�S�D�$�\s�Ҍ�^�IVyb��er�� `�J�x�6x�(���0>�&�i6��B"�'��xl)1��}0F���Jk$٦�'��6�8�I�����̦���4t���GZ6�Z���	�c��T�C�
�b���i`��O>U�w습��wa�<���>�k�0t���ȇ��8<]�R��ΖB$�D�O���O��d�O��$%���OrIb� �&~ž��ů!���`�O����O�nڹ_d��ߟ��	ß��'�^ #3N�0�nM��-Y�25�����e����'��7�ѦE�S�n�(o��<��U/l����L�T���0
)���2p	ƿ~���������4���$�O��䍳Y���Y���0!��dN�>�P�d�O(˓) ���,W��'���O(��JǸ�T@a䎡F����/�8�y2�'W�Iϟ�l��M�b��T�O݊��B�65*���S;Q=���u�ئ,Ɯ3���
�����n���H�OȄ��cO�
���j�'��`����Op�$�O,�d�O1���"���n�vC���f�T8m$�u��L�Jd��h�'���oӘ㟠 �O�9m��O�.iA�[#e�t��b�1q��ܴ3+�V��"u��6?O����
L�\=��'$�r�A\�ˀ� )��:�)3"V������O����Ot���O���|jdhǱfUu:℃�0/t1��[�V��։�2NEB�'����T�'ȴ7=��8D�P+
r�hQ��{���g'���-j
z�$��S�?�S��HmZ�<�&	(]%5��o�*��ٴ��<�U��3���D	��䓍�D�O���1+c�AbS�μ��x��.��|�I��4��џԕ'�7��"���d�O&�UK����e�1Z�Z��LK4ZV�d(�d�R}2�}�^	oZ*�ē0��y��P�A��1/[6
~���?a$L�/���J� �����$Z��_��D�$M۞�`����X��Gp�!�d ����@��Դ��.�����
��a+���۟ ��.�M��w����&l�"4�`��� �6.T�p�'"�7M�u�ش>QꔮX��D�Ol��ƀ��r�͏2%�CfL�
����,J�O��?���?����?���E)�pC���.��1���E�X��aH.O��oڦm-��I�`�I�?͕O�C� ��!��]�pw�=��削�M���i��7��^��?9��EV���"RB��q �D��e���؂?L��I����OB��K>�/OR��c�ܐ!ҋ�4(�0���'��7��$�Z�dKD~�Q�����U�%���M���d����?�!V�4�޴:6��cӐyA��.X��[0J� L�r� &��6rb�6�e���	��@��b�OB�T�'����k�� D�QR"�;&P���՛w��M��8O���dĚ\&A eÝ�AH*V�{@�$�O$�T¦�cF/RҾi��'(����#�4��t�MtZ���>��ۦyݴ��U
N��M+�'t��J�\m*`BV4p�
�j�I5B#���3���x�|"_�<�	쟀�	��t�S@�'/1&�;2�A�Q���7&�ǟ���jy��|��qB���OZ�$�O��'j5�pc�F0a���!J�bG)$?��Q��X�4Z1��-�4�.��ܯ-ՠ\����=�$x���G�|���s�Y$��)n�<��'w`�dO��?�)O�,A"���Z�Bu�B:h���$j�O��d�O���O��|2)O�HmZ�{Qh1t*5S& ����� 2���֟X�I���%�T�	vyHf��5�GLH�?���HhEZ��LҦ`�4 ���ٴ�y2��>bD��aj��?����:���27[^��E�Ǐ�TE�5�঱{�V���	矔��ӟ���Ɵ��O�R��kI�|B�h�(Q/z�f��Cv�ک��O���O:���dRʦ�]�,[���P�RH��i`�d�ڴO��b&��I\�<�7-`�dMA  ba��N\#o(Z�S�l�$ ����i�b��j��ny��'���P;���BU�Z�10��@�˻,*��'�B�'�剢�M�r������O�u����d����eN7v�H\�d=�I����Ҧ}
۴;މ'5�1�!�3+�����R�� ��'_���&�J�b�#t��?���'���	?�,�@d�J
2pa�/���Iğ���ٟ���J�O��5u�2t�5i��Yh�����:k\�`��[��'86m�O֒O��L;7�b��c�Q+E��!�'$�*��$����J�4LK��i��b꛶:O����l@���'�5�)��|�R��OԺH�f@�������>�3�5�7F��c�x$��+�n����'��7~����O���8�9*���!�\�d��,�vꂠ�JՂ�O�-o�*�Md�x�O2���O�j`��''�F��3焨9��1*���R�D�q^�B���L����q.�*� �2m�:S���a�I����e�6Ԉ������E��p�&�HpΉ�
� ����<_^Td!C`��X �C���y�P�S��G<�a(�5o!�|�0�ti
Y(V̞��B%�����]mڤǌ�;�T*`�n�I�^7#��D0M��}x��w��+%��� �؞J������i+���޲�	� 1k-��:�ŗ1�(P�Հve
@����]CDI�h��^F�acU'�p�<AH1�P$9���I%E1Xi*�'K"Ͱ�@��n$h�J6�D�*���L����P'P�P�E�1�W9pj=� ����?�H>����?�RHt}b��.�b 0f^>d�*��S�?��d�O��$�O��<`Xȋ���􋁉x�諶�B5yb���r�L.�7�OR�d�<����?�`C�ţq�Yy5��-ly��X�C�>LRr�{Ǹi���'��I-5���O|�����1H<z�F��wg��"b��moy�'��4��O���M�#��zJ����M8��@f"�¦=�'@����ddӎ)�OZ�O�@�e�,�f&L� (���N�*���oП����R.�����$�'��L<a&e��6<`<#���(�����C�㦥��;�M����?����2�x�O��gLD2]�.���n]�E�
��%o�f�Q�ϳ<���?!�g��?�'��?�ni�F�ְ/��h��
>r�6�'���'g��@).�4�L���O�`E��<��\��E4;���Lp}B�'."DIߘ'��'^�@�T<p#�M����a�0��(I��7�Oرs�Ax�i>���ßȗ'=h��OUZ@��"�"�`8xCBz���$&qB1O����O����<aĤ��{I����^1�L���3��=���x��'y��'��I���	�玙2F��kD��ʔLR��R�B�;�ߟ��	��ܕ'$�IBdu>5����KY�,$�4"%(�P��>����?9���d�O ��
/}+��$>��`�d�\'�&|�T�:� ��?���?i,O��V�D�S;6ȼ��"�"URН0ㆇ7�Ecݴ�?AL>�.O}�C�iB+�̓�_3��-I��̈G����'�rV�P��5�ħ�?!���P�գXs��c�6Z�KB�~v7��<����?!�Ŗ�?��U@�M�ֽ���s \3dzӞ˓S��s5�i���?Y�'#��	e�vH��k�g��(QU�.-"�7����'D	�E^���&���5�\#��؀R���:(��)u"w��v��צ��Iʟ��I�?1�J<�'��e��U�f��,�>2;@t���i���Z���I��3�	埔D�ڡIhW�;2�6��6$C.�M����?Y�k2`�ҝx�O�2�'�&)ʒL��:d]���>R�,,HTM�>���?��Gn̓�?����~2K���.�kHU0�>�sC�%�M��e��(O>���OV�"�;U��@��s�xG�4�0���g~"�'O�Z��I���@c*ߚ|��CE�A�w�t�	�Mpy��'�2�'��O�D;w�4�js��-B�b� X~l�a�I��I�����_yR�'�lt��ӟ��#���T�I��ȯ!�浂Z\(�	�����T���?V-�W��Doz%�+���8�mh���F2�eʮO ���O�˓�?��dD5��	�Oʕ�p�Q�3�HAJ2�P�>-Fԁ0�Ȧ��	m���?�bdN�="I'��;AI�H�� ��'{��R�EdӘ�İ<Q��r��,�����O*����U(>}`e��/xp�����<��y�>��P��nJz�S���Ɔm0D9�� /Ew�j���9���O��Z!h�O��D�O��d����Ӻ� bx��,�uN�pQW��8j��mPfZ���I�&(� A�<�)�S�~��;P.�;>�����(G6�7�\D���O���O��i�<�'�?	�,T�`�`��r���Q@�6⛦@J$3D���y����Oy��H�57��)�*�8��9�lJ�������h�I�I(�	�����'�"�Olq(�"^*A)�p���1?�J�$�x̓�����T�'U��OBH�b×<��H�a�[�r�~�{1�i��^�)/�ɟ �	ܟ��=aC-]�p�S�eV;(��W�>���9<SB0���(?9��?A+O�$����"l @P�KǊ��_�,�s��<	��?����'8R-�*��[�E���`lC�G�J��.@���Ol�ĸ<��g%j9��O�<@h4ϓ�+�X��B�����ٴ�?����?!�b�'�j����[��M���ռMP����@�On�]��
�E}��'��\���ɢG̖O��jމ�b<��o�
����C�6h��6M�O�����W(�ܫ�M-��I:`D�AꕽvV����ޙVZ�&�'�Iԟ,"#]I�D^�����t:��M�3�&�{w�F�t}:)C�}�^���t2�Ӻ�T�@Q�6��h´D�<�k`�V}����P������ßL�I�?	��u�S�	��m�P.J�
*�mrcZ���D�<!)�K��ħYD�����˅l��}ѕ���A>B`o�;{���	����'�tQ��ȟ�9!o�9*���xW�F�*� �)G�չ��$��b>!�	>*��0���͡S�H����$�,�+�4�?q,O���w)�<ͧ�?1���~R��*W�H hu�.DD�5	�D�./�`c�dR_��ħ�?����~Bg�<Op,��B�>7R�i��ǔ��M���O��LZ/O��D�O��d?�	'N��<a�o
U�H}HC��,\t�}��d��e~r�'��R�t�	(4e��)�mN <z1rAᎺ	�9���'�2�'�����O��Q�kR�R���,K���ksd�k��(:֖���I��`�'X��[#���
*a��TJ��ּg��I�=��'.��'��O^��5 
1@u�i? 
J�R�����d�/o�&S�O����O��?�T�����OR�C�h��1`�e�Fi��� J¦��Ir���?q
Wr;�X&���F���pAC���66CHQ�~Ӵ�ĳ<��-�l�+���d�O��	��$#��0@��N��4��BX%Nl�>�k�	�u-�~�S�Ĉ@9Q�e{�˝�)=F!{��ȸ���O�	�#��O����O����.�Ӻ��E�E+r���Z�T�{E�Gn}��'�z\�W������O_�))!�H,MV8��1+�*+���ݴ�a��?��?9����4�b��L�d�(<;�a�#8Oʠ��"�V�pn,CiZ���6�)�'�?���e����3���%b��z���m����՟����Vzy�O^"�'����	M�ƽr��5D80"��2D�e�<	��׳m��O��'���Q�"P�3-Dv#�R�@��&�'��!�_���	џ��I{�.[� ���}X��vk�U����'�Ե�����$�O��ī<!�k�d�@�J��� &-K�6t:@1b6���O��$�O$� �I4z؁02��04t00��s з\\��?������O�Qrl�?�![�x����]|s��Ђ'~Ӷ���O��d,�Iޟ��ī�!�7�C����)�joB��Dcχ�����vyb�'�x��G]>�����]0��)o\	������!m�� �?	�X*ĉ��@�-j�"�m@x�Y �d�n6-�O�ʓ�?ٗ@I��)�O�d�z�r�.�)e��+d'ϭrT��2��L쓸?�!�U'wXj�<�O iz����M,`L��V�R�:�Of��T�K���d�O&���+O�N��0Fܵ�w�ȠB�~4��Q�)��I���9�M[�8stc�b?�c0b8m�򎔞Z����t��`�P�OB�D�O&��럂��|�����/Y�EJ�
߰8�(���Mva�-7���<E���'��`�f��@R�hr�'D�¤k
h�L���O��DޗZ�b��|����?	�'x}:�����$i9���� qa�o(�I�"(l��I|����?��'�6���!��/�^	VgM�m����4�?Q�������Ox�d�O�➨)�<0}~�sNV�W["̒!�>فM�M|@�'R��'J���������� ������*��́
���Q�<��?)����'d�@� ' h@��<5*��a�_Hi�u
��>���O����<��'�*DB�OFn��4a�'@1R��R�iK���ݴ�?����?!�B�'�D	�ÍI.�M�^�ez��w��|���ʆ��j}��'�Y���	�,<�O����&v٢�$�[�s:�#��o�H7�O����	^q��a;��}AM��� ���f��4Sn�6�'����(��%�~���'���O��З#��br(+�Ҵ��dZŇ*������v��1/Ѹc��R�ti�:������U�'�".�M�R�'e��'���X��]
l��₨,HP^��nI+-��?1���
�ܥ�<�~�o�+��IC�L%4�j=�������s ���M����?!���&]�Ԗ'��`�ˁ(�� �p��<�`��WMi�rس��o�'�?���\�>@l�G��I<��� b$x��f�'�2�'E�􈄀�>�/OH�d��� �
�d��c��Uqv(���W�ib\�(
�r���?	��?��90�h��MS�`Ԓ h�-��V�'o1O�>�)O�d�<���{�hL!$�ܭ�ĂI=Fp��*c}����yB�'@��'���'%��noR�yT@F�a���� ª �d�S��%��$�<a����OT���Oh�C�搀eV��Q!$S�6�y��bKj1O����OB��<vQ�Y�)�.En<!b反�' �P�1`U�l�&X���IHy2�'���',���'����$I�@x�er#DB� ����jgӒ�$�O����O\�$���QQ?��	�$�V� $h]��F��r��)Q"��4�?�+OL�d�O��$��aG�IJ?	ǌ�VF����;`�Q����Ħ�I��P�'O��j�$�~����?��'ZR���'��n=� Kg%Y�	�r��_�t�	��H�Ɉ_ ���$�?��q/E -�H\���N���#A�{���S4t*�i���'�b�O���Ӻk��?A).2F%�.^�Ф��������P!g�ԗ'�"�I�I��C1�Wu*����ԛ�I�|�6��O����O����T}W���v�s�\��0�(e{D]��L�$�M���<!M>�����'�Q�v�F%&��"�N�?Ch!#�!eӄ���O��dB;Oeʩ�'&�ܟ��n�Zh�@+S�a�Ek��4HU�5l�K�I&v���)���?����10f�*�}�Aʐ�@<;��iB��*.$6�Ob���O��ćD���O��1��D	ij�8�FO��8�<��sY��"�g����ߟ���ßX��\yb��#�:)�)��8�(8i�MN��d;���>	.O���<���?��'���1��7B��)��fV�(��F��<y��?�����X�Y���ͧ$�Ɉ�mN8$�Ђ"Ɉ/!�0�m�`y�'U�����I̟`2��y��!�
Q� �s��T5a�@U�«߳�MK��?1���?q.O�]�w�Gp�T��5V��l��4�R����Z�O3�M�����O���O�XY7OV�'����N?2HV<kG���U����4�?����d�)y����O���'�����wn����c��aU�Sr�˼5�&득?���?��n��<�I>��O�<M���H�\U}�sa��$n���4���
� B�(m��h�	��������2�x���,T"�tF�p9�� C�i���'���<1K>��4�Pn�PT�d%O�s?&�{�'_��McR�Q
m����'�B�'�$"�>�/O�pKж(�ģ& T8~�Z��Q��ՠ�g����Ky2���OJmòE�3�Z����3*0<(�j����Iɟ��	+�X�ɭOZʓ�?��'.�3HYz�X���Q���y�4�?A+O�TI�<O�S���֟�3�BƮGb�9F�8$�"풢h�<�M����°T��'K�P���i�:�VZX���k� �����>q���<	���?1���?����D2|��,��̛u�&p��k�b}�Q���Igy��'ab�'2z	��L#[ux�Hu��hH�Z���6����O����O����<���Y����S��Uذ���)���0w�"Zܴ��D�O���?����?aӇ��<��8{�Y�HJ�a�`��C�}��`m������۟��I]y�F�v��맾?�1>R��U,]&|2t��$H�^/
Tmҟ�'@B�'I��Y9�yB�>�"+I�F�.���V� L<���Ҧ����Ж'y" �J�~����?I��,ix��e����I �Ӟ8[RT�QT��	��	�Ez�I@�	OJ��r��P)@Ϟ�LBhU�fNZϦ�'�n<��j���$�O�����*Uէu�4r{$���I̾(zM�0�
��M����?�4���<YtR?�	~�'f����AĘ6b�I� E�9v�elZ�ca*۴�?��?���=c�IJy��W�h�4<��)�Rtc�.{�6��?�:��͟h� �ؙl6��SF�����fW��Ms���?Y����*CV���'Sb�OZ09�3�E��_[̩z׻i�rV��k�y��'�?����?1Cӿ`�μyԇM�c����.ݗc���'�H� �c�>y.O|���<q��D��J'l[�L�0�S��V릁�I		�$�	ğ�������D�'�r���lŊ�D��NL�z�֠0�#.\5P�����OLʓ�?���?�eA�e�"D�e�I�p��Ä��S��͓�?���?����?�-O�`Q4�I�|⠂�;o����A%26��a��Dz�	�T'�D�I�0wm~��r�H=;�  k�26vQF�	����O���O��4����v��T�N���Dfة���"� p�~7m�O�O�D�O�m��D�Q�^�H�&�/�=4��-����'q�U��@D�֒�ħ�?���Y���d�D)b� l��*���q��x"�'T��\�b�|�ԟ��	E
ۖ����w�o2�hr�@�I�R�{��i�&�'�?���[��I��		�.V�seh��#*6m�O��D&&��#�D#�&|B��q��{#9\&ڨ�@�a����C�殮��ɟ��I�?u�M<�� !�ᢆBǟ?�*�4�ڂEP��q7�i��ۙ'��'���dy��'�Pdq���XU2�sD�-t6B�j�'q�H���O���G}l)�>���~r\+��Г��'6��a��-��' ����y��'kb�'�`�*� ¸|��`*1��	�Ӌ�ݦ)�ɀR�H�M<y��?QO>�1_]� 25�H��B㮚�>��|�'E���Ƙ|��'Z"�'���#;���*Q��D ��
�ێBm`TJ���'�b�|��'���8� 
yBq��XVp!�V�_�x � ���<�-Oh�d�O���BԻ�Q�|񂄵��й�
�.uM(L��.�I}��'�B�|��'���?�yR��IU0-�r��P�,
e���?����?!+On���p�Lq�ы���c5��3`�9�ڴ�?YH>y��?�����?aN��B�m�qiژJ`�K2�x�j����O�˓�J����D�'���l�>~z�)� c}JB�a,��m�tO����Or�:o/��r�@D	x�Ƭ���	�A���.�ߦ��')XI�5�h�l��Og��OK��/B��Ҁ�=h��T��o��|-l�����ɝ���n�S�'U{��8�5-�<�Jr�>l��lZ	@A�9��4�?����?i�'3ԉ��Ĭ�<t������R�4�	�\�g�6�������Ob�S�O�2%������'b�%��nL�i��m��i�B�'V�����'N�����Ugv����Ѳ3]6<��$C"c[���>Y�/�@��?���?�q��J�I�r�#f�hM�v� ,G�v�'�>�z�]�t9��Z��9���+EKХ ��!n�e��"�8y���'+*����������O����OP�D�ZX۠�/}����!S?�q��ʵiY��ʟ�������~�KPh�:��(;��ѹԮK@!9挊&�䓒?����?���?�6�^��?I�A5	�b�2��ʿm�T`[���&A��f�'d��'{�'e��'����<�M+6m��HH�6�4���v}B�'���'���'��Q��'@��'�@�fE�@����%5�����z���=��O��,vMHy8T�x���)e�I�.A������M��?A+O �!ET�$�'��O��;��[.�F�s(ױM�
�cE}�:⟴Ф��D�����R12s��)Vq� �υ�aឌo柰��)p��!��ݟt�������FyZc�@��c�V8�8�3�H�@I" ��4�?�@�Q�ǖ{�S�'x��CD��'9��e�W*{f	oZ�0���	���	ퟴ����$'?1�G������vc�1��_��MS��>'�q�<E�T�'��a0���Q;�4��m�+)���p�D�O��$%w2��>����~�$.N6^ݛ3�I�'x,Xp�����'�Ҝ��y�'�R�'�8��tNю��u�J�ye���on���dB0�U%����ܟp&��X>U�fԒ*��R��Pp�GR���3���<����?���$��T��}U��@8��X%I�Z�H���w�	ӟ��K�Iӟ�I��q���p
�%P,��QR� �2�I�H�Iӟ�	�;�UL�C���n�<�k ٤U�j}h��O��$�OR��4��OP�ąmV��7{C6��ą[���$�j����q���b�95�U�!�ݻQ� )�f���ZDD���5煵Pi>C�I+�F��1�]�i�t�E�mi���a��]�G�-(&�]#N�{1\�����2f�""C�>$���V��1ad�䌌)�~��F� �&��|�SǄ�F$9���R�Ã$%34dP�'�Zv����;6d*��q�E3�l���M32�T��¹s⤡�Ӡ���		�B)`��x��i�4*qP��5"@�XoЕZ���?	��1� }}ڽ���� !�{f,X�>g>���ᓣ�µ�)O�k��p��H)��}E�܏"E,�����ZtHDC�nѿq�A�)O?�DN9v�HY5��t{ ɟ�]X�s�k�O�l����O�>�:�r��V�(t��[P�R�BH�d�O�����{���5�J�9��!�D Ґ
����4����37���+�`V*l-��cu�\�����O��b�gɸ(�����OR�$�O�ԭ��?���{k$�듇�2�,�I���~����')6yh@�C� ���~F{2� ������J:�x3��={}��dE%)ѠUŇ�E�Y���hO(��p��+H�6L�)�Z��F�O�P!0�'����Gy�燛tل	�t
"Y�l2�d��ybIY*)oX��6MP\(sMX�gij"=�O"�	?5��MRڴv,L%#!��5L�����c�ʴ����?���?1#LR�?��������5��P��HLH3k�*z�(`��Mϑ:�DD�C����y������ 
�p�N���A�G�-�dƌB�*dnI�/�yeƌ�?�� ��I0aH��c�8���iWS�e���D.��9+N��B�v2��F��iڼ�ȓmf�c��Y�_{�}��a��ҊYϓI��IRy� ��t�.꓊?A(�����9���CE�n
���W��:2�L�d�O4�DYKюR��qLY�Ѓ�ȟ�'�D3�
eL�I%��h0�Fy&\�&K��/�8V�K0X^�#�.�(<h(����3v�9�J�7���Gy�k�=�?!���O^�H(D��Xm�` ����>���''�2�_�!>,!�f]�J�yB#�� �0>�E�xr,1Wt�ے�#�dK���y��@�-<���?�/�2qYW`�O����O�([7╌(2`�2��)pyRf�&BW�u�!�K7�:��Ɗȟʧ���?� -+����s(S)���ѐ���ANE�!P��d�${����0��7�Z1/��xG��?u|W� Næ���'�r�����O���nYWpI���#ܨM[�"O� ©Br	ԿH�Fl�̤f�AX��ɝ�HO�b�����̔l1��K����ڟ�B7��^�y�	����	�x]w�'�����v^$�� �|���'P e�䔮0�Ԃ�$O䴘d��[p0��(�x���O�a#o��UN,E�x8�<�v��_:�,*#ѦnG	�Q������OR��6���Z��zkC�D?g~��:�g���!�DDZDik�ʗ�&>��5��� ���FzʟN˓M�
�Z�i��U���ͺ�X8��Ƹ.av���'��'���^�r�'��)�#�r6M�OT��w�ԃW¢��0o�>:4����'�0T)pQ�����M4E��c?:�t�¦'-�O���a�'�27����XѪ0#�1t���[�F�R��m��4�'"���?�iGc�lw爺K�X�:�`2D��ꃁ�L��� R�!�4A�0�t�l;�O��l�hf�i9"�'���\�T�r���2�����,Ұ0>F=1�E韴����L!E��u7� �<�O�(T@���V?�H"�;�8tr���K�w�����퓅��aK��j��Z�NZ�Z�<�5��՟h@�4R�6�'P�S�D{��%&�R̆),�5Zz��IE�S��y⅀�{�`�yT�̬�}�'�:�0>��x²،@��ޛ�z��׳2���SH�h�i���'��VE�y�Iǟ0��(egȨV�F$D~�h�g��J�`��M��y*��<Ȑ%�Y��Ţv�<W��B¦�-5�t�����'+�u�i�<���@3G�Д���ڇ!��'T��:#|�	�n<���4�
�P�`%�J:vE0�	�����ɣ uvL��@�-~b��`H�F1X"<1'�)z6��#Y@UkJ"Wr�xwC��?Y��p�����΀��?����?���Ss��O���F�V.�#q��d22��g�V�]��$גt�>(���'T��� $���@/�Nj�3�'H�))��̹��=����C'\pC6�H�Zn�Xa�0�?	T�7�?y���?�gy��'��I1���:c �	k�Uy�n/L�VC䉵��xRG�%D���a�-v*�����ـ	�z�d�<�V�5o�[�w�����gcX(��Lԣ:z����O����O�����O���`>!a#j��Q;L�oڟ�q�� ��q�R��p��R4��$K�`-���v�jӬ�#	E<W�y�Dd��`�����'�X�_&� z,L���2����5:V6M�O���?A�ʟ��� ��: K���c �%B��Ec�"O��CaL
�fK�|�@!P�{�F83�6O>��'�	4J����ٴ�?	���T�US�����Ko����oP"dq��2E�OB�D�O&);ŁP�:.a�#�ɜK�	3 ��y�t�U*XTbE�,P30�F���J2�(O(�:w.��l �Ÿ��^� ��}ZD!�~"�c]��ȴ��'���{�mN_�'���	��*����o��$�|�P���)���cA�/��GG��?���9O\�r���?}4vY�r&�K��!�A�'66O��Q*�t\\��VO�z�4�AC?O\c!cV:y�����O��쟎\ZP/�O&���O���&͖9�n9Q� E�b����V+\��E��.[�0�pHoDl�8��O�1��)�ZU�����{s䱸a�>`�HD����F4�ga/Hp�Տ� j6H����I ���eɖ���w~ܴ�cB��7�To�IGx���'�.��D�,7��!�à]7.���B	�'
�!Q��B$oj������ e�	*��D�I�����'6�����z����(%"���'Q��ή ��Qa��'	�'�2�cݙ�	���x� $z0�2�))A��m�E��ؠ�۠]踝��I4I���Y�mء0��	cmH#�R��\����J�A؞ء2ЄQћ���0R*| �&�ܟ5�ޟ�0�43ޛ����O�ʓA�4�Z�ɺ8�he�I �M ���ȓU�j��wo֪*�H8�w-C�A�X`/�HOj�'��$K�%�F!n��=��o]�FO���덋S~���I����ߟ8�����P�	�|����2b�4nI�	 �K��h&͐e�&܄�	$zaVq�a�˦����7d� �pb�ۊ&�ޅ�#�O��{��'�6L�B�&u(pDur��dDE��ym��Д'2���?�P�+�`
�a!ra� �,D���(R�<-(!
!Ԙ���i��٪OP���娢U���	j�TK�23���Dm��ĔC�Qt�P*��'�"�'a��9d��@�j�	!�,�T>�8�"Ǚ[���(R�7]�la��L;ʓy�j=9V�ˑ�%)s�,g����*W�?����J�b�KR#B�(7�;FL/�`����	��M۠�	�=g=t�:f��}fV�@�/_B��D�O^��dR�4���f�ƋK��Q�ň��Z�a|�a%�� &�y��f��U�I?MON)�0ON�K����}�I���O>��t�'�2�'J<�"��g5��M��0-��I�r<������x�T實�l̈�ܟhb>��P�`Uv8��W�w��Lڳ�3R9IbE㊛��Rdo�$+�"���Y4��9i[�@�(��Ͽ�R�V�$��[�)��	�D�@� �,dj�a���?I�O���OD��9KV�ĭ݈�l��1O��$2�O,��)œlrz��r�)z��՚�I�HO��'��y�ϖ#u�Z��f&ڞB�����?�7FA��L�a���?y���?�v�� ��O��J�T�n^�4b��!Z=r��O��bу��]�`��'p�pJdL.*T�ы�k�ktE��'����J�-O��ϓM��D��h��/t|b���(\���M��(� �v e��Y�l��Ky2�C�5�z�@1�Ĕ &g��y��A+r=�4��q�X1dC�'D�#=	-���O�n�F�Z�;��U� �N�C1f�)8!��R�j)!�H&U��� %f�w@!�䃒p�X�I�$-w:�`:��άM&!��B��`��c��`1d��pd�->!�D�:(B���H�k�h����* ,!�T}7^p��
�T��	p��N�(�!��O�-��9��%
����C�=@!��
�1��L��d)f��� �Y�!�݈58�U��NB���\B	^�3�!�R�%�N��aH�	x~�Y�� �!��\RI�$�$�M�sg@���
,�!�䛁3r*]�f]f�j%h �9V!�=^0Ԡw�ڡҔX�%�D;�!��S>5�d<�􌏚;���+�m�!��D� X nذ?�!t�/O�!���;�&���-z>z�넊жb}!�$]D%��k@��&#6h �L3ou!�DjD|�$��1d��Ș���Z!���B��`���H�~��` �,׹on!��"}�&��w�$�d��"-�Py򡃘9RZC�ˈ]2� ����"�y2 ��J�H=����V�d���g˹�yBĎ�
l�Y4o2CD��Ag��y"@�. R`ɂ��
�){�0;��W�yBoنC��<�e��g����
Ǩ�y�ܳ�D`���1\�1ХM�y�e��sT
�(�M6"���@7EP4�y��F��=���Eņ:$��y��T�g~&�0��UTЂ9r��K��yR웦H��ts�愗J],��d(�$�y2
ԙn��x����&7�$�G���yb�U���Hr�/�@ 6E�6�͵�yR���:42�IС�N�t �ML��y����RT3 ��K�P��v�I��y�I� w7��w��
>�� ��5�y��Ksh��r��04р8�ֆ�8 ز0�I��@�'-����h��'`���b�#v�M`D��|k�P���
 Z�X�k7�LbX��g�)�hA���@���qa,B�P&�`l(��a�y��D
�;LҘ⟼�R`S�w�5"�G]2>���*!O*�i��	9_*z�����6�^y*�e�yͼ|�ƥ�>^�mf��"X� ����(�
�q�*|O*���0Ժ���oS� �����<<!n�*"�X���A�D^����'�K�*G�!���H�bd�2@_� ���?i�)�ȓP�B�	V�ʔ:$�q:�#L��N�J�%M�$�<M���	�w5�$mڹs!6��T>��.x�y�w��	�iL�F"б��ޥT�a�
�'?� '�P�[̫�,7"7pp� ����?�2aɮ>�"Q ��J��y顥A�j�����d �X�h�(t���hu���u/ax��T�'QP�0r ^�_L�x�mS2�Ψ��e��x�
��OY� �,HR��|�Ɖ�#�P>=p�{�*��j"I�/
�@�*�2��$b��L.2��sV�Xd!�a`tMP1L�P�S�'�&����.Җ|�W%�e�����"O,b��3��8�u.[~V�Q�� A��9����o�Š�e��;�,f��|ʒ���u��̻y� 5C�C�A� T,Z�I�E�\rh8��"Q��J��d��=�%�G>} �x k�2�P8��ӡj���uȽgrFD��w�*<�#�_ǀ�d�0 �px#�ң{b� �%r�$���`\xCc'_�ب��J��O��޵W�VQs�ɔ�Z->2%LS�e����
N�`̦D��×�$�r%P�\"�u
�d�O|DR�a���!��~ʟ�]!�d�	�$C��T�l@@���$@�.i�Mچ��Kd�C�*D
tɓbҴM���~�\��Ƨ��4����76۸��S��-���[d�Q3z	��s��zC�����x� \-6�d���S�W$�(�'��'���7�J�#SB�|���+}�K�(dti���ԍ0�BHr+���yBN��
�Z�J7%�71��G}�[�hF �``_$��(an�J�{�4 Q��*��w͔33��"$��O�	Xr�.�l��m���v��"ZU�y*�E�+"	۲�ɭ �^,�Q͊��d�!Ԍ���7NB2So$��K��б9F�ӈ�O�d��`��h��]\�è&c$%1��) }��w�_PMҔP��1���֟Z ��+��_���t2�_B�'GhE���-ʆ���E	q�,@�#iV��6�	�,T��P�'3j���6%C�E㦅����H�D"��8�VAS�U.s������Q2�nك�f�q%Xb��=K:X�/҄I�Tt��`Ն&���@y"L�@FT�}�Vlj��1�K�X�H���j�B�#����A���'��#=�O)0��q�:��*Ď����f�Q��)(F�C٨OB�jt��)�ְ��O��^�x����5(�V�0���5�qOrY��'�Z�0@��HY�~R��S���^O���E �;GZ��Nԩ{� �'���:%`��w8B��':��{���M�m��(��-�hCCHD�T4O�x˲��`?�D�'���ق�J�lk�)�A���}W��`�� p�P�b�#�`��s=O��	'��1O�����H�#����Ŗ�P�+� g� 9V�z�HME՛��xi8�x�al�IF�A�����Q���<QF�p�(O#|B`�K�N5H�0L�B'�:XW�E��iI� iDP���߭���	}ցSd�6^�E�.F^��s�ɉ�'��!x!o�?�	.0��Q���0%Y.�r[��Z�N�Rk
��$٪0YH��ƅ�}�b�XW�ڢ@"�
f�#1�h�9�&7��A:45O�R���^�I$A�q N�y��#�>�e�O�."v��
I�3�tZp�T�$�.�U��h?���M�.[��O���@@E�ajR�ٰ�7ul!3OTE�.E�M�hqQ��֡�p<ɶ$,n�U !�� $Y� ���Ł����J������ x��e�<�3扊�$��Y�hi�OP"z����
O`�"��=0������T��0��b�jܕ'�Rt�?��'�Lz�wT�6^�q�b�Bg�S-]3��i�:fyKׂZ C[�h��LM1�p1�ग���,��$���$�����n� �`��Y��m�д; m��a���/[�S�F{@�tmI�%b�'}F������%�~��O�XT`
s��*B E�%����AM�p'x�`]#�D���YFV@ a�)ck�@ʵ*X'����'F�a��cE��2 �%��*H`"�0I�ʧi)�ej�cA=dZ��A��\&/�.5�ȓ;�ā �F�S��aկ�?@T�7A(B�h�8�Ƙ?���O��5�r�ͱ� ��DM�H�찻1',D��S��e9�$���.$a�x!+�;:1�';��S����Ϙ'Eh� o\CD�'˚:g���3Q�֨@r�$3@�π12��q�[ӈ����D�wn�E�u	ۨIহ�GA�.HEz�J4����� �4����-Kڑ�GG#�b$B?9n��ڶ���]�x�s0�?�!1e�|�'d���ߊ]C@��tJU*Tt���*R��'�rt��F_�t���"�Y
��l�	V���L��'���J��h�$C�&`����t��z�\B V�����7��Ex�{i��[� L�x �J����$��j�Q7O	��lxʷO�r
��	�0s��;�Ŗ�<{�b#(��*�=�a�>'.U:�oܖYo��a�I�ZV�1fj@�Wu�L�q.Y9F4q�g�T8�g̶�'��%�' jO�S�b�6'R���p�I :�`q���'���*&R)j&�q��-q�\[ �I��y"fS�\����ٗ��Dͤb��	�o��d��a�I�}����&�a|B��O 0�0^V,���֦(�W�NyV���mр��O��Bd�4t
�%ǚ�X�,�Ϝ!�.�ZDIÅ�K#�ʬ6��\��΍G �}�1�����N`��1��̞�� ������a�� CKT���i��(�Oh�h�f_(I�N�W�+��5<}h[a.%-:����0Rs�\��O����q�T�Y~!1O|�hYe&~�֪	�n������D�O�}jX;r��,b���*�㞝��eڻ�9v�5|O�a�V᝭{��R���L=c��,����@���1R�����������]�Cϰmk��x�Z�%�|��qc��)���;f�S�5�<;���Gl���AnҸa�T3ˡ�8`F>��?��Ef[��U7�Qyu6��.�?,�n�KqD_|�#<�g�ߙz��Lj�EL,;���h���<�'�ަ�2�ca�T0vَ\���F��=Ț�\��!+C$���r��L��'JB���R ^H@�����Qlb�!�,D �8%�� 
=[�.9�y��B �@�
��ё�~�����R@NH!&�#�/�-�D��`NEd�ebj�"y"!��E���Oe ���8nԢIi�&I;*��d{�A&b*�$��r႔�RJ\�w�D�O�9j�NL*G��T����-g<��d.��h�����'���Y�.��`� VUJ���:'�fL��a����foD� w�d�.��Ɋ
	��gd�?��4�M�,vFu
t��=�R1c�(
�lA��B9Iu�T*#�^=.&C$b�
U:)چNYe����	7�.D��]�h9�� �/v���r��S�8X�4�T�����`����<׈�<��AFQ�l�TaҦ��1������=�d�G-���9��h�SL�V��=�t�#j�I�s+��~E�kA$ͱߊ��H��y7£?���We>��`�(|�K0	S1��xU �怈&ȇ�D0��˟� � 5�`�
5�D���m�s3:P��IF�X��P�@�;��<��AV����λmo~�j7�D�#`]P��y/�\����6J�
�@��<��ۥign�*��E��`\ L~$�
8ߦ�9B�$~}t	����K�'�r=y5@X50��L�w�	|��6]>��5���0�dt��� �`4A'��IK�BW%[5�	0evq��SCyR���Z nP�.t���C�+O��T`a�����=q�`����Û�h����/G𰁒�V%`�qP�����r0	;h�lt@��:C�<�t�O�'6d �$O�tPYD�"3 ��RiS��A�G�� -0H�/�u��O�7�t���z2�l��_�-�@�REEّB.���#��V8�� aC5%�
�:�w'�5p�@,U��3�-E]:�p�O#W� ���y�h(�։��
�(� ��jr���O~r��G%}���ޞ*��=�G�Hf�>��"��/^\�{pk�/:����K?E����W�ra!
�4C���@�N����81'4F)�M1�`��N��#|/O�$1�Dt�l8@W��8SX!z�`X2�N�BƖ#4�
�!4����>=��"�jG�<��=�4�K(3����(��6�x�Ç��3	c���6K����O|uQ�ׅU��]�Ta	��j�f�G�%|\Z1g͕���x�� ��n���?���郍I����ի_�,��8�$�K3+>ٚǓ>���ag�"jE�A���%P�l ��C�ru��l#�nx���y��K&��"r[�t�s�QN���VJШ�viF�>I��#�薅@z�>�a)�ZJH'*ʇ]���C�ă����;�*)�R�Z$_�(��$L��ɹע�B~"�H,�'kU�D�R�?A�'g�i"��
"P��R)�]��͑u.�b
��
?jR��a"���O�����'�01p2}���f�&���H�J��/�o ��k�cB�N�%�Óg��`y��Q��d����%m̓:o�=ad���͢L8�J�~Z�?Q��I�I�^h@Q�4Hs���v"�����)"�1ѠZc����`��\�R �7���/��o�	Q��r1h�ȥ����y��\�Rtؕ�ECT����@��T9saF8:���N�U9޹K�}iE�7fB�8��ݧ]i�i*�gU��'h@��U.�av��BE�]bdŁ2x�$��I:�Ɉ�O>ʤ�3�^H�'�lhB,�%V�L����<��1CDǖeL2x �	�6H
��G�3��O��4���T�5����Z��a�@[I�Z�Cq�Q#X^P	���6J�ay�ɉNY�U�'��9D��X�E�0�9��-N<ʺ����5P��:�S�� �?�&X���&韫4ZE�UE�(���:�/U�+�yRM�=h��8�'����17k�'.J�XvB\�[���@!�<)�j�)1�n��'��ҧ�s�f�ѧ�4���m�R��_�ƀ���oV�N�|	�p�W3/��HI?Q3�#� L���� C���Ɗ՟�H�8���?7͊V�`���-}�L\�~Q{��$%�l���%MĴ���w�IPf܆-q�Y��,O�)��s,�{sf�
��(�#%�ZV]9�X��
�MA<i��Մ㉞k���4��:Ջ�
�L=�軒�N+c8�A��@�8-��S�,O�e�'�>���ŊN �W�D�w'tX@���ԩQ*қS�,��ݿR��Lc��^DuB�S�ℴrvNP+�'v�!� m���)��iS�c�BX)^�� Z1͕�a��Y3q"O��m��#SIS�ѣP��+�"O~4��m�=-��,���y7"O±xE	/6�p �cH��>x|�r"O�M��'_��L�6A��K[�Dc�"Ot���kR�H��O� �,��""O1��.��.��Q�Ɣ*��Ɇ"Oty�O"DΝ��]��´{�"O~h�r�W z
�� �dL�|��"O�T(���E�������P;ıy"OU�'i��~��%*퍍;��9&"O��"W4)���w"��V��"O�@�&��)��!A$!	hܸ�"O��S��e%@��ّ���""O
ݪ4J�:0�fm�eo� >�~� "OzXA�́� w$$+��C�D�����"O� ��_�"��|(�Ɨ22˞T
�"O,ĳ��.D���єc١P�=h�"O�l1�Ȫ����P��F|e"O���		
�i���E�F�>-��"OAI���=P�I��(�?'{�E��"O� �dަI��-�)�au˳"O()����0m�@���AK �Ha"O�Y�����`n�
��F?�x��"O�i(%F��K���c��N+hU"O�Aa�!=~ �jҏU�#|���"O�9��Î3�q'P
��qb�"O���E�҃3H�s��>NՊ�"OB�jp������9��^�8"O�����̏��ZؙW���!򄟏�6L3s&U�q�\�)0�~!�D\d�"�A@S"$2�xA4^�|!�$��u�u�+,;J@���9q!�dV8r���x&��317�=��@ f!�@�dYNq
蛿2�.(�ՃT^!�D3UB@��g�u��z�'��Py @�9#��p���.x����b� �y��Z,!�
Cd�mZxp���.�y�+8%�- �M�0i�^8C���y�Bx�r�h�fסj�������y��F*��fǆzͬ	ڷ��5�y��E4c����>odȤ����yB�֔-�>��4��j�0 �&����y�)�~~n%�S'�e��8����3�y��78WP̳� �J�>�`����yR$ßSj��F�ҙIE�5�s@إ�y�JƷ/3^����P�pT����y�
��LO��� $�5��U�/Ҭ�yR��)VOt��F�Ж&`���V��=�y-���Z��M�-��	���y�ke:,�c R�(�xYR�"��yRǞ�T[�	�V-��(��Aѡ�,�y↖�8��S�/Ȍ����
&�y�FF)"����CiIv4�7MG��y.��Dm"��%��@�6E_ �yb��m%��A#H���t4��0B�B䉕+���c���Q�7/�5W`���A$j��#jC�#�=��K5t���ȓ�(��nP�W����@�/�@	��1 ��D�y��5#,f��&:
�q�gŰH�ׂ��<�|$�ȓ@~|��u`:@S&�%1�Fi�ȓ�v)�����_)����
��Wu�`��<`1J��.�ڰ�Շ!�n��ȓ!$�bs��HK4=��烠@ٰy��caX(����U>	Z�N�F��e��^���"�؍s��,��G&�$%�ȓ="�i��=~W*)����f���ȓ%#$�4#�1BRG2xp�ȓ_�e�t�Yp���gdɨHP@�ȓ6r�1����4r�2 x7-B>b<��g�%Q3���N�;P��%�ȓRK~�C�Jԙ.*`x��8 ���i����u��xbU�$i�����ȓ;2��Y}�2c0׬P�� �ȓ_D]Zs,�� �7#؎Csz�ȓ1��+%rt�d*��F$�j�ȓ}T�����"��0�ށ��N*U���^.�	��L@ ]�(���V���G"ԑ*�"�d�VT�ȓ;��Hz5O� N\�9ceG�2�6�ȓJ3p���JǾo�������4�ȓP�RMS2c߼9eȽaj��K����ȓD�t�K�l�~��@1�O�B�� �ȓ� ��-�1|��ǥC��Ʉ�S�? �4З��?8p�z*V�a@v��"Olˡ��!)�}�ی]+l(��"O4�r��Ag:�)��"l]9"O�=�0��PA�]ZTG�K�q!�"Ov�����7�h�%��!�j&"Oi�-�gmf�Sg\8(���r"O��B�֊5PV�@�f��4uH�"O8q�.1�2�A�^*Ȧ0� "O��@�,!-�`d�geO r�L���"OZ�C�*	/!���(W�F�2��p"On��VO�S��(#s�D'�y�s�	P��"���]⎝�Gi�r�9#$���@"��KXx���H�)*~��0��3�y�%A7(�I�Q͞
	�~Q"����y2抔R}����M��ܩ�+��y��W�a^�IP5I=3'�;掊��'_ўb>���L���VśO�;M�R��s":D�����q[�]��cԭ\y��0�l,D��0p�_�P�M��ő�
��lA@�)D���̙�uD5𖥐?&2�Aj��'D�|)��e�C���,�Ex�'D��6��/���)e/*>ql��1�0��E���'g������=w/�ivKԐ�����Z�����#C'���B��Y�RO~u�ȓrB���3'�c�J��$I(**%�ȓ�v��TH�8�`��n��'�"���q*��0/W�L5 �#��/R��xG4Q���3�VMr��ΓbP��ȓl�HhƇՇ΁P���b��}��Zi���E�՟+/��� �4���IP}�Aؕ&��b���m�@�f�Z�ybNȾe�|$�d,M9�L�k��D7��'��D�����D�q%c�6z��  C�0�`�"O� �J!(��:Yr�\ �ў"~�;#(<ےN	��uI3��p{Ь��PS���d��Ss���`T.4JR�ȓr��:.�1׃�,�T�"U��e؟ ��a��Uc����`��v`%)tXH�ȓ-��i������q��դt�(��y��e�%��j�f��d%&7��OD���n}���Sj��'�<I�ȓWNȘ������o�q(�ч�-�atȇ+Vt)dk!��A�<	�
����d�=D,ހ�&ɉt�<iEfA(��Ppcw�>�k�nm�<YD�V��PztN�5����
i�<�0�W$1��ύhL5���^�<��)B������Ev�x����Z�<�p&��i��a C��.��<�#��X��@̓	��,2e��D��!	�#���<!�u0��⯈�|�X��E�r�vT�ȓ��Ȓd��{�Ԙ�B�q�踄ȓn���Z��CZ1\49K�Uf�ȓ|�������*x`P�� L��%�ȓ���U���,p��ϳ����ȓp"�թ���!��;R�F�%���g�d�{Ư���Aʶ�ϱT�fu�ȓX�8�����p|�P��iʨt��m�ȓ=6����&�8��
�Y�h��ȓCBB��'�q�z���� ��)�ȓ��$`c ^")��I%�*/���������/����$�&��C�.�#�%W4<p����&���݆ȓa٘����pp g�	���h��S�? ��s�v�*M;�?
`��"O�× E�QSvXx��B�%ؐ�V"O�D!I���F�C�/�u �|�"Oj��A��n@9�S�M�{��xH�"Or�#��Rb��rU$aێ(�&"O||�`,ݙ]8N%�L!p����"O�Aqp�)/����1b�|��"O"]c�BZ�f�h�C�;���V"O�5 �.V��@a
�xx���"O8x' �1R���5�G0ktv@S���ą��7w0��zG� Q��m���X�e:�d1�,�@��,/���*�N�u1X�6M$D�|��ʉ �֬*qN�Sz�h� D��)��ȩ>�XBt�$o�.m�k>D� Y���4l���ۃĚ�lL
���N>D�0����;�P�*���7kd�h?D��!qg�=m�z'Rw���fl7D��: �,j��&�M7F��8ʷ�5D�d[u��=v\Y��^�[¦I���2D����,R�,���7�2E�0D�T:�E2q4��YC�!HC� FJ,D�\�6"EhP#K��؄�(D�0[�ٛN�\Ib�ݑyEl�se'D�����nY��9�e=,9��.$D��� �q�6�	�jY:�p`	&D��#��ېB�qR��k%� zqN?��蟤#@ �95�R��@��/Z,,��"O
\��ϋ(�3�,D 'CHс�"O�=�QY�6嚴�I�a"�"OF%J�����ܳÁ�>`aK1"O�Yp��2
��+/Y ��!r5"O*
���*,ԥs��'/�fu�6"O� uj��,���S�%�6��"OPH��ʛD�Z�[��&\�T��"O��P���P@]��݁�R�"OlL�3�		��AC�Ƚ8��8Q�"O<��v��X~R���!+��iB �34��
�o%j,C��N�,�hw�%��`����↳{��#�e�,���"D� ��,�f !�6����5�E3D�H��X�]~���Dk���xŚ2D�Lg�Rc��t�m %t=�'3��.�S�' �(h `��+J�,��𠙴	.��ȓ^VD�@��gf������]��1p�1��ۉ"@�v�
|B���V��sAT�}j�<���a�F���x�r����%O��`E/�
L�l��\bq�d�rض���X{���ȓm�6��6�ʞ�H�YB�.��Ň�V����a��}XF����@<~$L��ȓ����"R�Nm�x)����K���"��P��ȀM��U��D�8��܆�H8�����?�H�@��Y������)� ��n�u�3n��c�h�ȓ
^Pp� ���1ؒ��$B�F��ȓ7����AD:��%F\�a�ʓ�$i����h��x�� '>�
C䉱M, �r�S@��
�o�9�BB�	�b_�$���v`TH��#s� B�ɀa�
�A�C��c�Z$�a�C�~��C�I\�E�UgE�R�3%���X��C��8eQ�YҥJ��*!4�[���(v��C�ɓkV�x[rF �|QD�A�I˯��B�I�O N|����,~�l���7|�C�)� �I�DX�\3���Lm��%"O�٦��# ��21*�=O2b4�'"OV�ڑ�/hs$�{�U�'>��Q"O�9`�Ǎ�!B��GDG�&0�R�"O^��e�
����I���"OnIآf�I�.ʑ9�� S�"O��S@G�lFD�Ч툪(Ӥx��"O�Y�Ő�)��h1�`���&"OJ��P���l<��+V�T����"O�:�	MN:��S��5�xi�"ON���t�$����W��`Lk"O���(U�E�Dh��V����"O����.�VY�(�,�T-��"O�A9"
��G~њ�G�m��"O��j���6����F��4�H �"O\`ae���$=XǓW� �H�"O���؟SI"x�R:�L�	""O��#Ta�0��B$�P\�k"O �ze��(3`%��eN
�)K%"OhD��59V�@�0I�(�"OrȢf 5]>�JW,ݬp��1x�"O� &*0[\��C��p��"O�)T���R��tk�A�`M���e"O6�Y�� �����b��'1\��"O��c�.�P;P��A�d%�U"O&��'��Je��!���:�N�+"O���o����"[k �X��"O�9A��HET��e�_N� �"O$�*�'L�"��	�e��N.�
�"O
�R�E )lܠY��l!"O|! d��f���a�i�)0�P���"O8��M
.E,Dp�tƁ��pY"O<��g�M��"�d�/C�Hg"O��A�V2���#��o�`�"O,��"/_� ���2� �M���rt"Ot��w����(G���8n�)��"O"!��G!	���0e��4X=� �"O���"W�xΠ��IÄAV<u"O��逍��©b%����
:U��ͅȓ!%� ��ឮ.�<!�0�8F��ew�iHu���= ]�bÚ�ep�9��}���I#���6�l�*f��9j��x�����DD��;֐ S�cΜ!x���@�á������ࣛ./$�}�ȓUjF�h�E/A��`����F�T��Bo�(��اd���%��!K1�Մ��D�!���?�&�	v/2v���KG΀�p�@&E�d�9sGO0�6�����y�gĵLm���T��A��'>�m(EHٚp	ty	'm�7W񂄪�'�V�8&�́T<�i��疹LT�L��'/����-L�v�˵&D�?�z���'����@O�R�x㟁?����'ά�Rկ�����Qp�hAxyy�'��d+���rJ9B �M� 4�I�'��r��4�HaǮD�wb1��'V�����s���sgG��v���'�p��A�/(4��c�?�����'���#/ў �t�ranU� 6���'��@2A�?���k��M4(�	�	�'utY�,��f�x����]�M�'Y�ukW�%bn�=��A֙\vd]��'d����+�� T)S#O�̙��'�a���X���1zc�=|9*\���� ��J�䁹�R4�F�������"O:�@� �T~~I���J��a#�"OX؃��:��k�O>��]ze"O`��&�'��,(T�'�D]��"O��ː(�U��1���Y>�RE`�"O��#JN��#�G�8�p��$"Ov u,X������
"��w"O�`���"S�ic%�K";!�$3�"OT�noX;��m�P,��$����`"OX��S�B.n̎�A���
-�5Z�"O��2�ǀ�Lc��3�MB�'+�ȠF"O0�",�o'�D`Ѣ�3OL�"O�`�P��$Y�p\�Fa]�g$��"Oq0`'�pD�9�t������9�"O@�`f�̾U]���9e��B�"O�qs%���{�T��6�����"O\,��@�vC�X0e�>R��DA"O�<�ՆH�^2�dOA9�>��G"OکZ�m�+
�
� B��T��"O�A�S�L�'�(���]���r�"O>�	�J/�z��3Oݠ��\H�"O���ꋭ�L��t�
�@�a�"O�I;FϳԔ�A��ެ�9�"O� �ש[�ի6������"OB������+�F��D��d��mH�"O�����.@� ͪR�)sF�15"O����!D'>�Vɗ]4N\�"OBňe��I���<d)��`4"O@i��k�&q����vg��F=S""O8�(�.� ��С{��I�""ON5���J�,F	96�0=���+�"O�L�m%n)��ŉ�=��Њ�"O���R�ǜ{�6�іnV5?� ��u"OR����=dI�(��h�!�@���"O�|� fʡH���a��ff��X3"OH�'�9�F��n@��L�2"O��Z1��':v�u�U�,���	�"OJ1p�&*�l�[��%�l�p"O�<!�F��	�gII44��Y�2"O\� .])Z�  �ZsY�ɺ�"O�M�b�F�<;ꍀ��̠"<�-�"O z"��9L6����
VA��"OȘqb��y#դ*���q"O�$P�ZlY��W�Qk�R�BG"O���R!�@�Ҹ�� E���Y%"O��bd��7$�ȅ�Bo ���"OLp��	�iFL9�k_H} ���yB����ʡ�¨Q�����(�y�$ٽ?,���v�V	���!MY2�y2	ZGP]�v���D[d��y2�
�M�|d珐���#�+�y�h�1�
}"1mI7y�����
�y����tf�{��v��x�lI�y�O�Mx$)As��#�Z�"��X�y2ʆ���"B�P���i2�y�l 0cm(�*��X��XP�a���y2.�a衙2Ɍ�0d�"�ϊ�y�@҈L��`뉫s���cg��y�����ԝ�+hV�y�GR��yr-�K�<3�a��e�ہ��,�y��/{��8Ү�`�V��q�]��y��T+^zbh�akީ4��!	ݍ�y2�_2a������T�Æ�r+zM����#܃K6���F~��S�? �$˰A�%(Hm�Soޏ8��9�"OTt���߻=`�h`���2=L�3"O��{p	� pJ���l�j�z�Kt"O�@��8�^��%��c� ��4"O�`:�KU�t��e�e2F��J�"O��Y�E�3	b�)���13�k�"O�9h�/�D5Ƞ�N�!0���"O4�$*T�Fj4��F�u����"O��(�Đ"�� �h���ޜ��"O�|Sg��8��%*T�?fL��#�"ON���٫e�@	Q�!%/d���"O:���a�Na����G��6-����"O��s��$titFN��9� "O�i�q U���PC�Ԝ[i(髥"O�=��͐�$�0�Z���oLꐺc"O|�c6L�(5�R휮i�m�E"O�`.�}h � m�8H .�"Oj�+�Z�$��L��U1N8EY�"O�q���5oHqb��:0Z`�"On�8�ےf*�"���S��7"O����(�9p���F�z-��"Oe!d㗬i��pǤЖy����""Ot�����7E����dA�Hw�xA"O���.pն;E$��k��"d"Ov|��/gc��h�����$�""O��0&!�03%�Ȉg��!�Ұ#q"O��,ղyք� F�)]V�I"O ��匇@�ℝ�FM��"O8)(��߉g��	3T#�.q0"u��"O�9��m� s�=� �&�� ��"O*h�tK��Yk��څ�0qΑa�"O�����7h�YC�$��G���"O���6�̽j�욯G)�Đ1"O���w�PX�ì8=p"O�9V��#����ϖ)����"O��dAǅ)�H�㖡�)?'`�s"O|AsֽT�}���Ԛ\-���"O�������e}Zi�g�"�3�"O��p��O��ؠ��v�|��"O�@ժ�r��b&��4�c6"O0E�aZؤ�g. "#�X�"OBm���(?Zhq�W#Y*�^ĐR"OԴc3�<Ru���#D+	���D"O4`���c��h`B�X<y�v���"Oꑁ�kҎ�v%Yb/� 8�2�)�"O.�@埁���e�"&<�1R�B�<y�%��nO��jGmP$x+@EAbD�A�<����^d���ă*I�~�t�}�<�%��� �0q�&zYa��w�<�fcŜ0h&4��i�"j�uÕH�N�<	���8VkR�	sLˣ]�ze�TB�<q�NH���Ѳ�:̼k��|�<�D�hj�캲��9��u{��r�<�s�˺Eh��Z�)Y�@��٨a'�l�<	��wY~��Gَs�UX�&_j�<9T���� �Jցn�z�����\�<�7���D�1�D>`o��eA~�<I7L� 2@��5 
![6�=�ȓ8�Y���^S��	��m��O!��a���bC�.F�&�1�py� ��U���s��R�rf ����*�a��~>�0`aS�`6���X9%|v)�ȓ5Ƙ�"ĭRv.q�g�C`R��ȓl�<��J(���P ����S�? ���F�Z���8�iK�A���A�"OVy�vd	{�B(����d�<���"O�q�'�L(�c��"��s�"O�����i1B�F	SQ�d�P"Ob,3���p�$�`5)�+4 �Y�"O��1E)̳F���wǍ�E ��"OBE1㫞%%��*qf����c"Ofq�a'� Dx����`;�͠u"Oݱ ,Q�J鈉ٴ�&�a��"O~y2wDIw�6�T��&�N��7"O&Q�@���@�h �gJ�d��U��"OhX1 n!��2`��|��T*b"O��� k�����㟴v�>-qF"Ob�ZW��3�A�����3�F��P"Oƌ�2jڣR�b�q��_u�PzF"O.�f��/>c�%Ʌ�à*ɮIt"O�1�Q��1Y"�Ԍ�:�R�"Ox{��ѐ0۠C���T���"O��4iТ"��Q�5��8\�� �"O�m�(��I�zu
sJ�\W�]a"Oн��,O�]�x�J� ���`Q"O����L�R���I�1�إ:w"O�L`C�yb�	c�JX���"O��#�dJ� J(	�P���5�0�  "OܨqB@�G.��DE8��l�"O��!���Ph�p#���P�ƥb"OJ���O(�t�R���  t���"OzR�A�w�����h߻,�ͣ#"O�dj�MJ=C�ҬPdI�(T�<3$"O�Y�6�(_�y��'�3kL(5�"O8�҇�7�܈P�-��E�ܬ��"O±+!`τC;b4d�P�/�� "O<�PCe\,}�B!���B����:w"O�P��F��FE��-ى,���Yc"O`�D5`�s��΋*m�Q�D"O΍YשV����ǡ��w�u�"O�Y�l'a��峰���`�����"O��#���-Ҹ��S�	t�Q�"Oj������&T)�#�@�JVҬ��"O�Ԁ ��҄�0qy^0��"O��6ñ^�f�qbǆs��h��"O&M:���i�t"%GJE���"O��D��MP��AeG�6���"O��Pc*ۖ94�x�#�9Ik�ep"O���w�l��;3#F� k���"O� ��O�t1�1��!T��0"O��`�X��H�hR�Ίj�؃"O���&+åS�x���OB��A�"OfEД"��c�-P.�,�~���"O����D�7+A�Ap�#K��Q(�"O ���g��zc��P".] t� �q"O4A�B�F|٢�U48�ƙ�"O��c�B�&J�A�7��� ����"O���G�<0���� 	Ӣ1��"Oj�¢ �'t�fK��-b����"O` h�C��&���aC�mkF�"O���$�Q�$(H� ���g,���"O�������8XaW@P�j[nMC"O (�E�K�>_�5��΂v��Y{"O�"�'O)��}�����d�V)�v"Ovp���:Ǌ8k.û6$�""O$��ec�b��;O���zH��"O\��Q�$�d.ڄ#|v�y1"O�48�ɟ�4l��"�F.^Ԑ�""O� �՚W�H�0��5聏����t��"O����I:X)�1���`�<0��"O�Hx'���%���bR*�����"O@�4�0"��dkPO�b�=h3"O>la�C7M�8��s΀#(A�s"O�]��Ըua�!ya` 3W@x "O��� Kx8q����+	��
�"O�	ӕ%����ЈPh�� "��"O�X����=��� -"J�S�"O�����7(���U�N/a-�`��"O8�K�,�P���
���L�Xb"O�0��ȾG��XZ��V�*j���"OP ���t
D �����OΡ�w"O"))��Ј�n�bv������D"O��g�ԋ{׸��ek[�l놀�&"O���aC������5ѐ\
2"O��Ke	�+w�`t����4�7"O�z�&
Cs�(��lJ
S��zU"O\$����>�$hV��% �R6"O:s��R"G@�eEJ�atk�"O
hA��$g"x��ݷd"�Q�"O��ɷ��0^�xi4�?y��%x"OD��q��~:�0 ����I`"OR� �CA|�P9�`iG�y���X"O!Yd!_�����"ޒY�dڳ"O���G��'%-�R���*j[b�z�"O�T���9�H4C��pHpH��"O<����&t׾\H@���'-|a�"O@�� ��0r��@��
�ũ"O:���bt0��!�1!�2"O����Һ>B�u�׆��B��I�"O�,c��8!�i�cC�T��@b"O�e+E��)]��ȅ�W�!�|��"O�[�iދ ޡz�M�p�^���"O�p�	7nT�"�D4�4���"O�D�`)D%ٕT�E�g\!z��\g�<���P8d܆��7��5��YF�b�<!�b  
B�w�m�v�_f�<Q�+ʲ@001v��}.�����O`�<)t"�e��9+t/X xr�,I�'_�<a���/e \�(ULH��=�$d�c�<�b�^S��;�F@T�� ��c�<�bJƭ(\��D`(]���6OBD�<y��ɳi�,�b	l����%�G�<9�ŀ�Y�쁴�A�O��L!A j�<���O��rrb�D��8WgO�<�J9OmNU�«I�5|��`�l^T�<� ��#4α�V @�f3���A�O�<QcA&#S��aS��C>��0��D�<ٓ�7���g��"�X�㡄V�<�`HY��%%��E)z=A�nB�u�jB�� G�F)।[;��]j�-�C�	�4BF�t��5;5��b$9�B�ɜ0�p0tD�Y-}�R�R>�C��I�����s3 T�cQm��B�-"�v0���K/�R��Ҁ�0e��C�I�c���;���)d��D��RH�C�I(���:��f���c��A��C�	�*�h�sG�ŨqĹ`eFԽrnC�Ɉd?���I	9��"��Q�C�ɏv׸�z��":k��T��D�C�ɤC~\�۠M�=L�ʦ�E�"،C�I=|��se��H�؛`o�mCrC�IC���"��C� B6���e�>C�)�  ��e��B�j�C�,4�Y"O�łHM)UBS�̋F�lܪ"O2d9�H��5t�0r��/i�H�u"O�<ZQԷ+3hI��ԯg*d�V"O4����@!V�
Ha�N.z(�tB�"O���"��"4�@а��E�x��s"O�\��G�S��I���B�L�bT�C"O$�x��WSZ�Œ��K$E3΄Zd"OB$Dˎ�����g)҆��@[4"O�����F�n19s�T�xs�t;�"O�œ�G_ lb�!&�$N,Q"Oh%[%IB�qmH�B�D�4�J���"O<p(0��X$j|�c�3,u��q"OP�	�C 5:�thA��]W�`B�"O�d9,Cr�9�+]7SN2T!"O���p��V�JmzÊ�!֑�E"O4��R�ܶUV��a� h���G	W�<�$���  �,�dk�-P-���~�<Y��O�j2�ec���2� �'�U�<	S�M�C���U+֑�Eh�#
h�<����>m�4��o	v밍�3��`�<	�'�
b�� ���
h�`�$�S�<q��M�{����玺���C-D�<��)�70��!���H����aA�<9E�RN���P&t�ӣ�R�<�$��;r9b����(1]Xu� gN�<����FFڄBal	� ʨ�8�H�<1���ώB`F�&�8G�G�<y�a���P���cNd�6%H�<��H3
�(��~Bh3��A�<y3+��*��qX�*�7�"(�S��|�<Q�άA�p�(Ө���<ʴ��x�<�oK*�^9�D�1UyHtY�V|�<i�*�l`أ!�5L�T񱤈x�<qE�0?2Hl�q��V�T��E�p�<9Rm�Y�j�"��KL���kǍs�<Y'�P�K�n:0��\��"�K�t�<yF�n�`�3N�+ ݪ���o�G�<Ʉ@�nH&Ļ)H�֥"���j�<���
w�z)!G�4���C��i�<�pm�J����V�5�-�B��z�<�DMǖ���O�#�n�@/D�\R�!���|I{��ԋ>�Z�Q�!D�Ts����{��5�֬R/.P��� D�pi��_�\�f��x�A!# D�p9�KׂW���� ��{�"Ͳ�b8D��c'���T�@A�ݬ���E�:D�|�'�ǹM��H{�(��}��R��*D�t���P>%-��"��)
�咴-D��q�n�'.�H����߼3}$�;��%D��htH�&�
B�	3��1.D�ȃj[�)<�Y-��a�����. D�43�Em�ui������̓��(D�4�Sm��pԭA�o�
�t��l;D��6�E��� F�]!R(���h&T��H�
}N�� �Y,�$0"Ox�s� =���{F�=��r"O2��M�x�4� F�	�$�x3�"O�X��K�%V�椠��8x�`v"O���v�������$	+N8�z"Od�R�eF�8D�Q�>N��ԢA"O���V.��v���#\)�D��"Oh��@�Q	�
����/��Z�"O�p�"�فK�J��%
?݆"O� r��l����eOͅxePs'"O�[�#�`��s�$*p��*q"O�|qf��0pJ�j�� y.d�`"OY@Q�������K�%Ib!R"O:�a��Y6F�eFV�]4�	aE"O�]!�,�r�ڥ$�9��(�p"O��(`�G"]ax��5��6�@\Z�"OpE�kٽK�26�'b�+��yr�?|���W] i�~c'W=�y"h/8r��9��-v|�SF��y��N� �Z$"&�ԙ.���Bn���y�43z��e?.i�" ��y�/>���'�v^�HH���yRO�:�<�F���k-f�H�#T��y�/�/��Q��@�i�@P�a���y�%�-8��dB�\�v������y2Ɛoj����QL|%����yϋ�=c���� U�Huc�����y'A-��ѻꁸ8i���#��>�y�@	�|��ĺ�A� bf-�B���y� ԎD�B@��dʫc�20�q���y���%O�z$��îb�R��FI��y�o�v��yB,�>Pۤ��$J�yRgJ�F]���#i�F��)ub˃�yr M:J�@�%�؈!.5[DM �yR,*�ܠBQ�
��<����y�Ƥ2�bH׏��Y��5�yR�0����B�o���Ɗ��y�հ�@s6�G�o����狃�y�"Y+[ۦ�J�nF&hUH��f����y"��?�~��5!ĩ,r�F���yB�/��P�%EE=#;���X��y��-A��	G,�H�0�'Z��yi	+ ' .	��8b�Y��y�b��B�zy���>�bԸ�>�yM��$X�Q�ɔ4z"I��"��y"�Z*F��2	�s��p�5�H�yr-�(z	�K(���c���yr�Χ ɮ� ���j����!W��yRIڟ>��,X7���~��˥�y"b�BR��P��O�u��%���3�y����u�T0��Զ%�����y�i٪&���3�ς����f/	9�y"τ*9� 	����#U]�6�֝��xB�_:l�3��d`0Q��B��ds��)�'#��B�x��\��� Ԯ���'ߨ(�dM�xF"+ѠOy: ���'̈́!�a	R=��|Y0Ζ7mV4��'����7��Qg�]�͇|��)�'	��A@f�I��=b+��d)+�<�0CJ�Th"�`To��|��őz�<�BK�5x�Q3ul��Ir�	quK�x�<�CF�	X1���ڻz2`XPǗs�<�.I�E͎Q�&��M��ĉ�Bp�<I�YA��p�3%X*J��i�<��A�E�Hba ��S��(W�1D� �r/I#-����" �+j��!1D����M�^���1��QN���0D����ݏ0��Pa��Y�Ytn��1D���3;g��s`%41v,���-D�L��M#"N�T��F��dJ>����,D��;�ϛ-���K�'L�V���%�?D�l�r��q&A�ui	7<8&j��<D�L�"I�k�i��*I���A:D�� zL�ԆV|�@�ц<=��B�"O�"Da��3�%ѳ�O*9��p�U"OT��܇|�<�jd�X9*k^$�"O�*�.
"�� �um\�}L � T"O����g	�^NY�f��*���)�"O�����	4�p�y`�3op�8b"Ov�4�[%j�2�4�C�?6�""O��ыК]*��聎��[H��vO�e��ݷd ��C�P� �ؽ���O C�	�'��cQ�'*�5��c�B�	#&)Q���*t��׏C�7��C�I�'L8�BcJR>��5Z�m�=x�C�Ɋ	t]ᇧW�)��1(�,�	��C�ɏmnR��5$�k5��4��L�B�	?4�&M!��[58����O C��B�@�SnI&�RPc� �XC�	6f(M2��JͮT	��Er�B�I�B�Z!) 4�������@T�B�I ]X��s���	}�h�*
�kB C�I���P*�-@�`G-Fu��B�Ʌ:*ݠ`��0�"�
�䞷T��B䉄W�}�5닶)ζ���l"�B�ɤ^��h5��_e�q��,Q��lB�	�::�0�4�� a�ii��5PA�C�	�.w�X@�	@�x��so�BS�B�ik��C�!.�PTJs #R��B��(&|r(��Z<
�X{���?"�C䉹W�LB�`�$m�$�6b�
b%�C�I�B} ��F��Wꑸ�O�K��C�	�p�n�:3�P����	��C�ɝ+���)���$d�yR���3!$�B�I}N���D��,2��"b�˼x:B�Ir��Ӱ	T�3C.h�.�(ԺC�	�|�HeJJ�~}|3�C��u��C�	�6٭:D)|�#��L9^�̄ �'��twkB�am<�2&��]�4<#�'`�Y�GF�&�hMY1�G�pΈ!�@"O rF`��V����jǪ�ç"O��"�Qhf(8�)��y�]��"O��k%�K�� �h�.���2"OPH��IR�gߜEH��V�;(F��"Op݋2��7F uY���EDX�7"O2�aԙ�t�a�\���qg"O|�)E�bu0����BE���'�I��HD{J?�`6FH,B�h�����09���,D��r2�88�a"�F`���vF D�8�w%��o�v�b���˸�Y`�9D�$���Î�%!���Hx�,���8D������2��%�DH�df��Xt�6D��PPbV���tRD��"c��P��*'D��p	�Z5��K�x��q��#D�0�hT�����͝�qQ���,D�81#�C�J4HL��&(JLy��*D�4�#��o�$,[�nޣx$��Jh;D���!�1v�DKg��z���w�+D�<b���h�L�B,��l+��ia(D�(z���l�(�i!fm� �@C䉬G�ny8�eJ�n�d����T�PC��!n��ۦ�M-���EҧeblB�I�h��rjC�E� �+��R UBB�Ɇ$��HӋ�p��H�I5V��C�	�Kc�D���H�+�>�s4Ø.SM�C�	 &���PW��0��JD��"O.�;@���Zy)�b(0s�F�d�<� �e;3�]�n���Y�V90��![S"O������\5<b�B	�(d"O�Pb��)@Al<��- �G&�-Д"O,�0�H^ M�Ђ$��F|�p"O0\#�I�rS��gE��w$UH5"O�a����i��A�C�L�G i#v"O~� �'��k�h�aA�߅�����"OT�ҷ�[9�%IR`ѸC��"OX���â/�X��s �!A�J��F�' �	Ɵ��IM�3�I�C.5�éD���РdT�*pDB�I�E�v\�`fJ�/���!�P<#\B�I�{���2��ϜF�j��լP��TB䉲.�,�(�A��X�|"Ċ�7тB��+�ș�F�A4�X�.�7I4�C�ɠcf5b�y�P](�La��C�I�yhu�4�ßtU�k$�A�B�I�6!<h�%��;��"�N�rB�ɱ�@ZR���I��dP�HU��C��~$�@�(A8~��R'L�|�C��9
�����(�1��a`�� Im�C�I6S�>�p�BܕTn�a��Ȇ�=
pC�I78��x&�RI��� �Fq=RC�	 ��	�oJ3KΪ!��oU�C��r�L D!�x%8��e�"8v�C�:&����aa��Q�d�BL2�;D��	��31��8�	��U��2�n9D����T<p�5��IK><6θ��a6D�0j�뙭]�` ��S\^��7�8D�4�c�ǾyF���TH6rD	�&7D�T��`?*�蔢�ᐭ>�[�2D� �`K6��
�iκk�@�Z%D����D�:=/YX0g&���3��5D�`��	md��� f�q7�>D�T� Y7*h�;蝛\�f�C1O=D�L�w%��RN�$@gjְaQh��TG:D���de�""���X*�@03sm6D�
�� k1�$�a��(�4ӥ�6D�0!�	A(U��ٷ%Y�l�x�5D���g!
0�Y�"�V�*&�|Yn.D�@C.��JX��M/cg�tu/8D��%�Į}�h��u�'A��4���(D�0 A��Dպ�qP��7Z�;�d$D��
�B� ,y{#`R�<<��Ǆ!D�`q5]!jH�;�a��Q4�	Ƃ!D�vf^��.��Z�&��d���2D�|��a 
l�,�H�W�w|�P��2D���v*�J��T��I�Jר�)�`$D��c%۬V.�K�*�T���o'D�����P�<@$�7i�8/x�D��7D�|ѫ]!B�J��f�2"j��s"9D��	!/N���:��R�J��<ȧo:D��ђ$W<7�B����(1�D�7�$D��[���t�P�8��
#8����("D��-),j�p�FE�~��
!D����I֨~f���'�	38Ieg9D�p�2a �v7��3�D98�M[� 7D�t	 "ro��J �@��	�6D����O��/��"���7*��p��>D�8�gF߷K�$���-�\�b=D���)΃Mf�K1�
'���%F<D�t#8U7Z����N�0ȃ'D�أO�p,1󂉔B��[�J!D��(�I&f�~1��FE�.�٤�=D��h�"�.7ha�эD�$��2�- D�� `�9%��9���Q�*c���8�"O<���Xp�N�R��6tO 	��"Ot	�Ec˝5��<��BB2'����"O��	 ^$��TY&�V�<��7"O>��$��$�>�ψ�KnxKR"OvD
���*w,�)@'�97�j�"OX@�C�%t,��*&a�4TQ��"OD�ЍR��@+�bù'&]+"O����D� r*h(��!>S����"O|XE#Ȯ�ij�.C=NN��(�"O4�8���]��Җ��5B�<�e"O����ņc>Lx�rk�X�p-�W"OP��� }v�a�
ޞx�9�"O!ڲ��#O�`5B�hF�<c@���"O�l"� �$"n��ҧ�wa��%"O��:�I�n�t��@�L�]/�0��"O��V��'5���&��2%���A"O��.�,��5�O$i8��@"O����+U����N[(X��@"OP)��&XP_���L��M�噖"O���EFW|������T�&"O���#A��x\�C[&��`p�"O�9�d��((�S����N�x��"O24 ā�9ϼ���ߣ���f"Ol�*E�B7N`�1	&
�H�#"O` ���-�ҩC�֢0|D"�"Of�u�'-ض�g-Q� "AҒ"O0��BE�?KVv�ӕ̘�^|��P"OL`[֪�y��u��KĨ�
�B�"O����͉+d��i��Y�:���	s"O����엋�\!Bc�(�Ψ�0"Oā�Q��Ȭ:���$�(��"O~ݺ��N.F` �a/,2�y�D"O�eô��)Q\���m�S`X �"OL��ԩR�f	�p�&4P�"O4�C2�nq�!cS�ުdI�d�@"O�a҄b�,Ma�P�&Hu*���"Of�
�ǝ5w�V�r��
D���1"O@1 ˕�b�R�cE�QJ$d�B"O�TqBl�;Qߴ����ܢ'>�L��"O�i t�X+NP�`���P�$"OF쀇 k?4�(�Ē7!^��v"Oz`�a��X�pM�&Gx
�yq"OZ�b�ΘyM�Y����Bl��SW"O����+q�PÀ�6̘�Ӱ"O��� �&,�Bl�#/�$�M��"O��r�+5R��`BLM3<��=��"O��H�J�ܚ�d���Ĥ��'Ӱȸ ^���<�E��$��a��'������,�N�b��$hĊt;�'XaF�ϧ.<���0��W_�%r�'����e/�9P��{�i<T�
�'��Y@��K���"6Nȋh^�,��'��X��J��^Լ���%�].���'.��Z�U:�^= r%ܾU�9��'��	������sO8N�y�'�8�s�4_�x�.�:�b���'��ع�� v��PK�ME���
�'Ն����m�&!�I�o�؀Z	�'�^�	�:���;�F��ib@���'���@#��w���� 	�Zz��	�'sNɊp ���%0d�)˚�-D���fI��O���jէ��QQ�-'D����M<7a�X�#j�7w��0���"D�� � �6&O2-��C�E+3:�(F"O�#�O�P���µ�"p�TBU"O������(�L���aS6z�t�a"Of��W-Rj�L�g�y�["O��a�v`yу%[4ڡ#0"O^=h�.aS�,�dFF�S�4��""O"Ip%�,t��	Iw��`�"h@�"Of�@"��k�p�P�ߵ�*lh"OF�	1�^;F-�8�7 A�Ne��"Oе"�E݉8B`	A�lJ8J�4�3"O�Q��(G%f�) jZO@�x�"O��Q���P���b�N&�xq6"O�)S�=;gƔKA'R��4��e"O�aP�aC�t��� �6<F�\:�"O��(P�ؠ���R�S@d$��"O8�cpf�9}�8P�F��+(�Z�"O�tP�l�4=�y�u��".��"O��1K���� �z�IS"Oz�:�ȏ::�Z�����G�P��"OL�SM�5����fCR~���"O�
g��4s�E*�o�/���i"O%X±}��SS	�j�$M0�"O�8���.����G�n@��"OR�@wMMIr�J3�պt���"O��[��Y�3�x�E�t� -� "O4���*�FYX\��BϚ/>����"Ox�j�H̓u2�a ��s�"O8�r���*7Ǽ]y6�����z"O�Y�5+g�����Eҝ���е"O�Ys�T�c���1U)�=Q"OȰ�է� *h)���]�ljb��C"O�AxQ,�
1�vYZ'AZ ^^�$�"O6�XR�Փ#�QQF�İ|!�`��"O��K�O����$Ӎ	���۠"O
�W+W��]�.^�$���Y`"O�Ԡ��A�9�-��)Ag�\��"O<�QT��j ��`q-�6��j�"O�H��T<���w*��{lr"O�� �%�6u�J��qJ�<0���K�"O>tI�HҺs�V�"����|I��"Ol�j�)0w@Ӧg�Pz�"OAj#
�����3ㇽ�NL�"Oh���_r'�����=?x�h�u"O2$�ócf�C�"hf��J""O�9�',�:��8�&b�T	"OhL�A�N[@zA�aj�MUfI�"O:L�$�2C�Xi�D*�:7G@�"O�ٸ�#�~�l}rQ��u)�ض"OX!C��ϫX�2��#���$�x�x"O����s����S�|��mõ"O8h�0IāOJ�h�f&��S�`�1"O"�`%M�d��M5��	�ȅ9�"O� QF��Y�}�b�W�-�T5�"Oֵ�& ��>�1FW��� �"O0A�S�Ǌ���"t��R�i3"O���tm��Ut}����U50%�1"O����$d��a� ��=!��"O�%�gn�yo
 �@��Tu��"O6Y3Ɗ��y�å]�7��!"Oa*�Y�S���$���l-�"OJ��W�Q�aʼk��r����F"O�C4���n�:v����f"O�����>�
8s%Q�6���8�"O$�ڀj�;m�Д{f��K���"O� Є�%HD�Q�%�	e]��sB"OZ1k,�~}�0#�%�	E���"Oꈨ�«;Y��E�[�7D�(1�"O<���ź,���Pd
�lQ^5Y�"O��z�Jb%߸u�X�+�&I!�M���\� �Ύ����c%Z�O�!�D�>���H�HϒP�8\*##˾-�!��&�d�?�ܩ����!���1w�>ܑe�H�4՞��s�\�!�d�+t�Lp �/,�D!�!��o�}���a�����-�!�d�~"l�Q�ů>�����;U�!�dB|R����G��jBg��Q�!��=zB=3�- N̰�CgeH�P�!��	1>��*(��F'Ռ	�'�vaZ��J�,E|:��������'6�-�"νZI�|c�D\�n����'7Nl����e>\("g�	�j*"���'�89d�ӈn$�i)�OS0��
�'ئ�G�� "��9Te\^��:
�'Qt��5��$x@�X�c��RT1
�'�x� ���)��l�R��;���3	�'�hA�Ɨ�b�	��u�!��b/D�� �Eտz�8���"W?��M��+D�p	u�ȡ�ʍ�7#��6=�Q�@�*D�ē��ɂj�d�𧎒�+��1���<D��������h���JZ��je�'D���r�X`�xhbI��V|�J�A)D��B̝'��i��\�j�u��G,D�����A�;��H�F�ئ���	7D��2S�ٶ:N��R#����� �6D�T� 	�M����K 8���HEF4D�<�0��(��Z�"�9 �S  3D��a3
�B�⥺�g��8-Z�XWK;D��䕪k��Aa֏�A�F鉂�<D����#��
ơ9�ܙ��P
�l D������:�H�c6��,i��*CN>D��چ葨R]L��� �j��q�"<D��H�fK�ar�ү�8�Di1��:D�0Ig�͙=�8
P���{�-&D�0���\�G�i���Jv��Ua7D�,���ڜ�d��k(��:��9D�pؗ���z�� ��GW�R�`���-D��a��]+c�:�K�AH�������.D�( m,Pwl��C�:=���-D����E��EG�1��;F�հ!�-D������6(���Kg[4��1�)D�tE�_2̤�#�p�K�4D�̫�#�^���S�ɥaS�\��2D��3$#^��,����iF<�8�G+D�tQ�/$|�x!6`�)��p��)D��PѡO�3b��[��;l��Qr�'D���s)	�=��KF�G�@y���g)D�L(�G&Lx B�F� ��陖A2D�8�S��Ylx�Ad��wgҍP��"D���@�J6Ti }��Ķ{��
!D�P�J�IN:�a!)A8P ����+D��)$	�)`]������ ^��ix��5D��k��˵n��" C�;S���T�2D�܂��9s��T30`;-:%He�1D�`4n�e4��]���d�tA#D���W���=���Qj�c��P�- D���ب<NX�!�#�0_�P�=D�\KDA�;]���`DT9(�0�g<D�� ��x��^�-T`��I�8Z]й�6"O��{������H����PFt\8"O��E)̯t�N�*s Q&?���"OXC 	7/�j�0Aϒ	���!"OB���N~��C��e� ]z0"O��PD��W�~8���
�l�H��"O�$`��	�%¢��=J0H|��"O�"�N�	�F�[�Z q#��"O���2�
-�ԅ�g���"O�� c��E�x�;��Y�P�z�G"OR��T��<c|��F��ڀ�T"O���L5E����5jڽqF ��&"O�|���_"�K5�G=,�@�"O��k��e�^�32j^��+2"Op,��L��d�lA��k�7r""O��;q�>:�p��$��$����t"O�`H�(tLVY��#�I�P�c�"O9�d`Ђ��\��g�;�ܽ*C"O�(�U<�0�ufZ�a����"ONUP`�X�j��c��7���B"OHha�DzΤ��X4K�~!p"Oj�Ǝ^Lt�����͜Nu����"O�8s�,�@EF9�����d��`�"O���'
Mv����F6fj�,�"O>�H�c�;��Ĩ���$3eP R"O��(��:3�����+�p^�=��"O^�2��Iu�ث�J�?\�ц"O6� d��4J:%cI�/,VTR�"O����3#֬�A��(H4"O���R�W?]1��D���zl�I�3"OHt�@�ξE��IO.Xg2�"O$PJt�Ք�\�Kr(Ӓ(g���"O����A,z�vi�"e�"p-A�v"OV�����X��΀�L�C�"OH� ^�w\va���5_D8�2"OV���K��`�\�#�A�Z�	9�"O~�k���*&6,�)�/���r"O������|-Xsh�]�� �"O�d���PW��˴i�98�p�"O&��`Z�H�xj$_����"O2Y�K�L,X��h�0�zy��"O�U��e��&U%"�쉱�"O���K�t��EıT�L=@�"O�|)E =��X8%�<]ΰ��"O`�� �I�"���Q.�*8�DA�"O���wh@#FV�� �ƛ$EjH��"Ob�a�I�$��h��u\�9��"O�@ږ�=|��CN�;t�F|��"O6Mc�U3,`ȩӌ�?.<|M�v"OP����  �5LI6-�2�p�"O�Ĺ�R��/і~f�#�F}�<)ċŊ'"1����F�m��${�<IB�Ҿt����7J@1�t1��Oq�<1v.�{d�C,��s���YsM�Q�<�j!V�Pj��<�vI#��	V�<Q��<!h�rT`P�H������R�<��ښc����JV"Od��3��Q�<!bV#<��l�v��,�]0$�XJ�<AD��f�,<�%�d=�����C�<��d'.n�B�y[@�s�B�<���
5]�6C�k��F�R�P�_G�<1b�Y�w$j�b��(��D�sh�i�<��T1_��s���`���@�}�<Q�K��h��Rϒ�o�D�(!��w�<� .M��kϾoYذ�e*;B�b"O}�H`TD����4�,�'"ON	��
�{��كP	�p���"O\Q�i�"�t���(��El:tZ�"OS�B<r#�������٘�"O&�uN�M�&\@s%T�h�"OR�s��R
 �����\�x�B�"Oμ!��M$\:�yj���,:��cw������)�'b�.�z��D�5E,��U�T+-���ȓG|����@6��!ʉ�T4j݄�d��Ց��L�Z� �hC�� ��لȓ$P�h(�C�����*8�����m~�`�I	F���{Q�O�k��y�ȓ/�<�k- v��Ce��$���ȓ�$��`��C@�to�YO����v'�,�!;[,�cR�L>j��ȓ|�Zݺ��: O^�Qa8Y��=�ȓ�~L�p�X�f`@�k��EP	��X�'���ˇ�ދf>��r��[wߦ@�
�'E^��I��.�x��&��kl�i�
��O�]� ���;����t��N����"O�آd�T�#���IA�C�(���R�D.|O(9�e�(,�����F�M &��W�Ix�P�֪Kq��ՒػHʂ��  !D�01�dJ$t�i��Us:*��b;�Ox�ND!��ș(m�*�r�'J�'A�����i�'������C(��L�doת,��	�'U&К�Y�F|*�"�.�9�'~.�sDE�^@ �
��Jh��}2[��D�4�;�i�ω5.ot ��"F4K��l 
�'��	�0NޤBDu
a�R�={���'�ў�>��60O�l�vOύaB�PR\�Rh����"O"=���Ʈ&)~|A�/r�(��U�x��ɉv�*�!�'\,��h3�ӆ��4?�RK�:Zd�q%^"2�]
�K�b�<iH)"�U�F_�R�6�P��c��o���T��<s +؞]��@�MXvHqH�H��<�N���뉃_L��*؛g��Tr7��G��➴��!<<O.��2��gdİ���50�K�
OQ(�(�(���P3��Z��� �?�O��'@Q>y�w�?%.F�Qr�W�"��sj+O�P���^Y��.3����P��C!��K3C�Q�N߹��j���<J�'2\��=i��)_�#"���نiѠ��� \!�ӵ[��q�BH+�lpG��
X�!��W&Q.�� �ѱ��x�g�G�K!�D��*z�%�6�%RO������tFbc2�Ӻ��G"�2`y��֓pTI����<�a{��#�8�N�r�AO-x<q�֧E�?�C�	1��]"��1rY=����n��#?���	� �҃4qn@��C�Ŗ��D"��OX�X�G�6�Kǃ� �< 1�g6D� ��gìP�n,�!�%o��آ�2D�̋�g -�d�XF��>p8ё�N$D����*{隬B�#}�����"D��rt�w|�|X�o�8>�Zy8��?D��4��/WBp��	� D:6�ʷ�<T�ܑB֠a�y�V�V8�"��"O��"RE��4o�(Q�2޸��"O�-R*��c�@{��~�VI�g"O�tp��3���wN���{��'�S�)��Mנ0��������!�dD�Q��T`�ł;%B�r�cAz�!��� I&Lm#$gZ�z36`�'�έo���m�RY�y���� �mk��%�����y���9�"O4�J4�[6LQ@�T�$jc�]2�"O�p���PZ�z���,U�YM6��E"OLA����
�J�p+%5(&�A��hO�	�I&
�HêO0S��S�c�#t!�΋z���#�+vx����H-k!������&
`$�ba��W!��G�l ��zM� X`��?+3!�DA��p��<1(@ie�*���������;�IfVaa��'qTZ D�[r�=��+!�,�4
�$B2*��v��Gxr�)���)E؜!9�/���Z���e�<�'$�*zY�Sh�AJy��c�b�<a%�`O��b�&�\��D�`�'��?�	&�D�|�9I�L>b��� �x����@���0"�ci��H���h\^C��,-�y����`yl����L5B�I�7^~��(L�vV�B#�$����o}b�xRW�H%��]mi���ܭf��A	WHɒD�B�	Gn�a�t��T(UKBI�u���l؟���^2ϸe���P�
Ljѫ)��刟���B�P$<�R���`V��6"O���nN$_a����b�>Y|��0T� 
aX���O�>���4�ٙ!	,����s$;D����È dF� �ǢS8�h��9�hO���_!>�x���'@-2�YpdABxC�u�p%[Bȅ�t.�1�-@\<��hOQ>-�!@�*d��w�;R���eh$D�#�¹X~N��Ek�t8K��`��&�P��ɝ4��T@��P'g��@S$$�'���D�<	�� �B������P�<Yq�
�,�I���؅��0"�^�	�O��)O�Ϙ'�6r�l��Xm��2IA�L��'y���ʂ2�(i� J�Y���+O"�=E��BR(�(�d�E�{3�%jU	���yR��1���5K��`A:ըL9�M�1�:�OfQð�9I�h�#����3���2�	@≵;1��%�4Iˍ;��HǬS3D�~\"Ox82ej �'l�a
�K�hb���'�qO�P1�O�/��tX`�� ��lk$"O�@�f�X)un.�C���5j>mQ�"O��٥� H��#J�'s�2䱐"Od��1 ��z1�@w#��:�e�x��'������x�P|b2 ͳ=Gb|�
�'����,��)3�H"sɊ��Ԑ	�'��<���+���p�㖙EBn	��4�?q����iE�(� 
9"grtja.ֽ-Ԝ���'��L�%��(�x�db�>+'���'�x9�6"\�dƹ���(�e���D��u�S�Y|z����|LL��'�T��ɀd~�0��y�L}��ORVB�'�a}���n�B�#�"�����	�y�!�O�����A��Z��C�����$.��i�U��@"cK�&t�H�+�	!�dU�=��I��ɖ�:	Cd�Ԓ�PyB��}h��0fE4T�hi��*�=�HOL��$I0K��2�A�(0:g,�+9zB�| �H��-�4`>4t�D�h�vB�I)V�xx���٥{T�0#b���a&O��d[�w��@�B��@K !�Ыԩ#����'x��D͡լ�E2��j Ep�zQ�f"OŃ�Eѽr4Jh�vː�r�ƅjv"On���%��),"ݩ�J����A��'cў��'�`�4�N�I�. `�͏$kP�	
��� LiZ�`��8��& C4rV��ɂ��@x�$��ק[��M��]��b�yQ*O ��O[s�8��F�6ˬ�"O��Qp��0RX�B!�1��m��"O8Mc#ĸQb����L
36H�"O<�9w#	���;���=0@��`�"O�@R��%74���WEa�j�8`"O�Q8��̈\&d��$�R���)�"O�`p�=�$��E��ch��+�"OذSKN�{,l�PU��W9��"OHY��m�j�b�0����\�i�"O����L�Q��`{&aG/6)�@"O�L�!^���h� B4l�:�"O,���E>v`:wτUTب$"O���4.Zl�Np$m�P��(�"O���GGP�.�I�mгz��8J�"O���쎦6�d��lƌk�H<:�"O�4i��ݻO~��Zu���,�e*O8��@�G(\��d�߱nHT���'ˢ[ե-9+(�񣤃�e_l@��'U�h��V�L���r��3VU���'�d��'�I#==���Q%�Q�2�'[�Y�PF�mʨI;Xn&���'*BY���D1@&�\b6�B)S`�	�'���kd��@����-P4vj2�'IZΉ5n�=H%A��	Or	9�'?4uZRl�	R1�S�|��UP�'l�b�yP(�ss�Պb���r�'�Nٻ�'�?L}�b �� 0Z���'�N$MݿI!T*`�E�����
�'ȁ���ߨ�����T��6m��'T�`y�i����@�l�-`�,8��'X�!�ʏ)"U�����ӧ]1�0s�']����Yq�!բM�S�ܸ�'mqM�1X��ԂěF�T��'~���ƄR���s�j}��'�x`�@g,?�TIH�o��-l��S�']�Lc%-� p�� 4q�`���'"��:qK��s�i��A<:�B	�'!R�I�=B�0�а�.4�tІ�ə_5v�ra*N�Y�h,A���<l|!�V1N\FC�I�ph����n	3��s1��.1U�B䉤P3��jE(��:5X�s
�.YfB�&/\��6C�<�Z����[G�B�	�K�l��!��#L�p�fA]�6�$C�ɲ(Ȃ���R�4|Zq����.C䉯J<�����#����ЅM�>C�ɴ^��+6��by�E��Պ0�C��@�艛1�B�9@�$��J�9��B�I�U.)��-�-Mq�8��L3l?�B��4gb"l3qM�I�����$��R��B��!mh�mV&��F���)C8�B�I�/	HRW��"t�\Ȳ��# ,C�ɔW���񁋓z+̴8�	�g��B�I.a�&�K�Ǔ�^�웕.�J��C�ɺ> ���V��j������C�I�'\*U����� H�#��o�C�	+?mz�Pd�0U� �'˼[~�C��0A!�)�8?�p���I
`G�C�I�c̹�TO�6�"bUZ�'E|C�Iq��IH��'=�$ڐ�?TB�I�$7]2�`ݲN`�*!)ہc��ɑ�}�I�)�']�^�!���->��|��lh0��hN���7g�UвY�B��ڎ�'PI�V��1{�`+f��� NMѴk>�ı@`C�=E�Z����'�j�`�k�(+�|�X�B�%�����c��$��'�.p���"lgpX�!��%����b��S�ޣ<1U���na~D�Qc�'����J|b˰;����'\<�<��KUh�<�w�߼Qb%`�/�+lJ�:b(�.���a%W B�R���$-"���F��'s��zք_�m���'A�l�]��' �hY"]>kv�Չ�H�I�J�CD"��D#�����=������F �lE}�( p�͊��.+?d]�J��O�@�,X*쪲㖴C���(sH�u*8����w�9s�F�3RmL��R��>���ɰ3Ҹey�Ջ5�Q���ԋr�T��ۖ6V�@Ӂ�5{�D�g�ղ6٢Qs��0�E��?q�cD��B��ҧZ>izabU��~�<Q"NC�2@z�f��T@�q�&�$i�.g쑣��U4����O<j��/�(����O洉dSN��;�+	�bH�����?0&dz���o��P�Qs��OV�З�L5"��=2"�̥(,��� y��|s�ϛ�%��p��`�MS�H`�	ʙw�|4��.�1z�`�jv�L�`׬ǃz��'�P��Ɓ~� �Wφ�b�T��D��p�b�'�T-���3��ǉ��1z"�۲��#*Z�OԘh�K�db��'�3�t@G/�d J����u#�j�?{p�:@NG�a��' @1f�2�ӷ��-�p(6�@w��sL̈Q�t�dM޲$�8e�W��e?��ě�i��9���?�,��� m��E�a;s���E�݊*�^!��ݗ"�#g��2\�̽�8��I)�aC9v��0�կ�)�N���R	�t�T��G�B=2�΋>xF�2��O\0�t
��t}N��S*�|�I�EK��i�G*^�h��K�A�Bٹ.�<��+!O
4{Ǭ�AT�U�|����8��@�G�
�E�X���nq��!�J�θL`rEW<_�-�B34�(��F#^d��u��by�'�H���֪C��y�p�ހK'P\�1�I�[�8�V�V[�\lU�L~\�;�a
j�d!��.���^	���'� ���ב^�t� ��yZw�}��mW�0Ɓ#� �&k6���
P7�x�z��]�dFM��܌�M�a-�6̑;� 5�;aVx s FG�E�������v�iL�� �M�L��w�զ�S�	f��*0�^���7�F����
1�E�`��.Q���tfU�弐i3��$�z%�C`�ʛ3�mѰ(�V���q�f�撝�D-_�R�!k�^� E]��i����@�R�e���� I#-�ta	�~yҏ
�'������E'm:8h�m&\}�A%��@�b�� cÇ�f�1���S��+�*-	5&Xx0-�&XE�q��@�lՂ�#�<��Ȃ�0����٫8`t��j,:�"[�P��M)��4Ґ`�E�bXPv*O�橲@뎗b�Y��᜵_JD��S���t9��7y�i�e$E=;M�T�q���a�� +���&⟸�1K��QS�o���x�U TN�L���	]�����F3[ H���ԹH��I{��K���;ճPq'E�j*!�蕇�bA��Z,s[j]q��ғ�Vm�Q�W5�b�W`<�aH��r]ϻG��)Z����i4�Y�qn�M�L-[���#���'�6e�$�r���W��<�`��%L���W�P,|>:���Cٸa�@4	�(��R�G5��[`���d�jB/y.�'<x5���]�(H��	�> �40��2Cdi�c��h���"�I!h�9d�9�p�&)='��H�ן6KtE��/ n���땨�90;���RB�bDTLx���>Z�Ĉ#�#�o�I7|�
�9�]XN��s�H
��|�gp�c���-@�Ľ��P��ht�#nZ�7���J4*ݨ}5)(�G�?�!CڮE�ҕ����9�9D,?-�6qq��.0��
��'����r	�7�|��	.p�=T��l�hm!�O%Z�,��E��x+�d�F�&�m�%I�\ua�7��?i1��[�Y�>ē�'ч~ ��	?g��蹣���k�2�+�a�l���'��m�w�~�Ӻ�7�ÿ<���',�6$Č�� �<����@nHl��\!����(�(�c�\�� ����0(ܢ>�4b�0ha\����"�+�%�h�p��r��&��iS3*T=%v\$��\�/yP]ra�'&!��HAn�M������
[h\2�����~"���r=�o!j�p1`R�$ ܱ'-֑E�tQ��⇎8�롲i������.`#a�Ƌ���̻s�I�u)J!�1��G8�Ԅ�l�vɈ�I�)e���̃g�jȠ��V����R&�/
�� V�Gl�~ݰ`iK,o��� �M�b�|���Wo��x@H��i��Bp�R���9��4CV p���T���:�o�0IZn�RfO�5���b͙('�0�D�W�`��ya���)ڊ���ɲMPx�F{���gD�9ѡ@(~���J ���'��噕
�0/trA��T��'I]^�
 �"'��L�3	'W���ތW�R�)��94��eRU�?�O���B��X��͙�R�h4ɔ��3\'Zm�E���݌-y�HGK'�	���6_�H혒Q�j<��2��Q���Abf	��뙵����"O�99�����0i*�(])�j��#��4�m���s���-�n��	�1�q���%w��ٹB���=��5mZ%E&�a��ͺ1� ���f�v�,pAr$�G�ܨ�H Xh$y�����I�ER����{�0B�����zG�	7k騡���=g<�!��ۯqވl��ۨ6��������Fz��h|H| v�˧r�����D?V��U�Ƨ�a$�p2�n�>�X�#EoޗmxDd ��ʥu��Ի n>S��q�Fa�+L�@��1��ܘG�(B��Ja����#=�լ��hld�;��a�)ޑS&V�c�dAI�K�:lCÇ�;c/z!H����9�Ԉ��2rڅK޴$ژ����:a�y��FϺs��q˰���<ؚa��ē�R���Ԗ|��S�P��ؤ&�6����mY�*O0��i�Ln�uې�
���Q�ϗx�<e�&șIg�Dj���D��|�'
o���񔦊&��ado�{�4i�v(��Mm�ln��I����{Y\��̭VP�����	�|����HH��
�E/�E��IF8y\V��DL,VS�ܺql�	)xP��k����t�N�gDp,�P�f���E
�Z`�ç�1&0TA�3�6�	�cC�z�� R���+n�Ո��Y�;4���7�J"25��2�I����#ލ~��<2s#�O��T��<8���Ӊ�F-����|\Jga�?�b��A�1ʓG5���ͫ�dp*�!ڎ9�� T4x��:�Q�)pb��ŀ �:ݹ��R�U��w�0 �H�$!� %��+vr!�P�#��sBo�53��1aږxP���3�xB�Z5.��8Cǝ�eC�!�b�G:.�m�¯��7u�����9`Ƣ1i��E�( ��	,�ԙ޴'���`re�6?B�m� T;wʘm+Rȉ�$S�1@�	,b����Z�Kxl;���4V*�񊑀��N嶅aA$ƵvD�h3��/l��$��GnDsGD�4T#��FL'8�Yf!�il@�m�>�<��ҝ`�U0Ƈ%Cބ��a�S�'#.��r͙����s텤Z(����K(*ҒI��L#>�P�(��t#�A�{��tS1iv���j�n����a�¹M��a�S�C�s$p���'�ʵ�"��S�^�B��H�{6z�b]�[�8�8��͎Ff�t ��� �����Bg���x��Ά`ͤ��!B�\�*�$�En�Dh���(�%#�.ے?V
Ex������h)�	
)��y oP�an�MR��#�Ը�`bۙ�9a6FܴVm��PoJs_�q 'G9ua��i�E@.�5�?97N�'��(y���T�y%L&N����>�PyD�kX�D�t+��L8�a,�E��XȆ��'L��ȃ�d��pY$Ȯ��A��]��k���.�^��#�9k� �e ^�p��2M����<�E@ٻ7 *`h�&�4vx�5����e ��k�d`@hC��_�|'b�P&`�:5&$|Xf&�s�7�,�4K�F+O�Y�W�\�x��|P�`� ZazBn��r~4�[���
XpAr�ͯC� Ao-��	���<:��jQ������Ƃ %�D̮B
��g�QEjx�� �J8
�=zT��!��5�K�����=^�y�(Ѣ;�H����P=^X����k��3�ĺy#j��H� b�$��4te�'O�)�����
�.�Hܓ#@L�D�KXGDh
@	�2nx�B��H��x��ħ��,[��A"�Β�/j	!���$3�\�a�5�P�@b�,�����+K��h�3%�������伺��:2ax2ƣ5耬�*��8
�|����DM.R޸�I�dB"���+A�Qڟ�2ݴ;�`4���y!d0B��φ%�щ��
�@aQeΘ"9�`H��1\OV�#���?���@�-'�QI�c�i�*�*�㕼t4�ZR�[�M�PMR%[�n��N$ZJ�a��lG��,A��NF��T�V�?^�]�d���M4�z�@ax��j� ءN�`��q��L'�}j�c�L�0:�k��Ʃ��bZ�8���$���S�����ܛJ,�Y*��\�L�<���<!s� a�T��)L��~�aZ�'�Ԝ�&@2E$̩����P4���j�����V�t8i��M>""��8�f	����)h2����Fxj< 3���+�8�F|r��]XF(cE�Ӯv�pC򡋝��Y����U36�Rw �"����jX\ZB8K5���s�T����u�5*�vQ�5 �&9P�9](&�6Ű��^�}b/�4m��<2�'��K�tcु��He��)�"3x��dH��Z����U�n��Js�K�@;p�@	�y���`���u�]/�NܘV���0>�Ub�5A$�0���2%�Ȭ��dM�M��E�d����؅�I�2j�0m�E�2`BY���Q�DDn�T!f��@�(T*�ʘ9�J�I�q�����BA�������^h"<9ᫍ�J�,�ɳ���b��ѧ-���.S �𪣪�J���y�@z ��Md�9�U'x���g�#!�P�$�^�'�� a�בX
tp�$&�4�Zu�X��j1�u�F�JiQ��I��!81��[`\��е1�NE�D�ق�Y�5\��,
i�6Wp�����p�RE���''��g-�4/���a�$u���}�0}����<+N$y�gЇ /���ߴnR*�ᗅ
#G� ��4�"Fe��s�b��g�Tqڤ����'�̜���#�%�ҮǒC$���oԒY��l�щE��t 9t��/J�B)�E�˥�F(Bq�ƐF/���t/�Z��x�QɄ#����||�Ab9�wi�0��$�4 ���#B�	;\�awT�2�$`{ @ɪF2�uy�A��tT� T%&od��`o�z��QMF�ER}:RF׋�]a�ɚG� ��'K��w��I�1�Md��i��/y� A*W	ޖ���&(��C���w���r��}����� ���N� q�ʌM�m��BM�Gd��d��1a~ҁ�
�zؘd�̻t*�X��K�8���F�O(ʄ;��� ��pპ�j��t⌸r!�%@ ��y�ݦf�@X!�aՒA���s!)���p>�2��%*�(�y�Iم/��-�s��yA�%yDhY�EtXm��	�!9@��7D[B�����T-��1���	|K�94ș�����f����S��*����@�J�9��{R��/8�HQ@��^�<�$������S�U�b���4j+#tT�HS�H�����+эL���r�ǔ���E� Rf�ۍ��ƦT$��@�j�Hٌ�r��}T|U�wb�5��5���X�%|�4�_�8�c�Ɔ�SÌ]�6�U>k��2�?if��e�6�<�QQ�Tj!ӄ�L[£>a�����z�`������˱{��3p!��I�l;�i�1��0�WNK�
e҄ �7r�\Q s�
�}��s�$H�`�i�4��N9�N� 5�!ecb���|k剌�����4[��T��s9��D�-��=C7JB,@��f�M'"pْ�ߣ"4 I��Æ/i|5��b�+��z���5OH8d��O`*�i�/vQHBh1�~m����a����C���wk�����W:�<Yt- y���Q`R�J��u�bM�;��SB�M��e�0��5)��s���86) ��i�	��U��}�)�,dҶ,07DT�rR4:�d%+�� �M� vIPi��"JXp�����2��pBzq�E$"��Xa�CsA^��d�? �\ �g@��Rkh$)�,�:H���#P�EB�`q�	�Vb�?	�#���g�I�Cv�jÎ	T�5��4|TN�yԇQ�2� �8U��
-�u�g%��D�*C�P �!ː��6y_V�)DgO9N��� ԨM���`k��L���y�HMZgf߃]���X�ǜ'^�ve�Wʔ�rn��'=�0�r��9]-��oX�hgH�i�lQ��Y+���x�h��ff�d��鱪\�v�N�ѧ�W�mlR�6,P���7m�"Ӳ�B�� q%d �򎗮6t �@�[/u
�0�,�h��ןx�k�:?\g+�8	Q��!C!JΔm��L[_2L@u$�K0,����$ZƢu���QL �TB#I˘c���B!L��<�L�1zK�U8�Ιz��|Y��I�K��8��� ���w
M�D���4L�|G�E0 ����%н <�P���	�`)�G�m���A���#VZ��@�V��'W\����׀y���o ��x���+�:��MO��Q�oF�l���âo@!3>�����'�j��f�>(�(B##L�H��yZ��F�o������ � 8$DE�=^���BEV:.$ձ�S���5E�,�V�!��O���ɟ�Y[H�Ȣ�D���S�M �S�%
�[G\�	���i�`X�g�=AS����ub���fnM�K�E��ZDT�9�ތj�hT�Էiݚ�s�銛8F����d���SMI:5����!�..U��(�*�)?����XS����Py�!Q����e 2� ��L�I^@�!Ă2 ��sf�C6�ؘ�TE�fJ:[ �>d8��=�&3�B ��	��] ^���$m�v��-�2:�,�%�Ū-1Xq�f̆{�N4����]\��R#զo�x����1?5�RlZ��k¬�3n�e�ѡ)��n!�	3Fh��"$�5�f�7|1���y:p�c�-K�������qL�a�'�G8�Тd��mm� Gd�ug7�<�҆K[���ڢSb��V?A���ŉU����
 A�듫#�TTs� ;�8��A�:�'8�T+Eb\"g���e�'C8�ђA�Q#�9�!fI�Y�h��٭�H�j�_��a�쒢��A�C
;��t�ݴ?N�Ijt��:j�q�uӱ�֤��*i��x�A�&M�5a-+ ��ڠe�f6�{�d�T�H�"P�L,_l�3�4&ʭ�gM�W`!���F�5Zjqz#�\j?�=?ڌ��k3��'{z��&5$Ρj���(P�bO��qJ�4���D g�&��Ш"lOܐ�Y8d*���;������?A�֬b`�'@̬��K>i C'Aͮ��O�A��O�,�ڱB�E�$�I��ɱi&�B���V��<�vaLM��O���&��-@ʖy���<����'<zYQ ������\$'��Y�-O
�j#�²s����N��|G(Y#t$�8���%$�(K�lj�<��;h}H4��)�.��Jdlgܓ_�n-"&�3O-�"/�UJ��@D�#@H�9�"On�U@PMh�
󁑇&�9�3"O�x r,L�GtfRQ�x{���"O�X�RBF��aG��XܪuY"OF��B	Ϟ9��%�v-�"O�pq���)��l�eN؎{��)"O����<,��A�l(N�X��@"O<���
��Z؊��dϱQe��"O��fe�����c�-Yݘ�"O��w�G*���w"\�P��hl"O�W����ȗ���h,�W�D�<����"+&���0�����F�<iU$�)V�A�$ثiOte�G�v�<�#��8>#�l�c�l�� ��H�p�<q
/�)��ϪvB�����Uv�<Q�e*z�6\���YH�r��@�Wt�<�c�ǎO�J�Z���*~�r�HRv�<IfhԠ*#�!� M�h���"���p�<	�� �BD@H���0d(t6aV�<ѣo�D���M�2�h�f�V�<�En�\;M'/؆��qЅ&�Y�<q�I��u|:����8;l�7KR�<�u�S����O l��8���LH�<!p�j�v��Pχ�**2ܱe*�F�<�L�$=�(Xqk"[P�u��k�<���^�D�X0C�ŻCm�.��0��d,�a���P�PRŰ@獺M2��ȓ0��U�BR�S�2��C̕5~@r��2��耥���C�L0$�<�$E�ȓ.�HU@aNR�D.�3v,�4�ι�ȓ8�	��
X�}�}�����9�ȓAT�M��&M�.�ҧȎ-,�p����Pc�b�W�t��a���8>���ȓy�v@+e	ɦ`�B�P�N�ȓOF�%���H(i�
5�b��� �ȓ-��Tp�)L0VD�r�J4]yF��ȓr��Ȋ7O��7BR�S�_7O
��7�� `�_(�CU,_�j���C5t�����0�#Dn�.B�hQ�ȓn�V���NB.�kB*�k��ȓrB����X6�� #�	��t݆ȓRQ�ɐ�l_�<i���~��I��u���:��W?@a�eF�<LF��= ҵz�Ջ(�Dm��l�3IT���f@x�b����1��.��m��S�? ��O��z�
��6�JA���B"O���L�U�T�0S =�L��O��R�����O�>͚�C_�Z�4���A�-��pQ',D�K��XC��)�e(�c��	WF�<A��W!y<�͒$ܙ�0<y�J�&A��{�ՂI1�P��oX�D�v���\jV��$nķ<;�q�eL�2t�����Կ'�Npۣ�'zn�E�J�q P�j�G*�8���~d�)5�r
@�J.���7���p�Ȍ�Ao����!3!�X�B�2Fe��dLl���G 8�=Q�(g\v�F��k~�)��H؂fV�p1�EmǮ	vbkD�%D�	���� sƏO�nyi�)ݑ�(`�^ 6n�Рt�וR���3�	}��j��ٰ:�HQj��x}6G}�Ǌ�ޞ	ϓe�\��G'�3v��B��޷Q��Åi�=ckD͠��3Qb�e3% +�O�L�t�^�>���¢oO4H�4�'v�]�c�٪-���m��Hq�I�>Lp���?��ӝ~jn���K��W��%/�oq����D"L�rr!��[�d��@�3�DPb�.#�����A4N^H�!�OD��-H�A����}��,xH�t�LM���`
C`qOH4��H���OOByrLû;9R ���Uê��āX8����$�Z�}�ʘ�V�.$��G����@cfO&h����dF�VO�EcA_� I��3�̙�Re2�{�d=��Y�Pc<�;Ud\�3�I�dH: ��As�F�;Rm\�2T;a�T�HA��,+"��t�T)@@���?!%h�5t��p��T	��S�L=TDH��ɜW9*��$���ٔㅅ `��)�O��qQ
��H4@l2���S> ��4ޟ󎞉78�q�ӯj�MS�&T�i���e�tMcЌ�7��Ekç��Ys�Oۚ#�ljV�2��s�Ꞵd���9R��d���ySHJ�|z��[�'�x 
�J6��k��5b80!1g�T�F���9�� 'cZ�)�c�R?��LN�o(9�ҮY����'c�)�d�9`�hL�DnL��wCL�HQ�I���R�@P��Ď*}3�|�d%�w�R�:�j�nM���L��y�l�Q�Rt���5�Z̃��876����S"�u�a�=.�I+N��e"mF��p�x@N�M讱��h�E�v rW�<]�x� M�jk��G�O!ug����φ� ������J7�߾Y�H� L�in��iݙ�'�
$ >�τ�+����gk2��T����X�V��ۊ��V��I3Fp�k	FV�s�	H�&X5F(�M
UD��'�}�T  �M��腵O���`UdN�h�6=���v�Ԑ���Y��R �y�LʽQ��Ĉ��Ԉ�
\ ��CE�`�	M���ژO�*t�������1
�	´�[U�O�9���R-P�@|+�OA��M�C��YȤ	�Q���i����E�;w~˓{)�=��@	t����F�2k2�H��84*�v��Yj^!1K>	VnGZbL	af�0�$�s�­b�t���T�P(r��T�ͣR�@�r��2M�<I`UB��J��0:-O6U�D�\=2eS蕿R�^���J��ReH �8�K�\�x�@�.�:�6�Ӊ5�Pi� `��r�X�����ʄ���wR�����͑9��3 �*{W"�7��;}��8�S�2e乢g������-8#�t&J[/�h�a���+�̲���f��]��j�d�"�.Wf�t�ñRҾT1�M�sH1H�w�H�� �!D�R1�Q�Ňw?��!�'K1���f'.��O�y̓g$$�����:Y)�qS��� ��)ғ��H���&�62��J�� ;��q�dh�j
J|�n��P�1���V��_�%�Ý9P��qH�K� [��!��Ђ��'Y��� 9<ƭku�]�q4��Xp%��e���� U���Crd�D=+ ��_xJ޿�ē�*���=}MH�x��i�6r�I�W�<d���S��Ț� ys�'&~	��#v*�� ��	���5~�y���>g����缫׋C�Y0DM�cR5k��0�B���%#�!; ]���>E�H"S��Y��^�<}t�c�͝3k��j]^<i�F=����f�ط��&�
�z��^�j�u���бCV�d�𑱏&Q�O��#_��اu7�<(l�CR�q� �Ц�׌9^�u	��:*x Š@�Ék�`��c�^�5 Ɲ�BGQ�	�8�D}�AT�^��6J�.�6-�V"���'�XA��K
��*G�M7W�n@�f	����x��H)x���1@��z��r�i��b;"=� �� �����⍨bi��6�x��ϊWM������.���;#nȃ"�� %����e!�E0vd�%	�$՟��P�;T�"��w�L��n�)�� ��$D������su6TYdǂ��\H��/_�=�4qH�'��Eu(̃1OD7�셲�	w|"|	�ǃ>�H`�A����ʏ��
�CG�_��*����<LO����/�L�m���Q�Sv<� ���T�V�y � �E/�Eq�M{ JT�z�t�� O^�,�p$�<ړp,����]�qv�^=?%���<2N�<;/��sѧ�8K)�i!�A2%����#��;}6���	V�t�衢���4j��F�HR�~����'�V�qd�7̊�sW��e@T��+T�Aɪ, CL�<t-�t	�DT)[�X�!��
�1���#��M�gAP���whư;w 1H
�`P�
]�Wf��'����D	�5y `Z$\2M�΍>8K�Lc��'&D����;����3�63t:L
��N�_:a�Cnl����.��&{�f�a��|��i���4��IB�FhT���H7K���O�)b3*N2ZK�y��`��t��� �o�ee�����M����PU��6�Hp���^�������
S���H�$�RzX1��øAD��"�S�ԍ8���3�>�D �-��e-�
Wlp�	�9DT%�!"��V�ޥh%��}L๚5Y�#x޸1�P�����_�\���"��I<l�+ �ÎTmt�#�T��29J�͈� C�dI�)_���� �� Ոt
P�@���l��47�ZH	�$��S�	����Y'&�pQ҂�t}D��ȍ�>�.d%����H;=� xYr��&*VMz��D,�����o�'�x)�"�>پ$A��	g{�C��f$���˒dzR� &皲�!�B޻<ܲ8y�'�ex�{��c.�� ڈ�U-R���Y7 G3P@}�#���HH@�b���q`(�Qe�4;�ʔ�DdխS���qg�G�WLy��(MD����}hEI���o���q��	~�p��G�f$���
����w*ʓ|夜JU��%4���gΔ���&�*Rw�y3�c΂kp�x1�J�m���j��ܵ!=�4�&��O�<�毊�U{X�8E�������A��� nEPB	Q!�*ʓ���p[��,y�.�
V	p�S`b��r��1��J=
�<���HG=+�A�\�;��Ի�.r��+����v����ϊ<�,�� H�</Ё�wIߠ@B��^��Kqn�}��'��*�<;���kuOS<G���E�ܢw$���#�X�R�>��e��*�)��84�H�2hR�M���#cU�F��#_Q*����j9Z�rq>�*�Ű�D��ǀ,<��US����`�p�ULQ7,r���O\�Cǒ	Y&�N�X�u�R'�-?��}D�d�p�����A'H'[��mq`ŕ)C"�l	�G��r�P�u�_L��J�Q|��D}G	���1a	�D@�h�ǉ1es��˞����<	CG߯}qVlz�ЇR'�6ز8n���O�){���
>(bx!�T#��JRay�CU#X��P�G��� ;���c�|軧�g=�庠"E_
~�#�F�T�q8V�߯
%V����G<a�~��W%�O�� bD�Yd�sf�ڐ)�I���5��`�6]�BOmK�o�"i�ح CA�7.��� Q4�$�&+�7 �q jW���#�KA�Ź�oR����OY�aPR��9��QjQ��-8���a&�%��'!�%��g�sU�\H��I�=�:`���Z�Zv�Z�EH�0��,�,��)�=˕�-w_�l#�H�?�4|��;^'Б�W`��=��d��JC!2���@��zbT�s+�>�>*ϓz�IGG4#�Y�FJ]eh��လut`L3Т��\m�d��&�?,�a'��5+�q���j�����E�;���ӣ'�fyB����r��2�' ��؆L�J��]����>�����fкX��S(O���z�i/(y`�IV-K%_/6��4:O����'VZ?i��T&R�(J�tQA�D6;25ZHK)-d��ҷ'
oܓ2�P��SE�3*�Q�iыAXNe9S,U�<Sz)qC�[� �Je-� Kj��~�"I�4^��'���t����XM+�j�R�)�As����yݼ9e�>t� ���X5����K�2P��Ka�ʢ)���"��a�2��"�Xܡ�8�\J��Ŵp����R�E�&�ʢ�U�e	VX#��-f��Y.*,{axj�5X���`ƅL>1x�y�邜��$�3,c���3O�:H��3u���<��42~�e	���z�"U�%��f$ ��#JP3����6Κ�MQ,=xf""\O���F!�J��u��.@Q�V�ʹ-�xA@`�-UNR�BT��M�֥/	et�%ʈ�AV��`-�i[b� &A�+7ō�w�\�1̔{~\�Rh�ax�X�r\!sP�0rV�]�<}�A֝@��y��l��`D����R�gf�9To�=�~�1ƀ�[�(Y�!�@��u���W�<Q'�:&��q#���I d��1l�[�'ڤ�C�]Nr֘�f틧9�� �:9b�m8�!9�Lp���-9��h�bư�СLشĪÉP�b��t f!,�%�h���
v����mV�+<��Y��H6c(�-���[�~��cJ�!�d�B]"	~���uMW(9��a�	4���"��b$e9��	�)N�-�	O"7tY�	�r���Sz(4m{�◤j5��A��5O2����R�g/zE�F��v�X��$0i{BV&n?���;J֭I񥁅+P�ȧ�Hk�F���	>TAHDS�
�  ����'TK)4���B��Uj$�S#.��y@�ܴz>@HXT��rg؝�EA��&�F@�Gc�C��T`&��?����e��Z=����On�'������%~9����l<a�I�_�ޕa�"�C��AbaB)Ei��
'�~)8�H��'.p�2Tf�,v~ȍ�bE�ўPKg��$T��ѸCkU� 3��r��5usPm5]=�L�[��H�1�
}���U������9&8��"#��q}D}� "H<f��@��U�E&�YB�-��	)��3F�Nx����M
 �\�k��W �Y&G	�%�Dc��#�(��Ȭ���WVc�FL?f��)� ؖdz��]�*yb�	�e9�C�e�-RC����ت-�|�B��G@�"j���/%�t���h�|�2���!W���j���i�t]��,F�D#6)*���#�\�vV�j�l�jB�OT]ɲWz���TLA,m(�tr1�	O+
��2-�><�� ]�F<�d���)\���(Ћs@��\�p���he��L��P�AU>+hЕ3W�L�R�&���1�# �]*FJ�-�P��"���m�P1:"��$a�ֹ�ID�+��9��O��'(�A�ܘ)�F����S~V�����6�^Ay""\�G��A�'�O��0?YqA��$�Tu�$�	m�8��߅		�-T�I���v�M���e��Q�!�B}�a�h�Ɂiļ[�9|þEa�G؝f��\�C8�H"C�H!?���NJ�& h��W�FkLA��n�_����$u�x5xdF�>�L�rP�
�%
t:�ցCa^a���h}B�B�F��1dt�2 B	�|Q)C��D�]�����
ѽG`!%d��Z����}TA���c���9XF��G�O�B���H=7I����Ď~6��>!�ϷG����dkPf�,\��Q�^`pch?O�iy�iX��eGǵ@��ԳīЗd�"@�H�Xrz\3��Ȳh,$�A$��*t@�L�7�J8���	E�Bɉ�G�Xb�0�'�Tpj�o#|tԅ�G-�+�Ʌ*��s�\��'�޺�r���]�B@2GO!qЉ�wM[�(�8��w�v�@��8u�`AX�@ڝ��a�(O�!�E��jplx��!C<�H�����.��^����Ӳ^��h���3&���!,NH<1��a�r :S�!K��D��T��1X�87�ñ�~"�\�o=�� ��+J��� ��|
�m��c��PHb̄lW �ϧ�h�V	T#�T`�ƅ�>�"Q�Ј�F�ʤ�3��<yzȻG�"��aHT�͸8���0�F=9tn<�@�ZF��<����򍳷��$T5h�zf햧9Z�+�޺xIb%���b�pE�5����7`ЦP2b�2��W�?V� k�HˉL4���F�I�s�'i�����`D"Z,���@`��{&<h�lS�x;>M��E�Q��ƁB)��SQd��c�1�ȳl:���	��H�]0VN�rX�$�F�C-��51��a�,i'eI1h���c�-W���/�Y�R�;�O��r�Y�yl���4�0kp�)��*w���7F�?I�#h��*��5z����Z�>1�dT-�j!�r��'H��Ս� IN9���#.��*"�Y�*9Y2ĕ(�d5��4B�:q��eEz"$)��E �QH�B��Ҷm\R�w#*]|Z�%Eoꂢ���m�"�S
-#j9R�:� 4#g�B99{�-x�'�6-{��rq� 3ue"��#��!tH�g��cF�x̓�#��C�#,�3cc�6~��̂5�E� �I2�871e��N,_lDh��@B�&)�#��4|���]�0����x�����"`��nOJ�㷨�+�N�qA�N��^�!��j����$D�}���*Є��{���ڶΊ�F<M9�
<B��׉X(i��(t!S�`�j��D�~����Fn��C0Q9��W�G���gN�'1Gh=�@��7|>�0�l�P}R�Y5}���SA�+b���+w�'��uS g�=f��O���ٱfܬ3)�xpc��"= 
�p#Nb��Jc��0����"�-1����,2+�tP3K[�>'��@��ݦ2�51�B�f��"W�t����`k.L:S��u�U�9���a�?��K*
y(u#�0�*y�/�	t%.��k�#x@�K�'E�~� Ǣ2m�rʧ�;qt  a�Hܓ:� ҷ
�b�RIc&NL����3�aX�.�����g�!0HJ�%�ź��A`�^Uc6n������خ.�<X�A��>��Qb��ٖ�R�'���P�C��'tc��;v솈_(p{�
���)_��1 ��t����/�b晐�D��$s�� �>���"v!^	+WB�Lcݵj�|��M�GR> ��o��FJ�3����$/}���f1���iyRk-e�5��j�1��	�O��q�F*���@�
�t4tݣ��j��h�K+�lx��+��>U�;Y��%`�ׇaIp��%�5	;����i���@,H,t���F���c?U���Xм�e�/Vd��bX#6��R%%Q�ZU��zA%Ƌ(�!J�!ϬWW�g�'餩y��G�Q�m2P#�!��0K��Z��~2��f�-���S�9OΨK2iʱ&ꠡa�/B��4��@@$}�8�Ѯ��M�$@��c؞P↩� �����I�L����>���ǋ�lO$��Ę|��mM&��Ԉ�(i�ܒ��*&F��8s\��+K�p q�1�	10A�б�@R.]Zց��NE��G�2��1��ɝ,S �}x�"O�pI]�앹/ z�"�57��ɲV丌3���=��S�O�:�!�,�S���1�iW�l���'D�샱G�
N�ȇi��H=X�{"-�G����	�s2%���O�T�6�$k�0�B�	�]�6���kы=�Xu�k�#��B�I�	e���ǯ�6�:�ѲfR�C�	�^�
�� Y�x�U
֮Z��C�	@��h���Œ,�ՃA�j��C�;t���u�X��4�ʅO[�nC�,C����3�я̠�a�.AiC�5*L1��f��O�����ٻZ��C�*�ȱ
Յ���^``�)ՔO�rB�:����u&�b|"�C<r�:B�7���d�t���*׫Q�1�C�Ɍ,�0ԫV�ԥ��5����fu�C�	� .�Y"@����h4���_rC�	�xN����U69�j�����][C�iS6ȑ�ήG��]`�$��6��ȓA��g[�T�>���\��]�ȓXlt)pTJB�48��V�T�L��t�ȓ����=0�1�ǦW �:�ȓF2A�.A�H]�$� t��X�ȓv\�3��	g4!��MK�
��C�I�a���ɳL�"1����\�uG&C��BIܼY��_�b��r��SDB�	�yw��Q
��ht�q����C�	F��d��Q"���;t�Ò}|�C�	o%�Q+@M��st=ab��U����$�n�.DS�O:X#�`�&��W��0�VtqO���GC:���a'�0����}j@_�2u����!ɺlx�[%#<�� C�z�8 Q��M�r�f ��'4B��3#�Ӹ1T;�bc���K3�o�fy� �
b�\��sP4�0|"R���i��U�=���� �8"4��A����I��0|�ԋ��3T�K�E�3e5	ZݳL���#I�nH��ħN�F��ÍC�BX���W+�*H�&�Xy��)��.QZ,��UF�"���
�@���<E��Fb됹�%�ȔP?�����McSL=�S�OE�h��֑7���zGk��.1{G�ȶ �hqØ>i��O2Ԕ2c��?@��q3�!OlU�	7c�3W��$�|���Fe�0|���U�z7Δ�b�;Jo�L3�B�
+ZA�g3O����F��㸧�OJ"%	![��d�kv�� h�9I��Q"QnF:f�)��Edq����YݪQ��㇋H���AdV>�,��O�����TO�W��<!�ؠe98�Ur�:O7D6 ��)�~֧�� ��*A*��)��=cŬ���z�>�r�@/�0|��&I�C3ځ��	��a��ԡ1�OT��>a��Щ�'j� 2$�3� .�B5 X8%�DxӇnk	�4s4�O�-�'�O�H��X�.G�1��	*t
�^F��0��O0��M<E�Th�Manq)���2�(,p�+�$�y�VW�D4IHa���R���i3I=.�� xC�+;*O��Iش��b�b>k���n�nYxQ��79�j6�*?���p��䢍y��)��q@�9S&Z.c0Lʂ�� %;�$�ܟ`�"��S� ����D�b� �3��ԓNL��
�Nʓ�y
ç
�KS)�<���A8��䚄���q��I&�?�J��E�� r��ObPS`c�
G�F�i���e7�)X�"O�5��F�JI̒s$Ķr���S"O��9P� B`������< �"O�E��]~}�Ԁ'a[uli�@"O`�Q� :]D�R1�S�f J"Ozpp��t�*�rC�;)zL{�"O<T� ꛉLjH�^�	:��@"O$�� �C�B�rH)2�/*՞�B�"O�!b��lt"p�$��#'�Y��"O��JH�b�H��׍�Z�0��p"O�`[S+u�RD8�*���&�S�"O�p�C�1
�Zx�4�N�>�6�Zv"OlP�F H5B(�Ѧ�.r����"O��KG�;�J5��CE�U��A��"ONA��eD�"&�l�@c�J��!��"O��@�)B���IK^�Q�e��y���@�r�X���:x�	��7�y�&�[�Ɯ�"F?*n��U-M�yb��X�q3��ש<px�1g^��y��~z���E��ۤh� �)�y2�M
P]T\�����du(a@-�y�J��`��*��>W0���%�yb�Щ-p� J�m� �y��%�)��D">12U���y2�X���$�P��1j	���E*�yr+I�Pܔs0G�-3Dx*ׁ��yr���B#�Be��@�l(0���'d.��-ӈF1
�	����d.d[�'��� 1
ɨo���k�d���s�'�F)�� �ZT܍*v@�F<��9�'Ѧ��`�U�Nג��5D�DZ*��'	dx �i�N�>�u,R!-¶U��'.��CKF��v��$�� ��%��'��0�c�l6
�2G�UC)��*�'�n��j��5-FYI5ΗhS��Q
�'�N5R�G��;�v� �
Ǿc�pU�	�'��ȱ0��1:]*q�6(K�(����	�'����
�b��x&L�o��-b�'c�b'�� v�a�$I��4%��'��d�&���0��ذ3K(1�Y�'�¤� ������a�@�}��-��'�|Y�A�ĵ%~�����s������%�>X�Z�:�j�
h��)��,�]�<Y�eO�1�$�"7��c2K���Z�<�p��n���Z�Nǋ7Y.;�LOS�<�e� ��1#Z4A#� �M�<)C�ɍ-&jhA�#{�X�'�H�<Ig�T�6Z���C.�$�%OK�<u���驰 ϩl[��R��q�<!��ܿ2>Ցm֧s�L��@��f�<Q�*͹m���ʦJS-Ww����cw�<Q�Ƕ7�����Ũ<F���R�r�<٠�!h����M�n�1*P@�p�<�p	З}�D3N̠ܦ�2B�q�<��5`F��I�2�R����l�<��m���FD���1^t��.�f�<� ����΄�RU�r$m*��q�"O\�u�G9jB80em��%J(Ё"O>���̾J�zх�
� �"O���Ãثjf���d��6�Lq�"Od�r%�0[�fT 3ᅙ�`�x""Opաv�v�fD�t)�f�>y)"O��(4�x�hj�,g��9��"O����'x�0����\��ԣ"O��G]�5��rD��[��"O5E,�D6� kE�X�,�C�"O	``e��T�c㩙�]�x�J�"O�Ii'�ب%/^ݑA�B�(��E`6"Ol�h䬂�>Rn,y����`�UI"O\��II/0�a��֚#�ޙ!�"On+�AԤi�mWn�)��"O�ስ�ս�֨22��,A�q�T"O��(��P*hz��A�X.��"Od4��*Q�S>���X2*S����"O�aPF��)A8IaT,χ_�^�r"O��gC0���;e�6R����"O����hؽ֘�uJ�;`X��5"OX�� �vI`��iPu6�a6"OX�����z�豐�i��hn���U"Oj��V'�AИ�FnM9z�
M�p"O@�R�^�%���¬يQR��S"Op��T�D�W?�y֥ߧ]C� !�"O�Ԉ�ՋnD^�� ��bG� �"O=%�0P��ir䁑�oL�})�"O��R�A=�$��!U(��<�"O`�V��+Ts>���U/^���"OTY�R��Q���6Oå:r�Y�"O���ֹ��j���4|V����"Op�n�
y6�,[��NE�mhf"O���`0��iIp�J�p"O��Q���%lK����Y	xP�@"O���؎1*R[��P)dO4��"O�X��(T�.QP�+� ;����"O���`$ũu?�m���!K�IcV"O.�ZDoR9U.�: J�=}I08�"O,}i1̃�bY~h�%"	�!I>�"O"��tX�	�.��#씒i¸j�"O���g�&ԥ���KeT�B�"O���`�s	r1x�	\^T�"OHy�b`Z5x�ܸ����e\!�DBN;b8Ö?D�@���T'9g!�d��v�x�p�غ`�ѓ̛�WP!�d�F�M�b@��z�
�	/19!�D�D߼��w#Q�g!4��ߡ36!�$	�{��:4@�;j����J�!���U3���Ă,�(\��o�S !�Ă�0��l��K�"`Լ���Յ�!���W ��Kʩ܂1��X�!�$^�7:�	z2/����ӑ�N�!���!+�jE5�){�+%�%�*���9e 4�W��W����v�L�#�x���&<�20f��%���l�9���ȓ,�A�6a�L��F�cl���FIvm��C��,�-_��m�ȓRh6��3�C�( A�!)H���ȓ[>���B]8VY�F�RI��1�'�`��]�6O�b@�aTA��'閤�E�F'8��=�p�]H���J�'b,�a����{�LP:WN�AR�́�'��\¦a]�U� f 9� -K	��� �*��6t*��PKS�P���$"O�Qf�W��Hia���lc��p"O�8��5 	@�sQ#_X`�"O�8�2�K*V�����>LtEZu"O�)���9� ������E0���"O��z��5'-
�3�ef$�0в"OT!{�!|��!*ٿK����"O<l�P��29Qp\ٗNP4>����"OT��R� �De\�`1� L�x$��"O��Sl�> ��PR�,�R�Pi�!"OH��V�T�v����R	�~�2���"Of-0Λ"/<h(V&�5
g�=BG"OМ� /�8��`��Ǜqܡ"O�Tڇ�ϊ$���g�)U��0�E"Ot 3��������9+���F"OL8h��]<v�PE�ĭ��4pb�"O�3�	�	VL��`�	�$s�"O�H��X�F����` Y3$��X�"O@|(ǥ  r�A��������z�"OJ���2<\䐑��C�L�� �g"OҡK�@�hD����A�8�r"O:�{���M����c!�)nεJ�"OB���a�>y� Qp���8���s4"O����cT�7�(����?AJ���"OļyW��(�j�"A.j3 �H�"O̸���̬4�f���C�.�銶"O�� ����㣯ĶE��H�"O��2p'�m�<La��7X*2u"O���&�@�qPȚ�K��qNR��"O6�Ú� ފ8�3� A>d��"O0�Y(u�������t₇Ec!��D�H��)����|Ra�3C�!�D�[z���;�ҕ矦�!�$T%3>c%F���Ii�I�B�!��-U� 1z��Yw�ݹ�A8>!�䎍S�&�ӋM�qn��8!�ְK���,	m�`�QB�#(!��2%��jel��L��}bM

!���͢�dĆS�>��S�ȡN�!�D�P�j���?dbR�"UJ�:�!򄕯I�D]�� C�$�0�;4j���!�d�@^�;�U�<�e���E�!�D����@��٪�3�� n�!��jD�aAsB�:	�>��,�t�!�dC� ��a��N�*������{�!�[ K՜Iq`��4��� �g���!�$�_�IXwk*�:��$��=:�!�D��%��ɔb�(<=qTHT��!��C�8`E��D�/'�EJǇ�$!�ޅf���͈�"�N<��T��!�D�RhX�ƭ��9��ؤ���i�!�		��qR��ϔl��V��!��<�l8�r#č��Lz҆R�K�!��K>m�s�����ͩ�fH:2Y!�F!6E�%�/�8�j�v��/X!��C��*6�-N���(5�1nR!�/�D�%C
G}�]���D�H!�d
2����B�$�BQuR31!��L�)������M.~iz�V[($K!�DI�A��J�_/[f���\�^�!�D��W��d���E����C�@�
�'K�Z���a���Ç�D�k��'�>��ЪJ�qx��Ad�����'iJ�y# ��R2F�f3�l���x�<� ���B2�(tP7�	�>��(B"OBD�bL_lt�o3)9��9"O�t���^(�c��](>	3�"O�����a`���U���"Of�[����eE���)��%2�"O<�Q��v�z�uiK�b�%��"OT=x�A��6	�(R
���ړ"O�Q0�G�e����1%�%{����r"O�C����pqjH�g"��R����"O���g�<��<��� J��iR�"O�t����<N��9G�҄?6�ȋ�"O8������\��oö=�A�"O8��/�\�8�EN�+�v�"OTu�
   �