MPQ    ��    h�  h                                                                                 g�M=�ʛv�������`�Y g-x��c>oN�=�V�nv���LJ��
�qrQoEl	'�Nq	W��������2�)	0c"�#��������݇9@�h���O����D%(�>Es�����&��%]M�D����^��'���ɕ��"��l�z�Q��5XG���v79���D���.�i��~��e@�\;��rF��'.��L5�L�c7&&��fY��u�E�<tV~�:{\�=\O��+R^�z^1�8�qS{�o���8�\an��pIp�����H���fDD[��愈'$�D�|�5%��E1���Mx���Hv����r�]�
4���'�_�&s�R��_���9��n՝3�M9�<�H�G��K�^2$� 8VO�#&����1�h�T-��֑ˆ	�F5%R@մ]Sb��j6�>�{�D��w�*`Y�"�$�*�v�u62"�O +)(�(��6����`]k���⥖2-G��,�����QẈf�3�.�z2�e-���3���V��=���cG��\�r��$	��c�MA�h釨{�K��vd���H�S\�C���z	Xn�A>���uΆ����B���Cd���b%�?zv�s��c^�����ѫ���.o����p��r�OY%TLX���X�tA]N���Vꬨ����w��F �5���sܗ�^M�������<�V0:���R9����j����c���8��p� hH���J�6��n/�k(	��>&����ր��/�fa�Ob��s�\p`�� � 6�w�i�~��	��̓���*I�lC3_��j;�����]�H:�l ( ?"氘Ցփq�����Q��G9����X9��K��'�aV��4F0��������A&1�]y7�=�ꔶ	��zDq�P7� C�S�b.�M �&���R�V���!5Io|�X�֣"�n��O0�ã8;�i�i�p{�$� dJ�M�P�yU��5I�Ăt �t��ڱ	�ڥr86��i�:��f�����Y'��M����i!�ђ0hҮ�F�ͻ�-�{-�i��s����Q�	'<�a��K��^'�,��ע�\}�������[�j���䖬D|$�_�=��.���j]*����d~��/�s���J(�fG�S*=鯑~����}/��Y���ʷ��@�Kt$e�rL�����*t�k'� s���۱��w������7B5m;^�0��[�^�h��w�׸0zM+/�ч1V)a)��1��D��n��r�Z��b��L���JD�zbrR�xL��t�s$�i�yc��K~7X`�aZ%y��ө֠?�r�6c���n$U�^s<'�_�10.�ul������Fp}uy`4����7$�]"D��:m��|Ρ�o��KP��� �MXͺ�0n^2}ݥ�
�6��z �������m�rh܊B�P�h7��}w�"D�����LLQ�ޤm��7�R��KϠp�T,G��#��r�J0WP�ⴐ
�� �e�Y:��hL!��r��~tK@��(�m�A
�)[��kt�E��/�d)��E�6�����[�<�zh,�#������vJ��.�֓�I�Do��`G1��*@�Dc��UV�A�ۋ�� ��[R��'LX`R�}�:��Df��s�5�+ ��爚���"E� ���ȸ� ��̛m3l�	�/F����J[.����Wc��#��N���0��2�/$1qh�C�������z��g���h�����u�����O7�*ʸ$��`U��,�:E�[e����m�nF����wȓ��;�8���1frqM�XK��i~��b�q�շ�\V��Z���r�b��g�Qo�|X��M�� zhEt�j���!�f�a�6�_��F�3��r堕z1֑op��>E� |�*���� V ���*.�/��4��$2��MJ�X@�y#���>[�0	��Yh�;)@2�B4We��F�?>�����ݶ(�x�թ�u��GP� �(T�&Ŭ�W�.�ah-�}��Z���
#u ")sid�W�3c���@:_�'�r�P@�.ri%�x�H��a��EM�P������8s���,�׺��0P/��9�'�U�I �,��b�j�cI�<�!/,^��FZw)��Q�#ݫ�[-����A=PB���%��f�zp(�v��Y��'����x@�\����J�a��j-m'�������oҦs�;�b�$��B��2f�e�����(T����}\-)	�E(�����>�G� ��st���%ܞ��E܍��4�D��n���,ed�-蔎�Ғ����W��s����廾8�
]Yȗ0��5�}���U������ ���~ŚM��K�'�F�v�R������[���K�h��lK�ajR� �D$sĎXQ�NsQ�B w�[<�q�GxJPzS�-����&�l�V�4��p"ذHV#F��'��N���A��ѦfΟ����#���D�VB�*�Z��{�D�p��+ak��}�b�xS�Pg�R^�](��W|�5C�.�U���_�������W7��&��Id���8@a>
�q9]6��'�� ��2EHt��g8��Cb$ �q�	P=��(�TW*ˑ���y0zT���q�k�6�`���7�8/O;N����<ڔa�WN��I��e������j
m��L�P?��'��j�ٰ(/�U ��F�8���S�QN�`�D��d��v�r�8s�����o�x��t�]�l�h��&%!��=�}v̎>+���ߕ�$��:B�o�^B�� )��� l�b�i��?|)tW�8�NK�`�>NxS`'<�I�ߖ�P�9�N��D�Q���6V���j�,�sH���C�Z���k���Y~�M�@Ω<�*�[�*��:?{ex/��A��~B�d�&�E�蹤[�D��B�d�gĎ���W�I���d�z���|`��z	�`��ֺ�I^��k0P�aM���ް4u9�ou���j=S����H��l�fp��!s���%3{摒� ^�J�I�T�[v�<N�C����f=TUJ�R�@Bjh�Ĭ/ԟ�){��[�3ڳ�F̸`��b26{w�^���>�nְ����Z� �xg>[�6��6t��̥�Nb܁*�=����,Rr"*1h�B�ǁ�s4w�ߗS����r2�``,?8_:���� ��[蘓����4�GNp�����*�?���LPo���8&���Y��ua�_W�@�
����\=ROf�n+MCz�*�8�-zn7��к���a��p���Ù!��+�HqT��~B�_bw$�Y�|_����14�M3�z�c��x���8)�4�'��!�3R[��g_�Ҷ���<ם�9�gH�p���1�^��� 󦤓>��-y׾�����I�T��-֌|b	�%a�x�i�(!(��fH���S���S*_[���r,�?(����ucd]�� ��ɞ#A�6<�5�|Rgk�&Ǎ.�	>�Yֈ,9�ݮ�����?���Fm��ğ�����$��ר�������D��f��#~�F�M��S��֚v__����C��&��6�np��2�����68�$��܍d��.b�C�zQ˼:禯y�X���j�$,��Y\�p1A�rd%/��0�"��XN�$��Ԩ�����we*�F���&��2\�^H�}�;`�ʊ�<��]:h5�R<��XjǇR��c�����,�p�j�H�*J9���IK����w�@�W&�(ܾx���J[��͉Oݠ�N��\������6��iZS����#�82*�҂l~�V_33;���
]aH�� CB&"a6h�lDq$���y)5�Bd�G�X�Zu�f��']2��Ȇ04�ˌL�f�*�A���]�y��X�1����m�D���7Ν��Nb�U
 O����U����S��W�I�m�X�+�֞Nn|�0��Q�S)\��v��K\�_��d�N�K�����5��ĝM���ڌ����p'b��+�:�H����t�%��]����!8�"0td��|F��J`�#{H�u�t ����DDK<�&��,�����N��q��ZE�o+���ְ�߹�����~h�����]�I�͗T�W�n������!�9SE�B�y�~i�c�2�a/�Ӗ����%������t?��r�s��ZF��e�!�s.�����5�W��q݀��łPA�5Ht��k B�6k^�[����s(+J���f�VE��(�����n����l�Z�D�L�ЕJ���bM�E���{���s{����ŀ�X{��Z�cg��(�<��6^���������Wb_Tg�.�Zl&[cĘ	Fk��y�:�G	s$;�"�Fj:Hx�|	-o װKK�{�X�k086�2������Ձ���v1N�����h��O�k�7�R|�D,�i�YQ�G(�Q:8my�6�m����0lK�,Tg�:G9�f#�7r*�0��=F
X���@�QYu��h���mh`~�ϧ@yu��-_�<�B�:.St"O��*��)q͇E��x��}q���*�U��,��zZ����gJ��@�����W�������s13u�@`$��\`V�5�c�拭R��{�p��Co�Og�L�H����`����_�����9�h�;n���>���1�"�z�=zV��`�/;�m�Y	����,��~U.��?�T֮cک^�C+��q�m�$���
Bp�F�M�>8���H��u���Qܰ��ϳ�j�J��f3���K��{!X����E��j����i�;nAh?�f�N��;�ŗPvfM[%��pZ����~����͐�\q]*Z6��r��0�.�ɧ�у����5�����h`j'���U��	���EsF�e�:(V�P۔LNo�:�> �R|�p0ԕ�xV
��<��ꕸ4\�2f�EJ��0��t�-�[��%�e�h;��@MS�B�h��~��z��������W�i^�xZ��˥G�`V��T�������.#aÎu}L����
��"
xdB��Wv�&3^�����@�v"B��?C��	��i`X�x4m��\�펠�PlDZ���w�Yj�ݘ�,5`w���*|�9R
�U�w�Gw����>�t<ش�/�X�ʔxZ�6p�� �>�R�� "��$7AN�P�MS� �Ff߲W(��Ǜ2������z�{�\��-�E�`�F-(������%��ҁ�vH `�=��2�w0����C�&�v9}}7q�D�(�,ۦ�i�>&R ��s�[Ϛ$�����ȃ_4�V��i�N�I������Zw�u[��#��Ip߀uN��H
�h��R+Y�P︢�PU�16�A�� G�J~�u(u�q��!K�du��&v�#��莕b�.=w�#Vlf��j�����7��N���0��=q�ⶡ8�,��xec�z�{�-��K�G���DV�pX��ݠ�C6#a���[@N��0�|���d�fɦ��݈����D+�yB-7<Zzv���%�Z*�kɘպ��mx��P���R��U8o�Uy�Ь�.���*��=����}�W�[u&��d��J���>[}q����?z���A��2���t=ɏg��]C]W��K�P�p�(��*F�6���yk���s\l�t��ZA`X��Rq�/ʾK�֠�<PgF���MI�|IS��eٵ���y��_
H��Ln�?T7��Dj��&(�4� �+�R��Q�V8`z0(�_�v ��8�|_��$�����g���l-�]�P�!lN={̩jZ�|k1�4�$�w9�z=���B6H ���8'��䇍��Y)�܁8[{��[�{Nw7(Ҩ�d�������C��Df�������R%(���5����ĺ5L���~4�m\��H�)�"��O�E�Ȳ�WeSz���D엎_ &��=�t�g[�;�A*��?{��Ɏ��"�D��ѿ�]�֎|{rjz�mB��w�Ԅ��tˣ�1�W 9���戊�����=.��v�4fk-J�|4���o�3�s��y	S^rA��WK����v��~���$Ő޴Tp�5R�vjCO��j�f��Y{��ʎ�U�ϝ`��b}�LȻ�P�+�-��>Q��۰�@�E;��g�C�6��{t��}�@�tN�����R��,m�*��tB�jB�Xq	wP�S|r���ʋ`Ў8,-�:m~���T�����.��$=��p����0�?qH�;L��8��N�&��fYt�u��r�UL�qb�\N\O�|+H�zD58=rg��e0��Ega�&Gp7�>��Ap~H,$ƻ��_Q)M�:\�$1�L|���Z�1k�M�3��~������U4L<�'�΅�6Rc��gM��S�d}���2*9:�gHH#C��71^莒 �^�Y��������ޟ�Tc��ևM:	jY%�q��y���%ʾER���z܋����*�v�����Z���l�Qu�f�T4 a���6�[�7d5k�������ԔM/,�YS�@8�pK��ܵ��zV�[|��qa��_;�C�;��ۨ`���_��B{�|H]M�`����>���vZ'�Nl"�ɡ�C���p�FnK��R0	M�i�����Փd�u�bܜz,�r�u�C�≋�G��IK�%>pL!=r��Z%
Ҏ�k6`ЪLN�MW�[{�ch`�}Bw�X�F�}���R��<�^C����ӯ��i�<��:㮱R��!��.؇�	�c�j���]p^ԠHѹ�J��&�$�ϙᦺ�ۋ�&���i@�P��Y�OX�H)�C\��E�V�>6��i�G+�a�7�����*�|el���_ο;;�ܪ�e|�H��� ^��"����G`4q_���!��=�ۖ�0�X��ˁ�'�"�����4�d��7��A��P]��g�s�?���D�� 7����5�b��F 
^���x��C��r��I�~XUd�֙�3nyG�0a⃣n7��_Hs�&]���vd����F����5��ĸFf�jɸ�gP	�5����:k�
�kh�Џ���Cm)��,!s�0��n��L�FXF���{ci	��-�������<!��u�A���/��, �RX��J���Z���%y��������kר4@����`]�KT����TW�i��?�y��,S`=���~D�I�m��E�Ʀwɀ�A嶻itZ;�rBR׊5��̠&���N������G ��b"��j�5#��Ѧ��G2s^�&c�-\����+eK��'�NV�H�c��zv�n��F��,����6L��J:O�b(�h��@���gQs�u�/�
����X���ZnKn:��L�L���6Y~4�$���x�Lr+�_ϼ�.�_1la���3� Ff��y	��O�$8!":��:#(I|D��o��KFD����XC<�0S�2s�]��+��Ɓ����<�#2AhR"�ۆu�7I -�Dgsh��9�B$RQm�km4����U��A�c&TT��G�!�#z�r�w�0�'�C
�u:�9^Y�h�~��h�J~*��@4r��7���HMu�t�x��%<�)��AEn&r�����QH��0��,��������J<	s_�]���S�:�E�~��1nm�@�#y��N'V9�K;6�ȧ������K��j�L��ss3޶�ǉ�zƧ�iA*�CȬv|�������"�"���-h��F����*m�Y	4(q|7{���k.P ��c��������]"�̨�$g���a,١����6��Iۂ�5Κ^@����0�N�$�E���\���s��"�"l�E\�_�HV�Qn<oV�	��;*�ۗ�
Gf(e�εC�G��~��g��Km�\�GZ���r����i�է��g���^ҐN"�D��h{��j�)��f���d�ȕ�F��sޕ�&�\�g�`of�t>���|���0�V�d��ҥ��
4!�C2�nIJ������_Ȭ1[�h^�g�h�H�@h�oB*���Y�鑵�.���g�Ĵx�E�$�GF�֎�T2�!�.e�a-}7�� r
�?"��vd}��W��3Y�y�F��@���]�l�U����i���xϱ?�W������P'���.��,ph�p�%�9��Uq�<�b|��X����D<hQ/bsS��Z-d�r��Y���Q�w�BA���Px����f:�(A�M�2���ƣ�l�H�\���@�{D��-����M��w��\��������8Vk2&��;���^���c}ՙ��()�#��,>��� c�;s����D������n)4$���d8<��M�]-���ᣒ�ũ����V>2�O��x(
��F9�ka���:�U����|�� �~�p���،�\K�ʧ'v�D�YP5u���ǔ�����6Rl�~jH7˂�yl�eu����8��R���?�x��KzI8-`dɂ�آ�:V���&�	����#|��=�N������D�Mf�͔�8��h�lDF��B�cZU2O��(���HikĊ���x�'P��DR-X�2�����k6.{��ƅ�!������\W-�&���d,��n	�> �q�K����(��2���tx!�gnY�CX�Ē'�>P�n�(�*�"~�̓y� ��<>�g�Y��7�`:��m�/Eb5����<��&���;D�1I��:e�Ƀ����M�
#WpL>��?��f��8j> =(��j ����m���Q��k`<��Zj�v[�8�����e����*\l�55U!u��=6Ǔ�Ķ���:���3$,x\���B]� ���#oj�X�1�[�F)�8�Ǒ�VrTN�֜9�@Bߌs�����~W�D����l/�C��}+��B��wC����9����C���hؠ0�`�q�0e.�����y�Za&Q�$�/\;[�{��p�����`�B��?�6��푅|�@�z��O��8�Կ�Jǡ�~���P��S��XX��ǝ�h�=	s��M������ff����w��|�3���0^MX=��r��v��*���^�Kv0T�H$R�7jR����B��{��u��(���`�b��)�40���-�ȯ�>zT��f=����7V^�g4L�6��t(����V�N���d���,���*'��B�-s���Rw�ySw��(��`֓b8Gh�:�V�����@���ck��a����pm@��Wb?|Z�˲LƷ4�4
&��@Yϕ5u�r��ֲ�S�L&�\���O��+C�<zo}�8��8�����ɴ�aqbpҝ��ӆ��mH����������vG$l�|������I1�2\M���ܙ���n���C4��/'U6�$�R���"S�D���?�Ģ9uH�����]�^Ct� i�{�t���#�t�h���qT�2�ւ>	��%�3������/ʙh�*�����J�*�S�S�S�u��>�u�$��4 ���/ 6�k@���k9]�ǃ'r�� ����,o� ������<�d�ό�Χ��S+�L(���N�ޙ�����t��V[�� ��j�M�Ҭ�8P>�`�vU#�S�Єt#Cg���?n&8#����Sˆ�|���t�Nx�d���b��}z�j��M4��������چI��pg!�r�=%�D����E�7N����gâ��t�h�w[��F����S���h=�^>����f��@h_<y1:^H�Rʭm�����uc�I��I��p^cH�z	J/����ؙ�Ѩvb�&�\��.Sŀ�d���O��B�\!�,6�v�i\Ņ:hR1M.}*�FXl���_il;�����Hk�� y&�"W��"�Tq��怯8��8����IXj��˜|�'S3��~�r4�!Q������ A7�]<ە�K6�i�h��D"��7R�;�֣b?� �)�����鴭M#'I �X�=֔n�2�09Z��ev��9:�~f��d~��A�`f�S5F����_u����BFXP�Cd���:���&��Ъ�-Ҿ�a���u!�h09����F��iִ{~X%�j�Ǧ�����<����Y�eX��� ۚ�uŲ%����Y��;����_#UctАy��O��Z]�î�C^~�//�d̞�������S{��b~ɟ���"e����*�۠S�q߾tu�r�P����ۯZ�<����^3��E������覂F��5�E���(���M�^ص���ʷ�a�*+��X��ogV�l:������n�K;�"�y����L�h�J�.�b_{�)�`�EYSs��PO�|�X�_Z���I���`q�Cz�6Tn[���3���]�_J2y.]��l����Έ�FaN;yq#z����$7UQ"��:���|�oV�KA�q�1�X�,0n&�2�囦d�5��L�؍��~�hh��ۡh�7�����D�T���B�=@"Q�P?m� ��3��S�%�T�p�Go��#ufwr�=I0���3��
Nb9���:Y�v�h]|�c��~��@��u4�P�޺o���tX��� �/)'��E)�o��N��ʫ�~_,C���\���J�P����KU�wx�Yw\1���@�C��a�V��0��ɋ���qܘ�us��ōQL)���Q��{*kq��&x������B��	m��c"V����ԑ��%x�mą�	oa��ᖓF�.�r���sIc�L�9��8K#��]$t� �$�������9�k\�zs�9�&G9��47�@�����U7��T���PE7xE�<����Dn7�lʒE�ėq;E�y�	�f��	A��՞~�=�s0��'\�Z,�r\���X�"v���]|�����h�{�j���!��U�0��F��]���W�������o�/>��|7]k��]V ö��+d�`��4<��2\uYJ�z*w�ce�[�4�����h��c@�OB��a�4it�������� �+[x�::�ƝVG�y!��5Tm�v����.�ay��}�Rلw
���"��ed�:�W���3Ty����@kx-�5��Ϳ�{iֲ�xj��R�-�V�P����/`�4]���,�Ќ��?a �9/4U,3��}����|���pd<N;l/������Z��l-���t�X���R
�A�wvPy*�Gf���(���h����Z�~���1\��?�;���<�-��{�*pߺ!W�7�u��V7��3E2w���.N�ygN�l�}�X
��L(��Ħ��>��[ �Os�g$ϐ���q���>x�4���_���=r2�w�߈X�kP󪂷��S߶�绯��
n���Ȁ=���'��U�w�Q }�l~���+\��G��K*?觐G�vlB���;��	������g�ݙ��l���jâ���T�?���>�3���l"����x��z���-;�bɽT��=��V�H��y��#��>�No{��h���f������#��Da��B#� Z0q�����qk����s=�x���P��0R|���\t�����.v�E��t1�����\�W� �&z�dX���	�>��FqJ�썵�.��12�{�t���g	�^CS1���9Pn��(�s�*<��ݨ�y�҈�(b��G5�`���ӈ��/�%���T<�c{�26"?��I	�eO�������[_
�4�Ly��?��*��tj�s�(`�� 
8���k�
Q�~S`�g��U	?v��Z8?�%���E�֧
�<	lc�d�x!ОM=����"��r*��pҾ$G�^A�CdB��� ZA��>�5��9h�6}D)%G�8�4�Qr�N-2��������"��'D�x��76��<�����o��,��������W�>G�I�[1��{���1�e	pS��z'+�U�&�f����[/�ķ7�Y���y�?Q<�� �:ڔ�u*�L��|�.�zz���n�����<[j�����.�e��������d�=��vو�M�j��fa���2�L� 3���ox=^(�ќ���%skv��S�T ��.�T���R
��j��0���ȟ�½{�Am�D���w4�`�bsj���Ա�d�c��>uw����{��cmq��g�t�6c�tc+B�v��N
�y�;V���@�,�b�*�b-B����w���Srħ��[�`�w�8b�C:c�5�PƉ���d�]���X�p(�V��?�c,��L����&~KWY*�u�l��XB��'
r\��,O7\�+>�z��)8�[��+�[O�ŤC2aZ�qpmO���e��X]H�#��Ҡ�G����$�YG|0�l����1!��MdI?ܴ~�� G��wa4�
'�"�qR���xe�#�N�Z^���2G9��$H~���^�y� $Y����}�{%�C���T��T���}O�	 H}%>o��_���F�t�@�����M���&�*p��g]���D�b�Ru��{�� �7 �֐6M�����kT���ӣ��\�
��,
wF�	��&�D�v͌�Ba�QK�'��՟�y�;��5���r�H�[���r�CM�d��sR���zvP_[|�?g�C!X��f�nuz���R�3冝O�5L��	�d��bm*z�h���0y�JWt��c��5䧘�.p�A+r�%�ׅ���7��WN����KJ��o�s�w��Fl�=�����^^9���L����<8o�:�OR��i�	�#�c�He��g�p��H\eJ����ڦ��W���Y6&�&���\*�{����ѷON/��!�\\	´��=6�iik�_���Hm�E���*p0[l/�:_9m;�|�`H&*� ���"҆���i�q��I�Jph�3% �X%?X%|�˷	"'�cZ�Y�42]��]���A�F(]�;(����6C�MD]B�7�~��Hb��@ ���(���w�(�BI[�X�5�֏��n/>�0ׯԣ��?�UK-�ܾ�F�d�a��<D&���5�5����`b��P���޲��1�:!r/��a������9��[,�!�ڋ0�@���F?��̚{�g���}�gC���[T<W4��j�����U��; >�H��� v����@��$2���m�E�K���j��y�]�[Y�~�{%*߆_N��K�Rj=S����}��~�f��6� m�����6���,#�t���r8o=��%�YU�ׄ՛�B}�F�
��}��S��?5�������}�+^�d&��X-�!R+�Mk�$�V��5��nu찣]n�ŋ�}ٽN� L���J0.~b�M~�d����j�s�q��4��7}�X�}nZ�$N���5�����6O~�ڡ(���\_���.8�lכ��ipF\)�y�]z�x:�$R�I"0�:���|���o�nNK<p���fX�=�0�N2i���vAT�p�ӐG
+����2h�9�ۼ{l7u���:D�U"�*k�8|Q#�m����1g�7���T}�G
)�#pmqr;$�0CW�N�
�n���P�Y&��h�[��^~4~��@��L��I�-�ޕ�u�4�t�+��V)�"�E�q�3[��Gm>��oF,~�+1&��y�J�7�a�����0eW�41�2@1�o���V�V�֡������߶P��� �L�J<�O?�8�&y����0�_(�������9�SN��,	"���n����P��F�m�#	���`����.�����c+L ��� ���� $�_s���X�W�M�o��5�%��d�;�a�τ���;��w��ސ�E��0E�wu�:��n2�=%'5��S;`����ߌf���D�R�}�~��z��ů����\�yZ�'#r7v´�芧�����U�F����h�h�j�*f�� �M{����F�R$�K頁���v�o\m�>�!�|r7�f�QV���Mlv�;4WE�2כuJbpc�e(K�=�[� $�G�hlֿ@���B ]�
��+o��d]Z��/�z�`x�����6G<6y��T����WR�.I�a�r<}}����
�"��Dd�PWG�&3O`��re@&~�������͚9ei�x�Z�M�7���fP���.�P$�X�nX,��P/��69cq�U��i���Ne���h�<�.�/��>�Z�{�h��ݷ�G;-�-��A�u�P�>���[f�(�EK����٠�Y�,;K\Q���6����-Y"��Ev����Q���'%v���.T2����ȔX���}��J���(_སݗ>7� �?Hs�C%��ĞLMF�y��4ZK�Zb�阶�ӬZ��O����Ȫ]�"�̈��Q���8%
�V�ȃ�e���[��JUk�_���N ~�������s�KE�ͧ��vG�v�φ�k�]�����?-:�T�vl�;j>.&��O&�z�i��)}�.���/�]�x�\8z?��-�F�����}�V�����ϻ�4w�#�fs`�NJk��-�?��if�{����ޜZD|A�B��Z
c�0�=�+��k���ή�x?4�P��R�{�����]����.q�U�;A�n���&{NW#&Up�d�&r��R�>�R�q���p2�I��^I2nx�t�1g�x�CN�Y���tP)ʖ(�h�*�3q݃�lyG��r3(]M���R�`�R ӣ��/;	��g9S<D�ͫ :яId_e
Q6�{��u�
�2*L�9�?%y���j��I(q %�X^�F7�Q:C�`K���P��v,�8�Y/�(��[
�ւ^!w��l����!+h�=��A���X��9��K�9$����w�^B� �v�Y=��N�*�'R)`,�8,�8�L��N�5gL�ǃ��߂�b��w����D7pQ��"�����V�:�߼p�m����W��>$��9�V:��RW���{�&mse����p�h�PC&t襓n[J��]φ���zb-x�5&�������|�<�z���I�5��������D�h�ɰ ���ۙ���f=����%x��af\s(��8q��3�%����^�U�R����`v�0���L���4T�ƙR�J\j���;��x�t{�� ʟ���2�%`(�b�g��n��f���.�>p��bA�qQ����g*�n6>k+t�~"���Nڻ��#����,��c*�kBg%�	,Aw!�;Sm����S�`L{�8}>�:޹!��-�G���dh�����p�=l�8�?r���D�L<�I�j�&y��Y��uM�o�XE�z�\�ysO�·+9@�z%Pt8n ��g�����a�eup!��t�R�LH]Sf�������	X$���|�${��iY1|�[M��ϐ��dV*�|�4��'�e:�Rt������>�!���؝z��9�T�H����	:^��� �)㓪n�g¾S���bT4O�x��	{��%�ʹ��2ز;h�O���b�K6���"�*ˈp��M��`���!u}f�IYR 2����]6��K�hY8ko��y�!�y�:�Es,�5Į���_,��r��ׂ��bg��������̒�*���F`� `����M���
z�Ri�vK?7_�Y��yC<�G��,7n�����3���B�����ē_d&7b�e�z�pJ�&4���-��!�ڐaf�E?�p��~ra�%������{-�N��f��q��#*�CwQ��FG7h����ܞ�L^4Z���r����<S��:T��R���D;C���c�gl��e�p��4H"]	J%����ZY���{��o�&�Ӿ�o�6�����Oɞ{���\�C�'�6���i������-���$\(*K:nlj/�_�%j;����v�JH�' ��T"M�_��&q�����.p����tX�q��Ҷk'I���4F�4m�'��Y���A��]����[�����D���7�Ĺ�x�b��� ;!:�C���|�F�o�I�r�X&�֊>jn�i�0�F�!1��|Lη�K�ndQe��7�'+�5��p�	�k���s��*�>�y!��s�:|���Z��;�Ҵc�6��!$m�0o_���Fi�L {����`���B�v�0��<�x���B��R���A�VI����ۂ�����q�"�˅tH��������]qT�����Dg�Z��P�D�C\S�������~�n������l���ɑ1����t�l�r����ƽ�Q"�ru=��F��,1�xl��2U(�<��5���W�����^�3��>c�ך=+��Ň��|Vp�N��Kj�n�_8��X�	�;L��J�M�b�\q����{��sO��@9ـ��X�Z�M@���*��y��6J�}�5�m�����!�_@}..�l���x8FW$�y'���3�$m�	"���:��<|��Uo���K76����Xtn�0���2�\�Q�����*���dΏ��4�7h����׮A7�n�S)Dwݜų�3�Q~��me����O����R�&�TS��G��#k��r�*0�(�i��
D���dYa��hSzZ�Yp3~;��@e(г�=����p�&w�t����y)�~pE�}w�N:L��/]���=,�eg�%)��EJM?��ԛ�5�P�r��1�@��~����VJ?�OԽ�gM�gm�+#�;4L_��moD2�l��FѪ�˃�Ԡ7'g���T'��	"��)	��
���5\mz�	�3�M�����W.a���@�tcF�ۿ/.K�����YF�$8k��}�ٲE��*��P7��b���)ܜE��d�6i��Ҙ-��^j���z|E���Ჶ��Օ.n-����$�:�9;{�M���f�B&�Ex�O�~�ݞ�)�O�|m;\�%�Z"��r����3�X�{����ҡC�um.h�u6j�~hF/��6�f�F���ަ=ڠ<���n�o�hi>��{|��v�Y�V�$O����ք4r(/2R�J=�������6S[�,��xһh'Ϳ@���B�����ʙ�fKʠ��������w&xFo���'G�gr�T�j��� �.�a/T�}8���
���"p�d.�W��3J��WJ@�$�+�+M��u�^iL�5x�?��H�ݎ"�PX��I��� �I��,!�r��>�&9���U�nf�K��m�����<�A�/3�;��Z>���ߨ�-��^�pA:��PI$��Y�fK��(r	*��@@��w?�4rgd\�J��1TuU��-q��`�{��x���bY���}�)�&2-���l��ȯi��bK�}��[0��(��ؑy>�&� ��$s�?�φbM�'��ܴ�?4��w�U'���g��A�7Z�a�*�8˽�����ụ�
$��>V���w7�
�UF�x�-Q� �o~�!��Gؽx�K`�{����v"��
������U������lҳuj�ٵ��j�ĵg��Ug��)u8�"#,�3:x��z���-�U��37��s&hV����7�� #�����N%܅�h���ff���Ibt����D���B�5Z�%%�k�C��d�k� κ)@wx���P�iARrS���ǡAB��<��.l��Ɩ�P�),��A�>W�%&0�d����?��>�:�q �\�+�d����2I�t)�g?8@CIc>�8��P�'t(~3*2��^{�yW
v�^X�1����`k;�Ӿ��/�{�B��<<���hA�59I�i1e��U�8f�����
�P_L��?�y���@jOz@(�o� @�A���! HQu'?`�	�K��vl��8����Ccn��1�]�T��xl�Y��8�!�Q�=g�n�[(�hi��&�$���I�%��Bn�[ �`^�t�d��y���o)�1e8�m�G҇N�t��ă�f1��cU�����/(ND҇M��-x�T�R?���)���ĺ����+�٦v�4�B�T|�ђ���Fݲ���e�������➎K�&b���`_�[eTo�-Q���Vĵ��d?�0���+�,��)�|�j�zps��$;��pK��r���3�ù$�۝E���3���#=�vp��lv�)fWu���y���b3�ȏeg�^�\ʜC���[��v���
��|��Tܵ R �j��V�{���{�Q0������`C�8bi��};��<�l����>k��w$G�,_��M&g�%�6�t��V̬�oN ځ��>R�,٢�*���BB6��D��w���Sh���9l`��8��:Y��g�%��|֘���tw�_�p��%�S��?���\��Lwb���&tI8Y��u����z8�]�1N\:�OmI&+4��z��8)����Q��Z��a�mp��� ���<H�N��=�榃�$��|f�!��Y�1נM��v���7��˹��-48}['&-���RϞ S$��Y��P�םU��9& 2H�-[�֏J^T�� �-��v��rK��͞��8Tϫ��s�r	��%�Fڴ�%�����*�>n���>c��>�*&$��T]��>B�X�uX7Q�Eo ��<�
�f6_q�#�k�X����T4BԀj,@���GV��P����u���G�'��<U�K�vׯ����=���h�;���h�ZMc������^vF����Vе��CWL��\�4n�N��>�l�RA��U��e�Q�dA��b~�z��2�aW���L���������� ��p��r��o%v]=�W/��#�N�1��x��O��,��w�R�F"�"��9��^/�בឭq$r<n��:�ԜR[�q�$�Yx�c����Z��pJ�CH=~�J����.ҙ�#�G��&�w�?ϔ��b��ʉOD.����\ҝ�±6ӕ,i!Y��k�����6P*&d�l��7_:2�;��܊�9UH�� �l�"ȱ�ճ��qK����?#�)����X�����}'�$%�Ʈ4�3�Sr�+AH�]m]y����v;V�XD�.�7#��y�bP�: �L�^E����!��D*I�jX���օ

n崅0M���گJ�KΗΒ�v�^�d숚�2Rew��5w�o�$kS�V{J��?�	���g��T:ה��W�����F�/K����!_A0
J��@Fķ\�{�����ݦ'{�k�i<��ھ�:�񭡌���qT��>����\�FRl�����H7fj��b<���oT�]L���ws[ǆUA�:���;�S̽��s�
~��B�Y�*6����J,�쩊�
�t�g�r.Ԋ��̌�����je�����3{{�M;%��PF5�p�ђ���`�^�"����X��4�+��h��yVK���OM���Pn~A�3R9�ĻZL#=�J&�b��T�ک_��)s�^]���sX�%Z�T��ĩ8@X�PE6E�xΐ Ӑdް޳�_�R�.lM��ğ�FR?�y�2;�$�l�"&�i:�'�|0�wo'tEK2�B�3X/�20���2_���,׃�����}��@�����h>�O��7kc��٧DS�,�`�.T;Q��zm a����-���W�T���G@��#f�r�P:0���
������Y��h�M�T��~�&�@ �7�R#�"�K�^aټt)_���W)8�*EZ���i9��=ꜳD,��Ta:����BJ��|Kg��P�J�&���"1Z�o@gbF��Z�V�b
��4<����϶���v�pL������{������Z�U�$¯��b��������"g���<ظ%3��C�mU��	 ���y���b�.����O caX߿����Ʌ�̔�Q$Ӗɦ�v����hބk���u,��O����JϺ�~�1�H�-BH��3ڐ�Z�j4Eȴ���pd�p��n(1Tۯ��V$;�>��z4f��N��
����-~��^����7X�\�gKZ�Br��Ui���^=��7ΐ0�h�5j��cC&���j�S�F�^E��+���ӆ�oR��>g�|�*Ԝ�V񅕉M��|4�+�2�H�J�U���4O9[�XZ��}�h��c@ԹB���ū4��G���D���A�0N�x����|G2B��Tr����.���a�U�}�)N*q�
B�"K��di�W}G3EZ_���/@�ͮ����ߗ�P�hi��{x;��C7 �gyaPR
�d�)mT�$�,\�3��n���9VU]<����s�D�w����<�t�/�9��SZ�Y�^8M�ŝ.�=|��R�Au��P�)2�f��](-팛����	6�� ��_\����,� ���-���{ⅺ��������8'j#�$҇2�g�'���ʚ��ݟ�}~�<kW�(�M��ӫK>�� O)�s\_�B�Kg��V�4��_�P��N�I�,�0>��ܯ�i�BS߇�B��x�
�����"��i���P�U!j��h�� N�~���<���x�K{v�iv���E}����|������9,l�{�j4�1�f�����.����$�S�}S���n]x�Ez5�s-�;��n�|���V�|$�f�4#肦	nN m���
�&�f������ĵT YD�3bB�U2Z�a���E�a�k����)x���P	�eR�J��١|�ל�.g����`����\�Wh�&t�d	����J>�Bq[�č��P�T�X~2$҃td�wg�ECD6ߒ��P���(.��*�Ĕ�9cy��E����Si��X�`&D��ѣ/10�?�<w�1���0��I�e�X��Sq	�kG�
��$L*0?[���j�-�(��F [�Ru�#���nQ�+C`����F��v�ț8p���^D5Q���8fX���l4P�{!�Z�="��0'`����/ $���"L��B��� � J؏���D�S��ڝ)�VP8b:@�B2�N>�1���|�xI��[�b�jX<Dm���X���{��Z����cEB�|K���f��tI��/�
�	C،�-�̾&�Dxe��UK�̎F��&����K�[��з��ކ�(������܂�+Xц�0�}�E|��z�?��{jԫ�3��}��)��?���ǈ����-=ub��9�H�;dHfR���C���}��3�ӏ�H^��.�~���?�v�굩eEH�7HT��/R{�j�X.��s��Ъ{�	��UFb���4`^�b��UX(�wV?�4.>f�~����猧�2ng �+6�z�t���G�
N�UԁL4��
�,�ru*}�By��H wWa�Sc������`���8��q:���B����%\�5���X�i��pY���n/�?h@�7VZL��.��8B&o�Y;7u��Z��e��ut\u�|O��+/�zۢ�8�g@�����5��a�Xp>$Y�W��,H�;�#vr�]���$XyV|�_��i�12��M��H�I�Za��Z��4s]�'���LR*�����tE �˟��0��9a7HO����57^�IX U+ۓ�������h��/pTji��nB7	1��%o�~�9@�
��c,yo2��gU��z�*���?{S��<��ӄu3(��Q@ h�/���6^EW�ޜ�k�A��o��/�Ի��,�Ȯ�D�7b��P��7_����S���䆦�J���¬��M��y�u�V�f��4�M>ړ�$E���vA�1t�p�sCr�ȟ���n�렬y	HT�����o�F�5�:/�d\�b���zs�j���@��(���>�F����p�a�r�G%QPA��}bб8�N���ӤA�
��GU�wG!F�Rm�?^���^*&q�]�j�,��<��:J�R6~��㹇�c�c�/����p�HX�)JV��k"��v���-&�Dw��8����Z�#��O��dp��\#�]s�6ΊHi|�.�&���`1*��l��_�^,;�\��,�HW� �n\"C�cՎ�q�����$f9�i��XV�*�qW'?�<��e�4��N��czN=A�&�](8��� ����ND�(7���b��� ����y��r���:�I��X\_0ր��n@ �0���]���?�mA���d����-	��7�52U3�?���7mڮ�ND���^��W':2V���k�$ҪR}���!��0�-����F����6{�T��V���ȏ䦓<(b���R���D����W��+ײ����:P秓,��+���`�|����Y8��<�]'�9�/km����PĄ�W��T�S��e���~��Y����]
�����GB��]�<tႷr��1�|9�������U�ݮ�W�^��hAJ�25jid�͹��N��^�1����M�`+��S���V&<��l��Wny󥡎k9� ^L>J���bo�'�Ԝ��_sy����c�h�aXs�Z�����z�su͸�,a6@n��X�9��e@_6HD.�W�l����:�FMz7y������l$�	�"���:jw�|k�o�&�K-"!��p*X�/0چ�2�M��Á!65���k��h��u�u7�9�t�D����M)�{Q4��m����G���m��T�a�Gۣ<#aB�rL��0t,��r
:T.�b��Yד�h���O�E~�6@�A��*���n��&K��[�t�(���)���E��ԄXjҸ?�w\,/`V�n���q�J�O��k������Ūo1�&\@ƾ��V H�/O1��]~z��R���Z#L�
���d�0�Ws���ʪ�r�&����$ ���G�"�L����~�@���rdm0��	[���Zl�V�.���.0c|�%d��.��Ϯx$n�Ȧ��^�hb����/2������u�ģ�UO�,]��C�A(.��-��yXE��<�(K����n#��6�Ȱ�;��B����fov������NH8~���������b�\ʰZ�Sr���Y!���!��IK�W����xSh��j	�&}��Ȝ�F���\ݠ�����oͿS>B°|#�R�7��V�؉^�L�b4�N�2H�J����χ7[ܤ�.I�h��@��iB�q�����cl�5����$��D�x����2�G�+I�STY�R�(�.��]a�v�}�vjEU�
���"&3�d�CBW�_3@O��@W�=�,!�;�+߂i���x��w�>�����Pδf�W�jT����,�1)�!��.;9t�uU*,��u�����`<:� /i���Z�&��U��-F򸕅��UA�0�POz��Mf�E(��s�������ꭨ�H\"L��'|�
�-�n%��H��KңA��!(�e�A%2�m���Չ�����XV}Y���֙(0�����y>H�� 
Ήs1���|�������*�h4+`��K%�C���Ke|�W����^$�}�)�"<��H�
�dȴ����{� �PU�n:�q �R~�72����3�K�s/�|	v�A���(�<�l�w�x�P=^݅
ld�j����A �+�?��B��j�أ����xv�z��`-�ARɩ��ةשV~xn���w�e��#A|���N�Q�ބ��Tz	f�p����յ�~D��5B"{Z����ˏ��k�$s��¼xp��P$r�Rhb�Z�ۡ��I�r�k.b@n�L�p����w��W�ʡ&�%�dD�N�u�Z>�j*q��L��
��g�w�2�.6t��uguC?)<��Y�PZC�(I�*(���k�y��i�C�N'���j`�l���b/�s�����<��V���l+�Iu�Ve;!�n�'��դ
j�yLe%1?��*�\}j(L�W vЋ�����EQ�O�`VJ�A�v"�18+W�yED���,(9l�f��v�!<��=�.u�K �^(��܍K$3�6���~W6B$P� F :تb�ڿc�����)�O8�&(�=��N�S�}r+��n��N?�66쥨^Dn�ʣ��
&��
P�0d6�ޕ��W�Y�����*��K�i�Gt/��VX����eu�M?m ��A��&�+��V[�::�#�x�a�s�+VyIuޞ&�&����87o|';zf�)��ܚ��#pǨ�I��v�yF�Q��,E �w��=Pn��t[���ҿfM�C��\��8��38,G�[�#^���������v��Ω����L�T��R�!/je�M�̲~�I*{��cʰňc�`y�|b_ �35H���E����>aC��-	�����7~g�V<6�2�tO8���}N�ê��K؝���,c�*�p�B������w��#S^藢��y`}FC8�o�:O.��ŉ��u���}\���E�p����?���L휯�;��&j�	Y��u~��.:	��j\��?O��+*�yz6|�8���+ܝG���	aF�8p�U6��c�H��+�>�t3��\�i$�n.|��6�噃1���MP�>� �����5K�4�]}'\��ʸR�3��O'菢K�F�9��B9��H��w����^
�9 \���m��!��#D�@ERTG��i��	�I�%*���5l�������E��x��_���L*ܺ�������Z��Nfeu9��}� FZ� �,6�K���n k�J���c�
�����|,v1N���ᒓ$�)��RSX�=i좓������	ݳ�iu;��4���q���^��M��_�j�#�v<whp���+rbC����R�4nm����aW��}��۵��UF��,dw��b��zNH���կ��j���ڡ��vy�p��rv�%,c����X�Ln[N��R�.�����b��w�AF�H�z���o �^%�&��'׭�A�<�� :�'�Rz:��g��oEc���! p��Hs �J����F64�C"��}s�&̎Ӿ���g���>B�O:�{K]�\H�+��T�6ɟ�iסɅ����z�KD*�l��_p��;�<����H��  ��"�\��i��q��߀�����Ď�X��#~�'�e ��%4����',u�*A�[X]��Z���l&��"DI��7Y<�۴bX5 lj������	���PRIG��X�W��{�n���0��'�,��AѲ�H����d"0u�(��-�5�ֺ�Z���L�ډ���1J-9��U:�7������1�_�%z҅���!���0@g����Fz�8}k�{��ч��ӊ����<������c��2��([�4�I�li���Bh�B�Eü.���7��־5�eEg]�$�j~��T�K��a5q�>�S>�i!~fW���tlCM��\oɢ�/�r&t���r$)��W�:�>	�C����ve������g����5E�������=^�`~�O҄�Ș+҆�	6XV D�ūM�~=nt�f���:eELY�JlCbJI�PΗL�fs�=<�Q��#|SX8Z�Z�L"��@���V�J)6;�C�F��ڳ;8�_�]e.��l�\C��N�FHՌy8���d��$���"J�:E�|�{�o]��K(H3��U�X��50�.(2U�����s�\�萳@��զE��h���(�7a0*OEUDɚ���M�$��Q�9�m��!�*j8�#[�H�T�Gv�$#\ɲr���0/^��} 
�੽= �Y+h$�<�JY~L)�@����E��F�����t_N�
�)�S�E���ԟ���37�Rw�,jl�����YJ^�B�����6�[�����1��|@����ޠ?V[n����jF���6����*L05���(Un\Ӭ�#�Kv*�e���q������ې�"��Z��[�����m�'	�_[K�zj@.r��q-c��^���2��j�
�S$	N �纃�� ��[\˄���k�#����M����%��'8�����<f�86h���E~���cE$���n�Z����kv;�L��p	�fJ@Ф0�a����~�=��:�ͭ��\.L�Z�}r��{��if�)��{TҲ줐�.�h]�j����E��9(�78�F���޷��m <	�oH�>��|^�����V��������4Ñc2�u_J·��Q-j�M[���4hXq�@
��Bcy�{�z��ˠЫ$~�C��Z�xwc}�M��G(h��u�T��۬�L�.�Ua@��}i�j`Y�
�0�"�!dߕ�W�Z�3;Ժ�hd�@�����dk��i�DDxq��9Gy���P�7�Ú1�� �ڒ�,ҙR��-��_9Ϻ&U�7��;��:G2�;��<u;�/���6JZOv�I����E�3I{��x�A��P�����f\��(�ߛﱖ��d��{���\����"@lfM�-E꼱���P��~����]����2>ܽ�� ]��Ө}4�n�u?(�:��?>��� ŒsL�9���o���H�e��4�Q��F6��7�+�f�ْ�䘪���츝d߽]ͻ�8p
5T\�o�p����{�Uד���1M �v�~��p����IwK��5����v��������!�r����*�@�ql#l�j*��{��f�ķ&�*�~�3$�IF0x"isz+9Z-�gv��z:�D�nVy���H}�� �J#z�%�N��>�q����f�W�ZU���#hD�QB�Zw9L�M����k��O�:�/x+�P?&�R�E5�͡�耰�.]�nƧ�Z���7@WM>&���d��e>��q��\=���[��c2ګt�ҧg7wC:<U�I��P�(d}*������y�ޝ	IǞ�`����r/'���ĭ<�
�9�+&�I�b�e�����M�a��
Ej_L�^�?�;g��Ej`��(, ��k����Q&�g`�!?�<�v}�8�@���f�G\�����cWWlj�|�q��!�͝=��N�f�ٷ���$nO�F�y,!B�+  .��Y(�:>��}*)Lc8�3��8R8N��|8���!�	�nt6�����D�����^�e��B ��K1��Y��2+>�C=}����%�.������r��-eP�z�m�k�<��&s�葂[�ݫ����<���f��-R�!��<c���<|8��z�@��]{�!�`�C�M�٘��Լ���G�R��2$=+�ٯj�qa�fH;������h@3S�"�ֽk^o�Ȝ�Zb�,�v�$d���ŭ�lT-C�RqT8j@<}�p���yA{��g�H�b�`���bڝtbݱ�ƀ�j�~>\�ֈ+٘]Hx�\Vg6�
"t���}��N�Q]��ܝo�f,*s'*	��B�^ʄ��w��aSYA��Ju�`8�/8�jc:�sJ���m�3�#�k�x����pϸ+��w?^sj��L(����&e�LY�u9-�/���.�n]1\��O>��+%h�z�u_8Z��F��L���a��pt���A����HIR �Y���R��7�:$΃|7W�����1�.�M/Y�;d�P�p���4�}\'�C����R�����?�������	9�A=H������^et{ ˬc�O��Uo���>�{{�T�D��d��	�%�yT�P�Ȳ UjʻN���R�����R�*7�+�(,�����g�u�i�5�� ������6rc�T`Kk�s��e��g9�1�,p,��4����ƥ �mg�� �nqK��J3׀�q��F��&m�亂���J���M��������'v7��_��uC����"7nH� ��ٚ�q0��N���'�հJsd���bx��z)�˼���Q����Y���!�1"�p	��r��%���z����N{�����2�}�aw=�F��p��
�"^ ���{㭢 J<�o:@��R���0�*��c�#�k�p{8	H��jJ8�!j�~���
�&����PkE�"�l�Y��O���&<�\�l(��Vp6���i2vd��_��[�*��[lV�I_O;�<)���5H�z �"9��D2
q��G�Qf �ܶ���Ẍ��>�c'56����4Yeƌ$j�pZ�AY�T]����0���-p�D�D��27��W�<Fba�� '������hp��o�>I�wX�p��v.�n�V0~�֣+������#�7�=d��6�#׆��65�x�u������d������&룻�:�8����L�Ҡ������!��0��ۮڇ�F���8#^{ ���L᦮l����<^�����G��bu������h�G����j����÷Q�w����kS��C���m�]�2`���],���F���������S�����~A:׼
.HI������B��U�tr���25h�=���wΛӖ��z�dg%����(5 �r�CB�����^��*�� �����+"���9V��O� ����no��D�ٽ��Lt1J�b%؞�����9s�"e¬��ދIXSa�Zx7�k/��?���Ea66�Ρ�Ð�N�/*v_,�2.jl��3�p��FCP�y�a=���$٣�"���: w�|��o��K#�!�S[8X`q�0��2Є��'���B�N���;����ho$N�C��7�F�*+�D<��15�QQ�WmQUA�EQ����#��T?��G�D#Wp�r��0��
0�q�<xYM�vh�48�Ex�~��@Q�Ƴ`Nw�=X���D�mt�`�G�)I0[E�\�Ժ��ҮyQ�-	�,�ڕ28&��a�J��U|ߒ�()��Ǖ{�1��@8���s+V�H�;׋�{��S4����'�L�_��$�����d�7e�ƙ��@,�`��Zk=����"x=��W�v�/�m�	�X�{B�u�.����,L|c��ڿT-�Z��E��$��o�����P�h���M�洑�[�܈��ϋ߫"ѹ�>�ظ�q��S���EYY�_r�A\�n������&6�;�X��Of%*)�k����~ޝG��b�h�\I�sZc{r~"��ߧ�㧃v��w�a�h8��j���ԅ�tcs����F����S`�(a�$�EoÖ�>�w�|�"��m�V�hQ��S��s�4��/2><�J����~�Y|[Ҝ���?�h�(@%D�B�t�V&�R�ޠk��y(��A��x2e
�h,G�ĥ�aCT�G9�^��.a��}$pO{}"
v��"�@�dSWN�36������@ʹg��W'��B�i8��x��4���x?�PDڋõ+���X�V,"��W��@9*�U�e� 4��A� �<���/��B���Z�!e����-�]�t��A&M�P�������f���(^XΛ
mn�z13Ơi~SI�\X͸�$L���- �R��t������YS�Nj#��e�2�j��Xi@���N]�}�5�(f�ĦĹ�>�K| �wsgpC�r������ܠUb4ac�A{M�_��z�����M/+��r���r��X����H�
�c��*�M�( 8����U�ؼ�O ^~��kM�ةϔK���r�tv����Xr��m���V��+l>�qj��-��!ġ�����B�y�⎤!���x=|z��_-]�*�|w��LVt�V�8k���K#9�z�N��܌T}䊁�f�^���;7���D��B�ZR�N�W+��2��k�����łx�#ePZ�CR^�<&��-���y.XZ������*���PW��f&��)d���9D>�Eql���dЛ�m��2�H+tg�v�C5o*��^]P�ޒ()*����;yCW��yH^D��i�`W��*�/�Zl����<(Y�����!~�I+K|e�����R|��R�
 �L۷�?,���d*j�\(ªf �\v杻��cQa��`Rl�7cwv�#�8�Jܫ��:������C��Il���l �!�6N=S8́Kx�Tg⒫�$�Ɂ���t!�B�Xq �&��p$ڵ8,�XX�)���83`��3VNO�R�"�<�L��ٮ�����?D>&o�������U�U�f��Ԗ���r�~�E�E��� =���ؽ�^��s��vje+Q���O�'�7��&�|�L�v[Ѡ%��І��ġ��ޞ�ї���Į|Sclz\y�����\|�����O��/S��d�bW�m�=�$��ɸ��fC�"�T����U�3nf�Q�^Jx��/-6��,6v�qu�v���hTH��R��j޼�BMҟ��{���f,��d�`�YabU;鮢�(�����>W���mߘ�F��g��6��t��q�1�N���]A�*�X,E�\*��zB��0�w(R�ST�x��u`�m�8��:E�r��C��n�e�s�s�z�&p��u��?�<���GLc�ͤq��&`��YLzu��?J�!$C�I�\&�AO٣Q+ B}z�
8�at�=����<a���pY����H"�tk)�V��$	�|�3���Y�1C�MƉ��V�m�����t4$�o'��<� �R;HN?���ż��<̝�1!9�>H 8����%^�9 �>�1���ਾe�����rT;b�_Um	B
�%�u��k2�{+�ʖ�(*3��R�����G*��*�p��2��D�wuĺ=p6� 9X��_�6o���r:k��]��~��c��l�7,��b��O6�HV���Bw���D�3�a�I��7ͯ�}~��CE�����̴�����T�M�o*�Ռo�Y0Fv2�&'�С��Cô��Hp�n#�x�*r%���v�W(�k�"d��Xb��zx��M$���v���D�W�����`p$��rl�F%����C(�Ђ9�Nv�����;�w�V=w�L�F�쭄�)�ܥ��^��n]߄<��:��IRǫÔkв����c����=�p6�(H�BwJ�C����֙������>&���4��u��t:O0��;�\�F�.x|6�)�i�j��W���D��h*�K�l�i"_��D;�\Њ=��H��i 65�"�����{q7���]:���zCX��Y��'�&L�{�4�` ���Fk�A�&�]Y ��K4V�bi�e�D���7��k���b�x0 �;���+����JܺI��X-���qz�nQ",09*�F(B�7T~���-rtdXW0���'5c:Đ���B-��?/�����*k랝�:CZ��CN5�gp�)��}U�!K(0v:���4F0)Y���{;b����O��n.�W�<��}��Z���-u�ܜ�|Z�*�3�"���2�4�x"�ò���3�ЭY�鈪[�]�����Tǩ��A�x���^�S8>5�_(�~=>�E���n�����X���Y�t2�6rƒ��%�x�[�y���:��h�S��P�����6f5��~�;���^��O��~�T+=TŇ��fV��+�;�2�R+�njA���wz����L�m�J�.b �B����t�s�'
�/4���CXn��Z�A F���$ե���E61~�����P	WJ<_��.Zl9}X�~�F>�ky�[�����$���"k�:�&k|�Io��TK�뚮�OXB�0+�+2Kp!嘂$�������D���4�h*� �^��7W}�1CD?�2������QE�m<�`Ƒ�>T�ZTzf[G�>�#R7<r]*�0�!7�U
�Y���Y���hZ��@
�~�O@ؾ�{�nUB޷�qM�;t�E�����)�,EF����u�)�,��,�����!���RJĈ7�*༒�����Vaw1F�Z@Ӡ���f�V�z��G�����C�r
��b4Lf�����EI�����RG��A����6Nn���@��т�"����K������Km�v�	r�T�Q�p�.(���犘c��~��-T�5�̀�%$?���؁�y�����Ȅ��ǂa�K�6_����&3Z�����'t�rƂ�n���gME4p��ٙ����,nERGA����;ۮ�f^�f 4���_b���~�x���P�#Cd\d��Z�h�rY���Aꌧ_;��q���h!|���hS�jz-���ʹ���m��F����m(2����?'�o>2>ӂ�|Ԉ���.V�I��o�f�}/4�w2�"J����������[�H�?kh�~]@@�GB���1o���x���Zt�6���Dx�[�m�GA��msT
�j30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�&ڜ4�z^�27лXo��R�|n�?S4��{2�в��3�i��R����@��r����>x�<%Vֱ)#�׳��'Z[�Ϲ,@"����4����Z��mg�U�f��Go�����X"�q���D4�y���O|�:�G��oT.�t�U���8 N+[II��
U�v|#r!��HQ�I1���7 �dI -/�,.y��1#r�.$�����S�����ڮs�
օ8�9�$���q�|:]���;~"喢z��l��&[@	Z�H�đel+R�U��]��iu�V�>�5S���f{SN�:D֙��c0���k:�lj���n���L0T��O@�x�8���k�m��?"�]V0|{��E&쥆��kx���?)
�Wi�x�l:R���E9�	
e}AbP71��xS����Ҽ�S7Z������Q�,+��3�4dԦtrTF1,�ߓ�O�e:���`��r�Hn�~��y�o�Cʠ:���g�L�9�є�ʵ��/���S�8��٥9�B�a��:"t[��A29G�r&��5�$���O!�aT�9��ai3��[��/J;�If<�7��_�]TX t)Z��H������;��t�����zL�UH2)V��WH?�}m+�%����9��4��H���Đ����vh�U`=�x?_��Tp�KТ=0=���	S����&�aO��g��IAA�0�w7�ɢL���=
��p}���#���fm��V<ӷ�S=��?6�s�SI�-Ḥt+�bR�V�;�,h�>�����`<�QY%m��G=(4����w�<�}�僾�����RՇ�B�pq�a
ܨ��?!�}V�dB)(�O�S`N���W�{���L"
�]�ohw{Ҋ��{�7d.��Q�W��\��]����藷�1��c�G�d��	 �)�\*�a�������1/�v�m�cSǂ)�'�?�� �S�=��p����'�>��Xs޹=;���Ҹ�]�����U�p��&p�p���=Ta\�7��	���r/�*S ɇ�#`����0�t�qh��N@>m)r���m̄�5 #޺���<
�y5Z��[���2P��P(c)�m�+Z�̇� q�/^n�=��q&�z�*Kٙ�'.�*w�k� ꕳ�s�LSt?;�&G�/��8l��WYN���?!���s����[���:;�M���r>�݃D��\�?q������^�0\CMaY����Z���!'�=(�M8��gm?)�쬩0����4�OU��'j��,��
yS�$�(�-{E�½Q�4� ��xo���2�N���^��P����F�W^��w�RrFT��:����"��H�s��N�IA��>��A�V��@s^`_8%-�j���U��8��䦭���=�Ez:9���4^B&��#�zb�L�z�*�S�*�*M����k�aB搾��
�TB�p��C���赽W{�s����?�V= ���i�uL*��F�A�c�.��m���I�Wk0�iﴟ�߯�;1�*����CѪ.D�a�}��??�O�'�P�~�IC:��M׆�b�'T�����^�f�P̶�uY���㾓A�o��Ɏ����?,�c�:��j���.y��GŖx)�w�q����)�Gn.[�r���%����������bI�<y�y����y� 	���%�B8�u��^��T�3���ĉ5bߣ 2�"{F%�<��R4^��C�2?pT��Hvظ�e�Y/ur�3��0�5w��$���f4u�$�kX����6J�Eթ���AE�a������J�hW�EV��]_I���W�mK�w�$��x�Ǫl�)��K�_�,d�>���9��C�9C������lE1T��������]�p��'l�9
��~TFr@7����Ԏ�9��tѫ��؁��"�& ����C~�m�z�e)��$���{ {.�l� {|E����nd�hz`�@[R[_�<v��06��i¾�{�ǺH��uz�Z������+Z�o��>���/�M�+���X�(F�`�b���y�UfU1eEh0�.�c}�62��o���*s�I�C��{�B�|���.�h�ؙ@�_mKs�T߲)�&{�v' ���44�~U�%�����2�N�����y�P�S�>ò�U$U�V'QS&ܑ�/��;���⳻FG3������\��<*�]T�T/�d4"a�ī�����	N6(��\7<DrN���8~�F��W���,�V	��ZN�:����ZP�d����Uh[�+��{��i�,Ga�' �[L֑�4��gC�hg5��B����T���P���,+����#��u�J�K�+�w����<�O�(r���R��%z�@�J��گ�$,\��v���ɤ��� �5�2���	h��`/([T�q��2L"ۤ��jIc��6(py�I�r��_�M9qz{���GVC�g���/K�O�L��v�.)v��3�To/R��XӮ�� �[KY!Ѕ���� \\u�Q%\ef�%XIUa}w[�����I��	����â�%Or�6a�ofJ����I��q�����v���^�c��n�-����ȳ_A%Q����k�{�o͚��	%�g����yU}S�zf�U�ǭr��?�~�N��B�*�j$�致2H�f��aK�֒x�۳��"����a������8%R��\�=�p�1�V�E9�҆�3rYR�M����ZH�s\��	R��8_'�^y�Mg�����7�S�"�,����F�t�,�� �g��l��?������-�A�IQ�st���r|����`e����/��A��h���v���bI��΅_=�B����{����(�2�9����w� bm�Hl,v5k�v
�68��(X�M`܊�Ŏ��;����c�V�9�B�{���NO�ƍ�ρ�P�򛂁�E�����Gu3����p�����~2�[�i!2�k`��_���3j���܁����$n,�jM {06e��ߩ�c��2<q{��^��ڱ�\]Ä�e76ٖO�:H��Zgqb+���m1�1��c~�:C���p���],og���]�\?��9#"�P�9r�����$1�]��t"��/惥.��7���ܬ�ꌿ�O-*�2�1���DGڟe��7x�><���%\��<���{�B�D����֟��`�.u�@A��6�0�V5��;�bPx�%zX��p����3�x���Z�[}!�O'���~�vp_H=���6p��Q�cm���&��	+튈�X����R8�U3%"���������ǖ���� ��ROV��d(V���p�6	e�����;x��E0*ty��:�,ʬ�7;Qٌ�>_N���q��g�Ky�-꾧I(K�����bS_X{T,���]���t6�5�7���`��u��9S�\�حM���)�d�6�-�4+n�.�`�{��Os�f�Q6��;���~�-b�<�1��d�Z�j":������n�;̍�~k�A���25;���ˏ��Y\�{�M�j�;Z����qIݹ�~� ����MnG���'q�*��&��*��2��y������ns-�S�8΀�{[���@��0i�v<�1��@l��Pz~̷�Õ���a�ȵs��qG Z\Ϲܱ0"�v�ǕO,�ZE�gL�vf?��og��7�"O�c�6��4c�l�/�s|e7�����o�t�T���V ���I�{
X�|���!�$wR�!�����r&7��IН��ܴ��ve�s$�#"٤$IZHֆ�d�Z�W�y�:/0W��� �#3�;��^�uKXY4 6��a >��0%1�Uβ���2;!�e��J�k��+�����O<�ϣ��΃U��8,&X6����n�˜��;"�q�v�$��׽#��{�)S.�h�v�&�&r����kh��Env�$�Uȗ>��������#*���f���p���������>
�#UöPUTUoe�u�NF9mS����9vuݶc����eG���7�TV��1*N��y�,���ӆX(ez�^*�L37kc68n:?z[^��'2�U��W[�^�^��D�LT��m�·?��D�+F�v��Ю/��K}�)!/L~�>�J��:��O�V+1v�k��^�}��X^]j��~��4�%1٦��*���|��&���� �i��X�|�HxGmDE�<�A�͜1�® T|�%�c���o|#Z�0i;���ͷp���䝟�� �\���+�(���ZF�/c�l��@W�ԴseA��pv��p���h�	�@8�]ǁ�9�B�и��d�Y?R�F���%������o2��`�V�s�,SH��ҸǸ[�\��a�t�{ ��?
;�h��R	q�[�M����݂�l��/5b8�v���hJ+����P@�Y�n���Wx5e�����JLA��M̐�4V�FH'�fI�d<s��>U�=IR����/a��#�Ny���� ���}��wXL��;Mv����q�.��n3.�����[�:����k ��E6v4u*[�xq��f�������qQhaØ�H�y��֤�!~���h;�mذ�B]���b�b����P?*���hy���Tb�*�oa��n��w��>��j!*�3z���<��K��j'�5we�|ubɀנ �1Q<B;�櫄�2T)x��١��a�@��-?:��Q�ڼ��P#w(��5�+1},9�'�wUR�va��o`t8�������+�X�ϰ}�א<��!=b,F��8�U],o��{�)󱉒��s�Eaz��]��a��is���`�?������෤�	zCn1�qD)�/Z����71d��pP�J���~z��Z�;�ב�>�~�<�]`��F��9�r
u���A��(t��n�
�#��}\���F+�+��Xخ�wI^ڠ�M�A
a��k���=�_&���ƮmR�]������#�(��2��2�����^���}&m�!2�P?�>N}�GQMU�\T�W_��yz�� �>TQ��u^kGFNZLt�������!g���-�T��p������κɮ�:���!���f]��e�r��(�I�u�ήNNӓ'u5�u@�ߓ#hK�B�����|k"�8hMkb5;�W��1���qw�-��ؚ�;��ςb
{C9���z_��ثk�GM�����2E�0kH�b�̛�9�t�ԌC����ݚZ��%t�$�{��@Aˉ�J/o�:��a��N��-��D���w39F���8�/L[���ږ\|c��d<(����'�&(��GNP`pR�@��Xc�N��͋õ�+�t#}�=�G|~W�p`��qI� �paf2��m��	��=X(�c�2�Jg�������5�+/��ܓ��{u�o$`�9EG�xI��oçi�Wf��!��Q�a�rk�$�P�)�u��5����~�' ߻y-�P(6r���}B��˶�}�rW6~�,c���� ��x����9Ly�����C�P���"��{Q��2�F�i�#ؿ�����Zjف}�l��2A��J�p����j]\�wf�v��0E� �N�2񠳗 D����WS����x�cӝ򶃄E���Qa�_yYo�{=o��ͭ1.�_PV#����4�XG�UwYV���$K6+�Ū�l�303�4���X03�x����͊`Z@��|��3Q� �z��-�DD��N�M�@��ez1��"��1�?Ú�b{�6c�#�ǯ�����?�x�v�_h6�Z�?����n�0K����.��������P�9e�5xri\�����wڿ�晢��Q��e�ƭN0�<�m��ˇ�G����͢\Rr�Ē�/��N<��3�% `K�����I ��"� y����*�|�uM���h{���ͦҋ:�M̙���8����u�[�:�*�GE�PFT"�O��S��*g������lA7\>��}왰O�N�TB~ѡ�l��b�*)��\�!M�\xh�ԙ��͆�a��s�_�)�մn��G�b*z(K�sօ�I�������"��H痍��fe���d˙���U4X%3���A��~�(5Cg8�v �j[��K����-�A��ls��0��� �)b=8C�j�^�3�|	&���2ĽU`�Xjs��,�h�	ܮ�H�^�g]AR<gu���Mi���V��5��2w"b=ή����
.c����d��k<
Rl���S�<���0V@3O�x6�SzkF���e��D�|=��E(��Ex�^<�O��
���i�g"��E��E�E;r
�z���"[�����TR�>j�7���V�A�,��FM5�*��$��!q?� �����D��Ȥ,�Xiџ̌����:�¢0��WM���#>N��q�J���u���K^��$SkZ���x�������mͻ�6�`X�w%�~0��2����R�UF��,���r�jR��:�=�Yn���dr���[�:~1������C:*��t dLdU��S��ǟ�����,�$��˵��a�b["�Д���9�=�&�<�5�}0�O�sa��0b3��j�-�<;V�<�v��)�]�j� !a��Y)Hƴ*�q��;�o����0���L�Kz��V�H,��m�N�!w�9�/<�eN���w���$�k ��BT�������p�T٢�_/=��9{OSֶ��۷!>a����{�xAV�X��d��O.�+�����a�xҍ��Gm`MV�kƷ�=�ɦkO�=5�@��p{�8���/ҽV=��;��h�w���AӰM�Q�N��^K(����[h�&��}8��*�u���R���Be�����
I\��LB}Bv�:O��XNJ}�W�Ls؜C�
Q.�ouU�*���NdNC�jn�WԲ�\bj]�	���Rb1}͂���dݑ�	�*�����.�K�D����1��hvE�qP�w��*�§������+�ۅ�Ыg��1�E����5;_���F]�=���~��.&�{e=�q��d�}	`5�r�KSX����j��G��al,���/���@R�r�
p��i�4g#+>���);�����7�ĸ�k-R�P5l��ZP��t:�q��^���=mv&Pji�7��A���w�:kϩ_�"��s���t��&��<C8��W��o��?!�'sN��������G{tMs
ڎ��#���ť�z.e�qVߞ�_�P�=YwM���VE�X�#@�'�j���k�7��?6xE�Y����$�4���U�'���,�y���5Q�(�,�
��4|8����lƥ�	��m��.7*F�rӾL�R��0�$�ܢ@���s���SG�0��胳r����m-`,��-���Aŵ8�C�1��	ʗ�zg��ټxB���#���Zz5���@Z��v.��s�8MJBSk���2�T��?���y1H���V���Y�����48 ���i��*5���+Aj.�:Q����NWx�*i����,	�;U�K��C��3D�����E��L`�D�A'+m�P�8����C/	^����5�T(�+noz^��P�su�Gz�k�A��,�6����~��}���0�W���tNXx�yj��/������ź[�X�y��%|���P��[��I7�ň���ђ�͒�Ð۴ԩ>�c�o{�uȽ^�r�@���q���fy��bl"�n�G\�B^.��C��vp&���7��3Y� ��`�_0y�I��K���"� M�f_��X���r�]J* թ���J[��n!8�f�gJ:�XW�=V0�V_v��$F^ځRw�$j�����l������_��drXx��I���9�������l2s0�67�@-��Ʃ����'y�9�'�~�{�-C�4��g�k���+]�.���o/U �C���Gp�G�qe�3h$�z��(�I.)�� h��Eo���vB�!z�y�[_��c�F��\��������PH�QxzE����f�O��+��$��e���{��\g�����n�	X�W���p�bT�Q���y7C�f��!E5��.�ޏ!"��l����s���о�{*��|\.�����@���_�kĈA	()U�1{Ў �/a͡FM�A�kU����[Ȉ����L��py�������ÿ
\U���p'>�p&is�/����<�� N^G@o ��}����<]�9/&U�4�V��1[�Ǖ.	�t��>q�<1��[s��3׭�-�Ĩ��91	�\�N�K�����Z�`��â��"XƖ�Ӽ{��O��?
�t��H$��I
���yh4z�5���)�s������[{��R�
U����L_�J$o+�����9]������\�-�b�g�P�)Jl���r�\j����l��C�ō��_��U�v�d�(h_�q�r�2�$!��.qI�f�6UkBb����_��q'E��G�C�P;�Y6K�'XLY~e���@�1QW{=/��bX�4���)�K�֯�R����\�*v%	�fNX6x=}����FIS�������С2%�R����\&]�a�w�۸F�>1&�'�!2
ğ�c�`�6-���U,�Q���xTB��	c�c���������b} �,fk~�Ǻ�U�,76�y����j*F�;�F��E	c'	�'� ��M�DD���vN�\@��ezg��"}�1��w���L{�E�c|$��e��E��?�]�v��h6We��;�����n��K��/�.p��Ғ���&9e��xr������w���)��CD�Qޒe�|dN0@ʯ���}�G�ⓃC�\�ٛ���/Z N<73�[`K�#9��I A�"� y9V����|B�uM�	��I��q�ͦ�:�CF�ɓ�83����u�QF:��GE�FTX�O�%�	����g�X�� �l��\>�}��oO�D�TB46�����b�)���!�\x���
/��͆�������)���nٞm�b��z(�Qs�W��Y��%���49��%�CY��W���[d���J2U4�A%i����A��~015C�O�l	 ��j[K�ӄ�-�J��"��ܦŮ�V�)X�8C�j�y��3�|	W�q�Ľ˔�X�6��"6�h��	�$HÔ�gSvR<I��;�i��V��`5��w��=����Wc��d-Lk< �l�d�Sq����0V6�O�Րx��ى�k<���\�ߺ�|=��E(y���x��ȝO��
��i���� ��{�E;h�
�̥�%�XL�����
i�>�7Ej��y�A�,�Q�M5����Y$�}�q?d$���&�D�Ժ�~|,��7џ*��|0���J�������r>N���q
�J-�u�o�w����kZHΘz]�܎�ஐ��m�6��XL�%��u��h������U���,�� �r�`X�J�:���8���ur�}+[^a~1����8�^:*t]�tVLdKU�S�t�=ܵ�;l��"����A=�7[a�X�"�ǫ��6P9�sO&����}�bOӿa��0˓3�WӲ- �;L<�,��)A�j�1 !W0��H�*��q��;�e���{����L��r�ߘV5�H,M�m�Oq�!ma9���e�w���x���k���Bʏ������p�
����$=㷴9qzS�l>��-�>F0��d�{��AV[d���e�O�+����8�x3��=Zm`�V��緶s�ɦa���j�@������8���/��V=�;�	4h�m{���^�MQ�����T�(K&��ѵ�&��}8�v�*EW��ak���B[��ِ�
I��Lx�}�BvvrO�k�NJ��W�B؜�
Q�2ou� 7���dć�j��WԨ�\b ֩	S`褈�1}�����d�	�`����q�.~�Dj@�V1�~CvE��PB肶`f�$����ۻ�Ы]m��E�A��D�;U���Y�]����5&���{۠=᧴�d�	`�~r�}2S����������a�޶�1��'@!r��m���4��#+�N�ʟ����-�ĸJ�-ȷP5�&��ZPO��t��q�^��H=m,�&P���7G��A��w�xk�T�"�Ms���tM%&�e�<y?8��W�~��yI!�s���G���c6�G�xMs e��k��Z��.[�qV�s�_f��=�QM������#v�'�`a��Օ�7
|?6���Y�q���4�`LU��'��',�y�Z��5�R(�y�
v�4|�n��<�b��z��������7uFy�Ӿ�	R���$��ܢ��B�s�=��I��0]?�)��.�m
1`,�J-�g��w͵8�R�1®�����zg�ټ.�B�,�#�е��z5Cه@�ǆ��7��i8yBS�ħ�hYT�L�?YW�y����5�������êS ��>i���*5�����Aj=�.�:����Wx�i���,�;���KoC��%D�O����L��D�>'+#�Pˮ����C/���B��ϫ,T(�7ne^p�P��;u�}��a�A�W	�6p
���`�Ȧ��@x�W�F�F��tDx�/��ޥn��;���y[�'y�%|���F1�[fRI7Xe��3�ђ�"��y��*?�>��oqu�s�^(�@�2�q���ã���"���GR���?^.sjC�5�p���p׸���Y�6�`�k0y�����,���2��c�f�X9y�r��J*w�ٯ�Jћ�nW�f�J:��Wߓ�V0�g_v�:�$����_wPW$jz��ll�D֍�>�_��dr�m��:�9���ٖ�l2��l��@#H��_���~�'y�|9�?~�1-�G�4��a����b�a��.���o�� �����Kk= �G: e���$ɰ��(��.)R� h!Eo8;��lh���z��<[_F��c�w��a�֕I�%����H��zEw?���&�O��+������������\]���enK�X��P��f8bT�M��|,y7y�f��	E5k�.���!X#�lӹ���s܄F���{*�|\�@.����@��{_�!l�A�)UĞ{Ƣ ���͡�6�A%�U��ޖ[�ň���ۂ��y�n���k�ÿ@JU�Ͻ�&p'>-;&i�/������	� �sG@����s?����<x�]��(/&Ko4�Q�1�8����	�j��>'�<1���[���3�B�6����9T�	�R�N����b�Zݖb�Ø��"��I{�ٕ��5�t�s�H�I@��h40B5]N�)Տ���`��}���J�@��~��L�J$�+�歽�/����T����-��]XP]lJl~#����\j�����ֹBōQ��_��U��d4�(h��q�h/2��$�ؤ�I�X6Ua2b`��ߒV_�K1q';���EC����Yl�K��LY4���6�g�Wq�/�pX��6��_K����R�=�+�\�`�%	�8f�SX6��}0��x�ISk}��� ���(%�Ho��P�\�/�a���ۮ��>�l�'F5!h�ğ�ic��A-���3,ɌQ�x�����K�cU��x����ў��} �fk��Ǻ���,-��/S��O*F߳F䗴�ɜf�aK���xD&��9�
��P9a��k��8�#�d���Jgҍ�v�Β���n���)R9�"���;P#�������wR�g_�^�g���0^S�O��?,E ��P�+t��}�6�;g"�lr�����J�AS�|�7tw�1iN^�A��NS,�f�/#�1A�Ȓ��9���1��1�0�o���j�OD���
�C]�(�+������۠�Gm/��,��>�#��6�A�(E����:���&;��7��C
���kb�����x���ӯ�X 0��3b����
��t�8�%���������/���
,�%@zO���J)���kNa�x�N��-><?��w�,�����@�[����爆c�-dͬ������:�y��Dr�6b�^�eo�`7up�<�C�b���'��0�2��D����q�l�
�е�c�}X���/��SVR���a�b{u�"K7�b)��v�h0�|��xt���)0�o�=�{E!p�QB=�R�������h����!fjX���+�bRuܟ3ȣ�a?H���H����c썟�! (�]REE���d���M��*�K�>��&G��_$��|v0��ykM:�W�}�WQ6�H>\�-J`Sɏ�g��Oyrx��AsK����'�KS\7�T��}�N4*K�7ӄ�`uE�QS���JYƥ�Wd���-dw�n���`sQ'���	�Q�e��xFx�rr�-�7��ǐB�!�Z�Ǩ*�U�FE�0e�Kh��
��k�mPSM45�T��^���@Y��*���#����r�e��j{����8�/n��������wE&����$L2D�F��？��n�M$S�`��G�8��\�Ȍ�iEo�.]�@	`����̔M@�i& �~P-�r���"VZ��y�j"��S(&�̩Zb@�g	s2f���od��ԋ�"�}��K4�4��L�_|"u*�Tv�o��t2K���s ��eIvS�
"M||z!'�O/���J֯�~7��_IM����H������3�#�j$����ȯ�A>���,�؛�0=�|<�#0CW�78u���4�8S��~�>���0�"�U+�G��	!�Z���ґk����)5��l7��`K}�����5.X�Q��W�K� �%[�;?�a�aBj��׺�C���)��Mh�vu��|�r�mR䣤ˉ#�8v��Ues�>K|��,�b6���_���}�m���㌜�d>G'#2��Pғ�o����Y�9a�䋡:���
��.���ue� �3�����ֽ���*K���"5��c6�e�y�*��7(��6��?wk;�A7��W��n۪���8LU*mT}?�NSDo�����,Ћ':A?U�F�L;���h
�����G�V3����v^�I��Ej9�m�����' �:�P���[�?t�ל�� s
ҡ����x�rE��B���!6�_ �|��yʈ��AL]W���lYpl ��q90-`�.M&�t�e�G�����|��&kdJ^�����,~���"�O���rJ�ƽW�<V�L_�d���V��w�'�$�H���0%lp�����_7Y�d&ݠ�N�����M9$~����llf,7r��t��z���'-w�9��;~U��a�J��_5�v�FO��c�є��bUg�#�� �����9�6���d�e�*S$}X.�\��.ݶ� �	,E#����Dvuze�[bO�g���B�
�f�����z"Hwzzy��߫L���m+[������X��ǐ�̬�V���XK�š��Mb\�-T�y�6�f�:�E�e�.MI9���j��A����sP��&q{^l|&�.9_(b�,@ 6�_n��u>3)	j�{G"< :ȸ�������U�Is��������<�T�yj�������sAU���j'rԇ&7�/�@հ����T�hG��}�ر�]��<K<]���/Z��4�Kv�e��{�8	/���<e���g'������'N��	�x�N���/�BZ��������4��F�{b}N�P��(&��|?���)��Ԉh�ʛ5QN���캽׮������
4�l4�J�|� $�JXʽ+Dr��1��=˷�IYw��VؗNY���J�W����7\�����LŤ
E�A���	�q�k(	Aq�R82MK���I���6�EM�k�T�_v3.q[ �̡C�V��K��Lk��������C�/S��X���auvK��p�|�<��\60�%=]f�a$Xj�}��V�#9�I2m�+�铄%%0��7�l��������c���!B�[ױ����@Oc�/�:L)-^0[�<���w{Q<���,�9���F�>#$x����}�5�}Ԭ[f�m��n~��`�x����B�*�n�zt㴳`ZfC��K�xx�З�\��7�a6�t�28�.l�'����2��f�F�M�9�7�t�.Rmб}�Go��4���-�R�H�_H��^���gA���P#��m� ,yf��
t�pߕ���gV}�l&���OP��.=A�*�R��t�Y���t�.}Κ�/�$A�І�N�.I��VC�d��ʽ�&���6����(3�,�z����ˠ��>mc��,7�1�WA69>l(y|M�h�&��d܄�"��cU���R�|���oh���J���ʿP���"�u�Ŕ��C3�{8���������O��aE!�÷`�&����j�y�ܢ0Ӂ�1n�,M��"6�V��f<�����3��{���"+����B�Pʡ6z��W�H�v�grF��3�1/�.����՞���^k]a����a�(Jɵ=��"P����W�E�$���]�{"�c�/H.S8�7�h[�]���-�O�).�����$aDh�[eS��7ٕ?<�*�ƔF����gE���D
�~�U�J�n,d���_��'��C!:uV6��\&vb_ư놸��F&��=f��􊔰���\���16�S� ���Bp��=J2��OZ�2uznx��G�+J�����ĲR�z�3�2��k��<ė��G)Ɵuxa �R������d	�T��d�W��/�ǟB$줙	i�)cP0Μ�y�\�:�S���>�Qx�>��.�-��g�<�y�I����K=����S�|�T�q�q��I|���7�ȵ`�E��SR��.��e�Cd�<9-��6n��`�5���M���,-Q��H�ܼ2�V��-C������q���"g�P�*#l���/O��n[�k����yo5|g4t��Y�����R��˛)�@�N�O����n�{�������&�A�K�{2(�d�i�ͼ�L�nT�S�3‫�x>���i��a����@����x���y1�bi�֓��k�Zlu�]�"P\�7Cӕ0!gZF�CgmS~f���o�kg�A]"��0��JG4D���0�F|�y�8Joee�to{�@x� �TI�u
�|�D!�[�� ��z����7q %I����ݘ�����#��$�V��'�s�%���84����0x���`��#�\ɨL�u��\4�q�B�x>�O�0F��U���U� !tD��3�mk�|5����Ps����PDי��X��>��MF�/b����;#t����eT��XQ���t)���h߱��Tr��������vT*pUII�>��*�y����r���Ƀ�����J��w��0r>���#
SP6szof�>�o��9E,G�,X�	V�Wgݜ�& e($ۦH�%@t�ۡ�*�O��M��3%�G�e[�*�)l7���6y�?ۤ��%�����BW�4�?������Lu	<m��?H��DS��
�o:�����*�[L�\�Mg�e%���q���|�LgZ^ҭ��y�[j2C����y{��%�v6Ӹ�+ ׀t{ �*������欵xȦcE3��A��}���� u�&%���xc��� ZJ�;xq�͘㒵g>�Äў��w��KL(�Z��̿�b_ld�X�Ĵ��/�i3��̬�D��$�8p�؁���B�5ٴ�i+Y���F�v%6��60ioړ��A���t�^Si@���!�[o��\=�����F� ��?��h���	^|[8��F��~R�l�v'5Ct�v�Y�h4�ĥR���mYW��} �m�5F�)��Rk�r2;�#t�R� ½7K'y����A�s�U�$/a=�p����Ps�a����M��/0��Yl���L����T�$v!��2Q}��R.� ���W�:F%t�H���Cڵvՙ�[�1(�Έ��w���}@q��X��B�H5�w:>��gu�x���n6�c{���Db[[�-�1*!�@)�c�c�b��+o�[qn6�w?�<���*I��qQn<����L:I�#�F�vK$wd1�|����!@���QW�����)��v:?�����|}l?��Q|@��	��#�tݢ�+��,�1���=�7@���m p�8����6��++�X���c}es�<{�Mj�F�
08�\]mw��t��)t��4�\s���������	wd֪,i�@�d`?M
�Dl��Qe�t��Co���ә��MK��1z�p���z��z��-�\���Y�~��]�GFHx�3�'��O���*��6O
/櫓K����x�F�<+XڴX�KwJ�U�Ԧ�AK޻��cbU�� (p����m3� ��v?��Y��p|_X1ma�����)W:<�g���[L�@��%4ܔ�8��]�c�,����$�`&��a$��"�!ߔ��9&��&I���r��pOpa�����$3�݅�h�;��z<����;��Ӽ�d ���y�1HآA��Z~;Z*u�����M3L�U�CVڤ�H>��m
��ڳ�t9��~�w�2�N3�8��=��T&j�W�$�pp������h��BS�@���{�V0ײַf�M�2AhbW�փ���$������T���J�z��m2�V�ڱ����8��U+(�R���ʢڤY7VO�M;=Wh@eU���w�_>JQ8g��[�(��c�����xU�}�*P���]��wE�f��B�=L���I
[�X�)u}��EBH��O�s�N��;Wa���n��
ce�o�nn��)d-����WfoG\4�-������1����Ad��	�ή��N� ɞ�VNW1N�Nvb ���TH���g����-5��=�]��Wϝ�`�q��qU]�<�Q����&������=3���X�	2L�r��tS_k�bNժ�ww�s�,�P95����@�r���o�����#�K��E��X^6���-Ċ�?'�P�㜙�zZ"-̆Hqc�^-�=?�a&b1l�����ӂ}�I:&kᩳ�t��sM/Lt�u�&ƨT��8��Wx�䀾�R!q
�s��&�"��ژㄙ��M�3��_����k�oA���Kq("4�q�����hM�!�����.�u�;'T���7�I#E?�����@��24��?Ueo>')�7,Q�*y�eC���%�����4��S�W��Ʈ���������qYW��mF�4&����RQ�۶�Z�tK)17s^���E���P�Q@�5�R��~�`��"-&b@�Q{µ�����蛙Y*�z���َ�xB��k#0Q��M�z��Rܨ�	;:�u�W
nXBe���оT��^�ݳ�����2�D������a� �p�i7��*�:���A�/�.�M8ַ�Ƚ�W�Өi.�����;0�z��'FC�A�D{���Vw۞�Z�-s'��NP݂��i;�C�h��td��8�Tz)V �^�)P˯�u8��AAe<��H@5kT���>�i?����Ix��B���	R�����[ľ��M%�������-�BII�^�����$:���0��w��i�ZOu�n�^$h����)�s��0U��f�"Zd�٬���{^@�CO_�p�o��g6Ḕ)�Y����QN0K�����3����8���j����uiJ�T^����\�L������J�SW���V�ʈ_Ax������wqG$�#���wIl��N�*W*_���dD���,f�(,�9��9��$}lD1Mն��ҷ(ݘ����<'���9I��~sq	?����b,�َ�hr����o�B���_�A�� ����"����˘�:e��Y$8�a�.��� z,]E���EW$b%z�Ɲ[��^��lj��h��襃�f7n�yJH��|zW@G�I�'����+y������������+m���2X��O.�b&Ub�q�y���f�E�Y.+�g�s�d��%��	�s�jf�"��{�g�|.�(.�k 9�@^_�?��SW,)���{��� X��ͳM���MU@ߖ-�Ɉ��'�-�?�2y������L�&�Uc_�Ѩ�'P�&��u/[	��2�29�G��~�6u�{� <)&]3H�/��64���C8��f	�����<C&p�Km���ܭ���w����S	$8�N�����Z/k��U�I��>�����{ �o�k�&�Fn�Z��F��&�Fh5/���{���5j������>�
y҂�����UJ6�+���@k��[0|�'bȎ{J��p"�zJ~���J�F\�����ﳤ������ ��'��vG�(�
�q:��2k�����*IBk�6��t4���_��q�̦���xC�W«l�K_(1L+�^��-\�p@��t�/q�lX�������KI��$ɢ��\�kz%��f��gXH�}Vv��gbI%,%�	נ�"�%�0r�U���n�����V�m��Z�9@s�:�1�[c�FOG-���������oQ�3��+$�W��5��q߱F�Şx�I}�`�f}�=���پj|���9*�A	�ؚ��Rf!$�KQ�x��<�eM��,�a� ޳y��8�^|v[�Ĝ��p���d����'�R�/����Mג����KO�R���_&t@^X��g��4�n��e4�,�?�"��t�_����g��tlDo �-~��J�A�G�p�dt�F$�t�z2� V��x@w/u�gA4����U�4H�����+�#��"��u]�3P��+�(����lKm*��spmAE,��\����6W��(Wc�M?+7�������� �}c�<�xg������MM �l��@_OP=�C� ���`P��"3�z���������=�����|!���`;p���1j�m܀P���Jn�dM��m6���M���C��Q�{���婃ļ�n�]6X�=b1�H�g��}��1͈���V ��|��}�]k쑞��א%���"�"�����#�˃q�]l"��/�۠.�,27R�M�{x���O�=��qU��mDF��e�F�77��<!�W���ț�8Pm)�4t_D�qy����̰g�͞Ӟ������o�?VT�/�:��b��C�亘�dt��x��9�>;�z��J���=W�p���=(B���[�Ő����r�%���L�G��鞎0R��3��1�#����5�쿸��F���� *��R�辷tV�dgK����5Jl������礷O��m�0l��y-V�:�x���wQ�\P>"L2��gN@y4�Ǿ�D�K��ʩW�Ss^T�35O$�2��+7�i`��w�~yS_���L�e�C��d��-&fmn·"`����dlv�P
Q��ú������-�ȿ��9��c���I���	��H�ںr�Y�J���ʡk��P�8F5�z"��βY��Ҙ�<��z����d�s߹�0Ʀ�tR�:�nƲ��vh�i�@&�W�)T 2ƭ��ǌl���n�MSCiD�	�������gli����e@B�ϩ�����+�dրc	ȴJa�P��Z�{�<".R���x���Zd5gKif��o&����15"������4�3�N|�|d,;���o�G�t4���j� ]�uI8��
$؂|�S	!�(,aw�W���p�7�0I�y���ɉQ�R��#��$� ��*�Òu���&0VZ����#�>�94u��4�l���>�
0$bxU�}³��!�j͊�Pk%�u��]U�nx�Ϣ���b:���RX�C���5���Ek��%�;A�T�����|.��[�)��Xh}S�e�+r�r���I���lv�~�Ug)5>�|��kȱ$E��F"��D1O�ϋjd���N1>���#�'RP�D]o��{�MB�9�跋c|��e��5G��W�e�s��5Aǘ�ڽy/*�؉�h�d\���e�n�*颋7j&�6� ?9���Cu��Ԕ�Wv���A3��ILS�m��-?�v
Dq�Q���L�P^x��H��L}���)3��mY������ur�����%^����W%j��P�cb;����|�܋�t���מ�� ����7��D�x�v�EzT��Y���a8�� Sa?%��#��%g���Z(}�;���ء��T՟�F�;�~��(("fBZ�����.l�&�vӍ�rhի��?���7%�����8�@�B�2����Y$�FE��%Tk��ox���ƒR�SG�6җ�[�A\[���Z���8 ߶ ?)g�h�r	� '[��6�d�\�lX:�5��Cv�|�h��b��;-YuqJ�[�n���O5�<y�-.�I��7�X;�p����'���Wu�s��,��=(O�I�nq�a����~Kf���-p���C��鹮6@��r�v������@.�;<��։:�:æ�`�aT}v�WS[%���,6R�#�����q0���Wo�HS���KԀ�:�ֵdތ��A���~�b����K�5*���ǉ=��9b��Yo`�Yn�4
w��&�.*'C��;<]�a�jM�!��=w��|-����{_�pQ{�W��_��x�)W��cT� �V�Z1?��PQ�c��'<�#v�Ţ���+�$�,�q������-������N8�����f�+��\��&�}C#7<`�|��F�8�H�]�<��)�)�8v�qsG��Op��2�Y���Z�H5-ߞ�`]��"}�wy����C�}�pU�q`߫��*��1�#�p�tb��0�zҨu�::V���~iؗ]��F& ��с¹3>������a
�(��hF���F���+�;X��wh����A��
�*3������˵�!�m��^���?�� j���2\C@�H����e�7�mL�32��?���>-�1G%C��#����_P����%�TP�Nu=65GuL�r�6��o�V!��LPNT�C�ON��>F�m胮a�z�!�+Of|-�d��ri�|����%���>���u���L�߲��J�A�m���;G���/M�a��s0���p�-tIH�U��n=�b�C��iչ	ɚ���F��������00
2Xbi�ǘ��tNx"�������y�$��%货<���R@��'��e�J7�9ݧat�N\6�-L��Kw��̉���N
+[�zR�u�cl��d۞ a�_��zV(���Gm��pQ�b�|c�<;�l1��e��t�.=��~v�lp_�7�Pj,��a����h(�=��b���S�F�JCr����ʴ'�/Q{���T{�ZK$_ӌE&�/�N�i-��@xp�U���$����8��}_���#�~(������6��Y��TB��f�u���~daHc��L�?p���L4���y�ˮ�P��eQ����tX�q6=�a�ؾ	����j����� 2�����å�oj|�Hwe�vz�s/� wls2pr�y�D��v(ь�]̭Bl`�k���>���AmQP�Y���\�C����1�Z��Xp�泡JG5�Y�N��C~�+m���3�'4�� ��.`��f^�,h�2B�@�����P3���k�����D�^�GYNߟ@�7�eY����w=1�Hb��{Y���������K��5ըh��˚�jr������K��+�-��ρ��@��*��9�x���;�ǂ�x��=���Ն�Qe�\ N��{�,�
-�f+�����;c���n��hUN��-3(��`�y]<����Iߊ�]? w#�w�X��c�u�������
ͅ�:��h ��3�ynu�mZ:���GDCwF3��O׬[У��7�9ghý0��J�\=�]}�fOT�T���gl��b)9�x�@�\w$�fz�C��%�@��'Ts&)�T n�O#�auSz�72�Uశb��� ��WDc綣A�@L����#!����{U���$��A۩`��}#�5"�i��n�G�j�efK
~;�l�֢᥯�((�����U�8�oojB�ϒ��|H��ުļ���7р�MoƼ��	[��H"�����R[9r����i��xVcrU54�y���{ΑEf�����c�1��C<�k���lK����_0�h1O�O�xj4��k�u6�d���^`u|�@�EgzU�2$x�!ݝ.�y
^vi����m�}�
�<Ez8 
Ƥ��c���|jp預�ҽ�F7{x�=�H�`J�,��3M���U$�|�q�6������gs���,��*�~<|���ɝ�~�A��T��
?>m�p��J����4��Ա]f��]k�H�B����"�୨w�Lu���CX�׻%z���$X����t?k�+�����rg�ѻU:q��{mL���r�o�Z��~�[���=:����#DL�Ď�r-ݔY�`����#ጤ��ّm�3�EaѠ�"�7���E9�G�&vd��������O}~�a@ŏ�Oʀ3�:`�c�;��_<��eE��]� `=�ƽ>HŜ��P��;�S��q!��vsLX�/V'�*H+N�m�p��੾9b�	��,�[&�h�ڊ�z�AZ���v��ycp=ۢMh�Jj�x�yS�'(��LEu��_I��mA�����Ɏ31�J`���Wv���gQm�0�V(wP��g��R��͛?�4��C������V���;J>Rh�-`� �۰L�)Q�o��|(�
�� �����%}wP��I�-����� B�q��x 
Ȕ�뫊�}BWB���O�U�N)ݻW���;�
�uYoԌ��MX����d=��I=�W�],\m���3��y�1��e�$&d�	lh��H�!���ʾ�Y �1�I�vd�^O���ײ����]j�?��:�
���!���D%���*S���>3[]l��^���\U�&�]z�.=����#��	��+r��Sl:���N�>'�`&ն����Ⱦ@�?�r���|�A�s 9#J����r���(������W����P�,�Y�&Zo��s�q�O^Z�=�7&�)���ә�Jwޖ�Xk�>��uszt��&3�b��8X;�W�z��!��sۂ<�L;��G�2��M�C��J��i������%Dq��>���뻜�oMM ��fN�l�Ԅ'�z���'�ڶ�}?��'�|��4鍂U��'V�,%9y?�#���gD��).T4{j�����ԥ�)͎J�H�~�av��F9��ӽ Rޙ����`�AՈ����sk䥠5�(�Os������~�,`�`��-�B��^iE�w���P����$�V�z&R��[k�B��#=�ֵ���zT��?����e��]��nB����8nT.b��^|ݜx.c�nZя_(�Th$�B�w ��i�|�*Tv��[AI�.͢�����5nW׵8i��z�K@�;p��*H�C�sDHH8�i�l۫2����'JSVP�������C�.zȹi��NǋT��z�\�^3O�P���uŠ�����A2������MN,�����V�K��<�3�x��x�]ߺ(�3Q�[Lzx��%[����b(��-I��������.Ȓ�e�ښΩS��.ݪugW|^�jݿ��Ѱ�!ηR���o"��̬�
V^��BC\l�p@*���㸁71Y��`���0�&�y�Ƽ��R�qƅ��WV@�Q~CJ�ny�x �U���k���\JYNgW�?Vu_58��Û�Y�[w~S�$��5�3�hl�]���_�d݅����5-r9/�����Ul1�4bv���h��e]{�\0�'ؘk9�*
~��G,�
�_��g_��T�`��|1	�m����I ��{��3�� *��fey�$(pd�g��.He� g��EN�%�r��/b�zLΉ[����v��.�՛Ͼ��8Ǧo,Hb��z�dF�VZ���<+�L��p����:�.�̗N!�GX����~�bs�����$y�fA�EԂm.���|���B�"m�s�7���{�#|��f.�4r"�@��_ٟ��@��)4FM{҃! %[J� �[��~NU�x��z���5��s�l�yU�?�����U$(%'=��&H	s/�X��p����G����]��G�<g%]���/��Z4����'��&�t	:]��]a<0��:������g��C�(��iA	��N�����o8Z�C�����n���{ި�ƊǓ]Y�G6[�(\��SXAhӿd5����Ȕ���� ;��s�t`ho@N�����Zg����9	��N���ۑ�Z3����y0��H�.�u{+'����JĞ��sM��L�W�h
��5�8����҉�ӆ��l؈C��,���"�J���+�#����_mޏ�?r��	0�0`&��J���N܋\��������l5i��?��u�˜+:���P(���q���2o�e�nVGIF�*6k�@8���u�_kiq=E¶�IC!�2¯F�K�B�L/�M�1�8�t|Pm1&/u3bXV�~�0`K����(����#d\�k^%f�LX�A�}Z��
I)�*�&ٙ%u �Yt��%��������c�벽�xw_�ĵtc�ߜ� - q��i*Q��=��wi�ۗn�9�I�n��J���K}���f��½�B{��@ɫ {�*���\M���U�f��QKU�zxZ*��J��=�Va�V5���8�%y�dĠ6Z��0w�h�e���F�!ROj������	��yJ��+�R�c_���^\�/g#��r��cr>�,[&e�&�t;�N��5-g8^�lH�㹱��N��Ai�ct��t�?��3�8q�$-����/yT�A�ZG��+�S���*F9S��ΈF��� �<����(�ѫ�a.��%����m�O^,���9�76[<(���MC�غ�������8�c�����ۿ���������p!���u�PA����j��Y�pAB3�C �J����-���Uu��j!5��`?�ߩf��jD/�?C��|�no7�M��u6hX�Q�~�����UT�{o��ć򃟦�r�V6�<]f5�H�jg�� �\�1�@�$�� �9����]�R��������Lo"2���v�+&ˇ��]�%�"�5|/i�.�b7֟{����^"O��f��e���@D�B6e��7��<%�;�(Nzȟ�9�M�8��Dl7����S�P牵ѥ<�C��������VX��ib/��h5��h?*������tJ��-_�~����0�������p+�=��������U��Ti��]��o��˓���?R;<3� bŧ�ъ���p����1�W;* .zR��x>�d�3���$��c���7 �$�2��*��K0p�6y���:�5��Ce�Q�j�>��P�4�!�gR�Qy�1����K~�ʭ)�S���Tϖ�����6?�pL�7ٮP`;�<��S�i�P����d"�$-�^�nҐ�`9"��h���Թ�Q���>
[����-%���?����M�I艈LNϺ�����n�PKkЉM��5�z�D��A�Y_���������֢����h����ަc��>�nJ���zpL���&�1����)2�ѻK7ʼ�}nv�tSG5����je�R��i���t��@�SIT�HS��q�ք��85�T��ZN!s�M"�5��H��۪Zh��g��f"�o�F���x
"R����4&L��R�|�uɝڏ oG>t8����Ց a^BI�Pd
(��|B��!�fO�_�&��u 7�I�������M[��V�k#e�$�Z։�ػ������ލ;0�o����#v?^�=�uN�4���$.�>�O�0���U���7jS!��6��^�k)���o���ru��&J��fc��{�X�"���������k�	;Ex��'����� ����M)V��h��Ʊ��ur�9�io����*v6HUk��>Ĩ��ɱ�})���Q�\�ISN���>u��y%>% #�#�P�go��՘��b9�Fɋ��T�ݹ��[�re
4��9И����}>�*�4~�����$���qe=s�*�7�7�[t6�u?���G�<�X�WzԻ!�����L�Nm�5?*a�Du��yx��\����L�L���-p�G�O�����U��U�.�^�����&~j�ָ��ԩ���� ��\�ע�� 9��;	g�ȧsx���E������_#<� ���%���Z �� �Z�(�;�/�zuN�ׁ�%㋞?~�n�(&uZ�s���lFfzĜ��yկ���B�;�1�&78����d�BT��LJY"*�Fɔ�%X@�so|C�#*�Ɩ��S�d~қ��[QL�\_3�du��? cc�?-� hP	 �}[_�h&8��l\*�5%�7v�}3h��΍fZ�����YyT��	����g5(q��1�m���M��.��t]����'DF����s�}��[�=,)���r�ca��������T�1����3�������^�vJ�v��������.�LQ�*A:����*E��eG�v7��[)o}��z�'���WpAq4�w��U�HWna�_UԄ'w�Z>2ސf��ů���Ib=�/�O8�*�h���s�Eb�+So��~n���w!d��2E�*�b���<�ݗ�nn	��b��wF�/|0ɃYc^&Q�P���ڄg�_)[(XZ#�r���h?�Q�Q^�A�+�y#��|����+t_s,ܪ��z}�ى�m���-[8���$�+7���u�}�Rd<�d ��F�F(8e�\]D��V�)�K
���)sK�n��t�6��ky��L{,�"�`a�ے�π�{!��Vw�C�6���.�uj��/0��.��1g�p����\�z�%��W����H~�f$]'F�_�ձ���c��5{�9��
Ѻ�-;����F.-�+�/dX�U�wl�0�6�"A�4���I���4�b���%��m������t
���2��a�L.�G�;>3m�|�2�s�?c#>1��G��H���i�j�_T	�<Z�#vT�`�uA��G�W�L������s�s�Y!*�e�Pe"T����S���.e �qߢ����~�{!Y� f��7���rmġ�Vx���ǮQZ��8Y�߶T����q�%��-��B�Mn����՚]��m���\-x��ِ��r�b��C��[�=����©��H���6'�u-�09rb���ǜlwt�&+&��#���}�P�R����~#�@�g)�g�,J;,ż�*�ax�SN���-Pe��5�w�D��~NP�R{R[h�ya�c�d����*���w(F�1Gq3�p���f�cA��pH��|�t��$=��~z��p����T��Ce\a	�^�pI�l�B=���Y���-J�Y��b��^��8��/U���V|P{���$�tgE*n^��WYEi����D� �[첕�$e��΃��Õ�J�~�ď�����6��-×
�B�1a���]��~�^c��,�ì�����Ls,y�9��2�UP���eC���%�������B������j�)���2D{��@�h͖j��hw��Iv~���� {��2���}%�D����zAh��F�F�!5���9��T��U:Y2�S`�Ռ|S�1 �H��\/'�7A�G�SY���G�+�.6���q3s��4�#��[R�ۺ���<�6��@4�rភ�3�0��(�0D�v�q�N:@��e] o�e21�S1���1{]�w&����Qߠ�S�"�=���h٧g������1D�K͞_���)��e�N�K�.J�9h�x�W���xт���R��u���Le���N3Kί���U�jdp�C?��\�o�҃oN?u�3,z�`�@|z��*�I�ح�el� V��?+��	u���@�Q�͉�\:k��l��;7��}{:uSb�:�	ZG�haF7VO[CeЧ��gLZG�i���\�+�}� �Oؑ�T�)��댶����)����D\���jn��bP�)wҶ���X3�)t"n� ]��f�z*�?CY����uQ��x��HO�8�SvK������A��sU7q��l���#�d��[5&�ǢH�Âj^�K����B����_�I�����l�c8�n�j�ϖxF|̱�¿��@ޕ�;Z���żyz	���H&���*��R_���b!9i��UV�(�58lz����~�ɾ����c5�y�G�&k��lO�`V��{�0�O�|Ex�7���:kX���h����O�|� _E�Z�6Mx 3�2�y
�~i�����谳d�E�\�
�Y�g������6~��qM�A'7���%�d�=,0V�My_;z$�״qB���J�b���,:�vт�C�8A��n�0�[KK�?��&G�X�8ތ���N�BӇ�T�Y�wF�-%$<\��oH ��o��b�S��g5�[�)\+yR���(h �e3?��h\�	��[fN��4xF�,��l(�5q*`vz�mh��S�2���ߡYE��+!ã��/5t�O��V9]*���܎<�@���k&�'�P8�'�s���Ą=��%�>Ra\�ǠN�5�]п��8���4�R&Ǯr�B�*v�zZנ1����#.uԗ�v�X:����vI��1՘v���[������/��8�У};q ���'�PH#f�2��Pd	���\��I��N�b��c��X*��J����h[b���o0��n��Vwm���l*�M7��i<-��:&��w���aw���|�����>/��QK�<��ބ�;�)'\h���;��*�?i�~Q������#Fzעp�<+���,��c���å��}�^	%8[[�٤#0+Y`��WZ}nk<�OL�F�.�8�{�]�N�ʢP�)b90��se�����׷�����n��`-�Ȓ��G�����#C]6�@(�A�Y�{������1���p�����z�1��
�L�k��~9o�]�*�F��!��f_��w��Lf���
��-�y��%Fz�+��lX�/�w8m��N�A�{U��i0P6������ma�ۮq�`��3����2,JБdO�e�\mo
2��P?��,>�<G������<�]�_ �W����T �zuC�G��L��F����?��!v�����T�S�+��z���=9x�1�UJ�!��fL<}�4��r9G���T]��E��yD�V
���{߂����=7��������M�lj؋�����@�-D�i�%�b�>�(bY�Ch�Չ�ʚ�F�F��Q�˯��0���b9��h�jt���\w�o!9�I�e���F�w��rn@p������J��	@�aD�$N,�~-��]wb���,$�#�[T���E,�c<ۓd��17�V�(� �G=�
p!�=2�c�3��<��5p4tRK8=��~F�p/��� �l���aէ�ʼȺ�8==g[�R%������9�X0xʄ��/!`�ܢ��{d�q$/F~E�hO��g�6`i�8-�-J�`�e�a�,$�A������M�ٕj4�~����C��_886a�7����B�D��EE����~4\�c�?�_��g�ؘ�>y�X$�~��P[�/!��ܪ�Q�A�Z�X��؎�,�l��jh?�� �2�B,y񼥴��jL�Qw5{UvJ�zԥ� G��2@�g�I�[D�Q��Faތ^���������_\Ѡ|�!��Y~�F,�$����1�n��p��(a惬AG�YeM��W`+�_1��0�3�l4�a�	�˧�v��6�@�q �j�3�B"���b�|��Dsc�4N�W�@^ʒe)s�ұ�81R�Κ��y{)��r-Ҷ8���uj��/�,�      Ĵ���	��Z�ZvI�*N���3��H�ݴ���qe"�T�A (��џ�:0LՐC� ��̞~_�����8�Mf�i�07M���@qe
H�>`�0��ab��h�(�~#<y%+�"�\7�\GTxV�QM?J�d��?*��b�P�)��%N���J�y��o�*��'e8X���Su1 �Rs"�0hbt��M�6~���i����Oʜ�2���$3�2b��Uz���8|_��c��5���DxR	�J�'�*}�UD����:Jr	�g���%����ቑ^ �'�"�X��ݭ2�c�$�����'��!ExB�D�'�(E�&⎸9L�[fM"-:iR�G<2j
#<S��>��O�8��ɢ��O?Y�ܽ�T�J��Z�OVT�{��V�����cP�G�l�o���M��b%$�#<	����@D'�<W*�G�$,�P��>I�4=)��Hb8iXH�=e��8��oͬ#}�ݖ'��ExRAM��B�V��ՏE�e���DΌPov]��:�z�"<!���O�L1�Ζ;�<݊F&��n� �Iw�Č�O6�	M<a���NZ2��"�Q�N`D=���D]?)��:1��OH�X-������]3^mb��@�~x��IB�?>�t6-u��'���^wv���	ؒ$86��-i�x��t��9}qO4AB��d����'u��R4*0M�
Y�� _���.q~"<���1��y�!�]���1�J�5r����ȓ'�E   @�?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       P   m	    �  +  B$  �+  2  ]8  �>  �D  <K  �Q  �W  !^  bd  �j  �p  ,w  �}   `� u�	����Zv)C�'ll\�0"Oz+�⟈mښa�	"�L�D*�`��2	����%GV,#��Ù~d�(�C�|,nU*�ま~�@��	��`��z�`y��Mօj��7<��j$,dߴ�	2�M,\p�k4R��x�QB�u�,f���#%D柞��\�̤����{���
q%R�\	PȀ�#� 4It@�Io���2b�Z�g���I۴����?���?��58P��nټ Rf}���U)��H���?!c�i�.L�WW���	9?+�5�Sܟ����~Nd=�兖�u-�a:��ٚp;���	#��X�'jH@�&��Ԃ������^�!���Ll�xA�D4�ԍ���/D��y�F�D5��c�*Q(�k�O�Y��.�<3��%ZU����£�x��0�~��	�;�,`&�:	������?��?����?����?�����O���A�gI4ɴ-�C�K�+@2�'k��'W�S��C�4t؛��j���l�ş0����M9B�`_%o����dJD�'��gI�3@L$z��Ӂ9��H�tI�j��j��D"g:A�R@��M�5�i�V6��0ȭ;I(	�Х+dέB��A�R����L�#i�,�1P�i�V\����3��x$G
6���[ꆂ��M	�-n��Qm���MäM�O0���m6T��FC��Qm�X�ܱ��ii�6mZ������"e�\m2��ZI�l����8^�V�
0䞥^�֥�M�7�2-�Ai�EJ���j]��MK�iSr67Y�����\�Lm"EP�iZ�f�x1���M�zɌ�.X��`�(k��4l�`T����O�����s�S�p��C�i��SF�W�f�:�afD�>�~�Sև�0%K.,��i<�6�U�����?5�A+\; �i�F�Ο(�g��X��Ɓx��qG@N�<���+_V��r�%�'Y�>ԑwiFO�<���0<�p,���H� ��s�<� D��
�@��Ԩܣ���I�J�<A�"Րo�
m�F�P���)�`]G�<�P	"HH�s�n��bd(bmR\�'��鹍���SB�Ձ��S�H��M�!��ِlH���
�k��]R!#�$L�!�D�*�h�``	� Hid`�!A��Q�!�$=��Ҍ̽Z� )r�)X�J'!��? �rY࣎R�z`xb��j�"O�8��a\5� h7�˿dq�-�3�'�8;���Sf^\R#C��O�ZX��7�l���7�����/��U�-0֬.g�4���{��DX%��V���b↪w���ȓ�.����9����*��d ��ȓymL��o�k�P*B�UA�6����z�i#��}Y���3��:Yؔ'���	�N��ْ���|$.���D�[�д��g`���E�9��Mт���g@4,��2/~��}9ʰZ�Ʌ
�@k2�(D����λ��p���U�2d�v�*D��1���@鞍 �lT(5�	���'<O����9O��3~Ys%
(��y���1!`�M��I?m���)Qr�Q�|����:$`����LN�� ���	<�0� �ኾ]�h�T!Ê �5
�;��\=+LZ��I�Vh���O����O�8bo����p�@oF3!妑R�,�<i�����(����-�}�����eb"0��'����P�
�E�"e��,���F�^��]�i@�[ڟ����y�hN'j
Ⱥ���r����*���$U�W�n��{��	βCZ8��eJ*p���a`b+�	�n�@q�����f�:c'o�K�l�ht*����n�ܕ���<'?��|�p��^��1���H){��.Qy�	���	�v��{r��>q=��'�A�x�?A���;J@&����a$uBs(C�r���b��H�3�1�������jx������R��>o-��FS��0huH�:7ʚ���?&2dpF)��~ �u��KŴzu���ȓF~���f��y�Ԣ3k��@�ȓ䴐U��,`�0���` &���Ɠ}�UA�	ڂr���BH#@v4U��/Y�<	�]��(Pg2�Vl3�.?��AA#Gy<I�H��F�Q�[L��8)P�fG�����F�P�� O�e�&�C��Г���X�Iӟ���Kyʟ1O,�`�
��AC��Yp%�_�(�Ȁ6D��#!�	�p�j)[�*ݜ,�2bh6���]�	ly�M�yґ? ��\�a��3���|�L�[B�)O,�r��)� "}��ßP�6ز�j��
k���R�'��0ێ���f+b�#��j|�@Q$�s]axb���?q�y��
!���
]K��FǾ�y��yLL,hIX��QZ%#����?6�'T����O(4�"�����R�h��d�*z��̧ ~����c^b�qSaO$"%x��ȓ*Zb���DY<�@�1�%�|�|�ȓ/.RIO%7��v�	;D�섅ȓ �ċ�IB�� HSbI߳LE����
�6@z�)��JT*�c������ȓΈ��ٖ[��]�sn��z�r8��0cn"<E��ە3@�VR�PY�@���ofr���4eaɛQ��u;'ȟ�\lq��n��t1ehK �b�
�%Bxḟ�Q�j0�b���<�f���x�ά�ȓ�r���o��1������#E�<e�ȓS��3�D� >�=�c�"c���'�~c����6t�nz5�J�5�%��c�4H"O-1R����D�dP`�ȓU��3���,2���V�G��'�ZX;���e����&�$:��-�ȓY��y��O�]��T{FCW)l�؁����/&�I��eU�O�5��o�{bBC�I5�$�CUu=�}{���.��C䉃� zt�:�Up����C�8HVڸ��iα�����b5۪C䉺!
�� �S�:��v�ƔGm�C�<���y3FY$>�"���.�*A��=����A�O��ăҴ3���Ц�X�����'�v�b���Za���`�d��'Tz�ֈ:`xF(�p�C	[���i�'Qص��ȰIs.$�CO�1Q�`� �',>���>X�
��IY���M�	�'�8�'�!o.<���K0������Q�l�Ex�����]
^���Z�G���5+V'W5DB䉒
�]'�F�qޚ-��ET/iZB�I� Qx�%��)����=c�C䉸&'����LԐM.�S搼S��B�ɪ_�l`c��T�x�j]HOJz�C�	8;�B`��A��h�4SB�U�
��˓R\��ɊJr��%�@� �I�rc�A�C�	�Ui�	�#��KV�Mv逻|N�C�	<],T��'�)GrRQ�B˹<�C�	"oT�(�u�u/ ���ǉ�*�C䉊d\�
3�]� $�;�#T�',��ċ8X����W��kf��%G�h�{�	�!����0-��2��a$���$�!�̸j�rI��L9(�藁Ԥ5�!��D'���@E�ƅ��c�i�7A�!�D��1���e��qڍ�q�$�!����@`��# '�!jxb3��W�ў,�G�/�'�B=��"J�8?��q.X8hD�1�ȓR��܂3 YÜ��7Ű#H(�ȓ[�XA�+7}6���'��+��<�ȓ}=�y31O�H�(%qA���9�ȓtx*��"(�H$D:�P��ȓ���Z�*I=gJ&��0����r]�I
Ql#<E���J�K�(�����xJ��Ӯ��D�!�d�??j�dpH��O�����λ`i!�d��^�Dm���~��T��O�zG!�$֭XM��C�N��*�H�+q�78!��#�4��υ�x!*�ND�C}!����- ���}o��Z���剸8�
��D�	�n	�d�Z�IP�]���J�!�� dQ1��`^2Hw�� ���"O��Rq�����d�	
#�9#�"O4�Дc���pxsC�|�"O4��%
�r�X%!�h���'�x�S�'\ფ�!D�u:3��(��В�'�vk�J�u� �S�"ؗ)pB	
�'�����1,F``yå��u��P�'�N�I�`G=U�- ���_B�)H	�'�h�Gꔭ:��h{�nH.\>��	�'�Hm��Gp춵��KG8h�����-$Q?���m�L[.җ.J�jv4�wG1D�tQ�3"����&��,��r�-D�P�2�V��4Z ���[^�ia*9D���F�D8j�ހň�Ғ�cG3D��	"���P���q�O�=��U��
1D�����r,u�R�Om�ʭ�-�O{4�Gx�����!k�$1"ɠ$ɼ����Z@�B�	1L�\��o�l�r��S�ֱj�B�	+1�Y"&K�J�B �"b���C�	�u�����lX�!�p�p@>3��C䉌O�H�ie��1-E6 (2��x�C�d?F���/�^������`�?���~�
m*�$�ĝX �r��B�	�|�����jU4-�a��)ZB�ɇ��]µE�j�����i�7�C�|�����"�;k��M��g��sA�B䉢)k�(�F

@O8��d �L���ߢz��F�bÌ�XUb��k߬a <!�2Y6��e.ǫ2s�1!��שm!�Dұy�:X��G��IsT��~Z!�ڦq�(: dEa2mQի�x!�dH�a��T'ՌK^l��2K٨C]!���;@=8�hR��h�sJ�=cHў�B�/�'ml֙3r(R1:��&僟g< ؄ȓ�t��b��N�L�[L�0{���1��`�V�N
(�̓Mp��ȓ@v�M��a�>}��0��� $�I��U�d�']"D��YU��=)x���EJ�8';}|J���
D�E�I2"<E�d�IG�6ĉ��O�Q� �{a�M-�!������Z��x�v%��k��b$!�O�S��y�cC�9�� ���ny!���-0���k�Y�b봘�#L�I�!�DKc�{��Ҙ��Th
�/o!���1�qc�Ɍb���hD#[I�I6X�����[@��5G�	4�D�AD"R�!���:�q���4 �L2S���Z�!��Y1�Rm ֪��F�R�#%f�@�!��#+\�u;r	��Z�� S�x!�ĕ�V� %�,�i@�8���-xf�}b	�~��w��d�D���*A��y2�L����A��ȃ� $	�A��y�J��hT���P�9Ǽ1���8�y2��p���[=/N:l�0����yrnɷp�)҂�V��`�͝�yr�� �ءg�G�}��x����hOV�����<�[��[�x1��K'vm6B�!f����\��qlWf�0B�n\Ѕ��-i�Ҁ�4�@*�C�I Z�����$&��Q&�Ճp�C�I���L��aY�K~tzWꓹ�xC�B:`MA�F�b֎	"pg�2�J��	nK�"~�%��n�(�bW����\{� ]��yR�H�4�V3V� �[SB�&�y
� ��0��E�'?EC��A�[
x�8"O���w� P:��鐫�T�;�"O ��p��N,`9R�ĩlӀ�!"O�	���ɝ^�h��տ(0F�[��k�O>�O5�t�Q-b�j�k�c�y.x��p"O~}Ӗ� +F֬�`�a�E�58�"O�#���"D���p��>y�X��"Oްp��� �ju�$�;g:@�"O4a�&v�*� @�0d��bW�'���'�He�cnG �Y��F����':n�j��
 " ����B�f���'��#��UI?@8AP�%8^I��'��P�%����C���� ���'��ui� �`��5��ꗖ~~���'��h� �B�ʩ��!�޽q��$�x�Q?�(e���H�=8��L]ỷA:D�<R��xZn���<H��Y��%D����JhBL�'�[�ppu�R�?D�x�b2���\82t���
#D�t�S-�t	m�s(��$oPl�4 D������*I7�,i��F������OBQi��)�'/rL�xf%%}P��fшNh�Y�'��ή(~������N��)	�'Oj�X�%�,J��cu�N^�Q��'�<|�WoۡG���t�����'GX}��	s�H�b���ug�ղ
�'۸!a�	2tp0�)y���[*O�2'�'�|`8⎑�{�օK%������
�'[rK���%'J�Cu�.H� 2�'4���f�O�>	��ۤRg(tZ�'�m�b�-:	n�u΄Pʐ�8�'^hD1��@O�n���e3<]��x	�C�T8�o��{�EU�w�~�@Ê�p?��ȓF���a[�h&J@+5�X2T[0�ȓK�L���!I�k��	AjP/2Ħ �ȓ,�1ɔc�D�j�rf.AVц���Dȧ��3>���A蜫^F"�������qo�5�&�#��)h�B�F{�%^������	@I9p*I�6�̣O����"O����V3k��!���P�H�D"O�%8�S,#2�)AF�
R���"Ov��@�^h��Y+��mpU"Ovйf�޴���"���+�"O^шuCF}=�e t��1|��{��'ȚY*���Ӎr2]	� ���pE�M�:C@��ȓV�pQ��W>�|!ۆ@֘\�vX�ȓ<�(}`.�E��}#E=�$��m�����	Ղ'�4�@�)nd��\���+��3�|H�#�'v�H��DL����Wp�n�{4E��S�M�'�>,@�R�$�Ѕ��5~� c���<I�ȓ0����@��+,Y{��K;\���ȓ1��T��Ϩ=&`�������@��"������8F����ȓ$J�(o�O�䉸�N�Ga\����&8���	�RA$�����%D.\B2H�B�\�PJb��B2ŉ	�H�B�ɟ(�N`����c��b�<y��C䉨+*Pkw�B�}�ڴQf�	!w��C�I��L��5H���ݻ�C�I/VW�(�5�gtN� �o]�CϮ�=A!d
j�Oy���4A�Mx�!��)l��
�'d��QM�E&��
#0>n���'�%+�ǅ�u�Rt���E�"�B����� ~@"E�"Q����HX�b8��$"O�d3b��AΉca'�E�P��"O��aE�D�^e�y�7�ޭX��-jt�'�I���9Q���:A�\*:2Z��a�%`���ȓ����Fn]�7����FhK�%��ȓvrĠ$O�0���I�'�� n��ȓS�>����j��P�w�
,�Z���m">�������(�`Ci�ft�ȓN.�=�2��p2H��`&�����'�>4��tLlm��  �{��:A��iH)�ȓq��8� @ݢv������/�45����h� �y�^(��h�
K� =�ȓ*�b�1'���(�r��G����ȓ
x��3#�j�l�����Z��Շ�	�%Zj�	�� @��R!:Q0���N��C��7P�(x(a��7���NW�f&�C�	��Y�o$�P�U�����C��.㶠�G(̄\㎰�D��'HntC�	 ���#���P�3jx5��"O� ��m' �T�*�GĞ_����!Uw��~"d��&E��O�m�,@��Α\�<A��V�q���y�͏�����)�X�<q��q�E�Wn�	r�0����y�<��FH��ر�0���h6 y�<ivʛ-ES�����m:�`��GMx�<A�@�9g��@╭J�@�cfbɟ`��?�S�O�0,��O�#n^���f<Ɛ"""O��)��`�����ҸUJ�E��"O�x2TK�u�j��@J��N���F"OT��6�Օ|8�0�B(Ct�H��0"O�1H@���o�A��dʱ*�L�3�O았��E��"�ʁ�,*U(5Y��O��'���h�'��ig�!ȗaށwEh5��ΟA�]I���*>��t:h�7I:î�|���kC�}K�oU�@���3D�'��l	���1X϶�# ��9�S30 �0��ņVn�!�墘�#>Q�t��w�'k����F��b�<uC�g ���'7a~�a�\��0�4Tp�K��>�UT�`�t퐉k� �N��Y	��)vj�<Qf �<Y������I4)A��ŉ�{�"�$�ƕc�h�	 -N�ˤ�O�X*��X5J�[�OP���$E��xX!�d,cO�\ќ'�d�bK��5)&�傂z7�?��v�H
�<� �_7�V1��	r��`��O��$3?%?��'7��
�-?kN䈗��Jrд	�'����I;>����� )y�&P���R�O<28p�)�T	0�(T)X��PQa�\�8��O���I�^Pa*�EV$*�C�cܤ��C�	^S�j�n��	� �Hү�7 ;�C�	s�l�Bፕ^�^�aa��<�|B�	�t����c�:�+���p#�C�I���!�W�6�Z|+�ƀ��C�9l<캦��e�� �5�ߘM_P�$��~riּq�@iS��E���"-)�y��C�yظ�K����F���yb�
,<`�Ā��5xİ��J�y�.S��H��(P�q�3jR��y�,�Z��6�Y.���^���=���A�dD�9��U��M'(dH��)�*e�!��!Ek��B#D� � �#�!�$Z|�a�'�U�v�h�s4�!�DJ`2�A�.��2�@�i`��x�!�$ȡ_X��B�J/=��t��)�!�$	2�\��0CV0%O"�yp(]�0F�O�X���)�4M�E�q�L�.&�0�j�mH��y"��7%D��ao�7L�������y"I�1�0�M��>)�丁1�y
� �u�E��"Ĩ`'	�V�L�R"O(���J;%����i @��TH�"O����͒�(��@�%G�"�6Z���O\�}��,aĕ:�,�
�P�
�O�ڌ��/=F���Y473Ʊ�W�T�K�مȓyt�� 6������C�R�ȓ[6�T�Bʊ##����E���!��f�Q��l�BĒ��K٘N-��ȓ^2�!IE��6l���b��L xJ���-+K���I�Q�^!{(�fu����fɿR!��[�0Ѕ��C��T�4����!���bHcW��'/|�<CUM��8m!�$^�$��<h���Ker�谋O�.7!��FYIR4�r��"{|����o�i5џ�%�h���|�`�)[�$�i)��E��_�'f C��)�6�0�4G�6� 
�,L7:�XK @>�RT�jҨ�AU�(Sl�>��F|"
���?��)ǁ��Aс%\?{.��gJ |3!��+*İ�*�0�B��oӻR��}b��<��iܩL4��cCK@�.1��cU�fyR�'�"�|��)?�>T*T��;�0��1���7�ax��	�v���c����6� @d �'G���o�_�	w1��0�S�ё >���Y zI��Q ��xb�'@�ܩO���<!C�A�"�vU�遗+LD��ϓ�����O�ȤO��ӥ�>᧐��NT�eka�^�"�)�Y�s�F��O  ���h��dǸ���Q&�syf�P��ƙ�1�>!1�>كʇf��D��9T�d���A�{��)���Լ�?a5o_��*y��?�R�i�6z} �Ӧ���d��l��t���=}�'$}"nڶ����M�$U�k�~���C2��8�"�syB�:��:�ȟdq)��ɠNK��P�kʂHB��Q*�l?1rmGm�T>牯/
 �%h���&����-p�jC����DF(}���D�#�H�`0�r��!w8XR�	ڵd��,X��'冰��Mެ-��9O��Q��O�!�����C����n,�K��'�����4a���c6G-n���&9��C�m�LrB
�!�b���()pC�As��*�	��9B\H��&��\C䉀]e���S��F�,d��A�v�@C�?&����&��ux'�5e��B�6��(n����j^l�&B�IK���qCA0u?	!���"B�?qBx������JW"�Dt�B�	�RI���Um��xrJ ��B�ɴjV�("/�;'���bJ� Z�B�	�_9T���W*W*�(;��Y��C�:r��f}�)� �'��A��D'D��jC�W��\4���C�@v��AG2D��j�_���M�7FT=y �$��/1D���A�<���t*׽�����2D�,� f֏p3�rb��Slp�&�2���lDj4���~�iĈ-1��P�LE�H��:��U6XϾ�+CK-,yn�y��\�UUp5#�m��<(��b�f˂S&e��X,l�nxj�D3�|�p�Q�a=��
�bE�w4&8�� ,���ץ�6~��⁆3�Xb�iW6K2�u�g	�FW�	���:��Lx� �T���l�K12t��f��x�ס���ZqaP�[�Q�|ņȓC-T�C�HF
��xr��)u����ȓY�`�a�(6�n�(��Ρ'm
%�ȓ���JD�Y�8�28p�,6,d�d�ȓY��f�
�(���5e5'��ȓ��������\}��/®X�.��ȓv��;T�D@��QrI��x�@�ȓQ�%�S[�����ǖ�nY�D��;�nܰ㨃!5�`Xy'-�	3�bQ��9J<�Qgټ#.
����VFB���{�	����2R$Bìʇa�<ц�eԜ8!c�&��9Fl؞E_��S�? �A%!F2�i�$]�
�x�"O�H�UD�\-�۱�Q�R�H�'Nt��֧A*K!x�A���k7�X��'81�ǝw�5p3�imB�#�'��
f�Z;Q���
+PNp"�'��UP��ɀC��<P��Z(<͘�'�0kċ�
|�Ny�F:X�����']>��c��JоQq���&q��'X�|JA�[
�f�q��� T�%h�'���Q@�9����,�,{^��
�'�ʰkU�ʇ^�V\D%��
Q4���'�0��%ߜP�AS�����
�'0X���׵9F�*7-�9���ȓ35*�q���:5"ՙE�U�|l���ȓbbޡ3��N{�T�cɍlc$��U����R��S+���܅(�8��ȓc$͘`��3g����&�B6n��ȓ�0hr�W<-q��0d��%Q�H�ȓs��Mӫ#�p 3��)-����51�4��t���b�B�v��ȓo(dt��$�7m��� +�F;܌�ȓ_��k#��:/̼-s�ǟS���ȓL�ީGFY	Lc7e�%��0Ft8)nVRc�5H�(�y�ȓu�~�HE�֐P>��PK�i֜��|�� a�r:����P"_�lX�ȓ�"UCV���H�d@���O�{��!��@��\�b��X�!�1�G�B���z�S'��@M��Q��0\ą��H��A`������䪍�'@N@�ȓ_�2���"���� Sڢ��ȓs��ҵKՌ N,s �]m����G����"KK.DR$M�Jꘄ�$78�0�Ì���a;u�ħ`�@��FePA�D�L�7 �)Sm͊��L�ȓ��M��R%� $sD�	5�ȓS�(��!��wd�� ���<J�8qvn�:�2X{s��GT!�dM:&�"���M�!��u����R!��i%�؛�"HE��д���!�Ė�&��y�$?��9�
�?�!�U	 ��|���C$�D̢�螾9I!��U�ĺT��:&�`X����%!��R
`��P탰6�����A.!�B�{��&/�")���J�C�`�!��V�Ǯ�s��E�
x��j�CH"�!�d��W�z�P1�عb�$���)�!�D�H�ʙ�aA�K�<kc��26�!�D�!��a
'f�wR�q�P�e�!�d�,>I>���!?4�zs`M�C�!�Dۜn��b�	Ó��T�! F�]g!�DwȢ�jt��A�`��C��� H!��m8�,J�'";�(���N�-!�D�M��%L�B�R0�ǮJ�!�ͭiL���&�!g�ܝ�Ë�p�!�ğ�4܌С�˘8�H���$�V�!��'N��ܺg�M��xP�L/!��4�^�˵%�K{`�("\�X�!�dC�@�Z��@���$^\8I�ҒHn!�d�ߐX�F_lk��bc/؁#W!�E� �B0 'H&
dT�
7��)\/!��yՀ*���Ko�����@B!<���=�u��N�1�|���J�7v�Zi�ȓX>� �����(w�0�̱6��ņ�S�? li����*F��9�  �W��-ˠ"OBظ�Mc�*Ze=�Rɀ"Op(2�`�<�{���7"�D�c"O���գݳLbPV�@&�T�;�"OPXzR!}Q��@�Ƕ_��@�"Oؤ�h�~]45a��mѤ��"OL�
V`�N��z�N��@v��6"O��[�b�2:��8�%���x��U"O��	� ]�T�8|+�@Ӧi�\U"O�5n6"�i�wN)�؁bu�:D�T��υ_ɼ5 �f]���4*�!8D���A	'J)r��cNܰ
Ze
��7D�l`-ק0��������"�`:D��K��4����E��Md�h�U�#D����KW�d�j�U�D�u�'D������q����Ņ�S�T���k&D��Q��˗&Z�|	2��$`h(w�/D��h$�M�l���&����X���!D����P��e�'f�	9#@��#>D���`dE�P��O.\Tll���y#�?9��Y�ԙU�$�Ku���y2&F</s����M��Z�.!2���y��@BNU+�[�R2��r���y��<-h��ĀPo�����K�yrf�#~.��犓r�Ji�rB��y�ǎ;�P�b�B<m#�9J�Kͺ�y�	Y�6������7O��r��y��J�C�Ȣ!�߈���nS3�yb�[-ࠡ�D���|H� ���y�e4:1N@w�C�Of �b @N�y�%'OD�e,�BӴ�pd��y�]�&�h�B
;*��Zuֱ�y2a^I���Ti�*0�9`���yR��-sf�q��*��٢�T9�yR� J",�Ӥ��~�Ρ �b\��y��Ñ<D �R�Y.��A£
�y"��`�}��)�&�Q2%W��y���8j��9 �R��b4Ȁ��/�y�.��l���A&4[����BM��y�SZ.ʴ�f�CF�����yBA��j>x���ą)G��M:3OT��y�)F�g�>���C��Ԡ�^2�yB吗s��r�"��	�@���(��y��%k*As3��(S􉁐�y�� I4�KD��~QpT�b��y��h��C�Q3R(��"f�y��Q� ���A_�.�<��%���y���+�����G��0��	�W�Տ�y�A�3t�.���M�:�r�Zgk��yR*[��z��L�1e���B�y�٨/ �y��eܱ&�fIJc��y2n܆h�Ջơ�����F�y�	U�*���S��Vg:��/��y��@d�Ƚ���Z��&�ظ�y2a�h�l8�%~7D�"�`ب�y��ֈ���2htx����y���tyNўY'�|S6��#�y��d����C�2��tR�&�/ld\9��,�<$�4A�2r��V��.E����m�r\�!
%:͒�*�.m�lA��g��i�I��L0Ka)�%~{B��ȓD�@-�c �.b�L�rQ#")@ńȓy�x�b�+m�,S���{��Y�ȓ;ώe���K�]o*���"��q��S�? 8� ��&4� �JKQ��;"O>��1��*�j !Ph�2h�l���"O��A�ٍ4�n��ֲ8�Z\�4"O�!��O���\8��K�Jb�]�"O\�چbWu@`X�ǣ�:]p'"OV��	 %V��XC!�.�4a""O��c���!�X�v [���q3"O��с�� ƈp�a�v�� �"O����ʉ46�K� Su+&"OX�s�gѝo�R��U-���X��"O�U�G��i���Xb* mŨ�b�"O�P(�"��L�#
��L̀�"OR��d	��ku�ZdQ�	L���"O ����Ő�h�����]�2��U"OrM�� uk��y�P]8�q�c"O�H�M�<y�p��!m�
S!\T1"O�)F�ݛXD��kКW
=R"OQ���(S��S�)I�nM0x�!"O�hK�[�&`�pVb��tC
��"O�,��$�?$p�{�"C���q+�"O<<����#��$��K�|��e"O�-��
 ��-�1��1�Ё'"O�b·_ƒh�����d�F	C5"O\X� �>�p��h_RB�CP"Oj]ca`�"b��=Y���R�49ˆ"OL$�2�L�?a�G,F�3x4��"O��wB��c(�S*�Pz ��v"O�T�X0y���3��8fv�!C"O�,�p����l� �hҰ+b��(p"O`��rc�-a|)c�G��G\A��"O�ݢ!��#*(�@"�����"O�u��(!�pu�&�4���"Oj��F �"B��,($�G�J��P"On`��hXy�Pb!�ņ(�R���"O�D�gH�I�}��F0e.��@�"Od=p� ���
��_�<�̻�"O�Pb
�+���B6#�2MBB"O.���(
2� �Yӂ_��qSU"O���D'T6p��`�W�=�"Oy1r�S {�bܘ:�b`�4D������:2���!�4U�pQC�%D�d�D�ӑ-&$�x��~^�Y�#D�(���A�F�w��.씹dk"D�l��%a��`���W7�t��-D��󦥂%A0���ǈ�ZwbUS�?D�0���
�	�j����j뀭	&�=D�0��#t�ޅԥĂ� d�"o:D�X�u�ص ����G�����$%D����ڙS*���BB5TiН�4h!D���u�G ��K1ϟ�����$D��&�� Ԧ��iҶ,��3M6D��o��g�@D���� �2D�T˕�H�,*T�8��\?.StX�dk1D� h��VF�T"�#�t�ivC.D��[e.�n��!�� U�/u^�s�-D�����B*v�N�;1�Rn=3`F6D���'�^�(ƶ��U��x�
a�0�'�I�cŰA��-a��D0����B6�OLx����1/&T�C�+MT�[r"Ox����C��b%��K}���"O��Y�_�o�N��@��'�fQ�"Ov��iΕ\A ��?3��tr"O�]Y�f����e�i�bQ!U"O�T�W�60���t+Z.+�̸8R"O���6�\�f�P�jB���i0%"O�  E0DNG��(,�I�!��V"OFlKGN��&��� åښ1��	""O����fD5W"����7rsʰ��"O�JT���S�P�u�Z�Sup1�b"O@��ŎH�N�J�P I�c\
`�"Ol�	G��:P4l���ٰeV�ՈV"O��3�H�X ��g(@���"O4���:B�����ѿ��4�Q"O�퓣	J: nm�+�; �Apb"O&�Q�Ӛ@:a�p�Q�)�#"Of�!�V�#F��2d&*��LH�"O� ��
4{�v\r��	mZi�T*O�] wA�X�6i0u�@/#>�H��'����Ⱦ*�8U �k��j5�`�
�'�=����a1<XAcWh��AA�'b�Ļ�#�����B��֘Y��'��]��(�[L�kwG[�	��I	�'�� ��H�c7�YpVGɽ<8�P
�'���K==�F!¡%9l]
�'!*8S�@�3v�f 9�̀=n�t3�'O~=x�E�#S�:U:���f���'�н��eڒ1�B�"VM�/=x�h�'�ܬ�%�͌��a$�77J���'V�L���;Vda��-�,�Z%��'�h.ƒsNR�ÇO�7�����'���H�z�(m(�B}����'�0�z���#k<=�'aB6@�Z4C�'�������L�j���c/4���'�l����"����SKQ�H���'�4��BE�Y=N����++h���'&Xص`������t� (��'YL�q�Kn�%9��W�e�����'E����	�X���ţ�'iҬ��'+>I2����R̝���]�`���'h"=q�Μ9��d�ǅHƤx�'�ę�� O�^%�5���͵2ߐX��'����C�_�'�,�B��)�����'�Q��ae�P�V��\��M��'s���ro��k@���V6B��j�'k�����$-#p�N.0��'|�h�#�	�.�(ӥȨ4�011�'�RQ�$һjH
5��4�����'�P���MG�;Ϝ����۷,���'�mk�Q�h��
�@� �@j�'��y�j
~D<U�sC�k�Z���'�q2%�șOU�����J�7V^I��'nE��͞[:�Y��H'$�:)��'	2|C ' ��m8�)Q�H~��'� t��ɔ\b��ScK���`�'��US��[#$^XP1⍛�QYb�9�' �Y�Y����e�?lr���'�H����5|~��o�1�����'�Txp�ӂg��-�E�-�x0�'��٩D��-"�H�� _� 	�'��;��M,c1B8
��J�T��,k	�'���y$璊J�飀n̙M'�d��'�\$���X���X����R1$���'0�A�N'EN$I'LבFd\!��'@�Y$��i�İ�Ug	�xuj���'� ���aMO����@��t�(���'�`��gI�D�����R]z� �'�x���1,��B6O��M�����'Ȅ���V;xZ�<6��37�%B�'Fja�o3?)R�Q!*'+�,s��� ������2sR1 �@Q�@E@��"O����&�aZ��w��%�2\�C"O9	DJ�a�n �tB�w��Mا"O�����I�4N]��O�uO�@;�"Or\�2���1Rl�`�K����"OtrS�ڂ�L	���U�*���H�"ON �V��sN��3�^�K�� �"O�%XdC�'u�X�Y��W�0\e��"O �[���-
T��
P�w��;g"Ỏ{s̀u���dg�:�,��P"O��`��7�<}��g��&V0��"Ojt�r��:�і�ڒ'- X��5D��{�/$ LH@V&�D��${��0D��m�H��l�/L&U\q�e"D�pi#��%���9��?!Xy! �!D��8'�б9>���CD�=Kft�!%D�|���B�kV�A�RX+�0D��!�i�>@��6���+���2!9D�����,^l|�)�eĉ}��H��&D��CN�BG&���N�����e#D����$T���iq3�"�$�C�i<D�苗'ϘG�M�´q�,d��Bs�<!@ߓc4�u��-A�R
F0�4#Rj�<�)�e{v��sɂ3��x:3��f�<I���0���ٍV�R� Ni�<Y�)F�Z������R�c��=�gɍe�<$�/�&���:Yʜk�}�<�r��#�ʕі��6ln<�@#�|�<iŌ@<]��M��D+#���3J�x�<��#AK�l$�!'`t���B�Cx�<��.K��v��@�ٞz��I��g�I�<!��	oi�	��Fj<L��Kn�<I� 2��08�&�V�m0ūZm�<A�+��Q�va�rj�sF�����h�<y�B��4}��i��L�F���/Po�<٠ O/�m��_S����Un�<i�� yh�A�̋*�@��5i�Q�<%��A����S`�`Qܔ�k�<��,u]�Ne�@J �~�<�#Ȓ��$�2VF�"E���� S�<�G됀33���֡E�7��U�b`QH�<yR�L�S`�1��W\4&!��e�o�<A���n��9`�]A��\j4-m�<�re�
KNE�����@r�i�<q'���_xU��*�A �bRˀL�<��V�^����C���*�J�s�<q�BK�I��#�h��Bv0<����u�<q�C�ڊOP� ǡ3,$Y[�"O8���N��[	�uh�E0M\!��"O�1�4��V՞4�rD�L$����"O��r,�q�4!Pb̬W��1U"O�� �˚B"�A�aO� `rY��"O A�c�
D��+Œ:B� 6"O���g�s ���NϜrK�8�"O��b��F�Hh��Ԏ��\�,���"O�x��x1P��$�9��`"O4�aP��=���`EGL���"O����'S-",9b�T�8�h�c"O�A�
)��[�D]
��xs"O�Q�'���9 e���\"O����&Gl)y��e
 � ""O2\�3��i� ۥ���j��"O�(PՈJ�y���@��^�\)�f"O,i�O�"�d��S��]�1��y
� ���#�L��h]��F� >#jh�"Oڀ`�(�X��f�݋`xj!k�"O��C���=�p�F�� ?�����"O�%�Pk¹D�vu�#��{�	��"OB8SNS� ��~h��"O����5�}2�_m�hXA"O YQgd]�^��@ь2AaҨ�u"O�1piH�(�|�R���N��)"O�H� ��Bt4���ލz���c"O~����dI����L��:T�4"O��B�#o4�W�Ƭ+��tf"O���
��'� �� fS]���3�"O�lHD6:��B�.��S3|$��"O��r��Q
N�!H��[E��C"O0���BK�ν�2j�x��슱"O�1��Z�c�Μ�E���9&x�4"O�	0��'��! ��U�--jq#�"O�M#�
(Xd4P���	�Bh""OV�1�N�j�aV ��R���0"O8��ąl�bȩd��J�Ф�"O�""��" ,X!����i���!"O��iTɌ�ixL@�Ǖ�T����4"O�*��x�;�"S�N���"O�T�c�T���vdT�%��10!"O�(����Ml���MI4���Q�"O�aS�<�"��G���:\�jB"O@ q��@���k�@�~L|c�"O������j^�M�B��"pm�i"O�ț6h�;v�h���ǀ�BZ�-Ѓ"O�:�n3?'X C2�հ"O���t��h��)��Er��I�C*D���rN5w�2�ie���X-T��I%D�x��拰4��ES�+&#�
��&D���œ:yR��b��L�,�qe*D��L<Wh�|�Av�@Ec��)D�DX��Y�>r4���pJa�E�#D�Ph#.̜���bdꔕ'b�zd#!D���M�?;r|�' ��{B���+D��d"$�t�
@�.=��L�5k'D�l��BD�Kyd4h`jι��p�T�/D��"B������H=*!���w':D��%m�'BD��bvD�Bf�p�$C*D� ��c�#�(! '�"J�t�)D�`�C$�!G��	��Sdia�(D�0�0B�I0L���,8j8]�Ѣ5D�T�c�èf��HH3)C1n��]�a*2D��ۓ�F.{˘��]�1�Тc.D�H�q�Y���\&>/rIK��*D�trO+��0�3Ɯ _DY�dl;D���K�)�Ղ�%%#&fEЕ�:D��k�!�M�J�1�)k�^����2D�,��DT�^1��)c�2M��E&D�t8F���gYn�)�M�L
�1D���S�z�\���r\�@g">D�4b�Dͬ ��Eq%b��X���<D���T40P<�Gk�
2lm�g D���NֺBaP[C�H�6�.)���,D�|�h�(�$x�w��q=���*D�,ۑ`�N2�Z@d��tb��%D�h�t�W�z��� ڄ�x��"�=D�	��� X`Q�s�K�lxƦ=�5bv�b��@�F����R�S��O��jԡ�.1��[A@�o^�4�7"O� �'��12J�4I�^�6s���Q"OD�X#���Y���r���4bOh�c'"O� vy02�[�\p�Nв\K��"O\m�C���fձ oW.L�[�"OH��C�n�TqR&Œ��#"O=��E+�. Г�!١�"O���Oƕ�QG:1m`ԣ�"Of)�l��*,�F��2I�Yy�"O�h2�J�Tt��k4.�=æ��C"O�����Y�e.�i��L�8o�2�A"O�ԙ�@��4���F���"O�(j���q �q��%J<��f"OZuZ����4Myǅ�*,�8���"O�Tʧ��F����c�:s�{"O���`.̧="LXad��5X�I"O�����9 g:��d!֐ui^E�"O��hu�Q�vyƱ2Bޤ#M�ի�"OΔ����y����@V�8n8Ʉ"O�QIc�&X��5 �7d�S""O�[�T!g|��o��04��"O48"��H���$�a@�f�\�{ "O|Ȣ-�=�6��EO)���"O@ܛPc'f�))5��ޜ�%"O I�����#^�QB��|~l���"O�I`c[#<:t�r���5jg��("OR�G�X6d��`����Kp���"Oŋ�� 
�� bI��Q�"O�H��OB�1(��ڳhѢQ����6"O6th��9*�B�3W	�6���"ORD�ҩY_�h���+{��Um���ydF�$	�Q��D�OjT������y�%���4 �#�L�B�*�p��]��y�-]���d�":����$���y�Aɑd��B�M�<.��$b��J�yR��<�p94Z.��Кt ��y��H C�h���67�4a�U%���yR�ʘlK@�C��5	�+�A��y�eZZ�N��Cs��xb�?�y���+z�E�e��8lq M�����y��	���FL�)�� ��+�y�a������ ƕn�}Hg��y2�ۚ�H��f��Ct��D[��yB�Z:�sq#!<�`�)��y��RĐp)r�\�V�ڤ�f���y��߬
���B�$�f�3u@�'�y��'F)���uB`�`8���y�Fݪ *�Q�h�
UP��@��M3�yb�I3TG��sЉ�BN��ȁ�o!�'0 �ѐ&�"b�9ʳ�Q��JI��'�h��AKB��"�0s�ɚ� �[�'%���c�;.$}kDUx��=	�'��)�϶8�9�Bųr��]q	�'��5C�k�"ʦ8P�k�a|p�b�'����KX4pP�ԊPN�d��)��'#��`�m�26t�n�U�X�0��QK^�'����+�V`ju��d+D�R�)I00�U���D�v����w�;D�T�s��z�,��"6�J��'D��X���T~8m� �K#9��-0?ъ�ᓪb���L�¤`� �Z�T��C�I4l6
I�pb̔�t�` �֦ZlC�jP��#D�=/�yh�HZ�8�(C�	'BVQ��R1� �-*�.C�	!�����R	i@���H�C�	�(�t�B�#F3���Vh^%B��B��%+2"3��� -
�C�L�0Y��B�)� &���%�ܔÓ�@��@�f"O2�K�J-�̀�c|
�r"O@�dc� !iF\�wN�kc��)"O���1R&hӢ�D;:S���"O�8`� 2�5�Ш�X���a"Ox-��/�7`,����&].�|��"O�pA�̂�{�HM !̏%Z�:�"O�P�	�"�� k�8z�H�@�"O�;ЬY=�h�Y&��A]J��u"O��;��F�]�����
��gx��yB"O,�e�3?D:����07uh]Q7"O�@p�M�Sd0�h `��5|�|9""O�l�,�.UBlC�T�E���q�"O�%I֫�q@����nW�A��K"O��s���K�*��"`٫�H�sW"O��:r�YV9�p1��!G���"O��(ǃ��I��l�҂۞B��!f"O���Ƃ�+<h�b�Z��(�z�"OX��e_<�}#b�7,��,KF"O�����ͨ-d�A��..T-��"O������a6v)�do\'\����"O�i��]�OB~|jĬ�$��`*`"O꼂ԭ>#�D����zq����"OX�#����
���3U�a�"O����Κ�:J����ĝ(���"O
� a$O�KD� �SmP��T��q"O@�[�G��kW��#ĩ��'�Ј �"Oб�Ԁ5Zѐ�Ʉ�p�@�*D"O&��&��u�����>��Q�%"O��" C�J�&��� ������"O��r�F�:w2b�h!Oŵ@w^�"O}�L��t�0NǲD`:5;"O�5YdO��S\��O֕L��0W"O��� F�hs�Q�e�lFʌ�"OAJÉ-y'��w���a��"O� X�@�%k��Ac�	}�.(j"O��Q���${��ٓa��#r5��!"O�1�sÖҰa�@H�'���"O�8�M��o�2�YRH�[��r�"O`!��Ԓ*�r� �g/J�b  �"O�y�G�lhfR<	F� �"O0���A�)�6�ٲ��1d(�6"O��Q�CR
z๨e�R �q��"O$\�&��;:����F�,'�R�1"O�԰�"�.c'n�u�C7�� �E"OD����/K��Y�b�� j-�"O��mK��Z)v��1��1B�"O�hHeg�3P����Q��]�̊�"O ձW�ѱ8�� Buʀ�7�4��q"Oz��M�{�¨Q�(�h~^u+`"OTIKk�!�8�BW*d`5x"O�P��Ab'�i83	�"w�Xۢ"O�%�+*��BA�M�]j"�cq"O�-��dĮ

F��ǀ�)
Tޔ��"O��!ӯ��+��a:Ơ��{<��z�"O��6�å�� +ѐy�f̓G�<���AE���@�6�6���hD�<��x��&M������h�v�<� ဘT���:�Ε,��p# �t�<Y\�� �a��N���If�� <�C�	$
n�L�7`��ѡ��c�dC�ɾ��]��L�i����%2zC�I�V��^���0P����XʒC�	�=�����/[� XPI(��^�$T�B�)� b�3N�3Ģ�b�n[-cSRP#"O��e�*���M^5}���"O�\P�%��o
Έ�a�Wy��x�"O�X���!B���3Ꙗ
�1�@"O��� ��&�B�+ҋCM,��2"O��@Į�F�{�
ن7�,KP"O>e�&����	���"O�a+����q�-��]��i�"O��b!j	���9�^�˦�:q"O�����,��(�)��	Pƈ`"OnA(�k��<6�� �:x�t��c"O
d���=�Ȅq*י�
9�"OV���/E����Q�(ʧO@v�u"OȽ�$n�5,�S3���Q"�8��"OD��Qb\�k��3O 4(5��*6"OX ���� �Eq�.#��;�"Ofl���V�>�H��̢/X��"O��/ƚn.IYҬ��*Pր��"O�MD��_�H���l����i�"O���0�4�CQfRw��T"O^5���S�	���@�GM֕�P"O��했}+J�jdd������"O~1��$J�B�xA[èñd+dt[`"OZ���&�a:�@�&|l�p"O�0p�N�):��t�$�X9Kp��w"O�� ѺQ�6�b$��& h8""OP�#�E��_��hTAD���"O�D)G�	CV��m�o�4x�"Ohp����+�~�+���ZҬ�Ђ"O*0���D
)�՜A��D�r"OZ����:�nD�¢�'��"O!@u�[�x ����*D��:"O��#�ű>��lx"/�_Z���t"Onȳ���0m��#g��i��"O@��!(���mSD>n-��"OT	��#Jq���Ʈ�`0bx(�"ORuA�n@*C.0񠥎���-�"O���e��0y�^�!n��?��V
c�<���\�W����4��Jp�T�<I�3G�~��	D�w���
�,�v�<y��
�6-��!�fL�m���i�<Q��h�2F���,9~�C�I�_g���dM�V���:��ġK�C䉗9~�ٳ�H�_��d�p%�G�C�p0R*
�������n��B�	�k�Q��#ڸܴ��'���!�ҩ)6je���újb��h@c�V!��[*8'I�3d^ܨm�4]�B�I�L��0�؋a��ap�iDL;rB�I"z^�BN����7j\pB�	�'U��Ufp��
Emߤ0a�C�	�]tU�q��\S�mH ݙN��C�ɈcV�e���P�*�~�����2H�tB�I�A[��+�D�R�z���j�s��C�%�jp�\2;�b�CE�A>ZC�I�7־]81�Jz��(˱_ �>C�I�1�-�Pkַu�9B�C[l(C䉿\ ������椠�+�+J(�B䉐G���!�ѻ6`�Ы@��)�B�� l8���F->0�p�*!,k�B䉣rY��4�K:U�X�P�D'`w�B�/�0p��f�' �L� �:{hB䉀$�p<9oG�!6�X�1,�%g�*B�ɤU����e��R��ِ$c��Y��C�)� N%�5� �r,�fMޘ��A�V"ONP�Ԉ�y8$�Q�d]�H�"O
Y��Q��������(>���V"O:���a��`ɳ%�k9�;�"O$�!g�++
��G�7� X�"O��hg��m��dJ@��l0��""O�y*�I�+���S���5~��䡃"O�i{�,���� e$�9pA!"O�Q�G�4C�R����NI`��6"O؍C㠆��Pmp����?5�]�"O4!�w�ͳܶ$Ӄ�7�H��`"OLh�M�-k�<J4#�Eyʴ��"O,q��d�){�4���Hڲ4xDP�"O���Ư@0'�<	�Ǉi���"O�5��2��)���	�0&�`�"OHI(�+ϮkJ��@9=�"�JT"O���7�؆e�ip���*i��I�"O��LQtp+���F�2 �q"Oj�$f���s�O�-"p�sLP�<��Ɛ5uG��ʖfD0���c�Dg�<�����gc�x�Ry��i�<�F��!�L�+J�� 1��Ym�<9���@���ؒKe��`�"Tj�<����&MK��E'��(7`Y��%c�<	1$P�vҪ͸s��6���F��W�<�&�����S���v�0�ۄI�P�<!�K�dp��U���Y�b${.FD�<�%a��A��Y��9�V8R`��<�e��p q�!��[������d�<��.Ή	yĔZa@1cF��\Y�<�'n�KF���G
��+���O~�<�eũoi��8���%@��]SU�e�<!�B�%9\�lc��,>Mv�K���]�<�ck�=	1�EA�������Vi�\�<���sj@��ᒣ2)P��P��O�<a�M�a^�x`@gކi���)�w�<I0AK8��0�v�N!�8tybL�q�<I�<@f��I� H5 ĳ��Bm�<�D��e ȋ .�]�Fu 	�`�<I�-ڷ'-h<�LC�7�� �NZ�<�RM��#� �	eEB3a������O�<Y�R�Y�h1Q�)-��b֤ZJ�<�IY�VT�� ��N���EC�<���)Y���e˞_Hn�B'+w�<)���a�`�P�A~q�)��
~�<�WaжGvz\�WN��.�H�A�^B�<yDK	'Ɛ���%ԘQ9xpSf'��<!�iS
EH�2VΑI]|�C�e�y�<��AX��V$��	ZX��Z��L�<!��:Z&��'(�<n.Ȃ��DP�<���*L���EF=x�>l*�F�J�<ч���Y�N���Ǟc[�Y ��]�<
�;ޠC#V�B�Bw>��ȓL��@u�sQ�U��p���ȓN)n�aB%�2���:#Ǚ*u��(�ȓ2,�$	��t����M�%e-Ѕ�ȓw�Z|R��6a�8
���j_�9��z�l)�,N�(��1'MR]�P�ȓ$<�B�g
��Z�+���]����ȓPo< ���yr�Y�H�!�f �ȓN#��s�h?)y��萯�
����c�%)!e6( ��K� 8�ȓ\�0���N7M��,��eM�����N�X1r��I?�b\S���I]�u��S�? D�Ƀ�
;���+�����5"OX��皦|F��g*H<s�;�"O�%B��H�8^h�+W,�/9gNMZ�"O x���QƔC��H�Gi"�"OޘJ�İ /0:�U�H����"O�9Je ��yR|�I��S?x���"O�f�	\�,Б��-��	�"O��sn\m�4h�JA�Iʂ"O����(k�����L�U.�`('"OT�ٳ�H0��lY�kޛ$\��1"O���� �o�@e?1���D"O�-���|�X(bfe 5�� ��"O,���S�d�x!��۸k���"O�1H�JU�f"�B牆��`Ț7"O�ER� �������S�1B��e"O8����D�:x�"���=�ʹ�"O�|R�-��(�M�1Ai�8)��"O�X��jD�~���	>����g"OR�,Q�@w����=��"Ol���O�tX8���3Ԭ�"OxA&s��4�l'<(�ea�"O�=���ǻq��1��� ��+ai!�d�3o.�p�ꁌt�R��U��Z!�DכO���!���<j����6pG!�$E~:h�3�M!,�$d!Sf^51!򄈫\���HTN֘+w0{���6;!��X<,��t�$�(�h񣆄�P�!�D�P^u�4�O�}�f�(w�Z�'�!���0Ӭ�E�5��Q2�]y!�R$;E�T�U"T:�$�P`[i!��W�j�\$��MP�Tg��k&m�5i!�]�.�*����[�i�J�����tN!�$ʚ|�ūÍ����Ze��(;!�d��;h
	1%̈́�`��H�	�Q:!�$ �h���#�dQ�*�!����!��%N���嗚`6�kRHK?@�!��o܂��FU�6��r�Z�\�!�G\�r%���"A0#�	a!�D�5�8\�`���4T��ȥ� Ky!�½|G.��6�'"-��9 �!l!�D��"�$�� $�e�n��B�_�.e!�I��L�(�ϧk�v<8����!�$���/�v~�I q�82�!򄄟Wj�z4�A�>b"�Jr�ª-m!���,|�����6|�0�A��	�'B�8b�@  ���B�g�/���Q	�'X��
 �Z=y��p1b��*�P��'oz�3��fܘ��%W�b�U�	�'G8 ��N�&r, ( ��FLR���'�:tC��@8e���Z�E!J1*�'�4 t�F6~?2��գ�/:�(���'�����Y�fD��*@`(���'b� �&ͤ>M,0qV�\�-�uB
�'��Mc�p}&��U"��)d�X	�'.���a@�,*Ϥi��ɞ����'�l��vl��8ha�"�'B��'�d�f��v3`��C�|&tz
�'�L�0���RL
�XF��-A]P�@�'>��I�*D�w$���ǟ6D�4�C
�'�j�A��@3A�  S��08hҹ3�'���hB��!qT�"�(��>Ԫ	�'���Z���wU,P��Oݹ5o��0�'id�H��$BT��2A�;y����'U�R��+2b�� ���{xJ 0��� $x�T�����<���A�"O�<zv�*K����I�x�b�"ON��W�(R�^�!'W1�"O��"�b׿M�@lȤ��o֒��C"OnMA�>W �xso�4�T呣"OD	��`9\X O��md� r"O���Ӌƞ!�h��o�(y_�Ԛ�"O���w�W+J�A0�n'UO���a"O�y%!�� ��1��vB��g"OH$����:�j���$f&�JG"O污cMˎeYTܚ�'ϕ���;�"O�DZ���I�x��G��!.�:yiG"O��Yt/�,�,�S䖎��Jg"Oq�uF]�"�&8ۓIX#K#v�s�"OF�i2�1&.���'M1�-k&"OR��,�T����z�5�"O,=r�JD֤��%�'\X@��"OԄj�)�<g�THf
�6���"Or���S�V�ZPQ��)���X"O�ܨWK݆c�NE
���k��`
�"O}+gOQ�R$ԠaHT0r�L{@"O���ЃR�����FL�a�݁�"O��KD�$ҽ��	3v��<i�"O8��k]���y���>��e��"OA��i��n �d	`�]�;հ��"O��ht��p�&���H�Ț�[U"O�!CR8,Dq����3�$mQb"O�jWk&ܑ��ڗq�P��"Ox��Tb����1
s�Օn�{#"O�}�E��).X�C�D 3%����"OT�P��U�CK�(�,�/dj���"OP�i�jߵ{��h� ��=Xb�""O`��ضS�ܹ�)݋P90�`�"O&i���D�R�*L�uh=Z��"Oh ���"z�=��BHV��12"O�X��`JA�"-B`�ϕP?4yj�"Oh jh�?(��ā�O�%U� r�"Ol��t�}�����$S@5nAK�"Ou!��	X��X�C$�l�X�Sc"O�!Zg"־Y�|��BC�-m�)�"O|��p�B�+���u+�:�"O�s��Ɋ5"�C��ԂA�ސzC"O�}��។g� ��A�3Z5�m��"Of��0�W�I/4� ���)J��5"O@�@2�K	1D䠨�A�W�
բ�"O�����N�RO2���ML
}}X���"Ol|�AY5Sĉ���}x��R"O�c�,N/� ���M�_}��W"O�|�D�L� �)C�C}8Iː"OT@i��_�~��y����>f^M��"Ov̐�*��)�j�2�+X� ܐ�"O���d�� �	qEa�:3���"On���N�vr�	h�4J�h\X�"Ofm��ą�P{ ����Y+�Vq�<Q��_
? -6f6� т�Pn�<�'���dfH4��<�tm��gk�<Q��>
��8� ��;i�X�	�c�<�Ӯ�_�=k���E��0Y`��w�<�����Yi}�#+��R�� p�u�<1�]� 4>e�/U)Q��Ѡ筇V�<�`^�Pi�b�ѭp��a�r*O�<���ܜu�z�t�E�kX���hIO�<Q��	C>��lϭf��C�m�H�<�V`�_f�K�*�xh����A�<� �@�dc?ZV��fd�7.�ղ�"O:<BU�4}����X��<X�&"O�a#��Ͼ��)"bÕH���"O���Ό=��a8���P~�HB"O�-�����y�x�K���7x`�|3��	՟�k�B��m����Ɋ<*d�}`V	�|���A� -B�qO���ֵm9 � BήJ��HfI�Hr���O�.�p�j�&fC����G1o��U����>c7� RT@.a�� 󃔬l����;�8Y��C�4��\)�n�%&
eY7	�h�'�$�����?9�i�U?ES3��
�p��Ƌ���eQ��T4�?Y���d�x�N(X�Ns��������p>�w�iD~7�nӼ1�Fo+�={�aA:���`�O6y1���Ѧ��Isyʟ`O�$��U�\�� 
9��t��W'!���޴(2��"��]	t��I�g���O���;g�Tpb�F�F�����!B�F�n7 �XP��7��c.P�g�zI�� ��c>��'L�0��޽n�B�X�\o�6� )]"�'kj��?D��4"Q�+���++t����C��
 B�'���|��,�i;��i%�IL�`1�ǉl�(�<��i��'p�7M�|2شT�R,���G!Q�������&)���H�Z�؃�6�M��
|�zTE�-�&����I�Aޠ Cʳ}=�M��X0RT��KG
�D�RO�'�d� #�R�:�,]�S^�aF�e�b�H��� -��m8�fۡ����	ON��Pg�xǓ2K��a�ٳi���i�MU)p>���6����Od�b���	��'��r4k�ls�dɵl�0�BH�<��I�D����l&^>��Ch=],���#�i0�7�7�4�"���<���S$D������?i�B,0$��=QD�"�.X���<9��Q[���)�r���0�� >�B�3�b�_cJ83c�3	)�����WDJ#?�!%y�F�I���)60�E1��˜y଴b$!�6D�>+0%�S�l@���J#g}
�Fx�O�?��48���n՚ƌ\۵�؀c�t�Cp����<������T�i4���U\g6͸��H�$|��'���	$��Z���s���T�k$��Ɏ�M���d�VDoZ���'>�j���3o5�d���*g���sM9��󟼛�jxӒ��5ϲ>�Tp[unB�C�H�Ӻ]�� �Ñ�=y��L#
PV#=� ��>���'D�0�v�9� _(������ґOf[E儺]䜥d&ϱ,���Dx�Œ>�?I�9��O2��-�u\����K�W�f�#'X�E���?��O1�n�矴"�h2�D���cǻ+Dy��3�OF�lZ៘nZ�)�E��$v�@d2"cŨG��4H��i/���.�>�-Orʧ��N���0���C�za��D_2]�0��d���4=�}��K�
I �b��t�`P�}���ߡ����`?�	��@�8�JG�j�R��'�ΨYT!��p� ŀ4�	���;�*O��s�����:i�-i7�� �^钴�hӚUsS�'��&|� ��*�禡1SKPG�@]ۤK�>w�՛ ���X������	D���9<�5��Ϡ%_�a��4�GzҰi�7m�O�oʟ��SϺC#��[[�|��Dّm�DD���H>4��'�a{���z   �    �  �  �  D  �"  �(  g,   Ĵ���	����Zv�Ll\�0R�PΓ����I#qh��)J��Z�V�Y�XB��-+�H���D�kr�yr��+B����-BtEہ'�-cb��q��*$�y���Q�L�9��2"�V�~E#Q��^T�XӉ]�R�p�^~JA�!V�pT��'�x�$�AR�չD|�1�T�A*Cj+��2��W�M.,^�%���0��w �K�JA�Y�U���R�Dx$���O��d�O��;�?�l�8("@�2��r�!��>ݗ'�bP�&>e2�ɖz*�����	7��<	SIKN8� �%�C�ʤQ�����
�j�<�fm�ǟ�Ii�	ǟ4�Ij?��,צz�P`�cɌ)r�޹u.�^�<Q�eڙJv������&D�|`Ң�٦����4�t�d�<�0��Ϧ����"��̙g���]y����'Q��'��]ş�I�|r�C�ڟP�FF΢5�nm�� .s,�a7�Є��>y�@^\?�lG=J��M(!��-u����F�Rx���F��O^�#��W�s�b��.z���S�gC覡�	쟜�'B�g�S�D-�g%�	B�Ϳ5���e�<��(ެu�8Cg��ж��"o�a}�/f����<)���-~0��؟�'��#��7�A�&4@*n�04~���ǟD�	�ig�Ts��%�@�	�X�p��
��X"�ȃ9Bu����@1,�}E{�@�9����Ԍ�|@Bʆ\����-��@RDI�$|�>L���hO����?!��$I�����{S�T���Q���d �O�-� +B�ZP�$���#:�{��'ܸ��(4
��9z����T��!�'�v8�'��'V��q6ҵ�����iī �k���PA66o�1�1e��M�R&�?Ɏy*��O����
5uh���ʂ'=����'<p�p���Ӟ,}Z1��I�%j�`�o�^�I��h����0�)�'��)R�&�/+�&|r�,T�b�q��'Ѻ��+�9W� h�-X�i����p�O���jq��<-��BeL�9�¼b��¾6���� �1��>��i���
�df��#��]^�<qw"�hՀP��"�T^�Щ@X�<Q�F�zLb5͕f8(��b�T�<i�&M�z|�2H�.W=������P�<��d��c�b�Iǂ������l�<��L�>��Hɕ%q�@!��k�<���T@)� ���ݖD��[l�<�t'�V�Ҽ�Ռƌlz !hu�Xd�<��NO$W|ꀡ2�B�Sj�H����c�<�B�m���4��F"9QU��c�<�G�@V�E���V���S��y�<a'�R-.�ty0u$<�q��r�<ɔ�XI�1
ղg�Թ���L�<)��F�@~D"��Z'�&sN p�<���M"$�R���@�AY*╍H�<�Ej� Na&�ɧ��6�r�k� �C�<i�c� �nE#�	�wf4�K�c�\�<a���9��I�aƼH��Ls"�r�<�A�)z���S��51��BҡN�<�F��^���;��0f�x���L�<Q ��V���yD�=����`k�^�<1E�4i����U��,�����D�<Q���3������
�
��C	@�<���%$�t��'� e"���[�<�"Ǖ1wL��
�gT4.�.��R��X�<��ؽW�R09��
������'�L�<YU��,IP�;��̝8�����bL�<�DN�Bw���5/�L�2F�D�<�f�ה�&$1��Z�F�� ����L�<�ǥ�#i`�"�ʈ :����"VE�<I���l�U�'ԏr�a2��H�<���L-��yA���l�D�q�`p�<a�*4�L#	�=9��dhGΗO�<�pmF�1ܱ����Z�NeBlO�<��R-#n!�FG�:3�����<T�P��BS�O��S�['�L�zTG"D�� :��V���h�|}x��βs%R�H"O��1���jaR��EY�R
��b�"OF�Bvf8��խ@<X͐�[u"OHqq�䅕dʀ�"N9c08��"O
�3a)��© �C$�q�"O�PX�j��x@ ���i����"On��"�(���RI� 7����3"Op���K,Fd32j��+�F����	��p<����;���Z�R��ڝ#�xh<�f*@
>�� 
�ض)H5�Ǝ�?y����8D�L��ɖx"&��Տ���P�Y
{����7Y!�I*;C��	t\�-M�Px���0=��C�6���BɵXl��*jM$:�'1��Q&���B$�-�F#}ZGÂ�iva	�xa����]�<����<"բ��>��M3�c�6Q�Xȇ(BZ�����Vm�}&��{ab��rX��Aϑ6S4D�h%��yej[5>�R٦����4�$	�)�xU�"��-z���t_
�z���K:r�A+% >�Rq`	��0<ѕ˜()�ɇ�C�p,@�ݥvn}@�>*@�������Y�<I�Ƀ�cGv��f%ѣ)*A@Q
�lyB���-� 	U	3�d���ȱd>���K�h��c���!7�J�SV�>D�\`���-��d��D�a0��d��%F؈��@^�;�$!IC�
��$b��J��73��ʗ(A=T�H��F�8�O��H�LARX�W�ىkL�ʣd�&OH��`)��?�����l�|������#��4	��[&a�%���-V�џ��,�*.���{���6X�x�혁y��d Ǥ��V=@ڰGf��ȓgL�y��
�L��H�I	-�>M�'P2�0&)f��i�0�	�-��$���
rPٺ +,X|CĴG�"C�ɧ$�]9�I����
f�F}H��̵#��ҕ��(�pb2`$�3�ɆE�RS$�^�py&# e�\B�ɦ?R�!f\~*�8)SE��p��SF
�+Q����J��r�����'a �H��H�ivP�IF
 hf��!O��b����b���ܴT��A@e@0s�,��@_2FP5��&��-�g�O)Ϻȋ���DM�u�O�t���7^	�I�¬e~�"}� ha:�HW*�}�2�XT#�q�<iaɜ=,����G�R�Z*�×V����HlyB��+N���Q� �a`���U�b��v��H�W.:4��vN�Hh��A�����Ϥ!����E���=NՆ��2�p@���I�Iit�b6E��U����dB: �Lbm�>�,_πD+�m@j�`p�S�<�Dk�1p/L�)ĥ�5-1��D��eF4���'$R&�`@��$.�����B�FRa��l��M(f��;c�݃#�K�̈́ȓt^�����:VF��␮Vϰ��b���y҆S���
�*/��h�����"�i	0=R�٢��0��<��Ved]��bO�et����&���ȓ��)a���9g�>����F+@���ȓ���& <Q�bPI��`!�ȓ/���TLZ�[�/9�����Ak �Y`Ǉs֘��7'�3 ��)�ȓ269	��܏O������MJ)zt�ȓ#�R��T;p	��	�D����` ������o�8m.4X���Gv�<YGI�,2���&@ a�`�q �u�<ٲI 4c��'˹-�\��cVt�<Ҁ�&WV`�F���x���!P��s�<��D��x�b͊5��Oʀ9 �V�<��m8xi$� ����[�<��/[�/��K����A�D�[�	U�<�� F#����u!�6i6��C��T�<��bS��S�1ji�Ĩm�Q�<aq�ӕ-AH�b ƈ+�>�8cn�<�b��M��)��G1+}���"�f�<� ����*��*��9Ca�z�A�"O���#C��<jw��a�
�[D"O�I)cR�t=���h�Pފ���"O>�R!!	FUXT��/[,o��&"O����͝W<��a��
"�̌"b"O��ED�	�l���G�h����"On��eʏ38Z�RcΥ>���q�"O�	q`�3 �q c�:�j��R"OX1��{���Qa?97�#�"O
=
E��=nQf�bG�]*���"Oʠ��b]1'H���&�!]ꀚ4"O��c!
JX��% '�0i�"O�(A_?���sE��1y�0��b"OXie�Z.V�\ej�.O�A�\���"O8EK_>O�j�y�I�85���S"O\=t��.M���A"o�S �ң"O�����X�u�Z͑�L�p��rp"O ��L�i^���A��6q�W"O@�b&�՟Wt��x�#�*�!�"O�ly$�P`?��!�A�sQ���"O&�ڗ�I_
<r�Q p���#""OP�[�ȄZ���Sƍ��1�h�"O�+v܊%���k�����y+�"O��A�ى+��yA�'éw�&���'�$�q�!��,�� ZJ|�a�'�^�B��s?.t�%$R�jE�
�'*�h��!r:\CE�F�9`6U��'E�0��Ղ"2<i���"{�����'c<�TȊ5#�>���)x�x0��'��49��
�z,����jD*��
�'��l�$))V�J�X�2�d��
�'��H�D,8� z�� �=b��3�']`a��/z�l��i\.8rpY �'�!a#�|C� h�'L�Y��%�	�'V4Ձ�!ѫ
yz]����l`�'����q�O%|h@`�N\$f�}�	�'&�4�T�ĝ�Z8biJ��XI	�'|� ��� �X�p`�E�=@	�'zp�X�U�l@��3폌4j�dx	�'���k��T=�p�"A/�E��'+�)�atEȶ��4f�҄�j!D�@�$�ɲu�A�(ٹF�[�*D�T5��);>�9 �KIR:H���6D���A��-� ���$�
d;�6D����lW [� �Eh9>U�HS�A3D�x��N=�xt����(d,�i23D��0Ƅ#U�Pb����!��e2�#2D�8�ď�͎<@%f�K�����?D�лŭÒ7i^ձ�F�!
��M�Db(D�����Z�4�MZ��.H��cFB7D�t�B�Z�FÞ岆)G�g�b����?D���-C;+���3A��wPP ��-=D�x:��1�.���&<yp��(D��{�ʩF����קѢW��QRb�)D��,�$q|���gQ�Z�z�+�@%D�:���
а�*�jQ1C�:)�%D�JDm�"O����홴@�e$#D�`����|Cx��)�X�8ӄ,D����'�2v��I!��zR����)D�#���,�(��Dl��c]��K��6D�,ل�*��a���^��u��3D��J���j)��-��%>�BuI5D��г��%�L�Z7�
Fi�D�5D�\1�K�=�d��Y���k�0D�� $p���
.���OF>"���"Oа����ո�[m'y��"O(L�aJA�J�}R���<,"q"O`�D���I����2�*+i,A�"Od���5A��)��T-*Th�``"O�����̻ ^D
 R�u^�a�"O-�����^ⴵ�5�G�^�4@S�"OHYH��6�V�(�NX	�x�u"OX�ECI7U�L�L['#����"O��{G�B�L�Ĉ �ʗ!��i�"O��"L�E_�A�e�?~}�<1�"OT��VH`y:�cV�9zt,�w"O"�jpaC�*�`h�GZ�BlA"O����b��[��U�T"G9�6��S"Of��1.K�����M�`��!jb"O�𰂁�7A�@Ie�_�D��T��"O�hҩ�.�H�0���r{¨�"OX�#ßJ�" ^x��KG"O8t�aoĖ*������
�H���""O����a^� ^��yo��W���ѓ"O2�r���Y���Ʈ�����%"O��2��^�)�L;k�H�v�1"O�DCc@"0�b�̋0˨�1"O���%!�=��Xcl�7�*%�"O$!x!�fz�5Q�BE:�b��`"O�D���S&����A�E1{�"O�R'�խ/��� �A�(1��ܢw"O����Kӗ<�ؒ�g�&��H:�"O\Țg�Y�!P��s抉c�`I:�"O� �5�_]X��
F�ڑ.��ᢖ"Ox]ف!^�N��� �("�Ll�U"O�ܘ*)+��!��Җl���0e��y��s�@LX�b��F�2��A߂.� ����&D�� �`��>�8���a+jl Yi3�%D�xr#�4n�|��ɖ �Dj�'D��	�R�=�0B���P ��'D�����I�^��E��
.�����$D���3ら�rP��$��-��8�#.D�pE�E�Xp���#k8@���.D�t���Tx���E�w��A�&+D�`S�g�!�x��"�rF>��� *D����^�b�$��Njհ�%4D��ǭ͡:p�U�4�g$xڢ�-D�P!#�ߒw��@���."T
�Y�d>D�p)֡U-v�r���*<M�F�7D��#£�,�
̢��
5|mkpM D��)���.n�rU;�I	�,��A�=D�X��%T�`P21�����G#��!D;D���$j�zO���B�,B���R�m#D��ᠧua�$a#��G�|�x%B-D�l�K͈;a�]���?sl`d=D��k�|�;u�\`6�R��;D�d���U�[�\E�c��V�]ZF?D����Bگ��P�+Ed�41�K;D��"�N�j���b�Lǲi�"a8D��"T��/�	k��&n�I	��5D����eX|�U e��#q���gj1D�$Ё FDT�P�C@/Wn�E=D�P���0M��r�摆H&>�@�:D�X�v�Vm���a�ˏ�~⾹�77D�ȱ�oA�2H������-�q4D�8˗D�Eb21@B��\����$�5D��[R��:t����fMe�$�� 2D�l�j�S��ҤE��F�����=D�� $�IB���p$��%�5_`�ab"Ot�jC�·E)������*�Ĭ��"OLuBFZ
H\�#��(y|(�R"O���J�4OL�
76wL�q"O�����	M:='��$ag���"O��q��<SA�m#�jE�eN&qK2"Od�1�,��{��K��]�`E���"O�"EƯ<�B��#-Հ]j�"OV8i��?\�Z�B!�Zm�D*"O($x7I��1����I�d��-h"O��Ƌ�bP���D�?��1�"O0ؠG�X�4p��N8�J�@�"O.�ٖ��N��� �b�a�"O�m:� =9�$���!X�n���"O�(]*LL���U$bt��j����yB�2k�hm�T ,��1%a�%�y�G�Bl���	��$o�QS�I%�yr���4g<@����O���r���y�dV[z�a�.H&)>� ���V��y"�M0HԈt@ՕX��#G��y.5Wd��bAS�a>�ڥ���yRi�M��6�
�]�qr�lS��y��?W@8���̗Q.�"wf��y]�@�"�T�\
C�С��,�y���?H�
9�'!N�M�Lq�B���y�,��o�����
Ԃ=Oq����y�CU�wU�	C���,F��qa�"�y�	*HJ��p�ׂ��� �Ţ�y���5��J�NL�7�())E�-�yB��W��qB�M�)w�<���8�y�`O%ִ1"�R�.��a��3�y��D��4�:���)Ĉa(��ԧ�y�J����
�×�"�Ġ�iC��yRB�8�4䌳i�ipq)��yr�W,q&j*#�V!h��crl�yrP"$]>�CU��0�\9�q�N�y�B5?~�`�-9��Э��y2�ڏa�r�r����	K��?�yҠ"|�8����2Q&�뢅D>�y�X�m6�M��6�h����yc�P��1� #�4t`R�`��y�a��@O��0��;)�����ش�Py2%ſʘ����,�則c�l�<�5��I&�`����1�l�<	W�H�K�Z-��gŮ8]��G*�f�<@�X�"��鐊���@I�Ga[^�<ٳC�Qm�HJ����!� dyd��_�<i2�
=[,05qU$[��m�"�KZ�<a !@�`�T����`܄i��g�\�<�G�2l����';���Qo�S�<�A��eo��Ytb�tϤe��h�N�<���8YP:1N�{2@�-�<@���I�G�1I��:S��}�<�0\�dذc L�hhaZA��x�<Ig�܆5�d�0��l�����g�n�<���a�8���%tks�_�<	���:/{LP��
u����J�X�<��GU.|,k�^d*��Vj�o�<Q�J�64p�c �	5�ڕ�T�<���W�O	�=ᅇDS�p�B�M�<��/��"��p�6�B���O�<٥�"��4��!��ld��95ʗH�<I׉�
JOn�+�k�
����O	H�<i��]�XFB0��.�vмs�n�<� tH�Ď�MĘ
'A��*�8�"O�(E-ǥC�Mh��b�؈�"O�`�BP�Z�R��w���-��"O��!S(N���A녁"1Q���2"O�l &���,��#'*Ős� ��"O�$��L֪5ղX��� �J���"O��b}@tz��M�
X����"O�͐��;�2A��&ϓ ;v�b2"O�Q*r��34��Ř )����"Or�dC��<3�yӓDF)#V�:�"OB��DD�<5[��;G�]� "O��@�)�P�9�3,�0B"OZ�1����\(C��oE�m�f"O�Psd��/��H3`�	U���A�"O.٠ᦕ))4��N��u����"OD3��;5�(�'�V'+)h�"O�!B���v�$��ɸQ���u���Hv�' 0�Q$��")�ztX'µ��ݱ�'a葐v�57����a756����'r�QJ��4Hc�$���;d���4�hO?7��Kڊ���L���lX�r�<C䉎;�Ф���a���m�;�"C�'j�R���2��"oV7^`�C�	-O���KRQZ\8����XږC�ɵ_�2(IPm[�R<�	��ڏ6��C�I���!��I��6��bC�lC�ɡR�tSvk4���R�X�|
B䉇D�`{���[E| ��I�p��C�I�H5�`0JQ�pI��Ӈ` #��C�ɚ)\=@��4n[fY��
݄8TC�ɎZ��Qw(�<�f8'&V<sFC䉘@�|�P��-��<`gh�E�C䉘?T	S"A�:l� 1Z��,�TC�	�jA��Y4�9��$�Cf��5�VB��=��0��*<���!�n�pB��,hx" �ӣY�-�Q"��/5�\B��e�\0�kǥm�8Y27��$B�I+r�0@!DC�8jm�F��JrFB�	b<�EAS�<  �An�PC��T=z �bF����'���g|C�	5\�Ң�Ȫt*BX��G�G�bC�7DBNT/KC8��LQ.H0C�&S6pyҡڏ]���&J�A�<�=�A�ٓ�B30�(s�˛� �i��6쀙  ��>�
�J0@�&��$�����IE�Tj���$@�(M��B�4x���O�4֔󠡐��C�	�'j�ۗd��k����Sm�)%��C䉠dTT8��A�;����@��	Gw�C����aH��b~jyj���cH�B��C�E �(��;�>���0��B�ɇd�}Q�jL��܀���� bZB䉓X���s��I�<���O�b�\B�	<_�=PqB\�rtR����A�C�ɽ(�҉+��xkT���`O`JB�	#Qo��#�/B�-���	/+pB�	� T�"��3@e�5(Я��.BB�I6�H ������nF/*��B䉨.��!��	��u���)��B䉨I�l�c�F�&_�4�'OÕ5ˡ��W	R� �g�N2@Q�Q��`�"�!��Xv3~YvÓ'0Hz�IP�ɽ21!�$��Ԋa��êcE~�(0�єX!!��ۻ�Ј � W+.>u�Dm�"<!!�� ��36/U�C4���e'$pe�m1c"O
�h��
	N�⢦��w쐂"O�y�i� t.ʠ�U��v��%�"O��He�ѩhR̬�D��W�0�P"O�PZ�B�"x#�x�Qd�W=�m�"Oh���I;{ԡi"�Y/�y�"Ot�҂8Zæ�(��]�8+�Y��"O�L�w��Q�A�A�H=(�|�6"O��3����q[�9�Eȓ3���"O�l
���VF$��΋9e�B���"O�t��/��m[���3~���"Op��aػ}m�xɅᙎQ_��ّ"O~��㚢=d��B��?IqyC�"O =w�45��� SvH�[�"O��
����h�!��K�{� E2A"O4�1�[�'�j���D��4�6��""Oz	 @[�*x�#2�ھr���0"ORܣ�I޲7�����W+����"O$�Y2���1�tX¡#�_b��"O:h�E�;�	�( 5,mCd"O���!b4}O6<"�F]�>���"O^E�c,F ��4�u�4e�� ��"O^����X�,L�(6���"��M:w"Ot���"{N� k�bG�L3"OXՂ��V�
�\��*�̄xq"O0I��NЙA��[��K:&�ԤK�"O��hV�gT�(�C@�3�F��"Ozغ��#�š�N3N��	1"O\�(��N��ո�.C9�`EI�"O4X�U拶9�na��C�B߀��"O��
fQ:em��C��N̎h��"Oxad_v�^I8䠃�'���Y�"O������B.���QFĢ~2�zf"Op�����@�j�9#�˱V��x'"O�P���]�P,@���,uF�iS"O\b�Ż1L}�q��oi�P��"O��a��  �   /   Ĵ���	��Z[vI�>.���3��H�ݴ���qe"��A,<B�is����C&��k2�Ɲh3���a��h��6�DڦŁٴ8��{2ރuB8J�ڛ{��x�^,}�<������O
��ߴ]B��r�%K���0�G�:2zI�'w�x�bň�u��H-O"�g��>�r�YR�������wY̡��O�3�����Δ'N�q��i����s���1�X"��Ξ1���ԊL���xA*�48�`�&!L�e!ʾ�x@Gx"l�p�'���rU��\�b�r�I�GT���N$�$V�O��N>)����YY&�Y��iz���([�<a��=pLL#<�.�72��� d6��q��Ha���r�\��I7"��x��JM�e��&�av��'՚�Dxb��l�?$�E��fֹ2����B��mڇ��l���I�m��Q	d�"K~̀x@Lk��H��*�	%=����T��Hac@�)�Rq�&D�:u�0T!��<�­%�5VF����Q�F)�"�"�!0���iD�\�<_�dHb�ɮ���ȝ�6����M�Kn��SR�ڔݘ'��!Dx�&�D�+�z���f6�ru��	 Ϧ�	�����I:iD�Mk�$�s�T�r#܄Z1��d?}�C�u�n4���DM@��bT�;�6L��kQ�^�F�{����?_���'F��0�(M���b��!���GR≳<m� ��Ί}�@���L۱TWX8��+о�<A$�t��
w)Xr��q �ozYA�j"D����   �@��>$�=A�D�nkа�U��ğ��˟��D� �L�<�O��bg:@*ذ�#�<RwD�Ɋ�܇��?q�A�IߖiG���)�.�D�*ʓB0�`��F�O�0M6���m�� `��>tY0�'0� ����V��Q��?Aw��Q
�2ɉ'�L�m�a+���vg�B���;�'�\ ��z���$�O˧1�Ze���?������:��܍ �t�J䀁]�P�����?�y*���xQ�١,0��<D6 T��/K
4@�Gx���'�>����K.q����TA�{�r����*:�b���Oꥹ`)�c�� �!���h�c�"O�l"���6Y���ٽQ�y!��I��HO�/Y�rHJ��lψ,B�΂=���I񟈐!+A0?{�(������̟$J\w�w���Y��\���4��b	8g(2l��'���i�**)p���b4�\�c<�LP   
	    �    i%  �,  83  z9  �?  F  \L  �R  �X  <_  �e  �k  r  Hx  *   `� u�	����Zv)C�'ll\�0Dz+⟈m[k`�,Q}~�D�\Kv�Т�íM.QQ�T +g�4��
��f��"k�WO��e���E��� ��Q&���')w��C�j'����<� M;N��~и�eԨ!-�{�.E_�� g�� PA���đ�G*�e �(~cD���F�HI%Z),7���ɠ_����fnK.+�^h��4e8u	��?���?A�'��9�Ch��6D��"�%Б5��]���?a����?Y)Ov��å �J��O��$.v�v�huG�Џ� �م��O<!�4��Ƒ	>��i�����?�㣯����/\4R����}����oD$�˵�2=�}���A��F$�'��#��2=���Ɣx��%�Z���$	�J����(�?Y���?���?����!����c&-!PjDbso�mG��d�֦cش ���'�>��i�46m �E�ش�?	��X�~��ı"@0
�l�����y��Ŭ'V��� ��� �� �N���S��K��W̎:mW�6i�N	n��?��� &��cF�\
��`E�#)*��)J:h�\���f	R��d�R:֠� ��U64R��Ib�'�OГ%]��3W�9�����x2�ܘ|�bc0� �V9I��
���O����Ob>Ɂ������r�X�r��7L�<�����9�"1�v�Ԥ�H�م`�6I�H��	S�',�'$ڼ��O%L� �k��muC�A#iF��8�'�]Cխ+������fJpy�'X�DJ7�z���n1Xy���
�'@�,�P1p
��9.`
�'^�uA��QO8��DG�u�}+	�'�ȹTFS�PB�C'@��v5�8����<N�Q?ɉE���8tܸ$�ܡ >�irU�8D� yկ	.z<�h��J[&u��щ�n!D�`p�M؝&�z�Y�)٧"��}Ps,D��S�C(�J��n��4 rm� �7D�P�Ȕ�����Ue&(Ō�I� 4D�L�s�ج_q�D����1FHxJ��Ov0��)�'b.���t�Ñz�.��/tJ�Q��'Y@�� �i����I�9��'����D�
]�=Ѷ�	s����'���.m$,	Q#CS��;!�q�<I6Ɯ%������ve�t{#�I�<���z�hइ�]:R��HyRnL��p>�Ո��t�t�{�#OXM��
A�<�)�
\��-Y2f�8xpaj�az�<��!��"��´f�4f߮�I� �r�<5�Θ7x|��ǎ�	���Y��p�<�3p�̚� M�0J ��c�cx�x2gg� �'��H2���"dl�¥!I&(.��Ó4e��c�ݳ:;��'ris቞+&��s��Oh(Óf���h�R6:.�'9�e�����d@`��LE���u\��Ο����HZ�D�]=t���f�Hr�l9��|yr�'�OQ>-9Bh˒��իӥ�7��YJ��<�O4��ɕ?��Hvƍ4�%�Y
'e����<y��?����'z�DA	!�21�-׺m��y��F[��>O�F)���S�W�.U���j�:,�sn�{B�?��9��2�)�'2�E��hA�jQX�A�w �|�'8�(:���?iI~���4���iy�y�B탽�į73X,�Od�d3LOPA���]�W�ذ��d
�#�*�sQ��9�h�&�1��E�>I�p��'%�E���r�P�d�<i3n]��r���Fk�[w����k����Pq�,�B �<�6���hߊE�|�<��i����$H��V%@��@�\.�,4*O6�If�M�@a1�1O����8yZP����
jZ�5"��'��	�Ԧ��&��O����Oh�;r�R�$'��t&;X
x��3j#D�L3�\-P%d�������҆�<i"�i>���xy�HP5|Y@Y������S��A?q�h2�'�a|Ҥ��(�`��@:ht�}��/ވgܤX"�'o,А IX�TJ�PnL�j�
�� b�)�!𤒱~�zy�AC��N`j`���W#0 �@�q�'d!��N�t���gՔJ�\5z�oNVA!�L�'!89��N�TM�d#�-�gE�'�*7�;���6A�fQ&��#�H;gt��CMҸ.Z�1�h�O6˓�?a���?Y��՞nHb�� ƍ+@�MF�P� �H3Q����7�'+��l)�ɑi����bc�@2������_PR�'��'���c����300T�f&�_wP�1�Q����]�S�O�i���Z Q���r��;��0{�H��B�A��Z���B� ��I��?�/O�`����¦$?�O"7Zr���Kǌq�|ɹ ��L�"�'��Q�Oم9P�A��J�<E��#��jߪ�P4M�v��t�����Dл*��y�eg�)���2�7����8INBy�Ǐ�K~"[��?�����'��O�t[�+уw(t���D�X�*�HL>y��0=9��τ/��I�$߾S�<��F�\�'�@�}r�a��|i��1`=b�n �0n��40`�Sp��|Fy��\8����ev����Fe�$�y�C����Kr̞�@��;1��,�yB�Иe��y4�����:&�
��y��.e��` Z�NE�Q�"h]3�y�i��V3<�*fL]�B�T��P�R��y�d\��-03aV�l�=H0�Ν��$;&��|���3�`�XDc�W��X���y"�	�����b
�_�ɠG-���y҆�G�����I)S���z�
۷�y��l�(i�E.EV�a7F�)�y�E#q�9��a[��7C����>	��Ly?Y'�c1@��Ve�I���B�S�<Y1MڥB�bʱlT�0��ܠ���H�<��[�"/ T{�$C�C�e@�H�<�����������0.���W��M�<ɧ��8|�@�x꬙��e�<��بs����.�:7}���H�E�'��ʉ��Z	<��G�S=+$��p���S!�kl������`٫�^>.�!���4����l��t�D#��ߑ^�!�u%����'|-�I�V�@�H��W�`�[�O�00�x�@�l��ȓi�������c�Ţ7><���	!P0�#<E���.
�}���'�ؘ��7b�!�Ę�H����̺M��`��1�!�$�&h�`Ɣ?���Ço_�U�!򄄅W��8��҇b��{���1�!�$E#y�R,��H�6%��آBl\�y�!��̫h�1jr$�7h~L�Rٯ��	.!�����kd��1���kjF���L��!�D�5Q4����B�ad��P�K��G�!�dBT��4�Jʳ!O�)t��m�!��|g���R�]��D�&�N�R^!�ڟ�059##Ю Z*d*�̑5*N�}b#N��~�-���Ty�H;#����l�+�y2��+N��b��5s��@	ؘ�yR'D�>�(��&
؞&����4C���y"j�;,�����T��t�Һ�yRH�I/r]8��7ܠb�-���y�)J<�Ќ������H�hO��q%�����d�H�D�A���>B�INa����T�k��J�+,�(B�ɵ�H�cac�i���	�+%6U�C�ɒWB(��7
ΚvƆA�T耨T��C䉏G��u��eKd��K")�B��5D+P-���!�hؐu��9%�L��
�W��"~B� ���3��Ӝ�,5�d�̃�y�⒦!�us�CX����2J��yB/C#|"���aI�.%����2O��yr@(dD!�	��	�'���yr�W 4Р�;!�9 �P��)Z�yRHQ(@O�)"Vg�|�5
tGX��d�"Z��|�jD�]]�x�mS<�<@2���y
� ��z���\���b�0,���V"Oڅ���#k��F���?{F ��"O:�#���..)�aС�TR�=)4"Od�il��Xe�!�nժN4
] ��'�����''v]C��*Biڡ"7.�"�\�h�'f,�+EC��!@�'�My�'v:��d��	f6���J�'p�(��	�'�~`'��@ކ���s��'+B@r��$��,#�@l�]r�'��M��:C�R��qbЄ\��B����,Q?�Y�ۅb�x���
�
�pR�5D� !^�\�Xӧ��w�mS�<)�'r�ް��'u�̀�*V�<�Q&�)�ґ���@	\o�x�k�k�<��d -z\3�̍,26p��P_�<I0��(E�:U�ag�
�l�#��ןp�sG,�S�O��8�M" G�����y�&"O|Y��2�Z�`�ʘ�#�퐥"O�u�#@:xa�=��(�.#���r"OnDS��X4 �#g�"�4Q�"Oʅh��	v��¤Ņ�,�(�)�"O(�� �_J�Jr��%�f]����6�OT�C �Ҧ��0�B"Z $�2Ā�"O"8����1R��m�%�&GC^���"OD�=�y�"@%C�"Op;��ΥJ� 8�R�}N��"O�35��a�(��%�� ���'P
�A�'
:a�sXx�H�,�$EI����'3fPg�
)`� (�F�
<-!��'\��k��:��+�Ԣ/v��A�'�$#��
J�\Sac����Q�'D����ƈp2����ٔ!1�T��'#�\��Z8<0���I�6�-n�P�~���-d��鋗F�  ����I�<��
�t���B��j)3��G�<A*ںT.�D�vkW1JbhUQaEC�<����x�
�qt\*Y�h��NKW�<QCcȋ}H�@ǥ�25��`+XT�<�f�,G���a��[��e�!�ӟ4���0�S�O���{q����@��R�^���t"O�	�k��JN(��
��F���"O�1��m�=M�U��n��2�ByQ�"O6ػ��6]� "�hI!.��U�t"O�R�G'L|���I��¾���"On��Bŏ*�R��gO
���L��Q���I!�Ozt�'��z�A��n>i䁹�"Oع��Wv�t	9�ğ42m��"Odi�M�n�X�9��W���,�f"O������ "j�'텛BL�Lc�"O���j^�	x��R�k</V�Q��'Шi��'ĲL�D�%^g(QE�R�dN,�k�'�H�33kI)��/_���q�'�L���+4X�J�'�J$L��'����Ĥr\�0�#tYx�R�'�~`�n�3=��9�eÍ
����'� �B6Іgs�Xp�h�>��T��$�?AQ?��g�"6����e�߯
�+F 5D��
�
W0�8�O��Ro�%��?D�XY���O~B�*��N+����0O>D��!��n~�c�*����	/D���)W�7x��ɵ��7�k��1D������{7��-wM����O����)�'?V4lh��g䤹�c�R�b�{�'�P��D,�J�إ�oƐNV��R���  ��p�f5�r(��q��a��"O���HO{e�@�hH@�"O\M[QBU-x���@HQ>�b�"O�j�M��dæ�Kة�X��h��$�O"�1G��:m�@q�hD,2��"O�4��	j�I`�H)Ud�0"OL5�D CRl� ���$n�r<q"OX�;��hND���N ��Bq�2"O�Hq�F���ŭU�U��� ��'>d��':�I�.�,$�JIawgXנ���':�Ta���
1A8����7L����'턄
�mEQ��ɲb��5Lrؼy
�'�L}����>vt��ƃB��Uj�'����,AO:��0NܜF���	�'����+*���Y ��/�N����d� _Q?�1'� ���*�*�O��0E-D��b�D^<� ɘ�Z��t���6D���!
��(�b���"�^p����(D�(Ф(F�4L�3�R!0x��35/%D�0ȧK	;G ��j�G��Q�� (D�h���>����+�!jT�g��Ob��)�'g���x!/Wh Z�'ҔUU���	�'eY�h�,=�0��N�F�\��'(��i�-����R)�C�f,�
�'�q2�ʦX�`E"���n�V��':ʠᒪf����j�9j��H��'�L�����<=κ����x��/O
���'����� �, ~��R!۪n?B��	�'ֲ�����1_"���J���D}(	�'��U�u�E!\�\{r�

��\(	�'-������X6�X�1��&�)Z�'�<�Ȅ�_�?�<�Κ�Un6h�*����.��-`����6�����^Ň�G��=��`	-Q�4��`�#b�p�ȓZ��)��-EN�]��l����ȓM�����m��+8����ż8|���;Ÿ�r�kε#Q����nX"7������9+��%W����ʩDl��G{�`�����4h�eܽT"�	���)��8# "O�IjbO@�[���;%��>��I&"O�Y`S���>�0��S�1�v"O�Q�#N��p�su�0���1"O�����Np聵gE��K�"O�z��L�	hJ��B�v9�+�O?ɲRi֢rZL���� �t�8���p�<��-�#��qsM��i�\0��Q�<���͒6~
Q*�bH�Z���BO�<�d�M�NB��p�H��B��t�<!�
s����c�K~�MB�#�s�<��o��q�|Cd
��~~�x�u�gy��N��p>q&Ȗ�݊��0+��#N*�Е&A]�<	r��#<ncc�ˈCHt�8�W^�<�5ON�_�Za��L��xX0�1T��#T$� ��a�c^�o�,�4"(D�tYD%M @���sB
���e�N0�O$���O�@bv�
 2��1�mX3�n��'"Ot9�A�ذ_z�p	�
љ
/N@�!"ON� ���u�R�;ej��X)#�"Op|��`�GD� rH�!&A`7"O����R=��,�G�.����"Od=���͍8�� ��j�F���	�&���~B�+���;F��m�ک���j�<�f��4��b�%[�~��e��e�<Q�@7Xtj�&�Ԍe\�M�� �e�<� �X�j�%*��9I0�U�5x�"O��P!�;6;p?;X<�u"O��0���5��S�l%4J�A�՟����?�S�Ŏ�ؓX� ��o��:<jp"O21�� 	��0��!Y9d��"OHT��^�C<�P焼~�ddpF"O^�M�EJ0�K��� O��21"O����a^�]���M�L0�q�"O�(A��E/|�8�B��'`H��\��#4�O���1���fGn9��`Ubm6p��"OV1��h�
E>���cʺQhp"O� �G.I>2W$�
p�ڿ�t��r"Oʽ�0��nxҌI�MJ%3@�U�"O �2��;#8T�
�*δN�� ��'u\��'樌��Ȭ[<-��@�,=�x��'���)0a�u�,�WEń0yz%��'b��"�ܿ5��fOu5��8�'~�HP�˩-Q�4ڴ�mGH��'~@��T&^W���#�j�XE��'Ւ�K�߰L��,��^�t��d�
Q?M� e�$w]\��C(�=Dd9k3i>D�I -����(
�Ni,`5��&<D��F*�8J@�h�+kH	���=D� ��W�v	H�[�d�%�TT���;D�p�[���I���T
m��# h�!�$	� ��t�5σ�f�l
���0����O?�� ���( �O�5p�p�â�j�<��B�ylR�����e�>l�֮h�<����d�2��Yd�P7'Se�<y����%�x�qG�O7�.,�v�d�<�T�Q�e�R�z�N�`=�aJ6i�zh<��jV�i,�D{��Я#"��Yt����'��}�=J��$�#BrlX���%gc��#��B&������ܟ���@�
+u��t�ЁE6p���|�t�:(a�-��]�W)b�)�C Q�'�p���8RdҔ�6�哴�rY)�ɀ�4��}��^19�">�ƢX����u�'K���C��.lSh}[�^�1`
��'�a~�+�}���2��^P�!�����>�G\�КЏNY���r�+��O]�剓D�R]�	柌�'��⟈�	��$�1G˘����R&���II8�
W���?�m(�$T��?E�4�� ��	�f1��� ���yBo�y���ueM�`��F��'$j�փ
]� �7�ӈ��!'�.��O��S��^~"�T�[����7M:��S���yr��H��A��C�x̓�� �hO��F�	�K�D���]V��%��:	7�P�\!�韜�	ßP��Qy�O^8��L�I��2q�@�-h1Hrfȉ]�iF�'H҄������I�Z��J$�A(K=~�*��p���������˗�ڲE��Y ��#Fx��H=
(�l�z%Hɛ������d$4��'ў4��rg�=�X���˙�T�&x�" D�Ds��٩[�0��j�#M].�x���O``Ez�O_�Z�@�4bO2<�@<�g��`Zq�"(+�ލ��ן��	��Ė��O��ڤ�B&  %��OQ	n�p�M�:k�Nt9��]�8���� -<O�Ș3,С(����&֨5@�H��q�n��엠O7�=� <O`���'N�1�
��)�̢D"&h�V�RT�'�ў`F|�7�����m�7d��u�_)�y�)/1F,L�s�ڟz�(�%�C�������iy�"M�r�c?�Q3�T�}c���u��|�9���Zy��'�'zr �&��5Ǩ]�#&�+n��4�b�������&�Ϛ:�����,ab2BM(b��x8��QI��%XB:��a��4B�p�7+�'��O�+R�'b��5ö�W��yZn�	����&�	П`��*8 �J��%���&t�.��d�Yy�f9zmH��Z2$t���C���$Є��Tl��x�'8��|�	%3��5�PԸ!s6�`��)/���I�$��)b�a�5�E�Q�U��uG��J[b��0�,1�(�8dB�y"W�w�^�+��y-��8��\�O�z��Ff�4�X��)5]tͱ�'c��I���䧶�� �5���I�p٢u�mW�qD"OH=����;�t�"vE�?VKv,��I��ȟ�({�C+=��8����~�&AȇaQH�����3�{�Tpa�Q	4��7�ܦ,�*���H�I	���i�^5ʠ�#:UF,�ȓ
�h��V&ɍC���RN
h�ن��>���
�z� ����M*e��56ڄC#
^Y�P3��N�8���?ݦ!�UO�mn��5�MwU���&
z��$T���l�"K�{��p�V�h!�ɔ_+b�H�7��e��)�!򄉾ZDT �%�g�~)�D�$�!�ؽ@K����_<��1�Ej��!�d�c�@$"���7ʨ]�HO�w��� 5�Z�(R�J+XJ�a4ݷ�y���)�Yk�B8U��|y$n��yҨN.��0��JÓ[KX��C' !�y�,Hˈq�Eˡ���0A)�!�dK2I��yIuĂ�_���F8!�$ׅR�l�zv�_:t�@���P�p2�Iݟ$��U�)�'VL$䩁>}H)rB�G:+z����5��J2��ezFj�W��X�?)�Tc��s�' vX�w'�(��`�Z�t���'O��	5tXӧ�9O�	�ÿi�`]�d��Q��5Jq�ڦ>��'�J�'��zJ��M|�%b�����a!V�jŐ�b��[#(�'�(��v��y舭~�X�����Zm0��<Ʉ�H��H�dR�=}bn�~��'6�Vd�b�y �H��8IR�,}r��&�蟔`�wB�}�*��6
�jD0f�O� �7�>���>�PD�$Ǧ9��b�8
H���q�
�.�P�"�<v�V���a�O��:v��P�2��l=Sđ�����:��#}*��G3a����{��!rh� o����N�R�X��>)�g�]~��	h�O(�e:��1_�p�+N�+}�J��r \��>[p��S��'X��3�'pV؈�85�8����#G��;��P���$���(5�7��j�"<�!�8c�"=Z窞����p5��2J���'��'o��g~Z>7�	!t� �2���6� ��J� ���Z�IU���	��nb4ᤠ]W�P��DΛ1$�!�dʵv��)C@��J�#d��^l!�D�\���$dԯM��Q��F��`!�d� 	y\$�!�L�An����U!��MR��S�#��q�兏ah!��ٽM�NQ��Hw ��A��
/!��%����o���bw!$I$!��4�5Y�a���Ua!�&
!���48*49j��.C���{d��(*�!�DP�F��3�ͦz+r���N2!�d��S� ��BF �N}�N�;?P!���z�UZ��v�F)*��46!�M�L6�##DI�)��{2��u/�O�x�N�O�~���	C.���Ŏ��l�ThśmG�6���% �O%�~�7E¤f߄�k�^z�&���lɍA/ܼ����<t8����@;$Ѯ���C��k"Bi�`��8+Z�SB"@�Q�4��g���Bpi�#�H�\cFn4DB��#�	C�I&����J,J�0IX�Ar����&D�(j��+� 	yc"�x<����?D����	
��� �د x$�#C?D��@���uS��B��IHe�8D��%�]�)Z��RO�*YR�"�L6D��[��U�A�wj�8^]�k0D�9qEF�@*�;B�dR��/D�t��+�K �a��:2T��C:D�x����!�����CP3a�P�+T$4D�p6���1�¥j���:7�. �@�3D��ۡex�xHb�@���҅2D�@���N�-: ��@R1��)҅-D�����S�|.��	O���C�8D�� 2!��	���l�r ǟr0�Y"O�0�� 8Z�x��.��v�ik"ON�7"JBƸ���� ,`�$r�"O���G�t�JHc�OY�@�d"OPh��J~eb5�V�
�};��I�"OĘۢ"�������A�g�q#�"O��!�E�_n�H+�V.h"�0�"O:�%@�60���7H�^8fIq`"OV�����$�C�	ҖYC�"O��@!j��l�W ^�Z�(���"O,����*g�rp���
Ę�s"OP��g�ZU7��R!Hٚ~��8W"O�u��� .�X�u��C��U�"Oހ��%UP9N�p֎�\�U"O���N�'
@YS��1*[��c"O0�R҆�6r���p�k?t����%"O�|���	�Q%�ئ�=;����'{�@�5�:9<ܐR&� ![�:�'t����>J㸬�1��!�L�p�'����E��# ѱ��ǆ�|ܒ�'�,�Y�G��� C�45���';��F)ș#�r�Q0gW#:4����'�p��FDQ~a!#���5e����'�� *�e��U�:���c@�`vU+�'�qa��2��)\{@Q�'�h3�����ѱ+R$uP�b�'�DQzc/�qFq��E$mä��';�PbeE�������=]<�)3�'&>�C��~N�R�N$S��� �'�5F��e��3񅕩��x��'x��lԻ��pD�)�(4��'����2�C�2F>��,�4$�|���'���ݩ04y�u$��2n\��'�p���[���!��ނ�nT(�'�4U 2�SM���Beą��@��
�'���'H =����bK X�]�	�'��}���!P�J5A�����	�'�@*Fō�N{�r@�q&���'���7j��R��h�⛁�����'X�RP�S�l�\ѡb�E�VOz���'�H��IGj���@h�6�i�'�2�`�r�$���E�=�{�'p 9b�f�X��*���"ی���'����ǙD�+�
���D��'��Ѩ�(��I���Í�� 8�=��'���+��̖8���fɋ&�D���'��Qٔ��y\��T�؁��Iy�'l9*G �=״I�$jȟx�Y�	�'{�M�����ݐ� �y~r\��'
Rd�@�X�-U�@�n���2	�'���
�`��!��! էclq�'l�!��	�)^���G"��^��
�'�܉A
���Б �.Vt�
�'���P��iL�X9r�\�-�:y
�'�l��F#�>�p,��M�?�(��'yL��B��?$�l�U�6T� ��'�4ӗI]=l��QS�N;c7��x�'?���#�_Hhv�&r���'����ǀfk�|�$%�V�p
�'\ƈrP X�~�{e�ۧ�j(�'�Zmð�֪S����ShןM�hR�'��4�k`��ђ�BF5�~���'�"Ȃ�lD>0,-e�6Brkj�<�CSi���\�ր�GD),�!�� ���R?	���ө'>]��p"O6�q
�!�ڌ;0KV##71�p"O2]�Q v�zm��d�6�$�2"ODŪu(ܟ}�<��7`�
��"O\}�#F�d@���-&Z�����"O<��tlݽ� U�Q�2��a"O�5�բO�JӤ�c�,P'3�Dq��"O�=3T�ՈG���-�svZ(��"Oͣ�!�J
�5���ǋҤ��"Ot���g�
�*t"ה#|��"O��9���(P��e��;#�\(he"Ox�ZwE��.�Z0�Ɔ>1zj�	�"O�Գ��Гo�0 �ŞeB-��"O ����+&�4�#�-XT챊�'q&�6��*Y�����+�(6�r\��'Z��MR#	�1A&�	8vV�\��'�~5�1�P�&����pjS3l�� �'0�W�<'$���fޒ*�j�"<D�@�	.*eHIb��[(Ua�m���;D�(�_{�,�cE�y{�\� A�i�<1�@-sc̤���6�2=�m�<����!I���g�ܭm=@T�0��i�<!mY4st�(#0#ǭ8԰٠!�\�<YeC�"��Z']hY�a�Y�<��X��ȨH�H���!�V�<�KҴF�*�ye �{�L���Q�<��_UU.m˗�ͬYY��JvQ�<V����8�!�
%z����1	�b�<!4H���Q`3)�ja��Z���[�<ŧ��j��8K�1/tz4[� C�<�W�״_䥫2 �47��3R��c�<	�N@�R�hP�P
D�<j�aS^�<)Ɂ�:��#� �Bͨ��!�W�<"�Z���aVpA��L�<2�M�p����)�p��]` ,o�<��샆^Ж{�lՓp�zp#�j�<aNTYL�e��J��5�αp䨈f�<� �Ynd�"��	d�Bi�qN\J�<��,�#G��J��E�KM��J�D�<a�'�'IBY��� ��ܳ �E�<����:��=�r�"we*�����f�<�E�?�,�eGZVļ�ňMd�<����,I��}*��D-K�lip�\�<i�a_�{<�U�A�^&n��5��]o�<�Rc1.��pև��3lȫ#I�n�<����!rd
�i j��3A�h�<!b �ؘ�)WJ¡ `����f�<���,3*��S(��
�kѢ^f�<1B�
8RC��9�8ظ���d�<Y"GŤFʤ5�� ٔ4�$T
�bX�<�4��<y^艋��G	7&XM*f�^�<1�P�yI
(0g"��u(��9e��O�<1�`!=`�y�Đ�C�f��w��R�<)�J۩;�8�&�ѾŮ�!�g�M�<�����o�4���`�����A��^o�<��A�*?Ǥ����ԝu���� ��C�<��)5n,�d��Z1}	�.�I�<@
�< 5���-�ʡR��a�<�Ef�JP��9��
�ok�l���G`�<q�E�
�8�aB���}`9� �]�<��`�6jE7J/$=��I�ʓ]�<��)Q\��	�D�,;�v��EQ�<���F�;Qr���F�`�A�N�<�u!�`��{d�WMfP�+��Jv�<� ��i	ND�N�j�c�s�L�	1"O�����F������N}�H�"O������*�a�XNS��s�"O:����f�����^�Zj�i"O��sG��>|��0hm��C�A!V"O`x���P�Jȑ*.F���x0��b�<)�_/vJ��ؑF?&D�d��\�<��J$� �k��2YX��gl�P�<Q��-d�Q������mLh�<���&,��Lk�k�?+��8�id�<�!�(X#昨��^�q\����Wu�<��K�ϊ	�!��N��6�M�<��F�-Z;V��Q�71��`���	r�<Q�I�1s�r��ҵ�T��QL�n�<Y�Dދ�����^3��y�$�v�<	�j��f�}sN�/��Y� �s�<��bTf֞|� /[�Y� ��An�<��-T��Ո�-��-	t� ��[i�<�'��$k�� �w��^��!�ү]_�<9w���Y�>E8ѭ�oP����N�E�<Q��Gg^Z�!�)s��P~�<٥Ĕ�vգʐ�U�u�U��d�<�&�#\A��G9y��k�F�]�<a�5X� ��͎�F�@4k��[�<1�M��*��"�7��m���LV�<�6bϋ>�LZ�C�0^8�h�*W�<��x%�ջ%,E*dGX8[�AUL�<)�U55�$b��Ȯ:�\�*�!�D�<��j_�~g��j���p���j�h\e�<!��?2��<0ƣ�/$(��e�<��+��?C�A�NJ�D��yr���a�<����B��Q���RU��R[�<A�T8%�4q���K��l�g�DZ�<�҂��m� zg���R���E[�<QQ���N���Su�I I[@�<QF��'Im2l�/��t�`eE�<�S&X�-�.��%Cށ� �j���w�<���<o�t<8��e榍jr��s�<a��ٸd�~�C����ț��I�<1@nߒKQH��6H�==X�)�G�<�R'��&À�`	�:3�d8�"h�D�<�&�>V����kǁh�di��V�<�F��)-wF���.�#���ڡ��Q�<��f��(*q�նzd�ijW�x�<9�O;ot�5��/�+�L���dt�<�G�,Q� ��# �hTZ��@��K�<�$*��V�P(&�V"	�0虧*�a�<A ���'c�Y�t$S:7([B�\�<u���n�����A\䵂���Y�<Irm��t�|��a�!�fd��T�<���B)	2f��F bEl-r�e[�<y��9R�px�� 4���UW�<�S��>?�J�##N�5!(h��U�<&��7q�Xp&k���Ш�bLDN�<!@dU%D�f�Y'e�"x�p%��G�<*KW����d�p�IX2�N�<9�M�P��ƌ��X�@i���L�f�4���a΁O��-j:41�#!>��	�0� C�#݌�X��� �!�DE�Q�<Q��Z*	��	Q�LA!�('&}�T(]?A�J��e�p�!��=_�Pԙu��
��`�vc�(E!�Ğ�8�ؕ��J�s���V�GH!��W�U�V� 3�Q"����LK�6O!��

 ��� !��G��{@�K�U�!�� t��Ui׆
Cl1��υ�F("O>�q���mS�\�@#c�Vy"O�|k��ң<�l� ���m����"Oy����1�m��bs��"O@ܳ�A>8ٚ���i׎Gj��!�"O佀�N�<U����A��?S�� �"O�]:$o�,Da�PB�OC<6��K"O���G�E#�hjF�N��Y�$"O��K�䓼$�A��K�	�N��W"O�<*t�C�\�Lta��(.U�"Oz�%,ω�h0���`p�,�"O�y vk��Z�T�Xe	.O�؋�"OV���gM9@)�B�~LR�r"O�y
2��Vq���� �<2���"Ohd�W�?"�*\1�F
yf�C�"O1ЕB�@�P�$�أ)<�g"O$Ę�`U����� @�5B�!��"O�|�f���S��PK�I�t���څ"O�)�r�TȈ�E~|��;A(�(�y"Z$O��*��4)FȈxѦ�*�y�M`��]X'`�(��z�ጦ�y"�Ѧ=�b@�а��C�$.OD���'�^��A(_3tP phi�*��(�'݌�#IS 5�E�dA_y�d(�'���x*ѝ����������'�H���Ď*$��8�3ޛ�ź�'F���!'��3�l���'}X����2�8�@���'�d�Â�5rB���y��X��'�li A1LC���Fd�g�Z��	�'�^�e�H0}�R�2�e['1�y�'̵ T���*�R�@�+C@�k�'؎y�&錦O����:�
�';@ �3'��O�� ������'=�Ԃg�Q��, �š�>^	�'��r�E$dX1��J'6,�j
�'_b��F��
R�0�i�nK-;'�T��'s�1`ˉ"�Z��wc��}/PtQ�'	��ˇ
\�nC� �&bL��. �	�'����#�Z9�:]I�B�9�d���'��4��,6�� w�X�2Nx���')6��j� taR�j�/�)ܮHs�'� Ȧ#�/B+�I���K$#�H�3�'S���]:&�U���,YѸ���'�|��kV�}.�d�i.y܀�'d��
�#,E<acB�~���P
�'�I���3�D���=	N&���'[`R�cCU�nx�5K��D��'Z��a0E���22n�)7�J�Z�'�6�kU��
s���� �N���'�8i"O��y�bl���VΉ��'F��ەÔ�9Yhݢ2��(�0\)�'�%�ҭ^5I�@RBJ��	C�y��'b�٪B�6�q%kȤ����
�'��)�'�2K ��#
Υ";���
�'��$�!x��8�J�J���,D���Չ�1����D��"@a�r�,D��#��I13���`C!�=Z��r�7D�" �0u��]{��܈aø8�)9D�h����!,���'AZ�x�J�hS$;D�`����J��,{���t lr�4D���@�J�	��"���d,���wF.D��C��ʡA_ �(�ǆ!t6�ے�'D����'��I��ѳ|W�88��!D�� ¬��ʕ�q�����b�2&����"O4|�t'�/�xȳ�Ύ�$�tԊV"O�} �R}l�RÔ�E����"O^��@V+i.���a�+NYa"O��[��U�q���BRJ&sH
�J�"OTt���=b��G�y�t�Z�"O��C�M�^�X��Ѯ%��!��"O� c� :ZC�4�
�$��@�"Oډau�мT�U�'_�D��<
"Ob%��Jϥ`p��˓�L܈`�F"O�t B"�1-ܲ �"�\�t��"O�/�VHxy���7{�ૂ"Ob��b�-v� 3Ҩ����yr"O��w��+d��Lp��O�'+p��"O�ј��5z�ux�,CY��9�"O�M`f�ǦGK|8��e�!}10l¦"O�}���9==�T�"*ݺ+��!�"O�,���֧j��I�6�E�?z���"O��Z�g1A����`)�c<�P"O��C��w����a)�
�Ȋ�"OH��r,�Z�3鈾)�ε�F"Oz0���#��(R�֮t��� "O� ��7^N�#4�C�C���X�"O���G������?���2"O���Я��=\(4�w�ثCU$�(V"O�!��6?8�@�	߬CmN� $"Oe�PHP��͒`IP�� RQ"O>�1����a��jڴ{��(b"O&D:��u�D8"�
�/�"YA"OJ]{7B�;xj�eab/t�%H�"O���R�ԙS�<m���?�4e:�"O�:Ү��\���fծ	xt"O(�ӎ�~���:�KƑ�2��"O�ܡ$!��0�T+�+�
�B"O0� �X.G6z�6����LX�"O���'�	�j��pQD�U�Q8�a��"O��1�ǩ=-��30�Q880>�"O\,�d�ѩ��B���E��ɳ"O�p@6N������/n��q�"O|�x�e��N]y��ݥ.h��2�"O��S�g
�y�� ظ5(����"O��37�&�F�)tƛ�`!V|�7"O$A�O۟y�P�ا��\��Q��"O΁���:�$���*����"OfM��I(J�T(���ۭؔ�I�"O���Ǥ��;u��  8�!�"Ot����i�J�	4��~h("O�����ڬ4��B7�65����"O䔚�H��>�1����I��"Oxe��&
�M��]sU
�&�� KQ"O����ur<@U��&"���"O�L���z*�]8�A����$��"Od�g�!ll�9�Ȧ\�A"O�T�eFi�tls�Ŵu�b��"OVS��tzB�1h�`�q�B_n�<�*�
 ��d�mw�h�&CR^�<�埁#S&�I�����yӖb�V�<����0���bM,a���4�Q�<"�M77	���b�&	��5f�_R�<���_�W��mx0��"1x�8��X�<yT	�N�&Y`*� } �(U��J�<Q���:-�H�=���(s/I�<����	����J��u�����C�<q�l��H��S��P�bW/�E�<� n��M�~�x��S?�zP;""O,�"��-��=k��/~����"O��B���H�!�Ǐ	���uXq"O�8X�N+/��@��7븘X�"O4Y� )LF�j%�`Ŋj.d�AB"O�x @��)-~鋴�4q�d��"O�%p#�˞PY�R�4A� `��"O��1"/Y�&m�e���
��"O��� N:��@��K� ���[4"OV59b'�\X�#˓�6��"O1tK�~K�)�g��v5���R"O:P��� �� �Þ41��A0"Op%S�� 
W|�2'W4$�U�5"Or�������@�6M|�y�"O��Q�Z�S �9S�؉j~��#"O61y�D2L�~l�GoʻB��M8�"O��$�Z�1��Er�oS�\$��"O��,m�2� 7E�D��y'�yR�D�@�Ԡi�N��0⡳���5�y�GՇd�~���)�� 2���?�y����.d%�B��-;V�q� I.�y�oYd�)@3I�5�`i��L�,�ykC�q���%*��)��$����y⌘36����a΀(��Ms�ת�yr�V�:��Љ�l�'.���ō�yB�O�"�Ԍȓ�B�+o8e��e��y�?R�(Kv��:"�ԐѢ&]��yR���>�Ժd�ZA\�B�(�y"N��5�&�Bt�ѤO+0Q��\%�yR���h�J�Z
����o�!�y�j4Cu�@s�я�(y����y�Z�z�\-K#f�7ynx"�T��y���F��dְ#	�O��y�H�q��UI�"��Y޶m(Q�I��y���\h��Rnb$�'�?�yR�>2l�}����:�l
'薥�yB-uGRI�_'�-�u����y���V��˓6G)n�ě�y��2<�s@* �z�tȅ�ܮ�y"F�M��(`��=�>�u/�y�]�?t��'�W�f޺|Yuf��y��֐*`����N.az���yr�ӸhA�0���H4`�(�J̱�y��b~P*�ǛA~����*ِ�y��Y�!S��jӢN�n�Q#_
�y2�-UT�l\$`.����yB!��:Q��r��H���)�HZ�'�D�d�MS8(@���E��0�
�'�|�(P��4B�}�
�U;6M�
�'94" *=|SX4,N�;C�{�'i�a��+^�uJ�)��KL�H�'iహ�.U�Vˤ��ʒ�M��p�'��,qh�<-"�j��?Jk~a�	�'۠L�	�
�xZ�ɽ{ �\z	�' �u"��(�fq�) �ut�]h
�'��T36&ؑ�fX�v�,t�V�s�'�4�r�����1�J�	,���'P��yc�8�X��"ӫ�X)�'�HU��-G�)!�����	�'b��z�n�`(Pj7AJ�(�'`uk6�ہR������9jgp9�{r��A8v���hN�#��q�ac;�dU.FВ`��6x
���e�!�M0���
��K�$wB�h�H��Y�!��z��MxC'Y�%s�<C1���!�� J݉@K����Z���3o�q�"O��x�HΏ
4���f�HjjH;�"OsW'�[@�q�'eK&PO���"O�IQ�&lR�Q�� 1H��"O�A�6�.>�ӗcĴhKN�)'"O�$煎��ةX��޲���q"O�� �O�+�ȑ�P���8���V"ORY���R�84`��[�E��iS�"O� ����7iVm�4R��H�)D� �b痴�� �ǣQ��0Ҁe'D����'�,�s�8�h�@�,*D�\sC��C�D�� �3�NX+w%&D���Э��xP�Po�v�,� �!1D�t�塜�fyF�
 ��/$��ي�5D�\JCn�%~��j���Ks����.D��4�]/	-} �h1 e�v(+D�8�e*߶E�"��F�X!qE��>D��S���%]��l�ehX�*��Db� 'D��+�HG�$�d�gF�BS^��F�%D���&��HF�Z���%B)0}*�#D�(�`�Ǭt��t;��R�+�.���"D� ��.��+��h�A� °�B&?D�x�S��!1%��"f�b��kУ/D���t�Q
n�i��m�8���k�E2D�����9S�C�/!3[jL+�e/D��
+��Q��}��W�\,��.D����žKn4h�&�޸[�H|��-D����cՊFΖ)��0c'2�7�*D�1��/8M��sO�$|8g�=D����dLT)|�D�"Y�șS�6D�`1(G�"��c�.����+5D�pp5F����24�t��9�"
(D�ܫFŃ5[ڼ�p�,��!:�E1D��K5M�*IEBt�"�M6��cb
2D�l��Gh,�3�➙?��%{��"D��"E匆^��H��C�B�刡�"D�8��R�$��	�T��3v��,3��?D�t���:v�bq8��B���:F�?D�T�*��/�8I超�;c��"D�Dp�)/ !ib'��
�2!J�,D�����P 7j��Y�>P�M�*D��`�)��%�$�&��L��XX�&D�����!vPa!��${Z ��2D�����2t���ˡ��!�X �v�1D��Y<-U�4J�i"7䝢�I.D��ٱ��[�5�����z�'�LEE$�9VӺI r�hd�h�'8�+T	�M� �i�y����'Ѭ�8f��#����m��E{�'��Xi/f��};�o��i��S�'7ҍ`�O �h@�����W�n�i	�'�ع+�/z)H3aWTH�t��ǁ`�<1edR4(�4��M%(E�h���[B�<���'3�A��oE">U �a�^A�<�]0�T)��K�(5 ���n{�<iA%�a�py�`
$@MTP����z�<�@ܭ@	p�`�{{���Nr�<���4��+���J]^�ؐFi�<1!�'k��5�҅��o�lp����c�<1�j�&��2��֖#"��Q�DOb�<��C�Z)fl	����&��TKLF�<�C�3�B�	�Έp�n�sX~�<Ƀ�6{�tt��+@��СEm	p�<��:q=F��m&��{SNG�<� ����O�uX��GS�.��S�"O��bMCFV�cl�6c?��C"Ox@�#���pl�˘�z;�S�"O��Ӂf���8�c��4��c�"O�yAV�#/+�}꤃/�$U�"O�@b`7B	��"_�kL� q"O�j�@ىi.�J�_L``�2�"O��4�x�a�>vI����"OR�Cb�K�Ys&mi�G��}	@|"Oh�bI�[�H��p'�:I��:�"O�L��Dn��J )��X���"O�y���I'�&A��^�V�"�"O�A
���q�0BQ�=�#�"O 8b�.�7�$��φ,�`�!�"O.�p����"���JЭ����Q�"O�y���`s4(!����4�m�@"O�I��Õ]=*9��l��!,�$�r"Odɢ�Q�k��H�ī�B��"Oʽy	�)�գ���m�(	p"O�}H7)O�i�����.��]U����"O��h�V6!�|XEN�wSޝ�T"O,E�j�t��u�v-�{a�,�7"O��0��Һ+�@�0�*N�OAN�"�"OJ!��십1|��Cu*J8,B��"OvY�3�φa�$��	�%K�LP�"OĜy����2B��sf>���U"Ov-��BK�-�ԓ���<u�t�"O�̓�d;t�(�b1!��*�b�37"O����L���1�OPz��u"Or��3-M lZR�<*s�(w"O��G6>�hAaď�5=pBA�"OЁ:vn۠"��}A��E9<Y�{b"Oؑ"tB ;�&�hN��+�"O��! jM!�f�P���D� `"OLA�A�X,h�X�#�XX0>=
�"O�5��ĹkS0@�G�C�*��-��"O�yb���l�� �*C�:��"O�Y�։C�6V�ձGf_�z�Jls�"O U��'6!?��&R;$�����"O�(�A蝠$m�!�6ƚ���"OL��P�۰1����&D^y�Y"O.i� �ğ
����5b͟~9�A3"O�4��mͫq�j�Y4A�����8�"O��r�	�l23.�z^�\xE"Ob�w��$����'�C�KpV��"OJ5�HR'b^���l�8jn��"O (Ө_�0^�  N<R0�@a"O��ӷ�̦:�"$͹3V��#�"O�x�BǠ},2]Ð"�E@=!"O�9�aD)
�l�����B0�Js�'!�Dޑ82�\q�o��}w��2 �1S�!���6���AOP0(�^����7!�((~@ы�f�2z�8���˟�<!��DP�3�M��~�H$�Ы�4G`!�$P��6�`a*H�]ht���C� �!�D�*�nI�&��1Kva1��B��!�d���c¦IV5�r!U6�!�޺j�����&+\IufF�v}!�d�& �d���V6}22`��C�k����,�&\i��㦥�V�zC�~z֭cM��#�e�B)R\C�ɑ���&�>a�[v�όk�<C�I�z
$�j�R��LZ#�C�ILH�mr@��-q��u�ֽ
#�B�)� ��W�u���1����K>��z6"O�#d̹MX���NJP�#"O���F6*?4d� d� �F|��"O�!kA�+6�J�`�`� ���Z�"O"%���B�^Vf�5	P(E����"O���@抍:�5��
��-��d[�"Obd��/��.(��a5I]x���"O�U�'ț�?j�2���#UZ pD"O���f!�j��9
�0�`܈W"O����.�9 KP�䐬6H��2A"O� "&2y.�(�`��KKh�T"O�����)W/���1G|S�"O�� �DW���2]/6P���$"O���/�?����T9MA���&"O4�� �9#.<�s�.DE��"OR-�f��@��U9u"��T��Q�"Ov�Q�.L5�ƘkBBԡj�YD"O<�Ä� 2�.��e G
g(P6"O ��wF��U'Ơ���74U&���"O�yr�	P�ĸ��B�2$Vr1�"OJT�T%U2-�B��!�|Y̊�"O yp�!ž/^�[Ak
)G�<z"O| ��	9¦���A�x`����"O~$�AӚ,xB���˞'^h� �6"O�T�tEϒP����`�����
70!򤅺^�6��FjҠT��Y�Iц&J!�Dן$��:�kԆ��LP��[�I!�d"oy(h�L�)v�~����!�� �6�"�ժQI�E�p�N�:z!�d���d�A��Q	v2���AN�;a!�X�B��qą�5r�L��W���xD!�D
>o�DE���TJ����F �:e�!��/>�&����У6���� E޴t�!�$�|�6hQfY+�8����Ԟ �!�$��w�PAܽ��L��&P8%3!򤚤��( ���'�&���!�Ě2&�,9IF�1��za�{!�K�����fH�>�8�)q��>!�D���R��&C��`9�PD�8&!�3o�\�[��ОJbhT!� Ly�!�$�>8ș��_�-U�t��Oܸ�!�@~� �T�4n�}��/�9�!��ԅ'��8X�
X�R.`� �_!��!>I�y��聮DK�1��@���!� 2�����L�|]L�J7o��!��T�Q,�q��C@�x��e`�-̨)�!�*M�ԭ�#J �T� rMF�K�!��.c���9��28���9��X�!�$�?#�h����%�0��Z�!�Bs��5�e��:�4dS�(iC!�D7y��)0� s��I�!�.})!�$�A�����F�*�:X����]!�N(d��"s /��5���x�!�$�5��\X� ��-������ұ!�!�V ���E��,UÀy�@�� �!�۔a��ǈ�M*� ��zw!��b`f����]�Vt������!��^
mb©׉��:7ϑ)R�!�Ūt�E�У
8�T=��.R;M�!�_�5&�9ч�?a��1����Xu!����c�S(�r��'Ո	�!���KJ� �4���BGU
�!�DԣC��� �/F) �F)q�(��m!��1I�By��j�)�$�b&X�z�!�� }��*�9Y�V���C~�ӷ"O8�;,�gx>��CM�o8�"O(���T�Q�:$)��jPp�`"Oh�9�.X�w*� ��L��p4�1D"Ol]xf64ltY�'ꄣ1X�y��"O�!h���2Sf�P0K/��\��"O~x	%Ɔ3�b��0��r�����"O�m��b(/�� �.�.+��i��"O�@�ƕ�S#���4�R}��"O6��� @.�!Ћ�T���� "O�q���Y��%��{�v��!"O�`�CD�sq��'k^j1l@��"O`��ch\�%��٪U��( 
1)S"O��J�@��rEQ�ퟩW��)"O6HcW͙6GU��(���~*N��d"OZ9��)_&v�xX���S�zN0�"O���Q�R(��|�F�	$s0ࣆ"OfuR��C�f�� "�ֲ5X��"O�x	��3|ߺ���"��^��)s�"O$ir#�B1
S*5�W� 1|�V"O��a �--�8` ׯZ�#l�Iiv"OH���V#x8ڔbsOԂs�����"O� *�,��j�H5�m�V����5"O٪Wϖ�8DyB,޻ �d)Ӧ"Ox��v��)A����
[z�ҁ5"Ot����;h�(�UJ�W��HB"OxU3��V*K��ڢ��
�&M�b"On�sE
6��,b%H��j�D$�b"O6�Y��ZR*F���FD�/�F�xW"OD�����'O1U_|��d"OZe�ăWe�`Q��Krx��"O@��Ƈ��xݲ���=c��{"O�����^)T<��R�OF��T� "OΘP�S�f�Z����-T��E"OR\�D-Ʀ4�D�4"��K*�0E"O�l�g��EO2�d��TB `�"O�M�Bm��-��b���'F/Y��"Oh�	R�\/	�0` c�]<b�F5�!"O<���ȷX���D���G���"O���\$d��
,e *E�7"O���P
����L�J�uڣ"O8�����l��v�@S���IB"OB�sL�E�f��7��!<{�H#"OH�X�NεHz y��Ι<onXa@"OΌ�Q��0�vQ���%cD�2�"O�)�D�[^�6xz��_8]hX�"O��a�%�| ��PNp!�6"Oh
��36�X|X���<f9�"O�5
2�� XϘ��ӤgF+M�j�<�$(�\�b����fP��Ua�<1���	��ذ��L?ĸ)TE�`�<!o��$�1 �> ��B �SY�<�R���=b�5�ùS:�	R���R�<��GLTA���2K��0@�q5��c�<��mB[�,9sra՗>vDj4�HX�<a �I2Vt�$�Ӭ]�e{z|�O�T�<�Ӊ�:w�8�A��Y�����&M�<��M��<�F�a�ܸ��m�*�L�<��Ҳ".�1�\� ��B�<�����H*V�+���+`iv���PH�<	TB�+f:r�#S�R�l�j���"D�R�ͨ����ųs����
?D�t ���_�eG�3pp4�J�<D��;R �M��b��%>�@ţA�8D�� &��&k�!�b-�D�)���X�"Or�hkA�cPc���!GȽi"OZ!�A�A%n<t�ǲY�`��#"O��h%�-*(��+�zx!�"Ov�ҧ�ϵdec�6C8�y"OyA�-�vi�����*In@�Qf"O��Ӧ	�P����{en���"O��a�
3���K���5��� �"OPQ�@�G{THi�Ӏ�q�"�*�"O.̡3�ݔP�4���@Cj�VY��"O�isq,+]��� �~�J�A"O<43��- '� 0FF
	s�e�'"OJ=�.w[B�BV$G�Eh�%��"Of�c��B9Y`�"�*N�x+�"Of��f��� �� 
=c<L�ɠ"O�I;D��>�	q@�w��xv"Of��Ϟ�E��]�g/S&��h�!"O,�;��ǐw9�B��:�ؙ�"Oər��)h��AIÈ�'#W�\��"O\�c0�  �z0��狮/Q�� "OH�X��uj�gAS 7M̑ �"O�I��Y�>34��-��h��"OZ��g���� �Mӳz����"O
�#`�ޯBXP�3�T,y<ht"O4����X�c�W�t��E+@"O�<Zb���[[���f�5�$��"O� ��g��[�0�0�.N6|��A�"O�i���N&pm��;�nX�kD�Yp"O�)���ωh�A#�E*J-�"O�P� ��?|��ZdI�s>NQj�"O��o׻u?�xB���2�c�"OAI��,�d):��D�]��]��"O(ȚuF�E7&�	�"7Dά H@"Op�sSa̳@�ļ�ËE��!i�"Oٴ�_�,���bCLl��@I�"ONP�NH'X��YD��\�� �A"O�;��L���\��L�Kf�e��"O�X��B��%� BL�JE���S"Oօ�g#� ��3���3P]��cg"O(f�M�xv���H�wLH�c�"Oʍ
��9�0=�F��#9��+�"O���(X�z��5�7�S�9��t�"O\8+G��J�����H�=_�����"O���aGL�S9�7�V2\42�"O��`�CF�H�&�<28Y�4"O� p�S_��D��G׸�[t"O�|���h����v�I�Ҩ3�"OcRh�/q�]���Y�(8��"O:H�F+�f���HE�T$|����a"O�Ȱ�i&PY��㛱c�^��"O���B�<2����g@Q@**��g"O~MQ��H�0<�ms��ݦM��	�"Onx�ԀU��� ��k,�A"Op����I�+|��r� �*���s�*O�PBn�PmF9��
+m����'h,��B�K촃r�\�Yк�#�';���e)׃A5vTSG��ڢ�B�'��Ib��F#�\Q@�v�2� �'x�Y������ᝯq�>D

�'�HAcWnɰM>�P"��@2�}�	�'О�#$��[v&MR��ә�8<�	�'mD��͎�L���M��u��'�V�[q�Q�������$Z��'��q�B�'�(S7���g�С���� f ��%|�)�h��K�T� �"O��0#�>07>d��眑	�p�۲"OF��N�}� �K�դj�
a�"OA�KX5N(d���Ҕp�@���"O�4�dB�p�5�P莛/�H�"OF�$N�#G�L�`F�	�d��"Oj���ː�_U2!��>�X�(1"O���c�TR��A��ѹ�P��E"O�T�ե�# ^} f������y�� 	]�%'�ϡ�H��b���y2��JP�Ƥ���b�rܥ�y"��F9
�2-к!��f��y�F],LT+uڵ��%�Q���yB�.`ysFj��P�ܐ��@]>�y��� [�`ȴ �D{��i׀Z+�y�M� �nE e��,,�t1���;�y���p
�����9i*�S��L��y���&6�>��W�O0 ��u�@̓�y2��jF8PjQ$?n�. bM���y2�
�M6�%��jA�\#�En^?�y�˔p��� )��DtT� ���y"#��j��'
$7+��
e�9�y�'��BA.ݰYr4��y��e���9����7��@e�*�y�-T�>�����=B�p�A��ކ�y"b��a��QrWD7ӚaKׇ��y�	�\j1�6���6��E���y"뚲Y��A�*3AD�K����y#B�bV)B�Z:v���y'$����O��L}F�A�����ybN��ZH1��O!N<�p����yRf��v�iւ�
z��)�I��y�����<`�N��kΤ�q�)"�y��� �^����F�3���S�L�v�<�N�E������Osޞ��AE�F�<�&��#ETc�ʫ%����JB�<9fT0,����o�<jLy"��d�<Aw!�!Y��
bm
I��0��l�<��3U��LQ�Ǜ���&�i�<���*���Rl'�pFi�<iT�Ք����c]�~� �+Ff�a�<��gµ `h�
?�x�NVr�<Ac�U!V_�9ٓh[�� y���r�<�FD�h� ���Y�-�
���RY�<��)�,��MIv��M��,��QR�<�)J�"ٸ�*S͝:U �q��l�P�<����_�سө����H[��t�<y�e�ccz񪗨O!l\Z�0���l�<��Řha���@��((���Q�\Q�<A�M� be�����4@�z�)XL�<��,߱ }��h6��_�f�$��@�<��޺հ]�#CM�{�NEW�Q�<�%I�-�\0��1B=��N�<�1�I��x�Α?�,�#3!�D�<���]Q�$��Y� iP�[h�<��#f��"E�A�d��@A(�k�<�Gc�1���"u��Qx�}``j�<��c��s� �2�)�8/�H�Rd�IQ�<a�C�,`��h��[ )w�|"&
�R�<��䊜���SgΑ�;;,�i c�K�<���W�m:�d��X���4,�l�<���H+r��MP���/���"o�g�<Y���M�\�S�E�А��Og�<ѵ�Ű�\�7E�R���3D��e�<� �DFp�$�3�X�`�zA�0"OX�s'Z���ą�yr�H��"O<�R�i-e7¸�r╽p6�݊�"Ot�A���"0[�ؤ@x��"O��؇��%�2�e�;�� ��	ӟlqᮈ�J
�&�'3�X?�B7�O|ІY%>Rɮ�{2i�/XH
%���?)�/��Dƣ�M��9�J$U�����h>ӕ�K��q�c��V���+�#ғsfi2���s�p!�b%��Q�<���شS8���1E��~�*x�ER�ON�P���Nx����O�n��@�Ocn�BQU����J��?JM�7&U)�l�֝J��?�Bm�Y���0��%?sz,Q�@�A8�0:شl��f�i�NH˳�Ln	�y��$��q��'�v$��h�>	����<;}����O�6m��\M����V>�k�ߒ$�&���L�~�v�lڕC�xQ"�ޙ]���W���O~�Z�aפ�i�NZ^�=��A�ߦR��� ���m�(U�x;�JA���� �s�W�8C
��׃��ɠ�&��Mw��Ο�I��M��������E�<s*����V;�ؘ�d�P��~�'���)�)э#���!�
;-������T=Q���ݴo�f�|"�O6�Ώ/6����,.�����"�4�����KC:>y(�	�|��ğĺ_w�ҼihNi�Ɖ!G����
O3��� Y?L<�,`Z���TO{>=�����j���D�q�4�
e��''#a9�n�:]�N԰��N�dnZ�67Mi�$O�x �b�p�`��)J)���G�2��l��Ȧ>�sJAʟ��IT�	J��U���Bm�5TAp�As�=10�+�#��܆�I�5����`��8�d�A���!pX�h#�ii2�|�OT�$����R߶��Pk�.��1��o�R���o���T��П��I���	����I�N����TB�&<�R�I��)W��iJP ��p�a.�� K�i�<3k����f�G@A�4�Y$p��EPF�n�y�j��U@�4nYe�� )�&�
�HO\(k�'����!b(�����/[n�Y����C�0&�����\�?�O=L����|`1+�3R��Й�'�a"�L�.|���#��{����Ȑ?�~�o�^-nnyRC�-	����?1����&�
P>���-�T|�%������I�	�H�$�զ]�O�����u>e�T茭9�P�P�#��/l���+ғY*�w$[�dY�,�M�	6��{4#üu ��[$&V+�� �䄣6呫 푞 `�.�O��d�����Ij�dX�D��q�	�Y� �{���iƸ�:�)��d���.j-�"��J��Y{3�7��e�'hh7��Ol6�ކ#�l������^�d��.މ�D��ll��J���O&�d�|*d��?����M�5�ʢ6D�d��v�8h��̓�Z�
�#P��6QV�x4��-~��	�,Gy:*���it����T-^̬PC��}���B �M�gM�4vpu���@���C��`��!c����X��A*9���Ī(�BL)ôi��8x��?��iP��s���pDi4m�0q)� !H|�y2�O��)<O��4��ZR�P<������2qQN!Dz�iܰ7��O"�m���Sͺ3G�W*���u!�㎐�R@&s��'�a{B�ɰ   �   /   Ĵ���	��Z�Zvi˕.���3��H�I�
O�ظ2�x�ؠ�!ٴ�?I!�R�pi�yzvI��t���9�
��6�o�Mnڪ��=�&��9wS�5öo�F���En\?j�aDx��W\�'Vm�8V}�s�D�W����˓E[b�C���>b) �'O~Kֈ� ?���`�O�pr�狽cb*-"�K�@�Np�f�_�\�ܳݴC�=O\EA�F�u��a~bn�<#2Ӂ�N(bjraPgd�V��M����N�'�0�Gx����<�ʑ"t�����6���t�	�A���'�|b)Dm������)+U�,��钼�yB�HS�'%��Fxb��ג���E[ p�hJ��Cnu�"<1�M1�q�F� }�����W#w��`� �}�E�Oiю�$�Ҹ'�
U�7*���5��fRKn�U��4U��"<ѣJ z���ɭP�F�
$'�<#č�e%Q���"<qׁ+?���Ȋ-�v1�"�[x�AA�HSy2�Ko�'Df��?�`�ô.���OV�Qn����g�v��#<9�./�n�$���0]$伙�`�-j�΁����/�1O0�x�����ēdt�=���~Ԙ�NHk����"�F#<�Ud$�Ye� ��Ӄ1$q�"ZEw$�Ip���LrRP��i���HȜw�ĸyb����8Y�b�#hbm.O�Q��n���'�8�r��Þ�� |�	bѷbxf0 ��+.� 2�ѨW��Ey���c�'ɞ�B��J�,j�M��M
j�Ċ�'�Ρ @ ��Pv�U?@V�b��s����w"O��x�F/���	g�1g8X:Q"O�%Q�KP�L���h��C[p09�"O�]# ��+:��H��cLԒ��3�y�f	�%��!Y~���� 	ϐ�ybK� D5���<C:�����?�y�oY�y��{���$?̜9�g�V�yb�^<�u���H�4
V��� �y�f� f��m�p��!)�����?�y���]^�0�����@����yb!������*��)���8�y�`�l `9�P���=`��I"�yb�ϬcR�z�KǊ���D�G�yRI͏P�i0�.Ѻ=n|�1����y����JbT)Ċ�:.��s���yr$�U�r�@bC�X8����0�y�#^�s�����)Ѝh�2��¬��y�
C5_&���&W�bZ��ŊO3�yB���oc�i(�i��`�������y���5C�K    �    �  �  C!  �'  �(   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic�Iz�����$qX���b;y� ��bM��!�D�<�8�3'���|pR
қ&�"�S��M��޻L y;$��$�a��H�v�<I�l�H���ƍY�qId����Φ�?�Pi��1i4.��0��ې�	Z6r�	Q�@|qJ��""�'��#*1Q�h\��LՈK��4�é5<Pҋ=LT��`�'j\��6�^�)>@$"adXf�����"b�Թpueĝ0�|�J@��P�T	���吠p�b�i�Y�@��B�I�<-Z�����-@6 �e\���ת�X��� �h2~���Ñ�-�g?���T�Sֱ₨�nFH��Ql�<� l��R����უ4�J�c�l]K@��(A&�+<�>9H��T6J�Ԯ���O���F&>����M��RQ�Q�C�'��H�U"J�h�!��!^���&�r��A��*�?(4r�Q Q?��~��O�5��Y��fK�\k����'W�2��:~��e�go�O��,Sw�~Z��^=HU0��"IM|��i"h�F�<a�&%^ؓ�-��S(�ّ�B�!V�PT�iYrX;�J�=i��D���O>�1j�3',t�����m���"O�ȹ �٬i�|@��eP�c��u��i��̘���o��8¦M���2�4�^2��"|��w �@]b��ɬ<���	�-V�t~^	б���4|���CU��<8-][*XJG�'����G�1eO(8Rf`��,�@�!���x��<�ǃ��#J�Qr���j�3� N�р	á&~��W�[=l�`\��"O&hɢ��77�Ji�0���+ak��lZ|�zw���D 	���O?�I�g�xP�E�x�P���Ğ>�XC�ɼ����*�8 J�N�=s�P���+M!�xr���i��1��|�'S<E��OQnJDy�F]2eb�l�d��f��r ��K�$Ԡ�/��;K����+74��`�OjO5���.�j�{W :ғBPn1�#��g��?!4bZ�s��!�nF�Y�4����'D���p��H�H�q/E�a��a�� g�|��$]wRU&�"~:��L��x����<�xً�EII�<��m�8MA��V:&l��B�D�I�l�Lل�	:Z�Piaa�,�����9 "B�+j�"2E��A��Թ0���X�B�	4Q�1p� x��@�FUvszC�	�4�����t�v��G�0C�I�? ���_��$,;���|��C䉡���)ʎFm��C"�Q�~�B�>T� �MW�g�D�������B�*2��<2N9s����q+��tHHB�I�̞<P����/g,��7MO�)B�	��9Ȥ/_�=K�a�$�?o��B�I!;�3F9��*Ԧ_�QZ�B�e6�����=|��a'��B�Iy��y����sސ��'��A�B��M����B�_�eP�c���<)HB�IB��8e��-��a#`@p�B�:?��q@��� ���Ώ��B��s��ˁ�7��*�l�4=B�	�ba�d�rǄ�0+0���$<l��B�� Q���p�I-��1���^��C�-�R�A�b21԰�p��ޤ��C�ɋu�)AS��T���d�c�C�ɸn-�Q���"0��C�@.*B�I�AG�آ����0@�ek�M��B�I:�E��N�=IX@��@#!�B�ɁO?��zu�Lr�*Р��U�\�C�I�s����#����i����C�	F�<t�� k>���$�T��C�I��N|y7N�8+���(�n��P5C�I�%��Õ߳CơJ4�L�Jy�C�I�K>l�x!o9�h�0p�H���B�	+kP��iwe���*�NY{f�B�ɶw?���_�p�H�� \�PB䉹X��E��`�3OT��GQ�B�I�RZ���F��0l[*	"�ޮ�C�$�"\�Z�4<�#�;{2�C�I{h<T���$�Wb�=��C䉅tѪ%9��ά8��E�T�j�'x���T��.�@#�T9B-z	�'�~��A�ØJ��}9��:7����'ɦ����sp��t��F��$b�'�^m���EB�p�YU�JG7�h��'�&m�ĉ�.�@6f�{�Ќp�'0l�YF��b�r�j�L�;!�X�
�'-vق�*�+��E���A
�'^�� ��<�H���DW3v�n���'�jqR����km�\�cDF�o�t�0�'�)+�!���^U� F�j��X��'V�@��� &~��m� o Բ�'�*\��I��Nm�p����ҵ��'@� j�Ф6��G��Bf����'����
�رt�W�hs
�p�'��R��Z<]�p@��a�~ɪ�'p����Á)O�IP��֤-8������ �UH�fSn�c�°7G��3e"OJR�썸|�}ce��JA��)@"O@��f@�@�H=)+��<�ȩ�"O8�Vf���ш��
!���"O@Ԁ���!���A�F7B���"O�M�d��hH����	?͒�[�"O�ɒ�� M��p�A27Ȝ1��"O��*�	�CR���#� (��@ˆ"O�(��b��A�"� æEt((��F��?i��v,�_X���#��r�������qf٦S!�O?�vL�0Cч���$�a�!�Ċ|r�a(QM�`��p�!�!�$^
k���h���/O���`�z�!򤐡!�L�`a�صa�Y���&s!��ːsc�Tc��-�1��,U9j
!�Ą	B�brF�8��T�tB�>c����v鬕��ꇛQ%���!�&�yҫ�*�h|�C@Xu!L�Z��y����H�pl�Ң͊qd:l�Bϒ��y�,��!q4T*��d�2qS�����y��)p�a*�N�X��4����7�y��O</�)�(�4Cά�A�����y���-�2��<� � D�� q�C�I��6H� "��aj���O�p��B�I�=u��u��9G�H�k'ˍ���B�	v��L��
�Vxze��nL�r*�C�	���=�v�:X����H�F�B�I`�u�R�ީ�(� B�}(B�	�/����U�i!D��;a �C�ɮI���*�]�!f���'��B�	"!7Hp`b&�(
H�*V_�l�C�I�S�	�UV�PZ�3ç�s�"B䉥E\�pʖ�����7��NB�I�kbh|��(	 �ؼ� ��E �C�I�2� �ҭP�Ҝ	���&��C�InG�%�ӤF= d���c� �fB�- �`�BFȜ�T����@��a�B�	�5���%�B$ㆱ��^$D��C�6@�.��*<$���3�G�?VC�	F`�q,ёuڔ1��mK>`��B�	3����o�)`5MP&B�I>0*�pF�G/�t g�/N%�B�	(��UJ�ƟS��0wD�3|�B�3�1su(�=a�d�@� tj�B�I/�~p��?F�|����n hB��9k� G��˂1�b��#Z4B�Ɋ~�ab��$oY�P�'�V�0B�	�����-ä} aP���C䉎?��V���F��9���[3[B�I+<茑�G�ޒ�p���X�C�
w������5B7$ϗ-�C�&B8 ��ʜ!\M�����.#�C�1)n�R`��7'Ӕp[�=K[�C�	�xQ���7bDx&vL�`��R=�C�I]�8�h ��u.���p`ѱM�nC�	�{Q����=|%�ԉ��ͅe�C�I'\J��g� 9y�DXSφ��B�ɧ#L"��ǌI�"�pP���c��B�I�l3$%XqlW�`��ʊ�oR2B�4��|����e��/rȺtb<D��XF��q��B���| !H9D��S6��qz�(��M�\:F���)D�p��\PQ
!��=.4t!M;D����O��K*Th#��V�0`��8D�� ��[AJW5l��x"v�MHЀ�"On@��W�U�Rd�0n�o��]�"O�i���-_�(I!���U�g"O~�F�6��-��!^�r�"O�5RcLU�V��j�ן�B\� "O��(��� zr��t!�(^I8C"O� ��h�\\\Kd�ӈkPPH[V"O�l��"�p�4����3m1�s�"O��@v��"-�n�*rb�x-��i�"O�Ł��Q�Þy�G I8;�@�!"OJi���[t �o�5��"O�5��kL"@���� ��1�p�b"O*#圊Ao���BѰ�Ay�"O���ϝ!N��s`�rH�"O����T|�I��G�`!��z'"O`��&C�D04��Ů��p4"Ox� �F�O��K!H�+���"O��{$�O�n�$ r�B�$bD B "O< %H�7+�=i�8[���q�/,D�`�2� ���a�G�J���y�'D�Tq�ī;��y3h�VH�:�L'D���A�?�ĵs��O:7�����%D�H4�%D��= g5Q��1�6D�@�EQ�?�Υ�sOt��Iu�5D����I�q�ijfK��s�����l3D�<䞮-�>Ub��/WӨ���+D�$���s�VU�߁s����S)D�@@�>@���0�ǭx�hȳ�D$D�p�ոV~��A�E%3R,��/D��hd���\�j}2����8{L���/D�(����Q�!H�M,@p���/D�82L���Хr%C�3C(�8C�/D�dbe��An��Hc��
K����c9D�(���0nb8�S�H�P�}[C$D��)��������#qs��)B�>D�0XU��!4�P80�)Z�bd\aG�=D�Ă���
d:\�AFX�y1nU�W�'D��ȇ����Kq�Kzd$� ��(D�P ��/	�h�情+I)�!��J*D��H�;rQnQs�G�#����,D��JCOQ =�QH���`�$B1�-D�dC'�C���ʰ)��D�0�`-D�<��&�"Z<���.�\��5!)D��1�F>���`�@F�,C*��&�&D�ۦ��!S^>D�$D��� s�6D�h"�?n�X;ŃQ�*��I�Q�5D��*A�%��-K��L�aŠ2D�p��lH�z���.�%eOb���-D�L�
+[E(�Abf,bM8�b$,!D��Y��8Qjx��O���4�� %D�lR���x�C��V#)�
���H$D�X�˖p��7��G-Ƽ�q�'D���H���&�C�%���ꦫ$D�|�,�&3�p��uh�1;��`h=D�Ӈ�]W�钂̅Y�^D�Pa.D�� -E�G��3r�&�,��AJ2D�h�C�qܐ����ֈP @��.D���%kJ>0�S�@6���r`�:D��@��υJ�f���C�%���� ,D��R'�E�
K���㛟u~�(�J'D���6��2^�1ׄ�r�@� ��0D���񆅔4���Pl�?��@8�E0D���堎pRH�0��Sj?��V�-D���J�3�|W�V$:A�l[�h+D�� ��aFz�4-@�
V�[B���"O���J2O�fX��,ՈV�<y��"O`()"aЛ �~@!�+�%�
q��"O��b�?JT{R�ʎ��@�"O�0�2�J�6��(��m��r�p"O̐F���\�� �+~���1W"O��GF��TN��DK�2���f"O M"vM�7�b-�4��m�Ƞb"OpС5'ӟ!`��
�	�$
ג�"Ob(��kH�0�Ե����?���;"O�E���>�^}Q��DQ�tE"OB��@@%:b�8�%�G���A�"O�)j6��N"]��o_�o����"O�i�f(��U]�
2N�1%����"Oj�"��	�������\|ڤ"O�	!�:<���
�On0"O� ׾^ޔ��Wn���	�"O� �c�z�Dhc��?# �Q�"Op���y/>�bk�| ����"ODe��C�v/��!L[���`�d"O�hc�i��۱����"On�񧫃9 ER��e����"O���vM{IZ�jת��}-R��#"O�i[F�-@��x�R �H$慺�"O�����&U��0���8�ā"O�!x�-_�b���0J�}��p
�"O̀��	T�nɡBKV�~oܕ�`"On샢&V��`\+!�Y<a�0��"O`�& vG�(���9DM�u{�"O~1�sd�"mx�Z&�e	)嘞�y�̽Lq�����@1�d�#b���yRȈn[|�Q�@	/���ٔ���y�� O���v��*��a�
�P�<�&ܶEoLl���
;�H�u�K�<IǍ�W�ʉuG��7}�<;F��n�<�צ��Eq��.��|>Y�&�
h�<���΃�֍kê�jƆ��e�`�<YE�s2 �g݁W�ʱ3�#�`�<A��(X&2�J	�5��H{���Z�<����kvX�΁I��ӑ�	X�<9o�,���*Wج!�s��V�<)%��CPڱJ�g��u�	�P�GV�<9�F�P�aWd*)���PcP�<aGc��1�\:0�	-��A:s&�H�<�d�b�|�9VO҉?-�X�b��E�<�@�;n6vX ��˂wy�];�iGD�<��־H�.Re�x�E{4�d�<��-C jJ�x���߶"�t�qCTa�<)χk팤jף���n�MC�ɇE��Q�A��|�d�ѷ`�q��C� 3�.y�"�P�`����K6��B�	�D���#q)l�)�.4*�RB䉟D@�������D� �`G&�3.>B�IVm�T:'���c�DZp]=!�&B�ɰ2��(�fGȶ0|\ٰ`��%�B�"��`I���n�2eH��8�zB�	,0Z@�P�H{_�A��!q�DB�I�%����%��|�urQթ�$B�I���dZAف_��!�!œ*wB�I/�F�'E̡a��B��P�PB�C�	>C>6�Aĉ (�zxs��V&B�Ik�l�#��̓K�)��!=�B�aŖ��A�� >�A�!r:VB�=Z,�X� D�/��ɦ F�Y"pB�)� (a{���[��Z`���.b$�1"O�(����<>�a!�M�^-*Q�"Oڐ���ĨgqL�0!���-���"O�-��U�s�|�0i�;'�5YV"O��K@�Y-s
HYU�ю
*�k�"O�����PrK� h 0Ě�"O�aĄ�6���5�M*l����"O8p��O1���g���.n�H��"Oju���]1/d�jR��"2Pb�� "O!�a
���P8k&,��G9X$��"O4�q�/�F�vz�֫�t�"OF�J�����,�FjϏ_n>9��"O���#@Z�	���Mk�a9�"O�%"�	�  �P   �	  �  =  �  &  ?.  �4  �:  A  _G  �N  VU  �[  �a  !h  cn  �t  �z  ā   `� u�	����Zv)C�'ll\�0Kz+⟈mڃ	g��,Q}~�D�\Kv����0MX)���޺l(nIe�ڐi��q���)�(Yj�J�����/�T\���z�8ł��jHp�RíQ i��@�4������'��k�)/lm��� [ᦥ�׿��� ����D�`�	����N
�u���
J�<����E a�^)��V%�U[&L# ���޴zc����?����?y��2w����IJ%4ȘA���݊��? �ir`���W�,�am���SޟΓh:JR" �)�D���k�����Z�͕'gr�E1m���蜵����	R",�:X�X��v�X���r�!"D��I L�1{�hBg���h���>ɛ'�O�hRB�N#��Z����]�0�D|ك��.&����ǟ\��ӟ���ܟ\��� �Od�Ο>{���N\U
�I���;���O����O>�>�
hӬLn�0�M[��Ld%2���u��@�(ES��̣���J��ȟ谈��@�@�.<���S����P	X�A$K��*
6l8u�z�p	n�M��'a���K�3{�!P���m<��׀�8m�x�ww��l���ĭ=�n �S� �x�Y��?f�H�i�40x��`�D��`���5u�-f�͂e(�0;�\cqX�tj�2��ix7�Y�QZS,Ra�jy�n�"0̆���`��߬eV�������\qJTA�Ƒ,#K��fB��Kb��Qm��M�P��$X@��э�n�H�q@ɒ� 2'N�ҰtBR����a�d��ia(	'f�ԩ��J�0$r���'�r���kYIc��5̝�y`,dI`��/N=lY�4ki�f�o��M#���e���	����S��=�?�ϕ�yf�T�ڕuO���K�yb��9RB��v���;���B�F��y"C&,\2M3")Y,o�̡r�ó�y�a��}Ѱɹa��a����x�|��ȓEBF@#�+�3B�d!0OY%hcb��s���ss�(j�$�w#Z��E{�)CҨ���镬��E�3E[Ry�+"O�K�Ѱm��P(���Ox8���"O���¥O�?v�u����J�Z�V"O�MA�c��Vv���@��B�a"O�u'�ʋ-���he��}fT��"O��A�D��)�\ c�l�;K�5�'���b���S)�p��m�,��gU�l��݇�h��p3�a	�ŎY�擸g��e��s|�c�eW�U��P`�\5jP���ȓY �hW
�8��`�Ï+�"Q��F����p� {}\�X���	7^��ȓY\P̱��sP�Ur�%�e��'�2���Q4fEa����u|@J�c�/JO���ȓs�-�rh�=y�P�� 
�-��ȓp����+��Aޘ���:X�4�ȓU��1�-o�hi��0)�Ʌȓ�\)��٪q�A6��������ɻ�>U	�4�?y�c�D���N�r^t����}o��A���?�E�Z��?����doöi�p��mz��I�B��R7�Ȇ
������=<�R��$^�8(��aF�Έ>��	Q�sb��	<B��VNݡ
�����s*�Hvӌn����I׃]�0��u%�*&�8q[4I_pyR�'��OQ>��0.M,+�a��N9����A�7�O�t�Ɉ�Z%BD��("�t:���o�f�$�<��]�?����'�����)�cCB/fE�d@�^'b�	d�\����ӷ~b�3�,Ώ\M>����>�\�Isj8�)§m�ɨ��>�����VEh��'|�!���?qN~b��'� �Q��1L*T8�'G4���?i������� :ysi[�\�Gb�,ڧEyV,fO,k�ب�ǘ?V�(�z�4�?�-Ol�
3���#>i�bϓSG,�IE.��p��#��#�%Duy�[�V�Az���y2�>�~y����:�d�w�ӥt���@]��� c�0|�c>c�h�ႆl&�b��@*58�#u(�O��Uhp4�IF������$X�.Z�h+�7��{���3�m���y�+�mu�qGo�!hmT��#C�4��$�B����'G�I-$�	�c�d@�a�GI�e�P����~�d���=��0�4*L�!3%iɛ4�J�x�$7�,�Ud&u1,�`���v�<�I	p�(C��'w1$�����`{��qe$�{�tUSg�O\C��!
�pHV2s�0Ё��V��B�ɃG�1�f�A#du�}�r�x*��O\�og�	J�,���G��m�.Y$d0�M�ph>O��y�/]���J�� �������s��Ck�5��@r��'4!�'��c��8�O�,��]�-TL���cV�c��1���'��m���?����?y����LB4E@���p�SKǛ���O.⟢|:��q���0��{�Y�C�H@�����c�8m��Ɲ\�.h�d�F�RA�h��Vy"�!QB7�3�i�����r>ŚqAE7%nl����(A�<A�*�O���T�V"�Q;W��J�4\�"|r�Ϟ�n�9���$��� ���Q~b�A>c=a���\�?U ���.M�܋ӌQB`��N'?�7�Yß���|�a̧T�9a��ö/S`A�Ak�v9'�8��A���
&k�74 M5�ߗDC��8�&+�v��>)h���K�����ʥA�Ɲ�G��O�B#`:�i>�<)fLB5DI���D�#�dQ �R�<��F��Iғ���G�ݺ�J	g�<��+ō>A�����*�ژc�k�<��J
_�^t��E
6���Xw��g�<1egQ�	&�I��EP�1�k5�Xc�<��C�T�ԭ(��+���±G`yBM�p>y��Q߀� @�ڀ!ڔI2�H�d�<'\�tD<��T�#?mN���V�<������̀��� 4-k�C�Q�<��J�m)��rEFN�k1�ө�J�<VG.�����!a���ҩ�Ix�(!%F���M��]�zD�C�?	ޢ�i�#D���\�H�H�!�	Im���A`��yB���]�� �.?���tBV�yB�4��� �
׋9ؔ�����y2��
K04xPɆ�h�ej��y����J�P��D	�:�I�.ҝ�hOX\����L�&��!�#]��Q$��DCtC��(g3�#�e�q�����j�(�B�I�{�L�� @I_"�΁f��C䉆KX�$B���?�:���X�G�C�ɍ?H�L ��$.:�᎖�w�ZB�I�c��!��'ĺ#���6��QF���G��"~�'#+%�L�ɤFH2�.���g3�y��0p4�4I��!,�X�AE���yb�T�\�r5�a������u�^��y�'��s��	�e̝�(�V����I��y��Y�2��Z�[!Td,�P���y����<�&��"�����`�O���UQ��|��IHm\�cFSC�>�!���<�y��F�Nr�8���8=>l��H$�yBhU�.0���T>�>���B�3�y�j�>v<�p2`��Mhb�b$DJ1�yBg�).��h��F��P�	%�A���>��m�o?y��K2nc�YQ��\*�co�u�<qsk��\�D3���tFNMBc��j�<)fM6Gd�Qyt-8�h\��%�b�<��Īwr��Ի��l�E�S�<�Q�V=/��D�@�߸L@v ���Q�<Y���E:�4��̶J�r,I�!P�'�h�X�����#͆@�&޵<h���!F�]�!�E�Z+\L�%2E�;�Jڋ"�!�$�6
��(3p⋓�V���jӲ9!�䕔̬�HFo^�{���U�B�;!�$��MB �Q�*Ed���[Y�%!��_�����k�2<\!I�e��}g熏�O?9ʵ�Ϙ3^�Q㟌^�vI!�X�<!�mN�p�P��>"O� �KY�<	�-ɥw�ސJ���8j���ehY�<��&���u��e��u��PƩ�T�<$J��6�ⵉ�������T�<9��� \�\��A��3�훴+�Ry��л�p>Q�l�;Z$�d�u��H�V'�K�<� . �Ť��-�8 �D��z�N` �"OB��e3M�8�����l��T"O�Er�އw!�����<i���"O�E�FF��r;<����
�h4�6�'���3�'l0�{�)ڶE���Kݬ^�� �'Kp�����;�zP���@��x�'C4�v���@�����#d�'|��FK24
J1ꔈ�+�P���'�d��v����XT�d(U�lP�'adYr&�V�}p�ZdE҂ޠ����$��&iQ?�JG �Qk�)bI�>B.�
�/D�,����?]������l_�-�r�(D��H���c,e�FKD(/FT�C(D������#�(�(��R&-[ �$D�@)�'Y+'�6p����AE���/6D�����;\�-�'*ߞu�����O�@4�)�'<��}	 6R�\����.�(D�'�:���e�)R��h4���-�8A������۬|�8|²-R�JY�������V�q���DL9{�bB���Mն	6p�Y-<���ȓ=;f1{�@J�sR��)�D�[���'�0�:�w� �Nݕ
�T���O�otz�ȓ��"�΂fK�Iw��%#mRĆ�$K�a�n�̰�mL�/���ȓ6�!x����i[rFռvN���ȓ5j���ȟ��<�q
S�C� ���q�h���l�5r�ҋs2T|+�(Y�v>xB�I�B�Hh0�@(a�0h�nû|!nB�ɫ?-�Л� �I�� C�ԛ� B�	�2s����e$P�Ʊ��+Q!
��B�I{Q,�����`3kN�PC�+D�<*u'��a/vqx�I��\Z�l���5ړ)p� F�t �c�< �/TL�؍�2l �yrΜ�

`P��[.T��؁�=�y�GX!��T�#A�EY�xZ���yb���&�N�s!_=�� �*ٖ�y�K�x���@�Aް;�,�q��y�[�j�$�2���r ��&�?�wT�����)�f]+&�l,j@�+Bp�M(D��QV��(1����$�\����;D��x���*h�p܉2�x�>�¡c7D�@�F�+���D23*4�*D���,�H6\Xq�bA
�E�4L*D���N��$�Pk��̀�,0fa�<Q�B�@8�ɴ營c���B̏\B�����#D��Rq

*{����!V~2 h��$D��3D�)>qb���
�`��q��%D���RS��J�xRc�*!� l�¤%D�@�7��+Mz�{���S����#�#�Ozhb��OR���n� zX�yB�Cr����"OXE��h_� ~�P
!iĊQ6ԝ��"O�Q��JñJ!����h�s0~ ��"O�Qu�\'I��x���o���"O|��J�6"�g	�SP����"O�ؐ�BNll(5�����<�����ɰUɚ�~"7��~��䉓7S��u�D�<9��˓/0"Dia%݆g��ؖM�|�<Y��N��vH��O�P��k&Iu�<94K1y�21�D�z4�w'�{�<�"�ѥ^�Р8�e٘�~�e�w�<9a�	L��� ��mlP�d���d;G>�S�O&m�&�3A���ʇ��/"(��6"O�L)F�\�b�lܪG�	0��=�e"O� �8��M��G����S�BM�"O����Z�1+�&�2���"O�x�!H#�>Ő��G���  �"Or�9�gY3�1�żx;�9�\���+/�OF�����S(Ф;�m�_�X`I�"O0�3%)��#8t]z5,���\���"O,����<�6|�rj�&�$`I�"O��k��Ȇ6�b�p��F;�^���"OnY�R��-j�Lt��H��xTT�C0�'��	��'n<�)�h�'"fVUlH,��iV"O���&ҷ-��@W�I��Pb"OhDhbcQ-'{�,PB	 �� hF"O�������@a��C �ٝ%�(]�"O,]�Pȍ�^��Y=2�J8˴"O���0'�*V��ؠK�kQv���/£~���U'2v�y���{�V��%��D�<�iT��"�3��֭pv&��2�x�<��g�a�������%����^�<�̕%d��9P�
?m|4��
a�<)�Oߵ'�Pk�DΪ3=��6W�<	e�	h8Ja��*$�>�'�ɟl{qL+�S�O$ty���:��2�&W�2s�EK�"O�)��hYPRQ� �ß��|�"Or-��T)��,H���}y~8�E"O��C�	A��$	?e����"O����M� �z��7t��Z�"O���4b�\.���"�\`��+�Y�D�-8�O^Ѱ4i�epF�(��(�`<K�"O�a��2s����]- �H!*s"O�l��%ۅD�Щ�r%A�9�P}�s"O0q�tJ[�PQ�@Qqb�Y�t�I"O� ���h���!� E�@ǐ4���'8n�y�'�\��	�&�����a�p���'���Q�nk4����ح���'>��VI���Q5A�+�Dq��' >8`����ni��P�(�95��[�'��BD}��՘Uo���C�4D�[��BT���ehF�P��k��4�-:hF�4\�Z�d �T 7|m��C%P��y�����ˇJY�l0����)���y�V/h9R ��X9�%���y�N�QPl�KD	��P�� ������y�N6}�|P��5x�dJ$���y�H��(��Zba�Ex�<{R�-�?�wmDV����(:�KH�@VE��}�Z�k0�+D�£���Xu~T�F��p�
�Q�+D��إꞢ����v�ƒ���R�>D��p`g�"�\�󶋁'�d!2S9D�d��+�Y��sR�*�@Q���3D��*0�>.��)BEԀH.Z�`�m�<�Q��k8��a�S���3�b{:<x�B3D�(�tNQ��9B��&*�p�g3D����%T� ���$\�T!@MxAl/D��X"�K�oN�S��D}$#&�-D���AIA r@��SE��q��� I/�OB��O� :5n֊n�
���-[T
X�"O��ȣF\�`bHHR���3L�l"Ob���g�^����@�MOX �"O* 1`�Ǚm�����gJ�c2I��"O��X6j�;yȮ8aG�w�x�f"O���b��rb�� Ɖ
W$d� �ɇX�N�~" ��=<�a���GC�U��A	w�<y&G�*?�v�S,qb&ŠR�O�<�B��7�K��سM�tz"��N�<� ��6�
�s^e�w+�pa�@�"Oz;�jżBWpYc4j�s-jt"O@���%�0�QH�;j%�L
4�'���y���SP�V��r��
gjݱ�&Y+x�N���C�~�Y�i��C�(U��f֮���ȓ�`��Q�V�⧆)k����1����c������Ȅ�l ��ȓP���[�#R"5�zi��+;E�I��g���S��-#�6pI�>:y��'Ir�!��5�莏]( ���n};P�"O0��K�2���mזc1�l@�"O����ǘ��R���
H'4J�"ON�)ꇹH�Z�����B�<8"Or���18�t����\-
Y����'�n��'l�y"r��@����X�wǀ(
�'f �AtÕP�8�ɀ��w�L2	�'2��1�KP��j1�W1u���'0�`�c�� �8� �)B�\D��'4����D̰+ɀJ�����)D��3���'x+�lɔ��˪`0O'ړb� F�$AK�R�,��l���R!J��y"���U	
�#3����H���y�)��j����ۑu�����S��y�*I����N1�����*ǆ�y������m� rd�꧎��yBC�6=���9�@P4h9�,�wmL�?)EGb���������j�2�J�%=jP�aC:D�칒iܽ����D-E��k7D�H�7$�a�t �E�m@Abņ3D�$K��D�6�ذ��N��%���0D��2c�� �; ���B��k<4������<n2��	$�ަVI��P��<�Ol�'$�(q�On�'��활T�(k �˸�<�+�Z� �I䟔�	/�m��!�����ʢ�?ͧ���D<�&�en]��t�P�1� )�0�a��r�\9b����I	r��&j��	�hp���[�{���!A�O �1擵L�h�Sn�H}��8l���0?Y�"GQ9vp�1��%31�#���`x��.O��	gb߾b�hhW��wM� �AW��3���0�	[y2V>q�I۟!�	I�`����@�+��G#�џ���ȅN��a��IX`��S�O�Ԝ�f��"C���
dˍC~ḙ'b�{	#w ���#bZ�,��?9�tFN�BL��R�'˞au(���.o��2���O���$?%?]�'W�	�'��lV�"�┸Y�r� �'P�P��ê:f�(��M������k�O�.H�bm�m�T�Pԋ�6T��]��'��	�n�E�I�<�	������$��Z6`܂ �A	h���IP�V�2���'��D��O k�D%BΟ�\P�@�0qd�8x!HO�6u�h#)�Sc��� �&XP�/��g�'�4��̏�a��hh�I�q�O X��'��	�<�&�G6`TD��A-=&����UD�<�f嚹�(�pa�:K8�AqgN��d ��4���d�<�i�1p�r�	��ͽA��hs��ğ�Vܣ���?��?�)O1�D�#2���+I\Q�2���<��RO�4|�����,:K�=*S�Egx�T���T7kX����8dԪ�pG�:	��`��X�>c�"�kQx��x���O���:+Z$��Iδf�f��O��=ъ�$��8�5+�e�M�b��GϜQR!�ĕ�,�6�5M�@��m�5Q�	��Mc���dI.��A�~*�K�#����D�\���&������O|�$�O���O�<C�m��ҵ�?�'N���a�V�O&�БAH�eժUG|r���lUQ�0��6*[�x�Z>ic��K�390�J�"'��H��9�no2x���@�|ҳ��4j������I�P��� �ny"�'	a|���3a�ܱa�4w9��8�n����.O�HC���#G�
����J24��2_�(���Y2�MS�A*��d�|*���?Y�U4_�}@e/�3x���oJ/�?qe*ܚ`����A��A�~tz��,׈����Ư�0j�ѥ��J��4O꭪�F�M5 p�C�X0����ȃ=8.�q&�@�aLj%� C�{+��X?������T��� � #A��#N���j�c8� �"Oj�(���F���sS�\&A̤���I)�ȟ> ��5HpR{��ΥIR�0%e�O���O��P�/R���O����OPԬ;�?�vK��1�a��Y>Vd���@�5i��j �'@5*� C�;�^y�͟��H�Σ)�Te���.�R'�"�4��I!g.Q�r�Ӻ�Ο�xzw�N�er9�3��z3�0�f�1?Ig�t��o�'����+ЦQ:%�B�~Ur����&�!�$E�v<l���O�H�t�䁋�/�2,9��|����'�nXR4��R�a�3ML��
��:��q��I7���B�� v��w���<��C�	a]����O�'C�a�焕R��C�	  �$�g�
>�Qpq&P,��B�	#�H��V>�z��,���XC�I�W�JQW��* `C���n��?Y0���<�����:R(�㋱f
�����7��Oִ��
�(�b�9��?s�8Qk�kD��L�j5�ɜ$(l�D哙1��(��%:j<�"�����">9&���p��F�Ӕ�D`"gQ3ڒ�P�E�u�	��?E��i���h��N=+ ����ş:_~�}*�<ie�'\UI�C�ބYh�P�G�Zy2�'b�'i�Z�E4���B�0i�B�Ð+N&� @��o�'�|�aʲ)D��R�J�������O�,)򥇛�94$�Z��y�����d?1��OZ�T>�ɏt���:s�V.8T-�b/ڌw�^���͌M~R�,}⃌��	;�ħ�<Te�o	h1��iO�7<hع�+<}b)���E��'��h�C/	�`�R�`R�C��a�Bdφ��	��'T|�'�N�'n�$���P4L�B1�0ĝ(�<��	:���'1z}ʉ��68L��З�i�,�EQ�
xB��L�}��N��I�Y�O�qn's�D����l��)`�`O�{iʓG��O,�E�D �=8�؂�.�&o���zGN�~��I?ra�ҧ�9O�i�&���S�*"��P�P�Ԝ1*�0�&č/>��8nT�'�� F��NO:Z�ap� #TE��߲�?AAè� ɰj*?��y��?�~�.87��xb%	�P�a�
��?Y�*�O�賲�B:0J˷��+T�F��*O:�%��7ig����ݜb��`�ܴ�?�����$�O��|�+��J�t���Jd���,)�tq�AJb}�|�T�E�d�	��УI��Pn�4��.-���hO���Y�P�ߛN���!��'�8 4"Ol5r�a������⇆�w��k�"O�ܳ 'S�v�\8��K�N�q��"O4ۥ�ɶˆAA��N:M�ɂV"O�I���H�!D�he�>��H��"ONI�e�ʹMG����$�5kȦ�ɖ"O$ᢴ`MPzx`��k'}�
�'Z����J�d���{�
A?"];�'��Q���Q�<R4��+	��p�'-z�!��:wL	�p-��;
�']1�`D�G6\4HA�]�����	�'����L��h	f��tAӏ�a@.j���C����88$��ƅ	.�B6N]9n,��k����!�ti�P�!΅WP�V�ɟf:���g>,N8�2��5_�d,ȅ'�H�c���/?�	S5��JmPq��A7h���9��ěP��0
���� #�H���|��
>z��� �\��'�:H�§	8	g������ l���'�f��G%� (�4kB�L��'�9�P�ts�x��C�5�
���'� ��<y����n�.)n<"�'#B�I�Ȑ
Z " 
�.�(Y�P��
�'h8�I3g@�Y�$�3q�%p~<
�'�2e���]��	j���j���	�'|��$K5g�������s,�1�'�ʵ*e@���i*G���M�ʓQN0yu��P�����s�V��ȓ!^�T��y+`)$n@�qk85��)^�� �.@�T�n`������y�ȓi۲P�DgRD�\� 
��-����S�? ����;]$�-���X% �r"O��cRmˬ<n���	H�"�"OHxw��o�\���.�;*l��5"O��V��Pr�x��L�x�D��"O`�J�B�V��HI���b��}��"OX���Ƭ.���h��A����1"OVxbP�Xʄ��Nˆw����"O����.�9Z��x&Î9ei�1��"O\�0���<NT���ₔ
Q:���"O�z��Ji�$k�kE<�4a*�"O�I���!9��!�
�!+��U�`"Oj�w+^�0�4Z6i3��yC"OR�#i�'�0�ӧ�=AH43�*O�XJpDA	"{�M"#o�:���'S�P0�"��tѨ�����#_�9*�'G�������]�*��.F<G�.X��'�n�a%ʤ <h��D�=��b�'�zu��͞�
E�A��@R	l�5�'CBh��m� '������F����B�'Z朋�뇿<����1��� A4T�
�'�P� T�:0@��gŤI�.���'�u����2F4�a*C9�D���'���`T:O��L��.P��	�'�x��/N�b�[�&0$1�	�'���T,�����,Mx�	�'N�*&��zRJ��U����`r	�'��a�9yY�=K"m�.*��H	�'$� � � w�ȁ6)�����'H*�R�B�zX��@��}a�1s�'i���WI�@I��#'��*Hh���'BT�Ơ��I� ��&�1D�f�k�'� E2'�;<	�<�� �@�����'8�xൌ['=L��U&�3<����'uH�Q�Q+D��5��4q�
�'�Dۡ#E�i	��'�®Z4�
�'����,R�%sX��/^�|f� 	
�'x��*fhI���yCh�!Xxl��'�.U�� wd�C/G�`����'��J�-O��z�GBQ ����	�'����5�ʠ{��H�6��n_ڴ��'mց��`������cP�e�n�I�'�l$��8�҉��*�2[4D�A�'�ࣦJ!X��4���T�����'���:�)^"D�@j&QDx��!�')H�-Z�I%lAŚB9BQ�'�,t/�=7I���Gȃ90X��'��8��/A���"�/]� \b�'m�3�Φk��}�1�\�����'�B`ڰ�Ȃ=Ht���C-cT@��'N!�K.;n,t ��Y��8A�'�ļ2p�ݲ ��A	��Tzv0`�'E����h�/B<�!K�J�Q�'�j}��&E+U�6��T'��ȶl
�'�t�7�+� �j�I1����'?�dY��E9 ���FV>)��T��'hJض�C�z�E ��
�"tx`�'ֆ�+����e�D��L`�'��d���~�uQAV��n�Y	�'�:�Ib��Ԩ;���"u"Od|�GͪU���H�2=0`��"O\�JfEZ}�{֠
��;�"OD9&ݴQ��	K�hF81�{ "O�)[r�]=0�V��7b����Qe"Ov|`C� ;:d��W�ʙr"O� V��`C׉ؕJ�* _�~��"O�a�/K7 y�l�U�S�r=���C"Opx�a ��o��<��đ�-���s"O�p�w��(j��䘕�T�p|fx3�"O.0�*ܣVDHM{с�$X�"O�Q��2qdL�I��4���"O�2a��i�Hċ��W�-�����"OB�aQj��>��9u�ݖ
���B"Ox	�ej���l�j�k�1D��ݲp"ONٲ�x$Z\I�H�8��{T"O�4��ŶC��xc�I	Iz���G"O�����	�SzM�W"O�`ύ�	~D��G�?{L�
�"O��WÓ�,`,{�F�RK��c�"O��sCL�)=�ج���D�52�"O���c�"2"�|J��j�9:g"O�s���)��TD2
c���"O��qn˕}�	����wK���"O�bAiG�V����"�NJ�1V"OxTh�č�0�:�A�;r���HW"O��!�Ƅ��z���xt�H�"O(p!#2���Y��/	g��J�"Or�A@I3Gl^��R��WWFPv"OY�r��<����e��U��;b"O�	f[�>�ҍʇ"M'(C�7"O\]��)�0u��Iׁ�>-�1#�"O��ʵHUGQ���+�{Tع�"O���E�ؚ7 �a�k�ms!"OA��@!S ��3�]1qL�ɚ "O&Ydk��-M���_�^�r��U�y"�\�}��@�sdܽ:z��gٸ�yR��9�x֍ܶ,c�D�3.�)�yr�
a�Ra�R� '����*��y���>=��ۑ�X�N�t�G'�yR�l�D�W ðM԰H	��'�y2k�!*h0gL�><�j����y2G�"f+��
�&2J�i�m�!��
H�X��T@ٚ_z�:��Z�{�!�DX@%zT��%[ �"āL�!�Rtp~p*'�3CNjP0Î׉}!�dJ�)%v�C�AF @�G��_�!�׮hK(A��2+<��&Z~W!�S�5� ���H9i9N� ��,�!��+s��K��Ԃ	���e�D!�d�O耐:��%{m��/EI!�C$x���o�e �G�
H!�R!�
<�0 gIC�%S.5a!��ΰ$��mБ�ވ55ibv*�MQ!��'V�B�!SmF![* ���$D�!��ǋ�B���  {�(T&pv!�->�j4�'hE�9z@qr���qd!��Rj��$����	x�Sb@U�tN!��!Y���"al�U�"Ĉ0��/[!�DI00�	����!��8��ܷCr!��J'-BY�@���B�*T��T!�$c�����C�n�"�Y�b��!�d�Q�
�q��.-��@��vz!�d\�)�6`��_�N�d�b�]$f!��,
y����L�nX�s�B�DE!�D���)ˠl=W�J؃4��'-!�D��v�d��v��
~_,�2�jC x!�C~Ǡ$2�	�b@8���HU�mn!򄉎\
�P)%��h=�!��{-�ٚ&��>1q�ܒ�(�3 !�� 9��:�ܤ���L�lTJx	"O�@��O1L1f/O�xIp��"O�u�7������4΃<?S
�w"O�1ɶ̒�Y���B�ʞc��D"O�x����c�
�:e�,�a"OݒEgŭmu�T{ċ�;e`q�"O�r��W�)�
\X���1~����"O���w�M3l��[Pj> @��x�"OtA`v��!��=�H�2ɢam"D�����]�AR�%�kЏ:t�$D�@S����mHhPX�'Ͷ3SDq�3�"D��� �F�|�&hc�K�1p��;D���ga�
F܅��,I;[InYXҪ-D��i  ŝb�b����DH�&D���E�=6׬x��(�-;:���j#D��Cg��(��E�6u��WN D�pQ�ǁ9ly�h ��#]Q�tWE;D�0ҭ�+���K��(]p�T���:D��ⶣ��w�T���R�C����b:D���j̕a�ѻW�nپxb��$D�`Bg!�{�5;�D�>���V�#D�X�T-�[���#dD2�v|�TL%D�D��Imo:�C5C��bq2Ic"�!D��b5||�(ac���6���>D������3jJ��c�Ypd�:F�8D�x�b�^�)����B�e�mIb#D�|��E�0S�X՛1JՁsˈ�r�M#D�0�L�5Cf�9ie��"v"�R�"D������MIX��2:
�@�č%D�D����<������-�~Њ�`"D�8b̒@E����+�wH`�T�?D�ԯ��J|��#R������g���y�L�m�b�*�B�	��l�cះ�yR�_,�H�+,�r�K%���y¥%=Q�A���R4'��d��ۯ�y� 0K��d�וo���h2j��y�Z��Q�-�Y��PR�T��y���9���w�$7������yB�ѴR���Ir�K��xQI�J� �y���|�(}�R��\���C���*�y��?L�L�1P1RW~��۰�yr�׷*"R�t�UE/�(�(֫�y���91ET�p��@<<��� ��
�yB����h0B�J�&L����>�yB�ò8��!�i�T}����4�y�#�����΅�>����-N_�<1�&�/0ub0����V<��W�<�����U��#�m��(�ϋV�<�`�=����+���
\h��^�<��L�:9B�rOݤB=���R��p�<a$�G�J%�B���i�8��c��g�<��D�@�!d�˂v�v�`7�W}�<����2t(*���)
�g���Q&�x�<ɣ
�"� �rt��'<���Or�<iqLZ�uine@��Q�u��B�<�w��ZVQрBO�V�V�KC�I�<iL Lj��Qd�D&8����b�C�O6Ip��I#0 �aSA��2se��$�8@���'o�:���ٌqn�ɱ�K7D��#ň'd3H�
�A&.��*�k:D��ᘀ��)k�/˙0"�]
g�2D�8�SĄ3:�^8�CWj���o$D�lJe`В\���	��)z|��!D�\�',�� ��xJt��u�ۂ�!D�h�dB]]��{ӌoN�����;D�� ds�ဨ+��bhÂk��M��"O����Lږ"����%�3�-��'8|�a��P���x�}mn�	�'0z\2��O1h�0�9R���#s�X@�'GT�Z剕�A�H��'�M����'�eZ�-�$^���e�[�DdY�
�'��@��N�R�tMw6�H �'Ͱ���,�t���T�Hn�`��'Y�D�6�U�=nt��J��g!V���'���P��߭$/p��O��nQ��Z
�'7F���f�O�� aC=t���#
�'�Jeɤ���p_t��!A^�n�tz�'Z�0���'8��� 1�M�"�#�'��A �Ωm�V��P�
�*�'��m�eK�'q����$	H����'�p-b�oP� &έc�#n��'�P��]��,���5\��a�'}t(��.�
S5�V��n�\�3&D���2�|ڄ�:RXՑ2/D�h�. D���Z��M�_�V�b��,D��Hg �=3�.�r���X�>M���*D��	(äg9h��@�� ,ɪS�*D� kׂU_�#�41:U�2J7D��S慍">lm9�(��� �:D����A��jL��Aʙz�j4��+D�����#~3�Z@��h@��{�<��`��l�l���R���^t�<yfO>2��7�Q���A��D�<!�^_��(��TG�6�y��Z�<���q��V�\˒٩�X�<��lF�<4� ��fP��9o�K�<����p�9C���^ʈ0�ƅP_�<1�K/0h\��A��bᰔ�W��e�<Y#̽�9W�ٗAx�XD�G�<)�Efx���͛&ˈ�(�A�<9P�Q8�� �W��ԅ�X�<�Q�U�2R��5���X��\T�<� �L7V�zU8-E�iy�@��AS�<y�0Ӏ*�#ӬE�<��ff�<U��2m�؅�&�J�h���a��b�<q�ɒt��rb�%_�]ڲgQ�<a�C��iXг�#"@N�霤IQ!�� >�x�ug҂L�8D�v-�5%!�E�'��m!w�Uzf�.!��fG�a�"*��=�B 
`P=!�^��>Ʌ@��"�zM8GoHDt!������,H2�|���M&o!�қs�l8X���1\ö�j��Dp!��̅8(���Ak�4�) N:AS!򤄊6�ơ�c��<��8"�M5tO!�Dmh�*#�=o v��L�o�!�ص)�����٨a�$:R�R��!�䄆��$
�N�9�^ ;g	q�!���@���PQ��R�X��E���!�$lO�=Ѓ(�g��k�%	)!�dK|F���΄�x7`���ŝ�!�d
�t�Ra�~ƌ�z�KbR!�D׷g�V)A4�Ӭp��DJ �&Q!�'8�����
g��Qǉv!���,c2��%B]:%��Ʌ��!O!򤐁2
8�j��ت4�$dVÔ�6�!�d�V��i�1&�D����� �!�Z�jb�QcQ0^	�P��N9iF!�Ě�=���`U'Z"ȑ�f�+hB!�� �%�a���2��Td��8U�)�B"Ol�p�
@"(`�`�d�]8F-,aj"O�9�f�ܗK���ҏ��R,> ��"O��D+^�����-Ό�>9Y&"O��T.�4���o��HH�	2�"O�QTL��6���q(��hA�Ii�"O����K�R�	�A��.���r"O`|�7�D�rHZ�H�Q��R�"Ov�IտS�29��.ڄ%���Z�"O�8*7�
�:8�Xt�H"1N���"O‡���[|ƵZ��C)Z�����"O`(qAаJ��LYRj�@�ڝ�D"O��b�%�97���$�ȃmN� �"O�!��Ù�m��Aʗ�Q�S��І"OQJE��jc(y��ޞ`�t�A"O��r�F�R$�e��܄�a"O�ly4�A澶��~�"Od�g��
w� Q#�Y$av���!"O���Qb��aZ%䚳dg�U��"O>���'�#kFrc!ި��K4"O����hZ5O�r9
�
1"�̑c"O،8��t���X��o��8�"O�	vK�9W�$��ʔ;��r�"ON,#&�D<->�xs���M0Q"O�p{�%�D�ѱv�� b�Q��"O�b�&��'֎h(a�@�|��أ�"O4D)W�ګ?�h����"�Hp"OL+fLʘ� P;�W�Zt,�S""O��{jτ*�^H	�Y)6i���e"O$dbb+̻D��s�(��p��"O��`$j����1Id`�5�h�.���$w��]0TgG&@��Q���E/[����"O�YIąo����ai�<��4�'���<A&�	K�<�!r�"bʠ8 ��	t�<a�O�jb=����ˎ���F	wy����M[rD]vʸ��#/�$h�9��gKz�������'�V��ȓL ��y���&��L���ͭc�)� ���G�m�ɴh���8���b�3�\�r;�D�=Sz����
�
���KC8����./0n�92�_�+%+�߿r�>�IÃ�[������:|O!ڲ�1I�%�$���C��E��ɶ% �H� �$L��'
7�ɖ�D��,r��B��SU,$�yZ�P���
�hM/=�]�J0�~�G8�z�c��J�z�`aB%W�m�>1��US���Q�C	�-�ʧ�:D��0 Y�X� Ѣ�J=x��TY�A����� J}�ՁC\�E���O�OL<�'`�@Ƙ�#�8T}^d�'���2�ď 	�L]r���0�TZ���Dz|��������Y�EXa{��P�g�9�nO*,&°1���O�tNرk���f*�PîH��`�]�&7R&�*��Ŀ8:�HT�8D���dI:��M���k����#���{�dZ�`}�Y���X�
�j�,}�O0jB� �p�z�6��%�	�'�:,S�]-$m�l9�U�ig��ڐ��U���@�Nʶ3QZԙr.���g�zb��s#�,s: �X�A��Y�4���� t�����RC�d���#M>�$!��"@HZ�(1�Y6m�<<���'N���v�D)I�}�#�M,^���A���ʙS%x%���<v1x؁cq>�zvg�MU8�q+T�p��7l+D���:h8�ݘgJۣwf}` �<�rk�	-�X���8������8e~HҔA�k<(���X�,�!��]�bppg��%\:�W��T����`�F��LIJaaAj�g�I7K
�i�Ƭ�2j�-�`��.`C�E{89���O�yE
x�k�2h����I;���S�'��ʇ�^ ���G-��N�L�`�����C%�����>�X@��m׫
^�ɩ��	&�!�dK5PmB���呹3Q"�r  �X�qOR8@8�)��D<l�����z�ʙW)'Z�!�� ���pgѭ���1p�Y�%�Ҵ2�"Ox}C1a]>]�r]�6d	*u�Dxxb"O�(�0Ή�5�n̛�薂w�x���"O�HҖ�C�c����c٤M�U�`"Oj=�g �����S<����"O�mCT.�� ��p
b+^�"�Хe"O�1�1�S(Z4hD`�Ajx�"O��jN_�\^��b7��\�����"O�]��j�$��̙���_?zY�q"O�$rQ�D�v䃒�q1�|k�"O��1�B<r��8�����P�s"O�mK���d���C,F>+�0�I�"O�UʷBͺ4U� �n�&8�v��"O��n��M�F��-F�	&���"OV�@0a�z�ܩ��̌�(�%"O�}�D)�1-ی�:��7
y0�"O\�òb�-���v��+a�TT"O:�*bF&�\���WYt8�"O����S�.�n�רR!?V��"O�]��h �8���icjK'St���"O�,h1dֈ��Ѻ�cK2T��A"O
(a`뚴A�t�3��?�|�"O���o��N��5��(^5D#l�8"Oy�`��,?L���鄊d�`h�"OXM��)"��%��H� D�t�a"O�(8��
��!��aV {��Xa"OR�D�(;vdaZq�=<��M�"O���v/"x.���E�5\)~�"O��#d�&v��p��#V�p�"O<0q"�J61S����T�y�1C�"O�MBIMj\0�ZE�Љu:H�ja"O��Sf�G���#V�Ȃ+��H�"Or��K�(b,<����yBLyr�"On�۱�ƽxM�����/���r�"O��YA�7�~L�0��J�8A��"O����L��*m��`��71�V ��"O,L"���u�Ѩ��]���PE"O�8X��"5�`�f�C�}���*""O�\h��ܓ~X�8�ة!�,�C"O����W>U��q&g�)��)��"O�����P(���G0+���"O�%��� Ne$��u�*Oj�[PJͼA�f�"b�O48��r
�'��oE*(_
��IC�c�����'���AG!��6��0R$��V@��'�`Sr�J.s%"9#Ȅ&=� ��'ⲝ�bD��8:����(-[:z٩�'�n�Z���$xv�	ѫ�0Me�-��'��H85H�394e�0CΫ�� ��'���[�$�|��|�#���t9	�'lXȂ���4T\�
�#U�5p�'"�L��9#��er��Mxؕ��'�����
�?=�U�BI4kF]�'Z-��	�8EK���jR..Ġ1R�'�r<˧j�?��&�[."����'e.�`t�\)r���D�ۣU��s�'�����Q%��QT�]�N��0
�'	&�����|#�:I���
�'j�4( �@�v!���Зv����'�J8��!�EW�0��P��V�q�'�S�k�&��1Y�h�O8�	�{2M��!�n9�Đ|S40`������&��0A'�F���'��N���jt8��iI�[�B�`��-Pz(���v8hrƓ=�`D�Vf��i�X���S�? �U���Vt��Ǘ�~Ȁ���"O�MR��"p�k���(8bV=#�"O�L�vC���ax�G�3�rE��"O@q��N�L�tH�Ƃ�M�IkA"OP�æ�E1�P[tE�w�H(�"O��`�"P�Y�Z��8�`"O~e2�NzMt�0BJ�9$��f*O�u���m���� ̵8��Mx�'�q��T�P�I���a���$�2D� p�J�H���@f !�R`�W�,D��rצ	uk���t*�SQ XR?D�$���U� @Jl0��N�"�DECׁ0D�dI�g�7~�QJRv���a.D�l�b%�/u���[�V�m�0�?D��b�B::�PL��d�gp��0D�!D��`fm��f�sc�Փ4���C� D��E��Ufp0��/,v�ؒ'�+D�L@C�Wn6�{�ѵ;I�L��+D�,0Cf�G}�2t��:n�ڀ�4D� +0N9c��$�bS�cʲ|*��1D��x�$LK�֥O)8��0U�1D��83�Ń	i�\�>�d�j"�5D�Ĩ�ӠLj��{�,O3D��I(D�(y"&�8b"B5ht"��u�Zd+Dg9D��9C�΃Z�*� IC�y:�c2D�\�)O��ɋ�'2�� o3D�L��.�&Sʸ�dbR)k�,9�!$D��AmN�)�<[b%,� ᣷�&D��A���.hH�N��@�8 ���0D��j�E)tVu�p�H�H�.,#C(/D�ܱ�D�2&�:��R+�`�&�,D�����Y�^���e��R�@I�*D��u�F%`ׄ�� e�zV�q">D�̊�ǈ��4��C["k6��0�<D�0�ޕMP~HY�EV0D�5��;D� z7oO)3��QG�1-4F�Q%=D�,Q'��<N�p=�^L�ҍ*�y��P'~����0D�&�[qMU"�y�2@f"pj#"Dv��`�ĩ�y!Ğ6�\�3E�G=4��q����yү��2����E�d�M�qe���y�1:P�5Xˀ�`Ao���y�bڒbNҕS�݄"xy8��A��y�-<`/�<��Y'�PQNQ��y�K"kUFXF�<#-�ɡ�����y�'���e#@��~��f&�$�y����0:�nԫ  x؂�N��yr�C�!D�H4)�b�-[�Ɠ>�y�M0.:�!�ω1k���sȂ��y2#P:#c�X��k�:�T�X�J
�yr��$k��$�$� C�����@��y�$M�&�Th�U"M,P2(�G�� �y�
4k�M�4�Q9)�M�5@��y���n��1� HY�R	�����yb�2T	y�!���Pq�t9�G��yb���@��@˲!��� ����i��Y;ĉ��@�F��f�P�����ȓM(���	��y���пT�`��fl|\�A�,{H�@�JJ�p�����\h��9 �t�AVH�.d7N|�ȓY5�)�/£Dr޸*7@'p�2��ȓ$S�Hp�Δ/dv��L A�t�<���ܒZ�
A�c�R /C��A5m�n�<9ǯI��A�E�v�mY0�Sj�<� �\z��\�*�`�fF�t���!�"O0����_%*ҕ"4�[�/.���"O��� $�-W]�H���ݠn"��A"O(�3��H~����P�N0M��"O�AC�D��VE�#P(G�|G"Ojx���D'<��B�����1�""O� ����͓7���b89�"O�T�g%ӎdq���#O�3e"OJɸ�8KP���mY�K3"O�]�6*Y�]C���&�E>L�l��S"O�A�3F�?3�UR�@@�.q=Q�"O��g>8uVd�c�O�ZNMA�"O´�ƀ�.�V4;��E�v0�"O��:��&/���񔥓/c��Iu"O����J��+:��գ��v�xa"O,�#%��q��0��H�*d��"OH=�B���?&�=�4Ex|ʆ"O�H��-#D��Q!L�����"O�1�Q+�r������R0P`"O$(`��� ��4�	D��rq"O�uC'��6U�#�a�x�$k�"O�5��L��M��X)9g��k�"O0��tΌ>Av���-� cW"O��f@�гO
�p
h�V"O��jK8bD�r��_��RU��"O�|�'� ���@ �3���x"O,��'�ԃ8�
8;Ј��)A�D"Oj�Y�D�b2�P��Hϰ�%����y�%[o��4���$4,��Ʈ���y"O�1��z�&��9�厹�y��8Dt�+��W	��d��Ɔ�y�*!����F|[>U V���yre�m�>�:�bUokv,RB��	�y�H��.d���\-��RaA6�y�X@��)� Ā�TiJ)�)�yrK��<�*�N�P��	��e��y�0�pp�D�IE�-�aZ��y�\_9~T���m-�U�WM]�yR��/B8b����Īd�2!�B����yB'�9f�ْ��cL�8S�@	�y�-���4�
%28㡌���y��T�F��}� � }�~�:�'��y��'�l(�R��$����n��yr��T d-ԣ��%Y�d��y�Ĕ�Jur����Q���Ś�	M��y2'�/>�@̋��\m @Y6�Z�y��\.7�0x�_Y���j��WL�@B��2*0�fU�vh�V��x`B�ɌU4�����,3��Q1 *��4��B��WN~�C��W3���s,�k� C��	fj����K;�l�1N�k�B䉷{��`D��Q�����K�3`l�B�I�I�dRCg�1��y�B�C$�B�	�"x��q$��af�AI�jI��B䉲<rN���$��k��m3TKX�d��B䉩!�Ե��\7PS$�H�cՐ0k�B�I	1�B��ץӟ�H=8G��

�B�ɨf���फK�t�h�đ>L�΢?Y��)
g>��uL�.�R�`�a!�W�2���#3�1^[��q%'�*M!�A!��X�@���IZ<x�2�NM!�$�E�0�PÏ ;>Pi���Šc@!�DV	E�(1� ˢ��0Ys�_	k5!���K�r�G���3��h4��&!�� �p���	-i ���n�	��e�"O~p�M��h�<���lU��~8;�"O�,H�⑄o�����3�
�*�"O�X�#�59p��N�^�8|:a"O`�J�ˬz0�@�U�\�1j�Y�"O"	�e��Le�$h�K_ 6-�D9b"O2�s%L�-
�#E�̵t"P��"O���M��`_>Yj!ޒgv��"O^%"��4;���!�Evy�"OR�{�g��1�Ѥ{�x �"OB��B���a�V�Y�8J�l[�"O�۠�ŏT9�@����D백��"O�\�!�R7_��c� K0��"O��B䝮]4��ġ�"t�`�C"OZ i�Ȑ�@�������t<���"O"=X���:5t%ꀊ��NǶ�+%"O ��E́
R�:��U�L��"O�iU"�"E2���*
$���"O���O��QԚY`ß�V��J"O*@ ē�h�
-�3���P���"O��1'�X73��ȃ�!Ls�]+"O�@H���4+(�p�DYl�A"Ol�8S�QkQ�a÷��.��l�<q��F4Y����� �.�!*Ї�e�<�Fe��{U�m���P�2��x�a� ]�<�6�4r�I'�״v�L�a�s�<�v ^�Sa ��/��W�(��&
Qr�<��+��#i�ժ��6؜$QG�h�<Q�웻q�P��ǔ�����ƣ�[�<��&E�j��S�JG;~�@�G�@V�<Q���#y��7�Jݣ�L}�<�d�d޶�3��B3Rq�y���t�<y�Á�[�4 Y�#K-I�^�pb�\s�<�Ӈ˲m��`(�*��xl�E�<�6�d}�DE/�#vذ���\�<A��	"uJҽ�S�Y�k�p�q�Y�<�1��-����K�>��x�KL�<�����a���@#�=o�����b�<QP
^�rpY�f�8���E�w�<�4��c�6��0J\�\�"0Wr�<9��K��嚅H�2��JU`�k�<��-6Z��e݂E^<���Qk�<i��L!x⦅J;_������Oe�<�`�3^�J�K�X���e�<!�O�6�F�B5��� ���ZC�y�<�4ᆤW��E��%�?bm�XZM�<��h�;yԡ�$M��!�>���F�<��tk��"�3)��D�"��k�<�`.�'�����/(7x���CA�<��	�3��As��/7���bC�<��b�{��!FM�(�=؀��}�<�B�V(/�4xd���6�Xh d�n�<�&�1p����_|y�p�ƪ�u�<q"�ExA$|�D�هf�@��BkKr�<I7)V�=M����
D��ڳ�q�<q���5�@�w�=m'|rg�Pj�<�EN�/=�Tjco��y/6̡���c�<a�EE=%r�����p��R"�y�<y��L"�l<@�(Z�i�n��1&�t�<AcL��4�P�V��2��h:��Gx�<��� 9���j&�#0 ��y0�T_�<!�n^,	�vHP@���aԮ[Z�<�
�I��TK�J$}�YQ�b�X�<A�/΅zL��lB9V�:�6��R�<� �Q�'։za048�쟣K,&i�f"O<t��b׮};�pa#+S ���a"O@�t.U�kY0���9�h)�"O4�ˆ��,R��A�C�3��1B�"O��vIK&?/�Ղ���	1~�da�"OjY�e�
�RQz���K84t~��"O4@:�d�#,�؈8Ջ�&n ԡ�"OX�Ф���3#��{�m�1g�:9��"OHc�^l�F(�RC�?p��H "O����_(�jF톇ye|�HC"O�XDG(L�����8MV��[C"O��%�.b�����F�BH�%"OԴ Nw�+`%�,+$��"O&��҈Ҭt00hBWk�S2�cd"OB�S!�t��=���φ��xk�"O���3/K�;���@���#���"Oh���j�\}��� (�)r�L�@!"OnE��IJ�
��u"�e!���D"O�d�á�4\�R����ت��(5Z!�$X,#A�\���5\&Vybj\�qC!�d^�z������Z-+ �Iq� �c!�$S���x�ã�&��p#ņ�xT!���$�����)Xn61��G��!���<�"�	5DP(y���b��1c�!�DB�3.�[2FT�T�$d(�(��;�!�d�!FqV��V��IH��HZ$j�!�?_�X��a*�A��UII�6�!��J�Pda��?+{ �K#�ſV�!�䘵W��X�p� pD��/;!���!3���,�ULXvE�p(!�0vέ#��ʬmP�Sg��~�!�d"o�����ơM$���!_=8�!�dX�NB+�/��[��	ӀaI�Ou!�(���j���b����m�Ai!��A�g�x�� 
-!frmY���IT!��`�X�'��bl)H���z�!���$}�%�ł"Y:(z@/���!��R6@���&�A��p��G��)!�̤P,4\�&��.}*u9D��UF!�dׯa[�(��ڛZ�N��dfO7)!�ήRn�����{x�����iB!��Ĳ:�m�W�@5+g������O<!�$�3ʢ��a_�D���&��>\�!��R )���XbL�0@��SF�}�!�4��*��]�y�l "�M5e�!�;b����LaɉS�F?B� p��'6\�������"��
�K�'�@��u�^7�P��+L���!�'>�qБˍ�L0�ڳ�ЇK�<�`�'����qd� ����eB��k�4��'�|�ا��>6��a�P V/]����
�')�Z��ø�6�� �W�bT��'��U���]�i� �B;N��HK�'�(9����X��� G�G<az�'"�Ei�l�I5X)���ˏI�t�0
�'(۱��U�z`���瀲uX���'�T|ɥ/��n<�( �@Q$nJ6ճ	�'2���S�3�b	�'���"�Є1?��� %<.n{	�'�q!�	&��`eO���9Y	�'�{���z78<Ё��D����'X��+?��(�����l)�'F��1"H���f�Q 
�^"��',"-�@,���j���y���J��� 4�!�
+^��6�KL�,)A%"OdE#�J��nC��P��i��y)��<D�t�С1��q�0���O>�y� ;D�p;f�DLr�\:��ެv?F �ӊ;D���A�O$x>���GH�`"R�!T*O ��ӵX�F�Pq_�=�&"O��[�ʉ�k�ẕ7�
gl��
�"O��v��f오`a��&bP �"O�p�7�ΧF8��I7WV���"O�P��d�rFh�i�jK�Mj��	U"O�1QTcD�|����m_��3�"O�Ț�J"1��Y�f@�LW��s"OBp� ��3�X`��Q,I?��0t"O@�� �UU:��A#/�ĩ""O\94�(i�@� L�"�4\��"Ov� �� ]Hظr�ʺ*�cb"O���_���gl]�;��ɀ����y�ߝvZ��W�28��z����y!Xp���Ub� ��=)�'P��y�
X:h��q�~j�\A�	=�y"�W����q-za:6�ֈ�yT�pG���wu�F
\��y�� ����mj4Bq!�����y"i�7-��*#$Ƃc��� 
��y�V,'���Sk�	a>�h$a�ȓ5��&�ˣ��m�E��9���)�\���&ʠy�(i� rk��y�o7i<#�'��5?��!��y�
��V�xrLA�4Z�L��O@��y�&�Vb�@*D��&)�޵J��)�yb�3h�餂P+'nIJa�ף�y��۲'��-	���i��*F�y�_�P9� [ (g�@+W$R5�yB�H�� GGP`�f,�rm�A�!�$��[Ƹu�e둱2�J��İ]�!�E3S�<�c��K! Y"0�P�p�!�Ċ�P�F�b�nI�G�2X�Wٳ]�!��;�h�bo��8}AgAܝ&x!��<# t�U�'Q�ơA�3_k!�T2Q�uK07�
��@o.VN!�zBLeS�%X�s�*���gU�5i!򤇜C4�Ë
A�rak`��#N!�D�xOx���F?k,i��W>u*!���89Z��Ğhj���
��E1!�d��[��uH��Ǉi,��۲N�s�!��?t$���_"�<��!�*z�!��J>A���ր�1#U��k��!�d��7V�ip&M8N��R�T��!���$z�~��ҥ�-k3d=3�F�'�!�X�pRz�qC��g%H�c5�/*$!�d�ʪ�Cd�0�A"�>`�!򄔼W�MZ�EU#V���"#+O�|�!��V��bF��B�4���D�-�!�d�z��)�͇i�|L��[>1{!�t�U�`�c����tذ6Y!�d]�/aH�X�����Y��� p!��76TX�Tk�������	G!��.m�<��s��<r�"��-J�G!�M�.?�� e$��|��`�Q, !HU!��_<^s΄2g+[4�t���G�!�؟
��)��`�"S�4�svE8�!�V@�ܬ�V쑟vv�$�A�A��!�͢j�v�su�_�;a���wb^�V^!�$L�w�ƀX��9L�U���ǲY\!�� 2�!BGa�&pJӭ2+���"O�둆�h�4��#��&!�]Qw"O̘:C�T�M� �]��d1�"O� �'�Z�7'<�QF];�n`��"O��R�	��M������6��q`�"O�:gB�	�PK����p��x�"O����*�LYd�Z�`�ņc�<Y��F=u�Z5�2�>����]�<A� �u��]K�֒�	`�n�<udО50�3Ƌ|�QQ�"�l�<Q�	`l�ȉtA��fE
��Ȁi�<�r��&��	cܮ$���nIJ�<�kV,Ye�����������Vk�<��o��T1���1` aE2T���ꋽ=��TRs�դNk�1�V�3D�DA��L�] 
 6���Vd���0D��Ƭ��G^�M�!mͼI��Iq�0D������&L��s$�*R~ta3 .D�,��O��w���#DK�B)rȨ-+D��0R�ˈ.wX�Ȅ͉�Qs:�Be'D����Ė�!��4J3<�l2��!D�hi���H�u/;,`�E2�#D��Ȅ�B�N+�q*׌�7- �hc� D��B�	h�Q@��X- Bd[��:D�hP'#	$xlA�NC�4��@:D��ye"��.�v�`Q	ǜR�ĕz�m7D�8�6 �6&��%��iAL��fl6D��JQ-_��-J�Lש��ux��4D���S�� JX���V%wb�䒀,5D�D�P%�X UC���oZ��0�D3D��X�L@�#���Qb]�m������.D���1H!<��\����!Ȑ�W�!D���T�̒g��¦3~CX͘�*O:�+��\�RDp�
t�	9bn�5I�"O�R"�P%��B�a�"t4��"O�q�G��vL1 ��C=D�0�"O!3dH�z2H���_,~2��Q�"O��W��s��U!�D_=nn�k%"O`|����n�ܑy��O�]���1"O@l��.�1:x��p�ΗGر�1"O�5��I��U���.K��M�$"OԱ�r)$'i4��mB%G`�3"O�(�O�D���C�R�|���"OJ�Ӓj�o�^1��`Л�0��"O �g��R��<(4i�)Ъ�yRł�,ټ��l߅_6�A7!�D_�>�Q�mO.Q�~�����2!�$Y��`�A0�Rz�X���	�/�!�z؉!��Ӱ����f��F�!�ڪ�n���L.K�,�K��'!�!�W3\"��ZQ���.a�3oM<"�!�D;����,S�|�t���ܯz!��(V����R�ި^꼵�ǃ*	=!�䚌K�l�+P�H�@:�8�(̐LE!�ގ:����F�ȜZ7�|�`�Y�'Z!�D�/f���c����!�TG�S!�dW��zH2G	܃_�� �DO��!��ݞi�ع�C��@t1��
R�!�d�<(
��-��D
&hޭ/!��@�e�z	���E�:;�f�;t!�ǗY�f��-G�N��y���%Co!�DG4\�T��!޼{��l@G"=S!�$Z���VB�Q�n��h�N�!�Msi�8����c��E�!�� ���Ņ%!�r���Ա{T}��"O�,�0�Z�>>T��[b�"O@�Ӆ]�]Z��u��3!Gt�*�"O�Ā6#;M�i���=����"OpI�2(�� �VE�0fVH�%�����*����>I�f�'I��X?1C�Q|���A���,��0�3��T����?���-h�(
�7���R��+����`w>������8ޠr��(�X�`�;ғi�0u�2ʑ=���ǔ�X )�N���M�C$��`t��iT���(!�ft�'/������?�I~*�4��4"Â���!�g�r�y�p�'#�'����'&�b�́6AD�c�i�7Ԭ���'���'����A¤�#U������u/
/�~���'|6M�OB�ħ|��+�1�?a��M����>T�r�iTOT�KPB�u+�J��i�v��f����V�
j�LwYe�/�l��q������EX�bq�X�c+���u�gӲ��
��FZ��±J�)#���ഥN,6�",�~��b*>�B�� '[��Rc�-AAB�l�<B����Op=�����ix� �/&��`�%�WM<�i�'��U�hF{*�(i��>�83cB�j������M�7�it��ݚ&��@�]�ݸ��ԃ�T�����?A�ID�Ux�<X��?���?�7_?�m�*��\�c���[�2t��
{W�)��-ϸ	���F���M3��1U����G�'&i��N�977Hpڴ"4n��{"埆s�di���%nD�kg�%���V,V���<)�0w�j=X+M.����ҧT�2R���%�R�'%N����$�Or�B��x���OxB�
�m������IK�'}��`V�6|�|ًT�Õ'	8�PקC����	o�I=��I�<ѱ#�s0��R!`G�:f4b��4R#~�bM
��?���?���q�V�b���?���R`�dǬ#!d6�&���I�e!�,\#�q��H�R( s�V�6�#?	��ݔpܜ �ιo4,�+3�A M����A�#�0L�\���ǈ�-p��|�#��O87�ծ���8���Z��\���6�Z��I<���?��*��l×��17b�K�Dd���2�\���	�/"�
ͩ��V8p�X)��ʚ`����̦9 �4��d�!��l�P��J�$�8]�uFbS(3���M�8�@�ץ�O,���Ov��nI�C}~źe�Z�h�Bj
���eQ|&4�ƬB !ґdyEz�h��rAv)��Fި9M����O�+ �ة�擭E��5Z�bP=d�&� �gW�"=���V�(����M���	T8w�u���2 ��!c�L@��IRyV�b>�O|����5g&��f�LWdP���'��ƃv�J7EU�N�#���N^b�Q���*�Pj�4pi�TY���I��	t�b������o��pW������\¤p+�n��E� h��մ@(E�&L�# ���{�-�+L8B�n���O�kL=L,���AdƄid@<�4�rE]oڲ-��i!å�<IPջg�Ǡk�:��N����5��V"R9vuY�!V;(X�}�ӁC��MCT*G�,�I��M��߈���o�����cD�U�Bȉc		�~r�'7a}B��re$Q
f��"Iz�����O�~�|�gӰY�~
���u�A1Cq��C�Cv#̥���}>��O����+� 8  �   6   Ĵ���	��Z�Zvi��:+���3��H�ݴ���qe"���@"<A�iB���gC`�����Q�R�y��U�6��7�i�X�����f�TYؔ�.(�r��j�j�ቄ@2�Г�i��̩�+�>8Y�A�Ϭ\?�Y�.O����I_>7r�P�_��Rs.H=_��8�>�@��/H^.Mr��S��
�r㠞�?B�r��r�$�	�< �"{������
���[�$z���SF��F0��&�� �x3D��$oy�M��Li���R��8���4@x�'��Fx��Ba�I9Н�s�a�X�SE&,T��	69x�\��ቱ�PH���>��8[��P�<����ď��O��	�O��ҀK\lQ,��	x�N�i1�>��-tB�� ����^-:�0��I���!�a|���������O�H-�'!y� bf�T��jԋ�st�O����d����� a2�l���S.e�P�Е�	�ai�	9NF�$!7���(]n����@}ƴX��`��G/"�*��Z$�O�@s��;FT�kS����p��J�V�
!�<y��!ϬOF	�e���Y�I�(�n<b��OR�����Z��ē��D�,Nb�(jB�K��P��J�U��x��J�G�\Iml�D�9jE����'X ��j�-߃x�	j0��n�Q,O��p�O�{8�'@ \�gC����axr��S�P�k���U��C�P��s!C~�<CI>�'yQ�x B����W*W�~�.��"E-D�蓇�   �O���?1���d�O�Ȱp��'r�L���X��Ȑf5O���̈́�2e�4�j�~������`��-D4�c�b��\G�q�@��(�`T�I���	����x��yGeKT~���S��骡��X���O�A0�]��ڴ���y�]�Nhڅx�.�t&	��*��y��'M2�'���i��I�IRp����O�:y�4�I=b�J j!M�^��G�`y�O�r�'���'$�a�"G%��rlÔeNh���^U�ɤ�M���?����?)N~���r/�����ڷ��gĻF�LZ(�����O��d3��)Ò3���g���V hF ��ހ��#�~_�	>މ	�'��T'���'�ZMa�"��瘼CWvd����'t��'B����S�XٴS�x�Y	�̉%m�oz���@��8��!��*ۛV�D�t}B�'��I)LҡP�eP   �	  �  A  �   &  K.  �4  �:  )A  kG  O  aU  �[  �a  *h  kn  �t  �z  Ӂ   `� u�	����Zv)C�'ll\�0Kz+⟈mڃ	g��,Q}~�D�\Kv����0MX)���޺l(nIe�ڐi��q���)�(Yj�J�����/�T\���z�8ł��jHp�RíQ i��@�4������'��k�)/lm��� [ᦥ�׿��� ����D�`�	����N
�u���
J�<����E a�^)��V%�U[&L# ���޴zc����?����?y��2w����IJ%4ȘA���݊��? �ir`���W�,�am����ޟ�I#+	r�r$jV��TA5��(jA�I�8]�ԕ'c�"�=c�����D���%*��s �h'�ɋ=����L9D����_��
�a	3\8٠d�>�'J�O�a�Ū�ēd���^_�<<QFg�4S�I��Ɵ��ן��	џH��џ@�OS��]�8�:����_;��X��F�~����O����OH�F
�Vl�p�oڸ�M{�tQP�3�m۪2�B��P��؎�D��ȟ��B�+�I����,͜Q,�l c���TCz��D��-:�E����t��l�?MC[w��Q c�E�T��q�����@����25�)R�ӎ�C������;Q�ŋ5E:@�b냮R9��@o���Kٴ2כ���l��BbC�&z0�cr���h�@0���A�.�FMa"�r�(o���M'�F�
~�0ѥ��C6Ds�/I�M($<;s�ƾʄ�j�_�6�x�
ó;�|�po� ��43כv�u�E��@9`,��'��%^q���7�����Z�>#��4��	���K�U>�Ib#��?Gb.�Á H�?ʴ�3��]cp2�T�f���B"��V�<!3��]�NUa޴(I�F�u�t����G$�l'����O8��g)ߥs	��KCZr�<5h֯1D����L]:�d!�`�ˢ5�t��5D����푈[�6�qĬ	�&�hY�P�?D� �f^8�H���G�_�X!xT@)D�`�4�ɹg��y0�C�w�PA8��'D��H�%)nI�w�^	t'*�x'�%�h�,�E�4H[�`-̴	 ED
!��)4���yRmBpT;q"����:vD8�yr�]������G�	V �u�$�y��>;=p$�ӂD����
����y�G1J6���2!�*_�uz,]��y�D?[���E��,L7��iP��?I��Wg����l��se�����Ul�
�)xS�2D�� i��M��qA��5��	�_�!�d��^�
�0c� -����{{!�J�!�6N2 �2U���4s��5��Ig0��TN_:�v���/�Cf��	<������ ���_1<�H��'/Н��AH!��Ύc����Aǅ�� �ȓ⤸a��- �����ި*.jm�����#lC(p��=�U�S&a�`���:�Z�Cq�,��!v@�$o��h��r�4m��k�>F�~�ke(N�&~<����/\[��cݴ�?q�$�\�QU�O����'I�( l���?AB����?�����@�	}�%�����	
b�h�f��P:1
��čC�axȧ2@A�����d�?\p~�C�cߩB3�9���\0�ax���?��i�7��O��Ł�6r,*|
�,8�-�a�<�����(�Vp瘕,E^��V@[/�D%�T�'����:dp��� �?�6�؆i�.�B_����������Γ�y�h�,1��b�kϼh� �KSgJ���H�r�s�{��	��^��%@�[�9��d�0��.s��&R���s���q�1ѷ�@�j	ұ����!p���.���	ٟ8%?��|Z�Tx������
�q��(�Y������!@5���%(�	fqάk��G
f$֣?A��%�:��A'�9@��s"
�S��1l�Ɵl�'\uId�O�D3�ĮO��8��ބK���B��$ܐ$�'B�����Ϙ'�B��'��]��
'@%|͞D:oʑL��ɜ:�(�RQ�,�3�'_� �A`�gj���n�3L(��8?��͝��p�|�����I�`ah1�'�R+@MH'�qHb�ȓ��`��)��F02�C�z���'5�"=ͧ�?q+O�k2��kߤ��bmZ��@�����$;�OH����$>�:��E�����9��
�!��?´�Ic�\��y���҄L,���O��I#f�*IQ�݂�C�Q��@��@jO�ԫ��_�r2QE���/O��w"O��1v��[���*� �=?�R0�|2�e�|�OV}�S�d:/&���ָ� &�lTaxlJt�v�	5�	h�� �9��m[0���ˈ&vyT1+a�'��<$�C�e)�!�O@��RCΈhG��A*D)=bX}Y4�'sDD;��?����?�1�� 3v�!�C�Eۖ��%տ���O>㟢|���E�n�t��5�*�����}�� `�bzl�F��eJ�bP��>�b���vy��/"�6�<����H��}>ف��B�Q�% �� � Pc�O��$�:"�Y�C�9Xh���B�	���p�&5q`�N]߬�󁒟�qF ��]�4��t�O	��a6��9E�RY�
�S!�E��O.����'n��T��Ш]}PU�H�T)j�j�0
��'7��'a��c爼aZy�`L+ $�"���Qb�O�i@���W4^��cc�#a��c��K�򰣌��(O���v�_8��F(_&,��"O�!�'a�y��&��	
�5P�"OJL����@`J�Bŭ�z�~h�@"O )bG�Й�1�r�?��=��"O�cU��5�A��
 9I�PQٖ"O���©9�,U_|i@ i���Ę�j�|��x��H
D��@1�1���y҅00�6���+Y$o���$%���y�/YJ:~�` �����T�X-�y�i��ɪ�+�;��Dl���yR韊3�|���啈��)8��ҍ��>�dr?��D�w�b���A�����p�<��m�&���̎�n�D@*�NOj�<9(�<�8)���2	uHD�2c�<��d�e|�@�޷WB�0����a�<��@�/�R�BE�@>%K�t���^`�<1��Z4[�� �WEF�k蜂� �R�'�rUC��iýe�PY[AF�pM�.ܓ1!�D7�Z��+��"�&����]#!�Ї�-0TeP�����0'GQv!�$V�W���F�0p�Փ�^&P�!��ɼF�����(\$ػ$���!�Ϡ)?B$ʷ�KZ�͛a��̛�O?����Z�L��%���1#�Ժ�v�<�2�Ɣ:x��fZj!Z�d�r�<	�+�$xt}���wz��mDk�<q�K"�n@����:1:`�n�i�<���2ђ�1�J�+}�ЩP�@�[�<Q��%$]��3!+ &|UHEx���My"![�p>�m��	�t���[	 ��0P�ȝB�<��	IH�&�	Ք�PG%_B�<�`�S:d�
\k�Aڬ,� h賬�t�<��B�3�~e���a��qU�Z�<a�@�Z.������L���!/NLx��P����,���AT�0сG�9[���k#D�t�RK !x�
d�4��:�`6�;D����d_I�$�h�b�M̰xm:D��ar��%L�ز0����֓�yrd۳#$��3!J�W���Tkڷ�yb!��X�К�.�ְE�� �1�hO��3T���8�(r�O:)S\�Y��Z�X��C��('"\PP� <I��VJ�$X?�C�I-S�mB��C������X?$C��#'3���@��l$�[!+�*U�C䉀\�>M٣-�%��r�#�B�	�8;b��1`�.8���0�NPz��ęc��"~n�^}�Y�Ӈ霽�7�F\T!�dlW<���!�J���[^*x�!�$˵Nξi���P)!9��`	�5�!�䃩6u
�������0�$�K��!�K�Lzh���2
:ј0b��!�d����I��8��tb/%�剛:� ���V'[�P���Ѻp���`�R*~!�� �āg�	�bR�yC��ϻ�(�e"O�x)�év�~tA`fW�"���"O���V��i& �� ���#�:�"O"�󄬗&)!��a��A
 0MY��'�����'|�5���3L� a3��#�����'��a1k�UR��ŭL�	�2d��'x�TA�Θ	�5��&Ǫ����'g�93� �D��J����~��s�'���	�FUq=�IK�V�-��X�'!ֽ�A�WS�|�`jS����%o �~"�i�R��\!��jr��O�X�<yq$��<?��Raυ�-��QyAAZ�<	��C<G~��w�O�=f<�_�<I�G^�aNF�۵��z�J�P���b�<QW�� s�ʑ:�拜�,5Ȳ��g�<�([�!ކ�&��8<�'$���h��'�S�Oe��s���,z:^@bF�2٠ԫS"OzLqc��1�\x�GA�Q�0U�C"O�|�a ���	�+����b�"O:�Q��
h"f=��j�p�F�4"O}�&G:EE� +��1,��P"O.L{E�3�,���B�qŎ��@[�4H3�;�O��KeL���\@��&�*�8G"Ov!����x!4%B����nu^PC�"O��H)U� `�Q,&pb�/�!�@�7�r i7�ȶhtVM��:Y!�D��v}�ӢT1lv�I���#P�}�K^)�~�H�����.��f`H�����yB��ot"��=OP��l\�y2�˓X!4ZR��98���,ߦ�y�h_"_���j
)zi�+$AF2�y��
1f�6�-hmcuCǅ:��Є�X3���"*W;{��9[�NU�hD{R�	3Ĩ����e�ڄM�"r��K����"O�i3	%# ,=;�oG;��X��"O� ���5s���2��V�,��"O��ba⍦O%u6�ЏP��@"O,�ƃ<R�p=�$	n�x�*�"OZ���ž<��d��=n���T�'�0����p�}���Y�~X��D�KOl��ȓkB�6F��&����#�u��{�ѓ�b����&Ř�B�`͆ȓY�n5��^�8+H�@��K�b�^ �ȓI(д0snaŘ�PW���k�"���~p���@�0avX��
��Gw,Ȕ'<z$�
�7�B@JR+?`��+��$FT��ȓ+�H9�7��HЃ)�%I)01��=	8�SGm�2P�C��ǅc��=�ȓrh�DjB�5è�A�Iͼ�i�ȓ=����4R�SGJ�@Vh���
?���I�0�z��'�Q$ ��z� �(�B䉌D����k/Z��P�a �;�C�	X����LC�D�Fpx�'��!*B�	 M��lsׅƬb�t�%M@4j��C䉒$���x`�[�@ߐ��s
ܼzYB�Ɋg���+�n��D
~@G�
]�2�=1G�\�O�������)@
��UKR�om�Er�'�b����>R��
e�ׅ�P �'L>uiEnʶy\��A��3
�'|eH��ǉ8�J�Y�T�Y�Ah�'���  O4}��[7V�;����'?�1��l�T�;g��<�i
�o̴Fx��)Ī4+��{0i�o����$S��B�	�I�0��)L3	;�)k� ?4�B�)� �ųW#�?$�i�!��2"Obp��h�m�
�j �*3?B�"O���&�E Nst����3J-��g"O�z��N�~�,`NA)"+���DR���E�?�O<*�.��,,�%!"��?��ԁ�"OP�94���V�`��`/Z���Br"O��i�kW�c���"�nI)c�� ��"Oؕ)�FՎ~�N���gO� p|-�a"O���ŝ,^�d8��ra��/��}�IІ�~���8�����&U���{C�κ�y��}�L��� A�n�Qo�y��Q)	�l�G���>=¬�q��,�y2e�U���ōǏe�.tP�i]��y�e�2{���aܗ_�8�H�,�y�Ț�\Ъi�g��shM@Pg���hO��IQ�S� ��($O)%E ���(�!|C
B�	�d�(�bMG�n�(I���R�a+�C�I<4;�1dЩ���bO0!��C�I1}.! ��F
�bj��6j�C�I�]n���u$���a��;�C�I�ARD�C.�'�puK����Ԛ�Ě;A�"~J!Ձ<�|��!<aVf��C?�yR��K��$�����"h{DF��yb�S!}�r�3P������F��yr���
{�T	�oY4L��,��KU<�y�B�i�\=���H�BQys�N6�y2���aj7��%952ypc�J���DIi�|ᐊG����p)�5�LP3$I��y�
��/@9�0b�uY��"��y�FH�$��ȝ	hV�gX �y�΋% T<���m��M�2] ��Q%�y"
"+�8���7�� 7�J��>���s?�i�C!šP��F�Z=���]Z�<���,a�<-BEn�?D�qK�SA�<�'̀	gtH�3�.Ͷ%K�� M�@�<Q�-�yЦerƙ'{�4��vNWd�<I��p"X!����}�qhL�h�<����L�:$�UDW;*�}����M�'��Î�)�G�	��O^� |2DZ��!y!��0�
� '��� ����gE?-v!���p�,L�E�'@��	��nÌ{z!��s���mGo�~���BQ�2�!�ɵ�CU�ܖYp���E23�!�$�_ ��Bi�_:�1���y��Ϧ�O?}�p�J�`�P��^5O!����a�<Ѷ��3��7d<T�B!s�"�4�y�˴/'�1	ᢞ]��t�B+O��y�O�n��s�-�: ��$1����y�C���)q6��a
(�Q�y� Аs�Fy�uʇ���0d�)���`5�|BhӠc��U� C6(n��E��y��o�D��("1�XG��8�yŋk9���W�i�d��J� �yQ-^v��Cр�d�>)r�^%�y���6��� �e�<cQN�i� ���>�s��a?y��Т6d��9s,�����]]�<I�$�I�.=j�)�+&<�'��}�<��M�a��a�$��&oش�Q��z�<QS-L�Z��5��nH	EP��2kRa�<�G�V�M~|QB���z����f�D�<�e# �5���Ɔ[�;����}�'�$�����t���`@x��d
A˞�h:!��=��q�酥wq0$��	:R4!���X^8��L�sdTE	�!�!�� J[E�H�
^ 3E�] SV"O���'HX� aef�w��	h�*O*�p��%\0H0�,L�9��8�Ex��)�;7S����! 7��Y��k��B�	�b5�4�كfǨ�����5woHB�I:��BRC� �LuS�Z�3>B�ɿt�\��Ǧ�^����I B�	�Y�`�u�kA����n��C�	�hm0�����KW�C��@�F��˓P�Р�� J$���ρ/�M"��D��C�IX��Bd P�E<���Rh� E�C䉳��� ��W�b�`ș NS�s��C�I�4��-1�m�6|.b̢�+;@8�C��,T�����L�(�#qcU�r������=_�䌎�f�u�Dv܈���o��Lf!��T�x�4��Lm�9S�[�,�!�]�0<ܝ�� �M
� X�.T�!�d� �Yz���jL^}��@��]�!����s���(� ??'�D �����!����*p��w�����x�ў��A9�'
I��c�C�O��i�'Ǆb*b��U1�YU���
� ���=��' �A+�j��9�J\	%�V�-�6D�'�|ᰒ��K�1�N '��y�'�rt�P�UT1�Cğ%|h��'����̓8��Ek��F2�X�� "�uDx����A�<��!�A�|%�԰�@���B��%M��Ha���W���p�͊R��B�I�B@!r��U�?���1�˷-��B�	js䕳'KʥPU����Ȣ9@�C�I0Tv0i$(I�ر�4|j�C�I�'���Z�g�p�\����2)M��	R�d:}2�_�@�D:}��A	i��!��M��,DB�cN8J�֟���֟h��T��PP+˷;��ՠ��|"�DJ�H�\V��'a9.�����S�'tB��!�����7���r�Ӌ@�prB��P�YA��:j�>">A!��ȟ���F̧
����Q$ǐ����f� ��'a~RǔK-���b�J$>��z�(!��>�W���!��l�*�x�b��w��-:U�<�a��?����|R���?q�J�):�����@�98Y��A�?!�ׁKb8��c��Hpl�a������4�lKk�XR 	@�Y��i��:Ohe>��T���8�J�&��� �z��ԅݩD
�\S�nC�<1P�՟T�Iy~J~��O�q/M�H/�\�!�Ϋa�dE��"O�`��䄁^r>5i) �	�8 �s�	�ȟ��·	 �	�v%�$F.N����O�O0ʓ=�R����?����?Q+O��@�H�׍�2
�X���-���HWn�OX�2FV�%G�P�P�?#<Q���|O\+C!�=��2!�h���{zy��U�P���Oh�XU��G(�ÅI�*j��P��L���O0��4ړ�yR��Q��``��=�>0 i�y#۵�*=2��\0��h����?a��i>��	^y�#��H�m��x�C�DZ�����D5�"�'u��'��)擶:~<تCE_�4-K�+�d�~$I���U"�{P��+԰Xpϓ}{���\0 (�H�%ϒc�~`�ą,�F��5 � ϓ�F��	�7P`��J��a�G*a���Ij�'�����ׇ6lx��f2{A@�p0�8D����X�Y��h�3.
r�$��%G�<)U�iP�X�,ŭ)��O� ��Q�f.:����JD�`M�R���I����F���=�j �!��?�'R؋�<}&�P�%�7���D|r���L������ �xԜ���T>�ae�Вs�� m-�E�#!�6�,��͟��|�D�� # P�p�X�G����Yy��'a|�C˻B
���ր�05#,	�� ���>�T�ȳ�	ٷf/�ah��|�hI��<Qr��6=����w���|�T�O��*�'5G�T ��Y<Wv
u��۝�r��8�B}r�a\\�`m��	]�W?u�E)ִK���%P�'2�Sp�l��o��qܝ��#3�R��V�S�fߌ��Ѡ�	ւ�h@H0��	�~r�'��)��%?� �m��攏j�8���Ϣ�"��"O��+��$#� �`A)oE>bC��6�ȟTQ�U�\�T��Mep`E����O���O&�P�$R93}^���O��d�Ob@�;�?�,�Kݰ\P�&Yl,���-V�Z����'9L%�5�	/��KΟ��R��λSs��R�Y{m�ȉCƅ6S�0 �I�L��Ԥ�(,��g�'�k�ę^T�n#a�n�;M ?������L�'0�dU	5:��/��$��m��13!�I6>S��&&2���2F�=#ª/��|j��':�i���c�" 4dV7�f0b����Q����02Ijto��T�ޫG�C�I'!"x8��^*)̖ qw�$£"O�AXw�>4(�����YfBh�"OX��� �<uh��W��:N��!�"O�	�G�6>j���L ���I�6����C�')j�d����1���A��}hj�F|�y~=E�dE���A�cг~�Z���$ňO(<Z�G_*�(�8�����0\�ӳh�Ew�-+f�I�����O����K�%71�)�!oQ8/�����O���?�)�8�,�f�M��>P�S�@[}�i��$��	��PA�Ռ�1_%��%M�;
�ʓ�?��?��4��4y���
X�qq#�)�I9��(O��=Q���8|>|9�!�@0;�pB!Og��L(��%��~��1@t䲂#C* kVt�`o�H~r��P�`�=}*���D�XĨD0���C
�!n)A��N,?	��>Q#��X��RⓡS`L,���)#�ʙٱFM�41�2��>��O¢}Γ �Q��A�g5zH)Weӟ�B8R`�b��`���o�Ӽc*>���A^;#O�5bwOFAC��d����� G��)�7����ҰX� 0¦�� P��Y ��7��	OÜ�'xH6��+y��X�%S2J^��S���?��I�I���'��#�a��Y�<��҈��t�`���Ï3�dV�F��S��'M�9��O|����Ĺ|}"y� l	�NQR��@��-��I�����#}��i��8��L�Bb@uX�H:�N� ���On�ˢ����<�&�]?��H]�W���Qa��Mnm�̎��` �'�0A��-V4,C(|��F-l��y�'@\�aeƺGB4x��Pì�zݴ�?I�����O���|�-��9����Q��GZ�:i����Hh}B�|�U��G�d̖�K��U
�M`�`0�����ē�hO���	Z�)J�T$��V+{Dĩ#B"Oh��R�x�Hxz��B-D����"O��{G� 2\�T�u�1��`RR"OmZ2� Mڶ4��%۽OV�q�"O4�Yu*X,ЎܺC�\�2U��h�"O��EJ�;�x�g䑸4F$��"O�)x��JG�ɸ���A<�%ȑ"OJK�<9Cʌc��E	��h"O����@	f���6A�W�
w"O�E3�G�>Cw�+�oÌ���S"Ox��P�VOL�%2%�P�qw��[�"OH8At�r��8:�ǟ�=fLՃ���){tމHȋ�	��	te�Ro���f��*��(sa(�/6����!l���s��9�ʨ�#NL��~�	&!�I��.�5�,$��k
�&u0�B�#5�L@�.�,C�`T飭��8s#(�2�����E�0�b�a"�� �@4��O�r���� ��A�I�PP�c�B����W��(p B�ɭ/x�����/"��*a�f�B䉉~N-��HA�\~` �T� X�B�f}�m[�d*ny:�C@4K$�C�I�u�Jy�$Z�48��[�� �~�B�	9z�ڤCF/�{����H]2�B�?kļ���F#8�X��_�@��C䉳`X���Ɨ4c����`&j�C�I�rSV!��аo��	�.ҮC�I*������:$ZՈ܈t�C��5@A���{���@-ۺC䉳&����f�2l�EG
�8�RB��*	U��!�Z�/���J�½\�B�)� ��:g��/n���{��/�Z�"O�<0i܁jw��Z��"jZ�e�"O�q ��n�� r�=8G� k�"Oxe1���]�M�!iۚQ�|�V"O����b9+�"԰ŧ٠4��f"O��a��O�C���gE�*H��["O
E!"'5�� {��?O@a��"O �����1T����F5=R����"O����.���v���?�u9$"Or�p�E�L�иZ��,���"O^���ON�HR�8 j��$D��p�"OJ�`��/&f�$�U��%'@(Y�"O<-���6�rI�Q��97G���"O���0����%�!jȋe����"O���҆�g0�]��1o�&��6"O��vEB�1�P8��6ޤ�j�"Opйp��D�b�@S��	i��`�"Ot83&ʊi�-X�.�pZx���"OZ-�R!�V3���mKN6i"O�ă!�L:pC�તm��G*�e"O��2`�P��s��+>�M�"O� aB+�[���["̓t�v �U"O��T���h�H��-W�R��t"Oha�&$J�!�報L��]����U"O2p���͢IJ��n��3�X���"Ov���ƁZ���Ä��z�"O D��C�����xd��6�� �A"Oa@�>����7TM&�`G"OP虷ɞ�d�u���%I���6"O,�۴�([5UI� T�"E �ن"O�I�V`��q�������q;��"O�`IZ
V�2Y�C9eG��0u"O`�I
��vTHR�YU���E"O�Z�H�T�)D��
6���"O�K�
Y&>��)���~"TQA�"O(e�p�V�Mf�+_�����۽�yB�/J�0��$�&��kP�R��y�✅q��KdB�iߴ��r&~q�ȓ��e�!.��oh���5F F���`i)��. �t�!�ƌ>Q�ȓ[�ڄ��]#Et`�[�
PӴh�ȓ���HG�I����5��U���f��Ȼe�j����2a!�a��P���
n�=Z�d���������Q�* �Uz1�O�o����Gg��fۣn����GȈF$�؇�fa�T�ņN�N{��F�үCo8͇�E��d%�
H���@6��,"�:���@2�8��Fg:dX��[�-hy�ȓI
.h��~�J���E�T�)�ȓzl0��FH�;y(��`�O� 	M0y��8�P#��������^�Si%D�<�@oA�+&��ص�<Pz
�x��5D�\+�o@65&���ȟT$� �D4D��a'gՔi䑃T�^�q���HC2D�cA�C5#Jδh a=�t�E�1D�4bn�'�PA�q�L%, ~��b�-D�|JG�J lz��U�=]�8��/,D��yv�/l�� iI�gX�$ %F,D� b�QM�V�a��Ȝ�l*D��R�E�85�����?Bv(��(D���cD67�D��$^�?�L���'D������Y$8�Э݌j"FQ!K)D��'�ѕO��1Y��Z�m�T���(D�� �	����(�����ڛ{�L��@"O ��$_f��$1����^���"O��S�nȫF*������k�6ٸ`"O�As�H1���"���}���"O|��J=��q0�ȘF�>�S!"O��b',��8P���qk���>P�u"O�DabM�2,�4�!$ʝ5O�x�"Ob���mӏ5�T��L� ��$
�"OBu3R�����p-0~���G"O^y;Ń��C��ԧZ�ΰ�Q"O�0!�a�'3��)�b�J�d�:���"O�0J",�^\�Q�ѵ�\�r�"O&�Ʉ"��4Ի�*�*���k�"Oj�Ғ�O�&�����4+��,9"O"0��H܂Sؼ�P1&�(���"O^�q0GL� �
h��ʍ�~�b$u"O��1�z������s�X1	!"O~͛VjW%P|��$��5�`��"OV0�!�a� �b� "U�1"O�e�"̐)�j�p �!n�L�C"O���s��CS��A����d|�D!�"OT�@R&Sp�Afn�	t�(`�"O0P�m��a=�;��O�5�Y�"O8L�4���T�e��ލn �8��"Oh�R�Ɔ�.]p�3���g"O��q��خT<Ay�:C>�� "OF�����"<萐��^s!�*E"O<����7]�� {�IF�~�Ys�"O���4+��/���%�L�?�xp:"O�Y���f���Q	 P�$z"O�yq�e��B�<�r�M�:��e��"O�X(MK�Mn ����G�� 1"O�������EЎ�q��tYw"O<�y�E�Z��iH1S�CȄ��"O�m�����~4l����3�V��c"Oz���$LL�k�^U�$Q{�"Ot��Q�N��Y�3nE6*8����"Ó�m�?, (�!��>+)��g�<a�J�
W�P�c�Oyt���y�<�o����8Y �ır}��1V�]u�<�%���[(m�,Ħ1D5��w�<��A�G�Xܻ��O�J��ES�� t�<ab�ߓӨ(b� ����t�<a'F��ҬPÀԙ<�n k��s�<Q惒��%B]'4��)jÇ�)@�C�I1E��� ��V�[@��� �׮C�	�kJU;��۝8��(��ћ(*�C�	�hq�]Y��Z~�@	3@�+:{RC�IG�t:4�L�F�����+	PC�I7�\I�����ea���>@XC䉡6l�@��N֐�ڂ��C�fC�	�|����6}��#@���QC�I#g}.�I����l��X`�� �B�%8�2�rA�G��ѱa��iN�B�l��!�q���j��]�����l� B�I��4�CG�tA�f�W��&C�/J?BYQWc�,U��RAۉ{"C�ɢ �4�S�%U�H�
��E
O��C��	�V��g��*^@<M�%��1��C��>�x��̑Y�2�E�*f��C�I-d=V�!&��M�w�P�n;D�|�SϜ�zf���+�0~���Pb(;D�X���ԁT�`(�e���U�$%.D�,��&C�U�N�;%�7MJ�D#.D�� JI��C��� y�i=(�`�`"Ot	�1ܾ1��l�fȥD����""O�y�����4ۢ	�����R�Zآs"OD�k�*@+n՛�eF�S�j	[d"O2b`(�8;�|���G�f���"OBy	�rH=s��v�©	c"O$�t��)� ���X4sJ�y�"O��B��XR?��	Ī�PRb8+�"O�|�#I�H�p��؆��P�<�#G�K�xbCm�i4�� �kP�<r��
uɖ�(�oT�@��p��N�<16I])������D,�Dt���<Bd��Mj慇 	�,��&��Q�<���o"�7(٦%5<T��H�V�<�%�� ��0H�ˑ&|+D��b)JT�<Q�M�N��R!�V]�fl��VT�<�]��R�N�|S���n�5Y�!��4�(� �Lx<�<�CM�+��$Ϙ!�H�
f�ȹa|�Ѧ剁�y�盍���!F�R�r�l{7��y� �~�����m�)��-8�y"�[�Aͪcb��iZ`x�nB�y�j�%o�U֙u���#K���y"&�0"�T�&'r�6�J3�#�yR�Z0�3'���K~�rcƏ�y��_�@I�5Qu��?\N����Ĺ�y�_6/\�J�EF�W
��SR�ղ�y��6`�J�8d �H�BY��y��i��ḁf��?�n��I���y��ѠN,7�e�:|�@�ܖ�y��,3�Nx�T�b�����$	�yR�� W�	Q�Ŝ�] |8s��y���u<��+��Qp��C����y��N-+]��r�σE���
Rl�;�yB�I/h��4�[%if����y2
	z����t��bp��aE�Ԙ�yB��_֝���K�X/�|��KD�y���B���p�O�U�8� �퐅�y� A$r\ki�6��P�b��yr�O8}��@Ғ����Z-�a �+�y���R�� A��/Ҵ��'�������HH�d�V���1�'�2H(�mW25�l�6!T�ֹx�'��9w�l��EjF #J`ȝ�
�'�D���n��6��孕�Ee�@�	�'���aFܥ��0�5FI-p��	�'�:����M��$����W����'�j}�GN� \��@a�����'
�p'���'c���K�+ָm��'�l��,�	vf��S�B�2��8:�'�`@��ht �#Fފ-F� �'�,̃��N�m�  32����X�
�'��a&�,.�ڱ�ڮ+>�
�'&�T҇���&l�{�K��8��
�'g���ş|�}x�ꌤ?��3	�'�H����Ԛ[P�rwa�	)D�	�'!��cGd.n�U�GIθzը�3�{"cT�Jj��+�pppѨB.��v[ ��#�0~BH��O&)|<��,T�Љ�]=��Vd��8�݄�G����#��b0�=��/[z�d��N�B�"�¨=O��1aiJ�i����ȓzXڀJv F[�hIa=ց��Y�fi��
7&���lV��T$��Mqȩi��ێK�D�é�
\�(��S�? 0GC��Ѻ�S�i-d�"O�M��#B)��q1�͙�16��"O�h��U��P�
M"}mI�"Oe#H�e�-�p���;b��"Ox ㊑�sߖE;��nt��V"OX&���t@Y
��D��"O܂B� W�h ���O�k�zI1T"O��21nB�G�C���8�d\�"O�m��M��E̔�"��5���d"O� :V"����2V��]��M��"O����؆}r�ZA�\)`��yc!�d�:ٚV��c�uRs��vS!�d�4f�`i�4�ݑV����N��R!�E�hy�X`�#E��L����͍wL!�dSC��H�c$a�p�t��D!��י;o�		����T�9@�Nc�!�şg��:�^�9`"y�$ {�!�$�����Ԡ�)-B�1�5�T�_!�DV�F���k��90�
X8㊃�VX!��%/�L�Sâ���`ȺШ�B!�Ĵxt��։Qv/��.�0A!�$�2�DE(#eФB������!�D��+ʹ#',9v b��K�g`!��h�6���DXnI�c]�_V!�D̗h+�l�0	�>K+�{gB#�!�d�V'�$��e� w=* ��*
/89!�d�{�B�ѣ��>v#h䂧�ڝ
!�õAx�ɶ(B /#��!��"O�iJ��;L ВcCN�H�~}!W"O�h;��E�hs���Qb�//���J�"O��`Q��KGb� 灀(?���+#"O�[���r�%�p���B�`��G"O4Q�	Į�&�K����U �"O��a��3��	���fΒui�"OL���ѵ@+�!�!�M�'��l�"O�!9���N4	�G�7�
��R"OdayIB.E<az��I^R�RG"OAK��C�;wp���� ;A��p�"Od�Z�:��m�����6�ޜ��"O��3�Y�L���zu��/:�,A�"O��"�@�AF�:���%}�`E�d"O����KΖu;^�۰gP[�pIP�"O��3e�º>���j�/�0,��H�"O>8� ��2�6��!Qx��p�"O��g�I�#��P:,��a"O�E�R�_�tU��T�LQ��< "OJ�aA%��1 H2(�'/���5"O�T�O.�t��'(�_�hi��"OB��1�t)��Oϭ/��T��"O�HeOG6� ��M���@�k�"O�y�r*C,q	��¶U�_�Z�Za"O��@R���Wf��C�
�$Qb$B�"O�țAb��yߊ�p���C�U�4"O؅:#�
N�>H���A"-�"O`4H�J_�X.�)P��Z�����"O��1�8gT�Yɗ,܂8Т�"O�S7 ��� 9�m%*w�3"O���DƚN��q�l��,�p��"O�I"�A���L݈�cמ����6"O�8�q�Y���b&�M�s���"Oz��&+5��+�AP:H�yw"Od�Y���6%JH�G��P��TA�"O��&���f�N�R��J�n�bI�"OJ����Δk�*=c�Eּ<`st"O� ^�X�M�/��9y�KX|Tɰ"O�X�dR�:R��2V��6}U�*�"OZ�zGC��'ۂ\�A�W=(C�@�P"O�p;VÂ���� �͉G@�T�"O��(�V���z#��.�z�a�"O���ӧÝK�xd���9���!"Ot��d�-w8f�ŀ�!"���/�yҫa
� ��jQ{���o�y"�Q� \xZ�b�.EC��B��/�y���>Et�2B�H{�����!�y�(L,	g=��o'v�'f�y�c	�RFiR�۩f�ؐ"S�Q�y® "@��@8!E9��S�mA2�y�`U%NX<s@�O>R���
�y���f�j�R��93� ��'R��ybc s�V4��BX;~�*阴�	��y�,^n��$Z� P4���y�֊4�v�:�C�� !�)·�yb�Ƶk(2�{�зw������ybm�2{�A�S�."����W�ʌ�yr%R!4-�#�/7]�De�sę��yOɅ@��T���C�Je�;�G�y"HBi�Ҥ
L�D�p:��T��y�'U�1C���>�6�&���y2� �0�\��Պبq�xi�A���yb�I�<�X�+sb*g������y���},�hx"�N��%eK�!Z��eWHT�eR�e�h	�B�OkBȄȓ
*~�p&��9FB�bt,�V����ȓ*����Si�"딕����^̆<��/9����a��@���i�f��N> ��McD�K'17~XsdV�љ�'GU�<��i@H!���)(�x$�Wz8�P"��Ұ*���*y>����3F�!��(Jj���@zЭs�M��I#� 7m��/��������#~
u��Uw�e3��FP40�Z��s�<���L$��em�3P5ڜ8E�
��̕Cv�M��0Q�ݩSĨ�&?�4�E�@�Ng���!EJ�vJ�*w�2�O�\h�!R���	Q�F"S�XͨG�!D��#�M�PEn%01�Ŭ��=i1��'@U�$��+%�Xq���Xz�'���:�J=^(K�GҴ�S98�vi�R��y�Zq`1���C�	(+f���
E+h��p*��n���ɍW�P)XE�����t�B�U3r�D�DCe��SV�L���H�.���y2/!gV@��J��	(��z�$M���k �SIk�HQ
&�O�OR|�T	G�E��Z ���",�Ń��'q`�I�BA	��g�mM�����=�b��X ;�`��Ҭ;P�a{�nߖ>ʸh��أ�x|:V����O�l맄�6+a�<h��ׇ#5�m��foݝ�g��¹c��	F���G�*D����̚v�~�h�*
>����#b������U����@�>Q�|x�rn][�O�ԉi$��\<B�Z�&h�Z���'��s�F����[6�1Y�ⅲ�h�W�h��4�	�%S��a$N��g�7�J��4���	t�8s�1O������1�Ɣ�CnΆ*����Ҋ�P�����Wd�m��i-x�
�'9������3j2���l�H�I���ʶ&vΩ��Β��4"�.e>�(�l b,� �d�%����Ѥ4D��x� ��t���'ڬM4l��&��<с�N�(36в�b���<��^�m=�d�dEA�Ϧ8H�S�!�DV^v��8�D�.'� ��4㉁Cmd��a�>q�a�3C��>�O*q0a.[�V�f���7:RD�a�
O8�2�
�} ��I��S4&�����h�+��q��
��0?��f<�F_�\�pB1�CJx��NO�xq�'��Z��N'Jݜ�+F%��J�"��	�'�n٪A�Y�<6��r��r��x	�{�N���O�O8�1��dR�Cɼ��B`ٱc���Q��� L��G���	�Fp��eV�n,�"O�I�Fmߪ0��`�LT�BQ��"O��v)��m��M��A������"On�×���9X�ࣁ(��,B�"O ��$ވ�๻'Á&����Q"Op!L[.Y0e5A�Z���PF"Oള�"6L[�;���6l�)�"O2�Av+ʫ\�bB���J�\	�`"O�[%�\(rVBͺ�B���P��"O*�p!�Z
C���&����T34"O2�pT+Z.��% �n>t+Jy�B"O@H���۱UH��MH�9�T�"O�� (g�
p#F-dyt��"O��)�B]�>����"zr4=�V"ORa�#c�_���T�G=���p1"O~��U�4l��s��*B���K�"O����(��ղ��f�*䣔"Oj��@�^��[���N�ԅ 3"OtM�u��c��1��Ǟ	���T"O4r%o�U�T�AƜ ���!"OD`b4�¸4rF)����V���*O�l�%��;�n�`�-�e�vq�'ᒼC@	4����E쌳i_j͹	�'9���G:/�u/ڈ4G8�J	�'��(I��_\���i,&�r�']r���U�i�D��L������'�bp)�1\�< �h�����'I��)SKO�<�T���4��pJ�'z޽���M�$Z ���˒y@.�j�'+���
�9r�*p9c��q�
K�'4�!�ǵ$�D���Z$v���r�'���в�)��T�+ݐCpj���'�&mJ���#X��1� ţB�<0��'�h��ڴG�E��lˏ��S
�'�aB�E�TԼ���D�Z%��'�aF�>?��X`C��@�y�'��(%�5o�L:�b^>y��5�
�'��Ř'�h�ܰ����r;ڸ��'��P�C�V�'�޸��)cw���'�	���8�ѫ���'��M��')��:0C.o�Ι���Z�w�Zi��'��@�ʒq�0�s5&[�=�� �'���1���@���g���0~��
�'���T(ȫz��S�l��GǺ�
�';�$�B��;�N��j����
�'?ؔ�)�!j�HB���8�i
�'	�V��<�|$R�*�!���9D�� �� ��	Z.6�-���9D����p�&9"�Nܩ.��1�G9D�d������7)Z��pl���8D�<���<RE�����
M��@2D�x�@A�5B�zQ��	=����:D��"��\�x��af�3<p�(<D�@��W��%�R�K2�8i���8D�\�e�P�H��[�	M�^IIQ�'D��2�hA-Fサ:Т�*\�:Y�"@2D��@��,b�9�'%�57n��e0D�ȉ`�39)6u��!�-b�};6$"D��� �47�ipa&ͽe"p���(.D�tِ�Y�-�����O�k
 �z�B+D�X��\�3��D����EB�(�I@��!��
���Ԅ�0M@�ODx�#�5b@�uG��<v����"Oj�x��ѴaQb�˄��A�"O��@�O 5���V*�D\T"O� x0� ��<L4��k�^����u"O��	��[�%��L�n����"O��b�e�yZ����a�-ꮨ�%"O�a+5.b��AQ���-*T�L��D¨@uZE�&��]~N�YA�)D���/O8~�D5ؐ���A�(L �'&D���ҩ^2��"����	���$D�!EN ;a�9@@oBUB�!8N-D�(c�ں$M"����E�4�FPz�� D�ܘ�˙�3��yz���x�H=���>D��B �Z({̵I�aU/F��TՅ D�D���^�/H��abe�'n�р<D�`+C�$R�k7�R1��@���<D���P	օ�@1x7� �j��:D�d��E��2iN���	��a�%O&D�t���I^^u��ט]�XA�%D�(Tg� �bd�Z'>cz$���(D��R�KJ�1����#ث6���pC�(D�@��B	��z�̨���ϓ��y2��T�JA���Je�9HG�y	N�+�,�R��!Y:��V���y2��Ut\)�s�֑R\9lƧ�y��ŲoW�p���G��ɲ����yB'�?_\T`!��C�V���=�ȓH�p]J���uA�č'����EFU�!�F�5��X�͎7�Z��ȓQ2i�7�`庵HA`�,��Q�h<�FU������sYF��M���pR1s�& HP������ȓ#B�U@d�ДP�na�ƨԃ%z�Ȅȓ0DT���߆Kq��#-
�\L��ȓ4)"�
��H��G"�Q>F-�ȓ]�1����=t��N��6��(�����X�����bf�B|���_0xp$�5�P�ajA�`�ȓ���w��!e� 3d�/ �}�ȓkW��Kn�bpР�u �1۠���;�0���CZT`�R��	�����	���ٳe�j~�e`&���)�b��ȓ��ч��K����G+CI����܎\��jQ=M�Ό$^(X�@�ȓ �
����^WLa���Ѥ�jQ��'A���S�oP�����
J��ȓg9P�@kS9�ZA�w)N�M�i�ȓ!�Ƥ�M)���Qh�}�T���o�D\qp��,{� ��EÀF�x��ȓ<9*g''yԐ�;Үֽ|�FфȓS��a�AQ�3�e���2}���a}���ቔ_�P����03
���f92�;dn@�nZ��yp�Z)���y":���K�I�	���j	��?�̼PDGI� ɎxA��#��܅ȓk9z��i��\.$qg��T�d���B�`H�埛&	�	a@	T�����^M郧�mu:}��E�a�"��ȓE�`�1F m�RDce̝	!�Ї�Q� B&���2�2��d,�>%<VT��b�x�SV�T�-pP�j�'ۼg���8�$�2�Α� ����\�	����aӰ�D�B����#Ph_��ȓ��`�J�,͖�B3�³~^d��q�r�hd��Wu�l:�Q!��m��\�#��B@ '00����tȊ��?
�c��,>���S�? x���!�=����F4�""O4�IR��R��"���c!�a"O�!rBb�,=*������c�c�"O^<C�M]���hP@,~^��S"O=*u%�"h4$���Ku((��"Oj��'�_���сȐ�u\v"O�3����!<�
W�gn.���"O
�B�4d���"�T�Wg6���"OLq��c�(Q�<�C	]#Lbī"O����� K�Գ��ʟc3@�0�"O4��cJ�1�dx�p��\��\RT"O�ᴫϙ{�p#Q��p�p��"O�5Ѷ*��{�\x��bHĸ5"O|��S��U�\���"]�X�p"Oܘ8d@��e��"�d��^Xlh�"OL(�b"�w@�����kO�i�"O���S��&A]�|u��m3bɅ��y��Y
+O ��M�6�<�&����yb�v�tu��@Z>Y36l�(�yB��# �4�)gjC-X��B�)���ybOZ?
�DLj���g���n/�y�BǙF6���;
�fY ���y�DQ;_ʝ0sl$	j�({�S��yroɎ;����@�V�*����?�y�/ �M�YC#/ �V�i���y��XNc�!���,���eH��yRϞ9c��l�4L
|iVɘ�j���y"�E�.`����<�P�3
տ�yR��
,g��kpG D�$�7K���y�$Ӟ`9�	x�9H�ږ����yrl�;�l��%	Z#-ʦ��E�O)�yB
��芤��[�p�ԣ

�y�������@j|M:�K�)�y�O`�ހXq 06��uq�矧�y"
s�[r��4x�X
C���y�E�<���qo��d�V�&[`C䉔tAx%qV�@>a:��iUI� @B�	+wz�	�	^�-��z6IǆE��B�I��Bh�!��U>��VC�/B�	�J����60�4+���y��C�	�=���r/����
矴H��C�I/O��<1��>�ȕ"t�\/_�tB�1�x0F%S>Vb q��YaH�C��1��A��,�hL��G��o�jC�ɓG����a��!B	tiQ�ȻL�B�&tgr���'M�x!61h��B�u�C�I31�иE��T.����^�74�C��dg�p�%OC�|�>%"���*��C�'yJ���G�*N(��Wm�$~p�B䉥2��Ѓ���<�)Zqw4HB�ɣ �8�&�W6R}�:�O٣��C䉍�(@@�I�c�lY�M��B��@U=I�L�xb3��><B�IXŐكԃ�"B8�Uɕ痬(�B䉔�\�%.SI��G�A0v�zB䉣@�.=�P�w��2�J߯j2C�	ej`e`�KA;,Ű`�3�^�|h0C�I�Hu��R �8�)�s�܇�4�?Y��IZ��D�۽�urR'��!�!�$���UsËY�|<�E��~}!�dɹf}V�ڑ�U��.d�g	5{}!�䜶Q#v�(@����yS���p�!�D��A���[�7,��ue�4_�!�	=N4����o_�f ��D�ړ'�!�� t�1�/��>A�$�$�Z.x<e��"O�HC`��L$�'�C�b��S�"O�8[��n����#�F�%����P"Od=��E�6��`���q����"O������p�r�!Sʓ$�0��"O ��@�S\��az�'T<�&"O:!�-���YQX�c�KN"�yr�s�

���;�}�����!D�<3u�j)��s��
;��EǤ#D��Xu�)D<>Tp1�̔K�ųģ'D�(�7E݀A��iR�*;43��Y��'D���r"�=[�	HB�s�`�P('D��I@�
�M���De�b�yrK#D��a"BQ���g��0E�?D�0��&�1A�m`D��$�y�E�.QT����w��w� �y���]YB�(߃m���`����y­-(��K�g �bx�$�._��y"+-~��-
ц�D�l�AӶ�y�%�����JG�OF$���yOX�B4b�ʸI-�Q��ybL+x��Ap���1<�<� ���y��T5B�d[ץ�:30��0�G#�y2aőv���x��»'����w�Ȭ�y�-ѷ���!�Lvx�p�I��y����&tPRNZ|@\)b�C�2�yb�SX�,i�E�8bhp%2A	E�y2E;d�vQE�F�
��`��>�y�	�[Y^���ލ�j��C���y�m��Gx�\�VcG
?j������y�CU����H1�%X�̘�2&���y2NҊ{���ڱ,Tz��ԙb�E�y�&)Mp��`�s�F��0EG8�y�A��[� p��$��	7Ѩ�y��=w����Un���sAU��yr�6 �͢��ӝ@�}�P��y¤�sw�d��f�	<�<R�c���y2N֌M����׮۝8k<�W�ˆ�y��ȷ��U��Nϳ0��������y"%�7���A�)E�M�wş4�y��N�D��)�%�H���M��y�"�x$#��ޜ�A���y�C��t� `��U���h!�Iȸ�y��'B�y�wĞ�w��)�դO"�y2��
�s�hT q`e��*X��yB'��8�#��n`hب􀎒�y��Y)8r�ȃ��T/ݪ�Z��y�CI��p���
F�}�̘�'X�yL�-6(h9PD�{�TI22DL�y�	?}!��A���g���1��yRG�O�Rd!qL+af�y�LN
d,̘��H,l"`����-�ybi_0��@���ə��}x�&��yr��c�)R�n�5/ؔ���l�/�y�
��Q������>,˖9��o���y��V�&�4�3��� 2kd|���X��y�e�� ��=Ro�.Ez`�o��y�ⓠ_�n��g%X U�@4����y���5Xtp`���Z1q�#(�yji���t����8��-��yҬ��2���BW&�3��y�b,���y�vvtt�{ !��K�y2#\��ţU�k7Ve��O��y򅙘4= hI�L�!7ڢ!��+�y
� ��#ԍ�S���&�!=���"O.�1R���֍s��d&py��"O.�@cF��]�jQ��K0b�Y� "O��q�m�1$嘄��j
�B%�dз"OZ���-�\�`5 Y.1�Y�Q"O|�{"&B�j̍�/X5��"O�[�������N��i���Z�"OBȪ4�Z I�����̏X�B���"O�8�!�4�H `o7\��qt"O8� �F�+&xQإ�]�Mk0��B"O�,�QƎW ��K�K\����"O�a GZ@�1�bkP�s��u�s"O�G�һ{J� !WEQ?�>�I1"Of�j���;N�4#���Y�!�"O�kT�\wl)+BA��%o�P�U"O�Y�U�'xƼI@�O3T� "O$��%b�:` �@��Ң~`�i��"O�H��یZ(]PfP]���"O^`0����,W� 9qd�@�<���>x"- CѶ�r��y�<AC��=a+��K;c���;*u�<	�$Ą���Y �D2~ Z�;WlBm�<��H�Fs��CFD�O�N5�͒j�<�WJPLt@l���ZF�ES��\�<��ŋ1
� �Qd/�$�7�PC�<��Y(Y���m� �����H�<yv�"8WB݂aaվB��4�E�G�<�C*
R�vc2�	�A�-��g[�<y���6�I����TݐR�k�<Y���� %`OB���q&Fk�<	R�1�P䙶i�4h��=�/�Pybn"1�6��c��
?� ���Kc�<!������w�Ceh8����Rt�<��Y	a���D�#��)s�s�<�%gS�����L �8ϼ��`�o�<��&J3���&	4a'����_j�<acg�6��@"���0^r����Nk�<�3�[!�Pd��
�/h�2��vm�}�<���O���@g�/@��A1�L}�<!6*�707�PH�A�:���w�<Y�b�m�F�i��]�E\)b� �Z�<YC/�K:�����%@
u8f+O�<�3�Z�G�4(��?������N�<��*T5� ���E9#�����[N�<�4�­M�.�9��E5y��Ii��RL�<A֎�Po~�.GѤu���KR�<��I���1�u���I�ʝ��`�L�<!2�"erY��c�e:R�b�F�<qQ�]u\8�4P�\
��X��@�<��-!b5L����3\s�� �b�<a�C�D�T<��0|� ��2(Ja�<�d�FPz�y`��i����kZ^�<� �T�yzb!*��^C6�/�X�<�cE�/90�q��l��e�"C�[�<IK	�\��Dx��ȻG��Y���\V�<#��=M�dS�H�����k�y�<Q�$L��l����Եu�Lp�/^�<A��O�MH��2@^�1R�Y�<���6����k���|�Z%X�<iao�A����Eo+DRZT�#��y�<��h��'� ����'X�6Ѐ�"�s�<���O/�2Y���]9C�n%�*�k�<�t��&�JsA�/b("3�e�<yvL���E۳�_"U�L�q�IG�<� *l����$vd���aG�*=����"Oj�+#��+C�R��V�׸�{D"OP+�i�>'.�AEQӀ��5"O�q"��k`���l�|�G"OV��Ζ2C�����-�'¼S�"O0�i7�T2N|��Z3MߘC�V�F"O�8��M�:RpPrbX9\��(x�"Oޝ(�N�GQ\���KČF��r"Oh�CK���T�,
4��h2g"O�xWf1��Iv��u�X%�c"O,=1W�M��4rFK&�X�8f"OD�CD8� ǭƽ�� ��"O&�D�&mO���mW&w�R1(�"O��Ak�dH 	cK�d�4a�v"O<���X�o�E�`�	�>�fTq�"O
���B� ���G͎7r\��"Oj]�� M����GI>-]lt�"OI��@�3fU+���)�JI�"O����		�o��VC��l)Hw"O�a�,	|�c��	�u��Ź"O�EJ��x�*�[$���n���E"O�豦��< ����K�e>�˲"O��)���q��`�!�{  ��5"O<Q8�c_�@lkU�.1��aW"OhD�jn�`��K:N ��"O>5�#��>p,��;,�(ra"O�(E#��F�x��C���`3�ݺ�"O�h0D���&�@١���O��3"O2��C�B,x��7P����"O*њ�m_��"����՚%�81�"O΅yD��]
�f#��a�"O���)0w�و2�9g���3�"O����(��4��*UC�e�0� 5"O�i�p�EtG�:0�;",��&"O"��tbZ1VK�D�TBM���q"O�x��m.�5�r(D�8u0�"OJ��bQ8d��Q d��3R��E"O�}�Ӌ�R*rd1�0.�q�"OR�R6J^��P�܍��if"O^bw����"So �#��@�*O�(�6�ݪ1����鼍	.!��+l�@S3ɒ�S�FaEI]�-^!�D�Yd��"M�3I<A��(�	V!�T't�
0f�J�Z0T=*3�GX=!��A=i HlS�IJ�! D�З��&L!�QN��ۥ�����T�S*�Py� �
��\��A	&}�8Ё�I���y��R�|Lj����,uw��N�<�y�c�,e�$�^� �8�ג�y�;0����%oӯ"&�8��V��y"B_]�Q����:��%C]�y�Ƕ`Z�Y�*
�42%���A4�yX�r���Z�&� u��8qhK)�y��)D}/�q�������y2�ӣy)�ũR�`y�u��ߕ�y�嘥Hm�Õ�պDL��PхA*�y�.
^z�0AH��*�JQ����y2�	Nv�@ӢÚ5l|\�&j��y�m�&�JXz���8��P�F���ybeL�T
�"�Bb�����y���*+� � ?�Bᩔc��yCY�;�I��ؐP����/H��yR-�?0��-���2� �{�%��yr%ѶM�n1k�뉸R;��z���y
�  �
B��*>鶉X� *;�����"O؈*3�!b�ba��i�.Y��8��"O.��0-��F���r��Ѵ
�:��"O��)Ԥ�.`��ƅ]�)�ͣ�"O�i�g�ݦD�n�b$C�!A��|Q�"Of! lE$Oz�� ��Ϡ��B"OR<���E�b��s¢߸"ɖ0 a"O�����!��ۓ��3y���"O|���C5T�d� ����w"O�A#$�U��*%�V	F�<�*�"O�������Urަ��D"O �:�]8CV��lD�5��!�r"OY��B%d�
��T���Kg"O��s1���d/[:��TR"O6��������DP�L�DԂ�"OH�
�֞9��vDI1i�<�i�"O���3��/[��む$36�"OIy����u�=�Q��y�l�b&"O�� 7�ȁGT90���|��"@"OZmD����` ����'I�b�ۓ"O���Cb�Wk �I��k���S"O*�+��<^�p �H����a�"O����M�L.�fǆ���'"OJ�aEa�"p>�X�c�[�|��g"O�i�,τg74�)#P&��<1"O�}���ȱ��E7�(��]Qt"O�P�C�rQ��]�D�h��#"O\@J�O�;B(���� rJ\�P"O4h�a�Xu�9i�I�7���Q�"O\!ˑ��<(<t�)�	?2��U��"O ��cS�V��89�o�GC|
�"OV���:n|P��ޖ;�P�b�"Oh��s!��$�d�sI@)M*���yRh��j�<"ĠC���
�膧�yr���%��@
�ܵ�����y��7.�`H��N�g����Y��y2�W�Z�i+G*x�:���L��y��Tk�h��5O�$ph��	΍�yr��%w��a��_"p�B�r��9�y��	*4��j։4XE�F��y���S݈ɣ3nQ$���gd���yB/!|N��5dɤU���G ��yr�+��ie�ȉ"���c� ���y�mF�A;�ab�Y $0JA��y��I������*L�h�6���yr��M�$}�Ƙ�Smx5�5!"�y��W�k�J��F��9`��� ����y���<@�K�D�%�Mb����y�-�$'�� �0�H�K�(�yU�;�@��'�ס�*wL�5�y���17���c�=2�\B�. 
�y�ժqU��YvE��t���j�
[��y�΀�Rܡٵ�K0$�$	f��y2益^��P�dJJ�"mIB#�;�yRf��;�dͨc��G#��"�՗�yBoK�N��d��BJ�[�#'�yaA1{��mr4�F�&+н�Rʞ4�y2OS�rH����B/	�d��b���yHQ�xr��E�}���N�y�-�S]�U8J\?d���9d����y�@.
����ܡV�0!��oþ�yb��5(T<�J��\5;q�ǅ�y�+�m�p�3g����Ejq��4�yR��0��јD�5ur	��/^��y
� �<Ҷ��{��3n�v
���"OX��ŅH�P��Ƀ�/�
�6��"O1��%��4�R=��o֠j�4=1�"Ol��C�,bPiW��|L�AV"Op���9"rӴ��7i���e�	���g��r"�V�'���^?9��	;|�]�c�[0N	�@Zj�����?��xhN� d�R�%�}��\WN��Du>�rc-�E����wg£~|�hum3�B���2b"�v%�:-
|`!��ީ�McƧ�P���Y�Ʒc�*����Lb�'a1;���?QI~��4���j'��B��s����O�����'��'���'�^� Wg� �h���^2z�p�
�y6���'��&�I�26Z�ѐφPHD�Ɋ�~r�:c546��OL���|r�)�?Y���M[ ̴km (���[�m�08�ʌeF�:Ն��{�t��7 d����Ao�.���)b��EP�8���5I�4q�Hh1wi�&�k�P��ٚ�H�������>�5�~��3,l{���	.��Q�1��o�l�"�d�O�p��J��i���K���#����5ď�
�.,��'�2\�LD{*� !0NR���TW�$��剎�Ms�i;��]0$�L��Ĥ,b�l�!�S����?�$�W�5�,@`���?���?��U?�m�[A���ÅDE��-s���5�`�fb	�`R�9�ϔ*�M�5����Q�'���*v��}��e�\�|���d��X�>=h�|) ғ`C���	L�@��y�<�$��+�:̚��H"UV����� �M��)���'�
����D�Op�>)f���
1<0���H�%;N,��Iw�'>�1xDm'l���o[��"0X�G̦-�	M�I5��I�<�� c1�J�,G0�8¶.B�~1���#�?��?����0���?i�^���p�xǄ�	��sμYb�uE���7#��n��d����B#?1�*A7.��Ē�!�����:PN�[�8M��ǄJ�������4�$���,I���X���O�6퇂`R��geM�_p�(d��"v�~N<i��?I�*���:F�D"4΀-Sa��39D����II����Ll��:E��.�.؉ ���Y��DHঁ��4����Y��$nZ����E�DG�ty�Mk4$4������jt�����O|���O|� �!�):Yx��%�G,]����
��!��e��zq�R"Y�d�q&���HO���s��6��=���/Z��(1=��Z�,� I(�	��m�֍[�$�/�HO~-Z��'�rbg�X��~r��\�15�\�T
�XG�ju�~R�4�����G�T��^�%Վ�P��'m|9��I��ݴ�M�!�:�aK�nE�}8��_���6mK2JR���'�b�'9����l��'6GH�p�6��߾
�bTa�$
s��D�"�Q�ʏl:j��r`�����_>A���ہo�W��5jf�9V8����������V��ST��i�F���$���
��\c���&E�Lo|,)X6r��8�4B�\�	񟈨ڴ�?����i�>�2�CZ�t�,�Ё	�C�p\��'�"�'!�m�!�V�_��s�&��B�lB�'��'�z7mDF질b^wfpH�A�m�PԒ�#l�`�ff)�D;lO�(�  �   6   Ĵ���	��Z�Zvi��:+���3��H�ݴ���qe"���@"<A�iB���gC`�����Q�R�y��U�6��7�i�X�����f�TYؔ�.(�r��j�j�ቄ@2�Г�i��̩�+�>8Y�A�Ϭ\?�Y�.O����I_>7r�P�_��Rs.H=_��8�>�@��/H^.Mr��S��
�r㠞�?B�r��r�$�	�< �"{������
���[�$z���SF��F0��&�� �x3D��$oy�M��Li���R��8���4@x�'��Fx��Ba�I9Н�s�a�X�SE&,T��	69x�\��ቱ�PH���>��8[��P�<����ď��O��	�O��ҀK\lQ,��	x�N�i1�>��-tB�� ����^-:�0��I���!�a|���������O�H-�'!y� bf�T��jԋ�st�O����d����� a2�l���S.e�P�Е�	�ai�	9NF�$!7���(]n����@}ƴX��`��G/"�*��Z$�O�@s��;FT�kS����p��J�V�
!�<y��!ϬOF	�e���Y�I�(�n<b��OR�����Z��ē��D�,Nb�(jB�K��P��J�U��x��J�G�\Iml�D�9jE����'X ��j�-߃x�	j0��n�Q,O��p�O�{8�'@ \�gC����axr��S�P�k���U��C�P��s!C~�<CI>�'yQ�x B����W*W�~�.��"E-D�蓇�   ��L�;�) D�(�e���8Z�A��	�5r�Y�b��>і�6@�����;I�U��aʤ	�H��`��ra}�Ɋ���)� l�����?��j���#�.�z�"Oz0�seۅ6#�T�!L^�*�:=R$���z1�wm˥v�>	�$��._)�L�f�W
E���<D�th5�V�p�UұBҗ]����u�Z�h�Z�O]�4\�u��?Zﺓ�4]%��2�z��x�收#����'�O`(���C���ݹ�� �d�H�dD�-N�"[��߿�J���Ɣل�	?4Ƹ�Za�<n���n�T5�3�	�R#�Q�g�L����P� � >�p���D\1�	�`�r�CM��y"�Q6u�hu��9=
�X�ǃSy"Eճ����`�?O�k��V=r�D�?�X�#J�+V� ����$q�p�#D���S�
n&���0�G�7i�	U+N?|Uޡ�    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  ��   �  ?  �  �  �)  5  k@  �K  �V  4b  sm  �x  ��  g�  
�  ��  �  e�  ��  �  +�  }�  �  }�  ��  S�  ��  .�  ��  ��  5�  y   � l 
 �$ �- &4 �= �E zL �R Y �]  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+���6+\�s
�<4�d5h��'�B�'���'	�'/�'�B�'��(#`/�P`b2-��
�v1��'�'�2�'���'�R�'���'�APΚ<�z-�,�Ŧ�@��'�"�'��'���'�r�'�"�'�d=Q�n۶P�r�B�oM� ��+��'��'�r�'	r�'���'�B�'�ҩ�Ƃ��K��Y�RmɂX>����'S��'���'�b�'�2�'B�']t(�t��7���A�k����'(b�'���'���'b�'a��'&:)'Ƈ�S�d��R�k�ܵ�c�']��'U"�'a��'e��'���'S����l�/U$�L�*ĶI�.����'���'���'9"�'2r�'�B�'��l��Ѡ{h�1� �"PN�e)��'nR�'���'(��'�B�'DR�'`\|ؕg�
Ɗ}���sʎ�{�'f��'j��'�2�'�r�'���'hT�	���,8������=�q7�'���'`��'�r�'���'��'� xRP�ڜX0x �S8�D���'
�'���'J��'
b�'2r�'.i�B�{����Y0�ㆀ`8��'���'��'��'ZR6�O��$��x.��2��/_��0��ؼw+���'��R�b>�p��Fɉ�ʊx��j� ��%a��U,h]a�O"l�D��|��?�D�٦����ǯ�/V��4(�@�*�?��^�J�4���e>�#�����y�F��&�"6|�u@�?��b��Iiy"�S�JQB}�sa�!b�-�T6J� �+޴����<!����r��N�a��� BG�w��Mh���}���O��ID}���͈�2�F6Ob�Sel�Fľ$�p�3zZ-�6O~�	��?9��5��|��_�6L1� g��5�֩�TZ�,͓���:�$ Ц��1�	8�J����8xJ�i`��фJ�\��?�EY�����<���d�Y��m%�C&kͅi? ��'b�,Ú<�~�����ڟ �%�'�n8*1��<G*�}P�l�
^]B�:[���'\��9O@m�Uj
2z���B�/L�>��"3O(`nZ�!^�ڛV�4���r���^j�����V����8On�D�O���9W��6� ?)�O���镇=B��
�F@#NYE�J��zL�P�K>�.O��O����Ol���O��CC@�O��gI1
5���d�<	��i��<�q�'��'M��y����{a�8Ѯ�:5��<A�3M�ꓶ?�����S�'ؠZ�	?\�zM�f&	D�Ɂ�K!�d��'�4��+
֟�*��|�[�(�֍��C���XR�G�J�n�E�H��`�Iڟ���̟�uy�x�(�@��O*�IkÆR�09E�W�"�
���OlilW���ߟЖ'�>8��ܐ�l8� VT{ԍP_K�&���X1�ѽ�dd�S���i�g�ZC�Dzp�Y(Ŕ0n�`�������ҟ���ş��J��T�4����^�n�
3�ֱ�?A���?ɔ�i��@3�Ojbca�6�O�5#b'�;sR���ˢY��Eل���O�yw�1�4��$Z39v�lSV��\��8q��R�
�!�iM��?�Uk#�ĭ<����?���?��υ"�����b�����8�?!�����9w`ȟ@�	˟T�O6�-�w��#�yi�O�G9Ld��O
��'�b�'�ɧ�)@5j��c�R�g�X8@����)�D���Y8*捬<ͧ0�h�䙷��1�(mXP�Y�?o�L���ɠG�:����?a��?��S�'��D�-R0fG(7��};���/��X�V&śJt��I��l��4��'����?)�h��8�@ȺҌ�Fx1��/ʆ�?��D�ش�������l��l1�.OV��O3�2 F�z�ْ�;O�ʓ�?	��?���?������G�~���6#XNj83�)�'M���nڠC�d��'������;'3<���ƙf�>����.���	ɟ�%�b>��Q��ҦI��*BQngN��'��(`LĂS?O��D��;�?��$�d�<ͧ�?�&��Q@�
`閲|��"T��?y���?����$�Ԧ]�`o��@�I����`N�d�3����S�J|`|��?�cP�`��ɟ$������uf0�Sa���8MӇ�&?�u�ȤU>���O�Ķ\?�����?Y���@�88c�Һa�txj��?����?���?�����O��bp����x��� X�'d�pf�ON�m-B�I̟d�4���y�j��&7P�ւ݀2R�4�`▬�yr�'m�'��ˢ�iT�I)�(Ȱe۟f�����N�j���'�x��(�C?�D�<����?i���?���y�Νmq�ZfJ�^��gả��ɦ�Am�xy�'��}R��>/��jSގV?��wk�g}��'p2�|���V��T8��!M}z�ӑ��
GeP1˔�i��	�.�I��Ov�O�ʓW�%��aD�Q�R�`u%�!||���?q��?��|�)OHl��[e<���*�LU��/K=i4B
�z�8�ɏ�M���	�>i��?��N@ �M��GR@�	'%�/P�H�ɛ�M��O�D�BR������ �P(�R�7D�-����5A5�:12O(���O8�D�O���O��?�(��
m@1"��G�>F
@��̟����hhٴ0a��ϧ�?QQ�i�'�zeD*iA�Y�$�/^�Iw�|��'��O��d@%�i2��A�^u�1(P�5�����ND�X=N��f_����4�D�<�'�?Q���?���)~�,e3�̂�s�H����9�?)�����٩ ��@�	����OE,��f�:%0���`�E ~�d(��O,y�'�R�'`ɧ�I��b�1!�3��Z��3:�v0)Kn��B�i*�i>ᑳ�O��O��I�Ȇ!f�,`'ǝN�f���m�O�d�O����O1��ʓ!�֎�� PZ���G�]�����V���@�'�"gq��PS�OB��dlH�����
x�ycD��d�����OTA��Ӿ�Ӻ[�/7�*cD�<�@�>��% `� "F$鑭
�<�+O����O��d�O��d�O�ʧV�A���qB��!�M�l�`��b�i2�$x`�':B�'��y�z��n�"�d��.̢@0I���J�`]��$�OƒO1��h!�Hhӈ�_S�R�b�\u�s�T�1'n�	!5s���%�'}J$���'B�'�@�wΖ�*P��3"Q�F����'�r�'_�2ߴg�T���?���62��#c�Ր1ȸA�EϞUL �{�Ҡ�>!���?N>��	1!�f!����_^ K��u~rG9�,a���O�.q�	�gr
�f0�%L�$0�@��Efɸ���'�"�'M��S�������9�M!�2X_>�RQ���۴	�F�Q.OLn�N�Ӽ#�Θ����e�Bx`�����<��?Q�*P*��۴���6�yS�'f��c�6����dl�1M.�P� ޝ����4�X���O���O���V5%�� �nE�M�Bp�ბ�˓69���#�	П����IX�d:�lŏ~�0��p+K=k���ɟt�	G�)�S����p��+| <@[FJ�-X�N����-�h�Z����S��O��pM>�+O�T`�(�'#���x�BQ+y��<W-�O����O8�D�O�<�ֿi�h���'z�q���c�f��֖9�B����'1�6�3�ɥ����O�ʓ}�X`��#����ї)t���cC�M+�O�` .޷����!���שּׂ��)�
U^tx�vEϿqv](a<O��$�O`��O8�d�O��?�c	�E���ֆ+К��L������ҟX9�4$Nȍ�O�~7�+�$�(=iH=��I_����&L϶�v�O��D�O��^��6�1?�;iHx�Bƙ�D5Ba��'2u�h� �(�?T=��<I��?9���?	F�R~�m	�c�__t��S&"�?�����dFͦ�ç.L���	�ĕO�1�w���i�Q���Ǳb�<���Oze�'r���?�1s�A�zD��%��#�a3Q����Gqȭ���K���!'�|BG��y�<��P��o���C�6S�'BR�' ��^����4C-qJ4��ܰ2,�>L�T��+['�?Q�~��D�p}b�'��mq�0"t�!j�*8�����'�r��
%�������CL����~Jh̀4�X09�ǘ����jA�<a+OX�D�O��D�O�D�O��'!x�Q�Ɏ g1���⍑5K��!��i� }��'Qr�'@�OR�Li��A�P�	�bN���򆪂(PcZ���O�O1�P�PEia����*2�;p�!R�̈Z�]���	��D2��'�J$�L�'��'t���1��Z��dеa��[�Lig�'���'(�S���4Z��Z���?��/����C�[2d��*2K��[� �Ҋa�>���?iJ>u(��s�и����+>:$P��F~RÒWh>IP�K���Oe<Y�ɹ �"�0 �N�� B�@��Ӈ�����'P��'�S韐:c��*�8��G���ykꟄ(�4[hJl�.O�m�J�Ӽ��`��#��1�YS� ��nC�<9���?����,��ش��d�#�,����0N@�R��B!7��U�O"1Ȑ1r+4�į<�'�?)��?���?	7�!�(8 D%W�"����N(��D��%����ٟ���ɟ&?����Nz���	ٕ|�l��=b9Rp�O.��.�)��?�� �Ua��y$@*Lū0�݋A`H
X$I�'�����oF��T���|�_��
���L@x'�>QN�}�"G��t�	��$����sy�H~�K1��O�� ����&i
�:!�� ��\W2O|l�c��P�I�����ߟ�Ѐ�1A��ٵ_4Jf2T(&O���o�R~B��1<&60��Rܧ���r�[;R����ᗼXL�w͝�<)��?���?����?���cJ�7�h�!uhR1:j�v�
{2��'�b�|�^aSs�<	!�i|�'����Pm��g:\���ڳTb&����|��'�O"�蹕�i���-68p!у�!*Na��U�g�,���8�TV�	Ry�O�R�'^B+S22`n�	����G��1��Q�b�'��	��M��Q�?��?)��hJwf?R� t���Lt�E�����O���O.�O�S�\d�h��D4ny��z�FL�?::��E#��S�T��6�/?�'4����9��'vة��&q�p3hӏ-kzDp�'���'�b���O�剐�M��, !BHPUb�|���B�!e\$���?��iB�O�y�'�"8"%��������� a�R4r��'�P���i9�	od���O4�g�? �\
�.��C�+@���(�Ti�3Op��?���?y���?����ɓ!r	��8g���Q��+`�~��Yo����I�� ��f��r���w{��!��#<���̐"2�����'��O1�����bӞ�ɦ0xP�Y7':&^�M�lB0^Ҭ�ɛuEs��'�& &���'���'-�0�BD��\w�=`�&]5͘�+u�'Q��'}r]�\�ڴv�D4����?��2)\��ʸ��m�6#A>-�|<:��o�>����?�N>�����/R!�	� ^��L[V+Mf~R�4�B�Ǿi������'��C�,5�n�T�B��*�h�n~�'�2�'�b�Ο<j��\��A�3��L���Cd������40��qP-OR0m�Y�Ӽe��,�d�8�,�*S�R�cGA�<����?�|�HY�4��T�<��y�';c�LRsHUH>�''܍%$ �ȕ�)��<�'�?����?!��?�aK�w*ƀj�hG�������d���MEBM�X����0$?U��=�L�B��.]�`mzW+ɜJ�DY�O��d�O�O1�LpI��ư\�v��&�K�b�PF���<6��\yk�"
��U������E�t�y��R�4�KQ)I�`���OR���O �4�2�<���OT�C��=r��M���ٗG��0�f�nm���$㟰�O����O��$�*'��-�䌒�j�^�')S�E�fT�T|Ӯ�L�~�J�>�>Q��5��MY0��	�t�3֭�>^`�ԟ�������I����t�'W��"���v!b��*:��R��?A�֛F��6P��ɨ�M+H>ID皫ь=��/*��f/C����?���|�ƀA��M+�O뮑+*o��G�pz��6eԘ �!�F�Od$@M>*OR���O ���O,aă�@?��a�k�&�`V��Of���<i��i��l �'���'O��6�h1���a��#j?�IZ�O���'���'Dɧ���o�$x�0���N� i)!lN�mj�X�+��c�8����擸��)_`��A&\��n��P��e�e�H��� �	��d�Iܟ��)�[y�Gz�@��޾sҾ*1��X��ɠ����{�˓{i�V�$
Z}��'��U�w���.>��Ȗb�3I���a�'C��/W����a!���x0�D�~�bE��>*x�3�a˘X~*2�<�+O`�d�O��D�O����O��'��(Pjw�R\�V	��H¶l"�i�2]���'���'
�O�rcx��NYdjd���ĕK.�pf� E���D&�)��L��m��<	�H�k��H��sN�J���<�O��4���Z!����$�O����3�ސcF�ӱf���� Gޜ�2�$�O��O�˓����_*Ql�ğB�h�dֶ|�CP�9����6#X`��I��	П|�?�`R�CA~X
�>^�;�J�n~"*�%5��p���3Q�O��d��2Q_ۛxU����2Ú�ipI�J���'"��'���s���e���
m�<hèJ"�Rq@����D)��r��J՟���M���w����d��AZWbR��5��n�8�Ipy"�Ӵ2��������/��)��DH�V�nu��ې���� �D�nu'��'���'d��'��'����D��::5�ւ�-&�,��X�,i޴d�<5����?1�����<��C _ ��ʠlH0.^�Y@���x<�I����z�)��48�1u�ܱQ���%'�\�0,�S��=�'�s& ��g�|2V�pa'��?$A��U�=�<��sAٟ�����t�	���py�ee�`�S2��OH�`f+��<Y�r�ߛs�>(�=O8ll�f�]���|�	�|B��C�@�ܩ�/�:E�p[��/R-�|n�D~�m��k��F���w1%�2��v�N5`���hZȰ�'B��'�2�'-��'���L��n� s��Y�An�� ��O �d�O��l�?s[�ѕ'y�6m:���K���U\�%J�	���"�h�O���O�)ԍ�5޴��D��c��IЅ� �R��pI�	��"�X�i܄�?y��+�D�<ͧ�?9���?ia��M��=�c�$,�Ѕ��
��?�$���$J�Iє��?���ԟH���?���H
>d��$��*!��%��Go���I���$�Ov�OR�'�?�ig�-8���#9��īf�Q0�
�� ߙI�2Y�)O�����?�di.��<]���bG=W�>=ZR��W��$�OP��O@��	�<11�i�5����p"�0M�i����(�(��'|�6-9��6��D�O��2 ��	�h��g!�=���B�O0���)�6M>?�$�ǻ>��>�Y�S�y�aD�K�����n�ȕ'#2�';r�'b�'���I��؈���,!�Ej�@˿m��i�4+�ذ-O��D;���O�hoz޵K��0h���2�W�XT�U�I㟈��j�)��d�N�o��<1���
D(+Ő# o�@�_�<�@�J�:P�I`�I\y�'~2ǟi�,,���R�B�\�[�E�f��'.r�'I�I'�M�f��?Q��?�a�<,N��g� �@��n���'����?����V*�2�S�3{80��EQ3	*���'e�0aT/N%T���,Y��'�Q�Ƈʴp���i$*L�/0E���'P��'�r�'0�>i�	
;�d���H%I[>��M��:���%�M��ꇧ�?��G���4��%K`	�N������21&�)Q8OP�D�<I����M{�Oh,�b"�b`� $\�`�x���8,�.�Z���i+�d�<����?9���?���?��Pxaɪ@�/W2��R$�7��d
ɦ e*T�$�	��L$?-�	�m��P�NL���p�S�^ӊ�ЮOp���O
�O1�v���c�3-p��A�.��0���)�kb�<����\P�S+��%�x�ky�-N|��Y0@�W4\ �A�b�'��'m���S��@ߴkL�x����Tx����82.��i B�m͓}�����o}��'~��'쀐Xf�=Yr~�#$å+�0�J��MZ�������bԸ 'Q>��%Y�2��&%ʫ6�<�9WhI�z���P�	ݟ�����t�In��)M�-jV睽jizSπ� �N��*O�DD����<
E�i)�')&�놉�,��E��rʔ<X��|B�'��O=�Dk��i��	�I�������&h��K���|��b��ֈN�d7�D�<���?����?��� �M�BA��TD)��S&�?����ꦡ����T�����O��y�6ɓ�r/TMÂ��X��Ya�O��'C���?�Rv�άA}Z���5G,=�d+e�0��]+�0���ԀD��pS�|��ȫg��� �z���ѳę1{��'B�'t���X��ش,Ԥ)��[�3=X�2Úg�.H��j���D�Ȧ�?�2R���I)K�ft�S�Ē0�6���@JՅP�d�	�?@dl�R~��O�_����@�ɒ�jؕLׂ=�6A���-\�Ķ<����?A���?!���?1(�0ոǮ̰���3V)Ai�zAq��[٦�Zb%Uyb�'��6Dmz�k���(m�����
1rr���a	�����}�)�.� mn��<iI�R�"��0LQ��Jfn��<)5�E�d���	r��ry�O���T���02��%g�����,��2�'���'��I��M���3�?Y���?��J�h�H8�/R.F@�a V р��'bꓨ?9���Y�����ʜWK��Z�ݑ ^|)�'���au��>�К�������"�'�ځAF[1��Ʌׁ�������I˟d�	ퟤF���'�6q�����4�EMGpu�(XA�'J�7-�1F������4�]���X�HHkW��Jˤ��t1O����Ob��$7&?�u��2c"6�)M
\H"5��"�V��\�W��`�M>���?ͧ�?����?���?9�b�#I�����cN<���Ŧ�?���`�V�#6�S�?������?q�i���O0 A��A�7�2G��<6=:\���O���O��������u�R}��8��kԊ}J4��L���"�%
*B�Bɺ�@�(��KN�恲��T� �O�˓u,]�F Ke+���Ak�m������?���?��|R/O��o��L$����#Q����GM��N� 颡β$�t��3�M#���>	�����7iX)�o�8sD���Ld�R��}���|^9�-����J~b�����`r@�2r�|q�!�0j]:mϓ�?����?���?����Os0(˔k��?`ȩA"O�'}�H�'���'�d7�� h��c�F�|��R*�i�ŠƑG��|j¨��5��'9���Df]�rO�f��0����L>bA�t-	���1E�ӵ>`��ɴ�'�B%$�����4�'�2�'�`i�&�9)<����&E�0��')P�`��4J���i���?����򩃄$M><���'xj�`�v	
.5�I(���O���m���Y��V�k�*����"m 4��F)O�8-6����+��4������J���O��3�3X�b��T�xp���bh�O���O��$�O1�4�����8�:����3�D�"c[�?�v1�'bKj�`�@��O���v�l��C+�0���˔��>�����ɛ�4���F�"���(�'NI�˓P��4Ҷ�υmy��"ŮMd��(ϓ���O��D�O���Op�d�|zAH�k2�����"%S"�;�-	�tA�vnשu>�	۟�&?!�I0�M�;5|��\�]CU"O�;��A��?�M>�|"���M��')�\�Ԣ�*%�|<�c(����h�',�R�C?�O>�/O�	�O��Pè�#!~,�v�F��L�����OH�D�O��$�<�i�`�22W���I�ZF�H�#	�Rft+e+��8I�1�? W�H�	_�"�ܘ���\�!�b�8QL���R��'B(��`zȱ Ð���_럤 S�'N6a���%~�H$@!��\�n\�3�'��'���'U�>5�	�e���&�A-u�(��Ȓ"m����I��M��\�?A�ʛ&�4�p�B���,�0��G�i�6O �Ŀ<�U�Mk�O���&��B��>I��4�b!ڸqL����ڼN�̒O�ʓ�?	��?���?���~G.�+��Y=W��`�MG6z��-O��nڑt����蟤�Ik��4����V1�Cu@	�P&�xZQG������O`��3���X���m�3a_@�,�GN��AY�X��u�̖'Ӕ���|?�O>I+OX��c"�
@Q^,@SG؂]�^0"��O���O��O�<a��i`l�y��'��u�a�-����)U k�c7�'��71�I���$�O��4�T�B�Ԋz��9�
��֩�����7m,?Q�3_���D��ߩS�`� ƀ�����0�Q0�{��I�x��Ο��I����%T�,0b� �LŖ��(��6�?���?1R�ie�Y�Z�J޴��GL�a�FLm-ҙ)f�A9���RL>)��?�'y	L��ܴ���J� ����	�]U��S��>XX�!����?�UE.�Ĭ<ͧ�?y���?�G>X T�cE�_�v���!�H��?����d��E8(��4�I��ܔO� �P-��5��CFO��N�)�O&��'�"�'�ɧ�IA<<�2H�,Ы\ :�Pu�H�B�c2K
$}���n0?�'/���$W��VxF%��o޲��[�ʆC������?I���?��Ş��Dʦ�;�M�.d��$��&��r�>uS�eX�v�����,"�4��'-�듴?D΄S�Iz�����J���k��?q�>t�C�4���Ճg��$:��4c�.��󢉞I���+�	�y�Z� �I����	����IǟėO�Ll��-�{�\�W��J���n��5�r�L��D�O��i����$�OD�4���".ר]V����B�lt�}8��O2�O��4�����O��K��w���	�G�T�kCO�s�.���'8���ɾ6�+g�'y�$��'��'FN�Å,#M|�7�\ `;�AA�'�r�'��R�Њ޴G������?���@CA��G��J���;C��1C�j���>����?yK>I@m�Pc�i��5:�l���
�y~�Dk�<Y�����O�>I�	�)
�h���̓�-d9��R0
���'�r�'<��� �v/��"��ak�+4�,���G������4a�iY-O\]oN�Ӽ�� �>�0��2���T�����<�����䛦p��7m<?逎i�<I�S}�J�d!�m�<���.˨|y\k�|�^����ӟx��ퟀ��������/3wL�	�K�t�ÅKyB#vӐ}¶��OT�d�O撟�$޳&`��a�KrY\I� C��8�'���'�ɧ�OXX ���n>JK�݃bFm���b\��"�Oƌz%�N%�?�E�'�Į<9&J�/{���RƲYQz�ó�A#�?a���?����?�'��DZ���C��ܫ�$�x��)Aʡd�h�S��m���ߴ��'��듃?9���?��O:6@N麄�EK	E�U�4��!�M��O)�U��?�R����w_�!a�HO��� ��/G�x7��	�'���'���'G2�'��RT�ǟ�t���@�h�R�I�O����O�0l"�<��'�p6�)��4���b�V��K�m��@�O\�d�O�)[�7�)?I!Ĉ*`5BC�3)ֈ@IA"_qbpF���L%�<���T�'�2�'v���m��?������6�� �'�'�"R�T��41��yK��?�����IZ!W[>�[�IH�`�� a@h^*E��	9��d�O$��'X����f�ҋZ�P�	L�F(u�J,r�H��K3��4��i`�-�>�OX�e�ZE�x�#�H/y�)���O����O��$�O1���u���������D�{)0iX��iѤ� p]��ܴ��'%0��?y���:9��f(A��FIQh��?��-m6`q۴���O�q'�j�����B���T��`�\�1�n�U��ly��'V�'�"�'IT>��D��X�N,R*D7v�� SEٛ�M�H���?���?I~���Qe��w<z"���	����J_03G� ���'��O1���#b�R�	�Z�,�$�µP\,	dJ�%��IJ�*x�Q�'���$�t�'"��'���B����}j�|ہ�S�X���V�'u"�'R[�����{�tT�I�x�Ɏ4�|���b�:	ADXb�H�N����?9�Y�D���4$���� �V�Ȕ2Q�O�.= �
,?!eb<���ڴ��O6z\��?�b��M����&���7ٚ�%�?���?���?ً���O$�nʵ�i �پJ�e����O"n� i�%�I���(ش���yG��+0�	 ��@;r�bC��E��y�'��'��0`¶iN�i�mB����?��"�S� �zu@�+n�L ����'����4������۟��	cO(hPʄ53��I��F 5�:��'�l6M�Z7
�D�O"��:��O��+���lڔ`jLC�<�	qK�>������O��2��Ժc��|A+S�"�6��0���<"H��[�`�ԉ�&_/��|�Ify��ߔ7�*J�%�j�r ��(���'�"�'!�O��	��M��n�?ٵ�U,f� Q;��3y�.�4��?	ýi��O�u�'�"�'�����yꁋؑ[Cz�wgII�*��q�i$���%w$���S��)p1��yI����핃j��Qrbc���	�,�	�<�I͟��z�hʇW���A��A%W���E偉��d�O�Aoڜ7kN�럸X�4��/��Ux�H�;j*��v���B�61�<������oOX6-%?�b�Y�L�2�#UZ�>�(d�ٞ���s�n�OX��O>a(O����OD���O\D�w�cB��`רcn�͒ՠ�O
�d�<95�i���e�'
r�'��*"�1�E�L�8��Ee�^���1���� �	q�)�14 ��)�p ��>/$��6��s�A�#ʈ �����g�П��Ǘ|B��9��x��,S>�8yu"���'���'5���\���ڴ.A�h�4�I�8�2�c�&�'9@�+������ڦ��?	�V���	� �M&�R97�� �U�M���I�����B����u��R<6���UVy��2Dt�"fi�4��)�чĀ�yT����ԟ(��۟��㟤�OS��AB������e�w�A�R�a��٘���O��D�O��?E�������\7��P�I��U/Pa8� �;�?q���ŞZ,}�ߴ�y
�  ���	��E���Q#)*��(B=O���FHI��? �3��<����?��n��O�����L�0�p���?����?����_��aG��(�	˟@�3Ł�+F��A������G��u��d�������	_�-{�F�j2�`9 b�>7���dj�!w��#Rn��|Rga�O�����
���IJ�No����Q�Ҩ����?���?A��h�P�d��� s��3	9|�Csg٠�D�-�g�nyү`���ݼ�\}�Ջ##��Is�@ T���ן0�'�4u�5�i��I�4�
,Ru�O�\Aᆤ�% t@���Ì�K�F���YF��Xy��'���'U2�'.R.(kkj��G��,�h��"�e��I�M�EÏ��?���?����
%޾�X�*[n������� �>������O� �����aτ)x��j�p���LѤ(����vX�D���1D��K�s�	qyb�O5 L��@��W�&�2�����';b�'��O�	��M#�d���?����@jXʐ�3,G��('̂��?��i�O8 �'�R�'5Ҍ:}����5��dŬd:Y�m跈9�M{�O�@��AX��(���n�q$����Z�1�҆S:���O����O~�D�O���8�� c֑���ڽ��K0" >6���	���ɨ�MC����$�ɦ�&�ܐ$��'r��'o��U�� �O��p�i>q�E�ئ)�'6$��#n��K�b�z%끾s�B٪���"�Y�I�W��'��i>	�I�����ٜ�*�H�7�P���ˆ'�
��I럸�'ظ6�xOR��OD���|�5/����5�'f%B=QU�A~R�>Q��?YH>�O��R#�2�(� C"!&��hgA��-�L�C���>l�i>9C�'4��$��Z�.0a�������m(E�l��ԟ��	��b>ٕ'�7-p@><���Cg�p�.�1`��Q!d�O���H��!�?�N}��'I���ᩚ W�ܐl�i�Ph��\�L��L �-�'���r%�M�?m��_���C&��� f�Q9l��"�x�l�'�'r2�'�'H��5f��y4�ޤ1b:��G�o�4D��4H�Ѓ���?������?����y'��|IhT�G=x!�Q�X���'mɧ�O��q1�i���	0*�i���E1b+4�.�󄝦_�@K�'Y�'!�i>��ɐ
c���f�0'�������#!�t��ʟ���<�'m6�\taV���O���`�>S.�/b ��LE<"��0ªO��$>���.M"�c/��t���>C��-*�Ћ�|��3L~��+�O��{��IHu�+�<5��!��EW�D(��?���?)��h���*hR����־'��)��]!>���AݦqhCʄ��I��M��w�Q�
�=�d�L�|ș'l�'GR��*1қ6��Y/��_ ��DI'E�PGi��ey$$�ꔸpM�p&� �����'/R�'��'�|�#�m];&|"�p��R�a�޼0Y��ڴ#��	���?�����<
_�Q��5C'" S��73��	ʟ�?�|:�N��a
!u)��	1���EÐX��YS�`���D�C|1+�[J�Ov�d;��7�Z�c�I1g̅(v
i��	(�M�ц�6�?i�Ҕ
tB�OQ�&� �+����?���i*�O,(�'�R��y���BBTl�D���^U+c�H�V����i����A�"�27�O�>�$?��=�*ae�}pܱ8#f�$I2�i��<S���J��C�[�o����qe��0����4{�4j#���OY�6�9���		��(�B�:؞Բ�ĀK,�O^���O�Z)K��6-8?�;$�������}�b
�d $�W@	��?9��7��<��nF'd*i ���bX��@�>�O��m�7���	ΟT��H���AH���!�U.��B�ڡ���j}B�'m�|ʟ�С����'P<!e)J6hO�,�G�D17��W�2��|�0%�OH=�J>YK]�B���H���|���PC�GE<i�i"�Q�2lR!40�Ȼ���:�0�H'
]/�"�'"�6�0�	!��D�O�kf��+f�)��(UB��pT-�O���
� ��7�5?��ǂh�b��GyB��-�(42r��F���R��L��y^�p��	 t�����	ʨ�
u�(�&+�D�ݴT�dE1���?�����O<�6=��x3e�h�(�h�%z�\ո���OF��"��i�.D�7-~�<��M�2Tp*)�`%�4�X���~�(C�҆R��5�ģ<q-O��#�a���`R'
Z$�����'M�7ʠa�����O���M�:%� �K��(%�
��r��⟸[�Oz���O,�O��z!/;�}����sTr���4���%��D$�i��$��$�����`�.I����S.o>�`X�f3D� �6ə'����`ғVm����B\��ش{DHZ���?1c�i!�O�N�m�@����L:z�
Q�0��-���O����O�xH&Jwӊ�Ӻ2dP���ƍ��V�r�&S�2�4����
�z�O>���ON�[S�ʫfQTLJ5o'���	a���޴%_�����?����OP*����[�'�(q�Gp����f��>9���?yL>�|ZR(Ob�? z�xT��V�pȁ��ʶm®1�Y�B̨˓*�	3� �O1�L>.O�*WHD� )��s�*D�	s"�'^F6�X�3����2*����νt�̱S����2���$�٦��?9dV������]+1�\�S!��*Z�*��E0sܘ)%�@٦!�'��1qӁ��?}�&����wf���R/EGҘ`fbKB�BA�'~R�'=�'}��'\�Xx��=!��)f�>SORd+��O`���O��nZ�r����쟨�۴���,�CB�əܖ٩��l��<����Ŏ;�6�-?Ɂ�=#6�n��OV<�3�A��^�(��O���K>1)O����O8�$�O,욦��O��@�t�V/X,T���O���<AR�i�d8Z �'u��'�Ө:�ٛч�pW��1.�9�D�n�������)�E�ŉFx��Z���,�h���K��\��EEU��Mk�O�U��~��|��B;�J�{�D�>�F�6�L;�2�'P�'2��D[��:ڴ+&�ԓZ �*��^ r��1��M�bЋ���?i5�i �O��'�S T��4�'���Z%�4f�9{a2�'���{u�i���(<��5r�����TԜAٔ����l�[�ߓi���<���?����?����?!.� d*S�ĜM�Z�/�)v�P�[��H�Q@�O�՟���ȟ,�r��yG���r����G��ww\CF�ΰC�R��)�//��7�s��j#댇0�ư�Tg��)X@t�k�|i̹Ipb��W�yy��'��
FD��4��J��Kf�����_�"���'���'��	*�M�gB���?���?�5ǌ&%+JT�a!�$�T�VI����U�O��>��&(<=�0c�.\1��"�,I���]���soM�c�PɛN~�S��OZ����{��ĳ1`�'iaFpk�T�2���?!���?	���h����]� sN(ɵ��1�r%�1,�*{���Ʀ�:�doy��n����H��}�KV�P<���mյRh���ߟ��I�����Ҧ��'��iZ5�[Bg�B	L����tS-u�����aޑ�����O����Oj���O��DD�`��,F���P1�4hH�ʓ;a��e�Q�b�' R��$�'�P�(f�<
�2���.B����d'�>)��?�M>�|�^����"E�m��V*W"���B�J��M0W����2R�D'��<�7NA�ʐl���mG>|�V��?i���?y���?ͧ��$�Ŧ��R����L�T�O�v ����f }��܊Vğ\`ߴ��'����?���?Y�oM�1\���� "�\���<��$�ش����3(,~�{�O�O-M�!e�\�fJ�p3čPfDK;�yr�'�"�'�'�r�	I��-@ �W� ���Dɏ#n]��D�O`�$Iئy��k>���MCJ>qҭ�m����ʈ�h��DB�����?A��|�d�J�M;�O�t+@��"є�����Cw�7>ݐ�X��JP?�L>a+O(�$�O>�d�O68Y�k�9s��P�$ 0G�Z	�,�O����<Y'�i���\�4�Ii��f,h� 2LAf�P�ǅ5����B}��'��|ʟ
�1��4e��� ����	3T� C^+�<ks�!�<�'5���	T�!n�z}�h��o�8����2��E�	������4�)�}y�q�e�F�I{����#A����Lոx�D�d�OJ8nZQ��A�����4������B�'�F��4@]�D�	�g�6�m�n~E@�iѢ�����K�{����c� I"�z��آz��$�<���?��?)���?�,�(�d�5�X�q�������L�֦�[1�ʟ$�Iӟ$?-����Mϻ����p1�`C?e�4pj����	@�)�Ӓ!O��l��<Y�K�6!<�)R���t�~a���<q��*�����䓨�d�OL�$.|��8)�ER{�r}j��2~@�d�O����O�ʓ2�6��7p���'-��$P ���$3�d��⇊:)��O�U�'���'��'�l��䃄>w�����Ӣ.2� ��Ot1+�EJ�e ���&1��H�X\lD�u���.D��jR<'`�Y_���Ѝ}�:UL\� �`�Vmx��]�]�� a���>�vyʓ�ۛ) ��f%֭4��+V�	9�}��%E�wd �a0w/�`���>)}qOrPiv�ߕ=.b�s�hѦ4Mt�kV  5gA\��`�޻I�Z�*���|1z���GS���)Ǩ(u$<+�"�}\"n\�Z֮ȷ	�أ#�A�:�<�p����-2���6,.t�
"Ny"�Ȱa��)E�@8c��D�.�l0��,�ZY�w��.L��h�`�_��B��\�?�Ȣ�g��� +yIF��'��	� $��ؠ}�T�CA��=e���VMLG�t�RA	K>���?a����s4��G�X*v$Gꊒx���#G�}�S���I\y��'V��'� ����	�~=�2�VhĄ�[&l��}�B[��������ImyB��.e*�Sq�*B�#׺4�NiR��A�&6��<����䓝?���i�) �'`œ���J�<Ă�+K�{׮qJ�O��D�O���<Q��݇,��S�����ʡ���c� Z�l_�h�2���M3�����?9��'����{BoB�^�,q��A�o��Z2��
�M���?�/OIq%��o��'���O�zU�
���Tr�Fa-zl ��5��OX�dq�p�'	�,��%�	kn����F�<mZy�
��~>^6��O���Or��K}Zc�u�t��T^X���DH��c�4�?	�t�Ʊ����)I�+{T���U8"��p�N1q��v��E46�O&�d�O���QF}bQ���� T��f�Ϸhiպ�,)h��9�Ѽi�:U���'��'���ĝ�^�n��G��>2�(�B�V�|�`�n�x�Iߟ��6J��d�<1���~퍲V0z̊Ǡ� �~�;�
���'�ޡqs�|2�'�B�'�Z�%�N<q�xɳu�^,c�	�v���$�T���'9�	ԟ�&��X�H�dI3��1\7p�'T�$�*�I�H�I>���?������pG�P�k_�YF�9$M��H2���e�WJ}�^����g�������9h
\�'����x������A�Ͼ��'���'�2R�@i�������h�n�c���AT�kfCC5�M�+O���;�$�O��=o��	_�5�2D��b
�1�A�0�Lꓹ?����?�-O�qACL�}���'�9!�-Z�!���@��&J��(��boӶ�D3���O������9}�JϽ�q�J>�d9�����M#��?�(O�1��J��<�s��*�*s�8��J�"8�� +�D�<I���?AM~�Ӻ;��C3��q��!�S�8��U�Kʦu�'�"<�g�lӎ��O���O^���H�t��+3�*��&��a�l�Ayb�']��$��2��i�$L�U�l�5
Y*ܾ(�ش(�����i���'��O7�O�),hk�$+�D�<W�����L�I_��l՟0�I���%���<����Z4�ϫ�j�Q�$�)d�>hcv�i���'(���m$HO�	�ON�	�~t��u�3~D��d�Ҋ0�7m�O�O����D�O��I�\7@ݚ� BRZ6��u�L'<�D6��O�8Pj�<�$R?5�?�
(<�Q�&B�n{�	�[�1�'"!��y"�'�؟Л���&L0p1	�Z6,�d+�eǹN2m�'{"�'��O��䴟����^���fG% Tfq��*�D!0�$�O,˓�?�DI������<j8D��*�f���9&���Mc���?��b�'3�	��7�ֺBA�5N!�Ȕa��ޜz��I�$�	�З'��EU��O1��хӡ}3�y)��`�H]cy�:�&��<ͧ�?9M?}X�?�P�cJ��;R�S�'|����<��_Ƣ(�.�v�D�O|���R$q���nh��
��@u+�����x�'��I[��#<�;Q/��ڦ�*��4!�?"�m�Uy�㏒a>26�_��<O�dM#?Q��$4vҴ��C�	�`�A�զY�'�"�'_��R�����O�FIÔkF)]�邢���Mc�뗨�?i��?9��,O�SO0�Y D'>��	��ۇ+�fm��O��s�)�֟8Y ��%[&=Ҷ�إv�Z�0CL�!�M��?��'TZ�r3�x�Oq��OJ�A�JS�J�0���n�.�r�Ƴi�B�|�~��?����?I�/.,2�q%C�5���LV�k��5O��a3=�4���0��}���R`���
 � +6�'���IK�	ȟД'B��nPx���95��R�� %:����V���Iʟ��?A��~r,Q���ȧ�Ot�
��M	�M��/�K~��'s"�'!�ӌxo�U̧D�n�2��	{���C�M3C��o�oy�'��T�	�#��j��z���L��t�kL�pz��5�
3����O��$�O�˓*]:��'^?�I�L�p�3!.|O�T3�F_�~F )޴�?Y-O���Ox�d�[�$�O���
5p��9Tܭ@v<�)��6!N�n�ɟ���NyZ`و���~���?���0�IIU���p2&��BM�_���X���	ן��	�o�����x�'7�i��QM��EnJ��v\�Q���D'�&Z�j��B#�M{���?�����S[���"U(ФJ6�W�UQP��48�6-�OD��ây��d6�D*��@j6@(�2U�FH ����7mJ2&d��n���	��������$�<��a�)�fh��(_&;�ָ3�����֤I��y2�'a�IT���?�N�6�8�SG�=Yw(Բ��(h���'r2�'^�i��j�>�+O~�d��[�kթL�p\S6��0�|"Эk�f���O��dвi5�?)�I럔���Uؔ!�vT���m�.:���4�?Q�NŊ.���sy��'N�����k�j}���]��Ap�,)P����� ̓�?1��?q���9O(X�6��c��PbAeԹ�c'7~�|`�'��	����'���'���	k� �C��?��
w�O�mM��"�';�ӟ���ԟ��O��h+<�I'��c�.�S���:BT�����i����\�'�b�'����yrN�5�P�H׋��M���1���6��O�D�Ot�d�<�e탦{���֘&nt��+�1K8p����C�7��OZ˓�?��?i4`�d~�O�s�A�O��1H�ƙ��U2t�i���'H�ɯJ�Ѩ�����O���S�L�>q�%���E'������
��`�'���'��Ƚ�yr]>��W�uf1|F�"EbY�N3U������'JܹsE�x�F�D�O�D��קu�G�\��L�Cj�4�z�G�M#��?�F���<Q!]?�F�'b�\(F��T�G-;8<oښb��Y9�4�?����?Y�'W�	Ny���:��k�H^�sG0L���;_5*6���(��2�ß|l��
�(�&&�ܚC�{4�l�ҟ$�I՟��j����$�<����~�dH'>}��)��T$I]>�j���9�M�L>Y���<�O�"�'� n�$��LF@��@k����6��O��j�(�H}�_����~y���5� .��@�>?��m�_�9�l;�P���#�e�������	��IOy�g؃L/,��R U��B9��l:DM�t��>	,O����<���?���w� �Hf�3�i���A!ʝ�����<�)O��$�O��Ħ<A7/�
���P��j�0�L f��q��ԒX��R���I_y�'���'0(ڛ'"�a��E[!�����ԁ-���� O�>���?i����d�b���O��E��TU�FN�B�4M��� <f�6��O�˓�?9��?�P-e~��M#��fx$��D��k�zP$oDʦ�����'�aq᫳~Z��?��'#�U����MD�0  \���I蟜���4Z&�Jy��'�i�Z�¸2�꟪8��ep�'V)P��F[� ��
��M���?9��2�W��J����D�5*ʩ�t��3=�7��Oj�J-D����O^˓��O:Z�����p�B�:�@),l�rڴe���$�i���'���Oc����DYP%���P�[A>!kvmW1��mZ�AZ����'w��䉞;���O�5� 8�g
X:O�B9nZ���I����!,_���į<	��~"ǍcV��B"#���1��0k�4����OHL"�0O��ޟ@�I�l1㋎��I $�)}F&�A֪�M����<��_���'d�T���i����j�!p.-�©G3���CȪ>�1�U~b�'���'��Z��
���?�p*��L�H,6���C�J�O�ʓ�?�,O��d�O,�$�JI鶏Ɉj��@�S�ǆF�Eв6O����O����O����<��,Z%0�	�<s9Vq�0� )g��Ar捵w#��^�|��Vy��'��'�L4S�O>��ňM�s�.l��/�(Iм�i���'�"�'A�ɹ6K��د�����r�#2-?UڞYbWG9#�}���i%�[�<��՟����'�F�B�d�
�\-2Rj����T#Ӌ��'�R�D�S�X���i�O*�$�
�GʘT�<d�щK5,�\��RA}��']��'eFiX�'�s�L��-,��i�c"l8�i
#È�
7֤o�^y�&ߑ�z6��O��D�O�	�O}Zw�h�	D�O���c"�B4)޴�?!��_��͓F��s���}Z�&=��Ez �rC�DÆ���q�@R�M���?9�������^��&LԜHjiX�i�1-��n���c�k���?)��۹d�r,0PF V2��f-��/��6�'��'�t�Xs*2��O<�Ķ��q��T@�pEc�n����{�v�OHU0O�S̟�������T�ۈc�z�z1�8��hsJN��M;��@C���Гx"�'���|Zc�$�c2��90��N�602�p�O�m+�5O���?��?�.Ov��q�%Z����T��m����ԯ>�]�>	����O���O~ ��ǋ8!S
 �b��(H��A@�Lڬ|�D�<����?a����s�t��'�VxS��b��Q�7�X�@-�j�I���&��	���t�d?q�B]�R�j�g��=SM�P�Q^}�'9r�'��I�U���O|ZׁG0U����s��E�zx��-h���'l�'Z��'�ZA���'���ȼ�t���3g>E���:���lZߟ���gy��^�X� �$��輘� !\QE����S�� 3�XO��۟��Ih�0�c��qڀKM1`L`�b̜�T6��
�����'�����fӀM�O�2�O"n�n��Y@f!��Ƥ"�ň1;`�n�����I��P��m��t�'bu6�Ѳ���'�0�FJ:LxmZ_4��ڴ�?����?���KR�O8���j�3s*�@[�)�j(�W�Iצ=0�g �d'��B�_�@"�A2���v��<� 4 &�i���'��8�O���OR�	"��I2D�*P��0J	x6m5�����?a�	ȟ|��+B\hҧ��y�BT�C�"X�ݴ�?ѥ,D>��O���-���D��6�Z��8��6��m�Q��!b�🸕'���'��V�lp�e
����C�Ub��X��Y�9��
�}��'��'6��'�Q`��ڬ_FH��Ųj&r�'bY�kl�U����؟���Vy�\qʐ瓖_�Hك^���ٹE��`˦�7���O"�O@���O~5�q�OƑ����-4z���V2���(��g}��'���'��I�c�ZxQN|�t�[2�J&��'WڄPG�47��V�'��'oB�'�dH��'��L�b8�w��v���F��e:hoZǟH��Yy�Q�x�����k,	v<h�m2)JiCS+2ױOX��?��Zw��@ӱm٤�HB��ۧA���[ߴ���C޶ n����I�O��i�`~��*p�)g���0UQ�G����d�<������'pq6�3M�;��H���ѻ3
�$m��h��a��ߟ,�R��?y,O��� 4�I�����7���\x}���O1���Ē�"t����R�ذ�#)�.{��o՟��	ڟ��3��?���|
��?����*>�ʜ�3��5�X��O�+ƱO
,+��D�O>��O�|�	?4�xѣߪ:���Є�jyr+[��?9����O��O2��v�O�NY���!�X��C�-Yn≃eN���?i��?���?���h�6��dC| �ԉ���'O�-��?���?q��䓪?y�'���+����Ɲ�A狀R�<,�ش�̍�'<"�'0�Q��#��8�����[��3���v���������O���O:⟘�r�~� *],2�(���ϯ5�89wS�����L�����	�,��D��ڟ����[2�G�|�vH��Y6L�b`l���$���I{yB�ݱ�ēR��S5@�?<�&��!I��;�mlZş0��dy%��)�����$������O��hdb!+�+�!L Ӏ�@�	Ƛ���O�#<9�O��l����*s��y��HW$Qo8Da�4��Ę�W�d�nZ��	�O��I�h~�НV�vlz�-S9�^͓��_��M���?I��o���OM��a%Aw7����䇹H��I��4|6�%�վi�r�'��OO�O&�$+�JՀQV�=�8�!���8��mn<h��#<E�$�'�jԡ���8ҢyY��=A>8���q���d�Op�$_�tV�5&���	�X��7}��ئ��6z�)���Ĉ;��(�>)d�P�<q��?��{3��P��I>`��rE�V|���c�i)�d�M��'z매?�J>Y�қ^�D��/ҏk�ٳG�~�'(ډH�O���O*��<i҆Y�E @8q�`�b`U���	m2�3�x��'s�'&�OL�@����'_(�4�N5�­���&U��?���?����?	�L��?9`OK�\�ĀZTǞ�ISf�QoX�`~���'�"�'#�'�2_��TJh�<�scKjڬP�3M��jQh�V�P��ɟ$�	[y� H�J����܀�� d~iR7"*��͎�5��k��ݟ0�	
PDb�d���DR��iC��8b,�od�<��O*ʓ1�|�A��4�'����b.�8��I�P���3�A&?�DO��D�O�`	7�	}j�bߋ5��e��'�1�X��H˦�'���d�`���O��ON�%�H}I��F�C�U9�*ԁ{oZ���	7R�#<�~BrJ�E.u�VJJ��C�Ȃ��!����	�M����?����֕xr�'R�ㄨN�"-�e��#��X��-��){�H���)�'�?�V�T�d���r#@P	*P�mӛ��'�b�'�t�b6:��Op�d���ypM�5k���LǛbNAs� #�ɶD��c�����,��5=](� Ό�di��A�H��6V����4�?�0�	L�O��d1���L���A�JEYɧ� {8�	�R�,"*���l������ΟlCDj^�^�VQ��/�7�$psV��
7R杖'���ҟ�&�t��R?)t@�}TB��P���]n�1c�eRզ��D`5?���?����Ă�l_�Xͧ9�&�0���$$�t�� Q^�'�b�'�����iE��+	�(�� ��1?�>U�h֧Dj&ꓹ?i���?Y���?��!������O QX0�UG.N=�����!3�DQ6.��=��m�	ڟ8�'���bN<�S��4 @����XԵ��������	˟��'�H!�):�i�O\����k�1B���+1LA���Y�[ξ'���I��Yc� ���t�^�>X|Q�cۂU��M�4o���M#(O&� u�U������d埮H�'hB�bc/�F�l���h��AWά�ܴ�?I��}�"�Gx��� [%#$ ��--L���Q��?����,3��c��?lO��9��٪MIL ��E�,�D@�a"O��:���A�q�V V�;���1�l��Y�x����dH��Bh�i���{4��U:��*�Q�'��qn��M�(�VΟ�9��	:3%�6�2�q	�`��I{�J��9G
� ¯���Q��̚�-�����&�*�B1��t��!�!��t������#c0:5�7�� <ЈPn�O��$�O���ĺ����?I�Ot\�q�D�ܙp`���4�X��g��$�l0w�ٚ7���b��	4Ny#?���+
����A�F[P����.�欒�M�"h�\����i<��E֜c{t�BW`�tO��b5�G�wz�!�2{V\�K�F.d�R�'ўt�?I���<B�J �͑��ъ�V�<�c�ϸB�:�S2����b�Ȥ��K�sm�IXyr�|:�^��ɘB�=!1ă%G& ��,B�rs<���ן�R�oB����	�|��Bͱb�f����E�$��!�~��Q�	:��Xr"���x�KJ<oI4�`Qd�(%��	%�����O�.��:�KD�0����Z�>���'��I	76�L�ℍ-��p�i!24bc�h��	�}~|�P��#L�� `fgU4}�<C���M�G= C��R�m�]ǚ���Z�<�(O0%�C�W}R�'��Ӻ}.� ��l��)���U�b�v��c� <A���ڟ4��I5VV���F�[���|(�tL��߁AmX9h���3� A�b�>�"$�9Pt����gٖ~�Q?e��d�����ɆEP,
�ĝ�m-}�m� �?����h�>���!y���26�ݶni,���>m9!��<D�>��V�D!a�0����m ax.0�n�t=����rH�Q1���p�}�&�i��'��S�uL0y��'�b�'��wW��C�	K�a1�BS JFV�f�|"�y2E�%Vcr����/ǄD�t�,��'|͛ϓv1|�w�_�o�<�C��U�qin9�y�@U��?�}&�������P�f����5��+D��V�
X~T��*��:5S��;?QW�)�'Tp�aWC�-E�d{"���'�:���LCQ8�Z���?����?qG�� �d�O�擢:	� ��JӁ��2�!Y�Vf"H�$+#��3�O�x*��J��<{$�{����:�4B���z*pMi���6UA��z�4�҉�O8��䟇gL*f�<>ܸ)Q�ԍ}�!�d� ����b�F5;���v/L!d1O8�>Q��L�O���'���\�A���RB.	2g�b�'$X���'|"7�8$3�'�'nE��џ+��3�����8Ǔdv��?Q�dL-f4p�j�;aR � Ma8���@�O��OfX*6��)4������ �V"OL��0�%'�|��g׽>b�avO�9n��M�t������0�Z1�91��c�p
tg���MK��?Y(���˂n�O�5����S�`�Xn� 'n�O��Ø&��D �|�'6�9��^ha�+��(�ԚN��˗�)��F��Pfj�#e\H�E&�<�r�'μ����?�H~H~��B�j���U�FKX���S̓�?�ϓ&;��Ч�9b�U"$DُT�N���:�HOz��0�Y0@�Lp�2S4"�Щ������џ��<I6h�[�n��p�	����iޑ�7u?Xr���.��|�Fy̓?�$��I-e�5��?"n6�����|�r�P� /<Ob)�P'^0w	�#4G�A�BB!7扊C�J���|I�,!��G�E>i�^�)`DY�y�gϫF����BW�	�J1�b�ϼ��$ZQ���$e�Ƨ��7kH�@�Z!wGԈ�$HN.;.�ɴ��O���O�����s���?��O�2�JJ2pnE��į�x)�t E�x�G��"�h��z�d�
p'R����'��w	S"I�r���/ �)a��ѷF]��?���)K\0I�		d&Ēhת-��)ޑ�խ6t��yS�]2a����<���s<moZ��	<?|*͐�~RN89�g:j1��ȟ�@�Dџ��	�|�g��%�܀�m&�U����Eq��L�p<��v��������T�5�te�veڙ�A�㉏Q���:����Tۜ�����h��Zl_	�!�$X�9� i�c����I1��=^�!�ć�Ur �*${d0��ٓedR�-�	U�Z�4�?�����Ȼnh>��S�PDfabā�
|����	ۍ �.�d�O���(�O�c��g~�l�F�r���͈�c��)س���I���#<�z�@@�B���쀢)�h�m{�� EW����28s�1��Û�u�̓ U�>�!�dCG�ɒŪ(E��õo�(l�axB�7ғC�Bj��,BmR�X�F	V�+Եi&��'W�c��jGr\;t�'R��'*�wLj���ޝ?t0��d ��h4����X�9�yҊ%k�,����M[C.�0���۸'P��9	�� ��Q�56�~m
�i�/�R@�y����?�}&���R悆s <���S"??�8��->D�Tr�G�&����`M2���U??r�)�'��p�ˈ/(�A5)��6V@��X��P��oٖ|̼i5�A�h���T��sa��?�J}�3�ˇ�&��ȓ�R[a�\so���p$�?p��ȓ?�*(R�m	�5�VQ�Oƻ.�ՄȓJ�Ĝ�u�+{��fŀ24܍�ȓ)Fe:���@��m���,ƕ��$��y��-��$mD�I�̈́�2�X<�ȓ4ڐa�3"Ť�t�w�T�:�ȅ�a1�9��djح��dW�y�$���p��@FyV2�H�fsKx�ȓ ZlmJb�>�f\�v���c�0!����1'�;��8 'R����O�^��W���DJ�X�3T��C�	1h�Z�y��K�8�qaFײcxB�AO捃�E@��4�맋iC�I��iBGN�|D$��π�F��B�ɫ6m�W��t��U��� ��B�ɾB � g]?�x�x�C�O��B�)� �ACg�X	^|d2���Ť<�C"O@�c1fC�s��s��ɸ-�Э*�"O��v)�DZ�q�E��$!�r���"O89�!S�* ��Ӈʝ�2���"O^x����vH��Qe,Ҩh�<JG"O�+���'�ذ%ޛ8cJ��"O0�)�iN�E�r�H�%O3"�T��T"O��[J�LL�Icn�$�v"O<9���(A|,���D+j�&-1�"O,�F$)1ڕ(m�.g^�9e"Op��>~���K�PT��k�"O�1�f��B�TȻ�I�F��3�"O�!���I�^̰wg�%1�B"O\�Cv75�<�+��XH��"O؉��j��i�jѓ�	�X-0"O|����<_7�Q�"�6�Zt�4"OzL�GERG]��ȡ�EY���h"O,qf��t9�D:����z1x�"OL!����"�ʘ9q��#O�^�'"OAc�2}��a��^8����#"O�Py&�OJ,tk��%� ��#"O�j���D���(4	K^@=k6"O~���-Fo┥sB�J%�&"O.L�+^9[���Kd��j��Y"O$��Y�[K���O�'H]b�"O����#q/�<2���d0����"O���8!�͑A�Ոw��"Op	��HT,tώ�r%���}anɑ�"OHcJ]7dܴ�&�y`Xt"O�9Sg��*~Lb=;p�0D�,����&{a�>%?�B���2,���b�r�6� Wn?D�C�I�m�-`�M�6T����N2F������<�*F4C�h�zRP�4���� _�<�$�k�����cޑ��Y����Oj0����M���ّ	 �^��`���E2����fa-\O>2�!��$�q℉��'A<x�Ύ4Mў-{��)G���K9>Eq�=2�x1Fĥ��'3N�Q�&��8���DȔ|c��F)^HL	��'�� L�u�S�O�(X���̬c���z#ϔ�k�����"O� �7k�<Y��h7kOl�K`T�D9V�ܮTa{��N2D�J$xc��(Rܜ��2�
���>����bt�6�Hi(�1R�?>��4�eH @!��(UrbT��B��h�!خ/	�Y%JO��H��s�ܪ=i\p�&&!L��6"On=�4��H֩ZV��2�N}�B"O�t�e��D��2IL�_	�e"O���A��8۱h�$	B}#"O����m��`{������E"O���g�+R��� �F�4`?LI��"O8]`��V \4��c�Ċ5�ؑ�"O�{��P�ؓ�Dҳbg�1s"O��	-$�Hd�֝Y�"O p���Ȫ.��`Q� Aa�]å"O�� ��R1xě3Ő5OT4�4"O@��F�ѫ�\:'�[�$�L�pg"O$� GZ�=�$-�s��0�@P"O�$���ېk�L���V��܌8R"OȨ�fU19^��FmӴ�� ��"O"�ɢ%K�)�󇊐;>Ψ��"O�P��B�7M� H�˙6X��R0"Oh*�G� ����#���T"O��P.�����k�6
@�Z"O�QT��:oZј�H=H��PB�"O��J5 !5�0кcg�$�B���"O� �-Pe�&;�H��6�ߏ�=0G"O��;�aK�-�,��R@&K��-�2"O�Y�H�#!�R�[2���,�'"O�`!�+�Y��,��j�"O�����T �+��j��"O��ƔP��e� ��3}WF�s"Od����X.�eQ���9
]pu"OlM��+Qy�!��^_�`�"Oh�{�']���[�B�3
�ź6"O4�ѣǓ/�$R�*�J��"O�E;3��ܑ	#i�~�=�1�'n����͸�N�h�)ҕB��g�cb���ȓ|������"L�����kc�E}B�N�|�0�F�O����E���	bXR2��pw����عU��6��\X6\��A�ލʐ�%�)�'x14�gO�n�\�B&%�*�L��s��V��j[<a�6΃!)�6	�O�X��m��0=9a��4�ꐀ`���}'J��@ˋc���b�nwBUSa@�)F3`{e��'-�J�qs"O4��bʀ)N"x#s�"y"�2w���Z �,�b�S�+��PF6��B��5m�B��\�����Ȏ-`����E�v�ɥA~|!sd�O隱Vc�O� q�҆Ҏ�HQ�r@W}�f��	�'F�tB�m��|
��ٝq�Ha�J% �&1x�ƢT��Y����C*?Cđ��iߙM���pa���ab@��Pv� ���<q >��/R]x�{⭱��Cp�F�x�a|��Q�8F���i	fe��o�|"%��ybZ��9ۘ��Q ��14
���F���O ��p�΄2�2Q`gc���aEy��G�E�TB5#�Ni*�k�4	�,� i���y�(4@���B�U4�H�f@8!
��[��������Fɔ��ULŕ,��P��늵�y�ǇF���Cg�&X�=�fE��~�o�>k���I 1։�L�	_X(;�ӋSBa}� [���Γ-F�uX��":"$za@Y%V��ͅ�7�f��RX�>I��h��|l�EyB��3�v�G�d��DA�Mك�K�g�l5��MR�y�$L�f���ȍ0
r�:��`\a�Dm�ɸ���R����Ա��l��,Ѱ,�@+�,�y�8F%:s^'�Y;�M����0>!�h�p�%pRoR;6��JV�x�<)�(ٷ;��[Rk��g�Ld��/�Z�<��Jٹ�����N�����C�!�y"kߑL���h�&U�Q�4DYQ��y�G���db'd��Kbu�DG��y⥙ Q9�4�ubЂ��H�/ĉ�y ��!.����DȤ���E���y���)_�T#��	�xb$E@/��	Z?!�EA-���z�wX��QB7i��ᣠC���L��66ީ��D�^�txz��ɝk�ɹ������Z��u���U~B�A�j�}�'E2(M+��.��<��E ��D!F�F���ǕǸA�a�-Z�r�x��n�r�z��)OH�i�ᙺ[��=)��įjV��#�|"�ŭn^�I�'jnd8��ԮY�v�2S)�j��ĸ�/Q�H�jCa@ saB��V
&����C�`%z2A"�����>X�ٴ�y�8O&��M� ��|RE�ǄE�ȐSSn��_��0tdMG�<��F�����Ξ25�J�z��ܮf.�"��n�	���';J��)U�]�~2 	4C���vG�LY.���BT��p?Q�àdP�Р�K�y�n�[q� 65A2١S��O�%��变UW
aQ,�=z��Ҥ�Ik&(����)W���&�u�>�b�R�P����v틜k���Rq�V���y�����	`Z���a�!��7I���'2��a�{��!��BV�Z�r�'5 ��`QV2��AA��};p� P�<�M?�h�`�3St4��NHl�p�c�-!D�����"NLt��ԅ� (Q��K����)��\'���U
<�O�t��t�$E*�)� �!�EYB	b�A��x%;�'I΁���D&nz��I���{F@ބ=�ᤃE��0#��Ā�dL��+Y0�X�>ɒB�@�.P��.�W/D@[��j�'�x��n.� {�N�u�8�ɔN��v�a� �5w$�;�L]8Jeo�A�����F�
���l�/�pIBb����8 �}�G
"3�%�r�D�6>����718$�H��6%��!vT��c�]=�ubt"O�� �T;c���S�U�\��}��>�5��d1P��`�xk_�r�(�Q?q���ʾV��PB�_�z$�pd-�O����Q�;������(<�36�Zk~������}�dW����w�|�![�+2�`��[0o�:`����O���Ew̓hݾ!A�U��"�r��	��
4dLJ%��,3�O<I�p�9T�<��*P !�c�Y�P��l����'��p�rd��D	���'���3�L�`J�+�@G�A�Ƚ��'�T\q���,���Q��_�s����I<a#j��oR�A���O���ɋ#U�<(���n�B�d��|J���a�V�����NX��r�I�;Vg��9�"O^��� ����D�O�>K��V"O���R��Q�t���"O����+*���T�r�vY�"O(�B!c
��}BT��9&�!h�"OX�÷D�vMʴ�$6|�D��W"O�� ��13���;��U�~J(�y`"O�lb���&��BId0�@�"O�x���I Q��X���;%�"O@C�
�n�B43f�ܬK��"O�S疤<��\��Έ+r�z�"O,y�鍈}o�(ʖN]�p, qc"O��X�m�*��K�-ٝZ J��"Ov��fa�!:�hi��l��
T$���y	t��%��K��Yid�����y�ϟ�x����P5���y�i�?X�\P`tfK�Hc�����y� � P�|���DΓ�\��2����y�LU(0�e��D??�@tH"%�?�y���P�.��!��+�.��$���yB�]+Q�����C�Uzr	
��ڸ�yBd�8����`�	�R� �U�-�y"�޻#�~%�u�L�K�� puQ��y2��[U���/M�oH�|�4���y�MW.'-�䘀�31&,�����y7g��+�L"�YS�Ǌ��y"aI�=ø�8�Ɛ
�0��e,���y��J\�H+WƏ.�$�
奄 �yb̌�b����Pp`$Ղԋߺ�y"�ޢ>1�U�ޭe�.`I��M��y�d�
[��3@n��%�8=�%�ˏ�ygY�z8�%�Q/$,��D[��y�e@� ��KUǒ,Ʉ�8pfݸ�yr*N�H��W'�*>���IR��y2���]pBu�j�":���D�y�k�-3�ܤ�S(B�!>��[�N�*�yBnZ1z`�YH���s�e9�a<�y�e_V�E��!��i�dƿ�yb$[�Q�ʭ�¢��R 3���y�!�f p�+��z��E�R9�y�c�|4����ێg%,īCN
�y�r�,#��:7��t�ahJ�y�I�CX��ȱ2��[�����y"��mXŊ���
x�,���(�*�yR�A={����0m�r��w%���y2��	�x\� J�k$�a�Ƅ��y�U��Դ���^�z�r|��yJK(<�ȕ����sTBu�^��y�m>t�A!�q2:�q��S0�y
� jЊԥ�uT0r�^�P�)1"O�p�F�!\d&hᅉ��7PT�Q"O��z�X�qzpH+j�y4ʝ!�"OF��v�˫@R��0)��V(����"Od��������2u*ЬRHlx��"O����ؓB4�BW�%,Ј"OD�T�.%\5�"��V����g"O"��e��0Q$}�l�bV���"O�d��J2T�M!�d�?�	c�"O�R�mv��Ś!䁤G�B\9"O�,s�I�3C�-���җJw�X7"O4ibI�"L36隄j�F�"x�""O���.V"^8h�'��`�P]j�"O>��QDR� ;֥Rf�<�}`�"O��C�b]�/8�`�1	�L��"O�x8�.@�Y���!�e��	(��w"O荱VoY#fP��FR.f�����"Ot@�oZ��d�F�~�Ɂ"O"� wB����O�'tux�"O���q&��1�պ a�7<����"O^�ەɒΛ5�?e\����;,OT�<y���5��82
��o�y�`p�<	�̂fLfr&A P�c�l�<�eMT_(]�2�E�Uٔ��*B�<�D�D*L����``4�}ږ�Tv�<�Cސ%�E�G��1*d2��f�<�hݨt�X�"��N�+BR��d�<��9q&e"�Nc*N��� �u�<��#�< a�裲l�w܄��G/�z�<���B��y�6AK �Z����DM�<iFO׸\�P�Po�0 ��m�mR�<AW�.{#���c�<�du�Zq'!�7Owи�qB�n����F��!�ć�M$
\P�
��v�!u�I�!�dG�G�Tu��V�u�� ���:*�!��U\8�Սm��8��-ݱ ���Dx9�g}B�>K�<��SgT�7����'���y�IH�^�� ��b�D�����U�v�(�$�O|�[G���&pƱ Ef[�Fo*��"O� �g,P��@"#�AD����"Of���j��x` ������g"OPi��k�>4�����r��Q�&"O��q7�Xl��+�C¼N��+ "OL�@'FS�Z�X��@˩�T""OY#/C2~�j}0�4n#0!ٳ"O���e�ݖ:���#�ĎMA�m+�"O��j�Ʌ ,Zfm���GH9��"Oxl�u���+�bEQ�k̞D��QZ��� lO�Y�
O�nZ
� 8<8m#�"Oz�A`
ڙ_�~���v'�\°"O�x²�T�#$0�#��(��i�"OZY�D%�bY��m��6)��"ON�Io�SJ~��"6b��y�"Op����`4��aG!x��3�"O,A1"�_ZRx��m	�^>�
�"On J�Q�^8�K�p\���"O���Q#QJ��k�	.��U�"O��ʆΟځ��j��X����*O�0���#,��0Y��w��K�'�Qsކ'���j�j���
�'��H�,L;e��MI�k�*i\h@
�'%r���� 1�L�-Y��S	�'Cv`��-�6O�Cd�Q�AW�$��'���+�D5t�C3/8�p����� &�ل�Ԑ)��C�Eۼ\�5�`"O���&O�Y��5+W�+� <��"O<Lx���wiZ��M/	9��b"O�ћ��	�0�f3��+!6Hʵ"O@u����:��#kY�~>�5"O(��2%l�1P0�H�F�:�[t"Ol�c�HX��]0
�}h�K"OD� DI1-�ru1�h��6����"O����?�.�)�K	���"O�1�4ʊOm��pԧ
5-����"Onl��%��d�d!�Z:Q�<c�"O6J��`���؆�׻�UH�"O��Sh�WHT�%Nн[DS�"OܥiG�^�V���HEZ1| r5h�"O�`��$ �n�����Y�*M�i!*O�*5m��f'��q��GT�0���':8���H� ca5��� 	b.QZ
�'�(�(v琧 &@�AA(X�� l�
�'���RV��A�t���y$��
�'p��UIȣVf������j^����'%�����7l����L'0\�Չ�'6�}��o�<��d�3k�/NA��'a҆G?9Q
���F��-T���� ���y��Yl�B:�ʔ��(�8�y��B
J_�� �*��e05��yb
��~uj��!?`I�*��y�$����z��87r������y�K��4�}(G&�mz�b����y�S )X�(#�F��aJ��y�/�w%�u��#H�G�T�;��ܯ�y"�\�Hh�=6�͘?�<RdŒ��y��،i���6MD���I�r���y"AFtO��4ùp�R���eW�y�������9T�U�\�������y��7��Q�C�U(�����yB�N`{�N��J� ec�-���y��pf	9$�I!;栰���*�ybO�o��=H#�ʐ-j,�s�$���y�%�dEɃD!9��*�#��y�+�60_n�,�)�ԚnT�yR�`���
3����-� �yB��I�pͣ4Ę��*�hX8�y�dD�ty�Y&�8 �U �♓�y2)�1B��#Y8^�<
�H"	�'Fj1fcQz�`�kW(J[Ƞ��'�b��'G@�w�z���>�����'RT�p5!�*����(	�dj�'	|	�4_��d�5aH% ���z�'��9{��)���P��F�/,�i��'Ɏ͒0F�:t��a/B'>���
�'n����J�0�a��I=0	�
�'�ބ�#��6�r!Fx��� 
�'H�1�p��)��P�k��$@@m�	�'vFTE��^�f�ۑ��N��`��' 2�C��7N�n�Xnއ@�Z���'t,�3�&�L�):���s���ȓ�pTa�-� @h��G6u����
����F�(�(�kw���'�6@��\HN��Յ(P�HC�N]\���#�JA�a�ơw�}⠂��3p�م�p������0X�jf߇fꬅ�kR�F�V�tR {�.�rf��ȓC�����|1��V�=h6�l�ȓ.�Pu��G�z����t	J@��S�? 6|k���'M��M��D�1"��"O�!�+�;4��u�3�� X��!ȶ"O�`�p.�g(0�a�@�"��ð"OJ�a,�Gn|��MX4��kv"O$�yA�1 �0���ڷ#|��B "O�5��\�@�Cr�ωmP����"O 5`���D����Bi�y�"Ovx;��?o��͉&cv���B"O�Y�B�X.ܹY�(��M��"O��µJ�(�9D�N�z-��"O|�
�mDRq 	�2Ol���a&"O�!�S�+>l1�tT��y	"O:q�v�%	#ut��S�$��"Ot��FQG�x��I;dw�px"O0���ؼ:ְRH�$[�p1�"Ozt�Ca��0��SQ��G�R	�"O�a��(��]�\����	A��$"O\YS�㝆=��M*���I��M��"O6��aق/��e��&��j`�b"O�yy�	�}" �1��H6&����C"Oj�8gk��QH��� 448ԸF"O�L�ؘ�$�2�]�=�����"O��pQF���!8Į�p���z�"O0��7Ѻ ��0����1y�"O�|ڡn�,�|�{&MY�	\I�"O"T郁��w�����"{^��b"O�Q�B7)
�-�≌�T�x�&"OXM���0RIP��(�̦�3"O���a&����:2��'m� ��"O\��A���p5�ЎK��%8P"OZU�%b��>qpM���Ż��B"O�ňc��Js�d��6�H��"O�a��ʦ'����K��J���"O���dm�r�  +]���,�y2���<�Q$E�2��)�	H�B�I�aV<}9᧟3�%r �&\�B�I>k��%9��ˠtR�)�@[��C�ɍ_��uA���;|�&����V^�C�I�������^0T�a�A�׈=^C�ɲ}��JC+�u
:\��,�.k�B�I_�0|1��
4�x�:�,~��B��4��1K7�*UGpA�G�J��C䉌ixdm�b�H=(���>��C�I�2P�4�rfļ3��m��d��_��C�&�V$xe���"�5B�q��C�ɂ ��9��*C�@HभΑ |@C�Ɋx�B��$A)�8��3�̭�C�	�0�=�Qdž
��m�B�:U��B�ɡ2�⼊@I@`���G��-;fC䉑_������ ~��샦���z�B�	� �+U��QV��#�jO�=�VB䉂.0�R�AN+=�p ��
��g�B�I�% .C'I�Xw�1�bJr�B�ɢ3������
��vjF���B�	� ����?o�<x���
J�<B�	c��@�#����Q�H�\��B�	�YD�S�	E	]�K��T6�B�s�b���Uת(s��G�XB�ɯh"04�ԮL�vA��/A�t̀e"O$���T�H�l��B�#~��)x�"O��R���9W
L}I��q2�"Ox�:���V��	�d�ՃMs�(3�"O>�����l����2kdԨ��"Op�� )M,���㏒�Eu��	�"O� $9&/����Y�`؁?l�!"V"O�%�΀?{� �C@Lv<�`h�"OZ�r�.#� &��	/1���"O�e�'I\�)��	pg8G�2A"Ot���|�lC�F�|{d��"O��@�É�Z\���p͍|S0�"O�I�q	��v�z�Dȅ;��l�a"O������8��!3r
��<��	��"O���2.�V�m��n�,1��*@"O��q��Tj����m�Lּ""O0P��un�䋑MO1��D�7"Oh�c&
4AY���7m��B�H�Aa"O y��H��Ht�&́�����"O���wj �ӊ�w���>�hEȡ*O���2DI�Qr�SbEZ����'E�<*w�F�0���0%H�ef�q�'ڦt�6�ˆo��(P�ZKLĸ
�'�H����z����7��LZ:Hz
�'|`���S7��y@�Ē�t?��	�'�:5
�(���ѣ��:�,`	�'��d��f���I#�Z� (��J�'�n���FM�M�@���-IE<�X	�',f�KP�Z�����mG�3& Q��'�p6�Oe;W�^'+T^!��'S~iz&Q�9,V�qv�
%�̜��'G`uYA�b�~�X(�g�8���'=p�{�ֹ��(�B���[����'�.eK�Ϟk�ph���I����
�'pܜ��ڭ
���X�`N�ҙp
�'�6�) �A�
f�B3��->�4��
�'x"Hs�K\�f m��j��Mtv�1
�'VD='�P�5�<� U�Sn��u	�'֨Q٦�U���*J��|mMޫ�y��V9�����s���vd�*�y2IX^=V�NSP����yB��(w���Bb*5?�$�{�	ʏ�y�I�+9��aÃ�ۚ1��xj�I�y2��/+��Ս�'��H� l�%�y��*Fhr�Pঘ�u �C I"�y���roaբO*s��1S�/�"�y�n��4��4x ��i�U��yr��	vR��*�3k�ܐ��&B:�y�N%�R%�0�X�a�0����y��8 n5��G2U�64��d��Py�ț�X�a@�=J%B�7^f�<)#�\�����Ӱ4�ô�NJ�<�x�ܵ�5l�74t�4�L�<Ap��%!�YW*�+t�Da�0�AK�<�vڇe��L��nR�|
b��D�<���J�T-�q�֤�$:F�aaFHF�<aQ��+"����d��86
��{�<Rឈx���a� ۭ3���D��<�"�F<���+\�(�.KD�<)s)�x�d��g��'M�̸�)T@�<1��Y�1�ީf��L0�g�~�<�\�ՒC��"yHл�!Ei�!�_�t�|Dp��[	��բ$/A��!��'��[�A@�Cfn� �@�l�!�d¤jg�����5Wy(�o]��!�X�y�ꡊ b�	@����M�I�!�X�1��+�3|0���͒�W�!�,+2��
�?�V��!�!�D�{��񱏋�L�S�w�!��3%��b�Ȍi�.�p�lC�!�� h��Im����,��x�Z�B"OduڑgӶHR=p�,]�U�v�ڃ"O���P,.<:L�ckN����b"O.�#S)Ӻ���C�����.��"O��R��.�U	�E��EcS"O���-�+V�ѥ&�����"O`��VC�!��p�e�q�Z +�"O�q`��[(��x���P��4a�"OnU��dӄRK����L�m��Ш�"OH1 ƌ���Ș���l��H�"O�3��]�z�v<@��>]"x2�"O��i��P�K:�i[���sB���a"O�" �6[�T���'(��"O`��3jY>[72	K��T�� �"O�%��&Ǒz&�� MRwV�x�"O��`�0BL�����2#�"OP�Y3Gڿ.4��*FkB}N4җ"O�jD��2HYvtjQ��5n!�"O~ ��Ô�M�2��㧓�hɱ"Ol�4
�.?�L� �а��$�"O�a��Q��Mau�G�42"�ˤ"O�QR�QU���9s��B5��"O&�� !Ǉb���k����u��P"OD�{���Y���A�;l�L��"O�Ys�T�uab�s��H�Wl���"Od`s��?'2��w@�/YΝ�q"Ob�D�*b��)j^��$��T"Od�`�g�\Ȣ�ѯ�L��"O�Ix4�[.Qr<���WzDe"O����BؿZ�8�C�YT~���"O޼!7� !L>Qҳ��/F�e��"OD�E�ț
�}zt�G��D�0"O���@�,���k�N��l �!�"O^���NXE)������s'"O�0�V���*�,{�#"0� H�"Of9B�*BE������d��"O����A 7F�� �"��)��"O�� Օ1���h�*�j�	!"O��!�K�5uU���"I�!�����"OHX�$M�luukpJĐ3���23"O���_D>0rF�� 5.����"O�AyъB2`���C�HYH�r��&"O=вD�P������\�!��<� "O.��ǁ�z͊f��i�@��u"O$�B�� Z��m�I�a����"O�<8a�:$�	��@��rĻ��'B1OB��h-�	+B�� �4����=LO�d��%��N��rȼ3j�`"O����[p�^I�4O����)��"OM4�BW���
I2��ش�|b�'(�("E�+��	G�N�STz���'��t���n�ER�"+O���
�'bT�Z�@N�ul0�B��s��u�
�'^)`��Р}������ /��
����эOT8ć��P�z� �<�!�Pa�@: ��U���L�����'���{ƩN`�:p{2g��F451�'��XZf\#eO"�KB䑵qWޝ�	�'�x�;V4� �ˠ/¦W#� J�'�6���S�7_���w�~w�08���#�V�X���z�ea��=I<�a"Oٚo�
G��0�5�C�4�"O�����&xT��iUE�Z ~UY�"O6���~S�ңDM�> ���"O� rtx�&�/l��ė�N����"Ol��v�J���j�Hܯ
�Us�"Oy�@J��a��=��)�*	�t�D��&LO֍0�U�|���pH\9h��,�fO�]�5�=��� 4OM��,���<����yV"ЯF'��K�D?M���ȓHM:l�7�Y-/Lp!IP�!��F{��O��D�T+S�A�֐+��J/$��'@�u�f��h��C5�@�'��e⢀�._<�K��W�P��(�"�)�ĭB�b}P8�˂h0*M��P��y�(�pd��V�g��(0��S��yB��n�"�XQ@
��|�R�ۅ��?��'�ND��K!#eh��b0,v����xE�P���Z�GI� ���R�׺�yr��u�2�y��Q�>eJ�����y���?��*yp�	H����ybB��m�U$J\���#E=��7�S�O�l��Ps8])��<�H`�ϓ�O��惆)@���Y�TG\3�'��Ć�tBQ�
�G��y0��J?!��ʛb�L`�7��==$wI"b!�DT7Pk�T#'g]5��KGa]5!�	�"������4?�=����0w!�$���ִ��+2q�4�%�?f�'ba|"��'z>�D�f�S�4F8P�(E���'��o�'��}K$�Q&������d�����"O��z���_���)G�!=R,��"O��1��TE����-$��"O�������i�럎w�B̃&"O �S�b_�G�,qkC��<ZƠ@�'"O,3rO:3G(���V���$#�S��C!8�:����bբ��"���!��5@�# �-���g��#���?�5G5����E'I8��G@��yb��T�|��:H�h��H�?�yBb��F�2i�Dɛ+JP����y2h���b��W/5 ��1�mA���D/�S�O�V��vEK�wJƘ�� B��	��'�fH�B�%E��b�ι<�^���'$��2�Cӑ{���qpcYCax��	�'��T)�۾n38|� )���q�r�)�t-��~ Y�hغ�"�`�'���A��X
x�Sw%��'��j�'�P}�5.]�A��8�ؚ%b�Y����'s�>��w��ͅ�N Pe@W̆�*5��$�. ��H�#�F8�L�CP!���_� ���!i�D�c�"��E!�$ˁ_V攒V���
��e���U:=!�׻%�PR@B�k�D�K���)!��-��A����G���ˤ�8/!�$�-R]�Lc�"�D"�D`#�H�W��}b��x�/�-�2�SbO�!<l%i��4D�4A��'dQ�iuL��G*��S�<!-Ox��dֿü���XP�c��]"^!�$�g
N,����m$�@�BlI��'Ka|B�)Xv���-H� ^�����U�y�I�!�����I�Tz��#̜��y��@� ��E= Q���&�hO���O4�`5FG�}8��.��Q����g"O|����Z�^]iUjh���\�$G{��IρGZ�M0U��!-�PU N���!����j�9�o[-;�<�(�+]�|�!��z���TL[l�DB�
�f�!�� �U�`c*��<���
0vT`S"O�}�2�?�4��@��	r"OHqP  �7D�n���)	�D=�d�'#ў"~BЍN�dD��B�
M#8��Oݟ�y�� 
����FA�^�bG�L�yB���G��	4H�!��|{��ʫ�y������0 T�s�Ï��yrMսb�&��b���4��y2��{|��ZǨ��F��(y����ybl�v4K�,v��c�.
,��xBY�Q\�I�,ތ�VXS�����e��(��S�K����{�M��	��"OZ�8B�O3�@B#Ֆ[�$"O��o1��0�`�*pH�2"O̜�&k�9��xh��	�`�ؑ"O��x����]t�h�FۉIŲL �"O��b�F�L0��%�� �䘧"O~0!���xL���O/����"Oܙx��K���=h��ݖ�bb!"Ot�c�l�E�|����{�H�f"OހPd�����1����6"O�܂6j��n�Q˘��t���"O*��TG�Wp�X;Tʆ��r'"O��ѽ+d�A���e�
�X�"Od�"ת�
:`��A���N�0_�(���5���Y��J�'�(��n1Y�C�	-ao&l���>;<�;A	�7[t�C�I�}��<�u��4s�AB�C	�jUhC�I�%�$a�Z�u�Z�f���FC�ɏN�a�jZ�u��Q�j��1� �O�⟈F�D��J�8���B�x���{�@��y��[�	�@�֏l}N�Z���y�#y[�$޽e����V�[,��>��O�i*��"so~H3L��=�$��"O
 pJ� � c�*C�W�`%�$"O|���BJ'S�6����A�.�0�"Ol���/e��qwd�O�I�"O�Ě��8y���S�W����g"OP(I��|.y����/ ��`��d#LOr��1�F�xt"����>��p��"O��ujB�"ϔEX��\Ze�P"OČJQF\�'�����W����"OjdԅF�8�ź$i�8yN�Qa"O�����U�>]�Q�"H�I�#"O�x��������M_�vA�0	��' �D�O�<�BT�jŒ�#�1_U!�� h
�zJ�#��т'�N�;e�'�ў�>��DlS�/����� S(X��Aǃ5D��#�یK���!'�5XV4p贪 D��1��*�^�#�oR>�LC�)D��8��
,~�y'g[W��iR�C&D�������"� F`��Xqb"D�4C��	 �A" X�aꮉ�!d ����2擘r˶��O�uxP-��m�3OH@C�	:�������iW�ߑB��C�!>xH ���	�5��;&( 9�B�	�66$iBrf	����rС"3ӼC�I#[4��j���f��'O!"UtB�K|�I�Z�bv�ى�D��8B�I:{ڀ5�cQ��$|8VLC�'�0B䉩�(Tc���l��IfJ�12�B�I4ψ��rT/ml��(�̂D�B�I��^���)_�F�]���ͺJ�B䉞A�`���#c���
��(�B�)� �e�F�4"��P�k��W��!"O�hC��^*`u��L�@ސ
�"Ov��T
�B����Î%!�y�Z����I�' �aç�}���#n��7�H��d�O��*Q��aǏ�G/2��3���征��'ݤ����ub��8�k� �YI�'��qS6���S|zٰD�B,t ���'%�*�M�î�2��ð]�(
�'�v�+�%P�e<�P؀m��V+����''t$��N!g� @%�@V��q,O��D1�)ʧ	o�]���%!��9��.�$��ȓn�`���T�t�,�9`��%�ȓF�����U3��d��S�Ą�?G��Sc.ïKC ����D5\b�ȓ(Fv�C�E�q~0�0���H�ʵ��/y�Ѣ"�E1 �0����^�E
6E���b���˱>�<0�v��QT����Xp���,�y�Sy�޹�ȓz�|`�5埋z�θ9��G|}���8��L�/ie�!+D�N c�!�ȓt�xg������"�H�.F��ȓRD!�p`�9> Ⱥ�#T;\�q�ȓRK��2�O�m�xe6T�E�ȓgm$M*�(ߝ|\HK� �3�@$����x�u���<��5ȇ��r��C�ɼ���"dF�>�XI�E퓭7|�B�I e{ʝ;@�1E�0�(��75��B�I�=�v4c��CI��ٳϝ�hPNC�I2d�>a&�\�Ay���F��C��'LFԽ�aOS#\G4	�M�1	?�B�I�F� ��P${�d���%aG:C�I�$M��X��U��5�DwC�0X���jҁ("2�u�c��x�NC�$s���c�'��4�v�9��M; �.C�C��/Q~��Q�o�y�.C��	M:Tkqń�:�`���JE��B�	7	;^�y���^a��W�1��C�	�3���A���1c��s3dT�FY~��0?�!�пv��5�D�A��4B7h�ox���'�b�S�$�f��Mi�G�(EvZ}R�'���5�˘ .�%�`�P;
�.r�'f�I�`��'��\�С-	Z���':�P���3<�`(U�Vl��0�'��)g]58Z��a�@4yc�= 	�'֘�J�⟀C���i&��q��H>ɏ�����|Ub���7Q̸� I�<��yB�	�sN�4�u�]�$�m�VF��,��C�I�
 6����?L$F�+6N@�=/nC�	�;N��0K�7�<m��.�'>C��
��д �?)�1��	�
C��M. �r�3�٠h�<(��B��d�f����	�~(�x�V�f.�ʓ�hOQ>%�q�Ѫ@:�0��kKl�	��/�<�ߓ�y"#�)_jТ�	R/X�^0�%����yBD�/�ay���-Q��	Z Aِ�y�Aܫv��E��dΕA們È��yR���A��+���<���� ��y�bփ,N��eR6ybQBw�E1�yb(2�N]ha�^�E�^�!w�A7��'�ў�Oh���fB���s�g J́��>��p��CO��-'F�s#�`��"OTljr��S��pզR�J*��j�"OD��A��'��IҷD �i��"OP�ҁB8Y3�tfN?n��)u"O� �Ak�������# ���ͪ1H�"O��↣P�xa!��]�l�#"O�@�Єیi0ꠓ�ʺ)��M��$>�S��<.d�Jde
/��J�I\ W�!�$���-��A+<�N�#�Ƙ5�!��h��a���fd�aht�Zs�!�P�S�1�a��������-�!�䎩;6��s! ˗2����ď�n}!�G:S��9�pn�{_.��fcE�t�!��YN��5��*�qnZ��A�">�!��AlpPQ��*e[�H���;�!��@�OܐQ5ǁ,gU�`�7�L�z�!�3T(�A?l���;iH�!��{B�az��3�K�bܗ!���pu�q�go.>Y��;$ g�!�Dɼw��y��0V;�t{�O0��OF�=��zp%#δ�(x�!P�f��0�"O�T�A��/;�(Q��-w���"Od ��EY0Z��E!�ᐁG�>0�6"O������>a�q+�=5䬹:�"O���	�OUX��J�'� X"O4�U
ξk�f�)T0����"O����m���-���	7er� ��' �ă�&�VL�N�.UJ����Hy���$�(�Q����Ert���S�@�B�	�3@"劐�܆[��B"l�T��C�I1/�0m���� "R4Ik��_5o_�C�I�K��E��' p��Vf
�Z�C�� ��oZL��-q'�:LpC�	1}ҝ	sL��=>B��L_a}C�	����iߒ+�]p��ە`��˓�?Y���i�Z�~�����a���G�2O��婍2m)�]���R�i�8�1"O1��e�,a�����8��U�#"O��X0�٠����m�#N��"O�����1��M!-ɜU�\�r!"OP�+@DӺM4.���@�.o.�"O��8���by��IB�u��jA�'���'/&]@�DHZ� I�J�1:`Й	�'�b�ǁܺ���XפR,x�I�'�����/!P�qbF�^�&F�;�'HD��1�,Jž�֫¬iZ����'���%�gޑs�h�K5����'>��B�O� !��$jM�K(-J�'KpA��D�#�$u:a
H+
�z�'Yf�y��I�2a������tLz
�'#�q�"�(�\qG�"}�x�`
�'��(t��J�xi�)��vЈ��'��ܘ�,����d�6xE�؁�'���[DT`�f��R��% na��'9�4��bυZ�,4��%!|!��'�T|�@���g	$�s��<G��-�
�'��r񅈣&N�V�tHes#-D���U�� A��YD�&jz
�@�+D���0 �,$��\;���;�*%jf�;D����z�>(h���)����8D�T�T����Pf��)c�j��7D��p�!��ubV��w��yy�|��.9ړ�0|r� ,ʔQ%H=!��E�j�<!`Β��p��l\��9��d�<)��F�b�Zك3f�31[��4Nw�C� �rr��o�T!N��B�I61��Uě���!+�~�B�ɴi��!9�F�d��##��;�LB�)� d=�����J'bH�dOG84'x`qP��N�4�g+���'�G�zH� $�����2(��藙E� ,2t�ݭ) QP�"O�E�F�`:�R��ϙ02�"O~�It��}IL����d�"��t"OPD�D��tF����^!tV� ��"O�ٲe����D�̹J&�ݱ'�'���A�����bL�RĆQ�@ؠN.hC�	(x�m@/X�w	Pm�t��p�ZC�ɖ	1��I��� A�u��	m�&C䉢X�4u:�L	A��t���V:s'C䉧�|���!u�`#�1bpC�	a�c��;�(��tc�~&��hOQ>� �$�S��&K�&��8��*>D�\�5B��&����O�v9[�>D� �$�D$�Ғ��
�i3�#<��0|R�΋A�@�PdA����8�w��m�<qV�ǽik�!�!
Q4l�ZH�u�<�bF\�|޼9+`N29:�`�B�[�<�G�A� �R����Ip�KY�<y�'��8k��	C��`�BAĢ�y�<��bP�)����bH'������L�<�K�H(ЌD���h�
��R�<�p��V�SWH��)�p�!#�P�<��m͋O�����e�4�6Ab��w�<����t�P �FeP�@p��!�Bt�<�����-�E���/����DFsy��)�'-�PP	���>>��c�s¤��ȓdx�` ͟;t{0HK�JB.5~�(���`Ł�j�qE��RA���i6��|��&�M�`H��F@�2��9�ȓPD�	p�L��2(`(��t\�d��/a�	�JB�"�v���,S'|�-��i�p3-٭8'�i�Ti�#+5���#�JD�(I� �1q�a��<��|��VL	�.�,���أ� �L�&���	�<Q�^�V�H[��Z	;�H:�G��<1���6zf�����'�А)clU�<�'�?l�4aRb%� I���6 �b�<�7�,*�� o�:HX\�*'�R\�<w
͊`���H�ϸ6:�g�Y����<���ipˁc�0?���@`�W�<I�%	A�d|Y7e*BU\����QS�<��ӇIбh�kF�Rˬ0�d$[f�<	S�Q��\��k��v����KAGy2�)�'1����bZ� t7��1Rr	��G&L �� I�I�l� ���`~���L�<P�i�-t2���A�2|�Y�?�,Ox"~���72(\A2G[�}���r�j�E�<Y��5O�n��v�S��
t�G�[�<i5�_�YH  8u�ޜU�܊�!_b�<���:-q�)�����8 X�j��^_�<QCK^6Q���`�S�|�:��a�<�� [?��;��6v�R�%R�<f[z��!�S#AO&.�:�ON�<Y�P<?�:G	�!���c�WB�<�C���!E�1[tL<I�t��2�NH�<�uhر3�ty	#ą�\q�L�p" F�<��D��!Px�&ʂ-�JkB�Wj�'�a��F�Zx���f)�dڠQ�K
��y�-ҵg�F�+��F�+H�P�
B��y��\62H$�!��OM�8�c�U���+�O�\@�D�5<tL&�V. R���"O"8[�)pa>a��S
i��!P�"O� ���$?=
t���	��"O�(S0�Q�u����O*e�x)��'e��b�)�	�4p�mZ6WX�|�d��
�����'���0�H�J�6ჹg���	�'_���ǡ �/�@,	�G��w.�@�	�'l�*�O_�K�P�!e!��j���		�'��y�R��^b ����jx&p��'F���;��q�3kZ)h2���'���3�K�i�@�s+��g��,�N>1����2xD��p�iG�wq�B$ƒ�0�!���2W�Z �bO�X�,�$E 8�!�D7���`Á�r/�u:���{��[�<%�"~���H�8���%�N��a.���y򭄜�,� ꉪU�n�p�1�yr��J�Pn%=C�aj��_��y�&Q�k=��'.�C��qV�����hOq�����)E<WHB�E-ͅ�l51�"O�(QQ�]'���,���:��"OV	X��L�q�tP��)��q��<�"O���&%P�d�V�3��9q�"Or����v��qٳ����,y%"ObpyֈQ�	���x@CҘ�P�	"O���'OJ�,�.y���Xl�Lx�"O����Р.�Z�Ө�$�~���"O��@Ƀ�tp2���I�P����`"OPa���ϩ�Zt�EIԽ|�*g"O,Hpt	��R���*���8*��%ZB"O�qs��c1��ɐ�*x�Υ"$"O�c0��7s��p��\E!.tjr"O$%�PdI���t��'�4#����'!�DJ�~� i����F`h�C��� !���'�r̓�$�M,\�x�N�4!�d�9?�HDKGØ=)PЪv��h�!�䌏1#��BB�"f�����e�!��R������{�r ���*J�!�dڹK�ȁ	��2/� ��P��-!!!��17�E9#l��[�
��!O�m!�$I{j�%���"|�Q���OR!�$D�P��m�p�J����#
�'y2�r5AD-B�j����Ӛ	�5�	�'��H0�������@>	�	�'�Z@�}�y@r��$Τ�	�';,(�ס�t꠪ D�t�R�RJ>i���i�C-���M CJ~H#��>!�D�7V��#'��
Q>�=!$`�>,!�!K�x��/ґA����m�!���z��௓r�LL��,� ��R8O��;��*
3�ѐw�՝9����"O|\��ۗ������(PE�6"O$@���>[(\��+�9*q"O���l��@��	��P\�L�i�"O�� �݊$�eS #�
8Ɲ�P"Ob��"�[�~��#��^p��"O����2Js�e�s"�:9(��'u�����1 ������D��&�� 1ړ�0<i�E���a�0
ʄ�K�g�<��W�8��|B����Z�b"(�y�<��j�`��&��E��Nr�<�S-x�Ӓ�6 ��U2@��p�<�%�F2���c&hY�P���Y���k�<��R1��q�%B�����d�O�<�V�4��0(�"XP}�vG H�<��!�v)"p{!��+*X!���G�<����
YQ�%h�L_�n�`��I@�<� ��7a՘�<��E��9)������'LO���[9%�p��oU�QBёd"O�5�')�:jV=	�Q�\�d�G"O�TCI�.	���cb���'^�I",�ش�LU�L=��dg�ej(�O<���P�-r�#l))*�cb��d�!�$�-8J�Q�f�(�iaw�i�!������&Q&�v|��'�*��O���$П9IC�⟨<��c�ǫ�!�1u,�}Z1���4G4#�!��-,�h�q�G�s�nX���R�!���,Q������*�rp�"j�2�)�(�V���G\�z����4l�P9D���'��ѹ��$PM=b�'�=�v��'-Π�s��?�T�vD� >�%��'��qq��.E�DH�ꏿ9{ZA�'�L�B��\�DxGă*d,���'���2��T�@���@̾)�d��'�DyZ�$J/ y��	�%Ֆ���D=�X���o��a{.�"�JLP,aj�"Oj=K�)�%5Z�]ۦ��=*6��"O�(�ևX��l�a	V�	�$���'�ў"~R+��.<���B�?? ��N[��y".�33n�<��ɞ3e$�dV�yb���+c6�)��"(�``�櫛��y2�O6��J�Ƅ���P�!��y"B������׊Էn�e5���y��Nf�[�;�=�AG��y�@B���(��%��u���Z:�yr�Ĥh ݺ���Ii��`��y�C��E�@,�W���d��y�$J
IƘ�D�߰L	^��p'®�yB��e�
��%�U�n�2T�q� �y��r������nE��ҷ�ּ�yr�C�Yn@,�D耺l |�X����y�	;�`�i�Ȋbd�|ȄHZ�Py��O� ����F�"�6�9�E�z�<�4��.n�p�'���C��5�mw�<�q��|dV��ef��c�(9ҁ@q�<�V7w�B�
萪S��8�C�w��l���O$P�+U�Tcz��"?�✚�'hd8s6d�"�4�����-���c�'Ox9C��j\�\�V��PǨh��'�0��q*��,@ƨ�Pj�6�Ѫ�'���p�F�P��} ń6�9A�'̘���T�T�E��E\�{�8
�'C��ML�2�9��#E"�J�����*��Ӏ0� abU*ٞC蘭R�ŇF�4Ćȓ:��d��MZ�r���wI��4��QpX�0�̓Z�LQ �/0��ȓ*�H��'҄;���[��6`���fm�$�e@ԏXP�|�f�ގz�(�ȓ �Z�+$f�w�T���V��܆ȓD�r�.i�d�&�J�KW1D����H]�It�B�Z��3D��Q���G�飐�Q�S�X��q'r�L��/&�S�O�]9�)���� Ù�H�P��'vj� Q�Ϙ��l1	
Ht$Uq�'�n��2�аAXx5ʓ�G}�P�	�';0"3�;/s��aT�T-Bo
�'����*��ּHd�0,��{
�'�x�8�/���q��M	7:�p
�'��h��S8X��`����8w�GR�4F{����Wl�5Ӵ�Ƶ �*�聦Yw!�� �XA2Ԍ&��bңP�V|�"s"O���dC
�X��̢c�	#h����'��Ƞ6�_�ı����/5���'���s�Kӊe���!�V�:}��'6��I�8�T���D�	I|A�
�'���E�L�Lʌ<�7�Ј|��a�
�'p���P �rCF-��E]3*S�(;�'� 4(�&݋�p51��2*9����')"���oôtN�VZ�mR��i0�!D���Añ5���q�ǽ�D�1� D��Ri6S#2�P0	�J�(eK��<�
�r}�8j�����Ʀ�$� 	�'�x��V �K&\|�G��*E7��!�'� � �K�#4Y^�Q��ҟEŶ k�'&}c!��$����G��54�x�'�����F�+q>�+��d���'�p��`�9h��MF`��	@�'vhD�Pc�/c��+�ٮR��#�'�,����5�@��EG�+ZJ���'y,#�!٨�м�U��U��!��'�4�B��;#�(��Ǘ�E��,Z�'�:-�rHHy-�� 7�
"@H�	�'���B��Opߨ(�j�MN�H
�'���BG���Of=��MU\�ؔ��'ZN K�AG�d#R� <? 5��'vr��E�/ZM�)�AS�8��0��'l�� $ �&,�b�B�֣-��	�
�'�|�s�e´H�P�Y�ǟ� �
�'�DaG,Ϲa*��J���I�a
�'I���c��&p��n  ��9�"O����6vvB�ZN�q˪MӅ"O�r����6��ڒΝ�p `r"O8�:p!S�;�#3@����{�"O �J���B�p�S�ψd�ZX�"O��rϵ~�ѧgՐ�:����'�ў"~���[���l��L ��!����y��U���rGHX!�'���y� S�L�P"f�-/Q�-b�^$�y� �mh��n�~�9�wk��y����ܢB��ٮ)עQ4�y2/�y�>)�c՜}npS]����It~2�^� ��J�e��-�y�kǦ�� �C�A�%�t�K��yR��A��-A�cY�>����y�)_��X�����2�ʓ��fC��U5i�C�W�Z�DKY�lC��2[s�����d)��T�
�<C��C4E��G��d["E�c����,C䉬Y�`I3#�KKPD"�ʐg��B�	�c�Z��G���8�$1�B��Tۜ�� L�H� Q"'
P�D�pC�	�+=I��S.� � q��Dg�B�I6v���S�7A씝x��(}�TB䉱('��x�E/<$�%ғDM��`B�I%>��@��� ���Z'�+I�B�I�-��M�����RWe��`��B�ɳo,z�1���Y���k�W�-�XB�I�vTҥbU�{��h�!�zRB䉀{���gc�"L�d�+D->B�I1o�d\!���{v��CC�X�""B�W��PӔAN9�"h:DB�ɩZp���ʀe^�u�&@_�(B�	��"Xp���<w���"�^�gY�B�	%1�8M�!��n5`��7��p�BB�)� �����x@�PB�i߬/춄8C"O��e�^�Zx��g�
}Ш"O0�#��Ŀ܊P��=hZYA2"O�АIU3cی��D4OcLUB'�'�ў"~���®j�<m���J���gV��y�J%	xA1�ė�H���T�y�G"��굨ɝE��I��i�&�yR��'w�i�੝�N���"2�D��y��Jqo^T�JCL�!9�$��y���� B���&��5�f�1-��y2��NV��[(c��� ��1�y� ��O��LS��F���"����y��Բ>�K��@���b�\��ȓB�N����#n	�)��d�o�B��O!����T0i�2�Y���15�4�ȓRMN��Pl8	�4iY�Uݪ��ȓlP�!���-M	����-\��g��t&Ϙ�F>�T��HP��ȓkx=E+�-�~I���<!fE��|3ndh�TG�@��S5�t؄ȓ#4X��U�׈7��=p�@Y=l�湄������ӳm�Y��hN%>e =��B�f�`�+H7\5"��I")�Y�ȓeg�
��?Oni*��B*ȴ�ȓY�*u�A��<�ii�ENJ��I��JO
`*"ŋ����Ke��*� A�ȓT�ċw��44���"'jE�؆�#�z��D�3F�D=�O��	����ȓǞY�!�++��M����(-8T��U���`� |\T׫V��V����YY��OI�QHgkD�W�ԅ�3xb�i� ɷNxX���ᝒtE����Kz�����_�K�9�\��*+D�LP&�B�_����s��3}j�	�)<D�$A7��k��e���|� 0�ab:D��r�� oӞ�jS�߲�؅�ǀ2D��֥�/\��q���K0A&D��Q�#	�(\Tx���	X&n�C�"D�H#ޒ1H�a��A�S(8�j�J3D���h��
�3�gV�}Z��=D���p��d��@�D��R���a��'D�bG!ӭ3�����`>�E��;D�ة�m�`i�88T��m� ;sB8D���٤M�"��3�ʎ-�d@��3D�xY���&����H�!+Yzq9��+D��+gG40H�@�$D�
֌���.<D��k�D��ġ[�D�f<衡O;D���珅(	�X�;p!��fT�܃�M:D�0 ���4�j�RW�]�?���2��;D��q��Γ6����"�Yr�ٰ�9D����1Tw��q�
 �%�d�4D�,0dIP
u�6��v](�Fܳ��1D��1BK�.(ޭ���Z$7�V1��B.D�d!���
�~P���+@t�=�B*D�T�rD�#%��=�a�fo��J(D���')Y)-¤��C�_5-�p����'D����C��+NBr􅝋[�d�&�;D�\�֫��#&c1�;Oz�e;D��)C���p$(IH�����5��N8D�t���t(�a׏Q��J�5D�[��_�gt�3�˟�n&��8D� ې�W���h�aEعO2$��(6D���.�	���H��I �3�?D���X*����"ȹ}4�)��a=D�� R�eAO�yi�Ũ�bҬu����"O�q�%�e����\�N��p"O�)!���w�qkV�ön&p2�"OȰQB�p`�A%i�\��hP"O��cnԓ9~�m��3���I "O	K�L������+�����"Oڙ�d��Z.���F =�֜�"O�s���N�V�K5 �HkD"O�ՂU�W�&�MYc#Fv�R��"O���C_�X�׀T)(�"O ���B�1M�x�b��.�0""O6T	 ��`q�1��M��6"O�m��,Yk�����*}�]��"Od<
�D�A�����"��X"�"O81�'�8FĊ�f� i��H "OR���蜭���þ! l�"O|�Hq�5]�A3'�ǒ�2��""Ox��K��, ^,�A���u�vU��"OH����N7E�fQz�t}�a��"O�%��
݀o����1ʞ(a�4}�S"OJ@z1M�Z�����&j���rs"O��hP	ƎV�b̪aH!:9J��"Oy�A�Y�l�E)T�Q��ȈQ"Ox�صٚn�q�	
�+�&�9�"O�e��./���QHL�h�t9��"O����0aPh@�HD0��"OЅ[ �ƨe&HC��
vB28#"O��scnN4_^��X1�G�tZ6|�"O��h��	u��h��eQiZ4�Ȑ"O~��a��xo�����ZnY���"O�!��Z� <��䑩8X��6"O�(���<�V��@V�-9��@�"OH@C � �@��%��oC�TNl��"O�Ũ�k�m�m�T�� xIx)�"O�iI2`�hZ��!C���LGj��#"O���ժk����d߆�9E"O��k�X
��3v�C�(t@E"OT� uk�*�T�1аcl�ȃ"ORE�c�H=L�x�#�e�{c��g"O���v��R� cUE�#�j@j�"O.ų�Ō�^E�����v�t�"O��:��ݫQ���U�۬U��"O��3���`����G,~�.,0c"O�kcC5���Ï	��1��"Ob�@�ꌃ)�reI�v��t�"Oำ�X�lC�����)@�r@"O !e���w�^)�B፟c�Yr�"O�����
H"(Q��2cD�+d"O,�a���B���,p��X&2L!�d�%'3:�)�Ⱦ�x��fm�;?!��U�Ai�u딮�y=��8s��_&!�䜚X\��A��]J2���*�$.�!�D]��9�[� �-�@*��j�!���0=B�A�핋U�dxo�. �!�҃g��q��D�P�mS���'�!��V���P��"�$vUk��B�G�!�^v6��6��> 1�(���!�H02$�9�3�Sd[�`�Pȋ	�!�d� ��s��J� $�R��%�!�$�4sd�%�!��%ɾu���	�!�ȿ`��	R�lV�,(Rɠ�լ�!��Y�/���I��G�7T��L��b�!�N�z���Ϋ;-
]Y�+��k�!�$�/�������C:�$ ���A�!�� Ě��3u������F���Z"OT�a�h�B"	��]���7"O$�S❕�R���-dse��"O������813R3R��Un�ac"O����$��4��P���(:�P�W"O�ig�1kLxz�*̕
��c"O�d#6�:���@H�.n��B4"O�5��MӮ^T4Y�F�6�>(p"O�X��]�ql�疶�0��w"OJY�BdƤ!��H6F͜GM84s�"Oy;���'tF �b�c�	OD��@#"O�yCf���n�R�V1TJ��"O �jR��+���3�fH�
&�"u"OM��љ<�v�Q�FΩ�m%"O�A7&��؄��юd��i+@"OFdy�IL�Y�0p�U7g,��"Oʬ����E+P���╊;��)D"O�gMY��� B�Fu�H��"O|�Q�C���+��^�H8���W"O��Ao�-D}�����~�a�"O>A+e@E�me��:�`T�'��1(�"O�e�R��Q���a�ƳzM�%Z�"O�I�Y�n��x�P�P3n\I�S"O�H����,�>�:T)��M|���"O�a�!��z��ŃvG�W|��7"O8�Hl�3�A{$!ךF�8)�"OY
r��&$\P`F�Y�x@s�"O����`�]��Dź"�T�"On�딆C�qjD���&�d���"OhكҍɱH��Z���,�[�"O��
q�'d��#Μ)���"O��Y5E�p�M��_?�t�x"O�0�Ł�5��]�Q���z�"O�Tc���gJ�
�+�x�1A"O�,7���o�Jƍ��\����"O�`QpJ�����q�¢~m��#@"O�ى cYzZđ�U��VTM �"O�d)r��C�^p��ĬI��n���D{���?*���R�BR����ף��K!�DͿH� ���̞Qd������=X�O��=��
$�g�_�W��AdD�����1"One��
_a����c�%��ݩT��4|OT<���o�漘Lå�������<Ey���T�x���*F��ΕArՎ �"��q�0D�$�$Y�\ѡЬH\f �y��.�0�d��(O���C�`��tk�G����	�A��y�l9M4i"`@ ���{�l����&�S�O��!ˇe[���@�"�� z�m�
ϓ�O�E�r"I�5��8���
�0�7"O���b	�BO��p��S�@,Z@�|�)��>����#�V�ZP��"A%[�C䉏p%j����D.�������+Jx�	]�'��SG�'e8D9��螵K���!����_�2������p��^?%�(�U�-I��T��o?��O8T���O�TÆ��a��"��P�FS��Z�"OZ�)e�#"���T ���|`�1V�\����V�x1#ŬX�F��&��C��?���D�uk����Jd�����c�<��cؔK1+�J�DF �U�״��Od#~:��*w�X񘇉	?��l���Fn�'�D�G�d���\�~\a���B�h	���&�y򤖔X��\����0w)B)بO��h�O۔�b�L)�L���#k��"�'�F0q���[d��׫�6\
���*�g�? <��_�me\��Bό� �Br�"O�J@,b$BdٓNL��M�D"Oؘ9MS�7i�P�͘h�4�S"O� 9�&V��c'̄���!�"O,xqC/�x��bJ� �^�("O�ٱ4I��-�|t9Di߈%���"O�Y)��S`�Y��E�V}�h{�"O��Q���{؆5
�eȤ*M�e��"O��1JU���P��	�5f7,0��"O��$璂^B|k댹��W"O�p��o��u��jN�(^�q3"O.Ys�B����U���MT���;"O��§�ܡ!�lR�"G2Ky^�#a"O�l�v�R�:1���Ͱwx�˶�'��$�H+�M��Z���q`��	9T�!�d���C�ж�:-(���.i!�d�2��,�����N�$�I!���:P!�dD7ȣ#�{�`+�J��pB!�$�35�p�ؕo/}�4�rɆ�
!��+'Uޕ3��ՠ"x���P�PO�1Ol���ѣF-:��MiTr����!�Q��h�ת��)��I��(;.�!��Bv�(���@%n�0Q�?m^��m{�O��bd���`+4q���b�ȩ
�'ъ���*)+�`0rN9ˀ�l*�Iz؞(!���(It�����ʁTrL��B+,Ob��n�����kO�}eh���-P#�B䉸/*)R�$�*�";Gk\�Z�pB�	v��pv��,[��"�N�pB�6x���K��>.W��jdd��r�&B�ɬ}w�m��U�P��}ä�]5cG&B�:<�[�^���:���P��C�I�mrFQY3J�<S��8r�C�	�Q� 0Aœa��xBu���"�MI>)�P!��#�d�*2�6�R�$�
~�̄�z���;*�65����dGg���ȓK�A�El¿V�<I���C�f̼��>�O�"���O���!hW�'��T�Į���	��'hҰ��Z21�j��`�R(zJ괈ծ�|?َ��S�o��:B @8wf���@�19����L���'�΄+�ę�S��f

�thN�h �'�ޜ�F��PA����"��!x�{�)�	\�'��aP��d�0�b���(�!򤈤 6v}����4`��"DI�"N0�D=ʓ96�}Z��::L�\��� "@��QXglF�<� �R�����T &���{�fP\}�"5�O0$��(R[&�B���R@P\�T�'P�Q����?�Ձ��`�Z�B�
������<X-hGy���'6L��)�z���C�c~���Ó�hOL���Հxl�|�2������OX����;���#�l̥tm���*n@����>9�E0?q�	�71� d��� ����"K�<���6?�d���˟�w��t�C�K�<Y7HFC�΍8�cѦ(�D%I�iI�<Ia�Q��X����)�b�s��ۦ����)��!!�Ȗy5��ǎ�.i?H4 ф+D�|��
�+S]2cJ[�j���<�Od�j̴RӃ��j��S�OŘ$�����ɀ1a�ɶ-?`���
L�%3�B˱$@�C�	&|���$K�kj�r�)F�x�^C�	"_�� 	S��88�j4X֩o�vC�I򟸈"HǾ�f��G�āEF2��ӆ���E{���M�W��)Z%��&@8�I)�!�&M줵��l��*U�A��]r!�� :�q�bפg�R ��Q�#\���'���T��R�#�� �!I
.C�I-�
�0�V}K�񻠬E	1b�=�
�']��,��(L>R���{W�\Wd�ȓg0ؽ���*ж4;��(�� l�"��'& "}�'���9���;�~�a���;vҔట'Wў"~�c��TX~ ��@F�ۨ8"�[w�<��,B_�Vm�b�V-��9�"-u8�&�d+S*@�b���3dӋ)Y2T{wA,D�`�Q �j��LB�.RR��iC@,D�4+3�ٚQj�}����1��Ы�,�OvO��SR�iO��iŏpʰ;U"OXQ��_���Y�_O 2���|�'��$:�'���@�����J�>)��-�J�c�>��zW��}�h�')ў"}"���1u�U��
�N�|�`�Np�<�e�5i���� ?��	p�Nn�<����o�VܡP�M'o����@��h�<�pn�	
0� b�"�@l3d$'T���4�u��T�Eg	�X�1��hO�S06*V���?Дt��*��K�'��[ ����!�Q & u�'n�4�O8�,x�B��q~~ͱ3FC&yШP�I�O�<ѓ	M�8�v���!�#�:�*vj��<	�j�A��(�r���Ǌ-O���uHܧ3��q���',�^���#��+d#0l�!)�14��U�ȓ#>\1Kf��!~af`sN��G���'�ў"}�G=Wq�$��._J�Mɦ��p�<t��gu&�sf��Vx����h�C�I}�'�>�a�(Z�C-@�9e��R��x��?D�D)�*ŠJ�m`"n۔M��E�7.<�	�^�Q�b>�"@�w���Ҵ#��'�ĥ��:LO�㟄��₩�� �q��bV�h�"�@��~��L<�倞1�hz��I1��a9wM�r�<qQI؄KΤdjVȺ�Ԅ�5�p�<Yd�:�&�f��H�B���I�n�<y���1z���p�"ʈ ���0��m�<IF�S
vi*u�r��b�̽2�@�Q�<q1�ݾH��уU �&���� L�<I�jFs>�1s�P�6�ۓ瘅��x(���h�'&O"4XDEҮ�y��[2��^�Nό��c���yrG��v�x��҄åJ�����˴�yB�0x5� ""Á�r\�IÃ܈�y2`�?9��laU��|�{ϙ.�y��	���T'ֹ���֋�y�ę}����͟
�l�JL>�y� Q�C��aR��ۑFb�c��y���j��(��N<�J�j[�y"O�qf౒�d27�$G�%�yB�I[] ��N�,ϔ)am'�yr(^,p����
�(\�a��y�cY�=h�U9����x�gC���yҡοhX�ق��e��T"����y�;G�z#�lQĄ���dE#�y��̗h����f��FX��*�䅳�y�L�(�����g5����N�y�j��$&���u�L�+��;t�Q��y�n�|�Pq�篝�(\F��`i��y2b
O3H��)n���`"D��yB,͉ba���}�ɛD	��y�AȆ5�a����q⣦��y���g:t�g��zLa��dǤ�yc�:+�\)��l1�=��-G6�y
� �ujP�6^Z�y�3�@<&��`B�"O�)a�I%�riY�kN8
��"O6ha	@�<b�����ЇK�VpR�"O��2!� �!c�s��U�!"O ���2O�|{��#[e��r"O*�ѐ�EiCDd��Ȝ�cnd w"O�xt��o�͋��ז;X e�E"O(-J��?{jI@Ro\7A����"O��P��&���
v�ttb"O����Y8	��ɛӫ�<-���"O�1��ʎ��pd�K7C��
�"O���U
RR�9�({� �6"O�	ɠ#�N���`����q2"O��3�Ɩ�3D�${��ؑ[��R"ON ����kO�H�c�Q?"�	G"Oi�7��!��릭�w��"Ofl�4BC�p�@A�!y
�X�R"Oh�"�c/|��"cd^8�����"OH�In����Ǧ2O�Rt�"OȸHt�ˬ2h��"Ն�y/!�"O�4����6 �P��$�PXpx"O�l�b��|Є;v\L��"O�� �2Ӻ��fhD<����"O��ْĈ�/����;# (��"O>�1�EOUd`�r#Æ9]*��P"O d���2,�K���=)d��"O !��k�*td�c�:�����"O�q��1>U�0z@�Z�J��s"O��7��mK̼�P/B=.��)Y�"O��X`&̏)��Q����y�.ȡ�"OP�%�("b�mrW�O�&쫴"O<�2��j�x�bRǂ�A��=2�"O"X�7��*9�\�����4]��"O��9�F:~�`��/�B)��"O
H���R����!B��!��5K�"O�iz���6ڰ�iaCC+1,b��B"OJ�x2m��Mk�	�r��6�B@�"O�%i��5����E���:���pE"O(�$	��?Te��Ըs��A�"OT(��k�zz�h�S�E�b웶"O��Ct�+F~�<�u)_5Ii&٠s"O|D�ACĎ_�5	b-{A��3�"Oz�9bB��Au�4[�-��^L	�`"O��p�ٹ`�8ɹ���MLp�p�"O�ܪU�@��Ȫd�قD+�X�"Oщ�n^�#z,B$bW�N"88��"O���ݣ4N,]R����JuJ!"Ov��5M�g`j}f�Q�(;�"Oܼj��k澰�t��GXT-�"Ol��҂J'0�U��N#5|N`H "O����m,<bJl��G�vmRp�"OةT�ğ<���!��7G���"OpDb �Kc��8�ɉE�R"O(��c�̪3������@<E07"O�2�#�!r"��R�@�.14�a�6�'���X��[41��v�Z)-�`|zbֽ~��L�t��y�,öp=��ȵ�E���1�M���O�RGLo�rTÉ�)��Cд�����2W�u:6��I�!�]�]���X�+ܮLI���f�0-�ܱ�5�V���ڄT��F��'���c���&K�"H�4�5�:Ea�'7�@�.�ɚ��G�8 ���*��8A��L2td�ӓ{i�qKW#C�qTr-�&H�jT���I�(f�Tˆ��~n�yKK����p�1��(S�L�<�uG-��zw�n���²@�@��P]�r�kO\&b�[��� t2��T�9��4���� ��TIt"On���$�4�j�0��;Qr�M��*E
�!��׏Q2�Iw��~���! P����:��:q,Z��y��J2�((��9���@��>�?1�Hg
���
@
�0=��h �a�ep���F89uE����=@!
PP:t�Q�d�0�G�m����͛M��4	�'w��V�M&W����hB�M^�Pz���KH*�X+�-@�(������	::�q##�~� �0T"O��3e���r~}Bv N42����]<Rdn@lV/��S��?����J�X���\�I��T����r�<�#�6�D�X��ۏ3���*��q�<)�LG>y>�HuEU�$��*d�Sh�<ypi3ވ�`#Sb����r�i�<�c�I�Q��Di��ddra��)H�<��T�4�%IG�U!Ϡa(e�D?�Pl�:�㞢}���)���3$��$��(��g�B�<9��N l`�)`�+�)�`i�&�y~�FW%5WN5���'��Q��L.��yS�*�.�ա��h87g�,z�r�i�@�>�}@�/� k�8R���Ɛx�*��W���HF�_�Ԥ�2�ʻ�O$\Y�m��p����G�'RЕ�i�+~:p�
!���k���f���h���;gb�����\�`�rFK		,��`� Ih�$4�g?QSCn�����	�Ps�d����]�<)BE�g�m��I��ؓmޟ,YfMQ�$��P$M?�ay��z����rA�!��jѮ��=" ������EE��y�\̢�b�'?$�#bC��P쬳Ќ%$�����O<�|�bB�[�~A����,�I<���1�KZ�rT������O8m��G�=b���G�Nm!��Ӎi8 �)7.��ԠrG^�bz4��F�Q�wt^����+u�q(�����M�I�Wy��w@S�.�P��U�����؞����>'VХ��A�mcܹ�ci"H���S�O�I�fF��<1Û����H�i��
��4����Q�'1�mkp.��G�R����H-�	!&��7�8����W��r�ϔ`�0��:_�8J�%54�����(�w��<��-���)���,E�(�[%EI-J-Ê�I�9d��-��i�%z
�[�!5!�ċ�d������.S��=o�#�cf,�=XR�u�܀�P��~�5�d��V��b����E��a��~�䘳(r�J����Fd�!�@cG�_��(��کQ8 q{&�>b���>\O� ��ڠ\<TY� BT�G��m���I� ��P�:� ѾvW8�R�È}�t��
�.�x3�:~$u�ȓI�$Pg�@3t�^�pf芩~sTU�J ���Ub�1@SH�����'B���d哿-$U���K�`s���C�R?R�C��86`D�F�p��P��KsU3i8t�0P�Ǫ(�E���x�4��OV��aü�&��+Į�2�o���j�L�x؟L ���*5�Y)�Jɢ4��r��ȁ;����a�� ��0Z��,�lZ��>ػR��S�'YX��!�G�g����jE�0��-�N>��*ţ1����(?N�(S��^�P��S�ּ�X���i�����H�T	����-~��H����=X�~dI�^&�H��O���cZ>Z�h�-.��'>^�`Ǎ�-��(KK'F���B�Dv�(��&�r���C��G�y@�/U��B��i<�}�`n�ZI� ���%LR��	������0�>�hB@�#V�u���[H1��a��Ե���tϳ0?<�{��0�x��S<8��԰Do�x~��)}f���
�&�$[�� /!�Ԭ�W��\�4A�i�؅ԟdGyJ�����B�O(���QF$׋���R7�ݳc̉/#��� 3��ň�?�bң%����ħ�	�� Q��Ȉ-%(:�(��Ky^����
`����ͤQ/҈P��ȭt ̱(�>�Փ�M�Om,�*Q�ŀSH|��!���b�^�ӄJ�"-�ph��k����--��= u�֦Z`�\��ޢ9���Biy�d�u&Ͷ�1��>�|����9n�T����*_f�%[�(m8��su.�n�l�������$X�PS��G�xtfqA�-�E"�P��>�¢[d����B3_p��`2ȧd#z (7ꋞ8��O�L�8 �T�?sX��	҃t� ���8/����k��.�"5�''΁-��[�j;>i[���� 2��q���e4-���3�ę�g
>9��fHY���2-��_~�Riȡ=���pa�	��-��U�d�!S�����q��+�<	5|	Cg�3���_��A������S�g�? T���+k���@b�t��ģ"O��V���B���qpaSj p��EAѺ��j"x����x�Ǎ�^�<��B)k��=�0Mҫ�Px�.c�&P8�;4�zvcXp��Y�� ۼ���I�A�����N��UVˤs�(�bN\�%#0	���u\~x�'���K��S)&Q2��A$��8�J!0,l#2B䉡F�,�1��3kRM#�Ěw8r��1�<���U6$A�ѡ�#ʧu<��3��X(� S7<��I"�2/\�B�	&�a{V���� ��mĩ#��9��]�e!��鐯�2�L�j")��&�mG|R����k��hZj�p�⏀հ<1�� վ�x�
��LT���u��5)��P(0�^UK��� ��917(�p�a~b��&43���cb�\���ڙ�ē6�n��ς40�@����cTb�0�l
P��3x3Dy�(���iw��B�In@���6h���n�9q��Y�!��K[!Gl �5'��Ywp���d��8��t̓?������ZO.������N��|��BV��ӧ�{L����T����BGG�<{���gDH;t�Bq� �ϩvq��٣�IiH(�xDCH�:�t�Q`��0�����D�G��I6�N�h���oʵ%⤣��HVRIx���I]�-�c�:Z�����8;8����P�	�\1t)�~�h�4��R��ӚU��H�'�`^B��4g@��B�9DL͎]�(��J�5�y"m�	0*0��R��+^;�5�V��G�L�hcbª,B����_mJ�!����|R�G�V��(i(U�_�^MR�H�xB�G.T�51��-ep�T�d��*9�Mjwّ4f�"��ȗI�"-���'�<,�b^82�9X!�VZj�Ó�ʽ�A� G�4���kV�h��
P�_2ue�1�WX������xBO=5hM@Ӏ5lB��7����@�nԤ,5���B?3b]1 S�4n@�q����3K��*��R�Q��da�'ݺ9�g���
i�a��X�䌑�rI�yo��� f�e��1k0)*�&8�G��]���\�PP I��o�,��ŉ0=v��&�e�����I�o,D���ːU~���B4��,Ǚd�����OD�asP�8�f�V� [X,\�4��7�LD|"��o�����Gٹ����@�����֟g��r������$(��i�����k.F��J�R��f�I�yH��,��#��P!���0?�E��?K����H�'֘�C�e��^���jO��G 
�k��I�7i<9�:(��Z�y�̃�w#��c��C�M`R���o�3ft8���_&���P)*{Ҡ��*J�+���*U�TK�����
�����̮U�FQ��*ѫ)~��'Z�쑊09O�\Iq�S*$\���F��us�)���ip%J���<AN�J& '�t�A�途�-kЫ7a�u���@qpoڱ �b@C`�g�']�i�����mgf�"Rb�<_:Ji�.O���Q
I�s�r�8M�֝�VFL���+�)Ӳ���a�#D.���G�L`G��Z��S
:��DB��z�a~r��Xl�B@��.xX��wB҄A���'^���W�E&�l9��0A��K�E�}�Z`�P8��@���(Ҽ�ȑd �D[�H���'��p���8]�� �M�.N�auf��FQ����Ȧ�h�e��N�Ĝ���>E�ԥ�
?��<1N4mo4�Z��]��0<!�e	ku�asK>��!��w�l�Ó��q���3���(�'���#3�{�g�)*0�3G�;$��7'P5I�2ЧO�,�7�� 긧�O�\\�	�8H���(��Ȋg��X��'��3 !� I?yx�&G=[l`p�'Ɛ���Ii� ��szhm�
�'���/�`��0�@fدu�L�	�'(������5�7�Jd��|�	�'�44�-Űx��j�A�^�R�'��t��c.H��"�u��a	�'v6��a�c6�Ab�ѥi���'�l�Q&��XE!1�Z�t���2�'�HC�	j�N��ЏE4n�=`�'��t���R�]���)�#V�-9�j�'fD��gd�%)[������8��'�z�ˇ�J���y('�Q�h�	�'���&�MK�feP�+�:c�ִ �'�Cb�ƫf�p�;��_&N�$��'F�A�@�eb�l0��:�zxR�'�� ��8z{���ʂ�7�����'A��+d�.!�ȭ�gl��r�s
�'m��X�@/"�,͸6�hͲE#
��� �,r��z��Y��V�<ń��"OF,
�� "6�b8�`˄ 5l��p�"OP�CܖM�hH���G^y�""O ��׻!*��5�E5fR�m��"O�Y �$�Nڸ���(P7$-d"OQ���e��L��"ۿh����"O�ٹӃ�wx�(ƀ�"Qc��t"OH���Ҵ'i�[2�A�%l�8�p"O٪�7R�C���
nL
D�"O|�h���!�� reo݁3+@)�"O��km���V�J஑B�ak"O(�+�h�r��X�C����W"OD��,��h"@!#ǉ
����g"Ox�J�d�
H�<]�t�G-o��4+"OhP��P�	�$��ƫ�i���P"O�B�̜�Cc����L	'�4h��"O�D����)�\(��o�B�YAs"OZ��p�C����U8�"O���¬�n�0}�E�� n��txt"O�|p�o� D�R�Y��=t�!{�"OH �Jع,��a�G�v{�)qw"O���B�\��E  S�x��"OЅj�F�<�5Ѱ�P�oM��h�"O��(aߔ9�� �'C9�L<�"O"KC�k4��@�L��"O��(K�yͪ)��F��S-�R"O`���錜P�"���F�6�^C�"Oh,�Ҁ\`�8-
r%ڠ�V\��"O����2B��nԚ8{��6"O��K���q�8u�K��RR�cg"O@Lم�JD��$]��4IV-Lc�<�6L޵d,�ɢ���5@6I�Y�<y��J1����G�]?�q���M~�<ٖ���U�b�qS��(Sn@��!�{�<����
$.P�1�nj��k���h�<��i�|t���9>��X��E�g�<ɗ���=(U[�N��G��G�`�<�G,T�2�]��'X7$��}��H�<B!��LG��Q���kA�E�c�s�<�n�h�}���v��Nb�<	c.ݭ��Ș��L�}�D���.\�<�GLU�{��za�T�L@JD���S�<��=T!xI2.@�lJ^u�pbp�<�Q�X�b�d��bĞ
0���ee�q�<��\�F �Kg���`W�	i��q�<���$D�"�g$�>d�j�b�PE�<����n�Z\f���
�l�B�<�h�?B4f���Ƙ	5HE�[C�<1A�P�d䃓i�3K���rk�x�<�����y���iU��"L3���$��y�<Vf�;D[*��u+�Rv. ��cw�<�r�J�@Fj�S��]������'HH�<!'�[�u&9p"�6 ��j���O�<Q��,v
�������*"gDC�<�6`Q�|��M� �9�əC�<�c��sN@����� %¸�fv�<$C�+�*41�aT&9�L��^l�<)��ɏz�d �Ŋ�s^~�djF`�<���`Z�*���5�NuhT��u8��*��с"԰}m �u��/��a�X`C�I8u���"C��:�w"͖}I\#<ђ��*r�B��d&��B�����z��v�.�wl`�<�GK�G��,��/*�"�$�
t�XC�	#3�*��'��>��,m՘i�ei/�x�s��(��C�)� ���T��/(Jd��Ȋ'N�dY���'�2��"��4^��`´�'j$$S�H0cQ�A�T�.L�X��	�I`^ĢD�)`*0�̚���3�%^�A���C�y"F�Y#8|[S��&��<HR Z���'K \[ѬW�RlЖᓺF�(TM�OjD�F#@J�LB䉰r��x�a��LrqߦV��l��Z9�tǰ<	���O��Q�E�T.N�(vB�,:���y�"O2X�h��g��1(#E�TA�'�^A9櫜�4�2(r��'���I���#�l�P�#�$a�x�ߓ?�T*VlZ���AE@R��(i\��i���b��k
�'�@!��
�4;3�E��*Rga�dB���N-ĕj�����(�Vx��o�p	\���	_4�aR"O� �qMnr���b�<Bҕ��N�%���f�y�)�矴��#�*}"��
�H�#{x�����,D�T�3{���d$E�/��l���.D��KU��aM�e�K��^	d ���+D���� �#_�"�1ש@�i	FPS�)D�؀�	�0k��6�¡wߌ؈D�$D�� t ["T%`GN�/��Y��n��d �j�;s�qO�>��PH�{�Y��d	�L�2G�%D��Ѣ���q��Q�� v���kÎ"?�"�C�"�3�*��4��N_�¸�hŧX���ԇ�I�c{:��#o�98HL����9%��zO�T6� �zH<I��Xqł�5i�0OU����m\}�'Ҽ����ӳ%�%�e+2��-Q�����9��m
�r|�C�I5���@3m�4Qt�E�@�=�%��a�V���+?��@���h��D��p#�a�%E�*9�SdU;;�!�$W�5�.`���6 ��`c�DYRm��^U�HS��Ƀ1,��Ib��A�7"ƶj!@L2���o�l��D�� �	��JGd��Mz1�֬t���@���Fe\�1�F����x��M7w�R��L�&�v�3ǃ��'`�d "���k亍╅p�'vM:9���$�������H6���KgZ0RG�S;>"n����,f���� sX*��S"�<�D�r6�Q��	=�'���{%�X{-�E���ST�	�7LE����}�eC`�Px ��Yqh�!���G��7 ,M�g�ݝ���C9*��H�'ˠ'�h�Q#�C�J/Q���� �'{�jb�6u6ؙ���9+ �*q�/I0b��'aPFYQ"O0�B���a�tYSl��+Z06�O|�T�J�g�@�H�1Sx��B�7ҧI�rM�᫆8/oF���ήn����~$��M?b\� �g"߲)�,��W��0[܊���ͳ~*���k�n��qO���"_!h���J�������'�x�"���#{�m��A��{E��31��mb[�[����P�T�>����(j�9yqD(В���P8P�Q�x�Ҧ��K`��!mY�N��ciP�)j8��F:U��8a5oE�0�
XS"O��ڵ䐻FI�5zp�:Tx3b�O�%z��P�vܱ�`[~�j�
h�c�O�BM��$K�DC���v (�f@P
�'���蟟Y�<�0Ƈ�(��iŮ_�	�����M�az��J�\W����?)����!��ŝ@�vlB���O�L,�P ���a��
9�L�3�ܼC�D-��m�f7�@R)L�@���ՑI�r=AV�iI.�aG��x�����L@*xBhZ3���K'�ݻ��'���J%�ճ�'V�b��ں'	D�}����WD� E����`�߀�u�Ԃ���8�X���� a;�O6���jȑ^��X@��D@�3��S���DB�+T"R(I��9�%�����Ď�@-�.��l�d�6HY(%e�D���"cz����6k�I�CK��9XdHBC�S�2��H�Æ�8��\���$4�4�ySj�';j�]�#�
��Om�U���msb�`�]�Y�Dٓ�E��p<�EB] q�r�"%>?��4W5���끇t��T�	$tiKc���h�Q�i�` ��O4��<I�J($gͳ�'6H-l��'x8}�B�?#��~zTŎ	7E�D+���Ѷ�@�7VJ����"{>�jA��k��h�D&��2�޼\�EӶ��2�L�1�O�$�"n
�XΟvU �͚5FO� Z�'�Qs5Y�lL��hqσ�V�B�2�'آ�2�� US�������^�(FO&W2<
E�Z�<1P��d���Y"e#}���雀d��B�$U=x�������p<q��]�Q���;�"?�6�ҙ.`���<�Xc&�ii<�ɠB&}F�9���I-�n�9% ��I퐌A���&i�8�'��5)���Nזu��3� :t9��VG�˧dZ�q�Hi�E����TXd�=�p>I��"E�ƅ�6LQ+��Ur��f�R�O�]3"aPI�I�S���Fd�>���G9*�,�B҅8d�B��h<!�O�Lhd�q�>t�Rx�B��l��������S��@�0lH<�}�u�1l�pࠕ�	:'�%H"i�h�<���G�n��(cv퍴/�8�KՋ؃�|�O:�k�+�B�g�	5(2%X��Â\��A�/W�C��� �+��s3@��,X��!��:1�vT '�'~��v�H����`&q����L,9t'����+�F	�a�j�FD���?�fن������$�/5��Q�����\0�Oi���P�38�p�'U�~E�R�rT��ym�
Jb��ȓCT}��"
�)�)��E��W&@	A�UG�D˵0�6p���L>��Πv&�I�1��_7jĸ��e(<���7psT�d,+�
t�g��9"2Uc���3.D���DE����/^�TưsE��rr�xbDҾ|cxY�N�}~��&v�Y�I�5�(B����y��B�v�hڣ ��Bz��x�HdF�2�o���𩃑4w�$�.E���k��W~!��;z`�h�n�6��!B{&�+H>I5�N�~���'����whA���#��Ζ�h�'��@Ô�"�x�g�z���kfE� 3HM��ɤ)?,ECp�M�!���F�B�I
��[��y��]�AQ$��B�����K�D�
����CS?��B�	�O�D���,S=6�F�aD�_B�I��9��IT��l0W�%��B��qgZ��#��2y��A���MFB�	'��4@R�7g�x�7� !t�C�ɲ?�LL&f��VX�u�I3~� ��$�xv>`JA�6�"�A�Vyan�����	���h�B��ҝU��y��M](�e�G�֨�y�	�6*�ޑ�P!f��Ӝ�n1�(�CJ�`g��&���Q�B|�8r�&�DK%^;D��'� $�J�EɀM�@�S��h��͗&8�'?�xs�'�e�N]zTK�2����g�<1UIѬ^0ƈB��>}��$L2:�(ճPEW"�j$��/���C4��?_d-�!�'�f��̀9C���#�ְ��mk�*&}�ǌ�e	ԙ���O`���Fq��r�P� ���=��	�w���bA#j��������3��XU-ԕ_>t!�ƩQW�1YsnN$S�Bj9`�I
TP�9��(����Ͳ���*d�Uy P���ɠ4�rt���QU�O�p��'A�\�|ۃb�B5<��@���$Of���3��dF'(�5��n��;`8�F%�zo��:w���P��"��Ş67f�"Ї�"]z@�	*����V�"U���Ҥ�0?�Q"n1 �� v���ba7|�8I� A�)E�0�~���=���p$�7�V`�'���X���"�3콃�c >��?��&���A�4���uC�&{~��Q�@	~7��P�d\�4oB���)�'i
Hj��[�gi�P�%&�Txt���	;�)c���o�]�pE��50� +����Wx
��M>!���Vz�>�O"@�U��%�>|�DA�"8��it�>�"�(GGr��?� ��v_��3�!�1V&���=D��B1�H;�!�M{���u(9D��x0��"'cԥ@��
3B`$6D�{��	}���8�(��?u��8D��Ie-�%8�tș���%���bl D� "N	7/���abn��ʞiA�-D� �v��1b~�E�ǁ(l�~yHd?D��C�<�Rd�ׅ�~8��:D�$���� ��� ��F��	��7D�\�r)B��9a�%ټwfyF>D��#Ξ��U�Ex���K��;D�Ch�LXp��Ҭlp0E8D���K֭��9���]jkT���9D�����>N�ȄY6Δ�`�^l��j1D�\y��N��1"x�$Dz� +D�� ��P���;k��:���=����"O�Y3$ɘG�<�I$h�f�����"O����[z8"UG@�	w1ɳ"O�=�I�Y��,Y�ǚ�(Q�)�"O����S�j��(Z%��7i�A�'"O��!��8Ĕ�{�@TaQ({�"OF)�a_�[L七n��,Y���t"O���BB �� ϝg�p�"OX� ��� �ji�Ł�C�P��R"O�@1
܍zu�h��%��#��@�*O�`"@�~��1�b!ƋL�.�
�'$Xl27��/.?821��1���	�'����A�~\��p��6�f�	�'d���N��E��liuK]?(�H5��'�F�RB%�7u����o��"��9	�'c���wFӗQ��jt䑖h�l#�'hx�Y�N�[�$�r�-�Y	�'��`�m�(/�:���IΚ�V���'�8$�������`Ā9{J8�Q�'����k��3��1�ܳ*()��'��@��&Y-E���L��p+�'�@ݒ0慴U.������3�B�r	�'/��Q�㉔�x�u$B�~����'>�y�%ѹ�d���Ѽ{��6"O���끬���˧E9ς��"O*���O�~��4��$/���"OL�Q�J \�xxQM���0w�/D��s��ʍU&Z��ub�%U�I&�(D�dZb�F*���Ѕ-Մ}7���k+D���
S�g˲�
���'l��t�D6D��: o�'20�ը�+�,("�5D���B��Y�- 7 �]��aUc4D�Ș��2Ab��M�Y�B��P%1D�X�wIR�6��U��bNV�>���d.�K�?}�7�	vI�i�e�M:AH��fa+ғZax!�	B��eڷ�#0I�q�a��ēFa�ɐ��?� r�H�t���'���8�0ʢ���Fط8�L��	 Q�'�uwR?]̓t��Ӓ�KZ~�Q	ۣ,CJ@'I�-�P��G.��9�S>�[%c�$|�`�x��x52Q{# 8U3�I�g/G(�I5W0 ���Ͷ9����Q����@R�R��h���P9�~��ΆB������=���d�$芳g�B���N�t���'�$���	�d�p��CP�����	B�@���n��x���:}.�ڶٓ-o���dc9D�z���=g�=`��	E�t@0�)D�D��ʝ-F�|���R	?q�M�3a)D�
����{_4�x��<w�Е�A�%D�z7)�&,��ŧ�~S�	%D����_e	��s��^��8`7D���͑7\-@E��|qӥD5D��T��
Lɶ���!I
!z��U�4D�(�7���b�\���H2R���s�2D�0�fN��)���#+��cL�Db6D�D��MG:!!Lmɳ$ʈBiR�;�3D��j��/
]���-M_xP�g�?D�P��%�1񖤨��Ҏ=� �PG=D�8��+U�If	*��и)V��3e�9D�H�Թx- �d���z��d6D����6lVͪ)�5b)�`�.D��;W痃AV����]�{�쥂�j,D��N_�9˺%�6�Z�s��5P�A?D�8�qo�T3nY��+j��e ��:D���+�j �в����Zڴe��n=D��)�ާsO`YX"��Ur�q��9D���@��X�8G�ؽg�Hs!�2D�� <��"��6g��ꃋ� :Q�$[�"Oe+@`V?�P�;���NJ	RS"O
��#�%Ru��1'Mζ<���D"O�Q5�ȴHy� ڂ�q%j��"O��r���1~mN5��+�� �<��"O�D�"�ϧ"&^���
�:p�ހ��"O�}Q4o[� ���y6)ΘĲ�r�"O<�:�K5+��;�&�R¦1c"O�(F*�(������}�h�R"Oƴ� 囌e6`%������@#"O0�2��_=$�YCߌ{�2���"O��񂒺3���8�g	����@"O|�P�A�?F�j�!$��I7�*""OA���.��d�ek�`/�+�"O,U� �і0p�A@6��:j�!�"Od%�FO#=눩��!��VP�Ұ"O8�e V8sH!���>"�T� �"O� �b'��'IL C��0(����4"O��[�V.uP�`���R/sH���"Oj��Ł4m��t�U�M'�D}1"OvY)�p����=�t}#s�m�<�C'
qd�$�!Z+&�����q�<�����\�TĀS	Y+E��ت�n�<����V��q[���;@6���GIl�<A�D6o=�4 ˗9�(����e�<���N�N�P|��cΝC��j�cK�<�$�G�A-�L���%E�����nGJ�<����peCC�O��Uh(�L�<闠�]w�d��nM�>�@���`�<�g#7 Q�y(�������C�_�<95F�0��q�G,�]p�I�e�<���J7X6����҉
6�@�M�<i��_�3���A2�+�Iq`k�F�<��9[Π�H�� =FQ)"Ζ�<y����s�l𠧭ø]�<yH�
�@�<�I��/�H�c�4�0`e�f�<9�d�g�`���0A�`QaD�d�<�s-S������@0L���3@-z�<�Ѓ�.J��ԃ�Eܮ7N�k �t�<��	�R�J��և�'���2�	n�<q�&cڠ$8��%_Ƹ(� Lj�<�І�M<���cÛ=g��˦Ĉd�<Y�1_��9q�G����eW�<aLS�z�vQ������S�<cJ�a���$,�Ţ�{-�V�<�3Õp�l��ʖ�PJ��:��k�<�E�m�9S��!��	;�.Ci�<)�%��bpD�i L��B��e�<AV���g\�@�C2�΀j!	�c�<���E'fi��YѨ
g�9 J�w�<��Ə"?�ŋu�BY<�};�s�<I�еR�< ���5�&\�u_q�<��n,P�
l[6��u������i�<��E��;��aQ���-g�V�Y�c�<yv�-|ͮTBb̞2b�!B�Gu�<�	�C��[��ƂOu���$Hz�<q�NQg9`��BĊ?e�2ࠐ�[t�<��.�,	2. `r�@�� lXI�<ᑊ�,��W��.0jȢ���o�<�f��|�c��Z�XfD,�rL\n�<��c��r�V-"��\(A#�%�t�Yq�<qB��&~|���㗸���Iq�]p�<�Vm��gn���4C."l	���a�<�V�]/HS:�c
˧O[�\�&TD�<� �!��¯'U�* i�$�L處"O"���(R�<���O�GHt�X�"O����E' }ؐhV��<x�.���"O��j���y|���ƚ9K�(t��"O����H�
#r��tKQ��} �"O�"M��u}@P�߽sq�t�U"O�X��"]Ɍ��GKfXp-c�"OzX��ޡf.T�3��B�A|�$"O(}�4�&J�pT&��CP�$g"O(81��_�\F���P�ʀ8�P�S"O��;3��$n���;t���R4"O����	:*�т���v�y�"O�����Zn'f����3o*8+�"OF=2iŮ�P�8�)�%hp$]P�"O��V'K~<�s(Y]�59�"O�q�K&$dX��fؑ%l�G"O�<�,n{@5��ֶ8���I$"OttY�BŠj��IQ�T~$��7"O(i��_��@�M��0jJ��"O�I�j��+��<�Q�O' Upв"O^�rBoC.�LB�
��4]9�"O�ջ�iE>dX@��:�t�q"O��y�����:vGҚn��t��"O��� jE�E�(����������"O��!�2}>n�b�ؗ&u0$x"On��S��QB�Ӥ)k�S2"O�y��ݣQU�YC��آ6�T��"O@�0j	�"A�aZCK��k.���"OfVͣ	ZA*R��%lPdHf`�`�<!��^�-).��T!F�3θ*�H `�<�t�Ԋ'��y�V&�=�\���E�<i��}X�]бl�RkN*c��}�<���ޙ@��X�� 	(�^Щ�d�Q�<�e�6!��]ఢQ�A��|���IP�<a*�	�|3��A�?�x����N�<�vON��^� k\qr�r/�G�<�ve̟1P��(ǋI����'�F�<yQN�!;{���!Շ&<$9Pf��B�<Q ��F��t�vR&���V|�<�CǛ�5�De�:��W��y�<�@���T��f�KyD�����w�<y �N&����&��)$��f��<Qu�I��ĸ�
�g�\Ae/~�<(8P~d����Q�l�"���v�<!��Ʈm80sR
��j$�e@r�<1"
�+hKm��}}`�p	h�<qU�Ժ�陳-Z�ܒM2Z�<�
ߎu�����@@+�0rD`�<� ��2n�yt��?,�4���BG�<I�o��b��� ���>���A�ƟE�<q ��N�l�']�d�.��5�C�<	�Z�"t�x �U�B�l���B�<�\?n#�A�g�?��4 ��{�<qt�E
f[�1�I���$)س��x�<I4�
�l�
���ō&Hz��J�<a�&޺پ��H��l����I�<�D�]|���C�/U� �+�!Op�<��(x��� H�*�d�j� w�<���$] z�H��g�w�ħv-��[C*���Ҷ< �Yx!C��_"P��ȓ>̕x�� �6ך�G��FR� ��X���*)G1 {RW�P{Nͅ�w��l �.�"�.l���kt�x��J�T�ʣĆ��8�%�	ĸ���S�? ���4�^w =����7i"��c"O�!��� �xzT#ΊYFd���"Op�𡋾;�ΠQ-Y	X��#�"O& �&�D�V\�Bcǽh9B���"O��!g�J�	��}�F��4o1���"OF$�4d��t���ģ	���"OL��ƲO���¬1����"O�QR�9X��5 ��T�E�6$`�"O�iÑV�:�X}��V([��IG"O�ݸ�N�)*^(�p�,̖$
�`�"OL4s�n
$��=��� t9�"O$�q���I�|�cS�ž%&u F"O��`M�05�Urr�M �#A"O4�`�ĽF����� Bt��&"O,=(�C˨l ˚#�<��"On)��̀���A�DF$��b�"OҴa��]�7�~Y�3"óԖ��G"O�K�G�)2`��·Iќ �'"Oʕ��Ā�$��$Ȇ�^�'Ԝ�2�"O�@�4��-(�����7t��K�"O�T;/B4V�}�W!�1GtD���"O,=�P�Z�G(�V O�=����"O�T�����x׬�/,�hh�"O��1T�-{ώ��,P�? Pa�"O6$���ݥz2���O$l� Mȷ"O�����Q%|��7�B6Mk�h��"O��HA<U�:Y�$��>W�	7"O8�:C"�C���j̳Q�YR"O�bG�ؿR'�)*�i�7:�dV"O��&#Ѡ=�j�=3���s"O��+2dؽB��e+G*ϯG��A"O��.
�4Lp�F�A.349�"O�`ca�R�A�VIs֧3����"O����h�	.q��:�� 3{�d�0"O����;.+���B� L�(��""O4%q��P<p4�2b��:����yro&C��d�g���Y�ּm!��)|�`{t���'Z�=����~�!򤝏H˼p �&�%S$�<`vOB,<�!�$ج6��0� ����j��Z�mz!��B�_��!J�BF�-��Cዙ1g!�ć,KG�IdI��`��0D*štf!򄞝r��M��AE2nЕq���%6!��P-d�r��K(ǞyK��\0�!�Y0 &���㚯o��5��;C|!��.��@1��8}�����%y!�D�K   �    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   �	    �  )  �&  #0  g6  �<  �B  BI  �O  �U  \  db  �h  �n  2u  v{  Ԃ   `� u�	����Zv)C�'ll\�0�Kz+�D��8��Mے��<�&E�H�aM���vo�^;NP)�A+.wȜ�2��O��h(6e
�:��1q ����u�cY)��te+I��TK7�<��`��cU��'� 	������ѻ�l軷��!8Ĭ0������]8��x��ߟ�k��� ��iHF�фY��x�ul��f�	JF�� �?Q"�S�&8h���Nś�gvq��'R�'D�`T<x����D� |cD&;a��'x@7͐����':�ӉD��d�'u���#5|� qn��N����DȦG?�(��o��Iɟ����?!��H,?���;7��a$�^�A$�ؓ~F���'�~��6���9̐e�2�_M굱�OH�A�9̄e	C`3�6�a��Μq���L�J���'f��'�B�'���'�������T8 '��"�ҵr��{g�T柄��4]�v	�R��'�26MKڦM�ߴ_����'� $��Œ�A)!K\c�فU�	� H�>�Ӻl��1%�W^7�{���wB*I�v��W�ʰ�e��C���lZ��M��i���x݁��aH'&�Ke�ő��h"ehXb:z�Y4O�ݟ�ɴ��(y�%��#]v��$��+pʈ�$GX8�M�S�i_.7�z�h-�q�	�hm���B���:�"7��=��	��Aۦ��ݴj���ET	C�*ccHGB��9��E]�y��9�ʛ+4Ǟui�`ѹX�5oO����Bs-�&q7R����۴buv��C	�3��i���C�H��b�J��}����W���6��p��&�G:OJ���%�����-ƨ
$��F�t+������r)��ɅUd�a�
j�lZ��M��i���O��x�&ۑnQv��'�'PR�k��ϥ%�z@8�F��(��"O��#��3x֝H�I�.�"OnEC���T��d��YqU�"O��$�I�=�rĨr/ϲ��  "O����$K�a����KT^�X�s�"OF�bU�N��܂%Eȸ	A�3���$.���~��,��XAc2H	���U�<�E���I8����N@�>�I���P�<ѱ�5
�ֈf"R���IM�<I�+�l!�$��t-�T���RE�<�QC;i+L�����Cwj$ZN\A�<��GM:fny�lQ�f\��у����X��)�S�O鐀��ޚl���B�/"�r�a1"O������*�Da㠣�E0�["O��2��Z3)`���ǳh�X�"O.m:��,,D���'�D?�(�iC"OX5�bb��aw��	5Fأ`נ0�'"Ov���ɇ�<:���E��.�2�Z�3m(�O�Z �Δ^�(���M�wI�L��"OƩ2��X-�������C�<؅"O���0l�+z�CE��\�ze��"O��r&�U���eL�u�P�E"O����f��4�$��^�`�'���q�*�Tf2�x��Q�F�d��	�Du�����d�O$���O^���
�u��T��=g��=��	����jH�� �C�����Ʌ�h�W!��w����	�O�łk�t| H�bëܰ	��'�RX���/{Ӻ�dW���vI6�B\�� �z�˓�?I���iÁ*�$4��̈1KY|�mh�)���Ĳs �4�B�M	P*���?+O�Ѐ"�O$�?���<��	��,�,
��kU*\Y��M~2��%�`��=E��(��)����A��+q�&����ɝ��Ă.f��y�{��i)T+�	�nA�1՞��׭�.����Sc���Oʓ��c>�xb�t�\�w���u��y	��7���O����q��(C�X��С�[�����\�O��0HDt�����D54���i��R� {.��?!F|!�z���&�wм�#��TQV�ӤX�Ze	Uq�1O���:���a���l:��HǟP�"r+O�d��f	:/_1�1O�؋�(�TS�2a�Q�m�~I:��'C�	�e۰�D(��O��$�O*y+*�@1<�3�Y�F1ht�׎)D���`%M�D3����(�0p����<���i>5��Hyҫ
;Z��T��>�h%aW꘩w��r�'�a|���\`���Й�� 6c OY�U��'�8"��և �l��4E��X��x�"և��ܫw���D!��éX@������x��I>c�
�d��?6hV」��y�C�D����D N��p�qB����1a�F�|���{e���?�t���\��M��zi@qW�?���D9"��?I�O̚�8"ə+E 9�"�Z�@�j��  ç

�1B��7�R�L1��Q��/���"�@Wd�y٠U��)��-�u��(��<;�	�(9�-cq�*�M��V8y2�2�ć7�"�'��I/K��T�'/N2$X�P�`L�O�8LOޅh���N%��!���p����r�'� �D��E $�pfk�6v�0IbD�[%�U�h�!͒ԟt��˟��Ol��S��'$�W��rD��
�˴!Eu�p�'�B兵	a`��B\�"H���VLH5 �'��	�UD�l�2�8����w�[/=�ɫ&���N.�2��4$dA�;H��@����=��֝*��d����*5	��dO=xGx�V;j����G���'C؈P�E�Q)<0��JKnM %*O�
���B,��獘+N- ���_`�O�)����\램���4��Ԃ�DR"��r��(OT$��%U9'f�g##rrŁ�"O�e���R(tC�q���Q	4x���'F3�c�-��c�w6`��'���d�$E
��r���p5J@P
�'�jɢ6�Y�Z�Z2���t@���' ����(�f��A��;��1Q-O^=`B�'%�mR�K���JYPa皧}��Ա�'v�� ���xshX�tSb9��'u�m	w�8)���R�ad%�ȓˈ�"r�
�
�"��N/L�=��������B%%��Mfz���I2����17��<8�F���$��&�K�C�?�
P��j�i�"dqg	?J�B�	?�V���N��� �(�:8C䉾Q.���H��G��y{���&$��B�;P��pFƛ'�T`��״V��B��2\>,LŊ��jp0젷▦/��=�E�Hp�O��Y�ˏbpR����C7d� ���'5d��b6*��]���)Nz���'N�U:e��kaƀ��gQ��+�'�M�Մ�/a����a�׎ O�a�	�'��  &�(k�\tz��J��� �	�'�Н�cF�* �`� Ù�x�	��@ɞ�Fx����I��0X$�V.4����C�C�	2.Ӝa��F�<5T�p�_	4�B�I�\A9��
`�]�t��M�B�	*qy���d�Z�P��� a6VB䉳�8�A�*@SR�H�:)`�C�	&t��T+(�7����,�R���I�]w��k!$*b��ɤ4B�c�rL#�\�%b6u:"���-�C䉗r�"���c�'X�@U��ZC�	�(�.�!q �P�6��1�R��B�	/)l�yG�:K�����@9�H����e��O�V��Y#�
��X�8��3/͇M!��.l�2р�@����a�0!�䑏m�$X�pi�*K��j�ڠi!�DL�A�����L�Q�Dd�F�   !�$�Yx.��g	�r5�
�mY�qD!�Ď�"��pL|���Ҳ�B+9ўK�D;�'L|\�5Z�""�1r��\�\�ȓƚ�3A�0XC6a���
6�~��!@b�Ĩw��a�`�oB"1��*ڴ��B�9�R���ɪh���ȓz�8�3�@�Lhֱ�fF�%o<���ȓ,�\]W@DI_B ۢWE���	*��#<E�t働�l)h��@=���銺f!�D��	U0��F���X�燞>T!��'|�l� @KP<%��`�a�E�*^!�$�?HT��̐!�����d۽6N!��$͚8��@J� �p�^�>!�D�7��"��7� �� �則 ���d��#{�`���Z�9�`�Cu!�66 !�� �a(�D�t�(��d��8[��0�"OFQQ2��%��3t��;��"Oy���
�� �A�A�Z���"O�@�@��,��=����B�h-���'q��h�'Cl�A��Q����&'Γ>�,<��'0h�@��L�Dz�ܫU��64�`3�'���Ў��u�h���і;1LS�'$��Dl��� $gC>�d�
�'�B)��*FRp����7L�l[
�'a���K��s�"��@��NƊe���ę'�Q?-�v!� s*�����Ȩ���!D���T(���ّ"�Z�
l���<D����I�����0����t�:D����#�	U|����K�l(�&�4D��6��$ȸ�:4���`DN ��	-D�ȢKM�X<8"���2>|���O*�r2�)�'5���7NIm�t8�D��V��s�'�6�R�M
?�*$X�$����'B0��O�f��q�΢4x��'wZ0��F<K����)H*�|�(�'���B�g���sC�߶�
�'�(�:A�7t��!�cC�Be��(O.�Pp�'n�ʥn�8H�v�b��3P�-��'�$�S$����BA��F����'�
�KCFT�
����1+RU��'t��X���<]4���aS.(�@Q)�'#�c�,V:�t1��N�$69�	�[������0��2-�lO��N��T���ȓtɼU�w��<&��<�BB�?�Nt��g��d�т������f�bNJ�ȓh�Dw�	@;�|ÑIU>~6v��ȓy��8�dK@օ��HP1fH���ȓe����Ʒ8��P6܌E{�F;¨�8)@���Iu��V�^.C`�Q�D"O�hE&ۯ`p�h�	�)c�i�"Ox�!E]�z���T�М+N���"O�����.J(֐�Έ6t=��i�"OI��Y.-JN��f�&<�y�"O� ��J̻77��#/\ -�.0�F�'U:A����*2��|�cEƲs��=��G>a��a��BغAҍיI�x2:d�8���?ስ�ոn~깹f�X�x!�ȓ6i�$ÙH�16�O/L@>���=�jM��."R��V��,T�$�ȓHbL9�!k\�Bn�����(7�Z%�'F��B
�	 ��a(�0L���w�L
;}VЅȓ���H�}ض,&B�8����oǏ WN4qf)D�Y�؄ȓ91�����[�h+��x��)˰���,M��Z�Li�5���P�bd����i��I�{G~��b�;It Ȣ�LV>ĘC�	�<{��i)s$�@ o��B^rC�ɀ]���K U!T�%�Ce(�6C䉱k���%�<k �=����)��B�	>+
vX6�+���j6��W�B��f����ކ+E�q׌#|\�=�F)]f�O����旬[Bv��CPϦ�q�'\��ݾP^���в9����'����h�,H���"&V�;�( ��'-��Z*c�|9 H�&b�LmH�'��1�AY�T��ؚr�G�.c�d�'��(qɗ�.[ �1iW�-����mh��Dx���Ą>���Xd�
�M�L�0
D< C�+?��5k �@�d�*rfǊm�C�)� �=��)F�0����Ѕˀ"O�!��	���!IA�&�d��"O,- �M�>�b@Q�!�Kڦ@;6"O�i"�E<J ��҃�V�cb��dX�|���0�Oj@i$���)� ��W[��("O`Y1���}h�i�dJ�6)2!"Ody��O:U	<e��$(0����"O�=�&��za1P�F2���"Oν�G��M�W"��U6��1�'��\�'�fm�'(�-:�ThS@�ك_���'��m�pJ�2%0��(x��iC�'��I�Q+M/Kt��WA�^n���'N�qB�l�
4BdY��kR5O�h1�'y�!�Q��!�x(W4?"�=h�'4�9ae=��Ȣ4�	-b�������29�Q?�IPf� r!j��$�y>�U[0c"D�(�2�W3���A��l�H�Q��5D�Lb�&1��y�����%�B9j�!�R
U�~q9C/Y��>	��cu!�жC*pҫ�V�,x��&�!�d΂(�0A�u��;g ~u �ʇ7��̋�O?��&�B�N�Rq��,V+cpD-�"�K�<��FX�_K�2���$�Z���D�l�< �L�D<b�0�'Юu��j�<�gB��F��Q����j���QF�P�<)b�{sL5�2
��8<��	P�W�<9��
# �p�5g�
n����Wy2�#�p>!��Wjj0���t� ��DDT�<�u���R�]�G��[Е�h�P�<��ʻvj	��J$.lhE-~C��0����K��8�˖H�M�B�ɩgX��"S~��s�G2FB�����9��3NP�(�L��]r���%",D!�D]�:X�(ր\�ii�ejaҟ>!�S�|S��"��7x�|!��NQ�_!򄐈S�Lт�D�5}.%H��"9M!���!��!V��ic�ő!m�32!��x2���ԩO/\b�kjէsў�; �!�'`��:ޡ�"ϣp#���Z�m�b�T�`���J�o����'��@&�QHX��cfݞTꠇȓY=������{���ѡ� Gi���ȓ=��w�ե%%F�v���@PΙ��z��&�Y0+-�A���<�B����}f"<E��j^�#X3��?R|�����]$RA!�"k��!�q�ʴKu��)S�b(!�9e��QNQJ��t�%��!�ѭSp�\��%�<z�Ԁ#��N�!��W�p,�6B�mj6���G�!��ʼ@�:�x��_	g��`��ޮR�I� چ�����M/��P!G�6�|�+����02!�ݟn1���7$Ϯ�ˠg��!�$� r��ђš{���p@G)K�!�$�(]��l�/7|�	���E�!�dGZA����Bip�n	�5��}��4�~�mZ}�܉�̓4���b�B_8�y��O�IµI#F^�w�>�����y¦�G�ܕ���8r$�H�,�y�D�7�B�c�I�p6�8�h���y2)M�d{\����@9�N�h�n��y��=L��� q̲.C�9CgΗ�hO<�I���$ʒu�s �9Y�q��L;>�NB�It
1����`�
��#�ShB��9�^�C�
�,Ij�hޔ�@C�)� �,�����J�k���=4�p��D"O�
V'��0�D<s�+�{��i�"On);FI���dY@@��� ٣��'k��0���%���C�MZ�5��]2�`�2����ȓm0�]a!�*v6���k���$���1G�W1Z���Y��<z38=��i㘨�����H�hV�J�x��ȓ
�fxsfP� .��@�e�N����*A�T�F��N�,����j�.9�'�ĄI�tV�A���M�xJnx��oL ��!��a�j�p� )�܃%��*�ц�b���0tCӝ?����4,��`��#ոI��O���kt�ߦ-�J�ȓF��	�4��>0��;�` IM�a��ɸ6�@��8 Ū�R�m�.R��b�	��NI�B�I'�2��"���*6B�	�8���H�������Yq��/,kB�I4wi�e%"��
BA�;#	�C�ɘK�=�mӖM�1�Tǐ+E�C䉡<Ƃ���D�
�P1��N�3�B�=��PN�ODY;b/
<d��l�@�/9B�'Z���n�LZ`u���I�r�	�'�j�������w�>�bp��'ӈ��r@�L��� Oĥ6�
�'$I8��QRT�97��2C�qJ�'�$�k$�֝y���M�0B�R ��9-� Fx���ѕ8v�A�lB>�9��(�s��B�	=eS>ʡ�?��#%��'��B�əV$	��[<'��i�u���]��B�	�q#t�&F�fN�`:$�DB�<D�����\�1��"p��>~��C��;5x��I�f[{�� ӥ�;�l��[��+}r�ϥBK��+}�&Q�U�������|ı�i X��ǟT�	��0˦l�U@x�	�+�A@VI���|b؄A^�]���";@�I�b�1؈O�8r�.F����D3���'f�H9P�DGf���2&�(�8TF|���?��ϘO��	R��*:�.=���XZ^��/O�������h� �5��#�L�O��}�%�<�g���;�l�B�+�=�����Xy��Ǣ4�r�'{�k�t�'z��C&s�r���7'�[�@X�	B)M�b3��rèƸkF��r�O?����Rq?vP[cM�0_� �Db��h�Dʮ�z��-M�g �\F�4�w�T��㡈�tD����y2)��?i�������\�$���cנ}��G���< d�.D�̩�	�4[�{D�GJ��Q��.�E��?��U�T"��uh�a�ѹ��O��'2,80T�z��$�O��d�<��l�]Ҡh�/|{]` ��rߒ���W��?Y��0x%�/�A���dB�5l:t�7��,7�lrֆN�� @�O�EQ���=w$q���?#<�D�F�%���疈�Ġ���]t~b�ϭ�?���?��2>�����3D � 7���F�tIK�"O*5�Rk�>E�*���N�q� �.���$��|�����$�Rf�X���N���z��;>��M���؇y�X�d�O����O����O���u>����2˦��ׂL?��8�aZbs��ف�X�ne ���ئ�B����|�*�&����0�∮w�B칇m�?�|����7F@6m�=�z����	q��zJ<!��	џ<���¦��=�Uڌh�ބj�֟�F{��I+���u���D	Fb�Z�B�	�kY�K�g\����Uo� ?�����'#�	/9h���*�$s>鰱�Ӿ4$q�ƈ��Jp����ON}�D��O(���Ǫ������G,��'{V�lZ����ύ ~�Y�$�F�Q�`��T�'��$�����Ԥӎ�:]~��S�	R��Έ2|�16n�<�܍��n[�%)�AM�	7#Kr�d�O�c>�I� Jт́�	�3����'�<
�G�.p��
��n���\�LXXh������D6prly"�#�P�����5�ɽ@d���	 (����Y���$:o���'By��[�T5bT�SOt>HF�'q9٦�ۊQ���Q���tD��!�~"��d'\��^�a��A�H��Б���'�y��Y�TƤ�ת
���B�aR;��@7�乪��B��i�u  �C�J��R�fl���*T=��;�2�'��)���Ot�)� `��6�Ɲ:�N%���?cz�MC�"O8<�XnFm	eW3g���7�	��ȟ�M���� w�R�r�Ã�DM&)[�+g�����O������I����O��D�O*��;�?qB�� 5�=�d��e�0HPM�
9��@3�#}�.!E3�$������T�d3ZQà���e�>A�6�T=`H�PgY+�f@��MS�H�Ju��S���i�����X����1���Z�,[6j�Ĉ F�g���7m�.���O���?�I�|rf-���^Y�sf�:C
��K�T�<YB�d�!�(wO�DT*]I��D�r�����'81O
LaW��p��q[�oE0���J�'z&���1���0r�� :xɂl.tI����`J\�@�F6P�F��T�[��*O� B�I�gB��c\-W80��'��i��N�P	��dF
��M�ȓ(��G��'���G�O�H8�Fb��r��*@+r:��\#�#�En�x���<WtX� �'HRt�'.B�'�Pв�&�?Uy��� �:9"2�h����FH�e�u�ΎX���V4��O�Q�0��<ТUyc�I+��z݁3��ϝOZ~���.�)Fp��QAS�7&PЧ%�W��'hL���?y�����)b�OR#;e�������$�O���$��~@�T�K� g��Q�G#ln�}��<i$�
.{j�����T�z���Ry�'=b�'Q���w掘3��D�1��E�6ɒ����y�'*��à��'z�6��dg�&N�����ɗ����O�0����#1ܬ�Ӫ��?r�@��ba�N�D�5�X牑h9����On���O�����t���(F���eN^�E�܅X���ꦥ���������<��Wnz�!�ʟk,ݦ*
��:g M'/?�<S�@K��m��?�򃏧�y��8�d�O��)�O��I6��%#�ϖ�g�&�x���'Y$�IK�O��ąA��db�,�/�?7��h��O�hZr,Q.D��d� &�#EC����'�=�	��4RD����	�OZ�������w���%
�W��L(� wT<��		_����Ozp0���O�I,S� �s���º+e��5W".����^*ft�U��d�U̓8V����dA��%���?!�'�N9��D!Q��բ�ˆ�0���@��y�n��?A����N�OF�I/j��s�`1C�n�&=�n�t�J�M�`����A	2�b`n��<e����M���i38�i̟��	�`�O��#�B��Wc^�yT,�r�����B��	�<Yׯ
ş��I�?����<���|R�Mڐ,=TuK�A�D���)��A��M��EF��?*O��d�O1���$_9@�E�
4=�;����BC�I��IJ��0���WgN�M듎?�/O�$&>��	]��Y� ��q��L%Q*��i#N�#=���T?�U-҃+#�5���Es��퀣k.D� �G�W	X�2�*7BN�5�i,D� ��
�~{����g�V�t���*D�l{��-�n �F�\:hx�'D�ȡ�ƀ�@{��Ce�F	:� ����2D����{�p,��ŔV��褩/D����G�Z�T9�(C�ah�u`8D�� A@�)R}���(N��i*A7D�\��ꍆP�YP� SY�؁�l4D�$ɅcO�G�̊�QVT�*�'3D���ū��w:z�c ��C<,�Zvd.D�@���Y�.:e��R�GD.Y�B�I9����0��K$���3@s�b�i�l�:�:���?X�@l��Պ�.�A�/ $*l�, ��҂~���1���i��H�d�:� ]��i:�������4n�A �ߘJ�6!�e��U� ���b��%��4#�^�IT�Y,����X�C$�9�bj֙N!b� !U�ELd��'哭��m ���oB����wӼ Q��Ξq�J�{��I�HʤHj��Kӟl�I>.�@�+�. 9Qtҧ�i�~b���iQfa�K�7�N�RD�T�ɂR ,Ms�m�;��?��� 5q8@�4 ����'�Ni ��'���'��4��¦��W��T�@���D@C���O���ǥu� 	���.�LMcd��~�x��/�a���ć�x�[1DG�ZwZ��'}��'�~1ӢJ��2��<�F�r��K�'�^�I ă.�ع+#��r�њ�'и1�pʜ�m��̺r �):=��'��5
`*�5�<���, C�!��'��&��*N�P�񭇁%BL���'����RA �F���]�$���1�'�f)���T�(��{pcӯ"td1��� �в��1RF�<Xo݁<��b"O�D;͕� $�5�d��m�`,Rg"O��'ޑLf�U"��K�`�p���"O���i�9�8[���BQ�l��"Or��F�(~�Q�Z�%7z=0"O�b䃘Bg��S�)
�H��M�"Ov]�!�U�9���s���Zt"O�i�/M!�F4�e��y�	�1"Ox	�Eo�F`Ւ�̒7hj��C"O.
0"�GDM�`%Fmp�z�"O�1�7�X�h��<��Y1b����"OF�v��+:0���#C�2�v�b�"OHaD��+�D�GIY@��!�5"Ox R�H!�Z�����5� 5[E"O��Z0CP;1ڢ�+�e
�k+�"O�<�`��o�4H���ޏp�
)bc"O��;4��X�6��d	3G}�䘡"OX(
��/�8A�(	�����"O�8����$) Ai�(E*�"9P�"O$M��*U�X\�B� �j��3"O�9� �O�!Ybܽ2�] �"O�50$	ʈwψp �@F�+ @� T"Ol����5G���o�P\�B"Oy!�/��Y�l��gϏe���ɒ"O��1���&51� 0��x��"O�l����-0�t<K"%A<F��eJ"O�a�u�F�/�!�$،)}�,R@"O��K��	�5-�H��"O���a�ߵ{�P���D��"O���Ҡ��e9t速J�e��"O�0�+މ��	q��6x ��Hq"O�`���'Sܚa����A����s"O.��W�����
���4����5"O��!&�&!'x��W���M}��s�"OtUБh��y��PX�aHs{`�x#"O����o����醔k��5��"Ob�B�dA	M��aH�Ѩ���"�"O��A�B�>nq���r��Y&"O0�s��+UA����7P���0g"ObqഉED�"�H���|�Z\u"O�`kA���Q�)��(�R�De��"Ov�)
q��5S�'܉(Ξ��"O$�����!�fTɒHZ�T��"O��	��ױ!������4x�j#"OREhԮB�tT�"#�X�f��Jg"O\�˷ ��.iV��CH*t��+r"OU*gƜ4�R��bg�t(h)�"O,,yB!܈b?����
����+\w�<9������GF�ub6����G�<Y����:���PĊݪo�I����F�<���E�OT��㡕(P<�SQ�\[�<1'�֑�)�B����r�XW�<�� Ed%j��ݡ,�:�d�K�<���-3�@"�JtR!�aH�K�<��K�m�8e���yŴt!C�KG�<ѳ�.-h�#��?W��!i���A�<�"ޗtu�|9�Ĝ g�hy�v�r�<a� #��M�"�P�0�� y0��y�<9p!�
 �a�w�у/v��Ppa�o�<�A�U�{��b�kO@��)2�Fu�<��I�W ��`���"	.�#���p�<Y�队iV)�BM��
��k�<!`��n���v�`>|Z�K�h�<Y"iD!OW2DB3^@���Y&iQo�<� ��Tďr8r� ��5��9��"O�9rb�R-�>�y�D�Xtʔ��"OҍU��)������Ϛ K���"OX!�KZ�|���C�";�Q�V"OnX��%�!x�z`"i�!�t"O�0���� |^u1�
�,��2�"Oz��R"����W%0XRuh��|�<�c��-c$0	����|�0s�Ua�<�1 �1	�P��q��7�(h�Gh�<iW�Q~���j�@�E��[B��`�<	���+0�JMD���1�|UpU-�_�<)�%P1F-R��Rx�A ��^�<	V�G�޲p�Mũq8d''QA�<!����R:�\�2���N�:tҠz�<av[�W"��wb"r՚�:�r�<���XF�ʩ{%'��j.��qv�p�<Ѥ)T0d��E+#�B<�����@�k�<a A%B��`�V ��F� 쀥��o�<q�I��ESB5Q�-ܪ��0��B�<Y��[-Ұ  %�]�G,j�
F�g�<�b�')�};j� =L*�Y�Ta�<��c�4y�Ƥ�����u�<��;9��\�g�?���	Q|�<a��z�V��tNC=D�]���z�</��#m ����z!��z�<��h� ?$�����6 9�p��j�A�<	���(�Z�"fS�2�T!ba��c�<q3釐E��I�/��DU��i�A�W�<i�Z��u6�3����!�$$��=��#Ȗ.ڈ���!��<?�b,���4��ݢ�+G&4�!�$��A��U�B;C�	3�h�!��W$	v<`�D��QV�W��#�!�$[5XߴXd��'$�6Iȉ܎C�	�A��x���W�^04�bKȌGoB�	��J���K-R*0��+D#B�ɸ[���A���XقƉY�C䉆q�.-Y�咗���s���2��C��c�40�u�X�Uu���̞���C��/Y!����k�.�hK�
;�B��  Кa�P?#�X��1ă,,dhB�`��i��j����ŐRn,B�7�|(�e��.�><��+�0Q*B�I�c>��8A���>価����	FwB�ɇ	�����ʔ(J�g⁊m}B䉴M2�My���uy,|zUE��DB�Y�\h��E���d"5iH�n��B��g� �Ae_�޾�Pw�Ġqn�B�	�	�2�ba,�	����G�/T�B�U<\pF��ln8Q�	&�lB�ɒ~�Ir��ҝ16�2�kR8#`PB�I=NS� 0�ʼG@�����n��B䉾a��됬K�,�����(m;�B䉾J�T�z���/?��;�g��fB�	�fJ����������Jh��"�4B�Ib�����G�'Y�t���W.H��B�ɇ>l�+��)����fԦ%	C��/d�]P��h"�=�LR�$��B�I�,5�� �-X���7�T�C��8AS.����	i�V���ũ4J�B�I���%*�BE�^6.� V�D�nW~B�I����1+T�f��V�C�(�LB��:Co�c�ǧa�qС��\��C�	�!�4)T�ߪ8>�M��Ǟ)shxC�)� �+�hF�u%���a��'pF�`�R"O,��am�}�z��TÁ�o'�41"O��G��7QP�R�M&'�tڣ"O>�����* e>�B%��x.��7"O���@�^QE�Q@��fp�! �"O�p�F���1��׃4Ɏ)�"O�x�Cřt���BG:v%���7"O�5�SM�����;2a�J��s`"Op(����Y��A:�����(�"Ofu�0*ܿN�Di��Y8	@E:�"O�0(F�$��Dۛ},h�"O*�!�X�8,քJQ�;L��Q4"ON���:$Up�c���~�P�"O�`��w�vD�MDv����"O�X�׬�7��l�c��)shx�2"ON�Th��:��	��LҬ��E"O����\�K?P�AT��
�t��`"O��`e
d1"򂈝40�F�*E"O�Q1��)��̲�!{�L0&"Of�z!��;gx���E�Du؍�"O����]o�& vHǽA��Գ"O���@%�)r���z��� �
Db�"O~qg�_9��@�ɓ1"y�H��"O���c�T��Rt)Ӝuո)Xw"O���/|��!f��)��`�W"O`��?12{�%��%�S"O��i�.E$��H{�����f�_^�<����R:L���±$V��K�h�Y�<i���t�<�F�
�]�4;� �[�<y�݋"���y��!Y�yA��DZ�<!��47�F���u/v�#�O�<Y��17��0W�\�5[vѠ�M�<Q�- \`$X����S� 8���c�<��A
,U����d�P�����N^�<�G��/x�
��t�0U&��d�X�<�S%-qt�!������aw�G_�<9TA���A��O(�����^�<��#�HZ�+c���-�X]��FCa�<�4�1=�̉�)��N~Н8��F�<1U�]�&��`��hQ 	��D�<�kATw"8B�c��^����z�<9D"�&'F�t�ug�:����ы�{�<A0B�-"����
��#�)��#�x�<)@iӹ&>.5hv摡1�6D�4��t�<����()$���)j���6cֈ�!�$t����'�W:����*a!��D,,>�)rDG	)�H�H���!�����
1D�' |h�i�睭#�!���܋� �`W��#u�!�d��6~X�
�t�� ���^�t�!��h�&� �
�"Ӭ��ƮA:+�!�$��;H�R��>d�bH�uB��!�RV�6ћQ��(ْ�X!D��!�J&��!���K� �������#�!�dq�	k"�K����{֯��v<!���"��9���&�����P�N!�	J's7�ȿ3�.��4�,`!���^1��s$���HV�0R�-^��!�I3JD�׌DU�I)�m�a�!�/JRPu��D?��KqkK�!�$ %o"�y� ��-�P)zs�#@�!�"�șL�&�*@cڤ&!���e��`B��"~Vt� h VF�lQT& Ĉ(��cM�/����$G����U�D�`�=B�L�>0�!�� �Ѱ��D�E,�����6�`�f"O& t~
�R�F��F�4 �R"O���������RRFD��%j1"Ov,�
�2R�xä�|ńC�"O&��1��q�V�(c-U=Z1J�S"O�%��N��Y�&L�X"F@g"O(U��*ȬSĒ#.B�lLaa"O��ۣ�NMcf�AЍ
�iWrk%"O�AA��0,�(1���WH�Ł@"O��fgZ����sq���:
��"OƽT���BSΑb7��#�A�S"O��9#o�22x�Ã��~��'"Oεc���6<�lf��.$m�X.x!�Gv-"٧�4�*�E�Y,!��)�`22�˼X�d�#
Oy!�DK�6�0˲b��:���c�T01l!�D�"h����(��ƈD�T_!��*�<��wƀ/p��q��OJw!�$��\��"㈀�;�,�!'m!�c�x�0�M�L��C"�� Z�!�Ѱ$2�y0�,���ؗ���!�΍OS�u#C	��UÚ��AC�n�!�d�3� 9�/�9)+n8@��|!���fz�d��Aˮ~�4sd��
|!��K�~y	�%I�T�֫z]!�$F X��9!�F��?;���Kۀ"�!�q6�8w��{'��cǊ�"�!��J�fH���SN4F�V��� �!���,�h4�K�;a�<�#g��!��4�~�i�U4=�p`@`��!!�Y����:��'Z-BІ�p!�D�fB�[CE���*���)
?!��{������wĜiC�
̕L!�$�2�T(r�L�`�
��"����!�dC)x�R51h�b�l%�T��W�!�$�Q���{׀)�^� �OS�!����a�n�
5�f���&�:@!�Dٍ E,�� GS�>%���3&{!��PI�	�����fy �y���MI!�D��w��I1�/!!	��Be��x�!�䋧OqΝ�6I�"sq��q�睐�!��4�`K�l�=Z�>���%B����8.Ѳ����
Qe�zG�T*�yF.-`�ĻN�?��u2wÞ��y�F��Ȩ��cAH9�%	wI��y⁃�y��i�K*p��ɫ�JJ��y���*[Pt���.�����(�y��ڵl���2'��G;�h٠-���y�GE�t`�e�J�l��m!/Ǒ�y�۲s�(q ��aw����nS�y�ux��S�������3���yR@W�\*b�����p�ś�L��y��	j )�s*�<xݜ�%���yF�2W��X���8pGn;�+���y"#� � 9S��:C�e�ԍÍ�y�.ڳw�0hp�b�Sa���y��ھp�B,�D��7�N5!� Թ�y2�ׇg%��(A�����%���yN� g���8guY���-�y2��<kV�j�,�!e�A��y�'5clZ|�V�L	w�б�o���y"�P</�,�HTi�"4�7iF�y3X���l�&=DN`�"(�y� �T�Ak"`��铅�y
� H��q·	ylH�!�� ��0��"O���1L%zgP���1�$���"O� ��D����3�hZ�'�PJ�"Oj5(�bW2(Y ��g	к1�*$��"O��B%�iBV��b��IH���6"OB�W��&�r�KΒ ��Y�F"O�i�� �r����s�щR�
��"O���vCJ�&�x�Ҕ0�x9C""O@P{��ٓ8�&��"/�x�����"O�����2���am�,�d9�R"O@l{���h�� ��
��v��Lq"O�ݱ����w$��3I�'yD:i��"O�=��M	�2&�`E���V�C"O:��0	sb0��i~S D�e"O4�ۄD�5�>5�'�Ob�ke"O�-�M͟r��÷�ˁs���a�"OxH+0ǅ81:!�@=D���T"OB�E��MXj���]�W_<4�"O�,Kbj�c�(��-N� ��G"O�\���H48~&�S3OT�� �"O�(a׀�0��x�`Άu��AA�"OjH9�ƀ�O*�@A�0 �zUb�"O�m`ȏb�*�R1ރ\>�50s"O����A4N��Ջ�h��"O�Ube�޶I^Q+Ł��$l�!�!"O(����"\�%�S炔3M2� �"O�X�6�]�"\�ZV�\�
dv-�@"OIx� �c�$+E		8���'"O��W�l��Rn��{�@�Q"Ox�1�Z=�X9��g�!�"O��&$X�X�lh�"� ~*N��"O�8f��;A�3��$r4�"O�(�sfS�Uz
���D\�c
�aZ0"O>�-Y8�óK��!N:� �kI�yB��U��۠��0dTh)�cy��hD���Y�5�vX��KԈm�,<�ʓ,�>���@�ےp�  ;>�C�2t�e��aT��j��Ϻ&u�C䉊Q�z����_ϲ�:sǚ!5��B�I�q���u��Rq�t(��+K��B�	�~��A�7�� ��Hؿ}J�C�	=-i4���i$�p�ss��QI�C�	�������7�<c�(�O,�C��2V�	��+_Kb��R��:I�BC�%��-Z�fI1"M.�s�G��C�I
=�`J �^�3b��#�OY/�4B�	k��	���?��yz��>�B�I�7t�c�S�x��@Њ�$�B�I"h�0�iVc���q����J� B�ɤ8�^�s�/�;�l�@cE4B�m��lJ6$ⲱ��@�c^��a�ĠC C�*i��+H6U�����c]����/�1v��br	��-����ȓJƄ9)�;W�x�z����IS��ȓ`H��AŅ�?����i�9��r�VM�1"\�PI���H� r�^���i2za+��S�h�0Sc�~��ՅȓI�e��	<T�3�@�3}�|�ȓh'^�Z���s�xɠAi"7T,܅ȓ6�d� 5�AM=�H��p7�t����-^B�,��`��cá
8t��`V������}'�9���[=J�Ѕ�ȓBe��l��y̰U�V��2ͅȓB�ZU3��H=V�T�X�c�N��S�? ���!�ϲf-�-���S�ڠ��#"O���'�)Z��= 6+�:l�v�F"O2u�U++P��j	�hŮ��"Op\1l�N��}�B�
~R�"O 1��뚀E�ĸ8�N������ "O�d��ip�@�%m�6�U�"O�� ��%B���Q��0i?څ"�"OX����ڐc.��X4-�G2� �"O��t�L��Z�lٗ{�q��',-"� ݃b9���ΎX^p��'Dl8� �ݍ2C�lJ�������'�:����ֲf�B��E��<��գ�'����Q�3�F!U��;����'�j�)���6�<�"_"��@��'q!Bg��?|��d��U��H#�'���@�O��v�cD���R,�'�Z�"��|_.��7�PLjb�
�'��`-��Y���KgM�Aiji�'}��:@̊6+.(�f�L�
댼B�')pH�s&�$/-�DI@1
�Ԭ��'a ��`�I�}����A�J���
�'t���eE�:1�$\+TR0CK�k
�'�:p;�G�j��D� #��{���	�'w�qb��2D�^���΂\���
�'�b��UGcƭB�FӕN_4���'Y
4Ċ;S9l��BI�B�8P
�'�z�c���� yb��ҕf$Rl
�'�x�
0L9U[X M��Hx80�'%r=�u��!_S�@�3((T���#�'�^�y�
#}*�Ȁ�Ix%D%�'�*PJ &��-�c@fݠ0�'m@�#p7�b�R�ѐb"�@@�'�\K�#��2�.�	��V�`���	�'I���ܪe�4I)Ҥ��h�	�'"r��b�?Vr*�rE��bY�a�'���#v���j��qe���	�'T��(eٵc����`�+ҘP#�'T.ٷ�&�4i���\�2 :�'�ژ(��Y"^H T�0Y���
�'���: ��
6���XAS�;���
�'�j(�T/L!и�pH�	D� ���'q8�'��N�RP��� {���)�'�$� �Oӷ�U�&�}��i�o9D�dq� �N	�p�� �����,D�	��E�o����a�/?���U�)D�����
I�bm����9�����G$D��i�l������:~���
0D���gJ��􃗣�.Y<� uh>D�d�7�J
M��!ѯ�8T5��'D���P-U
���"�R��.���8D�P�d΂ 0i�lY��Q�1��m��"3D�@i�Ȅ����2����+!M��'?D��8E���Du�(�Q�K�0](G�/D��x5��@x~P�F͟&�@��K-D��A@�&�0l�ANV3g?�C!D�  FOY�M�F�ӥ��r@��S�/D��QUE��U���C��_�=f(rN(D���aK�G�n�9�=4Hє`6D�0��G,(n����g�����T�!�$ٿ	�H{&���16B�kA�!S�!�D��l��Q�cĭlxT0W�H;�!����%��BV�<x-X�� s:!�$Ŝ>����60�}p��V�XY!�N�O8@Kc#>)���c�I)�!�� N= �ϟ+�i���� Rr���p"O�Z��D�{�n��U�	�?�VH�"O�	�r(q�>�[�&�?Pv��1Ǔ��2�u�K�.���a?<O��8�(M�4�`�4�R([�p`9d"OvpӉ���csk\>�~(S!"O������,D�tЄ�W�;����u"OFQ)wL�&Iz�TpJF/G�f��q"O� !&D�Fl�uK��o��-��"OXؘc�EH,hᑢ�46~H�8A"O�d#f�P�F��tzGJ:N,	�c"O8���O�#cp�!��鎧��T�S"O�d3'A��8&\�� z�AT"O
T�/��B<p��&Ƒ+H�T�c"O�!*�-�px�13U >�0]�F"O }�5!����Z�xLܛD"O��b��*I��DK��>R�JAc�"O�I�V��e�l��"P5|`���"O$��7ûg���Iw@��t���"Oh쓀EV�I� &	�d����"O�)s/��h�*��$'���"Oi�0B��gh (VD������T"O �A��A�����M!};4�1�"O��@��sx�����Ի=?���%"O�Z����llZ ���%j�jW"O�!���X�$�(C�L�D{J(:�"O�Q�h�$��+�� _r�up"O�QK��RGj�|�N��uZL��"O���6�چB9�A�f�y@�I#�"O6Y� ײh���uhXYB%��"O]�"fY�C�����EB�AA���"O�!���(�X�2"�,�9��"OԤz�f�>M�`���P�ML]R"O���J�IuЈ��!�>�+k�<��Q�4P 3��� c��i�P|�<�V �Uu-<�Д��C�<���L�pq��s�gC�� Y��C�i�<�v��e�����E�q�D�J��c�<!@�Oh���P�#�4G����G�e�<!5�٬0�4�v�Y50~���!�l�<�!���|� �&̊m����F��]�<�c��S6��+c��.,�4�����<�(��0$R����*:�Ν�PGe�<�@\!CVIѣZJ��8�+IV�<�F���y	$-�F�]�A���(�Y�<�v.�+\gFhs�I~lJ-���T�<i�-�Y��K���]����Td�v�<I���>
�����~fP���L|�<	c���2I��^R3lѰ���n�<	�a�Q,��c��|� �0Əh�<�4��&�$�h�H�(J�:\�u-V~�<������`q"f��?�����Ky�<�ƃZ�=���/ľta�ѡ ��v�<�Ǭ 5?ؼr'�B?��IЇH�<��$�~�l�i��0>p0J5g�k�<��b\��	���,	�bt�!�Dd�<���CvJ���
��-���p�J�<�&�T�;N�q� Z3�
ɨ媙a�<Q�
�h��yxv%r��h�+�^�<�Q��M/P���j�.S�<��	^H�i�v��//,�:��L�<�j�6h���;Dh�JRfhR���p�<�ա]�}] �2��
��|d
�d�<Ya��4~�N�*p	P�`E:���N\�<��Y� �d��ܐ�Y�r�Z�<� �!KCIŉx��Ťߺ;Q�9"O�1j����xdIӄ[�� "O��g�<aPm[V�0r���W"Oj8�EN�3PЍ÷����`���"O5��
�_Z�d*1&��}뒑��"O&�ڄ)�\Q�7��4t|Q"O� :�M&ޘsi	�Nh�!�3"O�(�"W~�=v&ؗL��+�"O�T�U˝*{�[�%��?"2��"O.%�W@�0=��-9�$��!�Ƞ�"Or��0�U����ɞ�t����"O�@�W�)L-����	��i�����"O�X�G#x3�%˥FY#rh��"O�!S`��T¦��deb1�C"Oz�[��0)\Ds	Et|q5"O������s����V$�@"O8�
#ۨl��֗3���:e"O�ay�c�3FJ��0�a��ZĈ��@"O�9���2�=	�/����d;f"Ojm�C+���(Y ӭ�5�:�#�"O��z��бT��	W�V�L�l�b"O��ҷ���'���6n��"O���f�\��A�DF5A��s"O*���AQ�?'nԓG�J?8���S"O&EAv�͡MbQZ��`���"O6����:
�a`@�	U�u"Ǒ��M�+�~�S#���:� �X�"O&QK�Ȇ�&߼�Y�fI�%o�!� "O>��c�R���t��*0b�Pb"Ot�鷏��M����BH���@�"O(��V鈧	p���21A�4� "O��{��#W"�<����^̤R "O8͛�*dj���c�÷�t��"O��c�,��$�.�I�Q"O�H!�.�� 7�b�y$g�<�!��;wP��I�o���³C��N�!���<�R��&�np5�6HJ�0!��4j}੘g隹^]�A�;8!�Au!6�"Fm�ظ�ɇ!�� ]9�ܺ�É�Up=���r!�<D�Ga^�1�P��Q�U�!�d]	+�N�	`�\�����!,�-CS!�,(t�a���Fq�d,��:#!�è&\��' D(��MQ䍙�|�!�D<7����I)pfةDB	�!�Ğ��(}�t�5f�������R�!�D]%]��2�RoѲlp��W;$�!�d��l��È���r�@��/�!��o��IĨF-�R`r�A17�!��F&u��m�5�ͥY��{���$�!���s���͘)
�~I ČW�E~!��V9Vc`�;��G�Fj^�S$%L�u�!�d�	�D�8��Y^b2���F��b�!�dZ;&S|��1#�GC*M2�V!򄁎d#�٣��,7(\��V���<!�>=�jLX$���d�\7!��W�zQbx`�"�8xl1C�`[�:��'�ўb?���G�X����W'� �(�s�"2D�(�c��/*���!� � :8��O.D� �3�'Gw8M2��߆eJ���@*D����jϮD��=�f��BD��J5D����oH
��ab�	D�\��i?D����j����Ǆ�B��A��J<D�Xqr↕P(Tщ�{�āCQ�;D�� @�h�A̮��i�'��3�N��w"O�p� A�1�XB�'��:��0�"O�I�(, 2؟rd����"O�I9K\ g��1 MR�&v<���"O��q��K��I��F8i_�D��"O�h9���d��H�~�Z�b�"OdY�̢n���6d�`��p8r"O��Sg�ɨ�E�r���A�"O��c��߉^�D�f��e��}�B"O�� ��ЬeʺՁ�@��I `Q#"O�%XJ¿ ׼�� o�2n��p"O��儃�*�� ���Y���)�"O2�93�&W�����F����P"O�P�K��U@%�q�8�6��S"O�E���۲X�25z-L�/�.��"O�
S)�=8�lh� �ڜY��"OB"�cH�"h��e/�|IE"O\�PT�Fz��Ijɒ0�. �"OڠC&㊚BlFGF�5��8��"O��B`�Q�O$���c��|!�"O@P�4�F�D3"�D��;u"O��6JQ�C��!� �%U�HUѓ"O�M����7i�u��@3Fm��q"O<M*��Y=Tz��=�&��"O^��Ξ�rn(	���8G�d@sR"Ob�8�Ǉ't�*�j��9��4!�"O� /UL �"́�@Є���n���y�h��e��: 05��dh����y�+�HB��cU��1��D�f����yշ/�,�`F�uT��%� ,�y�RV�t܋B���h�t�Ц��)�yr I;:7ڤs`�oyp����K*�yB��x��g�0�AE� *�y�LF�A��X���^�N0��[��yR��v�I��CYB�xȇ���y�ޓ6��y�eϩG��)��_��y�ۡ�ƌ{�#�Oײ���D��yRm��HPq󢢀�OS����.Y?�y��-f�|�R
�W�!zB�� �ybhK!C�� ��_c���H"ˍ��yr��%w����-C�D��a��+�y2'ҭ
:����7�x�*����y�Ȼ6B���J�5,�p��-�y�o=l�@����
fo!q`F;�y��"dM�p#R Ѷd;�=p�)J�y"ib��X!���E�DM�tcҢ�y҇�"un�+fV,��I�(M�yB�R*I|r�X��B#\`����*��y"�^�s(�1���P�bxY�%X�y��ͳb�ItBاK�����ED��yg�X�P�Z�A3@��y��;�y�D�*AS~�����5�آ6�y�k��$�"q!��ؼ{j�s3�_��yR��2�#q� � e���kU��y�"��M���V��5.�,�`"��-�yRaR
[��M0��#���Q��y2��*s����P'4
��ae��yb��$|�P`)��:AYx���ا�yr��H�4X�C�M2��bgCS��y�ҟ'�j��R"(�`J��ҋ�y�͂������m�Jy�7̝7�y�� 8(e���(h�z'��yB�X�S�6`�`"X�Y����6�E��yR���|�p7(����p�n�
�y
� +p���_}�	ku&]��s�"Ox�XD�7-(����N!C���"O��㥥�
>�r���ƫ6v��aV"O�y��A/�`��&#�ĉ�"O d)�J@�g�X�R��Y>���"Ol)��	څ�,�� �Nn ڰ"O�����ƕf��:L՞(�����"O���԰i�
�\�������#�y�jIg���h���$�x3�'/�y��r�hQv�N�q�
P&�V��yB/W+S�vئ\�}F�4*��T�y§��z�q�o�:F�~�{�\�yBl�3 ��ˆ&�@��������y��O��I�5m1,:ԁ��y��1l7����)��e}�	��(��yrj��QV�%a	7]�"�h�J���ybĐT*���ڈW�[��3�yBC�cFr��RdWWe�ESa���yRC�.U
�"���le3��H"�y�6��,���#	>XT���y��J>�cգE�,��i�<�y�<3ш���ٍw�j�A0	�	�y2���[��y`IB�m��X��`Ҷ�y"+�*Y�9��Ll�ZU��L�"�y�� j��4�pb3`�.�"�� ��yf��^6��:�"��I(p,j�P�yRm �5��U1U�]�H�P��`&_��y�m�i�Z��̇�u
��@ރ�y��ق%5�����دmT4�#�LC�ybm��ܐ��*U�f�.<��)�yrI� Eo]�7a)X���Է�yr��~Y��p�DQ(�P�B��y�/V �P�G�	VH����$�yb�z��xsC�¡0������y�	ň9��Ҧa8R��u��)���y��P"��X��J\(-ymƪ�yr�B(qLJ8�4ŕG� �+E,��y2ڵ��Y�
��<���W
�y"�O9J � ��X-��A�.�yB���v� �!��y�P�����y"WB
����7t,,dPFJH��yB��8f�)���݀f������yb�H�8^@ D�̖ear�ti�,�y�'D� �bt�r��k�(�@�g�%�yB��'7bIp�vp�p2-ϓ�y��S�<�JA�t�T���\��y2�P 37� �s0d̓Rʈ��yb�W,3d��Ӂ�$A�4q&@��y�"�^f��y��K��������:�y���34"Jѐ�dV��v�#Uj���y*��GR�����A
{l��4#�3�yY<w  %�ǧj�1��!=�y"�_�T�v���mT2�zi�fh���y!��Ms���/N^lX���yb-�)Fr���ӊ?Z)kt́�y�M�?D�ui���2�H�S���y��%F8�P��
 .�Ik���(�yR��L��ѹw�ѧxÆ�]����^A���JK�wo41C��Ѱs�ʌ��1�j��tĆ�@��ԫ�ZZvp��4j��toR�^m}���\#�t�ȓiyp��$L��[�"- CԔW�\M�ȓ@�����<��������D��A�Zt�2O�0z�N��?TT��S�? �Y�G�P=�(i舁&բ��"O���b���S�~x��'�%s��Mҗ"OJ�`���1��`)�Z�:�|̹6"O8Y`/^"=�`���ƈ#�v��T"O��Jr`�87���d�H^ꝳ�"On��v���G����b�̐LLd�"O����U���KX�l3\A�"OhH��V/���kJ�Ɩ99�"O����J^®� �ME�g�Ʉ�K���ҁ���:����l�v�f%�ȓG��i4K�tQW�Q��ȓX<<���_�|�Z�`@*���p��~d��iF�m�`�M�$`.� ��9n�5!FFB�i�ݡ�+�u䴄ȓ X�h[eO;zx���[�Y�.��xF��sAD�(�2L�TeZ1���ȓb����-��jaP�IW� �O�U��.��X6M�'YK�\��+��eI�<��J�ұ�EfS�Y�a�yjx؇ȓn����� \�A��aDP�|@\��ȓE�h`eF�% �\�qq�U�b�����o��I5呶ox�T�2�o-�T��$ �AP�E����^Y�@��ȓDzZ����fK&�G��A���ȓ@����q/�{e~��T+ކO�J���yU��i��(����B���'ў"|�0N��v�By&a��c:���z�<ag�}P.�D�W���=C�H�Q�<�0D�?-�ChD�!%\p��
M�<鶇ԋ%h)��B�R��:�Dp�<	1�X<����bN�7zQ(�I�h�<a)�.0H4�r
�(�#���d�<)wL%&���+����W�t��!B�a�<�u�^��]їI�do�47��r�<a0fp���7���W��d�KSy�<�W!ݞX�H8a�,1"}$��r�<�@OJ�	����nV���]��/�o�<����R�ȓ���s��x4�Jh�<���O"p!��ɖt�qA�b�J�<�2�� A�$�"5�	}��X��C�<Y���%@bM�WN�+H"b�ׂ�u�<��Bӟe�����"��8CΝn�<��%Q=ӆ��teT%Z��&ea�<"��+?k���t�ˈ)5��C�*c�L���,�3�t�j���{&�B�	�6��`e)��?�<|{��\*|��C�I]J*d��(Y8"���x��C�	K�t�Ӌ�b_�	('��I/tC��:Y�&�J�섋�c_ge�C�I�vU2փ
�L��[?x��C�5&�L	�w݊gh��@���6-C�"%Z
ųB�V!`K� c̃�h�B�6���pq�X$R..ؐ��݈H?�B�I�.��p8��	:Rde�gg�fҔB�	��Du���+[ U�X9weC�	�uP�m	��f�T���B�I��z���f��&c:��b��B�	�)�L���̰.�bh�� ^��NC�	�m\�X���*�( :�`�6�.C�I;��x��L"���%kf�C�	-�L��wK�4.|��Ia#E�b��C�	�^��<���^ c��
Ī)ĨC�	<-�d(��ǌ�b��,0Ʈ�#�C�	�T	:l��kץtx�uɒ��@f�C�)� (�[�O�5/�`3�ÉG�J���"O6�*@��Nu�1	������T"O�cU��u\Њ���+�XX�1"O�4�7'��9haW�+�A�p"O��9v%�5𤰱#�,	�6Uæ"O�,�u+��xX�ա(��h"O�)A��Ԭ!`��\[b��P"O|�jVl[�qF��jPe�?2?�)�"O�]d��%H��1�$Wk(�I�4"O �ѕ��'0���bз:�r�"O9A��� N&�	w!�C����"O.1��"Nt�z�� F�)���:�"O�	1e�ݤ���s�%���0[�"OZ�+��������ӛ<�Yi�"O^��m^�A9F����G�:_@��d"OPI)�,ˇh�
�K¤ʵ_N�PP"O��b�/Q %\m��F9-4��QD"O8,�BdB>��i .���5"O�J��O?��cf�8{����D"Oޕ é�<9�Š7"([���"OT�ҁ��K�쀺c��Y�y15"O D���UA%&�1��"܊DK�"O:8`Q�W8�v,��kɀ+�q��"O`�'��Ld�,��I;
�(�"O��0�R�8��%I£ٚ`G6A�"O�ͰG�[ ���GB 0K<2��G"O��e6����1V�dJ�"O��E	N�\p%GC�+<|\Kt"O�H�Piʩi�<)@�ʨ�ۢ"OZM��lB�7Z
�{pH�-p����"O�%�`nޱ*���3��4g�����"OP�&�)fsD� '�L�@h�%"O ���2�j(����M�����"O��[��
.M���k����ԛ�"O*u�Wh��pM��GU*G��}`�"O�Hu���OG���gg��ZT����"O�Q�e��C�0XI'&�.T~9"O���BLN6+
Q��=|��5�a"O�u�Dς��4�rE)�b���"O�0�P/P�u��Ě�c	�h)�!"OPE�%j(�Q3"i�=Q$�s0"O��1Iܰ,�6Zf�y�� �U"O��;! P�ِm�C��.�D 03"OdAŗH6۴�խR� �"O��iRΓN����� �kmNh�t"O:-⅍L������.��"O���'�(�+��ީg�b%;P"O�Li0"_�r�%5�)C�`�"O,Eh�O�X>驰*M�+��)�"O���Ǫ��Cv��r>�izs"OrQ��Eɒ�*�ѠKU�@َ��&"O���;=��E��F���G"O�x�%&%Z�̑�I�����~�<	��W(Z3�h6��Rx���Æ}�<���>�$\�����F�n��+�|�<�eBĪ,>�����vlf�#H`�<���F�{G��H9��Ń�S_�<���Ғ� ��A�O�0������d�<ٰ���PH�H�+2l���ڧ`�H�<��N�E���*��ҵ[�BM��<QW-؂;���0s�-t��+7a�S�<y�E���m^,c-�嫳	�D�<�鞥'sVp{Vf��I�n��6�X�<�gkK� ~�|0.�:��}�"b�_�<� �1C�h���$�*�M 1W�p���"OV�S�Cz�D�w�g�N}J�"O��&�޷��{�fώ4t�2"O�ݳs���8�T���!*8ɺ0"O���ъƠV��[1k�9L�8�v"O8`yB���6-�`��<-�q"O��%� =n��ț4)�B_@�t"O����í���Jq��?@�I!d"Ov͹�K�7x��y�®�&W!�Y�"O$�!�ճyVX)�-٣rzb�3"O�H�h�(7=�x�dAN.�s��O��k�ʇ��M��O?�	(}��4���O�R��ږ���~����G?I�&�P��8_S�u`���I�b�>����M�N������*&��AK�i!)���T_���Cb�(h���Ѡ�o\F����՟4?���c���?M�TѴ(-΀8p�M��ꧩ�O��d9?�{��M��6i��y駈K%5��h%�]|?���°>��"ϟ�>�"Pl���b�+�B8?���y"�v�6�$;����m�2+H�eh�g�Dp�l#1b�&����mZIX����(QɆDv�_E�! �Ö�\�BYSV�ɜXR�a�6B��rU�����Q�D"<a�,�)$&F%��a�:"u`�'C�0<�2��䓁.ޭ*��,u6�a�O��tIcHي	d��hu���5⟜6�Z�ȇh�2-��pN��?)��?��]���gy��'��	�w``c��Bli�@iу=0���D,ғA�#gI����Ҥ�ɓdv9TN~����5�d�.�D�<�F�ϫǂ%��ė�O8�Y��?_wh�B��V���<Q��_5�c�V:l+<!��%�ĮQ�"B)<��D��{4�xb�ʖ�1C�"?�
ܼ`��@���	���@B�(��Q����:�� #1�i,J���cCRh�VW�O��P�'����Q�U�_��y"��v�*�����J7��O4��?��*�>�P��^�q �52��M\�$��S�LH<���=<z��eэ;n�(�d�Y?��jf	zܴ��ě�5fډ���?����X-a��D/O ���7��So�5��Q��Iԟ�� ��/����[2zU`��$FX2d�)��K�za�c���]�Fl�2պ00����⯂�~�ny0�`�iW6ܐ�M�/�.�b�IG7Q�1���Us��#G�	퐸��П�ē������۴�?a��*�1A%P��#�*1�p�Ag�ߟ�?E���H���̹}u�	be��&)n�0��)�S��M;Vӟ�-x�
��S����d�4B��O<��S���m�	yʟ�Ox�e��(�*eiխ��q5���y��DS����e��\HD�!;�-x��I��G._�@�X�2g&4͚IXQK��M[�߷6*ۧ��*3X���s���uL�����*V�\c{@yE,�1e|le���<��Pڴn��%����Z��i�(�
��ļ_F���ubN-M� l:�'-�'�d��a'x�9�M�EDM���d즁�IB���Mũڮ��5��+T������텍Q���'s4t��	� =���'�2�'����M��y�-R�H_�p��b�GѼ��=0k��q�&5��
 _����Oٸ�Gx�@N2����`� An�H3D�e*��R��4AchG�I w |�	��x�在 <�-����<��bR�TI� i�&yJ�9�))��O�&�b�'�6����D�O��n�%�(P�9������{��І�`�'�@HEM^9���Ң�pCLQ�_˦��4��|Q����䓙5�FL<# |  �   -   Ĵ���	��Z�Zv��9/���3��H�ݴ���qe"�$�6@; <r�il��aDx!Ei��K��+uň);��6��ΦA��4H�{�*S�.��LZA���A��5�̴��D��O(I��48���Uɂ�;��`�F,^e�R͕'�ڥ�۱:-��
,O�pI�o�s�꘠[������"�v<�F��"�@�	�K:�h)Sl�C?��'}8ّA��W��'Xj�@!�� ���EϝK^�Ը���hdpDx��}�'\lΓf=\D�E��.���q�I��p}��%�0r�+F��'�&]��@�N��h�fQ�-6�5h�' �Dx�j��'�Z�+QeI�|���f"��.�n���,�&"<Aڪ>�7� 9����c*�gx~L��M�O�$K�Oeq�{2�`�����]
�>�(W� �M�,/O|"<a���2/(iӠBA�4r ��#L��>A�c?"H��o�j�H�GN�P��m���X.R��͖'�BAEx�ȘW�k6+ӡ�]������	��ʶ�,�)�(#<�!��O���Ԡ^�.F����M�M��4���dR�O,L�L<A�TU�8s��6DV�r���G?q�%&*�LO��98[$"�8�f�c�C�9ϼ��q�_�$�"a��i��?-��I�E㟎�R��8�N� �@�]��}ʖſ<�G���;�D�'�,H��K�8�tO����L1;轰��K	��� ^�tڱ�ɾN���R�+�x��h�oǇbhje#�B<D�����   ��ƊI�X�8��%�<��i4���R�'��'y�O�A�1�`����d�#F�����?�����Şa$���C֨X�K��,�ه�>�ȁ�\~y�g�$|o|��,r��'n��A��|3v�
����r�\&B����럔�IߟP�i>��'L�6���ys"�dҏF=��ᶁ¸;P����f,Y$��Xަu�?�2W�����X��\�^��3��AF�� ��P��u��ȦI�'�B��6!��?��}��ּ�Z���1��3kZ�����?��?���?Y����O��3���
mq� Y������W���I9�M3�jE�|��sA��|b'[Q�!l�*= 9��.k~�'�������ݹt��֓���6ÜRX��ϖ�M���'��!��O��O���|"��?Y��N��u��j�u�jY~Ah����?9*O��m-b���џ��	~�d
���+Q��g8��P�Ϲ��D_}R�'�r�|ʟJ��
0��y�qH���DU�S����M��W֦�+O�Z�~��|K�u��B���Vs��Pr耥�"�'��'���4U�R�4�TY1�쟯�Z��\)(��@0����?��˛f��Vp}b�';����ȃ S8��w���T$�� ��'�Bیn��枟�:�%ȑ����~��a��l\�!cF�8r
��2���<�.O����O:��O��D�O6ʧL���02͇:���[�Ƙn��9@Ÿi
���W�D�Ig���,�����
��E��B�3�b]��Ņ	�?y���S�'0����ٴ�y�\�t�p�Wě�p�||��FV��yR�|W�%�I�9&�'Q��ɟ8�	�4
�Y�RۖIPG�t����Iʟ���ޟ��'7���u����?�TdJ�6#���շ0��)����'R�꓆?�����~�]�D�	�G\:���ć�`���'���x�e��6�tE�4£�'?hQc��	>xL����n�=�4��'���'��'m�>�6QVt�3��r���p �ԻBv�P�	��M�g�3�?q��'����4��+'�'����D
L���Q�>O����O���Ϟ��7�&?�ϻNl��ӭ83 TR'�G(8�)x�Nݻ\�'�,�'���'�r�'�2�'sέ��������pH(2�V��B�4hr�S��?���䧵?��%ºbrx�6(Q�1�"Q���2R��՟���Y�)擋"�]JD��~�\���A�v�E	�gK�D�R�w3L,��Oȥ*J>)*O�i�эC��e� @����H�e�OD��O����O�)�<A��i:d���'�ޕ�ٮ&�.�
 O��Q,!�'f�7M9�I<��D�O����Ol�8�.�5)g�A0j�1E�5;�H6--?)2D�\#��)$�S���$�M��0�g8i����Cf�P���L����(��ҟ��aB5D���fd߶N:�qE%Y��?q��?I��i��)��O���i�X�O���V>b {"m�'I.�V�!�d�O��4�&ԣǦl�*�Ӻs�� l�ӭ�r��ܣPK�u�j��VLB�?q��'��<����?���?B�31�]��,Pb EJ���?����[Цe:ƮLy��'���X�6 x��_0( >y�w���F�+Z��şp��B�)jBaҌSp�i��F�26]������&�� ��;�McDR��S�`���-�����LI�$KZg�� h��K�9����O���O���ɯ<!��i�愢�O@�p y+��:\��:u��
�"�'|7�"��!����O6`���q�m�,z�B}�j�O���	�6M;?�ˆ`x��Szy���>:ȉ[ %J�c����#̾�y�S����ʟ��	˟��	��x�OT�X����s�0�P�F=Sq�] pBs���ye��O����O(��������]�c(xHIw��_ǒ�*��Rb>�������%�b>��t����i�1?>h�`L�O0�9�Gڝk��m͓	�`�xt��O�ݱN>Y,O��ObQ�����M���it�M>�ZѸ#+�O&���O����<!�iiDd3��'���'W�ɳ�1[d��"V��&b�r0��N}��'$қ|�EԿ�̉� "C)V�BQ#B���dD�E���F@eӼc>�1"�O���P$!��m "+�4m�^��}��1�A�'�"�'{��'��>��%)���k�G�3d�}�0�^/~�i�ɴ�MK@�	<�?��� X�&�4��iD�Ƌ)��P��ͪ,�f�C�=O��d�O����<!�:7m,?a�*ø��=mT���k˂.��!�gO� Ff�&�(�'���'>��'���'��`+���o9U�� Ԏo"�k�\� �ݴ+��}��?1����O����`�Ѻ�������n�,	��>a������O�)��&z0T1)�&�~,dlC�ڔr�0}��W����F�kV�iVL�Sy"��C���kR��q�6��Wd�=ce�'���'e�O��I��M��LԱ�?�eG6��Xa�ӌ2��)-}�\牬�MS�R"�>)��?���h�:�䔛&,�`�aW�[̤e
&-�MK�Ol1��*�(����X8�s�d�1�Ck��)��O���O����O��'�S�i�� T��3
,���R7�U�I�����R�g�E�'YP6�+��s���9q�Ί�qр�D���OV��O��;�P6�*?�;^��8zG�� ��P�c���gӒ�F�#�?q��'�d�<����?y��?�拤IX�:�	<G��0ڰ�?����dF��hGg�������O�D�v�ÑN�D8���cĦ�z�O��'�B�'Uɧ���(��� � l��8�FE�2#Z�b�� l�7�Ey�Oqi���_t���c�W NuJ����!�jq@���?����?��S�'���qYQ��T���1&	�D� "�7MP�A��'dr�a�4⟀;�O�$�?,����#ݾ#m���׺.���$�O~�d@cӴ�|ep��o�?��'^$�����t��9�r蕬���q�'
�៬��؟H����x��c���Biz.�$ C'ք� ��<t�L6M
(j� ���O��d7���O�4nzީ��c�2~�.���OF/T�n��Ā��,��{�)�S4RZ��lZ�<��dG~J�a�f�M(�l��<��dw�ă>����4���d<_�L�#�҆���" ���O����O�˓lf��Nr�'��o3$ʮ���׏qT�吪��O�5�'
��'u�'TVI�%�,��� ��mט���Ozyi�!H�|�n19��	
*�?i��O��
��+�@�I7���fy�	Z���O>�d�O���O��}b��o�����ͅ�"�6\����Yu2���G�Vf	kb�'HH7�0�i��F�֊9����Θ�(qL�3�d���I�� �I��*dl�|~�(J����'n�`XX6
L�p���҂4t1�L>�)O(��OV���O����O��˂��"�P���T�Q	aQN�<ɔ�i��2�'�r�'����
s��'j6AJB`p-*�F%l�j� �³>��������'�B́Z0Dሥ�0ZA�(�X H�
Y8nRD��'V���f#)e����J�Ihy��&sȘ�O��� �d�'e(��'�"�'��O$�ɬ�M�D��2�?q��E8�����J?z_�6n�0�?Y��i��O�T�'t2��y��M-�����=w��S
�b�R)�i��	)Hx�iqdןh������QȂ5��C��S�����T���O���O���O��S�'	���@�H�Y��ak��A��İ��?��l_�f'Ө����'$�7�;��4���c%� Z�*��W)�D1O*�$�<�S����M��O�\��O�(][� �%H���'	Y�s�t����_�V�Op��?����?��\j
�YH�'C�u�N�V������?Q+O�m,-{�T�I۟���L�D�_�?�h��F��5����DG���d�}B�'��O��#,p����iS��+�Q�.9b������f�oy�O->|����'J �(��?~����H0�V�[��'���'�"���O����Mc�l�x�\��d���8/�YY��:2�<����?QW�i��O���'�R�ǻEi�Z�GI7�@� !�� ~5��'`i�@�Ig���[�f	�?�����i���3�|�0�ʛ�L��1O�ʓ�?����?i���?1����iߑ^z�h���,�0ai�"b��m�qՂ���ݟ<�	��ݟP����͘�)�z1 4��X��Q�c$D��?����S�'����4�y
� ��◃8��a����������5OLa ,_��?)q�?��<ͧ�?�CD
+o����M��f�qRS��?a���?�����צ��% Dğ���ş��`+ѾY����� �+*7��8��l�Qm��֟��j�ɑ5,r��]�<sB���C=x��myF�h���N�
 �|��
�O 0�)�|�7��Aߎh�T�Ǎ4����P�Ug����0!��R.��HE�6"	"b�'��6M2�i�ɫ������	V�¯:�J<�F�q��I���I7酋�I�uǪ�m����>���>�j�$�.JI2�$���'7R�'(��'�"�'F�]�� V��� ��=PV����42� ��?!�����<)�e�0�HSLT5	��Ts�TyU�I���?�|�ᢎ&t�a�h��*'A��]+'#��`���'�=����͟В|�]������J���AD����I͟��I��͟�Soyb��O��y��'	|T�IM=(@�(��0V�n���'�6�(�	%��D�Or��O�a��Du���&��7M�x���ʏ�C^�6m3?�fE*u�*�	������ڤy�����@����:���<��#�BႱ��0y���#�%�����?��P ������&�� �
X�<�d�÷�ñue�=sUj[H��џ<�i>��!��i�u7X*'���RRKϣUdx�(Y8I���bb�'��'���'�"�'��'�ՙcLبWC^�� ���2��`c�'�P���4'�B����?����IL�3k��4�ɀ-�������l�ɶ����O��D1��?mc�	�=x8P�CF��
h�H���6V��E�Feᦕ���E�U?�O>	���R��Ce�� �t() ��?���?����?�|(O �oZ�l�]�"�?br�Ǆ�B�f�Tk�����=�M���>��d�&���a�)(�)�ŀ����A���?Yu�Z��MK�O,m货K
��O���GO �9��a#ޏ&���'������쟴����|��b��LF8y[�1��Ȕ(3=��k��<<�6mY�S5��?qN~���K���w) Р*١����RO@�A������'*��|���_/nܛ&1O��QB��62���#�#�n
q�5O�h#���>�~|�_�4�	؟$����1v\!k�D�R\�ђNڟ$�	����	Py�CꟜ��v�'CR�'V4�����o���V̟?Ă���d�r}��'(r�|ML<$| pGuq:��&LL��'vT�`��S�B@��#1����~�'�l�ru��p����l�HT��'��'�"�'��>%�	��H�M�[ii#���oL���	��Ms��#����ʦ��?ͻ.I:AS$L
0���c�IѶf0�`��?/O* ;��e�.�f�xm;&c�0Ac��|�h\p� ��g�!��V������O��d�O��d�O���W)�P��.N"2m�D,��B ��@P��ۯbt��'r����'�v��,N�]"�p-@�`�L(2�'�>9���?�O>�|���L-G��Cg�=ظ��Gϟ�M��cܴt7�>z�D5�7�O��O�!T85��lۢa�~%2�@عX�����?)���?���|�(Ol�lچdp��	:���('�	$0���F�!q���	��MÌr��>�����L�4٨- !-}~eAO\�S�(���-}�.�q�"}3E��`@KJ~R�;K8ܩb���z0@�)�P�>��,ϓ�?���?����?q����OJ$x�VF,��%�qDJ�o	X����'T��'q�6-�KT�ʓ ��f�|c�-.������J�-N�h�C #9�'M�������Q������� ���L@D|�N@��W�G��<C��'N5%�,����'���'J���YC#2�j �1P{ơS��'�P�(��4E���A��?�����i�/Հ	��4S�Y!)̌Im�I<��$�O��9��?�e�$����ՐO�e��ϡ&�*K\���Ԋ�l?J>A�M�C1>���&�1W��]�5 ���?����?q��?�|�,O2�oځc�<�����Q�rQqd� Ǆ� ��ܟ��I7�Ms��D�>9�xD��0������!Άd �����?�7�A��M��O
��A����X��1�M�p�,�V�vOt<�Tmc��'K2�'R��'�r�'>�=k��G��VZ��r�C*A�^3�4��8���?)����'�?��yצ^�q\�Ҧ�Ǿv�Ŋ�iߐ��'"ɧ�O�&�@��i^��W�v�ZœХ1A�B�R���U<]�3� ڒO���|���E��	ٺA8̛��>f"����?����?�,O��n�,�9�I柼�ɤl�4��Ĵ�CG���~�`�?	r_�4�����'��ۂo�Nl2sOW��B��7�(?�df����X{�/O@̧���dN �?��LL�l�I�פ�4OF$�z��^E�<�M�!b�$����|Թ5�5�?�g�i�@5�5�'�BGz����ݤ~[@]���>�D��7�H�>�r������럤��������u��H�?��Ի�P-K5�
�`��R'.lB�&���'�џXh����
���iü0��`���5?i�i����'2�'��Q�K8c��{�N4(S�AAJ�G}��'�2�|���@%�� @LH��'D�D��_�T�~�D˄q~��~a�}B��O��9M>Y)Ov�:���.�`�kW�ֿ�r��a�'��7-��'~�x�r���� s����7  ��d����?�UZ�D�I՟���;�-��V�-�V&Z<����FHS��y�'k��B�� �?m˦���N��G�Ԑe��58VڤrP��4')�(`���_r2	#�'H!a ��S�Xڄ0X䥖;$n�D�ч�>3�� eB�mz�(W���v�8I�o��]P���t~�DL*pc�CGK�$0�8+'�\�Ԣw�<b�\��l��lި��FI l[�p��H�*$�^�k��/L�c�FSr����d3Rn%�0"�+tŀ�,L�g^��`fP��H� DVn��J1g=z>��� N2=-�ea%@���XD�q�U^8r�c�'^�M����?!��^�VV�@�'�"�O|0�q�9
���k���j��X5���O]1Oz���O&��ƭf�ݚЁǌQ��}Z�D
�+VJ�m����k7�����<)�����t�ѥ`2�yX%d�x��8yp�ZW}��&
x�'���'7�W�XK�+�.o^Ȋ�f�;Ԕ��-_%�ə�O��?�J>���y�ӐVlK�4�����J���!�.�͟���䟔�'^����`>��a�o^,�P&߂BU�5��g|�&ʓ�?�K>���?A�-J��~��۔V��@��f�@{���*���O0�$�OV�DKr�"#X?����V���9��16"v��BO7ц���4�?9O>���?iLR��'����L�*y0}���8��n�����IfyR�O6x���?�����v'Y?�6�@���6���z5C�37�'+��'>� b����?�*Go�*<�𡋝-�@��b�o���i2�ՠ2�iF�'��O�@��cԉW�J�]C3GP;�B\H6 \ܦ�������4ȟ�'�����R(@Cݻ��\ހ�Za��cU�����K��i��'��Oav���$֐+�bu�*��%h�R�pd�oZ)̩�?���$�'��	��@B�6��Z�2ʐ�V�fӈ��O����.�:��'��ӟ���4�jlh��K��H���L�4��>��Э�䓫?���?�����1G�؄l� '�� di_�*�&�'C,,`�>a)O���4���Du���%�H��d��3u��@�Z�两�K�4�'���'��P�$y��3�����J�6����	�9@�h-+K<a���?AN>i-O��M \8Z���6mg6Ru|�V�'���ҟx����'�L!�o>���䘬e�k�K�	7��rpǮ>���?�I>�(O�i�O�Ab�Wh����nL�O�Z�@���V}��'\��'5剹l|�-�H|JE$ ���\�&�݈+מ��'XP��'��I��D�����'��'o�8�C�Unu�3�L?�|�m͟�	Pyr�$A�T�����k,��t���U�ʀAWEû!��'��	П�Iv�s��~�0�:�k�1�@q�7L�#���?���X=�?i���?A���/O뎗�8���`c��D0�x��dI&y̛�'�	!Y��"<%>���%�oQ�I����������od�m���O�D�O��$���S��%?`��@�Pj9��l� "U�;�O��P�)§x~�	(�.�n(�u �PlaA�i�r�'�BH�"-�)*N�P���W$y���u�X0b�/�/\�V1Fxr�/��Ο�����kGK1�z�X���7i?d�m�����GOy���~�"]�I�00ՅZ�m1fp{�$���O�1��O�˓�?q�J����K�� �l�8$���p�)O����O��<�	V?���0�n�ۅ��gB���N��	��O'?��?����$��N�L�'y��FX�>�!��G	�/S���'���'H�\� �Ig��'ǈD�'B?u�����!$�.H�C�2�D�O����<1K�'��Or"�3�L��BP� g��4�h���
q��D�O�˓�?y,���$�|j�B_�t(��#��+o� ���ќkH���':�]��yqL���'�?����F�qlm�V,_�zD�@�S�	~yb�'ҙ���uǌє���kЈE:'� ��+����Ob�x��O(�$�O��$����Ӻ�0��2_Ƃ%0�A �;�j�Ŧu�	py����O�O
��R� H+){�ha����U�`�4)�KԦM�I����?ՒJ<�'_*�8Xu�f�`�����vttE[�i��'�Ҟ|ʟ�$�O(��&E�Z�bb$�	O@����L�a��Οt�ɳ	a�`��Ob��?Y�'I�92��׻P�t�a��=+p�pݴ��2 jp�S�D�'XПf�`c���>O܌(�B�|q*��imR��Pꓶ��O��?�1�0�V<Jx��bV*��a�'�ZDٚ'���'""�'��Y����Ɨ�_R�e�&O�NfR�J�dD�?6~��Of��?i-Od���Oz����A��-�CƽT���qQ/-e=T�Y<Ov�d�O��$�O��D�<��a`�	V2T�0Sp��y_|���J�pW�Z�L��`y�'"�'!6u�'���h�.%q+$��5M��jm����O��$�O@˓8��J�^?��i�Y� l����(�B�ږ:e��	�dl�F���<!��?��XV�̓��i�����2�*�P���`h���ݴ�?������-�q�O2��'��� �����6\�<�h�KW�3:��?���?)��<������?� .YA̓�.ʌ��<.�by0�i��I�{w�9rݴ�?��?)�';��i����!c-���`k��B��V`qӾ���O�YQ1�Imܧ#A>��c��xe�����dItPl�oyش�?i���?1�'O�IIyr�ܢWp��˅�ò-���.[6I� 6M��?���O����O��?M��~�̌�D�+Vh��rA/C-�5	ߴ�?����?-+���O�ʓ�?1�'l���f��#~�����!� ��۴�?!��?!�*S�<�O �'D"[)o��Ƙ�d��mY4H�bm7��O.�c��Ez}RV����OyB��5I3���+��K��@I������ć�o)�$�<����?�����'4����8J��S���udԩ��ɒq}�_�,�Iay��'���'�p�Q�✭�D$0�g�hh��
��yB[�D�I՟(�ImyG�/`���W�R�h��[���B6�<������O����Oh�ȗ5Oȥ���c
���u�9pR��f�]}2�'���'��D��09����$�SD
��b�N**\�ӂ�K.V��nٟ��'^B�'erI��y��'V�$�>��=�$�jm��M�2����'�B]�A�M�����O������kA��uG&q�6.�0?74���ab}"�'0��'��)��'��s���'>� ����}�0��g֩1��mZdy��>DH7�O4���O����i}ZwF֕I�6JČK�KM` �4�?i��r������O��DhBD�a��0��C5r�v���4w�� �i���'���O8����$E�5*1�$��g���h0�ĠSd>m�!$���	ݟ���۟X�*��DL��H�JTe�T����p��U��i��'��&J*
Hz���$�O��Ɂ��l�R�!U�X����:F�X6m�Oh�^.0��S�d�'�2�'������H)a�b�;�H?�N<�ce�x��բ|��d�'1�I󟀕'0Zc����N1D������841\��OdD��9O�˓�?����?1/O���@+[ZlZnO�2�m�B/#����'p��ݟ��'qr�'v��ڷ�b��P��� ���/~\�؛'t��'�Z�M�����DPk^,��')���C�8�t1�F�dD��n�@y��'D����x����$��h���4)��gH��x V-ȟ����OP���O��NZV��R?��I4]*�0�.�'i;<q`��R���c�4�?i,O����O���6Z�1���ßn7�����$����d�8�Ms���?�,OJ�����w�ɟ��nL��ȶLˏvI`d� �"C��H<����?��k��<�I>)�O�-9���8���I���B��0�4���G�Ot"n�����O>�)]a~�LV���`�ӾӶ�6���M���?Y`� �<II>я��#S+�JK�'�Lъ��X�M��	J��'���'�$,)�I+��T�JI>}��S�hP�m��)�شI�&�������OOLO.�Pd�e�ZX�C@!�7��O����O2hsP �y����	r?�JX�!HvPʳf�)���[�����'���u�ϟ�'�"�'"Zc�R\�#hw�{!YJ��ش�?a� ��,�'V��'ɧ5��yك���!W�r�(͓�I���'����'�����l����`�'%�I���&�.,s�mD�l�Z@�.D��O����O(�O����O��k���i4!�8<J�`��>D������'�	����	Ο\�'.��K��{>M�ƃ�g�()ඌ��mӴ�ɺ>i��?N>a���?�����<�A����S���_���[G#�$���ܟL������'�p��s�?�B7?L$��C�6�"Yp���		n�n����&������a��䟰�O䗯6�$D��k׭k�XPh֓�MK��?�-O`y{$�[��ȟ��ӻ6.��fjW;*Qv�rC(L}P1�H<����?����<yO>i�O�N�b7�^�3�Z���̌�F/�0۴��D۷Yg�9n��	�O���Fc~�\0|�ɱM�R��H2��M��?9 ���?M>ш���M�NhR�1q��H?@��Œ0�MSB��c%���'��'����$�d�Ofu��B`�)م��:~*؂]�m3�(�?E���'**�Jg�D�m;�B���%g�H���e���D�O����'�j�$��E��N+^+���0��//��ءpIW0b'���d�I��ڟx�	��Z�h�0����>n�,���9�M���y��x�OKQ������e98pʂoZ��� ,	��'��\����ȟ��	ry¯X.sO! �[w��d"d�
}��:wJ0��O�=Y�'N�iH5f�v.�E�G�0�^9�ߴ�?a.O�D�OD���O ���7��@�(�� ��-�4�KbD��i���o�����ޟ'����^y"h��M�5��&@�Ջ����D���Cw}"�'R�'�Ip|<�O|ҴIޑ�a@�
�x�0�{��ȑ|9���'�����wN��2�h��U!J�lɱӀ���MI�i�r�'wR�'�>����'�"�' ��O�0��㥓�>�t� AJީ�j,;�3��O�˓Pb	FxZwmIE僛}������r�i�4�?y��F��X����?�*OZ�)�<�1�|��g�t�y'�	
�un��H�'~��Ê��!տOV��𷆕�ti|=�pGH��Mۃ,�?K����'B�'C��ſ>q(��}���P7X�mC�^�q5^T�F���	d�'��'�­;� ��3-*w���D�аZj|Q�i5��'�R��b2��{�D�'"�Ng-���L6(�y0A�.>���Gx2�+�	I	t��zװ`�2��O2�z��5(�bH�ȓo�t%A��ni�z�#1X��̄�	���� %�V�<9�-�u�Տ0��
WH�2\�q�
�%ah-��"�n�4��B�1�����҅$4�@J� M�A읰�?U ֍��	>!:4pԎ��'�j��2,˜W]�@AR!EY�0���)"<��ٕ��+	j�0UL؋C���I���g?~�h1��'��#���1(��0b��BȠ��O
�J%��OP�f>�ZӇ]�c�2�c��t��԰1��<M%��#E��Q+������R�u���d�2p�F4[ �а88N$#I�(3F)v�F�-`=��.S�aZ�A��	K�'1��h���?�*O�`l�7Y� ��o�nRp����,|O�q��Iԣ]p�i@��M�<�iH�O�l�u`�����12�U���wyR�,=x��?�(�8%a%��OR����7o"�J�#��1�Lȉ"�O��$P;CH Uh�		�xi�=�pM�ʧ��)��C��\���W8*,�e��.l��,[��!7�Fn����H��$��k�M�Qx�b�
!��>��������_�ON���5�{Ѫ�{�v�F��0�y��9���R���rKֵ;vl�6�0<��	�M**4B�e��	Z$R���*�,�٨O>���Oj�7M�k:���O����O��>8i\�1�`��6>���
~0Vu�B�	������b��H�@�|b�I�h��$�L�$�U�ЫC��q��JKP}B1n낝�}&����^;C�xITkӾzT�.�|�'4���|Z��D�`�p�x���,��"q'@�z!��Yy��	aGC�O"�P�u撵bt��9�HO��cyRC�x,����L�>r`��%Ќ@ZI�k�]�R�'���',ם��T���|��#Q����Þ��KR���b��p#&�*|}���'��<�Yn*}i���6���4�J=K��ц����`�j	{*vH����b@���) x.!CVL�9ۺ�C+�O���4ړ��'�x����G%��#���u��,�	�'иm�W�D$0=3��ڷn��yRK�>A.O�(Y'��j}b�'+� xf"M���$�4��n� �`A�'6b �KB��'d�)��%o�x��"�J��1)� fӔHyBД�e�v���j&
׌�p<@�T�OU�R��бl_X��ٴBlv#�U0�Aud9o�F��㉕W=��D�O�˓U�ZE���՚qrP0�c�9�y�<�d�q��	6 1P�
a'�&؆���`�� �dI��$��e�>�P�Ŵ�y2�)�u���dCA�B@�0cLQ�l�@�ȓ ��H`�	þRB�)�'�9
��}��3o��sӠ�=l��(�C�=��ɅȓZ���2�D�{lT�*�g.<�BL��/�ƩЂ�ʑP:�5C�"��6���ȓO�8&�՘I��� �AdE��ȓ;����Ļ>�z�۴I��+
V��ȓ`���c�:0���9r�R^>�	��,����xS�L�C $�͆�	)`��EW*F�z��]�\�)��je�M�2��T蔋#DX�+�ޡ��!�Ł҅ՓE:6Y��ɇ8z�Y�ȓn%�y9c+Y�Uĭҕe��?�v5�ȓLt�BK�1ŮP�fO��������V fE�Vb�-ݬ�ȓ3�$����<��"s�!4��zޜԨpc_<7�0A���!u�ن�C���fL�d~pE�&�,�X�ȓC�&�0F�d��,[�P�Yᨹ�ȓL�j��EDB�r$���u�N#
f�l�ȓh��d�*$����5a�b���Q��KA��Jp㢦�3�� ��%!�y{�$F�OP����[�jɄȓ!�x`���B�L1����#��H�ȓ("�Q�B�&J�`!���[Y�Y��j���X�	+Sj�}�����5��!<� �	æ�k���<��̈́�X%�<:��E�l��a�*T����ȓmdvq@�27(C���}O���S�? R�����<��Eŝ�U
x\""Ov���7o��x�6ř�<�3�"O����5^&eIq$�rX��"O\��hD)>=f����_$�"���"O�c�Z-!Հ��E�4"n��"Od�i��AV`"�j�NmD)ɶ"O�ث𧈤s��	v�	�pZ�̸e"O�1��.*8|B2(�>mN`�Z�"O$���;<�= �&� s�0���"O2mɧE�T�Hz5�ٻ�Eȴ"O�xz'i��u��p3%�s'����"O4�8�i�7o�<�򆤘5e TZ�"O�Ta7F�Dj�"��"O֥��I'!����-]
<��"O��w
ǂg)`�S@f
�Wa�5"OX���,�2u1*H�e��52��`�"O$��@�h92�R�=s�6�C"O�0�)z����ʗ(sxBī�"O��k���@O����&�i�h��"O`�'$R�*>���jѶ
f�drc"O�Ekb#F�s�l����$`H��@g"O	�b��y: �el�?PC��� "O�]���)<��1 픨='09B�"Oz8��BX0>#,�PcƤ3�P]�w"O.�	�̄�;"���OByV��y򉀬's�1�$N��i�J	���ۆ�yₘ^�p�ĎXbv�%�e��?�yB��)6Yx��FcUp�AF���y�G@�s@G��/�SL�(�yҬ^""Ţ��Ձ��	P���y�~���q!�OB\��"��yR䕆U�Ɓ�в>�Ah� )�*B��/����w�[�SN���s���cH�?�'ޫjQ�<TA�ýa<�xI�C�h+\���"OH�STL�^��$䊹'8�E�pQ�D(���/�qOQ>�2�$,[�E��Kx4�a- T��s��fR���&E��ٖ�|b&D����剝���J ݐ" �9q�����$�����0�l^�2�N�{v&I
9����7l�
��x� K8*C`<���#x6<	E���0<Y��K'�O����KԶz\���a�"R�0��"O����̆�cUZ%Kpk=c�:h f"O���c:���e�ɵS�6�(�"O�$P��w�69��,�!'��uq�X�����-⺜(pn��6ZqS獙:������+S��I�YEn$���İ0Y�9F�Q�c��B�	�g�`tP1C->o��D-Фcڢ<�4���ȟ���hE�e��M�!Ih&��"O2Q�.Y� ������X��+�Q�X�O��@ʂ.����:�����#@^�D��J[�����Z &�(w �2�-�(]���('�G�ǐI"�B�`K�����f�40������	K��/2ax��<`����&C@x`|��' 2�x1�P�wT(�I�vn���'>���CM�zivͱ����N ��OR��%^5 ��Cƣ�:�?sSD�2/:�qa��L��>D�`���W�1m���S�^��H��6i����JD��꤈Ǣسp���g�'Sx`�f��*7�M�[hո�����>����u��a�P��S�DA��^�U*�P� n��]*�z��P$T�j�X�yp4H�CۆW���"iȽ+y�D{bNF3|͒��0�H� It�R�Y��+�.�S@�-s��AE�L$l!��X���r�_1G.� WB
*~O�# #=nZ�(�ڵs �IB��q0G�\c����1U#�`���_�"ئ!K	�'dl�6B��qKJ�*Q�2dnH�FJ��d9���r%*@"E����ј�~���Z��
�d���Ej1.ѡch�W	�|B���	d^$��N[[�? R$��уiA�-j�*�dm�p��(]�~��<��ƒf/2�	�Ba��?�O��s��F7ɲ��Ͳ(B����P
\�p�
�&��ȱ�ՂH����O�,%i�%��G'Ӊ'D)���Bt��>ͧ)˔		�}������A0q�B��q+�^X��e"��_���$*|w�@[��At�n���0�X�0���-nNz�%G�D)����>OZٚf�E�s�reI���a�6��/�D��ѴM:�\PV� f?AT,Z�%O&l�c���:F�˧(���4M��<��S=E)�t���[v���'���0>a3̟����֥�;%"�S�j�?$B����7
K�8�Q&�(u����/���s.O��#"@����V�h#N�I���`��T\�)c�tФ�	�Nt�������S���.���ӺK�^6��q��-`9�\;� � �y�'7��jw�؛BL�-"�\���{�	Ն�X����S��J��[�Pl�D��?����4��d|�4�-O��dXv0R��H�J�zi�C�	6�&M��io�E�P���p=������a��R,h+���)q���b�O�`E�(����Ð���L'-�@�	MHV<:�T�4 [���d�|l�d�S�0B\	0�����#]���s���<	u-��2v��|ږ�Y�����h�zx�ѐ�+&��)Dz2G���D�p��%}<�iJ�3��da(�x�H�:n4�v!��s}V1�^���HʥpZ���'
�E(�m0��$A@��B�Y�6�>����$����||`cM�x� ���(1�g�S���˗-h�ܘҒ��F�3�I�A<�؀���	m�,���	+�v}�F׮@i�pRk�/\𘲶d�7N�t��N*g5����q�1@M�S{�8Pł�/rB��@�,�p�5Hݩ{��S�N�5����0ݕv�"<��Ȟty���:;[�x��6�N$ڇD#"��"�t�9�g �`Q�x��0�<�/x%�$�<`�F�Kp(��V��	R[!0^E�p��D��,�y����t�j��V�٩bf�	 T
�)Hbl,!ј����$
�s���(J���\��ԟ`4���t%�:�A��@�R20Oh�KSʚ�C�t���j��p˙�p���)@�~P謡�n�.H7���}���$�ӓ>�1)y�|�'O�T7��qD�l?����	�_��H�w�S�o�`��Ɨ�4���	v@��V���S�� �S�J\#x�'�����,��Pҏ1�PHJ3�Z�8�����	7*���b$�	*	��YI/w��特V΀p����R�xBŎ�7Z��)a�.��%�x��	0Z}ZG�Ğ"F�ĩ%鄊P����D!?��D��N�
��L ~ZL��Ď�O�	��~�� "M�p�dQ8�����lb��[��#lO�:�Ԫ6�S2�a�D�*2�8�ĊvD�O��p0!8BŤ��K���W0�����o��HGL��n�P��d�dX� ?��*G�f��ĕ8b�x5�nX*��I3b�4�ф�!��ͨц���OzQ�ѣ	[��r���&2L`�	Ƚ+r:M���@i��kF)�$6�ݹ&�ÔP��˜��.ѱP蜱e�d9AB�4u>�x8$�?O�%����H�z�
��>A�A�O�� ->�H�(��q�#<�0(Dx�'z(�S��T:$	ؕӷ.�f�|8bw��t?	@���q�ۓw@d,b����S�6���C��0V��xL�6��'�qi�S���x�V��S�E�M8�ʶ�Z�v�iʠ̞l�<eD3����ς�]�:E�)Ƅ0���:|,�8X�r��&Bډ��;3����OWfY��Ɲ;t�̇�I$[����'�~�"�k�q��q��f�9��@��+v��ISbw�i>��&�T�>�l�Ӏ(��j��-��n�<4����I�s��_��q�ʇ3q��ŘA-��\RX��'���˱�;lO��+ӆ���0CÑ*5�F8X 剣�HO�������� Nf`���G@�%\C�	"0�hqr�ɘM2pԠ��Q�x$C�Ƀ$+�٢s�؈A
B\��O�B�C䉐o��(�Bф>|����.K�B�	�|v(͸ ��9�6̘�枞��B䉿 � �%ɇ	��B0=HB�ɿ'����%����ë́J�VC䉥9��w׾.4���F��p�6C䉗oa�����wT�!s%��>C�ɵ�-{5��:7k�yh���ZC䉻d(��+4$I#�������0�B��> H�p�-Y%,�^�"�����B�	(q� x��)� "(��]]hC�I�l�X����ծ0�V"��{�PC�I]�p�+Vk�U�L4�%%3��C�I�p+jew�7M*4X�
��F3�C�)� ����¹:{�,���Qo���W"OfK�
]�*��dPB�U*_fص"O�:6m�#2D�pHv��g�|��V"O��K⃔(o20MX�/�i�t��"O6�{ �ݟ�r�.� ��P�c"OE��8s��YA�gےtc&"ORm�`�+21��l9��Y�p"OД��´s|�YcQ� V�B�c"ODi+BA�;#���x�$�^�p,��"O�@���|�<8�w
���;�"OJP@Q�гd�L:t�`�R�x�"O���2�L�1�D�[�~���s"O��7F��8F������%]�jt�W"O,� cB%*UzM�3�'c�.�Qp"O<�� *���(�1�����x�"O��"�`�'sn|Cc�^�_�����"O!i�@�'���J����o왪�"O@��G�cɢ��-#���L���y�D
;G�xy���NmŶ �'��1�yrmA�T�m��^�[E9["	��y"H�m�@���*�8�Q'�yB���
4�qA�-q�~�Y�
�!�y��� �:�x�*آgu.�P@oS��y�Z.xd��G��?)l����`�y���<Z>���^;H�8a�. �yB���<#���q��cz��hW'�ybΓ�+�0
���-W��YW�I<�y�Kލq^n-��~���Cu�
�!	�'���x�Z�2	-a�"�fi| ��'������WO��{�j&`�6��
�'�X�ꂁ�P1$���)����	�'|�A���F�i����� #ْ	S	�'�`�U #�qg ��!0�h�'��ᙇeٛD�(���,P� ��'\��r#�D��=�������'~�#�A; *�0���5F+��Z
�'K��RTh�3H.�Q���>k%0�'����m�g���x�$_�/|Ѩ	�'3� q5�T 9��!cQ�;$%��y�'H�i ���.% i������
�'˄�j�MB�,-d��.P[ Ě
�'�����%�7I�Yj�͝$�xy��'��!aQ�!1�H@;�gB�!0zT+�'SRY3���R�yE���X��'"���V�܌7�����@��h�	�']���	������b��adi;�'�Kn�*-�R���L:	�'n�k�O�5�B����o0�а	�'Jj}J���,&S���U�d�b0	�'8�ܫ�AB�$�ӐjU��a!�'PC?G�Z�C@ A~��=��'��D:�lŉws ��$��g?6"O���1'�Wϸ�J��[���U"O�3�%Z'2v��%.R:e�<9�"O���`�^ ����MM�l�$�k"O9ɥ#�r���O�!����"O��I��QV�<�wL�%�F��"O\ňƊT`]C0솘�r�I3"O�0ȁl�>Y��� Մ�4_����w"O��r��,����@FJ{����"O�p{Y�t���JEiF��f"O��H�ȊZ;�:�$����"OxQQ@Lݍ�|s����6�By�"O��Z�5!9n�	W��"H�@�� "O� 2�ɒm�
x�z�X�e^�H�~���"O�QW���~����FىS�*��V"O���B���7��2A�ۗ	��� "O���J˅kĴ�2`�.w���"O����^�.�v��VE���옠�"O|[�,J@̀k�%� b���"Or�z/5a��S�F�w��Y�"Ox4��䔟L�V]8vk72L8t"O(�jq�n�ZL�4jU6�:��G"O���C��1-���zI�-)���
"Ov\�1�N�R�H%�R⇜F�@9;w�x�)���F�G �

2�Ts�M�CD
B�	�64:�T��\��ԋ5Ɖ$+�B�ɝMWx��a�L�qM�p�n�2[��B䉝F~�q@�.�"�|�
� �9��B�	 @f6�9GiǺ3�|���)��B�'%�pV�L�QN����9VDB���ɂ P�g����矕!�$B�	;e��a�p�ь>��1�����y�B�	�%Pޙr5b�|��Y)'%B��':߈�c҈��\�6� g֘B�C�I�l��s�B2}�Djc�����B�I�0�*��s��%g���[4��ڬB�	��"��B H��`�3���C�I�&��Ix��Ю�<�3@΅�=aC�I> vfܿu�	Z�iǝ:B�ɲg����m��U�>0��P�'��C�	5�z���$�B�c���N��C�I�R���Z���D6��� �0.4�B�	�={>����[*��:��ܸC�	%U�8�S@��!O��t+��C��C�I�Nȭ��&�%{��$u��'h9�C�I6("�Lź*�~Dң��9V��C�"�IrP�7y2�@A��3�"C�k~B��-�L��l���ȶb�B�i�X�鎁|$�A��"�v2��+1"O,9*U,W�?�r%��`������"O����A�礜���h��"O	P�ݡQf�-�g2|���"Of�T'C�t�=���
U�໑"OԤi�� 2S�"L�T��[$H2�"O�� �� �|�����7�A"O��0��&+t�b�M�C�x9G"Oޑc$��-`��3�*J�X�tpx"O��W�=K�1����Oe���"Ol)Q����z\DgȈ(7n���"OJ���ρ�b}pH(HR$�4w"O¥�G� }��I���9&�r�"O�Ё�ڛs���R���{�Aʒ"O`L� '�r��q�G��k�L���"O|L��K_������R3{�e�"O��+w�Me��Q�Ӡ�;�BiA�"O��I#�N�%���@�V��i"O ���Σ.�x��/=[W�\��"O�ĸdC�a�fl�.\/E(b�q�"O�����+����FmށB�R���"OJ1���XE$`���l&�X�2a"O���.�>Y: �!�	��f.B��"O̴��� 5z,=bV�R�H�ћ�"O�Ȑ��;��s%�P����	�"OR�q����-�����I�0<�̴)�'��ɄP�ށ
Ң�gxj�3����|B�>( ڠ����o�.Q0��߅ ^B��12������r#Z�st���)��B�)� ڼ�VĢ"2p��JX�O�LdjD"Od%Y�*�U��2
ô35�pD"O"�Æw�؝ ��+��L
�"On�P3dK�v�i
�*�ؽ�"O��!����A�N��h| �*"Op�j�\;A�ݶR�~]+��'���:N��y�V�֔���בZ.�C䉉y�b��AW46A��{f�Ե	q�C�I+	:ȴ�/�(_��ya��	2�rC�ɔ�ܙ�7L@�>"�81�I�K�lC�2Wڨ�[S�ɗ0��V��E��B�	3Q�f!��]��Ҕ
��%%�B��sr��B�
p�H��NB�ZX�q�4�?~�`�Ƌz>&B䉄?�A�ࣄ�H�"�C�l��C��("vH�n��>D\)եC�YV(B䉵`��	x�G$��T�߹I��C䉛M���b�%=����v��".V�C�	�F�*��_���F��/3��[�9D���u�P9M�K��/�����-�!���k_L��s9>������ t�!�Ğ0+J
b�b�0'������2�!��0hC$��D�;ViJ=7Q�a�!�@kL�	C���Fu��)�[l!��J�,� ���׾n���� 5!�d&
ݤ\Xd�ϛwe:����=g�!�	S���0�M�O�X c�+%!��q�^�K`��k�VPQ��'+�!�7<RN��!�E(_����H�!��E|r�L͛*��H0���n�!�$*R�=������ٲ�!�!�D�!:����,�e���#t!��˞Y}r�x�JNF,y�#6`!��X/\21���˃vrPI� Y	Kl!����y��I���2�}����Di!�d�C��Ɓ��eKf�ʴ��-�!��v��������� =�!�ۨt���OٕO��A(��˗G�!�dW�c_���1��Q"�����&S�!�$ЃCM0�ЖG�!DP#Q��<�PybJ��b,�(2�˗/%Ek׎�y`�<O��@�Z��a)��y�
�<b���E�t���P��>�O$��$�ރ=��ty���
˜��"O����H��L�����+*�jB��7Ka�IuIH�#�P�!_vcLB��	d⠊V��9=t}Ri�-V0B䉠i��X1�O2�F�c���4#�C䉼9]����%�&�MiS�Y�C�	([>e��� *0���%S�Ai�7�$�S��M�%�8}Hxݩ0`ݒ)!
��s�<�����Ja��V�>U����!�D��.~�0C�=S.)jF�2�!��K'/�4h�� �%��e�7�X�p�!���+
�T��%C��3���	K�!�� �$ш(���F�њ �R�خUk!�$֊#+DQa0�\�If��5̘�m+!� .L,	jo�/Z~�p`�)3�!�D	 �P!�s�Ÿ J�<0vI؜cu!�d�(H�&iVx
�}�`�@�Hj!�׹
�r��ټ�4��ʆr[!�d�+OF��A! ��I,��i�XY!��K�rVl:#OK�&�I�F\<'!�DP5&3�IH�� �[cF�77	!�� �k�"y���(% S�(R,�i�"OH`A�CM�L�莐Mp�0"O��X1��%?�����̙�b���"ON�Cī�--��TD͓�^-�"O����\41B̴K`�yu��"O�����=Ig��bN3/p8���"O��ʆa�# �A&�W��
�''��a�W��� dK�Ѻ1	
�'c$�[���/�����HT���a�':Ҩ
U��Aθ�a&�G��%�OA�<��Z8.�qUk�.mJlU ��z�<11�#Iq*���.�.R@P!F�x�<�+F(�bI�%��z)0`�a��~�<)��N��a��Q��!���z�<�g�)G2�Xr!<>̊ Y�AFu�<Qq�A	c
�#ch�P�V�`��Vo�<�1G��&8�qb��U�<�A	��%���hQ �5`��p�l�<iEJئ{,(L�	\�L��dg�<!�B����� ���`����K_b�<�g�N%)(�1"�̟3tG��2o[�<�2�N�P(ܤR��{�@�zU#�Z�<y��������0Rw�*R@WX�<	AA\�ͨH��đ�L]n�4&�n�<�Ņ­ǘ�R��¿bL�` �c�<��ۮY��c�;vfV��`�<�a+�&v����C��u��X�e�v�<��I����8��<�(��m�<1��<���K����q3�lHF��g�<�@��}�qK�� U �vŞh�<��Eظz |�����x�l�3��`�<��V:Jc`u�r���K|��Hs@I[�<�$&��Yk��"U(����Y�<9�H��0j�2'�F�s� � �.�Q�<��E �0x���	9��=b�	K�<�7�	/d֜aA7c�j�u{��H�<�Q(�DT�C	ûcٞC��I�<!�,��S����(��)M�a�a\K�<a�N�7�D��L7�JL���II�<����7��=!�o2K�<�v�G�<�����f%2�p����D{��CC�<��P{:E3��D���"�@�<ń͎;r�Z��T #iF�j#*Bq�<馥�*+�Ģ`��Zt�b��w�<!%�\�H�@��B��v}`D���l�<)�@a<���m��q����N�<��Z{<P�B��5|���DL�c�<Qg�˾M	��ĄvcD0�t��[�<g
^���NG�n�{�r�<��aH ��(Wn�>]�&����p�<��ԯ)����R�:���ؐ�Im�<����=v�8� �&��8Eh�hKQ�<y��+��$q��2TzP���J�<9u��o��`�㍪����0%�B�<YSm�^�H�cg �-KЕy�aZd�<i�bI�O��J� �4ay'm�W�<�')�5K������ژH��Yk�<�⃏�!M��;q�D�T����h�<�6+�j�F,)t*HW��KլK\�<�#G��<�l(�.�ޔ��o�<iq�Ǔ N��iudBI��Ů�l�<�w�W�r�vi�R;R����	�\�<�V��ޡ��e��t&��C!d	S�<���	�NM�&I�/��X34��i�<� �E�7�'~@>MJ%��n�E#6"O��y�`U�2�$P>mZs"O���AӔq�|�6.Žo[��"O�C���"}<�8w̞�q�D0V"O �;�j�8��(b'�	f���T"O���ϖ,6H!h�l
L���"O5x�����K���!b���B%"O���ӂ��6 ��P���h�xs"O6X�����oZ��A�DNDW�H�"O�}�S�Q�`�,����\$���"O�S&���*���9`I�~���"O���c˗-,�IE(P���H"O�� 2aK ���#�ҩ)H"���"O&�J�$�{�PRd��,nr�"O���� !�\u�DC_/"f�"O���P�
���q��P�j"OH(FE$<�6�g��-����"O�l���j(@�ui��1�@�"O�5��F�Z�9�%h^j�	�"O��S,T�V��0��=El��" "O��b�D� m/�0bwA89���G"Oe�@�#i��F*޶k�潁�"O��# �;x��]SҨXH��D#"O����J�zٔ�SЧϼp�Ĺ�Q"OvРڛL�p�:��fz��J�"O�ƍI9�N���I��]z� �"O\��VE��Oąx��q xh�g"Or�h#B#ra���͑#���˵"Ol��c 3[z���@���_�<�7��$t���x��/8�t;�%YW�<1�C&XӀF�[���Z���\�<A����X���X0h�|�*�����]�<i�
�t���[�m��v6iS�Z�<�W��4ׄ�3�˛B����k�<�`M�B
D��F�6�.񀁇�}�<�C>%���@	�n+�p�w�<YpK���HD�@�Z�zp�9�e�[�<9��	z�|#�n/���xe��~�<R���5�hi�ݲX����o�z�<!���	<NT�^-�H�AN�v�<I!"R�~|<�2��ۧY���"Pv�<1�ǝ=i�� ��J�$��Rt��\�<y��~�5��G��b#ԨQ@ʙ\�<�!' ����:��Q�8:��Q4$�Y�<�ŪҪ ~���TJ�0�ڥ�-�Y�<��F�c�tACoñr;b�b�FU�<�q�7J��0)�-gxN�颭�Q�<ك�n�zuH�b�+0)V�� f�<QV�Y?b��A։WbBNI�b�<��ݚ4jf���K?��C�@�Z�<A�$�=��@�Z�N����Gb�<��&�Y.L�ÂS;^uL��J�r�<��%M_�|`��N����ӢMk�<1�$�,$���FKcF�"��A�<�C/-hހ��N�	8��rb�Q�<)�m�*HI��i�[�D��*Iu�<`ρ+`�v9uO�	n�
���h�h�<Y��b�F��Ӯ܋w�v=��H�f�<y�R�@Q�
���	|�1
�
c�<���F�3�{�D�q�)b�<�b��2x�l��W��2��SËw�<B!Z@��8�!��G�pY6�Jl�<�#jO�5�T1�"͆�9�HuR��Uk�<9q���o��Pb���ws��T(e�<� �,;�\�m{�,�A-*ٜK�"OVa!�o%Z�,q�Msv�p&"O^e!M�;B�I�
Ll	>�i�"Oژ:�*�p[7������"O8yw�ˏ'�6�9`ST՜��7"O4�x$K˻p���Cw$A-�` G"O���l��[���D���dHa"OD��q�}�	Bp��J��	`�"O�8*'�#N"Q*B�A<4Q"O�h����X:��A�(�*S�0�I�"O�����D��)C"��@i��"O�Y�oԴyVr5��>����"O�@� �2
�a�H�U��}Z"O$q��Iϥi���2��I��*��E"O��)�"ղg�Vl��&R!�����"O�,���N'o�t������h�0"O�����-]��{p	V�<�F9*�"O4��Kշ:Q2m
V	N8l!�ѓ"O�����N�@�����*<�""O4x�`THΞH6"ל4�Q"O���f!�
�ةj2bύ5�|Y�"O ����0Qh���Âw �m<D���We$��!6��88����,D��x�@�5Q�B�����`�� C'D��p�.
i-̘��+�_�n�rbD2D��6e؇`�ŃR�nA6�F�.D�����Q���*En�Lp�2R .D�����19Z��)�iJ�YA!+D�T��FU�z�4�7.͕���K�F)D�����(�0p2���* 砅u�)D���Q������_�V-�o-D�Б �s���+�㐙o��@�@.D���� ��8TQ���Ї wV�xC(D��p�{[��`!��#X� ��f'D��z�Кg
�m�Q�Q�<[��*5)8D���M �Z�nQ��MG��y�8ړ�0|�'��e���ƕ9(,h!��u�<�tD<~�4�H�a�)yr��l�<IB)��w�΁�r �L.��hfHSA�<��Xl���P�2]�53�A�<���?W� �lP3�=���|�<� �'~�4p���cV���#E{�<���%k�����͖��T!��y�<Wm�=4E�l��n����R�~�<ф��pm�n��:�-���F{���ݮ`� �����67�ă1�D?z��C䉨<�rm�e�Ӟeg�`�-û.zC�	kȶeׯj�z4R��bnC䉹C�IJ�U�K�p��&e�B�	L�J�P���Y~Tؑ�!�a~Ғ��zVf����eg�ya��B�9D�  ϒ�x����'A�D�2��7D�x�MX�Z<�@�@7�X,�0h)D�����G����2�C$k�h0D5D�$�'ߐ������<��5�0�3D���F#]D�L�Kcnߕ{q��ZR=�O�牵G&x*�j�S��L+�咟 o�C�	�]t���W�J)?�z0Q&���㟤��� �����"SWP�K1b����O8�=�}�U/�-%�<��OB?�xɠ@�p�<ɲ�*}��e�'j��@��x b��P�<)%��q�ʍH�<�ht`�/I�<��A�vD~�S�O�"v���b_H�<�@�-8uz��CO �bD�<� �<w�Z�z�N�4�R��$���"O��R��Y%� �e�h�������5LO��:s����v|�W��-��	�2"Od`1`�S�Z�h,+�"k��u��"OhqQ� �_N"�{�;U���P�"Ov}�P�F�sf���a�k����"OL�1FkF$[#�u�r/ˏU��q�d(�S��^�>(9���ZS@]�ڈ3��C�	�+��E�d�H�5��� -0vS~C�ɴ�ȅz��V�T򝳗���pC䉟�����]� tu'+9clC䉃&۠e����r��&,Ԋ-"B�ɰQ;�|R�k\�]��Y@VK�#[NB�����3t���T�����ľ��>��O��Z=ss,TX�m1+В͓�"O,�x3%��LP�C��w��"p�8LO4����6e019� �d��,KR"O&9��@{�l�sO�/+���"O�q�3���btb�nĝ`�n��"O�M�Cʇ�i��L�f�N�E�&��T"O8�tE��(�8�-��#�0 sr�H�l� J�@ �	.�\r��e�"D�ܸ��vu(T�8L��f6D��S�E�!�zI+v�[ EbnQї5D��r@��h5��!GC�! �`�K3D��"��q�P��J�_I��"q�֨�y� �}<Py� �H&X.�+@�]�yB	�)�hP�L��j�1N�y��|�D�h�
	�n��pF���yR��y *Q ѾnC�P#�����y�+O�0� �;�!H�`��Â(]6�y��C1:�+P�E
*#�� ��3�y¤��8ֆ��@�ףJdP�r���yrˇl�m�Q�G C`�%0Gʭ�y"QL�j|A�M\�H�̔��yMR�����*�	T�(&����'�az"�\ B���p�.@�|?b�vΊ'�y��S�;*��eѕm�]���&�y��ʛ��|��Ѿn����Q5�y�&�>m����J�>�4��d�á�y��F3��,
u��0��x��V �yR��C��I�e��&0{J�CJM.��<���d�+p6��K� ��$A���P�O�!��/.�8pC�A�͚ JFG�eC!�Y�)#vp5�"�Ұ��F�z-!��
IRU�k��C�΍�2卯 !��V��=S�^�K��)atBB�!��5�h`� E����[B��V�!�D��;��IK�J��V�4=#��L+,�!�>-ب�P#�23�����Z�p�!�Ǭ&�V1�0B�	��M�Q�,�!��Ȳ�`�����Pua�"WA�!��\p�D,�$��||��Bֵ.�!�����ИV˸%��Y;���=�!��=]D��O3A?�q�e��=[N!�G�bj�e��X$���t�ֱ+MўP��"hȎ�	;Y<p��F�4�C�I��2lI�`.:�t���Z���.�S�Oҡ�Uΐ�I���AE�3�Vx�"O�͈� [W��Ab Cf���"Oty�PY��4��!���"OTe�gźM�tBG ](K�ڑZ#"O����	�ڶ�I��2m�B���"OY����)�8���8'�Rd�"O� �M[b� Ru�;��@%ْ���P��E{������1 �2��4p6��!��M�J�es��1��@:���!�ąr���\B��i��` %�!��Б=v�%IfmG�l�=� O�Y�!�d��.|���LI\p[�nO��!�$Q�V�N-5m~��r�_U����9�$E2�,[�v7�������mG"OȜSp(O�/����Iͩ�����"O�5e,��\kTb-Xy��B"OX�P�:q���`@Mlt�� "O a����@��(qj6 {"O
����=S����$JTto5��"Oqaqh^�@9x}EH�[_<����	y�'��`��N�	)Fth�	�<&E��w�|�)�ӛf����bKӛ3�����@�Pt�B�	�,H�=Pl��D��@HuI��u�C�+�0��eY� z�S��ݾ;C�C�ɓH�(�!�,#�:A �! �jB�I2�,���_�2���G����B�I���hu�3M����'
JVB䉨���'	ՙ.�l���ڠx�T�O���d�<�6�A�+~Y��7���
!�0b�$�P�����b��R���"O�ɰm��,�XE�/P�I	a"Ol��` ��) �R�D(��5{�"O�%#  U$�}#d� �0x�0�'!��_r����Dm?���J��!��
�֘�1��(<,X1YԇE1�!�d��a��f7�6)Z�!�D�o������;Th �A�P�
a!�],�����7WՔ��e�Q� y!�$�L�t�*��ʰcXF�����gq���Ҁ	欨�d�00��0��;�B��,Aˈ�Z��[7'�<�!D�� ��B�I�9 L�!CX�X �D�ֆB䉡9�\ɨ����rw��Z�A-n`B�I��8��H�l��X�C�	^�lC�)Ue��{���y�D��7	O.k�:C��svT����_o��̔QJB�@��P��ݲ)�U��ɗI/�C�	IͬP���U�$���ł��F!YD{"���<A��Ё\B��P�'N6*`$�[T�]�E{���@2J�Ȭz�L#q&z;s���%dBB�ɣw����Hμƒ���@@�=�xB�	�?���C�/flD�qҮ�,�HB�I�J�v	��r�F�cFG�g>B�	�]XJ�D�N'����'���ڒO ���I�q�S̞�lmL�hT��Oz�=��$����6Fҽp�>��\Q"OF�9%��?m�$��C�77�����"O6�i� C7{�U�r��B��	[a"O�U)�P�D٦4rS$y���e"O>9R��.([j�p�O�?=:�PW�'`�	=� l���qlZ%��a�D�N�=	*O�#|�"�ݢ6���E���4.����B�<�1���a�>�{��X�>��a�vJF�<�2�HSʾ�E�,4k�����X�<A��'&�[0AҨ�a���YX�<��O@�b��
�y� �S��S�<�@�5W��@q�͗�v�����t���ϓ	N4Sf��ku LNa�"OZ)���[vy�Dπ�M	0mA"OB���C��7tȝ�%��k�PP�b"O� @���M�Ja�C&ھ�h"O�i��j�0h��Z�/�){"O:!���B�,��@ۑ�-B^Lr�"O�ɒB)pc4�2��#C4H�0"OB�Ko>���`��:)��!q"O�Q�ā�D���BGχC���23"O��J���;_��9� M�"�L�k�"O.��2ɍ-���Zu̌���j'"OJ���̾.)J��B���R�X�7"O��
�1U"�(�. ���0S"O<ٺ#�N&L�l��r�B v��HAc"O��:`G���A��Z	H.��"O<U�,�)P��s���1qY�R^��'ў��'o ��D�Y�W��F�P�Q,Z��'�N�x�L)lN�R5��=p���'9<�i��אS��pٔ�ɦ'�8+�'�j��Q�Y�5��w��t�'�"��Bɟ4��	R�h�rm��'{�2���=�\����\��9�
�'�9���#�v<r��H7$����'{Ԡ9�OӬL�1ЀژϘQC�'� �PQO �<��a���O��'}ܱ ,�1yj�ׄK����'� ؁n�qP�C#�A�I�'���M�>u�R����#  ��'���P�o;�9�Gˀ*P0T9�'��Y���E�a����g��'-��J�'9�P���ɐ�˗�q�
�3�'S�=�ׯ�58> �R�H�e����'NaB�h�,[F�#An>\B:=��'+�@����)���cN�M���'>6���6.�@���C�,4�4�
���`-׌X�&̓����F��Dzi.D��*��BTŠ'�B�R�l�0%.D�T�f�^�$(�Z�F��[t��XV)*D�3�WH \S�LT4!�T�ó�)D�k�K�>J{�hI��_!B`�dF&D�$1�-�;� ��n�:��u�7�#D�t�T�Y�n��4:6�Y� �1��-D��
�F�4A.�r�H�:xh��A�&)��0<����1J�;�(J+3`$�D�D�<y�Y=`����Ύ�n�B�Q�h�}�<�E�g��k2J^��͓�o�u�<yt/�zܤl��B����1I�[�<15ď%um���U�۷c�-��cFX�<���>|T��폴M?ZU�M�U�<���ф[�7f�.Ɔ-y"�(T��[ȅj�4�2k�3|p�h D�<��+��c&���:���q��9D�x�rn�;V��*�! C9T��Uh3D�(1�ڡ=ňr ̙�l�v���B2D��ZF!
+B�p%�:b�J���h3D�|��W�Fa!r��R6d��c�<a�j��OY���E�=�Z�tDv���0=��	n�xI�Čɟ?�]��H�m�<�s*��p��̘#�[;B8�c�%�j�<9c��_�ؑa�^�̩�&�TN�<9e
Ѧ4�
 �qm�"���+ZG�<�tD�%F p�bƎ�3U�zg��y�<��h�*U���B��b[J��P��zx�XFx�(W��JA
�&U�<`�#���=1�yO�wh��s�/�M��9��Z��y�̭����C��F���	��y∁�ZI�U@�F��@<��Qqb��y
� ��e�=��HH$As��"Oi"uf�4U���#��SX��!"O��J�G.4����7#V'y%��Â"O�tyJ�<It�"v��X>F����i�x�#�3"Δ1���F-h�v��g(D�Đ'�LwD�y�Q8&1C��9D��bt���i�����[����'�8D� ;�#B�h�T��QhۙU����b�5D��fK�[��υ�<Rr誃F9D�@�E���!z]37�/�F�bV"8D���uaƌc ��P�b�zl�� :D���K4>�|���P�>tBCTH=D�Tˠ�S�>H��a�� ��.�r�<�gK�_I�ȉ��V0f��m	��W�<��g0P!x����kaRh��ju��7ۂ��� ��2�Y�H
�iB��ȓ3�M�E�>N�Y����C�	���M�Ǘ;@�4��"��8�'��D{����R<k.�z1�R%l@�e	���y\3bL�2�J�"\��a��y���q�Ψ#bo&D��Ɉqn�;�y�%�E:#���6'L}� L��yd
�3X<mʑh02�q�7�P�yb�	�)a6�9e)U�$z��#�.�8�yb`�2-�t+G�F�op��X�DS��y���VsF-Iw%�#��$j�̋��y��S�'�� �tL�	:abƅ�y���/|@����Ҿg���㖸�y2)��F�V�:�,-����'eγ�y�l� aqLI+2F�0$�bAJסO��y"��0��c�ҟ��-��"���x��J!b�yy�����U0�����O���$/6�|%��D�"ust��#z�!�D��!��h����'>׌�А�	�g2!�_�s��xt��>�����&�s#!�$D8�!q#́�i�ɻ�ER8!!�$F� لd�5E��ܹq��o!�Aְ��
>��;�.�("!�D�4G�$% �� 2�Phe�0�!�$�8G�����L�OБ�3�7
�axR
�(�OH��n@<8�G`��J��0��"O�����J5��j�-ً\���3"OH��C��0���Q��W�*d�"Ob��@ ��>� `�D�>O�l���"O� qtaC�G)t)Sv#�>4�JY�P"O��ૉ]�^y+�! =M��"O��`B�P9_����t�L`���BV�'��V�0�4 5#C�
���@%���y2�Y(<0��R���0f��h���y"��k���HvOP�#�4i!#* �yrJ�"a�~1�B��E�V��э��y�n>z2��r��&D0���i	�y��L�Yp<���@:L�M�Wj\��y�%բ&w���%#/���m߶�y"�Q(��9�����ZLj&��/�y�A٣`c���B-Wrt� M��yB�͎\~ft��靚[��4J�hW��yr'@:z�P0`L�_4b��7CJ�yR��h����ZLH�*�#���y�+��X��O�p�:R�+�yG�9x��5I���a���yBc+M���X3@�]J�Lޣ��'ў�O��B�[� �B� !`�'�\M�A��|���
����<`��� ��jQ�W�n@ {5, 0�h�"O�Ic�딀f|�H8��D�B�ȹ�T"O���.F{�`�R�$޺�~\�F"O�Q*���d�j�PھeC��a�"O��&DDkF�a����Ud䘖"O�,��Ñ�`.`TY��N�f���� "OʤS�ٚg�حy�F
�� �q�"O0�3�l�K����EÂO"i��"OZ�!2
8zb�e����z��c�"O����˼gnX|{%������"O��i��!�J,{�f
�B�8qQ"O(!����Z"8�B&l�&�YG"Ot-X�)Z:y�"�7�1�2�j�"O�D����$X��Ω����"O^�GN��:���X�N4Ԁm�"O���+J��v�	"6���bB"O��`��D��̋� �o��8��'��ě��[�*��œ.,>aQ�� D���G� X���%]�/�4}�3-$D� k���<?�y��(X�L9V�,D��L�)h<Nբt�Q`�l��C� �a㴯�]}�hq.�K��B�	>y��Cw�J�4��=�U��3_H�B�	�=~����M�҈;�,k���=�	X�4�%��W�xw���`<�PN7LOBp@�.��a��i9�KY <�5P ���C�,Y�"O�pRѮV�1Jԃ�kʳI��ˤ"O��cV�q�Z]	��	f�н"O$Ĩ���.R�zdp�U9E
p�4"O�@z�	��P+�f*t(�1Qw"O�Ih�O�	F��!$�=�b��Q"O���C(V�Q�1a@3��
��'
���hj7 R(��d���D!^�Y׎=D�|2D�oҮ1��v� ��0D�L���0V�j8rSb��4���9D�p�DR�G#�ɪv$�$:�	ڲ�3D��@��O�8�H�KޱE� �b�a1�O�cبz��Y�����d$��g��D-�S�Ol
�J�[�O�l�&�̞SZn8a6"O����]E̥�5l�F�M��"O8�+([�\Q�s���#��*LO�E�dmA�g���թܕJ� yr"Opb5�ME�����B(.-�Ѳ&"O�I9bɏ�q(�A�_�~��&"O0��"�:0"�d+ŀ��Fip=�"Oʭ�phѤn�:����_�@�"d"O8��EeO蝒S.��f�0��f"O�1P�����5"��� SNӽ&�!�DI�9&�U�c["0�!�lӁ.�!�_9Cmf��fnR�q���\s!�Ċ;	��Qr���� �ϊjS��d׀O3�A��o����X�M_�5i�B�	<?�"hr�۟�Ma#&_{L$C��%tY"i��O��;��i��G"Z�BB�ɼw������(W踍Jc#��{dB�	�?8�)�W�Z�P��؋A*�PQrB�	�/��R	�r]��ˣ���T�C��/5'��iI�H��Qg>!*B�	��4)i�AJd�*��gh�_��C�I�(�10��G#T���8�gQ6 �C���Rr�&����ǅ����"O�����<6�AJ��@�f�ze�"OR�@n��^�0Kת��0THD"O�� a���:$�g(���Z�"O� Ь��NO?e%^h
�i�_�X�V"O8�ӄe��\f����)�Ai��"O��3�ǀ���㑺UO���"O���@�w�"��1%�+$�x�"O�<:��v~e���1-~���Y��D{��I%kV�D��!�]�6��D Ǐ�!�&^�:�0c^��^P$ �'p�!�����R�KXp���EO�!�D���J|��K�6�Ƹ�4�	A�џ�F���E/��@�P��Z�D��y��O($ɵ�̚G���YՌ���y�ɚV���؁n��rL�3��۰��'�ў�O�Z�@�3}p��:��O�$�Z
�'�X��D@��S8H��`H�=���#�'Rv�D"�Qj}��D�41d�s�'��0�G_� Y�a��Ƨ<�Y!�'�6� L���l�:�6���'�q)��]#G� ���薱�fP��'��@)`F�;Ib�� �%J��}��' ��JOt���ycLFrq���'��}���؂'���ؽg+6���'��Ґ�O$n�i��R�Y�J���'KU�Y0>��P�L�}n�Ҏ�D1���s@L��<Ц�sB����"O
X���S |���GDd��� ��1LO ��@��c�:}{0F�ds�� ���}�O�-�#�߿fZ~y���'�>ъ,O|��0=��&�5
@�A��T�r�����O]�<y7�́ 5J�y�g�(��x4�@�<��DMp��M=*��ȗ 0���<	���O���@���$t�A��#�(A�E"O 0`U��3T���(��� �ܠD"O���ץ�?DV8�`�R�<jP"O��9����z�ϑ�l���$-LOf�*��5^��<×�O3D��%��"O�T���1A��I'�V*��{@"OXr�ȇ� K^�0���̨1�q"Oj$� ���c�<]�B��MP,���"Oj��u�>s1�CR��/K���Q"O��;`C 2U�A�A܋{O챀��'��� )���wg����@#�"��h!�Ā�92<H�+v��t� ��_!��Ƭ	X��J���S
��e��7oo!�d��?� ��=j#��g
��
T!�����T)��R}���4i@!򄖮��uѦꏲ
g��H�!�P6!���{�!�������Ҡ�.��N'z�H�� ���Z6E���U�"ʓ�0?�ߨV�xe�I$�x�J'�W@�<YBh�#|��R��q3����R�<I�nH�}�"��M��nn\�Cd�O�<Y �_n}\�ƢȰc�-��RF�<)E"I1Aa� 	�`]�'Dbla�H�<Ɂ�4L�d�F�L�$�94�L�'џ�
�f�04U
�	>��q1��gy��'?��CdA��Rl:�(D�]'��Q��'H�)� J�'��99&,ܼLr�|�'����ٸ���sRI�5W81�(O���0=��J�'tZ���Ƀ�Ua�9z�HD�<��D�(��j ϗ
}z�	���x�<Q�W�j{^�񳡝Xl�bURzx��'=�a��N�#>t.��φCTq��"OB$3'j�zKb5*�m^�k�4J�"ON<Z�c5C�q#H�b�)��"O� :�*�ȟ�5��٣׏�a���Q"O�E8 ���:+T�Y�N�dI1�"O����4,��B�/�,u�A�y��)�S !�~�@ �� �,���8j�C��ޔ��ڿL��Y��؈��C䉖>z����Hm��2g��<�.C�	�66F c�K�LF�e�R!�PB�I-&zF���ǽhb]��P9�8ʓ�hOQ>y!�摔	ܵB�i��t�@=�d''D��ʶPV�Xe���	O����g ړ�0<�w��	&���!R��8�H�"�Q���0=��m�04��
���6r����O�<�����<�(5��"πX3&MF�<��.�#p:R[#N��[�.�Z�<y*	`ĸ:�$�Bn���V��`�<�����8�Z1ڵ�����P�[�<!�H��P%��J@�
 ��$����\���0=Ig���y=�qJ�KJ�?��Ѡ��C�<IU
A�_�P�
��_�l�z�D|�<	� �&s)�컳�Lt��`$	@M�<����O�&Lh�޽y`xd�@��P�<iW)�R�b�sB-
O?�-�P�Oy�)�'V`F�r������V�X�m�'�f���ÝHh���K����ϓ�OZX��o���ḿ.PVy�7"O�1z� �x�>�
�
Y�m鈴"OV� a-B�u�'˛�p��P7"Obĉ3!�	ˆ5��CĨ83���b"O�Ex ��k�:��◱n����'W�D��B/�;��M�C�����\p�!�$ًQ>�1g m(�K*Kx�!��
����ch�u��ԡڡ�d�>]�`"6��-A����y&��v�D�Q�$(�`���Z�y�#�oB�5�A� �R.����x�M�BK�L"���cNuHb�q"O(۵,ąWSv�Ys䉣��3"O ��QʅR��9y'������P�X� y�@�!iR5I�o�6�"��C4D��j¨X�L8l���/7�<�P�2D�x��yh1 �ʧ��ꂅ0D���ʛ�Ι[�"T/IA��7�0|Ovc�DZ�
T84�`X����}�%��,|O�b�x�A��^t I#��9΄�&D��[%�ֳsSAI�hF�3�D��$�IK���)��L���� ��(U��z�L	! W��$=�S�O���Y���d��ikp䌢5;���G"O�������b�0Qj��WJ&I�"OF	���D�,�F�3)��xB��c��'Z�ɔ-�,��˂F�$Q-��rR���&&A&�X�ŉ,-�&�InH�zt,��ȓ.]��wc� U��P��!_�X��g^ ã�vF�u(��^�W� �ȓD=�]���P�S	P!��H�^p@��m�!%&M��v��al��"�b��=��U iF�ȓR�VUK�B5 �`Ջ��Ǘ^�"1�ȓC�h��� %o��)z4�ڭo��ЅȓI�h� �"AQ��v �,<���	B�'���2�B�4Pp���	�i�
�'Ϩ�ҳ�O#G��� �F'	����'��2���4m�|@��W(����'#f�y�	u�2����H_�r�J�'�0LI���G��p��L[�Y�d���� 691��N$�(pj�#s��s!"O:����@;K
��R��n�F�]��E{��IP)G�P�&��JI\0�� B�<�!��[��иu�ٓUf�ș��M�!��;_s���	��=)�)�x�!�$_9@Ӹy��Ŗ-e�2h��=�!򄝊���� _&�~[�n�.&�!�Fq.�Kc螛W�>���o�!�dO�}k2����D�����ǟ�O�Op�?�Q��Z�B�ōG�&|�R��G�<���)�IAL�C���'�@�<���->j h���Z��\*���x�<1O�|͆4ʵ��>�)�ӆv�<1Ri@�G`�p�jI(���1炘z�<1��$p�l��DeC2q����7�(�� �O`gjF1V����S�6&=�Z�Y��G{�򩒜JX��Qwm����9�C͂6�!�ݖ9g�u+b���bHƅ��L$(�!���Ҩ0ҧݡx0��s���t�!��;�bq	`'�%d;���GIǵ�!��4f�h�gb�TL^�yA	0^�!�W"8� <�g�X4�e0�Ȝ5~!�U�}M�hY�L�(!ӵe�Eo!�$�]t6%�1,(u�%kڡg!�$X>f�h��D"M�ba`1�P�tL!�=uh�"�mV�?.QKk�/x;!��/���Gϯ<�� �L�r!!�7Q��7
�w���Hq�.�!��-r�ę ���` 9�锹�!�$Ӷv��9�qN�7v��\kE� ��!��J\�]�g�	��������n�!��F���E����=Ͷu�6F$�!��NP��8��+x�� @ƈ	�!��rx$	3�i\�0�1��\5j�!���>b�҉)��6%������Џ4�!�Ld$Y�˒�d�P� �o͞wq!�DR50��a��\�R,�"-�&���$��+�1(!K�:ÚAVU �y�LI���͠i�-|o�X����y"�P����%�|���S"�y����M$(2AN�$&�R�J�y2@ÔrT�M��@!
.1�ȉ��y� ߱$����-T�Lw4=�w�K�y��Y17�n	�c�VI��%)�+�y"-N0�~�*"ǟH��9�+݌�yRgD���آ'��.Dn��ɜ��yk��`��8��O)!��1d@���yҏ	�U�1���qL�kS;�y2J[]������,�Ŏ��y��Iw���vB��4�ʡ�!�y2��>�ZԠ�̫u
鋠mU��y2��^��]H"S  xP3W�G��y�a�/:o�aR ��t�@��&c��y�i�)��h�w�>io�X�րN+�yB�Xa[^D���_��q5
[��y������!0]�(�24kH��y��ú$Y܉"G@�	q��Qc���y�D�(]�y�s`׷Jx ���7�y��H0�$U�DX�B`>(
��y�� o���!��%D=�ׇB*�y��j@6�����;sgB���'���y�@ؿG�5"c�Y�t7zP����y2��Z�&�c���1o���	U�H�y2)�z3���fI+8���(TnU��y
� �5I�B��������p�B�;"OH*��7G�r0X���X树g"OθJ'��r��)p1�*
WDi
r"OС����mC�ت�'Y�&2�(�"O��YAHL.iqʀ�Qa�8E,&���"O68ڵL��u6�cB^!8�5��"Oj���54�Ġ�d�@$#$@YE"O�@��bĿo�&h��o��L�� "Oȩ��d�1����J��2"O�аl�!�`9�AFzv�H�"O����&P�:��(�&%c��m{�"O�@`��
)F#
�B�� qƨթ"O��X@���B���i�����, �"O�8�"���/��Q�K�b��,8�"Oڔ�a^�}�t��`�M�DEs�"O ��2J��&+|8Z�oB�y	��H�"O@@S��yO��Sn�U]	q"O MX�B��N��T_hb���w"O��� B�t���#B�H�1�"O��0e1P{ 9����x�"O����f1H�Z�S��B]��`��"O���OB�'	8�S�nŠM�Q��"O����
]:gmV�/���"O�1qD*��5`}���]�c�P�*D"O�����b��8�Sa��#�����"O�D1���;��r"#�
w��h��"O�u�%�1br��Aߩk���s�"O�h�tm۵e�n����H�6߆QB�"O�=�t&� I��$�DΌ�N�t�� "O���o��uJ]JdMJ���6"O��ZcN\��wm��Xb�"OA��IЖf.D5Kլ
tl�3�"O��6�2sɼ�J K��0Ya�0"O���Ǉ,[Z�p�<g �L�q"O�a@��0e�X��t˽6�B�@C"O@u��NI��j�/�z	���"O �K�*X0ݘX�H^"��
�'c��%� &����dN�D�	�'bb��Q�U�^�$��`�^*N����`U�Ě�cʚ�K뜧.�l�ȓ1bf3C$HXtܠ��${r�8�ȓ��h7�_(fz9��?[���ȓ|��(q� �/0�7D���)��?�­3�,܇U�<�rʘZ���ȓR��a#`��(J�(�c�(�� "��k��Eа[�z��L�7JU��g� (��-���E衪��BOm�ȓp�u��.Ӵp�(x��@T�yઈ��u�4�)�5��i�KK
Ea�l�ȓLv��#�B�>DRU�b�ƉL6N�ȓM��S,Ϊo�v ���B>|�4�ȓ!�!�����X�-T�Z4�ȓ_� ��� �8I�PI�� �A�ȓp.����� X�]2!Y����ȓs��]��`˙ %���=k���!�bP�I־t�V���ĝ�pTPA��8��8��c�ɂ4�C*+	�"O�9ف��s����U?YVQ#�"O�yڂ)ƲZ������+: ���"O���P�^)��X�W˛'u��i "ON�!w��;6�8\�c@YJ��"OzL;Qg�Z��8sd��y����"OΩ�4��bYv��\�9g����"O���AE�5zfau�AG\�z"O� ��#�(�x@qt�F	=Tc0"O�LXR1m�X0�X96�.Uæ"O
�2�ŠiֲRp�8����R"O�i�#�$�F4�v�,�4�(�"Ob�Y�d֮QY��+��&n�>�"O
ؘ1jN�LM�uC��@�/b�Yq�"O�LyAES�8-�����M�ڐpB"OfE��Bc��]��7�8�"OBȱ�kۚc���f�5�Dd��"O��C�6f�(�����2�9z@"Oʡ��ؠ\F�aG��2`��Pk"O2}�'�	*+F�X��Ǚ�t"��� "O(}
���>��lq!�c(I�"O��x�-�`ې��F"wg��"O�T;a�	5xY�P R	5���q�"OD<{�@5\bl�'!��p���"ON�1��H0J3�ƅ�;(���	�'� X8�*ڽ�z���m�_o����'��8y�ˠ!=na���Beݦ`q	�'�P=��#49����V�P WU��2	�']��07KN��A��Ɛ1xA��'ܪ��3ǌn)�)	Z����
�'��e��v7�]�AO�$�n4�
�'{h$�Իdq�5��Y$1_�[�'W4�"Ӂ7 �@u�ɟ*�8X��'8⨸X%D\1:q���.��s�9D�`�VA�"Z.�1Q��10<��K=D�j3'ϕ%���T�K�|�36�>D����q���V��+�>Pх@<D��@E�ߡ~Gp�{bM�@㇃5D��0`�y�h�!��J����(Rj/D���U�ת'M2A�f��T��}�I.D�����ƛ�8m��+�'#�hPh+D������0��sO��^%��".D�(��HF�q�@i��@J��Wo+D����*;̴��A�L�HaH =D����%V5L�L�Q
sҁ6D�L���&m,�x��${�4˔�?D���6�:I��u��*	�<�S�9D��3b/��]b�e͉�t�P0�j7D�@p�BU4*��dI �<6 ���"D�tw�("v��Ѫȑ_3p� ?D��0�Lo�Sg��(fg�9)dK)D�X(&�U�l�z�т��.5��݁4�(D�D*r���/�H�YtC�W�b� W�4D�ȑ��S�.�\�ْ���P��ئ�.D��!�D<���BR���L�-0D�ԑd��1b���aN���8���,D��X�G� � ͊�+˩1�`���>D�,apO[?��E����-fxz�'J?D����H'p:	H1��r�Xq��)D�D�Ō�;f�>��,A5���V�)D�L����<H���
^ ň�R��(D���6OL%c���@��m}��A��&D��If+�&�6��u(Y�C2���U2D�Ty!������6��x�z`o=D�D�8b�Z�F�0eBr�C� CRlK0 �`��Az ,�9
��C�	30���0.#z��A4��C�I�j}~�v٩*nd�ˑ(�RC�ɂĦ�8U�>K��}��+�{u�B�	��� �� �"��5��
v��B�ɛl���s"O-8���#�ز#>�C�	4+���3G��<:C�����֥'6�B�)� �q�W�
$��1������l�E"O��)�_/~ʂ`�dc� �8a!�"OJ���A��`"LB�11f ��"O�L�E���\�lS�@�*��Q��"O: TmR�7?|r�q�h}[ "O(��3J
#�"u�4��(�P�+�"O�c�A<!2̙R!�]�5�Mp�"O�С�ˆ�'�Ε;g�B�%��"OJ02�J]����!�ؤ>��m�q"O��Ȁ%�<4}��@�dʚ���Y"O�ͱ0-�$k�eS���J8�R"Obxi��L�|1`�@���}(��h�"O���F@�TtD̰3,S�&��"OJA�F��`ۧ*8<pcT"O~�Q$�ԕ*b���#�>0AP�"O:]�6�D�VB��U�-.��p"O:�&H� t�[�kX�J�Cu"O�H�`9PG���� ))��|�A"O`�*Pl�>s�8��ʁPA��q"OX0 s���	u�T�f��!�v�P�"O�i&��h�NL�SM��c9���"Op�O8�\�Ȇ�9{4�&"OjEkd��,Z^z�׈.]��8P"O*�j�� �,\��
�yz�u	��|2�)�SzX@���΍	D�Ո��MH�B��S��A��V8������E%�JB��6h~����(������G�B�I�P��jp��ԚFf�tE�B�I�B��䒝NYh`��Z?L�B�	6Gnҭd�	h� ����7d�lC�I�oc�(���L�ֲ�@f�o�:C�	=/��CtKI�Y�0��C��6���$8�D��V����6n�@Q�A��}!�Pc��2�� dw��3J˱q!�dD�	{g+�uf0!�G��1n!��c�0XaW�+X��c�͉ O!!�d�B=4�b�U�M�)��m�/N!�D�k) �:D�B*9���QL9L1Od�ID8��at��4|��$�"! � ��	��<D���cǎ&OY�0m�-����l�B�	%$���2�ܮ/���!`��{\B�I5]����F��"�+pOړXB�ɚ<�8�ҩ�"HC���"ꋖQ��O���dݙ/��y���cǂD2�(b
a{��x±i&:�#`�\
��Ӷ�ɚ`����g��p�O�ҧ�gy2��^�$�*�(T�j;�Db�!���<���DA�T�t�:5	ʾ�#K"=ډ'W�|�BW'Zj�xp�b�2U�B �?�'����ɋ(08P�T��BM�a��'Ȓ=cTI�,&T=84`�gq�a��b�`���>�O���K*
3��Y��'x�P		�'R��{�k� �ԍT�y�(�"�'>�H�Z�~��a�aL\o�e��'�Ђ �H�"ș�F�J0[$К�'KH�p0��p=�PKs�3VЄ��'zt}0����-��T������^�<��O�7����k)q�z�"J]���u��7P�p�K/Ct�[�	M�i��B� d#}��ְY!:�i�.�!f���/��?�q+=k�� ӥ�(f���VKLd�'�1O"U'>�� �H�V�U-�N���S�,D�fG��oi*lY��ݵ^�2�)�hO��6�XM��vJ��2�D�/1NC�	�-�N1X��۫2�иd��-k�bQ ����O� �m��]�J��|Q���#���"O,�r�Ƃ����+�B�Jj��`�"O�F�"f���GY�P�����'	��٫�Y�n��4���U!q�C�ɺ֦�*�&O��Ф�.�E��B��?B�� C��
t�TЦ �se�B䉥Mf�jsʎv�|��Ϛ3�B�	��n�#�)�<���H�=0�B�	#bJ^�iS�P4?����c�M�=ݪB䉵>��t�N<�]{$�m�@B�I+�9	B�m�H�{�ˑ�mZ&B�MQp܈!�,H,}�c�E����d����ț$�8@I]pܩa!D��@�+�+���Eg�+IY*����>���8ړP���7��B�?9�NɒTf�/�y�&�0����2�(.�i��	[��y"�i>���.��S�]Xx� D�(b�V-�3��()��#=ً�T?���댐:3��k�Ӿb)�L�E6��d������^:+ﺙ��"̡O���kx��=�|I�(�����"��?ʦL�4D��Ӥ�%B����FZ�*��Ǡ0D��Z��S����$,�..{���/4D��Q�- �d�|�@�%=N�*�c3��<A(��Io>� J�%l�Tɱ/�G�<����6��=�ύ�����MRF�<�AI��!/��3��$v
���%�z�<9���j2��$�̨>~�
K�<rB�E���Gm�.<:��~y��)�'#L�ĉ$��.b-Tĳ�E[i�4�ȓLp�	��֨:��E�$Lؘ&�T��	��.%I�g�t��qx���D�C�IG���C�'C����d
�im�B�	�&�0�Af�Ce^���	�	�B�I��sC�ںjzX���gU*?>XC�I-��Ԛ��ئY��e��M�R�ILy��'���Ӥ=0��h�el� @ ��?tr�0<O��O<��H9z�غ���<J%C��I\��Hv��j��2�3^V���0D���2Cԏd�>���l�|h��fg�OF7�4?�*O�#~┊UU8�P��L�~�д�e���hO?牅񤙑��1lM%S`��Ag8Ez�'�B|�`D�M�E�RIFN��Ax�'~Y�vF<h�ؐ��j��J�����'�j�R�J�3d��ܘ���ݚ|�'�Ĝ�eϗ0��;񨟕H�P��'X����L�)s�4x�!F'�M�
�'���A��n(*��FC�1A�|)
�'E�XvGç6;t2uR@l��+�'��3am�*
���:��>�݈�'J� ���)���sS��:�.\I�'�$����,K�(�;TC�,H 1�'���6�3��h�J�,:�	��'�8Z� �WR`�����0q�����DD��Ƙ���"l}�m{�f@�>PجZ�"O����nZ=J B��"��h�"O M�s�K�I�2,� AS
&HiCe�	E�Or(���� F�CQ�W�}�j��'���֫9�q)��ͱ���ɋ �y��)�o8HD��
����	};L%��fIP�gb��E.lՀ��r!�O���DNq��W>3,��OK�~��'�ў�|��C� $���bΙ\��+§�S쓅p=�F�I�`�!!EM�..�-b�#�W�<YC"s��<a�.�L�vx����{X�̦O� h��$��"j��]+�O/f'�}�"O���g�@'o<z@X��ЮU!6�za��U�����<0�i3B�C1�M`A�U�@S!�$[ ,7����ʇ? �e��	(f!��JK��ֆ����=	�/��kS���ēB��µ�5$xT���h��]W�Q%��Fyb�$R�8@��S�&�@��w)��bN�B3O$�I���uR��P��^n��R"O� ���u)�W@Z�+SL���O΢��XHt�|��	&*4����E�<��
�%&�4�~�mY��\�'�?�)``�)?|�XrhV���y��,D��"#H�;NF��@ $��P�(T�|�叝�.~�r�@P�D��P��"O�%Q ��T�
�b�(���"O�R�FZ�ڀ�Q�$ݡi޲@�b"O:�9�犱"�P0˕.CA�j��"O�`e�T*�BH�l1<dAq�"Odl�P������,�,hm��'�8���W$+� �1em�� ���'�����L?@���/ӛ%}��;�'�*5���vY�� H�9��'
R�btΈ�E��I��eyH���'- �!t$�@ͬX3g�;	NL�'fv��A��98p�eo�Sr(��'2<ag@
�ZJ\��cX�JE<���'g��a�c�:W{�>:yrY�'��A g�&2�1qO���T��'4��0�/�?�.��P U|J��s�'�`�����`�ޙ����{��'�A�JԪL�h�+ŋ�-v�I(�'��@��K�1u�W"n���'S\��Ю�)P��D쒝^8j���'��eR��h��sQ�Ѹ���s�2D���Bo��U����ƍWv���j0D����RP�Z��H��>�7i1D�䨰��>/L<볎LH��0A�.D�؛*J"H�vT��cY�c}���!D���eG�*7�p�p�:�T���)D�ؘS���>Irʖ:UN�{.(D�L?��L3hr�ł��[ ꌄ�[�$"� 	y��a"ìˌ�H��ȓrXh̢�G/��� fC�^_Θ���>�k�M�j�<��BѬX�F�ȓy3��h�nڧׅɘ����E~�<q셎p�����X<�l�
�Kw�<��o:�ڵ3%Y4Y�f��"As�<���^���dΰy�Y���Xr�<���Y��������"%���0�Eh�<y�hc���a`�)R�y䂙c�<Qk�o��pVm�'+�8�{���e�<�uA�4^��r%��.���W�^�<�) "]$P �a��PmV��`M�Q�<Y���.p�pX�B�(��]xG�P�<af$(v�@LA �-Y��c��N�<s/K{�����1�A����a�<`ܓ1i8	A��W�bqS&EH�<1B���l	V$�k��Z�p���<��);�\a�?8@jhpG�{�<�1
�3t���f�$Q�R܀�%~�<WGU:�lB`�69LX���=D���!�&#"��A��0� lऎ9D��j@+��:ކ��'�V�N|Y��5�I�Q�P@! 	T)�|D����x=c�LlRi>`	��Z�\��s�5D�� ���T �4���řH%��"O�<N�2K��I�	�{Fh2"OʴЧ�T�o!��� hۄ�ހ D"O���A)v�*X;�Ұ8��A�"O�� G����j� P��9�����"O��V��5�~�s�f\�.H7"Or���ͤo_��YV�Z�2� �"OPȪVg]+�`�1G�c�:��"O�c��#
J�Ћ"�S�-�\�i%"O��Y�'VV Y�agF��&�Hf"O2d�Q.�%��q	�핢��m�"O�@kq�]�m���k����;L\��"OxU
�eٔ԰Ԃ'`?c.�B�"O��8􂟕( ��� �8y�u��"OJ�s��8|�^�+�oL�Eo"q��"O%ۇ��	9҄i�%�G88J�"Op�V�Q�./B���i�B��A"OP�Sȑ�Sp	� ̝^]��5"O��qW �.x���(&�ȦU�X���"Ot$��a�'(j�H�$�N��:p��"Ob�2!�޹w�{2�w��z@"O�i�3 � �AYC��r0���"O����G܄�$F�{���*�"OP)2MO�u�~�z�d�� �%�y�/�M���C�isd��"K���y��W��P�����x��I�D�J;�y"�ݲ�<��(�x�&�de�y�kU�QШ�
h�ɨ�eG�y`4`��}�1��\������y�gݹ"i����M0H��L�e���y2�[_���镄K~LP�/ %�yrK�sNd9����p��#�0�y\�;��(Ʃ̹8�H�GP��y2ʒ�s����e��t` �z E�y�F�!�V�C&'B�b��K��yҀ�3e�����C�=[�H�[�H��y�_�(�ȋ��ݼV��!��ظ�ye]+V��(�@�p��m�f�ɚ�yB۷w��D�!�8z~�6�I�y≁��T5�!�I){58���ߘ�yr��+P���CK�#�v1+�K$�y�@�K�*�z�E������C��yr�` f�PG�J�QqÀ��y2�փ`�)9	�d���E%�4�y��Z�o1R��Qo���}�����y�)�20�x��C��G�"��׉3�y�O���``�18� ��,]�y�iıb#.��4�f��M��B䉗o�L�q�d� %��8[ሐ��B�ɽE�a�('��\��eJ;/��B�	�z��	�iJ%}t$���&4 (B�	�#V<CB�4zh|�������"��(Hq,��FE�c-ϊG4�	�����ē#s�)��cː>��@(����l�F|b$N�guvx1�WVܧ'j���b�,0��Yh��Y�{���5��}S��V%j# ���톽w�T��7t�dI�F *�jܗ������&d�6_*l�&�V-�0`)sI<D��"r&O�I�`EW�> Z �Q��<�U�\Q�@р���0<!�d�0;���ӿ�t�+�+D��}��]*A�Py�L�d�YG4��4�ӊZ�`-c�O�\�#� �	�U#�#8��ac�	0��8��h�o�x��|�E���i�.���Ez��`��	P�<�4�X7j���
�ʟ�22������|��
گF���xSCQ~y���۪s��� aC&0�C#:;B�)� H�pШҀL����:�QP��;4$�U>4����@��� ,�(�R�é�x���:,OhU��DI�M�O��i��4𨘪hEJd��Нx��5@�g�����'�vA�T��+���hCW,Kot��OZ�c�NF.Y��4�dET.j��Ի ����O��={�n9�I�F'WO3�P"
�'��D0��ރ0&:c��6BM*{#�Ȅs�5Cb(2f�a�$B���'Qf�t'�@H��3[��t;��
K[2����$�O��)1�Q��,��D���\.	�Cm�GK�$�h�L!�us��=ք�����Sx��2��*�H9���4\Q� �,`-d����ʕa~4Y��%Sx:�Z���[�@��T���P��y�^X(y�����^\�Ju��y��R�i�FU�E�̣P`rt)r�[�]^"q���4ޘO����R�$�8��#�(C1R���'��Y�F�\�c-(\�h��8;>5��khڽhv"b���F�c�Ӌ�H1"�OLy�oN#7��x6
ݕҹ�%�B��>����"s�M@�l�8DꞳg�Xٵ�\�J~ȸQD�G@��	���Ԃ,�4H|�"?i��%��	�
��Ds:\�`�f�'�9R	ƃotڔ�m��
�:hYB�P�3�J1�3��3Q`��r2��F�@Y	��:��4��I%c���M�W9deq£�O["����J�)%� 1�ͩ�C&e�����Q3jqaJ?q�`)[�%��s���q�&x��(�H�<����	4���#Ƃm������i�(�IQ@�	��J7AW���D�|R�̄,�u�g�>����->QJ�(ٓ�0�sVLOx��k�Ў_���
��;P8=����I-�#�Tci��������$Бw0�|c���YÎ�që�6T�X�!�n�H�=)U喱`k��rg��&^x���$QRj-k��9�(�k�?K�� �&V%J�Z�㰇 �O��2�K�W�Z]a�˃7E�0B&�'¾P�O՗� �	 b���2b��T�TA)1΋C�i� E��adFbP��2G�i 
C�	S���P�@� �I��$�>�0a�-̳q
ٴh�����FY�t�o�:�q[� ���5A�b��cT�j�X�r��*�OH��$���{tTS!�E�6<"}���'
d�y���F6�P�S��8�8u�`��LOaxb��3G~��kue�b ����%ˊ��O\1S�G߸S]��f`�.\����F^��R���i�����P��=��p)�AZ"�]Y��x�H;B.����q���J�A�RŅ8�ȟP)Ad��bP��Q
��HQ"Ob�8$O�m=�p�&��!��x2UMF�B��	�	nN	ud����g�"�`�[���Zg��[n����"� 8���:`����ݒ7���`�.%b+z!�#�!�Op� IM����dd��A�'�����Jl�I�cK��
��	�j4�!�A�Q��C�	sa�r��ֿ9�lĈ���F�B�	�&H&@Ɗ*�P2�L�-xB��S�\�8a�W�3�Ĺ��m�"a�C�I(>�y� /��]�
ɉŁٺa��C�I=E�"�jL
�D°j�'ow�C䉐45��Ӓi��S��v��A��B�ɿ]�^В ���lH^�EY2w���ɞ�F])��R.Q�D�K#%�G`!��0�n(A�F�#g ͈���RP!�$���~�;�ꏈzC��"v"W!<�{"�]/c%v��3Oؙ"3�AR�،0���#o0^Hr3"Od`�N�|!�P�?�;%�DA�E�D]�U� %�h��Hb։�T���}�|��W"O<Ua`�em�=�Y�+��,�A����a�f�Sy��FP����0���l �ց��)T4|!!�Ii,Hqm !q� ڰ� 30����Ã�Qr�`؞p��!��
|r�i��]�����l+\O|���֭57��-nӴ�
�H�?k��m`�.��ii�Iy�"O�=� A*�.	��S1
6�C�_���6M�N4�P�ԼrC>Tx���rd=��I��H�T�iT���C�	*0H�p�b��U�F�.^�@�����UQ#(�JE-�?2����+.��Dy��؃c��5δLP�N��7P�~��MFw���g̩|���qO��:��Q�ǄB
|΄
`ʋ��Q��'��[��W"��M�Aa�"vT�=���ϼl�AH��5Z7%]���]���2���wan��(V�B�(P��e��g�#PNaW�6�<�I�<�����
������T)Kհ�}� �d��B;Rm0y��'��s�8�4"O"p�S��2uj0�r7�B�ZH;a`��;g%C��ud��X��D5�g�� >�1"G�;��d��i �K��4��I�;
���cF	w<@H�� F2���04���X�Op�AQ��(����m�x���ca�I�ZqѲ�3�1����X�l4hPbLQ�\�� "�"O&���jߪj��5�˖(�*db�OT]��O�[�HL��}�tl�2q��8"+�x��JXf�<A��=S�~��W��
 군���~�I=J�C!EYO8����):����/�s|`!�n.�O����ٲ�Fu���1(,ڝr�Х[�$s	�'Ղ8qc%��Q�431��I��A�
�'3�qB�,5�܉%�N<F]���	�'ےՊ�N�� ����w��d�rB�+Eq��f)��Q7�$+R��C�Ɏ`���'�
9Zհ��Q��4B�ɒ
@���C�	:�r"aDQ(xB�	�Ӷ��e�R�+.|�@j�TUDB�ɛ�tP���Hz%R���`B�	\�1 ��\,�t�Q�M�7��C�I���X��C�#a�
0��旒<6vC�	�7���b�+Q@��3ON(VI�C�:a��m!a'��ҹ��A�4C��i��ZU��)
h��q���B��2�Z@�PE��F�\=P'�N�B�ɭO$H��-S+$8�0K��+��B�	6!���`�2��(�G u)�C�I"4a�� _�)A�����X�BC��<�T�d޵sʦp;��\-3��B䉛|R�:5U�HL����ڗDL
B��{.����n1�D�g���^�B�	�C�`��K��'���S�C� �x b@��'g�|�tN��n��B�g�1I��C����l�׉&D�PW��+M�D���-٤�j����#D�t��&��d��-rw� �txxV�=D�TW(�� UK�,Ҽk6�XS�/D�Q��6��{pmg\ĺ!L'D�`��C͊E߸Qb��:88�g"D�t���,�rP��z���S�'D��Y�����m�*��\��	��"D�����^YH-��5\|,%��&*D�س�یj�E8ǦS0��J�J?D���,8��ݙ��y��:D���e�(+�x 7`��7�px��	$D��I2oԒj7�,��J�7Ƅ�0�O%D�h��	�L����(��_��Q�<D��@�-�;[:��ص�^�&jN�&D�����ί x8��E�S�SC+D��2��"(~�����.D�l1`/3D��s/PG^t� we�(�����C$D��h7c a4V]�g+R+����g�$D��;N�3��5�Ĥ��lUؽ�" D����^�Z
���B+0�k4�?D��Q"���AzUa^�dҬ�sb�#D�p�vdWz��n@l���Uc D��r��#y�D����R,��9��!D���E��[x��p�DsRJ�.>D�3�IT�V���PG�y�d�U�<D� Ѧ�Y�� ��Ű2P̐�1A$D�艆�Ż�Ρ���'}3�X�5o%D�@q���wo��8� P�Y�*�Y�m$D�0�2ǜ8z��l���Éh>�5�"D�|��ǌL�Z�̌
�y��(>D�� ����;���X�L�2��"C"O4|`t���h��_�,�Tp��"O6�:�c�"j��(���νC����c"O.���hU�J%27�K��I*V"O�XQp�5-�X�ہ�$˪	h�"O�֬P�k��↥ʠn�$$ӓ"OԁptD�>�^����εBMB��"OX�A6.L�u=��%ؽ4=~ux1"O���GdǪ��'%A�DT{�"O����ǻ-�aK7lI�5��"O����(���'b�"8����"O�U������xTk�4��""O�db�펎ayR}�cJ��B��"O��s�Ĵ,��uJ���|��"OHl�[��0�W�Je���"ORI�F��^� �rFЇz
R�)C"O����%�� �$L넨���X�a"O ՛�YkؠĈ��єH�Q�"O:s�.V<Js��Q��0@:���"O�l��7{��Ag�UN�  �"O��Bd�ȧA{n*���%uB���"O�0 )��ZN՘Q&&He���"O �i���z?�h���VS:�+a"OQZ����`IN����;Cbh�"O���VL�oJ.iQG�	a����"O�<�f��Ws�\0òQҪݙ}!��Y>4��u��!�[��	3(�!�$��Y&�����Yu����ё	y!��'D��xAɻBX��۰��d!�J�Xzu �K�"��pgeI��'$�܂U��N&R�Ak�x�l|+
�'L�A�A�D&��/��
�'c(a�ۏ!�蜳ck��'B�4��'<��Wǃc#�(�C��o%
�'�nU+ȓ@ռ�"��/ư���'����&oP�@e�\{R��Q�� �'�"��D��{/Z��N�0Vz"d#�'����W��<rk��HRn�7E��tP�'g��@P�0w����GR:�Ƭ��'lD�bb��o1�%��J�D�
�'�.���̖g�PI�."&�X��
�'�@����چ|!a�����s�'VjLke
˕s�tx�aO@�2�R�	�':T�5NJ.	��`*^ 6Έ �'��Ke�"U��-�(̉(���Y�'��0�E�s ~IQe�N
 ����'^�!�娉�G��铧Ǉ�T��'�:(�s/̬H�Y{֨�>V��3
�' ���C�R���E��QN��'�̈� %��I<�(�Ţ��{6@z�'e�)c�d�j�"0��������'|���&�^ %jKC�ź�'����J؛R?�m��k�-"�AY�'*���e�S�By(�ض�t�H�Z�'T|9��(D�)�V�@&J�b�t�y�'����G�h5��r�LRP����!+�X2��L���UĆ=��)g��H��'��;��Q�WN8��_F���r���_�p�6)�!bJ���O3p�{dM&qܐ6/Q:t�r
�'˾|��j�.n=,�u��;h�h��x���ڦ#� Xa���+O?œ`��g��Dـ�Ir �9r�Z`�<�!�P.v2�C"��6�<9 ��Xy�	�B�P,�R��Iaax"�P�nP�}�G��.X�(��Cͦ��>	��M�d�5��]&|^u�P� X>��Pa�[;h��q���� b,XJ��)3qM+{f!����2����� }�FT�|RaV9p�0|�2]���pI�m�<yu��
&��{�j@*z �\�4.럸��Q���w�OEy���ED��!��?z֘q3!!��p$,C��YT��fү0�q!V.���ʓH��t�f�ٻ�l�Ó3�bx��	
u��g'	�q� ��I�p���F7�\��ψ1G�I�$���@ŚU<y�ٳOs�<��Ϗ����ΛS�����L�&;D�X����XBQsOO�b+�HC��+!�!��������&�����H��D@��2��#f<��ӡ��	5��[ϸ\��&":TpB�	��h�Q�[03$��y�D�-_V�n�Șw�!lO�0yEg@2�.����A$Z�Q�1�'��A�Ô'���'ӱO�4@C��$L�]���5D�蘲��:m*��d.~J� H'h0�t���j�8o.��D!��"%��<
�)��00��$H�_��B�	�t�xڶFC�W�R	Q�ĶdYG��ha JU�a�E�)��<I��@�@�f��-PC��q�R�<�Th��,᢯O3'u���r,�N$�m���+��#"G_�*��e�3�]7dC3��c`���P�M Ԅ�67栐I�`<��c�/r�H�1'ޣ�(�Rc�/6��w�4�OPq6m��z �ԋ��D�M�z'�>�7݉5#��!T�)H̾�􏅓|�ځXK|:Ĉ�Nᒘ���a&x݈6E B�<I��ζs������y��
�mJ���\C'MM3D8��	��pخL�|�GI\ r���0q�����ޞw4D4�b�κ ,h���V�w�,���- �8;�&"��2T Us}�ȸ�@��b,�Rj�*E\1!��d��"�xi8���4(Z��F�'I�џ�����<sذl8�nV �4I�E��?���"�7OAxu@��׶�@0N/�arF�u�9!3��"7�� �����Č�A�츗cD=A,N����sH�P��A�ħRP���D��}�����ެC��3�Dr���/UT2��L)eJDp���&s���Ze��8Ь���E�=ؤ�(O�l��;G��)���*~�~����')�p��bU:]&l�؁T/aVPd���L&S�N����L�v
��l"��'�����gW<b,������d �����^�l���.O��t�П&db��<[��Ac��.:,�8��"O��;r/_�K�d�߁3���G[����| �4h⧟�"�?y��(q[�����N.�T�*D�����,�\ف��#�-��!~�"�9��a"�3�	� TE���@*T�e�6@[	=VB�� �c��q�܄��.�??��ق�OR:W�!�$O�l����7GH�*IY�*�H!�D,"^�(C��Э%&)��(I.�!�T�^\h��LN�@7�#�@�!�$F�E4~5�%�S.P���#��9�!��I/�t9�dG)y@M9&b]o!�M5i��8AW�a�}3P�8&B!�$�iӲ����_�](�G@�B!!�ϭ{L�3cB�-'
�2Z�TY&"O�dB7�S4�(oE�L]D�XG"O콩�AC�(]Cp.C�,D�M��"O⼘r��&E>�U���W�OP-� "O�PU�β_��ʴ�гX�h��s�'�
5���>���J�p,}V�L*���c�[�!򤂹�V��"� 4����NX;R�O��3�.�b�S��)�Ssj$y& ��=�,�#��J�!�$��Vy�S���?8�y�� 2Q��4R�g�9V�jU�'�@�F�,O������@2�OY��� r�"O�H���8=�	!��վ=lN��5oЋ<`��sF�R��ɧM�^��#�H�'���uꏅq� �����a�p����ݠC�27-��^d�I!d�_?T������;�!��7	xl��'�a���䀆Ac剟]�-�bhߑ�9$C��>5!�M��x:�tّIN�UǞh2ы.D��% ��%
�v���|�`��rm�=^�h.+��Q3s��P5�u�Ɩ��}B�ҝn�\t������� F��p?��Ip�� ���"��M�`���5�|�g�ѻ)�Q�Q&	�����	�I��̙$ W5CH���t��%\���>�T.̞Lfu�Ĝ<N@2@����?�u�iF�l���҆*��E[Ȁ����y�bǶ,�����I ��aTD���~�lU@Y�(�� ��H����h�E�r�;5P"�Ѵ�L�|(��a"O
�C4�!n�� x4�KiV�i2���?E���&� Ed���%[�~�g��re�(�|��Jf���X�T����%R,\�U	B�,��9IЏ ��,	�L֒X{4��RO�a����2R�T��`������Q���	Y8 ��E�4;1�0���K('�m8�`��i	�A�d"O��j�M�rE�d�J��W�O�`r�ˊ�@)��pH��}��E RS]��D�BL<�3t�d�<qT-�.�j9���A�d�f��a�	� �2P�6��m8�`a�ш^��@���%���ҧM"�O&hq�MѲ6�%D*=�,�!HC�L�&$c�'Ѫ���K�7hj�� G���R`�	�'x����fC�J2�d�&�^�r4�ā�'�VłP�ǽ{�V�"�	u����'(B��C�Z�<�,�S�ΩG����'2�XS��Ԍ%��Y��.tM��:Ru�P(Xc	QBbI�@���U���t'M?8�4�8c�Xh~%��&���ǖ0����Q�ަ%���ȓ=�>T�J�4��-K0�=Wd��ȓd\��S�;!�0͚��˛w�`�ȓ(B"ICUi%�  ��ŕ�g�Pi�ȓ*n�"2I
-?��C�V;R���K[��&�C�4�Z���֎C���ȓT�S��2K����lӎ	:�l��@ɪ���)ٰ�c�#�'tN�t��
��!@��)��ɝklt�ȓJ�L�����L��c�aX@����02�k�)�:X`�#�kw:���C7���悝(�<u8A�Hd��I��7��U��[=���Aϔ�yN ��n�ީh�BX�%پy&Φ0z���Zd�a%PZ\���� o-<���o�`�g�o�Bts���#X��Ć�33:���̂[�l�k���_��}��J�	��Ch���"��{܅�F��h�)݊Q��H���&[�!��&��X��^(�U���!<�h��"Oܬ��+ɞ>^<���֍f%N�"O�
���#q\^#u�@�.����"O��!��C \)�0-Ix�B"O�Y�e	I��؋!+]4{�x�"O6T��Mܳz�h��1
RBhb��p"O��dۊ�2d�gj�K�v�W"O.�"�!t��=ٴ`� �����"OZ�qҌƼQ��}S����L�z�*�"O>P��L�]z��� [>R��$qf"O�=`mX�m��Jp�]��,���"O|xCsL�,r�~@ @�G�� �B"OlȲ�	U� 
B%"n����q"O*90r��,.��՚�憸Dۘ�"O|=+!	��]��eɮ5�{�"O��q��1<�R�{�jEl�]5"O.��Ə�)Z{���JE�v�DC0"O�A2 �r��A(�"_��B"O]��KD�h�d(Y�>\ �pp"O���ǆ�u9�DZ����r7�s"O|��7$�u���4���!"O�4˃&�/ P�tĎM$�|"OP��e�
���#�\�d�0��"O� :T���ս^"��Ġ[9$�$1H"O��g���d�i 7-P�|�"O��Rd�Jb��-�S�>$�w"O<�kԤR!<SB��ժ���@�6"O��r��\�]ԲpxbI	,hnn@�"O>�ɤ��w5H����F�i�B��"O~Y��](Lu p��)��o=J��v��Bh2T�ӆ	V��������$=�1O�`��c�Iy�'X
{�|��"O��҇��V�({���%�,t�d"O�!�C��
���Jf��n��"O��"£Z�8�Ę��RHJ4xp"OtM�F��`<�b��I'ڠb3"OX0����6�=��I�8-��:�"O.�.un��RD��5mV(X'@�yB��/=��p��$-aTI�����hO(㞬�t]�p��ul�	A�R��7dkj�+F����8�'��ЀG�\�gɧ�O�"e��ƛ(�\m؇
���(!��o����}�Bҧ��<��B��Lߜl���X�Q�P:�ӈ/!Ƭ�����򟛎�dڟ����ěg����ɂ!���I�>OL�q�4�"9Q �_TyJ|&��PP�	� �`���N�H=�s�ۋě$P,Pb��蟘l�`�	�i6�5SҢ�"v7t�Qj�
g�ԓN<�d��L>Qb6��mJ\��!Mɢ(�6�H%I�f��EPi`�j^�?�ȏ�I4qF�U�%4�
��I�\Jj�S\�=�S�OSpXq&eP�z&69Kadq>��'SQ�wB�3�Iǳ>�~b�MJ�+��fDY1M6���a\�\QQP\)hG�[�DS:z��ɵ�U��a��2W��XC�ϋ���qA�� ^]�%{
�<���E��y��i_�K�,@��M֝b��L�g����'�4]P�'� ���i��ɀx�ҍ���-J�Hd�`c׸N/C�ɀl�H9)f�� ��,��d �C�I,�Q*v E0e���d]�YL"<!���?�8秝<Rh�20J�"�zQ��"D�d��_�-�@H�I�,a͐H���>D�\h�$��A9���*
+TZ �w�:D��j�NY"g��]rS�*�jh� �>D���
	S*س�*R�8Y��6D��r'o^0g�D��
DX4��9D���G�2.sF��H� )��&'6D�| &ɜ{N��S�ڡ� ip�4D�TpB��A����4�&;����3D��c��Sa�D)�!��R�x�q��#D�@��-!G"f`��	
~_<8���"D�h`¥�%����E��8' D��҆�B�V�:�q�k%&���
��?D��#MK�s�r���M<���	>D���q��,x�	����j4�
;D��Y����ܼ#�!��8��#�F-D���OC(7���BB�\-"9D�D�v�����$�2N��l �*9D�lC �S;i����I@�p�!��:D��W��K��a�Kd1|���F6D�x�`�^�^���js�nv��(D�h��S�]Vh1c�G�{�TD��%D�T d�'����Avf�i��$D�˵�	t��I�#�����3�0D�@�3?ߐͺ3�\0��2`N.D���D���i�$`5��'Ϟ�o,D���
�+1$��%H%mkzE ��/D��#R$�T�j�C�%ʒQ������ D��`���^@S&�\�n6�i� ?D�l�)�6�jA�nM�R�XQIv�>D���W/
8P��X��J��,YJ�J;D��3p�ښA�TTDG��Mx��9D�P1c�h(��/D5:����h$D���指�s_��y�iD��c$$6D�� 攘vH��7a<���e�i��\D"O�Y��]��ݒ���W�z�"O��1�M�~�ع�d�1>�T�c"O��p��]�A`U�ڟ�X��"O�ՙgZ1$|I c�M�"O��׵;�$Y8$;td��"O�y�E
��Yd�p�a_�,�, �"O|1�cϡL�� P�V+��"OT}B�������Vʤ�"%"O�Q��
�?L&nx��͙/<�xl�"O�Y�5Չ�J)x��E�g�L��V"O(�bj�;^P�*Y�Fi`�"Ox\��K>>�jmy��� �*�2 "O��*v@B.g�t�8�e�;'|� "O�!Ӱ�O><6�4�S�Z����V"O���iNr��t�X�"�R���"O��O��Jz��]�
̾�8�"O�8��%�y���#�`p��"O�}�u@�K�N�ₓI��=`�"ON�KG
KH���jٮN����"O���F�F�@|��z�;x ��	�"OzUS���9|z!�6&U/�!�`"O<!�@�b��pk � �s�]B�"OjQ��j��,L���Q��u�R"O�`@R� �,Ղ���F��L�$"O<�S�'��+龄�$a�L>��Ba"O��K�F]�t��1B���-y~ЕW"O�A$ǽT��t�O7wMs�"Od�Z�hӈv�䓰� Ymȭ�C"O$�83Mۧ%�0m��R�D� "O,����@�B)�A��x �"OH�!LR|X���/ҵ|[f�z�"O�Xpb�)������0>T�ҷ"Oh�q�r_�,��ş
��e"O��X���b���C��R#U�b�+B"O���B��dh���ǟ�5�U�""ODXa���4JWr�v��0�dI�"O�`��
A�:�(�K���8z��"O��K�ν8'tU�4���qV]a1"OHM��D�$J���O�5�^��s"O�Y��Y�HaR�I0�C�U�"�I�"O`)Ӂ�"K��z���2`d0D�"O�!G�drB8����SA�5��"O�E�%�\9*6�)t]�"O��!g��b�T�0���~tXRe"O�����X .����p��#� �{�*O�@�6oݥ_��	� �M�o X%�
�'1Nl����.^�U�"��:*^��
�'�Ԙ)@bܽ5���hR�D4&��	�'4u@��Y�~%�$0�,�&"圴��'0<I��j�3!`����,N��y�'[hu�2�F!CH8���H%H8 �k�'�̩Ӧ�<��:a���@��\��'[��Fc�Ö�R%-[�=�\��'<�X6/�:X�x���5	���'~j,``�2f� $9cn@,/�Z�b�'�n�IE(��"���")X�(�z@r	�'Ϭљ5$ÍT��m�r�X I�OK�<i3I�;�J�B���$_��x�]G�<�"b��B�r�������JX�<��F�p��1���<�>�'ÞS�<1!Ŕ�/c�����N�p��GZx�<�'T�Hx�����60����K�<�!-γA�`}��
�q��!��J�<� 2�K�Ɗ-�E36�ѱq�,��"O������$�D�f���Gk�ə7"Ov���%��%0G���L`���0"O����j�)x8�U�MRJ��U"O��(B`Չq�+Կb$N-X�D���y�j�	���M��^��8��AG��y��#p=��*CE�W�Q!����y҅׬B�x�J�	!I�`������ybF�:��آ#-O���b�݊�y��O��f����;b�@,�%:�y2���օ��<n�l�HQ�W=�y!ȅ&Vу�$F*l�^�bPi[��y�k/`<r�`��i�vl�GŒ(�yhJ+,��Æ^�OyqЃ���y���"�(�0M�L�çS��yb�E� ��v�ZC(�(9��π�y˶;�J�#Y@���C+��yb4E_����&MWऺ&��y�nH-��T(��U F�T�(� ���yC���Ez$�+N�rMRE��>�y��ri�����,6�D�6ɀ��y2oA6Z`�e���3cm��&��y����-{�Q��f�]0J@�5-
��yr��:_�v�;�.N�N�3�K�y�${��hYpb��2jRУDFħ�y�F9U� ��C$1B��@C"�y2"�'p�%Q��֮6:�;�@��yb�S�x��
GϏ'��%[�� �y�O�4<�J�F@�̠�D����y���  ��e*��׃ �4���Ç��yBҐ0��cP�H�����yń$[t����WO�<a`���y�:`>�c���Sm�YR��y2�\�iT ES'���L���Q&ݔ�y��A4Z��!��ϲb�aA��^��y�l�
nDT��v����͈�y2n΢�re�&K�;|�R)�1�y��N�A
H�	3�D�nE`T�W�F��y�Ʉ�rR")J�V�b*�v��yB���:$��X:^?�E�N��y.Tf"x #"Α+4�Y�����y�#�[��0t�X<uY�q����y���3���8ő�q6�A��y"C3^��k󀁘]\,��쎱�ygC�G��d۴��X�Pa�����y� ;q���w`��Jd�
�A��yr��2-y�!'�K��AQ�l��y��#�δӁ ?VȄ��N�yr�Fs8�q��)L�v|#�-U�y2�S�_����VᒢF���ѥ��"�yrM�A$�T�J�<s���`e( ��y2���b���a� ��5���y�+�	R@x��4n���D���K��yB��@�B,�K�Uj��"
�y�d��L�z!mWl�X�w����y�&h"�)�f��>Ԁ��X5�y2K�0/| t��W�ڜ�����y�BB�S����e!פOsHMa"���y�G��I]rPAH@|�
����y�.�+P���X7��=?�!3U��!�y��źW�����k���y����yr��o�`A�q
Йq���@�$�y��U��>A�6Iݘc������%�yr��(�Y�ǃ5aN��`��y
� ��Y���c����U�Ξ1̬4��"Ota�J���9���W����e"O��@�	]�Ab��堛�Z��m�"O��2��.6e�,�D�B$����"Oh�xf_�5q$􁴡_!U됵&"O��� `II�$HB!珁��7"ORh��c�'9����'����""O��a�Dg��=�vN���#�"O��z�
Q�>�(a��Z�Ru2"O�I�g`k�>�Js&�;`�$)�"O&�0f��I�����3���"O`�bb-����%c�$S.=�M��"O��C�$:����4��OЌ��"O4%��1]��]�CP�4-��!E"Oĭ�1��	I���1Q�͹&���"O���BX�0�t��h"�0W"OJ�P�ʯ
��a��\��T�`""O0��@����e"t�tS"O8�#�J�<�	�Ӂ�4��"O.
è�5Xұ(g@^+b�B	�S"OUȶkD"d�!�S*-;l❊�"O@�����F��2g�*`�q"G"O"<�3�WF��Yr��R�٪"Ǫ�#
'7
P胆�אE��"O��t�		3Z~)K�ㄬ]��%�"O�d��.�8R0(Ɓ��-��I��"O�tQ�%��yZ�iB%*��S�V��"O0`Bc�ӵvTTC��]�$�R4cp"O�E��пri����;���"O��*E�!6���2"�rtr( �"O�iq"�>\�G!�Ob��"O�ٛ$
N�F�t�ԏ�&j󒕫�"O������>���M^�<����"O�)&Q�M^t�Z0LJV5���W"O<9�J;d�|���Ŝ>��{`"O�غs�����h$%ǰv�I�"O9�5   ��   �  ;  �  �  *  �5  LA  �L  X  �c  �n   z  ˁ  ��  �  Q�  ��  �  -�  o�  ȷ  E�  ��  /�  ��  G�  ��  ��   �  d�  ��  J�   { _ � A$ �, 5 m; nB �H �N �P  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�OT�y�G��l���"�R
0��7�OVh<Iq�\��`q0Rn�
��Ku.�X�<�g�D�t�����K"5fX�8�Cp�<�!����uM�J!J]���l~=ODc�"|�NV0z�1� ���vOC`�<ic��?n�봠]�Qݸ�
�A\���=�BפD52�[�O�9xeR�J�e�T�<9���%��u�E-]�T��4��bIN�<AKCu��i3��	w�ʽ��d^K�<�f@��dl��ց	�q�s�l�<1ҍہL�u2S��<��\�C��v�'<ax�-��XK�m�E�9O�n�8C���yҎ!Q�~��2��H�H8e)�*�?	3�IK8�Ȱ�U���a�6���� D�d"���=L<�GE����q4D�$�MteE�PƋ1�M��5��0<�׭�1�|ɚ�aG�q1 ���O_�<9UI�?@>`KT*ɓ]���ܟ���]&�!���H��ዒ<|J݆��}��v��@ �+����6O��D��Y��4���_*w�i��)вA�q��G�'����dZ����Ae��uג�'S$�����I�Ɛ��+<�����'�n�������C��Z�2��Y �'^�sPbF)��
��Ղ�B�'���c�#޺[�<���֨*"���'��@@�F#n2��᜕%Β��
�'zn-���~>qy&��8K�
U�
�'+���g��*�`q�O(Dߚ`k�'z�!)!�'mCB�dJ�8�� �'	0�@���Y�z����	pY�'��XE� �H:�ܓhAVX(�':~q�����X`��ǚ(%P�z
�'����M��i
U�u	A�,�$\�	�'�8�f��36]���K�5B<C�'��PMLN����U�R`��'i�tBDo��_iZ��	T=O)����'�T��F\<f)$��w�Ѽ��T��'���K�+�f�ᡧ	�~]v�h�'��<�P��Fܞ�c��D z��Q�'���L� m">0�*Ҹt�Pc�'�2X��E,�>����n��}�
�'�8���_n�Tx���Ba��)S
�'���r�ζ~�
��IC.�yb�^(\�4��(\,{0MFI�y�KH�|�be��n��~#���y�`�8_���p��w��}��
�8�y��T�S:����ўoߐ �`o^��y���2�n������x���B����y2�/]����%Z��L�q��5�y�P
�4u2(�?TĪ��R���y����L��Y'C�Fp�0r+M��y��
����7���)�X�Y!���y"瓠[���(���W���IO0�y�J55�bvC�"���
�(ɛ�y�
�XFF�jr���.B0ؐƈ<�y
� �}K �G>$%y7��"zF�ʖ"O����H5~�TJ���J��B"OX��3f˸Bt$�h�K/J�@+�"O��Pe�
}�����$TI�P"OZ�Z�mϜ{`E�#+K-m�h*q�'���'���'�B�'v2�'��'����4���4�3MӜ1NQ*�'���'�B�'���'�R�';�'�8��Lj���H`�X�&���Q��'�2�'�2�'��'��'#r�'� y7f�8.���0��>10�Ļ��'|r�'�R�']��'���':�'r���$�=3j���� U��t ��'tR�'�B�'�'���'��'z���U��2B[3q&Eٟ��	ڟ���⟌��ϟ�������۟�����:T\S���1.T�2T�Vџ$�	��	�t�I����I����	ԟht�R�I"J�VFD�&	������՟�I����I�@���|�I쟤�	��<+C#h�"b!K���J�ߟd���h�I䟰�����������	��0��}7��"�㋻r���i��\������ϟP��ԟ��	����I�d�0`�)o�⽹��|��) �[�d��ԟ4��ß��	�d�	�� ���\
5뇮j�vu@�F�%�NmR�C쟔�	��������	�,�IʟD�����4z���U��o����M�̟��	ԟ �	ߟ����L�	��M����?ic*�8K=�FHȫB���������I�����������yo�F��iR#C0�p��)���?��f�4����O�`�G��,�QŇ4`��҈�O�ج*986�'?9�O�|�i%��"�e n�@���&�"զ�7��'�V��D���A�f)b�cL#]ڎ��4�{*�6��tm1O��?������2"ϑx�`HXp����)_�0�,�$�O<�	b}��d�՝\ڛ�<Ol���o�9|�f�`�h۲E�aIW>O��Ɍ�?QDN:��|���)��F��dŴ��U/��FuD0ϓ��D6��ئ���<�IU���/��F.�����L�@�?�R������͓����4��ʅR0\Ͱ��@�ږS}�	���uA��-��b>��e�'������]�Պ��*/ lĨ_2nd��'��	�"~Γ*�l����C`8Xf�8%J֬�*�ff�?����U�?ͧ��E��ėsLj]��`6����?9��?��H��MC�O�擇�*-׉w���㝈�m�j�O�p�O��|2���?I���?���6x���x��C��S��,�*Of�o8h��	ԟ���|��ԟ�
"A7Tj��B�����0��H�'к6m��]�K<�|R&AƤX�FqB��fA�fOR�;�4=��iT)�?�1 �j�$в�Қ�uW*)}���Dy"+�*o`0A�b��P�t��2x���˟��	��STy��e�0�:��O
(Kta�CBܘ��
ϔ
���!��Oj1m�X��#_�	.�Mƿi�7�ׂbH��t�T;>����A�~��I��\��r8� �?��'�����] ��.'��D�C�U�L@&e�2�|�����X������	៸��7m09�&A�Dծ,��2��X��?���?�P�i�B��Ot�dj�6�O�D"!�ѿ�B0�j^�<�RacV��d��,�MK����$�_�^	�F��0�F�䰐r��R�8�Q��T!
����!�Oʓ@�R��	ӟ���ǟ,�g.�s<�s��h�x��!.Mݟ��ByR�o�
Y���O�D�O��'{���Y��VK�@�GŔ���Y�'^��x��fcw��'��'%��<���D��X(�f���CbI³ܲ� ݴw�剓�u��w?.O���@A�6����6-�9)_����Oh�D�O����O1���"�vG�j�ҬȲ���ds@iC"eF2cg���'��hvӶ��-O7���Z�M�R�yvゆ	���nZ��M�m���Ms�O��z�������U�Pr�k��u�`����ծ1�~!rf+��M[(Ot���OZ���O$���Oj˧ mv�iV�Ey���)��<��i�~�`�'f�'H�Oe�Nu��.]�.?.]��NI�}�T��Y�l�R�l�5�MC�x��DGыU�v=O"C��֎{��@���I5:��ʂ>Ob����4�~"Q����4��d�O^�$��f��Ya��
Q�IH�Z�-z�D�O���O��T��n�#���'��f� ��;��tͰx�-J?m�OD�'��6�Kئ=�J<yf�G-&���S�6qy�H]�Γ�?�Qb6G�l���4M��I�u'	�l?q�J�����³7�L�Y���*cu�!R��?���?����?�L	�A��yG�ҝzV�oé30��ӂB�C�R�}�@�Rd��O\��F�1�?ͻ"*tt��R�9\�)�ӟ)������M��i�6mZ�`�6�l�4�I�9��(��ܟ��bs�@�R`
�
 �U�'��D%�<	��i��	ʟ��	ϟT�IΟT�I&2qY੆1z(|r0����|��'��6�-'Ť���O���9���O�B�8_� V���dV���bdy��'&�VD$��OE��O���*��O��\3���+nb��1A����f��<!3��AV�	ayF`��^Px�`3�Q '��G�0��	;�?����?����?ͧ��ȟ�����O��s�D$_�f�c���-2D������O�nN������M���iE�7�@�̕����~��}X7�2}і�P0.y�d�.˜D��F���>��=� �3�EތD�<EH�iM7;b	�&;O��D�O����O����O�?�EЫ9�8`�:Q�<Y�(�џ��	���"ߴo����'�?Q�i��')����B��5�!�4�T�I�?�D�OR6=�N�sR{ӈ��Ź�J,�,��_Q����4��<fZ��D������4��d�O����+��D�f$JM���GT;#���D�O��p��lI�xa�ß��OsF�B�)Y��h���A����O���'�\�B7�r�)�N[�8�V�@�o�"�T�����t�''��<�������l�A�|�dAvD��3gK��AQ"��#׬wc�'���'���W�$hڴ5�$@�e��oo��@FƱ_�!����$�ݦ5�?�@V�L��4{�v$p�@/P���J�G$@l�1��if6́�T��75?���\���)%���P[��g��]��!�S�3�y�^����柠�	����	��O1X���._���`u�V�e�L|!2G}��T���<9���'�?�S��yǡ���P���M=z<��8�ƕ�6�DꦥqK<�|����.�M3�'��[f�	�(ɒq��*_�9A>A��'#���bM�柌��|]���#e��n�ƴc��Q9NͼP��F��h�	��IDy�es�8����O*�D�O�
��
�v�ȱeg%�ĕjg�(�	����æa�۴q�'}�]�3F�-h�(#�k��L���O40�B���Z�V�٥�IF�?����O�j�)ކZ����l����T��Ob���O����O2�}���9u�`�c�����d�_Q^������&̑)_��I �M���w�h}I����Iv����,E�U��'j6͞��ɫ�4p^�!R�4���^nY����*�9s��N�P��`*�-�*�p4�1��<ͧ�?y��?y���?�6dM<L�$��?Ȧ,� V'��$�ݦ�+�GQ����ܟ�'?�	#�B�(U�՟�Z�[�έ+H���O>�lZ��M�U�x���IK,#�Z�9��W�H�yЪ�6,�T-	w���U� X��b�=6�O�˓E~��qf�YH^l1�7	|�ƅ���?Q��?��|�/O �o�4G�� �� y���$��c�"����E�b	X	���M���(�>�йii�7M����Fɓ�7�$��F��S�^��q}�5l�J~b�P��M�S`�'�A��g�����eO֡�E�<Y���?���?q��?��DD�|fv�9� J�N�ؠs�)�GB�'�IeӮp��<�'�i��'H�ENۖOݤX�k��^|C�A!�DC���i��|rà���M��O* H��|���艝y�R 0w���~-����l���O���|���?��e��Ihd2��2���27�NA���?�*OX�nZ��&��I՟��IZ����'. huig�C���d�#���Y}b�'�"�|ʟ���r"م0*��ڠo�"�rĦ<'rҒ�Eeg0��|Be��O���N>I�`	�"��ѣF�\+c�҆C?�?����?����?���Q���'��
i���	x䨚7�S%�&��l���1�	�\�ڴ��'e���?����?I�d`1�E��1��S7�?��i��L��iN��z>!�����T��D��"�<y�b
�bc�X+�L{��'��'��'�"�'���i@���Μ6/Є `�!Γp�	K�4Y������?���O��7=��h1���P�*Da��@1L������O���T�)��$t��o��<�פ��U@"�hS�=�4���Z�<I�ʉ86���v�	]y��'���(h^H=r@.D':$��%צ*���'���'u��M[�	V��?���?��
D�i�x<;��T�S0�����'O�꓉?9��R�'z�1��4�
�H�H!A)&��O��"ȡ8�*6-�L�SBt�d�O�e�ª�JOVRd����Gi�Oj���O����O��}�\ ������(��)�5I�4=����V�اe�剒�M���w?(�yQ�Q� #���p�X�2Y�ț'u7m ߦ�3�4c�h}��4��$��!e��9�OE2 	'/��U�>�ÁI��&�O�����O����O�D�O*��Ym��8M�A���pw��$p��@�F�A0#2�'j���'>����O_3V
lհv�C�Yf����>QB�i�>6-Jl�i>��S�?�c��
.p�fx�`M �x-��m�7+���L!?qƃȂaU�䘂�����	��� � W�H��4C��F��6���O�$�O
�4�@˓)��Vn��OK�"B*���A�DYM[XQ���F��yr�|Ӕ�Բ�O��$�OX@lڐv*�e��jپ,�bɺ�K����$��"�ɦ���?�ӂ-�^��lyr�OF�)�kp��	�Ԡ`ڸ1���y�'���'���'"��ɗ/�J�{��Ҭo�����q�t�$�O4�D�Ȧ!��Lp>��	�MKL>	���1%T��e@�**��\�Ƅ[�1��'������E�:��&���q���*�\X���<,��M�>N�����On�O���?���?1�:�����HL��}�B�iC����?�)O l�GhH���͟$�	t��*6�4�3D�?�mpnܼ��dVV} |Әln�$��S����o,bS�Ů'�uـ�	,� ��DJ�XĲ�O��J�?�eg;��a�]��@��qN�|Z����9;����O����O��<1`�i`P��없*�|��a���Q�BQD�L<<��I��M[��>�U�i���T��m�Z̃1.�(>�T��F�~��o�`�LmZQ~2���m�X��'��� `(I@ᇀ$J�y����-w�ݻ�;Oz��?I���?����?������C">@	7���]"�Y��eWh��<oڑq�Ĝ�������D����$�����!M͒hQ��0	X�fb���u�2IЛgj�<D&�b>ݺg̜���ϓ%�&�ò&��U�H���,X�l̓.k�顕�O��|"[���ğH��OڊT�LI��Q]��,���ğ����T��sy�}�F����O���Ob�"�#�>Jab4Z��3X[����6��
���O7s�~��##_ m�0 ���N���Bڎ` P��t0��|�` �O$��p��q���:�J<���J��T�����?����?����h���Dͅ+3��S��Z
T�c�o�a������EH�iAjy��`Ӏ�杸
z��3dk�6�P�k7$I-LG`�	��M��i��7�	a�N7�~�h�I�wؒ���Op�Yy�*4��-�f�
O���Ʈ�U�Ky�O���'xR�' 򡃙	ژ����9'�̩�j�_��'�>`��fY1q���ş`��t���'�P��ˎ�x%@C��x)�`�>)&�i��6@a�i>���?I����"��-�We�6���a�X(+r�;?	7N6j�v���7����ė�\�2]�UFK�X�a��̄#a|"�{�~�A�OT)�5o��^-F�
 DT�4�#Q �O`�m�j�az��0�Msg�i�6�2��R�A>..��d	��5��nb�H�&p��kS �?�%?��ݐT&��'�]J> ���^ :z�	x���Y� nn��E�M�"�c��ޟ������4W�f�Ou�7m8��6ɆI����+x�2�ڏDc�e'�p�	̟��9:�l�D~���d���P�N��*���KT#V�a4$���N?�L>Q.O.��bq)�ow�-�c�)l	�-�!-D�F�<|k��'�2\>��&�g�l�h!(�?{r����,?��S�L�	ϦyN>�OM�%���.gЕ���0R�y���}'V��¿ih2��|ҡ���@'���Z�R��A0Eh�)&�V=
׬�؟ �I̟���b>�' 26퉆*��%h& If��уD�f�hМ� �۴��'����?QA]�{^fi�MV{�U���?���U� ��4��䟗j��A�����^/!Y�Gץ"��H�,Ȭ�y�R��������IΟT�	̟��O�:�����"#��Zl�"@nL%	�l�O��"r�'�"�'���y©v���ߺ1V@X:�dA�!�X�&��l�|��O�$�b>�dO���qΓm�FMQ�ǀ,�=��eH�얥�tz�ȲA�8%�̔'O��'Er}��͐*��1��jK1ol�P"��'��'�bT��C�4HDBa����?1��lE��������W�N)x0�̊�"`�>���?�G�x2ʅYx��णG�@\|	�����G�T��ei�l�,�'?qӂ�OD���<z� 5��D�z\F!`pʆ%���D�O �$�OX��8�缓W��.��4a�Y���1�$�?�@�iԒ�r�'2�b�<��ݽ;1��A�2z��b��X�����,����M���M��OX5as�H����Ɇ<��0���������!��'����������I��0���;��SG(B=}$E��?Ze|�'x6-�� 7����O���(���O
l1 �Օi�V�٧�C�~�=��R}��'�B�!��)�3:j}šW��Xi�v|����Ql�Jԗ'
���f�O?�M>!/O�hjS�dg�Sâ�	1 "��O��$�O��D�O��<�E�'4��:��M�,m@�eÊz�d�E�C^���J���XV}rKjӌpmڤ�M+�6?�|����F�b/
|�!�ͩoTy�ٴ�y2�'|�m;�i��?� �O������ze�(*EB��4���$U� 9O�d�O|��O���O2�?U@��؞I�4��
I�'m�P�DKZğ��	ß<K�4:΢Mϧ�?�W�i��'Fx���5���CLb���U�'�$�ئ�ܴ�2L��Mc�'�2��qH
9s��?=&N��੊W��9*��r?yK>�*O����O��D�O�i�uIjt��B Ɇ���j�Of�d�<!ѿiT�t�p�'��'g�.Bў�D��3(����k�!Sk^�t�Ɂ�M�Q�i�hO�S,$�,�qn��?��-0� ѓ<�H�B�A�|��l���4�z���'
�'��7�OW��@���V59<���'$"�'��O5�	�M��L�+��<��N)��x`m�3:
����?m�i�O*��'�v6�͛f@.�c��y�j��B�^�m��M{RS��M��O"���.����]�H9��{>v��@����`[��`�@�'���'R�'���'�哒 ��n���,}-�V�x�	�Ѧ�h�J�`yb�'@��lz�Y�Ae��u b� "*P +����r��ş(�IM�i>���ܟD����U�_�S�	�d�J���ߎw�p�̓0�,`�O�O��0M>�.ON�D�O�s�HV�2�P��"A�T�$�O�d�O8�$�<!��i�[��'��'gn����@(QƼڴi�>6�F���Dl}��'���|2���Z�(}a�)�?f2�B�����Skt%���{�6��Z-��~����̎p�PjPc�!}{t�+X}�Z�����?����?9��h����� k��}�f��8DYz���V�i}��$V�����KNy�b�x��� t@�vM �BA�U����	ԟ����x2�@�����u�����G!� 2��"ߙ<��phehN.K݈�i�:���<���?q��?	��?A����]�6����Nh�Xf������0����	�%?�	pZ^��@.�>?nى���3���O�m�%�M�@�x��tE�Y����ېF�:�E��_8�
rā���$�=�2|p�锓O>ʓ!2��ϮA�:â_3z]<�8��?)���?���|�,O6�m��9�Zh�I�0	`��4a̳S^�ib$�C��	3�M3�⣳>��i�7��ئ��l��%a�kL.S?L8p��œH�l�{~���a<0��m�'��k׫3L!���6s,}@���<����?Y��?Q���?1�����<a3n1�h���� �^� ��'��*p�aS0�b�dꦥ&�pi�E`��� �RF`�-F��<$��1�48����OWjLP��i�d�O�40&@>%bnK���t����/V�4�.�k��QH�O&��|:���?Y���pŃ�.^+�̠	Ua �L%���?!)O��mZ�v����?��'��K��&`�e��=.pL�ӡ�w~��>���?1J>ͧ�?�c�W{�����!e\�����3'f�5��m��M��O�����~��|��ܙ]���m�[�L���Ú#W��'���'���X� ݴ%|��e�Y��n��C[]뤰�,��?A�b"����FLyҼi%&�J�iT�.�>�P4l�&)>��Q"r�&�nکu'�en�Z~b)T�.�6���c�	E�-�^��J�s�|	��#�<����?���?1��?A,�����_5!e�Y��W9����Q�C����`�	؟'?e��'�Mϻ�=V�OFBtJ%�IQ�l��6�r�h%�b>]A�����)h�A��6?�hqCB�_0��͓"J�`���O�+H>9+O��O�݋��V	G�v a㎛�%_���O �$�O����<6�i�y��'���'�6 �Gd�T���`7BL��qy��Dx}B cӒYm�
�ē��I��N�\`8<{��%7#\I�'��z�*ڱD2F�Z��tK�Z��'���a�eW�k��N�\	��'/�'ir�'��>����/
 s���:�L=*���I.e�I"�M��`�)�?I����4��)���, ��U�R�o�=O<�n�M���i���f�i3���_D*�!#�O�@�P�˟�JP�R&_dRbVd��gy�OH2�'�b�'����c�"�㰊x�l�҇���J�I:�M{��Ӿ����OT����d~/�	3$�*�@E�����9��}�'V7��U#H<�|Z�oZ RT�S��E#X��=ڑŒ50Ĳ��WDp~�#Kk|�y���`��'y��H���x�c�
����N�|h�Iǟ��̟��i>-�'p�6M�?��$U~ļ�Av��-�����a�d�T�ߦ��?��V����ğ�"�4E�)�pj�h������Y]Q�Y����M��OpE�de �������w�:��gQ�x�
)�5��->Bh��'x2�'��'�Z�M3��/Fw��z�c'L�x/]����'l� �2��������%��ʤV�n�TJ�7Yzp�B�%�(��~��f)}���U�~dd6�;?!�	�܆X+����.�X��V�`���[��0%���'M��'���'�Kτ>Nla�N�/h��c��'�"P���ݴP�����?����R��~ ���B���y��a�&[��	9��d�Oj��Gr�)R7g�}Ĝ���.nv����5ts^)@�J��MDY��Ӈ;Q��;��:f�:�ů#wޥ�w��&�����O����O���)�<��iL�s3�Tl�B$D�,�P���Z�1���.�M��$�>	�C8��4�ʾa1T�"S�ԏp�P!1���?Q"�M3�O����k3Z��Տ��ɵX��X�.J�+��L�t��)��<Y���?)���?���?�)������g��I��e�{�(���P���᥊�uy��'���enz�	��NO?5��ej�����J��0�M�3�izfO1���'ky�\�I�i%.�Ł�j���)�ר*F��ɠ[����OԓO
˓�?��B�L臠<G�V���H͈�?����?���ӦUR���ay��'D�	sfI�>~�T\@�A_}�����D�x}bo{��lZ���o^Α�Y�$A4]�AC�$BXTq�'L� �¢�s��V�2���~��'(�-�X8[j&B�T ;�y�c�'�B�'�r�';�>��	�1V�6HT#-�hPh���	��$�I��M���[��DǦ�?�;eF����bA=Nj��( �&i'��.-��cm��lZ'E�np~2`�M�L4��Z��a@wbO�x)���s�X"!�~ �O>�+O���O��$�O����O-`�j֖"����,�
}j���f�<y��iM����'���'H�O��ώ3Fp6��\E�x�c�Q 1�꓁?)���Ş!z��ViUg9�JT3	�s�ȖX�B11,O�$ U,��?Y��9�D�<Ab�Л~Hu(0艿:!؅C��E��?���?����?�'��D�٦�᷆ӟ����z����I�W_ƬkF&�ܟ:�4��'u�듵?Y���?�r��_�ƥ���5�F�"�d܎[����4���H�\;�����t)������2<N 8jv*�(@��|�
Бw#�$�O��D�OZ�$�Ox��?��������0.$f9�V!Ҭx�:���ʟ4�I��M� �|J�O�Ɯ|2�^i�ܥ�vcL]���0Dg)4a�'�B�����L�����^H� ��Ǆ�2�����σ%N �i�D^ �?q�h0�$�<��?9���?9p��ݪɢ'ӹSh�8��S5�?�����ڦA2�!E͟�������O�BH�S�.%���'�Ⱦ ���O���'���'�ɧ���'À�w.�f��ˆ"
A�ht0�p�qqF��;p`��?5���'����<�k�14�JBl�p؜jr�ן��I��D�	�b>ٔ'O�6-�:T��Fȉa�D�·�U.2b�qQ��O���{)Y���Em}�s�j(c���������W@}@ǥ�U�ڴ�6��4��Z\����������`Wz�q�X>GK��p��[�V���[y2�'9b�'?��'s�T>E�(�:>�a ���M/�	��o��M��h�'�?A��?�J~J�c��w�b�5�/�ph�%��\x��`f�Ɖm�=��Şn*�d�ش�y�,�U+] '
�Z�� �E�]2�y�B�8 i���	5]%�'k�i>y��"�0I�E}�<�3�o2�}�Iǟ�	�h�'_^6-�w�^���O&��F�I�G˝5�NU j 1_���OAn�#�M{u�xro��"aٵ��G��l� H���GE��,蓉M�8�1��<���2���D�>p��v!ϹsZѧܥ_�@�d�OV�d�On��:�'�?�P�-��-�0�� ~��Ъǜ�?��iN`���'��l�0��]�P�(y8��V
~���ȇ�
.J&�牟�MK�i1�7-V�H6�5?���ɕP�X�I%=l�P�`gW�_�n)��$H��f$�K>�/O���O��$�O���O�=�HƼ�,�1�"$R-�"�*:��!݄�"�'>���4�'��������z�L5�0m�B��<A��M+��|J~�%�E���g�!W��Zq��, -z� m~��̐YZR���;~��'Y�	e�d {%̎�1Fl���"��q�*5�I�(�Iǟ��i>ї'_�7MƄf�x���=(��h������k2���D�,�$P�A�?��]���	��P��_�De��I �h=<�4�?!��fM����'��x9&���?E���T�w|�!GgY,��9�7)�Vk�q�'u�'���'[�'��Ɖ�L�2|D*��_�{�F$����O ��Ovoڸ|U���'�.6M7���{�Ś�F��D��h��ЈnP��O����O�i�&Wv6�1?��V�`*l[8lHJD赊��d�n-	��&�?���-�Ģ<i��?i��?����>n�2��T�Y��9��+��?a����$����P�Bҟ����ĕOJ��m�p3���/�?���S�O���'�6MM�q�H<�O������;�zȂ� . �sτn���pӱi)n��|��'���%��JGlۙ:.�IЇH�;��`hf�����ܟ0�	��b>E�'�^7m_���A `�F,<"}�c��$F����3��Ol�Dæ�?��Q�<�۴IPP@ �A�A�@��k��O����i&7��dؤ7m,?q0�[$M�H��UyL<\��$S�XTlz�B����y�X����ٟ��	��	ȟ<�O%:< DIJR�*��^��(=Swfk����P*�O���O@��������]�B7�U�%�����˦〥X}���I՟�%�b>����I��!�
�`���,��̄�[eÌ(QМ�KɖP��O�8�H>y(O0�d�O<u�g�U�x�$�A����\�M�O����O���<A��i�|L(d�'@b�'_|��I,E��0`��԰u�5ɇ��_{}�'L��4��r��"�I��� �QG˄]<�	q�!¡$�˦�J~��㩟t�I!Q�0ᦈ�ATj��6��6��	��͟D���t��m�O���F� 9S�M$\Xt ֌��wf��z�j\C��<�T�i��O�6u8�B"�:vg�yu�=k0��O"�$�ЦEA"Ҧ1�'[��;���t���->�zܡ&�J�]�P�b�������Ot���O����O\�H���:�T�=�Ԁ�6�RG{�ʓsۛ&#�=��'��Ok�O��}z��H �}��R�N'���5�>���?)q�x�O���O���G���(��$S���#�ՆNw�6�<�H_�<��k��ny"#&2ۊ�)�l�)�J�jS�'��'�r�'�O��I��M�Sn�
�?�I�"��q(�L�UI��@���?�V�i�O@��'j��'#47M�:4�J�XS�݌v���i��d�2��Nz�8�H��Z���?�&?��]�@0��*�F�����M�����������|��Ɵ$�	Y�'g�`]PU��V�Ȥɇ*�H�ĭ͓�?!�^�V�.���k��f7�dX\O�q��L�NN�Ę�OA%;V��O~�D�O�	ϲy�6�.?V�ۓ<M�����Y����DV�r�������&�h�����'���'{�t�N)V���S/zW����'p�\�Tx�4yK
̓�?�����ɟm�P#1�T2jaa	C�]�+��	����O��d$��?�ᧈ�=E��L�C�Op�R� �~�(� �σ����d��~?�H>y�%ϩc1��E��x���m�?����?���?�|R+OZdlZ<asb�w�%+������&Gy^E���ڟT�	��M��b��>���%?r��'^#N�X��̿oV��Z�!{�ֈݲj�f�� �S�Q�P���<�G�+n��j�/�z���F���<�.O����O����O���O�˧?��!5"�#k�pKe�_�Bn.e��iA2�#�'���'x�O�r�o�����YR�ēN�@$3G��?@����ON8%�b>%�)�˦��S�? H��Ĕ�Gr�p��Q�JD$�!<OH�Z&�҈�~��|BY���	П�BC��67 �Lr�#�B���D�V�@������Ay"e���s'�O���O��@� ߲�D�C H|�(��j.�I���$S�U�ܴ$C�',�<8�d�lMҤ�g��F��O���`���⌊��镟�?)Ī�O`Y!������D���4�S��OZ�d�OT���O�}�� �P}�s��7�P�#co�P!~�a��a�fJ��qg剼�M���w�F�@f,Ί!�Q2�Bڕa/��'r��|��@o�8��nZ�<��������@ ��S<D�|F!1aݞ$·�Q�����4�J��O���O��d�X�lZ7f�8�3(L l5J�5:�C�	Ab2�'i2���'�r����:EC�`C�oY:��8	�F�<��MC&�|J~"��f��sG�F��m�f�јR��;��D@~���1����Ɍ y�'��I�8<j H��;;�����Nl�d��؟����x�i>��'�����Y�R�]�w&r�c�����T�C~��Me�x㟨ȩO<8l�M���i��Ax�˖ :s��Q�*�<丸��H�� Ǜ֔���m޵~�d����J�1�jE?CE���W�Xo\|X�=OT���O��d�Oz�$�O��?��W*2W`���K�y���$��ޟ��	��h{�4 Ύ��'�?�`�i��'�����!�k�:�V��t�X�*>�ۦ�ش��T��)�M۟'Fr
��~-�C�c�Α��c��\��(;`�Pz?YO>�)O����OX�d�OB�Ё��(2��1���ʩ���?������򦉐�&�ly��'��7>w� xw#Q�`�KX�0ƺZ��L��O�n�MОxʟ��[ЩEA��T0W�
#I�pdd[�_���9n_y��i>ms��'�Q%��:��2q�9�ǪM�!��H�h��D������	ʟb>��'�6MھFIR�y��R:�Ҝh$�J%wD4 نD�<�D�iR�Oʜ�'z�6m� J�nyz��c��Qt�6n�/�Mc����M��Otq�����L?	zw����pS�@�;rr��Ĩk�(�'���'���'K�'(�Ӵ48&��� �l�dpVK��y�Dzٴ)�� ����?Y����<�&��y�#�;
(��B��]�P�Թ�##֏%�p7U��qO<�|�BMB�M��' 
q�ҙ>ل廄A�j\}��'�(��lX?�J>.O����O|<JN/M��Q)[�[�FI��/�O��$�O���<!��i��t���'��'#���
R\Nj� u��� ����d�x}� r���n���c�q��bJ)7)��`k�(�h��'kR�����v�1��R"�~r�'rZi�0�M�p��B�Ā\p\u[��'���'���'j�>��	Q	�+ƈ�b���"�G�6k����Ms�S����_즥�?�;:V���K�7X&�'"M�=��@͓/`��.k���lZ)%��\oZ_~RnĮ`b�'�0���eZ��'�-f�]�J>�/O���Ox��O����OF�B�	g�x�1���kNv�;Ti�<y��iݞ<z�O��� �Ӗ.��J��H�/cHp �G()�r�O:���O��O1�ltS���@e�D�(AWB�+y�6�??���Q�j���Ih�Ity�μ-ne����2���AéD�+���'8b�'��OD�	)�M�¡��<Q��Oa �B&*1��*�N��<)#�i��O.��'R�'ar�S5\Rd�1Zmf>TiV$P�3���;r+Y����'B�@#F��t�O6�%U���� �:[��9�+�y"�'N��'���'���I��f�^��F�r��)���@����?)żi^�(�̟�lk��X!8�L��9	�>�d��H<9g�i��6=�����`�d�D�"f�X-=�t����(pC㦒�l���	�Iwy��'��'���F�e��!�Xp�����B�R�'4��(�M�� �<����?A/�v){�I-%>��c4��.BXd���Tr�O��d�O��O����!`��z�v-J �Ÿ{V(|���8%Wfeo�`~�OĖD���>n��K���93z!IJ����{��?����?��S�'���ʦ���n��$@�P��.��c�=$���ON�v��MW}B�'� �{mTp��ͮo����'*�cO26ěf�����Ǟ��q�챉�l:c����/@���b�2O���?!���?���?�����)�$b�uX�D� "��l�?VQo�S����Ix�s�dh����#��"�)��P�>Y�Hh`�S��?a����Ş��|1�4�yB���.צ����1D����B�.�yBm
�;�,������4������O<�0�ăڠCvmR�Ƭ'��$�O����OXʓ	J�v"F4
��⟠,�|*/�@�Xs���n"~��?I�\���ɦycO<1��Q-J-ȴc�l�*'�`!_`~��ٳ//��"B;ܘO4���I>\���D�4W �!U �t��h��?��'c��'�����L`���5��՛�&#/\~؁
�ǟPk��S?@<�'�~7�:�iޅ��En�dRCT�"�:���c��@ܴ\H���hӰ	pՃ}��\G�t�e�������J�gX��?hR�C�·�䓍�4��D�O�$�O>�$ƣ4,f�CƊҥ1�$q������kћ�
ײD�2�'>R���'�:)*uiS�z��H	%X��Q��ı>���?AL>�|Zm�r�? �a!�U�%F�[���0w��)bwc���'�h�*�h�OHbM>9/O�e镬W��x��Ў.�v�I��O>�d�O��D�O�	�<�Էi2�}���'c���"+`�U��H'���'�t6m-�	����O�6m��]b�.	?�6���:YF�\6C҉ .�m�h~"�!I�P���~ܧʿ�D���;�"���P+$�H����Z�<����?����?I��?)����1j��mЂ�٠>ȺX�����2�'��hc�Й���?)��4��~T�Æa�kuDE�l̫~;��g�xRGxӺ�lz>�����Ѧ��'�������*~B��#O7T|<s.#wPB���o>�'R�i>�����ɅgY:�ѥ㒴$�� *�Hy�����ȟ��'3h7��@��O�D�|�e�ÿ`8�,R�퓋z�Ȑ1-Q~���>��i9�7-�N�)���
 ���醟��\���	�"���
c�F��4����8|�b�N$�q�	6q����G�F#��'ER�'��tY��iߴd� �W!��zr�"胞@�
u�oE����!�?yX��o�\;j�³���:*E��GL/���4Xz�V�l��������� =�D�~:GNn�h�J��$�v�P�<�)Ot���O(�d�O����O�˧"����o�=�H񫥉F�7��X9P�i`�����'�2�'G�O��iw��֢EA��æ�t��󆈟�ZQ��D�O~4%�b>E!�ۦ�͓���K�a
ow0	R��W����̓�F���P%��'Ur�'���� U�C�z����.9����#�'T��'�Y�Xp�45�U���?q�K��[F�S2{3F�S�.�=�
lь�h�>Y��?A�x�CM�rP *G����u��`8��d�<;H�h#�s���%?�z��Oz�đCf��~ɂ����۳5�t��OH�D�O���2ڧ�?�c��!�����iN�v|�3$a��?�i=�Y`2�'��b����=D^T)d)Ol-� �f#p��I%�M��iK�7MĂ}�6�"?q��\�"�����{k��ڢ爇& }��T/z��&�x�'�џdZ�S�L��K�L�D�Ќ�T�&?��i5�}Ks�'���'��4q"���?��D"�eA+��1���c}b
r��!m���S�'Cu��ҌԶ@hy����⭃Ť��M�U��`4b�&��"�$�<yld4�8QdJ�~�L�h�hG��?)��?I��?ͧ��d�����X�6(D&-����IH�.�0K~��Iڴ��'����?شjۛ�@���Ii���f̴�'fʺm��E�¹i��ə)9�]ءџb�����7���@��xI>,�v��(x��d1�O�l��	�0*��a�M�:S��ɴI�O$���ON�n�(�4�'F`���|���Z�����Ҷ]3��Q*��@�r�O��d`��I�6Z�7M0?��O-n�DH�rK�/��b��7��!VΤ��%��'x�OH���x��o��p@�� �)ћv�P�!��'�Q>u���6?��B�>bTL�e�0?�5T�̳ݴ>����/�?�@$l�{��H!���N�n`���MDֹ�1���U"+O��Vm`y)�n˺]C� P�ዹW���b�,]i�r��g��H}h�*�C�#���0��1mڰ�!�E�|!�h"0.VE���r�j�f!���U��"�,��P�<�োY�J����E�Ф��O��/e6:���JV"E��z�D�)\4�(e�=@�n�I �֏H5{�U�e�icUk���V�(@�S�=t���`�+l��(��ە8 �պ���6���{�A|��k�a�.o��Sph\�]/\�&j�,�ր�<�����[S�.�z��7\v=��D�#V@��g
1� GZ� �0�i�>I(Ob��7�$�O`��B�LT@=�gM&ڮ��à.C��0�4���O���O����Mz�O����q�F�x+ܕ��0ZX��4���OƓO`���O�s6��s�ȝ�*�t��Y=n�>��H�>��?�����D�Ж��?y��Z�w	й0)�;s��ݣ���*'h���'%�'O��'3��W���d�8	P$���i�j,jw�ʔ(Q���'�"���{U/p�d�'��O�=�"-
�5�E GfS�� X`�:��O�D@�n���;���?A� �ߞʄ�������;�c���<��ڴ�?���?q�']]�i�!z���L��<��lN�v.D�I��aӒ���O���Q�%��sܧDQ��*�C�.!��)@��iD�-�I�/>��n͟��I�4�����<aV�Ƶe����#�U]�DYD�::+��U��O|�?�	�29 ��p�Ҿ.r$��3���W�Z���4�?���?�w�S���~y��'��D	c&VQ���H�)�&�I�A'~K�O�����?�d�O*�$�O��0UL$	�H��%��hfTQ"`cJͦ��	�#�FA�O�ʓ�?!K>��)��p�JCD1\�b@��5�PI�'� �|��'D��'��� s`�	�+�2z}�I"�H-��1�&�Z}�_����F��Ɵ������A)6�2`�f�L�
2 9œ�"��OR���O��#?�	����DeɉH<ȄHv	޽.���b1���M)O���<��?���SK��O8~��&��e��e&���1�O���OJ��,?#�Ф��I�OTy*@�������(v�����ɦ�I}����ɨS=��=ibD1͐�"�ό(4P�d��Φ���ԟ��'�nѲQ?W�����$aزl��Ydz�9R�� Z�, G�NK�I�\���=�H��?��π �pKfJ~.��`�e
7� mq�iH���ݖ�o��0�I����� ����VeR�!� Z���wE��7�n�p�i+r�'i�̨b�'��'�q�-�ׅ�^5A����X�i�X駇bӼ���O����$]$��S�.ئ�z7@%;"v��!�lBش�?����?�J>��y��'����b�S��\����X�X��G}�����O��dL&���'���ȟ|��@�Ĕu �I7���EIo�ɟ�&�������O����O@ᵪN% ����j��m��PDF�٦���*""Z�L<�'�?H>�;��#��35jY�E�L�N��֟Ė'���'|[�h Aص2j� � n~P�@��Y�^J��0K<���?�I>	)O�omd�I�k@R*`�k!�Y�"O�6�'b��˟P�I����'�.Uъi>���B\``"�����G[�����>���?�J>+O���O ��!��n:�˕���^M3'^T�	��'�ҧ9l��������j���u.ѰV���#�<�M�2�'��	)yO*%����2ML��;3��XF8l��ia�Z���	5i�@�O}r�'t�\c�������J��)Zp���M1�JK<Y������:0��ݓsG0 P1-;*h�U�Q+;���?ٖ�-�?9���?���Z,O뮈(C5�Y��� \`��t��:��v�'2�	D�#<%>�c��4So���$j�
?y�XQ��ӼQ{t
�O$�d�OD���B�S��A%\�(�є��4��}�����]�6�{)Z�Gx������i��\@E۳H�Aihln��I���MMyʟf�'ힹcA	V�R�'Xf�>�#&�����������Iq@���A�+O^b)�&�nӐ�o�<�w�Sh�(O�<G�M�$佪�9k���#`�x������O���O����h
d`��)�d �aťT��|���Ħ4�'�r�'j�'��ɾ9,�"$\(�p� ��GE� ���@�'�"�'�U�@��aJ���$b#%k�)����4�_)���O`��'�$�<��Ŝ��?	��@�$�m�֥R�B�PK��]I�	��,���L�'6H=#�f�~��$���I6��,FF-:t��p]�ǰi�Q��������	�]��	~���5�`R�eߒL��܃�&MX����'�Y����6��	�Ob�$��@T����S�֔:�.K�@�]I�`Vd}��'X��'C #�'m�s�����,���X-���ˀǋ�:[�n�eyRhٝ<��6m�O>���O*�)�Y}Zw�d=;�Sr�۵dU<�p&��ڦ�	��s�dg�X%�t�}r��N��{P��;+ľI�F��J1�	7�M����?���"�_�|�'Mx	�+S�1J�U��]�z���Q�x�i�4O~�Oz�?����L����@��!�*���YO[�xI�4�?����?�t&�S���EyB�'��H*�~q9r�L��ȤX�S�aɛP�,�	�3���)R��?����r�PC�%x�"��
ۚ @L�!E�iFҿ~�^���$�O�˓�?�1v�Z%�i	S�Q 6JL�Cs�����.{���O~�D�O�D�O|�p~|�h7�!F�~$XAHȨ'pT�d��
��	HyR�'�Iȟ8�	����C��2T�5a�,*f!��xE�T�X���	џ���ߟl�	���'�):Nv>eSu*
X�����F\aE:�A�(r�^˓�?�*O\���O�DR�9��T(+���d�4��5��b�L�`n�՟�����4��@y/��u��'�?�1�x�4��6G��:d��h��Qn؟Е'���'aB���y>���c�rD{T�I20tJ	@�g�ᦅ�	ß0�'N�ۇi�~"��?Q�'0H���1o��@cr��K<� �b`X� �	̟��	- �	a��'���o��(u�Fo�,-��O�"���]�\�O� �M��?!�����_��c�fIr��E)x�(mQ�_�7�(6-�O���+a�?��8�:���+rD��~��С��-"�6�J�GD��nZ���I�����į<!,M�fkJ(���BM�`����p�i�����'3"\�8��Ck�rvO|�=
Ҡ��L�I��i�b�'@�J2�R���D�O�ɐ39d�h��:R�שN�9�f7m�O��L0@Y�S���'�"�'8d��D�_%�\�.1RB��/b�
��կ&�"(�'��	��'�Zc�,|;T΅�NN�	�V�t���O�X�r9O��D�O���O ���<ya��f��tI��X^t���ٹe��(��Z���'�rR���	ܟ��	�}uB���DRd	ځ�[�0ƪqX�m3?��?���?Y(O AE��|BFA��'��9bj�'ml@������'�RR��������	{���I7����D��<�V��=&��îOj���O@�ľ<�Ǣ�'d���������j҈���C=V�
x������M�������Ov���OBLB�>O���!"�-ѱ��L�5��{� �lw���d�O�˓����X?���ޟL�S�D�>��BIG�,�����8,u��B�O ��O��$0I��`y�۟p�hC,ϲ_��akÄ
:SN��a�il�	�6:��iڴ�?!��?���BN�iݍhp�*��x� È�HԎx�i~Ӭ���Oz�zT>O&�Ob�>:���}mr3�%,_� h;�.~�uФ�Φ%�	������?!ɩO�˓9<�T�&$ڍh��,�2d�4{R�౷i�23�'W�'��r�$�P�? ����A3G��Y "=`2��i�r�'
b�^�L��b����k?�iN�m\0I[Ï�?bM,iBW�Ҧ�%��g�ħ�?1������O(��U/�A��J��M[��� U����?!����#�I� 2�J�+���	h���d}��I�yB^�4����T�Iyy������-�8 �*,��JýohB�X�>�I�$���	K�� K�e�7YP�z�p�jԖO8��wy��'b�'��I�D��O=�Z��\-S�-j�n�7ZJ�I�L<Q����?Y�J �ΓVK�i�K\�X�8D�TD[=<~Bm��W���	�����_y�	�Hu���c��g��5(�
HA�q`�"�}�	}�	ȟx������w��H�"^�9S9y7&��q�]5Ny���'P2_�Ċ$Ŷ�ħ�?���"����;eN*cbP�!��xB�'�b�y2�|R؟P$�h�$�s�ҫXH�X�i��ɭ?�\M��4ZN�ʟ\����N�d�*��s��a��I�d���'��I[�j7��|r��H���3�K�X�>��
�<X��&��/ ��6��O ���O��I�T�I�̰d�7�2@C�X-81��n�	�M���<�I>Q���'Zܬ!��^�9�d��HV�*���:WFm����O�$-b�:�%�(�	֟0��6oD5�5g±8����-�'P���nZh�I�Ko6Y�M|���?9��Q���u�	�c$��b5mŔ{z����i�r�I�[T�Or���O��OkҝW�Y[e��m��x��kW�0���[g���Ly��'��'2��8d�@�gKmh�Q�-^�#�d�r�f���'���|B�'�b�L9���GA�	y��IX�C��u(��'�ϟ<�I�X�'a� ��b>�"��B�y����"�ўS�A����>9���?J>1��?��U��~b�ѱ#ڨ ⧉�6>?^�X�/B����O����O��l��5���4숉���2_�5E�(�K'�7-�OD��?��?q��<�M�D�'EJ98߸�1d	ؖ�@% t�����O.˓C�������'w�\c��y�� �0 T�:��B=h�T<��}B_����x�Ӻ#���,j��1�#�ը>O�#F�ݕ'(��pRKxӆA�O���O]��>�6�h#�Md�@|�섡A`��'n�AIz�|��4iV"C^����'�C=&5`b�Y=�M#ձ�?1��?�������?a(���q�� z����B�V��\�T!�<	MY`���ON2��Ӻ(z0	�0`�:ii'Ҧs��'�b�'90X3��!�4���d�O�u	�Y�[�P�vN$nZ6�f%�A�h.�<����?���g-��P����A�����k(��i	b�(%b�'��맫?�I>Y�gG�q̼-	#)�&P~�9C��].ɉ'_��OF�d�O��$�<㥃)o��0;f,��n_�рg�:cf��2���Oj�O����O�IŧA�&��RA	������z���<����?��������'j|��餍��X��99NG8e^X��'���'*�'���'��:�O�1�Q��5a7t,sP!��WpNl�BY�d�	ϟܖ'5�����)�Ob �R �0(Z�	�5D�9Q���Ŧ��	J��My�؜N�P�M<Q��Oz��A!kE�Ep�H�d���E��}yr�'���b͟B��zRe�bRI��;	�衤O�;a�'�$>�H�d�=�~�T$E�B+<�rT� L4ܴ� �]D}��'����'�2�'���Oj�i�2"g��rd���ȿY���2a���w��@Z0B�j�S�3�6�aF�W�6����3�6z0n�m��t:����ٟh�	����{y�]>M곂^�
`��T����!��2��ă}"�b>����
��Ae��7����oP57Q��4�?A���?i$�[�g���w���'�R��e����dC�|:����#=iH>����?I��X���+ L��rf��د+Oz١��i�BR1��	<����OB�O��e���CA��C�^-!�0O����>�1��)��'FLx��+�:Q��`y3�ܡ`����"O2�R!�Q�T�6��a֊!~�����I�0eb%��$p�p��+2���A��i���U���=�f$I�$�ν�C�S�Y/���{Q��2�H�Z4u�M�؃hK�@���CB��7;6�r��K�h5��Ѧe_�p�����$}u���gF�U�AF˼1�	�Th�0GU:Y����;8N4�1F�?_G:���G!�=Xq#�hIȵ� �L��?����?�aQ�;]4���C��)%��T&�S^��EZ�'́t��]1ԯ�[Y��<9g�iܬ�k�%�D�
��/Ql7��ޯ���1��&�Ըc$Q�\z���O���"��o�y�-U�Z���8��]���	Q���z�G��U��1c%$��-��5�O�%'�<��"FR�<,�v�C;AR���WHf�� I�����O�ʧ)Mt���?y��9_�1����(���h�W+%C�����!����r��"A��	*��O�\�h��(�Z�㓇؄8��H�r�ʱ���qI�'.4J����E�"~�	��l�*��&o��083�T�\_A�˖埤��O~J~RH>���E�%�������b# �$��B�Ɏg.��B��}�� gE"!��#<���)� 
0�ńC/Rf�$v/̥_ڌH�s/�O��D̥x���1���O���O��d�ź;��?�U	O�fl�qJ�<S�\�'�
�i�˫,�(IK6�ŷLspD�g�'�Ɣ[���Pɨd�t�Ŗ9��}�S��O���jǍ\����լ�����,��H(҆�E���p�r�����6D��'�ў�'4��4'�(�D}�$摢� ɋ�'F��Ǯ�R*����5|>v���?�S�dP���Ti��M��%�v$�KI�cX5	�K�1�?	��?��� �����?��OH��@!�ܹ~;­pE^,@[hђ�N�L�2�R�®u0<as��'���ȡ�&BV|Ar1i�7���i�#X��t�q�ӭ%�~� `�'��t����?	��ޑW*���	[C&|���*�hO�?A���"ǨȚa��b����]d�<������>�� �ڡiEr�#Q�M�<�U�,�'Q���B*{�4���O�ʧ`B$�"���'i?>�T�ĭ^Z ȔlM)�?����?a�%H�}�
2���5]^�I�$�i��t�����1��0����W��<i�'�	m�8��B�����O|:�A�%AV�� L\�V���H�b�'��,*��?0�i�2S>�(�bS�'�(8��	�6ڭbt ̟��?E��'���2v�ƍ�Fe ET�!��m:b�)��6�M�]?1q0���L^0��%��Zi\��&��<%1;���P�C�I�� �7@�G�<yQH�9)`�Cf�IC詳U,Jh�<�k�-Y�С��,�1OL-�� �O�<)�Т����g���-W��j��N�<���!42-@��λ�����O�<���,O�ܣRf�2j����AL�<�w��gP��ƨ@��`�
�K�<q%lכx�8�[�.�%d?��(���~�<9�
�<"\0�$�ӹN��pף�w�<��@�~�ⅪG6!	��v�]�<�D�RlYF!�	�/A�YH�N��<�v�߿q�����E�uM�1�Ee|�<	�L&�i�����}��eQ��YB�<���N�r��ŭG�@�"3%J~�<�b%�?t�M�2E �4�Ҡ��U�<� "2X�P��d�80'b�J�h�<���҂-iz���	HQ:,��`�<I��Ւ�X��������#U�<Yvf!5G�0�� Ǘ23�m3��H�<	��7+� �:5JؑWb�J�TK�<�4��" {`�bbj�bEd(�wmLD�<�O�?p+�0��NObrY��Yu�<	��v`���G�mW�1�`'�Z�<9�c�� �h%[!���'��s��CV�<1sk��)�|��hK�-r|���o~�<�%�H:#�)�ŎB��Bŀ�G�R�<I�GF�"g�ԩo�E��Nv�<�fM��֑�JA�,	�	P1�_v�<a��B{�|��'5����":D���q�"==H��k�$�"�7D�X�$$��F<���< �Z��D�1D�`7��B����,�*��eo.D�0���Zc�����d��찉#$+D�`�*q&洲'f&Q������[�PP�bO)j�������9\7}!�䂯��+��y�b�@O^��4d�0[���Ճ[��~r��%���2/o���s�͹eR>��C��7j�J�y�O5�O�jU�=Q�L�chU�<�@bFK
y�b�S� \.�y������*s�	s=t��eC��(O&�3����F��G=_&ɘs��k��/���y��8Q(�Zjb���
ݖzj=P��6��e%�"~��%K6�(�a <��EH�h�!+�B䉔J�𼚠��T����ڽ|4��!�ƀ���	��p=yS��7����@���0�b5Ӆ��W8��UL�{W�t��eG1PF~��F/]� ��)�E�U�\a!��M����͑����Wş�iQ�h���I��Ȋ�� �E�s��(�=�ƈJ�/���`�"O��AtG���D��sƁ7o�PM٥��@����N�8��S��?���Q22�1���8��dK�)�O�<	q"J�3\d�H�E)=�`(��LO?���G ) Z����'883V��%;&��(F�b�e�6��(���e����L�Pdذ�Ԙ��0�"OZ�{P`߬Q*,���oُ��	Q�"O�)��^�q�p(n�5���7"O�'�Õ@:���5)���0��
_�|��D��i N4-ψH�e�<1F�S�-�ZaxVN ��M�7$Ӷ��±v
h㟢|���%�98�$C*pX��bC�w�<���ߘiCT��A�>c
j<���m��<gz��I=rfy0�&g�	��k�������^?vnT���R�J�X�3��ڡ.���
�(D�lcS���0�#���.,��lC�:�C_������ v��i��	H[N���	M� �!�DM�{
l�F�
DG��THϻQB�	�/| #<E���'"XupuO��y�D:0�ٙ�y⥂�ޭ��)��2�h�CƓ���"���ɽ��@�s����!��@��cy����ɿ�Ȅ1��A�j���Ya���a2D�8�0��?m.MI��^"��0��^���D�� �@0�8Pe��,s�ȉ2�jJ�y���8qt0[��C�i;���F��dD����|����a�׀��z��ЊF*"{!��;!"����ַ^�yF��8$j1OY��I+K����h��F��ot�VB��^�2��U�Jf�A��KLB�I,>Ԑ����]�s# ��프�TC�IJub�2�T[� ���FE��VC��0R�R�pv��x����@-D�� �O�ɠ�-%LO�ɸ�AQ�r���`��p"!9��'���3�	�@�^���$��v�P����I�!�$�>��P"���)��Hb�	�9�џ�r	T�O�0�av&�:[�0E�BC��#�'yq�Ӫ�9=��Xv�@;E,�A)O�H�c8�)ʧQ��E���  H��&�[�؍��B\����A�(Go�Hx���.Ό�$�h8���d��XSHġ!��p���oX�Z!l%D��w펯S� (5��
{��`Bo!D�,a�*�_���Z�:,v��(�>D��P �D �@��Q�AC���3�8D����,�nPk��QV�~���4D�$Q��|; \���$��1D�D;3,��6�҉ �M�Y��X�7�<D�0���[6��x�i�(inQ��;D�ԓ��S${����H�&�b��4D����E�J�v��'&�.�.�2�/'D�Hk/Q.��8C�΂{�����/D�x��L�ox0lQ�サ&����-D��#��\*�h`#�@�Q�]�an&D��.m��}��B��rTDy��ϛ0�!��G�"�h�Ig�H�>��,����3U�!��M]Qp��a�C��d�oF	&M!�ۭH��L��[2�xXT,�O4!�9]@���4�7b�6Q�#�:!��M���1C%��$Y�fL[��!�$���(6C��5�
����؄4�!���@\��e�:p�����Ù�!�͹{u������'/z��P�h���!�C�lD�y��b�����R�!�dX�*7�Y����wv,�s�j��!�D_?m�|Psu�Ƞj_0�$�yB!�� pM��͔ebC&FŲj:��"O\	Bd��6P�6lzvE�=M��r"Oƅ��lH�d�0�c�n�Gn(�;#"O����7E�Q��ض���K�"O�IQ�+U 3�� �fgB��R� �"O�d!4�2?0�L�`LF�-�B���"O��ZUbQP<XQ��)	�@����W��bA-ֆd f��5G5����ʦ>��s�ה;O��'uX���3��?]�1�޳wV�ڷ�+LID�r�l�:�o�>d����H�y���� �3�2,˗��'��d^[��ɰx8�1��X�9#���(/}b�w>Y��Lm��87��>�� M8�H�æ�Nf| ���"Kn�Տ��QZ �el�'2�|�h2�'}R�h>�@�l�o�	>�@�qkX�zX�l3�-�����H�e��A��8?51D�����a稄1K�L)�Ƥ�F�*���O�X`cB�f} 5�	ϓ��Ѥ�(M�q��mȁSyLl&�8���ڒ�M3�!�1J��(2ƶ?;t"�B=��.?�����H�QI6`-��C�I�7�~V �BM��'{f�h�C+ǻ.��� 7&�1��6��>�y��צ4�V���?�G3�<���P
o� `�$ܔ,О�2�O��c���d�@���j֡C�F�Hr��6O���;Fd���~r�R���Z3��Q�I;*�6� �O6=��}1��z���\�,�Rt�f�G!Z4�4kA�ɖP���a�.O�ơ���G�X"҄�'�Z��1��/�zĄ牍=6@�6a��]<��'ċ1�
Ox!
6�_�w�.����c�m��O�B�w���}�@)��ց �p�*�O�}���戀bh<1��J�y2���&�w�xQ�F�L3.8�+۸Y��x�5.L$1��Z�S�2����yb*y���d�I
&�)	s"�<(	<Xp�8�O@m��fŶ(p��*u���@áM ��q�Pd{�X��]�4(��
b���(r��l2�Cŝ|rd�Ny�(
�c*P�DU��ȑ��O�q�wNQ�]SP�"�'N�94��~�@���j��[�Pщ F"/vZ$��?*V�!�H�T!�ϓz��Y#�?@-~��'"%����9� h��Qq(в��U7=,����|��]}�p�a�7"{�p0�e1%iL�1�fgh<�!LN��C�S�:���Ѹ]�ra������'���`�9l&t�3B݃�yg#Ǒ(�q����-j��]	�	P�p?Ќ��\Ǣq���]�9y2u��#=�`�+��=�)00�B�^n*�˗�4\��O֐�/H(y��Pk�V�J�\9ه�	�<�B��S�J7�U(���$��6��L	��̈́>y��-* ��ʀ逐\L��O�K^���olpd�P�_�"�$�P��8f��ɤ*~��")�x��0)ᇝv��"=�u"�6&q��÷�W����@A����xr*������A�G$igIơ'b��ņ����=Q��!I��X�u w�%�0f̜m��c!�3:��|��c6�Oz�H�i�8B���E��2&lȰu�=z�*�!��|r�	�~��"��3eK�M�	�E�T�9_EL���fMz��\y��$�*gK3C��[W��s��X�4u<P�n�2�<��jJ�C4P�O��iP����;������[
sխS�b��Ɇ���Pd���.�9���o����W�O�PY����}c@9�eM'�!�$M~#���&�C�ay$�*�
Ҏ���3*X/R8U�I�2* �zT��4$�D�	r��l*«]2t��բ�/�����>dd��u@+vdT���ݕq����W����`CNՠ��\g<��<��N�1���{t�ʹj��(��!�W�'�8���σ#�T��L�NI��c�4~���( 쏱y���:�k�"uN,��'���p��o�H�C OE:= P�*�Oy9A"8�����G16ot�C���O���RG��'J��ˠ�24|X�'�t]I�gJ%|��܊d���i����Fǵ4��U���ߍHƪ��$�?�䧈�')� ���r��Ks��
F��b	�'�D�*�V�p`�'�*�u	�'��Ejqk@;M�.���Z�x����'���F��oN!��g�	q�z�k�'7(���EN!\F��y��E�3�t%�	�'FpY�.N�V�V���Ɇziɂ	�'FDm�ѣ�@g�8�r�Ο!@^l�	�'>����Q�]�0¦S�b] �z	�'��(3CB���)Юˁ�DT��'������
"���,�8�����'��e��΃wÌP�n�1M�|Yj�'�>*w/B6�|�HJ�r�X�
��� b43E��Hm��!Q5|�hx��"O���7ƃ1$e�(I�ǉ�.��Q"O�� �BS���15$�+��ej�"Ov��/PV^�x�H�#�ʑ��"O�-�cĔ+��1��gܧ$`<Ñ"Ox���%tfp�E耷y�,��f"O\�0���~���X�(B�_i6��"O�`��$W��(1�倞�aRq��"OFl)���L�L�R%	 Y�pi$"O(4��,ȁI(.h�6�U�WQ�q�"O���&��*	Z�c��ڂS��`�"O�л7/��Xl��;W���*�Є@C"Or���bT�!��Yb�ϛw�%h�"O�h���PNP���	�X �"O���ӝC����̕u�\MR"O�4�$�H&����� Z��`(�"Oژ�Wi�
�m*���C���"O�ࠧ�ߔh��(��͹'�t��C"O�Y�ï�&����M*2��L�"O*="�NL�����P�Ф��l� "O���T��lӒ�Y�h��$"ODb���-*�lph	�t��I`"O̹�Kӿ���&ע	� �c�"OxE�0�_D{�l�q[7n�B5"O�Xq ���??�L��� dtk�"O��kӍh�l��e�]�����U"O�-�ghP�%'(ɣ�oY����"O&	1+������(w���"O�M
�JY?*��ӷG��k^�a�"O�4���m�hu����Mni��"O�A`7�^ `!�,0�FϷ<\�[�"O,�5V;	M��X�(�8Ĵ:�"O�11��DTS8�8C&U�> #"O�H�t�zY$�ӳ++q�(Q�T"OV����WH���@�Y'l|e�"O��s�"y����IP��9�K)D���ں'���#D�I	��pg@(D�j�L��D�&/z�T(a�E8D���s#1+��(�j&.
Q�l)D���D�ӚB�@�aS���)u-&D����ߚN@� � M��=�h(u�#D��*�S8��!�d�X���i!D�,pB���a����Dյ�A��>D�L��AO��8�&咪P�Aj�/D�1���[ @,3AN�&Ō�E�"D�`ZSgU9Gy�C/Z�fI�P�=D�T0 �C�7�����]�,�0���<D���f'�MR6�Jo�(�Ce�v�<� C�/6��dk��Ǚ>T�����q�<�FJ�te*�i3��6��,TS�<�R�E�,_lۣ�h�ƀ	!ɄQ�<QT��kt�ӆ����b�c�<	fG�:Y[\���g�"f�,y�w�<QM��lx.�@M�!�,�@ӭs�<���V�}A�$3�n��@��lPI�<�c ��?�Ȍ���C̈���E�<��P��4��b����\�<��Z.(
�%ZD�+%�J�9�\Y�<��b�nI�L��n�$pp�x%ADS�<%��t"�����I5.��h�R�<	Q@�:J��ʀ�.$�I�0h�R�<	ЊB<M�����P0:�04h�+L�<�f�Ț�Bc�&��� A
\�<�6ƌ�Wp:�â��2�ȽM`���S�? �T�s΋5?>D��C]�xh�r"O�!@ӆW�~=jG��7��)'"O���� wn�h@FEʊ��EzD"O��&/�w��T���9g)�w"O�����Ցc�2�;p�̺g^X��"O��ypk��g:+G�W*�҈U"O�*�oͶq��,I�*� �٣`"O\��F�8IX��	��Z��"O���r�]�^�|�`H�n�I4"Ot�`��8�Fp�mI:j�6��s"O�=yC'��XPʀ5[NP@"Ov���'Y*9�<��V1I;�Ihq"OJH��N�dH�ـeO0I��`
�"O��"�C}�6$q�	r�H�a "O� ��E���sG��K��yc@"O~�p���V"���IR.{���7"O�	Y���#��asbϞ֎ٚ�"O�x�$��1T,�l3�"ΗJr���R"OBt���_%.��ڑ�.eB4�5*Ox�A&�_�f���/u����	�'�0���e/!y���D� �D��'M0�glP=l��q�nZ�;B��'���v�U� ��HG\<6,� �'jr����
�/,|ah�oߍz>2tY
�'��FEEo6vbd�[�A�.�{�'D����	�Z:.�р ��4V��a�'%�Q؇bT�
v�Sag�&0���'vX�mO7f�a�K:SL9!�'��TP�6` �1iO�zwhUH�'�p|RlǴ��X��iLj�
�'�6����. ��&�,'�(h
�'�� ��Z,�D)p�A*k��
�'�� ���ɋ'���j6��x.")��'@&�"NS�w������0w���I�'L�����@����?t��T��'��5����2
T�q��I�f٦�q�'��0Q�a��xB�H��� `1:<Y
�'|���2O{�����qP
�'�:(����
D4L���}�|�
�'�$)����3E�a37E��r�T)
�'���c%H�I w.m.�t@	�'$�R��� IB�Ɇ��c��'Ԓ��"�	�gp15g2���'v� � &��5#���� IL4�
�'��V��9����4�
.�T�
�'<r�!�]n��,J�d�4%\��[�'EFaمH�.e��D`B��_����'b���@Ǝ��� aA��*M޸�Z�'��R�B�Qrb��Q�ȓ@��|8�'��A�F�
mԒE�q���>�f��'�y����6�J���?;\&y	�'=r0
CB�<Wl���F��"O�ȸ�-�96j�nF<�0��$'LOԍ�`M�K��ē��Y�;pe�d"O�9Ң�R ,1�H/��2�]A�"OZxItǔ?V������i��Q���'�剄J=4�k,�3?�<�B�Ѕ7��C䉠+`�����=:n�����T��C�	wft�a.^ %��!v�^��C�,/u�BIA*S����T#3��C�		s6�d���a���E�%~�>C�I�$]���í�<5�\�i���#D�6C�I�(;ԛ�@aL0 c�#GH�B�	j���2���6�|� ]�{N�B�)� T�06ZzV�1�ץe�F����a���əC�������-���J�k�!��[K��
�Ь0�P�:�o�!�D���d��צ� V`�8D�Ͱ<!�D��`�HlEn�
]X8p�,[D!�$��^C�� �#R�d@�PBWɦs6!�D�M?tYMYO�(ن��=!�ĉ�bXP���#�DJ��*����e�!�!�Nd�p�؉&�}H�o�&"#!�$��,�bY3�ĕ�7����!�/�!���Z�YPB�5fи��͖ m�!�qV��A�6' �F�˪!�!��\���&�\4|�N}3�j��}�!��$DqF\��N/U�������n}!�$��n�Fq��%�2}F�����bO!�$Ԡ$Glq����[�Vř�	�!�f���d�qY��A"��i��D:}y��ȓA--!��V>޴iV�Z77�x����y���Nk��b%B5y�x��ȓ:m.9cg� }�����݆ȓ1���@�

T>D�f�Na*ݦO��=�
h�x�~t�-Q?Yb�#w'�f�<a!���DP�`ŵ:� 4۶��`�<I�E�m�&�Ѣ�[�|��\��#�D�<�"	�����&P���Eg�~�<����-(����G�N\�a�3��y�<q�+G,LK�� &%�9��r�"^^�<1���~`V���W�x�(���\W�<I�!�,0����s���]��-p��g�<i���D�t��)d�1bbL�<!�I,#QR�H�&�"vN,��o�J�<��ˊw��u�1��6�8��QE�<�M�"&=��P��ݺ=$F���@H~�<��-THy'M��w��9HĀe�<�'c�."���7!H9''&�� g�<����=H��H�hN�Nݤ��3�e�<	���?��t�	�+XL��ɓ�EW�<�6!A2$q���p�&h��� Q�<�
��qH�͛s�s| 4��K�<	3O�)� ��EB�^��H�b�A�<i���&"��!keBƎ���#�e�<Iv��/�d 2¥�/E�(%*�K�d�<	%՝?+��s��%�X��E%g�<�o�,t&���O\(g����f�<�g� K�&� ��� ����f�<q������v)�.CzБ4c�_�<���I 8E��
2\�{gl�Z�<�שװI&���L�!%�}���@�<�΅�~5�Dj�m��T�{��r�<)�f�,�pAӚ�����c�<� ��3/:��N@�,9y�-\�<���;�fĪBGڕ �@TS�<�R/O[
��V!�6��D�E�N�<���ǂg`p0A��	@�c�p�<1�K��:�vI�w�3:���,p�<!�"�:n���+��
�k��h��l�j�<��':E9���ӡ�E�Je��n�<�0NKJ���x'�� nqX �Dm�<a1��=JxD ��(t��M���C�<!3�Ƌ^�4HrÅ_ q��sfC��<���|t��"�iU�E�2�SB��c�<�� N
bnj�3���$DM3�Ɠc�<I�G
>�����&\����
\�<9R�۱Qd��P���=L����A�<� �UP�eb�D@3�N�b͚�� "OhM���8����eHB�;�h,Q "O�A�CG��_�����h)v��|8�"O��B��ǜ,�f]ӉƵ[n]hc"ONl��I�y�$�S�K8+1��"O2�5��Q�� O><�yA"O�V��<S�B	�v���~Db�s"O^|�ÂW����B��?"]"O����%Κ;l��R5 ��~~�RW"O���;$%�\ڠ��"bB��"O�t���0q�6}`V�:�d�V"O�\i�.U��b ���[�@0xdz�"O^-jX&c�@�J�I�;e�v���"O b�BֱIP��"��M)F��5:A"O�����'\�^T)�&%H�vR�"O~��(�#z�hY��E�E��=��"OH��6e �wQ�d�W�C�~�~`J@"O�۔���	��'�VHY��"O�Ȱ��2F*��s��;�>��Q"O.�ؖe ��k0�ŹK�dl��"OP�r+R!��aZ	T�����"Ox<6��1c}�}h�f�85v�Y�%"O���ǣ\JA� Q�$ʴ<A��:�"O�1�M�@_��b���=
��)IT"OXx��D-9��nG"�C"O�l�C�Ҷ&<�1�B�7Mݑ�"O
�p���,KN-kV�ŒK�(�Â"O�r��٠\�25��R�,���"O��bk	$,ۈٱ��G�3+h��Q"O�)��³G����Ձ_,��"O��`aM������R��@���"O^,Zd�2�:ٚQ�I/Zȍ��"O�8��G�r�j0Zr��J�̒"O�L2�� ���<�bD�,<�m�"O���gDАEٚ�sQ$D�h�Au"O(��6 Q#"�,�������f"O.�HbD�a�yY���4���""O���G3K�V��&�9u��A"O��A��OI�l�pDH_Zy%"O�"� ��^'"Qz��!t;����"O��d��-�ta��H*�L�a"O>��s=J�XaKD�.!��C"O�spn":1h��4� U�N�[G"O�=�6���oJؑ	��^�<Y�"ORLkaP(c��[#`ɼ����"OT�#i	H���R!�T��-�B"O�\jE�[�O�����4.�Jq�d"OdT�֧ ��X�اg�d��d��"O6�sC�Z�D�K�y2�[ "O&�z� Y�%���Mоp,9`�"O���3��!faHìU*@6̉�v"OT|`���8/�<-�3�K�^.�䃄"OHE�!���ش�儇>I�`�d"O`H05�\LZ�p�ԁ�[��l��"OlF��-��'U�>�  "O"��c�.A��BG'2ҕ�A"Oڐ
%���4c�ĺY.�h�"O�\#�]�=<ĢEѯ}ؔ;#"O�Ѣ��Ki���1�CH�u�z�j�"O1��$ʍ#y�������8"R"OV	:Pɍ7aL��0t#�!<Hs�"On�qd��Y�X/w�2݂�"O ���8!�$]rԊ�R�j-:�"O�q�bĕ.U.xq�����"O� `Ct(�')�t�X�f�
W2�y�"O��k9|O�d���-��ź'"O��VF߁j���p��[�L��"O,���ӦZ r���,N6�ƈ�"O���֪[�:���M�M��bh�<����.��̒G�z}�yJ"`�I�<���a�������h����E�<��l��9���k�J���ɻw�Wv�<y4i�w�|`ˤGߛ��A�%N�<��I�.��MW�Ľ{j�UҔ*�t�<�WbHm6��&�<X��!�.�W�<�q�U4l뼁�& �59�5�P+�V�<�f�Q�I�e���0р�qP%	]�<�c푎Mb��'�If��HVp�<9��:��P��-�D�¬q���t�<A�܏i> ����O��T��
J�<� i�#Tfp)tj5�u�5mD�<9�F�� �k���|a��Mg�<�kQ�~���
�/�l1)��]`�<Ѥ,]!�f�'�D�F0�/���ymH-M�*PI ��#]��q�a��&�y����0� ]��֭#QA�-M>�yB%U�<�p�"�F���QIފ�yb��*�.�	��Q���	B��	�y�j�P��d���
C�Sq�O��y���89	�*�&��|��j��M�y���M\��"`ׇn��׋·�y�љ^��(C֨f��T�2��'����K��iW��>�8���'�=��/�%�
(�7�B9=�M��'

Y��a�Q�L�)l z�'�6p��َ$KB�Z B8w�fyR�':��Um�0Ĕ4�iΛvT�@�'�����)��T8�!��pġ��'.�����G�"\r����|�����'<�LK抎�?�(
�)Y�!p853	�'Hr`0���=c�*e��ٻ�$��'��˔Oִ	�Dp��@�b��5��'ݺ�s�.�m7��B�	X6[�H��'�^Ѫ�ESX-�u@F��ON�H
�'����Z���0�-�99��X0�'H��jrf�2�8ɂ�7B� �'��] �@Q&n�lRe d���`�'o,�!��?�6mJ�Y��=	�'4z�� M*z`�\c�l#։�
�'�4m�3G�>�%��Ol}�X	�'~��Iv��'���3��&L�|��'y�q���б�À�!N���'�0��(��R���}φA��'�\�d�ǁ@`��p�Ü,hE�-�
�'W�	�p��b�J񮅨^i	�'$�j���0sD �+�-� D�U��'�bh�q���-�Щ����P��	�'�D[s@SGh�ԣiȦ�\(	�'KJ�QnX�S� q�L5YBŀ	�'%Bd󆫄�1�X��"V
`<I
�'����u�X+NӰ"׌����$P	�' .�+3���x��̏�p`d��'��U���]�b�HDiVW�����'�С�#d����Ӌx�����'��Ae�ƑB��	�fE ����'�h���ȱ|��転���|
���'������.��h*Sˌ�}phlx	�'�jp�t��9|qV��b��D���x��� �Y��:s8��V�'V\ �"O&��c��:�ؔ�-m���"O���K�.
H�S7]�����#"O��2`��y���xQ�\8�M0"O��D��+����LKU�
�7"Oΰ�F-҈_����&Il�ܐ3"O6� ���S�Ř�)G�q���"O��r$��.z\(��G�?�Dh�"Od�f-��A��߰-,f���"OX\�+��Q����1$ڻ�✫w"O"��c2Y%BT#;7�04�b"Op +lB.�5�0�n	�#�W��yR�^�.IQ�A颪ޔ��H�ȓ`<���é�8v"P���ܑ��m�ȓ7�(���]�H�����؆d��|nbd��ŻF�yB�O�\�������⡏WPR�N��葇ȓ><pD+!ȟ9h̸ڇ���\v�̈́�~H��SQ����p�%sd�]��Q(=
�(ܺ}y!QHp��w�A�`��}�DT���ڜ<���ȓk�&��e"���hH8�oد�����؁�eϨ"��I��&:%�-�ȓ �H�B͞19u0ثI�3����ȓ}�p��ʂ;<��t�'	 ɆȓH��H�B��x��� B��ȓZ@���ؓ�T���	 ���ȓ2�D��U�^�<pK�nJ+Zt�t�ȓ�0�2+���ĺ��ͨȀ=��3)H�H� N:D9	�<5�
І�2�¸�M��<�b��P�Z>c����ؼx#��l��3	O%�@u��8P�A��ϡo%�|��	)^�e�ȓf���ز쇧׶�r�Ȗ�'N�<F���!n�p���Ϳ*#��@�D���=i�-՚�jW�gкI;'�_*( �ʓ?~l�$�I��Q1f��|5�B�ɫ_\H�2�Ӯx2~M"�×=��C�	�+0���Bń�Q:�;���lB�	�|������2�z�r�!_�97B�	�|ZX��nMB���$O�Up���7V�&H�у[ޕ�u�Ӛe��L�ȓ1ڴ�D�E�(�q���R���_�����\;;U�%�@��G+v,��v>h�"��<D��kЏ^E��\��:��݂��@W��laghRQ��WNb�p �"M��� Ɩ�%������T�:tO�T�.8�I�6���ȓ�:�ʐ���hh��Y�aT< ���n-Y�#� �z�#�?nBz��p��Dh� �Y��s�o��R�L��ȓ~��!B� U'�����p�����b��4�P���m;�	� �^�ȓU��`��鞊[�:�+0��/d�^��	~�����u±FʌO���S�"i@l�J�. D�<"�I�}�]�"%�fV!���<D�XF@+(����Ĉ�MX��9D��R͐�CH:��*,g
��9�2D�����2<#���j��F(Cs�,D�@y��[vn=�G��ȣ�*D��+��M=.�8"a/"��Q��+D�0��פ��d��ѹQ������<���D�?)�6A�/VAg�!ZK�-��7D�<�ȥvvvA�CfZJE�����:D�� R�9�酨J��CE&D�`Eh�"O@p)�K,�$rg�ˬF~C�"O�h�"��,c�zq8�LQ6G�
�"O����R	L���˳���q�"O�H�F/�#I"����ʒ�V���2��D�Oz˓�O���e�Rg�������2Y��Iy>q2��� ��=S���1o�,m�Wb3D�@��ES"^}�D+ßi��`�#>D��P��z�l��H�L�.\25�&D�L�F�KK��K��+,�jLY�?D�,�\�%tX�k�=wn�Q��7D�@�����T)Ä�0�lQ��6�O�~����E�3L'Z��O������\~�fPS˄��w�ߞ	
��" �yb���D�*�2���7y�"�C����yB�M�P��ӓ��"	΢�2���y"n]�1���P�Ȍ~+h4��j�y2D�9=K4(s#z�h9��)I��yίP�r��%�Cpט�C������O������9�����ڄG!�Fb�� ���3�g?� l��3&�,�qIÂ#>`d8 ��c�<��ň2�t5[d�B�=�0LӇKb�<�%N��G,#א��,XU�<�T��f���J�/M�8���ÅDg�<���'^�<�j�M��V���_|�'�?9h��H�"�*d�@��BL)��?��:�tes�k
�lG�8�gF�1��a���'��'��)�3}�g^��	�2�ʝg�>�s��֩�yR!�?y��b �+N����h���yB#�F��Z7m�&A:����y��C&l���ԩI�d�� 3�yb��3K�:�h6��z'|�p�3�y���$i�,���l�)���s5���y"��F\p�s3��%��s�����y�,V�|Q�䂆!�z@`FP�yr��91T(	��M(�ҥz$oǬ�y���)v|)9��T�fHp�����yR�L4F,�ڑ�Vd`<)�'�yBb�4�Τ���\��PD�%�����O�"~:u#�T=d`��! ��[1��K�<�q��95�M�7��^q���IF�<a��wknQˠ�Ϥ�ε��j�g�<9���`�"Poͬ�� ����<�@F^�C�`���I��q3��|�<�D�	(ZI�xp�k� Q�� @�Cs�<��-�M���8���nEX�Gs�'�a����l�D�F� ( `b��yBԔN��`"�-M)��vN���y���>AQ��[6 �?֠�f�y�I�"⾑����7�\K���yr.S�]!f�3�.4���xL5�y2��v��c��-(����h���ybN�9@�p���V,%�T]�犈��yR�H�q��Agm�?@y'�^,�y�$��c,����j�.��iǯ�y�/ݼo^jh�g+ә��A��n���y��ح~�) cH��W0���ʰ�yr�A�
�A�R��V��D��e�y��mS!�D�ǢK�(��a��y�H%�"ɛ��l<�4Aa,Z��y�+���lQEd���QhP��y�B13\���Ɛ�]k�pr�C��y�n�)�� ��U1��R�^�PyrNL�Xrkū}�=x�a��<� �I����^T0�A0lM�	���"O�u��h��%�v�#�D �L!{�"O����Y{o���\���"ODUR�#ފ,� �@I�$�:q"Oԭ�!6d�԰1��Ϗ_^�4c"OȜ(�n��Zk�/e7���"g%��d�<����0|�E �&e.�P��B�=`����/�^�<Y֨V�b�h`{����0KPlHW�<qcd�g56�����T�r�����{�<�F�ΆA-T �ߦ:V���Nv�<FdA�%�y�䈁�"y�YF��q�<I�lѕ6� �(5��Zx5*q��j�<�� or��䄝Ŕ���O�<Q"]wqȍ�G�1;�L#��b�<�-�*{ֺ|J�B1R�ܲ�H�<A��:>
E��bF'�̕"w�ZA�<�`׷}h�Q��9�<�K�{�<9��Ӄ��$�ϙ�c�B5X�F�tx���'u���ҋ�!;�.9ib"	�Q����N>Q���)�	5x�5��(͗Q���ꘋ(��'�ў�>��ᖾL����\j�0z��"D�xH�Ȑ,��%"ч�3H@P$3D�T#��
9�x`���)P�l	a�2D�l���L���ё�
-p6��l0D�h{5a�!jr��B4E��Y�(�O��8�UPy��E�嫆�W=��ȓz�w��<��q��@-L��u�'��y�)�O6x�3g! �b8�%K��m�F��"O~����m��݉��5*�v�(�"O��O٢RJr�s�H��/���C�"O���A�K�
�F/L�8��"O�P�:m��5����	��)� �d?LO����Ci�J�K͟d�<�BV�:LO����� L�5�������Ɨ|��'��Oq�F�ޚp��1"R��\�S�"Oh<�e�ݎ��<*3M[:"�����"O�8�� ɍR�6�@
�cF�	3"O���M�ZXU�2I�0iDZ���"O���2�B�"^�5�0r�RL���<LOX�2��(d�ҽKsj.7����4�I]���'��q��9Q�F�u���t�+D�l���׼N�<�rem����(�($D���1!J"+1��7e�M:�\�"D�3V%όz��"�Jّyɰ�
C�%D�x
�"�xۀ����	��@�� D�и�fw�)� .P.^�j#�<���0>AU"�Xi���O�gG�hIT�|�'�2�ɂU+ޙ�"�յg�v�`��
V2����@�~�$�Z�}�p���S�]�P ��/���)��*U*��"�s��<��(N�O.*J2�k K���Ƒ��C g�U���	 <n���C� ^�<	�C���Ю�
V���rƒq�<1�G+mm�LY�/I={����!Kn�<�IHUX��jС	�8��s�m�<��Ĉn�� Ι�i�"��%��@�<�G��vӞE`"N�5t���~�<9�oD>D���J�eE4/�(�k4B�p�<y��ջ Y��zv�[2���r��a�<��JT66t�9Pf�!���`%\�<�ӊ )J�yע�J;bi�0��Zx�`�'�H�0	�:s"Da��`�f/V]I�'�ڹ��bV�WH���Ï#\`��y
�'�����׵ RP�hI�B*, 
��� d�!Dп��� V�/kHh��"O lZ�Ԯ0{��PP-�D=sU"O��K��V�p�BĊA�N�-��H"OZ�mE;��<|LH"O>���HD$\K���i蒜k�"O^�A@R�}�^\�S��;]�,qf"Oԡ�3 ��}�i&�Q �ưÁ"O�Ur��[|0�Xb)��D�4pY%"O֔��R�}�0�3�n�'v��y&"O���PA� 6>�#ż
DXy5"O`=���2Y���f!�>?TP���"O8$�@�1\zf��R!�)N49�"O}���U�@��Qx���+4�c"O�%��Z��~���tz���"O��"�O�bH��xe�[��rF"O"�qɊ�� ��Wd'���ID"OΝ�2�.K0�X}�8�"O��f..l38�ʇ
P>-��u�"O�QXC"q0��p��?���"OܱrG,�3ha�4a�:�K0"O�,��ᚹ?��쁆`�-2��lA"O��#�_��@�˔L�	 {��	�"O�	+s�s���j��ϺU0�Ac"O�5Af�WV���o�:�T��d"O���DaO�&����j�"O�����G� �\�C�ުS�zT�"O�)�� F�	;��BâV��`���"O�` �NRWB< Ea�(>�^<�"O�ѱ�!͓j�x��
=~ ��3��U>�&Β�<�� �$}R�Bf�0D�B�g�"΂�ZH �Ql��ǆ-D���Gi�Q�R,��D�mӨ�T@>D�����{���H�O�_^n��n)D��ŅD+U0��zP�c��Cdg:D�  t,j�}�c�M�#$*���M:D�0KQKM�@FP�*ը�'0<� #������O"��`>�ѯ� S/����7gӠ��g�<����Ӳ,�ȫĉ�7c�.a��ʉ�)s�B�I�1���bE)ߠE���D�`VB�	�O�	�GdOE�X�vƌ,v�B�_Pb�K`Bםf����7BLD��B�	(:�"@{%P�t|��C)@�a��B�I2��ł�Bܞ  yk@+\L���??���B�W�������  P�!���g�<�5*7T���ˍ���hY�j�<) �$G@�!m�	xQ��Q�<9'��7Oc�pɶjF��VQj��������jzT�3��f�@ۗ[�*��`�ȓ_A�)� ;;�̸�u��2.y��qjbdC��&6 p��C��%��8�xX��H�8x��;� ��2�'��F{��$C
6C�i����cXؽr����y���:\�e:2-�"^;��B�FO*�y�΀�cb�iP���3\��U��g��yR�W�t*�mLTB
c����d)�Oj��ĉ��HNݑ H��1Dl�B�"O�qr"k����)f�@�L��8�"O�e��ʑu���zG㍼g�E9�"O�sd��/cl�$RYLS����!�Y� ���I7'���0��ڒ7��{�󄒛s�,�j�d�VS�
���'	a|�b�.[�b%�@�V�E��ՠ��Z�yB.8���Z����f��BAަ�y��#��|�1�_=��Y������>��O� (��+ѭ}����s�p�7"O<���./dY�� 1��R�Bq6"O��!P��0o��IT+B�L���[1�'����@<���fҾz���kc�4i&6����?���O���P��M�I�����H�\&8�L>q��0=I���:S���e@-x�bؒb�w�<A C׊ٛ�S ȵ v�<Y�R����"d=�� �@s�<��D�0h��Ҧe��"����5��i�<�@	�(���q�U�wtd�	�G�dx���'2�,�d���p(�'��'���'�F���kU�iG�y����t�npy�"�'��Kv�B�G�U!���`f!�
�'e�A0#�v[-L��m��X�Zݚ
�'=\���H��Y;�E�9�2�Y�'V9pVǆ�Q|�P҃K�5���'�,e#E,ɳ��ْ�Ί�*�L��'_$p1#�>����TM�� �y��'�L=
�3k���g�����M>	��F��hӁ#Y��᧣\�;�Q��3^��"ծhȂh� #X�(<�(�ȓ3����Ԇ''��h��*]�
��ȓfmZ8z��ż.��!�L/+�t �ȓ[�6�p$�U=v�tĂ�2+!J�ȓ`(`��KО,_�|�A�E/b=�l�?����~�`�C4MZ
� � �5n�
Ђ�j�g�<y��͸	��u��.f��0L�a�<�A&^=)A���V΅i_ܑ�t��a�<��,�A��)"����%��T�T\y��'����^�: dp��ǿ>_�(��'"��I�	%��5+�,W�3�h�'�����ȏW܄L��&�ּ	�'"6�a3��%d`�0YՏ�+�b��'H��H���4CK�����	�}�H�'�����
R,y������E��ܡ�'�����-O�B��݃WB֗:S�4+��?��#�J��0�0`��� �cֈŅȓ}0� �*K�K�^��T��k�a��w��`�LP+G1hA#��l�`���l~���1
�,�C�^e�#'��y�F�O5�r�X�}�����H��y���X���E�r��Y�޴��O�#~���ln,��Ë.I�8M��a�<�q���� ƾ �� "��]�<9vH����S�A�hob|��GZ�<a�D���"ڦ}��p腢Źk�X���!�	.�4���'��Ժ#��+:�2B�	u����H�1t)��c �#4C�	�����/��k߼m�t�5E*0C����}a%�[)w��%�#��|����<� 2Ϙ�ql��#�1WP��F�.D��`7��9����kW;EljH��2D����S�p�����攅R*���"���O��؈���� ^c�h#�/_-#�Ab0"O�����%�2��M��]�}s"OFT�1�	�k�"���`�`�A"OL`��B�;���b�$.ָ�K�_������^N��� ���G$��3�h�<-�C䉟C�ذE߂L�du�T�?+C�I�)$<��g�B\p ��q8C�!6Rm�f&�u��R��
G��B�I8Vd��V�EP��iK‟//�`B�ɃJ�&IS��3y��cH�|2jB�	;`;�٫�fD�X� �X�n�p2�B�)� j̲e�R�O���r�P���qv"O�KU	�{�l��M��cE��[�ԛ�(�-"	���!�F�RB�XCE �Ot�I�>yX�{��ZPL���[�O�C�	�2�r�i���S�6��C�+5	�C�	�h�j�'jwd �L�-$C�	�;����G����e����W��B�(4/P0��F�J���@#i;C�I' ���E��D�H�p��>���D.��O��?�'���k�%��2rܰZA�T��'m�"d�0Y�aW�ԨgY�ua�'D��	� УR��*E�.X�A�
�'լ-R��S ����fK���-r
�'�� v�ӗ
�
� �;;�|u 
�'��Hk#�ס:Y��
Ǯ�$�����'�R��� ^*IS�l�V����)
���?����S�O=��Pcō�؛�bX
,-��S�"O(��l��3ʆ��e��qly�"O̍���P6^q�I�ǢA1*h�S�"O�����9T\F�J�-ZY�&"O����=1͜Eq5��z�q�"O�E�&
֘C5n������֤�s"Ob�8��<AӶ��F�)3��\�'�O̢}��<�(ᩦ��pJjb�EƝp��ȓgb�C&�S�9 �Sg�6h�ȓs�f� R���sZ`�A�g����s��m������uq�)Y)�%�%D���/E)cO0p0A+	.2�<�A�Oz�O��S�O)ƨ��U�%�|)4߫-�L%��	���G�4�B5~���ϊ/��a��(�y��	���	�,�(w�@ba�X�y�	;M����Z�Ξ�` -���y"k�
#XP��A2�"e���:�yR�]�J�Jw� w}�Ղ�ؗ�yrbFwj��a�Bo�4��pg�6�?����?�����>�'�>/@X���h�C�]jA�E�'"a�ԭ�P�yґA��`TyPt-�y��ã�051��YdL��@����'6�O,���O���E�p�LT�z�P��E\2B�	45l}9�)�<x��e�W�kPB�	�A��d:dj��d�xB$�p��C䉤?�6T���׀Y�"�lƛX�B�	'z,����S	fd�����Q��B䉅\u�	[�.�*�~�P$���DC�B�.�@� 

h�PZ� ['t�fB䉼:qRm��L.U�Z��A��"B�	=U��jfD�D�C��J�)�HC�I'G[���7�$3� ]� !��
pBC�	�x,$�F��	.�0!yw�Ű,
㟸E{J?ՉI�"ӄ-�gǒ& A赢�:D��P@�B�>��t�'��u���D�4D���e��H�kD,Q,6�%���4D��y��;`ʕ��H��1Cr�?D��ӥ	��08�#� y)�!٧c9D�(B(OK;�ˀ��+"�����5D�tÑ�Q #q<Zg&�5L/�43��8�O���(vq���eE,&%jT#A�x˔��D4gh�8��H7>�
� 7��>-�-�ȓ8��Xr�Ȍ�vl�Y@�E�b�0	��}i0يb Lg�����͝ ����C�\ĂL�5&\�[�p��d��씽�JS/�2����D	PA����$�U�֌�!K�*Q�`�UPl�'�0F{��$oB�U����J�?b�U�˜��y
� fȰUJ��R�h)r��W
!L�)�"O��膇&d���d�,Zi2�"O�@���M�qJ����B^ ?�	CE"O��9a�C2�vՋDKE��ـ�"O�@��(ܯK�3�I�D�B�@""O^��t`R~4�@bh#14�d0�"O�iE({e��*`n@'̕s�"Oܩ
C��9dQZ@C���|8��"O`�z$k�7L��MX���&k
�$��"O`��A�D�x�y�-��D����"O���o�)T�=H�m��aΨ�u"OP=��ҭUZ��a$��Fy�Cb"O.�re�0�	� ��>gn����&�S���?Z�)T$B4��Ś6ɂ|��'�a|R�8{뚥)fg�Yy��&�y�� �v�V����&c�M��_��yB ��zL��8a�."�u{v�M�y2'BK�t����)� ���"��y�J(%kv���ՃL!�D���y���4�z�P�.Ն��h�4���y��,XN���� kHd��C@���?)ӓi���f���)�hۙB�h����B	���!���Ԓ�����	
���Lҧ3�x\b��JO8`ć�e*A L��nu�%�a�qm>фȓ90nEiW&��H *V	A���h��gb��Ã		(��������&����K��P�v��)5��xU�5݀��ȓ(a H�6��z\f1��Z
`���}נp
ũ��)�� P��=�VD���`5��K<$�E�� ��c|���+���rN�<���F.�/!��ȓ_&*�	��
|�f9"Sb�
��q�ȓ2���e	'mh>�iĩ�=*Wbh�ȓ�""��#K�T�K	��ȓR�Ht�ߖ$�=�qG�粙���D5��đ1_���`��S�XI��?�~8����p�(�H���(e`l�ȓK�!��A�l�ր���Ur~���s\���&oĎ|*�= �� ?��@�����g�@ϊ4��
�)x��w_�%���;Nv
��bxkT��ȓz/�E�&nA�]�����-C�'�b�����y�OQ2�-s���D?�؇ȓ3�P�K��`�Py9B`�l�����d~89���J#q��Q��π:�t��~�2�ꢣ����ef���.,��=� 	����B�B	�OPz 8�ȓԢA�4�>�����	�?[��1�ȓl' m�Ƌɶ$�Rhc�*��)�*x�ȓF�N�r�b 8B2\��푿W�R͆�j(����ų��и��n�L�ȓ&7�!K��xܮ��	71�2��s�0:B�'���t��cԹ��D����4�1@�Eb4��x۶���;m���G�Bf�9��O�zXTX��]2�(P%d�A�8��/ǘ,��̄ȓn�"��mЌi���u�0��r]2�h�·
x����d#�}Ԝ�����R
�,u``�ssGJ�A��L��#mXd��<�.ɹ�ͮu��)�ȓqA�E�A'��R�:�AGm�,E1 -��`�
dfE	�U��I�kکL�:@�ȓ\�`�dV�s�N�wH�1m���S�? �-2�坡D`��1s��UKȸ�f"O,�9gb�=]�,`$'��>;ZLh"O2�V`N4/P�8xu��>
3ԁ��"O�Iq!RQb�ׄ̐#3 �r�"O���� 5.%
��'S���pG"O����
��� ���P�f¾$�"O xإ���\�<���ן�R���"O4L��L�>wC�5sAh���¡�"ON�;%/�<T�x�e�����"O�A�u���*�0�ÓG[�I7���6"O0�#ᅀF�5�G�<J"l��"O*	k� �Jn��P1��6hg:���"O�\	���<��93Ė9[�6H�&"OBȲ$ ��;�(�b����t-Z5"OE�e�� #<,��p�N�huh�"ORY@���T��TR2��.5wlLkQ"Ov�G
J,�pô�ĞC\҄�1"O
p{0B84�f5�bnT#d�,4��"O�Ϟ77h�\��Ǌ~�H�Y�"O���M�+'��pǂ �Up�"O"��	��DS���@Xv�`�"Oڹ��$Cl-��C6't�y$��`�<�3�ßw�%;���34�n�aE_Y�<a�h����a��,�� �C�p�<q�鏦V�4��똠Chl`��T�<4��=F1\d��M�=JLT�v�O�<���΅+�D�#��� ���p��H�<A�͔z/�Xs�J�Q���{��D�<���>#�Xu�kI#��ms���Y�<	�H��J�m�gH[NVTK��T�<9�m��b���V�Go c�OOL�<r�=�Xuc@�?l,�J1"@�<)p�X�M��F�"=� ��L�@�<!�,%WJ ��]#n>��(Q�{�<��X>�H���N�X��NOt�<���J���y#nU��Jp��F�<Q��Q7x�~)�F��RvA!�Sz�<�unǺft۰IK�JTH�ʦa�<IS5p������J�R��D�PY�<Ѵ��d_n- $�Bf8�۰J�S�<1�BшD>�	���$��H��NL�<	C��()�!)vDU�	4�9Y��E�<х冑-����c��=�B�A� �L�<���;_��A��m�1��}� .MN�<5J�i����Ùd�<��HG6S�^����~�Jmb���`�<Ԋ�"�8��Q�K<|����B�<�u#�+)L��MX�e&�{5.�<�ud��вv%B)�h����x�<��䀤uO1��N�{����'Ďx�<�")gʾb�댺+u�}Z�ϝ~�<���0��1ԯ�B�Ny�7�v�<��"��O¯8F:y"��
W�<�`$I>(8v)SD[;�.Tr��T�<	�A�)��iC��
Z��0� �	Q�<i7�ʍa�^��Vʟ�M%�@�GF�J�<)�Fo�US7��4w|��Am�<!���P����/�Qi e�e�<A�bдf���%e�`�Q��`�<����\���N� �TI�Sg^�<�@Xs�d���&�����e�<��B.V.�2�/�/o��A0��Ia�<�#J�8'S��%���Sdi��+a�<��+�<���X��	�8$ir��^Y�<� �e����5)f ��.�{�6�Js"O��at��m�x8���]�(h��"O���� K�_#�=0��C? �b�"O�|�"U�p��(���{jp�@"O>��m9&$bE�2 �1Lf>�p�"Ou�*�/w@F�ʖ�Z>%x�"O��:�E!+lx[%��7�<��F"O�82��/i�����Z|�i�"O��jlӂz��У�MU Q(�"O~<iQg��n(<��֣����ps"O�Y+0� �#1&�P$��=����"Ox�קZ(_�܅cE�@g���"O������r��9 s�[<��A"O�Xg��}�D�#�\���"O��'-��T�Ţ�
S�R'|��b"O�	��iG�rH:��f�Q"Oܰ�ЊK�2�d����ƂG�8}Ä"O�sAF	N��ћAE'A�za��"O\y�ш�2g� ��I6x���y "O�Y5���C�G��Y���S"ON �)L�Mp�ԛD쉿|;^ԙ�"O~|�6��$w	�s7J1DX�TI�"O�噷+B(D�x���G�!��"O��X��@��J� Fʴh�.�h'"O�)�NT=��y�F��)�p�:�"O�����<PT�I�?c��4�"O�h���3Ö����\�ot�*V"ONA��lYsYk c�-g^*S"O�(9���$h��T*' <QV���"O֥ʣ����m�`N=�����"O�L��Z>�j|A�:�.ye"Ol��F�/5�!�T!��\y�$Q�"O^`�֍�N���9���"J��C"O���gR�i������ I0�c$"OH��D�2N�t��
J31�"O4�iq��s�l�`EǡI&��`"O���V,�4r����t�]��i��"On$���FWƩ����4򘸺�"O��:0AC�E!PC�1.�����"O��%��n����Ā�N�buKa"O���D>F^	��ҡ�􈋗"O<��cg�4%��EK�i��� �"O
�W���: h���SH�����"O�4{�&V	�N�b�#�'`�|�"O���2���B/@ ����.~!�Ua,�=r��#md���_8-y!�S�:���Q�g@�Aʔ�-!�d��J��ՒA
D/�)Sjԇ/�!��>k�x�@�Us�����!W�!��4xs"�Ϝ#ew8��fR�p�!�D�O��CA+T�F	�%�Q��C!��¤C�6|�vI�#7bz�{���u!�D-T8�ۅ�*Y.i�b��4d!�d]0t�l�V(��+J�5*����d�!�DӨ#��7�
�
6iz���!�䏴ͶuR0kZ8'��GJۉ]�!��ҕ'�`�c�*R�}t<H�*�G+!�^o�.زS��
�b�@�i�J/!�dB)8d��+�ܭSVG@C+!��$����g���B���f��h!�D֩U��xG�	]�>�A���/w+!��!
��S�П�8d�&%ţ{!�d�,�DPjr[56��![��Q�!�dJ�}@�1�l)x3��rg�l�!�� J�c��[3�i
��K?_@�[U"O2�C$d��J�dE���O�uA
�QU"OX]�T+�05v&)��3$b%��"Of�2p됄df΅���[�vJ3"O��3f��/�4	g#�_�:$W"OX��S���;��LG��`W"O�E���qȠ��r��5E�E"O֬Ҷ���
[�ɲ��G3l�x0�"O��4��W�<�"B:Z�d�"O.�2�*�G�	�RC�q�YB�"O�iۗ��?��{sE2Z���q"Ot ���?g�|E��FP�zA�c�f�<�V�ɽ6���
@X P��z�<YGd�Uװ�{jPV22� �Ru�<����<2�ƀ\�f���H�ep�<���D ���֓D,��H�)Ai�<)4�K�Bk�\#`�(G� ����l�<1�d0��	 i�/Vl��@��i�<10�S�Ⴍ�&�'.*�yq��h�<o�nݮ����S�D��0/a�<A�GKO(F�JΜ�Y�q�BI�\�<I5M�*�z�Q傄=\u�8D�@�<�DL	( O,�)�'V�y3����_a�<bO@0��$J�o�4*T��&��E�<i��[>,�۲$Ո+�����
�f�<a���]�(Aj��)-:�*�+�_�<1�#JX̝25�5C%���B��\�<��#<���a�;<n���E\�<�d�ƀ�j .��+{:�0\Y�<��d�.������n7���*^U�<9�%I�&l�)��	`�PہP�<�+OX��tc�f,F���K�e�<�D-Y�� c��ݦl�QӅFLd�<�h"b�ĤX�A���8�jǉ�a�<����0),4��c�=h��(KI�<مI�7cV �ಧ�-z�Z֧ D�<��ݙ(o�ͳ@܉p.��d�I�<�a���ʀ��1^B �רW\�<�OE>,$@�#ZD}��A�h�N�<�3L	8%�0�å�w���b�J�<��׿q2�q(c�
z.(	� �Q�<��]Q��|(#����3�O�<�*@?d��]3�aT3P�t1�t��o�<�S&G�9и�Fʓ,3���!-�d�<�0k�({��u"�L.+z�Dʕ��d�<�gܷ5���Q�E5m�\W�k�<Y�B@�E��AA�k�/?�8 D�g�<iP�n>��� �W�����
|�<�L�E|�V�ĥ~2��`(Py�<QN��QU�ɛt≤g�V	� ��N�<��#�z����"<O�����a�<��)���4�E��:�j}K��G�<!f�� �\�q� �wjL�s�B�<p�іryd�%�iLC�<0l@<�`�
���zAh��S�A�<�G[�\���Ѽ`wl���	x�<�c(�9O��
�@�T��yI�mN�<"���\n�1�N�0_�.da�)�K�<q�(�!}�J(�u#�BƊ�R��H�<Q�jڿ|�e��K�$V�(���F�<���F9[Q����'AY)\����B[�<1��B�Jk<�)"�P�}H�@ 2��A�<�r�Ɖ=^8�B.���49�C`]b�<�%,S,t
��ao�_��-��Z�<� �X��L;9�ּ�$��x�L|bR"OD���FB�y�$$Z�%4����T�<�diO�M�4�3B ���3�&�N�<�F�	aB�!���X�����c�<ɖE^�0�X-DM/r�>4�j�`�<�@��>�2���A)`/6��	�`�<�Q��l�� ��EIl��F��S�<��#G6>�|qI��&]����ZQ�<�!ɞ#Vz�ek�j^�P�ޅ��.�I�<�l�7C��a8q���S,��~�<���>�!*�O+)����w�<I�b<<�rD�P�I��}"�Gt�<YTgͥ3'�cc ^B���(�J�<Q�d�j�"a��^��A"D��H�<�'mO��PI�+�)v`�w��^�<	S��$q���`�%Ɨr��Ct��W�<Y�i�5&S�(��Њ �ӑk�Q�<��,eΪ���j��u/�0+UO��y��N�~1�F�*y�ƐZ����yCT</T4щ����[��I�/��y�&ِ#�!!�@�T�ک�
�yA�9*����˚-OGn��c��yr�B���1D��*�2AD^5�y�H >%����xH�8�Ę��y��[�`ף31`��V�q�!���x(�Zd�	&q ��v��!�!�D�1U����e`X��5� ����!�D�
k)NĘRK�0�8`FZ� |!�$]E�&<�. ��|m��J�&p!��&)J8��"��/V����J/ �!�D�gf�C�a�)9BA�0L��ȓf1ȀK�R�*k�AYvkؓ�X��ȓK�:��^.^q��¤n��.Y,ԆȓW�B)#BoA�^Ɔm�,�2��E�ȓI�IR��˪�4�O�`���ȓk�9*1E�&�&���R){����$[��1"��:� ��$ЫA�0ńȓ�����N. �FK�d��t���\�y"dW7g����&�4�����R�0X���9NVUK�W<�P��U�P�(�� ʤsB�"MW���ȓ'<z��A�CC�x=�ua�c0���igйR�S$�P��J�>��u�ȓ*�, 8P��3&zƀ��(K�/@��ȓ`^~xH��G]$	0��)4ײi�ȓ0��S��X� 	(q�%��<�Q��Q�����̍>�^eѤk�R�r�ȓy
�i��J'
|���O�@$���$�����ǊT�,��8� �ȓy	�U�"�M5pP�d���%/Їȓ~���K�o��yYB(�A�L���1o��OAbp����5|�d؆�F� �Z0�R,!�I[�FL/J�<��(n��U��� w�	d��ji����K�$���h�%z�����5{@N���<��Tr׀�p�#�ծL�d�ȓ.��)��!H1�	��b�-d2�-���q��8+~�|�����S����<�0P ���u����.����ȓ
���f^�����#<F&��	�0�ض�N�"�ͳ7�����;]PD��#��j��s�)�J����8���H�2�V0�v��!-���f�<���n�bkP�"�ܭ��S�? ��Z��̂� )��B�6�V1�"O�e��ɂ>-ܴ�BCuzr�"O,���h����!_�T��"Oh-;��2\�H�� �J�X P�"Ol\����Duڐ�F 	]oؽ�#"O��ē�J��Hh�NX<�-�C"OҩS!�I�cO=qS��47�r�X"O�Y�vk[0Î�`'Q�	c����"OX�r�e1��R`�S$;b�i&"O:��� ��o��t�&#�QY�[�"O�KG�MTy���AL��"O�hkD��kǨM����#�`���i�l�Gy���iݔ��9�		/O,�.�	�'���B Ύ�,�n�jv�[���٩�O"���?��w��,�� :M�U(�U���I:*�L��H���p��_4.ͲX[7��d&Y�ȓ(�ҔBɤdU���ӡڶ4	�E{R�O|�[!a�N�Vh�$�ѱl�X�	�'"�$ReY�L��L ���h1t܀	�'��c�oD
��|�LR�%��@	�'�(��H*� �D�8	�1�H<�
���S��ʱHZ8y8r��
�e�� @MڠN��i���Z�k�(9����ȓL����ނ	e�!ѹ=�`�Dzb�O����A���E\�1P(���O�1s>$���X�5+��Y)�5��ʟ�Ia$�mjy��)��,z��D��,w^"ݲ�JO�m�0��D�>I��4�Ð��t�2Dse�K\�<�e��4A� ���.~�W�'��?�jY¾��I|j�|%�&D��s��>��xR�,N�����J&D���Q���sk U)�o��A���!�%D���ס�0�*�R "�:A���82�!D�x� -�e��A�	�|�{�:D���ֈ'yfq��b��c~n� W--D��N� >���B�J�w�*E���&�����'E�n�GIG�~<��Z#lD ̄ȓD p�ÜG�|�R�)�c�h=F|�	�|`˛�K� \ҭK�qg�< � �_�<�����YsGlE���<HEI	Ϧ�Gx��O.ўP�B�8Ih�$x��E��-�0��|�<w��+��c�+\�����dy��>�O����%x���!�',���͋%�B�8I3��)r�	/����Ȇ1y�B䉺+LtD���_�6#
������B�I�V;��K�d��M9�F ��^B�I�<�|�%��7���r��W�V"?Y��Ɍ1D���� �}ZXhPa˜t!���qD���Hؙ[��	".�"!�$;1����7�P<����#ڵd�!��h��g!R2�rPz$�X�R�!���i^���n�n�1E��c}!���m*Ib�9?b6�Y��1��Ű>I@g��2�:59��הz#� ��@GL�<Qt��1M��IѫP8-!DRb�^�<����iь�Bp���>c�A@�Z�<Y�-��L�#B��)�"X*���T�<9���Y[brI0J��E��X�<!0���D���h�<4��Hc�ky��)ʧG�^H�Q�?\j����' �p���%�����H`!�O�j����N�t�B�	��2�C�&Z�.L���W5f� C�)�9+�m۪Uf��+GrA(6����OTP����|nZ��1�Wc�6*� ֩4'pB�)� ������9;����ΠJ��A���i���PX�L5�rdL637^�
3�i�a{��Fq�$Z`ڜ�C�	-v�Nh����5w����h�Qre	�k5��.�G����0(8D�h�%HP�F�
��g�Ĉ.�����$6�o�?A�k�L ��k�H��<ء�w�2D�P�tN8V�0���̄y���aC���D{J?ݥOjL�t��~�88��5.n�r�"O��R�F6����#SoH}�ו>q�V��?�J?�)�صoM*���6�v8�j+�O�������n�'ql�j��DWW����+����ʅ�p�V�� �����Vh�ȓ>8�����-�����P���ȓ7�,�Y�k߽���V���Є�^^�9�
-z�E��	Mk�N���U�D�',�
P.dx!ēI��)F|2���>�`A
�!г?"X��`�OC䉹a>X;4nٔvI���E68�B�I�|7 �ڒ�	.b6ڙ�0�B2?�B䉪,�4��t�I�/-���Ŭ0+H�C�I�r`�@c��Z�*���\!��C�I�K6�5�M�nd$ ���N�8|�'Zў�?Ua�E�#5�h%��E\�ҼȠM#D���f]?���xr��Fd�(�Q�!�	}؞1���`8��W����P��vĜ��=����$͘� !"-������y��zB�D��J�<��A�O�f� ��2>��@E{ʟv����K�?�&
�(5pݮx�"Oz��b��&��������h��"O��9�ᝆh�
 BS�)#�pc�'����9E
�#���:)]�����8��m���17c��C @��ЉӮ%;t�sB3D�Dj K8�Zp��
_7_T�Ð�1D���Ц6eczAzV-@�kV�{��0O�"=Y#�K����=J\
�/�s�<Q���"6l�f-`��@':�'�ў�?%kQ�@���1Z
�^�(@ �?D��S`�s)�"��#DY2*?D���臞K�8�E��Bu���>D�����k��"jΊj����=D�`Pp�7w�PP�h�?��"�l?D�ԣÂV�t���N'R�� ��;D�x���ҺP�b@��� �N,�p):D���&rk6���NQ�z�.x�6k3�O`�ɍ:'pq�a\�	�LT�`FB4C�Il�\A���H�~<Z���O�c�,�'�Q?��P0��g�&�1D:D���qI�.xS�90��V���B��O��=E�����|5[�
��#�Q���$!!�d[3�nc"
�q����q!��npX�������y��� es!��[?����jϳD$0R�C'e!��>L������ëlӈl�'��gR�|��x~�c��u"�U�b@n�)c ��yB�
�	1A�#_2~�#
�����\�dEM����(	�~ΰX)aF����S���0>Y�'_�	�^��@W
2��a�uᘘ@�\���<)�'�phק���D�@�<ջ���C�4�(Q���`�!�$�F�uӒ��%||���΋|�%����	g�0�׈��+���p�퐂p�����9�ɹi�fEKO�xhddL�,��B��Q�U�2A��0������G!_��O^��ô-n�`���@�>u��)��ۺ�!��O��B!Q�PAAF�e�.�1@"O� ���ƒ^|�]��O[�1��A���'���O��s����c���H)�0�:���ȓx�,\����lĘ�e@7$o�q��	9m�\�~i���I�Y'J���i�f�{6�G@S@�@B�X�E�8�ȓFT�+S�N�n��@5�V���ȓ@R	p!(A�!�u��&�-�J���`)���
O/쉰�iÕh�r��AH���w��)-�T�'������ȓR��s���H�rqATAW�$�ȓL��%뢭ٌr�H9�OM�m4���7>:9��'��6�ja�v�ӆ}7JM�ȓThX�Am�_,4���H8A�*��ȓD@�a���L�H3���� ?��-�ȓ#�`�a��.a��{ց�}l�ȓ]�0���ס9��"�	+(�I�����[29�j���&jX��t�H��J�t̈qGQ
�<%�ȓ.1̽j��W�f�����oK�A�x��<���nB�v��P��A?����=ά��㎥7����6�H�A��͇����#����^�iĨV�i��a�ȓ]���r�K
w��u�TLB ڈ��TۤQ�7�%/R"��:1��1��b�0�Y���
r� �{�ܝ�ȓr	�-B�[�>���!�� �7R���ȓ.���ѵB�"Q��$f�X�V��N�fq��>����d
����ȓz�}	��P�N	��O�E�rt�ȓs?��[�k�+l�D�e@�
d��-�������3�MS`�<2�4��0���8�(���ix���,h=�ȓvS��Q�]8+	2�� !�&(�Q��X�q4�Ayx����:����B�zl2��į�R!94��+:��.m�E�G@59z<	e-Q����ȓ]���S�ꂐw��(V�͂D ꀇȓ@��*�&�>s�N	��o^�vF=��FSZ�b�"�mp�� h�2��ȓ�D�P�j�(�ܘ�p�F�3��q�����悉7:2A`�H�R�����O���)t�/D�ڄprN�Ț4�ȓA�&�ঀ��	FU��O޸L����ȓ>YLs�״ox0 sAc��	�'jıgD\;����W#Wlj�]��'=`�xfj�7cʀ, M�!x��9�'��AKV�	��z$�G-_�y2~� ���53B1xqG�W��Y1"cJ#:!���O�,�Q��?�8�$�)!�ą�YH�Y1ȕ+���W�̞3
!� +X�U�0��9�nA;�!�ҬQ�A,��B/�)�O���!��W\$<�"jڮ,��Q�ηH�!�$O�d�p� @Eĕ.r�3�MU�8�!����L�g�@���LI��!��� �R� � \�|�� b�C�|�!��^�
%�mk���|�x�zQ+�DV!�ė+wfʽp�F�D��)���0!J!�U�{�jSC�G#���x�:<!�$��QP�h� E�}��4[E��&!�d�^��(q�V��6�"c!��՚���q��� �Y!��ʵ1� ��jǂP�HYbW�\P!�ĉ�BWj�!U��y0L�y"_�QH!�$Y87Hx��TKR2������H!�� �|�Q�ן �������`�"O,�z����IY�!*AÐ�ℛ�"O� ���4L�}	p#�j���ؤ"O�<����&��U��C�`"O�����],Q���
P�l��"O*yh���S���v�['J�R�r7"Oh�@�����:��	Ta��h��̑���@�&?�;���&l���09(��
3�X(���8�'�p�r)X��,8>l2Q�is����>��>��OS��x�/�"�ܒ�)Vd�<2�¯���h0��xBP!KeK�# �(�ځ��v͐7�'E��'�=<C؅�aV6nqR��w%|��5�ڞ���4w|,��h�Wt%��K����ȓ~�b�(� �Q��\�B�Sfr��=1�I5�d�C�k�H��%��T? �\5��NR�ʒ"O̡[�!��Z	���]�%@2,�"�9B|1�@	@y�lK}���D=P��%"��*Eb ��!�T��!���u��P@I� t��S�� f<�xW���=�'�p=	#�	V�j�[���$�Tp�FQ����,H7V���!��u'���P�w�N��ؚj5R`�"OJ�2��
*�����_�\=�ea����.��,��B�-�X@�g�iĕs���S'Q�"H�B=f!�$˝p�,�B��Q��[���:fA��1���/��!E����sF�<iU$׼n�<Mp��8k���[7/@S�<�R"R�7���󠘍��d���('*m;�Kλ8��X���\�ay��r&��J�$8�8�J��4�p=Au�N2H�
Xƍ_?F��	S���8��QE���������1�x�&d1ҭ�G9Jnix�����'�>�#5�Ew$�Q.DF?��`-2�F\����)�&W�ZUk"O���1fG7$2�˷�
"n�$��@�9obh��yl�(�	�x
Q>�hC��Z�@R+3�d-����2S�0��BG���] L�r�*��/�̌#T�P�/��-��)��g ��1�'Ū�&Ǡ]�HY��.0Ϙ�hדRT*��v�A�d'H	sSQT��R���z�ih�̟96���Od��Ë�p=�e/:LL��#)eԐ�U�{�$A~�ٗ=f��$�G�~�+l�b�S�+':
�R�A&9��������!�$�9��!�C�*�Vm�&,����Κ? 8\�"Y�`I� �u�� ���:�)r+X�1�fy����NҔ�"O 0؅�\X� )i�nԁK���X�i���k���&!k܅�O?7-�GW.�
T��%@� g�09A!�G�D���-��$��BP�� 6�ɇn�� ��/�y��[�q�����
!S-Tػ&��;��>�'��/q�Y�a.�� F�����7>�^�y'L[$9�B�os�԰%dȎU��| pl
�o�@"=1W"�?Jr�*b$'�S�`pl���3zI�@� �G5"��B�ɧf�
�򆆘Zf��r��F��6��S��,3�+���)����F�/<�y٣�K�K4,�3d�,D�@k��rh��I8I�x1"�!�>���N@�a���1<O�9���N(~`IHO�M���'�ۂe�=#�T��Ah�-��������"��"�|h<!"�HU���v#ȉ�����\D�'�&�'�J+�zm�B�
�n\��Y�<�Q�5�@�<Y�$˯wgp���(4:��X�ɟ�j7�W ���&�"~�%A�Q<���H��LQX��e�5�y�E�a��s#Q�0;���!��?�H;6q��#^@~�Osc�#��)r��dY���P��@�>D�4Qs�>ihd�����xl@�z��>Ac��$/X��kד[NLp��E�j�$��m)c�%����i|\��'=������S�鈍lyrP!c�Q�%$�Iv,�9O�d��`���d�J�3$� D�����en�M�s�Y:;4��KCm��(Ett[�昕?���S�_;6Ў��F�gn���|�<�ҁI�Nͨk�TiX��Q�����'�|e*U΀8I�օmڍzFAh"%�,���dQ����'s*4�AR���$���?<�,�3a��p1O��P0�S� NE��w�,�D���F��(Y!���Mk���Wph�a�Ȓ�|*�m�o���d#�6��%��㜆2�����N:�\S!I�r��� ��ptiB�W���fɗ�n[��@��B�>�9 eZn�x����P����XTٟ�d�DK_����B`+�@�Q��)U
|Q'�G�Q!�$�g�`q��W�W�����(D9��� F�7[fe(E���]�^���o��b�zu��O��bT⍞��C��J'
N�{fc��9�l�c�@���=��/�<�<���J'#�aS�A�a���,+Y�,��6��"�&̐�~��1�܀�5�Հ5d���<�C�ׅ>h�!������1�o�?��ܲ��ݭy�$
��5$����.��d�vl��T��.�>4���S�y6�)��W
H=V%��C����6E�#|(�7�,mj����DC�lU!�'�|�,���(C8��e�?��V�6�T�X��\��S��>�`���qNpl�NOO�<I�c��\<�0��!CxDT���G�1&`��cM�):�I�gd���� �o�|��'"�dHDcg�y��C��X�U.^r��XK�.1�O�%�Bm	;�?1g�5H[|���*ߊ~!б@8��A������'qh-�v�KN�'� !㗃�r��A
��T�������ĕ��Ub��OzѣDɨ`+\˧�"P�)]�H����OR3D���7d�YH��Lf�0��'6Yw��cfXW� q��'pvi�U��z�O���8O
�arFȨ4`$�t��D�!�L/!��i�jI�oGP����%^2����|��e؞ q�Ú�|?�h8��M1
�򸲳G)|O� � ��(=q�4aݴ!j���SF���J��G@xJh��ZƉH�W�m������i�d��?ar�_+��+��9ҧ�����	%t���P�J�]��G/2����0#6�Ó�>S��H[�b>- ��虦��F�O��n�$��`z�Ǔ|�"�3��!���"n~�"�i�yh����!/�~%
����D��M���QyZwlv�bT)�d��XuqS�T�4nq)��Y�����I�3T�}�kI����H'{������7r��a��Ն�~��J�����ME��Dh1-�X&�HJ�l5R���CE7c�����ږ��DZ5P���S3�Wжtb2�ܖ<٬��6�Z�f�H`1+���xr"	7!���d�9aφ8h��۾X'�x�1≟�����T���b1d�H�L�u�<��w�+�·�����`E�� ��'��B�̪`U�q
�ˍp�v�X�؀/S°26e_�"����	�H���/�|������6�d��G!zC䉼�8��H5l�VC�/�4�S���1߀D0У�i3��l3O���d	
^f�b�նg��7�'�޸hՍ�.��eA��$��P�waD5�>�!@�)0�d��A�U<I HM�F��d!��4h��Q���R̓j��aԣА��88t��H�H~2�4#�E���ڵ#dI�%�H�<�)�%L��h��	:Q��1���D#~��q�$`�3C��#�ؓ
KF F�DQ�h3DŅ�r�v� �˜7O����C�(D����C�!BT1�ո:��yJ�̒�_9>��$D��@��#HY&f�*�Gb�
|G�2` A$!&�X��Q��0=9���>F ;�K<=�D��"��-��@�Z2y��t�BQ7)wfA�
�,D��c2U�k����D7v��<a�F�G?b�S��<5���_1��'o":8У�̱W�r�[�Γg�t��W�-+ALO�PA3g�lI\�B�`Y0Ȝ���)6p��}˦D�n�O��I+:����,��{!�Ł�$��<�ZC�I1*r�����&Q��اČ�W<��_�t2DJ�əyB���A�q�'���ᡅ��zU�숛.��rד_VH%��J/`��B�ǞZ��ܱ�`�-:,-���	6h� ���l-�@V��$^8�3&� �~��N#��I<�ds�[�.����B��0�1��1�dѢ1vP�H�!-����"Ob��E͌. V��ƨ�,l
(��;^���:��i������>�Q�]���ɽy�b����O�)`�y�ȓP���m�;)3n9�� Б{�No�BV��Swņ��["Bo�I8�,�1l��Y��hX�!P�>��\��"7|O �����4((z=�,G#�|�K�mI�*�&d��#ԝD�Z1��'��J�E�.m��jȸR�*�(���C��R�� ����8�B�:l�!�ÙnvN��"OJ�+4N#5`jx2����:}���5�'�64Z��g�S�O��<c���H���y"��<uHV��"ODquŖ}?煁5���"Od}��oA�X���B6V���"O�}atM��@���G=6UH�"O���eI��YS�b�X*l�r"O� �ق����?L�ܠ��f�`��"O�k�)U Q�tY��ϻ��b�"O�t�W.�d��G�ˌq�l��"O
�yba�=H����NӼ`����"O��Sr��4w�.�Q�m�S<d
�"O����V9F$�#�*

��x%"O�a8G��7�E�PB:E��"Oڝ*�"=���&��>�bQ��"O��/%���)�'��>gް��-�9�ybɂ
y�p=�I�zb}�6�I�yB�HX�PU8�gǁgWz!���^��y�ib<� ��P �`�Ͽ�y��*y��$����C���u���yr"Ǫ �� 6l�.F�֘�$j���y�e��=�N�7�<37��r4j���y���[��jC�]�����N�?�y�+��4�J��P�^� ����ybF,�yےM�g-FD��揫�y2���>#�8��Y$#�u�I&�!�I��$ȳQK[�_�>��a��pd!�$�"	܀�A�Rg���y2��?^5!�D����d 6��JVĉj5�Y/!��Ljj�*�]3U�.abb�A5!�$]h0����UX%�R�' !��2w��F��'΢����7O�!��^7��ps  <;PJ���F�e�!�D�#rh r��bչΚ�We!�$��-��#�E
X>����q�!�$ۄ���a��*A�R!^�p�!��N}�r���/[������	 �!�d�����u�]�W�����,A�Ix!���k��`�S*d#@*Y1rl!�D;KGL �D�M���2cW�^I!�dP+BR����Cl|�ZsLӠk4!��K V褉¬	w_� �і`!!�D
�A�� `�/K]X��'E$E!��Ǣ�N��gF]�4^�-��|#!�$Ȯ@�0p�r`/0F*�A��[�:%!�$�	A
n9R�CH�x��[2�Ћ&!�A'Dw��Z��ά&3� ư[!�D���H]�6jN��M�g�	!�H�D�8���@1$�a���M�Z!��U�f�!�C��B"�tڒ���
�!�� �!�@�"�	��$�h���w�!���(C�t�ct���pMA3v!�DF�7-�܈�e����-	-���"O@�Ca-T�9`��a�D< �"O��6fW�S�DAq�J� ���*s"O�%��2����.�1����"O��#"X"}\�`yR��>-1b"O�,��]�"M^���K65��"O�F	�3xÒ�Av�]��r�*�"O�I�2(C�.��WH�0H��y*�"O��Q�@G c�A��gL�C����s"O*p�G��;�6@ � ���,�f"O:8�Q	��P�c�OUm�$A�$"O6��`���b4i�͉-v�zu2�"OL�`�W�_��$�ƕ�6�Q"O�a��W�z2Ѳ�'�b��iBb"O��A����~���(�ń�f|�ܳ�"O�R��$�`�\�*o����"Or}a��O�k0�� #�M����"O�%�ah�y�`�*����ZK��z�"O�4@��!�"X�a��h(~�Ҡ"O� X!��OC����">$�P�"O܂��Y�~>8\yAKM�S��)�"Ol�Q��v�� �Ȟa��h��"O(p9`CԳA����\l�A��"O���̨M4ɡ���J_���"ODh!��ď\^QD	lh�*�"O �"�cE�HI@d�s�3%#^X20"O�W���H����u���m�D�<9�ʡx���G=i�j�H���x�<a���+�!��̀90"pXC	�t�<��#[Δ��WAV�Kh�th%
j��@iPUcǘ���~�hQC�>P��Z��&$���"O~馅ťaL��V�48�����fl_RH:�D-}�-�g}��4j�`��rC@�r���)�!H��y���&-�&DP'���� b�Ɉ�wz\d����5r,�Sp�.lO���q�^� �l:�R�0@��'������+@tsB�i�ӈ^�-a
T���R�}�f�a�'/����J��pZ� �o�@��{"'�2X8l!�4��>5
 ��7Re�}sn$�n���n"D�P�w�5��Ԣ���(a韷~���1��,���%�(��T��a0@c�vj�d��>���'��āw���D����*X�%�&���	�{=Pɩ�DK�K��q���(,�icB�IFm� �۳Jl���F�R*`�V,���J��w��${�,I��\�T���)���y�� �<��o�"C�2yYs����'���	o����-��!���O���G�W��달'*��'cV-I�H�V3بS$�A���U�gW���c�G@�D�0�(��I7^�lM	�Fք`��T��� �`9HC�I�g�(Ԉq���%d���ghߦ>�h�HB��D9��
�}��}�	�%%*0B7�
 Ԙ0�'L1Vwb��뉈7!�i��Ԟf����hB��0���0V��̊1��5%�LI�ēqZ�\P��Ė1Q����Cį"Z��=�qד�P���dC�j,������,2J�b�r�DBP���+5d	 �y�Β-s��'aI�g┛�,�($���^-v��Cv`�OF�ʉ�Y���Tm 	60h���]�0����$D���#g	�S����=�B��@�?v��j�� YG�y�a+��<�qk8(�� ��خ�\ez���|���3�냠T�R��A��Z���Ɂ.��e�r��7�CL��!��O�_}�KԼxd��VO�x��J�~tܱےhɓ*
c� J�J@:\-�BՋ*h���&Q��U<C����
H���&�#*N0��'gm����%NX1x�T�(��RP�\CxqJ�ĕ��$�1�8�2�kS���'�yw �$o��ȼ��z M��yr�D2Yڔ��鉉8a��;p@K�M[F�K�7:$Qg,}���i!Vm�PMo� �F)�5��uY	�'��LPъFy��p*f�x� lH�O��ӔR:6�V�sϓ5k f�#���3K4<%ti��	�j^ت4�#ar�m8A˜4{n (�g]�tZO� �C�>�5@�7@��xp��	wV�E��&^�j��`a�@ �ҌTqbjJ*����"O�	���?c���I�Dq��F�iC���6������>E��4�f�q�E�@ >��e�݅�;�6�� ��7=���i�
U2h��4�'_��9�MR��I��I�E5��Ӊ� o���ǉS�P@H����=����7h� $�8���6�Ҹ���Q	1��R�' ���To<"i�BH�?d���������pa��-����OX@X*� �w,�ċ ���e��)��'�$5K`�f[��mJ�C^��P��b h�\&��S�O	�Q�V��<!͒�ܪ��	r�"O������t����%X{�Z ��'�^�[GkL�p_����O�)l�3���a�I�^di�F�ςr�&��ȓTN���t�ԛRY�)c�C8U����'�ڄ�"LH2�zRk��'�&kPb���d#!����j�*�1��؄	��RH?���e[��1�倗�P9x�	�(
�6ǄEK���.B��8��3E��W\�HB��P1ULDA�o z1���s��7O�$�F�S}�O�$�=� `"�#�.\�D�LS��'xD�qT�5vdn��o�\d��
A�/��<H�I�&�8���E�*�����0!�A��t+�dY���_b1O�lS���R�0�b����;~����$�.V�(P��fT�M�p���RĸŪ�|�S��R7:�A��
(��c��<G�X����&TH>�0�'�R�����	�\�p�i�l���*�����H�ЉU�'�LY�ʛ��\���O�h$��Cu~��C&G���	f��7��1�+�y�`�J�>�3�*�,1�4�rv�B�@�Ѥ��;d���*SO�e�::d IN�<��'B1����Y"CݢG/v��hISl.��Q�]_��|�����)C]�IrL�@O֬7��C�JDf������r�P�P?1b��:,|<���W��b�t�Α<,��J:f��!4�#��4��U�v!"{<p����s��	 #�X�|*�(����u�c���5.)@2����*�j��9` {��2\O�}��8|q����M��N�9��!��c>��G�_�<�.4�� K�i�ӟb��F��&r�x���{��ݑkK�`pW��G���'*D��8w�?s��uk�"_+���!H�v/�3��64
>$�i�88�Q��~�˓�ty˰4��cb���Јb .3�����'-��`�k�ǟ�0�D\�.�	�!���H4%3O���"N�y��Jd���'"%ғ6� ,��ں#�ni�Otʤ�Dx���h�H2�'F(��ԧ����B��y��q
�|Ґ�·w��C���ӯ:���SA��6;ܴ��%Qw�4����l����k[�>i��x�P�L�� M���ȓ~WN� ���>�p0��0���I@N^԰s	�"3�a{��@�ӆ)P1aI;�=��Ǚ��=��JQ�(f�!��`����#����S#X��r"O�u[��@�k'(pie�Ŝ6�H�����jP���_��H����P���d��<qw�ި,$@�"O�d���6��$��M];xj9@EG��
�t`1s��B��.�g?y2(� Y�������B}�I)��W�<Av��V��`�CO5 ��9��֟�Z �	S2�L#��'�*U�&瀌v.���Ŗ�F��iZ	�\f�QT�'�(7�0��k�DW�^�)`&��.!�U�,��kW#Nz�Y�&�(C��%�C+2-\�G�tGמ2� Tq�c\�B��ZA���y2�D�2d]� �ΙO�4"1Ѭ3#J\8cP���������7�z���?��9�7���y��3�Ia�!��+�DD�w.
�y�(ȿO��S%�>,6����y�dP(&�\�jc��V1�EPJQ��y2�\9;�Tm�$a�7M]D=iSlK0�y��Q�h��q�Q�Ň9ݚU�B���y�C[60�W`��4���n�y2�^5�t$�*5�	R,S/�y"��}1Ć6�4��D���y��(xܲ�P�-	&	����+�yr���Z�ۓA̹VjB�;B���y)�&}Q0UCJ?F��	��'�y���,�pt�ɔ5/KB����]��y"c���H�D9��HW쐤�y���2G��D	��$z��]�#�[�y�*��i�&�N$F�2��Rϐ��y��
j5���C,�p�"�L�yB��<��P��f�0 t��邬��yB"ȯ6�đ'�Ps��#rc1�yB�;�\�g�F@~�RWoX��y
�(�6�Z�.�&H��s'���y"�ڽA�2!k0��H�R�C1���y�J	%`�*�y�	�C��h1�D��yBʘ!��X���
��)pf�8�y2hP�$���c�q��@P��yb�Wl��&皉P��|��#R�y��]�"�e�2T(y����yR!��v8�#_hpa ��yb��KĀ"��޴yA�S����y҉M�~U,)�����zŨ�5���y�����p��Y~춈��� �y
� �uaK�-���:�\�2��W"OlE�n� �Xs͘�~�Tq�"O���G�Ɓ����,�d�`���"O����ET�d�l!�����RD��"OB486ʊ$���C[�*Ę�rb"O6C`�M�̛b���i���Ys"O�0q�ݶe�
��%��/����W"O���g�*g=���o�'g�)R�"OD��V%� +\qsဂV�20�U"Oz�ae˘�m3�I eG�rў��Q"O�)�e�x����������"Ox���NO���ɥ�&co�0�B"O�$�L��i�x��,Z2��"OR�tL��x�L�ygh]6�Rl��"O�A���H����ڷ�HS���"O���A����=�#��:j&Т@"OR-1�(�f��d�QȅE����"O�ԑ@��<m� �֏'Cxh��"O�z3n��ښ�0�"*�� �"O8����#�]a��8tՈ�s"OxͳG1?L� ��#Z�[��r6"O��C��O:ld�E��W����""Oxx%��nlz�p��J�T���x�"O��:�%@��TU�f�L�%ل"O*D�d0=�
����_�])�0e"O|�Áf�Z�!���>@R"O�!�-�V:ڄ�bo�EH�"O\�����1D���!Z� �0"OJ1�R�߸z�`�@��l �"Ob��� �+9I�d�C����"O�qPPj�S�4��;B�ly�"O�l�Dh�~S(&�EL�8"O�U�G��n��E"� _
֜��"OzD�G � �*I��]1��l�"O$l:�/��h����^��<�!�]�`)R�"R��
s�> #�
E�va!�^%�h�X2Ƙ�EJ&Ē�iM�W!�$�o���QԤS�(T��NY��!���s�	V��Q����Cv!�$�1;M�9���D�J� `�=h!�d�&u{",H���D��<�P��OW!�DŅ[�p��u��$a�����~�!�5'lpy��{\���
�s�!�D�{�"t�i²<�"��뉑n�!�$��~(���p�{�<(�E\�l^!��R�T)��b'G���Z�%���!��![�]+ƃ�/S㺩%d��8*!�$�"T�� ��SC��\��ev!�X�_�BY���P�XH�&g!�䑿&��BE,�F�� K�Z�qY!��
�s���v�H#m��8���^�'f!�DU�%jhB6���#�diq��� >!�K%"��Q������J{@aݽ`�!�d�"�1KD�L�>��􆂯,��N��Z��dRN`6Ĳ���-����f�a4��W�|��+�N7D��cP�7J`����2+����4D��)��4���J)�<�#-D�@7�Ǟ��Q+�斜M���h-D����y�z�W'Z�tUˠa6D�t����*U��		6��\�B	"s�7D���#�Ne���N_�~DQO(D�,AQ��)X��&nY�T�Yf&D��u�F;+ ��F�"�l�w*O䘠5+َ{}^�9��O�]y�3"O� �=��눽K��Ԑ�����5{�"O���W�ߘ�m�V��'w��c�"OZ}��AI�7�b�����_h�q��"O�iS5�9U����;>z���"Ol���d�"+��J6��M�^mY6"O�<*�	zn��P��	m�ڍ
e7O��
���ض��<E�DX�'�H4@��� xA�p�ڱ��PsR�t~x-��W��Sa�*�\!R�$�!���d ������eM0
AN�H4�	�>!�a���-(�LJd��,4V�e��#^݊���$DH�RC�1[wH�0
�' v�Ua�ɆX/$ ���J&\�pdr��v��h��bB��`�E*V>Yd��14:kF�(�٫�IEǸ;�g�!S�d�����=9�"|�/��ru[77��L2��N�Y���J� I�Wf�q{#h��#M�`�5��/
��;ҧE|iH�*ۂe�f)!4� �4��0�(O��������|���O�ve��G;q�ơP��$v�؝'n|�'N\�%a(IrW�"~�Ub؛K3pa1�Z�1��+�Q�<��*y��)��eA^�NM �\c�<yF��~9�y�!�^6����&��V�<� bM��8;�jD�
��PԞB�ɯ.ߌ]y��>@�
T��Ye��B�	'~�����Q�=��\fJ��@B�I�=iR�
&Lz��C��VC�I�p}z����/E�~\��-C:�B�I�=�r�3���+-�d+��M�|�tB�*&Fܸ���U����(ʟ��B�>������/�<5�i:A�nB�	T�x`�l��^R��wK�6�B��4�����6ܹ1dF�>e�B��1���;$�S�S�L0s��RMHB�Ɂ��4��£W��e�>�*B�	�O���b
M�U��j��7�
B�I�r|T$r���hQ����_��C�5b׊ك��F�t�zi�`�5l�8C䉚"�6����P�TzPQ�d�W C�� n(b�'�Pjm�c-Z�B�I�S�V�£�
���RP�[$J��B�I�)|���Ӈ�C��T�%�S!(e�B��+��6��.G�D`s$@T",�C䉾|�=!te�Kܸ/�`��C䉔֠�SUh�K ��@	�$
��C�I-��6�L,<p��AѾ!=^C�	�w;
YxT�L9�b�:��O�u�@C䉥B����.�1	l��A�4b�8C�	�]��H#O'9�iI3$��b��B�I�AL��ӄʕ[��А���UǞC�I�}�8L�宍i�B��q�ĳp�B�	�'�|�d�%!6T�VD�	�B���4sӢ�{�4�0$��\O�B��8E@h���K�B��و�фHy�B�I�X4��i�.��KU��a򍎭�B䉧x@���D/_�~�X������b�bB�@3,`�%��
AV���݀��B�4�أE1ٲ��ϗ*N$B�ɺI�y�4�RQ��Er�����C�ɃN���D-G�h�pɃEm�>c�`B�Ka�Lpbf]�n��Cl�dvB䉦:N��锦G�<M*���ZV~C�IVjΉ����~�,ᢔ��&C�I[�����Û�o
����<�RB�I�M��E�@+���
q���
_�FB�I�!;J�0�GK�L�:���d�
f�xB�	�7b�CV@�C	1*ô81�	&D�dj��d6|x��M�k#���o&D�x!^�'פ400��d�@a�6�'D�đu�E�j�D! �j̬)ajt9d&D�� ��g >��q���1p�,��e"O�[�O�n�hT����?N�"Q"OF��N�$sX�W#V*YR�I�"OH ѱ�&~ �Ԁ�Q�M�hp�"Ot������C����`�.�R9
�"O)��F̰E��Ms4  �g���m8D�D�����Y	�`��V���d=D�L�m��˚����OD��U�<D�$[�V�MY� �x�f�4/'D�#qI�bs�%p0��j�.1P�i0D�,S�"�	���3CM�>�y��	#D�0���˧<j-ZuoP!<�x�B� D��(�j�pd��t�Re��l��E4D��´@�["���C�Lzr�cr�7D��9S�u�����ͺD�p "V�)D�$���]�h0�taË�z��s�%D���D��<X&�H�\@[�D"D���S�E���b�/y�&���%D�h�p(>e�©��KƩr� �Q5�$D�T�F$�yG�q��F�K��mn�/D�8��-kt>}s#
CCjAJ!,-D�(�6���#���a�e�)lV���"�,D�D��̅�8�q��-vde�d(8D�D ���O�>@QÃ�9ye�0 g D����UÄ�#����e�Zj >D���c#޶6��` PLL�B���t�:D�$k���&˾ӢM˭=4��ks8D� ����>�B��*v�|��J D�T�.ϓ)��a���',°h��>D��h��(~�kU#^9LlN�6k>D�|��8p�<A��)Eqp]��:D�RE�ȖV��a(`�_�3�0�Yb�:D���(�<��٥*F̌��n>D�$�'��+���&�8U�Lhz�C<D�d+)ϘK�\Kb�\�/Z�|*5�>D�t�qEѿ��%jQ��V��:s�7D��0�GuE:�	��Ъ&3t� �5D��{$��|�	���-����&� D���A�R27�B��O�o�*�[�`<D��Bp�˰}!�(�!G3;����%D��R���.f�@:���G�
��k(D���B�702&����U��5z��$D��9��L�E;����#� O��Y�D/D�@�3k�8������5h�5�_�C�I�]bl 0�";d&xQ2dM�x�B�	8k:j�*�b�_."�P��B��B�	�n2`16,��7y�Ȉ$�?K�B�I*g��9r���bh��B�/PN���'�Rq���L�;%`���7Z6�us�'���qlʹgr1�"��Zf���'���3S���|%K㊟+.Hl�'�ڹ�Vf�i�:�ӑ�0><�
�'�a�SP�`�@f�ɪG���
�'K\p"�G�2�u@g��%��a
�'k�� � �����Rh�p�
�'lj�kE�. q6ԓP�� �'��4�A@�oǤ<�� \�+9��0
�'�64�&�u9��r3*
�c	�'���:���|R���|���'�4���Iρ}y,բ�IR��J���'VSRiݖ%�؂T�����'��X �ɻ�8̘�mŅ�6�<D�|�UC�-����cN'8��b�4D��
��':D��V�
<r����=D�� �lxD�Ţ>4�Hh�_	C.�	r"O6T����S1p1��� 	y� X�"O�Љ��[�a"�d�p�O�7�Q�'"O*I�1"[�a��0�BO�*��"O��p�+W�&o\��Rd0zD���%"O8@�@!О��hC��ɍw@��3"Ot{0	�LRVY��aO�#���"OHy�F� �_�h9�*�-r��Z�"O�MX�aΦF>��p
�e^�9k�"O�Tz���-[ؚiSY(q��"O���ˇ�R'��!'�G�9Z�C䉼h主p�[�o{����"�VODB�	�Mk�x���Tc�+��B�IO#���)o��<�bo؄�BC�	�4��Ի�H�XjplsGL�5UC�ɈLȉ��j�8*�����%��B��<BL���G������k%�K�EΜC�	"+W�����Fw4�:�I��bKZC�3/��y��.?7"EI�k�drXC�I"=ve��V1(��p�Q�8D�C�	�<��b(� 8�V�S�A"3�jC�	�������OS�q*��]�B�ɑ}	�er`��?s$:�KP#?�nB�	��� �� ��	�LX��L�&anB䉱M[R)�'a�,d�\	�!W!!3,B�I1��z������eƎU94^B�	2R���{�H	�2�	e�2��C�#*���xC�^v�"LK�ˑ"3N~C�I�r"*=��C�l�b�1@jQ�R�PC�I
Wvx(����'e�����h<"C䉁;O�|�W�
v=�Hk�(ou C�Is���2� ��nE�DJs��b�B�ɻK�LU1N ;����2 ���p����Ý[O��8Å�1mb�0��z�(�a��ǩb�l����ЮE��ȓ<�haT@�3s�l@se��}|�9�ȓR'P���G2L��!���L���T�zh;boЍ.O��c����8фȓtܐc�/�:|�����`���ȓ':Z�ar O'�vq�Q�J�@�� �С��c�6C<�i�f���'m�!���n�`�ņ ��A�_y���^��h�O\�D��у4�[�$TՆȓc�䡙��Vy����O=jH�ȓS��E�������!S�[|��ȓ�	U��4"��l�� 7IwH�ȓl#���d	T/a? SUOZ1�ܕ�ȓ=��DjAl��@Z�z�n

���B��ԣ�e�>b�l5'-R��:�ȓ	)�2Q"҉ ��t�X�a*�Xi�<y��D�y�B����&D=� �d�b�<)�Ɩ=LY�L�LΤx P�\a�<IŠ�R�%I fH*0����"`�f�<A#��,�6��w��?!�,�a�Kc�<�U!N^�P1��DH�.�`���t�<Ĥ' ��PR�D�/Wę��Tq�<Y���,<<XP"�+�����o�<q�(׹v���p���/,T�+�D�<dQ�ҹ��Eɗ-6����I�<�'9z{HdP�L�+NnR�� @D�<)G���H2J��]*l�� "��T�<���=T�t!�Ɗ�Cn����(�h�<�d�
�j�8�k2��wP�A�Y�<	��րlq�	r2�[�s����F	T�<� *�ć�v��(����E\��PE"O~�iTK� ����V��<{X�-1'"OFxF*�.]�d�kk	+HG���"O�1�n.Z�b�'�-5E��"O�8�*�:3\H��D"6 P�"Oޠ�n^4CV����d��[�)J�"OZ�$�@!�X��0ʋ(Y$421"O�M���4hw�P��8Kg��"Oȃ��\�J���>K8��"O*Ԣ��Ii�b鸁mJ�uJ��X�"O�{Eι����6G3��"O^w��*�·�W�|�Wb�>�y� S��,��%�(U^"� ��[�y�Cv���K�Ƅ}�.���!�y�OwlJ�C��g�D�Q��%�y"Cڽ=���D@�{�h����3�y�!�3LA�db��0o,�U�P���y�΋&8�� sL�=k�DS L ��y���+���7\N���Gk���y��\ v 0  ��   �  a  �  �  8*  �5  �@  FL  �W  c  An  �u  ~  !�  d�  ��   �  C�  ��  �  B�  ��  �  e�  ��  S�  ��  �  T�  ��  ,�  ��  O @ x � � S( �. $6 f< �B XE  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" �'\1Oh�����[!ҰzEn��
:�"OF4��� \�lq�\:�"OL8#WB�"�̣��;�� C�"O*�3"�h����&e�X8�"OFx)��6z,��
2��"O�T�0���9��젴+Na:s1"O����"M3蜻UA��#I���"On`��j����2���1\�ć�	�M� �7�_���4AEM��h��B�ɾn�^����y\���
�a��C�)P�� #s�Y(;jѰ7A$&�f#=��T?��s��3{4P��ӵ �RK?D�HY�!��BQ0M�ƈ� R8,D�s�7D��
ј>�b�����_F�3�1D��1��~<zxS�σ{?fe�O�������lhQ��Um�pЕ���c�"���=T.d@`ƞ"%���an�
W�P(���&{��U��Eq��Ŀ\콇�;�#��a��E��D��?ZpЅ��؝��A(dHY
t�?uZ,ه�\� �A�S:H��nI�^`,�ȓW�y�)�"�ݻ#!
�*�>L�ȓ(�ݚ��RS�. ӢY
aٔt��+� Q{C�2>`�+RǄI�>��ȓ:��i��1� �E���A�<ц�p��u�4B\��|��ł7g��ņ��BeR�G>/l�Ԓ�b�5E.�la�����V,��Aul��1�F����<�y2IWڒ-�!�)o��L��@Υ�y��<T`J:�,ІoI ��ú��ē>����s���b����@@B)$t�Pg�˜�!��;1��q5 ֓p:.X�#)�~�1O�Y���'��'�F���ܼ�h�A�XG���
�'{���r!�N� ��#�I�jQ��OX@(�JU��t�Q*��D
���J��ȓO?���ՠ�0%R�g��4G����S�? ���S��rX�U�J8V��M*v"O���4�O3(�x���<��V"O���I��$�L������%��Jb"O�Do�7P�#��8�YJ"O� Q	�6U�T��.�V\J�"O��p�I�NR� j�k̶}�Zqs'"O	��읈��=���C�q�v���"O��3F��3�~1a���g?�U��"O��T+	NO�p�E�O(U`y�V"OrqS3@�1Pv(%@J4`� ��"ORР��F�n�4��.�'_�)5"O�M�!��:QX`չ-�+KxР3�"O����W�K��Yi�=i��t��"O��(èTe+F@AHǤFTS"Od�*�I�t�x4��%�+4�M�"O,��2�� .�R\1�k�:ؽ�e"O�a�Íۦy��� �� ���C��'��O"�ɶ�� }�����%ƒ�P"OV�f���g�U�%�O`����u���)�Q������G�D6��aY�wA!�ă2��YcfA�b�0�!"�\�y;!�$�;� �ЍدS���Bu�؆Q�!�X�9�d����%�Ne���K	1�!�d��T�TA����z�$���/�-�!�� �]��B%�� ���P�#<J�!�]9!,hIu�{�$8�,�%-�!�ď�BF=P�.p�j'K�!0:!�ݻ$P
<p�
�-[4:	"�iݏG5!�dɞy����o[� �����/hO!�$̫T"�X֩ם���ǈY�fG!�Ė)��I�C' �hmRF�Q�!��9���$�`��G��r�!�I�"v�!@$͖;�`�Ņ��+c!�^-uΨ�cf��<} �c�EJfE!�� ���Ǎ�����.ԯ�!�DX��<�)cEѩ8w�����L�G%!�dy��xy2�C<^hY�PGV2s!�D�i���H�ˉ=?2�%ǈ�! !��
�h!��囕%?n�rd���!�ؐK{%��OK(�"|�Ѓ��:O!�Ĝ'l�����Cşoq��3AO!���wj�����ϗ}K�����!�\��v���&��tPN��C�!���X�F��V��$5�T2���!�!���W<*��p�4@%�p�U�F�!��ϸdV��&oE03���Hp�^%�!�D	t��aj7m	(������!�DٖS���Ȋ�|���V�_�ko!�$��h`��s1#�7q.5�a �,l!��\}���J8����M�!��5[��z�1{�:��0ԁ�!�d�1�h��Y
"i���λd!�<	����̌u�1C� �%�!��	�U ��H[Z����U��R�!�D�!�@6I��؀�� ��yH!��ǑI���F�П:t<ŋ'N�-*!�d޸���V��i����_�W!�C�@��XCd�*f�à���`�!��#5����J
Z/����)�ZE!��v� �s	[�|$*����T� T!�ČxY��)�1f�3 ��7!򤃝r�"�0ȃ&�D�����E�!�ٽ&�Va�D,��P�vP���)!�J	l><�#�0�X|��/q!�� �	��\[|L˧�\�hb
��"O��Y�bȤ��R( Q �!�"OR-���N<\���[)A[�At"O�=�m]�V&~h�J3H,H4"O�(BV [�lj��/A�l��'���?y��?1��?���?)���?���?�`��	..ȃ*�?h�
�I���0�?����?Y��?����?���?��?IS�oj��h�ϟ"��|���
�?1��?���?����?���?���?A4���@aX�!ޜ��p��`��?����?1���?����?Q���?����?�áW"0P{�EαY4p�Jun�>�?���?y��?�'�?���?���?�a�^�0b4��c�+y�� ��A �?���?I��?����?���?����?��G�4�lq��2"C������?9���?���?���?���?Y��?�b��=h��u(�-Ū!%
�$�?���?���?)���?���?����?�0�U>�̜@�DҘ=�7E� �?���?���?y��?����?���?i��z���$A�n���I�?Q���?9��?����?a��?���?!�bT;.r��*b�ъ̶�(C�$�?��?��?y��?����?y��?i��^5f��퉰B�� ���?����?����?q��?!���?q���?���RXl �@����N�w�T��?y���?!���?1��?��@��f�' � ��x��A�"F}����&A��ʓ�?+O1��	�M˲�¿vMإ���Mf�U	3gP�\����'��6,�i>�I��4:5�|j�� Fj��]���Y$�G��I�#Pl�nZ~~�0������	V�K�xK���"ID�Y�C^)'1OF�d�<����A	*�f�л *F؋ѹ�;���ĦՋ��$�C�����wcZ@��%� 1�(���#~E��?��'S�)��{��]o�<I'�@1Z��,�jեu��YS.S�<��'�T�$���hO�	�OD��H�I���h�N�dY�9O&���e	��K\Ę'���)1�2+��TR���IP^�@��o}2�'��2O|�#�0=ڃ��($�A����=�Y�'\rRCW*�ˏ�t&ܟ��w�';������RR���*;��Z�S�L�'���9OV�s� �,Ү8�ABR/Y��M��:O�Umڭn^J�S��4���/0�evf�+u���Z7.̽���OF�$�O�
4~����D���\���K�^Q\��N�7nF�9#������4�V���O��d�O����fK0EiG�V5��,f�-x�l�v3�&O�[��'�r��4�'6�	���K�q�ee�[�8�ڴ�>Y�����O�v!KW�ϓ:���W��3F�1b��H��(��\�Qv�� 7�Da�Jy�bB�C�����B� ,��qdF�?7��'N�'Y�O��I�M�����?�d�K��x��n��e$ܡi� ��?�$�i��O8�'+�Z�0��	�b�"�����#B&�X˰
�nH�m�o~r-C'x�(��ӱ,1��)��z��q�7L$s| H����F���'�"�'bb�'��_>5ñ@n>iE���C�� �t�كi/�y���J[y2�'U�7�/RU�D�O���*�Đ#�:;�D�-��}�P��!vY�d�\�@���OB���O ��ix�&����r$!�,�t�K����1���ÄR�n�|�²�O,�ON��|����?a�x�D��^2��%�&/��,#��?q-On�
�H�I����W��?��ݣ��"h��s�`L���k}��'Z�O��g0)��q���r"55;\z6C91�vIOTHy�O��d�	=Qh�'
�@�O�!G\R9�D��M�� S��'���'���O!剔�M���81[�W�Ι��1"DݽL�΅3��yb�iN�O��'�BC ���D�Բ �$Z"̈�ltR�'�|`C��i��i�e���?Z�X��F ��d<�2FĔoNX�s�v�L�'R�'�R�'B�'��S�0`�ђ���WS�+f�͋_l����42� ��,OF�d6�)�OD�nz޹b�O
*hTv����K�!��<9�
�˟���H�)����m��<��J�T�����	�;�X%�v���<I�Ga����f�	qy��'l" ��U�����˂5��L�vmT�V&�'�B�'��I:�M#�i_��?����T�z7�x�@`� s��+��'�$ꓺ?y���ch)
@�:8᱊I�;�`�'��p"�Mj�,้���M͟ȹ��'�ڥ�\2t���y�HLwR��H0�'[��'�2Q��'�?)�Ӽ�SMɡH��aZ$��s�T�j���?y��i�.��C�'$��zӒ�d�<y�ӼKW&��)hÃ]�*40a�D��<����?��u�J��޴�y��'\h�`2�Ir�Rz�����ј]����ET�����4�����O��$�O��d�W�^|��n�Kjz�NM�|[TʓUQ���� �'#"�Ot�����'%�-�r�m����Ȝ��GØ% 
���?A����|��?�A�1_r3��!s�`t�0�M�z�d��4&�I�Q.��d�OޒO�˓z_l$��Q|�yH��(U�4���?���?i��|:-OdlZ�nW��	�.�n�9 oKo\�����C�����M����>��?1��zU�}@��͎)G�$(��I�h���k��ͅ�M��O�9zbN�*��d��� ^m�r�����E����d=OH���O��$�O���O��?i�〉�<���a &H�W�"�9i�wy�'�27m՞h��in�|lZn�44�����K�y(D�T�[�T�A'��Iȟ�1>��dnZc~Zw倔��%��6���;�����ڭLYh�c�Ily��'�r�'�bM�8�� e�L�!h���	L�^�r�'W��1�M�U�� ���O:˧ ^�M��Kޡ�ѸĀM6�$)�':���?	����S����oܬ� ���l���`?�� ��Is:Ը�O�i"�?�q�;�dȬ+��X�M�?Zh[��/J� ��$�O���O����<�P�iۚa��� *���s��Ha�|�3��,���'6�6,����d�O4e��M�3�P#♐pU�y&F�O����HQ�7M??aS�Ă>���Py�ǉ-EeP��f/�9pl�r��À�y2V����ퟄ�Iן���ӟ\�O�m!�(N��Ȫ��Y��&͸Q�|�8��" �OX�d�O�\�D���EQ�DU��l	ug_+g����I���'�b>��`�妩�Ks~�c�.!?�h��2�R�J���̓6��S�O8��L>�+O�	�OX�K�K$�"�1���je�O8�$�O��D�<!f�i1̙$�'�r�'�ֵS�l�G���8���._�XS1���O}��'xr�|B�S�o��(�n�)2��`P�I����ݴId��m�0%&1���֦1Q�'t���QB'R�.��V<6��9@S�'r�'8��'P�>��� 7����'��<hr^� 7��sXX$�ə�M�F���?���}�f�4�uУH��u4�ǤQ7d�'2O ���<��
�MC�O~L�t���u�	&Jo��� 3d\9�خN�@�|T���ן��ԟ���ş��4K��b�ɒN��l�T�O�dy��m�<�k���O,��Oƒ�.��ըvoPr I��	���*r
D��'���'�ɧ�O�Ա��C�#>���2ԁ0�*.+.əg@M���$&}\zX���G�H�O~�zoHR�H�6<-"}���z�-���?q��?��|B.O(l�,u���ɛ��Q8��L��X"�M�X6����Mk���>����Ę-@��a�4w�D�����H���g�~�<.HcFk⟺@XM~�;}[�l����$W���#r"��sS�9��?����?����?1����Oޔ����/y�h���Fvx��F�'�R�'t�6��+b�"�:��v�|2 ��N~���:/O^�x+Dg�'/���$B@-*a���� ��JP�%V��<~�\ȃLK�5c�ɣD�Ot�O�˓�?��?	�=���� �Ϙ'���ux��N��?Y����bѩ������'RT>����X�|L[�'?uzM���3?�]������'��;�& ���1�0��	���� E��lS�l�h~�O����I�Q�'&ͩ��(���zg�>h}��
�'TJ7	<wd��3-�,�6�Q�Ą@r��s���O�ꦹ�?��[���	�9���`��_�k<���<x- @��ϟ�C�Nɦ��ug�_�j�t�ny҇V�<N��a1j�����w�O�y�T�������	ן��	��O�&%`D�E=WI��W���m0@�z��t����J�O���O��?������C���x Өb!��c2��$���Iߟ�&�b>E��ɦ�̓6�XI��Ҳ mHlD����D-����O���N>�(O���O��T摤��Ĳ㪎bh���A��O(�d�O����<aF�iOҔx��'Qr�'t遢��v��	H�av��t["���Y}��'��|A�K�ؙ�B�9yc*�!4�V����d�6�ȗ�hӦb>Iء�O ���!�
){��P�xފ��B�ݏV����O����OR��(�� �I;U�n�P/K&�%�[U�l1b� �O&�lZ"T��}��� �	f�i>�@��c��TŖ%�+�"g.�I��@�	�HaSQʦ���?$
Q�B1����[��-!!g��n�k!m�/5ax��M>A)O�)�O.���O@�d�O@�i'�>���S�2]VRi���<ᰱi��Y�¦\�#��'G���Oir�'-��$ ��f| ��f��-n���9�U����埄&�����	N��e���O8dӼ]y�Z �x��� Φ��
�X<����'��'V��;O0�b�L�	s�fz�O�V� ���꟨������R��󟐗'��7��/{���74B���E���p�W��$�$B����vy�O�V��?����?��k�cr\A�ǆ�c�����J���۴�y��'o\���Y�/O�����ez�$���A��&%��	u0O����O����O�D�O�?�`6'TswJqh �үx���0��͟��	ğ�;�4M:�0�O<6�<�DX)EQ��R7N˪Vv|� Z0$M��O���O�ۢt�$6-;?VJ[�aᬰ����+���E�  ���n�O�xH>�.O�	�O���Of嚵�ژMo"A���oW&��O��Ļ<YB�ipH�S��'�"�'�S�]�$ls�cK?|R`!Ƹ."|@�O��'�R�'�ɧ�i����1'�@�
����m$`���rȋ�:#�� C�<�'$��������}�`	��n�$#'Pb'�
���I���?���?���|*�Xخ��-OD�n�:-�$xխ�2���˚�L3�H�eMßt�	2�M�N>��YU���P����L`��T��<~%<PrC���`�I�a��nZ�<���e�`���	�@x�*O� �48@a�D�(��c� �X�4O$��?A���?���?	���i�Y���#�*ӛ@hs��ܞ"���m�>jRm�	̟��	n�S̟�C���#0�ӕm��S��*��2��Z�?����S�',�dTk�4�y�k}��AP���, 9�Dr�H���y	e_����&��']�i>u�I.n ^A*�K4Xψ<����V�����T�I˟4�'�f7-@ER�d�O���̈́N���ʠ��7H?�9AB��68~��D@�OJ��,��5v���z"�W:��kc'e�d�t,�5�!	
;hʴu�L~���O�u���,5�Aq��>.L����M�r���?1���?	���h��8
4����L�����j�o�IB����򦉀C�ҟ �I��M���w>U�塒i ��$��o��1J�'��'����f��+�c���_��x�� 놪[ ��pE��yj�d�sO���O����O��I�O6�D�O�����/��3F �f��B"�˓�~I���d�O�Lnz>�	㟀�t�0%(���IE�\d
�� ��2x�%�	⟴�Iߟp��P��'Ir䟤5 �z3��%Ґċ`"TC^P���)���D������V���O�ʓZ)B(��K�f�>E���.��`��	1�M�S�K6�?Q�HV!U�������G��T�գR.�?Y��i�OLi�'�y�ӹw�xp9���p��"�L�d|����i���,3����4ޟj����.��*d[���]���0�mǘe���O~�D�O@���O�d1�S� �h� �)�̝�fZ$�<��	柨��.�M�����|���U9���|�O˼�̌3�휒��
� ݒB��'m����c�l�������2� �$�pqP�	~$i�Av�QC��OڒO���?����?���N�|L�bO��xZq�G��?��%;��?�)OРo�-m$ĕ'�S>���&\�;nu�e�'Sܘ)�'*?�Z�(�I��&��h�.0;�N]��T衠�Z� s���,3IZ!s۴��4� q�'�'�����m�4+�t`�L,����a�'�b�'�����O��I��Ms$-A����S*/f�o!�0��?1�i��OVt�'>�(Q*.��Xp��M)D�m��Ƕm�I88M oZ~��7 ڀ��7)�	�^�2h1#�ԃ<д���㉕x�@��Wy�'i�'`��'ObW>mq���5:f�8���Y��LS�� �M�wF	��?!���?����-s���V�ኔ	A��T
�P傄�����O�O1��)@�nӆ�I��^ kD �!����A#�X���I�FD"y�O��O���?���d�a� *Z�&2��'�Έ���?����?(O��oZ7\�d�'i���8"�����o�)�v�cn��"�O�!�'&���\����0.�����Dt���-V\4�Sf���2 &?��'�2���?Z��a�Pf�Q��L�$b���Iҟ�	�����Y�OP"�	�-���RNY�a��@�����r�b�O$V�'	�kӎ�杈al]x��ܙ~�l����0����՟��	�+$"�ݦe�'��`v�b��ȋe�>Ę�>�\q�G������4����O���O���R!),���,
=H>�c�!׺I�H˓V�8��'��O5�s���C��m���|=L���`���d�O��������	�,P��_�H|�P�+�6 ���X��^��'���p ���z1�|"P�����h��@2��<i��b3�Iڟ�	��(�	�I\b}�	Sy"�i���y�D�O4-)�֖X�&�5���?��I���O�im�e�i>�ڪO�$�O0�tw�ǉ�t(Jp��1ZY�!���fT�7m{�\�I,d9�� ՟����������F	!çN	g�^|��?����?���?a���O�``g�שG�P�7N�'��s��'5R�'�x7�Ǖlo���O��n����'��*6	ͬiB<�R�M��������|��'w��''���ie��O��W�3,,1G#R5�"��[;A"���'��'��I��������	�x)�� ŊB<30����N*k :��Iǟ��'��7M���0��OP��|�g�ڗu�b�x �'Z�R��$X`~"`�>���?IO>�O�$����#d.��d�3{(�)CIB-�~�ҳi���|2�c��8%�DH��D�������ۥD�ԟ@��ݟ,���b>m�'I~6m�hq�49v/�=wn��TK_�-��!�g�O���ڦ��?)�W�,�I(�RGo�&0302�Z�J�M����ܫ��צ�͓�?)�N� Hbl�����5/��؈4j���zE�G����d�<����?Q��?i���?�+�>|SU�� ��`�c̘�^��z��H��W�sr����h$?����M�;0F�-bS ��eg:����0G���?IN>�|�G��'�Mc�'JR��dюn;^��Ğ_�؁��'A���UI?9O>y)O����O,�C�E@/QͱL�CH����.�O(�D�O���<a��ibJ�TW����}���WJ4�����@L,<,�e�?�V���Iʟ�%�$�� ��H%	ׁ8W6�XE�#?���x��C�4ؘO=���?a���~��As��- (`�y@Ҿ�?I���?���?�����O���4���r�XT�gВe�O�nZ����	��(��4���y���(k�ᣢ�z�"	2h��y��'J��'4|���i��ɳH��T��џ� �`�Dh^�`�� Z�2W�A��"��<����?���?A��?�#Ɲ=|�¹d˾N{<�XR-���D�ݦ5
bDDҟX�	���%?]�ɍ�����i�=
���_W���O��D�O��O1�.j@C�3����T�[_p8c%j��guXM�����p�OԐ?�b��V��QyR#Q���²B�0�"5-	�g`�Ւ��?	���?Y��|R+O���	�D�l��S�r�rP�����2 ڷ���
�>���ᦕ�?�AY�d�	͟\�I�OX��F���u�©
 �A�c�T�cB�馭�'���Se��V�O�'	�p�����ϟ�F䙺f�	��y��'��'=R�'����I�!����%�(*�KX'1���D�O���J즉r��q>a�ɞ�M�J>�!�A�
w`�{ťхj�2�+ˢ�䓪?1��|���ة�M��Ol{��ߪL���j�l�/�aB$��&�ҩ��'�'���ğ(��ݟH��,��P ��xx�Ӵ�VL9(���ʟ��'%\7M�*+Xt�$�O���|b5O1B�J-���j[�@SB��<1�d����0�?ͧ�?Q�k�
f �JB�ʽ2ТG�7V�Z2� Ħ`9+OZ��I��?-m.�'��	���0|��#(�	W nh���'���'���O�剻�M���1c���#�)��͚��ıI�X�	��?��i��O"H�'r�4A����k��a�^�P��HY���'9,)�d�i��&l
z�RV���9!�D@��ԝw,l:��*|��$�<����?��?��?�/���ȃ�I�ZF�y�,O�����	�ş����O.�d�Oʓ�,�	Ϧ�ݨu�
� `��2�Qc�e�B���I��&�b>��dO�̦�̓]NyP���B�sL�.�>��5\�� D�O���K>�(O��d�O��R�o��,ZX�"�#��E;���OF�D�O��d�<�G�irt!�SU���ɤq��@��OĄv�%i�Q$_SVQ�?��Z�@���,%���-:����S ՝Cahq���5?�ŧH*;s�Q�ٴ ��Of䈣T�'���EA�( ���E$So���b�
�z{�y���'"�'O���)�Oޥ����O�L����(t�6�3�'گd> z���O�PnګU�H����@�	S����]�Rr8]�m�
�|=�E,zո��������ΟlCg����?1� 
_��qϻR�$� )p�*���a2�#M>1(O��O��d�O���O1сU��+ ���H�$��<��'.�����?)���'�?闇�5.ī H�"<j
��Q%xj�I����n�)�Ӡ}
�����_U�y!į�'y�̽
��Xf�D�'��}3�kL󟰉��|�[��Q��2E4�i���3v֤�#�ҟ��ȟ��Iܟ�By�J{Ӣ�B��O�pԉq2Z��cҩ������O�LmZH�8@��ğ�I��,�IQ�b��E��ҩÃ�\$ ��YmZk~�"s_�a�Sfܧ��C�k��Q���BJ�o0X�j�<���?q���?����?Ɏ�t��?H*��Dўb*5��F�_4�џ��4_����'�?��i:�'@,Uz#ɋ�������*J��Ab��|�'g�O˄,�0�iu�IK��P�0e�%$M�K��b1@�H���P��8�d�<ͧ�?���?�!��-��J��S'��I'�2]�!y����$ᦉ�7ڟ��П�����=��� ��u��N_�e"x�8�	#��$�O^��!�4���F_�y� 	�!�9������d��4�	l�/���6�8�'��'ЈD�c�A�B� �\,�M�0�R��'h��'$���P� �۴U�F��tG0y�<R��ʫ]{e��h
�?	��e9�&�ĘJ}2�'	@49R I2"O�j���P������'�� D��搟@���p��d�~�F�=}-�|����hҴ-��<�/Oz���O��D�OT��O˧c%pt�4cE?#P>����q+���4�i�@�7�'<��'��O>�g��Ƌk� Ya�8�H���� /����OJ�O1��T��r�P�	�%���r��Xe���L�W���/7(��(�O2�Or��?Y��UՂdb��5��`�6�X�^9���?9��?�/O�Al�.D���'�r�:��@N<V5�1y��٪��Ox�'��'=�'�8`�*�^���cŜs ��h�O��?��52���O��%���eRD (�g�� 06��j�/%MR�'
r�'��ԟ\�rDӔT�bW�<�.B�m���0��4.kЄ����?�F�i�O�n�B�ڕ��HI0*��١�M�5���OT�$�O(TZ�gӒ�tv@h����#q딽"�45���þ
ڮ�S��I�����4�����O�D�Op�W�_�+��N�g���x�d��dZ����4/������?I���'�?i�.��R��ĳ�����͜ �������Iv�)��w�tSw� 3��)fO	-b���Ye�*uMn�[��s�j�O��L>A+O�pJ�(){���2��&s�օj��O���O����O�<�պi~R �D�'�i���n3z�J���^>UX�'�H7-'�ɡ��D�O���O܅�t,R4V*����q�´ctH�G��7�0?�סp 4��4�S��9B �I!9�<PIQFW0N����Ƨm���ҟ�������柜�2��%D2ظuƟ1@�ɪw���?q��?�ֹi1��r�OO�nӰ�Oޅ�W(ɎH"�:D	ѽ�� $�=��O�4��K�$l�v�ӺKU� ��J�iC�Z����膎(PҜȳ��,�?�'�$�<���?!��?I�g��K�(h� ZaC���H��?���$���Ss�W�����S�?!𤉙+v� ݐ�N��$)���|���I����O��$4�4���D
9gk�$���ĝG(`a�+�+��s��H�o7�~y2�OTp�����?&��5�	(���FA�r�����?i��?��S�'���Ħ��j�fd-+��`�2�>��:$��O����ꦭ�?��[� �	�kB���/Y\֝ƭD�	T�P�	���IbZŦ)�'�@�JV"�C*/O
�&�� ;9����-����t<O�ʓ�?���?����?Q����i�(
��� �eȗc���J7|�Pn�8��I�p��W��tq����df@�3�T)�*	�����D��?9���S�'$�A��4�y�"N�@������!�ő�-M��yb��q	�=����'�i>)�ɚn����"YET(�6G�
~����؟h�	�8�':�6�+^���O`��
�p7	S6{ ��c�o~�تO~��O��O�	cQƁ'c����k�q���c����ך�šaӒc>�a!�O��L/A_�A
r�K��n�0'�x�!�$�,��Q�oA�C�"�CpƎA���ĒӦM*p�Rş���M��w4bQ� 鏽`�]�UW.��k�'0�'��ɨl�������.�����]*lșEzx��4hٹ%)�q��|X�8����<���p�I����I�|X^���'`�8�GwyhӐ��#�O��$�O�?���V�F�h`	�M�ut($1u-U����O��b>�9V
P�y�m����9JP]��^����7��tyb�C{g4T��3��'c剟6[��0�U/d�$�(�͜ �$��ԟt��ğ�i>ѕ'K�7͆�9M��M&W%l)����8Ut��33��|K�V֦q�?�T�D��ϟ��	=�lهd�6�j�����ڄ��˦��'B\��/��O��іj�$�ȅ+�KJ��eĿ�y��'���'E��'�R��d��i����^( �+�*N6���OV�$Ϧ��U�i>=��M�K>�@�� S��W��#0��� g����?���|Zge[�M�O�ΠA���$h;3j��1�cSK��pp7��O�{I>Y/O\���O��D�O\�a��V�3�H�FN�bHDR��O*��<�s�iX� ��'O��',�Ӹ��ej��
���b�����Oҙ�'�2�'�ɧ�IK^5�f��.�t鰠�	K$� �d-@��7��|y�O�j������� b�-`��ևM�j|p���?i���?Y�S�'��$���s�ƪj�5�%��d)��B/]|n��''(6�+�������O����ې5���@����]"�{��O�����'fj6�1?�6d)w,�SJy��A��b�X��Cx��(A3���y�Y�L����	ៈ���8�OF�Rp�T' ��P�f��򗭘.t���S� �B�'���T�'є7=�.��4�ܡ:��*-�e��<����OL��<����(6Mf��C��j,̱v"Xf�Xӊq�ȫł�k"Ҍ�@��Yy�O�j׺�>H��/�ca6A�� �J��'p̭���'F�I��M�1��1�?���?ّ C4xr�Ѫ¨U����E��;���?�,O`���O�O~U�0 �ވl�������[74O�����q�̼Q'�Q�p����?�q��'����I�x�����Ɋ5����d��"���	̟@������`�O��\ @�i
�ISz
}�SB�`MB���%jS�<ab�i�O�n^�*��C�ά�[��l��$�O`�d�Ot���q���1��m!���?��M�fw��y��.&�P�TC�	Qy��'"�'��'Cb��3#�5�W��/�.t�b�E
AZ�I�M+5NB�?���?�������O��᠑=K$jU!�dI�G-pm�ֆ�<�������i�O ��ZST���n=�{a%��7<Dsq�J)oB��(��X0m�O�	QM>q(O�Ex���|�TS˄�g5��b�O�$�O.���O�	�<y�i�F�G�'��$3b�#1��H�C\d��Ѧ�'�Z6�8��.����O���O��0�:6�N�ِ���4�p�U�k`6m#?1�E^�J38��[������"f2p)֍3RMس[s�AȓN{�$����IΟt�	xy��Ԯ]�������	k,�eۗj��ܟ� �4j( P�'�?�C�i3�'��\�c�̮7_]�"iƫM�PU�yZ�M;)O�1�{���KEB�)�&W�X#2�H��^��H�ퟪix��S�䓗�$�O~���O*�0#�Ш�ÍtQ>���&ڱ_A �D�O�ʓD�"F�hV��']>�	cV�7D����'��q�T@�:?��Z���Ia�S�D�Βr�&tp�"�!G�´#K'`5��)g	��b
q]��S'2r(�g�I(��h�w��b�"�C�[�z�����	ߟ0�)�Yy��g�4-�A��m�����J�'L�-QAM�@���O�0n�s�+���ğPȱO[)9<��@��\О��#�ퟄ���q�ڡox~2J@O?0���v��9� �6gғ������#���<i��?���?���?a.�N�[ԨX�=��8Rd#��\u�'��s6�џ���蟴$?���(�Mϻd��*4�hʀ�xf��+��UI���?�N>�|�� >�Mӟ�� l�Tb^0r���AK��8��=O�u�!�
?�?�@�!���<�'�?�����nJ���T�!	l�&��?9��?�����ߦ�Xď�֟P�I�X[��F��,�@&�8N*f�����u�=��	��y�'%�Q��GK��Vn���7"6�����1,΅�|B�E�Oڅ��l(N�KB�����	2f�#qi h�ȓ6ƺ@!���%I^0�B�P%����{���@��&�:O�7�?�i���4���\��h��I�,P�V
g�8�I�����o�0�m�P~ZwT �&�O�؁)׍�4#w� �`�ǔ���*QJ�ITy��'���'D��'=�Ζ�WQ��r�H��8��'8���?�M�p��1�?I��?	M~Z��x��!Ve����,��!P���Il�S�'{y�}��	�'KR"9YI��r�Lҡ!؜d��'�wy�?I��t�	���'��I�~����P~�؁�!�����Mæ1�b�Jɟ� ��6(2�Ų4��v��1$��<�4��'֠꓍?���?�g�Z�_h����O;Fڐ���)T��XKٴ��dK����'.�t������;aI���Eҁn�ޔk�c$&���.�O��`��db
��6��4��x��O:��O�ho����',�F�|�K9B**Yb2́+"�QX�O�6-�'i������Z������/B,J�;D�[��q�b ��Oq��T��\q��|�S����Ɵ �	ɟ���+��dֈ�@�7�&��`��ʟ8��_ybd�fX��O��$�O��'�L\AG!H+i�b���фd" �'�v들?����S�����{�x#��ȼ7�f}1#���Y�0�7�R�a����K����O��(<Ov����v��u��
 Zh����O����O����O��,	:����<ǵi�,�7G�@~ȁH�1$��2�yp��'Q��'P�i>��'ңޛ���a���B�*;r�'0>m�&�i���O�!R�X���s�ܘ�ҾE�VR�XcR�aN	�y�_������(����T��ߟl�OZ�iI��0x=$�еȕ�t�*#�y�P�b�O����O������]��$h��g�]���-�5IA�T��H�����%�b>�c���ʦ��b~��F�ҹ]�
�Ca.K�@d�̓h䮝S)�� '���'�b�'O�i��1�*��oG5?����'s��'��R���ܴn��J��?��W�\��$�S�6�iP�p���:��N�>���?yO>q���E�=����=\�4�eA~rOͅ17>i��iRL��Bx��'o$G�X�km%-S�1��&{b�'���'����П�3��S�_���B�E_��y�(���Hܴ�&����?�W�i5�O�� )rG�C� dIʣ�Ư~5��ϓ�?�-OJ4K�Lq���<���w���q�h�8r����"��T�5�Y��䓫���On���O����O0�d�2#̽PP M
�V@�WA�z���6��4
_��'�����'[��h��ĭ`20E`��Y�c(Q�f��>���?	K>�|�f�{.&�S��H?4w��� Κ�I��۴$��p�b��O�O�77��:uJHH���[�H@�d��4x��?���?y��|:,O��n�<+��;G��QaVc�K�&�B/i�������M��>������j��a�8i($���	W^9��Og���$0�e�h9N~��;E\.��sa&3rqҕmS4S�p��?)���?)���?�����O�$r%��g�x��,]�d=�9�c�'s��'��7�
�1~��a�6�|b��4���ʒAV�}�JMpԨ�+;^�'������M���F��\!C&MNs����3����㍐O����t�'0�5'�蔧���'k��'M�ܨt˞�e&�c�_����B�'�"R��s�4(��P"���?i���i�dL��,,j	<��w�ܬ.E�	�����O�� ��?�S�S0b,��,�r'칲D�H90;:�B���ۦ����Z0A���d�A�ȕ����x4�鱦d Y���҄jD�ɨ�`� _���@��Y=�e��4���0cTVC���g'��Dj�i�Q�*q��3��3�r3g��+���D�,YE�D�5�ݳo�0�"���P��2@��}"�힤�<L@���?� �����,t��z1H�J���э�$l�0�D蓾��k�3?Q��N�<Q(y��/[��&���'�icL9�Q�0���p� �e
LqvG��7	���е+���ҁO�Z���t,èP%>�rĀ(s$`xP&��'JcR���'~��|��'��Z�i�dh���Q!�-��ሪ/$�\x�y��'��'��	�DR�0ӛO.�vG^�=j�:&�	�4у�4����O&�O����O2��쾟��O-A0�,Z���*8���c�>���?)����9��p�O>�O��Q�tX�M�b�T�b�Q;�6M�OP�Ot�de�@c�d�@���j���@�z��D�r�&�'�X���5P����Oz�$��B���ME�řG�':rB��FLt��⟀�	kG���?	�O��Q��_2��)B�OnVJ��޴��D�9<�}o����	���S
����d�K�F�~�<*��ɆPЄlqD�i(�'�,�K2��8�S�i��X
�ւ;8�8�K�,Jh��"�.Kt�6-�OF���O���W[}bR���'�3F��`����0��
��M�֍��'��@���g���$��8�\<��iT[[,�n�����˟��d������<Q���~
� P8[��.6�>�Q���8�SD�i
�'�9ڷ�|��'����5v)�! ���z��"~Š|GI��M3�zal� �_�4�'u2�|Zc۔��E�&��ؗ��b��� �Ov���'���OZ��O�ʓWq,i�P��0mbY���]F��<)�Ǎ6h��I|yB�'��'�R�'k���P��-L��pqL�Qy:�!G�8p�'I"�'i�Y�Ě2�����J�m"�l�W�[rV"�X�Y8�M�-O���!�D�O���O� ����۶m8��s֖x1�K�A�b�"��'���'Y���� ��'O�~�B���$
؈;5+؏�*pI��i�r�|�T��S⟨������X�@�8+!��p�8m�i���'$�I�\��p@K|
�����LzF��g�J�h_��
��˟-��1%�d�'���'��yZwސ��F	f�^���IV11$�Bڴ��D�52�$�m�!����OT�I�X~b�I^�AӅ.������ҟ@�'!��'g�O!�R?q�iӕhș8���q^�����O$�r�Dɦ����T���?13I<�'MW^�	���ػ�����9Ӻi�2�'���|ʟ�ɮHC�h�e�ëW�R�j�"�
 �)�4�?���?�J���?�O�!{� h�b4z�!T�{k<t��M�'�Fc?=��s?�TN4z��!Gk@�g��5��ᦥ�ɧw�j	�'�'��'q��c֓7q&��g����)%`.�$�&H�1Ob�$�<�:���#�ʎK�>�s1(ʅg@|�Cռ���O��$&������e(����FEc���F�B��mZ�,�$c���eyr�'x!ߟ�v�ݶj��V'
)*�Jѳi���'��O���<�&������Iع$�jx�lK�RBD94&�$�O���?��k���)�O2	��(
�}�~���| 0ֈ[�A�?�����d�k�'��Qä2!ł���B�0���4�?����d��<�xl&>����?��HS�����e5v\J%�.+�J7M�<���?����?!H~���� ߷0�`���H�E�`�g!��'Ox�9$|��Osr�O
��it���Θ�:�qEH���n�����ǟ�I�����<Y+��v��:d���XV��d�� ��M��D�R��&�'X"�'��D3�4��؀��Ozk�蓍�q���OW�6��O����O��O�3?��ǂ�����X%�xJ�j�tÛ��'���'!H��^��'��*p���@g?
\�1�G9?{pU�����Q�ϟ��I�����i��+�09��jX�Px��	 �M[���k%�x�OF�|Zw�5�d)�8KX�#� L *.6�BJ<I�����O(��OVʓReb9�U���A|��zc�I�VO ��aݣ&�	Yy��'^�Iٟ���ǟ<��*�,}�^U�E1R��q M���	Uy2�'A"����́4�:��'Ւ�
׭Ӯ�.���h��7��<)����O����O�İ7?O�%�q��a��#���'�H�e����I̟t�	џp�'�$����~�����/#h�P�{�iU7k��
�Z�����NyR�'���'��x�'�r�'��Y�G�g���R� n����dӆ���O�˓B쨁Y?�������I'�@�%���M�|3� �t�Jeb�O�D�O��dG\O��|B���d��:K��LمmX�{y�Bȸ�M[/O�P�����������H�	�?�B�O�n�$�l�Ps����\���ܜT����'k��y��~���O:�<���$�F����J>[���ܴ.{� ��i�"�'�R�Oܒ��� o|����gT�PE�rm��f��o�
���Ė']����9C�:��Qf��G������A�uo��������󄭃��d�<1���~�NF.�̅X�Lɖi`A������'@)9�y"�'<�'l�8p�@]�&t��Z
oU~�S.w�����m��L�'��	ɟ��'�Zc��3 IB�N��A&��:ivH){ݴ�?av�<���?���?)�����B	|N�y�K��..;��A�1���g�X}�Y�H�	Sy��'2�'�mX���/o$��(��T��'���yr�'���''��'f�I�D9쩳�O3��k�I��H� 3�eJ�M�/O��d�<����?I��T��̓|��QE�� M`���B�ۛn�ji��[���Iߟ���uy"'S���'�?YE	�\rd@�29�4�ƇJ-L��6�'��I��d��П�çb}�D�O 1�fmƖN��Ӷ�$M~��`�i���'�剺J�ب����d�O��ə5l�J1��B\?WI8�R0_4�
X�'���'��GŇ�y�|bПR��T���d��D҆]R<���i��	*'�0���4�?���?��'�i�i�����8��y���J$n���I&fo����O��9O��d�<ɉ�4��$�28ӡM#"�$�j�-D�M��&fd���'���'M�D�>�-OX$1�D�;(|�I�	ڳA]�u7ڦ�ee�H��vy2�I�Ox�zvM�I�hy���ı^��hP�(�˦=���ɱq0�i�Oh��?Q�'�Hdk�L�X<�(s\�p�aoӾ�Ora��6O����d�I��`k�W�SvN��@���@Lkc/S��M�D=�51SW���'�RW���i�m�"�S�(��fi�� �t�xӰ��D���OL�D�O��$�O
�`��0�z_�d�CM�<FL^5�a�>t0��^y��'��ޟ4��ן$�� <$�@!�{���X%Ad��s���<����?���?9���D�.� Χzk^����֢UW���C�|�n�IyB�'�ɟ��I�����b�����p��K�Mf� ��3nF����O����O��p�C�\?��ɨp���c�Y�H��I��Ȳ.�Q"�4�?1.O����O��I:,;���O.�I ����%�P� �3r�W��r6��Ot��<a��P"[������	�?��r�/$��|���˜{� `��T�����O��$�O(ԫ�3O��O���v�J���1nG�-1c�O�/o�6-�<��!{�f�'��'��>�;]Ѧ| ��X>�JE��f���m�ԟ�I�mۺ�3��9OL�>�⡪G)S�T� F� Q ��+!�j�ޕSw�G�}�I��L���?S�}�1�>��6�ז*�����]0Z7M@(��5��3�S ��a��[+�UJ �Ү|�f�a�EH��M��?���.�*	��x��'<�OrAr ��3
�{�K��Zc^�#�i	�'D������I�O��D�O�(�.�`�! �`,}L}87�O�A[�`�B��?QK>�1?E�5 �ȗmV�x���T�e�'B��[#�'a���X�I����'�*تa���s�`"�@��o��t�� S>�.O����O���?!��?�S��r�"HP#y46�h`�.7`�#�����O���O�ʓ&.���E3�R]�V��>_ޮ��B�VL�nS���	ϟ$&���Iϟ�Yq&k�p+G!�hrvhӴ��(jqvjR����O���O���D0"���#��X9�ҿ��(Z�3z)47��O��OP���OB9�ť�O��'8�1�t�8���y 
�1':l��4�?9��򤓽4��\&>	�I�?q�l��f�z�՚}�Pr��!���?���.Rϓ�����K�-P��A%H[�u�hц���M�-O~���S���{�������h�'?��[`@�Pd��h�F"^�x�
�4�?���!�VMX���䓟�OD~�i�(ڸ�j3�P�޽	ݴw|�A� �i���'nr�O�"b��ib�V;E~��%�q��i-�M�R��<�I>a��4�'�T���>��j�AoZ"	Ȳ�s���d�O:�D(/XF}�>��~���P���W��YB�5����M�O>������Os��'r/Ԕnl��0Dm�1Y�j�-W�0D�A�io�B��YJlO����O��Okl��7b��2�jT$kC����f��m��']�]'�d�	��IMyr�M��Ո#ꗢB/64 �ǌkn��<���O��=�'A� 1D��}�u!0$�4�0u�ش�?�.O����O��d�<y$�W��i*@>�K%�C��T�Rs唰qu�	�E{rT���ɮg�%8Tąz�$D�%@̯'gֽ��OB�D�O��ĭ<y��݄\��O����`)z�i��ҧG��I�r�x�=�)O��d<}"OY����v���?>(ᒆ�M��M���?1���?A%c�"�?Q���?����!�I Q�� C��O&p���H���ls�'��^�t���'�ӺKD
$w�Hmc&��$oɔ�
��Ŕ'��B�	w�\�O���Ogv�c}�MQACߵ/^�`��.D$�@07��}��&�p)��I!un��ٗh�;G
l�a��j�z�#�N�OV���O�������D�O�'^O05ɷpų4[�uD<�z}"�A�O1�����h~�U86�֝XM�Q0�*��l�&}o����	��D��	]`yr[>��Id?���:8ٔA���Z�vU�Ur���	c���N|R��?1��J��p�n�%J�\��3)�p��uX��i�B�W�S� �@*��l�Ix�DM7��2w(�/N�h�[�J�4+��'��'��'���'W��U*K^�	OC�8	�T%�g���ːU� �'���|B�'��$�Cd��b7Kıb���%	؛�g����	�*p
�!�)�4�3q�pE��D���Т�8�yBf����В��*�����T�ϸ'R��
P�1�&� �'7 �B�ԦG:$�8�����%���C��;:��aW�3��=8S/Z�6��lP�B��f}��Z@�О	�Zu����B��fX��2�y�)W�!�eaV�}ٚ�P1�H�0.y��k�Xe9�,xr}*�o�D��D�H	��9b5>�`�*c&�X�c�"cH�̀U�H?`��Q ���?��a֑lZTts�i��)�eʿ_'d�Sp��ā�/@�@Fpՠ�n���n�\�BMP)/hT��dc�1 ��t���$�H�lP�;�e+'o�,��	!Y6��O�}��wK��c@fE�6�=�E�ձ��۲��"%��A��S-ت~�rQ��I��HO`!��┐�^�y�N��q����#.r}�'i�@�tz�cq�''"�'�w�ԥ�6/juP	Z6�����G�QMrA���O����h�1��'�:�h�5�����m��3�=�l�)�4銓��O�5:��P���K�2ف�#��_��*@B�E��"���dD���O�ў,9��F���I��"�d�P��Ff2D�\A�M�7:j���� 'b,�Ȑ
4?��))O|=2J�9��$b��!.f���hC�xr���O��D�O�dº3���?Q�O �B`��g��lCv�<"���6�D�0�t	�Ɋ�T����$U���x�lJ*"���Ƌ��R�������j$J0�Md؞�j�� �u�b��c����딏h�`bc��O8�d>ړ��'+��*��\	T{
=��
���	�'��	��Ns���"���;�d��yr+�>q/O�mZ��VN}�'k`tAF�_����YS�ľ\x����'4e��5���'Z󩕬'8��[�Mȶxi�L�D�j�8���Q�ȥ2P�e�b途�'��kdM�8.ԝ��� 6i���=r��cj�@���h��҇�p<y�������nyr@"p����&"�$p��6�'��{�cͨ
Y`ݢd���Zg��xb�r������Mw�4h��_ݜ��<O˓B�4�{fX���	B��fΠg����,<>�$J�D�:ld�%8�(�Zh��'^�bՠљs���׀��0B�T>1�O%`�:4�3!�\����Y_nH�L���`Ԩ�9H�i��E���]-xx uZ����#>�� �'���ɞHG<���OR�}������y7��'P�v4��`E2w��܅�2�0`k�.�06��b�*Ǳ>�̤��4�HO�z�,ۄp+�1r(�[�x�A'Q�I����L�	�f�̛�C���p�I����i�!���I� dI��	)BG�	@*�9]
�5��*��?�"�� �$�|&�֓<9��-j�IS�K(�el<e�~I�n�9R����H9o��yR��L>�FnVv���E�U������V��'�����S�g�I��	��&�X8Z䁉�!�C�JA.�#��19L,�vi:q��ő�"|2w�-Ν��NUG<=�VΘ7;��]���?���?1��,���O���q>����9J�> �Ŭ�Z���ۓl݋h�BB�	�}�28�P�D@$�cE�A������/�$�P��=_��l�U/F�������ǫ0�P�$*�Oĝh&��y�(EcK)xH\��"O@iqSC��k��D�7Ѵ��2�$�Z؞��fŒ����X�dC�Z�z���=D���vMJS���"�� @PY+D�:D���3Μ�Vl\��ϛ(`.��,:D��:5�8~6�)`��=(��!sB6D�d�P�8��\�t�U&~i�H�5�2D�ds]/ܼ��+S}	��rWi/D�t{E�T8:����A�[v9z�K-D�XC��R^}��T*_�&<�g=D�0w͊F�����#v�u#:D�4��BF"qjtzs��,3�p��,D��D��A�����+ U�a�vM(D�X�'��MzP4BT�	�aɥH,D����!��{�@��b�>~�D��/*D�taD�M ;8�P�D��i�0]��.+D����M�sf`�-0/"]��-D��8�oV5A��%�Ǎ�7DV��4�/D��YT˅1�<�	@�̂42l|��H8D�R5���brr���9�9��7D�H!�֊$�V��+�
�r��p4D��b#�Q�#�3��Д#� yҧ=D�`S4�@�qXM	�̏�	� {�	!D����'�o�RT�LX��иm D��hV�t��pC��F4�Lq�$D�d�ċڡ6�Y��'D+G,~,��-D����� + ���!aN
5�VT8�*D��;��
�I��e���%S
h�#�;D��D;{���AȔNʼ�y�'4D�$���^;/#��@n����qi2D����f��7�^�c�kO/�DT�k*D���d�ѠF��e�U�MYR����(D���4�E߬U ���.)��0�"D���V)Z�5Z@ �u��H8`6=D�t��!ߡtR��ض�E�]�:qz�:D����ЌP�2��VD�>(�p��!�6D����6�8�y%mX�D��`4D���3��%��Л�a�y���ק6D�`����1|�L�bQV�ECA(/D����IӘ��aC��7o,�c�.D�� �<���YIKx��!��4�,�p"O�D#ń�;�<*�G�!/1��"O���C�2��gE� �3"Of����W�q���Q�>Y;�"O֝��'�D>4��w����p"O�qEh��i� ���N�l���"OB������`-ї���PI����"OR4a�,�,|���c�aL.Z/����"O
�;T�N�w�2���= x�p"O��恍*_N�)oϲ"J�"Of�[�%\r�,�!��B>I-##"O��6dʤ8TD�����h�\�*B"OT�IV�O><�]a���'�*M��"OЀᄆJ�g%V-����<?� ]�"O�9S �@�8R��޼+�� �a"O001��z s聖l�ι�"O�9��˂
;<�IC�g�"9����"OtM; o޺T�>0ǎ-*n �Ȥ"O��U#�$-�6�#UF�6y�Z� "Ok�+ȅJZ��1�^� ޠ��""O<U ��-O)��5ŝ�j�:���"OH�` ��N�����	��a"Od1ʍ2Z�՛gO1�*���"O0�ɠ�O4Fh�A�R��;*�`��'� �� �H���cEA }��Q�w�zB㉻���	=��b��L�/	�?��L6g,�b?��BO�R����­�u]İ��H,D�؈���Vb8�� &��dr-�<��d�k��➢|Q혍7DL���R�)���x��P�<q��PjH|��Z
�t��uE�O�I�d����'��T����$�B� �Nh�F�	�'��t�'Ɣ�I��2l�#�^q��3tj\C�I�$��S#�rt"e�W}ȣ=!�/9�'tf6Q!�F�$D����"F��ȓ[jQR���X	ë́%|Qn��u��O?�đC2S�e�}S~ي��P�q�!��J����
��ju
�m�Q���
*p	�� �i�W��\(��9!���U��ɁH`�B��O2ѩ��0Kfs�;;��|�"O�A�T���	���F���pYǐ>���<�:ⶆ�h
��1�E���OP�9{�!��SL|�+��H��'�z� �ٽJRD��焴Xk�e��- ��ܩ M�9�?��nI���O�NI�O(��T�����HM�ٚ�O(�ͲPĞ�i4K�]�6�S���c_�I��Y�3D��!b%(�2
�D�Pt؄�O3��-��)
H�e���l���� gP�X�HPBv$��:�9�GL)?1��	�0��m�ʸ���Z�Ԭ�d(�,���,m�DݺA����T�ؐ	���J.Nc�)��/V�V\�Q�����A��2��B�ɽr��d@�	��G��LJE��/E��)�_&���%��Y�O�	x��ބ��qp�1�� ����Y�U�l}��	�+���"���\���C��]�i���!	pec�Ô���8�͌�;I���GV8�Zs�������D�����HO\� ��*��y�ڈ��O�}}��ܢ%��s����5��R# ��,��$�f�S��5i��B�~b�oZ�dU��fb��fM2U
�G3!�8ӧ�����m;�� eF��^�:��$�Si}��*7b�|�"R9j`�&�%J:�%�@ě�p�  ��x≘u���6��A���4,1�$�Oh�r��>^�i;�Oc*�����'ٌ�F�6Z.\�2ч�<e��\���;���~��	!��ò<g����S�?n��g�̴� �V'F���1�X�<��Ep��$�H���kE	̍�����k �p���>?��JT ;-$J\+�%�_�L6�ډd��`a��x�ǟ�w��Fi����P�(ȴH�X�80#�x�ya�.E�M���U�C�By���g�IH�޲�ч�R�gv%�#G  4=��%�=���;�lNA����W c�R�FH��7t��ѵ-��app2��|��	��6E�4�`��{U��%� ���� ��l+�(;�O(#�nK�Y�(�� �(��W*�.{A��J�丩`���U�L2R�,�\2򊞷_��sW��C��(��Aֺ�*�M�'7���Z5(%�+�2UO�t#Qf�0�@8�'s�P�%i���;�Ø.��6��8�fJ�+�������*E ��Q�%a��Ty�=Q2�*ӛV�I�@���H�JƹC�kj�y����<8� ��r�	A̓@��ӥ�$h]-�B��Y+4�
�I
=��@��)�2q����$N-*��jG%�KUjTPR�B� ��ՠ�)+�&�ɵ
u�(�G%[ y��Pڰ�S<	��yu*��_Vޙ� �]���>1eI���6x�#�	>��`:2l\�\Z��0h 3#8�O��� >vdx������1qrh��ҀAL��`A��9ʚp���3L:���G�ȑ��I$'��c�i�6��Ѫ@��<%͸��V��Cb�����W�ڂC�L��;&�ݦ��"��p� ��	���a7�a�|�I1".-0U��x=D�f�D]Xd�qz�r�(\�/��!��e̓	CN�p��L����t�K���-�4�('�JeK��)Ǹ���F�M^�i˃��B$� � }uh�����|�h�#P�'ў�'/�� �vf����꟪&d�9-%����*�X1��㈱@d��"`�U=QB!h��Q{y��2�L���/ZȺcÂI�0����q �R��x`��:U��݄�	� �֨ r�O���Q$�:u�|b(KTڐR��_�^��	��,PkGB��|�Ū^=b�➐�P.D4!Jȸ�i��0wް��j��[TJֵ������$kH\***�P.,]�2&Ţt�!3OP������%h�R-H3�q�a{R͎�cm�2��M�X��!U�i;�.��p<!�.��@u� h���t�O*4�n��ΏZE"���W�b (Bפ��wq�� ����di���)VQ��"ՠ��3�����Q|dh���	�iz��%���أ ��q�t��℣j�T��Q��5�B�N�^�r�H}��2�^�R�~�"�_�)A�		6�/���i���
V�$�쎰 ���6�N�~� �}r@�:hW�Q+�iN���a��㏿�yr��UJ� 6H����sH���O�JV�-8'D� _ �@�n��$�����JQ&�%��ɊTYv�i��p�u���&@O �J�m��V�8��D�6�A0"t������ . y酤�
K���0�<�O8�9���Hp����=5=LSI9�nxR���%!�XP�s��u�LWY#yynyPֆ>����	��ziC&��&g���	�68qL����kZ�y�.�c��%M`~Ԩ4)!O1���w�CbH�Q� �W�
R�S�9/.�a�}�D�<�l�:D�U�©�D�Ʊ�OH�:2T���Ɍ0�8ʓ|I���f���T�T;;�P+�N�.�Fq��Ǐ��X��O�2Z�x#P�J�>Z`=���.u��(���~�'�(t�/OJ\K�O�#Y�P���5f+��v���\�:�
ly�X��y�O�4�VeI��J426��������~�\��?i�Q^���-����������6{t�K��$Z �0�%'��G �B�	=zݖ��ǅ��y�K�Y2�|����L�Ruᛱ0�U�!�ط-]���ϕ-Q�c��ӵCYXU^�B�؛U\컡�;O`T{a�& �Us�疒/zt�R��0|s`@�'s( �Ȓa_�࢕�W�����O�4~����!i�R�#�A+�$�'R>��C���5Q�虂�ߒ���~Z@��6d�����S��a�+�X�<A�aY�D�� B>R�C���8t��TJ0'�J�D�!��O�b?2�$a?Q���kZ�I�Q�*����r`H<)�)�<�6UBV�%!�Ԝ�'����eC$�Q�E�?2��T'�ĨOy�)$��Y�1%��/�<�q�'�X�5-��F��=�uC��	�ljP�ΞY����$KѢH)���HۆF����I=u�H�A���E��y�h��DR(c�x�`���(�Q����wcz|H� /^RZ�M�N�B�	�(xg��m�Dy��)-@�~`5���0�' �F�,O��b��ؑ�np`I]�@�j�"Oh���>lܕ�C��*ypr�{C0O���2��|��Y�w�C6Z��"�
�p>i�k����wKF��%�X0���<B�!��-�*݃���R&1"�cAT�!��A!]�\HtkB�a�8!����!�$Y��-"3�9Qf�E�� "O�=�ƂV=4�x���	�AȆ"O��H��be6D�f([�5I�"O���BB�we�pb.N�J��@�"O��8���2�>ABQN���s�"O����P*ZT���BL6q�~�07"O|�za�>1�:-�t#-��� �"Oj�ه�Ш������z�����"O� �9��� f `PǢvzH�X�"O�%)�c��^J4������X�0"O2�#��J^�"ј�,Y���A�"O� 6GO�th(���1j%� `�"O�E(�-5U�`HJX�9����"O�\��"[r��@�i�����-Do!�$�1Aߴ,��iϞ]<�P�&.�uH!�Ğ���R1#H�U����r�!�V/@^��.�b`��IR;#_��'�� $��Z	>�ar�_�ݫ�'Ҽ�S"�5	���E�3 ����'"�A�6�������1C����'�:la����o����!��1z��
�'���gC�c�ȩS�n�%/քp!	�'U�=���0!��x&�ͮ*DΌ�	�'Fp� O�(�lK�G��k }��'LT�g���	�%�4c�.(��'v�0xg��$s�<S���bjl�'&�aU�T�c�@�XS�PlYI�'>�Ȩ��Ӄ/0y�b΀ A���'������"+�V���+�t�P,q�'�.0Г/��L����B�q>v���'�d=*b�Yҡ؃�ăn�����'�z���
1)PDܳ�i�<a�4t�
�'z�H�%+�:GV��5�R�Te�I�
�'�J\J��T�D��u-��`�(�
�':0q�|�=�d�-
ej,��'�$99#U����[$�^�wW�L��'U,���G�3\*~�y�b˦r�8�)�'<�ua���u�t3CK�.o��h�'j����PH�1!2�\�uCJe �'1���&�,�b�ha��E=h��' �PkR@� 84��0K` @�
�'���E(�dis`m��0&耑
�'4T]p	܇^�����J�|$<E�	�'x� ¢�ϓFGVi`�n�ޘ �'���x���[�$�*�?
i��'L6��d�!'�Q�&	 '/,\��'9�!+b�H�Tx��\� �<X�'�>��W)0W����,ü)J���'�-+��$�Z��-׵\�0#	�'��%�B�>r�E� B�: ��'�F���J ��݊��OM��I�'W���v$V��^T 0�A���'Qf��.Xb�<	�7��	�����'P��s\�8bWOýS����'��x`�0���vF�9bA�� �'xfAA�Jڅ'+��y�*�$Uq�P��'�v(�VZWh�i�d�=�J��'@�8�jʺ8[z)���T� !�ų�'�2�k��5|�1 ���m��'��D�p Ŝa$�=��l�>� k�'���6�όX#��Q凙�[.��	�';ղ�F����H�l �.�	�'�\E�6H�?`^�<��X�~�D		�'�H	i�	���B��C�to��	�'��f�3������l�¬�	�'�"��F�@]�E���Rä���'V�|������Z*�PZ�,+�'2�0`�6^���cZ?E(Lei�'$�ԡǒ!/�+d@.h�v�J�'� ,A���G��� ��"e��k
�'M��qcߢ�93�cޕ`Ŏ�Z	�'����E�X�$��Eڙo�r�#��� ���(�
Ip�W�i��"OF��`� a���"�́�J��<h��'�Q�X��&`u��� Y��0�$D��"��8/�8u{�̌�N��rQk.D��j����PQt�`�o`�&QaZ�y��Z�V����7d0u��;ԢX1�ybh��N����%CD�iT!���y�HЊ.�<�#m]*�(�cc�y��RP*�O�=3Z�-���yr�?#{���A�]�:��cg� �y�+�	��٢�՗5jD
p � �yr�	-�4`AB��)��tA��y�cׅTx3oS�O�MP��Q��y�)��|�`e�ԉ/T��:�̊�yb�@�'"t�aY(����3���I�'���� cG4\@��(�6���'��y"G��
��T+@�.���'�X�H���wIH������N,
�'k$�g�֟n|
̩#���8�q	�'�p}+���*t��u�,QL$+	�'���HE�9�&a�Q F�`�'�8�r	����b�D�* ����'`��:�bN�y��h2��
"|ej���'̹�a�F�B������W�&G����'T& ��lP�t��#C�� +N!P�'����E�EPzղ1��I	Fi��'�| b�&R���{�J>DƘ9�'����s�ʋ`4E�a��>��t!�'��9��B�q�h�+
�9����'O�D)�F��y�~���F�N(��'�*�H0Lºq2$�ۓk��	�'6�f
R� ޴�Y��$U��T��'
f�+a`C�_΀U�5nV>���'��h�B֙($V�2`��A���
�'\|!��F)K�V]�����o$9�	�'1@��ѧ֧l9 �.ek��)ZK�<�"��`y�(�EL�?@f�`��F�<I��Ѻ{j4X����0iTB�<�F��9�z�1��ÛD��uxb��e�<��[�V�2�1vHJP�L���C�X�<ɶh ]6ƴD�n<�$��Q�<A"�W������ے5C�IQ�<���c����4~ ��Ԧ�u�<��͖�*���Ď:T��Ji�i�<��e��Q ���^:��(F�c�<��
��c�%H�  �ӠKf�<Q��Ȥ1w�M+c�$J�ĉ)�b�<�4FT�i����e
:-&�jF�\�<�%I^/ iƤ�Ej�`���K^�<q1��@���%綉q'*�o�<�s��.,�P��C�+~�Jh��%A�<�s�^'t��5��JF#%�s��>T��	��N�Y�t�$�A5�L�:^���	6MZ��:��V:Mu�
���fA�C�	I�X��O�'_�1B6���2��C�ɻ{�D1CG>2]�%�C4 �C�3jy�gBZL�ժ&k�ήC�I	�z��,�r��̓b��oôB�I�}x�x�a(��Q���K�*@��B�e� � ]��@+2�[�z#|B�	&=����ӅxC����Y�ӸC䉘 "N�1���F�vi��&�k�R�'�a}���M��׎�
Zӌa�ĢA�yB�~��0ڗ�N<p�@c@V�y
� ��V��t��툻fk�� "O����Bs�\z5R0b�"O����/u��qѤn+%�����8D��a ���T��6$��=p����5D�8�WN[;{22eU���Yٲhxb'D�\!Ј	Vt4��G�X�7ֵ+`�7D�0�F���P(Y�~�|����5D���AJE1H����U;%��4Y��-D�� td:��C(7xL��d�+D���t �����,�Il�cu�'D�D�Ou�� �Ps��sg�1D��*&��7-zZPjB�� VP�f�0D�L�LQ��x���!Y� Ɂ�/D�Drs�T�*l8�2��u�x (+2D�\�b�p2����F"I�,�z��$D�<�SD�1!�T�	��5>%�V�!D� H���!��% r�Ǻ��҆%=D�4� Iv�z�#a9G�Ψ�u.8D����͓�R���B^%{��ѐ�"D�� c��q}6�;6c�@��c!D�p!%�S<m���6"�@��� $D�(�.�5ush9�K̢E�$��/D��t�;q��0q�J6p��y��"D�0㳡
�}9bm{�g��(�]���?D��*v�C`dd�$[���Xd*>D���$��:�$9B�-#|�Ɓ1D�T:���>F3��럒|���g*D���0�֣`jJ��b�Yr*�YYt�-D�@�G`#� ��T���`H�8�%!D�$"c �!|�-h%-�\
p�` !D�����OI8��c�3mU��C�4D�i�噭[�PyrF�]�.�ĉذ .D���2�� r>L�T��.�� bRg1D��#BF�!�� ��m�o3�����mӼ�=E�ܴȔ���@)0�m���;| ���cvJd�s�] 5���*���ha�ȓ6�P���v�jҢEK e�ȓ �J���'��<¦�B42��ȓEu�H��ܔ9�0	@DØ2(���ˊ�!"��]7�a�)	
Q�Ѕ�
��뷮��!�L�Ō�q���Ezr�~�ި��:��$H��x ���Z�<y�"q�\��d٫?�`�����]�<aB#3���S!֭C>N��O�<�1D9|��6&�\�nU� )GF����<!�̀�l�n����m:H�3���B�<y7d+]C03�4.O�%��h�J�'ў�'��Z��Ů12V��c��5U�48��4ÞT��ˎ�x�:�.�o܆U���>�S�"\��i�J1)��ȓG&h���&���C�$��X��Tb�"O�����7[�ȋA�z����"O2��Fϓ���w/V.}��i�t"O�A�e�R��
nY%��a��"ODt�ѩ(kd�)�,�j��\�t"O��	Ƈ�R����*˿\�@,V"Ob� %$ٰu
��Si@8:���B"O����aҢ=p�$xFɞ�o*��V"OX�ɀ��:`�`5#H�9("�a�"O��rVB ;Ȫ K��M:+��pR"O�Q�,��r���/��8����"Oʈ�b��,x�B���'�D�[�"O�e;�D�s�mr��,]u�1z'"ON񩄏H�Ê��g��w�:M��"O� 
EL�'K����bE*7�R���"OD�ztDL���p��7"��	Y�"O��3��?M����� a�3 "O2���%�7\�xl�r)�@�1 �"OTE d(H�!Bܩ�רX�x����"Oڅ��0F����'A�K��j�"O� Sr9(�,u5�δ��$��"O�mHP�Z#��3�	�+Sd��B"O�L�`� ��xx�B�K @�4"O�13��>:�6�����{iށ��"O����Ѡ;�(AiM�~H���"O��`�7v�� ��"U�.���"OfI�k̙87X�P�g�N��ˤ"O��a6����z��P������"OLpAU4*+.�@L�: �0l�T"Of��eN�fT9k��~�H0� "O�\{��F�7�H���)��6R:��"O4yw!�	�H9Rq�H� 5\h('"O6��6�*I�+�"ދ/��@�'��j�l[=AꞐ��m��	�p���'��!ڷ�� W�eؐ �+W��')|0+q@ �:�p��#S���3�'c8B��Bm��-а�8���'�z9v*��5X����B`���'@b̓3JF�ؔP"
�i�����'�\�H� Ю$БJ�䘆Zú�X�']*pX��8�~��F8$뜅��'�@�ђ�
?b$B�y�"W����s�'��Pk�"ɄZ�H��	��hּ��'u��b���${%�U�)�J�'���Z7$On�B����E�%mޠ��'d~,�6K�J	� A�˴#���'�мQUOB&WY�l���J�"����
�'�X�1cH1frR�"�nCک�
�'��HT�O:c��e>`} �*�'h>t�nŬ.�>H��%�S�B�R
�'�V��o�I� ���_"Ƅ��'�X�b�I�(Bh�e���Po�F��'�v�aX	��a{�/\�Qr<�[�'s����ɇ$8�#J�O��)��'�z}�t��0ȄR%*M4I�f���'~BĻ��ی��l�6��H��'�\��u`O*�&����3��]��'��\��蚵�:��u�؉2�F5��'���S�(Hd�Hq��B(*�d0�'�� ��N4U��XǃH��%#�'s���P�F�/��\�&�E8m�'��C��FN��5W�{y�B�'J0X�G� <a�����.y���(�'~�z��? ��P�� m����
�'Ē��ACNl���oN9z�*X��'��(��S�t�����[i���'���X�_�x�v``��W{��y
�'�&��N�=���gC�zZ,�	�'q&�jE(̉4ӶM�W뉲b�J�@	�'Y�@PP�I�lGh؂fĉ�H�h8	�'�*���¼P
��o�W#`i�'����G�o�b���:y"��'��1��FC�6�:���%1Д+�'�4�� W�8�8�.�/x��'��$���6G�2�{%�D)S��#�'��C���%a���Ԋ?4�����'�T��T���wm,�[3\�|u*q�'�1�2꒗7��r�9o����� RY�B@�oL�(ruB��!�&	"OB<H�*Y,����'��?�PiP"O�x
�NP�M���Ҧ�XX�`"ON�[r�<�^D``��8�Tɀ4"O&��T'�4}����W� ���"O��'/��c9�����΢Ը�3�"Ot тi�&@gRXc�a�	��X�"O�у�Dճ2�9o�d��2"O���5�{KDkE��&>��\*�"O0$jW���S@BT�"�\�VЪR"O����< `��9,)��X9&"O���tm&�b���z<,e��"Oz�I1�E�v�D�I��M��"O����3��]1����B	ۓ"O\8��"�K<9��7����L�<�r��	=J�0�둘d��B�g�r�<!��VJ
:$�㘎e�d���x�<�hIv�D aɤw�R��@a�Z�<1��5�}`��_�������V�<ae�����P�"��K��x��Fl�<A���mƵ�pI� ���A��C�<1Đ�=C~U�q'�[Pu"��FA�<�`�Z���:�R	����e�<����!4�P���E�!^�0x�g�<a�4�c�ǴH�9�t`SW�<!�g]6*���P �x��$�Z�<9�@�%>������s-�� ��AV�<��ެ)P��3)�9����P�<	\�G{dPB2 ҡy���3���w�<����x�>8w�4	G�8�!�v�<����p�r�Y[
y��
Z�<��m���f�W�6��dmPU�<�7+\�8�P���T�t�k�R�<���J�t��J�'��q4@j�<Q�� 5Fbp��𥝐e|�I:���i�<�@�?����H�'X��I���z�<�c�@�J�Ȣf�F�i#�EhE��s�<���ځg�$���e� 7N��G�Vq�<���>�m��� u��R�jVW�<9�8 �6qy�Ǧk�}�w��z�<Q��]F�ƽ����CƔ"uĕL�<���W2�x�+��M1d<��Ie�`�<�韞#��X�.²"�qs��R�<�"�Y�,=�a��'_��%N�<Y� L�d��R o[�\�=�.�J�<��)_bXXJ��^�xm��l�<97��7	�����'�VD�A��<�"!�]W���"�$Lz��0�~�<�ֆCh�
�{r��u��=�o�@�<Ɂ�BoP$�s-ΌP^�)��y�`I�t�P�c��(�
�bP�A�yN�G���rϤ*̞�k�oH�y")�+�Q�I�(D:�����y�*Ui�!#���
�&�ڏ�yrĈ="�^D�%M��L�����bA��yA�7w���c�;Lg��B$B�3�y�B�s��M*<�8���'�yr	ʵ-�H9�F@k~d�3��G�y2��2E�\�2��<*0�F�ǘ�y"��6=<a6ǀ�^%�����y",WqmU��v �h��J��y"c(?��Zm��s%��a��E��y�`V����hRI��?�ڼ�Ă\�y�h�J��<�բ��CT��Ч��y
� �zb�&ED�҅�5"�Ҁ�"Oj���I8U�H(�Х�+�&=ZA"O��2��;(��M�ņCΠ�@�"O����NN�@Ћ�!!���g"O��i�(��ػ�$��VE�"OX�S�%Z.��t�+:�I�"OD$3�ŮK_��H!���_I��[�"O����䉺nu�=�0����6|��"ODH���S�u��/^Y�ݚs"O�,�ӧ3)m
Y@�V1,�d��"O:]��C���q��Ͳ2��$q�"OH!� ���Y6�B!&"j�X�"O���`�#}���v�yd��1��;D�\ #!�cp�a�L�5s�%�p'9D�@�B��I�J�ƃ�` b���9D�4@7���A���B���0JFaԦ$D�p�Q懫vt��9�/�>_L����,D�b���� l���]��8�f)D���UG\�,���1&ʺu��T�),D�L�D��_�p����	� ۶���6D�� �,�87�l`�B��JB�_�!�E�|�R���o�/|]"PS��hx!��΁Bw����¬+T*X#ӎ�*r!���9��K�l[,Rz��ㅍ�!�dɍ_��ˁ�Y�=,����̀!�!�R	B��}Cc!R��e�� K�!���,a����"� ّ�Y��}b���2a�S�V�UO@�<,(��M8D�Lwj?r�
@�bH̶V
80�A7D�|�D��6��8b�H�|6�A�%e!D�x�E˔;'X�z��G�R����G!D��pQN�;�8��w��]���;D�xrm��&4���Q__ �P�;D�`A���%uFܩ�.��3�ؽ��>D��B�)э<0jhj�Ə"_��#0D��cΉ�96��@'M�)%��ѲB:ړ�0|*�/لN��aiS!2��ћD��n�<!GJ��V��0s Z�!�ÄDB�<�ŗ'�ȝ�6jU�6e�l��m�}�<I����N(<T�G�{1��b&x�<	� ���G��0�D��w��u�<y`��V^�%��ſ],�y���nyB�'tjy	!0*"�)��ϻ)���C�'�N��7��<V��d��i�"����'Xr�x��Z�O��l�`+��+�p�'�)K�D
�H�$E�PK�%�Z9q�'P���7� u|	Q�Ê!\,Y��'�PB�Ti�!+%�J�i�x��N>y�0�E�0;�D��$�:zr.|'�dF{�������eٵ���9���r�m����<y��$�n��:֣֩
X�i"� �!򄔂4d�4��-c)�-�v5�!��L�g�H؇,�4�e�w��(R�!�DX<Sh�5�ZQ~0��8�!�D��x��DC���bL�ܢq�Gf!�$�5|peq�H�;`@1w��4O!�D5Yi(�Aw/W({+~$ �5_/�'mў�>��F���Y�����W�E�J�D>D�@z�&[��#�g�4IXy��;D���j٧xlڐj�#V<5����(9D�����'%N�`�a.��h�3d!D���rJ�t`�P1SK�I&���A |Oxc�\�6�5h��t�U���l*D���'ʈ�x���!P�����S�<� ��#"�(T�L���ػ*�xX�"OƉ�n�)3�b�2��(*�<�1"O��Id�)���ìb��`"O�����Ǵ8z���`�
[���"O:-:g��.&*4	�� F/?�
�å"OХ�tM�g��*�@��2���Y���IqN�uI�KO�y��A*S�`�N�O �=�}��ܿ����r�t%�ЈK�>C�;k���
�۬Y�X��d�8`(C�ɚ#��h�)�,R���swg%*��B�v�ر�@L�)�@����!1P�B䉜*�����@�U����Jv��TD{J?��W��j˲��$EV�[VT9O&D��+��*u)X�����Tv6Q�":D��PB&��.L�8��OS0��A%D�h��B�d��s��:�D	��$D� [��&K�*,r����m�E$D��*gd7��A�Gs3�%a@ D��B���19����xȰ剗�>D����.W �㓢פ6t�
T 2D�4���6��3�LT�~�| 2��-D�� Dn�a�H�[#�V�d�6��-D����&�M�N��d�Ԓ`�� ?D�� 7l��i�6� �T�8�8�G	+D�ت���Y���qF��9h�����.D�(�z�� BDe�ZI�@*D��
�NY5JM��8�-:�&)�Ao)�$:�S�'j��(��E�I/6�lK,_�Ry�ȓB$��h�JƤi$��Q!�l���ȓY�������{O�l��-�Y$�C�I�s�rAQs�]UJh)�#̇-�FB�Ʌ6A�����,-���k��DP�&B�	mပ��À/������	v[�B��)3fL4q�.�&v~4`q�^�Wz}�ȓ�=�HN�,��צǞ�V�ȓ=Nu3��.TP���mX��ȓe�<��DIB���`0ED� *�ȓ�ԙڇN�u3n�H����RS����!��X��A�~(��R��K�Bp��q�V0�D�A�5-��'�M"��T��� <k���2�\�!�={�X��x<4�c%�me���@�@�	�&ԅȓx��(K�AP&XQF郳df��y����b$F�!id��t&[�7���(*x����)O]�X��Μ,�,�ȓ6�0�sC�&-V�k�j'yȓ3�ĝ���֋4_T��>0���h~�n�����Y&\�25����yrcQ=ʂ��e�i ��t)��hO��ID�4] �C�"H�@�n 9s�M	$�!�$�5���)3��'�&%��g�o�!�D2�6���$j8A�QBH�/��9��7�hH�% � �8aAT���\���E�c�.k0�D!6ë#�؅�<wh�Bf��#(��c��ؙ�ȓ~!p��ѧˎ|��5%�̼�DR�S.e�\�m���C��^�<e>B�	68ֹ;�.׬�ȡ�'"Q�B��1@���h6�T�`Z��rQ��3��B�;F4���536�����J3�jC�*
7�̳ ��8E�Z��Ծ_�B�I,Ɓ�A�AS�)O���'?U$N�_q\uh��V ��A�q�<y!���)� ����Z�@��dk�<� @�r���/�>L��l�E؈["OFm:P�]<������ �PQ�� "OJ��#OD&t���J])��"O����kĆxE�kg�#�n�<���Xb��Q0JB��a�h��ϓS���1���F��8�&Iеf�M�?�L>	��D�_d��3&hܵ���U�i�!��ZH��YUn,P�}y2'P)W�!��=P_�4�(�/X�y8��!�D��L��8��=���s��˦<q!�"Q����waS�~:M��(W�B䉕�� H�j[x;��׉�"^��B�	%���M�9Д��FD{~L��hOQ>�3��.�j�!������Q@>D���*�q�� `�Dgwl��:D���!ˢ(8�x g״�B���8D�h�C�I�C�P!�m�F�!�!D�P��`ɫ_�Z��b��]ʢ�Ps#ړ�0<��oD�W�9�30�B�w�<!B��k�RzC͇28l��%��q�<�s+�L��M��DۭA�pyB��q�<���=����ȅ-��0��)^i�<)�˴y���-��\�� �F�{�<ɲ,�B��T�f��5xީ��m�<a��o-2��1��l����g��0=	7.�w�D���kN� S�r��X�<9���agD4��ŅsQ�����O�<A�ŵ6���R��%+�B�)��K�<i�@����λu���he�p�<�@��S�yfcܺv�p�h�+�n�<�� �B~(ᰂ�ݲ%�`�Xl�<є�֕�`�z
Ӑ6�<���J3D�̛�4^B�8C�Q�;�z�Ĭ0��b�'����z���;"
���@c�&�k͠�O���hO�)��A��C����5T и���p�!�Dƹi��hc`	7a��9��X$�!�Ė�=�L-���F�>��9I���,�!�$�5=X�!�ז0� h{��I��!�ۜ{�(B���-��A�3A���X��(�:uP�?+m�V(L���{����=i�y���[��	)��B�(xb���1�yB&�W^rɸ7��H�Y9�#�6�yRˁ1���R �@��EyQ"U��yR(B��Č�����;\0� �E�y�+w��q�օ�.�*4z�,�y�Xp�9QK�5o<��������/<O�˓w)~�iB�G)I�zd��X�l�.��	�'S�j�D��o�8#ʏ�`���	�'�Լ�휷ܹA�
�#����'dv�� O:2送X�&QZ�-��'&�U��چF  �x�4CâT�	�'�h!�v��<�(w�?n�x���'Ҫ���	V*lԕk��32�T\$�X��ɞ>V��`�
ۨ�@�ifB�	�@�T��Gh��6Fd�1��:TB�I�Nl��IA��} ���ʊ;FB�IL�8���$E�P؂d�z��C�.�"�0�mN�
-q���&��C�	 b� �k�̾f�Qa���C�	6k8X`���" p�ٰ��-�XC�	;H�>i�Q�~�`g�V&SSzC�I�@kHJv��(�R]8&풠zLDC�ɽutDm�BkM*Y_R���ʒ��"O�P! `L+L��W�N6�P*#"O� m3a��3�S�'�Y4�x�C"O�X�wDˌx�$|u����a"O*1�oK%VD��$f't�U��"Of�r��M�*J�Z�$[Q�|�Ð�'���\�)�y�b�/@�P�:q�G���baj�7�y���:H9fX���rm��� ���y����
�H�C�
X�\B��P͌%�yb�O;�y`�H��͒�)�9�y
ڙP�^��0,�8�ȑ��-ȃ�y2I�
�B�*??h�ʒG���yB݈eO� ���F� 0��F�yR�̕PZ��$��7E�pI� �ڌ�y�B>5<@ ��<Tlݢ"���y2��V���y$�U�ʱ�f��y�˦R�$��gS��лu���y�K�Y�$Q`�ҏb��p5D^��y2iF�3�&H�`F:���$���yR��6zd���ִ�R#��>�yR��+4��!�A����MH��/�yIP,t�ҝ��H�c����&�y��9i�Tr���p��7ϊ��y2O��/�b�r�h�|X�Œ���$�y�H�M�t�͔�m <$A���y��\����1���^B�}��V�y���%8Q,���E4S�Țti��y�K�^Z�q1@�G5I����s
%�y2n�P���Qf�ٸHF��'���y"A�|���h�ˀ�o�T��@��y�
2Fh�R��:>��zѪ�#�ylC
qK5�Ơ9ܢีL�<�y���g��i�7��)i&��"e(J��'�ў�Ow2��1o�O����#D���C	�'v)��DE'_xB�)A�F-@�,Uz�'�x���Z"=��홧�\�a˞�A�'�Z���(m�J�-�3^��L��'�9���^z�l�@�\Ā �'�ni���Y�%>F�bЇ��]�����'����C�c���	P� �@��'�b��!� r��`�M?�Q��'`	P�ո�|��F��#G|q��'�:���e�'j�dӡH�� �]��'0�!�!�Մ#?`�{�#ڽ�jeR	�'�6�ZV
�
g@]�F���ܝ��'L&�؃n�J��;v䞣�`(�
�'���A4�	<Q
H�ŀ��J�B��K>ь��	�?=�&��af����3��Y�!�$�&&��͠���0�I��m�!�ę��D���%J�0�P����!򄑙*bj��GV�lz�&�!��s��9�BO�"P��. !��_7R��!�	З:BԨ�`�8;"��D8(`���Ơc4���ڂ �B�	R�A��IV ��Q�tLYx��d:�l�"��4^e�t���/�^���8D�`��['w��1��oǀ�0��(D�� V,�#]�q�� lJ�h�(D��a�)4q@	�8�����3D���S�LA��V0$	*��6i5D�08�+cd ��/&ar�8�b�&�IG���S �8+T/�,|]0��2%��,hB��D��D�sN*;}{�� �DB�8U!��P�`�p&$}����1�nC�Ip��|�T�C/7�����V yrB䉙O_>Y�qϒ[/䨸���S2�B�)� ��W͕5z�ma��M#L�e� "O&@�;Z��w�K;��5V"O`��D.S�]�����+.&���cg"O��r��/{|�yRAIz���"O��cY�A���Rbƌ"=mR4y"O�Eȕ��GO,m`�$ɇS��� "O\p��^�0�k��B�dJ�!��"O����MX��#�Ԩn0�`pW"O��S�b�Z��IF�M�>Rp��'���!&ӬM�0my���.d�� �(D�Ѕo^ /)�ЅCg��d�sb&D�D� ��rk��� �,q�pb�/%D���$B9*|;�Fރ?%L5D�����4V��fK[!��1I��4D����$�����bw��:nx�M��%D������'�݂�fZ�	��Y1��!D��H1�\�I족�`�-���b>D���ʖ|4b	�C������3�=D�L��]�M[����$������:D��BV��a��t�Q�ͻ
� �PM#D���FA9%[��˷��.3��TH#D����&?��}��oM6q�z���'6D� ��ċ4x�ȄS�=)"$x�# �d�O�⟠�<G�h*p&����I�l��<�J���d���"�n�n���/�w�<Y�+���ኀL^�N�D��gC]�<	��B�~��,��I�/H��2HYY�<A��r�H-�6)�)IꠙZ���U�<�N�1?Ɯ��
�Y��ij�!R�<Q��N"�eq���?��@�6��Q�<���Ӄ:3�T� BH?Q�E9 B�P�<�$��x�NḴHMY`;�͓Ix���'�@�P�E�va��%Q\g@�x�'�F=ZP���tb�m����Y�$K�'/��Q��q�2��J�.���c
�'S4H��[@��R�l�Bh���y��M���`Ѳ&O�u���憃��y�jû3p�P+
��k[ޜ�f��<�yb$X(j�B�����8v��)K���yb"-]�JX��.Wn�Ρ�$�y!+���D	�Z
���t�Y��yBNLj�i�0��.��l��@N��y�/T�h���k0�į��z�gK��y"%AR�Y81��!.6����y�L����@�v H�G��yB��A*T�#��	0{Hru8G��'�y��!��P���ګt��;e�0�y��C�N8�F�Z'�y	f�@2�y��+nH�xa�X'Tq$��y��ň{�x�	�h�[���S�
*�yR�Z+^�,�)��Ecb9��M���y�C�)��w��8�������y�C�#��3$�ߕe�n�9q`U��y��Y<ycP��E
YV].��קС�yRE�PĞ�؁h˟T�FܺV�_��y*F�+!�M�EvZH����y���/ ]��(�O�-�U#�0�y��I����D�T!FÖ�yB\��������=��1 �A'�yK�����eڧ^��A2� \��yb�XnX��3�
.�����\���<����
�zGM9B�J=aC]H.!�F6՘pP����0�����!�̕#p� �+B ?Ch�x�A��#!�� �!�%K�f(�����;	*��"OR�J�):_ H�KB`q�YA�"O����G�5$���O�zU"O���v"��|̬rRGݧ+H���"O002�6	����צ�T|��"O�٫�J<;4<��F��6ClD�"O�LI,��5|�BV�y�"O΀bQ�E&��i4�C�"�� gOv�� �ӣ_��c̹�jl�tj.D����(��7'ք#5��6�*h��9D�D[7�QD�$�����W�9�I`��"<�|ʃ#Q�5��(�REߨ9��Ba��b�<��nЪG	2-��	 &v.����V_�<)6M��D�f)��H� zRe�S�<Y��/^̶0(�̅�\�AP�Z��?ɉ��O��
Đ$��}�v�A�I(�)S!"O�h�HX�L$�A���޲qk�E��"O��H#NPN�ry8V�K�?�((�0�'���(�~��4�'q'"ݑ�@�(~���`��ʳS�nP[
�' �l�Ɖ�)~h͐���a,Ft{	�'
H�4d�	���S7��8[6H�	�'6��Pw��[s��[e\Wd��'�͘�h����u�غS+8��
�'3�)�#�J?����D�n�1
�'B�VM��.4�a�	��� �'ړ�0|2��ѕ<��|2N$ ��h1q.S�<���[�@�J�h 9:F��s�L�<yW*�6����a�)a�I�"Oq�<�%d�	0��2E����8�lS��Zy��?��:<�i�Ɗ� ���iӮ2D�����/�rmbthş,���0�1D��քӛF�(�1��V�(���/D��J5#�l*�v@��-m,���3D�0���f5�=: �_"����2D�D넌�~�x :�h�9��5�
1D�����^
���¾�=���.D��d�1�E���ZRN��7�9D�,���Ք���D�#Z���$8D��	q�Un��*� *��Y��:D���G��qz��6"Z�S��@��8D��!���1�n�x���r���C,D�����N�|��(�3��9EI��!5h*D��C��B�o��y��D��6�a��'��L��|�``Z: ��%��d@�c*(���(D�TYÌ�l�	)�&��btJ )�	%�OR�Gx�ʁ�ԃZۺi٦��?/BI��I����)��?=6��@�> 2؇�"���1���j6�5pS�
�P�d��k�4C3�Y3D��Q�INV�ȓa���0�-&u���l�sg����0%,�*�LS�W;ع�gҭo��ȓac������3��YUd�$u@���r� �+N�oJ0bdo8X�i�ȓ�&ekR�Yl��9��1.�V��ȓ]��������ը��qH�E�����!���$G%d�ȁ�U�R؄�-j���w��	��6ÄSCĩ�ȓ6�h�Ќ̐w=�<Bn��Sjܱ��gNް�&��C�B@��g
�(���OhU@ҁQ�v��{��2u�`�ȓE�ڭb3�5|��2��2`�����tAQ�(C����3�*z����ȓ?��d29r��R�S�(�hP��lD� �$W.�}�T��=�Ԅ���<� ��ҭD./jBi�`%F�X@"O�� ��1f@� ��0ڤx�"ODX�L��yW~��7 Y%i,:���"OҴ2��#�8���V2%N��5"O�h���S�"1,�-�/SJ�ذ"OU:����NoЕ8��	SR�`��"O�s��
��J���ˊ�|5f͉w"O�ӡ��C�x�)��B��h�"OL�)�ɫfQh�I'S!�5�"O
5JU��,�i���޽@���"O�Y�a�h���q�+um�4"O�Ġ�f�5#����OQ�s�X��S"O@(���Z�l1o�(��!V"O���*g����U���V���'��Ii�h�q]�Wb���n�;t��DA>|r�})f
�"x�z0iQ1U!�dK#<Ú���8=q�eP5� (G!��F�B�P$�!���B	�i4�8ڣ�'��IH�)�'dx5�v��07�x�pu�B�PS�'$F�0O>Bv�ʤ`E��8��'=�@��:K�v	��Z���'�'O>��P�ѡ!����w$�n�4��7D�$[�K.�l�ȧH	�h�4��e1D������`�_�@Q��0D�T{񭊓M�����-����,:�$/�Sܧ�p�q�@�N�̬j���,j�Ԇ�?��p�fŴ]��4ʤ �2S���ȓz�6�P�Wr��	RJP�b\���F%���rh�VH��a���@�tX��w��bq�Z%0��J��P�ډ��o�����
Vm�T��4�-��0�X0�G"D�DQ �D0P�z-�gɋC�E���;D�h��	��Vy��#�?,�)���=D���炌DUl��Tg[�9��g<D��0o�=@�e���ݽei�Q�g6D���B͜*�>�Qr�ތ@^]��8D�x�/�1t����!��8�P�e#1D��I���0f��. .d�0�S�#�,�S�'S���L�9����0�4@	4���'Vu��AEX��@��>�6���'�P5���կ:�6E�A���H�z�K�'��I���D�sL�-{��R!E��ٹ�'�a��Ό�kO��[��6�Fi�	�'Zrm�D@_4Gu���AnG�1ߚe�	�'6:�f�ՄN�ʁ�p���~�#���'��i��$ �h�q�
�J<��(O���d�Ґ� �	�aB�eW+h,F,3�'�f��잡 v����]<2�h�'�(9pJѵ*��!�DQlu!�����,��Ӂ��[���"	]h,�S���d�����S�L�:RfRc١r� ��ȓ]I�E���Y�Y��큷Ͽ&8@M��v�:��#��[�`LK���)�D��'-a~2-üHˢ�$��/XP�o���y��	�I��yS��/V�}{�Ɩ��y� X"SgpD`����W�T� �]��Py"Ρ� �� ٍ�
�3�|�<��J�s ���.��Q��m�N�wx��Ex2,(L�rw+N-4�P���o��y�˝/V"�}`,��lƠ �Η���D�O\���}�4� `�`��!(���,:!�D��;bص�㐸V�lg�>!�d8:��8	7I�3����B�̐#џ�F���	�l��B�O�����`�(�y
� 耋V�M�(��5""CM�s�F����4�S�)	�}Z
 �F[
,L�k3��*p�!�g���q�l��n�HA����H����\��h@E↬H�����&RyKH�R�&D��yH5i�E:I�cm7E�N���'T���(=�ZX`�ML�T�]{�'L֜$�X5ygs��� zq#�'&H�2��=dz�-��fy-�]�I>����I�$�-
�f�q�, �"�֕xO�'�ў�>�)�e � ��11&:E�е2q+)D�T$Oǀ^(�1���u�p�)'D��Ο��#�㐄@"��U�%D�P�q��>t���G 	�\-�lq&	"��������0&�u���\e�H���"O�)(�/P������ϒ)���y�"OS��E"f�6�­;q�)@E"O��
��S�������Q�F�h�<9�jK�n�U{6D�C.2��Ve�d�<�T�/�d�M%u�be��ƀd�<�&=\V� Uǝ�cތ8CF�b�<Y��4@+�)
@�Ʋh3t�Δg�	`����#*�~a�@A���#@�1D�0mK|��`3$�� �����j1D�	�M w��A2�H�{�~!�@ ;D�t ��
XF1��d(8�Har��>D��!��p�H�
5�R�gB����A"D�X��}������\[=R��E�>�	~���Y o��	iE��gNv�2 ;D�tx��XQ� ���n=����<���哿%�F�H���,�b���N~B�I��Jl`�-ŶCp��@��8G�C�I�F(0�)VK�ZH��HTC�	�)�伲5�\�te��r6��6=;fC��<jb�MH0J>Y���8p��%�(ZЦp��ѩ�O��rh�$��O�C�I�QV�D
�O14�ȤP���%i��B��. �h�C,S%g���*��A�l�B�I�{D��e��$.�P�F�@�d;C�I�+�H�!�E	y%B�Y�ߒKVC�	"l�P�3V�ʈn������n�B�	��:���D�>���K��[� ˓��>���BB�í�+l�r���yr�� ���C,�<xy�r�ne���(�v�#T�j6x(â�C���\�ȓc �m!R�E�8�b"�]�Q����ȓ�b�
�gA^1����/i����`�t���V�3���4� .SP��0�Xa� !<�$�"������ȓN)�@��-c�ј�!�B�=��a�0;E�ʻ[z8���S@��)��O<�8 e�A��jQC�ƒE,�ȓ�9;�%�J��
C�)�hͅ�)�4E2�-Ŗu>PHq�J��w1��2��8�Ӯ'�	�!�ȭ:�T(�ȓx�<�B�Z`LTmH�B,}��ȓ8���A���kL��[���l��\�ȓVU�83B	�wS�M1�i�0RG���?O�ݩVA%mlX��B3}(C�u��8���N�J{p@D)�$1tC�ɔLRD��)_'ʬ�)!��)pC�I�2Un��F����C/80=�B�ɅQ�0�bQh߼w5��pC��@�B�ɪv^$L"�g�9k��t� G�?2ЮB�I�6�b��Q�N����V�Wt ����7� � ���M4&<��$�%b�j���"O"���NC�5v����l��4f"O���sGJ�9���J�A����"O�A;�+k:������`���6"O�-�P�D`	�.���Pac"OlT��F�#F�,�2-�9��WU�\F{��隨O"ժ!͡#�B�a.�kRџ�E�d�ڍ9���I 
D54����s#���yr�	a�	���V�.U�)3�
M�yүT\�z�Jb���ER��٨�y�;�u�@dVa��!!�@�
�yrE� U�{+̨XS�\[��Q�y��V�����E�]a�x��C
�y��"�8���	l�����&�y�d�,6�L��3�S�d6��欁>�yR��b��{Ц�Y���vƚ�y"̓�v�a�S�D�}̀���lM<�yR \�6�)!�R�uJ�%�n�.�y�[���s��,c���`�j�y�M�	�\}��F�V�P;1�J��y2Đ%��ժs�B�:K�H���1�y�n�#'�"P��I5&�����y��G.���%Ƒ�2�ri�5�C��y�X��D@�5�F�$��X�%���y�	Q�B-eY�A�}k���2�yB)ʨ;%��Y�H��q{�-	��y"��ȶ8��3.y�)���y���=�@"��� ��q���/�yҭۄfо2%Iұ�����I�yR�����)e�K��d����\:�yr"S� �bS�ɓ!"a��U�y�%�i�|��@��sl,U��ܓ�y�d��3��r�Ql6j�`�N�y�a�h�@�D�ӥa���ȥ�N��y�D�p��5:�JV�kv�H3��9�yRK�|�ҨH�D֟c�쁷�^��yB�Uhu
d�`왈Qm��y��ƷH֢3 �%���g��7�y��_�z�
P
q���j��	��y�掺n5
�EOΆ���J�d=�y��J)8Ԭ�c��^q�M(+A��y�H���Y�{����P��A�!�L�$]�P���Q�8����ė�x�!�DW�m*��Vq�ș� a�!��D�Pg����-I�������!�F�|��}�����iYȉs��<�!�D�����	*5Kh�$�/�!�䑘w�E���F:\� �pl!�T�B� Y��+��x@��ce�.Y!��Bޢ�%*��H#�CѰYX!�M:I�ڨ*@�%}�Q���K@!�	ur���q���a��X��[!�d�&Z|.CVDV�_v\D[G��")o!�Z�s(�	����E�k!K�nf!���$�lO�	�q mLSH!�Dү`3��9��
0s�0��*\�g(!�$�H.�X'��1�JQ:I�!���F?����J6>��8(�B�.�!�D�#E�L�a���
�X�a��p�!򄕄mv��j��C2��u���q�!�dW�#J�A��@ݲ�+�S�ck!��-�N��p��6;�U����!��O0dLӣ�zS��
G�uk�!�Һy�.@���jF�9���f�!�� �tcU��;���b�i7�Y�7"O`Z�+K7{2�E:��ҘG�H���"O�h�P
S�����ѵ}�8ͱ�"O���u�ɂ���8ff��Sj���g"OXd7oёw�<��E^>~L��b�"Oz��t�S�c���y��;EN�"OX�ro��MZ�I�r�i���g"OHhh ��+Z�12��=�����"O�y"S5O`���s���>�2�"O�	����Q���S�朰E��8��"OLQ)@Ù��Z���$׫znB� d"O~5�_��J� W�Vmx��"O�\��>�V�r'�� X����"O0�yS-E"T$�M��.Y`@S"OX@+�bV�Z&�0���\"4D�"O0�R�*�k��� !Ĝ/�̝��"O���bŮ�PU��!#�J�!�D�84	�H0���\iR��~�!�DUl���5.EON��J� ړN�!�	56�p�Q�lκ-���K�!�d��+�`���m�"��b���x�!��}X80�c�	:R����Eːe�!�dI%>�Ԉ[�}DJ����)6�!��f�*L�)�C��z&�R�!�d��aj��ɰC
��n� !��X�!��$Db^�z���X��b͛kz!�d�.w$���h�w�  )�ɉ��!��G�.�Pef�$`xxuip"�Z�!��QVp څDԤ8d^O�!��"a_�Y�6��
gɐ�(��K�!�S�b���"��ĉ�V�!���@'�=Q��Q�h �X7 !�$WT�����Λd��H��3+�!��
�PQ���e�4�1y���@�!��!E��(���B�2���{�B���!�D�3 6f��BI<VNVd�F�A�!�dȻ�>�-��{��y 8d��'�mQ�ٓ?��n�s����'����N�e�M��?z��X��'Mx
b�]�(�f5G��%lJx�x�'��Y�S.�z�nE�C��i�8u�'1�1�U�A'.I�@��ቘ^�����'�y��fߣs����#�9��+�'�z}�KN�@,p<�3�
�	:&1S�'w�,�E��|IH|ڥÑ4�F���'+b�jP�օ�H �%��3Z���'G\5��O.hn��RO@�0[�i�
�'�6����H(l���Z�V��(�'?���tH�pB����P]wJ�*�'Ќ0Ă��-`�1�@���'��q��';��q� I3�#/�&H��p�'�.����oL�A���u ��J�'�8U�Q���Z�Z؊PBm�p�X�'��H�L���ܐ���4���'����"�ԔS��&�:���'EFDa6���o��z��Bg��yk� �����M
/}!4�ABL��ybk%$(h�.�u�>��ŀ�y�V�)�<�2�@�o�zȘT&���y�l�w�6䪰�L1��dCG���y�mN5B%�黰���*0��!����y�"_�O���1`�-���S�y��;C�p0�KA$o��u��ƚ��y"�^�d�i"+cزX��V �y
� B8���>U��`@B��9�xx�"O�00�'T)�PxQ"��2���"OTQp���#���#Vy��c"O�[5#��f~e@!���n�a�"Ora�Ǎ]����0j�<�$"OH���N�7.���mw�P�6"OT`��j�	`�Q�u�J,:b<R�"O�0�r�9g¢Ĳ�gPA�TГQ"O�!�#�Z	]��-J�&�b0z�R$"O�S1��>9
��eƅ���32"OܝDAR�lY���<K�tз"O��� �M>#dll{7N'�<��"O�����:B�X�D���"O�T`'��/�hH���'e�L�$"OX-C��"6@*@Ѣ�R]���@"OP�3W��=D����ң�_�$x�6"O.��SOƳY�6P5�M�y�b�$"Ov��B����J���*):=�C"O>���H/d�FXR�'K;jx�{ "O"u�D�H�g3�M��挛Q�F)[�"OH��wi��-+�*�Y8;��y��"O������Yz"LA�
����$"O<k���6-�HhD�֒@��"O`�B��S>s��`P������&"O�u��-{��Xq�HJf��h�"O@�� �Y���3�_/T�εk�"O����<�S�m"?�Ea@"O�)�O��5�8hptnA*�Z"O�@)��}��y`TO�08�eK0"O�����Y� �8��7"O��sw��;�V�(�틢��(qe"O��"�3�rբV��>�8�"O��� [( � �aL	x@"OJ�R��/����B�˗^��zW"O���p��UQ$��+.F��쀦"O�8#��H��T�P�{3�)I�"O���ǔXW���^Ū܉�"O�9�S��;�RS�M��9�:8��"O�9��7kBjԛ#V;,��1��"O�l�e͘
}���D!��_�D��"O���R��'�^��Z�l�a"O��Y7�T	-4�1шL�r��"O��aE58�C$
������"OyC6��Q,)��Q�$_�D�3"O���3O�����I�9tb@�Bt"O�-yB��6ZǪ��s���dXT���"O������!68�0�]��b"OVa�e�_nBD� G�
 x6�P�"OT<0㆛Bn��	�f�!l�u��"OZ xV��hf�}�υ�T�<0�"O�� �|#xL���!M>U�!"OBY��̗�Q"�Z0��u����"O���@"':����[�@��"O�Pbr.�"_�0��s�s�*��p"Ox@��+��c
�B����~���(�"O���͐7�x�ڇ /g>��Ó"O����ĕ#��0�NK3N5:�a"O>(���!]J\��W6X�(��s"O�ic7�Ѥ>����$ňVÌ�x�"O���"D�=�(8�a%��R�!�"O��Xp�6�uK0� C�*I�"OJ���֠6�(����7�r�"O =�DB�=�¤����3V��I�"O�	1 (�#{K�d���&�����"O� :�3U��- 킼r'�X.E���1"OLU�P�Z�/ݮ��)���(�"O0���+@[�������> 3�"O:��$��.n��d&��z���;�"O|ASgD�*�R�@�EX�\�L�#"O�JVφ<[��p¶䕂��5��"OP�ڐ�G��~ ���ybHO2 r��j�LP�I��DȦb �y�Q�0MpH�%��l��|q�� 9�y2G�~H1S4ȞQ<��ڋ�yb��AUxA
�e��9�ƅ0��ʶ�y2OۛL7��3� S> �%����y�N�%(P� �;쌸y�	�yC^ �\i`��E�/VR��$��<�y�ň�3�dxWJ)m�=S�����<9��d�Z��	c��/t7��A�@�B*!�DӒ�PA���сL3ޅp��K&!��Ưk�~�;�aE5)�� ��ς0!��̱&p	�bJ+Z(���MXn!��,= ���V�)��
0!�E6C߾�з�V�h���j�!~!�dJ�zl��G;dd�p���!��[lp�35�B9Lu$h+W O�!�Y�� �1d�Ԅ:f��D��#��9�O�Y3r�	;GL�JE儷u�Ayc"Oj4�# _�;��qPv
�'LZ�pЅ"O�Q�!ٛS] )��e>B)H�"O���T�M: Eq�g��t:�"OjqtG��A�ES�KBxP��iᕟ�����������GE$�[�� �C\��"O�y��{+:!���$T L���IC8�P�3m�g�$���Mx2��<D�|c�!�'IJ�lK
�$0�UX� :D��a�K�&�jmI5+��}�xpp-}��)�SSs�図i��>|���P�(^�B�I�>IČ�b�\�k^$ܲ%!'L7� �dw��P���Is�D tf`'cYS9N"�UMNB�Iv"H�s0�T�[����Ѐ�~jt��'�ў�}jhԳ+�}Q�M*q��:U�%D�0kUD�#%��k7��֙YA�$�$&�O2�y�ՆP���W���||���|��I	�y�S�L�J�Zq.��iGQ�t�7D�D���lw�0Rሿ6G&��%M4D�`*��J�4��#��6u��<�q-2D���5+�c�F(S��EwTI��:D������.b�Awf�������#D��Ц���Qɕe�j��ps6� �IB����N�I������J�
TbV� ��3�JB2s�H�B	,��qF�- C�OrZ4҇���.�HY$�ט4�(����s�l���ݼ-D���L�2�,=R��?�O��B�Y
� ݠ!J
��gD&Q� �nVab��	4|�S�B�s��	{�`ï�0>O>���i�$aٿ6��Qg�`�<Ia"E�X`�1IAߒ"3��` ��hO�F��� ̦m�*�@�����C�ɣ�� 6h
9d^�(�� 	?5�C䉍^򾔈 ���>�"EJc�T��C�	������&�=�ެ���?{H����>yӅZ*8�ez& �Iu�u�GO�W�<1J��/�1r�i��z��,;�+P�<	���SL0@T�-F	#S�K�<��A_��5@F�&R��(
#E�<�m�8�Z��F�W$+)Nt��Eh�<� ��S���	9V�Z��Τ.�|2�"O�x@�"VG�6�A@@��Q#��0"O�Y�WAC�\�����A��HU"OL-��MbI��k``B���ڤ�x��'���g��*R�2�	:��y!޴�hOQ>�Γ��TkZ�3b}p���%����Z@a'��.����G�i�D|ҷi$�D-���D�rQ� �Q�DWyz!�(Q�����(}Z!�X0��Z�Q�uh���n��d�'�ў"|���h���"���E+���EA�}�'ў�'Iz��打�nw��C���HCҹ�'��~ҎǜB��U#GGFp��H� $�y��}����T�1hp�d��1�y2˛�>,����ʅ�*�,d�Θ'�ўb>5rt�I2�^�s3H ]���W�;D��0�/V+5��S2-p� �ҧ:D�ظ��ע>R��Y�A�FeF�f�2D�8YdL
:L,vh˃��(K3b��pb0D���(\��$êb;JU�A�1�ʈ�HU�ao�G�* �C�j�4���"O¥r��z0@`��#�E�t�Y�<E{��iIPT쬹%�;{G�E9��X�!�D�,W�0	H�(�aY��"Uf!�$O�lnX&,Яf��-q��ޗT�!���1��9��J�%y���Qqdˬc!��*k_� "#��w�b��F�.����S��yr���-��Y�� E8w�f�!$V�ZW���)��$C��v&�_�T��!��E8��>�'�S�iA�H]>qyc��P��jޏh!�d��S/�KƉ��3���!!�J�Tўl�r~BS�,�'i(:T� �.$��Wb�Gx��)B7.��X�"频��}DRG�Ao������'6~�J�g������Y4,�)r�'�F��f��sA]ƛ�/�h9�',�l�b)P,.��ԁş,w�բ�'v���w�J�x:\Ԋtmq�UX�'J�0$)��.��@ꔸ7�p�`�'�>� �"@	 ���H��D�y��'�&dk���f*�M�������'s�i3��H�t�^�{��@�S2��
�'s�� ���P��T�2
�xd|�J�'E�d�tE��U�2 ��p��'���JS���;�R�k��z����
�' pA���;-�4zd XC�TC�ǲʓ8�����.	
x��ꊝ.j.p�ȓZ�ԥa@G]��� ?4���Tר=��_�%�t�@F�/�H��IN?����{�0!�fq��lO�hO?�,R�L�1���ܝq��׈�8">9���Ճ�تr�_�5�t1�l,�!�"<���('�
��r����ɂ}���.�S�O��A@�jn(�uU�_X�e���)�`{��e�ފ��A��c�X�b�'�XF{���7it$������x��̄��yb������ 0Pt�tk@�y�X	JN
 yp�0n�l�'����9�O�P;eę����䏚%�p���'n���=j3ci���@MP�Ub�܇ȓq��+�'��=�8c�bP7�l�ȓ`�z��t��D��,����5n�J�Ey��'?��V�ވf$��hҤ`�J�*O��=E��o � �JTbގ_�԰s�O׺��B�	�n��\�0��!ʂ��"I%
0D�Ov����F��-a��B9���rP$�$41a~�_�� P<x��3g�����"R76}��"O L95��uRZd`���1[����'��	�!d��03OD�$W��r C�/�B�	�>�p�GH+xV<z�͓�R&�B�	��$�r���)7j@H��M�=��B��9RN�� F��l�X��g`�C�I<R�60 ��اv/z�a�	 1s�C䉻($)�R+}\H����I�h5�C�IC��l�eK�/b��A�\�UފC�I�Hh��R�X�igB����C�Ɇ[�&��#��M2�^!�B�	0��YZ��	�j�ݓ�H�7al�B��7wYH9���š#NԽ[�#X���B䉴
��ေJۺMu��V,&�B�	���&Y�̶���,�=A�hB䉕cB��!
§=� �gl�O�fB�ɪ$�(��.W]����_��ZB��,��6���ǏՓL@�P��8D���WK�0��S�녜�����J)D��c�܃W��(A��?X&�`�F�'D�4�s��8D��#���]k��B��!D���bAXo�p�@�a��v�;&&?D��z�CќyIx�A��7+�v� �=D��AS*I,޺ъ� >LRta7D�(��ǌ�^Pz�rE��"�"liti5D�(Q��ɶޘ���H��qy�	6D�D�W�ř�t��@O�f{�ա��2D���[=�H�R0��	�E��yJ�)9�D��d!��M��M���y�,�g2�Y3( �}����w�ɨ�y2
�(��HA$��C�x*�˙�yB��S��-`�lV�F(b�ghB��y��'+*0����)7|d�b"ã�y"�@��=�4$L����$J��y��\3T��w��p����gW��y�%�1_��Q"G�6|�j��F�#�yR�ܺb�Vԡg�Tvs����y��XH���V�f�p4Q`N��y�%���<9S��d�^A�`EP��y�*�,{@�cL��_*��j��yB��W�nl�W�H�[.�}�"ڽ�y�cŘjz����ٮ
i���6M���y��^�S�
�X�L� �%�F��yb�-K��x궋��~�L�{t��0�y"��=>`11QG��q=�2��ybF�|��hPOZ�搡�*M:�yhE7C�`���M�|�~\3)��y�.�pP!o�+n�6�#�(���y"J��f��aaE؂`�8j����y"�X�&�<�#��
o�^9�'+��y����vQ� �E�g6��� X��y�O}ztHD:uAl�xCˇ�ybBρJȀi#�����y!�
�yr��|� �2T@�����q1���0=Q�!��\�ބ` �F*���.<X�85(�[Lj%���Do�<�a��!�ʙ1GX6O|
�
b�`�<iGϕ�T�C����G{�����b�<�A+��};r�C�Z�TtXIw��c�<�da�!$?�ɥgF-'� U�r�<��\�D��k+V�K�H��+T�<�Qi�/S���r�	å\�i@�Q�<٢�K�e���'�9Y8��� OH�<�7�\*u^U�6/ʿE����TCGD�<q�C�&eءj'@S7,APyP��i�<� R=��Z�w&f�y�"0�c"O�E�Bl�w#�)�$��8r����b"O�pSA�J;�R1���JݎUS�"O���4�ҍX#p#c�9o�>A��"OV�hN��3����Ě8bj�$"O��J�JA�Z��sTgˆ^@�"O���JV�lFAk�L��cN�L�4"O����΄`?��Ґ-0�U�""O2�ƫ��^1�a9�!�!`\S"OP�&O�Rj�0�Fomx��sS"O��c&���V���@�?KabXu"O�̨�܁5�4��O��02��)�"O�51�c�m�.�&D��2F���"O�y�׫Z,��H���,@9�"OV�3�Y.l�$уu�s*h�'"Oz���F�9��x� ��c�Ȝ@�"ONL�a�@�0�R9�g�&s��|��"O��&僿)�V�r�a�7m<d
A"O��!n̗*aPS��kX�%�a"O�ᒧ'��qc0���g��I� "OeY��ԁ!ڲ��' �B-S�"O ��ǈ�#|�*�:�Föi����"OԬ������X��d�4�,'"O�����&m�0�a�m] F�"O�Y��� �Fl9J�!R�T}�E"O��3i�|��4�iȺe����"O�)k�F;d�M�V'�bz�i`a"OR4A"g��[��zP�@bJV)�"Op�8�M�
�$�K��@N*�)�"O�yz$A��4[H\��fW�HG�IQ"OR��Łލ]jNFZ����¹�Py2kA,K��tp�Ͳ
��r��"�y�M	"O���B�
�|��F�yRA�8�؃ŧL�c(Y[rF��y��#BLi��<UŮ�H��=�y���>�~\C�
-U�ZPq��E(�y"��4r�>�)n)r%�}R�y�c
�f(K3�W�9�D C2�B��y§�:]�\ճ��!M:\hIŮU��y�
�")HUY��5�0��c.�y� f�D���F�"��ɂ�N,�y2�@-2u�5%!�^%����y��ʚc��D��� #�D�H����y���ETQ�D�Q�%��y�2Jѥ��ɣ!I���%�bX���S�׬|8�APDSZ� ��"�O��+��x���g�\;��hِLB�f�j���Px"'!Z����@�Pu<��ëٞ�hO`�a!h 28�,x!4�=��A�A�+��K���)�B�	�3��|@�O�-mBH��M*t�����Bpf�&:y��S�OB�f�B,sDB� ��R,0�"O�*�F��E���� xQ8�1E_��*2l;8�u��g�}�܂) �u�v<bĦ�2pF9�):�OB-! �.����
�M+��)F�ۉ9hأb��,��B�I�;R�����XV˟�N�~8��4j<b��ck"a��L�|�бgH���g�5h=�9Rf��O�<Qd� /�n��Ȳg�D�2��Ο�2��{2�;���ty�����
#�`c&�y�L�FFE?s�0B�	�@�x��T�TR�hX�w�;t:ʓR;B�M���Ó=�H�F��n�ޤ���8.����IP�����?R�� 0����QأN��k��3U
O�=��L��Jf�ݰ���}<������Nπ��D��M�Q�qRc�_(6�AKFR�|���ȓrNl�3va�����Sd�,1TT��9b��J`���ه6�L�7��0;w�|"�+Z?�y
� dQ ����1jG��/g�Y9`R���T(�t�x��	�?�6T��oN,1 <hԌ���$���ѳ4�`$� Gϴ���p,��uR|b��+1�U������x� ɛI,�y�Ⱦ�%��*�O�xa� ��2� @J�nM�����I�n��dz�h+P�W���l��O�!ۣe�0>!VǏ�pj�@�9a�E4��
cp�dZg��㒄+�.�A2�$?�֎�4A0�0F�i�ƭC�\�q����v���J��'<�iS�[
��`R��z>`�E�>�2e�%`L ��)�w�_H�гI��Y���<���� ���N_-l)$�p���`�X��`�Y�J��x���k<�uS���*a%2��'KZ	�<��#�=���Z�ة.In��+�<���3a+Y*�?ᲄV9�(�����O����=*�s�J�;�R ���<��u>��t���h�}���_�g�T=hO| ���8�إl�&G�x���� !h�a�N�	^�jtZd׻��<9��P�q�x����M�u�)�����FQ{��F�|z��)� �28=�u�Ow��Q��݀y����!�A�`��B��5B% �)7�S��$2O�X��ȳA&�[��H�LY�		�0zb�S�S��8�5,��!Ċ��0 "$$"�P�	���'��0`54��h	J+ZMJ��W�{����c�Ƹ�	�����F Ou�'l�IK#�%9`8����� ?�Z8ҕƘ+�����&����Ņ~������H�\E��XJKZZ|�w,X(���O��(l�7hµ*��p��Ԗ2�X��'ՠ\HF#4V\�H3Q��#��� J�c:�O�Uc'�%Z��ʓ�W7%k��"%iX3p"x��
�:�hQ�fȫS��xRnN�:���P�T�F����;_��x��@�.��H��:���˭�V|q7H�(|�ʁP���w{<���BH�]y`ț��V'��T �Į)���$W�K�)�Yq�q���	)�B1i"BA3� �EG�����-�#.3Q���ܺ����R�:��0�[+�� -���OV��-f�P7C�4�������"s�6�YV�Q�
ɪ푀���9!F 	'ꃜe�A��I9}B���X�X�ɛM��)C�
����7	���Is�,���	
W#����A۞. \cK����Reb�N�݉ bC'5�X�A�=O���W�0źc�؂~4~�Ȧ�D�?=Tl۪O\��D+N4f���"�B�dB6#3�V�*�E{���&ڻe1�B�I�hm�P�H�s���G"ZF�O
�� �&SRm�F��$<���!����	��3�'�3p�����Z��y���~����僐<>Ll���KٵX6���I��]8����F:x��M���L�xB%�g?��Q�M�#X��;� 2D� ��L/��`�φ2;�p��]�*��p���̗�`<��aOgx�i�!Oa��*s�L4n @�;LOl��EIJ�24��-��~AP��H�Ka�DeH�g 89#�m14�X$C���zrn�,�M�d�,�I�S��`�&�#A�� �� V�]���_�E~�T�N	%�B��=m*Ra�#�0̄��JN�K���ÖBՆ~3&[H� E��'��|��K�j�2T�A�%��R�'Ŭ��,���%�D7w^
�h�5���ق�0>�B͍�g�:P� �	KgfЈeH�z؞�)!I���J��']Ј!�ڢ"xs��4�M��'�<��mݤO��|s��UC�L��{�jǆ"M(�(��)m�>aqf�Q7x{��As+�-YTx;fL#D�L�%�в9��B�ek\R�B��҆_�;�ΰ��D��(��I�E�>����W� &�#�%�7��B�LW��k��>%��XuZI�h�$��P���3BNL�԰=i0Ś,��Zv��/Q`����B�'�(�zw(YA�P�Y���1ED�;sn.��k��햪qO~�ȓr�Hh���zD��2��'4 n��'�b �s���2�a��G	?J*����VY�qxf%���XI�H�*"���>PL wK�-i֪a�B���� ��
B�4iߊ�8�#�4����X2�.Ɇq� ���3"�~"g	D�r�R�ؓZ�\1��,A
I.$ �Ȉ�%Ӏ)�%-������'ne#�F� ��#u!��L^ޜ�����qe<�h`8S8<�E͈J�D�Z�d��@CD��IF�p��*Ǧ�y���]�,@R�'	'=���@�Ď�~B�R39E&ٱ���&r����n�OQL۳d$~؍8��&V%.�*
�'w�X�� N~d���'B�Fu)J��X��N�:0p��r�'�6�stb��)7���m��M��ɡ{���D.ؕ�,tK��л"Le�"�9IÒE)!Op�)�/����(C�N%��L�����3����-aT��P "���c݁U��,[�Ł.�!��R9 ��e1u(=|�r�����, ��ɩB�������D�)�g�? �dD��5�jhp��ܙ0ư+�"Oڬk��^*�ktǃ�'#���|b��&!���3��T8�f�b�Q��HĈW�2C�ɂ�؝Їo����)t��e�C䉿-��[��|���#o #f��I	�' D4Y�!σn��M�r���W�)��'8��Em4E�d��1��I(J ��'�d��N���8	�)L`��'� �2�o�ck�]���M	�܊�' �(�D�	5p�9�d�1����'Ef8x䥄0�B��3*�J���'��%;VDI�A�N�J�쇶u���'�^(��Iݦ|��Bu��5Q����'4izbF�e�l��d$Q�x%���'-�t�6�Ůk�b}B4H{G�)�'�����з>%�hh�l�zK�S�'Z0�{�xtqׅ��t|���'�󄆙�;z�a(K%n�TeC�'iVѻ��K�p�́۱��nk�U 	�'r�b%]�q�	�蒰Li����'��ԉC��3#��a &�K�X���'~���m߫AY�<f$�	� �	�'������#R��D�O�H�5�
�'J����gϒd�*�ptb'Jp��r�'��h��c�}4�b���\qf%j
�'|�a���Ma���է]}<}K�'Cr�	p��d�4b V��x�'��9��~� =�4$׻t�
�'�\��Bړ;�b���=F�n)H	�'�0<�僘�e
f䙳���^�Q�'h�H���%oeZ#���xP�h��'g	���!�&B%��t����'��u���ټ�Z�Q1mܚ`��5�
�'����V �%#�҄� �--�)
�'��k��ۘt̮��1�.PP�:
�'LA���\�\E��M	�����	�'4hĲ d��YE�9y�Usp�"�'���!ҭu­����p�'�\!�Vm.6�U� ��l���*�'�]@��{�RM�6O��1�N ��'K^E��G3G�Ѓ㈨�TP�	�'͠yB��/��(��C	Nw:Y��'���hC��u
�u�狜9��'\>���@�EX�m`�-(< ��'k�)C7+�!��_�"�@<[�'c��P�CD+jL� b�wH���'��{ l΄^~�rp!C#�Ƒ��'y��o��J���� 6P���'[2 y"�%v����D�:��''r��e$��{0T��R�{��H��'*�Xpb�q_�\��X�$�>4��'� $�@� D�� ЇH `���p�'!�	iRB��-(�w���0�;�'nҠ����J�\����(��j�'�u��E*(�6���9{�x��'m2�W#��Gbb)Uȕ)2����
�'��ȑ��N���A� 6�:9��'߬����� >����+.ٴ�(�'�*	xN�<h��Qj�j�8���'�ƽ��)[%r_��2ދTXt�'�l��Ŗ�F�8�2(��d��'��E��;Y*�&�@ʉ�'��Y�RC*].���L��o$Pɡ
�'�8T�WF��~�^j��aM�lk
��� ̹Ғ+�8FB��X�Ŕ%M%��S�"Oz�@�*�j���a�z ʕ�w"O���V� �t�c�qؖ�V"O�1��)CM���� �2ʼ1�"O ��)1>��*�I�/|H\��"O*9��n�:!������w^��a"O��	w�͓*�d`�ߥtM�ؠ "O�0��C5_�\y���,J-�x@�"O
�+@�Z�/N��T�D3Fd�"Om;���#.T%$ y�v��"O�Ĩq�Ӎ<Wxk2�A�g��<c�"OFђgn�;�0�r�Qo���Y�"O,�
f.W:)�|���̕�[��H�&"O ��T��Y/� S0$3z���KR"O���6lJ(G�́�G�j��P�"OJ�	Tȅ
KD�]h��?Y>5��"O����,�1i0�iAZ	{)����"O�tB�o��+BXhh뎇f 4�k�"O -[��G!ph��h3(��d�]0 "OR\ #�Bdx�K� �z��v"Op��h�Q����&%J�e����"O����ӾtR(j��Z&��Ĺ'"O�8B�C�*V�r����p)�"O���FD�p3� �@/ёnA��"O�!�1M�P��t����	��hu"O�`r���y4]WAC(p�6ك"O���QCJ�/���b*]u���!�"O<�񈂶4k�̳W'8�:г"O�$�A��&XU��S��=��"OTXQ�D	(|�r���)��@r"O�L�2΍�F�S�&��v́�"O��d���[$�E9t�My�"O*G���'L�X�D��}0j��"O$��aiɿU��L�S-ʮh����"OD�rF�D,J�`�p*� s� ��"O8� u��G�2i 4J�2zN�C�"O�����\�Q���,7zM�c"O0l��#ƍd�Z�k��r:.08!"O��O�b�Ʉ�F!r��� "Op��%L���U�f�0*j��b"O���#�GC0x
��C5+�����"O����Hī\�6����& ��!"O�Lk�Пz�ґ+S�O(b.d�e"Ox]ha)G�blHhc�g�jϞ���"O�u����A;�T�e�|����r"O�MK� �T�$�I�W�{N�A"Ob��b���]��E�79��鸑"O��BӭD�Zt�ǡߟ]�{E�>�4�ÿ>��#���}b�K;O�ve�B����>��	�P~0EO:4Xr�!x�}�P�^� #z���
O�x` �	vG��Ö��+�^����I+5�Ard�.ഡ�|2C@�YMT��� d�֥S��JM�<q��c)�Ap�d>M/z���m�ɟ���RA�ɓ�"ny���΢PG��$:O�1C��={ B��3):&p�� >v�p�z�MZ�k�:˓y��y��jP4o3����_�@�b�mS�\ ���-,	ER�����BF��e�լ�Y� �*C}�P�C-h�i1�U<�B5��Q�F�$��c�R�'H�҃���s���I )b\h���͟�Jb��o^�N!��'�v�h�ʕ�+�`�������B�H�"W,��)�'O�<}�_0%��!��&��?�aJ�'鞱ȵD��n�5ä�__AHh�'+��J��S�}
p1��'g�M+qM�� �z��-߲z��5��Y�ds�f�f�a�߁v�D�b]}��B�H&�� �B�C��8�=r5�9zdi+7�	+%>�񘃊�c�� �7�2
�4��!L<�<q��Kv�}!��(DgјE倝gP���� ��Rd��ӗ�����'�L����Eꈬ��?�r�A#�o�P,�1&�-����'9�h����0p�z�n�!c��ж�C&qd��@�ˎ+�p>��Q�8��3�#;S^�� MC�������`��٠�%�����H�+?���vE��SB�\Q�M?�+(���)��,Qv(q�m
���K��8�1`F�#�615FS�乇ȓg� Ѓ��?��5���òi��l[!&�	1���3j��J�48���v��~�'�9J�>���L�7����o^��y�GN����2bE�#��[4Lĸ0}��Ho[+&\�|X⏎�@�P�;[��OP����A-0@j4@f��%��d���'����@�q[�|rRm�-Q�pX����4��̀C9`�6U�T,�>`#�'|��j�"��$�@�"�)G��L��OA�ь�Q�f��k^'N�C���X,$>ɋDF�~������ I}���5!D�\�A	�b�z5�QE!�}���A��x� �FA.T)�Ԃ['+���ytb&���ۚX��P-�=3n���n�!�R![�\��)�FOx0P��q�,ʔ�b��6j����CTAْk-�E~�ń\�~���.�0%��=3V�9��Ov}Õn�RȚ��7Ly��ޯ|���" 6T.y��Žm�<�ar��-�	j��GT�T��G� !!�b�'�Y����E�X�����W� ]��LkB��z�P��xuz8
�/�#7&�0"O������3���%(Q/%��Jbd�k�)�`�O;Q��b��!A�O��r���:JGV��yV�ڕ}i�`V�(�O��
�
��w��f�
6���06�Ǹeޤ@+W�Z�b��pc��'$l��ب ��hrs�	Ű����d��a�����iM"V ˪�pe��l_3-l�e�J2	�ѡr"O������K5Ȱ0�̼c�.X�����!�Z{��Y$�"|:Rl�,ʡj�H�D��Jcn�\�<�`�P6:�9֢�"A*]�_ܓ�*iY��/ODU�F�R�v ��#��fo=K�"OR�Y`�3vE�p@� J�A�Ѓ�"O���%Dc��ٲ�i�L@�q�"O^��b�<s�r��'��"6"OR����1PH��cD�P�LD�a�"O���sJ8��mz�cp	��Q"O��uÞ;S��a�5Ȱh�"O�!�UFE !��Ic!�1V6 �@"Or����۽v�
�P�	.>L.pc�"O��)��G�+�0���?<�t�0"O�������D�Ae�߽~"<X�2"O���v��&=��̹����x�:�"O�\�ރo�L�kGG�$R���kQ�'��5����wua|�eҷdV����E)Z�rT+�4ϰ=����T�`���)k�\�`*:A[th�U :�X�"O��c���H��}['��8������D�D��UQ3��*m�"}���s�P����Sb�L�KW�<A2�f�V��Rı{�p[�� ���16h*�剛qBQ>˓��=�U,�?����&��`�"O�)p�d�Ҭ0I0�@<,QZ�9V��UH�ћ�M�4̇�ɨx���;uIMt0b�"�6#�l�?1ƮT%lZ �aԈ.Ԕh�ej~�I�^
J���ſ��<�J&D��[��%���8W�;&�� �J�>���8 b�9�G@�S6Ɲ�+�O�� �A��	`e��Ȓ�1��'�C��]�	Z�3$�N>"� ةPa3!S�e9��ռA���2�����k�@U��qTHZ�}qLH����e��ن���u�}�fF@^�Z�-�.�|����L�\��o1b�|�b��K؞H��-e$��N�B�"���D0�5]�鰒�	�@�	$�9?I ����pYb��)(�T����M��B�ɇE�"��f��:]~9��DՇ]���ɷAc\�2� &�:�ZE�C�M?����15*��ǃ��qFxl�S*(D��07��+cd�H�P $X |Qw�;}��L�ED�p��N�w�����NHR0���+u�P�`8�Ol(F�Ơ�� �����U�v4����
ؤ` l	>/!��]�MkdI�e���qttQ�@��\�Q����V[1	W��4q!2�U'mo�K��h�!��P4s�@��AB��p��Sq��(f�:U��s�)�'p<�1@�(�%a�6�H�Ɋ� �0���'_&%�� �y="	"K�3�"�'� H˳2�ay�H3V��R�Iөd`(�r�@��ya�@!���Ӧ+�<��mՋ�y���-t-��%̞<�9� ���y#D�0 ��
!M%t�@�N[��y�B��G�B�c0'OE�����Ò�yң˄NdȌa�l�-5�p�GS�yB���r�.� �e�$cVIQ� �&�y�Φ~�q:С��r 	3m��yF����%�-	e��rb"���y� K#���ۢ��X1@��y�+_]�Bp�
� �֬@Sm��Py���)\�(W����BYISJ|�<	f �gqH�AVT��=����x�<	�č]��!x�		 ��hf�}�<A􊅳1\TBF��iD^`@�$��<1@%�m1�!�� ʽ<�(U�#+Ay�<��왜s~ar�]�k�@(@��y�<QQ(P�qd�M.w�h�x��q�<�5O�+	���£�+QD�)Q�eQm�<Y���Eє����Κ]�$0d��A�<�4�G�x&�b��A)uI�̐���|�<�kιպ���*�v�������p�<1��(I��K�+˥$�>�@$es�<�+��t]��q�/w�dPeǊo�<	b�H�z�:�aŞ&/��%ذI�i�<9RgQ!th0��0��A�.ɳ��Px�<yb�[��ڤ�Q3R�e��a�{�<1�&�U�B�
�4S�����,Fx�<ѥ)N�N8�=��Z�H�ga�{�<�Ci՘ �tpQÄ9j�^�V�u�<A��t8;���j~AX�ĝt�<1��[(�H��߬|�&�[u�<I�f�J̘�'�$X��@���v�<i�g�k�h�x�JEӮY��+UO�<���Zt�h�X'Ø2�	�6��L�<�Ҁ�!b�u��-Yd��'L@b�<1�J#��5*�Gǲ,�"��Q�<�F�X�=�X��79 ��kW-�S�<g,M�0*��Tc1:6`�B�K�N�<��Vd�2�׻�F,b��N�<G���[�.Mu���&� p�<��#/p���t�*Yvt��`�q�<��̜;c�eh��ZhAɦ&�l�<�1l��\^@y*��u[�m�T.�j�<�Ƈ;)^Qy-aΕ{6�a�<�é׫?V�i�g,P+���(�c�<���4F� x1d��D���ȏ[�<�f��+vik6�I�āY��D�<a������W�/S�2�S4dq�<��(�7�@�6Dϗ�&�St�l�<� f܆4�-�T�ê?)ڝs�mGW�<1R���?��	�t!L�n�9���N�<i��"� �����LlF�b��O�<a�a��]|&qz�.E�Jv�Rw�BE�<)4E�9�r��V�VĊ,b�b�n�<ɢ,��1v6@���.�����L
o��t�,�`a�X�e��b�¥�``�� v��h��"��;�D6D��A��<.NQ+�����Q�(?D�� Ѐ#����$0��3x��Z2"O�8�s蒈��pv��p4��!"O���,N�[�@=�HlV`��6"O���a�Nmd��A�w%�mq�"O|Q���YR�$���Q�|"�p�"O���{����B�q���D���(O�O�n�3��w0��&e��"�����'�"����X�)�f�E]��}���4��!��Q/\<��V�>o���I���bX����O���IGR�Z�bq�٣A��1c�b��Ov�(���&�9���Fx���������$��-���-q)�P�ӂ+I� ��z��/Oa��o�?�`)ӕ��>&��#��o��d�+6�d �:�a�lf)����(������;�8!&�x2�/w�uJ�'����G�'#�f����6*l!�'G��j�C"mVܦO�O�f��X6PN�`)u52������d�� HQGC��)�'xIYj4��5"bj���s5�����%F�h\+2�&}
ç %�a!3��zxf��*��4��B"[�2Қ�P��p�af/�h⓻;.���Q�6`#�ɆV�꼳�R���Г&Xa���y���H�ݟ����~�� [X�Ca(�m�L�,x������M���:-�����OZ�>��2HXdL����:P�WƮ>�2Cڅl��4Xġ�>2w�)ʧ0f.4�A�ʫ_�0!��;$0�$�	#嬸��h@�Jj������f���'�&�Bg�4**bp�6�Ϯk�Lp�J~�N~��
�xH|��#H��D���D_�<�%��	8���b��S����s�<�1
�oo*�Z>r�l�)�Cl�<	��
�N�����]=:�L��1�l�<!��]J� M�s��4`���M�r�<���ðt�Y;3��
z�uѷ�l�<٣�[���V�0]��0	�A�M�<��[4��9aP��1<�,%!&�B�<9pDǬnK��2�'��~��!1�h��<)R�kfH��v���d`z�؀F�O�<A�[�Sq��3��R�'�D��!�D�<񗂘7T���UL�%}O�,;���y�JL�1���34Hx�d������y��G����QϬ�U���y"��Z�Hh˖�ϯ}�	�Я�y���/w�jUi�Ɵ^����FA���y�&�dfP���M	#w.Eqc��7�y"+܀M� �i� w��"�ܝ�y���r�%i�Z��sg,m�C�I/!ڈ���M;%��
��ϖF�vC�=E本�)�&v�|�t�Ni�rC�	�Z�Q��BV5�2���5n�C�ɗ1LR�[b��&h\�bV�ο\�B�	�9�Pa%�:��	�7%�	v�&B��?:����)V�[b	�?bC��/����j�], u#@'��b��B�	��D��LK'P1М�R�(�B��/2�4�
�,։b��+&R�Q̪B�	&"�\D���4�љs��a>�B�	6�������/K)����شC�������d�:ƥ�:D�DsdO1��P+����n�H�.7D���6AC j�LP�ȩ/TB��k3D����!�|�r�c!�=:�>���i?D��y�'ɩ��H�m��q���2T�,un]� ��=
�n��?7t	Ru"O⨹��

<̀�#�m��W"O���H��:݃���Qإ)""Of�!�.�WD����D�+c(!�"O�HS�� 9q(��a�M�h^�u�"O��z�Z�t���riAt�[�"O���� ҕ_ۦ��d�-��Rg"O@�8�Y1r.`�T�эt��1"O� �4�CE+}��u�B�T��yS""Oh�y�gCSm���/�n�6�"O�pY��%����X�OC�c�"On�Ss�X�=�"U���L/P*0�y�"O�=@@o�uȘ�Ye��9)�"O0̙e�/56����D8��"OP굆gHPQ�,�1�~4а"O�P#��7��a�fтJ$"OFU�1��N��5i
V�D��"O�1��1n�F�BEh^6����"O����g�Q�g�08�b}k$"O����G�L���Ir��4����"O�dX�e @�D ��  ��YZ"OȀ�n��el��Q��%dur�P�"O��P��s�Ih�J��[lf�"O޼��Η����ש��<W�ڠ"Ob4ad���y#�M`ԉ�8�X��"O��!�CF��6]��GJ���H�"O���&@�%!!j��E��'V��9�"O(�sd: v�eQ��Y��
�xe"OV���̈.G�4��P�� �@��"O�Q�OP�_H*Y�p�
o[ 0�C"O����72�����NK�YHw"OVM�roԥJ� m21 A:M! m��"O�Qu�/�����ˬ��~!�;K �uБNF�<��0�'�q�!�$	�.�$<)�Y9��3'���!�dF�[Z��Q��C�U��S&��.B�!�Dg`���f��6��!w$ɖt�!��$�`ͩ!~���+��#*�!��7�z�5*+P����¤ͨJ�!��"|HPxq+�S��SA��,#�!�$D�8c��1�!v�"��`��3v!�$�QX��i�K��x�d [�`!�ċ�0��i2�$�����y��y�
�'ҕ�RF��%"Zg��i"��y�EI����!2+�-H Tx��-�yr썢W�4�aF��75E��0dϋ�y��E �F̰��R<_�0�C)��y��G�o-��p͂T����RO��yR΋2h�45��ݭ|4hM���L=�y©� U~����J�hpW�A��yrmZ�k6np
�B��V��Å�A/�y�!�`��$W�9@�ٷ��yr`��,�F1Ϝ=1-88�gE�y�͌�S��{����]���Q���y"��~1��Xu.�Si�kd����y2cY'n<���.7E��r
��y2-+Z�x$�@a�C����S�y���qެi�?C���B��(�yBN�VeD���8��(�rM��yREΉ5TYs*Z�;�>D�R�ʀ�y�D0&��ǫ�#<�� (b�!�ybρ�,`�H�.DFdDs�C��yr��9|�Zvk��,ê��k1�y�O��~���&B�M��9�nъ�y�i�001��Т�(@���Zt�	�y�JG#q�"�BMD�A���ԄC��y��~nmjV�#4�2�Kq�y��!"��y�aC�5�8� hX��y��ٻ&�<�J6CO�Ap���{���w�Rx�MA�.�4�q�D �X��/�. i��@�i]�y؆�E%'���ȓ`.��!�\�t��iĠb؜u��S�? ~�bS�
_F}�`-ӕ!����"O��(�)�0&�>T
�ֹ?�
��"O�Af�5K-�M��O-�.t5"O~��۫o��:�j�N�D`z�"O�lj1玠RvlUk�Èr�~X�V"O��a^8|�ȸ�2����x�б"O��ª�!#�,=KE�h���"O�Q�P�v�ܻsOW7)� 9"O�<	d*^#�^�[P/�>3�%'"O	[Q	��'r8����4t�
�t"O�ŠP��0�nХ��*b-��"O~�Y�&�f�ܬw�U�F7�dz"O(���[�}��-�a��?MM��"O�]X6@@7|�9��d��!
��Â"O0ԙ�c� J�.�cb#Q���I95"O�<�g	��r񫍇G�T���"O��� �CH��}�J��E��Ł�"O�(���	t3���띲3�̵�&"ON��1d�y���Vj�/�@��t"O@a7L�j��U��j�����"O!�#��>(p��	�{z}�@"O༲�a��9l�1s�ּZή!��"O:�k���_�r�sK�h�q B"O8u���0lJ�W�|��p�v"O��GFRH�yӤ�)}����@"Or���EO�J��@9��P:}�%��"OZI��N�Q����& [�wa|��"O��҃��G��Cd�00�"O�D�1d�:�@Yчb�$U��Y"O�4�!��>�2�"ܞl.�-�Q"O����%�)XE�ӷ F+Q,���"O��KS/=�88c�� t �K�"O,�y$�"mtP:�х&}�MjC"O΁�6�8Q��R0(�/Se�L�S"O�8���U�<:AA�FE�L^�#Q"Oj��@��ep��`E�[Iʘ0�"O�Ț���7v��4�T�M/J�
�Y�"O };ViF�;J&h����@�:�*!"Ori�@c��T���5B&[vB�R"O�{�d_1dt�B
�h~�m"O��r$�ى$q:=�R�Z��B�"O�Mar�c~*�BC�A/!�9�e"O�6fG�uH!��� .���"O�a�]H��҂X�Yڶ"O�ܪ0��%	�jp`p��)<���"Oօ���%+"h�[�K&�8E"O���R�:s���I��٭=#�(XG"Ox5;��2] �[��D�L$]�1"O�)CU� �9�|�b1üJ$�PCV"O�y�R���a<v�(ш��?$,5�`"O���b�V9b�� �w(�#?n��2"O�E��PL(0�&��=!:|¢"O��;��5C��88���� �"O�,9��0]���zgkU$j�
�"O��Y�◜�T���$�q��@:g"O����cD`t��b\?|[6��"O`�P��7r �g"�!>�b0"OLT��.�2Ă��=l(�	��"O�h�ƎP�'n�(�֑��y!"O����HD�<��ɲ�w��H"O���F��MR��cC&^��)�w"O
Q�Q��e/�a A��-9��ѡW"O�i�e�����e�����B"On��e��{�$X���=i��� �"O� ���2!�
yO2�:�/�K��=��"O��&$���)ɧ	R�g��P�"Of���nYN��7Ȉ�`Q�d��"OF{��.��(k�P�856("O�AB�R%-���D��=~,��Q"O�)����r�TPE^�Uw [�*O����[Z<���,1�@(��'�,(&�I'a%���M�8pH�'�4A���T$���V�6�l���'���2R�x��H�R���.�*U��'g��â�� v�Z�9��)pE^L��'X���%�W�^�Q��v�����'�f�dąiN��P�̕g�(I�'q���i�2�#���a%�a�	�':����T�&���e�0QR`�q	�':�p��`��J�|¶
�U��\
�'8l��g�@@(�d��g��Sc��H�'�ֈ!tυ	���{3JE*W�6���'�$P#䏟{3
a�"	�Zt�	J�'�	g'0I�A�Q�>���'xn@c�+ ���G�C�IBh��'R�zS
R�6���bg�=�.���'�"=J�	��T�Բ-M�5S�'���Fo�?>��G�����|c�'� -
Q� Y��![0���'>����3�N �Έ� M��'�~F�M�Qx��'�ç�|���'L���  ���   �  ?  �  �  �)  -5  {@  �K  �V  bb  �m  �x  :�  ߊ  ��  ۛ  ��  �  -�  p�  ��  �  ��  �  w�  ��  N�  ��  �  [�  ��  � y I � � w& 2/ 6 t? EG YN �T �Z p^  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h���)�S�	N(2P���W-MwR�pu�
e5lB�I�d�U���5��ag�=v�C�	�u�ҵ����r:]am8�C�	�S�A�O�9v�`��%V�r��C�I �,�aw�0�ȸ`�n՝mbB�Ɇy@h �"�5��,��NרS�B�I�|9�}�1�7G����ӗ(%�B�I�q�# ��Y6D�)�iVf�C�I� `����>S�N�T�5;,�"=y��T?��V�B@��(cȄ�L�x�:A�*D���L=2�0< 1��zj�H�6D�h(��:'���R�ߴt65C�G9D��zS���@v��ѫ�	,n���6D�t ƴTؖ���j�J�^��5D��wր#}x	"�d�:p��5D��c�O[
Y��,����O�Y��>D�<!W�
�#�U���H�!��37O(D�и ̍f�V�(�"R:�0�%D�(A�j�6*��H�.E�v�ܫ�?D�8b$�R;y�lqy�9?��#�d=D����d�r�GO��a��Ģ�L9D�`��%�6U*��Ə�ݖ< �5D�@@�l`*8�e���d���m!D�t�'Ċ2F���H�9�HHA�>D���4(I&u+�Q:ӯ�,/��H0�"D�@b1��55If1p�n�$L|�$�'"5D��X��̚2��!��
C}��K  D���6@�	e�P<��'��{�\$�#�=D� ����(g������$c8�1�:D�TXfJʻD�1A�D�>C�"��G-D�t�V��Z�t4�`�[����3,D���vݷy�$�Kb�+���GO)D�t�L��%N�-�w"]�F�d�3D��0��ٿ�:(�7�Y�0�Y&�=D�����E6XJ�@��5^�ӷ@:D��+_(7��q	���0p8�A6D������eqHTqc��}*�u�u�6D���F�@�{�X��E�H�|�
 �8D�0��� +��P&G�>I���6�5D��ɦ�L�=� ��a�Y���C&D��(�A�1'µ�!���]	0��v�$D����Ցv8,P�`/:�^�s�H!D�P���;xr�r2C�&
~6����?D�D�Ū6J�E3����&$`�,(D�����Ni�9Bj�G�2(!��$D������R�D�`��09�6e�a�%D��+w��33�x�$@��\c��#D��G�S?/���6g\�6yά
��&D���֬(~52��Z-����q�0D�T�VoF��iہnX-uNH{%O9D�0 ��_��@���=w ֝`c)8D���q��9"txlZ�eY<{�j�"$<D���Ɲt�L�;[�1�A?D��)�A�w���2�c�[̘�4(=D�<r%_�{�Y�݆1 ��c'd>D�@��W�P5� KZ ec�,�r�=D�� ��p�<iR����Z6a[|�3�"O�YVgϼKUX���!�&n(�ȓ-����n�%]@,��Ɗ98��ȓd��@�ɐ{?��8�׀h޵�ȓ��h�V���PQv�!X�ȉ�	ȟ��Iǟ�I�����ݟ@��㟠���.`�.&n�Nͫ�C������џ�	�� �Iӟ��㟔����]�,"��F�y���8v0����֟��I韘�	̟x��ݟ��I����I]�Hu0D�T)�b��``�gJ�L�������ʟ�	����쟘���d��9;nL���{��a�0;W��	�(�	ٟ�I����IПP�	�����@n���'��	)�#R�.ݾ���ٟ��I֟�������IɟP��ɟ��	c��I�6M�j�^h	1��1afe�I��H�I؟�������IƟ���۟L�ɸ\Q����L�2e� �B+T%*��E�	ן`���@����d�Iϟ��I��l��G���:�&ދ6p�r1f�r��IӟH��ҟL���� �I���	ן��ɐ0�v�A�NS�y��A�ς/�$�	ٟ��I֟8�����̟P�I����,Y��Ǆیvk�M�$�Q�P��E���8�	ڟp��՟��I�������l�I-d�<[�^�Z�9�b�;��������I埬�i>y��ٟ`�	����I��&U��Ŗ{MЅ���W?_�����Ꟙ�������̟��I��x�ݴ�?��4|dɁ�X;7�����%�@���W���	Zy���Ot�o�@p@t)5��,-q\u�&D��
=ze"$?Q��i�O�9O��$^�q�\�h���w��:��B�wb�d�O�IXT�x�l���������O�L��$���/�O�K�h�*�y�'���l�OΊ,q��
�f,R�($��.4'��とb��q���9��M�;�|<ѧ��
���1���6F����?)�'��)�WP:�nZ�<��$σjLR���_�r���0���<ɞ'���dL��hO�	�OLE�g�"$X���d�9%j��0Or���?ڛ��S���'�(�%�`0�D?v��{`��a}��' 3O
�#
 @��!_VJ����X��rU�'�i��g���r��I���ra�'f2�Sӌ^$\D��M3�VTCqV���'���9O���M/Pm�ͣtD�3v0���2OP�o	n�I훖�4�Z������㰴[��	0t���0O���O����
$6M,?��Opp�)F�������R.ڈ��l�k�PI>�/O�)�O>�d�O(���OP�+!�Ү	�%s�N&$fb�E��<�i22I8#�'���'��O�b����rA��6@���嗨�N��?�����S�'fK����T������0���J�H�L�,4�'�m�u
��ph��|bZ�l�0[,�)��%Vg���	�H��П4����wy���<M����O���N�7,�-��L�xR6O��mZx��`b�	����'�0Y�����Lw�z*�2�`	ٳl@�y^�&����EgO8M���!�O��ߙ��
��bj��7�ި��z������IɟP��۟��d�]^�(q"��!�*�M�3���Oo<	<����dQ޴��/'TĊ�,�br�!pr/����<q����D��-�6m6?�r�C,G�h*�ۛ"�pmk��#	�H��Q�O��aH>�)O�d�O@��O�i`(�*�rslƾ�8� ���On��<��i�0`4�'8��'��^ذ�]'rl�"C�S�|�E��I؟ �	M�)��eT�r<�A�҉Y��h�thؖ8Z�5h�"�s}4q�/O��?��I6��K k��Xx�j��K�^�×�L����O��d�O����<��i@tc��R,[�T�i���CD�v�B�'�7M3�I����O����V=��m��^*]X� ����On���! ظ6m<?�;��e��'XXN����Ӣ�u��y/��h@�ԕ'���'��'��'�S:B�4�
Mp�Z,�@˚
5m�=!ٴ2������?1����O=�6=���(S�A�r��(��A(yZ��!�K�O�$(��]&@�6m`��;��n}��g&���ܫG����y�Kމvp��I�z%�'r�i>��X�L��O�,|�Խc$
�<3�q��ǟP���D�'XP6��`�@���O ��D�9��Ѷ�ӞG8N�Q3��L�B����Ox���OF�O�UR3�!�B�g��*רL�V����S�Ĝg������/�Sg�������u�d�"�Q&�a<�}#@�ߟ��̟��	�,D���'~^����xEܙX�
F�g����"�'��6�� jR���OҜn�b�Ӽ��@� �����BܲF4���?���?�SO���M��O�� �,S�����7� �e��a���f�'���ٟL�Iџ��Iџ��I�*�|�%�ϰ��(�յa`Bԗ'��6M�9�����O���8�S@����ÈO�\l��@��3�@�O��d�O��O1��� ʳ'�<��+ۥW+tp�@ �uf�7M5?����I���Z��Gyr��x�
4�0IM�9u�=��
�+I��'���'�O��I��MkEE��?�$L�:A���C��4Y�#��?q��i�O��'U��'�"�4�<dA (��/���*U�4��@�i��	�T�J����OSq�F�� N���iD�-���Y1 m���1OD���O��$�Oz���O��?��3��@�胣�U�k�p����H�I���:�49U�������۴�� �����\ f{�!h��S��b�JJ>i���?ͧt���۴���%4g���r�ʘ3����`��q"�Y'�۝�~�|�]������៤���UcA�q �B��wR��R�P�IBy�
b��p��<����	Q�\rnL�`��f#�Y	��Y��:���O���'��?��	9�P�y�疞�*l����Q�;�e��1���ΌV?�K>YQŃ�3��٘� ��l�A��?����?���?�|:*O�l�:�(͋gncݮh�Blȭn欝�ã�}y$k�l�\��O�D�,�p�M�.G�I���F0U�$�$�OJѻQFi�N�Ӻ; ������<I1���6@8a�F؍[w <
�@�<A+Ol�d�O��D�O6���O��'N|~a8���G߮���Li� �Ʋi�aj�X�T�Ig���<
����k�����ȝGL��*�?)����S�'}��Q�ڴ�y��C*Qʔ2'��&d�J�T�y�L�7s^�I�DI�'�	ҟ��I+S^ �Ad�+6�	@P.-=,���؟��I؟��'$�6\�TB����Ol��SD�p���I������.�x���O����O��O�=Ȣn�; W�uC�N�7X͆X������ƫ�xbų��8�S�|"��� �
��'�\t�1 �._{ݻ@Wʟ��	ݟ�����4E�$�'R��#)^ f� Ƣ_�1�����'��6C�)�\��O��mu�ӼÇ�M�B�|���	�'~�D,��Γ�?���?I���M3�O� ߀�2ӯ�)9��k!(: ��(��nү?8��O���|����?I���?���<��ȟz�̩F�H7$��@(OdMnZ�#�)�	����I|�'`���v��+N��"���Up���P���	���$�b>��)R-X�G�E�f��wK]=<x0 "u6?�%�:py��������D=x�t%����#���ZE��< �����O����O
�4�\˓��C��}�b�0\� ip�X8SJ�r�/A�|U�nӤ�\��O��ī<�R`T8yBFL��[1&�����M=�(�;�4��D�6,E�0�'Ӕ�����2E�T���3!���.ˎM��O��D�O���OT��;�ӛ�JHq�� �� sn�#����	ԟ����Mc`���|���Y	�֖|�c�!�hěfM�3��b��;�'����To6Fx�D��Op�B2D sR���� @C��A�$�ŝy�^�'I�'.�	ҟ��Iϟ��I���Մ�p�����I�4p��I͟(�'�r6��b���O���|���G6�ԁ"��j�	9B,Ti~rD�>9������ΣX�*��	��Ւgc-:��<:D�[�9�)��<ͧj#��� D��h��m�&�c�(�&U.]J��?����?��Ş��	Ԧ!{�hB)_��v$��`Ur�Ys�:W�$���ڟDJ�4��'����?Q��փl� a㏄�Yʸ� d���?���JX=Yش��Z,RX���'���J��L�%.x�"�*��!}���Ey��'���' R�'��Z>��Gӄ]�D���U�{�<����K:�M[��Ĉ�?���?M~�s���wF�DҰ�MN�h�Q�
�@�a�'K2�|��ԄA���9O�iv�J4
��@%�8��p)�6O�Ds�AB��?�0$��<	���?���\&xǬ��n+�d����?���?�������k���ǟL����Z�⊖�V̊k�!c��w��a�H���Ɵ���c�5?�xe�dƊ�N	� ӆ����$��zx��,=F��|�e�OR����{B0Pa&�H��L��

8>��8���?���?��h���d߻bC@Q��ZiMt���gD�����y ��IΟ��	��M3��w�a����fU�9����@}h!`�'KR�'2R'Z������xA)��Z�$!@��p`�O����EeS�Vu%�������'A��'��'��p�B�%U�!��@ ����Giy2�q��-��<Q���'�?��⎅q�DX�ud�eo���#��B!�	ޟ(�?�|R3lR*;4Abt`���qBG�:O{�`@���
���	
�,�m�i�V4&�P�'r�I�4F�=eehf�Vp1*�#0�'F�'�R��tU�D;ߴ>~���Nx��t��:gάCVCA�i����F���D�E}��'�r�'�lXR��X�6��%�P=Z���V��#!����d��,������)��Ԝ9*ל��x�U�:���#s6Op���O�$�O����O��?��N��i�W���w E�d��|yb�'�~7-�	y���O�oZs�I<G9z�re-�.�>q:�Zi��'����̟擗{���oI~2�Q�|@=@ހN����A\�'�VM�&�$�Ę|�V��h��ߟ�9#���J�2g߱Y}rX��ԟ��	dy"do�d����O$�d�Oʧm�`Ԯ� ܁S�B�17�)�$����O�d�Oz�O�S�6Xq����9 ��k�N��/
�=�o�,
\��� 8?�'R8� 0��wH�� ��	%m���2�>ݶ�Q���?���?	�S�'��$Ʀ%0��¾V�|���H)o|$�fL8s"*��	ޟ��4��'�T��?9C.��/�~�so��2� 9���̏�?��@A)*ݴ���
�E>����'��3� dر�֋$E�,��	Z�J��2Ol˓�?���?	���?1���)�!#��cc�8O+�%�C$�6~��lڊg:n��'�2������1Z�9����``�1���R�Б��{�S�'P�jxߴ�y�*M(�ː�������y2�/N�M�	�!�'��Iş��	�iD�lK��DMD`�:4b�K`M�O����O,�d�<A��i�F�*0�'*b�'��Șf���G
&���6r�����LZ}b�'J"�|RȖ�E.���&Ĩ(�N��������M�qQ�U*r��<5'?��O�Ĉ�9C$kA�L�zeڑɒ��*��D�ON���O���+�'�?��	[,rX;�f־#�Ԭ�Q���?9B�i�]�W�':2�rӜ��])4+z�K2h�;����ѣL�,�	؟p�����
P��٦�'��(`�	S�?���͊#s$�A0&�?�h� �	q��'��i>y���P�Iџ���"T��'��D}� {�F<f
���'9�7�34����O��/���O�`a�� 1!
�j2M�*���*�!T}R�'"r�|���� �
��a��00��J��=wX�r�ia0�g6h�#Њ��D%��'^ԁ��J:Kh<�D�Ğ�}�A�'�"�'������Y�ث۴Hۊ��#�8T!wB�2w��8�S �{!9��/����I}R�'V��'�<*w!� aen��-��~��}��BH�Gқ����k�.� >����	��&��#�><�2�H��0V�dJ4O����OZ���OR���OF�?��Z=~��Z��#F���w��쟠�����4��̧�?�5�i��'����� �=�.��2���i�@I�p�|2�'B�O�����i��i�鐖bսy�:�Ï�)�V�Ҟ	?R��I x�'=�Iޟ��	ǟ@�I->��qq�h��?�^��I�U��0�Iܟ��'��7�W���D�O��d�|"�
K�V�����ӾH���K~�d�>���?)M>�O�&�[�m���U嘍6.5�l�7!�x`���J���4��������O<�v��.Q�<a3bK|0��)w��O|���O��D�O1��� _��IȕsH�3RH�	����	�|��0��'��m�8⟴�O���ўo:9�ԁV�f�P�s!��(��$�O� �gt�X�M�u �	����O�<t�4)>�2q�Wd�7dn���'��	џ��	��p�I��(��\��A��V��VO
�'>2\��lW.X��6mM8Q���$�O��D6�9O��nz�]�R畗9 ,*��`�"mhc��x�?�|�[hi��4�y"�ܗY����w���̱���I��yr*̂�~h�I
i��'��I����Iv��s�����92w���j���������	��'��7��:x�x���O\��޹G3(q�M�&�b�3%KU7����*�O�=�I�}i�5�ǡ��X�l����Šk�����r��$�\��O~*2)�OV���: H����εkA�Pu��h�@93���?)���?���h��nZFȴ�JR r�,u�5�Z�G����Dߦ	C����X�	��M��w ,���Ā)Q� =�b�Z���'��W��Rg���'!����Q�?��a�8gt(�w�Ќ-���bEř;o�'��۟D�	ȟ$��ܟ`���>G��ra�,v��,�§O�H�'�x7�tD0��Oj��7�)�O�m�I��B��9A6�,B:���.�d}��'�2�|�����jqJ�hVc��M��ؤ!BR�֫Dʒ,O�ʊ�?a�&�Ī<q�# (υ6s��5���Bj�����?A���?Y��|
-O^�l�+y@���'!h��!��گ��l�(J�<�$u���M��>����?��@t�ى2��j\\0rn�����kJ
�M+�Ox(���Q��(���Y�7��9����#f��V�:\\���O.���O�D�O��"��CB�Xi�lȴ+��燛a�V��	՟|�I �M�ч��|��b_�V�|��
�e�XX�v� H�Be�ۧ��'�����t#׻oɛ������n��Og��P�I��6u<�hDDܔ*5,,�$�'��%�(�����'��'��UR��ב%���2�fě��9# �'�]�hR�4q��S��?	��򉛈^��)��B�L�9� �X`�D�OJ��?�J>	/� �D�Iq�`,�7-<Z3�B�NR =!����|�Bʪ<��'K�X�D���0�8�b!2�XR �_�M������?����?y�Ş���馵��*/��1SP�ϓh�R\�7)@1A�P��I�L��4��'D���?�GB��V(�P��n��y&a�v����?)��Dt��ߴ���
"���Î�4lˆ), ���P����p#T��yP����ğ<�IɟT�	��O�:4y2 .�J`#.*�`�hѪi����Ԣ�Ol���OΓ�j��Φ�]�7F�9sF�-K��IQ��""�O���6��i�Z@7-s��'�������e�=Ld���o����o�1]�$�ĭ<	��?����"�X5SU�L|�^ypo�?�?����?���d���! ���h����9vmÏ:�TyA�M�iHڬs���_�~�����Il�I�I1��A0��2q��X�0G
(��d��� �H�QD��|B0�OP�����|��W�U�ؐ���`����?���?����h���G�*La�-��2��M�v�������ǂ`yreӦ��݀8f�z�ʁ+���۾T�f�Iٟ��'<�#�i���00	��[e�Oc�� �i�f��8�Iq�NU8'�,��46��<���?���?���?��B^6K�T�Cm�7ey���#������c͗Wy��'f�O�B�Z0���p���)_��Ish�4����?����S�'�t�p,�2�ܬ��#[�@��s͜e����'�<�Zǚ����s�|2W�̫ �LBȵ�t�(,78I3#	�����џ��I���SWy�
a�j��O�9�F僫No�0��)N�cpr��DO�O�nZV�
��I̟�������U�ޠ+ڜ���Ҿ(����D����Ym�u~�C�""�p�G�$�w-����
!n��h�L�6+�t��'P�'���';��'��A�SꓷM̌�	ȅ6z�"�"�c�O6�D�O�(nZ#|�h~���|�D�;v��׫V�8�\�;և����'����$
κAk����@:��:up��� W�@��l�`��0Z!��[G�O0�O�˓�?����?���}
��ҦH�*�*��M��n�By���?�(O6mn��[KpA�	ğ��I�?9�4Fj9��m&��x��&��	ӟ�'x�|�[>y�	�ӲH�G�'f�Q�7�˯U+z�)P.�,6�4s2�	gyr�O������&��'F8��l�(��z��>.�j��b�'�b�'	"���O6剒�M��j�e��P���X)Ub�����?��H��?���i�OL]�'���1����`���E�y1�E���'>��%�i���:|r>�`6�OT�'HTL�Dٱgt��wհC��̓��$�OP���O����O��$�|b0���P��c2eM0H��ݒ�	>%#���#{O"�'�b������m7�	�#�	7�p=����	��}�	ϟ�$�b>}��PѦ-͓`l|����Z�Bb�=�%��(��R�<��n_Dc���`�by�O��V޸���Q"�f�[�O_�v��']B�'��-�M+��N��?����?)֯�iߜY�����1f��u��O��'S"�'M�'�t�KvN۽*NYXB��%O����O6���*		��i��?Y���O�:Se]94I8��c�B�R|�#N�O����Od���O.�}��h6H]SF�Z�
L���Aĵ�l��@ԛ����:��'�|6�1�iީ���H�c2J��C':���z�bw�d��՟��I>�~�o~���3b�����#\Ry�S �>Y���ZprD{ҕ|RU��ҟ$�	Ɵ��Iğ���#j]���g/	v��8�"HVyB�q��@�,�O��D�O@�����:vo��H�D�|�T�G
ɡr)r��'���'Jɧ�O Ȭ�`솋H����!�c0��t*K�
�l��P�H�PÓ�-*�BVR��lyRNC1��y� N�U<
�c������?���?���|�-O�Tm�����ɌF\"3���!4*���`ױ9e ���"�M���>A����DP7U~@!�<|и�&��I�0�QGl�r�:H]B�`�Z�O~2�;�:"U��t�6��8��͓�?���?���?�����O$�$@楚���8t�L+G�� cR���	��M�!���|��sI��|�Oˢ�% O>�T)١<T�O>����?�'q��!�4��$��m����@�mn�����&�(�S����?�v�6���<�'�?���?�1Ȟ+!�İ0�.J'�N0s��ۨ�?Y����mJ���ß,�Iџ��O�0��*V=8b���NW���O^��'����?���ť��͉���Q᫙9YLP4
���� ���dh�ӟx��|�Vs\0� �F �*�<�����;'��'M��'����]��)ߴn74ik�dQ�n��������|���ڶ�?�� ��6���o}�'cl�A�#O�ƥ2����#��hy�O�<1�֕���3�E�p����\eyb�Kt�y	ݔ4l�V�	��yrW���	Ɵt��ڟl�	ʟ8�O��1+��9r�<p�,L�PE6i;5��On�*��'���'��O�"er��nJ�+�ءdڧq� {�i�9�f���O��O1�TQ��Hcӈ�I�n�$�H:N�d�APH�3U���1A����$�O��O���|��3���QĖ��DDq���7A Ȥ���?A���?i-O|Tl,4l�,�	����B���Њ_4Q�b��r��:DXz �?�X���IT���uP5f�I����d@�j���'�YQ+N*7�1¦���k�$�6�'���/�1$�Ib�ϕx���'���'�R�'��>Y��3N4LJ 	�()#jD�g�ͧ1CR�	��M{����?��l�V�4�Nعt� _C��b%2FU|�XQ?Oh�D�<Q6C<�Mc�O�!�U�V��tcг��aPu�Ԓg����v�Q^锓O�˓�?I��?��?��J��pbI���%�Ӝ^�m{.OΌn�'h
�L�'2����'�x}j���#nP l��e̞8��X0���>���?�M>�|��X>Y	���2��/j��u���/ָY�����$�sB�P���?��O��C� �kb�>�愳���RP�p��?��?y��|
(O��lڝq�n���Nb>��	�O���0�7�I��M��bj�>���?	��CRv�Iq�7o@�����3}���j�M;�O��3�fҔ��d��4�w��%S��J#o,x�����MH^�h�'��'���'���'����dlS�/�0�"HQ,�9ѱ�O8�D�O�l�x^��S�$!�4���`q���Ҭyw~y+�B�q�,0�I>)���?�'o즴�ش��F8p� �S�T7!l��j�p:U�����?AB �D�<�'�?����?����Jz�,b(�*�uЄ��	�?����Φ��t.Gty��'��<BtڝMxwH��� h������O��D�OޓO���t�J��Х��$^J��ϔ���J����BN��KB�3?�'���ċ'��)=�A��g��\��E�2^l�{��?���?�S�'��Bۦ)�*H:����q�2|l��4cV%	�����ϟPs�4��'�꓊?@�H%8L��,.I"���Y)�?��nV�L��4��$0����l�4~�%R� �"R���J�Ӈ�y�Z���	ǟ���������O<h4��g☰���߼u `�2��l�@��¬)��d�Ol���(���O��nzޑf����hs�F�(���b��%���i>U��ܟ��i�Ԧ̓�d�K�*X�m �P
��Q��$��%�&��O*��J>�.O��$�On�R�;5p"uJW�Jԡ	�O����O �D�<���i�8� 5�']��'i����V��U�4�c/�01T��T}��'���|��l�T�JbJKD�PŚW�K��䔖��\�v�˗+w1��X���.w�d\1]�D�h0�$.���q 7tRJ�$�O����O��:�'�?�ГRUv����Y95af���J��?	W�i�	"��'Pr�b����5,Xtȥ,�0B��]0%o�
I��I���'!D�Rѳi���Sěf��� �*H#%�aPf�	8��X�������O$�d�OT�$�O(� L��H�;t�y�p�
�L>�
����cU��'������'���Fn�1h�#�6mr��*	k�	��t�	R�)�S�V ���o\7`�<	�)M2iJ�T�;���=R�d����O�a�N>�,OrE�h��y�ޅ"#ŗD���8c��O
���O��O�<A�iX|����'p��12���P(� z�p<p#�'�~6!�ɫ����Ol�D�O����C?[��}���#�D]���_�7�!?u�y�n��7���)y�J�1_`@2��j4�e�qK`�0�	�<�IܟH�	� �ґ��)i�1y�i٫b�� �/ֶ�?��?!$�i�ЈӞO!��r��O8!%FMy�jDbWHLD�ސr�J!�D�O^�4�b`��k{�|�N����-hm]@�Vz�<P	1)��I@��Ty�O���'o�k�$)Wbԁ��	"{A2M�G�A6T���'�8�MK&�۔�?���?-��P�B�@�
��@����8�ٳǟ�p	�O�$1�)҆,
	���i���[~�R��m�Ρ ���A_���*O�	���?�7"���H�����i)�"'r�v�IE�'�r�'er���OX�&�M�b��= HD���Zo,\�%��tV����?yu�i��Op��'�b-�%x���9�G�e��=HC�S}�B�' ��F�i��I%cUN���O�>	$����1i��4k�k�o�6�ϓ���O��d�O����O���|�� Сb�u��m�	<}nq�Q��;}\��(N���'6����'*6=�0Ѩ�mPD��� |�$��G�O�b>=b�	�ئ��7S�@hvǗ,w0�V��{ܬ�fw�R��O�Y�M>�*O~��O6���DZ�w�<�
��3�>�;ci�O����O$�$�<Q��iD�I�'V��'�`��@�ޥE��(v���o��Z�$@}B�'k�|�I�(niv.�>jY�4�7�ª���\�jԢ���,`�Lc>m���O��=a����C�&k�*\め�*�����O��$�O���4�'�?)ӭӴ:j s�텞P�(�SW��?�a�i���S�'�"�z�f�村0dΙ C���u������%sw����h��ߟP��LM�q�u��� rp���ܘ��i0ŋK�.h񻷤2I�L�$���'+R�'["�'�B�'�J�X�T�%�f8K���U�a[����B���?���?	O~��zoQ@۸�-*Ԩ�S�$wV���II�S�'"x��(��R6"%&QB !8��ة�mG�� �a(O��c��6�?�$�(��<)G�[�`��m	/G�0�?I���?y��?�'��$�Ŧi	�-�ɟ�:�)��E�B(�V���V���ڴ��''���?����?�t��g�b �T��:Rl�	��m��h_�P�ٴ���ʷn0Y������А�ħ��`I�m�eP�,#�5OH���O����O�d�O\��H�+gl��bA �H$��=ْ1�C Rj��?!Ľi�z9��'��'�1OĄ�w!J�{��=��̭�>AH�O�d�O���Op��kg�0�	ßHs�߿G�"�"7ǔ�OP������kt�'vL�$�ԗ'&"�'UB�'�I�D��/@^�S�o���F����'{�V�<��4Q�4�����?����)���L	�_C�|��r�F�������O��$(��?�!��/֊e�%�̄3�.8���>v�C�%��Zؾ��|J���O�}�H>�]����3W���adзlP�,����?���?Y�Ş���_��qZ f�_E� �Ud�e��jg���4��I⟔�4��'2���?�W$G9�V���.�"�d3���.�?��ZsT%��4�����*��矢ds,O�x����W�T����xѾ,�P0O˓�?����?i��?������ɿ!鰴�!^tш�F��n
V�>Д'{"�)ͦ�2N!����K,JG���GhJ:q�!�	���&�b>Ց��
Ħ��S�? �yT#ІLƔ�7��;Ԥܱ�8Omơ�)�?�Cm#��<����?��#V1 �׎�7Uo���ЃL��?I���?y�����Yئhg�cyr�'I09�Cگv�J=�S��\D���d�b}��'�қ|�G�;n���$ODfI���"��d����!�I@{1��%��E{���Ţ{K2m Ȟ5pʉ��JZ�E ���O���O��d"ڧ�?	��Y$٦�v����$y��3�?Y��i:\=JS�'nbl���%V[���B^h �F���ȟ4�'H`��նi���&\�80�O^l��F0� K�
� �<��B�d��_y2�'Z��'I�'�""ǑR�Y�b��4k�yc a��_<�	�M�5 R�?����?������v�E�Ẅ�_3��b� �R}꓂?����� �x!ڇ�w��l���̰�"ʂ�p��+Oh��&
��?A$'�D�<�5�˨&��bL�uj���]��?I��?���?�'���֟,���?Q�'�zI15Ȇ�VCe �斸�?�b�i��O���'-B�'#"l�
&��)㇫�8���%�Z�����iG�	�djj5ӂ������M�2ݞl)�j̐"\t�Et���	ޟH��؟����(�zԧ<3m����a�u�V@JK�"�?���?9E�i�b�Z�Ob�
b�Z�Oڍ�c�Z�Z�O �kq��Ӧ<�D�O��4�H5R�njӈ�v����u��>�E�b��*u���D� [�4�$P����4�����OH��D��}+�.�m�Pp�E� ;�����O�˓9P�v`�/Z��'%2S>m�R�:�@G�0)!�e�pg1?�^����ޟ�%��m�D쁔�·5�r�3��7R���Ɇ�_�Y��j��4�V�Z��@N�O.��؈+��aA�M�; �B�� ��O����O`�D�O1�X˓hU��/E�
*pp�$�,hM���v"
F�����'K�n�H��O���C9x4!I� h8��7Fg!A��<��i_N��a�'��X��@�?�#W�4P��Y:h��}S���	;P �|���'%��'<"�'���'��� d�}K�C�],���,nv�ڴ	?���(Op�$!�i�OHylzޑ�3��M��� ��a9������L�)�5e��	��t�hA�L�?;�`|�Ԅ[=5�	�t����FKN�d8��<ͧ�?�b�ۮf�4��ƕ�a�6��W���?���?�����D����B�uy��'��e� ��&f�&]ag�>8G��R���z}"�'
�O�UkL	3��15.]�M����p1i�/�p5�d�c�.�2��<�%@��5F0����_�*8��O���	���	��hF���'��C�	u�=��-� �0� ��'\7��Jָ�d�O,|m�U�Ӽ�`a�7S���EB�g����I��<1���?9�Z����paY~b�ݷ#�:Y�S�o
��JP�>B�y!ٶ�*4@��|2U������ǟ���џ QP��e��
|J,��Zy2$h� ��B��O����O�����5'����T)9��<j3Y@Dq�'dB��i�%b�0��*�.%b�h ��0K�lȢ��L3M��;�@��+�O>Q@H>�)Op ��v�le��dBq6PV�'Ub6m�/���:�t��`΃#<���卓�A�.��Bզ��?	�U���	ǟT�I9�A�CޔZ�f<��]c�޵�C���t:���ֽ�ǃ�`��H~��ABH��`�:.��p�i�9��X���?��"�B�׀��E�f�3�?)��?Ჽi�ΡhΟh�o�U�	8)����0��}XV�V/D�B�'���I���Ӈr�y��/?�;"�fx�C;>W�����x��@�^QP��Ε�����&�ɘ)�p���\&>
6%����1["<	$�i�l���'�B�'���)��v�N.�L��u��1 ��W$��џp��~�)B%�=+*�j��\4=V0¥��<Ub����ʏ*Uة�)O�	���?1�f/�d�U��0�	4�Θ
���G�!����ƶQ]�A��$T(-,���-�*WNhx�I���ڴ��'��ꓕ?y��T�� 8���j�B�Aԩ�?�����!���A~�A�<��'��K(�q8e�k�z�J��	���<ߓ D���ǀ.�x���؞�e8B�i���ؕ�'72�'�P`lz�	����}vm��A�)�z4�4̎П8�Iv�)�??���4�y��j��K�*P1	VhQ<^vdX�/b���aQ`��*��<�*O���ǖb=��T� � �J�'��6-�3%jF�d�O����AQ��8L��5\�)�e!�5 �⟘��O��D�O�O.1q���gf��pF"�	{0��R�ʅz��V �w�{�� ����tmM�r�$�0Q��/	���(D�ȑ��=\H=2uT"I��*c$�ߟ��۴�Ƅ���?)��i��O�Ν�[�t��ĎEu7���t$�?+�D�OX���ON\Ťܔ[}�i�;ҍ_�?�2�� a�b����H�G�@�k1�V'2��'��e�'o.����*QLh�����>�T�O.�m�+v��x�	۟���V�Og���p�S�6���π�]L]��V�\��ޟ�&�b>)�Cb1� :� ���#?o~�H���IQШ�b$�W�,ʓs��EɃB�OH��J>�+O�t��e�o�J�  E:M�U���'or7��P��DI1*�mp#���״�1�X�O����ĦQ�?�Q���I�,��1`�Uѥ�n]x�
ËRsh��!�]�f��RИ&��!�J~2��T�p4�	?"fU ����iM�Γ�?a���?	��?�����O�e9@ �	K�@��$A*�
]q��'��'�6ړO�˓y(���|2���i �)�J�њP���ѽ��'q�Z�0x#��1V�iR�E��'�<��vA�	1��q���Y֦�dS������O��d�ON�dZ4h+
�k�U�,|P�rK�Y��D�O����� ���'5�U>�a�N�C�h��`�<L��X���>?A�Q�������%��'<�4q�ΈMD��QA#Au����IġT�Yv~�O. ����+4�m��%Ц$��e�Q%�=A� k���?����?�Ş��٦}2@,��#������3#j�����ՀH����I��Hsڴ��'Ō��?���-1Z5�)
Eb0���͜�?���\���Ѥ �]~�#ƠF�<)�}�	T36P&PX�A	v6|'���<i+O��D�O���O����O�˧2�D�R�I�4e>��LԌ{���Q�iz�P�&S����X�'p�w[���1�� -c>�5��6q
��'��O1�j�H��D"N��D��	Ơ"��BX��h�$<�D*	:���)Ap�O8ʓ�?���c?��7ƒU�FT8�GZ����I䟬�IJy�of�2HE��OX���OXd��,��D� |(g��\4 �2�%�I��$�O�㟜 �D�=4K9jTmj�MR�<?y�h�"w��
�@����'u����?a!$A!OF�IJ�(!Jr�����?���?���?�����O�T�0Ț�O�V`r��ڈ�P!$��O6Ilڈ)�H�	����4���y���:[ẖ*X�uJ���`j(�y��'���'0��Z������$��>d) �O�*��R�P����6��.{��)A�|R]�T�	ß��	�L�	�tK  �.b	b43��z��Hť�fy�f�p�w��O<���O���:��_/v�$��
�tӸ�����OD���'4��'_ɧ�OM���@E�
%|�	e-+i�)�gfW@f��GS��"��]9��/�D�<�`�K�@U���F�H8xY!U�Ơ�?���?!���?�'��Dڦ�"A�ǟp�@�]"S��X֬��TM8�`��Hr�4��'�L��?��Ӽ�@���>7�D��C�<L�ę䅉#��(Ac�z~"������䧉����(�F�A�,@� ZVpA&L��<����?���?��?I���a݁��R��y�B���D٦l��Ɵ�	�M�B-��|��/ʛv�|"d´DP��˲OnF٣����O>1��?ͧ
�d�葧�Y~2d¤D:Lx�(:q*��&��$�~(@��@?�J>q)O����O�$�O&p#m�K�T,B�bR��xR�'�O���<��i�X���'l��'q�Ӕq-2B�O�	�:����3y��"��ӟL�I`�)2n�)B����QN�~jq�,ƲS������[,��H�-O���Rͮ�J�Fz(���+�#+ʦق�葧 �T��0�вz���{��"&�v���@� }�J�	f�y�"ꚱ�����ݨN�|1:#�<��2g܂Kg$ n�/@��S��� 5[���5$�I�=�^�:B�tzh-B�o]>"�yF�&�nš1G�I�q��Ή\<���hP_�!8t��R�쨁D�,>�ޥ`�B�}{Fњb�Ó,$�}C��O�0�xu�@70�h��Vl@]R���RQ*w"���sĩc�>tqeĊ���.SX� �J�_�ʘ���"f z ��m0h�|���/�7Q�� ֆ����<	�����?���6]��d�2j���L���9�"�����?Q��?�.O����V�|
�˄�g��A�&F�!�Ź�������'�"^���������v8���#�������*��8Q��h>$��O`���O���<�S��㟀�pAS*QC��Z�OF$,�A��MC��䓜?I�W�R=R�{��;)�aY�E�>�И�%f���M+���?+O\��E�@H�D�'g��O�D�8�!�[�=ؖK
�%���t�<��Ov�$Gnq4���'��q{e�7i������
	�(oZzyB��>��6-�O����O��)X}Zc���y��m8�pʓ��V!�q�ݴ�?��l���Fx��IWV�>�9q�ӕyj��E�ƫW�ƅ��6��7-�Oz���O8���u}�[�t
�ƶ01�X����%gx�Q���M�Rcȅ��'��8�D\{��M�3dC(��͐g�":��l��|�I�����f�(��D�<1��~2�$�ҀJ��̬K���Ӧ�M�O>��`٤I��O���'�2	��x��(r��v+Ę�n]�da�7��O�ei�n�@}BV���	p�i����IÙy��Ǉ�g�a�n�>ad�T+���?9���?Q/O��C�̞�
PY�K�*��xö���"�|��'��	۟t$���I۟�iO�;C��5bwOS�J�6]���_�\L�'����ğl�	cyr�ā~�t��M�e�S��,P�+�hֻrr7�<�����?��j��t��'/��U�W�!�l�7K�8�O��D�O����<IeKѭF��ʟ��% ! <H��-��~T�8���!�M+�����?!��N���{""��@��0����{&fXXf����M[���?	*OT�x�E�`�T�'��Or�C���7��9q߰Z�Lk���W�Iӟ��	�B�$��i�IY� <\ʠi@�?�.����ߖM[ �´i�.�����4&L�SߟX����DC��~�{UM�Y ����G.��Q�������rI|�M~nZ	���3��!���1��.wAt7�M�1u�lZ���	П4�S���|j�(J�"�PQ��	B
[X�J4I��y��f�'[�'�ɧ�9O���%Q־�A��H�kx����.��pmZП�	ßTP4�_����|���~�,�P7�x�	_vr9�d#�ɰ6��O>�O�a��yB�'}��'�B�ST��H.�=+��G1����6�g���ę�H��$���%���3�/z��� �� \�h�S�T���?�I>����O��`�g[�0V-R��YR�*��q��|���?�����'b�O ễ��	T���/ɼf�XC��iH�i��y�'f���Xv�Zr���@-oX�cΈ�Q�����ۦu�I�?A����\$d��F�[�U(x�Fɐ,b^�M�u	C-���?9/O��$��`�f˧�?I�j*^CV����#�`L�!�'m���d�O�˓iQ��%��
@@�/���T㝊cVf���vӞ���Oh�G'�`���D�'n�\c4�ȃJ;:,�3׮��Fz�PL<�/O.���O�����tIb_�9���*��w^xI�X���I 1�p��ݟL�'1��]�֝�'��QR�B�&����d�|�@6m�O��X�DxJ|J�͐�1X�3v�>�� u�Ʀ���C@��M[���?�����x�O�L�9&�߃*�\�! ]�,�42��b����O^�D=��?�i�v���Ϛ��`İd\*\�ȉ�i92�'��`@�1��)JJ���k;��#UA�#}��8'm���OZ�'>Q�I���	�Y�p�`���@:�TIX7k�T}�ٴ�?S�/����$�']ɧu�0Y"���Í?�V	�����?Q+O��$�O��d�<�~a$���^�0|f�9��&g�<Ԫ �xR�'�b�|BV��}!RaEp .e���N?o�N��|�v��%�d�O���?��.T7��tN�)PA��r�$_�D�}J�!ӛ�M����?����'��	$j7M��Z#��S.W_�D�iRc�/���֟��I��l�'�h��a��~��Z#B�z&�,���R7�	�{ bç�i��R���I����	�;��|��N�~�5X��7#n&٣���|����'�rT�,7�J�����Oj�d���i8!�+@�
���LT�(�}*��C]}B�'��'�yÙ'�'��џd�b�K�3R�]��Rt+jyV�i��ɞ̈\A�4�?)���?Y��W+�i���5���N��<�&��5%z�uD~Ӥ�$�O���yB�'��IZܧVBq�u �&x��2t��{�pLo�����޴�?y���?���#��	Yy���Y\@���<e8!;`�ӵa>�7�B#��#�D+�����qQf�'�"���fI�H�(�r)��M����?a�=���C�^���'��O0�w��|�`�	S�.<"��i��_��tmi��?a��?wb�j���ĉ
{k&p M���F�'~�iH� �>�(O>���<���C�)T��&�����;��H���Y�!�	�Z���ݟ0�	柈�	ԟؕ'1H8R`hD� }+`S<Q�D8�Õ�~@�����O�ʓ�?����?��\� �e�Mʉ+���s��
�t�Γ�?���?����9O̭����|��J��bd�"�#N%XEj�\⦅�'F�[���	̟�I�0����(/�\q��oF1-i [�@o�d��O����Oz��<�7+ Wn�ԟt��D֟�@]��S�3�KV�|��Im�ǟ�'���'��y�Y>7����p���'J�0cFȠA<��'��T��h�@�����OZ�D��b(:DD@&,t�8qdĕ4<��B�d}��'"��'����O@ʓ�����6���!bŞ=+��	�����MS(O�
�ș�����������?��O��XJ����B�]D�@l�#"d��'1�N���yr��~�ܸO�vd�F$_�L�����Z�Y=BJ�40�s��i��'��O�2���$�5@E\��P��b>�q�s�;�|o��/\p�I����'-����̯X�q���d�-�A�Ȏ+�)oZ�� ����R�`����<����~�Lѣ1�z���=AĨc 
ߛ�McL>�T��<�O��'z�h̔H��Cs읬)މ��$�#�v7��On�p'E{}�^�X�I~y���5C�xl�!�c�ڳj#ʙ���ƀ����d��$�<	��?�����8�LeC�@[�E[�tj$�=e���hA̋v}rU��ISyb�'8B�'�"���
R�R�r��@�'-��sT�V��y�' ��'�2�'��I$����Oj}��?���$�\q
�Cݴ���O���?����?)����<�1R%��`&Y'��e�i!Tb�/�>���?�����d1�*@�O�� ʎ�C�DGvf�G�E�b6m�O�ʓ�?9��?!���<�O�8�`�V9�N�{��_>K�ݩ�j�����O��n3Py�e[?Q��ҟ����Z�N�y4�2) N`�Dc�"\�b��O��$�O���	B��	Fy�ڟ~�)-��K�,=��	�[�i�w�i$�	�/¡)�4�?a��?!�'H��i������B��q�Uh'f�v!�kf�~��O6H�8O`˓�?1����R5����A��yL��	-�M�?I�z�l�۟��Iퟀ�S1���<	��U#v��Y���*o��1a�r�f�ܵ�y��'D��{�'�?�f� �i�tL�M6$Y�b)ƴM/|]�S�i�2�'P�Ɵ8�����D�O<�ɿP��ei��RY���фA#-��7M�O>ʓK����S��'���'��M21CD�vD\,��`ѧnc�a��o�d��ֿ�!�'Y�I����'XZc�҉x�O����6iU+a�)��4�?i��<)-O6�$�O`���<��KߖX$�ɒ�s�8Ce���IdLi��P���'��\���I���	�<c*%S_{B�����}t�#��3?��?����?Y)O�@����|�q��tD6Q��H :����ئ1�'!�_�4��柀���E0OklmI ���1j
���NѲ1�*e��4�?���?����d�,���O�Zc-|}P�x�l�ӮA�&�9��4�?)(O8���O����mV�i>7�߼�҄90��(bT� cCO ����'UU�t�#J�4��	�O����Vl�@ �B1 cD>t,�i�&O�B}�'"r�'<���'��'Y�Iz��0)F�?�X�Xfb��V_�4C�����M#��?����rgR�֝�_����0�|U�TnX��n7��O��
��$�m��'�q�8�Qsa�5/ԕj-��=��� ��i��t�(`�r��OB����'{�I��4a��R�TӵI��_���4c����?�/O��?�I\�h�6��="���z��F�8��4�?����?9��P�db�O������U�R>1U��q��T�RU	nӦ�O��!�8O�S������P���MR��S%*�7P"8� �KF%�M��|���21�x2�'�r�|Zc��P��hߥ4U|�KX��~�q�O�86Onʓ�?)���?�)OH!������[TK�sBVD����<�%���	���'���I��t��B;<����B "L_��R����	]y2�'���'u剥(c���O�Z4��Żw�:��s�W�.��I<�����O����O*	h�7O�q�#V�U�M���ΠDI��I}��'�"�'D�I.AC�uYH|��� �,�r,q�	�. �p�eɟ���'�'��'z���d�* �|��0LW�t"�w�V�'W�S�l��G��ħ�?Y�'�h� �Oc�zi萃��5�2�x��'$�)0=2�|R՟d(fI����3hW9ӔU�i���I��m��4M��S˟�ӈ��DW�"��s`��b�g��0�F�'����yҒ|��)�-~��]��X
B� ���h֚4���hX.k<�6��O"���O2��Z�	ڟ��&�$h`�ms1�X'q��-z3�K��M�`e��<�L>�����' ���cQ(e�L�F۲P
j��
t�X�D�OJ�D�$����>Y���~��_9mP�}�)RWnR��-�M#O>q0ܹZ��O'"�'��IK-L2���C��Q���ƈN���'�����3�$�O��D)���*A��ׄ��2a)ɝ!�H1r1Q�0���u��'�"�'pr�?�#T��M�H��W�b�v8�B�Y�v$��>q����?y�H��x �ׅ[W,ʥf�=g�\��ր�?�-O��d�OH��6�@�Z����Mrz!ku)�X��#�k�ē�?O>I��?����?	`�F6|m���N�YK.<���J�jc�	�����ڟP�'�0�i�)�)_�`�0�tKؐ��1�r��� �mZޟL'�D�	ޟ��ĭ���(�Od�j�JՙD�m1n��2�^���i%�'#�I�!�l�{M|
�����JR]$��2#@ :��
A�K�@�'u�' `x1S�']�'>��ʲ4�4H��	C�/nd��1`�L���V�8!�>�MkY?]���?M�O���k9�h�Ч�)|���2V�̕'�������G;��ꚒB?�e��L�	�M��CJ�c�v�'Xb�'<��" �4���9��zAP���J� vUv�Q/j}��'��O1�@���n��-/j�����yx|nʟ���͟�a.�KybR>U��O?�N	�I�2��&����x�@��r�4�I|���?���% -A�o��X�XW����i��怼��O���O���5}b�;^�$����X��7F���D%N1OZ��O��d�Oz瓰-���3b��< ��u���^�q6`�ȹ<Y���?�����?��'뮡*׎�	�v0C�EѱK�$ݴ+$��'���'ar�'��)�	��i$TؾP�sF-%��M���� Su��Z����s�Iܟ��'Y�y�4~��@r��K�2"az�oE�&�4��'`��'�Y�8�3`F���'#��I���2\F�C���@VY۶�i���'��Oڈ�'��Y���A�e*�t��Ƀ�Ƈ3ߛ��'���'xb"ԍl#�������?Ř�j�<3td�ou2��7�Ӊ�ē�?y)O~����i�Af�ȍ*��S��ؠL֤���wӎ�b]Ha��i)z�'�?���FR��7
�
ْ��Ŝ_�f)j�F�"+6M�OT�Dދv1��}j�"[>e@�	��F	@������.��M���?����$�x�'��K���@eb0�D �̠�� o�JI�)§�?�A�{?�X��l�0"��`ᢎ�jh���'�2�'�hI9�b-�$�O�����ԛ�	Ҫ��Z0���	)�9���=�	c���	̟���&H�ܹ�G�ߐN��Y�$�T�޴�?�w@�D�'/��'�ɧ5�.� :Y�傰�v
iZ�k���dC�Ib1O����O��d�O��B�? L�GY�;�҈���|a ��aߤ���O����O�O������[v�XE朋1�"-u�zuK`Ӑ����,������	QyR
�)W_�SnIx8�����4�"iK!o�*��?	���?��r�����?K{~-��\<NK������Bo�I��$��ɟ���|��!�g��'��4a0�$x�*˳{@nxq��D��"���OF�*�` $�����H	y�̤@�*<!���cNbӶ�D�OZ�?��� g��t�'��ġH(g$.���9�8�q��<K
O����O�����~Rp��*:���f/�pQc%��ٔ'/��s��kӎI�Or�O��n��q�FY�aTY�+1���mZ��,�Ɉt"<I����B�W2Y���Bw��yE����Mp
&4�V�'}R�'��i"���O������Ebz��F�d����v�Y�y��"�S�O�r���l|9bD&M	_  Q���3�07��O��d�OҽH�"�f�Iȟ �IL?��N����wS:XP����L�G�8:��<���?���8y���i��)���i�l�
�i��挸%��Od�d�Od�Ok�ݜw�F��gL:L�6������z�	n2*c���	ϟh��]yr��9� P�L�9(��G(_ a��ܓe �I��%��	��|)P�� {��ٱ��r���,�	$b���	ߟP��ߟHͧD82��� 6�Ma -����rF���v/FU�ߴ��$�Od�OR��<Qq Ʀy�r�Th[(���>��	��b�>!��?�����dQ&Qnl&>M U"�V[���4��<Ь��?�M#���?���CM$��Ob�iӴᅶH|��X��Gj��h��4�?i��?!���6�����?����?��'e����R�E��:`��nG�f�ҵyÞxr�'��+mь"<��~h��T�����4CUE�$~~�oyy��#*t�6��x�T�'I��H(?��ᗟS�5��嚮����A�����I�̑ D2��O��Ic���
^�c5��">0��4%�z=�u�i�R�'~"�OC(O��d�-(|M	��ح&��%3G�ڌGH��nW��"<E���b)L��%h��={$�n&�����r/ʍ�����G�'BF,㦄^�)nt��	�?b�b���1^!�i�a ��_�2$�SGW�:5�MCU��*zHZ��E�"I���?BQ�#��K�b���ER�mr-���7k�����D(��x����Nsv 6-ô.P� �B��	%r�Ku�9w�jKB�C<7�8C��XL�P��Hٸ������ � h�$|��$�Ot��O"��`�O��D{>)c��7/J�щ(n������x��#C�!�J8���H(����$Ҫ";r���U'V�!�6K��Nf	�sNC >�֬(�ϓ֦1X���ceg�09X�S���:c$����t�GaB�#��F��y�X�VnWZ�'oџ�Y��8��*�B�0/ئ5�3
;D�d�E'ՁnNҭsq���aQH����y���O������'Z����p��b���.C��ܮ[�~�;��͉P�����'�R�',| �����X�w���S��E�[�y("n�6j(�j7����dK�`��tH�����}�RH�9A��9˴��)EkI���GQ�'~���?Y���%��^p�o�,L�:D��Ǌ�yb�'fPD�D�*Y(:#��e$��^Љ'5��xWCC�a��lB�mZ�rL��'(���(�>1���iV�1H��d�O���ʓD�X��Ūצe��Q�HOt�|0W���m��.8(,ק�7��O�M3#	�,F�
�9p P�������ڠ�pḦ́J��ѪO?�DO�;=������0�t�#ń���C�O��!?%?�$��2�ùC���Fۡl�v �B�<D�LKƄ�*�>q�pO�thؒ&�.$-���?�&��1�ۣc�TD��É0]r����?i��X��Н ��?����?�������O�iѰD�T��3����x���O�#C�'4�8z�c�Y�搱�aJ�U ���'�x��"`���dW
|����ɍQ����$�R��	B���X�L�X���b��q�,��!�,D������\��r��N ku�|qe�ɵ�HO>��C���M���MY�P�dۙhr�)�n���?��?i��2
z)���?��O/�)���?	`L�(8�N��C�&'�]1u��P8��ٴC�<9P�[<t"�	��6'֜1s&Q8��xsF�O���F^NRv#�	I�dQJ���
�'�B�@���/F	;C��V�H�		�',Z��%�ш:��TQr�ƔZ���R�'m�b���g؛�MC���?a,��0J�;Nly��,у�0��M�9p�����O��N�\�(�|�`�X�4�]嫈16 ���s�''ވҋ��C�(�v�jP%�w�0X�ĮP}�Q���L�O`�}���O/	���Q�έK���qՈ�h�<��Lɏ-j��!�K�2߂д �P�hI<� L��
F�;��{e��!b���4O@�� ^ަe����OJ�X�5�'�b4O�hu@��-��]���_��6�B"I��y"�T>#<)r蚞�l�k�!֨�0��v�"�l)Dy���'��+�䞮2���T%�
���qM �b��'Z�韘"|�	:eJ]s@�	0%:X�Qh�;v�P�������	�E:�4C�A
6+p�0N!�^#<��)���AC����Cؔ9&�yuA��?���-؂��%��?��?Y��8���OT��̕I�fD;G&�s���XT��L���"��}�	 64I��ї �5Z�8l��b���~BȀ���>��"@�|biKA�4� 8c#�Mp?�SK[˟���	�>˴,;�ȵ~*��a,�K�HC�	;g ��qr����1�a��~L�����4ڸ{ڴUU:��JC�cplD��W #���P���?���?1���?y���tdZ�?�<~)��&���
!�2�ܰ(�݆�	D�j��Ȭ���~F}��-JY�D؆�I�*]l�D�O�`��Q�y|֐�k��_(n�ڴ"O�e)"�F=bnH�Uh��&R+&"O�����]�s�R8��H�4u��3O&��>Y!�ҙc�&�'�bX>ݙ 蒥h���h�1����-{t.u���p�	�:��L�	g�S����'`Z$��ڧB(B����(O���Ӧ��ӧ4�z��%����<Y�*�6m>ڧ-](������Q�Ԩ���J^�a�ȓ,�5�� ښ)���A��T�v���-��;���F�X=n
�B�� �ϓG~��iHR�'j��w��%��ΟX�I2iX���c�V8$�I� �a\�e�t�Vٟ��<��O,�ʆ�j�|m�qGkx��ë#zͤ"<E���e���
��%C,\��B���8Y�_��?	�y���'C�-[卼�t	�1�S9Dr�A�'�vt Qj���5H񢚲$�`Ɋ��$�S�����!�����22�ҽ���VH8��D�O怈vhŒt\h���O��d�Oֹ���?�;��t�C��B�@0��j�PM��1������A��@qF�~�N��@��UZ��IfP��Α7�Q"c�L�R�^��Ò 
��d{c2�'��q�$���q�^xz��I
	�~� 
�'Β����R�����a����#�&�S��y�J]&8V�1����7j����y�^�'�D���K�Q�BЁр�#�y���W�<z1.�&4�̈�P�,�y�KԋZx��̟]�yeO˛�y҉E.3�ֽqlB�X(�@z��W��yroP;���٥G�!��I��N��yr�������N�5,��yR�?@��Q�I��}v��D ��y�Q<O�X1�m�q�,(��I��y�Q8^y��.	fJ�x`g��y�6;9�\R�`H�Z0�t���y�!U�(�$$�&"�5&&����і�y" {\	g�E#��x���E�y"N"$0��u���P��*�ɟ3�y�j�� ϜA:B��
r��>J2����W� :�
G�a\)1R��}I����Zú8yª�-3"n�Hr�C���ȓHN`�9�%P&�9X��B���T��x��iJ���ԕ��NU�l�ȓR��%
�u�����Ş�hȓB��-@��O�$���\�Y��ȓS� T�A=$���gO\r��ȓC��2֧�"[�e�X:�V�ȓchL�!����#��H҅G��<����%kPD�`��d{*�	AM#9,���N�xf��N�������Y����R�ƈb�D��RV�L[m�L/�E�ȓ(�pp�D���)8�*�a�"H�R̅�C�f�`�.F�R�woL8M���S�? "�ؔMҝ8h�숁@&�H�"O�
̆�됡ᓪ�3�ԡU"OJ�q�.�r� ,�e)�Yܭ�C"O�t�� ��A�pIՇ-����e"O��{`$ �dx"���>�:��"O�I�'�C)W��Ѐ�*Z&[�&�Xw"O��2��I
��[���4q��"O~4�e+3,H5YR��y�,��"O�1�pNy�b���U(2�ƉБ"O�)����/�V�5�ı���\M�<Y�Ǝ*!�� ��Zс�H�<�rI��XL�w#�(���K��	G�<9��Q�af�+�!^%EV(KƦE�<ɥ�O�m�1�+�`:� ��FQD�<!`i��CS�hG���a���<A@�L�z\R��&MԚS�@P���YT�<�rlɥ+��S%�6f=:�O�<����U��Ň\`	���V�A_�<�0$"����U;�tԱVB�b�<a1ɜ-@��-YU�������_?��j�/k��O�>�b" 	B`ti�7����Q2U*Ox���Y+.��T(@NL���BԖ>�Ѐ��2����L�~�h��A8(�� ��w5�~��\7YJؑH�$[��h�S.K�V�^D��KF�<1��Γ[Nܻ�DS;`��9���'4��%���O`�q�$����a(�>
��N>��(�<�Oq��	�&OV�z�ޡ9�zm�R\�@����1�اH����M"SΝq5�Y�"�Z<�cKOi�K%���L���g�L50a<����N�(S�̠f(4���Ƈ�+]T�[V\)�	�|�\|��җ��?Q�%�"��8��o=+L�QBI ax��po?/D�'beI��>���#��ǩ���'K���D���rڡ�#o�2��T��y�o�0�b�b>�� ��oܩ�磌3�� � D��c�g�H�z��V�W�/���T�9D����E6�=��բ+d� �$*D�`p$\0n<�F׬|���`�($D�(R������,Jk\�C�L#D����y��`�7%G.6J�9�"D���j��'7f9� G�.S%:Y��3D���������B �
%���,D� 	�H�><Ȣ����AJ0q Qe,D��p��8r �;S��!q�Jm�3)D�,��
D�U2��N�6�&��qB!D��*"
N���eQP�_�ibE�bn$D��4c@�<:N4äƞ�:%"��m0D�D��MÝU�P!{2�\�G�t�A0D�8��c�8a���W4�Lu��b1D��HgF�7ޜ�r�.U�`@%���-D����݌Z�Bx2���;f�!�R�*D��s��[�}��B�D�I��q)D�p2��%�fH�#	H�M�%�4D�8��Q92���#*	l��if� D�J�*ՍO,�8Hac��d�t9��<D��ADî<]������lTt���9D�D���߉Z3�)h�ƂPT��B7D���儋q'&E��gL0�l����4D�d�u�	P��u(bK9�bS�b%D���6��4h$���+G��X]���#D���j̥��!C��_XI��?D������+i�0�{v�,�@I<D��K[�������k����e,D����� �zE�av�O�g2�A���(D� qfC�?/�ЃI҈xh�2�F%D�� f3�K�R�ȝw����UH��'������!}«D�4�� ͘3�8G)C)�y%2}�̳��H�x�(�р�0�'F�(@az>m6MY�_��C�bOlFf1�A>D����,<%"�)p�HZ:\�4���"�tZ��<�DH.B�0��s'5Rٔ�R��TM�<�ǀ��9�,�@�T��V1�Qc��xh(����H�� ����6Z1a��ӣ&�Haa��,\O �t��3��$��>�;W�Y�|b6\�B)ՐY�!���^I� �ݮyT���r���qO�eyT���0|"r�T�s<�2F{��3$d��>)�C�	�i��5:����A����Z�4��&︟p5���M�eM"�gy�m��!�,����c�9��N+�y�"1~1����I#bh�CU��--�0��Cڒ�~�^|)���5yRD9A&oH�x`|u:�	�R������J�(��}ZT������ �X� �����	?�>B���T�cP@�8C$�J�	O�f���@��,шy��r�0��� ;�X� s�(��xB�\L��,�4��\I6Uk���@�ܒ�M3� Ք/����?��톈2�|8%�O4-�Ʃk��!O�A�1脐~Q��OtP&F�j2P��椘�=!��3���ڜ��98�4&���B�V�V>n-)r�,�̐�'�Z�����-.0]1�O��\#�螯/6��$�"̘YJU��
��uO����*�${�X���*m�؃ϟ*���ڷ'HTh���>���I�6ޮ�<)�GO,:W��C��~�h���O��|�ī�>}1�Z�0|��m�S�Ʉ1b�)˶B �e ^�۴isZٰF-�)��3�@8�����(�KƵ-�$���-s'@9�񩑴h;�+��K�y*��.�\��\,l�T}�':<ep�oµ69� u�'9
��͓R�άhf
]��3�'i�=+�ܪ&&�D�������~bJH�pd�`M�5w��xeB�"$-��h�W&N�!��|� �� ��y'��PViL�%���'����<	d���T헒
���*�w����獰�*=P�`��	�85��,��G��5I��T}�X��r�N�i��E�'��T`o���l(��?7�R`;)��e�*O��'O�`ؘ8�7��%+Gp�z��	�w
	��/_� X�9�3��k�p���A�5��)T^�a�ԑ	�t=R���
��F��9f_@��C��@F�!��	X��E��zt*}��h�2g�2�d��
�i�C��
�(q��?�<�d�Ӧ:IVi�!e�t'"h��B׽.�<l���'�L�a�ށO��{��-rrj5��Ƅ<�?�P(̼��'�
��	 d��h�5�H�[`
M�xs �J���'�(�v��*k$�,2f�$Jq֙[�&��&����H���f����X�*�H�o��u�����:J���K��E�T1�cP�&Q�"<��,Z:1�;gg�(;�f@����S8Sx�<qEmʇi�R���e��]3���3T�}�r)Aeɪ�Y��U��x��Jp�ӅB��Hc�/	�g��5BS�K�p�(5Zi�V|���~�<��M�0k�9+��ȗ!tF���M�<�0BI$6BT�A��x�p�"N��E�	<jp��w�nx �R��Jg (�;�>�y��)y�T���8HR���%g��@����,'�!��ʢ~��TC�Ē�g���z�c5手c>h��	]��-���Xd�qOJ�z�!�L��z��_�A��� ���3R�V���S�}^4���� 0�I+g�����Z1J�$�K`k�(U��Lyऔ?l���ED6��P��'�ir��[5��񬃍:Z���f�w�t2UKZO:٪���>�b���~:��'��ɣ�-�2�hO�#l��e�<-O�\�:!�K SF
��T#՗/�y�A��sЬV�:�>Dy+O�qd�X�>j���U/~��\%\�0�
��7E,����U������]1G��a�pM\60�@ CR�<���˳�S�J\f-��i2p�E���d��i�{]�A"KB�|P�ȍ{rHӳ<�Fx��!�"C��=�Sn����'���'n�O���ڦL
$��W�]���� צf8�a��W�.���P͎�@�6li�O1���&iʸIU�zr(9�������, ��MD�u������MK	8� 6�{[DuZu
Yh^�����@#.���?�q���1�� 0�#i.b9P�fKK�<i2�=?�#�*^�Yn�ip���f�`�B�ǂ "��%��B�G-\����	!�"N���hr�����ү��
�̡rBMQ�nV��G I\8�DZ�!d��i%E_:1��p��{�h	w�بAr􄱕�L�qkL<I�+;�\�V��.Xv�Q�O���H�䜚O�ў$���*t���U�=;��?�Q0BS�u�����b

�p��i���v�\5[�p���'�&p�u�Y1}c���N����'G��3��lP���5H�*&q&>�Cc��S�m��� �	��_lfٱ$�ϨBDb5�B"O�H�¯B7r%:E{��w���{�m��n|*u!۴(�0����1���R�^�j�Z�'kxͻ}M�k�:u����d��$�Lx���)/{>1�d��9X��J2"Bc� %���Ԅm&���M_�`�2�sN<�%���FE�O~n��bM�S��l��a�ԥ���?�1%^���D��C��t�'Zܢ)��C�>[(�e dhn@�ȓNS���̈́���ո&���4�$p�OF��uEV)s�H��a:�';���j���0 �X�(�C6�a�ȓ-Y���ҍ�;����� O.���ڎ}��W	<<��S3��-]ily�ԢLu�8�ȓ#��	�򃒐P900C��q�20��	3�<���ޫc:��X��˗^X4��ȓ ����eL�z	���*ʒK�N��Q��Pc$�Ӡelr̛��;�� ��T&6�� ���tǢ<��Eh�R���k�.܉f̜�JuV�2�Ȍ�nLN��ȓ|l�չ㎄7���F&�L����8bl��F��%נ��"��u���;e�9:�Ng�sc"R<o����(D����Ny�M(2�K?&@)h1m;D�,�EkK�Ш@@�K�.��7�:D���U�4��lBC�&t?�b�6D�H㦈�����f	�9\����5D�8J��Y�d�<��̙�KM)�6b.D�4�jГ=�xq�dإy�L�a��+D�`�Ј�f� t��
m��3+D�PK�N�lZxD��A؟{��d�# +D��"�AS�y�Tu%U�X��y�+,D��	� �")`���7q��)�%D�$0�lG	B��5h��Z�1L�LX'D�p�*ֶ@?t$ᢊ� �nB5#D�8)�'0\��D��N�@�� D������mWޙj4���3:\@b"�*D��@Aa�>D�<�QK;j(��H+D�p�CĈ�+^p�`��'.��; �6D�HU�E�W5��ʄ!Hq�~����?D��	�aY�����l�"�p[`*D��+�g����AC�&�>0HV�-D�(z�sƲ��Lۅv9�еn?D��Z���i������8I�T!1D�T�d/١L PU� �~�b�-D���'e-��dE�p� �C�.D�($��7,E+W� pXԩ�e7D��CƠ��>����]5L��u�Q+D�� 0�܈0#Rx)�Ϝ�V��a��>D�$�w�܊!�����k�Tp���7D�X���gN��d���3�*-�`n1D� sd`��<8�Ń:?�.�r�0D�CȈIb�8A�C�p̩�:D�<;���g7�, ��J��ak#/=D��IQ�ڈ5��m�r+/=ЈI��%D��z7�R�[��dc���=<"Y�1D��볨)�j�Y>��Ir;D�Pj�l�"i��&�0N/.����-D��B��^9n�
�`U�[� ' &D�3g�@�&,�b��6����R�/D�x#�a߃z��:ł����#D���Q�R�o,��QE�9�|h�d�?D�L��	� ���ъ��V!F\?D��PG�Q��!�Є 7Tlr ?D�t�n[�A 2�� �6Q[L��L;D�H�T+��A��ĩڪl�$ZB:D�Ԙ�U��%���ܫuV28q��8D�(Q&&� v4(�4�9V��1��;D�� q�Ӥךe�� ʃ�'�r1A"O|���`�� 
 �CB/�|���"O��+$�2f�Dų�.�'!���*s"O^�i ��>0�L���Ɂ�Y�"O:=9DeJ0B�)�NE�,��"O�3U�MzE����k[!!G�h&"Oh=p�G��~־#�+�990B�"O�1s� E�!�Ƥې��U�J� s"O|PH�g˂����BaU6e�N�+�"O
�8��Z�P�b��R%����r"O�� �J�X��6��"���ۇ�~���i]�Mj�����:@� a�D	�!�D�"��ű0/�4��|�%�e�!�%\���1&b&Rw 5���+q�!�$��t�4�����fe�맄C��!�$��C�:py6H\�Dd&awa�D�!���|hnu�t F�QS�t���� �!��I�y�ڍ�0힄)H�{0�!�D���l��EF������!�DL�(�Z�0�ŏ=���JV��Kr!���n$��W�pἑ)4؋fp!��@��h��Μ�6�`m��m�&T!�d�;v��`I�>8����L5OH!�$P�0Ь9E�?ZH�h��F!�C�OD��u�3g������}�!��8gGP�y�F(t��ȴ㜓:X�'�ۓ �ĥѕ�$m���� -ʖ`f4��ɇ0=��o�D "�P�BM�G��1���ԻzĂB䉽C��8��D4��iT�d��B�	a�x�xv�_*�=A�A׶,VB�&x �BщGa�X-�/�4^ZB�I(_vR��b'Ko?V�Q��C�I,lɊX�p`� Ju�v�\�
��B�I,G�t�`PF &x�`��PK���&B�	�#)�@%F�o��g,�*�C�	:]#�K$��EL�r@n�6=
�C�Ɋ�t����[$��)4ň :a�C�
�h�`R�@�v�|���ٙ-:��L؟�Y�g�0A |����(D��i0D�d���)
J-qe�Z���4�0D���AL�&�Mh���h��4���.D�ӱ��5
6A����
HJ5�� "D�<�Vf�I�,|�jP�Fc&i�a!D����Ē�"�Z$��m�:lq��sQ D���4�X��9�S`�O�8s��1D�㇣Sr�,� 2��N������2D�pq2m�<�$i�S��\�����.D�lr�.�N��=�M�2���{ �)D�\҂ř?'D�{��(�ȴ��%D��Q��B71����BK	�X��#D�@��C�5K���K��T]b%�#D�xjd�;�y1M[2"m���=D�$@��ޢ`��+�+�/��꒎.D�8��Ĥ5?\P�g�),Ę貅n2D����˅�2�X8��!e:�x#�g%D�,K�פ)��cĊ�U�Хp�&D��A��^����u�M/0l^*�)D��PV�s`�!wn
"<u��R��'D��@�nΞ+�X����R�2q@�+;D�L� kX0
�>�*�m�	C���.D�\�Àd��h�6�~��Ï)D���eD�+6�d)aʁ6G�^	�6K"D��e�!&��0�2E�:~F9!��*D�Ђ�
[�=d�۲
F�8�!%D�� ^�yF�h�֐y/�5;�2�0�"O a4�sȴ�GHQ�}��ՓP"O&��Pr)�NL�Oz����"O�I���7_�p��$�6`r!��"O���5#�ǂQj4%^�91���"Ojle��)�"��qC�'��A"Oj�#��:.ʝ	b�~�"}�&"O���cN�;R ��D2";�1�u"OJ)���4��X�蔑!B��À"O�A!b(<<͚�!]	1���V"OrxX��.v<|��˝RN~��E
O�6��G�h����:�C�n�&H<!�Q�VȊ�I�&��o��Z�́$g8!���!5:Lؑ ��6,&�\"�!�d��y�I��'4x,ҥ@�$�5:�!��C �`�/حm���m�^�!�D֖r#�d��+ӘF]Sa��!�!���_E���(T7G~�if�Kq!�Y�N,�GEL�Gעx
�Я|7!�D߬=/L@YƁ�*
�:�`���v�!�Č�k����@�Fm������P�t�!�Ϥ�d1��3͚Mp�g�Y�!�D�9C����&\�9�~��f�A�-!��!p���d_A.��aÔ;v !���j���s�E6��i+ra^r�!��ƿ�2�Sol�J��f�!�T� �	a fڮK�I�G��n!�Y2(�e���KN�+]�jh!���<��-!k
�~�Ӳ�'Y>!�d�r�ԉY�H��`�@��=!�d�.$��aY�v����2�)H�!�d�%D2 ������y��'OG!�d�++{�\�A�8�j�7�(r<!�dX 3���rn�rm�R�55!�Ā1r��{Q�^�ZTe�`��<;!�D<f��YӴ�;@R�	���i2!�X�n��xp7gؚq����i�!�$E9���&")�2Ec��R�.|!�D"2� QD��~b`�`l�3�!�䊹d��A��AI= |x�X嬟�]�!�$�$Lo�{��Z2u@�a�]!v�!���<NF��.��?����$�4)!��@<��d���Z�k�°15��T�!�ĄO��Q1qFڀ5��B 'M�e�!�Bk^=p��"�fR�%�*!�d��7�vUI�$Ⱦ@�rI�pgpL!��
}�����(d���T�1V:!�$�*jh��QC�]�l�3�K�B!�D2cX���B���A��a{��=!�$���H�	�-u�Ѝڥ�G.7!�M�9pȐZE	�ʉ����-!�:@��l��I�+%kLd���D =!�$��M��ݛ1)��u{���%��":!�䟋f����#CW�o>Ekc%Ga9!�5<�6��GEF�c�PD�daM�*!��րn�����c�2�59�'І�V���\N���d���,N�j	�'b`Ѯw�<i�,�N��z�#D�(��Mȥp��):�]�S(.D��Q%��.y��I��xղeBf�,D����ϣ\�,�y 'Z�`��)��*D���p&�X�z� �Wx����>D���1` �S�%�1(>r��e:�e)D��Ԣ�2�z�ig &~6�C�"D�� �X��߂�
��N3U�0��g"O��
��Y�?K������B��R"Ol��e��ov��b�P�����f"O��R`ʡN���1�%9l�hKD"O��31�Z`A1C��ig>�B�"O�yǤ�+�.X@�虢eV���B"OX�qE-��hn2�0�h�H3�0��"O���C��-ش�k�瞴w���t"O�0��Hl� ;�#5�6I��"O��Y�A�4�����S�3A�"O��� �Q�8��c�AA�[^�5��"O$��E�c6���:!��j"O�L���O|^,��CA�<Q:���U"O�` �I�79�pY����o�L�w"O��#LE6P����1�>O����"O��+��U�
��EAc��n��E�v"ONlѳ�;ռe�@A-u���U"O���$�B�A�88��#ʉs""OL�q�NB��d(�iZv����""ON��� =�ţ��6e���)�"O�P�玘
FPp����C��&"O���6쒞i{5�ۙ!1�PZv"OL�ٖ":N�>Iڒ�3/�BX�R"O�`:�o�$
�`cl�,l��@�"OpE���˶q�<��[%����"O�\3v�קI���Ф  2[�
%`g"O��A��ʰ=�(�`'��kb��)C"O�e؀GO�!�ܓ��:��ԣ�"Ol��¢�^���IȦU9�Ɉ�"OX�"P��B;��bH�22�Q"OZ�� F��mY�'	��+c�%�y��DdV��6$'rm�U���y��ثҬi("�"�	�u썟�y�d�6&B����֢G�zm�$ϊ��y�J�\��e�qf�hO`�K�
��yB��fb 9b#ě�[P	��n\(�y��&`SȬ���Y4is�_��yr���R����J״�3$ɋ��y�X$b}&�P����w�x��c1���P,Q�4��+��(���ȓWb8&�*��b��.�L��U�ZK�<����B4�X�G Bp�������H�<�&�?���i%n�5-K�(���KG�<��Ӄq*\��3ȋ0w�h�##��A�<�戝;r�IQ%Ñ9�,�s���T�<ф�Lv�R��W&�6k~4C�R�<9��C�ܔ(v�3� ͘r�<��J�`䝛�'պl*�"�ET�<9 ��[ֈPA$LH�"�>��š\x�<�0%�e�=PK-B�Buzf�m�<1 �S�}e�B�Оe�YZ�A�<y�/9+�`��5-ZjU2�)��Q�<� P�����OT�,DanKb�<)�E�&[�,B��Y�[Q��  �AD�<���)I>�U��N�})��hǀ�X�<9%灺<�J�K�f�8E�i�Ԯ�Q�<�pg�;>�:�#�].�a��"�O�<i�C�P��� ϫc���@NT�<y���%X�QC�2#�6�;s�J�<�+V�J	�� (x��S��TF�<Y�n��6��2,#p� �G(SE�<�5aKJ�Rp�"���>��d��c�K�<�Mh�ph@���	k�2X;���C�<ɲ@�������]�9+֯G�<� �����:5��S��%y�(=��"O����k�1 ��-XW���0�¡"O4=���E�0ݑBg�8�$"O�Bv�U:4r�`rU�K6��X�"O�Mp7 � �<	C���]��)��"O� C��� W�tt9��W'T��"O�ȫ��Y%h �R ��,�Zظ6"OL��ǵUXTI2\�!�~�:�"OށraQ+(>����K-���F"OĨ�砙�e~x2�$Zz�x�3 "O�]�U$Y��
M*@�,��c6"O��Ҡ�	�t|������ƨa�"O"�X��\K�z̈� �7�8	�"O$�&���N"1ROK�l�v%�V"O�<�Ӎ�(YK�5=tr]aqJ^��y�@���찥��3���4�y�F��xa��D�<)�P��R����y����mĦ���iL� ��{���<�y�㈍Q���A��_�&����-�y"O��'��ѣ�$��*���/�y�c�*n@*�K`l�1���be´�y�!
���<��ʗ�ʎ)��,���yB�L�S��Av��"!��4��6�y�-	�=�K��V��{��y��#. 訳�&%B�[׫߃�y2�K��Rc��8Zf��˷���y���J����F]�Bq���'W;�yB� w������R�$!�s��y���)���Y�M5QL�s�n��y2(O[�ލ9Tc��2���R�R�y�b˴a�ʙ�'*��@w4�;G�˜�y�
1�Lb6�J�:����Va�<�yB@�<w=\b��3����쒗�yr`ĘHH�ñ�/E�顥L��y�� ]�d�օΐ#�hm�U*L'�y�oS�x��5���^j��7�y�o�*�:�B�ݰ!��j�b���yiӏM	$)�
[�QP�����y2��h 
l��G{�	�2B�7�y"$�0�"�J���m�����O��y"���T[�)���[�l���PG	�yBfƙ���x�A
*T,�� ��y�G�+n�M�k�b�F+�jV<�y"!S`���X��T"_"�X�F�yB&8#"4��b��
�N�/g��Ņ�1�f�Zƭ9y��܁$�H�A�v���~Ԓ���:��`	�ş�God��A��;�W�B��1�̯7�����z��V�ۭh@\���.j����)�����P3��b�
֎c-�$�ȓ��T����`� �����x.��
]8��`GJB=0��&͢M�ȓ[y�)I����:K�5���85&Ą�Y<�-��������WN-}U��2���a�(X�����N����:��ۥAɉJ�N��O΢�(��k`n�i�#UF��@g"���GRzزS��I�^�8�+��s���ȓ������,!��RT���@�08�ȓ�j�"����@�ɱC�N�P��X��)�D ���61*VQA&��A��ȓ}{�M	g.O�Q��(�ͅ ~�i�ȓD�@S��	:C>�uo��r�ȓ^S�9P#װ(�N�H�� �t�h1��S�? �a82Z#]�lХ�K����	"ONm�q��9ɼY���P".����"O�Њ�ec���#J�/H6Hmؕ"O����:neA���*�8�W"O8 �7ÄY�I�j�4$�Щ""O�	�E@�K�|��G�8Y��"O����ǮS���Av�͒3s����"O$��#G5R��Q��^!`�`Z"O�YE�##������&RQ���3"O �[�CU�^���4�υ17fТ""O$��mZ�i�&M���)r�D���"O�1MU��m���jw8Y9F"O����#ݏT|��/��R��驡"O
<JƨʓQ�z�:���,!=@A"Od��#�Z4��C7�!,�;�"O��MȦq��9��ARJ��h�"O:�(�	�R|�y�f�!|�4�z6"O�����!�0=��œ?�`D3s"O�D۱��?Kapi��σ��|8�r"O�ea��R�6N�٪b��vc�]i�"O�̡�1&"�
���t�s�"O����$	�jJ&h���L2��4	�"O|9Z��MQl��jֆq͖P�W"O4�Y�� ��|������ȑ "O� ��#��*/�L��̫PRԤ��"O��"��
\�uZ&d�>���D"O�mcDHR�͙��׼`�Ę[""O`��4�ΞI���Sa�&��<Y3"O� ��˙qb��@ŕZ4�E*�"O��W�Ԏ� ��b��1V�8a"O�|T�D�
�UĀ� 6����"O$��Ө�2d��i�A�-��x�"O�U"@�;|�R�P�Ȃz���#"O�9k��\�vl~�(%�iah��"On�3��@�n"6�Dk4�\ڴ"Oع��l%5U�Mk��..=���&�I}�O�͊R#^Ŋ�C�a(CH���+O���$ ����b���UﬠU	�*9[!�dT�0QVY�3k�[/��01�MU�!�d�)}+fD�t؇+�!@�R��O>��F+�8�
%B��Ձs���""O��Siѳ`~��k��!Z���"OF��D�֤:�q@s-�#Z=��r�"O�r�"�H�(���k�Z6��c��'��D��H� �xИ��	?"�8�PI'D��b�`@T4@0t�̑��{��"D�`�c�س8L����E}�M�3D�0"��ݺJ�8`j�(IoR�k�I1D�\��N 
l���$��L�5{F@,D�<)veX��u��ŗ1+v�-%��&�Sܧ/��#�!�2��(��F?��1�ȓ(�|DҔ�ݙt� ѦЃѢ>D��x֭G@��qW/��h�x!p>D�t�檔Q,��ht
��E�f�y��;D�|�b��3X"��`B�c�V�YŦ;D� 9dFȆ]�0�S��1X�T��uD/D�H����gԶ��h�=;m�Q�<Q�%@^����μM� �3�Ny�N����QyR+� �[�H҄FL:\�U+L�
!�?=�a��oAS/ԉg���!�$���I3��O["Мز2T �'2ў�>�"��D���3C�������8D��p�F�1[0Ja�Ǣۀ:��5�5D��DX�FBz����1=Ԓ�­<q���3� �i���O� ��1�$��7Ê�Ö"O��w��dpp���L���"O�����**�y�unƖH�����'��I�<���	B� ���DU�� �N�<ÀB�p��x�gʇ-���"4�N�<ٳđ;�|�� �C�,n��jQ��M�<�tgM?p��@(�+��T��a
�'�G�<a1b��A�b�(�X7Cl$Ԩ��x�'�ax"�؝g&��D� c��EX�!W�hO���	��z�l��kH�W�~�Kg�̔��=)�yB��'���ctƅ�T�"�-�yRj�*em�ؙRm�6/+�a 2�� �y2#e-n�	Vu�X����y"CУ�
	0f��P�અ��y򏗞-v"`k� �6@͒�Isf��?A
�'���Z싫8mҐ�ጅ�f\;.O���hO�J�aJ6kQ-��!�ŀ�6�<%��Fz}��nH�zc %p�߹;�Q��,��(�Vƕ�r���I�bӲU։�ȓ0F��p��,���b��}��H�ȓ\���� �Z�)��ӡ��}��8r44���?Z��yԮ�G[P	�'�ў�|�F���j�C�$_�'IҹI�
m��@Γ:Q��� �s��8�T쒦6�Ox�Y>��F������e�*LtȄȓphaZ�F'=F�Cq��*�ʡ��w���k6hѕ6?:�J�PB�܆ȓ:D��	�I�N2v�(�ڔ's��F{��'XV��Aɧw-D�Xp',&���'�N<s��V�2:V���n�uV��R�'��#�"-��Qh��@��f�K�' ����/����Ԯ�>l8 D0.O��=E�d*�[���J�t�kH�yF��y��bmE�WU��b�]��y"�	k�P�o�f;Π(��P����?1ӓ4Q��!B�/~��j1�	q܆1�ȓdh�	RU��P����ahJy����9��#�M�,�e�&��ȓW><�H�g�<��d�fj�848���ȓ�.��.ǤT�j�:K�_ӈ���'��ɄC�#c��|�&韵X��9��#~��v�UU�8�pG�&����	l�'q`HQ��*	 ��C�Q.�Nx��'+��gi	���#���qF�X����ɔO:��"EƸ �+�K��v�q�'&����g���y����V:���x��x����,
�	^��Ɓ2�yBh�v�>��� |b|�@��W��y����Qj����O�k�L�d�0����d �S��% ��1!W9���8��D�<�ުOM����@�N�i��k�A�',ax"��<Ў)��ʑ!��#�"��y"/�b�NU��-*��6����y"�]W�ap0�T�f��M1zC!�K-Nu0d��|�b��'��J!��׎���0m�W������ZI!�^�ԉ�c��	Z�*��Z=i��O��=!�OX�0��C��X�1�W8*���"O�tx��5rc�U�V♣d���E"O�i:�*�c���BU/p�P�W"O`�`�E 8Cjp��W�y�.��"O.i;�\�	�L���9䎌�"O&�)f�V$�X:��&a�R%R�"O�e���%rd�:f	�GmF(�1�'W�)� R�j ��fM�أCנRZ"!r��q�����1w�`�Y"�X�c0�D��B)D��)�¢�.Tx�'T'q���ū&D�(C�J�H��@c��v*d4A@�0D��i碏7d�XCκW�!�� ;D�Q3�A8fkz���f%����,7D�l���O�D�"y�dÃ9��Y	�C?D���u��
`�Je�3-ƊA���ȳh=D� �F�'Rą2F�s׌AC�1D��1eD�4��6�C�/ʞ��&�!D�$�TC�K��H�#@�mZ��#c D�ȓ!��?�l)�so��h-�sb3D��hCKܻbilm@ �Y�X�P!�ׂ$D�$
�5V��	��MY�9d&����!4�x�c�/`n]���%�@��3�ZA�<q��}���3��"zB,�a	 V�<Yɝ�8�TD���ˈ*�tcsJWO�<H�7���$X� ����LN�<�Rl��J�l�×�P%B0i���OK�<iG靮MI.��%�'xW����/�ß(�?���I43I�I0Z�Pi�3�ѣ��C�I�N.\x�� ��-� )��� ��C�	:Y��pG[*>�>}�PGW����7�e����߽\�"�'Ѯ��ȓ^��=���J,�$��P.�l��7` BVf]�I����$/H?�����o,��I�N�H8}���OQ<��8{���6
ڱM�P eK4$��ņȓƀ)���Sgi�b'�`.�	�'a~bJ��O�5sP̍Xj漰���yr/�Y��E"�	���z�Ď�y���;(�����|�4�����y"�^.��`���rI@}��6D��y +�0��5	��(�8�5D���'��1��-�$�
m��1|ODb���w$��9�\�#��n��B�"D��c!��:�����f:>�� )�b�O�=E���T�h�Niz��M5x���a��B�!�!�a� �	o�E���	�;�!��V�ڒNQ�X�tQ�o>�!��Lm�xe���	m��R����d�!�drǐ��7`Q Q$*8w�G?h�!��LZЀ��g��-��7�-7o�O����
���fɿ7Al�k!u��ͳ#"O���ө���j��P��(���"O29YWh�E~�	�H�%K6)"G"OL���E�q^EI��^�}X� �"OR�@���Z�VA�e٢+*�"O��A���)\,�E��f?}�+�%�y��U�*ӆ����* �M��Ό=�yT�.�p���A�l[v�S��y2���sg� ����"ar�H�H���yr	W�u���ja�F�p$\`b�K	��y�؀)l�#�g�։�f��y"��YJ�Iȇ���v:>�x�'��y"dY}[qO�2F� �E��)��x�%͟�8%
��՗:҄ЊP)�<!�̪P,ȶ.CB��Ũ�rџ<�	xy��?���C�^��xH6!�-��)�E�=D���vD�~#Z��0cS�`
��4�>D�h�UHT�T
��.Q�Fy��FZ7�!�d�.~�-�����@ 9�@��(k�!��<c�>��g�d<\�B�@ܐv�!�d��r;A��њa!"�30ꒋP����7�g?� ��ꖤ�-x�v��f�2l8�	��"OD\8��K�BH���/,�01"OL�S�INC�X	���H/� �٤"O���A%~��!I&&��IR"O��H�Jč&� %!2�Ƕ4˸�h"O8�!"
jA�WDך*��7"OJ�0���K��,���ݐ%�iY1"O��i�Q�2I����F��>��g"O�|sP�
:e�X�p�Q�Ot��Z"O�-C���`��Ȑ���9g49��"OT�ӠM���|�* R�8�G"O�+�".Y\�E Qo��4��"O��X6O��`W���Eѥ��y)�"O� D�X���C�B
6��f�'m!��K�c��j�@)wȮy V/�!�$��O2����A׈W4��խ
�!��;N���τ�Q,&� K�r�!�$J'?�x��E֥:�(S��
y!��=e���Q���r��ԋ�ٜnY!��[��\H&��|����� yU!��
X���&GƸX�0���ꞛHG!�dV�Pՠ�!��[<8�*���)=!�Ò"x���%$G�	(ҧ&V!�L���U�"�//ʁ%E[-F6!�L.W^�� @�
�f5
�F�>"!�D764���ea�1r߰!���!!򤋆V"�p:��Ɗ��P���_��D�^����7��*�Հ6�V,��C�	7wJݠBIܑU\UA ʽ;����:rk�T���`�F@
�T53оɅȓ|n��������n>f`�Hp�'��Y�tS<M�H�#$C1`jd��'-� ���_���e�q�1��̃�''��(4�3���I�k��l!
�'�m�����V`��:�Ȏf��p���hO?A�#��E@����"�j͒7��k�'�a�4IZ�((`�yV�YŎ��y��A���Jd��;h�$��J)�y��7g	N݊��W�r�X��u

=�y2 ��?�R�S�b��d�Ԑ
���y��Z����`�� `���E��yM�3}8t"��$ǲ ��U��hOf�?!�+��*�<uZ!m�6tZ����F��=1�y�c��^����,�n��A����y���U2dx�'R�a��1�qkV�y�%�2Nƍ���O�F�8��GD��y��!;���c +�*<0���y2�Aoi
�Xd��'8NlaGH$�yBÅ�|f.�`"/Q��D�v� ��D,�S�OS���K�I?ju��B��`N��N>Ɉ����k�H��GD9J�lc�ɟ{�!�dD�x��ULNCk���hI�y�!�����`�ǯA#6_��Q��*�!򄆉w�xH	�N�Rf��I ���!��)�
�i��)AH.8RA�ͷp*!�;|����R8��2�N0F0!�RZ����Ѐəu�ؙlJ�d�Dʓ�hOQ>q�0)�>!3\�2��y.zp
�!.D�Đ�ǚ;���^2�Y��Oέk!�dĚ(�@�C䗕(�~A��m�2o3!�P�4���P*�D8P#*O�:2!��U!{c��; !�[L�$�Z!�CgO̍�g��iL0�ї�_�!򤒯#O����ɍ�aЁQ!eD�\�!�� ��y�Jw(���W4l���"O���duP��g��o��3"Op��֢{'l1"�C75OV��"O�Q3"d��&��-
��ɸKB�@"O�P�bn�3�kď�LNY�"O�E+6�{+���OH9ьtp_�$E{����3h�$��v��R�T���A�e�!��hL(�SBZXX�!�q[]!�d�>8�}���٬&Tf�:v��CT!��h�>���y9���3!�.J4!�DU�S ,�gЩA}z a�OM�!�dV�\�P��E\5 a<$phW�%~!�*4��x�F�!.%�(�%@��=y�{��$�'
LI�[=�\,
%m�7F��}R��h�h��J�4x��A�\�ru��6D����Ρ,�����-'H�y�j D����i
y>B��e��6؊с#D��n��%S���%���G�C䉉d<<��i+.���A ��C�>D��a��tP�Ag�2�tC��/l�LX�5.��9�Bt!@VUO�D%��o�O��DLGޠ�a@�zPI@ש,w�!�䙻>[NysT
֭dd5�Xr�B�'�N��	�f���b�:L���9�'瘠a�C?^��a2cD�?F�6 �'E��A�ځ�����*�p�z}z
�'oR���& 0e�䳅A��;6��	���?Av�ݵ+d����"B�U*�pȲ@��y�eю^�÷�7@����A�ע�y�U�܅#t!=��%�Р��y©��7��p���-�4pw�!�y"�%�*e��HĘ+%T\{��I��y��H�(�(�f�R!)���"�ye�l���`,�}u�yࠟ �yb6�
 	v��	�e�'�(�y���
��`ܐ+*`�%]9�y���2�4P!�<?��Z�h��y��J244�A�߼��	��8�y2�@�L���p��3�>l�U���Pyr�`Ć��Ab��T�dEC��M�<Q�\�2 (�ۻ&�#6��M�<	��Eo��X00#^�y�䔺�� F�<�ĬA(� �q/��r� ��u̇V�<I��_�A��1 ��B�l�8�fV�<�s�L�(e;�JC���P��U�<����8YϢ�RpB��v�}�1-y�<�w��-�B9��#��v�r��cny�<Y���ԅ�a,P�.#�QY��r��t���O��=����J���ĕ?q�d�
�'�NѸ�"���6�RFeF�lX
�'X�����<vB��"�ƉH��	�'w� 9�KZ�W���0�!:�֩K�'�4:�$�D܍#��1���a
�'��hkbAGbʸt���	�'��8B�'��8�b �H 0Y@��H��T�O>��G�y����06�2�����@(^%�?!���~�2I�9W�=��âx�B! �*G�<�3+&b��ʴ��� �+��K�<�cC|WN\�#mU@�wB�]�<��@�D�1{� ��,R#�[�<q2mP�[3��".�':��	�J]px�PEx�`���r1��G#M�J�V�X!�y�X��,D*5�A%R��Ik�.�yb�̀���;AeIBFj`���.�y
� @,cF��A��lv`��b	���"O4e��	E@q�)+����V�x�"O���<��!JPh J(�mjd�Id�4�㮞0+WXɫ0�A�ut���#D��Ӏ��8&�$�*��ۜlb�9�$)"D�t�AH�7�,�3A#�}�0�!�$)�S�'>�"��T�һ?Ӝ+��µ{؄Y��;���GԻn��	˰ʄ�<**�����MS�l�M8$�R��Y@)��S�C���8J@Pa�b0��ȓ��C�lZ�7+je8Q�;Nu�I�ȓO�j�ߡ&'���Uf�7n{�1�ȓ=c.|��D�%h��
`e�)4c��ȓ��P��t��FeX%
�$h��R�M �K�=qȨdq߼!��)�ȓiN04p� �:UXN@�⍙8<�T4��T&d(�0#X̶,��%�4a���F{��'��D��)
�]�'e��f�����'
�<�c H�P�������@�x�'RP-`�'<Ŝ�����[�Vɛ�'��@��nմ0�� K�i�0hJ
�'��`ca�A7<Mr���.b�����'��H���V�)z�e�b\�^EQ�'
�q'Q�D����Q�֒_K�#�'��h�f����@ �M�^,ta �'�ޤ�V�C�?a~(y1눈@:&	(ߓ��'0�1%�i��ѱ0�+
�p��'\�ukW'�d��� �&ny��'���΢Pt𥱆'�����'I��S`�A,�<����:d�Ƶ�'7����
� Q%�Ģ��	/������3�-@�T�#�0gR�ʥ�B�k4,�ȓA�H5#ɩz�*�b��e����D0�!a�"�~=���L26��<�ȓd�`[�N� Y
��R| %E{��'��0����.tF�j�h�hP=	�'��aa�J��B=0�R�M@~,a3�'��r�:ut�i��~���-O�ʓ��S�O�B��C��<�p���//v��9��'\��S��E�c1�9�%-T�fS<���'�t�BT�p؁��[�kј�"�'o��I��I"��A]8r�6aq
�'U2��g)�('�2�3O*�24:
�'+�p���ƺ=���I�o�%��:	�'�n���L�+H8	�ѩy� �'�R�:$�
,�����9_xx�'�:Q0�∡!Ch�a������
�'��u�3��u�|sEPw2$�c
�'�|Pj��,�������"�DajH>Y����1�%�ԕ`#��ae�� ���	�'RZ�C@M3V!�����.�j	�'Pq��I lJћ�G��d Եe"On��3��!#��@�0��
-�P�6"OD KW�G�B��i6��"g�-(S"O�,22J�*p�ZA�
��>�l��"O�Q	�ҸEa��J�	��&!h�'F�'��)�3}�'C5g�Y��:n�&��u���y�lG�*�fK0C�8Sp6d�uG�y�g�
��Tр�6L\l�@D�T��y��Vc�$TC	��a�@c!�y"��Hbyy��= ޱ��*�1�yR(%� �pE�	0zr|a:vdZ�yYh�)���qiU{E��6�?A���4DH���E3a�Ba�
¨.��T��S�? lu�V/�#:\5�6��Jn���#"OU�QL�&���q��.tc�D�F�'��'f�)�3}��9�l9���џ��LB�yb h3ȋ����.�3CB,�y/��B�jH�
H
x���7 ��y��)|q4X��n��k'�Z(�?	���>C�X(���4x��/ɌD��t��IPV)W4F�� �v��7q$�ȓl
�w�_��v%��jW�T~Ņ�9�H�%"p�ܐCcF�!V(�y�ȓ#�t�3�j��;�$R#x�����j(1���F�&j�U
Fgќ֒Y�ȓo,���#�	"�X1�T4`Ą�L	�E��A�r�0� �ȓ'�H��˛w~���L��	[dՅȓ���䛼p[b��G�IG���ȓY�\Y���F�e�>�SNu8<�ȓG�͊��#P|{wʘN`ńȓK?���R 	%�b�PQ"Ň![R-�ȓ;>���4��qp���(�+`�29�ȓ�*h4���(��P��+8YB��ȓ@����!�
J��sa�L"���ȓZ�t��K&?��*�üE��ͅ�J�m�H@�6��Y���=^O���t��RRo�3_���b��
9(>ɆȓDO����̺eT�"M���ȱ�ȓwB��QN�Mj5r!�F�=��e��5.�8�L� ^�>�!��KS=���B�,%�5� "ZV�r�]�q��X��ma�Yj'���c��E� �ȓ?̼��B$ѿM�P�j'NB?E4R�ȓǰ��5��^l�I��;3k�Іȓ<0��φ�{&hꂀIf��dFR�|b�?�KA.Ҏ�z�ۀ�N�hw���D1D���3�ه��3C��9�����#D� C���0�V`H�sO���4D�4 �h�-kANl˧�:$���S�?|O�b�<�rc�5�"�@�s���`1�>D�h[ŕ-n?�9�2ID3��X���=D����>K��d�+ϥk@��9ԫ:D�xi"m��`q,�r �I�(�n�
A%7D����U3e<	���_~ju��%6D� K!�!JV~��v�D#0��M'D��@Q��/�H��
("i۳G$��0|�# Z�-��%��� ��:be,�c��y��ߘm��<+���0i�M�f�?D��kf��$L�J9�u����a[uN0D�8k��o,�ɳ�9	Tv}R�.D���c RA��It���
2���F8D� ��J�|���� I+\��(3D�  b��I���cZ� T���0D�ؚ䦇�^�Dp����G�B�b#�/D�4��[*��\�g/�5G60�d!D��z��A�\O��Ç�V�����?D�������M�Q�5�o���9��;�2�O+R�	�f�ቕ'5,Ĉ�I�"OXy�*�2��s�h�	1��屲"Oژ����a�1;P�ÐG���CV�'^�L���M�Ќ �d޾S���C'�OzC�I�QҸXfρ�vX��׫�B�I	I3X�Z��Б�PԸ�聲(`B�ɺV7�Q�Z�Y�P(�mޱ=�B�ɱ��Mr��T�7���B��>��B�ɻK"4�bbᚵ�l���팡H��C�)� �5��f�^�t���E8��!�"O� �$�B�L)DH����p����D(LOzLzW$�z���)�h�
DA�-��"O2'�K�Z�b��c�l-��"O��
 �һ$��e:jH�9�"O�9�1�O����cd_����"O�� m_�+(�P!I�~�B�#D"O�9J�	���Hq�ɒJ�VhI�"O|�P�כ{�	q��D=^�@UZ`�|��)]����	(ľ18���	Iv�C�I]ݪ� AIяjM�Ux��N�=[�C�I�F��$*����r�IćPQ�Ѕ�w�I�1�ưon-��d�3.q4C�ɞlʤ(����b��|�q�I5�C�I)hw<š�XS׌�P$�
�C�C䉅X>�'��JM�S�ܠm�C䉓x�xxZ��G�K?��e�>E�TC�	$C�5QU��^�K@��~�$C��%
�rY�5Ô�/`&Y�r���tlC�1���CAY��ZԊ�k��H�4C�I"��s�� ,�&�ƣw�0C��JC|`��Z-c����G���(C�	�cl$J��)W��A��j��C�G����Q�,hLd&ڣ"��C�	3_"��
�����e	F*Һ:_�C�	�\.�*f���<|�r�k��f0�C䉳, Z��4��g�ms#k��d^�C�ɾ4�^�1-q!'�֑i.��=D�؋�b�0NP(ԝi�H�e�9D� y�L��<w�$KD&R�|�`aЧ�O��=E�$L� Ia�����Ҫq�vQ#SA�H�!���5I�TY��HO&���jf��0�!�, d�}13oH?�%(�?3�~a��'�R]�shًKtdB3����'����.�9W�-�䠊�|�U��'�T�� ŗ�D$n�y�&�~��)��' 6ELĕi��0XaoK.V �!�������>���ݢ�F�P��;;( ���$\�<���z�B�p�*��M��A��*�Y�<1c"&�N�P�H�zk��#@�V�<Y�_g�6�i�,R!$���gV�<�pJ���,pq�c4��srjQR�<�� ��^d���$��v��N�<��8r�a8���
d^�� M�<!�)
�>�ٺf)I�st�q2p̝a�<i3φ�9=p���&E���bW[�<)"խf�d`3m��u �8j��\�<�g윇��Q	����*z��Bp�<����~2�\���q�T��Ad�<y��ؔc��P����	Մ��q�\�<��IN=c�д������xt ���M�<Q�L�3�渀UL�>� E�P� A�<���^��h�B�%A<��d�L{�<�S�:b=VU��.F�>�°I�B�t�<������QW�#�ZT�4�s�<Idg��	��I�˃YӒY��F�<AVBP�F��e+��v�h�x6�Ax�<�qj)L�$�s

�❘��w�<1�����!�3d�4��x��k�<IS��8���3	�u�4Q��+h�<Y�G	���d&Ap��80O]�<���W�,5\��u��<���#6��Y�<��ǅ�FݦI;$�U�QJ`N�I�<AB��+$�zW_GZ� �6MKCh<	
� pi�#I#o'���s�+S��p7"OH��痒X��If_���z�"OH��j� IX���IzKde�"O~d��Ǝ`Q��`Qe��f����P"O2��7g07"@���Zh�"O�P�"�@6M��pӣ�'q`��v"O��#v��> �x$����v!��"O��(���=ܰ)F����4̩�"O�0�b�t�l��e�>�.}[�"Op)z5��9J�,��'(�:&pAڇ"O��`e矑M
�t��26Z-�B"Or��_�`lR�(�'�PǦ	e"O"�pU������� .B�"O��Qcԕ~Y�h�֯�jn"ON��uK�dafX���/LĆ�6"O�D� 	q���y�_�4�� �a"O*��c��0s�t˳���Y��ܓ�"OХ��ƍn�(m)p�y�֙i�"Ofu������8psrmG�H}d�"Oj��gC�~�bL���%tʐ�$"O&Y�e��5+TPs��-nb :�"OZ��a�\+za��I�I�/Ya � v"OBՃ2�^�}�I���H�	� "O�m"qd�j]P�Mǃ��kq"O.\��HF�]Hf��7lA�ce��`c��#LO4:�ZI��d�qjݧ$fp��"O�)#��S�h/~�s��A�X�"Oz���P
��)�#�;(_�P�"O2��*Z��z�1!�.Q�H@"O����Ic����B	5�jS�>D���/����+-d=�@=<O^"<����.(y��-�9��Q�G�u�<�eA�<�p��範�1ZX{A	�z�<��a֋���3��(�d�J�b�<���ȃ ��q�bC�*(����o�g�<�5�fe6I�3�P"#�Qe�a�<)��ɶ,D\
�g��bA$_R�<1b ^<�~xqP�؃o\x�2'D�d�<����,�p�J�	_4���A`�<i��Vp��8�5%7NN��U�^�<�p�%i��wIBYɒ�QT �]�<qա�T�)rU��?�t���h�A�<Y`�Y�.��|�@YH:�%1�JX�<�b���h�f�;A��D	��8�EH�<�I� +2�yC�''Zbu�J }�<�u��i*�b��ϸg�.!�'|�<�� ѼG��2�B�.���G�<��HM&@���I�%(�xC��Is�<A�̀?��\ a�)R�
|��k�<Q�,
2CCv���V�/�H��iM�<�r���0N���*ʙP�{�HBd�<1�-�><p��Zv�ޕ{�|%
�a�<���g���f�1P�$�Ǉ�[�<6���EY��j�^�4�h�y��|�<���8�቉�Q�M��	�`�<��'ӿo:QS�	�|�35K<T��Ң�չr�D��#�i�z�`��?D�X�ʣ	��=���\�<}�b�=D��jD9W��B$�N-`�&��!A=D�\j'�B�"�AhvL	= �Y�ь9D�9�"�.]��3u�L������<D��*�X��DI���9eʌ��Q�%D���S�2�H�@��\���(���7D�컦�R�*�Z5�s(�>Y[f���"D�� �Yuo[�I3������Q0�"O�\"�k	�C����D[l����"O���ĥ3�� r�E�>!�J�"O��2��<7Qv�!�MS+t�t��"O^u�E��'i�� #G�1��T�1D�0zē�zx ͜#�����;D�� ��H�8��cͯB� D�T*4D�T&'�R+���L�
�����3D�p��M'T|覇	�PnDiai'D��I�M��3�deꅉ%u\\z��&D�X[��Z�PQkwc��/���/1D���6��x�R�7%���gM:D��(��䐭4a�
Y�pM�0�;D���uM�G���C�P$XnA�� ;D���D(#F�PA��L:�^11..D���F�#�R���	S���q���-D�l��͊U^PD�g�΅R�R���!+D�d���	k&�TB��xB ]S��(D������)=p`T�ۮ���{�9D��ґ[�W1*[�N�&��Lh�	;D�T���\/3�֘P�I�V"p�kӨ$D��bn�<Ry����p�d��2e"D�bs�ǀ>钄peg\?P���=D�lX𡛢�n�i$J]z"A{�):D� �K�m��%x�\�0�EJ&=D��dΠ�.��,(X�2!+:D� 8���E����(J�M�e8D���o[�XK�a�!��d��,IC4D��{PFM,�B��I����>D�h�LY�G��p�%`�Je@a2R�;D���7��w>���ȵs��tZ�9D���#A�u�����4OQ��Xr�*D����� ��̐�LC�#�l� U�)D�H[B
ϛK����F�B�8�����%D��+s���3��8�P����#D�8��
1
�d�S�&`*0�&D�@�1d͜6\ddZ�]:��K��$D���@��شa�C���"cm/D�(���ڌ~��uPF��w�`L�3m#D�Dp�+���eek�+�H�b�%D�����{�v@�c��
(�S�J(D�XD#+_�5���H s��U��)D�Ѓ�B�&��UHH���H�
+D�P��/U�h�]���!x�x��N)D�8�&@ל��#j	Y��t��G)D�$+2a��M��`Q�F�
HDM+V)-D��8�
]�ZM�$'F'�;�o�<i7�V���S�,�u8�KAT�<Y��rt�1��L�\Y���J�<	ai��<t�T"�ŌA�����AI�<�*�,�����+�&8q!a�<�։R#�N]`�FL.�(� B�A�<94BK�2��R�	�"��1��B�<A� `d,h
�D<Y4��5��U�<�E�/y��5��2Y�r�!2�FO�<���F��ʆJ�t��w�E�<�t�X�\������*P"���Az�<	�n�/mT0����UZ,����m�<Qu���e��4���,B�KVh�<ѵ�<a n��0���A�˞f�<)wÏ.$b�hD7I���a�e�K�<U�#��@!�Y52�0đRoJ@�<����:��[2H$0�"�<9$�ϻi:�Q�ðlr	$C`�<� �K$jS0S��t��NX�@
�"OP8�f)x{��;�
�:y�����"O��T�8M��5��DD ��"OzD8aM��hb���7hD0V;���"O|�P�GB�x `��R�74��I�"OLL�`����aE/K4X��"O�r��rh�E��"�n�p�v"O�l�T�M!^耽a��6+ap�"OR�zp�e�f�'�̭tT@5�"O��uk�,nu���E"U����"O`�2��D����u���@iX��"O��A�O��h���d��s�"O�á�Ϲlid��ōVd�Y��"O�%*�ƥ}XVl���m�h�4"OD-a�K�	p�H{��U�IW�Q��"O���t�v� =��G��@ac"O����ڟx�%,���F�P2"OF0�dNR�Y�$ՋWj� fF��"O� Qd�!]�x�@jM�~1č#q"O�t�@)��f��Y"�$�P�"O4�L�2��AUCܢa��yA"O
y@c� (TZ�����@T��W"O�P���݁w;����Ļ94b��"O���Q �Xd�CQ�F�
/�AJ�"O`�0�d?nB�D����\� ��F"O�IreEϛ'���I�X�"O��R�,U�fe�$� 0BY�"O0�������Z%a�$ɑ21��r�"On �Ef�`c�$�P×�M.*�1U"O<u#E�\�~(9"�m8�Z�"O�$��m	xb�h�![	=v��"O���G���nĠv���~ZM�S"O^}�4��%k28�F�VV��V"O2�+�F
�)�0|R��g�����"O�a�Jϒ:���+ۏ(��ԃE"O�����D�Ĥɏ�{`�@�"O�8#�O�b;48�m��lG� ��"O���5��/�
�R�=(A��ؗ"Oh�� �Z�x �$Y�a�2Rz��"O�x$�0�� i��A�P ��P"Ob�"쏬$��W��U0�:E"Ou�a�Ki�4�����)?&H5ʇ"O6|��B�8k�Qx@�8k�>}�'"O�Ik� ,��q���ǹ!{$��P*O�gCҥc8���$Z�G-b<��'���Q����A�h-�`J	4{�m�'�DLC��BB-�*�7�x=��'b�s��-M7
��V�ʛ)��p��'	fU$�0F�9
F@��m����'֔����&W����	F��@�p�'�$���C�"�<E1�kX�}����'ب�(W�&q�е0�/�z���b�'8�!��]����$�:��8;�'�LSF�(m�N���
%5�����'�P�C��,j�^e��.a(]Q�'B���#�N(�Y��*P�\(-��'/�\��>w� �!�JC�SՐ�!	�' �Cb%X<����*�I\K�N�<I��[�j���Hۇ/��HX��p�<1�h܎I��u¦�#7�[]f�<i2���V�uA@��9f|�3"��z�<a��o���"��0>v�dk�e�p�<	� 'H��%�r'BVE;�k�o�<A������!R�əs?�h��b�s�<�  yd���<�k��>�^���"OH ��H�p�l	[JBf�8��"O<e�P�+GB�`/��� �"O���gf�Y���vn�t��`a�"O )�m�t6��P�Ix��a"O����"ьi��=�&��[6c�"O�hb���	
��$��a�M�"O,��墆(��)򍀶�j�#"O<ܸ��[-(�.8��	O�h���"OL��v�A&c�F\s��+�r�hb"O�x��2��,X5̖�}�BѢ""O���T,x��h�j*J���q�"O<���䀧j�A��hn}x�"O����I%U\ait&�D+h��s"O�|���20t]"���(+�e��"O����E�:�򈠃'�1B�Q��"O,H�aឨE�hH��R1f�H�"OK��ƈ�a��~-��z�"O�����@-ޜ��p��9��"O�)� �#Z�ּ0���e�ó"O �#tC	6$�2�ˇ��9=d�Y�"O>5)f��Ia:.�M2n܀"O�L��U*����MH����(�"O�����=�t�b�� t�`<��"O��w��z�6i�1k	_�J��s"O��A�H�*q�|� �M�M��4��"O�hZ�X"D(@�Q�_Ev�x��"O��e��4,,0q+�/eYN|9��IFX��Z�J���(7��� !�6~!�D��M��y���&
�����������(��x��3p��c�D؛d5���"O܀9�㐮G�y˵Q=5����=O���d�=?�(-��&	�uy��Wk��y�N�<�U��$K$�|��PX�#@�9�j%��+iW����G0%���/x�X���$�G	�uoZr≅	�Q���t�4�O��+nÏ&�X����]l�<�%�2�D��L��f٣���\�'axbT�'P��i�aoXU��@	��hO>���	�a~@D�ԥH�L�86:{!�$W�`.V��pd���MR�d�V_��)�'G��[��C,�(p��A�^��
�'h���1BӸ#2���m�=r�����N?a���Op�qȃ!(���Ő2K�MbDG$D�LJ�%'v�Ti2��62�5ӷcߤ��Dv����+�4���T�*����`#72��C㉙d8��Q'ǁJu�IR��S�t��	�ȓ���i�bA?jt��Adhԕ\���ȓ��pp���	-$ر
�Y���	A̓jFD�y'#B%�}�P�sE���?����~Jd�V�RMx�0?6-@pnWo�-F�<�|�@hO{S�}�Ʀ�k�V<rcll�<ѥ��P�L���ς
x@�
��@ܓ��'p���])��R�r�$�sG"�G�<=;"O��(S��x�q �"1���Y���?�S��1�D4*C9o�T�B��5��B�I�,��I#�Q�[���w�e��B�I��t�A�e��Y� ��nB�!Xq*�'�U�n��y���Nx�B�ɟp벸��@_�8��;��O-"N@C�I���u��/R\I����P�C�ɰ/�v��$�F(�ɱ��#SX�C��)�Ѫ�m	N�g,Ψ�C�	<f��t�7�P�DM�! �?wZB�I�X�R��BI�)a4!ZPCB]iDB�)� �M�"Р47�$�ƭ̎.��3"Ob��1C��a��Uh�ZW���"ORP��mi���Fm��*=L�q"Ob��D)�419�����ބz%�[��',qO� �6l���҉���,�1��"O�����د����)�4Z���"O�����"f2���;Ƞ(xr"O�ٔ��0QmF䓔�¨w |�Yq"O��D�ЏW�](���9t�C"OH3tg]��h��#GĝZ"��G6O6��D�dnLy��I�[jP����iX!�䂳-�D�т8J9�yZ5���!�"R��%ѥ��(~�*݊�cM5u�1O�7�.�S�'\0�jV�D�r����F����	O���Y~�Thn@1�T� �Ż[�D=�O�p�7J��u��0�G
�k�����Ic쓣�'L�X�Cue���I�E��D��Q��?��;�Ζ��{��~�T��yTdL'M�8R��=�wm�Z��ȓ�,x8#�����@!5��	pj�ȓB_*5���6%~���Ю���ȓG� (;��6в�9f�)a��T��U�������1�Phi�H?+q$ ���K���#P��ز����+>���+_"O�,C�Î.��0��!�!����"OB� H�&Nl�@o�~�
)Ҁ"O�"׌·8��xH�.� W� ;@X�L�'�\�FyJ~Bt��P1��e~(z��Fn�u8�$�a���*���Bq��mϛl.����5���<1�@� ,�Pr ű8>���Yr�'��aG���0D���k�N� Iy6<�N0����'�����J��T���^�D�s�'�ў�}�s�
	�0��6.��ѱ�`t�<�d̩a� %�1G�08.2���y�Ud<�<��������0��oҙ%�бY�P�E�!��`A_���pG�F��@��	,��SЋ��G?���r�[�|��U��ɺ-���D;��V�8 S��qՄ�B�D�n�qO!aӓ>�|�COֲ
T#�s� �Fx��?�lZ�wk��A��Ҁ,����NO�RC��("&yA ���a8&]RTO�b�����5JY���7�Z)��l�:�!�$[�!�(��G�K�
�%ǘIQ!�dǅ.���� N)	� aK��!�d�#U}t�&fSy"�}��7k�Op(
�H5 ���i��+�^<@��ĽN�����N�x�	��̴N�&A볅H$U������`�K㒘����=3�����eW:jO���I{N�O\x�EkԴ�6���E]�Fx�"O�E�-�d;��6Fڝi�
 ��"O�t@����ie�lA�z;�Ź��'��'���	�i��Q�µ�Q��7"�@Ղ��d9,O�������2�L���l�<5z��Q"O�i0��a5J�F�-"Oh��V�ԉ3	�icꐕ���H��'j���6�,E�Ay�knQ�a�"�.D�y ��F�%cӕ-���9��?�S�'`>D�T�-_�Va�7�^�w0�X�ȓ?lpْ�"�)Ä�6��|'���I��0=��	�����#�1���B� �p�'5�y�E@;? d��LU��$暭�yB��F<��C�k��5���K�.O��p<y����'Քx�dN�?]u18��F�Z!��Mʾ�A�#�7dX���ӊm�!�� ��.1���㧃S�.\��'E��x@���?N��i�.��0�p�Ə+D��!f�eqpA�r-�F�TpzV�	V~�2O��)��<��J��,�]����0Mkj8���]N�<a�l	1K�8Pyf��)����4d�F�'A�x�aU�6gvoK�H��qWb��y⩚;����D5>;��������yRȊ8��qBk�;���Ea��yR��]�d����!g��icm�)�y¡U4�`ɉ�S��ј+�&���3�S���>!A!��G�^�	ӄ�'&|z]��R�<Q�H*& TH�BE�S3�1T#�N�"�M#�'�qO��p���٘� �y�54v�H���7����z���':�|X���X��hO���Dŋ�XpG߇V]��Є�B�Z�ay�I�1�)�R���Q�P�˵8	�C䉫J}��3cΔGx�ؔ��)M~#=��0BI"Т��h�N�P�	�z��G�D�FbĹI-�p��`Pn��lE�'^�?7��:� �L]�&���K0d�8/!��T�H�����V���!�)i.�d@��(O?��v* Q�fՉ�&P"!]n$YB)8���*�BPl�0u��ˣ��)1v���[����=�'`ȹ7�
�t��8sft��BO�<q$�0�PUK��>F�lX��ZO�<�'�԰$� Y֎E:��y��kVL�<��㆏J0��!.y��(��H�<a�f](�0[G,�-PT4���@�<A1���\�!� �=/d���梁c����'�
ȣ�* A�6�=��pP�'*i#n�$n�xA�̆'� �'�޴�5⛜�R0ɑ�5�T y�';�5�����t� �H�>Zz�� �'�	��HO�no���@!D�a4n��'Hؑ�������0%[�F'N@y�'��@2D�[y�(s`*�7[���	�'▉qTO�H�Hڀ�]e��	�'�(�;7�������(`���'�J]IA��tmȘ��G�8ʁ�
�';LR��
>_�\��)�$/$��	�'mnh�!T@���T"����I�'���c-��H��΀��R�H	�'����ʕ�r�ģ�+5� ��'5�]��!�@�fq4@�,4�0 ;�'���j)SK�Q�`8� c�<�P)նI�.!��B�8�����\�<���O<�>M��Z�P�>m�djU�<9�$Ϙ~$&�Hb���M+ē#�>C�%t(�H�AL�>�J�Ͼuc:C�	2<�xx:g�O�b��h��e�*C�!8��5
h�".V�IwE �[�C�I�O�����Ō^�l�2��ڄC�ɁV�v� '��,����B9i�4B�?��3��վ;"R�)��0v=rB�I?��Jiћ0W"Y�w���C�ɶ;W��iV��h�$Я��B�I�'���1�NX>JBF�RI�S��B�I�ܱ��C^u hi,�	BB�IW�L����5�,�96�3��C�Ɏ}B:|B��,�P�pk�j`�C�ɰi���s�D1&0��ia��)��C�IKFY��259��a��z�C�I 0���F�1��8����p�R���˻{��Q�h�-J <��W'T.LLb1�'Ԙz�!�� ��k!*��|���ԍ�H���"O� ��A5]sr`�E�'�&�r�"O�`X`�I%Q�0���,a�Ay�"OR	��NB	o/�����3b�F��"O��S�(�NP6   qk���#�"O���EI
�* �k��%N��	�f"O���E�l�0��<8�vT��"O~X��ͮ,�����As�q�5"O���u"ƈ&���F坂��q3"OF�ICn�@�`h�*!(逼yq"Olm2�/��P�r��.�Bya�"OZ9�����B���G�H`�"Ov��O�6T&ڀ�=���d"O�3`M�w6jhr�V3�� �"O ���#e/����ʕu�` ��"O����)y���"T�*� Z"O�E���@+r(�T��dߟy�tD�&"O���&ZV�E�R�[�F�
�'���'JQW��a�f,^x���'^X�mA�J�����F���݆ʓamH%	6fA8��3��Ӆ�N���giv��pcR�1E��+�a��^\�x���U��O�,hCUOɊFr�1c"O
x�נڊe�e!#�_�|+Txp�"O����3�m Tl�{x�!��"O
� �
�o+$�m �!f(�Z"O�|S�#d��4r�'�;H>IxB"O����J�~�:4�7�ʨS9н9u"O:��ɕ�g�2}ysFNH�"�"Ol���*�r���F��".h�0D"O�!�F�Cs��qᱥ��f���"OB�Z���	�qz ��[��u�A"O��A��U�Va�U�\�k ܑ�"O
����&l�hrG�R�N�8�"O.���!j�����3>����u"O~8��.ě9w\a�6���s`"Oʁ�SÚ=�FQ��Ѝcڈɚ"O��sqV�M��Y��ǰ(˘�h2"O>���52�>!RU��!�,u�6"Or雂k
6:�~Hq@ķ�nU��"O���eZ#v?�}�� [7�X��"O
Hv�J�`�u�fN�aif@��"O�A���*C��#Ql^�A6~�"O�A@υ�	�Ƞ0׫ߐ9�&�s�"O����b~�%+Pi�X~�1W�')�����,I�'J�10�nh ޼H�ǐ/ �|1��'�r`�#M̩A�Xz�EN*8�eK�O�%���Vx��N�"|
�$�Z��W�0��c�m�<��o@jјr
�7^���Qc�:dtU�'�l��fY�ϸ'w�dstaՠDwr|�J��e���{��6s�D#�cՐ�x�����T�I�;.2B%ٱN��0?��ދY��I�'[�*���K�'-lA8� $�xIH�?��G���:p���Ѩv���Q�-D�L���ˊG�0@�7ɏ<}f�����<�P�^&9� ��'�0|ʔn C�>%1�DjNj\�pB|B�	�K-�mI¨��L��D`��y!l�����<!���v���M~�=	ƖD�D0�!�U�Գ'�e��P*v�O���ȑ\�Bv�U|�DY�Ȁ���9os�d�$��/P����`�� ���?I��u�N�b��1��Iʇ����&��e5U#���~!��Y0(������;*�ɛ�j�1ly��?s^��g�Չb��S�ϥ�ϧ3���8&`Ԯ Y�H���^�<�c�:9�f9���إkFT��'i�:�'GP��)[�g�g�d}��T���+d�!N<�B�)� ���⃷T�)k�+� �6��s"O�i��%�|�Ǡ��8ɑ�"O&�S��ܖ%�0�"��. ��!"O"Yx^
��M��o>,���y�e�����GJ�d^Ա���:CZr�(�{�(a���Ğ�s&P���C��a�j��{!��J%#6@Ka��Y�`%��_-=`�\"�C�$(����"8�iBbI�	�~�0�S�cV�x䉉$�*���-Np��"~
��r���JP�E�B��5b?�C�	 EP�Ѳe�_3��c�#��;�nDKUƗ"L��"��ob�C!ɇ�"2~Q�A�O=(�zC�	�����U|-~��g�ͰB|��A�)�~��?i�	�S���{�IښrZj<��G�'f� �"�=��?��ژw�`��Ϝ� B�a�#E���ǀ�h��Q�P`$�Oq����Q�6�����$:̸��	
xuPɺ`��8h���V?-آ`=vU8����6�rͰ!+3D��r��%s�����١���v�`y�GĔ"�UKjZs�^�D��oV:f(����!1�t9�B��yr��5y�%��͋(HX؈�+Z`E���=޾��`�.���(��y�#=��F�2a��T��E,��;�n�~؞��(��}c�	˧A�>0���6,ݹR���s��^�k�l����<i�؍;��'[������~0f ����T7h�{R�E�	���-�4�T�A�Ѕ�X��OD��,�<�����7@��qz�'�ډrW�J�6JyQ�# ��l����*r͠�y#���9�J��=�(�h���@���J򔭑��R�5쮍��s^�b�$��oL���B$�9���EQ*SAܨ�$؛/F��3!H?s\�>�cӽ8��`�)�3h!�B��xbE�͆].8��W�N�naH��ۖJ�bS��"K㐁RQ�����}���rP]�B_�4��e��V6żd�=�'��dR�5�ӪB�`�n�)n�	~��G3��"�Ȅ�9�T�0"DQ�Ն��	Ó�о�&LKB�$Ht�b��28� ��`�B�"�"h��Wm�O|�	�Wj�0Id'�aZ�-AQ�ĩb��C�ɔv�*8�%�ٶ#���(D�$�PI7_��}"���9�V�)�A�v�R*Y7! ��&��C��C�J螜�ħ/eL�B�-lO������kY*�1�@WHm>��e�
�v��ibEψ�Ge�<�$f�9]��6��1O���҈,,O�<(e)"Y�X)p��-���
��'QR�2���U?qu&�(Fa�]�PC�Dђ���Y(^��E
¬�K̭WV*A!:)�Vh��C�P����*[_��%�E��yP��`��	-@(�H�H���0Au\��2(�/D,�t�C�	
3Q��X�k�0{N<
TI��zz�|�h$"������%e�H��2MĀTLF�)��D'F�PyV��,�J$(�E�QlFlZDN�T�'RiB�'��<K��ΰJd�����'<�4���Ð*��6α˸Oj�5��H�>2]��Z�@��TԀT�Սڿ��3õiI�Uj�/��Y���*U+H�� ъWd�c�](>y��B�bĨl
�� 6}�O��P�៌����)S'\Xڃ�E
(�^�; MU�z����Y$?���Y�1�T�5	�E��d���T7���B-2B`���C�y��0�rS��a�4��%y��H�i�y@«�m�����'T�}�d�$hN���2ǌ�g� �`B*`nV���D�<9!Ƌ6>�:�&%}��)�����[��\�U�x�5Y�Q�X�)����{��ӔB�������Q0�5{U�čm��2�l�;V�M������F�����P�R���˲"��0�0�;1d;O�;��>�BA��O�D Y�,�C�Y!���ls��H�0w�`C�	��1�UB�)r&�4e9Z��Z�X�cA� ���G�w	hŲ��*��O9��%����݂��٪Q*�u�
�Q(�}��#m�|<��e� �Y�'?z�Ͱ5�'Y�ఁ[�D~ O?a�$��>l�A�u�0L���b�G�<i�(،+�$��Ƣ�P�Ը1�cU~}2!���L�R��'U@��T`�<`�`I@4&o,Ip� Ӓ��T!ݔ�8h��� ����>�:pA:D�LC���;4���������a�<	rC�=,�ć4[��D�� ����X�a�.Yo��!���<�&yK�"O���-�.)�H�j�E=B��@i&�X;�V��Ʌ-%�V�;Ċ��g��XO�c�,q
1�Pa�	�07�ة��1�O�ܹסу�8� �{���h
e�:��@�>	����7nJ��N�h�3LO�9�s�!O���ٕ�y���	.!���#�&S����p�L?��b�,��� ��aPE+���Ó"�Px�Q"O�p��$p�񚦥\�r^�xz��i߲�Tnߡ]Ժ��NK�Nk��D�3J��c?�X�{~XH �KŬbF؉�bH��B�I�Ux�Ǐ7Qp���\�f]B�2� фTx�xSŇ�ZFڵS���?��c��+?1On8����<[��� a�*`��ag�'��mK獜/�M��&4I��y+ç�DA�m�cD̓~c,X�di�0y�]`4$8\O�姝��bͺ�G\7<��<aቒ&Ϩ���ιP�����I9l{%i�l�>�uǤ�"u�i�7`��N|�)�v��y�ݿh|0��A��@j�0I��ܵ^��������aJ�p��M��s����C�o���B�Ҩ �:�f.D�P��K؆+}�B�"P�G��53Ճ̈́\��m���^)p'�4*\�V7��F�'��I��ޗ�<��i�uB�N��+"��}ꜜ
�����J*0[�h t�%x�4)��$m����I)*����]�y���5`L	F��#<!��>Q
x���ʸ*�,)�e� ��	A�@,$����2g=�ՈX�G�!��ف@; P �!ܷA��Y��g��r��(����M{��7[r�׈Y�A9$T�~λ3*��	�3whQ�S�D����	M�u�28O �5�@�wR� pC�ȏy�J�QG@^� �I'%H�3m���g�Ńr��vW�<0�{�Ǌʪ0(宀� ��kբہ�OX|��Ȏ#��G�R���L!V�r�я�D���]�oR �&��.@�p�ěs+���� %LO<�(wŜu	���e*ъ&>pBe���q�^�i�`Ky�I�?�g\�$*j�j���
�D5�"\!6���B 猞9"y�I՘b4��ȓ����MI
�X��˛Y�j�o�2] �������uYcۏq+��ۑ
�]�P?Z�_xu��#M�c�����#L��{B�L]�����æ�� ��7	�-��k�����a�
���s �?q�d��̏+��'ݐ䡣��֧z���J3JCk�1*EfKd��O�xQ �\�I�,��M����`Y:Y��UZ�%\�6/�)��c�0�>�q+��W_��@����6�)QsJSZ���1�b0�|j��G4&��Á��/��A�#����ɷ]6��slFN����F��q2�U�㚾w�T�e&�Jn�X&�86���ȓYj:S%�ɵ*3Z�АB9����	0W��p�ԍ� ���=Zm4C��/9J���T���ZH�#�/�����M�;��=a�Ocݪ�v�z�ޠ�#�[(��!8�g,R�H��ʍ�9w���7(���)��<�Qz4@��K@`��r@��k�'�)QuhW6%��>͛�;O�ҵ"B�/j�>���|���c|U��W4��y�e����ғ˜�'�b�p��F9:M�(�=E��,�� �N�s��dQg���?8���ȓ�~uy��ݾ-�$m��Oƨ&�9�ȓ���{��o�&8	�)F�M�x��ȓc@ʵ�P��C|��1�+-�@��ȓ`�x���Su�dhT�R�q��Ԇ�sc�`����Cg�YC�x�ȓ3����/J�@%�T&z(4���o0��Y �Ę(M���B(����]�Ҁ��S�n��~��mh�#�e�<"(YĒ���ԧK�$���[]�<y�,A���B�h�:#	��.W^�<�$�j�,��l˨�p�)�+Br�<�uJY��8ت�*E��!��Im�<Id�*Q�� _&-�$UЅ�n�<y7	��JD��:�� Q�"A\�<�� �%�j�Q�� <��I���\�<Y��ڦK���e�iq���Tf�D�<��AV	P�dH!����A7)C�<��!�v���s�+��"��7���y��P�`��i�Bh��a^�{�
!�y���y*��05j4�tĐQd�9�y�*L�VY�Fɛ7*��Q�T8�yrm,�5H�Ȟ�)��%"�b�$�yc�%O��p��k�|� ī�JL�<���7f^LQS�YT�r�X�/DM�<ɠ�Ru8�9��b46R0XT�D�<	����T�hѲǃO�9�%qe��@�<�s�Kg�Vђ�g��X`�8a��<�&ƛ�,L���11���@2&�z�<� XQ�
Ʋ'�3��H$L9Q"O~�vo��D��*®Y^�8�"O����X�2& p�m��M
t)�"O � �훣m�H{���o���!�"O�Q���T&V_��b�HS/ɚh 4"O�Q��Zh����'Fֻn�l�:�"O�D���-�A蔥�J���"OX�J�V|,�$
R�6�6�b�"O┛��\&y��#B
��d��ܘw"O�q���%
��3&��w��+�"O�@
���]x(�P�hP�Gb��H�"O��������h�G��A7F��G"O&ՈEzT� (]%�䋥"Ox�c�BאZX�a��J�(�I��"O��A��Y�}a8��A&ܔ_ ��(�"O̵�v���q&�(ivG�����"O��$*��z��31C��1��-�"O�	�Gn�%QC@d�"/�nQd�V"O0 ����\�l -5?�f�c�"OB��u��Ka�Q3'�7E�~xk�"OP�v�[70��rH����uX�"O���bE���X1f�S�{�`�"O =Q��C�N){歉�PҢ�5"O@�Q���<��܊fL�E-R�A3"O���C>
��`@j9_���3"O�t{sʉ	lXl9�iU�G��Hac"O0(p�K΃-7�����	H�.�r�"O�p��3qF���ǫH�@�PiA "O��S�H3*p^s�]:q^A�"Ofڰ
��X��yPB�$ɫ�"O�[�L(v��p3�Ĵ���cC"O.hq�$T<��C�C	=�,{�"Ov�p�U�L�$}Э�0C��Ka"Of���G�&�R��C�>� ۆ"O���0G�g����'��~�<q�"On��pd��@��ЮE�R�iS"Op�S�GB�}q��z�h��%�n$��"O���`P������?ZٶI0"O,`�[(y��A��r��"O�)��'Zp��qWA���5r�"O�ҡ���<�Dh@%!I���g"O��q�.X*|�J"WF <a���4"O�p�HΒZa��Z��[H��m�"O�l;�A������+V�2���"O�<�p���MΘ��1�ʱv8����"O�|����O�$����H�(�	��"O촓p�×
���K��Y5*�T�R"O`L��	��;�r�ه(�2��b�"O���֫-s�U�D�*������'����w�R��'�~H��
��D1��`C�֋O��H�
�'Լ�
u�Jq�)�kفU����O>,s��3��)@O�"|�4�0<�L2wjݒ
R]z�'�X�<a�g*s�)ѣ�!ZL�=�7�%x⥖'�l%��h�ke�ϸ'�0y�ǖ��[(ɱ<����
��-�<Y����1c��dK�����4Ӄ��^EJ5c��L��0?i�-�"S�"�Ζ""9��9O��6��y�<)q�("��Q/d�&%��k�%V�Ls1�s�<q&"cH0槗+E����el�Pyb`X�[�
�R�KV07Aa����fpx4�
�	[���b`��y"��<J(3sJ5��-�����s(OP�l�5n��qO4aW���$!"�O[�Z��}���',!�!P��@����q�H�Q�����:`	UH�a~∑� ��p#%<`
]����?��O���"M#��9 T�.U�J%5���SB®8�F�Q%�h�<� �	x�EةG,�#��1�p10#�� H��F�=gd�rp�>E���N=Ux���d\�S5K ��y�A3]�VYc�@)]�ϊ5�O�4�
����NT�
�'�>����7G��^�p4�ȓ8�����&�p4�@�U�26 �ȓ&��p�۩d�l⥫��-�`��,�*\��`ϣ<~�8
�㚎+�&E�ȓ9�2u�K�<����g��A�܅�f1�!H��̿9KXP�A�[踹q6�^Bܓt�آ|�'�N����
r��#u�S�y�z��
�'�T Ae�
\�D�����t�" �uՁQL��U�'�Z@ �#��.�0�h� `��{�LL�l@ #P"F��eH�O�d���@%gT0[RFț'-|h2"O��Z�L�f�=�H٘_
���w��`k��ѳ2�  C/��ȟ���m�H�D)��e�4@��-�4"OV�+C ]>A���K1(���zD��7�=�0Z�Y1��V!��g�y�PĀF�%!�xD�t`ì������/{�@�8Հ����@�gS�aY��ju������`�'�*�BG�N+H��V�Æ'-P����D] 9�8�:P�Y�	��P��N��TDˌOp�ḗm�-a9��ђ"O0���5Ģ�1�Κ)@�҇U���F�=g�P�J��?}3"�RnhjX���	C�h##�&D����T� �� �ѣZ)c�Z��f�);gB�
��=��
�.��k\ ��ԑ�HOL�[u�H<U��'L�3��	�'��Y�3���"@�x7��V�� J[�d	��k��B���8�IPr����I�����jV�$�F�:p�̲@v����#�fI��-/T��9�g*T�:d��G&(��6l��ebD�1�f���C�I�4(ād(��8���s�E��CK���{� C�8v� �!=ʧ�����*�b�@Q�σT���⋏t�!�$��V̌��4�D��2�𡂪 ���H��I;O�X�ѧ��� ��Q�h�F}� �4�.9CcN��@���7+���p=����,���r�m�����Q�^K����	��:Y����OC{�-ɕ�'�y�!!��QT�F�:�k7	����'ީ���ڿ�6ɀ��Q*���.��'8ȳ�bE(90bp�R(t�����+�=Yv��O/&]����jl܁�Z�aq`Y꤂R�z��ؑ��y�On���	V���3�n�L���8t���mSJC�	�eITi�s��.?U��h#�7H�^�{��7>� ��S%�4�H�T�8eKO�=W��$���#�%o��w�L�K��1���>lO�I#	�?$;Zك�,L�ȼ*`�o����k56��1��	M)�h6m_�53r��1,OJ�hq�X�y�JR e�P�`@1f�'����a?�&C
1'`�1^�H�Hd ���Ő2�*"�*��;%�F����ɲNB&��I����d3��5!�@7$�B%!L��	�O4����(EF i"�
s��ʰD�!Z����U�(J{�8�q�@�Ee�T��'�Y#�'`P)�m�<p��T�ԽxD�����X҄�g�A3H9T����?=�p��|���4}��9^!�ql�c�rH��ѿ�(O�;��<V1���T���Yk��e��y
�`I�^<n�����^�^��)���۷-Cw8��Bo��-x�Afϕ�>���5E ��Xƙg�Xӧ����e�X]�	�[�D�q�/
�HrX� ��|<��'W|�"��
O�A�ƕ>�I�a�*���B�O���H��Z�0�'�¼��C����O�	
�GY���
�C�o�k��|"�E�hض�ӲE�ڔ��ci@�?���E�����?�������]��ӧ���h��U�4$���-��/ty���	�[��98 �Ԛ6&>I�Em
yu"� A�	 ��a�/?�c��.� �6O�H1Gk��s
�b�d�7�O�qg�L!�I/p�di��>����\<U��B�)S�|>BAU�ܠ_�,e�v ֐�0C�	�S�@�z�(��$��D��FƳk!��Ec�1	���$���?��9:��)��O<�
"L:v4H<ӂ�A�(
V1�Op�80����M���"zd�!��e>���HEџ$�g�N; .!�I<E��+28{��?M\� �)CH!��&\R�����&	��!�)�� R��\�$a��La��P O2~�Q'�
O~��R�(�O>U��L�@h !�xC�N'>,VEzT�B�(ÔH��ϔ(ɀ���,-�52�8[w�\GyR�M4ŀ ��T�O02�q @����Cʸt��l���� �ɪa�ƦxD�08g$�@�a�,Az\�D�qt�S��?9gI_�vq��D��l!Ca��k�<y7 � "��	
�#�����.{?A�ּN_�4��M=LOr	ĥ��,���=��j��'��\C�+��Dy9dHB�J��P��cJ.,J 5��A[�<1��1_j�([્+	���� �Y�'��qQ�3[l� G���v-"��tH#tn�Q���(�y��9-�v��Ϫ��d(0-�Z��2�א(��I�"~�	�l�f�p.�)Kn(�h�n�B䉙���T吣a�( �&�>p��*��g�� �p=�FAH.j��Q@�<���.�{x���6nE;k�VM��y��O�!HxH�Sn��y�$�'5���b�ʄ&"\���C�y�Bƍ$(ȉ9�b�&(��#B��y���2aY�K5m�W�ސ҃(��y2�=|�FU�E�����r�	&�yb�@%{�:�*�,W�@ac3��1�!�d�*m�Ä-K�m���#$���q!�DV�cL0�"�nF=��)����
7�!�DĀS&|��a�\�2�X��"��.�Q����D�R$x�E�4�֥D����-T���9)a�\��p>A��1s��	-t��x�芮�H����=Z	��R��Y
u���:!�>E��'C���s&�:�1c	-� lJ��$��Ol����,�'I]>h�0l
�fJxyw�CBE�Ɇƪ�S�dW�r"T܄鉃 �`���N�0YD0ۣl�!@�@1 ��>K��K��&?�@�GX�F�b�2p��,0��8�c@�G�D��$�=`@�,�ȓ)H��D Ů^y�b��r=�ɈBBĊ���.�X��P�а/D�xT��lyJ?P��|!��T�^|�pb��6|O�A���F#1b	@�4�D�ه�AOF�{�H1ej
�j`Uz�ԡ�Txy��D@BCڛG:�|XF"X-��A!�2�I�*�q�@�G55��>������g��M��J����9@l�O�@��ۧ|����1(9LO�%����3�.���3c˫��~N�͓6��&	����U��9��&�P�w�]� $��gQ1���C�y"��Z.�2'��GD���tÉ�?��%R+v��A��	L5�p�Pf�X(�j/O�$T�l�!�I�[(b-��[�::u���y��a�%U���I91�����B�\�^B���$ܙPM��Qc+}��9O$ ��a���S�O ,7N��	VD
<` ��Y�OlI�)J�WZ�U° �Y� ��'P.��r풆�a{�j����c��ڑR@�$PI�(��ı��_�Ƹ������-�|0c��
8�� �̇��y�ϛC�AAJ�0kX@��C [%�y2!P�# HB5��ai:I�!	��yF�T#��;�l��k�f��PF��y2M6��QF��[lv��� �;�y�N�3��H���CWQ�<Ң獚�y�N$>(MA�ԐO��x�a�á�yr埿c��Qg��&=	ԁ��iŻ�y��M5���c��D�[ъE�y��� #�jqX�&��i�zz��M�y��HW��;���1� ��Ɓ�y2@ΫQ!��h�G��I�C���y�BE:jX����*��lp��:�y�/ur�K䔿"T�ǦO �yrmN�ْQ�`F��A��C��y � 
��{��-n�X7)��!��S�I�h�P t�*��1욢'Y!��Y��� ��i��<xR�T�$�!�$*Fq��2a���UwD��#,�!򤒙Y��O�q{l)t�Ҽ	�!�d�I���Fd�R"���6�!��> �Pe���)[��bg�
9h!�еh��tH�)~D4� #E�	�!��9�@���L�D���TCK�c0!򤆲FGܴ󳋘@zlC�T�|!�� ���(9�.xJ����E���3�"O|E�:_�L+��rZ���"OШAå��L�P�gޅ��9b"Op�GO�W�f1{g(X���,�%"O�D ��x��<�5h�,O�$�Q"O�����.[�ݱug�A7RXs"Op���L��W� d2ed <-�� g�'�p��uKV6a�|��	V#����GF�j�k�'�L���Ѐ/�t�I!�Q03(\��'�H�!U�#p]DMѰm3)�h��'���g�,ԁѦ��+T�k�'���'J=�ƨZo� <[����'�����%$�A�+�!�Iz
�'��XQ����z�b��F�L�x
�'�����}��K�a��%-Rx�<9�Ƒ@"ι�v��C��ᯟ\�<9.�#z�نGĨzE, r�Z�<�Fn�6SV-E̅(i���S@ɖ]�<I�M��@Q��H檃�/D@q30�s�<ٱb�%��KX=s��)��Gg�<�"ER�9�2�C˶,r�a��,Xe�<����c��U���P��6U�OHi�j��!�'K����*G�{��y��37w`E�O��� �O���0�q����&�? �������2Ю�Qn���Z�:�(l]ر�_w����'�$})E�N�1��A�֪U+N%b�Ru� s�\4k���X�R��~�*�
Y���uMذ���q�\�.����k(]ֆ	��O���)R�7�p��t���$a��@.'� ap)�Mf��5p=y��IS�)���`����ɁD��Y�%���0, *�O�@t�ەq]����;�b�}�*M�`�� ��/2+X1��ũ�?��.�!��*���c_\������m#T�W��Ј2��h~��-��BdxQ��OA(������1�>��7��%HU���,���J �P&��q�T$�'�N@���	�|��NL�bAp� 9B�6�𮖙��'4����~��/��G*��;5$ܵA��KKU�<A��)ƀks�;QX�� ]�<I�޾#���z%,�::EB�d�t�<�@��oc��f	!JR��I\�<����%j؍b&^6@pXG�HY�<����nF��d��&~}�e"V�<�q�Z%�z���@Y�,B��h��}�<YC
��!8dY���q{�H��x�<	�BӺ0��(X��-�D9���p�<1FΌ=*�Hd�1�O6C���'Fj�<12 RM�h�E�8xGp�Cu�P�<!�'��R.�KD �1Ek�a�DN�<9��N�Q�l�DD��#e��fa�N�<�U	A�����*��)�c]o�<�t(PE?f(s���>�����li�<Q�,%h���&@��޲A˗�`�<A1�D(I8���%װ�YC%ZX�<	ģ\� �9scX<��1��Y�<���Z5�<}۲�	�<s��:�/EV�<�0 B��֩kӉĬ�4H�2�Al�<��ML^Q�C�īB�
ܩB`�`�<IV�ǈMg�<��L>7*����LZ�<y�)�7"�A���B�H	C�`�<!��ǅJp�AeI�z)��h�s�<	fІQ(��w�K.�nUH"n�k�<�$�H�����v�t@$��U�h!�ȓj��Ƀ"�·M�� �㉖7�~�ȓ79ЂGCŶ.���"A	_�h���'��y¤ 9 ��à�H�<Zd�ȓD|8�ԊO�hs�`�uE@p}��w�T�Y�gҜ_�dCpk�L�u�ȓ*�!�O� +*����R4R����S�? ~ec��<"�T�s�酒;�vy`1"O��ui� N�A��yږ`Cf"OV`�a�ӏ@3��[ȃ8����d"O��c���'!"�\(���>��\�#"OI��b��
Z��I/Ƌ�����"OFu�!�@}InhxF��=#V��"O��G�9c��!�tl	�88���"O���T��0Z��8�>�bU"Or���"
T�(�Z�J��oy>��"O�P�b���Ze���^���a"O��	�!K�IqبP�ˊaX��sC"O䌣��. |�M�WZ��
�"O r�Ҍ@N��a^�/��q1"O.�Y��1��F~��`�"OXIc�,�X�n�q�m�(&�@�T"O6�����X��|��&��0|b��"O���!�����!'G��h�8��"O�0�S�ƭR ��[�x8�"O u6R=#4@HuǓ,#��i��"O:܈��
�GfR�jRĉF�t��S"O��LG��(�"�R�e�Xl"O�|��N�^�R|�U$.���$"O�A��W�ͤ�8�H��9`"O � �I�F�~	IP!ߕ���*�"Od����F���1��]˒���"O>	je�3d�}I"h�k����"ORX��� @٤�B'�,�Xe�F"O�� Q�ؑ3��s��
�"��P��"O&�xsɥp6��(�dI!od�hI"O�l�P�l(���Wf=�w"O��J6��:6�,`³�&n�#"Ov���ĎKj�c��9jd s"Ox0VB��R2lC���7�`P�"O�@[B"�&�����ʁd���"�"O`rV�׃, ��'��pӢQ�"O��6��!ڞdH1/�X�jd"OҰ�Vo�+|��	�N�N�N]�S"O.8I�͘�@��*��zi�� �"O��؄�"L����6N�I�İ��"Ox��\`�e���CaqգE"O�\a��4`(ܪ7N��uZ�j`"O�|��RЭ��K�u#֤�"On]����	&��U�O����"O�} v�Oj�9����
�P��"O�@K�/�6d���Y�E_ .�<�"Op�p�뚕OA"�b��5�l��"O�h��%F�Om  ���M5�u"O��b����A[���F|�R"Oށz3-G�v ����
]$D����"O��9񎘺|���2�h�7�Xu"Of�����&J�X�˄�J�d���"O6\"��:T�����K�h�,�h�"O��ȇCB�|� �{�$�2f�<=0"O4%i`	�1�:|"7����<P�D"O�����D��A����<��K"O`@� d��ɱ0 �9�\��"O�4 ���4s��y�Q��:ɬ�Q�"ON�J���9���GD�q�4��U"O�𙤇��`��5mD|�@���"O =����wu�c ,̤t9)�"O�S#gB�	���LC<p���d"O"h.eD�1e';P�F�B�mǳ�y2
�-=�Ƅ���"P� ��6��y����'�p8��[${�Jw����y
� *��2,B�M� �d�W4�X	�"Op�A�"��p�)xS/�bf�
�"O�E�e(B3
�(�����RXH1"O�30(�sC�x�v�F�|Pz��$"Oι�RO�@�U[5�3%<R(	�"Oj5��Gf~e���פ%r$"O��a�M�8�V�$	�	�T"O��S���	����^y"O�=��F��:P��g�E�Dct"O��f�׭+��|���5A����!"Od�r�Y�tŨ��S(Pջ�"O��V�h:�ö"	>l 8IY$"O��u 	=:T�x��^7�x��"OڰX��<4�2��G�X;;�#"O訣��,�Q�$.�QsT�A�"O�$*j�8������*n��ڧ"O(غ��T����H>n�:��"O0l��(�*]]�yQ�╺d���b�"O4�S`&�=z�(y���*�<cV"OfHS6n�H0���`�<T|�[�"O:�h�=g>�����J
!��[a"Oxj�A�ub,�^�a��)"ON�sY�b<��-�c��ձV
4�y�i�$G��T
1�M`\Х��A�y2Œ	��Djv�$X����5�V�y�U�\�|pv�_7!��QV��y2��H�0i& E�B���5�-�y�f]�#Ų܀t�<�`x�j��y�@424�d�7
Z�3Z�}�$D���y�ٕ+�\�@k �%eF(:�m�0�y�A����\2�ʄ>H"�[b"���y�M��V�"�0��Q�Fk<8"Ql�Py�&��sr&�V��U7�0��X_�<)g�V8�@�3g�F.�R�Y�<�e.�<B�������1Z��p��Ya�<)1c�60��\��+n�� h^g�<!�����R ���0,U���_�<y ��{�쐉�HQN�Z�Y�� Z�<�	��Ո�R��a؊&�S�<�C�N�0ș�M��k��x�f`�O�<iB�z����
Px�d�0��Q�<�qBɞn?�} �k	x���j�SR�<��սg�F�x�A�p��K@�QO�<�#��Ccؘ��EE�l� ��e��H�<���1����W%[?,�Z"Õ@�<i�W>l���3�b�9�����Ac�<9ċP��^h�[B�5p�D\�f��B䉕0�ly���Йw!�Q��+�?m@�B�	�{ݲ�S��>)��!�r��s��B�	70�*L�uJJ(&��`)��w��B�I�@��t�����L���� iK-�JB䉐!���Eq�Pmh��ƹH�`B�<5+�1�2��?4�,��iF
hd$B�ɠ94��a�K��3+D�8çE�i�B�I(ow�ԋ4B��+�ظѤ�/�C�	B���-
bG�-yeb�B�ɄF����2��Z{�}8 )Ыa�bB�6P�T�G��:p*����C��C�	�-(ȳ%`O�T���g�M}8�C�I�a��@ �Ä�]Ŝ��Ԭ�'4*B�I<T�<�#���X^�͐�`A�5k�B�I�:��!zbeT}�T�Q �C��2e<B�BT���V	X�H��d�~C�I6Rd��
��Riؠ1&Z�H1�C�)� �����<�81���ܬzWh�c�"O2)A��K�\�BE�![��X�"O��
�Zz��&�(CMб��"O��Q`�,z��(cт�,n/\X�"O�)�p���J,�����"OX��NCh΄�dB�k� �"O4� �H�.�n�Ňʭ}��P�"Of�4�? ���&H�<R�T(p"O��C.\/&��FEˠ=<%S&"Oy��J՛;`E�bmN�($r�i"O���4�\d-`NBV���s�"O>ᕅD K�(�:�	�e��%{�"O��
ǩ	S��
���9V��ɠ"O�Tpe-�>N��ѻ�EVr $�"O��A��3̶X`���02P��&"ODq���>2u�r'-KrH�V"O� �aE%V��2K 6�P�;�"O���J6 $�|�PC��M�6�p�"O�e��V��*(G�L�Z[�"O��B_�����ǻ�6�"O�؀��l���r6�]<,l�R�"O��1W�< �b٨���a��"O���X�F�\u�E�0[KB��"OV�I%E 5kX�����ǭ=z P"OX��W��oO1�J׀@1�m8$"O�pA�F�b��)�=6���"Ort�%��Z'b��GnqZ�"O�P3��z�9���ȅ]�Yۢ"O�!Ԥ�����S�/f��"O�hkp���NN����$"O��"O��f�F�Z�!԰Mڀ!�"O�F熩߆���n��D"O�A�2Y��|
%m@ն {�"OR�3N>��Qb��K(a�xܫ�"OH�e%#&�xk�j�-C��lB`"O�q[3o
�~.��rήF�5iQ"O�X�   � O�  T�  �  Y�  ��  ��  D�  ��  ��  >�  ��  9�  � (	 � ( � $# g) �/ }6 |= �C �L V �\ �d %n u a{ �� � A�  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6j�V����2�81�8	q�G��Q�O/�yRL	0���(%�B��a�B���yb�'nP(7'�7@��*T!�/�����'�$ģ�ȑ+�&4�3iйڐ$��'��HSB��&-"m��+�1~�=��'縜P��5f�0r��
�g���J�'��P���Y�X�kG�`�6%X�'l�e�&/oøBu��@(�x�'	|x
��P�2�9���-o�h��'g�$�e�|[z�Bd�)j�ҥ��'б���͆;R��І6`�6�1�'IBk�ݚDA¸�`-�C6`�ʓ!
���s(���@F ����J�RT�HĆR�B(��h^0*rB��ȓ`&6�h
�;5�Q��Q�1�ȓY;��2j_���d@.6$����a%,����7&���*��S�p�ȓ�dp�Ã���h�E����@ ����c��!z�y���=�\��lb�����'�:X��W;x�F؆ȓe"�� ��}�K�d�1T�����IAę���݀}��3\ib���"O����AB�X��S$�P�E��B3"O���C1eB��7���A���!"O �`�-���ӣA�w�h5�"O�R�ļbi �b��=����"O��S�H�]ں�a��ޞ�Hx�"O�eq�bֶE^�%�5N�$bv(�ȁ"Oʐ��HU/��؁B$�#��m�<a��ߔ$�q` L�	\$���d�<� ��"U��%�kR4+_�Q13"O���g��H�"���	qx����"O��#Ukܔ.T����=Uu ]�r"OT������yK� җ!�"\h��"Or]ѣЗq��Jwa��pZB��"O�c���#}5r� ���ES\9�"OT���,�*v��x�A�m��`x�"O�TSp-μ'*qB植�w��Pi�"O���&�H�p���f �U?��P"O��Ň
d��J���8B6ta"O"u����
C��ҷE.G�����"O��լ�"M�����$�}����"Ox���X�l�$�����/Ѵp"O`4KR��^�d8s�&�r���"O�<��O�E�08y�B���"O�J�`C�;���_.J�H��"ON�3��&��HT��0�z1�"OD8f��J\�eȜ
p��Qx"O����Iƾc����� %�:��"OFPAw�+kvȰ�ߍ.e�䊰"O4Q����M��S&a�*2ƍS�"O��HJT�c�x{���$挊�"O6)%F��
z E�cϔ-gxK�"O��Y�nˎqC��Co+Bʰ\H�"O��J��jENUz�IE�:�`""OT�PC �t���"S���P���"OȊ���9���b�ɛp�D�0"O�����oh1#�)�&�>���"O�܊aoO?���3E�V�����"O�pR�"�[���mD�-4(��"O ���ꞏ]�\r'M 7�@�T"O8����+L�ȱ�ʐ�$�$��1"O��ۗ$��,J�ç7+�X�"O��"A��Lk0P��f_�Y��ɸ�"O���*�*���'L��$��=�"O�ua�i�8X�*����^=-M���"O� �e�P�a_
҇�KX��u"OX �e��:����X�a�R��"O����ظ
��q�B� z���CF"O½{�m�V5���A�@�T��"O�t�cI'9v��*H�gK�PC�"O���@�sa5i
�#�¤8�G�'!!���}j�0AO:[o�t�Q�]f!���A�⨘���TV,�P�I�|!�#c�,����_ � �&Q�O�!��&~�TC��Z���D� �!�dPG������
��3�&��5�!��U�^(v��x��)p��~�!�L�X{�iJ���<D��!QE�1I�!���mƬ�{��ց%d)�z	!�	�U�4L����M���U�S��!�dЗM̅8��	��j��	�3 !�D4@@Z'E�䚵`O��!���<j?��������DK��kV!�pW�Lʀ�֝{�:P2QiI�n!�3DB����_Td����
�C�!���M͉�I��p��É2�!���Ȭ�e�`K�(��c�
6�!��(= @�`��?|�6���@*4c!�$�6�,0�'� B��C#��qV!�	rl����3>܆�P��fU!�dE�C%<\�k��
'R�q%k�F=!�ĝ�2���Z�kƢG%�iؔ�?M:!�dM�j�"�Z�H�,��(gl�I!�� �=�7`�[����N�T$d���"O }��(�4��p:�)��c	�tj�"O�af-ðTm�|`�(:.آ� "O�t�4��-x�b(r��[�ʁ#�"O�����$0�0Řu�A�@%�e�'.��'���'q��'���'���' �m��m8VddP:�l.-�N ���'b��'���'�r�'r��'�b�'l�M'-efb9���&Cd�%Y��'���'��'>��'P��'nZ�MG/
*\����JʤN\�<���ϕ�?����?1���?���?!���?����?��+�
��ӧ� &ZL1 dN	�?����?����?���?!��?Q��?��NM��Ų�ȣ � (� 
�?����?����?y��?���?���?�1������S.[�|����?���?���?����?��?I���?q��H.ZA�EI�N�H>��b���?Y��?Q��?Q��?����?����?)��N�m�"�'��?C%�a;1J���?!��?���?����?9��?i���?Q�d]�I���6�,�Up0�(�?a��?���?I���?y��?!��?��	V}�ųŇ�UZ4�3��H��?����?����?��?���?a���?��j�d:tH�N� - �'��?���?9���?���?���?Q��?��&���ҢC7c!��S��?)���?����?���?!��hb��'rH	69|�A��R#8�4m{p�R.' �ʓ�?�,O1��� �MӰ�S�x��a6J�&]OƸRì�?u�2��'��6m-�i>��|�JշF��s��ŵ�\:С��(�I�"��jӎ�����韞�O��Qcq��-]$�	�.�{�~��y��'��Q�O�$���U�]�p�i�eK�T �c�u��M����=�;�MϻYb���$�@�!(���-
%d!�Ț���?��'��)�S�0l�%m��<Q1ϔ���Bt"� ݤ�1M��<��'& �d�!�hO�i�O��ì\�����E��g�,LA�8O�˓��Vq��B����'�`���^W�*2#T�wK�(kc���X}��'b2O�SP^`$���+V�`ɲ� /���?Q��^�%�|R���O�%a�A$X&I�#*�]� *=+��D,O�ʓ�?E��'�X���Кr��0��mv���'�t7��V���&�MC��O��{��B?^��$kƃ']�čQ�'��'u�lT�撟�ͧpb�d�n�p��"�٤V���
B���u$�������'���')��'2�c�*U�~�` �'J���R�p�4�p� ��?!�����<������i�MˁS�
5��h�3`(�I�M;�i2O1��uY��H��ѥ�.�Z���"iy@&g��Q��KW|��ui�GT)dt�n�q�	���$ ��3-��h1Ȗ�O^�`�$�O���O��4�<�v0���Z$2��cݸ%��eU _2��y��R�F��{Ӷ�D�O��o�
�M���oK`*���5�,8�k�oa�١G�.�M{�'�`�-;˚�4�~��$>���;H
��롤���Љ�ւ@�'�����?���?!���?����O��,*%RH���Aß9bvU��'�B�'u�7M_�|\˓;ƛ֗|��� hd��5J�~X�a�)��'�������3sp�V��<� H�^���14`M�|$�ӵ�@7!�&q��Ox�O�ʓ�?����?��z2��4��+"`�Ԯ�#e���?�����d�𦩁VC쟔�	�<�O����M���S�i�ijFDP�O�)�'
��'
ɧ�I[=H���!�E��!�$�MEzL�Ճ�^
#�6LGy�O�@���Q�����
$:����1	\�H���?	���?��S�'��d����+�x��m�#Gw������]����,aܴ��'t��?��L�#�����R�.�F��(ߵ�?)�/�䬪޴���Ȧ�,��O+�ɪA^�����d�b\�i����`yb�'"��'���'�U>!A �� �`�QkX�.�E�f�D �MS�P��?y���?YJ~�7қ�wLzA��%
*6���/ƿ,��(����Oz7MDf�)��d1�6Mn�d*�&JP4�0mP��Y�d��a�o@CiB�J_�ICy�O�rd�,��Y�\%-@]-S#����?a��?y+O%o�~��-�'2g��h���yƩ��--ƥ��e��fu�OȄ�'@�6��ۦ�O<�r�2j݀�Q�)s��
P��{~R�ń y����1טO=
e�	3WPa���y���"H���c�V5��'���'B�sޡ�b�9[�0=�pFX,,�`�a�ȟ�Rܴ+
�p+O.xm�k�Ӽ[V��;!D|h���ۼqB\@��M�<d�iX�7mЦ)��bЦ��'�Ԃ����?�p'Ŕe]0���X�jK��B
�S�'O�i>�������I������Po���-P�<8�s@Ւ-n�'�6��:�����Oh��=�9O� E�V8D(EC0�
�V��eK'b�K}�z�h�lڷ��Ş�xqE���蓠�6>5z��2jKaP ��'yj���ןhz��|�T����[�g�ꤹ᧙�]��Hs@��T��ϟ��I��Sqy��pӂݘ3A�O�����	f�^`�5�ʯfZ>��6O֙lZJ�j$��=�M��i]b7-@�$��Y �S":�PCBDC.Bqf���l����ɇ\�`���Oq��� *�x@��@FL���-IQ=,��g5O�$�O��$�Od�D�O�?%��l��=0d����>"x�8�.��$�I؟X
�45gha�OR�7�2���y�hR��M �*A�a�80$����¦�'H�x�nZP~�����AS����8H׍�?:/cA��؟h!!�|b]��S��$����40�B�e��Xa��)A�舳�-�ʟ��I\y�JqӦ����O���O�˧$|�}Ӆ&B�TD��2�c_�iH4�'������o�d�%��'���b���$��@՟�U�1Ȟ�M$$0&Am~�O�`��1Z��'ڲ�q�m5c"��bMP�5��K��'�"�'�R�O��ɤ�M��;I�9*�MI58z͋B�J�W�z��,O��l�T�38�ɋ�M��lA4jp1�s��rLa�A)�#ΛFm�H���n�2�h0 3��d�Oƪ��1BX�jG��bq΁�zF4�S�''���l������ş���E��Ϛ���M�1u��f艘Ȁ6��;3��D�O�$1�	�Or5mz�%`�hL|n:Q� ���`��)��BD*�M˥�i\$O1�J���mk���	>1�䤲���z�`�a�T1J�\�	+{� ��'�'�J'�������'���2c�$J�@����T	JC.���'��'�V�p�޴.�����?���+��L��I2N���a�JCa�`��k�>���?qI>��F�>�Q�k�a
V����D~�F�#A� �iQ���4��'����o]\0�ʂ/1
��Ӣ����'���'�)�'�?�#K�nKZ���FP?Y,��zRō�?�t�iQ���w�'Ld�(���8mƅ�Ȇ<W��@���4hpZ�I����ϟ|�Nܦ��'>P$9r,]��I�*������ͺ�Y��W������O����O���O���Y�V̋�����H��Vm,ʓw��R!(��''2���'�M��:y����JJ�$S���C�>����?�J>�|��e&K� ULŶT`ВC�Q�XZ��4!���"�2��r�OB�OJ˓�|��N�(��P���S�jx����?����?q��|z,O<n��Oo>��	�3�$���E����̘.&�FH����M��R(�>��iz�6MC٦1◌R�j�fa����;�� ���$&#41n�|~bD7���t�'ǿS`FT�/�"q���ʁq��D�wl�<���?Q���?������O�s��,�d=٦n�')�lA���<��x���d�$���QӦ�'�,)VC	���S�bMY���˳Aڐ���?���|ҏ��MS�O����J@���A�L�&�k�O�%G^�DQ��̒O���|���?1��vl`Z4c�z��Hӳ�I[M��*���?�.O��mZ�l2��������o��nۓ2/
�cc��w/pe`�`����Ap}�*bӖdoډ��S�d���e�կG>z�,ȉ$S��#pe��kjz���O�I��?�W�:�dյ<��	dԌ�� �{�`���Ov�D�O���<��i'�Y�%��UJ�ٺ��>'=��)_!剗�MӉ�>�S�i��c��]�8*��c��tD��a�~�d�oڿ?N�mj~r띖!,���r�)C+�H]B�K+a��t�"$܄����O����OX�D�O����O@�D�|B���K�d���*I��1aS.Z� #��I		(�r�'`��O���P���i�Q8��!�$�5�Ǎ&Z��&��?9ٴ ��I�<�S�?���+uP��m��<a�٦��p)��z��p�(I�<��Ǐ:�F������䓻?����t�'�mRe�1^�A�a�K(}��2�'��B�'�Dy)�'ZBlw���LF�?Q��՟p�vBWI�A�f�&�
��s�t�ɻ�Ms���y��'��6�i� �v�O |qh�;*|��f"�z���c:OD��,4&܌ a �:2����?�9�� ׺;�'vmqҫ�N��H �~4�)���'�R�'���'W�O��M@�
˳6�HM��
1x��D`�P�q�Rs��E���O���O�O��4�u�O�#[��B��+�"i���Od5n�)�M#ײi#��rñi����O���'	|k,E�e}�,�4����բ��״i`PN>�,O�i�O��D�O���O�Lz��R=ou���I��2m�7��<��iʲ|���'k��'y�Oi�ˎ�/Y�=����""�Ф&����dl�&lr�Ĭ%�b>YR27ay�pI����Hf~��Pb��&$?I!JW!"��$O�������5I�a�+�� J(8�#��>p����?���?�'��ď̦9٧��� �S�0*����c�G�b�`��ɝ�ĳ�4��'Ψ�hǛ�-x��m�u�FK�
=Bk�g�n j����e�'�Q���C�?��}���r����Ŕo��� +�k�Z���?���?���?1���O�Rt	�)^p�C��;z�j��'"�'��7M[-sq�S�M;M>���� ���jEDC�r�H�7cڡ/\�'%�7�F̦��~��ll~Z�p4LE$��H �ڲa��a�A�J�O�@�Č����4�����OJ�Շ+X��XcfI&"�t50D,�Lu���O��$V���֞,@��'��P>Uƫ۱=gDXٖj�:g��k�H.?I�]���I��'��yr��+2�=K�q�Gǎ�=��H�'��<��T(ߴN��i>�9��O��O��$��?.��\6�Y�	h@���O���OZ���O1�˓"X�&.ZNr��0��#3�Hq jZ���tW� ڴ��'?���?���}, !��X'k��������?��2Fށ��4��(C ��O��)� �)�ŀ�&�r50u�~p:���?O<˓�?9���?!��?������ a��H�e�I4FR�rf&ވ+��nZ	I�1�'����YȦ�'=l� ��#Y�(�z�i�����4��F6����p��7s����.ܺQ�΀�v�K���֊t�����km��l�INy�OQR愨` �ZU �Y���@^:5I��')B�',�	��M��H���?i���?! %�>uق�j1��'b�:#Ŕ���'X��5ۛ�*|��%�`ӔɃ
2��\���p
D��' ?��O�!`b�DP̧���DF��?Q��6Pw�ĬR�R�:�	δ)�b�'MR�'��S����fmԍ��(�B��M��!�����)�4_|�9)Oio�_�Ӽ�E`1?�\��@fU�g�p@K��<�a�iQ�6���q�%LŦ�' 1�i��?�"&EI!>��rEX��@�[Fƍ�^S�'��i>%������͟`�ɇ7"��Y'FV0�a���76.<�'D6M �eԺ���O��*���O���}�*%�Y�8�R�a'#Q}r tӜ�lZ��S�'	�]�4隈N�&��/F�x}�HSцO����'����f��ޟ\Ù|2S��cƭԓa �XRjۿ]t9"%@�X��؟������Ay�/`�̴� �O6�:���<"A�1;���t�X�B?O,�o�u��T��	П��IƟ8H�J��Ux�80 �*0j��t���b�o�p~"/Ӆ[���'�䧅��N	%=���0�W�#��t�$��<Y���?���?	���?!�����1�چ���*;t��9Y4��'D2Gg�|C6;�r����%�`��.\(<�*�j4�ɥz��kv��f����d�i>M�c]Ʀ5�'��
���q�x���0D�媃�G��������d�O��$�O����*ܤ�j ��� �ӂ�3�2���O��w ��b�n��	ß��O��DءF�>K��@��ho�ш�O���'��7m�ئɓI<�OS�-��W�Gj�aـk	]���sd��I
&q����4�"\��,Zr�O|ЂG$�'Z+\ h���k>��p�G�Ob�D�O��D�O1��ʓ;��VeJ�lm+�&�?P&&�!����I��MS��b�<�ڴ�J�)��#Tޮ2u�I�u�^�81�i��7͘�Y�6+?AƎ��Xں�I+�i <�`����<1�}*���y�^������P�������ɟT�O�6�P�AL��<#�L7u|A;��d���
�)�O���OH���D	��݃[�ԌY��v�(�`�;�`=���?aI>%?�R"ZѦ�ϓ`k�� b��5e� �����$w��!�Y�N�O�M�K>.O����O����~�T-�A$ڵ_�`����O��D�O��Ĥ<��'����?���e�I�n,_���@bD�] �(�RH�>�i�L��(�m���k�|!ty��Ɖ�;��I(f�B4�3 	9Q}t�%?��'wt���6)�p):*)p��Å )�\��I�x�I�����r�O���?fZ���VJU0`�p�`�Π��!mӂu��<��i�O�.N�lM��bѫa
�bb�� #���O��I���C�ئ]�'jٱw���?Y�V�͜2'txjR�	
��������'�I����	�H�I�����:(��4R�gj�3��vժ h���<���ivzܢf�'��'��O�����-���7�%��i��<}ל����ӂ�'�b>���c���lp`�ʻ\jL<R�e�'HO։���.?Q��ݶB���$ӝ����DS)!7Ɯx�䁹"&��*# ���O���O��4��ʓL������h�rO�;6'Z9׫�$��۶�Ʉ]�B�u�b㟬h�OH�m��M뇹iKBѻrS��9���P�v��3J����X &��R����)���:������x6�U�	箩#=O2���Oh���O��d�O��?)���٩�U9E�c2�"w�X⟄�I֟���4P�Zϧ�?QS�if�'\
��BH�9F�xj���0�,�B� �D��A���|����Mc�O� v�O@&���J\.�F����W�"�i��e�ƓO���|���?Y����г#̑=�.H��	�L`�-����?y)O�qm��N��'�2Y>;2�ˮp�H-��@_#|Hf��;?��W� �	Ѧ�O>���?ղ1�ҀuO^���OO�]�n�ˣoW9'.��C�9�v��Ef�O�� N>Q�`�4U�d���Y���-�?���?Y��?�|�(O��l�)[(���RM�(d��T�<9A @�Ɍ�M� �>q��iZ�U��E\VGDBf�c���Ч�zӬ�o��s!�Ao�a~2\#V^L0��T�)��,`��!%=��d�K�'��d�<!��?���?���?�-����WI޺,�4�0운n�$Ԡ�'P�����BџL�IƟ4'?I�I��Mϻ"��0ː"Y({X�T���db�!(���y��x���`��9y��4O�����J�T��*��m#b�9O��8@H��?�6�8���<9��?�AC�99ĴBB%�9M�����?���?Y��������W�˟���۟D��D�1�$��WkN�HQhf��
+��ß��s�ɉyF��Y4��f}��`���R���l�zۃ�:�M����&�L?1�J5��ҕV>:�(X����#6=����?����?I���h� �d^�>U�7Hޤn�Ա  �[	&H��DZʦ�����x�	�M���wc^ac��B�3c�T�j�:�'�"�'$BH�_Л֚�� � <��� �L@�.j��.�7��m�eK ���<��?����?Q��?9f�_�:�6u��
K�G`Fh*B����$���I�`ȟp�Iޟ�'?y�	��P�Kצ� I��q�5R#, Z�O���O�O1�2M�Q$���+T��]`v��"�	
X`7�Oy�kQXR��������-_Gv�7��n^P�2�H
p(���O,���O �4���������۝�|B��"��D�pkN�[2��aӮ�{�OLPmڅ�Mӡ�iI�S�g!��� ����h��
ѐtΛ6�����N�i����i��y�4�	:j�rhs�gZ!zPk�<O��$�O ���O���O��?�J��B������(6�X�������Iʟ���42���O�7m=��F�;"H��CЃ"r�l�V	�j�z<&�`�	˦�D���l�L~��0�L�c�Y!���зcܭV�(��� KƟ�R�|�P��ڟl��ןL8�H/�3 �_"5�я�џ���iyB,a����<�����)U$aeL�I�:Ւ�2ԡ��A��2���ꦥ��4`����߁9i�Z�"�p�a9��?H��8�&�*�|�����Ӑ^Uv�ɈL�=�ĭ �8��d�c-�d��ҟ�������)�ny��t�l1S&�T�`����#)���c�D�YSF�D�O��n�^�a��ަ��C�\r	�>3�<����J��?yٴ=�.hڴ����� ���n�ʓ|�U�N�_�V�j#`�������O*���O��D�O���|
�%�1I��K�)C���L!4d���K+E2�'�"��$�'��7=�v9��$3,���B�bÔuӔA��M�5�'����O��DcE�i+�d�K��P����r��`�*W����%D�y��e���O�ʓ�?�s�:H Rf�q�� Jנ�p%hA��?1���?!-Ojdm��8U�'��a� \���+!އa*�Z#���O̕'��'[�'���	�a�t�e�K�7����O��9c��gl
p�A�4��@��?�A��O�����+��]� nFތib
�O���O��d�O�}λ�2����E�R:�Xه�ʎ3ݞ�r�N�֧E�+�R�':`7�3�i��aS�?[N��r��kĜu�hj���۴3\���z�
-2@'x��Ծ8#�������3�ڙ�ȚNK�	�D�R�����4�����Od���O*�d�I�>ۆ$\�L��a��
>5��T��M�'Pb�'����'J�����"hqm�kH�KQ'�>����yR�x�O���Oм8b �8�:D.��=X"��瘹7��b!����d�~��$+��F��O��&�~�B��D� 0�bU�t~����?����?���|.ODHlZ"c�r ��6'���T�Y0:��kT$!7�:�	��MK��g�>���yҶi�Z��O�&ɴt�qȵ\"�a�cj
 G�Ɛ���&f�'W(��I`�����kJ$}�`��1���?�v!�Iy�@���|����������J󃌆e���u#���"䂧+M��?A���?�2�i�D@�O�2�fӤ�O�Ȃ�O54�LM�� �����(a��l�	��M���J�b)�MK�O��R��-3 �J��q� 	�&jTA����!���O���?���?a��R<u�'�X�p�ԍ�*U�2@Vi����?�/OX�m�3ظ�������IX���I�m1B�qei
Y(A���7��$UH}�Os�6<mZ���S�D�S#VB� �K�%#X`����c�8�`��*r�dQ�O�)$�?i�@$��˼Cl�̺'�δO���&�X5F�(�d�Oz���O���)�<��i{�2���TgZ,�p�S�%St��΁�c�R�'�<7�*��&��dæ�Z��P�>���Z ��(b��z1,���Mk��i�`+0�i�	�?~�z��Ov�'?����^�AC�Gn�':������O��d�O����O��D�|�tO��T}�G!�D&�0Re�J�o��66O���'����'��6=�.���X�C_v%x���%�-ٔ��ʦ� ٴY���O�� ױix�d�>(Oz1#g��tĪ�Y���11�|r|�p��P��Ot��|����01�R����H�`	�;4��Ep��?���?�+Ovdmڔk&��Iߟ���3.W����
׿Y�}�b�۳MV  �?��Y�,�ش/-�vi*�䆼$Wz�B2��4w��M��L��`��ɂiu�5���:K˜c>]��'����I$!���gB�B�zL��G(2���������I��|��a��y�/.e��X`i@�l���I� _�BjӼ�J0�<6�i,�O��W�N�C��)oQ�M��o����ߦ�K���McĢܹ�M��OU��S��*�O�?/��l���*c�V|F.�9w��OP��?!��?���?���&��(���N�p��v��5B��*O�0mZ; 7����֟��IF�֟��
*5Xh�o�!D�Y!�f�'��^r�֤�OtO���D�ie>�
�d���P(�R�@7�8D�fb�e�˓-��� %�O�-�L>�(OB�e�	ҍ��c��L�Q����矬�����	ß�S\y§t�x�T�tޡ��^�5��i%�T΀%�%;O��nZ@���	̟ �Iꦭ���N3a����2,S�oNf9{��Gt{� lZA~�왈a2��-"4�Oi��ġ*��<Kæ��L�%���yR�'A��'��'����
�p����j
&#���P�@+��D�O���Q��U"�GUy�Ne�
�OȔi�)��8�L�)�A�2�"�����Y��M�@����nD
V������)��3� ��w�?.��E�d���V�>ŉ&͚0�?A��:���<�'�?���?9 '�!1r`hlA:���`�O6�?i���ċ�	����۟ ��̟P�O� ��F���ӈ���t}��OJ��']p7����O<�O76��U��v�>e"i�%cLY�c�aA��4��(�� �̒O����>A�#��19�B)(3��OX���O����O1��ʓY��O�=�0��E�F�;!&��em)C���*�_�H��4��'-&��M� �z!��C�	����yZ����a��od��Y�a�|Ӿ�|#�틆I����O�Zc���p��@x�`�:By
�h�'~�Iß����	����IV���3e�4�I�#���@�syB6-ջZ!6�D�O���&�i�O��nz����j
0mb �(�Vy�W��%�McS�'���t�O���iWBW�V:O�И�F>���Q�l�
/wh�y&>OnD0bh�?�r�?�$�<����?�pD�1|�%8�#�/�0��gC+�?����?�����Цm�1�̟ ����"�;pp]SW��*����w�m��$���	�M���i�Oz��3�U�&&��2ª
{�U*��D�%������.�S��RϟL���oˠt��d����e��GM�����T���� G�D�'��@�2��=&���cD�N�v[�ٱ1�'��6-�V���PE���4�n�+sG8Z�-Yp!�u�8�w�O6�i��m�l٨�m�M~��\�Z��S�;�*��Q�=Ю�@���/,�n1��|�Q��Sٟ���ӟ�������X��Ʀ�v���Myy��}�\�{���O���OH����ܸ:��vƈ]}<�w�C�����'�D6�ӦU�H<�|���o���bCY_(Й��ԋp�܌�Ѐ_~bߏ�&���>s�'��I�9�*a�q!F�fEz���$�:���ʟ\�I��i>!�'�f6M��w�L�Ю+�����+I(v �jV&V�8�����=�?��^���ݴ(���(w�X�!$�8m¥iqEضv0�:%��(}6�%?�Њ��`��'����1  ��<m��3��[�L(��r1o|�����L�	��x�Iޟ��bT�U %��5z�I˛q��(�h�1�?y��?A��i�x�:�ONAs�T�O©9��݈g���Co�E,��]��Ovo���?���Y�B�lZm~2NM�'�NŹR$�A�g� �>��4��ޟh��|Z���I˟8����Z5���r�� �㭛�Pa2,p��\�����fy"Dr�Rt��$�<����Iׂi�s�ɱ~� �U����ɜ����Ǧ)k����S�A�
�0�7/��hZ6ܲ����o�� H:A<���$Q��Ӣ0�b
�V�	�!R��)�$Z!�����1o�y�	������<�)�ay��`Ә0���Pz1��l��I$5���	-e�V���O~Qn�`�@��I��W�0i���VxrQF���?	�4g4\�!ߴ��DK�)rde��'<�8�H���-�m��YV�T�B��IΓ��D�O~�$�O��d�O����|r�扳Z'�| A�Ěiʮ4hch�#T�V��%�'a��'R7=�D=)e�3L��EÝd��i�F�O���4��	Z��66�e�������|����&x$�p�l���l�(	��.�d�<���?9$�SѢ�1'�ىb��%:7Q��?I��?Q����T����r˄���	̟��7�� 1PJ*l�%�3,�x�[��ş�Iv≐h���"`Id�U�n_�o��4���+Ĺ1�PH~r�k�O�)~�P��c�o	B8�5-Q���?q���?Y��h���d�$oDX=Ѓ��6Jz&M�%��.���̦���k�埀�		�M+��w��c	�A��)m�	9�r�J`<O,���Ot������6M$?�uB���S�y�vL�.	�  �'v�P$��'��'U�'�r�'�����J/�Nmi�F0K�v�Z����4��]/O��4�I�O
|�W8;mX�r��E�tTc�KGg}��'���|��to��i��I���#�b�a� �(Ԙ��ihfʓYp� P!���%��'SL��A �)�@Ekf ?���C�'m��'U�����T�p�ڴZL����wDm�oG4+�~���dxL�8k���$G|}��i�`9mZ9�M���\^�P��BP=vlƼ�禋9R��c۴����t�r���'��O"��֪��Ta���t��t�r�8�y��'�b�'���'����W0D*q�կ�4آ,s�!R�p�x���O��D����k�K�oy�z�0�OL��*R|���7�B�L�k���z≽�M3����T��C^�&���Hg T�t݄0���Nč��
� �fyjw�'8�$�p���t�'���'�n�r��[,)�B v���d�'��P���4O7P����?a����	D9sN`�kR�'��x5LD�Td�	���d�O�7�A�|��ʛd�`u1�-��$
pY���;0����ɋ�x�
���l՟D���|B/JB4������L��+؈i�B�'J��'����X��j�450J�"���th2�Ї:Ĵ,S�� �?���j+���D]J}��'���@+/%�֌q���=����e�'�-)K������OI)5g�ɽ<��)�=Q��lS���KB��<9-O���O���O����O��'��-��/O�7s�}��?���M+�
�?����?	H~�� ���wB�Y-�f|����˻(����$�'���|��$��%T��=O� d0�f�	d�����5LjL2v8O��@4M�8�~|rQ���	���V��]���y�,:t���5�����	ϟ��Oy��p��U+�Oz���O l��� �jF@�����")��P�O �	����O���?�$J�9�L貢�;%�~,\��A�O�S�.cض6-AF�\���O�����H�9�K����A���O����O��Oң}��.|2Tab�I |"53b��9H_`Ձ�� ����2fE"�'c�6� �i�ݪrj�y������o�p��q�8�ߴh#���{Ӏ��F�m������xe���f����7;�*���ͮK$��#ʛ��䓏�4�^�D�O����O2�Dک,ײ]	��'c�>����C�!+��>��v/:��'�����'p���n�dh���3�EWb�$���>Aa�i�\6MU�)�s1g>�&T
�oY�h�(��3�߬�r��J*?��^?T�������$�f� :�k[�c�P�)�Iu�����O��$�O��4���@�F.	�Y
RS��� �0�@��	�y�h`���
�O�hl�?�Mk'�iY��+s�E�]�xH��+�}(�Fٻj�曟�����k����i��(0�!IӼǒ�a�CĆL�dy��:O6���O����O����O �?����^-�7�PC��k�O������T�ݴj�J�'�?��i�'�Zz���'2�9k�H�,�،��5�	��Mp��|2U	���Mc�O����#P.�����o����&��#?� R�5.*�O���|���?A��(���AbĜ/�F�zJ۸/�L�0��?q(O,4n�O����	��	W�4i�d�\pB$��[KLİa����Q}MӦ�m�?��S��ȹUi8}ґ���:8xñ��e���Y�+�:tʀ`�O�)�2�?Q�d'��B�1\��q-�*->���F��>=����O|�D�O���)�<���i'h�ɖM�.t���H��^�"u��l���'��6�:�	 ����O������aI�c�*�G�,��Ģ�O���I��B7M6?!GjPL����wyB�T_ժ,��k�Nv�h�����y]������4�	���؟X�O�V��f,ܛyz!��Q�"D�i��rӔ���A�Ov�d�O�������]_��<`�)E��pcĭڢ
���ݴG���%��iK
M��6�h��y��6&�f���� sV=*��}�xcba�I��`�c�	My�Oib ��<,J	��L])t�
-��DwQ��'��'��ɜ�M�6�Z:�?y��?� }�T��f�:X��r挹��'e��S|�v�m��<$���gF�ri�xI�"(74Yp�3?�l��bަx��
Nv�'lݨ�DO6�?IWƌ��� �'呴C����'�R2�?A��?����?��9��Y�fߠ2�ƥH���4�u�v��Ol�n�{t�'��6M6�i�I��Β@������>�J�Cc�g����4s�F�oӺXh�$v�j�@2���&䟔�閤�Mx�9�`�^9>��� i|q'�������'��'���'w<���#T5���X��N*0x��V���4Gl�qJ��?������<� ����Вl�2~ �[�g��0��l���S�S>(A0$�jZ�2נ�qǠ0����Q�^�$�b.88;���OTI�O>-Op�9GgF)S�0ڔ)����P�&�O��D�O����O�)�<���i�X�p��'S�T�%]2g���b�

�6���'l�7�9�ɔ���զu�ش,c��
��Eb����^�PK�<�A'&z�� �i���q����O�q�P�.޹��e������h{垾B8�d�O��D�OJ�D�OR�d'����@�d�0>[�8� ��4�|�I�$�	!�M����ߦ&��*�M�!C�
$M�t�@a����h���Gy���Xn�D6�"?U�R���\��b�7$p��y�#?1իE*�?	�-)�ļ<�'�?Q���?��W
a��1g�)�уԅ��?����$[ئ�������I֟D�O������]<yp�aG��좹c�O��'��i�ؓO�S�1Xq�K�	_��H��^hx�۠ʁ	m�fSPe!?ͧ�$��˂��W��("��m(�P��)���y���?����?	�Ş�����Rw�ĲS|�BTC��zt(R��/y�L ����j�4��'���fJ�T�)���	~ n���V!�6�����`2a����'�E�q���?�&>���V27t�yB4G4���2Oh˓�?���?����?���;>ժ������4�/.�HoZ(�������	A�s�<����+�鑤a���p��1
�bek����B�2�iFܓO�O:G�i���!�����͕}\��H�æ��O]��P���A�2�O���|��j�<a�$@Hp|饏�
�0�����?Q��?�)O$��	< ^���O��`��|pw��.D����@ܛq)�tk�O|��}��$��3f�	t�<���#�&�9��??a#�@�yr��#3B�/��'}q�����?�R�N	t!\)6Ҿ! du��(���?Y���?���?ы�ik>=h���p^��s�� ��,jB�O@1oZ:l���	ܟ�kش���y�@V�l
m�dɻtܼkĂ��yp�,%��ۦ�
�%_����'}�Tkd��?m
ч	%cD�0	G!�;����s��e4�'��I͟d�	ϟx��˟����<�i�f��+B4
�k�J�V�`�'�p7홞,T��d�O���5�I�O&�S�\ ����Y]��Rp�EO}��v� �Io�)�xl�� ��E��&׾x2�@G:!v�MI6�U�]e�����1e�Ob�!I>/OJ	��
�X8 ����K���:3��OV���O�$�O�<i"�i	PUa�'�]�PA�>����]�B[ ���'!P7�7����$����
�4Ǜ���cV��b
AtZ���HU�
���i���"U�F@ZR�O�q���Xt�����lj�XI )܊ry��O����OB��O��D6���T�����T�t��fl�5{�D�	؟��Ɋ�M{�#A]��du�B�O&�0.��e'>dz�$ VE��i�M�����lz>Y{4'J��-�'ht
'�E<h*PbvK�
mF�+���3\���'f��Q�앧���'���'dJ,�Z?9:qh��=����',rP��i�4=�x���?Y�����10|��h�4\��U*raY2v��	���d���ڴ ]�����bAD yS&*G��R��
#_�2����;@)a�b����v�R(�;P�'���e�9O)� j�D��C	B�2�'2�'D����D�'�Bݑ5P�ȫ�4H�tH�	�I}P��dG�\��@F�
�?���?�M>�������%�2��,&��ڣ�E�YÜ|	`�0�M��ic�1 �i�$�O�l��g�P-�̺攟4�&D�IF �M�/x̃CMo���'��'Eb�'	2�'��ӽL%��H�"
�l������7��*ݴ,�@���?���䧶?aѶ�yGG���,a��Ҭ�'FA�t��$l�|�&�����(�nr���ɺ}Y�����E*LӀE+ӣ=A*�I�:@\��D�'7��'�����$�'�0�Z�)�.c��s�Z�]Q2D�'�B�'wbQ����4~�=���?��7��+5��I0٪��_�]i���>)�ib�6��H≥P������Ty���T$xK(�#p�J�W�1��T�|�5�O�T���`��=b���#z$�3�N+2]����?���?��h����M�8�r!AY��@	Q�G���$���Ѕ���I��M���w�l�K�>/X��X��t�'P�6��æ�#�4?b����4���193�-���5V�
A��hP���B�	˸�*�B%�d�<ͧ�?A��?���?1�%�1y@��ir�Ӯ4��y���H�������������I��(%?�I�-I�}�!�u�`	+���^�ɪO<�o��Mc��x����k�"��EŘ0m�B�5��V�9U$�)����3N�:��V���OD˓gfx5	r@��,Q���rʃ2~����ɇ�M�v�+�?��G�FfKJ6>�^���*�;-:��/�M��Ȭ>i���?����*��W$_�hp��@�Y*,��U$�3�M��Od���
ĩ��d���w���3��@��'\�]Bl��'��R�R &��Q�
p,�r͋9n0�I�q޴7��u�O�6�,�$�'ws��R�DÉP�r-K�bU�|�6�Or�d�O�)�32�7-0?���՜S~����j��$�6,�@��6	&����� $�̖'�O^�*�K�6�^�c�F �*w�Ɂ�M� �����O��'�����,
$)q��b���d����'m�ꓤ?1���S����*BHK������\%,
�\��!��%�<�'t�	~�I�d�2ȉ�bY{�T�@��G�BC�	��M{0�B�*5Tő�!�2�N ^X\��o��Ċ�1�?IZ�\���و�BA��V��,���Y�qC�)���`+�����9�'�P����bJ-O�*`-�'mʍ8Rd��$��9q?O����=���x�L�:��Ì�@
���UP�����[b�Iß����yG)��m1@p��c^0e�($��"5_��'?ɧ�O��}�R�i��d܄���U/Z�@�h�r��Xp��*�'a�'��	؟���6Z@�0�`E�f��/�Ow~���ǟ��	Ɵ��'W�6M�~�6���O��$�/:V ȃ��J18��Yp�KL#G���ty,O���xӆQ$�\�f-N���`�D�Ό4.�:��"?�t	
-�|�r�U�')��$�?)DgJx� � )L].|"��ŏ�?!���?q��?���9� ��m|~��
�9�y�ׂ�O��mZ�
�`��	����4���|λoY���"�27T6`�e[��ϓ�?q���?���*�M��O�س�����f��V�
�*�kZZ>h����l$�';�Iɟ��	⟰�	ڟ��I�R�T��ŋ?B!$	e��x���'�p7-E=���?�O~�]X��K�a�/����T[�Q�U��Iȟ�&�b>eP��Zke��O��o.ҍP�Y��|4o����D��2�1��'X�'��I�60�9q���h����%'�N��	џ�������i>��'K�7m�9l&��D�&�Շ#
' ^��a��.r�p��*:�V�|�Odp��?���?a'��Q�� ��+JV�A�c�WOZt��4��$�5n�i�Ol�O&'�*U�$q3��8N0{d:�y��'�"�'Yr�'���)P�B^qX%f��=0�����?�5�i�����O��r�p�O���'�}��q ͂K�4Ey�8��O4�4��Dswӌ�c�&�鐺��Ql�8&���� ZO1@��OT�Oʓ�?��?��!j����Z&���i�h�`Y����?q)O0�o�Z�1�'�B]>�1��ЎED�i�0�ڤ-�0`�G,b��������O&�D&��?� ��H��Ϧi�9��F5(�8��a�
�4F�!U�cӞᕧ�$h?�I>iUB,�F(��&�2 (B|��]&�?!��?	��?�|�*O�elZ�=��(2��T�X����U�W�u�ƫ���I�M#M>ͧ8��Iן�Hg�I'8��xC`�ݻk4\��.�ٟ|�I�J�@��F�=?���e	��cy"[!�YP���x�P��@\��yQ���IğX�I��I؟��O_�H�W�\4
�������+^1�3_�Mk�_����O���.�$����2�N؃���!j�<3aBېY	�-���('�b>]S3��Y	�	�HG^)���,G��aU/�/*W��ɢK�`�2�O�O���?i�D1D���F �A������]�p�������?����?�.O�LmT8d��	�����1�0c�Ȃ�G�����&��?)�Q��s�4=��f#8񤇟hvŁ���<.e��+��/�Ɍy��dy����x3�b>	YW�''����V� c��²L�-�\�I��,��ɟ���O�O��C11M��C�S�BHP��'���wӂuxgJ�O���TǦq�?ͻM�@��
SZ���4gQ�<����+��F�|�6�m�C? `z�8?��G:0��������4:g)�j���E�L|	�H>�-O���O����Of���O�x0gCN�zA\��ۦo�8�ŭ<9��i66b �'o��'��Om2�G�zj&II3���Np" �GI�5*�~���eb�8�&�b>�p���=7�ԭ#B /�&;7�'85*�{sm5?v��Ct~�d�*����D�G����@^�B�Y q�T�i4���O��D�O"�4�D˓A*��'Y"92�Wrt<آ��$� �����y"gӐ�V�<Q��M���i�
���!U�|��܈`țsh؈`�ؤEP%��O���[ ���d�w4�qBtb��I%jmB�G'�N�Y�'&��'NR�'��'�<�D�H�� �3�	�8[Q
�O���O�`lZ�gqH��P�4��{�VuK`��;˺�@��5!�����x�h`Ӝ�lz>�ta�e]��y�>t�f���re1�ډ(�-�P�a���U�����4�����O���]-���� �c�\̊��4����O"�2���PM"�'"�U>yv�J�#G�y�C� WM�( �8?	�Y� �I��(J>�O�>A3+�p�H� q����|鱖�c�N�$�Ĉ��4��x��a,�O�d����'�����ٍb2~(�d�O0���O����O1���e�F*��v� BpgJ�Z� �#H�$��aa�Q�Xz�4��'�Z�"���8$2��eM_��@D�n�6MGæ�r��rr��l�+�f����O����d&�;�J��SC�?q��Þ'd�	͟������	����Ib��(<&�P5�Ȩ<�L�6e�#Ɗ6��$6� ���O���1���Oؤoz��*�Ɏ%{�,:�߾RNrɨ����M�C�i��O1��|15lt��$@�0�s�>b� L��Ɍ�*��� �fw��s��S�ΒO���|Z������-^��`9:�I	���Z���?)��?q)O��oZ-e���	ʟ���f� �uH�@z��c���1W���?��Z������sK<��LʒJ�nY�dc�y��㴥�k~R��1��AqeIK��O��i�Iw�ܑ%`�Y�#K� ��D
�@Cr��'���'R�s���!��Y!���n�����O�0��4 �qi���?q�iO�O�Ή�r���j�dX�H���d���-�ٴD5����NE^��O���|��S�a��X�Ӄ�-�5�T��%��EQ��|rV��ȟ��	ޟ��I���`p�@�g'��d�"m���h�IFy�d�vh����<����'�?y!�N�Ҋ��Ԃ�f�R�)��  �˟�oZ3��S�81���B�C�|��h�/K8���A(+/<��]�U9���OPLiL>-On�B�e�[�BE� ���t�8�,�Op���O��$�O�i�<��i9�[&�'��<�$̔�9�'.+�Y�'�Al�⟸ �O��d�O���Z�l�tiR�Iؒ3��U���H�UM>��`��&��I�n���ݟ����R��u�b��$j��U駡��n3���O��d�O����O��$9�S�F��P��a�'��)˔�8�a�'��t���8�.�$Ʀ&�T�uNº?���A��]>59nd����e�I���i>�Pf-ٝt/X�J�NI�W@O><rU����m��D���هw���G�zy��'���'�ҏ�?n$`g,�?n� 5�L�.�"�'��I"�M�Lډ�?mf��$�|*�]�J`٤ D3Xr��#@b~B
�>����?�L>���M�sL�6��Z%cǍB���D)�:$�ؒ�*uz�i>���Of�O���$O��v0	T�̯>�i���O[m�Ɵ��	�b>�'6�6�Z)DǼ���^�p;�і{�< el�O��d�5�?�!\���ɬ��ˣ��&�F%�P�l�L�������/Q�
�B�{yԠ��ĳ?��'�de����;;ب8@�J4�|��'�I� �I�������0��w�4��e����倗>�Bh��J-
6��B����O��$)���O�]mz�IBɆF�
�{��̧L���Ċ�����z�)�S)G����b�$��ԜTDi�G�x��@���h��IE�В��$+�ĩ<����?!��1-����� E9D�	�7���?��?A����$���2U�C۟��	�hh2��^��p��0c�*a�n�D��3P�	ޟ��	p�)� (���̔�4Bx����$�5�g�����ƤXw�QbV�W� Xs���O �(wNҊr_�AQ�٤�r�t��O����O���O��}���<�F�@�kͫn'�J��3p�y�����֠Q6Q,��M��w�8���D|f�04ʖd�2�'�b�'�r�ča�:���O�Aِl&���@�T�����T�3������R��'����$�	Ɵ��IƟL�I�j���Xp* ��Q�K�(
�P��'��6�	I�N���O`�$4���O� s��~Hѳ(�
��aI�r}��'�r�|��T!�)�>)�%f(&v���ƞmK@�cɓ�x*�	<;�iq@�OƒO�ʓ��a�F�W35 ��d�~!�M��?!���?���|b.O��mډEȤ��Ɏ)���yCi��g!���rm.���	��MC���>���?�;�B��dG+R���+ʬ�Z!L�:Hv��'V�YЅ�RIbO~����F��@
\"������(>�ϓ��?Ї���Y�$1baL&�����O
umڎd56�'*I�֘|�ë8�����Z�M��2� � O�'�������77G����O�`x��37��	�M����mk�͗M�.9S�'��'��h��9E� ���I!j���td�7�Fx�eaӖ�c�<����i��h>��W
N1>VV��$��$cE�ɓ����O���3��~��B�?��H�KA6+�({��'^nD�۲fE~��D����O�[?�N>����jl�(��ގ}�H��ՄR��?���?����?�|�.O�oZ2
/� Ӧ/WsM~�!��_�g�V��5�J��	�M+����>���2v�] d-G�x�8�AŞ=S��@*��?)��1U���'���	V�Br/OƔ�� )�$l�5*�^�B��5O���?)��?����?����I��d�u ҃e���� :����Ld�p�B�#�Or�$�O���D�ئ�]<�n�0��,$�0��:H$�	ޟ�&�b>�1N<:���2rL��HĊu��PC@���F] 牬~�D�Pg�O��O~��?��d5�a�LF�/xP�舚��(���?����?�*O���	�y"���O�( �by9aU`�z13��:��$P�O�}m�:�?iN<!�G@�6!Z�C��E�:�d5�M�x~�f��&}�a��&Q,�Ot�I��$Qer��z���'mΤK|�h�Ê�I��'�b�'��ퟬ0�!��a���2���0YN~��0�ȟx�ߴlqƑ:��?�@�i��O�ʤB���R͆2�~U��!��l�DP���Y��M�e.��%�
��'�(��0�Z�?=��!VG�ҁ(�=m��J �ܜ/V�'n��՟@���L��֟���%�tY�!3o���4�A ^VL@�'ʹ6��}�l�*���O��󄜞RP��o+��eHsO i����'3d6mƟ�$�b>�Q&ˤ{a��[�����`�]�#x=����iy"��w���I�F��'�ɷAF|k�e�.T�.)(#����ڌ�����i�n����~y�'k�,���f�O@kP��<���*')-7�J���#�O0�m�W��Sh�I��M+��'��L�1e �u �F_Y��QC��@�����X������i���F����.�.��]�'�[ ��%�V�A��$�O����O����O��$2�S�^�5ѵjR,��)1��V�EhR$�	ҟ��	�M������Ǧ$�X��@N'�t��Р .�K��%�ēa ���O�4�P�Y���O(]�!Ǟ�%n��ڝob�5P��՛P&�E��2�O���?����?	������GD�=�H!vk��H:���?a+O�������D�O���|GOI����J�$��`uZc~�n�>a���yR�xʟn��@��w��5�p�ϐG޵ 4�F4���#��fn��|�&C�O6��K>	�e��B�j���+k[�h����?Q��?9���?�|r/OЌm��H^<I��_�C5xxa5��#�6)Ia��ҟh���M��R��>Q��i���QI�D�3Q�&P4���D��O&6M?S�\���H��*�G��$	_y�J\�E�	ct�}��!�i-�yRQ���	��	П8�Iʟ@�O�~��񃀉kq*���A�;.�i�np��p�bM�<i�����?�Q��y�X:{�r�!�/��~��n��%.�o��M�7�x��D��(*��,y�'�J	�%EL�5l���N�R5|	A�'W�X����)E�|RW�����JR'gOr��VAN$iࠆ���� ��Cy�H~��	;3g�O�$�O�J�S�%\�2d��N�@<�a�0�ɇ����צ9�ݴq��'�L1�ɝqK�ఀ���F'X��O��ea�1�
�x!��Q��?)!��O�B��CJ�U{%��-#���5��O����O:�d�O��}"��v������;�v��vAE�&N8��j0��Q~���'4�6m:�iލ�#��.�%�[*X�(X��������OT7�¦�pC �?��,�`� ��0P�l�7tjHY�ŋ�T�z���a����4�|���O����O��d�'E��D�3'��Z�H��w*�j��\�F�F S���'q2���'�xd��:l�9j����S��PB0j�>Aa�i��6-X_�)�S* �,��!��q��$�,N'��4 b�1HJ�L8
�p$�O��hJ>�(O�h�1K��*u�!$�95Nq�(�O>�$�O�d�O�i�<	2�i3��
��'#�d�U"E��p�� �D���)�'V6�6�����������۴g�� ؀�IWr�s�����=rA)�>Q!��� {T�R�1���	��ʔ"���0AxT\`���%�2$��5O^���O ���OP�D�O��?�d�7?�Z�8�ՐZ�)�T���d��ϟ �4�Nͧ�?YP�i
�'n؊g�ĩQ �"en�)�djb!��L�i���|�φ�;�F��'k���M�64@yh�)=�H=��؁�q�	�v��'��i>I��؟d�	�lt��Dk%t6TP��^�#�P����d�'�6-�3��˓�?�*���{�GM
i"R��s�U�v��5��X
�O6�lZ�M��xʟ
�*�J�'!H�T��!x�mB&@/?�f�	4��DD�i>��c�'��T'���e.��Vh�1$�O�V�kcO�֟��Iҟ����b>��'(7-��A���9,�-����%�Q3.��̬<a&�i��O���'I6�D�N�DU�B��WI��y�O;�Mn���Msw��m}ޥ�'�.4#AL�?���&m�󦓅PiSB: j��57O2˓�?q��?��?���3G�ʡ2���:i6)�,S'�u��i�bQ�5�'���'���y��d���\�[��1�a��P۬q���lU��n��M[D�x��$���m�`��'W8U �F��Xl�G�н*�ϓb1Z�pi�O݃H>1(O���OX��$#E�,�hjE:M;�i��O*��O�Ī<ᒴil2}+��'W2�'��8��Y9tn�zE�Zt[�d�K}y�(�l#��NV�%Zd'�kxhMڕ�[�'�L�'�𼘤j�e�5���tSٟ���'�|�C�@�0(<�JT$��Ģ)	f�'X�'��'��>��I
4\�l����bOS!J��I5�M�S����?9�j�&�4�t4��'�<^褠���b9
��=O��o�<�M�D�i"���ٷ��$�/98�3��jxB<���Д+�L	�`f��m`f����J�VK�0�.�9
�yF�<W�����%[��a8⃖�yH6�t�M�Js�9`0J�<>�DQ���m�vp�ϔ8�,B��LϊQD��$��e��2]�H���@�[�恚���4OD��A+�+B~�T�ݣP'���H��Z��C��U�5㚛/�����N��Dn֨d�=X�e�7Q$���eJ6��
όp���8Y	D����=W���M
���s���Q�l�0�&����Q�2M14�pd�s���F�,~,}�)�)dZ�8�T��v�4s�̙7-���'���'��$	3?ٳi��H*� ɛ|�[6��I�'kP�������={���"�BT@Y�b"דp���	&?F6m�O��D�O���H�	@����,�<���t0Ȁ��:�M�fku�����$�
y\�hKDH%FW��3'�)&, �nҟ��џ`�@��ē�?���~�#�)T>�]r!��uĄ�@�F���'���y��'+��'�P���!�,X�t���~Y��k�2��݆y�>&�p��۟�$��؁E-T���B��蛡{v�Z ���<)��?	���H�@�0	�M�WH e�1�N�wv(���
P�ܟP�	\��\yrC_X�2ĉ�$ĕA -�j�|��1�y��'���'J�	?��Aa�OE�����#�dI3���Z��M<���������;��	�"�6�s�슘�f��V�H�|�H��?����?y.O��a!l⓸�XY�֍�Mm�NB�-D�eP�4�?������<	�O�L��O2���/�\t��m��DU$ɘֶi���'��	h��)�I|R����G�I3��RT�W$1ٔ��%f�)S�'c剒��#<�O�H�B�k��d`2���l �<p��ٴ��#J��m���i�O���T^~�	�Gx��Wg�e�%������M�/O>�;��)���*>x�G�	 ��e���{G�7튵s�H%o������џ|���'x�귫F�X�"<{��S�\�h02�zӀa�6�)§�?qT#ޭ^8V�X"���<��,�-��V�'J�'N��5I7�D�O�d��@���(_F����ł}�83#�2���R�&b���Iʟl�	�"���y��܍	@Jl*`��8Dw]��4�?���)�'r��'sɧ5��Wk�����m �6"`� �ʠ���əsY1Od��O��$�O�*6�r|�m�DFP����A�m�,���䟰�I˟$��N�	˟ ��A��*Ï4h��cW��F��Qo�.���?����?�����<�?9����El]ҥ��5��a��*�,5��'�R�'%�'�BU�T�!�}��A荓'Z��ˤ��9��P�`���\�Iݟ��'�ց�Op�&P*�F�1H
E���c�	��H��7M�O"�O��d�<bb�d��]�}z���zʠ9!��D�Z��7��O(�d�O����"{��d�O����O���#),<I���¯)�ٲ�+��%�<�$�O0ʓ0���GxZw�$�ȡMV�04е�����1"tP޴���1lZן��	Ɵt�������`JP)K�;A�Ar��6a��=���ib�'��b��'��'�q�FђWgӼ��P�I�_^�dB��i��T���a���d�O��D蟆8�'��ɰ:c\TX��@	5�NX�DF��4B��ٴޘ �b���OR,����$�� ҉̎|3>����¦��ܟ��ɛ3W��@�O���?Y�'`r9S#g�q��8�$�j�����}�cG���'b�'5�L��|��sv��]�F0�cؿ%��7��OQ�+
H}]���\�i�͘�+�
����B��.@`q+0�>��L!�?�)O���O��<i�Ѓ閡q�'(t�F�`V	�#fm�9�^���'M�|��'L§9� 
�ǯ]�V6԰��͛�T��P�3�� ���?��?a-O�1
Q	�|�!'ԍE�)p�˗3��y.�ܦ��'�2�|�'����O�����$�|ИU� B�P8PtL�)��������쟴�'�H,�æ�~J�$�����[�Kմ�����&$6P�&�ibB�|r�'c��ݾNPqO�)��@�]�D��a"8�Sǵi��'<剪.��Q��p�d�O��IV�(��^��`
y&��$�P�����z��8���4�.o�����C64�L9S�@��M�-O2��vJL��]�I�I�?�R�OkLəG�T�#��S^~D���.=���'b���sx�OJ�>�1r�צsY�QQ�ԬG���@�"d���f.����꟨���?%y�O\�{�f�Ab-�9P2ii�	A�������iN<�d)��ӟ��@��i<��枂@6�%�7���M����?Y��|�ZYb_��'x��O�}�𫊾DPz)!���:`�lzQ�M>����?������Ծa�tՈ���
���ռic2�=9����D�O4�Ok�����j$Dh�Hj��U(f_�		�b�d��֟��	ky��Բj�3�EG�9�!iFjՁ��!j�>�)O��$0���O��d�7Ry���H�\=R���K #b����5���O����O���^���3�Fa���{���DlT�?��4�CU���I���%�ؗ'0~TaR�'X���Z��(���L�)��:�@�>��Ӗ�6�'�>l*9K|�gM];I�ָ�ڝoRp��"K�@��&�'��'��I�����_��{�<�A��9b���i�ad<6��OPʓ�?�V����i�O���k,��D�5��x�	AS�ǵt�'���'�����lW*�����E�4B��IP#b�$�x@��'��	ϟ�w/�̟���ܟ��	�?͔�uWaP#̴BU`%=��t*�5�M��?y �1����<�~bЎ�(	&�5�� ��8�$�b�ئ�Cv���t�	џH�	�?�����ȨFQn�����d5�S��\%�6xm��9~FͣgC9�)�D������C��(�QM��B� P��i���'"��� ��)�I�l�dm�8O��,=T��)������'�
��.8��O��d�O��uk
�Jy�e3tI.D����E��I͓u�,��M<ͧ�?�I>�;��	�m��'a��*u��ts��'(R�*C�'7�	����	��ؔ'������=W��qb� ,��O����O6��?�*O�͏!Y�1����"��cԁM�Š�D�<q��?�����䉶r9Χ��m���D&2]�0�d�] ��L�'&��'��''削F�Q���m�v��iG"H8	SO9+�굱�O6���O@���<�b'DSb�O�=
��5�`g�2q̉�E�m����&���<!"B�:�?�J?M��֘|�F9{!��f�����y��d�<��i��� *����OT���\�#��9�P�*�fF98�\��xB�'q��)"�i�y���%H�5�F�����q�f4p�i��.}�����4O�S�<�S����ݦt|���H���)c�*?7F��^����#��1J|I~n�o4X�N���X�)#ig��"bӜ���%F��e��䟼��?e�N<�'@�2��	"r�ǈ^?u^��i��(���'��^�'?��pz�H2t�R�z�Ċ�6�m�a��M3��?��'�H�מx�O��O��tkC�%p0����3��AZ��i��T�d��T1��9O��$�O�ЭP�*ݸǯ��7r�������q��l�<�e`N����|*���Ӻ{#��.ta�]Rp�hq� O�z����P�����O�d�O����h�NA�u���3�-O�ص���Ƕ�'��'>�'��	�$�h{g�Ԉt���q��9\�)�QG��� �'�"�'��P��RT�����I��+�N���e� 2��\���9��D�O���2�d�<q�jʸ�?�t�Q9z�Ѝj��2D(�5�ŘG�'#R_���	&eVV��O�"��y��=���N܆�0
��4��78�	����>Eb��e-?��C<cU:$Z��S�7��J���ʛv�'��V��Bw�����O��꟬UY3D@�e��ySg�F+dP��P�-�k}b�'4��'N�,�'�b�'	"ӟ�iS�w�r�ę��n�$�M[+O޹�t	�ᦡ��؟<���?�+�O뎔&Z�b��
s5���L]fڛ��'CjV��y�L�~Γ�Oqpрd �#a)z��".M ��޴q8"�A�i�"�'���OĎ���D�pUحJ7�վm{���'�!G�!o��b���	W��{���?��-A�� s�2LtM8�1M��v�'hR�'�z�)&&�>+O��$���j�C�c���0R.�A@ĩ2��>1/O���g��������֟�P�(�#d�x��ܕ&��쁐��Mk�f͎�{�T�h�'��[�l�i���BMy6��0Ç+*��>��NA��?y��?Y)Oj!9���\p�A�fN 8�b�2%�9o�8�'{�Iӟ<�'z�'LlHO�Xu��qΑ���,^�ؼ�O��$�O����O��h\��Z�6���S��ä<P�`��Dd6����i��Iӟh�'���'L���?���������D��Z$KV�S53����';��'�rV�hj�ɋ:����Ok�gt�pa�Q�<�j�!S�ſrp���'0�Iٟ����0�pe����y?� :�I6�[�$]{�j�? A4�#1�i���'��I�H�脀����$�O��)۴_lb�1��j�T���ڌu�v�'���'�B�Ν�y��')�	nz���x\��)�]�� R��̦e�'����2ed��D�Oz�d�V�ԧu���!� ё3�I���;�L��M����?�&n��<1����� �ө1��� F*�F�ط GW6m
�Ho�֟���՟��Ӽ��d�<Ѵ]X-�!��(-tu�7��).���d"�y��'�B�'����JT�1�a���� �-*G(�m��	؟�Rt����d�<����~ҁ�#nS�� O -Y����M3,O����f��?��	��x��#n�n��D��&0�@�A��0�Iaڴ�?Q�&�t7��Vy��'���֟�ز|��܉��	H�.q�uJPA���Eϓ����O�$�OH�3`�M@�� ~�Z5�*����!���4}w��jyR�'�����	��h�c�'�b����I۲���Y���pyR�'K��'��	-}�"a��Od��3���@[H A�iƦ�@�4��d�O`ʓ�?i��?��+U�<�gh�
/������
-�52�+J�?������	̟��':��XaΥ~���/���02�X)�t���a�ʄ获�M;����d�O����Of���?OR�'���c�X4L��I	�d�9K�F��۴�?!����@�\w���O[b�'��$���i�
�X'.����ڇ(i�꓀?���?Yǯ��<!���D�?)�灨�"� 0�F�'嚭��g���Mh9��i�|�'�?��'Q��	�r�m[�O�V�`�S��˕5R6m�O���I#Y��$&�$0�ӱ;9��c�-Բ,JR���l�= 7�G�L��nZǟ8��şp�����'=�@�M��}#&4�q�	)���djӂA��<O��O��?)��;a�L ��ի|`^y�rڅߴ�?q���?af�L�'@��'��Ċ;�I#0�֗ ���� ć&I�&�|B�?r����D�O����EQbFB�9=�8�"jɊCpo������G���'�|Zc���+�D[഼{��	}���Oт�5O@��?9��?	ɟx
`əa��Y���P�jQ�� �͌; n�O����O��O����OJ�/	�r�b-�R�&8u�$��e��+���D�<a���?I����	ƾ-{��A&z�@��] `!��F�J�O��d7�$�O��$-W��dG$�E1&s.� ��_y�'���'��X��{��E��ħaQ0��0J
���v�Y)��ʀ�ix��|��'y�	�y"�>�E���O��ݳ$�ݼu�@i������I󟸗'��5�b*�)�O����&RlM��GU�I ���\?AH'�4�	�����ퟬ&����L�����F�~���!'�ݦ*4�n�^ymϥq307mWo�t�'���l3?Q�7A��[&�U�j�l��#Ҧ��	���"�&�͟�&���}z��� 3�T�z��N�K���ɱY��	xP!���M����?a����x��'L�f��̪@(Wh]K�d=�+���w��O�O��?���7wԔ@���]� b����+X�;GZ�i�4�?��?����E�'B�'�����N���4LR>&��D+�2+���|�X��yʟ���O�ā�1�Р	�jE���
�⑩?��`mZڟ�������'"2�|Zc&��##  ��X����S`a(�O�h2��O���?���?q*Ofi�$�1:�@Z��S�(H��D
K"d$����̟ $����̟X�p@�꽱 ��c"�4�7�6a#n�IZy��'���'h�IdX���O[ �G�Kz �x����q�ɉM<������?���.Ȉ��u�]���<X�P�W����R]��������zy�j�J��� �V�J�R���ǉ1T@������	n�������4*��=y��,H�8�qw�
'o����]��a�I�P�':���!6�i�O�	�,d PqsU�� a*ʙ����{TX�'���I��yb�a��$���'A����EԞOk��%��u�4oyyB�ǲx6�p��'����'?��F�r���B!/�vd��/	B}b]���I]�S�S�-����1��CP�%�`���q�6M��w6l���O����O����<�O��c �ۜ^Fe�0��b��Pa�zӮ��g.�S�1O>�	�n,�E�Ր
thaäj�!pt��Pٴ�?���y�FGh)�O����PR��T��ŃKզ�Y�&I!lO�$�OB�dv<��s�CW�X�"z��O$H���o���`I\�ē�?������f	<#9�gcH�F���AQe�o}��U"��'v��'t^�LRC�){��U�Vn8�eA�Z�(�J<Y��?�N>Q���?�ebD�&�z����B6���
r�z��<���?����?)�O�ܠ0�Oތ��FƋKL�PQ.J*#��ݴ�?i���?�M>a��?At�J�C]B�l��Z'b�ru'[�f@R��/��|ꓥ?���?/On@B��J�D�'+bU��Oތ�8��.L�HD[RdӢ���O0�H��7�I��������`J 3��b�h6��Op�d�O�����D�O���rG^i��	�C� 9��;��LN�'sb�'	���b��ʘ���ͣS��Ԛ�lT��!0$ &#�f�'��g�/=��'�r�'���'yZcn�93p��+7����Š
I�dߴ�?��4����Vj�S�g�? �HD�P2զ�)�,X�3��a�i.Jls�zӴ�D�ON�����T'��/z��e"��
8�>��b�3d��(�4'$)[���Ϙ'pb��Q�
�#�ݏFmʉ#F�N-Za�6M�O����Oh%`Bk�<�.���d�����`R�hM27�۠a~8���2��'�حb�	.�i�Ov��OLR)F��`�J�4{����ئ����S�R)�N<����?�N>��~�Z��M�z������Q�c��\�'"���y��'��'��I�����OI-r��(�Tnν]XX+��ē�?	����?��*<>�IT.Y^�h�T�P��Ȑ����I̓�?a���?�-O�yRB��|�e��9��x�g�J�{]\��du�I͟�$�`�	͟�hp �>Q0��6�����P�=x(@��b�r}��'�B�'z��|�b��L|�s%�1c*�ɉgvNAPէW՛v�'u�'b�'".�s�}B�>�!Qr�N( X�$@V�A��M����?-O2훐aYM����(��3aMǋUTn�����D�)J<���?	��S�'e�i��a��)��K�C�*pCfEZ�d˛&\�| !���MC�\?E���?��OQ� Ą�?���ۥ
}��ib�'F ���I�E�������ø��q�<Q��&��0"�6��O~�d�OT�I�[�e�
�AO!-��Dk�*��(þi�Q��d$�Sɟ����(&EpKG`اI��Y3��N��M���?��7���&���O�����p�I)5����t��W��c���BK?��������r��ҳM��Ha��M�)@�ՃqDE��Ms�]o�� U���'�bP���i���G�-l�����h��/H��Ia�����t�Ġ<��?�����$^*1�L���"[�Pɰ�m��9�0 B�_}2Z���ISy"�'�R�'�� �H"a�@�B��^=�uȅJ?���?9���?����V���l�'z�6���N�4�^�У��$V�&5ldy��'��I����ӟ�B�v�d���`*�b���l�Y;�*¥����O����O,�Gw^=xER?y�I���	�
�.�*� \譢�M��M����D�O��D�O�$Q�?O^�D��x�dM��2��
�&,'�5�lt���$�O��=��a�P?����H��1W6 ;MJT)v��>+�p"�Ox���O*��ʃFD��'��?�"��T0t����3��yh��S)g�2�1��+�i��'���O]�Ӻ3�#h$L:�I��δ�!�ɦ���ğ��u�q� ��Zy�I�381 �th�J�~t M�.`�m� ]7��O�$�OR���a}2P� �!���h��*��C%U��u�ڑ�M��<�����$-�Sߟ(���H�!dȟ�P�x�hʙ�M{���?��f�=�wP�ؕ'�R�O�I��*�55��2�*�%�@�i4P�P0&n��'�?����?��
#)
ܕ�����JܝH�6�'�hBo�>�,O���<����Q���Tx�gE�r�AI�x}�E��y_���	ߟ�%?�B��>UKpS��K�:�JH@�ꐃ^��	H�O�˓�?�(O��d�O���K�>m9	¿��p!�R3p��z�<O&�D�O2�D�O��D"��a���x�®B�3�$�(&�7rQ�J�e��M���?���䓕?�-O-���iL��P����o8�!
�4��L
�O���O4�D�<�aiF�C����Ps��T1��2���7�V0X'���M#��?q���';qO��(!�&��]��U)�ZLX��i�2�'|r�'ª��q\>�'��T-�7
���D��#㤕 5�P�.O��D�<!��Ko��u�+��A�5#b�ܰ*Vnύ�M����?Ap����?��?������?��/F����^UZ�q��(.#�o����I�"U�#<q��4k3pUqF!L_��H��S��?����,��s���0=	�2�Fm3��V�"���[�<��`�5?���ԭ
�.3Y��[�0k�	S� L
Aɂ�J���.I�թre�?+9�t�U��2t�2Q^�$C�����U01�`)��DV=��՘&�>LpU�����ZLuq��X�2P@�P:%�0��a'Q!ܠ5X�� *d �#���[4:��g���Px6�Ĕnv��k�
�?���?i��Z��.�O��D|>��A(V�S[��	ďRI��\���N�8C�	I���P��͘�-A�k>����D���N�� �D�e0�� ��ph�/T�.NH@���Φ�#��9-$!4�E���@J<y6hFW�¨넅R0��[2�G7J�(H�	��TE{2���M��A�14Ԕ���bM/'!�֟pt�-;���<<���Ȅ�p1O4!�'��	D=�aB�O �]�2mb�0��+l�$1�V5^`�$�O( qi�OH�z>�I���9'�ڝ03�خ�~��'�2�Ѣ�"o^ � "O�p<I&��}��� ��K��Ӆ!/�k׃�}�����a5H �x��]��?�����d�am l��/�;M��&T�	�1O���DR�
n��0��F/�r���9�!���!۲�
Q Р�0k��~a"��̔'�~����>�����	��U����Q�KG�-�샞q�ƼP d��X<���O�`��)d�AI��ͅ0�?�O*�S�4mj��#��#�!��o��G��'�
7	Ҋ8�i��  7A�>)����'`�n���՟5H��d�)}b���?���h���� ���R �\x��נJ�<(�G"O�9rǃ(l%�1�դ�,��P�'�#=i��Ɉ!�Ȁb��x�0/��W�����@�I<M��T*aŎ����	韄�i��F�c�N=b-���@E�_t$�A�^�L���@�b>�O6�@��*2�$�E�a��e��tc�+�O6��Ɇ�и��a�H)���D�A�,Igɣr�������$ʒG��O�ў8���?np�⠅�l�ZCe=D�7e��(�jm#D$�.��kpM??!��)
/O&! #�ǰT��<�1�D�9.8��K\>����	�Oh��O��D�к���?��Oz�Iᇏہ;Zd���̆�]�D� ����x�k�&ɠ�x�E�)8������*F��@	�'Ψ��vC�3H��Dާ���@��!�?��o1t}B�N^M8��r��	o��)�ȓc��TKQ��p��(���X�dS�`�<I@�DP��l��t�I2Y=L)z�J֓x`>�kƪ	#"z`���<�`����	�|Bq�����'����^��YK�O��1��$O��� �Ĉ3m���0e*T~�1���Y:�x�C���?�N>��X�C��t�!��?D�����J�<���O'	���
�o�\�z\@b*�_<y�i�x<YӣI�_X8!B�P�"�,[�yB��&�듓?A+�������O�����0-q��;1�[I�=1�	�O,�d�*$W"����S
#�:\:�f��$UJ�O���*���Ɉ}�.��v��;F,�'����+[@x����٘*�>�PBI?�/2�X  ���U ,�LG�<kD�'�F0p���?1����OJy8$�D)7��$�p���F}����"O$�ڷfܫy��E�D䄽d2	S��'�"=��ɝ"i�)S����>\�V�M�.���'��'�H��)N�'K���y��N���8�cd�+ag �*�C7.1O�%K��'�(d`d&�/&�v!�eGZ�xM�{�� ���<����;&�p��)�="6�P� �.��'1�P��S�g�nM6T+&ܠD�!�kֵhC�I�9r@���F7w�Q:�+L���ߑ�"|"u�T�Rr*�c�I��u��c���72�+@��5�I��p�	ݟ��_w�r�'��	:*��:V&�#����1Ό@!����Onu[�/�B�6�{t�~���e�NM���'~$�G�֨E����#��Q�� �r�@�?1�Z΍�wE�C
z�3��D��ȓ`ߤ���v�9��ZB
"�I���'t�ŋ�m���O�<��	�5�L�5�F�3E(�%��O���� �|���O������'�W�+JXy:���2'�4�A�/��x�E���'[jE�w�ϭ���� #L����<�Z�	D�ɷM�x�It�˵{��HK!\�M�~B�I�( 8Z5�V�3YPc�x%�B���M3��A��0�⦭4 xٓ3��P̓UZ�h�#�iM��'��,s��0�ɯ,�|��6dI7N?V`Sb�w�^��	ן4���<���D�!+�@���*u,��P�o�a:2�Ex��A��uIJ!�ߎ{|�Id���ɾ��<�)��&.#x�[��� _,Ż��Z�;a�C�I	
��ȡ�����2U0!M������r�'�Ѱ�+U�4}�<�u듾w��J��i�B�'��n�[Hؠ��'d�'��w��!!3��:��Ų���E�<Q��i� OP-�P���_M�S=*�1��'Yl��RP�?���U)�I&�����B��	��ȇ�j�T��DU�����X�,)	ׁ�?�`y����'��"�i���'^��C��d�'_��'"��'t�T ��|@$"��F䰔btO� �4ƍ�EFe����r(�8T��p1��d^}rX���	@�t�CΙ^��q;5!̐\I�D0��şD����L�I��u��'\r�'B֙(�0f�pxD�63e��cT�z!�DD+W�,H�t`�]e,+㎗�(�4��F�y'�ؖ��h؞��5� "l���5�ٯnx�X�Q$L�R���d�O&�&���Iɟ,�?��_�K�
M��&�Hwh�`�$�]�'?H����0I"r��#�pd�%Q�c�6wfx�O|\m�Ɵ�'��*�ê>��[Q�5B��D��l�@���Z�,�i��?��b��?������n� ;B��#��h���#V�6g2��S+<�,��K�<����9%������)?� ��D��:�p�	�D�6z���b�1�@x��'�0����Uś�>)�N��$��Y��҇w6�=�� r̓�?1�S�? ���CƘ*
�D��jͩ4�Y3FOulڮXq&��$߮6D��RE,E3A���IG̓�MG�,O������v"N<A �D%�$�P"O�e�ņ(yL�����15���"OZ�r�$��a8�b���x���1"O^��s��PH���	��dF��2t"O،���^e\4\@R�ѩT1�t�"Oԙ˵B)s"&c6-��':H@�"OV`��S�eX h�Ǭ\Cx$z!"O�<b�E��3��\4��$�@"O�s'/�b|	��j՘||ȕB"OT�"�ч�$z	Ɯz�)c�"O�T�G.�k'd`Sw�;<�v�t"O�Rrc+C=P��Wf�)��u"O�a�'j ������I�6��"O�أ��, ���)]ְ�a�"O0X�H�)�(0"�b��X�.�+1"O* �H�.0�%�Uo�"P֬��"O�,�S		 d��W�ϮX�"O���0$�7/`�}r���"� �a"O�]��C�$<�1��D f�2��T"O4�$f ;S���9��o͊�"O�Qu@�)W�$�̟\M��T"O6(��mE5Q�d@���_�7O��!c"Op�m�%K�(P��W(B�y�w"Op�ǁO:䒼�"�B�����"O����ȏ,v(1��O+/�nXk"O���d�V4V����wLJ�#�Lec�"O�`���%P�� IE���X�"O�5ۂH�.m&A�e��4+�8Yɦ"O]�&���u:�ad�V�z��Qv"OhIg΍�M�:a��]'f�D�D"Od��+�K���%��
K��2"O�� v�
+/Jؘ���٢g���0b"O�p�/A��MJ􉍢~��̱�"O��Rg��
�p�@E��#'�n�$"O���� ��Xh������+y�]��"O��#�D�'��S�PE�x�a��8XD;B���t�/�g~��ԗ�tqr���6G��v@W�yB[�&4�&c��ID2�9�. �wL�e��aCn:f���)�����^�*�@Ra�L{bͅ�	b�J 鰈\�9���ɣO��]R�E�d�zi���)K��C��/�(ؤ��G���",o�zc��ӄ".k�j� �#�'TޖHB��)��M��Q�S2���a¢�ys�Plpeh��A�`g��R�,ۚ3�q�'��@3��0�^�Z�<�7�*$�j2D���[�3��+0��YN:!��͹zr�x� ��;�����$Z9򜃗�/vȉCr�4:=az�Ȅ?���s��y��C7L� �K�^P i����y�&N`�p}	�jL�fr�-!��'�v%2%-#Ed��A��IK�N@�1%,�.����C��x!��˨[D��EI2޺ЊD��<�����D\��'zq�#|�'��9Qe��c�J�����y �i�'j���ŝrb�����Ml8s#�"�N�i�F�0>I�!I�}�4�E�8x��D�T��И"l�	됩�Ek��p�i˝hٮP��`H�M8]:�(D�����&�R�Ӂ��	�LXj�*��
�\x*e�˃.#~�Ă	>R���j��c���X�o_P�<A�b�74�� !0�U�/
����J�<iF ��V=� R��$!}�t#Ch[�<��NѨN�كa���5��h�L�<!�,�0?�`(��D!cT\y!��GR�<)#� <�j��D��Y�a��L�<�tE�>,�5�A��!�di�'ɌK�<� \=K�?l��ّ�X�����"O�aХ�N�Sp�%�I"p���Ƀ"O8aևI�[~��#��>���q�"O�]�g
^�����w��A�Q"O��{dj�:��P��>�j�C�"O�pf�-|!�,�3�_�����"O=�p�^8M�R��f	�	�|�R"O(ě���m^���V��4 �����"O�M�2�	q��Y�b'�"ai��� "Ozܚ���8�0��֏�!gNr"OdT�Ջ6ɞ�Z��!6(:|zW"O|8����"��;p4�U"O`5!��S%`�@Han�Ct��0"Ob�Z�GX���1G(z����{�!��%A�����#cK���n��%q!�Y$��X9Ff��:8�����\W!��ƞ:��1��ȝS(n��P'� ':!�ğ�#>2����ǜ#
���f��O)!�D�-0�fH�Dʅ�;Vnd��,!�_(���q���>eCr@	ep!�d�M��ˡkI��D����� ��<����'pB$��!O�P�2�b���8CF�
�FL��I�=ƪ��aًD'����Ҝn�z����&0��' ̪����z�)����w�ъ���^���J��I���p0!�I5x��q��2Vt�O��2�4�)�.�ꎾ R @T�])��'�=@!�)�'v��CQBʀ8��TQ�Q�7\T�!�C�T��'�D�G�,O\��go�7���BEQ�Ig�D�C�O��A�O�צ����M&�p<���ԤJ���a�M+�ʄq�(�y+^l�p��=Q��#?��&�B���qbB%<~,}�ʂ<�l�UN�.,$t�c�3�D�l�$u�g��`,,��C��m�ԟtȠ���?�@9�Y�!��y�D剥Ld��3��;�`y4�� fe ء Kc �-����#ȎbR�]��e3
�|O\��S��cH��S	il�)b	S,X y�̉6[D<����G��M��	$g��)��@�`�ɽ{骰ZS*-Č8��I^����u%�� EĘ�[�`֝5fw�EyR�]yh���A�&�2�5�B"����ƈ��pq(�(��\>�`J<�T�A96}�Ŭ
�\z�)�#Ư^Kv�:�����	����|�pݨ1l�s�#<��.!F)bAS@��d�!&�\�Ed�Ȱ)�c^�+��f��O$��Sd�+pL��i����V�6d@�D�I?��O�>��-υN�����W�:��,)p+G�T�X�u��?jq>T���iP�>E;bA��U�+6!J�eF�Q�'��0�%H�M�Bs��q��ϻS�MЗ@њE۬ԱF���Q{�!�y�4�Ko���10�w���S�v���ω1A��lq�G
U+ 4���'z��d�6Wop�R1��"٫&d�?c�@��'�3>�t8qNў,.�#`)�|tr���A��͉b�_9�RO���t�7Jz9l̘��jM�L@�O
����֬)�:���L�$Ty�#<�*�6.+�����][����-�|P>���!
Ypu�� 
��O����QTܨ��ڇ�:�"@Y�擛>��P(�	̒E�7Óc��p$��Df��RTjA�4��D���I1��DnV�s�-��_2y�L���Ѡ.dft;s�"A���)�S�yW%<����A�T���e����5�*B�}���	���a�X��;��99���d>yf�т��Оs���_w��D{���1�Ä@[;Q�e�M��t����'�z��/ڲjB������	F�9	���.y�x@*��#�z�\�)�p���r1�Ys�X�����*}=S)�f瘸r5-���1�R��1A�b�	��%����ZF�R�3�\��J?����6 ��`�bS5q����u�#�ts�MCҀ�2"&uS'h:���45��KSi%k⎐�R�5N�PM W��TUP� �oe�PD��O�Ă`&N�"(�a�2N��VІ}���OZ4�ʔuJ<�¶��%�0|!L����1V�k$&q !Ц�Y�#ɅX���f��� ���I,R��x���SQ�!r��^1��b�(�������K�¨�ם~r��3Wx�R��C2E�I �h�\z��Gn\!� 4��ǋd��p�cEBæ(y�M�3
��5pw�ÜZ��Db��C����^����*Ҹp���� 7d�d���2qhNt���S	c��E4������Rg��*���(�NŊ&�^+2	UV]� �D���R+ԭkt��Q?�V�>����m�fś�������#��w�<Q��/+��X�㜘�>�xd�ͦ���m�{���5��U��y���T��&M��3U� ��=1��	!8&j��D�g($@;@��KT�R2C���Ԙ�F24�� ��Z������W��8Hz�Ѓ��_�X��@c� �Q>=I��Ҹ$����*"��J�+0D��� , �U��ev1��a ��>���'�Ȑ�q�D�i@Ο��|���.o���x �'P
8l����@��,���,{�0�P���B��"ѡD1*3t��w
RQ7��=E���s����W�9���1f��E���G}�`���nً�dD�zdQ¡Gcr�kea���~��9b�8��4V�x8��IMƖ1PK�u@��	�j@:Hr6�)�)r�K	�qH�牪s�q����.Che� �ə\�.B�I	U��@sgπ`� ��F�/>��'� a�aA�Wl�k!j�X�S��mC�\s����ګZs"l�$�3�p?�aLK�	�b�X�R0i�:C�Մ-G��Zc���a8<%��0�)���ґL�>?S��:tj�,S��5!���ͳ�%�n��VV͑�I2'J�zA̀5K��'����əSN8�kF�Id}8D���I5X;�mbC�"�)ڧ~:�8�߷,n��˘%u̸Y�ȓ
�\zu�G��P�C�"W'�ႇ	@>���	�E�Z���G�hND�+a��
�'^�������"�R���+�,q�� ;�'fv�b�$]�h����e�y���dF"X) 
R���'�lQ!ІCZ,r�*�1!���}KS� � �4 (`Cb$9�'��%�0ɧ=ɧh�<��%�*����W�U�l��"OƩ�l3�И:���Vu��>q�]9 3���
�Ƕ)�G�Zj�F��0���y�@���2T�L<�&ܑ=b���L��^�Jĩ��L��=��)k0Hɵ�߈xЮ�	��L�M-�mG}2��X��ȇ�	T�Sឱ���ɫi,��mH5V�!�$��2��W�XF��cs	)Y�^���r�x�rrG���S�O���� P)p�z�C�k	K�f��'�&�@s�O;F�F)���.G����L<���r)),O��Sv��(*(��	 �$4���U"O@�ʃ��S2���(�ho�t�f"Oș���ۋ"dVPr��� ~�P�"O�Q)4�[�p�A���Z�$5�"O,0�)"<q|�*r�� 9�D"OV�� _��P��BEy"O<�iea�F�8x���-?��k�"O 90�
�(O\x@��D�Hks"O�虷�K�?�|�/E�b�0D��"Oz�:�a�$���{���T��t�Q"OjxP�Ł�a@�c�1y_��0�"O���C�Ι0���p�ၑ==	�"Ox\��AT�tQ́@7�7i6���"O�)�RKD�SK=Q�	
��p�"Oި��k�2"G�p�vZ:u�f]�"O�m�F�ܙn�@[���,��Qd"O�0,]��Em�)���Ӣ.D�D�r(C�D}��ɘ8QG�e"B��o1n�{�)��]������00*B�I�/�Rq�X!_��mawɞ0k�C�	8����W�������G	S\~C�ɻ9���Q�aG�Q�%�6G�$�<B�ɒb<�� à5�Vye�8B�	�Js�M'�ef��`-�' HB��wD�p%��6 c\���C�	�4ìLja�M5z���/ �L�C�3i �� *݄8��q�Q��0��C�	��q!Dȟ�
v��H��r�rB�	M�h�Ǎr⒬���)T�B�	�^�:�J���Qt4�#�R�|B�I�^7��teY�]�b\�Nsj�C��kP�@@,R yh8C��:]_zC�=)L���I�0AyX4��*ޫ�NC�)� ���@�ܑ��â#6�2�`�"Oj8�d��R페@6��dXB�"O�M�`E0�l@�J�d� "O���4
�:ʌ��AN�'�Q�"O�����7k6��ʇ��x��q"O��3� �GS�U)�oCYy�TrU"O��b�-2]�	�0�7re�s"Op�j"$��<�F�R��13T|��"O�<�Q���4V�P���P���"O0H��Ih@�rb�>oN����"OL��.�= ��t
�730�}�"Oj�[���{wx���0D
L�2"OzqC��/:�(਱�7` ��"O�XG��-�<5 FB�%gc��ks"O�4%"�?
�$��!�ULX��"O�Œp"��xPRC��1o9����"O���u	ҙE��a��
�9.\�f"O��(�[�NKV1�Ώ�62�[�"O�Lb�a� _;R�{W/�g�HĪ�"O>l��Y"el@�$�&aʮ(�S"O"d9N��0�*���㟴���Q"O4$s�;N��ɻgCރQr��A"O�1� |$Lu�g��;3``S"O��!r�3HVl�J$]���i�"O�񀐍X�kz��n�!�,��"O��N�3�Ġc�]�ov�s�"O>�!��B#㦉����-/B�e#S"O(Bnۛr/�c�a�1.��"O�S��רk��	�2.���0"O��2Vc�!f,�ŪH�&|�)[�"O�q��۠%
ƀR�A��L2���"O��cj>-��3� ףN��k�"On����0�-��i�4)�"O����� M�L�M�2H����"O^ ��΀�����	
!&^J!�"OH,1Ѯ���F@`�EP�)�Z#"Oܤ�U�\�O(��Ņ�&hj�kD"O�Y�M���t{���!:hx��"O�� �␎K\ �f�Z*&�N�S"O��J�,�?�4q��A����8"Ohqc�S�^���`W?d�$"O�x�����O� ١���]���"O�HeB])�6題|M2�)E"O��
U���<3�`:
�+/(4�D"O�|�weǼ9r)����A|r���"O�U�fo��
���c+�o����"O2���mUy&��R� :q���3�"O�pp�#r���E�9,戣�"O��	4͏�1/$�Q�HסW��A7"OH�x2G�RF�zH��kn٪�"OJ\�7*��&�6<���!#�t��""O�$3�OF�{Q8������t�H�is"Od���k�
vX��6/D�v��Tk""O�x�P�?kҶ��d$�7�tYt"O P歃�t�X"�?+�R��"O��[RM��"Y��$�ɉ*�p"O���x�۔)�w`�]5"O$�KqOP&<
�B��	DXq;�"OJ��U�rpNp�I��<�m8�"O� ���A��� �1ba���[�y�䂁)�.�8�&��Y(�� ���$�y���CT�rD'��
}�qG3�yR�
I�s�
�|���¥H�y��	:"/�,�$C���@ƢG�y
� ��C��ĸ,���0(E1
`41 "Ox�C��:%j<m2���;$�
W"O�XC	���9p
DZ�h�t"O���Nz��]2B)�q
��s"O�3�j�SԾt��g�D��9;G"O���!0ڨ�{�EƂGڒu��"O�%���Q*[���n*݂�#5"Of�p�?�4�A���>�P��f"O�a�` �BJ<Ժ��2�K�*�yrc�]��@�!�CLO5�N5�yn�NKF���)W2i�jW��?�yB)�3���a5��3"���Q��L��y2��6Ks��agH��T� �)�y��%S4 ��BhpՈ
�yB&K��`�V�G~�Eߨ�y���Ju���/ܧS^��Y�.�y"�����������g	֊�ybۖ(cda����:s������y��, vy٣gŴ�BD��cS��y2@�D���m�Z�+w$���yr&�(<�HؕF]?R� )7-��y�o����i���B�6@�*&I��(O6����_�^��F�S
��s�jG3G!��REIv S,�>5͐�P6ʕ�9!�č?E�|�WjW��vD�b/�� *铨�>!f�_*��-�čD/K�8��U��C���!�����A�l ؜��)K'-��eK��:D�4�qṀ;A���`�
�s�<]���3�Vb�D���l�(q	 E�${�,����y��˫B8��5��<"��r!��y���>8��W�7ޚɃC��=�y��4��`P��߅'p%Ȃ�� �y�, 
SÌ! �I2�� ��yb%�����*���(2k٫�y��Tl1�A��}� ���G_7�y��΋*-��Y�HEGX��Ј�yl��k��X!�!��:�^�!@Ԑ�y≓7X2`��7�`��JI�yr���}�Q����e�:	��<�yH;z�< ђK���|�ae΃�y�j�����"HL�����1B�=E���X�RD�����L��X���z*ȇ�[�8[W�E��V��g��\ 0�ȓ[!6JB[�iq�ԣP-ˣk�:̈́ȓ/���gZ�V�p��a�H}6B�	=}�͙���p[��a�bB]B���>�H>9P#�' 乹!�3*^h�r��f�<ф�ٹ3��=��M���|��O�L�<��/Ϡ:�rp�peY�
�� �H�<Y��B�pM�uPHL�Z��M�`��\�<��2�e�!j1:0��&�>Ii!�Ğ<	�.�P$O�6,0��C��0Z!�$��8Q��A�'��M��vH!�RQ� �P�ƛ`�����FWU!�Da��oӷaq��&.��*J�Q"E"O&�Z�	X�_X80��N�*6�,�"O�͉������M �h�T����"O�U�T�S8v"�H��C�S��33"OD�����;|n(�!�'V�(�u�$"O�T¤�ŜH�H��a����!�"OdC���kǠ٪S��
��s"O�b%G��|t���i�l�B"O(�`(`-�QѕaP�:#�1""Or��p��*��u��Y�u&���"O� �YE*�2�X�*F�Hl�*��"O(�
��ªS4`B劇��1J "O�Q�'���ޘ���ʫ[���2�"O*���	&7��E2�q�� D�4��)ͧ0Aj�zgG���͋�1D���U㐶�
}��R"O�es�@.D�8���E�G>b-�%ύ=ahA+B0D���e�Դ`�h��P�0{I�{�	0D�h���[ ��ZƆr�fQ��#D�d����FB<�1���w�2e��C'�􈟸%�2�<�� ��,wi�Q8'"O�!K�\O�u�AB�T���"O88���=a i�b]�zQ��G"O����_���0@ŒjJrTk�"O���0K�����$��+���'"O(}k�L%3���h��ք2�"O
����̔Ȁ�Ѷf"K���8G"O6��g��U]� �F��HjV1i"O��g@w�(���GT����x�"O�Tb�hV;.�����+f�Z�q�"O*��7K� ���N��C$"OB��P�@:k,Ը��Ԝoh����"O�\6&#T��TP�x�ܠAe"O�%caE8XY��4n6e�2��D"O����aFA@|�7#:� � �"O:`�C�
@�R�ʢ�
5Ӡ�:��'$qOZ���n]�]�U���64�0��"O�P��L>M6�8b�P����C""O�49w)���Y�p"����!"O
i�dH��z Z�Z� �6� ���"OШ���:�@����B�C����"Ob́��QgZ]Ҵ��� ��"O�xCMڧ`�@x(��B:W}(ɊS"Orp�<v1ΌK��P�ko�U��"O�0�h��G�̳��(ø��"Oj��$��e��)��̺e��A�w"O���SL��#�m�d�\=���8�"O~Q�%���d�%�Sd�0��W"O9���=+D1�r�Y=7o���b"O��ࣄ�5	�0��	~��aU"Oֽ3 ���z��#<����"O�đ��ξL���j ǖ�S��8�"O�سU�lܠmHw 
���b�"O�0��i�I�n�7ŀ}���I�"OԴ�5�5�`0�aD�S"��2"O�,; :IP���+Qr�*O�����7'h!#�W�l:���'����ȷ_��Ih�MI&b�b�Q�'�Rl�t��,N�PA���D�nՋ�'��h�I��8���0�N�?����'���%��@�d�W��H�Ȭa
�'�X�:��߄����C�4>��x	�'l>�P#�V�6�q�S):�Д��'���s���M��a�@�~]~H��'�����e\Z 2��'*A�h��';,h�#��;�6�zЊމJU�� �'���ۦ���lȉ'�F2H_�4��'`m����{�M���Z8:��Q�'��lZբ�U+HcD�(:����'���D���M��!˳㉯�����'�ڽ��b��&LZ�k	�b��'�>�i4E\�Zid�P�Ǖ����
�'M���ł 2%��� _.,��'[���r	�3ߴtA얬\�t���� �5�HW37G�y� ��<AF"On�	$K*.n�S`n���<���"O��+��ƺ����#@���"O�tS4@҄R����֢Ąe����"O�xĎL�wb���2GշM���`"O���a-�#"��-HC��J�b�R�"O�%;�&֜!��Tsw	ʃO��3"OL�b�^�5�ٲ�(Q��T�(1"OR ��Wh�) M׏@�
d*A"OxM	�HK��Yu���F�(�"OJ��
(i�̬�G�U&`7
b�"ON�9���
@4*�%����"O���%���"�(X�Y�k"OF�aA�V�n�jx�G�+,����"Oޠ�W��3$�� ��;@�
1 "OJ�VÂ=Ft��Rb��cj�:D"Ox��7�^�"�q#M1�t�f"O��CdX�O
j�A�{ (3u"OP@�S��*�|���oJ�VQ�!S"Of<���F��f�a�]�/;�( "Oz����V�[Wz�ϝ�:����"O�P"�ͷ~��	K�`�!Yb��"OnDR"o��$�m
���8���"O^I��Ь}⁮;�X""O�Y��J&n��ٵ�ɭaj��"O��)dj�1/(F�8q؂�,"�"Oi�t�O$�<u�կ]�T��Q�f"O0 (����U�(�� E	R����g"O���֪a��!j�i��	{T%��"O�F��)���A��Ra^���"O�8����-o���B"
D�^U"OT�TM�,&�(�LU�љw"OP�pu+�4R�T�S�A'C- R"O��� ��7c|qk&�R�b/��"O@XY�,�!g��1\�9��I'�yROL�F51�ÞZ��i�#�ݛ�yR��+eT@9"�`��4 �m��y�AW�M�f�`��:<Pá޷�y�#��<kX�)�D�.)�>���]7�y��X�+i���@�'&�`B��J��y��ɨI@�-����dv�� W�yrE_ ,!�Aa�HO���x[�e��y���Qd`4P����ea��y�9�� �g�6���b���yҢԸ_���,ٴ4*��LK��yB��_��x���TqB��O���yR���X�A�dҵA� g���yR��%)|r�1���n "i�����y�a �v*�PdD3Z,������y�lٕ;���j���"�
=�wB�3�y2ÙN���+E�0�\&��	�yb���K��H��FT	*!^-Pf���y�*ӻ2��p�/ε@�Ɂr'_�y2#�^��@{��@�pQp���y¬�6�(g��x-`Ur����y"�I2����DtA�Da� X��y"�K�
��͸g��j8a����y���mJD���'d��E�cd�<�y��
�~��q#T�U� ��ӯ[��y�B��_�ހ!S�$;�0��#`\��ymBQe,$���U 4��a �����y���X(�\�����(�,mB'o���yR�,a��]s���v�['��:�yBj�(V/�%0У�K�t�y
� *	)F��(d��p�A��J�@D{r"O4��j�8YC������c!��"O"��� �%�Ȫ��Z��q"O|5���h� ��#c&�a�"O��0��� `?J� "�ѷx�s%"O����_�@h��0W��N��\
V"O�<���Dtj�`Ɓ��Ai�"O�܁q'�.:p�a����~�ցk%"O����ܲ)01L�'y�p�Q"O�p�RKV`��9CP�Çn^|�R�"OF0�7#zmZ�,M���a�"O�Պ3��"�6�q��O�I�1z�"Or0xe�W9.�����xÈ��"OI���?I��4Ӵ	E3O����1"O�=҅
�2�"v�V�OuR`s$"O:1�n�T6ʘ���c,܈�"Ot��a�O�>�Vaj��WbO^�� "Oʌ� a���,��%W�����y��G'O���G�)o�}�!�D�y献Ae9IW�Ϸx��@rE��y�,ֿ+pT�p���p>��1�S7�y'�#/��rDjR�?j�������yR�ޒa�؅�H�!�L�����yRBM�Yh��{囂�z�B*�5�yR��(7����Q�g�~ J ��y"-�C|ؑK6m�P�ے&ت�yB���Kh��iH|�t�P���y��U�Ҙ�e�oG|4R����y2�D�K�T�r`��c̘�&)N��yBG��?�"M!'�כ[1X��e(��yR�_�f������M|6I#����y"솽H�	Q��J�7L6�Sa�\;�y"·8	uhذ0��\L��˻�y��فsL�1��G�O�ԁH��ũ�yr����;�ܝE|������yrϟ�wI���"�!(?P9��
=�y�+G	W^qѢ�P>�x��L^��y���9�,�[���+Y��l�R�'�yR�*E��y �h���h��]��y���>t��	��%�D�kO�y�Bۃ%2�a�-�6x�f�a���y�fA�YSȕ���r>�|Б�ݽ�yRO�FL����P�=>�A����y2�](Y���jA-�>@�i�G��ybJ�&���Q�֫=�F�'��y��D9%���x'���.�dAF�)�y�+�9e&��(�.��e����yr�6����hT9O�`W�е�y�
�>=�60����)%0Ijv	Q$�y"� Gת	Z�c�(v�I��g���y�F�)���@j"J,�{*Q��yҨ՗S)�=���6h�.�y�@��A���Aa1�����y��+f����.��4T��g_��Py���"E��SG��
��Ɏq�<�6f�%(��"Ň�0V��U��V�<9�[
#?�a�� �-$8֑ pHy�<�1Ϛ�1�-Vv'p��E�8D�L�U,��r6|iqa�ҁX�Z<��j*D�B%�C'-����"�	u�	�4'$D�X!���<	 p*���2Y��D��>D���G-��Q��U<ڸ� �:D�X�#�E�|��su�s�LP��9D�kwA!#�9"�ʰ7S�@��9D�� �xs��N�48b��p]`<:t��"O:��e��0��P�S�FJ�"O��Y���3]���E�3Z��j"Of y���&�t�A�?NC�@s��'��$K*&>a��`s���&�)r�!���(5!IX�����Ы@��O:�=���T��,I>	�1p��	��,j4"OD���@5$��<��ƀa�v4��"O���b̛����xbeܻ(3��c`"O�@q�Y�;�J�`Dװ�d �"O��)U%@9�ԊAC�9I��	�"OR �f� 5����:C�AA�"O��RӏG�z0(`�I<:0�	�@Q�h����i����/O�&�
\9�mC"9�C�ɧ\
�Mic	M� 0q�v̀Q�C�ɬxZ<�c�f���z����B�	!D�MYP`_>#&-����'I%��O���!LO��Y��}�<L���x�� 9�"O�tq�M3�.�:F͖�"����"O�� ����L�4H
0g7J��|2�'�I���:X	���5�^D^�Y�'o,x���:!��UJEj�����'���ۀ@9(5�
�BF���y�O�M���p��%��F����'�az�U����`ݟr4�-Y���yR���-R��7i�<B�`˟�y/�<Y��J�%
+a���aN-�y�L$}]�X $u��Rh��yB�	?C���G5O	�<��&�Py2�^(�����$zH �6�_t�<y�_�XUn	ib�����p�.�r�� �ɹdt���`�JpA�i��"J� ��jF��{DOY�G�����k�,ȆȓD��@�@�!�<��G�T�5`��ȓW�aÄ\�h�l��gkM�l��=��^Yʕ0��5�$A
1��^?��ȓP�@�f���wHdb5�%>���Dm�HW�˛UeL�"Å %5�� ��W4.�c��W�<�.$	�&��U�$i�ȓA�u��������AK�+ ��'��D{��Tcd��	��\1�.�t����y�J��`��6Pp�հ�y��R�e1HHc���-�,lY`-�y��K�#}�!d��<<�a4m��y"��+ ���!p����=ғb�	�y��B�g �Bq��'c$���X$�y�U	H�,i��Fºc!T�jC��<A�����P���Lد$!�8���3LoV�OL�=�}2�-ʬ~D�R�� Kl�$�I��<��E�\_`%�'l,���D�<�W�ZJ�����#CyT�zd|�<Y��O'c� R�lãf�\\��Ba�<	�͚Y�Pӣ"*e�tC���G��4�<�D"��Xʬ�S�R�$����	A��T���OP�Tz���"K�-��!�%��q����5�b�� DD1��i7MR�E]:\�R"O�����_�!N(@f�PQ�t�R�"OH�QB�6zϔE�#i[�d�"O�а!�yM�p��փo��8��"O�+�6'Hā��"O{��C"O��a��5Zr�M����ٸ)��"O.�(TeW?���'�4��1��Io>���2$�f�V%K=kZ�ukSG7D����G�$.��sɈ!sU�e��:D�� �]��	�e��b�@ǻs���:�"OF�ʧ�ٿf�x��V�	
f�"ݠ%"O�Qi�H�@���)!���2�L��џ|��'[�h E�=G~��*� �BT��'�&PcD*�wB�I����w0��ڎ��7�X��j�_�6�I�!R�5~@P�A"O��	�`�4%?t1"�n	r�L1�p"O�U��D]�e���&C # �����"O�%;�`O??&ı�g��`M�I�B"O^���ʇ��KS�\%��id"O���Ai�z�8s�d��\�"O��@�
)U��
*@���t��U�O!ʵZ�`QR�n���!�� �.O���7f�^*�C����T�1 �f�!��B]+��Krt�ݪE�!�d �t���@ /��!���I� �!�d6��8�]�3�@#�K�XG!�D�M/�u9d�V�O��!��Y#�!��-v�$u$'I��E�5	O%n��'�ўb?�X�b�M�>L��"ִxV��g\����I3I� ;�9o,#V�pfC�+&WȠ0��PL R�r&�8
�C�ɉ^!h�P�M ADؠ�BP�C��B�ɬ%n�9���>2X�q�N	"RB�I�1�Z̢��H�mlTC�
�&\ B�	�_$P u��>`H rDG��bB�ɂV��q�2�F"6���"�)��C�ɰ �j@�	�	7��YHr�9$�`B�	!S��6����&A�p�@�m�2�=��'@����l�zL9�E�B;`���FR�����@-F�tٱ4�V<�܆�wv��WJ�4�����̺Z��0�ȓW��TJ�		�JSd��R�R���ȓgE�x�dX a��-��P8$��=�ȓ~���aea�������1^��ȓQ'$�kҨ0(rd�ThZ����ȓ����1������Ŧ��ȇ�B+�1ah s�b�H�`ӭPJb��?��,��q��B!N�@x�ç/Q���ȓX���I�2���X�&Zeȇ�;9��R�C�@�Tp��g�b��|�"�)D�J�)^,q)����`B䉗nY�8i�+ɋ7�
a�C�{�|C��/kG*�� h�B���:nZ@C�	=*���4iy ��	PHӍk �O���D<�z�9�+\�-A��q�(�ў���	�z��ar�ǄS~���smJ�\�8C�	h\ Ku(W�L�H�����.�C䉘N����[�[y,�HrK��r�C䉲W�ٕ���u1@d1�(� x�B�I�`�CV�V�6X� �7D�D�zB�ɇ��-+��?bM� �Xq@`5j���'��`o�<�4�rŤ���ۈB�)�df�Me@��c�'"������'��'+��'9
�0:`�D=���!>!��V�g`0#���-�,��F�9-]!�$�*@�nUa�fX#͌�x�&�%!�D�7������1`���d <!�d4e�4�R+ʕP�1�6���)!�d�
ir�����˙&BdMS���)K�'bў�>��N�z�`4�2"�x):��A�Ic�O�"H��K�	70����CF���'rN��a*FS���؆dX�'��U�g�A&Z�x��7c�<������ �X�so�sd�)%@$i8�X��'����0����#ԉv��x�u�X�]�!򤋞y��A6J�)�P!`�C�1em!��Y���#c�_�TH��o�<�5O�����=,�Z��v�xq�"O���@V�J/��1+�>�TB!"O,�!�
π|�.� Ӓd�X���"O��ʤ뜬UT���cE�N�`I���'�1O��qBӯ(�՚XY&����ៀ�'�ɧ��N�"�
��H���w
��/��-<D��١� ?�����f�	�G�44����C^�"o� �'�R� 3��b�<�#]�����_Y��RP��Z�<9��1J.�q��"��C!z�#a�*D�|����7 9���b��40���1eg)��䓹?�ʟ������P���@&�f1���S�XG{��i�U�Ddc�T�j�D�b����*D!�D�4��JcG�..i� ��34!��D�� aAʖ�(V�K�CB�9�!�DQ� F�$�c
�5
6��S�@6O�!��V�]�����Ʋ7�I1��#!��P`a��+N
tVոC@U��O(�=ͧ�y2����%�T��v�`C�>�y�F7X�Y"E�K�$��!�n��yR�@�~.���WGK3;�X�+�l��y�jte�)PBfV(=b�8���y򩆻X�|5c���D��A�����y�/��.Y,YX��֍;��Qe��y�*V�w 4(y��I:,�`�����䓫hOq��i�ݰX��e��4M���J�"O*i��;��u8oH���T�"Od巤Q�@� vhbY1���y�*Y�� J�P�A�ZX��gX�yB����.P��$��9�d����y"�_T��qjB�9D�0�cT��1�y��Y�`
Z0�/�Xi�Ç���?a���S�q|��� q�ȴ�Ӫ �ގ&�Ԇ�+�ruӢ�_�"���D5
�C䉺)#ެ)���k��Y���fǔB�IV5P��A�Q���l�O��.�lB䉎u�2YH�H��QO��ye �r@B䉣xك�i�"������(qu(B䉃0�z�� �,n�	��\�p^�C�	*�#"'M#���\Y���$�O�����/^Ǽ����Ӹ	7� �L��'�a|R��	ejH !Ő�n�L	�Wl�=�y��S(��ժ�!�h�i����y
�lƎ<�bC��K�bQ�v��,�y�!A�CJ��%�X
lc�eI
�y���c�X���/B�܁�ؙ�yR�	(g�[g�.@��:�/\��y�-R.K�,h����<KF���y�*�Og�����-J�q�&l�y�D�(;��ȃ��Tp�!��H��y�˞%�bH(�`��`B�І��yRn�2Ud�s'�'�Xd���G�y�f��F=5�
߯/D��6Jլ�y§ 3	$v�!�G�)�,щᇇ�y�*�w:]0gG	� ��Õk���䓓0>1sJLL�v�[ �H�5Z�|JG�WC�<y��B�6PJcn�[���1�o�t�<��d�a@j]�C
H:usNHie��n�<���K{[ެАM��=x�t����g�<�@.�$�|kB�[P/�`ąN�<� n�Y��)#W��B0�Έ52��j�"O����FO��8b��D��h!U����	��:�BGm�@̘9��C��B�.-D��mL��0�b�'Z�bB䉪(pHt�C+��,��b�/q�B�I�JlhUXg#H4x�h��L�=!ĢB�	���%�C%]��e3�/	��B�IV�,H��aܖ8c$lK�ύ<BB�	zd0Д�Վwd��'�=��O ��č	^L9ka��=T�ft���	U�!���n�2,�@�ߵ;��H���u'!��ܡe���u(I� ��Qo!�3:4m"fm�̨�n�)�!�	-4��=a��s��ô$n!�� 	�<rB�@�:�\q�3+�!�D���ӀfT�j5�P�PI��[�!�dӪ ۴�"7�E�! �=�u��	�!��C�lq��A�
e*��� +�!��Ty-�A�M_f�b�c+�5"�!�䆞>h$��ʛ=��b���S�!�/ڎ�r)�&4{h�[���3��O���$
�Np0�a�@�"�E�D�!���J�P�K�zjT�JS<
!�$�Y�U� Ύ�+WĻɍ1H!�0��}`U�Y'tFRp'��-�!�$o�1�'�ەB�r��匮f
I��R�jT����3'�<t��S�eǮ4��0ղ��Ei�.P�d�0l�� t2I�ȓ�b-����	"��f*F�O.XՇȓ
n�}��C�n�D�QL�ȓ>��4�K�b'��3D$!5���V�.�� ^:O�x�Uc�:����8[n����0{DN���0mb�Ԇ�:��h� W�.�,+rH�ȓ�Rl�L�H^���E��������IC4!
�,q�Θ�	��ȓl�z`��%�S�m�Fn�#�nهȓ)����jtN|=�aUV�4u�ȓS��q��!��JP��@)ev��ȓ��h��K�����j˧=��цȓbr�e�f�C�g0 �F�P#]k�U��m)X���;QpR�xª�E�q�ȓD�M�V,�C���4m�'�bx�ȓ(�.��͐�Sd�u�I�F�*-�ȓR{�t�sa�V�����"�h��iԒ`[����h�!Jǁ�G�����G=B���,�y_������Qz����>i��LFS|���+��_��m��,��A���C�/�QG)��@����t�������`iH>'!�9��ʞ��툤�/D�H�6��*�<EH0�����UA'�-D�P1�HJ(Y$Q���D����CQD,D��B�� �`�X$��KD�w�iJ��*D�,J�#H.���J��Td�Q�s)D��"Ro��A�6kxȪ1R`&�O�����UѲ@�C�me�yhp/Z�Z�d4ړ��OD-jb��L�H��+�,%�*��"O `���&�N���B!Y�m	�"OД`�(�<z�zh�ǡ�zS�"O�1�$Ŋ&�1� V�8t"OʝJ��CJ��Ю&<�B�Z�"O�۰aw�ꔘ��	���-I"O@�
!n�4ͺ���ܘ�:M�#�'��'
ў�Oļ�)ŀ����M�S
�b��� �#sH�1�H]�w�#�9�B"OT0f��J����ܡe�""O���7	�� �  ��)��q"O��׃@55�QǮ��Y��Y8�"O|-C���";Ă�����R���'���ߡ��9����,J/N5���7]�|��)�d�T���8�	_�1�ޓ�y"㑼^.@pB��L���� #����'9ў�Oufm���\�͋��UU��
�'TJU0��ޒ{����.��U#X��
�'{:�� BC�!��KS
?v2�
�'ܤ����g��� 4X�/{�� 
�'k4\���1�x�dAǶ[���Í�'0ax���d2��x��I�Z�#H��yB,�P�P�ޜEX���a*Ѫ���hOq����w��i!p�YÖm[�"O��2Ĕ*���0q!���8
�"O|}���*{G��Q�{�xY�2"O@�	�@�<\`*0H��k���H�"O�	Ѓ*
���RAG�[��md�'�ў"~�1EƼ}��є$�#9�z�yG�	���=يy��.<C�D�k
�C���2tό2�y�X�*�ȥMT�)�6��>�y��Ģe�>Չ�& !��,x�����y��9L�J�� �Y1����y�(�����F�X=JB�A5�y��*[�!��y$�����?����S�v{ٻ�f�)Wa$�A@[�j@2�ȓH�������<��	��M�.�=��W�l��Bb�7�V��I�*x촄� �2\��枎8_b�����L����ȓ#��49���?�`��\Y�^ԇ�.1�0� �T+�2%�0`�T���	��)�a��͜P�A�X��8�?��.\�y��K�0�q�ë�o"  �ȓrR��c�� 9�HP%�`e���rz��1#DVzt�!ůs��Y�ȓ���jS`�i �`$)���F��+�\�#bK�(R@h��F)�X�ȓt�H��9&Ʃc4G��cptȆ�|y�Ԛ�L�8'h�SӅK%%`
y$���'��>��4:�N)Z�����c�O<��B�ɌY&ب���� �.��-F�B���x�r�`�+���:�lZ2hfB�	�,	�l;� _!=��`3e��U�C��:Ԯ���M�Pv�D�fA��ftC��<2�b=S�7����a �~\C��^a�����܂��[B�a{ C�I�od���"�!xt����H�HB䉵<��mIsg%+X�v�m(� D{J?���	��S�:\�U.MX,���H D��QFL�6Up�i7�xX�=�5�1D��ca�U6E!��aپ��A1D�@���y(���0%( ��q5�0D�P�Si�>Q2�j֋UlxQ��d�<�H>�
�'L��h��P�[Ȁ��Օkv�A��x�N�Q�o�Ojv!ڠ*�_N�?���~:d։%l�`��+T�"�ӥ��d�<�s$L�L�h�'�&aT� i�^�<)��M�#����gG�Ei`X�D�N�<)�nG'f�(� Cl��[%\r�'�@�<YR%���C��:���A5F�ПhE{��IY1K!��X��"em4����H��8B�I�N���AE��u�8��%�G}6^�HE{J?� ñk�<S6h`�GFd�1�"O�С�lL?U���b!�&W3�@�D"O6!�w�є^�4�Bd�W l�I�"O��5�K�%�T�$�ڷD��b�"O�����R�a���_2G�^5��$�OF����-�=*5��*J�`ҡi�=r�b0O�EY��х9��ě2ٜ9�`��"O��jj�	2f�;bwD�B�"O�,q��
?�8mP K/Xh��1"O`�Zf�D��ur��4FI0��C"OzH��'m�P���P�YLxh�"O�$볈J�~�v\7h�.,�͑f�|�Im~�e
�`��T�c �8�xU�p����xB��V�zh�B�SV��훳 N�7I!�d(J����!Z�c�t%.d����"O8��@S�p0�Q��H�Q���"O�x3qH�55=\�S�m�4�|]��"Ou�$ͯ��eyb�d�l�1"O&�4�		1�~}�NN��\6�'w�'!�)�L~'��0��ɥ�@�
&�	� F��y"�ߧIIZ���0f� aˆ�y�����Q�S)(萣�;�y�+ЍG�*-q�l�R�XM���M��yb��:T
5�$�C�0������y�)֔P���e'G�,�Ѷ�W�y�V;�h��7D+`�|����D,�O�Y��fQ5<ײ,s&%ОO�V$�0"O�0�_�g��\��M<h��`�"O.��D�,�l��"J@���$��|2��5h6az�CPԆ��Aa�]�9����y�E��`q`�Yi�)�D��Q$��y���9I^��r��3�Hz� X<�y�*�>-���E��9�>���Ɲ��y�E~}�Cě�3�.C F��yN��.^b��}D^Pq����y"�\&(mQ��1w<uI/��?����D�<a����5e�Ԩ��-�PSE��!�T({��b�̻~��ј�,��!򄛑F�9t-�##MT����!��K��er�(��a�б�rO[�e�!��-)XP�0��E)�ʍ�r.�<C!��
	Z=�� ޠA5��hӔ^���M��4���̰>A�����"�,�P/#D���G �Y�c������ #D�8��`�&>-����e̮>�p��$D�,a��(���y��ԣ$�D��&%D�@{�F@2Bh}	�n�3�M�QE=D�h��J�?p8������ "�%H'�?4� �2oI:o���h��'H~٪���H�'ya|��ߊ&wf��Ӂ�$q���Co��y�g��R��H� @��i���*��3�y���sfz� ���a����(C �y�%6g����Oٖ[ ԼRbJܦ�ybM���B�jG���V+�I�Q��yR�߮+�,�"L�G��:��Ż�yRkOi��0���̀Ft��i��+�y�̓�%+ڬ
����f�iY7H��yRnKd� �3F��¡�f.���y��h�.]��u3p=�jψ�y"��E�%s�L�n'�!+�
�yr	�8��܃!�	:��p&��y�j��-n�����V�8z�x�	�y�_L*��҈�5�@�Z���1��$%�O��d�-8�Ĭ8&�6"U��9�"O� dDzI|�|h��\	5���b�"O(QI��!&�e�FG�7f�<rb"O��C.�%3z� �GJ{�=�""O��+����_�ZV�]$U̸�p��S>���A�; 8�a�G9�d�G�5�O��uP8��`¯>�j@�SiH.W��D+�������9L��U��"�6�a�8D��r��0����w��U�t�"��4D��6��.��Y�c�B���$ D��:�ڲPM�؊`c	
,ތ�uh8D��aө�#9Y�4l��]��)�Aj�<���#}*�(�(\�w숵0w�^h�<��U��} �ϝ>2F���f�IX���OҐ�`�E�b<��'$'9fm����dЬ'?�u���H��>��'V�^>�IJ��\�'%W)x��&ޠV�@`�J2D� y@,ʄ(�PbdJ�ޤ}�A�+D�X{욇37�t���_H�\PGf>D�����W� ��ز���;cƸW�8D�L"S͆-[: "�J�Z����7B�OT�=E�dC��'�$�U)�kj(�Lg�!��"gҜH���̆&Wb�
H�*�!��:Zn�I��O$%�\���� �!�DV:wJn9ڰ0 ��$b@�~�!�D	�'Z��a�ă%Ŏر���pzўL���+q�6h	���A��+�H,ZO�B�	�\Ppəu��7p��e�:R����$�S�O��`��N�<JƸ�!E�M�7�C��Wl�x��l�@�j4	��{���ȓc��1��Ȁ�!�Zy��*�;>��ȓXġ#���l*%J��j�����^~�s�@��y��m��-N6L���ȓ`���cI8\0��p�Ҷ%L*��ȓ2��`͝ 0u��:F�I�&Z4E{2�'�$z$H�1J"@�jE7)t$�����y�C�gH��OE�|X
R����D3�Ov��
ܡq��K�/V�e86"Ot1���ЎW-0�0W�WI�lB�"O�хJ�/.��6G�&b6`���IE>)��3@T\RA�ֳs�l����3D�0K�%ʍW�8W�S�q{�$	�
�<���Ӣ�^�#����5���h.B��D0?���؏x��\�%�7d�v08�kRAy��'�����2dI�&�١+#:1 	�'����)���͠v�L�o��!��'3VhxC*�m+��;eoʋZ����
�'1r���n��eQe\�=%V��
�'j��Y�T�;�p�PR!��O�%����hO?�p�.��V�rVJ�
�}�a�Hx�<I�̌A���Ǌ ��`ht&i�<���.m&�a��+��/�%ȷ��d�<1�(�
5"2�P���QCRd�2�K�<��ήr~h�"�T�]���#KI�<95��b;��C"��Z���І��]�<��B5c�N�хi.�\�e�@y�)�'M989���K�p�j�R&EXC4�ɇȓhfh�gg����ӈ>����_x�<9��ͷ+�V8�CL`�~ YŎ�u�<Ѱ*o��Qr+'|�<�`��BX�<�%�()d�&.81Zd��H�J�<Y��5]�D1KF2v�()B�L�<�	�*�5�a�	��9d[J�<!���
�	+�.��L�0��HyB�'��c��x�0)�@=�(���� |a*BO݆�\��ր541�"O�8�gL�	�����.����"O�c�� -�V�QɄ�.����R�'T�	n�)�=qBΆ�?ST �񄁟��*�	�l�<�P�\��`�A�8��H3�g�<�Q-O�d�>����ـ 0h����b�	I��`P	�x|M�n��!�tp	$D���4E �b;�=愁�;&�K��"D�8+& %r(X�_�B��SaE6D��
��X�d��v+�gG��P�A�<��2��m�Ba?8jh@ C�KL�|ՇȓS�j��g퓃f'*��؏n��݅�i�`�6",(��˧hY��r)&�0�'��>��*V	�!��B^�^�е0�k �e*2B�I 6�Y�� �̮i�d����yBȌ�d�B�&�dT�@Y����y"��ow��mG�X$��;�G���>a�O� Di�=zԠ,c�ȅ�^:��[ "Opܰ7-�7�����b�h�%ZG�|r�'�az"� �Ӡ$���(4І`_+�䓑?��D1?A�f�D�16bPcy e�wM^�<���Z+�� ��?i���@�`�<�eo6u }B�"�����@�OV�<��/�vb��Yr"Q<b�HŰ" Sx���'�dK�P�8 ӆ��$ڨ]1���hO?�	�.���P�S�W�h4�}�bdU\�'�ax��ޜ\��x�M!-�t(��ǜ�䓉��3�SJP���Oʠ�JW G
1)�b�<!o��4{���M�M�^�q�[g�<�A䜬1�)�ɓGݠ%H2( J�<1�/F�
�p���ʔz�(У�͆D��x�<�S���@	��"]�uk�˟p��[�S�4�'��	A$��$�T�K����CY�1�LB�Ʌq�8�����~���e���L�B䉅%��@y�k G��Z��<\�C�ɪfÆ]QT�&<?��s/ӫahC�Q�v�;�e.V����!�mVC�I�qcl��@���C��1�N�'(cLC��7��`�H�8}�W�̲C�ɏq�xИ��ԁR� Ŋ�x���2�S�O<����ތf���ZW蚶gq�d"OV=�U�V ����Z�nWU��"OD��:��yq�KE�8�H��"OB�(�cB
FJH�3%��o��T�S�'��Ez�٢F��ly�:�jY	a�L<��'H~ɩ��I L�h��dĒ�^�-(�'����	��7=YYtcί |dK+O����S�L�@�����P��OC��P �h*D� -��OUd�YUN)3.�ܹEm#D��%�]�m p���*@�.m��.D�0+vN�)���ˇ�4h��P��84��	�>Xr�ҐG
�Z.�t�Y�<�"��:X16H�ON�_������K�u���O�\"ыD�YI���C��b]	�'��"�N�K�R|�Th���8X��d(ړ�y�NY'_�"]����q�h�8�h0�y"J�+e���:� J~dp���ֲ�yB"۶"��HA� �p� �"����>�)Ozd��G��e�-�ʖ��C�=D���!J]
tT�T`��att�" �ON��!�)�'	�R�`q���t�T
E���Ѐ�'k"Y��o�$���)�l����$%��.���k�X	J&"p[��Z�O|�<�炂�56�����ڜZK��Y�B
u�<� ���	�&l�2YB�U\�2�"O���cD�2)i6����&gJԨ"O6|�F�x���P�M-N�6C�"O2����
���⠁�bp�X�6"O�DȤg���Ȋ���;G`��7�|��)�ӄ'�PU�ˍmd��˷�H>�(B��,yθ�ɖ C�L���ʀG�/R�B��7�Z,�� ]!�켺�H0��C�I�	�Rp��NT�|�h	c�:]r�C�I%\��y�"~�8�@�dv��B�ɡ_ hA4��`�J��QHS��B�ɶIT��/�o�>5� B v�<B�	�Hd��l��mx8�IF@´B�,k4���� (=�T��,Q�0C�	�AB���T┦#$4,2�nY8#�0C�I�_�}��"Z$7"�ZtN�e�C�I.8;�k�)L�)�K �n��C�ɅLX���7�[�G�|y��ž|�!�䙴z���2o��߶��vD_�m!�M�;��(Q�/:���_ �!�Dֻ�R���
[ͼ%R����!��ȓY	20��@>0^"���,�#F�!�ײ�x�B�8cpvh�lTG�!�D � �"f�~*��j�!�d@�`��BT�З#FP�2)�(�!���MP�����LKx�`��!�!�NJ�0����$�n�i#���`!�X�<9�h$�˶��R�˚��!�ĕ��45RI�Gޢ`q�
�&�!�$�X�8ڒo`+��*
9B�!�H�o��
�eC3(��HY��!��������+^*�!2���-s!�Dډu�Q1���4%K�N��!��u丼�$�ؐo�h��C�xm!򤈪N�j쫇��2~>�j�@�8�!�ό~~%��ס-f�e�P%�=@�!�d�(S/���T�XIv։�q	p�!�PA���5�,V^�-�d(�.Z�!��G��P�t�L�JK�5H�5<�!���d�w�}W�TA�aX
u�!��,���
�#F/g@�Q:6�_G!�$W��"��A-��s���;G�!�*���(7熃,r�<QnR:�!�WY�����N�8h|\գ7�>YG!��	Ħ��@�[���+���Y!�$��!
`4RS!��[B�����X�!��u,��jǽM���"f팅#�!�d	^6�<�a�@�`�;s�(+�!��
+Μ�"�_-8V����	�(�!�$C7*XZ�e��-	p	�эݡk|!�$��@��j
�,;0-Jti!�M�x���փ$|���=|!�dB�4�t�@)�He��&Z�6�!��֭\hT�%���Y�-Q�nʩ5�!�$ϳ]
�Z�з�.���U�!�D�;ef�����$8d J05+!�D�+��}1� �'II��CB�o�!�D��<٪ �E� 2\H��n�iD!�d@3��I�^j�]"���Z@!�`3�H#0�؎�̢�FK
yhB�I�&e��
�.�H��K�ƅt�~B��C�f�G,q�à
DX[�B�,8{*P�R$��M0�e�r+xB�	�z�$�A�K�F�}��e['EVB�)� N���H�:��h������"O��)�-���6�Hg��	n��T�P"O�9A�HN
�u3��ݬD¤	b""OTA�@��-hb:���K�X����B"O��qG��:�R�h��b��	�R"O0�`C�؛*��1�8V�,�W"O<\� d����B$��zF��a�"O�]�f��S�l�9�A-Hu95"O��褢�.�(���F�Li�"OBura']4���=��M��"O�f,X�6�Blr��P�G�|-��"O lYW��4� ��|Ժ�ѧ"O4����o62�Sd���M t"O�5����5�@�)qi���~|�D"OL}A�n�EHƅ2E�F.*��u�"O8$�Ƥ�-���ɶg5C� ��"O$�82'�.L x@iB ��Q�"O���g���BUʂ(ƅ_����"O��RKe�`乲�Lgj��z�"ON�����2X��+�	E<Upp�"O�q��`��}�tW�qq�ѹ"O&I{����_��-��G͠jEb�	�"O����I!~�1w�V
�"P"O����,�5�Fn�]E"O��q��>i�*�X�o:]:n�K�"O���2�ڤ+�}y�i�*R�*�"O�� P��e�(�JG4�@=��"O�S��̰ Fh*R'^<E���E"O�}�ǯ�}�fb&a� ���2"O$�9�kR�0�Z��Q�_M�X�@U"O�4��/7GT=����`}(�c�"O�(��o�A��M%KӶ�y�"O��'�� ���Gɱ%s���"O½ࢊB�/�`F^�I�.�!�"O:���AڢP 9:�NC/6���@c"O�0�ͅ�-��(	�-�U%��1�"O���5.�H1�����QD"O ��EK?=�&Uj#�G|���Sa"O�� $8E̪����4�9�"O8�)u㊕y��ࣰ�I��.�D"O8]@�݌Oa�ͪ���A�>�K�"O*����L�?��1&K�q���`�"OR�@�Ӳ+�0)`s]�!�"O*؃֚S�U���?I�$�s%"O���7 D)9"�|زe��|�&ك"O��bC$T.XQ ��&d���}�6"O��b�e�2wn~lxg"5z�t�h�"OIs��A(%��Q5�N3o��c"OX�AS���r�lXC�NX&H6"OF0D��-�����O����T"O@���a�lo&(�����x��&"O6h�H;���tm�R����"O�Ɇ(ӳ>���DmUf�~���"O��FC݆L�ݘՉ�K:(��"O*�3��H�*j�Z�Iӿq�D��"O�4�5�ʖ\.*I)p�ٰ��L�"OL�їG�F;�Z���\8��"Oԁ����$�<��HF!t�1W"O�1�"R eR8���۠I4���"OB)��ʨ[�0��Nߞn���qP"Oα#��
|���3�-ܢa�XrP"O¼��kP,�-��ٖ!h�BR"Odts!�R���,Ʌ�� ��i""Ot���>j�^���U��)��"O� ��hǄG�`	⣣��Q\�{@"OT��K:����@�ĳ/C��"5"O:��i��"ul�ː��+p B�"O0���K���1Unȭ4i��"O�K&&��+���آ8 -��Xs"O(����A
9{Z�B�@�r yI�"Oh�[�Z[Bp!a(�?C-4!�"OzI�!��8��+3.˱:�H�S`"O"-	��.�* ��N�n�2�"O��E��?��T�SȀ�,�`"O��qCg�-���`�F�VL�"O0ui`�T��d�J���+�☰"O|�	E��"H�:P��'
?k��9��"O0��! �,bx���f�>�9�P"O��:sOQ���$V"s�D�"O�)*�$_�2 $yQC.����"O�	�v)؆r6��C�R�u�X��"O^��S�β%p�:Go
)$w�s!"OF����:@��1�R��]ї"O*7�8(l���En֋oΝ &�#D�4��gΨH��� �T%>< �Y��#D�8a&F�7d�D�4+��'���5�4D���#*�#qo���H�3@��x�3D�̹�)7<�`,�h64�|aiw�1D���I� %���ĤslAS��/D�\��(̄I��I#�n�wN����-D�4	���c'�#aFB�f�$���,D��Qr�M)�F�7f߸$;�X��+D��GJ�"%ZDx�E$��rA�Љ�e(D���SF�D".ɰ�D�l܊5��� D��O>,�ƝXC��:�x���*D��pCLS�hz%��I�mV<ͣE�<D������	��b�/�4}��<D��37ɂ�HT�� T:��%���8D����׍Y\�m��hΚ8��9P%h8D��s�(��A��p��Acg6D�d��
�����5&��5
:D���w�͙��I�a	��t�U�E�;D��@ԫ->���7'�qb�IZ�%'D��CǏھ!�(i��ɢ/�}:/&D�\��ꕝI_(�*�j��#@VB䉏D���rFK�$��90ϔ�+�B�	�J���� `�	'P�4j��H�C�I%K~��F��:d��G�Y3�B�	'X���m*A��j�|C�I�#q$UZb�W�}&�1	�&��<ZC�	�ob2Px�خv�5���E`�C�I�E.p�yV��&_h��Y��B��4C�I�@�j��\�FN���_�r3C�I�ަ��7�Zl�t�Ŝ1F��B�	�\X6|`��N$Z�dز ��K�B�.h�4:��Z�{�zl�E�[���B�V졻�O 4�HT�b��N��B䉔�@0����7M�:t�w�V�MڄB䉬��f!�Be�?y)L�Aq*O�͚O�!�qisD|���"O��Pa�Q�����U.ظj�A��"O� �� �/EҰ�%C߄J�!�!"OJ��(ٕSR�5ءaF��h�"OVY�b�ϡ}�n���@�$��(�"O�%�Ң��\��p�!7Q�<��r"Ot�h�ܥA�H���;q �8�D"Ohĩ$"�3��!�C����'�qO��/C&"�X�rI��1��A("O�  �(���m����2���`��'�L��'�b�٥(�A�����C5�=Y�'�9�5O.���H�9�|*��d'�S�Dʓ�]\&d����A��h���y�#S��9�TZp�� �T�/q�<���O�(�-Oe������n�H���I ����!�[3Q9�Ţ0�׌�b��Y�hc
�1�2�4��=[��2@�)+y����Ñ��'}}�'|��#H$T]��S����z���H�'�&-�\��؋&q�Ɓ��OTY��O(�	j�Ӻ;�O��36+�3I�h�b戅�3_l�[�'��U�s���hy�!x2œ!F������'�ґ|"P����ʑ!G0|�D
U�SaRh�cVh�<���E3'�$){��&~��x�b�Za�<� �&�,����׼cK\Ը��Z[�<��Ƃj7�T2���yl� �,�Y�<i�E¥BP��Q��8I����eY�<)"�ҰV�2u���\</�B���S�<aL�%����9i��;ui�P�<�f�dl�Q�v�̭8�:a�$!�$�	O�$aA���T����)��k�!�DK`I� o]�h�V�2!�!��˲=�R��Gtԅ�s�\�j/D8��hO?M��9N�$�H�BѧMڢ��U�#D�p	�Ƕj�� �φk��$�!b7D�D
�gH-�y$���G2����*D��e$Եv0V���@C�sh�ʷI)D��Ĥ[�3��(�fj�L�d$�s%%D�p�  ��sž���6M�b�r��5D�H�s�*�`*��b  �))4D��ҐD؟+|���ߞ=�
 Ò�p�E{�����pB� E�:�Ą%-!�D}���c�ϥ9��y��IݪW!��(h��d�3�&��&��N!�d�6jB>�$�&j���0���n�!���g
�51���,�rf��X�!� ���ۦ�L(x(ٛ �ΏC�!�Ԕ|�i�筇h�����,^�	s��0<�I_ʺ1Pd%	�@
��$k�<�% �/\ph�3G�H�U�0R�e
릑���/�T�d�J��N�Ť=cBiF#C�ZP��6�q��VP��G&էg�D�'��~�#w��IF��^~�p��Y��d5�S�O,�A�BG n�&��B�L�a��Ep�'��+�ߓ<6�|	����T5����>Y��	��t|p��PdY>Ti�V*�	F�!�&�>,��gڟ�Kѣ:��p�ݴ���1���O�@A#��a� !��Ȋ2�nM�'F$ы���1�����gH-0A�xS�'�д��	
��uA�`ԛ'�LJN>����~��tR	�0,U(H����ȕ�y;<\�� �K�j����RKD��R��<a�O�ܣϓp��@gٖ���9��$Yݴ��=t��ifjݝ_"�-H�	�yr�Gx"�'���X���1���ׂ!H��4���d>��UeC-Iش8O^3	�(�0Pa6}b�'SP�zg��G���ж�M�C�f�9��?	��:1�ѡp��5ͺ�Q�g��k�!�_�z���j�$�@`�4p6�N�+�ٟ�'��;�Oq�
$z�H�]��dCr$P�M��=A�"O����♎>��<k&�0,��,;"��3LO��x�
�+I}H�Sdl�(%l�q��"OL�l@�Q�dЧ�U�`ܩ�g]���I�G��ʁ���fL(�Jː*��C�)� vh���ùl�����Yk��	tX��Y��[7D(�(&m-YV8��.��1�O�� -a��� qo�; V)0! $�\�f�E�^��p��Q�H�Kc&�z��D�?�e$څ|^x�K#��2�4ъ��L�<�#�U;]l��@E�,Z�D4Z��dΓ�M�O>E���d���B��H�&�2���J��'�H��?�͟��J8jYP�dj2
M��֞~���'��&�'���3k�u�q
�͉���a��>�e*�>�N|n�?'v�,Sp�)!�U�ƍ��l����ēMj�H���؀"N@@(�nLE���Ml��u�=q��T?��r��.�
|�&g�g7�A�:�c6�I��P�p�圜`��xT����84�x��)�S�9�ؙb���-�`���	��b@>O���۴�ا�O���t��0e�`�+�23+�y�O����5**PK����Z8�D~�Gx2-�'�?��w���d�ЀII�58�Bʇ:��ȓ�6�8����+�@D���T�����p��>	��3�f�r��AM�Q9D$����
���ȓj�Z�q3�
�;fE�p��_	�@��O���G�*�(Hb�/Z��O��@u�u!(�21��/����Pe3D�L�� ʗs��yu	��P"��#0D����P��8p`j��a��� /D�dY���Zc��` �]&t���XAM+��6�SܧVJq13��};�B��5A\Xԇ�A�&	��d
��J�ふ�(�Gzr��d�O-��i"���x��2�@83�4��'2F1÷Q�h�x��B�G��4ճ
�':*��'��,}z�;�A]�t�މ�	�'��U�T-S�$�z��T�6Mq��'�p��K;3�Vp�қ@�^5��'����%�ʢb*�<�D�)@�f�8�'ˮ��D��i�z923 �iD�Q�O���$߉j�X���l��&�.�Ԡ,�y$��asCnJ57��Yc!��~R�)�'n:T�b�J"�� S�ɫb�BL��ID�k����D�Eh	�eXe�$(\(�ȓF���c�<A7X��`�Y�"�����hO���`I�/ԨxS��������T��DR���'�(��`�پJ��5#�;6 8��'� �C�Tٜ}:E�92.`x�'�*��1ڬW߆0����[�s�'��,	�)��p�왻������0>�N>!WG!�H�3��	W�F�zg��<�'�Ă�-��؆C�8��S�Oq}g?��(�9$P�-4��R�S/0�����"OP����L�o�D�������'��<�	�O�8{��H�cG���Fįw���/LO"�`�ׄJ�[����&�@px�� ��>1��-�b��$'��3��C�&T�J����8b�H���$(=��ښm�TXb"O���QMX)?�`�6nC�U�ݐ���d�ڃ��D�$@q�%Ŏ8`�Ҍ�S�<�6`�F�8A�_�$H�-�t��<Q���6{�Ѣ��
2R~xx6NO'��c��D{����P"a<8���?�$������y¯�+a�� V���r�|�"&���y��/qGF��'X:w���!gk�%�y҂�q~���T�E^F8;�N[�yr  ���3�IF�T��X٦ ���y�!H��#*�Gk�A��V�yr+45P��"@L�.D201)5g��y�̖�r��a����>%"T(J�7�y
� ���#�uZT�ħߡQ�����"Ox]9�D��b�C�ĝ-F���""O�Ȉ�,���1���N4Xa6"O���dl?��(d�9�1H!"Ot�S�Q�:��eH1�P�U���"O��y!(A�4����0�-\�r��"O�����k��P��B��zG"O^�S KF�Uw��KDIQ�?� Y"O���G0�[Ղ^��ڰp1"O:��ЯJ�j�`�Ȅ� :��՛�"O2e*@�B�\ܰK<�fl�S"O�]��!W�/�0��-ʭ0��<�"OACU�^m�Hs$���1���"O���U
Ĳ+H$A!�ю� "O�e�"���DIpӬ��VÎ��u"O�]��'�:F�nX)�+P�nI�"O$r���j��݊�)|����"O����:��H�$�)cy� '"O�b��E/4%̽�6I5p
�"O���Dbϧtd\*���5@���"OB�K���?A4ؐtȮh*�At"O�$��˩Gz&�j���v� "O.%ఊ��l�\���j!�i'"O
�§�˘24v,�hF�r�us�"OD`�
�z�`�f�C�~�xV"O���'f�.�0hӲ�&O����"O��6���e� R�-=��B0�J�<��
H:`�h�@�pN���G�MC�<��@N�?C�$�I� 3Zt�v�XZ�<�#D�>?~��*�o�1��bX̓`��s��;M
���=w�t�<)U�S "B���^�xTx�Z
Q�<����G���-�#
U���T��O�<Qテ&ݺ�`��5����f�@�<a����Ҍ��Ѵvʍ���@�<� ��&�{Ӈ� <�āp�<���Y�B5���׳*V�e�3-�v�<�v���p攕P�Ƃ�wvL�ѩ�K�<13 �/m"&P��NZn�! fN�<id���Ԥ�>p6�Q�VR�<A��9 �:��\�2�����K�R�<�t�Z� �����y�6u�4�QM�<�C��T��K��K���{S%�f�<�d��P�R���Ki081[P�Vg�<��E(\��}�D��tJ<3���D�<����$$ �X�B��r �A�<��N$(��SpC�P�� �`�Yj�<�
ߣ(Y�@��@�
�y�g@e�<A���VTllá���r�J�a�+�a�<�剓>;W����Ȟq�l@��"D��3����$�3��pVp���!'D��3`ڕN��r��Ȉ	�Ppq �%D��W"Ҭ	�n<����TB�r��%D�Hy�o��#ΚQbpmF��v��M/D��"�%K!Q�TZCÙl�^ҁ�0D���Ug�m��� A+{B"�.D���Ɠ	2m���9o~	�I/D��F�V�H	���� 	Ap;F�-D�$��+D�g1|�q����&�[��*D��������Ul�#m7ܬ!��*D�[TQ/X����.߳2��J��(D����혋u�8ys4�V��`�A2D�0$b��+]�a��h�H��ԛC�0D����(=7�yc���7IJL��0D��`��w#�1�u��.P��D�,D�� ����C�%8tY����L^�iv"O��C��Q���� ��_�`�( "O�)٤�&S:�q�`�4	���"OR䠳�!�Ψ*D�*���H°iv0#�'��	rC_�cd�rǋ�\�Lu�(���2a7?�s,[�xAXݑ�GК~Dp�+��Vz�<�!!Ö9:�<��	v �+��X�
��9�c,��A&�M5.��TrA�;u�=�"O�TQ��]H3��b�!�I�"81�䈗V�qO��#��Y���DNݫ}��"�$�)ۨah�M2D��ۆ�M8l�fbt�+l^�X�>lȨ��6�O���*� __�D3SiR�m���'��H�da�A~��G�<z�Z��O�tP�'�Q���x��-��!��l��	��a+�+f��Z�x�FV�cU�O�On��b,I.A0v�v�T�# �9#
˓]�n�S�.���|"�  !(�b�P��R��'!�$]-���@n��1�a�F��%���VhZ�[6qO�����"GƷp�`<J��m�PE�V"O�(�b��Ey��FI;d�%"�,�	��-)��L<�Q�H5>��k֮�$�f4(7��vH<9"-?ԨhI��M,Uba��E�9ɖ܃0�*�O>��d�_U�`	���R$���Q�'�D�*�K�M�I �j��aD<1U!�$�!XhDC�	�2�\u`a̞��l��
�&��O�`��J?�)�(R\�6��[�M����P+B�	6Zժ�L��A򋝷V�B�I�^�F�ߺh���5↔r��C�I����b�S��";}�C�7s!L咒(d���N�(�C�IKe0�KV��0c8t8׃�G��C�	8��{@A�� ��@���C�5kh�Iq�
6�8Y�	,A�JC�bX�{'D��q��ATIG�#-.C��ol:8P&l�j����BB�I�n����ٱ��	��ЂS.bB�7�P\[�J�1y��ce �׊C�	�H�]0�Q�9!H1�Ԃ�Yo`C�	�.�o�;FR\mKB��e)RC�	<�h�aԈ̕e�\�8dmA�(C�	�7�\̺r��t>���� ��B�I�9a���ҥѤ|�{b�"'�B�IC�b1�FG�-OX�������4�⣓�5��?M{a�`y�,�7��5�|]��"D�Db�(����Fه"x��`_��ؠ0�|rO?�g}2g+4J�D��?K񌽠'�,�y�]�)��񨧭YA��L�fD�ڽ���yܐm ��N��0=ɳM.^��e�Ee�"~}�|�0�Fpy�-��T�����|ZwV^5�wO�`��ͮ5�4�i���+ ����'�҃0�P�'��t(�"E�k��+�/��h�!���01V ��%����X��T�8'�b�qq�]�<&�=A<��v��S�	��/F�9/a|Х|3�Q!'^�_Z�)�E�]{
	ӧ�Z�t��Ј �T&UP��2~_��a��JXT��e�~�B�x"E9z�r�3gۿeI2�6��э,��ں��<I3ޱ�'�^�&��i���	�@�	?q�&iʠ$S�R2TԠ`-F�s7�$@*�K����<)��3c�D�%/ "D2���	�0��%&n�5[�*1B�d�Z����3a�l��/�!&N&�ɵi5��%s�?����u�ˢS8V�(�*��u|R��Y��(2�7u
��T,��t�D�Zӫ�u�RLXs� /L��1��E�6���׈�4r��,͐r�L�3ًs�@\`s� /q���2��G���4bU��#x����D�~��@N�|�BE����JJ,���jg��qPR���v�m��D�;��0��"H\r'Ϛ&KL.����	�g����ٓ�I�a�ҹ�N�*V���8$FX%�c��9&�:n��zg9�L����?E�D�Q�e{HQ���_�,�#�$\2�y#6g��:ޕ�%o�?F�|�UcX�cw\M��A^� �sԛxr�'��lذ%�"k�n��&�J�Z J@2 �]�1���:k�<��'��L�e� h�j��<+�n�1��Af ��VH��Ni�b�	Yol�(4��o���)�$ΐ��,3L�"ׁg��,�PC[�_���2��)ql0&H	�7�����*,1B�B�A�g��,l6� |��FQ
>ԙ�'�Qf�P�=]�6y��]x��@R�^�^�:m����؀ �	Sd>�6	�B%B�h�|t�B ��1D���h2-^0doZ�[蓦ɾ5z}
&�
�o�\��0� �?qX#V;M
R�4.
	p1�� ��!�r��fl�Ojf�j�'��nEr���n_>GAP�I���)ts���D�y�ըH+0/2�
�n� ���.?DF^��'1.h
�m	2*�W,�/.�LM���Q��0�B����铄5$|"�k�W.*Xh�#�!_d�5	W��	���Ae�1*)���]�s ���o���k� �6��j���%���'�Zh���]��)�'�)�^�n�;,�=nG��AS�V3{]���G�-��	�d��k�(a��pE����i�&}��含mV��OI/|�d�4F2a�� B�0}r	��f�Ʊ[�D�}����o��1�8�P��vܬE0wBΩ��yK1�	�5(4�����rڤM�~J�G[�X�`0
��S�G;�Z4�̌@p���%� G�.�P�C� D����Ox����<���&��ƍ�9�z	�Ѩ��[�������+ݹB�:&`[*t嘨��g�-U�ԍC� ��f	��"���-��J��'�X��w�@-V}�%��5ΆP�'`%(p
ʌ/%��Y�>Ap�T�XZD1LI�P�H���L��\1��y�G���(��2k�I�b���5���E�S��~	���Qي��c��1���A��ӱ��bL-a�¥f9f�R�9~��>`�gّtVdk7H?7*�x*��/ʓS��80g'X�|Zt{���o	n�r�@#@�}��,��G�"��L��.�
0
t�WoO�z�D�𙟜��F_�xE3Ŝ�ed��"�)h�=Y�n��PWƑP.O?��Ӓ=�1{�!K�?Ḅ�gMZ:)a�#_��8�s��}�d�5��U0@��a�C��6 ��)�J�>���X�\� �l!�	�]�(���9T��z��0az�pV�H5X�|�`g�-��(3�'W�Y�b��3b���a϶~/5�U�Z$6�����V�zt`����8�� ��׭dl�ȰgG�|��&��p�N��T���x�@A$Vu�<YW�-F��IP�I���@
u�j��R0e�,AQ)xO�pl�����y���Z�:��+�(�DA�����y".�Sa,���
�UG�������j䜰	e&+R��`h���a�Ƀ��T��E��f.����&�?h�bxc�6A��~�2K��pA���q�"R��X6�,�B+�u�<r�UZ
a{�<20&Yڔ-�+h���ܩ��O♡ai��n�B@����x�ZIZa��������
�$�g:H)�"O�=��(�"��s��nz� Z�<��bL�2�Y��`�mCr1����G=ꌺ`�B$*L,���C7JrB��*@*z�(�a&��UJ��@=0�b ��A�.O����Y��xgOٽ:�,؛a��� �:�Z��%D���$M
��s��?��0� a�qՔm�@�=����,`�vKƶjWh!��Ľq:���C�4���@lڗH̙���ne�<uK&eJjB��/$�2��& \�̌L��M��-Lc�h��K�G����@���4x���_5���A!�z��C�I%^ <d�͌7
�Ip g�%+�R]�%��&k�ΒOP�}�j<�c�lΩ�8`A�DN:oq@����Li�f�U.,*�q��;G�*�ȓ"�(@�@)-�̵H�FF2|jnu�ȓ � qU�
M��w�W� ����ȓ���Z`�zAZ,���1>�\��O�T qO,�}��l���*cx^��]�TI>�ȓx�%9��8�J�#�O�<+��n�%�
`�B�i8�P��D�a���-��A	��25b6\O�ac���}�F���'��b���1$�������Y8���'A��9��_�x�噲��َ�!�{"LɀhM�8J�MA�O� �`��;Uz�2 *�� �'�����Jҷ)]�F�ζ!����e8�*i�J�����<P��̆KT%^,B� ���i�<��NI�kw,�8򌒠c?~�  j�X�'S�&�"��(��(�&�ްDA0� `V���A�RM�Z �E��y���in�9`�W?R~��0��N��yU�?�.J��L-��K����'����Ņ<�b�E���!���(�/�F�Z-�pjS6�y2� K�n}�a�Ō0Qh�{Gǉ�rL��OV7���b�Q>�|�����b����;Q��хȓ~�����kd�P��1'�Z�mZ�bҚ�K�!�L8��b%�\�i� i�BJߎ�S ,|O"�ԭ������=ZsV��`�ζJ�	��}k!�d�5^1��Ǉ�q�M� *K"o!�� �8"��U+�RQ��r�n�3"O��� �5�TXJ%�M.0�8bC"O&�A3e�S^J	*�͕�-���S"O��FG�|�3%0�*�ѥ"O6� �j�!�`�wn��@�@"O0�z�o�;�] ��� i����"OJ�X�lO�/J8T��� ��L�T"O�dK`(^K�t}��Ͼ4��,��"O�Q��S�Fs��9��5�V�а"OT	�����ĈF��0�d�"O:U��_Nj-���y�4���"O&���N�M��V䍐C��-j�"O��JW�Gk2�9FYAR6��S"O*D��5p��	�@Kj(��"O��z�ƀ>"B�����"*TC1"O*x�
*D4�i��3"�|<��"O�a7���x�ɑ*Dd�:�*!"O�-(�k�&(���Y��w��l��"O�l�f��&(C℀7G�&�\)� "O|\h�#�b��� ,�|+&"O ��2,�7!S���
��8|�1"O���`�1-^޸J��d����"O��� ߁N��E���>��Ԓ�"Ob��c��CN^YH坫Y@�i�"O��@"�c��l�Cˏ�G��\��"O�Lv*K<){��Y���8�����"OL]�]�n5
��掹1����"O�ܢ�4�b�H���!G�����"O��H����>�NE���7BK�؀�"Oh�Q�.���d�aOF)S�m(�"O^)bU�N WVX�2��	onµ{�"O$9�7�O�J�}f�8]f	i�"O�ap�cL�5��H7gԓH�B�H�"O�%#�H�>L��Q�2)P��|�{"O*�9�+�~�ڐ+R�Nº��R"O�pF)f�ȸ�/�@�|��"O��3�R1+#1S�v�K�"O�U1pBD�FW�d���N�bx�|s�"OK���=�ѠD�ie���"O��h��O���H�U@^@����"O�dH�`ћr��lbA�N=v�\�Q�"O:�r.W�����H�;�J��"O�D���i�@�cMW�>���Q#"Oƨh� ��~:­��L�>�4��"O�Vdݫ)%��j�?V|�S�"OR�q���G��H��
zf"Ovq3"��	�,�+bi��ڂ"O������7>|�*&���`�"O�9�5�`a�	9\�:��iW� !�ě�B�f��eG��.���v���#-!���)��@�C$Y�ڕ���7!��H�����>d"YC�o͚C1!�$��6]H���JW#F���ڝc\!�@�GU>x�qo��k]>p(��!�ą+,|<�b��:Ui��+�N5)�!�䄔��ɡ`�V=,��-ΚE�!���4w�xCV���b�LqslƎ&�!���}5�����t����Gh�!�$ܷ\�Б�tȄHF�D����`!���Mt k�A�H7���u�!�D�n��ʓ)�<@֕c�c�: �!�� �2	��)F�i�*��0���!򤍴�Yy�N^�^�H�[��Ȩy�!�$V3*0��b��D&�E2�(�6nS!�� ��!��-�.� ��ڂ\K�"O�(��	�V��2	��d�s"On�� ��|����3��6~����"O\d��i�N�hr�$d����"OԹ�>�� s�D�0S��"Ov,(ԧS+eu��j"�W	�0���"O��#S��Y��$�#A+5��#�"O��	Fa��X�ZY�'"O���r�"O�x@�Ì�;�T8��8Eyv)�a"OT���Ɔ:-)�n��;f�4�"O��ycj�9	���.�����"O4�+�C�y%چF�X�.�:F"O�p�r��|碥��o�7�$���"O�H0P�Z<�#X�4��䁡"O�Ly�Díw�n�����6��M�"O ���Y�S:�l�˾���"On�1���� QJČ)(�^�p!"O�H(��2" tԘԬ��+��\�"O6<Q��¸�u�2��%�>�"O}[�a@2z��P��	�/K�*��"O�m����g�X�4�
"{��IZ�"O胣�ѦO��5`�ۖ>�<Y�"OX��pR�e����	��LUc"O�9�#�X�%j��G�3�N��r"O
q	E�G�A���# P & �"O����➖@B�q	���
	���"Ov�3��F9�~,�A&�
�i��"O�`:�[�,c��S�/L�u�T��"O�L)�E����Ϙ��{4"O��G.�)^����qM�:\��"O�5�vFF��0��NR$��"O�IPӌلPUً�ʄ"!���"OJ��6%��M�|��B�_���Z3"OT8��Mdܰ��s�ǲ-s2�R�"O��˛/@��ї�_�
KDd
�"O(|4��0�G�U4;�X�g�<1g�"S�H2˂7�l�pl\�<��ŝE��3��KM�T�
���f�<1���dk��g>1kr\�u�FH�<��
De�t��";�b����p�<ADf�5QVLK��`� ��͟r�<1����z	jE�PH�$��Ēw�<Ib�Q���X�&%��+�F�h�e�<��G3q�h�pD:$�^L��-x�<�7��!_�$�U+I*[����⇂u�<��l�ր���ռl�d�f��l�L�h�ō9�'| ���<�TiAN�',!^��Z�a�U�%��1�	\f�v}Ұ+�^�OtuF��O�q��o4;pp)`����jr"O��z��Q/*��ڴ�K�%�V�&�ɨ&���Т��L���K�'�0���>Ro���V�D̴.OJ��f�9N`�O�ۙk���L�c�:	��\*2����FH��X��QЫ��dP��d
��Hg�ղy�c�\;y�$�"%�}�Ƈ�:r��e�"��&�+r�Z�my��Cg�x�}X�-9x��e�C"��`Ä-9�O9x�G�&m�20�f��p@B��*X� r@$�Āԗt� QI�$�O���JB�DI	BiaWJsEF�O!�O�𱳩� |���ǇZ?Z�Z��R���#�SD�$I�O���hM8��P@��9zNu�5f� {MA��h�7(���'��&Xo�=�$�DX�4�F�^3:���C��Rj��
n��)��-�g1�hI�AƐyШ��^29��IV���W~8���k���¥�X�D�<!�BB�j�j!I/]k���ȗ��IqƇ�2�@��v+G��t)�N�btVCp��)k�`h�����Yq�1 �T���F�
�k��Ұ u�˹k�HR�.ٕz�����'H�9�r��7�V��j�&(�ja�!R�Rd��#b:vH���t6=��Tf�23���Ľ?��R�Y~�U�UP�}P����,*s@^���'�� ��FB�R�Za�Wq8R���O��:v��($�]�U��?64ɱ��јoӠ���Q]Ǭ�S3�-3����� ��9�NU%:�"�3����$,~%��*L��L}�S��0*�z���9�����$>�6�s�BA���N*6{P�+"+�'�VD�`��(�I��酊'�(q���zǼ��ثD��ث��E�6���w��?h���
�H=;�^tP�I�zŲ��FX�D�����)4���R���c�Z]t��;0�o	�x�퉹x����lC��9jDHEdH1py�m����9-i��s�F�WL�<S�޶t�Â6O��x�*��X,P��WM8�۰-�{Հ4�?	P/Z$ ,�P��i���̘c�	��E�
�f�L�1r�"���~B @7Xa| ��k�U�hᠯ�V� �3!�2A���������0p%J �9��S�O=�x��	�uZ�BS&ػc�Ų��ƃ~tlPJǰij�cW�\�ZU���� 	��h`@�$�d�����d,�	6f4Yu�F}�	28�!�i5�|X�'���X���6>6�p��"d�r�	��p>ch]�'�0�I�m�iR�h2�S�?:,t��Y"Ym�Q��}���n�U�M	���[$e��1xx�H�뇻{��k��I�D�9�%�5~p��~Z�)@�Q0��-.s7����gګ�1�E҉}ڼ�槈��䓄9�ƕ9`��v������7p>A��,]�:01J�y���'��fL�A��@�D��gΜM��'�کC4O�&B�Uc�L2�Keg��JC";��˗�Vp�:2|z�!�W�0P�}�@) ��"��y�f	Y�hL=e��[sM,`��I6|O5����.�|!a'm�A���c��> ��lXՠR�&�R�\���M����GB#��O�2�a�&7z��p�D�X��q��$�$�&�1bf5y��b?�0�ժe�9�Ӫj�:�e��z�L �0 �lj�G}���iY���� �),�p�*��y�f��
)\	���2A��M� �S��?q���֩���"�N}�aO�Z�$��F<J��v��0<9���&��&GڄLtL�*�DR}�GƱ;�,p�#�i�'M�=iaA��7��Q�Ϸ!,ԃun�*���(c@�y�����/�3����gEi=I)v�д{��0�3+
l�'}\����g�E��H�<����'%#� �H[%r�0�C�^��P������mڇm��I��@�1��t�o�0D���������
]��F�d@D� ݶi�6�A�-�H]+�Mг�y�L�a��� /�h]��)��w�
���'<�����W�]�N�PO?��>�F獏'�4Ec��;+{��2 %�]��LY#��49 I�#I����{@,�*���Z �Ѕ8��(��ڽ�*ń�	2�6�i��:0��"�b{d"?��i�"Y.ؑ�_<< �S#�ٺ#u
��?�v�]��\����P�<�b��N�*ĺ�k���BiOy���6R��#�#
&R0���|�OӴ+g��0Y-�ɲr!+@�xc�<�S�^)Q(�k� �>�2��ݨ=Y���<db�u�Q>�X�.� 	o�.�@�EQ4�p�ȓVݔ%��e�=4��@��#Ŷ�0h��ٳhW��#ꋅi<a{��;CL\Ѵ�W9<��a"֤�9�p=�u��9t��)�.п�MCu
�����(^�l�lK��p�<��
*^0i�C�74*\Kb�Pl�WŚLD+S*�z�}�����r�L��W�e���"Rf�<�c��q�r��3Kψ0�F�`� A ?4�x	goN�	`��~�ւ2�-Z���
+�F�7�y"5{ �u!Ӹe߼���O=�y��Ԟ=�T�pf@�f���)� �0�y�	Ԕl�`8p�;_Q�墁��y)S�,��іo?R��`���;~�6���?�I��~"o��|nmK�愂���BW�y"��H4�t/�7@�9�ɉ��M[#�Ad��Y�)m����F�%8�!��q��=��	Oy������!~��ی����S�	Y �{G��O�!�-z-� �m4<,V�N�9�qO�gQCld�{����QN�����
mk��V�&!�d���`*$a�f�(�[0�:zS2��Qa�'@�u�|�'7�rt��-�\�K�Ϙ��C
�'N�LY����{t<��=n(�(��VQ�5��ǁ2�0>Q����,��A�%G_	e���W��Q����'����I�S4ON|���@�\hqa�/ѯl�J��"O*|g�>�"���A�6s�d�w�$�8F�l���!�9����:�	��,x�®^φA�G#!D��+EL@���P�:0~��#��8Q�
L�J>}b�x����Y�)����a�ԝR>�y&�ÓV�!�� �Y"�F)a�t(�w�;i��iE&� u�$��|"��"u���F'�H��A˒��=�d*Xu�.��t��g 
��9��!�4I����ȓ�(}���s"r۳KN/T����8b`��o5hY*����]9�݇ȓv
U� ˠ/'�����s\���Ny�غ�Gܪz���;e�<RU^��t�BDQ���""~��`C�' cN���x3�\IB�
�u�n|���c�|���9�j� �❍v)\��H���ȓ,��]�p��7�l�� �F	�ȓ|��h�ML:=D��Å�j� �� ���r��z�J�@P�
W����D���� �	q"���վY�bD��S{Jx��,�Q�h�G���ȓ5P���j�*mzI�	�"mqn�ȓ2�1q��߶?�P\S��"z�dI�ȓL���Q�R�waɲ��X�EGh��ȓ�4���ѓz :�b�bT�^��_�t4�b%ATb�E���,4*�X���F���R �x��ce�,���Y�'���xT�ΚS��5�A�(�
�'��J�V3_G
��
ݦ2�� 	�'���蔣�jd��� -��+�'����qf��T�B" �/ ��	�'��X�B�3}g�9*������
�'�d}����i�<�Ï�;e`�Q
�'zq�r�Yj��8aF��zʌ	�'��Q�A �E>fa��EN�D��'�����L�\����ň>��9��'�<�y7Jʹ
ă�҆ �a	�']�`�פܛo.��УK*��3	�'|p��9�n �S,��w<�0�'�A���&[��3dS�����'o�AhG����\jqkW�p_d���'�8�)�扎p���PNޫsh49"�'�p���le�� �a�l�@Z�'?���+c`8ya!�0}�lLَy��O�z�rp��ϋ�<�A�fR���'Z��Q�|,�i !�7r��Y�'��ᢢJ.j�<��R	p����'zh��e�G��\=*R�����'�D���#p�+��J�4ƐH�'�dEz���Ta�Tb���g	F��'*�s҉[�a����v��'t�*);�'��Z׬��m�b���ɲ_�$<i�'�����;u@��"1e�Q�4���'H��BP�{�$+��V
Ji�MH�'�D	 'P� ��!�劆��x��'��"=E�@C�4f�0��>�
t!���gg6�Bs�Ocy¥�6#�����-KE|�ʣ�އ13L�X���{�xݺDT���q
�
�����O�8�ZF�?Q2��K〉\�����'I���1��M.���]U>�YR��	3�ݹ&�K�%ņ90���%��� ÝkC�|��)�q��b:`�8�d�m�����^�~m�%(�#�CJ��h�����������,k��Y!֬ɉ,
�T`��>�R�X�=�����/,r�9���4NҪa��'��	�h��Q�6,�)���5����g�I!B���t�:qp��+~W�*��<�)�'h��mA�6v�6Q�$mR�z�J��ȓW��@��3"�d\��������ȓ��0lɂp�V���ٍ �5�ȓN>�ٛ�
R�
,+�hJ�(5GzR�'�tӥ��?� �E	[�yg��'v ��`J�	�.����Hz��xp�'� 4a�f�4��`(�A�'r�ٹ�'�lKd���#6����HПǪ�	��� r��l�`"�Ѓ�{$�h�"Op<���=J6�0��"k
��R�"OL�4�Ű �l��'�#h
�uRP"O��b�ր �hb��خf����"O��btJŊFX$��C��f���H�"OVec� ߒP��P[��)E��D4"O���D	JMA��K�
�R��8"O�	���GT4:u��F}ϊ���"O8��@#�&�VI����&dv"O��
��'�貴�D�+�P���"Oh\9�jCb��5��G#<::���"OZ �c�]�0Q��fi� " -	u"O�	A'f�$-{E�ԑX�A"O$� Fē:�A��Q�`��Չ"OL�c�A�T̀� ��.;��۔"O�u���� ��4�0C{X}��"OS�&*^�P��"Ɓ.Xx�"O浑B`�2_�,�+���Ie4���"O�R��k%�ͱ��P';O�p��"O |�jIx���A>=��W"O:��t��8YÜ<i�l�+U>P���"Ox`�ע��ę�+P�x89�"OV
Q#�x�������"O �D��i���ҷ+�1`~���"OlmS��1}�� ��.p�dV"Ox�����"$����(��6i�d�#"O���&��;@�ذ��GIPf ���"O����@�6I���#���dW�@["O�@�Fd��K^�!��D�3cT||zG"O�x�u ��pz�!�<���R"Oƕ҇bU�~s��"� �O�N�y�"O"������i�/�d�	p"O�h��B|�H��%�HQJ�A"O@u˶j�>�N���7�b8a�"O.�B�&�yV�b#Êh5���"Ox͒���z���*tC�-���S"O `{!���^dꑄ�=>��"O�����#���$cEp.Ƭ�7"OM�È�2p��ⓣ�r�
"O��3��ri�+w�M��D1	�"O�e���P\�V���O�C�蜒b"O=���ڑ�����@]�� �"OF�b�4��������HՑ2"O�!P&"t�$spE>P�|4s�"O�x��iI7[]r�٣������U�!D�t� &?K�{`b\�R$��u�2D���0g�\����Y�k%���2"2D�����4�(d��'V
o�Ыa..D���f��3�-i��8������)D����C�)��mYↅ�.1bQ 'D���&��^ncf��:~if�0��0D�PQj��=�Ed_#f�D�I �.D�\�@E��WGd�w ��oO���+D��R�/N;/[>I��YQ0+D���a���7�ѝ��rPL�Z�<9І�j�����/ra���}�<�ckS=�K���d���fN���C�ə D��:��;MaPE�aI�8��C�	�^s�Sm�(J:Ł�-E�M�C�ɬ&�� ��U3E�R@#�	�D$�C���֐�pmW 2Ft3%��$��B�	%Nm�šd������F�T!�B䉃}��@��Ή|��cP��]L"C�I=3jd�򷫆t�����k�6x1(C�)� ��	�*!�j n+zy�@"Oj��s!� p�5��ְ�T%�Q"O�81파E6b)q�9(�4�kQ"O�-��.ΆZ&LT�}��U�g"O��� '�wj�²����8F"Oք�6�.�*��؜��(C"OԐq�6�yF)zZEС"O��x���!L��J��Z���p"O���p��=&f Adb�w���f"OL���A?:0ha;�c��i{�)�Q"O ��oX�]��<�C��:9�Hy�P"O�|���	O�8�c߾n���yw"O�遥��C�.T�g�Ό>�xf"O`�H�B
39x���H��t��"OX���-�68��B];H^�"O�x�pgC!n�V 	�CʰTiI"O�] GㄚJ����U��i��"O�$��\�c������)���4"O�Qy�!�'I� U���Y]�t`2"O+Í�;C��Dg6����"O
���M�9�,ܐ𭀻�|Hx "O���cD8)¤*���\�T��"O��±j�%b1<�{�j��Mf2��"O�	��i�2gbtY�L�Fk3"O��a�ތ{	�������H�8��b"O��x3+�Rw�L��Z�s~�YX&"O(�seMٖ �B�BaB� %��a��"OR=����,1�K��ŘVX- �"O8T�ՎK%Ny�5��䄨p9<=Z�"O
��ꅰAD4�z��S�+
pa"On(�S�:L����!	8��� 7"O�@�
ɽ7���x���Yf�k"O��藠
6�T��6Ep �"O4�󳮜�JIĸ�w,�+]-&!1�"O�\���\4J_�W�^�#]ó"OB����>/WN�9�,��&x2#A1D�|Js�Îo\`�˗�8a�TX��-D�t��	����d��`��1Z�+D��'N�RA�YАg��T� ˵)*D����T�2��礃�l�����(D��)V�3}�l$��hC x��`E(D����A��r�3�\�#� p��(D�����Q�i�>�k���:�zq)5n%D���1��n���
d�9$���-D�JW������-�H��(���-D����b��y�6᳖��h�hP1�O?D�$)1��2	�zLZcE�!�|Š5(?D����P�e,|��!R�d�zq��=D�t����*q̰c�
�%]��y��<D�|���45����������:D��7A��II�����[$����9D�8;���68u����3:�k5g)D�Y ��t�ְ�¬�<fQ��0�:D�|ɡ��.�t�$M��/���#D��xujɈN4ܫ��[�d��4�R� D�T;e���,c��)���cP�>D��Z�-T� �T�#3XP0�!D�8ٱ�W	�Չr`V�uzu1��1D�xB�F����U�CZ`�Q��3D��r��ڗ>;ne�fL՘GU�YZp�6D��C'O_N� �̔���M0u�0D��;��E*n��Z®ђ���@<D��Y�)���H,P�Q���w.8D����%AB��⨎<ƀ�b�;D�� �̳<����/<0V�\�"OV�$�#�p��͟�NFJ�{"O����{!^�[nY,eǖ�Ce"O��ᢍ0t_���Ae���#u"O��f��
ٞؒ��Uhc^C�"O�]�i�/`��"�HX�,q�m�P"O($�iH�E��y@���>7P��""O�!B#H�W7֍k�aUH�8Qa"O����K4>�
y:��\>���g"O�0q�	{�d�"����+xx�"O�!����jk>y�㘌}�:��"OȘR��tL�"�a��~�쳥"O�Y���[dd�j�a�!=��H�"O�8�6� �S��z���!"��q�"O\q��*�8<[�C�Tv�!!"O�	2�
;��A��c����"O r��.6r���,�>���Z""Oq37�@"zw�}@�j�p�b�S�"O���� �9�.��(��޽��"O�8�2�UWu�`��L�(7٬�j�"O�Y���E�0���O6�^� �"O>��3�M"}�N$��m����"O,)D���xAd���ǂ��"Op���E��W�L�ci��U�p��"ObD�aL�L�z���U F�y�"O�q�K^=pO<���ܲ.��W"O,)Ss�P<_�,Da�7+BM��"O�����4/�:;�տ<�0��A"O�ܺf$OT�S��Y��|�"OX�3*X!�V��EV9,���"Oz|��K�b�� D��X�A��"Ojt��3׶��AB��w"Oz���	T��pA��r� �"OHX� �ʭ6hJp�r���@��:Q"O�]�1�d��u"jv�y�"O��)!�^�q�t�����A"O�(�"D!z��i��C�6��Sa"O��ӇF�#qp��C�̿@�Z�iq"Oΐ@�DT-V���s���4)��̐�"O�M�c�R�?q�(4"��0�(	��"O��R�aĨ&,�X�A��<<����C"O��P��I�m<�[B틏7���T"O�Ԁ�F	�xW:3���[�䨦"O� b�h�1]�|H�l��)t��$"O� 2�'x8�Br����'o�j�<�nKTj1�A'۸'dD@�W�A�<9���:m�e�B��t?�,2Rf�A�<�W�Ʃ-��YIQ
�Z&�av�}�<�!�IgM����ĎC��KVgv�<QuLC<��,p�49�-�r��z�<Q� �"d�B �R`��#*T�<�`�J�rb�D�"�M���j`��_�<y�fQ��DE��F�<$�fLҤ$�^�<)�F�>���1'��Y[xE*��V�<���ڤ����Y�NY�����N�<1��N�m�4A`FO�)3���I'�q�<a�ID35 ��VKJ"����D�b�<�	Ծu<d�b`�K�l-���^�<�C矚]�TQѥMΉpv*��e,�~�<�a��,}�,����̉!��2�)�{�<�cR%/��a�"�ڼQ�0P� .Tx�<�6EU��~<��f���ybH�I�<��D�$H�H�r�®~th�G�]�<qA�Z�&-!헬 �̱� J[�<� x��K1M�!J��9Gnm�"O�Tۤf��!�̸@�<��b��>D����9Mf������x��C�d*D���u�   ��   �    b  |  �)  B3  �9  =@  �F  �L  S  FY  �_  �e  l  jr  �x  -  �  ȋ  �  ]�  ��  �  %�  f�  ��  9�  ��  ��  ��  u�  ��  *�  n�  ��  B�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�VO&}��a4/zY;�#m�����#D�D1���'�01Vo^w:,�U�!D��1G�;(�x���n�$X�6@?D�P�$�Õ�ha�v�C�y �a=D�t�+�p��xj�N9N|�C�<D�:�K�<M�N<ca��*�Ĥ8��9D���������%� .�7Ẕ��<D�L�p-��h�u W$�[Ri<D�������e��E��V).�&9D�T*� -5��dKq�߾{|��聥*D�\�t��J�9��D,~|qR�&D����O�RtN�I0�6S�L�jUC&D���f�a�R 	!�j�T���$D�d8�FD�p��a���t�L�b��&D�|��揺-����e�˳I$Z��A�7D� �Q��,YX\�;5M߾[~X}��5D�p2'����(��R�,�^)#��2D��"�V��V��7-V,�^�QEF#D�(!�c@�x��V#�FP�-&D�\:�英B>��aι�m��#D� ���9SO�ؠE�l��В�'D��x��̎j=*���?�J�A&D��Z%��.}> Jr`�89wQ��N>D��TBԖoƾp�1���HIF	!D��-�$[� ��T���p`��1D�d����S�����K�,t���h%�/D���Cn<5TP��޽2�x����-D��[#.1S���g]�?�d�Q��,D�,��'i�踰�E391`�֢/D�@�OH=�)��ƀ�M��4�,D��8V"J�Rxv&� +�4U��*O6�E��#Y���d�Ѯ8�*�HS"O�H��E�<X�b��hF�U"O�cQ�0��s�;-�q	�"O�P���,�.�8qe��N�% �"O��HE*UR�����]U�T#�"O���HIi:�֧�\���"O��[����d�@��2�"��"O�kҎ��.����o�-|�Q!�'�B��P��B_�TQ j��G�II�'<VEZ&��9/<Փw�׳*`��I�'ސ�������Щ� /���
�')�9�#�W�cp
��
тTx�'.ıRV�A�Ws��id�D�o%8���'�΀UBDE7�³j�����'�@	�W&ŬI���K���-!س
�'qPȻ�+Ӽ	��E��
.�R�
�'(�D飦�"�`5 W:�U�	��� �<(Ĥ�
N��Y��KUR��ۣ"OvtSqJݲ>,8�&��w�2|i�"O��S��^�@�
�5/ɬk���2"O�X	A� ]1앪1���
1�(��"Ỏ�F�>�`y��-��He�'@�'2�'R�'���'��'N�
 �A"t��I��޵R�0�{��'���'B�'���'���'��'��������)�/��{jP{Q�'�'���'�b�'�r�'��'�Qid&Ǹ Ub4�^�l'邑�'y��'�"�'���'Cb�'-2�'w�td(ګ6���I'Kx��G�'�R�'���'���'~��'A��'��%�B/�K�lX�5�!?�.8*��'�R�'�2�'���'�R�'�B�'�V�A���mО);�,ӎz��Ybt�'��'���'�'���'���'��Q��L1�tT�����.̋W�'�"�'��'2�'���'���'�N�Y�D�%�.A9 ��k\T���'���'	��'�B�''B�'ab�'���4��%%%�!	vMIx�J|��'���'�2�'���'3�'�B�'���X5 Y��N�3ӭ�`3x�҆�'<B�'�b�'���'���'9"�'2�p��f�_��Y{��JZ,����'rB�'���'r�'���'P2�'|�Ju�ݤi!����늏"µ ��'x��'�r�'X��'�b�j�����OtUP�GN)J|�!r�Q9���`&$Ey��'��)�3?Y��i`� �*�Ɣ`�@�,kx�С������O��<�'��A��`:�#M�Ι��l,[��'G�����ia�	�|RC�O��'J��}�f�<ܴh��FԤk����<����$,ڧ �ԝ��@^iۺ9�F��!\r����iH@��y�i�O�.�rP(�{fb��Xz�X���O������O�	U}����b��F7O|*ĩ�3"�L��D�Ew
�H�9O"扔�?Yt� ��|:��k)����� t��(c'w٢��p�X�'d�'�v7-ږL?1Oq� cH�GԸ��`�2r�|���0�	wy2�'*b>O��\"&!�2,[p?��S� W)�+ ?a��Q���NY̧Q���N�?A��W}~P�&Lܼ3��Jb#����ĺ<A�S��y��!�9c6O�3qm2��b(�y2!r�Ft�4��h��D��|2�IU80=x�h��\�* �	���<���?��-)ݴ���i>�0��U��u�3��O�E�5������K�=���<�'�?a��?���?Q��ۧJ(<�pwc�"s�h�ivD�;��٦�RM��|�I柈'?u���0Q 4��@A(�)t"�:*~D�'�7��ᦵϓ�H�����eZ�8S��@��jx����6Q�d��X�����ç&���I�Gĉ'.HʓPL�y���Ig>�ˇ��n4�{��?)���?Q��|2-O�mo�0T����ɽr]��6������部��;b��������?�+O��m��M��Ee栙�J� OӠ�Q$��B�n��+�M��'@��km=\b��I%�ӽDfk��-2T�PTm�-h�����l��j��d�O|���O���O��!�S�A��0�Pȏ�w�@��C�*0Τ��I���	��M��F��|Z���?qH>���~�6T{�Hξ'�\l`�R{��'�R������Ni�v��싧�R�(wL\K�E��;�ޑp ���(<���'K$&�0����'���'�	SE�7Z�(Y�F�*l�Ea�'tB_���4h�������?A����]�75\\�bh�n��T�FM��e��	P~��'��f�:�T>U��g 8y`ezB�� 6[�ѣ�]�&5��(��'�P��|���OH�L>!��N4
`���U�@�9�!eL(�?����?����?�|2-O��o��HH4m�qϚ��`�8�^:���PaFyb�'��OZ��?q#��xy�B 0�T�c
"�?���i" �ڀ�i]�	�L�P{q�O��/b@' RnPb���K�ϓ��$�O���O���O����|����5c���V���m�(�����ϛ&*��V���'3�����'��w�l1��g��H��I3I	� ���'���:��)V!ch�6�e�����	�7`޴JeE��N,x��{�M�US��DQ�Iny�Ob��j�� 1իS�Q�����0W��'�B�'���/�MS����?Y���?�폦z䒘���M<:=����mߨ��'A�IݟT�	���L�b`�
)p[�IC
C�]�'�|3��\,���[����ٟ�[��'��y2Ԍ���$��s�T|��'���'��'��>��	3fA$X���B&�ң/��h�ɣ�M� ������O���k�a��Չ;�m��g�s>�	ޟ�ɤ�M�+آ�M��O �i�B�RG(U���jA#	<r�����.2�P�O���|z���?���?I�U�X�a�V�h鶸�Q�Y7D�\�j)O��n/\ɸ-��˟���u�˟�ңˋ1�HP�E��iW�I�"�KyB�v��Do����S�'�^}��c�Pp�3��/� <�靤);��'Z �z�ES��L4�|�U�xc e��Il�9b��M��|��%n�����i�6��O6�4�.�ep�6��/-�BX��2%V� 4�v`O�$f�'��OV�?��47��O�|�̜`gBC��^�y��!�sW�i0�$�OH|��b���������� ���4b�.v>:ak%"ScZd0�$2O4���O`�D�O��D�Oh�?a����P)���%N�1	�����Ɵ�	�hڴ�j��'�?����;&9 â	"���S��3{������x2�'v�O>�I��i+�����w�R/r��C�YQ�z��B�_}�R�K{�IUy�O��'tK?J�镊¥`����u���'��I��M�Q���d�O��'V���ua�`t�:�I�?i��u�'[�ğ��I���S�4I��Ӱ�k�'�%�6HKr�"g�ԩ������O� �?u)1�$ˊ}���3V���;�%�f ���'mB�'y��OH���Móh!tTL�F)�J���#!H�|�NZ/O��%�	fy��p��#pUc�:��U �80�V-iv�����Z۴�ة��4����9����'��S/Ns�PC߉Ch \ �@��6��}yb�'��'�b�' �S>j�C�"�\,��*.���xY,<�nZ�^$��꟤��b�'�?�;PX)�ɏ��5#�
��7�i>67�g��֧�OTlP��i����o
���KKd'�Q#��\���A�����!�B�O���|���yȤ���F�N�⭹��S&4�v�����?y��?�*O�eo�S�Ԍ�	֟��I!#,e���@��
�2p�P�s#��?q�O(��f�J$��1�A�!vÔ=K�T(��08d9?Q�B)=�~��t��E�'0�j�$��?��ٴ�FĈ�=mpR��M��?����?q���?i��i�ONbf�� !���z$P Lp,rR`�O<@m�>[����Ο���F�Ӽ���Q��lU��m@�Mحz���<�r�iҺ7mæ�	s���e�'�`Ye�B�?a*"�ʿ#h*5#��:<vuځ�A�T#�'�i>�	���	۟<�ɷz��A�@�?V�ش�5!|�N��'��7-�'@��$�O���>�i�OX]b� r_���e��B?�9��<A���?YƜx����5w!�͡�nH"%FA+��ۼ"��ɒR+���]�QEջ��9�ԓO˓8�8�@�W rE�RVog,�����?���?���|�)O��nڧE�\���2� �d  �P[#�Ӝ�$��	��8�?�O���d��pl�%I�Р��И|�l4�f�E�Bl$9UJϦi�'
�$R�?Q�}���P�H�s�ҖJRz1q#�_SwP���?����?Y��?����Of�p����YNVHq��J2e)�Zٟ��Iџڴ`��D3+O��� �DѶ�D*W�ߣ:�QQ�HH%he'�8�����!H���mZ[~�h[�����李p�f`�Ug^�>���Z��̟�'�|�X���՟����D�D�G�=,��c"T/4B�43v����l�	by2�r�A���O�$�O��'j�z�xw�]-y���MY)�T��'i��M�g�i��O��H�eꎎO�bAx��!,�}�t�=�ʴ�4�-?ͧt$���P���*xU#�-

�V�H�KR�؍k��?y��?A�S�'��Fަ�p�[�}��Ѣ�7]@�D��9���<��p����O�űG�55�J���D4`�B�ODQoi��m�s~������Sc��H34���ǐ�Y�Tѩf�ȦG��D�<Y��?���?����?�˟�hE�V��.����̫x=���AbӨ��#��<���䧎?1�Ӽ�A�-"���֌I,A�=�tO	��?!�eω����'��$��o�F<O�;� �%+]���3�6X�~��b0O�\2ЅY��?���'��<ͧ�?�`.��Q	�5�� ���(H%��?�?�cυ��?����?a��LZ�.I . ���O��i��|��ޑx��9YW��DY����D8?���Mk`�x��@7����B�R�nX������y��'�*u�V'D�=�8݊�O��I��?�]
��_�M���&gV��)i� �'m��'���ǟ�H��5l�v1蠏J%h]�< u@�̟<[�4n�U�,OH�9�i�Ia���Vq���yZİA冡��lZ%�M��i�@���i��O�s'�+�j�LĒi��E%�	�Ԗ8z�T�2�|�V��S��`��ݟ4�	ϟ(3��K7GIFqA]�Z������}y���*���O��$�O�����dD[��	K�#G �����Y�dp��?y�4cSɧ�'q\}����i*P�0�J��N'0 B���1��'�N�BT�ş�!#�|Y�@3�]�t�Q�D'C.PZd�F��I�� �I��Dybil�:	XVc�O$Ͱqi�
e-T�0ʔw�\�`�O�$4�	f~"�'Ǜ�)f���U��ou@���C�"o�P%Ǝ�H�7-5?Y�`;<Et�i;���iʐ)I�.�j��w)F_�h��z�`��� ��ퟌ�IڟH���b�#�P�#�̅���
�3�?A��?1�i�رi�O)R�'%�'c�A��̆9�PHRX�rU6Oj�2��ֿ�\��\ǖ�n�w~�7KKv���R1U^t(j��I6J�f�C���ꟴS��|�W���$�	ҟ(��WrS���!+D�.�� t����p�I@y��z��z���O���Or�',e�AHЍav�0�!M/H��'X剞�M��iE�D ���_����n�͎I�gA��)��/7������ˁr�i>��՟4�0�|�i�i�,QH݃xK��W"]6w���'�2�'e��tU�Bߴ
>�M0o�I匁3#�J��Dkt���?���?���V�����0#�7x��%�5e`�x�	1�M��ʞ��M;�O����<��J?� �%@Ü�?�|��+	��X��6O���?��?����?�����I�,�$d;��a�F`���NRx�o��)z���ɟ��	I�ɟ��i�����)T��ҁg�V�����(�	��Şk�i��4�yr	]�e�:9q$��C�b	��\%�y⮓GrLD�ɑ��'v�i>-�I�3R 	jgꝧN� 2�S�^�b���p�	�P�'�|7݅/g>�$�O��3O�d<�!E����w�N��?��O���d���&�,2��J�]��`��9j��dj(?�"�S;I��c�i�g�'A´���'�?	�T/,���Ƿa�&]J%V�?����?	��?��I�O����X�h`򂎎��\@�e�Oftm��I\ܕ'�b�4�|%;3�.f��E���2�::"�Oj��x��mZ�'��ul�O~rL�L		���q�ViX�B@���yG�Hnm"D�|W��͟ �	۟��I�l�@�4,U2L�3#O�w��0� �WyҠe�b�����O��$�O4�������>�<�� N&A�ؕ�4��*\�ʓ�?a�h����O1�F^�~�*�84'?%�5�s�N)"��1�OL�� �?IB6�d�<s�PI@�pp�Z�y�������?����?q���?ͧ���ň��؟dZ��qn�Y7.�*�¸s��柌��[����զ�a޴I�����'LN=��h_�
�ҕp�B�=1�y�u�iL��.
-�@S�Oq���N�:�F�sE��t=�V���<m�D�O��D�O��D�O�'���~K
9�(�\��X�%}���I��	 �M�G�|Z��?AL>!)�t���,��X�U 8F��'�z7�����o;�lo~(R�3.v��f�LfO�|rRg��~B�6��)h���`��'t��͟�]NR��?A�Rp��mU������˥,]���%�H���?��B�@z�����ɔ����<]�Z�ZѬ�g�l��O�1�b�	ǟt����d��ğ�Jٴ\1&$	(���$˩d���'M� @�h�&�{u��t�]")��(ԓ�(��EW����B�'zU�gi�e�ێdɎR�#�1�?q��?���?i4GŧDǌ5X��?��2����j�)"����&�@S!R�T���O���3���զ���	^���I�!��[�O=���"���Bk�˟�Jߴ
�� ߴ�y�'��9��Ǡ:M ��O ����ܼ?Θ����i�"O���%!W%=,�A+x���B"O����a�#Czhk�����%xR���l�t!��h�MQw*]�1��q�@c�)W#*�+7��c��Ÿ��� ���d���h03@AT�2l��#�m�x��q�@	4 l���0�N�)����8�s�BS�.T�\�0o�l��Zt�C�2�㕮X�"�p�[�6r�C�-%�5�v��)�2��%-�#lC�T��CK�'B�ҍˢdY�",v�`dB�0��	�4�߽:f�����Q|^d��I�-^�m#g^�6&U �fG�PF�P�0j�qIB��ee����u�%e��N��ץ����ގ�J��	��&P�'�Fn��) l[�Nz�\j�ΉJ��ɀ�}��I2D�8��^�qO\����چ5٦�{5D��B5ʍ�R��[��U�)�S�,-D���p��*�D]S3B.
p��iFA+D��$��\M�9ѐ&Ւz��hQ�*D�DĬ�1IǞp஖�9�yQ�-3D�X�������X�!n�3%�8Z�
-D��Q��D�	w�H�K��� "%?D���V�H+DA�`��M�l��.>D��*� _/i�E��&H�5o�(��<D����k9[�i�c�ӹ55&<���?D�����&d�:�*�HR��-!r�!D����,B�HHY�M?9�έ[BJ:T���D��P��h���^02���PU"O"��@I�|f,���܊330@"O���'!,~�Z�dG�[2$p1"O %c�bY�[��$����/>�:!�b"O�ѱd�0i���uR�c��t`@"O���
S5�2d��m���c�"Of�)�,�/|x��`ކQ���p"O���s���d�xdE^.w����"O~Y�c$C�EPj���@E�>`(pB�"O��#F��>��}�7 ^S^���u"O���ۃ}�	hQ�߉g��I�'���q��EV^,��L
3�
��'YƘ��	�f�J�C���3��99�'���ao�5K��j5��1��};
�'� $��c�m� ʁHȗx��\�	�'bB�8��=�����4:G��	��� ��h��HN.��#�<Zd��5"O�x��%��2�Y���4_WT��w"Oh0�!U�H>��gGD�ei��H`"O|�A�lS1'�"�
�H-ޑ�"O���*�vq��Q���:�x�f"O��(��8J�q�$��@(�x@�"OTԋ��Y$O�\T?~�x4`c"Oȋ���F�a��k߶y��3�"O�٨7As����
�F�*Ò"O�E�¢�:P��;JI+*�n�Ђ"OX\Xo� c*lT	C� v T�X"O��DN�E"RX�@mZ=.���2"Ob<a�υ� z�1Į�8�:�'"O:M�@,�J�ӂ���̠��"O�Xi�F��B�l!6�E�1���e"OZ5�2� v�8�B#2z����"O�[�
�Ky.���C�5*�,R�"O���!a��Z�u��	6B"ObEzClʩf�T8RLJ�$]�5"O8�z�F� j���re-͉4�ƥ0"O���k�M؂x�5�K�Z��!�"O�dA�MEL[�M�"���zz���"O�x7�߭ �ƱY�i��9`��`"ORx*p�BLl��
��k���b4"O�mbw�5�>d[���9�N�Y&"O�$���^�l#K��8�i�Q"O����G�e�Iа���u�Z �"O4x���[��ؠ��L��,a´"OΙ��Id�P���;O)`=�"O�=�f��R����	O�V�
��"O�]j�G֊<�X��-"����"O"����0|(@ F\"䠀%"OI�ѥ�8\p9!vcܦJ6��s�"O�)�K�%J�RL�B�,nX��"O��â����'O�Jx8f"D���`�3��H�G*̫q�(���>D�����G"[S�q�`$ʾ,E@q2B;D��c� n�
�C#��31���P�D8D���#M���܋�B�U����N!D��a�)f�����L5Z�e��!D�|��.B%<��S�ꈬx�0���=D��Se��#"�mCq�2�V�68D��2�(A	O{�|����;c����C)D�1���`X�ܙ�b��Hж�z!�4D�L�LF����3eE<i�ޝ��.D��!�A>F5��I�-W�{��)C+D��97��=	�N�(ᓛQ�D�҈6D��P��M�o�lBfH]�A��
�5D�haT�M�?�6��3`��7p ���3D��X	�"�f̣���:Y�څ;�n3D�h`ۼYqd��2(Ŭv�Z���TJ�<A���.
-��Y�H1$5Vy��l�O�<�'�q�^�AU�ޭDÀ��ML�<�MA�

t��&9�1���H�<��ꇧÈ� �*K%���#�
i�<Q��M3��*v��4{z1�Q�]f�<Q�m�t�� 5�����P� �^Y�<�wJ�2hX�"�Tk�d%�T-^V�<����J4�A�7��3aD�ٺ$�y�<9���`�ly1���� �
��u�<C��qt�SuU> d�X�PLk�<���9M���[�|�P�Q��_q�<��	�rÌ1��6z���Q��EU�<IǦێ^�&�X6!�-���p��O�<� T�JB'X�+^��dQ�,I�@r�"O.MA�L�E�0h�� IH8Ĵi"O> ;�k�<7s �S�E
�C$- �"O�ёG�>{��a�v�Ȋ�*ܛ0"O��ڰ�8w��qa��[6CےA�w"O�]p�"[�_Yl�2�bH
^��"O��1�ϨGR$��@�E�)�����"O���"�txF�Q+ݍx���"O�ԛ��^_�jƇ��J00r@"O` !�:obzyr� е+D)��"O��#�-A+dA���nF
W�-��"O���W���qF����mh| �"O��x%OQ,;��m�AI�P�j�"OLI���}P1B��\�2E��)"O�e#����vp ���� V)�es"O�$��%�%v���Iط}z�X�"O\�i1g��&l�����^�@ȁ"Ox�B���b��Q[�w�b5:�*O��(�@&�j`J�rKx��'z9�G
�*���yg(�;�9��'��mIc˚ |�\�f���5�؊�'���P��L.��G�<����ȓh>��J�фG� ,�7-<�<�ȓC�Z�@���'?� �q־T��ȓ}U8AW�4�J}�2�S7$�2d�ȓx	���_��D�����H��؅ȓ\wvQ���ϰ�6(��'<[�N,�ȓI� S�����9@d���ɇ�^�,�3/�;B�,�Ӥh 
sHR�ȓL�� H���4f`X07ꑃlA^��ȓvn���� �gȄ�f�ת���D$����L�_�`)�B�t��%�ȓ9O�����ߠi�����Z�K�Ĭ��~�nժ�Ő�DY2��ğ1w��ȓv��Ps�!�ɺ�/	!�|��E��j%�΋{�j�``��G@Q�?�@3,O�pr���U(C~�ҽ�On�+�B�'
��'�	�R�%1�d��B�tB��+Ho���h���ܨ�G<3����$�$���<��BOf
ze���q!�X�<i6dW�L�̐�MO,K���i��TL�I)j��?�}����^�<]c���bDnA�҉�F�<AQ��3Q2$aH"��$.��g�[�A�|�q���2W ��v���x�"_7C����Ɠ 2� [��ͬaP���ώ�b�Tma$��e����ܪ-���sA�F�e�4�EN3Ű<��ν�J&�(:��2t+�M@HL:m��-D��{c��5_��pc�v�����7�x,�4A�{����C�z����Ls��Z4)Ö�y"�-��d9�K+f��X"l4��' 	�9OVQ��̘*h<l�x�ҀzBO�0�F䓦/����BC�$~���4G��h��C���0�Aǎs������9h-8U�剾}'
��=�ͪ>F����K�*n� Ӕ�j�<)�'�����&�;p����Q�I� j0�}��D�]����Z�p�2��fdɍ�yR��l亡I�#c���P����'��U03�3O��s�̈́^�5(��H���rO�q�O��`�2�~�����a�2�pu��~��8HFM�`�ej��\�b������>PqO>��qK��А%
��8;%���y��"c����S��Д�й�yү�v&!�s��97IB���C1�y�,Ҡ}�P���ɩ6K���OL��y
� <���V������4��KC"OB�bاjiX�pA��cP�� �"O �2%B�5r��1���AG�g"O�eiv@�6�ptr��ܼ55l%��"O�!��/�$l�� ړ$Zu�"O,�Br��9gL7��-hv[�"O� `͙�I��5gX�nHJ�!�"OZ�i�   �l �eO�%���"O���DGۂn:2���$H�V	��"O���o���D�n�"O�,a�[=p՜�����"H��"OR�� �Ɏ�J�(v��cҤ��u"O��� ���H�i�����"Ot��V�s!�MbvkU��Xб"OV|� ��!O��e��D�/_Ў<y6"O*%���Tff��W$;�J9$"Ol)ҕ@C)WM(1QS"	�+��{""O���T��$$ \��?�<��q"O|�36/�w�T���*s��R4"O�
�DV����1��ܘ!��)�"O* @A��-N�&���@�4AiR�3�"O.�
/����oB�b7�4Ya"OD1� ,�&OXi+�O��d̰و%"O�5���#+�r�;�Q�t�<�3�"O6H�及,Y#Bݲf����+#"O6�[�%�7Z
$#��
=;�i��"O��x�`�8@֐�1�M�/����"O�uj�/�SGl��e��>fp"O�]R��"fCꙑ�dݫz�:��4"OIHB�ޝ7v~���T{211�"OJ�{#��=����Ꮽ/�H��"O��8f��p0ѣOC�*���Y"ObtH�-V��y��ْ>�:��A"O0l�Î
 ǌ�:TÂ\��X�"O�����
��
_)tX�Cϛ��yr�3�%�6㟎W�8TSoV��y��O(c|�[a)S<xk`����6�yb�
-?��!5��s��u*a-G��y2f� bQ��G�L�p?��p��!�yb�	�@��i�P5p.�H��,��y��R<}(����7n�(��+���y�.N�=<e�wC�z�n!��ق�y��5�0i�@�qז4��!�y��V5jf$!5�S�\.�PgW+�y"`\�o@X	!�Y���!���]��yJ�>��MhT�Չ0��u*��<�y��\!����4.��)�� ��ϛ�y"@I�W��q�bַ�^������y��Ж	�f����R ӄ�L��yr�K%���@B�l�T��G<�yr��<< |���b ��.H��O�y����푅K%f8���eլ�yO��n��(b��>uU��c2�M&�ybeD ;h���� 8mJ��$&��y����V;�lC#KZ!d.��3���y������!	�0,-��Ϟ�yBH͌=bT�)�F"���v��(�y�Lنi�uB���/W�m!����y���X���#$G*f��`V�y��3=�}h���(�jZ��4�y$�*�v��B�I5�VL���@��yR��"a�x������)���1-���y2M�
N� `�o�+*r����J��yGQ�G<Z�J��Z8��0���y
� ����O!o��ia*̜0��]�"OJ��A⒞Yx��B	ʿf�<�"OT,�卐.6��=���Qhd�3�"O�J7O� _�\z��ƭSMV-9 "O��b 1 �z��'c�r�J�"O�X�ǫ�|��MRv�],	�\,i0"O�	�׉%�Vx�7���">lġ"O�a�dF1CP<� !��"~���"O"��F�"�.d��۵f���0"OHd�w� |G����Ȝ�^��,*"OB�A�C_��\-١�Fo�^l��"O4���046bU�7�C�%چ��Q"O(Y�q�H �д`#GL�r�F�V"ON ჈H�h�6H]�.�Z��"O�D��d��>ˤ�ё;�&�q�"ON̨3"�5BP�av썥�\��"O
�Ђ��s�i�Z0y��h�4"O�0�ШyQf��#t���"O*}2��K�i��()�
�^Ҕ��"O$�ʄ
h�����ϲ4Il[�"O� �C�>,]bt
�#Z0ٰ"O��k��$5����k��a6���"Oة�����c�Ԕ�𫕺&=ʵ�""OT,�Q��0���n6�щ�"O\��4�ȼHQ~)�@bҜc6()�"O�����D�*�BG>;
�+r"Oj`���v�x1i�ҰB$(�;`"O�1p����j8"5��87�e�"O~���Ži@������:/��a"OV{DO	W�b�F�8or�`�"ON�c˓N��ūs�F�
x��"O�Q3R��3n��č�x���"O��u �&n�����E�و1��"O
�#�L�D�R9�o�3���h�"O��C��I!Yl\���Ң!��\(�"O<w��o+Hy��R�
�^t
b"O8�Q0��+6칀\.�1�*O��*��X|�-�@F�;N�{�'p�eXd�Ҏs�!���1�� J
�'J������|���Ө<�V�	�'r�x�cG�X�� #���0�h���'jtA��P!�"	�Um�"��e��':���ញ$X����lU2���;	�',|��7�M�5b$8���'��-A���V�U�� �6kJ����'�eNN9YV�AEB���,��'�ֹ���|!���b-޲�i�'vص3%�hǤ���6h{�l��'m����숩 p��QŌ�3dF��	�'��� c�J�i����>`�f��
�''�R3AC�� i�@�+� ���'5� h�GHP��E�N�v�l��
�'��A�&eά"4�Q�9�D��
�'�V �$�
�V����/�&aP
�'E���K�t&�X�ҍ�>!v���'f���N�A�B9��'M�2�[�':�u�v��/r~������?HX���'v���		�A��4��[ NeJ1��'���p�܆Հ�)�i�G�0!j�'{\�I�O�<bߪ�ۇf�1G�!��'�8d��J��4>��W�8�R�'��<qG� jˀ�PE�L>Q5j\�
�'@�	�t !g� ���D�#af9�	�'�.e�S�Yhֺ���(��Q��H
��� (܀w���H�ք+8�`U�"O��3H��8HI���g��+r"O��p�SgC�EQ���}~����"Ot9� �݊!9@��ra��\$��a"O"�c�J1���P��3@tlJ�"O�	����0dj����20�Ձ"O��IR�Z<xB��o����c"O4�#D�0V(��㊤M�h���"OҨӂ�U]�F��b��b�~�(�"OdT��!�b�R���[��\@�"O��4Cbp�3'��2?{���ȓ���2�)ȩB�FX93(��-Hz���t����F�0m
��8e�@�n�6���h9����i����u�uS-r��ȓ2�8���Aĉ%r�h��8d��.@�ه��Z�ҁrQES�K�Ḋȓݰ�*�	N�O��0��0_�`��ȓ��u�w��'l9����* ���$�ȓE�=�@��>^��b�ɰ��`��OD}`�I�O��Q��%?�|�ȓj�-Ζ)�vɠ&
34�H��3��Ti���6=��b�`ės}�̅�Nk�����I���		Ɛv���I� 1)���+q��r�A���Ą�L�n��F�!+,��� P�Ȇ�q�Ȉ��CŀXƐ�g6+�̘�ȓDF��:�4g�U�1H�0,6�ɆȓK�4#��:VI��wCҮ7r���f$�]j��-�n�R$�R�d��͇ȓT\m��8~d��BT�H�0�ȓZ-�	�Bj�/C�X'+Ř`���ȓ��}�P�!Nr�J���6�v��ȓUl�����4^Ȣ���K܆�ɇȓ�m�ᮇ�<�6h�%�+Ha�|���6��j��Dٞ��7��d�4$��5:� aPV?@�a�C�
$O:�ȆȓD� %p�&X�6NZ�0C�;Q�Zp��4�fܫoܲd=��l�
m��U#�'�hd�!bN9Q1��<���',lD�p�U9p���qR��zȉ�'t�q���V�����P�{�z�9�'>�#%�R�5�xā��={�����'ي�bTD�c�=���r�\q�'�R�����-)�P�)�唝t,
���'����F�]80�6�s
��e><Q`�'Z�!��_(`i
���eA5]x���'�N���U�(G�P�B��[���

�'n��u�^8&8��eT�h���'� $�q�����o8f�X�'��X��Q8x�~[�.h�PQ��'"`Y�N��v;K��U�غ�B�j�<iq(0x�R��&�z7@���_l�<�g�����tꏀdօ�D�WP�<ipa�?z�z�*�댹�8XB�V�<Y�씘4ĭ"���5a�8
� ZU�<�'�H/Y����ώ.%�b���O�<A�D2�����OձQ��M��B�<�q̄�FMbq�w�\�����FG�<���(\��@�J���9U�ߖ%!�$ūf��@M�%g��B�c݇>�!�$���Uc��M5~6��R�e�3t�!�C�Mz�$���ͽ(�\�+���!�D�m2l�;ԆM;Ant��©�?!�X<<�d����֏kc�8ȕ�^+�!�� ��VFL!�؄i��L�}Yv��"O�\Cr
���ɂ�DYH�����"O�@�$������&C>#�0<��'�x�3t�_�5?�II��T�]Z ���'�A9�^7���Ջ��j`q�'ΘYS� _�(y�#���x�6@�'6�bt��9X�2(�L�i���
�'f�m��h�>��BC_�3j��;�'�l�;p�<Rj�Dx���C<���'g~@�T���s�$�:��<��89	�'������|z��V
a`�%8�'yPh��L,tmNɻB�L1�J���'� �h6�4���2)C�3�8!��'F�a9�ҟE�x�VJG��iI�',J�$傴L+q��J�,D8���'*N�n	��!�\!��C��0��'�i�J�-��}�^�O�0j�'�% W�V0W˦���
ǐM�p��'����%e:��d��Lpr���'����-/�@	���R�KU����'�� ��FS��i�R�D�q��'&c�!�)U&��g�/@̙֔�'�
%kԏ֦/a�Y��6���2�'��Aԧ$g}@�8�ߤ;F���'.X�� ȝKkf�3�C��$��'��(�蔤!���C� �#F@}k	�'�J��+I I��\µJ�7;�����'�Ω�0B-0t�����<�HU)�'���;㋕�¨��M\̩[§���yreߎc�P�k��L�<
�ؼ�ya/x�|9 �nޖ<�D�0��ǯ�yr�4�V͘�)�$?H`��y�]8$`.�8�fΠ_U��[��>�y�%�qh����0FHeivɞ�y2B+���խ�7���� _��y2aL�U"p�c���+Ln�ڣ��y2��D��(�[�*��M����y�k�G; 4�a(��(k<��C
,�y�%��~X��0��j����QJ�yR�@�`���3vc�j�:��I���yB�ؔ>[� �A牝Z>�������y�(P��@��CR�X�D@����y����J���s$� �X�ẻ��y��Vq�$��B�6u����dë�yr]�����OJ�W���/���y�	��r?p<e��%(���M��y��yK�@:g�Y���}�a%�-�yR�-$y �$����q�&
��y"��i�rh��j��A2y+���5�ymF9d��*Dr�vYs�#O�y�h��[��� �V'l�D�ٴ�ӑ�yc�oT�yXE��%j�,��D����y��@�_4Hp�L�c/0K�j�	�y�� �%`�jA[t>T�����y��� �F�bs�P7B����bgʗ�y�*�[)* �Kʆ�3gj�/�!�d݄Rh~��0w$�Y��Z�!�Ă >�cb�W6kl�X�P�Y�!�D�/�\	�R��-`�y:deC�P�!�$�*}�$��%� uu$��I5P�!�$S1jd>� w�Y��P�"�ڧ�!�d�"a� ӣ��7�2B���!��N!�#$ �t}��St���q�!��[?�>}��e��(zD����:cT!�� �c��A�k�dUp�I��A��A"OT�Kҗc+&�Õ�=-լ���"ODLـ`��0܄��g�H%nFlB"O.���ܓGH�0��pZ���"O�� �t�5sS��H����"OL�ٰ*F� ��Es����)�t�"OV��M
�a`6�)¬C�l��I""O0��a�m���J��?ݶ��""O�Z���Ű7����4�NZ{!�D׾#�=)��e>� ӊ�Dg!�ĝ	_f�����D��E��^�J�!�dT1<�-z�.@A'�ȶf�!�D��1�Z��Z� pK���3�!��`,����!,|ZfO?5�!�D�7���.tX���v&�)I�"O�ث��K�.�q!s�H�( �;�"Oū�h	8�5K�!P���q"Op,��̚�{
���Ə&x�Bqy%"O�h2B�5�E`B"���bi�"O¬�s��(�������{�"O*�s�P5D�����:m��4�q"O`!;�ʑ�h{��s�� 9�"O
���H!}I �wc�$F+!��
~��<f:����W�g�!���8D����#REYԂ�8�!�d�*!��|�J�Yg>2�S	dU!�D_�"�@�b�I4Y2Ĕ�"�L0!�D̗ �	���ۃ^�,�ۗ�҇i!�D��IzaF+K�e;��^�N!�d�iR��SdE�lhnqoA�pV!��4A�fH)E�4?^4���9_C!�DQ3x�:`�iE��˒��+a�!�Ā�zz��ü3[.��PV�ԊZn!��خ!���J�<5lD����>h!�$F$�21Q��$G���ڳlÏd!�$ �9K� � P2A���R6
�!�D�,T�T(���í���C�-	�N�!�ݹi.T�W�y�NP��l��.�!��B�x,(�KL)�hE�S�X4Q!��7f1�E����q'<�@�^*6R!�81$Z5�Ṗ0~�b Y#>L!�d<_x�˖,�9m�U��6F�!�$��)g�E�Q��<hj�A�� �!�$F2<���dH,��d��7-!!�D�_�m�P'Ӱp���aa��!�$JW�Q�s'�����%R�!򄉿~��`��F�2"�R ��!�ݒ42�T�@W����c��LM!�V�:$(`*]9&z@����:L!��G
>7(1r0�Ѩ����H7:<!�Ƽ��� 1�H8�bV��""!�䓁b(���'g��G���H��"!�G'
�<h��̇�ް����M�j�!��#j>� �B/ۃ}FYٖ�_�j�!��ɴ;X�G��<Ci��h%�^�6�!�3n(�b��ΨUJp IWG��Py"␽T��t*ŋ�$=*�&ߋ�y��H��L�ڤ�Ϥ^�(��T �yb˓+k�Ւw��'�n��N��y���u:���w��`Hb�R��y� @3�
\�CL�3Yv�〉̦�yRC�'D��A;����ـ`�L��y���#VZQ�is�p��W!�$�T1�T��oT`r���e��!�� Ȉ��㇈Q0Ҽ@�K�*
D�t��"O�X��*�&�d|����8)��kw"OJ��ϑk A�˘�=�9�"O^�u��3�RH��i�(9Mb�r"O|�y"1q����/W�?��"T"O�����}�n���58 61j�"OV5�I��k�*M`���.�kc"O���`��F�b%��.�:hp��
@"O�M�'	-"��+f��7CzF��7"O~�"��96�G�oj�%��"OH%��n�fM���(NP@�S"O�i��֓~�u�U�^�Oh�|� "Oz()da��-��X��Ң5`\��"O
��E �f���ц����"Ov�#��PPd��SJ��zS�"O�����X���1z�ƈ�zIB"O���$Ⱦ{v���v�Z�L�2"O>�Q���5�6�'��e��"O � �һb�t@�1�V\��"O������r�j����HR*��"O��i3HX�_����b��jE�isU"O�<��R�ʚA�`�!)�䙆"O�H������Z�����I�"O4	�P�� qč*#�I��ɢ�y҈��<H���$Tgn�!�M6�yN;DCҠ�R�W�A���)1I4�y�
�e$�	���7��L� Hͤ�y�d˫~2�i6��,)�`� )��y���Y�:%�2��P�`�PG��y��ٜfP3�ܹIp�㖌U>�y�_�*�"���B��"N߰\�`P��Y_�(r��Ƚ^_h�MO�"1�ȓe��[���Q}^D3����Q��ȓs�bܑ#MKed<��V�$`���[��`�v풓S�н"+Êc~@4�ȓ?���w�O>5R b�
.��ȓdf0� ��#���W	+���4�������g��"�"�\ �ȓ]�����!�?V���˃k�.��������k�	;�%Q�AS�Sb܄ȓZ\�ɸ��[�l$�MH�B!:�R��ȓCSإZ�!�~xݳ�B6T���ȓ_�1'��009IR_�2��Ʌȓc�����O����w:-��x��p�H5p���V���`	�Q@��e E�V`#|Qa�K��ȓLIF�#R�[
m�0�@����݇�@�PK�������
uG��q�"��ȓk?�Y��-ź�>)�s�F�[PZ���m��4��
�5k�,�a�L�[���C�"�y�W�R�y��N�d��<��BN�%�'m L�f$*4��%e��ل�k�4\CWa�7�A��%O$.M4y��RW�XxS煵c�I�!gK!H�T�ȓM)�\�CL�N}�4��Xr`��	�"�7.J	.<H�GY�U�8���&�}+����bQ�IC� ہ\�H���jO�seܲ�XE�vi�8�^1�ȓ1j�Z���x7h����1������� �@�H	*#�	�2
D(j����p�� !�*HKn(s�J=W2�<�ȓ=��H���H�dph95��?J+
y��d� 4�S�7߈Aɗ�;�z��ȓ%�T
����lP��V�j�����S�?  :!�E�<x���*�3��Y"�"Ot��"�������c�'
] �2�"O�@�O�8<xUC��;T��F"O�)x�N
`�a���8͑�"O�ѓ3�>I*��[��5��< !"O�ݫ����eބ\kE��/,HA[�"O���OV�s; 5�FI���\�"Od�QA
�e��gF(9r$"O���Jۮ/�(Pr�'_�mB ��"O|MpDE�l��f�!N�#"O�i���W�kr�Y����>��I[%"Or%Z�,2cx��W�Dzeᘍ�y�@�:l3�d�U�F� �"��T�]��y"��"� EHĉ�8v[U��䝳�y�ʈ*��J�I?l�2��bQ����hO���<�ňٯ����I�2W��q
�@�<	"%�:#Z�ԲD�ê,W
`*c�<	!ܦ?�6 ˶�L*PL0LCԈK�<�a�-�6��6��Sþ�`��p�<	nR�<��9�E��v&�P֤_o�<A�� ;�JA:��.-���Gk�<yf�!����-dN֬)��e�<�4�x� �B�U�~��E�Id�<��Ā�g#R	4 ��h��y!lZJ�<ɶR�7{HT1�J�o88���D�<�&E�b�\<y��PH��D���<�䄝�d��=��ɋ�v�� �#O}�<Y�D��d(�YU��1���p�KFA�<�2gΜ(X�@���-)�!r��F�<��R�0��@�#�'W
yX��VB�<!`
;^�x�� V��Ś��e�<���0i��gʃi��Ē�*�l�<�e��WtݑCL�d:Fb�e�<)fj�,A.5��mF�W��t��b�<a�ɥ[811��=�"<+���^�<�5� &�\kQ@H�A(Nqp�D�<q^zH�bv#̵U���ó�F�2B��"K��1�f�9rc�$Tč�VOTC�?����/Z������%���Yh<y�ՐnP�up"�^�gDu����\�<�G%HC�l���N�a�F�@���^�<I� ��1=��q�鏇_'Np����Z�<��Ӊ{�fC���w��y�f�\�<i@�@"b8����ʆP-nU�cE[�<)���w�@a��*�7�N̉�.�T�<�".�9�pU���{��Q�͎U�<qv�^�@�h]As�.�l�h�L�<��"%&C�eL�V��h1�I$D��1w쐏`t�-��A];)�8�Ej%D��"W��Vmr(� D�&*�̑�o#D���`�ϴMF���$U?zθG�?D�4�1�8e(��[@AD{�8���;D�Hz5(H�)=���B��*v(3�,/D������	9Rs��O�{TH�Ņ!D�,�E�BH���/Μ=T�*"D�(`2 ����)Fi�q����M*D��!�m��6�j�G
�
C ]xV(�O.�C��zC"�l���K��	EQ~e�ȓ]���JR��?>R ��Im �ȓ0�)9�jϡ%�2	� ՅFܔ�������ö1��yҔ
X>S�����s��D���ŧV�,�KE��^��}��-��DaōN}*�KЬ�i���ȓrU��3�M�p+��#�I�tm䀆�S�? ��
�!$�n�
���1C`0Qw"O�(����9�>ѫP���[a��(v"Or���.}��tZ!J<ZHr���"O�S�J������$�?#\�H�"O�����p3�4`��v'n��c"O�Up$LF4��<h �_�;3����"On��c���	�`�A���i+�d�'>b��;\� �!��{�a�D�O�h�p��ȓ2�2�����,�n`���=a����{k����!��Dm�%��Y�Av݇ȓ.��Q�v.��Js��Bƒ���ȓfe�,�`ΘB_ XZdd��ˢ���1��m����3 �0r�66�� �ȓ=��!�D�<� ЂAU�T;$���П�'��D��'d����+��q,a+��=�$���'F���n�+�*1qF�e3�I��'�c�Y�$61�D�LX ����']���T�_��*�E���y2�]F��ȓ��A�@AD`���yR��
3�f��1���$�lt��jS��y�CK/_�@�ʃW'0������G)�yB���R�Խ��-P%&��e�2ꈼ�y��)G��|(&៫%=��3�Q��y�!ħ#�BL:G��I�Ԥ�Ƙ7�y�˛�h��C.I<<9��
�
�y"�,m�fYId$�l�X�C�ݓ�y��O�f���)%j��Q��J�y�C&g2�y`��<75� I����y«�D��pS��!L̍��+��yÓ=Ҧ�CB� .� �ή�y��7P����ՆpR t�GG��y"��	�]�������OP2�y�!�h1��ţ��p���ǋ�5�yN��[� CG��sz5	��y���6�V����@('��91�]�y�$$�j�;1+r�ub5��<�y�b
��5z�&Jm99��\��y©æZ�J�[�Z�d�\y1��ُ�y⧓�N��9��e��I���qD()�y�'ҹz�V�z#k�42V��9%Ɛ�yb�7�؍���5\\XQĢL��y�.��/*@hJ�l�9M�
��yR`��5t��I�3=�t���U�y�O�d��z�I�ľ};f�\2�y���7EI�����M�P*�yb`܆]`�BjW�Ύě"�J��y"�� 7���a� �5���9�y2/���q�T��<Y/.-VDɜ�yb�׫�J�̭Se�R婕#�y�E�<y&2	� 'U�L�X����yB���_��Ys�G��Qc���y2b]�g�T�K���9�)顯٥�yr����AQC��CXVa�A���y"a���XܓD�?��2��yb��S�8���ܷ'�rT����y�*ِa���qh��"��4�vk@)�y�LN7����DW�(6�*�y�چzt[7��:9�Y!&`� �y�,_(z���9��
.�p�P����y�M\�u��{Ƣ�)�����y"ņ���Ԓ�iŐkO�=���L��yBi��|�h�%%^�e������]�y2��wH9K�c_ /��1j���y2��|`�pR�71P��� ����y
� ��;���X���&K΋@��p�"O��)QO�t	�yz�iG>|�LqR"Ob���ɞ(o�ұ��(�$�j "OF��f���t$��Ǔ�F�:�I2"O2�K�f�WR����R�&���!�"O��:Aā�!v�3d�	E�.Ԩ#�'I��'��
���7f�B�1�I��`H�'nH��@^�t��5T
�53��a��'�v��5:H���ş(l4�!�'�8Az��Ț)^�5�2m��T-��s�'�ʝ0%*�}�6����/@O0���'\���c�q�S�M��4�L��'�^�Ɖ�-6= T	��1������?Y
�D�|Ys�Z�W@��q�n^�H���A,�pC#�J?*d�hG�O���ȓl��Bv�4�>�����~@����ް�RQ�P6l��'J�??���ȓ|L��x�&��<�9� �ɀv�x��ȓ:�(`2��ʦ	�.a9�e�>��ȓq�p���)��V��h��޾NIH��ȓĒ0 ��T�B� a�5ϲn���!��}iqiŰm�J�KP�E.��Q��,�p��gV�
�D��2O��;�4��-�:���C���������^��ȓad�X���_�v�kP�`x*��ȓJ$6u���\�$�nHo\���L��'H��q�.#A 2���|�N ��'{�<b��8��y�Wg�80�B�	?+�$�h�#�� ��a
±��C�I�}��I�d�R/bW�������DC�I�0:\35�!rx���
ܾ,i@C��.�q�AaH4�,"ai�1�^B�ɯs`�	(�I�s� ���Nػ~.rB�	�j��@���͐��t�󇙵q�|B�I+MX CG���,Hr!�p�U>B�I-��r+��P/�x4	�:��B�	-+8��𢎐D����>)P�B�I��!��%|r�
��B�f�RC�6`��hS`	�$U�� ӪG=�C�Y�h����
�u�bD;p�ۃa�&B�=yf�@rrƞ�gBjLc����JC�0l�a�&9?NdJUI�/) �C�	�A��X��FI�
r��xR��M�C����س�(E_3l���ܱr��C䉂 �X��7/P��� A��C�I4Q���fe�y�&���C�Z�C�	�Y1RA�7c�+pMX�w�ܗA�@C䉰F��EY`@��4Y��nЩ[��C�I�3֧?̶=p�
OxX�C�	�.�h;E�z���H�ΰ��C�	-yj�(GΓa�\s�96ؠC�I0&� X��  ��K���w��B�I�d��BF�ȸV�0�M5(	�B䉵!��i��K؃ ��Ti�h�c֦B��1[��d���&Ln<[t�Z��B���zi����p��e�'%�d3VB�I��NQ�cW�-g�-q%ġ+��B�I9kŒe!
1*¥YQ��N]�C�	�0�Vq�"�Z���\ ��3=v�C�I�B�,�*!��$��K�W�B�I�&(�4[��G"��଀8n�ȒO��=�}���2��ǌH�f��0��HV�<!��M�O5�<P��)�4�ub�O�<���1;x^P��f$�<�!`��K�<� X���a�4e���vG�,gČ�"OJ9����w��<��GM�\6V�i�"O>����R���i��ۮ|I1�g"O�%���$�:��6�̋;4���_��G{����Z����iF �����f�!�$ܦ@�v=Bum1>ɮ4hݽ<!��� Hz= ��V�TP�!��*�!�N6z�}�iG�^���u�O/)!�d]"O�I�Ѩ�s� ��/ԋ!���SX� �F/
���U�!��Y� hip'�����H ��'�ў�>�3�E�"$
���-Xd���5�?D�\'MS� ��'K�G���G�2D��S!/t�1" �n���E�;D�TR��?U"�y��^�#M$�I�N4D�����P�V�X�o�I��kq�$D� ����4G<i��J�
XSZ����,D�l8�AY�d=pay���5i������*D�H���ܒP倩�"i	��P��N=D� a!�/2d<�Y�ܼl���J�6D�D����%@���+�hL���(D�t"� H�L��&ưW�Z��w%D�(ð�:w��y��O}>!�#"D�X�H,v�"�2o��5e��6�-D���ħD./߮�B6�Q�&�ٷH,D���1"ޑn|�+ Đk��[�+-|O$�D2?�b�"8�|7$�Kεч
O�<a��=h��*�MռZ&^�!�$�M�<a�F��x{�h"c�:E!�g�D�<�E(?��i��H m���a4bY�<)��,Ly���
}
�d��T�<٣'�b�P�r�BYKF�"��_Q�<q��I��J�jZ�7Ϣ�"�I�O�')�Od�)��\�\�@|S��E�0����ȓr�j��/��G���jU�&x� �ȓb
�����[i���Bv'N�Q5,��<?>� �4p	�Թ�'�t�5��u��=@��ڦk2x% R�V�8)����`2�A���EvX�cU���\��v\t���HfN���M"AZ�'���Id��DUg����]�w�U=��a�5D���E��cYB�Q�+�M]�Iq+2D����)y85b��ԔW�֤��5D�H��EB�W78URD�l�b����4D�@;�,ԝfblQ˱� c,@�rA8D��*��V<��K#�ޘO�n�0 �<����
fT���ա�R�ҙ�Cغ[�<�=)Óa!8E�i�/� {�#��D��w��A`)b�"c��R����ȓ2�Xly��#�r��������y�BT�1I^�G�,��1�ֽː��ȓ{U@�W�EZ$u��F�h��!A�����R�;��4M.�F{���<��3XG�tq`��0{���3�^�<كG�i	Tݒ��U�:@m(�CW�<�G/����a��,ew�H&l�O�<A��įo��Z�����ț�A�<A�xK�@��C:�P�3��r�<q#BY�1�C7�ۄl3��"Gl�<������t<��O�>\�q�l쟠G{��ɞ	~�h����B\���E�F���C䉟I{^%���T�*����oD�k����0?�p`��itT��m
.fQ��h�<`"\+~�p�) o§LYJ�g�<� PM#��5�؀!�O���8G"O|��*	i����%%B��Xg"O�9�ת�C�pը�*�+><br"O�˓�ǅ4�F 3��yq��{'"O�|(��
0z�<D���Ӕ']l���"Or
�+���z��ǋ��W�<�""O����	�\jD%_�@D�p"OHrt.\2_J|�ˑ�py��4"O�Hyq�Z�*<���#��L~�#g"O& ���	Z� Ѩ$h -�R"O�<[���P�FP����H��1��"O�yQtbA�C��`���=[�Z2"Oe!îӊy20����̱<PBRS"O��+�ur\�ZCMK�a�U[�"O2���Ef�٢�J�`qQt"O�X��
-=d�%zw*�)&�xQ1�"O<ا&B�VP�Ǣޕ#�:�{p"O� �b-�<�$�r����:%"OdE��BV3Kh�h��a	������"OĀK4(U��@��&E�W��x��"O�y�Q��/kUD�	��G�#�4��"Ov�eFj�<���ގK�$| b"O�E�b�X�i�:r�i�{P��"O�9���R,WVl b�B]4^a��Ie"O\,rGQ�(�f�xᄖ8]�a"O�f�1J� ���Bi�F铷#�<��nnD0&NО,�DЧJ���|Ş<ó������a�-��ԅ�'}t!@�)�����gP){H}��V)��S��5P�+u�6 �`�ȓ�؉�g��zT`S""T)F�(��p�B���H�6
��*�bG)M]ƹ�ȓPSd
e�1^|��NĥVN �����!g��.�D�9D����8p�ȓw����M�"z�h`�P�]�!���NI�lSqA�8��If�в4!�D�����[�I6AVV��E�ӳ�!��1Z�*e��g���1�9�!��qÜ�ۢ!/�\����Y!�d�A�L�R@/Q�.%��	�m�!��V��:�"��w�lв��;�!���r�����ϴ�,�c��Z,�!�d!⺰;�L ���T	�M�!�DN*؜H�e�6>�@ȚVl��]I!�$G.$(@)v��79�Jy�#�BPQ�2�)�dk�B���#��W9O���C"B]!�y2����ɐ�Ј���Xt��{Ј��SH�UT��cf�愇ȓN�������M�X�d��0��D��P�H�Q2�	�u)���g�����8h>�aCM �p��ӡ[�$4��u.A����tw��(���7��?ɉ��~�ч�Kq,��$��4Ct�jՁ�D�< ��=:@i��+�0b���g�<� �]��2l"��_��P��u�g�<y�b܄K �P'�?O�1���b�<��"G�7]:i��:r|��J��QT�<	ã�9��T§B��Rx�����V�<I$/� v5�X�^�1��y��NQV�����n~�  Ӝ!V��'`��,�q͛��y����Tb@$���Đh��� ����y�bŨN���LȨ[�n0I��M�yb��VN ����҈E:�y�m���������"m�t�٥�y
� bȻ5!O��hԋ�g��E��|�F"ON�K��K�2�yr�Ha=08�e�F�����J~"��FҢp@�M�>�L� 
���yʛ ��1�°I��b��y��m�@-��.M6Hlԡ7Ő�y���t�ƀR�%�%=\�ؑ�W��yb�%�-R��Ҕ4Ѿ!�ai�=�y�AY;vI��S�cW���1���y¦�7	���#c�(<@`�/�y�͇^���
"���_��p�gL��yr(y�F��0h(�� @�б�y�����0�+Q����n��yRJ��yf�`�����H�� )6"ƺ�y��kۆ�Rq�į>(�pJE"��y�!�*K�l��./��tp�ŧ�y2DL s���Q(�<��݃����y��D�Wm�QI��`��M0@�N��yRM��;�(�3%_�S<�����I?�y©�.$��B��M>�:A�1�y"m@�n^D��K?3����k��yr�R M���Af@	�U��X�Cͅ��y2.ӊuΈ0D�I�EF&	肤α�y"��/I�t���U�1��ZK�+�yr��$�Dm�)"�� Ӧ�؊?!�D%�e�� ��5z�P$ 
w�!��:WC��95a����b����!���EPh��Ӫ?�l �BH_+b�!�$_��4�Ⲋ�1��|�'ȣ)v!�d�)%��ջ�(�z��"��#Ov!���
��R�Ԇv� ��C�X�^S!�$C"h�x��ԦD�2�(�2��� !��J�q�th�F$�c�<�4
M�L!�Dҟ~AZm�L��
"V0��ȟ5b !�d��h�e����)Q�hH�ö7�!�ĕU˄䒤�ΦJ'|����In!��]�Io�X J�V�j�F1g!��U-D���
�9A&�+EPȹ�"O���C�Z a0��A��#|;�.���"�O�5���Шj�z���DW�Z�J�s"OL�r�Ӌ5�Ή�2Õ#}���@a"O蹲兙�ok:�R%dH,IX՛�"OV\�i��8[x���m˫26��J�"O|r�h^.PM���K��e��E1�"O�T���!�|����͢#ll �`"O�X�!�� ���K'�@�4�X�i�"OJ��L� _�6�����3j9��)""O6��Ũ�.m�R\x�kG�*�0"O�d�G�����C"%N�cr"O´*2j��IQ��Ӗ*g*�J�"O�S뛈.% *Sp`s�"O�)궉�m�l�T��+YN��{�"O�#��P�H�H%
7H^5��Y0"O>i�F@�b�����@�*r=`p"O���q�X�Ty��R̶6�8���"OZ�hƤ����Ƀ+��yZy�w"O
����["�C�ަ.u"��"O���e%`�I#�F�q�#d"O������v��QVF! Y��[W"O<D��R���B%��<Gj4��"O�
g�v���qoG�4aH���"O�M�u�G_W�\��+I�Z�d\��"O��4o�;R�e�jJ��(�"OB43�b^&�X�
�fF�j�±b�"O�Y(ՊW�j�Hb���R�~�2a"O� ��c�ď�(��W�LĀ�"O�lk$�^T4`B]���l`�"O0��ހL:B �V�e~�k�"O�x
���^F���5�ާ>� 9Ar"OX���R�B��"U�@�X#hiH "O���q�_�5u���gcWs� x�"O��x"��X�9p�":R���""OF�9g�'�@kUŢE�\rgO�m
�U�q����N[�� �	9�!�$8��(c%1x!���i��u�!�D�c�L9C�Lb~�XXqIA)2!�D�U���gE�.Ey�,`r��-C!�Ę�v沘�l��?b��i6j�$.�!�$�$�fxR$�V+-�<��0��/U�!�D�5T���*���	���L����
=,�^����.Z�H�9��E�lE~C��2 	(����7�PP�PJ�7�hC�I��R�Y&-TWhѱ�O �O8C�IN��93�ߎe�6db]g'"C�IΠ|����a&,��Hk�B��81��}"`�K�b��l�g
"
A C�I�sIPhʠl����v�4B�Ƀ\��DБ�F*�Rl�'(D	Q�B�9g��=��T#VU:��%�C䉟s����� 6+P��^Q���	�'�Da�t
Ÿ8~�t�%M��Gv�`
�'&0����+(P4��Q&T�P�'��Q�Dj�-%���J��ũ#f�T��'���@�bQ*l��-֓RA
���'��A�TNJ14 ����@V��-
�'ӆ�餦L�wL��Q��*Lk�U�	�'��u�W�S�:�Kq���IuT �'��(��tf�BKΞ<5f�(�'LȅHDE�.L������7]��B�'�����E�h�p2�1$"�	�'È塑���� �v�$\+�'3�C&(ď ͠�8��B�!$X��'a^43����u�����W ���p�'n���!���M��oT?��'k8�2�� ���X�+� �ɩ�'��|�ѫ�%�dH���	<aJ�y�'3��p������!v�@�D"���'���u��>A�}R�#�%�h�<i�_8���Aƌ�1nҒX�FLN^�<�b�JJpz��TI�91�)�X�<�%*�mR~�XW�B�x3r�(��NT�<1&���
<�v"$eĚ���n\M�<Y �T�<1��ag�["9�8b���E�<���� ���:jX���JI�<)ABnt&zp�� �%�o�<!�G��1"�L{��LS�N�tʐj�<a��5\�$h'D���Л�%c�<�u9�z��R��= ���y���[�<A���$'b����P�x>B`9�Yl�<����<c R@S��-B���@��I]�<����n��<���Z�=!����S@�<�p�σ ���1��+����\{�<�$f[�b��,A�#λ;�*��v$Ax~re���0>Y�K��`�����4�^,�P�Z�<�S���.x���ڂ�h� K
V�<a^ɠ� �-*�p`8�gUR�&=�ȓb0��ReKߊ5H��A �$��ȓX�d&b�%n���1��A��$��Vs��;CJ�}���e!6r��S�? DT����D�v�� Qv	($�|�'�֥Ǎ[<��;hR.���9�'��0dg��r�
�Bч�9d�x��'�r�&�ݒNr��b�L5E�q�'��ۡ �8x�F=!0�n�j	�'�v�C�\GW�H�ܳ��
�'�$�;����%�J�+��,��E�	�'�l�W ��	�ō
՘}�	�'�>A�ɏ$8��m�  )�|��'4 -���^�?�V9[�G�3��<��'��h��X'�`[1�_�G�N ��'��ih �Ą-����@ �@�����'�^m@Xh	G��)Sd1Ӄ��y��&>n��SgDF���eFP��y2�*e��&O��Be�X�����y�C�$2xa�"P(;���w"0�y��i�<e��<7�9��+��y¤O<b��$�3�؎?hcg�֦�yr�� �.1��Gl��h)��y YH{�D �-�J�t��yR��o�,=3Qj��4EV�j ��yrb��
�($(��Y�&���y� ���yb���xID3��E	Rm��y� 8] �Y����2�4���́!�y�i��X����)���
��yBA�z�T�*(8����F�Z:�y�Î�,�h��߭-n~�`�*	��y��>gv�2�������6�y�,jA����!H�hѭ�y2`A:!�jꆦJ9r pS�J�yb"�s�8�E�U9����RLH��yg�	�	KW	J88r���y�E�Dv�P#�}�.�x�bK��y�j�&4�fi�U��3y��r�m���y�Y��QRĎth<q
s���y"�؊ -�pk�,C�oe��QŮ+�y҇C8_|,paǭ�np�����y�M&D�0��DkB���R"�ybG�x�X���^�e�D(���y�*Y7*
���� {��B!���y2&חK�HL�֯h-l|�kQ��yB�04�Uɋ�c�@h�'ſ�y�g�7r���E+?Y����邬�y2��%]�-�Ɖ��x�D�S��y�	�=	�v�^�jp�
�S��yH���U�	&�<L�f���yB&�d���c�gB%y���y�̎O�b�����mJM�V+[��yr���M�*(h��H�8{ ����K4�y�L	#�����>-4�r���yrn��o~���N��y����f��yBȃ�H5 � �PrԨź���yr�ٹ!2Ȱ��_�e�B�v���y2�	<�6�C�@
�
��)+V�ė�y��(_�r��6d�����s`�N8�y��]A)x�*2ɐ��ǅ�y� ��+Ȃ���΂vl�d��'�y��G�3�uB��2_�����(�y#���aң��-;�t1��+�yr$�Z^}�G��P��\)P��y�mB�4���ؑ{N�P�C��y"GզW�X5�3�ìb�dLpN���y�H��@>��v��]d6�7�W�yB!��|V�u0%�\�9����y
� 6urH�p��8cg*ߘ�H�A"O����LѓM��a��3O��I�"Oh�kQNص/؈p4%�]>F�A@"O<qS'�ԭ%���:U�͂!=l� "O��)"��N�	��u�H�""Ox�YM�2U����W��2�a`"O��ȟtt (
S� ;�:yZ�"O���v��Y��1����u�L��7"O��Z�$|ԙ�o��~#�]+w"Oy*�(�2�L���c��~,��"O6�����.�ؑ���	���1�"Od�ِ�/w��)cb�J77�~��"O��(�A�(+�� BŮ��6tr�"O\u�u�Y)^�R� 3.ɮ~ָ
"ON���!B�b����wLX�=�M2D��� �A���B�V 4Z He##D�Pi��t2����g 6�R�/#D�l�5��8zR���AI-D^��"#D���5�3D���YwaF�`�B|`�&D�h�Dֽd�"	S���rB�� E�'D������&T�8�#��7p֬�6�!D�|Y�%�8��X�c�vqtY�1�$D��+�$�H�^`GX!L������?D�@R�gO�Ͱ�BJ6?��eQ��>D���ckk�Fׇ�pn�@CO��yR��v%�e�R��@��4J�o�yrIQ�j5��(�ȋ��8������y򅛨c$M�u��z�x� ���y��<y��F�V���f&%�y�Ϥ�I�(���!�!��y"����`ǧ �"��߀-?!�DV�MX|H�%A�9Ft��d,�=:/!�DO,
1�Y!�F�OG��23��"!�ǁ"��ኴP��KBbA!�D�'b{L}��X#`��ݢ�˙�Xa����b���J������Blߵ�y�������̴X��U�Ⱦ�y��L���,��%@37�3�I��y�%K8.ɑ��&-�P��埞�y2�(}q�C)�Q��X��y��T�6�D���eܙ"�(��FN��y�m�F �m��a^���%�Љ�y���Lڑ9�
��4.N$1����y��P? ������\�E�wN�y��.���[��ǲ���q��3�y�c�[P�E�Q��y���4���y�Xo.p��%F?�ࡹ�E 
�yҏW�}���Pd��l��%*�M@�y��D�=8�� �ߐ_?�PC�٣�y��ѐ}@���o�7n�"]3����y¨]�uj��Ύ�=mnihݵ�y��E�J���I��Y�:آ(��A��yRL�Q�Ӎ��>a� ����y2EԺ�,T�V�� {D #�_5�y�MI�A��R�kWL鱣���yB� (�Ĉ�닂3��}h�&�yoD	8$qB� L,��aa�� �y�bʂ:H$�+�c����ph��y"�>;����Pꅦb.�	G,�5�y"�Ix����6�M�q�F�N��yR$Y*����1�S�F
y:��/�y��9���qō&l�(=�%���y�aTt�+R��f�JXFcQ>�y�n\:_���2/�\wH-9tNÀ�y
� B�A����,��A���L�v4@pv"O0�8%4-$~̂��<<���"O����M�-߰�Y�7S:��"O���V�6CF��i�m�4�I�"O�����[5LƐ�Wcʔ@)I��"O��� �H!|��Tb���a��"Opq[5H�2c_��q����SΙQ"O�哧(��Q�|���@\�=PF\0v"Oj}I�
T�v��٣!fJ2-�AB"O��A�ה�n�C��U��`�"OPq�ʙ�L�)sd�(&{ U��"Od��0�,mJ��[�b�:���#�"O�uh��7F��S�/W<�r�X�"O �)����;���w�>�Tyic"O���E^? ��Y�.�g|z3�"OV%@A�T.!�����1~cN8��"O�)P����<�WO/V&��E"O`! �bP�2�iFC4ZC�{�"Ob�ÖfY�/�$p�@���>�`��"Or5x�K��t�=��K�BU��sT"O>���iK9�.yYa�������"O5�fK�\���T�T?>�V��%"O <��,Z!@�Dx���V=4��}��"O"A�Q�AzJE�� N�R�Ę��"Ox1��]�;�|�������4�� "O��I��g��x��ݰ_��=�"O����;]�AH�#ތ|5�"O�i����%\�̩C c� �
"O�H5I��
d$Ԉ�h�E�"O*�aa�^�����ao�?�l�"O��* S�X�p$��x�"O���a�J�$�.%�jL0�`)�0"O�!؂@1Z�`(�D��r���� "O�q����!��)�'�^���"O��3�P�H�r���HK����"O��
tʀ)Hh�b����4�d�z#"O���`?,�A�"��n;�9q�"O��Kf�9��Y�&�Hd��"O4@*3��@f�(8rf�9$<1�"Oʨ��"�A�fhɖO-:&(��"O�����/K]�qc���6�1��"O-2dܵd|�5�îF���A"O�Y�"����qbb�H��- #"O 4؂hL�s�µ{$���qt|�"O<���cOa'4��10T�ia�"O��у��|���g��t;9�"O�H��_ %�ph(�eL�&/����"O`PQ�]�+t,�H@�L11ɼ$C�"O�@��30��*a�EL��z0"O���e����hȉ�d�-����"O�`�K+ H ǄR+08����"O�u"���W��p���?5�MBb"O��z��8Id@��p�_�h����"O�dC�N�%k܎p�S&͡*d<���"On�˞�a2���o߬((�)�"Ox#s% }�� 	��N+e4�hr�"O(;��
#.R�Q
<N�`��"O*�"`��G~l�!�����P�"O��b��+�𸻴j_4�ؼ�"O@@�����L�+���84M��v"O�m�#ц[ʑ����&����T"O���Pa��`{�M�����('"O<<CR�Oto���bB�'����"O���I�F~�A�&� :'[����"O� >�C®w��h ��/,Cƌ# "O�k�f@�k9����F c$4!��"O(�I�C�I-b,S�O=$�H�"O�rD�a��U��q��i2"O^������L�9��'��� @"OZ�����mr���T�x��I�"O!�eL++��<���f�abr"O@!A��I�+���"^,�:QR"Ol�sEN8z(�ș�.��C"O��@�Z  ���z��8J�R�"O:}�5��59�`�ő�P5Q�"Oԉ9����Y,��D�*jp�	"O��X���=�(Myu�R�Z�6�yB"O`: �@���\D-�Q�*<�"O�T,�,Rp��߈K�v,h�"O��ӭ�0L��jʨF���V"O\A�RZ����,�&��lҔ"O��*H�:`��!G�~�J�bu"O�E�W�F�W���7�y�"O8=�"lݨ` ǭZ�^��8��"O�}�bfJ�y׺�HmG�h�t�؆"O�$Ja\�P̜�)qO�>����"O��[b��t~�Q�ɓ3k�����"Oȡ�nӃt��YU	ƪA}��*�"O��ǒ4�u�P�Ґ5�b�""O t�Vŀ4J������U} �Ҁ"O�a;�`U1T��q�BT(|��4"OnQ��N��Z��'�D�E]()�g"O��AW?!��/����	�'JZA��D��U�g�X�kL����'0� ��AIf���Jg�]��'��$���_6^t"0�b�O1gt��'���2AǕT�a�g̯2����'�>XZcZ�Z �J�	��i��'�ڑZ0֝q��4���F 00�D��'��x:U�~ՠ`G�QE�Y	�' ���cǾt}Ҡ�W�8����'x���_�A���r�H�d�j
�'��; `�?>����a�HWvL 
�'/�h�F�Y�5!n$kae�Dx�)�'jt���$�%e��Aa�Z98K2 z�'����+�DٷK�1m�1@�'"Z�ږ��$r���G��=,҄b�'���)�dtÃ�b�ذ���:D���C��5�U D�هM�h�7D���F�2Ű�� 7���H �3D��q&d�3m���b���IȐ��0D����d�$�@�#7e��(c\9٦�-D�L3�җ;�#�ɋ�>%�*D��b,>��I[g.�{d�`rpc5D�Py�˙s�fU��哢)k����@7D���2J��J���MB��i�m4D��C4��J �]ذ�(O�ܐ34�4D� �"�!T^��� ܠe%0D���pcH	2��m�$+�5׋.D�D�FK�2H�P����$]��F*D��ڦa�����׏3�xu��%D���p!N�^�L�A2-�p�d'(D��80�ܐs�tP3�@S�S`�4�%D������
��Qz aV�roj,�FD.D�P�sʈ,[ru#�/U�w�x�Q!,D�j��
�I�8ȩ��:d�/D�;�-P��p�ʄO![�1:�l1D��f�O
>��ICѦҨZ^t�9 i0D�� T��gOI5��
���J���"O68@WY�;G�-���I9�va�"O2��$(�x�V�ҦhD�JP�=0C"O�<`�ټE�Z�*���O��`yU"O�j-Yrx$��dL�E��ݻ1"O��!��y-3U%KA�N���"OLM�fɏ �x5���e. �r"O���:!�Y�F w&P8#"OP�Y��X�S�]�O�!c�P�"OV�k�b�x8ғ�ٙM�es�"O�\ӑ�\f��9��L�'I���u"O�qp�0@� ��%M�V	H�	e"Ox���u�\���Ƒ#��"O��3���'��IVňM&:#�"O�\���A�{� ��B�"i �"O��	��B#?*n��P
X7 R�c"O�t3!M�.�����e^���"O
՚w�� FD�e�ܖ�:5ҧ"O�@ӑN��4b
XBRKC'��(�R"OB��a��lhD4bᚄN�v���"Olz�`˷s�z�[E�]|��2�"O<5���?���	�9]�ӥ"O"|�dl�!+}��za�C�!�����"O��K�eҥ)d���Lc�"Y�u"O m���ޑ �6�{ׅZ+r�0��"O�`8#�  ��9��L�&Ҷ�"O~��J�6�"T�#�P���Y�"O�YG��
^�����E�lU "OT���gղ6{r0��b���¸��"O�]�S�+
Xd��KC$x����"Of�HU��:^����G�M[rq�"O� ��u��@��L�	���D"Oxe�#k�2},4@Ѝ��f+��J@"OP���jН2�����B+
�`"O�0b��Iz�؊�;�e��"O^(��$æ!�g�Q/]���g"O�<XUf�0Y`D�p� R�4)�r"O��qE�#��Lٲ����R"O�9y��N6>E����(@+u���
�"O�]�Ԃ�TU�$:�}��(�t�3D�����M���Y'i8�xY�`2D�8Xd�2��]��Y)?�~�3�4D���'n��i:pI�K="�b��$D���jA�!L�	%�R.O"��2i$D�tˀ�Q�*-�R������ D��HA���%ې��%U('!v�{4�>D�`��hM�lS���z'dmr'H"D�X����~5t�q'�
�*a{�'6D���0͔h�T(@f��n���'D�|�qf�13�\�#��'� i��9D�4�Boӥ,<�t�O<�P���7D����7WVvmQ���,S�X!Qp 5D���-K@`�&�'LZ0���g2D��rl��-o\���@J�3-���.D�L��ٽM~`PÆMI?��H�
-D��y��AP�B�Ѵ��x��(�3� D�$V�* �L˷�E�W���d+D�,�q�@��5��,z���*OZٚ�ꗬI�$i�F��=���Y�"O��A�i	��2�*Ҥb@���"Oj��Pd΋c���,&���'f�\��oY�p�♑��G�*`)c	�'���h�2ZV�h����6lh�j	�'�bUb�ֺ�2���LJ�|ʬd���� @(*A��
���I��ބ[ٖmC"O��)��ʥ}�0����C�Ԉ��"O�)�VG�4IJy���vҾ<�S"O� @�)e�J���#[�E`��K!"O�XʧBP�.y����I^�rs|!!�"O��( �p��5�4OS'©�"O������*~H��'X�쀀�S"O�������S�F	����(}f%��"OZ8��ª���jg�G5=�|���"O1"TG�n���yF+��^�PA��"Ov�1����
Ba� 7\�Z�"O�\��Wn�<��E
�z<��E"O����H�Vs���Y�1�hf"O~p�e�]+_w�h��唟|)�E��"O�dBU;�-;'��>?ò���"O~�W���6��L�@�R�5"O$x;�m�;}N��kX�pR���"O�i��ۥm%�؃���-GKJU�q"O�i�r�ߒ1V$\ g�{,�Q�	�'��')Ԣh� ���X��ح�	�'�8��Ꟊg�dс2�V�_
F)q	�'3.5�H�7[�������U�<��'�ƹSpR�M�n����2S1`!��'$U"w��?@��A޼M3Ե��'��i�#&_-Z@��Ȑ,E��0	�'}�D�AD���d�P�X�tez��'
t�*��57`��`�]�e8�')�L
Ѩ�*_�`�7)��
����'~�Ac��*B������7�����'��l*�g�7E� `�7@ /:D��'�@̉�Ǎ�Q.�Ap-��v����'w���FD��\r�`10�ۄi��I�'�^`3��Vצh��/Z{B�2�'F���O`R��g�U�����'*�sa ���lX*��"dx��'0���F	�s���	�_� R�B�'ɖip���b���@�B�
���'���A�ԱMpbmJ�&�	@"5��' �Aq& D=�F��ѳ7�J5�	�'�� 閏]�]Y��"�Q.�&�{�'�0�/���2�@=R���A�'-*���X��L�y¢��
�'�Fmi�X.q }3v�U�j�dP�
�'ξ r J�<�ځY�7t��*
�'�X(A1 ш)&�C��:��4�'��l9�m �"%>-)�mЏe2��'\8�Xq�#%9�Bc�<s�'ꎘ�'݄/D�9!��X�P�0�'�B�c2 ��W��@�N�B��h�',�A���2 ����#PKX�x�'o��J� {:I
"mV"E�B�	�'�d�c� Ea�(����5���1
�'�
�O�ii ��b葤,"�x�
�'���%�Z�L��c�!��	�'����;lnyHb��(yL}��'`rX����ʸ����.�Ԛ�'Y�8j�0A����']޲�j�'����Ǽ0���'O�d�
�'ټU[��\�G�$E�?���3
�'�N�x�MO	A
�`r���IRZ�Q
�'��lX�I?T�n���1����'��鋴���Fl�\)�c��n� �'xFm*�b֨^���C�H�4Td��'^x��@�+
!�DR�h�x�
��� (�6�C7~�4j��N�`�q4"Opd���h�|(*bcZ�t��#6"Of����c�|! "̑�.���"OU�6���8f��@�\=�\��"O���RGISn2|{嫋�&��T9�"OhL[�*��%��A��i�7k|��Q"O�UJ��o��鑪��7�V�C"O�M�VFF?g���3H��%+V��F"O�9֥�8(�����	�%��Q"ORT���<k<"PAa0��h�C"O>`q�g�K�����@��G�<e"O�iDf�&+���1�NȶL���X�"O6m��c�����d�:
�� #g"O�9�`kD	,ۂ�(����QUt��"O�b�P)(��a�1-F�VD(9I�"O&|qpd�6*r�(��757�!��"O,;6$�5_��6��"&긛G"O�UѴDΘ,�"�9g,��5
�Xч"O�<�4��>/���&����L0�"O��a�ꕷХK�@�<-�����"OT �e�.޼�#���'p�}�"Oα!�j��/�a��EI4V^���"Oi9�Iڞ� EQC�S)&}D�'���I�H�嘧��>�0G��G�bP��y`�|��h*D��`Z-�P�z��[:$̲��5ˤ>���
��-y��'A��,�!<�6��%k�,�F5"� �<�*�HܑD*��H7J��b��dPP#Ҡ5M"���"�Oh<�U�*N�:��(�"8=bt����]�'���#KȲW�m*5�1��F�T-A孂�q���ҧ`��bu�B�I%:b�X@#�!�5���P�:�X�C���P8��Z�mQY��,�g?��̤z)JH:ǁ�Hb��u� \�<��BQ9FWl��
���\�7��ݟ�{$%ւ/����} h��D�1�4k�fL=_����t�N�y�F�=^������
�H\5� �[�H"�| �C��$r΅��D

�Ś�'�v���S�N?xE�C#Mܲt�L<���F�,�}і)�\�BL��)���O�ơ�uK�x�V!��A�?�U��' :`�e�(�H�Pǭ��"�l�j``�'[-"��A�Ռv�v}�����O���'����&T�{���"f �@jԌS�'��Ď۝qu I����V�6IgΪw��!'�R�mq�M�
�wp褆��2id�Z� ���!��a[Xz�?�s�]��HX� �mov]�a,[�;�c��w�
U�%�<iSl5J��x(<Q��^}J\;��-.�՘ �yb�Џg��l��C�w�B��#���P���P5�q3�� U���pc���y"���.1 �8��НqL��i7nՑf��<�£tb�1�d	r�N)N~
��[�$0z�Ĭ���ZL�^��c�54Qa�FJ!c��y2�.��E��i@�AZ5x8�
�mK�%�"DoX��q	g��r��x�j��9i"\����
I�}��A���O���|w$��g�{.�r
�"::�m9��N@.��b�&�t��c\V(<���@��[�h�;_n����{?�%�By����7a��ɫb�\��K�韓^n��;�E��F~�P����!�Np&H��s&�U��#l�G��y�b�:h��#@Ś	5��h	��~��`
4h�e��18��d��pe�H4m�,��	1I}�����������ؗt�0��A�:�R���\-��I��g��g9��ǓN�0��u�	3 P�i5��Ul��E}r�]�{��\�V��} u��K� �(�/R�~��a�4��?	/h�4�`� C�	�H��Y�Ǌ�mҔ�{��L�H����?T�L�fl�(Kh�iz��Y��[%�I��OAb�Ҫ�i��5�<� i
�'$T����Ȳ��1�0-"~����;jy�0��H]2׶	�G�ˍ��S�g�e'�,��(�^ћ3g��Ih�0�O��	��O!$p��� �*"IdI�EC�qz�x���ʪ	���5CY>��'�)G��� �R5�Ѥj�X�b���9��u)V+j�*EK��*����eG�U�n�KQoD%s(���e�a�<��M7���[ �ǧ�ȃR�Py��!�^B@�
 1CxMy��M��(���6'�>w�z]�WBO��("O� R���#$Jh�
�(�~�� f�ŁK��Ɋ{���IAL2�3�I.s\��c�)C5)V��� X3[�~C�ɹ.�d49���#Lu�q����#�H��	ƓBJ9��Z>���L80p�`�$D��.�Z��ȓh���pr*�	}��)��6l�%�ȓ@z���hSos2��&a�f\��&"�|���_+o?@ ���
����ȓ2Rz'���T�L��
�� u(��ȓ/h�YV�c�Dp���SNh�ȓC�<�i�J�N�� e�
;]0�ȓQR��� YqR����U
�n���`��-c$��j���ځI�$�ȓ<�)��GInހM:p-E�Q�ޅ��M<�0��J W��	jdbYH�L���KqD<y�+	�'V���5��v{楇ȓr!4��dB-���GC@�����8��&ɤ91�!�e`B�&E�I�ȓh>��PN�9�ht���z!B5�ȓ.'<�cJ�2��5!7k�9��!��O$������]��<���O�A�,Y��	%R�Vǉ�g^��3bJ�	�a�ȓ^N�UJg��[�d����('jT�ȓ � =��bE [#:X �o�?>��d�ȓe,~D0���&~�@��f@�K����:-� �,�g�}�P$'> ��Ge��BROSF�\�p�S<3\\��}�s�5E���S��'�E��j̬���1Rz��s`X����AA쌉!���>�ȤcJ��)ޅ�ȓJ�����N
�2B:����%��ȓ{nlM�b�� %���*���8`9t�ȓ9۴u�E��$�����9,����"�'���!琴q���2~޸M�ȓTl���VJ�"G����'nI|�f5��|�P��a��w��ԋ�,]Bn����?�L��	��
gL�^�P�
�� D�|H�i^� Və�}�@��w�?D�����[����xEO@�y*�!�vO'D�x0��W9$�t�!F)��Z��!#�/%D�l(GjXR��0Xi�-��-j�a#D���2���D3VM�n��I�&d4D�����R�0L攡��*3�i�*2D�La�mJ��{eg��xָ�9��.D��jդE�������'=���.-D�dȥ��VD��u.��R���N>D���G�3<��xp��E-?䖸i��?D��c�aݷ]��R,��(��5��*O�(#���:TӶ��@ ��_�P3E"OȠ��Ҥv���r��I&��h�"OV�K1�56J���E�� �"Od��s���Q���ԋH�u�-��"O�<�-\!Prz|X�
Ƙym���"Or�H�B���L���D�4��0��"O���`�)������3�<�2s"O���F�5�*���8L� �0"O��Ѝ�l� �e��$ ���"�"O��Ӥ�]�.-*�+
|m��i�"O�1�s��q�t�آI��^m��`�"O���Z .π��P�Ո%�$A["O ��6
IjwN +�S�`�dA"O�^
���% �c�	�&!�y⣝�a-:��a+���,<ju�B��y���-@t���+R�b@J4�D�y���v�\�����0I� $��
��I�" ��*,O� �@�dN�-<n�E1sƇ��~�`6�'<�Ų2�R9W����M�XuY�O�>#h�I\<���%z�p衧O�M���[Z�'i(�v	�%^r��sA�v�� X*�Q�c��R���$�}s�B�I^l0sF�0A�" �>^W�7��g͠)(vH�[hM����}��M��,K	��u��'Z�~\cA�Rx�<��X�$�l��IW�>�
��Z�҈��M�~m�3M��rG����HOJ� �;��˰̓d���pS�'_�Ւb�4C��H��I����0��jX��)ɯp���I@�NL���Z��t����L�c���C'% �uQ
�jc�P�q���Cq�a���=�hM`�c�Zl$��wC˭��L�ȓ5� ����+�����CٶQ���RqK�{��b0�>	4�q+UJ�-�h����:��%/�4-�ZɗL\# �!�dA�M�<:VEĿ`G�Q�b�P}��t`�aPH�C�D�,�VxCU7�Ԣ=��[zYkcɂ�0ĉ��^��ǁ�=��<�6K��r��Q�r/�l�� "��F�xp��4.��M���a.6)9�
��k�@y��[�53n"<A��,�H@2���!W���JK7��6�`@�&���
O%!�Ĉ>q1�eA5�NB�k"j�����3GC[Q��`���#������(��s �� D�r��F��?����c��t�<��ꂑɨ�CP�ġ���S��.]�&���9�\4r�L��0���'�hO$�y�$�+`�N�i��-b����V�'�lˤ��7^��B�[:/j��0��
R<�ST������[
��}+)s
(h��L��kѳ�(O1�P��(w 8��ѻ D�˟�c�:6,
"P�0x�MG"O���3H�7�^dI��37��I��	�>�,DJ��D� �:,C�Y�>Q?�$�0|T B�.4Ρ�Ȝ�|!���B���F��$1T�G�X�R��rhD����#dL=St_?#=���x�4�3�4�`��gqX���	ϯ`^
��7�T#Q\X	�d�z�:�Aц�(QF�("��U����`^jT�h�N
'�>H�7k'��(���fܠC��)��
4P��1�)D��J�t!� }��)���) �ti��ID�]��ΡNH �K��)�'M0,C�<d�BC�M�:����.��(��	WJt�"�n�3b��t%��*�Nճb�ay2h��T��?2�J�"S��w�!��6<hZ+�<rTLzr��'?�M�ȓ(�8!8�B*W����4��!Q���ȓw�"$��	�����N1艄ȓ)�\� ���/"���y�EO<UF������T`O_�pmAQga�z��ȓ��h3GI|�u9e��>F
��ȓAtJ��3����q�"-�>�ri��hĐ)��ۙ6h�qqC91#D��ȓT}� �����"��?�����8g���?�Q�u��-ȅ�_s� �q2I�Ԫ�'u���A�"��'R�*�F�`奐�������6H�fX������j���J˺"U�]�#�X��E-��'���ȓ ��ћ5l΀$�B!�œ�B(�ȓkS h(�%:LHIF/ϋ%�$�����*S,E̕���	O����|�̬2��B��(�z��E?OLr��XUTq�BHG�w��%�I��f�Ʉ�%8j���i�FH����qG\Ň�IO��2�+�lնuT�W��*���zEtla�i�*;�ꙛ����o׮���!�ʝqS%@�BFf}s��v���Q�Z��'�F-򖝚@�V;h�̇ȓ5�f�i�"L�i#C3d��ȓnR�x��ܠ��!�60U�L���J2����	Jqr���eصHN�H��u��}Kcc�#0�Q�V��
/� ��S�? L�� /��Дpp
Ax��Q�"O��i�nΘE
D���85�52"O��@q�N;�@����G��'"O
$��J�"�d�T�}1"O�0r0��4��)څ*ښ�ر0�"O��C��+����vN�p/�%i�"O�\+�W�	�֬��ښ~�@AB"OMR&�ǁj�P�zB�۱oh�z"On1��%2z�p�{�cܩZ#j�p�"O"apu"ז@�6�+���3 ���"OdX�4�%&\b�(� �s�
�Y�'�y�$�9 &t����.%t�`��'f�}Af+V�z��7�ȅ�t�1�'�{� g��\��	�(&���'��d�A��P4�bd`!�,K�'8�աrc@�^��4�^*�hPx�'��< o��Nv�@���
� "�e��'?d�s׌��:`ī"J�F���'@����א Wx�6�ɬr����'h��l�2 B��D�]�dVĝ��'A�$�@'�<-�T`� �ޡ^�ua	�'�x �%��"|DꐅɜJ!.)J�'�j�['�]
#o�q1�A�ek	�' l�!���E��|��n�A�����'�L�i����p�(�굣��0���x�'@dᅞ:CED	��H�y
��	�'Cx]`��YF�;g�M�4�C��V<�)��E{�S�O�Z���'�� ; �2���!@"ObEQ$;)wةP�'��.	t�R�@��΅�=}2xYӓ&UKG-*��	4f��N�\��I$�0�Be`��E�BD�a(�^��8���t��!�6n$4��臅@� `F���.�;2�As%N1�i��1��� O̜8��I��lAr�f��>0>�`�>b�!�H*�D�`��9ghX�n��0φ��@NE��ڸ�F�y��ʧ	L�dI$x#t%?`ȉ�U7D��ٓ�E>Y^�p"'I0�r���A�O^軕%��"y�(���G�[�x��ЄB�̒�.K���� �+��<��ϖ.J���RB�ڨe�i4� ϒq"�2)b墠g�
l���G~T��N��|��zCÂzh'�<���+ :�VhN	P���
�/�cܧz��ؓ�B�v{��!��0��#6�HID_�:��ғÔ	o�c�AM���CG�)>?N��v/�aܧ��OL��QvD �B�^V�9��~LT"BL�:�F$���,m�e����!����� \6B���k��=���񤌀Et��$��la���Dmџl��Ȓ\J`�m�-N�A�@P�����뉔a�XD�7,[)pAB}i��>��j2��*�J��\�S�4Âè<!��w�X���lʌ&���a�)Q��%�}���0[,e�T�R����HFg�<�@�C�1p�D�Ve�*x�P`p��"pq�'��o^t��g�I�+*�$?��'�)}���)r\��{c�1ra*��t����?�⁒P�&QR D��D�����oޡW}�X�� S�OJ$3��I	��12�G�4�p<�g"�v�� ����h-�9+�x�''�XQ�K�H�b}�&�4�l���L*��E��ȮXk�,C����4�Ro?�,��Y�E�Z�����y�1�bO��(j�B� ��T��l��|�ȣ��S*V�@��e�=	���Y{6FX�Ē�y�i�"��[B�¯cbfQ����X]S�+;"�>�26�WH%�,�I?Q������IY,Lmڶʂ�MV8 W�B�6��䐵Vv�X�ưW�\S@�׻xD��'j�0|/p0/a�H4K:)��#u8O��[Ѫh���7O�\�ȗ�	����ض�P;�~=AQ�	y⼀�JL�Vm�x���?�V񃔍Ǩ&�Hb�'�H����@�be8X��S#h���'�S���k3��z�ԄR-Zٛ�@ް0��>uL�=5��m@G現`:V�	�l#D�|t�ŔB��り��Y�6X2�D�VP��9-��I��	� (&�O]Vŋ��xR��-\Ozl2��o*(-�� ���p?	���D�biCD�4��`R��}Z���lδ`I�$
cA�%�rU��eQkx�� |��ց�X�@1���������60d�tj�S(���휆6:�h� ��}�bGE^�VL(0dh��yRB�L
����샘f�ԡ#'�����g�5�2GV����l�n�Q>u�qk��a��̰�K�D���Zs�.D�t�`�ƃ2�t�7Jɰu�t;�O5j�`8�H�6�^�g̓=��0��16���-_NHx��RM�u�PF��B����Qi��F��"�ݗg�1"��'QP���ׯgޚ@C��qn0��'��H�w���Z�!c�� �rM��'�ĳfC��8#����Bi:�]2�'BL�ͪ���RgI�m	Vp��'L������,D�H�`�Tp��dJ�<�Y`4\0�iӺn�V�Ff�M�<DV��hmx�e�9���ᓁ�J�<�0쓃m庄�t��:m`��z���}�<a i�?Z�� ���>/�)Z�b�<Q�k�"9�y"�Y54h{ׄ�]�<��ɃF�P����6�dR��G�<A��޵s~�|z�nG��u�p$��<I��-����� ���a��~�<�`1פ�aV�0���Z}�<q�c�(�^�c��ܼ*�(0��@W�<�Ƭڷ��)2Ǚ?�>�+��Y�<�Fϕ�Od��"S�@�Q�[b �U�<��n^ �6T��%Úg��![���t�<�tiU1I9�Hc�` �YT6}[��Ty�<A��@��L� )�f8	��@y�<���95�Y��l��I۾�_�<�!��RI��b�6�"�A��A�<����P���Co�h��t�Sa�{�<�G�+`�n��J��:p��ąv�<פӎ.��@f�^��`�w%�u�<�6�˰5
���ғseT��Ev�<Q�K�D�<�,
Yv�=4�Yp�<�Uo����Q$Ǥm�ko�<��'I�y�0��l���jW�^f�<Q�N�h�����B/�Z DOW^�<�#\�x�R�� +khũ�Om�<�e�A'xDBB���&��eqM�<�ɗ�\Le1 뙢]��)g�\�<�k)1ZG�xcx4�T�TY�<����6N���c
*��	��A�P�<a�!��QS� ��e)Bˑ�M�<�3D�l��2w�K�G���փO�<Y�$�	9�nI؃�_�d:A	�K�<9�L� g��@BHW<��ҕ��L�<��nK<W$�Q
	�X`�
��a�<1�ۢaj�[6�8g���2u�
]�<�
����6Y�#�&^B�<aǡM��&��l�0B���K2̀v�<i��B�[))p%`�]��{d��q�<A�+�3
�hi�qaܰ�.5µ#l�<yL��&����A �,i�H5m�i�<���(�}�M��7fACV��L�<�uF�7f�������iI:�
')FM�<�BD�h���#0+�+N�`��GR�<�U��)$� �	�S��D�W�p�<QR��6~|����mZ�;]@�H�Fo�<ѣ园^�r�2EM�pӈ���^h�<R�T�LX�d(��W~6U�H]�<ّ,�.>�xhaL�Ɉ�a�X�<��N��Nx�􋀻lwL�+�aWc�<��dEQ]�s
�(�1��p�<yw�ą}�n��ġ'9��dK�q�<� �=Ѐ�èk��=����`D9�b"O�䋤-�k+Jp��\)�xzf"O����ƶ6������ʼB��C"O���&	�.!.����oӤ	a�"O��pJ]�9���A֭��0���5"OB����il��!4�(�p�h�"O��քI�Il@�dK�_� ,�"O� "�e��J�'.�F�� "O$�&�)= ƀ��b�.3�P��Q"O��Va҇/���r�<�n���"O<�h1���~�
,H )[��Y��"O�Q�v͐�5����B�5�4�(#"OB���{�l��Aʡz�<Hv"O��	����Ĩu���:�$lS�"O�!y�&��o�HaH#6@�0�"�"OR0��0����Vr��R"Ov�QW�%<E�Ad�xB�hG"Oi�{�H�A���6�Vؐq"O�9�'�L�%�@yPm�<f��u{t"OD��*� 3�F�x6M��\Xd)��"O�{&�^*[�d㠌�HF�D"ON�s��\7%Sh|�V���nl�0r"O\e	�؃6���j�G�$F{����"O(�"Ø w���rS� c�\X�1"O@�y�֫+���/�_䔂�"O ���/@�Q�	S �C(}D�"O(�'�=H���#d�5nWz ��"O��K�a߻Z����]=��	�"OLQ('2��3Ck��Def�r0"Ol ��[�.�bJ]�jf �'"O�t� ���a��ɛY�t��T"OP��G�98��,znM?k�ڱ�"OuH�h��sMұj��3"O~q	��Hu`�6���zDJ4"Ozၔ���u$�@pqiD�i@���"Oj�i�'p8D=���B?���d"O�A"YC �* Ǆ�<��$��"O��27��^�i ��\����"O���?!��L�$�K@�4Ҧ"O�H���/5}���wm3e1��C�"Ox�Q��
C=��C�L�n����U"OV����>y9���PACqy<�#"O`��"�D3���O��S��h�"OT��5��)�]HA��K�<�"O�d�E��j���4'^���R"O�d��B�:CA���o�/Xbe/x!��K�>�X�v�
tr�"T#:1�!�_�/�a����?Aȱ0QBG�0�!�$^�fk|�9�昣]�`�c!a!!��l�2�@�]�(�H��Aʠ�!�O1������Z���r��-F�!���<�W��6��s2N�>�!�1S��-���@7%�R����Z0sx!�D�*ޮl�� Q!x�0�P��k!�DY)E8�-��������<|!��߾uZQ1�LK��9���!�D�F�� BF�M�p�ڦ�Y�"�!��J#"Y��\�J��AOS
|�!���R%⌂��t�l�z�/�� !��>.��ۤ��1yL�S��; !�S�h@�쌉^{�9��.��,R!��}"l���M�Z\�A��My�!�$N�؈�c��+k�
�L��+�!�DSJ��Z2���Z��@+M�8!�� ��[ +L;8��۷�	b�� ��"Oҙ)�l34Ȣ��b��&P�g"O��P�%�L24ы�W ��"OD���/
�+�r�y�MˈET詓"ODE��mG�=�.�n_�7�"O��9���O���H&�D���t��"O^x�a0w��l�&(\<���h"O����ZtT������7T�\P`"O�Ա��CX|��H�;;�X�*"O�|A�D�Nl{� eFܺB"O0)�T�$X"��{�/��1��)�"O�,� 	�8򔫴�Wg96�|��)�Ӵk/L@�Έ%ݚ���Ś!i�B�Y�z�Z'�S���4��珍<�RB䉥J�`�hg�>R2�����y$B䉡>lܴ�u�_-�<���O�	�NB� 
�r0��!MV��1Lƌ�B�I�D�P��;���@fI�f"O 1��G��E`� B= @ի2"OH|b�C	r�liU5߸�ȶ"O\ �Ƥ(LL��C��0Ό�b"O����^J����ՆZ���)D"Of���^#Y�lLR N��9j�4��"O��X���=6,�i�Q�ٙ)�T-H�"O(Qс�ڨ�Fmp�8pl��V�	��� �"AT�n�N�#�.f
����������	�N�;$҉��..)H:�XA�x���\S�O���5��V�[(�9�o�,89x�V��J�If��|�>�u��?���E ͶV��2��Zᦅ��7�S�O�F�0���
&��y��،uD5��)���x�!h6E��'ʜ]��Q4�ϑ�y"�d�$���jIc"MϤ~�}��,��s��_6	bdKǠ�q�8��OGP���߻~��	�FG<Y�
�ȓEs5c���!?,���gLL�%��%�ȓ�(���_*Kb���f_a�~��ʓ2m��f��@kX�i1�.e��C�=hMJX���A�88�c�|C�I)u5GZ2�c��r� C�	�j� b��J�u^��v�(,��B���d`�EH��4	�C�<0� B�I�ikB�`�æ~1�ak�6N�B䉢*��Cs�p]ا�ژ��B䉋�V8�,�n-*��ֆV*B�ɮ~BtX`f�Ĺ8��:���W"B�@����t/M����&�W;~N�C�ɺ�[�K�+B�Ⱥ0)�Eq�C䉛HZhɳ"J�	�=�H!w�RB䉘[𹱷cŮ9�t�#B���ZC�ɝ������9~�(��/?PkB�ɔjl��
�f��	���Õ��'nJ�C��$":	��(R��A���C䉯V�e �� ��#5�4?B��)5x�I��K%bݴ�3��J�B�Ir/�@(AG�Abr*:O��B�	#(�m�P�U��!�t*ː<|�B�I�l�� qR\�)��mk��v~B�I�m*��u�U�o!^��r��=�BB�I�jU�ds��I�-�~W�v*�	�'��E�Ū��i'R)۵��Zh�
�'.(s�Ӑg��I
�o
��|�1
�'R���.Y��Rh������	�'�2l1��(ڥA���԰Q
�'���H�ˇ/>瘈 %FE;t���@
��� �H���re<	٣hMe �Q��"O�$��$ �yBm�HӃQ�tTq&"O�H9&c�#$$q{���j��7"O
(��L[,���c��� [Hh��F"O�<���%T5� �@L3E0t!�"O6�)S�E�==^�����%!?F�:�"O�8d(^/;��u/��}	���""OX)؅�sĞ��v.�?dKz�x�"O�XU(�b`P3.��J��5"O$<�Q F��]Ґ�������"O�,�5�ߔ�&���*RQ�*���"O��C����	�mq4�Ì}\����"O*�PE	��q �Y"4���&r�#d"OR5a���Y��D;�(OJj"OdH�Q��P�d��!.�髆"O�%X�ԟ@����a�(Z����"O���GcI<$P�+g	�n���"O.��5��jѪ<󐈐>�z�s�"O��#F�;��Q�Q290��I�"O҅��̓G���ʁ���F�z��d"OzD*�hU7'�2P ���<���9�"O���$甥muʐ�V��f�����"O���@aԉ��;�'2s��{�"O�(�$o��cV@3�JW�� �"O�86j_�)��iw����@��"O @���ӽQ9�%)1�Ñ-�x}R7"O����\�B�V����R.J���#"O��B�H	d4�+�Á=W��@90"O"��b'W�)�=����*�c�"O�@! ��
8  �eBI�Kt� ��"O�`Zc�L1�n�p�
��8$�E"OⰨc*[�i A�0J\��i�!"OZ��@B�(3DA;2�}"<��"O��Yq�%h	C�A��Hܢ=��"O�����Oj3v 2�@��K�6;�"O������g���B��<X�6�i"O��`�	�?��
֧ol�MXB"Oܜc�휧0�P(�cGM�syi�c"Ot;�ᚵWU`D�f�>�f���"OL�cF��p���_�-Ӳ5�c"O^���"]� �	�� �,�s�"O��`�$��wi\"��6J��@%"O�1{�EA�55%EV'F��"O�	s�+�/U%zU�"�H#W��Ѱ"Ox�X��H"���"�C�4)�"O�@��ɒ����3ŉ�?���#�"O.iAa��[w%Y6h�2w���*"O�Y��
�z�|z�AS*T&H��"O(h@��8>�CV!�?8��!Z�"Od�z���C]�t8�	P�0�r��F"O��C����2��T	\8}"�!s"O��*�Zmޝ��Ʈ��PR"O�SQ+�^��=��>���J�"O��1��! �1�Ƨ>�6�
�"OX\�J������Ƽk~B-	�"O(�*a�OȖ%@�cĴEi&��f"O�\�� �-ɦ�`p��;Ng�C�"O,�V�N(}inQ�u�U/-K@�X�"O�CM]/Z�J��o[8.�$2"OvI�Q%��U?�l�W/JF ��"OnyHP�R�x�kƺ ?(�˷"O2��G+Y�T�\C7��;,�]�"O$R��*x��{JZ
't0��"O����G��Pr�p���cH�I�"O� v ��F����a4�[=m����"On��1��6:�����"-�y&"OĈ�R09�tP&�=0��Y�"O�	)q�F�D�6�@�f�X��"O����(R�h��$�>1�y8�"O��i ���x:nM�ctUkA"O��a�g��b��d�$c]����&"OL����W��$�TBO�[c���"O!�R�N�&QBR!�<���d"O�#�
2]����� U�t
��H4"Ov`��F��I�t�s5 ؼܙhW"Oj�TO��<�bd�� �4�(0Z"Oޡ{�NT5馤���_2C��#�"O̽9FƱrQ �s�73,��y�"O��OJ�� ����аaC���Q"O�8{A e���еaݪe'�8�"Oh`(�BZ�qGU%��>�]r�"O(p�Gě�f=@��P�a�"O�)0�F�p��%blO.@jrģ`"O.E1���8�X��Eןe%"O"%�mӇ8.�:���F�0I"O��q�F�%n(�����r�H�٧"O��&OP5=Iθ	Fc]� �q�Q"OT=�CFl�9��a� -���`�"O8�s�CV���5?H���"Ox�IƟ2i�,�c�A�5.�Yjt"O	�ĭM�h	X���K�=y�"OfQ�a�,*���ɧW���Ӡ"O蕸�傳<�h���=.�5��"O�%����5 �N�=�BeB@"Oz�9aո;]�d W��'��TC�"O i0t���R�lBS&͝R��p��"O6)���_6Z`v��SjQ����ç"Od�y�m[�u�uz�
N�^�N�� "OH�K�G������"��IW`� �"O�4�Hܫ	�0�V�9I�@X"O((	W�)X0�L�� B�� "OB�@�Y'e�5�5"J3D'�}�D"O4قR逭h�Ȕ�&��f�b���"OB��gb����uP%�����!"Ort�'�
�.M�9�Aʃ.��JS"OH|A�o�Q!��K����~m�7"O�-����6P��`W�U��j�"Oz
!J��ؐ��.�J��"O�i�p��|jH�)U�X&6q��"O\�b#�
nq�w��;YCrH��"OV�@j:Gj�h5!��>���"O$�ʶ��V�$;$�h\��"ON�xU��:sT��g ю6_@��S"O�1�V��8�xI���O��(b"OzPZ��H�u� 	k �|���T"Oj��*M*���s�jڼ=#~��"O�x7��nt���&Mm�X�"OTp�Ej>oR8��'�k[v���"O@�� �G�����iQ3�:� "O���F�J/i����/,9��؈a"O9���+5�L��}�ZUkQ"O ��nTM��:1�;^_����"OZ!9G�M����b3�/N�"�9�"O�9��,H2+�Z�R�L�uMX�;"O�u@E�֝aSb<�r땬C>B|�a"OhQ
�g��u��,@C&e%ʠ"O���DaH��2Ɵ� �l��"O�@�� �[	��"�d�uѼ�U"O� �� �ސX��P��:�Z��2"ON� �L��X A�\!�"OXh��I�z��\z7��>B���JV"O����)4;�R�n�34����"O��I��P<jZ�Y"nY[²���"O�!�C�	l��=3c�J�#Ȝh��"O���D<f��*�kVf�@�""O`ɹ�'�;a����"Et���"O�l��%C%V^n����8Uy�$*�"O���:m�N�p�ʉ4Ds Qc"Od�x�L֩Z�2�Ǝ��5s@�l"O(-�n@�o\@3ȕiF�@�"Oh�3��^�	�Ua�m�U$$��"Ol� jD�� ��j�g�`��"Ox�8�G
�\�N��l�9vu�lb�"OJ��.��d
`�#����S�rp��"O��tGX���Ѩ�*!	v"O�-�l��N�b���Fy�q�"O6�ѱ!T17lD@A�Q�a�̩b"O"��J�-6�.��ĭt3\r"O��aI\��qGT �!8"OȘjMW�D,�0���=t�Պ�"OR�i�+a��X�@���>�~��A"O�!S�d����Q�g�����g"O~��áҧo	�E�T���L�y"O&ъq֏�¤H3f�(\�@���"ONX��R�T��恘H����"O�\b��0�� ��\���	�"Or1�Ud�9<��1i���G�<��"O����,%RP�BᇔRؒ���"O�(QEBrvR�K��D�*L�"On����Ў;3M�%�:�╉r"O"�s�' ��DŅ�
��x�"O���r���v>�{��G>]��)��"O q����(��9zT#� ���j�"O�k��ΏA}�X�C�'l���07"Oȸ�   ��     ]  �  �  b*  �5  WA  M  �X  �c  Fo  �z  G�  k�  T�  ٤  Ы  X�  ɾ  �  q�  ��  ��  P�  ��  P�  ��  �  ��  � i �  ^ �$ �+ t2 $9 ]D UL �R �[ �c Yk �q �w �|  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6j�V����2�81�8	q�G��Q�O/�yRL	0���(%�B��a�B���yb�'nP(7'�7@��*T!�/�����'�$ģ�ȑ+�&4�3iйڐ$��'��HSB��&-"m��+�1~�=��'縜P��5f�0r��
�g���J�'��P���Y�X�kG�`�6%X�'l�e�&/oøBu��@(�x�'	|x
��P�2�9���-o�h��'g�$�e�|[z�Bd�)j�ҥ��'б���͆;R��І6`�6�1�'IBk�ݚDA¸�`-�C6`D~"�i��>�a$�3{��t�D)�� 0� �V� D��:'o��jA ���i��H�珹��e�)ڧ,c�1S�Ć�Q
�2���<k�xQ�ȓ	X�@#�mU�or �$)��1�I�ȓd�ۥ��eM����]5W�a��MCu/�
�`�����7��-S� V�<�т^���h�0mےY�3��i�<�t�Q��T;� �:t��HtBP{�<)�#�Y��ةUa�7v�0!�P�<)�JAeZ��g��qtX-�� �W�<Ae%NO�)�¥Ê�L-��k�<Q�e��BAIo�1f@)���h�<��Ö�zgD"�M� �V`�\h�<�d�(/����!:x!��}�<!P@߉0<�h
ؚ\��Q{�<��mudAcPc�V+�� �l�<����PD2���$�%k��ceYj�<�p���!"¼"��e�jIx�c�<� �Az�.�4;�р�EՏ:�8��q"O�XƧ��=y�<�$ՙ-�x�q�"O����ʂ銌�1c%|p��"Oj�� /� _4 9�&�A��X�"O�4jV��8����SM�\L.���"O�h�gF�/\���ǆ��(�b�9F"O���'OW&?���Ku���H�a"O`X�}N���:
ƈ�'�ԅ"-�c^�9���f�<�!�D�`t���+V�ss�:�+��Z�Q��v�d�~R�.�5^f$�1˜�--����i�<A�-��~Ƣ8�w,�0��TD_}R�)ҧ ��S�aW�73���#���D����LuTU�c�E,$���B��~g���ȓe.A @�$k�L�a%G����2a4��o��8��9�a��	
kʘ�O<����+[py��hX&�$��AM�V*!�D6;��93�E��d�i�R ;!�DY2@<�P�u"X6w&��ж��h�O8tm�L�S��<q��%�aS$%��Z7���ȓw����D%X�M�����:f�X��?i�=���G�O�`/���E_�X�X��ȓ#��4�7c��<�i�f��@�ȓW��D��$ލ4��|�#��*(���	p�#�� HЭ T`�գ)�!oa�a��K	���u&K%*���[�ȵTbz���a�����P4��Gmմv��D�ȓy�FݹPK�	-L\8 C�J�pGyR�'e ���ꘈ��D?
\�M�'�j6�1b�� B%��M���%"O
}���?��1��C�q~8q�"O^�`Sˀ��W���1k�"ON)PA��,zΕ{F�!s>0��g2D��Bh��%6lt5��`��Sn/D�hÄ�7L@m{F�۟g����5�8D���"�L8:p�U��\a�,c�+D�`R�KG96�V`�d�3�p<��%D�`�䣚�p0��Ǝ�B�(�KC#D��×�e������Ԃi>�����!D�p��طw�q�F+R�Z�P���9D��P�*ϑPpd��� B��M6D�D�*�l��PvdQ8f�(�g�2D�D�A`�pOPM�O͜iն�J�<D��0R�1o�R� �O�7]ߦ�m�m�<)�+	�e,\�wk�F{��� Da�<	US���$-!�(H5��[�<����W֍��xv��C�+�[�<�����1�@"����v�Bp�<Q2�n�8$IJG���bD�h�<����,��BŢJ,>,��;e.�a�<�ԫ�g��iK��R�_	|���ƐX�<�d�Z�8�  XG��#X�8cVaV�<EC��iэ��Tp�QYש�h�<�B�-��Qx7jӍwE�q�&�M�<�'F�ȰѷU�9��"H�<+�^%��*��s�R�9&@B�<iVJ\�6;
Q�t�����ܐ��|�<�s �&���$��kR �V�Fu�<	�Ȃ�+���qBЁ ����$[r�<�TIH�Q�J�p��7o�d�k��k�<���%�<�jܫKf�H�so�i�<Qԍ0'PF=�f��;�0]8a��j�<(A.4�d�P�T�H�'��~�<��)����U���]9���Uq�<� "ȣ��
z���+��K33��AK0"O�T�� ��H��q��	��"O �F��4|N��Fџ?s�{"O��a�S�^0���妘�Id2�A@"O9C5+L#=���Ȕ���ع��?!���?a���?a���?1���?���?Q���W�FXS���;/c
�R�L/�?����?)���?Y���?����?����?��V$ƽ�g�� ��t*�L���?���?)��?a���?y��?y���?��KΏ���A�˒�F:d"�n��?���?���?����?����?q��?q���Ƞ��H c~|�t����?���?���?q��?	��?����?��ҾX%����@<Ǹ�y�K%�?q���?���?����?���?)��?eHp���"�\A�8Ѣ�e,�?���?Y��?���?9��?��?�6��#����V�ު9S^�*ɉ�?����?A���?A��?q���?���?�BJ�0F��"���&���Ы��?����?����?��?���?A���?�/�R�X�{`�F@&$�i�,ء�?���?����?���?9��?����?�����<��%OQ�U�
��QGL��?Q��?q���?A��?���?q��?��i"X�`6ڛ,�x�5���?����?���?����?����?����?���P_�4B��>=j�����Ց�?y���?	���?���?���bk�f�'Z�j��rrC 2`�0C��	#F�ʓ�?�(O1���	�M�R$�����hghZ�E�$�ڠȏ�Iy��'M�7M#�i>����t�w�E�b9�ؤ+xI���M�@�	�(t�l�g~�=�0m�R�)X�'�̙�7�7�4��O֘j1O6�d�<9���ւL��(�E�8~�|�bo1GY��l�.{#�b�������y7-]�4��q���US���F��7S��'T�>�|�c�I$�M+�'�.�*�EV�i�T�ȴ��2R���ٛ'V�d�˟(#��i>!�I θ]B�=|��2�)�`J��Ey�|"$n�x�t�M�9�T�`FѲ&�L#�GM) ��⟰ڭO��D�O��In}Rn�294z[7��o�b��C������O0 �a�';'1�0��;'��$��xxN�
��D�Y�@(�`�2$ ʓ��D�O?�配�1��9i`�$1�nb����4C1�1�'��7�<�i>�� ��&�duA@��S ��5m�H�Iǟ��	�@�hl�D~b3�p���8�����JH)���VL@0�|�V����H��ן8���ȀQ��qv�(��L�zݫQBHJy2�v�L�����OT���OL�����O��d�F�QT��<"�*��[>���'�6����I<�|��i��y�� �K6av��B��Τ{��5�R��8�?Af�('��]�\3�u7.(��RqyRG�Koz-� ��<�t�U
cd�'L��'��O剒�M���1�?1���lT<��Ds�PW��<�аi��O�M�'H�6M������*@�^�8���!�|uR�(���4�����Ik� ����_�V����������q�zAcCd��T�['m6%��I��T������I֟��IH�'\�Ҁ��c�&�4���Ƃ`�Te���?	�g��&V1��4�'�7M9���[�$aڱd֕K���u��&p$D�ON���O�{  6�0?	%�^�N�R�HQ�Wڪ��6g۹-�`$����'�$�'���'{2�'��=i�$�L_x�rR�5d�d� ��'b�W��4P�@0:���?I���� )]�=��F�07{w-Ɇ^��I���$�O��d;��?��aJ�0:����F.�'�t5C�%��tIabl���.O�iH�~�|rB��t|�6ǁg���o�e2�'XB�'���T]�́�4� `�*5+�Eb�d���B��́�?��#��P{}��'�L��¥�o>�TW�� t$�z��'^2��W ����|���
0���<��<n�rD!aU7PQ�S�R���$�O��d�O��$�O,��|���(QBt,�T�@7s>�;��̏#ݛ&c%��'"���'��7=�
P*R�A�`�C#l��j��a�� ���o.��S���nt扪@.�Y%	�'_Vi㦥׺���I�%�dXR�'Nz�'�t�����'�)H�ʝ�Ҵ�o��[�^�
��'���'��]�d�޴�tP����?���V����W�f�
 ��)r?�[�""�>���i7-|�	�o<� Q��)n�0A�2Ɣ�8���P܌`�*T�Zq|��|���Oh�
��p�x	�f��.B������._��M ���?	��?����h��.jr��M�,w���L�0�f�D񦉐�������Mk��wN�hs�C�R6�+��͟)t�{�'86�Y榁z�45�Vu3�4����rS�0@��m����V���ꜤG�h��Ҏ!�d�<ͧ�?����?	���?�%A�P6~E����h���M:���%y7�O�������'?��	--T� H�n�����.)�ɡ�O poZ��MC��x����Q�% �ڳ/�l^�kWM_�?p��\�na�'��y+ b��� �|bR��+��1.N�\h� ='ҍ��aJ����	П��	���~y2i�p�B"��OX�L��]|������Pw�-HG��O��l�M��@&�	��M���i%�7�	l�f��#��v�Pܚ0���<ԎUJ�J�~[�I$Q⨱;��O�q���� �����T(2�)H#��0p��<OH���Ot���O��d�O��?!����O_�=��+٬bu�6��by2�'��7m����S��M;O>i�j�/K � 2��,G�" ���[�B��'�ҵ��FY�P-��� ru�68�,t� 5Rśj?$���'��$�����'2�'0��fH	�Ub�ՈQ�Z�.0 `�'�RT�+�47۶Q+��?I����i5Bb��EB#-���#�|�	���$���S۴\�����+6�P���L!FT��`�!�b��_����ᗟ�S�b+�H����I�UOK�V��9�&%��Vոy��͟ ����)�Sjy�Faӂz���p�Q#�G�M�
�cd&Z�
+f���O�lA�5�I��M�� �)S"��;��D��<X�B����
d�|����p�j�U �����O>8q�E�2X���ۇ'��[���x�'_�Iޟt��۟�	����It��H�8$�H��H��r�����N,d��7M�b�d�O ��1�9O��mz�-�SBNjE�.6$���՚�M�'�i	FO1�f<�f�pӜ�I;cD(��A�'hT�Â��=�T�ɚ>qi��'��'�d�����'���6 �p/�ً��3j�~��'%��'7Z��Qܴh�2�����?a��Y�0��e���-�.ĩvߦy�n���R�>����?�N>�b�;Y!���Ø9Kv��umO~�)��1���`�i_l��d1#�'��
C����fBM>Vx��`���$z�'2�'��)�'�?i�E��=�t��4!�j�YcdP�?���i�&L�v�'jB�qӾ��.@���!�3c�1
t'�8xD�	꟬���E��¦I�'��H�!_��i�*��(�L��F�%R��]�����D�OT��OT���O���Z-u��q�N��Rt
�!`��7f���քʚsE2�'T����'z��z$��B�*��ސr�(x��>����?�M>�|�@gڽ2v�� D�8�8��CJ��-�v��4oU�	RR�5I��O8�O��_8��!�B�e� �ף1S�4�����?���?y��|J+O=l�5M�~��I�B���A&\�Z`�ѣ��ץ
��)�M��Ʀ>�a�iW6���� �X�<P�Ť��`܂	:RꌗUZ&oZ_~r�H�3X>��tܧ���!�y�j�����9Zu��
c���<���?���?�������-�LZ�K�ki�@$JR46����O����ͦI�!�&�`�i��'u�Q��+�3�h�!��B[j���'<���Ol7=��	�j��8��x9��?a���+���J���iAE�
.:��$\>����4�|���O���Q Y�IIW��*7Ԥ��'�BtN�d�O˓j,��$:}��'f�X>����� ɞp��d�4��0�.?�\�X"۴a��k(�?�@@n>|Nb�8������EU?hP ���K�P�6r1���Ӑ��cK�D3H��t�@ �B�Ӑ�J�X�z����h����h�)�Syy�dwӴ��PK\<Sb�,�?Q�p7̇ #����OX�mZC�5x����M1�	Q����k��K?���h��P�bj�pD��Kd�J�S��2��럜�O�<K�hE�tF����:$�t�R�'���ߟp������ğ�	}�tΔ�a��Q�P��?}��:��ǛH�(7͘�,ʓ�?1O~��N#��w��c�"�ı��gI9u�I9'qӶdo7��S�';j����O
�<���	�PX�g��mb�p���<y o�%tEF�dw�N>a/O�i�O[�둆Sn��*KR:��$C�Oh���O���<��i|��I�'O��'��ò�� r����M���Y�0�f}����!mZ5�ē@";Gj��Q��Pa0��~3T�'��ţF4�d,����l������'"�iP�H��p��R�d�$%��'&2�'2��'B�>�c��������v1ʧ�ún��l�	�M�얮�?Q�K؛F�4�vYI��9��yz����n	(��60O��l��M�Ļi|�P��J2��d/#	����aK��A�ڃ#�(j��IO�d-Go8���<�'�?����?���?YDၣX�t��C���O�:�������ju����I��%?�1k;
��U�ȗ8�R��5+Z c)j@�O~�m�5�MKD�x��t��?Q���@ �A�)�C����`T�H���ٌ����!�� ���kB�O��3�Ա6$@��h��%#`c�)*OH�D�O��4���g ��B��4e"�0;ռ-��dB1"JZ�r�d_
�y�xӐ�d�OԼnښ�M�C�i�4�[fh,c��rP��*$�p�0(��{<�V��LÅ@�&��D�	���ztL� Q�@0��zB�R8O����O����O����O�?1ٗ�<5����/;Pv��q��Sy�'�$7��Mm�ӎ�M�M>3��)�@Ř��àc�L(7�U-5��'&7�D��Sd�� lx~rfT�S��p�R�U�nؐ6GW4qG���7�dY�|b^��ӟ��I��0*�LZ	<%�8�N�-3iLqsF��h�	Fy����A5��O<�D�O�˧�(e�q�̝
�4T���)؈H�'Ө��?����S�D�J�@���P���l�ʭ��f��CU��
��&�����<�'d�@�Ik�I�UbL1���L�D�d�EJ��t��ܟP������)��qy�$s��  �A]�<Q ��S*G�p�R��Ԍe��d�O��l�B��!��ɟ�'�ǳ(C.U*FR�,I�4Xsm�џ4�IuH^�mL~�,ʀK�������� r�*�-�tP�����7NL��2O&˓�?q��?I��?����	�& �h5��<����D��
3�n�f{<��������i�':웞w�����i�?A'��0�f��nRЕ��#m���oڋ��S�';�lPbߴ�y��)`�F���R8L�P�R!�G�y"j��}%&��	-��''�i>��ɓzv���O���2�JC�E�̍�	ߟ��I��'(�7B�C�4˓�?��̓�Z;��ɧ
��@�c����'�`�9��}�,&�hP +	� �5*S ً&�(�D??AT&V�%�\i�TbKf�'(�H��I��?�`,�#*���甩]���Cqd:�?���?���?���)�Op�e�#N��SUʔ8]	�u���O��lw�H�������޴���y�@�A��Y�ȸO���xpaM8�y`�r	mڭ�M k	��M�Od�������b4`ӶN�
�	V,Y��P�$&_�4�O���|���?���?1�E̄rwf\$T;$2w&��=��m .O��o��ZfQ �����h��'���3F�B�pG/�A��)����ۺ2�O(�mھ�?aH<ͧ�2��V<�C���V��I��֛q��Ӗ[�$��+/O��%��:�?!��5��<Y�d��V���'���>�YP�Y��?A���?i��?�'��$K�	�7
�����r��Kq�m�7�ʺ&w��K���ݟ�K�4��'".��?��?Qr΃��@l�D��kU��'�Nb�X��	^~�O*T^�i�'�䧧��I/�[�A�pG,|�掃�<���?	��?���?Y����K'�6���6W��i����}����4&,8��OH�6�9��30=)Sj	����!�H#J�O��O�ɇ6.���K�8`"���,	��]e��Q�J��fa�`�Op�O�˓�?��?��$U�X�����U&�C�z)���?Y)O��oڻ*TP��Iʟ��Ic��*�[�qڥ�� i2`��Ȕ���|}�h��o���S���@t
	�AB:�� �X�R�� �!�@�D�g�ý��4�����qqf�Ot�:�&LX����"k���D��O^��O2��O1�H�w����	!tW��Q�ނ#x�X�
Q�xKG�'�BMd�^�H�)O�6M�3}�	���9:7ڜ�6&��c/�QmZ��MC�	�M�O�����8�"N?�X5�	�tK���
A�U�Ex���'-"�'{��'��'��^#��X%�U&`)�T���88�� q�4����?I���'�?!��y׋�ˢ�g84]�:�!F8,����OR�O�O�\X�i;��qj��hQ��r��@<5���ʮ&�Y���~ޘ�O˓�?Q��`x�"��چG�=0!��+�������?����?I(O�lo�=a���Iß��I�H��h�N0~���4'ׂ&��=�?i6U�4`ٴp��xBl�'^�I3�b_���c�Ʉ�����4�쵛��	�������̊����&^`�e#�8��tk�)�~$����O.�d�O���(ڧ�?a#��]r��*��X�;�Æ�^��?9�i���4�'���}����ݲ%'̖2"nӖh�=5ϰ p�2O>��j��oZ�tp�lZA~��gR�S3y�£B�*G�����\8�ʆ����$�O`���O����OV��DF�9��K�@�EG`M�Rf��7���hb�'�r���'1(MA$�QF��24�ܝy�T�rO�>��i�7mj�)�Ӳ� i�sʋG�p��w)�6e9�%�!M�$;sf�o�����O��pI>�*O��/��M�ש�9�@�xGk؂GM�'�B�'��O��	0�M�4,���?�e�Ņ37 \@���*�ָ� ��<i��i��O���'Ԇ7mئɢ�4o��!"� 'X�,x֫�"/��p1��M�O�,����(������w� P9�@���j���R�Ѫ�'r�'%�'��'������I�\��BU&6�d�W��O����O�n���H��'��6�?���9
^$R%*�,ERthW���'�$��4"��OX%���i&���s�@��I`EFTJ-v0�!ВH�b t�IRy�OP��'|g� w��Q�!�M����@�0d%�'M�	$�M+3!�;�?a���?i.��\rЅ�1,�.��s��-i4>�k%��D+O���r�8'��i�,�z���	#5�%�)#�J�ʘ�-ZX5#��HRa���?�J��'���$�����]�?@�t���N�jLQ`7�Ɵ��I�0�IПb>i�'z�7M���Ȥ _�u�L�)�z���Q���<)ռiG�O�L�'��6m�7ݦdR��ӭ8s�9b�׫^_&poږ�M#!�ڔ�MC�O�l�Ь��K?� ï���<��oMV��ɠ�m���'r�'%�'qB�'f�ӳ)p�x+E�D+z�H��hM�l
�4��H���?�����<����yG�ߍZ�T�39%q�]X��D#d�7ObO1�Le91�b�J�	!R�Rta�E�G>*X�f��c�D��fX8cD�'���&�,�'���'���I�+P+?���`� [�dE�'���'y2P� �ݴk&����?��IZP-S�G=A7�<A�2L��4����>Q��?QK>�5oGC�T�'�T�q�D�x~"O�1���ְi�ⓟ�u��'���(3m���E��{��=��0B�'t��'"��˟tQ�#Er����<G�����Kԟ$�ٴc��<����?�D�i�O�O+n�8��/�T�2L0�&;c���Or�d�Oҽ��uӨ�L�i�N�?� 䰐�G�3^{(�P�HX�Ep��j'��<����?i��?����?aS#@[��e�p�͉7XՉs��$��DH٦#0�ݟ����h$?牃8����@P4(b�Q0��``<!{�O����O��O1�������H��;�(��������7�My��ހp��������䂌B���I��
6����`���0>�b�i̠���'\�>E\1ůʛ<�������ğ�۴��'����?���?1C�D�0P����⨬�5� 1 ^y�Ef~bk�>r��'�䧱�{�ф)�N99tE�aZx0��-��<���?	���?i���?)��4�I�O�Z��'ɘ���@cȜ!N���'|B}�LHK�i�<�u�i��'�@ Y ,@4c����\?�a��|��'��O��+E����d $3'Q2hi��YF�z���6����������O���Or��/E����(�%�d��ą�wNL�$Uwv^�=L��e_�W[���'9��O����E�sB��Qp�Q6���1(��y2�'��a`����O�O�I����j�#�#�$0�F)\�!*�[�Ĭ[:|ɚ�HEh�R˓��+�O��O>�g�9=�g��qd�}�u�3�?����?����?�|�.OXl�B����p�	�5��ֆL���f(ZYy��{Ӝ� .O�7���Y��I��P �t9���B�:��	ئ��(��e�'u�LQ�H��?5��^���D�a���`��QY��p��v� �'���'"�'x�'f�S�!��pk0�׍aUN�H%)w~0E������?a���?1N~�1�w~~�h�*�o`����>0�d����gӘ���^�)��_�Pl��<y���pA:1s�a@�Q>&]q�G��<��S�$ӕ������O.�$N/C�*uHG���@r%�*|h�d�O���O�ʓ����F#v���'?b��3�#R- A̴L�vbH�>��O�u�'r�'[�'P��(rF�c&�c� Z �"!��O(L:��F�I#�D�#�)���?A�'�O:8:�ƀ�v��Y�/8�I�"O��v���g"���̷�lb3/�O��lZ�	�T���ٟ���4���yǫ��|�(�[t*�E'H|X����y�'�R�'Y��s�������/�Y�O�b�ɂ�D�` D�`��(Q���	��|RW�h�I����	֟����D�$A�S'j 	��^�'R���HPy�ab��-����O��D�O������H�~�A7�S7}�١C�����	�'|�3O>O�i�O>�iI��ŗ?=�HH1�li6fg��|2��@ĥ�t�O���M>�,O�J5�43! ��BÛ�AgZ�ٖ�OL���O��$�O�<9��O"�aI�j'"]9�D��h�P�Қglɸ�5S����US}��'/��d���Q�lM�aB�Lc��: �ء���"t�b7-$?q�
L�8v �)���'��k���D�E�r.����Q��<I���?!��?����?Q���k�
$��X��C�-ݖ�-jd����?���Ey��H���ɧ�MKL>�C�����<V$ y�O�8Y�'�46����i�=%T7-2?�OD�{�^uR$-�<���##"��\��w��O��[J>�/O����O���O�hc�H� ����ܓ@�Y&��O�D�<E�i�ف�P���	}����xd��D�1�~D�Q������E}R�d��Im���S���3(�>�����cA��Y�X;$َ聲D=j�(y)�O�	�+�?QR
(��h0�p�H(_?2q���"D��D�O��D�O���ɪ<��i�� �<��b�?PT��ƒ k�u��[�h�ݴ��'\T�UқGM'+2Š���,"m��
�j�4v��6M�����
�	�'?�eIF�?�����hUed�Ή9rK�Sw���b=O^˓�?q��?A��?����iP�j�|����=B�^���Ó!40�]o�	Tr\�	ʟT�Ib�Sʟ`����[�I�*����͟,x#z�0���e��Vky��|'�b>Eb�ަ��G]6Y���(c��2�"�>_���z`��a��O��I>A*O�	�O0��D!(��,Ɫ�����"��O��D�O���<�e�iάQ��'�b�'���ڶ���%�n��q��W�D���DX^}��h�X�lگ�ēRa�xKtV�WάEI3/��,e�'��5���C#w�*pҏ�4���X�G�'��l����;>aNH��ϔ!m�0�KG�'���'���'��>睜LG<�� �p�\� gL��E.�O��l(Q�^��	Ɵ�:ܴ���y�����c��'ڜ2Uʙ��y��nӢ��	ۦ�GJ�⦙�'}�t2���?�)�gJ*��p�g��,�)��Bm1�'/�	̟��I��D�IΟ8��Y�,��t��:F`u�`Ċ�j}|ݔ'�|7�Q�"W����O���=�9O��#aAZP{�-����_B @�BE�{}�Hi��Id�i>��S�?�(��D�4B���#$�v�e���c�fqI��Ny�iO��E��Kq�'��Iu���2j̯�)���a�0I��ӟ��Iݟ�i>Q�'!6m��b���±F
\�����RA�bʵL�&�d�Ʀ�?)EP�D����o�5�da�눂|,�x�b�G8�	�P�Φ��'�X��f��?�:"����w�j(�F�Q5��p�b�*T(`��'���'"��'���'����`�T�
�YT��К�/�ON���O��m�Z	���X��4��p�"m���q6��uのk�(|KW�x�fӮoz>aq�@��9�'�.��� r�dU�8H	�-\;6� �?)C�4���<ͧ�?���?������H�8�U��@�?����$Y¦�c-�ȟp�Iߟp�O#�{���@�NMa�h��mz�E��O`��'��7m�ަ�K<�O@�0�1N^�5��	+���c�fͪR$��|i�#�5��4�8p��aF��O��qFȑ�^�|��3䜀I��n�OT�$�O��d�O1��� B���W�a�H��#���  �LI��z���'���hӜ�4�*O~7��`Z�|���(nH��W�͘q(	l��Mk�BA��M3�O�t@�,�)�"O?=����Q`�K �/$���Ac��'�B�'o��'��'���+�4!f	A��{׀*�HٴP�*%h��?Y�����<1���y'��7Brn��4!�R@��Ӈ	;}�:6M�͟�'��S�?�ӛ��lnZ�<	���-���:q��&h��H�@��<�򯌮Ԟ���䓖��O��DG|�(�*u(�BmȔɲ�[�+�\���O����O�˓-��VA�76|��'"���8pHx �Ļc] ��!��?�O�l�'0L6�ɦU�L<Ya@I�tP�郢�ԩ/����o~REK�Sʅ*�G���O­���o*"k�|t���%�S�GR�;Gŉ�]�r�'��'N�S������[��P��8AP��L�̟D*�4&�5��?�ײi��O󎗓e�j$�R��w��j��DM�D�OF7M��%�1�k9[v��|9�Í�&��􍞹	c��H��M�CA⥮J�G��'�P���D�'B�'Hb�'�(HB$��x�l)!gnA&l� # X��#�4U�T4y��?������?q�LU�_�x�`���d�怙A�J'��ɬ�MK#�i;�O1��1�eX�3�t��w��-��"��F*/�T�h��P���pS��'g��&���'!�}JB�?�±r�&4|ԋ�'"�'8���DR��ڴo�D���-����V���N�΅k	��M��X���v�[i}�r���o��Mc�)M=:Z��ʢ#�lY��i����z��ܴ����'Ъqr�'�O��I�,$Hg��CVm�3��y��'J��'2�'��I����A���Sk��b�M���7�O>��榁�)RZy�e�(�O@L�$���%K$�;��Q����D��M��ii��֊�̝��'�"bB*i�p��4N�v1�5���pZ�+#j�ܟD`��|Z���I�������+`�ĺ,����#�<1# }��M15xy��f�F)r"�����O�����%�ՍL#���rG�C	L:��4O����k}¦o��!�	X�i>U�ӷu�z�r�c�#x�r0����QphZǯWČ�wMqy��O<JH�I7-��'��,C��\���8ŭZ;A�b���'@��'�B���R>}�'��6��#�����S�h�kpH�)8�!��Ol�DR��I&���ɯ��n����SaF�Z���h� NÃ�٦Ձ�4��rߴ�y��'1`=�D��?)q�\�Hⵆ±&��e]U�&��d��'T��'���'��'��(d*��;AOUx�
�r#Вx�d���4E6��)O��D5���O�oz�9 �g�*������>|�|�0i����	]�)�Y��l�<9�e��*#��A��u6�9��\�<�2��_�`�ID�	oy�'�r�N�*W�9�c"�օ����HI��'��'k�X�0I�4A���z��?����D��3/ƺN��P���ð#�4XA���<���?iM<1r�J�!)���A�7*Έ�5ȑ~rk�op&��e�N�Oy ����NG�����6�5m׼�[��;4�B�'���'��	�O�NP%7B��!.g�f��կϺAQ��æ��l�my��r���$�<��Ӽc%�&#�p0ВP�k���S%@��<1���?��iLv8�i���y��'� �#* �?��4.Nt�����K�|��Y`�]���'������I쟸��۟P��5D���⤋��[���:��F`�d�'�
7�	�^�D�O~����`9�l�<G�
� ��D0g(`����x����M�b�'����T�Oy���L�!�P%��/En�C�D�4�Uゅ��T�DQ�'O8��ԟ$Օ|�]�
(B]��D��Lip����h��ݟ�����S^yboe���N�O�xjqfѡcS�ɶ�B�I�V�?O�dn�_��C�����M[7�iY87͓�j�µ
�G�1�Rؚ���/+~4��ob�>����9����*�>q�ݫ$?� �0��f/\�y���Iܟp��柸�I㟈�IK��s.�`$ �)�D�����jw��!/O��DM������l>5�	%�MK>)�ǣY�`P@4)E�,ϛ��?�DOr5o�
�Mϧ{&.���4��D�:��#	�Ntxղc
$��T�����?ID�7���<�'�?��?�֭_6|��#F*��.�J���.�?����Ӧ9�v��Ny��'���$A�xM����E8�IL�n4�I� nڶ��S��4A�@��aP�@�1�PA�FKؐ����=���O�<�?i'=���?bF�SQ�"g��]3r@�<b�����O����Ox��i�<Y&�iߐ�0�mC�\	���U�A)HO�x:s�ϖs���'/$6�(�I:����O����pJ��H�K�)p:�e�O��Ĕ8�n6m"?1C��i!��SUy2��:#$L�����`Z�u�E�ޏ�yR�l����P��ǟp�	ٟ��Ol��A$��d��A��M�"V^D+�#n�8�*���O����O������[̦��$A�}rtÄ�S<j�� �<d(D������'�b>]�GL���S�? �݈�(K�@���p�ߚJ�1O�t
6,��~�|�W������zw�H�=2B��/��\�r$3jF������p�I`y2!i�D���"�<���"E ��GՄ|eP�
�`�Jʎ�s�2��>����?N>)�qEε)g��+"��)3@��K~B�%W�J�:�iM������'�үO�������Q��)��^�-���'���'�R����j�\�X�BĔy��| �f��p�ٴuJ쌀*O (m�G�Ӽ�s�6G��H�gO+M��)F��<q�iI�6M���͠�M����'���í�?�6�E"gj�uu'H2S�I�CSR�' �i>��	۟d��ȟ(�Ɏ�Z1�ܓ#�z0� �ƈ.^0��'�6�Tt5@��O ��)�9Of��tB�V��a(�-~A���O}�Jc�bl�-��ŞD���u+M q#�#�/N=<� �3"����'x�"�I��7�|�Y��!o�0��1��
r5��A��ʟt��ݟ��	ٟ��pyb�zӨ!��A�O���@O�g	>k@���^������O`�m�E�;z�	�M��it�7�G+S4D���@�E��Yr���z�A� |Ә�H�T2���H�>����s%�p*��P�O�x�V��cM|����䟬�I�0��ӟ�'?M���H��9����qk�`�� �r'������M�&�P ��d
̦!&�|��C��}�sA�����Çϧ��r6�F�oӬ��̗��ݹ�3O"����z��Y&ץ�4����P�g�\�!sG���?��l*�Ļ<����?���?��f?�zY4�<B���CvEE4�?����S٦AD��ПP���8�O�j��DLM�?-�%�f�ȭn�A��O���'��7��1CK<�O��rD���(�Lq��+�"~�rd"0�G��x�c�5��4�4���n�t�O�qqg %	�X�A�9\�*,S�.�O��$�O����O���vd�'��6-ʸ{}p117�X$���id��n�ҝ�Ǉ�<�0�i��'��$�>If�i۞�B֌K�t�Ε�/�1gܰ�#'�y�umڶ#�@)�v�u���ɳ.ґ#��O͜Q�'�č!FF�	}�&�yt�4f@(�'`���$�	���I���IQ�����z@��ʌ$j�@�B&O�N7�J; X˓�?�H~J�|��w����K.Q��}�Յ�%]�\�Y `n�~emZ1��S�'m!�5��4�y� g��׊��p{�ѽ�yK@�y������G��'��i>Y��)g5�y&/�3uϾ�Oϲ!�p���ޟd���l�'.�7��L^@���O���H�A�|H ��U��s�Bw$(�I���D�Ǧ���4;��'΂̸�fT� ���6'G�=����O@	�e�ǭ|?x8���	-�?���Ot,(�j��NI2�:fG�T���Ox��O����Oڢ}λ-��ق1�'y;b���P�SS�%���1a�&!��b�'�7�,�i��`6р7�:�p�m��{��j�43�f{Ӹ����G�q���lg�����O����*�8Tp����L_H���8p��o�IOy�O���'l��'��e�# ��#�Ë l�\iǖ�^G剅�M��	 +�?���?YJ~
��|(<�.�J�sQ>i��Ez3e��6��(oڙ��S�S8+��}X���8bU����p�>���a�ufX���|�å�OذO>�+O�}��!5dI�G�vm�e�C��O���OV�$�O�<�#�i�d��S�'�8���CC�A�;c����'�6�!�����Xæ2�4
�V��I5 S�bO&h�Ŭ��
��3A��$��$Y�`x�{�'̸O!���CX�Bi�%a7�|�%*N�yr�'���'��'E���D�f�h�H Ȝ+q�1�%��J\Nʓ�?��i�b	�O�vӲ�OraZ���/�ȥr�*�8.��\�'�f�I��McQ���d^�@�P9B�Oxa��i���Y�����v�譺�@6\,�8��\;ؒO$��|���?���`�2���Ə�{-T�p�+@O��H���?�-O��mZ1�n����Ia�tGO�,Ɉ���h�_"X�Ӆ��I{y��'y��(�T>�I��
U������K9Q�ĉBֆ��N`��Ī�~��|*���O0� O>Q1!R�:XF�R���+N�=��*	��?����?����?�|�+O��l�7}q�a
��T6(���e�.-+��wyr�d�B�۩Oo)Ab*0�= @
)vMúSO��4E�6o�1G�]��O�q�݀��N?]K�Ē�@z��Pl\
&\�7)y���'(b�'�r�'���'�S���}��j@�'&�#4�A8Q���شQ��	0���?1����'�?Y��y�N��s�8ʣQ����d(

,����s���$�����4
;�D߇#�PA��x��E�Ci��q����XĨ]��9��O���|j�m�ʠ������l��R�i�@����?	��?�/O�`oZ�Hl���	����	��}��nK+�)X�/ؕ$Hd�?�tU���I�<QH<��.��r�
"�5C��Хe�]~2D޴m�	j�kK&
[�O�!��$
�H����h���n�d0P��~�B�'�b�'���S�l8e�ʎt;����G�];���3bğ���4���(��?閻io�O�n��3�u�"@��M����%Z�$,��צ�Q��M�BK�9;θ�'��4�M��?�i�`Ԙ�͈���`����@�.E�'��	џ���̟@�Iʟd�I�V�� ´��
G�@�;�NF�Rd(��'x7-֠u3��$�O�%�9O2M���b&� )��;�.X�KC}2�h�"��	@�)�S`4<� �9���<����H@(=��髶DA�6=�� ���k���O��pI>I/O�0;�F�5mk��K��[���� �L�O����O<�$�O�I�<Q��i���s��'�l�D��0_
���+[����'	7m+��3����M�ڴ~�V��:b�>�S5@)f�F��5f	*�` �͓����̪_Tx�a�'�O!'D	�6����6\܎�yč@��yr�'��'���'wr����#��pr�I�//�� q��=6,˓�?� �i5���ɟX�n�F�G�^�e�iAZ�u��Z�`L>���MϧZJ��3-�S~��њ�\�C.�a"��,�!6�]b&������'��ay�O��'�2ȗ@�(����,z���^��'V�I5�M�W�L �?����?),�$�-VpdP��T����2��D�n}�q�d�m���S��ŕr� T�S��8/�����͌�e�Y9P�tH���D~�O�H���	.�'�2�KV��9g�ׇl�1R��'#��'��OB�	��Mk@KM����D�X;%����D�"_z��(OAn�U�� ��I��M+�도Iw�U��;J���(B�����n�z4���&���:g*�B��OF�K�P����D5�D���1J������D�OX���O8��OD���|zΒ����)��|RF  ��-ӛ6 ��;���'K����'�@7=�d�X�"�U5��k0���>A��B�͟�mZ���S��6K�E��i���l�k���V��ҵ�tM�$��&��k�� k��My�O��U��@@
2#��w�Y�?�B�'���' �	��M��ӑ���O,���c�cS��ـ�=*�H�J��#�����d�ަ�۴7�'���Ί�75��i�*�tw"5q�O`h���S�c��@:��I�1�?i�n�O����^x[*(K`�Юx�pu����O��d�Ov���O��}
�� ����#��=�]ڗ��jc�8S��v��F])K���1�MC��w6F���)T~�|�d�BT��'�6͓զ�޴N�J�1!Bt~b$:BR��YTj4FBQqX�����;b�2ձT�|�T��՟��	ߟP��؟dk⇳I��C�.��"�kgyIjӐ��u��O0���O���2�D�$PtBb��4{|٪2o��X5�'��7m���K<�|Z"!	j����ȈBE%�V!�9G��+���F~����s�x�����'��X֔s�,/{E����)��5_��������C�џ���Q�/�PL��k�*c<�%S�����ڴ��'���?I���?�wcȎ�&��6�9:ct��d�-=�rx�iBG~Boɼ[�l�'�������D��k�`ƈX!���<i��tI��*��)Lj)�
<x������?�����m	����Ԧ�$�$��AU�b���W��_�]����R�؟\�i>���Ǹu��$\���7�04b�ٛR.*D�Pȉî0p�h��F�Iyy�����Ġ���&�U�ŃN	�@0�4� �;��?���i��/�ڰZ훧r�TIKv"�-%��I��$�O���-��?2�,��n� �)��W�j���d�!3�2LH�,�B��e���$ r?�N>�Voқ�r -M5n����V#�u<)t�ijĝrU�Y�O������:P�1[�*�W ��'&�7�*�	8��D�O����E҅w��v���p�l:���O ���:�$�K0��D�� ���	�<IPG�>H�4��C�2�� ��*�<�,O����rҨ\��"� ,��P$d^	(���m%ZR��	����	H��;��w'V��G�_�UP��Q!��$�X0�v�'"�|�����7�Z0�'}l�������UiЊ	/�<�R�'�<!)P�\T?�M>9,Ot���OL ;$M֢p|�s��G���*�OR�$�O��<闻iy�Q���'�R�'��b�&%���7F�AЁ����}y��'���%��C*br���C�4hA�) `�#
��3id��s)�3R�b>�S��'F�|�ɊQ~F)�#���0��T	����ϟ���՟���G��y�喤R��p���ח[��iK���[R2llӚ4�a��OB�$]�	'���i�	V�ˊo�d�x0)�-i���[! a�,�I֟���>�xV�'?�%흖{*�S�o�)�B)P�nZ4��F�8��%� �'m��'q��'���'{��@��LA����.{ي��T�T�ߴ�����?����'�?y%�E�D�|<y%�^����t*����˟���d�)��"> �-p�hB�%ԡ�K	}�n�2CE��7���'$���T?�M>!-O�1v�@�3�>� ����^ex���OV�d�O0�d�O��<a�i[T �58O�	��N�<v-����B�<�Cp�'W�6�%���O�i�'�"�'B�9&��PQGG�#۠d�� ׊ؒP����A�5���O<�OQG�[����
�8��&��=�yB�'�b�'��'���ݳR����*7�@A!�[X�����O(���ݦy���q>��ɋ�M�K>���E�0�l0a�J�V葚������?���|j� [�����'T��I�&� K�D�����.��TJˀ8}������M����?q��&[P���g�S����gF�]�p�����?�,O�uo�.4�����\��n��=;��a�)[�d�k�,M�yB�'/���?	���S�� �9��^ov��-��h��d̚`R�K%�Ժ@�b��|�寵��'���c�$5����R	�`Cg��럔�I˟,����b>��'�6���)vpQ �KFb�>�y�]j�hu�q��Ot���٦�'���ɤ����O"��v�V?#�@�g��Zk(�3*�Oj���.m4��������d��,���<Q 99<����Fj>,�	GC�<�+O��$�O8���ON���O��'Xh�BD)ҍ>+PIrl��|?��!��iHN����'JR�'��OB�$d��nW�y�ĵ����<X�䉓@@! L��D�O��O1�Թ�s�! /���m�M0���]��A�P3G,���#X����'	�'r�	t�I/
lP�����>~�	���"3L8�	ݟD����' 7-W�8��O�A2z�ջ�?d��� E�Y86�� ��O��o�M[�x�ԏ4�u 3�;n]�`�'T����,��`����:�1��p���0����]n}�b	N�����3��d�O��D�Ot��:ڧ�?A�hx!~�xG��TE��[p΂�?15�i'jix�Z�8��4���y���V��i���I��Ź&(_6�ybih�6uoZ8�M���W���'�������?m�0ς�P; �j��ҁP�F�Vo�6K��'��i>m��ǟT�	�L���m%NasEl�mI��+U�=�J��'g6M��q�����O���&�9O�8��OU�B�~<��G�<�>� �T}�y��m���Ş+�0�e����hq���A����"`֦J�B�'�T���@��
��|�T�(:�	K*~:�O^c}�p	�����I�4��ڟ�by��~�8)�OB���B܇��݀B�ƈoB��B�OPl�}�w�Iȟn��M���ΐ@a�Mהko|u�U��O��&�i~R�/U$P��S{ܧ���5�Q&h P�c��J�R��F�<���?I���?y��?Q����&I6Q˅gY�%Ϧ�Z��@��'t")lӒ�R��<�U�i��'�4K1�T�+�"���L���%�!�D����B��|�%T���'��IaE�c�P�2�M''� �Yt	�[M���I*3��'O�i>=�	�L�ɚ_�jH��1sX<-#�G�
��O��<�ƽi$~ѣ��'�r�'��S" ���&K���O��H"�.����m��S��J1�H��	�
U@u!�o�5k�����+4N�P��O�I��?b�*���:!)��H#ȑ8MI��I�L����O&�$�O���)�<���i#����]v����5(Z��17f��r�'P6M*�I1��dXڦi9��0D����.˧vX��B�����MS��i���K�����":j�#�'��S(g�<�"1+Q2�v�x�씔'<��Ioy��'O��'��'5�V>�g�-<���+2`�5<8pe�eI�(�Ms�'��?����?�O~Γ/���w����Q�ҧT�^�cB=����El�*]nZ���S�'$*xxu��<2�E�l*��Q�Ǥz�,�'�V�<�Bޜ�d��͂�䓙�4�����;=,0dC��2g�|c�J�l7�d�O(���O|˓+�F@�@��'�rɏ%/n���ӌ�17Z��5�J��OJ(�']�i?^OV�Z ɋ5I��)3�۔#�ܵ���\�mJ*&k|%cL>�,$aBM�ʟD`@(S#Q:|�b�H�Ziy�K\ß���ߟ��џ�D��w��Xs�}&�҅&�L)EIH/v�$ԦQ�0��Qy�k��杁<��mD�m�<H#�Ķw�"���M+��i��6� MK\�� ��|3SÄ�u��D`�$r�xU
���#�z��0BA�&L&�������'$�'"��'5��S�DY�%��V\�	�P�Ă�4u�8����?a����<� B� 	#b^�2&��ZqI[6m<�I���lڈ��S�
7$	�  �g����ڑ2t��+��ښ��!e�)��O[H>�/O�t��ć��a���_:H�`"��O��O�ٴ�?�'��Ēߦ%H0b�՟����#M�J����#"�Dx��M�!�4��'�4듇?���?����c���R2�ɉ\{��x�&�j�P�iW�\t~�fM:z����'��'Ϳ��b�N���9�CM+F9�����<���?9��?Q���?ь�$#L:S��`���~��f�Ƀk7��'���aӜ�c=���D�轢&�(@��Rj��$��柬{Yجs�+B���,�i>�
��(Ll8��]��� Q����)Ǆ&�b��2�ُ�h��]�	Iyr�'P��'9����bm�"�g�9̹K�W0D�'F�I�M��.��?���?�(��qۡ�J�k�m���"c�1ے��<)�O����O��O���>��X���=03DX`q*P �h��C��z~�h3#�Wy�O�������*2X��`9J��|9��p���?���?I�Ş���ϦQUL��8��8Ak�7�hq�H�9O�X�	Ο���4��'f���?!u�,v�i1��-G
��RJ@�?���S(رc�Pp~�Ŏ+-����'�򄝀v�8)�7��r4d�#���$�<���?���?���?q*�^Ez�g�y=\�PQ�P�\C`n��M�Ɖ��8��ݟ�&?�I��M�;8�ܜ8�L&|��	w@�~L�����?�O>�|�FK�LΓH1���W��b��3%&�e���%�`����%�L�'b��'�B�2���oadxȀ�	��Hf�'�'�"X�L�ݴ$�`����?Q�{�.U`�dA-J�4�����`)FԒ�r�>a��?�K>� �L߀C�a�r.T{���s�������=#ȐU[�d@m�#����O�$��Õ�P`>c7MA(ZX��ӓ��O��D�O��$�O6�}���H��Py���8��)���x�����)���ʛ�e�2�'W@7m+�i�Q*b�*^�|�;e4.�8 g�P��ן��I��r�"b�"?y��Υ���-��|�@�Ե![F�zU`�
�LT$���'��'���'jB�'�� D=F8��#3	�`U�Hp�4g�Ɲq���?i���'�?�ţzY6����'-N1�t�ߛ��I矼�	g�)據6�`ur�/+Z~�u�b��#K���b�G����'�,�fN�'��	��M؂Wn@�s$&�Y�l0ٲ,�'WDY`@�ʙ�"�㇦x���Ñ@��i@�N'.V8*W�M�_M�9���ǃ8`�c#䈸Da�[Ŝ$pX�q�j��F�T$��`D=q�$���Ł�j݊t
j��gL�=AVt1���N�||����<q�,��Bf�(�6ʅ�a�0���I�c�H٢$��a�tx�ƎP���tX剌�>
H��̈�U��uCF�_�ਘ!"��U���OL�:�q2��o;���`�;6�k�P�@n��wh�|��F��{�1�W���G�n�p�m�8a�"AT�0M�e�1t�rq!_��۟�&�d�'����O�1�l������ �ĝ�CW�d����X��^y�$�^�� 9��E+ dV%L�"{^�[3�ئ���b�ayB�S��'�`4і+��QB��l��]��4�?�����D@�e1Je'>����?��V,��%y�9e돘Zr@Q�ƉJ��ē��D��H|��v �K��K��5 B���a�ZpnZDyB+�zz�7mg���'D�$�9?q��Նo�f���U?)d��PGߦ��'%��������8r����n��g��T��I�=t���N�4��7m�Ot���O<�	�z��Οx�c,�d׾��H!^��=��!�M�3G�s���2��@2c�#�a�#4��Ė3X��oZƟh����x�V$���'���O�q����$���eO�V4����,1O��OB���S���P(�Q��-��+�+wF`oZݟ$��O���'	"�'�i��AEA�"Zth�z0�H�⌵CV��>)-�O̓�?���?/O��3�#�B`�����d.��b�$�H�I��'�L�'��8�T"ޛc(��[�'J�4����'�b�'<�R�,z������,�qk�΢"��a�H	��$�O��)��<qeQ}"��;���EE���l�#�R?���O(��O�˓x��H����@�#�,����K�i�4��6�O��Or�@���>!%Śa��6�C�Q~>��w�צ���Пt�'�x��,��O��ɞ3c��k�*�?Z�6aa���%zj�&�h�'H ���T?�)A,�5�ȵR��H!H�fX�Mtӊ���E��i�D��?���]3�I��4�'�!.l�RR�B(��7��<�F�D���O���`��!q��CLy��5Z�46�Α��?���?a�'��|j�
�:Eq�؛��%p��Y2�����	�Z��"<�|r�cq�!�F��4�̔��݁�����i���'����(vn��G���'~�d�=G��h0�Kk��#�ʘ�#��$Dx��!�)�OX���O��&_q4K�:
�t
�
�զ���]0 x��ןи��6��9�_�vuҐJ��̮e�2��#�!W�ZQ%���8?����?���?a�Oژlh���	��d)T�X?x�T�ֆ��$�O�$�O^�O�����B��f�X��>���m�:0��%�����Od���O��:����43���AŘRTI[�aX-�t�!ҷi9�ҟ4$����ҟL	��Oӟ�}s �"��<�\Q0�&5�Xd�'&b�'k�R��x�����)�O�1��z� pB�d��U�};��@����L�����I�g����=q��	c�ډ;#�ɱS���)�����I��<�'����G�~Z��?a�'.$�p�@�h^Z�+0;j����x"�'w2%�'�O������Vn�+/�rT��G��2�7m�<�F��?ni�F�'�B�'x�DA�>�16r!x鎹Q��P�C	�b��n���	�
i��	J�IB�'pdd��1-{�Րq�W�w�<n�r��y!޴�?���?�'K��	oy2 S%M� ��ĭX?�d��'l�~�H7-�-aݲ� �b�x��@bc!�"&d�l��$�e&^�s�i:��'v�f˻w&�듦�d�O
�I�f����`�|�xQ!�F�c��i��O����O��D�':x*�!W)N�`�a�0�:�oǟd��������<������DP�X��D��U\�Av�q}��M�>�'�2�'W����b�;s�:i�3&�@�
�81�N�pl��(�O���?!H>1���?�V!h&q#�h~�t"t����<���?����dP$� �'2z��T#N�F�J@�WOE�]io\yB�'	�'pR�'��X��O����Y�@!�'�5.�.�J�Y��	՟��	Ry"	 ���'�?����{:,ƦҜ*iX0*@Q*I����'��'���'�z�A��B�b��i1����'_H,0���<����'��T���w�O���I�O��$��ʙ'G�xY£ٕ{�X�f�F�	���8f��?i�O�Dx��,F�r�@H7S0�(�ش���%C�n��l���0�3����f�4U��+Q鄿b�L��R�i���'Ǌ=0���$�3� ��:�aP%)L���把=p���C�i7����i���D�O����0�'剅��Q�㒦G��|r�n��f�zx۴Z��l����I�O�(p'I.i��I��ʥl��D9A���I��ҟ\�	�ayʡ	H<�'�?Y�'�q��
��1kv0�nƑ �l@��4�?�(O��w�D��'�2�'�ҩ�
T�ͫ`�߈E8*�B��*H��7��O̵��e�i>���t��=C���(t �
7	�5B1N<XN��On{�o�O��O�d�<!��5�8x�AF�,�������Żt���Yy��'��'S�O��D�OL���Î�x�0,0�WTX`�PV��
es�D�Ov˓�?�����$�O#E7dBӮY�J�acB�-�F6��O��(�	��I�<���jp�T�x�]1�a�A#�+׌e�&�x��'c�۟x�(�O���'j<����$�6$��A�"9���ib���t�I۟�[� �f�tO�I'B)$�����ю}V 0H��i��W���I�e����OGb?O�\c�ڤQ�폨D���X��)��-N<Q���?(�K�N �<�O�f�8���	I�.)����sYāPݴ��d�!1u��o�����O�I�y~�o_B��j���3��	����M�)O��c���O��&>1'?7�Y���NXhf��gM�=�Fh'?�26��O����O����F�i>�Ȃ��]"�C��J��Q�:�\o��$
Z��I0�'�Iy��':.Yu+!{����c����z���D�O���6LS,T'���T�f��D���X�k�f��F̿D�Ȁoҟ�'�>��~Γ�?!��?�Z_��q��IF�`&�T��V[����'�A��$�4���D%��))�ļy�@��_؀ �2l�5)����'C�����'N�'�R�,��-�x���mFtx�#V�lUz%"���Wyr�'����O��%k��1�3��L����,e��O��4�?����S�;$���'u�R�H.u�������'B��'�'C�� rᖼ���B�Yy+Ț?��!V,�7SJ9��O���O$��<Y֮�HǉOW^���H-�ˑG����-Q���'�'-剏o�T��j�)�bb�U!���e� �5�:eA���'*�\���vh���'�?A���pˏ�P��;���e�X�6.^Ŧ��'�'�&�8�'p��П��s�M�m�+_B"c�c^�G`�(#QnӺ�Ma�8B&�i�ꧡ?��'a�w@x��Q8�ܥ"�G��%�i�	�D֨Q�	2�ħ��禥����	�~U��GϷ5�h���j��I
&A殮�	������?)�M<ͧ' �%�SG�$lDl �ƀ<'��y��ia��F�'/�T��%?�۟����X� B"%�h�H0�ٓ�MK���?I��h��=;�x�O�B�O����OI6. P�CY�iw����i��V��:.چ������IS?AKI9��Q1g[`c^Q����a͓O�h�'�����'K�0�G(�2QBP���!®�˦��>Y\�1�!o~��'���'��	�U���(6�	E@dm���j�R̀E]3��d�<����D�O��d�OB)@�卶G��P��F�dl��$'�d�O@��O����O�ʓl��M��9��qB)���{��Z�o�t��'�iF���0�'G��'��H��yR�RQb��
�/٫f��4:aR�[Q�6m�O����OZ��<��33h�֟֘�[����΄:�M� �(1�6��O���?���?�V�<aH���^'D%D8&gS,p��*�Ki�D��O�ʓhDQ*4_?���ퟄ�Sx��:t T,|F��K�c�
���O`�d�OZ��A*B��Iny�ҟ�y:�,�����<wRzxr�i&�I%E��q�ڴ�?q���?i�'rR�i�}�E�T�� J@�84؈Q��pӢ���O�3�Ij�'5�X ����6(v��K�_N�mZ#5���4�?���?��'?���WyB�
?��e���(��&.J�3]�7��s���xyR���O��[F@�f��L��Z�f�)3��æ-��؟P�ɒ"<D�c�O���?��'�ڼTh�� <��C���`�\���<	C��<�Ov��'��)N"]���p��]��RIҡC���'抰k2$�>�(O��<������ �2���A�P�4kJ4OL}B����yr�'���'���'&�I'C��y��^N��]@���M��ЙڮO:ʓ�?�-O8���OP�D�F�ثw�W`P�h��d�� Hq(>O~�$�Ob�D�O��ķ<���&���z�
țq��8|ĬA �%^&l��_�d��|y��'2��')J�+�'��5	�H�rs Pwhֺ?� E�a�\�$�O��D�Oj˓}l\�{[?��� o���s��;��X�T&��hт��ߴ�?�*O�$�O�d@�d�d�O����Tn��`�7C��X�����En�4��Xy2dV�7x�'�?����B�c�|}q�LR�a�F�"&N�c���ß��П��+x��';Bܟ:�@�%��7�FСe�Z�
��ҷi��I*f�P�4�?	��?i�'v��i�)����y��p ��w, P�gj�~���O�!��:O��O�>:zT:�)P�'�&U ���U\6��f�nZ�@��<�����<qу)z,�\B�E�U�D�
�c˛v ��yҚ|r���O���f��	*E��b�I�7e~5������	���ɑw���;�O���?��'j��#$�J�y|�!��]=�$��4��-Ӥ8�S�d�'a��'�� ��
��Ŏ��m" �E��q���i��o�+M8D�����OVʓ�?�1-�&���͋>e�Y�l�-v	�U�'��(z�'���8���@�'D#��0B�6Y�"g ��f=�'�R0������OFʓ�?����?	եB�dv����W�_�fa���ET4��?����?����?�/Ohi���|2EG�T�ґ�҉�$f��Ȇ��M�I˟\$���	˟l��f]��萎�4V��0"r��6���IW���$�O��$�O��F=<�8���4�U�H�0���(��@��
W=��7-�OV�O���OvhhU6OP�'P�h��: M�(Z��&O����ٴ�?q����$�=���'>}�I�?�h��� ^�⨓�S�mG�����ٯ���?Y��/n��������suj���^��8�h����6�<yi��I�~R������� B��I0z� �2�ەJ5���ek�6��Oq;D9O��O �>��q
 ~���!*`��cB�t��$
������I؟ ���?O<)��1����@�d�DX�SOԊh�z�G�i	zXh��'|�'R������y��	�P���C-I|��Yn���	ܟ�`�؁��'Hb�Oԁe��:��8[Co�0t5F��вi��'3n�蜧���O�d�?Z�'>T$h������SJv�V���P��`'����ϟ�%��;�`1R��/3�)*�+z��4sv�̓���O����Olʓi>�Q�΅.}R�w!Ђf�:�a�	�O��d ���O���Ȭ<�Bu�GޮFi��ăݭ�`Ts��O���?1����'F9bm�f=�|�[3���	�D �_��йZ��xR�'8�'B�';�@A��'j&H�Șv��9b�
��7Ё2�F�>����?�����`��%>���O;rȻ�W6�@YV�\��M#�����?)�?)������Ɋt/�-�'^�N�����.�P7��O��Ĵ<id��c��O���O?�-��F�|'d ���΋7W�5��/��O����Z������
�1�Q�J�2sFC�`G��M�,O,��!��������*����'��}�`D5l
]�S(݂7{�X��4�?��q� J�����O��iVO��sΦmj� �)*��$�4T�\M�E�i�b�'���OF�O��$O3�,�w���XcP�Dpw��mZ& �d�	T�C���?�����'g.�y�B\M< 3�id��'���G�`�b�,��C?��ʌm�d*�Ŝr?���'�Ѧ�%��¡e�8��'�?���?9�Clʨ̩g�UHBD�f�� g2���'EzXi!e)�	ɟ%�֘� �4A1g�U�[�h�`����s?���|)�O>����?Q���DL(�hpР.���x�aA�`�����G�ß��Iw��ß��I!R��Ȋ�P�R}ȕN� d| V�h�̔'Q�'�"S�|X�eƽ����3�]Х���	P�K
����O�=�+Ol���j����E�;��'�^S@8��'+B�'��	֟�ie^�����L����qԄX�[db,4�aط�M�����?���	�Rt�Sz�ɃE���Q�,�76HK��_`��7�O����<�̌";i�O_"�O��\93�~5�%��A�s��ࢬ=���O6��d�%tX^�z�E�g�R��[ W.��^��s�T/�M��R?-���?i�OD��7�D �*HQ&D�
�n-���i���'G&DɊ�$9^���;F ɢ?�[�)U�T7MA���-m�Οh��䟈�� ���?�fǜ�@(�S!P)H����b��6ő��Oh�?1��
|[�Pq�y�� ^e���;�4�?	���?�Ck˿�?9����	�O��	�I,�8Wf)~""��ҫ�V�J=c�y�m1��<�d�O����g/hj@��$q"�8a�K�Z�FLm����	i�����T�D�'��>���S�U��d��/n̍YR�Q}R��$��'�R�'�r�'��i��I+�%8��"���K���̛�S�8�'���|�'���ߜR'&}zd�E52��$r��
$v�p�Ȇ�����O����O��t>�HÎ�?���L�M�z�0�阧_"`yI�DzӒ��O��D&�$�O����-�l���iJ�Lsu-��+<va&��9"�vDR�O��d�O���<QD�.X��O�\��`]��j2�'�"[^�b�Hn����O��|���)���^l`�Q,�l�T�Ø_�6M�O����OH��S�i����O��rbC
I<���cw�|
�T�A͉'��'Xz ��f�!����	�(ZAؕ�a�SL\Ф$�=��V[��h����M#\?���?QR�O�P��S�����d��OD��Ʊi+��'-bx[���钙n�P�I�x4�9�qc �1
��]�]ج6��Od��O2�	DU�؟�90�W�'Z*s �?�(�3�\�M�"g�T���:���;GJ�ɒ�����pm�-K[�QoZ�����ҟ��f���'�r�Of�4�F�jt�����Q��w����/|1O:���O@�dҀp�HjQ��
�I��@��eY�o�ڟA������?!����;��a-Ɛ��L/%Ȱ�`��s}BCЦ�'���'��]� !Gfh��QK�o��W]�$� �'��1��}��'��'���'�ZQC�ƝV� խX�tڱ�1��'�r�'�rU�� 7f���� Ē�C�Z�i�e�S�K�
��_�$�I��&� �	��h볍�>�Eʗ*8� +0J�"]Sj\�JT}��'�r�'��I$�F�@L|�%� ~�T yu�!T��[�k�/���'��'��'I`���}2��75J�ݛ���>�Z��T恉�M����?9,O\��C�FZ����35��t���D3�^��"��55K���N<1���?��"LA�'j�)�/!�D8��Ӭlj\X���v���i	�ɚ.�J۴�?��?�'&j�i� ��׾-��,�*�`i3G�z�p�$�O�HR61O�ʓ�?A����(0��i'΀%1�MJ J��M�0��3K���'���'���f�>�,O6�Ѳ�D�@��{�� ,��/�ܦ��G�O��$�<9����'�L��C�1<�JI1�hh����Gnl�����O�ĂF�8��'���ݟ<�KQ���*�& ��Z���_̐mZ~y��'v Yx�����O���O��q���&I �z�cQ�j�id��Ϧ=�	CVp�q�ONʓ�?+OL�������Z�8r��0�i��h�R�$���x�\��ޟ����\��uy��Êp(�}�)��'(�[%�V�>�4 ��>)O��d�<���?��$ ��"'����è�Q���re
��<i*O6�d�O
���<��(�.#��I �Q������d��m�4�ݔGA�vS����`yb�'p��'��P�'2��P����I�+��k/0e��Fe�0���O>���O�ʓ˖ �"R?��IP�"��M��P�pCD�~�Jٴ�?a)O����O,��u��Oh��0�&U+GǞ�3��xA̃6	7�On�D�<�E�O���SΟ����?͛�kŬ�޼���6'6f	�RȂ�����O��d�O�:!5O���<��O�5�d%�2v��|�q�&(�4��4���@ߨLmZ������+������ys뉩3���X��G�K3��0�inb�'{����'�'q�.ՠ�B�0tR�1���.T
��౳i�p{��n�
�d�Oz�������'���#�@���0��!��Jќh�شr�8�ϓ�?A(OV�?M�i�b�#!ʊYk��0\D�@요�M3���?I��`z\*O��'�?��'LVEYs�^�|�:!�'�\�+N2m�2�*�R��O���'�eMLx��)�aK!D(�Yw�J$/ 7-�O�!����E}B�~����?�H�h�C-��+�.��L��JSJm��.�$;���Ot��O��$}>�q�F�I����<c��*�� ����O���O
��=���O�ɮ9����JٵhCʽZ�����M��������X����ɫ1�h]��Zn|2�I�!u� [�f�!IO�@mZϟd�I���'�`�	���	��>�rM 
(�>�����K2x�13�My��">�)Y�a�FG@�F�d/�%7��!��/�l.aѳ����'F�UC��G�+�F��d�uɠdhS?��
�Sl8�0e��P�CH�z��ePA-�]p ��%f�"Sܔ	�Y�s�n��%E��|!��÷+��4�Woļ�EJ��}�x��%f�k�|����1�\�9gĪSvn=�w�ʪV{@18�����q��Z3KnnZ���9�JE����)xN��!P?y!ԑqP�-�<)R���O����O(4ˀM�Ypp����0�:x+��@';�FD�Ś�\�	 ,"~ڈ��O�1�w��?
fd
��	.�d2�aW{W�AQ0�˽0>������Uc ��(~�h��BF2|�Q��'Λ9�Iҗe�\������pⲕ�`�'k򒟒�6�Ob�Z�f� ygv��C�+.�d�k1"O��h ���JBc�Ԙ=���k��ɯ�HO��}��ix�+�&.)Z���O�a� ��ȟ�2��Z/Y����ٟ��I��\wPb�'�ȥyJ�
j$�, ��Lb��'R��j�����i�E3O���p�Ek�� Kam-rL-��O:�
���{L��r��\8�8��Vk8):ҥ��4ap촟D;���O��$/ړ����F��,r!����%"-]�z�!�X,[�(��Є\J�(5K �م2�v8Ezʟ�˓��u2�i�h�{ �N?�Q��n��k�Ea��'�B�'���	*���'�iV�Q@cM��#����n��&l��j�_h��D蓐\�����eX<�.��x�pu�J�R��X��,U�^r�%�R	Ɠcib��ĕ�^Rr�'wlx��Y:B�9��� lRbx�b�IQ�'�x�CU�rj
I�Ѯگd��\�'�B5��.ٹ7�����&��3�'lꓴ���7�$��'#]>1K��~F�1s�l՘tN�;&-�V���	�����K�zu�يMf��Z��'dGb/H����:4jI��gY&�(O6ك
ŷ_��� �HܧZ���Vρ�>0|�i]�D^�Gy2��9�?	����O���#��͍w��L��;Ҝd	�'9��A"S0@�r#�׏T� 9 aÌ�0>Y�x2,]���G����8�o��yIIz0�6��<a/�����O��d�O�(Q�[{��Ua#+�T���zdL�"]r��>�|Fx�%"+����J�h�(�+�� ^|����)�矨���Z%1�1
�5 �,���
����u��f�S��?Q"�*s:�����b<����@�C�<a�M�j�J ��:d�Y�D�|�'Bj#=�π n���n��Qjǝ�:��S���OX�$U	kT����Oz���Or�D��s�Ӽ�7�K=�|hP��]�Њ$˔b?aŎSx�ܰ�ȓa7�ź�� �pL�`����«:�Ov�i�#� �H���R1�4� �O�0��'�{���t���Pӄ���e���˙�y��X��0�����h3�擁C'v"=E�ĢR܊6O�q�"�C���7E��+QB��2���d�O����Od`�D(�O��a>�Re�{�.,v)�.!d�;q��-w(ܜA���,�(A���"##Xe���Ƒ6����օ�v�)Պ��a٦aÇ�Y�!Y6/څi����J�'9z�����?ich�k�&`�1�Ƃ�bQ�U���hO*�? �ߊ�buX0q�E&��DN!�d�,����`E��v���p"/�zL�$a}bR�l�FiS��M��?�+�HAℋT"oð������ �R�L5�^�D�O��d�#� ��5�|��
˷6,A2��SD�<�@��f�'C�ٛ�����\�Ղ�AYHer�l��"�Q�db(�O̢}��ʞ,FT�C�K(
%� gFEX�<)�+Г~�p�hWK�%@�}iV'RW��!I<Y@��3 N�pvaP�Ur�� wLM�<�"[e���'��S>9�_���'k�I�b%� ��剽7���[T �
+�J�'^1O�3h���� �
��82&b
�
���vJ
�O?�䜷$r��X�/}4X����Z%�ek��O�c�"~�ɾ&��p cY�<f
@�U�]l*2B�0c�ucC�11���� �[x]B#<Q��)�I�0j��J��\�Y�5eK!�?Y��x�X��3f�5�?I���?	��^����O�.�:=3��̙�K�E��ִK��D�R��}���#" �2��Cn,�k7(]��~r���>�G���I�
��V�U/p�Pրh?HG���>.�Ph��ґB�fQ,�:�B�	�[hd��ÁC��4�2 a	9aR�������ͦ���G�k�6��q+M�Q��A���ڟ\����	$} ��Iǟ�'r�p��I؟���Q�a@D��.{�E�%�O4PTS�H1ы�/b��t��͟,���f$.�O�RP�'DR�?$۸5�$�W;<غ�K�aG!�y�+N&Q�vxR6G�o@i�ǂU+�ybH�1+�x|P�A��{�<8�m�.�y�f8�I�lI���4�?)����ɑ�	��	Y"��z�bx��$��"�+�OF�$�O����1b�<��p�Y.O�~�)t��|2�@,C����f��]d�B�I�T�'˜� e�7p�\!�5�O�j��*�\�K�e_�K8l�����5K��I��	�Q���ɦ��I��t�O��H���N�XT�vM@�A�y#��';��'�������'f�AR�,͛r���Ѯ�'_����dIq�I2_���%��C������&y�n�Ʌ� �8�4�?����D�!}F���OR�d�����H�$S)xQz�E�7J���b-�O0�O��g�'��
���=172XZ��+,�d�iź�e"p!�<�maէ���ED�E�)@0�t�x��NG3w_BY��'�"��<��P��?�U�P�L�� HĢ��lmi�Q�<�����>qD+�,W ���Ǎ9��i�$}QZ�d<�I��M����h��P�D�'Bz}��cS�H�B	J!�)4�dڅF,Ǣ˂��eіm�'%+D���M�N�Ā��=}b�S�6D�d���g�l �!Ǆ!� ����1D����ȶP�V8�Ѣ�3��<��b$D�[�2D���vH��VDܘˑ%#D��X#�y!�5g�N�D�@<D�`��h�(��(�Z�Ir\��n8D���W�@*| �	�!˥b �2i6D�HP��4K�E�3釀��*��&D�����Vo�$S�D�71@�f%D���ʖ!��0if�"��9F-(D��3�M����L��
X�c�N%D�,R���T�FtH���L���$>D�����1�@��OB*O���2D� �#�ݥm^�t�Т���l�`A.D��J����V\��	�/�JâLj�.D���%���CC4EӔ#J���8Q(,D�� �X�!	�r1���Ԭt���"O�T��hq5���Ä]@Z���"O�iC`�7�y��C�d��x�"O�
U�̒bh2�9��v�i�d"O�a�����Eh�nܘ\d�ap�"O�P�@ƥ)S��QD	5<L:u"Ov!�¦�UT��)���|(ڵ�%"O���mR�w]Ԝ����q=b<�F"Ov�K���F����Ŝ�7@��!"O�����O�q�W�V%B�"O���pN$ ��<Q��y�N�S�"O�)�cûL1��Ӌի,��K�"O�93`bԆ 3F\ɥ�Xk�@H�"O>%3gT�|�X9vM\�r�@<ڳ"O�<�%c�	�:P�hP��"O��Iq�T Zx�qc�e��TC"Or�:a$߱j��bϑS�b�v"O�I�uK�<8��`��\;*�#�'Z�1B�O۬_����čn��h���J�!���r�Oɳ�x��aN<ݚ�k%��ɁJ#��O*���̈�_{l�@!�L���ⱦ�+@2�HqU%#T!�$
8-�jI��!ܺa%F�R�M/�󤗶^ҍ[�b(1��)�uܮɀ��{�����@7Y��P�ȓqpSP΂YxR��� ��#��'��� �� (uO,0��%
B�"�-�Q�&�wĆ8/H�8��� ]�������ƝY���P��L#|�T8*�K!�Hx�O��i��%�W+*���Ŧ%��)���T�`�zE�|r�g�\��{�#Ƙ*ԝR��l�<���1&��B�G�
���t���<!2++`t�0���~~���NW���2��*3d���f�!��Q"G�x̨%��/y��mѤ�>w�I	[���"I>0u���D�;F7��1�`4��'}ya~Ⓖ8:��!Q�S�H]����7�-�e�֔f* ux�'�|92sg)� ls�n݉`�|����$�-Cn��b��iF1�J�bD@�c&4H���(B�f�1�"O�Փ�'��%9 Y�Do�NǲYb�;O��J�6]����"~rѫ�
tx�0�J�E��Uy#��l�<�rmܶ5fѳb�4��4��Ŝg~���%`��)�/�;�0<	�!\&^ZX��Pf�T\��8��W�<Q���8R��9
�27�� C�H�<q�@�lO���GPȽ����X�<�0(�L�
	Ď?��5�U�<�a�Hf�Kg,�~�	�ՅV�<�c���UCRtÖ��x� qRǪ
V�<٤ȁ�9!"ٰD]�,� yP ;D��E��P�c�� ��Ģ&D����R͜�� N��0r�$ b�8D�p��C@�!pv��U	6WZz�Y5�7D��'�V�
<���jȪG�dh#'�9D���o@.!G^Ԛ���&ˎ�� !9D�Y��h1Zy�`�ə6�xu2D�\Q2��+M4��{��ū�Zea�).D���ւH>=�����G��#R�*D�<�pmMB��c���=4q����"D�����[�x��L�#�b�Ю4D����
�^���ȃPQH�K#D(D��Bq��*K�$�s�ɐS�VM�B&D���!(F�9������QDq ��)D����*8{s"T���:3��Y�"D���"L�"���#��rEе9Eh?D��A���1~�
H���X���5J��;D�Lʒo�0�8��v!����[�%5D� �w�Äi^%R�aE��4�%�4D��A�Z�rT"��]�Y[����2D�� �01D��C0]h�E�J�;�'��!AG0}�D�]��[҆�:.i����߮�y��nH�	sDn@�{�tI��h���'��`"���r>�3���*���򩗷(�����>�g�ߒ���H� �J"ќgH�����,s_��ca�p)qO��p��Y���D`�"2���4��Stl�#&�dE3Ͷ��Ǆ�h���''���y�gP(/pl�!̀�ݰ=	a��i��@���߳n�`H� �)t�y�gL$��O��á%�m���>�~���j��B�>I�l$h&@��Or��N�sB�)ы�T)�=gmP)��ɭ.���R%ޭ��_UZ�Yf�J�_�:e�g�S�f,�}�CE=�J�Q񠙰R˴�k�j�Q��e�e�\5O�)�D;��D<U��w3�� J��%.�Q bDW�Uq�[v�����h ��+���f�R���3��з	���ۄ�̖kVv����|��dB�-hHm�`i�H�'LԸ0Dkȡ|�6)ju동V���b�G��6m�$A�~�qK<Yv φ	J���.Q�)l�[���AO|��M���Q�&��#	���0�0\]Q� �UE��
� qӦ��!���S�?��y�aڎhS)+��T*[���#^�D��@I)<%R�($L>1�=��a^�ML��Q���iɶjha{�k�@8��7�_��~�ڑ[K�$��(�M���4dZw�O��hsro�-�Jl�2Z�)iB� �G7ց���݄# U��"ı�ħm��A�2-�<��IޡHF[פɴ��zvJ�?��=ʔa��uE�l�7 ̬c�����m��a�sHYA5(�k�\(���(9�DA�bv��n�JA2�0�H0��)��+��M(����ـ����T��Y�G�$	v%:��É'��Hp�OXI�D�5�4mA�ˈ$����K�	^�� c�Y38��#�O�����`P�m��o�R���OA��$�R�r�kR�i�9�OD���o�6�M�`�9�E�qdD6�YY��"v"��rK_	Ph\Jwڇ�b�I�_�Z����S�?�.�P�k9U?�:W�T(PWH0�I�	U[���Q���3�N� q�L0s��	�J��OD�R��Xky��2-�1��h�?�f��AA�8�@<aS��M�g�Ю� H����O��˂�9_��%�G�/S������QѬ0���A��~��6��~�����O,�a'��$f�Ȥ@v���X��O4��&p�		44��.�K��Y���"l��7��NlU�!ʁ�e��9�g�s(�q:��&O\�@�8�Q��+gᨤH�(T����$/1rf� �OF�0��G9h��7��J	pUP X����đ�CC��RUΒ�G~T����!;:a�u$��4�<8Z��i�	U�#E#A�m|E!��K���U�P���'��Y�L|���A4x��1w,�AZG�АN����AZ�i�F<3G�ql-��N��l���6���a�gͬFutd�ل*���ʥ�	�w��Ѡ���0I����ꞁ{��'�z�	3(&_,��Z2J��s��4��A�5�.Z���O��[��A�p�@�%�8ل�;P�i�����K���[���2]@!��mX��7I�m��V	_��I�cBn�ˋ�Mi+�	����K���f�$ZJ�j�#)�L	�째ϭ�E3O",�Sw+��PzhɁ�{��U*9��`�֪�
)�YF�� X�Dx�B)���@qm��an
����P�7���I-TW��J|&M�|�	����;�*�`P�W�}�J�*- ��'�Z��`��X�R�P*!F���u�N����l*Hv�f�*����DR�AJ�0b��ǳKd�hB` ?X6�O,��ʂ1`ģד�i@,O��x����e^�j�v]K�oC!�$�� �x�e�5k ��i�KT��2��v�Y��Z�F:D�)ʧ?���԰3���e�ƈV"Dd!��0���:3�E�c@9�f�Ίr��Qn�<�V��O�����ͺ��O���ēP�䛤#��4��9I���M�h���c!�tZ%i|�����@0+
�б�nŧ	댠14��:5P��H=m��8K����ɩ_+�L� OD�Oa  ��a�� 
v�ޒ<�^�Xel�%8�R}Gp����Ӊ���� �pdD�� %,5���d�� B�ɆpHB8��B��5����w��LJ,��>�(��J�]m�L1W���?9[a�����43��0$�  �a�9�Y�&�<KFxC�I	"FxQ��.[&+ņJ<O�R�Ѡb�1� �B1e��Vd��� #U;M�VY��P�&)��:?I3�I?4�T�K���)^2T�!��e������6k�:�t�B�a�������k垸�`!��c���BЋZ�زR���yr�L�{�����Z�lЩ�`Q�)=�,��$�1O��a, �K������
���֫ؒ����	��	~���EZ�g�f-�R��.��8q�F-Q!�$�"o�>4`A̡azt�hb��{"��R3A���O��f��11'�/>���t矩�y�*O9�TI��J?;�|�'y�L��f�q�c�6k�"�o�8)Y*2X�AP�X�q��2`��  D�Z��*?qS%�? L�6�d�����-
r؞X� �R���EC�Z�E�d�*��"��t����]+���f�[\!*Ɔ]�|��۱
H�(�џ,�tD�!����E^��|�R�(�c��sn�=lr�%��S�2�El��Bi����|�~E[+đ�-8�%�v��� ����HZ5F�
�8ǪҥB�@����:��UcP��3,*\(���{	����@JUy�O��$λ����a�,�bqīM bo�%��P��82D�*��e��B: Q��g˴\�U�p�tT+$�,�v��7��xy⎠<i��3�$���/գ(gTT��l�_���u(�ݶ[���>��y1�LR�e�N!�w%Y�y@��[%��7M$TY��"8ג���Y��ʢ?Y�g��v�	G�X�+�d��5��\ܓS�X�Z�M� 9��l���XZE�\{!�D�QU�-�ߴ(�}�"��{�1�X'J4K[4OC>|����X��ԉ�ڥhy*q���Шb��h�ՋI�ll�\����
�h򃝔5�Ջ*O��/�y�	��FPz�X��)>������$�y�e��i��0Y���o`b��u%=ۆ�ٲ�!��ʓ8��m&n�:8D�šG���f\�'(<U���F�Z�aB�ɠ�H���I"̊,J1��-�<T���C�f�h52�g\)U�$kU:&>kb�F#��q*A%2V�a��	�*x�Є'Ρ;n@C��]I^�?��J�x�	�%�F�v${���*^UvHC!M�jS�ȁ����P�Wm��xr���O����-ƶl�"՚�	�HO��;����h�-��	��A�LŉsJt�d"O$�£I(�AWm�s;��S��'��U������I�c��?N{�y�@K�4vx(�ȓ}�B��G�ȃ=p>���F�5RF~u��>��lQ�m�w� �#��'s@�ȓtff��qe.�� �'$֤.Vb,��'� �A��uwl0J4�rm��ȓL��	@�Շ/�8l�ևԇ,��q��_
��l��L�A��.xܵ��|gD��r�M�7�i�q�*-Ą��	��`�BK�<�J�F�8Fzy��T�����OL?��<���B'2\���q|Q�`�:Q�0��2aQ�Hx�5�ȓB��msQ��..洩��H/�ل�VP|�֫en�8�i�;k):Ąȓq��y� �6C�@���D�1��A��D�Pq�#�A��*M9%R��3��VhX	���봪�0"�ȓ�.�b��2��p{"
�'*�n��ȓJ�`����q�-�_��ȶ��P�1;���d)Οn�|x�ȓ!�P<3C�O0El,[i�; zA�ȓ�Z�s�����%K��7:����ȓdR`PIu O��=�b]�+�x}�ȓ(��	16+�5$��0�b#�7~>�Ņ�kW�Й�!��h����mǵ_� �ȓt�F)C##��@i[D��d	�0�ȓ��]ӑ�Z�u��2@˩�����&���z�AD�)p���X�q�@��ȓ-��ǘ@��u�7�O$�.هȓ("���%���U�L�56�E"O��I���C�.d���s$��A�"O�$�<V��
R���L@>]C�"O�E��i '	BU�� ��CA"O���p�|�kF�0V0��J1"O~�3pI��t��B��Ͷ��Mx�"O�d�GM��H���:���Uf��"Ov)�M^�����3^$j;�i��"OLT+m31%l|j���9��"O���dϙ6F䀴�;&tr�"O��θ/��,B䡟� 4�C�"O�0��QU��"��70�� "O������,� 'O
�p��)#�"O*p���IS� q,:{�F�`@"O2Y�@��=N@�0�)�Z{����"O(Y���R=6h�� �鍇nt���W"O��L݋lL�@Pg�Ǻn`Y�"O��R��7��hr�UPb ��"O�4����6,^VH��BՂ+��-��"O� ֝@3�J
K�D�3��y6A�"O�D=T�����F�v:h��a"ONA[%K.f�T� N��X����"O
�V�5\��u����=pwr�h�"O����]$i�%P��U
T��%"Ox9
���
�`x
�T����"OЄ�7gQ����Q�.�� P�i��"O
�W�^P� �k�.��<B"O�U:�#S���fM�-@<p%��"O(���H8)[�ha�+T(a�"O�e��U�j'�H�U��� "O|�3ak�:������9�7"Oh�QBD7�DY4���:�h��'"O��Rv�ä�<����4^�B�s6"OK� D�<���)U=)kƄ���y�eO<x����A Q�<��\�u��yB���M�v�+D�)A+�+�y�C��R�=�b	^1Bl�9f��y"Ζ->�U�� JL��U��Eլ�y"@ߖHv	��M	��&(��$F��y�`�2Z�ZU�q"N>Y,�6n�c`!��Z��uӲ���(>1���B:�!�*Sz���6GK��0 �S.K�!�#R;�`� ��:��(Z�7�!�(F��)�a$U�Y�i�@gB�'�!򄌤2r"�G=D����%�<F!�$�O��r3��(-�,P
��[3	!�?��RT�̽8�"Pь��{�!�>V(�(���?����A� �!�ҝt
R�c���e�m���	!��a�^9�q�N�0��H�s�^1!�DFY�.��V" �.�Nk�a��_!��T��`��F��Nb�m����I)!�N�6� ��C�q|�˰/�m!��]�<���ɗ3d�u�6�߼gD!�dW6�4d�Cf�%���M7�!�ĉy��L��AN� j��x!�U�{w!�Ǌ��b���r[��lU)#!��Q�Oq��1��>W,]9�mӔ!�J.f���$"@��݌{!�d�%l~��ti��v��Łp��O!��)
ê� B�5*VT�Y����"O�-k��S���%ݬ;�F���"O*7�5O��I��H��"Z'"O�q(Y�5�y��EY��)�"OĤ�l��3�肤�] B|�"OԸz�(426XYg�U,��%"O<PQ�͔-z�Ȳ(1V�><��"OH����<]+�)�P)�v�x�XP"O���鐑W��q�(� 4����"O`d��
�Q�����;:T�"O��#�BŎTCι���S�Z��"OT@u��:.7���,ŖD_�"O��;#�/4z�J��G4FU�"O`�ҳ��#;��x��ퟦ8���P"O��B��RB��l��P�t��w"O����es���0LʶRvP�"O2)k%@�G�=*�>\�F"OP%a��.� y�p&̮�\(8D"O&�R��]?�* ����$$b���a"O\U��hV�YL��.�US
m�a"O��J�"P%\�(]���W;~'0T�'"O���a�92�|)Y��
�3-ƽ�"Oj�ᷠ�%?�����H�1o<�Y�"O� dYP b�+V禨"2g�+4�t��"O6ʷ�͚m�r�x񫖖LI6�є�'y�I�$����G��<e��I�Q)�B�	9a��EC�`�<njp����B�,]ŉ���DX2��������,�	DÀP"���8�4N�,!�B�I.+n�)6��J�`�rs�G�K?j�d�ǣ�{�S�S�O_�3 H˛H�2@�'  ��C䉯~�TH�s��y�"�&@(WH�!C��d�{���$&}$��[�	ݩ< �b��I�!�d�=	_�LQ��A�l����K�;j!�d��m��ā%IǊE�v��B�N�!�D�5�pd�� /�T����!�D��jMЦ�ˬ7-N����
�!��D�r��H��A�lɾ�3g/I�!��ͨf����I݇��`� �X!�d�4f�@͚W㈟T����$�P8%I!�Ӱ/z�%*qgT!q�0��ҪJ1�!�d�5�����g���Q�V��!�$���4	$�Оi�j�'ϼ?�!�Z1	?\E���F ����Y7ޡ�Dw�Z|�E�6�ft�P�y�|4��"O�H�1��N�-��İX$�e8�"O�0""L�<���0��?S$�Q2"O�%��d�(�!@�~^
� r"Oԁf�˥LR.�C���SB~ij�"Ox���4W��22A�55�lKu�G^������]�A�IyҢ�0s��6���y�2 �����*U�<r�F��y��ԮE�|U���H,A� B`U8�yRn�%��a�9�^���Î��y2A;dd<� C	j�u΃>�ybd�i��)'&��Umf�ID�G��yr	�)Xr$����Rm�4)am��y�Jn�H�唠N��ь�y��B�/}�b���Fٸ�9����yBaVb�i	E@)zX�B	6�y��C�P�v`o�0Ou4���]�y",�J�0�(W�xd!Eƽ�y�Z�G��`��]6J�z�Ak�4�y��R�d�����Y���G��yr��Y�f����_�Z�XP��?�y"`ͫ�6�1%,]�IҢ�'�yb�WeZe
�m�5M9���dJ�yrh' f����)G"L@!��yB�=�09R���iO�=�`�ߓ�y�&�=<�n����g��U���O+�yR�P�(����S�F�Xi�`!�[�y]3*�a6��P��`7G�&�y��[�5c��ځ*F����M3�y������
�>o쀺���7�y2�B&O�AQ5�^�2[���Q�y�%A�H�2�hAA�)<G����,�yR	@�(ѐO��=ڲP�v�4�y�ߩx����D"0_��i6b���hO���G9ON��cW:$��JC�>�!�d^�ZI�tr��U�@�W�!�d >"�[�h lrE�D�E�R�!�d�'5�@  e��	���g�� 1!��K�xi�!�Y�o� =R�.q3!�D�*Z�"��2�V�bĭ�9A2!�D�r��ċG�Ͳ!K^��-	<~�!��!KH�a�K�}�~d��F��!�]NLl`�I_1e�����ĕv�!�� ���/��1j޴ ��W�H�5	1"O�Pa�m�*�AY�!T�/��u˒"O�2�V�BqR�!"b �)ڶ@�%"Ot�A�d�8��u��5?7ֱ�R"O�!�I\(=�>�� o=3� j0"O�#�
WH��	�E�6H��!!"O$D�d�жW��cd½m�Z8{VZ�HG{��)Z� �A�
C U���˪�!�DG� �=��A^�y-^@HbӘ]g!���oB;�`ڈx(%vE3
@!�D� #��5�ŒD�uz�� �8!��&zɎb��+��YB"�- !�D˜i[\IƉ��"Ju� �!���y<N����b��ʓ�0|�!�dK�g����#C	7�$�Z�f��h!�D�$jcF���o��Dц�A��^�"�!�D�,Z�y��ԩsb=	vl�!�DO'[	Ш��e�oaBвL|7!���!�P��,i\�|r�Il!�D�)ߴ�2�j��5|��[#8!�$~�L��E!� [�,� $k$G%!��T2 ��䱴ԙW<�|���O)!�d�-T�0�H���C�@�F!�d�
X��h�b�ݓ��@��oK;
!�d4'��-(ۉl�q�@�#�!�D��Lw8�ei^&5$.�xf@^"7�!��Ց*X�ȚR��aFe�ρj�!�ĉ&���P0�0��E��e��!�DN�G�R�Je�,j�F��FJ@�5�!�s�bt:�|���
<�!�d��pp*��2��q���`���!�DV�!���R�G�(�Wm�T�!�$ǌY��T)�J��lsb,P3	�!�d?/�f�Յ٬d!� ��!���16!"!�e݂k�<"�I�`!�Ȝ�"��+��*h���@Ok�!�d�.%�tI�(�?E��#G�X�D�!�q�p�8T�̡M�~܂��Ҳ-�!�dȫh�6��3�5�Ɛ��A��!�d#�V Q���"�дJ2� =�!�d{�<H �']Lg��u���6!�d��|�ع���:�2I��*u2!�Dۂs��kS�Ҩ5V���g�6E!���k<�\�$�Ԑe�-ꗦ	�]!���d����e{�50gT!�$H�)r<�2#n��La��I{�!�䞂=�f���EE�u�euOB@!�DO4��H��&��XgVQ���u�!�$T6]�6 ���-O���v���!���_|�Ѭ�7-7�-R�*��p�!��)tj����ɵj��Q���P8w�!��S5ܱ7��0�ab7�2Q�!��O�"�ȳ2 \=^��ĥ]�\h!�D� m&b�;b�J������"3!�p����$��-$�,,��C
>�!���9�*铃�.�
X�#"�*	�!��\6*\��Fr��� �a�.L�!���M���bk�0{�u�s�&�!�d���Z����٢d�$Xu��-�!���T�
q;�F�Up��Ya����'}�l�ԩ�k�D�0	�<#��'���BNX`D�h������q�
�'�4u2�*Ћ*Z�}�����D��'<)�7��&:��5�T������ ^��e�W*(L��Cq�_+��"O�̩w��ŠMHD��n��"O0�eㅦ5-n�@��_)l��-��"O�9�����t��b�j����"O�9��E͢<���r�6[ ���"O�!�f�ߗv�n���%�2l�"O��� ���}��L	1�K�����"Oz1:����N�Tŝ8Rv�ŋ"O�u٥�C<U
`�A���:jr١"O����@?,�
� ��;`���""O�`9�B%k�� G �?/���W"O��'�6mcH��d��{�Ш�"OJP�`l�a6���|c��Bq"O�]0E��b���p��ի>32ђ�"O|ڗ�S�;��Q�7>S�x�"O^a�ʓ&�B]��E2a `���"O��(�)щ[���СO�	�� �"OZ�k�燏eg.����)�za#a"O�=���C�p���-��j�x�"O��hɧ_�䘕RgR}j�"Onɓ�h_�O���`���`��"O�<B!�6>�\ف��&P�"O��x�ᗪIv�J4�A�}�0(�"OXX�.Q
 ^�H���t��6"Ob���0 }�� ��4�J¦"O��C�XN�]�C&�?n޶��q"O��xGL��z���+dܢ��""O����L]�/tQX�;VӀ�%"OL��"�n�=���k��}A�"OI�#HүO��!#���
���b�"O\1�DiA�F�&y �b�Y�Hu@"O�u��A�h}X����	&����"O���P�CNjab�]��sS"O� �r�P�}L��`Q��0�`�"O(l�rD�)y�h��.�j<ȅ��"O���	!}8A��Mۋ�0��&"Od�!�|��I[c�[�h���r"O���ӭ�+�����X#V�4�!e"O��"�dF'�<q�0`����,@�"O(��dQ�t!��;u��5u��5�p"O�m��MK�eJ���,V�}�x@"O���G��d��vk^��i)�"OXyZ�DW�t��Ck�+)�V���"OV��ĀIt�tІ�mΑX�"O %�U��
�A�Vm��TW<�i�"OdDA�C?3��Q��;cl��"O�0���C�9n:��#-�F,�Y�"O�QC7�F���%E����B"O"U�$&�8A�: ���?t6�(K"O�x�v,Ә:�=��C�,4$�ab"O�$q��ٟC�H����'/	�"OКU�I�:e�Y&l���\�"O��
ê��
J� �\b�"O�y�"��;Ԃ5�u��4H�^4m,D��a��Ҝ-�(G�K+
\I�#'D���&F�E��j�(ʑMx�P�,%T������-�x� e��TǶ�K�"O����P��I ���}�L\�2"Op�r��L�nv,B2䃚� )s3"O>�"��T��5q�#J��A�"O. � ��F�P,����4��� �"O�=������0�d���0)P"Ox�(��X�OL��c&Z�'�V���"Od`�� �.���Q���e\��IF"O� �� .�J����5��wh��P"OB��`L)b�V� |�Q�"O�M�W��6�[SFY1g|��"OLP1�܉J�VXq�  _7ZP:T"O��Ӡ�:3?�	�T$�,k�Ф0C"O�ĘW�D�.�`A���y�J�[p"O蝠��ҧZ1�] �K,��H��"O֬Y���#nZ�d�ц\'[�(��"O�hY1�2����OG HRB"OT�[�glhL8!n�LŁd"O�U;T��"!��Ix���ml�Bg"O~]1ҮK�TH$�
s�Ŗj\�)�"O��s��)h ��$�>P#�	y"OĹa��Q#e��cI�Ih�"OxfM��r��Q��AG�W�8�"O���cf-�&	���3fSZ)C*O�����Z�q���e`�1�\�h�'����c��{�@i ��']bT��',���T��6402�-��	�6���'U�壅^�q�|��Ga4]<y�'�|Mx��w
R@���<E���'�p�Za)�rs����CE,)���'�f�V1�vyR�@C!g��(�'C����ɤY{`�32���x��'��yʦ�!T���;���wE�t�'�D�r�CN/�=Q���nH�M��'���;�M@��������WP�<qg�N�!�Pa��+V\\j�+��K�<���I�>��;�푽MI$��EX`�<��痡P���0���V���a&�V�<����tT��d�!{�Y��#S�<���ڌg�4�T�ޖU6��`��j�<ɔ���P&�Xb�0�g g�<	G��p�`J�Ŝ�qt�9�-�e�<YWҿx�&͙��5 Ѣ�3�"�g�<)Ǌ��+����
z<bZq��w�<��O�yn�qivk�-,"����ENr�<y�&���v�a�U �<�c�kFU�<)$`��}���AO�f�̃�LQ�<�S�1e��'FȋEl���L�S�<��$uѲp�s�E=;B�����P�<��ބ!��KT"��xH�8�q�KS�<צքL� ��� ^9x�乚��L�<�i���({�`7�΁zЂ�G�<ْI@-~t5��.�mf@!Z���E�<��.V5o\H	�`�/G���*��z�<��jD0vR�h�3��0�D�gÛs�<	�a�.#pp����C�F����K�m�<ɇ�E�q=���VEW8d���j���hO�0/�K5�4�Z[�e
 bՄȓF
L���Sf�52R��	@r�&����%L�����([�P����d�RC�	�	�� 8󏐡T�f%¥��MTB�	04��3p�ӮG:5i�B]4h|C�ɧA�M���R�FiZ�S�c_i�zC�n8D|��Y�d�Cu��L	RC�	�~]"t)7�55y.����֌KU����.�u>RH��B[7pK�Jt�](8�`�ȓe0��%�:.N�Y�ɟ%.�,��ȓ�z!X�-�O��%�-@&aOn0��+A�qZ���&�,"��ٖ-������'�<��s��11���p#C_��b@��'���A ��C(9)C�>4/ �
�'�����E�1h��{��= ߓ���� XJ�D�'Ӧ�q����J���"O�2�D�c�Z9i׀�	p�6)[�"O$�a��۴�b�i�BU�{ź�3P"O�� iJ-m��a�~P����'W�ə4���4J^�(H�c��1Z� B�I6]�&��d���R�s��0��B䉱Sḽفb��f�9�昏p��B�I�"
�#�	<ju\4��X ~�B�ɼk����"�X�f?P�+D���X �B�	t�4���U	l��a��e�#)LB�*E�t[�})�B זc+�<�""O�e�󇍮P��mWLX�2����O����L�]ȬS��8�X�I��Ƴ:�!�	Xh�H��̜4��H3�	��z�!�DD�m�VA�5��8ߔ�"�fg!�d�l)�}2�MI��<��OģO�!�$�i0��%i6bйΝ#%�!�5.�Ue�8R���&m�Q�!�D�?3�����$m��}�!�V"Q�'��Y��j��#E�!���5`J�A毙�>�z�H�m��n��`�a���8�S �U3)ݜ��3�'D��&&P��zA֨W+ItU���&D���cbS*B�@��AC�S���4$7D�$��
��8Y����<(f�3D��A�,kI���=M�q�v�˦d�!�d��ֱ2k�s�	�B8L�!�d��nIɡHW��8c� �/��O�Xҗ&�Q�6� �_�k�iQZ�̆���h7*��'dR$[P�x�d!<~�C�ɍ"ߞt[A��2$q�t�j�|E�B�ɯ8����PK��,j�� 3D*]G�B䉯=��w��!S�UH��Оr�dB����,Xh:T�ٿR���@�<a����q6�u[��beVMyL˛~�~��0?1Ô�`�|�c%�:"��P��]J��0=��(B�t�H<2b�:p��-�#A}�<��%X� `��=27P���C{�<	���#�~���� ;*X����b�<!T�H�{@�ŦP�ऊLU�<��$49o�2v*٣+FD�*WER�<a�jۦh�`�+�NU�5b�g�K�<���PI7b�IV힒gB�cU��G��0=�q�݄"�����%J�𑢤�F�<٢&Z���,�s�R[T�adEB�<D�΁ 1R�bJ
�+�~��7-[z�<��@��Ȍ����lP�8)���v����<!"ズ/q�%�]��9�!�IH�<!EQ�W�dYz���!��KC�<!�KC15�}�G�E��oF���0=�ť��^�|���
�L��Q�A�<Ac�^	7�|S���;KR����Q�<d##6�j���
�!'������WM�<Y���
WlH(	�N�8l0�
+T�<���&(5�ړH<�ѳ�S�<��*վ2��JC�[�N������QX�<�E�Vߒ�qēe%XL[���J�'M��Y�']z|Qq��g�e�#�<a���
�'K�P�1k���u�DH�V�\��	�'c�p2Q�c��BB�VH�⼉	�'��YU�Br��u�qH �i�����'�P)��G�c�01�\�i<���'�L��s��jo���1��[��-��'������D
����®S�ʥ�(O��=��� �`����+#�&��R��	�h,�@"O�zu��:O'��H�+ڷo���"`"O�y0LU5�4XR�Ȇ���p�4"O�j bC�-�PL���Ŵ0�1yg"O�-HW���Vt��%b[�,�\�"O�]: OW���<�P��,����$"O|�Y��_>̂�#���s�¥`"O��[q�m!�W'�"@X�"O&�y��#\���0���)h�y�"O,� �ʋ�CaXQ�Mً\
�kg�D+LO85�,��F(p�,U�K<���"O�9�҄��@�}�j\���bE"O����U7G���d��#|l��"O�"�ߴ	&�"�!��$K~�:�"O��Q�"e�r��Տ��+�i��"O(�yG�'��ݛ��Q.4~�f"O9x�\*����گ4�	�"OXq�Vb�4\����ǡR�Y#��'��	�	\�o�!32X�nU��B�I�b��$A� ў�Tbb��iM�C�I7c��}p�� 3Hd fHB�#b�C�ɴ�I�&��>b� ���;A�ZB䉚?�Є2��)\�@,����4��B䉭X��){E.�2a&|I��(s�B䉨	�\�yQ�ѿ_94Q �I*/����� �fl��� ̈́!�U�!ʭ�|���n�\�,�0^�0�	��΁p�~��P&D����� ��j<{D���]���#?D����Ӳ9����	M;��l	w@2D��p%D#>��E"�o� 2�p`�#D����a-P_T�H�h�ãM#D��h�(lԈ���Ԃ�Lp��H �O^�K2��;�dN*������if���ȓ �N��1�Fa��*#._t >9%�L��2 h��G��L}�:4��>Y��D�O��$0��?���G��`�R���ٞJ5T�)c�%D�D�V��9(8��Bw&�kC7D�\J��OD#���m
W��;�5D�4P�*f���I7e�ިc�4D����KF&9J`���[O��0�s)>D�t�� �Bu�R�['Pe��ȡ<	��H��I\�h�L�"wmS&m��H�	nyb�|ʟqO(tr��}\�L"֭�  ��h ""O�j�I�${������Z�Գ "OJ�)Љ�2��I��iQ=J��Qa"O�;������j@�J�X�䥋�'����"AO�8T�Y�0����cA��w6�A��-���֘a��0*��oGJ=��P���§,�>2`<�+`�B��rX�?)���~2���6�,Z��K�5P���7#�u�<���N4W�����I�6Uܙ�ʞV�<���1���{qE�X$q�G�g�<BG� ,[�ЀtG78�q+W��fy��)§"D����)��,D�w�m���,O����Z�Y���W�u �"em!�$����[�I���ґG�ʌ,�ўD��Ӣ4��L �F	�h����)�B�ɂP���I>`נɳ����B䉈bZLh���K�����2Q��C�ɽy,�d��/8��=�p�<{�˓�?�����S�L���/ю7o�IzǛ"B�r����O�C�	$t�U˗L_�b��GU&^C䉱A< �����5���P�L=�:C�I��v����v̕iE�O�5F�C�)� ����ؤd��`�S�[,-f��&"O��@��hڌE��h$Q���Q"O�U!T�ɟG*<0���Q7X:�p���|��')ў�O���A&=e�Tбc��!�dM@�'���P�Q�Z!�A`H�!�Є��'~�e�s�^.��A�Z6��C!_�<Y�BH�?#��F�6�x���EA�<����;%�a��n�"ߺ4�fbz�<� *`����3n�6D����t�<ygO���<y$K�� :J,"�ny�'U���ϞA�n��R�8<���',�tS1I��&|�����%`P��''���s���EM�A��`�:��
�'��y3� @,�­hE�2[�J�;
�'�Pd�FV<:Dv)�+�L5�$��'9����@\q����עB1ī�'z�ٓmՃf]D��4`A�'�1O�n�47��
��׭"k(	�C"O((��ԉ5rĠwȁ�fj���a"O,��	�K�nQ�0g�9s���"O�Ys��&c ���EY<c�T���"O�p2�h�IhD�q"v��Upw"O����W�I�*�#�!�{F@�22"O�bT��E�"۴`F�b	,�c����PF��ϗ�
����ͅx��E8 IV��=�yR�I�n*x����ԅ �ꠈ��ǝ�y"���#�]`��з�&,c䀀�y�B�X�0.P0RTp��.�y<=�e��`��H)�/_�y2���yc>%����	g�ѳ%G�>�y�)"o��i�y�ؽ��b���y2O�>o<�J#��ket����*�y"(Ϸ8�.l�jT lq��u%�%�y�	E:#s�L�ѬO�,�T}{��[��yr���J�JC�M ,x"b�í�y"b��i�Х|��u�0�y�H_u�.Pp��Ύ=�Ƽ� ���y�%�>1����I��Ibx��ǂ���y�bɏ;F��A����;wc���=q�y�+�Z:	�uF޼�@�J&Y�y�I�Q����#ӥx�ݸpJT�y2�R:p���!���aڰ$� V=�y��"�hi�	�F[����\�y���1/��3�(�#];� (�yb`U1��"ߢy�>	�����y�dY���M�b��k���"����<���$� r�٠êۤ"�j�3���F�!��Y;BTZ�h��2�t	���Y�#�!��+�H��p�<w��.�9?+!�~j �tkG�U��� #j!�U�-���H�!�%gT?&!�D��9����@�S�Ȍ��ϓ_!�ĝ!_�VLxs @C�Fp��B�~��{r��r���c�(����eA�@�!�d�}N�;�JN2�!�q%K�!�ă�hE�%N�f,bt"EE�> �!�$�=s�( C�H7L
��dELo!��^[Mء��"��M8@�GCߥPe!�9+�=��EW�'窑��̐�!�B�Gȩ�oL+X޸9�F���Q!��9)�:�r 	��Bjh�����T+!򤚡nE��T�@5"�*�a��J !�D�P��ID��r䰭�r�Q`!�Dש(+��c��"-��Q1�[�.)!�� l�ZBhL�T>xb@�
 	�<�#��'���*	ra*#��z�� #Ӄ%��C�I�.��UB ✙&5��7��H|C�	3m�|Z3�¶!ʴ�V��!
pC�8r�N��w�&=ҭ�ݞw��B�ɺ87���[	v��%� f�7ÎC�I01��86 1 č�f���{�\C��J���17���P�����}��C䉀sD�Y�V?Gd���qN�$a�fC�	�j�L�shPIM���W4HF(C�I��h=	c���~�,��1��z��B��֒��Ջ?���)WAB/m�py"O�H*aA�Ē��Է��M	�"O�wi;)<h�RN��I�
�"Orءc�M�(h��҂7a��D"O�(X�d[�0
.�� 	/an�B"O�z�%4�:��!�KZ�C�"O>� G�U42Z�Y�q��9R�a�"O���3�($��т#�z�`"OV�i�Ȓ-	��"g�����5"OR����5l~�9
\&>iT��"OѠ�H�t��)�X:�5"On]�""�QH@�_�M[�@3W"O@e����T���T�do��1"O�8&$9a�F���J�#8�,�D"O�͚1��A���#G�	6D��ASw"O����:Y��ԫq�J�(����"O0k��6}���(N�O�E�"O�xX��ؕZ�2�IE&�!��U��O���#�
���҅��~����/%D���P�ěh��m�)��ig�"D��+6i�H_�ų#+)M��d!�$D�ˢnE1PDqɂaV�� ���!D� ���� �R]�UA��`޴�R�h?D�TC��Oz��8L�c(��`1h<D�@���'hg$�w��7h��HB�9�	ϟ���~�O ����*nN��T�Ƨ
�=Z "O�M��	���� ��c��\"O*]�2ʖ�cfB`�Tj%tt���"OLt�T��A� d�viӁ_�ڌ�q"O
�p�#м<���4���Ҥ!7"O��"�Mb@䳂b��Hy�0"O��d��ek�Tᡐ�=*��$�IN�O�8��tKH>`�B�ÄcQ�M�ahN>��MW�b�B9Z<R�J�b���$��s�D �G� ����y�R��ȓP�A�7"66���˛�4h�5��t%v�c�`�# �1�O���ȓ5�a�`��/�>���&T+�J(�� �N1�
X�f&�ICd��n�?!���?q��	Wvn��"I�
ݒ��/0�'[a|�
Ѝ/�1��YhR�0`�RNB䉎Eˌ��qcP!]ش�����~��Oj���=`�T��T��,0X6�En!���%� aHeĠ�����ԝ(K!��E7dZ���ԋl�F�`&��?!�d�;q���[D�� Ov��3��6T�}B�'����7�<�"7�Jl�����O�!�Ā-6t�� �i��Z���ɑ��/\�!�Ĝ#?$(�0��ȖiE�R�o3Z��	D����v�
$j�рAɐs"�Y�Wg3D�İ����.�<aG��Eh���L2D�q�̈́0��LZ�bO}p�����+D�H�Wʑ�[�z�C�AL�EP�;�o-4�� b��ʞ�V8��0+ '�f9��"O<ĩFC�D6q��ɝ6M�N�xP��E{�����fH��W'q�1R� M�!�WxAp�jF��TQ��ɂ�O�!��#4n8)v�~�haY�)]�a�!�d�CS"	ã�Hgp�;%HQ_!�$Z#u�ԛ���)Wu�3�[�.)���҄|Y����b	S`@�7D�(/�C�	bbJ��4JE�=��B��G`�B�I�8�(e P�L2v��s�:=�B�IU����Bn9i!G�ɐG��B䉚;G���@oԓsMV�Y�͛�n_fC�	.�d�"̡$5�#�۷l�XC�I�]v 9�D"��%��2���#^b����+?IbD�ԅ͐������ݮq
�t��*
�u2��Q7w"<p)GM�) ĭ�ȓ}*�����^>NX���>1N��ȓKIp����7Eԉ[�Z<zW����:�Pd�c"��IF�@��ϹS:rd�ȓX%;4���BW�_0)\��/��ӷ���������'W}>=����<qgÜ&����nN�K��B�$FJyB�'RX�2�%�<� ��$[.B���`�'S ���Gւ>Z r��P�8)j�'DQ �n�5����Q�5d�k�'�&���	�S' �۵	�c��̨�'16��ڢ4��t�D��U��P�'��x��� Fz�y�ĭW�y���9�'�H�F�P�L���;�ĒcF����(H�肯m�ڙ{ƨX�/��h�ȓU*q\�m�RM�-M5bT%����p��}�to�)>I��wF=-tB�IisN�C�]D\�h����N�B�I�U�ȭq��K#=�p-ýqV.C��S���i�F 1��� ���C2C�	�)�dpqNd0l�B�,���?��%LO�]ztOG���(�bU��U�"OP�m'M�GC����"I&v0\sי|B�'�Ҹ�t+�<<��񹢯� 4��!(�'����f	N����#�=�DXp	�'�j$�I;6�*(�JK-�&�z�'b��DA�KUR�	�Zk"e��'��hҩE7%�b�9�*�S�����"O�D	E�V>A��C�5�X"O"�:�֦M����yp���ђ|B�'���fŉ;i`Y���I�-�l=*�'�����'ʏ��m��N4t_BP�'�&�s0�ND^1��J�+h8�p��' `�K��ȵv%��-�h�zt��'4�Q��"_��iۛ�^uHJ>i���0=a5�E�RW.Wj�ez!/6z���G{J?mH��|���[�!��Lm��F#D�hk�� ��]����%k4~a��d,D�hs�+@��� �6T�>�"Bk)D�0
�j���6Dڗ%��]ٖ�%D��˔Eːj�@![e���h�i#|O�c���2�8�LB�#�r�L�1��!�/�S�'lT�|8�EE	S!�`�b��N���G{�O��ٓgH�v<tL_�'m�0�'�,I
��/3lqǉ:i%�	�'\�x8W�9\�x 	g*�b�8��'� aD�ȕV':�a֩�4_�v�'�d��1�R�9b��;�(Fk���0
�'�|�@g���%z���#�!L�,M[�R����q��O� ��[w(��G!$U��� �d�!"Ȏ�e$!? �uJ% ��)/�I�"O,̫/Mk���b.�?>�a�"O�A��/W��s7GO#F�v�{�"OB���J���&�a�^,j"O4���-Χn:�Ԫ��I���]�#�'��X�!m �D���a̦ ��  �.D�\�a�V2p�^�kT�J�]ڜx�t�-D�\�F��#	or�2��I�?2b�ptj-D�H���G=+,r���y���  �)D�<����E ���e�$�i�AL=D�xڡfZ��m �DG8J�͉��'D� �d�G*���C�`�9Zf!%D��@���bgv�8P�΅DG�� -"D�8{�A��^�Ȳw�Цf��\��>D���g`�4E7���G��S���*)=D��c��F�cG"�#l͞iAfl!�@=D�xʂJ�6~*�Ps�Ʌe<�[��:D�$)QS�S-�q �f«���Ӯ+D�D�a����J� �h��{�9[A))D���r��0�j̣��ЈKWl!9&D�`)0jJf�(1�,%�.� �'<O�"<C�Ogq����C/��|���Xd�<��W��Z �%!�Pe�t�<a#둸"��f@ވ'��q8��Zq�<�c�Īd�"$	�%����!�o�<iE�\�tX�`p-	���u�N�m�<�P�ټ{لLj�-�oi�@��m�A�<��d^�R(���|뀍�}�'��R���|
��7����1z ��B�<� ��be����욼7ǔ={�� @�<a&A�'2��P%��"i
Mz$a�}�<�'�^������I9�$�i[|�<D��e����ĝ����1H�x�<�$̔64Q$'ٗ%�r���Z|�<�� ��p)���`��=>�t�Q���M�<��.#�PR�Q!%�͉@GGB�<10�%+��������0�dQ���E�<��~��� �,K��r1!�B�<�%�W(w�*4�&J�$sF�*��{�<1v�Y�]Ḙ���Ʃ��P*�o�`�<�V�I�\����ǋ�����&�]�<A@`Gb�+@��=`5�Xx�<Fx�c��F�'����'(��y��5��ȹ�o]����yBbҼ7��T�#4V9�I:V���y���8Q�T�wA�Aπ�Y��A:�y������E�M�N���	��ybOA��u�CV��1���]$��'vaz�IL�yW<[� �;Ml(�` )-��'W�I`�O��	B��V��k��Gfp�Y	�'�|�б��� 4�8Pam�>��'n�-��
\17��*�hQ�yP��Z�'���pWdݽp���8���j�^��'��3G�^�,?Y��ďa��$��'C���7-!b��!��
L,;�'8�h��H 3�|�6�[6�a�'�z�`��T"B��Uxv��.Y*v�
�'�<��&lՖ)wD�`!��YL����x��W I{�쟫7�8��	F�yR�ў�<}�FC�_l�˴���y���9:~���I�[�*��A ���y�19���x�g��M����ஞ5�yb�*QL�Q3���I�~h��	��y
� ����nN�1�$ذ�HWo�f ZaY���Iw���O;�lA��C2p��-q��)vI@�'*|L��� 75f� �G\?r��k�'=����oi��B͈p�D���'2���ߔrŘ��2�^�3[����'>���ֱC�-;r�ޯC{�Q���'	`H؅��	^쉸!�1zP�
�'%"IkejW ؍a��&�Լ��T�8��I:�t|� �M6{��5D��M0xB�ɉ���e&����WAU;
�C�I�W+䈪ď�#^�FQ�g� 	�^C��W�`���KV:~���',]�<:C�I6�\���n�8 �A�W�[,O2�C�ɩ'��I�p�V	T �9����+ �����n��Q���xSO��Լ�e�/D�D�6J-hm���O5P%��3a�.D�X�#���u�~�8pgҸ�LdI$� D����@P���y�d�L(�E���)D�LZ�'\1�U�!�֌��h��<D�H1���7MxAt�S
;P��iQ(:�	L��@��Dҙc]$D�1o�_+N���6D���c��,rZ@��7%0�b��)D�,�$Őgpi�@`I)�$!@)D�C0k
=�h5 ���Gh:D�tڠ��56���8si�Y�()�@3D�`�q�K8A&�����`M&9�U�2D����I "dq�X�F-U�EC�m0D�,�C/�^��a餍L�k�UJ�� 4���׈��Sa|��5g��%/��뤌TWy2�'��\Pv�Ŭ���&�L�6�jT(
�'|v��S�(��y��d�Xz�'�N]"��'$]�U̙m��4Z	�'3U#�e��	�L4@E��h�Y	�'ꡲ���Q�ց��Q�`In�		�'%j�1'��5y�\�M�x�5`�'�p���lԒ5JJ� �*��A-O����ɽ O����!�tp!����C�!�K p�T{&	�Os��@�\�K�!��N(}eP�y�
VCbx4���N?N�!�ğAW2)��,�ȸ ����!�ױ���fͬV?�0x5aF�x�!�dF�@�R���n��a'	�Ɵ��!� ~iT�ۥ� (DXZ�*�J�'��̑��ڭ���0�,ߺ��'0��Rb�
R���$%\�;�$5I�'0~My��j��تaB.�,���'�TA��Dڸn��i���O�rB�*
���qT��BFMU�$�p ���\�g=8Y�	�'�,���I��X��*CX2����'�(l!C�r-�Y����CW`���'��D��lռr1N���J�8j0���'�X���n�+Sՠ�YG��/$�T���'�R��ԯU�u��!3�)ΒoІL�
�'\��ԀDOՒ��g�o����
��OB�e��p��Rn��4�ȸ	�"Op�Ph��|�c���Zy!"O��w/ۘ;-:ph!��=-�	�!"Ofq���<n��)�Hݗcl��"O8Q��6�t���Z�T���"O�|Ï3JCXia���';~�3�"O~����(p8axѧ�h ����"O)��[�X�'�>*��D�|��)�ӫ[�ҵ�å?�P�e^�*x��D�O��@�&�Pv�ݱs�rA"T�\u��S�? ��ӒDR�lƮl��#B`���'"O�,�Df�<c:x��˔hO��2""OPu�DL�=)�s���|��qV"O ��s��Pj"�Tr�O�)L�ȭ��.L>8�A!D?��z%4-�D�O�=�|
�/ �]������8䘀�7����?�'7�Z��U//�^t�"eٔx�d�"�'��q�c_�3w,i����$��a��'Æ-���ɬaVt�f�ԏ"�Y��'b4H��_�yd�ݓ��s�@��'p�xke�^< 48mr��*4/�E��'��A(�K{�Q��O�2�d$A,O�=E����F��d�`IϠn��Ѹ���d�r�'����Q��J�JO��B�s$ĨTx�B�	m�nBé�9�$�!��k��C�	>���A��!l� ���aH��dC�	~.${�
Ό%��Y�Ǆ@C��Hm|�r�aE�?���P�`M3v��B�	(�*-���X���xJ� �]	�C�	�'���O	5#n�cE�A?�NC�	�!oZ�1@��.} ����a�(��Gm0=��S:NUw��0!� �ȓmFM둈ܪ\'�[�-i����Z���rc�O �B��B),U�Շȓ��c�j9g~��1�A(_�:��?��0|��@�I�\��� �~�2؊fcS_�<)f�E)������ 輜J���Zx�(�'(X��U�&4^����C�=��Mc���x�"�8p�l{��\��(�H��y�+�Фӓ�У��j�����ybgQ��2�תK'~����Uh�	�y��(3�x\�3f<z���#&�;�hO��	�ɒ�� o��8tİV?
�Y�'	�tX,�81�$	ySm�\�t�.O�����4'ZVm��*1^�<�]�!���:+��I���sDͨr�Bt�������+Ja&$����
��`�ȓ;�(HYѨ_'������)|����q�)�;O���$+�l!j�%���'Oa�t��$  ���#��0_5���� ��xRc+_<N�ۦo	���'�H;EE�O���GP&Kآ�j��Jn�؀"O�������_?*9�aEl/j4�"Od���j Pr� ��)���D"O�ű)ޓc�z)k��E�^�t�b�"O��r�N�)9c�+����{��px "O���W�-P�7!�8 �.p"O�A�W�3"�e�r�Xw ɑ�"O����5q��j���`�"O�0#RK�Jа��Ì-9��qӷ"O ��5@[$6!��6H�t��g"O�|�0*@� *�����:\�|y�g"O�S��0b@�p�R���%��"Ov���kלUO��(vh�1̱��"Od2ef� �z<�F���A�"OЅ�o?^��M�c%�r֦X+a"O`�"�ߵ�]0!�^�r�xB�"O�)��A?*8�v�
	S@�=[�"Or(�B�R�}��qX�`��E%��9�"OFEH��H�u&p�E`�$ !6�z�"O�!����[�iY��
�+.�q�"O|9��'Y�`p �'��,�a��"O
pQr͐[����3��M�V��"OP�)�g�4��To�*}�^9"O� �#�Eƚ>�N)��g
�T��"O*�1BխҊi��&�6�`d[�"O�za���(5��J���6y�"O��;�D��>Ҧ�:�
rw��"OHl
g�#E����I#3e|��S"O��񇀸r� 1;�
�OP���"O��2��\�5)D���=u@����"O��4�/\�b�A�MR� ���"O�p�v!Х7�����n������"O
}�2��,����-C�F����"O���t�&�����U(����"O|e�f�G^�qB�L��F���"OL�pP��1)�4.!�D��@�&�y��΋*�h����qf������y���<����S��hB�`Kv���y�IE
3�P���A05� e�#O-�yRa�;�FH�F���83B���yr�Ѹz��t��e���yn�-wNb��ӫٹ��Ik�8�yR@��M�2�3g��2A�[qŝ�y"�L���`��ˆQc� ٌ8!�dV�̴�qP"���@��.9�!�$X�T]��.�o��u-�4D�!�$4;8DB ]�;���¢���!�DD!�V� �$tϬ�ء�ٜ*�!��� w��P� �̈!�Y:<�!�$�<�H���9J�.���-C�w!��0-�X�X"ݬ���" J�
	!�dG87r@B	�e�p"��< !��
 nKHT���
L��0�&C�Vf!��H8%�C*A�zf�I��HV�O!�_�ȓj�V
��Q�A!򄎳%�����,S�{�"XRq�#!���5B$��2ʕ�:6��K̘�!�$I�O���Ԧ��|.0�H�-W	�!�@+o
\�ՀL>>�Y�f8!�dE��t�q��G&IB�F���v
!��JpJE���Hp��H!�nD:	�!�Ě;q�R�PF�t���B1���!���k��zu��'g�|�%�u�!����Bc��Y�J1�!����':!�&\_��X��Ŀ�܌Y�O�YS!�σL���k��F$��!H���4*!��N�5�.�ȇJQ>��2���'b!�ā�Dk�k���)U��v#Ö!�Q o/�QKD�Bv<�����9!�DU�d���u)V�*8��)V�M 6!�d�'E��9i@j��MP$���T�!��E8R��Z7g�xy1h��}�!��s#Z���ӈY�4;��B�!��w�.`�H܏8�0kvFM�2�!�AӔl9Ā�b�ıa�v�!�DM��9�
	(w�j�	f�w!�DHCJ8�X��P�`�zfDŽA�!��C�prj�bUJ�8��'��w�!�d��X�D�v%�9o��P:2�^�!�$U�T�r(���<, `��ꇅ:�!�DTXn5���}�l+d��'>!�U��b�d��w��b�jR9!�H��z����&SYr��̕A6!�$)t܄T[�i��wR����J��!�ᾑ	D��x;�i�*��G�!�dۉAƴ�6@C� �"��	g�!���-4AY��>�f���[9i�!��  ,caIN^������;�p�{�"O�qY ZRjQ���A6!�z��S"O�a�*,��ч)Q�E��Y9"O�U9s���/Y԰�_�A�.)�1"O
aȓƉ1�\	m��&y��"O�D���ZT��'��%��20"O�9`sD�z�)���/S�H��c"O�=��\%l�s(E�� �(�"O4tX��ٝ4h��ۗX?ņ�b�"Of�8iC5{����t���"O�1�c߰j�@�Kƭ�;M��=s�"OB�kգH�{�R�����?x��Е"OD�R\����B�ҽ'�x�#a"OЈ���ÁV���xe�J�SĒ�U"ON��b#�'�(�#�v�"�z�"Ov�[��]���	e�>)�b�iu"O@��%�5-K�� L��`�"O���+ʃ)R�Q�t�G�W�6�	�"O�����y����u���)}��E"O�:��3�`�L��K Q��"O&�
r/��&����X5Q�,p��"O(���%&�XS��=�4�C5"O0�C�9
�v����G�4� �	�"O^��у�0|�2�B��/��L�"O���.��G�F���A
���@"O}�G"�&r{�X�`�؈9��Y"Ojx���t��e�E���$�hu;�"O\��f$՝Kq҅�R<pGh�"�"O��:�d�*�h��d��R�b19�"O�D1\B] !`�%�VvexU"O8e�3Ĝ�K�N!�cJ�mCR���"OzQ�`l�#M*���`ĀQ(g"O�� ��l${�H�^d�kd"O�x�Amϙ�~�YMʩ+��4��"O2L�3J�6�ds�KȐ�@5+�"O���RiK�D��XƭЬ'}����"O�9�2��>."�Xa�m�)	Wn�jt*O���l�?O�n� ���>�]x�'7x`��O FQ$Y�f�C�<jd�ʓp�Za��%Љe��k!��1��ه�A~*!942-񤉨�E�y~��fn���o	�\K� ���g�ŅȓO(TR�F�^�6�r�^�E����� /����� �JPr� �`���a��KƤD�r9³��q���ȓz}
XP� Q@�����{��E��_]2D��M��	�D-	���A��:��q��.��C�o�d�m�ȓ=�����C�������L�	�*��ȓDqH�� 	u,��2�-f�td�ȓ*̲�:�A[�
8x [r�P�b�����!/6�S��jLtM(E�^�T{�C�	�c���#�_�K$l�B�̸%^HC�ɼ�.h3�ꎅ�`Y�
l�'D�������*)���֞��ҡ'D�d��D�*,uɅQQ�2-P��8D���Enڌ�X傴��5B �I�8D�H+����q,�s�j�1�=�	6D�8���CH4�zY�ΜXra���!򄀸�6�`�#B"aA�B�!�N�$$��r�b�0&E���Ҍ#!�$�&t�*V���z�Sp��!�H�3�6�(gd��7��#�F�8�!�d�%C�mc�6���`@ZM�!�� l�k�[/]s��rb-�?\�ȉ�"Oz�c��_=����6(���"O�ѨI�<@�qP�71s���"O�8a�Q�1|�"�}"0H�"O"�x@��e�r�3��	R�4j�"O�`I!�G=d�"wASH?�%J�"O�x{��X+J���7�#��A"OL8 eRm�����G���"O��Bk� ���iգģAΪ���"O�=��NW
L(e�,7��	 "O:9`�[�#	`�P�L��t��b"Ox9��ƵP0�'�߮p��"Oƹ1��6tE���d�]�@Z�"ON�S!ID7�L�@��7���"Od0ه�?\��u�Ve�6:ײ�b�"OD��Wg�46P�gβ1���0u"OF���Ѱ{HD���5&~vy`'"OB��d�1h�$���AŞRk�-�"O|���NΊdv�0�sg_(���"O�PyE��09jQCw���@R�"O�YжE�_v�*ĥÑ?��ʴ"O$����2
S@M�E��{���"Ot)�Ѝ@u��Ѻ�� �����"O �3hB����z���G"O��1���6BkV1��*��1��D�R"OH8�0��1dڍBTJ�08+$���"O2Y�� �Ecz̈���'!��+�"O,�� �&u��$����X�LL2�"O���͌�l�|�A��*v����"OA�N�3<|�3u��zi2�	$"O���'�9Jn�%Y#��-e_��!e"O��ZC�M�k�e�V�Q�"OZ7�ȓzP8��$ވ\(�ѹ�"O��[��K���Q�K�D�H+�"O2ɪeûm�l�r�V�}�
��D"O��B%&S	-�`��̛&6~��"OB-Q��D\p��A�-�h
�"O��	��D>r\��Ο�S�� �"O^��E�q��J�J�W�,���"O�a�b(K=<���錬^�i�"OT(@.�6 ��ek3�CY��;�"OHY�V'�Qކ��Ӈ��M��a"O�����xV<��.A6:�z"O�� Dމ
a�T��@��:-�]��D{����,Jݺ�HX�y���3�!�T�*����4�͋f_��7K��(�D�<������gHH�m:�%��l�.5�B�	=1m���FK��)I��. zL�@��<�0�c�ՐA;f���2����Mk��	e�xK� �/!N�&�e�<�!�qAp���l�Ĺ��[�'��`�� sS�ܰ�z�s�I@�X.)�*D��2d�Ӭ!���ŌQ�&"-�uH�,e��DAa��(�8m �
����a�K�q�n,�q�'K�Y�=9�D��=4�zUO��4�!q��Eܓf�7�<���dU���P l΃)���+�J�(����'�������9�EH,�=v�"��|X�0G��'�t�If�O��5��g�6 �<���'��k�I��;W����ζ~,<���'�(�1BG'9)pQ�D;z:¡��'N�x�B��[��À�Ts;t\C�'%�kV��9# ���"� 57<�
�'���S"ׇ4L(��`��!'o�1�
�'�`��u���&v|t�`3�0�I
��� "}��n5F)t�E��P'��"O�e"Eb�%7Y���A�N-j�zȓ�"O��X���%`����i�A"O h(��Ǟa��`Rn�v���2��$4�@���@�t@����	���� -D��� �,))�É!�¬��(D��S4�Ďx򴨊�Á�,+#�&D��hu.@�j�<���N�.�<�9&b1D�xI���
�X�U ס$�m��4D�L�u���ji�L1���m�ܱ���.D������0-IpdbG���D��e5"(D��Kq	���H������ђw�Gth<�6��.Y���� �*{?�<j&�_�<ɗ�SZZ�a�Y&:��J�-�Z�<!$ �e����%=��AQ�C^�<6g6k�Z��#�(F���b�<�e�O �B$@�f@B���RdMS\�<��_y\�E)'��~����JnX��<i�'N��94}��� F�C
�'����TȂ2o���3��OE ����>������ �?m9�`�F�[q���"O �䍍.q��<B�K.dg��2��'�Q�,�1M6yo��6��>�(���=D���p���q�",�&ƌe�1A�O�B�ɍ`-d��I??��xsA#��=�B�I�82 ��@mѻ|�\�S�//��D2�Ia}���O��Sg
�|Y����^��O.ԉ gA�Nl��څ ޷RP��W�Hy"�'���JW�*n��!��d�"p��'R�5��n_�Ae�qiJ��X����'���(Ԋ� �\pHA)ބS � p-Ol��hO��
<} �x�X�z���"���6�
���>I�h�<9Th0 �.l�ԫ�l�
��w�Gz�<QR!�=�c��<����m�x����'���c�� �%8=�7�̎���'��d�fD"��@qwo�^n~X�}�D2�	@����U��n����qI�gX^|�ȓm��Г�@��o\�{C����>�����ħE�(2&ŊZ�F4Q��ؽ;(P8���A�'��ݘ��b�<�a�e�(w+��P�^�L%�$s����M�׬�YWf���Cc �}�����T���2Ge���!�i4D����l5Et����9d�vi$�/,O��<A�&�1l2�وL�4g�]�f�VW�<���'E|pPD�p �Hk ĚR��L�'���b�N��x4`��F�a)r����'��q�N����;�#�7[�<�R��D<��xBথ�U�&�ض��f�X|G{2�O�aq����o��1�Z+���'�ў"~���kIbi�$��k�Ĝg�:C㉅Kߴa;0&�g=(:�Η�in%��M��/�T�Xs�Vd����c�=Z4=�y� �a�'	��u�4�M������X/&��'�Ґ�IJ���=�=Y�"�>���'rJ���)��
J����G��s�j���OZ k������Yxl�@�7�,�zG,E:]���dBd�iL�}�%��S1��C�'�.R2`e���S]��p=��#I�\:�T!P�K LW|�P`�R����	����Vd������rA��Iح7Վ ���Bf���R��H�pHD��ȝX��� �Ԝ���>qF.gӠ#<A��͒*R�
"p-�;��c�� .��?G���]FO��rwR<� $���Z��!������?�|�m=�0�1��r%�pj-��'��O��'hF����l�:R�F<�R'\%OX&�e�$�S��y"�U�;��Aw�G)%�1�ヅ��O�#� ld��iX-.��=`!BGzXp�"O�Dy%g�?X�z���>u������`>��c��$`�ȹ�a��47F4��:T����$[�p��|�q R1B��1B"O��s@���/��H��nYD�4HР"OZ�Z�"�~���U �(#�|�0�]����	�jp�"";��Uؐm��C�	Qs>�"��̈L�}��o�4f�c���5�'ML3��4��)���^�S�v���'�u�&��E(����ȬO=����'P���I'7��BE/?V[�ah�''�!�� E�ZI�5�d� ��y�� �����#�)Q���w����y2�«o&����C�PIV���0=�rLؔr�y���;8����?�yB!٥0LP����?(h��%N���y��ڈ������̄�4@Q�<� C�I�U�r)�'c�9WPh�p�ʒ�5O��=E�$��4r��)�B	�aన����0<����\~KS� ��`��$��!�1O�����n�j9:e^OC��r��K:󄐣�(O?9!��d0h�D�8j&�����8{	!��
q���� J�Y�P����2�axb�	AD�0v%�U��8bݽ	��C�Ʌ^�� Hfb�./u��0�Z(�2��hO>52�%QY"�C��]i�)83�<D�,�T�\��$Y��'��S�Z���z��]DzR�I>{2]�Ԥ�>7���aŔ�;Vz#>a+OR8��i�$�"�W`G*'Y��(�g+�!�&:W\��	N_<��E���8�Ӻ����&�P�*�,F('\��Ԁ@!򄝿eA2i�kM
K��e�@Sݑ�dF{���!��\8;^X	��1� 9"O����G�!������1��A�dW;2�y2ͣ^��(� L� �`H�y����f��CB�!<AÙ�}�B�93��+����(��覂�V���>�V�S'{=|՘�Q�l�~�C��R�<��ϭi �e��Y�HC���z�<�O�K��H*T���
��Z�^��C�I�a>�P��Q�%c�x� KQݪC�ɼB�8S�S�/�biԊ��e'�C䉜/g��k#�щq~�Ac��*�C��>F�l1�D�a~x��$`
+��B�I6fH=Y�Z����YO\!"^�B䉏b��]�$[���)��l	-D�(�e�ɔQ	��
��+?�n��W� D�<P�J;PJ~M���>P�r8#��?D�L{q��%y�r���P�-�{�?D���A
S�Rr֘X�.No���'`(D��N4H|����&��bbj(1�%D�0���5H0q`]22��s�]/e�!�d��BJ-j�
Q�����A�)L!�4�R�j'f��M_���NDVF!�ٜ6Xx��B�q�T�3$�+*2!�� it��\t0��'!�%*�p�%i�8c|T���= !򤙬7�xع⎖@���P�t#!�P�s�V�(w.	14��S��M�6 !��+O��2��{��ZB���>�!��C;*� �h\��ԜYҮR/ !�D�.�à��q���@9!�䇪s+���P�~��I���]�f�!��H�>lʦH;6�^\{���EW!��  ���#B�
.�T2��rU��a�"O�ĸ5&��W@�������t8��W"O$����:sd�0t���J�ȱ"O|�jr��x�N���A2D�A�"O��I����q���ǖ��C"OHQ�� ��BfN	*�|��"����!��#aTl#��D�:�]���n!�$�N�2����P'v�	獃�!�M���
!�X�03F"����Pyr�
Ȭ�� '[i���c"�y��-6�0d�)Jip5q��.r�6� �3�0?1��@�{������8Z���aWr�<�RĆ�w�: #� >��(x�`�r�<! e�5xx�U���΁wŻ�lw�<y���r9qd�P�H	��l�<ɶMN!YDU���3|�Xa`�XS�<���)|��q��7N� �f
O�<���5]�F�-Z�L�S�WF�<At�P),,p��O�&:�Cd��T�<�a*G)�MrWLܶyx���i�U�<����P:8��G��T�,�җ��R�<��ܾ>L I��Տ7vm��$T�<�6�C�:���Ef_�'�[�CET�<��K�u�f)[����ʅ�KR�<�1�YЀ�p���c��-RaLS�<q'�۹Xnn%.M��]9w�\W�<a� ʸGd8�L
�!ɪ��C��Y�< �E�"�4d V�ȳW��`۠��_�<9��7�PAhPO�+"5�hK%�w�<��$VH���y�åSi�u�2E�p�<�k9Z�аzS���e(���6	m�<�W*ľ?�ð$��b��=��ǟA�<y'ƀ+S� �QALP�6����e�<����&2jJ�j���xiG��h�<	F��*U�\8T���z�5�ҤNo�<鴅�0$~}25� �l�f �5H�A�<�ƌY� ���L�%}� �DeMg�<)�  �F`�BӞc`�0��lCa�<A母9=G�B��J�5�L�e�LD�<��
��*sz�`&�S8I"0PW'K�<)`�9 �*�Qf�2x��2r�l�<ɱA�f�&����_`�U⅊A�<9�,���������5^7*(�a�Uy�<��@.���R��3s���*�ēt�<᳎�S��M2�ĳ8���S��n�<�fP<� ��B#ɨ,�L���w�<�1�S9^�h��d�NF�"t��s�<��cYC�:|���85�:�j4��`�'ɌZ�����e�6�%H�����R�)C�(Ė��&h���y j
+�0�	�C���(��0���0M.�t4"�OX�C�I!D"��F	K�P���)�4s��'-P� �œZ��(�F'��S�M�mC��p�i8�OeBV�ڜ&��(Iի(qe�-��G�i8���'�U�!���Di�P�) ::,��p�����I��R��	��>�B�����0�
�1�eߦ�!�$>k�b��M�>d�դx{��L���xʍ{���"��t)�R�B�Pi��K�ƣ=�������l��Nמ%R<����'oX��r�x��N��z�D�&�l����[��7�̃�MK�#PR�"~nZ�{�X�4$K,#qdi���@ޤB�ɑs��0�fE$vV��œ5���6,6�k�j/|O�q�%ˇ5l�@t�G˕�x((�oX�ԋ��)>��D��Rv�9e+RZ�`x��jU��y
� ���ӛzVx!eJ!�f�`�ɋ3�����퓋7Dp�a�6X�&��/�B�	�%���q���"�,�RR�ԖY�7��>I�eC�{���i��Ȳɚ91��!q$B��GR��K�'`j��ܑ5���h��T= �-OҤ���1�O,p��i14Pd��Ǝ+O���"O	#+ǳJQ"A��/'n/xm
�'����%$uhG�E�]�X��'Lr���޽�!�Q;Q3d=P	�'y��Cq�� Q��2�7O�h*	�'�@TYw	��Q1Rfg]�Q���a
�'�t4��!�0Hvl}`sB�N�6"	�'��D�bT�PR8�ز��O�y��'/���Ϲ|_nKg��/rT�D��'J��4��lT1C� ʋe�ʽ�
�'&T�{FEV�A�I�"i�9E��	�'ޞ�	u*�:Pvh�(ѪUF��	�'�<)R�埜Ξl�P�ېGY�'��@x�DKF�S�O:n�R!Žu1t:5���#���k
�'���fW ����'\m���.O��b4jRq"���:���X�ᆶ{}T� GԷ3x��ɜQ�0��Τ<$8H�u�G�Ml�5h�u�؀�v�$^F!�d���rq �
��D����.��'�@��#��~�>�aq�W�B���B�(�On��O_"Ũ@g�)RR��D���<ʚ�{�rͶP��A�-��遢�d���I�
#[K��rn�/�q����Vj��$�
�(��$pp(혵H�m�eS����1Q��WGZ�Ȕ�m�6Z�SK��{#���3��S�C=@+8|��/�:6��P��=A3*�+���Q�T1��W�z-��(rf�2������Ozm���X�&o`As���~+P͓{/��8R׶0��g���j�!ԦW kB�:��?o���hT-�Ahr	��lz�m�g��h��Ę	{���Uc��B��7
Qnׂ���kJ�^7�! $ ��}�-m���diYt�G��"�� 'ڠ�ݡ�<C�`N��
x��F֠�D;F�dI�';�]$BC�f��ӷ Mb0�1�Z�������n�"lp!
]�g�j0��f�=3���n���;VIh��S���k�.|`ɟ��	.k���p��B�R\���tn�P����&�N2"�;�%)I�N��ίh���a�<QV���.�S������C)0=��C̏�A.Y�qA��sv*�Z�X�B��Z�Bp�Y�?A�
�M�``t���"d��b��ߞrd�ʑH	�@
�	�J,v!��y�@���p@���$h��:��ql
��Q(�B�#P�> 'ܸ��گ&Ĵ�fѿ�V���V�yKZ�1q�ѷYB�	A댣�u�Q�kQPh�+�,>jD�Wb!!-�&E�p����æ/s'"�8rbPlZDP��/?hL�*7�B����f%L�| &��qƇ�7f���
0��dO04�Q3o��2X����f�����&���,�2��aׁ7����#$Y$�}����w,q�.\?m�d�%�Z��QW��2��ՐcF�~R�'��a0�c@.h=���AT�__N	҂�6Ĳ��MP��eE�#(��I�#�.i?��4�T^YT�w�1Ӳ�S"��%��Hb�Ib�3,X2mrܐ

�<i�Y�u���HqǂQq7,���zpb�d�	[3h������3]Ɣ(W@��h��<���	yjӱ�̉r���F��"m���0�Q�[��#`fw�����O�'�ݓe�[�'��m��M8��={GGE(K�!�1	=�&'��+��yZ�-  jw48�C��iq84���'� �f��
5���'â*����59g�\M��9u�N��!�F�A3B���j�hږ��5�`�����k 4����٪��\o�5���҉Y���7�ܭzօ���[� ���j�O�ъ���	j�X��s�X0�T��� � Eĉ^v<)�(�dD�\|(�c2�J�I)&F����	A�P+��D�#W`����5 ��ȏ$M4xA(Q��I\�I8As��X��ϕ1���CS�E�Q�&���`�T��T	s�>)AF�Fx�R޴1���Ss�EP�"�����V��TRe�z��Zģ.J &�Q�-�%TQ�"?�h��8zE"��<S팖@�ݲ7��8�II��D41��`D�i��m8a'ԡ*����42Y�ST��t�	z���m �^��e@�z���I#(;}���9��!�?��^*	��@r�A;��\��A�9]�����$&��#*H7`c>c��i3���{�ISAOӅ����`�֞3�$i
)O@sS�޸��T��A�(�n�f(2cH	�,S�d��ɛ�M�|,���'�<1�񈟘q|���T:
T�U6��y��h�O��q4�[�WJ� hћ��(!�� �m!�h��
1j�%jQ�x"ĝ�(�=Ad�
)/��I-}�嚑���[�BВB�B���n�.�@ eD<u�y���S���t��C�8$�(�t \�H̐�'J"MH�i�
��=1��tU���)X�R�����暍Jj�h�I�^��Ʌ4�bXh"��|��[Y����� 0vv%�����xq��E�<���ܔk�^�>�'Vh�C��I|�hJ�c
4h����B�ܒ	��''6=���D�7f?�hsD�f��#R����e�#M�D@`�@�)�&���d�>F]��	�/f9�H[�%�9ڠE�x����N x[������ 6h�U�̨M<�����Q�n�������ORV����È�d�@E��bh����70�Xؗ�|�O71�Pȇ�m� xR�N+�\��ř�=(8b7��!����N�jZ��ʣb�#w�FD�,O�`�5,�кLzP@M�'�>鹒�I0
VOd�'oH���0/N Q4�أ��I.1�J]��d����4B5�=h��:3(T��O�t�ү��8K�mZ�N߽���&^� Q	ȹ~�qO�.ӓu���e�@�sc4Mч�I�Z;-Z�h��cu�A0�K�&<����0�Ot�"��g�A���<�E�|��7�> �5�Ǳ-��*6�] �6u��)�A��aڜt�umT By��+�
��?)��V�d�LxӢb�$&
e�C�L�aِ!��Ķ/.Rer�"Q5>���"�MY"�J"|�'���*��Q�8}B= ���]������Ej�����C��K�½��S1�~�ٕGU�Z:�Y�Do\�}<Q(�k֟[vL���g�'��hiS�S)&�pa�D3�%�OV@J�H"�)��Q�xV��9D��>��Q{��3AV6Q�K�5M�D�s�'qZS�#��!��M�enx*���E�#�,�j�	QO���X.�0�C�K$���#�K� ]�!�$G2l-,1� �׾	ɔiW�n��D	�Z N�����'N���S�O2�e��+�%�6CDGH��'��%fVh $��U%�=^N1��>Y3+
�\~��B@���}���9M�b��7HSp�i�]���?���\9���%㌄G���QA�`������	
�x2D�r}��Φ'��x:U�ؿ�y��ʙ��X��(T�Y�����Y(�y�F�D��!��94-�� $G-�y���4N�6$-T�8اn�z/bm��jˎD�aV�+��ٴg��ix��@�$ldC�ɣ��2��	Rπ��M��	�"?�Ì�K��r���$� ��Y�+�=��.6�y��`)s`�dZ��uK@�Y�-��'�Ji�J�X�ɦO�>�w �Q�FH�J�ljŀQ�=D�`zQ��P|�ժ�
nI��;}*�&- �Ҁ��w��A�kX�H�DU���C rĉ��6�Of����ܬgx�:g/�iyv�i�	�3a��eY"�ߩ�xr� ^*^Y�U�d>x�5W�OJ�bT8�^�[��dH�k�����ӥZ��Y���	�y��I&N*h�BPkH�-� r��~b׃_OJ\�ࠆP��S<����E�R�[�J���
D?\n�B��jy@��!�1@v��"nA��'��j!]"����(��E��o��?}j�̎�3o����L�/����/��I��L���ԣMB�`+@�J�xђ�'qL��G&S7r�&�c,6��P���<0�����8�,O2�ty�Η�1P��s`�p�B�ɬ212u�K۴P�&���O�5�˓m�F��T�#�)�'I꼔��M�;�:=Zp��L�>�ȓޒ���d�;ðHQ���!��8��:ı��.!�AG�%[	�<��G�$�C��;��ɢn�!R�� �ȓ:0	�V���P�zU�ܘhl �� ��@(��RI3dĄoÆą�U��*�cF1C�&���g�\�|���	����o� ',(`I��mܸ��o�vLQi�0��0��"�6!X=��)Pd��#�q�~��� �����ȓ8B�@��ōpB�� A�r�,P����*���f+.m �	�7i�R��~o�0iׇ�
Î$�B2MIjl��\,1ؑ��Wn~���gN�@}fЇȓ	�&�f
�9Nۦ�e���4�
�����JB*�$H
Р��~B���r������֛+ �`�N��
۾��ȓI�,]*#`%3e�Y���z4����AƐ5jQ��V�0���w"�E��N�V�)�	2� �
��f��U��#E�萦B\�x�.��gO��Ԅ�S�? ��Å�Y#<�t2�ꕀn�v4c�"OD�`s2�1�GРN�`�p`"O֤���%�z2@�;DR0�"Ob�aAK�ː�2E6G��E"OȰ:��1�-�B�ٯ-�<�"O6	���6A�:�"�D7#��"O�( ��.=>YˡCY$^��0Y�"O�c�2}���@���?$DY��"O*�K���r��B� S� ZW"O�a�BA�~l�p0�J�dd~�qF"O�@����&�p �l��+B"O�����ySv�X�J�L�,�P�"O��Y�.�V�n ��B4�T"O���� ��7P:�Y��i�|�3@"OdB�MÈr�.�j�`e���w"O(Q�5�4�t\q�O�$�XU��"O
��F��M��#0�&rP��"O~����]�M���
gAӑw\�"O� E
˓t^"υ�(Cl�q"OVY$�S�a��� 1�	G_���e"O`Z�Ɉb+�qC �88���"O(͚�$��E����Q�W����y"Ζ+4��\
��KE���/�,�yr+1K���x�˘D"�d"�M��y¬�qީI"M�0j���'��y��6b��l��	���}Q��R�y"dD�^u���"Bc�@�CEL��y��ܚha�Y�IQ�X�ȁ�a`R��y��Х�4\	#,ϳL���B�/��y�+�-��Ԙĭ�w6Hh�rԊ�y".�D��!
S��p7l���y��S�9HU%ň<�01K`�R�y" �54<�a�ԏ)��A�����yBh�[���
t(Zj�)��ΐ�y%��4��<�m	�f�YBjU��yb��7i0����~a��'&֤���'	F|�6D�T ��,��I%~�k�').��P��d_Tq)�;A�¹��'�*�@���y���0�̔�s��D��'���Z4G�:Yj��ru`� Q8�'S�ݢ�����u���D.$�ɹ�'�f9����8�da�4&ɑC���'_�� �A�|dE�d �?/6���'���j�u��BE�BhDD-ʧ�yK^+nz�dM� >8EJ��yB��D�L�Xץ��>����2
Ē�y�뀂4ю 
��U6�R1KuJ��y��,!v��S+�.}4V`+(�yb"S b=Z|��Nq���A'���y��c�
�)���Bf
عf���y�)�0���	��� G�2�(�4�y"δ`l�]���Ԧ4��m����y�L]*,��p0mW�7A>�y���yb���y
C
��80���ao��y҂ۏ'BJ(1$��9����ࢍ��y��ʊpel���¾.(��fP��y�hʺ5�䈲�K�u5PYKR�H6�y����X�������$���y�,5!'�a�g�}�L��� ��y�ķ �h9�Q�_"w0�тuŐ��y�@;�� N���0Еb� �y�f�� 8b��S�8�����y�HГZIhH�d��
{~�Ռ
:�y"	Zо��׋�6��s$�ļ�y
� ��B؝r����#8C�:$"OR�� ���Q��%�tO�۸��4"O$���\�2��9b�O�k����"O�I�,:R+2���.�����s"O��fY� P�]�e�F)�j�a�"O6p��瑈Kp�Y南�*��
E"O�ؒ2/O#o�r��uE�~�<�"O�4"�iK�.��P��E�Z��\�"OD�9��O�ddX��փם;S����"O��WD3T*����R�a_V)�4"O�h��$>��%�S.�[*`P "O� ђ�jU!v��5|���K^�<�W�4kR�:(�.JEڬk� �Y�<�%@�F����$̀�lj&��!�~�<A�@�z�� �b�`P��C�~�<pc^1c���t���n,�E[b�t�<Q���.e��tRRO�ft�36`�[�<�g�R���4�eܛY��8��h�z�<�4H̶\%4����h��a�@��r�<i��M����$��Hx
���/AV�<PoN2d�F�#�`^M`Q��eE�<�!O��%O�hC�n5��I���@�<Q��ۘ%*��/��H@ i��� p�<��A�t��h�f�4���4Ņ[�<�螊�@q#2��1u�ԙ�j�W�<�f�2MH�X
$�A,9\>��*SO�<ɕ�
) ��k2�7q�$��2��r�I7p� ��"�'����d�R�Lu�`��==�b%�
�dR ��͂�-�^'L��e)��}D$��
�'�"ū�D<I_�\��G�;�������<xKZݫ�eI�z~`��ɟr�0QZ7/�|9�@��+ϐ�ٷ"O,����J=حh�`ʺQ���y��'�����܈��;K^�U�.�	�K?ܥx���V��)�+�=Ct��X�a{be�!e���Wk����6�H�<Q���)��Y���>le��q0��%�4��R�l{���C�'�ԩkӮ��Q`��z7�l���O��.�*3�d�1S�^;vh���ObT����b�̕#��QmV��bk->�t��� �]���Ju&�=-�R������ �P ^�􍛵�Xԡ1H�����9[O���0L	������[��㕄����i�0q�*�PL1qb�c�abX=�Y�p�w�r ҈_;u|1!�V���AK�h�"�⁫�GVh`Q�0ힶq�j0{rh:��t+�i����$F�H�L���8��I�50Xp�*ٖG��X��%E^�Vםl.E$�9's�dJ�R���aF�40IX����'7�p���*Q+��%S�\���N=a�����.�A�@��'w��v�U,r>N$���Ūl$n��O�p����7$DA[Qˀ�L��|�b(̾_NڙRP'��*���T�J�-������'��ĠQK/lc�"5#�� ������F��Q9��٧(�,��؈q�/mf�JU#�z�L1�;h�d	O6 �n�\����k�,B,�b��x�!��A�6lY1J6p��u@6�'G�������Xs�l_a��d�Q�i���6r��]@G��t�be��f�%^����I�'=��÷k��3� ��H�H���-n6d2��"���	,2V��"�B$"CV0�q�� �?1c��4lb$%�9DLhr�],)
֡1�Jk�Z1�'�f]a��MVzTS��#��3�,��.���Z�R=���I�i@��(�oG�5�$�s@��@�&���	�6���.�C�
���-�	���O����E#���xCK����̍o+I�OP,5;Y3�@6͞�Q58C�6�D���D�l�nm��͇2�d=
c�^0*��6�V�{�~���E�C�W6�M��mG3�b-C�~R�	�"}�]k���gbڐ��\X� ���A�\,���Q�@!��YK�.�A�9�=��Ǝ#*���ܴc1F	�� 9$6��E�t7O� �F�8�
��� |q�fc�"��I� ;��@-?F��F�:
�
	�wK8zޘKU�ī\[Խ��O�a'��T�1�1O�Z��$Zv�\*!��!:�̊$�ͣ!�6H�'�\�kj�gyFKuf���*�D(<`��]��y+�'���d@	�s �C�r)P���f��R#��2F3�h@7�ś��'ޥ ��vd)��dɕgv�%����9.Ȉ�2׃
$=b�x�LS�n�[b���(��	!Q�
� ���tbL����+`����ʰB�	
S� �14��7OmF0b�j�Cl^-��$�_r�'�Ҡ
�H^3������Y4�	�JD��!
�nx� P�#��a���0ud��+u��|
� �P2V��~���LR���f �'gC���'{@!��OC�g����)���ܣ=*����.
�r�b��/��!��B\��\r�ޣ7��8��D�)X��G ]`�! #I�P]J D{���=�9 ���<��W�v�J�q�ؗ"Ϡ��EVX��:@CL0-@�Q�[� Y�e�e�*t �CI�?yn1��7�I>����K	/�?-��@ڥ(`i���f�<y���8�䄋g�8q���8��A����e�Ĺ�7�:;�`�3��=m�4p&�z�*���V�2�Q>˓z����b�ۊQv���&[����0D��{��ݔ��<���x^��  ���f��e� �LjX$m��e���
�Gb苛"]L��1�p����E5�p=Q��ܩu��Pm ,i���nJ��P�ʃ��'Qd����\:8�L��x0�BåE�`S��"�$�qQpt�=A2/J9+?�y��	+'�-˒N���'Y
� �� :;��*e��ꉅȓQ���Pf�$;��:t�M�o^N	:V(�;����j�2��,���>�Pn��g�i��i�-v���Z�<� ȫ1��{C�0�.��"͙�<	��
C�Y�6&�aPcӿ(ވ��3�&��Px�K�_V�r�`B8d������<y�$��aW�j�PUk�ҬM���'�Y�L�n�����u؟0V.V�+q�L�C�<6��hcEm9�b�n��GO�=|��sK|�ց�2{U�Y�w%ӯj�2\Q�,[b�<����"�m;��&8iY�\?!�[�_�>�Ѱ�K���퓩=�M�S'D�pj:3,ƒ�B䉷~}�0bkSd��������|�O�Y�w�K�<�%>c����ak�M+��2 _z�9��)�O���\�᫒�C2=zbA�ȁ?�J���h0�<� c�;j���(�L@T9�̠��$D�4�������h�OR��r,R�E4D�̃�a��H��0'-��Q�J��9D���dC@	)0�8 �߬M�L�6!7�Op��D 9c��[��'Y�0Ǎ޿662�;�'�N����[Ѐ-�$�:i��<����̅$=�Ȣ&L!�"�lĘ��^,C:��B[�'B�I&h�pR���B"��ք�0������	�`�U�'��S�OuD*�.��>@JĉC!&j��'�3Qh
=P��u�3���P�M�`�Pg�
R=����'�9�F�B��Bn�)�Ȝ0�3"x4f�Y|PQ6D�,H��0��#�A���G5�xHf_R�կ��/��S�L;�e�p �����[�.b>�F��!u2*@����h�T
�/9D�����$2؍����c[��[�A��(��.�; � ��>E����/=�j(�G�S"n, ��C��yBoV�K���a�M�S��a[3��8��*��5�f;s�ax�ōr�B�D���L�8����p?���0��7��*��a� ��'~Fp˵,���hC���h�b��R�C	j�qۡJ�#  "?�5+WBX�����I@ԝi�H+#�D�pGN�&�yR��%������R 
|��/���
�K< ��{��i �B �i���D*.`���%q����zNU����W�<�g���y�B�%8d�)�d˔W^!kaY��y2�P3u��ł�� ���(��F��y�Kжf�bL�7��1c\��"��y��� d$(y@�$3�\xR �?�yR��D2\��B^� ͦl@��^�y�d�������/'�H�t�#�y�-_�(�\�4a��]~���'T��y��-��6����\�wf���yR&Z�vŔE�wL�+|��=A�����y�c�5G�� �%�اp������y�ꃑ1�HX٧#�0k=��F���yҌM�^#q*��*jw�Št`��y���*��h0���Y?j��Lə�yr�I?r��(�kJ�T��jׄ�
�y�W0[n� u���N��(h
��� NH)���_$�Eѹ_S�92�"O�,��a
ĸ黒��
?��lh�"OLLA٣:�����Y�A�����"O�5�ca�,[�4��%Md��r "O`�ye��
�P��H�`��	I"O:�� n��v��8�ą�x��j�"O(Y���Y��J	83�]?1i�ed"O<y���3}����LφO��%��"O ������tS�탸/��L��"O\�[E*K�)e6� JPI��m��"OD0���.hP-�7*C�r��Kw"Oj���	��*�6���y#(x�"OZ8�6lÐm/�H�h/Y|r�St"OX���U�'�ޔ�LR�6[���"O��hC~��#UJ�&q��M�a"Opٶ�<zqb��W���E�Pi�"O�@����e#<��Fh_�r���B"O܄#���h��-cm!H��ae"O@pi�J�1D⺴)�,ۆu3����Z ;��'��ۖʌ8U8ੑ�@O�~��S�'�걛-�� r�!`����A�'�d-���%[; ]r��������'�x�Y§��09�r/ uQ|-��'��I��#J�J��dC�D�@n�8�'k��㯀�b4���1`ґF\Ҕ��'��(x��Z�Ek0	� �,B� ��
�'l�9H���(c XqطD�l�,	�'ٞ�Y���8�Y`�^�M`U�	�'#����+<��2!�E�:�x0BKN�'D֝9�>I闃�
.4�ˇ��$d�%÷����_:���2�,���ȟpp�v޺n+ʸs&Gg&��aE#r?QA��38<;��N�����IX�A:�\h6F_�b��lKX��	�#hG���#A,y� ק�X���Ϩ�zDi��I>��Z��~+��������0|z#J���R#�6�,u�5ϒ97�&�2��>Iu�.y�����m\-r#jT�$8 HiU�kںd�'��� I$U��m�'�H��eZf�ì8Ŵ���,W�lIw�&�M��ضzB���J��?E�tn�,<b�	�tFI	h��0.�,+����3f� Kf��( �Ȧ��u%<�܉ C��/@�����N�=a��݈2%���d�Ϧqx�� '����@36P2YF)x}Y�m��C�0k�ea&����ݴ�0��OW�D��Wml��{ek�(b \-1D��I~�\�%�X Vd�𩒤O*�P	҂Q�(�iD��:���N ,J$u��FU❢��OǨ�{��
1D:�a��̇ h~d�d�Z<g��S���F��x�S>i����O�� ���0tBa@Nu�Tب�5�)����yVkK�`T��6f.D�82�������TA�%���:�'D��P7h@$�zuJ��T5 f9�b�!D�,�ń&kZ�35�L�E1&]��.3D��S�MNB�N��F�A�lPEf/D�DӐ�� �h@��j�����Ǉ,D��q�/Јw�@ �q��Ƙ��f!/D�4��/��~�)R&i^d���A,D���C&hG�((d�A�2�ë?D����̒Y����p��3iC�,=D�l���o82�2#<|��ܪ�g:D��;3͓�E80�[��]��HQ��#D��a���m�$�CC��l����O!D����Zתd+儇��4�B�.>D�|�t�0�L���E;o�d���d0D�x�j �[��� a��Hf�A�.D�<i�uA����@���z��.D�x�����l�a��I	U�2� �&D�`�F�E(��
���u^�	�$D��@���P���U+���� D���p��G�(�v!��8$�B�)� .HR���"Qoza�P7==Vm`"O��xpL�	�r��Q��;	.�!"O*,��܆�3�̔�-��r&"O��E����99���g�h��F"O�##� �>�4�C���I��:�"O �&؀FT�E�E��&xӎ��d"O���Bb�46˦��O�I��*#"O�XdЛF��!nߖK�>\u"O�D�c�
�K�@dO+`���W"O(���喐m	L��c� ?V�0G"O�����(WZ �D�b+B��"O�!��@��p58��<t%��"O����^���I���}ex�`E"Od$� �"s�b%9��/&d�`��"OF��d���*@�UBU"#x��z�"O,USNã[�􀙇�J����"O�MY��1?K�Y
��I�1�P�"Oja��_�=e6�ʧg\�M4]Ң"O��#�7%0���4++|�g"O"X���"��0�],,J,�#@"O� ���&=P�0a�,/����"Oj)RƤؔs�,\�vf&?{rx�ȓ'�h�Q &E8�^� `ņ�;��Յȓ9wZ����Џ�^``!lS�~�Z������3S��=�>\X�J�&�Ri�ȓ�ȍ2 �)ii�-�r��;����m:-
�,�T=�G�H:�"|��:$�\:!��:����ЎI?x�`�ȓD�$�C^�;i���� �5�攄�o�X��u'՟bٜ�c�� P:���-�I��T�dˌd��A$�N���T8H�:l�*R�bdS!��|��y��w�dYkR�M8�,�A+NI}���ȓA+2�U��_�:��MΦІȓ
���@�����!���(��ȓ_&"�����1��]*Q&S�j����O0��&X�����/s_����;��Xw�;|���tV1hP`-��¶|���x��(�ǅ�
��4�ȓl쉊���>I
6h��)u�Ć�9�K�CN��z4� �S`hu�� 4D��B��:y�q�1C��>�V�qR�?D�@���]���(7&���I��6\!���\��(0��"b�ur�)��c!�D@L<5�գG� �E���wJ!��,9�z� �d5C�0�2����v�!��jĘ�J���&��|ef@H�"O6E�%��=x{v��4��~H`���"O���3�^�j������kݤ<ے"O��ꁣ�Dm��T ι\"�E8�"O��36cE�J�����`^� m�ɺ�"OAp�$�?%b݊�L[�U�S"Ot9p�b��21�]�T�^�gBv9f"O�lZԇ�&�.y���
~@fE�"Od�ANUF��)�@El���"On�����3k�9S(ɶ"	��[&"Ou��nޫ1��-k�˒0ę�"O<m[�E�X�`�y���9��퉗"O�3v�\�`��+(ל�"O�	s!A�;0�0��D�8��-j6"OBq�K	3T�,����,W�D��"O�#�	-w\!Z����BX"O�I��a9�ި@V���f|r1ٲ"On��.�t0��r�×K���"O� �|���B(bU�cE���@�Z 3"O�ѣ��rȪ슴�J��J�R�"Op���N )=h�K���w�����"O�@��O�H(��'���gl)�t"O�)�� <}k�mD0;m��"Op�Y�X�m��A1LW�a�}z�"Oḅd� U3:���%�����B�"O���i��P�����ل7��4��"O�z�ق>���"0�9w7�,�f"OL�@�[�j]��)C%Ĕe;���T"ONAk3� Q,���Z�v��"OFܻ@Ù>k,~�'?�0��"O���f�W�HhP�u�ۓb%�"O�eQT�8ml���D�2'`�R"O�Z���=t$����ŒM��R�"OL}X4
� r��s3��'s�M
�"O��sd#T� �rxcdKG�}�#"O�����>so������xD��"OF岰�Јi�h�SE�E��ЂD"O����E�w������+mv��A"O�(!vdO�q��1zю%Ӹ��"Oʕ1���Ye�-�E.8��q�T"O�rE�W6Im8�qW�Їa��P�c"O���쀰{S8�(��2qA�"OUkB�ԝ0���G�'.~L{�"O�hB�C�f�(�G�wΡ��"O�q��-X	jX|d,)�"P�P���y���/��p lі.�J��whB&�y̑8q�n���^=&?bE�6l�3�y�M�������g�&�DX���y2* �p ��]2�4)@߷�y���[�D�Nu���*p���y�d'',�)5I¬#$J�"��۔�yB����P�E<m��������y"�S�.����d@Z�/$�ʏ��y�Ô9;h$�R���.)F�� ��yboG*�<�0u��[�@��y2C}��+�� f�X���ҥ�y��D�M?bQF�#_�����yR�[*����@��^� �¨W%�y2l�	ty	��.VubX��	��yrm�JNH`��"ԥN�v�X��y��Y&,�6��ՊPp�.��C ˝�yB�
$'>��Ս�2P����G.�y�[�k��8ӗdA�:�l�R�\��y��25������3iN����y��ӊ:��P��H�2��t�N	�y�L�VH�s"��%�r�XCB��yB������U��,�m*��U��yA�c�ڈ��� �W��y�)�:���kV�K� ��L�BR"�yR-�,�&��p�^���mJP,Q#�y"Ɵ�~f ��u��C<q�tő(�y҆"gX������1K4M�3I��y��S=}�ʩч%�#~
����A���y�B��dǔ�1��_-hd�Xc�ר�y�,�`JFd҂���^^�q뗬�y��֓zô�QkO&Y0�3�X��y�'�J�~9U�V��U�ON5�y2�E�PSv}�gG�9K򚈫��]5�y�}�tԉUb�M <�q��yb�]1LT;v�Z1@%��-�2�y2J��O�eڠ&�Tp`�@B�yB�V���s�ɪK���b�&�y
� V=Z��!YP3��O�{�P8��"O��)��rhŰ6CݵK6��J�"Oz���n�+�,�k�4cy
�"O� �s�W?v�kV&ul65� "O��k�d�>����$_�:)	&"On����1[�{�hO�G��h`�"O�xȶf�/
��	�r<�D"OP�6�ҽg�a@kT	�����"O�!ǔS9�I҇�z�Ĵq�"O� "o�Y"0����l{^a�"Ov�3�1&�H�# DjE1�"O�tA�f ;�ƈ��Q,�2�"OD���$;{<�Q3VJ��wB�d�"O��;���6?U�����D�D?d6"O�M���B�~:� s�ԍ���g"O�S��7uެԡ��Q��Xy�u"O�T��N�o���:�aW�B�2��D"O)���)l�U�DA�k�F��"Ox���ݝS�vZ`Ϝ�Xˊu��"OZ���+\&X��oA�$�VY	�"O�d�"�َ//����X C���f"O��蒀�8n����W�
ȀAB�"Oލ*�	�2��z�+N� �u#a"O@�����(G̜tbJ��;�Xxqp"O���E
ܚ;�U��N\���z�"Orp��a�za� �˗�6({�"OJM�5��P'2 Cː㤼�@"O�H� N�� .��r&��S��e"O��dP'DgB���J�.q�hU�@"O�jrϋ E��aAi� y�"O�@�'�@�J1R��"��+l�pY "O�����ڭy�	@��^ W�\��"O� %EX���Rnzh���"O�e���Ӧ(���@��ns4�G"O$0#u��!\p�hS�m���b"O`�y��y�D�?"c��Z�"O���O
�1�KX�=}F)3�"O������R�B!:7�ų3��d3�':Q�ao�T6)�d@��`5�9z�'�z�RB�P*�$G��VZL���'(0st!��}*"�B�]�pM��'�b�r�OæI�����ɮ>���'>(�;��FO�,!R-�O�xX�'���u�ݬu�p`��l�~�e�'m�3���:O��`�)-s���'�l@r��NGα�-�V�*���'sl�ëQ,bd����
z
�'O�)@$�&u��I��e�����'�T�  ��