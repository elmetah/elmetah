MPQ    �,    h�  h                                                                                 �I=A�?ej��i�n$�� ��N/a�� wE�zM��J��`tr�����R�1��͕�ZJY(׆��p[�ioRB�����U�t"�� �ݟ�@�����#.u�H�.�jJف���d
��"'�yd�F.WY(�3�VH��38@�P�����,��i�{x������C�Poq��@�rvӾ� K~,�Vфb�6m�9�zU�����⠘��a�<[~(/�RˮZu5m�������?���A�wP�z��c~�f���(������m�ep$�녗��\c(�ވ�H��9-+op�W]c��XҤ����T��v2dO���Ȧ1O�9�}Zbf��)(q�H�/��>��H ���s�/�]��$��Kl]4lOE���h�*[�����8ZŪ������c�ٻ��
[��U���T��U�{��@ * )~��+c��9BKW}^�]K%vٿ���f�}����Ϩ��ӗ�&q�lɞ�j�#��B�8�L�з������k�Y+ˠ/B�x��<z��R-���������;�V�d��nZ�Tm#���e�N��[��uc䕏f.����+ID��SB�RZ������=��k�l�`�xuuP�p^RI9�[kB������=K.ß<���
�@���8�Wu�b&�I�de2����Y>H�q7��B׏[�oX�2 �|t��g��AC�*w�o�AP� �(
��*	���qMy�򈄝.����4�E`�[pӵ�P/��b��h�<�3P�����+I��ve�C�/����AE
k�'L��?7��<�Bj��(��K 7��G���J�Q��`]��ޢ
?v��Z8�x+�:�o�%Z��I�l���W!�f=~a�����?�>���I$T����c��>�B�#� �C��k-ڠJ���a)2Ȋ8>�ȶ�jmNU�q�ǳ��Om�7S���eDIxW�+-���ۚ(p��}�����X9��)2�PIˋd̅���ꤰ��|�x��evگ`L�'�Ў��v&�?��w��[\�ٷ��bN��LƔ��g�����b�����|���zG�Z�۽��%��Ο�?ϐ������j��"y�X,=Q��ٕ� ��f�w�ǋ��V~3�:�<��^�mY����Ҡdv�fr�AM�œT�3�R�Y�jf�f���M�{�!-�1j��\`:6�b@��4���C��ǽ>�T ֮FE�C�g��5g|0�6�H�tp��#6�NW���(z��U�2,�5t*o��B�bR��mw32�S��X�pQ`V�8�s:0����2�灘ӣ�৮EV�p��"�J*Q?ĖmxL&>�|A=&�_Y�u��q�X����\��QO�a+��zz�n�8@��r
(|��
�ago�pe���x���H/�t�������]��$��J|�Z��Fb�1�`M�Xn��ڶ'x�6x�4�* '���_dCR��jŽ�P̰�'D�P�9�t�H+��-f:^��� ��k��A��k�\��2��a4TF���#	�Y%�5����Z�f�C��H����]4,�:�*]S��j�����/�Cu*��� D{�a��6:���:(]k�8���k���G�[�,���V�����֌r��`r��������&���������x�2��??M0��V��d/�v���*��^�CNA��3�fnn]�նR0����ڹ"�Ֆ*�d8�Eb��zOn����`��kR�
��"�]���p��-rW&d%-����btЍ��N�(��w�f�#�ew��F�t��߀ܰ,�^�n6�9H٭�r�<e�:�0R�j�C��,xc��t��2�pa0gH4��Jw��G J�dL����&-��vČ������SO,�L��\im��9t;6*�#iX�m��c���v�*��l<�_�{�;����fH�	� ��"�}��j:�q�s�������Ed�X��q��y'�ק��Ӈ4?���Y��>�A"]�����N�M�����Dj��7���&ub�� �j�U����ŭ��=Ih�X8�����nT�0d�"���G�"6>�I��dcuq����(5��0��)�-��ڊi~�F��#C�	��:�Z�n�<�����%�Ȫ�!�&�0���@�lF�+8W�{�Cwײ�V����e�<_��E���\���h���h�m.��ݧ�烬>�`�l\�ثs���#�F?]1���t�������⃓�߫}S�0�Jl~g����v!����	0Z�#:u幡t��lrŒ�X�%�#VW��#�9���3�.�J9��D�n���5F��)���*�C^ �=���2��+�WC��s�V�8�����]�Xn�3�j���ǻL�J���bK���q��� �s]U���	D���NX�AgZ�,���é�&5��	�6��)����{8=�P�_���.�il�I���F��y�l�'$�"��:F��|���o�;YK��w�y,WXFg�0���26����c�}����3Z ^*��{�hU�9��B7BT�P�D�:�����Q�Om7WE��F���I*<T%;G�t#���r(�j0�7I{��
��u�>��Y3��he����f~��{@7�m� �\��+�Pt����h��)o�Eq���`��7�S�e,���+���ɊJ��b�t�GN������o1�SZ@�ډ�?�NV܃e!���+Z�@���`�$�Lq���T������Ȭ�龪,�%�fP��� 1t�<t�"���C/�R�mlm�	��	_����.�S�~�cXI���!���9�+L�$J+٦H@x�DRU�����b���L����!��n�%�1����]�d�����������G�EM�� .��9�n"H̆���;�D�Q��fK,R�Qa!�*�~D6�����N"�\�t�Zt��r�楴�fܧjM>����3�ǐG�Mh޶Bje>�P�Z�I�x�eF+���8����ʡao)��>�|���ŮVH�:����O 4�M�2��bJ�7�rݲ���[8MM�
��h�I�@���B��^�|��8�%����2�g�xMe���G	>Z��T���cb.To(a�b}
�n!�/
�W�"��d ��W�!�3�������@��q��}�}�ui9�x�e@���֎��P*T��[�E�P���w,����V�h�c9P8�UteS����a��<�X<�Q�/E��Y6ZЂ�u�@��������?�AV�P[ ^�^׫f�a(Dd�������Ε�Ƴ49�T\�8*ރ�� -�}+�rC��c]�c�4�n��{e(2��>����ʴ�}5�!�U(���*�>$ň fs�R��O���S�܆v�4�϶�m=�+�`���'�9�������p����]}��@ 
�h�+D����\l�U� ��>� �'!~���s�؏��Kr���k�v��o�ܑ�'$�ӵ"�,yN���l��j�\��(ć���g��{�������|x�4:z}�-�'�;�؅�GV�����U�����#���GN�$�:�1�0c�fu���εk�D�ӑBk�UZx�N�=������k�纻n�x���P ��R���6�Ρ\��N�.�|;�(n����S�}W��-&�{�d���Q�>CC,q�����i�v��ӬI2۠�t�gggQp)C��N��YP�>|(%o>*������y):q��}�7�����`=��Д�/R#�ԛr<�O�z]���GIQ�e�?��J;�BP�
F��L���?҇�7��j�T(��� R�%L�P���9QGmk`��ޝ�v�6�8��U�(���b��.l�KA��l�!G=96 �'ʺv⸧$�J�[�,��s�B �� ���؆q��Nk�~�)m��8�C[��jMNu5ٱQ���\�O���2�6D�O��&�1��F�������:��30�d���`ˆ�'�;أ�@�ù���)eQe2�2v!���&����2jk[w���\�=��ć��%n���ѽK{���|��=z¬�����B!ǄR��:�W�U�5��r����('=,L����貗%f�9b�z������3�{���^p�8����m��v����y��NпT��RR�jA�ܬ(��%�{�y�ʌ�c���e`U�Sb��Gg�l�����>�w��	ɕ�����^�g�X�6��t�A�̾��NR�S��'��;�,��*��B�E>���w�7kS�Tɢ���`�9�8���:�O���MU�T0���C��dS��Y�pp9��ep{??����LIz��&�k�Yr��uھ����o��\1oO[*+��lz��8�ur�����옟a�ىp�����v�?�H����U�r�8͹$�}|xw[�AD1ic�M�����q��1]��] 4
��'80Z�)Ra�J%�.�k�Fꢂ����9��mH��(��^�� l���	 ��g���m�����T�w5��^	h!�%�qҴ���Dʼ.�U�����5��*����V1��ص�ª�u�=V;� ߮X�\6�6�[9��y�k����FҖ�)��R�,R�%�Q,V�n���g���.�ފ�WE�o�*�������&����G�ML~����M����#����?v�ϽL�ЇQoCi�.���nI����<����ϛ�}���Q�<dS��bY�z*VL�3�P���>���}5��Ґ�p�$r�I%���)QE�(�N���
e�!��>��w
F�VY����KM^��摔���C��<��=:!�R�۱�Qg�k�c�課��p�HOwnJ���"�m��[�Y�k&(�p��ͼ��3����O�{'�-\��v��Ձ6%<6i��҅=##��l�*���lw0�_LH;�t�c�HnT	 �;n"c��E�pqہ��G��{�t���KXmnC��D�'F���4z3��e�8�4�A���]?����ƃ��P��ÊD��\75����b�� ȗn�p�{�I�r�pv�I�g*X�d\�תrnw_0�ǣ�F���G�$D�Xt\d�X%�$J	�c5I���6�¨&�eU�ۭ�&r����:i#��)<6�8ҁ(���A/!1�0�Ʈ;w)FV���nc{�R��-�g�� G�=�<����@�u�?�[�؜��՚���H
�0��<�����N�Гٕ��e����q]����pm	V���=����dcS� ���?<~BA��+[H��It�~r��t�t؜�r�㶊3���^����q�4���
���_b��	Z�5!�L�dK�����^�(�+�s�ds]+����e(�V�=�!�����?nЭ���p8���=L5H�Jx�jb&�����(2>sX���-�S�_[X�ZYw�lk��
��&�6��W�"#��63/��_$6.���l*_ı�~F�i�y�ӕ��?$�M"x��:!��|�	o9�K�x��ԑ�Xx�0��]2���徶����K�����!#h<��ǚ7���++)D%<؜r��Qk��m�}[�E���B$�T`+,GR��#��Qr��p0���t�
����Yn�h ��榦t~(�C@�%8�!�u�F��K3s�t;3��cF�)��E,��{��ҏA��.͗,�s D��1�J:yL_�b)��xb�|9w1,�U@y�:�V7V܈��F���4yŶ��Y�HgL�_�O��1�vn�>��i��T��AC>4W���F`�7=`"��L�7t�7�5��:`m�<	������ֲS.Ng���
cs�?���*�[�e�f��$�;�C�ٟ������}���b��\ܩl���
0���(����XDx�)��`��EZ�Ὶb����nz�m`A���;�[����f&v��������~?�����	�t\
w�Z��rۦ�'����O�רCҎ̝�
�h��<j��Jճy��Q���vF&��ޓ�G��w��yo��>��|��KԮ2�VC4����եc��4�2�iJ�-ތ��Fm�[39)�eh5h� l@�*BhY��W���s�_��T8ڕ̶ª�xӮH�)�3G����S!T�yլ��.O�a$N}��	<,(
W_�"ݣ�d;�W�;Z3�И�D�@n ۇ=�.h��CiY�xM�$���K��+P�V��v<�l�����,.���F�c�9�z0U/�6��a��I���<�D/����Z+�0�G�� v�糥u�AGT�P����YPof8��(������[Mơbt�+\�i��~H�Ba�-�����Iź�&��Z\7o��9
�vt|2���:{����/5}��=�U(����%��>ި !Z>s(���S���������#4�Ҷ����o%�ʔB{�.�����F�O�ߙ:����
ز�˅���¢�a�U��P�:\ `o�~���?��J��K��w�S�av�?|�ݍ�ك�λx��>eݜ2l��oj���Ĉ���R�vT���ڠ��x��?z�S�-^�M�@��� -�V�|&�$q0�|A�#�y�[�;N�p��u.���Vtf�x�6ei�&/�D�B�`�ZS׋�xm��s%ck�����x��hP��R?���K�N޵��V.�y�ƃ
���;�n�pWkׄ&��d�,(��!h>>�q�{|����KN�L2��&t6 tg��C�0�%LPq|@(@d�*��P�ˠ8yd�C���������`��;��t�/�5����<IpÔ�k��_I�1eR�K�e��~�
!�wL�_�?mh�2��j<�$(c{G mAq���|KQ�1�`�j�ޘhvY��8B,Ыp�������k���lF�����!s�a=�*��B���5�Zⓦ�$�$��m���B[� ]#�ء�aږ��Y�)�rR8tЅ����N�65��U��W���z$��ܘ�<&>DG=�!�_�AP1�{R�'���������{���ˁW}�P�^A���nٴe,%�8�]\j���?&O`l��r[�܉������3���8�:��}>��
�OD|Ьz=~В���}=���ģ5�Z򰌛�hΖ�#���NE�=�����M��f�����O�3/�A�2lu^K��P��t�v���Ş�	�nT	�(R͞�j��c�j����{����81�z�`p�\b6�g�-�I���FF�>��T�dk&���m��gr�J6�؃t攈�Y��NM� ����˳,6�*e��B�H��Q
]wi]�S�-6�&��`�=�8�I�:&.���������GԶ���|�p+�����?���	^L��&�ڝY�;.u����l!�J�s\G�`O�K+�(�zmA8�7"�T�g��G8a�c8pP�)�������>H�5��5�J
}��'�$*��|�t�<�1�2�Mg����ڬ�h��a�4EK_'ӼUz�R��@�0�膦��#���93�uHa�#�^A�y 'd)���*�aS��f�o�׀�T|�|��P�	�q%A͙�,~��\�Qʗ4�Ks�����0�a**~����s��%�ru�k��  z�W�/6�j���#k�jv���:���|ԍ�,�t��L���ɐ��"��Iz��o��J�L�X�[�\Ԩ���r���Khw�h˞�5��M�s��i��8pv�� �CZ�BdC��}�)�3n$���K�Zf������'�F�dn�b��{z^/�nʔ�-!� j^�ز����p�DrM��%�?+�d_���T�Nט��eݨ�e�Y*�w��F��΄�.��G^|�������Ϸ<�ؖ:���R�䨔�)?�d�c��G�pף�Hjx�Jm1���ga�ڊ����&#y#�,�̀~���5�kO��V�\��M�oW@6 ��i8��3�jxlp*��7l�u�_�4;������H)�n ���"�h� �<qX+Ā-�.�v0����LX(dY��Z'�X��|s�4��8� ���J�A5�4]�v��_��C�
f΢D�Fv7�+�Ȑb=�� �����m���,�K,�I���Xn����VanҊ�0ڐ���y&������d�\���d_5�8�QM6�#���@a�5~����M:Ĥ�����(_���ﰅ~��!l+0��D�6�bF�d���{��]ר������x�<:�*�;{��������k�-o�#(��S����}��2SQh�N'���j��<p�]�����l$醢P�����U=�S��)�@3_~�*�f��]������ʯ�/I�t�w�r�!��̙�6����/�x��q���,�z(���D5�\�џy�`�^TO��0t��s+��Ƈ���V����\���i~n�Gš JC�Q��LP��J�eb�B����c;sS���c�:�kX/0$Z��#G%u�E���"6�&"�}R���ME�_��=.[�lZ**�LϩF�d]yoߕ{R�$��e"�:��t|=��o� �K>m�/�X���0��2,�qH���M�*��`�|�h��F���78aQ�bD`]>�cD{pJQƈmm���!c���r��+T�W�G�S�#���rޓ60F���}$
��-��پY�;�h���桘�~��@���<��+�޸��n��tּ��^�)%x!E�GԖ� �
��	��,l��Q�J� dؾm�}�_��ؕW��1g�@z�5h_V�Ȇ��ًab���¶s���L�t��J�i�gu)|�
.�"�x�V�oŖ�6|D�2&�"T��qK=�R!�c)�m�^7	-Z��J��f).������c���w�_�6BB̡4$�"զ>����+�r񠄘(��B粚7)J����g���~Ѥ�
$��.�/uH����E5����4����nu,<��ȂY�;ÒؗG�f��ǋ��`^�~:��q�O�ė;\%��Zji�rZ�״b�O�����SD��ֳ��_�h��j[N�s��YȮ�_F!Q������X� r�o՜>ԁ|�g6�I�=V>uo��%3��4��T2�}J�CZ��_�e}[.E!���.ho�@_�B���2P̑�yM�G���l��a*x�0��DK�G��+���T+a��:�s.J�iawq}�׈WЈ
҆,"���dv�hW*uU3�=����G@)���"s��ͽ؇i�zx莡��]�Tc:P�y Ñ���r�1�,i݄3V�^�]9��U�^����R����<Xv/{b���Z�}��ٲ��pH�
;ХP��A�r8P��+�T�.f�mF(�ˍ��K����|o�
�\4���y���D�-\����o2�Y
�5u������|�q�2u�����pʪO�}�M	x.*(BU� z>�� ܾEsC����.�o����t4=�L���Z�;Ԋ�~ܔ]bQ��Y���,�O�C�47���@+
lgxȆ �k)�Rw�U�j��u�8 ��9~�a�)���K�T����vj�شRHxN�������#��W�Wl75j�e���X���N��qE�j���`5�x;MzJn-9��{�ػ�>V�8���D�7�S#���\Nm�Č����fj|f�b����ĵ�`UD߅�Ba�@Z.󘜳1��&k�H�qq xBK�P6�R�_��_��������.�����ƚ�qNm��%�W��g&x?Ld�]��vS>9�;qHc��s�r���g�2���tq��g�� C��1��^SP,�H([y�*zP�ݦh�y��j�U�����E�`��7�u/�8i��au<�>���hM}*tI��e���;�8�C
���L79k?i�-��j�[�(z; ��B��iEQ��`.�4ޓGYv���8��ȫ�~�s;֥ߎ��l�ؾ�Ƞ!��\=�?��]>Yʰ�
�nś$��'��=�B� � ��ؼ��#R�4�k)�w�8}H����N+vUO�}���E@��Q/�w6�D_D��I���\Y1�Be6�0����8^����!FT�|-���>�M���I���4,eۇ_z�I���4�&� ����[�n�u8)��O5���h[�x���s9�
tP|/�Cz�oM�l�5ԸygǺ�+�0�����#��>��Ɂ+=��p�Fc����qf�6�0+4�
=33J�o���c^&rǜ�b?��fv�m��R2��ğ!T$�:RHqj��`����[��{�(�B��5��`�db��3��|�����>��ֿ-��t�V���g�	�6aPTt!h��e�NHЉ�9☝�L�,!�*�UB�kf����w�3S�&���i`Oa8��:�,p��J��"��������V�p�v��\H?5K���L��l�M47&�i�Y(�YuP�&e-��c%�\�O&O�H�+|�ez���8q��='��TŢ�a�p��!�����z�H`���P:�����$ej|�&�7�a1"qM"���2��'(��ǆ�4�M'n��P5+R�v�������㜝�_9nv�H�L���^��e �T���=��^��ACe�W�T��ֻ��	�%�H�Gqs��Ek�rZ�TS�.��+��*n����J�R� ?Lu�<���� v��R�6K�Z�k}-k�3��<�����8,�S��Gp��$�6�����d.����/�%�^�²��� ��
 ����jG��f�M�EP�1P�5�8v�?��"����C�u���n�s������z���Q�3�a���d���bO�z��b���,�ȫ���G��3P��H�p ��r��V%�
���C�^J�N�Am���O��9�tu wG&Fj2ԄL+�܁�^wj��J�ݭ�.�<�:��R�P��mˇ�/c�F˲�-p���H��J�u!��;%��è�%$&�2��@��9���P��O�z ���\�
�v6��ii����G�a�J"*n�l���_�A�;딯�;�H�I� �;"�1��X8q��:��s�q�_�Vc�X�y��5��'���W�4�	͌���ǀ6A���]�G�'꾧{A�*D�7kyR�ɘb�� >�����?��&"IjYX	�k��"ln-�*0�G��"C����\��%�Ό�d4�5�z2_��5�c�lƨ?K���Q�\o	��}.:F������C���w��Y�!��0R�:�1�F1HO��{ќ�#.�e��< <�,b�6s!���$�d�������t��TD�H�T�1�I`�sN�	���菳��8�]�X[�<���^T���i���6[S���Fn~�&���*~?���ڜ�4C��̬ts+rv�#�����Ա�U�o�*�e�D1�{������5�5�������u^C����4�چN+k�[�xV�%|�����.Pn�9�{C.���Lk��JnY�b��p�"��^��sN����t����XJ��ZOl#"�e���\ߢ6�v��ءѐ��&�E_��.6�l�J)����F��y�{*�6q$�'y"n�':��[|xPoo�(Kz$2���[Xw�\0�62�n��tLc�.�Ð��(̦׌�h���:Mc7���,D��8��ˆv��Q!��mh+t�<���ut<�\T֣*G�'T#�;�r9��0��̦�
,��ϵVY�$h6��未�~�Wt@h�x�W�mk�#ޓ9��2tqf��Y�)���E��|Ա��҅�T��,,<�'�	���a�J���Q������n<��2�1�\�@��ؾ0ہV��R�d�|7��*J��N����M�LB_��E���d��$X�.�A��������S!��� �-/2"�]�,��m���7&m�<�	h� 0i��:.��CZ�c��4��C�������1$N��9�
�Um7�-;�������'�]S��8�#�y;}�u�	���ɐJ�=�V�sE���5��ފnpap#��=�;�陗�H�f�i|�Q����7~5֪�̥���&\@��Z���r5%9��wק;t����D
�x��h/ވj�O�S���^�I� F���I$ �?Y��>o��>��|0N���myV9� �K��ْ4���2}�J`yf�#Q�|~n[)q5���h*.f@MfB^���1���u��;��c��x7{xI�[�_$�Gz��K�Tfh��΀.EUa�t};�r�Q
M�"��d�ϹW���3��ق�$�@�o�Ǝ�3�͘��i�0kx�S���o
����P[�cìP�b���l��,�7I�΅�Y�t9a_�U�n��L��z0��%z<G�8/����Z�*��2����إ+��A��+P,ц�O��f�Ey(u���f�Q�2�W�l�S�\�*��t0z�G�-j5�õǺ�H�����o�-�l��2�H��o��6�%��}�15���(�L	���>5q� �C1s^�.�I���J���7U�4�U?�����X����xi)�$D�["#���S����
�^�A���]8�ͬ�UiOH�_I �^Z~��/��e���K�1��I��vE?���Ӷ�ˎ�'��=)��tl5��j|�̂���86�8�ΓlV���,�q�x4�bz}`:-y[ɶ���V��V�<�����#0��Q�NHr���f����f�	ʙ�Q൜��D��Bܙ(Z	/v���BBk�����"�x�'�PQ��R5W��F��B���B.�� �9�u�,������Wa<�&SѣdQ���"��>4�-q�j.��0�D�W2l��t��)g"�0C��=�ې�P�W�(v�z*�(J݁Pdyڃ��{��e��>V`n���!�d/y\��e��<�,�K'x��Ib�eȚd�����;
�Lr2�?���(�j�H(٘� ���m�D.Q�\`�a�ގF�vr]8�_���_�w�րs�5�l|���j�!)�7=jt(�x
�+'�IB$@9�,jX���\B5� ӂ���6�ڌ��x�)�j8�I���*�N�Օ
2ʃ3|���%������f<D������D�Ȥ]򭢫����x��=���w#8���ԭm��]�d��e��ZL���W䎎��&R�c�[ȂZ���������8K-��s6������ |JLz3���G��՚�U�ʣ+k�f٧�ޱ,�YG��D�=���ف���#�f�?����,���73e�(��^	w�����>�Vv�Z��������T?��R�c�j�5��ٛ����{�A_ʝ�,��&G`�^fb,߫��������|E'>�����/��
��gh��6<�tt\��̏`INC利A�,<�"*[)Be����&rw��S�?��=q`
�"8���:K_튷��˘}U*ʰ���#p�Em��?�|BwL�6��o�&��Y�8Eul�A�5�i~ �\��OP�+w�kz#��8,�lX�?���}:aS�qp����Y�P_�H���k�� �x��:|$�?�|I�o�2��1z1M݃��M�ڢ�	��{4��n'	l!KFRr"�V� ���R�xO�9�a�H����>p^�Z� �ew�("9�W�T����MM�T�P�ֶ�	yr�%�䴴b�6�R���M���U�����&�*ɀ��Ek�)P�Ru{-g D �	��M�S6���&/�k�6Ƿ��w�����,#RȮBBL�����&ӌ�
�F� a����ג���
�w(GP���☞)x�+	�M�7��lKK����v��[]�
и��C�)���n�Ǭ��2�)Ȇ�G��,�Ղ�d��b��z����0�cV��E�ڎD�kOp%wrCt�%�Y���p��_qN�
'��B�R-��nw�BFE�i���-�o^r�����t�t�<�d�:��wR~V����<[cꥵ��kOpM��H���Jc����/��PI֨*|�&���⩍�����k�#O*��s@\U�ش��%6�Vi�&�n"_y(bE�*IK$l(`'_n�;�T�t�|H��� -�"�����Mdq�+�c�o�l&MX��Q�P�\'�Y��2��4+���6���ֲA��]p�0�B�0�9��D#DVs7���b�P �����0���ĭ�8ITOX�����n�A/0P��=��<�εƋ	I�d�Ñ�u�C!�5zgQć_c��X��ز����Q���k:z��Z�{�^G*����4�]!�0��,�HFg�
v�{2@dמi�@�5��t<p�1�1���P���gޜ�a��H&�١)�Ɉ��瞧�	,J	�t��"���s�2!h]oPA�w�b>�����Nyd��NmS/1�6zi~��}�ܯ���S�ɏ���p=t)��r��k��6&��f��%�%o��4�64]��>�zVz5�.��(���3�^RQ�<��@�+4\j���Vn�2�Ң��Vn����\���L�|�J鸝b�/��]���&�sI)Z�>[���n�Xe�Z����f��;=����6���3"�g��AYo_~�Q.=klЊ\Ă>(F���y%����o$��T"�w:�$�|�fqo
FsKu*Ӛ�X2jW0"
2"���OG�iT��`�]⤦2}{hA�d�U��7.�B���D��ƜCT�q��Q|�m#�v�W�1������T8G##���r� 0�����
������Y
�h�V����~9��@#��r)��z��n�(��t0��T��)ې,E]ϵ���T� �v�b�,wf�D>6��)�JKoN�����ȕЮ1��@J�c�+n`VH���3��,���!�)@C���4L�i�@Q4B������I�=��|���J� �lG��(X�"
f%���[����Yf�mx:�	��{�I֖�.)._a���8/c�a�m�N��s��$����4|^ٰ��[��J��8P��,�Zz<ϝΠ�tű��|ϸ��H�em���łE눰�pɸ�S �nk� ~�q��8';�`�=�Ff� �=6���WM~0�q�'Ņ�:�5\[=�Z`��rzʴ�g���kՃ�	zҟK��3k3hJ+�jQ@�fS׹F���T�F��ޤ����y�6­o,]>���|kTh�;�V4WΉ�Fn��>.4��2��J;��^b��w[$�e�vjh�d�@7[@B�m���1H�$�E�}���z��-�x���z�G��-e��T��y�p��.@7a-(W}�P3�x�
�5["nH�d��W`H�3�w4�Uq�@�G@,��i�o�s�Ai
npx8c���S�
2P���
$݆��Gk,��i�ST.H9�#U`\z�1��Ò��}%<��N/������Z<��a���(q�� Bͥ�JA��P����J{�fI>,(0�-�"��̈��2�J%�)\j���oԌSk�-�������OC���5 �O
��ga�2+���*(��-��ʠ9}�51�O(x���U>��I R� sy���čI�%O`�r��4s'����h���UL�������NE�6|)�Ů��j������
"�c��Uj�:o�HWUDT���� 13~�w���{VZK�.z��-�v �~I���������N���D+lP�xj�|��uI�s���)�g�� }���̬xO��z��-�~:�����V���5�M���w#KT?� !N##&�&3t��4f��L�G���W$2D�[BWf\Z�#�)��D�k�Lm�'��x�$Pl�R�n��Mb��$�����.�0Ɣ�P��=���{Wܞ�&.�d�����>/#�q������⚂��_2GT�t��g���C���6�P��%(�*p!y�\Xry����r*�o����`)�[�<խ/��_�@�8<�:ה���s�I���e�N���'��.��
�i�L�K/?>��#5�jM�I(�� �#E8Gc�7�Q3>�`d�މe�vjp�8s)��`����['�p�
l��T�!���=%�H̓�Fʦt��$c�${s^���Ƈ6Bl�� �b��.�xi��m)Y�8E6�����N�T�Ŝ:�N>c�;+®~����	DP�z�dR�R�s���x��&:+�����P���W���r9�p�؏.��/Z��K�e�Н�O.����O&`��ٞ[�O�k�&�����s����w�n���)9w퀁U|e��z��˒"b|�.R��𠡣&����/N��ӝ�t����Z`=��@ټQO��f��z����v 3�O��b�^ܿ�gx�٠�v�g-�k��:�TZ��R>v\j��%�9R��dn{�2��^Z���/`�xgb�<�{ڬ��L?��>�CV�uY���%�kg�:�6��t�N#�*{�N>�0������,W�*��B@O��w:��S�xe�7��`��8{�:��Z�eŀ�@���F�Ŵ���p\4���ȵ?+fZ�L5���K&��>Y���u��\��v>��f�\��-O��+r��z~m�8���s?���r�X�a���p!z��lG��coHքջ�([{\���$�4|�)Q�-�1�`�M����hz��s��}0�4���'�s7FR�|���]o��ԝS_B9�l�H2��^R�^ X���Cj��ՠ������c=TM.$ֱ�#	�"m%r��}���R��(G�v��d_��!oH*$\;�B�0�Dn|�uV>�B,t K�ޞH@6�|�� �k&�2
>�RY��>/�,�pY�=4�����S�������uʢ�S�	'=�-��Z�����|���1����MaI駘Z�k��v�/s�y�s\�C��\����n��)��/�7�͆�[������=��d��LbEspz�5���Y�� a��c|���혾�4p6�r�@%t�JД�@N����vƵ�A��k�w
jF �����
ܷ�^m��� 	��/L$<�ڒ:�wRY���=V ��&�c�$ܲX�Ep��H�;�J�^���C��ؼ���<&�d�=3>��F~�%O����2|\�0��@�L6�Yi�h�)b{!���_�*$��lc�_���;�4Ǌ�ْHZ�w H�"9dձb�q	�À�e$�g�:�X�XY4�k��'
��S�4f`���x�LAF�I]+�~�]�:�~!���D�9{7�t��+�bN�' ����ܶ��5>����I���X?�����n���0ǣX�~���Mΐ��D%dj'&�p�du��55�Ģfز��DHǊ������:�����y���m-�ݢ!��0�'k�F�)��={Mϳ��$�h��)�<V��,�=�1�G�(����|���?���犺��/�d���Ǩ:���)�]Jhw���[�3���Z��I����SJ�)���P~��O�����^�����H�`4RtD�}rl������J�\��vΛ k������k��:��?W5�G�P\��1�^�,�����PP+Om(�Q:-VI����t�d}Kn��4�1����.L�x�Jd8�b�����˗��sD�q���k^�X���ZE���x���q����6�v)Ύ���"^`\+A_��].��l����{F�jy�Ё���$��"dn�:��|���o��KpPP�@g?X���0=��2���*b遤���'��y����h��9�pSL7�����oD����SlDMQ���m�X�r}��k����TL��G�.#�)?r�f	0w�Y�
�$}����YZ��hlՠ�.E~�Z%@�XJ��}jaR��I��<_t���O�)6M�E���;�{%�� ,��ߒ���J�V=	�q����d�B���v1�K@�X��&!�V����?G��A� �����4��Lx���;�c���Z��d�!����­N/ В����#��"e�m�F���t�ԴmSX�	ޅ�fJ���BS.����7.c�7ʿ�V��<��R��$Q��/[��ʎ��._��*��4���$�ܕi�8�v�ooB�+fu�D׫��a�L��EƧ��ý��A[nf+M��,ȳ�D;����Kf�ݓ�x;��1�~+6ձ�Q���h\v�dZ�Y�r�x��q�ǃ�����v�� �he��j�P"AsA���f��+Fs0��.y���Qo���>e�u|�z��)�V/�w�L�O
�4]*2��JE/������[)���U�h���@R�BBT_��R��_�O��.Ʊ��.D]x�u�6CGp,�@ëT�֭��.;9~a�i}��^�|
C�"I��d'T8W��3�D���X@Z?�G� 上�N޶iEˉx�<���9�eɣPѡ����?X�3�"8�,轄E�O��9ĞUjn�L� �+���� <�Q�/L�����Z���DM�C!0�{����AA3�nPb<%�EtVf�V_(��Û7��G���y�`FQ\l��j����-��p���j�ʌH���[$���7�b�%2����as�H����}|Y�)��(:z�(K>�� ��s�W�?m� ܭ�!4�����L��+���q�y6��?� d��홻ް�
}Չȷ0N�U�N��w�Uy �&� ���~�2�:���6�^K�K�?�kv��δJ0�s��j��݈5�lk��jr�^�d�iĮ�!�n�+�b؛�{����Hxj��zs��-ʤ��,a�،�fV�,��B�h��#f2�G��N��^�a��7e�f����W��FD0�B�R�Z���d�;��߁k������9xsA P��BR+�}t��:'��U.��{��+����ڢ�WW!Z&	U�dǡw�X4�>*k�qYو��'��$�:p2"ѻt"��gX�xC�����U�P]��(�x�*�9t�7��yP�׈&���M{�VY`�/��W5�/o��zB<5i����nřI|�e>"���r7�x�
���L�o?�*5��j���(O6� �Y1�@ֵ�_sQn��`�؋ބ��vŎ�8.K�܁�����6����l���^!�>�=�=M̮��!����^$�ʹb�#��\�B��� Ib&�-ڂRG�ū)�G�8�B!��J�N<�v�'σi �߶P��Yp�('D�e���p���_�N��l����,�zX�������mo�e�J�*�J��Ze��Pg��>��ע&�!8���[��K��뷆�q�ĮMr,]��i�;ф���;8N|�H�z)͒���i�ǋİ�!y�����Tӈ�p�:��=s�`���t� �f���A���;C�3��j�J�^����<�t��v͔-�c7���FSTu.�R��Pj���O��,ɐ{���SV��f�<`ܲb"��V��5%��Ĭ>����4꘥z�@��g^�6�w�t�!��ŵN9N�Jj杷֪,r��*Q0�B�k�=�Ww�3%S��¢�`���81v�:�a�@�s�{~阳V���R�gJ�pCk�쮨?���5�PLp��G*&���Y9�\u��wx�2����\3�oO��B+mP�z�f8��2���
��3C�a��{p�n�����*H�4����p���Σ$J�|���(b�10��MS��܃�ژH[�X��41O'?�A&�R(��̇b�����	�"�.�T9��Hͤu��^��k �U�^���MAپ�s��Ù>T�+L֬TK	/�%-|ഘ
ղH	 ��;7�&������"*We����_����u1o�}xX �L�CYh6\ۭ����k#OǭVז-5��y�,Y�B�8F�50� *��
O� ���6�D�p�ȺV� 7%���7�^��r�!�,M<{���~��#v�&!<�.�9C��L���n����7�������e�D������dڤ�b��zq�ܼZ���>�D���y�~pQ��r9ۖ%OKG�P�'�/�N������t@�$w��F�kE���|�R�I^h���[\���
�<q�:�=�R4Hf�x���rR�c��>��H�p�
Hּ*JY��iwQ�Ƈw�`�M&a����΀j$�|O��n�\��3�۝�6�iz�΅���<�X��*�>Ql���_S'!;�4=�*��H�m cF]"��Ռ�LqD�ր�=��b�B�g��X{Zˆ�~'}�R��2�4�;��l	%��?A�B]�0�x�,�/�V�9dD�e7<"����b�1� o@���|������CI���Xڟ�־F5n>x0�+��s����kh�!4d���k��Э�5��zĽ���XڬЭ��-����c�:0�L���sД�)��Mم��!X��0#H�"�FVY���{h~�הn��I%�d4X<���'6���͖�
vU��⍲����?���%���QR����:�>�9�L�(R^]%����ǨtΦ��H
���A�Se�N�,A$~�o��RIO�를�El&��t_$3r�[!�z2�̅-�&硛���U�x������pI`5h�>ы���ʠ^�C��)��w+j�.�̎�V$q�HA�����n�Ａ��/�=%L���J�׆bm-��ӆ��/j�s?���C��&n�X���Z��j�L��1��-��6~&d��O#���w�_t�.��lFk_ĸ-�F���y۪��g):$!_d"��y:h$�|)]�o@�Kk����l�X��x0Xz�2qQ��T��`ߐ����J���h�&�ۋ�7$�drh�DL"��y��g 1Q26*m�h��Q��8�k��T�HoGYb-#���rJ��02BW�y
x�/�`	�Y�X�ht�捠~�N@�5�����I�$�HZ��tB#��J7�)�)8E�~4�b���M_�uf�,��iz{���J^����[d�߄i��)o1S�K@�8��!�QV��������vK�s������o��L߹�6mo�2�l����0�[�y�����
P"�V6�]ڊ�� �O#�m.��	-k�v�.��tV�c�-ѿc%�̍��$�n�*Z��f���^�&���.9N���O��x��ӛ��j9/��o����厒�D�E��b��ݶ���wna��4&��n�f;/��3��fm�7��`����@~&�Ա�c<Ͱ�\�a�ZV?�rƃ}�N����q��?��U@�����h�%�jG�V����9i�zuFi��Z䵠p�l�Do�>@ms|��jԵ6�V*��\穥
��4&��2�pCJ������M��[��,aVh[2�@m�lB�p�������*�����S��z�xzw7�o�G�`�VT>���Z�.6[=a�ʽ}lJnà
�d:"$V�db�eW���3~1^�j	@W�b�_�1�) <i�H�xTa��|7����\P�Df�����v��$8,UpƄ���J#9r�ZU֗��g�^�����^�l<��w/�I�LrZ����H�^����z���An+�P��h�@�f��(�ޛRxv�¥<��f���\�<��e|	�-Hv�Hx�E�
ҡ��ؠ@���]��2�_���c��ʖa�}W��dk�(��6���>F=k ȑLs�ӳϺl%�����SC4�*趉+g駥!�}M��>⒕ó��f�;9�ߠiλ���
����r+V�p�U�>�U��$�a�� g�~�-�#	��A�K�d����v֮k�>5k�6����N�x�CF�l�]j��?����ŷ	�N�]I��}ĠL��x���z�c�-���gb��'�NV�h����ְ#�+#�0y�c�N��G��+�����f�������gDKj�BM_�Z���<�zޥk��X���Wx.~�P��*R���X�̡uI[����.�Jc�J��]�_��a*W��m&�Fd�����>%Ӭq�@�_z����]s2�mt]��g��C}�ɒ���P�(��*fr;��~y��N����KО�`���r��/���l�<p�Ӕ��i��IsdEe�������$G�
h��L#�C?t��=!j�-(
�t ��E.Zu�ը�Q��`�����v ��8�T��¬
E<���|qlMs��!:�	=��5��.�ʜ��ڀ�$�G��N��Q^B"� �I�(���L�����)�̥8{oD�{
\N��;҇��"W�1�2�4ej�c�@D����ZK���EH���YŢ;��U�{�Ʈt��h��I{����e�K���BesFt�7�d@`���&bk�PQ[lP�aU�_g������5��d�����5���|��1z�u��؃�Ԥ�m�&��0��w<۰ẅ�������=N3Q�2�n�T�+f�e/��pV��/�3�79��QW^��&�w����v�ᩩ�#�Ű�T���R4��jc�*������MK{�)�ʮm�!�m`�bb�W1T��p�>�M�>���+w��`�[�g��46�o�t/�`LN4�G����r��,��*�c�B�6��x�xwp�eS�J��`;0i8L��:�fu�A����֘N�������p�q����?!y1�EL�����@&���Y���u<9��i lG����\n�O!�+h*�z4��8]2l��,�xA��Ea��pW��ޖ��a��HL���q���Z��$QR|���#��1��M4Yܞ�d�>��3Z�4lL'��<a�R����ml�x4�%=�	߶9Z�HhW��
�^K� �W[�yZ�������n����T�Il֧%o	��(%�w<��}����I��1�r@��P��*�r/�y��z
�lu����� ���>��6�!��W�k>�r�(ü�1:Դ�	,���3xᐇC�ɜ���>�{�������c�n��369�����&;���M�$������Lvz�vn��顛C�䟐ynk��r@�m� ��a����Pճ:\d���b;�ezLeP���֯4�����ڟb�4e,ple�r���%*��������`�N�%=�,7�����w A�F�i��8P���^czV�������K<"'�:��R�͔�����cۂݲ�rp~tYH�]�J�Ǉ�D�U�W��?�&
���?�%��EOx��I�\�ϴv�6Z�iգ4��A�W~����*���lٯv_�!;�TO���Hд� ~��"�cG�g�q��45��]����X��ˡ3<'�ʹ��2�4�6h�l���PA��8]��F�7��w��D&�7�����bҸ *�\��.�++�����I�Xuثֹ��n�C�0�b�����P��Fi��=d�N��f�Z+��5�L����C�Jڇ|�=����8��EM:����(�Я���c���j�!��0��î��Fx��;��{�M��!L��K��q�<A�0�"���a ��/)�%04�r�C�jH��z���92���p=h�����Tde����] ���(J�r��VM_�2��X�S��\����~drC��j;���~�ɠd���tz��rb:��U�������w���3����g�t��>��r�5C���$+�g�t^�>��Mx���-b+��|�GV�t7�����*�n�)���h�����L���JZ��bH܊�`��;7s:��O赀��X���Z;֚��ʩl����6y�:�DԐ����/�_�Dz.��l�/�S�JF�+y6�ٕ"o$<\�"Z�-:C�|d�o�dKf�ޚ���Xc|�0sb�2�\o���/�&�1���CUhr�pۦ�U7�1Mn�D�����b1Q��)mTW����a�AF`�T��G���#���r��V0�8�C
�.�;e�Y�/�h�2�2V~J�V@T2��ÅWa�������\t�L3�E�)�%�E�z���q�%�P,(�R����A�J\����Ɖ�Z2<����1�}@8T��dVY$<>[:���Z�l��������FL�IT�1+WS��<��
���	m�c�H����=hC���"�~���٪4�ʱCm	�	T�d��ܖ���.p{��/�cD �����}.��ȩ�$�<!�%y����������납]�~l���@�n�*�e#x��a��`���$�B�8E|E$�!��$%n\u�z��)x�;J��r�fH�����g�~!p�8�G�km;\�#�Z�D�r�8�������ԃ��MҰ��d��h�҂j��V�����ȵ<�F޵�R�+�#�*lo���>x�|'��PdV%����燥�|4AC�2W�J̐8�V�� $[a����ph�@�E�BJ�!�y�*�զ��N�z�U���?x5������Gfl���TRŒ�A�%.1�Xa>LA}'�a��
9,�"��d�X�W1uG3y>-�f�@Ў�}ڽd���i���x���wَX5PGZ��oN?f��1,��:��E�*9ͨVU��"䂠d�x\��9E<3��/�����ZM ��ը�y���q�3��S�A��P�'��;ƲfZ�E(a~|�mS��=���tDָ\\;-.�`�md��-e<�/�����|�cѬW�O"�Xnc2<B��[5�~:I�6�}2�J�(I�K�<J>�� ���s�o��5����L�#>Y4D\��������}t���ڒ.���I��v.��;�����
36�-F���e���+U�"y񜠔 �~�O�}jج�3K/慧5�9v��X�y@�U�|�����~���v�l�_�jh���F��$�ݷ�bi�Xڌ�1.��<x��
zi��-�P8ɢ�9�� OV�ĸ�F���	�#�NR=E�N�����W��m��f��=�X�ϵ�9�Dfs(Bȋ�Zu^�����!k��X�8(Vx�ڤP��zR!uF3"ꡰ�%��
�.��ƥT����ANWM�&�X�d=�����> [q�ύ�3��0k2�*�t�1g�m�CxBƒG�sPӎp(�¼*�����/}y�P�\rI�i��h`Z!ӍU�/e*<���<�% ��4?dw�I�lce�)��i��5�
CC�L^W�?L�j^(�S� &���@��(Q�j!`5�3�z�7v{+b8�F!�$�����9!�l��~���!�1e=V���z8����?<$,�=�0��f�B}F ��p�CS��xg��{_i)
r�8���v�N����d��D�߬�l�z��g�D!�1���c�� ���f]��듺0�K�j<�(���c;l�����px�����P�VeN�8����y�z9=&q��O�p[4O]��X��:}��$�b.<�_�;�:{��,|�đzT��D�߆q��kw�\����������k�0��=)��m�<�f���Q���<33��o�yb^m����������v�N��0��kV�T�,�R�m�j>}Ŭ���b�{�aS�	������`�[bF�ݱ�����>���ֆ�̘��v��gT��6��tH(����RN/�� e��-(I,�6S*G�CB����wߞS��q�H_�`��8g��:����
��W���2����Ap����"�?�b���L�G̤T��&��Y�tu��z)�{�lRl\�KpO��N+c$z���8����� �J�� a?AVp�q��[���0�H�@��}4�[��5�$��|����b�1殹Mɮ�ܹ��ڎS]�B4���'uJ�7�
R�KGBs��(5C���#��Ni9�N�H*��h^c0� ��ē�7�Cx�����9f�T��֢�	��F%������>֟ʹ������5�u�C,*5���s Y�����G"u�0@�p= �О9Gm6�P�6�kYǣO��L����,���.�H��7��Y��!���ݢlt�亭���m���P��x��6�
f��ӒM�>��X@�<Tvu�b���Фt!C&%�z�nF�r���Th.��u�����n�zd��b�<�z'-��}��@X��}W��B,��M>p�eBr/�%���T��e�~N�n�懟�><}���w{�*F��a�s)܈��^^�ˑc�`�U<=��:~P�R�����	�c�a��i��p9�gH�JO�_�?*�<Fi��w&��N����$���uO�'&$/�\A�_��6�Ki0���Z��r�No�*���l�_�`�;Ҕ���7�H��� �*�"w)��Ba�q�����L��X���7�X��s˼��'s����Rm4R�����n=AWM�]\�쮏��%1���eDBL�7r�֮�b_�A ���- ���ц�m6I@ �X1�ִ�Gn�.�0<�A���M��A�!�/�y�d;4�a0��5f.����.��bH�x �c���G�:�LI�F���ʗ���<v���!�8f0Y[�r�F����{�<�׊�1��mU��Ό<�a�+��5x�ߜ@
������E���i�[�~���Ju��а���o)F��]�o��c�?�c���l�n7��S�1R�"��~?�e����[��w���|b�?�t�:�r�8�0�(����\(��W��B=�"/o�m��f��5R�����^��&���:��g+�`�vVژ.��_��5�1n���B罳m�L�,qJ�v b#�i�I��e-s5��ª�ƀ��%X��Z� Wi ��P��cnV6t�Ο��S���a�_j��.}�l��2���F��y��e���$Wy�"�O�:��|��?ovPKa��Q��Xm*0�j�2hy�r{�U���̠��eᦞ~Hh-������7��(��D��ɜ��<]8MQ�L�m��÷��[�!1T� wG�),#�~�r Z�0�E�STU
n�y��Y'sh=����~��?@O���9�Ҙ0�ڻ(���tx�@�@�)GBDEI���8���2x�+�,c�O�P �Љ!J��7:��PW�����y�1ɕ�@�W���3V�����A2瑄q������LI���,	�7Q�Po��j>�m��>g}�����]��<�"v�G��aʸ��P�E`�m�q�	��/7��>z.�n����c0zW�Y�=�XW���S$"� ��Ų�ԋ�:9�$��Y@��F���	��`-�<⧸u�-���"��C�EW���\r���nWJ���^��w�;e}Z�)M�f#���)9�ʔ~�����s�&��\�ZLj�r|��h��B�����z�[h���j=B#Ғ`�2j�P�F�>��O��<���{oZ�>���|W�=��-V �]�楀-�4\�H2|]�J�f�J�;�ٍ[-@���*h�@��9B����Tu��C���t���?GQx�����ADG����T�lC��W�.,��a��}��9�HW
��"��Fd�
�W�n3tkx���j@��P��U�#��wi��Nx�
�r��vO.P�q�33�ɼ�^,��s��S*@z�9(˒ULS���2��$��<nk�/���HgZ�m5M�l��@���إr��A�ǹP3���6[f�_�(���NT��B�ƞ�b�@\�=��[���8�-�s�J��;)�W����v���S]\2�����șMʌ*h}�B�I�(䍸��S>� >�(s�+ϰ˱��J��^Hc4߭�V�]��8����l[���R��#��C�������@�
�c���Ҡ��\�4�uU������� ���~�#-K��g�KJco���Rv��k��;Ŏ�e��$�ݹǃl���j�j��� l�_�i�?`|�S����ՠ�{x�MIz��-[�W���I�]igV�@�ఙpp#��S�F�N�&*�����Gf�,���ѫ�C+D���BC�$ZP:��0���;�k�Դ��y4x�WMPإ2R�������&�F.��� ѽ�Ӝ��+@�W�h9&��Kdx�F�)R>qjo���N����72�etөg)�ICs�~��l:P��(���*\C.�ȷ�y�9��\Y���g�`�UӨ�/��]��� <泠�R��_��I)�eo]+�"|�D�
!�L��?���j�o�(�j *��$�7���
QU`����u!�v֩�8_���-�� n��6�\�(l��z�<D!�ڠ=\����ʒr
��$g�p32Y�vB�/ z!��^�Z��)�V�2)E7�8�(S�q�ANM����e�����'�S�ꮨ��7HD������4��أ��䓽�����k�<EX���5�^���K�{q5������Ve)<s�i�{��u��&�BR�
H[ORr�W�����_���F�Z��ѕ&u�l|Ѳz��ْ�%K��)�\�.���-�h�����D����[=+�٨��芌�f��T�RS(�li�3�����^H�����[�EGv���t\��&�T���R* vj_p� ������{ι��d�R��4<`-!�b���MN��-����>����[�փc��g��6���t�[�̖%1N*�ρ[���.,æ�*�*�B��a��w���S��â�7`��,8�':�����<��,�l��H����x�^pH/��=!r?l���?L!�Ȥ�y&�c_YJ� u�4ȫ�b�yG6�\�.OW�+^>�z�8����({���ď�az��p�#���@چ�\H�m���gF*�X$�I�|P���^1A^�M�I��Ԃ��	����,4�,&'��27�R9&���L�C�z֝��k9���H��� \^�5� D����ʺ�C�c�X�t��T��֝'�	@$�%^π������ʔ�y�;/�����[*�	��.���&��u��n.> ���4�I6m��͇}kt���k�����*Lk,*+�)<n�F�
�?6[���q��G[~��o�יw����TC�h�7�%�e���M��o�a���gvp��$�v�_g�CA\���n!������G����U���)�d+�db1�z(�a��j�����U�V��V�p��yr��#%�u�C!� �.N�׍��'����a�pw���F��Ǆ�"J�#��^Y�\�lʭ<X�i:�	2RŢ��)�ۇC�%c�`ϲă�p��:H' �Jʰ����ΙwU��1�& _������Yn��Onw��m�\|�㴬b�6�c?i�� ���̮�	*���lOں_$-�;��G�;�+HF*( ��g"����q��G�j�(�S�x�TXE�f��-'���y�R4R�.�=�:�dA��]|���t꠬~c��D}��7�"�owb�rJ �u"�H���!���H�I{q�X���֯��nO:�0�/��7��uSA���P0��d����\\A��A5!0w�=B��=4��g�f���i:A���"��5�Y�f�{x!	�0�ٮ_�F.�k��X{�KC�棦���LE<w()����O�3U��[�h;�� v�����8���z�����k�;��滋�J]�q��!�E^���g|��r��S�0��['~����| �G�ܐ��V���L��t���rXW���Q�6�������;C�f������7��%�5����<m����^�|��u|�<��+���=L'V�����;��W�n��}����nRaL�pJPvb��8���ŗ ?Ks0B���׀W]SX�a�Z1K�D�]��%���u6o��������ȳ_�OG.XUl��jĉ��F|��y��1��Zh$r�X"P0�:��Y|ھo��K\(ޚ�<�X�}0���2��o�7����g^��֦���h虷���7��rڷD��<�J�Xt�QC	m�3!�޵,�WM�!+T8	G*��#���r[@�0c��n=�
���|�YF>�h���~��~ �@ʋ���EM��޵�+t ��;��)�~�Ev�S?%�g�V��k,�aK%W���2J4v�a��:���P��T�x1΃@Q��-�V)���=������pg`� �L�~�'�	��F����ª��Z"I��ss��K"ѯ���U0�au��.�m��	�*�ҌY���.&���r�cK�ֿ����3���>R�$��.���w?����UP΂�"�44�܁f�Ϥ??�[W��Kθ0j!��	��8�#E2cw��Z�Z��nR?�E�ȟ��;��L��G�f�D��d������~v{��A��ᢞ\�XZǯ�rWs���L��!������f�Q��7hь0j�һ�2�m�h��!cF�
Q�kĬ������so|5�>��|�SUԆ:V���mHĥ;yD4w��2��WJ�\����G�[��=C�h�V�@���B@e��/��K����������"x�<����G\^g�28T�3Ȭw	.'��a���}���͐
/4"���dݦWg�W3o�?��@F^��E�Boͺ�,i1��x%���m��fGP���N�@DZIY,��pCl;]n9�U���
��nt��0<�^�/�<���Z���!l�gj�MyA�ePΒ�1��f�,(ץE��i��3���y�L��\qn�V��a-y���e�����Z�2��G��g��Nl�2����ш�ȴ���?2}�(Oi+(�}��Ϲ>W). ��ls ��++�l�Dܙra4zʶz���T�͔4d�ct�};��x�q���ʰ�
��bȣ�F���\���kU�L��� 8,8~�^�����"�Ke !�+08vg>#����厦k�_��t8�l�O j^����MĚAj��}��N\n����}w�x���z_�-6|�&����V�����U�T��#��|3hNjw#�M�s�fړ`�H��<BD��nB�D�Z+6��P�8�K�"k�m����x_��P��RR�'�O��&p���}I.���[m����@�F_.WCk�&u�d�	��Ff>˨q�6���2ui� &�2�StB-gČ�CnH��^API��(�*��Yݣ_jy<w���gA}���3`В����/[�k���<!b�����Z��I��e*��=�M�r�
�<Lԩ9?E�C
��j�(;�� Ers�f[�fC�QZ�<`kG��p��v1H�8��HF�{2\֢����Bl7���!K��=�PH�s7����k�$�v��S[��B3@ 5���y!z�n�7�1�)��8L�>�l
�N���l�����ߢ&����(DW�����C�#�v�����墍�+����w@��^X��Y�GZ{�6�V��2c�F5Ce�~��R5I��p�&'����;[ju���Eu��Ě����U�����'S�|���z���i&7�U��������ϰ@\Q��=��&�=�����T�%��f|����ta�'�	3��
(�^#2G�("�����v���Ϩ����yT᪛R���j�`+�;+���{�1vʿs!�R��`H�Fb����!v��CY>�R�<����q)��,gJe�6^�t����1��N%�]���䝣�w,�6\*=�lB��>�)|�wA
�S�u��/%`l�T8��*:������gc�����L��p��X�?����PEL\y��u�&���Y�.�um&*��S�D]":@\*�O�v�+Yx!zE�58��p�+��V�ş>�a�5p(���E5�rYH}3����P%��u�$��|����1�-QM?n��ڄ���F4̀'�yo-�UR� ���"�^����T����9��H9/]����^[_ �iēʲ&�9/��>_����TTb�֘X�	�t%+i��s�4#p�o�#��k�y��*�N��ͨ������)u�rMi�� R5�/�b6ȴ�����k�38Ǚ�5�����e#�,��X�$��ᡛ���2��!���쪱�"b!�0R��4�����QJQt�#&��@Dǚx)M��-�����r]Yvk���z�C\Ɲ��Mn�]�#ɞ>G����t��:��䳃dF9�b�Pz���Fd��������ڰ�e�p�Řr%)+%�Ve�<QЛ��N�`0�=�v����1�wq��Fg#���;ܾ�^T
���!��EV<s	:t�R��%�d�T��@�c�"��Wp�q�HB:JE���ՆC������#&�H���ҀV����O����̸\�\�G�6��i�@g�ЀF���D��*k�ll�{_��;�t.���H�� ώ�"m����^q0-+��u�N���kVX �����$'i\��T�4����SG�z�A��]������Hd30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�*ڜ47{^�6H�?�q����|�emHW'wNn�㣔��Ld]�m�fh?���D�����xо[����9�nL�/l�Z~��p �G��)P�A�U{q7^���h�j����%$�59�����w���׏c� ����h���u�xW�kE�V�Q�bͬ�)b� d[%�G��'kf���Z�Z�;�H��^u�Ĕ��S�l�ҧ;��(�6�Z���?��l���gtǴ�'���t���s������=8��m��GB��2��6�YOf�F�V�%�����Zo)ξ�p
�ƃ�=SX�����[��\�KOq<d�'� �@/?+�h��	-�'[��G��[8���	l	o�5rv�v���h#Lz��-��`Y�~��)�gDg5uH{���Z^9��]����5�,�'�Bo�(�s��Kw�=Y�T���h�a���/�,�^o�Բ�Iӽ��u�&ka�a�Ҷ�8�\j�&&�<Y�|2��a�&�����"�7��1��	Ū�H��+���|R�F$�H��id��VMg�5^%b`�|F@$�/���$#�c����E^k�)�luê<�.�-�0HO�p�xp��bk��p��3����u|F�EQh�\��x2���Ϸ
H�wi������?���EEdp%
���M>V�*T�\�����'��7%e��'0t��	p,aGM��;�o�$��Iq( H��ٽ�m3O��=, 7)�(xH������G���������u>�R����J�p��I�۵��o��kcS �,��%����Ɂ�j��@ Xݹ %����l7��,��&i��q�U�rQR���p�:۳�%���Fr��*�~�W��Eu�z�:M��}L�L���(��ubc�
؇zF��r����:�&a�(�"
��g�69]�&`у��s�f1�O'�Ra*�զyـ3
/b���;ȡ�<�7�����s�� JY��VHH/[)��];qT,��?��oY]L�[~��VQ�'H��ImA}����9�bآNں���ڴ�U竬�����pg@<�n��F��b��S_��Di�����>��DtKA?#���_��xw�tó��W�*E����m)w8V����1������W���wCA2��P���jV&�;��[h���*�P��`9Qo�m�r�S(�d��j$z�/�4}ar��s��՝~�B�x���c�
2�V�U!?},�NB��Od�NӸWx��e��
:��o~-����MYd�Y��"�W}�3\+e���0��#1��4�N�dF��	X��2����{��-!�ȣZ1��v�m%�E��?�7k�i��ͣ�Hh�ԋ7��ڞ�[P�S.d�o�hɻ]�����F3<&���U=j
 �~�	)-r���Sf��&S�9c��������V���@��+ru���&g`�]r3#t��3��J鿦>ā����P>əC��Z�&���p�q��^DC=6��&9�<�@�ڙjP\����k89|�4ysd�ut�Y<&��E�L8B��W�����!��*sŷ��v�ű�F�P�M�ݐ�3&~��I;פjq5�H���F�mM7�U$�
�)�'�'kCy���� ;??��삪��Fϧ4S�wU�|'@0(,H�&y�d��>�!Q�1�S�q4��َ~���v��#�����(�`�[Fc���'��R��͢��kY� ��sd����y���챭�lLl�Q!`��C-����|�a��z����`qSܕz�مB|�5#�F��Ez~T�
�@4�����ZB<(اǌ�TLM�l��:׽�ƏI�Д~��ʏ ���iΰ�*~'2�\��A��.��I����W�xi�e��u{�;�����C�֮Dr��Ӎ��U��mv�'t�P4Ma�P�C��(��<��V�T1:�nP^]�fP"�euob��,A\�=��Ë��J���H����ׁ�D�2�S]x���>������[;���t%������$�I ���&�ѻ6�SD-x��2v��u���^�!~�I�Jњ���.��V4"��Ϋ�+w��e^[1CUp*���޻��]�YExʫ	�D0BV���D-�ɵK�<��Ư����FR��{�J�!ɩ�0c3k��w.���tfJ�c-WH��V�_5���5]�j/w( $�K�]��lQ��a�o_�Θd;��O���q9�g�"�dl�)�A���9ݏ��ƣ�'�y�9� ~����󊽄��B��� ��K�&��W����� ���Yc��E��X5e��$�d��Q%O.r,< �1�E�ȋ�\�Y��z���[h���4�-&ȿ?���.kǐ(�H���z. S� c��x��+���0��-4��15����W�X�,{���b� ��b�Ky�t�f+3�E�l�.3�*�ܡ�l��L\lsE��Yi�{Ӻx|%r�.�-��H@���_F��_�)ޱ�{�du OY͊�+�J�U׾��"�PB��d�MV<�y�n�1���&U��*H�y'��q&�/r�氚���	cGI!���p>��^�<�c�]j09/ϴ�4��فI���@�	$�Rʇ�<��6��z���ݭ܍��o[�B��	��5N��d gZf��l4/����s{�@��~ǽ�𱐠����=�Fh��5`��25����F�J�?�A}䂿K:���J�+�?c�ש���Aď~����ܗ��K��JU3����\����d�U�?����|��7��/�M��(q�vq�)2�T�A� IyD6��+}����_ˏ�qP Z�ag�C�y����KvO�L"�D��v�'�j�O�/��X)��6��K/���ڒ��C�\���%2��fY�UX�S7}�$��$ID6���ԓ�{%%Y������Z�������y2��*�G�Ȼ�cG	moX�-3�w�����Q�А��]��A隬�Y週}q����*}��fTq���7�U�b���*�i��`�Ȇ~f��zK�xm�V�����sma2$����8���M���Ssٍ�����n���IyR�o��?�$X����H��a�R7��_}��^�l�g�$@�eM<��,n�=˙�kt۱����g�H�l;�U����B�A|��?t�(M������Ovg/,�^A˹]�6Pc}}�+�����߁���4��X-9���$���:(hdf�ON;b�Р���m�,�k��LX6��`(�z�Mv-M���y*O�ן
c��f�dq�C�Ǥ�$ƣ4�WόP4/��t=��l䔃,83\����������T����9�!���`�C��y�j�T���]���u@nWM�66��͗���4��'Y{BGD��C�2�y�e,�6/0���H�_g���/+�1�%V7�S@@�4�],X�0	f�]�R�ϟ"��_�Ϥ���d��:a0]��g"\R`/<�0.( �7iKy�r���:9OC�X��=���gD�9e(�c7N�<$ۉ{��RQ5硵ҫ;rD?(��*����X���I[�����L��&V����b4�����!�[&[��h�I�P�Փ3����fgn�(�C�TM�p�T�=�8�L.��'�@Y�|��<�^���NNR�G�3;��ź�݊ɐ�Cp�/��8� !�SR^���+��d��\1�j����Ҩ��������0#
7y�t�:6jŬ(�Q�[>5��C^��g/�yˆѾ=��KQ���ɟS5,oT�]&*���r��7Li'`���7JSv���C�I�AJd�8-�y�nE�`Nj��l��g& Q��z��穛�6�-8��@G*��U9�����7�?�{�I�U3�c,dkC�_�['5Q6�w���TY�ó�c����0�^�}�#6���1��n����->� �)& �U��E�2�ɱ��/�����n�S�Ȇ��&��]�%��i�!K���@O-�U���޽���O��T�
퇨;Z��v�r��"���Y�%��Z�l�g�.�fU�~o=�/��L5"�]
�LoN49���:�|����NEoچt+�c��ʡ �PI��F
�,|H�!ȧ<(Ǘ폀�ȸ�7�.LI�~��r�� �!��]�#�46$�0���ֻz���-RaQl0��5�#	m��0k�u��46���7��>�`0{��U�W���zE!��j��ߕk�9Z�������b��<�Ι����ẌS�p��~[&;��g���1:�qדW���W)��h4yޱ�Ńru��<�̉�Zv��aU^|>d.��W�����4=M�/
��$���۬���P>`2�#kۯP+oqo�(��n�9���z���a��`�}�eE���Ef�ZrZ���*$���PS�;x�Ӝ�
eP�*`.�7� s6NM?P���:�h��W-��4a>�\�L�bm��?��9Dhc�������>ڿnLԽ(�`�8�ڧ��wĦo�)GdA^go�Tj�5�z�����D�S���%:��E��[ V��nt�[yx�E�c�W� �r���� �^�%�̒��$�G5Z�M�;�jF͍;?�J
��yƞr��bS(��ZWY�E�VlY0�����3��	��V�h�.�x�_�W8ő�����Bzb���(�YU�CF\�}%K���o/#�6��	��S�dg����[��\R��ǯ�� v��?�8Wh�r	3,�[�)<�[���3n�l	58QRv!դhi�j��Z��&ԲYl-��2��m��5;����-��ѧ#x�gy��r'�(���h�s/[Y��=_//`�@e;Kac�x�5o�$|쪤]�S�;����MN�i�,v֟�ׇ���_�.�k��٧:�ý��X,�v�.�[�\�������J�*ezqgg��n��HJ�����7��mE��P�И�x���b�4��B�o*�1:~Ɉ�Xp�bo�so��nx�w��1�%�m*��W��J<��Q�����X�n�K(Ow٨_|!M��h�XQ�;? ��:_)��G�[���G�1�?PNlQq�!���K#�T���­+D<,�!���ҜÌ�/�����88��+�ƭ+�����/�}K�<Ђ�FV�$88��]Bh����)�H��ls����ʩ
6�>���"�ߵ�>`T����.*a�i�LC8U��^���&� $�!�1� �pf�O�o�#zI�쑪ȑ�Y�~��g]���F��F���+��H������u�
�ғ�q���F�T�+�A�X��w�'�	J?A �0�Acyw(��])����m(*���ˠG�p�>�2s���?���l�\��U�m��2TDv?6�>dpG'���d��dzR_$�Oˤ��	�T�but�G�L��i�6g�&��!=w�û�TY���s���
��d7g�8J$1�!l+�f��|���r���� ��{��S��=%0�K���)1��|���m�R���� (M�]�Q�խZK��-�-�C��l��e�&b`��CO���P��n%�������W�_0��b@� �O�/t�����{��k�ݰG��ڴ��)Ѩ%@W�P�z�9J�w��!�a��!Ns�-COQ�]QwIw����_��&S[�%~ڬ��c���d�`8p��=�u(Y��G�<p�����c�@��c���<�t9'�=�4�~�%�p�Ze��	��a�����ZP�d=.��M;u3k}vGZl�T�ʋ[/*�i�g{��$��E]ΣI�ci������'ӄ��'$8�E�?���/��ƥ~��4�����&�6��j�B)��ˌ�w��x~;J�c��w���;�/���y�"���PP��h(�@ܑ?˥X	���<�������j��8�8�2�^!`�U�{�2j�]�w�B�v�nUk� n+2G �0vD�b/�튑����yH���W��Jѧ�Pp�YE�����O�%1D�&�$�O=7��G��Y,����g+j�+�N37�4�t�殁�ˎ���̹�9i@�f�ђA3'd��F���.�DZӮ�d_N�]T@�e�~t��v�1y*��ڟJ{��9q��]���sǜ�U���L��h��Z�rr�����D�K@zd���V��%�!��9���x��V�Ҕ����ք���|E�':�e~S�N��x�2w���Ԙ�ū�٧�rw���:��f�N��L3���`!���m�^��I����� | �N$����0u#��t���$�ͼc2:�E�_[����0��uf
|:8��G�arFji4OК��"�g���Z���\�G�}�Ok�T���>ZP�xv�)�k��B�\�`��Zq�����f�M)��.no���Lz>�[Ib�L��刉�����|��-�~&�2�ʼ�:��}��U�'�;�
�غ>�r�D5Y<����}Zj�Z�K���=A��:a�2�N���O�8٬�j���I�	|�5����U�n��d�8���B	2`hH�:�=�RҠ�52'i��Vz��5+����%S`�����qz�c��z��kZlB������
10,�Oşx]�n�Hk���[��5�G|S��E�C��� Vx�E�e��
u�.i|��DZ����E�o
=(]:V���H�T=��A�Ҕ�#72y���Ŏ��T�,^MK3)�{$���q�cY�����&G�\F4,��ѵ��$��������.f��fW>�<�Ǻ�J'���K�Ԩ���܅kp��ْʷr�7���t��|*X�Zr%Qփ��tt��6���e���@�GLr~j�Ѳ�~:H�&2Q ���5rg���5~G�i�rj{��:�A?���L:����aN�b�����w���R�hj�e ahI"W�t�T�:9꼉&����f���_pO4��a�G��"3��)�C�;�-�<IA��Ӏ]L �3�=��H�釕<;����h�J���jL��8�2)V��WH��mκm��:�9YnȢ�_���@|������ �����1�p4ɭ��f�S�״��Sl�=�1z�T\��>�zkA�⠀�3�%�j�����Wt������m�m��3V�^��̛��|��y&��»�驣J����nV�xw;�^h��w����H�Q�����p�(�� ��:�<j�}أ��6'��9�*�bB��|�o]�
�1r�b��}مB��O��N`nW�J�2��
��Co���U#�^b�dq�O���RW�&�\�X��_���>�1S<l�#�d3�	�1&�_�����y�����{K1�m�v�|��>�����|W�������Ё�$�!�2��e���,5�54�]C�ޅ���&S��d=����: o	���r�S#��*��ie���ض�f��T@�Ner�:�33��
�#���� t��U ��o6�N����[PK�L��K�Z�&���z�q'1�^q|�=ߑ&�壇M�(�Xs���k%�s�8�es��t�5\&
aR��8���W<��0�!5��s���Cf�U�]��MI��U叀 ��3H�u�q��$ڵM��Sa�M�"q�Z�px9c�'��^�`Eڍ�?L6��/&����4@�'U)~/'m�J,e�y.��K����� ��4�<0�40������p�!���5��QF�ʇ�GGR�����;�8#��ms"�)��6!����٣P��{m�CrH`�O-j6���t���������H�z=���R�B���#�1�����z�60��6�������+�ѫB��Q��4zT����Ղۜ�"���j�v��K��B� �Yi{��*�~�I�iA�ڠ.�P��AB��`W�@}ir�P��Tb;ts�aVKC�H�D?��@?�b�!7'��P!��-�.C+8Ȱ�5�%%�T>�SD��^�qWPqu�<����A)4Ѫ��͋.��e�xhﭱ=�ѻi�J\wx�Bk�4���ؼ�θ[�|H�3.%�
��������I��X�����hSZ�e�1A|�T���Eu[u^�?^hd�VN��G��E�ȣC�"b��¬��$^���Ch�pא�+���ثvY҃T�6u0y�P�ֿ̼څ����Z-��1݈ĂJ |��o�F����߅<
J�!FW5��VF�V_Ll �R0!w5��$@QcêMCl>)����_��1d�f�p" ��Dz9���o~�l��=������\"��3��'�w�9��~7O��\n�J���~��H�7��3�����9s  ����������he쪙$��D����.�ے ��E�K����&<*z#�G[u(M�9��z�˿,H�*"ǽ�EHY��z�d�U�%U+=�n����d�2sH̎6O�.�X�����w�b�� �OEyM��fXR�E�q�.o��7\�BZa���s2����{ �|��.[�e�q@��O_P����	�)k�6{�=5 X����F�W��U�f��񓪈=�(��2��9yL��'���ftU��,�*�'��&�q/�`��g�9�vu�GV���z��?�,<m�]���/�$�4�!i��xS��]8	�?�Ԗj<����qV��	K��������O�4	h��Nl�_�Q�Z����^�与q����{�ע�����
������XU���]
B�%`��JS�
��;����}�q�Bg	�O�\mN{ƎW �=���
��o&�kPګ����d,6��XaW%�\Ӥ���e�U�i1N�}���=d��%	����ړZ՟�"��}Up�1���v6i[a����V�ZW���Q�ڣ�b&�|ڸ�|�IV�_���f��m�� ]~����E���&�D��Q'=�	��	��r-�7S�v2�Ŭ���=�rپ�/��a��@|�r�����/�9�#.��.�7p��N�R�)����P��C�돓ZA�̅��qB7�^�E=�ׯ&����蒨�g��h��k����S�/s�t}�f&E�m��8�ɘW��'��t�!Pi0sm
i����Y���>MDD���)��֤�N8 q��y������=%M�r��+��˪Tz'撨Z���'$?�}��*a���Z�4���UD_'��m,�%yQy���wg��,��V�4����6���mi*��k�\q��˙��F����BlR0qj�u����n��bss�ؠ�Ҡ�! 1�*'��۾��`�hF-����˃�	h��"�H����%z����-��B$O#��3���z&��Q�G����4u��x�B�§o��T�� �0���+/������&$��T�? W��ivw*&�o���A��!._�$�>.�G:�W)�[im\�Gg;/Q�|KVCO��Dh��{�2�����?'�Pܵ�H�~C��ȋ;��`ӋT�|?��^�sP�qu��a1DA2@�ǘ����Y�����h�l��qt����xg���oϤh7�ō�[�h��A%��}�j�^��*IȂ0�7���c�b�����5ϩoP����>u9�^�>���o)�B���ף�d�"9�}��&��V�^���C���pҰ��������YY�嘫��0������\�q�h���U�W��i�7ݣ)J{l�Jд��$�Xͅ7ӣJ+�W�Va�_ǧ*����k'�w�q$;�����l��h�	ы_Ti1d��V��3���}�9�T���IPlC�������v�7#��n�'*�9���~�EC>r�e�+R-yw4��r:�������Ż�`Z� �����MSX1���Te'ݲ$zV���K�.(� y��E�N��I�>�z^$![N�4&;��I���g�E���8�H4O�z֬�ߨ�� `�+�8���q���	ǭ�~�i�N���XH�,����bE�N�
�Lyhr�f��E�t~.�/#�ҁ��=3�����s����j{{��|͡�.�R�_p@�t6_��z�R��)��G{dgs ����2�����U�іL����ܭ_i�f[y'>�Q���p��U����'OH�&�&�/ ��B�Q���G�RE�u׵����<(�]��/w/%4`{Á���x��	�z�/f�<B�|�h	΄������U\���Ca	c8�NǡT��Z���y�>)�5{_�ި�\��e�C�Y���zA����eh�A5��I���t*��ss��h�Ⲃgf���J�%�+A9���n�zEB�&Q�^T�k�0tJ��%���\;�_��Ф�[�ž5q��dÜ�W(��v�(*�qy�92�_t���+I!"�6����n�p�#_s�q����	��C�j���K
Lʪ��,{���= (�/��X�����&wK�y���o��p\3X{%ڄ�f}UXG�0}5z;�@�pIģ��BN���%�w(�t�/�m����^�,�� �����ҡn�p	c�$��Y-�h��Y���ïQ�]n�)�ٖ���T ��0�%?=�7J�}�e�f�=��kZ]��4�[�����*w7��V�p��f���K��nxY�*P���{�a�O��8�8R������$����΃������čR���:�̜[�1�׍�p�R�ޛ_%��^7�g^G�����j��,��A��t�[\�g/�gs�!l�^L��a���k�A$��HMt��!�_T9y��t���20/��>As@H�ޫHN$���#��v�qO΃i� ���r���40K(]���[{
R�P�Tm� �,4S��ي6vu�(V��Mc��C�F!j��ԽcR����bĺ�I�L2�Kr����P�~�ю�r^a�+SS3�3��S{�c)�����ԙɰ!0#�`�]
�!7,j9x���U�~#n��wM^��6cUS��^ƩX���psk{�������3Ȅ�6����\H@��g�����e1���K�8�>L��<��ܰW]��#�ؤ���*���y"m�~�w��ꢉ���u]U�C"�/���.�m�7N|�mꊇO������ћ6�~DEq-e���7�G�<��O�#B
��Z����SO�D����*R֋�]�l�>E}��I.��"VsR{�9ǫb܂�����鞚-T��=Ұ}"�ϙFZ�@y�О����p�L=�����%��Ա����$����y��=n�R6\[3�?��b�⊾|1��:'��l���+� ���R��ӈ�d��	�Ҹ�4T�ͬ7ܟ_���V�[�^�0�uyl��:�mh����Q��>��V랪���g�Pqys�ƾ��K�+�ʈ�Sݖ�Tj���3��
+�&7��l`���e3S9������d}��-e �n�/`�>L�Cr��� Qtײ�9��S�i-�Q�����bn��(��ш�����;�,��#�k�X����5���9��]&�YZr��*�`��slf&�˃릞#"��k�nE@��J��&�֬�(�2�o>����@8<nq��S���H}D���I��x_ii�V��S`@�&cN"��u@ȕju�֟}ȳ�X�/�nZ�����"��[4lߕ�i�Z� �gJ7�f��o�u�ut5"Mz�� �4�e��m�C|cꘝ���o���t�E��� ���Iw�5
C�|���!p���=�7�p�p%f7n03IN�Ď�S�e��1�3#��$�РքX�"Ʃ�հ���40UŞ���#�ߤ��29uI�%4�R��sj>�L�0#\U�=��r�!1�`���Ik����*�]�ϡ5j�A�&׶��Xt�r�&��,F/�&2�;`K��9��}�;Bgܹ�G)Q�
h�Bݱ��[r����𞉄juvq��U�z>���vIg�c�{��8��z�.�d�)Ќ=8�>�m#�Pӽ�o�L/�L�9�M؋"}w~�ݴs+���eŻݦT���3{�X��*�!މ�/��L��DF�e��z*��7i	�6�
5?������F�S�OW�&D�'�����LR�m~=�?ed]DN�t6�l��B-��g2�L|��#wނ�!�D�̦�<����2,^��V��j�4�"�W�c^��rK�s/��@D�׽�� ��f�K���|���n���g����b��W��yU!rf`r|EӒ�.wi�?ߓ�J>;�d�s:����{_�|��.c���|{@�<�_X�N����)s�4{�m� $�����ڌ_(�U�Z����E�&������yT�@�1�݁YU�4��'T'�A�&�I�/��|�o�~�fG^$:��D�G{U<u
�]��D/�4��܁�b@���	����ܣ+<����y�6��խ����".��WO�	p�rNt<��Y�Z���67��g&���{�򨷒������g��r\�h�Gx5{hG�GL���������4Sv�9��"����J�n+��佌���'��sr�K%(�����iJʅӯ�<\HE����Ԥ4@Cū���=�S�����¹B(��q���27˾�6��I-163� p1�=�5_��q�3����C�H�w:�K���L�T�����<�5/=�X����k�Kd\n��E2�f*A\�K�%��;f���X�l}"\����I񴚲UyǓ� �%ڕ��!�������:��:a���A�?��}�:c�ad�n-ȄN��Jʎ�Qf���/5٣H����Nqe���� Q}��f��"�����
t�iRS��Ń*dWr�$j���	fm�UK!x"kw�ף��Ea�B����8#�¹.�h�{�����0N*�c����T�Rz�g�2��b��QÍ��XR��p_r�T^$_g��:����!�]O,#?����tT�T��g �
lXV�y���dMA1�<�tՎG��1ƽ0��J����]/A A�L����X%���;��$x�P2��m٦�-H���(]������}�`m��6,�\���6#Tp(�O�M�h���BN��L�c�-���\=�fR�Ǚ���8M�ό`P	�k�La����8
x3�%����P��ωBr���!�/�`3�.�ij�m��̡��k8�n7l:M���60ߌ�"1�e܀�Ɣ{7�����߃g#��:�6�=.��HM�xg\��$�N1�:.��!��9���?�I��]��9���u�RYW���:"�]��ov�o��O5t]bV&�/%m�·_sD����#�tD�^0颒4�[��<���[���~��VCV��	Eqb���s6���a��jD��ݾ�M�`�i��ލ���������pm�=w����]ş>�{o���������J8�z�R�|3�!�2�|�����(7����bͪ ��R� ӷ��/dv���y�r�|���/~�&99�V�&0��ly<}�:��׬�.�Qg]Q>�0C�Z��g} �yC����̈Kɉh�X��S���T:�����a�\���7�p�`���5�kS�ػ�򥒳dM��-5j�n��`�<�*�ߒ�QD�˺	R�#�l-�k6�>��2<J���T�Ј����q�����Vk�|�d:5��	�
-�]Y*ژ۷���ࢨg�Ӽ���O�nE����n��ϥ��xn�&������2ug��V|x�d�nA]�Srb̀����oȝ�7i9�0�s@z"��X�Ep�:���o�ȃ�	��5;ZYh��{�"}�lӕ�clZS4�g��f�\o���E>"�+���4�/�=��|3hk����oR�%t�z��m�) �w�IG��
��|���!@Z��c�4W�@�7>��I���_���Ś��#pQ;$Wܭ�Tޔ��)����0%��ѭt:#�����=u
�4�!���}>���0��U\�g�B�$!D+�`�ikT����t��]qt�q���W׆�XDԊ�����ޜ�ۃ;0/u�r;��!�Tm܉2)!��h���t>�r�i���TR[vAËU��y>� ��F���39[������x��a]���ߌ$�>�1#�MP�׵os��Ր9�ճ���YG:�݄�����
e��6�$���е�(Hh*�s7�����R��e�?�*ؕ�79w�6�2F?ȱ���GA�#��W��D������ML"T�mN5N?5V@D�yC�D�x�<9
�'�7� LLe�����Rl���$��S��-'�\8^�P<�&��jj̔���3ۜ�˸c�C/Ӹ>�׍�\ ��͡�y���-�xUE�E`�϶���'�s "�%e�ǒe��}��Zw�k;Ed��d���A�p�����y�(�2�Z��	���Al�PBe?�AR �Z�2��Y����`��+E8={`�	FB��S?,Y͆�FԆ%�5�co���)]Ɓ��Ss�F��[\\ʡ/R��� ?Phh[yH	�`[%����������l�ڭ5�Q?v��1h�(���P�Y�8{ª{���M�5�����6����q��|���F'F��fY�s�Z���v=��Y����6a�8H��(��d@�UU�o+�1Ƒ�Ų����vN����w�@�.����u�r:��?�54	��8v�f[T0�;����KТ;�q�����H�yqg�fԯ������{/0��a�-��bH����~�*N|U�b��8�b範o/��n�qw,�h��ƍ*vr�>��<lk�Y�I��~U�õwQ��|����N�H���Q�9�Ǵ��5y)I�'�g�oi�ީ��?���Q�?x��x#ER�O@+p�,Gݼ�E�������B}�	8Zsك;�+#�� �}�m�<H����tF�q8�"k]����a��)��a��svC�^)��!��׶S���,�-��`̯�q s���Ϥ�&�C|���?�� �X�:��䙱�12�p�E��'Cz����	1�J�j~���]nr�Fu�8� ^�.�K�L����,
|8A�8n>�-�F�N�+%�X&lwW�d����A�-�WB鉶�-P�P*�m�����K8��4mŶ)2�W��8���u[�f��m[�O2̻F?�[�>ܥ�G��p�j؉��\�_U��+E�y`T�Eu�AG���L &1��؞�!��h�;#�T����s�9߬�ܚ���h�t!�{!fkUI�3):r$��a�o���q�ؓ�>���;"ߡ��æ�����]��-tM9 �����%�K�\�?l�-#Q��������bخ�C�����6���l��0��0���>0y�b�fP�ǚUt�2(�n��(E��]aԴ�XIS<@ϐ<��ФJ&LG�H\a#��N�X-���\ �w�h��	���=V�[SDp�$��c�-�dJJ��
����U(њ�G\ɼp ,ܷcL����۱��}�t��=E�~eE�p.i����N��at��;岫��=��@qeK�9~�K������ga�޹/�����s{��[$.�E՛q���}��i|s��o����岀��$���ɷv��tȕ	�L~w1��I�J���6�����B�U��0�̀��~���c&�s�NӮ���ؗh�yuج�=^sP������	�ĥ�89�w�h؍˨�K��j'
��z#�2��7ť�jkE�w4�v)���e �&2�b��xD3A�ej݌]�`���@M�S�����	�Y�_�K�.�Ǵ01��?�(�����PnGB�@Y�́�2��+��ۜ3~s4'@��&������;��!i@K_�IQ3�����	���`�D�TtV�N��@]3�e���p�1����Rʐ{�q��,�լ���mc���F���hDu����@�n���K�)P���+~ä�Y�h�Rv93�x 'V�J-�3�N1�0�L��N�e��N��ï��K�e�Ue7�Q6��Ԧ�g�W�=SN
��3W?�`�P]+8}��c�I�;O�p$b ����&G�
ԡu�{���K
��@�4�_:*��ח��6zuނ�:�;uG��F⮳Of���;���gI�qR�z�\��}z�[O��TP�5��D����)H�X�/�{\Fw����c͔J�i�c���)�F�n烯�0'fz���>��s�]c��,B�f�M�V~�Q�B���y��4�U�2��P�O��L�O5�Y:�S�K.�8j)%*K9'w�{�����p���H�f�ݷwl8Q �j����K|WOs�Sċ
������L��vE�	��HQD����RJ�ĭhii��V�nV5�!�E|��aL�T��~c���k��l�4�!C�H\0���O��nxմ$g��kc�d���z|ˤ!Evd,�!P�xk��ݕ�
�w�i�IfҼ��9��E��k
�O��l,[�/�� ��d&�|7�Z��L�w�Ot�,{$�M�zF��$�q��!����.���]C,����-�$�C���!�ц�����v�g�{�
28�	���}~���i*uS��E����FDFd���-���n�Q�`8̅GKE�ڴQxƺ�V\�W��-dm��v���z��,�Xx�뵋�u�-0��̏�k�"�M5����a�UY�
ט;.�=�ˢ܇L���Ϩ �"������n�C�����,�@&̮R���n2�X��
�ۼDrVn�1PS��N�̨�9�Q�Bim���3�|@�$	����y����u֣�:�7K��3ZL�rE"1��8��Q�Z�$g��wf*�oi���y�~"�����7�4e]��q�(|�����}o�Zt�X��!�7 ���I�0�
G�;|A��!t�nTG�;n���7rϫI�4Q�,pL�;�5t,#$!�$����k��&)C�Ytn�Ӳ0�y���[#5�����u�
�4�8��c{m>�D%0�T�U�F��>k!5�H�_=k������Pf�%r��E�S�:�Xx���
�0�B���g;d���&^e�׿�tܽ�)�Kh�!�(�.r!�	�h�t���v��AU
��>���z�`�����@�[��2�i��Ox�A��>�a
#�NPW�o�̘�S%9�*؋��{� �8b���}�eI[��X!8���g�\�X*P�0��!��g��Hɵe|i�*��7�ݤ6�o�?|�Z�桵��U�W�m8`O��L�.dm�f�?�jDȸ����p�Ƙ^�k:L S����8��HO������m�o^�d��U�j���/�g0��]�w���7k��H 8������x�o�E�d>k͞$�[� �7�%��C��{�fZ+�;y�4͹E���Y}�$��x<�-��(�D�Z�Tҿ�Al����Kn���Վ�ҧ�iZ�������d8q�y��ҋB&��FYdlF�
�%�/U�o�T�bg�Ƶ�@S���z{0[\�����G@� �o�?L8�hh�	��{[� ���_Xl��5dw�v��!h�Q��E�'�R0�Y��^>��	5ge�P� ̵��C�OஐG��''z�g\s�_� =�E��"�sa�����CF�P��P�.��e[ծy�F���v���3�*��5�.�KL�)�:�$����I���v���[�	Ɉ�`��FS2�V�Rq��ÚC�H�U����ꝙ�ޯ���İ��a&b�����*�*N�����b8�o�aZn�rw����H�**ڻ�r|/< 1�ۍ)�������web|�b���Y´Q>sX�7o�f��):��ۃh�����]n�?���Q��s�J��#���c+3ة,{;���!��8������8�zٷp�+����T5�}F<<|�2?9]F�8d��]����m)5:����s���3��U��jc��+����p�` ꬒ%�u��""���,C�7���T����w���l1���p�$���z��@�_��~��~�j"]���F)On�4�@��.~�<h<�8��
�1���Ԕa�nF�+o+Y�LX��w����5�4A�ؓm�#����9����mT�+��O��s���
�2��~��6���:cۚ��m�[2 ��?bZ�>{HGS.Ȟ������_��f{a�Be�T�3�u �GH�LT��9�^��8�!iy	�oAT���2V"��B3�u�d=�F�!���f�)&�烱rL�W��(���E�в%��i��w�'��P�͑W�P(R�~�a6M�(����٠����-Wꊚ�[����b�+�C���|�2�����j�d�=�4G�0���blW����7t��E֨�"ř�\�گ	_�J�8��@�|��2�JZ�r����aWPN��-���=w�W���W�q�I[WL�XMc���d~�ddW*��m(���G�IZpԡyE9�c ٨�V��h>t��*=�]~��p�c�3=�
[a�2��L�˴�=Z����*��J)��ܝ�+�aʷ��/���ܕ7M{��i$��E	ՇK���ci0����j0�S����$d������G�=~+�K�}d��Rk�6�2
Ö�B�vb˸w�̴�~~g��cZC��!��I��K��y��.��8P.�3T�p�=���4����:�A~����j�9�ɮI�2å_�\���j�e
w�?v];Gcs )�2s��܎)Dː!�~Ɍxϭ%���2̈́��k����t"Yq1G�5�{�1��)R�!���涘fGvBYX��f��+�-�����32s4[6��x��:����>�U��@3B��}�3S���󈅯�mD��
CN.@�;e<���$�e1%Č�o�{��qe���	�"ߟL9����x{�hxG}���Q�t��p�=K��i���~�lb�z���C9�Xlx4Jm���삹���5�d�S� e*��N��t�����b����q�f؛P��q�-N�53�J�`M�}_૨��I��ț$P ����z+�>�uOa3� 觨Pc��h*�:ޝ@�.�����)�u��:��5G�n�F�O���F�3:��g}���?0���\��D}�5�O�b�T���j���$��)�3�c2�\���I��ā/�Ȏ������)���n����z�*u�������K������ٶ�R���v�f��)��U����������&� n�5�[��b'kj�9�Km�u�/�[�.�Ư^Fh����+��8�B�jE
����|�G�J��?͗�ҙ������{�	^�H��7�i�R~/�a�=i���V�"�5�K����謑�u��c4ȟ�&�k>.�l�R��'�|�0X��O�9x��1��tkL4�,��a�A|��E*�
�U\jx^�
��{i(Pb�p{��mF�E=�N
�Ofs���l�l٠3_���&7ޱ�� ���hk,/��M����$A�]q���UϬ�F��F�,9~�a����8�U���D���>��͌�>�����KJ�n$�wo��T�����k�͘%G����0��/��8D�XV(=%}Y��])��4+�)���
��]r����^Hb:tz��%���X	r�,ݕ�~�%���
R�:��|�6�Lf����i����C���$�G�ٔ�5�ea���"[���2�9��l&���D�#���vO�OQaæ�r�w3#�-��-Z;!v<+�@��,�� #N/��HH�A�3��;���$?���L�B�Ÿ�VJ.�H�n�mz���#�H9�ݢ��i�����zڭ����Mk���J��Y|p���J:��{�;�S��]� �������FA�1߀FA;�Q�y�m���7\^�:@"��m0m���V+
�x�Uɨ�8�tI��3>|�z�:���qڿV���;���h��ׇ#�C��%�Q�<:��H�(C�N����b�}:�^�l
D�����B1+�'
�0���} QB�]iO;[Ns8W���ޱ�
�d�o7\K�	}�
�d���,sW�B�\��ߩ�u��f��1���G��d_�<	Od�����pzs����$�1�+�v� ��73�x���(�ξBmԣ�rZЭ�n��V��V㹌�V=�S�ᙾ]o�W�^��]O&�]C���=��%�f�	�M�r(�Sψ�����2�V������ȿ��@M��r�G�ߋ1�6.)#m���L4��#���������6P��k�&�Z�F����q��	^��=��4&Ұ���'�C�޹�$kQa���_es���tN7�&6���]8��W�̀.[!��s����S��J���	�FMu������L`��Ơ0�q�����\���UQM����6���%'İ��+&tڹb$?���[��?|K4l*�U�Ծ'���,�ZyBc���;*���L94�ٝ��vQ�vF�]��M ���f+9��F\^3�@PeR�,��&� ��&���'s�0��p�rd��ˉ��6�o�4`n��-�a���hc�:���s���,�O�zigo��(�Bo�#������Dzw�܇4�y�:��kz�BՅ�����T�sF�Ɗ�����Q����Z\����E�� h�i��_*w3\�uA,��.q�|g��8}�W:�#i���np�;��Ϻ:C �QD�є�l�Z���F��'m�TPM���ِC1#-�\�ɕQ��T��p�j^Ve�P;�Bu�ˋ�g�A�����G��2P����AX��ن��}6��v,�x8��`��y����Ԕ[4H��t$%>q��U��p�I����H֎є�?��@] ]�q�u
��^��ɿ�sn�񙿣o�x"ʠ�IฬaF�^���C��p����1�Y~�|�b�=0����|�Z��`0��ƨ�m��"T�4��J,h��Bu̫��0�q�h?�J|�mWa��V��_xĠ�f��\4#w��$lߋ�V�}lj����_�d�亱����9����;l���El��BJ�X�_D';��9�F�~�z���׊��M��H�r�cj��Y�0�A��P� ,�����h����v]en�$���*�,.k�� �CE1��
�5�zO�[!=��eXU�&���X-׾֬2��m^H�4z���߹U	�Q3�+�q��I�Z�f۽�^���:5�5�XYȘ����b����{جy�D@f�
Ew/f.�D��4S�nH��E��s^B#�b{,�|���.�Ȧp6x@�*E_�X`�ÞA)�}{�c ����#�Y�F	U�,���i���4���[y��O�B�Á=U��A�'��&+�P/��F�?(⢘[G
���pn��Y�<���]��S/(��41{������	�I�ʀ�><�-G�A%�5���U�z�F������	�4N��}lQZ�����
e�d��D{p$S���}ǶȮ��^�'�6hv�5������D��%��?7 �X�Rz�����J���+Ruܽ������a��)a��0��uX�uoJ��ٵ\l77�]���XK��O�a����ݿ�涁(*h.q���2�e�Z��I� P6W=��S�aw�_���q)H�Z��C�r�K���L����}<��}�Y`/�?�XBb:�o�K�l�ДZ����\D�%h�fRƑX��}�[����`I�-��y���2�%��l�����f�#���R��˜���a�d�ġ'cc@�=��-lL�
Qn�uQ����:)(��v���zr����#k����}b��f�$�|�.���u���*焳H���A�f��K��fxFa	�{^��)T�aD6���u�8#���쾍��r��l���~�催nR;c
�����6�B�����R0o
_�{^��cgB�����s�{K�,G��˒�Rt'ׄ��(g$�Vl��$��-����$AU���Z�t�-�+J����G]��_�/�pA�m��/|��d�v2�&X��t�����{���Ğ(�{MɈH��٠!Em�[,E�2�%Id6���(ǚ�M�P&������p$�cc!��rn�
-5ǽ����`5ϰ��P�U��p�j�-��\�3Ud5�6����ϭ�Q�j�!!5B`����R��j��𘱁�n[�EM/s6TȬ��/N���?���+{[�k�0�R��W��ޥ�6�ص�NiHqOYg ��Hx�1=�(��p�l��q����]�'��)��v�ȵK��"āH��1��n]]��6"U�/U#�.ab�7��`��Ƀ�{~(O��0��0��!D�x�ea�97��<�A������P��<Ҥm�DX���c!I�<t3�=��/���!�߸V�1㪐�bmz��T������G�����|W�����/�a�5��pn��=�����-� д�,W��ChXi���Q��R'8T3���œO���ė\��Ugi�Cxl ��R����cd�W*�����:�=3����'���w��0�_uy���:/�/�Q(�>�}��{��g�-Qy�\��6N�Kj;v�}�S�F�T;u*����h/\��7E�`'r�S�	ؼ�}����d��i-��pn>q�`%o��qI���=QE�m�*�d0�-��9�n�� ��a5-Y��0��⾘=���<&�k<��0�5���굂.��YK�јZ����H�)�iw�ȹ\�ܦOx3��Vn6R����+��)�&��+�26s��7 �dZnb]�S�f�yc���K�>��i��t�`�>@{�?)m̆%����b�����$T����Z:B'��]�"�AE�����Z�.�g�/�f���o��e�Fc ">CX�Y4/@Ӿ�|���F��o3{t�>���9d �?aI�__
��S|.[�!����iY�a�\7�I���k-�9ƚ���#Q�Q$X���uD�30��]J��0�A,�n׼#b<���%�u:4��C���>@�0��MUI��#�l!�t��r�k�{�[�
��T�t���ʠ�gK�XE��	5�=3�W��;������s�����܊�C)BT}h����)rn�p�U�y�v"��U���>�[E��8����K�-0��H\�������p�>���#$eqP0do�`���69S^�ӟOH�;ݥ��ǯe��㦥
f�s�R���*}e,���.��@��U�2e):�*Y�T7ڍ�6��?�������D4�W��}��tL�{�mQ!?�vD�L�e��}M�s#Wڸ�CL�<��7��3Q��L���� � �j^`j����j+J��ӵ��4͟���ċ��Z�q|u�ߚ %�̡�(r��xV�1E��,�=�K����� ��%&nQ�FYE�~VfZ�L;�<��fDL�C.͟9���ҧZ/�(�wiZ��ÿ�[8l2
����ߙ�9ާ��Ь������8~�h���UBsX���%Y���F�Q�%�\?�o��,�}��|�S�"�N�[=5m\�9P���T�� O��?� h�9�	l�t[;��ؖ��8l�'�5G�v�=h����-J�VY岍��5�&Li5H������:@�|����g���'��`���9s(��r�=�T��^�ޒ�a��������S����lt���^��c���vooa�@���ty�.��:Te��6{��U�v#�`[��i��i��	��Cb�q����rH�(��g���,,�F���v�б͈����b)%�����*o��7�ݝ1�bh��o��nDjKwَ��Wr*���r�<������ �q���CUw2+)|��F�o���g�Q�@8�Y�S��)��'u�p܏�ʐa?	�QJ_H���L#�~��0+`X�,H���fa��E��Yz���m8����D\�+�[��!8�}�b�<��)�d1FO_f8Q�]]{'�B=�)�6�� �s��p���ʢ�]�W��ָ
��|`����7��熽�B�4C��;�ଆ�d��$�Y�1S��p�5�H\�zBB���J~�;c]o�@F�(�Ao4���������%�e
=N��<6�.F�+f��X��iw�Q�"��AYt\��v���N�X����mB7��'�`8O�w�.2��ȑ��]�b�ۧ��m�k�2M@�?Op\>�N`G�H@�k�Q��ٳ_�v'(uܫ���T���u�zGu�L!t�����p!�_⼉eTr8B�����B|��Yz�ѻ��!Eg�f����pzr�_>�B������=NE��r��$���"ѐ�������bv�.;MZ�c
�UՆ(�D�����-��F��������b� uC}�)���g����<���G�a�0zc8b�Ip��qt}It�Ms�&���D �>YT���jǙ@�H�S�/J�X2���a�ֽN��>-��}cp���D�8�]l��S����T���u�GI^�Lu�Ιz9e�3=�!�	����TF�	��5��+��1~+��jq>�!�f@�q�isr-sV�����>c����J���?��vG����1��tˀ�a2M.�D^�Q�ZZ����+-8*������2_b�k�C\B��#��|��_¦E%��5��0���b�H��\�-tQM��ˊ��n��=��'Q�kfn>Z@dv��'i�J�꼼}��a8N6N�;�-�Q,JwV��>����|[�b��9��c��d�Ь�[r�J-�(�AG1r�p�޻&@cJm�0����tF=f=P~:�p��w�cj�|a�@��0�n�,�F=ۿNFbG�
G�/��L}�����/�s�#�{XZK$�ˌE�.L�-�7�iqX)�;�����UY�$%��̼���|��^�~l;���]��8)6U�H�W�$B��6˹���1~���c��������[؀�
ry�����0\PO���\�ܞ�7��]�Lq��T�`��j��j���822)m�W�(4}j@w�ev>n{H\� ;B�2� G�=tDL"��:@Ό�ml����~���J��c+TY� ���<�1ю!S��N���7�Gד�Yم.���+W����X33�.4|��˛Il�p����@��8�^�Z3T�ָ�P���xDg� ���N��@�Wwe�Z�%�v1F�ÚG!{���Ҫ�u�`7����K�y�h��̚���Չ�����K���q�O� W��b��(�9(m�x��Z�ߍ�Z,R��.ÙEd!�TeKRN��l�?]�N|�*cl������B<����N���3�"`��9 ;�K��I�GǛ%�� �tJ�6_���u�\��S�CX�IY:�q?�,������=
0u�\:�H�G�}F�D�O
��g�+{n�gޚRl�O�e\��}���O��T����������)}����\�h�*� �Ũ��Ͷ^yV.)4�n��I���Cz�F1vF0rA�R,����ț���zw���W�lg�)�J�SU��H�#݅Jq$���s-5�HԢ�#��
j8=KΘ�ݰ)��ϼ�}�{�+�,ˀ8���j���VG|�X��>�� 5���1l�����W�	�wH�?	��bR��"8�i~�
V��#5��:��`"����\־��c�����>k?l�lQ�4݉�0���Oe;�xJ�|�tk�>�(���F�|`�E�����x����"�
��AiIp�ұ�P���lE��6
��'��p�P��;�T���q7?/��=�$�e,�,�M�'����$b6>q)˰�����?���G,�<i�B9����v�v[����>�^%�N��>1��˴NJ�V��xS�uنI�(k}�1��!)��&���$�� ��9�ZXw�%��/����@"��8���o%Oo0,r�dx���:��*?���;7.r�{��c~� <��A�s��:�h���sL�k��6�;�O���$1Ç��T�h����w��F�aL�"�+��A�9w\&��eQ�@�JOAU�a�t�b�3�ʀ���;"��<L}����Ӎ�� ��e�ٙH	1���;�{�5ԍI�*L���FLV�1�Ho��m[��$cf9&���(G����)$��N}���樛�� 7�pt�Hkk`1Ѵ���S�����3���!#�ޡA:��[����ъ.��fj�����,jmÞ%Vl���٧��)Lf�Ǜ�o�]4��;楤�
kV ��;��h1����[����Q�Aˣ��^(d�4�D���I�V}��tw��l�շe�BCj�<y(
��o�}�*�BY�8O�	N��W�}����"
��o���%F����d^�i���W�6�\�n{��m����1 �H��Wdd �	0�l��y�ՑM�����N1?)Yv(�v���Y����%Ig较� ��2�.�:�n��d�mw
>܄��]��"�M�<�&�-��X�=�͂�g��	�mr_��S0�h�S꭪ӑc��򛶡���i@nըrO���@�Ƅ��`#���Cb��� �>���TlPX�l����Z3I_̷�sq��^���=�_�&�݇Zߕ��A}�Z�k�����s��to3�&w>_��8�6�W��l����!���s�+��ŋ)քj/M�B�����J�����1'�q��(�"?�`��M�'����P��@@'��L������?Y��܃܋���4-vU���'�&	,�V&y�Y��X^�O���L4�V٨���'G�~ߡ�����B;��F�ן��`R����'�����f�s/���y�տ� ����M��puQ`��x-׸N�"������������%mW�zjk����BVwz#�ѵ>5z;Ї�ĝ�Z)̏�z'�4B?1��~QTr�G�"����.4�2c�@:��z�� �`�i(��*/�6�:A��.Ȥ����y��W��i�P�;axO��X�C�D����R0�o3��Y'�
P�=�-C2\��}?Y��UGTKܧ�y^�f�P��Ku�����A����,��)�\��jW��
�^u��wG�xY����u�چ��w��[�kw�;%���p��||I�:҈�n��jS��	�����Ėr*u+=�^�!�c�J�����~�0� "�ҵ�JNF��t^�{RC W�p�a��xf���[Y_1$�c��0ܽ����f��k�����I>��~��9J-�5�<�b ��^�駊J�W"l�V���_y�����	�9gwB�F$�8���*#l+�^�{=_�
d�V^��W���'P9sM+��X�lu�s&3��C���)[Ơ�D'��9:�X~�&apL�ןE��i>�Ƥ��@4lر��RK �݂�s��~񘪛eY7$������.�l ��-E�޲� ����z���[�����fo�ǠT�ா�� ����H&ϰz+��鳌�2�+�aS�
���G7U�_�'�[�15X�,M�@��b7���<��y��af�SfE���.��O�DjR��)����(s��s`n{-�|��+.���<@O�0_�{ƈ�l)�"�{� �x��d�s�daU1�Z�>S��*2�~����vy���~J�⫢UT�#��'��R&�%/�չ�4������Gc�{�'����j<Zǖ]�x/)w�4R�L��	���a	~�Z�!M�<th����Y�6zZ�v���j��\�	��N�Zx�>�IZ�����j'� �[��{�z�\Q��WQB���b��P����h��i5��n�L��&�d�����d[D���wᯍ�J�iT+��1�U�lt�X(a����(S���J/��9�\�e�����{��0;�b#���~�'�(��&q+��2|2Ҥ�CI�y�6X������Pu_��'q�uK����Cέ���;uK���L�xW�^r�AP��~�/�.�X%��P"jK���е����\���%�w�f���Xy��}��c���I�u�����%�t�f���<p�����kx��D���O�D���" c��It�-MZ������Q�1���?��HY֚Fߩ3?���1���'}�M�f.$���ٯY6����ͨ�*�(�I��b@Mf�� K"�1x�%+����<�a%7��T8DM�'��mu�aI��u�~�H���c�R<�ձ,�	����5ݍ<a�R��_W��^�e%gA�����7��v{,�x��3f5t�R����g%Xl�`T�ޡ����A����t����&떾�H�)��/F��A%细�(1=i�Ee34�y1ε}�r�g�$��&�(B���i/���C�Bh�m�A,�I����	6h�F(��DM��غ������\�c�O��i��	d�~e�ƽ�ϱG!PΚR��k���>���A�3�Q�������Ϯ�ԋ��!b�`��ӷj+rܱk߁�>�n\C3MP�6���"�
���b��{��G$��O�����6	��3�gH�_(g�2��	��1�����e���-��N�B]\)t�ʱ�7bc�,�"�i
���}�T�r]��"���/��.B��7��u.꼍(O]�2�bM��'���=r.Wɠ��H#����@�x�����>H'�!z)f��[�ǌ3�~+��ԫ�����@���\,�R��X�|(��Bb�������y�z�ff�rE�UG.�.��k�PS�g�s����4�{�|�ŵ.�����@���_�Ɉ%,�)��{�;� �3ͅ;\���YU��_���_��Y|�?����yŽ⤎L�#��U�;�c*'""2&�:�/��I�5m����G�H,�{��a<�q]E��/
�84S�F�<��+��	�hʢWt<�*ῂ{���w�g��-=��?�	v�~N:VL��C�ZA���B����|�^{�6��1���=��,4��a��x�h�:�5���l��@��a�3����k��o��CfJ�+�=���s���B���Ʊ��z`���E��JPί\$�\N֔�t���**���w�C4���~�Hw(�4lq���2��祿�ITN69?�����y�_&�qkO�|)5Co�½A&K���L��`����N�;E+/�	X��Y!Kj�wж�n��Y\�k�%��ftI7X�K}h/���B�I�q���p�4�%�d��]�@AV��=����>��+���ăR�cbwy�~-$X�����Q�/͐��٩cߚ�5��e��X}K��N�}�� fO��z��5�/4ϫn�{*��m�*>��c`�f��CKc��x(Җ��������a��ˇ�8E޺H��ĮJ���K��������$��R7&�-�b����~����RR �_�0v^j$�g���� 3p7
���,)�˴q�t��d���gl�DK��z�\�0A7�ct[gͯ����岝�Jz�/� �A���Q��f����	z�I���������x���]�(�8��*���nC�C��m��,�D��N6�e()�/MQ<���H\܂�>c�����,�H�6(�~Τϒ�Pϳ��Ҥ��%���>G�3wܘ����Ϗ�ԌA�!��`M��4��j����R^���gn=bMQ~`6�nF�_��ke���oa{��U�Ҿ}�m�� 
�6*�8tCIHS�7g"������1�SV��FL���N�C���,]�r��K'��؇I���r" ��jX�����˕g�]h�~"w[Q/��B.�7��ȸ4���,3O�%����{���qD��e�7�_C<����v�cȭ�J��v��PD��~��T����_>���0�������V��^�$bz��6�������ფ����
�������|돰*p�y=�7c��@�����Z��`��)�0��R�0�3���u�6�1T�� ]���r�%�� �S�RYB[���d�a�Lma�=e��:���I)���x�0~hy�5:Q�񬑬VQʛ$>p;~�}��_g`�5y�;�X	K�Z�ʻ�@Sp�'T]�(!�r�Du�>D27g��`�����=S�K����!id0-xD<   Z   Ĵ���	��Z�RvI�+�� 3��H��R�
O�ظ2�>��j& ��ش�?A��[$���(�E�r�c2��&��s�}m���?	CY���'��6O.���.n_8d1�I�TT��k���A�p�ش)iqO�a��d��Móg�$4�H5Ѷ���=�
��F@yB�@A���#^��$��yލve��=�(�*�E�a2����Ȍ��X���=3��<�A�B=Z�'�+G��� (���p��n3ll{��lV��
��ۼ
���.	X�|�T���I&c��8�DʣWP0{Ŋ�- �� u'�i���K1/Cc�	3i|��c֒|�g� W|�Z\E�zͫ����	$�ɠ<]�Dd�I�(@���Q#����I����q���DJ��O�I�OZ�q`T>��5�B;02R5���>�W�5��➔
C��#/�u2L�?J!&���z�u�����"�O�x�#�] E5N� *N="�`��o\�a5�O����$A7��dD�)KNiұ�%߸���T��	=[��������`dH�i�Ĭ�G�Ëm��Ȑ��dĝ�OH�@��E���l�/��=ha@ĘL,�T�<�f�;�x��O �(��C�rR&�!���#�^6)��((���8�'v���>����sM-MT�逬��\[l�D�Py�0�pi���i���������� ��%�"?�$T�tCJ�s%�$ w��<q�M ���$�@F��#��O�<�'�Q����34Í6~-��H�_�x��?o ���p�_]H��O�#�(�ñ�3D��u�   �                                                                                                                                                                                                                                                                                                                                                                                                                                                      P   b
  	  �      �(  �0  7  [=  �C  �I  =P  �V  �\  !c  di  �o  �u  ,|  ��   `� u�	����Zv)C�'ll\�0"Ez+⟈mZ�YL�I07)��Dw�����c]f^�aPnӗ[��9� l��t�(�iҢJ�1��ݱ��׏X<X�;t���'L0+��PD4��gŃ\�^r�e������٬8R������.^�Y[�&���hq��|I:Wj��|�D�LE��H��������N^lq���ɷg�*ٯ(�>�ش'�����?���?!��L��m����3@m� �p)eY����?I��iU�ۂX�p�I*rY������SP�[��6v�PU�?ȵ���(�'��'�BcB<�M;7O��T,2kB|���U�"� �@B�<ғڈO�7mI�e�T�"'����.Ы?��p�'Y��?�I"-�����xҨ�~C|]�3���p�f��)��?A��?I���?���?I���m�1���N1�0ّPK0Zt۶o�On)��ڦar��M��xΛ6�kӶ!o��M[�}M��1c�����9��V+Hv���d��ȟ�m�bn2l��h��M	?Z}�yC�ڤ*.& �����ЫUy��Uo���M��'��G'E j�PqІ�PՔ���G̋�&}�)�n��kJ�tG�uzq"�O��x �����@��%�p7�Y��۴Pi�Q3 �2Ɏ()�A��W#�A"I� ({P�ʒ.�v�d��Tn��U��#eI%��.�����*!��nP5k��ٹ$��$dd܅b�Cx�p��ΟKz�7�O���شs)�]Ce�%Y�%�E�z����'����hhz�$�X�E[�j��U��� �D9�"#�V���eDן0�?I��-��H�/ƦJ��L#J�?����'�2ðE�:7�,��`Ѩ�p0�Fa�'u\�+�OS��Ȗ'�2�'e"JoA�d��E��'i�&M��d�H�޵e� !
y���7�/)]ax43k�Ѱ``Y,)`�I���'*�0҆ �:�x��T��dUn��
Ó4������'� yC&*�)Q����ەW84d����?A�����(�����
L�"� 9�������DA�'�p��L,X7j��	��h���1�r��A&'O>��;Zǀ�%P�Ve;���z���ĭ� N�Z��v-��9��@���ʵ��j��:�P�g�G�lײ����a�Ӥ��#�6`Ss�W�4����ȓMp�paF+.�&Et �ȓL|�9��!޲^��*s�G�|� �I�&�"<E���{���@^�26}b�W�Z"!�?eǸ�f��9 Э��@��*s!�$W=E�� pBb��s:~y�O)W!��϶F�����Y#څ�c�Ӑ5V!�d"0T���㬁�K	ڀJa#�M�!򤏯m�F]#���V)��M:b��Ii����s>|Qr���(�hħҠ<�!�D�& �YHW�B2i�,�ۂL�!�!�$S�_�na�@!Q|���7�!�Ċ�Rv��i&뙛qc`h�@&T!��VC�<�;�H�}H���fd�l��yb��7yJ�7�(?�TE�`����^1��`�`��t�'3b�'�Ҭ��yBv������t��XBaƅ)���qk!��ǅ�<$�0���� ��)�1L�8)9�����$=C�Q#L�~d�(�Düv$�@*T�,2�DH��D�DW��'B�'�P X`J4=���&"��
vX��^�(��L�S�Or\�	w��$����ا4,������ D՜��7H� 8�v��B#��?�/O�\�q�̦1�I�P�Oq���'�̘�f�[#���adf�'%H���q�'��@�wN�Ñ$�.+`���FW#6�PX����i�it�=��,��Nf.�#S�\l�ɤ��+d���'6��4�á*��"���L�j;B�Q����*Ȯ�h�Ò���D߃a2�'��OW1���SӈSʜ$i6E� 22�s�|2�'"az��0�~�&�M�����[���O>AE������Hq0I�r�xQ!��8}��V�'I剾WM����ȟ �I៬�'3x-�"�Ձn4rh����v����c٢3�����O��2�
$=Q1�1O�+�J��KC�m�X% &L:-}�!r�G��~U��Y�R�t�����y"F�,NXB��Ȩk�^�3 *B<�?��O*��W�'1��'���2�b%��T3`��e��F4a�!�$�^��}�0�
,x����%��	�HO�)�O���<�ڒ��;��}��l%5���ǃ�,h���'9�8�ag�^	��բ�M`�J�ȡ�x��lѾP�gG-�P���� q���	�'ֶP��	�t<4z�,pI�4��D�?�	�'6@!E�2J�S�ą�g�:EA�'�R��� �*S@d�xRc!p��XJ>���i��'�1i#k9�ɋy�l��S!4�BѳТw�V��	˟|�	xL���I�cԾ ��E�'�� �ᙳ�
2h�	�jR�q*��Rb�'V�9���a�
�rB♏?�6�Ț��0�A�g��X"��4ax���?����䕀C��Hѵ�C��9� 
�,��'�R�'��
F͕�~����V/	1d.!X�l�I�
֪�˃GU�U���g�?a*O�H2�����&?��O�BA��2�C5һr�x�Y�n�8��'�1�4
�������]%��uBE�ޢbΦp�J?�s�/ݨi�t�z�ύk��e�ՙ>��d�-� 5��Z&O *��S�dKb����8�t,G���]��nE<>*���M���$�
y��'��>A���(�Z��1T �I7I�4b��a��|�hb����P��郮ܴ�8DFRf2ڧ%�f����38Lj��@�	j���I�'@��'���� Kv%� OR:f�5�AIÇ8�$�Q$�Y�>�����?��b>)���U�	��$N�[ɾ�2�_
e�JPbRLX*M L���1S� !��k����������l%J�'��e�anG�l��8s�����`h�i8�7m�O�����O���䟎��O����OR�Z���a�nY��"Z=-�j���a'T���c/�XrT��͊e"`��]�4���D�ϦE��Iy���~X�`�A�\����@��%׀�:����'@r�'xP֝����	�|���HM��u�[;���F��"�h���B�H�d�Cn��XĆyX1�ɯ.t�E�S#�6X�IH��`�4���IS�	G��GF�D 
�KJC���O�E8"h�!���D�B��h�����'��'���'��O��h�cǀ!Fؠ�MȻ9et(D�$D�$��I���K��^���a6#%�$���-��[y��[~��7�O �dW%9ՈXg�*��a&(^T����?9�CL�?����?)I��O��h���<�w}�q�Gj���:P����+�TzÓ{wDm9�c�%\����3�� �jPJ�̐�D�^�Z���lz*%��,~�,����O����ͦ����-�R�G].8A��b��
,��ؗ'�r�4�Xb�@+�%Cr@F`ڱl1a( �4,;�OLoZ"�Dq�GS�(ԫ�Dǅob@[ٴ��DuK*xo�����	y�t C���Eō��!���t�nX��A�H-R�'�.m94i�=l���Ot�'���F�P���P�jM�J��0aP�x��	
�`�2��(n�,u��\++Ô#|�ң1I^�t�0FR�I�}(��|~�A�$�?	�_�f�'�O��ɀ+z����ď��3����t�'��\~r�ёX��0��I�9IT��*����M�³i�1���Y���ZdL���+������'b������Q��u�O_늅(��P�SV:A�բ*D�����2�
�E	o��8�+D��Z���>��~�0�3*D��:���$p0iP��߃8��0���2D��{��D	�аb�^���p)2D�����ߦ!bh:�B�<b��s�<qV�t8��`��"gJv��eA����-D���Rn�;Ni�7��un��{�?D��`3�Y9KAx�[�ܳk���{G�>D���Q�ǟ��9	�����F&;D��0Tŗ 1<i�	ˎG:t�
�,=�O�	�E�O0 �0����ce�$V$�})1"O$i���-i�@�x�e��>�!!"O�]�a�N����t�Y�e��ѓB"OB�r%�Ǡs��Ҍ���4a��"O�0#	�'�Z �FP�B��I�"O��a�G�:\s���4&�+����L�f�~��g�@x]Y.ЋK�̰��La�<����bS"�hv��/�dta��YQ�<I�c~, �
50��R�<�VgF�XaZ����CFڶ� ��K�<�ТY��AraQb����3��C�<iKQ��ah�-��[�b=�PAٟ��N"�S�O����/ �F�Zmؓ��Sg��H�"O����(� Ht���1DLt�{"O����sS��	�B:�c�"Ox�Isb�~��m�e,ΉJ�L1��"OP�acC��2����.4�:���"O$5�e�#� ���H�>'��6U�Ly�	9�O6!x��4W�e��	ŏD��T"O� <Bub�c �$���� /����f"O&���8i��ũ��9��1{�"OI��_�Xo'b�	9�9"O
1��EF;x��×Y���`��'$��'k�PG�4Q�Px���syt���'),��Sa�Z갼���	5gy����'�Nr��	3�	�@Տi��p�'�0��ƥ�I�|�^�t���
�'o�����;k\ à@D�6(3	�'q���$�Lv���2#�4S�p�ʈ�Ĝ#FQ?�[ꗸw��a��䎪pmFU�Bd3D�X2c��H_F��䍶@��
A1D� ��H'4�����/ǔ<����4D�XR@�߻v|�0�,Y�_伈���3D��qSco�%�U�Y�_n� bW	?D����P�K?��U��>nE�`��O��C�)�'C�hBc�^�q��tB��ڌ@����'����@˲��$�Oś3j���'��R$dѪ_���!�v�lU��'y�] J��o��dX�M��j��A�'�lM�k°W���Sw�Q9a��)�'i��j���)�x�%,�|-O�}��'O��ViTM���Ql�}k����C�S�#�l����+d����_�ҕ��E�(("�S%=� t��J?ʝz�H�@��%3�

v��ȓ����a��&%�>�bsL�8�p����9Gp����W�^���@�o����. �sm�B�I4�u+���>��M���^;ĀB�ɻ?�!��j\�P�ĝ*��Q"A"C�I�y �Q�Nt
�ՐFN/D�FC�I&��5a��Y�NCn5e�̪\u�B䉈!0�#&�pcP��w�挻W�*ړU�x=G���]�an`Q����+�ܙ!%��y�DP_���%L�(�.-P�(ʁ�y�'�3�H�h׊�B�Q�L��y�h��W���:h�5`.�A���
�Py"�
1M��eq�NB�C�d 0D��<i�d\�� #�<R�1�d����ʗ�1�S�OQ(�HU����<�~���"O,tvA�#9h���V�?��="A"O@���W�s���Sw���h�θZc"O`͛�I��#:��1��\�z�s"O����Gq��X���*}b�Ҥ"O�8����j�,�����k�CRy�a��p>��ǸN�ՠ��7�L@#�o�H�<a�힗R�
��g�3_��h����H�<��Ɯ4aLZ��"��9x�AAD�<�S�Y8^��%���-I�*XR�$�A�<1���jU��L�x6ԅ��@ASx�x(#���T��C�U�4eaC�o������'D�HM�K60��OG9a�	�w�2D��
�&T�~"�Q�cÄ:y�Ԥ!�n/D����I�#���f�ƅw֢<��N/D��@���_��Z���	"H��a:D���PǚS:ֈ{�Fj�4�ۃ.ړG��)F�D�
�q�t ���L�n��Pqt����y"��LyԦ�m���*c!��y����]�aDB�^��A��]��yR��4�y'_�1��A�a�/�yR�P'M�j$K�
��k�� ���,�y���`��\C��gS���r� �?�1�J�����mY��X�A!x�sJ�`Zƈ���#D�\��Ei�ܬ�u"D�s�+�.D�� �A�EֱU��D`ƘQ[0$Å"O, )�瑍b㦍�@qX��!�"Ol�W�Ca��(Ɖ[�g��4)�"O|�!C��|XX[�)�#[�	 �^����>�O��A�됨4�Ҩ���a�-�c"Ox�+��P-vZp�0g�w�L�w"O틓b��?H�̘��X�>��B�"O@���"g X�%���e&�H��"O�1+�.��1pv���ݙbsƱё�'�8L*�'KT��n�*@c�"Ї,�@�
�'���e��FY3�Ƞscl4
�'І�8����*�χ�E�l�x�D(D��-C*^eh�Aa
�hȄ�s2�9D�`�N�6B�\�&���!�"=D������A�Rp��L� Ύ-�D%ړj��YF����/Rj�a-1��H��I-�yr��4M� 9�#��)��V��y�J�U���q!P�N�uK� ?�y�bO3�� Q�-?G�ĕ�)O �y"��q�!��S�<u�a���y�Z8:Z�A���1e���擌�?YT*�[�������v" �Q^
��g�L2��,*D��Ń��&�x�3�	-Cb$��qk&D�ڷ@H����RmȘ��u�%D� ��K1�� �i�Ym�-#��?D�4����䦰r�i՞Eˬ�B��"D� ��%\�S�uY�cѹ%D�� '�<�!��q8�4Ȥ" NGH5ѷ��+V��@�8D����)O�����:W���0h7D��8aF
��]�Rhˏ��pR#D���c�.D��@9�(^aj��!D�$pGi��O��n:�F���� �O�H�O�T��%�Q�n�Kw�	?n\�"ObX�r�	 ��8
�`١sH� ��"O��I���V�А��3>3|���"OZ��&ꈇ��t��x|�!*A"O���oK3=*�X�5v��"O�Lۢ*�#�̥�4C�J[�I��I�B,H�~���C
q����5FG*b�U!��}�<�$����]s��Y�U*�!KFx�<����;/�	;5%��/�|�Fz�<��cӇaT��b��!+J�#Ou�<����Bn���R!֞E�f�;��r�<`�����@e�Ș�дf�d��g1�S�O�Hz��U���2�D�gEPHXG"O���C��$�}K��>�l�Z�"O��A��)%(�U`�-��B��w!�D�{�����f�24��Pj����!�8���Q#�+�����x!���_b4M�v&
J�D�엗E�	&W������<9܌��T�ӱ������!�$�{W��Z��d,�+��":!�@$l�L˶wa%&�&x���3�"O^|�"*K��$X �Õ8��Tː"Od���`Y�Qqڙu#U[�Ȁ�`�'c6}I�':���S@B�Zm ��/�90w�Y��'��8A��P�(t�JW \��Y9�'릹��+ѥ��	��)M�!�'�:`Ra�!ҹ�	�Bά5Q�'�"̈% ϐ�|9*t�.� �s�'���C��� ���۳�ݡr��mS����ZZQ?ѡ叉(=YL<��p��!Kb'D�h0��9w#��&�	�gL\�IU�2D�� �Mꕻ�NȊ3�DM��k0D�� .��ք۩_� ��\4c�� "Ofȫ�,�~Hd!�'F���f"O�԰ fی7�-��o0Lߊ��1�'�H0�����]��|�CN��1q��;���*|�0 ��M�H���
��	��Ề @�j�Y��:�����%� r
�"�-�f�p��ȓ#x��!N�'��: �W(y�E�ȓ�.�����O�*&��%�n�<9�bY�I4�`F�}�(�C�-�ly2mƖ�p>�r�'M��b lG�DHE;s Tf�<�� �%��Pçj��2��'�X�<aq�L-%�q��@�ov�z��W�<u�ĺ[ٖi�v���K ]R��O�<��(ȫ1A��+��,� ��b�fx�D!���� 0q���qQ��#D C�{W���r�1D��� �QW-J�sJ�2�`�0g0D�<���^[̸!Wf���..D����F�;�h��`hA�d"��*D��)D��a|2��_�]Tr|Ҳ+)D�T��.��S(���F���7�(�]jPD���R�,�����#T)2�X�'�!�y�b[9~�T�V S+V�b��C��y��5U�8Ao��R���!��yB�^�	z�I�ŋ,C�$!� AŲ�y"�O���	�><Y�7�y&�HQ6�rBA�:L�S����?y�L@���� 1�
�� ؀�)�h��l\���6D�4K��>m;b8[�ݗj��3w�2D�8ڀ�@���1��ݤ}��E�2),D���Q�ҁs"h+W�׭"��k�*D��z5/Ӷ �i�V�Ӽd�X��&4�t��FJiy,	A��#���2�G�ǟ��O��'S2�9viX�<9��OL��]NH\�fJA�$ZrQ��	�ln���Ob����6<FP��$�Z^�ŋ�ߟ���Ɖ2PN��	�0-��x��#>a�D#gj�500�ӻqpt���|Dיm|t����Q�$���a~�'$��2��?��4Hȶ_����U��8DC���*���O����I�"a��]�!�|8
��Bt�}rL�<)r�/R�n�#2�:?%����@fy��D���'�Y>3��Oϟ|�ɷ(rr���G�|A��"��	hl�I�F� ��bD"�4�E�@r��uџ�c>���M��ag@pp��*&T��4�b��b5!�P�t9c�͢}����JX��H��H�];<¢�s�KB<��A�?O޹�S�'�Ҝ�����=���
�h�:��y�aHн�H��ȓt�$�(�61�<A�Wa]�R�
 E{��"�'qVL��������×l�pڦ����?���;eXq&�U8�?���?9�����vqj\3d�
�]�Lh93D�G��9���5tq� ���,���ې���XR�0�p�4 N�%*�� $_2&m��p lA�k
4��!L�<,��R�DR��.��d?������s�����R-���䬁�I� G{�<OZ��hؔ�(��9D6-Ab"O|q*g� � AubY�g��e�!�'��#=�'�?�)O|�c���L9�)؛x$n�y��9&ڢPR���O��$�O��$�N���O2��� ɒ(�I�&��B�S����፞^����UKޤ/*�@p��OTHWC	�J�|� �����Jc���f�`�B�&��iЭ��&�G~�g���?'I	��pu �	#���K��L��?I���!�Y��t�ӫٰ@��K�"`��ȓ3U��0ʌ�b�8L��Y�~��d�'qt6M�O�ʓǺ1��S?!���|�I�9��t{�iƾ^��Lz��ퟠYƥ�������E�C R2��J�ˏ�i��tB�\3F��.E7V洌�%T�
Ā�iW�a��䑅�Q�F�Kdf� t�q+sk���u�Y6t"�S��B0}��5)�o��шO8���'���)�����W Q!n� ��B�*���@��dJ��#=S*@��M��I��2�ON�':F<ZƪH�P�a#Pǝ�'$`��)O����Obm{2��<-�����OV���`��Emp���
:r�b��/�O�8"�!Z��p�1{P�����O?�#s�!�Π p�\�Ak-���a��`���7w�e"]):��hF�� ޴ �PD{�iE?Z�Cd,��y"kE4�?1�����䘟� �8����PD��f�ݓP_	�"O\	��� L�\��N�<�"�I��ȟ�HW�� ;g^<@h�?#�VE�@�I;�����3�ـh`�҅\�
�C0B��:e��%4�hQ`�h�F����ѧw�h��ȓr��$�����d��rNN/xi��6(l�;�̓3j(����Q�Bܚ���+���UMZ������%}��d����3TP�3l̟F̅��.N����$^IJ�H҇NXiI�v!�]U�4(���%$Юpj�f�2d�!�$�.Z��bB	ù0��5��eak!�RxS����[��	"X!�D���BK�{hT`"�џ��g'���MKK>�ǫ�'1A����� 0�<�c������O����O��#�� 	Ip�)e.H9|����KW�p�@�kW?z*P��4-6<�P蔻^�Q���&�&C*�i���O/8���sآl��y�V�A�l1�H�!�r��3!P,\�Q�����O��Op��p>�:�FY�T`QN=;�"���e�O��D'�)�'e4��9��J�*J����sP)��k��	$.@��N�G���b�Nª<kx��?����?i��4��LR0k";����S�I.W"�����2O�=q5 �`U*'��*gdT�C)A`��M�O<	�,5�ӕjf 0��R\pTU�`�6n��8�D��6��S��'h�T�ҷ1�`�!T$��f�)�&�x=I�O�OL�ƙ>q���%�ԒfE_ I�xTs�)��<�Oz���h�󤈩 ����ga��R9��4$�$	�Ќ��>��>qb�_z��RK�4�U�{Z�]PT*��i)��C�$Z��?���z��I7>K�?ݣG+֎6n�:r.[�h��qd�ԟ�(s )}rC5}rˉ���I?�M˵�P=Zȃ�}&|�iGnky�OW���ɬ�ȟ\%�@��'�=��IǊ/�\����I?Q�͙i�T>�	'+��:����U�@6/�h�(��@|P놫K���dРIl���Of��=O c>�R��Z�A�F�
��̆()�D�O��A�'��p�O�s�0)B����C2�3�Xa����*Pyp#�O� [	��2xp�&"԰ �<d�FC��~]�����|�1��n���;fV"¾hlK�.��|��=��B�
$�Cო"��K�ꓑ?�)O����S�DNG�؀�MC�L���1�ē�hO���$���>2�]Yh�:X���"O��z$g\�N�!�a&�2RB�;�"OvU�T�-n�0豤Q�b�EPS"O��и�M{wᗑ�P�*�����y�oņG:X
���-�j���yB
��X���0va�. :�p�	U<�yr�\�=��E-sD2�i��	�y�@@��se͌�eL`"�Q��yrΆ$>N�((�O�N�X�l���y��6S��q�2"�4>l30�
�y"+��z,�ނ��r<k���y�P!x]"��~�lpH��+��'h�QuD��V�ڔ�81툕@��[[�}����9�0�3����9��Dv6Q8S��>]v�z�,��)'�@ "����r&��!���92C,��y�n &�uA��C5+����� C�@&���"a\Ju$��Oc예w��g*�`� �,�P�OB��JU�8���4N�7,>�	Cv"O�\ ��7�m�sB�/>�=�"O�! �F8�4bڴm��4��"OLm
u�+��r�C1+�>4Q"O$ՁpO�$!�R!xT�Gk��P�"O�� ץ�
�"|�3o z}R��2"O��3��x&B����&j��`P"OZ  ��A��P!M5U$Y��"O����L,�h�D*�1��8�s"O	k���]�����ߵ"��`��"O���+ГI���AE���v"O�;��L�P%��hM�>���)S"O���a�ܬ5��@e�:?k�	��"O� �����54�@�����|�"O�uc�g�;��8"fe��Yc
��"O��I�$F>l_���1�TI��B"Ot�B�iM�4B�E��#7���5"O D2�#��no�يQ�E�"L�"�"O|h�F
�E|Q+�A��2� {�"O�@��Ӫm�H����!^���"O��+��4%G�р�X�$Ĺ��"OV�i��	�
N���O�1o숝Ó"OZ0���*v����NU�V�8&"Ol����	o�,`SO�jCf	�#"O��!�	�|�.���V�/3��C"O*�P0���G"jc�R$v$v��7"O ]�#Z-[��4JT�'G�p�6"O<�At�+�\	A�a �y:b"O�	S��Ї4	R�i"�ҏY��T��"O��%�њ`H�1�.�05����d"O���l͵Y���t-��M�QӦ"O�8�p������+�$y&0�1E"O$ ����$?���&���h2���"O�IQ���YDNu�f�Y�T0D�8"O� bt�D?sL<I"����q�"O�����/dkn�{e	܅D�t��"O6��ҮX�7	��J��#��U�c"O��5��*�Z��be�(��&"O�x��+s�&e1�Ę.���Hu"O�� 钑uZ�e*�"ݝ���R�"OF��+��<�0���cW}��x�"O�D(ef�))< Ib݇
l\�k�"O� c�F���TA�
J
5c��"O�
OZ�+nT1�o�of����"OH[�A?2��"eOt!�"O��3s�߇/V\�k#m�/N|���"OlDQ�l��W:4]��k�j[���"O��	q��7��x�#ʁ�=@`���"Ov,`1I�)%�j�9vf�)g/�q�t"O��ap�9���X�b��_%���"O����H�/�� r�!@0�}�W"O$��Rh�+{vD�p��O�l��Lj "O$L���;eAf0kR�F*o�h:�"O���!W�Z���Cƙ_�d�V"OH
���b���{�"ӥP��aa�"O ��5(�aH2D9�At*��"O~�c7}�0����5Pm@R"Om�l�Y!|J�����	�"Oଚ7�؄n�~|��a�`��kB"O$h)��7����P��m�u�"O0�s��ZEƺP���S&��(8�"O�p�D�	D~H��3��%����"O�%�!�b��h�b6q�Ƀ�"O,|��H߼
2QKJUt.�s�*Op�����9}pB�� ��BP�y	֚OK�<�m�&[��٩A�ˑ�y��8^+^E���U�F(:�o���y"HC����J�0M=ļ�0 ?�y��!'�%�u���@=�$�(֯�yR�A�pd͢�lռ4>�l�G�	)�y"�(C���Cߙ(U�� Ĭ��yR/�
c�4E9�� di���y��>w�}q։�
�c�L��y+����d5e߲5�@	 s��yr��Fl�ڵB5 ڒ���1�y�$U�><��/æaqb�S��S �y��-.��\a�D��\�v\����y
� ���$n��Bh�Z�	H~��w"O�dxң�29.�LY���ߪ9�"O
���G�)�`��@K�8��0�6"O
!�)ŅF�ș#�i�a�VH�"O4D�7T�({R�Wnܲ�H�S"O*��"˖�~@$ ���V��a��"OHm�p(ڟ'ݢX�����F$ZE"O���G��3=��!�%K��)�"O���s�˶3�� 
�#� ���a�"O9w� 	�����/��-�"O�H��B��P�P��3m�jE#�"O,�#)b�2���b��a�Q"O��(���>qD��*��K�/�2`yS"O��Co_�]8J-����"���Ag"O%ѧʊ���"XY��h`"OD�ɴǍ�p�&;u����P��"O��ې���0Cj�Jp��=���E"O���Q�� ������;g �-�`"O��`�Ò�+���5�Y(���9%"O\��P�14���L�,E9�"O�l�$b�=F�@�`�ڬ(٤�Q"Ohr�kD4aF��j��"O�izF�G�uH�E� <96�0 "Ob���Z0Nq��cCǣz�I�"O�P��<1�" �5+��9p"O�b#BJ0R�{ӡ��F��y�"O�Qh3�Q�J�D1�7�����	G"O@����V*"��9��)�}q�c�"O&�ۆ��?'x8`���fcH�7"O�ڶ���8xR�@��I �Q"O�ظ!J	r�|mZŋ�2���Qb"O4��S�L�! ! ��M>��"O�!���s 5
�,mV�9��"Opq�
Pa2����J�W�dxq2"ON��T*�#q�&ph'Iۇa"�K"O�L %.��,"�i��IZ�g.$x��"O.A�e ���^5y⑈���"O�-X���.�A��_�J�|yD"O(��$�8x;���l1x׊Y�"O���O	��Iх��Պ�+�"O☠�D���
D�Gj9Ϝ��&"O�(��C�B��bʆ����"OT�;4��~����h����Q�"Ob���+q:m�����:D�a�"Op%҅*�?mJ�	�!D�I7"Ov��􇈌�ddaD�G�f'��!"Ov8�+I�=��x �gي?�X	`"O��aNQ;@��F�? ��C�"O����f_�
�;&'N�45�"O�]j H�(;�V�i%%q@�5"Ot��0+�w��"��WiaK�"O���+�L�z<:�`�4	��m3�"OX8���VN@b��:>�<}��"O
�I�f[ /���4d�(�h��"O���"����mseɝ�Mrf�
"O
E���W'�Q1�U�en�	�r"O4�B蝬2��YA��`fp3�"O� �G9Yz�� Oy-B�;�"Oʅ�i�~<L8@�@�5*t�*�"Oĩ*���/9�DP���-'N�c�"O`QB,
�˞�SG ٛ�L;5"O@uB��ʧ#�`��o(Z�p��f"O艂�ǁs���0��v�ڜAw"On����HtTLq+l�+�Y��"O� ���Cm��S�R����Tk���0v"O�<PnG$��s�ɒ$�r)�$"Oh��Չ́\��c闫#�P髕"O��� C�67�U����:��A�"OZj��B�fb��4L<$r4ѰB"O��r����x��b��ݸEc8�"O"�y!�,reXq��h�<'���J""OĀh�
O�A��	Y��E�o�4��"O�u@c-�Kju�F���V��"O�Yx�%N�Sf��ɦ�!-f8���"O<�X��+m\��� ЖD��$��"O��	�B6y@��T���u"O�ȳ���}R���p������w"O��3dO��j��:"��{~ iaE"O���a�'[���[ �Qc�9iF"O���1MFe�4����f����"O(�X`FO�`�t�J@�N`���"O�%H���	�tq���&.8�1"O�sW�V-$vͨ�i�J*ъ�"OrD�Q�P�O���(B9Phy��"ON�H�@�P���
J���1w"O��T�M��j�be��x�h�u"O�"�ZIN�$�O�`��KC"O��s� 0֢�sh@�*L�8"Ox������o�#�][j�Z$"O�9B�G � �ZMJ�n�-%U���D"O�Q����
��a��ЅDv�*p"O2IJr���k@�Kv�Cg����"O.!pA[�P�V��u�Y}�\jG"O4�j�#��^X�Y��"|�yp"O\z�kAZR%��C��xNA��"Ol ��it�V��V@����"O0)��(�rzD�p �5`�ir"O�5���;-J���͓#N��"O�!	�� .��SE��;�i�c"O(�J X/`�
Q� �I�p&�� "O�`j�OҠ#�(8%�ʌ[r���"O�A����a�L݈uiˣ?S��0""O�@T�Ĝ�kp��j@8$Ӈ"O���'�=4�`�;���!J;F;�"O~]rd�npI%O�t6��@"O8�!���`���3s@#`���"O@�3�^8<t�����P�f��p�"O�X���S�!�% �._�
�P7"O	s�Ҙ���I ���(L��"O������P�V� 0��Gf� ��"O��`bѧ(rn�Su�¼(Z&\@B"O!jv��CL1s1��IEÆ"Oj0W�B�#0����V�v"�ac"O�Y�MмT�(�j4KQ�'jy��"O�)!�C�9e�(��$�.X�Q"O���k��AR�RB-��Tf�р"O@�d!Xo� 	:� /`� �"Oܥ��#(KW��!���.T���p"OzI����=£�ߣY��i)�"O�-�H����@�����,��"OĤ���Ԇ��Q���܅J������J5A�ph�%"�,�t���-M��'#�Tx�˕hUڗG31sJ)
�'�pq9eZj>�Y�&�(	�P��'A�y"��H!x�y��
�w��@�'hP�Ól�.��-��⍿pn����'J�lp3�
�7f�#��S�t�r��'��xQg������A)؅��'�@����&�`ti�6XL{��� �a�+8�F�`��9W�~�d"O|���� �cg؜����%��ʗ"O����͗{�h�3፷Y�j�"O��arØ�2��6�J��6�{"O���a6�)���s�t�A"Or�
��ٵ'��G�;JҸ�e"OZ-p$c
�X��a�f�.]*��hR"O���nQWo��ZD�;y�Z��S"OH��ℙRl��s�d^+���(�"O��Sb$�o�*Й2�Z�3��!۰"Otĸ��E(���q��y�l�*�"O@@�T�%iظ˶��$�J���"O~����ZTز1c���$pP-kB"ON��@��)�����Jy&��E"O�t��Ɏy��+��L(!��"O��SÆ�k��9�-�;L�fm��"O��v��y��I$��	��qh�"O��"R"KvVF���DP�T�yg"OL�K���n�ec��N�a���"O��٤���②�*�l(�"OT��� 8�հD�,���Җ"O�'��GL��ه�d�$Xp"O�$�P$�}TJ�J�dȰ7�����"O,PE�ҡS2&P J��6�|�X"O:tZ@�µ:�D���7�� �"O8�#&.ەc�P1��]����@"O8���W1@����ڣR/�]�"O3b�<u&����J�;�P��"O*Uö$P�,>�	#i�fGX��"O���STA�H�h�NF�80"O� 24f@�k(�ےA
I���Z�"O�I��"<�	���V��[�"O�7�=�8$��!A\P���"OXsv9�P�j��zN��"O�q+�!�9��V</��q��ME�<��.�Tbz5�!苭q� y!be�<��ň	�Juʁ�Єy#@�2���{�<�v"��;��\�4�E�(�WgEz�<1����u�B�ӓ��@_�[�!^�<Y��(���#���a�2у��TW�<$�,%��Ub�εe0D��S�<���Z�1�|I�G�k�AE��m�<Y�(��5�<=)S@נ�q�ek�f�<!G�3aQg�H �^�T�\�<	T�	FHJ���Q�xū�e~�<��-��@S�ѡ��ĵ]$�;e
�@�<�g"R�2����$EJ�Uk~�g�]�<�0�&eP�b�,O�B};ᅌp�<i3@�]�B���I4���`�Hw�<i���-j&�7�  E�y	U�g�<A���1G8��@'����%�R��e�<���0a��īS��"-��%Ib�`�<a�Y������ό�jѮ ��C�	+`Sqx��
�J�N� Qy"O���c�D�ށ�t$ɠ(��1�"Otݳ4iK�3�<耓�JX�萃p"O�,���X��b4	^=u��͈�"O�y)����6ܓE��g��"O�D���]�a-��AA�A9'���g"O��臬ċ2��a��b�0ez!"Ol�xD�
�L �O?fĞ�v"O�"��$�2�JQf]�1���W"Oz��	H�oF4
 Ý8.q	6"Oz$A�Kծm���
EG�2my�xk�"O� d���	��9x��G]=�t"OT�7ƔL��`e��E�!2�"O^����M
h���Kc�D�$T���"Oj�r�hĊM�H�;E!��MX�"O�lb���7�ް V�֣d�0�X"O^xF@XN��e�^�(�j�"O���j�-d9���TE&�J�"O"d�
NM,���E�
L��"O�\���+I�pҵ	�I���r"O�u:�*�fR��'�Կc��I��"O��2U
#Q�� G�ՓІ02"O�I��$��0oT����Ʃ�]1"Ojt�e2�/V8k$���"O�h
6Á�jJ� ��
�\�Z���"O4mӢ�Ͳ l��ǒ�DѮ���"O�q��NLU�Pa��H�w�����"O���.L j��D� !�|�g"O������7�\��s�\����P�"OXY��G�,�Hp	@7`����t"O��cPfҪC�P�h��z|Ҧ"O�!Y�e�65���YV�4�yE"O�yy�ܼP. 9�ُG�\�"�"O��D*i�"�X4��2h��m3�"O��jI��Gb���@�b$b��g"O�a!Γ(�PR��\z���"O4��- +%�|����w��\i�"Ov�pC�';��(W�J7:``�"O������2�� F�SU�M b"Oʘ�RH�q���(��l^��"O\p�4)H�2��a*��Q%$�8�"OF�O��o�}��aZ�gon�I'"O���$�
i�d Ȃ���uj��"�"O�A��ȁ�A�թ6$C'�6�Q�"O��S�Z08O��1Yc�d���"O��K�L�\:.@WJ��_܎��"O&�z���R�T�*�IG�]1HԨ�"OF���_GƦ=K�JH5����#"O�A�M�3wo���^�Y���7"On�q�\�
�<a2D����!�"O�L���M�,$�d�׫��*���4"O�a�s�T�C/l����Q�j��xc"O�ԩ�`Eg3Fyj@���PqH�"OD����!EС�E�$��v"O(�� ͼi(�`� n�&��X�"O�(�' ��C�ވ<�H@$"O*q+��?)�;�x��	Y"O"�xP"�2��U���Y���A��"O�Lr��"~*���	ٲm���"O�	ᯐ$\B�X"�i�"+�ʬ)g"O,�3�7x�^�����;a�j0hE"O�����(/�*�h��D�6�"O� ARJ�0If���΁nؖ��"O�}��$m�:�y��Ws��Q"Oh�������'c�� w��5"OB<��{��3��kH��"Oz��b�/�	(� �N��k�"O��J��H&p��P��m�q�@��"O��#�(�8-nā��&�X�\t�"O�<�Dnݼ)hL	A�%�>1Ŕ�`�"O����d�dڢ
� �Pݪ�"O��j���>@4<cf�1Y'.�J�"Oh�@��p̚&i����+�"OҠ�H�?4��I��Z�vxp�"Oj-C� �yW.!�'/� 
<��"O� Dl�gK; ^�s�CJ=e �$�"O�$��钹DlV�s��� Vf |�"O���ц��P	r'I�-� "O�+�(�r�a0 U����ڣ"OT�[��۬v8�吧��w*H�=v!�ē�C۸�pB���>cm�7�Y;�!�$O�a�$�� K�UU6UI��W�!�!�̟lU�t`�1&q��r��$#�!�D�~M4�a��7	Z�I(���!�ą88d5z0F"i���z��ٞA1!��J�h��C_5�J��c! 	!��@���
�c, �T�27+!�DM��quBμ8{�ܻ�k�&j !�ĝ*El� 9��[�0Y��ʞ(c!��1-V���Oz�h#JF�B"O�y�)��|unPI�ׯP�q��"O�ų��͌6��i��G"��"O@	0@h�$�z�Ś!��s"OZ4"O!bM&�*�eD�gdv�P�"O�|z���'S�ĉS�	�yL$9�V"O�e��c�*[DJ!PǇIE�hٓW"O��vB�>.�5 ��<����"O��p�"H�kڀ"V�J�o"n��"O6;1�L��hP�t��Y� ��"O��%Mؖ�b��beX.yn"=YQ"O~��v+\�]�q���dUh���"O���m0q����S�h��"Op(1�I�t�8y@"�I1E)���"OJ���˗a�����#��/��c�"O��rA�][��sA���+�"O��2�]!A����ˉ0M8Pi�p"O~��jB=g ��h� ]�)�	�B"O�eRk�=V�$�ՄQ��"OH8���Q�]V0��F�y	hr"O������(b����'���o��2�"O�MBSJ��)�ݡ�Ăxj�Q�"O��&�G�N]*`5he*�"O�i��JL0� @�π�8�>m)�"O���D-2 ~1�g!(Y�V��"O05��Fڋ}��m����v��hQ!"O>$�oI�Q�jS���.*��@�"O`m#��Ϟd%T���۝a��
U"O����>�rѹ'��?)��e�g"Ob����/$��E��ON�i��d�r"OBة�2B*� Wn�9d�dE�p"OV��D��2��\��'�&pJ�"O̅i�(z���e�d�\�H�"O��NW�6����e+b�5��"Oj��=K2��E��F՜]��"O�)��ñ#$\X��
u_�s�"Ot5`qC�9}q��&�&{|��B"O��AA k�ik���?$:Q�d"O�D�%��|8"�X%	T�}i:A"O45�EiM�G��I�^:F$�"OV�x��'pH^ٳ��@'H<�XQ"O�IY6!Q��4 �DW� ����t"O�q����ʴI�,%��=��"OV-#4ڗU6�)�	��T��u�Q"O�k壖hƌ�`�)l}n���"OF<#B�À\�>�qǪ˅A���"O������
!��;���:���O(���D�>���ђ�_Y��'ʘ�◂�^q�=�4j��D16t��'������T�Sܦ<;$e�8���'5��"��mx���B`ᴥ���� �TїL��] N���Dɲ5O���"O<I�c��b�4�Ȅa
?7t`+""Ox����wo��&�3��$"OV0���}�Hr�N���>!0q"O�I���C|}�0����q��p�"O�q9�g��`wR�jg�Cg~���"O F�C�)�荂�M%7|����"O�h�İt嘒��5c\��k�"O� a�Aڏ;k��Ihh���"O:E#PGޑl��ȣ`/g"�CU"O�a�%�j��
P.�XM�4��"O�%��C�42��JO�Z��{f"Of��L?A|Y����O��0�1"O���]��F]ibjq|z�C"O��d���;�ʱi�b�Yi�P8�"O��B�ŋ2K�6��p�=I0j�
�"O ��V/[�H�I�0L~���"OD����O�g����V ��D~HK"O���׍
�~��]�����4Q`�Ȳ"O�"�D�u��(�a��>N�	��"O�|
v�Y1�,��艹eX���f"O�t��H�R��&'�C@���&"O$�3w� 8S���i��(��=9w"O��g΀.`��� p��:6"ORU0S`�N�(�h0%α=\�$y�"O(��T-vglc䙀 O�Q�c"O�����/%j]#�$<2Bc"O�� �	͖pM���R��B�4&"OhMP��J=�*��@�
�;�"O*0�4+H4��R�b�0K�Q��"O�-�@��3^�Z� %@N�n���"O,Y G�W�1
�K�E]1)�`�"O�1��u�eX�d�{�XH�"O>���c�����%�����"O���
�,8�B�A��ݷnV����"OT�xw�E�3*���k8!Eh�#R"O%S �YN�@�S�ʔ�x6�倳"Od��	��3W�:��Z�[.�b�"O0���F)e�H$R�kԋ ����"Od�p�+!�:�d��� �Q�C"O�x�ԉ		O�i�E*�
X��Q�"OP��p��(2d]P�b	�w�x�e"O�t��%�0d2� ��[�����"O6a�a �-t���
�HE|�Z�"O�q��bՔ 
4f�'rRx�0�"O^벅ҙ6�m;A�*."�8�"O��3c�F�OW �W"O�
A�����c1-��l�����"OV�@��R$���k� �a�"OL��,��*���JD�R����#"O�B����W��9�B�N /�2qI�"Ob�aM�B�hXQ	��>���"O��uჅ*�1;��W�A��%"O�YI5S}��dLQ B�:L[F"O��C�ѹ.u�0
��{�x�K�"O���@cǐ:�Y���g�<"�"Oz��1KN�N=�1qê��]&<��q"O�5"a�C6j`И�&���'.H�"O<)�3�S!1�5��@�06$ ��f"O��zD �u}��k�`β]�"�8""Od���FJO���w/N�a 4az�"O����YT��Xs
�^�.�p�"O:m�d�'c�Y�q��
��"O��ju�˘5��X�b*_�	���"O� ��Ņ�6�*��i�2d��"O ��AȊ*��̠�HPD�sD"O(a�G�4��e)D�O�7��(��"O��M�����d��m��D�e"O�ЂF)N�eBZ)S���;j��W"Ozrf)�Yr�e�@�L[�@�"O��:+N$��u�H������1D�0`�c+Hp��� 9�b郐a1D� ��S=i�9�#d�z���y�g;D�\� �J�1R2@�dMQ2(W�4�3�&D�,ȢKR�}Z�(��Hю:~bP85� D� ��2xnbT�����j�$D��qB+�e��@�^;4z�ڠO!D����L�+tY
�x�F�Z�P�c�>D��	��H46�حI�D? 
l(Ą)D��Rl��,%>��nVz�ҝ0QF(D�|ؔM��~I�F�Ek�m�!H"D�,A���<p����鐅'8�aX&� D�����ҳ"x�!!�&J4֢Y�A=D�����~����,��^@t�%�%D��i�/�A�j4����1�1Pb�$D�0�d��I��ق�cңp���Z�&/D�Awj�0l����
W@���.D�� n�&m����D�;Zr: ;��7D�%�ԭz~��s����}^�͑�*8D��W��8_�0D��Z�
4���1D����J^:�ڜ?�� ��]�<!c�^�'��8���4&󴥫BDBp�<)�F�E?�DѢ
ǭf�rY3��Gh�<)Ua�� [�Z�J�K��1� c�<y�n�:(X�A�cY�e��P���a�<	&&@�TV�}駥��#j �K���_�<�s땓QP^�A-Q��E�AG�<�ceW�:_քR��6��Z�n�j�<�$� q���C��L����jm�<Ip�S,�| ��fʹ�R,�]�<��N�V5Y�Eq���� �E@�<�ѩ_�K��y�Ĺ.ZQ3�{�<���+�*��ͽ�
L��fVu�<�W(M:m_ ]�`�W7tB��j�f�G�<Q2g�*(>L�+g�^�z���p��Y�<!��� 7V=I�፤RP�p�F��X�<A�oӊh+�Xs�JWMP���	EO�<�G��(XG�P�� ���{6jGK�<��ӭL�V�W��7��ˤ�I�<��.��0��İPX�Q4�g��G�<�gk� 86�a$̄0	�,��k�<�E�[N���ܒT6BY���Gc�<�c·�]|�X���4c�zPej�c�<A���:A֒�� �Fr|��$�e�<)B�J�OJ�u(��
����Z�<�ehȞ)�
E���ҍ9ɒ��L�<Q@$�/��L{2��	%���A5��D�<���ͫZ���q�P4�|1)�Ni�<��Fֱ�:}���9c<�p`��c�<��&�$�������2I� +D��_�<��m#se6=�Dc��DA�A�<)v*A�:�R�	6�d��
^@<!�9�2`(K�a�P��� Aڽ�ȓ�x�tB�?"�ơd���ȓ}~u��fP�1,,��"]�T�z����Ժ���݊�c�8^&���sX�@�1�� �ڤ���)�bt��@��T��/��){(�i�ܦ��)��S�? ��P¥���n�#���
��$f"O�D�#i6.��xJlA�E�tT��"Oe��J7a����%��-�����"O�t���כ5��!��̂x��e��"O���E-_;6�F���
ܞ�ҩ	�"O���@��>]9+/S<����"On��B�P$C���jS/T�
����4"O�1����b�U� ��
7� ��"Of�ꅯګ.�x��A␗S�:�"�"O>(���JT�\	��ʜ>v���"Ǒ�����F8�Q�^1�ް�D"O<�A�G۸PW@��� ގt0���"Oΰ�p��n�^�8���~L� b"Otɘ��;c唕9&��v���c"O"0b���;b$F�R�ɂC�-��"O��tBN�N��,����4I�nQ�B"O�!�M�E�pͳR�	�w�`��"Oд�ңOJީ��P?dq01K""Oʡ��
N@��['��,Slf��"O���k�?s��-k��26�U�R"O�  F�
 @l�'ƕ�j��r"O��Bs�ջ|�b�[��յ,���ۂ"O�թ���`�`<iE��6qptk�"O��vGJ2.S~e�N��EWH<2�"O؀C�	P����NK��T"O,Գ��޴ZT��M�V2$I�&"O���&G�"4�p�f��t"O�I�"G�R��-��`J2P�T�t"O�@�ԯN���!�)�5{�RT��"O��rU(S�r�B��S�
=+�if"Ox�0	�#RذSg�R@����"O��pQ�{� ��fD�d���$/D���R��G-d ��IV2�T �W�.D��0�f��(�,�cIJ*%�PT�b�,D����l�	Kn)�ôlB���o+D������\ څ��d˅8Ҝ�ȷ�(D���QD�#�4��g`�h���9'D�Ћ�aHs�DlC�a��"�z�9�C&D�$,�?-}0��gE�)sF�� �#D�`H�no���#��f^T���?D���%*�Q-BHq��K�E�Jx:��"D�<���Ҿ1�L��Ń� 6��,4D�|���LT�H"�aATr�Iu%.D���qZX=�!�g�X���*��-D���o�tKZ�c�c-pq��h D�x��A�7B&a�P(��1��	=D�����^�Paʂ�0��EK��;D����� hPp�7�$N\����%D��K�^�\����#,�B@�$D�,��U���ل�mL���#"D����I2$���"�U-F3֥1��!D�<� �cŲ4Q��W$
X�]1��>D��XsQ�p�� @g��l���A;D��6�AoY�p$$ٵz����g�+D����@C�'�H{��յ]�9q�i4D���F��~]��!����|d90�1D��F@���&-���>I�G+"D�T EBV�9���k��@4e��m��/ D�́ҵ����	ƻN	̡�Ə�U�!�]�v>`������L��ů�3�!�C6�((kpg�l�"y�t���f�!�$٣?"R���I��;�5�� �!�Đ$LtTkN� '�(���!�dT�*�B�Y#T(��ƣ[�o�!�� ,Q�1Á#��q�AQ�M9v@I`"OZ���i�Z���ۤo�<P:���"Oj is�ƕ�F�
H�-�a�"O8�rP�	YxL�a��h��IPE"OD���I&U�:��S�E s��B`"O*l
$��y�xr���n7V"On ؑ-	��ΐ
ԀX$ ��"Oέ��O��Q�"��u��"6�ɳ"O�xc��ɕy�]�vE�?� r "O�䊲�غh���򊒅0B���"O>�U�0ܺ�i �"���u�<�WhͭM$�A�H�<A?FX���Ax�<93B�*z���G!�D���y�<)U�鶱��D:C�����p�<	d�Z�8����HI�6J�Ġ6k�<��\+ �Z۫V�D����.D�\Y�D�_$�a�Y���4�2D��c��ŗ��f� �k3`,D�D�a���o4���R0bu�l+"�*D�'��(:�!x��\vi|@��e%D��	U�ս^����u��
G�h8�'�$D��DB�ళ�/DS�0�{c%D����,J ���!H�*���;��!D�$�T�֋4c����
�1��T�*O����4(���K��Z,Gp�pV"O���$���Ơ@/\e����"OE�#GG�ʤ)[c��@�л"O�L���dY(l�1m�\6v��"O���ܪlȚa��%�5.+x4J�"O( ��+>f������UV}2"O>� ���`����ϛ�&�З"O~TYp�U+5���"��"JϦ�{"O�4��Ú���,�>�t"O:�H��=4ON��fßJ޸��T"O�E1� By�u�Q!2!8�7"O
��A^�n��B#�nP0"O�� ሜW��sr�<��u�"O�,���r%,(�$d	&u�PH"Ot���/��cW �͝�xt¹��"O ��g�!m�<��S�X*+d�D�"O.��"W�^���X�j��9X�S�"O�@�"bF>**@`2p�A�qB�b"Oq:��$���S�S�~RX��r"O�4��D,l��#c�N�4t"OF�BsF��j�0@K�k#�=�v"O� s�Ȱwֹ#��ںzLkG"O��(BCE�b�<9{�nސs�T9@�"O��y�,�:w9�ݳW����2�"Ov����Рsn��@f�/����"O�1�&'�"|XS(ö/>F�"Oh�%/t8p��-��Y(���3"O���CK��	v�����Rs"OhA��X�����K���i�"O���йB�e2�	K�(�Q!"O�8�l�%�B$���yӮ��"O~@C�&[Yl�X�9��ӄ"O�mS��g�P�ҕVB����"OVP�@��8:u�icP%��2�$L��"OL��6)�6��GV�/!���"O 	��l��(�8�juBN�垜�"O�,�aX���l�%��(��d`P"O@-��#��;xj� ��XK��@�"OX�ȒO�Tc�e��N�R4&��y��ä.�NP�$���7KP�/AM�4��S�? xպs,B���lyuC�2w@`��"O�|J���-7kX�U���w�.t{�"O�|��DO�%��Ћ�
��G�=k"O���� �6C�I�NZ�Y�Z�J3"OX���Mͪ'����O:��$�"O yY0$J%*�d�K�ݦ{ٌ��"OvY(7*ߍz�
����
�u���k�"O�t;$ي�0������;v"O��!��h0�\PA,�>N���HT"Oڼ�s�$�昡1�[38�rp�"Oz�B*�,j������u��XP�"O^H�Fሹy~�*@Eљo7 �)�"Or$jF-�J�0d��G�cU"O�]KS�ߎ��3%�O!J�b��"OlR5�%c��~}Рj�"O,<�#�U�/���x��4Nr�DY�"O�d�0��64tN��R�{��c�"O� �'��q/���GU�n��1R�"O����Ń!��-�L�V��J�"O4t����p`d0�	� a�� � "O��6F�RUV� �JˣF�LѸ�"O��1q�D�gh1y�
Xz�� �"O��d"K)'�I(a��&hpU� "O�Ճ�jZ�q^~�1���7Iإ�E"O��a
^�:�b�ZD��2�q�T"Op�����#�y� �M�J�sD"O�[w�E>w��J��@3%�F���"O�q1Ń�d���ǦҹnDNma"Of<A��Z�LQG�/�eb�"O���ʇ�D�LA�OQ��pE�"Od�5�0$^�@04A��1n
\Pw"O�y��Wx2&��EEH^ܕ`"O�1#F���P{��#bBUTP��z"O�e�@�! ��0��7k8:[4"O��Y,P�B�@!#oV�����D"O:�� Gsy�ȃ�mз.��Q�"O�`�th�"N�f	i�L�6!��U�"O(��ئ(|*U��Q���"O��3���Z�ʝjBB�C�d�3�"O�p�O��yBtP�+�%I��a!"O<ěp*^����G7.���f"O޼@�"Y�xyx��ŁӨ=��"Od�ihg���cF2Ȭ���"O��s��E03�}�4�T [��As�"O�)���+B��耳J�w� �)�"O�-ӐG*aj �dD� c{jq!�"O�Ŋ��ڝ+�dR�S,7��r""O(IY�)�2�6xI����"O8X5��u�򰲠��8j||��"Op����ӿm$�� ��8k�n�)U"O^��睄0P�x�@��d�f ؕ"O�T��a�q�L9;�[�n�Pb"O�`	��X�B<c����^$Y"O �V��7Zs�=+S�L$���C"OF�1Uc[p�R%iQC�2f��)Q�"O.�j썪}=���ʝ?+�+�"O¹#�n�#3�0YzЂ��C"4��T"Oȉ�F�^��QfAO�,��@�"OnY���C./',q��&�0j�""O�ݪT�P��$,������"O�\��'I�`�Dҋ+tt��"O�xx#�C, &z3U"уAo8��C"OV$�r@L5�"�jW�� T[xӐ"O�����)g$@"��ΧiS����"O� }kR�K�y&^5�GA��X�"O�Ȳn�b�*T,G2K����7"O��I�X�����^�:�Li9g"O`��B͈+5���@1�!~�-+�"O2�	�=[-�S�ց#q�]b#"O��Z -g4������cl4�g"Oܭ���
`k�	u���W5`�b�"O��ypJ�1E��S��H8p!��
�"OƜp��|f0���%�>�Ji�"O�]C�T-~"�|�2��x bl1v"Od�a�@7p�c��P��"Oz�
��>=�Q�D�4^Ҳd�5"O�����W�h���H#$H�F�VAP�"Oz@&�7B̲���ߐR���f"O�e���? 馩�W��tQG"O6�[�ü ��!�gcǅ&�z�&"Ob��ua��i�t�q��)D�*i�$"O*Z�	�n���K"gmF��"O\��b��Sa�`��]�rWF�pa"O��ғ��#�vT!פ�@8�=�"Oz����G�NT�D��$98,���"O�$�W��>LR�]�7D/	:�a"OA)0�W<�RI*�D��� @BV"O��q%�����Ѳ�&?���
G"O����eE	�&�
��-K�����"Or��4���{H���bZ�}
�"O�,Ya�"J�<m��nA�|JV11"O����.��]J�`�2��s�6\�B"O�@d�D9	L�)�K��Gw�ɲD"OR�(s��8rlP��c��f��9�"O�<��&�7��tH��2�l���"O���MK6_��T�m���tI�"Ob�����|����l��d�f"O������;Uj��K��B�Iv�s`"O0�;2�9D�� ʚ�|�~�$"O �ۧԆQ�89���M�g����"O$]����"M*���2mZ�{���v"O���ShR���p�L��6Μ]��"Or�U��5y��PkW:���"O��P{��S������"O�����B��|)�
�5� л3"O�I�&!H4`�0��2�r���1�"O��8�*�#���K�T�y��`�"O�`h�g�/J� x�N4���"O8T1ȓ�^����1X���"O��dO?���`�T�|���S�"O���p�A�#@hb��O�jdƌ)"O`��N���a#�!u�yK"O��µOZ���
?d���"O���iN:���F暁'Zz!y�"O*$��mA�����=!����"O,:�.�#�ڑ8���5
��`F"O2m�'�Q��yP�,W%����"O�T�]�ej�x��k�5��͑R"OT�ca�ZH�։b�� ^�!#"O�S�פke�q�i��{����"O<Y � ��n$�&�Ee$hqa"Oh���e+��pu^�%[� Z&"O�t���ăD-*�s��X�r?��B�"Oh��D��%i�j��Q��t"F���"O��Q(��Jn`Y���e l��"O&��5ꄄSذ��m�c��"O"��#�Yt(iӳ.�<q��-��+9D�́�N�,.h)�������R�3D�� ��TI\������O�=d��P�"O�m�g	+H�����)6��qё"O�2�*�*m`2%S��B�~��}�r"Oܰ�p��o\����FF�JIJ�"O�]0u쑒Fl�%J�@־a�`HDxR�'蚸h�(I�5�~��)��#lt0@D!��*�b�˳�}��?Q�@�(})X���8(d�(f�^Q'0�?N]�4�O�&�Вd`�Z��#=�i���Ѻ�!ܕ!(���3�@-w��$HŤ蹥�+�J�0ǆ�~ؑ���F
�O���ͦ���L��*�;�~��@
n���X��� U���d5�)Z�}bNN#<����oݷ6����Y��p>�4�i��6nӪ��U���}�A���B4ʁ1��Ot�a0 ������� �Ok����'��i��4� ��Dj򮁃�j �d :s� ���*D���8X�L˛Nr�<��OR��?e�1&�8yHV��Y�"!�E��/"��n�76���+7����B=�t�Ӏt;p���\�r�hc>�X�s� ¥��$�zsǕ�s�7-�@��u���mZ��pD�ܴ;( �C�E�D�s�/̨Y�L���?�/ON���&OM��I>�N��f)Ɇ9��8o�ԟD&�<��1��p�P��7!
��˃� Ah<ҥ��uyR�ۛk7�1,O�k"�ua�:rv,�' �*���P��M A�w���+��(^�"<�t�N��d:b���o����L^�Q@��&���U��
F���O�#<I�'^�&k�٠)�B�&�A #��d2���2Ob�\P����I����'ʊ!�O	���	��Fۗzx�����Vh�@3*9w>��N�=8��S�JbӚllO��4�	�<1�#K)<TТ7 �'r�`uزO(1�x��v�-�?I���?���~/�ъ���?���1��	����YoHmJ�ן1S>���CҸa�,:g�H�D�Yh@��8S�#?2�\"+*�k�V�i+��L��i�A�ٱlV�Ha&֮$g@	��͗�-�j�<��V���n�Zz$��1�)[�[J�x�a�i�RV� �IIy"�	%�2E{u	6;P �i������hO�:TYd�G�a;� PS�/$Ξ�yq��՟��ߴ^h���'b.I	d�7M�O@�$�O�EP�7G��@�weVp�p���2[T%�td�O��D�Ot#��YYtp��+EAJ��0�M����ə-C��bD��n7nP��K��HOl���Ď���0c`.*_(q���@N�����L&0�VD�A�G�S�5���s��r��O���N�ܦ��ĝ^��M�"�Z�&�4хMH��?����i�>��+�`F\���CV�Ns��!�J8����4TE�ֻi]c��%���F�>���'�$ ���y�N��OX˧:~ҥ����?�4v	�UɦHs^b(xFi�n�Aa�a��U�(�G�W�}��LpB�������2֘.] 8�����f�쪰�'�z6�I&޸�h�nXo5�E�GgP�o���q���
<�1�k\$!�̙�ƌۿD�$�RB�ǧ$1�6D���?���i�6��O6����u�C>Z�R0&���G�RQs���p��{X���
��tXp���p�D1&�nƛ6�u�֓Or�'R���'f��y%,�k�b֭)R�p U�|��'�N`X� ��   Z   Ĵ���	��Z�RvI�+�� 3��H��R�
O�ظ2�>��j& ��ش�?A��[$���(�E�r�c2��&��s�}m���?	CY���'��6O.���.n_8d1�I�TT��k���A�p�ش)iqO�a��d��Móg�$4�H5Ѷ���=�
��F@yB�@A���#^��$��yލve��=�(�*�E�a2����Ȍ��X���=3��<�A�B=Z�'�+G��� (���p��n3ll{��lV��
��ۼ
���.	X�|�T���I&c��8�DʣWP0{Ŋ�- �� u'�i���K1/Cc�	3i|��c֒|�g� W|�Z\E�zͫ����	$�ɠ<]�Dd�I�(@���Q#����I����q���DJ��O�I�OZ�q`T>��5�B;02R5���>�W�5��➔
C��#/�u2L�?J!&���z�u�����"�O�x�#�] E5N� *N="�`��o\�a5�O����$A7��dD�)KNiұ�%߸���T��	=[��������`dH�i�Ĭ�G�Ëm��Ȑ��dĝ�OH�@��E���l�/��=ha@ĘL,�T�<�f�;�x��O �(��C�rR&�!���#�^6)��((���8�'v���>����sM-MT�逬��\[l�D�Py�0�pi���i���������� ��%�"?�$T�tCJ�s%�$ w��<q�M ���$�@F��#��O�<�'�Q����34Í6~-��H�_�x��?o ���p�_]H��O�#�(�ñ�3D��u�   �R]3dcct���*��C����n�>����?	���d�9T8�(�O�rcմ?�Ei$�[��x�fZ_|"7M�O�˓�?����?�4���<qK������&��R�"|�ūgJk����O�˓gBܐ�\?1��������f�B�Q���'u���//l�aӮO��O|�$[;��|�������:��=sdl<`��M����M�*Otq�5�U�e�	ן8���?U�O�.�J�ā��j^�T�Uc�W���V�'���yR�'�"�'�q���`)��Q���)�>�jtyַii���Jj�|���O��$런D�'�	K�`<�En�ikŚ��:��@8�4N/������O)bO�"�����7{v]���N�6��O��D�O"\A&��U}U���Ii?9@�Є=S�dh#ɩP{�-9 EB�	��Uy�����yʟ���OD��ЄR�����# �C%�:���nڟ�땠����<9����$�Ok�^�]���zv+&At<�r�S�
��I���I֟P�I����	ߟ`�'��AY$c�)v���{f$�a,��{`OSE��듦���O���?i��?��JFLDXIVǆU�z��v�Dd����?A���?����?i.OaS��|2/P9*�E�G�,81ڌ�Ѕ���%�'�W� ���H�ɤ2���I�r-��g�G�l��tcH�L���
�4�?	���?�����I7P�O�B�]�5b�9æ �*�^a ��P8]:���'��I�����\y`nh���M�7nT��)x�+o�b�//�|6��O��$�<Y���%��O���O�rIi��7[u�l�䨑V8���G�%���Or�DU2fp���.���?9땈��X��|bE� ��0���d�˓��`A�ifL��?	�'jg�	 ��)i�	]�
y)�B	�\_�7�O��d��h�P��+�D;�S�&g2�+�P�oSԨ9E��k��7M�)I��nZ����	���ē�?�� ���'b� ��hRE�c�f����i,,|��'��'��.�$�$�� ���؝#z2���gڪ�F5lZ���	������'"��O�,jƛn1�V�C���[2�i��'�ސ`�d>���O���O��q��˃F��X�C��#�$�瀍��a�	��t(*H<����?�L>��:�������["�(Oʘ�'u���'�ҟD��ПH�'�����x",r���~H !uʂ�8�c���m��ߟ�ɀq*��E����6�	pDd������'RR�':T�0�cD��d�ܐ~4@	#�ÒPz�A�@l������OT�0���OV��ªmmX��H�4��3M�	z�\z��Z�B=�'$�'-Z����X:�ħ"´A���ɄG�����ۻVp,r��i��|��'�2�66�>ɗ��g�d!bcշ3���k�gYӦM�	矤�'��K!��'�?i��>D�8�ykJ� L�
u���C�xr�'��$۫�yr�|�֟y��GH4�=�b
�n����is��_(,D�ߴ`��Sڟ��S���d�%H��Dp�O�0�����3���'����O��>� �i�/s��*��S7|D1��m��,��Yݦ��Iߟl�	�?��K<ͧV�0�:�O�bV�����ʝb1�I�0S�X��Aya&ҧ�?�+��aj��ߝG�\��$�Ұ�&�'h��'>@���'�V>}�IO?A@D� 1�g�P&wUR!@���{���9H|���?1��uN�C�(°�����V�Z&v�3�i���pO��'�B�>�7� 9�Pw�٪R��!P���m}�
���'���'���'tL9gN|!����X�R!23cZ'M/8){�U����͟8�	S��͟<��3�(�w)W�ļ��f�J�N_�n�(��?����?�-O���EM�|2�e� 4sL�'�T���
h}"�';��|2�':rE�������\�@�S�_�	;��^���	⟴��ϟh�'ВX�5�+�	S���c�K�y�̓v���9�n�8%��I蟠a��'�I�od�0�qGڒT��aA蒄$$7��O����<RN�7FE�O���Ot�|���hfT����	�ɘ#,�d�On�$��A���'%|P���C�ThC��I	Hq��n�Oyb�ըl�L6��m���'.�D�$?S������.������������� ��?�S�"���Ԇ�W6�'��?Ln�x��X�4�?����?��'~��'�P�yD�����6��+��- 7�Q�K�"|�J,��F�)A�ʢ��.L�	��i�2�'Z.ӱa��O��$�Od�	�mlm���	/U	Z�`Dm�*b�H���%�Iҟ��ϟ��0�$U�2 ��?���H�"��0�'-P ��/�	ӟt%��0Į�AthK)�~�h�YN&��.��<!��?����~��ʷ�0s��0�u#�;bP�����a����$�	e��� �	<7ԥ"��O��ΑjB �
pL,t��	9�ڟ��䟠�'2.�P�z>����%���el��:�H��>���?qM>��?YR��]}� ։J��Ȅ���s��Ϻ���O��$�O���&�����D�R(2�D�r��1%6�!��7�z7m�ON�O6�D�ORl����+ n\S@�#E���G�S ��V�'5����,#t͕��,�I������?Ap�F�ޔ��b�>d���5��3�ē�?�+O����i�M�����ki�P#�(�!��­NC��^�ċ��2�M5T?��I�?�H�O�������t�R撹�6e�C�i0��'����F�%�u����9t�(�ٴ)w�ـ��i���'��O�O�D	�D�ZA���1����i�p�P�o�;*��#<E���'� ����'h��a�Y!��dpP+`�8�d�OX��!N��#�)�On�	sN\J7̒_�b���q�J-ˎ�d�V�����	ڟ�9�	љw����\H�91��M3��^n����O`�Ok̕�$B����&<��b�;���������Iky ��A�6R�0��)؜l"�Cp�=�$�O���>��O��	�k��@�����jmI���Q
c�H�I˟���^yrkM�Q��7u qS���:p�� k҉N�hB6��?���䓍?����r�':�²o� }���K��+l�s�O|���OZ�d�<��H��	*�O������|�8��Ω4NdX����� ���O�$�� �O��@�R4L.���#�8$� $�i4��'0�'I ���'�R�'#��O�Y�Q��3	����%&Q'DRA>��OL�+`�GxZw���j�B������/K��|�ڴ���Ym�Tn֟��Iٟx�S.���ư�ŀG�H����ϼ`��M�T�x��'�ў �OF�I�dZ�x����0<�	c��i�Z�ô�'>��'/�O��I^��ɬ:k����"B-��c���y*�'I��Ex���'X⹢�A�:�6���㈾��@��mӦ���Or�$�E>��D*�	�O��I5q���`�@�o$#��]�>�.���dZ�SΟ8��ܟ|j�L����ᰖLE S�ʉ����M�� ���S�x��'!��|Z� `9(��R�$Z���%��-�E^�!'6�	����ٟ,�'����1D]DԢтd���>5y�O���Od�D�OP�Of�d�O���0��Z,��w,؟8 ��Ѩ0A1O����O����O���G���$��sݒ	q�Hu|(6�ڳJ��PnZӟ�	؟'��IXy�h�Mc�W�w�朩�냼��!Äh�[}��'$B�'z��(P%r݋�����W8�bY�����K�1PV�ymZ̟T�IS��?�{�Bѝc��%c̈^�݋J��M[��?��?�4b������O�������c/m?���CA��`Sfu�@@a����Ȗ'��� ���&�C0J��C&�������xR�C
R�52
�PF�=����x����c����D��=A�e���ŌI4ҁ˖E3=��%���5,x� t��fE�A3#]�2a��AZk�!�G9)Έ�HR�;fqXqp�.4;�NL
@hD�L	茂U }�Z�Ұiơ
�~D+��-R)��&+"��J�jA�X1�lB�y22��w���-���\�t�~�K�8_�x`�fy��R��h�	�|�I��u��'��,^Up���/R���&e�Za����-"D#�V I7�����hOz��pk�a��� K��@�@��qo��@`ը̀<�*A%�X0+��퉃l�Ɯ��sYy�aN�by��I�<�4���OȢ=9+OVԫtkܭ\���ӄ,�kl��H�"O�lr�
X�"2���J*)�")�� Y���)�<ٕ&@+�F�v���*b�+gr𰣅
U}q"�'�"�'����'��:�P�F"m8y!�<9���#ٰa�s�Yw}�Q�p�=<O8Q�@�gN����T�̬���Y�#���Х_�]�
�F) <O����'�"�X��4�J�i�+NP�ў@F2�H�dz��n`{N�GU1�y�
' �5(�)X�+>��n͝�y�>�(O`hr�[˦e��̟|�O�p�Ԥ��Z�:U�qnΔk�:���!^�JA��'�b.K�x(]��T>��
k'^�+�"�Z�n1���*�)kdh:6�SP�R��״]$�fV!5\�<�AÅȟ�������I`�D�̺n����w�S,y&:D���E����s�d���l��u ��ݦa��4� � �O��$����»%+f|��m\7&M�@x%,`�`��'�M���?	-���!1�O��$�O��(W���V%��)��,'��`�NB��V���2��E��\ןʧ��?ɓn	�c5�U�5���A{n���F�<�T,�U�T�n5��0�a'F���'��Ayg��@��= �%��rY�53�)��w���'Y��H"|�I<P2��"i
�~�BE˂���c������X����L��}�#N[�?$<uCQ	����"<���)�D`Ҍ~<-Ig+F��u���7�?!�i2�4�q�O��?9���?����OT���7���ID�{.�p�/G�p;���v@�}�k+=��i1֪G;���ͯ�~��Ƭ��>!2��C92�����(�4T���ׇ�?	����?)���?�gy�T>�Ɉ+�wD�~�Z�q�م	.rC�ɲ
�����,[�nD�)��W"�P���?Ք'H�+��bӨ��6(�(Ҏ�V(;���O����O�d7hY����O��*��+/�"�ban��H�P�	��u~]��1!�F����[�_�������i�Ȭ"qʍ� �`�$E�E�-(�
,�BmX�ї:L�0#��I I�����O��!	�pS\R�
2x�2�	>�d�O��i*�)S-��Q`v��EV�CA�ՊA2!�D�4%�rQ�i͘5�9�����2 ��o}R�)�Ӕ+X�0Z���L2^C�����VB䉨	)� :���={�:�R�0�tB䉓k��A�G���t�rH�/[
`�C��*}����p��+24J��,ZLF�C�I�9�P�)@�DH���b�E�`.�B䉭AhbE�C��8*W��[J�B�I:0J�p&I��&�M0����BxB�I:o�-�%�8Z7��z���5_�\B��9U��|��A���K��^�n�C�	���	p��R`�P�ݍ=5�B�I��(����ر��%��f��B�	%\�ъB��(�d��d̝�k��B��"�e(�W[�u�3 �BB�Ɇ0��٫�@S�I����b�9�C�x�̠A0-�TA��ʫV~B�I${����6�ۦ
��9���Ǳ!RLB�I��]�с���}�v.�+��B�)� $�� ��j�t��u��,XH@��"OXM	$cױ1'�C�������"O��S1��r�V���e�0P����w"O�k��!�z\�bE�+�f�Q&"OD�sSB�3)����Pj�b��L�6"OF��v�*&;��$J^+Ӷɫ�"O����PQW��[��V
@�J�ٲ"O8�t �z�p���%!�\��"OF���S�a���w*�C�T�U"O*=�Є�.ml"D�2i� )����"O�L(bBmf�ZTƈx�z�)�"O֭c�A(w�����$7�`A��"O\\8�"ݼk�*�0��E�ԥ��"OQ�B�0{��(�U��W��s�"O�찖�Y=��jrm�&fG��;3"O� �D�G p�Ԓ���{bDx��"Oҙ��!Z0=@$x:��@�p�$@i�"OȨ�+�N�k3�=b,�b"Oι���Ӝ�� ��A�h6�@�"O�X�Х��A�,��OA�xNr��'"O4q9v/��BY#��D�pe:�"Ot�F�1�佢 ��=Z�4�b1"O i`�&�,!�Y�tm 7J|Au"O�)�ԡ������5��}���ps"O$A���1b}2�l��c��	r�"OZ%�D�]�t���C&�=7�i��"O��N�C�b���zٰ=J�"OH9c"]���q��-jШ�:�"O6(a�g�5)�xX�E���.�q�"O�3�b�qn� �0�E�4��T3u"OH���+ۗa��T�%���4M��"O����߷:Q��o�+��X8�"OFY�T%
8�xmO�}�f��"Oj�!ԠPFv`Y��(dq��Q"Oڑ��*W�0s��f���]�����"Oذ�'
��F�0����/(�Q�"OnL��k¨Q���ʲh�4q
�m@�"Oĳ�ş�:���نʁ),�:��"O0�� �IFFu��ʇ�y��BA"O�ĉ���73>��p�JܸJ�P�p"O�Lڣ�1��-r�
 Q{|!��"O��hQ^:c�BH�B	Ƈ���{5"Ol9#��S�+�j�V�X�~�l̹�"O�6͍6+c.Ԛ��N�9�d��2"O��3��HT ��� X�l5�R"OpAB��T�qb�%�Fe�*s���8"OB�qa�!=��հa��+��ģ%"Ol��Ϙ�+��X�5C8M���P�"OLD�4d]�2E�������t�z""OZE�F#��W�
k��E��"O�ّ�TK:�$��ɡk�j-)E"O�|A�BQ+S�𠸰hN���`C"OFx��ʎ�U���Ʀײ	e��C0"Of\S�O��h*�1)�f�8Gd��	d"O^i�GC�'���#��]!mIm�"OA�$��4I�\xǥ�'�BP�"O��3���<]SV��g/S�ƨ9 �'k�<@��'�q:�D/	RHp�1�Û6���'(ji����S{~���οK!�u�v�K81e�">	�Oҽ�h��!hR�&��-
��;p�\�J֕>�1�=A�CڂZB�j^�\cPf�b/\��%eQe��1���F�&1)���]���Eӟ�S�&�ͬ1N��1ӳ��&���f�D"'Rp�ȓ�ơ�6oP��� B�z>:�A�<��P�JA������	��B��� ��,Z��y�;x�upu��0.4��GG��4E��ŵC��n��}�*T�#�4\;�� �� �.	��훂 N�(d8 ��h: m2��DȜi��ŊF� zv�	?I���>I�Ҏ
<����*�r8sg��C?�T�=d��Q��˙K̜%	be_<kŞ�Bdl�O�����Q� vKC�ҏO�<��a(D� ��}�L��t$.�����z&�����U7t')���=3�	�a��9�uBu�2z������:�����U?�p�9D��.[4H�8"�,ϰf�P�` $d��}�h$U�D��HK ZNl���4�Q
����P��^���XpB�� ��y�M[�`�ܠ�,9���J0t�Ɏ>�b�#c �y:�%j4�|X#=��bW?;�̐�5�]h�4�Mjl���O�&Q�F�bdՎ6j�Q��$$le	P�j��>��0�DJ�V�'!N=GƝ�р"G Z�\ڨ!�0��x[2��tȡ�"��< Aʅ�u�*Ȅ�:�L�5RIф@§{�|��c��"�U[�)�4��~��Ȯ}Fe�`Đ\<��Cѫ�<y���mL�ZA���W�|1�cO�Y��'T=ɑ�wT��"I:n\����E�b�	�<���z��7Qվ@��lQ�63�cg��5����'�*���#+K��D��*ߠaj��R�y�R����ϺY���-&����XJB��p&@�*�����$>��iDAX�x���O꟤JQ�)r�%A#B
��˶�21Y6UH���d�H�N�4P�"��'2p�!ԇN!E"�D���^0C8`9�'��P *]�(�T7��C�p�#���K�[W��1jE�N6����L\�4X�d�qM?s)FU��k^)zF�$	�;��I\���e�{��S����[:���@	Xض��牁_*(�@�A|P���k�3\���CS�����-��I�a{b�?�$qąV�pO��Z��ĈA�m���X��hOBP��+�c���q�b�( ��"%75�h�&C�,�(PG��0#����&4�-Wd	��KC e��n�2�ޅ���I{�b�2{�@��8r�dd���##&��=kH �cgDV&Np�Hy�j�;7@��2N�	2�<�(�'[�9�J�!;��7-��g]d� i�g\R�1`O�B䑟��r�\D�:u�QA����$��jG��B@�B�^�d�:)ܢ
�����|�8�1 ��5$D1b��֞z�\l�Ӏ3lO������Ip
\�ѹ`*R,>g�
c�ע+��|�U�`j
��z,��c��쁘��Ӿ
j�iVD�/y�h����O>��{m5�6�J�:Ҥӧ��Z�~Z���jڿO��c�O� ~,N|k�C�'r���(���O�R<�a�G� >�N}i�K�2R�	� N���ѺJ�n-�$���B��L���bHG���B�	ЩY� 5XS�͏��es(Oޭ0ElO7c�Ԙ㠣E=�&L�B�'D�u1�D�N�Z�QmҴlDެ2�y�'LΌr���'Kx͒b��f�45PEc�8*X�@��.i6�Mb�EC#�FL�'�2O`d�6��f&�x���� Zt��CV/S��%����+[��)�b����'^�d��(iT*9`a֮�D���l����ē�J��.�^�37C\�.Q�L�Tm3�Ru���D7;�V%��M���"�fPHy"&S�h�&@�����):\�v*��F�Z7b��B�r$��t�xYG�c݊�%�@ ��,�a���A<��f�Y�c�n���)�>�T���#�ryr��8s@���túXbR�ȑ��']��Ң�R�����' ���PM��#OA p5J7ME�%.���P��z��J��W�8���_6���=3p�uA��7�>`�Ah�O��1�+|O�����_}��1/+ �s�hl�b���B��d �
џ1� ���xBZ��n���T*��#��cb�?9����N&� (U�Y�'�K2�X^�h������'���u�LΠ"�F���ہ\m\��J������c	�<Z�y���:\�x�g�!t�H����q��fa|��l��k�f�R��#�x�<Q��+c��y2�G.1Jfȸ�f�H̓D����̏�`d�� +;�u�O�9Z@�A_?I@���AO�y#��� �����N�<�	QҚ<!Dl�zw����n�J�$��3Dv��s/ɼ��<q�L**Bd�	��5K"lr�cm?&k_�w��Xؔi�Yx8B" u�'\Ɉ�Â;Q�@ɪ�f\"z�OL���o˰?�������1�D�i���hu�-�Ǡ
�~0JXX�D�[�R��4S���&(��ԛ�쎚$�P�#��/M��h�ŝ>��O�$�
�'6"\
Fk`�H�@͠k-P��teC�+2��=����5Y�X0X�T"D�\i�JEE�+��Ez#m}.8�S�A4W42O�|0���A?��Y�����y5EqA+�9k��a�D�U羍�#�è^�ҝ�C?6���Rq�˘x�8��1"�Ix�\�t'5�Υ+�o��x�yBn��(P�.\�y �����32c.l��� g�ۋ{ǚ;�z���G�6$"�BՋA��yr�$~��͒� �2&��m�C�(>�N`����eF�_��M���ޝW���g�Dݼk�O��pH��h�瀸X�=2co�\������=	��`���C�6�Xu�>'����:D��x0a��Q߉'<�h�D��i}bp�d$ʲM\ps$->gF�E}R'5MN��D�2C�"�3�d\�|BU�^9#�1rVg=��)�k�`}B���z�(��	Ĥ�x2MÛ7�<�k �3X���ɑmΜ�ga^9Q���� fډO��9�Q��?��#O 8w���ǄC�vކ8��'D����
�I�(��7���F�r�G	/����4�c���bC�ʦe��ʚK��O2��;R�^�H�%T/Zx��q�����+�i��:S
��������&�HO?i� �� 
��I�j=�2�ҵP��1�"OtH1TBV�� ��/Z%1�`"O�P���Q��X��'5W���[�"O��0��Y=�8�Q��![��m�d"O��� �<� 5���M�h�D��"OJt(fҽ2�нcD��(h"OTx b<ڵa�!�LT�"O�(# �r2��d
[.G9~�0"O��S�\ki�7Iu!����"OBDx$�N/�6�3��I+@�X�%"O4���CK���j'OM�3��):�"O [���..���cN�=�jq��"O���&ʪf �ś% �~���"ODM�S�
�4j
hc&�>C�h�"O���&�,D���fͮQ��+"O���$�$3� ��FR�Qꆔ�"O�PrJS�lpΰH c$՚h�"OQ���RO�&qw���{��� 3"O�9����1R�j�qV럠|���"O��⤂�h����G�݄!l"I�q"O<(�TB�P�܀�I�8s��1f"Orx�@j,L#^�S(�h��A"O�����,�~��g1b� �"O(l9�`�(A�	
��#[^�*�"O,�	�Kܔ~MH q%�5m�RF"O��E��r"�����Qj�U��"O
��0{>�����C�"M��"OdX��ȝA�$���F>�mIE"ON�(p�N��U+�'��Q&b�("O��(�hI�Ԯ�ca���6 L8'"O*@���~R��ED"f�R	1�"O� @��] ���0%�Q��"O�ʲj^�<<�#J����k@"O��k�A\�Q������G�:T(�"O�����6�*�
9�8ز1"OFu�#��'o� ��S`\�Y�!Zg"O���D���su�]?���H�2\��#�xF�tkn�"��!�ȓ3T*Lc�'��4cDC�<0<�=��%��`㒉� �	#���6j^�4��/7.��#O4��-b�E44�|�ȓ7�x9#��7?�����T�!�<��ȓVA������;?���+��\�D؇ȓlB��G�:2d�C�"�F���ȓ]��9;cH�� �9�qh�Ai2@��`�e[F9J��%�S�!�a�ȓ+�X���h	 ����gg��A��Ňȓcߞ�(�(H�~������
-U�0��B�p�C��� {���s
�����tǢ��C�H���ĳg�Q Ee�ȓ0n�Ը�l�~�*�cf�;#EȆȓqö����ߖ I`�֋��n#�Ć�l��EB%��9 #(T	w ߣT�����`:d��6�,q�,R�֎�ȓ�&Xҡ��R*U��R�BT�y����!3&��n��J�
~�L��ȓ p5QуK�O�D\�

��4��<�:< ���<^9��{d���S���ȓ-&�����
�SUMMS0~��4���
E�A4G�Fp{A��)l8i���.r�OR�!Tl��3@B��<�ȓV�,���]�a�ЬP��EJф�g�����B	�6�N]��-H)��~�,�`DD�A,�$�����d��S�? ��� �m'jA����<7�$���"O�D:B���dS�V�y�.��"O�z�M>C��<
reO�|���	"O��y ���YN������3��9��"Oɸ��؃w����LX�8b�Ӑ"O��ؤ��:z ���ȃ2�����"O*ey%d�Q[��"тy/ ��6"O���+�x����A��D��"O,�c����%�P�ϞQ,��0"OlY���l
�]ۗML�ThAK�"O�!�F��4i�eH�Q��`�"O�SP/��\L�fL٢�z)�"O�չ3�^�ޡ����T�ƙ�g"O"ق��_45� ���\(y��1p"O܄��$��u0b�A�h�3j�,�f"Of%t.P?[�%�%GN�88(0"O�Y*p�ƞo��fE�	�C"O�t�t�ۉVÂā6挽 �hh)c"OB"SE�o�d����.8�D@Rg"Ot�H�IB�h��8IN�(��"O�a+��G�"d�L���S:\J����"O�U�BE�1;�ܠ���	S�����"Oj�ZB�B�J���"#/B��jqZ�"O DЄ$���y�NF��|��"O�\H��ʋz#&�#.^U}F�0"Ob�yW@�02F�#��,pS`QZ�"O��X�l��x�d���L��|Qh�9�"O�isbhU�1��"�Q_|c"O�p`��RG����J�L\E�G"O�U����<�z���8 ��E"O4� �'B���pc�BaIw"O�H1w+��O
`���I���s"O4���葵8��r��:R�\��"O�ͱ�¦T�f�	��U=��ur�"O� ��*�8\7��0��9��@�`"Ov����=�<���I����4"Oؤ:%^�V����6NV�l��	��"O���g/F��`Cu�7;P �a�"O�,+c�Bo0bu:��;E�H0"O�A���s�n,��ݭg�򙘢"O�@J�딋>'��kg
T45~=�s"O6�gdA<j���i�hiY�"O��:����3�<��r	��4�n���"O
uK�c�
p)$sC&H�8z��v"OvЃ���dj��H��jZv�F"O�L胊�,�� w�H^$�"O|}���At����q�ڱ��bE�yB́�k]Fk�l�(<����i��ȓ#@&Y��v�Nؑ7�L�h�ڠ�ȓX����(D/w}�PZ�e��(�lq��O�z4��h^"tz�<�ƥ�^��|��LW���p@o����o��zv�$�ȓg��9J'sҘh�n��d�>��v�.Ԡ�.^�i���f�CD�t�ȓA����2��t�f9���A� 
9�ȓTpt$�U��1m��Wl��t���iy��c`E�YG�Y�i^�k_����8
��hR�0��fB�%�(��)�DJ�OO�C�,��/��,fr|�ȓj$]��ߒP)�L�XC��F��:\�흱=�z�H4bؙ!hC�	�y�#��K;>ZL���Vv�C�*R>���'̯I�<�1sk֢�\C�I_n�I�o �BT�7�ћbZC�)� ���Q.1�N`[���y��"O�=PA�{�t�i$&��8
��"O�5A�F�6B�ݲe惹b�p��"O�*%�x�b�0`��V��y2*�#{Dp ��1�:��ğ��yb�P8������i�)�(M+�yb*ٔj+,�85@�
s4(1�e �yB����й�d��Yu ��y��{��%���ʼkV�9�C�(D���/ԛ���F&�~��4��l0D��㪗��@��$� ����
e�/D�<�@@�'�̩҆�>A�d���,D���+��2L΂l4l94�&D��@V`M6n28��M�/w�A��#D��8�&H7t�
��݄ao̵���#D���㚬N@a)�?\:��d�'D��zw��=�{�A����� D��f�ȣq| p�����Ok���V=D��!g��,z t0&O����s@�9D�(r�o g4dl����X��4D���!��a����Vq�Q�c�0D��Rr �t��h"g/h�ĬB�/D��:�B�v�(�?p�*�"D��B0�4�t�u�m[v�k��5LOL㟼�0�Ʒ�8�w��-R:hs��4D��s�S�0��` }���# D�D	4o�1(^�}�"c�j��)P��>D�p���^<s�f,�)a�;�IK���r�4~���B� �L�2�aD�;D��Ѝəl�p�۵��B���"&$D�@����~wX:�D�R�x��?D��#��Ʉ3k�Uӄ��?:�V̻�e?D���+Һ����j.O� ��Qn��ą�ɭx�PWd�?	�:�� BLB�ɊI:Pd;a�?N�BX� �]�}B䉇O2��fH��:�����ŢQs֣?	��Ʉ�7[X��rN�i<��qq`C0w�!�,�Z&BPΰ�4I@�k$!�d��%4b}sg�2n�4K��,?�џ(E��).J%��QT�Z�z�b��cض�y�c�4r%��/�r*��9���yb"�
���i' R
iHx]H�Dȇ�y�+�.v�r���e_w�! �*Y4�yFǆ���:��ޓ�"���
M*�yB�A�B��Et���B}��Cq�Է�y�)_4��<[��D���I �
�y����d����$̟�P)$$��ƈ��yB'�+_��Tʅ)�6=�q�Ѧ��y"IN�v��sn�-V�qq�ܾ�y2EáY�t5�%J\2 4�i�_��y⩀�nNh����5��KS�T�y��� \`�J
ťv���G��y��M��6�Qs#�\v�[����y�Ɵ�'#bh���#Z��2��Σ�y���>�f�аC�"Yvx(��c��yrb<[-<<Q�Ƨ��i��dR&�y��k��� ��W�H  �Γ�y��_;.����p�_�A@X���ƌ,�y�O�p h�ik��0�s-K��yr&_�+�ŀ�`���cI��yrNЏ9@"��r#«\þ
����y⠛8[:���J�(Pټ��BH(�y�#ƾ	���Q!�� ���Ң���y%�d��!a�G+^v�zK
��y
� ��H �P?uÖc1D���5"O���5-պ1��*#X�q3��Y�"O�<c%@�j�@Ly���9��"O~�Af)�1�<Bȼ.hx�B"O��Z#ʓH���P��4�x�"O:�x��Y���XC�/l����"O�J�K��������t�b�x�"O�e�����#W�l�� \ {�����"O� ���<� �s����8���`�"OR������P���խs�����"Op���Ǆ9��Qbo�!��T��"Oj�B�� =f+�c��H%N�x���"O���re��#v@Y���&W���t"O*��q���,�8�n,D���ɡ"OT�u�>jP�EB���95�����"O�x�6(A�d��QA�a�8,��"O�"'k����� ��3��q�"O�ݹF�рT���S	+G���J!"OB�1��r��	:�H�u�R<�0"OD���m�3����r�H���"OTP�Q���9����(��E"O"�0���6�z@V�- b�=C�"O)au��i:(P�dI*�H:p"O�ӣ�ӲA�^谄�[���["O�`[W�V�C���w�
f�L�G"OL��� @�P�$�*RD��,FZ"O�QjvHB�7@bl�7#D�k@]��"O��T�H,/z${�AFs-�A�s"O����-Z�X�p�D
&r��T"O�Y����'=\����Ȗ}D ��"O�`���� ���I�"R�YI	�'ˤ̃@ IY�D��"��}
�'�W�ám�����_�Tp��'�r��%A��'Ӛ��,MM��z	�'��d�T���z�"g�(>$��Y	�'b\�/��F�X���O:6�ֵ	�'I`�R�+)&IұQ�E�1�$`��'��0b 9 F�X+ �ʖ0�tj�'�����ιe��T@��+�����' ,�H��rČ��.�F�'{��.�'Wy��1��)-���'RBD�3��33�F��E!��IA�t�'�č�ӊ��s��X��jCH"��'� 4��bqN��A)X�:����'6�1AL�Щq�Ѻ+�bH�'�0w��\�����Q(��\��'i@�Cdş.�HH�7�C�M��y��'ޚ�@�)U�Д�(tz�Lp�'O:r�*�9����lm�d�
�'��Q�7Ʌ[U��%�C6z�h�
�'iXU����ޅ�C,�F�J���'MV�x��OH��a��LA�8l�	�'��`	��Кu�� '�}�CF�y�e3,�i��t�C��yreU7?����*j(ÄV��yR+��u�E�o��r�����y�.SIIk�*S��$Y"g��y�JK�'���Ѣ���w���!�6�y��À|9��^5v� ��B�y��^(�pȐ���!�uE�<�y""�	
�X����7��E-���y�.@�m��� �n����C�'�y����P�Q�U3 �~����,�yrE�-V��pU�v�U� �-�y
� 0qb��/5���qMA83�Bݑ�"O����T�&����3=�0ѩ�"O�py�8Ov�}�/V#E�v�8""O��8eN�,v�<IZe!;2�@MY�"O8		�
�N�� gI��P�!"O6�� J�(�D�pd@$�,��"O���Fi��X/��s�)`�z$��"O���E�r![AD4����!"Of��S�W���H!c��Q�L]˳"O2���`� CX�"���4<yT�)�"OvI�`�G�9�����ǙC^U�a"O�*�fM/�=�6b�F�L0S�"O؄�`�\�O�����@"O�@1���E_�TҶ�̓D޾UQ�"ON��e蛐�*�Շ���p"O���\6L��˔�	�Bs�r"O2l򁣃!J�v�:�ieT�u�W"O�X��邡g�.p��n�>iQ�8��"O��(u
R0r���µ%����"O�T�I+b'э �ms�"O��B�*>�ۇ�����"O$�h���-0�Q	F����U"O��1%�>��R��60�*�B�"Oy��N�%9�tS�'ݫ~����"O�[��C)me.��p�ƲF����@"O4��5�Y�:~�`%�.<�1U"O��S�E.��=Q��<[�D\��"O�:3BIz̍	5�]b���:W"O�$�I��"b@=b��@�Z����U"OV�B0晭9MV��m�4gь<07"O�T9��ԂS<n�k��,��C5"O $��BZ+ŀ%��� {���'"O�%�ટ�#k"TC��9V~LY�"O +.K�J(� "&�`�0��"OT���&N�8ЦY��C�	�j��"O��y�JQ�F����V�6����"O���G =OPH��JENG"O|<�����A��c�GA� �"O�����6#�p�RI�"b���"One8�E�rCr���!J�rE��"Od�!'i�'輥P���4P�m:`"O��CK	�b��\�W��(9�X�"OV�R`�{֜�jR�F�37�ي1"O ��,�4bz�����"OVMX��^e�ɡ���7�ځ�"OBܠ`j�1v��Bt'܊trbM�'"O�hZ��`ʜE*u�!h<���"O:uS���j1P�A�tR��"OD�2Q+�g�0L�`�T��]i�"OLY!��3'�(4���\�j���"Oʥ9���(;jN �F?d��I�2"OD�8�.��|>(���*�&�s�"O��)��WB���C;>��EQ�"O *V��8/�F���d��-Q�"O&���.��@RD�P�h�"O����a��)�ΝȐC��R<x "O�`!.���X�	� �X4"O��#ᢜ�������v��,ۓ"O��itnVLz���&~B�d��"O�PZs왑
l�+�L}/lQ��"O���c%�y��h0('l��hR"Oҁ#��z7�}*aF����( "OԤ��$� J�4��g��4��A"O$RC�"R�떆�ony��"O� �����\�-3L�"���E[r(��"O�ݺg�o�Hm��fJ�Y�)D"O(\�cKԠa�pg�?SKF�!�"O2t�w[9�����V+��X"O�|��+AR"��u�(c�� �"Op��b�Z�F�V���OK,T�B�"OЙ���w�0��0!@�&L��P�"O�,���.D6� ���:d�t��c"O��@��mA���b@�9��!p"O�p� �C~ ��D��9�e"O�L����Dͺ]"�&
��k "O ���Y
5�|��>0���"Ol�;`oU�FbH�`�J'S�q[r"OP�9���R'�e��bA2a�H�"O}���#��=�Q![�e%�,�f"OX����*>�Hl�pO\�Mf��Ȅ"Oh r�	�5@yڕ@�<a֜��"O� �9"d8(f��p�*U	"OP
�쀣;�R�{� �.� ��"O$��q�=e�j�sb�L�t
D�"O؅����8�. �V �
w�5�g"Oļ���6yN4ኤ�
1�H�X&"O�X�/��M�VL9��Dy�,Ҧ"O�)��ku����'QM����U"O���ː<=#b8`@G@QA�P"Or(Ƨ���4`��D�!p� ��"O��8���>eu���ć���Q�"O�ܻ�L �<��bM�	Kt"O:X`S��q���U���2����"O҈�l��FBʠ�g�*c˘Pq�"O2�`@��8w��-P����*�4\z�"OP�V�P
n�$�b��"9��!"O�3��ukL$�&�B�^��"O��!0��;A��%,S ��8(b"O�D2u�ۘ��@R2+˜�.B�"O:��R��w� ,�U	�o�4��$"Ox����7%�(uڃ&����P"O0l�A-�>\��1�L�i����"OeH1�F 5�k�D�4���!�"O�X�r��_ �)��U����K�"O�ń�>���Si�= �ڄ�"Oz��ʇZ�`@�V�B�*��ESV"O�,8��EQ}��W�ߦB����6"O��FnRDɒ�E$�L�ض"O( ��%C����X���1"O���3+�\�ᴄߴf�й6"O*D �[}J� ���:ei��A "O�=��l\�%��	�׬[�c>�A"O�ՓG�
�%g(ty#�2}�d�"ONIdg�N,jT�A�
k���'0�'�b�����[� <�#�b�^����3��a������89��E룬�Ϯl�� -D�@�dD�
�. 2��7E��<��+D��K��*��8D䛄9snH�a�*D����&�I%DY �\�s'#D�q�"N���p��	�HH�O$D�(q�/^�Z���G�%+��$�R@(D��xeD
A@�b�ퟗe�x8��%�����l��l�8o�6���mC�[	�y�"OX�Q����)Z�/��{R =D"O�)�T,K {6e�!oE4/=���"O�0[��é9Nl3Ȓ49�hq"O����AV�sP�՚A��Ȅ��"O�lb/T�,�d����>�>��U�'�ў"~�� �U1�ӿK�n��#��"<n� �"O�a�t�1cj�ؑ�$�>9H�&"O��D�3�J����hr��"O��ځ�C�/.���[�	�����"Opѡ�J?<RTRc�`��(�"O,x��ğ�!�b�i�B�xn.]i�V�`'�����25�iS��8�L�WiH0}�d��5��q���,p� I�2��Wkz��&6D���ǝ!hO�U�U�<Glx��'5D��1�.�������ʫ^`b��e	3D�Lb�H�	�]��[6�6���=D�(j�kS�;��Q���{�V�i�b:D�ܘ%�ɑ[�A�2ʇ@���� .D� S�OL�H�xy'�Ks����#�,D��R(�C���A
Ǣz|)R&?��'�Oz�kG�]�+� ���l	<_w�(1""O�1����'G�$J��Q�b�%�b"Ob�KP̒�k������1�j�Q�"Ol$b�B4?�F�[��	n#�}��"O25KSg���"0���y���D"O�!ro�5�ƸҲʥQ�*�c��'�!��̱6pq{B%O<��H��g��'Tў�e~b�S!q�؈ #
�� 9��	��y�d��q��|�(
�Q*���y2��#5��آ揊���]�L'�y�Ǖ�p��-
soǤ>��2c�0�y�#Ǩ;������:}R���ҵ�y�ǘW(�9���6�>j�-	��y"��y᲍{RbR�8�t�I����y��è�f�AS��D�ޥc�%��y�G� �����cӦA�`�5�i�!�A %�|�@���(l����!�$Q�4|���3kH�qPz��\�U�!�=t¼��j��F�_Z1!���2�ృ�lE�Na@��p�4
!�DI��ބ���
 n�d�ݯ2!��ΏL����kj仇�]^!�t��o�EK�80��P�u����W"O���g�<���1�#ګs8$��"O&\�E�c���V+$H��"O�L��d�`�F��1 ���g"O���Ab� E*V� /re��i�Z�`G{��i���k�#4z�V};��K*��}"��ĺ$����Ȩ�
X��3-/D������+6
�D��x��+D��B��M2sI���%ҭ~2$�ņ+D�����Ӥ:WLȸ��� �*D��*�եs �AI�$T|��	ho)D�qӢ��*]���Q�W�(D�0�V��'<b������?���H��'D�4*�j:4����e�=h���xqn$D�k��8o��,9�'zר�r��=D���햵<�U��/��h�6D��31��X��M#F ��H�h�1ړ�0<�Յпr�>ݹ'�U"k�� ��jV�<�V�=1(�Y@'׃P��lp2��\�<	��E-��YDKM ����JNcy�'��qYc��+%
5�D�JP�����'�ep����(���mP�t�A
�'������4��r+OoYཡ�'��$����:nDʢ\�m�t�(�':��z2�D�y��(#L�P�<
�'�(%+�$�d�V���ނ|����'�ў�|�b�Ͼ-}>��%��r�� J�/O�<� ,�2FcK�z�b��w`��\\���"OF�Q��N)��l��\�(!|�""OI����_gɱ@n΅K�F�k�"OD���e�@<zE��l�;z�d0���'#�[(>P�)�r�߫=��ܙ�iE"8��O���ҝ�dT�E��!����G
�e�!�dS�)�.�qee^yh9ʡ�̲n��	A��(�R#�)b<
	���-\����Q! D�$�T�W7�~l��(�5��A�>D�(S�E�6v#t@ �bL�?�a�+"D���$�+O{��pC�,�"Yk!� D�l
v�@�E��ԃ0�H�)i��Z6k8ړ�0<���ۋ��m�B���"��n�]���O�~�8gI	I�j��'�mv
ar
�'��E�ŉ9fy���A
ļ7vf�	�'�<��N__>��;�� �~}2h��'��= �H�!7��h�u/?z�*�
�'|H�0�.�BVyV��j����'AD��-V1O��4�0�S{�J1ˊ2�'x<��%\��d� `C�"Z#6 ��'s abщ˙Z��5��c�j���'(0D�'@!@t�-F�.�q�'0	R�џ � 8T�Vo�e+�'��ly�"'f {㭍&=���K�'��!���nt~��QH�0�\`�'J��ڲ���$E��OF �"O���DЛ*�C���A!�Y���',�|cZ�e�z� �"$*(<��E,D��C�EB�8x��LP�C�MB��+D� ���>&O������5g��uA�)D���dHʀ`��A��əaI��7�$D���u�WP��#[7���Ĭ!D��
�L^_.J���&^4�V�)ړ�0<�pJřF�hy[��C�iĶ��&�HS�<A����C�zP�E �j��E�Հ�U�<a�FU���I��V�Aځ�Z>bB�	3H�v�W��gi�Q���i,B�ɫSH��1�Q maŢ��@�B�I�	�Q�YT�В��c���D>�S�O�T��p9��)��M�:0��r"O�$� .�(As���k��n'�TC�'�ў��D�'}F�A]uk�������BEZ�'[�]83�o;⡈��ʃu|�9��'��Ti#�$x�I�#M��:Ȓ"�'����.�����-�!`�4&�E�<�t)\z�(�׎	4�mH�@�g�'�axOS*!Bژc�!�67 ����V�y!�6'/h#�N/�|蒤����y�L��k�j Y��R�(f��2��A�Py�@֚	FBP�g�.�~I�P�`�<��Ɔ,M���X+A=m���`"T������>9�6e!�+^�y/84{��&D���#+�[�6U2QjP\G�,��a�<���z�PaF�<�����N�?;v0��	���с[1�~9y��B�:`]G{B�'ў�_�e��Q1��h2��bi�Y�<Q��T:�MɑE�w�0�����W�<��iZ�AVġ*���Z�<���>�p<2�F+Jr��T��k�<��!U?U\@@c,�&dƲy�Fk�\�'�?]��l	�6�p퐬��hzo?D�H�UgIH`zx�6��7�\i�`N?�OJ�5v� ���E�H|����C�	�cg�CC`ӎP��=����p@�C�)� ⨲'Ɖ�C��Xq��L*8�}��"O����<M[��. �hQ"O�-{�Ø*5�Jd0�)L'3H�I�"O@�0��n�P�Q�<~�ȣt"O���ψ3(zȴ�F6jB�'^1O��7ʛ�|��Q������,ZQ�'�ў"~�n��q�Z8��߄���0�K��yB�H�nUxy�|�Pk�$@�y�JX'TDI ���73jHSRb���y��8X�@��ԁ�5;��C��ڞ�yRh3v ��b�J�&�t}����yRʐ�^}Ρ:Q��,!ɦ�{�4��>��O@(k�1i�Xk��y4�i�q"O8����LJ ���e��`B؝�C"Or�0���A0�<��+U0�Z�"O�s!*ˎT!�d�Q⚮Z�%#�"Oh$z�c��mB�aR�W�����Z>YH�(E�g��HԂE����!(D�$��m��2\Q'"XFxh#��%D� �w����r�)�#��}m��J)D����B$Ea�]��&��	��%�1 ;D�H����Y��"�.T�$���a�7D�0I���9�z�ر�8fR� B(4D�P1LV�6���Gd�&�"�X��1D� ��)DjX��E¾W����g1�� �O�(S/X�,��q��n?hl����OBP���9����*��v���$�3D���3�U�~K�,�f�~�>@��H0D��hVD�;i�Z�i��/�f}�a�!D� ��K�m:�L�R�{#�,D����4�Y�t�W�-C�=�r�>�������R�}�B(�5�@�7F0r�l��/�!�$V7
�b��H;Ȉ
�͊� u!��4]�� ׌)x�J!����1�!�X,v�L%��o��)��^
f�!�$�#��$#_Fy���(�7\�!�d^DD�a� i`�����"F!�$�L�L%˔��*mc�YF�L�<!�$�|��`*�cMPDZT�� 2.!�V=GЬQ�B+O=$��U�v	S0" !�$ڼ,��P��
!	㢙��O4V�!���5���2�
p*:��/G�!�dW�l��I��۟'r�Cԣ�4}!�]�gZ98��V^h��
!#� Zc!��.eg��2��Ӕ[Pi�q�B�oR!�$�"�1�g��(,>�I)W�хL�!���5A�L����\�(�eb����sK!�d�9`Dd�##ț�U	90@�M6!�dH�q��3 O
�AA�	@!�U>�h�p�M�=$!3���'!�D_�p2���4�� �U"Dl_�X>!�d@:�dCPdG�{F\q5�Y=8�O��=����qu'V�h�Nc�"�T�}�s"O<ܲ��3�&�8fℋ|�����"OhdY�AT�gW��x �Տm�E"O Q�ACڞx �؃�՘BJ 2�"OX@sQ��$aa���Ԫߔ'	�}G"ONt� ��
#TĘ�&����y�W"O�͠���0$h����6t�"O䌹��vo~p�Rb�u�q"O��@ ƚ	+��l;t R�$�0��"O�U�'�!I���OY�V4F]˲"Oh|i#�Jn���`ь 2{"O�0��m�D�Ƒ��n�u	
��"O� �4{d�����Cd��qX�A�#"OR'��i�X�d��Lpe�`"O�%�$��p��D8v��:��͈�"O���pAU��Zt�2�׬D�H![�"O�,���FXP����Z'�L}C4"O�PCRJ�u�Y`���X9r"O:F�(u@H�PiE{Z�Yt"O�p"��94���e��+m��F"O<�*0�ݕe�(�c�>U��
�"O�� �Kw5���#A�]T�%YD"O��SW���� �a��_�,��R"O�q�*�5@~��;��چa�m0"O���1�=f���e�ĝn�&�r4"O����<Y�PqP�+=w�t(G"O���w)KZ�3�+6"��"O�Tʵ	
e�"��Wd�!���A"O��V)��oi>X÷�Z�M���"O4AQgf/��}��,D�k�	�_�<!!�*Ybr���M����W�B^�<)�����w+H�����F�@�<�6	RWEXm � 9��)�R�<i�)�eL[@��h�q`R�Oz�<�2a�$}a��;��B�t;�̘�(�ny�)�'u��Q3J�*Y&S�k
J&�u�ȓs�|��'MF*SB:���V!gL��'�~��w��G�@�4	X9{� ��c��H饁T+�4�)udď	�$�ȓX���
·+oZ0׏ՉQ��ȓR�h���L�F�#��B�R�l݄�#���Q��.KЖ���Dp\8@��jRX�Bg����D[֋��F�V���.^<!p'T5So���HD=C�R��4
��'?&L�q�A&�y>��ȓVE��������eΣr�l��&"O�|"a�¢F�[wE �8�SB"O$�Ci��xhj�cϜj;B�0"Odq��i_.P���ja�@,Z�[d"O�S!��$m'� z�.
|�t(�"Oh���S�1�G=}�|"�"O��p�&��vPU97�H?8=$�:�"O�ࣦ��Q®�a�O:j��%a�"O�ف��^P�X�E�7jZ�P"O�X`�oE�O}8����Oo�Eb�"O ��� 	<^lq���_,*n���"OzX�6-�|,��cj@�N�`��"O>m�2.�Z2����ޛ0��aA"O�s�⏯Q��L��f�\��"O"���P��lQR�]�Ė�{`"OH�'�8�|��2Ǒ�G����"O�hz��UM��E���14D9�'"O�m��
�$d3�(i�+P$� �Ӡ�'�1O��w��4K�%1��N�e7Xq�D"OH-[�!G�Xq�Q�U��!J'���"Or�Z��O h�q�LO� ���Q�"O8�E�P
z-uX��̠%H�<ˢ"O@Ԣ��J��PJ0F:P���"OH0�"M{�X1�",�5V��!"O��!���Qf�Y�KS>Ov�SE"O�Ś6CW��(� �?8,śt"OR0�`� �f[�� �n�g#�5�G"O�Y��4HyL0�.�h{���"OZ��������a�K�jt
!�a"O�	���j���î�|Y6���"O��)�J��D<!/i8b�!����y
� �)��M_]pw.��"���Hv"O��ӓ�3`�~�q0�=�Q��"O�a!�HW32ښm�e,bybm�"O�"�*��%�a����\k��q"O| ȴ�őhm�CDK�PPC"O�EZ`��OM�Mi�b]2:8�"OPMK��3a�`��F�$)N:$��"O
�p�9Iئ�3�D�yb��`"O��0�h����s�Ɍ�T��at"O|�0o�1-�R,r�jP9!P���"O�}A�`�"-ɈDhc�ϒ>R��E"O�TP�<Y�<PDcK�3�����"O��cF�̲s�	� ��0�@""O���s�3q��]� ���P��u�"O�{RO/w���*@ K���K�"O�{a��*]$��"�n�(�jI[�d3LO@q�f_9L�Ц�-j�D;�"O�P��E�VSr�֚B@9"O��ӎ��#fyh2,̞*���"O�D�v)��v�����)2L�3�"Ob	�r�1 �aJ�	�	4,��Е"O��5H �85����ۑ=>�#C"OR���8z�eK��If� �	T"O��Ԁ��JF���܍.]�I[V"O
��iX �:#��7T6��ɰ"O�	�v�͟S+zE�߾P�I86"O09�r*�-�
X�g��0f�H!�"O�q�����C��thqAP:|R�X��"O���$��킣m-[5d���"O>�p���1qB�:Q��:Q'���"O����ċXPDK��D�g�$�� "O�8ɧ �$ ���m�>=^h)`"O����V�Jq*'?b�R"OJ��'兯C0v�;��+1����!"O�����ȑ5�X�k!��*�ę�e"Or����!i���h�N[ƌ��"Or&��))$|��th�!+N���"O�IbC�A+5����UB�Q3v��V"O�dzQmT;;��)+�g	 �!�G"O�q�q�p���E��FZ��R"O�(Q fA>�Fl9�d��.��p��"O��P- �\��*�G���1f"O���EŵM�nb�����O:���ApL����H��i�j�]T!�Z"g���J��H:@
"$�a����!�+Ϥ���(��RhEa��>�!�$�Dʰ8�յy+Є>E�0*�'�2�ؓ�Ӓt;`�Q B�GF
���'��HWGW�O�$q7(E�C8"��'�����@� L��c��@��̺�'��-�E���9�l�+/iBU:�'��RMP'�.Ӳǉ>&��l��'�6�`�#�i��=cg��U9�Z�'�0�vo8�ؕ��5���'A�QnG)^̅�E%D�����
�';������ s�5����1C�'{jp�B,A�2�r�䗘��a��'�z�X���,Y-���Ɠv��M��'��<
F��m@
l��̄��	�'�� ¨�:%�ɚ�F�QF���'S���K�n�%
�"��M^TI�'b"�3է�6�> ���\�I{h���'L�9��Z-��P��O0v���'@�+��j�$YgޱH�@P��� n��2aܗvӊ<�bc_?�p�%"O&q� E�0�d���J,L��	��"O�Zf+7�>1�o�KK,+$"O�i(e�X�oO��[�-�L��<{�"O� T`�(��%��̴+�|��6"O���s皪z��'�U�p4�"Ot�I`+� i��z0E�S��hЄ�z>�u��{��ʡ��!;�x��#�O���O����˵E7$DhcCY%x]�!�RZt!�䇾�A��A�w ���DC!�Đ$t��Y�.
� 
1C@!�SrTTݢ��&�½8��H]6!�#t�BƩ~���r`͵����ȓb�@��B�A�P*���IҳG��)�ȓ��)��o���N���
�\X�Ib<�v�V!5���� �2+_:4��h�p�<��m4r%Ɓx�B�l�����X�<I�j�!I�����
K(z$ ����K�<�R��,`�A!��(8��bZN�<PM΍
kV@� ����\�J��@I�<���M+�Uz�"�e�p�p�b@Kx���'EN�1���.R�FD�$ d��[��?		�S�����k�([��{W�+ �� ��x<���25�CC��v�T�ȓk��1��>�d�9�@��1D�L�ȓy�lX �-V�'��u� ��<0�*��ȓ$⠼E�[��ࢆ._�<ߖ��b�z��=%�(qB��;s�hi'�0�'��>��~~V�Q��1"�lqb��8��B䉣�t,w���H@��M��lC�I_y�ɓ�_���%���F�I�NB�I�
�J��A�:!]�}� �^
��C�I�jѺt��|���1��q�B䉲Q'�8#��߽H�ȀK7��6%RB�ɂ6*lIFgV<Xz����L�C6(B�	LK8���%�+*"���wdB�	�N]�d�T|ޜ;E��.-�*B�I�v��nY|��$���$��C�ɭ2Z�
#̋9XB"y�QJ�,�B�	&R��Ӧ��HY�,r	�B䉧s*乴�F3hǮ��s�[ vC䉸u�IeLǠmz´�W�[�m7B�I#p@��c���
lS� E�)g�`��ȓ	T�+�cV�Q�����D$
gpD��V�D5Xg�Y(/���c�R�����R���{q`�5�u闀E�]c$�ȓx��Y �',(yt9	#��n�4�ȓ5F�5)fb�<ֈp��jY*���[x�-�r[�p8L���Gŗ�T��ȓ:Ơ����=%�0�3`_(U���	p<�r���[�n��6�:1����Z�<�d"��%����B�J=~���J�k�T�<aٞe�H1��5Q��qІSv�<��i���s��X�pTFą|�<�G�2K� �9��7C9
��cAJw�<)�G�Ych�pN�2]-P)�`��Y�<y�	=?`!ʲ�6ӆ,��(�ן���W����� �T���ȣ8pb�����u���� -�srg@!R�.M�ȓC�lh�NN-Ll���u�D��ȓb �)c���"����#ER�mV�ȓ_L(��7�T�x��h�^�ZȦ]�ȓQb&����B��v S�1�L���)���r��U�f���AC��`-��	ҟ��	�<� ���E&\�� :��̱V)Mi�"O"�j�m�=��O��[	B��&"O�eʶ�M.+PL�B卄!��
P"O�5�#�$���T��jU&� �"O�H�BS�2���b/C�EP�< �"O��f�Ã4V������%X$1�"Ol(b��X��*6�\'-R��'��	�<	�(�=����HV�Aeʱr��v�<a��ˡ �Ƥb��
*x�`�hq�<��lO�~�V�:�"��?�bX��d�j�<���]�L�C F��)�8��ǅ�l�<a$�P�A�٢�3��<x��Vf�<q�e�2Ux+w�Ҹ*�򁳐i_�<�q��n�6`��5��H�� U��d�I�ϓ6�F�(�DO @�r�nKK�9�ȓW�*U9�AǛe�"U����YX���F��PA���Ѐ��o� .tV-��!6���c�@����#I�L�~���bSd�Q��9_pH(U���x⁆ȓX1DRP�N�<�%��n$|���|���k�55��ӧ�B�T�jx��s�,�Cfꂟr�r����I>;���ȓ?PIaSL�T��-��HK[L���@����������i��E�ȓj=�����X� Śȫ��D������S�ۓ@��X2�@"Pq>���o@�]xV��8m6E���� \��@�ȓ����̇{ �L!�E´��ȓ#��C�A�)@����2�<��J���,�;aU�	@��8��q��!��p�(��\�|�����7R �lE{b�'=��*�A	Ǧ<sӪ�u��;�'�:<`��f���i�"�p�C
�'����⎓>r:��SL��r�ͣ	�'�$t��)���j�@�� �kX��Q�'�X4�<FxF���`C�j�x���BT�dD�������T��5�`�8v���hOZ��D�%��(u���p �"�8=��Oj�3O�Y�#9Ѵt�.�	6zU@�"O���6k!Ʊ�2�U
"�j�"O��R�F�[�&���B؉d��"O8��`��3�����&P"^\�\Q�"O.EJ�X5~�d�3%啜D&��A"Or(@�"6`0XR�� ��"�In��S2Ώ�.\���F(`l��5D�3�aNW:�dZ�R�#5D��yD�S�/�X�n�<�HE!��2D���Mk�v��a16YB�l1D�xB�" ��i!�b�.}lI�Ɗ0D��@�m�9V�$hc!��}`A��,D�������
��6Ԍ5�<��+ D��ɗ�T�J���ҥ��"7�ftqǀ D�0�э��izm�e�O�o��l:�J2D����O?���D��s��l�ā0D������|49�fV*R�^�{Ej+D��e��1&y���Œ�"�`�*D��C$�]T�E�#�[�a�����+D���En�>
�(�Z�Ԍ<Ϟ8�'�<D��R�&W$iJMb��^P&�0�V�6D�ț1��:a�H���j[�nt��5D�Ps�Pv�c(�1U��&�lB�	>T�dY�0`��h8�tAwB�C�ɸx ,�`2a֎&�jػ�o�>E�C�ɝS`peⒸ��� ��XD�C�)� ���RBC^��1�&��K�:K0"O~��"�ShpF�9 �Ly��"O�UA��[�CY�]�k�S�*-"�"O�a�H�1)�����5,�n1a�"O4�0��6Nn1a���Ru�	�S"Oڐ:�CLWF\�ꡈC�"t�( "O~X��� y�"�q'Դ!O�!R�"O  �cI�.6��ؠE��a5Z�0�"Oй�$�9H�P�&%U�]ȩ
"O���/X�`-�q21D
��q�"O���� �{� �D�J�y� ٸT"O>����}c�|s�͓/�J�"OTrP��MJ�ձӫ�8~7*@!1"O�h���	r�z��3�C�,���"O>=2��^*&A��k�9'�Lz"OD�3�lU�K\n��`
3'����"O$ܠU`�$?E8XBe)ܳ=>\aB"O(!r�U�{��s���;0����"O�+�j�ip�t�g�M�$t �E"O�P�$/�"���4��.�A-!�$�/�6�X�)ڥT�
�C�/�|!���X����6���>ӘL�FM5!�$��0�4өD���|%!��U2a��ȉ5Gܑ��T�b(VH!�DU>���E��=�Й�G׫e�!򄞜_ݺ!HK( �̹�'�]/!�d�sذ�!���*�Ȩ��
�S!������\R�g\�E�hhY�'m1���G��)�ˎ#kvt�	�'���S�N) �ly���_0.`0�'�:�Λ�u:����߮ehz<h�'���rE� "^�!G�HZ��<B�'s\���-U�T�G�E�Nj�3�'i�p��DuPV�̊}���
�'��7�ӏ:�
��V�Gq�L���'���Kҕ6��(F40`1B�'�i;POA-%��{��ɉ��̀�'d�d��
W
���/��tr�'-�M���hwbH��܃
�n�9�'F��I�e�@������'F��`�Z�'�`d���S�{�H���'�~�I0O�l��a;ƃ,y+h���'���SM��$��&_��}J�'��J)S�xR%�ė �P�x�2�'j��3�*	o�p�@�υDaҌ��'>�M�B��="�p����H)"����'��	q�ʔ�He`�7	Xo�XX�'�.t�u�_s�]+�J�Q����	�'}zmS5BC#[& �C�H7�,`	�'K6��K��g���b��B*���'�|HZ�@�@ܙ�qCY�f4�F"OA8��ۿDg*9�'���eP����"OX�y7g�a�pT� ,
B<�a�2"O�2J � ����3MG�%kf"O��1���6x��X��jS=%7T��$"O<����0{Hx&j�)px�v"O�Q� ��L挀���h"�""OF�ۓ�I KI,�3�W�l`xR#"OR}T
�O��l����Ou��1s"O�y#i]�_x��9��	91�)!�"Oܴ���
4C\<�w�A�x�v$�q"O,�{0��P\��;�n�5i^�f"O@G/��.P���B�0��QC�"O����`��7�h]��G&x���"O� �@S�y��5p��L|��%��"O>u:������h3"S�:�2m�S"O�<���PL�B5�c) �;t"O:e���!��R`@� @v���"O�P6K��t�|�{3"<�G"O��s6��f�L@M�10���"O� � �d�Ѣ3�3�JbO,xCb�%�d�)�B�+'Zn�"�m2D�L�1'�J9a��Q/J�TX�`.D���ר��W䖕�R�R�����b*D���"'ȝ92芴D�f��C�&D� �#GT%/�@�3��(���
WE&D�x�6B7EmxE�1��Jv���Cd7D�l�&'Y�s�`����}%���5�"D� g���(&���S�tP�J?D�D:�.�y�������$(��	+D��m*@Ҋ�ؖ�E�
Yi��,D�x鴣�q��9`ǃ�hd�йb*D���IN: ��"��>>����.,D�����o�$�祜�D 8+W�(D��xS$V�F���'��N��}rso&D���E/�V?�}�u�
7=	Xcm*D����MCu\�"啺;$���j)D��3&�ǎf�0���a�en��G�;D���r.901~��� G)sV!J�c$D�hq�%VK|���o�a�D��#D���5=h��X�R�I����$D��8w��C��dV'&k����Q�-D��0�'�^պ}�F���<'ޝ` ,+D�܁�ڴ]��*Q��0gr��X�,(D�F�U0N,B7	��QH4 �&D�H1D-��S]�h�2� Y�2�2pL$D�\Q2@,)��X�R�[�.����	!D��iΚ�Z�vL��CY�zZ�Y�s�)D��A���&u��B蕆i���S�+D� �`܏}����sʒ�V��!a�)D�8�d�AF}�9�+�G��h�E2D���GS>%�e�R�'Y ��$	4D�0�Uh��q� ��6�Cf9$�$f1D�`����7m�M���n��4�b�0D��U�U�|pY�V�H���q�0D�H�� �/$k\��W�=���f"*D��(�U�d��lzã���Z�f(D�lY��	B'PH� M�-x\tq@`9D�|k�\6Dr�ᱢ�FL9#B6D�l@�-��Ȑ�K��ʗ0҄i��4D�0s�� �u�C1]��D�v� D��+"JϪn�H=��H�g����&<D��qaHl�Ԣ#oĶ*�J�Z�/D�l�
K�����g��O�X\��+D���'Z/(��!�L���~d9�)D�d���Y�yV�a-e�|�[�*O�\�@(5�"-�f.7���W"O��� &Q��m	�k'>��"O^lA5�
I�zdqVE��=n�p"O�ūR�̬B9n-�W�=[д��"OX�Z#�Ίlh"i�di�7!���F"OX'�ݵc�����i��Hs�"O� ��nT5O�Z��a���Kr"O���B�ԧYH�i��f���p"OZ��Т�-Z�>����]-�xX�"O
����5�B�Z�G T��k`"O� ���>���1G_�'���S`"O�LЖH�;g����u& ����"O� �p��Ҏ)z-��oԡ� "O
���iJ�d����X8$�v�"O�S�J�'����@�"�.Q��"Or�B�`ۿ)�J�V`�(�8U"O���F�-v��|pv$ܲ���8�"O~����Ń���F�Ǉ�L�2�"O^%�+J1@���t$�=���2�"Oz0��>I���IG߁.��Y��"O�ec�e�
'�E�� ��|����"O~aa���B����eK�4�p�1F"O�@���,;��p�wd��8��X��"O x�7��.�.��Q���9�bՠ�"O�Ad�
cغm����2��xA"O�-y3HR���E�K51��$c�"O|�2ӎ�p�:� ��:w؈��"O��i�m°?Jα�a`�;�����"O�e	�	�&T�vΒ�z� �b"O�r��6*S�����V�)����"O��#�V�}#QC"F����"O|�,N_ި�SB	hB���"O���%��b��H��'ΊW����"OLQ�A�_�y�0Ȑ��?@J���"O�Q��-@Rv�����
<Nx�T"O>m���Òi^Z)�c�	v���F"O永&�X�"�B�	�1M�@<��"O�u˕�ʕv������А)��U�5"OF��L
EX©�[<R��m�"O:�pS�ؑn��"�LմQ�();v"O��R�F[g��cѭ�.i�F"Ox��1�� ,PZ�)��)c��� �"O�T�Ît�C@� �D52"Ob��� Üv�Q�e
�N���W"O���`��=<�P�g�W�VuZ50�"O�PZU���E>>袴/-jHarD"O���!��A`�U�68d6L�"O���bO�z{谧��u�L}�F"O�-�3䄆e���T�h�,�kf"O�l#�n���Xx�K'td�kw"O�k�Е4y��AD:x\|	`"O��P�F��� c֊TE��Zr"O���c���]�F
�c��yr�"Oh��a:���ӱ%��-����e"O��[U�"/.ڜ��#�w�P�K3"O9�Gl��G�N ��!M�b����"OҐ�d�˛RSD���I6����"O���C��<J�U�Jޣ`�!@"O �F��n��ɉ1\���e"O�A��k��&h|�� -K�\~���"OX<
ݙ#D��+ë
���x�"O�}�bO��]�`3��8��(R�"Ol��K�[��e@n� C��-�V"O�X���F�����H\�i*�"O��B�'e�Tف�+�D��%"O�	�d��^'�	�W�Qm�FB�"O�
^5d�����o�ne�B"O���p��}�&cbi����#b"O��Ӕ�:8n�(�&M��@چ"O����ûaU��K�JEit"O|X�횸*��%�V�B�`�p"OȘ�d�Ȅ1�4A�c#*pAt���"O2��S����a��؍J\d1r�"O����o���y�1�Ҟ,L0y�"O�0*�j�0N��:&P�R<�܉"O� �`[�~]�YɖL�VΙ��"O� h�X��yJ�������7"OX@.��1l8���I.��}��"OR�1����Es�HH�5�P�� "O<IQ��##�8�`A���^��s"Ov̘0(�?w��1�؁��4�A"O|�irŒ�=#7蕻3�I�@"O(4�b$�i��DI$��~��Q3�"OD� nZ�-�p�Z"%�F;�D{�"O@� �$��b�S"&q&"O���ù#�
@j�"
g����'�i3�&}z���)��M@�	P�',� `����&�P�nC(���'��� �ӌ�*���O9q(=��'4'&�$q2��T�!8���'��4��ސa�H���6�TT��')��+ҫ�VZ�����50YP
�'ŸAR�*[�wfԡB�ߴ�����y"*ʬ ���ׁոA��yb���yҬO�L���ka�L�O.̣r��"�yr
	_D��o�'?����bB��y�+:;�rH9�E�7a��Ж�X;�y��z{���X�`'0܂A�L��y2�\"��0�"��R�~��`)�#�y҉���\�R	�9X3�BU�Ҥ�y�M̕L���N۪P�����N@=�y��
`�EB	�F�����ų�y�"�;���Ң�,���ā6�y�
��d�x"��'r�(N��y҅��\����ḇ�J��&�P��y��]�{��0���g�8�em �yri�d�abF��x��0+�D�/�y"�T�h�xh��	m�R�� '�y�ʅB��D�����]呒�y�*C�=�j 9��9#��Hpm�=�yb-��(Fb��@��66�=
D���yR)�%�#��«y��%)���y�#G�q�2z�kǗ?�tT#C��1�y��^�:SP\
�I�9q@ԫ�ʃ�y�I�* tX��O*_�L���V;�y��ޕXB~�ꦎ�_�I�6&R�y�`ǣWR>�� � ��X�K#�ybʞ��Bi�Qj߂}ц��yR׸c�"���]H�ӧ:�y"��.�Djw�H�J�Dx3д��y�J��i1�AڭD\^�a����%�S�OϪ�9u�ߺo�2����
<Y410�'�|�d� !K�8J�1�� �'Y�����iD P��d[�H�
�'���IHU����*�lK�#��	�'y�9��K��0E�,�d����h��	�'��axv�\�bx�R5$T�	�m��'��������]�}4�b�'�d��e���pX	F�@��'~t"�AE����Pύ90f�����xR��@�b	��uG���¢S��p=y�}2�K�M'r5��س9��X@�C��y"g@^� ��e�.t~H����Ol"~��+^::K�}I�dMH�M����iH<������ѡ�9)?�d	��-��ɚlQ��|�`D��hU���1AF�y�#WcX�,GybB;Dp|�𲮊�X�n��`�������<��yR��i.hC���|P��VB_��y��^�s�<0!�R�yPH�I�cX��'�az �\��B҅J�z�&����'�az
� &�Y2m�7|jH��P�D� wO L��é��Pt����%�uL�����=����8�I�p'��2��^�w-�-ze�& n���U3��'~�\��R(+
ک�w	�	P��u˔�|��)擞
��Z�H'��ɡ&�=G�.C䉺K"����0XWP��(�?b����!��'t�a����a�V�s�Ă/Z���'��|Sc�I7'lΔ5�U�/�p�JA�k�<��4J��P� ��x�Q���Bn8��Gz�+{W���7��3�8�G�G�y��P6=;�mk�휧�\xc���	b���O*���iρ���ֈ�Ú���'�����$f?�q�A���s��	��}I�*�d܂2{yK�a8S��Q�ȓ.R�ԍK�8�J�P+R� l>��ȓ/K߈GK����R_�E��E5D�����({V�+$Å�����0D�t{wf��@�B�cÅ�jÚ�`��#D�D+��� @��F@ �g�~̻��5D��z�c\;y�l���"x#�D���&D�$�ʏ�,<�A��-���rC�M�<���%�I�"*p�D�L6_�I
#��8Wl,B�I�yG)�q�ֽI�D�B6��9{LB�	*�M��I<'N`�GI�A8B��q*Ԝ"qj����03��v�,��p?��H4j��xc�n+��hr�g�<��"Z�6p9�t���U����	`�<��M�͔4�0fǍU��te��<����$�Ot-
I~
�'���O ��Qt�I��(9�'D8�*tfD+M�p@3�?<d��b�P�ЧO�D��O�T��+Z�vv��[����Z�pY���'�Q�L�.��q,쉙���d��XP.F��y�d�R�H	����I��XZ�E��yҎսNżaye�Pu���MJ�yr.L-Et.E"�#V�t	� �����=q�y�L"9R���WŘ�<4��W��yr�S��@B�š�R�k�K���'ў�OK,�*�@2+M��{p �1�\��	ӓ��'$`"fF���Pp`�&?�Pش�y2�)ʧ{q. �e�X)>�외��5\�-�O�7m(}RU>�}ҐiZ����v�Ņ_z��	���I~��UE8�@��+� j�1x���,(��͹$e�Ob��ԧ(���kh_�>�<!ʖ��=�VU�ĭ�-[��B
�'9Dq݈H`��@�	$^� C�R�t��X~�@�k~���I
lxb8Bg��̒�Ȁ�y���-:�bP���ڭX��ȋ�����5C�1���T>�'�� :片�qOJ��t�Ȏw��+H>������85DԼ3����h�*�e�!�$͖I�����Z�1����c��5/�O���O��ɝ��-+VaЊ�޸x���.N2B��c��	�vEƯ\��8�����N�'�ў�?�cqi)S@4-��B+�Y�+!�O`� �'1���J6L���.	m���y2�'��3�k�	%)�1k2Y�hol����?��u7 T&��q�G��NѴLq�ꈐ�y�߹/��8a�9=��T�yR�;8�h�b�D��)9��Vƕ��x�ő�@��mמ"f���k
�!�D��Wy>C���,!h%��E%!��
��PH���0$ ��'�'|JqO���$@�4Ϡ���=o��X$�� �'��#=�}��� v�Ęp�!�9 ��0�X�$$�O�|�d`���R�ԳTؤP���^x�j6C��c�4S����h�-��:�O��d|��� Ф�W$[�C܄�h��=V�$��"OA��֥u�^a�r	��i6ܱ`��';�O|UA *�(&���GطU�>aR7�;4�����[��Y�� et<��f;�d��(O���	�ea�ot0�Kb��X1�a"OZ(�Ц�*q|d��@D 'ԍ��>���&�	���Qca�:~B� s�ǝ&D�1��1D������0݈���
����"-�D;�du��u����$Sx��Ս� 2m��hV���y��);�r�sѥ���(���`	��/�S�Oҍ�T��y��!���.W+�ێ��7�'��y{q��:Z#ZpJ�#*8ɸ��ȓzU��	�,J-5�H�f(�$2�F{"�O/� [t�̊x����F��X~��B�'a��A�o\�*H4��i|�&���x�S��(O~�=Ab^�}|��a��%�H�Ūs�<��(���B���E���Q�C��r�'��y���C�`10���*|���1E�š�ybB�3h�`!�PnD�nd>�Ҷ־^�':���'��yzp���!����d
�tS����'���ʗ]�z���FX�X��5��'VĨ�%�O%L�Ѩ3�V�f���X�'�h��!M;�����ԏ0�v��'&V��U�_�*��a��A"t*l�A�'1ў"~B7��� X�H�s�N?j�I��r�<	�@��a�&��!�=;(L��Qd�<ɀ��*t�| cV�Z�2s�%�e�<�P�Z+8�r����ܔb�^_�<AC��4��QQaJ٥ F8�* �]�<��ʯh��S*�#/�0t��m�W�<q�O�sM����^#6o���F[�<!���5}Ӏ��ǌ�tň!����\�<I��4��\��/ˇXT�"GU�<�S.\8�R�����%�,����P�<	���_��Pc�)E�8�:@@w����x2�حsp�t����_��y�
gp������i��M���y"�[�Ii���$�;eN^ŋDjY��y��\�
��XZA���X4���G��y�)�7G����R
[�W���N���yB�X:]DV��3i]�D�`��H���y�C�B�&1��7�A�#F�y2�¤skԠIr�-+*��A�)>�y�ɋ�g�(��i�R ��d���yD�>m�u�� AX�31���y��" ٙ��H!Z���-�y�-�8�bM�C�Ǌ�2�#���yr�Z�?�����M �,TD:�#H�y���d6�j0�X2��W�y�� Z �8��� );�C�8�y�&�P(Z�+�#0��9D�
�y�#˞׌�k�WĔ9I�@��y�b�.m���Ӱ��4�X�'���y�H�����ʋ�֪%���@��y +m��ɪbʕ+O�4� ��N��yG�>�$ՁI��?R�]a i��y��P ��{f퉗9�N%��c��yR�ʎ70l��t̞/	��`e%'�yRG� Xl���k����)ܒ�y"!��Jjp�pŖ ˬM�� ��y�QML�
6}�=��#��yB`�.$�s�E u�FA�/��y�NZ�f��E�h��衴�?�yrB	E"`#v�S�f^���#Kܥ�y
� <k��9Y�bA7l@	$w�][2"O��q4�A[��X�G-
�`���e"O��(�"،<�\���#��L��"O��j��|���R�
�~��K�"O*��E�@ [��	��ڂ,n�]��"O:���/Ò��e�$�
�c���"O��)	�!�|��4���~S���q"O��Sg%�OYq�Aa6S8�D��"O
M��D�:q��u`��+�y�G"O�I�Ѵa�J�2�l[�&xYJF"O44Zl��}(xd���ևfT0q�IA���jG��>�� ,A	)P�ɛ)����K	vl����8$C��YھM���Q<i�V�c�7�lC�ɛv�J��JS9*���T��&5e`B�I?`��ᘴn�RW��HwbO�&�B�I�w��bZ�4��%��NٖVY6C��'p0iyEaڇ|�B�PT�ل@I�B�	�~�~E�M�x�NBa�=�RC�ɑ=r&���MHr$k�덒*��B��]\rB��*,$X��� ��B�I�_Ң�#d��ps2�I0K�-WlB�I�?d��{�"��YB�)��I}PB�	�WiJ���c�o��۳&@�#�B䉽OR=���ܰeĂŠ��ޕ^�C�Ix����fS��Ƚ{����C�	�\�"g�kN����Y�re��dD2p�&,h6+�3#���s(	�b(!�L�BCx��%��#iʸ�GfUD.!��*D�(��_�-X�
�f�9!�E1_`�Ғ��~�J@�R&W�!��Z�r=(�z"�6��!`�&)i�!�$9*�� vG^5oJ�"0�I�Q�!�D*]춈ʤ���FS�8Z�Û�?�!�d��x7��ǅ�T|]:���_�!�؁cM6�Fi\�9h6�+���n�!��c�����I	�΍��cJ,C�!�$��<%�@�4�Y$���ke�X�}�!�d�fq�l�P*�;jQ���;�!��Ő'����I r���堞�0�!���Ȳ����z�]yu�P�!��JYH	�vX)��4����	t�!��
0h#���M�4�N�J3�W�h�!�
�"( ÆʉW�1�p�kb��ĝ[�p=i��|�x���y����ȁ�̀C������D��yR�8+�P���
 r$`r��؜�yba��g�U��׍]��0Ca苢�y��˿@�z�2��8�ʌ�`藾�y�,P)ij����J�"���T�!�y��z�<t��Z�;�@{�i���y҄�f�DI1�0�����<�yr+ٟx4�q�N�v� 8aE6�y�ԧ|n��w��0�R�_��y�-�+\80�!�0��)X�O7�y�b�GHH��dЪ�p���舐�y2�88uH��QH�p�P����ċ�y�R�\�v �gN�?kz� 8 �y�J�87.�"Cl��e��#��
��yr��w����gѾYk�!b��N/�PygT$uh�q�nQ�@�ı2a`�q�<��ϭ<c��(�N˝>���a�<T�ьh���jEcЭ.���Qa��G�<)�d�o���[��+H��YY�v�<�.� )�����H&M%�\W��j�<� >�Q�m�嚹8����'G��"O��hq6^�^qh&��6�"OB1�1K鐥s7��#W@=�"O�#@C��>dh�BƇ`C:x�F"O"���$D�W�w5J��q"O&��&��;���D�<=6$��`"O����F��@8`U�J#4՛E�'"6ѓUGOʦ!���V�����W��$�FL9D�`�6ʓ�8cD��u��	#[h|2�I+ʓ#��l��S�9aF#|���;bWf�Q��/���&OS�<y�LهFpX0&����T0��WȒq8!� �`�!c��O��}��"�j}�&D�@ܮ�r�!������5�E�%)� �Tp�e�Y�O��mZ�i�"��[/2���� 'Qd�x�h@�;�H���C�D�4��Ў��=���$�6�CQns�S��d�('�;�^I�a��Px"
P�;�89���=KV�@5�B���'*R�:1�U�Z�1����>����|� G��M8��'m $����Co�<A�lYJ`袯K.leh�G�&˘��TA�*�ɂц&3zdF�,Oz�R$�
i���j�hX�X�#�"Or�����4�bg^.))(
�̵@B�s}���R�؃`�p�?�c�2C�"i��Iy���p��b��tQ���T�ZT؄�65��Z%/�5<�Θ+�%F'� (`�+W�X��ɞUd���j�;v36�(6�c�+vM^)<��1���;������q�T/O*3�
�@s�L#K�D-����.b� aA��@N?�*I�t��d�(C~H����,8+��Rhi��c�:(BؚF���*H# 喧�uw���q��O�
\��IˏP���!��nPN���@;%$
��S�4D��+e��v�X��i��t&�a�w�=S"�,"��	�:��Q:��{Q��U�N#p�h�Cɞ$q,�}�7e��?�҈��d¦���	��|�B�.LOF���ٽ:|j�'B�%R�ʒ^OZ̻%$ md�@Ag�#%���U�Ľ[FȀ�� v�1r�/j>śE�P�o6�l`��66k`���1X1OhҖ�4T���RJ2u{��a>�8��Q�i:Π�E��2����2~G�ႂ��Y&�%�a�ȟW�:4�W�'�
=A$��B�:���vc���MPBM�ix�䟫vR�8p7F��k�)y�d܇H�*��̃ui��&M�E�.���"�4EW�lYG-Ǘp{��k�'&��"��P���p��Ȝ�:����d�#�	�1�&o����so�M,��ZR͐���X�vH��<����O.��P�ۋl�� 9&DH5�V�3	ۓ$Č�Y0�������e���>a��AKÜlZj�����Ll����Fɱ�$=(�P����S'���l̓L���� ��l�2c	�;yL�>	ѥ<���OÀRX�eڟ���\�����O�z�&��%�֣ а��Y�,����[�f5���e�B�.]j `���}�"�+���*�F1�r�bx�������J0QO�|���_%���N��A��y��A1��� E\/���c"O��K��V�2����|��h?y�*�u�� ��o�2<V�uE��d��iJw����K���ɀ8̞���N��Iv4�C�؞ ��}R� ��ۑ@�R�@=��,�Af��1p�)
� s��Հl�6]1DV�D#p�4�g?i�YX�23�h�&~��qJv�'Td��d� c�'}��Z�O؞Dܰ�q�-�2��I,w����$�
 �鉊\��Q@�hX',�"�N�e�������l�:f�_��s"3��	S��`2=���2D���*@V뵠��@�$���+��T�"د�)�7Y���Pӈ�#+�)�t�ϟ(�H�ZA�P�Wt��PD@ɀ�0>�#$ƣ O4����Q{0�1L�JdQ�z�80A�4��nJ�Ed��ߴ�ħ(�1O(�(A �%h��2dO#CX&��q�$K$;;�M(1"����'9?�E8��z��1O�=G(�K$���R�֡�ߴV8�q�GH�x���D�")`ʽ���:d�*�����8��5Ң�]�^v䤧OT�KtŌ84���I��iat$�F*t�kL��0��h�ƆJ�T80�=8�!�V����S�_�R�� ˗eЗc��,�>C���+5쌳��ɴ�:ͫ�jY��'Q�,L��!ޓ^?��z��U�q]�m���'���G������ҍ�)�M�D�U�I<��B�'���!�%�\~�%K���c3��P8���5�͕
��lARC$�x�U�<���	�O�``гm�2�f%Q#�"�[.9bN�zrF�
*���{Ȝ�"V�"�B�Pj��
�'��|���T8kɔ���2��=����5\����?p�ê�":��`�@ U;nΞ��O�N�E��m�f.�*pC�f�9e�a��&��}i��RCN����pԸ�pNB�2�&�8�Ũ,�8(G��F�&�ɈA@���O �bL��:���H����/ ܽ�B�?�A�hz`NY�$�*p!�N�`�dh���?��<�R@B�lJ���<\�<�ci�O")D�''>2���S�? �ș!IӾwt�͂��XB��ۦ^���S/�*ɖ�PF_6tk�Ę��_�9�hY�r蟛���8=�d�j�%[�D��D�F�8�ΓcH<�c
����D%�~
zQ���=����)� �S��%4)d�]?9��G�6� ��Im��]�n98��6(WX��Ys�r�����3D��Ͱ��ܰ)�p�C��ݤX�����I� f�-�k׹|�Q�����Z���00��Ot��,W�X��'�62�ˊ�r�H15`�:+딜���$��`���K��R�6M�R��qH��țA;@� �c��`פ_�t���IģTϟ�0Љ�sG�}h��'�^�H�IE�d	���H�7��y�'(�9Po�<A����+r+R���b]��L�C��O��b7D?E�5[�Ⴠ��9��S6I�#��s<��_J�)��@�A�24���"sz�݈��!:Ĭ��^8�G�O�$y�� �D�*�@����������0�,�?�Tl����f~"�'�p�S�A�G\J���"طF�ڝ;� _�15؜ 4%�.(-�q�i]�s� #C��BVZ���bضE�εk�����D��7հu �+�BO����MYlQ�,j͛�s����+zܚM�� 4��Jul��a�&\k%J3�Lx�E�,W�x�(�,B�4W�� �Z��=ͧW%��˒B��~�����I!��'P��>6,�I
�����UQ�U:�N�٥�MK%�ؿDږpX��V�4�`D�u�Q) �D�{�-I�hO?m�`C_'����)i ��ehf�h;BkE�S�<�#`⌣�����0"�D0y�8*�Z!��̼+sf�,?޼K�D�>9����v~��'#H$0��C1��D{' ��/Q���ŀ <>��H�s
`��e����^B��C�x�_h(��͈�h�`r��>�0D����8ʐ됼8FY�7k�W�H�aWC�0b`�����6{��i���Q��͹�	�#D;���AY{o��=!��Ի|v�erfHP�s~U`���~
�h֛-��TCR�]&�Z!h�d�<iw/�{�4ـ�Ǘs����C�<�'j��
|h	�ʛz<Pxg�S�e�h�'�5n�0�c���B�	�3p�!��Ő1+|&�u_�Zw�C�^B�Ĝ� ���~&���C��{P�1g"��J�8	�B�74�|)�a_`�����뛹t*^�p��ؤS�����|}��)��W����&Ϥ`���2d��pr!��G 9��yđ�~�%n
xqOց�H��0<1f��(�P��H�.x�ЩK�AZ<9F,��2�����r��j�2���s�<��?9�h
ps4ȁ��H�-/��Z�WA�'���P�; Ȳ�$>�����`� pѡ�W?B��1E�5D�$A��B1����C��M�9�2ð<�O�Z*ZI�$*}���%K��ŀ��1qM���,�:M�!�ę�l�����@2-d��q锘���O^�Xuc�*7+��qOf�'b��{�t��v�ǛS�z$qp�'Ul���"	b@Z�r�O:e�	�⥊Z2l�pvUi؟�bR���u|З�̕J�l���%�?#�i0�޼0R.���Xw�N���D�L?~̀��"O$�X���k�術�����*�]�����<?�2��S�>E��%�(�Lb�B�.r�60�E*���yBB ^�z(��fjyt�{�ƃ�^&�'���J�DM$��ϸ'����4i�%���G�!
�]��'����E#$_JX����5g�^�J��SX~!R��'�:�J#�X/���[V/O�CY9!�b7����N9�=)b�1��lL�T� 1�N}'\B�I�g6Lpr��îs�����L�0B�$E&ґ*0*ɲ��0
�=Q�B�	}2uis+˩E�h�$��]�B䉒$���'$����JL�B�ɗ ���Q��li1Q��ON�B䉂LX�C1�$��c�푰%��C��:iNq�aOU�E�x�5@��|B�ɢC�	"Ƅ�?�v$�E�4B�Ij���鱣��'�F$X��� A�"C�I�&*����¸&a�R3$�+enB�Ʌ9�ɹA�	#j�UY�
[,B�	+u��4��T���8�r�
HU&C�	�TA��c��4��`�
[C�	� �I�a�71`�(+򀛈9�0B�I�7�|��o�#$m��C�lB�I�q�J����0S�x$�Zd��B�)� ��CQ�̮0����P-GѶ�r�"O,"@�<y �ᡄNKo�y�"O^e�J^f�n�A�T+;6�"O�}���'��E	�ٷkɎ�K�"O|��D� 7��̓�
4 �NB�"ONM�� ��q�쐉�`��L����"O������6p�r��
a�}	�"O怚��G;�6	&ș�V�fh{R"O�p�a��\�f�Q��C�|/~ub@"O<%�&c<{�T��fv��Pa"O��Ф<���`����PH�5"O���䖞3�-!4�5[B��"O"Aٵg�<�Z���ɳI6 a��"On���8~�6PQ���+$/0�;�"OZ��u��r�jT6'C0���"O��z�k�5n8��B� ��e"O�i�U����C���{.�#"O"�@�\ �����Zu�%�"O�9�Kߙw�<���d�?'$Q#�"O6yk��4AW
��1I�On�"O��0�#@?����[�i�T�"O����� I堰8a���%&T�3"O�7DM-�r���j��0?j!�d�/O��<)�jF)zÁG��!�+P��+��g��HB���!�E>'e���˃$�P��@K3�!�� nj�h����]�N��S!�!��U7`W8Y�]6v��yb�Exf!�$*8:\�[�ċ'Y92���=4�!� �.��e�ٹ"�Vm��9z�!��@zx�i�6�A/`��D��,��!��2%0��*��%�(i3�E7�!��-0$��Q P-Gt��ڃk��!��֡�	�g��`!��(��!�DK�!0nY	�PjD��(ػq�!��
/�bM���� |�4t�A�Ӡ	�!��}��� @灴=�BH"�I̓:�!�d��qb��ՄS7 �jP��+T�!�� 'n� \����Gɢ������F�!�$���ip�$"j� �;B��8
�!��O!܅���B
VU��Q!�ȵy��$H���\̼J�LSz!�D�<��k�CQv��ŀ�=x!�dF�H1�(�T�`�"D�T/!�$� �e��(a�M
���Ga!���,��$
2��7b�V�k�̎6�!�䜣 ~��ӂ�<2�0@BaKQe!��;Ll@#B'��1�$|��AȪ�!���$y=��#ק�@�tpk3�=�!�J?v��yL��9�6<��@W�5e!�Ƞ����D��4F�l��<2�!�ѲjWnhF�@=G��A�t���O�!�+.��s@ÇY��:b�*:!��O���\��cƙ*n ���;{�!�DV�U�H���J�/�\�qsKπl�!�D_�6xP�k6{�����V�&�!�D��<"���Ց$��EcNߧm�!�䉌�Z��+�@<mSW�ۨ"q!�Ę6x��;+����o fk!�d�5}��Ά(>L�DS� 4Z!���ODV�V*�% [�%��ŐT!��E�t����2`GZ�ˏ!��P�<�z���	`:(��W͌�h[!�dW����[��/���ѐ�W�^_!�� �a�2L��+Ԕ��EK�;�REy�"O�XXƇϒ?�p��E
�+���B�"O�qr��6lI!�	�*���W"O��	��@�s�ڭs�JR�`�6@R�"O�%b�ϝ/q(�9ؑ��\�X=�"O�,r��_���R"o�"UpQiD"O����`�,����@٥X�!k�"O����f�n��1�V/G�7��m��"OD�YrI��@�^�8��/]�x��"O��� �@ u�,�g��D�<*�"O� P�W�+tPBd��	lBLZ�"Oz���aM|���9�nU�_�x�$"On ��
��E�Bq��O��v��"O�HbwGW,h�P�d-��|�j)R"O4(&���S[4Q7L �o�v�jf"O�`�@k��A`p٪���+$��S�"O�\ �+��@�Hae�9Q�eJ�"O�9���M"<R�Q�h �X�X`�"O��f�kh��H ���^���I�"O.qB��ŜĒ�F��R�.���"O2eR�&�5��cgNاRwX�X�"O*z��܁���"�֦F��h�"O���O*n�<Pj�l��A��!�"O��ߒJFar��Λ'�:�#"O����ɛ1�f��¨э
�y�g"OT��f'[yܺt�b�ą!G\���"OLa����X��hf�`�!�I21�Hi���	�O> +f��l(֔#Џ���iKcØ0�~�朁f9���:d�,I9�@]�S��@�#�3sy,�S�o�
б$���?JV,x������l�	���h�d�ұ�wdL�,q����>B�I�,��\¡DU}	������*�(��O%NPaЇ��|+T�B)�7/��L�ᄕ�~���BA%����k�8k�ă�k<d�ƅ@�F��{��V�oV�*tΌi��9z��J(&\t��1h��6l� 0�n�#ϸ�2bEF�FP9c�q��1r����(�y��!5ڙ1$ʎ�2<��i���'52ѳ��Gf���dd�)Hx � 0��6J\yk���9|����Ф�s���z���6�@��g/ݟ�0=y�&�_7��Շ�;�>(B��5nf���#M�[w���1i����x��ǬZ;�(��'
;�4�$�j�q���R� ��!�)A�~�So�1DB�I�H8���
&a'~ArRh�]_��$��Y.�x��"�ʀ���ȃN4�!��B%g-pi���^Z��Pst����M�,�.�˰���v����c��YA�V|l�K��?��<Y��!
��1��B>vL���Αw�1@��0�(�s���?�C��D�z;��C�֐	���3�D$�OD�`��C��x�{6�/"��%8Ř�^-ǚ��Ð�.�ڰB@$�q�b�	�4 Eh�+�*azB�[+��i�HY����u�%��ʚ'	8h���1�yZwL�����D
"maT,�=Z����J��[uo�1�,�T����"OX3���@��߯y�`����O$��;�r�%K�$q���W�A G����=Q��hB�ODV]K�.�<X��mS���z=��gҀ��Ƭ��5��ŏ%L\K�$(Ѹ��aA�gV�Ty�T�L˂O-�g?�녹w�d RC�l|���Ǡ�D�'�ڱs��M�'`7�<��Y>���K�D�R��8�I#h9�e�)ʸ1I�ȇ�	�F��@�l�!F6�q���e����D]����;ȉE��gl�=b�PY��a��Y�rh'D�p��@"�v�jP�Ҕ%�F���������ԃk�
]�{,a  P�];�)��A�EfAh��	�;�b)@�+L�0>Y5�A�\dJ���H/.����?2����\P�
$LĪI*"�#�)>1����\n\n�j�S4��'��@���@��)M7��@Y��^+�>��tGBH�S)�:��d�_+|nP�&)�J>��%^�c���n�+�.����Ɇt��z�B�iC�l{$�%M�`-rN�%_-�<���̴D&8�'�P�B��n�Np�ܴXI��V�׊�5,3}<���L�67�|��`Ϝ �y�g\#pmL�Ӫͽ����@M�1�?���<��ܳ!̚M��,qB��烘t�Sf��g%�)�^�iC&�y����8*{J����7���+0�󦝣_/�ұ��	;����I>?qw͓p$",1��3OR�;��»k0H��2d$���\���`�!ϔ�p`�����О����6c%�-��ܒ)�ě�+�2*��顁���J�%�IZ��ҤG�h�Z5A�
�<W:���E^(HP`,�v�Փ�Kş(JD��/�%+4X�>�{�? D�A-]\Ox\��G <�S��'�Z��#n��Ȩ��h�$	�veD6E�&p ��*X��y�Pʆ!SFPhCdKb������
�| E�>Qn���I���@	�%SS��[�'�p�O�"$Z���X��,w*<k.JQ[�Õ�?~^(�%T33Bxԛ��T����'E#yWN!#3�'���r�	',��1�i%H��ݱ�O$,Y�.O�J�&U�ů�c�d���B����$��M�,�.��� �O:yP@���N��ԛ!�9$� ba�P
j!:��'ȑy�\�F���~�i�>9N�D�c哵Y-��H`Z�o �@�D=O�����$�7BE�Eɐ`�~���^BP��E��`�t)#�@Z�>ͳ£�^RT`)��3��� �?-0^-��'��iĆz���@�H�� Ŗ4r�ZĘ��C�J�G}R)�
\tyC������©t� �h��5��ᆬشn~�J��B�i'�u[a��O�]�fg��aa$�0<ɖ��;� ��U0`i�Ph�gDs?yF敍c��=+�e2=#�m�&.�ekH�8F�X���cBٴj��WF��o �s�N��*7|봩V�r``C��/uAv�0���Ѽ-It-S"zx�B$G
���mڒG�&�Q"G�/tDx�Pa�Ѷ)��R$pv�]5Y�>u���߿_ļ9�R퓁w�b������p��T���u*2���� =v9Ī� ���Hx����@��dA0@��_V,�s���N���1��D~�(�>E�bްt�H���*��O.ȩ��(a�c��KV���ÅÝ*��)r�ʕR�f����4��o[��R��/�:b�n	s����0<�ԆF�h����%���^�NH�2HA[}�L�C���7
�A�D:�C[7B���B�ɭ{/�D	�4HjfHs��U�݃ŉ�'�x�����4,h,��#���B,�����*���l��3�֠���Ĝ�%*E�п	B4 c�L;�\�!��[�T�әw$� L����s̝�36�y"	�'x����"/���A�0d^rai  9O()��N
+�{F�֕��I�wPdP٠�x�����j�C4`�-���!�Cy�a}��fȦ���� TMzE`LI&h슶䙥�h$"$V��*e��M1T��RF�(2xR��G�W�G���D{B#S�W1@���-����a�s��	$U�
oK/:	��1�=�yBG�4���Oſ1�|�闏Ο�y� ]��P�33-}���1dg>�X7�=�3�;uвu��/;8��хȓ:��L�gN �8р��1��@��/K$��ɳb"V����L<)T�.2P0�m�3�B|bc��mh<ɕV8|�4�bt���;��c��Td������0?9�	�Fa0�o��`�詑uF�y�<��
H�ĩp���;N\i!e�Lܓ'����'D&O<L���0b­a��;NQJ�8�O>D(�R?>�%���ս{�3�ʽ5M*����:�Or̡�a�:���� �Սg^��W�I�I��*�cñW6�OE�����C8:uj�ƅ�M�je�'A.`+P&��
�2FM�-F8���.O�D��7X��N��|��$*A����� 0Ō���Cq�<Ѷ�2*c ��菪;�����o9�Tr���ጠ��g�A0Ṯ!�ԧ4*P�T%�}�da����C7@��!6q�e�F�M�ح��ɍ"fv|;��'9��懖U2�*�fEW�a�����PNA�DKȚ��'i�>}�ceE��8Bm�m����I�$�WᎿ,v�x1O�\�'��|�ѢD8#nT�OQ>U�"e��̔�D��)r��I@"O"D�(��Q�6SuB%E.x�բ�
���	�]���5#T�3�	�{@N	��G/J�pT	ǀS
�B�I�zDD�qԣ��F�a�R?Cz>�'��E9�}���R�썡@E�8=V��׬�M\���G��P�y��o�
�@���43�F`h�S�yB���Rt�e{5��.q�y��B��y�+׏lf�9P���ht�A[Ҡ��y�f�&'��Ggɤk��(�A��y­@�fR�9�!� u�K�
���y2,:��M�g����@l��yb��1�.D2GB>a���yR��&&0�r؅����>�yrD��~P�T)T �#_��鎥�yri !3�bX[5C(@����kڏ�ybn��r�����q�TrN��y2��yzi{(�/wux�8r���y��?lL���R"2@�	�.���y
� Fhr֥�'M\��!�%41l�3"Oļ!�D��-�tq�m޴,x��"O�}ʓ"[�$0��D]8��"O�(b(6��!I��V*����w"OvA	�O�&%ׄ4Yd�7D��Ep�"O�)n��[0�131�����"ON�!���:E�H�*da��{�"O�ds�'�� aF�Pd@�8�̠�"O��Y���wؾ�A�@'w�Nt�"O�#բ 6�x0C��F~�@�"O.��F�%��\{��<[����"O"���_3������M@��"OB���
'X��d!1h�6xOT���"O$��s��R�(y!g@�M=� *F"O|t���L=}��,y��H�}8$�d"O��C#��lD^%+���hK�"O`�ȥ�kؒq{�ƆV�l$�6"O��ґ��3Y��X $�(H��xc"O
p���(w�0�0��<7 	Z���,���O�ax,�W ǧF��I?g�D�0L\�	�|8��Ƞig�C�I�g�.$Ӓ���j��1��q*xC�	;�)��b��%nۘwΘC�Ict*$P���n��d���"�fC�	�n�P��"�J���-)>C�$���*��>?�Ub��;x�2C�I%ӈظ�+����"���72C�������=-a��93M�)q(��HOQ>��%/
*<�������ovZ��"*�Wt�4��#\:
�h�ɨ*�]xU�~:����O��8c��G�Q���a�`��L�aY�m̳Y|���6$L�фX��I4�'w,rA�W�V�g�U�a��* ty{�w��s�.�:��b�w��S/:F|cf]"B�x��0C�:r�^�Oz�� c��r�1Oq�,6h�)3�2�P�,@�Ml���Q�¤b�3 �4c��|��c���1�*N�Z��<!��D�(i .^�p�qOQ?-RE��5$,$�ҍ� >0pɒ�U�XK�{rY?��'�O���3��� �1�dN"�>e��O�3Z���鱟<P�	[x�S� r�OM���V�HA|VY�'����{Ǥ�o� m��k�&��1�Qp���`�O2�A�6O�dJ�� ڼM4lx6YԦ�a��	7�D������?A���#8V0j�m�*�)z�-���M�p$��Fl�IGcE�EN�Aۊ��'JR䋆:�!�Cܾ|��ꂚ|�c�>�Oq�bL��O&,dR�qU"�u�\	cQT��Au�5�Iֺ�?��ٕ;a���)W�`����`�v�<�p'��n7$p��(D)Aܐ��c�t�<�q���M)�a��	�y7��brFI[�<c��,P��$h��(T��B��|�<�e�T�?�Ę��� �"�p"���v�<1!��o�~�2`�S��Zt�EI�<i������7�M�mw
�+�`�<Y��}�4��UJW	 P���wdIr�<I����z����l�![x�#u�Mb�<�,X�q����c!���.�cr?T�0�� �<%����U�9r�)q��6D���f�#'
r3)�c��[El1D��@�G �(�`3F/7F����3D�pc��M�yX[�V�E�3��$o4D���e-�3ԠD��L�R`�1� D��Жo�"=��4c�#�;�b[e!"D� q��4B��H�󥄤Rg~���5D��
N�*:A8��R �5l�E�� 4D�hk�1���� /H�҈���7D�ԋ�^�%&xY�D�Sڍ��e8D�����7<�	a�I\���-qU�7D������P>�]�ժY����r�9D��ɐC�[K����
T�w���f9D�`�$� ��z"mR8>�J@z��� >@ڇg��J�J���[i<���"O�x�FE�\��0d�M�H+�"O�9�G
�� ��Q��ˑ?4Vջ�"Ob �)�zp��〤�� :d"O��b��P���Mz��I[�ԁ�"Odܻ��S���U�ӣL��h�PA"O�l�AR�q�S*c2���"O���qc��*�`�W��%)@�q�"O԰6�ʴ�x���� �Q�"O��"2��X"}Z�J�#�r)�1"O8�;v��by92Z�&�`!���y�/��Eg�aQv	D9�^�aG�-�y��ƑE���V�� ��@ 2�y�%F{�`��B�fa�U�^��,��`���
�*�	���� ϯUXJ��ȓ^��x�
�#����.}��ȓ"P��0D�@~NM�cl�EK���ȓ[��e�F]�6$��bFF!���/&����Ll1�	b� ��x=��84��8E�ڰ0`�A�.�(6���J�} ��sK�a�(E�@��'~>��Z#�L��G�3NP1�'���r�m-$�t���/͍/���
�'�ĭ���!E!�Mi&�3*��C�'�F�%N� �S�K).T�z�'j:�9@`�3Q��l@A��i��}i�'%ܸ�ug�=��:6��L��,��'��M�L	�g��ʥ�!=nʱ��'��؈�m	�_�8i��ě�2�Zh��'I�0�Ķm�r�t�	q:y1�'�B8x�*t�0����?R8��'�~�)� %������3aF}H�'�J�10�<c�����N4-��Ё�'�4���mF(�zup �Y�%n�e��'�rX�bBԬ|�"�j0�F-�Z��
�'��]��K��D�k���!�V��
�'C�TE��d(؃'摧�0a�'$�UG�=Y�]��B����'oB9��*�v)�+�	�9�����'�����O����V�,[�\��'� ˶�Ϳk���2��U."`�h(�'�n}���ȴ�pX)����4D�LA��0s@E$���]����Ï<D�hʰ�"(^��Ê�p���*O��)��ץ�ʝ+��#D����"O�-3�i�`��㯓�H&�Y��"O�@�A(�=,Kj� �m�!Ć	�"O�Y�d,��9�V-��-̥
�hs�"O�q�e��/߄=I�U4SZ�*F"O�m�b|n|��+����5"O�!����'���� � [vH�qw"O&�[W+��8
���F�:sR�I@�"O6�"U#۽Ƃ��s]�<$�DB�"OV��s�P?,��"��A�ld�D�#D�X�� T��p[��z#�+Cm<D�ذc�y?B%�t�Y� �,�F�:D��t+O?.bz��-�3j�A�#8D���b#Rk�� K�k�!�� S�a5D�܉f�݆Z�r�����^(J�ktc>T�T�����@�X�:�BM'k��x�"O�����$H2�;#B���H���"O�� �-�1I[F)X6���<�"*�"O������ 34(h�p�Q�"O(=K�䝵hW�q#��Q�/��\B"O� ެ��Ϛd����݋N�.�$"O$tg'�$/K\� �J\�$� a"O.�!v�Y9)z0H����!���"O��4��o7x�h	�f!�|*�"O���t��Es��+wf�
"O��`A0��Ł���+"<T�s"O��*Ů�&�,�CeJ�I��� "O��JseX�zU�!뀁Л5ʾ���"OH��+ҤO�����/$�h���"O�=�b�K�G�sa��;���)�"OZ!R!h��.���ZR"՗mX���"O�	��GZ��.Ÿ"�& [�"O��;�n$mk�\��H��"O�	I�d�:D"V�B"KH9.�ъ�"O��b�Z�6N&09t�ҪF�d�e"O*5uB�<�*4C�55��mx'"O��J�N�5٤���M��Y�%"Ode1-͘*��K��8�zh"O�5��Cԫ=+d���'[D��V"On�)2�G�5y6)��R�8�"O������F������?vcj��"O؝I �� q۬��B/ߪ%Rֹ�A"O�$��bROU���C�Y2�p�"Ola����N�䑱���:!�,��"O:�R ��u����u
�4o��m�q"O�� BJ�L�|M`��զ?Զ�"O\T��(���T�#p	����H�"O�@F��6Et���"�({r��"Oܔ�����,(��̲A_PDp"O�0h7�F����ID�,�`l�T"O����%��f��ߑB� ��"O���s&ȣ%�Lа��=
�mJ�"O%�#<i�ppׁ]�S�|��B"O��3C�q�@Mc�b\ *�����"O�|A2FL�-⊭*cl����i*�"Oz����*3.i�I��v���"Of��pFY"dL�b5���U�V�f"O�Ȋ�%J�E�d`"�J�b���"O0Q�"ʐ�WHViy�CI
K�P(c3"O�@��b.m��Pk��8q��tY"O�����X_v`AZ�e��M��y�!��͛ � �%Ұ���Sf�D��!�$֌v4ʡ��o 7�6(�F��lv!�d�7������=q���g"NWd!����q�	L2!ɠM���F1`{!��4n=Rm`%���	�����@߲]!��g0���#�_�	
�$F� S!�D��&l`�eBt#�{D#��$A!�D�v&���l��XAzQ�D��~!��H$2t��T&�Eˊ5�r.K�7a!�$[�57 �	���=z��(T,�
0w!򄁇{��u��o�y���1f��k�!�<r��]i�G �R�@A��H E�!�䆔%І Kg�>i��ᵁ��k`!�$��(Ƣb7AP�W��]9ԭ[�^!�Շ_�QǤݹP�`��vl�%!��B^���$�$���t�F��!��E.4�~9�����3�=��I9�!�Bop����Q0Bn��r.M*d�!�(�⣕75�a[��|���'�h�v�<t"2�*�`r
v�*�'����n���ܱZP����H�'����Sf����f���q��'h.��׀
4K60�qt�ق}�t@
��� R�Q��<��3aA&(��IS7"Ox��Pf>*^�����a�"Q�"O4�9�lز����h 5rL�"O�����֦O�A�G�#L�n�aS"O���ReU7*���@�26��-Ä"OT):e�Φc��(�#`�5sX> {�"O&�dn��]���'.k�~q��"O�Ȱ�ӎj'2�+%h�i��8��"O���� �7L��1'���)K"O��i�����\����"Ohhad��.���A ДJ5"O���M"k��C� \�@�f�@�"Oցc&�Bj�"�.D��pf"O�H2�A� ��1p�Κ�J��F�V�<iC ח<�R��s��>~�,=��CEP�<��I Fp��zW�>09���E��O�<I���=��\���S�^�FT`�<�'-ã+�\�H�MLj�xf��_�<A6$�?,�j� "��D�5:��X�<)�ғh�t�b���X�%���H�<Y��&SN�RУdֹ���{�<qTJ12P��Ė4�Lp�6DG^�<Y��P����ꃈW�d �6��R�<�0�3q�F�@�^i��d�c��L�<�D�p���p5��Al�1����K�<A��N1NG$M�A��Q` �c��b�<��J1��<B��9�i`��B�<q��[�
�du
�JI�]yQ�S�OU�<��m)h9�)�@H#vLd$9ҦDR�<yUL��b5�cR \O�A(��r�<ѣ�q[p���MRżu��p�<y�Fܳv��qɤ"��F�KDoZG�<AeIBr�<p�]�t�y�@B�<	Ң�@� ���YN�q'�T�<1� -$�EB���-AwV}��H�i�<1%�1>�|x�ñf6@P��b�<I�H����ѥϒ2Z���My�<�r؈Z;���a�H6t��+@LMt�<A��	;as��"��c��S�̘J�<aiJ���Y��:�^��� r�<14膢6���F�\l��"��j�<��IX��5�����~Cp(�ld�<��C�h-Ii���b� 5\.B�	� hl���L����r�`�=)TB�	�X�r�����7}Ϭ�B6hī��C�I9y�L�%k�{޵�E&k2�C�	�C��u�hQ Yd��3����+,C��/�*��2$$��%�r%�f�`B�	�U��@  �P   /
  T  �  j  �'  �0  �6  
=  eC  �I  �O  EV  �\  �b  i  Po  �u  �{  g�   `� u�	����Zv)C�'ll\�0"Ez+⟈mZB%8牶7Zn�D7sF��aH�-똅�#��n^P�Ĉ.~�� ���DV����	��o&U{��	 ���'o¬�a dW�~����
��V�
�[���F��vp2E!B��a8��4��R�rԁ�&��*U�0��I�u�݋3���m�Z0#n	%ye��IG�Fh QCڿLh���4/�����?����?�� &�-�ᬌ�\��e�)���j��?�'�i�7��<�����C�'�?��>E"U�v-�J�5!�A�=\E��	���?!,O~���<�CĎ�a��'CBk��"�@�3��@�8�I��#h@��DG|2�ieʅ�Ԋ�W�:9`@`@�r.�x@Ǥ>9�'�'U�� !��)a���r��w*D�)�����'���'��'��ٟ̖O��X�;��p���޹G�l�C P-%��h�^�o�1�M#2�i�"Fi���o�!�MKV�i�2Գ]sj���Ɏh���e L-�ў,
��)��<dY�q�I,IV<UoO4>�ֹ�C�����Ȣ�Q-�6-P��q�ݴ�R�O5L��T*[B���Ǎ�j'x5 �j��f	�D��'��� �eH|@��)RN�]�$�{�ː0� �i=�7m�����%P7>_�u�WMV�D�PQ�@hJ�M uP�D^��f�R�4V��f��|S"�`�}S]w@�]�uI��F66�!a�El.M���%*V	��H�*����Զiw�7M�ʦ���5Z~r���H� �(�*�K@�n
x�����=�te�FA9;�T�޴!$`02��Ю J6, G��>L
�Z����E�Q*�aVM�%��P�"�?q�B�'�ҏ$rM&7��O(��V�	�j�!q�%^��\5aH"G����O�ZR�O��Du>�(r�=��X��'���=;$�7���6�Q*f���U��Q�|��&Y�R�rb��3�P@o�<��\ѷ�D��,c���
U[.Yʀ�C�J���0�e�OH�$3?�oI�o��\�S"m�)Z`�W����	��?E�TCX?��x�0��:�D��o����?���'��-�G�%�F����YW"�S����'t�ܠ��iq�Q���0��l��!��#a�k"D�!��(o�J9qN�z
�Jk D��%�����g�S�|�ȑ!1� D�X9�)�0#��,ڱI�7S~��S>D�(:�j�]b5iw�� o�H��`C/D�,�0"�8I���wAǙ}nX�� �O�phC�)�D��d�D�/' `�({q�E��'(�|*�ߍ��1����)y�`[�'���cW4Th���ϑ�?6>��	�'ˎ�iσA#ʨS��;�@�	�',�2q/(s��l(q��.@���'p�����z�*� 2%�2E�(Oҙ�'��:��a,�BVOȖI�83�'cf��lP*+��B�
��|	��'����I��L�!&�%:d��1�'��${ ��p�$��%���0��M��'3Z��"eB�C�`5�ul��.���ϓe�Tݠ5�i^�'aH���jK���p��X!pn��x5�'�"o�6G�2�'�	A#���c�lV�V@yeF��f�Z��E	&��q�dL�!�4%H!EXA�'k ��7�_<J8�DM
�
$맊���]���� H ,*�╝.Ť#?���R��I��p�I�c�`%p�(��nn��Xr��� n��'��S38n���P��Ē�{揍#�t����̟�H�'_Τ�Cj�,\���e�O4�3f�.�'�y7�
1H�(�;��J�y��{E�>�y�c	~dMA���x��������y2��P�&��#�	u'68I1���Py2e�
o!��D!K�'�^-��MNt�<A�ۓ`'������I׶��E_n�<Q�i�2Xx<�
T\V���(�Mc���?��xӂ����̀�?��?�ӿ[�EJ��Hɡ �+.�p9� ::�� ����8�rm#�a�� ;���F �C�hج��#��d�BŚ������ׅ^N��%����(����It�2\�^u�r��6&�A���%�'��ɴ ��D>��O����OF�����~t�<8uD��<�8�&�=D��X�		�PY��ԼY^�wB�<���i>��IFy)4i�pİ����c�,=p!��l�@S�+�1;���'B��'�r������|���ܸa"I����&�L@�%%N�����.��{��9�zȩb�&iwdH�!�[<AU���d�r,�C?��℆��3��	J<�����UB؀����'oIv�h�EP�<	q��Q5�x+�o�p!Th�WJ�I��M�N>�(Оs�ߟ�1fi� ^��u����**�F�s�ǟH�I%iyΜ��ܟ�ͧw���U�H2��]0���P�6�� ¼i��c�a�uǍ�s��'���6��&����2,4*�B�rӼ���@/�2��VO��0<������	m~�ȓwPZ�j��° �&�RU�����?yӓK� :U�ƍ_l�(�a�T�Z0���	 �?9��QrWj�ۑ��氹@����Д'�6x��'��>�ϓi"��k$��M�A��k�a�,�'����8��+ËȽ_�f8J��2)Ӣ����J���&�^P���ɽR����w����MO�k��}����b�1�G�������~�nG-�����*G���}*��Z~�U�?�t�i`x6��Oʒ���iե+ʉQ�j�>B�,���Q}����O����O.��D�	�1��Y.$�ʅ���n�џ<�����Xlh�+ǏI'zc��(��9���?���*�1G�,�?����?��{��,�Y��qkf$:UƂD���C��œƌ�>�?M&��|�<Q4��^b1#�d* 20r�Ovc�5�6P�@�gݲE��b>c�4Xt���)�� ���q@��"$�O��d�O"��O�c>˓�?�"���Zt!@w��*}�iY7�^:�y�J����11�)]*}`��&f�0��$WX���\�M+-O�qP,8G+�-)s/̠���K1�Ȁrꐬɳ"�O����O��H������?y�OPazQ��;ZU"q0'��$�*�p�b�hi�<�6#�5���=,Ot��Eˏ�mϾ�kpj�N��=b  �X�$��*W5"ü�J7.�}X�T�/T�vƎi)�� �!B�Ae���X��d�O���:��X�O� ���/���B�jRh*���'0*��i�j��t��J7`��(M>7�i��_�a�-�8��I�O��0�OC(�D����@�� ��O���c/V���O�擼)wF�P����P��uQE� ��M��M\ 9\���A&U:��i5gX����&h(�1�����`"ݴ
�r� @�^�_A�
aNA!�x��Ɂs���O��E��Z󪉿HKm3�%[�kD�M'�8�	[���a���@�44��.V�]p��f9�Oh�	�J�5)D�>�6��Ҧ͑5ھ����'gFA���	s�1��Y�>�(�;u�����s�&D�@i1��[���)f�Ķ`S:Z�'!D��2����	�0��j��E�`���;D��*3(���r$��z(����7D���e���x����B�X�g��x�;D�����@Ÿ���D�mT�โ�O^T��)�'h�L 1�%�LH�d�����'>b1�E�D�NV����bʺ`��1i�'x�
Q���B'z��W�,C¸�@�'��4��T�OaLm�ǀ��:�Ƹ
�'� �Ō�]��[�B[�h�	�'�`�"��"1ƍ�$)�>�L	R)O:����'��`S�� _T�t��N�1�h��'2���j	��l����=)�FpP�'4rD�T�*�PV#����'���cvGV�L�p ��L^+}l�)�'?R!�P)�,� �T>��\�
�A=(��gp�K��O�n��P��q�j��9�f|3#�		|ت�+S]�(1�ȓ=��yK�ސ$&h�L�3*��}��Ub�����^�L��	ϯAj�q��'� 5�w�\9���±?04���W�:�s��*T1���I��PE{�*
��p���?u�|���@���M��"Ov�ѥ�ȞC���P�Ղk���"O��p#["�����G+fj���"O�������Z°��e.2�<�i"O�đc��^\q��)<���a"O2�	cN�X3"����$r.�r!�'��z���&�F��t`�GR���2������ȓضȳ�dڅnHb)��KX+`����Qh��qE��5���&i, �X�ȓl�h�*BL�3$f��Y���Ipa�ȓD 
�;�JD�Iް���.#�\��e*���枃���"F'\|�&l�'��Q�SCX��ȨeS��I`�K�6�\t��S�? F�Xsiܯ:�,���F�HbZy��"O��IU�M!̩����-�
E"Or�`rLE�����R�D#	T�9�"O౐�.�,v�����M�ji�'"����'�E���[^�\@��l�X��'�����!���u��`��-�'B�jE��r �1��U��h��'���V��0�)PF��s�'�YP��_�V�Ɛ!���4���'�D�A�dN�s�� ��������b��i6���%`�8wp��7��!�������n��=8����!�$�VM0A�v͚)pLe�LY��!�d�%lk��r%�N�iT��k��!���:uj�B2x�)��U6$�!�ۉaT|�
��g�<U�#,�7Uq�*��O?Qq���B�ajUX%�I9���T�<�,F?9�hTC?L����R�<�@̧F�d�%�ҕu�<bgBJ�<y$��()|̂v�W�T���Jz�<����	#n�x3&)��VVLz��A�<���_
!#�[q�6d�j:��ɅO����+��]��)rx0l���Ķ!���$-X����E=�X-$��5�!��f�n�a�֣ln���.־:�!�%'n��B�Gq]H�Q@�)j!�?�|,ĩU1cJ���A^�WL�}���~��
'J�Q`��OVx(*�k�y���U�m���V�E*� c7���y�	6egLp��Jt�n
g�ӑ�yr���¤k�ֶj���S.�8�y��.8�$��Ӌ1�p!B���y­�i=vhB$@����)mXK�ў�!�3��lE�� �iZiP7��#7����l���A�$:b�$(Yʸ��F�J��bY�t'$�!��?v�^�ȓ-[Z�r��}o
M�aù)
f�ȓ9R���JӷS�fu��
g d��a&83�e�%�����ZێD�I���"<E���:]9(h(� W.M�^�s�+a"!�D˦��d� o�"0�\�x��9p!�D�E����҉Y 1��uC�� }!򄂌Y�V�;�i��y����l#;_!�d��S���\)4���DPZ!��-k�̕�� |�rf(\ d��	�'���$+�p�B@�����-B?o�!�$���YX!ѓ�-�j���	�'M6Uz&�E`hb�3�iUQ�� 
	�'
��
T��&����A�S- ��p��'F* k��?��	���B��"�`���B�f��"Z4�n�)�c�ai�y�ȓ{��H���:y`!c]�M�ȓ��5SF��S�x� `J�3քe��hb�U��A#	w�ha�-P9G�؇ȓ �U�,F
x����R��0�����Q��qf��s�z�R�Sf=ZG{ң�+����@x��Ⱦ����юD%\���#"O�ȁ�-��F`���� �j�P��$"Ob)��m��4B�X�# ^�"3BD�E"O�=�ЋzȌ�"4�D'p�"O:عf��N؄�Y"�%��Y�"O� ;�  ,UX���ρ�N�L�yV�'���;���w� �2��:r�R�;��U�E�V9�ȓW���+���%g��8�*OS�h��S�? �t�A(���څB�r���A"O���&f�=�P�KD,قaR��Z�"O� ���J�+2�\�B�D�l�S"O�-�$�>4Ez�*��=����X��+�.�O��rb��87�!"R�H�+���á"O
��E�Uo�u�#f�'qj�"O��pk� R���V��b%l	��"OT�@UG�W��ɹ��W�)���"O��g��=W(x �ȍ���i`�'6���',r�X#�^�!i���s�U= Px�'��:S&\�n���oJ~e)C�'��u��܃&�@z�/� r��i��'�$ s �@�R���U!b�"���'��}��G��14���%��07��Q�'&����W����*Â.�������]6G�Q?�rE ��r@����<�<,�!	"D�`ô�-RHy�T+�;G�
tZO!D�8s�A�a|Pp�d��ع��>D� vF�U�<��J�@k� ��>D� (�)A�&xLs3�	
%���T�>D���s�	6�~P���@�j�X�"�O"m�D�)�'7���B���:FdDW��|��'5���+ �f�)g�.KzHdc	�'*蘀�  !�zhVn�7G����'�p!`@%O�a1N��u�B�C��(��'QdH�f�-0$��F��B��l�
�'+F%��+�',�p��єI�v�H*O`M��'*0Y�'����,|�V���<s|��'=������&8x���ɍ�0����'E>թ�h�>�Y����.6�C�'���t`��
� E����ȣ�'�,U�Ӎ�duF�[��H(~*4�������dJЍ�F�����9UA��rT�d��EH���	B�ĉ��%^�k;�M�ȓ&����!�8 � 	� =X���*S�:�@	4�9��8|
���mz�4"�'%��鳶d8�b-D�ܹ�E�Qb���D<@�6�Rtm(�^���F���2n��(��iX0.��[@���yZY��Ȣ�K�.G��Y�IJ�Y�VC�I�=�b�a""�//���
�=�2C� 1�\��(��u��L�6L=C�	ni���L�%q��SDț8�C�	4>iT��fK�'2&h�O"����
�I�"~R�mQ�* ��B��-�d��.^��yrlR'Rt�1�ˀ�Z�2ͪƤ���y��Q$1L
��p�B�B%���L�yr^�WCL�	cd�48�v�1����y	�m�=���+@�̢%ڍ�y�E��FX(��R��y}� �`H�4��2��|bI��x���(z8x����'�ybM�]B�����q~,��7Ǘ��y�UT���PFbRmlꖅ7�y��J]���HB��Z�#6��y⇄�R(ĩC3��5��ek�^��>��*�x?�Ŋܺx$tB�j?>M:���P�<i#�
Va�L�E��[츀abL�<�$Ϝy
$�����{�z����`�<є��94��f�ق>6&�"�^�<��$@�A��+7N��|	�av��n�<Is����X�g��'HD̑baWn�'F,aJ���[Y� Q���^�<��{�+ �!��M'TB:L��gT�R�.=a�	,E�!��J<V�]��Ͽ��p��(��Py
� � �N_�#1$Qb�kF7v�Y �"Oؐ触J&}E;$�U_��P$"O��2�T:%h��0l�Y�M8��'\�X�����(c���q呇��b�Ŗ0n��@�ȓMf>q9G��GrR$
�YS��ȓ>�q�'<���/�,{  0�ȓ/s.�h!E
	T �#I$@v�t��U�i��"G!3���u�ß:�p�ȓ2�������v��"��؞s�H}�'m$\����<�wI�k�x52�dG	'�C�ɏ5���4j��A%�X��ɴh�tC�ɕ9��Q�p*;7�,i�bI�o�hC�ɳS6~��B��#�x�JCD��/�JC�IBm�Y��#�5M3�i��T��,��$�f+����{��ɈTo�2�H�鈰y!�$�T��!�WꁟM��%���=yd!��T3E_|������+D،"��\#V !�䘺E/�� ņt��Y���L�*�!��z[h��7 ��T�!�Fi{~=jcf?@YP��#u�ўhxf�%�P��c A�vH��!CL5��m��lhƀ{���*x�>�s�&@����)s��x���a��]�s�D1T,��cF���G�bg]�F@S~І�+zDj<0�$�"��`Q�X�ȓ ���RÓ�})�l��$�T9���V��"<E���ܡ0���q&���Z6<=H��Q��!��6(,~)i��/ �x�G��;y!���$�a'C�
f���&�k�!��f/R$Qw֕HR^���+cv!��T�T�P�I�C7����%a��3]�@)��5�Lp����B����_���Q��D)/�N�FT4�'v�uRGc�&��pXc:*�P��Ą�t������(
�d$>{`MC�L�b��f�K�Ye:A
��;�I`D�1s�����8#��Ĉ('r}��m�&π=��Lѯ��O]q�'���V�(Ze�"-�r2��23��ay�	u���"PG	�*�X�IG36bl�g-0�O��'� ����*F�ѱ��R4��,O��@�2OH��0�3}��ƹb#bk`+��y�����y2Ǜ,2����AZ�aV��S�O2�Z=!�0�;�F�'{�Nȝ'+��|v��h kڥs��)�8mHГ�@�M�L\��@�~��ΓJ��Iٟ��䧫�䖷sJr�B�_�~Ix4�Q�U�w�!�dծG
���`� �uR(�kF�Y/�ў����iA�M��pր���VJ�nB`m6��O����'7�2(����O����O^�$к��e�*%��	�<Rx]ْ��G����.�H�[	�(wʺ���I�n00�Ɓ��W�V@СHhUXPkr��ڟTc��+�����!)FxR�ͰR���5)0q@����d�7jS��'Sr��h>� ���� �+lN���'�!���BB9j'a�C=�A �?���+��|�����U�1��*�#I%R�q�'�����@�@W)9��D�O����Od�;�?�����f�nגe0Qh�@H�@&M+*��Qp�.]/ ��(��S��	Ó^���y��"e��@
�U��l�T�J�W1 L`-G=���2���{���A�O��P&�8lҹ��F[Y Ř��O��d=��z�O��㡠	�f��� 
n����"O � b���c�ѓ�Ȗ}�db1^��C�4�?�.OL0�nB�T�'��	�-m����q��],�QE��-���J V��'tC6W!r��ˀ{]�ק��%3�F����52A�hE��O���GR3c�Lؔ��{�SS�d�"�02�H��UPR�#>1Q*Vş��J�'b4���Kj�����M�{R��'[a~��^��\��)ݏ~ޜ@W��>��Z��b�(ܞ&.�ܠ2���,
X%	�d�<9%��&�?i��?�.�z�	���OD�$�<kk��5��6}hP��Uǘ�$T���)g��Ԣ�Ĉ2K8NAA��[bdz�O)1����DOW��}�F⊢"���V>O����S�|Kb�B ��o�n�Aש�A�Ok��렩��[�
y�3閿
uX���'�<���?9�O�O�)� ~���a�u�4�yB�/r4�7"O�����N(�Z��4)T�&�I��ȟv��b�N.�
+�$�v�P����[%V٠���O���w+Y�E�d���O��D�OR�i�O�蒱�V���s�
� u(����
�){���(տ7�2�{Qe��fj�'H�O�Q�HɉE�ly��_�E�0��5fR;�f��)чv.mZ5�O|�����'e0� ���Vؼp����8-�^���O�u��'hr�I�<��ǔ�d�@,��=$�1�+�T�<��ɻ-�؈$�%u��hAmYԟ@ ��4���D�<&�vU�I0!�A%N�ܹ��I	#`�5A�-�j=�1��?��PT��O���a>̀��Y2lQ�"��w���R�De��� H��i�m$��ٰ<��^o}����9��tp6(W�J1����.��Y_�
Î T�ay��]��?!�m�FnD�S�ԗv�&�q�c��?�����'��>���*�r�a:]��x����z�<��eٸf��4�"C4F��q�My"�uӢ�d�<��FY����ӟ4�'غh��Q/P
6�p��9���>@"���ڟ\��.�RLzǄ�0c*�-`c��$XV�c���%�T��d]���Ҩ6"z�	&tǶ-{1��[4��C�B��J_w @ q���7�pu���J�B`���� 	��'@1�r���	�y��d�j
pi��_����I�L����O�f�v���#TV���d�\yr��)4����ɐ�9j�䁂��D�O`���O��?��'�� �$Ll�x����&�2��hO"4���0AnA!��7Z�j��d \��'#��ұ�t�Ӕz���ɦA��>���摟 ��'��I���<Ѱ���Ϛ��q�S�|�Yp(�w�p@ �Op�OP0cR�>!Ԙ���?>D �#ALI�zt(DPRC�%լ�O���h��d:����p�ۢu�mq�ǉ$eê��c�>�r�>�+r��R}�dgQ�dې,޾s�7�
�?�@��I����8��?qp�ߴ	��!�K��NR�I�MH�P� A4}�&}������	�M�vj\�������6��Y��cPSy�Gٞ��	��ȟt�!� ���x�a�=0<��$Fd?u��g�T>片w?�����x!Aظ��`��{i��'*��-�I?z��ʉ���Oa��	+� Vw���M@�R�U��q�$��'i�S��'<�ȣ�'+x�	��q�����ژR6���"�������G+�H���/zh���.B!�$�7&1�)�<p9!��PV�v�'��'�(�g~P>7�����1Z�CO ���%.��?��	[�]����S�*Zr��0ꄊ�����!�䈍RXU9R�c���EA�2:�!�G&`������M��J���*+�!�ʅ2�f�Y�K��`�r�=�!�$��ܬS�!�W�C�D�/!�d��֬%����q߸Xh'N�"5$!�۶h1V�yцh��P���>#!�䛕^�Y�e�_ 3���`�-ҏo8!�Dɹ62�B�ˆ;C���C�!�Ć�X�zd��gĮuW$���L�A�!�d��I�2�ChĵV�I��)�!�dß;"�P��K� h�%#�B$n�!�H'a&��SfP�?��]�f!�� ��O.,�Q��F�d�M#yo��#Dl���i1 ��20�(Q���͟5d:M��MD��c������'�!�����$�������ʭqJK#� 9"!�S������9l&�%��ʁZT@J0�4상�P�7(�(���4|qN|��hL�%��&�(Ӗ��x�^�K�a��j��eB�4D���'�N=pg|1Ҳ��	����4D� �m:N��ۗL&K�IJuA0D�̈¢���
C"ٕ���`��.D� ��;�t)a��Vz�3�:D��Qr`�z�4��"��Ĉ��8D��:�BX�J��N�!}*��G�8D��(E�Uw^ 
pjޫ4HX���6D���BᘞQ?ƌ0�F׀@���e+4D�Hk�!
�A���b��i%��i3D�`(`W#m��s���T18�S,>D��AT�s�t �D 	!2pC�.D��B�̀�- p�a3��W'Y�L�!�� �ԂsG�4TR�|��ۀS=D��"OT�6�]M���1�Z�q$$qa�"OF<���ӃVq�ݒ��6.j��"Oȑq��=����,#?>�A�"O���#��(8�ıZ�����\z�"O΀�4��+l�X��OŜ�nȰS"O���ff�!*"(V	o��p�"O�ӒOUD�~��`�,Τͩ3"O�5�d���R�@��+���"O<er���
�J1PҀ�C���"O����Ψ	�y����~��g"O^�+��Q<y�����G�<;d"O��#��{��QQ�"08����"O~�"�nC������u+�Ȁ�"O��h�*��A�^�k櫆�>��I�"O���w��;��#'
J�Ij�a;U"OV �wJZ�[�*=a��S�<_�AJ�"ODM�Q��,��J
4Ȝ�"O�M�&	(t���!�J��B�"O:ez�A	�&}��B��C�Su"O�=;a�޷}z�y��L�>�aC"O�M��dȠh�j���^�se:���"O�D��oϠw��� �,��r"O�<AG�T�*c"����ؓ
�f�g"OF���Ff"d�a`.�	S~ʵ[b"O���#J�xO%q�
�yhx��d"O��5ܜ�x�B�C+xh�0"OT ��莎`�,a��i.���"O�S�K�,C6L����O�m`�,sE"OJq)�@�>B!Ι
���-tm�ݹ@"O6T�#�N�Jڲ��RL	yv"O���J�?� �$F�%<<���"OR 	Q+�B���E�>\�z�"O~�DQ�i��,���K	8R�Q�"O.�9��ko�x �@]��!S"OF�0S#߲x���{���:鰅��"O&����T1ZŢ�YFŗ"�P�Z�"O I�A�=4���e�^��a�"O-���c�ʔҲf˥cI�u"O�-��h��4���&��}4���"O�5 ��δ89t�K�o�R���A"O�	 �#.�r�smɇ1>��&*O�}�T�ܻoL��Ri9n��S�'3�%�c���$l"�Ӻ4[�D��'�tt*T��+I�B4�0`�B7D�|�S+R���Ŝ��$RG�5D��ó�B�@�V D�%dVt[ע2D��Z�ɶ>e��B����*Ъć%D�����ʊɤ����=P-�=�Ɗ=D�({e��"0�OZ�@I�ݫg�8D����
�!R�X�J׉
n���$�3D�4rCB$+uИ��LU;/��$Pl2D� K���0�iA)�,>�����1D�2�V;�*-cQd�
�<�)1f0D��c���=j~e�Bw}l��蟞�yr��_:z�{ �M]4<8ê���yR��2�٠u��B��p@�-���y���%�Ɖֵ2�p���6�yB�'^�d	�fI�1Lj�X�M�y�凵#sV�#�hA#+KFѨGh���y�m݈UvV��J[V2�`�M��y� QL�l۲�Дz�v��"	���y�I� j��5�%�J`h�)�-V��y�ɟu���P'N�U�̐���]��y
� j$y4��r�(�i�T% a"OaI�o�5gT�7�8t#Ҽ�D"O�:���_����0	E�>��2"OdpZB�:���c�(סD�@"O$�٧k
���a� "�m{s"O�U���C�=� �B��ۗ����"OT �ԍSE�F1�P�{0ؒ�"O�;�
C����RՀ"
��)�"Oh��ц́=!Zy��@���
AA3"O�D�q�
s�u��/�(g�X0y6"O��Is���D.A�a����"O�	8u^�]A;�,NW�> `"ON��Ɇ�F���V,�6���(�"O(yQ�-@�dY(4RǫB�0����"O0�Y#�P�,T����Z��ޤ�H�<1��҆rے0���3<�1��,N|�<�$��� ��C�č
e����NC�<Y4�џq��5+2���/��S��Vj�<�4� ��0/�?dg�a�"��d�<���)��K��g��Д+`�<�jU3J�b<1��ɱ8渹��C[�<�����.��=)Ea�8ke%���Q_�<ypc��Z-$�"��ĞI��icŇ�Z�<��͈[ڂ "jЛ7]� �m@[�<I'��	�xG�H�t��$@��GT�<�p�]Xs�U�ǡ>I��}�V��v�<��T1��)�d�:;�9ks	�I�<QQ`օ.y�0�� V�j��7ͅJ�<��$�>	��c�lG�,��2P�l�<��3'�T` �@E7�����,�]�<��/4?0�1CW ۄM.�b
�\�<���_1X�j��[�&A��� Gs�<��ӫ!��'K�r���r�n�<��B�9U�$iW��k�d3��i�<wAQ{	��BL�������b�<Y��_5E��pAR�^��##�\�<iC-�D�<+B��-$�!L
W�<��kF�Fx�`��b�0�<�˰�Yh�<I���?�M $f��$J#�a�<�/��qx6�[�#��v���9uO�_�<�4�Zs_v�Y�(W�Dg��'
P]�<�sHQ���v�x��_�<sL]<��%�3F�č��a]�<�4t��vɛ;Di"�;�ADW�<	Q�K7Ͳ�e�40��2S.�x�<ic �kj2,
RH�� #"��3�L�<���'S�^�iA��* 〉�D"N�<!�N�r��h	){�pA�Q�AG�<D�ҳ	�֘z"C�;/�x�ƌZ@�<Y#�:O4hA��݆O�u����<Q�!�)@D>��5S��B���
S�<ѳn��_�@E{p%_9r��-�Hg�<�M�� % a6aɩ2XT�Y��~�<�ǁ�=g� s%�p�f���}�<�v��1�M�6dR�8����&	|�<���C�z��Y���>Ⱦ�Y�z�<��O2!�0p �D�0*��|�A�L�<�2	Э7cb��Q+�0L	8�0�h�G�<#�A�^N�9fd��HC�bOJ�<�ւ�2i��
Q��G(���Ԩ�H�<dm�3n	��'��RnJxX� �B�<��%#̠��uCԝ6��/aeFB��5/�]A#"��d�<C�(6f�^C�*8$"X�f�Q
s����,X�6C�)� (l	�Uqʦ�K�%_�1	�A"O�塢���9n��1��(��K�"O�Ȋ�g�7I�̡�×N��pڄ"Ov0*�ˏ1|���7��F�����"O� BK)5Lt�J�]�y"OV�2ĉ�]-u	��*'N`�%"Ol)CeE��D+1�'4=.�j"O|ha ��_�V�3]��ۢ�Њ?!�dϭ%e�0�*��:��aܬ}!�$=Pڊ�3iD7!ܰ*`�W�k�!�$�%��	�F��I�ިx�dD&o!�dPhݰɸ�#� =�Ȅ��$!�D��hq�K��y���e�!�$1,���*S���t���¦�B3h�!�;kr����X(^��k��U��!���
W^��[`·�`\�2r"��!�DC���X��G�Y�P�`�`�!��/u4EY߈Omn��S�7ZC�	��,l��*�����5m�Au`B�7��l��U<EZ���d�YbB�	�N-�����:c��HÂK[7)`B��Q���1��	:�ȓW)�c>NB䉝�޹h�d�7}�p��R��^��C�	<p�:�)�(�@�j +Ցlu�B�ɻ0|��g�ѭ,	(�!�aN:k�
C�ɏd���0�Єe���9qB�A��B�	3^�
��F�Y�{�{�L���B�I8{�� t�W'h�����A Al~B�5}�T��ɝJ2�J� ��-,`B�	.g'�1��cJ�j1�TK4�?V\nB�	f�v�1��ވK����SeA��TB�I9q�8�e�!h�lp��oDn<B�8�Y�E�G-�h,��i�5�B�I�r�U��m��e�u�O��C��?WѴ���=0���h���;Yn^C�#;��b/�?8�Q�Q�^�I|C�ɡ@�����4fUЁ�rVC�	>:��0;�j��G�"����;�C�I�VnjT��%ΏQ�P�+q,L �C䉹 ��I�Y�)�$�ۓA��d��B�ɂO͐xk��s
�Q;�*Jk�B�ɧ�Ψ�So�:"�`�� ��B䉿�r���=:��́we5�B�Ia�j� ����t���H!+�
��B�ɀq��Ȑ�'�'ʜ���FS�B�)Nl<sE����@%j�X��B�ɮ,�8LzsF�O�\�)E/��B�I8(�")���:u�.!a�0&|B�I;3w~�  Ȑ�=0�کiKzB�	)���2��4(%ܸ��G�B\tB�I%Y��R���V/�U81��kcB�I:8�H8c��/�����˂�mc�B�ɫ]�L�9U�F�8Ĵȡ�
�Gq�B�)|��WǊ��B4�0�V")��B䉅$�p1rK�����d��/&JB�	X�l��iW� 
�J�	�B�IEJ�=�U��'FL�� �$�"$EV�u�B(S��I�2����0���\N�ZQoB�v�D82�B�/4d!� �8LRp'�]?R�ʔސ1D!򤘂M�bL�� U�]h0;@��>`�!�/[oDH�b�<O~9��a�=�!�D�_�X �q�]M�bA!��`�!��J$kr
���	�&�r�&�G��!�$�E�
�	�cѢq�$D����c�!�� PL*GY�(h����ɖnu��`6"O�!���&�h��R�XU���"Ot�f-��~=�4��.Tm+X�@�"Oh�aTB
J�����8$��4"O�p�˫hh�`� �֯)-�i�"O�ZUAw�ڼYS�,(|�"�"O4[��QqsD��؂>w� �"O8h6G�?d��(���mj�i��"O:�{�AP2NHbL���F0fPBHrs"O�(�S�J���a�� '��+�"O<�3���?c��,#��"Nih���"O����dɺ<�8�H�LZ�=�%"OZ��AU�N�ll�HJ�zH0��"O�!�R$B!B:� �3�����E"O�̰2�A�w��X 
W �d�+%"O�P�G��Y9�i�2�Z}"O�с�/�?��3�n�q*��B�"O6�X�kZ�n3�Y�����z&����"O4`[wD<C�D}��m�&K�y�1"O ��։�.{���gG��t%8"O�M�ckN�9Xv)��%D'6e�M��"Or�[�O߻NÒ��5EV�3ü ��"O� ��IU4nQ)���X7��u"Ot���_rU�yBd�^�&�(�p"O�(#�U 63�$���	,x.�o.D��@�fN�#�r���y��*v	:D� !�c, l��%,�2C�Ь�f5D����M�cCt9ç'u��*�>D��e杉
��!��ݨ4�R�!D�D`���C[�`�7�O^ʵ뤇2D������o�tx�lDo���x&D��sS.�?@
9կOe)�dE/D�4��i�s3ʐ����=���4�+D����B� ��D�ƻ~[i"+D����j�D{�ȟ7}�$k��*D����R�/,�R�(ޓK����H)D��ɷ��7|f�Ia���[+D�$)T�5Ri�u�ņ��}�f5� -3D�����"w�(�`0�G� �����A?D��j3����,��*�#)��Dr#�=D��9"�4k�<�Y��IY�p�A:D�$��߽-��0[O�%R_l��6D������P�Z�1r��#{4�w(8D�̒�(K�WK� D�ڡa��9ħ%D��@ �G;�՘�
Y'ь! ($D��J悃l2Phu(��|�R��%�-D�p)ǅ��`1��a�L��4�RPA)D�0�$F|��NӀ8t`:D�(D�pf�,k�tT�Ф!z 0�D�(D�@q� %*a�I�q�&��0���:D��3� ��?������^�I2�P+e=D��q@%�H�\��G܈Qä���:D���ݜ:-����^=�����$�y�$�3�r� An�n����Be
��y�c�'lu
�;�E��p�N`�RMӘ�y��^�T��uP�A�'h����u+�y2c�=�� (��_/uL�Z����y�L4`LI��ř-ZdrdO��y���3��`���:�bm�Wg�o�<�1+�>z��RrI4,�^����J�<���e�L��LY,h�K1BN}�<yBeec��� Kh�ň��X$�y�� 5�CHO�D�<h��c��y��РRtp��@�>{r��2i]=�y
� 5XGB$v�4�:@�O�OF�=&"O8
eL�.:�������p���!"O 8+e
�WDҝ­�!�J�ʲ"OΥ� ���#R<躓���4�
�3"OPm{���t%B��囹C����"O� �$�ڤ:;�5�.�J@V"O�52Pj��@Xj�'P!�D܀V"O@(q�f���0�ݠ8���g"On(8���)>�X8	2얙l�"��"Of�Q��$⚱x0#�p��P�"O��9�h	<Khx*�a�&G� �k�"O2!��;|�(�0�ֻF��ɰ"O��z�F�6.�����2��lk�"O��Ǝ	 m�|XT���A���V"OB���Ha����L]Cq���"OL(�Ȟ�U`��"邔g�(h%"O\z�@45!֕��#:�j�Q�"O`�@��1�yC���O3̱�"O��	,I=��Rs��0'�A"O�,"SoO�sC�\���*Ƅ��"Ol��CE\8��=*ѩd�D�z�E2D��k�9^b^:@�
6,
y��`>D�h�'N�;i��M�7 �<yR�A�?D��aɌ@*��6�I�S\"� 2
8D��@q��'>3tP!U�Q�`!����L�<���\�V�DYJ�b̰<F�:A��@�<�����L����0j,��q�Y�<���_�E��!��w&���@��M�<!"Z�Bf��af�0
V	xEI�q�<��E !;uJ� �垉���iǬ�r�<�QR�5̸Ro�ǆ\	�-�O�<ץ�'JB�*F7Np-�tHN�<�kE�%��YPpꏰ@�T���G�<a���#���5��	<��P-H{�<Q�)Q: �i�f���Б��g�R�<���5�
�8'�Z^K ��3�VH�<Q��N�\��� b-��%>��3�G�<y�G���-IG�P�#�hdS���i�<�IW8Ҥl۲�UIɈu#Ai�<���
X���PoN�mcx �n�<I�e0 �{�*��j�42�LE�<�S�V���ԢcA. � %"fƗ_�<� ���J�D`[A�8� ZӁ�D�<)��D�w�pɣ��]
d�!��@�<� ����Z��s�ę2u�a�<��S�S�H�12�Y�D/V"b�E�<Y�mܚ~�<���H�Tcv�+2)^�<�p��egR�C�I��� ��\�<�G��'|��T��<H}�ɻ���o�<���H�b\���'�Y kd�+U�f�<�FjT	~�h%���>#`5����~�<)�o�3z6j"�B��S�b�p`B�z�<	"烀5�X���Q�L���'��u�<��%ī(��ѡǷQ��):7�Vp�<�25r���Ve³g<8�K�<9gG�f��`��(��>	��E&Gp�<	����͊b��kD��Y�
�Q�<9 �<A}�qh�a�d��qGH�<�f��,yr�0�f�Uy���n�<� $�'�����ϼ{@��"�g�<)����x��gR�4"�4�K�<�1(�~�htjB�"�:!����J�<��F��5��
�x s��TH�<���^�S�q��1`�ebMH�<� C�K��m?�1��C�z�|��"O��xuG�1B���7H�#r��ؖ"O���ŏ�X`8 2�':���8"O��+�.QށF-R�X�p8�"O�p�@��->=��Ð�gV�t��"Oha$lT3��iY1�K�B@���"O�x2�V��������u�"Oh$�f�Y��4h
��]�&����"O,X��X4h��]�EB݄}�ʨ�c"O�Q	�`ۨm�x1��Q/-��x "ON�2AL��q��D��'P�y
"�`q"O�5i�F�/a���Y"xޔ��"O� wi
�(���;��7kor���"O�4���_-ae�M%�\ 8��"O�m���	�e� ��\���"O�H���]�����Vp�b1"Of9�CG�{���y�ܲzO�1�6"O@e�0���Y��Y�fg[��r,��"Onݸ�Jֳ�b0�D�,t�`�b"O�L��iS	Wx��㡤�!L����"Op���� beV��k��64r"O������v�=���R)����U"OB0z��<71��a�(;���7"O�E�À{;���0O��v����P"O����SN��]��L&�$<¥"O�����2\7P�p̈́-P3��S�"Ov���FW&~ߤ��C�#Ӕ��v"OZ�j�'�T���¤ǒ/7~-�"Oj��D�6窐�qğ\ūv"O�m�G*ԿR%���v =��iU"Oj��:~�n�2a ԯ^V��"O�]��
�;7�����S�-I�iۤ"O�P�lU�!I�4x�"C�̠��"O����8.�C�@H��ZUs�"O=K4iM�	�zG.�&���P�"Oxa��̓���s��k�r�q"O*�x'�`)v�v�!Zܲ���"O���j��q���5�A��H��"O��ՄK�[Р�������P"O�K@���ұcŁ�`�L�hc"O05��Ax2H13�R��0m@�"OJءqc�(�m���$��ӡ"O@�Ռ�
J��ad�/���Q�"O҉A*¦A���(��A��E��"O,�A��r(}ؐ�׋� �;�"O�91�߹4!4yK�b�*:Y�=��"O�q3Δ"�ʑ`f�����;r"O�=RSIΕRB#�CR��Lir"Od��l�Y�3�hU�]Ĵ�+t"O,�i���Uw�s`�Ȓ/�l�"O�M�6���S�L��󋅪|��	0"O�M�F)z!�M̓D�:�qT!�2d�!��ν.�(����ڟ2��I+4A϶]�!�ܶ2y�Ǐ�iZ9S�B�;�!�d?c��	�q��9:�6 ����&�!�˞)�d� ��G�4r(-`E{+!�D@�G��(��	�L����]�!���C�$L�a,öbM�(�a�BT�!�)��`B��O��M!0�̥`!�DY�k�"تǎ�r��)Xj�F�!�D��:&�:E��5�r'�>�qO����
@r��1��9r��S�|�hݲ1����i�7�"8x ����y��	̩�	�2px��L;�y"�g��1��Z2#���;��R5�y
� �bS�jXĐ�#�׹�(@!"O��)�@�9?"!ZB�ӭ!�l�!"O���Db8
���ѫ��ͤ�"OP��w�F�VX4��C�O�!Tj�8�"O,:��<$����		_^�0�"O�\;�J["`�>]�6
vJ�}:v"O�$B��-:� 	��O�Y�@�ys"ORUPH9Z,�"��"8�0"O(���Z�A�!��8Q�j��"OX��G��83��1/}6��`"O|�swƜ�>��	���!_ԍy�"Oj�qMG >�	�q-Ө}X����"OR��P��@*���
I�YF"O��ڦ��	2<2��ߚS,�2F"O��p�_v�V]�OA�N�v��"O��"UA�(g�1�����aL��Y�"OB�J�jN[�j�x��SQ�i�G"O)�t�(�l��/ڥ>L�Ыc"Oʌxଋ�t�4���.V�&L�"O*TS��țs�P���M�N8Ep"O�U��/ҡDX����!�4�RK.D�D�"H3o�݉c�^�0�\�$�9D���c΍*O񒬐��Bpp*�N,D��(�
Ų�xё��<U�,l��*0D� ��P3{�2��G�G)x�0D���ƇU�G���6`ō\���C�N,D�D�s�/2v��U��2:5�E�%D�H��bY�#n���&P>h�1��b#D�`q�űp����K�!s�(#D�tB�BC(&�5�3ę�}G~�`� D���d�����3|�d�P$=D�٠ڵO� �Ã��c*2�5.D�����,+��%;d%ϟj�QC,D�8sdă�){@�$O�8J��cS$=D�`��%S�Ej���3�X��h*;D��Qd�xY;�`I}���/#D�X��ߎ;ͨѤ�J�iߢ�"S�?D������&��˄�2JԵ���)D�X0e�C�2F�0�8-E^���N5D���afߨAP|x B�4k�dujF	(D�@0@�V(E혠�V�V/=����!%T�d�WȞ,β]aj�;<攱C"O��XdAӸf���;ↂ��T��e"O��
�=�Mib�ؙ<��A U"O�Ը.�		YVeȻeQn�z�"O�1���	P�6|9r�{=� �'"OH����2e�&����.%��W"O-�6%]���D�Y$B<�Y@$��X�<9�D[���ׯ�#?~q �n�V�<ɦ�A�ΐ �iC�_>�pd�w�<�t�/8�da�"&JD�>��Ƭ�s�<�sC�>SVa��ț^גI����U�<���>]>�ӑ��azT�UD�N�<9�NAu�BIy�.ӕD�0�d�K�<�hɂVx&p� ��K��+��O�<iR Uyd�С
� �f��P�L�<��ъ�D�1 �<�R=���F�<�v����ɗ�ߍiv��w �@�<��AO�sh|��� w�p\�ƦYb�<qV�`M�d� ���>S"ng�<)Vfʁ0p!C�D�Gq��2�l^�<!���:LG�xeGA�o;ڼ��ƎX�<�R������u���r������kM����KӚ �Ti`���;H��=��S�? jX�e�f��H�`�Fr�K�"O:�J'�z�-*e�L5s0<��"Or�˖ ��vT`�9 ��:$:4(:�"O�z1e�(cȰ8�� �*?��"O.Y��F�Z�\��һ%v���"O�u#�"]$rxd0	N�U<(��"O�	�dmM.~4��:\hT�r"O�hB��D5��	 F�|
Z���'���r@L�`L꼐�F�Oa��'����L�\��D#L�l��	�'�p:D�[���j�*��1)���	�'a`i�c͍�Ed@$;�e��~ۜ���'Q��ٶn� j�@�-�z�ܸ�'̰(��FA�k�8D�䊈�s�i��'L�0�f��g�J(p�'��:����'����W��J��+�@ 0z�4�
�'�, ����X^�9�P�č#lq9
�'�h�b�
�D��((㉜"�t��'��mr�C�y�6U�f��=0y ��'BΉ��@+ux6�*&뇯�6IK�'�F�ekS9?wĭ��H[�aSl���'�Tm!s�W�Y'vmPF�>U�M!�'Dq)��2Y�\�%�H�LLd���'ٴ��W�S��0��+�71/��Q�'�X(��f �r�#W�˒(�V��'�Z���.I P>�(dX=!�ЕB
�'�p���/	�d.6���ӟc���	�'�b��U��"���/ܾ#��t9	�'VDrǂ��6���Y��sȘ�r�'�P�	"��|)4ِ$�=��]�'�� ����1*�t��c ������'��ĎݖM�lĪ'L$u2��q�'BrĈ�-A)hfy�#���3�'�X�Q�+K��C�J_�j��'Ȣ����HS2I�陒R�Е��'z���}d&�R��	b�0 ��'���7`ՠeǼ��g�9*�ظ��'��p �C�k�*���Q5 $B�'�2Ũ� F�=�(��elCk��Y	�'<�-ɦ~�Phu�M�z�~ur�'�b�@��) x�<�3�ǎgF���'�`��M���q��_��a��'�R���瑜\Q���)M�dm�D�'�4��|�t�XB�����.O�!�B.Q�F�a�+ߏ]C�uY��Tm!�$W���(`�F��3�.�RC	�!��ӻ>����W G�A���	B�bt!��M�@�㠀B9֬I�N,a!�$�Vef���D��M�d+n��B�ɚ�H,��@#�2����G�i�`B�I�GX���Q^
K@�ƻd:^B�ImV�`t4r��E#
(B䉢L�>��r�Y�JBB�B���)ݰB�ɏ'��I�H�v�ĉ��LW&��B䉩k���ˆn�%�1��픪QF�B�X�&,
х��so�Z�R?�B�	�k �� ΐ>��у��T)aN�C�N�jq% 1q�v :�'��P�C�I�b$���S�r�R���"~H�C�	_�%��,Y>ej�� 4鉮	���)ړ�v��w-S�����G��޽��k3`(�ᇀj�r�q���� L�ȓ^���l� B4�Q�D�U��lvXC���,h�T�c��LɆ�S�? 84(��Wv�l`�#��1�I�"ORQ��.�w>����T�"Op��Q�b���8�^s�6ls�"O��R�/ŧ-˒��/X;D�6���"O���*�nh�h"�G�{`���"OTT#1�YT��,
� L��"O&m" �i�)����_�
؊�"Ob�2�C�X� '�;D9T��"On5Z1��#M^���MFnJ�!�"Odm�e�O 7����4��3&1�"O�9���r)TC���<c���#&"O����f�;,,"�D+?v��!4"OLu���֯>�8Q �T*����"O����H�K�D�7_��js��`�<���N=O�x4eT�B��Q�TG`�<	�bYC�����	��%'�b2�X�<��Ɏ�g�j0 G�Y�#5�8q5� T��x��U$Xb�  a�do�ᢂ�(D���DXU�i�èՠab��+(D�,�uf�
o��@�ҽ(��es�
(D�h�2/�T_0�ui�9Cy�M�q�9D�0�#斲��Q�MJX\1�D�"D�x�'x��i�A��3,�(��"D���s�p��P���TE�\�!�5D���'ϊ$�
�$�k1��8q�4D�䒁�u���HE��mhZ<�C�6D���7��$��Z$h	9n?�Y"s�9D�ZgL��T�� �-����}���5D��zc���1lZ0�dA47�ba2D�4BѬ�%INJ�I�e]�q�L���1D�Hb�j�(*e�d%�"g,a1D���!j�&*dD��j�T.��pF0D���c���%E>��1!����E�dB/D���Iɢ1��F�	�<}"�D�!D���T+��e����Eۗ_�ͺ D�|p%١M�JpY�3�N���#9D����C�5<-is��Ԉ�Ä2D�0�W[ 9#�9����c0D�x�e�#~�!�	��W$�� $#D� ���?�^��FŔ��br�<D��V�&Oʥ`�lP���<D�����W	��B`�nY)rG;D�`Bp�M+JN��§Ĝ�L��)Ua:D�x��)��43�5�c�� h 9��(+D�	�㑺�v�Qun_%1�&XCGk4D��CR<�1��>����1D��7M��_���v��7���k��<D��r��ݯ<cL��!ZbI�3�;D�����_�U=<����Ҕ'�|<�f>D���c`مY$�r����-Jhb�k'D��{��
cZL	rcLZ�#�PK�&D��Ư,�LU����(B��!k��*D��@oT'6`�������w�%ᓠ'D���@ߏ.@��4Km�f��&D�L�u��7p%@]âI��D7�Ҥ�.D��r�ND3w=6p�L<g���Va,D��N-C�2X�A2N��EK��)D��@���/���%�9[�\���3D�\��C���p`��ilVx�0�6D����ʬv4z�A�$�(8	8��6D��S7"�/8߾�K�ϲT�`��Um4D���2aX�@I��/�U�$lj�.3D��� q/ �8�
��AI��i�+3D��5
�"##>��@�
=��U�6�>D�� ��X���GL�{g�P4�TxI"OhABC!ʬ4�0+6I�%�X�9E"O�����sR,I���Q�S��\�"O�X���NJ�ԡ�H܂]�P��"O���hӹ'ٜ��&^��P�R"O�([�J��hY�ާ2�HRC"O�13�ݑ$w�ܺ�%O�cz���"O�l���Рis<Tcu��1.���"O�,js�Blr��c��
[ifd��"O�-Y��#'("�b�E[��N�a"O�q�� �7ufp�$��>dQUi&"O�$��c�l�r�Ň�J+�ɸ"OʰJP���0r�Z�$��D"O^8(h8(�H-�d
y����"O�s�N�L���0L�oF��Ф"OX85'%����*F�h��"O�{�'A�T�a)� d���"O�y�Q)[3;dIS��-xr�`�"O�E��DK��2m��I�I\�в"OD��*E)<���B�$�]7�!�"O�T�SD u��)Kp���A4x�#�"O���f��A�!
Y��u"O����c��+��(H6˃A�6���"OD�Q 
�.A�b��%c��P�"O
1y$F؅TY֘栆a���%"O�P����J*�Q�5>�8���"O��#f\튣'��"�D<�NC�<�옆3����G�$
��)eNW�<Q�,��5�t �"H�h	%�R�<�&�]�)Ef����w�6���@V�<��-�s���¤��L���r���O�<�Q�;"��0����=��$��R�<�����YF��E/	_9�13��d�<��␁�.E�i�	�2��4AY�<�ߋ{���`0�c�a�cNK�<����
���+u��Jt�}��'�B�<��CO)SU�y�'?�襹���@�<y2��>��hd��<H!\����}�<���]�]j�iJ���[�:���HR�<�BR�8�
t���n[L����U�<�!�?p�QXDCx�ХQ�<9R@M�v=r	r��#IrT�DKMJ�<�d�:%a�1 sH�:��-����D�<��lH$nejl���-�j S���}�<q�Gӓ]��A��eߊw;�+��OR�<y�ş{�x�Ǡσ@����Ys�<Y�Ø,��XS@�� t`�-�$
{�<108��TJ�ۤc'F�ÒM�u�<9&ƅ��x�$gZ�a]� �Bu�<�a�d��'T�"�����u�<�qi��G���S�Y�9�<x���Y�<qv�L%d��;"���P)�f�S�<Y6�D p[0�Z�s_� 5)�C�<�Ħ#3�n]�֫C�[��0�΋~�<)$jՅkRdr3��� ����2`�A�<!qI ��R�����(c����i�<y� �S� �X��*,��1�o�a�<�n���=�0�$jbh)�Pa�<��[;U��YY1 l��MIE�<��[7u������:<��A	6��F�<�æ4JS*MK1Hĳ�lԸ��IC�<a�/�Z�
P�S@�V�4�H�JQA�<A'D�
`��h{�i0Wy�&g�z�<�Z�C ����a�)C�YX L_�<� <șԂM&@����!�	�E���3"O�ͩ��+w/脒2��V�pYC"OtU0��rg2h4�^*�eX4"O�-hQ��u�l���ՐY�-�@"O��#b��j�^�B�-Пn���A�"OT8#��s��ZM��n���`"O�����7����+��lv:TC"O6Pb� ��F�jأ K�`,�R "OȤ{��h �(�$Ɉc'�0��"O�y℄�3Vb�����<���F"O�uX�-X?<�e:D��4����"O�v�϶;��,���]&�<�RG"Opi��fYNR��;��ҥ%�\t20"O�,	�cD�Pr
C�g�J�ف"O���&�-{�j�\6u�h��"O�(�S��!(�J��)�t� 6"O�0�E
@����C;�R,q�"O�\I�Ė}��8��X�"��f"OP�!S��{�X�����dS2"O�j�l�Fn �"���[o���s"O���Ű�$-�e U��Ad�u�"One�b�Rc�b}	 �ܖ*R|��T"O��#$��2�50ÅG� +Zݳ�"O��xT��$s�T��@$�6-h\ȵ"O(Q��j3�+��^
��d"O�h���^!��A6�<�F���"O�����84�PbT\T��4�"OD�ri*mc��i���p�
"O�X�ΛsR��p,�&Lf�}�Q"O�X/ݷlӊL�a)I+l�`)�"OR()��P<Hi~a���;�
Lҳ"O,���K�+��I�DZ�>ɒ���"ONPR��"	�
�h@l���B���"O(��c#�;Q#�XQ2��~�v�`�"O��a��$
�B��� ?�A�"O��$Oa���SiN� $ڡ�4"O$�"%i�����F�?�-�#"O���G!R4j�!��4�T���"OB� 2�F1�811��IC�"OK�����H!*������Ȩ�y�L��7&F=3 ��4-�Փ`Iډ�yb�$)U����G�	��#����y�(JBI&��-��jn�2�̈��y"!�)�di�I2s�5���yrIȨƜ���F

&j�p���yR �L�������"}�(e���yb ��+���/��FD `� ��y"g�{�X����1*#����y�䌀X��a+sF5`����!�y"`ԶH����ك,8� 2� �y⪈�m<D�r�GG�?B2�+�%Ϋ�yb�B8g�Z�;Сǘ:��!m@��yB�ƐZ\8TЃ��4V.�p$��yb�?{�4Q��F�0��ѹ����y"iV�	&��Uo�9t�LH�#bC<�yR�4lO.��c���mߊ��h��y"K,�|�PiލRJ�,�	���yb�A
[���� _L�(�2���y�GW��d!���.~�Hg��y�KUb��L�B�ԏH���Ԡ�yB�X��P=���KX�pc$n"�yŭ}f��c�CV�8�b�'�yRŊ%���7&W<q��x��jZ��yR��&�(��W�dz��CL�4�y
� pQ!P(�Y�$%Z�l�"O*�zF@S�"��炚?9w��!"O蝛�� x�HdPV!	/��� D"O���)H��
$"���@l�رu"O �z�� f����({]��@"O��A�T���⠓�0O��b6"O���Ç�z����W�R�10*G"O��r���s@�R��u���"O�y�#�V	o�XIX�E�2=����G"O0��C!�ws�p��V'l�c2"O�)i3i��!kȂ¡�q��LP"OFWJG��ڸ�+�) ʊ��"O:@ O�5Wh���H�V��i��"O��ӀK�p�0�ԻqAZU"O���`�7�°��ؚ.�F(9�"OFY��,X ���e�-��À"Oh�pӠ�Dm�aب���IR"O����B6W>���%�u�vP;%"O II�$G4f8<	Z��S.aܤ;e"OJM���ބ<���wĆlX�s�"O��(F�U�=�0a��c�-R_4�#g"O�`�l
�u:Y[�(�")>�� �"O���E��2� �AW�O���"Ov`��l�!m��=��!^J����"OH%c��ґE5�9B��P1?�.�xT"O�`�@Ԛ"(��Z��6j��5h"O�	�Vd�)#W��9"�ӑJ��y�"O�сv�DCҌ�U.�<�E�5"OZ�آ��D��­�Cx36"OZ�X��G97�d��6͑'�9Z5"O<Y���;es&E��	�(�ZA��"O�ؕ���M���ËR�5���%D��w�.@D5@O�pu�i9��!D���"鄈G𩻶A��:�p���3D�,j �N=X�J���<IL�d�dl.D���GR&��\��7km>�V�0D�,��-O"f��d
�4k� �E-D��Q!� �uw������X�cF,D�Hѕ�o�R��������n+D���G������bUH{%�6(_��yҧO47�� B�"G�w���⠃ؖ�y҅�z�:����9XN��a�=�y2��)���p*ƬG���#��[��yr��>�D}�oJE�h);��R��y�%U)F=����N�F:������y"G�U�&�Z��̑=�
��Bٖ�y���D@�ѣ22���bl_�y��QA3|�r���-�n��G
9�y�ȞH����*,���9E�Ǐ�y�ڡg ��
�Ň�(d��C�yb�Ku�m`�� z	Qt�S��yb��q� �Ȟ���L�Cb���y���n�4`eN���5�_��y�選w��{th�}!�,�5@Ʒ�y�g��&�����#L��$����y��p���c��)B	<��dž�y��z���c	�9�2����5�y2�ۨI���au�*��Ha��yBbȫj�P�"Ą�8���Hq��y2 �����f �>GV � ���y�B�09����G;#�ؤYS˒��y�lVL�⸳���!*X����@��y�ˇ= 1eh����.�%�d�ʛ�y�_��j�c����!�BA�y
� �L颮�<���;��ÜN���c"O|i���j���s#2S�pt��"O�����+�J4slƦQ{�a�E"O~�ZՄb^�mS#�&_L �b�"OL�n؏2�t�0�A�A<��b#��ҟ���d2m���)I�2�ܘ�S�@�86-�`�aqO�dB�9+V ��$��ZV �i�Ν�[���Op&�زؽ*b�I�f�Ôi��]���%	��c�Z���آV焪P��m�'-���!��X-�]y4*ɵhT��Fz�m���?���Q՛&�'\�e�<у�@��`B�ܣ����q9������I8�	<&�����8-���!���>����dKǦ�`�4�MS#
�\��T��
<"Ւx�E]?�	�X�F�'+�i>=����!A�� �&IE�eKbo�>��1 �M |s�УW&���� j^�/q�J��w���ð��A�[#L(H�6B�⦭��fH2���j�Os��������H�k��������˕�n�)��Ħꛆb��?q�e���'�?7�� q���W)�#m̱�����J�$�O<��5�S�S&g�Pp�#����� �hxv�<q�i���ig��]�-(5�`�V�����F;�LʓyTFX�c�i2ayb!$TD�&�ج��ӈ���H#0��y�b�nڴZ�+�D���Z�I7�/��H�	O5U�E`���<i�X1���ԋn��T(��f��D��h��c/��ZP��Z8�ze��%�v)LM��J���t������8�ɬk���<q����Ĉ~����f��-��ʴ@F�%�$$��bV�� �:Y��_�!h�		6)n��6R��$�p�O��	�7�9��f�&g�� p!,(��d�/$��M��ԟ��I⟐�Re��x���`r�D0/ud�[��U��zW�ـ:ԑ۔�Ǽ>k�xXvm�;D�p�AB�I�eS:p�g�*Z����W���@�6�I�@�B��r�L�5N��tO��">!D��Hn��F��$��gĬY�,\Y����K�i��[��IJy���*7
��T�N'6m���t�!�D��B�b�b�.C>Ah*0P�3��D��5ܴ���o�Bmn�$>X�d�#;=����J��<�6B �!�	ޟ$&�*\e�f�4`?qx�G^�7b�i��	�ډ��-T� � ���+� �HO�H
�%�\����e��xd.XP���|
 O�h�Zš6��GX hdnx�' �8���?���T�i���(�պ�(X;]$Y����/�?)��O����0�B51��%#P�Һ9J�A2�"�O=l�M#ڴ���2H���!� m����l?ц+ cԛ��'0RX>iSvGG؟�����鉂�l�={W�qerh�Ƙ {<T�5�ݻVI�G�ʌ�9@q�?��Oa���j<��-܇It9:!F�w-f�{a�i|lQ��7WV.,Bb(�{ZNe1�dT���k�ѻ,�!���B�Q�� �/X��E\3�?���3�6�'�?7M�.1�̨#Lɍv��wNǍ18���OF��$a�\-bm�+t��Իq�I�v��g��'�M{�����I܊[��-�3n�|S�)%�Y�Guĵ&�Ѕ��9� p   �    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   `
  
  �  "   �(  �0  7  V=  �C  �I  6P  �V  �\  c  Xi  �o  �u  !|  �   `� u�	����Zv)C�'ll\�0"Ez+⟈mZ�YL�I07)��Dw�����c]f^�aPnӗ[��9� l��t�(�iҢJ�1��ݱ��׏X<X�;t���'L0+��PD4��gŃ\�^r�e������٬8R������.^�Y[�&���hq��|I:Wj��|�D�LE��H��������N^lq���ɷg�*ٯ(�>�ش'�����?���?!��L��m����3@m� �p)eY����?I��iU�ۂX�p�I*rY�������Rk� CC�N�L�l5Q�l�;UѠ���� �'�"�'�bÌ��Mc�1OX���)��( \0�x J`
�'b��"=!���n��S��/ #���f�}�5���YX}�7O*⟴����!�':z��t�ݬ-�$@�'�Wat�1��?y��?1���?���?�(���]�>7.�8'e�$G����M��x����ʟ<n��?y�4�?��i�v7��ȦQ۴�?���+VJ�+3hȽ�*�A��]��hOD8��iT��нp#jM�~td����#�6�2�ډ7��$�Gg@X�6mW���4�b��\� �bBˉ4���� `�{�޽I ΂�G��H�i1�
�7!�[t	A���)��b±P��mp�m~��%lZ�M� K��((��e_�6����∊�gK���3��1_��Ѫ#�i{7�Ӧ ���z�h�9��E���n3#)����?�!�B�� X�3�ǀK����np��el��M+!Bϥk"��1q�RN�� Dƚ�`���JT*���J�2jp��icn�b� O7C�t���.�\2��'l�O�x�oފTdR)i����d��9O�����ğ`Z�i�&�M�͟Č�S�V�%.�ɨ��v�@I��'������	ǟ�og��R'v�xb�@�Dr
��`��s�������B�C>0Խ{�:��H�Zy>h`��]�?�GGڢ FR0���b�a"�H�� �_��'$���!�����Ϻz�>ճ��D�j��O��2�)�'Dz�,co_	8�:��vė�Ml���ɇ�?�D+ܪ{�"!9'���Q�v|S��[�l�?�1f�G�O����J�ν��$Htdj0jF��!��7��e#�+#1�D�յ�!�)2%Hd��&Fe�UƉE	!��I>)�N,�/�Bͪ�Q�i�;a�!�Ĕ�<��T���:&+RF���PE"O��ׯ8[ <�q����'}H���S?w;��ծÁf��)�#��ц���l(D/K�o�t�aV�	eV2U��O����&+M�X�����K�5^��ȓ'�^=Ȱ�FE�m���4�ȓscx,bgAӴ,e�I1��Y����Cl�a��@+���z͕�l\��'R��	�����%�8h���D�#b�J8�ȓ ��vGT�kBd{*_Q���ȓC��q��nA�Q��3W�������3�b ���x�nY��L���A��BJ^���Bp���B��)�^X�牮_���ڴ��D@�w}숃�M	B4!�Ӫtx�V�d�	̟`�	�����DB +�A��,�5h:m�u+ݦE�lH#�ė<���oӒe#�$�P���a ��
n�pb�ʯ[�v�ǥ�n\:�1����� %lrq;��K�Y0ң<�#�֟���ϟt�I�@T\Ѡh^�@���Hd�F�6h��'����g��=kt,ۼ}�>�F��Oں��D�쟄+�B�q�9⠆�eԤ�"��Of���x���i���'���`���4>�N�(U"S���P��F�Hf&��	՟D�*��9��E�%>�N�V�.?���(�'�(o�<��aL19�Gr~��?hPcr�G�_4$Hb���l
c?A[��_@X�r+�!U���:�6?)%�ԟl��k��@�'jb�P�#eA�-\,��腈q��&�P��L�����e�ڸQcVX1	�tEb��4�F��>��U�ȅf�qk@M�^4�̓����oy�L�o��d�'���'��~+�4h@I�U���C'�)�x�[�B�1��ah��s1̏c�g�,*`��IG�\�w���`�Axa K{�TYI��\f�<��_�g̓d
�h �t��S2�L$]�	d~�$Z�?y�����?I�Kly�,	eH(�V�ڴO��)�'a�I1��	�$e�J�:D�.O�MEz�O�"Z��c�O�`��}٤.�c�hZ�Ŭ@�� �4�0>1������C_Q�� �%ښ	L±��%k:p��쎶.�B�qOJ�n`�D�Bj<���79���脩u�a�@�]=_<��B<I��Y�A66���I����� d�<ɤm���u���2L�j���a�ɍ�MO>�1�ҡf�O�jPJ��?�x���ڐQ|~9���$�OD��O���S�85~�h���X�h�ҕb�t�? ���g|��b[E9�y��'��-Ҵ��'�R��.¾r.7M/U�kd���M+�K�Gax"�X��?������E,B��5a%:���4ȶ^��'�b�'�
�
�K�$q.,)bE�N�"y��� !���
�9k6M��j�Ѥ���?�+O�MӐe���'?5�O�B���8� �H��r��E�#Q�R�'�*�X��
6^5x�Zw��E��p!qiD���`CO?�A؀=F%h�+�{5�8�cm-?�⢙5Z�*@%�Ӄr�ʬ*�16)>�)(���I��ፀ�@�]�E���$�;�b�'1�>�ɥu6`Q��螡+�`4�CC(odT��j�D�z�M�T4��Jc�
'ML�DR:�'r\^uCg�F�p�@��QBN9;v�L������'��R�'��l���;9t�99уV�F��@r ���?.�@e�	#O�m$+�"!�b>�*'i9�����֜�p�ͭ,Ǫ`��5||�飌@ �
X[j�w��`���� �g��[�'9��*���˶�ũZಐ���i��6��O�)Iq
�O��I��f��O���Ox1���L9��d�Uwv%�s�.D�2eh+mM>Y3'kд8�h1�T��<���'�M����D_�b��a�ӆ�"���ա6I3�HI�J9@m2���OF���O�q�;�?i�������L��2��YY |9x �r#�r�5�9)���0�`�iĄ2��j5����&њ ��$[ ��`A�N	��Ph3IďX/��9э�S���t�U��5$�h��l��Lr�A������O|�O����O\�\���W�",YKV��th����{�<�Aˀx�@EX�!�/}LΰA�/�a�I��Mk���ė]��l�ٟ���d6�a�b)�*K��@�6GU!/���	��r��� ��ǟd"��	�gZ��U�y�x̻[��<CV��>-~�)g�ܚ
OLц�ɦ`8���FA�5��aa*�5FXY� �6<Ӯ$��#�p����'O�噦�'���|�~�D��5���x V���Q�H#Ֆ��?)��O�1O�!3���+�́󲇚(d ��w�'H�7m��tK@9@dl�E. �)g��k`-oLy�jM�3"�6-�O6�D�|�Q	�?y5(�1{Ev�Z���%��Hb��X�?��}5ȱHM�Li@��'��S{�d�=��E	���*K�)3"�ɰ����.ePZ<+B�Q�>cq�-�>!�����Ⱦ��+_�8�n8`V�/?r�埤�ɬ�M;����'��D��!O��{���[~��b�b5���?����&?���'s],9!�D�`���$��^�'a�7�[Ѧ��|j�!]�2�y�++c�dp� �՟����N��Fy��xP��렦�!� u:1lԃ�ybj  #�.�S�,íI���π�y"Ǵ$
��Q'�M>M��x�d�C*�yn9n,V9�W &O$	�����yR�5E��)�ϔ#xU�귢�)�y�T#!T�¶k��j|��I������|�C�3QG&��aT�J28<b+���yMNe�XF�?�(���C��yr.W*#O<1��O�Rj�y����y"h�e�,y�����}aԄ��[��yb,�*QV�I�'.�t�4P8jм��>��C?���D
��f*߶Y}�<�g Lb�<���"���Y��,Ѱ� �c]�<yq�)AH���p�-/��y`��\�<�����V|���]!?kt���� t�<��A;Z=\�UKÝ���z��o�<1Q��m��q��˕ �f�;U�d�'o�����˿ss�����RXK����r�!�ߗ�cA(W�C��k�\�p�!�dD��t���?"�(�ReI�q�<��l�&���� �3�d��'�h�<�U�L�=�ؙF�,-���O�}�<9��օ%��-�RYae�W�L��-p��"~��F�}�
xy� A9]���P0�yB�_�A�rIr�!%�����GB��y2�MZ�x��쎢z�J��/���y�H5o�� s�D�'s�����\��y�I%]�dj@�kj�V/J��yb��1t$�ckʽm�Ј���:��$QV�|�P<S�"�	��u�ڌ��D��y
� ��t�HXu��BM�0����"Oʅ0��B��rt�T�#!X�K"O��S�ˆ8D"`�92i�p"O�I;��T�`*.X�RB��e�b�BU�'�Y��'�B�AtGݪ�����.m��K�'<E`�L0?�H1rp��
t�'B9�"�	+��M�'�^+���'O� ��N/Cᮜ�1�$^�he��'Z"([6�->&p�!��'[O�5J
�'��EP��P:5p1���V9j��I���V��Q?��p*S�(Pʌ�� �)l�hAY�L,D�@G�vtE�`Ē�^Ϡ�� �(D�XzujQ�hag�ޤnID0�dH:D����ߧL �E�e�H ��t�R#D�JFi\������v���&�+D� ۲�W�f~�R��C t��A{��O�h���)�^��) æ�b��ԛp�ʃe��h�'3 a'n�:|�x;��(_��m)�'h��h�I�+oӺ�(UG�#S(�)�'w�|"'���Z=K$��
D*�4R�'u�h���t{L����g�Zu8	�'�~	�!G�B�X=�� K�/�l8�(O�l��'*(18�G��.���˘Q��'���jq��'?�a��ΘkT�xP�'�nq�DN?���p��i�lR�'���k�Y�V��X+ʨq�'��b��x���Y�O�d@��0K���_���ʖe�'v�
��F�xF�e���x�"��7�B���/��`�ȓC�d��2ł1_�F�b׃Jt�܆�RkfXXKK�@�̭����5Ai@��ȓ~�V�1a�κ,|n���02����0Y��*�N�&)�:�#�$��DF��F{R�)ƨ�v�a���1�)�d@|�$�[�"O
�P�!�#r��"r�F�>a,�*D"O�D�%��˶���O�LC��8�"O����=�����U0.y#0"OlS�i�(W�yb	O�|v4��"O����)�
d\Yj��ӡ��(9��'`�Z���ӧx{��S�	 ��i�!�7{L*Q�ȓuو9;b$U T7"4aN������P���8pl�'K1���荻g.�5��m*�e@��Q&"�ũ�AT��,�ȓr���*��8`�l�h�9_�^���n~*�AWm�9mP��8��6+oN�'J��	�)�B�AE�ޑg���!EC��$�P,�ȓR����b�̃
�}Q�IƮ0��L�ȓyu&t�G�Y$f�*S�)>6�Y��%��;��3e�6�3h�0b.b	��`�pT����#�IB�Z/y�(�����I����nT��áă-��ݢ"�U� �HB�	$�D��J%��`��N׹<>B�Ɇ)iR��fAɂ��,+��WH�B�ɝJ1�E P ����`��f��C��1.V�0�	�-��}�7�P9=>�B�	�C9�� F/�#ת��%�8c��=yt�q�O���C*׎g�¨�%�J=/���1�'��1阩Wb��إ��%��,(�'�X����4XqJ�B6�0[�C���y�mO^�`ܓQ��`�����c��yb*ޖ,4Bp;b��XG�љ�燭�y�D
t	0hpMWL@h1d��?�`��|����Ѝ8ӌ��T�Z\z"�4*�@��%D��qԥ��v��0�(WxD`��L#D�� F��l�B5�B�"�B��e"O�XB����~���y֡�(&�����"O�A��M��[� �Z4â:@R{d"O�0�p��=v�Rۓ1H���\�$���4�O �:��}F�1�#���N ���"OR�AْN���ba�}r��[�"O�$�t�]�af:���oâ"ͺ�ȣ"Ob���J�WF|���&����"O�в�����B��	�t	�'%�O��Q�O����M�{uRq�5��9���`"Of	�vGԧ\Ob�Da��O(�#A"O�U�A�{v֨��
K[���Q"O��SnF�^�t0ip\�-�ٙ�"O0�#1+��0��0S�TI�6xc0"O�(y���F���5�Ή�,y�/A��~R��̓2S�H�"l��L���q�I�<1��CIX��#�2`��mq�f�C�<��f�X�1AW�T�!GH����<!�T�*����X `<��H��Iy�<�Eh�gq��A'�8����_�<���W<T�L0�ؙ�F��s$X�8H�
3�S�O��)�
s��p�F&M��xa�"O�41ăGfl<<A��L5?��L0�"O�*�L[�bw\�%[\��"O��iB�OMl�ɖK1|Q^	�"O���2��-L �C�ˢ2��Pd"O�8� �	+7# ��N�!H��#Z�p{Å;�OhY�1�5gp��"k��I�n��B"O��Qf+!�Z�j̎=�Hy�"O,�AcK�(g�&I �	Q�&���"Ob�v�'a|�Ԡ3�mk�V�C"Of	r�Ҵ$yL���ԎL�ftk��',����'l���wcN����	�
Y�k���'9bA��KQ� �t ���q״��'ڠp�cc��,z���[�hܨ��'��!8&�B��Ђ#xhB�q�'��cυ�i��8 �\�E�>`�'�R��ơެ"��!��f��k��DVk�Q?=�G��b|$8 �[�^**�P�(D�jG͎�4m�\P��/i&�J�'#D����S�S����fE��H�މ8bC D��ƅʖ'̝����搽��9D���d���,���Y%B��d����C7D�,��I�5kA��ȇ���So6\���?)�"�o������&�ֈz�.m{�K��C��M��2D� )v��1B�LQRk#�Xb��=D�\H	E���(cgH
��ti�E>D��Hv�I3�D0x����:8¨���0D��C3OQr�~�A���0`���b.D��paԳALj�ᣇ�	^H�Ja��<Q�hPa8���H
0iE�-�����o9>�)�`,D���hV�4�LT'!��2I8d��(D�F��+�誢��*qH򐠡-)D�B���X��Ȑ��_�	�ִ*��;D��Zw@!!+�݁�K�QP�䉔�8�O
rc�O��"$�)RL0Գ�$ʕ,��qR"O�����+y&��0��b��ɓ5"O��c��	�	|�� [<a�h��"O�-���W�}+�&)ֱO%��x"O:�Ie��&��G� �@���"O�˙��ĭA��U�����I|Ɯ�~
�/L )n�}�`�X �\ĩ���d�<y �E^P!�U�D=�%���2T�k3@	sEbC�A��G��i�0D�� �m���ӺB�T�Yr�U�N��M`E"O:,��*�nV|QE�/rDXkG"O��x"�
�l���Ϝ3`�R�@d�'=�]����2$L���ˎ[SL����ǰ!�jh�ȓg�¬jA�J$��B�#n��ȓDs�3�?P�J��F�Sb���#	d!H�);2��am �01�ȓ"���
�3̚l�m�QK��ȓX���,��(�zD�	�b��͕'�\}�q#&�K!�#�dk�_��R%��9�<l�Pc=]���Z P�v�T��&�` �'�B H�Jð�����J�{�������ܮB�\��ȓQRF��
�,��U:���?m�҈��	�,��U[L-( �� ����ۃ1uhB��n��p�Ɉl�(�@��'m(C��52
�B��&k�h��jGzA\B�ɼ+$I�/�%g왠'��gZ,B�I��b�1C�J�-.�UBE
]�H� B䉹{���!S���{�ق�l5B) �=��X�OϾ��Q��0\� Ӆ�ј<V̔j�'U���)�zT�bb��'6p�Y��'a0��ܣ^^��pc?,����ʓEt�X�A�Y�q�Cab��pD�S�<������8Dt��_�D`C�Gj�<����'���rT.�'wjv��V
矀��#4�S�O����GT#��%[RF�Yr�a�"O��aII�w@�"¤N�8P���"O�%�5��A����1T.�r"O8��R�
W��S!O+��Q`"O^p:��͍v]d�:���2�$x�Oz�� �YtAсA�.X*�P�A�O��'�N˓��1h�+r��"��'��T
9}�x9��ɗ %a@ �T�]RBhB`���'"d�!D��T�Lş$M��	�&�O�I�Ad�D�#żJ��1��䔻6�d;o��>�<�֍%0F s�j>Y:���TM��B�L�^�l�i%*�HDY��ݟ��|��X���׉	.n�v%�Sy��'�a|B��0�-Po�=SD������>YfV�`� r{R�xW.��S��]n�dyEGy���'��[>e�����T�I<\����G+�*1��X��{�|-�	U�*	k�
>#=���T�W�o�04��ݟ.c>���oW�+��U����K����gm�T�AO�.y����n�}p��h���H��Y;P��V83o�&s�X� �'�(�����?9�O�O��I�_�1�s���F�B6B��7u0��ȕ?Ƣ�y��*=$�=i�ӻj� y�'D�f��P�����������ɶZ�hi	4Ğ��\�Iܟ,���?�ݱi?4т*�2)�0��\[�|�
��M��*%��76���gK'F��� ��'��`�1$��<��hH��խ�V%ږ�&.$�X��#�]n1���]F�U�س`L�6A(�)�iK��'j���?Ɍ��s�tzǔ:Y[4�з��:�p-Z�2D��.)r.�*%���&�nA�d �r��=��|�����2J��� �[�Ei���@Pz`x�͉s����Ot���O����O��Dk>!��A�:�����Y��0�w�$Rd��>���F��0�� ��$[96�L`�"�
M��0�#
�k3$�rP"́qD�)��"�3Wl`5�Ou�'f��.8��B�o�PI�,{������hO@#>aB� P4T�QSZ(ċ���_�<�妆1�@�j 4�`����\y2Dr���$�<��o��"��S��xͧvuFa��Ҟdm��KZ�NsB5�	�#�.���ҟd�I�^�eA1��W9��ئM�-}s�������k�)2 �q6���H���2g�ɪ+B�QH����$�I)�-n��P�Zw�-9�'D3�0�QؔX�FX��d��%���'1�rT�"G�3*����Œl�W�̇�	:4�݉h<���G�К=��#��'�b���4bTAY�8`$�&oZ�z�`0�'^�A@��'[XxVQ��O��D�'�D�����z�� (Ι�i��Dac�'�,�L��"�P��T� 68���F-��c� ,�割��\�b�5򜼃��Շ8V�)���KO�O&�����:� � rf�"O��y�'}n����?a�O�O��)� ��{6o���QB�8@��}�a"O��C��)u�`������T`C�퉨�ȟ
Xs�H�H@��ӋI�F8��V�x!��(�3�����u�Or8�D�/¬\��G3��S1��{�(�aV#̀J��t��	��P�2Î
�$Q���TT*���sۚ0�Ub`E����xQ�ȓ_��1y��I-h�d�{�������ȓ��-@P.��h�|Ż�
T�K;��	�{���C-^V�r��U��t�	��0D�!��#t�,E��皩~0n�x3�Q+�!�$V�&T��@'�7i&`QfC�z!��5 l�{�+"h�Hm�¡�7`!��T�Ppn�[\1?@�� �@�)Tџ�c�@���MJ>��E�k�jI2�!�/.�ր���;��d�O��D�O|�H�V�c�>�9��ϵ�"���)&Y*���(مY��< �哃0�8�8��[�Q���ɕ�`�|�1��W�Ҿ1�`K�i����O7ð<	�R�#�*d����Q�֔��?!��?�������N�]�tm�
(��p@��&�?��������:�dFд�vLg'uV�K�&�O�E�'u�3�H�F.}K�d[�_lT��*O@���Oh�%��o~rȕ"a*քQg�@�B�z���=�0<Y����>=�1Z�������]8(�Oj7�5񤉿��O�Ը���$�v�2rg�L���O���Hh�O�s�l��&���i�rM��;���@��!Dt0��'uH�'`T��K���K|���6T��8+ ��!pD<<r�'�����yr�}r��b�::c�m�4�!5��(H��J��Vj>}!�~���_��̀g��6���ñ������!}��X1��T|K,�X���@���!���Ѩ�O�a��>A��>9���R��Z٦a��g2}x|K��)U���#�<�QY�DZ�O�Ȑ%/�w��	Q.�8d<2�������2}*��DD�M��,]^�������z�=�,�9������
kyҀ29"�'�8 )�'1�dx����Jب�3�����'+`t�{fڔ��9O$����O�p��\�.,@���N�#�'��)��I�I��|���҂���a
'/�B�	�^tcD��=y�ҝ@s'� [{66!�	���Oy�s�
����D�w�>�s-�]jI�r^���	QybU��'��S�iB��F6r��J�
8A�1'��D{��4�N�W,�%�t�6��Cfe:�y퍩[܊! �eQ�[Y�,7h�!�y�� ^��E Mx����Ē�y�BÚN�vY"%i��F�mYc���yb�,8��#��WD�Xa����y�h�@�ڤ �S�V,�b��y��͵_���x��R
���
:�y$T>z���j�+;Hl|�sE���y�!�=BF��N600I��y�E(qF<�A��Ԗ+��<��	[��y��^wJY���L@�h����y�"ߤ+at��")����k*��'�r�aUo��M^��@'�Mvx�7�X�n�{���2��a��B�"�VA$���Ӡ1�M�G1<Yr��v� �(s�����WD�8!���ɧ���<�p�ːkJ(	Īd�&oD���$؀��iU�42 -H��-�;ai��;� AE��?9�n��u���-�
�OP���׊P閴[f�p�ĥ#"OB|T� MՖ%�C��)zV���"Ov��!��Av���ʑtoN�R"O8�Ys��c��uр��9l��P"OZ�QM '��d�q/�R�"O�����L�GT�(t���]9����"O�D�4&�4=��J0�F�:<DLڤ"O`�S��TM��d :%�|iR"O�)��9[ab��^y�'"O����DڿqU�,z���hr� �$"O�ev�	�ZӘ��Sb�-Xt=&"OvȘ+«:�R!@B(�M0�P��"O�A�Ri�b�nq��^3k,����"O� ڤ0���8��G]M(��3v"O��aU�C37'�P��&�g	�R"OP��v�
�,e6�"���8Uh-�"OT����@���W$X�BG~ś�"O���LU	I6���fڜ<N��"O-���X	]�t��&D!di�"O<0P��r�^-��Z�~�@���"O�|��$��*��x��`�����"Oș������[���p��1q�"O�Up%�<�H���M�E��	(�"O�����T$7���Ō	O�x���"O���a?!};��Y�(���"Ox0b��T�E�̄��"��R�0k�"O��@g#L4Rh��r��E�x�"O������?!7��E#Λ�v<�'"Oh��⩇*u����5�޽���"O����N�,�����bMk&"OL\;�CT#�Ɯ:ń q�q6"O��Z6���X���Z#N7}ߤ�k�"O.���E�dI2���Z{���#"OH$�H�
E�Mr r:!s"O��
V ]I,0�!�V�]Bܲ�"O2�z���<o�dIPlǑG�\:�"O` �K	/`S�p�®yE
|p�"O�0��)2@ %1���`>���"Ov���㍭C��ј�ES.)2<�B%"O�@�F�v'VQ���%9����"O�y{RO@�W$�1�J!+iD��"O�H[ej<T��ى�b�
FPx]HU"O��SCI)
�͒�G�@�D�"O�9#�KU)���Q(�b��,1q"O��[��C�G�("�Ӑ,y��(�"O��2���%A!�D2@�Zj�}��"O�5xG�ʺ�|i�H[�xZFXI�"O��@����r����"��&Cl�	�"Or9t��P��6 F�=	�#g"O�DC+�%M�t��ªr��3"O����ؚNDV�R�L�k|���"O4� vG�
a��C��(�-8�"O*����J�(�tK��Q�Pxa"O�E��ö*�$�b�ͳpU�q"O���V��/o��#Dm	C9\i��"OZ`���U���XIa��q8d���"O�XKD� �|E���G9@`��"O:Ј�ٷҽ��I����"Ou8 )�9�I �T�6�
���"O~�JE��6\��5�R'D
j��"On�ʤ�28~��k��J��Q:`"O�A�7�ΛU�:4�9r�N�+�"OfQq K�=,`��e�nLE��"OPIڗ�6�" ���?OҸ��"O쩉�KB�uJ�FCR�*�z���"O����"֛l�yb�AA?C����'"O*,����S���0�e�&.����"O��i6Iɓ\�J����	�w�9E"O(U�7"XNqE�@�«Igt��*O���P��ky�0�Pc	.*�j)��'��](p�Y�E>���!��&Q��'�������Ph�a(	T��'�,2�+�U��{VD5��A�
�'0^�o�KJ*�臷Z:t��'S�-K�\���2��%)d@lP�'+μP�h��q�Z���	c�8	�'��,c0&O���b��Ǯx>����� ^�2�d@�l.:,+1��L�@�s"Od���Q�Y�E�AB�
' ��a&"O��J0l�L�6�G �NJn䃅"O��-�)�"3��"Or0H#����`�@!��jdc�"OJ����D5��I��#m09!"OҬ�T�n�ȉ{Seߎzl��*"Ottx��̢^�:U䐧kK��i@"O��S�:w���EDZ&��"ODYV�ǳwF�̪��טLD��P"O�9Y���y�r�"#M�qH���r"O:	1�ʊ2H�>P!�@
&|�p�0�"O�)p���J(RR�Ӆq�Z���"O4�Ƞ�>#��cEȁ�(��-y�"Oܔ�M�Y�41�FîF�D��W"O���1[� ���G�o]~q��"O��k��z<��b`
%_R�0+�"O<�:+�+tYX�@`߭OFaH"On��9e�>� ��N7.*��p"O��R�R�K��t×�"jN��"O�y�A/[����y��Чs��1��"O2l� @UWҾ����r�n�W"Ot�Ң'�!��S�/��Qs!"O�\Z�'�X^ܴA�iv��""ObŊ󎐷E�R����ǼMkRu�q"O�iR��'L��d]���4"Oz8񷮌�A ̼1�.�
�H�6"O� ���vu�����7x�e�"O�z�YH�mX%����D�*lj!���~��m��� �.��k]�!�DÌaF�`(�q�~�3g��c�!�$7� 3�̈́���xWҵ
�!���^�v8i�'_�j�n�`/ , !�6	��cfCL)>���T�Pc!���&g���2��;}�sd�]�!�D4\�����ggp<ӣ�W"A!�$�(J}��œ"INNq�.�=1�!�T�*��HXdL�X9�h�u���!��'�
,�s�ǌ_U@��A9(�!�D��X`+ā��R�d(k��	!�$N	Q��ŋa
J�;��i��/�!��|T~�c�_>�\��bc�w�!�,F�B��em\@�x����B�!���rd����9���3@��e!���"Ek
��2���;2/ӰI;!�d��B���Md�&Yh7��!��ѱi����A��8I��"n!�D²@{�9���"�\i
���6�!�.0�"%���M��R������W�!�d� ��&�.zR!zR��*\�!��ü17�4Bi�9ؾk5�	~!�D�.p�-�pE^�'2��B�DM�=j!���R���W�$��V�Uj2!�Q,�-�Ǉ�_���!�d�48��Ą��b�i��ؽtE!�䋼d\T�s"���N���,,[>!�dӷu{�����VJ��$�wiE�0^!�͗~1^����06&²�W�i�!�Ė�.nzAQp�0}�F��%=%�!�d	*0��Fx�r������!��A$h92�A�4MT�"� �N!�'i0���T��NU���ϖL!�W�=s5Aӑ#���j@�A?F��$ &R3�,�5*8}b�E��#��y
� �MА��"Ѭ�)�ޜ-o��a"O�*`޽3P]�6$�(k����"O��BRHۿ6��А�@"aX��9�"Obl�Sc�434�8�g�?W�V�҇"O.��aHP 7��e��$���IA"O���hP��H�v�dyڲ"OPI���(�\��#�	J�j8 �"O�X{�	UK2I�$�� ��ܘ�"O���Bc�w)da0�� �H�1g"O��E�q�yQ�;2���"O�����1�����-KkQ�"O`�����L�<����"Ob	����[�~$��Ā$�x	�"Op�r%�蠴���n{�@��"O���1b��#N��D�Dr|Q"%"OV�Hs�N�BĤ��Ѡ;Y���"O>��`�?K1�dfN�Yv�Q��"OԼ���׃=�"�V�}Y�	z�"O�H`Ģ@�~�y���[ N2�D"O,A�`Ԣ68��D�V,QX�"OF�b�kA;Y֘h���(s��A#"OnQڂ)Ȃ\��D@���d�b"Or=ӃF� ��X�!��|��xt"ONY��ٳ\`
��b�;
�M3&"O���� ��-1�ӕ������ �"O�L����<A�XɈ� /gz��#"O2�5M͕9��X� ��?.W��`E"O�����=h��.W|>� ��"Oڐ�6 � 	�EyBL�K���"Oz	��&��'D�Tö��b/�Dy�"O��04)��Z�� �JX�:z�&"O�虇k�-Csx"�k؂4�Z}�q"O��z�͎+y ���`�,��H
�"O\���EN!`����I*Dt�ED"O,e�Pf--�6��q��?y����b"O2=�$��ѴxF��W����d"O*�OL�b��k�JJ��>ԓ7"OP���͗M\H�pd��z;L�2"O4�����Ú��aS-R7X���"O����E68�YVGE�@L�"O�����Z �������t
�'B6���L �N(C��NުH�
�'������� 1��� 11c@��'� %9��S��&�;�NQ�*Ϭ��'�r]��$��P�����$a�S�'vȱ�*Q�#s�Q� !3gX(�
�'�>�q�Ȋ����EN��l�_�<�DJ��i��m��l��Uа�BL^S�<AR)+(�1ه�
��!����W�<�BH�z�>\)��P
W $��jJV�<i%��]5�� �`U�:�z���j�<	����CX~$h`k�>Y!Fu9��h�<�t�6� �Gn	<T)�D�j�<��ˇ�^f���ჴ5����Af�<�R�-lĲi-b_����c�<IdIX>}E@��%CV+P�H�@�I�<aЀ�R˞�k�-N�*²�`P�A��� �&���[��V#M12T$�,
��'$�"LU.M�:����0D�����T�0T �F?����a1D�Ѧ
F�_#��t,�d�v���K0D�(� &�+5�8�Ղ9����0D�	���!� yc��S:p�F�*�n=D� �-Ş�By"!��}:�4�.D�xq���kI*�V�v�����?D�� N)��d�q;���JVbS���"O���F��FX��7�HxR�m!4"Odr�;(`�i1d��8���"Or�[d%�KR�0D���./�q��"O��+(�5�vU�7�۱t�01�"O���'֑r�0�;�m)FW^�	V"O4����,�Y�Y�"TX � "O�Y�wȒ?w:��e�7�#"O>-��j��J�B�5��P�S"O�T30 ޺(0֨��� u��W��yǑG��,��͑����QL],�y҆�.P��R@jW�P"�BB��y��˰P����ٚ8�R���_��y�F��//>E�p��&^�n�a!�K�y�F��Xt�����סR�L�����y2�\�(Ј�Y5F�Cײ�+�����yB;F
ҥђ&�'4�aW���yRG3[�T�����_Qn� TB�&�y�d�?6<Jy%!� 41�6����y"�F
�����e �8��(�y¥�x�~��QM�
)����	�y	�P]�e*� т��I�y��=�4L�u@w��mU�C��y���xk��A#F�����/'�yR�Y{81��_�^������y",�+5����ǜ�u>�l�,��yb�_�q��a�����k!"�;�y"���P�f��&c*K��0����y�����`K�͛'���e !�y���o�<��h��Δ�B/�>�y"�5�[$�m� ���@��y���X���3B֋:� �H�(E�y"��?~���V��0<��q�� ې�y���MAv5ZS�E.69��!%[�yJ��a��2�(5�L��fT��y���?U]r���<�`��/��y�j�s���C!$.����HU��y��9Z��Y�hɔ{����*[��y�8I��]0�FF�Iy��{�ְ�yr�E�E��U���0I�`�h����y���)L�Ơ�'E4�.b@<y[	�'�h� ��Ո�p��K� A)H	�'l����F>\��`�c,�+�(h[�'�lɁOܼ+�T��3�+����'� �x� ���BxІ���7�l�	�'��|�g�!cz�ɥh?3��2
�'C<Ű��A�`
���Ԣ'�a��'��ѫ@W*?�B)!T��#�4:	�'ղ�!�W��n��a
�lL �'�:1��Hn�;W� ��I�'�r1���E�Q���P��\��I�	�'<"� rDU$Y}D}��ě?~(�b	�'�<<rG�� �d��e8��l;
�'Y� `a̛�^����h�Ҧ ��'��6��S��ѐD"6-�̰	�'x�K$�OQ��
�d�*)��eb	�'/�����X�F\��"T�K�X ��'�T�h077��s�A�4K�`���'�JaP-גI]���s�¾$H�'��x#�Z?] NX`Da��uU
��'0�<���HbUH�jȨ#����'�ʗf^� �Ti7�ZMm��0�'#0Yx�@ɼS��jO�s���1�'�,��Z5@p�)qD�0[�α���� z��Cχ�
-�ِ2Q9���ن"O�S��3i�V�PU� F�
��C"O�uZ�j-A#6l�f+�>,��"Oʍ�c�5k��P�kΗQ�	:2"O04�B�G�(!{1ʝ�!��h"Otd[j�7�R!�)�!+u���'"O���
9p2p��Տ?Hz��"O��pEC.:�-�/&�����"O����A�5�8BD��{��r�"O
I��d�vU����n��:ݠu"O�l��B���A�m�Ln��A%"O��E��yE,��ƕ�[_|-�"O8DZd�H=���r+ě&x��z#"O��� Տ*�x�)4.Mp<!��H�]	�@.��t[��QY!���|��y�F�|�
�2!U� C!�SSZ���@��(� F�]�!�$�`�� :�ג(���H�;Bf!�Q0@j<���T��Ab�W�cI!�Q�iRi�"�����ۊj�!�D��4D\lD�a�>���P�!�d�9C� u�f�Y�~<*Ű`H�??!�$�w߮���K��N��0h�%%!�!S~@�Z6o�p`
����7!��0��)�'Jd��C�N �$!�d��dND6g@�8c�Pt!��:sO 4#c0R� ��3O!�D܍.��ɪ�%�x��p�ӶW�!�˓|X%1R��8e�@��`���!�dR8d�B|hu^�d[ �! 
t�!���
;Qr�H�J ~+xl(���)|�!�D�=J�zX[��ɅM"��k�D�!�E'i���	�(��|�d�
ʓ!.�!�$ ��@,�T��+�d��A�_�T!�ɭOo�Y8��>PXT�T�C�.!�.5te��L*�N�(0�!#!�DP0k~ȩk�d�01���'x!򄃔T$��򇠈� ��90�Aa(B�+`Jt��%�
a�$����'�8C�+K���zvH�(l =�3�C>C�9&�F-p�߄?���0s�÷>�C�I��lżh����'/B�3ޔC�	�{�����
F�VR�5{��¹b��C�ɓ#z~m2%��">�����c�+NlB��<i����� �4c�x�p�jY�{�lC�	�d�n<2UiؿR�J� DV6C�I	>�p5�VO��%X���E�x��C�I�*r�(��HBa����՛BN�C��F���UW�L4q�`��Yf�B�	�u6r�2p$�7+��E�y�^C䉪
+�y�C0���kc��O�VC䉴w��)R!ה���KA�Ұx�bC��5NM��%��?~�h@��A�4C�ɝ6�h�K!��22xtpi�����C䉙pAB�j�ʄ$�b�&B�m~�C�	��x�t�<h#T�?f��C�	*�5�P��W�`8Q��,w�C��cFr���FG�:n)�G	P
OrB����2�, F�,���\B䉨Kv��zSɛwZ�h�ՇA�BB�	~)�xa��J9 �N���c��/�B�	�^���xJ_ @�$��#D�s�B�	�V��݊E�I�<<����(V=:��B��
0���q����f������Q��B�)� L�j#N�;��@���N�a6aa�"O���琿z�,���}?�Y�"O܉��'�9q���`���F>�:�"O�a0mΧ ������Mkt"O�ň�a��;~��v)ŕO�J�"Op���G�x�8-�ɞ G8D)X�"O0M�W��4QV�W=~��9a�"O��q�mK?j]�IRC.'2p���"O`���c�b��S�	6Xj�3T"O&�
���O
v���l�3`��}kV"O6q)�C�)*��ԉ�	U!�5�t"OH�`bsa�(��U���U,N!�Dɢr;İBrd
�%��
E֌8��'h�eʕ�,2�DHV�C�~�qQ�'��i	�#+cR̸!�zh��`�'�|��U��3�Z9$�m��)Q�'3ajC�ܗ*o�Ѐ��0���'��;S �2�Z`�*��Yl���'��L(�L�.��`�ժ�Y�1�'�J�b��H�p<��Ē82A�	�'O��J�&��G Z�1w�2�ച	�'�̨�S&�2,��A��B���J	�'w�1�dkU���.�t9����'���A��C� �n�Y�A�h�$��'\�"���
�b �� �%��'&��r���h �Y9���Xya�'��X�GnG:��yJϓ,9�n-��'�`5� �=��`IE��8���8�'�8pK��������$p^D��'�T�ؠd�E�e/J��2"O|ez왺2�&��cL(C��py�"ODy�cQ�$PF��ĢD�N�N�ٳ"OD-�%�sR�;Gd�,<Ϧ�""OmK�嘏r�x��A�//�p�@"O�9���]�6F��	6�E	 ��,i�"O�yx���> ��3�F��/m�"Oh����;e*f��S��+epM8�"Oz�['�fNJ�!97�<<2�"OXĒ������kć�/��x*#"O��U��nn�t�S��9$�p)0�"ODܫA��*N�$A6�K�3���"O�T��k��C�����1��4	0"O0ͻQ�\�J�t���7]A� �"O��
�_���y��$0U~E��"O
������<Z����^	 �"OڥK��o"q�C�#=���"Or0oQ':q��	���w=��c2"Op}�%�A�
��e0�J��0�"O�I:�K���0s*�=%�9�"O~���i��)T��5įX~d��a"OB����t^�Q��b�4o��P��"O�U�威�A�N��V�ڜ&�\��"Ob� J/rF����Ms��1�"O�t��F�\�$E)�n�<�N���"O|��e]5w'�c�֦S����"Od=���V�A?5��.	N5�%$"O��ѩ� %$��m�ֈ�$"O���
�R`p#��$dRpL�0"Ov��ڤ_�h��[�2D"��P"O���I*qK���D�r"O��u�_�t��1����y�!�PV���b���3�Z���`��,'�' ������#2��cM�			�'��ؠ5���\!���%G3j��'�h���KN/:��l��,��J~�}r��� �t� o�:W�!��OW.'���ya"O�x�c?�v�QB��/y��"OpqP&�_:ĴX�L&v8�m;`"O>�! �E� �*��D�N??4���"O����X2a�<�@A-'��"O���S�4�r,��]�G���y�"O�<�c�A:H,��6�&0s�7"O� �]d��AjA�S�	�kD[�<A�ʆ
<���"�bژz�|X)r�Q�<Yt�ϛe�N���H_qfIs�	N�<Q��̾9ʅ�BӉ)�r|���L�<��Dݗv	|1�e�ROh�q��E_L�<1 Tz���JpX��a	�J�<1a�P
y3ҋ��%�p�F�<1	�-bCh���G	�6(�\a��E�<9מ0oh�ꗬ?���ٲ�G}�<	Q슉pP�#N�;|�٘�g�v�<I��0J=i@���v�J��0�Rp�<W&܀Swxd��(\��}���@�<�DCܢx�x"�اt�f�i�`�<����lΞ�Q��]�	����f�<�C$&��u�֝'@���%��{�<� �G'dj�Re��{�N��'c�|�<1�^z�8KW�E�4O��+u�Xb�<)�A
�c"df��z����e��F�<����<: ��q
]#Y(d;�,Vm�<���J�[��i1��LV���m�<���7DdJ��5ON��ÒgTl�<�@-�+2�Ѳ-�5:�z�c@A�e�<�$��z�،J��Q4$PH{��z�<y'f�g��x�#�$f�
{!KIu�<I�ѥ&� �g�"_JD�
7 �s�<AQ��;�&B�g��1ZT�r��u�<I���<sy ��"�ʤQ�9�,^}�<���� ��%����
ID�<q��LC���EB ("0��H�~�<��n��݁R�^y�H��{�<�a�@9{�@1�H7i�-�o�<i�h�"Ş�3bc��;�r�W�Qm�<adfҼXJ,y�#�1r2�ãg�f�<��=&�l��l�	d`� �M]�<1��E�?�̜`�C��J��x�IBP�<�1��,H�R'�8tF���IL�<�А'[$!B
ZefJ�rEkZC�<Y�'J�h�����P���ř{�<i4��-h6�l��ˬb�����'�tF��f�ѣ�`�J�x���'��aVϋ�/8`���oNJ�J%2�'���G�$8<ܫ�Ayʤ��'y�(�*�5�ʠ���#��'ULervb�'gA�JDf7SZl��'�4��
j�. �dƼ���
�':� �$�V=|K�53�.k�Mx
�'7x��4$іY4��HE.D7��6"O�UJg�ئ J����.ӽ`Y�%�g"O��c�Z.L��}9��8a-V:v"O|t!�L�
2V8�CJ�*(YK�"Ol�T�D�$�ЄO/7��kd"O�A1�ŕl�"}���Y_��Ȩ�"O>�p�_+��黶a��[�Z��E"O,3�%C��>lӇn��i�Hy�"O��3����M�A��(���`b(D�4Ђ�:r�х�'͜����$D��z�J>G��z�@� �h�Q@(>D�� �ؙȅ+T�R'�\d��}��"OV�H�Z$7�I8C�AG� �CV"O�D�����3���^�LqR`O��yr�8�u��A��i��0WGU�yi^��^h�S�4�<�se"Љ�y�	L�w�v ��:(�vI��D��y��}.@�#���6c<�
t�L��y"�W�#�<����10��tx�#�?�ybc\�ږ�x�C��~rp� '�R��yR
7O! �	eh��$ܞ��㚡�yŋ\�t1U�\�mY�xhA�N.�yj�(���3R��8_�P\�0���y�m >�F�a �+(k�I��W��yb/��s���h���)w�p�B���y+eبؒ���$鎬�*��y���k)���E�A\�R⯊'�y"�Fr�+5�Ӟ#��y$�Ƒ�yB�ݵ{=d(�AN��	[`��&⇃�y2�(9{>�q�D~|��R6$���y��!l��9�'�q�~���#Q��y�J3��q�-A�t��U���y��V�{�
�ѱ튾i"���̑�yBFނX8a�6BC#W����&cC��y"LLSL�|�B٨M;���Ed��y���r<��W 	�I�!��m߶�y��
;9��Q@f�D�*b�[t�«�yR�!@�ȰP�.թxt��2�P��y£	Q��� 6���R��0�y�� 0A:���ڒxZ�q�S �y"ō-d@�%�a U(&!��W��y�e�4k�zȳ��_� �����:�yB'�\�(��F)/����䐑�yH:HD�c*[d��1+2����yr�
�,H�1-!	�B�a��]�y2�KCC|��JY��:���f��y�J+͎��Xq�٣2JE��y"���>/�IŎ͝bD0	�`��y��Z�[��c��/�fL;�,�-�y2�߽1вt)Wiѩt,Z���Ǐ�y�����D�c���n��8��͵�y�� UW����n� dҥj��y�Z�
B�ʶ��`޼�"���yr��l��HD�GJ��{B
���y�a��2RH,<_�`�T��9�y�,N�&�0���]~���4K<�y�
�"@ h�nW��`
�J�$�y"��`�T�BQ�B�����y��Njd�X�Eɯ=<�q�����ybB`��	c�J;}h�[p����y�)	�1�^`���rz���$�M��ybgq�H3�F;gM���щ��<C䉆D�g���fcĉ!@ �-P�C�	�D�,���E����->~Z�B�	����Q$j\]��oL�0r~B�	�t�y{�B׽8�t-3R)K2=�8C�	�6$�Q��N!�G�I\C�ɠ7|������7�D��A��8sL.C�X<[�!-\M�@�F�"$C��˟Á�;	���O�8�\l�0�*D���T�]�a�*y�%+Y�F|�!f(D����e��k?49��k&w�8(Б�*D����V�?�2��!S��0�Ȓj4D��8��]bE2�N\�_�H� �7D��Y�+�9�n�٦�7;���±�4D�� �����8!�B�+�D
	����"O�����53XP��B�(��Ƞ"O������XH�,XD$61��ha"O����mQ�PhY	5"]� �d�� "O�,S3B�r=Z�k�UB���"O�)
rbW�TA�<Id�Hc5"	W"Ov̫䉐��> jO����4"O��a��ŮX��	��G�4�t��2"OJ���
?a��Q�#�b�8R"Oƌ�NY�v��I��a���S2"O����K
Gxj��G�r�t�+'"O�hH��]�Sة� V�%ː���"O\"����=� ��r��ئ}!u"O�:w$��/j�l	2J�E�V���"OH�i���2�\D�������"OB�h�4 �� D(M�6q��"O\4y��D�K�^�ⴏK8T�[g"O����O��B�$�:="G"O��9��N�r޸�PcӃ}���HE"OE�B▹rcA! #ԆK�:���"OtqrL8��qb�W���"O:<�&͵�������-���8�"O�$X� �4�  ��I8����6"O�]��%�	dX|��[ah ��"O@@H�g��%��̫�M��%�<�ȣ"OpH8ƈ��F%��Ip)
�h��y�%��4��l�GO/��ѷ)Ϩ�y�F
&�ycd΃3��\t�=�y���h]0�j%�;ؐ+�O��y�/S�$��k�F�D>���$�'�yRI�"��DJ�Bɾ��J� �yb" �-�T���&V�f^x�tc���y�á$1d4�Ҭ�.a1|0�c�y2��H�ڴ�%�+Sc���eQ��yB�_�J�ޝ��OOx�U1�Ԯ�y"�ҍB��,:���R��}�a'J"�yr�hI��Pj�FD��ғ�yRk�#g�P�тų?6Z��Q���y�#�q2�7ʝ�6�z/�yŎ�l�(�6n 9P���	��y"�޺mq\Xi	�3�H�� E�yb����h����"��|RP����y���6�b�bk�!B�����8�yb�b�H9r�D��T�NC8�y���X�C��!���
q`��y�Ş0e� �h�"���F���y2gͯ.�}�BkQ�MЅ@����y'5EV�<*G�Oz��`"�<�y"Ní�
1��4D	�Ɏ�y�m�8t�8*ڔISg���y�ŉ w��冇 �Bqy� �?�yg��;�  f�G��!Z<����M>U:���<�<�������Q���!�C�Bm���0l�=ۮ�ȓ+l��Tbw{(��,��~��ه�ZC
)keGJ�j�����JWn���"'���s
C	{*j��"��^dxX�ȓm�x����0a8L��,^Z:t�ȓN���(�(�� б�l�4�<H�ȓ<]����	YBJhy2�_�2��ȓr�����B;�عi}t ���@�Բ��9f�T�ٵȎ��\�ȓCG
ɸ�FL[ZMP��X�;%���~tⱊ��_��髐���v ��S�? ��@��

�U�a��b���c"O�a�ȁ�9B.)� 럆�Dr�"O��+B*ˀs)�T����!�"O�d��M��QN !��� u@�"O~��3m0��YS�΅�u;&���"O��0��έ�ծ�� 9�"Oℳ�D��!�b�*&ĕI�0u��"OR��GB�n���C=�F�"Onl2#��U�`�t� z��z�"O��K��ƟߤY��Z�
��i�"OL1CV�I�����ؐ�2��"O� �fH���Di����hq"O��Ip$GJAQb���=�<h�"O��`1�A�4�0����*w��[�"O�X��fM�5V��RC���zu�"O|�	��I���D�B���1w"O0�s3��|�0��'����4"�"O�-���*2��'e]a���;�"O�H3�b�\PT$�WD��F�~�y""O�t2���O\�@��(/g:ez�"O"Y�� ]�"`x�2H���<<S�"O�=�H_�E_b��%b�<t�
-kF"O�ň��8	��U�w�O'?�&TI�"O�t�1BX���ihF��	 ����"OͣV�VG�БǤ{�|pE"O�]jrțP+x�s�O�4���G"OX�@�SVT(3�&�:>��0#"O�<�櫆.�Xps#T�!:�a1"O�������n6�Y�F�P�j9����"O��h�0lB2%����7� m��"O~9��k�3:$� r�% ku699V"O�|�G�ޙL����&P<>���p�"O܍x�O��h��F&eO�"O$���Y�~�ʠ��L�:��	�"Ox�أ �;��1��	z$X�"O8)���)b&ĢO�1	�%�"O��Y`�������oG4#_���"O�,��A��8n����5{�2�q5"O���Sh޷v��@�%떋nK*5#"O��	�	�>FA �1:=R���"O�A���s
�8Z��Q�����"O��a���c�`|{��q�nU�6"O� �؅��ARO��s�!�D�d*�k$o7*N��k���,d!�DІ*#np�V��(>��Z�욤~c!򤓀1�\U�Kÿ
4 �뱫��FU!�F�@�R0�SΚh�j"jL.F!������â�Ǌ9�LE�_�2���R�
4�Az�|�a�!�ine�ȓu$��ӷa�=	��šQ�˙r��\��;�`Es��V2����Id@}��Py��p%BӅ1��O	������4m���; �5�c�ta�A��=8X$�w�0��燚��j(�ȓSߌ�R��5wb����F�4���j���+�ǎ6��pE�N�n�ȓf��{��RZ2>m��$ǂ$gА�ȓ{�xH� Ɛ�X�sb�.��X��/�H��٠z�~ �I_Վ$��	��Q��
�y=��4��v�B���'�:��D��,s&�hW;Z�4��,L���")`hBE�4B����R�ةA&&b�������f����ta�����?7�����N�tB�ń�S�? 済bɌ��4d�`���R��"O���cƺO�2�e�sJ(��"O@hP#��-V$��#�'*�h	�"O���&�g�t��b䈎N�"OvUW��!YP<X���+�d@7"OY%nĞ������0�v��"O:4if -Ee\��4�ON����"O�}���̾;�l������	�"O����R�xeę&����7"OZ��n׀\ab�h2%4����"OD�X���4不k���/G#��{�"O�m�ceJ�!뮤ɢC�?0Xq�"O*�s�@ӄmZ�t�a:�����"O.t�B��: ����&[	5�d��"On����f���ʐ,�E#D�Ɇ"Oj�xo�>C) �ȁl�p�D��"ONiPι+YIs
�p�~���"OJ�rq
��t��գ��-�d�ӓ"O��#���Y27�����`��"O�MQ�n\�^�:���ƃ���"O�TS"
�	Y�^$��ߓj�r8��"O��PFY��m3����r��"O�85�,r�M�E�G$1�Lm�"O�J���|v�����q�m�"O�a�g��:}~������<J���"O�I��+�� aQsA@�1��K�"O�i#4,F<��X9���SJ���"O���b�ƭ4���cPh�J?�R�"O���KX��R�폆,7��Q�"O�u3#Dė]�����Đ;(6�a�"O�DS¤&����| �"O2H��n���ډ��蔄{�9PC"Ov���HӶ��)R#��25�DX�"O���B%<-4�Ї�k붑[a"O�}[���}���a�&Զs\dA�"O�E�ңX8�CҤ��z����"O�ɡ ��ƍ�@%�&]x
q��"O$ �t	qFu!��ru�k�"OX���GKF-� �'a��~{�@y�"OČ!��e����sfM�Lq���"O�`��n��Z81��&o�R�"Ot����'H8�8�+��Y_RTڑ"Oj�ّ��(�����ȫBSFŒ�"O���Æ/h�f�3�ꖶ��@�%"O�d��,ʱ�&(�b*�45�0��"O|!��Y�@��[��ǭx�İ��"O@(
(G#Q�Y0a�X���9�"O�(��
+.�p{Q�
E�Z"O�5R�c?Ǣu��^�2���t"Oj�k�e��d�8|��Oٮj��{"O�Xi�m�S:)i��HT[�"O `2�m�Z ��ƀ33݀uˑ"OXdx#Cܮ3ipC��d�0i�v"O6=SBo59$v��B� _���)�"O�Q���\j歫� B�J�L�8�"O��zDM>9�n��Eb\5d��{F"O�0Ad��%A����2�W�N�r���"O��j1㉕4
�L�G���LJ�"O(�ņ��5���G\��>XJc"O�D+�ȝU�43C�W��PE"OjT:�@�B�$�0�$~�����"OH�p�)N�mdF�� ��0vה]h�"OD��HQ���v�I�-��4� "Oȡʢ������	إ#�f|�w"O� �)��s�2Y�3IK /�2��p"O�����$y��CĈw��y��"Obq�@��x��hȟO��Y�R"O�;`L�?B:T��LY�$���"O�r@�7yR���!�6s�9{�"O�W���i � �,԰��"Oni�E���� J-]:�q"O�8�"-?q��P@���%����'s�i+�,F"`�r��`�W=|�q�'��pSh�-;���!m�.���'���h�<�=��&m�)��'戰e����bҊ,D$ȔdWM�<�Ţ�%_v��V��$���c��@�<� �_#	>� �O6~EN�xPL�|�<���6-�P%�R�4.�(��kP`�<a��h1��%J�@8���[�<��͓�t@i$hiE��@��
4�!�$۹� I6�
�	�Y�a�!�$ ��1E�[_��L��,S�R�!�K�&���նL�Di#Ԋׁ0�!�Č� ���A��vr�Y�JZ��!��s\0�r`L��]c�Gi�/r�!򤉦y�>E�����:��	ɥh !�DR�C����5�L�4q>���(O7�!�Ė�*NZ�XR+E Gk���� R=�!���>+�[!F��9	59�@J�2�!��P4��cbT8������$!�΄t*J�S7L��B��蟘 �!��^,W�p1 C�Z�t�B����W�!��P�u^y�O�y���4ꆞB�!��`�uY`���U��,7�!�d�d ���ǇU�fp�m)[�!���4�p0��JZ@�c�J�0�!�dՁ�Z��.�/1�dd�Q	�9
!�,O�|��G��
@�J!��� !�^�a�*�8a���Iឈ u��� !�DB���� �NR-U� ,V�|�!��sF((�u�]���ЩGD:b�!��*4�|Q ��_�~%B�#Q:!��Yr�$�TC�]}��(�"�)�!�d�$P(�q�Ԓ��`"fbH�9
!�T�)&�)p�	��-5�\�!�d��H7,päS�p�$��A��^�!���#eo��[���:0|����]�Lr!�dT�e����B�;�d˷愵SN!��T���(�;�.h�Ȟ�=!���Y$���!lɨG������Ǿ�!�\( Ε
QK^'2����CLQ�!��PU��XB���<���Ń��2�!�d��Vv�𓒡��"5��ΏL�!���
{�C�$��d����X�!��5��1��՚O(���V�_�Q�!�DV����&�h����h�!�� �Wh��C��>[Φ��Ǩ�>�!�H��܈vM*�z�b`ŌZ�!�D��G�D�V��WN�J�!�dӿw���GdY� u$�t��N�!�d��l��	�ӭSXz�!�˃�j!�$�����e�]A�h��T�!�$V�Rl�P����wS�K� �n�!���u��s���1D�#2�� !!�$�?��ē&��@� ]"�G� !�4u<B%�!���>����Z� !�0c9�K����#��3�(�J�!�� �0����7Te	��� �0t젱�"O�[���3^,3/C�0�X�"O�	��X
Kː\�M�*ݐ��"O <�2%�5�n�pAO �D�n���"O�Q��۲s�d�m"*���	V�	���s�%�6d�6�)����P���4l��]BV� �n'qO,����%�R(p�
3}ll�v(߫Bq��J�Oef�Z�&))@`8@�47HvP����
&���f�ߍ(T��K�A�;�h�'Wm���ӡ�7#�b�a� G�� Ez2%���?I��3�v�'���3~���GS�Xh�(2d$�^9\8�������I6��)ȽKF"���&��h4������9��4�M;��8;^Гp���\kAŗz?1���jM��'�V>���M�����˦�:0�X�K�0��	�in>�[��)`�'��5�t�"�f!R��A��b�?e�O��t��&��D��j��(�NXv ��XV�i?d�b��3"�<	���������#�}���\cy��!G%!?����(bX����Ħ�)G��O �n���M��∟��l�+$��ip ��m��</n����?A+O����H��xs���7a3��Ŕbב��l���p'�� F?� �B�$Z3���"U)TH�<yf�Nyi� 8@7�),O|����S�3�Lx9��;�Ȭ[e��+K��Sr��M��G�T�*�'H%2#<�+گl���3���,�ufC/[�l]kE�ĪG�X���^<UQ� �OK�#<�㎟�,�@��R�	�]KS+:���O�<'AzӶ4c����ßէ����8+�ʅy K�R�FC�B3�ONO���ʉL�|�����<:��ɣXp< ޴d����|�N�d�*OX�ca���F��Y�J�D쐹�J�YX4��`�O���O��D�.����O�����a1�����4��B�Y��DJ
�"R�)sNS8C��U�+��O���1H]�F�V@���3����Q�_�Ҩ��)�|(��*ҍS5%%��	�'�(O|b��'ɛFE�(ʠt)�΁�=ۄ�׍+T��m�ԟ �'��U�<�~ZuCъ9̶��G��.�
�F�N��0�S��-����E�������x$v��"�'M^6�٦}�	П̰)���M{��?q��߭ۡF�2��H��c�8̙�cܺ	�@����?y�1m�#�D���h ��\�8P0�q>��d�D�[�`T�P�C�3_�b��8ғu�Ȫu$�4pUj��Gȃ/o�%�Ɗ�={C><с��r�v��eoX�"F��%�_�'�`�Q��?13����i;�RU��2}9*h �d��i�p۱C�O2�"|ʨO�t�ڐ\R(� ���B��B��'j�6-æ}o�<T��0Sצ��aP=!�*���L��6t��ش�?����i�*O����O�7�Z4F�����[�Z��4k��I���_�rA1�,ï6un��g�q��	�|����5&�TPB8�KS	�h��	��M#�i~�I�M�2h�@6����bLq`@�J�����Q4� �H�nD�&��h���֦5���O��l�:�M{���i%��i���ǰI챱℁��f]A��O��(�O�m���(Uo��
1c�eb��j �	�M��i��'���2R!a�ğB��m���ŻfR�,�L>iۓ=�~9�  @�?ݬK0p *X�d2�%�%s�qO�,\ � 7�حsbJpA� �]�$��E4H�{O�H(�/��V�h���F\)n%´�|�'�T��`!�B<�S�Y�/�@�K>�ӆX�'�A�G�?^��R"�x��8u�����P�2���E�\���c�"�?)�`��є]Á�^�8��)@��@J�'`�5��;8��rNXZ(9!"���<_Α�G�	W`�T�ʀ3b�(I���l��IH'�O�``̐���$�%aWDHz%c��!FF(�t�a��	F�IA-PBlв$��8#8���$��� !�v�$�c�3�)z����y���@��% NNQ�,k�A���D��<(e��{���-i�Q�G��ݓU�^�������L��Wn���hO��É��d�a)�Ȓ�����O( �2� ����.}��s4�|��*u��s0N�" ��)��/��|�VX}����w�@�p��<T_̡�!`���?YuO4K�Z�A���]�ƨ��ȇA�'Y�p0JDu@@�3��
�_z�Z�����` �pf��I��[&�QU�ɅH~��C�߂i���rl�>G��]��o�/q��챥��۱��a@D��A�a�F�%ф&T���Naʁj�w���	�K�z�(�*��1�"�k-O2@��i�S�4�A�9-f��(
�B������|1.Kў�F� �$p�@����t�̄I�Ȣ� �#͇.ԮmQǆ�19�(f�,��3=��	yR|�E��65�=�w�"!���挳F��/{$T�˄�Y���d�+���CJU��Z@�q��(R]Q���Q 5}�r�8�T�H�Z������֩} �DPѪ�����P�ēv�`��'��8jv蝚:�ܽ�)ɼ%�b���Ǜ�&ި���**���9�!Q��ܙk�Ӏ%�x��vB�S��;,O�㷆�U���'-��3��dHE#��Ą��D�1�0Q��'��eJA��L�*�q�I�,�*hcV��(x���G��0ɰ_�H��	�J�h��(ێJZ��A��� c�Dχk�T)
���)m@����;O>]��BA�L�Nhv�^nX�0r�o�2b���WNO�h�j�"�<TR-%tU��^�6��H�Gm���O�	"a��7������I���y��xR�2iVT�� ����Z�??u� �4eMYOҍB���wFM�o��L�Viߍs&��'��1�a~r�F1��qG��B:� �"G��~Us�^�]���*���I2����_%g�`��wK��� �&O�[~Tq��Ӂ;ݜ����|Sd�R���S��y����x[�O��2)����3�S�NN�y�T���
��HsOH/{-���d�7kլ�6!��T7�1�C��Fx��'���%��::eN���$A�W��9�J>�E$@�S�qOz�`�(ԋ*p}�S�H�Q�$j����)1M��H!�.bF�iǄ��r�1�g��aК�>9�M�t?����+P!�j�r�bی��'������!���"&�C� E�5�c���Nx�mS�(��|�!�3U�褸g�X/DL����d݇�p?� ��q�D� ��ܝ4���JGT ��'���x��z`���7���w Н��n ^�	��.�T�*���N��#���bC�I��zX𨈏s�<0��P
E�亦��aG�;�h���R 0§T�
�	�fT����9y���x� τvZ�B�I�0N�}�5�ҙ�.��cE�^�	� ç:c�����;\���C�I�P�Q�@e*@7}�����,ݲ3Ox�I�&\Of!I���#z��G��`�8����1~X<�P剘�:=9��[�,��$�	g�D�rFD��P0d�c�!1)��7�p���.[(�P�1砏;�2��A�`��G��  l}�"�371!�� $m�4�V�C��1�r5�=��N�6.#�$:RL׍q�~Xb�cȳ-q����Oꄩ �(.�P�D�ŜA܈�[�
O�tЃoQ�<.��C)I�cb����5-p�d����YT��6*�
��X��ɘU]J=�viرi^�RA���%�'�>-y2�ڛ���������S�N�@Qa�ɞ'�9V&��P�B�8�lSܩ.� D��`2B���3}B��b䄅*���J�8Ӊ�(��>!�@�@�2�pI� ��u��耔�0D����[���gLm6hqǦ�y0�)�@A�F%��G7���>I�I�\��,Uy�E+4� 3��b�*$���ш��=��:�O��1��ݚ1��6mP�0g�y3�E�w��YǓO�UC`��@�ލw��<�f���ɝ�p����'<U(����]6�x�#KQ7eC���W��QH<9� ׃v�x�X�s�P@�WY�<p�50����ő�G��I�Do�@�<�L�C>4�0-�;c{�Yԧ�v�<q���3{t tn�@p��I�q�<�F$
ʁćڵ �x�yAo�j�<!c*�7 T��Q��+&@=�S �i�<���9.ڤ�ӁD)W������q�<ac(����eh$I�h5K���u�<�T�P�x`�ʢNP �'�x�<A���V��9��F	O�1��c�q�<��喞m�F��a�ĄJ�V�8`�p�<�f��6��@Í��Bۼ�j�iX�<"�TZ�@9#AWj��c���o�<�����2�ԝ;�,;.,�P�d�]W�<97�x�6$�Î0^�Xm�FE�U�<	���	#7C^51�z����S�<��E�L�"ݳa�C0;-�ə�c�N�<)�*�"��������l� K��K�<�ǋS6t�^4�&�[
b (�T��K�<Q�ܸKϐ��dǀH��'��B�<1�,ƾ
Q�x�Aj��(�U�Р�{�<@�8k޺l	&B�&1��*1�S�<	�d�	42��1�� ���1#�N�<A1��**�o�U��:7���!����@�YD/ۦkK����D!� ���0�J�?SH�%�7�\�t�!���) ��9��m�=	�<#aDP"n�!�$�Ք��G�yD�c��6=�!�䎌�$dkC�LJa�)��!�O?|�R}JL�b *a�[��!�%L�И���$C���
s.��S�!����5�ѥ�[��UZ��K�(�!�ĕ"4cb;�� �$�t!�dV�h�����0V ��%F�!���q܎��r'J�&D������,}!�
�d����$ș\���C1�q�!�
�1��aA�F�/��a�5��r�!�DS�{G.=�B�I�F�&��v��3V�!򤛖SVDȀ�+�����H�a!�d�	4����BٞfD9Ks��G�!�DI	�"��$
�|�@�= !�$�H$�`�ݶB�Z]�A�6HK!���Z�䣁L{�X�@J�BK!�E9L�L�h�'YuRd�s!�	D��`��a^!qN���=&!�dL�6 !��/�
|��E�Nf!�D�$��iЩ|�JP��_2b!��X��;Pe}aMM�*6��d"O@H RF^�V�ԼT
ڬ����"O�ph2��5�����px���t"Ox��(�'�`���[2TlJ�x1"O(�U䊐*r��K�&W0(�Z5"O� v�����1S�&Y��^�G��u
�"O��x��͠9Y�4�u'�8����"O�����\.>�p'g�<���!�"OPAr��f^D�'O�<Bn1"�"O̡�a�"�")d,6d �xF"O�3��20�&���-&�P܋%"O��P��I�p�H(#AT ��	@�"O4(��bO2&���!��V��(�v"O �If>p"u�P�ܴ"�Ի�"O�D�e��'Vg:�	�%G�Pj�BC"O�Q�f%ւh~�P[�	Ѱ�ptH�"ON౑�b�t�zʋ�C���R"O~����ɞ��T	���
�C"OF���S�z���nY�x�
��"OʘCd�F�x����-�4;lp"Ov�'. !���ŇΎ@���"O� p�'��j��Y�A��,��ش"Ox0)4F�
*.�"F� 2k���*"Otг�,^�s�������\��"O$x���P?#�*@9�n<W�"(1�"O2��P�30��Y�T���{�:��"O|`%�"v��crk^�|�4�v"O����Z �Z���Jſ6Q�%x�"O�<�����r�i&�?J��I(u"O�`�b�.�Z�F�..f� �"O��  �)wSd��%NMj�a"Oah)�$���Ӣ^�	�(w"Orĉ4@�\�A���г.�0a�"OH!�&���]�f�:�A4"�f��0"O61c@e� ,���喟@\DS�"ON�j�KŭtWl���EI"y . ҵ"O�ya�>
w��P��V�y��\��"O�EE�
G�8�׈�A�Э�"O�l�e�^�,M1�1�<y�"O��*O�\<�� �"w2-��"O@��P�F#xz 4� �V�v�1e"O�5�pL�"JNA�g�M�BZ���"O����c�Oml]C��'Z�k�"O���{!U�Q1LE
L��"O�P�wJ#{k�r�ՇB=�"OR�Xڄ
��x���D7Zt�T�'D��g��<8��'D�?����%�0D��X��G1i�^�SAK�$uv�3�+.D�xb��@�nP+�D�*(D<�7� D�(�7��$ \y��8#H���M!D��xA�_��`��ݔG��툕5D��{Bb]�K�$�cV@���w�W��yBM4lb�� � ��>��s�y����\����r��ãN՞�y¬�T�p�SC��q����"i-�yB�#_L�1sA�9c�t���ED�y�e#v�`�Q�K-:bp �hK��y�%�)Ye�<�[�8B�S	@��8	�'~2��dL�%:�����d�T��'��Y�g�>A��2���(U��i8�'� T�%� -3�]��K3KU����'
��e�ӗM4´p%"^�E�Nt��'���y��:1-��˴�Z�,�����'�B�CH u{���$攫�ޱ�
�'���7��$�z�GC=ek���	�'F��ZC&�'oJY����?X��� 
�'����Sk� ,~�-�V��'���(�'à$)ǩU�e�M����0� "�'h�CN!+��!�&��|��1��HO� �t	���:Kb�����9�F$Q�"OtpHr(C c�S���64��\��"O����	B� ���%N�v�X5S�"O�����5����Q�>>�X�"O$�f��*����NN�F(��3"O �IP"]+{8���!��a��"O���d 	*���%�	!*�,��"O��z�aT�~��0�Z�Z<������I�Eִ�RgO�"�@1(R�J��B�	�sV��6FT���!;�"9� B䉁#�P]0UM�"�(M�dѼd�C�Ni�% r# �35��8B�P��C�I�#05�AȿsF�}�%��v�C�I7Z���a������+ B�_�C�I�3�,�T�!S$zT'^[B�	�m��de	�$��)휇9B�I�-da �/
�a4�a�'�F�P�.B�I6������� �|���CY��C䉹5�2��"�l�2]��H�#q��B�	�"\�H����;��}��O��$��B��t|�ԢscI&7��@�	�Sb�B�	4��Rv��^�-8�䈢�\B��5qZX�J�ʈ�xq��:-B�ɰ3d�A���̹u&��j��""�BB�Y�$�	�o�_6�X0�	a2B�I)Uʐ�r�_�0s��"O �#%(�b��h����ѹ�"O|l��@P!ZLf�S��(��Z�@�!�S8o��Q �.��g_���D�!!��>�jp�'�ï,<��&�Z_���;�O��8�L_9��L�ĀN�|T�	&"O@;R������h�/8���[Q"Oʰ�4%��2s�0s"h@�,���"O6D�ǂP/9���5'�=fٌ�d"Ou���H!4�
V���������'�qO�֩� "���CF��dU�D�)|OZ��k[�m�0�$M!L\\K!"Ov<�A�Ʈ� Eۧ�� W8-р"ON
�%�f���vc�xn�Ye"O y� ��9y`���AB��"X`�h"O��)Dk����L��gŷbh���"Of��C�Ꚑ�fk]�e
��'��ɱ/�6Ւ�̈́�d$┢�	
�.B䉍	V!j%l����|eG;i<`C��!=#�DJ�i�b����_/O�*C�ɛQ*�P��F�dŮ�A�o^�t��B�� ��ǩ�2�0\(TL�AdC��
{ר<ـ�/L�$��Y2
��B��?7��)0��x˔L
UHSXc�C�I!	V�ֆ�eؾQ��Ǐ�Z/�C��:�uz��Hߨ�	�B��Z�xC�	�J�	`d�	�!΢IɃ�1{Z
B�	WSL�����a�tգa��F��C�I 0��-����$9�0�U�Q�`��B�I���dqb�=7���T�Ι:��C��/H���"��G�,��,��B�-�C�'NP���Vy<��amM�TK�C� cV�h������=���K+w�C�	�KS��c��$2g�5�"L4�C�	�`~9����+�F�[SaV�+Q�C�	n��A����x
��a(W�-�hC�ɒa��mvEZ�f��U䔙�LC�.ń bB*�.Q �0�ӍHC�	�h�¤�8��`��(_C�)� T�j�A�JK�;'$G?}�$ x!"O
E5)�g��IK�Ó�{�
�"O�5�Q���c�H`т�8j�59"O��y�H�F�0����^W�ղP"OԤ!% _#b�U(7FZ�O\:0��"O�5�q�����ء��1X?�L*2"O�Aa6�ås���
�Э:h`J�"Ox��Ul��8�K�$X�H��	�"O�A�U��+\dxy��I1`�6	��"ON��R@L�?����e"�3Bt�Ź"O\��U�˜u���+vf�fb��X3"O�|���VJ�(�t��"?�)B�"Or�����iJȠ��0r�_5!�d׫f���A�o3�њ�jH�G)!�䁪>���pTk�L/X����M�C!!��'��mD+�5{d١�
(�!� [޺<�3��:aĀ��)]�/�!��D�|��PɈ�eQ�! !�!�$P"xt���MWg1�TC���p�!�D 27r�(ackH(_��*/V�]�!�D.N�Q��.Ϛ:!j��5��>P!�$N%L4u 6OߘF��$��N3!�$G�4���*:l��@�,�;T�!�H�)!�� �+_�t`�q�K��f�!�DE�@�GO�JJ8��f��R�!�I����֥5xh�0��NM�C䉎C{8e�c-��VJ��'�	��C�	&�"��bR�`�ҴS'`2f�C���ِF�'���gE��{���	y�&)X�e9yC�d�u�F:�!�E	d%2��3(0�(e��a!���x�j�J��'*,%{��/U!�.�Pڲ��K;��[t�Q'T!�Ğ���Jc�I;\!���O�P!��y]3$	�*�Ȅ!5��RF!��=�b�Ѐ��:���*��I2!��ޏq�y1� ��R��L�w!�D�;Mb��qUD�l!Z�+�r!��0_�
����C�n!�d��R�:�v���D�];4CV��!�C�<�Z�-Xw�%k3��h�!�d1r'�!�% �>Y����;B�!�dU	�n�HgH�k�6�����t!�d@$U% ĸ� T� ��r�͠7Z!��L� ��PB5������CM/dO!���,Q��	@C�H���hFB�Y!�$֟d� H�-B�w����(�i�!�DL�A@P�p�W"Lzn�S���&N�!���uF��+V�N^[:1�7�)z!�d� N8�|��ʂ�G�2�ȅ$P�x!�d�#)pb�RG(�hΪ9CQ�^X!��].�!�S���p�M�#W!�$�?1�`�a���(��0H����oT!�䀩v�4Q9҇��W 
��t�HD!�7�~�qd��?m�ۓ��2!�H�<�zq�B���m�c,��w0!�$��z��	X�X��|�*� ]!��C�Zkl��!�r�X�(Q52Y!�1W�N)�5g�Sr��Z�P�wg!��}��@N�
��:�j/g�Jy

�'mz]S+__R����˵Zz�C	�'�N������/�}�f͟� ����'��A���'^ȾX�en<BQ��'b*y$	{F�H�R�ļ�N/�y
� *��'�	n�D��@���r��b"OTԊ ��=�n���U �p��t"O^E	5ʓ�C�m@L!/q�	{�"O�I	r��5C���*�3d[�4��"O����S[,$�Q
�	@Z�a�"O|ui c�Y+ƱZ�"�-a0<;p"O����o��A��{A��"O��8�ν��G�ߞQ�p%x�"O�!��){�.��`��S���Y'"Oi� Y	dP ������@�����"OF�
� *D�@��&���"O&<iG��2J\^�"FOV�k��aG"Or2� _ m���Ƨի*0훓"O�x��FW�S0�D�QF(Vq�q"O�A��N3]���qD�+��x�"O�RbU��Y�e�0u<-�7"O*}�DϞV%h��ga�u<�,""O(�;ԍ��]�ؙ�v��S*���"OZ=��i�-�eӣ��X.bț�"O$%q&Y�*����D��$"O���O_GL]pRg��xt��"O0���ᖈ?�R���凇9m���"O���&@','�Ez`�ė@O�(�"O(<�{ځ�Hܸf�|���"Ob��m�$Q@�d��)�pঈI�"OB5�&i	#O�؁v�])eü�Q"OLd`��F??Z��F.N�Z� �"Ot%jG��8q�#�e�e�.Y�"O���ѥ��2�J��pOb�9�0"Oِ2���&��ha"l��*e"OZH�5 ¸����d��Ĩr�"O�y����Gs�Y;1�2c��C6"O0�s���N���qp!�=p�H�p"O8�)�O]Wp�	ƯF�F�JqB'"O�)W�ʞvL* ���%B����"OH\��l�0��4A���?P�N8U"OɃb��7�=0���t�"l@5"O���1��.�pQ�"��=%6b�"OPp ��-u�T��P�ҸsHY�p"Op��b�?ydJle�T�{�H� "O� ���<?�^TCѯ��sֺ�CV"O�	V/�lڥ11����I��"O.!:�
�>y�b�£��\YZe"O0[P��R�$4`f�,J�P�h"O���UmS�n��a &]���S�"O�(�a&/ؽQb�ū
��ࡕ"OZ����N���*	R���q"O��E�����SI����c'"O���"�cxl������y�(��s"OM�@���L��GF�3���Ҕ"O� gP>6�ZD� �7p0< P"Oꉊ�j^�#���(6�<
�y�"O���kO!6�"�]�w�6��"OΌ 3iȂ3!��1���0?�"�*"O0�3���|��-(5�"�@"O������V�p���̦2��0`"O���$�H��:8���������<�Ǡ[I�	ٵo�)>���:%�z�< B�6�PR�!�-`8��0#IN�<)�ᙖ&NY� B*^{^ DD�A�<a�F4"��-��Ɯ:-�H�m�z�<���ϝ*�z� tj�i] `�Zp�<Yd��9�D���ұ~��Qq�<9�� kG���R`�&1�#Ώi�<� x�{"�R.���`19�Hs"OL��f$�3J`|��K�2�P���"O^-zc�S4G�X�A����L��@"O��d�@Q�t���-���҄"O0���|���#G+��Z���"O��yj����|��T�&60id"OR�8��.X��Qb$�EF"O�q�Ei�,id�
.h򊴊�"O`XR]�X��ua�ϗu�t��"OQ���B5g]� g�9Ħ��"OP�1V�&1�����g�3\��Y"O1* B�:DN,P���4M�D�D"O��:��]��lcG���q����E"O�!�R.ρd�Y��ѕ~��� 	�'Ȱ����uƄAr�b7o����'7�г�Z(f X
�C�l	B�`�'��I��Ē�c.ZkD��b\t	�
�'��aN$]���+^;Mw�9z
�'��@���=��R�^�J�$�	�'/�� �<+�t��HA�����'�"�!��=jFp���>.x�[�'�n���لX"Zْ�jѯ0�x��
�'�P]�dmo˞�
 (ɂ]e�E9
�'I�US7�M�tE+$#�Yݐ�{	�'qB��+\�0C�9}�	�'T����ֿ4(�ˡ��:��Ѐ	�'�#P�؅g�1��/xi��'f�0�N$h�*��HX%)���A�'I��Vb�%w� ��N�P  P�
�'�����zWt�%��y�����'�� 
�ː,�@�-ܐp�z�x�'4��pa2���d�T���!	�'����`���#���tݱ�'L��H��GA��[쉽r����'�H�0$S�:��a��#V 9{���
�'��0���Q���e��b�T1�'��jƊD�,�je@�,�VԮ��'z�DA��R:
\4� �ꏆG����'A�e� iͲc�h*�8KQ�8;�'h�y$�ڻ�VȨ�'/8r����'J&Ps���r�ا-��ZG��'�n(��*���₹TT�I��'^���R,dI����L*N�$���'<��K�F����C�[����p�'<FpJ&ĝ�y>��@�נA.�'�r�2�Q$����_!W�� �'���t��>iLm�W�A�w�p�[�'5��i��bL���2p��Y�'�0����/	x �懜��.Y��'� �Y�KS Ux�r��I�6����'-���o�#=;*l����50ZP9�'F�XaQʆ�:�6��BX"<���'7�YP�25�.������8KFXr�'+d���A� ��5ZR�.3��)Y�'��Qs/�$dF m�֡B�/&M��'����3��
#�~���Ŧ``	�'���J�	"z��F�E-<)���'�bs�Y�C�ГU�A�2}���'��u�3��8����98!i��'{
�
�e?UZ��i��4tl��'�`���2a���� P.4c�Ą�Y�¼����`~vz����!�t�<qE�O����4B0c�H�K6��r�<�7�Q�<���q���P��t���q�<� J}K�N!{ɚ�Sw�\�>7��C4"OD��r��*A���+Ṕ!�l�"Oʅ�T�ñB�4`Nߧ
�2d�"Ot�Q���4RZ�y�OӾV�@�"O�I f �=����.q�b��Q"O6X*a�ٗ]Jt�xC�T�����"O�u�P�O���w�Z%v�0�"O()�¨���
�KÉ^X��'
ly(�ϔnĤb��|�d�
�'�BHʃ�I]�l���0$g��#�'8��i�b�
"q��0��
�'��
���\C�-�$+��|i
�'�*����ϸj�4�PRG�(��͸	�'�*�k��:-y�u*��W��T)��'���#�4�Z{h���J���'P@89�l�)$���@���DA��'�,��Q�օX��z�끠Z����'Y�5���^3�eC�Q�)���Q���/O�r�%A^��ܣ��_�f��KR"O��(օ��x��Yp�ZK�q�"O����Z����� #V�`��"O�abȖ�y+ez�K��̚@"O@;f!V<6��D��a���Z�"Oq3��R�8Y�0q�@��P��a�!"O���cD�*1 ��1!EQ�"���r�"O���vMU�N��!J �ƀD�����"O�ы�{xDŃ�V�{ʗ����hOq�$�2d[�QLt�@s̉�h:M��"O���$��O:\5��퐄� "O���?�����VQ�"ORl�A���
���U�AK@^�{�"O ��L:t���q� IT���"Oh��� @x��\���F	��S�"O�
�fÛxz^AXX	s�-" B�Y�<qu�.e�n����<SEj�qVA�o�<I�1l�"�KB
�(��uk	j�<�d�G(#�6=�$N��*~���C_�<�% ���� �^ش�R3	V\�<��ȹ#��2'��egkW[�<a��"8&�[e��TcD��#��X�<Y���NTFE2�	�{�Q ��TR�<���Ͳ�] !�	����D��J�<Iq�Y'�l`F�S�h%
�#%��E�<�B�	�B�����3wkV"dŒ �ȓJv��aP�n��`"��˜z��ȓJ>��j�q���E�tD{��'��� VB3,J�����w��F�NL�<A�����&1�� K<
��q�<!V%	'_��1��L��*�!���n�<ag�#2�@u����� ɖ`�<��c��f�nyMK4�J�@\�<���B���(@�τ5�L�1�m�<!CD�gi��x�8=��!"VK�a�'�axr�9t~�:�HF�w?�� T����y"Dл;�h�"��lv�2��T���x�W�O&�P�wc�3�z�'�*1!�\#gEvh�VLR	{Rj	⒮F�Py��E\��f��?"�U�S ��y�/�*rV��'��'��B����yR+
��r��G&E�B-(����=	�y�D�#n��9�#�/2�	���y"#4�D���GF:[(9Ѓ���yrh�v�dJ��͢%���3G�(�y�`�>]D\�����5�q3�E�9�y
� B�j��
q�V�[G�5z^F�BP�F{��2,n�Ui �9y��cS"X�P�!��Θ8����Kx�1*��.�ў��l8�I$�Ƈ^5 M ݈m�*B䉺b�.T���Ԁ4��d�voE�C�Iu����i�)rt�xf�����C�
�лf㜹j��Z���I>fC䉜v�VB�M�~"���G�4C�	�}�Tx�!�S���0�kX"C��;R��GK�"ܼ�{gB�6��B�	 @E����!T!`��ŅP��B�ɵAU�@匜j�\���OWt� G{J?)�h�
`Ƽ����cx|m�pB"D���1�I(�a(��=q�!�3�>D��{uBR�YK��h�����:���O���>�ѥ,U�NPԳKT3�3�7D��R��	5D���%p��D"On@ZTFY+{ఠ�7��D}���#�(� �Sܧ!�N�ʇ�;6رJ�hV�aǂX���^yR�Y�%t,`�n�H�A�aD$!�d1qd���j�-$�1�nݹ<!�dX%bL��'\:u
|����53!�D:JȄ2(�'�����F
AyR�'p�|���ܲdVaAND-u"
u�����!�@[jX�bƇfvR1��"�!�
se��Ss�H���J�@�!��lW̤���p�YB��j�!�d��A$59d��.����E��]5!��ΐoQд@�DA��|]�,�"g �}���0(�&ժS�B����� y���Q*�<A.O~�OQ>Փ���U�(�h�g?u��)�k6D�{"�ŞjǮeȆGM"x㴡r�4��hO��$Ï{�HQU����c�ՂE���d3���z��z�
R�Q����VGM&}&�1�ȓN�Ω
0��C�Bd@�=K�����5��X8V��F����֥�8Ur\���IF�')���ӢPY>-˻d�0,O����OH�OQ>��C�4r�	���y�f�1�m-|O|b�l��/H4�R����410@ʶ�<�����M��d�D�Ď4ظ��AԳGU�B䉔<BD���k�`�J���7/�|B�	�vDY��V]6`!��,dB�	�S��Q�,�p�S���d��C��!�LlC��=c�<� ����O��C�IX0��F)��5\6���ڼK����"�&�
I�"Ϸ1�p|��-��7Э�ȓ~�"��eʹA1"y֣M�4��!�Ɠ `�]+��.!�,�+�b�D��8��'�*��f�lv���q��=B�,�Z�'ǶH1#e�q��Aqc؅J���(OZ�=E�d������"�:Z�����y�m���m#�D*A�}p#C���y���:٪p��µ� �9�D���y��C.i�����(=R��
���y�/U�so������$��;�i��y⦁.T�����}���LD��y�� &��ㅅ^�j��hFi��y2��.��e��%�)P�ȱ�hV��y�'��3����&�E�o����'��y��Y�pSTY�w�ڸgb@�f/̂�hO��D;�}�j��bh�,w��=x��\]��`���hO?e���JW�����3;�*�Q�op�<�@�� ���xT+Y&�*��a;D��f��8T����;4���Q�3D�� ����!`�����n�9_�T'��G{�O���:筅�b#*�Y���<�]
�'�:=)���M?��0��@�G��ٱ�'Q�A{f}�����D�%3)h�Q���1��+@�Ŝ���X�N�nQ:d�2�SV�<�@Ȃ}!>�0F����!ƁJ�<�d%I�4ԡ���Qr� �d�����#?���/>	��H'�BbY��ӥEC�<� e��衢��qb0�#Z}�<�#�(dzZ͢���\����W��Myb�)ʧ"�j�'CU��Y	`�J/1�z���nnD�ʆ ,�u
F�\(2�X�ȓMz����
{�<�{V�*1��ه��8L�`>u�hk��K?F���ȓ2��%bnK)А���ʏ�8e�?ӓB蠄x�H�%����.;6�ܴ��{	�� �*]�[T�AQhK/I]�x��j�P��% �:tI��!�ȇ�Y�(: �M�j�x�Qd��c�
@�ȓ}+.Ha�ǈ7�B��+�V���F�P�s��8�ّ�.�f�� ��v���������{����<J��8��0ړ�hO�ɾs݂��DC"v��̂��/�C䉎:�<-��Z� z�����?H���O������p@�Pc�R�x젶�дo��j��TI���=DV�4Z��a� �'�y�߲9hxK������b���y�IM.&m�#�� u@t��Q䔕��&�S�O�굃��(�������b$�i��'�J�k�Ο�Ma�����[��i�'B0!��Ș!r��!m�@�1�
�':`,JwlE9�1��IAH@
��yB)-��j��	,��fC��y���BN��fj�z��\���4�y"��¡�djp	 �!6r�����������Պ+,�)��ϖ=G�bO޸hR"��T��f���p%�"Ov��b��\Gԍ��˖L�H��'H1Oj���'H� 6̋BC;S��qK�"O� 0�DV;{n�T�C�	"1�����"O�`B��6h��� K)����"O�2�V�1�H`�%��@<��"OYj'�ǵP֊Iأ		��xy"O�xP���
aڹ��[��D�b"O�l�r)��o��#�&F�6�|"O��x�`�"�� �PºHP�"O�PX���b{�@K��J�c�0�Q"O�ѳU��S�m�v*�X� ��"O�(9Qn�	8���"D�w���2"Of41u�E$���T��t��h�"Ov�S����[$�B�LB�9@"On���HY�!���z��~>�|Pv�D&�S���,%����1�֫0��CQ�!�d�<O49��I���h��j9 �!�N)��A�G�z9���ǁ�!�ċH%W&U�g� �`�-j��� ��Y�)�'o��]+��9f�.xrW�X���$��劗�	�I��B`��h��
2P����>	t-����+(�F��''ў�|�dӏM�S�>�r	Ы�[�<YD۰e��c+�	4�dЀvJW�<��Գ@^}'�Y�@�Lå��Q�<��N̡nt } �Н2n���Bx�\�'�8I�*Abm1��[	b��`�#"O� ����[���ٛ'�0e:�"O �*�5�P�zAC7���J@"OI�/�);1����ۣN���a%"O�tz�L�+1����'��FWԑ�"OH|�5 c��dr� 0I��"O��Q��@	[����j!9Ʉt�!Z�������&��|�&[B���` A�	2�u�もb�<���ڔ<�`I�I�����᠇S�<��ϋD`�@��K9��H�1dDR�<E��)t�5۠h�L��Eb3�R�<��C�j��`����a�V��� \y�<���b�@�yw���qj֮�y�<1g�?�|�b�J�ZϘu;��Ku�<�%�FX��UP� Ø{��Q�C@��D{��)�#�<|cD)��[P\���	IzB�ɿTq(+��ĨAֆ�ZԆI�vB�I�gjh����)|�,��,^(8B�� O��2�^�(�n��Ӊ7Z�B�Is�40����0Y�P���ȈK��C䉷P��(�/uO ��#.g��C��<@� 	W.��H�ՙ�=�
ç\��D�1 تSgV�u*�%t����,��i9�"I3U�����C9��ȓT��i���y� @K�)�ڼ��B��y{����g�"E�I�F���ȓ � 쟩Q�|ք�:�:��ȓ`5���盙&�pP,4(̆ȓEo|uóbQ�=��4�w��|�
�&���I�GjZl+B�:<?Τ�
�<] C�<q($㡒�q�`۳-ȲY��B�)�jE��bʛL"ƈ��,�,>�B�	$n亙��A���L�n�=#v`B�"=i�a�f �[������̓P4B�It� ���,/�EHf��:9�B�I�(I��K��e<`kE_oHv�=��,&���$��T�Ĺ�A�
�`�ȓ�v8��6iN|��͔�|��X��L%�eKŮ�R򖥨V��8=^Y���x��6%��ӄ�����ȓNN�=���܎q�xP@շ	�H���%��|;�0�Tl�c�ٓR�Mth<�T�L��|9�+�8p�
v�>�y��8uO0�+T�M���XE�G'�y� ���&���&��d�P�CX0�yI�s�\i�ŚpP�W#I���'掭 
�O,���O9R��hƈV��-��G�.�	G���|�TyK�i�0/�|��ȓ?��tf%��D����&ʖt�ȓN(`0�#
�j�#R��[�ȓ]""l��O�9z@F٪@ ����ȓ�#0��p�"�Z����d�H����vAJ%�ٕ��¢�eqHD{"�'�B���D%u��I��;lL�!�'��W�']>8��ę%�2�'�xM/}�\ᛒ�K�KǬA�� m�<��ٹ#Q���R�ܜ�@;u��h�<)�/�*`*�b�D�-	ʤg@P�<���	YӐ9`�]6K���IN�<1��T�pY0����Ɩc�Z�Q�lDM�<��Lļy���fD�3&�+ ��S�<�@�U�O(��镫H���5!O�G�<�,Y
t��H�+ˌ	:�m���|�<�b�?4��Z�*�|6����<�F"��g����J0b#�	��O~�<� �,���F1*����HN5->]c�"OJ���hXu�	�g�cL���"O.�����TƑ�c�T	D��0"O��V	��4U"-Q� ��Wg�y� ��Hpv���ׄ50`�n��y!�Z���q�N�]̀�VO��y��DKN����2���ӄ�R�y�L%Y��Q35�R� �l�r�m@2�y�o�J2�u0�4(�.�����y��k9 i�,�v���� �y�o��<�(��IT�m`�[@�L �y�D��?�8!2��u��Ų7	�yR�ςunlyQ����f=B� �����hOq�<�n��7�R��V�@�;��a�%"O�� aL�g�R\J��Y��p&"O��2��'6~�L��hD� �F�J�"O�I[�dT0z8z�;�-$��=��"Ox�@�Ѣ/:�CDN��;sD�k�"Ozh��AZdw�!C%��V"%�3"O0U�P��U��e
]=DyRc"O�aP��Z�> ����T��"Oj���@ܽZ�|5:0 �p� �"O���i��f�R�X$5(ܩ"O�a�3��~r�3iG!֘I�"OP�AA�[�UU�5��W�,��UHV"O��P��pwy=6�@ģD�'61OX�ȱ-ɱ>B��S����k"OV0��� #r�̣1`��+`±�"Of�����j�*����nk�Q�"OҸY�b��D��`���+I�1O�!��)�Ӛ��i��g�a���ȱ��2P�C�0^8�V�d��q��Ђz��B�I�SNhz$/�T����EP�A�z��2?�5䕠r"�b�D=h*%P&J�h�<qdo�ry�$1R������${�<q�h
����(T(�94�\b��Rz�<1A�IPąP�=O��Q��m�`�'�a���!�e���V>l��� ϒ�y�A�=U	D)���ˮi���5�L	�yB�۠v���Ѝ] TVj�U����?��'ǘ�KE�HsJ��ˤ��$W����'�X5Y�IC�:i�K����'������=q�Jz0��l�h[	�'����(��Q�����2Q]Z�x�'9Vx�׃�8��a`��ъ�D���':�|[4螣<�0�"�"�<	���'��9��J�.*��C�GF>�"����?ٜ'�4�F� f^���2OH]Nٺ�"��%�	-9]tà���^�R��6^��C�	�,��h�'�Ƅp��T���C䉥p�Re(�ʒ1K=R�q�ڡB�6c��@��#�Şh\%���#Ʋ�h�叇`x4̆ȓWd�qg,~�0h��σ|���ȓZ�֡�@��Jq+�j�=|'���ȓq� }�Gt�րK���.�z����=B��=�d[��68���ȓG��l�@@�!|�J���-9o�h�� �)�&@�#��H�U
 ���'��B���Ӽj��m��-P)��p0j�Pg�B�qH��J��F9��0I�c� d�B�I5+��,��g;�ڸ*�"ѥy�B�I���@I��f�DY�UW4B�ɕ�l���P�o�L�ҡD	� B�	����Z!g03��ԒA@¥��"O� ��q��9H����Ǟ�|�ɠ�IL>�9� �P���6�˴D�޽���6D�(��iG�;D���	��i�7D�|�EĎx��a����>{t�0un4D�<C&�� rs���#[, ���3D���Q$E=��H�
 ��l2D�4�HRK�Vͨ��҉F��a��2D�h�S�оBA�aѣs�|0�l3D�8	v"G���"�`�	�lB�2D�\�S.Eo�t��Z� x֘1V-&D�t"S�@b*L� t�&���т�9D�85JU�l@Fk��k��8�$D��k�d@�E�� �r� R��&I.D���w
��C`)��!J�;�t��4d,D���tBH��(�+���<)�!J>�����1(6�3�G<���pB�r�!�D!JHh���IMj�Հ���2��\��y�n�3/�ej�m��yr!�;ux�I����P�d��*�y�	�Iּq�D'���=���?y����$AK�4��	¼_�x}��Ly
��:M�9���(JF��H������'�jqs������rp�0#]~��Ǜ*��a"O��H� ٽmq��EH=v�V9�1"OE�EF$#�>�`�#S�-:r"O�T��j����91
�6�&�"O�!���W�+�ڗ�J:<m�4"OL�r0K:WNZ`)E�ƺD#���W"O�j�IM�T1 ]�]����H�hO6��$�%,��*c�P��]Z�j;�!�$�+��k&�@\�أ�"�!�d�X�𘃷�ɶ���[�aD!�d"x��8h��UD5���>i!��S00޴� ��1�� ���h�!�$<P_zE��IP�+u^!�d�Ԋ��3�E?�����F�?!�Dt�H89�,�/@�%�'�^!�_5K�YDd�6��1��M�!��!��0�@A�P^>���=�!�jN�L@Ӥ�����ض"� so!�ɛk��RGBڜ���0'�:a!�$� oĐqS`I�3x$�%\-k=ў ��S�W���°�Y(�C�mcVB�I�%���傑��
���;�NB�I�@Nt��AB����W�_�B��!~�6q���׈Y������و4A�B�	-�ڭZ�)[�6!V<` K����C�I93�0oH:l޹zd�4p
�C�A��p#P&]мٶ��B�	�I�`4��鋾9��@ �H(m~�B�ɷ4PT1a�Hڵ��ȑD6�B�I������bO�0o�AB���G��B�I4N����L�g!�@� шg�~B�t#<��2��*/�1;�j�	ȡ�1���4�eW(��!%� =!�D�2|q���jS4��a��Y�3�!��̧6�ܙ1���<���bE!���Nu]Z
�\�Ή`� G��!�?;�@l�f���|���1�ڦ�!�݁i��Z�-J~��ic�l�05͡��Q�)p�h+vU$��U�v�ڶ�y����>��'oI/6(-��Һ�y�kݪ4��Y�6ƾB]};D 5�y������	 �F�j��q
�n��y
� ��&W�a�H��5�U�A�|1a�"O��t��1m1>ܲ�N��LiP"O��c��mlTp��(ٯU�R�"O�<#�e�ȸ�5N�7C��z�"O0T��E��B��f$� �ɿJ�!�DT$%c^a4��<�����E��x�!򤗶�0��$��Tfyq��$f�!�4g���TO�<L6]P����@}!�d�)B�5�g�(Z� `2��T!򤂶I��-a��9tVh�L�(p�!�ܟV����Bo�2}��ɻC�L3/!�6}A&u@�e�)9����Dى!!��O�g����`��0���J�$և!�$P�h��݊���V�~n㑘O!�$�=e���7ɒ�N��}��J�#E�!�$�i�z���>'�����}[!��JbX�D[7x��B�Q->!��C��ܒ�'� X���1$O&!�JnPJ�$��o�T`G�Չig�A�ȓU��1��^$x��ɱI��I�<ɇȓWr� ���9h�N`��Q(mB��ȓM�.}pc J�XwtX��v�`�ȓ|�R��D�9C!-XZ�e�R�<A�*L�e��S���1%}�T8&�v�<�j�`�؉�UD]�	�>�E	r�<	�'7�!H����,"sLq�<9􌑶dtvY�W股Xi�pP5�RA�<	t���:#��i-G�sS�{��Xz�<ѣDQ?y�5a!��t9��1�b�<��"��fb�i	��U��3�T�<)DF�i�a��v�� �ՠ%D���e�H&ġhMô��"D���ӈРm(�@蔅�%1�*l�s�?D� Z� ԫ�d@�ѭ�!�X�>D�h�`��Y>��P,��DN�K�0D� ���d���hB��,@�Ʃ:D��	d�٧Wo�����o�
����5D�`�"�q�V�*=��@@�G#�y��1S�L0���(@p�(<�!�ǆ|4��B�a2�LiE���B�!�˷wM�tB2��2<(.��W k}!�� �vL��Y
5�����C�y!�$ǆ��h��NAI�z`0�-�c�!�Ɓg9 ɒ���m�ȍ����J!�ו
$���^��h9Ԏ��'3!���^�0�� �U��(�[F@߬�!�$Xk�x��vT\͂Cm@�M�!�$U G~�Hւ�+��ղ����!��J�7�h�6�P�#iMbg���D!�ϴ$7>yCa+Z�Db0���]EJ!�$��N��P���R:�,e��	�Py�'Z�3|�@��EW�Y�e[����yR$�=8��-�7ї��}����y�7X�\,1&��#,h�ۦ�yrlˣA/U��[�v/&�J� 	1�y2f�Lj��S���n�u�r��yB��`�$y�D�i��ْ�׾�yrf�:�5͗L*R�Brj���y�+Q�{JL�KOBJ��yb*�!&�jP���=�lE2&���y�Ϸ@����qe��R�c�iK=�y�eJ�Fc��1���$@��I�`FM��y"`�l̀a��c�{��%�y"쒘RF�q��&�$��X��.��y
� T���̕e�8���� 4���:�"O@Q�$	�ld��I�\!�ܱ��"O�FҦ��s��P�(̐�"OHAɶ�M(
�"�c�+>b}� I�"O�*I4�p0�i?D}L��"O�������B�)�i�M�N��"O�Y�f�� .��*o�{Lf�0B"O��y����*kn8@�ę,Cl(�"O��	�
�
!��ːj[�,�w"O�:w&_0�< Rv��+<2"O�=���ј]8�o� RD�$"O��B�[L7��Q�;���2"O�4���4��P)� Z��x�4"Ob�)���;��GO�+G�6mI"Oa���� 0�5�? ��+U"OFY�S"%ά[��*\���0"Ox�:�/�X�hiH"��CF��CV"O�P�������&���p�"O�y��P�
8��iժA��QT"O���`�.k�8c�.7�|���"O��a,�z���U�{�HH �"O��	G*'4�ɃK�[C�!i�"O�$Fl�b��,��)Ϊ@�p�6"O±��>�\����,���"O���&զrGđ��O׳E�<Bp"O��C��}XF5 ��!���"O~a�)N q;&�2mÊx��IP�"Ot�	���^��+W��Q��s3"O�M2"(�	V��Mq
�4��i"OpX�- )#��,O�hhY��"O�-����!/o�,Ó�(f�ȃ "O�\�e�E�rp��C+D����"O
	{rB�-���A؁,;�!s6"O�Q��O#��"2c6JȀ��"O����ѱ_�����\�<�I2"OZx�".�?s����R#�/�T9�"O� !bO� ���ɗ��MH"O��PhFb4��S!,�@��"O  K���4�d�d�t�.�C"O�J�/é5�(���Zf�02�"OX].5	.��b.܍"f&l�����y���8�c%H��
�"�o���y�Ƒ�[p:}�1��,]���1�y����i�j�W*�(3�EM��yR��-N�d(E�݁K�\e!�M.�y�i �;خɱ���I_tQ�W)�9�ybؿG��!�46Ek�����V�y"��&e9FE�M�%�g�ָ�y�/{��ܞPeF�'kP=�y����pm����(���1vn��y�OZ/AEv)"pdZ��� �#�:�y⥙!s�怊I]�:������#�y"��4��hggL�GWz%#�š�y���L��{&b�27��"$�(�y
�e@X7�NZ�}y�,Z��y2�� &��mC��@%K�FT���y"�ҽ ��A��PK
�,� (���y���L�\I5cD�Nh�y8 j���yR�5x�̱"�Kلl�JG��yR�Av�<����{ify��GQ��yۀN��i��j�l�4M��H[��y�OV13q��P-h���쏹�y2c#Hr�ЁaA^�X0*|�����yB�I�Ѩ��'ծ��Fl=�y
� �8i#i�U暹c�B,��͡1"Ob����T�JzY��C��U��"O�t�rNԔ}��������p��"OB��vOתSK�+t�A�X�jE"O���$M�
�~h�����p�I�"O2�-�t9��+��1=��)�"O6ձ���_����[�#�dٲ"OĤ
7wx�� ��ƋmUZ���"O�im��d��a�N�p��"O�]`�#0D�JQ���/`K��[B"O�ԃqdZ�<��1��Ȇ`n�y"Oz}ab�ӏe�� 3A	�f��!yA"OZ�L�m��=	rV!:��,"O�L�6M	 L�RAi��4~��� t"O�m�0KF7}A��j�:�f��"O�` �^'%����	���H��"Oj�S�<��	��F�T�0�k1"OحB��x����%_�^Z4( "O��X�Ǔ�dI��D�!iJ!r�"O(0bi^c�L�҂�>8/Ԍ�@"O���R5I��JA�ۄ`;�1Xv"OVPJ������j�똦h�� ��"O�l��jY�R?@�I4��<�>�sq"O4���\bB��������D"OXd{#*P �0��7�ߢ��y{!��֓=&VZ�� �I-C3jǭJf!�d�<6��H �H�rFv�bEfT�g�!�DL��|��I&&�n iÇZ"2�!�ӵ	��@��`�)�F(�a��j!�M�B�rS���d&� ;�*1\!�Į�t� Ӈ�'1"��CJD�n*!��D�l�^�z$j�<(��K�"!�� pƠ�E�	�S:�p0���*!��F�W�$� �A0!~��*΀D�!��Y�2�0��cK�HxN%O�K�!�$լ#�`�=qvĝbPNP�>����S����E�N;k,LiuGͱ�y��'y�^]i3�V12��w��-�y�Z�N(r�Q�&->��dK2���y2)ǂsID�b\�m�Z	�Qc���yr
�	h����cݧ|6Ĥ��g���y�+ݗf(�Z�'^�G��q�L�y"N�#X�.���'*iR9�p�Ӌ�y¥��%N(j�A̠!�IТ^�y�@�p��4��fL�˦)ig���y�˓J%�}8�Γ�1�����J^�y���6�j`��N&)�V�xa�^��yҡιm�0P3C'DdZtBQo��y%H�Q�Li)1;xXZ��AG��y�ڟW�9(�D�AxN]�0F�yB��9�t�卉@N���F[��y�ʖ2w�ri�I�mRRpc �Y4�yRɕ�Q���⍘b2�Q�fL�y�uvNt�������^��yRi[���#��j��9�ã���y��9�Bq��D�\�����"!�y��ů<�F=��H&N��9�cf�%�yR�F&�骣�B�1�ְ��	�yr���(TH�JGb�<����%D��y�.J�D�4e�lH�gz�����y��V�,d��V��'g�h%2��	�yB�]�W4|iJʌa��M�����y2��G��j�N�	��%)����yB��� g֑�юŕO�"��>�y
� . ���=��%(	Y�7&f� G"O�<@�V%�]���a%B��"O�Z�� �1sp��숝C1ht�S"O��pIT,rv�5��D�9Hq �"O��Q��=l��	�� �Oh���V"OXx!��ڎJ�P�R	GO���"O�t����7[l)IW)˲@9����"O��(�F��N�� "���l+��p"O2x�`�m�T��K�~��"O���fHw��ffժ9q\8B"Oޜ붴�z�N�X�Dؼ\l"s�"O��04��
j4F�{aFA�"O>��J��6#ҹ�ɔ�R`(I2%"Ot�IȕZ���z��)<��	%"O�e�,�C���QDf�$94Tx�"OT��`'!8�Z�$(3�(6"O�M �<�%��2�iP���y�8xҴ#�D
�
��p�]��y"MP�����d���O�y��BKrI���p�1F`#�y2ψ�+�d-�� �J&4���F��yb��
W�a�>+��
F�y�΀������I3fµ:�ߨ�y�e��J�A�A��&����QLW��y��%�j�R
�� �~@�Pʑ��y�/�2r 2|1�X��� c��'�y��G��xaЁO ��(����yB���0�U�6(TCK�a��"ם�y��X�Vi�2���5oȭ3��(�yb��ېE��MǞ~{f$�@��yr��4fxv3D�D�y�N���h
�y�@X9{�0�Q��w� �YR���yB�*Xal��W�g�.xĬM�yB��:C�Yx��)d��4#WJ �yC��#|��	`CɌY_"�Z��ו�yrO�<~��Ȃ1b�>cx�Ɗ	�y"^iR, Rs#D�6<J	`�e��y��A�ZᚢA�d�z��5�:�yB��p��U���(O\�<�"���y"%W�Xft��F�!F�1����y��Ր&K@�з ȏv�����g��y2��z�(�����P�R�ϊ�yb �<&Ҝ�2��C���T:�'1�y� H ��}��Iږ7���rJ_4�y��V%^��H�!í(#�9
�e�/�y"c�p�m��H�=R� ��C�N+�y*	<('J8#��]X��5��fļ�y�B�.}+�@p �ȨZKH4h��֒�y��1b�m�-M��#CC��yR��k����c�FZ^�!r���y�$I����M�@h��h��y�o.'����"8d�$��hJ�y�cR1��@���K�gs�������yR�<d��0��R	W�F���Ϭ�y"��&�Ђ�������yR��C��@�#��|p�[�I��y��
��<�� ;{U��ÔǕ7�y��P�\Xb�o��t+��[��ּ�yR���u�x� ��>f&8	D�	�y��-4^N�2� �[g���S���yB͑:;� ��rC�	��y˃�H)�yR�ɑb�TŲ�*H;S!~�R����y�	�I�ᚵA�b��;�����yb��$pT�}��ᖃ[Q�ͻ����y
� �Ͳ���W�4��a��.���G"O,-��Ȅ�q'<�	�ڝ*��\� "O� �ݮ	�����"p���"O�qA�����r%+U�-�(D�&"O:�ؖ��J>�5u�ƂN�82P"O�X���J s/�� ��׍8����7"O�s��E+b�d	B۞.��ɹA"O�@s�l�
A�d�P�E��Q-�yR��l��%�@�t�Zyõ����y2�ˈRT��6�IhEJ�30˒��y��>B�=h�Q�[�}+@W=�y��4-���d��C7�,P�	*�y�l�z�0qVaPw����J��y"�¶2�)YN�?=��Z��ղ�y��E
9r-"�h�6W��Bk�%�y2M۴�� �Sk��]7ƭ��@��y $Y�zUC��X!V��f�]��y��>n9�5�"j6]�h1�H2�yr�W&����q �_� �:��N�y��T�@�~0r��^���������y�a\p�Ǆ�,��yh�A�y�C
-�vp������������y��۰A�ʔ�uED�T���k��ye 7�H��3柲RL8;����y�2]����a>O�Ƙ0qi���yr�3�MҦ"�	H��{�g�yb��
n���[B�Ȫ<�B���'�yB-��PPq*Ġ��5��k � �y�g\%<!2����|��"����y2�B `��(x�A ~4�P'��yR�[�(��2��]�*39�!K���y�!�"6�:E�����raK��y�E׸'�Աc1���ȑs�'���yRA!3�d���F,sF�q���y��G�=f͐2��y(v	��	!�y2G����Qi��C�o$8�	_�yr�8N����+gJ�@c�y�
$FTy��JE�-�1 vIX'�yR��c
� �0!L88Dڀb���yrX�xX���KL(��1��e���y����z4$��ـ��9����+�y"��n�d��gI��"<��eZ��y�&}"�XjBhPil�W�B��yRL�Z, R�C��z���7E[��y#J�]n�C"ph�AP��y�k��m���ч��X�4�]��yϏ�h?@��cϖ,�l��-\�y2�
0��Z�ˈ+!�|ɸ4M��y�$S�O���{��).�%��i\-�y�iR�(r� qW�HT�����y�N%2��1�`���@�H��y�fΒU�x�bg# %]�ش��3�yKC�a	
����&��E�,!�y2K��2�r�퇨� ����R�yRo��L�L��Ĕ$+�X�)��y��2�p�V	I�TtlǏn� B�ɣ;�\���+�{�T|{���&4��C䉁#�h0�F�,�I�q��8]��C�	�2w�蹅ϑe� [���^��B䉈?b�I	�"J�n��p��n�#�B�	�Qr�h9u ¤/Ȍ,9c�B���C�	�����e��&Hpd�T��90��d�+"R�{�n�<���o��J1!�ƻe�3�@
} �����P�!�� �E��>U��-S!AQ'@�X��p"O����$�	e!�=�1��_ք|Ӣ"Oj���5�D����Hb�P�e�|��' ��El�TF	'`4!�4�@��,sr��k�ɂ�	h�!@`���y"ǌ�]�]	�[L�d�ǌՆ�0<y���:h0t�֒��\b��.�!�d؍j��S#@=G�JmZ�nV�O!��2yx��#�
6�~D��G�D�!�d�{H��Z����y��S,]X!���q�L�����h��mFGE�'Aўb?	�юǉ��� E��	~3���_h<9��H�4�r���U��PkAk�G�<��d�J�:�A0�B�. p�+�,�z�	h���ĎٱE��W�fdiz�6�O���.\��ಃط<nZ��f(+A�C��㦩ɐ���4�ƴKbD�%h��(��E0D��E�4R�za��&Չp��(�p�+D�P�V�,x9I$˒�X�$�*�$q�|G{J?�PED	r�}@qn��H�De*g�'}Q���<A�}�o�%yM���i�/5F��w�ѡ�y'��A?n�J6�6� h�����0>�M>�A�um�-ۤꔘ�^��cO�<���7-j�bMM�YZp�ɡ�Q�'Y�"=�O������.Lʔ�р	��16� 
Ǔ�HOF�B��/J0���RSx�k"Oz�)q�F�tXBYcb���zm�L�AiM������N�F��!�A��
  �ō(:�!�DF�d��\��U'bP���2�-�I&�O2����5T�}�ճ��ݸ5��D8��'���fd�2!|�#�G)hyy�"Oz�dh��G����ר��\ZX�'"O�9r�>%5�]q�^8��m���>��'�0#=��t�ҵ�8��mp�)��ȅ���'\�ɏl�L �d�ʔ]@��@��RS��=�	ÓU@��n����D�*�2��� |�,����Z*�=1*�#o���	p<Yu� j���g%jvpZ��KB؞$�=�1b	�C�P��&D���:$̃|�IV���O�$�z]j�q�#�/K6��yyґ�$��|�"�_"�a� ��*��ځ�K�ð=��O�-���x��TW:�ك T�ɠ��WF��c���f��٢���g��=�ѕ�(��	U}�j�
�;5d٧[�$�J�Ș��0<14k9ʓ$��3 �?&q������4Ё��/֕*�@�>���˰�	/@ֺU�ȓP�<�i�=�$X��g�9�ȓ5 ��0���ph�iC�!Ζ �=ۓm�r�XvC���^�z�l�J̅ȓ+�~���%X�6(<2�kQT��	s?���A�
��ō�>O�9���~!�d�{�:�R2F0{�����O�V�!���!5R�̳3��4&Ղ�ꣀ&cz!�d�O`�4�Kj��m��,Ԣ1W�����.}��)�S%O���u+�8,�P}��d�?����#��6�\��o��Q���֬D۱O~��6O�����Ҽh>ha#JI#Z�~9q��!|OX&H�#5�$���~��i��i����^R�>��B'�5=�T��G��g}azB!p�@�OfT9�^�?���WIQD�D�f"OB��L�m��$����3zt��O�|��d�XIaJ�"}��E��@P�f��s0�
P�U�O8��S�p	㖋ӆ���zpd?0��'y�	u�\��؈_d��PF[/?�L�1C�"��ȟ� f��� n&��-�XA�Y�"O���Wf�F�)���ݜ5AF+��'��&��֧����/.��� 3	��ɪ�\��!�13M�,ia/J=���J6�A|t��0?�VNL�d��6W+���תY��y���%!�cr�!��Pe�y�'�95�$�W��4R܁ ,ز�?�B��<�a�
�a.�`��+K�! �]�<��!�-\̈�`�I&&��P�&e��<)M���'Ή��-�D� 0�Z25�l9z����@�ē-=��1
D<$ ���@��$wLp���Ԇ�I�2��y��]�9���4��'*$@���4�!�B�3���Ӟ�`�m�t��#�O6,��_6y�X�+͂�����|��i�)$�1�(A7$-b��� e$��*��!D�`l2�"���V�8��A!<O���x�IL���ළ�T��5��m�xɘ���O����w
�]"�aCz�<%�$#� T?!�DVu��J�"D�R�<y��;'!�D��]԰u:�mY}��ܺqBϏx!�d�3>n(#@�Ӊu�8�c��J�!�d%e�DQ�Uc�����	�a[�B�Ih���ԋ\�@j0"�)w�B�	*'���V
1x���Su�؄}|B�I�I��S6-���
�־%�"����I@�}rv K��v0'�t�B�	��(aOΤG}>m�6*�&C��~����	*� ��,?�"]�#�Z�QV����)
rH�{ ���FJ�1�C6]�nݐ"On��‖B@��� �������,�S�'t��6䛪7�(Ir��n���Ѭ�`$\Y��ɤ��t��t�ȓ`����$!p��d���F��.��ȓSh�ifiM<w�t���O&PQ�P�ȓ���0��ܒ,|fHڤ�� �F��ȓ	�xae�خg�T��ۄc�^��ȓ"��UP5T��
����ȓ;7`��V�G]�L�B��!r)�9��(�h	f�I_4�#1�� p6��ȓP�`T0ơE,�ҵ�#b��v��ȓ\��k��пN2*�ӶX&,�ȓv�
�{ā�$ ��ؑ���4�Їȓt$@��5�N�'�H�	��d	]�ȓm[�`�C�B/R���Ɗ+G^!��~f����msd����#�����/�(lZ���<�Ԭj���;\(JD��	�	YW�G�h��� j�Py����	�
�?0QҜ�q��݆��ȓ1�����Q3<(I��"�;6�l��^I.��(�h=���J9:�N���K�P���Si:R�Q�,
�,��6�v�ŌyO^,A烃��R��ȓD#�� �-[A��"s\:�ti�ȓUn��LE$ot ��3oЍI��4��,mp|��ҡ���Rŏ�Ȱ��u=��A�k��i�Z�b��L	;)f�ȓZ�<�d��Qؒ�b��S�O0��ȓ<�BdzS�ΓG��Z'L�?,Ђ���S����3�E�
[m��8�����$3d�� �Q/�1����d�"���A��d �n�/%Қ��a$�z1�)���`S��Em4��p͊Pv�х�O ��qn�^��`���ЕVjͅ�9e�I
ԉ�/j-˲G�u�����S�? ���g݌[҅P4��^>F��S"O��d���5�JU��h
�F!���"O�|�	׹H[�I��G��L�3C"O
�y��(,80P�6�;ti�"OPek�	D�6d�y)rE�8��*$"O~]�A�[ ��$aӪS�>Ͳ��V"OF��$�M ���&�8A����"OF�ӓ ��<���X
%�����"OD:t�E?^܂h��D�-��Xc�"O~��sc�'m�tL1R#$\}��r0"O*K7*��82by ��]�3xJ"Ob8:��J�W\L-��kƴ~ ��c"O�+u�L�M�ހ"D�I�0��pq"O"�d�C����*�,L�L$Z�"O`4���]>��|��jQ�p�b���"OVhroE���T"���4���r�*OЋs,ƮLT�द�7PD�A�'���*��p�p
��E�����y�HʾH��ā��G+{�d���y-H�c�4h1B@D=8?$�Q��R��yrfN:c+�`�a��0��m��*I�yB.��<��`�S�� i�DӁ�>�y��A�_��(��Hk�D4�ц�yR��%>���b��`bb��y��Uj-��2���$٫c ���y銾ٸ�C����۞4ʂLU��y"�Ԓs��*��Ƒ1!�E��y�KE耡�ك� �T��y�툋&��ijw#��
��p�Ĝ�yF��r�E�8�b8�b1�y"L�Nv:�q)�&-�ޕ��Y��y"+Fj����,;6�:tV��y��;�����3!�5�����y� މ^E�X
�lƨJL�Ks&��y����)�TN;JҠ
�	�y�M�,�~����4K��8B�F��y"cY��qhU����( ��V�"=�)����0?AuM�AZ�tK�5�mh!�f�<�b�E3���I��@�}�*9h5.If�<�C'�8ǌ�+�)s�z�@�TY�<)S�$�&d�P(W�Q7���x�<��B�;<����`�.Zќ��p�<��Ɉ_c� +#�4�b��e�o�<�qh�V�2a�!�t��I��G�<���q�z�n\
�~��]}�<i�JTGzڕ2��, �2�(c��z�<aw��D���Շ�"}�9AP.Vh�<ْ�M�7���u�HH�C5IIP�<�#�����SԤ_4PAd�9�f�<I�)݃U��f�6�Ȅ��BYh�<����_'ni���^�0��bʊo�<���E37�L�R c�.<Q��NN�<�W"��u����Z�
�o�K�<�4�*L�b�(�v������@�<)6� a2�)��*Hx6q��jU~�<9v	�D_~���Փ}|6���At�<�AF�H�`��Gg�	m���Z��V[�<�b�̋'�!���ڏ}R�rׄ�h�<1���6:��B#�G�� ��Q�<1��իY�dX�
^!v0|uGL�<�AB	�%�A(�E�� rs��H�<)�)�M�uQ�`j�V����M�<�d��&�Ќ�t���s��(�b/�a�<qǄJ�V>4� �]�4ա�QX�<� ���T���"⎵q���*i�E��"Oܪ���/�"�$U�%�����"O���'�RBi�SMۻ9� �(w"Ol���M�u����ׁ'���S�"O��3�ƎM$�,sW�Hm6���"Oư���\�4֘����L:o���"Ot��Ș
 ���&�Z 3�Х0"O�Ae�J�@�B�"%�/=吴�"O@������.��eQ�NK���"O�����F.B�nd3Bb�"�i�"O��CЉƢ԰����J���Ya"O ph�-ϼ@�r�b�`����`��"Ob\��e�u,�X��9f���;a"O-)B�H��S�� a,���"O\��A��
"�`$i4(E��(��I{^P��鞗pU�8��J@ ZX"�)ڈ^=!�G���x��g	�1�ؕ"!hO�q(�䓽>N����4��,j�� �H�<���� �B��!5���ٴ/�>a(������J�}�Z<��Ъ=;b������S�M`X�<�'hF+<;a~#���L�h'���x��eپ#�h���b�Z�D%��O�ڸ��M�'x��xб+�.!�&�F|�)�r���t��]ܧu�D�SȊ3�ڠr���$ ��Oo(��Ԃ0�(3υ, �rEΓotF�0��1�Xҧ��6�HB�FY�\5�I?.J=x7"O���ġJ�c��X��P:�j���(���Ȇ3�h���'�6�Hp�əK;6��A��Bؔ� h� RIG -b!�C!��O�X�6ǒ�Gr�D�b6�|�ʟ#>����`ញ;�R�SU�>�/^\�K��W�.�>�;C�#���Q0Ü^ f5�ã+D�8aU*	�4 y!梘z6~}���@�AhK����'��}����p��Œ���//�z�ƢA�<���)D�(Ɔ�:wEإYt�?�'t쎸C�|Ŏ�[���\��	�����ȓm|s��� =�)P�MA<6<��ȓ.��,��в�n��C(G�`�FȆȓ#v�(��-�*7�Ũ�"�*��&�D��+Bf0�qk܊&���ȓdJ2<�M�"6a�� E�X���I1ːlh�Q8�$�!'=@o �`  H&>��]
ˢQ���I�t�t���p2Q�����Z�:����~³�,�0 '�X��f8�%G�N�<���]���L�PL�G��`1v/ �<��LM��pY��/}��)μ#^�Ah�ZG�dK�ō!�DH�1�$da��2;��{ф�.L��Icf��W���_��x�逮]opx00-���fY�����~���h���X�6&���q�P��bY	AL(N�\�+2'Śh���j"CL��z�f�<"��� S%İk_:X����С� (J(%�DL���u�'Y4@�'�ک�}b &Q-h�DRD!4d�5Yv�K���i��k�L���<���K� Ę���)Q�&q�����]%ug��˰#�6,��Dܛ8$�e2׆���)�:l\�1��d�+hQ5� ��!a��cv�@���%ЁJ�<BF+�:e�����k��~rb��x�d��T�=:�H�G������
�x| ���O \JX@c�^�}����O��W�LU��Gtpn��W02�n�4^=`tw��td� ��,bl��P ���l���`pa��10w�5{ӣU�_�.aؑO�y�O�S@������S=`▣��vI�}afN�!�Э1 C!k>`�Dy�CtL�mqv����!Kv̎���&��+�+O�%Rf�Z@�P�lL�l�Z��'P4�O0�A��.B�'�v�˕�2c�$q�O�5I���.̸���3`���QMC�8̂�QSdXӦ����	�\ႃ,I0O�H��-�Z����.:�Q>�	����h4�SWV�sr��38�=��,}5�9��4��c�| u	f2p�s���.���A�R�N�XF�W�t��Z�L1O8�+��Ll���PiO3R[8���'�� �dF�
��<�O�'=�@y�4�#��0J�a@�y<��'i"~�̝c���fB቏~T�0�&��O�4,�E�4{L�ʓ64�����8��99�㟕/�A+Ac�<���>�)�H�f<��
��RT0q��'+��p��Oƀ ��x���&s���`�>�N�*�C94���"��4²ر�E�!��=���'�,�iX+�'`�Ҥ�Yk���� �3�L%��{2�A��{�'�,*� ���	YU�Es�'��C��;/�4�燓�a���		�'�:E!��Uy�h[���.	�A��� I4&y�rh�+�(�&���K�ۖLc����G	 MXb"O�$!��	˦��ELɀ8�D�Ɗ�3�@���J�_Ŗ�I8�H����N�ap��o�|����_
[��B�	- ��$@�"��T�$%R�H�7$��
��&.�-b�#w�bpK
���£Gр#,�t���C**��I�;�b�Ȱ#D	;L�2`�E�)��5��&w8dP ��+\`��vw�!�v
�)eI&�������S�J![�@4ꈀ`��?ǀl�)Բ$@S� .�&"�H*�x"��y��x�.~��[5d�u��Q;�IQ�/�`� c��e[��hEkB4af�9�B@�$:x`օ�W�&L&�R�g~��=٢9 �[���������'4��e��
9}�Y	" \wܧ=¸,c`�3>8D�gjU!#x�-q�32&�s���|�F	�'^��0<�g�(�$� �H�8j$��G��'#|֠���̐蜼���O:�'$�y�g�Pa��d�R�h��?H6�R$D��e��dD�Xf�L��ɼRNB}9sD*)22I+�f�L�d�0�\���R�$���!�N��UC^EQSh��,> q`ZMj��'l�xȪc�A,W�͉!�E>���I�x�)$@�k�l���jǲ ���©��;��A�U���[�`{ ���%�³�_#����Z>uz�HN�Tt��'���Y�$2a7̄jč�({2܍�B�F�to^�is�Ha�d��O3ؙ+C��V*�#!*C�6��H�L b�����a��&�����2� (B&��/,""?��B���%�S/���yK4
�c�>���,� ?��Q���O�K!u������U+�Z�d�:�r�E˟Gy U���E>�8{Uo�0U��Q��'�(�8&NY$B����\�����o�D���1�C�]�R��F��f�uzܴ42B`@��_h��׍X��@aa�@-s���d�¬�0>�å��)n���kƬp�����-��^%j1�Ԏҡ4>�3'j�?8���uB�L� -R���0���Y�&�����N}���D��� ˀ�H�Q3���(Oj9�����E����Ob�Z���p�v�#̱9Y���G/lOH} ���:v��%�J�t��dC�xD~�-Ľ{��ѠB�s�h�KI:͈O����OS8Z�H n\�Kx5q���y�ܠ��	�8\,���ܵ0?Ը;0jMi�2��ě�L���f���2�@"�<�~R��4~� � �I��`\�ٴm�cXY���S�՘O�.Yr W8A�0hC��	9���'7����#�C�̲6�^�y V��T
�?:�$,��o8���g��,��)��Z�r�OΩ@��?�= $&êO�d��'|��s�ū�N��Q�Q�9�~���\�%�T�X�ԛ���c��(�����-d� ��Q��g��=�C���t�>I��� �@p�'uR<�Am��?9����EL��*�nV�?R�	�.8D��@C'^��ҤI�bU��,�>�����$�"}z�"Q�T5jI���t(�4ʄi�<Y�Cϸ>
�i(/T'G
n5��X�<�R�X?E<L��a�fF���M�<)�KT7�b�+�1�(��N�<A�*�b��_�"yn4��O�<YT+�7�,yv+,��0�eFH�<��>h ���03ފ���F�<�QE��U�\"���)�{(LZ�<q���6\N,�x���&w�0=��V�<��(�Z��D�!	�533\��%QJ�<��̉=S[@���Źe�����bs�<�'�
�X� ���G#&v�li��An�<� +�008�D�@N�P�ԏg�<�A�T�M�����/EAtv�9q�]�<�#O�/6z�x%��VYf�z�jq�<f�qMd(��O��0��F*�Z�<)�ȏ
�<p�'�¦yfBi�P�<��Ij��Щ�A�:�i87m�S�<)ǬQ�>�0�$=Ŋ�#@��G�<�&�>[PHRP���8L�TgUz�<���
�r��K����J�z��"�u�<�0B��6 <9&l# {L$�HMj�<�&��&w]���U��+[���rӫWf�<� \L�'M'>���1���d���j�"O�X�%	<�*��#Ǵ�{7"O��cB�BeGr��4M\�7�yZR"O,�K5m���� uCӛ)����C"O��9�`˼���2蟕k�ȩ�u"OH���]�JS��x�����؂"O�9�8ў� � W�O�:�b7"O�����V�(����0�M�I���%"Od��V�W�v)��nK&o�H�9b"O0��B�i��9b�ą
�ZBA!��YT"d$�n���2G��!�0.�:�BH�'/�	�,�KR!�D8Ud,���U��I�I݇H!�Ӹ$|��H0g��K�-"eJ�hK!�D�.d\�B[�k�����<5!�d��8�¹��C��}��Bw$!�D�|�x�֣Ёg�\}�7�	�!�$W�C�у@�Ⱥ`�z1��R( r!�H�fv�:苄Yy���iQ+!���8� �`�\�N&�S��!c!��)#s��C8-��bE�&�!��?;��-�GϘ;l;p�4!��!�Ė�3]�!�Ë_�f��`��Ɣl�!�d�RU�@�NZ� ��؍W!���7 �nуC.��c�~�b�� }!�$ݓB��D�g�I/���J*	?K!��>�&}c=`w,"��[�(A!�D�]:z���Fɯ�܀�0BĪ6\!���b��8�'�K!�ܘQ�H.;�!��:l�d��L �ĘA�D<!�䖅52��H���S궘�"�:t�!����Vp����<Є8cs޻5�!�$Զh����CDװ4�@E0��' �!�h�z��Mרw��u�Ua�<!�d� �8|�"R$^V�A��!�x)!��
�?ڍR�B׿hL)�P �.+!�[�X����(�UBP	[��. !�D|r,e*U��h���2/��!���^a�R�v�<e���ʻi!�d�*B센A�/�:C� �H�#Y�}o!�W��9{%�T��y�Ul^[!��ގ\i�\�1aP�gߜ��L�Tg!��W�%4&��[	��9K�`S�Q����ȓUI^X�4-��tOؽ��H��!��������珌�4�θ�V�>V� ��Uڢ��0��jj�G����l��h�zG�ʌQ�����AI�|���jT� �¯Oq��ˑ_d��4T<�ç@|��I#�*k)��ȓ/����f#�/� ]���V�R6����yP�9�e
P����
@��@���:��MN�GO0�*�O�z��؇ȓ���b���G`$E�Kԗ�\��8�.�r��O�c��ju�V(����ȓu�=arh�&a�� ��ȉJ��}����5�S-N�3i�����m�]�ȓo��1,C����Td_./{T��ȓ?�@�G�I�j�T�S�ȅȓ���'�$����'��6�R	�ȓ8 ��L�0�tH����	P����yK\8���K�|7�� ���L�r��4Ұ}"Wo/"X�D��L̀n�< �ȓ_!ZDPc��Lqt�q�lI'>��ȓe����#eW
�g�c�z���S�? l�2�oӥ#
�x�(���:���"OR S�F� O|n��ǃP���8�"O�$��&?:*��,�>��XP�"O�����"$;�q@�5<�<uh�"O�袁"�|�J��eH���HBb"O�MD��N�Q[�g�)OD%�6"O4B�,`�ڰS�#���(V"O�4��]&y�XH�V7JtnT�B"O�L�'�O�:s"i��A.`S�pj�"OJ=�ƣq�n�)���r$�Q��"O<}�D�R:��R�a��9�"O601��0@�L�0U ��Y���˔*O�5
��Z�K?�]�'bË_~,���'��y��I>RZ��(�ƒM���'�����F��Ħ��\:F,x3�'��:p������T�\��xB�3D�d9�'892����h�C��g>�B�I&7�<M�e J�hxX�� ��WdVC�
>�Εs!S�-Rt WF֝W�#?AV��	���?��0�R�R�B�!�ž�r�(�D+D���Ƈ�@�0!�C�Y�R�H��m���Ʃ���^�&��}b"�C�Ġc��B�N>�xzӫ]f�<i� ǭF�-RcE�Z)y�� ^~�h��)�\ ²�Y@8����a��x���yg&�O�,��c��&�9��K�-�صҐ�3r<�������Px��V�pG2I�g�*%4.y������OZɒ�nI%/��B�����25���0Ek��t8 �͔�y˭r���s�#�*6ܪT���y��>b4̙r�@m��8�&h�2�P	%:�i@+��GˬC��&��l��▖0���0���%ɾ�,dr5C���mN�����,6�@DH�`[�<�
Dٰ$=v�a~��:u]r��%fΚV�V�zc�M{�)8��K<`d�LeBUR"�/+j,��q@6+NDD|���I�N��5�Eܧ{��A0�e�����u(�,jp%��l.p+�ȥ<�1Q&���0'���oF&�I�	���S�Oq�Ȣ��A/x�X1�ѥP��@��'����4�*�h�'5��q�K<��"�"k���D��X�D��S� Tx��R��Py���<�� 3��)J��T�����y�ۆ6L�0z��^~B5Z�ꑌ�y��^-|,�i�D��W1hY���y�/B�|�ӗ'��YC���"F�y�K�� .��acޤ[䀤�Ƈ2�?Y&�8vN��P����j��h��H��44�����&])�	�c�����$8�:/(y��B���Oܴ��#jт��3�ȏ�p}`	�'�2$��Nޱ3
��s ��~��)��'��	���>��O?M� �E�C�g�C��f-��$D����3a�j8����V�T�K!?a��XF�(�2�a6Oz)ai,Q�٠�2V���S��Ob��"��7���%<ғ)䚕�e��p{�	y�A��(V�D9#���h�0�G8\O�@S��F)X'��9v�[�ti��@�N�nw����з��C��d��wcě���O|Л�K�	a��k�Ek}�\�O�P������4/By�z��S�L�xnr�?�rU���-�q��%k�n��{���@�1�@��>�|��X�P�"�WB��2��-�&/��G�l��$�r#��x��Z�j�V 94K�` ���OZ�C���q[h� T���PŐ�؂!�K/ d�1����w��%BB�����?�����1Z���I�0|�D;���O(�)E�3�j �I�6P��#<�&��>0�4H�V��P�1ҥ���%b�C�ݢh�J�0aE�!Xp�Px�>�O��钠*s���Ru#	 D��1Be ��q�/�#S�h$剁G�ENR����vN�$�my�@Վ1dL�'�^3te� P>N���e�##㖭�é�AU�C�L�to	�.�E���1Gָ�R�H���0$1�{J?y�|G��@�˂:0F�(���-���е��D�<�#�c�fR�"1hȟ(h�峟�	ѧă&�&�h��5r�^�bh#ړfL�I1 4J3b?�ҥ�<0�p��̌�&Y<��� �O\�+i��Z���P�%C8KB��� �]0��ļ#��1�%�?xӔi04�'x@�{�h�1{]z��O�'��Y{�AP�jF��#�vն5i��v`��٦C�> C�Iu�F�	�T��[F/�4Q�vZi�C��<*�La��2Qh��pA��<I���X��O4�8 ��[x����'��h�׏�#؂}��㐳	Q��(��L�4�Ր�O����/��T��ҥ~\P�k��I�Q�����S�Q@ ��%G.wv�<���ƅ
�nC�	S��C�%B!V��ôeG]�`B䉠Y�p �5j��'X���d�&y��B�	!�&�\�(	�5�	�r >]a"Or0���X*[z�dsŃ�#21z�"O$�"�P�H���%�+7�u��"O`t�띈טIW��,?�X0�"O��CTn@:�h�ۡsj�b�"O���r�88UЩ�AθM�F2�"O8쁔`O�].��f��2��*r"O
����߼4C��΄�4�͉��O�	ҭ?t$���ea�M+3��f��P+���6;�!��	9u��A��32ĢГ�̄ �����c�F���F��Ah<��#�4h@��%�d`v	�F�c#(��%�oޘ�%�+��/)��i{-�o�PQRbݏm���9��G6A�ax2�R�yӊ�Y!�A�zIV�r�F��U"�ɗ활���$���F��J@�8���I*���S�$�q����LϞF""���_r��yw���P0�����;�'	r�f�K���Hy����8K�cd+\����'p&�Kw�܁cb�YqB��;|fe�1�'vP}��W��8�쀇��p���NH�x;q�F;�p���v]2b&��22�ӧu��6�D���^��a�熽��!٦a�&u���ҥ�8���X��,�(�}��k�]?���$؝E|b<s�cB�p4(D����

{�8�2h�|�.&ā"$J�#�#?	t�tW��%�OJ�|a��ıB�IץI#Y��HЄ�O��`bӞ<�e�+�D�>
B�	���[��� �GA�,��|��$2\[~��D�:�X2���
1'P���'��¾i���
�F
9��I�'�PRE�inN��c���s6���*�B7
�#}�Z�!`CX��s�jN�,� �B���A�:��L9��-!�]�'�ɦ��
qje�O<����ڨO�a1�]w
�P�GȻ(Ϭ����-M��i��v�	�Y�ֹ��"�+|�i˅�s�h"�@�A��rᗟ��*A+
��1H��IY��YA�E��Iz,�c��%�">�r0-� )`	/}�֠g�*1��.I�9�p� �7#׮T�!�H���O��~c�T�鍝2�(E*2
��yƈ�k���y#*�d�d��k�4��C��kR�l���0R��A�R�Hs!�䈈3jF�@b`V�
g&� pCS�Kx�I��d������x�mU� ��}�1���(��U�����0?q�J �m��X��:n��Y�aD��f��P97z>Bቍ,�y���o�pp��@_�b��>���Ѷ����O��j�`9�R���`W��yBÖ#*u脙�nݣ�X�����Lt�X�{���!E���D
P�O"����!�D(g�h1�s���2(���$7�!��U%� 0#�����Z��&��!�dޡҒ�SPI��� @��� �!򄟛Q�-k�(�/C���a��M#;�!���:[�Np� M+{�4Z�&��E�!�$�?�  ����E�U��Z����
�'����*h��u����1Pm�u�	�'�P�Chyu�tx��$�$�q	�'�> ��;I>�-т�	 ���'M�sc^*��l�!����h�'�r�3D+�2T�~�H& ��Zn�`0�'�����2�0�zfH��Wg�Ԛ
�'��{�Z�9�0E
�[�,z
�'����dh���^	?�r��bB�yB�[]�,���۪6�n�9�@ �y���f�M(��A,��@c����yr��@Z�=��A�&it$IJV\!�y",ĒG��XV�	d	xDYv�X�y
� bt���ҭi��X-XY"O0��L�?6��Q�B�v��7"Oj��7fM�j��@���r���"O���Vj8�(��I3x�<�"O�����<���6e")\q� "O�c%%��F8��:0��<$�b"O�X�N�"�����Gϼᠵx"O�q)�鎳k�`C�f�$Ѵ�ك"O~���_O�D	�0
Ȥ]�"OJ���Ɏ�J��b�	�d���"O��J�J�@����a��TWJd��"O��0��T���
)ڮW>���"O��*%@i��!�+E�HC�!�d��.���ĕ�iQ�AQ�D+0�!��VF�����L�Xs��q�(̟�!򄝄sk�1+�E_�\�H��	9u�!�dX�j� �F��FY�H-��L�!�D�<akӨ�)0Zh0���TY!��Ӂ]i��q�O��/� �"ξ:�!�$,g��!�	JՖy(s X�5!򤛥����F�H���3� �4�!�\(��9Q��� ��oɚ*�!򄓈aW^}���7�,�s��Ɓn�!�ժ�N%0A��2p	(�m݆*�!�D�N�ژ��(ݸ��ek�В !�I&"���rW�=k�Xd�G��4�!�ğ-��܊�ߟ
��f߈(�!�d�M��Xa�$l�8��GŒ+8!�J`/:�8�d[�d�u��@�J!�l� �X�.�:?[�50$���+!��&F��(�p-oT��$ˤ^�!��<_����*H�DJ(���C�-�!�Γ=w���DF�<J�	�RA�1k`!�DZ�fPD�Ae�ď���iT��;BP!�$�Al��D[)s?��@��"i!�h�ؤ�_� USɌ8nC�I�fԱa-^�`�Z�PlC�ɽlJ�l@D;I� � �i\C�	��b��ڳDj���b��-�^C�ɐ=�a1�O1-��`#���+�xC�ɉ
6���L�X�<P��d�fC�	�nS�����/O]�x�%G94�hC�I��|�KƊַi���6	�(�bC�	,�4�Xd�&��8s�e�?	�C�I�jt� ��'�+��L�r��YV:�ӶɁ^q���d34�P�e(�>��<rcj�V�!�D�7��)T��k�~Qp���)~!���L�� �قt�P�+D
`�!�D�~t<�8�RթT�V�?��M�ȓn_�ؘ�kݮx�I��-H-��ȓaQ�!�#���8Kܘ`��2td �B�Ό��O��	j����m]-������P+*����P�x�g�!VUd�á�|ʟ4�����y�Iɿ�-�5��?���LK�A�'��<3�'n�O��#T���Z����:�&TU$�5J�+�yB�XPdV�����?�����e�~�iFfT+Q8IxA�ܼ����2�\��i���?�9� Ƙfb|�zP����e�`*:�y2�(,U�!K�����	çH:t��\R:԰����;�l���HTA�kZX���}�"|J.��T"q��19Ĵ"�T9�B���`����a� #L����;+a�		3Q��T����"2j�% �7'��4�J	Oi�(�0��\�y{���t�S��,��s Yl��q��W.�q�`��9�˓_�`�çYw���t致d/���6��U5 ��egH^~�M#'�hD2K~�O|n��b[<�2�c�)z`.�����97���]�ꅱ4���ҧ(�<Y2j��pH��K!-��� �W�<�\Һ�Bh�m�)�'w�,��씖^�٩�O�c�­��S�? (1@��ו]VE�@��,Ry�\�W"O�� �%m����"�O�\��	R"O�5@6I��>����F� YC��p$"ODE)t�  �@E��$�1:ٖp�e"O ��Q/�a��U�'J����� "O���V�P�1��6�<��"O�����z�
m[�r�:&"O��8�"�R�1:�d��W���J7"O@�0��=D�v�4JZ<��$�#"O�,�w.R`{��i7�WY�.�f"O�%��\���eQ#׶A��"O&p�4��	2�N� ä��G�蕓"O��1�u�.��A�V"O9��Ȓ�X���<BQ"O|��l �P&��I�`�:~����a"O��7��X�z����Q�4M�"O�`� �:/ZQ ��W� w�T�V"OL��j��}#��2g�0�"OX��O	�%s���0 �1R2=�d"O:��q��@:mI� .@�v���"O4���D��fc��p��RO���[�"O�q����1)�Ji��XN���"O�1����|1��(��6G�pR�"O�pA�g��2��
G�?���"O��c��Ҝ>�xZ�h�K�H��"O\�V��Bh*�"���G�!�"O�y�&@Ȫr�C���"OJ���E�8�0ت�H&u>>H(�"O>��Ƃ�L^�R���\���j�"Or��$Y?j0�N[� Fd��"O�M��HY�Wr�	b���Y���P"O�LHTȍ7$U, a��ޯsB֠Z�"O��YDm���� #�0T*�t�"OH�����B�`�𠆏�<��"O2\iF��8��u��OM9,�D��"O�9��)�R���k�-��D�L9("O����|���+�!p�X�"O�hpO���R!�'h�jp"O��0&Mߵp�n]��ET�K4>Х"O�Q�J˧^v�p��E��!F`�t"O0����ܼp�
�4fêdکk�"O~�a�5�J�Pa��_n�1hc"O,�s�ۤVT����X�c�r���"OB�Ck�'JR����!T� h5�"OdX	1�Ͷ/�f�9����~�YR!*O�U�3AF���� O�=$j(-I�'�ZP9�a�+T��k��,$Q�t�	�'8��Av�{���rT�ܖq���P
�'5��rӎxe���Ȋ4H`���'��@�gR?x�b�dD��ذ�'�d�	�P�ԭ)��~.>�)�'�$��O��� Qc�S~@P|��'x��0L�ӾA�s��}���'z�]�a����0�lS�n�@��
�'q�h3 ���H��U� aA�N��5�	�'4T�����m�z��@H�B�bA!	�'��IRH�"��ѧ�.��(�'��8놬V1~^ �'�)���	�'�Rذ�툕e��-z�eR&*Qa�'c�x����g�`�����`�X���'��q��N-3�L<YsA-\i�q�'�A���]"q;\iq��DY�N�)�'��y�*/Vi�);�	��D'̙H	�'~n���N�; i
Ĭ=�$���� 4M��snX1:���:]OhXR�"O�� GI]=&�Z�%N;�d "O���"��PA@�(�%��6��YK�'(G��	
x)�r��t0���'���*�Ô�2b� "#�4hHI	�'90ઓm��I���C#�ۉv�9X�'���aBB�b��<��K-:ɮZ�'��QhD�Vh����R�Z�"R<Q�'��� �+�9�ʸ�"腘&�DL
�'��pA�̦6 �\3�$ޅ Ґ�I	�'�0d�a#08y>�CqO�:kZ
�'�Zar-�"d@���fD;-P���'���#����ٷ���\c	�'>8xVj@9GIP=i6e���p��'�4�2ȶw���P��Ը*�'$���C��E�!�g��+x��Y��'����B& �h��ǅ"��'�&�F�4#쌱@�B�H��S	�'>�|`dL3h0}{V�@ D�����'I��c�h�2B���0��"Bڌ�Q�'�� h�&)\N�Pc�ؕ+*D��'4Lq �`Ɔ"&6�X�B6r�Ƽ��'���*sN�2U��v�\7�Yj�'�=;�gjO��*�L�!�4 �'ۂ�4�ғg������P^<;�'2d}ÕZ$G�2�k�S�-�@��'��1��\�:Eh� ��$5�8��'u�m���
S����!܃km$Hr	�'�(E���B�(����![�`��	�'��QeaJO�d4���6	�(H
�'���3`��V<���P
�' ����!��,��R�څ?z���	�'Jh��ҍP�xԀ��
�LZ�%p�'ޱ�Р�
Q��'�Z�mBP�[	�'�zͻdg'$iX��P�8���2�'7��P��3B�=�398=�p�'�X���/U�^Q�3!%7*��	�'�m�CKиy�6�H��^!|<x�'�p�k�⑧_��m���6ph��A
�'�v@���>��㦅Vb�2��	�'��T���5$؂�qsm�Vt�q��'�B ��]b/ˍxx2Y��'c�d�Ĥ��|��g���Fg��h�'�H)�ÎH���� ��+A����'T�f�ǯlN�Hx��:F��B�'�҄�`&X�w!�  %JL68Y�5�
�'�v�0��¤���I6.F��@	�'���2w/C"I�֑Irm��,x��z�'R����;f�>���d�1*�:=��'���C�/�L�+����R�8K�'s����]z	J(�W"O
!�4K�'^��G�t������4���"
�'�qs��@Y�6	B�Jո-�9a�'8����H&$��ɉ刚(t��8�'l`����R(-� �7
���
�'1�u��D͊Iwx�֛֡X;�\�
�'᠄�G�9�إ8VCӛ (fh��'�H����]��$�E�ٰu��<��'�4����7\B��%*Q�m%�b�'s��P��A�H�U`_�i�v�R�'7Zᒰ��E�z( �T�IV��0�'��	0���mi4���'�N�,���'yrm�!h�,~�RT�	L�j��'+��!@�Txt��Г)M=rR�i��� *i��� �y^�x��F�>CP�G"O`j��_zNT�kEf� &��"O�ps ����������7P�ސ�d"On]#�)�
H#5C1�G8f�j"O�)	䓙�\p���S�,S"O湰�h�<����VH�i"O��a�&�V��p�'Yug�A��"O���`�a�>ٙ���Mojؒp"ObtQ!��Q��,*�D$b}��q�"OZ����ДJ��*$�C�8e�$�w"OVA3��ϹP�*٣!��.c�	3b"ONXۦd٦x$�V!=q���"O4zQ�Țu&H�2�N+,��I�1"O��Β�_�>u��.��E� ]+R"O��i��2@���h6k=4d�	z"O�L�%/XE�X5{��mM��`�"O�U�3W�=Ԍ�#u-(���"O��J�ޓ�f��a���C)n��C"O�}Q2�UpN�ᛢa��T�,T1B"O@�j�*�f$�� �ʥy	-�3"O���	Z ^� e��'q�$�"OZ"��M��%��B�?��I*"O0��Ў�0�D� �C��[���
�"OY��{K�H�`mۨ�<�K0"O|mcĲ$!��(�	�$Gl�H�"O�س%�N�tTH�0H�!�Vq@"O���LT�w�$yR��j�5HQ"OΩ�ˎ�^@@r�(��Z���x�"Obx��/EH.xQ���H�N8�"O��U�@�آ3ĆB�[s���S"O ���3��A�Ř��Hz�"O��#��0X�ډ(�B��~�s�"ORp�$*�-�Bq�T!� E����"O��C�B7"Ϥ(�6�Ϯ(A�"O.)�2�H�^������Ґ�\`�"O p���2/J�a��흦a�>M�"O�<�s�3}�i�SNǈr���9�"O��`�l�
<�Q�!R�>���&"O���f-�*�4a�\,ej����"O��Ȓ�[$g������ţOɌ��"O^��r��]}r퀆 F�����"O��
f�J��"�P#oj��=1�"O���!%��t)�<�4�Q94{���p"O�����ܑX���ktIL�Kp"Ob�Q �[<d�����]=C2�`�%"O L��еp� ����7�X��w"O荘�%�W�\<����0B�:R"O¤pS��5n3�#c�|)�"O�@6FԻ`wZU(gce.� ��"OV�H�N�X��Y�BΐƮ�!'"O�|�S �&
�}Qs��Rd"O�$�6�)��#�o�S�� U"O$3&f���%������K"OĔ��L�J����c��@����"O4��	Fm8$�Vƒ�j�c"O���T�Ifi��D�,1��L��"OH�
`�-J:Y�ᜐv�����"O��"qg�z������xľ͹�"O$*%�	u$X��σ�|����g"O������Vo��`�#K91�t��"O��J��S���a�� (��Q��"O|] W��6Y�<!pТ>tz�Q��"O*4:��3r���"��ד?X�(��"O&\#�C�-�"q"��eI����"O� ���6�eҐm��]+P�8@"O@��%�ՀK�����I����g"O��`��#���RvƘ u0p;b"O���7�� �-j $�A�e�"O����N9Cx�B���3f��k�"O�iw��")0���g�3>$i�1"OL���G	p`K����R��Y�"O`�H�d�)�5fE$Z6�R0"O�i��̈́�c.F�3#ͻ)6̰�"O� 1�no��u�D�¶M�ty"O��s�	   ��   �  �  �  �  d*  V5  �@  �K  �V  �b  �m  �y  ��  ?�  ��  ɝ  +�  Q�  ��  �  e�  ��  ��  G�  ��  4�  ��  ��  %�  ��   c	 �    �# �* U4 �= �C CL �U  ] Cc �i �n  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^�+���������Q��_�P��I;Tf�����a��3�i�L�C�I:V�Ł�
Ӥ<��
�f9��C䉼R��Ӷ���a�f%y�ϓx�:C䉢G�"P�͍f`��{QK�E�bC�	� ڦIAVe��y�$ �`N?hŀB�	`j4��f��W���d��"C��?0��C��|̩#�]�z,����>9�k['	U�H���#�~X�V��C�<��
R�2��*6a�#" �]�q�z�<���%T���2��>�&պ�Uu�<��Z�},L�TTT���Ze��e�<���[7 �:ӧ^��D�Ej�{�<��	�4&�Faz��. L:W��px���'U6��j�4{HIi�J�=<���!�'@�<5"ށe�L@�B&?K�y��'�AC� ]�h R�d�2v|3�'�R���l�2#�{��L"5��`[�}��i�ay2��L����kh��պ����y�C�@Y��c�o2bX<�ْ�Z��į<�K>���U?��X&o��@rJ#@�g%�1P�'W��4�� �$��򌓈2��Bu�=}��'�6䲓k��_�,���펫��t�	ۓ���w�\a��G�r(]�~x�
�b D��*�m͟&���d�-p���cѤ>}��Op��S�O�.�@�,��(D�(�Ɗ4p{�Z�'q�&�ĕ۪��fh��e�����C?)Ց��F��'��-C5��9ND��h@�	�0���3�'K����KW�("4#���Qb�	��|�h*|O��C�3e,N}�ڕ���>щ��~��'�`�PuE�nb.� � 1B �
�'�~�re�0̖y�P�	0��)A�}R�)�Y�s�2�s���O�Q��a	�|n!��<J��AS�ϴ6�2��aP��1O|��dA�9�#�'�65�nd�q��v�ayr�	��&5��=nv!��&\[���y��'�A�E"4x����UA�|d�(��'��EIO�Bc��$GU,{ ��'k�8�*�I֚���j��{���y��'�,Q�߰n/������Rщ�'�*q����� �C��h�eO��� �=Bo�]��nJ�$	.���'˛7O�+�h�d���Q���ݾ+0���ȓ,N-��B�����FhdZD�>�U��$x�����[f��Q�+R��pǦj�<)�ʂ�a�(q���¥c�D�bH˟�͓�ا����`Ԋx�L	{�,���\�bL%D�����+ApbC�;`�����<	�S�? ����-ϷQ�<=Q cۚtu���O�u��D��^kr�[p�W� v~�q�K G�<���@�B��H�fD�?T@x��� Y����>��T8B8�b��4��(�t"�Q�<��/��L1��*��7X�*����<���S���l��J���髴AT�Q�B�IS���4E�82"�[��E7^���0�S�O�ʜ3&��^]A�T�W��@3"On��I��L���򭞠,�jPc�"OԐ��b�>ZҁC`�N�>�X���"O�A��P�޲�$f��Ѩ�y"O T`�*O6/LLI˰E�M���w"O���Pk�*ˈ�Jq��X�)Є"O��8�,�/f�P�Z�.
�:H��1"O(�D"��2},)T`΀,���"O|-A$YO��9�v��R���9�"O� X2eb�����,�I�4"O0|sȐ�H�tZ��L5x�"OFÔ���($J��1J�Vb4��1"O6��DfC�Z��Ƙ_G:�Yu"O���eP3*T��p2EX
n0*Đ�"O~�%�#�Y���G`��"O~�@�h��x�sc�0b(��"O0���l�) "�u�۴-X��"O�x+�O!�̨���TT����"O�%3�	�1�V�q�-ӼVb��"O2��"���!T�F:wG�,�"O.pB��/E��c�m�@0��"O���d�7�^ #',	�w*�L8@"Or|{Ӊ؍6Q���<}"��#"Oz�X�:^KQ2fkD���˟��yr�F�c���F��q���@�R.�y��')��(2��'l;JX����:�y���S.8h�ČM��x`����(��,HG�׆%���X�`� a�Q�ȓ{��2�h��a�!�Q5E�Ta��TJ&���.W�8��!�9����I�D�˳+�|�4����Bо�ȓa��(:�C��(�+ǳ!�܄���|6�ڰ]����`�
"���ȓW�� ���*P�	��*&����J՛���U�Rt�K��f��\�ȓUn�p@���Q�4�C�	��*�� ��K��ѡ��ml���7��gN%�ȓZ�*���!���YF��La�s��i�(P�t��+M)�l�ȓ[V�Tav
N.l�idZ
!� ̅ȓz��%�ttQ���WB����ȓn�
��Ո)cW�;s,]�/�̇ȓT&��cK99JyK���1Y��ʓsՈ���m��y`�U8�j�8&RB�	��f�y�@K�{��c���*J�bB�	�i&0p��Х�=^���(��yB"M�v݀�� �\=�,���"�y"�T&�9"&E�Us~Ȋ3�^��yB��>/�-y%n�?G@�@{"լ�yR�K0�r ���@%��bf�"�y��J +�n Pg�5/���J$e� �y��'::��! �ܜ"����s+��y�◜f�x@óⒾM.����I��yIC�d���I�X6�; %�:�yR�)6|�!v�Ӷ%�L|�흉�y��Q�WH�q���K����y"e�:�ؔ#�o��`J�b/���y
� ��K�cд� ���&W�4��"O�P��_>(ލbV!�0sy����"OP��ƃD5	�# ��wb��q"O�����:�Yj�.ăzO ���"O@)���>bɖLz/ԫYN�sE�'��'���'���'��'�"<xŀQ�6:.�1�dJ4S���1s�'jr�'���'���',��'Z��'d~D�ǄI�H6:����T�C�h����'s��'�r�'[b�' ��'��'��|����Y���ڥ����~����'a"�'�b�'���'���'r�'¾}B@��m�thg�r�Jf�'�b�'F��'j��'R�'���'��E��/��z%9E&D�THX�'���'�2�'�2�'�'L��'�T a��S[;��S�%R-5d�����'er�'a�'�R�':��'nr�'k��)�f	�s�Q�F�|p�����'B�'��'���')b�'V��'/�q�ݳ9�Y���z�2`��'9��'���'1��'5��'�R�'�DA�逯 � ��a��>ċ���?����?���?��?����?����?)'gٕ,�5�`�*EF5�S��?����?���?����?��?���?���.zvZp�g�SIh���)�?Y��?���?Y��?m|�`���O���܍}�Ăbi��	]�pĭ����D�O����O����O~���O�lZß��	�1J�u����nʡ �	�>>��+O��$�<�|�'5�6m]$Y6D�/J-:�����zfV͙�����ߴ�����'�Z�И�*��l�X��F��g?�<��'��E�0gA�v���Χu�4�~B��%[��HA0�<l�@�"�d�S̓�?)-On�}ʒIJ� ���&�"e�,0Y�D�����_���'X��oz��1��	/T�Y 0�OlU�m	'�U͟����<ѮO1���P�/oӊ��x�f��R��)����F�?`J��I�<�"�'`��G{�OF2�NA,Ё�@�Z6*�Q$@:�y�R��$��!�4z7p��<)�dRH���˖�E_ˎXI��1��'���?����y"V����a��%��Vh�'A/���`�5?����a���Q�'������?9�I� ^����*T�+��A�Ԫ���Ħ<��S��y��S�9`�7>�x����"�y�DxӒD�՗��x�4�����L���}�D(AA�ҩR�K��y"�'���'F�T�оi����|�u�OW|@�ϐ�s��7�R�,:$!�Jd�	hy�O�"�'���'����=�ځ(a)*Q��+e�!Y�	��M�����?���?�L~Γb2���O6�����.ݏo��X�R��zߴ)�&-#��)Q-e��KRNK���;��Ԋ �f9�&-�=8��ٿ9F�hƨnҾ�]��?�@��4
,OR�a!�J.��CB�i������OJ���O�� ~1�5�N�<ن�i�BDy��O��P%/�u`D�A�0-��Q��'�6��O�ʓ�?�W� 0ܴR��V�'��U��O�Sx~ib�g˒$fĜ�Q�˛�4O�h���'6b�;Ba�4���D�H��ݿ냋����ܻ�@�>o�!i��<!	���4������4hhR Ñ84�����?���N,�����˦q&��G@X��i���F�K�И���ē6��FGz��iņ3� 7�;?!1Κ�o�R�0�@F-w���H��ۃdd ������&��'��O���F]��i�D�7������I+�M#��@�?q��?�/���9�g�!-@�xp�Џ¦�B����O�m�?�M�f�xʟf��Q-�#l��p��
�eC��w��ʁ�sӎ]����PO?�H>Y׎ʹG@�@���&K�v1�2(�u<��iz}��<pn$<�A���J�m���S*X��'(7#�I���������.s��IG	�3R,�k�"E��M�u�i����a�i�������AQן~�=�pX��,ه� |�r�Ҋ6�����$*|Oi)��Я8{�����#z���̛ݦ��tN����џ$���y'�	�qY�\��iȊ�
FŽo"�6-[ݦ�H<�|�)�M��'�i���B�d�Lc�.�*�l�a�'O*l:���u?�O>�+O�˓_����Ӂfʁ#�����U�ቊ�Mc�cN8�?Y��?y(M2`�r�ȶ.O~Y�Ђ�&��'j�/���bӼ8%�t���#`[�G��a�a�Cd,?������ߴE�O7����?��.�Oy���ؠv����b�<�Y�Jm�ĹŅ�#5�f������?�i��Hy��'��|ӆ��݇J���!� #W\DbL<�I!�Mt�i��7mU��7<?��n y&��<�Y�C	@�&�ȥ��(v��4&�Ԕ'�b�'R�'���'̺���q��4S�A2j_��0BS�0+۴z)ZU����?9����<�w!�k\���+-�d3R��z��ğ�o���S�^;�,�n��Hp���	�xIa���0��� .��J��O���I>a*O��hT��P4nг���?�X����'��7�� �����T��l�t圉7H DAN��<�d�Ц��?)�U�@��4yx��!{ӆ!��ۺI��h��c�����(��~�6`����?iK�ӟ^ʓ��{�? �l�W�F��ҥYQ"��@�X��=Oj���O���O��$�O��?�$c*%!���X���X��L���@zشkϧ�?y��i��'���t�F5��.ޒ8a�|��*�$�����|�'K�
�Mۘ'��L� ��
L��br�O)K]���6,d"e����,&��6�+�D_zy��' ��'�Ү�(I���Y���#5.��$٣C�b�'�	�M����<��?�(��I���o�噁�G�/�$���� �Od�D�OV�O��G�\Zef =|V��N���<y$�79��xm�P~�O��l����!� M��F)/�A���(��I���?����?��Ş��B��Qsph��L�b,�����DyS��f������A}��'�jH�rcK�`�^�s '� K�8!��'<��3؛旟�ز$�1W�q�A���fR}ʓ�e_��01O�ʓ�?����?!���?q����	�3qv��h���A�E��2�mڶg��	�	џ��	S�s�Б���3'�U�=ռ�I�$Ց�F��$&J9��z�Z-%�b>	�sm�Ϧ5̓/�*Uj�̞d�4�A������ϓd̔H�&��O0��I>�.O�i�OB��:G��"%��	�=0��O�D�O���<��i����'��'��dx�R�N�4-A$t�m0�|��'���?����tӴ!$�`�e��[ⴭ��O���p���|�d�	�Y(�0�-�Ҧ5�(O��	Z0�~��'�(p�S"[�j��u�,N�q�9ȧ�'lr�'���'��>��ɇ(��a�U�H�`�"z�Y�I��MC�AP��?�FW��|���yWO� -�a��H���q�P�T�y�@|�­o5�M�Lج�MK�'�r��NU��k�t�@�$g,��ӤC�D}�L>�+O>�$�O��d�O@���O$�A�1"gV� H� ��A�ĥ<鳰i*B�"��')��'#�O*2���R|Vn!1c��S� �<=��b�6�h� $�b>!X!腨c�\�T�/ڰ��EcC&@J\nڪ��-sr�'V�'��	/
��
�F�<[��&����؟�������i>1�'�6-·w�$K 9F�����m�Ȫb�X����e�?Q�Z�����H�	2	f"����x��H�b9���'��U�'��u��|r�;h,|k�)�F�L�Q��E�?�<���?i���?����?i����Ox��:4A�j��by��)y�'b�'{6�6��I��M�K>) �ҧ���9�GЁJ��ecҥ�2�䓚?a��|*�� �M{�Oț�I�$- !��z�8#����\�nHr�'��'1�i>�	ݟ��ɐgc�͉SE��Z��5[bϯo�8M��	�7G�*��'��7��"�f���O��D���ND�)X��R ��m��<���O*���O��'�"�'vɧ���'$x�"�ԈT�B3���?5E 0��42�:���i��	�?����O��O=z �M]�F���-n�����J�����O����O��<�6�i��`"fM�t�x����v #ŕ&`�	�Mˏb�>���iT$�y����c�ˏ�l���u��z�֭k��dyb|Ӕ�l]��^*�T�~�80�����!4���<�(O����O����O���O<˧L٫%e��;��=c��B?+ݖ@IҲi��qU�'���'��y��x��n�V��0ɓ�2��52���'~@F\��Ӧ�IN>���?=�
t�Ul�<����M����ጨr���'��<�D��R��ߡ����4�(���>S��q�<f�ڽ�$�.���D�O����O^�fO�&&*C���'�R�	)2FFd�����C�](�*��f�OB%�'�D6K��QpO<i&�μvB�W`K�P6�2���y~���6���c�G����O�������R�Q�T=�A�Ӈ�'�����$�j��'b��'V�ݟ��Bǡ20�P���8��}�� ܟXK�4s��y:���?�S�i��O�Ύ�qÜ�� ld�Q���!��������4n՛���#?J����d�6
W	F�I�ni�PA��+��		1�l�K�m*�$�<����?����?��?�Q��7�.)X�K�H��][!���ܦ�)���˟���ٟ�%?�"!\u��i	�#� R6�M��!�O�m��M㳙x�����#y�f@
�G r����'$L U�X,j��i�2˓#a����ⱟ@'���'~*�`�J�#��Q�'ױƅ��$O��'���'H�OI剆�MbG�?�w�+H
1�i�&��@KU%�<���i��O8E�'��7-զ�3�4,�����LTR�0�	��'�4i���F�M+�O�L2��H�������wHԺ�M&�,@FlE�4��'R�'���'3"�'��2! �*�2m���ˉzd� 7;O����O>Hm�$q�d�uۛ��|"b��;��ڴE���yãńi)�'�����R�Rd�����G�6 (�R&��q�]��x2�Q�OޒO���|���?���j�b�	�gj�QSdCZ6A: j���?�+O�YlZ�����?Q,�>ha1*�+}"���e�Zv$�v��|��Od���O��O�S":��#+ӥ����aY0f�\)��n'Z��lH~�O�j�����Z��}�e��N��3"��^�B���?9��?��$B��O_剸�u�*�<�Z�Eʒ)�8�!V��#P�DXݴ��'f� *�6��4��K񪀶/�n�R�K�"�6�
Ӧ����	͓�?���E
[���}y
� �	9po��\"���f�Con�H?O|��?���?���?	���iϚ:l��[!�ȇFF��3���
~ZmZ%j�f�I����_��83��w��e:���u�6�H�H��`�]+Sy�|nZ*��ŞdKD�ߴ�yr�ƴw�`�2���z�r�p�M��y�+>�i�������OL�R�xh�1
�	Rv�0��,Z4�$�O����O0˓O`��h��;F��'�Rf���4왂l� �.�p`�C�n�O�'{��'��'F*m*pa�* B� �QF��gV�a1�O� �qʛv�*����i���?����O���c��z(wHK"9��i����Ov���O����O�}b�W��b ��o��8hHM4�T�+��vIًn�	��Mӊ�w	t3�Άr��,ɷ�h�d�h�'x�'�¨�M�搟��A�����e��y�$��7d��{0�S�脀�pc>�$�<ͧ�?y���?	��?�a�/A��-��n6R� 9#1#�0��$\�Q1c�y�h����&?�IF�>u�"�q��T����q#����O����Or�O1�X�7}.��CÓÄ�ˀ��y0�6�2?	���zK���e��|yB.��\Sf̐-#��I��E����I�����ޟ�SIy�oz��B�1O,����I�{~�1�X�q��y�?O��m�m�#m����x�Iǟ���FE*h�"}1��I�2�i���ۄ �4�oZ^~�Bn,�E�t�w�H�T(���Ā�@�H�b�i�'���'/2�'�bZ�b>�@B@نI�V���ĭ��X�Qx�t�	韜��4��'�L7-<���+L=L�S"^-½�f��S�Z�O����O���Y�>7�8?)��_�TD� 3���Vp�!�n�� .cT����$�(���t�'%��'���fGP0?A@	���O��5���'ebV��
�4hO0Hϓ�?)�����fB���/�$�D��"�[A�ɱ����O.�D5��?IR �Nq�.x�1�L�MH�! �	A$����AƇŦ9��d͇X?M>a2/ 9I�y]��)�+%L� L����?����?��Ş��D���]��jT�\b�t �`ڕ"TTŃv��.Y�D���ǟH��4��'\�ꓝ?�[�6a
��a�ɬ`Pj����?)��,(6�B�4���L�,j\z���@ԍ8�1w@B4�1��ܦ�y�S�h�	ퟬ��˟�����O0���e&V�I�@��K!k���+c���A� 	�Op���Or����٦�݁X�葱6�Ӌ*粘��fF�V��	ɟ�$�b>M����禑Γ	���Z��$_p�+
�=���E�4@�Ǿ��%�Ė��t�'ǈ���#O	+��1`�E�
=p�I�G�'xr�'rR���ڴ��4����?���{��!��	W+B~^�ۆ
�0�p��b�>���?�N>!���))%~��d@�7<q´1��P~�� op6y#Ӿi�1��h��'2�(N ��u��k����I7�y���))�� �a߽]��r!�>a�b.n��d�+�O&��Zɦ��?ͻ�ƄS��9�Tru!��P:1�5��vg�ZYlZ�-s�(nZB~���"K�d��Sl�$S
׻]�����W�d�TpO>�,Oޣ?A��7��@a��#���鴧A~�Gy�N�z�'�O����OR�?�@d��W�\�r�'×x�6��_������ߴx����O������J�7� s�2�|a �Ao-�v(�<a���o��	t�Ivy �"�ya��I���8����YS��'9��'�O����M�����<�v��`�����H٘u�w�M�<1��i{�O��'Q"�'��M�,i�� �*!:'̘�����]JҽiL�	D2�ۂ���H��9R�$<�C!�%lf�8�c����I�G(��V�	A�,w ��q�T����	7�M3�\�d@sӺ�O~,;��
�=R�`́{x�ѳF��r��:�M�R���t�U�v���XVGՋ��\�P �"�����_0��� ��O
�Ol��?Y��?���(A"Gŗ;�Ebt ���M����?�(O��nZ7�"��Ɵ��N�4oj���H0��!B��!б�D����_}��'S��|ʟ��5�^#km��b���-Bh�:�どj�~��1�o���|�租�'�|Z�蝉z��m��Á\_�Ի��&�$;�4. l�PWk]?B��)`ď]NP<�! ��?1��E����}�g`�"�&#iR�Cɨ��<�o��{ю7M�즅��&IҦ��'�d�P1b�i�-O��9��J�4萩ӓ@�߄�P%?O�ʓ�?����?Q���?9����iױs2Hz���^Ҫŋ�O�3ڭoZ�Xx�������Io�s��!���[��Ԕm'�9� (*��x�"�ɾEB�i�O�OQ���G�i��?����S�M������ ��D�)d a��dК�O��|2��C�ph��շ4�x�H ��64<eC��?1��?*O\�m��4b�IП�	�/z��󂁂(甡q���I���?ѷQ�����%�4���R�R �[AmY�{ !#��'?��B�2ZV����4�O��D��?�W�C҆U��L���L�"�t�<���Y�܅ʡo۾(�$�QMY��?�3�iY�5�W�'>�n����]�yX�= �/��7Z1XB`F�X@�����m��M�"JV��M��O(�6�� ��� 
x rk��;ʅ�&G� �Љw�)��<i��Dɏ[`$��
�tK�,��K7)���)�M#����?A���?���ԇ]4���m��$�"��!�9s��?2�fr�b&�b>5�d��%>,^�E-�8&�X�Cp
ĮJ�=lڱ��D�: BQ��'��'��=+���ՈŽ_Xnd8�$�t���	ߟ�������i>ɔ'P6m�|��D�S��"�f�( L��2֮�I�����I�?�s[�\�I˟���:C	�Tb��;{�x�:����{� a�#B���'�T�B�O���\�5]�}���Q'9���RO���y��'
��'���'	����-.�h�[d ':�@R�](+��d�O��撚�1?i@�i�'�f��0	Q�t0��R� X�B��ӝ|��'�O���cU�i��I�.�2a�P���@C�kC�Z��K�jN� �$:���<ͧ�?9���?�@C?[��x�É=��x�ɕ��?�����$���Wyb�'�ӆP߬y����&B<�g�as��J��	�l��u�)��$��z}�k�iD�j5�ͱ��L9	K��OH�n�R���Di�џ�HG�|b�A�n�J���j�^�kS�Ӄg��'���'��O,�i�w���	��MS����H܈�@̯P>�-c4��1�b���?ᑳi�"V��*��D�O|}��E�$P�������HQ��;2��O��$�%�6-w�x��*Iƺi끟~�����L�?�,��v�Џ.�J,�����O����O��$�O��d�|"�O��W%�ap�@Ҕdհ���H9כv� �l��'����'��6=�Jqц��au�)�2 2z����צ9�ٴ`���O2��jӽi9�Ĕ�9����t�H U�
����T�'��$�׼ ��J�O���|���9:F��B��4V����%�</B(�����?9���?�+O&`mڮqO���ݟD�	�A�X� ����j��$�1��p�~��?��_�L
�4gԛ�'񤕡V�|d�tM�[D k�HX7���pe���P�X�)O~�!����	2J�"��rH�:[TlL��,�% �X�	ԟ���ϟ �	y�O��B�&OVL�!�dP*El��T�'B@qӺ��W%�On��ܦ�?ͻ���[�)Q�>_^!ɕ&מG��Γ����k�t�m��B���m�G~�͚=��������V�[g��%L�e�K>�-O���O��D�O��$�OL�X��[8B�M�;bR��95K�<�׶i������'u2�'���y��E	p:�	��>_����_?J�n�w���y���'�b>�Xp�V�b����c�#-|��ruj�=$a�+��7?Y�jðwI���/����C&����C�.v�@��Dd[�a��$�O����O��4���1����_��ybÁ`ː��n��N��y22�V	�y�j���C�O��d�Oz��fB�)D���n�s P�1��o��A}�(�G9�'���2��3�������4䪵ӵk��<1��?���?A��?i����7�,R#'.+�� ��µ��d�O�mi���>y�6�|2ߟ9�̙�����<����R(�'����$Ԡ{��������aN�P�l�2rNN��[�)�"�D� u�O��Ot��|����?y���h�0��m�@X)Dˆ�&�6����?Y.O6(o�+}6���0��R����3���v�.��� ��$]}��'iR�|ʟ"ՙ��;Ѹ}9�ʊ����FR�z����wӌ��|z�⯟\%���F��X`�K�aȚ5�*7��ڟ��	�4�	�b>��'s�6mV
FIv p D(<���A9w;��S���8�޴��' ���?!��;1~J���%Y�G���B5Ɯ�?I�{��i0�4��D��a=h}y��TIO3N-B�h�g9J�+�N&�y�R� �	̟��	ٟl��ӟ`�OS��c�oٔ8㎈��ڥ@k^�sR �$�7O�D�O�����ͦ�"���׊�>k��+uj��2�rh�Iӟ�'�b>m��I�E�)����K+���2��ӱ�vΓ>t�S����$�ԕ���'��Ru��W;�|"6eUѾ��'T2�'p�\� ڴy�����?���c����FF�]�8��m�u�Q�R�>��iӸ6�w�%⤙A&�K��Ш*�B�'*�@�\��e*�T"!�|u*�O
!9��{�<��D?NHʰ	��-<�E+��?q���?Q���h�����<$J��C"Q:b�d0�c�����¦u �b�Zy"E}����];q��ڄ(f��ǎ$i� �I�L�	����G"_⦱�'��	��iZl�E�&B5��3��F�)������4�T���OH���O8���*R�Cs��m!0K�FX1x���������y��'hR���'�и�Â	S+�T3B<v=,�1V͢>Y���?�I>�|"Qi/]�D3�e�'5�tyVWO)Bu�ܴ���Yo}r�8�'��'�����3Z?b��XA@#7~�����'2��'�r���V��bٴSvU��>����_uL(�"I[�|���r�F��Z}��'YB�'�T�!��^Tݬ���$��	�A���oP~�ț��V���]ܧ��+��ڟ��Q5��59�^0�CCC�<q��?y���?���?����̍;E\�Gݩ\�T1�udAm�2�'|��p��PY���<�#�i��'��kagʷQ��9�o
M)����|��'��O?`�q�iH�	�Z� dE��6*�sJQ���)4%$�?��"!���<ͧ�?���?y��Iv�|��F��!q�p4�,�?������ϦY2���0����$�O���xCW\Jܡ��<$�0��O���'���'9ɧ�I��4����ӿl�֜��Ϟ%�) �*߶+R��F���<m=���Z�5{��H&���S$�Ace�ƃ&�.9�	ݟ8���T�)�Sry�d��UM	�'e���3n	�\
�]�S�8yԒ�D�O��n�x��#��Iߟ�@ӣ�$~�ܒ��5>�!���ӟl�ɲ,���o�D~�I��(����M�I���h�b��E�3������7��<a���?����?����?�+���3t��n	>�x� Ęu����C�����ǟ��Iߟ��C��y�4`72��#*�� ��Xc�`P r�'�ɧ�O���0�iH��JJ��ÇEצ�K�k�h��ԏ
0.xx��A��O"��|���҄���0(��Q��v�=���?���?9.O�1m�8od���?)�D��"\�|#�$�<";`e����'�<듒?!����
�ܩ���}��`�h�B��,�'��E����)�6��]+�~B�'����Qg�>Pר�@�H�8=�"	Q��'(��'�r�'��>���T%�Y!'&C�:D�C Hp��	��M��-��U�I�?ͻJ\�ą8ac&d�3�A�`d"�	����ܟ�B��
���'s��h�L�?����ԏ�9[D�� �<�:�KH>!-O�I�O4�$�OD���O�嘕��%e�X�c�-P;C���<�'�i�fQ��P� �Ik����p̃x%�"&Eǖ/��@��.���O��d'���_d�%��芅0+(��c(�)V��}{�.M�~d�	S�����'��X%��'Fd�U/I�YL @��Ŗ89<�v�'���'=����4]��شo(]+�J��05f���P$4S;hΓQ{�6���X}2�'�b�'O��#�K^�X8�%�?[2B��4K\	s֛����Am7�Q>1���gN�#��ڠP2(���B)�	����I�T�I��	t�'F�Ɣ�d�9"�� 	�(sf.�y��?���(���� 3����'t6�*�J@O��G��*Q�E��G�Z<��O8��O�	��7??��Փ%^�S4Ô0d��U�����5k��b���$'������'<��'L�q�n
�@�#&�\:\0S�'�b]�(�ٴ@䪼̓�?Y���I�"E*$�G���$��`��XY�I6��d�O��#��?��@�Xt�ar"D0B��{�����O��%��tėw?N>9��V+H��Y�$��n2�B�@�?i��?A���?�|�(O�mکh6|�'�M�
ܲ�;'���A��{DDgy��Ӡ��;�O���l��N �D؍(�fp/�����ORԹ�oӔ�*[�91�䟶�Ol�}���-��d�L<z|D�:�'�����0��ϟ,��ҟ\��K��(>��zB��/M�J��V)��	׈6͆8mN,���O2�D0�9O6�oz�yR���U�n�G,�>�bd��o��?A�4b�ɧ�'E�`Xٴ�y��+<n�9@�:�۱��/�y��F�#&1���
�'�i>�	,%�VQ�RHA����b� T�h��	��<���P�'��6�[(IA�$�O���
�,8p��X	e����� S���L٬O�0l��MK�x�.�"m9A��^�"����K�����=D��4k��ϗPy1��0+��Zy��D�0Rbp$S�Gѿ}�!˥+R hL�$�O<�$�O
�d �'�?Y�j0�dPR�IݣQΐj�)���?�S�iB��r�P����4���y�b��)���kH73�Fh�c��y��'��'����ĵi��	���d)��O���b��؈A�U:�L�NC�p�G�n�^y�O0B�'i��'��'��y���K�Ei�:�	�,4y��,��k�
 *��,$?!�ɑE$
��f�-tڢ���I��DǶ$��O(�D�O��O1�X%�Ht�<���)u�	{���RP�D)Gg�i~��*z����I�S�'�則(i�s��p�`��3�� �&5�	��H��۟��i>I�'8�6��U�:�	�q<R�	�)Qe���2�Q�|�dUܦ)�?)�V��I�� �	���pA��?P��´�VI�� �`�Ц�'D$A�s��?��}j��j��U���]�f�1s��J�"a�g�ԅ�	7ڦ��G��6�^���ǖaCj`�I�	��M��M��n�j�O8�x���*|���i�&���O�ɨ�Ms0���ďC�9��V��d�я��X����������m��:�Zp���OO���?Y��?��c_����IC�hKs��4*�(����?+O�o.�I��؟��	W��D�g��лE��6,�(��%�%��DW}"�'	�|ʟN}7┌2�1��)���yW��'g#�Ǩ~����|zWL�� '��PԀ�rv����^8	���1�Qß��������b>�'xL7�H�OV�y˖� ?M�h���0#w��jve�O�$���?��]��I-�12S���I��-�ub��(x�4�	�<�Cɦ�'��!@��?����`2�8Z��a஁3l.��qu6OJ��?���?���?�����ɖ&F�����)3�����B�+4@��n��#��\�'��������w��3�┴,㪁{��͹`kߴD�f+��)�V:7m|�� �##��9bS�ɺW��r�	��1O���3�٬�?�!�>���<�'�?�vm� �֘iBBDlM�+L��?����?i����dL��8`������⟸хO�\xz�;���[�`��3"�x��h�I)�M�`�i�lO�9B"霈.��}`���a��I�P� aE�:-Z��*�S��������K@�<-����$F��n�����������t�	П�F���'g*!�E���h d��:Z.("��'&7��?�Hʓ4��&�4��0�u"��7����� [[Jhs�5O�Pl�<�M��i�p)�q�i���� 
���f�O�N��ŨA�[L��1e������˃؟ȕ'S�i>���ʟ�	���	r'd|��O��]U���2�GN.4,�'.7M_><��O��d(�9O� � .t���Y���	�t����H}r�'02�|����j�~�	�eV�6⼱(�d�6|�\���i)�I����z�O����<�-O6�3��9���F/�]�XP ��O����O��$�O�	�<	��i��D���'|RA�GbΈ?-�3��L\��x���'!�6-%�ɋ����On���OhL�u &Q�zp����-GH���ʹ~!�6'?)e�֪|�|���׬̢��0wO����V&��Γ��?�pV2P���#��L�����"��?��?q��i��˟��l�s�2S��P�qO�+v�3����$;M<)u�i�X6=�D�k �a�$�g���Fg
�7Qd�[b��2<�x�$"R�gu���@�ry2�'Br�'�R�ћ	^�P�ǿ]LV��W!L�@i��'��ɐ�M��*��?I���?�(�� �FY ����a���tpA��8�)O��DpӖA$��'K~�����%� �;C�I4���G�/{��[޴/�i>	�#�O̒O�A2���.BW�0�/�;q�( jFi�O2�$�O@�d�O1��ʓY����Y�%�$�ۗ蒃�����A�P"�'��al���DثOX�o�|��`��I
U�nxh����7����4�����(��f���h��	�U���<��*"у�2�( ��P�<�*Or���O����O����O�˧ot��� ބ+P��8���.�mJ��i�T��0�'�B�'��O�2�c������ Eo��Ev��2���doډ�M��x���?�v7O�Hإˈ�TR�݉f���x�2�8O���#Ŝ��~R�|2^���	՟(TȪD�t�Y�U1-e��Zeʍ���ʟ��	}yR�t�, Ж*�O����O��2�`iN�")'\��+ `.�	:��dJǦ��4u�'i��	�n� D�F�;��Z7� ��O�q* qD6m]H�S�@���Oh�	�	V  ��IWj�);�=� ��O����O~��O�}�;b�|A`�}���s�� �8k�-���i�s��'� 6�+�i޽��Ȱ x��DF9n�8�������Iঙ�޴`�.�[�4��d\7�M��O|�X*f��'-�FU��ֆV�0��T�|�V������@��ПT�Iǟ����	b\P����INY�!�Sy�|�>��c��O����O8����(O�ư(��Ή��С�IӣWJ|��'�J6��ݦyrL<�|���ϥp�����Tm�� [aLݶ�L#�-B~��m%(�I3�''��4} ~D�UnոgU����g�������������i>�'U�7�K�7Ģ���9miHi�Ӆ�)Yzh�i�+��Ĕ���?A�Y���شA����|��D��"F!�T�8�Ɋ]X���E?n7m%?A���#3к��$��߭�"�J&H�41����7����q� �Iٟ�����	؟���i�
xq�؀
���p��+�&�?���?�b�i9:5��S���ݴ��r�`�
��� Foa)Dfaj�� ךxR�l�Ġmz>Y�O�¦��'�X1H
�n]*�R"h����հ`���K�p�	(%��'N�)�s���U	+�"`:��U8���t�4���vdӀD���'�2V>���B�o���0ĝ4s�e��L>?��]�d�۴b���;�?Aҷ��,��a�nV0i�s�X%}�^�!֦B��+O��O��~��|�$F�@�L�ЫF�v�桋���3�x��c�X�:`�R(BIt�)@M��T|Y8��H�"��Ozym�`��YF�	��M{�i�!Z3X�YV�̪����3���g��vKfӚ	��Ns��Y2���F`�?��'��A"�J�,[��BeN��-����'���y����hZ�2����E�-�<�`�	�Mku���?���?����r��N�' -������6�E=m�Ll�M���x���+GA��V8O��aA�E��U��G�)r�ъ�5OR��`��~"�|�\�����`���G Qq���5��ܡ!�����	ݟ���UyrBgӘ1�tL�<���B��+�m�8K���rrI��P�ص	��>)�iV�7M�e�ɱK�ȅ�Efݺ9^	
�%E�?��wsz����y��|B��OȽ2��*�)C��"�B"��|�9B���?���?���h��n�C"�`7爬
�8Z��@x���Y¦}�3C!?)��i��O��$j���q�g�]�xQ�������O6��O��3h~Ӿ�=^�����?�y3�X�.r<iQ�ɕ5�x���]��Ty�O7"�'e��'A��"=,5��/&��Q�������M�U�P�?i���?yI~�+b����G8�� GlШBXJ-�bQ�`�	П4&�b>�f):� 䰈2â.54ِ��Ҋ��}�d��-k�I�/�� �'Q�d$���'uv�Ӏ��p઱H���?9�V���'/"�'~�����P���޴&��l��-�^�B�fՈ+��Z���NX��v�&���[}��'��'�R�Ӑi�,�"�A6o��"z�T�M(����!� ��T�)��r�m_�d(Q����(C�9C43O���O<�$�O����Ol�?5ؑn�p<DMy�D �U���vf�Cy��'�7�O����O�\m�t�I�|g��Ӏ� ��Qa�L2���%���I��擳 �1lA~&�5^@�A�]9c�N����Ŋ9Q������3��|�S��������ߟ 1�D��3_�,(�S)S1����G؟L�IIyboӐdɰ �OB�$�O��'F��T�։{)�E�E� _�}�'�b��?a���S����1��9AƧOu8B��Ci��U��dT��O�Q��?�t�.��
 ��ec���b�04-�5���$�O���O ��< �iUJHBb�![�q��8�LL�ӉH�$5剛�M;��>��j
��9�D�d�.!!"k��4b썡���?�D���M��O�9Z��6ʸO��	��o�.�
�:��/
�Y�'���ϟ$�	����� ��w�T�[�K�4�G*�#��q��#c�7-Q�-�L��O:�d&�9O>�mz���!��'{�=`GHrOnp���M��i�O1�0eBf�r��ɚFr�����;g�2� v-1::z�\ �ċ��_����$	��U��D��R��-e��)[�И��-SJ|��!("��Eխ�Tອ�u!�2aJ1C�	U�j�٠�)�7gc��r&6�x�IV��`�j��$̕r6��&��<s,9�Lӊwھ0�gf��g���AF�e�$�(mJ�xi&��F�]>u<a�v͐�x����V�1�^L����9��dHӥ�	�2i#�lǡ#ݒ�0mG�)�hQ�+(���[���N�	P��/�	�i�&/|��z�% :�$��l�)7>��I�m���$ �V�^IÀD�?bP+"�:�6�O��DC�^��уÄ�Ɣ�g@	�!�LnZ۟P&���',�y��}"���O.�H)��\�5R��t���M[��?(O|���g��Ο����O���IAȀ0,
��P�4@p�u�N<�)O&ѐT�~�N��IE@(��\���q�d��M�'���T n�-�O""�O���m>�yJ�n�9�ni�p._�rԸ�oZyr���O��X	��̨7��,Q��'l��Ժi����u�p���O2���&�p�	&uۀmy�@�$B��#ƅ��p޴*�Dx����Oм��� B���A��>��Q���WƦ�������|'T��H<���?��'���z�-ۃ 6T�M���d��}b�8��'�"�'/b�P�9	AlXSk�sՋ,:6�O���pjc��?L>��:܂X��d��X�^��4�$Q�D��j>��ן��IƟ�'��)j�A���>����?Z��Y1��7V��O��d�O��$�<�*Of`��@ߒN5tH�c鞼�pt,G�Lg1O0���O��d�<��d��h��ɐ)Ѥ,��F�e����"װ{��Iǟ(�	~�	Gy��$�����*�jd�p�Wm+�k�"��{��I͟��	��ؗ'�,�##%�)���x:�_�b!�G����n�|'���'��蠋}"�M%}��  ��jE�h#��$�M���?�(O2�"�O~������S-}����I%YFl�����j� �N<	/O�h��~B�JМ-��,�e J�* \ç�����'�F]Xэz��M�O2�O��,�R��7΂�aCH��G��W0�-oJyBcN��O�����qo�=�P��;e�����i7&�xӃm�\�d�O~����%���ɧx$Y�#B�oj�Q*Ɯ�Bxzt9�4z�TtEx��I�OF����K;%��W�Vx{L��f��}�����4)LQ��ǟ(�OGB�OZ)i�m[�b4��2_�@�d)�aHJm̓ 
�Q���t�'#��'����;��3��	k�e2�k��扑Yw��D�O�t�O��|�C�5� P�.�7�0�D)� /�Oڜ���� ������I�t�ɿb�6d�7gA;��U�ǈ�q��p��c�RyQ����V��ޟ���B00i�]�u�pa#q3S��nڹY�@�?����?i���?�� �"��䬈�sqPqS�,q��t�U� �MS���?������?�.O����i���3�_5gQ��0A��+�0�O��D�O���<��N�i%�S��3����1�2ѡ���؜�1��ۇ�M�����?��x�H
�{2���cU�d�UÁP�E��,T��MK���?�+O�@G@q�4�'��O"�Q����Z���	��-݂݊��"��O����6a����'6����a-M]�lIF�*@�^\l�zyrj�0R7�O��D�O��i�j}Zct)��n	�~1T���Tp�ش�?���]#vHY�b��� ^@�B0��8oK��x��9K �FDǮX� 7��O����O���`}�T�4�P̂\J|)[Tȱ�ɋ��x�4Sr ���䓎�O� �%E�F���Ȏ\.H��L�+�"�?Y��?��& ���{y�'#�dY�Gk���o@)efy��.��f(���|"a��P�P�d�O����SЙ���M����7�U�A>�=lZ��������<)�����6!�9n�N���b	.gM������[}"BbY����֟���ey�ؕx�Xzf��l���1�aR"x 0�M�>�/O��D>���O��DG_�? ��P���-��&S�z�	�So�T̓�?	��?I(OzH2��|����3@7�Q!��|���B���%�'Hґ|��'I�d��-j�˙=&���������0�Е�ڥQ����?9���?�-O$�����f���'���#��2(b�YQ��<0�0|��!hӀ�$(�d�O��d��"��dY���k)B��ޚ>:�U�`�r��D�O�������_?���Ο������0��������#^
b���L<���?����?�N>	�O��@�P/�t��5;���D!��۴���1!Ϥ(nZ۟T�I���������*1�s&%J�IK��A;�����izR�'Ith��'��'�q���1�S5 b|��i!����g�i���k`�����O��$�� �'C�	�)��eB��A
Ff�y�(H�%����ܴ�QX���i�O!{�K��I�L�;��1�>QԏR����ȟ���5�q��ON��?��'C�4���˒$�D����F�xI�}B��'B�'�B�'[�HB�c�Y���E�FǤ�eF���h6��O��+��ET�i>Y�	K�i�Y۲L�v��hCB[[����&g�>�c���?�/O����OV��<��f�gE$i�~+zQ�w�P+��:a�x��'�B�|�_��S@F_$l\4[�gK��\� �z����yyb�'M��'��	l�> ��O@�*r셮$}�m:��.}�	�Op�d�Ov�Or˓S�H��AE�����ݣ�.8�7J
�'��� �X�0�	��IyyRk��'@��0S1�N�2J�M�!���kC-�����i�	Xy�F�H6R�~Ӄ 19���	��(n�L��� ]ݦ��	֟x�'Qj����8���OR���T��&-6*�<U�Sj�?��8�ՕxBW��h�!���%?��'b:�[u#S���e�@�ZmGyR��(�*6�@P��'���"?��M*>�~���AR�HH&�Lզ��'�8�*�'N������)�F���H���a˞4���M; I��?A���?����b(O��F%��j�H��8>D���߼yAZ-aشyG����(Xw�S�O�Z<ZC��@2��Z�).-��JS+tӈ��O����Zhh�S�D�>�a�y����o�Ԫ����Tf�1O�}3WC�d�'�?Q�'`-귡�<xÔ���T�M�۴�?��ؒ��$�_���DQ�*�R�y��M7V\��@NF
G�J��'pV�R-ڸ���O����OfʓH��swʑ�6s4�xC��u(�s��9��'�"�'�'��ItIܰ	�$��%����p)�Ft��1�d�O ��?��%��tH�-��#��%U�6��Q��4�MK��?��r�'�R�8,�۴qL�S��W�l�i���U
v��'�D�	zyr�'��}K�_>E�ɍw���0��+a����$X���%�޴��'H��'G
%���-�ē {҉bqe,t.NM� 훖#S(QoZ���'��K�=��S�L�	�?�X�(5)���/��M�(Oj��Or勖��Y�1O�
������>>��J���2����?�`���?���?���2*O���*� i! �Zﶖ?�8�۴�?�X��,�x�S�H�f�����@a�YK�/Zj�4�mZ���{�4�?���?��������_d�B�Y���Qa��6��$�����O(ʓ���<���,�Њ���+"?����L��Z<�58��i@R�'�҄�./pO��OX�����	��ʄ(䩂 ��XB6��O�N�`u�R?�ß��۟\2`�˯h�F��R�̜Z*E�p���M���(�Z��$�x�O��|�+Z�#�pqx�!Ӻ6�b�q!�ܡx�0�6 �%1�����O���O<�7x*� ��Ɓ�r"�)aox`�r��&��'���'O�'���3Ԃ�;E
�z���3�KK78Wz��0EV��T�'���'�B]��S0�ׇ������$L��n�d�&�JP�%�M�(O���<���?��c)d��I��a怌8��`ƋC>��Q�$�	����IDy�e�$~만?i�`�!��\�.H�G��pj�v�m�ȟ��'���'"�I��y��'��L4g�(l��%�1dP<3у��ou���'Q�\�8{ �	��)�ON���U��R�6�c���(fB�`D�_}b�'/�'���OZʓ���Z�e,J�����P���L�M�/O��ّj�Ȧ��	������?-�O�.�G�4��(�\� c�CV� ����'����yR�|��I]d�n�a��%v_0,c�;���M�(5�v7m�O����O"��n}"V��C@�|863�進-�.���]��M�����<.O��$$�ş�gL��52|�/$��L�
<�	*�4�?i��?���9=��Iyy��'i��K�-����1- �X��`�OϏ#�&�'3��'�иq���	�O����O�h���`1"<8��?s
�i�EæY�I�:S�]��OH��?!,OJ���4 �㖃q8Թy��G�GH\��iC-�<�yrX��I����ayA	b8���重V��]S���,t�+F�>A.O���<I��?a��M�=��	�*9�9#�M�hʀ�p��ZI~b�'��'�BU��Ee���t��ki4Ո'�}�d�u�?�M#)O��D�<)��?��~�R��cƣ]><�*�@�/��k�঑��֟��I��ȗ'J�E��N�~����W�D���§T	|�>�z�@VѦE�I_y��'��'�`q�'�S�? 8���EH�.T�	����DmR��5�i1B�'@�I�l���󪟐��O���At����D.S�Q�X%7F@�`��'���'���ɼ՘�y2ӟn�j�ƀ/���1t<Pv�xR�iL�ɥF��e��4�?!���?���P�iݥBn�5l$��0���BS$�c@i���$�O� �:O���<��l�9M�6YY���1>�c!����M�n��D��'�2�'��g�>!/O�i��aj��h��aF�X�a�H��
�y����Vy����O��Ps߅i�prD� N�QdVȦ���؟���1�,�O�ʓ�?��'=�E:�D��\`��V�e�4`�4�?9���?9����<�O��'��������O�.�i��ݠH>$7m�O,�)��Zu}RS���IqyB�5)�`�00'iN c.ڭ�S�^��M#��jF��̓�?����?��?+O����=v+v)���L�d��Y�@�:.���'l���'m��'
��'U���Z7�-Z��}�!#�v�L���'��'��'�rP��0�݌����%MZ��7lYq���т�H��M�,OH�Ĭ<����?)��`���L�x�z��ۮM��+�eO�e�E�i�B�'�R�'��I���񑭟z��������(X��#�1iv�iz�Q��	����QZv�B�D ȷ(�IH�+OV�K�̄�^�7��O��ĩ<�`i	�sI��џ,���?}P2�#��'�y������d�O2�$�O��?����΋z�TH�"Ğ�H�l����ӄ�Ms)O���r�A�u��ɟL���?ѓ�O��%7��A����`yN)�3J��A����'iR�[�yb�'m�p�'z>5Qa)��"WjAs�$!5鼹n���.�+�4�?I���?��'��Ihyr�	i��xA G�^�`4��r�z6��!2�<����O��Nu�rY1GA�S�@�`'��i.7��O8���OT���!e}BQ�,��`?Y�C�M���I0����QC �_ۦ�%� :�ok��?Y��?��gʰi+��X$�P�tm�TQ`Ĵ��&�'��I���>)(OD�D�<!���2��:=i�l:B�Lb�\P�	����I=5�D�I۟$�	ӟ��Iԟ��'��Z��Ҽ��j�g4iy4!	a(���D�O�ʓ�?1���?��:2w�}A�X�E��V՝AB���?����?)���?i)O���a��|*��Q����{5��r �idFVԦ�'�2P��I��\�	�8F|���1s#�>J� �Ǆ	\/��nZޟ��Iҟ��	uy�j� �'�?��Z���1��
X�/�8؞�l����'���'����:�yX>��%�\���1ZG��?τi	���ȟ���̔'2�"W��~����?���N�Ve��
T:R�5F�:n���Y�����,���IGP��j��'��)�+���G�s/\Qh�˖;�vU�ث��� �M����?���ڷ[�֝3x��0�ݖ ����T�ESn6��O��F7����M��'q���014�.� ǃ0;���1�i7�(�։}Ӟ���O����ʼ�'v則�d���<�v��hL�tn�ٴ8�\��?�)O��?���-L@���ID8q�����N��Msܴ�?I���?�a�	���Ixy��'8�d�6�����&58i�ᇏ����'�Ɂs���)J��?1�6�,�a�^b��l���3v�b}jS�i9��<m@ꓲ��O���?��G��u@6��N �4�$Ѳ5����'�v�c�'������	ڟ(�'��� vH�V���ǀ�>���U���`�����O�ʓ�?����?�'�A-�fa�u��+�l��lF�2�Plϓ����OB���O|���v�O#���L� �0)(���VV�V#��M#,Oj�d�<)���?��� 0���'ʊа��A`��@ b��ISᩯO��D�Ot�$�<����k�Sܟ԰��>A��MsU"��|�$��Kݚ�M�����O��D�O���9O���O2�M�K#���V׀5����iO֦����'j�%���)�O�D�m��	�07p-#�eѽV��Q�&!�m}��'���'�Xy�}�����\LL�D�N��qɴ���I�/�Mc+O�d��K��E�	ٟ@���?���O�n�1s��G�IY������e�v�'���
��yҐ|�iS6�i0탹`W<|��UG�v�I�-��7��O�d�O��)�t}"P�x���A&#���y�lƣT�QS�����M3"���<iL>ь���'�� 9�e7^�4�7A�,]4�u��x�,���O.���2V.'�H�I˟�r��ʶ](�vY�&J�.Ug:-�>�u.S^��?���?�+69!T�U�q��t�b.Gi���n�ݟ��'�P,�ē�?y�����F�{�(̳d��T� 0���d}b����yBU����⟼�IUy�W�ljH�z�ɸ\H�@��@���&�4�D�O&�d0�d�O$�D�MB���)S.ֶ��ɋ��X�@4O0˓�?����'#�@P"�3���@�ɚ�O�P�7iA�vU�%J�\�h����'�l���|�!�z?!U�6;$��ׁ���8d!TjVl}r�'���'�剂S�80�L|r�-�[�2d���,�4��Q*(��f�'c�'Qr�'�dc��'��|X{��CY�0�b�ɍ	���m�ğt�	]y҃�,�������2s�F�3�@�B0Θ�E z�����@�����I�f�܌��i�S��B]���z� ͮ���5������'���Fx���O��OL��%�L(��
����`�!;�X�l�ɟx���"���Ij��p�g�? ��0$%�5o�*����&+e(0�G�ipv}��yӞ���O����,9�>	$ř�E�α!P��#�Ԩ90ƈ:]���T��yb�|��I�OH=���D"o)`)KÀ�"pldZa�զ}�I����� ,�J<9���?��'���@�Go��x���<]����4��Y��ӕ����'�"�'6��gF���p�i�
U�]^̍��c�����0L���>a������gގ_O�1x�M�8F�ԂbA^}�.�f��'���'��W����J=6�$`��L�0��\`��з^�F1x�}��'�'��':d�X��x9�����%\�8�1%��y�S�����X�'��������^1+��L�)E��(���$f���'���'U�'���`���ʄ@g���7�_8	������D��@[�6�iQ�����&]B�~B��(�H�p�����b�B1b��M���䓝򤅤4%b(#��x�d�/Jx4c��O�P���-�M;����D�O�##�?��	�0�Φ}P��[�p�� ��V��,���xR^��3��J!�c��eNL��q�G6���#&� *��o�Iyr�Д�V7m�OX���O��j}Zw6�X����
E ]�F�/R.���޴�?Q�b��ϓ\��s�P�}��O�z��.�-z���R�E즥!+�=�MS���?y���rS��'@�� b���o��- P�H8<����gu�D��;O��$�<���T�'w��$�رP�b��m��
2��!G����'���'6��0d�>�,O�������%ʌg��i0c[�8��ɰ	o�F��<9�D��<�OB�'���>L*�� ~�"S�C�IF���'��\�C@�>�,O~��<����D�Öb����7_[j��1�̦E�I%���	ϟ�Iɟ��I۟��'4B�*T�� �*8h��S7@��jB]�����O�ʓ�?	���?�0�L�_)��P�rL\��T�L�x`����Ot�D�O��*�`��C:��0���gO�M����.\����5�i���䟬�'���'�ҭ!�y��O�<��8�G�pa��q͘�U�<7M�O���O �d�g��ួpc�'�bk�c:`���T�RQZ`���cP6�O�O�$�<q%��I'z�U#��~�N��)"R�iC�'���1.4�H2��2���O��IK9ye�,:�{���b����	l�T�x�>�,���
�K�e�������;zt�m��d��Qd�<�	Ο�����?�1B�0�-�9gg�P�Ӧ�4nRr(lZß �'2X�h����`�^:��:Ǐ��L��lH����Ms����?���?!�����?�(���n��6���.<�\�C��GI}BF���O1���ڕ_���H6"��8�Ⰱ�3%�^�nZ埠��ǟPi�&ӕ���|���?�bH�xzx����s��@y��W��O���'���O����O��� F*GZ}��k@�u�"u����@zE�'�@�'�?	H>���R���àj��L ��D]�'f����O����O|�d�<Q�"��	Ԍ�t'���bT��q�L.���?�����?��0� i+*ѐs�1�
FERV��I���?)���?�)O�t�3Hfj�)�?3�4�E+ �T�!k�>!���?�M>)��?�pO�w}�I>���r���(u*�4A��'�2�'5P�@	�eP���':|Lt��
S�`��h�2�]�P,�ҹit"�|��'u���*��',&	��g�7OB��)�G8����4�?���$�:�Tq$>��I�?I��LË��r*&@/�J�$� �ē�?9��Dx����6&��2!�!��!!M�e�s͗�RHE��d���ǆV(��Oa(�O�̩(p/���K�@��"%*O�\�5��f�^Aq�A�/*�@��3���Yl���vk-��B�֍0G���D[�u���1#C�%>�0mh����E�0%XCH�q<z��C��d6�xq�]�?E\�{%�)7 aۀ���E��FC�]d*m�<Sx\���Z�#+nY�S���,-ifm;*��g��DX�����Ҷ�'L��'�2ft���	ן� 49[谵9�j�6E��1�q#�=J���DQP�Y,�����(O20�D@�?�p��'D�%L��E!���L� ��+ʇJb:�Å�t6��D�'����6*��l��E�3@� }�d�:�'Fje����?a���<�t,R��YH��B�:��e���O_�<	��7F��,��fn<x���4O���'��7���lZ�� 9A�Y�?��+�e�Y�\���П�����P�7�ݟL���|�G�\�O-h��I�'��c%@K	C:d��FD��K:XX����<i���)H%z�i�N5c���	��S�^b���N�x��:�����<Ѱ�N���I\v`�B�!F=S	8L���o��D{2�ɴ3�|MS� ̖�.[��^�?�B�	�[�j�2&��#G�٢DdG�M?�牔��ĵ<a��_
(�����O��T��lR�`s°[v����� �(O�2�'���Q{b�0�%�^�D  �L�O�S�h n���A�OΒ��%���P���<��M8_n.��&�@U�N|���ʺ)���f�T8\6���S�':�0����?q���#^���q;��aOP�S�@��y��'�N�����e��Ju���0m|������� ��פY�
јH�`JC�rB���0O���Ήt}�'��u�L)�������7C"��%�^�ER�R�=B�H<��d�f̮�iW��7"�`h�S����'��2�͘�o�~�s�gC CQ��3.49�R���)˷q�3�#�O?���~꨸��M<.5;�mO1;K���n�O4��4?%?E&� j!�Fv�*$2�N�.#�: �2D� ���l�D҄��B�[6i54���V��<���'nhd�$hx1*"�����	 f�8=B�T����Iϟ@��%�u��'�B/�_v:�a�/��BbtQ�+Y+o�<����܄+Հ�!�P���hOV��UDE?�3����
�f4�ЬX%^,�ty��+D�ԁ���
�?���ɖ(^��X��	��@�ie.ю��	�OM����O�=I(Ojdcs�F�";tP��oė(Z8=rg"OJ2$�$3�6��'I><�x9H^���i�<�����p��h�
V;��9�ѨD�8�`!���B�'�2�'.�ɘOr�'��e�f�%�(dAl�X�ft�s�P�4Y^����ߩ�p>�'�KV�h�zva��l�;�.Q�r�0��o��E���gW0��Y�ቬ|#l�$�O �iP*�R�2��E勿_4��[Iئ-��gy��'P�O�	;$��BG�7tV x��1W$��>�ųj�|��)�#:��,�2뒼_0�d���bܴ��D�1Aʄm�쟠�	v���1C8Q��.$Qp88�	�ap�P��'��'��yU�'I1O响2<ԉ�&�/�"}��%Y�C���<&�T�O=��	!CM�ӓfʽ]w �@���T9��S�X��b D��M[퓞J��B�I�����C�ڻ^��1�&`�P����d�J�IPgܤ3���94|mɐ��![�~��!39��4�?����IO�a�����Oz���o湐E5QU�d�Ua����ORb��g�'Y���`�0
Z���@H/`hE �E;m�"~�ɗ�:-���ܕz��Up�&k��|�1����<E���/��B�?G_`uK�����ȓX@PRN(J�.�Xi�#e�lhDxR)�S���'h,�����!A;b�qsm�����'�v���!7�r�'LR�'?`�]����;^�4RgQ�d��qc���G�������DK�OP��W�[1QX�PZP"�#	�D��L��}��ON.�M�ehϸ"%��`�K �~��,�?�	�S,� �
8����~����ȓw��Hp�I�i2��@��V/G�����)§h�,m[G�i�T����L�(&xؒ`�S��]�'���'�B��a���'i�)�	e���'�
 ĂV>1��ȇ��!���[�]c^|�'�a����b����դ��!�d�(
�Q&�X�I!PgO>�d8��	87FI���9D��h�	�>O\L	�Y�ډK�7D�<��;5~�Qz������w�D��}���r(6-�O���|:�������31~N������,�7����?y���?��i�6N�BQ�y*�Ȑ��$]֌�R��b�������x���=��
�韲��84D_�(��<��M@�l�	u�����a� �P�&* ԩ� oR����?E��'���"K�0r?j���9��(�s��'��)ئ�u��ܺ`,��e|�y�'�zQp��|Ӛ���O�˧V�\`��?)�3B$�ҀmOM=��4͇'����S��6�?ٌy*���j�.�.K0��啾LsJ!�D�.��xGx���'�2,�c�	̐�zT��2RĔ��ó8r"���O�4y-�4<�P�)26 ��"O09���8�@����>/0(p�%�ɺ�HO��&f�qxRJ�
p���.��T����ҟԓ�i̗m"��I����I���Xw��w'n=	��ؾ>ɨ�eB�3�$�K�'�.YB�f�*$������<�Rl;���y���)�Kk��$Ӳ_i4��BB�`�̆�ɴU���2�9	����H({� D��. � ]��ş���t�'[���Sd�WG2a�l�(�*�ږ�=?a���<n��ՃC���e��B	܁��ٴu�Ɯ|ʟf�N.T��׽is�\pA�2R0t5K2�3��T���'6��'3�m�8kr��'	�iޓ
�>9��A��3��Sc�W��EÌ�0��P��e���'5"M�7Ɗ�RHE� ��d����D+ؤS�̘�kR-:��8��' �̐��?�B� ����@բ*�2��d��?����s��xg`D�H-�1�P�ZQPK�k*D�D('c�0+L�F�)A��St��ЭO��Q�ڠ遺i��'��3� ��S��*p�0D�T�#� `�`�M�n�N�D�O���:���4�|Br'��(^9т�	2�r��^�'��]`���TS�`H�r��iQh��'`KpQ���G�OL�}r�lE�<�h���"Ӎ9��h#���W�<aG̎n�p,�!�G&uNK�Q��RL<��jSu��h�c�2���qfC�<!B*R�1=���'v�S>I��oß���şP���Q�qdd ���
6i�H�b��1h����I@�S����[�Uc࠙TEp�QFLA{,Ȧo=�S��?��x��5��e�}��h�̗~w @��֘���"�W&?o��&��z7<�s�$Ʀ�y�MLh����yq���GO��O Fzʟ��AĊ��\FF�@`ʗ�m1����OR��=r�Eb��O����Oj�����{�Ӽ�D!ՏO�~��+&�����]A?a�BNx�T���S>	���;�Bv��h$g��T��
0�O���T.�(U?� c��$tR�Kr�OH���'��{ҏ�t�=�0#߀T��kG�2�y"EQ�y�Fl3��T�n8��[��"=E�DC�)����6@� 4�����}�$c�)���'=b�'�����'��5�L��g�'�B�+�f���+T �yg�2�p>1�`�Hy�A*^(Tx
$-J� v���0�p>�5��T�I�7���i�"R���]u,B�6y%�E�c@�$}�*��#�+B�I.8�u�@��!	� UKǦ�	JT版��'4�q5�}�
�d�O>�'j_`�� ̈́*b
1�ܾUÞa��"�	�?����?���=^Ҕ�S�|��b $�����ǟ�*�h��T{�`s�Y�H�Q��ȧ�ɂo��ei�G�b[:���?IA�]"^� �`��B,�J��.ʓ5��I��l�Iğ�O���Q�5*s8ij ���x��\C��'{�O?�	9~�J�����d��ATK;X������_�I4�z�!��B��#� 	8B�D�ɠ�2���4�?���)� ג��OB���#@)VYS�M�A`N�:���r� {W��O�b��g�'G��q ϑ�A���gb[4�sD� 1��"~��.+�ε�W@q�ղ򈔆E���"�\ڟ �<E��*H�*3(3�<��W��x��a��r5Qqj��*H��ࠋ]�R���Fx��*�S�T��8A��ؔ��*.�L�+�KC ,b�'��8
!	�����'!2�'�N���]�T�q#�@��14~�4�O�J�8�{V�iW� �� ��f٨�zF{�E�$V6|UoԥH;�&�I7��o>�4=�+κp.P�aޟў�pR��9p�Ԣ�k~�zlb楟�+���O`�D�Oh���Oe��H6־9�p�*">��
�'��I���1M����bIҸ~�ܻ�''�S��[�L��̎��M[�j�@Z� ��ȚkTj$+���?�?���?1��Z&����?�O�����?9���)h�:�*S:�5ΏC8�tiδ<���جq�@!*��H?H �D��w8�< ��OF�d�&��`�T���Rf��4e:�(�'�0�	q+D �����+&���	�'M�"D��_�l �L=����'�Jc�|ɕ(ͮ�M{���?y)�@�!�ы$a����MB�f�8����.]�d�O��$N~t���A�$,d4�捃��'S$6=�'.�.[���'���u�v�EyBk�jPv5�T)Z>5^ȫT���Z"GX�ܓ�Y�u��yJK��(O�@;��'<��'�BZ>�W�O��`�gE>w ��0�+���|�?E��'+б�p�ǋg��3Q�Ͷj7�)
���'j����-����-�eqx�ˊy��'��y"�L����R���Q�4��E$���y¡�4h�AC�Ϡ ��p������y���i�� �*K��@Ȣ���yB�T<y�捪���%&�)
g�_+�yr.��Pty��&KZ\�BÌ��yBoV�K�`Z$��u����w S�yb U��h4�ED��n>�E"�"D��yr@EIp^h����!7[��H���+�y�%�Wr0dI�D�Ѓ��y�D�2����,�O�ժ���,�y�m��d�3�Z�N�H,3�&4�y2NP�=�*���KZ�[p����y
� ��+r�6�*؛e�ߔa��d��"OpYa��E�'��n,0)r�"O��CDb�����z�&��n�HH�"O����$f��8#%��G��tW"O��i��fɫ j�/+�bf����ybaP� H���׆!"XN�Av�Ƿ�yr.�-�P'�X%Ő�!�B7�yRO/T�.e�G��
 �6H�5T��yr ��x|8ĨT�̛rl�t�e�E��y��T2� �:�j�-r�ha	���y�� �_ �\�+;hRL8w ���y ��X�;�xʴ�I	j�x0��'���qb �G7�q��_�R���'��h�>I��9:��U(e���
�'���1�ϩC��m�(Y�0)A�'�8]����\�����R�Ze �'�*����30���J 6&e�'��q�A�f:�t���V�*�vI�'r��1֯P2��qc E�(p���'Üdd�Y5p�!�N���*�
�'ն�{a+ŦA� r���� l�	�'~AP�םQ<�=JbÃ%FU��'��|�W�\����j&E�t�i�':R�h�YT�4��)��mԘ�9�'ƨ`U�Jf���)�. Џ��U��>]`�M>G�C�_�8���� D�PdK�y�:X�C��*XB��T��p�S�O3���%�&_bl��' ݢyx�1
�'�f(y�B � \�p
wɆw�^	�I�ȡ��O؞,)��D����rhੂ�%�O�@;1�e�P@���M <{<ؘ�J�
�,��"O0iyd��Z�c`jE�~10b���C���D� _uDN� g��4�-'��yrM�9�p����.�v��eh��~#�z��O�>�� ⓭B���F?]H��G�9D���� ՗<���{��� l�U{t�$�$��E�a{� ��&(���ύz�4��R2�yB�	0�i����$�x�beN�y��ߣ	��b1���"Rq�a���yr$�7C����O�NC�	A#W.�ym�R���Pe�]=FD �u铄�y���fs�2���9CDP�u���y�/R	+VT�d�N�6��(���I&�yr��\�
�Cܶ(Q4��@ƀ�yRfD�frm�0���Y#���yRC��~*����
����B�T5�y��ٚ/ȠJ��
b�ʵS�$׺�yJE/d�����Y|QKG#���yr)�QQ,Q���M>v�Ц���yb��N�]���G�t��\��iU�y2�O=Jp"��T'a���ic��y���*mp����')��e�h��y��&�$�b ����T�DE���y�&��]�t���՜��|��@N��yϕ�K������؀���� �y�_/R��=�G^��NX�¬I3�y2M�!niPm0�fԄ��,���L���=��ʀOA�4��n��(���(�j�3�E	T�d)��y�<+Ag!�\��(��X�.��?��+և<�D9��Iݔ)����$j�*]tl)�"+�}�Q�l٢)?ڧux�m@��:Z�|����<u�,��4�&�D��'�(� ( �Id�iI���	�\���'	mb�}��O>�`7`� Պ��b�50�Ȑ���Of�JЭI�.�hpC��{x���c�ʿ*��`���PGm�<a�'x�O�a���Px��@�Q���� ���E��p���b�9~��G@9�OH�c�w2ʘj��جR�Xː�C6�<�'���fz��ɑHq(E�Cѡ=�ڹh&�ɞ6sX�I4���w��\��C��~���&��8�Р���ḑx7�O����~5P�jG�K>�V�b�%�'K_}�N�qXi��RƯ
mhp��+⟴��찟ф�^�N=�<0 �4e�eSré�T���@Bܓ~��(� Hҕc�E��i@PGDFz4AZ�*�=� �� �4\���a�O�u/ �5�m��@�CCT/��O��͏6ԊqV
ų5�Z�r�xb��#떴:�ҡq�J�bFZ��I�c��%�×m��c���f�x���2�N}��%V
&X�~RdD�~n~�(B��Bz�d��F%���Ǩb��|b ��tHv�Rh\����+ċ�7&�z H�l��y'Z�!p<�cI�
3��é��0?�TI��B,!@�X!)�Fi�R��5wPZ݉Gn�F\5��l��%�\r�ݍX��b��IiFh�V��7�Z܋Cf����׊��Ų	�e��H0��'�4�J�S0�7%��Pa���!IF��ק��-��M"�qԇK�w�FH "R�Q�)9�(�,'�8�{�e�4Br��>)���2P��X*����MD�<�`/75�����~PD�(��?H~2Q��H
\i���A\�BL���T� ����3aިC����ȫ-5�A(�#(�OD(p�\�)3$i���HY<�)�G�"W�T�6K���<��B�Fp�)s�D�I�)*�iӢX�� ~�x���	b������LT�%O=�O:��'��9Y�2lr��I�%&Ҩ#�녊h�� �%�c0���L
U���Q9O�E�dV�"�L�SC��+UQ>�C��O�� �"�v��lS���"�d����7�Bd�P�_�i�B�aP��lvr]$Տx���C�:x01�����5��D@�{T������Y�Я8Q�dJp��7+�h�B��K�
�q���j�X�҉*@C�$* �7~��eHt��kh�@��[�F���E�`�W���}��PA�	��8n,��T��9������SE(a��O�DX1��Y�"n�2Q�6���@F�7W0��i��V�r��:d��,r��V���+ĩS#^������@X�t�xԹ���H/��;��	=c��	���'?�	�Oj�x�C�Wv�Cӌ�Q?!��H�9슴����&&Ř	ȵ�O�'�N8i��L�r^`U���A9�U�E╱b@���p �(~������E6��J� !��K X�m�TlS����D}����)vڄ��ރ`��92sA��y�L�%��JB�w���Ɂ���i�څ��Σ <�80�OP!��@)?�]��l�IKbere�Y�
������8��G�`@���
�*!�p���X&_>E��T;�w����B%Sb]h������9��MH���ƥFm�,�F���yjņ�=�hO�p��H�Kx�Щ��֧>Z�ca�O L���@:�|<Ӓ�ؕf�~����'���2�뉶D�5��܍m�&q�H#64.��`Y���X�GH��?aG�	K����S�۬U���zXC�'�^Ěd�C$q�Qr���H9�}"	B�;m,�y�O⭡�A�dB�S��)&
U�<̬�C����59᠎2!"�~�)�:DyX�fJ�$^�);p��;R���I�g?��Fɡ3����I��?i��wOF���a�	�l�#��ʏz���+�'�~�sR&��m��������MK�/?�ky�H����u��Y�D��2ޟ��d?)"� �qʹ����(�Xe�l�'��4Ѧ�X�`i��k�)2�I"�*�4Y������E;@�P��H�zw�&�?U��j`� j�(bU�^��OD1[�E�:N3�91�0��Ӏ^�p��ř)MX�8z#��&4"��ɦl-}J?���V�H����E���y&�<D���LC
8�n	!	n�\���)jA4����0��Q�t�T*wMBO?i��V����03��-gD�93��Wb؟�H����*��!�Gď��>A2�*6�PȢ��:����e�c�ʡ`G�:� D}�b��&2c/Ϯ_���*������O��2�8�v�@�F1M�Ԕs5�i��t�ԅ����xsՏĄ,��,�rB^����RN��J ��e���ϑtR�'��-����?<4����X	gUp$�M>�O�.i)�h٣X^-A3��<C�Բ
�'���`f�HJҔa�
P�H ���T��*&V��� E)��~���B@���1��A!w�Q<����$���(�Y �'��@#s���d,�����y�0�A�gŔv��I�,�$��U��d��+	+~�*%��H.�I;�l���i��Iu�y��ɚ<!��?��k��As&�����f��
�FQ[�ب�/
4J����L�J�����xҡB��į*��%��I�0��R�@.T�^��V`�<p�*�=�T�VL���;��Wb��0Lҟ֝&`���2�X��a��3!"B�	�\hѲ�ӫ'����ǋ�*%R��ĕ6m�:�xVCY�8<�P&��L����ţn�� �A�ɲ�&e2�d�VstC�I"GU
�J��'a� �b��9�n$pP�P��^p2�
&��-���6�B��	�F�����;���u� �0?���ZINZ2TѢ�����7TD�4H<1`�$A%�;?�Iy�e���4���or�cd�G��=q��!o��Յ1]T�z��v`9��.�6AX���#B"i뒁Ҵ`���>���0D�� Ԡ�pa�1�]qfE*f��GE8�?���5gFP�`2���<�Ԁ��a�3��'e���ݢ����zs�]q�j�J�`��T��!�����$�P@S<3�~A�(��M���� �1Od��g̓!*\�t��(2i%��l�1V��h��I�GA4[I�qqǋQH80x�D�����%4}rA�$U�� ,|z�*u�L�/ (\8��%xv㞼��ا�g�"(tjH�H�Rw:+AH@�H7D��nܓ����
�cN�
vG�#�O��ю�Y�(��Uy;��"t�Iw�xIu�%D�x8Nպ+i�X2R���=�`�
��b�Љ�%�W���;bQd��`�J2"(���"D�0q�Ö���	!�ZAϴ!K�!��xD@.u[h�"�;˚4�1��z6m
�Pl�Ob�G���`S�P7��3��
�R�c�����&6Zܬ;@�d���l�B��?J`��%�^)X��p��
�%� p��:�(bd�.���Od*��ɀٸ�����,ϓKS��w��KhE(0�p!"�O6D����LE�L�X
�6�h�"*6�I
S��DO�c"qO��ʝO�Nt"���
<���`�� ``���'/*1H�ID.+1>�2K�%(�� �딙`���%���'*b#}n�:X��|��d8T�hX��.A�������Q�@��y"
(�� rL�
�XCs�F9�yB���پ�P1MV>��	�y"�����	څy�"쉑J�24���e���!��т�>�b��|�8�Se�l�qO܉�2B��0<��HB>p.Ta�(�f�0��#"�AH<��3�����L��N�Se����qO� �m�
^���GB�\=��X�"OZ�k��D�O��6�$<��f"ON���m���T�*$�yp"Ot�#�.:=i�Dl/_�0�"O����"H�u�@��H���Z�"O�-�d��7�BK ��x��LY�"OTA�q�A�:+�<�&_�,8�u��"O�I
���7� 	� F۽A5dK�"O�����=�2a o�55�["Od��Q F���2�̒4B'���t"OT=hd�_�]^�M��Y��:H�@"O\�SqF(m���E��4��	�"OtLs��ԑV��놏8=��A�"O��b5#^0yd��[�d�{xLi�"O�iI���mh"���A�r���c"O��x
�?.�b��7�L�o��#"O�:���>P'����@�&T,ӵ"ONu��H$ �U�/p(؉�"OJ��cF��s�"�.e�Jpi�"O}�dHU>FP�E��\�|��"O�A8�/Q�0�$�]<�'"O�	��h� W:��#^N��!"Or)�OޣynV�:��h�Pqٔ"O"�T�8I���J������ �"O�3Bh�u�\Ae���$��={0"O(�R %��z2����AE��c�"O�]"u�Rm��,9!d�)���p"O��%��+{���r[,M��Ip�"O8��'�!n4�A��ۨy��e�!"O���ϴSW<[q#n�N�q�"OH�{3� ldA�d���}��S�"OK�U	p�1�)�T����M2�y����lp@j�C�v��b�ɸ�yB.�$'�m#Vn^;R����"��yb�ԑ!4F�3��E:� �YA�����FC�e��  �p��ծ��H��=_4�(�4RKF��7�X+C�(��S�? ��K#\�֤��4N��I��4"O P"�!���C�nɄ4)�]�d"Of�Qǥw,޴��M��'A�MjW"O���p���7���S��*#(�i�`"O����-�� \8�&l���J�"O�	��E!�R�ҥĆ(�@��q"O�a�5h��M�0�η5�Z��"O���Bu� �b�D%�8s��{�<Q'b� WH;�A��O2�a�P�b�<q���'I���f϶b�q���c�<�g��=/v�� �K4So�yJQa�<q�M��+.�h�� Q0eV��#	XZ�<��ށɺ(�F�?j�1���_�<鲅�4K�ء1�D��r"nA80�\]�<�N
1��qZ�FE�4?�����V�<q�ś�G�"d!��S�f_��C���V�<a1�����D��c�H�+��TU�<�V ק4b���7R�0i�R��\�<!#���8"05� �J�~������B�<��j�|c�e��4��)����A�<Ɇ�[$U��*�c�)�@��؇ȓf'����jW V#@�P��7���ȓRv��CVc.�h���6Wrȇ�V�P�ku�K�	G�p!S�R�E�d�ȓ~��1Xq!�q5��y��'�T�ȓq�<�b#�$q�l���@�x��y�ȓ*~d��(�N��iѓ�P"Q씇ȓP�N�s�Cx��b%���w�����̴��+@�G�}r�m$D�n��ȓn�ěv��HC��Ip ˇ��t�ȓ0������iaj�	���`!�'ў"}j���<vl�w� :*���&�w�<���ٷv���i�cQ�o
�i���w�<�d�N#.�tܚ$	���`i��r�<�D�X�h|���<F���#�H�'^axb�\�J�\��E x��
R��y�c_L���h1a�%� ���ʃ�y2�v{�|["&�?0a�	��ybd�2r��sn�����c���y2l�r�m���T#:����L���y"FU��DM�"��?;�Kķs �͆����6@�`G^�i�H�0|��C�I.w�xp�˳	*���Rl�$�RC�	�cw���4 D�Ta��
�q^tB�I�Mm蹱�#E��SF�E�n C��\���aJH�zf ��mD�J8�B�,�bK��[�T�5eĦ��B�Ɉ$W�� ��?Uo�a嬁84�hB�M��0��ܚ Oޜ:D�B�	)mԤș2���H��q%�^�B��>NA8�j��(8���3ǔ���B�	,i�<��ʉ�2h��8F�Ѯcf�B�	�:�,ӄ�<�����i̴a�C�	C!��q'HԄ\�$����2�rC��>J��Psc�4\�R{f���FC�I}|8Y1�H��2i��R�kBC䉭R9ȡr"�Q�{ ۟k�F��hO>1���"z�vDHbd�! H�94�&D�8��G�${�tITM�)*���"c/D��q@�W�p�*�/ߥ|ʄ��  *D��P�
�7]��tq4��9DTP��$D�+!��%(K&
�?5��,;c�5D�8�"�S�2����c�W<2�J��.��p��(+�?s�R)���߈4�TY:�-D�� �آЃ\���p�y���"O���RE��{+��!`8d�����'0qOx��T�[5*���a�n�O� s"O\�!�ˈ�K��6��?~�4�ʴ"O ܡ�o��_���#T���BՀ�Ȣ"O��6$E4G��(���S��#"O����38�q�CH�ȡ�b"O`����ɰ�L�s�L�8��] �"O��@3 �0l$���y�ٱ3"O�)��ؾX2��)@�U1dL8:C"O��R��/��@����yJ�p� "O����Z|"�������X�W"O���卟�7{�U!0�� j|����"O,�m����X�N[�@��E S"O��Pե�Ju�6�B
B�H4��"O���;=�\ytk��c���C�"O��@n��r���qa�e���1"O�HC��&����[�$�b!8V"OL��4�! s*�bN�R��q�e"Ox=:U�_�q8���cK.2v�s�"O��3Vm
��>��sS�c�1i�"O2��K9q��)9OC����+�"O�0ڀdQ2hp���D�m�,��"O� ��lљ>@aD׎k�0���O��dU�7�j�qH�%N�c��/�!�dYU�����Κ�?��X�&��)�!��
��x���B�V<�{ aA��!�d��W>�Y"2�ܘY�X��͌�_�!��F�BYr�˷懩1���q�P>4=��)�,��IK��
�-`��;C۲(�RL�ʓBּ��[��P�� Uy>U��r<PU�oη\Ixp�OT�/��y�ȓ&<��k�� o�^���Ҕv�4��ȓ#��!�.�`B�l�U��,-��J�Ԕz�GP?}߂��⌜Ezd܅ȓ ��#"��MvJ���>k4��h��Z�d��ۈAK0�#�%Dp�<�P�N|@�j�B:��`���l�<�qOW&�֘��ω�kp2�Z���p�<1F��C> k��D�7�桪fA�i�<I�%��⬐!�������`�<���V$h#�S�Q�`Q�)O_�<�Ah�:ᘥ��A�F��Q aNv�<�$h�&��C`��'��Ҳ�n�<q�Q;PI4�!D|��v$�`�<9v���*�ctc�3�2�`��[x�<��9<��r�� ^����vĕr�<Ɂ�*pK�MÍ!m��"DU�<A�U,4����Fd=Z�k��SQ�<Q��L�r�Եz�1f�*�cV��O�	j��8䌈#o�`�*eBQ5(� ѻ�	"D�0�ӱ	�2h2� ���=D��0Ej��x���%ہy�� �K/,O�7->���2�hP����X�q��/n��C�Ɉt��@�o\.�vX�E��=�=	�'~h= ��
]� @.�?b�m��Rx�37��IO�L�glC�8SDe���������O�A���}��P�ɺo���"OP�%j��lHW�����"OX��W�I>oBM(�K8/f|�2"O���'�NM�$p��ϥ����"O
�jB�J��f���閮�,��$:�S�S�q��(Ô
Ś"�}��ǙrD>B�I�/�Z]����o� �	 �?&Wr�O�=�}� v�!�/?��H6!�U����W"O�Yòb�!in(Vχ�hF"�R"O�馡��o�1�U[�0���'���c�V4���*��I�rnT�#���#"O4�!ׄıiAP�h��T4wjRd���'\d#=�� �N� ���g�%��e�_�<qD�˫I=�P"���,���^[}"�)ҧ�z���F���5�]�5h��,�D&�ON�c���=��l���!���"O��U�X�D� �;M��d�"O��4$ǭ"b]3C��:�²"O(��HB�!��r�c�z��K�"OV���ʘ4/ne`��La>�Z�"ONı�c,X�P���g�J����"O�#' �
���HS'P�2�`��Q"O:�a�B5j�D�j0%H� ��ݳ@"Ol�q�e͹?}��0oU5��4�b�i:ў"~nZ�Kth\@e' �oꨱ��hB04H�C�	&b<��P��%���P7`�4��B�ɘR��-�1ڦ����  Dg�B��];V��'�I�1It��c�,B�I6tRU�o�.8���w�� )�C�	�_� �� I�15L�t f��{��C�.*��c�("<�L*�k[1XU�C�	�QA�Y����
T��C��C�AI�C�I�?����ub�n��`�B�x�~B�6Y�F4�f��.��A���E'x~B�I]�~�:7��}���է�ƲB�I2vtt��� Zpj���8B�I�/��Q�cF�&6� �
6shC�I>U����Dȑ6a�uc6(�&C�IF�4�F�K��"E��&A�
C䉶4���NZ�qx�E�e��U�C��
_���`hB�!��ԊE�^'<E�B�I�0N:}� �	*fh��,ǿ��B�I�8�� �� X30��"`��;b�C�ɥY��� ,EVD���I8X�C�	�I���j��>m@2E����(@��C�ɛw�ؤ�f	}�"�+J<m�C�	�^����JA?\D��k�e��:�fC��0Ր��EC��U�0ʛ�Z�ZC�Ɏ9}T���Y4+�*�A�1"O�iL^��R�����,�0��"O�p���`o\P�&��]u��3"O̭��c\P̌ YDƑ�^i�"O�q���1.��#����}#"O�ْƩ6��B�䊋�^:�"O^@C�)�=)��Q�N�gϊ\�"O���"+�;���[# ļ51�"O��$D�%$�l;���
��P"O�;�O\M��F�Q(�T3�"OH	z���+�lGD�B��!򤝖,�\��H���O%m��ȓ0�� ���A��Ր��͟q^��c�t���\�b=Ad�.	@���A�E; � ��f��iҗ�N��ȓ/͒d;T
ОAF	��}*T�ȓ]��D���H�C�CV8n�X��ȓq)H���J��4���cͿG��$��Hڨ0���	�����FZ�И�ȓ$�bF�Q$:�勁��[��q�ȓ7E(���'l�� {a�2&˺�����TXт�P84�E�ЮP�:��ȓ0���hgC<^�-#wa��%��e��S�? r�y�)J�$��E!!�	��* "O�9`d)7?=v@�&��Y���y�"O5�"ˉuK&�'lh|���"OP�W�>_�mxC��Re��;�"OV����VI@څ�Uk\�O��Bf"O�`�SFޝg�|���+l3D���"O���������P[��S�b���g"O�H��&Q2F�{r���9�"On]� �ξGpSH�]br9a"O����&^V�1K�aIwU���"O �Xg�B �.�s!��J@(5��"OK��z��5H� ӦiبP ���ya�;nh�Ȇ�ɯ~|��@��#�y2)	Wk0D�3E�s�j�w����y"ȝ!�\�3 Tnh<���+�yRʑ�b�z�g� 9B��E��-�y�LS.�pA��䉌�d\cU+.�y��n:d�f텀C�|�q� ��y�,��=�sB79��08Ԇ�<�y�/f9�,��ӄ6s��H�Ey�<�e�H�4뒤�qn
�|Z�8�@(�{�<q"Lb0�x��I?r���:��]u�<c���E� ��c�>ǂ,Zc��x�<����"sV�a��ݤF��5�GBx�<Q䏓�$��)�i�"/�h�0��w�<�4�3s(	�I�F�x�!H�p�<!�RVEna�i��|��U�NS�<��֚N�����4Ȉ9R�y�<ag .\�QS�_�=v���"@�<)fOJ&f{j��� �)�A�A�<q%	G��ʵ�7��PT�M�% �B�<I� �8ǲt��g�H#�Mp��FU�<� NR<9��voFP��� �a�h�<i�bm30��E�hIS���5
�C�	*bh�0ˇ ��x��U�Ýj�B�	�b��� �K�(ٔy�,�7_:C�+:�*\�)F�`-`�9R�{(�C��i����5@rXu ��ں8�C�I�J�� $��R�bGA΢�C�I2I ��NV�d��	��B�,9��C�	a���D��1-X�MP��>'��C䉱b-F�� ϖ�-��5ȇ��k�C䉸o���k�H�4�UH�%S4SB�C�	&�P��_�aC���WE��m�C�ɾhjf�K�@ނ	Xި��#��*.�C�I�k�J4i֬��ր�f�u�C�I	1��ZU�	5c���Z���'_��C�	 t��\�d��[(��Ŏ���C�	6r`�-	A��64|�ٳӯ��4�C�	?H���S�(6m��R�J�8�B�Im�U
����xqbc��+5v�B䉿d̛u�Z/K�@�x@�A��B�	�C�����A6��X��ȗy�rB䉌(��\Sb�;H���"ǖ�.��B�	�
�X����ƍl1H��@D�Fz�B�/Jڮ��Phe\^�E�Ĝd*B�	:?
.��HN9@02P�
��	,B��(L���A��g0	w��l��C�	�r5�Q��l�@���	S}B��=`�$X�5���f�(A��Z�	 B䉡c��)��0\6�$2UkZI��C�	:f"M�4@��V5�Q��NЮC�ɪM�DS��`*�T�;6�C�	�4�ba��DطG�*x�`�Qh�C�)� pkuD��8I�ykf Z�A�����"O~,�s�Z.��!�F�h�"O�a�/�Lu��+��F�KTf��D"OL��3bG\������	B,��V"O�Yh��=5�Y1�I�<�M�r"ON�󀀱Q����lL3.�V"O�!�ը���s˗%EW0�A0"ODa�� �@HȁjeL�z��9�"O�m�&,U;� ����${����"Oz��mػ#{*�r,ݐ����`"O(�ya�ωb�B 1fK�$`���"W"O�0bզƚE�:E�UE��)�H-��"Oz�V�_�S��es�yú�Q�"O�` ��kb��6�L!_�>- G"OF�t�5?z�� �b����B"O�Hk��R�����@��{�"OlYz#�̱�D�"��>�T!�"O�]�@Hڝ5���` �x�"X��"O�QR A�cl�5�I0B(�=8�"O:8�4���Ut	r�ˁN
��P "Olͺ6�'��e��g�t��V"OF5��!ۺO�������&;�"U�"OB�wiβS˨�q���|u($"ONl�SE� f�	��JÖ	�fir�"O`뇌F�s!\y%�	 k�����"O(ĳ�F�-�	�eGC*�\bP"OF	zG	��vːl�f����@	�"O*�Y]0�ʥ;Bk�f�x�"O���P��+��9ӯ�}p��R"O��qM�1,*(�gĜ[p�Q��"O�E�D��*�8A�&�'Bq��ѕ"O2�F���_�H ఏ�#8o��QW"O��`�ѣoq��#�.^/6�r9�E"O����K�Xd����FFR47"OL��E��5m��В�n��(�R�"F"O���4?:bu��m=�z��`"O �k b��" ��UmS�v��"O�36�
�>y8'�

�R��"O���F�/P�� B�!I���ˁ"OT�Pr���nj��cg�ܗB��4;�"Ot�NQ�(`Dhi�+� C�,�G"O$�b�
��_��PQb,J�H��a(5"O��+�$ծ|>��SLJ

����"O`*��u؄+	^�q��bW"O����U�E�l�K�<�@��T"OȀ�mΗ���,7m�:�"Oh��UM\���!!��8�ހ��"O2�*H��UO
��2@�2w&�""O���`e�;��a���� ~�����"O�E�3儀i�l�"���:F]�,2�"O��;�dC��q�F��3eYz��"O~a�牚�sJ�axK�;'"O*�+�폼)/p9P�`�&/��)�"O�u�r�;�����	A�G��rs"OZ��c���E���0�٠{��:�"O�h8C$T*X\xA�Ry��2�"O��p�@R�16�pك{����"ODX��OQ���b��gJ �YS"O���UbU�0(�k7h��>�A�S��F�O^�i�N�13�R�S��^7��c�'����a��雒�-(d`K�"O���O��րХ/��u
�`b�"O� ��
�<:��(�CH�^	��"O����#Tq>�)�� �0�T�w"O� $�"DEȍ"���`d�Ϲ;�$�b�"O�P�� ��]�>���#�98 ���6�IL�O�j�Z�h��J_�Ѐ�I�y�"��'yr}����Ե0%�ru�m��'st)����>#2x�b�	4ĸ�0�'�`�sM��-V*H(��%��\#�'c�-:�n���싢˗�t ���
�'.��0Oܦ(�� `R�P��`�	�'���tLѹA�|���%̐��m�ϓ�O1Z�M:T|D��1bݝB/��k�"O�BD�T͙�&_�*��Q�"O��g	�79�d�X�FաI�r�[�"O>����,��1X�fT���aBA"O̝A��5R��Kw���Q�"OP����Ud�.l�C�\�_�x���"O��g[*v�� 8�<J�6�@"O�)���
�.{B�
�H&g¼Xp�"O, ��A"XY�C�n�p�q�"Oz��B.|}���S�7�N��"O�p�B�37C��r#㝾�8��"O9BvM�89@�q���A�ĕ��"O����搇$��6a��~9�$I3D������?"0��#�T���6D�T"�����xys���� D3ړ�0|*�� �j�Y O�.-Nyˢ)@_�<d灠a�>��ъ�*��C���d�<����:��k�,@&a�|X�rÈa�<I �͇aD }�畤)��i���\�<Y�V6	�<0�HC�;^P5�5M�O�<�t���O��y���"���
5� L�<�$	[�>U�3���J|J�!r�<17$�� f\ �2�[(�̅�u�Go�`���O]x�#�Y$O�AX�O
�A���
�'�8yR$l6T�b|�ᯀ�0Y��	�'_rDcW�ݪ+?L��(Rڐ�	�'G�z4cц-�$�p�
K\61 	�'5\�cC_�w������Cʬ|I�'�|�gx#y��Ё���J�ў���S��
�Y�B��PP)���0�@G{J?��mLxVz�D��4;W��" D���çGe�ze����s���E4D��aVI��j1 ��	f�޹Q$/D���Ŗozx)bo�����0D�@� K�i�X��CٵH���� -D��S��ذXw<��s�R"6{�U�5D��㡍F�A��&�07}<Q��4|Oc��iBC�#)w���w���z,��b5D���b!¦	�
	�q/M5q�P�Q.D������9`4���y��=�K*D�� �h45_ȰZ�)=m�tSe&D�Tj��	V5"�Ha��!X`t� -#D�dA���3(��M���ʗlV����!D��� ��.5 ����!& �G�#D��4.X�]��!M8Eh��4D��2�鐿&"r����M�h��1D��#e�X�	����ݍ1*�ѹ��.D�k�������˧+� }��}��+'D�� An�Y̸�:@�D�^�xYb��%D���W�_&�ra	��D�p$�03.#D�@���S	V@�	*��C���qZǆ?D����oKB쑲@A�L�Y@�7D��2ă m�I�矅Q�v��� 6D����'̬#��"�.R�-Ƭ���>D���r$\
��-���f�)�!f;D�� 2QB�55�D4!�C	�R2"O���0�W�{5���7f.R�XU�"Op�"G=:��P�ǥ�H� ���"O��FF��u�q��ڙu�<���'!�ˈV@�R��G %����,�8�!��I<+Ö��Ƃ��c��	c��gw!�.}�aÒm
�u�D�
t!���J�`$r��D:Eo mI"��_!�̝���RUcOhU��q��	��!��ż?F@K��uT��A��R�q�!�7L���`�I@� ��t�B��>L�!��?���B���:�P�b!��'Z!F�pvnęU�cCkâU!�$�Au� ��o]�A=�jA�ܣ);!�$[wJ4��EH�U7���3+� vT!�dX�z�B�����.V�\a��@V�|k!��B�(N�D[r��wm6Uq�M)%V!��,i���wD�
��X
V)̎zF!򄝣k6@T鏀[�$���Ř��B�I>i5b	�Ҁ�'��	cd
W^B�ɐLh�B �^y'����#�%C-�C�	.;]~�0dG�ǀ�BR�F<^h�C䉇u@@eŹ]-N9�B�_���C�%Y� ���>1�g�2zpC��eג,����^�`F��yRC䉱����F"	d�B�5m)�B�I��LX���[,nB %*���}@�C��xU��իGXU91�	�D��C��%HZ�0�ě�To�Qh�"
��B�	3)Bh-�ˑ�".�l�"���EՄB�d.��[⦅ zJ5;f.U�(B��/�
�[�C wHi
V��Q�V���??��J%:��1��d�f���EA�<Yգ��Z���ZWl��8Pb�{�<Y��C���2�mǸ��)Y�/D��Q��Ň%�����(�z��5�2D��x4��bjhpQH�?Ct�t�1D�h��'�'SE��� (V*><�p�2D��!�d�&Na:�aA�;:�
,!�/��(�Sܧ%�z�@���6��Y8%� _�b5��.?��)�/-�蓇�<E>����T�"�f�!s�,X��![�\@��	� ʓ�OO �1�k�=�j܄ȓ&S���&ظf9>�%,9M^����G��p����%C�q��o�*���S��M+r��?q����hqqv�V?0P a9��5?<1sW"O@�r#M�s�h���®4V$�"O~��Z"K��@$�U'PX�S"O\<��KP-E~ � �d`���"O�%� '�PGh,��)p�ۂ"O&�����j�2g�5ROd����IڟPD���%Q��1 Ɨ�C��Hb����=Q�yrÆ+	�!u��@`�8���yb�_�?S�8W���J�|tk1��y2�ɷ$���৑5B=T�h�yҥ�	F>��C,�9�x�#_*�y�牨h�P��4�5>9^������hOj��_r<2 ��
<dt, 3��M !��47�ة����S�TY�*I6�!�D��Q3DI��g��%��-���B�!�!��n���Af$�9�j�8է>
�!�d[�g��*GÃ^��������!�˱0eRU��-Qvu�p�%��(y!��_I>����' �P%j�Eלlv!�� ⥒4ݦ5�X+����r#�I"O���h�>��K��Ŏ�2!�"O���#��6���l����8�"O� �W'YY�4uӅl���b�"OV����6bнz��\�Rn���U"ON��W��a!��/��EY*�a�"OJ���j�2U��A�^� N��k&Ozy�)	�x��]��F0v�Yà$D�p �@7!A�<[U��{RP$Y�!D����*31ȜCA�7q�p訓�!D�,:S!Fj�H2�%�;+W��+4`!D�lr��l�"	���g�b����>D�D�v�!|�: ѳF��6s2��`f'D�8�2DG�2)r���<(�AE, ��?���ɔ�K���FG�Zž�#��H�T�!�d<9h8��d'�v��}�U�x�!�d֕ݠ����7$�J����5c�!��?H��t�F��q�� "agʿ
��)�C��lP���C���k'C�d ��'䬐�!(M�b�4��U;z�nia�'��1gϚ%@8����%B��eA�'����S�z DhwD�@��<�
�'7�1��l��{/�)CR!�
br�U��'��ib��?�L@�!J�Bw �@��hOx�=a���xy����I	ވ驃 V����O`���S��'7̹+�"B���3�	ʓRX��	�'�գ�H��*lZd�uK� ����'2�� %x4�Q�5�! ��@��'�BT�u���]y"U�I�
�����"����)U.2 �\��%���^���"Oֹ��H0��9�$ս�x�¢Q�PF{��Ƀ6^��`Y���:F:��o� ��Ty��'�Z���!��g�8=S☤2%��'8�`��I���ŐV��;.�a��'��z��Ӧw��-��!:Qp�M��'��8� #�07�\�З�H�J7:9��R�)�D%U�$SV\�r�0|�x��/E��y�OX�!S���Ɖ>>�2��6A���'���'Z?MS���!�>����It�&�$D���H܋,��L���!���-$D��R��g2����'�-�*\���!D���vfH*҅hDJ��:*25s��+D���`��&8'��Qȝ0N}jPc�O\�=E�T���<b=�2��?(�����W�!��ƳS@�<:�� &� u(�"/
�!�d�}7��ѐ	Q ��t����ў܅�I��̃DM>aH�
�4.��B�I,�P��� FTix�U�G$�B�I��#ŉ�)�JA":$�C䉆5:t����1y\��d���Y��=�Ó=0u9cL�Q�>��d)ШL �)��m�
�J!���%@$Ar��U����ȓ.�̕h���e�VѠ�*˝$y�=�ȓl04����J�E_�a`�EΛj�ņȓ{������-�ͺl@�v)�ȓR��PQr�ڊ0l�X��(v����pP����-]���B���7^Q��,������RR�j��ԁn/<Єȓ\&)A�O!��s�R�q��l�ȓS����.�4q�� 4�����f J�턓L:��h� amPi�ȓ7�^Y3�g�p��d�	0���ȓO@\,8�&�4�J�� aN����	v̓X���;C�.^���"�D�i,�̄�S�? �	S���s�T�qi_6h��e�"O���4D�?Z�8�q&�o���s"O*q*1D 6�$q�8}_PE�"O8�1�/];S��m���Y%�W"O*`㡍�5���צ#�����"O\y�lZ����$�`���g"O*8QVϕ�u��q���(v�0�d"OZ�D�.�HX����cmj�"�"O�ѻ���+v�=�M�DR��)�"OPu���h�X��薢86�h�"ORR0��-+Rd�zv��_@`�"OJ�R)�"�B�H`-8�ͣu"O��`�	�3*yl��S�[=�ܸi��\F��jN�v)�̲Ǌ�<��!&
1	�'�� 1��%W��4j��6���	�'�t����ȴԂ���L��O��h�# ���ȁ�D�h �ȓN(��z֧ �Y6��HS$^P�E�ȓ\V�!i"�1\AQY!�L���i&X�Js�޿<`��P�Ff|��F{R�'�?�zU��wIa���Ęhް��l7D�X ��Q�XxL�g�A�e� p+D�x�Sb�8B�9�FA�K(D�d
�Ɍ�8Ra�"B�}�e2D���G�K�AҠf�0jh�|���1D�0�Àtä��l��F�qb�9D��hq ��.���̕�p%Δ�+3D�X��W+w۲��b վh8,y�*3D�\�dP�{�*���!�6�S��1D���Fی?0� 0�ВH�$��D�/D�`�U��(:��[1/O��P��.D����<5�� K̭#�*	��.D�, �&J:,n���7o�)�<�!p +D�D�BI�=����Hۇ�塢�=D����^X5�I`�X���dcdc<D�`2gb��<�$t�U�H� ���
6�8D�`�4�X�_^N$cPʇ�x������6D���l��Z���P�ڕ0ac3D����÷+�,�	��
A�(��2D� ��%Ix� ���\�r��Yr�+D��ā5|�,չХ�fQ|�"�-D�\	BΑ|������-Zap�.D� pb�ݓB:
-��FhX�DH(������Aa	�5x�R�j�i�=L��S�"OjUh�O��A����JCT|f��P"O6���I�D�BH�щ\�ik6t��"O���WbU2mh֕؇O�?H_���c"O��{��7mF�҄��m�u��"O�1ҢϜ(��4j�e��E/����'���2��@�B����Ȏ�&���'��	�
	]��A���9#0���'�"�#��^�5� ��,U:s,���'C�ؑ�V�_�<��&��k[�T�	�'6
C&j.II���K�4c����'m6,�� L^��Ŗ[�6x��'��T���no܄����Y�����'�0)�S��O0f�1E�� �ʓW\�Q�����(��?�,��ޔ!a3ƇyL��D���������H��Q=A�%�Խ�ܘ�ȓL��ԫ��9O�@�Ŋ�t�����Pw6}I�]�unt�#�N�g�r!�ȓ��b�B�K�P$�����FP� ��T�l5�+��R��JK�-�H<��S�? ����E�4#TZ�i��f���5"O0�:r	�U
m��GJ�t��(3�"O�A�Ǯ��l(��kf��\�q��"OP� �B	[�ޭ�@�R5;�]�"Ot�/!7��iAdT<Fɢ�"O*��5��FJ�8&d��&JL�"OV����:WК�8J r4��+�"O~���'_h�6�-r���*�y�̃@�p�Ǣ̴��{�f�y&�"���aR,�?�Y��,���yb�q~.�a�@ 7
�IȐ�A�yR&�v,�ـs�8��	�#ֵ�yr�αn��
!��7�l��� �y�[9_�ޱk k�0�rq���	�yBK-�<��rn0bd�摓�y"��'c��qI�Bz���)�Y��y���88���0x�D0#�@�y"���l�lĳ�"�1�F�A��y��9�bFaM	���Kk��y��Lfp����oreh2a��y�e�U�$(էL	�mKR/��y�G<�M[�a�� ��c�C3�y2B�V�,��+PsFz)���yr(��#e�[` O�f!x�#�*^�yb��}���3aJ�6Z�va�So���y�M��+B���	�(^n@���ƈ�y�E�%\����v'\t�Y�S�yB���Y�<� ��x����e�;�y�NFf���)�fעnbj�pe�˻�y
ʹ6�*Q
FH��z�~����6�y��,)�BDаu����m���y�L�)'�	k0��=l?�ȁ���y��=(.�!E쓳2��9�C[��y"@G�K������b������W�y�c��\09K½TD�\�#%Q�y�M�N�������6�YrS�<�y��1�t��#�f��t�.��y2HŶ����]�V�ɀנ�5�y��,%9������$=�<�(vM���y�(����@%:6��b�I��y�D�z��R�:�HB�%J��y2E� ��@P$�,b���$��.�y�JP�#���Ō۝Z��M�JV�y���hknD����d~ys7Hț�y����z�
)��V'aTh:'�	�y"��O>h�!mǭјhVAM�yR�N�1F�!�3��ݳ�'���ybC��ɱ1�$�ܐ�o�8�y��o|lD��c�;(��1{%e��y�&΢�Lu%�2�`pU�G"�yr��PK�p��	�eQ��S��y2��)&z�p/�i4�w��y"�;H� Pѧ$�Qb�]bƢ�yr�� #��X2�Ar���e☆�y��*��JF;?�3mb!��3C��;���|T��u���uK!�d( ��ID� zp)���H�J8!���.5����\�P����%U0!�DƦtA,�{�M�T���V���K�<is��KJ�{!kz<�B��C�<�W���j��C�lA;1�,�� �[�<i��K�W�ұ��N'����T�ZZ�<��O�P[^2�����ܥK���S�<�1�^BMh]��NE "��Xkk�P�<� �Z��$m3� �|�B=��"O�����1K�]Y�e��C���(�"Od9�V�](i�8ѱ�b�/}�X�@"O���!@���@�2a'T�wfu��"O��i.Y�,mZbe�
j��@��"O�u���p0�LSQ�ٓ.���"O5B��AX.�g��K�}2r"O��w+��4�2�z���y��Ls1"Ohh�����T�<¢/=7�H�a�"O�ZƠ>=��й�-V�k�r��T"Od��a�j8^�K�KކY��}��"OLt� ��l4의�t�0�8B"O��h��X��(��䏾�*��p"Oإ���bPb���jD�`�Lʁ"O(�!4A,~8Z�C�J��j��`Õ"O�z#��?��)R�'��\�@t��"Ot]*F�?m{4£���4��2u"O>tz���1~	��r]�:���I�"O�|�g ��l�R���W~�{�"OHX�څ�|��mV��W"O�1���B�*�/�	Pa��c��'�ў"~z���Y� [�W;jh:p۲�ؑ�y�E�ЯĔc�8�
�%U�yh��
����a��1�����y��[�=���P��W�n`Aae��yrg��zݘ�zp#-PHb��p�R ��?���H�,x�2f%��7�)"d#	�'�XE!�eX1�4�1�%*���'�P���.'^ ��7�d�̨�'���$�Z&fd����#m�x��'�����@�h�(��[~��'��=����/&��)�i@��B�'�­�$IϽX��i3��T!4	V���'�Ը�歎0W� �N�'vL���'70@R&�xԐ��xUJ�'�s���}�-r�)��{��uB�'�� �J
@R�x�s�+tJ�P
�'p��B����-��z��'}�]��E�(p�|Q��te��c�'("y���rh��됇A�c�D�)�'��)���"�@���dc���J��x����e�,i��lʆQ��k��y/�07sv�C���!2��#�?�y�(.3�-!)	�'�B�b�]/�yb��x�>Ypeфwq�	�O�yR��dˌ�Xb��h?�y�щ�>�y"��{~���f.�� ������������m��g݈j� �'*a~��{(v�Pf��r��ً�͒��y��ĐVnҐ�7�I�r��gױ�y� L<�1�F�o�v��`i]�y"X�)�F�:������K� ��ym���4TP(���qcNi�	�'Y��!�D
�����@�g�u��'AB��Nζ�zlIufژXȖ\��'�!�$�7q��Lbf��B��څ�[� �!�d΃B_�M+�ft�7��-�!�� [F�a�B.�,�)j��3,!�C�PL��d�/�����	+!��8�2��Wk��gMH����O!��B�v�t&	:���@��89H��2O�S���>���(yeTm��"O�T��l�p�i���hxp�_�tD{��铴D�L�ё/C-T����r�ޝ=�џ�I{�π $,�� �?�r@�"��e(yv"O|�y�&�:XְA�F^�k;0���"O�A�F��7��1ˑ�{#�T)�"O�K���1h^lE�c�3�P��"O�a ��x�x�Z�+%+<	J�"O���"���)�@�OΒF��yb��(�\��5�A�i8��@Ǯ��y��P�ޭ�D
߈v��Ƅ"�y��~�� !,��u�)+!����y"l�UiJ�JblA�pڤQ��y��<)�\HcG��n	D��F�*�y���T0D���Hi�L .!�y� A�Y�����8����D��yr��+���$�>b�2ѨVCY�y" �b�e#�_�S�P�bqK)�yb$C�k�, Kc�M�.2�#����y�`�5l�f���c��hq�gû�y�lY�V�N��6! 1go�}c!��y""Qb�T1� ��X���{��@��y"��:�B�h���E��y���9?����
z,�a��jW+��=I�yB��GV���mR�jӺ�+�����y� �@hQ�Dj��`���ȶ/��y2��[�b�℣��X>��6
�y�KB�cv�؛X�v�xŭ��y"CR�o�����Qm��J"��3�y2g.[/�����HV�0�ѥ���y"��+H\\�a)G
��Br�1��=��y�$M:��͐d�$&"��gP8�y�eK4(t�Тo�.k0����W��yb�̲%���;6�t�\u��B���y�؟y�r��� ��=%�%9�+���yR㞍D\���d
�f�|�2T��5��'�ў�OE8<
�H��Nv���U��,A���	�'z((H��T(
O���u�۶h���s	�'f��� �9�ܤU [�_R؄�t�N�K���-}�:X��n4
	"m��ZҖ]b�\9o�@�Q����!���ȓ3Ֆ�#��3���ҵ�'p�H���p�����ۇ�^r�Z��5b+�n@���8��Ո��S��3�*���nʞ܀��|"�)�10H�8r�$L�^������
e:D�O��=�}J	�qi@����6�n!��a�<���6��hdF>Yf�E���r�<)��4C�j 0��$bq�9XH�<Qr�H�d̨آBI�x��[s�@G�<Y���6�Y�A� �mv��lAx�4Dx�����Փ�)�J���*;�y�Y!�0��lM	jٞ�C��)�hO��𩙀4�	�3��p����)i�!�d]�{�P�0D��L���E�D'{�!��C느�1F<S�	����g!��2f=2�`�>"���mU3L�!�D�9�^�Ó�_	j �Y8J�)5�!�$���L��d��B�ʡ��od'�'a|R�T�?�����l /����g%���<Q��d�UT�����Z@�P��W0!��ҶRX�@	"�V�e^L�k��J6<�!�d	l��K��7EV��#���!�d�>.�3�'׿v�����Iş�?E�%I s�q�o֖H�h���Ly��'E�O#|rr�V�ri�Lk�D�a�x�9��QQ�'�?-K7�V�8�@Y�s�[�H� rs2D�Ti��4J�nA�p�1V�Ji�c/=D�� �<��q�졂�5'r�z"On0�D	nh�b&�"{.A"O�eS��L 	�(_�xhI���|��)�ӊv��)�d^2+z�Z��1�ʓ�hOQ>�(�m�J��*���l���B��Ob�=ш�	J�p�ѡ�͇�{P��bW���!�� ��ʕ�
2?f����ŕy�!��
Z{PL�e� R����D�ǋ#�!�dS`u��x�1-�4p��ȝ$c!�d@<�D�h��X�)��:��Ϧc^b�)�'u8�C��Jh�p��B�.���'��"��B�kUL!��i[c8<�
�'̶p���P)'�ڠP��T!���'K �1�Ŕ8[�	�� ƁH53�'M�I�۱h)�XuEҜ`]�q(�'��K5�S"#V�@K6[�����'�xu�� X�
�E[@�j����D8O�A�D�]�y�h�3�B&|�,̀$"Ol�2$��?"�0��rk�n�@�;�"O�Q�C�?#�Ȼ�`ș!�T���"O�:��X�F�D��r��/qE8�{ "O�YFƃt�h�Z3#].s�5V"Oʐ�c'�7!;^A��`ށC�X�c"O`��Q�&Ȃ
����&��+��'����}׶����q��1y�C�ɸv�,	�,6NL�v�R����þv` ��T�9� `�wHթ%7!�$ʭ[�Ʃ��댤<�֍0�F��'5!�$�>%̰Y�e��&|��  ���/,!�d9c��0�4F��aÉW�M�!�D�(,�8%AU��s���z����{���B��d��b�<	�H6���s���)�Y0��^����'ϙ�9=D�Q�'-���b	��Q���P�J�C�ɢ�'g&�St�PV�8-�ЎQ�j2���'�4q���{Gh��G��dK$���'4�� j[�,nlmDB��U|�-#�'��4�W*�0Ქ`�EH��E*�'t��9q�OF��3���I�����;O��Z��CR�4A�M
^Jr"O�H�̜�F��,��8�w`�
Q�!�^攑����?��`cE��?v�!���v{��qբ�	 ���Z�`�!�	�^���F�d�V���M_�f��}��'�d�8K>�1��m̑��-�ROU�=h!�]h���wK�'[�u�m�ў<��	��Q���6��eq Iv��B�IM��@�Bق	������bB� ��ph���(?�~��o�`�>B䉚cZ@m���x�dE�	%D�NC�	}5$YGn�j��#3��ON���g����AA�-�ƕ�����i��f?D�tR`���kF���Ѓ/��h�>D�H�r��}�V�c¦�)/�t�p�;D�� g�UM]�m�� �O�t��R�+D��;p�� �lI��K����rJ+D��bS�X>fv�i36,�!N�]zr�'D�()ĊI!Y�ٻB�Z*$�M��'<O�"<��gY*�N"�o��#�����J�<���ծ6|t\��fѸ45h�RB ]�<�sJ�U��-���7e�* �Er�<1�Mgx��i�ŵ[�)�K�k�<ɴ�K�j+����	.yvd�A�`�<A��Ykb���Õ/k��Z�BX�<� $
��G�_Bl�ѡ��7�Fh{�"O�=(�Bz����3@�B|�106"O�Y:��I�1��;��Ez�t"OB���-�k��M�,�I�"OQۡO^ ��`ss�@8,�"��B"O�i{��̊	b�%��n@��ޤ��"O�YƊU�w
N	�P,�ܵ�E"O�ACFLܑW���3�*��h*،��'m"�'��I?������C!Hk���w�<���ȓ}�=S7�_'~ �ElɆ,{�ȓB�y�7ǳ9F��@�?aX����|zB�e��<���G�Ȑ �~��ȓ8���:qˀ@|�E�ԍύ#���ȓT��QSv�_;�EB��[�H�.A�ȓ	y�����!�"t��:$���]�����V�7��D�7g�Ԍ�ȓ^���á��ȉ�!�3^"�(�ȓe0(h��A� �ҩ� �ڮ1� ��ȓ�VA-̜MѰ8.�<�s��k�<��E7qV��H�o��@-�e�G�k�<iJ�Ka��`��X&
80��c�<q�C��p��D�<��[�ɐb�<�4�Ԑ8P�e�5��6-���a�<��/s����'�0!�Ry* )K_�<aK���hzP�8!Ė@:�b�s�<a�O�=�h(���$J��h]q�<�B!#(i57n�D�Y�!	j�<��j�5 ���ǫ�(5~��P�p�<�3�����#a����0�l�<9�N۳w�n�2c�dv�R��K�<!!2lЉTn��K������CP�<q�%é}���3��z�ȁJv�N�<�V(߹Y�" A��Rx0!��I�<!7	G�k������V��(X�@~�<�4�X)�9	G>ϲ��rGIp�<y"됸�W�4(�$4h��p�<i��M+Ƅ��FL-iTXA�m�<����%s(� �� j�*`�sn�P�<���
tּ�����:��٨���v�<i��^ |�]��MÕ(���[҂J�<iQK;w!�i����%�t�F�H�<4�F/ာ�Lε$�B�E�<�3Cի2E&$�0��;k�@!�A�@�<�D͟	�髰��f,��3K�~�<ᇉ�TU�T���Y���#�Ld�<�O� ��`z���4�,���M�k�<���Pp����IHv�]���f�<`(T )���f���� �A�H�<AQ��	"T#�&Oplh �D�<�QH֦\x>$x '@�b����!�B�<q�OԤh�i�ŋ(R|�k'�|�<i��V��mȣ5S��� �y�<��EtH�k"E���@��eGs�<af��+�6Er&댉���q�&z�<!��o�6��2��>G�(���}�<�c�Pe $�F �:sL�0$�|�<��b�����Ra&
�r2�I�fv�<���j\�XJ� V.k_fـ�,Fn�<t*C�)�`{��-KS�EZ b;T�삵e�AN�< ��U���%L#D�����E M�l +��.">�p�l#D��S�ՉE��	�1�?v�TEӢ7D�X[t� ��0YUo�	�zX�(D��r�n��NuXx�wDF�-xʓ-$D�� ���aB"!�b��1��	o��a�e"O�联`J�`Aژ����n���k�"Ol����4���X��Ӌ@~��Ja"OJd!֡� t� ��D8nh��U"O��	�D��Bޜ� F�H�V��V"O�R(E�ij�c�o�s�H�Pb"O��seo������
N� �"OR��a�\��y�e�݂"�h�bs"O�h�˯f�t�Ε*-9��"O�K@G/:��Ս�!F��"O0��9zoX��2�
J����"O� ������� )H1iW"O^0�N:�)� Թ!	��Sc"O&X���7v��q�L�d��Q"O-����|�����1+:�zt"O���[, P\�A,C=P��8�"O�y l�'[ <��+B$ �`	��"O�-�B@Ϋqi�	3@�T(_.,ڷ"O�}�D�v��0���2\�"O:�X���:R讽�i��A�vr�"O$��P���7�L��(͍ �:���"O�M� �ߢ,��(��f�_�@�"O��ЊZ���[�&4�v}�A"O�R� �m��J3�_�n���S"O�1�g�mՎ�IE�/��pt"O�v����g7p<ҥJF ]�~�ȓgK4��!)�2y�H�c�L!Jd���ȓ)��5�O�;�R���l�X��6��e�šf�"͓�gJs�⹅�����kF�qjݰ��^#M�}�ȓ$~��w+�O(�h�)�W�(��^��9��9i�a�v���$��E�����$Z�`�aYw�����b�
�J���-!:YH�!��Qu ��D�\��O9%���A�d�؄ȓq����CG�w� )���.��ȓ
B���C$muv��p��	f�D�ȓ��9`J\��i���1�DI��PH ��.RdmA1GR.G T5��q%¨Qem�8p����#�1���%�V�
��W�%G�#���[��l��}��ˠCZ�&R�2�莓�,�ȓ'��TA�$��OmZE#4J���<��|��� �^\x�r�j��E ��ȓAWF�QDضh��ȊEf۟�$��ȓ$�`b�e�C���甚Id����<���H��K/6�0�G*ܼ8\x�ȓW�v9V'ǘR���`W������ȓF�t���}�@@�3@�ņȓ>K�H��L�pt��1N�Odp��ȓ�.�XFb����`����Z��+�" x����L�Q�w�<J�1�ȓ޴���N�j`rQb�;9�����f
T�nˢ�
�ҁ�5�h��%�	۠O\��f��A.�.$��ȓ`� ���Q=�����ԧS�� ��g��8a���*I�L�B+YT��Q��^Yh@S ����ô!�
s����>=AT��`.�$8�!&WR��ȓB��� ���4Iw:�kV@�*x�̄�	�xa���^�+�㈱Y�)��4��)���+?.lP�d$�O�,D�ȓ r�	��$w}�!�Q�u��u��(�Ұ�%S*6Y�Ayb�?@����S�? ���Ț&r��0�@�_�Lr&"Oh�B��J��τ�|u���"O�\��fC�\pZ�AsMV4Jt����"O,i���P� fX�0��նLnrM{Q"O~\�/ؔ�� �*Q� ^��#�"O���B�I�4�8"$�,hY )��"O��*B��c�T�D��IK���4"O:��C
��J���)@�\1R�B�"O�m��b�����@��f���"O� �Gh� +&��)w�O^B$X"O�;b/�&�lء���9H�,у�"O�Li��('��9Җm��/���"O���Q�՘T��kQ-��v�&"OƘ��H�x����R[K:�1�"O�-;D�2�
�j��_0Lg���"O�$�f�V6K>�p&'�BNh�)"O$D��N�ip�HA�W	f�� "O�y���~D�S�U���!��"O��D�+4X@�"�9� ��"O��%f�H�PdbW���y"j��"OT ;�N߼g��t@ꘊ\���"O l�h�X���@�d�� ��"O�pѶ Y0��臯�c.8��"On�������`G��9�`M8�"O~���"����G',�¥2�"O8��(�! ��}�Ɓ�cᆠ��"O�����t���y�V�8�F��g"Oyzc]�d4�p�����t%�f"O"��'��#'��p�LĠ,��1A"O�i�/H�@B+F���2"O�E偏:x����R�	�~��p�"O$p��J�-3� �B�͊��-�6"O ���n�+�Y�u�'O漴��"O�MÃJ�02��a�GM<�X�3u"OzX��W���Kܴ!,+��_�<�!�|�����E��D\��q�<1+	�M65�H�7m��p�T�s�<A�Gӿ{�Е�VG�v�X��gA^p�<I�*	I'��8�mӑy��Ҍo�<�p���w�z���`]
ښ{wOi�<��L�v/*��"��h��0�Rj�<TI�X`�s�=�����i�<)���TV�
���"8H�ȵ�Ig�<�!�W(e����l�\�&�HSĎf�<a�/T�Z�PA��G�aa�h�*Vd�<)5��E��- #���PED @Ī�a�<1����-��1��s�@��#�]��X�>1�C"b�lŲa㘗A����T�<��b�<OЈm���F�&�.����QHܓ�hO�O�bP�	-dNF�pt�M�#<�p��A.4�܊���(rGJP*�M.8�&%G�nӨ�=�'0��O�С�`�3 ���F��V��}#�"O*y�� Ǔ:�����"[�bxH9�BW�DlZo���O_�QCjR�vS�a�� ���	ۓ߸��$ґF즑:B��=2���f��S�<9��Ex�Y�3�:��i�F�'D�?�X�Z�[�jH�� �R|�`�N"D�\*w��d�v|����ZU��Ȣ-?D�x#&���*�Avn�..�Y�@:D�lq���K
- ���U��7�e���O��Hkk�;��!1@�6k�$Mq�'`����4n@:ի��&-L���d-<O�SF�Ӫ��J���!D<��@"ON��`@��ntqӪW3U*��"O� �0�)Sάݸ�ŋ'�5�"O��('�эk�	�'/%�3b"O�qІ�N�}����SA˗]l4j#"O򱲁D�?�ZБ'#�$]MlX���'t�b㊜')�E/EN���I�C�<�����1�py����\��E�ì�?T�O6�=�}R"(R�r���!~αAm]U�IN�P��ɟ�-F��IB@��`���R��3�Xl��Q�4bp"�CB�vB�I!s�0qr���y���k����>����ie}r��غ�<	�1���<	�JY"p:rԓ@>G��8u�e?�
�(����c탁PPS�h��v�܅ȓQ�h��]	k��2HK4%���H��l�umB�F&��:��4T����/XBQf�>Оp�BN7z�p}��7�pl��I�#ko����1{�@Ʉȓn�L�rю@ E���f� ,i�2e�ȓX���ܼw`��9�BS-]���'�͓�M��'�� ��ф4�PeYaA>|xG~��� ��o��
�1|*�j��$8�:��U�O-���<�O��zх%�xx˛�;�`��r�-�I���p�SG��	6�΂t4��tֆN��t˪<)�MS�]���#��Т�Y�`�Q���<�۴��훶��3��'|db�%U�U��|
�kX�w�J� 
�[��P
:
^���ֹw e�a��S!�xAF����e\9�e�rOQ�����8u� �S�J_�5���튣3~B��5��h�Lݢo��x	�I�e�B�I�\���Ђ�54n|��oƨ#?�B�ɲ=���'(� yMJrc=O�Ft��%C:�D�B�F ���i�a�	]�����?����4:�X��(H�zNT`�I���M�?�����Iq���`����V�"٘L1U%�[��b�"O8Pbf�ִzr佐GK�����V"O(${Sg�	:�*)�ƹ��'w���=	ߴG�\h9��v"԰�ץ��n/Ԅ{�O�8�gZ�5��#���34����>q��X t�O���i]�T�f�#�ON*�tX�"Ox�W�Q"!��0�d�� ��T�|rΔ� �ў�Oa![N� ��$��a�&]�p�	�'��5��(̯HKXe��.������$D�<h7o �:��LZ��&Q͞T���8��>��>9�'��3$�P8S�/��
1D� ��l��|� 5'�
@�݈#a4}r=O�c���~���Hq֐�m_9*ٙF'i�<� �L�iE� �VcPv�5�tJ�n�	P��Gyb�x��=��U[b ̩ ΄2�	^��y�jO=5�ԑ2�%/hH ��ȜҘ'>ўb>9����(z5��v�I8ĉ�c8ғ�hO�>I������08�9K��|�H#=�;��,Q��%�������3#w8H��[�>I���I�9��1M�ڠ��J����A�{���C�@�3ܰ��B�VȢ$dUЅ��5i8��}�<1�J�.���k�7�)���|��hO�O�����Bݏ:�@i��D�vY�)��'��b7gK/+�� '�-^�����'�b���n�eq8x��T�l(�'z�4o�e&j��E��>},�'qZ���&G#~����1���p.��
�'�������\�YA��@E5`
�'��y[���AJ(� �=5��i
�'���ʒ�J�8gԸ��nL W�Y��� ���q���Vzl���A#F��""O�52�@�>sz���ˍ4?�h8�U�>A�'�O�(����2����!	A���`��*O�(���g�` �3�J�B���Ӊ}�i*ay�hB�d�,A��Q40�:U��n���p?��Oд�K�$�z�c�<���;"O"eǎ#&��v���M�������OT7ͷ<��O�Ӎq6��Ea͞f�p`� \̲B�vK�([L$�KE�.6�%���Klܓ�hO�O�pb5%��T��͑a�R�?�%��'Xɐ��d����IA�/���M)�Ĥ�TG{*�<�b�)
D�&���ȏ:X8!0�'�Q�,J�G�k!ޑ�F�B���A�$D� �0�?�*�DA��mz�:�l"D�ġ׋��MW��U�"JLl��g?D�Ƞ0�֔2�&��2W�0�`�<D��`f�B0xM|���H�C?V���94�hy��j�Փ�KR�#0�L"3bOB��Iq?��{��)�?SKB�e�%/<�Ӷg�)��yBa�q�R��Y"��@~(<@�� �BqFx§<,ON!��"��GU�榖�20Д�A�O��I��h��Q
v��9HZ�	�טF]���j�M؞L�F��$K�ģ��ݐ�0���%}�]�%������GT�4�Cv#��ȋB�Ùl'!�dOV�t��.6���"�\86Q���I���)c"�� p�L�K1�ǈK
*B䉩K�$�i�E�R�rd ���U����'�~BN[�]���z6h��Yd�B.�p=��}r��N�P�֯�$k�y���^��y��w;d�t�� |� FDǦ�yɄ6!� 5@��A6��q��y2D��D���ܐx�B�qVk��y� �{���/Y�p����y"�9}�(���R�i��4���.�y�T>x��1�A,�a��C%b'�(O@p���ԟ&�r�f�+�
G^�w�!�1"O���S�m��LC��Z�$S%"O�����!P�� �N�3o��u7�'�@UDx�8 �!K����v%���C%�y��O�Q�n�c����r�*@�C���IN���O�L)#��4�ا�]�y���'�~Q�ƀ\�l;�	G�0��&����'�R���	�t&\��+^�q���?x>�B�ɣw�i�&ƠAطf�n�|B�ɓ$8�9�Ci�6NjU`3"�)^d���,��'���Ȇ�G5ڰ5y�kE,'��	�'~U��i��Xiƕ(e�B�$2
`�'S����ȩ�����E������'n��e��"s2���i7D�Y�'�r�
`
�	�xq�R�ʝr�Z�y�'	p��І�:��$�fCO���I�'�pd"�*�uJ�;C�Ԧ
i(��'�`x���;@j5)��Q����'��`�r	�c��uCe�̶C$�%��'bL�kU�f��X�d���l�|���'�,	B�§|��sD@!]�h���'�إ�,�	cW�m����$N��]	�'{.���<=�0Rc�Nr��'����gg��G\LB4���n<��')��9%��3�����ܹ ��4��'z�Y��	Ϲ5���\%Fu����'Ɯ��ԧ �x ��M��pJ-X�'��A�!¿Ov�������o_����'T�# 
E��D���K;nn����� ���𦑰|�T˶@�Y�Zm�g"O&5�`��.6��a ��Y��y�S"O"{dƉ�wv�X�����h��"O�mSe30Zy@.�T.`��"O�mx4ɒ�R��Zp�Ѭy>E�"O�����X�8�}YBMס|�%1"O�D+�〯\�bE:-�:.$�f"Oh��hM�y,�"�͍2��Ӑ"OX� ��3��`��$�`��"O��2�� d��h�*�����P"O��I�o
Z��!�pc���"OJ	��_�F�̕[׀��3�!"O��6W��� 
J.��p�"O T���ÜB9 yӃ��{�tI�"O�s���n.NY�G�>W���*�"O��Z"��)G٫��}���w=O4��$Q>=n�ݢ��ݹv،�"��ɧ.V�a��.@�Ҡ��/�
A�C�ɼZz~Lsv�,���TЉ,o�C��pd1�F%~�i�5�N�@;�C䉐/�e�V&1Gxr�F�N֤B�ɑS����3�2$<�y	�!E :~pB䉕e�"X�K)�v����1l�tB�I�U����D#}��� QZ�B��?tZ�ls�d2�� ��7q��B䉤g�6��X��p�mL�]�`B�ɏt?���������A��C�<X��!͗3����#�H�:��C䉂P�pP�f�+�|����Z-�ZC��6"�e;�o����2��V�/d!�J>4堶��%tf�C��1&i!򄙔�����)L��뇦�"I5!��ڳM��M�L�n+*p	+���!��T���9V�B�vfѸ��,�!�DA�SHD��T�ڂw��3�P!�!��Cxx��t㝄��d!�?�!򤃑!֮5��L��rm�Q����!�D� ���9f�
d��gA�%`!�$��}�n͓�&=w����w��B�!�d߄ �ơJ��Źc¥��BF�[���0@k�~�OBɚ@K�pB�\k���|��
�'e6E��C�R�0���n�4x�@�I��B�<➠F��'�U*@*�Q���A�P�)����'����+]Z5x��.-�X z����M/a}r�2FLl� �<R���di7��=�Q�8L���/���c++��h c�_�A��!LŪ!aH�Mz@��2�[g;h�?i��E"��
ٱ-��Ԛ0"�-0���ڕgS_�<�;d���X�ݧ#X2���2���s���+�g?٤�֊� p�f�J��~qJ���y�<���Yf ��%�U���y�O�ҟ� ��Ɠ\a}RK�<��}�6��%.�����%V��0>Ve\���´r�t�	 �qҢZ�L.��	�'Q$E��Po �C�Jl5N�h	�'�tQ���И}�,��Q#�#Yx�ܛ	�' |1�f��5Ej	!'ڞ*�r�����#j��#}b���"�F�#PB��Y�Z����HY�<�w̋�rb�b�LQ1(}jŚ2��<9wƁ�e��"~*���h�a��1+��m���[�<��H���~�#4C�C� ze`I~r��(����ɣ]Cna`����*t@Q�Q�T��N��$�f(�:r�Q>UD�1��
8��1V���|(!�D�?�<Ab�M��-�`��a��.e�d�G��KOQ>9��,�Brb�2��3{�, ��!D���pJ�8T��MU�:p#�}�0�3��03�qO?� X �ԁ��Gr\�%@64�hA��"O
|0��3,ơJp	��;�x����>Q�`�ڰ=A����b��%=�-+�J^|�<�Ё�(��H�&n� �P�K{�<ѷm�2������D3�B(pq�Lv�<A��]�wF$$�כ��u���e�<�!%	�4H�"%�/N��L\�<�t��01*l�s�Δq�����Z�<tǉ$vn<��B
�MQ>�C��N�<y�C�4t�X[fFԉj�-h�\�<�$F��O�<=9��J�N~�Ax"��C�<��@FA���˗E��K��} ��U�<����Z8¤
9D*h�V�I�D(l�'�:���e�����-��Q
ד~���sS�E�v�����O�9f/�=a���tR.l�J�s��9��Z@��[||�HFF�=��Y���"�I�<��M�� ­J���G�	eg�D�K|��e��]sK��9ؼp��E�h�B�ɧ#��Pq�&�=��	"�$K�`B��tkh4�íݡ0+XL�č ��H����  �T3sC�pt��l@�C�ɓd�`�4��6��<��"�	�$qKƍ�J)HE3��K";-t����bޢ>�w��!Ǯ|�УMb�i���mx�t �AѠKn��	'a�~opI &��9���@e��;��d�ٰC~���Q�*�)��.J$rǰm�/&�d
�qͨQkr�`�rd�� ���PGL;
�i��t
��kF�A�V��b��H�<Y��NQ���vB�>^����E*Ʉc��tp��ɾk,�ųE��]��tP��t�ר!�.��fPu�`	߁G�l��J�<J���dC'��y�f�\:X0J��1�Q�l��}Z�.\�l
ҕӕ��O)�6�_&��QF{R'\'���Ȟ���h�3/۟��'w�m��r?�5h8��X��oZ!y���e@
1;��;�(�{��"�-
�8��IA9R��}��)'�{P��	~�z�/�	Z`9�2"�z?���!X��+H���H�-��<F 1ü��׺z�=x�����i�
�Q}���2|��O�>�r�%)U�N1�𮅤��1�E+$Z��*�n���Bx�A��[��z҅��V�@)�Ў�?��rM�O\AǏ�.&k�!Sr�Եrw(��`�>Q�(�!�	�%PiS��<����b�hH5c�T,a����%�<)&N�Q9�	���H hd"ꁒ`�b�h!�� c����Q�����AY�d�IXw�� 3�<���f�~g�`	�5��;>�(' �.��aΝ�|1$�fd[&x<耨�Z�$*%��("��bU�7�O�h��F�+N�"Ѻ�cW6z���ٔ�OZe*�IW��~b�R����9���H�$�̻;���H��Y�j�ң�B>��A����$�7�)sb9�Yl�`�-���A�C^�Wh��~bdV*e��R�мG��|���INv��'C���I�=��� ��
\M�6r��' �����\]?ɓ(��Q��֝�W\����m\����q�I�î�O����#w�b-!�N�?�$��)2�D(R�K�R�D��	�t6��!0�A<0.�H�dOԂ1��9�
��!�%J�{����-ɻ���Ӌ,W>�+�P������1���>!y��w�^����(1J_S���)�KK(2�5�0���x��i��G`���2S�i��Ȥ�?OF���0�%�p��}���:�y�FV'{njF��'`/�Ya&��p?Qq&�\��-I��
�
�Sj�2S�D�{��F����I�0�� #��r���ܠ�p�8������)�to:��̋J�<a�Wd%�?�\�y��3�'L�������I(p��kѢ)qέ�h/?)«��DW�sI~�=�$��3�����[��G}� �q�O�XS��Z�q�R�@άr�؋e�Ѿ
"�ˡ�0?	!fݮ0l�!���PV�
eh8������%@Xy���t��p�;P�B	@�*%�Cf(D�PCg�)V��c�ż>�}IL;}�g��|q�)��v>	�p@�zSh�D��(ዑ�;D��B��;N�UNC
3bYbTM�#1�'d ��H�O�g�1Z��eǙG{|8Dm�4O�XB�	*�dJ�%�w�(�9A�-pd腨�`J�BP-R��'�����\O��A��$Ap��sQ0��^�Q��7upˇ�B�G�mC��� [�9�ȓJ�>�:��*V�����@T�5�(�O���AA)ym4Yç�J�PP�O�Q�ʅ
u��K�6��u0�`�S@���Z|r��N(Q��Mp'�/���(S��Y�~&�@7�ЖK[��IpH���0ѡ!4�JSnN�>8 j�!�7 ��Px!�ϼ5�������� �� l
�k\�+ �H|x
��ޘĠ��Y��L���S���g�!&`]�$'EyǢ]�HP<��_��95��"!nI���F�T��9���\5$���d8au <����9I��x���jNzeP�-ʮ4;�O�y�⋍�4}�8����>h
��]��m�֟BHy�_&@�p�c	U�Υ� "O>���W�B�k��?C�4xe,�B\Q�H�:#��Ă���S�(�9��Ġ���ug_�fGڹ��+,1��Ƭ�q�<��U�xX��*l�ł�%8�B� ��F�QNv�qf��Ud��o�	�l�<��'Ŝ7]<��A�A%}�2Y⑮{���J 	^�J�l���yv�r�+O#�4œ�&M�6;�/�.B��0�=�p>���"�\Ԉ�O��~G����F�nܓ"��]S�V>4�� Q�B�U��+�̝����͌X�Z��\K�q�e, �!�dV$�Z�ےAն^M��K5ˏ�fru!2�8/Pa��Ě<U��sf%�^�˂U�_O���s��΅�N��mP��T&)!���"H!��*W<�pӫ��;Ő� R�B�j<�R�# 0� mA I�D�O � s��9�1�r�a�Kظ)�X+���
� �[P�'��5�rL C��ϓTm�4(3�òM����)V��{��	ß(���[�=Ǽ\��x���D��mV���Q*<M�1�Z�f��Ov��F	Y1$�c>7�R1e8XL��#�3cH�izb��O-�`�H�c6c䘧�0?1O�h	
�s�L `�̈��;r�PĐ�0O��/@�Mk7���
<Dg	�F������y�����tI�
ݛ[�T�̉��y��Ѧr��m!�! m\����X7-)m:wH_j(�pfDT�u���B/ðy�v�+᫖5YtP1pƏy��Є��v��Ԁ��x�j������=�b��M��7�VMa�@+ʨ	��`Q�'Htl��H�T,��kr��{'� ÓG���2�^�PrB�Q�!0&�B�� ��T���%^4�A��@Cxz!N�e��X�@BG�x�4�sg����),?y�N6:LI�Q�
D��`�O�%}�P�1Uv�T�Z�&�y" l�wT��1�%ڽ�yR�"q<��p���4||����J7�d!�c
�E�F\�G�G�Zg�p ��aXc�t��rq�\��/�7e�hta��%j�x���st�t�E�}b $؂-���GEդY�h�wFb��U���<𬠊#�|�B�2e4O�r,��.<J�!��+�I2U#Зt��Sٞiq�l\�L�Z��UG�$y_��	>w��5�22	#�ݛB�A*��M����`��&���������S�O9(���"ފl��P�(^>��(�����(-��l ���B�Z�Y F� �D�@A�|�	�>	bǀ�!���|�<1V�!�n��#�Uܒ8�0*X�<�J�?�n�s�)}����)XRP�b�؞W��%P��EXL1PS�Ŵ*Є�q��W%��� ��b �`�L�J~\T�'� b�՛"����'��B�H
��'����F+J4>=�XZ�0'��@	�rF`�Pu�C�|�׋�>#�Ȑ�u��p� ��<)cbV"J�b?mӓ��?
�:=������T3p�0">����y�]B`G*�5i���(&'�7\����1JdB�I�o��1�%(�½�ei�*r牛.xh�m�Z��S�O�(�y��)�<����n� !�'O�a�7�J�b,�B%G�.,a�m#�O,LP%�O[R�4��Qq[B�A�b?| 2���OJ�P��	�'@<�J��Z)@��""'�F�)#�kƳA�6�*�
O�+c��cjxD��Z`�(r�vc\�!�¬�q�T�A�eI�x���Iw�F�[�"O����:iR�т��wdj}�;OJ��F�ܬ+�*�qO�"~�AƉ%y��͹����0��f�<a����Kp漒�N�)=�^qD�j��4Q&�*¨<,OdY`4�5(*j�(��_�f#�lH��'h���(�!��y�񋟪�P���8 ���t<hPoV26�D�s�U�T���~��
b��(�����E�FՆ�4�V����	� c��2z��ȓf�j�	J�r��$��Z]j<��j?J�Ɯ<u��2cj�&l�|��X9y��O�C��P���R6�ȓO

�B9/w��5� rxņȓVL��*�l��cR�y�G?����ȓl�l����&'������F��\��S�? ��z��&ᾰ@t����T�0"O���-��B����3C�$#تi�"O�hj���o�ݲ`P$nB ��"O,�r
��k�(�9 �bCp�(�"O*� F�*��]�rC� DI�XR�"O��8+%#q���'A�%L68���"O�A �,I{��}����Y#l8at"O�e`��O�G��|j�͘%��QS"O&���e#�D,�@��4��a)d"O���FM6�QB�+$�Iې"O�4{�n4
T�d�1O�'+\1�F"Ov�ˁ�ߦ]����sn�O�\p"O�T���?omN�����R�zr"O4�)B%�G���R�l�#L����"ONU��-��H5n���ƪ-\��"O�}��Iԓ
4j��ɕ���6v!�D�;f��{�b��l�
l�$ʀ*!�/#�̌2b؋P�<���ai!�$½�65�b/֑`�����C3&!��}�J5�5b,&Bȑ����-�!�Q����a0�U wf �@�H#�!�׆YU^�eD�x^�1fa!��ju¤(�˃9''�d�/�85!�d	&{d��Q�Q8;��KT+�6!�ۧs��r1�� �� C�#x$!��Z�M}�ԯ�8QU��wm[�9!�ې%�T����v�D��'��!�S�1��iyD��y߮���D�i�!�dV�_�"�34J�%(��<B��D�*H!�D��zXpIG�$9�$u(�B/3!�D�a0���bO��6&��x�!�)J#!�$�`��s&"X������R!�w�x�i�D�5��pU	>!�dNH��,��Ӕ��PҒB�5.!��.W��R���"؂(��a�/F�!�D�(�>��t���P
�%�!��N#S�F�9���*D�L�[!xS!�Y*Z�Z,yC >$D�`Q0.I!�$�Y��6�N+hf��J�<^!�D�~X�J .ܿ;B��E&HK!��ĭU4����Ⓩ>>
��%��<�!��-��Кc�3|�u�*T�d�!�اv�|t;Rώ� A�+f�Q��!��!fN�ҏC�&f��8NS�~�!�D�+�\%�R�q8�LR�,�>jӴC�	��PA�@/K+-l�'i�H��B�	�f���ʥ�{t�`��ܵv��B�ɡ<{��cWK��*K�+@!�8E�B�I�A�%�HI
��7R"B�3�f�r��m���/W�$�B䉳7�@�KB�?�a�$�d�B�ɠd�N�Жd���Nm3���-�:B�Ii�aR-t�R�!a+�"��C��)Vw�}z[�Q,��A��C��C�ɠ4������z�a��Wx�B�	�u�=(Q���6lq�cc�#\-�B�I��z�]�=_"Az�)1Ib�B��`MH%ѡ�'/�����7�tB�	A}��5�ƨ#� ��M m�BB�	r��L�q��>O��
b�޴E#^B��&.S�Y%�G@XȰe�ҿg|C�	�.��H�H��WY��Pdm�g��C�ɻ P�%���=G�fԀ��)]�bC�	/�t��#�ҝdɛ6ȍ<�.C�)� 6�	g)�f�,�Zp*W/���;D"O�����N�PYx��6ݓ0��r�"Of%@��3"�.��U�تl||+"O�\�5"�
-W��bP��/^���"O@�a���W���Jd(UR��C"O�1Q���n�\��gC�r�f�"OlЂE��Z��h�U��	�daCV"O�ؠ�ӫ]��B�Oc���"O�5�e芛G� �*Tg����j"O ����N��%�'��Q��"O�a�����t�]�U&��$�d"O�mD�#!A�����X�|�B�q"OҜ�Ĭޘ ����So��8�\:�"O<��l�KӚ�*��Ϣw��њW"O�B�i[�hl����˞)*?�iQ�"O\ݣ@$ܭI�9Q��~�A�"O����H7c��͂p�מ+aq��"O��Q,�v�Hا$��k�:I"�'�!��ڢOD��I�����/=G,X�׃�#8�C�I7��X����
�9
!�	�Q_Vc�<aAI;SZ\Q#.-�^5f���-�L�M�fBN�!	@���bS���ό&Z��Aƀ���F�0[��`��O$$M6�3}��*G\�Ј�lS�OtH�����x�hp�-�U��
pj�̪tHyY��p��X X��0�*|O,�FhF�)oVy���i|(`��'m\e�uk�op0H�G��O���'��Q��i�	���>�Q7"O���D�ӣ~jF�jU	��y���C��|r�I�|���#S��K!:�}�&V�Y���1��ԨH0"�Y%l�i�<V���5��gT�G�tEYC���g9 1�0�"��d��I.�?�'��i�$#��=r\��O���2�'�08��ǭ.6<�t�1@,�9§���h�C�8C2����_.92��4RLآ��ʱxe�OpU)6�-�~"��5QB��SkK3{`�d�)��dcq�ׅwi�4)�hD+-�!�$G�[ ��� Q�H��Jf��Ppz �U�̝�~�NP�2����3�@l�T?���wy�1G�\W4`�����r��'�$L96��?{G&စ�V+����b�1OT	�oBaմ��Ē���'��ZU��r����v̔��L��ד��=c��*a�牛$k��"d�` R��Ŭ��Y��-G\�P�b\�.��7iJ�|)��L�S*�	2���qO ��gȇ k��]C�'/D���HM~�*-5���o��	��`ݎ�yb��4��ZV��)F	�e8f�@.[��=(Ӂˬ�~r�0nf��=ͧ�b�]�D@
Q�!VW�0��I12٬B�	IAF@��m�dH�І��[���%��/H@"BB�koL ��dNl|H���OA�D�N|؃�(.��z������ G
K�<y����Wz�7N�_��@hU��W8PP9��ƻu�0��%ɈD�����
�cD�Q!"�?J�r�� ��$� %q �!EU���9�49�O�Tk��;*�c��ތ\��|�1"O�h
VeC�Y�f٪`��."Y��Q$��'bP>��-O�l)'�QM��|Z3�����cT�d�A�%d�I&`�Y$"O(�g\�L˒��3D	9;8����B  |�$�� �T��?�	7nS�e��g?Y��î��Qr��b��t���y�<�ԇJC��J�ݺ7��u��;O��O�}���z�g�ɾ*$���CޣO�9��E�'��C�	Jt�P4j�0a:\� ��:��p�׉F����'^��S��Ą,�2tuw?5�Ǔ���pE�pv��,��JR��ꥯ��l��܅ȓEex��˪|��!�"�ڨi4ħO��{�œ�W�$|�ç0�x0��R�g6<����˱I|�чȓ,3��(��3o�n@R��.&�͛B��M�d�"VTT���L>�`��y�x��R��"	Vj<�!��x(<!1�ο��ma�e�
4���Q�/k���kZ�U^��$]=.�z�Cŉ��UZz��eč*S��x���&�BA��
Q~��?�7A�?|2^R�j�!��:�D���ӑZ$<��N�9��#�B``nI|qx��� �PR�D�(x�2�¦�˗"O���釧^#��(�/�O)�(���H��O+�<����x�.�zhXk���u������؋��xr ʶ"�����eU�?�ZAP�
�>"�d;2+	O؟tҳ��kx��H���-�g≷;�����H�3�ɪ�"5������y�Gϻ0���z�� +�(uB��<xP��'��#��I+dE#�����<g��yCn��l9�P�V��<��>�u+�����ْ�̻HRH�E��Y�S.$}�ux�
�V�|�p	-��B�I��,��.��P7J�H4��$���HH�9Ꜥs��A��b��.�'��D�?/����:`� �8���� �'�ڤ�7H(u�4�R�E]�~�R�"��M�}� ��S�FU���Ʉ/W��"?Y��S�Sئ]3!��e�x�S�e����w!X/�ֈ���-K#^���M	�[�>$�c���"��e@ ��9ٞ���I2[v��D�{HT��5��^ ��2��H,8������#���{��,��k�p�ɷ-Խ8�aA���!�d�8=����s�IK�)c�kB�,#���Sʈ�?��8����7�&�Bb�8<����c��J�-�s���
)]r"�*7`��,���
��& !�D�d�N!K����U�`F"�!a6��1��n�!H��X��O^	@����1���z�GQi�6u �D H��l��'�!as��)&^B�ϓ'�(��c@29mi�VFéhu\�K"�� ���P7jb8��&'�x���$A�^�db�`�,��!ۄ�
?)߱O4)��xc>7M��jԲ``DZGfu�!� %Q��+����6R���V�0?�C!���8fY� /6� �_�>6��1O���"��M�g�V�.���L�Px��'�y��K�?ϊ̪WL�
@2���<�y�A�v-UbG�ۣ��(��E���{�b�'p��°�˱I�\ˏ�4٧B)����䜚G�^84R�ɧ�&�����b�V�~��!Gk���ѩ��.n���)O�p��(q/М"D��A�N�'&���'��Eީ�I�<@|���0�l�P��L�
�!���d��Q�-�%{3!�=0���A钲������r����H9Q�v3Sq�@yTJ+?1r�>`��P����YY�W�!���S6j�W��N�(f�8�
p?�<HuK�8�y��Q̊�pAA�i9��B��64�@�숌���Cήs�BU����/q�FQ��\0���@��<R:\�c�4�(����]5�ܚ7��~�.��1��q&���X�~^�7�r�Dp��bN$�2���+����aҶw���R�UH�ቐ���[��VH����l�+O�H�A�d�?F�8!��I'%9,�ɐ����b���<F���mˣ���.�m���5/��S�O��$�U� +Y6U���H)gu�����2ZJ��E3�f��h ���6Kk�6ȵm�.A��>�w��n�}�|�=aAM��q�0�a��M�5-��37bm��
��S�u?��HÒ>E���E4)D\S%�KUVL�1c�0δ �4T����	1J>��+и&���N*���p�@�I"i�?P�J�
��W"Β�ē9Zİah�b�R����J�R,��ɥJ.��b�N�剱P�@�����6$�4P��#�kS3#�qO�����ϖ�k�^)B�)�<e ��a�	Q����m�G�q�T\[���>o�(5�#�3!��DxG"O��ɂA�c�L�Jh��6_BaR1O�u �M���yK�"~ꑡ��������"c�!��YG�<����= EV�h�ɋ	_\6,�3(�t~�S��\P��|8�D�M3t�X�Ѩ �_���9�O��b#�ók�\��u���kd��/_��S+�$�Pxra�	Wb�q4��	r	j#�ē��O*� a
�0'�j�2���JQ�>I�d�K3toX��dV.�y"�X+u��aC_�\� ���N��yB��1�I�E�@@���*�`!���6+Z}�p(�.*H4C�	:m~�
��5(���$!�3y,�'Q���Bf/ay����a�'C�v3�I{�덹ư?9�h�058���7�R�CTL֕4�@T*W�#4�88&
ٳ_��h��<�4G/D���5�O0������C��P��*D������~��a��EK�|j�����)D� hu�Hz�\�1ǟ���1#qH%D�H�!	'V|�TE[�d�D�g D�� ��Q����9�A/L�;�"Oȹ�T@V�ei�P� )�-�2\ �"O\�8�+E�f��WΛ�aKEP"O�`H�g֓*)��L]3�.���"O�Az�i�%�8x��K��k����"O�T
�׺>`n�r*D"� ���"O��9�,�>t˖�2��Qsl@9v"OtslR4���P	0@`�]��"O�1����+�h�"1'�4�r���"OĽ�B��:)��@c��.x}L�	�"O�\���&H\����֕ZS��ib"OhUH0n?o�pM�5E6ld� "O �@�+�!%��(�k7'E֩�V"O"�A��
<UBHcJO��Q7"O�E��-�z�.���I;4"\%9�"O��E��.U�8�)҉ؑZ<Z�`1"O��hIZ�za�לj
�qp�"O m��厾5�, èJ?Q��p�"O�S�)Z�4V�5CT�J7�@��V"Ob1R��.Ş��p��V��Be"O>U˲��	E��]:���AǨ��b"O�Z�Βi[�=��C�Iˆ�:�"O�Dh��A� ���V��P�S"OB�&��'=o���E�h��9Ov@�f_?_D((0�@�~�\,���	�h����>w�� %R�)s.B�		$��^ԲP��$�HA�B�ɪb~j��$�#v��MM�w*�B䉪-M�dh��\�	�x���$v�C�	6+h�a��4k�P"�/+5�C�ɉHO�!*�l�=�r�q"�,}��C�,'s����H_F�Qc�R�t�rC�ɾ`��2��B�z��w퓬��~���>%��)����!�̦Tct�!"JZ5��*]���hJ%f׽#�%������L���;�B|Aք+��)!g�$+�<�+	��dLĸ�)ؒrpa�$+�r��%�T�K�%���3�gA2C�%"�"M��PB˙�Cz ;çO�����$v�,�0Vɐ���Ԩȑ}qnIjwc���!�Q[>M!�hȨB���f9���$��"����1\�am$<�3��QM ��?qH~�hN�|:d�q�^�9dj�ZQÛ ��0������S�.�2���ӱa�Mµ��,�i[�哽q���4I�Ԕ��գm*�x�'�Z>���nC�����.����J0*��d�&DO�Z��Bi�����	��E2 �r���|x��*W�K�i�R4#R���$9_�(@˟�6-/�S�#��X�D�}8&��'a_X�1r�
EIv�ؗCB~�Q�  ��U��c�2j���рһ$V^� �x9�	��!��BF��ʉ���q�<�%×0��գ��(`��	/`ལW	G�Q����)�h}���	\�J�F��!��Q��y")R-mD�aT�->@r�����=��y�&
}�� 4#�\�H��֘�y2M�5N
�) R�N)"��d��
�y�ꂽqg�]���X2)�p@����;�y��U�\l��TC#�.E��d��yb�MC��BJI�h�.�;��%�yrLF�H�Ā81`�5��D#�	�y�d�k�T��E�'�Ȩ5�C��y���.���K��dq,�)cF@�ȓ|S� ���<*6%�r���]��a`���8�$�(��	uDĆ�O�(����%F�LE��'6_�^Ȅȓ�J!��"#}Q��BC�i��1�ȓS���W�8�F���O�Q��U��V�$!�7P� �P ���>La���b����(-��sda�6�u��<����� �,�P�덖{�BL�ȓ5P��:"^�И5�ƣ�!�����.{n�l�@"�;T�˵C�����S�? ʍ��e�3w����7��Kt� �"O +�bX�aS�T��mݿmOd�E"O��÷&C��h!`mT�~�&��"O��1��I�0eb����V�k�"O)	''�<=�Lj��@4}Riڄ"O�d�"�:R`B�����q 5�U"O�X���K���GX��2�"OCo�(�V$	�Dւ7V�T2�"O�e��+K$*P�A)�dJf"O<D��j�j(j��8I����"O ����++�8�qQAK�z�i�"Op���S4�� �(Q�v͒U"O�)����ʦ�3%��d݃w"O�)ڶK 9�a@P�N�J��6"O�]Ju΂��x���@��7��TX�"O��`��] a��� ��{��<�w"O�@�&�~�"!�t��|�����"ON�Q �g��˷��k'V(�"O8�i1��3�t�-^�z�D<�w"O�A��ʛ;M��d��1���D"OD����7��(�'��)4UB���"O4��K�;#ț�M��o��9:4a;D���%[�<i�mU0�c;D���
{���A�w�
1QsC9D�����ՙ.  �[�'߻%Y����7D��G�ܙ�@��3���t���#��2D�����\�ka�IQ'i�*ef����/D�I!l�K�(�1����=0~10� D�`0q�˩"�xUT��:_�N�S�?D��+���$m�s!�J1Ne0U!TN=D�h�d�۞(������/F�B�� �8D��)qNA/0ה�%�B�9Rը(D��
G� T91�n�0b�Ea$�(D�DR�FG�y*��r��]EbAJ��1D�dH��˽v6M�Gi�&4�2��.D�\��-D-B��5[��M�Z�MQw(0D�`��B�qۊ��c��f�Ҝ���/D���Um��	K ���P~��v�:D���HJ�f+�u��e¶
]�A�&9D�T�Q��*{ǐ\0$����a�1-6D����1_���S�����=ˁj3D��ʧC��n�98C�uz~uE2D�hR�%K��]a�
PF9�P&,D�T˧�² �p����:$ur�*+D��)t�d�ʱ�"��-�8�ǀ+D��q���Ҁ�K�Gԍ0�0�V�*D�,:�b�M��tq'#��$��q �n*D�Աj�t-���W��6^�!���'D�,En�2��`
lۢE+��%D��x��V�E�0I�mڕ[ے]h�+#D��
朳0J`�� UIb)�#D������(�K�.m Ԋ�!���:*�Թ��\'`�qq.Q�J(!�d	,x�T��@�MoPZ!k�;�!�����SQEJ-f>M���=~�!����`�$�3p�p!Q����!�Z��y2-S?S�R��� kX!�N�t�Q(֥�p��Ks�^d!��	�����'Ͷ<x���4�!��/m��bQ��#���WJ�!��UFl�{�D�/w�0c`�ZT!��޻VCݓ��I>�2=J���z!��%��M�q#�U�~p��Z�P�!���i�d ��fR6r;&PH�5�!�� f�FK�\m@Ѫb��7?�)�6"O*���-:dlU�F �C�$�Q"Op��sE�<��!+��H�E.= q"O0���Sc�	�AG�5x�I2�"O���т�(8:H�4��%G��<!&"O<(Д���X8����A�=>�)�"O�%�W�ܭ|�Xy 0K�?mج}��"O�a[��	p�]�W(�6a�&��"Oh����o��I�`爲e���
�'�4)�a`�%	z`�q�hP�'y��K@(ɋ	�J܊�',�8rPh=r���p�-4hl��'�����@�Y]���GD�9	���'�=���
?��"0&���A+�'n�!c'F�y���C���\�	�'n<�$�B#EgNXj�"O�~`�9	�'���p�9Q���1�R�u�|܈�')Ū���?b��=�pɊ�$耕�
�'�Jdct�J�C✘r�E\?$Rh8
�'b��' ��v��g�K,2e��`�'�y��EK�8�⨱� �>$pB�Y�'�"�� �:|�%�3����:5��'wd5�1���*�d�0�<͓
�'P*M�s�FE\�MK��/wZ�  �'k0	�u��$E��S�b�!n�.qz�'��Y�s�L��]ir끣����
�'�zp��/^y��U����5��N��yb,ɕer*�8p���7�ŋpaQ��yr`��XŐ5�Q#<@Ѧ���ybIɠ?�ʕ�r+����A[�ko�<��!ć,Xn�;5!���gL�J�<CG�<��*H����h��A�<�p�ɇv}�؋����8�WDe�<�2쇛Ip\zE拒��G�c�<�tj��d���*V��%c����k�]�<q5O�-̖"��<����Z�<ٲ��Wє�{p㍓FZ4�2.�q�<��N�����B!Ì]p�T��s�<qf	�'o/��0��L}`����u�<!���>	~M0DȎ�H�H$;�Dk�<ѓ�G���o�4c0��qf�<v�H�V9+ N�3U�-	t��j�<�s�R�j�`$�� �qRhZ�kDi�<Q"�S�Qе�B�SI�*���b�<��-P�`��C�N�[��i�y�<��OA':��L8񯂡xcBe�t�Nn�<�k�*u"��j��z�фnLk�<A�J�4���jf��9
l	Hv�e�<�q �.K� !��F=1�\��0�^b�<�s�m�D|�@P�S���*�_�<��R<t���i׉�6���'G�]�<Q�IG�H���/Y8�]���c�<)��YsD6d�4�\�*X"�
�Y�<9�"�	]��l�aA��7�:MJ��ZR�<�$�2�tT��)t��9Ь�P�<	fR�14T83t����Y���Bh�<!��ϡ5JX �O�0�8WI
c�<�q�X\�Q���L7J�!S�`z�<�6���3�\Aj�-�y�<a���&\�r@�W��P�"��$r�<!d�9~|��Ř< �e��dg�<��e�00��Z��^���E�g�<�b�q�BP*��O
A��4����a�<�$��!Ca�\�Ƅ;��q���E�<� ���cO�q\)8B�ʺw�|��"O֕�W!�XU�����<h{@�(U"OB�v
�/=���GJnfHm�A"O�����S�D(I򨛾?|�X�"O�Y"�,�P�⇂"LK���"O���-�M~�={�'K}�|�"O�,q�eΆB�����?� a�"O��hK�"9�,�j�opDT��38��ϰ �
�a�H>>����ȓ-��8{�@ P���H
�C��0��p�PtJ��X�M���[��
��ȓd(<�����!	�U�W�1}/ⵆ��8HzC�1�r�sOX�VA�x�ȓjʎ]�6�Χ��˴��+YvM�ȓc(F����"�����j_(n"P���zF`�٘"QN�:�b��Klm��ooF$se�m���U���b�ȓXtԩ��B�|���1R'�'O�D�ȓf��I+��#!�x8� �W�p��bV�<x��J4N�d�ɚr��`��a�E���F?�f�@V��s~|�ȓy����E��d�H���d�0�	�ȓS�ؼ���@�+�r���ݡga���ȓsf�7�M��M��(3u(��'բ���"�]�6P9�M�)�T�b�'���@,L]�![ �T0L?�,y
�'5��c�gT�~1���ԯ�r�l�	�'�H��$�(�:,��AR�n�*�S�'�J���Y��X����([
�'v\�I�R*|!qJ! �#��5p	�'�X}�vk�!4��u$�g��	�'�	!�T�cTf��Ŋ4!?��Y�'�J*�IʗJ��ɂ%����J��'�nxC�C�ht4<y0厶#�`�2�'�x�����w�JE�G,J��x�
�'�B���ҿP0��դ[�<'L��	�'�a� ��#^4���Q�֕4%ܭ��'��m�/V�D��ѡO�0|�9�'�`�)re5Oa�$�RK�(r#�'�`�C` YR�B�r��8�Ƅ{	�'s�-�.� I��3у�.d��{�'1`�e�Ǐ/k`��@ɔ�(Y���'����ҁ�X:ՠ�!'�~�k�'���FDʖ�Q���.f�k�'�Nxs�N*&��1� �?!;��'�0{�'=^V�5p�ꇮDb���'V،ـMթ2�����R=+Y��	�'���"Q���zXT�{���=.��0�	�'x&(�s�ڟ_8l9��ϰy�����'�*r$"�u����)�8��'����n	�i�p ��(&�]�'�Y�gjL $��%� '����'�b���^���1'քP\�h�'����  ���   �  Y  �  �  �)  M5  �@  �K  �V  8b  �m  
w  �~  �  H�  ��  �  '�  k�  ��  +�  ӻ  L�  ��  ��  9�  |�  ��  �  C�  ��  ��  ) � + l �  �) k1 �8  ? ?E +J  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���CO|EK�T�!�UjA�Q��Y�	'D�X����(�ت�H�H����g!|O�b�c�e]T���`�lY��!
��y"�ݔd�R®ɜQq�d���ɡ�y£-gnm8Vʙ	P,���U�W.�y��^�Vlh�'���U�F0U ȼ�y��-���h�bU�vI�����y�Q�lI�Vi	{*��Ӯ�8�y�,>%I#�gU�����A?�y�uDQ)��F�J_
b���<�y�'N�9��� D�ni(�+w$��yB��22��,���H(0x��s�]��y�� 	�1B�\u���Ò�yr�6(�4���\@�*a�W:߰?a�'�j�'ѱle&�S)A%
��Y�O�Ԅ�	�`��9Q�K�i���Q4!-7fB��  \6�i��@�L��,��Y�b��B�	�/)|G��:Wа��f	��B��.Bf=���ȂS�(H�g�/�B�	�Q��1j%��2Z��+"f��i��B�I?,�T�: 	Ҋ?/p܂�ON�"mrB��)�đ�N�6�ZAO�_e�C�I�k6���o��{���J}zC��'CGQ�F����T�V$ț�B�I� �X1�&i�FJ�����A(.�4� !���~J�D��]�!z� ��&|rwjN�<Aa��-6��%r�)�[�n��C�G���0=	�,]�ћa`��e~��.@�<qЀ �:�Q��W8�H�9t�B�	��a��g�O�Nز$���B�I#����`�O���H�f��pC�^0��6��? ^������.�ZC�|(n�kB�
=O�B���l�L{8C䉖;��A�6�]>� �uB�(�L�=�.�f�$��,N�tЃ��[0@W��ȓ02(0��h� ��g�I�IF���+]�T�Ge*`
$X���ҀL�޽���^İa�_�S�q���0\����� �1���I>��� "űq�D�=!��)��̤r���9�֖��Q�vJI�Q�!�Ƭ@�͑t�>�ʔ����Vў���)� ���p���ҷ�C�<:<2a"O��xC햭w���@��;��tr "O $��*E�gD|���-
<���)�"O�@��/ư!�"��6�߰A}�11c"O���ǋ�.�n�������{�"O�u��ΎA��@c��&q��H�"O�\���]�J����;=�  c�"O�!!_1	�yB�ŭp�bcV"O�͐��؋�ܪ�i��>R�h�"O����6f�]2��- ���"�"O�e�V �T+��C�֗�Z��"Oe(� [�I�.��5��D�>	�"O�}2��J`�؉%(��$ߞ0
P"O�!bT�Wi��ӳ���1 Mk�"O�S�M�T�RY*�[~���q�"O0]�
5%4�৮���\�2"OPi�J!lUBgN�9���г"O�P�'Wi�<՚��U�(l�P"OPhy������P��`���e"O�c�쌋S��c���~}���b"O�Y�a��W�!�CE�=	&Q��"O��Ki�1UX=ڃ�Q	| A�"O<�*��	g�vm�FC�m��u�7"O�p�4���-U�v��v�xs"O�D0�#V'��=H�cOV؈Bt"OV�ȴ�Y�k�Y�V�<]�0�U"O: ���^8 ���8'g�5V�c"O�)2U�u��`#�f�;&��U"O� �^�pYRl*��,{ʍ�U"OX+�bޡ�V��6�^�zw��j%"O��QCf���ka�0v"O��1�V�䃤�ߚ>���z$"O�I��v#Bx�j�<v䠖"O���6"��^����օ1�N���"O,�:�V��^�����a����"O��A�d/#W�� ����':�Ȇ"O����L0pZr����$��8�!"O�sE��0�01�ׁI�,X:���"Ot�Ib�>�X�a�@�\U���7"O� ;�H��Gp ��%��}�~;"OҼQ��&!o�(����/d �p0"O�A��L˕:������G�
�	�'�Z|ZMNˌ�AҤ{����	�'sZ�˱LOK).|�`�v	z���'�8ٳ��
��x�eʱnئ0r�'Ap�D�K<Y^����ŝa�`���'Z�}0өٮ�`(�E��-�	p
�'yt��T`_�>^*��DC@�N@	�'��tГ/Ҵ�,�C$ˆ!U����'P,��BIC�$"C��N��m�'�"4���/^���Ȃj}T�5��'�]����.°�K2��2u,�z�'��1�d���f�a�c��#U �c�'�e�s�+&�J�����f�`�'�
	�p�T�qb������2b��|b�'I|��a�У\�hA+!�&/�Z��' �hJ���i�!��,R�z[�'�fb�.3)HL@�ǂ�V]����'f����*����+ŐW�$���'˂�� �՗\f��
W$E�nF%1�'�TЗJ���Xq faP�M�(���'͆����pID�[�F��I���Q�'�v��[+4��yPE�@o,xK�'��0�kL�T.�(�M�`��u��� ����ӧj�P̉��1Y����V"O�`�����lN0�z�ϟ�Z�m�"O<:AY<Sn8����A�ua�"O�$c�VF����lكX'TX
�"O@dT�b�JT1��@	����'$�'��'��'���'��'*�d�V�L�Tn�p�]�V<[�'�2�'���'���'xR�'���'�^8�3�92�l�2��3D��͘��'?��'���'���'wR�'���'1�p�F̄1j� ��/(����u�'~"�'���'���'9r�'���'pp��A%��t裲�C�U�8�u�'+��'�b�'���'���'_��'%J��!���l��	Y���;���Z3�'�R�'3��'D��'���'���'�U�#�z7�Bt��؇�']��'(��'o�'�b�'�r�'	2�
�BA ��Q�+S��Ay��'�'�R�'�r�'mb�'�b�'L��`U�)-T���c�חlAЕ�U�'���'�B�'��'��'K��'�j�� ��~V����-���W�'O��'���'��'@��''��'A��8ң�9?��sg
�FH	��'��'�"�'r�'��'��'мjao�3i̜���T�-���R�'���'��'r��'��'��'県�`J�K�80���C�|��90�'���'���'t��'<b�cӐ�D�O6� ���B$����ׂ;"9���Iy�'
�)�3?���i�)	#�J2r��Hƈ@G*��2F��
����æ��?��<��sڄ:'��W��Ǐ�$SE�t2��?���Ŧ�M��O��S���K?��銾�hJ�ʔ�yH� T$3������'��>���qݮ���\T.UYbc1�M���u̓��O��6=���͍[4��j���cD�?i��yr^�b>�	Ѧ��h���X1@�(bY���C	A&/�&�̓�y��Od���4���� ykx4�2�B�h��M3C�Z�]��<N>Y�iT���y���#Z`J�C��R_��C�HL,\�O���' B�'J�d�>I7n���E2V	_"Q��y�Si�Z~��'�ba)C����O�`e��!��b�|�����n����(b�Y�,��{yr�������D�<�����V���Q�P�j%�$�����??շi��O�\.T��U"rϛ|�+�=#�$�Op�d�O~"��y�Z���T��R
���$���i1߹B�<xz�$T����4��D�O���O����r�m�@��.-״A���`I�ʓD��&�T�H�2�'�r���'ݸ5����&T�6��%��*1Έ���>)��?�I>�|�RF��I�j|�W�B�{�Zq�)ܹH`|,�~��'? �: I͟԰��|RP�D�փ�6h�c!G��8M���c��ß�����D�	���SPyr�k�X0��B�O@8��eJ�_�M�p	]?6���f/�O	nb�,��	⟰�Iʟ�jQbB�Y�����������P*\=��n�W~âp�X�D���w,��B�4$*�Y��bM|Bt�'���'��'r�'�}�D��߂l�񭝆A� ���O����O��l�B��'� 6m;�䄢Q� LZ�$�-s��ۍ�^�O����O�Η��7-=?1��Ҵs2����<7��A(���vLmk7C�O��{K>A/O���O��D�O���'ð]c�%(���S�,�a&�O���<�r�i�>4���'��'j���:9H�՘=1<HC�	 ���Yp�	���B�)r�ن>L`pk��J����6O0m���Ē���d"�ȟ,0@�|�+-�С�SH��ʈA|�2�'�"�'���D_�0��4CN�G �&zo4�[��π���$�.�?��+��ĐF}"�'�ιpSn�
A�	��&Ê�nQ(��'�"I� @�f���]
U��S���	�h?��:��!_�!c��9���oyB�'���'�b�'`�\>J�:=��~��a��d�L��aشN����?����䧉?�7��y�̊�(��b�z)�`�C��8jb�'Tɧ�O�r�!�iX�dԋ5��HYE Ң9E|	�B�	oZ�D��x %��*d
�O��?��e����r��2$q�x@�nĉ!�P͈���?���?�+O��nڃDU>��Iޟ���=e,���� WN��C��0�*��?�pQ���	���'��2��߉ld�X�#�</D�m�bH0?���C}�[۴՘O�0���?��$"9&5��I�>YDa��F��?i��?����?�����O�ql^�
�
yHU͐�Z'2\i���O��oZ�=��	�	ƟtAܴ���yׂ^<G��l�v*Z*f�����J�yr�''�.y�<ql�i~����{�0��=G��Ĳ�o˴2�����	�tF�X�c�|�Y���I����I�	���*�Y�����H���EV�Ky��w�bAx�l�OP���Ox����|�NMx�!'6/��[�kL�@f���'��'gɧ�O���2��C'�Mj&H�8v�	u�Ѕ0x>L9�O��*B!�?�rF0�d�<�
�m�*�d�]z ,҃h��?���?y���?ͧ��$�զ�q�`����ƙ�w62L �k�@T�D����"�4��'Q���?�)O�y!VO��u�N��_n����Je�ܴ����6\�q	�'{R������ ��(t��U�P�bj����['1O���O����O��D�O�?�!�/P"gd.ԉ���� �t+�^y��'6^<v��	�OJ�lD�Ʉo����j��N-�skߦ;�E$�,�����*��<l�c~"�8�dL�cI�Onl!��CYbA!�j�E?9I>Y-OL���O����O:��F�S�]��)1���ָt��O��$�<Q��iז5*�\�l��u���+z���5��~�!PFb�/��d@k}B�']�|ʟ�TQ��.@*��! �[�=HC�NMB�V�3�i>��!�' f $��1e�Y�^���!�) A藠�ҟ������i�l:��IyrDq�F࢒�:$4��;T���Bd0V`��X�͛V��q}��'��,xrŅSxvt��.W�(Y4h��'��"�ߛ����Bq�X���~R�I(e�r$q Ş�m�
���,��<I.O��D�O��D�On�$�O �'UV�i��	J���c%j�-���iL\�Y�d��B�'���w��L��Vm�I� �݇C
d���'N�|��$�B4R=�7O� ��$�'��t;� �Kܗ�y�Nhv����f��'w�I�\�ɣq��4P �A{14h���UyHr��Iҟ��ן �'L6m�%5��$�OR���Y;d�(�O�08)�$+�-À�t��Od�D�O��Ovu8�n,��<��a�KA�������yP�"3��oZ���'En���H$,vK�e��v�h�EI�џ|�	�l�I͟`D��'�di��&�/�4k�\h�'x7�M+=��˓ ���4鶴��Hŷu�NY8�GT)u+��=O����OT�D��_��7�4?YU�ۊ/6
�i�#r�i�4���Ԥa�D�/�H>I-O���O���O����O���0G�ԉscC[$7�D�r�<��iL�(��'X��'���y"fΰun�Jw���D`�w�M��꓃?����Şn�M"w
2[��aVI[�'"�BТ�:o���'M�����w�|�Q��!���&�h��ƔMh����ٟ���� �	ǟ�Uy��v�� �g��O��ꅂ��D��S�H&��)�<OPlZH�l�������� �5��
�q���v�(�Ǖ4�@El�i~R�
W�`Y�So�'ƿ�W��<V�����A4�,ġ�<i���?��?i���?Y��4Aj�b�Ю�a.����+%��'��e�p�h��?�0�4��1�p�#Fŀ�q2�t���+|�XK>���?ͧ4}���4��D�6��af�,<��I���58c���~��|r_�������쟜����qj��,9��i`�C���	`y$dӲ���*�O���O��'wg$��%��#P��c�X�Tj4�'p ��?q����S�D
QtXC��+���cl4}� ��:�旟�S:��D<��D�z�1�HVq|,3�S%�����O����O��	�<�бi�r��^8ܑN��x�=�_�9�� 럄�	��M��BǾ>q��zt0��i�b�P
<�"(����?A�뉋�M��OԄ#�ۺ��J?њ$A�`��i+��$su���Gu� �'��'�r�'�B�'d�S�W�ҥ/��#q/� V8�ܴ|�B�I�ª�?q��J�'�?1��?ͻK	XawEl�v�b�㐂A!�x����?�N>ͧ�?��%VL�ش�yB�I�[���S��-J���hF?�y�@ۻ<�8�������D�O����x�>��\�}��HӤ��>vvn�D�O���O��rC�&+F4b�'��� ��mJė,;�HM�` �%9��O�I�'*��_$:�D·K�u]�Y �h��4ܺ�{��"լ�&?�k��'Ь���^�
͊�m��w��=�b��	����؟l�IF�O>���p%*`ɝ(�~�Q��"N�R�r�|����O6��妱�?ͻ0xI7�W�f�H�/C<B��HΓ�?����?q���1�M��O���oQ.���"�.�7&@o���"g�SO�R�O���|����?���?y�h
We�:�rA抆�<0K(Oto�1P�v��	ß���B�ß<$Ϊ#�\4Cg�P�Y6D�"�!֧����OB�$5��Ɂ#=x}I�߫4���%'L�
�"�ߗa�h˓1M�D����O�!�O>�(O���g�\2{�
a�1��,{�P�PcG�O����O��D�O�I�<)�iz�ĸ#�'��i�Ef�$l����d�F9�#D�'�P7�-���OЌ�'���'���Z���@
�L(�H���IY����d���?Z�e�e-�?&?���:c� U��?5���B��<�r��ȟ��Iԟ��	���	E�':���M�"��!���n�6l����?I�(�F����'��7M*�d��$>9z�bD4C:��ҙ#�"�O����O󉗥i#`7M-?�`-�d��L��oԂ[��<0��&o�����	wy��'c�'��D�L��a�ŏ��&퐶G��B�'��I�Ms�&�?���?��'�r�ON̰�Bo�+ �\��ʐ�<��H���՟8�?�'�?�b���>�H�b���@���F	?6-�	�C�V)8k*O�����?�� �d��3���j�@�fZi#훫�����OH���O���	�<i��i���¥��y�� )��Y~��A.,Xr�'6M.���O��'0�I 3h�cW�B�q�Q҇AȘ,_�'�r0���i��i��bƂ�?y�U�� ��r�b��� ���hq�>O���?i���?���?������ȗ*��J��	9Y��u��HD�\���mZ�^��)�������R�S��������*Dt��x��� �N�V-@��?A����Ş
j���4�y�-�2^�;� X&Xdy 	G�y�Ũ3�y�	��'�	����	0� ��60�5�GAڨ.>��������ڟ �'�b7�B+�����O���̺g �
�c�SF,��k�(���LH�O �d"�I/-�XM��M�jJf�jp�R�6Ɔ�j��� �E�zm���O~b���O����@��A`������%G-& ����?����?����h��d�3Db���%��>S�*9���V����������S�\�Ɇ�M���w�p<�$Li�� Ci�k�ڡ�'��Q�td��!�'�� ���]�?)��,@Bbؕ'R�@F���/vX�'F�I֟��	ן�������	!�<̹�Ọ� usF��m��'�26�Y
�(ʓ�?qL~
�8����éh� ���-# D���6S�D�	̟ $�b>�	u%�6&��)�/z݀!Jd��w��Db�	+?I�H7��d��䓵�K�Ve	AE,O t�5�DN���ON�$�O*�4�˓m�VD5��ݍw���z��W.~�"A��� �y��nӔ�|�O����O<���W�6�Q)DQ���:<f�j�x�����tg��P�>9�ݸk�&�ӧbݕH�xQ���͂nbt�������⟼�I��<�IR��W��I2BާR��⥆K�E<�Y��?A�CF������$�'d7M1�DT�#/R���]e/�T0�B+&�@�O���O�M�a�6� ?��/��3��#1��K�� bΌ@AoW7<r�$D�	wy�'���'�2뛗|�����XT
*]��f�(Y���'��I��M�� >�?q��?i+�*)�S�5q$���I�,L�ZTsԙ���OZ���O8�O�S�N����g瑝_۪�Vh�1��l�5\ �l��4���B�'�'&aW����нZ3k��Qb��AG�'"��'�R���O��	�M�G�� o8�*�@��)��+���r&�.O��l�Y��)���Lj�͐�K�z�Zf&_�8:��3�ğx�I	%�$�n�z~�������L��S1,t��BA���R�B�((j��<A��?1��?a���?Q(���f�� I�J�RD͟"m{Ĺ�EG��5���ɟ��I��$%?��������<��L���B��\u�dbp�D�O>�O1��	k��kӖ�I�,.�Qs�.��]�p1�c�٨�|�I57�ұ�U�OD�OZ��|��,,Ʃ�SG�9�T��a�2�%(���?���?�)O�dm�8}�H]�I̟$���_��+���`]"�c�G�.m��'�������$�OD��<�ĝ�*I�E�6)E;/r�%�1�\0!��	�v�PaCA�ڦ�2M~
�����	�����1�޹�bT59������	��Ia�O��a\܂���<tH��D�H2q®m�F�H�΢<Q�i��O�N��)��T�#��d̔���Z*$���OH���O���l�B�2�~a���?Y1!(܂Dh>� d9+��@в��G��yy��'RR�'���'G���*B�Z�	�q���z �i���+�M#�L��?����?�L~�d�ҵ��V�aAn
�C��M�`Y�4��П&�b>�"�K�B[V�y$��g�~-2�O �@�)E�Jy�Ȝ>���Ac�'�
��83 _�n�
Wm�F`Ā�I��������i>��'��7-�.c:�$�Z^6�s ΍U�	����c��H����?��_����ɟ��ɳ#a�*JU1��p��	&`hL��f ���'�P��H�?��}b�;[! �����-���I�*�4Γ�?���?���?�����ObP��ad��g��xS各��٫c�'G��'oV7�?7t��OL�o�X�	(D�ZE>9�7�(����� �S�	�X�i>]����1�u��H�~�P�P�!��aѺ`�g�\������'�%���'nR�'��'������K	���C)���\�s�'1Q��2۴;������?�����[�;@�R��R5g�z����[������O��5��?a��>�b� �%�'m>��V&\��XfJ� Q���|j�L�O�@KK>��ҁN�)'їN�Zp��-���?����?q��?�|�-O Hn��K��$���1B�y�V�6����D#Ksy��t��㟬y�O|��J�5}�x�Ӯŋ �Ԭa�� !YM����O� ��g� �Ӻ�.G�2���<ի� V��=����7\L��`�<q-O���Or���O��D�O�ʧQΰE �!�::(t����j5(�$�i���S�'���'��O�B�g��ī������9B<�@�DA>q(J��>�)��t��tmZ�<�V$��kD�vj�dJN�� d��<���Fm�,�D����$�O��D�!I�X��nG���j�8���D�O@���O��F���-K�~�"�'����>�<�Ӈ�
	}%*�a�,Irn�O2�'���''�'�T�Z�@��-�2��p��	N\�	�Oe�C�Z�C4,6d�1��$�O����� 0��qv`@�
;����O
�d�O"���Oڢ}��=�2���`��}��	f_�ŉ�	1���81��'�<6"�i�5�bg��,3�Y"Sk��"i���c�j�������	dXbPl�n~���rs�T�g�? xt��M�g��� �f��;�'���<�'�?����?����?�6'� LXr��R�B<L�B9sڀ��I��M÷.�3�?����?�J~���3j����A���Ԫ���N�<y0V�t�I͟|&�b>ź�m]�[�x��P!DL�զ��B{�H�ŀ�uybDԍB����*��'��I�w��4���Ƥn��C4-�#A�0�I��8���H�i>�'�H7M���"��.���	y�ʵ���
]���V5�����O}R�'���'�|�wL_�/$�1 G��4}HόF��f�����%E����+���{���a�`��+I�	Hb1O��$�Od�$�O��D�O2�?9��ΎA}�(dH���k"��ҟ�����{ٴ	-R��'�?Y��i��'�x�bم�1��*.�a�@�|��'��O����i/�Ɂ|a^��  �E$��Pe��n�� �`�)a	��.�D�<���?9���?�d�-E�AǎvN��ac-=�?����D����
 ����	����O���c���>���Ƈ$?8�A�O�P�'�2�'4ɧ�Iʈ=�E�ǯ¿}�B����2g'����׈w���ל��S-���h�	�	����!Ým�"`��sn��IƟ��I؟��)�SPyb�g���0��W�|���?p�9x��O�x�t˓&�����}��'�derh�F9`�T]�:e'P��dG_�M�'�����!��?1�%[��"�f�Ja.�iы��:���x���'���'�r�'k��'u�S*�=D�iGn9iU�ŀe#�|�ٴW�x����?q���䧢?��yg��q_�k��׊KϾ�kM	R&��'�ɧ�OX����i��׽	lٰҢ��H���C���-�t���x?v�O���?���+�K��;Bd0t*ō=T�p����?���?�*O�ul��8v0(��֟��	!"�8 +�7��Q�$ ƾyi2�?Y�_�8�	l��>�&��m�l��Q��ȟ!����'�E�6	̟"fCT���I�ޟC��'Z|}��h�/tjsōO,�4�@��'�r�'�R�'�>u�I���h�7E���� Ӣ��;4���;�MsR�ۑ�?��z<���4��ڔ��>���I�_�x�6O��D�O`��ۇt274?�!��u��S�f�8��՞gj����!/!��&���'�R�'_b�'��'~V�$�Е
^`�SCFo>тU���ܴv>�}���?y����<��>q�t1��Fטlm˳�w3�Iퟴ��^�)�SB�$9sAk�*��9BC�cJ�Y��
+����'�A`F��ş��֞|"P�Y��;�� C����M��Z՟t������	���~y2l`Ӱբf��O.����X�´���e�<Z<���3��O2�oZt��d���������H;�"��XC!FJ�S�d ��$���l�P~�LHN݌���h�'�3��P���b���#���<)��?���?���?Q�����v�X)���P�?*:��0��	UB��'��!v���)�*�<��i�'
�Tx�A�E�0��e�$�|��'{�O�j r�i/��8;��q����j�j���k
��ࡡ\�7��4�d�<�'�?����?	������C3�ܔ~�]�׷�?�����Q��=`�/�ޟ �����O��90M�����ˤlH�h�N��OPt�'B��?e�j,r��Z��1�hق�`6��qa$����R��$���`KU�|���B�:H��,�@���$e³&M��'�b�'t��T[����4b��1(�C�ۘ�i�eŜOhD��U�X�?��+W�V��W}��'���A%S5I��c<���F�'\���>V���tɴO%q�V C�j�F�zuCF&�_�3>OD��?���?��?	����)�"�"5h%�0+���Ė�Lɾ!oZ6�ƕ�	�����{���������#k��^��E�J�`H�a�]��?A����Ş=��!�4�ybLѠw�LB��L I%��0f���y��4D������d�O���Jv��ebΟJv�-�6o׼A�����O����OL˓ ���#	�;��	���c��\P���N	I��iS� �x�a�	���IH�	#uj�����91ȪPZ����>�rb0U�@D=>;z��|.�J�䖭�?�る�2��ǡA�_�.��Do]��?���?1���?!����O|!�ă�'?�<�!堒3oء��@�OF�n��K�X�I����4���y�O�7M��9a���ʝ�����y��'f��'_��hP�i��ɿr�&Qi��O�4-�d���_z1`�̀��(	���R�IUy�OZ��'H2�'V2��u�>�5!�)h�n� ��Q���I��M#��T��?���?�H~Γx<��A�D?hy���NN�Vg�	qS�������&�b>�QSM%5+2��M f�@����=6��SFly"���sc����
��'`剰X����L:kĎ��|�x�����`����4�i>=�'�B7-ѽ9����?l�hH�D�@y���T�o��$]֦�?�!U� ��ɟH�	�?����*�;7>(�R �<�*��ڦ��'�@2����?��f����wL`����[��wm�vp��K�'���'�R�'WB�'��f��AŖ6I��Z`�K"3�����<���0��f����t�'7--���x�,1�Q�јl�6.��FN�O�$�O�)�R06??q��e�? �H'V�#���)gL^�H�iu��~�|�V��S��Iϟ�)w�	@<�\
@W.�n��3��П<�Imy¤jӮ�{�d�Ol���O��'C8.E1�E
��XQr��CVH�'�^��?1���S���g$.�q���2G��΍�N��y�Bir��i�P���xg�Q�	�l&�:��K�b��)�D�,Mh0����D�	ן$�)�Xyb�~�.Q��"��c��ꗀ	�r{���I�u+�H#���J}��'Ov��F��k~�m��
�9ͤ����'n�O�_s�������욚t_���<9�J�R��2�1E����uE��<�,O�$�OD�$�O����O6˧b�R�!�o 1w0mP�@Qm������i%4Q)��r��'���O��'`47=�ĥ�c��qzl!ĥVL���%@�O
����	�ʐl��<Y'(�L(>p��?TD��"'X�<Ʉ"E����T����$�Ol�䂗q�"��G��|�N�zwb�����OZ�D�O��=���L^r���'�֟L^P�Qgs�����=}�O���'|R�'��'5l8���Ԫ?�֙K�K�	@#���O*��LΜ,���[v�/�	L�?	v��Ojp�c'��JJ�,PfK�
9h� ��O|���O����O4�}��*�X���C�XG�<�V�N�(�t���UЛ� �'��'��7-5�i�m�&�� ���u	�Q6���g�X�	���ɸ"2ԨlZE~�o��mxB���r	���οRI��0eF��_L`�E�|RV���Ɵ@�IܟT�I��
����Ѓ�R�h�lu��hy��j��}3q+�OL�$�OR��H��_؝ A��O���r���,6�"��'<��'Fɧ�O����K�S�����7Z�Hj�jH%Ū�s�[�`Y���� �B�Q}��oyRd�&΢�b� �.\oT���3S|��'b�'��O��	�M���)�?��,92Y�픭GH�H4�K��?q��i��O���'2�'5d��F�p�N�R��頏-�Qb�i���>v<�P�۟В����y�f��2m��t&ְ�6 �	O �D�O��d�Oh���OL�d=�ӝ�v��T)���J&,T-���I����ɥ�M��F������̦u&��b�A�R�.3犨��钰D�B�O
���O�V?�z7�9?91Ĕ�2��IPAcX�${P��!5-~p���Ob��I>�+O�)�O����O�#��ܪ,W�	q��p�R��s��O��D�<��if2��V�'���'��S:,��xQ^�=���q��u�I埐�On�$�O.�O�ӂ��91�J�$���� (8q����UnZ��4��X�'��'�,��-�Z*(M0�M�ryXY3%�'��'����O�剧�M��˙=V�*x��@�
��x���&4Y��{-O�QnZf����	��C#X�LE���5��5'�`g��ԟ4�ɲ1�V�o�z~�(Sl�t�SK���$f��+��wu:�	�
�f��$�<����?y��?����?Y(�@�q�+6�ť�5"1(��dk��J�6-̻w�����Ot�d%�9O� lzޑ[fe������Y�d�"Q�PCٟ<�I|�)�Ӯ.��n��<I��պ؈	�7I�2T�*-��+[�<���� s�>���"����4�����{�u�Ǩ�2M^�� �YV���O��D�O4�{�f�&���'�Mξ@�|�QK�,L�!H�'�!"��OVi�'�R�'��'�m��cשw}�C�X�}�d���OZ��<!���@C��<�?C#�O��C�I�f��q�׵
y>M���O��D�OV���O�}�~���F��FtuRuh����S����ٴ*Dpr-OX-3��O��ۖM�J��3E���Y�Oŭ���O���O�%)��t���Ӻ���G-��T�)B�̻�(f�0A�k�o��O����O�*ጥsO��ԑ�SC�����4,'�����?Y����OR��x����W.����LL<}�4��!Ⱥ>q��?�L>�|zv��h�.6fK�w�j@1��B���i/��a��
 @���$��'%|��	4q�p�ӛ6�z	����.�7 !2�žP"�azk; �=S�%M�y��{�f㟼��Ob���OB�Y#��]$f��W��|�0ĭ/���3wnsӖ��
��v%��J~J�;Is�p5G�]�Z2��W�L|���?��[��h���#��́	��B��?i���?aQ�iyt<�͟��lZJ�	?2R,RD��Ȅa��ȮT�l�'������擭E
dnZS~�O����Gy�xpc+,�e�⓬}���������/�	}� @!lK���MRk['S�#<Y�it�@U�x��g�ԁN-Ab�bw(ǣl���B�����L}��'�2�|ʟN]�F��?�����R��4�Ǭ�E�z�D��}����|BU��O�3M>aԎ��`; �4Z[4��I�D<��i1��J�
րl�Hl�G1~
��۔�9$���'��6�!�I��$�O2i��BW�i�S��9��-Q�'�O*�d��F�6M5?��c���oyZA���6 ��z�Q�"X
�y_���I�j���OL�J7�	p�/��B��ߴkPČi.O���(�Ӣ�M�;1�`u���(B��R��?Ҫ���?�H>�|�%�K��M{��� �d��	תl�j���.��l4�E9Ot��I�8�?�f:�$�<�.O|	��ۮv�b�b�L��;�����'�.7-�+ZϬʓ�?��h��=ی�"��,H���K�FƷ��'����?!���`��he�!<f�h
@a�4 ^��'z�T�$E@j�@�R���T�ǟ�R�'u"�ᡦ�B�z|��a��R�'F6��#M�.p����!`���Y��'�7���K��F�4�L4P�����I��ݫ�C��yB�'\B�'��x�i��iݵ��A�?�Ȕ�1P�u)�Z�D����KU� �'��I@�'Xrt�E%�|�X�p�TF�d� �O��mڥT�Y�'Y�����N����T�j;�e �ɏ�m#�T�'g��'|ɧ�O�t`p񍙗QAD-�ELD�Mx��dY�]�QQ�P��9�IO�d~�EP�VynY8"�
�)C`P�I�p��&�̹�0>�E�i���1S�'U8k��ׄ]6�@�d�*i3bp�'�j7�&������O����O$�{�ȟ0:
����c�Թ�C���6m"?A�
�C��������ɿ�ժ�6���I�
 i��P��<i��fE.`$D)CKVE1�A���-B��?Q��:0���)���
Ц�%�����}��Y��Vΐ�ᐡ�[�ԟ�i>1��������'lv}A�#'-m�I�� 2s��4:I��'+p`������(�I�76��N_�TU�g*QW�"<��ia<�$�'���'��d��	���%( �2��#��U@�	�H��Q�)���=a�8�=y�z ��jř.���9��E��M�[���m(�d>��R�c��O3!ԼB�ËHQ!�dTᦱQ�.�<�	8���)[�  �	#w0\�'��6m!�I�����O��$� .H�%�slh@	���Of��əI�
6�&?�;H�-��'m��I���(�t���U�\fv����7|O��1dFL�E�����
ؕR*.�a3�Lצi�m�۟���\�:2��y�o�7,��4m�>>�� eR�:}r�'�ɧ�OVy�p�i\�d�!F�l��G QK^b fo�0V���:X:���'r�'���\y
�/uf&	��H'��]AbkW4�0<��iBN�y��'���'���G�ԚCF���/�MЅ� ��x}B�'Zҟ|��C�Jb�`�#�#@�"��'�]����G>g���Ju�\�$?e���O����)_�6���
d����(X3�j���O��D�O��d6�'�?!uo�4N����L?��E ��0�?aŸi�Z8*�W����4���y��
4g�D�Tn�/	c���yB�'�r�'�|� �i���	As�d���Oڜ��h�!2� ��@[|-QQ!�n��Ey�O���'R�'���[�#i����GN�yXr��%j��H%���MC�͂��?���?�K~Γ��H�%Mh�VYs&+�'BQ���[����۟0&�b>����1h𝒴�Q�'��:��'se�41!&:?�u�H���M4����ϱj�)���S�1�Tazp�f˸�d�O���O��4���\��Fie|B��g��<���c��4q���+�j�X�O*�ēW}��'\r�':\���!V#3�*�c�č�� ��v�
�K�����(@��7�t�Lg���ߙ�򇑹B����1�5��uSu/w���	�,�	�������� ̠yj����AN)S��sQ�v)����L����M�V��?���'�MCH>�B�l����1/�$jd��;b�����?9��|�c'���M��O�v�;1��YX���% w�MF�� $��M��yB��3 PX�r�+Q֡�V�q���0Z5ᄫQ��횑΂�A��8b���(*�q�qD� f��{7�>\��ia��"3�b�0i� @Ɵbi�3 Dp}2�ƻ^�ҡh0!�3`�	��fܯArl��5�݋c�[3w|��eF�R��͈��S4p��ӆ�&CZ<�tm8o� �j�N���߱{�1RM=c�n�@w�2_4&��j&[�̠��l�	b��S�ԧo�^�D�@�9�����F�%l5�Q�ކ�,MS�Sʆ,yÅ�"M��b�;�M����?����21@�+ḛ�& F�Gp =�r����'���'�����D�?��+?��)�@̈/�j��q�`�`�*x��i;B�'���Ok����� ̖\sfŖ�:})V`ަ���ҟ������%���}
fm��P����� �P���%¦���۟�M���?A�����_���'t@(�	�Z�QTkB�!\\��j�z���3�IO�'�?�FL����/�V�AՀ�1 -���'D��'Њi9�ȥ>	*O��d��0@Vz�6�y�kƔ*�<��e�@�Oƕ�W�J��������{�L�'���3���g�H�Jq�i��dU�\Jh����O�ʓ�?��>��@�!�	z]XL{v��&�
��'kީ��|��'8�'���$��\��Ųu�m�FȌEP�q�Jɇ��ĳ<���䓥?���.��U���-����K$z{$A�p*��?�+O��d�O���<a0�T�}��C<lY��11
�+�x��q&��l���]���G��ɟ�I�>��`�)H�� �^�d�h#�	Ǖox�'�"�'�[�0����)�O��R���%�W ��e�O�9�Ir��ߟ<���O����u��փ\p ��� D�|�� ���#����'��_��c3�A�����O����2�� �M�%H?��� B����1�xr�'3`�c�b�|2ҟf܀�äa X�0@S-c�8�@��i��	�e�h�!�4�?���?!�'S��i�E`3@�;"��@`_N�����v��d�O6�-wM�O��>]�a���La���/ �%����iӼЂ����!����`���?u��OʓS|
���h��C����%��,?��A`�iO�T���'b�'��p���#n��()��V�PF�9�qi	&�n�՟�����̀�a����<����~B�Ls��у�*�	���C�HA���'d��|�'S��'L̕��T;a������\�O��` &�o������C����'��	ϟ�%�֘��Q`�  �=���˘s��I��N>����?������3�¬�@(Z��z0�-��I�)Z�ҟ���b��RyZw� P�`�ʀT�>5�QQ���4�?q)O��D�O���<AH�u���ٸw4M�5#� +=.�0��[
}��	�X�Ii�Imy�O�⎖q:`�����Z�;�B�kw&��?A���?�+O(�{ƣ�K�Ӝ�\{ �1k�YB��9o��P�޴�?9K>�.O�	�O��O����Ҥ�)뜔!)X�n�����4�?q���d�> ̾p%>����?ט��x,s��v����C�Q��Of��?����<��X+�m0v�Nz�y�F��h�osyR� ��x�X�Ou��OȈ�� Y⒩\�r��E/Z��loZ`y��'��e;�)-��i��Q��� ��0
Gd҇T��h�4~�pyJ��?)��?!�'��?Qӂ�Hzv윞�F���E�����"|� �</"V񰦮��s'D頡��5E~��'���'����X����ɤ9"H��'�1'u���+�1��a���\�'�?��'��'�0K6�����%/����4�?����"��d�L����8��27�]�<���@�	Z��$����>?	��?�����d_�i�����TB}&�sdHÒB\8� b��|�	Ɵp�Iy�IFyZw��Zv�
�8�VD�'c�NX�ٴ�?iK>������O@���B�?��T�<� ��E��T8)�a�����O:�t�	Gy�f^�MS��Îp��y���!$�1 �l�s��Ο�'"g� =�S؟`�1���u�8��)�9��q��H��Mۏ�'��	�zB�Orl*F�N:b`P��EW��鶸i�bX��I+�4�O@2�'��\c6�� �ֳ/�͉��d����L<����߹vI��]�GE���Q�ؔR؊�b�E�*�f7��<	w�E;|	�fm�~"�������|�g�A�@� ��Ƥ!���~�N��?���@��O���M��"�}�48���R�W�@ER"�Ц�ѭX��M���?I����P���')�X��C�b�F��%(�<R0ֈ���g�,c�9O�O~�?��I	�L#v�C>4��A@Ϗ�]�05y�4�?���?� R�ZL�I~y2�'���0_�%rD��mH�գ��M���|"aN	�yʟ��d�O��׿o�9з؆P�N�X6��m�XmZ���sHѷ����<�����OklY�y��R d�C���T��"eݛ��'vN�1�'���'�R�'�Y����O�X��0��A�6N�	;��%b&����O���?�-O��d�O����f��:sDC6c9��ō�7V]�}F6O0���OZ�$�O��$�<!�K�\�I�V9D�!�َX� �E
�m\�FZ�@�	kyR�'"�'i���'�r�R��II�t�		v�,])�'v�����O��$�O�ʓ
�0���T?��i�ň��	�TP(��E)�Ę���iӰ�D�<!���?��,����ܴ9�L�8Ć���<�m��s�5l�����	\y�ʚ�qN\ꧽ?�����ƋI�>1���
ZV`;�՞1�����P��韸jS�l�@��y֟@0X`�ް%F�d�����fOJ��i
剦d���`ڴ�?��?Q�'`O�i�Q�3i�$(@T�*S'@_މ)�.h�$�$�OD�k<O��O�����i�7
Y��|�`�#�vѾm@7M�OH�d�O��i�h}�R�Pwg	~�&�10�R�<�{���!�MC�^�<�,O���$������J2r#���
C�B��@u�C��M[��?a�Hʢ}�Q���'���Ov<�e��[��@�b�I%F��e�s�i�b�' 2L��yʟ����O��ė9J�h�4���Q������"h�l�џ��Tȕ����<)�����Ok̟�a��Q�<������9��I�(�p�ߟ���ɟ���֟��'�L�!���M�*4����[��	�2��듕�D�O���?����?ɷ���$���牃�l��9Yѫ$� ��?����?����?�/Of��\�|��� ���IJ5`e@�#K��1�'32[�4�	�����0x����3�ʀ��؛�
y��#�vxڴ�?����?q�����בg�l�O�Zc�|� #V�~� ���0M�!!�4�?�/O��$�O�$ѭeB�$�O��I�R���Ϧn�J���aF� 7��Ox��<I!�v*��l�I�?QH1��y� ��w��%X%�C�A#���O.���OΜ���T�'��)�;�
�@��G�xH�]��_����*�?�MC���?���2S�֝�s9�1�:sM\ᡅ�s�:7�O�����h�$Zg��'Nq�F�i��[&.R}� _+,x�aKոi�4��ĎcӨ��OP���(|�'X�I�� ��C䕂s������3��lH��i}���'�Q�����D���Dc�*u�0�B+X��H��?��?���܁G��zy�'���p;�E��'V�����M��f�'���29"��)���?Q�p;�2��?x�H���5sjv�jw�iU��)�p���$�O���?���؄Q�g؀8|�1�4�ԗ"���'W����'��՟��	v�]"��!ã$Z�͹�m�=�N��p���<1���$�O:���O@�����7b��1��g�I`��˵��s|��O����O�$�|Γ{'xi��0��8�(�9~��L�P��,�D��ði��	ޟ(�'���'y��V	�y�J�v�b|��Σ0��qBB�ޠ��?����?�.O@TH�|�t�'�b �5���Z{�����W����m�D��<y���?�s!b}ϓ��O�u��-��I�:l[Aa�*h��l������Ay�K�u��'�?���ʷ$��e:j!�aėk�:٫Dȁ�l,�Iϟ\�	�, �io�Ԕ'��ݟ�mjv���]��K:nJ��������Z�mZ���	ϟ�S����5	�>{hL4I�Dtzd��i!r�'� ٰ�'����y��č+�$3�/�ݪ�FV/�M�F#�=���'���'i�$ȼ>�-OXAt�A'0���$TE���bI�̦��v�c����Ty��	�O������m�L�z�bG���a�&��ƦA�I���I�!��T¨OL��?1�'�8,�UK'(^�H0��.v ex�4��1���S���'9��'Jd�i'B�6'[��C�̂rw`UX�y�F�d]h	hT�'��⟜�'�Zcf�a�;4�,т��
�JLr�
�O(��:O6���O����O$�D�<a� �1�H(�o��X�i4�ܤ[-����^�8�'��X�<�	�\��V�Xh:�$�!jHxf��{�n-��`��	���I���	`y���9[#D�^6�]�e-4yھ��6�B/�,6ͧ<������O��D�O4P��5On`�3�Ͽ2�����:�X�@E}��'vR�'��I�i= ê�B��ϿmB�0���LVA��F؜
��o�ɟx�'���''RnU)�y�\�anҾRVl@ ��ڝ5Z��s �/�M���?�+O��:&i�i���'�b�O�J!6C-!� �)�)�D��D#��>���?���w��ϓ��9O&�S?$6p��+ܚ|G�$���N3�
7��<qu��-/t���'-��'�d�>�;<>��ٟ�8Yf��Zn��4�	�Lu\�ʟp�'�q��H��J�"@]G��,"���i/h]aQihӤ��O����� %�t���X^�1��H�u��BՃP:���۴�� �����S�Ou�
D4%��v�ԢO\z�� ӻ	�7��O��O�pr'!_{�IןP�	z?�[�`?��cN�%�`�9�B�Φi'��������'�?����?���c)ve�E�J2R�@P�G��	�v�'�\Aƅ#�	�4%��	 �zT��S�&=`% �.�"I��J������$�O���O��z8��A��k���p�I�EQ�m�N�bW�O*��:�D�O(���(��H:p�^?q�,���Bדm��ّd��O�˓�?���?�/OD)��n@�|����%A�f-��`�/J�\k���\����%��������(SٟT��"�S;D�ó�[1,%+Ղ���$�Ot��O��~}�%sW��d�T;[��"@�I#��PR�ؾ:p6M�O�O>�d�O���2O@�'2尵G]�&��5$���MY�4�?Y���
-���&>�I�?���KEw��|yr"��N���	�`�!�ē�?���~gD��������1Dd�h�pg�)ej�K���7�M3.O2�A���aB��<�$��^��'La�UC�?F($!�@t����ش�?��%X��������O�]�3A3�����ތn�5�ߴ4�LW�i�"�'L�O�b�@�#��#vw
�"���F�^�M���$�?	M>q����'�؅BF��~蘡�$��l�zղ6�fӠ�$�O��D7p�V�$����ğ��T����#ب�ҔS��ʕ��i�'�)��.%���OL���O�[ ΁�g,F�䪑� ���%o�Φ)�ɔ�^�	I<y��?!K>��: �-ٵJ	�r�܃��Hv�a�'� �|�'Y��'�剹3{4��d�R������,�h���@���'�B�|R�'���6'����2�_a&��+�.iv����'���I���'����w>�
�`�w&ik��V�Q��ʦ�>i��?�H>a���?	��<I0�P�h(��0-�Q��)���׿3��I͟��	����'�~}˱$3�	�	¤hy�fʃK�� �'��2:^�m�D�'�Iʟ`�Of\`���H���f�|�D��t�i��X���I�3g,8�I�l������'D�����}*�ӂ�Γ��I<�����:[��ݩEZ�I#�KR6�T�iD�g�7m�<A1m�<��'�~���
T��x�W��'��}�3K�qgZ�C�/y�H���O���P�	l�'y;�$z���n���z�Y�&��ش�v����?).O>�	�<�O~�1�PE��%��N*a)�H;A+�>aBS���O�r�P�%�\�3�+��W����V!��
md7�O~�d�O��iF�Rl��?)�'r����󞴫"�@,Htq�ۓ�?9���?�G�E�������8?�d���M�*[�6�'�,�z��'����d&��8� $b��W �XJg�P7wݞ���Iԟ��	🼗'�bxywnQ�X�f�2vn-U��L��C�wO$���O�O&���ODK�)ԃrw�]8E+�OS����K��1O����O�d�<Y�A�.]�i+ʆ hsGW%M"FiH�B4*��	ڟ���V�Iڟ��	�	3(�D�|��cn�  �����~^�t�'���'!b�'��Ē�hB�'S�I�2Ԋ��H%�E�0bZ,��F�'F�'YRP����=��c�*�����2�Ĵ1&�ē.z�6�'�P�x��ħ�y�'k�20�4g��X�1av��*'d���i��OB�(���?7�۫y�e��h���=��`)T!�&�'~Rn��'���'��I�?�����֘�� �ga@%4^T�ZG�ʵz6m�O.ʓe�P(DxJ|�W��9[�%��'s��������yp",USa}� ��i�$ȩ,תJ䶬�Ɗ��y���'i൰���-W6�k"@.cH�)2�]%��҅�F�0.�0���-}2��#��#K4F4��C$w`�rgoCS~�ɚR�ݵs�@�۔�Ԥ'�$����'I�����[�&���jFGV�i���ڻo�0 �P.3�N��do23����OPF� *ٻB��Ђ�_ A��'"�'���ԟl���|�@ą�6���/XaV6ŐWdئ!6\�-˶R��aucӗJEn�S����[-�����
_|~,ڶ���u~�d���T�(H�8��K9]k��� �=��O�IA�G��g�h�mڰ1a�H '�U�L\R�'�ў��?�t�>zfx��6-c�����d�<y����XGLA3 )q ��J���i̓���uy" ԫd���?Qw##O�\�8�%O*W|X�Bs�J��?q��'�����?��O��D1�H]�h�ː¦����fIh��ѻ�����E��1O i��	�(k��H"�L?�Eo]�1���	���yI@���a8�@b��O����<�ķM�hi1��޷c*@cQ�a̓��=�"�)��Qt��[�$d)EϗX<ձi 8�;�G��k T�뢋��t���'c�	-l�.�өO����|B�/�=�?I�o�Z/� ���9�h�c�D��?��� ~���H[6A t����]H*��˧T�)g(9@�@� k
�k�h�O � �[`��Q`ĬO9 ��#}��J�2d,�L��
��b�i���0��'(�>e��5�N�u�$0X��ҏZ��C�)D��C,h��'�����$Ga�'D��	�7V�\�p��i�l1{WD�>Q���?��nU(nr��?q��?ͻ@�pq!�Fe�JuR&䁪9�*]x�� ���!5�'�x�pn�����c;��(�:ݾ�[Ո��$� �AՅM/�٠�'݆���U�g�	r��0A�O�2j���CM8MԠ���O~򍇚�?ͧ�hOF�97L�1)��R] x'"Oz`[�B��7���)��b�L�u��L8���?��'��ʀ��|s��Ӵ�V4j"�p� ��4J��G�'�2�'��x���I��H�I�bf$���<{��I ��$j
�%�g��+Ϫ�i3�O
좁B^.�,�!g�Ɂv�� N�A����9/��p� R�\Taxb,�4l;t�6J��p9�x��(t�NШ��?с�i-�^� �	M��"p�Jp�E
�+�	(U^��Γ�xb�����,"2J�/Uތ�R.����*˛6�|�2˓k#H����i���'��k�h�HS4^�l�r-�џ���+w}4�	埜�'�b4A�+m��ţ�X�MEE��J����=l�X�a�I[8��S�/%ֶ(��m��l���")��L^(hµ��d��Sl ��D�2y���'L�	h;H�1 0r�Z)�d�܃fb�$���#8���S���L���$Z�d�(C�	��M÷�V�e~��b4�C��y��n��<1���08@��:�l���e��'N��C�ɫˎ��%�φ;�|a �	r֜C�I�>ܞP2VmȌ(7��Y���d�tC�I�RV��Ac\/�L���P/x�NC�	�H�|�zԫ[�V�@C�	�)q���g�@�)�n�s� _vC�I3�*@��,�>*D�K����NC�I�[�@��TK܇7T%��I�:@C�	�b|�����_fy���X�C�	'?�~5�ЍH:If8�s���.^�B�I�;��*�N��Gkvx��E0|W�B�I��±j"�կo�b��UI^.:��B�	6wA�T�V!G�N�śP�$��B��%AL!g�K��2|��o+:��C�	>!���`7��N9�dc��4��C�)� <�q�h��-�H@�c�56�<M�"Ob�@�,P��J���6�\�p"O���"�&����`��Z|PHW"O�����L�p���j;�蔈�"O>ظ�cÀ\�����@�q0"OT)��M5ht�2�A�_1$5��"O4�3ՌT$)�� �S���K��s�"O������O#&=��ǽ��U�s"O���%�
_&:�X�@��2�ҳ"O� 4Ɩ�԰�A�V�;ˈ��"O��ҋX�,N��kҁ?�0�i%"O��Y e�t_6Q��JJ$�<�86"O⸁S�A�JYx��gLO�$�e"Op��G'�9k0	�d�Er�{S"O��Ц�{���R%�%D> A D"O"q�'k�#	��Y�s��aӞ�{"OPiC@�N�[�n��0�,v�t��r"O�d8�F�$i,ȼ� �?d����"O��p7�RP���bJ�!i�RÁ"O���� �P��#G���b��"O��"	:�tR��T�]� T��"O��f�A1^O��`�ŕ!�ڱs""OV�sj�"�����Mz�Pj�"O��@
�E�Ph��S
P/��I$D�8�Fk�!R��	�i�o��q�g�&D��1Qj�3"()#��3HS�X��&%D�L��ļK�HX+B��$D{�l��'8Z=8�MI�?b��,Z��d��'j�}��%(8鋅
�5�
�"�'ژyÏO�o�̀u�U����'�t�`5��M��������F���' ��(�흪un8be� ��'�ڡ����j�D�':�`��.b��L��	i��dE�m&��BF�4�"��b�݉-��~�b
�ś�a5x�D*Є0�t��E)��?QփF3L����g "�y�(\| �-Rz��C��D�1���	s�����B�����(Z]��bbX�&�!���t)���@)�>9[����@�.D��NI��	%�H0y��S%C6��x���# ۮ�bA�[�JB��t���#��K��|3��\45J���?�?�O�5�~Ғ~�?�6��Njd�c޼�8�W�҄�p?�!���@xdÇ;`v� W�D�jE�"L�Ol�CvaF�ܰ>!!�]b�1eJ�,RBA���^��T�'��Pl)*���9����!�b�p�'��+aD�����H�Ez���
�'�(��D�)fz�1�<	6��������'R�>��BKYa��Sm������nB��u %	��O�C���Q,͟7�T�QUB� ,��9��(q�"�:Y|,�"HV�k|D$���|-�&@F�+�D%�]`���2�[H� #G!�T^6���]�N�[a��4#uHxc�䝑L��U&����l�c`ĩ���	����Hj���3eh�6o� $y��"O�ݪd��mOn ��#ڊd���l΍
=���⟬jD��)Kq��'�{��U�� �O�f�rXs	�'zy�Gru:-��|�${E��[���#S�Âx�(��C	?lOnqB��ȼN�;%F̼�=!��ɮcs93��8qsr�X����n���؁( �W�4Q6<�d�����O<uPq��h�O�P�9�.�di*��2
��H�0E��O�UHmu�`�Я
q?��ȦW& a��S+@����,��L�>��T
�4Ef��T4)��3��z"_�tq؜CAk��1�����Pyʤ����D��#���fW9]�hp#F�t�r��cf�d�\P��O�;��^+][����ʁ*��]
�E���бm�Ja�F|�_�Oi0��'\<D� -%+�h�B�Z0~bjD�@�Rk��P�
�&hd��#�V�O\<E��>	�O�W	�'f��!� P�2Ql���K4��'
�]Ɇ�T�O�<0� ����i[3P�Bո2#Zed\ �fڮ/&B�)]�s���|�	�4�.͋�T9Y�������i&l?���X#k�@H(أ��'K�������n�1E,t[�-�$}`�۳�p�>�y��@��YA��}na��'��Z���5$�`���<��㞰�燛36�h�)�ā-��|���O�#C��N@�d׷oQH��ዂR��o�?}���;���E��'01n��T!F�Ъ<���X:�,x ��-�b��I�r��t9`[�x2.!	�ʀ�U�
LK�(1�ȍ'@#B����;�Ш´`�#�\x6&Iʁ�Q%�$��h�J��CΠ[�G�RA^v�p�����?I)��8$d8�I�uh�{.�T x���GJ�3�4��R�i̓sZ4��V��Wa�`J��){�ds�fP�x�a6�G�T��5��L4e㞬�O����g��~���d�1W\�`��Wi�Ɓ!7?n��b!��w�n��j-6�\��u-�)�qO(��'N35�"�rh��<��6�'s�S(� F���Ǜ9�)�2+Wq2�	v`�_9<��2E��
�
Qp$�!�&u��_Q�j��d� %�| fcB7p������^*@��'3�5+SÙ'f�. ;�I�|ffL�0E�R�xa���s�E�gb�$)��4)Wˉ&)�O��8�/L�r��0��H�F��S 7d����S�hp8��"I�m4�1H��Wf@6�'��$H��.D�6�+�(��LU J7|r��	���>q����n\�cS�y�	דc�|����$!�pɳ�/�X�R���P�N�J�Asޮ�ON�H�I,3^���q"� Y�A��D��(l�i�B�Jp����&g]�O�x��I7�"����+U�0�)őx�KK�!i��t�X�e�:ء�G�8<�E�N�� ���X�a��x��F��V�����H�U�h��G�7x�DYe��{��UXч���ax"�E��l�0ODc4�T	d$E�14!�I�J&\��8ED�ă���:��٥�Ic#��Kk|�̻@��y��\��|C�D�	�~(�����.�R@�t �H ���0}��x��G3
1VM>y��WJ�Vj�$rlL�
���iܓY8U�pK-Bi�A3��$R��%�I�	��bL<I4��j�n(�A ](�~܂@��W?��E��J���I�h�4-�p�*���YŧD0(�%�"D#\Ovћ6���`��=Y�k?u�z|��4Ohy"�αQ3V�Q#��7y�vЙ2��$r"Hը6! � zڄ���Qi��ф�Im���`��Z�����=/��MN+{�F���E�F$�e�V���CK^;WF �3��@�B ��hK�T	S�܆&�L�#'퉎=�0���4�5B>�� E�'= +@��1 L>)D��&u�0)J�+I*,q���Pܓ#P8|(@�'j�Z��io��ϓ9�Dx��4�]39Ǡq����'�;p��u�H�e�܈(�08v��C�^!Xc'�T��t!�cT	4�d� 2�[�V� t�$�n�p�(���.R�v��fC��T .��ɨ:<�u���9[�&Us�G 2g&d͆�:H�q8e��L��-��ۙta��̓68�Ȁ'�K���K./z��p�)ʧ��g+	c�8T+�j������(pqCA&9\@��h
=����"W����y��t�B���Un�a���f2$30�ą�w8���G.`!�W8/ �r��K���ܸy��:�	� N��e�� �|2���� f�#r�u��?�(ONݑ���f����]�U@ƥW����6��hC�\{2����dߤ�!�$�<#=�ؖ���!$N��Ã
����qV�
�-��Fꄏ��Q�%"��H�7�
2>���&l�5<ưiQO� �y���=k��\�F`�i������� (ݱ���.��Y�2f_�����O���<A�HA�}�@����Ҏ9�Y��B�V8����*Eې$PT�Y@�L�i�,�P.|�I�%b���0�D�6M¡	�.%���*�$��<@t���ڰDyb��*����"�=dh�=Bp��U��S3S�H�"R���G��9��C�2	�zB�2�l��햝���� ݜ�Z6рix�f�'-e�1J3/њVJD�\ccĐ0nF�)�8��eޞ>�����'���bǭP��4�cW�)9�Uِ#J6\Jʓ1���Rm3�3�	�$$0	�p�2,J�|�pJ���!�=i�l@&N�QGD�`Q��c�!򤋽Urbux2��)�d����$E�!�Ȑ*NPe���P/�]Q"�)Q�!�$ރe[j��҆�9���
TJ!�D�?n90!�[}��%8@�VT��=��I7�э5�ɢ�^�a���ȓBhD�9p�_+�tL� �Ȳ}�����m�T��b��2|�Ir3H[�,��ȓ<Th����Ĝ�"kE�P�40��AC�@5�H�L���%��a��e��>ΩH�Q�t8�(Ч+��?L4؆�S�? z���J����[p�¹ 8>1��"ONxҲ�N�μ�P.�*1\��T"Oh|����_�d��5��?5 <��U"O��1��:e�RU�T�٢=>��!"O@<Q��:Uup,c'�C!(�����"O�d	hY�})&���N�����"Ouɶ�b��0A4^2-��d�"O�]�gԩaM��*��G7Hm�"Oꔘ�.[��=C�#�'S�luA�"OZ��L�?L%�)��%J}�<�'"O����L��=��a"� "[l&"OE��P�0�B�� ��ta�r""O�aX�L�;8�Δ����VWd��"O��heK �6q���<@U�h8T"O$���E]��%�Zi��]���\�y��DT�<Кs ��I�y�c��yr+����ذ'F�I=P���'�y���\�D8Q�X�R9�.޵�yb�R
^�pR`"֑F��� ���yr���H��jp�Ԉ>��]k�y��Z�'�����N�l���۷��5�yb�Y�1�p�a�ͨh�qJ��<�y��A	y�!�%S._$�1�g.�y"N,@���Q�[�f,�+��͢�yBH�9���)[\m� �b		�y��C�UǦ�ZT�V�_����1o���y"*�L|����"[ښ9(��Ɨ�y�$��E&�Q�M�X�:�k@$��y"��><�(
� EP�:�#@���ybH�_�����
P�5XW���y�,�dIb�ϔ��-
��yRJ؝@T�A��Bvѐ���y2lX�"�@��I��f��!���yR��e $����,L��<��*���y"�S�H����Q�8A�ȝ����y��S�,�u"�̆d�,��q`��yB%��K�8��D�Gd\50!J[2�y2���'��{��b��S��p��'Z���"-�PӃ(� �q��'~*q�䅆2D)p�l�,:|)�'���&�%��H�ˌ�_r��'s:�('��Iy�-B7��X����'�`zE��,e��#e��?��Ek�'|4ĪF G�*����82` ��'�`z�#�.^�u�_k<�
�'�I1(C	/��PG��jYx��
�'�X�KF!ڨjs%���K�
� �'-��qe�V*y�(H�c��%
�'brD��@�TD�@�a�b�Q�	�'��\)�
 E~��h0��|?vS�'��h�E�u^��kǊܷ'�8���'h���g#�b��A�'���b���'�L�K"�[�_���cb�� 9�4�
�'pRi�ξQ@���,AO��r
�'v\�ӧݒ>�t� ���62�D�
�'�0"�D�I�"#�O��c����
�'ɰ��ʃ���ذt�\*ad����''l�ȧ얇�
m
�I*�M�ʓHx��銿bX�p����\J��ȓb��mz�fM�AZ� Htg>i���ȓ36�r2��/&�H���N4@I�ȓ\[�h�u�9/���%hL���e��n��a� D�JQ|EႨӽ��Ćȓz+\��uB0L��1��=_:0���S�? ~�:d�"Z;�D	����5��"O,�IM$\0ƵAc�D���õ"O�Ԋ��X1�H:���3'����"O5�3*�p����t��9n�t=xA"O(*�@DL�6KTh�7I����"O0	-ܘ+�n�ѦF�'�,e�Q"O��C��?�(��`�8kh�9I"O�$aRXb�����o��rU"O*��ة5@�<����"s�4�V"O� !�D�l�����ͣadP�!�"O�H��ύA�]�D�5%7���Q"O���aR�0�0)@mոm%��c"O�M�7�Y	W����T�~,��"O\袇��.Wp&tIċ��a���b�"O���fA�pҼI�v�ծV���Z�"O�D�J��N�0�ʕ�J�8�xrb"O�H0�Q"-l��򭎳-�ܡ��"O�D���֟8|آ@�WK��ܐ"O�ݘf��"Z���o�� �u	'"O�`2%k�^x��%���T��"O��)ӊ�S�'pz ��"OD�(u�h�1+�^�(Z�7"O@��r�
8�������N�9��"O��	��ʴPoV�ӄ-A>+��"O�t��G�|@�$c�E �)
�"O�R� �Zܜ\��c,~��T"O���(�?c���_ ���!q"O:,DɃ8x:�z�k٭�p)��"O�k ���3�"��'�Ǒ{���1"O�� `OC�Tu �o�~�hb�"O�HS���\j�J��W�w��A"O����GٹZ��4��%�`�ja"O��*Z$�b,����G�f���"O��b��ǜ� �<O�x=��"O��������;�D�����e"O*�7��*$�@��nE�'�sb"O����O9G�:9s��1��k�"O*$00��1Th\��l6:E^eȇ"O|@5 y LQ0�I�A �Q��"O�@���oi&��P�T�F���"O�I�v��"f�����N���S�O���ȉl	�!R�f��`/f	����&�!�Ē�"#��*�'N?��1��F!�DX�[���`���	��W��?h>!�>w��P"��A�Fh}{6ꊶ6>!�d�@ ���g�ι_��� �
,o=!�DD�|�L��p�>��e��g�[.!�$β7�!�@���\c`u��2�1O��=�|��&G��c�	.G��d�$�]�<�C@�od�4�1"�{�jQzƠs�<���,��X�&��'3����Er�<i��Ε_ ��ig̝��B5
�b�g�<!%	��\n0�h�D��Y�fe�<���!k~�1R6��zF���c.e�<i���d�� B&]�H���:�n�V�<a!��#!�2����;D������T�<a5��I%z��5(ӳJy��1��l�<�4o]�$�r�b�wMf!bS�Fi�<فDq)��aF��0�d��@�<i0 ��FL�+e��0n��(�'@R�<a�*�-x�j`�p�+9������\t�<�e�P�S�`���ADP��%�p�<�'��>����, db:� 6��o�<9���$�R-��Pm�����"�m�<� �܉��͍a��}x�_�F��]4"O�u����/S5�D�$S�x��"O�1
`M�ga���@�)l�H)c�"O��P�Z��x�r �9w�hx�"O,�H�OQ�P!����F�A+��y��7lxL,8���V>�i���ڠ���U���OF
t�m��B���ȅ&I>yl
��'j	 �j� PHqT�
`��Q��'Cz�L�22:�BAA�-�����'��bˁ��,�#�o�4��5�
�'����"�T�4L[��; d��'���c�%�\��ؙ�Y�,�ȚL<i�'�ў�'!A�]�gJ,�<ȡV�\�SlY�ȓ L�Y:������3	z��ȓ;~��E��S�iaKCA��Ї�0!�"�Ý?���衧�I%F ��h�x���(ܡ]P^� q�\;Xr�Ň�q �Ȑ��@�R!B���}Q��ȓlE0�k�R|�9�mѳL�IDxb�'��Hi���3@��-��N���i�'6�����P����J;�Z|*�'	��P��F�v����3_߸q	�'���e���QEBC2g�H��	�'O�|A�F��B�VM����&���k�'3�l�uf�+L�Ҙ9t�P�R��9��'O�Zea(o�L�scV<K��|��'���X�ɇ�| $����=Y�Z�'�xJ KӒ07�J�B�V��\��'�B%�����+�懊S ��'},E��gS&�\a�A#�X�-
�'���!l��VxYq�[�{� 
�'��=R�b�������q�ȹQ
�'�r��(�06Ds��øm�
�'K������C�
��#[ވir�'��P��(�
>��!��I��\�
�'��@�e|���q��$;f@tx
�'NT})S�8Z��W��𶬄�; Ĭ���$4rtA��S�dmf��ȓZ/�)z�Ԫ+
���� �|<�ȓE�a�C��0~~l�bDQ�L����CB|X1�M��
�L`�ڋ.���ȓ����l��<hC&

_����f`��5�H6+���b,�c�
��ȓb�f))ѱ�aW':Yi҅qqD�f�<�����6��rD�1=	�ѢϚc�<u���H�z9S�&1Q�.�p#��`�<Y`F�O��`)�G[�'!��%U�<A4 �f����̒+sN�l�F� S�<)�L��1�D�+Y��Q�5I�M�<���.eNN�
FEռO���)hF�<���n��ES�E!uSd�IҢ�~�<�����T�@]�2�@SX�,�Q�<Y���RƘīݝG�M���x�<��&,;��i��K!Te$���}�<�j]�A<��� �p�7��C�<A��|+n��⓲C���"�Z�<����kPRô��+b�4d����m�<qQ%�*]�s#��k�ӱ��d�<�h��9���Is�8!bJ	��y�<9R��g{Lɘ�K�4#��|�mQ]�<�W��oRR�z�fγ�>R�Mr�<Q�P	ZfjH�3*md���c�r�<��C#���EDޫ&�E���v�<�F�L��\넯�-�>�)�`VG�<� ��J��-�F�1�� AkR�h&"OTh;�4�y���8��5�"O��K�Fǭf|2�Hb��&��h��"O�z0ʩY	�ِ���6~�B%��"O�h��%Ŧ�J�#J�fx	3"O���h@ ��t��
�O�2�"O�I�%j͜N<�aÑE2ba+6"Oh`��������pXV��$"O��d��\�FRИx�L-�"O�4R`
��DE3Q!H�&��SW"OH��ۺ+��(�F�n�����"O�q�PiJ�0v���@�ǩ�2�34"O�s'��/O�ez"�#d���z�"OZ��ƻ\,���W��V���ȶ"O�!����n�������a-h�q%"O4�s��29�"h���.(���V"O��+�A_�0����r�P&`)ĬP�"O6Q��-�k� ��PAU����%"O>T!G��<x���ϝ?[�P��"O6��"8j��C.��LM�\��"OH0�0�Ř��,�nv��R"OV,�t�ωw�)����R�*�@"O�]3VBZ<h����P��0��"OD@{5�EV̱�hY_���"O���fH��;Q$�@c%��W�h``"O������ie��8 b}�:Y�B"OTzrā�^W������>Mc $"O�=�b�։S�\�2o�bH��P�"OXY�"��EH�"D�4v<�"O2������^8��!�T2�p"O��Q/�6p
�i4�K9#p\��"O��4��zG��kD�d�8U"O��{_���4��D���@4ď��yr@K)�\�c̄S��!D�D�<!$���E
��:�h
#�\T���Tv�<����:�����]Khx�A�g�<i��U���C��,؃��c�<A"�� pht��۩����g�Ib�<�c�� [���
���%>�0T�@[�<!R�a�Υ~�b�zA)�Z��I�ȓ2�͑Sd��Ű��B#�<����*		�b�P�hA��h�*F�����n�I%�G��^���M�b����i0�����Y�i L�Emo��� ����!e�L~��c0��Z�͇���ъׂ�1Jm:mۅJGh,��<�.�ç�Z,q(�(��C�+�>��ȓ$�Cƪ]?|�p�� jyP��ȓ��X�ˌ��@|�1甤H$�=�ȓ_� R���wCP4��钥�i�<9%�O
\�A`cX:S_��q
�^�<�V��1?!q�k]�;���R�<i�dƱ�
�����Y�Ȓ@(�P�<�a�^�T����XV^��X��_A�<�윪.- A�t�ș���P���@�<�&L�c�¡�a(�5�����^}�<�b͈HA��b�� x���M�<YF��G�F��A�޴"�0�d�e�<�'+��i����MQ�����b�<���̉K�"��S8.��ynz�<i�� yWT��&�R27<���_�<��Ȟ$Xn��&ݣ�.qa@^�<��Bu[�yBT��Mn���r�<qi�|O��1C"qrX8��NE�<� ,����\$��(=Hbb��"On�k㨎�1`B��D4"qڅR "O���c 
�n��i�'Yb\�X%"O�`��Q������/E/\j"O�@{���#cQ��"��S�}��ik"O����*�"��������M�T�Z""O���@�ZH�ͪ`�nJ~5ȃ"ODL���� ��iX���RZ���"O�,��*J�<�d�iӧ�+@�y�&"O�@�FKM8z��M!X�+,
��"O�haŤ�wV��(t�)l� "O��y�MHF� c �7�"�H"O00���4���c􅂅0��G"Ot�c�.S/H�]J�$_�Y��)��"O�U�kG�L�t��\���	6"O(<�&�<'c�c`� �E���1v"O\$j�E3|UT�s��$j�	3�"O�14%�.R[��Pv�9@g�Ŋ�"OR�2��E6!���'��#��%�"O�� �Q��4K5� Aj� Є"On�����:������2
��	C"OTU�a�ؔ^�`m�@i�=2|z�qe"O:�xp,p��ͪ@ϡhg���u"O!Cc�2Q�T�C�GG�bx���A"O
X(%C>�.���F#��e"O,)��ߴIm��hׅF(�4x�"O$�`��S��~�(��H�D��p� "O6)�ciN��>9p�I��^v�$"O�4���ߍO4|h�IQ l����"OP�)w+_8��H���P
���'"On0��숚
�PlSFaRE�|:�"O8��6��!{%�� ��^�d���e"Ox��⣛��}+�OT�9���["O��D�
���T1�yͬe@C"OV9rFc�hPJ(�	U�z�4p�"O�DS6�/9�FY��Ew��	�"Or���h� ���QE�M(�+�"O	��eǕ3��Y"��z�>��u"OZ�P�&����qE����@q6"O`P�G[0Ye.����-	�� �"O�I�Cl��iiCI�?J�
"O�=����Cu
��'�
2�D�[�"Ox� �$Y�>nV��AΤ9[̬9�"O��Xs�يc
�ҎKA� zS"O ��E��g�zY#E��#!��� �"O��ҷ��!2��j�C˓ �r���"O������+w�*�	����m萹�Q"Oj̐��Ă[ ���.N���J�"O��R㫛�-��y)𩟛��m��"O������x�Tu��i��L��U"O|Q0�@^5l�rLQ�&�l�,Q�"O��9'�<E �)1f�s���Z�"O�5���*M�X�NO�W���ʃ"O8�z&���n�D��
'b^�QV"O�t��!�y��� 9|��0"O$�#uo�;(V@��ǉ*���"OT�Z�aݵRN���ک4�N�"Oz�g�ġe�0����Q�E���p�"Of�q!���^&�!��Gդ���"O�9�K�6-��| �/���Х"O�I��Q�L�b �ud� ��V"O��H��Ж d�J刃�B��Y��"O����A��4���ӡլ3�"�P�"O��#P�P4d�RuI@Ý|İ�s%"O� �h�h��p�-�o��l�x��"O���4�� bR��I|1���"Ody�'a��Q�h1S�(�	|���"OH�r�J�<;4��a�&�2Y����w"O�B�I�[�ʑ��%����C#"O��J�?e�"U�5$P(/�б�A"O���E��N�+���-&DՓ�"O8�Ê��_�Q���9,l��"O*$A��W�Yz�H�� �tJibU"O�x:��lF�z�΢�f�0�"O<E��( ��v8K��^7&�NHX`"O�!� �T�j���E�ܰez��JT"O��(Č_7H6�H�R��}\,�U"O<!)��S>���� �zDnժ�"O.cU� F����a(��(E"O�1SG��`J��1@�1<�����"O��J��
���ȚE"O`$ځ��LhQ	F�>|�e"O�1a���(@�.��цR?J� �!"O��֎)��S��>��E��"Ox�� 55c���1+G(��1"O6�ٵL�"��Iru(7B���'"Ov V(�
����H�'sm��bd"O��� a�f��q��#aj��A"O��R�hI�,�7��jH����"OTh� ��[XJ���&��}�LY	�"Of4*�ßKu"��$D��!�ڱ"O~�
%+_��y����>�J4�u"O���/U%K�P$h�a�
DӘh3a"O�@Pp�G�F�<\P�a�1#%���b"O����؟p�~	� K$����"O.T���_�3��9�#oW2oДYE"O��Dj�gG�Y���'#axM�"Oԍ M�^�1Pw��-np�|K�"O��q�+�[c�mc$L؎	>iD"O��*Ε�߮\
pMϠD.^�"O�xJ��W4b��!�Q#t,t��"O*PC�NG7EO�$0�*��v,"O�e��B�$#��p�JZe�<)�"O��0@-6�0�S��cE����"Oʙz�y3Z��b,�/+䦝�d"O�8�pC���`	�kI�m@��e"O�(�w�69$k�?R|d�"O����/ ����)͏�@(��"OV���M�p�E.�{��b"O���hT0�j�Ö��(E֮QC�"O&���ץi�D����I�J����"O��j#^(*�0S��l����u"O\؂��\$2>��"äR�?]�9"O���ȊnW�P0S��4�:���"O�1%��75IPF����q�<���3&
����,9���W,X�<��£*A��x�ɗ'~��d��`�W�<�O��rBVHb3�ߟe��T6�i�<��'<�Θ�"�X�41�©�g�<�s�0[�"��wE�R�|�����d�<y�D�z��9"���&kt-��+�`�<��:JĈ�q �����#c\�'�?���D&w�tۥ̠#����!�>D���@&Mx뢱��^{{�`j�=D��:6��{4萃!_�L����'�<D���W	IFH�� ��ȋ ܄e��'D��w�׼r�6� ®�0p(�3�$D��aìZ,Ľ� ��o/�$p�.D�� |�RႥ<��ա�停}o�\�5"O4��_�SnN �dE��yV ��C"O|��'�i�` ��jB%m:xa*W�'4�ɮ����Ǐ	�i4Ր&���w��C�I!h�*�z�IH�N�2iy��A�\O�C�I�o���¨���*��@�B�o�pC�I)O�� � �8^l�D��@���B�ɘa�(�s�V�2�\h≞� ��C�I�&R����\�[~�� p��"�C�I1� �C�i�+X�����Y��B��>��@����0���o��9(B��44�H���9<6��W��5"V"O����Nì,D:![P�æk���"O��1gI�+H �����r�A'"O�x�O��~���!e(�:D�����"O4�pd��{T��2�f=�~��d"O�h�aI���sU�������"O���5,ӏ@ɖ�p��Rb���"O�p�f M���8�j�  ���u"O蔹⇃�#u��O]5TK���"O0C�n�1Xxj��w P!H;L�(�"Oi1�D܊=U���w�X,Q,���IF�OҌ�Q$��?BF4�m�% `"	�'�(ە���¸�c!�hܻ�'�����*ʘ#��� s�(|�`I1�'% �`#S�q��<y�`֔xb����'V����],1:����X:T�y	�'�d�3"k�0Hox�� L��(��P�'A!���?5U��i��u ��b��d=�'Db��*W�pu�����3T꼰�����1���9_+�a8rAY*~�U��p����9:���ч����q�	V�����(�eFS }��8��C�[N>	��9D�DcgH�~a�E� �EN!Rf�8D��i,\��)֦xܠ����4D�l���]� ��U�6��yZ��1D���U7E2��p+\>H\9�Cf5�6�O������\C ��{��!�c"O���b�'�<Ȫ� "c� �:W"OF�􂄸Y��2U&�u��@�"O�!Ə�C���b;���iR�'c1O9��6�&Ac�"��VqX"O���s�Ȏu'Ĉh�c%Zd������D�O�TM�2��	��I�F݃*�r��	�'.jlA�I7j����#�J	�'�jكRK�m<������*�JP�'��T a�[�[��Qo��Qk�'�J��u�N�E�}��o>7�L+�'~%+�
�x��ɒk�A����'e�3W	-j�b�+r%��|�����'�,JA����;э�,z)�p��'�X`Qӈ�?m7����qi��
���y�s� Y���C
�����y����Ip1'L�J��KN��y2�+.
� �$k}�@@B$��>y���y©\3�|��1�n�F��6@���y����ݣr��4b$��Y��;�y2�J3uQ�cV@F�h�(\Z�G��?ɍ���/?��K &����H[/2�ډ��#�N�<���\����5��/�^�	tiIΟ�%�\�����IR���Wm��r���f�޻F
C�I�B"zl�Ģ}@�|��	�X2�B�	�wAsd
�$m����Ř�*%�����OB�$c���B�R�l_�y�p�Y��`��6+-D�� @�0���Q��:�CS�ju��"O���l�I؄�s�
ƫ���"Orl	`)̂L�*p{��[&�b�w"O����C�#V�%����
;����"O��aH� ��ň�0'VDx@"OX�B�9�J�x(��cZ�bS��'�	zy�5O|X��aZ��ܙjQ..=��"OT�!'ꈦ$��� g/V��vO:գ��]�:i� �L8� 0a�l�O|�`D��'i6q!@L�1��<�"ʓ�u(0�����?q�B�I�L�����"L��S��/0� B�I�\5��l�8F���9�-�
.��C䉽|���:!�Kc��0��#Mϴ˓��O"�D�On�	�Q�������PnԡI1�^�@�vC�I�&�jE��|��a���:�OУ=��y�cL>>���ʌk�Bq�NS/�yb�C;3�`�yGA�.^����L���y�N�&"TQ��䕇iZe�C���yb����a7�v9�4���.�y�S�H+�h G,�%@��j�$� �yR P�KL$P02�����D���y���4RX\A�� �T�Ð�	���4�O�B�鎅/���8"�ӈr�"��#"O�E2a �5'�&݂�M� @��['�'.ў"~2 ��?��!�fSQ�̐�)ƫ�y,�>}��x@�X%P&��h%i:��=y�y��+]����VK�!>olL����y�W��\ ���4q��{F�֢�yr@�72,0P�4-���2fP�y��I�4�\1�;2���S�D7�y"�]�@<3����!1��<�y�<=��L�!8�(])�J2�y�I��r0Q��C=&c&�+�C��y"���;"\Pcc��h�0F.�y2I��`!z��N;ž�P�ԁ�yI�!uNd�Z⁜���;��ɝ��O�#~�BhG��X�����lj��ۘFU�$:��?)�𤃁o#�t�DI�9��8��*j!򄙽\Z)⤨Z)+xE�w��o!�K�adtD%�٪}&&D����6I!��O�M�2d���I�9��Dk��ȃma�'�ўb>a2��2A�l�v	B�e �H[�X�<W#	�Qp��pP����<S� o�<W-w9 �!��э3��=x���b�<�b
��CZ�1��=�Ntqn�ܟh$����1W��e�0V�F �$O�egtB��+O�Lف��F5(�b��:g��=�	çHV��i�,�Ra����mh\�'�	F����`��;��� ^ Ta�M>D��B� L��dC&!-�>I�Fd<|O�b���U���q�|'��-$8�r$j8D���H��K�x$�g���/YD�`#D��BNJ�^Ց���.���B�"D��:���J1�l�S��3d�-���#D��!䇿h�н5��i��� =��0|�!�:d�h�{@,��y�i�l�<٤a�"o��<��5:b�p3��TA�<��T~S�(��N�8Ȉ��P@�<I���#G~�W����p�y�<�V�B�M��Cd�u<�nޏ�y͏�`Hd�rK�.~AZ6Ĝ3��<����-aI,��0`ʭ@h��a ,�g�џ E{��ُ �;�.�9h�EB�(\/5�!�ę�~昹+���z����ǔp��I�,�?E�� >%���=�\8��2��D��|b�)�-�d3�cPvL�5r�闰O4C�	��q���	�x�`����vgnB�*#pdS�
%J(2�YÄ��M�>��;��90��r�%���y%�ѯedC�	�q~rU��a]�S���EaJ�.C��>Am����׽˴4ȥM�'	�*C�'8�9��5���bA��.E�2B�I(f�E�̐�M������&:<��=�ÓxӼ�Ґ%�a�@hW[
Y/���r֩q&�͔Y��#נR�ȓ!��*�xt�=x�n�("q�e�'g��f�)�Ou��L��:"�,S��ئ[��X�D"Or��O�+Q�}*�D�,�E�"O�gk� k�t%R��]���z�y��'�M� �K�T��GMl��a�'�0�Y����_KbHR�hŶuP\K�'t)�@ʴ]�4a��a�@�`4��'���X	�Z���6S�P8,����������s"�D;	M.��
�E�Uǁ8{"�[�
�9u9��ȓ!�\(@W��En�J��̎O�F��������u������R�4���6��D	�̀P�(q�3�
2�����̮i��:D��-�1ʟ�3���ȓO7�Փ1�L�@��q��4H����E2�Y1�C�&#�}���O�����!H@�؀X�V���aB�����<I���=n~P2&#�h�C⏗N�<���]�;���CQ�X6F}���J�<a��X#%�$,ip� #7"�|[�mGI�<a�̍r ���!
�G�AC�WN�������$�(Ru�A#�0��Ts�H�:Bj��ȓMfe�ϵ?��x3�e�6K��`��QM��1���uFPY���
X����Iq�`r�4r���8u<�i2��S��8�ȓ"����g�?&6f`��Ϗ6�$�ȓ+�,�:FL�j�Z`�V �B���sO��7d؛��X!�i�r&��ȓs �xKT
Ě/ژG+=F���	c�xy��L�$��#�X���ȉ��!j�.9D�\ɥ ߞ?�4Qj��!:�n�{�/)D����m��j�(�C���t�x%�)D�XDƿY��
7B<rN�0��)D��2f�ĥ�qI_eb`���(D��{v
�hR����[#�� 0d:|O\�$�O@��@Ш5S�/�E��}+���C䉨?^x��D��du��M�a�vC�	wZybg��J�R	�0J�\E�C�	�	V�x�W#äa{�`�n�>��C�	���qS!W�O$��x��M.�C�ɗw�DQ�H/����E@�IڰC�ɏ ��)z@���8q��*��C䉵dw���@*�E���bD��;0O����1mbY�U�4�d|��W�HP&��.� �
a卧=�� [�n��x��ȓ`v�qʔ�ПD���ߑ,Xm��"Ob4���U�-�$��A�Q�dh$�80"O$�aQMW.<�|4z��[&T�06"OƬKf)#7.$����1<#R���"O��[���5�~��b��.ܬ��OLѐS/��#�A�A��%�<4�V`1D�p�.�]h�� ��¿6}
,Ȑ/D�4�!���F\eA��D� ��g$7D�� 6�*7I�;ϖ�ǋF�.p�Y�"O�`�f����:4-*j�B�"O�Y��R,5V$L	���.G��$B0"ON�����_�����dǉg����1�S��@�j��K�ǡGE�U	R���!�d�=i@���M�E;�e��^�4�!�dX'C�tQ�њ-v(3�(M-!�$��y:��9��f1���U.F�Q"!�$�#'��I3�E�v+6II���@7!�Ğb��hr�٢a��k�\K1!��&A��͈t$�%UQD��:�џ�F�ĭ�/p�(�ե͂x�P��֒�y�.\�,�Y�q#*e��NW��y�Ü�(�*,�1AUo�����O՟�y�*ū:�6�P�Ռg��QP��]��y�9#��f鍐r��M2��6S/!�d�*�ڶA;[�l���Q�P/!���0�������&q�h�"�噻((��)�n�4i��BߩT�̉��4�*	�'��t8��?Ul �{�K�4"�k�'��SjA#N��E!�iL"�.�X�'����cKO2����3�E��'���a��U�z��RB�2^�1@�'�^�g*��?��`KO�/1V:���'!�e�P�Є~�^E���;+�HA��'�$l)`�Ƙm�H�c�F�@��'���	�mB'?Pp�3�L/0��P�'��D+� 0G�40�M��|���'�~`0�>���S�h�-��<�'(�I�D�K3V\\�Y���xj24�
�'���� J "��d�J#x�J�����h�<P��)�+�N�\�suo�i�<��$N?'@q"���4���"O��c��\�#}�M�!�O&.<ȣ"ORTa�B�0#�u��0� �V"O�B��ƚYX��R�nŏ{�Rɉ�"OҰ2��p�|���L*k���j�"Ot$����c'�}H���3�2�0"O�)c���W�L3K���P"Oj ���0M�\�æa�<Q�"O���
92�jQГԜ+�z��E"O�Ɉ���
K}~�qďR�e�.��F"OVS���])d�YEn e���*�"O��@u��Cڄ��G� �v��1"OP�a������t�f¢\��"OL�E�:��hc��=���"O���C̑=�T���ܹO��\�"OHy�'�P�le�ir��ȞE���`"O6	X�,��1 Af@+zz��#�"Obу���I�����	
Svp�"O����H�p��A�s�Q�WȒ�"Ot�bJ^�,�d�[��R ��X�s"O>IR��B�ȃ���7�h��b�'����"�kõ/bJ�i��j��B䉝��U�a@�a��hi'�W
��C䉄KaJ\��i[0DE�����
#&�C䉁M�%�cE�6���+C*��NB�I�|�����]�h0�4$Ԧ`�C��<k�zŨ��5VQ�&ж:��C�	 �*��冩-��ı����	�B�	>HNT��!j���ҕ��8�B�	�$�� �N1q��8�0b�(Q��B䉸�Ь��@�8Ǝ4 �"��B�I��U��˕#�|<�%��5�B�)� ѹ��(dpЀ7)Y��3 "OH�����pt�1�H�J���"O�x��K *�=���@8&�T���|��'�pd�6��_�z����=b����'pHW�U�Ԩ�#�B:F솰��'*�!3`�X%MTLH��-<M�`��'���`�9�i"��Η-t�a2�'�ly����*����/�Y� �!
�'�HIxd됫%�T��#�Q��8H	�'�t��"ρ�56.<�5* 'Y�D���'���T��TĠj5%� ��1�'<�9�F���?����	�/��`Q�'LB�����F,Bi#r��2O2�)�'�HX�Q�Zd(8C�	ՊN�|	A�'�����0cL���S�Ȧ4r�'r���5@U�_��B��Gb�X�'�͚��F�7�\�Hp�߭L4JQ����?O�����a�z��A)\�!{�l�T"Oa�ԩ�xP��x�E�<Hi�3d"O~q��iW0��-�ŀ�egf�B%"O�Y`'G֟K�Lt��O�c��0"O&��E�ʞFv�P�Ta�(g9Z��@"O�LzÁ(8 88VA "s� �"O �8�`��<�V�Ǻ��
k����O�=��'7�PÆ��o�h������H�.�0H>y�'m~����� �� S�u���ȓ]xf��c�x&�)d��'
��ȓB����G�k�f��Y*J\�X�ȓ;L��C�)=��Z7A(&����c���C�	]A�Ց� ؤ�^���z$m�Q@,J`�=�!��\T��SL�eh�+]�Y9�	6j���b͆�E�Ⱥ�/Wӂ� d�Opj�ȓ2.�p�g���M�0@��S�8���`ߢp�E�0�`�{��E7�"�ȓz7��ɣI
"xS )���U0p�N5�ȓD��T�DG�jK�5rP�_+Qn�`�� ��᩵��(1I�����.�݅ȓ}v@�T�K�`���ɐ�Ǽ5�ȓ�B��㣎��q�kF�����ȓYH��

�X�� @�����ȓ~cVIp�H�a��(�1|����=@��Q��T4%,5��a��nՆd���|iI�W��h�!��MԄB�I9�t�H�&µ-�4`�@Y8�B�I�O�&1��]�5l�(����E��B䉺�R�b��Or�;�l��
4�B�ɮQ�|��+Q�v:�� f�N|B䉪iZ0��q(ͶiJ�!*��c�B䉫�81���'[n�`b��>)rB�	�A;�����E�I�V���B�Z�tB�I�HQ��Z��X����w��-y�B�I6�3���c��) ���"VF�B�I.jz=&DI�r�!A�Ř�,pB�	�
�\���ȓb(�!�2`�79JB䉙s�H�v�G�Cʊ-�V+v�8B�I4Q�P�GX��}R1Z�<}NC䉞�Č`o	\T]Z!S�m�BC�I
8�Դ���N�F}1G��?f��C�ɪr�T����!>�S�j9i���d)�
 ��%�F=����w,��Q�Du�ȓ��8qD� �P���֔P�֩�ȓN[8�����Cz�Ѫ��E,����49NDb��>��'�Hv6��S�? B�1tmZ��"`���4FJ��"O �{aӡIX�葮ǧT�6e""OJ4B�(�̽#d��[���"O�l��K�)'~�8L�d�Tx8"O<�w�Y#9��4��̢5�ִ)�"O(�؄a��$�$�����"O����+c���i) 5"���"OLd�e�>���8բäQ&q�4"OR5��!*��QLE/?���"O���#���[�P-�˝�y@���"O�9�@��9�,�����#'�=�"O�Q��:h�d (�*Y,ò���"O �!f㋂
0��5�Z�a��4�r"O$`R�4d��y#��:�(��"O�s���88r�XJ�@Ʊ9�d���"O��P��@+ ��ؙC���6l)`�"O���Ʌ�/�V��XN�t"Ojp�LR鼘8UN��fr���Oh��6���Qb�ڟ8����n!D���Tb�$w3���w�َo��� �1D��6G�6s_�Z�ח�`e�gK1D��pwk�5Y��	��$G�T=� 3D��p"�6!D�#�=l}�|`�&D��z�n`����b.eҨ�L$D���2�܅0�|U���%-�� �<D���G��-�P�w��y���;D�,�v� �`�d��sA�9[�8D��*�(B�gTi�&�N� ���puE6D�<
�k����Rڎ,�����.D��9�*ùQ���2BW PL��ڕ
.D�8�0fO�uM|����<k��:�&D��jd�	X7�X�� �:֌7D�D�s*G�g��8R /�N�H%-4D�L��L��:}�E�q�01;d�3D� !4 U;�A6���h����7�.D�h{���0jr�c�^�+d@���N8D�@4�XU� $��D.�$���7D��R&c�'Nl1Wb��gf
���� D���A�"r�Aa�
���b�?D��[��(j���I]�k���w�;D���BĄ<b\�A�G(pċQ%$D� ����7~"��tlJj\\!��!D��B�΀�w�����l_�\0HG� D�h	4ퟹe�b(���9r��8E#>D��2��E�P�"�F��:3��ջe�&D�lZ�AζaR�I���*�LA�w##D�����<V~@(r�tQ���T�"D�Dy`�X�4��Q	ûy���O"D�@����Pv�-A,�T�4ۢn?D�<aRZ6]l�3�Dv9��C�=D���� �(|��yW���>*d��K<D����̕����.���[��:@"Ojd���9t���x�0%�1"O^m9g��,��G�S�Y�r��"Oƍ��@�o�V@yċ�.7��"O���$	"V�H�d����9�!"OL�cԋP��6HK��[�3p����"O���؄~�<��#�/mJ��1"O��j6c�/+Z�(%L]5Ei�"O��V�!�Y��� k.��"O++;�n�Yg�K,�(���!�O�<Q�.�'Q��.pd��Q��K�<Q7�U�$�%��u$K�`�`�<rŏ�6+N3����/�$�rc�CQ�<� �}G&mY�
�d�..�X�;�"O�kcd��'1����[%_�J���"OF�s5�]�w����JN��NMI�"O��K��^��ex��!n|��7"O��A@F�S�N�;P�ë���7"O���WfU r&b�餤_�����?!�$
3���cZ�U��1��%W� !�$�f��4��Fh���re�&!���>0�ĂY%}��	�Q%LV!�,CT�17��l|�ӵ�APA!��<`D��r �ŔR�� J�=!�$H�>��I��H:=NxIC!�d��_ 08�b�m\� )� ��W-!�d�rZia3+Z kL�|'�>{"!�$B3@��Ԅ�^2v����@% !�����q�Hx-��
"�%f!�2_iH"W-�#i'J��0��;!�!�D�&*�u�a��:�Mr� �?!�$�X&��b�F����@@��
�'�\iCd�2GL�U)U%d�84r�'�P�a�X�z�(����cg�%��'��:1H�"}��J���/V�!��'�6��S�γ|'Vmu�=`�f�[�'����p˨,�܂��ݼ[sPh��'�6�aO�S���(DAѭMn0���'��ek��μs���83#�\b*��'e��6�ѽ�(�a3)�	[	<ER�'|�� ��]����b�]���m��'r3�C��Jp|��"�\8z$��'���%�0>L���Ӑ5�FH��'����LΆ6�^�H���<!P}Y�'������5���ɵc �c3��S�'��P  %��i�$��t,8Zq����'V�)��-L*��=��(S��셲�'8��jG�Z�22�BC�3�0e��'�����J�'jR9��`G$};� `�'Z�e2���4q|��w@�:{UT$[�'�T�WI�AcȠ�/C�D�0�
�'���fiāѮݰ�'X'<IB%��'�&x��J�y�8("���=~��<S�'�p�Ef����YV�Y�'��(D�@�?H��@��L0F
��'�`٤mËt?|�mZ?/��j�'�*�ku�"7��]k�AG,�p�Z�'��Ȑ�&Y�Y��d*%��"�n���'�h�k(��XA,�Aq�:%Z��'i��[�JE9r^>���)(vt��	�'۞9!SbE�@���8W���D9��'�6 ( ���8`��ږ��.����'�,��`�K+&�����̄[�'��yq�S�c��!����v�xA!�'�$@�D#*��-�Emχ!�Y"�'`i������z�+	��P��'��� � O,#���[DL8k��@�'?��(�k��Q����ۼ��%C	�'��D�aڊFkR�	����J�'ö͠���?��s�.\�d�̹
�'A@M�s
J`Y�4hU�i��'�0QO�,q��q�G��|���'�,�Pe�ЇTLp���*��#
�'����2e�(y���S�#�::
�'od5�"��q�<]sv�!�z���'G$|{ҡL1��������	��'ނ0���ߕ��} E.�_��8X��� Xm��aK����B�͐9��U�a"O�;b�5�L��f�J�+��1"Oj����W�.1�&��-ZT)�"O��H�b��]$:��C�\�OXQ�"O�eQg��F�qU��/nE��#"O��P�� ��X���&b �q�"O Mj�e��Q��3��/W�٫�"O���Q��<s�`��Ng�ճp"O$D�!*����3��>#[�̐b"O�bPf+H<��kB+S�,X �"O"�W�u�����@�A���6"OLu����$j�LG��0*q�2"O(�����)2��Gһ>�8�"O~�Ѥ��H�Nq �o��w� �"O��D�bɓ5⌽E��M��ᖇ�ybǟS��W!?e���1�y�j	$�f@8��X�	ɂi!p,]1�y2	�\X��K���t[��0�y"�>q>�y�f�O 5æ���yR��V�jIƍ
���P!
6�y�� �3��t��C�	�4(�0��"�yrAX5$�|Z�(�9r�<]A��ޙ�yR�ҵQ�p�i���qӀ)+T(Z��y�3Ղ`��ąb�����cP�y"�*d���oɗ]�.�C��9�y�+�r�������<V�ms2eՍ�y�&E�b��೗^�L�ʍ��6�y��:Z��$@���>'R�Z���y�G��x���+b[PQ�Gj^��yb玠V�2K �6S��\h�N��y̉�v��D���]G���r��V2�y�/1_�թ�f@4o�T)�� <�yr$�0Q�N����]�8�1�L�yR�V�^�"͊@��X@���j��y�C��)?<�+���5r�qC���y�+`V%{��yr��:����yro�(@���ʄ?x�����7�y��[6!>�×eUiwZt���"�yB�ǘVJx����"sØ��*���ybcp�)��͓�3X��fQ%�y&��W�h-�f�̜9���j�IT��y����	�\�s�&@�8k��zc@�yr'�L�K�ě�@�J]��f���y2�V�)��ʊ,�\�����y⤚5x��J�:ˌ�����yR�M�-uсg�ɝt���P����y��W?Knn�A����lF�ْ�-�y�N׬>8�%�ռR,�d9&NN��y"���D�X�4I�U�pQ����yB
�"���B3fW�Д!&Û�ybǉ�?��`)բ�=x�x!�h��yҥAv1���?�`)4д�y�'�#)�������R�(P�U]���e%<II�,]�	[t�'f[�O1�T��_��8 �'�#8*x����H"��q�������X�hM��@�HӼl,��e�B	�!���d~0{ҍ$f�]�ȓ7p��s�	!��pk�Du�XQD"O|EY�N��zNr��
��܏	!�D�"C�!�"��R:��r�C�:!�X�
՘T��	H!s��i����J�!�dJ@�(�q萨v�B4�צ��c�!��	�/2�`K�Dq
�I"&]Ar!�T�!_ld��o�}2��2$A,QT!�� ����� ��s�ҍ0Z6S5"OV��Gdޞ3�j0��Kɗ$4�tʇ"O�!�S�$D*�lR�@P�kh*�"O.���<:�� �DD���X�"O^t��ŝ<^��3��F��Xf"O�Da��`I�ȴ��5J	�I��"O��X�HʪT�ls$��7>�b�3"O�9 S!���R0d
3�l�"O"U���~�4$���@�
�YT"O���©G�b݈	��:�4=*"O�QwNͯΤ�hj��1��E�'"O\u����{ >̚Ab����(�"OPI�cV,#�>���*>�h""Ox��flڇJ��b���KM�eA"O�tA���n��Y�F�DL�ڦ"O��H��M���'\*��R�"Ob%�T�L8D���+p��@�"O�x�e�%3]�X!i�?xV���"O��"
W�26��j���$��Hf"O:Hk�BO�	��S��Z%!��"O�u2��.�$�C�ׂT'���"O���M�|(����9mb���"OR��5��~��Z���tP���"O��I�DO/��CA�3J�<`8U"O��*F �5�BY��E+Z5"O���?M��t��<H�q�`"O������{3F\@��Z�+ X�c�"O�qr��Q"�e�4LL�X� "O��#B�B�B���$�\��"O�S�	Z�p�)�4>��R�"O��4 ��w�K!E�F�;t"O^}�Ge��<$���eH�H���`q"O6l�Ř�����E���R�0X#A"O2�����S8D"���D!T#�"OD�0���5� �T��D��"OV���>}c����G�PN��w"O,a�"��>*����<
��T��"O �����4�VDx�kS���2P"O~]H& �x��I)�� 
]=T�R"Opx��#ʥhw�bՋ39�H�"O�вPl��%���	�H��F�̕��"OBd��	Y#5xti.��>-�1�"OE�g#=�xu�a0L'��2�"O� ����"�S�n��6��5"O&aj��:���y@��/S��2�"O,�3n��qJ �@L�a���b "Ohy�E�4G�(�AŦF�t5)6"O����@:#)r�	��A�}�V�"O���2��4jZ��%̓�8�@u�"O:)pAI�fl!�#W.��7/�!���U�:�9���4P�)��@O�!�dFv�Jq��i�9w����BNU!�Ӂ��A��[*��baZ=!�q�ve�D^:�����4#�!�Ȅd���Dv�\��k�,�!�ߓ�D����!n��T����e!�
�<���K'�;Ķ�
��@�!�d��|�ơH��[9G�,��6E�S�!�d)uj� qeځ?����#�j�!��	rH�3�R�F�� ��Ș�!�d�T��-�Do�]��c�k�<
�!�Dϙu��H2%^�����J��!��ë��hZ���
�^���h�Y!���r�`9:T �-V��
�J��/�!�� (<��ؘ ]�D��.ضK��]��"O�|��6�H�#]-�^iل"O�Yg����f< @Ȍ(��d"O��#�2~^�Q�H@;����"O�z�a�<P���֞*-��w"Odx[��І*�h�1F��E)�А�"O"���C?Z�B�┾ �`"O=�	�k�J�g��\��:�"OTd��T!Į�E�<yx([�"O�(ʴ])K	4���B�|���"O�Q���X+�,@K��9���"O��*�%�f�!��4Z���&"O�}�G�E�Q}LE��H�scz�;�"O��Qၻ�dh�w(U,G\��Z�"O���c��a˒��$���A��z�"O��{(W�cS Ef@-H.4uB@"OB��1�e?�%{ ��ww�0�"OJ9��$]9$�����ۼN�de9�"O�T&�-[ZTd:v瑱u��LQ�*O68��b#kDh*D+��Tg��	�'���UC�;�^�2"/��E�b	�'¼i�-�3Ġ��π�jZ�5��'�V�b׈�<B0i	'�iE|]A�'�}�5e��]qڑ�-H�-��H3�'PzA��O	0|v��E�
��T8�'��`�f���z2���Są���i��'��U�'��dH�(�wF=�
�'�f�Z�4S)s��~� l��'d8z�� z�La�bJ�"�Бz�'#@pp��"z�&a��!{���
�'���s懖�N-|� ψ-bF���'�X�]��V�xgA8c:���
�'��Ԑ��մ(�J�0�
EM��
�'�j��0C?�z��X==��q��'���cv�D�B��Sc���5YL�2�'����V�Y�w��ibF�3,�u��'�j$���?
3|�
��ߏ#ެm�
�'A�T��Aȝp���Y���(	�'�^|k��;f� ���� ���':�����@I(`9��*��
�'�*�� ���O:�Y�� ��q%��
�'MmaUfN�T���U%	-�T�	�'��Z3�
#(����|ڜ�	�'�����7i���������'9��!�NK�e��4��&Ư|rX��'B�K7	�(z����u!�-�h*�'�����	�H�a���-A�\��'$�h�ݦK�<�a�n���'(����f�2�D�zYH�����y��̫D�R@)4"�-9�@4�U@���y�,��%<&�����=8s|L#o�=�yB+��`�p=�AD�+����t(ܳ�y��η+��k�휉0|�4jG��yČ�7�����'����c�G��yBeh��r�e�\���0#	��y��ǔ7F���AS.Z��#��_��y2%P�?� (�eGY�uYrOI��yB�
-V�ԁ�g�0?FT�iT��y�B�G؜�avL�
OR�\��-�H�<)��-8Z��bD͉LJ%2W��L�<	  B&ˮ�h�Q�m����`!F�<�d�='��a�Y�h�䐩ŌF�<I�g�	`�`� ��M�h�"��E�<�ņAL�xA�ލVGX!���z�<� ]���,)'��&�ț}�����"O�!ö�K(h��sK'X���"OFe��͉e���2��j����S"O��b�(/�AZ�铳7� �*A"OⅪ�W,�d�1#	�	T�F`��"Opj�n&E��|)0.�k�\]
�"O�ȂkټO�>��qk_^���{�"O�ᩱ�Ą3��uː*�o�=�!"O�H�U�K"A>� �虣�L���"O��P�2���
��U�:e#� Nx�<A�I��
�q�'�͏!ti���v�<��.�"z%bdӰ%���@��u�<�@IM���RD�^�=���7��r�<����2hH��� �Q����LS�<!��Rr$�*�ǋ<�azDo	P�<�,J ��1he%U�fJ��!h�R�<�sLOWh�9� !K�3~x�!�I]g�<������^��@a�48� 3sg`�<��M��/�0�J�� s�N��q)�_�<A��~�v,��i���e:S��_�<	�%Z0V�{�Ϲf��a��[�<�WA	*��i�V�H5��Yӧ�<Y !%;�`y����^Hk-LA�<I5,��k� ���
'z1�b|�<q2�M1&��4�ڹOLP�Y��Dt�<yCL]��41�����?�zq�7�RV�<��]Z�D�3�N0�ኁ�V�<�D�\&{�uI��	
!��j���S�<#ża�Je�b�*6�X��PX�<1 H�lЁ�*���e[Q�<�d I�N�藺Y`&*�M�AZB�ɧ4]V 6,��/����|B�	�/=j�H��R"%Z� ���R*�B��d�T��%A�� Ѥ�:8M~B�#3}��!wC	,z�ʰ��Â�V@PB��?x��e�b	X�$ ��#J��$�lB�I�-$�1��I��aZ��B��8L\. �ǍP2���p��,:C�I�@|Y��ڮA�`�sG�M�NC�	�-B��k��M�7�d\�D�8ehJC�{����,7mFkB�W�0C�ɫ=J :@�� ~�h&9X�C�I+KY�dӴ�56ur�����0��⟀E{J?9�ô?�� �������H�O+D������Mq��8� �V��zE��_�'M�>�	0gi���N$I�0����@#�C�	P�N͓�2��)д(ڡX�f�I(ð?	�X/HsH�q��6Rd��@��^�<Q��C"�D`�	�.1}���l[�<�Ӌ�&b[:L11iϟ^���c��@�<��n�-9]N�ط�W�KWJP"2��|X���O�4hU�:~Ex�0���,��,b�=O��=E����*�t���Q�M?�������y��/N��h$.A�	��@�-]��'Mў�Oت��K�Z��	����`®DZ	�'�L'"�6b��Lhq*�
El�4����-O`8�1[&Xv($`1�х]�J���F^����"� �u�PQCãG�5ij��ʪ�y����\��4ENa�$	
wρ��'�ў���<��FS4��r�4$ X�c+Kj�'�1O8���jRi̢'��\ ��79�Z4qD"OF9�C.Hw3�!� �ӹ�j1�Q"O��s��TP4�f	��,��D/|O��WZ�w���v)̜FO���O 0m:� �Mq�OB"4 黐�P�o;�9��"O�����S�4	geE�7A��0��O���#;��EH$�=N1`�E⍸&�ax��)�5���b<bh���#�ɐM���ȓy\p�7��`�;f�[����';�"=E��o��3}f�8���o�f<��f��yb/��c ���*�t�5�⅜4�'�a{��Q�+ a�̅ o̩*���,�y�`�G4����,q{�:����'ў�'&@R� p ���d�ʵKP Ƌ�y�l������EC�
��P��(O �IP�'(p��R�Z���q6�O����R"OV��ԁ� �h��~Ѵ���T�F{��I	.A=�s��	 �yC�+K!E!�dWL_ā��hʾ���(BɁ�v�'qaxB��@��g��@q���22"�5{� |O���?)S	ug�h(�O�d�� �W�'2ў�'?��͚B��6��e�V_�:�t]�>��[��ҏ�	,_��Tbcb�|�U{Pl��4;�'�ў�>YB3*��j=�q��ę�j�BI��i&ʓ��<ya�ύP��%`��sJ�H�aT�<�T�7�O|=K�o
0�~�����6x6�!�"O�Z��r�X���Ή ,wލ�c"O��C��C>0l]:�OZ�Y�`U1���Y���IC8).`�S�O�����{!�$Ӌ.��e�%���f9&�!�dH��H���MO��I�g�K��f����b?�a���IT��*��{�вEE6e��z(�%�:�p{ (ѰEH��ȓ{ۦ�3��K�d;&��-m� �������O��}�,�à�D�A��%��p ���N7f���G�5�1�^$�f��<��'���T?9AgȄ�O�4���P's	��'�hO�a��=��X4E�>(�� ��j��hO�>�9ң�
�p|�!.�QaȄ�*?D��bP�N[x@ȴ��" �*G�;?��i��{ڤ8x�R6�60�0�2�߇q���hO���Wv��]�ވ8(śF����C3]F�D|2�%>(�ͳ�%�&�Ι���A�Z{&c���'�?�d�����c���Q	��Rŋ/D�ԙ���3w��a3�o�u��-{"L�ϐxR2{;8���0>�Ʌ/����O��1?�b?�"�D��4jPk�7Ql�7J'D�8I��ܿn����/ �V8�9$#d��'1O?90����W���`��0}�v�!D��IvG
O�E�UlD�iL����!D��csB�4(np�G�E�L�ʬ���<���?���@\��v�^�v�ʶ�έD�ў��ɸBN~mh��:!׾��-n|"=IO���� �YL�5�+�g�䛇��ȟԄ��k
"��5|+轁�V-��%lZ��8}���i�|�pc���#4�����'Y2�mHF����	
�z���jJ�(��[����'8 �X�Ԯn��6$mFT��
���DD�S�&ň3��#-�����N�"?qOZ��$�0K 
�B�6�Ғ-Ύ!�31�(Hp���T�*� VK�>a8�J?yۓ0��x�^�M��9qL�&T� �@�"�����'1�<�j��@���1NҫAC�ɼTh=�`�)yr�u���8<�C�7#a�l�6B8<j��Rѥ���B�ɺ|	v�D��Wb9h�03��t����P� ^ر��]��L�w,�59!�$�)b�F����S:D�D�C�[�i=!�� ԑT$�{7�u`$��IqT��	y�����R�1���3so���fH�#�!�N�.a7YN���t�8<���'*1O?��?@g���CC��qC2`�s�/M*!�?YY�e��\6���F�ִI�ָi���F}bD�^�A#@1v@�z!C��0?�*O|���n��,�8�9P�((r&��4"O�Q���=�^@:� خ;i�&"O�ˑ'
�0�&a('�r�!��"O~!1�ՌE���j2��"O�$�P�B�(H�����h���d"OƅK�iN��a�!鄢�N�;�"O�쫱��6�(��A"G �-;V"O@u{ud
&@|4" ���Z6��b"OLP�������U� 4[�p� "O��S���7`B�ATm��iD�QC"O����H�4BRb�P��/�>uA�"O�d{s,Q�A���2i�-UT���"O`�G 48݈��p��(C�&H �"O��z���"qPQC�Y�I���;3"O�u��Q\v��aC�V�^�%��"O8����"1Q�ڨYC�9 �"O��d�.R ����I��#!"O~%2'&޿Fl�����ʔiV�(�#"O�dұj�^�.��\5Yt��S"O�ՃU�F�6x������ZB��W"ORQ�O
vH�K���,Q,RQ�"O��;S�4���Iׂ�l ���"O����Ȉ/�|4���_�,�:x��"O>�ґ�ߌ&�X�4.�
x�L�	�'X4d��
�Xh�]�ƜxT����'E�c� ͡%Yʡ�5d�����	�'�ܽ�uV64�b�r�տ SLT �'�=;e)�M��qEIЯdЙ��'ʩJ�F+�����1"N�2�'��$���6�0Y�
��.�B�'l�L�"LE0&��k�� }��\��'���ٵf����f+��{o�H�',���	[�8��,�F�>{{�]	�'��ڂL�)���U��<�ؠ	�'��
��C>��C�E^��� 	�'~�%Z��BՊ ��v�@�<)�-G�1fF��ǲr8���lAy�<QE�/z�v��&ᐮ'*`�2 �s�<��l�`�N�u��"p�H"Ad�f�<Y��ŧ}�d���CӠ�,��N�e�<��*�tLT��f�K�	7�);�f�<��I��� I�4*���,�E�x�<�'�̟aJȕc&B��nlӄ�_q�<aC�~� P�*��g�(4H�a�<��g�2qN\���O�
,\ؚ�W�<���99 ��`�I	st:D��+Q�<�Ñ#a��HiD�y.�\2��TT�<q�ĥm�@xe�vI� �]M�<���¶zx�"��8j]�T�I�<��(���bHփ!j.��BC�<u��`��90��N�	/L��!j�Z�<���@6[e��R5��6
D8�P�^�<�cGX'(E�d��C�4M�\��uE`�<W%P�"B@����@-d��uu�T]�<���Y�T�\��B��C���(KV�<��,Yl��QP��&�>����T�<��b�"Rd��sd���w~�����N�<��-�-+�q�/��%>�-���GG�<� ���+Q�0Kб��
9|�Z�s"O0m��@Y� ⬄;d@ʟl1|���"O4�H��I�T�����N�`�;�"OF,��G.��PB�픕����'"O�����"�`mʃ�b�FA*�"O��s�h�1G�ȝs����ԁ!7"O��Q��8X@,��ǅ�p�b�A$"Oh�a&'U�f_X`PvFWJ�M�@"Or��M�/�I�q�%QrL �c"O&�� �T�`4�T����"OJ���S�Gx�*ab��p��1(�"Of)���2+م�ׄ<t���"O��:Q��������Sy��Z`�d�Tv��"�j*ڀ�)�jY��1O���MY��$1'GG�`ev|�&"O�<!1�܄X*е0��
Vi`tJ
�'� m�2*k��<93f�;5�����'��Er�
7qX`M7�K�/^�T�
�'�Z�z�A�m�^D� ��S
��X	�'tFt�ЎK�bn��37"�1��
�'w��r ��[8�a[� ��P�'���A�֟��0Cn���PmY�'�N�00i�:p�f*#&�.*�!��'�*x!�J��"x�X�0~Ա
�'W���BC9��3An[5
3�!�	�'h
�" �A��D�H6���,�z�'�@�4�	)]@,XV����^��'�hq�eBW�$h	[5*�?u��`	�'X�=��#s�$*Y�tDB@���y��]
j}ti�0��aZb	���y���"S?������7M����f^:�y�*�T���sDs��:�K���y�̠%\}���6&zJ<i��y"��j��r�
�$�qG��y��G�/�X���B")~~��p&��y�h�����{c��#R��
��y��'���]�28^��FȒ�\���'�>���4Z�~�j3Eކn�8P���Uå�h@%I!h�*>�U� ?D�P�/�=p�H	�R(�m�F�@#;D��"���61Qhtr��O��1��<D�x�/��KQ;���cr�:Bd!���UK,��I��4ؠ�@��/Zq!�$��sYH����?d�%:�!K�x!�$ �rU�w�$P���ߌ��| �'���a��^�@�^����ɥ��QH�'���E�9y|<}ڐQt ����'ᒙ���р-���$N�[��m@�'�m;�	��A�u�çG�Ih����'�8T��#�%4�(�pF�Er��'�a��i��`٠�AK��b
�'�PA� i״�-z�-ϟD�Z	�'���҅��p��sꌮ9��T��'>�"��D� �DA*2�2�Tl�
�'���C7��5�*e�B�͆?[ʰ��'�P݋��7TϞ"n�@��	�'g^�ҳ����٦�?G�>�ٴXx�5��;�Ot:�	� n�ЊuL� k�����'�f�dhZ<f�I;G������xxg"�$?��C�("S��Um?.v�eLڎN��c� �5�M�Ν2"�ӫ6���`܏e���5�L)�C�I�ZG����38�Q u�߹R��-��D� Z��r�ZUG��O�L����<Ø�q$��!&���@Q"O0a9��[�2��WJD(�$�DES ;R �%ɓ��p>�D-"�r�3��$aZQa3
M���� G�3���1��O� ����U�\$�@�Rc�[P��
4"O�iP�úY5 �i��x�����N�{��-�D Θ����:Ņ�~�Xi��
U��m�C_��G{���T�bΜ��Lo�>�T@��5�Z���&̨��	6%m�#|�'xY��$R7E� ��f۴.�`<�N>���''J�EMP�� [4�τ&,��f�DS�
�� Nq��T#��e��T��-P��ѓ�F	�V	��I�>m���j}�,�sUؼ���8�C�O׎��O�]E�E�!4�袆�Y P8 ���'��T��,*�	^?����%@�2/_%o�ެBP��<q�)ʧN}J�ba#v'�[�(�->�=A4�y�s�7�'CB<��Nӛ9�|���[�'��0&���ߓ�$�@�˒�X�00Ӏ�7.9�����F�*���O�u��,�����	9]������Q����7`�Y��B≨~���bHA�D����Rj��Z�hes& �>+��bTLω-��\��	�.r���Ћ"��홖c�a힘�K�vM��{l���և�$��K��}،s0�Û	z(��u�!s��X��'�2�H��C�4˔@I�o����&��6�*}ta�3M�l��jk�>�@��R�A�b?5*SdLd�j�a�ѕ?Q`%���6LOv��
+�PR�'�=�2��8X�@,�'J7 ����X1+�N�S��Fq�$Ò�ܸ��[B���V���H�������.Vu�<�-�+BU�e�;�'[@��y��]�֭�eF>Mh�az#ؒ4���1 hXr�����&63�%Y��i�$��ڴ��V>M�t��^ƒ��C��|�̙����H��E�>!u���|�K�WVr`�Vϙ�W�y��i��W�X��po׽J�x��☯I:�yS�-��tٻ��g�.K?�qsM~�<y4cC9}��(�r��8~]����ڳF68��')�+q@��W�����¹x���"�$r^c�M)��N�vLX��m�:SC�@'�q���B'�ߔ��?�b�s����R��8���2x�| sqg�p��xq�D�0z_��W�Ʊsp�7*KER��3{�h(#�Gt��Ddu��3uU�6�<�8`��0���Be�)�I0���ŧ>Q�Q>�+5��9��J6��z��跩��^LR��c@+b�`���
z�2E��D>��D�
@� �O�6ʧq����ݗ<LB<ң�Hc�!!g�lB��'�´s�O܆����bKbdc�i9#�(}�1�J���E+�bʳD�l\���������?Y$+F�>�B�� ���{�+;M�،���U�;��x��V�;�@��,��=X���
P�1ti�3+��L�ؔ˃�5�T��)r��X���W�U�z ���~�����6nu:���l���pcIڿ[���<}k� �-�}M�e(��)w�������D^�#����g��B��y���I%dI��ɛw���.00��e��G`���'�Dݱ���TB, *�k�cSD`#����y=�m!�C�W�f�"v�71-�u����֟ j�F�aP@d�Oa�`����	6��`D I�څǥ��<9�fSh�)!�I����$�W;:�Ah�Ֆg��]�H�f�v��`��~��'VB�$���y2�M;lpq�C�6�M�Wn�7��m,�A�O	lE̤I�mΠ��Om�i�Bלk�& H �ϝ<� �k�Y#pɩ�/���a}"����wN�z_��C������a�	�}���I�Mn(��O
�P�ˁ�v�0a.;B����"O��ې�ìzlP�"F\��5�͏��8���f)s`a|k3�\R��(:<�M����,��=���$M���[�`�˱� e9����&��	�ȓw/"����׳�X�K`Q�g>؆�d9�	�(5=|��'�z㮀�ȓĠu�7�*N�
U$�!7�̆ȓC4��eJ���DR�'�1�ȓ �,�B8K�P��a��<x��a��j5�qҀ(I>��ehȲ�8��ȓ<<��R��ym�4��T�b���hr���f�C\�����f���O�sQi��$�t5p	�'ugҐ��.�=l��@����{�`��'}8YSW�??b��8��1n�H9X����ĔH�������?*�t	R��%���L�8>��ҭ�<-��*�LS69@�D�Bb�2w��,
���A�:y�S�dy�hH/a�%�=�O$����1�ܴ�c�Փ]�0-�����,�h "S&�SGzEҬ����!<��)��ѣ���a��ˑߔ�1�/��s�D"h�5A�����X��#�<�7��P:tHV��?�L�' �h����|��MR�#:�!�C�Un�>�Z�j�Ɵ(�Cؓ:�P����'�ѳ3fV�m�D�T�:A�r��J��8fb��$8Z�)z܏V��Ot��#�W��7M(i$d ���h����sG��e�R��)l(t��F	ǫ8=��CM�bT�m
[��T�#������o�ܰ�����'T�e"�i�� &q��'C����p�49[r�t��,t�E��oBw��t��^?)��m�h�&i���ZZĐQ�VH��-�6�S>��I-���#�-�&~�OXLx�ʏ)���b��3=q*��T�p�vK����ؑ �S�s��b!��	4�Ӏ�\l
p� 
t���aI�~�Z���'m9r�׺��=AW��2||�uH�/wҮ|�toR�v�t(#+O�U��R�M�A�ɟ�����}���z�B���"]´�d�ЏQ��m�%>��c��6KbB�RTHZh���k�@X'8�Pä�)E��	æő����2�@!�'�a�SO6J`�]�wlX�*8-��lP�G�^��T"Ov�"ΐ|�\�Cv��M�
�������>��IS#�)�C�_j��nWz��cM�y��h�C̸@!$��I<M`����&�!���{Kao�!:@��Cm��A��Ĉ�y���	���0��Xό�H��uRL��<Y���pXX��ao/�(�,�;���F�zipB�49J��ȓY(��&� D58��@[d�`,Lj��'���������8L֘�� o��]u �	R�"D���6��f����瞫$mx	7�A�nA��IVA_���>aШ�2�j����ǻL3uj�KD~؞�h�)F�OL�Ig�b9�H�1�~t*���:%�C�I37���k�^@ZD��`���hC�39d��蔃ɹ8�x� [�C��B䉡j�|�!H��Ahv�r���J8VB�I�۪�I )d}	���m�.B�)xz���t��-nࠠK˾<�
B�I%��a+�iUS�LK��(IH�C�*2<0�A��MQ��A���`f�B�	bi@AB�S�*T�9�n�61+�B䉪�nh�'�xR9Z�Q/3��B�'0�TU UF1�� �� ��a^C䉘O�0+bgӛ`9���g�RC�I��y23K��s$Ґ���"C�20��
Ec�|��$hu��<��B�	:�T��`/$!O� !��'{�B�I#Oy��6���(SF���B!��C䉔8�ظzFa�&b�NY#j�n��C��-v�����3J�,�c"QxXC�	�c�0A2��S7Uz�E�ǰ�`B䉟{�����W�,��'��m;�B䉉R?�8У'��8]�(fn��m$�B�	6��)��	�`���cҪ��B�	�"����0"&.ʾ��vg�DW�B�-~�����a��#��H`Q	��7�,B�I5h�v��w�!%��#�-l�B�	b&�y�%k��-��H�� 3E��C�ɖTTx<�sL��8�p�	A kB�C�I:R����{L���r��7�C��"}��=8��R�k������<sܦC�ɩ~�z|�&��4=L�gy�C��-�^���%ۂ"s����U�X@C�	�R�IJ"�W�@*�rr,F;q?�C䉵fELQGo�T;��r��%�C�I�j� 4F]�	��z�H�9lifC�	yx!A�o��Iٰ���PC䉕n����g��	���f�'Wk.C�	�n��h2�h̫��A�&�	%5zB䉋+>0aK�N�2��@�
G��B�Ɋ^#���د;���r���:C��5yV�=��@�=R���[ �;$B��-�١0��>]f0� ���Y�B�I0
��	V�`�b	�W��C�	�N|���A�g|��ua�{
�C�I,j�"�UC"R��򵩝�[Z:C�$N���k��e0�4�SCU�8p�B�	��Tt*�+>s���֍�xjB䉘=���!������*o%LB�)� �E�++! �)��ĺV>��Jq"OT����[�v��ɊPKɦfN�PK�"Ozቢ��1G��s+E�	�dh�`"O�Tp�@я /��JQ�OS]���"O��ڇ$�#k�v�@�&N_��"O�e@-ݳ'*����ԕJ;���"O�mBb�.�؈���X�G.�EAV"O�xJq/Y:O��8�n2wԱk'"O�A���$n�p:��,H��V"O`uX�o����hA�;���"O4��� 2�A�%ʜ0�\ղ'"O��@�� #��@J��O�T�zC"O�xjb�7\����@ �0P��"O^@y�E���u��@�ol�(9�"O�$ 1m�:e�"�`pN�D����"OԄ���p�=�SB��D0"O���#ҘA`�-R����^���"O��"�l�>�aoLḤz�"O�d�vg�[��M��
��Ȃq"O"���-&A:v�;SL� x��u"O�$�S��$� aC�K�L�$L
`"O6A��Y:N�9�E��V�����"O2)�,�k��b���\�a0"O*5�R!� ����f(բT'�q�"OԈ�A)���)#�	� ��U"Ov�а�\
t��T�υp�1C"O����RT}0�*���'Wm�u�"O�"��|��agi��(#:\c#"O���I�n��q��j�:*��p"O�����8r��� �.�	ehX�"O�%�ؕC���e'��+�J�"O�]@��ѴB�l��m��5�X��7"O�5�F@Cl��yT���d�"OJ a�X9�� ���h�u�W"O~q��R)jB�$��ԕ+�U�d"O 6��Q2�Q�Ƅ,�f�:�"O��kcFJ�|�Z��'��al굻�"O��q�Gǻ{���ū�(`l�@�"OddNM�&����pjߎ5�X���"O�D2vL�u0�A�����0f��j�"O�Ặ�_�vE�٪0g�IA̤�&"O�m��o�	�@��1� *O����E"O��9�iz�1�&�؞/j���"O����m�
I��S4��2m� �5"ON�B�O)0w�%jvn��"���3"OR|�f�Oaz�DM�M�(�"O8uK�@��-�а !Kݕ9����%"O�Bb�!kـ2 �K���t�d"O̐��ǹyhR�k��*1z<��"O �cU#!I:a�%��)Q��s"Ox4Ӄ�I���3%-hd�|3�"O���A�$n� �A$�H�mjDj�"O|(3A��1%W.�R#�њA�X��R"O����g������v�B�"O����~$����

���zc"O�`1f��V6 �Y R�XW"OP�e�N�g6m��Ϋi�9� "O�T0�b�d�������|	�"O�yt��#;찇���S�Fɋw"O�HUd�b�ԊՃ@}B�[g�i�.H��Lx� :�iC%_��P2�A8&����*\O��P��Έ>2��Zp����KC'�D�C�V�(}`Q��,�2*��*>.��`�C�o���<�@	�	l����#�J\|a.�� 8ک��ۄ/,⠆�S�?  -���o�LA�c�֤tX�Y�IS zq|H�N����(2�g~r%����{��.NHbuh���yr��,dȘ!��Lǽͺe�%�65��F�~ԇ�I4z�2��w�ʂ���H��V%8��ė�fK�u:�'��~��T#g@U ��ǌ��`�=�yBfV�p|��"�-�h�PCץȘ'�b�ː�֦Mcl=F�Tْ.>�mR`�T�&����3D������H�� �w�II��&"Z�Ę>��LD���$�*���cیX?�ȗE�7!�D�%d�z}!2jҘe�e8&D��6UjfL�!�,�Q�p�����$�+1a2�[s#�m� ��	�M���`��u}RjL�f#&)��/Áxy��[G�˰�y�Ų]�B�A�]�{��H������'�����k�OE���~���Q�[Ҫt�
�'IL�����RT�:�#)\=�]{�'7�p�n���T��.S�,Dh	�'ۦ]�T�H�D���үס��I�'H@�)M�$N������.�
�'����,A�xa�|�%��J	�'� �c�Ғ[+,,�U�ݦ���j�OҐ?�qOd=E��O��&�8&%�d�� ���"OX�B@�z�ؒ�D4E�]�d�%`�w��mX�h	�唘%t�	�E�ts����� LO����;:�����'Ovh�e,�Jϸ�x4�1إ Tf�<)��ݬ2��+DaH�5Ȗ�2Ԋ\̓4̚�bt��A�ڣ~j�fQ��fi�f�)4����aa�\��1Sjh!���B�8O�"ꁅ4�n5#�I#&�@�z FL�T��x��6}��L����ɧ5�x�p�F��� �A*RJ��lrc(�&q�$HP��D'��D�8¤I&��#)┹��:S𩸃�['b��(�428��`G*�~�Zcq��(W���S�W�ѳe�� |�x�R`Z�gs""<������%�7����	DM� H�-���'<5<�S5�B��$��Cua�����_�t,Y��R;W���6t2t�rr* >����Z�2b������_�"tc��.wN�zf�L����hĖ �t`g �+da���� Kz�RpY��JsH���M��Bp# �ȖU0���'&G3B1�dڰ�Ķ�dQM�4�䡣|�QlT=43�1��$�>AD�~jH�5�Ю���F�	A�� �W ԟ�ѩ[fh�$?��٧�ў�N1�D 
.�LLZV�}���jԐsO �زNŧc.��O��'	s�	(�A��=��EA�f��0�Cᦒ�<㣍]a|����Sl��x+O2��Ǩ��_F�0�R���L��A��|� �O((U��"t�	cV4�6Ƀ�Q1T��Sm��K�v�dQB 5:C�	 i���8W	5Zز	
�f>>״���ȏ�u9�H���[!SiJ���K�h����ɴXڱ�hL@��='�>@���/t��D�V�'�6X�rNP-p��L�'0@���(ՠ23�e�n�59��TG�8�V	�pi��)D'Rx�g�Y�9����WT��S7a�l�� %��Cg��o��4��S8jEZ;@���JI�腄Q�P�|�b핰U���DQIX����0Ƥ4B��K'�rMr7(�Y�'�Hbw�$�g~r�	|���Q�
�eZ�h�ڝ�y��@"zs�Q�*�/dh�qEP��,�G���0?��� �
���U�hi�Bp�<aQFA�q2�����[<ܐa\d�<�2 �A��P�3H*)zi��g�<1��w��E��)Tl���0��Y�<��IA��Ԩ�Ջь+��9�Hh�<�Ǣ�4��{�G"3p\�"7�2D��! oE�:Q)���D�&�p-D�ؒ0�ӈ�4u@W,C�%i�,��6D�XY��	) U���+�%G�l�7�0D�@c��dt�iq��'�
��c�.}�D�)L\�]>	��CS<�ق7L�/xY�j�o*D����쇠5_���P�ݓv��X�@���`y��].g�h�*���yRB8[����V�J�hU�ۄꀞ��?�t⑹X+��G#���<��6�Q�ONqb��0x3�0Ӈ�<A�ɑ9����'�4�R��ˊG�0�э�L��8Fˑ+!
����52�:��O.𩛃+Ҁx�4�(Ͻ�`a�B�;;�(�ǐ|��9Oj@�/"K�0h���I>��M:1[���Х�� ����-���%TO�1h�_>� ThZe��~T�FO�rN�X���'�lԑ���<e����	� ��M� 띒
O���Fř�%ٴ�h�(�%�~��7.��	�&�@ⓘmV��k�
��M�W��Ք��PGC9V�TQ�"N�y����'⋗;�a�RC�!�����f�n��ΐ�,;�8��OT$��k�&6 ?A�,��?{����
~ ��7-]�ocڸѹP����K}�e�Z�3�Nd����u���� Z�� ��	�
p�*竘�P�� �����,3(�@��A���'R� ��^�"�#:��%a-OV�;D��K4�P�'�����M����A~�[�O�I�p���w�N|����E~j)�����oE������L�4K��"s*R� rtA�"$Ƥ(��@j���<�u�J��Xi-��J�&>8u��r��
�O��8f��H��Ǟ�҄�1� �@���L�;�O�<a� Y��ڋ�ȑ�QkD�s��	ʦ�`���]&��')�� ���Uc!)��X� f
�H�0˶"O0l��/���RQv�)wnd[uei���@�����5jQ��K��O�d��/Ӊ-`@�YN�J�Ʊ��I�2'�bgǖ�L��d�|�N4:�S���ء�޴d��Q�/�<@� �8���e̜�UB'��5a���<Qg/�0k��3@�3�'{z��lú���1�Z�����O0����6����5{2��[���B]��'�`���hq�+�
K�@3!.
$bLD�1��)D���� Xcj�^b�ek���y4�'��>���\�:��頧C�8q;1�GC�v؞,.�#g�剬H��A�R/�s����'��S��C��,�5��.J�/���'���oL�C䉾
L��l�.<b�����o�C�	
0��5)��G&�w';#)�B�ɪc&M�T�ܳ ����	;j�B��;N�[7g^$6�ᐎ@+�dC�%r�1���aU��ط���h��B�>�tI�M�2�ֽcVF��5ӌB�I,v�@d�B@�Z�Ja!�.�)��B�I!+�0��4J�>�6q��)G�B�	�
�ʕ����B�켰��"%�B䉫"����Ϟ�9�҈ٵjҧMz"C䉦'�ĊR �����o
6�<C�	�t���i �ƌi�h)�N�n�(B�I�J�iS��E��h�*�Q�B�I�2����s"U;3�������!��C��`^�C%�� Q���Q�K�0�PC䉡;���� ��e��=�Eƞ$j�C�	�[�"a|	���39BC��j��;'-b<r(2G�PVC�	�|���	c,ʸB<���0�C�ɿS�lţ�Eٮd��=HaI?�B䉕U��( �Ȳc@\�{�'_�{��B�I�b
(�t�$K*�id��PD�C䉥<
���S3;�H�@�N�"n:nB�I��X���'�8hR4 Ā��.9@B�iլ`$���l�
yaCP��=	�'�D� *�I�%kA#B��N�z�'�h��2e��I��aP)h2y�'(��p%���v� E�w��f��(�'b6���!�B�T��7j�\���'
�izC(�%��H׮�l"heY	�'�h4p���L�zU#�л
����'zz ���L�R����)��'�`<��;]n1�+·m�a
�'�d�&D�E4ސ�6dV�k�	�'>��z��!H���3�^d$}��'�>)r(�v|>�b# сY^��
�'��x��������掸�����"O�ɛ�猡/�4�C6G���5�D"Ol�[#�_�~�	��r�^��3"O�4��' �e��1 �Y�O2��{D"OȜ�n[)K>mP�@Z�����y
� �hr��4�ެ[P�@�i�A�"OL̫V!�-:A�tN�!>$4k"O4iSb��V���"TL"'����%"O���æ(@��a���6z����W"Ota��
0`(z��P�X��4�%"Or��1o-Y r�  %}F ��f"O�ĹUcI�u�XDY�!`Y"�"OFt��d�[zT�ٝ/���&"O�D;Qg��PUIa��
lDa�"O>D�V��+�Q#O�w�B��P"Od���k-s�xɈ��K7~�\���"O�A+A*�$hG�U�bK��Rc��pW"Or��4G�>bTI�u	X	r8���"ODL��-Y�6���.�7L&��"O\�c�xGLAcԍK&E\��6"O^QPÞ�
U��	AMU�P�"O�����G�j0��� c��E�G"O�Ԉ�h�:C" b"�H��AI�"O�$��d�-�U��OF&�zSq"O��iC�V]�|2��r���Q"O��3LE�8RҬ@�K�V��2�D�*L�H���-ι6�*}($j��"�1OhM ᯑ:}��qS�ê_q eB�"O\�	*O�X�$1�Ŋq�<"O��`��e��8����f�A��"OZ�{0d��O�X�h��R�vI"O��$.�;rx9#t�U�6�V"O����F��0H�	�c��(�E�I�x�,G��' j�q�+�}��&2R{ �|y,Yi�'���,{���ccޫ�,�'�� m`ԧO8P�o� @������O�aу͇wS�*S(�ˤ8��	 2��5�'a​������~���Z�Z��1X�ኡs��SΗ?n���+��yX�Kyb��I�6
�LM	Э��H|飃.̢Ӗh��'.A2�k_�t`��'d�:<��Ңd5�'8Fܼ�I�")��`3y`��q�[>j�`X�P������(������!&	��u���Z����b��۟�|�ԟ�2�G y>�]`�Kƒ��i�Q��sy���C��&�f(�1mߖ�a�Ԡ� ��]	��U��Ri�Tǀ̠��Y�����M3��
ⱟ*���+փ��/{��
)��W��0��fN<b<����Oι�4����0|R��,p�Ip��P�)I�����ٝ��B� yƪ3gva�4L�6Q�"9��� ��aɃ������A9\�˂'�g�)�'5'F0�d�������cܗ����#�"ah����=�6��6#����*V�R	�l��(�u�<12�M�@c:��l�&��3q��n�<�$�Ml{�=
�7�9`��^_�<I0)@/q�(�$=w����O�\�<��j�	���>!��Bb�[�<1e��\1��;��X���p�$k�<��ʪМ�I��:#�2�kR{�<�獃
sjƴ��d���B�Du�<�#Q�!khъw��&��@s"�\�<��N��Z�R�Jpm�	"��h��Y�<�։X�|�F2�iQ�a`S�<)���-�jYC�CɈE�t!���O�<�rcR8=�"��AaS-,�X�(���t�<!��O)�&]�#E�&gJ80ag�p�<�(D�?� �0ؽ.?aR� VW�<Y�%j�V��/T/ۨ�1#RP�<q#♉Xt\���*gm��KT�u�<a7%L?{`�H�n�' �P䋒�R|�<!A���`��Av����h����A�<yk�	�d�:ҫ?$��:�aZS�<�1��tk4�@��;4�� �b��F�<i�h��C���xfɖ:�R�Y�D�<��/T
ƢE+`��DT�,���k�<1b�Մ�z�ǋ#�H�P�	f�<� �!��ˆ=Z6DX �'U�K�"O�`�ѣ��t�x�����,T��2"O���M���V ���Q;#"OfE�v��M�� ��ȑ,���Z"O�7��nX$��E܉�
Q�"O�ԈWIˊh������f�Y*O�D��-<.��1���Z<���'�`��@�tPH�cW:V����' ����O�i�����,V
h
�'��!���C�"�+�k�0z&��R
�'�R�$�O#����"g )I��k�'l�EB�-I��=�D�5wށR	�'x|�Q�>vޕ8T�݅e��		�'M���ԝ;<�X!�(�V���S�'"�,�ԇ��6�A��B�c����
�'/x�c�4~V�=��(�.hR�0
�'�J {w�A�7��5 w�.o" ��'R��r�M
�E�6Á-�����'E>4��#*+���i慓"Oo�4��'+N8i�F-�"A�E�M/B�5 �'��Q�)C���0Y�?�xI�
�'?T�A��,��d/�I0��*
�'u�}C��ظD64��Dƪ�z�J	�'}�IblDKJ�C4`Ԛ;r�q�':�(��N-p��C"`���`��'JzA�����D�x���Q�S�	K�'i2�g`1S(p3s�����
�'!N�y���m��ْI�T����'�����6wa��'��	TÖ� �'�,zmÀ�*�W,�!Q�p)�'���PU�D%�f̓��Tk�X@P�'�b�����)�Б�C�c+�0��'s��{�MM�U��K2`��W�����'��}j��!OJ�pS$!�g��;�'%�9B@��?q����)D�O7�xb
�'�������Mfm��j�D����'������8 ���p�D�q��	�'���Qel�40�@pzᥜ��6D�	�'!���AbD�0��Dçʞ� <��
�'WlI�&W�*"4�Y4m:qt��'�@��2�Tn�ơ9J�&qޠ]�'���#q*��5�$�fY_SjY�'��EP -�0��=s��ͱU����'¬�0�Z�OJ�Y`o$���'}���,^�bi�F��PH��Q�'��p���	)�`�2� ¬q��A��'�����6 ��R�O�W�z�'<|��$�N��]w$�{����'S�Q�L�L�|�AMʄk�� p�'��%�!A�}�B�����9\i$͓
�'S ��w�R-Y1�A1�*�=@��k�'ظ�;&��{e�4)V`v�* C
�'�dM�$�޾NB�$&�;����
�'���n�i���H	�6`�	�'�P���O������RIt��	�'[�|�$oE�"�
 �c׶v]t�9	�'�A����<(3ĉQ��U�XP��!�'g
 �Tn�F�z���?y�5�'(%q�k�i�n���C����'������_�F7H�����#cN>i�
�'��(asHҙd/�Ȋ1��W�☪	�'ی�Ѕ� �͚3��B���p
�'Md��D���ȩ�	\%3
dL�
�'�~���Ϋ�:C����05�
��� �����iΰ�HG��9�d� 1"OL5z'��Lk�`˓����.��"O"IC4n�$��>y����'�x�0$�|��䘕�БG"��'��H�i�n�^��ʍ�D����'��i25��h�:�Cݣ6Irp2�'͞0[TKŦ1�n�c���#(�'�l�BE튖?���i���6�D;�'����-)!P�±F<z��ʓ���	���[�r!p4h B��؇ȓG��$k�LA� ��Pj5d�u�ȓ1��s�g��O�V�;�R]�m��rKd���o�e����G�� }ZX��p0�`�"@��N��)��`��u�R)�vg�!#��:T�d��ȓA����j��u���G$��I�ȓS���Ԣ�&6�CŨœ`�����Y��h��!"x�+�~f>���jx��7���a�F^�!��a��i�P�١W�$87쁽l�<@�ȓc����L��5����8pL�Y��n���aM�62y�=bwG�6sXFH�ȓA.M3H+Q��Q�'�(���ȓL&��B���m�t	b!r�n̆ȓQ�d����,V��QR!#A����7P�3!�D�B�`��)^����:rX���.
�;�ґ��#��7��ȓp pؘQD _zP�ۨj�����b�4y��:�PD��$�l���E��؀��%��q��B �5�B��}��p��F�/ExNa���#[�R���PYX�`�c��l���ԭ�Y_x���&A@ͪ�(��u�["�3��m�����ۓ�r[��S�M�R�&���a��u���F�\��1�DJ)i�NŇ�z8\�R�lB�!PpܛE��%'dM�ȓ}j �iߑF6B�k���9W�Ԇ�"�X���ʦ*��5�D�B�&�(d��i�Xj���8<�����15Q�i��S�Y��Ă�@����7nN�l�ȓs��٨e'}P�� � Z�����@h��;B��d�,� b��p�,U�ȓ���qAn�xE�)��h(^��a�ȓ/��૕�ItL@	���n�����*�$�kM�WTh]!FMSJ<$�����u��O�*FxPwZ
îч�7H5�5雫���A�A[�ve��<0�)[Ŏ�^���@O� ~���TwBEk��Q�{y�ฤȜ<�����1pe�;<R��`#�T�����J6�33	���q7c	�s�Є����� �(S�H�u����7�JQ�ȓG�D��:X��)� ����l�@m��B��R-�f	��t����ȓJf&��O��v�R]
v睬����ʓ�H�{7	>N�l��4V����C��8Z2���n2�	ۤ%�-$2!�DƑ,����E/x$��e��os!�D�@��h�AR,'(,Ր�n��-Z!��ŊCDD�	um:Ljb�B�͗c@!�dوS��eCwL(Wt\l�RC�(g�!�I�h���(��;_,��$-,!�P�
"͸C�ϑ4OL1��� ��!��=E���%�*I��f%@6!�� 
Q�hV!�X�CH�gHV��"On��r�E����~D��J�"OJXCbL�I��0Z��ҁ-�p9�"O@��Ѷf9F]� 
�7\b���"O��A�۬8��P�kH�C]j�I�"Ov탆�ܷ}xx�B�J�?c�"��"OF�Q�՜�d9�II�"����C"O�hXހݨ�ᗕ'�ѺU"O.0�a���D��E�AL�X 37"O x8U���I+�T���L��j�"O:U��k]�]NP}�b�ݿ$���7"OR�� "J�j����@���eif"O��u���Q���#��_>!��`p2"O��pdJ�	&�FI� ۷f�R(��"O��$�
&7��q[��-'�l�"O;�FǡM6Pt�1]K�L)�"OҌ��jZ�{v%!A�	jU��+T���1��cXVI9p C9FʺP��&D��hr)��9A�}�B-��w������&D�|!��ʦR�P���@!O���A�$D�,{"�?!0�x�f���L��H"D�@��셝G�4�q�=Z�2AsQM?D���$ �J�v8cdJ�^��YaW�(D���@H:���0Pp����0D�а���x'(8k���4�!D� �C� 4Z�AI�N;�<��"D���Aa�	U�4�K�*7e�V=2�*,D�8ජX��j-�M�9�BI��h$D�Rs�B5gt�=��þq���3'(D��JD�6�8��N���H9�n'D�L)�C��%x������BEnt`�0D��a!��+D�\�tM�5��x9Q�"D�|���Q>	<Hi��P�+e��y�i	�I��x�u��"L�9ۆ���y"i�,�0(`c�=�`�A��y��ɈE��h�g�	,kN��:��H�yH_���5z��10�kč���y�B����tϞ"5(z��46�B�Ʌ@���b`o�7$+�}
d�L��XC�./y�!�P�U��x�AX�g�vC�	<F.��F.-x�	���C�B�
C�	<�tȡ�E˥y�Q��V���B�$uޭ���9YVu����1v$�C��+����s�,*�$�PA�Ԍ4V�C�?x����bOw(��Z���r�ZC�	1�.1�W�6#�`s&/9�.C�>�b�� P�fC�h�f	G�69�B�ɭ!�	��/�18��Ż2,!1vB�I�}���ɀ,U�������,�C�I0��+ ��*KS걀c���Iz�C䉪q8Z    �