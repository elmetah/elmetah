MPQ    �|    h�  h                                                                                 �B=[��u�������k�M~��|��z�.<��H�,���A_9�Qa��i�/c(#Fo�nLA��H��7�R�%I�n^�����9���u���09����{��w�7p��D������p���!�����%J����/�yq�(=e���o���fQ�:�w�(P�u��+�&.�5��0��ʙ|�[z�	a�Ξ��Z$ʯ�����QbBu (z���ɚ��e?�����_��7�����r���`�O���Qy�5���cQ�I�/��Z��g�5��f-��{mU�MW����:�h�����.L�l�ܙ�Q��ڃʒS�{�յ��q�rK1r�mm-�G���ё ����F�R6P\z{8��d���.��4��<vs�������U�3e�ڶ��=��_P�������ϔ&�7��
�.�	�C��|7]�$����wD�Y�^[� ���S5�q��;�~Y��"�q�떻����B���t/�Qr�&�JW�U�9��L����%�,�|�S���@�58u��[?R��3^�R����ۊ+:ﴇ��IV�5n�������n�B�\���K�L���J��b=���K��r�s�|��� ����Xk}-Z��V���Ը��96N�ι�V��ߣG��_Dʇ.�fl:�Ĉ�TF[Siy��h�7�x$��y"��A:8)�|��o��K;)�kYXx2)0(ۉ2��>��q���f���F��z|h�}��[7
7�EHB6Da��I��7S]Q��miFl�]���S�;$�TWW�G)K�#o�*rJj09=�
H�n�0NYe7|h�,��]sw~�8�@i� �x�������*��t�2��)a&E�N�������9�EK�,�_J`3����J�*M�0|๜<��I���Z1#ԭ@PaM��6�V�n$S�+����k�g��t@�?��L��)���ȉ����O�M�����X6_+���r[�����"��O�-�˸�0|��{m���	�=��*��)�.崳�D��cʮ��3��r��]-$��	�����6���.O[��=����{�s}*ܠ��ϣ�C�:���VL��RY�k����Eq{����Y��n1���@�>��;��y�äf=,"��_����W~��Ʊ��l̀��\a"Z&*r����w��c�����%]e�y��hP�*j,��5�������CF��K�*��@�9<�Bo�}�>B�|�/�ԅ�V�I�,�A��Lm4���2V�J����#���[�磪��h+YM@=�2B���nΑj9���o2�
�YׅxJn��@�G�s|���T�x�v�..�a��}<��A�
��"�jzd2uAWf$E3N����f�@��v2�/6����iP�|x$���L�ێ�M�P\�n���<4��٠,%�E�o�7W�9BC�U����7�����N�.e<��/��v�_>Z�_��e�.�?��ó��EA>!P�j)�p�f��((v�")��p�Ƹ�>k��\p�	�5/��Y-t���ܺ���q,fg']��-"2�pu�p2��3ڍ�f��}'b�4�(~����>� ��Os�ϊ�����ܸ�-4y3�YN��w"w��R��/��e�Y�����8�pB�����
�1��B-�@�	��U����1oA 7^T~��ie@����K����ynv��"�������L�����ylVx�j�.1�`�Ĺ7����-���:Y�;
xU��z���-u���7������V����f����i#Q1|�~�N�Y�l:c��f����H��^?D;BJ�Zj��o��J�`k��j��#�x�D�Pr>5Rv�V(��E�S��	�.p�B��ڈ-D�����W�N&�+1d�M��a$>�E*q�H�/�@�B��2�"�t-(]g�6�CM2����@P���(�n*6����L�y[u����\^����_`o���B��/������<@�S���9q�IC�Xe��c������"
8��L��?DDv��5j���(�[� �0���F����QyuE`j-��O��v��8��«��گ#��~���l����!
UT=k�̙O~�l���J$�v�W��t�B�` Ԙ������W4�pZ�)��8KHնK�Ng B���T�G�q;����3��DV��������]��~ꑢ��X�%����M)�]	(�8X h����5KĲ�]�eC�ͦ�4���O[�&���d�[�D�1]φ/�Ĺ=+�N͞4��ѯ|���5�|k�qzt�:�����t������2a�G�l��m��z�񊅞�=x���j�$��f[8��l�����3�؀�i�^b�ٜG����<�v��橎 �ŀUT`�R�Bj3�ͬZR����:{����~:?��5�`�M�bm��	 �@L����>o,L���0?+.�g��6���t�3r�0	�N�́uD^�B�,]��*�^�BƋJ�H�w@ Sl-����`�8B�:]1���ey��F�� +����mp����5�?�����L{�D��K&xh�Yd��u��b�z<�[aS\>kO���+8}Ez-�8-y�y�U����&7a�%p'�\��1I5HX���0A�8�*-1$!~�|�*����1[l�M�j�n���l��)4<�'��M$�RS��W$��>�T�x���g9*�[H8а�ڂT^�7 ���I�P�G_�}C-��^_TS���w��	Z��%�΢���Დ*�ʮ� BX��ji�繹*���舠�JN�\ �u�4��� Qm��Ú6�~-�'�Vki���o��uJԄ�",�Ƹ�KK�`����c���߈�K.�a�8�O���3�����	���0���{�l;hM�D����qX�vJ�>��й{C�(��`g�n;\_�B��=Ѡ���4�o@�Ճq]dŪ�b��z꿼e�6�狷��or��lp<FGr���%���[ukК)�N�.��s)�S�����w�$F����fܽIb^3-%��ܟ�u��<��:�Q�R��̔�M��"c�Z���pN�H��yJ�2)��$�ѵ���xI&�=��R���V��>hOH3g�2\���F�i6�|i� ��oX�'o��#*�M�l��!_��,;�G��UECH��5 Ni#"�>
�7!'qOk��4�-JZ����X���qĂ'�u���74��V���k�+bA̤|]qa�c���zP�}��Dה�7�8��p1bԎD �`�����u��b>�I�-XE�e։ŭniР0Q�4�^���Ok�����Ldp7e�6х� 5{C�Ĩ��Z���W�p���*�v:[8�[�n�4��3p煕�!c��0�J	��G�FH�4�{S�h�߫w��0R�o�!<X���_�1������p=�B;u�:�V�JP��b����r�ٲ���$uʪsŒ]�|���9�߁��Yi�/�t��_�SPb�wϐ~4Ǐ�]Y�ޗ��a�p����YtJP}r2��%̐U�����E_�-�7'X��g����5Δі�%�7/�^��p�Uø���+U@q�n�V�9��St�jc2n�|���ݽ��vL��9J*�bqv��?���D[s
���e����uX��fZ�^&�<�޸��6I���l��h�b��_�.r ClQ�0�#~�FV��y¢��%�$�"*:#:��|4��o���K6�M��~�X3�0C��2c׊�̺���La�w���hB��v
7o|.DW"z����2O�Q]>�m$-	�x��1��mT�#�GĞ�#j�&ru��0��F\V
È����Y�hr��X�~
�@$��&'��ϩ�e��t��5�7j)�"�E^�A��QZ�A;.� �/,�L��������J,R9OC�����*�J�n;q1^̏@�`n��)�V)���u�����斏��|g�z��L~B2�>�#Q�i�j�o�Y��3�f���1���uR"�;���d׸�[���|Cm��	$W�lD���}�.@�N��;�c�ĕ���E�M#�̘8�$W�*����ّ�������>�y�N�N1b��"�>�7�5v,��E����2������yELڌ��F��-�n,�_������;wɗ~}�f6Ĥ����7��~���0f�;T#\|�rZ�Yrqm��Y��w�̃�M[Ҁ��4�thkcCj�|)�.��3�ȅ��F��ޅ����"W��oV�>�L�|앜� �iV�������X�4t�2ѡ�J�5��ߔp�9X[�V�Wh��Z@XF�B���Iib�����sb��:��-�x��뛙KG6���XT"����.p;ay~}��D���
	�{"�!3dmW�3I�݂6@�%�M3��HJ��fhi�dlx����G�'��$RPn��9��Q��i,`g0�
�w��9�E�Ua��R�C�H�C�	��<�A/R�M���Z��b�r�I��A���g��AyؒPh�����f*$J(1U�=����Ɠ���w�\���03S4��-�Z�������L���;�����(��2��+���N����"}�Ko��(��׎[>q� S�ys�����Ӟ��1��l�4eY�T����&�M$'�����8������F-���ܻ��o
aQ��,�[&'����U�W�lo� �e�~�˹��-�|�ZK�v��z�v����I�?%"v����yk���olq�Tj8zv�����#��t�v�(=C�돠��xp+0z9E�-P�l�r�ؒ@V����B���0�#lO�`$N�j���f��=��f���(R�X0�D6D�B�v�ZE�������Jk����U�x��$P�2�R�/�7��:̰[�8.k���uQ���+��ూW�&�=�d�(�^Vv>�ͺqߔ��S�b �G2��zth�Pg^�5CH�ߒ7�P���(���*��lݽ��y�o�,k�W|X��`�`*(h�]6B/5%����i<{.���*4ZI��de� �����o C
h�L.?��[��j.)�(��W ߦ�y.@��Q��r`9��J(vKc8t�=��t�U4ּ���j�l�"�%D!eޝ=&�P̴�O����Ԟ$��h9*�hBM�^ ����D�HrX�K�;)�p�8���F�ZN���ƃ��o,�|֣�߮�n6D�]���ǩ�3˷�T������g� � �m�����+U�3��t�ؐ���PC�� Y	e�	m1�D�J�P&A���[�������
"`���2G�/٬�
�,�|��?z�!��@ԯ��ǑT٣�	��OA����<͊ {�=���=���V�fVڰ��~��P3�|%��3�^=�7�����zvv����,��;�|T{��R�|jbV��O��2K�{��[��q���X�`��Xb�o��u.�{T����c>j/k�Vv����F�Fg$6x�tG��˃gN��с��۝�.M,x�*�dB�N5���XwۧGSg�3���`��N87}b:��+���z��o̘�p?�3�����p]gQ��[S?l����ZL��:�$�&s�JY��ruǉ�}����<�\y��O��+3w�z_f8��t��J�2#Ź�^ap(p�z�~����H�
.��n��fI�G[$\�M|��B��T1���M���܉Q=�^.q��S�4w{u'E��/R�h*��ź��0���S9e�	HӢ,�ըJ^3� Yo��dcZ��X^A�	��T���ry�	���%s�0��A3�!%ʉ�}������u�*;.�CG�e����amu����� ��	Ji6�����,�k)��s:ϖ���Կs�,_E����B�Ek�T ˌ�3��V$�<���\��������du��}�&���:��]M�#��(����(vE�����tۮC�R_���@ny@�}G�ؐ<��WH��R(�>�)d�Hb�g�z��q���!��9*���h�ʯ_��T�pWFr��%�e���C�5��N�Q�W�
���}�wKZ�F��N�C��XJ�^.Aȑ�o��0�J<~�:N�:R��Ҕ�1��xr�c��b�9��p	u�H�o�J/������fOx&���<À�k���O�b���,\�N��	g6���i 5Յ*�rB�z!*��l�g_Y93;�������H[�! i�"G���q�{+����(U��SMXZ}qˌ1v'C�3�nW�4��=�rg6~}A':�],�0�~�)����X�aD�7B&X�Tb/O� ����P��v�=��I_X�I�ք1snĻ0��y�u��\*���ZňDd��1�V56%Y���b��G�2�dH�o3�@�R:�yz�\SК8�Ү���p��!��c0)�Ů�F���+d{n���Z~��|R��Mt<�\8�흽�dFH
�K2��X���􅸽�+�I��:{E��Ѐ�D�?:��-�]����3�jz\��T����g����SkQ��j~ꟼ��&U$<��Z:�˹Z�a�te�r�X� Ӓ���f�,���	��Nͨ�� ���U�6W�5�F��G���J;^�P.�x�2�Q�+p�u��#V�]h�������n}�f������L�M?J���b�?C��$�56�s u�z)��lMX��'Z��9�U�wO��3G�6Dٞ�o[��#u�}"�_:�X.MEPl���ľEpFQ��ya�����$'
�"���:�*|or�oF��K1��!�X��60^�O2����G�%\t�������n;�h�T ۑ��7����8�D���!-k�Q��Wm�3J���u��v��T�.G_�#e�^rж0x<#%�
>u��%xY�th���S��~u�m@�����^�S1ު�@���tH���N)?�EE9��FҼ������,3ZT������@J��E
v����Z��I��1��@��G��<�V�3#�O��QB�a���e�����<L����~�~[WJ��Kz��gM��4��E��&����"F=�8g�Ħ��+m���	_���R���0.�{��2c �Z�)~��(L���|$�p���:k�졧����
`؂�n�)j�V$��!��0����ԸE��-��~gE'Y,�,�����gn'm��k�ȴ�z;5n���W�f�_v��	��Ң�~���c����p\��qZE4rLB���7Y�3U�������.�︒h�0$j�#��v��@� �;F�G8���{���hrCVo��>�w�|'�Ի��V�����Y�P��4,�2L�Jw��&�S�/[�_%��d�h��@s��B���$ꦑ�Q{���������x����G��;�+�T]Ka���.���ai�}����� 
�Χ"���d���W��@3DW���@[}ch�%{7ͯ��i�!pxZcY�Bz�F9P�P��tu��c,�/O��|o��9�g�U�i�m���O���<>�V/����[�Zx�_���dҹ��m�B+�A��xP�t��f���(��؛X������n���`)\�֏�+W�Ed-��uL��d�'�7�/�F4 �#�2g���E&�i\)�\��}�Iv��6(����H�>̼6 �s�L]π��aߣ�.w�4���O8��-K����]ߒ[�T�r�'�B�ߦ����3�
^��ȸg�v��s�U�܀񧏓 m��~�����7d�K�ڧ��0v\�(��
���,�{�<���݉N�l�(�j�姂����/Z7����#���\�F��ҧx�~�z���-+{zɭ��-��V�s �q=i�i�
#��2�a{N_�̌����hZf�/!��.�"�DQm�B�yZ ������k��"�c�\xt{P�FRlǻ޽	���8��<1.f�����m��3�����W��)&joMdH���j`>�u�q:<����	�+{�-2��&t��wg�LCC�Œr	jP^�4(ͨ*,n�ݘ<y���UR���7^E`��j�x��/����|�<��|�"SK/c/I���e?4���-��p
�E�Li��?z�Y�w�j�|(P�� �<d�e�[��Q�T`�d��E�v���8/}������H֗�H,�lS�o�z��!���=᢯����b�3�`��$7��;"�`B��] J8��.��ì�&N�)6T8���A�IN߿�n5��G���[�����OD�5j�Β*���Q�ʇ��$f��f��ۜ{��h�nZ�.d���p�K��k[r��t7e��CSTj�ÎE��&����ڞ9[�B�'
���W��/ E�_�*��e���<CH|��5zj�u�^�j��7�,���� ���%ְU�$���{w�=�o�x�6�ZE�fQ��"�M�<0w3�@2�_{q^�������лv�~��DYt����T�L�R��Cj�C��lQ��T{�,��4�W�g��`�ahbcM�����|$�S�>eRFֱ�J���#apg�Gj6SD�tSz*�f�N����+�����,���*�%1B|1���wv��Sb��st`���8R��:S���a�����T�k��q�H�pּ��,?����L�*夿��&n��Y�u������2;��\�	O'I�+.��z��B8�b$��K��Ŕ$vaJ�1p],R�c!��1�H���u�7Q�����$�H�| �����1��MT0ܤC���c"�8�4��I'�z^�$R	C��O[����J�m����9�xHn�����^�"�  �+LȾ3���DkT�-��m�I	�O%.&C��􌲉7��d���z�������QW*`�&�����'�R�}u�6�+i ��s��s6=k,��~3kD[x���z��ͼ��*�,�������,��֧�AN��p���R�i k��0��Q��85!��5��b�BM��k�c����!�v@~��x�/�C���Vb`n�Q��sp���*�%����L:d��hb@zҙs��`�:�E��.��%x�z]prf�rz�O%�� ��17��tN����dl�ɦr戜w��$F\ꢄ~���j ^)u��<#K�뭦<(ta:ɤR�����5���c�㧲�`�p�?H�P]J���ʗy�G���F�&бq�yE�k���¶O>���\L��|k�6͆�i[i)��M]����*`Hl��_��;��	��+H2 ���"�����*qū��:-��#�r�H��XS˧�1'��`�I�\4",y�
�y�sA���]���hB�p'3oxDM 7�3���rb�/� ṕ������%�J�IK��X{�r��Tn�&0�Vy��8y�En���?j �;d����,_��M�5�&�����Pu��y(�F����<�:۶���е\��)���K��!�Y�0ĝ����F���C�{�����p+�W�~����<G�n��U�������+EϚ8�A����@���a����?�~�;�5�Z0�i��]��9�n@bW��O����B��S�✯mV0~�, ��u���ؖ�sc�&��Z|t���r("������[�Ǒ������6����M��<���H5��5����m��^��'��Qb�8&+�B�V����}[점nxP1�mh0�>�4L�ɬJ ��b�. �T���GKs e�����'t(X�RqZV���$0���6?����j���oz�t�_�*C.(��l�z��Y-FL��y�וh�$BG�" �J:ɘ�|�]mo��K,���|)�X��0y�2Y��f❁`RQ�7�`�9���� h��۬7eI��~�D�(��b(�;Q��m�Z/�����'8�̖�TnG��#`��r+�03�>�
��ٽ���Y�h��V�N��~�%@�R@�ɮ�ޅ�۳�t㈤�Q�)r{nE�5�#���7`����a,n�~Y��d�J� r��;�
;�� HP�$U.1��@!�ؾ�ozV���-Ջ��O���C�@����L�w�����a�����l�O�����77�C<����Q"��s�^,{������m�4�	���%�~��.��d�upcQH���I��a��$�\���G�!�_U�%�ۂoqٚ�A�Q���tx(�+�.�g�� ����*�.�E���g2�*�Zn"b6 =�o�V;P��tR)fΩ8�4���m�~�h�����ͱ��\��Z���r'7g���ǧ�ʕ�CF�6����h��j�}�}7�=J�Ȼ�{FΝx�;�Ơq���oL�6>���|b³�VhfV���=&���4G�|2�ΡJR�U�O��[�K���h\}b@���B��������T�j��O�j:�x{3��ѫ G,I|w�T���G�P.�S�a��}mw4�m�
��?"��td㋌W7�3?[L��˼@�����Ͱ͊��i��x��l�=����3@P�S��Ο���^`�,���@l��9S�/U����>8�����<y}�/�5��	Z�G(���S�7�,�ΡA��P�[�{cf�4(�|-�s�����IcjO\Aw�&����-II�5{@������EDr�Ϗ��2�ۃ���ȄM��ש�}��p�ǅ(O�#��"'>'�E �Fzs�(���e��<.�i�U4J(D�J�B鈏sãܔ�$V��m��M�l�wv�Ax���`
�Z�s�'��jZ�h!U[�#��ϊ ��~�!�v����I�K5�����Cv7C���U�[g��v���/ֶ�D��l���j.qł���j�巪�p���ⷫ}�Mμx��z/�(-!��d��
eV}���X̰$�#�����N:쳌��s\Yf�����t���3lDl��B�/XZ�z�� �!�S'k����	x/��P�z�R�~�d�������.a�l�+j7�^[���>W�&E��d�������>�=�q���`�$9Μ�@�2^�tސ�g��C>�h���^P!�(�*�T�s�y�݈b`uM���{H`���ӓ��/+��WZj<�P?���c*�VIT�e�����m�e=�
�CL�h�?�o�kWj��)(�� �^o��68lQ*b�`;��@cv%�8�p���cK���rOfg�l�o1�u�!Q�=�����*�ݼ�;�$r���\��}�B�\ �w�I��>E���)P8��<��Nx��<y�����ry��8~����D'-���}g��?,F`���q��]W�����G߆�.�7�))*h1�谆�%��QeԻ\~Y��;�@~7&��a�J[:�ͷ��y�����j0h�l�%Qy��~x��y|��Sz�U�9�D�%�Q��{\����X+�S��]���x=�`ٳ�Z��S�fL~��}�t��|�3�$����^�FĜ�����I�v�+Ω��hű|tT��Ru=�j�E����h�D{���ʏ@�"�%` b�J�����Ĉ��k�>`����ʘa��|�ag��6.��t�����N��m��L��s �,��*��BW4[��j;w�}S]X/��l�`<�v8mS�:�l��|.�7"��q�|[H��$�p�d��(.?b0�qE�L,�C�Z��&iU�Yugu=�?�M�����[\�UO¯�+)�Hz9G8^��L�Ƒ��o�}a�d/p�� �h��B�1HMJ�ݜ��[���$��d|��:���1lzBM�ܿU��T��=�4�R'{"{���Rd=�����.���Q�j�99�#cH	����T�^�Gp ���&�	�߾���!�T$� �h��	k1\%�ٴ���nQ�?���;d�;����M�*����*������D�um��9�� "0����6�L�X�Gk_�i�r�i)��5�,��׮��E�q��������;c��eT��v� �*Y���uN����Q��Mxg�y��B�Ov;*�O�����C,���,n����p��������մ�dJQb|8z��ż����8���Mڀ��5��p��6r�#�%����@��kJNC��N��Z���wAW�F7H�����܎�s^$�b�������<C�i:D~$Rp��4Z<����c�)��^.p�HR;J@��Kܙ��\��\�&˛3��n�&���ݢ|O�!�a�\�B����6�;�i��}���,x����*;lZ0_��;�g�fc�H�{f �Op"=�����Fq ��Մ>�˘����X�H���k�'9Z�$�4]����StGA���]���� C���,z�D�gh7xaJ���b�/) +���37.�l�n���I�!�X[�ziRnz��0�푣������0Χ�);a�dA��'�C��5�H���f�����脼���i�u�~:l\������РҤfC�&D�!�$0_w��� FYD\<{^{���P�W�2�,� hU<��<��-O�B�	�~?�F_���)��â���t�a�û`������Kk�u$��^m]aD�����qQ�JS	@n����S��Я�I�~ŏ�4��m����ɁJs�׽�t��0r�`ʊ��P�AQ�b�C����5�h�>�"ZK�,J05���G�����^��]�. R�Ǳ+��V���,V`��]��;Wsns�W��A*���iL�e�J��Xb�=����Ηkyws��]�0���X��BZ|�����w�i`?6:��%�����_��%_0��.��l{���4lFGlyqѕ#��$]��"�ې:���|�h5o|��K'���׮�Xd5�0�;�2�Y��A����h��҄����$|hs����C7�����vD&ݜ�@�#�QnpSmU����Ա��v��sTCHbG�Y�#[��r���0��Y�
4�꽜}YQT�hC�+�I{2~+>�@U����H�"T�`~���t~��)���E��4�>��Ҳ"T��,����r����[J=���;�%{�UU���1un@�"����V:x"?+�	�%�W@жT��+��LOB\��7^4?��H9��kG�ʎ���������q����"��*�@�������mj�	�b�=�ۖy9�.Q���0�Qc6�]�������Ie�$(hݦ�٢>\�6ۄ@'�������܌T���$�&���ݸ�e��v>����Eݶ;ᢵ���r�nw�p���*�6;k���lf��o4��~�H��n�lTx\��gZ��rL�
xj�H���z�Uґ���eD�h�*>j.}X���x��V��F��ޖ�q�,e(�
oǫC>|-�|�������V�_q��er��;�4b�b2BDJ-������'[�W�h[�ht\@�P%B�I��K@�V�@��=C}�4���x6����dGG�%+W�tT�����4.��?a�}(����
z�C"`�d~8W�J3:Ƚ�G�[@ь`���@��eLSi<��x���8ʳ��jgPHv��9Hr�r��9��, )��{���9��U��䣀P�@����l<��|/#����PZ.�P�&��R��Qإ���A*ӠP9A���2f;�(b@��U��~*�$��W�	\�Wv�!��E��-��P�\�wz�ݰRx�|�7� 2��\ٯȟ^��R�
}��; �(���>�5 ��Ps�$;�v喞�Xܤ��4��E�����~���U�Q8��(�����n��t��3�
��.=n��<p��}�U6F��0� �<a~�|�i�حO�KPN�v;#v�o�����9"�q$������O�l�X�j�ς{�ĥ&�E����4��Ux��Mz��w-��E�#���c�Vx��'�ϰ��;#�i�~ĭN]K�X�@�p�f��9��eD�UB	��Z֖�[!���k�+K���x�w�P�ΝRbV��+ѡ1��,��.\�rƆ&����1iW��& 3�d�Bz�/��>�%q�ꎍlcT��q��29�tIcg/u�C9>ǒ(�P�~�(��*"�y�N��yGYS����H����`[��Ӯ�/��3�2͒<,v�X^t%�yI���e����({�����
�a�L�A�?����Ej?��(Ɩ� 0Ɂ�4��QeF4`���;Bov\�8��G�3XƁ��M�S��Ul�FK�p�-!v:�=W��@4�X�E��=$��q9�z�x��B^�[ �WY�d��ڹ�����)� �8�:�7=�N�=������+�����p����D�D�Ĉ`�D�F���Z��g@����������S��$����Q��Y������Xe��.�����;�&R`��Pi[U�`�7u��#ĥB��ў ���j���Z|��z`�a����`��b?��N1�2@��4Ј�'�qЯ=��~���R萂�fG����{���q3�(��Uj ^ν�3#��K�v��h��]�lt�T�
�R�uj�gQ�F����{�<������݀�`3�bYh�m|ڱ,-!���+>[�0�g]���O��g���6	�t�@3̜��N����9��.�3,�ǋ*�l�B2W��4��w�SXQ��)�v`���8��%:Ik]�W�߉r�Ҙ�"w;��g�p���C�W?�y@L�4Lg3V���V&d�Y�y�u�֧ξ�(D	�"l\*(jO]6�+$%zp�+8�/�cAqR�J�ua�!p��'�����H�Ȼ��-���T:$�|VN����1�i�M��0�ڇ.��.��ob�4(\�'�O�ODR�W�C���I���@��Ec�9�H�ڰ���U^D�K ��6�����n���uT�Ho�c�	ơ�%����X�����l.|������ie*���t�v��Ð�H�"uH�Tt�� �{$���=6��+�� kz��䟶�D�o�p��,0���RQ�̹P��_��&�7���͝��;�ןs���
�uj+��d"�+T��X�MMS9��ن1��jGv6r���Х#CG�Z�Lݣn���.0 ��`��0��IG�o�'d1�b�P�z��g�Q�گpy��ʊ��'ɘ��wp��rp��%f~L�Gn��@&Nz�w�hկ�?.$�~w�VF����3��)�^=Z���v�aKK<^��:�w[RK��o��Iu�c�A�J}�p:ҌH-saJ��	����2�7�&ƥQ�/����iQ���SO4����\����/6��i2҅[������b*5�l���_*��;�ϊ��H�� �1�"��գ��q;l߀p���6{��RX�^ ��8'�w��v�4��C��oC�A8��]]$�ϸ+�f~,��D��D7�����b@P  ���N�n���í��I��dX���u5ln�=-0=�N��4��;��΂!�v�Fd�a�"m�g>5g������F�T�ð �t����:����GbY����N:�Y!O�s0�p̮�;�F�����{�:��˵�x��[%�<}*���%���ya�a��.q������6�����ö#�V��б�䨐I��_'�]<����MK��E���c�ข'S���c]�~�q�I&�������¿�A�t�||r�������|:����������n�#�Ӏ=@����C5q�т�|�]�^��������K�+��3���V;���?\���=9nn�ڡ#;��L"�JNb�lJ�ʨ��s�N�6�����X�Z�J�ʲD�(/Ҹ�65i*΀鱐T�h�xV_��.�s�l=�0ď\~FB��yr���|�$x!u"��:�<| �Qo!YK"gt�2T�X�:0���2O���xA�֞g�m�@�{ڦLdh.�g��-7[���j�DCg&�P�-\Q�k�m���������T~�
G0-2#V�nr��20��t@
��G�wYY���h�%Y�D�~��3@,������;�QX�t�����)(TWEJ�8�Y�=�-y��,�A�Q�k����J�/+;��@������1J� @W�#��5!V�J��HE�$q��Ҹ(���$�fJL�,���u��<H��F��+
�ER��=R4v�y����A"Wb��s/�HX����mE�	��؆Ėt�.����v�cQ]���*�����̄	C$Óަ�*���V��%�[���e����@b��$Ϫ�y�!^��+��v:�������E�����o�`t�n�@ˈ���M;�Z�j��f����*����~�Hϱtm��'?2\�,_Z�u�r݀״EHA��Y?�u�!���=� ��h�Wwj~��3�0���B����Fĩ���;}��e��+@oB�<>W��|�n�Ԍ�CV��1���>���4}�P2�{�JM|�˙$�G[у:��phҊ�@�>�B����,����1���Sx�U� �Cx�V6�>�G""�2oTv�}|p.��az�}㰴�/
�D�";=wdY��Wm��35U����@�D��/���G�@.iw�x+Q\�3"p�W®P� �T��
P��Zo,LH�v���9	��UM�M���4i�u�6<�Í/�J��{Z���N���=�-�o��s=Ae�P�F*����f���($c�������)��L��W\wȍ�����-�[�k砺|�GҸ�q��(g�m�2xN�ӚȺ�/��2�}n��[f�(�:���6c>�h ?0sAF����+���U�4�k�@�v�>x9��� ܒ�"��&�2B{�w������
o^����ؠ�..�u�mU+��X� >İ~��R,D��hu�Kk+����v�B��5L}�,a�lj ����ݺ 2l� Wj$�ĂVF��༞��aK����m�k��%sx�7z%��-���^�t��{�Vs����r���J#�q�%�N�풌�Wz䩣�f��m��a��D�^D��B�h�Z��`����Qpdk���tZx�T�P�B�R�M�o��l�6����.W����ˈ�
��LnW	[�&��pd���h�>�-qK��^�oBw�;�2KtT!'g�T�C4⒃@	P���(�T*��k�)��y�<��թC4n�Ho`�����/!�G�`+<g!��} >�I
�ep�N�C��[�?
�yL;'?K��гOj�6+(�� K��eT޵��}Q�J2`q�`�6A�v��!8`�ӫN9A���(W���l$=��k��!�C�=�$� ���;���S$�.����s2B��Z {?�`\�4b���z)�E�8R��2��N.�������M�h���KB��Z7kD]|ƿ���4��뾤l��S�8�l����5��d�z������|����cD��Je�qp��u;��6�&�@%�G[pL����|�v������iO�I��vuT�mG�|�=zۧ����ԛF���"��ӥ��i��6L�a��,3=e�m�)c�+��fB���3Dc�mvE3Mɏ��^�T�n���朲v��U�Q�'�|T��Rk�jz����韞�{����E�툘#)`N��bԥ�Hiɱg���$k�>V{@��?����K�g�g�A6�VtԵ�7��N� z�<G���Q�,�B*@B�A�o��wG~�SSj���m`��8���:ĉ��2�!��TR�%�rJ�Y��pI���^4�?X��'W�L����5�&_��Y+\u�0��O?����fL\e�RO�܄+�zˋ�8԰� %<�p:�%�]a��p.���0��~�H�	��Ke���q�$Hh�|�ʓ��Ԇ1"y6M������y�J�>�J�Q4c< '����*nR�����d�~��ם S�9Q�H?-�����^�� E�ޓ�C����Ѿ�	�����TZ��^}	!2�%_���
�ʲ�:����i(�q� �Υ*qh��/"g�����ç�u#���� XQ����6N����3�k��8�_�F�Aԫ�,�O��$��'˲�@S�'�R���4����v%D�:ݝ���PЦJ�i,)�F���'%M.+���{�x?�v1�Hz��`f�Cb;�����n�,��ih�D�܆~c�6���*�dLTzbr�NzcZ����$���ȣ�6���7�pÆ	r�
�%Aq
���OСU,Nu�@�ý���!C7j|w7� F�c �/���Č�^�m�M���ʓ<y�::��R&˔����`\c��߲���p��YHH��J�?�[���K���&��˾�!������ےO�`�`v\�дMP6�1il�&������
��*�~�l�I_�+?;����yHG�; �3�"3Z��~�Lqv�؀�����Y=�XF����%'/����4ӝ#�ޱ�j��A�ω]������Y��]D���7��շb��� �O�i���b�$��˘I�c�XL��p!�n0� 0�z����s��b��]¸��ZdwI��$�°�5"��/yX��J�ڞ�T4<n��
�b[:"���O����ҚU���!�p�0��i�Ԉ$F���Ji{کg�FT�����<����=Q��N4d�|󖚩���=�q����dñ����lG����%��Q]H��A�^�@������s�S��ސ
~{�A���z~��~��7[��M�tї�r�=m�lJO̷C����ϛ�Y��G������XF�"��5Zj�ѽ���>�T^��}��q�=#+ܵX�~�fV-�z{m�qDWni~��~T��o�L.�eJ�o�b_�פ�H��<8s��6��z��X��XH~Zr������cdA���R60�;��X� ��*/_&�.�flx۲�*�HF=��yͅ���bN$���"�<�:Z(�|[��o���Km$���X��0�+�2�P���r;�������L¦�<Fh郇��	M7�l�dxD~���1�Q$��mˎ���p���<�])�T� gG� #Q]�r<h0d�����
*g�RU�Y�"Uhy���?�8~� �@��d����q'������t��O���)���E$A�t�JҨ*�gV�,������\�J�����@�[����c���1��@�>ݾ��V�<"���?f)�MQM�у�����L�7���F�Y�G�������5��zG!����=���"�e���ϸ0�%�m Θ	K��sgŖo�.���Ucl����/T̿�c$^���v��X[���3�v$���^䚕����v�E<&����x�f�1/ϐo�y�VE���Ju���n &}:Ƞ�;��R���f_G���r�>	~�h��ό'��I\��ZZr��״�8L�~Q��p���G;Ð�O�h�xj��׹����ȌbLF�_b�L�蠢�x�c^o�">2cG|u��'q�V�A�N���<s�4��F28�J㢇�����[��y�Ҙh��<@�LB��r��-���נ%e�s���{�Cx�5�"7�G�>K�TI(%��.�a���}���5�
p��"��d��lW�30��P�@Gn��k�e�0�i�VHx�58�.�Ȏ�9P�W�o��M���),��ӄ���9d1�U���٪A⯱ �PAQ<*�/Y+�ӂZ�O�	����R��X�v3A�o�Pol����f�r(�'D��+��t�Z�ھ��E:\Y��'���-z�u��M���@ғB��@�b/��2�fS���I�����H�w}I�A��k( �ͦ�p>8� �ԩs!}��lD�������4=��;�J�q�ҋ�;:�G-ܪ�/��mכ��뻋�\
�-�Ȥ�g��@����U�/,�P� �k�~��O�>|�#�}K�(
�l\Fv����p�^,?x�g���@��u�l��j�Ӧ�1���s��{߬��?��<#�~�x�
�z�:-��QəH�ؙd�Vn����j��Ur�#�ŀt��N˞���#h�D��f�����Ƶ�(~D�Q(B�4�Z�.}�ѫ���.k�/��+Ox`Q�P��RXe�JY��es�b#�.R;��<�������g�UW��
&�vGd4���e��>�U�q��qM���g�2�o�t�geT�C/��ޒ�PJ�(9=�*�)��0y�?;�3@�>�����`ѳ^��6
/�6H��4<�@���}ǴIe�"e+Cp�^�]�ֈ�
Z��LUT"?��A�vj�	(<�& f�?�-����Q�n�`SW�1`�v�q8n#�i:f��$��
l�S��fw�!,m/=�5�;��N���nX$#��o���n�B)Z 6�(ؚ7�گ�B���r)��8��-N�=mYZ���z��î&�앇�D�Ӳƺ�����;wᮤ p�����G\������������;���7;�������")ee|"/,iֺs�1�t&AG���[�ϟ�䐆Qo��j9����Ѡ��(��|��zV����]�����ǘ&ƣ���i���AX���Q�g�=@�,�d���?�f=�s���*�(#�3(�v�K�?^� ��'��vJvz���JF���TI�R��jU���!�9b�{�̫ʠf
�S��`i
8bO�#v豢]����>Q�Bʘ�1��l�g�)�6�c6t?�����WN�ʁ�t�*,���*~3�B��\��Evw�SN�����`m}8��{:?�e����f���mu��NPp���y�"?�ly�Lݻ��+��&ZbuY���un��?ͨ���\��O���+9�z&e�8����|7��� �5a6��p�2��7.�S�/H~���.ҡ#;��L�$�]�|�g����1}��M@���Lm��y��%�4�<�'L�!�%TRu��&�W��6���b�9��_HڟAƼF�^�w"  #��$�z,����7�0�T��4�YK	|�%U��%E�u�n��Y��?h�=E���*�CI��h���ߢ�>�xu��^�- �µ����6��+��k������"���b��GL,f���}��������B��-lG��Ko�g���f���dx+j�$4�a��N�M	={�O��4�v,bo`����C}��Bؗn]�w�����.�y��������%dg	�b��z>y���L����#���ڑ�f�|p�&Orf��%�8��*@�<�*Np����5�R��w�·F�!��j��_-^^����0#��h�<��r:��MR{A���lc�� �p��Hc�J�m��6'�31��m`�&�����W���.':O*0v;>!\8�Ҵ�1c6�Ci�z{��������J*���l��_`x>;���w�~H|� �U�"����Y�q����K��lt��G<X�>�3�'������4Y��y��e�A��]�������\U��Z5D9ZZ7I�z��b��� \�������<����I75�X���k-�n�4�0�q�� ��1��8���"d����g�5�m7�J2
�<'��yhYo# :���:}�i��['�!-M�}l��(�!�b�00�~����Fj	:m��{�8f��z$��ۘ���=<�S8��u��S9 ���mԚ$��\������2�ì	�H��'�����\�Uu]�+��Z͉����;]BQ^��.�MS�bݯY�~Vx���.[\`����ɒ����t��,r�P�G����l��3��Ƚ��P���slh����55������ٴ�^��g�?ˡ���T+��Ň��uV������k�ndx��ٍX�*laLI�sJ�|b:*U�@t�<��s�]�A���s�X(/�Z�g��4���ĸ:�@6+i��6�P�ʚ���_���.��cl�;i���F80�y(@A�Th`$�{R"�+:5��|�J�oM�$K������X��10�Ӝ2E���ҍ��LkN��� �=��5M�h��+��t7Qc�?��D�Iu���X��Q�}m�5-���~`8��T�wGf4>#L��r�v]0����
���-q�Y��h��:�~<��@����5?4	I���r�|�tOo#��)ެ@E�kMԏ���#*g�BȆ,Z|�����D�JN�d�S��v#�>m���1�="@��N��{�VKOp�ŋZ{W��	>��K���l�L b��Q�E����H�;9��U�tȰ������K""�P�J;��K���|s�m��	��hޖj5.b�aT�c�鎿�=c�o�����8$�J���U,ٳ��Ks��幂[C��p��=��+���������C�(d��+aEn�[�SD����nv;����[m�;�!ӗ`|.f:� ������~Ө�*��͝t\FZ���r�J��H��iɃk��Ң����'hBjt������)���'��F�5ާF��]Ƕ��do8^�>.D|N�S��^V�⦉�FX��>X4�&E2��sJ�#�A��Zm�[�;ժy�ahH#@�z�B��I�kNO�?0��(n�K���xg���=P�G{M���T�o�����.㛁a0!�}Yj�P�W
�3�"�
:d��W��l3+���X�9@����W��Q�i�xa:��)2��ѝPy��Êv� k ���,�����j�k�9��YUÎ���of�*��+��<e��/���fZ?=Đ�����#c����A���P
�&�힆fL֔(�K���Ƨ��ŗƵ�uϰ\�	��VV�-5D4��ӡ�r�e�n�^կM~�
kf2.���&���Q���;�}$�|ф(�'a���>�{C ��,s<ٔ��#'�����U��4�.��6�������"y�V����W\���!쨌�߭*�����
%��_m��r��k~jU�T���q t3x~�M�XL�� QK�EJ���v�²���qg�bV���+��0�kl�j�t�K�VI(�}�
C��#�Z�9�9x��zl�-r�/��)&�4m�Vi�g�8��yT#���H�N�o2�	
��j�f�r͙J�P���aD�~Bz!�Zg�i����k��:�*|xn�P/��RӜ�%@��g���l.M�mƗ_�J:����W�?!&�H.do
�� ��>ҝ�qaU�L���6���2��St�1Kg t�C*L�9�PX�(T��*�������y�b����>9С��0`��U����/�4���<�IӔ)�vp�I�{/e��y���Q7
5{(L���?�H��{�jP��(�R� ��['���PQ�J`���,��vmށ8�W7��[�7������Sf"lZ���a�T!���=����V���:���M$^N�
#�i�Bo�Y ��ص.0�*���m�z)<��8� q�(�N们(佃rO�^�4�̴����D�KƵi��U�2��;�&�IY��"�r�3H�2��}���������e@�Dj��q̎,��&ca��9�[�rK��갆,E��V��Ժ���c�,����|(:]z�*���ލ�_��3J�ɳ���5 �����73ފ�E=�ٟ�4�aΫf8F���f����3C�����^_���ل�pZvu"�;ŝ�T�RaGZj0�ݬ������{��)��]G�ɼ`�D�bʀ��7��%#�Z�l>L��xdJ�M���g�"6�;ftzZ��m�N�������_#�,�h*�FB���#rw}��SI���:��`(�8�2:�&���V�#�[��h+���{p��s���?NX��?L�Ƥ��&UQ2Y�Qu)Dy҆���^N}\�ŠO.��+�Vz�^8J��6}%��N����aqͮpd�m�����H9I��Iyf��,�'��$�r�|'$M��Tk1���M��+��@O�� ��4�\~'� �@�R�f�t����Ɲ֒]9�Hu2�Ʒ,^U �s[������t�z���k:
T���T��	ײ�%�0\�@Tǲ��;ʫ��߀<������}�*'?b��3��¹�eu���%i` ��R��/6�K�D�Bk��v�U%K��ؔ�!��,�'��(���M��,��]�⊨Ƣ^�����T�pó�A����C�|�����xM�ng�nL��H�v'
2�����k�C��>��n8�y��8<z���t)-��`�ՠ��d���bhZ�z/�Ј�A�w��$j�쿓�!i�p��|r�q�%���������� Nk���y�ըpim��w-�zF����������1^Y��魒'<�":0$	R�h� +���c����[�CpkO@H~��J��[��n�����&��Ծ@T����I�IO�s�\skɴ�316�O�i"OЅ�V��0� ��*�r�lFs�_���;����Ҡ�H�f� �")E��4�q�|h�A#]�
7��r,X�_4�.`�'%�8���.4I4���`�,AIZ�]��X� �V��p�z�|Dt@�7�W��w�bQq G^���a�X��_UIr&�X����fYbn���0n�]������N�d'��d�0���x=�5�}�e·#�T�-�*fՈ ��:ء�x�d�<�/Ґħ��_u! u0��ʂF�5�(��{���<������	<Ng�������[��������77T���T���ç,gʆ�����x\��@e]�c��� &ˆ6K�����,�Sӱ��W�~1[3��l(�ep��������ÌZt.�r��@�"F��-�п΄���AD�����T�k������5�R�3a��t��^�J��������J+�z�t�V��ٔ��짱�n_���4�ҽ��&Ld�J���b�¤{�����s� c��΂�XC6�Zh��[ ũ�.\���6&3Α�А�5]��_��.ol�S�`�F3�1y�<���$�Xm"��:( |�՞o�NK��CXP8�0 �d2��q����p�>;U�N���}�h_�S�3P�7�y%��D��z�!���Q��mA�F�5����+T/9<Gh�#G��r��0�F��{�
 �(��Y=q>h����5��~�C�@Ab��P���@���Y�?�t�xo��A�)9��E{�]ԪK�Ҟl0�Zx,�I�"�{��L�J��1lF���m;��"�kEQ1�q@(�x��NV��"+b�u�M�C����3<�PLL�������r��Ȭ',ê�\��0M8���J��ƴ�"hV�Ϝ�f	q���m�)]	������eI�.���sAc��D��׎J��5��$��2��T��������%��Gh�K���xј�{	��\��.�p��x�C�@�o{�EI��^�19"n	��Ŏ�-�;��ۗ�Nf���[	?�t�Z~�&��+��X�8\9�5Z��urn�h��x������f����/��Q��h(��j�/��6��d2:�eF�+���ߠ(Y4So�ٰ>��|��]�]lTVң[�'���*A4ΉK2.oFJ��N�|-���8[��L����h��@əBw�L�F���B�=�[�iC!�1
�x"�~�X�3G�כ���T����N5.޽Oa��}��k�
fۍ"̡�d
�qW>qw3&�\��I�@�+�
�KJE�ѓ�i(1-x�^��$�M�h�EP4ApåpM{����,,��N�G�X���9�U~���US⥢G�Qv<��/����O%Z�J�I�����߾�d�oA�bP����Ef�7(N�������j��Ɛz�Cx�\H�d��y���-����y^��\��IT�>����2�c��H�����>�}� �D(V�L��Dp>�4� p~�sWU��b#ڞ��ܐT 4Q@E�1�f�O�j�j�q衒=�h��C���a�H����f
�,"�h��X���U��"�	�l �~�(}=�\ؙ�hK��R�b��v~����b�.�]�����u���l.9�j�
/��Jđ?��:X��V�~=����x-�z��,-M>��+]�ϕ�Vd�c���˟O#)�j
$N�`��D`�z��f�yי����ul	D�B�-&ZBF&�G�h�"Uk���.�x֪8PJ_�RN� ����ɰ���.HUd��W)����KcWz��&�:%d�7V���W>��q\�׍����]��2�� tj�g���C%J�����P�5�(oG�*�	ݺy3�s�iu�4��Y��`Ge���/���ؕ<�ڔ��g9�Id�e�
@��g&��}
XL���?�F�j��(��) �a��@�}dAQQe`B
��'�v�R8�a�����S�ֹ�*��l��#�\�!�$=C?��q0l�D�{₌3$������d�`B�1Y �	��Efڥ���H)�)wu�8#-ö#}�N?{<�E�,t���R���z��\D.�'ư�����1�,[�Vӥ�����{a�n�
�5�4����ح�Ѱ�?�}��e���X�v�'�4&���<��[�5��	݆;dđGuo�X���чWO�k1|C�CzL�J����Lb�΍z��j������X�R̲�]�=�V��X}��|f3�F�D(Z���3^y	�A�/^:���R����vpl��f0�X�'T8�Rܙij/׬2�6�oK�{��C�Vu���˼`���bE�ﶱ�����>G���Ӧ
�-���g��E6u3�t�M6�^:N����M/Ν<�,5��*tzZB�"� "�wo�SDu`��&T`�b8���:5����TH�^J��$qco�j�Gpz���?��b��LSĩ�a�&P`+Y<slu���:��x9��\�Oɐ�+̀z�w8�QY6-/{Ŷ�a��pp��t�a��	�H�{�d@�p�|E$��~|� �����13g�M�p9�F�LڻDh��5�4��'�H��{TR+�/�r�q�,To���.9\H�2Ʋ2^��y v�/�!|�p#(�U�����T+���O��	2�%�,��[�Q�k^ʆ����B.ۿ�*�Z�`V�"|U�4�~u�;)`�G )�'��z�6_1,��,k�1��Б���Ԗ�\�,�;���Z�8��q�H�x G�#���9y�'L���	��><����CV��Y�D��M��c�����I}v"Ґp�БC����8S<në�ѭN��o�e�GS��[�3d�Ӕb��z���=s���㣋���G���1pǒr\Ue%�	��3g}�rVNfЃ��68�+���k�w��IF~�n��X�ܕ�^MQ�^�O�MF<���:���R��>�[�� c�}4��6�p&�YH�7�J|֫������h���c&�c�����|\�d�O /��G\�E��Uw6���i}C%�G����D{Sc*�l�X�_�q;Ǫ�-��Hxq� &�"����H>q'm�����"^�j�\Xw�m�I�'�y.�k��4�/Ì�yc[[LA�Ϭ]I�=�;���R�dU�4D�F@7%���b�� ��I������)��:m�I�7�X6��a��nA��0)���6���'w���d8b��dH���	3�3i5SцĀF�2@��/���Q�p�뎨i:3Ã�3Յ�W�z�,O�m�	!;�70f���/�F ���q{+��׷�i�y���GZ�<��-��Eg�	%e,����G��ɲ�8�"��h_�âoI�l\Н�s��$�K�!]��'��S��ņ1Y
ُथS(cn�O�1~^T�5�i��ݖ���H���~�Ft"��r
y<����h>�iכ���X�������K5���n����^�����GB�n�+-Ix��xV��o�+���B�nZ�~��`-����LR�JN\b�g ����rQ^s��������X^]TZ�Y6Ze���pO�6!���fp�@��:�_�K�.J��l)\r��:�F.Fyy�w���P$�UP"��:�׶|�o��PK?]��)�X	�0�2;��#ʁ·�ٸ��b����h7 �N#�7G�W��2D/�����
��Q5��m���PK��	a���?Tj�G��*#BRyrM��0��&�$8
�l���YYxHqhJ`�0�~��@�^��kG/�Wާ`�=!Ut��3��!)��*E6[r��ʢ�υ��z,�65���}t�J'Y����y��F��16�@��Z��A@VԂ��V���ڃ�b;��RS�LV��٭��qAx�f�Bl&�1�}� l>�e��]���=�"��?���ɸ�44�rp4m���	��D�X�`��.���ױWc��"���x�%�w�p��$/���s�i���������قQl��&Pdܳ h� =�F���Ƹb��^Ӆ���E$Q��ɘM�̺�n�&79���;�l�V��f���N��{g~Ɉбશ�*�\Tu�Zy�rI���1ɥ�O�3�a%��X�Ӑ��hCL-jj�P��5�����]J�F�A	�]�k�Ө_/�)o.uZ>�#�|�G�����V̈́�_'r�m6�4�Z2�U%Jtd
�����~�[�s�/��h�%�@07�B��{�!�ɑ}����d�2��`�x���s��GT6���T�]+��v�.��ya��}ϣf�& 
᢮"�X�dE�W�J�3!�:��x@xc!%,��\ͬ��icνx��\��z��_P�3���h�q��v,8)ڄ�Y�9u��U9
��*Z� K����<��/*�j���Z�w�:"��!�����??�AQJuP@���� fgY(	���]���"6�k��~AZ\������=�-����?C�h�4�$y]��� ��2������&�)ʹ��}�dcG#�(񔐦��,>I +��sr���B��^���>e4�qG�,[���o%"`��oI���o�\�Wv��C�|��
�[w�Ղ�37��a�U}���D� �" ~�#����TL�K��"���uvY��!���6ΎX��Q�ݦ6lI��jVՂ�q���U��L�� E����I��TxHDvzy�-(���JL(�j�V_W|��A����#D����N\q��Hj���f��� ���0>uDBpZ�Z���񌏽* k�����_vx��PeS�R�k���-�X��3`!.C��M�������*6W���&gL,d�?�6{j>ȍ3q�Oz��i�۪رL2�Ft@�?g6C ����I_P{3�(��R*�9,ݕs�yn	��@4/�E���=`�p�5�c/���y��<SV�_*Q"�Ivl�e\�����G��
��L`�?�i��ÑjD�(mp! �׉Qz>�X��Q��3`���"}�v#{�8L������-�(֔�(�d�l�W��W�:!=�n=��:̌|~ʿ���]K	$�b�@��_��B%�X gV���|$� �-�#��)�%8�y��]�N�Z��Y�G���T����p�F8Dɚ�ƫ�C������q��?���;���b!���"��qLȖ�h}��(�c���Me�\����e�"$�&�����[����W��P����
�6�������YbA|^�Rz�-3�[@�ԇ���i�(��A>�z��r}�m�ϊ��9=��J�@��K�f.j:��	��Y�|3y��^��Z��R��vkٴ��%�+�TS�hRWj���m�x�
�d{{�ʱ�!����`�9b����\f�S)���0>B���.	����<vg��46PK�t�`	̣�oNט䁨�L��t�,P/*�͛By�O�[@�w�TcS?Ţ��K`�hQ8ָ:�CM��ʉ�9��uF^Ӟ�Ř�p5]����?Də���L��@��c�&K�`Y��Gu��.U���
S��\Q$?Od��+�z7��8���lU���ő�^a�A'p����&�dP.H�r�'��:��ݕ�$4��|]�f��T�1���Mq��ab8�6Z����4O��'�A��nR��.�׏��.�꧴䝌RP9=�QH��oƭX�^�5 1uh�<$L���Ǿ0����T�<"�J��	��(%KH6�vZ��T��aK^Uc���֢ۺ��*ݕt����=��¯��u���a� ĝ4��R6�����:�k���K����hԗ�,7�`�֬��P��,�}��T����@4�b�5צ�ȳ�[�<���U�m��OY����M�2p� �m���v��qW=�L�aC�#u���n���U�S���joZ��e}�=!d��-b^�tz�pD�x6L�w��� �ڢ����p/ǐr�X#%�|c�n5����Na=�/���0��V�w#N%FY��2��0�!^aՑ��V�<��:&7R�uŔ���PO}c~\���p�B7H��YJ����"?���>�S&��M��?�����ˠO�^��:�\�?����56�bi�Wz�v�?0���*]�5l�]l_1�;zh���MH3�� A|�"���꼙qb}Ȁw2�� -��&�X2���d6'���F��4�JK�J��V1HA�d#](��V1Q��0[\D�la7d~��b�u ������+�N�"��QI�h�X���\�n��/0���Q����hf�Ʌ��d�J�	@.J�5�Tě�­|]�
lG ���V뉪&:����A��r�-҆�b�H-�!v�J01�����F{��i�{F���2�ަT�䂷�<����ݦ�d�W �B��}��ĺ��M�]z}��Ý�2/r�X�A�㳪��]�3���ZR���,�8bƃ�_>vSC�ʞl~��pI-�B���ɣ���9��t=Drr�wD���̣�?��	���9��S���Z�Ğ�#<5ƍ�ѩi>ધ�^�H��P���),�+H���j&lV��Քf8�ݞ@nU&Ρ��g�[Z^L��J}-nb�6n�񻮗C[s�Ǻ�R���D�Xy�VZ^ߤ��OyǸ��6ٚ�GV0��ʴU3#_��.%�}ld�Ė�F)}y9/�9/$�r�"}~�:Ƨ�|GL�o�*K	�}��nX��06��2����c������tV���:�F>�hղ0�i7����;Dj�B�W���Q�4Im��f�k))���ɬT���G7/�#=9�r�i�0PJ���
Y����pY�?xh�>e�+ǖ~M�@�{d����z��ނ��x#t �o���)E����i�ҔQg��݋,D�X�~�x�OJ_T,�@��a��}F��!�1q&�@^����TV\F#����z��9�ض=c��v�L�{�ԋiVp3i�]�q��5���yۃ��S�Ӽ�U"���{Vz�����im�b	7ڙ�)��[�.s���c�+)��E� �̫�$�M.�Ȳq��}�|����Ղ̰�$���OϱVJ�P���Y��B�y�2�ezE�����}�g\!n������Ȍ�;���ѫ1f�.L�ѳ[���~�(�;J��δ�\oWZ��Ar$i��l9���o}�\�"ҳ�Y���h^Oj��z������,�F�wN޸�W��I�J��o�0�>�N�|���ԓ��Vȅ���G��(b�4�p2$\JO:V��/�+7R[�?���?}hyܮ@K��Bm���p����t��3�_Q�����x�_��[�G��y
�T5+���.�a aA��}�p���
\�;"�/�d��FWtD�3���i�@3��@{L��U͇w�i��bx2���C�W�P�����+q���[��,s�}y�T�9��U�wq�E�������<��/�/��K8ZP�&���<����:��lA�(�P�Bf��I�f]��(�v�0X��`���F�l�*�\~�l���g��-fI��%P��������Q�������2?��𾓯�Ae��4��}���"�(�{,���E>�3 �s����X���9���I�4����'�s�����Y��y�3�%�J��Yl��~ ��w3�
6��Ȑ��Nɽ�ܞ�UX��� EJ~~>��g=�dK�\��Xv4�ƴ\�.��E�S�x���b�aT�ld��j��g��L���]�����]�4��j0�xc�cz�/P-*+Ʌ���G^VZӰ�I��AM2#_�P`�gN7�J���(䰅uf�矙[�q��/�D)60B��Z����H��Xik��g�;�CxL�CP�g�RD5�t���.��	�.>��ƨ0��{����)�Wp��&B~Cd �<�я>�5Aq�<�}����Sߓ2[#Jt{:gђ�Cn�JP6QB(���*��p�Ey�����*s**b���`����Pw�/����T�<��E��2+�IєVeR �ʝ���30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�-ڜ4�{^��T�b/s�C�5}��lO��e5��G���'�}�0�|�b�3��0�t3w*2�E����'��q6�����d@nw�	U;JS���-�a�F"N�H1-2-����w��3� ���4d�[*P��
�c���d�{�k���(z(�l�GSިp�Κ�
�c����R���Evt躴=2>"~\arpꕶ�"�>Ea��bʒ����=���h�Ļ�z\���R?R��m�4��[>� �e|��|�}�L�q�y�*	H,�&�ԙ���%���#sк�l^br��$��*����~T���bQno�^nmXwV0��8* by�(�<��$��5,�z��� �w{�_|�I���Bx�Q�� !&�\�)�ݧQ�i����S"�?��6Qw;����#﬿�9++�,e,���k���F��"K��8'���J�����4��
rӐK������vJ]�Q2�wl9+��x�ii�B�l�}�F�(Ḇ�,�e�vN�7����M���I���K��_�]�5$Nu�3Or`��#	@��SI�*
�h�z ���Rˬ�u����*�����,�:"D?�Ϝ��\'�Yu��:���G�Fڍ�O^o%�
��~0~gA�<�k��r��\�}r+�O�"TH�\��س��¤)@F�'k�\>G=���4v͌���a��{j)�0n߬��(oqz�(�d��X��U�{�/��^7������:���?Y��yU��q��&�H��G�D�5ɐ��K�&�5j!��K1��s�ˢ�"?����^p��o��8IMj�m�Ϲ{0|O�?ă2������R�n
�	�~�HI'>��6�RBiĥAiazZV��o5�^�=X%üؑL��᲍cx5
���k��sl�����@�/0���O�m�x�D�_;�k[���FG��F�|��4En��9�xc�e�՜
�]�i��Ҵ��1�E��
�����SV��FԠ��e�8A7��`�Dp9�GM�,s]M�	>vU$��q"V�7���@m�̮,}���%L׾;����ۆ�<(�{*8��h>Tp�7�3J��ӻU��j��L$k�
p�I�7��
��t�V��0�|.oX[M%���KQ���[N��`=R��r���"��:�	��*��ȩr�E�!'
~��ć��6�:�/)���GL���Y�V��k�C�������b�Z��a�>"�����9Z��&��y'.�C.�O�S�aG?�6��3gR$��s$;e�<�y���.N��i g�_�o�H�����Y;���n^�Lp�LDN�	=VV;&H�m>�3�g�w9�~�+~s�����'��q�����括�Cd_p�IT�K������Sܾ�����1]�`�.�jA�6�
وɕ z�1���{ġ�>�.��mfZ-Voͮ�<ؐ��V�������@ޥ�~�7�5�9VW�;q�h�H؇�;W��Ql��c("�G�w����}~���0/>�a�/՚uBQO��N
����N�}I�aB|�O`�N�\*WLآ�
(o���ŭ;��:'d���s�Wi>\h���<G�*��1�6�ld�d8	V=��>��4��
�?EX?1�UvK5	��<|,*���߾�<�a*�����9(1�P�^��Z���]������cn&Ú8Ajw=g]��"�	fL�rb��S�H��қ��q�'ע���s�Vǻ@=rRh
ף�O�z�#1�̐��팩"�CR�ľ���P��c�`�ZV��:qAq��g^��,=s<&����s���b��}�k�F��s�6tF&zL���8_j4W��7�r�!�1�sb����MŎ�Є�)cM�����x��M���\�t{q\�S�%L���-WMT]h�dl_'���'-������U�?�r���0���4�6U�r'�<|,�5�y�I��q�n���g4B�uً�(�b��!�������ʅ}�jF õӄM4R��3�jI�ܨ��ݿ�s�l�<Q��6M��IU�i� ۳DD`28�-�d2����~�e�7X�O�5P��z�����WBYv�#d����z;j����=�)p�>ҴB�z�D�T5`-�E;O�?��o���ȧ��B���� ,��i둀*;,���*,A�ީ.T�@"��|�8W��Ri�ޮ2�;�|��ʉCDK�D�����X�Ұd���'1�TP����Cu��� ������T�:t���^�P�Yul���V�A�dq��t�t:  3�a�����A������x�⬪��t=K�:�S[��D?��%?q�_���a�OI����=���В����{��h֖��iu�r^��x�ƪ�ѷz��.ȣ�+�"�v���nT�%��^��iC�4�pG녏�(��Hb�YBI����0�>��/�F�[�Y���ls�X	���,Jp���ߠ?�	���N��WNJ@�W�V�&_�^��*�P�o�w��T$����׍$�@���|]�f���J���●�
e�eJ!�E�M	�\_Y��Yۤ��bԻ���a�j/��C(�z�q��d2.i��I�$^6���w1{����_��q��PIC��9�.��KBE�LnJ��P��sV6LK�/4�&X������K����g&���\��%��f��mXk~O}٨7�d��IhƲ��]�%�%�l�he�����6�`�P�I�S̊���v�Ĕ�c�";��-_��}ƃA��Q��Y�͍�ٺmǚ���%8��ə��[��}5�Ff F��g��!�e`!��s�*�$��钴~�fķ3KT�x9�ʗ�y����aWrE�\48���ğ����S�'+�:s�K�R����N�P���ˀ����R��u_I�^��,g���豳���,:'�����t�e��~g��*l��y���|�Ml�AH23~t��i>�]���c`h��J/xS�A�9{����/ ��w���o	+�?Χ]c��o����{�رb(4�ɛ�y.!����m�H7,�9���36[�(z5�M�A��g��Ł݂��cc�Q����]`��p����1�#y>P����� �S�O�3�:������� H5�=��!T�q`>�&�E��j݉Pܣ<��".-n��M26�I�Ps�|���9{2=�CHY��vX���o6���e�Hd�GgSѻ��!1P���o��cJT�����5�]���|�W�)��^+m"��؁Df���ˆ�]y�6"��/�i.t75=1��@a�ϴO�"G�Ԛ��ɚDi+�et�7B<d�}�Gn�Ȟc�������DO�v�\֯b�����bU^��^1Ҩ�V ��]I b�I��ǟ^��:��!Ń��a���^�=x��2�ϙt��� o�pA��=��s���e��E�Oa��H�k�N�*����5�RZ�3���ņ�bvX�i-�h_P��r2 m&�R*kٷw-�d�����-�]U} ��hg*՘Ӡy���#\M�k}�/�Od�:T�K��w�6��ӊ)It��PZ2\��v���>(�5奶*�8dTW) Xmn��q|�z�B�DeM�q_���E�gW�����Wı��W3<y���U�8��%`�Q�:p%��J352����E��ԸjꔩK���|顢vׯ�_���1����*8��jR"RϢɎ|X$.΃h��#O�G�;�]��c�	k�HH2Nܑ�:<Rk����2ui��Vs�W5DP�����Uɢ�
Q�c��D�S�MkV�l[tg�v�)��0�ۄO�$�x�0�`Uk��,�tjýn��|��HEw�2�B	�x��'�>
n�~i����}Dճ1�E��w
֙i��b�-8z��ם��B�7���MQj�pO*,�cJM$8�ǳ�$���q�巰t*��O���:,��юէ�ĭh��:�Q�Q�d@����>}�uˀZ�J q�D�w���p�Z�k��P�RY6�Xw�8�\�P�זX�j%��r�4C�f|�;�m�prw����Q�:��w�>v��ir Œj��~ �X�k�H��c:����vL���낒�	T�p�݇�.���_�١|�C�a�b"�����9�@�&��D��~O�FaP�A�_Ow3�a'�l�;��<�08i��n� pp��R�H�ӱ�`��;������_��L-,J�eV77)H;�{m������9rg���{W�kWO��eښ��Q���������pM���N����'tS�n��"-�������*��A�P���A�ɞ���Z�b��9�g�����m{V8���%��Ո��ON���_��3���V�8�;Z��h�������\}3QՅ����G(�7�$޴�z}����Y�İ�c��6�B������
�C��l}R
B��tO��N9vhW�cM�K4
�4to�-�����vd*-�Y��W�(�\�{����*�1̒�4I�d��5	|!��Xw��6:��8W.�F1-Hvt+F_�т����I����Otn�J[5�����T���
�ːN�B]|�Zn�(�lX&����=��ժ3�X	a�r+��S|+������p=��l����@��?r�b׌����##Zh�ٙ���1����g>��1�P�=��i4Z��̃I�q �<^jݝ=_�&�h����ƙ���ަ��k�Wr�(3s�Pnt��@&C���8h��W�/΀�Pj!żs�݀�\���W*���I�M¦4���р��8�IK��zq�B��Ki��&�M]s+
<���-'��-������?�D���	�,ɿ4��Uz'f��,.�yO~=��cwל�9#@4�p��h��@��&͎Z&H�NU��*FI�u�ʹ�R�"�����Q������s{uQ�EKF�_��蒺��i��<e`�� -���n
���~��`��蘯	��7z6��k�7B"� #M�"�
Σzd��O����]C��8��4B���-��T>E��n�����~#�o
/�d��R�� gi�oo*d�e��JAY�.ݝ|�-��E"W�li��*�[��;-w[�:1@C�~DX���y�vۻ#J��T'Z�bP������C�I7����^��T�����^C�MP��3uթ���
BAB;������]_�(��.d �f����CM�x�RѪm'&I�C�2[!���;/%k	��+�
șI���,�ၚ�����-���>8�uw^�Ʌ����6��A׵E�TbKR��q^���P�h�u ܥ⊆'AM,��0�)�(�mSQ��l�Q`���>1��C/x� ��kO�C5�n�[�ʖsFF%�q��1�oMI1x���Rf����O�շ>�x��$�u���^���z����q�i���>"B��������4�^(G�C7�Lp{֣�Oz��|��Y��?���]03����V��Ģ����� 9�Rԝݬ�PJ�W.�� oDY)��\��*$J��Wو�Vjx�_���ކ��
wYq^$�������l⓵�mp_}��d,�ұ?���L9j����l,���4=���݀^���'�91�~[��'�ɊnHq{|p�h������WP�ب���)�. ���
H�|���-�e��1$:���.�  b�-E��޲-�~J��zǓ`[�i{����쎿Ц2�NU��a%~H}.Kz?u��1zc���+a�+��Ft��{��n�̲��h��X��+�7�~b�[��A�yq�|f���E��*.�Y�[I������!s֣ �
�{�z�|,�.�%��B�@F�S_tcB�;�d)�\{�e� @t(͛"��{JU(�֖"����ƭ��'~�yp�+����cUKv���'8Z�&�u/CP������*Gz�~��$�cL9<�8]>a/�x�4��;�+E���	u�k����<+g�ᕩ�έ���,�����s�*	��N������:Z1�=z`��x��q�{� ��SD�.��B/=��t��|�h�Z-5ߞ�c������	�з�����7�Z�J�P+�Aq�(�ĂC�[�C��gy���̷
��Jf��2��\���ջ��\z��SΗ�CĜE�^Į(�$�q"�w2S |�ҡ+I*9�6τe���|�_�t�q��2��\|C���KG�L���z�X*�ћ/Y�X�[���/iK �����ɽ\���%��Zf�h�X0��}>|��i*IL���֓
Ͻ%v'��=s �V��� ��U:!���P�!��[���K�c���  o-�\W��pn��4Q�������?�Q�7��>�.,	�`��}ڸfe������٦�z�+ƫ��Q*������Ҵ�;f	��K9_�x�lO��ز���R�;p����XV,�ﲾm7k��wڠ��T����2�J��|M��5��GBmڞ�2+ׂ?��>��G��.�I���k�_<uF��m��T^<u`�G���L�G��Dn��=e!4���xT'��f��8P�Ż+7�o��HTT!cT
f�=M�r�r7���`���b���'�T��B#� `yX�{�;����쵀�kM�j�h��դ��"#v~�e-B+�㹩���Vb�H�Bf�?V�ʞ�e��Eτ�"���X��N�a�32�h`��L�Jb��ɁI�`Û+�Z ����A���.u�1˶��9��q�͏e:�Y˙�j����<uD	:K$*G�4F=*EO!���-����g$�Q>N�ԋ\}�}�ztO�L/Tk=�1���W)����x�\A	�p���˂Xͯ�޶��^��):)9n��V�+��z޸|ƪ����ŵ���fȡ��@��yJ��	�m����U}�W�k�݋��ѮG��5,�=�X�I.Zj�vK/Bݶ�����������>O�2=8l@�jŐϜá|�]�H�!Ć�4�AaϷ� 缑p�	%�sH,�^��	R�(3Ĩ��iĮ3V��o5�7��U�j+��6�քeCc{<v�M��kE��l�5��g�#�70���O+xО��ջkb����(��|�uE��놼�gxf���8�5
�W�i!Z�7it��	E�s
P<����V��SN�'!҇�q7���&����\,vo�M�b��$(��q�>m����͉��o w,���ш�S��)��<>�,I�^
w�T̓>����:�vJ����~���;h(���`k�v������bu�w���Ve��?��X=��%Dz\�.�a�F�j��h������[�r����E�^:;r�H�A^vrz�:$Q~ꇥ{9MZ:skϟ�6�L�8"��*ߔհ��j(��ڬI�.�w�[q2=q�a��"j����c�9�9K&��x+d��O�e�a����ٛP3j=*���;(ȵ<*w�r��Ӯ| ���PydH����ZX;�ڡ���Ս��ML'ƂL��V�7�H��"m��o�*�)9�ۢ���eK�//��r*��>����Uhp�R{��"��-��4�S����U'I�#�����&A��ɀ��{��Mϊ�e��~��a�D��m�IV����/�,Z��	Ƈ�[��A���X�V���;Tfh7�퇊���Q�NV�ҟK(*����}��0�}�hϾ��İd���XB���V
�<�+R}��B�OcҹN3�iW�~���V
�G]oޗ����q�d��t�S�W��|\��R/���1�I��d��V	vR+���[�W�J��r(��1E
Pv�I�E��+v���R�	�٣D��4bm�4}�JU���Dv�ț�]6;�hv�i�&f��D�=�$g�m�	�F�r�=#SvW��Y�)���Y�*�X��X��@4|r�y�׆ℽh�#�T�̓.��$��:I���hv�IP������Z�H��=�q�#�^�ɓ=�҂&�K���%���� =mk���ϱs���t5&�	���8��FWO���u|!�s%�+����A7,M�S��h0����m��7Kwq��ڨ|}��n5M���j�b�q�#'�Iv��GڀYo?��R���u��ѧ4�,xU��'��u,�� y	����r�R�³�4E3����(�%=�D�K�������FáCӇ ~R���-���K�`<su%���'����L �̆�vן`U#�-]���h�����d�R/�vqzpsf�嵪Bܘ�#GӵD�`z�6o�	9��.��(a��B��B�'��Tx�����V�B�	�xNK�����ކ���" �i.��*��蜼|-ASq�.�Ic����+�W��i%���}o;�^%�4GC=�D�:��3۵�;��'�z�P���� �dC8�)�CFV�5�T���d^�`�P��9u�<p��=A�ts�2��W��bA��ʎ� F.��l�}��xfª'�: #��}�1[�1�B�Y%eP��"�(���;I��x�����5Ԓx5c�[��'-��x��u�ۙ^[�����#��t�XqS��"����P҉�Hy�^w�Cf�bp�x}�>^��KL�Y�2V�i�G0�(@�Cc�)�템�w��y�!���[��J3��c#��e��x+��
�J��W��>V��_���M��#I>w���$�A�ýTl���{�5h(��q���Ȫ��J؞��P��_Y��԰>����J�"��̙h�I0����5kQ!��q.���r�Eژ���Ӎ�wXK�n%2�H)���(��A���C$r��$�S5:	�v7���Qr����E~��z��áG��:A�a�kD�L;���
�=��{ε�L��(c��<% �)���,�ai�Z"x����9K�&�
9���O��a�(���38���?8;vZ< ��@AV�a� ���^��H]^���;�^�	�2��CLL��J�(rV���H�'�m/}��xI�9�Lp�|P��Z}��"���K�|���T1�pո���J�4�����S�^g�rV)��\�q/��zAm���{���&���PX�L䍡��B�?Obm�"V��9���v�}Fu:s�� �1����u�f!VT�m;�6$h�9q��>��7�Q]�;� 4�(8������
S}t���R�2&7ՋIBb�c��M
`
��C��}ڒCB-K�O1�=N��nW&���Q�
h�ol�+V�k��Ud��߅�	�W+�o\��_� ���N1T+����dt��	M���7�ed��[R�_�1��tv��碨�-�2�c�۾�Z����Ђ���B���ɹA?���e���]��c���@&t�I��=X)O��z�	���r���S�����|��7�u��g�@B
�r����[���X#�9��a�(�}�D�T� ��D8�P,���\Z\�TXq�2[^����a�QW;\cE�9�9[og�����\��O�qz����.[Hh�"���ʪ��`* �V�-�K��Ȼ�bC[���!*	�*?��K�b���oj��new'����
e*1�1�Ydf<���4������^�;wLU�|�[��	�M���Q/��lZ��u�)��:"�R��"�d�8?�lUQd�.����#�N����Y+zvn,��E� n%����sX��8��$�Y�+���{�S}Mi�<cg�zZF��8� ]U^)�\O)\��!3s����J������֒{��(�`'��,2)���G�\�CWӐ�zd��P��5߫��" 1��p�y��b�:z�(��D����x�~�3]�!F0�1C������f��� 
m��36*��YyF��+@��X�c�w2�C��X�A3͂���J����w�k�m3��k�Ǡ����Q4%2�䑑VD��>�ہoUm��.2�?�	
>w�G����� ���h_� wBZ!��v�TZz�u�"�G���L{�ę@�ع�Q!0I]��T�����4���79Q�k�Nİ'!_@IfF�i�n�dr��y�\W��ޟ������ʸ�>K��|�T�ީ����Ų:��h�M��|�r�ՠ�*��zQ�-����߻��8pb��GC�HG�C�[���ϧP ����ǯ{��0�*fbs�V���.t�
��1������ç@�X��q_�t�@��2�mbJ���CNVa�sN��-#�w܋}��~Z���[�U�ڿ��c�y�d��kA���˶(LlVG7ʙp[7���cG��6҉�o?�t�H=�a~@��pi�|���It�a�Ѱ��1�����=!��L��(l��ŭ͝<�R��ʾ�/��i�\Di{^�$iV�Ep�%��i7�"��q���7�[I9$���R�C����dlO~2�db�&�6[Ft�8�B<���=x��Z�~n-�cA8���f
�a����Ey��87PU{Q[G�$l���B�RS���4c��*�j"����F�2�G��	�n�hjF�{wo��v���.U A]2z|���h�D����@n ��\��L�;Ǘ�Yp�ڵA�E�Y8�&c9�?�1W|��-��"��/G]�'Y�M�+@�(�3yC�4����v�!���ڢ�t@�����03�3t��󅶦D�Q�ѵ$N���@��he�}�k	�1L���S{�Y�,�Ұ��&$F�h}��Pfh��8���|�[b�7�EK�/v�7H�c�T���͑9x�=�ŮЂ`�������5̆�eQ��N�m��Ł1��1�0�+��j��!�b**���wNŽ�3r�M`h�?�FI)e �k�8 �A큮(�%S�u�������-��E�:%&��2�+��y�à�uY0[:���GNвF}��Oa���m��A�(gdW7Mj�U�k\G��}?Oޘ�T�1�qm��)�1�
m\\������W��Į�$�]�
)z�#n���k@9zQ"����G̶���2B�����_��u��ݍ����P3�U��Z�)��/!*�O��k5lpܢN�0��j�y�KT)���v���M��1ҮC��r�,8�T�jLa����H|�	,�#��O\健�������	e��Hl�0��R%�D��i3sV�5�� r|���b����c�x�dSk��l
b���c��0OYOk�x���k^���.�h�V|�'�E�J��*x�<��x.V
�#�iOu��wE�TQ2E�
�����:���_��Z���ǝ67ų��R�*�,��EM^A�$h�sqȚ��<�s��º�*,�!��ȶ��>��|R��K�>�. ��yQ>7	y�zV`J:��Ӿg��{����Nk����շ��������<��X}`�%����n;K��ψ�>��5<:�zr�D�х��:{ί������r�w�d�C~Z,���ya.:�&�[�L-��<_#�me��l�y��n�;ٛM�}� a[�"�sO�`i9���& �k���,�O�	�aʹE�P�3�ye�V��;h�<R���?���g � �m�H�E��\N;gE�;���Lg�-�]�V�k�H5a�m���j��9,i��Ã��Bo��T�?�K��.���Fap簢?��}�aS�Uq��3rg��c1���A�=*�-������Z���Ρ�舎1#lm�]fV2=�_@�o�Kl���I�����D��o�V�پ;�o�hw����k�VqQӚ�� (j�.�
ƴ���}�о�밤K��=�BT�ԡB*�
Ҙ���?}̅LB_��O�NONs��Wd���
���o��Hf黱�d$�⅓?W�J\�k���l�MRc1F£��g$d���	��p���Q՗"�͛hr�1�6�v.d1Y$���pO�z�I1�U�β��:kbo���\zt�=/p);=�Ƽ��q����7 �0�`S�l����(�RBh�3oͳ�n�X�J�o��l)�P�̟�? U�)R#��_�!d�T$e�$�@Ғ�8w��k�Ϥ�����0W)�yxz6:j&��j�U*޲���nZ�m��i�����M��628 �d�:��'�`��������?;��о��Tm�4!>U*_'��&,V��yw����>��>�ao14�Ҋ����pT��FX��K7�)��wFq�d��-�R��
�y���pzs����m���$��۴���X�d&�`P�-�v��$쵯�F���*��x���;z^�ٓ��BJ�#uoA�2՚z���wo���Əړ{l�B
e�Uc�Tf�&�U{��.���aJ�����z�E =yziǟ*���*p�A�ғ.I�>��m&WQ>i�3����;U࠺b�2C��`D�m�����ㅧ�h^'�T�P��.��C&E���F���K�T������^k�P��6u�� ���AjCC��ց���P���V@��q���wt�k��x�����N��k3.[Iuj�D�%�7�����2 �I�L���H�	�6�&G�L�Ubٖf��u��^��������Q�$��"q��>����;^���C��px(6��q���hY���W��0P������WX_��� ƽ:����݉��J!�������1��֌J� W(�VG�b_m���8���Uw�$���kl�l ύ_�WdI22�ѡ>�m��9g�t�0�li��X�7�9ݝj�Ɣ�h'ԍ9.�s~���d�e�Kv��e�݁�Ƙ4p��$oإ����� �i�������eM�<$`Fퟭ�.��� ��E�ڲ��g��z���[�Wa��ͷ�;橿Ԭ�+*��ޕ8H��Sz���ߎu���M�+�ڀ��`r�����S����%�LX.�T�4��b�<��0IyN�|fy|�E��.��^}��T�Z��s����n&{!r�|3!.��nEeE@C4�_�4�xٜ)le@{
�x ](��XZ���y�U%�S���׈����J���y���w�L�V<�UH>VdB'uU&��m/���������$G�G��i� a�<N�/]��,/$�4�������^�	r�`ʕ2�<h�w�r�o�*�2���{�\��D 		V4N-t��2 lZ��e�����s�O���!��1?PvP˟$ì<i�^�|CZb�p��g�2(ظ�T�Y�I&���0��q���q��[����Ѳ�OaJ��w����@1�˝a�c��J���W�Vq_�Xi�AԜ��bw|��$g90ñ:�l%�*����_���d��}��K��3��9�'��v�0loHl`����Ej���(ƚ4'�$H9�6x~>jwj�*���~"I#�uƞ*[�z۸�+q��k^ �����H���dF�eS9�$&8%�%c�.�$� �4EL&�0q��	z��[����`����2п�����d�qH୲z�3�T^��LOz+D:��Q������`x��|+"�X�;����b�T��6j0y6f���ER��.�;�~�i��栤Ss_���{��|y��.��w�i@ɧ__Wuʈ~F�)2s�{�P ��\�^ں����U�t��f�$�P���`*�>y���}���#�U��;��'{��&Fr/F�p��f��ݻmG����N��F��<Tk]�-�/�\�4N)��5�$ȵ	��D�ۮ�<n��8�%ΰ9��0D�������]�	��Ns���8ˠZ�0�@�?��U�{�!��&��^����&=X�Y�hQ��5������/����J������C?�i��J��$+�ͽ�k��&>�R)�
(J��Oem�J)7�U�\g����������j������r���!'r(��,q���260����I�ͦ6ҭF<����_��q$~����~Cȼ�6*�KJ�ALv�|�XD�{˼Ta/<`X�������Ks[�o0�d�\��%4f�0Xs�]}���lL�Ip�0����-V�%��� O���Y
�>a��X��[�˲�Yv~�9Ĝ�>c���C�-�����8uI�Qŕo��"��£�� y-*��rd�c�}=4Mf(�����)~
h�R���l*#!}��k��A�f���K\��xA$1�ր����a_[R�d>�8�g�!��ħ&��!?�/�+�Bw�坼�R�v��!�����݀+���R��_Q��^㽺g����]�\,B���t��ĕ�ig�X�l��x��!X�U1�AP��;)�t���F�e���k�}�#_/���A�'!��x>7�Ӓ���!�3�sί���D��� ����(<+�ɣ�i6[Ӡ�7m�$�,��{� ��6"`(�ՎM��a�obd̈́f��Dc�6��㍰�e���x������+�4P��Ղ�����ߔW�3�	���e�����(��E��!\k2`F���M:�j��ܫt��*g�n�r�M
�v6�	!�X�J������{�C�K	8�Y���6%�m"�Hl�0g[8��j�1X��wi8k�=�'��]�9���ѯ�1yյf�|"���#w��΁Sˎ�]��z"�.�/+s.|aN7=������:O������n��ȿDq�e|�x7"�<l��O�Ȧ0��kY��?�D���~��ַ���XJ�j�k������V/��e9tb�:q�ϱn�HM���!���T�����E?�:��|B��(	wpI�P=�(��I�����W���P�s���2�����Rb��3��oŎj
���p���� uGR2�T���d�p)�_ͬ`vO�X�F��F���񲶖0wa�y��%:����.�QCiK>	�~����fgY��y�\Ǿ�M�K%&��4��S	�CT���c��=@kWn�7�=`��AZSJ��ؗ����wd)��-�wTn���`����;�Q �U�e�ܛ�݃-+�������Z��r��fͺ���T�7R�k�m��F 5�{egl	��Y��혷�"��T��t�2|��w_v��t���nqY�ρ�����z&t�гTX�2Q7��G�욞n�o�SN�C�t���j�5��f�i����|;@Vu�zF��!�V��T
�KD]��D1��=RZ�`����"�i������.Z/��gv�yf��/o���!��"yv����4V���|�X�ado��t!'��w� hEvI�
��|�>�!y�������֜��7��IzDz��0��o��BK#�ĉ$3��ְ�M������� l0�;�щ#ݐ~��	Iuu`04�C����>n��0O>�U8e2F!�Z���ܣk0�'�VnM�9���̓,���2��5cX OҊD�G��O5�Rq�;p��Η����g7��e�)}�h�8x��oUr�����0V�v�B�U�j�>8���"+ñ�T��5̓:ځ�U�����>4�#��eP�@�oO5�x�9n�N�#����&�bxqe�v� fT�.����*��r�czA��F���,e$��*�b�7�߼6���?$�y��"���W��[n�,L~X�m*Ŋ?��D�p㑠��W�n`���XL����Jޮ�c���K�C�g^�V^�q)��jF�M�NC��
��'ó��$�lO{�i[ �d���]�/�?x1�)E��!�(��Fd�J� ~�%A�l��|��Y��Z�:�;!��a�V���$�̰��ƞ-�՝�(m��Z+�U��|	l-6�A�[�����6/4�*�嬂���3�G8A��{��B�6괯�\Y���F0Vg%����*�o��)�
G��]��SrW��"j[���\�x������ JwT?�4Yh��U	��[�����I�?Hlc��5�Zvu�h=���������Y�G��f-����5s^��1%t��[Z:��[�����F�'"<y���fs���-*�=��4�4�}�a7[�������������'`C�§�!*f��B�v�����2��o�.p��D3:o�ÑGĬ��v^�[0��Xާ�?��c�q�@��B�H���΀ԋ{�A��W���lZ�	�b����5�*���@��,һb�t.o�3�n_y�w��d�y�*�?���<Ƞ�5�h�,{P��=hw�h�|_� ɪm�j��Q�
;�Ĥ��h)��z����Kt��$?��QE����#�7�+ �+�+�,#3ޡ����P��T�GYү8�C��_�+tz߰�%�}�r<$^)�H+F�8�`]��jʽ��)�RU����sRɘ�j�����%��ӛ�߉<�`�*������-I�=5CX`K웑��!Hߖ�w�uHk1�}�p�`�C�6z�&�eq��&�	~T�]J%vF�����7���`��u����
X�쓔�V�	a9FU��+��X��~w3�͠�8UAt��W�]J;|,+�N��N۴�lmi7)2��H?<�>*pG�"I�8�u�j�[_ͽ�՝��,zT��u:!\G��L�|�U�����!�o4�	��T_�N�L�"�G�EŪsv�>�S�!�I[f9����rfߋ�o���Q�����c�����7�o����j���ذ4��(�M�n�2�3�K����Q�-q賚�����Pbf�8CuV�֎P���Z���y�~(����0Gq bF:��tt*���y���ۼ�v�`�k>���h׫6@��� ��J􁐼�7�aq�KN���-��K��wA�����z�[��e�r�c	gld�>�a��(ߪ�G*�#p�fu_�*cZ<��$ɵB�t���=)�3~3E�p�b`�Me\'�aB��������=��?S{��C�jೝ�Ō\ʑ�/΋E��+�{Q~�$�n�E#���~TK��i
�8�������Nf�$>�j�췶�{���c~L�ߗ)%���6N���p��B�8l�}��N|~A}\ct��\�:�T��%��y�)~�K�nP�_B.T�W9Z���w�E9q�����Y7j5���H�t2���&��*�j9Ǔw���vwA���� ��2M5��; D%���3����Fѭ?�N ~�!�:ѭ�QΛ�Y�;s�U� 1
��[/�����~{G���Y�֔� 
(+pp��RS3�ԓ4��洘�Tf�I���:@�X��x3�'ĸVzA���6D 1�d{�N�D~@�TreVO��~`%1�DG��{ֻ����ң���y=������
Jh�x{7��G��_�K�-����t�g�>�g�9�`�xNM)�X)�S%U��F%�~Ɔ��\e�eN�>߯�l��'��#E���8�W�u*�tN��"3�Aq`��_�ɨd�Iܴś~ǧ U��TŁ�XD0u������*v�͂�):8�"�������cu�*�:~�G���F0_Ot�����g�N��GM�Hl\�G�}ȗvO�uTc�D��>j4)Vؗ��?�\Զ.c�����b�3��+��3)y�n�����Lz�D�Ǫ���g��e� �t5��s�[,�����X؈���U���^��"���J5՞�a�?�_�j���K��$݉A���C�8��w��'C8u�j����4|e9�{:6����4R�ꍿ�D��	8פH�����>R�;�3i���V ��5qr���Y�bX�ַ��c��@գk���l�s��[��.O0�'�O^��xcdj�M�kq{��F\�;A�|=�E����3px�(��+��
�p�i�d^�J#���-E��
�!�@x��T����m�Қ�T7����Z���4Q,	�MM�T�|$��q��Y�of��Zʺ�,�
�{6b�Q,o��ʆ���O<�'��>*C"���0J�|���@���v��,yk6&��_B��S��
��Io�Ӓ��X�-%W#��b����1�w������vr���8�:N~!��Y���r�z����~�3��	~�G:��g�P�[L����/�_�hq*�]���-�ˌ� @�nC��Da�a�"���ZK9�O�&l������D�O�<�a]S���3��V�	�;{?<ŋ��{��FIS }���|KH"3��M��;$����� ���L�#:�TV��H��m���}�D9�|M��6Ӄ�kB^��G{�
���2��Y�Hpz�g����ߴ���S�-��7
 �)�v��WT�A���`�Gɫ��u��J�T���D=�m<��V(��������_쮛��R�F��?{���V��;�7�h
W+�����cQ�|�%��(�m���O޴ }�F��vɰ��#Q���]��6��>ڊH��[���R��+
X�u@$
���t�J�nR�=��a��;N`'z-��4�wg����	��=:[�H����cpi�d_��e���
A�(ƈuG�u�pUZ�5c�� ����iO�t/=X�~���pc]�����a������v�=�ˡ��"C�{+Gq��ʸyd/�����3{�'$c��E��*]��[�i1���N:�MZ�]�$�vcɌ�ʶ����9~,�Iߞل�K6t��	Bv���yI�̕�<~h�c{I[�C���\T���yJ˲�PJU8R�^�u)������ͷ� �j�m�ɏ��2�̈́-�&��.j �wi��v�a.�� �%�2t\b��G�Dn5��Y���O��8M���h<����վRY���������1��{
�ܱ���G��&Y�Q/���+A�b83�j/4<&%��d��[]��0/���@�F{�z�35���4����D'��K�N�ʔ@��Ye�b�����1V)�=*{�:z���j�� 31ޢk��9QhY*z�������@���"KMa��1��S4���5"�La9�QxU���?k��0s�v�U�&�~�n���� ��U�V�P,Ax|@�T����J�̼ )�a�SN㏎-�`�T�xw�����T�5p�[K���c�zdB������q�(��GT[wp�8	�^cD�c�өԵ�
0t�4�=�c~]O�p&�_��SNF��al�3�3ꈫ���=���i���=�+s�Ϯ��%���Z�/x��,n{{��$&R�E��%��u�ithe�gK���g�xl$�TɯF<�C��xi~o�n�A�J�h�6xش��B��M��v��x��~���c,ܐF�'�~s�؏	}ym�&�5%P� ��e��퍥x�!�o`؅��C�jA��r9�2�LЫ���jc��w,�v!��n� ޜ�2��{���D���]4z�U断�|8B)�K�I��Lxm]Y�B�C���5|1�J���*�������G:�;Y�'؞*x�+ڣJ���3v��46��qU�����3X@3�@w���A�}3�'^��w��PD� �N`�N��@Ue g�h�1��8�Jo({��>��@���T��δ���缞*h<ӆ�ⱌ�8K���JK����_jv���Q���(�9+ayx�Z�B�\�}E�FlU�(R����+e�DN����!��}M�'�I����_�5��NF3Oc�`���#:t�Τ�I���h� M��#F�p�u��d�������#�,��:"�ҙ�M��-��JQu��:�-aG	MF��cO^ ��
i~{gA���|�r��\_�}r�xOۡ�TH:������賜)@W	�'�<\>���f��͌:�a�X{[w)�A�n��N�(��z��~��'�	/�U�;� ��^H��(��bO�:D����B$U��r�zA�H�FG.D5���Ka�&_j!jK1y�s�Ţ�S{�����^ᠷo3�8I�j�>mϹl|O*��Hă�{��P���㩼n��	�O|HI|��G�RB��ĥY�ia�(V�}5�=)*íw�Lݘ���cx���)vk��l��Kh�@�/0���O��Cx͕�_�Hk[��������}|���En(�j4xc$���
��i�EҴ�ϳ1��E��
����=hS����t��2�	J7����D���G~�,smfM�x<>�$L�q�(��Qo���a,}P��%��;�)�dІ���{��>T�d�7�J�ӻ�J���L��k����I�;��;%�tޢ��	�|�X�%����KB�����[Ou��JRM�r���"�":��N��2��ٯr�v�!x�~�P]�����:� ���{�L�!��Y+��Ҽ��������k��3�Z�a�F"���^9Z&��"���C��O�D"aGP��6�X3g�5���_;e�2<�*�������Z� g�i��H��e���);����[�LA�LD?�	N�VlH�d�m>`1�g�#9�/�+OG���9�8��q�v�H���C�p����K���δ�rS��=���Ģ�`r��cA���
ʘɕ1��1���{^����ގ.vmf�Vo�E�<���gf��+�:j@O'�~]�5j�V(t;q��h�Y��li�0mQl����(���GZ���w}~��0`�a�H՚�\BQ࿡߾1
�?��?@}I�sB|7�O`M�N��NW��آ��
��o�x�žλ�kd�����W��\h�)��#�*��1�G$���d���	�#���b�4�2�
�\EI�1��vKf@V�<���G�xG��b�a�����@y�P��X���4]�����}�c"&�˱A�=g�檪�|	f��rb�~S�9a�㳪��(�'(��޿VXt@�rR9+ף���z��#1?>̐K��n�C�\ľ�����P����`��ZV@��:�#q�f�^�_�=s0I&eE��d���sr�}A�k����^sZ�t�E&zP0¼28_{PW��ՀrWc!���sbn�����Ŏ����"M��;��N����̥��Xt�8q\���%��wMTn��L_x��X�'���qf��&`?�c]�Ћ
F4�p�U��'��;,��y��0��b�n���K�4B$�ً	��ba¥!b�����糧�}�F �xӄ�]R�C��j�Eܨ�	�ݐes�	�<b׿6~9�Ik?�i15۳�`2��-�5�����~��7�$�O'�Pn�z�^���TBYG�#d����z;����=s��)�>�Bb��D�T5q��El��?:�����Ym���ቑ� ,�i뢦*;]���{A�Ob.Ttr@�6�|a�W���i�$��2";�
,��;#CD�`D�����nH�ҡN��'1(P�T:�C�Cu.a� Z���0T�+���z^�P��ul��Vv�A�m����t+�]�������A�$��?�x��ɪ��'=<�:��[�R?�h%���_'��ap�I���׫��������h���Ԗ�86u�#s^�í�ƛnѷ�m�_��|�"��n���!�%Nj^��C�%�pG����Y��H��YBy	��d0���� ��F��Y�`�l�������)�Jp�Y��Q����@��h~J@�CW�i�V�r�_���*D3�@�w���$�d�w[l����^�_I�dx�U����\��964���el��3	G���N���ƣ�`'�d{9�{~�X{󓬊��G�'�,Ƨ��4�t�&�u�z p'�E��:p��G|8�[��΢���+�?,�jA��>�äx����[8����#��+�f��"}2O*<�	�+mFno78P�P]Z�c�M�)��@�/s������OP�Vn ֗�����`l��B��F�Ф�0�C����G�L�چ��9�C1�́p~;1���.za_��h��ty~�8n] �FH姠��������q�$%q
��؇U���F�P+���X���w���!�|A83�Y)��C���|����m@$��0	t�_� �V�-2�୑W��������m�z2l�?Nm?89��/Sq"d.�0|O�I_7��n� :�i�*���P8A��:."�V���ʬRW��i�{��N�;2MȺ��GC��7�J��ϻ��;4ݰ���ĸ�F.A,7n���ؾu����_F�Bx��u���K'>�����)�J�<���7Ԓ�>�zHk�P��9�\>��.0T���Ӷg`X��e%{T��E�í=���+6�'L0r(`/ќ9�:r���^i�8��rQ-���Y~���j��
�:�ә����L�'�ӻ���\<�KЇQ"��ɡْ �T;ar"Aw��~֗9T�&7����Y��nO�"7a��F���3!w���/G;�K<iu� D��� ��'�1HF�?��oA;H��R��|�L>јC�V�d�H�l�m8_3ڡle9CՈ��y�|}�&�������iu�v��}m}pz3�5��2�����SV���[M/�U!w��t`A�:5�jR���u��G8�5�l�����h�4m�>BV)A`�6�p�&��#A���+:����ä�w@V��z;k��h.-��a�,�͹�QfP��IԬ(��?�1���%}� ��t���VՔB�ZšY��
ɱ���G+}���B�%�OZN�BWO��i
�Io��a�_c�H4Ed�����WT�\���2��$X�1����?td]�'	��	yծ����%?_�1<��v����aq�6pB�Wf�S�@f�[�X�+0���Ş��J����ɧ]mgU��+�&=����x=a�����m	�ڜr]S�]��P�Y�p���ၞ�~�俐M@�w�r��ם>��8s#�#P�J�*���}-�8:���bP�q-��αZ�����O�q���^D}=훛&�?凷�����s����kO?����s;�]t�<!&4Et�H�8��dW&.k�,�!���s���-�:�H�W�� �M�?\�?��Jz��� �Z=qք^��E��^�M���[�[n��='B೨iE8ڷil?��������}
i4j�`U��x'��,���y@:ɸ�Vf�S%�4�Mjمj�Ɯ�����q�KC��	6��"F��q�>�lR�~ۤ�4�"�ێ�!�s�� �v	ݿ����K�cF��퉡`�$�-�����'���������	�dJ��z���<�B8#^�A�;Ϊz�����oa�7<�c��r�B�@"�>�bTo������[� ��5���C�� &�_i%�**�S��sA�A�̿.���v��6t�W�WCi�ٮ��;��O���C~��D)?v�j�i��e��E'�҆PKN7�t)C�~�Ț��O(T�I��^^��;P9	�uf�4�`�AG���O-�n��Y�������&��;����øxv�٪^97R�t�Y[r>�2�%��{��E%��U�I�7W����
�O)d[���r����:uH�^�r���!����'/L�m�)"��ޫ�Q����^�R+C}�p��� &�I�Y<�ѫ�60����z㔼@'���5b��D���X��ШJ���Y�!ʰ+��&���{J�UbW_3sV�sO_��k�ZW�w��z$깔Ôˡlhd��XN�_���d��E�����V
�9p{U�YFl����
���0�FϺ�]��'�O97][~!a���q����ґ���a珫�0�خj�� *Y��P۰����ǩ�e	�$I z�/�.��� �-�E�Gز3l��
zM�9[�|��H*�d�k�V5����f�gmHCw�z����wW����+'�L�G���$�d��\(�xU,�*}X]��=&zb�J��y�y�XfFE��}.�W���������s\�]�P�{��^|ܦ=.��.��@L�L_:�T���)�Sq{�E� U��!y��tU.37���%�g(�[�-�y6^��@K�?�UQ���'�̈&�8/I|��Qb��#�G��!�$�&�)�r<���]a�/�J�4o�+���q�G�	{*�ʾ֔<�%[��8�γz������D~�����	�mNV1�{��Z]���C���Ж){.���Y����t���9����}�@ch���5�����$+�#�e�}A*�V�8PS��}���iJ��_+�`�.	2����厭���ܸ���J�ݡ�x��\�-[���6�V���a������Ւ���p(�d�q((�2�8�XDuIp,6����S�_�_B�*q�z���,�C���{�KM�L�#A���6��0�/ �X@J�-� KLJ��)�����\�>%���f�NX�:}�!t�ox�I�Z�w�D�P��%|)�uB��;W�ዴ�[.��V���� ��-�Ҫc~�z�`�V6����JʅK{z`�0a�I-�������J=�����F���~��	�ycB��I�/����#�={�r$�Eװ��B����i>�}�q}���Q��$r��ɹmU�NKɕ��h~9�O�KeT���6��ä�B�.z�F)���c~uc(2����*�$��Y�Nyw�0�ynP|6b���]ҥ�$�����O���M7�jiG���.2�N�څw�5��j�w��,v+�:�c hV�2��嗪G�DYc����&-��F���N�Չ���1��Y��^�N=���1��^���I�����GD�mY�@M����+�7k�� H3�84��������t��}��_@Az��KJ3���
�ᅽ �D����4N|��@�e
�Ҳ�91s�,^{�,����W��߭����!�K1h�c�����B۬��K:������p����HD9�q�x�w��K>���>�2q��exN3N�Cs����[��׭ߓ���E���)��N̪23Ya�`۲R����^�I������ 	+6툲���mu����nX�^���6�:lӴ�Y���=�u )�:2��G��F��cO���ДH�>gK�:S��P0\Ζ}|�+O%��T���x����Y5)�����\�����R�P��޶+��k2)AS�ni��K�z�����Fy��w��RȨl�'Mb`��D��� �r��=E�p�����N��/�Acf>�Ώ��;�Ã'q"�wͺ�s�?��6�b���$�( ����W�߀�@<�m��,$����n6f9S(F��M㙺3k����o�jcB����X����j�<F��;�H��O;P̪��o{��bFV�9�3�0ܵu�S����*�ԉ�! ��`�5��}j)'�o4�ns�n�"MN��6S�ȗ�&�Hq��`�c{�	���@��q��P6�~|��H0qag�k���1���;!�*:��E��Xp]��Q������Y���"]��g����Ҳ�]E��"�i�/���.�}�7\b�
9��zѨO�]���?�&D53Be���7�E�<�_<�|�����V$�C��D�b���8�{��\���.o���j�e�Vcvq�)ifb�b�����0��Gn��/�mx�ωZm�����n���*p��z=������ſ����:�����6�-��R&V�3�w>�R�8��pN�۬▴����G �fKR���ðRd��nɶ¬$��͜��OB��F��v80��y\�O:�AO���bQ���>�|���zl�g�X�yc��լNK�m��x��S�DTZ�����RyX7�p�`��aU��S�����i���ldm�{-U�n�-M`�`�3����>Qd��)�՛C��-�'���~l�R���_�thj��ӿ����ߖ���8k�����5���)�>M"YJ�����a��m���0�Wy������Q���W�n5w��ź�ᘊT&�:޳�k2��X�v�@�0^naLS��ƀ8`��N�ȽJ�iY�ɻ�a5@���>l��e�!�Z�0֏�Xȣ����*Zy�D�
lK"��$�y����Zs4g:�f��uoը�e &"=����4����]�|S����s�or_�têZ��)v �/�IgK�
3_|�2m!`���N�'���`/�7^x0I>�j�
������!�s#�=�$wL��tR������m铠0E7���|�#���Ȟ]u9��4�9A�ϙ>>�00��U|���b�=!!�i���~kt�Z����}1�ϑ�Z�1N!צ:!Xd�P���NМ8�;P���nA�+��ܩ"�)A�h�:?����rj���"U�t��vaO�U��>�4�f1z�S�����^�ǜ 
��t��-T�>�P#��PÓ�o��8�<+9����˕g�Gݤ�����Te����D4��4�H0!*�_��+/�����4�Ke�;�*��7Y�6�:�?�r�����CIYW��z�͚��[jLB��mn]?U��D *�d��\qf2�
�W�kLl���2��r��4��(<߅�ٸ%^�0��FwAj�4����S���-�c�۸0�׭�c ����O��ZxuU�E�*��N��
S6G	 B�V%�6%��-��MZ�,�;e(�% W��3���i�
K���{(���Z�O��ݪ<l�,����a�]�z���E��`e����8]sA�?FB
�s�Y펌F���%�����[o�ف�E'ơ\S6��fҒ[|E�\�Q4O��3-# �N?8�h{=�	�I�[E�@��X���2l�25Э�v�Ļh�_�1�R���jY)8��o�Ɖ5����<�8�.���{�����
��'f�PԆ�&s�z{���=�����&�f�a�lG���� ݪ<�����Q�֮�~n�0�vnV��#�3�.������:��Z�U �����v"��[t���[�ǧ23<�¿�q���,H�	��lL���O�2 ޛ�.�0:4�Mݳbh����.!*n0�˝�tjbp�oO��n�U�wL0o���]*��;�^��<�Ǖ�y�Ą�b,���wqQ|���n�4�Y=Q����ǝ��9�)&��G���y{����?�g�Q	�{�6��#e'��o��+��,g�e1�$���F���.8z��٣ +8�+�@3�}���<h���lF��8І�]ڽʁ�Q)!d���>s�;~%;�A2��֠d��n�M�`�?������ƣ�C�C�w��_��@��Z���a�1R�%p�}S�d�z�A��)���j��~�]�BF���� j�N%��(,)���
��%�Xگ�M��FCO+E0XF��ww�>����A��K�������Md��p�Bm�6q��k���X�����23]��hy��|ۆGm{��2��\?Ο�>�m�G�S�Ȋ(����_�-��.�DT?%�u*�G��L@�����aؾ�!����[�]T�=����Y���*�аo�'n!�^f��)�S�.r8L~�������<����v���wI��H�9���<�F��K�MD�MY���S�E�|�<$_P�-C�������b���C�^���S�m§54֦P����:0��b�z���2�t<�t1R������H���}+�6�i��@�H5���JF�N�(�KaCn�N])-���|T�w�@n�)�a�]��[s���D��cdj���~��յ�(�G|I�p@�_1�[cl���kx��Lt� D=;a�~��rpN��Un��a�`��[�-��!�=��8�%K�u���<��8��#�6/�S��u{���$N��E�������[i�g���/v�G���c$Ч���O�, �)�K~�E��iUN�yD6���	B��
�$�@̠�d~��'cF`�n����Q�ط��y����]*�P�2�\S�)�4����/ح/;�k��jG��ɚ�2/-m�/���j��9wT�8vI���� �]2��<��/�D7O �
��}�w�p`G��s�>�?���A%Yݛ�kt��x91��`�tE���i�"$|Gb	Y�(U�R��+���C3��r4G0��F���&��[�A@�O��i�>3�$>����u$D��(v�N=�@}WNe(�ҐO1�r�d{�)��������t��ǀ���ohd�u�
�Y�`g���yBK؉�������y�u�� 9S@�x ]�j)ׂ����n���P�R��Zve��N�~���X�9��u�q�
�����]�N*u{3ww�`���K�^��'I�����p� �ߣ����*,u��V�,:��$��T:Jjљ��t&���ȮYu���:�;G3�@F7�O�=��2K��(�gi�q�k���B\,�l}�|O�KTpĴ��x�h�)h���O�U\f�@5�P�0R'ʹl���)K���)#�n�W�P�z����*����}�&�7$�Ȇ�����Յ�b�Hҭ��ſU"�~�&��p'aor�l7�5񁇢s�=N�pjI�WKY_[ݛ��RC�ʻs��	a��`X8q�lj�U2��hu|w����sī���!η�����5m	��Hq����p�Rj���l~i�cDV��5�1�e�H��b�t���	ڛc�A�ν�&�y~6�u����u�a��(�A����N�0�Y�����<�o��������C�xo���|φ���[
=��*%��r�1���s��IOs���KѪ-���?"󳕩V�D����u���^*hM�X�щ���zq��f" ��_�7��^F`�Cƣp�⏭f���bQY���x�s0����	ɼ��_�+!6�~��p��݊5�JB��b����~�JR�W�|tVH�y_���<nZ��w7�A$��<�,ZMl �΍��_��d�Ǳ2Pp��*�9�����IlJ����X�F�����c�'�?�9Ϩ7~�%E=��L��*Zʧ���̫5�U�F����k� �����,
�_He��$�h}�@� .Ap ��E�<����A�z�n[w�J�{�Ȳ��ܿ�<�,�3���H�	�z]�x����gmc+��F�������`�t�� ��(
X�š��<bl���&^yOEf�JEM�.1m,�9p¡��;��s�Ż��X�{B��|t�G.'c�g�@䆓_�7z�YX�)m��{+E �G�͹a~�Ym�U�>��st4��y����?y�h��ب{�� �U�HmW'V6&���/᫸����8��GX����</e]��/>�O47:�I>G��ۤ	~�V��<I���s��K�$�+�5��#��Q�7	��bN���4�Z�������:hq����{����x�ǌk-�`��a����>hL"55���A�㽻{/�P'���<�d΂.%a�d��J<�E+�V�Ƣ���X�-���E�@�2�0hLJ�����\��X�3����ť�	�w�i�m]��|1�(�5*q�G2��0��mxI�~6m�z�E��'�_ڃq?v;�0��C�'��q�K�$kLq���c�67�oD9/���Xأ���{�K�k�j<`� �-\��a%!qf(��XN�}�!�� Ik���Y��׆%L��+/�t���yH���}��V���?;�9 �ķ-�c���-¢V� rVDQ ��������2}�{�+�Աpg���}8lf�h�Ҧs�D��]���@�*^)۳^{�D�f'>�K`"x\�4�Q�;��قa�n����8�5�||�b_u��q�Ϊ��:����:RQ\\��]S=���D[��N�R��_,m�^�Kg%��r�k@_Ѫ?,]+��hk�t��y�N3�g:4l����30T�PAk�'�]"t����Z� ���f��~�s/;�A�#���W���6H��.y��
�g4���H�[��(E(��D9�W����0mG�,��;k6�/G(]�XMCd�
ʲ�߁���c�<��JϺ���S*��2I�ƕRP��������PY�r�I3+���̀��J����W��@�!�{``��h�tj`�܆:�e�nq M^�6�D��?�����	�{�b�������l���]�6^�J(T�H���g����ޅ)�   �  C  �  �  �*  g6  B  �M  oY  .d  �o  �z  W�  ��  ��  F�  ��  >�  ��  Ҽ  �  ]�  ��  �  t�  ��  1�  ��  ��  o�  � ?	 � � � �# a* �4 �= �C `L &U �[ b Yh �l  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+a��6 \��	�<4�d5h��'�B�'���'	�'/�'�B�'��I2w��5Kk����e��U�D܃��'�b�'A��'���'}��'��'�>��5�\ h4tIR �>���'l��'��'���'2�'���'b�Iz�k�fVЂG�[�x.(���'���'/2�'��'"�'"�'�^�qs�S%V��c߁Lb>ıf�'��'@r�'���' ��'h��'J����b���@�3MTV<q�'�B�'�'���'���'^��'��`�$�͡9Ql�#[�=�"���?i��?����?!��?9���?A���?P�Σ9<�x�
�&�+K[�Jъ���O<���O��D�O����O���O��DLw�eȴ���ŢW�2(�'��O0��O���O"���O�d�O&���O,���ƏX���K�8�n͊���OP�$�O��D�O����O����Oz���OL,���0�"&�:3�f�j���O����OD���O����O����Or���Oؕ����JT�
�G�Oݨ��Ԣ�OT��OF�$�O���O����O����OH�0t�ʰ[O�XbQd|�^4�G��OP�d�O@�D�O����O���Lئ��iީ�ć/TF�U�ՁN�:�Z�34�ڂ����O��S�g~�h���%k�2�8�!#$>=�B��PX
`��	��M���y�'a�S�)� @���@-\��r���'�R��5Ǜ����'r|�Ę~��!O1*�E� � �͛z��?�.O>�}�1�A%��D�(�����6뛦����'5���nz�)����Kp�D��ě�D&�!�����	�<Y�O1�N��ƌs���	�3��2�,yp����	�>���	�<��'�@�G{�O�2eʝ9f-�F�@1�=�3"�.�y�Q��$� Y�4+�(�<ɠ�L���(�&K�	H�JU�,��'�(��?)��ybQ����J۔Zx^�`��F�t���01
"?���j�l8�aB�ḑj�n�d���?)V�Ѣ�lG�M:9��0���#��D�<9�S��yR
�M�Q0EJ�h�*A��-�yR�|�8�[��`�4����4.��";���1��3B�ڰ�@:�y��'�b�'n!�T�i����|*��O�l�b�}-bCVBŕJ�(pن%�f�Uy�OF2�'b��'��lS?^��U��F��X�f�ھY��	*�M��J����O��?aQ!!�(AV��"�#E�>9�wI���d\Ц1�ܴ!������OQ��#�S��` `�&{�J����Ӹat-�A��GDҫ�N8��������@≾��?;hdTY�PM~n�¿葊D�'R��'����P�\ڴd��Az����P&�Z��ya���"#d����1d���CY}��iӌIl�M��4	x�AҫA�K�^��TL��F"��۴�y"�Q�R����@ek:ظ��'��t��0
B篂�E�X�S�ꑈ!����k���y��'���'�b�'����f;��5I�:}�HL:TI%^q�$�O����ꦉSrn>��	�M�K>��]69yzѦkڞ.Qy"3���+3�'P��Bb�2��[�j�7-������12�n�y��@r��1}�*��C�rʚ@y�%p�0��|����?	�x"n������{����Ęj2>:���?-O)lڍ|D��I�D��u�4�$9d�͹H��j���bU������T}R�t�Ȧ��N<�O��å�ކV}�#W�
�T���S�)�/\M��3vF�2���º���O��!.O�N O��A���c�a	�*��w�f���O����Ob��i�<���i��AC̈6䈍� �:PH:t�a�[�4�R�'p@6�)�I���Ē���� �'��	Q�Ƞrl��wKÿ�M�ճigܘ���i����O<��D�
��c��8���3^ra���Xz ��g-�Mc.O����O$���O�$�Onʧ9�����f׃!�*��D�j��P��i�f�sT�d�	^�ϟ�R���+r`�&��y!wf�"u�iQP�ƶ�?!�sd���O�\�0b�iY������� �t�2�C�$���M/	,�	�>ʓ�E�ey�O���8�t�bA�.�p�ĉ��Q��'s�'���!�M�bM�?!��?	�
� |lMJ��L��b���(��'����?I����'V5{Ei�-a0��q�²)7����'�����١B=��$Iƺ+���O�A2���.��r)�ezDd����y������?����?)����F�n�������1� �x��\R|�'"vj���ͦ�8�� �	��M��w2I����- E*�懌x��@�'���p���l�
�lZ�<�7<��;p�0|!D��G���z4�>;X��Ǚ��D�Ԧѕ����'��'��'���F��yt�)m�L 	]�0�޴c��m����?����O�Bp��-,"!�s�]!gj>���	�>��iw�7g�i>����?�ط��,Ws�� `�,5y���喽Z%~�r��/?	�'�-p�@�d��ަ��'��t��U������9Q�E���'���'}�����X��0��Z�8��\^|}���2R�FȂ7Bњ@g�L����Mc�2��<���M���i>~0��͕!l2%��
>�h��q�ܪyk�<O��D�>T�H��.C�I��u���� �l!$K�Y�Q�t�Sh��2O��d�O\�d�O����O��?��`l�$���#֊ 
@#G.�ٟ@����؉�4f(���'�?��ir�'��M��L�����Sd	
er�y�|b�j�R�n��������!̓��a��٭ho&����+���A!$бg뾌�F2A�֑xƻ<����?����?���Кl�B��!GKG��)A�G��?����$
Цq+�L矀����0�O�02Ŗ0l����N���O"��'���'Tɧ��y��ჯG�8��-pGCI�w*z����:�>����[p��y�ɃHQ�0���\(�`��!Ɛ ����ş\���`�)�Suyb%u��V�[rR�u��FږM|pt�BN��E���d�OFim�O�o[��֟�т'�='�r� ��	�����mџ��ɰ+�f�l�<a�xN��07��Hi�'��a���*��2BYf�D'*�I����I����	̟���b��MÏ�Ƙ:��ݗ���,/�D6�C���d�O���;�)�Od�lz�5#ǟ�Hl�3��J�Xp���A3�?�����?I�S�?-�EE��)ΓQ��g��8�����
/�H�͓}fލ�p��O0��H>�(O,���O�q��`h���E~��3��O�,#�i�O
�d�<�ǰ��Z�$�O���O���A���r���cJ�S8tq���(�ɱ�����}��ē*?"���
�Do p³b�Lah͓�?1��&;`Q�� ���D������ب��A�H���+u�G.h�Ѥ䈦�4�d�OR���O���'�'�?qe�Ə8����O���/߈�?qQ�i
 ��#�':2�f�P�杣]����V.<Vpz]E�ž<|Z�	��M���'��6o�>��6��Lŀ�8>s��,� ���֏֑ H\Q�'��k��$�D�'(��'vr�'6��'�2ԋ�g��	2�(Ade��Bk�pP!^����4SH�z���?�����Odn�j�/۩l�|��R�ò"�[���>����?	I>ͧ�?y�%z�kQEC#g�~��1l�\f�eЖĎ�M{`X��2�(4$t��9���<���M,JA8�!�6W�u�c&��?i���?Y���?ͧ��D榅SE�@͟,��JS`��oW#�
�!w�S�8�4��'HL듼?���?	T�R����`J9�!�Q��$b��A`ܴ�y��'
	��PIR.O�i���|8�ㆊ(c��b�ǿ~���@A7Ol�$�O����Oh�$�O�?���"!-���AB�'����˟�	`�۴'����Oy�7:���~S�e� ׶k�Z!��B�NF�O���O���"7Mm�P�	=T���)��E�*=ބ�����:'-B�r�X�]y�Ol��'AZ���Zs����X�C�̑a��y�����'�7�J�n� ���O4���>�)��o�ƉscÅ�`<��E.�ɔ���O���<�4���d)J� �I�(m�����)G	(�"6t���F��X��(1��W�	S��Ţ�gH�W�Fx�FP=qw�Q������I����)��pyR�s��%b�ɬjں9��F�<eZI0��k�����O��o�k����ɛ�M�2��)q�c�.ޛ- �����9��f`nӆ�Q�n���I͟\��(\�v��� eyr���$���(*��m�ZaJ�Γ��D�O^��O����O��$�|�'��D�HU�0��*4)����-G��_
B�'���T�'x�7=�QS`C�y���6�K�o�ʨ;�!L���������|��������M�'�\�����8-A
�"Ĝ~�Ș'Ɍ����pq�|�U���I�X���ה{"�H��oE�%�R�ğ,�	ş���yy"�y�0�j���O��d�Od�C�R�I�A��� �UC�n'��+���ƦM����3�0��3"k ����W�a,�'@� 8���{�d0����X0p�'��0���Z ��s�����'f��'���'��>���!U��Q2�c�R��8����Q��(�	3�?ѣdΟ|�ɾ�Mk��w�p�$OЇeF8�e�J'mn�,[�'2"�'t򼔸��4�y��'0�4ӦǊ�?�Ħ�8��%SU�'Mh�=+�/m�'k�i>���ޟL���P���c\œ��J|�&�y���1K��̖'D�7M,^����O��#�9O�M)\@Yk �\��Zq
��I�'�x6mY즡�H<ͧ���'&��ɠ�˝�r@��b��&(��+֎�M�ȁ�'HP�����蟸E�|�]�p�TJR7l�Y��K�rnx��K��0�	ϟh�	���Iy2,b�X�[1�O�8�3�� �@8zŃI3 '�-zB��O��m�ʟ4%���O�<oZ��?a�4|4MStO� %0f�ځM�0�@a*(�M��'�b���b,�S�l��?����3����4��}1(Z�K��I����	ݟt�Iݟ��I{��,�,�Z����Y�C�������?y��	�V������'y>7M"��=X�ڰ���
"������Qzx�'��n��M��'�Rq��4�yr�'8�A�p�A�&E����M07��Q�!OڶK����<n(�'��Iʟ\�I����	>)"�a�d 5g��4s�JE)o*��	ן�'T�6��^����O����|��j2>��#��"9�q��k~�+�<����?�L>���?�+@ج�L�Fk�h{Qm����@8n��'����̟��R�|U-�@�T�@=0��(@�îw���'2�'o���Q���ܴ&s0鲴�S�^��m &�L=\.�xk֢߮����ئ��?Y&V��`�4~\2���u��ip���1*[��Bҵi��7mA	M�6�h�p�	�y���G�O���S�?  1؅#�l�\)�`��n
<S:Ot��?��?���?i�����ȳ B�q�EИhJ��jE�QE><�oڤ��'�2��4�'�86=��۰�J0t\�|���9N
*ac���Y�4=]����Oj��H�8��F;O6�[�����5�?�@��2OJH��+� �?��(�d�<ͧ�?�B)�2s)rt���N/|MHh��>�?����?!���dPĦ���������ӟ`B�ۆIdp����A�|^@A����B��V�������IL�;P����8f�d�gML7N��h�c�	�Pr�ԣ$?���.����F��?��j��FL�)�u Ι�ĩ�@@��?���?���?Y����O�@Ҵ�ԙ2[:D)6LN�z�
�G�O�}mZ�NH����ϟ���4���y���BK�1���U�G6��H��y��'��1O@a�¹i�iݩ`��Kj�޸B*��`�K�D��{a�������O|�d�O^��O��$V";c��cJ��U"إ4�Z>/�˓U����q���'�2����'���˵�ұ_k�5rE]�e��xҀL�>Y���?	L>ͧ�?��8� q��,!1|͑2OT�q�EBE���M��P��#�.�*��d(���<!T��4j� ɳ�҇n�b�
���?a���?	���?ͧ���즭��k��0��)Ţl�:�����A�V�1�����޴��'����?���?q�l\Y�X�y�M֧`��r1/�/Yz�Q�4�y��'1���LYx:,Od�����0�Rd�%� ���s���8#4OD���Oh���OP�D�Ol�?M� �Р|&���lϭ[DV����ԟ�Iܟ�{�4WG2tΧ�?9��i��'@J�xmΝ.J�\�IS4`�B��$��){ܴ�u���M��'�R�D�w�B���O�~Gh�x!����^)ZJT�\�g�|2Z��S�4�	�DP�����h�(�I5�ҟ��	[y�#r����`��O��d�O�ʧIv�i�	�#�șX�IN�dq�Y�'c��$p�6�nӊ|&��
*�٤ꄹW�"��� F�)�����2�ր��i�H~�O~���I$v�'i��PŃ0FtpPs�fȏ|�n3��'c2�'J"���O|�	��M�S$�UK0��W ��ut�U���F-"���A��?�T�i��O���'��K�{$����$�����W/r�'Dh�!�i}��OD�r��J���W�W�WL�k�nȠ\e���n�\�'���'s�'�B�'-哥:نUp���0^R�`D��Ed<kڴB������?��䧟?����y���H�dh�!
��Vd���A���'�ɧ���'���	N#�F:O5�F�F������)d�:w:Oh�`��x��I���'u�i>q�I���E�Ɏ
(TB�"ƿe�����<����$�'�6��  �D�O���F�a�Q3	O�&�u�Ga�� �~�XٯO���OԓOb���M�I��/������=�y2�'~�}�������O��)���?���OD�Iф��0��F�	�x�H@p���O����O�d�Oң}2�]� ��ܟ}�*�s�,�1Zt���d���u���'��6-9�i޵R�*F�Z���)d4AK3�m�Ъڴ,*��j�,dpaz�j�IğH��OS25d���	m֘�hC�]���,�'R4?(�$� �����'�R�'���'bb(��7y��q��G	��8�R��K�4R�P��?Q���䧗?)�:9�t�S�U9�@�`�W< �	��M[��i(O�����ɕ,l�A�$�ܐ.��������b������Hp�Im^65)w�'���'�8�'+> P�J�0Ju����O�9Be~i��'�R�'�R���X� �ڴZ�H0@�:�q�6h�.U>U��X�V�z,���V�����`y��'���GcӤ���k� O�4�pm_�	�TQ�4��6�f����#*�,���O�h�����3�b�+hH�8V@ES�B� /�b���?����?���?y���O�D�h�I�
-�������nT��B��'�b�'|6;��I�O�mE�	�rJ4M�E,M�l(�LA�݊y$��:O<���i����O��y��i��	�r�4IQ�-�;�bUb�B����v�͓7����{��Ry��'c��'Z�P5"�JxH��G�]6dţ��3|V"�'m���M��
H�?A���?�+���R��E�8�-�b��/w��"����R�Ox�nZ��?�O<�O�F��bE�BXΌ; '�((����mZ`&�����B:�i>��0�'�
�%�D꓌��)�ܩ�v�%*�\}"QO�㟰�Iݟ<�I��b>9�'Ȋ6ML
"~nL"%�'H���
�%tO|��g�O.�D�%�?9�Z�x�4�5��c� ܁�
(UX^I3żi��7ʇ]cf7Md�0��5v |#��O�@��'��ܳ����R��ң/5X耟'I�	ϟ$���t�	���I���A�J�Όa��k13,K�l�n6M^.����O��=���O|amz����<1��)��D�g/���J�ɟL��^�i>e��ٟ�Ce���͓�άX-I	�pX�r�ʈ5:�Γt�2����O��PK>1(O�i�O�%XXM&(m���~�>�.#���'���'��I��MS���?����?Ɇ%̯O�6(�W.��x�W���'Ҁ��?�����'��l� ��$ �����WH�H͓�?Y��S�U�8��4h�	�?�J��O���ٖ@#��֭_� �@��Y���$�O���O��D<��[�k��=&��e�A\S:���%_<�?Y�iKZ ���'�b%w�D��c��=:��ۀN;��7�Y�^q���ßH�	��p(��¦%͓��Ԡ�^s�� ��2���NY�b�G3/��a9��"��<����?����?���?Ѳ��`k2���U� � ��텶����զ�ZЁݟ��I���*� 9	��]�U��*̀H	��,l��	�����`�i>��	柌c�/Rt��BFL�g�.�ɒ�Z�r�J�o���N�[�B�k�'��'��	ۮ8B �%Ml4Q3נ�&��I���	ݟ��i>і'-�6�\m������5��\�Q�m��p�,R��lJ�',6m-�ə���ߦ	�4՛V�#x����Y%8_ؘ�gӬJ�P)�i>�I�M(*1*1�O�q�,��D3~!h�;-4�!@�՝w����O"�d�O*�$�O�$0��1��v	U7��ysb2Sꌕ'~"�j�X��A7����ۦ�$��#�ر"^��Ɣ�:�`�C��O8��w��He�J�i\v�|7�d� �	;J�ac��� �i��'Ԍp(�7�O�Wor+�V�Ipy�O��'�bA	��,Uӡ-G�,$�cN�0< B�'���/�MC���?y��?/�Ќ;�/�5)2���Ε�C��3�����OB�o"�?�N<�'�ZFGI"�b@��7t��G�N�lt�%b�퐯}���3)O��)�7�?9F�-��5;a�uyaa[�X{��PDĻV����O��D�Oh��	�<I�i#@� ���6|��l ��'hE*52NA�R���'��6m(�	,��d�¦e㠄�K��ð�$ N�E���MC��i�ʜ���iC�$�O�,�_�
,�<94��5!��Ђ/-I���"��`���d�O���O����ON�d�|j����78J����J)^�-r��/:��vd,U���'eR����'�6=�8ʱ�6����ҡn���a��s����|j���
�/	�M��'sH=3���C��q`a�
=*-�y��'\��3�J�ğ�B�|�Z����՟�۲�46)b "�y����I���I��`�	Zy�j���q��O����OL��\���y�o�52Ҹ�2�4�	�����O��<�dKN
he�QŖl⨅c@�ٿb���O�%�K�N17��Dy��OW�|��?y�h� ��8*� ��4UGi	�?���?	��?���)�O��Ұ��+:���i�����ְ�?Iq�i�tF�'��v�^��]:V$��-D:�E�l��I⟸�I�$җ��馥Γ��4C �l���I�y��M���T�:�d<{��7 �Onʓ�?Y��?y���?��%-ؔ�� �m������<��X@(O�nڙ�~��I`�	v��TQ����p���b5G���U���	˟�'��S��h���*j�a��³s�ܨ�WLX) �B8���ɦU:,OLyb��~�|T�l�a��?����rS�VZX����˟d���$�	���Cy�r�X�+�/�O�Y0�/.������ �Bzf5 �M�O��n�P��I��IٟL�����S�� d�B��D?��P�5X'��Im��<���g�������'����wS�\����S,�$[�凭:s�h�'��'b�' ��'�p-8R=i�l=�	c�K.)����O.�����0�Ap>�����M�L>ID%L��%�-ܹw���� ���䓧?����?�˴�M+�'���J
����T� �� Ĺ_���u�
͟� �|R^��͟��	����m��fa�]�aِ#F(���ߟ�I`y��hӈ �$/�O
���OHʧ3�~XBAظ94��	�"R*�M�'��?9���S�FQ<jD����+�(��Ř6b�B��27����O��A(�?y:����=���X�/]�D���ȕ+T����O����O���I�<��ip���!�Hz�D(�2�@�Ȇ��80��'��7�;�	����O���BH�>u��su���q*�I�v��O,�$	6X�65?��O��'�V�)=�b��QJԇ&1S������y�Z�H������I埤�	ڟ`�O�XI��D�v� wK*�	�0�r��q�C��Ob��O"��`�$�����$ih5sd�L�sﰁ��J�_LL�Iӟ�'���������Xl�<y���WD�1�@C
?3���3���<iE䋞	>�$_,����4�4�dR�:���7DE)�� ޜdu��d�O���OJ�1ޛc�{;r�'��m��c�PX8`ύ�uJ���)0���|b�>Q��iV�6M}�I�2I�{��/6������&]z�I�l�Ҋ\
6z�hr�7?���o����/�?A�>m�f��8,�����+�?y���?i��?��I�OĜ�E�C�X����[�Z�ZU�W'�O��m<�}�	�|0۴���ywM�*tJ�����1O��E8e����y�h{Ӑpl��MK�ׇ�MS�OR�St�Ӎ��N\H"��Z1��� �j|	4��T)ƓOl��|����?y���?���hK�6s,&D&$�d�"My�g�2XX�@�Ob���O�	�|���mhR�*��?�2u����e3�V������8K>�S�?����>���
ZTi���9�E�go�H�L�Csa[4/�OޙZH>A,O��i�"M�xj���#ȸArSF�O����O*�D�O�i�<aƼi֞- �'uLAG+�7!$t�v��&ZT�YG�'��7$�ɯ�����C�4>�f�N"M6$�G�F�d�.JcbV�YT��	�ia�d�O�̒5�ݚ�;^����?U���W�(�����wz�� ����X��۟T�I͟������	V�'>Y���bJG�:���ħ�5Q�d���?���eD�6������'Bv68�����u5b�y�NU�
H�� �[��M#���.ôh�֖� p#n.� �5P$��H>��wkG�&���XR,���?���*�D�<�'�?Y���?��	�SS�X �J�3i���Ñ���?���?���M��E$E��?�-���lz>=�e�;n�a�s�S�U6����K2?)�W�(�ܴW�f�;�4�D�I�8j�2V2Ch�œ�L=*��`�Cɸy��%c�����p�bH�y�	�ntܠ��	�����'�8dFQ��ߟ���Ο��)��\y��x�@��(ӓ=d@Ę��:/,�?(l5����?ɴ�i;�Oȩ�'p�6���;�@����Ts>��7��>U�z$n��M��b��M�'lB���ɖ��ӿa��Iy�`
�ڗK�Mp�R�Z,��	gy"�'���'�r�'�RX>�A6I�8�����5M=���
�Må���?���?�K~��9���w&�H���B}P�cs�E(Km�D(`m��\�IR�i>!��?y7%U̦�ngDLKg'x��xѢ*��ǮΓv֠pjGI�O�AK>I/O����O襹b�A&(���R�ֶ6gd�+�g�O8���OH���<)�i����'���'r�%��e݊v�l1�Z4���c��V}�}Ӭ���u�?��#g��/!l�Ǆ%��������V�}&�,����my�OU���	�v����ҝ�2	�Z�z@n��h*��'�R�'�R�s�%��B�#��y���B֒��2MП��47��%8���?���i�O�N��$���eK�O,�sT�ӥ3���O6�D�O8ܹf�{��	NWi����� �)4�-
�J��<+�dܨ?A�'��	П��Iԟd�	ԟ��	�|ǐ9�eT���Q��N�A����'  6M�)9v�D�O��$.�i�O���bA	N�J#`�;v�˒d|}R�'��|�O��'C�YS��^)6�g�#v�j��R@��RC���<�U˖���{�By�F�	)VK�bp���e/�N�B�'���'��OE�	��M�r�A��?�@��=a�,a�ܩ#�*Aqv��<i �i*�O���'�R�i�6W�����<��0`%�C����m���韬�AR(�$�-?q��ݿK��Ո��̨C��v���n�<����?���?���?	��TCŝEOF�" h#ބ3�f��E6��'�2�j��P���<�'�iD�'0@be�P�L���0�+H��s�A#�dL�!��|J�e���M��O����GH�,3Q�@�w�Z�x�6��I��?aE)�$�<ͧ�?q��?᠊��ID�ժW�E?t��q %
��?�����ڦ��nF�������(�O������N(KVX���ӕ�1?��R��)�4v�v�.�4�P���,'6�T��v�M�vI�.��̪fc��*�T��A����S�R"�q�I(�
ZQ A?��=��O��������	����)�|ymӾT���?e��Y1c�u��u��kݒnK�ʓb����A}�Di�|D��E�>0`��G<��F�Ħ��ߴ(���ڴ�y��'�����?���O��K'MX�4�hS�`F?¨��8O���?����?���?1�����Y9S����bG0c��T�@�ӧ,uoڳ&�X���ԟ\���?��OQ2�s��	�O�6��3�Jz�0G�ٲM3P�d�O��O���O��D�3gdT7-v�ti��֖\�32	�s����j�`9!�N�#��$>���<���?��(�JZ4p�Zpm��U��<�?����?�����ܦ�a�L����Iʟ@����0�L	Q�̄�%�yJs��E��qh��ȟ�I~��\C(]��o��B��U�ϧx�R�����-Ė��oڊ��埠 H�'jbV��l�0ß�t��9i�׶�R�' r�'2������A͞F�Di�a�M*X|<(&��۟���4a&�i��?��i"�O�N�m>��f�DJO�d c�U/z/�D���Y��47�v*l��;O�$�t&n���'j>XI{�ˍ;PDr�NL`�܍�e�<�Ĭ<!���?���?���?�po�u�f5C,�3gFb�JA�B:��$V��9`C�W˟�	���'?�	WҔ�Z0-m@^�`���\���y�OmoZ��?�M<�'�:�'"�xtag�]qQ�Ұ5즐-^����@�Ty��62*����W�'.�I�:��x�ǎ�	������u�~��͟��	����i>��'�@7���j�d�$�������o��Q0��}���d�y�?��Z�ܳشw2·iq8y�nٱ$fP1�)	j�p@�eE�����$Á�L��,IS����	 �A<fT}���"^���x1�w��������؟��I�L��G�\!x�JV�{�j �?����?�s�i���	�O�/u���O�asP�R�i�$�A�
�6�A�8�D�O��d�O���jo�&��~S�I�.y�mӠk�c����`�!ڈ��'B�'@�i�MC��?��H�z	��@��;�8D�dk?mImB��?i*O�m�{(�x�'��]>�"`D!?�8߱ri 	��6?�Z����П�$��)��2�����\E"Ř��MN`t�7E��?�h�5e_}���B%��O&��H>�1+�37B����Z]�Vt�R�؅�?a��?A��?�|�,O�,n�#Ğ�HD�Z�)�v�F�	� �R���˟`����M��2H�>���(\��!HƄJ��Q��l�+���?�����MӜ'���K��SQy�!�j 4�&˘4O��;���*�y2R�8�����Iڟ�	����O��Y���r^ڹ��͋�
K�U���}Ӏ�QP��O���Od���|���w%�4�5�>KFȰ���
��XU�h�f�l����|����®�MK��� �uA�&F��%sbAFD��:O�i�����?A�@$�d�<�'�?���KpH�ps+W!z���&fC-�?I���?Y����ܦ�K���I՟����f�*����B82�E+"�~�VD�	�M�R�i��O.�p`�5:>� 1`Fi�X�#�;O2���Nf��$(?G>�	�?���'�|X��'k����`ޭ���pK8BP�I�����ɟ��I`�O���W�J�,-�gO#�<�c/�
���uӆ0�`��<��i�"�|�w;��` 8�0�Q.C�+z,��'�6-զ���4�&M��4�y��'�6(�2��?�`�*����S���F�r����B�|�X���x�I���I���$��S����af�>ĎD봮W[y�a�@�zdd�O��D�O��?��w�N�_���Pn��v�@�)������Ol��,�4�����O ��A��'-1�J��w�ى��T�jPm�P��8� �-(�`��ly�(R2^�:s�b��TLs�*� ���'2�'��O�剂�M�E�Y�?ѷ&�5�P��ꄾ6	Bqrb�	�?a��ir�Ob`�'�"�'�r���bȠ���
y��ȫ���`�qJ!�iV�D�O����S����ߡ��N��@j����?2��I�u������ ��̟x��������(]uf�a�	�-	�:,+����?����?a2�iX���O�GsӖ�$�<!qg��9!P�ެ���������?����?����M��'������=�4��+�Ѕ�zv&mꡏ��x$���'2�'���'���[dH�g�ݨ1!��^��$�'�rU�`�4s��(���?����i7��x��X�zf�S֠�9)��.����O���,�4��dX�V�N$6�Cjh��%F�|�V�ݭ2��7_yB�O�l�����w�j�����n���4ȹ�()����?)��?��S�'��Ė�q�%�"b6 �td��~����7u�B$�'�T6m.�ɦ��������‮MH���Z,UD)1�m���M���i��u�'�i �ɭL��u�t�O_�' x�|J�Ӡ1���Q�nW�,
�1ϓ��d�O����O����O��Ģ|ꕏ^7]��j�9'xщ��-r��f��� ��֟�&?��	�Mϻ~uVQ�`���p����O��q����v�i8���0��iLq1.7M� R�!��eSa"�bk�����y� B@��)B��X�	py2�'��.Ԯ]9Z���KH�4}PB���e���'��'^剑�M��]��?���?G�Y�CZ�d���? Bf�pEh���'�
˓�?���ēe�,l�I�q_��T-�3Ǫ8��?�%�=�ذ�pL������VH��*��X�l��lƶ䚼��] ����O(�d�O���1ڧ�?�r�I}~��� �ȌD5�A<�?)e�i�L��':��j�F����h2�j׀
�"UqgF� >��>�M{r�iL�7�T�F��6�x���Iv�l��O��,5&�5|p��fO������a�P��sy2�'��'�"�'Q�̓�~B�� ��N<8a�y",T�&��	��M�G���?y��?�M~r�)(��a�W�C�`iQN׌L���؂R��	�t&�� �	�X/�x���j3��ڀ�K*P�m��B�7C��U�Zj&��O�[J>y.O��HA��Ͳ�Ő�j����qf�O����O*���O��<af�'���Q�S��1�$�� i)GkL].u9��w3�F�D�L}R�'T2�'yX�`�
q��+��{w�T��GM�p�6Or���B[� �����	�?��])�4}cӪ�`�I�ǿ|�n�����Il������	U�''��q�U�=�XX��W�h.pR��?���( ���������'p7M*���!4N8���W*`M,�J�U�{3��O,���O����&9�7�y���'��)�z��DD[,Xnx�&���~�|�\�D�����������*��y������/(���1��_ɟ��IoyR�k��8Q�<�����ͨ<���ɗ�U�\5��D�9g��ɰ��D�O���,�4�r�d�T�9�DgX�|�~D�EcͰ/�RP��-	�rU�w�����J ��O�&~pH�B�)^	r��e#�(��1��������l�)�Sy2�xӎi�@�Q/z�d;5���7��{�h��H���O��n�^������� 9��ÐVlP)*�g�l�����ܟ��I���al�<�OP"�ן`�B��jP�[$)~�����l]���d�OD���On���O���|ruc�28����-?��E+�B�{��^|'�	���&?��	&�Mϻ^3J,�pk�"��)Pr��:
H|�����?9J>�'�?9��B<��C�4�y".�":��F����Fj}�	�N԰����OړO���?���ohP�0O�JiCi¬��
���I�����^y��jӢT���<���h�$Ӂ�z{bI����)S �5�����m�ޟ��Ik��HtDj_�ųիR�W�v���'�6B�J�{�,�FyB�O���	�R�k.!:l�	�d7p/��%A�B�'�'W2����ks� �2��E�hm*�2�n�ޟ���4�v�����?i �i!�O���o{�C�m�A��ɈC/ֽ0�� �	�ݴx0��Ϟ8D��?O��$�|�P�s�'h{.a���%)����W�f�h�{��;�D�<����?���?����?)Ak�)y^������0^>�{�g�#��DԦ�����꟤�I���&?�����\t�'��wM��,&��h@�h
D}"�}��(�	F�)��@zl� n��g�P�d"e#��{T�kGI>V��˓b�D��N�OF�SL>�-O`eceK��w���VBѫc���8���OD���O|���O�)�<9w�O�ԩ��ߎ��G�	.M$>1H���)�����D�����e}��'3�'K��"�B[�y��0���Q�s���C�m������n(���4����&��k۶O��J�,�$K*4��&=O����Od���O`���O��?��Q�I)+��lʱcT(�i}y��'�z6�O�
����Oz�o�g�I
~<����h�{v��AE ���$���Iğ擕9�Em�q~ZwR�țO
-C�mI��'TQ�-G`>Y��D"���<���?A���?a�*�Ft��Y/���3N�r��	��'�H7�Bx�$�O��|25Hίa�����U)T�$�PD�L~� �>Q��?N>�Op2a�sd��%L<A:�ğ=��3'�>S��"�i����|�2���x&���E`�i�����2a���;��
ޟ�	��`���b>E�'= 7-�"(e�DX��H|Hd$�`�B��P�Af�O����a�?ɑ\�t�޴��i�eՓ$>)1F�-�<<�i<�6��'*�7-;?�!�(=�	3���T�7ʊ�9�Ĉ�e��lP�aV��y�\��������	���I�X�Oy,X���@ pT�E'O({z}!�eӶm���O���O����� ��]�Re�vm��s�,�z��Ģu�VTPٴlқf�<��צDn6-u�l�B̄D��5!D(y/li�F!x�l@D�ݕC�R��v�	Uy�O�2(17є�[$kUy���ׁ@�P���'�r�'U�%�M[R��?����?	R"D�=!�P� �e���C���!��'p�] �-|ӄ&�ܲ�$��~�ĩC�u�L�c�~�0�I�H:� Dm�9�����qh�O,ѱ��^UB�D�)I��U��0��P���?����?1���h�|�75T�)@'-,Jf�9W*8�D�ӦAr��\�I��M���wd���t��mO �p�jU�%C�r�'b�'��䎄x�V1O���ժBK�4��'T���	;y�Ҩ�0G�IJ���Щ:�D�<ͧ�?A���?���?��c�ŀ�Q��\��Q������d�̦A�����\��Ɵ$'?Y�Ʉs��0�D��+�w��7*�1�O(���OP�O��O���',rPjת����W�%�q�m�"'�I� $ /�?qpB7���<QA��6*��WN�1[$�
��q���شHk�s�J5\u�#��(,5������α���C���ĎP}�'�b�'���Aq���b�Ppc��@�&mY�m��v����Tc��pq�	:�	��6%1E��;G���Kx��A�:O���D��-Ɉ�x2���h �(��Ć�.�����O�����+M3
4�i�'�뀘�"C�a����b �!j�	ß��i>)q�����u�?}#�a`'m��^T���Pa��_�����O^�O����'�蔐�߻J>���PӪU����A����j����	ӟL�O?�ä�
����.T�a�l�s�O���'���'iɧ�)���P��Aɒ��)YQE�<o��n�3�86�Aey�O������}JD��)͍������{J^���Q6�v�� ��y4�kd�X�'�P�x� ��'�oӈ㟴��O��d�0�����}��P@  7Stv�d�O���a��Ӻ��O����T�|�1E�o��D���U��ڽ��`�X�'��{��Š&i20L@�JW͸å�z,6m�����O���)�S�M�;�~��!\�l�� ��8��A����?�I>�|�����M��'� �	��ȍDW|�B��\���`�'<�dI��Ag?!L>�*O
�K���RF�*6i�36�,�ra�ቀ�M�$*�<�?	���?�qƙ�0��X�%#��
�Q�Un7��'��듐?����!�\LPAb�z�>p����%Q���'�P��V�D9E/��K!�釉�~2�'߈�hE#*2�� �3��ͣ�'@�x����g	��c0��A��+��'�7-��;���OzDmZD�Ӽcg�X�ed���g�9[P�֤ �<)���?��b�t۴���������?�Ѐ��&KDĬ��-s�]KQK_�IRy���!3�~|
`��LԮd��$�/	 r�'�b�iÈ{#�l01	A,sH�K���j̈�'�B�'ɧ�O8����]�V!�Iک~<�)B��(u�����<9�AC'�@�	s��RyүC�ya�ܰ��&��@)�#���0>��i�Ͱ��'�L b�ڤ&��MXb�A�{����'2�7m2������O���OhI2B�ːv��Mp%D�:PB��$Cٜ7m ?�K��]���k�S��E����b����Uf��G$��jd�e����� ��<p'�]�p���h�HZ:P���ß��	��MC��VJ�D|�ԒOzP����7,!��[
&��"�'��O,�4�\�s"i���Ӻ۴cڗ��A�a�.`�@��`��:��y��'��'��	|�l^�L�<�(	��D�>'��Ex��cӴ���O���Oʧ`��	��P+^X��+Z�=���'�$꓍?	����S��  8�цWŤ����_�P`��n�gn��ɤ	x������$e�f?!O>��O<GD�8��:鸸��nDz<q��i$���X�Z	Z!��.�)h�xCmĒjE��'�@6�-�I�����OҸ� 	����%E�B�O��jq#�O��3p7�9?��5��!�O�"O��`J.2P10�	q�<I��?	���?A���?Q.�re:����<����JzR�zQ\��r��,��ȟ�&?)�	�M�;6�t���m9�Z��S�y�r�bF�i��D=�󩃦B��6d��:��ֳ!�6�ƌX��ؤm�,RbÍCoR��X��Ly"�'��cҖ'����b�0��s`M�$B�'��')�I��M����?i��?���T�[Į�b�cLb�U���Z���'���{ƛ���O�O,)+@�J&m0��n�����\��&��P��Ih�C�w�R�rC�埄��aJ=S|@(+FiȤn˸Ղ���`����Vr����1�'�?�m�"?�~�A���Z���tK�$�?qa�i<���'��o{�N��]23��A�0F��\���dT�#n��	̟��ݟTh�I�צ-�u��-#l����D�!���l�t0۶�^d��O~ʓ�?I���?���?q�'%��چG�-g��z��H�{y���.O|m�*9�������H��W�S����'F��ԃ:6�	�ɋ
7j�%دO��D�OR�O1����Q�^��Ba��"���TQ����6mFzy��
u.������G�QS�P�����K���q@��p�a|�
i�(-b�+�O�M�!�]���|8�L�xd����O0�oZX��r���ܟ�����XD��>����e�EK*��P�Pm�}n�U~��ʑCY����䧩��'�G��@H�I��9&�Q�<q�@#$0�����7pȘ{��W<7Fr8"���?1�xg�����IBܦ�'��z��(e��x��j�40�Ĺ[�h��8�i>
'C���u����Z�V�@�Iߖ�+" Nq����Op�Oʓ��'Br*e�+;�ċ�D�{X�PC��$�Цɒ����8�	Οx�O�%!��TqjK�rჇFH~�Ŵ>���?	J>�O�0qU�M��H��^�f����
Wq|+аi���|��+��x$��S��aڊ�J�(�C�d�3j/���ڴVf���q��,*�ٍM�L��G0�?�������Il}��'����N�%Fr��~��B��'����旟�ݥ%I�'���,^6�� g�V}\x;.�2n��Ī<���?����?	��?�.� �C���+�	��ܨ@���[!Y���yeG�ៜ��ԟp&?�����Mϻ
bL�I�*(�B4��
h���?�J>�|�t�
�MÜ'���qH�s�L�t��2���r�'��a8� �ş� Ú|�P��S��bH�?��-z��[����l�؟�����`��_y��h��D��M�O����O�� �N!��\`d�@�nV�42e�;�	����O��$ �Ĝ"?Fz]ؤ!�)&\t��&ۙ&��ɊSdL
�	�3G�b>MA�'M���ɩ\.���Q�
\.XL�7*Ӗ��	�����\���O��`F@��d�V�M�v�P�VOD�sӜ����O���F��}�?�;#��3���1I��$���	9r	����?���?醬��M��O��@���O�1X��������u�@�0���#gf�O���|���?a��?�����9����h�q1oS�4�*O�o��z�'����$�'^�`�t%ȒTNB�xU'��+� %H5b�>q���?YM>�|*2�
�?Z�hP�M�B0k�Jɍs��7��o~�����\�I+_�'��ɇ�n�JР��ch"y��L׻�4i�I����֟��i>��'�6�<}�:���M�B!��J����Q�Yr�U T�'�6 �I+����O��$�O�����I��d{��G�T��q�&�)�N6�!?!��WmBb�)3���U�3������uǉ6m4jD���i�$��ݟ �IƟ<�I���󯍋%}f4��n��a��P�J���?i��?	��ib섻�OL�j}Ӑ�O6�3Sj�/-斄�B�ךt������3���O<�4�丣�L}�L�L�l�
�*�oH�Ҕ�c�v�J�J��X��U��䓊�4� ���O��DՊa���eѻU�2a��jE�=5����O��9e���0�r�'�R>��.Ź��xi��b%���J#?�V���	蟌'��a�.D�@�Ҏ2�,���ʝ.�N���H�&�B�9��o~�O[ȑ��%^@�'�<3Fn�S^<�DdER(�˰�'���'^��O�I5�M����!�r��E9T�a���	�Z����?�&�i��OHM�'r���H86�*r�(�Xb,�%���'���90�i����M��0W�O�n���Ά�&H	ʃ����E+^�D8h����J�(�A�C�8a�̃�;v�ɅɄ��bA��!{L�Ie�&?�t���`�u���$Fـ^�V9��T��(���WVν��K��"�q�Ë�G�!�Ŵiv��L�h��A�͜8�9�p��ܼ�av�M^���!#��SP� N�|����DΛ6&�����
^�\0GQ�Gt����Y2d$&��y08��4�D0Z���\���g`�g@9uEB&v�QQ\��C���m
"0��kC'1#z��@d�A�4]t��6�4	�4�?	��?A�'Gb�O��( %��f.� �֌J���ݦZcD%�S�OAB�1� �!Z�n�O� �c&�c%���i���'|rj�
V+�O����O�I���@�5E
>1����į��{��b�P��o0�	⟜�	�x�#/�:.xڭZ�ƍJB���C)�>�MK��e5n�1u�x��'Kb�|Zc��w��;��}�t�)
�䚯O��9f��O����O�ʓe��8�ް:��L�h�p7D�˓��'���'*�'��	�Nخ�y��!;/�%�sj�(���`��7���,�Iҟ�'C�0z�m>m�1��,?�r��a R�+ 9@@$�>���?)I>�/O���T��"�:o�`�b"��9Fļi��>I��?�����%L4&>�򃟁?���M�?����,��M3������$%Y��OΩ!uJ��
�
$C���6D�Uz_��L�I˟��'Q,|PÄ4�	�O����)I� �+i�����J�2wBd0	a�i	��tybN������s�ƭ�.�0RN�A*�i�2<AHT��i����ڴ!o���h�S����M.C|��hE(h�Qd�H6'N�vX���h*�S�'B��9�d�1�Tպv_�%"mZk_�� ޴�?����?���zǉ'ψ	o=�9���e~"�����)S�n6��c��"|���tɕ�52��Yɠ�@�:��Uɑ�i�R�'Rh_.*�Tb��It?!��?6D�VOϺږ�QL�D�V�jt�<���?���86���ńBXp=���!a>����i�R�4��OF���O.�Ok����S Қ�>ѩ������I����	ey��c�<��)һv4��3�A�'R�9ƥ3��O���/�$#}�#gU�0.�|��3mK�����}��'���'��I%FB�X��O�P3 ��J��Oӵr ��h�4����O�O����Ot����Ŵoq*H�C�GjLE`sh�>	���?����$ݦv���O����xI+��e_hE�v�Q�E�7M�O�O��d�O�t"0k+�ɛh~��)`�ahN�� �+�06��O:�$�<Qc	R4KF�S۟(���?y)b ҰR�鹖'Kc`�g�ˊ�ē�?!��	{�M��ҟ�u"أJ��(H�h]+c� `pP�i��I8Z �4�?1��?��'d��i���6��+Bav�U<��m�����OZ5�$��O��Oh�>!;AM^�'Xx�d�<W04�q�~���Q���˦	�	͟�	�?�a�Obʓr��QHg��ag\e�ˇ�g$�DI��i9,Y��'��'�����U�*Ab��#�h�"�聪U�o��p�I͟\ A�ʀ��$�<���~�g˅^�8(�S�UO��F V���'�0���y��'���'ze��J�s��m�抒6�}�4�zӒ�d2��\�'v�П%��X�O��=a@��Xo.���_���x+�Y;�����O����O��$t:�㌓�/q��@�:sM��[�B\(T��ILy��'��'���'	�E��/3�ƨ��� 3!;�-�cM�~��X�,����	by2��?>B�Sj ��3��K=>`���d]���io�	��%���I�PRk��X�0i�;o;x�h�Mߢ�,=X�#6���O���O��PCL��Q?u��;o���aB>ao��sk7���P�4�?�N>	���?YA]���'	�%2���*3���@��)\@8��4�?�����Ĝ6{���O;b�'�������),WQ\��Ϥ_����ƝxB�'��|%��?��OϲT���,(��IC@+<;�p��4���%��m���)�OZ�)^~�!�/��+!��*2L�%f��M�)O����O>�'>�'?7��)�ĕ�1�rZr��#�k!Q�iRP�"	hӖ��OB�D��%��S${w�e��J�yܠWA�%&}��i��qSe�'��T�d'?�	ݟ����� $��.֔��@���M���?	��>枌�x��?��'�zճ ɜ@�{�A�V��ݴ�?�)O4�rZfb��<)��?�z���d��>db!��,ݏ��`hD�i�ң��d��O��'�ɧu7�ʷA��Y����;�aǟP)��_�(!�����?i)OP��֚'/���Ʊ7�ZYsC�:$p�����<����?ɏ�'��<-P��h�c�~4������`�j1��'�2Y� �ɠx=>��'^����&X"��9J�H��8���o�ٟ@�	f���?����4�`HڦA�IH6�#�) f����8��OV��?q�ʸ����O�A �[N~�0�AT�R�]�F�e�?Y��?�Ʀ]�.���'��ÁƓfKDu(�FֱD��
�r�H���<���"��(�����O8���8=�3H_/o�����D�#Bp�@�x��'G��>s���y�����CN��@��F��*@���_�X��,,��������ǟl��XyZwe�Q`�`M,_1씳��/¬!�ݴ�?�����ҬGJ�S�m�ks Ϭ &����I��@��n�="`��4�?Y��?q�'����4ЃO�
ႁcU�R����K/@��ș�V��'U�	g�3?q6�
>V%K�Me�a�@$ϧ|{�&�'��'>0���_���ɦ�"�*U�ގw��}`�)�
-48���y���-�������O��U�JP�(�//l��RW��6/(Z�o���*p����S�	N�I*���� �*xD���G<V��tk�O�:&�O��Or���<��a�� `Y0��^5���a�E�dzn��S�܅����O���'�����	�T��6��>O����吠g�n=���#�c�<�	wy��'�&u��ܟ^���b�nv�QQ*�76_Q����?I����'��'�<j�b4�M��j¼R�bt��(�/6���I}�'[r�'&�IR���M|�0�_s,i�f�:]]�U��
�f�'��'?�(�`�Id�iW8ی�OT?E �0��d���'6�W�$�E�
&�ħ�?I�����;$P,;�$��a�^Y���}�	Jy�ą$k2���џ�Z��N�Z�E��ܚdܤ&�i��	{�Ԡ��4J������ ��dF�3�h+���n9����
��R�t-�̟L8H|�N~n>�� +�?�h���N�%d_�7mЈOD8���O��D�OV���<�O���S��E�l������	)���5g�$ț�HɈB#1O>)��a�q6B�'8o2���C�Vv�!`�4�?����?Ibn�1x���gy��'��DW�p	��!�4[)&@u"�^���|Rj��yʟ���O,��(4�ݡ$�8��` -�z+�9m���\�Q��=����<������Ok��IZ���R�׼顒!C�I$;�"�?Y��?I����DF�D��TmҨW��i��� 6�����Ni}^�P�Ify�'�R�'��D�ɾ�����N�  
|��K�#�yr]�d�I៨��uyȉ�WR�ӽib�<�d�F+�Ⱒ��ÆpeJ6M�<a����d�O.���O���D9O��q��S/0��Iu`�>i��8��jѦ}�	��	؟h�'�Z�3��~��O��L{1��V�P0E�f����iNS�4�	��<�I
R������jd����3E��PG�ڌcP]m��$�Iuy�C ?Z���?������T�	/�ЦĀ�b��iH6��G������	�\9j�d��qy�؟����I)�����2i���9��i��ɮ
���ݴ�?����?���C��iݑ�$�.W�DB ��=�bU3v�p�����Oj�C䐟ȗ'!q�԰xQ���IA�dܽe�v<�%�i�܌�aJq�D�d�Ob��$�'��Ʌ����A�5��uIf�ޑV�J���43�*�͓����OR��7/#�2�EV6º�`0�Z-o�X6M�O��d�O�x�-�K}�U����N?1agR��:��B��ȰⶤU�A�	Gy�Ь�yʟ����Oj�DR�eV��lN�S.<�Jv(K�X04`n�Ꟍ�%��$�<�����Ok,�c{��BfF�0��<8�'���I�D��	ɟ����� ��ݟ��'g`��Eb�N���hgD��h�"����Y� �����O�˓�?Y���?��œw��H��d-�К���m��?A��?Q���?�)O0�j����|�"�J�%nlyR��U�����ئy�'u2\�|�����I�a�N�	��!{ş"����� w�p@�4�?����?�����D�C�,|�O��5d'd�)�`$#iP,�@A�x6��O4ʓ�?����?qU���<QH�l˱�֗��`��!���e�e�6���O�n��v[?�	ȟ0��Z�p�Q�g=tlp�	m�����O��D�OJ��L���	Vy�ןz, �m�o�X�I@��aoej�iA�	�/�$l`۴�?I��?���qo�i�	���Ǣ��Js���\4��B�wӔ�D�O�#9OP��O���,����e�� �;o����ǔP�D7-� &��l�ޟ��	��������ħ<�LM?���5%G!HK���3$��J^��yb�|����O�ܲǭ-g�E�N�F�x�笙�������������(�O�˓�?1�'��CK�H��5��%�5>���ڴ�?Y��?�VO��<�Ow��',�B´%}*�����>BV�*c,!Bf�6��O�)x�GJ}�V���Ijy���5f�ʕ06rĨ2�ːl*`҈��A+0�$�OD���Ov��|Γ{*�5�E���"�i����yA�#$��	y�'[�I����	П\�B�_�Z���Cb4�Ĵk�m�}7V�	QyB�'���'E�Ic�D���O�R��b.�$NR���h�*�jڴ��$�O���?���?Yq�L�<��N�"J�aˆd��e��#
�v%��'���'��^�$��@C�����O 0��\4�T��ձ��#�Ħ�Iny�'5r�'�^�A�'c����Ѕ���&�L���ix��o�şD��Iy�P�l�'�?���*RC�l�X:dk�>@�0�hj� 8����	�Q�$��4���2|� !��N �dǇ��M[(OnX[�`E����������?M�O�NK�8�IÇE��Y�/" �v�'hR����Ĳ<I��4�A�Um��!��+A�xh�띯�M# ��d'�F�'��'����>�(OJ�:�jJ�C����P�n�0Q#��������w�'�@�:�
՚�@��l���ۑGݫu��m���i��':�B�$m�����D�O<�	��l8����
AB<c��7�O��#����S���'T��'�lDA�eYU\R���Hٍ6����zӴ���8Yv�$�'��I����'�Zc��)h�KC�L!��a���%��M��4�?�J��<�*Of�$�OP�D�<Qe�0NbMjVc�@�h���l�����T�$�'��X� �	ן��	�xB�%���F�)S��Ό/
��ce ~�$�'�2�'��T����L�����N�����<I<`E���M�)O$�D�<���?���Q����'���K�a�)�y�
�G�t�Hܴ�?����?�����MR��O=Z� �qp�|���֧���a�io�S���I˟��	�-]�IO��.��q(FaQ��������= 7�O���<)�bA�zىO?R�O������Ђ��ҭ�tl��!=�$�O �$� 5�<��?�Z���au�"c�Q-<� g�{�V˓3�-8ֱi��맸?����O���v�����l�R�9XXȶ�i���'�P�R�'��'Rq�T�3�)Y�m�"��$D�����w�i�@�`}�<���O��d��'����8NO4����H.��9�Q���?�`��4|j0 ������Ob�G�o�s�����I`�`\Z�6��O��d�O�|��@TT��?��'?����
^�J��a���<��
ݴ��v0�������O����OkZU��Pwɀ����g�î����'�V(���3�d�O���<A����@(D�H��i�#8�J)d�i}�)��aZ����D�Ihy��i���7�T:12���B&A!�Q�F%0����%������ث���	a����jDHhr��'F=,�	@yr�'���'剈x;��y�O!~	7�ز@A��@!�0���B�O��$�O��O���O�!�51O���Qb�
6Bb�zi@9��1��-P}B�'-b�'��I � �sH|����T�贈�,�(g�����k)���'@�'���'y�p2�'7�04dI��Aèt�AY#�J8��8l��h��`yR��Z������DI��-��Oֶp�J�<;�\r��A���L��9y���W�	KB��	$���`�g�VR��X٦=�'��m
w�@p`��~�����#��|
%� ,"y(̐`)Ț*L:,ӑ��f��O������OޒO.�>�c5�l�~�N	�7(0�~Ӛ1)��ϦU�	ş �I�?u��}B�?r�$X�烚�an0� �@!�7��A��d-��4��ɟ ���\�r� k҂�Y��XT�ʈ�M����?��{�Q��x2�'���O�]��'C>[���PK@5"nX����i��'ު�
B�%���O���O���ec&z��!V#N�w�����G���"Ih$R�}��'�ɧ5օI�v϶�#!A���#� �����ȥx}�d�<A���?����^�zĐV�M�Z!�Y��Gǜ+,�Z���L��Ο\E{b�O��Z�o� @��� ;r�;#�i%2Y���ҟ���dy�훽u�b��57��Pa�X2�m�@B��,Y>��?Y��D�<	�?Rx��gB7d��Ѻ���~2�U��Z�$���P�I֟��	�j��	��p�	<�⁢��  �vHJ��"+��3ݴ�?�K>���򤍥Sb�'�0!�,��G3���KŶ��M��4�?������AR�'>}�	�?E!'��3&�ܙ:�jZ�@IC��M{�«-����i �l�e��,<g�r� x��+�4�?���J� �"���?�,O:���O�������$�\�85X܊�9ŵi�2R� ��2�S�1:[ЩP�)@?CK� 4(�Xg�iL�YwF`��d�O��$��>�'@�	t1$!h�͘b��u��e�>�]p�42!�Γ�䓅�O-ҡ��D~�(�m
�,2< {�耉w6��O��d�O8%��n]B}�]���	~?Y�a��1�V�;�&	�_}�-�G��æ���0��>J��)����?��eND��9q����b:�2�p��i�"K��JP���d�O�ʓ�?�1��x[�m7�J
��39 ���'�v���'��'Q2�'nbQ� �ddZ�;P���P�
4-+,� �ȏ�;���O�˓�?�,O��d�O��D\#PĐ�ꀳ�����уT�h$�q��0��ퟄ�	ٟ�'/��c�Mi>}q��R���)-�-��	͛��7-�<a�����O����O��9rU�D����X���C�� }� ��G|Ӝ�d�O��$�O�ʓL�X�a�[?��i��i�j�y�^鰔��Mq\H�0�{Ә���<���?i�h�(ϓ��icB��֔�~p�c��~TD��ٴ�?�����ď��O��'��$ �Jt�g��B":@	�B�#3^��?���?�PN��<!/���?)��	�\L�t�K�k)`�y�(c��ʓ�X�6�i�B�'���O,`�Ӻ�V���<���0��Of�H���d�Ȧ�Iٟ�*�~���������_�']�}K`g](y&����ƨ8�n�J\�TP�4�?����?y��vI�IMy���=7� h�	�!���0��'z��6�� '���Oʓ��O��
� ��\��GN�w ֠�o�7��O����O:l)��u}�W���	y?у�Ӆ.�z@��Y<w��'��Y�	ϟ,͓�0�)����?��O$isS �W��e���Ӛ:$,�бio⋏,L��꓍���O>��?��?{v�˧@I�;��Рk[�j��m�̟4K7 q�L�Iޟ���៨��t�4E˥Q�h�%oX�`$�@J]� (� �[���I�$�Ik�	� �%:^�аi�zS���,�.LM��m�a����?)���?/O�qs��D�|2fĄGkZ탧��<�&�E@}��'n��',�O&�[�]?i@�%�(�r��儀h*��k�&�>���?���?����&�����?y�'Y�@j���NmAE��#os��ݴ�?�J>A���ԕC�'k��A�		2��*�֭���e�>"]�O��}� ��k �@�M��Іȓ�H�@��ԗFjN\a2�ݸp�l��a.��G�\U1dFE�!s�œJD/�z��4LWIJ�ysdY1c�<��,�F�? 0@�� ��d�h�JS@�#��eɀ�	~:X��	�q�<Q�Q�����!&��P��Ћ�E��pŉ�V���$��4X�*A�}�f�!�(� %<$X�І}�����P)w�X�[���?Y���?���u�[�q��E:��M��i�f�9rf�f	�����oV�o�.l� �;擒��I1H8ؐR��ȃ,N4C�ٵZ�����D�5�Z����ȯ*�����4��w�|i��'� 0@UH�L����/�R��(2��'���$�4�4��=q0qF�(��Ȏ_ђ=��N\@�<�6�@I��,B� <	��� .My~rI>�S��P��b6��!�}�K֭8�0h�"�#1X\��"��ӟX�	̟|�I�u��'�5�d�ж��;*iFy�&΍#���`䌤*"F �c���g>X��ɜw ���w�@q�5#J ��ғJ�Y�c���=Ab�Z7'6� v͏�+@ɇ��'s����ޟ�F{���2bưtc��9c��4h[69�!�d�
=A��
A�>[j���\g�1O�%�'*�I�k  K�O0�D#7� ��5Jk�9�qgK�_�V��O0%I��O��di>�i�*��K,�ˠC��~���b��+�Xm^@��-�p<	���4g 	H"�#D��DҋJ`&q�w�9�&�S��".��x��߉�?	�����/a��Y�nݱ%�$@eF�i1O���$�37�i�B�I�)�$���F-g�!��\�B1	�)m�D]��oqU0eG"x���'xd�ʷE�>����)֟l�`�$�9���*D@͗0����3b�6:�2���O�<pp(S���2���T>��O�f�J�a��f��w�	*2�CL�(�t�c,�PVLZ7먟��@펅���1�*3<}y�>�Ac Ɵ��IL�O�?h�Ԭ�Eӯj�8�p�!�y¢�t���җ�vx IJP)�0<����<RUv�Z� �8ts|�0��ٸ.�(�#�O����Ol0ApfʇQ;n�D�O����O��ʉ7 ^�P�H���n,��JO8gpy�F	#���6J�&8�p�*�3�$[�c�i6��7��Y�DD�(l�9'��P
�-�	B8������|2A�Ey��K������٨!ҝ������O�=ړ.�����+uwf\X$��h�I�ȓӞ��D�x��Do�x�t�'�#=�O�I�G*�a�E��8����7Ac��@�W�dL&��f�'���'d­g�i�	��8ͧ�L���M�E ����,o�ta���12��f��XXdXkE�!O@t9�E>e��\a�i�� N������*0d]b�ʅP�Lx��3�p<�E���n��	?�P�c�/ITH6����M�w�i��O���~��J�$�� �-[J@���j�_�<y��J�RB�hI��NÈ�{�g]�1��Xy�P�\&z7��O���S+); ���G�y��iy�gۿIWJ��O:�! I�O����O"��-^�V�x�`V'~;b��M�pS�Uy�#O6
z:�z�F_J1�xB�^�,��haC͍�IE��`P�		� qiV�O,,8�W���XÓ~b���۟h�ܴ�?Y7N�?ɢ�AA���j��Ig.ъ��D�O��"|2�N�al��
�C�~��$d�hO?�޴c���Iab�� �8��֊G8Mx��hOV�=9�#]*=���0T��FD�E�&#�E�<�V)�7j?��h�E?����*�B�<9���*6F됢 
��\r'|�<�F��&$-��i�B�d��A4c�]�<i�'�*;Ϛ9х�A�p���o�E�<�b�.:֜{����Q�x�$��}�<��O��������W��В��R�<	�1Hl:(*C-�2�l�p�P�<��NI33���j@� ���E)�J�<�Gkߕ[�ԍ��)_�},����C�<��G�It��Q�`�07�~��Q��B�<�	���
�!��N��,��a�E�<����L���AY�a+x�õj�C�<��*&g,	�i�6�-Be�@�<A��g��q*T�8�!l�G�<9��-=�dD��k<0�xQ��f�x�<9 ��9�"{��^���:�B�q�<���;��u#���~I��j�*�E�<9&�Un�}
aD��� �P��k�<q�ܓ1W � a�߇a7�}��Gf�<�5k��	�;�`\-j�܊DUe�<�'I�8'@�-Q��ʭI�����|�<� �g �d��Kt��5EkB4�2"OF���� 4�l�"O��t���06"O�I�gƼ>��{�nD"~��`��"O�`�Ǖ�}#J����{Ŗ] "O =@e���L�S@��P����"O*)�A��ꁻ��[2^L.�0�"Ox�y��V�����`L)aG�y"O8���"��N��X;�.3#nyR"O0;��j����6
P\Kr"O�8ѩ�w�p\l���Z"O�=�cJ�'!�� X%��"�<��E"O4!��Ή�fF���
��4���"O�tЗ$J�a��բ�]�)���Hq"O0�)C%��?[>�#ǩ\6q碀�D"OL)C�)��]����K!�*�
�"O�P��,G}�n���U� �8�"O�c�E�g�]�G�W�?���"O^�a��Ҍ�<�Z�`K31E`H�"O��LH����p�N�v/��"O����/�=~��4O+�2��U"O��b��L����Ĩ� �`p�"OXYyW��o*��.���A��"O~�x�@�q�uY�-�4l�\�ap"ONQ�0���9��T9B�� �R���"O�<�B��)S��ۥ��c>!iG"O�H����EA2�9��A�P�&0u"O"q���%]�� Rg
�)�4�j"O���S�Y�����#t�H<�R"O��ZՁ8�h��L���u"O�\K�Ƌ�t������S�"��m�"O|@�,='����.^��7"Oz��Ҏ\�PBn�#rl��j�8?�y���M<�x�c(S�\��ixg`���yrg�=̮lz!%��BZvl�G��y"*Y=n�����h�$�#����yI\�F��:4f0Yi���%�+�y��e�fC%kI�JH�4 ң�y�h͋2}�lz�';9:Uq���y2��z�صjBZ�-���vL$�y�D�23J��u��z�+P2@:*������39��/�B#��e�<)��2�Đ�ǥx�	�'Cb�<�¡
3zO��*b��v�v�pt]�<ɓ-&1�����M�cJ\��e�Y�<YЏ�0\&�I׆ϵ�r=�'R�<�J:���'�'M-�գdI�W�<٥��� �v�kdr��˄��J�<�1AB/��D���")	&�	r�<���n��-B5+��en8�T*	g�<��<S6F���Ǔp�Ę�3�e�<�F���t���!ɹ}����fă#j<)
�}b���U�+�z��p��46�p�y�9D�����u�8�b"�� ���)&��OzpW�R/��>�Ag]�e���0�%e�@� 3��h��pv
�6��	�GK�����%B���b0$W�W�B�
#��8(�n�i<⁩��1�⟼�f���4��
6z��"$K�<`��y��"O�<R��"'����j��Y�A�O ���)�'�$����ö�SK$>u����'��BO�;j��u�Q�ӠRَ��OƉ�$�5lOf̹�"�: g"٫Pi� lؐI�g�'��yڱ�iKFE�Kk��[��_��5�'h��@o��V��H���@:��FK@�y*�Od�7���'P��47�H���?E���qg#P<s���d"O� �2�%.-u����.EWF�05�@(7Wr��?����.g)�6���*�S��ʱ~H���"Ñ�]��09�M@=�0=�aH٬`b�������<郎&��� \�e+N��r�ί>(�@�F�<}��%6R���'|�1J��˿0�.���ؽl^.��<�e�ٿhV>��@ga��<�;h��{7!�;*)%�G���*iΓӲ���H�d���d�
^�l�d!��A3�Y9'��)S`6����W:D�	W��b>��B-3fPM[�gw=h`5�� `��"1��B�I:yy�C#�*���2�Z�l�d���90������� FN��� ��>�O�xD�8Z�bEz@%�>jT � "LO2��a�
=:�8�1O�TJs��)l(\�* T�L�l�Q-V�T�ȹ� Ν��?����P���'�Ҷ�T�o�,���ވWYxP�y"�ߊSQh!so�"�(��,4E��#KJCȺ��`�*�@UȂ�_r$Es��=�F���L�z��WƏ�x�8}x�@�)�����tm��2
[6�ӛ0�|���˷w�p�4�T�:�TZf�[+�F�;�+�P'\��@"ORQx!́�XT�U����:G���/��h�ŅZ�\�p�l��*5�P{'����M��g:��1���ʊ�?�|�g�_8a���DݝP��sF/����d� K���Ţ�5_��asC�$H6�6Ȁ>8�JX��4,�(���9�3�$́���C����r��5ពc�1Ob���។g��<0�ӡD+�����;8�!���*%<5�V>a�,�Їo�~���ד�|�*�(]#-����G��_24���I����p�˗*o�iK1숿QE���]C��C���$ֺ|�	�'~�l{B���cI��(���&hjH�N<Un��PՓ"����0�����!M� �h�h�YZr%��j�d�!�Ćb �P�iαM��	��@���&

>%]f��'>���>)��D�PF4�I'��]�����Oh<IUN�#�АB � 	T(y�Μ�d�$7�Q-z��a�.�:�p=iG��M��Q�bö%�ЄťW8��@��Zl����)�ꟴ����F �m�BC�	����QV�fP��s'�>]4\B��*q�t��dKP���;�]��'��U
f�	S{�%�͞�8;����'���37�Г}��a`A����J�	�'Z��3��	W�"�����0��P
�'V�k W"�<T���%&�<a	�'���2W�ʔg]��Q1�H4�	�'ƖQ��G� ���ql3���yrj�O�	{P�C'�}:���yR英QX̸Z$M xw �C��'�yʉ�^���E��>>;J��ϙ;�y2-�?KEj$�@?J�h��p)��yb+�X��Mc�%M�v֞1�P
��y"�Q):��)�ƚo�I"�6�y�R�~� L�8m�.�E�ɏ�y2ㆀ>t�h+b��d؊��W�P��y�ă�8����oĕ&&�|pW��P��|��� h)$d"a�=aA��D+X���'b�lR"�L	��B�χ)l�z<(����q�O24١������I�.���)�"OtE��c\���M���	���6剞j�deË�I֗h1@�h��4P_JȂc��0�!�d�����ɦN�D  �J&%�6��� ��ا���	מ1���ɟ#Cb�*Ud?�yb������R�L%V`�������d�^ma}�O0g�XP���
�$$�{a�ڕ�y�k+~�I�f�h�|݁0��y�,�����.�<�vlή�y"�8"~T�bD� tB�H[v�P��Ċ���|
�5p�<�� ȴv�T�rp�u�<�',چW���)����P�,��Oo�	X���ɚ?<��f�������$�]dR��$Ԙ;4��r�A��^�tI�툅&�6��P4D��p�I
x��v*#y�I:T�=�#!�]P��	�(T&��b�ѕY���D�!�dF�����j[&[�Z��3�剨i�|��?E�� `4{�+V<�:`:�*��[�z$"O�u	��=\�"�
RJ��	4
�|�J��<azr�	%Oj��@Ч^�O� A�PI̛�p>A�aB'5g�}9���?ð0;��0g2f\R4�� m�(B�ɫ
�b�I`� ^�RT0خ�<q �۩�r#~"��K�� ���/oc����D�H�<Iq�C�~jhL�)خX�����H�o(d�'��F�S��?�����ۑfM4a_|i!b��(t�C�	�u�n|�t���X�&��R� &��I�Ou�䢷�'��m� n@�IX9p`��������B>v��R�v��%���@i2���HE�`_�<���5D��v*�79��(��U��z�`R#3�"="-��*$�NF�H��'r�$��g�"^�x$��/WrݳQ��*"IE!�A��
t��%�?}(��=E���jRD�V�H�9��9�gԓ�����T�����d8EB�< �l��~E����&"�O��A�;4���3���)��'o�a���d�P�O�}�F(s惝:T�0K'G$D�s�ŖRB��1<|����4D��5��|yB�0ʜ�t�h��5D��SQ�R.ٓ���9����BE3D�4�c Ϲ<�F�C��>��xka�$D� r� �i�1��ܥ}Ǭt��"D�$�2�۽U)�����d�%D� �4$� 9�h�Z_]z�jg"?D��P�f�K��t	�Zb�"�%?D�,�q��}��]�щ��o,ZH�<D����@5T��̀Q�ѡU�d�9��;D�,����&r�"$)��>IzB��SL%D�(��X w�@�(��4�t@�&� D�8��#�2uET� D����i1B D���#W� q�`)p���2R�>D��+��D�T�u0t���U�� 	<D� S��
D,����l�6�۶�Q?�y��H�^�>;���\�\����yBK�	QF���6�A�M7���S���y�%/GN�Q�
/JI���RM���y�a�qT�A�b�%A�\XX7o��y�'�f�HX�i�=��lJW��y�E_e0*{��
>Dˠ��M��y�d�h��M�$�Ԇ�t��%��9�yR]�m�t�u�N�6�6�x"�J��y���(0� �
.���e���y�l]�nn�x㴧M�Ü4���ް�y�,֊M2��1f�J����d��y� ϑkm�Q�f�.%�k 9�yb��2�b�jṕ� HluO��yb��5y�<���N	SX4%J$K��yb�)Rn��Pp-R�~�>�&+^"�y�O�Pn�
1
Y>Lͨ��V�M��yBnSM��dXJ�;IB��RcmB0�y�G�6N�eb�Έx"���=�y2"�]4&=�1#ոwG��ID˻�ybe�mql=�b�Ib�.X��W�yBȜ ������Y A�R�y�OT#']u�2��R�a�#0�yB�{wl���\)`��mZԧI'�y"�I�K#���z�B�o��5�ȓX�"�@�c��Q9�(�����E:����8���1A��Q(N�B��Q~>���8����F��1�ΰRA-��0)t�ȓyx�)����W�T��'�%D��̇ȓ+���;`�܆+�΄�7�P$V��%�ȓ_����)]q�hY #�U@�����S�? �QC�朮yJ)�2&	<.u~���"O�Ec#��yX�Ɣ�kӤ�2�"OҀ@E��<������%O�J ��"O@�8Gk
9i}b �nˁu]��"OF�C�MJ
F^z%�'G�p[Ҽ)�"O�1@�U?L��g��EI�S�"O:���	j��5�&搓j!"�"O�<R6El�N|�ŤL"Lz���4"OH�LO<��$�c�5b��	�"Ol��c&d8P�8�M�j4T$�"O��ꁭ��� ��S�3�`&"O�Xz�LY"8� ����8�"O13��dG �s̛6q0Y� �+\O�e�w���}�׉�	���2�"O��v J_F����A��j�;�"Ov#�ɇ;�
#�ӯ�d��"ONݻeO@/1��PeA?8z�"O�EcЂ�<=ɪ-��O��ӑ"O��q�`@��@h��
�s"O�Luo7I� ��J��)V��A"O�3���#H^�c�H'�"��7"OV���2CP�Xh��"<�l\xA"O�hRe�C�:8�F@��o�`%"O�1P�M�A��`aq�_!�����"OV�;��B�i�AHT'ͤaM��P"O�9���V�	�PQt��?��XP"O�  ��N:�j�p���\>��P@"OJ��%�B� �>��v��z:pͩ�"OF��a�B�&���Fђ	)D���"Ob@:��3R��H[1@�"$
D�"O,	Z@�U+���Qn�3}�~���"O�0j���w=���0�5K��&"Oz��%�ߎs�-�S��"/�X�"O����ԗ����3�C�K	.)�՝|��'�MiS�0i �Ie^�v?�(��'q�Ȉv�֧JQ���"�ʠ^�%��'�Դ�N�>�١�'K�nQ��'$���� �m�)�� 9
��D�� ����
�3{V ��ȴM����ȓp}$�1VS�R��Q��� ���Pj��C4���d)@���F�~|A��oY08��c)%vD]A$�	�ޒ5��TM2�D�2j�}óCʜ�b��"�Ȑa!�_�*P���E��)��̇ȓQ�@];F�%)1t��3��1�:Y�ȓ@{�X�)F���њb�#�dՄ�`P0E!!��r��
��G8�̄ȓ8h$����( �FԻ�g��^� Y���]i�H�-���y���j&r���u�0��t-�e���k�
�{����}�މ2��F�Z�kV�/#��y���t�M�|Jtͱ��-��Ą�U\�꒱���Ō�>U�@=�ȓq�X���0;6�`���7�X��ȓh��b,�B`
�f�"�^�ȓb��8rW�Y�5��m�#� �}�\%��rf�H�PV, �.8�f*�r9�ȓX�.�_}�(�S`�4$��b��y�C-t;�R�
=(sd�v�<�δqZD큃j��f'���
r�<��&�3$���f�N�%�l�KOp�<Y�ٝn,�.C G�9Jǘw}��)ҧE��03bO��*�$���94�P�ȓ93�`bdX�̔;�Ѥ ��S�? X:A
�,���۴*�MȆ��6"OJ�a6�V��u�QɚU��P!"OX�Y��R�QOp�9�Wx�|���"O��vk�6X�0,�Ь'��`2�"O�� ���s�n�ꃱ�R��"OY��G^ C?��p�,9Z&����"O�9*e ǎd=옱ա�{k��#�"Oh����0=�����ߑ�$��"OT��#�[��I*��=����"O`\D�� /'T�*�E�?�b�C@"ON�aP�՟F�2��n�Q��u+�"O~ {�QA��kW�@> ����"O`E�$�I�P�,�c�n��2E"O.�҆6��{�׎/8Y�"OR���Ƒ6���F�ۑ#кE��"O����E�NZ���rI�"��T��"O�Q��[- ����Ԋ]��F"O�Y���ɗ'���0I��U����'�󄗰`�� �!�t�^�ؖ��~�!��)#��A%A
�3~j���&K)�!�D
�nR��c�ڀb�ѯʶ�!�䋒*�nql+m`�%I��r!�$(Jz�rd`�!���c�H�!�$��I��Ȕv�*Lq�aZ�S�!��M#��s
��	��К��F-J!���
r�}Kn�|��U��/��XH!�C*T�$34@]�,Ue�&,C!��s��E��4K�������^Q!�䍨^K�� �CB
m�`e3ĀG�Nf!�A�fX�B�0mk�`{���HJ!�ē�B��sB�8|O�$�2<!�ă��E�D�Quj���Gb 	7�!��6G^��ǥ\�hb�󃢍.+P!�D� o�Kħ˺Hy$Ă��ݐ3!�D�	$�K5��L��m�揊�_!�K,r6���Oėac�Ԭ�	G�!�J?h�~T���^�^���3�A�*q�!�d �v��Rce9C�A�'�C%!�	�\^���%D-l�]��c�@}!����B�.áGј�k����l!�:2R�B�!</ΆH�+[d!�D�0/�6ѢEo�nV�J&���t�!�����fgM�Z��L���5f!�Ĝ"_�>cQf�4
 F�;2�!�DT�u�����=�X�k��ާ:C!����q ��ǹ
2@U�G��Lb!򤖮ClX�8�f	xY�@9&9!�B�j3(���Ȩ$H0�#4�C�A!�d	s3"h�Ƌ�o/&1���H�x!�$��J��p&Iʙ[L����)"^!򤊝O�e��oZ���d�ư`6!򤔕x�b��'K fƉ����)!�D�AkZ�Q�eS�e�D?
v!�D�LMx�j���' 2�!�	N^!��ד��jb�
D��	As��mz!�ޥ��E�"���{O֍�"�v�!�䓢Q��hd�R�\�(Hk%� �P�!�$ʲ3V�׋A)o�H���J�6j&!�dN�oHf�S��	<�ĝJ��g�!�dϠI-DE��l���԰{a	֧_�!�DJ5:�0��-�.����nԶ�!��Z%H��(�Q�O��I`��κLr!��~$8iF�0?*�X��M� c!򤋾\s����j#jzn	(��E�'!�� .E�t�b���4g #7}Z�"O�e��M�&W��T
Q�Q+(�I`"O�U0��Q3%�ąQ�ԭ3�؉a�"O�9�H�B�L�A�ݕ[ޘ�B"Oh�ň�Kk�Р�l��B��v"O�Pv/�bN���0kFx 0р"O$�� Z����d�d�P����C>�[v���I�R"³>�Z�;R�5D���`@��F]^�0tK_5x�<u#��1D�t*�đ7o�,���b���D%.D�����ei�y�T �B��0��F0D��
�Gڲv�l�J����g��+��3D��c�ƘJ4��ʲ�R8Y�Z�;"m�<��y/ mj�������O�
$FV��}=���/�4��:P�G��x��B�����A#v(�@^b��Ey��'�J���+z��p1��98�P�'�f-K�Oߢ:˦�P瞣 �pI�'Ӏ@cF>�xQZ�J���0�'�F7]�ޅP�N�#A�4��"OR|j��PKH�Sh
�G�h��"O*`Ŭ`�({�'�%7���"O`����2)�*1�tD�.���"O8Ui��	uRp��F�r�`���"O \�E��g�8��'L���"�"O
\ 
���,���^u���"Olգ�▔*��y��ݹ
��ӂ"O��(�e�*$�hQPc��Kf2���"OT�["���)Tx���#˿0S�tbs"O.kpiM�q:JEbr�J�[M6�3�"O�́&$�>YRᓇ�ę�"O8U2��N�6����-����'"O�T��B���L��1C	;?|�x�"O�ġ��6Ph�	X�P� "O�p���D�z��q��1r���pp"O$����[)tg�@CgM�R���"O��XWdB f5	�eV16rd��"OxY2��Z����D�u
�)�"OF02�Ϩ|�p��ף��5�ĵ�e"O*ERg�4"V�[#�#f����P"O\u�6CT:]���0�B)b�l�{U"OЌې�^�*�h%�D`�t��y�w"O�1`a*L1y��cpȋ� ��"O(�q$H�</��Q�U炔GV�"O���]Z��WOb��� n�#�!�D�2@�" 1�.(�F	�jQ<,o!�D@%0s���F�O�-z��J�9i!�.P6���JL�"��ƛ�'�!���1Q(�
V��}j��^&'%!򤜰g -���L�.�aƔU!򤏢]��k4�E�8�4`�ʏT�!�Y9tw�MQg�'�(�fJю�!��@F�ʦ�A(]p4�)`ό�j�!��� ��xܬOj�͚�DDC�
OZlt򢟈��X>Ή��"O�Y��
� 갭D�Y�J��*=D�L� _ "N����3y�H4rl-D���O[.�l��FVj.dH��'D���Dǒ5�t���!ԑX�����#D����O�[-��; O;sVƐ(�=D��rnO�-'Ft1P�A'>װ8+2e;D�095�üV�|��#"��v��D�8D��X��@�;�\�؂%��
٬q��7D��ke@�}E~h��
C�=��91 5D�� (�w�A�7qde�a�&I��-P�"O"�#�$��2�p�)�Fۅfۂ�Q�"O�!0i�,���
����SӀL�"O�� "��$1�"�_

�Ñ"O�T�r�/V ha�V�C��!��"O�屠�q�:���J9I��"OJ� ��V (�RI�"!��ᓤ"O�I �^p�(���nx�@"OR�ss$&T*U²e�pn�[�"O�%r�O%2������4ZP�E"Oܵ��J,1bx�e�٥{g8��2"O�*瀖�C �⁋�t\`1$"Ot9� �T��2G�W�x�8��"Otș���sw�8z���03�H-1`"O)��Z<?p���g���?mj�.�y�b�'r��2ӛ��JSG���y2�ƾ)N�����|
�X3R
��yG�a�t}Y��ؐ���BE��yR.�4=�,R�FťiX຤hم�y���6��-��b/�@����;�y��
xp�X(��\!��u�L��y���9�600îC��P�����yԫE(��8��P8��U�$끱�y��}��'/Y:y~h��!T&�y�MWJ�*6Ɨ)$B�2¬��yBAp�J]��F�yH�%I��8�y�HHSpR�.qXB
�.�k�$���Z:M��k��S於qa摍*��Q�ȓ��		�ۧh��Y9�O��ȓ�� 3��O�kEi��lƂ90t��1(~VQ�Uz��u哅�A�D"Of�3��!x�2TY�U�$"OΔ�C�!gy| �c�ΚKT��2�"O*���d�Ǩ�+�(W�YBr�*"O�1�oE�$�d�'׋v�z�y&"OT����'��h�(� �xe��"O�d��Ԇ4ƀ�@�`�� 
&"O�<[�h�	�^�����28^�c6"OZس�A�*�.b���rۈ�[�"Of����n�xm�2�T���8�1"O�X�RB���$$@S�IaP 4"O�x��M߉6<J�0��,sB�@	�"O�M���0I~�5�tgő$�a�"O>��
��-:��]�$&��PB"O@�	"���$`�Aכ%@-�"OR�!��E��2�fd=�X5�d"O���	[	_�R@ա'-���"O�bf�K� ���1iK;e&�$�G"O��񋈵i�L��.S�E9r"O&HP�e\#G��0B��O�H�Kd"O"t��G&|$���C�=6¤)R"O"���j�<|�HH���*!��2""Od$�wN�:m�s�ܸ"*��`"O�hJ����W8�yBW�2]�(��"O�@w�j� �`��=&QpzU"Oh�!R�^%O����@._NX��"OP�*�GӥmF�h����=18	��"On�����iQ~��ʟ��`�C"O����L����ǟ%K��4�P"O���2�R� �X�b��3J�u��"O`;1�P/q,�yqAG1e5n��"O�9�0JPD�X��闙S"�A��"O���0���/��C�46���"O�ԑ��0t�[Щ� � h��"O� ����fا�H�!���Nڂ��"Oi�lL�\�u 5�
��1��"O,\R6��u�tm�uX��)��"O���rG��0����%�r��U�"O���'cΫG؞R��K3 8zU"O|��9:�vM6��$E؜!�"O����E�����S���-��9�"ONY��B[�T�n�q'�� ��"O���kF/t�8� s�6��"O����+��;�I�1;b��"O� Qʍ
Et	S����+RK��yH];*\
t[Z��` EI�aw$C��+9�b�R5�W3p>�H0�Gy �B�	
;�Ќk7#RL�6�c�F�͢C�	(5��R��7�jY���	�]�DC�		�@hQi�X�R����O�C�Ʌt�d0�V��9D�2]s�/�8	ЌB䉇$��0��!{�j\ G 
U��C䉕M���ZP�Z���"�[7zB�� N�4�����;�.�;���7qT@B�	/w��pX���W�FU3��,"�8B��AV���,Ƃ0&JPx���"B�b jY���7n������*�B�0��c�ĩ8	�LB�R�)7�B�	.���Y�$ұ�Ag�Q�|B�I�Z�ڤ1���3>�d���k��B��(V��`��U�@��� 4@U�2��B�	)Rʬ8b���/gA@5��>,�FB�	*@��P��FٚF��R$j�D�B�	0E�����3�ٸ�`بf�TB�	�C�<à-		���sJ�|�HB�	O�dq��(���  l��B�I�l*��`U��U�[d�8B�|B�	������ˏVޚ䪖C��b�^B�I�4�P4����,�D*�扰[bC�ɺ+�ũ�)ٺ�n\�W'C�q��C�	�T�`�i�n�g��x�� �C�(�NA+���.m%!�X$nC�ɆT�v�ؔs2`rC�p���ȓ�t �%� )b�4R�W8mJV����k�mW����bLA�ꬅ�e�l���G
{r4k��ˬ: q�ȓ4d�
A���r�Ȋ�*��8���ȓ!Uj�pA	 �&��*�n
�s� ��ȓD��a)׽Fڰ����VX�&��(�a���^��J��P���Z[����~�-��ʆ"��q���W2�	��Z��qѢ�$H��-�����ȓPSV�����f�hTE��0�����?� ���Ї6���&�?5X؄�)�4�#�&�4X�r�$��p)��?����g
u��=`�'�$j�ȓ'��W"��n�;W��s�rԇȓ*;8]�@�N(iPԍ�T��2��i��-E��9UȚ,M�XI�g�5.�^�ȓ^"`Q�J�!R���L��1D� i�Cن�/�w�Tt��ɊV�<3��5\B���*�3p��|��LJ�<��h�A�|����R�y��zy��'Z����T�kl �{%�IO��'���`�8d��H� �*��y	�'"^̳r�Ʃ4�lE�� ͝#j ���'ʺ!aWk�>��i� �m��'��p"��6��[�/,qf���/O���� ���C��Lp��S�$Ť@��"O���3,B���i6m��v��]��P���Id��a�_+�5��ƙ�v�6��C�<���0>��ơ*�tb%H��~!���p�<ahV�wm�%�T3�Ig��p�<1ӌO[|���䂗Pոiy��h�<٤�
�
Ѳ]��Gזf�"9��E�Ly"�'��`�눜-{"��Q'l\��'#ƀ{4��o֞�ȳ(� 8\�O>��%��;Ӗ�Be�ɶL�4`�Ì��$�˓�0?Q��B&>:��A�<}F�9��v�<Q�I[�D��P4k0b Kq&W�<)�H]����Ɲ��v��J�<i� ^����d�ҧv���BE~y��'j��x�c�|�waH����ϓ�?y�yBDC�?����v�\1w�<��J���y���"�hm�pM��r�r�ٰmɶ�yb	D�~�*ذ�Vj&�� 	#�yi��ҾC��M�v�H�NϽ�y�BK4Nv�h��P�
�l��©��y����m�I�m����!�"B��y�';+FMP5�Z��te���>��=i�y"M�UjTF�&��M㭊�y��
���*Z�L�]�w�R7�yB�M�vw4�;�!��X���i2��y҂��x]zT�Y�V�� ���O��yI�<S��ېGP�YQ�}yD�
�y��f4�3g����p��g�8�y�Aݝ�j��Di�'�lb�$���yr*�&f��J� ��R#���y�CY�/bp�3��׳"� ����=�yB�:0_T�!,�8����J�yB��pCP����µ� ���;�y�#3al��b�d)Q� �y�iW �|Q�"f�;��͂���S�ѹ�V�[��� b	 ^�\����3K��vp����툱�ȓW�R�@�B؉B���*ѵ0�L`��.g���QJ��1��L��͖�J���X�|�`4�H�2��<"t�Q�z�D���0-r,hd�p%4ɡ�O�N��`��[����#�D(�t�,M�	��(�ȓޅ�3*]P3x	n��u"O�X(7'��v[b��$ۮ����D��I�'|,m�0F\+r�� t�ٶH�����"Ov�I�n��AQ�@�K�5j�{B"O��R�6��ɦ�({��m;U"O��{��Z��\���L�HIa�"O����	m�`��'��J�W�P`�<�R���]�Si�.v�b�����\�<��]�|9��x'���W���{p&ch<	C�*FB��*Qn�����8�?��'��y3a�͞e�v1p���>%�R�;�'����J��H�p��5,\��'ØEJ� Q/Wj%�M?!p.�I�'-$���[6#8\"����`��'h�Pc�n��zHp�#�9��y�*OX�=E�ĂӟuI�Mc#O�%�<kė
�y���ġzᎽT|-���ۢ�y�c�9:$DP��	@�)pa1�y�h�#<��lq���!c��iI��L�y�!X�4�8�'��Y$��Z��y2�^'0G@cW�R'%!,��yr��X+E���
�h�����y
� 
e��H�2w����X"x��`B�"O�B��1OAC%O$<��U&"O���[>m"0�qa�::�&��"O���S�W����-��"O�A�d�<��M�R��R���2�"O"���^�
�����ss
mۆ"ObDHWc�M�8H!�2m,�����d>m�'��	��@�iG�b�����J9D���aK�a��r�cB�;�Dx2�*D��sΈ��[o��Y�� �
,D�t�QJ�_��L��Vn�,��+D�t;�- ZD����?{I���5K)D�����>�sQ	V�"�̋&E2D�� ��C�/�
Qc��3`��0�;�I_���S%�� j9@:tyge�:$H�C�InGH �!k�f��(���Y�k�r�O�<LO���*�Nz<c��/[��t��"O��q�ی\�:���M�#�2��S"O`��4��G~�(�M�B���"Ohd��N\�T߬��ҎF?|�؈#P"O4����Ѿ}��%餬��O�� ��"OZ,x�ʕo�Ό8ŋ�3"l�y��'��n �X`��҈_���V����'�a|b])��s1 E�Z��M� ̓�y��ʂ"�����I�K�<,�!ҷ�y�ÔL6�І"�H��§�yO�0H \;�J��oBH�t�2�y��|�| ��@6p���j�D�y�h
G�P\��� V<��z�gH���x�/�n�꽓�	@.d|�Dɷ�Y�to�Ip��`�K�!z&�#'nC$�\;a�5D�� 0��*e�4ĨQɟ�IV�8d�&D�Ȃ��ō?���7���%�@a�`(?D���!�ج5�����F�*�+�=!�Dɤ�D���dx���@$^!�$Z�d��C�
A�u���u}!���y���;�ԃRDa3u,[�a�!�$�.�bX
��$�K9J�`}��' ���0n��&�6Qr�ǌv�t���'|I�@���X�qe��V�.�'�8��B�I�B�b5ʗ�%��Y�'��P ��R*5��Uؔ������ߓ�?��O�b�#Ք5� �)窆,u!Z�B"O��1DF0���/R4CmpA�"O`9��ᓠs#����D�6]jt"O��u&ڮe���G���i� "Od�A���<�գ'� }rޔ�C"Opk@��-3���!v%W�OY�I�c"Oޔ2Ŭ�o��|å�I2;���T�'$1O�9�o6�f������e�1"O��#�!1u4�@���\��=��"Ol�r��Αe6��F���P̊�"OL�-�.<b�xx@/ʬV��I�W"OމR&K�3����P�K&�� jW"O��(�ԕ����b\	y`$�AO�T���0t�}���F��$i�� :D�(p����-QW���Z��t��7D�䒱�� t���'FD.K!z 2�"D�\i'�
zG�q�(mc�A�  D�@jC� �S�*����!F���1�M*D� ���ҔF�(�iFA��B �wm)D���㨜5s5��8&)W�;�2L�Gg#D�� �H� byz-chէ6״����>D�pc�N�d������{蚈�>D�� b���G��ZB氂���9U��%��"O�x �w�p0��6��	R"OL���/�]�z�k��LX�y"O�4si�s����a22���c"O���1GQ"�h�9��Y@P�90"OB1���Y+0$b��:�I��"Of��A�M����΃TvT"O$P24� �L�|;e��N�Da5"OP8�d���fi��O�|�p��"OBɹ��Xha�t��5�zT�a"Ox���qpdM{�m��V����""O�8����#U��P�:2Ƞ�a"O\�(tKa����(�"��q"O���h��K�\c�-N%<���	"OLIt�<cr<�;�I��J&p�ʑ"O,�1��7kA�c�N��Y�"O�D�Ů�r16}H��LD< �a"O��!wO��;��9[F��N:t���"O�,P�Z�<�£�ݞb &=��"O�P���>6�h�k�o���!Zr"OsPH�q*4k��K8�|�DR����{�"�9ᜀ,��J���'*B�IvO��JS�Z)hb����C3��C�	:��L�D��^�IȂn�Co�C�ɐ�(��A�2��钔��0�B�I(��#n_�hw^]�%FP�CΰB�	�6�8�7L�2�4x�͛�A��B㉀��A�°M3�:v�Q8S��'�џ�<�	�9�IBC�n{$K+d�<p�9`���ۄi�1�v+�`�U�<�&"�6fHH�$�8ʸT떃[X�<� c@�V���'
:XG����V�<�Ѐ��$�A
ҋC�V ���m|�<q��/ӨQiSCp�T��pl74�p��`K�[,��BE\2r6�� ��X��b�'P�L�b=b�j�;�hP�,5��i�
��ta��3���F�3fi���b�ʹ��	�^�V�("-�N���ȓ:��=M�>~qq��r|�y�ȓ����VJZ�!<�I��ώ��\�ȓ��}""D���(�!!@��p�ȓ:�V�2�
��ci�E��܈�\�ȓl���&*�t��S*C�ǒ݅�S#عk��Z	u�,�z�� +�P؅�mܨ9����<��"B�t����C�h�����,�Zے Μ0jI�ȓo�@�S���#k��,�q&VC����ȓ�hy���)�%�1'��>����0����&�۾'v�Z�g�&�|���u��h��ĕ;.�"�J�N7C�蔠�d�'N��I[��H��O��Z���kƜ�r�"x��6D�0��'O��	�uj�;S�Zi2.1D�tc#���1���b��Z�<�F�(�0D����&L3J/����AD
|2m)$/D��b蔃v���I������k+D����șP����� �`��Y�p-/��0<y#��#r�)��k�M�б3w�I�<1G�G;�>�ç��c��1�#��A�<���ej,T��KݏJ�E`b�~�<�5��<+s��`��H'tNZ�#S��`�<q2%��\z�
�jȹG����"��Y�<�n�>[�Hi��aH�f����W�<�'@�i�2̃`� +(�L�ua�T�<q]ڈ���M"�k�OƎՌB�)� �����
mt�a�aG	f,fH�7"O$��6� k�� Wm	�(��e"O��bti�v˾D�R�O~��lSB"Oĸ0�X�2�`l�Q�,��9��"OZL����0��<0 ����� 7"O�����A�#�b�s!
�F���Aq"O���̞;`9����� ��8C��-LO��,7O�H��cM1_R�K�"O���+L,<��(��ǫo ��P"O�lI�!�;���A#I Tk�H�%"O�YI�e�8]�B@�v`L+j���"O"��Ī��y�Ibsb�0W�eR"OL�i�\�p5� 7UcB9�@�'!�$��Xy�צ"pW����'!�DͲv���9P��[>x]�	��J!�d^��,�%��,p�՛p�],!�ɽ3����ŢAq��Z��2�!���9�P$ta�2R�U3�P�E�!��0�H���ӌ6̠̒T��:W�!�$PZJQ��-�,4�P��%ّ/��}���,�3�	�JT�"��(�t�3D�@�Tm5W��u�`��}.�dI��3D�(�W���F���sgK�?@*�ۑ�<D�,��iF�A��1.MˣI;�O>˓@�f�k��BVi�5+�i��J/$�#�'�x�!�̥,�x��c�S3 	�'Iv�c2�ý>�va�C�S�xl$� �'��5��%2!.��Ӎ�sgT���'���:�L�{�8���˟�R�Y�'��P�b�>�p噳X�]m>H�
�'�\� �N�	���u"WZ��8���?ye�r� �L	}�<)E�ǵ\��L��'�ԈW��1|
�tI����Sn�<{�Ƙ'�PCAI:o�T�L�W�(�'�p���*�LiA6σ�W���;�'O(𘗏�q0����8��E�'5���c�m���� D�)W����'ɰ��g��m� yp���*��
�'|��	�G+���'��	*���	�'�k�$����r Ə/l<��"O6e���Ėx�5��rQFds�"O� 3�c�N�J��[HOj��'"O�����S�y���T9b6Ĭ)�"OmK��Y�f=~�J�i�:xm�p"Of$:2��27a6����½=(t�H�"O��S��= �fi��%�;`1QU��,�S�i:t��A$h�R`��@c07�!�$A��0�dI�	`��oF!W,B�ɢW�H5 ԌB-2	�$���ߛ �C�I�"�Ha�N-p &�J6��
h�pC�	 >�f㕵���iA-HY_�C�I���јėu@��E�]�C��+�*U(A�E���;q�:GO&�O,˓�0|�wD�A[�w�,�N��bC�<�wOݟKTؑq�/L�a-�#֦�{�<q��ND�� �=x�d�sK�9�!�	t�b���#NO$�q�,��s�!��&xf�,(��q�&X2Dk���!�߆ء@uGQ�1�xUb隅y�!�$�:5����.��9���X��@�l!�dŏ0�QCED��A����F�/U!�d<q��p�A@�uWz%#��ST]!��ڃ����cE��h��T�9�!��M�tA��7��,X@����g�?]�!�� ��S.D�8n�e�g����!d"O�ym�1��ӅᚑR�T��"O��B�V2T����AL�x�8�"O��У_����:�B�=CQ$囒"Od���nZM��Q�r�̷�%k$�	m�O�x�7¹R�&���І	�>��'���pq��/[�r� 5��JE@��
�'����w�J�4ʖ+�nĎC����	�'�� 㰎�l���C�A܂A����	���' �)�m�'6�\���9H����'A��R@V<�b��@E;9V�)I�'Ȩ|�D*_�c��@���2-n�C�'G2�1!���@�tؙ�O�2ٜ4�
�'\`�2�C.BD �;����*&~p�
�'�d����@�J�7埲��[�'k��V/Ȫj���hvK��D���'�j��v�C������ڄ�H+�'��fC��%�hda�H�:F(i�'�����GĂEI�G�	�0$)�'�����Lʍx�2\��ҽte�0+�'��y	�.�*�M���aDʠ��'qL���춀�+�j��\�Ƅ �'J����-�$#�nh�aF��Q28�!�'Ҙ�@ �" ���	�Nݪ1��'��3��R1xlz���t\ݘ��d?���:S�M�)�Z��g`IuN]�F"O48�C�V)a*A�6f�3k>@X��"O��1�N6c�I�OSa'���"O���"o۩U~�����V�%"Oހ@d22"�j& N&4�m��"OXAٶ�
�?1��:��	��bq"O@=P��FJ%ЖA�j���	�"O��HƎ1p�j�8�o3y���;�"O����C� �n����S����"O*�X�,ƁL`v@�C<[4�c�"O@��6Ƃ�i=�B�!K6,"Υ3"O|1��Y�u���)3'A�FE�$�'��ɱ{6����P�d � Z'��k�0B䉱^#*�q��M:$�X��Y/2��B�ɚ9��PX��2���[� �B䉂&�H����w���B
HC�I0�lqA6A�e?��A5hW(C�	5@P�L�&G�mw��d� 
��B�ɟdt �Kv ��&d���oZ�p����8?� .�8!8�I�gP4_rB<+�mFM�<Y���+ �XA,Ąd��-sŏ�I�<A� 'ix�k���y�6M�bA�E�<�)Ɩd�Fe�1�<	�89��Fy�<�(��p)V�`�66��dq��Lr�<���Vw%����H�X�����k�<����8e��! �}��Ҥ-j�<q�Y2�@PIZ3"8��JP�<����[�6S���2c�4*R%HH�<q��e�D\���-$����$*UC�<	Q�V]�9˗/G5	h<�N�d�<���r����`�z�Q�q��^�<����u�Ы�DEL^��Cc[�<�����<|�Ah��m���T�<9�|0�z� �g�ֹ@F�O�<JO�.��b�d��	e�<�Ǉӿy�C�C�V�,�+�� d�<q�֝kb����
F���i��	�^�<	�o�8~>ݳf�Ǩ'�e�b�q�<���D�5a��"C`��w�J܁0��m�<� =��BM*�`;�k��3Yr��"O.ݙG�
��@��*�FX��q]�З'0ў�O.@��@KI�c�5j
J))v@�x�'ǎLcS�@&x�1:VJ�����'����X��蜒bNP$���'��� ��S�|��J�L̜l0�Q���x��D�&p��Al@+oo�`j���yr�üq֎-�1 Ϙ`:|��iP�y���t���(ƻb��y��O��yr�-:���:&#��A����X�yߌXI���A"آM�0���&��y2&ٜEު��Ԫ�Jnf!��k ���'~ў�O��t	@�Y( �N��-0Z����'��p�͈(,�|A��ڹV�A�'-����s�E
����k��Qc�'�?��j]<V��q+��@,<K�x��$D�4ze��=~�� ,m��kы-D��Ök�
� \0��\([@��7�,D���Ѓ6]�v�����{=V��a*(D�@�C��Yw`%;D�D 3� ��&�9D���FӢer���0Pi�a�;D�|�&�z�A�!���\A�"�$<O�#<�P�ȹ�n�K$�ЛR���y���G�<	��Rh���N�u\�7�h�<�V@>:� �'��h�V�R�l�<Ɂ�L�1����^ k���R�<�DôM��x��X�G�p��EO�<	$/�3T�h����bA:�D�t�<!!�I�4/�9I��]�4�Z�g�Jf�<Y7��]���3���fIԁ���ܖ'~ў�>]80#�B�Z��Ũ9X9�D��1D����z�0�ԀCE:j|P��,D�xbp)^.C���ns���J+D�@���O�6![�a�@��@��(D�d1����UzT��I 
����&'D�|�wkZ"jlPr#&CC�ZU#ҁ&���/§C�x��A7AL$a�	�bT������	�6\¬(׵?�\�2�K(>B�	�O���M�3.�6��`	J�B�,}؊	pC�4�l�Y�Q�g�B䉓%���q��|�ub�-ʇɲB�I� 2����6�J�`r�&�TB��&u�ؙ�3g�W��dQ��I�a����$8�w/�C�k�2�r�H%gr��E{��'���97���X��R��4D��=y
�'��<QOP=SI�]HPC˅_h�9�'�N�)�&~g��� ��0�l��
�'��u��ɜW�y���*U�l�
�'�<���#������Y+�e�	�'���au�8%�Dj �T�](
���'%~��&�):�>p�'��7� PQ	�']J0�0m�z�ĩ��P�!�\��'(���I�d<�F����,���'�2PSqjD�J�,�P�&'	�x!�'G�Mhq�O�X��8��EV�y�p0�'�&��IE�W��$�ta	2[tm9�'X��W��b3�D!�
TI��Q�
�'B�Y3���st*�!����r2��z	�'l�aKr,�5t����qa�W�pA��'�`��.��`��蓯,�8E��'x�l�d����RQ`c����X���'�ڈ�����p�"�*���'���c'"6}&x��.lx���'\�<��ؚu������L3������ E�C#In�<pg��IM�h���|��)�x5��5�<o��A�ʔ<�XB�ɺKfp����F﬽� bHJZ�C�ɻ2,�H�f�ܷg�vY�w�ǆh�C�ɓ��\K ĚdXv�i�K��C��T��a�[i!����/S��]�	�'��y��n,Q� �1����'O�فoP�X"\Đ"�-{��p�
�'B�)Y��F:e�v�P�F�l�� �'qv�;�h���*��Mg�'�O�%c��J��ѭМ���1�f��U��q�Ɛd�(e������k{�X��"�ܹ���	<���>T-�u�X	U;L�ʄ$x8�m�ȓU�Ry��!��QY��$>+�`�	˟��?E���7�F
�� ȷDY�w�ڥ��"OB�Z�o�!S�	�C[��4�'�ў"~�gd9h0�yj���:�x���y���E:�!L�s'(d#$͗�y�"�>ֶ�"!d�#��e��o��y�E�'-� �J����k
S��Py�����^�qv�Є���s� Bb�'��'t���Hr�BX�ҁ��� T|┐cK�wh<����� ��D�iGpc3��?i����O.牌,��"Q���s�ˉu��C�I�=��!$��#!� 0�d�$g�fC�I0Z���A0�L��Ɗ��HC�I�PެP���9)r���E�*G�LB䉽9�ЈZw�3�@���[9zv�C㉂�ة�RCL�K��]�5��Næ���n�Ey�fG�1��#�r!����'B��C7b�7�Y0��š#<hL`�'�H��/îZ��mkaHڡH�'���S+P4B�������ƕp�' pI�!g�n�bB��'�}��'�h�H�N��L)ңG	Y^,����y"΂�O^rH9BJI0&e��
�'R�˧H��)P��e�?�l����'�P�#�s<��3�{�D�s	�'j��`"&Nn��S�C?�j�'u.p#���~ Hd�+f��S�'�b�j$o�T
�öˍ+���
�'+����O�v9�!�$�L�
�'�|�j&UL��K�k�Ji��'l�K�B�>ʁ`���*�q�'�bh�d;�zԺ���7[�����'�� ���J�.D�pg��R��u �'�Ea�ٝ�x\S�N�Qӌ��'"p]��-s[���+מr���'�u���K}�Mq�b��
�����'¥I��V� }>��,�r�,�����'h`�YD�фD���s�
��3�N`��'�$�w
^oA
�Y��S,�ذ��'�������>q���f_��X�'�p�ǨA�}r�53��T��S�'��|{�Z7r��Tj�� Y3n5��'jh���W	!�^�[3��O3����'�4�SCʮ4P�A�g�үC>6HP	���ć�K5�q�7�T$K��qP&�g}!�&���&�� >���1&M��!�$�����"6AǞo% l[�))�!��2S���R�h�P��)�&Y�a!�d
7�$F�ϘU`*�y"�PFP!�$�0C�V�@T/_��4�vjХmc!�� ���Soq۴���t��l�Q"O��×��2����ȺY�8��"O:uS��W }�vi�� M��E"OD��.ǧ.��<���Ֆw��#@"OD�h�J�b�B%i��]�q�"&"O=�.Z�.I����9Ϡ�Z%"O�A���ƕ2���D�8�j͘�"O�us�%>�X{���b��Ȣ��'1O�I G�9*�@��	�"O<�#T M�F|~�Qe�C���"OLh�b�ׯ-|���%*�Da��"O$��T�	�!�h�AӒH�6u��"O�Y��ၛ<���xѠ!0����2"OLX��#� <���ɇ=+|&��"O��*0	��s��y�����QE���q�'�I5K�\����	6KanA��#3>jB�I�!�T����)�0�9'��GDB�	�%�\���R�%Z�刷.֮��C�I:����D=wM �7o��C�ɨF0�PTi�(J�P�eFTAw6B����sc�َm4�(�V��"B�ɲr�,�*!�Q�kXE��Ɏ�p����d�O��	&�(
 c�)B�"�S�΍�#��˓��<!�Ob�� %�=������/* �5 �"O ���K��d���@'�?�`X��"O�ՑDAO�a/,1uc[�C*��"O�x�A��)qg�4!'�I �����"O����IN���r�ڥ5T]��"O��ѩ������G��Ҁ"a�'�$Wj��"Bg�+f��Q _�qZ��'}a~�ꔱa\J�hc��92�0H�����<�O:�Q��K����E_k��T"OQ�C�_C��Vƕj^E{�"O ��`A�4{��ChD�	UhPg"O����m�2�~��'R;RȀ�"OJ0��X1J�8 VA�N=���U��H�O�}�%R� ��aC�;@���'��'�J�H����@j� ���^f� ���?Q�vB!���6I�!��i�Mg$��|͔$*�*M_L��Ytc�t��ȓH)h�KH��C��%��/@"la��H�lm���S |���H
� �Ɠ�@̓���:G��Pj�BJ?�İ����O�#|�`T 0�r�^�:&�4$��������p~���n舷b�1�\����� �?Y�'�pH�wJF�c2 
�Ճe�L�
�'q�H#��+t]rT��nU�Xi�'�QQG��s�tи!��|(
�'��#��Ͼ,j�[��X>4	�	�'u�<���ãM��T��F�<sx�S���O�˓��DG1,JQz��3i˾��5O˨f5^B�<a8�!�ŘX���*�!��B�0>���ʄ�ӻ ��=C�Ǆ�&C�!��q�����FقA����5K��C�I��:��J1Ti��mF�D���-\āf*�$�<��؍��}���G�^��PA�!���XS�{�<SL!	P���F-��O
oF!�D QC��EE�1��}r�/�K/!��Em,� ��<M"z@�!�G!��/��p!i���q�l��?;!�%�ܭ����&	�"�L�.r+!��F+t^��tAֈM0�����&�{�D�4; ^��bn�
*��eBğ8b!�� ����Mƪt?��J�܇D������'���X� �����P��Q1Q	$>�!����};Ɓ88�" 2��A'>�!�$�0��J��Bm8�s�C��!򄟗7�ZP	6n�.[N��2iA9[�!�D���g��N8�l!�(�2!�!�d�@�v+E�6.�`5�G�=�!�� k�4�"#��l�:CEԞ`�!����P��Ȅ�h�9	�m�}}!�d��c���i�_r��aR�!��D��4�h��+8��(%g�!��V�d�P����v%�zҦ�$�!�$�4b,�EM�[<�����R�!��������*3�b�z��ߤ|�!���/��1p ���6��ɘ2d��:�!���I�B�ى&��Iq�V�!�Đ=o��\��Iřh%s7)Z�r�!򄔧RAR��&���JX��iJ�3�!�0f�2����Kg�P:&�Ȏ5�!�D���2�*��\�.�@X�eٮ!� �?�)i�nF�x���+7�
T�!��NJ�C���N���ӵ���;�!�$\�Q�����1�b�
z�!򄙍T��Q�B��/s�VI��`��!�J�NR�q�ѤS�c}Π��M5s!�dZ���� ��%}��D]2k_!�D�8wp ht^m��%E8ci!��x�4Prf���T 5{��F"c!�D�u5��pc�=8�	���(!��
�<�braР	�IP��"OP�K�m�5��](Q��6#t�9�"O|����6l���.�:���0"O�@�瀷d;�q����d��R�"O��3��9�\��%�37����"O�Y��t��=�bDG�B� ��A"O�ih�`�?�� �#�Q#Dؘ=�"O~bdڌs�*A�%�8E� �Y�"OJ��LO�^�ҌY�� �#���� "O��O�@�>0&����E�g�<��C܆;.tS*O�NQ��h�Fb�<��&��?�0T��-^��l�T�Qa�<�!ܢ���8��2([�<9$�N�h��-�VI"�"�Q�<	f$�%�zu�W�%
��.�c�<ieJ�o|�K��
A�\� g�c�<�3�D>t �E�0-[�V�t��!HW�<)Ra��7���DJRM)���P�<����|B7	�/R�Aц��u�<�rɁ�*z��af�ެPd��X�<�! ���½A���L�r	J��U�<����_O��S4���I�t́f�TT�<Y0	JPcp�ue��ϲ����e�<!㊚�2�.�P��B�\>��͔Y�<�f���"ʮ�;$@Qs��	',U�<�N]2\�����B�?hp-y�N�<٦c�2ܴ��t"K����R�F�<�&�@3tz
��󢖕sEp��p�~�<Y���5����[���P�6�\��ȓH"@�ԌU�&�Zth$�P�t_X,�ȓm�V ��Z V�l��A�
[�p��"/^�#э�8�(�5���MɘM��b�V�����U�E�;:�ڰ�ȓ,��1�aBQKҰ ;𧝶CV����}r�����>�$���}�⡇�S�? ڝ�R�J�sS�$��*N=+��`"Ol����+D��+Ӛ�\Y�"O܁yI��Y䴈q7e�3f��� "O����Q mx�Xq�#ݍ�B�S"O��� ͌�����j��-C"O���g�X��H� Ę|�bT�"O@ͳe �l��p��N	so��0�"O�i�4�مL�Zu ܽ 54I�4"O�� a�j�� A`�ճoޜ�R"O�e+�cձh�\�D�څx0$26"Oh���O���34f֧�(�K$"O�8!�F?0(P@U%8`�p���"O��1�Β�8%0��Չ%۸��"O�2��J��xH4��:u�"OȅA����<:�(�0^�*��""O&�a���e� �(@@E��"Oe�V�q "���S0#�6��"Ot}��lቝ�&o���V"Oލ��mY�O�$��vI:u�f��V"O�
T�D�RMY�H��g
�H�b"O�\	jܥL�!ز[��RX�b"ON�%!a�~�X�J�za#�"O@D"�R2OO�50�������"O(�����1�j]�ť�I��	��"O��"/�7X/&�:���+X�N�*7"O�V�؊��s�L�>�0BC"O��[S� 9��AM]���A�R"O"$�1��I��M����)�ֵ�P"O`��Bϊ���!�C�y�0X�A"O�Lq�3u^�) *�<�\ �"O@��(��dr�Ȱ�b29h���s"O8�规Y#P�ЁO��8"O�L�%'�$u�Aڳmڞ({�"O%�Ff�]���z� ȿ:��Y��"Ob��hV8��ysΙ�����"O�9���`�`�;���G"O���Wcܳ&&� �1���Q�F"OLp����z%hUeD�3s"O�qS*��h�,��b��xGV��"O�i��×,d���x�[+?b|�F"O�m�BN4:UY�	;%��"O�|�p���r]b(����^�r���"OD��L��6��P�tL5y՘A�!"O���g��T�Ѝ� *T�#�|Xx�"O�5�#�ij�Yቔ�o�N4ڄ"O - 5)_%Z�:�Ш�0$��`H�"O�QFnT6,B>�AA�t13f"O�M��h�:��E+3a�$i����6"OH�XЎȯ{�p�	"�ҷ1Y�}��'�6��d�ƑA�r93�b]�LH��X�'��A�։^&^E ��sJ��H��9�	�'��@�2�)��D���A��-�	�'����aDL҄�.;����'�����-��Q��	#jR�c�'�<m̒s��|!@�
�Ni�}"�'Ě��e��Lڼ����T��4��'��]�������R�>�f���'~P��@kؕO^j�Q�H >d�q:	�'!&��N�5��� S7?.=K�'��9��2��EAB� 0����'S�<��W?E���1��T>0�')i!蓡d�.Ա�
F�D]�	�'���$߰NQ���b'OE�!K�'��u��l���pP+���:Q0MP��� �H(B�^����'Ꮃa�h��"O��Se
A]0��� T
���"O�A�I�69m���O�"�2��s"O���i��g�Y���'�]Q4"O��� KD4F��2�,��	�$��"O�ɂB\�CX�9F�P�z�n�"O�i3�Vm�YR*���<" "O����n�,+2�PA��6l�����"O>��W�	A�@́�a١-C��sA"O����͈#"�X�A�/�2PC�q+ "O6	�P���8�s�H�/6L��%"O�I�R���L鹐^%7@J��"O[k��,O�2�R6>7�c"Oz5�3Ȟ�=�p&��Z/��S"O�z��"CV\�B���$Z���"O�a�C����0bh���)D"O�����b���{��1J�>��"O�Cq�܃�J�#al�"Q�i�"O���,_ �*���I����"O�-�ǊV8#ˤ���N��KB"Oؐ�S�Ŵ4����N�,���"OPX���g'iʴ�O�!&���"O�!��Iz���K_	�E#7"OL����
��Hb�A��t.�:r"O �!Q�8��ɱ�%SgZL�"O<�IX�|�bp/̎<Y:��E"O���f�>t
9���	7#�Uц"O|�B&N �}�����Ta�"O�C�
i��"�5`�Q�&"O�)Z���1٪���K;Y�B%"O�����\�H�L��FEB@����"OR(2nI�j�"���A�;M.y��"OZh����2�t��C�I���	�"O�y5��!x�iB'�9�:�"O�˥���%E�A��&m���%"Oh4�
�b�J�U�%���i�R~B*��<ɍy��������Ɓ?�n���NN[a!��ъKu0A�_�R�S�� /+�5��R��cAH@it���l�
�� c4�4$�,���&�R�Buh�.<��)���5��Y�'��	�%�1��|�S��@�`9*	�:���䎁X(��ul�
n��)���("�!�d���\��cג|U��`��1�� ����?��O^"t¼�Z��(i��d�;D���p�Gyy��2��բP����&,$��{؞(�3�]�Sl}�w��mTȻ��6�Ov�ͺ��L�&ڜw�_�FP�ȓc�:!�'���t����aA,h�TG{��O��I�LS�!l:�A	5L5�%��'@�D3Vn̥ �ZDk�C��2K�e���'q���S�0���N�*.��{�'}�tXr.��g�$��͍��D-��y�Z�,E��'�A�PH�&Q*gJ�0�!��'�B�1p��CU�!���Z\~ ��'ߐ���m ��q���֕G%|��
�'�L� �T���aE �B)0a�
�'�h$"��=��M�O��=�. �	�'�>T��H��zAj�A���l^���'yDa�qb�O�
�y�I)rT��'.Y�Н2��0��P_ ]�'�ܘy�nן@����`�
�n���'���R�#NP�Z�8��7Fк�'�FIv�/��Lꣃ�H+<D��'6�H�뒑�$q:��3M�<`��� l@¦�]�y~x8P&F,�8��f"O�"G���;�M�1pq�(��"Ov��t��Ԙ��M�*Z�q��"O(�8qlP+I|-B�Rx�kU"OH���!ڽ}�=�@���%P�}I�"OD�à�N�:a� I��x���a"O�L�lQ#9t�g"��,Y�"O.�`'��u�а�A�f�ܨ��"O\��`o΅&���r(Լ9�@�KC"O�a�Ӂ\3R�NȢUh��K��]�$"O(3�+Ei����2-��@D��(O?�Ɏ~bj��+2l�����?C䉠7���2wI�w��)Qf�&m��B�ɉ��5[�m��@%
�`��B�		h�H����/K-ԀA��ȕQ�&B�I�X�B�
�� ��g�iYR�<ٍ�T>co[�>RT��*�e#8���m8D��@��^��b�䘸kM��1e"D�D
��W�B��4#Z9ִ\c�@>D�iŧF�@�P�3�-𰼈��>D�|�0��82� ���"��%�rh1�OBʓj:�)rKĩ6�P"@�18fX1�ȓI�@C��V?@�mF눴N�� ���������Qo(�����L�ࠄȓHX&�I3�V�t9�$SU	X�H1�ȓ1�v���FU�f�t����1B,��ɨF��:|�����dڝx:�]ے�5Tu�B�I�?�l5����E�|�@� Τ+��<q��T>�XfO�,c�`�&b^=�4���'D��#4�;BLd}#��֢ ��p�pFF:�(Of�}�� �*�z��T�r� b�^$�xD}b���֜�����/Rt�p딋�E�Ksa~GJ�d�l�eY41���#Ŋʵ���=��|�0�|��$���(���/����ڙ�yb@+Y�1�#�ٖ1�~K�n���~B5O�b��' �h�9D���ipTQ�E��~��ȓx�$i�X�P��ÇݳA�>-��L���h����f���A��Š:�JA�˞G�ay����.h�ޑ1�����Jm�#�^ C���yO<yq��>E��'���4ȇ�l�Jx���C�.��!��'L��Be�h^���IX\$�����'nay"i΃4tmiM��m��U�1��
�ē�HO��D�|�����9�T�i�V��ce��yb�Z)$�����ϛWE�8p3������y��d3���/��:6�)�J��t@�NZ B䉣.jm ��/�TŃ�ͳ\nC�ɇ"�~�Y�^�� cq����2��������ҟD�#(��7ՌE ��/v4@U�d�,�>�O����da��c  �u���ە�I�1�O����9dH�����$|�q�G�V�<�JB�I�qN ��w�P�9��RDB�V}f6�%�Id?�O-��MS#�XA��`���)�T�"�C�<@FE	�F�ђ�Ш/�r��vD�<�������b��b���Q����P��#J�!��"O�,c�LޙMʘ#,߸E8�q��$1|O�J��+��ZVJ�0�l �8O������Q��$"���1A�Pka���zRnL_̓kn.`���
a��=��XM�Zą�iܓdX�Q$��hj�li�-g��>	L��F���S�&T�qcN�x���1��y��Ô9��@b�m�p�e�R������6�S�O��iɀ��O���)g�q��Ě�'"�%z�DE5^[FY��ɩ_�m�'�t��$�$.QH�[��H��`Y��� �Q3 ��wIX�a�p����"Ol�eL �BL"A��@��HȶOL��T(kt��d�� ����aM��J�#�'21O�32C��7É=d �F��t2���]��~��)ŗ�h���`�t�e �R���p?)�%ҢX��	�/��\�~@�f �Z?Ip�H���'<��|�g$�/���O�.s�����5�O���OP�A��L����d�q�.�S��y��Q��м�cdea�%@��+�(O�9�c#2�}S���Fm�.b��ۣ��}��t�ȓ([�=� �ɍ;D��A�D��4���E��k҃^R��]�4��(�(0�ȓ{�hE��&��?�ʵr f\~6P�>y������ة�*|h�/�X��)+�C���y��ݨu��1ԀۜS_��q(��HO���Іr��@��Ϝ+N�����M�A|!�IP��[�I.}B��0ˉ}!�+B���M�!0I�TgSQ�XG{*��1;7l!.f��Qw�طޞ�h5�4�D3�O�P:���*d~�rn_�(t-��L~��H���I�zh��	¡�`4�vc�HB�I�u$Y`��N)I�<��$��<Ki|� �'�ўH*�5jt}�UA�=}�����P�<!�,���5��@�0����P}�|ri(�g}�-D�2\��g*"����3��,�y�`T(a`8����ݹ�Zi��D ���mX��2擩}��%@r�W�Z^�xk�#>D����_��a�0�V\�X�o1D��r"�)*��	���F�,T.ES�c5D�(��U�N��A�n�<7  %!�	5D�Ĩ뙏 U���9p`�9�D5D����ļi<](c���R\JC1���	�0daC�.XLU�$A�\�$���� 1�s���7����$Z$���IZ��(FH�8Bǟ�U|��fD�J�\��JQ�gD�f��䅁�f�)�ȓN�ș�� H�PB,c�b(Q ���M�&|3P��(U�|M(t�F�O���ȓ|�xYBA��jS�'/��?�	�� ��]��!J1g��;`�����P��x$�����7p�X� ��v�4�ȓD�����Ҹ��5#^�PE����o�e(�dM�.�l��%��!@����ȓ&E4�ć��B9j @�	�ȓs��$�ׁ�.���Ig��I~��0f(��7OLîUS�a��8��ȓZ<��ɖ6/��B���^�|ɇ�O��6�#!/Ρ�$�X#z�N�ȓU�����K�@��PV��5�ȓt�D�hGN�,������
y����pNI[��P
����C	���ȓ@�f�����L���Bڰ�ȓcC�X(T�
Z��pTh�8�.��ȓ	��`������=)�9�"y��z.ݸD
����@���A���	=���ĩF�O�2����<&6�ȓs�*��Λ;NJ���� BF���ȓT����$��O���f�S�W��ȇ�1;\	ZR .�$����+r���ȓ/�j�j�グ8� ��U��~��$��0�tl���-� h��I��xd��!{:�	6-�C�\0��I��C�L�ȓR$@�U��%m�fl��'�A@8���r�ز�ʆ}��Y��A7!����S�? j CT9L=����|c�h�1"O��Pg㉡@�wH�&=Z�H(D�x�Ӆ�)$�$qp�Ϯ�#��;D�(Ĥ� �A0��Zq<�A��6D��z�-�4D(U�qǜF��h�Q/D����k�>9��`wM^=QS���@�,找V\�����)o���`�؉q��c�@`�L��.�'���'��Q�b(D�l����Ld�i3ÚI!�*�$D�t�0�זU�Ƹ)ËL���1�g#D��j��4���T��3A�-��� D����`�+Q�$�qٮv��uG?D�,�sdW~ ��v�ٕe���S;D�\re��+pޠ�q'�!y��5a�;D�,���͈9�r]�dg*.r��6�/D���D ���-�����v�"�'+D�\���a~aSVA�#f^Zٻ�a/D�t�te�=F{|��`D�[���"/D��iw�	�tq��>P�Q�J/D��`���'rn.��$�ā\��(7D�����m���M���B'L7D���t�J<,���%^��ԋ�D>D����a��hߞ�yu�9n�2��+D�D����	�>�Y�g-�taE�)D�L�'��G�s�EZC��l��#%D�l�w��=F�d��f[�lڢx(B$D����,¥����&(��{3Z�˶�.D�d�q���z��DJf�Ȩ�:i��(-D� �G��@�����Ia>-ӵM*D���Q�Q��`}��j[�R%�H{��>D����~����غ��lÒ�#D�H��
��S�н���> �j����#D����aM$�F��L��
�id�#D���f�\�
�D<��ˉ|=8<0�i+D����g]�_�f��2"yd�vo&D��+ �,c^Xu�#�͘>&�Г�2�ɟ�X��?%?e�w)H�H��$O�0T�R�0D��if�ΕmD`ɢfM->0�:���d�qOl	B%�3?��B��ҝ�Ӂ�R]��[焚T�<�"�W�l�\aI��I%Sƚ Z���+l9���5�O���ug��+ƪ�V��15��D��'�qSs�[�D��/h�Lxv���uΠV�Ռ=�!�$�$_�Z��%��b�eCQ)�)`�1O�y�i �ḧ�O~ ��C�'t}�Y�ud͏F��B
�'|��GC**1 N�6��]��a�zܓK�QD��O ����4<&eO�4J��9W"O��N�*�)�d��?x��.
�b��I Kfd08�A�F�X���KF�����.rh�.�eP���2��$@�c�%�!�ȓ�<MxG��V��]�Ңϊ � �Dx2�ځ:�qF�Ώ/]�%! +�=O��� �)�y©�	�j`*�C>9 �0�W�
�4p�pI�f�S��y���X�Q���:z��ɔ����y�����SƧۗ�t%�ㄞ��y���bw�m���-u�|���*� �b�Y�����^�.�`�'�2��oV�2|��5�w��}q�'Y�Y1p�˼d��p�!EH5dh �H��DM�μl����ʨ#���z�J�-$��UA��!�$�?1rb�� Ί�O��J�.�<5���cG�J�S��?�� /��h+$������Fl�w�<1�@�QqBtʢ�޾[��(c��K�<�dm�kw���Kڿ\x�:�g�B�<�De�<��A1F�H;1J@͢��Gx�<QG�� NrK��f� d��|�<�V∋q��P5K�48��	�x�<� �X{g�ԱB�M�`)��<Ȣ�s"O��7���BLl�r�W�=�����"O��ɢM�+4�2�@&�x� Xq�"Ob�"���i�$�+dEs��H�"Ot	�Ѻ	�|P�㗖(���3U"O�)
�՚\�" �QD �J�$����ݥA���&m1�'P�d�d+�(ҢJ�G���ȓ�J���
1�nt��lC�>!�c�	��b"z�'|F9��x"H����jr��'^b�|���74�LA��T���1Q B@?g`��9G���D	�Q��% ���I.u�\E����
��t�6I
�%���D��	��\��	�&��	�W��ڷ$��a�H �-	���B�	�@D���1K�(5�qْ��a7��O�e�2(�g;��1d+���5�l8�' 2�Q{��N f-(�q��� ��[_r�$���bt��4���5�HEP��'�^$�F0����X�Oi�]���ș(Ҹ�(v [�>1�͹GL 4�q&�1���d�U�7�� ـK�e��!C�M�DP]��Z0�A,��P��P�'��Z���d��S��� ug��Y���h*�8�E,{��(��#m��B䉃�Ryb���ejR٢��d�OPъ�фg� Pp5��P
0!�"�Lu�0}1Ǝ�v!򤅤h�J9��@��Q����V�7kP\��(3��I�k�"|�' �r�NY�@�q�?] Ľj	�'Rx](-�
����3*�+O�ء!��D,��J)�I��F(�����
�:����=-K"��2'�U�!��3fx��Ш�AU�iI剘��9���	d��p=Y׉�1Q����jE�<ce�5��E؞� ���.��a��Γ�mh�/�79N5�a ��.9r��h<a�x4Jٰ�I���8�"�Pئ��B��i}2IL.v�IA��x3Hՠ�)̏7�e�AT�;�<���B�4EF�z�I�-`��'�����!���6��I��R�P�A+9�a�����$��(���7)�I��Z\Ҳ/ްjw$�d��78a��  U@�ʄ#<L�P��Kx�$�AP���<�lx�'�� ��IN�"!�tFA!4�D�b'B�D�Y��2�	���ӡ5�N�Z�bC	�E��R�ט �Ad�K��D�C>7'v%@P
O��s��ۡ ��p�T�ț[�s����TB�520�'䊰��
Q�C�����[� ��|�D�D:.��\j�N�g�ʬ����7��z�b:1�.��'B�)Q��Nfz�!a��	O�mz���(�Ć�8И������O�� ":�bH�3�u6)Ҏ	��)��}�B*f�>+� 5�I~*2���$O,��2�ֲvY*��b��9�FEk�$B*�rG%-^t��sN4O|1�3*��p���� �����uZ��[en�����O0*��|�$r�#�2V�V�2���� �7N^��c"2z�P�?�O���gϟ�h��Q0���;*��tYT�V�z������� xܼ��.�B|p�ڗ�.m��M ��)��lqt�v>}��������g�$k�`��7,O��ɏ?bK�8��^�Y�Z�%G�yT�m���E&��uGגeUn ��E�G(�SDےX}d5ƥ�b����mJ�	>5[r�A�ԑY%r��7%�.5���d6�L�u�W�T|�z��ٿ6]x��IUZ v�'e��D��㛵#��됅N�X�V 0d(5�q�M�R���%j�@E`�:H<a�	���9�p��d�D�`�|�4��O�xУ�.H�\�X�,�N���Q��?���Eg�h�d!H�u�A�6���!�ȇ-<��Z�R�@�"�����A�6�B��,�|3�Q�#��! ׏N`{�a�!L-3&�[윀s��@Y�Ǚ�`���#û!��'��gp�IkV�ͯ|6"�s�j֥������cW�0۶�cZ�|��O |h�f#�-~�m!�ڞGFl��v�H�"Z���r�+*�A��E�r#f	᥯��$�:TX�Sf�T��O���&�9�n�����AS`�ka�`BG�s�ֱ��b^�6j ¢�MI�0Ez�$�9/�	[��`��)��vk\���$EY��K��I�sz�u{A%ŭYLT$�� Y=f���#�'w�g����g�<�v(3�"�k��X�Z�HĉJ��n+�bs,Ӹtx���+ĝ<��ͧ3�*�C�'�F��[/@���7�	U��@�ӥ�
'�,p*#嘅27�c�@!&�LM�S�TU,[ʄű��A�c�9�g��\فլ�>��k���|Ӣ�ˡ�U�YΌ��SI`�>�[���5q?�'^T 9����UzhV�_�yȢ�'�p��c�3����Mh�1Fq��4
���F��e��kT�Q�<�0��hn�>�O��awC�_2�� ��ͼb�j�+�|��M�c�f�d��w�Q>�I��";`�92ER�^[>pq ��{�LArC!Qa~��(PK���Տ��_"��s�g�*��~���D��{���"`�\~2F�<D����נD1V��P@ʹ�y�H��1A"�Ϳ\K|�s�bM��?�p��% ���D�;Q'� :K���~� f��P�Qd8�}�iޯh\`�t"O�<)q��@�
�j3'�c`�	�2�L������C�%+�3��՚sY��i����	w&���EƏ4qOL@��ǈ���Ԕ��Ԗx�|�i�+?�丫QMU�&gDq�gk��0?q��ܡ0o4�Je	�.tVT���V��K>��iq���T�IU|����>�����5*��;�ɜ(3G8����\hh<��l�q:�g��Ϭâ�տKʼ�!�A�?rdb�CЌ�0-X\��>�Q�ϵ�l
�C[i���E3<Oh:5�l�� �O,I{A*C*̦%Q�͖�ER*I�"O�Y�5�і&�͋u+N�n���[7�|R���k���G*E�Oz�ň�d��j޴�����~��B�'�b���
�rѳ7ؾl��eqF��/O:��'�a�"��>!É	v0���)��V�pâDJh<�%�Ҹ��`�hL��%��?|dxr�	(��o�|� 0�2O �!!�A2��'����ТT:B����X�X�P��	ϓU>N��w�Y�[�T6M]^� �iр�f�4 �����P����:7������r4�7LO���C)K
\!�f����*�|�&���@�
�Z8p��� n"��qI�+���CVV��Yd�ګ/_�)Ja�� >fC㉠�nT���Q�x��t��гBb ��5*u�^�K�hRV�B����Ѣ����!	�<[d���Z@}�R�G6�!�$��|��:��,l2���CS�wJ8���߮4����VA�\3,�)�$ӫ}��*��O0�O�H�b�A{�v(�7����|�9��'��T��@d��@J���V��ؔ�|��ώ�uܴP U�N����<˥,U�MеC���Frџp8�l��Re"h�N>,��I"���AGl�bʟ�R`�h����&��	�'���3���JJQz� 6����*O.uũ�Q�h���K(&��<�U
�F�'h{�AYW�ȗ: �%�P�C��D��
^�z�DD����H�
j:*���E� 4B<�!���O�����c�[�)9��'&|�B E]	W�V���
���
���2bG�^�� ��A�h�|��MF�~���(��J3;,�VȆ��t��',�2W��=�f}X��,!�:d���d��J�����F�:�lZ, �6x��b� rn�HrG_��D99�"���O�@����m!��0gΑG9p���i<V��mE��)��'��Pё
�l ��k��)vj���E�G/i��h"�e��`!�$��9@�=�G�M�H��*࣐�A�^3�̀�4Iݣ9 1ԧu�o1�qOn7gY�n@��RKQ�	?z�k�O"�Ox��g`�\��1��ĉZ�<��"�@0tt�:,�oN!�D�,"�>�R��T�$��v*�\����2խ�dR��j/��~��g�L n�DC��.��C�I���� D3:{�-!��n���@.>T�3����)�'O�X"�
�G>��f�0�v9�
�'#��I�b{B�� �N+R��*O��!զB87j�@˓q��!�Y7������
���	�}�� ���P�z�Lc��/d��Ya���P�Ɠ<��2�A�+E܂��AP� �E}ң�-2PE���Q<7�
���Y�R��!�7)���y".�=#�向���UP�y�ƀW-�yr��e���ر�N�8����ǡ["�yb�1]+FY�m�=�P�P�%�y���#���e���6P�w'ߓ�yb����a��-��'Fm`�nG�yb�ɤ�.�#����m�J�۶�1�y"�I]���R`�(MX����M��yҧhVh����<E=>uqP���y� }a�	��@R��`�ę�yҥă9@��A/»JXi��"׸�y"/�@6�cǌ�?P�X(7*2�y�l�"�Ys�S~T����Ɓ��y��Wڲ]k0�[�t�����ɨ�y�ޞljm+�
_�u9mh��*�y�oڒ�d�R� ^�>#������y"g�"M�nx
vE g�Mx��9�yr���X-b7��o�T�Ң���y�oBVLū��9I�1 )�y
� ���H���!//W�r�"O�����y����&(�	LFIZ1"O��'�-���͑3mJn0�Q"O�%�ꑐ4�>[�[�#�D�6"O���%`��k��u�Z�8��٘t"O
�)��>T*�EC�%�ά "Ozq� ��.wNY��͒.?���"Oz��5*���{GkR"x+�]9�"O����)�"�� �A.'�,Q�"OB��HU�E4�J�'�#I��"O��r�*�m�'�"���"O���t�ڲ$A�j����pT"O$��Y'b�6���׏t^Ĺ�"O�Ƭ��T��#��@��ۧ"O�yy�A�� � ʒ�9I<y�"OH���&�dt
	Pd�͟g[>%�"O�ȥ���mf�!F�@Gd�d"O��`u�Q�0' ���O�@�"O.�׈L21�*�	����Xq+P"O�5�$��9(�����o)� x�"Oj��a ��@�`��1����"Oz��0��h�RM*`K�NA�"O(�襤��	\�ЊF홗)�Ĉ��"Ob�"p'��4x�g+Є� s�"O���S��$Ir�U�2���C`"OD��O>Vv!r�Voj0�3"O.�PbM�JD��M��M �H"O�Y1��1�$��˄�H(�f"O�-��oF�/RH%Y%�d.����"O �؃P�~�f�he(u0.�)�"O8�;%o�0���J+Y)B�)&"O.��cꙵ ��- #Û�<,�4�Q"Oh����z��Tza�_D=^��&"O���施9�NXxWMM(m-©P"OJ�c���t����T-�5P��[$"Op�Cq,ފlw�X�T�.s�06"OM��S=$�|��_	ʥP�"O�:��_5af,���Gc�~8K#"O��@w��/{P��F��>T�M�Q"O8��b�@%>�D�hǂ�:l���"O*�)�jU�Q/"y�ׂ@�7s� �"O��q�[1F����ψ�N% �"OĴ��ȷi���eoʹM����"O�Y(" K���Y{D,�.8����C"O�t�6σ�S ٫�f��~��"OV�R2�G�\�����%��^IJ�
s"O�9��D�zyd(c���95$�Z�"O�e��
�>�j�޵b���"O��Ѭ���@�c
�F���c�"O:q�'΃�'Wd�(��u�,��"O6��T��%(P&�@7ƃ/(�2(��"ON)��OU`���ֻf�����"O�����>����"O䩀I_�N`QZ��޶+���H@"O���jf(�jE+�frD@S"O*���n�] �+t+D�H�"OY�j>
�@9h1C�>U2h@�"O-a���A���R� �?^���6"OL�b���!j��m�8K�@(�"Ob|(U���D��8�l�EO8�)"O�٨E���CV�P�k;a(Ղ�"ORmqҏ:���B��Z%>�i"O�1[�S�(�9
 ��8�^���"OxuC6+O �$���G�`2 "O� ��;F�dY4h�b*Ώ~�$��"O�4rG�
RF�I�[�Ws���p"O�i���0w��!�$Lakd,a�"O�l���T?PK�պ4��;sS�](�"OZ�C�HR�v>� RA�N�[�l`"Onh87��K�pm�6HXZ3d��"O��׃T3�� �琝t'4Ht"O.D� AԕQ1^ūpF��}���`"O���KݱK}.D�#O76�r�"OL} N�&�N5�d(�*�����LH�C�#�Sdd ��:@@��qSiP�yͦ��ȓw9X��g�<p�v���'Y j��R�#ř{D�'��1��P�b��jJ|S�,�9�x1�&4�h�U�*c�a�Q,^�5N<�Q$0T\�BF�'�桇�#_;����D�����BOy�V��DD����[CNz�R�I�/u&�3ǟ�
B��"�8�BC䉛R��-`�Ѥ�4��v`\p�8�O0����]v� �=�R�n,`6h�/Қ)�Q`-a��Յ�a֢ R�`�?w���2����i��#`
�P�'h���>�5�¶��Hhr Tk�9���gh<��*ܛ6㎙�©�|�L��^>*�̕	�n�:(�����kj8�2M�.'�0�S�&Ͻ&����I.%� �ffN�"����D �AJ�f�s.%� �FRQ�ȓ9k�Ձq.��L`�p��i��M��p%�t���N��l���]�O�@��A���ԩ�!���4 	�'V� T��(&{�����<��0�O�B���O�q:��3?�BB�kB�ԉ%͗; ��HX���H�<��*�!�JA�7���S�8 �j�i��"�Ba}�+�C��4��A�U���'�� �y�L�0c��!w�
�Oq��"��J��y�)�gƪ� W%�Vf=Rq�M��y��݂pf�yrkߧE��S�D��y�'�=����H�P�1b�X $X���ȓ(��ai���5KT
u)񅛵LkP���v�h=P�NN�H{9!�&�3H�V��ȓ��E�AiY,H�t��b��*Ʉ�:���aa�UwJf�`t�( '���|�����̑X�Ă�
�)��\�ȓk(�(t$
9Z�.T�m֍WbP��ȓv��l ��x�:�Ȁ�U�q�`͇ȓ��Q;ᨕ�_BX�v)��HM�ȓrf\	y4�Y�����<��`�ȓ&��jq���N�K��?h�G2�E��Z�&�`�+B�B$���ְ�� ��d&|�1O,D��GG�;:.dAU�.SE2q�%P���1�K+`,r��Ov��CV�R��6���*�Y^d���E�8�;O^��d_�T6�,Dm)nf��A¥D�J���AEcɲC���v�&^H�%�Y�#j[`j��/�x�`Hʉ��q��	��Dqڼ��ɔ���d��	��I��J)�T�%�.�.��nڌ�Px�P�H���d��j;V@a�C���O괉fg�������>�k&�>�ūی/z6�3���5��d���^���'p�l�#��S{���K�k�jP��`Q����G(�Oꖂt��a�4�Z*(�,�5쟽}�uwO�L����Bi�[������u��I��Jۨ+�,	�-O�M�M_��2��ʐ1~A၍6�Y�ƀ�9Hp	�ǌ[��q��±/�(���Ŗs�t���4�2��Z��Q����yb�@� \�`8�*Үn7Ĵa��3U�� �d1O��(s-:T�|Y�]Fځڄ� �Ȭ"��>��hbR��Gt )O��#�ȗzX�q��d��G/�8H��ϸvh��@�*J��p ��xGK/R���WŕN��1w�|Җg]"�h9�% �I&���@4'�~h��k�_����\�Tt�H�\��4B�b�;��)�E�5�|��ejO�/�i��:�V|3��7��}�琧y+��S�$U��*C�Ɉ?Urc7M�q?H��/	5���s��G�uԀ�p7#�y���x�(�9v��j��m3�Fѕ��I��W�T!��>7(�K`� �$aT���	pydD p?䌋2;�� Ix��3��P%mg�#�d �1���L�<R'�HQiq��'�2�*^�y�Mr����n�T��K>y��>l�Z����Z��(��	
� ~%Xb�ܧU0��k��t�\���V�#�ar��'�Z9SA�B$8�,ŭ�+�x��b
ղ�,@&����O(��0�+kºU�'��uѴ���x�VI���B�.��<��'��=��Ĕ}4�bC�r90��8NHqp�'��5��������F�GL6�#^U�+����T��Q"O5�׊;��,8у�/�vD{U'т{��Z��V�/�3�d	�L�d`�IX�!�E�󁕢PXqO ���
Ѩ����l���� ��yb�%W�lR����
IV9`���0?i'k��NY���Iv6�� ��t��1H>� %�S�d��)�^\���>)6���!���ʿz�R��w	�Ah<y��A�o|�FH�w� �ٳ�_;{��!�&�0sm��p�K<I���>�HP,ą��ЈB�c��0fH<<O����Xf�� �O��8vl�0K3��a�@�!(+d��"O�Ec���
h|LEa�\p��w�|b�LYh���t�O`^��4�Q�v����A�R�~:PS�'���ęb�`�Eh�7y��}X6
M#BK��'�(�p��>���W?J;L��7m�Q���+"DErh<��L
�b�lT���T�I�4���J��Ȫ�I�G'�N�l�&^�\� 1O���D#W���'�z-x��a�`q���:��8q�`�lQ�w�9��6-د�
,	g���f��q$2,��I9���rt~6�Q,|<��a��1LO��(!n��9��D!��[�x� �|�D�X�v��p���2��Ӫ�AJT]�u,	e�� .�4s���Č
z�"�D�fS`B�ɧm�,�c��#+�rq�Cʇ�kri�6�b���K���,kzD�0m�K�vq�!G�}�����yG(^t��ŀV�H��-��y�낳 ��  ��N�Vt�Cb� �(83"n�1�h�٤�ŕ8(�90���!��(�'O��'��T(ƂM< r��fg�"7�|\����|H���/[O~�;�Ě�ilZ��j@o"Պ��91I�Y���*��y2��/(�0���U�Z��!� \���O�T��
�QSdm2w$�uq��耫�g�F$��$�*=���T��\-�Յ�U��&�7v���J2�^��~)�'��%��kH���m���:h��!˒�=��SB���P7<CF�ir�S?�B�ɩ[/L�1�I��DQb���*ݎ���b�V���9���t��<��M(��`(��!!��p���8ڸMR�㇗a������0LAz!��N����C�ܴ3.�f�[>G�D�Ä�،?�U[���>e ���	�/{����j"N�h&K֣�<�=��@K�82�t��M�KQvd�CGA�'��!��'j�F\��k[>B�!/����A��-��,k`�R����[(|�Q�"ϳ�~⅐��@��0��D�.����9pU�d���F�2C�	���%4F�U�p ��aPSG��	2Aa�1yU��JA �O���I+�'w�x���5wPh�S�(�8��	�)�6�с��h�9tl�'S��J$OL������ $�� ȇF⊄/�qq�B;Fjў�1t�@�	��	!'�I�{9��U	�X�²@�S!�$�1m����`��p�d�TN�(D�
��9
� Hg�@��+x49�&C�A�xl��4��0���2l{wL �|.Ba#�ϑx]ą�'=��8�m\>D+�q��I�I�P�B�R r�r�r���d1���Ѳ��Y�ʂ`�H�V�Ž[�
qz�j@,w.B�ɿZ��%z�oWF�^E;�L�$O̢>���ܢF�t#|e��:bv�Z$�F *�V	�4"[�<��93�����M!
h~h�k�R�<���S�JslՓ���" ��pJN�<Ѷ鑷�����F�
�4�(c�
J�<�"�޴��J��.sȠ�`D�l�<q�I�y�VI�ɩZ��!X��k�<y�Ȋ^ԍg�9�Z|����z�<!H�>i�:Z���?��1
Z�<ɀ�Ӵo<�� �)ԲI2_Q�<�e�Ƽ3O��(#� �Δ�i
�M�<���x|B �"a��%��!)���B�<��cχ6 �#��x?^���N|�<YC�#ɰ�Ao�8r�>��	~�<��R%^���*��ɴHT�X�m�~�<Q���-߲��Q�˳#�8, skb�<� X"E��`�D;`��O�v���"O��`V$dIs0
f�p�'"O����)�����_�o��A�"O��KjƸ0���ƀ6�P��"OԬv��{��xքo���JԞ�yBF�2�V�'k��`�� ����y�C��K�V�8��.U�N�� �Z��y��;^! 	1�B�N�� ��*�y2� P�:)����B	���w@ӝ�y����1�b���
��1�\s�!��y"��~iֆއ+��qg9�y��H)8�<���$��5Yea�?�y�F�;g�����o���h5�C��yb��7@Ĉ��@�70*�4��/�'?4(���m	0@{�l3.���ybk�A��b�i�'w�,����yB��b�`"���Y�M�#�Ê�y2�$�\{V*:� 9Y����y�P�o�e�K�]gV}9E��0�y�)^�`<jAb(тM��T��G��y���b|1��R�=�:�!PC?�y"	^c�(��e!��8#&u���V��y��KbP�f���D����^��y	\�,�r����Q'�tH�����y�8N@��0��:g�@Ɗ��ăP��(����f#R�R�&A#BC��ru�)o7 Q!U��[�	X�m�#r���Z�'��n�Ve���0}��k�F���S3ae���tT�-���ξi�"�'� S�gW}�A���gUbh���%\� 8�ጘX�R�>�.应 ��fɧ(���3��ִ{��9ʴ��<\�,�`�'�nI��#L�ɧ��x��P
�&��8KWk_��a�HūƤ�[���b�.�����֡�:_���H>D���7HشC�~��I� Ov���h<D�|�.�8�qAw+A,x��`�.D�HK!�B}�M�&�"H��Pd:D����`۾G��*�=U���##!8T�H�I9��rM�~@�DK3"O��:P�U?muh��skD�+NM)&�i���iQvG�8*�,J(�R!�a
�j!�D�2NS�iHB�.(������.F�!�dT�-���)��P���Dt 1 �'Y��AH\�z�6qkc-��65��i�'���� ���X`����ލ-c�@��'�4 ��=Tj\��oD�!�̜0�'�h��+�4j��c�!S�W��'��Eۆ��>)�� &T�e�LK	�'$���b�.�y���4�DEj�'���c��?#�ް����F��Z�'�`�# �<"��Q #]�p�����'z�����Utt	�Bp�Z��
�'�u:b%��?�j P��ٝZ����'v(�#�4e���V��L� Q��'�*��8���5)C*B P=C�'xLe)ǎ'4E�4����NHAa�'�<<��a�)T�x9`��-M�By#�'Vy8E�ܖP�@�S&�J�K���	�'G���c�kH<*�F�oS���	�'t2���Ս��iBƈx�B%��'ݨ�J��D>H���k�����'�
�[pM�-X���aJ�_3����'�0���"3
&�0,G� C���'��=�'�'i��W�	�Y�1Z	�'J4C��ɸ5|�L�7�óy����'E>���|c�(QV�8!��k�'�v��%���C��Ԋ��^�{t0���� �0Sfd����a�jX^S�I�"O�А�M�A�b��a�<4��e"O�a��GMs�l4�4�D�8���"OVi�d�4N���؅'�z��dI�"O�H����(�4����+�t4:3"OL���Ȳo�`��T%2>�L��"O,�*�b>Z9"��ř�٦!!�"O`���� ���d*�t IS"O��)��*H[V�����-�9R"O8�b�gӧ~��X�g��v�%;�"O\�C�L�3b��teΎF
�A�"O6�c�ՒF^$T:���J<"b"Op=A1쎒%���{���H����E"O�}s`�ˑHP-�#�f�:q�A"O8�(�֑+�d��vg�(��u"O����F�R`E�F�Q�m��Y"O(9�ލA�>}sq�3�\("6"O0�� ۸W㦙:`$�!w���s"OQh"�y����J�"O�X��H�z2�h�C��rN6a��"O֐���M	1����,����"Or!�v��JF��K��!����w"O�M`g��P���_iƭk�"O&9��D��m)c��fV� �"O���9L������'>%��Ñ"Oj|9q �?j�TZ���_ <�`"ON}AtG�bhq�7��i�"OČ�ƥā]��CE��xl�0�G"O&�z Oȍd�ڭz��۾O��y�"O`Hh�5nfblzÆ������!"O4��rON�W���� Kc����"O�p�Q9�DY�B�$-�8a�"O���O�:p�T������z5"O�����R����S#D#"҅r�"O�t1��\>a<�Ƀa_6� ��c"O��ÇZ6>�pP�ے!��d �"O�|�B���6���h��&�r���"Ot �S��Pvh���@���6�[�"O�CU�X�p�9�`��<�H4�3"O2l="��#��R)x
R��c��'�yR'��Z�(��CK[i.�1f�-�y�o�O�RD�� d�LJ��C��y��ߺKѢyj�AL4EFq���1�y"O�<���J�g���`�*��yr��0s��f�W�	Q�,��J��yjU6Nn3p �{���R�(0�Py�|��u����4(�6EP��j�<�FB�b�>��C��B'�t�҉�Z�<����P⚽���ݭ��); �Jm�<�fdح(A�4a�*
�5���XM�<"�E"�%φ�Z6�� ��BL�<y�(�� jb����6(\�HBI�N�<�K��8!�D
�J�.}���z�I�<Q�� V�i���#O�8) ��Y�<��E�i�
�.Ü1_�}�G�<9���!(U���T�<΂���|�<��m�*�:��q葻{q��c��]R�<� .�-��u�I7�mS���s�<Ƀ>=�ɨB�0b�ܘ�"�t�<�/�tw�\�4�.E���*�"E�<aAҔH@�!E��!]A�iR��D�<�� ��ő�"�6/����r��x�<���9U�؉��i�?9���m�]�<����{���P��g*�E���D[�<� :��wA� 2��R�F9J�� "O�a���'(&8 +��>װ)p�"Oa�3���ga��&���(�� �'"O %�%��r� T*vd�5|�j �"O��!�(!(0�p��S�t��{"O�=��CB%�	��Ndb�l�v"OB�Y�$�{�p| ��CW��Ʉ"O�5�v菈$P\��&�T�F2\ �"O&��:w�E����2A��o,D�hPSȃ�cvРc'|�r� D�ܢ�Oo��}�4h�7"���#�>D��h���"*�pȣ��
#,�iX&�<D��S�b�*��!y�g�- ��ɶ�<D��A@ЪS��y#A��!�E��L D�����Ϋ���U�rɺU
2D�4���xતy��f�8�QB""D�d�3E�Z^���!`W�Ip  �?D�ġ�l���d�6�±=��Д�7D��A�M��G,:a󆀖T.����:D��h�+ňV;�Ԁ'i�2\��X���9D��P���
E��8�����c�
:D���M��H��,�#�*�(´�%D�,pa�_V:� e�#h骐��#D�(����QI̞,}�81aԮ#D���'どSyp݂g���xB�!���!D�H�!��#��r�F�=��A1��?D�DyХ̷IU�I���{�
�p�,+D��o	��r�����'
g�H� M>D�xz#�~�e1Ң�5Hа�V<D���FN��S�!�6�|:�L$D�X%)_$C�(�CE�x��b!D���U�Ƽ|�\K�D�Ò%Yp�;D����@�I��c�T3Y���'.;D�(
FF�L�+3%^,�`��:D�sAf�
�8I��hϭtS4y�k>D��#�WtI Q����2��DH2D��A�D��I��18��@))��K:D�p`� ҙ,7��Ӧ	]84l�����;D��I���-����f��*G� Q��9D��C����R�Ύe��P���$D�p�sO�j\�9�dM�\2�i�� D�Ġ'�s�ƽ��'J[9���	<D��ŉH�5��U�G��6 ��Ym9D� s&fF�H��D�	�$"��Y`�7D�8�'�u�T��3d�3�T����'D�L8��x�	�JI�DTD98b�&D�Բ�n_�m������ž@yh�$#D��
C��:(n�i�Ў�Y�z�%D������J��h��?d"i @�!D���O�+��d�dBG�"9H�z�;D��1��P�c��U�E=%<�1�9D�����E�+��X&��L:D�pX�n����a���9���q�*D�,��A�0����Ԯm���#)D�y���
6���H�w�`4��O%D��* �N���Ҥ-|�6��ҥ!D�h�1��?��H1��
�N�$�8u3D�T��̒NzƸQ_�$�T4W��C�I=[�x-5�։j"�=z���p"O�8R�ͼ
J��L7(��"Op�*�F	T��u��悖$:��"�"O�;�E�N4ά��/�O�F�G"O�!�#�V�&9vL����&m�hb�"O`��@&E=*Q҂c�b���Z&"O� \%�c��*"�%�a4>�@e+�"O�I���p����p�jL�g"O�0��._�;���礐�$.�y�"O��7˘J�m�D��J6��""O�L�h΁���7�7?|�"�"O�b&�wP����� 8�DY�"OV<Ɇ�\5`����P���r1"O��THݵj����Ј3�N��"O^-;�G�&�<��û&��!��"Oac�oG�J���&�
|�:�k�"O�mÁNY)Q �H�\ 3�2e�"OP%ipg
q���2$ڕW��=A"O�@A���8Ed	VC�f�}J�"O�AQp���#�СT%qH<S�"OrS�T��6����TZb	;�"O����֙_���y��1I����"O�|��5�6�h&	�,3�a)P"O�(r�@As��`��Q)�Y��"OJ��BdZ�7Z�L��o��>��0�"O�l�%�:t��9���ƀ`�f�#"O���ƣԍB�0��Եa�:��v"Ot,@w�O�L�$I	��
$�dL�@"O�zԫK�[f�����B�_�~��"O����i9L��0z&��,���Kq"OP}�+	�` ]`�O�&H�t��"O4)ɱ�֓*^�	����j+>�au"O�x�ՎTBT�s4�޺o8`q"O���Β�d�����#48"�z"OT#b]1L�^�����/d2@���"O�!�!� ���k��QRn�B�"Or�
�Nʖ>���o�&�Q�"O�%B�!S@��A��a)+�a �"O�� ��9��l���T�OR-��"O�%!�!��T�*幕���oZ��SS"O�Pᦩ�|"Hi�A�.�`D�W"O��q3�V����U���r�=�5"O��RN�m������'mEP�S�"O��`�W�S�A���R,�吳"O$���G0.�n� 1f�4v���"O�i�wE�>��b;<����V"O��;��ˊt��W�#~b�:w"O�2�(T�s�P s�E�5z:Ĺ6"O�� ®�L|�,WG��Փ�"O���G   ��     �  B  �  m*  �5  yA  	M  �X  ~d  7n  �w  ��  ͋  g�  ��  �  o�  ��  ��  b�  ��  '�  ��  ��  '�  k�  ��   �  B�  ��    �
 � � �" �* z1 (: B J OP �V oZ  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p���hO�>U2��F1C4ӡ%B�>��eW�%D�����9]����"8�
mS�#D�th���*��6��4��$#D�\��2~F��u
�!.���sA D����ýe������[�<�����?D�@�w%��&�f�SS%D��8a!�(D�HY&N�1V�ȥ���V&D�A�`!�	�#��yr�C>s|D劥o^2;#y�Qk��Px�K�{�T�:���(8��+�#$����>iS�'lO�m���KTѐsF�W�ճ��'�铤�$ũN���rć:5�@3"��)rm!�P-s�h3eH�r�xb⪙�j�!�䈾�Bl�*ݎzp��a2c�1Y�!��8$�N9�%�D#f?��
�#��y�!�$R*l���2�Ɵ�1���8cǈV!���+ D�
�dV�e"⼐Fip!�$�8p�,�7�֐:$��`H�;�!��vM��­�@�0��/Et!�ĚYゼY@!҃&���K�f��l�!�� ,.�T�%rd$�4�]<~!�䛱���kah�f\삑�M<+`!���8�e��2G,%s�FS�gI!�� ~��d�)b4��ci��.�2�"O�a�L�I��=@Dg�0��TP"O�1���F�nؘA�5^�
���*O��(�NB4)�xt�θNy�:	��Ms�O�ݒ��hҊ�Q Ў!�ZM�"O�������@K�ux6Q���{�O˦�l�+E�x�Q�đ2 Na�	�'٬D9e��91��p�X$>��a��'�б�Q����i�&D ;? $��'͢\"�b�^�@!`�A70uش�~"�Pc8�@SD�?(31���T�j	���?\OB���$�`s8�Xt�����I�f�!�D_�)��#��R8�$=[���F��'Mў�>]@EÜ� ��9z#Ï1�̐ .?D�X�h�%;��hK�ɚk���F D�*$J�)" � I�3*�q'�9D�L��l�K�d<�7�1<�5xү3D��q3O��%pafӀ)R��p�/D���f��J������Ib"���-D�L� R.أ#�	�D�*u�7@+D��8R&R�2���B*^,�Tk�k5D���3
L0�,��f�1(��xC��t��=E�ܴe����Q�0�Z�(�N˖|���ȓ[��}(�h�0"��_�Y �0��j��s&�O @�B�I���@p�P���F~���`F��%�^�7��H�ӳ�y��9P�����:Dql9�F���y��N�'�4[�IE�%ߘ��E�̥�y" h�^�ڇ��5�-�'�yR	 ����P�S?`*y�����ySc8P�{��`���'��y"�U�S$�R�$b��z�K&�y��X�rm��"��\}&�I� +�y�)>1��E���O�H���؟Ǹ'�ў���a"QF�D�A$���;�"O����7��<�2��5c,dts�~����BAH�8�YPg�rhR����y�$�ޘcF�U�n���^��?qQ)=�ONa����ph6��F좱pe"O�e�/���Ukֶc�I��"O���茰+�j|����vp�d4�S��z��X�W {E4�(�&�DhC��2z��iH4�l%��7|�\C�	l��2�利@��MR���z'HC�I�)r�(z���$㠝c��+�FC�	�L��<�����Wl-s�D�$2C�I�]��%��� �X!�BE��ybgH�(�L�g�� �&�Prm����d*�S�O�<��� ({��Ar&�T
#��t`
�'�<M2�g��h5�����	�'�0`!�(��&��`ժ���� 	�'%���7�L�RE�Q$FB��"�'��h�Wl�B��	�qO�+K��ea�'O��Ȱ�H�j"�y��W�>��z���'*fՉ�Q*y������gӄq�'6Ȍa��5��Y2nϤTTh�8��Dp�ޣ}�qb��T�6(��Ob��u.P^�<a!��Vp��ᨕIF��S�GbK$P��O?��B��*h�w�ۿm U�6(Y!�\s����?s��!��$�����>��M�+�����*@�Rm�#�e�<�b�5q�������1�|0'"O4t�2�մer2�/�(i���"O������<4}B���M��!C����2<O� ʅ���^#7
��bQ��];bOx�����&PP�,[��=��( �� $���`8��2����7Z�����>+��;W�=�O��A�'^�}��(�d�X7��<wR�52��HO���&��&X+�c"�r��$I�"OJ��`S�l�1O�
���W<O��=E�t�܉k�Z(ˉX��0Bd	�:�y�: +d��)ɰ\�`�� )T���Cݟ̇���	7G�I�<}���������<IR.��h1����%"�&���n�p�<�u��0Am���4�D�e���yĊ�e�<�W�J�I%�a���
BRV�١AF_�<aTE�TԤ)���=0�U!7�x�F{��逯L`�!#$�˯[�&e��	�"|�B�	j��e��޳�-SET��ɧI��I��~��hO����Ǆ�$L�rs�<8oڅX�'�d��'�4��b�d0Q.Y�f��n�W������m� `�z�nZydN�V��0=A7�%��$o��<Rŕ�,��K�肍M��듚p?���	c����e�E�mhb`а��}X�ԦO�<q��ѷa�pz�X�L���"O<p��C�	R���y�-*g�|B�'��O�c���Tyƚ����Z4�����0D�x#� ��@�:��������d1D��!�[����g��r%p%��/D�� ����7x���ʕ3Y����&-�	��Q��O��좷��'>i�`��o"��	�'
�A4i_�f�\ѓiD�3L�ّ�A,ʓ�h�����t��|f)*>z���t+�m�!�:�1gI�>} e����)�Op��r옺i��h�&ԠXw
"O�p�A/EJ��E&��Wg�-i"O8���R A�	&e��d?N$	0"O��C	qȜ8p�!1`�V"OlUAR �;I����.	�(h��"O6�$�ܻZqd8S4�L(��e�F"Oڥ"`��?bH����t�(5�s"Oй�&ǝ5n$�`vkA�"O2�Q�!�Z�|�o>1���"O� �r�E�1ಸ��͔�/�1�"O`,b�m؜��H�&��8�`��|M��jȞU�ƍ���Ǿ^o�8�ȓRBL�j��@>A>qKv�N�pńȓP�0Z��E�
C�s��!9����ȓ�Tڰ�š<����s�T7R���ȓ-ъ�J0�O,B4^�#�a0|�ڴ�ȓ5� �+�!;ЌS0e��Smf���G�\���
U���dO��&�h%�ȓS�Pe�4DTJ�Ve����*p��m�ȓa@�����[��q��G)�,��ȓSIl��+m{B�ѳ���H
�ԇȓm*�U�#�>;�`p��S�y(�������Q@M��}��-S%ƻ'*Ra�ȓt8����������P�>� ����@�A�A�7#O�S7D��+	���JR᳢G@q`�[��\B��ȓR��;�n�iP��J�:{ņ�?x$I�6	E���L�ES�2.���ȓk�`��3Oĉ�7G�p�4Q�ȓlA���Mլ9�ɳB���$4l��l�*��T B�Rf�P�̇+D�$Ņȓ[z�akFk�7tv��C޲C4|�ȓZ��5��^;d��;A��+��|�ȓ���G��%Lժ���[vhɅ�S�? ,�T��5M�<���"8=�"O���Aٓ8.�ᡧ�7B ���"O�%�X�F�+��B�/�F"O�T� �/f��\u`�89��Q"O��(q��uJ~�	6k��&���0�'�B�'U��'�R�'�b�'���'arP�$@�[��9�,�95����'C��''�'�2�'NB�'���'��lX7F����ȣ��ͷn��H��'+��'���'�R�'���'���'�ik��4+*��'C�|/8DF�'���'���'�r�'���'%��'�t��I��[���LV�+-�?A���?q��?q��?!��?y���?q��ؽ�����K�MX�O'�?Q���?����?����?����?)��?���N���p$̂�s�:��D���?����?����?����?����?q���?�B��*�~�i��Z+Z�Ő�����?9��?A��?����?9���?!���?�S�F�)�d9�C�ab��A�����?����?q��?���?1���?���?�0E��g��A�Q]0,-p̙q�� �?9���?����?A���?��?���?��!3,KHI�4��/M.������4�?9���?	��?���?A��?���?I��=�X���R�;rr�$E���?y���?a���?q��?����?����?	P��)n��LS�ĕ5>F���6)E��?���?9��?A��?���aG�6�'n�x.�3��|��p��@�-8���?�*O1��	��M�#�?q������¦Fr��,/`,4��'�6m0�i>�	��p�v��.E����w��`Ǐ�����-��5$���';��đ>�R�ӂdY��N��Tf̓�?�*Oj�}�0�^.8�����֘{78�R7m̋H��$�'��'�Hnz�5�Т_v�x�ĉe�n����Bӟ��I�<A�O1�����<1.� ��Y���ؑ���<��'^��D��hO���O֡� Aհ_���xZ9��2uʑ�<Y-OX�O.aoZ�,2b�4A�DZָ�b�뜂&S^Bo S��Z �Iݟ����<�O�4c@o��d�lS�_�W�d\ ��	�6�>��P�>�'Tl������dTC���i��
����]
�,i!Z���'��9O��Ђ/�?X�ań�.�Xh�:O��m?Ϛ�3|�V�4�8B�` �j���H aDc��R�9O���Ol���2�6�Ot���J� Ҹ;��I�&˔n!Z�(�B��}�"�OX�S�g̓W�� S�
*��r]
,n(�'h�7͟Z(��D�O��D*�Sxê�q`l�8#�jyxG&�	 �H��ODm���MC0�x��d.Ёx
z�h˕��\�f!P�:�p�B)A�7�剄@��R�u��|BR�T�e�O�m��}K�/D�
jK	�*Da|�a�}V$�O�t���^�l}v�k���9|�Tu�p��O��lZN�u���pnZ�M�It�4���Wt�L](��H9XZ�K>��R�1��^�S�ߙxr�	g�V�"P`#	�0��Oe�����3g^���W�=F��peC�TRj(��ϟp�	�M��AM�dBg�t�O4����՛@2DmJ�+�
'
�:�!#�$�O��4���3�''���4=b�G	�Y�����k�iM�A�"�P#|��IO��Py��d�/Rʦ�:�A��pd	%�� N��,�ܴ9	X,���?�����	T l�
l(#�
$1n����l�62������d�O��� ��?p͚���-Z�͊'+vi[����YP*�ş�����D�i?QI>!g�S\:�\��FU�C"�L�1�?I���?����?�|J.O�5mZ�[��DC.0A�IGA��@$ND_܆�$�Oڍn�F�/��I�M�N9M�ea@AE�S�d�	O�i�Ȅ��%3��œ@X^\0�'w���B�N�2�c��H-HјV��	ܼ����D�Ol���O��$�O��D�|�D(��r#.���̕c���u�ˎT��V�G P�I�t&?5�	�Mϻt3�E�ǋ�^x���Y�1��H"�i��6-�g�)�}���'������ wP ��ֆK���ٙ'L�A��&C?�N>q+O��C���Щl�6�i �O@�̄�I1�MK�d�?����?!Sb�"7��+�蘔)�.��@?��'� ��?)���J<�s��[�x�0�ȇm��)�'6������1C�t�E?���v��ْd�E1=�����������?���?���h�����|��ֆ�+��`�'eŦ]���d��e��۟��	��Mc���4���Y�Zφ�j��� AV��g��q�d�5�4A�����?X�Iퟴ���\�P	��B>9�,�W#T�x���ȓl�)a��O����O��xcaE�7�|K�-�JiP��0&i�n�r�'""�I[�p�P�����l	�@Ґ�'%�6�Ц��I<�|b��<ک:� 1wڄEJ�>,������/{��@��'&�'A�	<��T���*7.����N�f��ݟ��	ϟ�i>��' V7���F2v���C�pc�$F�&h��
E�g2��d_���?A�]���	�0sشp��U�7$��]����Ŋ�Q����d�,��Q0��w�����>��=� 4�y��^�d��Rd�T�{�2�+`4O���ć�K���+�gT 9@C+-�t��O,�DU��)�a�3B��i��'3�Ы��wP`���ܨB�Jt�(�d���� ��|�G�)��Ax�s�l�2T�:��,�z���O:I��ӟ�����O����O�dКk7���T�`i���w�W�\��O˓)��AC"C��'��V>uQ4HC<uhe��bݪ(3 �-?Q7^�����CO>��?M+��Ohf��wb	,k�v�x�eL�b�̓0���"��*��O�.6�D"Zz2��@�},��SC�Z�P���O����O��I�<q0�iC�pbQ�x�U�e	O,-�m�5vR�'.r6�$�I'���b�P���l��=޲C �0o�� F+�ڦ��ݴC��1�(OP��ޚk����	�0{�b7�=����r��O���	hy2�'92�'���'n�U>�Q���%f�8)�N�)*f�œd�ې�?�� ӟ��I���%?�����M�;rߌ�bgd�fL��צBTD#��'u��1���tꖎ{��I�1&��F�΃q����աbgt�� j�� �'X'���'�r�'��l�!�T�4⣣K��Mˆ��O����O�$�<���i ���'���'4.��k�=+h�{���;S�D ��F}��'�"�|r�\/D�*%�qZ�
��DT"0
8��f?�4�H<��'��NײO�a��L	�V�����l�"�'���'t��S�����'�0s 6@�&�6/|Xزg	�ޟ���4hb�����?��i��O�� ]Yܙ���Y<I�2�@ڄW����O�7-�A��ÝF�@���O���խ�.T>��q�)YO��!�Z͟��'C�i>�Iȟ���ϟ8�I23�(B��8~�bM`����Q�ba�'��7m�'z�"���O���<���OD��d��YЄ�tO���D�*Bx}��'B�g2��!j�����e�Z6���n���(�1�J]���	4-[��3��u��|P�P���="���'\�0lni� Hɟ��ɟ �	���pyBKo������O,��W�#Nm�'mD	O
����O~<o�A�F��������ğL��g�&"�ht�S�ը��̚$�*>O��'�bo�<k&��`���� ��/ N9���-%�9��;>����O��d�O*���O
��,��@�R�	�p؄Z aH�#q ��	џ���&�M��C�|*��!z�֙|"A�_������^�&��1
g2@O�o/�M[�����,O �����$��ԭYA��x�v*üZi:��5E�+�?�h'�$�<����?!���?��I͸�	���J'�@����)�?����d����#v@\Ο��ßt�S�?�V��QI��H ��<@��1?�#]�<b�4cܛ64�4���ɒW�v@��	(4��Z2#@�,���V�L�M#���ch�<Y�'"�.����O��C�ǝ@r��[�l�&a�(�ON���O���O1�(�*]���U�l��Pa����v5B�B�:0��f�'��E�X⟤ۭO��oږ�B� 6+_%��U`�gE?:��ts�48ƛV��\$��柌0F��$��dfEoy�Nٜy�Y�s!�nQ��x���&�y�]�@��şp�	���ӟ�OO4T��+�&a��}�f� fy��1'`�,U86L�On���O����D�Ц�*2��(!O.g�j��$C�K\b�)۴{$���9�4���i�����d�<A6f�'BK���� �I� \�0�	�%"l����']$'���'�b�'Զ����Y�]`�T5i�~4V�@�'#B�'�rQ�|��4C����?�����)��/�4*&�I�4����H>y��Z��I�M�i�FO����F�N%�ƨ�8����8O�Q��4Aa���O˓���<�I�q9��rC�¸i��(p�@�,[��\�����ʟP�It��y�&�=Oն�1�ɓ8�,��d��`�h���O�$즥'��s����]�o8��w�J
oT�*vOf����43����{ӆ�y@4���7N�0��'T�}�c��FG�q�"�M5<�TRd�9�d�<q���?y��?����?D�Mo��(�I�t�}�Q	J���$�঱�'ŃLyr�'���^>q��H��IR��K����+"����OXn#�M[��x�O���O��a�g��1�&�[���1;SNöm�RU�<"��L����#���<YAZ�{��piEzH�!)��=�?����?	��?ͧ���ԦA�C����s��I��P��Ô|J`Ѝ��H�޴�?�J>	3Y�H�	֟���15({P���0�����:I��D� y��'�$�[�l�E�+O��I�Ԣ�%P$,��qH��+�(p�78O��$�O��d�O��d�O�?tm]�R��J-+���������ٟ(j�4ydyϧ�?���i��'����S�m܄��h��ƞ|��'���'���X�^�0�'40��b�O&[�n,Hf�&h%�Ɋ'"�-�~�|�\����������� ����?�;Q�/N��ek�����	~yreu���!p%�O����O��'+M�=�c�
��ل{�(9�'����?������|���_���A&�f�@����q\1���4���O���M��D$��S񆁠s?���b�Σy�Ib�A��D�Iԟ��I��b>��'�b6-հyT|H�4��[
�/A�>����SE�<�զ�?a�[���I"0�4��B�6$�
0۾e��t��ȟB��ny�П������?͖�� �J+��R�M�싽;vL�x17O���?A���?Q��?����	A�ߒT�$,�a���JgfW)?^h�nZ'�U�I՟��I@�՟  ����3�"Z5�|�B�(�CJ�?������|���?��&��
�(C��b�Ꭺ&��$y�b&.�d�*��z�'��'x�����I(��h��DU�|c2=0Q���T\ @�Iݟ0�	ȟt�'IN7��D�D�O��$H���0���!��<��� 
�xH�O���O��O���&^�e���[ÇQ�~$�-PĞ��鷃O;�tZ �>ͧw:�����Č�~�JDy��gyt-��?v����O �d�O ��.�'�?�'��:�t��-g�8��2�G0�?Y�i�� h��'_�dhӒ���q�:@P�a��LH��L+�~�	��`��ş�p��D�I�t����O�:�`-���N�[�h�`�ny�O�R�'���'�RJ��y�~�a�Ԧ<0�T��.l�剆�M#����?���?QI~�� @�T �Ϟ
g�"���[�5�tq�P�������%��Sޟ��	��nXP�J/BN��We�3�ZM�PJ�
��Yg��
��O�7��<1�ΕT?��q1��/|@����ׄ�?����?���?ͧ��$�֦��qLȟ �iP�5�Pё�Q�����Sҟ�P�4��'��ꓦ?1���?)DJ��h��p���2.��CG?+%�M�(O���Y�"�z�'���?�]"L(,	�ًkV�b�䍈#H�ҟ$�I���柰�IO�')ҩ�"���`�RЈ�U]X����?�����& ޜ��I��$��:F�<^ ���S�p�xb��h�I՟��I���Lny��'�����ӳp׆(�U/Y�F�(@��kʄ7n2)�	�[��'l�i>��	��\�ɰy9,}�oX<}�8�4%	U��l�	�T�'b7mP�3�N��O��d�|rs��<Y�T�g*��!�4�H�a�O~��>I��?��xʟ�(��A�0R�2�8�.[9x����"1�dP�����i>m����u��|�M�~l|�!�Y^�����U�1��'��',��Z��۴j�X��s/�7@��:p��-5*�+SHΊ�?)��_�����i}R�'��9H@Z�����A��^N�"7�'?�7��%g���?Y -C�|}T��,}r�ӱo��y�s���L�
�P�yb[�H��ȟ��	���	ȟ �O�te�V�:�^E�!��?I3I�/tӲ�"Q��<�����?T��y�%w���ibm�
0T�ك�G�R���'ޒO�I�O���ʀQM��2�>��U�)t�l5��ĕG�ϓ^�����o�OV�yL>�/O��O6E�F�Xp˶�$I�Z{�1�J�O��D�O��Ŀ<A��i. q���'��'��㳧ߙ3w�2�Z.�����ĆC}��'�b�:��σ7�hal�2tp�gx���Ox(�'D>�p�O���Ӎ9Zw2�AK~��Ʈذ,���ä,�7I���'���'�"�S����a�T rjP�E�(|c^)��OʟԪ�4Z����?��i��O��;/���ȇ�
h9P*�z\�o��l�1�M[恏����O�R��:�����E�`��[dIsQ(���UK>Q,O��Op���O��d�O",����x��X6��_� ;q(�<�g�i,�4�'8"�'��@�"b�}�Q�C.˜.!�{e�\D}��'�2�|�Ou��'���ÈؗEے��%jRj1�A���V8*��U�Of�d�-�?�;�䓶�d5a��6�W�o�t�(Ѝِh>D���O(�d�O��4��ʓO0�v&ƣ�R
A�3�B�h%HƵg)~��b��� l���
)O|�Dt�^)lڒ[B6Nq�}8�Č� ��J�m�S�I� ��}) �O$q���.�i'���ᣏ�:MP �bV�r����O`���O���O��)��?qT�7��D����ԏ՟y��e��ԟ�	2�M��*�|���<ț�|��&)8�a����%����l̢Y��O��o��Mϧ"��!M>�u��0��S�nZ����Պ�#h\Q2���O�%�J>*O�⟨��\4c,E#q �lgF�x5`>����U
r�"�'�2S>	`�EO2��惀 5b$ 5�=?1$X� ����('��'��A�"E�����6,j*�낺�dq�����4�FԂ�' �'5XL��S�D� ���c`�q:�'*�'����O��I��Mۗ�Q�;�.yU��-�*u:�n	�U ���?��i�ɧ�4�>Y��*Tf
`�z��1�
 @F� Y���y2��
��Ӻ3��ٹ���\���D��~���(�֫@v ��os�T�'���'Ub�'��'�������N�i�$�*O�b4R��Wf60������o�S�8"������Ir��Q��,�h`��@��?�����|���?1������$��\`=K�l�0C ]�"��:L0�dֳC�b�'e�'��	ٟ���r�x؁"��q0<l��� `���ԟ�����Ȕ'n�6-\��d�O����<i��[��$�U��j�5|LN�`��O����O�O^�� ��A�Pr�M�
���P����L]�.�����y�1.����O���B�#�6�J�Ĕ�LF$�p��Ob�d�O��D�O,�}���0���Td�ȡc���J�h��[ʛ$�;��Ŷi��O��X�B$�'(���yRA��$5��$�O��D�O��!H�<I�k���H$��v�� ��@��T9�^E�Ď� GD���.�$�<ͧ�?����?����?�"�Z/|�y�4E��tp��k����$Ҧ�B�@џ��I��l&?���9'�̨�*�.�\��V�I�y<T��O����O�O���O��䙐4���)E��D+�"�xd����/�O��P>���K���$�ԕ'�(���C8������4���ar�'Z"�'Br���tW���۴m�p4��`:�{ Ϛ<eVX`"GcO�~�+��ܚݴ��'���?��e8��\57�ءx��ՍR���`b�����|Rb�
�A�SK�'��{#h�f~�P���I#?ӄ�i�j��<i���?a��?���?����ٝ)���J�֣�e�r�ݎ/�"�'��#~�>d���<Y�i?�'�b�Hq�[�"��`E���`����|B�'R�'D�*�^�8�'&)|]�pΐ�J�lsԣП,D0RR��%�~ґ|[�p�I�D�I埀��Rx�<�`@A\?�9�M��t�	my"x�v�d)�On��O��''�N �Gџ@���`�� �J�`�'2�듊?q�����|��\��A��R�6�`҄T3~|P���Ñ.��L�����������'M�'c(I��)����� Oh *!z��'��'B�O$�ɗ�M�(KDȔ�ՎM�l�dY�M	�Q1܅����?AW�i�ɧ�D��>�ir��R�P�?�VTi��O:"�|�)��p�zn	Sح�'�2�І?�TD�'��̕���[`NC:O���⃋/[L�D�<q��?���?A��?q(���1��(<fb9j��]�0 U��\ަ���l���I�H'?���M�; A$5w��¯�I*�����?	K>�|
��E���ĉ�nMj`LP�U�D u��>7.�֤5�@�j�'G�'��i>��I�O��S+]�;�1p1`^4]x��	���ʟ̗'��7m
�@�\��?V��"g욐hՠ�`�+���.���?	�T��hߴ&��� ��*:���`'��(9N(8��D�W�IQ�r�*�噠j�0�%?�2r��u��'e�R\tZ 5(���)���y��'�"�'���'I�>��I�~x�qJ�#�2qoD`��&��y�I(�M�)ƈ�?I�3���4���S'�/'O�US��Ҕ��<J�5O����OpEm>K<0�'$�)JX^1��:���b�#֭?�r���	�O�D+�|�W��ǟ��Iן(���x�I	d��82�߁7n
̓W�cy"�oӞ<�G��O���O���d������ƾ �� q�'T9Mi ��'�7�JЦ�"O<�'�*�'"(8dSte�[�I��Ǩ�W,D��?�/OphؖC��~b�|�^�8!�ǘ#"G4X2�Ӫ���w�ڟ��	ş<�I���jy2�b����N�O��Fgӻ8�*�pf(?bƴ3=OB�n�D�I��I��MŲi� 6�ߕQ��!@vC�		���qƈ� u%�P�*�<1�Lp� g�?�'����wj�Hq�P�l�{DJߩZ�}�'��'���'2�'���䁤��1~F���-Nd̑p���O8�D�Oʽn������'�\7�<�$
��(�d���2���a��P�T'��mZ)�M��'(1���*O���
�jϨlY3��$j�����Y����/���~R�|�T����ܟ��Iڟ`C�$��-�� �0gÌd�����Dy��hӤ�҆C�O,�D�O�' �q���� nQrܫ���(_G�y�'o ��?	�4�ɧ���|0p���mS��ɞ�&�FQ�8u���[���p�>�Č<	gDe��\k_Ft31�
�+����O����O���i�<ђ�i��a򉞤tǾ�c�͒&���i� ��&�B�'�R6M>�����Ħ��s/=*����E�
�TARRk�2�M�W�iw���0�|"���4ڬd�'���@4Pak�.��7.������t��<����?)���?����?a(�.� �K��	�F9� b/W�����lE˦	�Q��iy��'�O�R�w��n�Rtɸ���dn�P�Q��xͦdn���M+`�x����*I��	�x�F pG�G[�)�����I��ps��O��O���?��AB<��⏬c�ԁ��_x�a���?1��?�.O��l�E0�@�':�-ϝ*(�xFEM�I^����"��'�$�>Qc�i�6�K�pФ�EF�
 I6�(�ȑ7 b.�@mh�J
8>@�\2I~��j�O���O���F׾R�9���J�a���8��O2���O��D�OҢ}λ}���+^Z�9��5,Ҙ`Jwa������4�������?���i�ɧ��w�Z���iKL��K�m��X�5�'x�6M���eܴ"f�HK>�&�U#ʈ�i&A��a��`�����4J���^�YN>�,O���Ol��OL��O���V$S�q�X�X��<� �i�l�OB���"��T� ��s����̙q^�U�#l}��'���|�O1��' �	k�Ô� ��,��`	�.bv�U�6Q�'avm5&w?9M>1+O���H�P~biK�Ŗ�!.t��PJ�O�d�O$��O�ɤ<qջi�M"%�'|�i���&C8H��)�#%����t�'�,7&�4��\�'���'Bn�$�r���<��eQ�x�X�0�|�eј딹����'r�"��0E�:
.���q$�8e�е�I	�O|���k�<��[A�찙�G�0�	!�'�6q���K�/̸:��!#0�Af��@d������-�l���rzf�r��S�<aX��C�ί82Z=�G�5?��ǘ�]w�HsG�=[��ژAN�eٱf�3}p� X�D�O��]�%�]�_����f�4�ߒUf��3c�%р ��Su�@�,��A{W�-.Ş��B
=["4h���a��B�o�57`� ��G�0͠����':��	�� ��oO�TkvcH�Cd��C�9����i���'aB�>T�����O��Ɉ*,2H)7��z�D�p��LNxc��1ӦS�	���	�ȰN�|x���HW�<VP�!���M���%5 슥W�<�'�"�|ZcDX��'����O]$	4���O^�8%��O�˓�?���?y/O��!�ǎU�u��o��r�@E8D \3���'�	�P'���I��@v��:/���F�@��5q�-�(�$�����x�IKy��4KF�S�>Q��ҵ-�W;6���A8)&6��<�����?���?���'!��W��E�&�!Т̙�@�"�O�d�O����<��Č�E�� �G-�5�P�@GDˎ|��dP���Ms�����?y�
� 5Љ{B� %�>�S �ڙC�<1�W��M���?1+O1q�]R�$�'���O �Hl�l2l�!��ͼkq�qq�&-���O��H�
�㟨��3p���%=A.L��خ}>�nZAyr��p7-�O���ON���n}Zc
�}
Q�]��V���]S�LE��4�?��y��(������:;��T/M&}ؖ}�E��//țf�\�7-�Ov���O���R}}�[��%I�u�Q�e!�?u�rH�j�M��K'��'T��������bdW
h�&�L&c�>�l���I͟��$���D�<1��~�c��y�	k�g

v�T!�0	Y���'�D�Xd�|��'�b�'��u��hԹPT4�h%d[�z?v��(l����U�a�'��I���&��؇#6��PAK9���ZPh�=Ȭ�A�yq����d�Ox�d�OʓA]����1F �
� B%
$�1�&gJ/U�	ay��'��'��'ި��F�r#�Q  �F0L�x��J�sh�' �'9"R�@�ˉ����C�!�
��'�
u|�z!���M�/OR��4�D�OP�Ē�8��0�޸s�BN��ҡH�����ꓖ?����?�-On=B"��z�S�7�����SX�س��0G��ٴ�?�I>*O��S��O��O6rl�F�'F�
�IRM�}���4�?���dó+8�@'>����?�؆p}����b2|Ollq�^CRH6��<q���?�qk	��?	H~����aπ	��!@WMD�=G��{@�����'��i0r�}���O��O���gޤ�ɱʣm-��H��E1Pp�l�Ty�͋�&Rb'�i<��iy�Ȃjԕo��$_�V3�5I�4S���2ǽi�B�'I��O�O��G�9�0�6��91/��	c���t���nZ>3v���ٟ���ߟ��S��R>Ya���N�� �#�����hۛ�M#��?y�Lبis+O�Sv��ma(�e�̆:
j0�C��H��m�<)Em�7C�Ow"�'\�-�a@��V&F���E�� 8��7��OH-��(N@�i>���ܟ��'�)���%�v�`f$єpm:-���t�<�$_�k����<ͧ�?�*O���8�d�b��=�Di��.��b�o�<���?Ɉ�'b�i��(��ˌ	`uѕ$�=D ؠ��P��d�O����OTʓh�,%B�6��Ly׏\n�}��@'PRF0PtS���	�����by��'��! �" ��s޼,�U�N�$x%eH0IN���?9�����O�s҉�|���h^L*u-�&Q6��C��bU�БB�i��O����O�rB��9��'m.��EC�A�>��B�
-X���4�?�����D��&>����?��	xqv�# N�0ia�-v��#X7�<��?I�E���?IN~���C6[��^Muf�o%�hJ��Qަe�'�B�"(sӒ��O���Oh4�A9��gB��`A�S&@':7UoZ��I�t@T��ɫ��'�(����>v��1���X�m�>4cT 
9�M!�9?����'�r�'��d�2�4�k��YP�!1�ω�e�|12G�H�DK��'k�'��X������N�2�A�����RQ4��yo��8���@���Ҍ���|����?�vLU����4��Ri��!B��Wś��'�B�'I�	3��~�'��'�*J I�pk��	)^�"��A�i�F�$N�S��5%��̟���{yJ��,����$�F]�W��%t6��O��9]��|��'��\�XX�(�	`�\�{#"��Ԁ�?~� �I<���?Q������O~��QBv�� ���I������ӡR�E�G'�ONʓ�?����?1)O
�!v��|�e�]�K�FX��+��s�9Y�fBD}r�'(�'�ɟ����9 "��ie\H��G�l����B0Z�؜��*�>i��?Q.Op��:ns��'�?�ҐM�i�D�E$1-I"fJ������O~�@6"�:I�xR�[8�NP�p������C�M����?�+O���-�D�S�� �s�	[a╕zzݰ,C�N���17�!�$�<�C%	�?�J~��O����B
I�0�ֱ0)^0��O2�DO����D�O����O��)�<�;l�
<3�ʑwRtJ��lRTIo��D���N�D�u�5�)��|G�d�A�F� �̠x�I)U�7��%\<��l�h�����S����|*��+�s"�	aa����,D)r̛&O[*{`��'��IN�4\�x����tC��8�b0k��K Q0"��ݴ�?I���?IT
n���xy��'�����eJ�h�A�5(�rU�wn�&Uۛ&�'��'׆���)�O���O�)��cת��2��N�%|q��o����	w�<r�O�˓�?�,O����� DQÊ����p{#f^�-���a�i����y2�'!2�'F��'R� x�.����>Af��A�ԅl��E���°���<������O,�$�O]i6i�)���aj����lP*6���OB���O0�D�O�ʓ^��[�:�v�b��&+k���ab
Ѻ �iU�֟��'Tr�'[�'��yb��1�Y(e�8.�����W�V��7��O�D�Ot�d�<�6�Cc������<�:�I��1X��%5����7��O���?����?IwF@�<!���~⁘����!ȒO���r�A��MC��?Q*O��2T̑D��'y2�Ov"� �aš@˪���4�v��!"�>Q���?��v����Om�IH�QjK�V�J�mǉag� S�i̦i�'j�P2�oy�(�D�OT�D� קu��P&a�ƠCf�ӚW�,y���M����?�F���<	���-�ӟbr�� HW�V�y�rE�5QX6��<J�n���p�	ԟ��S7���<ɒI��8��ńL��i����֏C�y��'l��O���?��Гr����a�Ǚ}ۨ�CFbR�9 ���'8��'��#�h�>�)OB���4pg�Np�,�����yd�2�`����<���<�O��'�r��9j>��s�]�B4֭jc�v��7��O~��D�z}�[�x��wy���5��E
1�~�����gc�K��,����T,���@�Iٟ��	|y�k�hdr���O�0Y
�I��E���F�>�.O ��<����?	��S�!�����Q���ly�H�<)��?A��?i���$˪pF�1�'F�œ6g���ة��B�6v���lZ{y��'��	��(�	��@CM{���WÁ?RӨTã��211�Q'X��M���?���?!+Oz�hrjDX���'�H}٤�C��Ai��N�^���O`��d�<a���?Q��&S�@̓��i���j��B%��t:���+x�^�r�4�?A���L�в8�O���'���ɁD�R�RuGS� ����4�~��?����?�����<�K>Q�O�	HU.ř9��G*��o)0ݴ��č�y�HqoƟ,��ٟ�������Z@B�k�v��l0&_6v�z��i���'l�@ �'��'q�X�k��)����g$)�v�j��i3����Os���D�O��d��I�OX���O��"WMV!��;���>�h$��n�˦�A����p��͟ s�������^�]�^IӐ �8-~Ъ�4T�n�����ϟ�pT�
 ��$�<1���~����ov�y��. �@i����Ms���dɢ:�?	��؟���o�D�������3�D'CzX�"�4�?���A��ky�'��֘)f}�)�5��I��iЁ~���F�����?����?!��?�,OԼ{!���֤��R���	���b��>�,O����<���?���2��"`%ܰRn�)����QX�dꄦ��<!-O4���O`��������|���ʛ�j��?
	�౱�Aئ}�'>bV�x��ٟ��I�`~��I�76�-j5�<�p�g�4��0[�4�?I���?�����W
���O�Zc���$�
�3�~uv���@���hٴ�?9)ON�D�O��d�b����Op�Ċ������.��r�pcw���dZ*�n���|�ICyBl�K�h꧂?���"r�J(�H�ʰ�
T!�iـ$	*6�	Ɵ���Ɵ(���z�@�'��֟\�cUR)�@2�NW3zARb3�i��Ʌ[�=ڴ�?)���?���[A�i�A{�A9O�$rp&\�>)(��Gu����O�0OΠ��yB�	�t���	���%���
�j�����%2��6��OR���Ob�i^}R�@S��L�1S��C��E鹄�	��M�ah�@~�W���R��vc ����#�� b#O�C�^����i���'M�ҭ�������Op�I�	�����H ��6��S�$�6��O˓w��S���'ur�'�� 0W��4H�r��7�a4jx����(\~��'���۟��'�Zc��a(�'�
N�x�k��?ɲ��ON5:O��d�OB���Ox��<��	ǐZ @dE�Z��@��Vo�iBQ���'��U�����4���6O��@�1`�j�nQb�:�
`�c��I����	���	qy��2NR����p"�Fr��)Ë&?�7M�<Q����d�O��d�O�ыR7Obi��V�F�\��B �d(\Ij7����	ԟ�������'�S�n�~2��+��m��L�1U��p�7a��9�	QyB�'��'AD�'G�s���P�'����@ ��&z[�9�@�i#r�'	��d7n�����O��IC�p�K7#�;�����F.syR��' ��'cr�������#�0�y4��+A�$Z&7��(nZFy2h67�O"���O��)f}Zw�B,�K��vü!X��Y6=S��i�4�?���S���ϓ�䓅�O��0���p`�g�N�4���۴&|��Xưi���'���O3b�� �!(T���Ͻz��}+�'��MKD�<�O>)����'ц�Eē�\}�1�f�	�Iz\x��m~����On�DM:�H��>Y���~B-_�[X6��֛7��cI8�M�J>q���?�*O��d�O����TmZ��D�D,Lh�C.:h��io�I	5xO���OH�Okl�?��e�'+�-���2��?��I�4�i�	ay��'���'���r��HZ�m�/�luva� <��Z&�����?����䓟?��=6Fd���)/1����q�*�2�䓊?����?�*O���@��|
���%(��`��5ne��L�h}b�'�|r�'��h��$� ZuX��ՍO��Z��%i�x�qY�d��ҟ4�INyr�S���t���ЁF����a�}�Bm�Wn�ߦ��	t��	�����i�$A<���2�ݷI�x4���qu�f�'"Y�������'�?)�'�d[� �	,�����Px+���f�xR�'���߮�y�|�ݟ�,K��7"P�B��M%j2��i(�8�v�0ٴXJ�П8�����ÑzdJ}���B�@����&�G,(7�F�'��%��yb�|�iV�J��pI�CR9i� �F�(8��( �.jp6�O���O��I�N�I���B�n�z$�[%"�d�XŴi.\<��'��'�Z�$E�֮5��oW:-����E�8m����	�����-��'�R�Ov�ꖤG\�  & 9eX��ӳi��'���b5�'�i�O��D�O��'&U�8Ј����G�F#"�Ǧ��	#q�:���}��'�ɧ5F�Z�J�q��/{��,٦�Ǯ��$�2+��ĩ<����?�����$� P��J�>Am:�a�50���1��j�I����Iy�	�����<ruC�%���w�99���r�v�@�'�"�'�Y�0�1�$��$��5U��"/\����C�����?�O>����?�ъٯ�?���B$9<IC�л_��Pr%�+�I�\�Iß\�'`�,sw% �i��F��P��$̠|��@�bJ�?A�doD�'�g)m�B�'N�$ْLЙ��F�e�*՚��$13���'�\��fHI��ħ�?���ö���`rDE�k�5�\0bǧE쓗?)C�ߔ�?����T?�%y����h:�>e!G��>���rA���ʟ��I�?���u�]�Bm]�MIq)G-� �4�?��Lݸ�Q��l�S�q$�M�LմN����B��M|�o������4�?���?���OӉ'��m
�j"���/�#���6Ɂij�7��������	�9�v�ݍ{�04q�f�ZP� RG�i�b�'JR'��DnO����O��;��M�fg�	�i�^]0c�ЊFJ0����ܟ�ۆa�A�T�I$*Z�v�&]��P��M���X�D�,O��O��|�iP�N�T�!�NYe-X��.q2�:q���v/�z~��'#��'��I�V���*�ڶYF*Lywd�$J��m�4+�����O>�d�O��D;�ɹ
�6dy���VT������@�D5@���S����T�	؟��I蟈` F�C��O+y�F�q)�e��}��'Wݦ��'��|"�'��E`
6�=\ Z��f
ܞ]L���&��$n����|�I�� �'����3�~��\ ؐ0r`�3N�x���9*k0u�s�i'RW�T��ܟ��I3D��Iן��I�� ��!z1�i�`N��]X��M#���?�(Od)���H��'{��OB�A�*iT���OA�a�	�%�>A��?���V����9O��ӵ9{,9߻D��}�%W�6M�<��-W����'r�'��d�>�;jP&xC�L�}�d�!�"^}��o�ğ���u���	|�Il�'G�������E�,�AR�2g��n|Az#�4�?���?���g��dyR��!I�P��$fʜрӫC�xl7m�%���9��3�SП�Bd�v����_�a��iB���MK��?��i池�_���'�r�O��	Q���
�����HA�Sp�"&�i'�'ϸ��S�T�'�2�' 
%�B��]i!�/t:H�b�
b���D��g��i�'���ڟ�'�Zc������w�H���47ڒ�!�O��h>O���?����� �e	$��+u7���iT%!� !��<��Ify�'j�	��	П�ap��-f:���ڗHrƜ���
e5��	Yy��'��'e��'϶�1�ҟ�y�wi��*�&�X���7-���E�i�r�'���|b�'���\��ݴ���3�i�P�z���&H{8��'�R�'U�Y���/0����O����	�Tt"1�Ye$��`��@��?����'��x�&�$]�d_�����Dku8L�t���Ax�F�'�r�'�"��l���'��'�����(Ⱥ��W����@
���(��Ob���OҬ
�(a1O��;�Є���LaK:tH��	�Q�6-�<ɤ�*XO�f�'���'����>��u�f̩PhÑ(p���皍m�To�̟h�I�nט�ԟ�����0�}
���� �ڜ w��>r��8AU�y�`��/�M���?I��:rR�X�'7�������@z ���
%eh|�tӢ�<Ov���<y����'�4f녺K�H�G���r�2���&u���d�O��_v.��'K�I���;��Qi��XA�ă���rc�4n����'�x�����)�O����O�Q��#Ρ?WVx*�
4r�Lh�&JEަ���a򐠚�OD��?�-OF��Ƅ	�n]�Mu>�B���5hXpek4V���oy�\�	���	ß���uy����^��d33(��Z�~p15A
>��%g�>�.O��$�<���?��"8L��[2.j���Պa_��٥�L�<�OB�8 F�
I̠��ooj	;����BlV�:��x�	�;�U���+9|(��O�-���"]͂��U���������K
K��q��n��@4��l��k7T��l0�.���H�_�(J�+ؓH��:��י��	�D��j��m)NQ�5ŔMx3M�?7|�e-׍t�<���ڃ9�<�Q����4��� � 8�4�
#"�].���SJ�X2�P"�j��1N2i@��� �PY&�E:��{�N;dM'�"��A�E��p���m�X`R�'N��q��
����W �j�r�X�.�� `ts�L�-%Z3�� �z}Y��>����n�I˱D^^�D����T	*�CC�~2��ƚE�P��Q�Ӷ.��p�t�D��m}R�'4�>��>	|k�$�J:�"�F��=��C�	�]t��Af�	�����R�r�h��$p�'�V@��`:�6�X;�*��ei�>���?I�BS�>��pQ��?����?ͻ �����H�} e��ѿ�@z��:X�F����&P�g��83� ��Aj�7HC<Ds$̀v�1��.����:���|�� �~�%fX3=�BH��Z8}�����O�	=ړR���vbZ�<��	tEW:7?���ȓ*K�Ĳ2��4Rc�NQ�;����'��#=�On�ɶ�*�zs�۬2�Q.SZ�Y!w�*Q���Iڟ ��џ�z_w���' ��b��C[�[��Q'�]"{6|�8��K%JQxe�׏݄A,��ā>p�D���C�-��
�cD� XJ�g�{��t� K�24W���{}֍Is�]6�V�8�]�=`(���'�r�	}���Y��bT?d�5�WN	'�8�ȓ�� ��=)�b��ë��h���<)4T�Ԕ'd�x�HhӮ���O�<��t_����AN��Da�`%�O��d�����O��B0�m�_�"6	BW�n�4�;��B����$T�'�lc������8Y:��1��9�E?O 0�4�'�rT��" ��oDP�`��,�k��~���	ş��?E��a�[�*I� \1�qrwJE�xR�~Ӣ,h��_6�@x�$��*%�AJQ9O��?T��Q�|�IO�4gŷJA�(қo�@�DH�V0��I��I���'P$ȖEV�D��٦� [���T>��OH�@!���",U���T[R�r��H�b�í��}s��F��/�Myt#Q A�"h{%�����ɛA�P��O��}���X��p��ؕ��]�%�O�S��d�ȓ@
T��"F�����oֺ8� 0����HO�<S��&0��� �<8�@�Ӧ��I�|��.~�yR�
����	ğl�i��C�LX�
B�K'` �]dFc`7>�\c2�	 Mk���I(����|&��1"g�=D"���Q@�.V�de�O		>I��� l��Z�[?{�X�>�O�)H�� �`��oǬ?�"�#�?�	�=�*���|��ī9�,`�Z�q&��`�`���y"���e��	@%�,�9�V�������8�t��cM�Y�JVW��\�^7Af��$�O��D�O��dB޺S���?Q�O�������=2�:i��j'	@9���O}�|��Щ:[˸�3�}Ѵ���I��m�L���X�*���qB�X����p�M	�$E�q�A�@A�p�'%��6�"ؘ���-%�����m�e���$!�O�!�X+y�6DhCJ������"OF�Z�ĵd���(ЭQ������R�*�PÓ�i���'���e^2~^����.�#0d�����'NbڑM���'<�	*O�j7M<��V|"<��'�1a��}p"j �_i�x���Y��O�A�W�Ǎ^��a����F���"u�'6x�����?���?iwkʱUD�p@�,��I["�W����Ob�"|z��T9T�q���A�p��B�n<�`�i:p���F�a����Д
�-c�'��+kP�ش�?�����[ �`�$�#D��+��F4� @�O�&ky����ONX:��O�b��g~�r!���c �j(f�������	�C��"<�*tnW��@* ���dF(��'�S��@.c������~ԉxu��b��T���ɯB!�$.l�~8C�^�b #̘6.axd?ғ��%��ףiʐy
0ş�j�YгiX2�'1bA"-x�H��'��'�w�J���âS��a#�
c�-��
U��yV�en`��%"&X��ǝ���'Tr��ϓ8?�`��(S65[������5��yr$���?�}&���1B�w�LE@v�#	�hX�0�<D��&U?,V	Ѓ�@�^�[#�4?���i>}$�T���@�r�P���o8$s��/.k0� �@����I柼���u��'�?�6��B��8D�����՜y �xk㄁TN4���'�O���r�*s�p��'.ؕ����QcL$�'�pA̡�A'QTX��hF)б�B��&?]8'��u�
��,�O�iSPOB��15��	�����'w�'B4�BO��n����l��]~���yB�p���OꄹaJFA���'��P��DO+>���I�,Ȏe<��3P�'_2��D��'��)�3�r�K��ĆMYNz��`�p� � ��m�(�	AD4N�jP��'p�7�Y�&�x��Rk%kV�� ��������wB����#$�'C����?�)O^���C�;�� ����m�|[6��O����68ƅ;l�*)��qr��+H��G{�O�7�D�#��Уu�ݵv#V(2��"0N��<�f�Ʈ}@�&�'	�]>u�1�ʟxX��=5�"caD��ȩk��ğX���w����z�S��Oڐy�%])*OpAi���[~�)3�>��ȍN���O�� R/[���eNoo�٫N� �j�ON��O��� �ӓ��1���&�h���p�c�X��ex�hK�Ď�Y�,Hu,�}����<O�1Ez"Iӧ]���Fcý+rp�w��^�66��O��D�O.�K�4�����O$���O�N�y����˹e9�L�*�2$��@����v�h��4
�uSF"�F�g�I�0 ���B���f��s-9`?�: �=D-���i9p�l�h�g�I4n'���E,��Oǘ��UhV�i���<�hV̟�>�OȜ�Ѩ�+q�bU@�d�<|��t"Olp� ��dG$�K'Cˌ�F�w���Y����~?^� �l\ �N,�f�+sH��A��Ň 8�a������ݟ�^wS�'���]�!"LQ�Cn1:��l�r.���aO�퉐��M��� Y�)��(���!�d�M�N��B���jS�,+ᡎa��y�'���-��C�Y��suB�y�o0E�����ѡ8p :V�[���'ǎc���!�O0�Ms��?--4*\[R&�:;&�)�a�A"�����,��\����|b���+{����b�ȹ6sb�HѤW��#G�Xr���"���9 l��d�"T-+�4q	h���F��<.��hi*9��@�-ڕ=u�m@�%5OF���'@�'*IC��	@�bSń*tq���'>,+тL61�kbLǰ�|��'��7�+|<�,�cݤ-�aj�"��u�1OV4�t��ʦQ�I˟h�OQTp T�'L8�S��l3�Q�w�ݪ�����'�2"�.MCb�T>�9iX���̏�2����"oF 7zrȥO8Q��)���Q(�)�N�=E����#�_#.t�'�����Θ��O�.��cZ	��Ҷ,͡q$�'�Ƶ��nI?1R�%�Q�@|��A
�
����KUA�k��X���٘/ΈtK���?�MS��?��e�q˖B��?����?��Ӽb�Y�S��[f匤y2 @Ǐ)��'>� ϓi� �ӶT�܉`�	�Tm�=��	^x������+�f���d�p��m:S �G�s��}�)�3����c=�(��/�(�  �ߥZ!�$8k��DA+ׇ)�D�ؒnY&2
���HO>qj��À;�� ƃ��a���^.Y|x��Ο|�	Ο4��q�$�'X��C�/\R@�e��!1��Ų�A�:u�x�Ɇ�)�O�&h�#!��3Sh[\:�T;7��i�<��r�ݡ�l���'�^}!��!��=bh��3� ��	1�?�2�id7��Oʓ�?ы� ,�0���QU<�a�Z��Oʣ=�O۾�P�F]�e���_�T8�����|�i،T�7��<���	�A���O��7i����0+T��͘w�R��z�D�Or@��	�O6���O���C�K�C��O���0䘘t)f88)�K~\h"s�'&9���V,sal98������'ǊPv9P�C6j�d��Q8�D�� �O���W˦Q�I.aE�l���Y�F6��En��_�<��'����SJ�����Y8?T�x��]�-�T����O$�n�:" d�Z�L�4��`A��G�j8ڴ��d'@,8n������b�D�R�[�t�k�oD
0�l3iͳZ(��'�� 9R�'�1O�3?FթZBR�g雁E�Z}�CmZg�d��2���?59�� �
�h4��:w��I3n/}�Ĺ�?a���?�����OT�qi�OV�Nt:)H���.(,�ˈy2�';�y�h��\1�^΢�E�՛�J��ቆ�HO��I<%[��ht�+�����Z�e����@���I�h�)� �՟�����8�����r5L�a��F!� ,L���k���)D�0�)�l�g�	�Y��M�톫"��5(�*yV=!N>�B̒Cv��>�O����lԍS���j_���'7�����,O<��=��F�N�uŶ�ʴ-�-aTC�W+jq�Kϲ^V�����������?I�'���c���>( J��$�[$K6dr�@�G����'��'�x�	�I��<���D�� �奇;T.�Hk�b��1��XQɓ�e~���ũ@A�3 m�/'� ���S�]���1�C�7캵SF��f��X��h��p��"u�N�HH�a�D#<a3�7� �����W�t�ʳ���z�D��Dg�O��DW릱��iy��'�����Q<�Y�'J4 @ׇ��8�)
��H�h��h+�'w��#]�,�&��_��H�y��;�,X0ņb�P�dTL}"[>�2��)�M����?)$+��.�n1���Lui��c��H��?i�P851���?i�.춵aS�i��'⢱�ק���ڤK#*Еm]J�zǓO��4B�� �P-|���O��X&
�%� \X���jʌ-'�'�Z������f)pӚ�DL�!zh�U���s$3��!>�ʓ�?����4�'+��ED�P�j�Ȳ�Yޮ��	�'Ԯ68i48�E B9���qs*�	520�o�[y"�]�{eNБ!�'ARS>!(&HF� z��� 6�
�F;�\����^㟰�	%I�)�,ؤO8����0t|૭���'I!f%�$|1���KJ���O��rRL�3B�A�2o
5v���B�(��Md��gdK6V�����<V�'����l#���'w����'>�z1�u��if�H�eت��'���'p��'&� @��ҽ�Vg=R��a�=O��FzR��%UН��&�3o�@���C�p�z6��OR���O�=��I�SJ��d�O�D�O��;|Ϟea�Z�1e�P	�� �l%�s�yrB�_�ʏ�D��<
J\R��	6&��g��.!�Zc���J�& �q��'*�Xj��ÎG�*�
�!�ͅ�:G��'��aZ�:�)�<1��7�;�)�,-@bJS��b
�'�U��.��}��Y ��2��p�O$�GzB�AZ?�*O�4ш�D6��"��Ҽ��J�ݢ9F��O����Od�$�պ����?)���̒B#(Ť%��B5)'*pC�'���<��+p�1PÌ�N
�0��R�~��A�4S�8{���g��uR/�E���b�=(�l�cڂ5ڊ,�Lɭj�,�$�O�	lџ0�'���D���|�tjW�L�n	ī'd��*�ODyХ/�z5���������6,4��^��j�l�Ky"�M�1�םퟬ�ɶ;V�2���>lg8��*T�n�����	������|�b&����z�*]^�Ԥ�4J�d����Rr �C�#*h�	��6\�����؁o�b$�F�����Q�I)	,4�P���]p�4���:O ���'���'��ҳj�Ё�A`DR�&�8��T5L��ß �?E���O�LM#s�_�G���-�xR/p������()��1�᪖�Fk�s<O,�R�Ցb�i��'��S:/W���	�@��� W8E��!_R�
T�I؟��wgިB:v=��)ML~*�@ʧ3tހ����PYb&k��(�bQ�O~����*V>�ŢA���r�"}�U��� �|LXC�$]���2g�Jl�Ĉ;H�"�'��'o�Dly�bI���Tԡ��o������O&��8B�$CG�U�}�h�j`ߦ�ax��&ғiq�Qp��Un(�%"3�F�-@�\�'V�}R,]	g�2,�WF]�/�ثMN�y�m�dL�f�� 8Ā	ǎ_�yBKBJ��%�3���[���3�C0�yb��}&��zO��|�d��R��y��Ғ^�(��"��� ����y �)>�I�5-Cy�qF�=�y2���]��uB�oW�Nf~������y�d�b��ҝK�r8��k�<�e��(A�ਇ�!� i2F^u�<IT��L��u�R'w���cǞu�<�@�N�ꕁ��H:���P�Yi�<��  B���9tA��J�~�<i��ڪg|�ӆ�����a�x�<�SA=w ���s�߁~��s k�<�udJ�Gt��1SA��P�$��r�M�<1!]�&����`J_	"`�-
��F�<iP�ӟh6��.���x���@�<�c��	��M����%0�(QI�o�F�<qKοyDUi�-آ-8�@���w�<��պA�H`�r!�a<]����r�<Y"��4V�} �L��8�*ݠF�X�<�"G 0{+�P�$%B�Z�������N�<)D=Q�\�Go�
{N  K��u�<�"�\�q$J�䔂^՜�Z�L�<Qp��=�^��d�N����W��M�<iGN�9=���(T�0L���I�<� N��E!A�6T��/Ir�y�"O�lÇ�D&�xi�Q�ǙX�T	�"O"}�����r�D$�J�'�x� 7-�j:9�'>�����O�Ϙ'*�@4�U�3<~��e�M�/L=Q��g�T��@ҊH�.�rբ�7��"��1'g$����zxs�&[ʠq.�6/m�t86�Ś#��G~R��0a�xk��Ñy����ן~ ��؆�H��L�h��
�"O�8�B瓔M�r ��cI�(1N�!1�O�m���_��E�q��Y�]G��%P%��f��ՎlI�*1�yb���"�`���G�x�<�kT��".�Hh�8`��S��u�-�媘�&�p�э���Lyp�:�㝑2 ƀ��v�azr�Ɍ� #��Q���dȥ��4���� ��u`�K1�V:�L�5}�RiKU�'�2]H&�_i"�	5n ��x���y�n��hỗ/҇`j�*Z�caɴ��?q�$�K%<؉P]�R�d�I�H�)�y2�6�� s�F�.�S2/V	2{ � í2�h2�.B e{r�b7�-vT�O�r�`�w��Lan�k����F�.�
�'�20�I[=l��hjw
��'D �X#!;��r��r/�{D��U�"�7IZ?h��b�����M�����ewV�#��0LO�UI@��?��税� hP�� � "Ϣt�փۖH�.��s�0j��!�$Z�*��l�דT����&hA��"F�ǡ|^���<aƆƣxV��i������`������عBԸ��u�Й��=JF/T)��ywA�U�<g�>�ژaӠl�H,�5xF`����+R���0��"zAo�~��O�����wFp���Ev�M����O�DY0
�'b��B�έn�`Xاj�6+�U�J�>h����� ��"Fh�D-D%/j�ϯj�px�=�qB�{D��ՂȈl��9z!kAO���*�dE4`���5���w��M�@O�k�\([R0�43Kє!�t�pǕ�eՀP��'��l��j� ^�f��42 (H�y��0:�I�x#��
䩙�ֺ�J'�����;�x4���{����Φ=�C�I��l��vy��eOB�D��S$�A?���R0 ��M�f9�#2�Z�8	����'b*����n����(�%ޜ�s���t���+9܌��AK�?���|皕h�q8���!��1;�`<���X�R4�Qc�8b���38o��*A15����'��{���3M�8��@�[nP1�%�G ��'�4�H�@b��7�F�~�Ad�Z	���D�>zm����F[���k���-D��2O���q ���:!�I�������ɩӮ���MоYW�tsm�~M
����K�(�͛u�]'qW�i�Ӭ��_S����E��9�qOz�i��E�#�:��`�X�B\J`�Ǧ��F�^;ƦӉ�p>arfԽl!��p�� w5ԈpOf�F���*��L��,2QO%�3������m�Nĳ{����ҡ 3>��2|Os`#�<�:M�FT�&o�X� ���J
�"�H�1�ax�Κ$ ŜUP�� �R��� "A�w�r���?$�h�k�m�&�$�G��� ��Q	(�6�b�D�d�P(J$�P.U����]��@�g�H�Oq:hiv�<)m�b->�뤭�= j5�1OD�'��qħ^6�xH��U\|���]Ct�E��')X����^�<���s��NE��yH�y2�D�NUPa��Ό0N�& �wJsN��P6Om�	��	;&���! `��kd:)������aF?F���®��MS6j�ߺ�O*C����Zc}ܰ��eB�w��,#t�9&p>�;�'��c ƵG
XA�AY�T�T���b���~b֕�X@�II�|��.q�|��ʒ�r�����H2uMVAS�y��h{e,��f+�(	�#� xAcЅO����!;Q�8� tY���"�  4lD\�@��x@aԍ_���'(�P�@D)I��PX��3��y��sB���R(E�D��	���'����,��:Q���v�ɐ^(ljSg��~M�9�M�/'�{"oK%,?�I��ݗQ�r��FOY<9r�U��+�@�|��9��'#`䔧��c�� DY�!�#��c���C(<�T���sR��p�aK�&��EЅ˚*2�#<QA^����-A3_"��a���0PuF�t� �ƍ�4�U���%�)��.$���t�Z,(h�-C3EQF� x�e*$ @�H��zt\ݲ��!}���}u蹸a��#���@��$��'dTX�]�h��u�*[�1F#�O���v%E�"�b�0B`��J+8���'_Bdi򘟼*Ճ��(8�Hr��W��D٘#BӋ�X���7�|���V�my@�f��/#Dq�"��-aj�ے��!F�Y�6�'���0��OqP�Z挍++TQښ�y��GeB��@V�ytt�ڷ�V�*�!��7�l=wl�j��pY�O�7Chh(5�Ǳ5O6X�Rf�Qt4�9����V��t�'m�q[�G�w�hi*�O�B$�O�u��1�C�T�U����I������P?'�h�d�'IH �ELh��E
穑���g[R�T��N柨QЭ�Ey�1�M<�=�Rd����v�ԻJv�]�6��U~"��3���DeZ	k܊�0��
��M#���=5��Z�n�eS�������G�ŚO����6�M!�zx�D��==�a|�J�e���#ŗ�
���r�.-�(R2�^�|�|��ϓ�y� U��Q 0�
�H1"����HQOT��Z�9a�4hcZl�Z��v��H��2�'�5jkJ5,Z��r��`!�Rb^8^#2��[��Г��2U(f�Er�ؘ
�n��H_:bJT��1�����c$ұ7|z��邟h�(rT��	}���X��E��M��jN�]�#���Dy2m3<�p!fiB�����õ�����tr���t��4�2�� ���}���K�i�J�&�VX�$3oo���i�&*$m���:<8���r�@��b	�shJ�G��`�SFq�O�����>H����D�z⚯o�8�����������t�.}���V�yv=�=��F�^�v<�0OlPK���7K����8�% �E3���Pk��WZҠ�%��U�'D���NS�=�^hK��x��$=6��e���;"~Ͳ��W�]˲�a'�Mv?�`��?���|�<�Q���h��)�Dٳ\ff�tn�L���'9�d�l�3}��3�vU+�K�no��	F�D�D�Z�@�dG�?$����M~���]�BVz�f< \���R��69��7�:���<��H��v�� ���Tw?�ӥ`�u@ᢕ,1[hё���M2�$3��,Od���H��ܸ'�ȅ��!z98�C�MP<�ez�)H�H�����tX��g)���?ex�w�2%!'g�X���s�P;4x�J�O�L��������T�ߩJ��&䇡Hr���у|?ϐa�E����u��Q��Z�;yx�ܪ1n׉��@��a;�ɩWF�A���|2f�|�rcY�[�t����Cj��ap��f���DǏ�x�;�N=lO�N˰gf����e
�����$솃��yJ>� 䖣B'�d�I;hۦ�)u"�Ο�'o4����(X'E�����E��R J3�	697�^h7�� �(���o��%rV��흋P�.��gU�yz�Y&oE,\޸
�ү>�V��S��y�h�5~��Qcs�>+
���j ^vXᓄ6�n�㷪�;)(F ���e�D3y�,0b�ݳcMp���#
�?����"c�<9���<��ם�SMў�9���&��01���<)��y�@�q�{�虼�?i6f3���Ӽ#BG�.qK�u�ӎ˿)��$㊜b�D��,J��hO���gZy��� c=��Ѹ� �C��,�ݖN�����'F1x��ڲ�l�O�1`��#��*H*6�n	d"V��J�cE�U2�؀У	Rh�r ؁ҧB� �b+4�D^dc��J~��}$pB��_\��0��"��$�+IB&]s�r��"�T?	��� l�UZ 9O�չ"L�IB��5l��`�H�kB�p�  DzhQ��f�"r�O�-�ED��Q;�b\�r�8�(Ѓ��e��?Y��jL�28�*ԋ�B����s& hT���e� Dvr<�5��	=o��T�I���yc��!Q��Z�`P<�B�)E�?8��(���e�"=��8�Ȅ�W�.?��nѰU{�M�UDޝ~�̍pbϓ�2�'����ۦ�9�iʂ!+����$'h��kנ�*c*��#)�	�j�*��+��1jMp��Y�6ZA궦#?A�i\�DT0ūҀ���4F�k~�V�qODUrA�âF����0N�4�z���V�!r��Q#*���iX����ja�G�4��c�8{���?˟����C[}�< qd�R�#O&�p��|b�B�c�&�r�+����Dӣ�2��'�Ƥ�!
D��Fx��֗/x��� e\
��'��>�I�՘Ł��E� d� ۥb���xT�I<Z\u
D���qO�Ӑq�2qϻ���$+w쉷M
�F�h�����O���{��}��6b>(4��E�YfH�ӌ��y�1OH�ׄ��9�a!�R��t8����\oA,}��jӕ2�^(��΅�Q��y�bõrS^)��ƕ�u���,G� ��EpjU�gLؽ#/�$U�rU��O$'!V�{�b��IP���?���`	�x�D�$,h4Li'Kݡ^<��螧T�I��FӴ62����$ˍEQ �p��F�7��t�al�+���Z�DWAj��>�Ą���&�u�'bJĊG�N9-�\����0xj�#�T�8���&�U)/�.��=�O��� P?��YK���-6�䋃M��O�^�"a���d���`w�L�xXy���Rf���O��PS�k�*\_Ȳ� G#(����/�I-c�����u8f���M�+�rc�<�E��l@&�pB���q�z4 b`ΓQ��l�<ӣW#`����9#P�;��F�`��(��Oߒĭ�9���+R�n�
�A�"*z�,K 薼S~�xR#��>dV�Y�GQ�}��(���0d(���5����/�)�'(rpd 'jV*�=i��Ζ&�:e�㉊��e��zۚ��	�O�8�(�Ν���Y/;�ڙ;qI^����e�̉]����{*�j�1s�b�����]4��p�@��F�\pȷ�!}�=x���gQ#�޹E��F6�l�ÅD�*=�މB��zi1OވF��:��aa��V�t��w�ĜN� J3,C�Pɦ��	F�y���� ��tC�$�'���A(��dJ"ɔx,�h��bX��E([
R*���gy&�B.��z�Z���(U�"��ys��'��` o:_�1�I�)���GS2Bx��a���1S�@�Ƃ��4$!����y2AK�v�V�9$��+E]X3W i�铗�' F�{���+�X1S
6�y�ρ�`IV�+C�����97)�UV�$e��6��H�'g��]*i$,�ƅ��1*�kW:g�d�DàjT�A���F:v�qRGF�?-�&��'j�$�3u"���tt "��|$���#����%EW'��	'�?� ���J��� 䲀O�H]�͸v!�p*QOp$L��Mʬ+��I��A��� O�T�S+r2"���	G,	���sF�ޝ!���I�=pŐ� X'$�S�?Kd�)žith�R7�+!q�9Qt�8)F}"G�5CN�/�3E��郗j���Ϙ'αؑJC�;J�1U�ì' ưX�O�Aa$�Ƨ�@�c5��;3BI�=Y���]qΡC��l]&%�,�v���Z���@��mBH"qF}R��yg%�B$���kX�6���&)	ֲ�"4AC;��c�l�T���!��-�'D�$�-{b���dS��|�y����#>�aG�Au�m�j#�S�u�������Ov�p ��ϔ�'��H"��(+�f����|�uH�~]�"R��<���<���5>�"d{��3}��I�<>c��c��)YH�k#ɉ\��ϡvn�{����	Ь����-��鉠!�4��g�L��IS��<)��
r����b�#۬e*B"�b�������Ğ�,��٢�	�4{��CvW!�D<M����p �+x��T��F!�$I8|ڄ�[=&�|`:�%R9K=!�d^�%M@lkW�A&L�y@1CL�E�!�č�3�֕�K[�0�+�G� %%!�H�F-hD���y�8bU�B5);!�dI/lX��X��ıyjt xI �!�D͊њ�ҧ%�sc���! �!��
 �Iz�MN����i���MY!�0sY �ф� �z�@�b�ƞd7!��d��X�(�!U%���R�Bg�!���0����� �.\""�ԁr��C䉠>���3%�W�F���e�?VFC��(_ƹҧ���v�t�#Q�˧��B�ɯH�zY�'�ץFVJ�b֝��B�I2jݦ5!pJ	%&I�H��һ��B�@�NVR�@ L0㣞$��=��'u��M�;P�'fG;�H�'r�k���|�1	�Z�2�yr����$y4L��afe���>�y�ϚWS��7#& �:��1�yo�$:�R|�Z-!� ����yN?i�<��(\�D�nH�f(X�y�'�2��i{`"�9�� �T��yB�͜e�,Y#Ç�$�pq�b��yb(�Q4�Ԉ^��Xly1���y2)�(K�fG���D��s-�y��
�]y\e��!��h��T=�y�`�*j7����l�j��e��y ���Ȩ����^�dA���y���0P4uC#�� VIЃ�D5�yB^�N�F���@�p���iC��y�$��O�L��E�Μc�y�s	�yүD�dļ!�dj��X���S��L�y��=�����|��$�B 	��y�dN/f摸e��:{�q�򭑭�y2DT�,�R蛺)'��� L��y��YR�*�H�"�v8���4�yr��	�F���K�o� Us�̖�y���U�h��O��|�\��R@���y��	�&v����\�r4����Z=�y2I��o(杀��"m�ƙH�چ�y��
�`��q��bܘQ8��	�y�Q��1"O��H�%�����y2(L�X|��JBC9N�����mė�yR"���V���_[��$̎�ybO�eޔ�5j�&(sR���S��y2�Y�R��:BM� �d�Kt���yba�V� �"p�ˬGҰ�j��J��y"�M2B� ��@��iA�H����/�y��Ɉ0����3���54`Q��P#�y�%*��t��Y$��)��͈�y
� D���B�Kz����p�T;r"O�Z&�0-���P鞗o�,��"O }���}��� ��Q����W"O�\�q��(D�����w��E"Oʠ�䯗�� �#7!DV���"O�Y�s�W�Nfh�����>*&"O%����q{��S���$D8h�6"O�ա�����e ʕ8#B`R�"O`���#2)�}k�,v��cA"O$q��*li2�K'lh�\����y�n�2f����%@m�9@�П�y"��d�����$�pTcB ���y�@V�.$xh�Y�s�J����yRH�;��e0!�;3�}C����y�J�'
	Н�!G�@r���D��y��o�ڳ��"1��1��(���y��=qL�c0�_%�>��@$��yr�Ɣ�^�hdȜ#����e�&�y"�/+X,io�p�t��H@��yҫF�9�q�Ҿ~u���	�!�yR�H�g$�C��R�w���dg��y#�?�|L�V���&!9
����yR��	i�tS���6zB���Ǖ��yB` /ZS��)%�ě1�1���4�y��9KIҥ�'��<$5ڽ�����y�� �Ʊ���Ѿs��bDE��yBe֯*0�%Y��\(�u!���y	�*[�֡�D��#N6��9b� �~b�)ڧtZ�`�E�"�Iҵ)��~�P��=9������A�NDf��3M�3�+!%����R�t�8}i���|.=��Ɩ-!�d��� ӃǍSQZ��A�@8!�QPd��P`��S�PKR#n!�D�;B,�LǪG� ���U�!��=��Ȁ�[(������q�!��-�ASbə4������;�!�D�~����u)(�ڤ��a��!�DR�d�̌ "��x��#�b��!��.�N�RH�R�����L��!�$v�i��MH�;�@ȑ�O�	m�!��3d
.��߽|��H�CC�B�!�D�8a����׬�Ш:em�,F�!�D�C#���e ˶c�p 6�[�Z�!�$+f�����3|�G�8
��*�S�OZ|�1��t>��n�D#Fy�
�'�m�T�9S�<��敕D��̳
�'�N h����{-2E���8*c
�'*�`cM��G�zd�G��2&��S
�'݀�c��)D	�	@�2ŀ���$+�r��(�x�9��E�(,(AQ""O:I�3��0�F\��₈{��F"O�˰���c�4��p�v�
 "O�����L|
��1�8X�P�"O�����2A����M;���Ж�M����ú>]�0�U'@�lN���$D���'GR�݂���R�t����'�d3�Sܧl���M�P�,�bΕ�|�XL�ȓah8{�H
k���S"L�����ȓt����p�ƥ��I�D솴e����<�* {�팈��x1�@������X��0iT+�R�:Ԯ�0( .q��	�I֨#<I���]��I6�űM��В5��_�<)�bص#@x�HS/YIx���	UyB<w���Ӟ|��)�Xo|�9�BR5F��Icҩ.I�!�� �� S�[%:͊�2�iĢ1�
�zF�d�z���C�G� Q�N�����D��UG�+D��)�(��ؽ��Y�mz� G�.D�P87��&��M��-�0m�k"c.D��HU�N+b�D�	�Ɨi ढ1m0D�,A�с;~�j6�%4w��f*OZ�i��R鄘sc�0/���t"O�)z���Q#�t�&��&�q��"OTLɆ'7B`~	砗(WiAu"O�yI炙ȩ5b�w$iAG"O��x�h��C�K��A�$*�"OR�R���-&��ka!�!�R���"O�m;j_9�܄����-?�<ĒB"O��g�$
�f���F�-x� ���"OV�c�jD�y���s"����@&"O�DC�l^�/R,!�%"۱8��Qr�"OL���~�T�aR��1,�����'#!��%J�ҹ)U,Y &�hi��	�!��	�AT��l�3	�n����v�!�D��0H(�S�G?,��ۑ��Nz!�77h��ǬR�N�~:�B(�!���$&��+��yY�a�Y�s!��^%X� ��S5x�`p����V!��*A�R���Rp$�x�C8)F!���1#
���`y���(��ךW�dB�I/Q�~���fՈ�¸ʶK�(�NB��0w��$ N��h���ϐ|����hO�>)0Sd_8e>2a
ɺw��Xe@.�O����5�M;y?��h�A�7m��ȓ=��9�?|�2���ȓ|�p)R�f�(\����M���JX�hC:�����ǁQe���x���hp�����k�M�1��Ia̓=9P@��6|�t`ۡL�)z܆�V3R�fж�*@���ӄ	�����ܛ�S�a� �z�J�Mn̔�ȓgV��	�-!��vAۊ���Ol�=�������`�B�5(v#�]�<Y&P�v���	aę=1�Vū��]�<�%$ɫ�də�K���rY{#���<�*���L]�u�ڿTtNȋuIU@�'��?��yz}3G��OފU[�>D��"SD�h'~e)�.^*4�hU��C���F{���_=s��QCu�U:"8��S�[�lN!�$���֐p
H�k��xc�Ӑ$!�$N��=
��@$p1ˤ��z��	h��H����-
��y��n7�!�v"O��rPi�xr,I�l( $�"O�X#2��<����	.0�#"OHM�fՠD� +�B �=�L��"O�6�N�&��;��Y>Ӑ�"O܅i %	{~�C5l�JWPC"OPʗ/Ɯ3'*����M�sT�Љ�"On!c�`��pHx����ZS(�b`"O�#%���d/��m4LJ�H!�"O�MҡI^?���0F���N8�&"O��{4C�h�8��=��"O@,��-��N-�DIH�X���S�"O��b �Ԋ  �T�a�ƹb���N�<I��_,��x���R24���b��K�<1�}hB�#���9/R�Җ�_P�<@��>���@��;I����kQ�<����#�����X�3� �O�<��ʛ�Z�����Ψ��Pw�d�<� m��j�:a>&	ۓ�c!ƍ�"Odth�/3�P��A+܁3
�ػS"O�̒2̅�Jr�Ջ�»2�B��"O&H�A�9%�B��
	w -��"O�HFȏ	 ��8&�Z��A`�	F���i��1� DҲ�!�����	 ]�!�dǋn�Ҁc���8A�~b4a��"O`���+@6�u�cD�ߒ�K��y����^��S@E(!*���'���yb�]�"�d�'+��r�y�Wo��yb�GP��DcQ�4���b�-�y��\e�ᙦ'ŗ~=0�I"���y�΂�z[��Ҁ�$qU �k!E���yB���.�Y��탻j�:]Y���y2č ����rW	�<�A���y�F�\��<xw�ðG!���B��y�R�إS&��Ȑ�A���yr'= :���I[;|�b��yB W0R� Kb.M�)��!�GH�y�JIDz14A��~T�ȃ�y�H�6��}
g)Y)�s�F���yb�Nb�|b@v8`���ylFL��H�V�6��`'�,�y�W��*d(s  [��AW(�y���&���"j���zqB��̞�yr"�
SG`��#��f�8TLI`�<1�oqP��`��ˁR�f�iv	�M�<�``��3}@��f��@��R��M_�<aB�ya7�s`�i"CH�AJ���2��t��;|�[�mޅ>ȓ_��<�3$�5$�p�YL��~��T�ȓ�4d8��T��Ixģӽ��m��\���J��''�r ���:@�hD��JB�$̭ k�4�(ŵzhZ �ȓD��x��b��[�
dC��ȓc���H�p/ZQ�ABY ά�ȓf�,`[�@�6WU& �6͹-|�!�ȓJ���q硆"&δu:&d��V�Đ��F a�Cc�,A�6�`�Δ�$5<�ȓ?�V���n�1�$	�	����C��A9���h�VY���S�+�̤�ȓ'��m(�Nަc�&���A�[�L�����ـ6D*hsj�27�DTK�AZb�<I����6a5�[2��]�,�v�<�U-Ørb�����Y�8 !	�^�<����M!������+S�U�%Z�<i�e3$��ts�A[)��4�HZX�<q�a��J�*p�c��%��:eόi�<Y�ˇ:p�aB�L�!Є���M�j�<��hX��n�*�E�a�ޜ*lD|�<� %�f$jj��__��{��\�<�!�.~ap�k��Vp��j�Y�<1$fU�^I�e���Y�p�v��'DM�<م�O�z��ǀ7n�����E�<P���(ǆi�&��4��1�� �C�<qԥ|����̖!fw���$Rv�<�A��2�x��h�c�����X�<�`��(���P�E1XB�)��c�X�<�i�7�<��a‸{HдeWT�<�E�1�}2��_����V�O�<a�lGt�X�ŕ	+�XT�@/�G�<IaǲT�ȸ���C:ӂ
���E�<��I�OO����%AzX��P~�<��C�ۂ�(�%��#��mIT�{�<� .� �+���he��WKS�X+'"Ox1��KIn ���!*�',B�!qS"O��*�+��g�X��G6++�-b�"O0��⊌$�=�d���iA"Ol[��?VXb���&�$66��2"O�A�mQ�]�)M�m��B �>�!�d=>Z�qN�2~��py�Z?}\!�D�#�`��Rl��B�����C+\P!�d�.qZ0��HE�[�@pj�V�?6!��J�?����&��%�Xy$�L�.*!�$W�∹3A(+��9��ܦ !�$Q
A|��p��&!���c�Ǆ!��֚Q;E.�B����!Y#!�D��K�Ɗ@���@,Y!���0d��ؐ��R�4��xH��U"�!�Ӕߢ�ƅ�Rt�r@E�.-w!�䆹W�@4��e�zM
Up*�`l!�$�~9�������b/\i�j[$yh!��ѹW��X�D. @#�i2iQ#K!�d�@*M�&�P>-��Q�NW 
1!�$��V�X�k�o�<b����ؙ'!�Dϭ����k�$�t�v�	!�d��6�Ѐ I�f��<�iV�%*!�Ċ�S�4YҡŀM�Duا(��R�!��[�8Y�ɖC��i��@0g薵&M!���VONA��8t��P�u爡qC!�$Z1,���@kmb���+5!�Dܗ[�|Uh��#O���/xO!��F�Q�rD�ud˵e� ��ƦFD!��]y")Q�-
�%|h(H�ʈ�3=!�\�Y��h�턮;g>U�Dǐ�!򤚼0x����j]#+�\!�ǙMe!�V�bz�uˀ�¬}8���Gғf5!�DV�\�@lS���"��E$��"�!�D[m��p��ίJ��IjD,R#4�!�D�J{r��LYP��}Q���!��T>)���:����X5!�d��VNQ��K�' $	"j��z�!��K5F`0!m'f�8�wBM'!��A�t`Y��;b`jq�۶�!�D�j��!�'�N�(����!�8Gh̙�l]�p�ʙ1��œ1�!��>AS�8`�:h�blxu�9	�!�$���H��]>'�С҅��!�bݎ��&��(c��E�n!��/^�Y��!��;$+h�!��L���� �	�88	����,�!�D��/H�,�-8zp��JD�o�!�䈕��0�$�B�%��X�S<u�!�ǞIQ�M�����'aD�Pn,|�!��X���f�ݟ+X�چ�џM�!��1�)����BK J�F�c�"OD}+�4$BHCq!�8�h��1"Ol�9f@ϲ��ԩ�@ r��A"O
��'�8|�H����J�h�"OȄ/��80�E�Zv��o0�!��	�(��9"�ӭ$0*�$��O�!�Q�Lxt��fG�s�|"CMY a�!��|{�s�@E�a�vI����p�!򤋞
Ș� Ö(2��t�7�^	�!�[�j�h���	o,V�� ��,:!�dD-� ��J�	 q���r�!���:+TTK�O�Y�`ɰ�M�S�!���|5LHdO�#�&$Y���!�� ����q�ظV	Z�N����t"O��*�&�	7V�T�EW�i "O�=X��� '��E�ӊ�O�Șt"Oօ�U��lf�)5�X9z�d�u"O�h�*��'v��[L�L��Ȁ�"O���c�M� `^@�sDɉm j	iV"O~\)�(M�<a�r�b�`���"OXc�w:�$�c����y�"O,d��`V?1!�	�BP�[T2	%"O�h�dY�dhʡ�� ǹ=���	�'I�%q'E�,���� @A�',h�Q�l�h�"u!�yx�"�'�d�¥ꉴE2iP��`��
�'���bC��$ h:`%���	�'��h�@t�-���V�h��'� �� �_�h!uŖ:#����'i$�P&:����Q9�<��
�'�T����.�PC�!a���
�'g�|����|Xp\�C�Y�J(֠�'A{Ã/mj�Q6�<�� �'ڗ��q��� 8%,R
�'�]`e�]";E\��B9-�"�	�'�$Ԑ!�W���h�--j�,��'x���w�I�XfȁY�+��T�r�'ٺ]�2�]�[f��a �7V �"�'��SȖ�G��t!�POA "�'�da�B��(��Qg�"D���
�'rbx�q�	`ܦ���<���
�'������#�)��)�.1��'
�4��	F1�p8sFG&�K�'��TH��Ư7���s
U<�Z��'�ν!��tt���mY .�L���'54`mX+�����6r�> ��'\��Q��,30L��%ߊl� q�'��!�D�F�Ja�H��W�/5Li��'�l��Y86$<3�D�-/^��	�'�2YK���|���f�s�&H��'#l�$%Ό,�8`FLÇ6ZE��'�>����W�Q������,yJ� ����Op��0§�
�ۣDZ:<|��
Г6�T�'�2�'P���O|�J%�u����"j������.28HC䉺E�R�͗]7�(�GeD�BC�I==Bpiu��	���Q/�	,�(C�	�9&�z�@ӊ͌ �F-��}"C�ɜ=ٺ=bq�Nt��OǴ)��B䉮a��h9R-��R����'��l��?A��iO�B`�c�b]<���"I$E�S�h&��gܓe�F�PT,�P��X���	9�ȓd�m��
�GƠ���5�Ň�8��%�g��#ae� F.�&kyR0�ȓE�>��JU$8���M�O�xT�ȓ�=�fÓ >̱2��rWb��ȓV���8E��G���Y��jJ���T�����؞�i�@\<"EL��?�ӓ^^��5��5�
-q��ȓ\� Ȑq@� x	p���>���ȓ`:���Ț '�\� BJ/M,��bu�pv�Q�3�h��4G�)��(�ȓ���RE�Y�8<3�l�4����>�l���H7�DQ+c-��PӤ��FL���"�Ё�Z���<�'����Э�0@�0h)���)`�C�ɮZ\"�[���7�b�1��[x TC�	�	!	��d�>�)Q�k�tC�)� dX���ȹV$A�q�ʶ�̲�"O�|���YT= ������ʵ"O�`��G�_��)�C�/����f"O2}��j�uN��d��={�4�C"OT�[���`
�[�Ⰼ�Q�^J�<�!�]mAP���WrNS�TE�<��oՕ;
v}(�/�e4�]����|�<�w�.{��L�%��<H���s�d�p�<Y�e�\��9�d��?lV|k���m�<�A��k�z�CF����n,#e �O���,��@>y��%F4?J�=�"��Y�h�"E1D��*穕/L���k1�[13���P5D��P[���0,�4[U�HQa�0z�,C��/n�@X�\�{̼��C�.O�B�I&���(��t]�M!�,5�B䉃|R,�pn��!�Y����ra�C��	9�����O� #�œŮڙ'^⟬�	D>e�`�z��D�Dم=m�\ۀ.1D�4³�R���E�w�ظ�ĲRD$D��I�J��(򖨪��*2D PQl!D�$�u�� eU�2\���
���y"�2v^�Ԡ$��O~5+�J��yR���%v��X�H?2��HEj�2�y�GG�6��qCNY��q�gDP���hOq�lI�!D� U|� ��e���C�"O�dpQ
@p:�X���G+P�-"3"O$"�+�\
DF�0���X�"O�UB��X�R��ɂ�D��]��<��"Ol) �l�)f����������X�"Of�c�J�1'¬�T�Z	
�~� c"OR�����бo�Ќ��Y�xD{��N�R����Bo�L���9��]�!��>Q����Մ��fy섂�KڂZ!��S���:ce�qL�A�j��!�$� V��ѐ�Ί#$:"�7��7!�$�1d��VC��<�����U�Q!� k��``N���
y��־�!�D�g�.Ӏ+�)"�`��A�P+�2�)�'E]0����@�j�,�#�%Q����'2��⥝�'��ccOW+6!X���'U�K7�0=B�$C9����'�TMec�X��9� �95�v�!�'TV ��e�0b���۳d�+.�����'�r,a�"Jb@H�83	Y�z���'|��.@�T��D�c8n��'���+s���W����U�9#&�
�'�z�IQ�Y�r���3���7�zi�'/��W!U�v�PLE꜁k�� A�'`L�HA���>d���#{F�l��'�	2e�g�5�H4��GaU��y̋&/���hH�Bj�Y�����yr��6N�F I��Ǩ?�I�G��?���'J��i�^}�� 5Z���t!\k�<A�D< O�-#Rjͫue^��7D�c�<9�����n�*�o�L���&g�G�<Y3��2[�8�	�5P}NdZ�A�<��B�q��tG(c{"xB  {�<���A���	�,�����%�x�<Q�  �-�$������r�(��q�<����bl�xp���9��4��E�n�<3�Ͽ�J�2��-C�����j�<qe����!׭5jK�bK	f�<�"��;4j���¸iJ��V��V�<�䪙x�Hu��1��ݺ�.T\�<� ��" FP�9�Ty�5l��w�b@ Q"O&��$�� �YzKF�(��)y�"O�|��Oլ��Lq������Q"O�$22�ݭn����� г/D��J"O@಄�>�<pzr��?"��t"!"O.��P�̅#
����ŋ:�R�a�"On�k1c�0hOh�rg�<(��(1"O�� ��V`��&�\��"O���dl0%ۗNu6�iY!"O��h�0o�,+��ӏ ���"O��"�L�#h"��K̠X��YV"O�5c�PE��H{j^/Y�Hc�"O�pxl[u�dhPF�Q�*Ժ�"O|,R���o�4���G�����"O�u�D��-�@-	UB;8h��A"O�`Z�aEK
��D���3�
r���O���2���"!o��5v�1���ص�N���%��i88����N\��m��P��Ș��53\
�����X��!��y�t�D�֛	�B�R��*)q�-��:j8��ƀ�<d�d
�.'zj�l��'���Q�K�2M����j3r��JP�!��h��D�93�oO�d��0�?�-O#~��XK����	t������H�<Ib��Eh�Q����B$4���j�<�צ�y©��͇�l�jۤ�EQ�<�ȃ1B���u*�1��ݪqL�X�<9� \$Ei0�y8�z���V�<�T'W�>
ʵ���B/lI9QGJ~�<�C�U
����A�M�z��$�TO���?���ň�b��cO	�T�A�'KE;�&��"O�i�D��
.������[�]��Ma�"O�$ѵ�̥d����H�A����"O�-���Ȁs�J�s2�89j�"O�!ff��.���EC
Eiy��"OΌ�U#I�_���C�֒C3teA�"OV�J�"�"%��<[Ċз	-�`f"OR8T�6Ÿ�Z ��2�P� "O�Ak��K�|A�D���R�D@!�"Oܜ���܉���Cd�$�g"O�H����(u�\�s�E�vn	��"O��ë]����b��N��Ʌ"O�%-R)%=H%���@Y���;�"O�9�qN)q�9Pˋ'0l�aA"O� �%�2�-Ѕ�];�N�U�|R�'�az"'�,ph�V�����p����yҤ�$/VP�Q��&�|+����y�-�I�d[�E({�YY'�;�yR�J�{������ku6]oJ��y�g�JN���s!ɏ]n��S�	ŵ�y���25V�1�B� \NZeb�-�y�AX�4tZ\p%��#D�ROF�䓥0>	D�7���Qև�c�x|�uJ{�<W!�{j�)v��	o`���'Xs�<��'?i�!�4+�-	P�@ K
{�<Q'�v	��(S�|w�(H�u�<�se��D��p� [������J�<i���:̜D�A@Rlơ��A�<Q C�kG��P�gV=Byv��`�	~�<�4IהX���Ygė6k�B=c��{�<iH��	&����C�6F)�y���t�<���I�X��h��m�R�ҐH!+ Z�<qA�+K��X�Nź��a((�q�<a�Yƒ�w�
�bڌ��Uw�<� ���	\y���z��g�2%��"O0"�d�n	���GMkJ��v"O0Aڂ(f�ɲ��>DёR"OF�DE�6u&hS��R�Ftb)yw"O��c�/Q� ���k,L-
�q�c"O�H���!���Q�/�����"O��X��
�>�*M1ʃ)��S�"O��8 �0/T�J��E7t�Hp7P�,��ɴ]�J�Ƈ4�l�сF!��C�ɉYU��{����pe	c��C�I�O���XbH"AX�W�.6^zC���,��� ڼu9�����̄.��B�I�6��qq`��#d�9`l�,_��B�ɂd���c���OT�����"Y)����g�(*�����ćU�%�h��8D�,ʄm�-�:���KR�2�` ��5D������2S#2l)u+R/]���hp�&D�\���{<q�&!\�?3����$D���hG<얥&�@Y��$D���  �w(��#,V��(6 !D����M��e�`�q@�, ���
?D����?k�l�!6I�-�ހ�/D����)<(Ķ ;�KH�}�l���.D�X&�ٔP����c�)
�����-D�<;a�2բ|�oF�R|xz��*D���U���	yn�H (EBh��b@,D����Q�U$���- �A=�}Jm4D�<Ah�4i�~,��X�Z-���&�O��d�i�B�L��@����R&�	�ȓA��0��N_8]X0�;�C�,��ԄȓNDzz��C58q$�;p�~U��+�Z(є�?$��(��7hm*U�ȓit䉻v���Qx�����X5���ȓ
�]��,B�+��3E��2cؐ�ȓ:RƸ�4o�l�Y��g�� �����I����I�<�6���p��(hf��We�B��I�<��L�$����g���W��l"�E]�<1U�ڔ~c�݁�n�&R��Ѣ.�\�<)�a�V�&0�Ԉ�1o)�I9��m�<�EgK2p/�����2A��!��u�<!�CWd��L��'�08����&�q�<��Z���pht�N$j�b�B	�Ex���'��Pő�:X����gO.Z�^ #�'{Z���ǉ��(������W<$��'X�y�tCD��\Rd�I�b��'���蟶9��T)�([�x���'Le�e�RD�PX�cC�Ԩ�'2�����t�U�GJ��R���'4D I�A�a*�X�%�$E�Ɲ��L�H���KP��z��W!d��݇ȓ�xq�s��ee�ݐW HqX$��:�X�2�#�~$�V���{b�Є��.� �,���S �	�t@��U����h�Ly�mS�h�`�ȓb�EJ�&�U<��=��ȓ	C�=
��I�v�*'�@�����ȓ�Tإ��u�TM�@�d& |�����c��	k����W��z���$��,a�R�n�"m�v��H����Z&�;'W�d��ʔN&M�JЕ'�a~�Iϛw����O?`ϖi�c昚�y�g�3e,à\�OjL��3d�?�yr�Y��lk�A:���q�@��y�-\'A& ��b��2�b\y��E	��d�Oj⟢|� Ɓ��d/y�@�RԤ�-�,*�"ONR@��,4�3��CY{�	�""O��cT!>�arD��Ef��"O� �� ��%���`,�o�����"O����@1NڒD�kg�`�X"O�x���+)V��L.`�\�R�"O���S��2))�	�> � x��D>ړ��D�3xX��ڄt���yA F�Y4!�>桠�
�W��p��ˎf!�d�^n�k�&�?U�j�Т� �.���'�a~��J)C��أ&�� E<�+V؁�yBc�%f�ډ���K�S?40q��ݷ�y�չ&�
<`T���PӞ1걉��yb(@�1���`)]�EL �с�A��hO*��I��~�5	��	������!�d�
8�K0�D�cLa�v���!��8d��L`r��.�^9�p&��!�D��L��֪M�v�.T�4��+]~!�M�!���RQ�Eln���eC�/�!��D��8"�i̝Wax�@�ݸ
n!��[�_�	i��K�riq�8 �Ox�=���
5���v�d�mX�@�VxA "O���2�������b'.�ȷ"O`U{��OB�E�F\��R"Od��¢�8�U�-Q���ʇ"O�-�Հ�%
��d���VF���"OYZw�Ƚ&��#�f�*T��I�"OD�����L�qY���_�D�#"O�s��Q�<��l�7P3`Ⱝ��"Od�q�O1.2-�W�-OB>��G"O�}�g �)����_%z�c�"O愻$i*aP�¡N�!rb��"O"���F��>Jb�rB>8S�la�"Ox�ke���U��p�a��w�8�"O�q�<#VV*�O���y�"ObX�G�E�2x���Ņ-�`a�a"O�V����������o�` �"O�XfNԸa�X5 ��.��Ы�"O���+~,����n�1a����"O�IQ��>K~d�Rc�L��Tz"OX �@�0 H���ޜU�r�C�"O"�xw�C�-˶���6�4%��"O�(S��AD2Re�ٽd��0�"O��A"]�h�� 9��)FBE�"O�!�nS�9	��B���8�my�"O���+�zh�#�oTA H)k&"O�S3���=��������C
2��"Oƭr2�٬'/h�p%�#e�� ��"Op4�@/�-[���A��%Ҝ�
�"O�S�R���a��D�1"OгũW� ��|:��σD��h��"O��Yd�����w��0�.��"Ot�;�Ǉ�1�
̀���?Y����B"O���FA)栰PL�Ny��&"O숑d�!w$��q`X�5[$���"O���U(۹l7�0&m�}<�Ix�"O��rf��,�OKֱ�r"O��p���Lq�3���f5�tXV"O��rc�l۲	r �C�Y2lQ8�"O*�[�o�s YKi�0"2mJ"O\�ȴ�
��@��f��>�#7"O�Z���+e&"I���
����v"O$���n�<1Q�1Q��Xjt"O�*�g��t�f	;�#�<w@@�d"O� Q��g�V�� ��A_�qY�"OF,��Aڲx����g�*+"�x�"O��9惞:��P1��@��^��"O>03f+�*m`B}��Ř��D7� D����W/����H�"?l�I�m"D�4cU��8H5�C�XÚk-D���2녫b.���@N�;W���ɴ�*D�P��E��y;D.�9rFIե(D�����ptj��]��%ʜ�#!�dԺk~ )�@�·dFN�HQAQ=}�!�I����A��92J0ء@I�-�!�d�o���W�ǿo� ʗJ��!�$D2J�*)F����R��!�K�4�f����W�=�f�r�	�!�D	�F)���	�w���8�LD/n�!򄜶�n-�W�G�G��D`r�˱�!��Ly@.���JX'Wm�(�Q�[l!��"�R�dؠQ\��;b�]�!��@j��@�L^!ONH��5�Y�[{!�(	���%4���� {�!�M�F�xQBCމu�n1��x]!�ĔJ��h�#:���#�V'Z1!�dM�kҌ��.L3_��-`�&�#!��?�P��D�c���Q�E &!�1��+Zo�n�бNR�!��>�:1P��Ύ&R��Q�l�-�!�D�(���4��'.�m�Pl��X�!��s�p�D��L)80�Ʀ�!򤛲U*.�"�.u��x���=MX�C�I1.$�أt�@	aw�5cBØ�_��C�Ii|�=j��Ԍ<�!�'"�?�C�I�E����u�x���߲V��C�I�u �yQa&�|�F�����1U�B䉫!_���.qL��Ǉ�dxrB䉊H�
t�E��<e:حkV@�>�lB䉌O�.�
��XS~ĽK���oJ�C�	5rȍx7 P��^]sc�˷Nr�C�-c2J��I�B�2�Y� �&^�tC�I�='b������N�X�Z����q�RC䉙\���&	N�$J]ʑ� &2fC�I}*B1�#�D��x��BU�JjB��
zT��%��[�P��"O�RN�2?��$�%�7mD���"O��s�jֆt�Y�'�E�j��b"O� +�
���`��@
�&hXM:�"Ob�0aL�-���ToT�R*t��"O�A�Ҋy$�`QTI�~b\�w"O2i#���B���(�G�>B�]R�"OJ��_�2�p 4FK�uX���"O�!�P�ZR�=q��R��y�g"O�9��	�t�����!z�l�؆"O�|�s�]�|V�G:N�
��"O�p`�IY�}R鐧�A���$"O��0J�:o��a�GVi���2"O� ��jS�+Č������`��As"O@�Ґ$B7b)�5�0���'���*2�'�'�B��>!a�X�<(�0�Y�1~<2E
�x�<�SF��j��Q��2���#�u�<��	&yx@��(Գ+O����V�<yf
��|�,�EN�/�@!�mSO�<��!K:v��erC���[�x��E��D�<��J�y��R�٩-�\���
@�<�J*wr=P!J�;�v)��~�<Qs�Xf�}�Ɂ;U+<񨇅�y�<� ��+Tc
������m �=���s"O\�8t��9=�ᰱ&�,<&P�k�"O�qq�ZB���AS�=�$"O�5B�,�S�~teɌ*.؄��"O|�����:S�5�v�K���2"Oh4롊@�Lj%H�r��3"Ot9H$�ˤ$δ`
Pi�/L��څ"O�8�'����D�"�K'�( �Q"O����!]7�QÇI�R�"O�)2�Ĝ�^��5���&K
�ٓ"O�бc�����F�_`����"O&��BÏ�g��u�Ȑ�A6%��"O���5��1���皱w����"O^�sCoY�Yz��YUg��HFY�"Oj��f��a�f�a��Q,�!�"OX��"ْ|�� ���*G;ؐ1�"O.9�ǖ�p�ū0��0���"Or)	5-G�tMq�%��G"O.�;5̞J�"���ܠ)i�"OԽSĭ�=<�����X (�6"OT%��d�CV�S�쌸j�= �"O&���Ϙ[1���j��y����"O�|Ҁ�h��*�X���
%"O��Ti���T����[�A t"O>���_T� G,�&��II%"O|�ja䁐j ���ʇ�D�j	y�"O��2F�ֆg�Ȥx2G�0�(�Q"O��AF���_f�ak�*4EJ�!�"O(,�*:&�D��P:
�@X$"Or�+����#M"�8vcAI�zEr"O̴8�O$P������1]��Rw"OtU2i��ZR�D���A}�zD�"O��ҋH�[��:��T�Hqc�"O�qPP��=>ߘ@A��)�N	��"O�t"F'O#w��[E��y��D�3"O���DҤSB�i&.�dv���"O,q�
�*-j񀃂CYj�q��"O���T� `b6�[�yp��ۓ"Ov�"V)��.p�5Z�Ŗa!zb"O`ui#\{&�k㪈�bRR��"O���cDJ�^��#�g�3@E���"O֔[w�=ԁ*cF��WAưK�"O�ЛhW-�e�d>6�D�'"OХYPV"\y��r霅"��B�"O��TeF@�\H���Ão?���""O����@�"9&DrV�3
���&"O�Y�Ӌ�^�P�����&в5rR"Oެ��+�,5V`C4�)�d� �"O4!�M (�j��/P<�8���"O�A	uF	�y�x�2,�"n����q"OR����@�X�	S� ��\��"Ob�zV�I_V��������7"O6�� �$eEV����J�^� "O
��C
�Fp�`�Mӓv�p|y@"O��ѐ@�Y'�Չ��Q�KEr!��"OʙӲcZ49|�T��K6_�%R�"O�țB��*R���pNI[Z|1�"O$J2m=X�4I��qR�T�p"OD��4�ɹ��E�m�6:H�� "Oȩ�6�B��|i���J�2��0"O���"N�ܔ�eB�)HՒ��V"O�9�%N�J���c��9�f}i�"O�$3ǅU�c���p��	/�.g"O�a�G����9HT�#j���&"O� F0�m�i.�h��_T�@aI�"O�tP�C�ď�A�Y�e"O��b�.J�=��+a䛡5qP""O,,R�J��-����0K1��b&"O0� ���Gr=���m��PX�"O� Cs���;pd���Y|@D�#"O.�c�%{�xaS5�� �U��"O�Ē�,�Mv���!$A��"O|D��,i+ !��w�ڨE"O5��$[�+䦑*ԏ$d?���"O���@B$+��Mx��@�A��� "O���H&?�05� �(8+F��"On��D�ǥB'@����:z�H�"OHZ�E�m�HX�H��Q�	��"O�fG9	��9�F�=.���"O�Eu�G,Az
�d�@/��0�"O�E��lQ 4�N"� �`��"O�I�G4B�<��!մ���"Ot�Д/U-$��]Ɂ!�:~$"Ov%: 	M�|�x�!���**�J!p"O�𠲨�q�����7�8 �p"O0HǮN =��b��պ
�v�"OZ%{T,՛5(��rƄ�@k�T��"O� ׏�!z��c%�A>���"O��B�a�(l[t=�ă-(2�Tau"O���� ~ִ;�Y�!�zR"OV�X0%��ab�-9�]8;/����"Oδ�T�5 �jG��HoJͣw"O.0��#u^�dn�"md|�q�"O���u�_�BUR����	|X�0"O�%�n! �u�q�%hV0Ա6"O49S`Ç�	�&��_C4X�"O疴�B��IװZY�a�"O^�S��2-�Xq0��H�=�%"O� �g�X!Ct���65�Zt"O�1g�-�4�� ��.(�"O�x�ĦC���
Jt��%"Ob-�$I�3TJX(p�I���C�"O�D#�# �*Q�G$��t�"O ���	;v@-Pn�����"O���edǣW���Ҍ�E��B�"O�!��ںH�ܳU�'"�m�"O��!"M�p�pykSǮD-�U"O
0�4�{�Bo�L�"O�Q8 ��	0���j�m_�A�b�H"O��X�W� '���$7M(�"O�i�0g�&@#e�ˢV�+"O~Y�0�W��)�U���|��=�A�|"�'g���1�%'��	�ΕMff1�	�':���qȕ&F:����:V�$�k	�'KP�7䆪Ob�4���0R��]��'��SSL��rN0'��K�.�R
�'s�ى5��(s�<��Aqx$�	�'���� �*.p�]rT.�7C�5 �'r���r���@Ϻ�#�/�?���K>�
�c��ܣ�K֎��FEY�[ ��3>��U�ݽ����̀) ���ȓ`��I��1m�j�"B�?u�J��ȓe=�-�$�?*�Mqf�>>��!��p��Y��#<U4���ȱ� ��W���b�<]Ԅi���)U,���Ed���d�Z��yi��ܧ�d �ȓ���Z�@�q?:$�DdԊm��(�ȓ\�" v��c���@�炬r2���S�? "�P�'Y������#Ϛ=��Ī�"O�	��ْ���RF�K�/C��t"O:UZfm��n08�� �v6���s"O�B0�K6�٠�^4"�3�"O�pG�W�Q���+Q���I5��"O�����;"����KׅxX$2�"OȽ�#@әH�N�P��]k�Yk "O�3h�(0hY ���<<�qzV"OB��&n�'�rdQ4aW�h��d"O8�@�-a`�Ж��5-"@|ك"O�ap�H�7���vN� �U+�"OJ�3v�?42�ӊ�\�4��"O��P����a�ԧ	vø�r'"O�}Sw�F�x*�@� T�"w"O������:��1aۀ[R�e�"O��b���8�� ��^)6���"O�(�5��Z]2e�uo[z�@"�"O���u,A+.\������Ig`u1�'���q0�-�.ē�7 ƌ���	3D�(���9?��&�ۜ �e�1�1D��C��F4?�%$�s�1S���	�y�&M�.>�@XA�K�RD�rv�1�y2Ak �u��'\�N��@�B�Ɖ�y��I'B��kH�AT�ٳ!"�y���+@��X�k�&=�h�Cϐ��x¡]7Rp7�N:d
�Ea��&�!�&N�TPVa�� �)ai*`�!�DH7T�݋��X?�48�h��{\!�$D�f��)0P!�?m�<��)9A2!�NBw�#e�׏Bp�xҳ�SF&!��t�J��%kX�4Z֕!)��!�� �{�<�g��::jh���x���1Oj�P��O2v���I�o�0��"Ol�A�&�8{bp(�(,B�)(�"O"t끅��(���bK%K� ��R"O�|#��S![��@Xfg�@�N��"O���D
4(��`�����k��3"Ox�l� �qf#ة	�Ԥ��"OF,b���⎽��"��u
"O��JE��2�@�	ʦhQt"O0�����k9А�ԏK1.���"O>���Ρ�	��OE��m�"OKF�>���3�E�d
��K �L6�yR�Ɋ^^^�K�e�]��%
��y�a��xS�nR�b�3�cK��y�؉�TCw�}�2������y��V8bNw����_ �y­��l,�g�oi *!�L#�y��O�R�����jG�Pjp��ʁ�y�D�t��H6GR6��A�W'�y2�˕~��"���'��ţѥ9�yb
ڼg���X�
�	B�۠Dߎ�y䖌?*p4���ܜ_z��`�!�y�W�9����u'�+4V�� �@�y�%�0� �0ŏ�niq��U�y�4	���)q��H��,rɕ�y2�� ]���aJX�m=�q�v�C��y�՚Kb�|q��/\A�( ����H�<9��`����Ջ]D.�ȓreva��� �h�2���)Ȝ��6����Z6j��f�w`X��ȓ����`#.���Ĝt�8���iVʕ3D�ԖX+1� E��d�ȓn��U@��K� �G�G�����S�? �);s�ىR�FU��h��	%�Qȁ"O���iJ(ZX�$+�ߧf�!R�"OF�Q��z)N�[�k^�s�VQ��"O�Y�#�̋@_��j��
>a��b"OF��@��W�,Cb
Ee�����"OșdF.��<BlS1^�N�t"OܠPs%W:xh�%!�l� ��c�"OR�` �Z
	�H�s�I��r�,�I�"ORՒ ��k#��ZT#�^pbذ�"O �`]���yyС�:j ���"O�1��@	+l�@g��b����"OYW�O�R��yG�� �D�*C"O��� W�JB�����ԕQ���3v"O�p���)X�%J� P .�X��"O
L`�K&J�
ШP/Q'��j "Ox�U��1pT�MX�/W�&�F��"O�-���ݼ4P,�D��mwT8B�"O��ǫ�E� Ô ��[P�X"OH!�vj�36�b ��(ƩkCBI��"Ot�%̘�9s��²g�+jasA"O����^,sZ��� ���d"O���P._�fgi����H��"Otʂ��f��p��S:/e�&"O�-;��[�n�|�C��l��1��"O�8�"#\�m�ހ�oE�v�t���"O`����F�p�C��C����"O�1�j��������\N��)f"O�Y�cK!,=�e���\��}I%"O�`@�_h0`+w��Y����Q"O��ض�؇Q�D�чF�s� ܪu"Ol);&�� /��5)�̞���"O�m�%fL}��Gk�- R��"O��H���i(6	 ��O�<��1w"O�±�\1o��ɸ������`Q"O
F���w ���f�4���s "O2q��#Ǝh��I�4c�Fd�Ҕ"O������nX��9EKW�xӲHJ�"OX�U�Ӹs�b)`
�Ϩ�0P"O昂�e#6e��3cT*_�م"O��3�IF�F�T���Ѝi<|d�%"O��� ���U��4��"Q"
#P"O��F�c�����f�B�X�"O�-9��Q-aFH��l�J�:$ g"O�l����HHBv�օK֌�05"OE�����h���Sv��j�\̨�"O�Z���4�fu��/��\c�"OTU P�'������ Z�6x�t"O�9��9+���ňBKL}*�"OⰂ��+�1�3:�3�'���EF����,�P�(>�<��'�u:W�ȏmc�Р)X�;^4�[�'�F�SA��S�)s�!�=5��ɚ	�'xj�A�^�h�u�;+�4��	�'&�����+�$�H&e�>L���"�'ʄ�d�Դm�Xha�LB�Iun�x�'����K�~=�Y���A+^)�	�'�R�!Pj��5�ޘ*���:.�J���'+��o�Q�[�|TKa��U��'/���!�E�!�ry�'�Dd���'"��a�L�Vic�/� ,�|�
�'�.�T�UnUr����9�	�'�̫� R�r}��uGHuC	�'����d^�F̩��I/g'�ث�'���B�+82��X�)��Y�@�8��� �|�+JT}����٠m�င"OH�X�F�9�vMk��Ro�x�`"ON0	Ł�� ^��#DB|�|��"O֡����@���C+�:�Ӥ"O���c̥E�Z�׆Y'."O�`!��h]���2�\#"���V"O�ـ&/,I�M���,X*��a"O8�f�ɖ5�r9ZE	J+ބ��"O����0��gƟ<;����B"O>��. �ri"0����h��"O�9 ,��'���"c��8؈��D"O<�C���% �D��s���,�$�`�"O��KA��c���QE"�=	P��"O�Yr�oE��s!�J�
Yiu"Oy���X)oj� �7!�mި�Q"O��y�J�E��F"�o;�98f"OjX��f��U��k�斋 ��	�"O�����
c��J�.p8�"O�@CE�Q���@5�Q'89#$"O�9�u�V�+6�Xۥe�?i�!)"O����l��T����ì7�����"O�H�$I���y;&�����s"O���ă5�֘"@���v�r"Oށ�d.]�x=�D���!7��z�"O�l�ԗ.�2ԑV+��>�X@�@"O��X�*N-;3�k kB���:b"O����a?F�����D\Q�"O0���3uO,���.�Eh�"OT�5"�4&�dL�6G�w�Y��"OI�+\�ѷ ݣ0�
�i"O��3iD��IpT�N`n� jt"O�x%��[����Tm�.Y�"�"O�y�$�J3�T��NwT�i�"O4ɠ����LL�	V�*fj8I9�"O����xӨ�YCG>��� �	1D���g�Q�as�U2C�!_���"��<D���"�G�/y"�9ϕ=�t��ą5D�iF�6yjĳC�)Z�r�j4D��B�A��J�!I"K��E�α�4D�@��`A0I���`��Fm��%�d<D� � J߮*�ȸc�����i��9D��:�nC�~m��w��71oؑ�b7D��A�4��1F�Bs�U:sG3D�P�4mٻcì$�2'U�d��jq4D�4ɡ��)}�B�f�my��xw�0D�@���? ��\��E�'*p@ Hg�4D����BB��^�a1*A�B�>�2â%D�
G�ݫs�N��_9�8�K�o1D�8�p��zY�T�^)��Đ��-D��#��ӷ3�4���!��p�s�+D�D;�ʷ7͌My�΃-?h�,/D�hxv��<}P�ܩ�L9� �kD�,D�Љ�b��I�Ƙ�PF����U�D D����oU�)�T[�DI�E��UR��(D�`�¡H_�Xz�b�2p�\�J��<D�@Q2b�'��q)AJ��~  ��j;D�$���'.��1�u"��F �1%/8D�8[�
\f��ؔ B''��ca�5D��!�ʍ')�6\��!�N�Jp��I/D�TI��a��iP�D��>�:��(D�x�ꈿJ̀J�<Sg�X'�$D���an�)#��fG8.=*�s�"#D�Ђ�\q��蕦32�&��6D���	M�j#BmЦ��}_^���(D�� ��Y�A#n������GP8�a"O�)bQ�E01���j�CN~��Q"O%ꇋQ68�^̉�a^5i�� �"O���W�he�B�P	o��ܹB"O�5Sq��9R���H%����<D� +��L��t��ѧp�P��<D��s4sV]��O]0*�����&7D�`�1��1BN\�G\)&����J*D��8eFM<-ab-+�NZ�2�d!�)D��ūW�^�eGbR�l\,�;1�&D���c�	f (Q�5"�_j��� D���b ��&���r��0|Fc�"D�l{� %A���R3��#�J��>D�$
�hO�`��2�@��s������/D� ��85�PT҄拣L�ȉ8g&)D�����H�z>�)�/�4bU�A�'D�|Sb�:2�%��2P(4H!D����G��\f�L���0���4�,D�$�`�N `n�(T)F�*��̢��<D��y�%Q�(�9�G�sa.�q�<D��9�!դl�=x2Ƈ< ��k:D�$8�GB�\�ȼB�*
a޴�4D�i��Y��6N�o��@@�%D��C0J��=� �c��cN�QN!D�$I�$͇6>��3$R�/<R��#!D��Zplө�6�$�ĭ%�hQ�w+!D��c0$�>ɔ19vLC�3j���t!D�|@W��n�RM���b�(0 �=D�$��i�l�h43K#�q��<D��4�n(�UY)R� dx��>D�p�4(	��lx���Z���ҡ�;D�d!�-�d�L�����B�P!�7D��R1� �����?da�qs׀;LOH�@�7��34�XQ��A��sF���v�;D�L�A��)�  ���@�"��m�!'�IF���ON��XV�N.\�*��W�P!��'ŢMX����zd� ;��N�z��M�
�'��]��/p|d�A6���\_�,��'	T���Y�IdA&Є[�(�c�y��)�ӑF:���CZ�F=TX��M�-q C�I�k?$`�	K�LP�8��)9��C�	�IE�9�qL�|:lY��lC�ɸR�࣢G��e���{"�Y9�pC�ɭ�pYqU)�.�m���2Zd��'(1O?�	?gr�2�H���9����Y�JC�	�m�j��T�'S��UT$Ԙ�<�Ip��໔ϋ TTB5�
�;]��� 1D�T1�o	�t��؃��g���e:ʓi�xˎ�=���9��� K������y��]*v"�M�|�Y�с�
E��i�|FlA��&�1e�֙Hg�"��	I���,�ɯm�-�Ӄ�@����󄁹b��B�	 /�Q:�c��բ$��W|���u؟�i�����=�1�����)5�'D�(V�j�Hw��,Yt\�P`(D���U�^3��}PA/U	v�ڰ$&ʓ�hO�&Z�����X�X� (#��RB�	/\\�Aj�
Z$D6�Cb�ϭS�����.�DJ�L�
 D�92� ���u�!�R�ԤI�+"]:��4:�B"�}�'����+�!�&��'a��%�x�� �)D��(���~B4ق$��zl��E�&D�abΝ �|l���J�QMh�&�/D�8� �_.���֕7�F<yv,-D�� ���2դ��!��t�"%i�"O�!C
�[�.�z4*B��
<$"O�[�aԾ'�d)׈*qX^�8��'�(�<Ad���sp�P��	?|��8�HF�<	�8z���@��$(����JM~'?�S�O[6�	�A�^�r�ƋD�1��H��)��<��Ʊ�΁�C�K:sn^ ��RB�<q�ᔚ�^�Q�+W�I�A��ʔ�<�
��,$8�Z@.���bcم�FX�$�O�3R�K�)}�5�%E§Z��@��'��'�i�v����`�`cW)F� q���'�S���C9K��Yy�E��|7�Уa�X��OF���k�-�d��fj�@�|�q�DyX� �O��9U΁�0^j����p����7"O�%��ގ+��	��NNF�4%I�O&Ͱ$/� Fn�8���70�yy��#}"�'������,D��݈��++�X���O������}�j'�� / �CP�D?C�a~U����ꏩ\+^:�H F�Z��v�>�
��P(&$��7��dB�"
���g	�p����'l$��'���
H���ӮeH&��[�PE �[4w;0�ȓTAf("V���/j8`���f���'�a~��>mP������qT��а=9�{r��_�i#��ݰ,[���D�	��y�b��+@p���0k�y�G�D���'���FyJ~UC�0`c���R�����`9&�UV�' �O��'źl��"G���@���WB1Dy��Q�ܪ��%���`Bǀ2Yݔ���g���?i���CRU���
Ul�i7�X8,�V
Oޅ���?#�V-#Ü	Щ�|2�)�Ss �LIe�j( ��z���'&n����|m��:�,J�}, hs�y"�'�,ѺצT�t��E	{��k
�'��X��1�v4��ũ:N��	�'�>��6�L'h�~PZ�C��5�ޡ��'0��@"Q|�4{Ҡ֟*8%��'������YX�P���ة�	�'A�Q�#�.<[�0��w;d`	�'�`�
љdxȅx���Eb�{�o�'<�'�� ��N�"8�
�K)"��
�'�D�(�#�#y�(�_�Hٖ�u"O���e9>���ҧ3*\IJc���'�ў��,!A�<F�
ё%���T�RX8"O<1���x�&@s�Q<Q�T=3"O�ݪ��-3[jX��F!z�޹C3"O4p�2��7 *a��F0e(���"O�h�q�S�0%KkL6y���"Ox�)�b�1V���P�I�;θk��$8|ODZ�(ג(cؙ�È.Hn���"OM�5�οc�\a:#h��+�yqP�'�	D
4��a-��%�Ш��iN�*����q���qJ�5��{��]�g�ȻM>�������|����0$� � (ɳ"O�i�'��*3�`1C�X,m�*�PA�6�SⓥS"�d�a��Q(��Q#k u�jB䉰 �>�u�SM��yc�n<�C�}"�i5>�C@��V��9J�M[tM�o)����f?i�� |��<��ů?���Q��M[�z�Z�RK�4Di�Ӹx���_�O�h[�j�p?��j�d����,�١FN�e����!D���'͈�-pʥ�QbȦ���C�=,O����Is�
W���Hءe̼8�p5�M<�O�Ϙ'�����%X���kg%��7��MQ���1�g�? ���`��:d�� pQ�R�a��٩�:O����� �慪e�>����&+�44y���$>�ĝ2$�+ٽ-�2��K�[D�~P�d�fعl|X�s���'�L=���*}��'�6�S3V� � ��]۩OVc��D�T���lU�U����8�#�eΞ�yR�T�s[>��eC�-��)���'�ў�	�䂔��y�B۠_��"G"ON}�!�Ʊ?����4��*^0���	g8��A��\��$�!ԩ�Ah�c3D��ذ'
�p1�y:��71��9�2�(�	a�'�N���'֒�܀s�Q6=��,P�'�EyZw(�'~��P3��!�S��km3G�!����`�v��I�r��w.E�l��I.�yR�/ғV�Pa���(ƈD��-WO\$�ȓ$4&��#��$r�V��)W#�6}�O�=�bE��(�Gb�C�АbJ^H�<��:`�Xh3���		���)�o�Fܓ���hO�%;F��2����L/x�O��Z�b9�X��.�E�"����6`�!�D�51I�SFD̢m��LPw����'��'��?I�Dd�"�bAJC��)&�aT�.D����d��b��AwANh �G�O�7�<�S�'��^!+d�2�C[�xp�uΕ r�!���`��0U�?�jq�U5=��o-�|�DؖtoH<�a��)#�y� hӶ�0?�,O��1@�Z���X�.A�W6!��"O���-�;+����gKD2(��+�"O�� �'l�}k��N.
�f0" "O8���LUdy��̐t�"O���&C6��5��J��b�I��"O�s��T�y�9s ��e(���"O��sASB>4�!��S1C� ��s"OT(gl��\� `¥�7�Q��"O`L)2�/aH��Eg�&���"Od!�W�s�Q��E�	w,}�t"O�e��Q7)����پ���!�Ó\uԩ�fɑ�)+�Y �ժ!9!�$���p�I�`O������˿3!��=��@R�J��߀{�,��<!�K
{6V���-�*�}SҊ��&!�$�CJ�k�	I�P�0�)���q!�ѹ+&�	ԠE&D�
�:D�`!��ϫ	�����#5.ʒ���<U!�$���֌�@�E)t�.�ʆ*k!��;y��H�R����ZL;׎4cb!�-p�qu� �<�ܥqQ(�7jI!�d
`�L�����$�28�pD(:!�DZ9:�8p�!��{��t��E!�dA�Ww��J3C�1O�Xc1�	�p�!���;8�����;]d^����D�0�!�dŪM�p� �&��uKv���
�9.�!��N	P����/eI|��)ġR:!��@v�LBf��n�\�q��<_�!�dP�`Dp��Ð_� Չũ��!�D�7ij��)��A�PD�v��?�!��'>�[�D��S�� �Vh�>W�!�d�9=�M�#H��w�T4҄M�2�!��	1Rk�5���	PE�����H�!��9��)���i;�t+u�	1D�!�d��Cdlu�B��>u�V�7�!�$Wp�dʥN#�
�Q��%J/!�H�Ʋ�����l�FY(�g��9�!��R;êm*͎� �Zh�F��i�!�� 4���&:rVѹ�LT�!jp��"O0�`�䕃l&��+˄�s�N��P蒌AF@��J9%�R�A�'�&�PnU��"�5a�.�@��'�*��4[����eQ�����'Ȁ�#�
ϫ�N-�U H�}U��[�'h�Q��ނ\��6���jy����'���"��5C������:g��9��'�1�V��&��!�^�g�T��'&�������9qV=i�ԜZC�I#��"��^|!@�̀��C�	;3S���F�A�%��1m�� q�C�xo�$�GW�:�=s2/� 0�^C�ɞSY��s-J�NΑ����7�C��0����BtI�hh�NI�*C�ɒN�0eqehAL�Lp��:*C�	}�ܐ���˨:�oʔz�C�I�s�b1됎��8�$�¡L��C䉿Mf��� ).p�؅�BڈB䉯(\P�,I�d���P��(	�B�Ɏ����Ǚ�0:��J7�X�	/�B�I���Ī&D��c��ʦ�ܮY^RB�I0���2C�=Cf��#�e�(.��C�	2�x�g�ʚJ��'F�8��C�8��Ei��ܤcq�2�K�	ntB�I�d>B)y�j�h� ��d�/�C��&8v��1eT01�Ԡ��'��Ms B�IZ�a�&� �`��NB�I�p�j�1GM6og�l��`� !�$߼pݐű$�֢5|�i���fe!��'Rc�)(��3|
����Z�W!���7<�� 5+	P9K���!�DM�i�x���W�,�|���ϋ6/��~���5��q�!dF�OS8�9C�.s�T=Xe��u�<IA��4PTL$+n�=�E�S��Z�'jV�rmԕ���~��L��p���m.N���Ya	�W�<1�������+kRl��b�#.Lȑ*\_z����Y?E���[��@�,#[@U�ҌD�i�Ʉȓn�HA���H�q�dh���.Ԕ��:��8���'I:���� ͉��O��(�-��O|0*`�C�S=�H��'��1�
��N���u�hY�Cʌ	B�M��oXI�'+�Ȩ@`V.t �lK�"�#��I�r��"�Z��с��X�H���\�Ӑ8$�u�S���M��a*��B�I[~X\:#		K�t����葵G�7�����J�&U���+�g?1��x(��s+�':�p��L�<��%�$Bm I+#k�
\"���B XZ�D:��R�6�����a+,,��;��O�|#�o2k�*�!A!\76c��'24 ��dg�ę��޼�rE.ƥK��]+e� =?���Q�ȠV��~��PxfHa@l�u���C��4��'��1�p��J Z�����r����>�8�Æ�E*'�NKA�Z�G��B��?=��ZqT2�A�5�� _U���à)\iQ�N��\4��UE,�'�~�o	�	BN��㜠G-T�Z�n���=���X���]�ȁ�7�G�{���U�	:������(~�v4�W^���c/�̺+���ã�؉q����]�eA��D5sKqO��s7ڸ'�]�qq'�ŷvG"bA)��4V<QK��8?���q�)� 9x3E�5�p?�򈇇}��xz3`��uӃm�#*�v`���<���7d���Q^,"���Q�n��hs�8�Ī�"Ϫ0���Y@��0p���SG"O��{do[=Q�����b���ŝ?F���u��<I0E`f�
)]��K�/�?T���˟�D�4u:����$ljݐJ�~;azrb�3�vx�r�?i`�u�jd0��K�̬{������A) Z�t�`��Ե5�ϨO��Rb�
�HEZ6��-ߜ�{���E.Մ�d����	�_�-q�h�5YF�z�n�S��1;S)i�9+�G�U쀉��	�$��DBR��1�
d�5ə#xX�)&��F1��"�$JM �����?a4��B�4J��}����<Y�
=��cRk�<�wf�6x��,�vн`,���n̸yb@�׉�o��� �Rk?�@�>OHh�'���S�? �)"�d��3CoK�f�d�I��'񈍑�Ř2B�Ҡ���2�a5�6�� JZ!s����'�`��3��h����	0�<��ФI�z(vu���['���\¢ʒ]�,��z�+X�0�>�@�'���vg�;V	�e���9D��R��Jnʰb0fU�%��A�IW,dJ���=ф�<�`LS�[��Ijâ�3X��8�5D��H�)�)w0� �Dʂ;=>�9��'�K��W}B�P;��9C��CO�<9e��1�d���:f����@��H�<)6�,lhP^ؔS��/`c�!��b���+sC�UY��XKA$;#FA��p9��%�B9�Ó@�'@N��ȓ@�|m;uH��|���#7��2������R�`q��j�x��	��,2Uy�#%�
ap `�!�YÊ{"���c�� uX` �ޟH!wI�;IQ��P�ᖩR�D��)D��C���:�>i3w�,�us�q�ܼ�G�&o��7��9a� [��5:��S�S9i�ȵ��_�-��A#������DK�o�T���C#�ybOK�����G�� ��{�+[��|;���~�ʓA``�|�'���6bʠS^*!B�χ
�yX�{�gC�(�"T�Ht�O�p8r ̞v0�a��a�e��NǢd��١ǀ��t��d�O�iP(ׇ0���ٕ�"���O��09��O�lj��V�mf��T�i'lz��F�4H���F�����y�'���:#��*�@��-�VSB�-p:z��� ]��R�T3#���:��<%?5��l�6Z&q`��¸	�t����=\O%����(���q�'" 1�$�6wW�ٛ����{Z�y�B��D�IC7��<�r$9�gy�_��8�T��33�Jt�'�����''2��@�Mt���D�DJþ,� 1���+~,p�1d�\;�6�� Γp����"7lOtac'���t��U��n��'f�	s�׷u���[�߅z��d���'{�^,R2&�3`v����S�T�	`$
e�T�� � X!�Đ�B>}1j�67�ZŢ�nC�"�F��&-&L�æF*Z��a�t�!V�8�O�i�O_����j�#-R$)��Ϥc���3�2��D*I�pX���EE��IبD���4+���9F_0vV�B��!X�ԲS�_�h�qFBC�^�=�3�/��4��7�����%�܇y��LI�@!$ވC�	�Ѵݠ�I�)8�$��T�+�z���y�\��ӫ���)�'m�.%���a� �r�A��6��dJ�'g���	�
����ï�&�tC-O,�{3�μp�h˓0�~�C�k��Nd	����'ꖡ��ɭL`��	%킑j��V�?�H�&�	d�ʉ��NX3����SO��sꛭ �*�r�A'(���*Q�x򂃋LU�ţE��9kZU��X$��O�ԍ$���0����,[����	�'s�|�fo�"}��=R�B�c��TgK�i�1�'H\�� ,�.�¸O�'k���(͖[7�W�.E�.�3B�,�<�sc��rr�-F���o�8O��A��ߟ(O���@d��<�����8���HB�p_69�R�ZAA��"qh�c|����	h5y�� Kd���K\�LOڤ�S�@���(
QE:�C֛��Q�����z�D�@T �b���H�D�!�4��ɧ}� h�Ֆj�>�ڢ�S�?VP0��dm��ɔ�o�RH�gA3D�t6�C�	`�/�FL�wC�(-y���>���WV�d!�k�.
dqO�n
�)ڬQ�n�;�j��c ��S����n�v!����A����O9jN��*B.��תE	���q�jҶ(D�D�M�Ffh��I�w�����6�p<��M�9$��!��.?9r�Ƞf�Dh���Nv�D����R~B��>��x��4\��dc:���H�e	�8NO�œ�ċr�O�ӆ#�mZ#3���C�T]©"C�1	LxB䉕	�r�ڂ�	���8g��#L�JP��{b��&d'��vј�a0+��l���@19���ȓ�J4�6�ޟB�����N����'�F�����yWl�b6����@9����'q�����<To*��UďE@jP	�'��Z�՚$;�p��dC�9V��y�y��)�J�%��Dߠca�haJ�	�C�	JZ�(Q����L���Uƅ|#<�ϓ��]��F�$7�T �h\Z����S�? B�Pvnڽe��˔ �k���@b	$4����=>�2D�u�U�iz!F!$LO���r�� ����'�QS��� D�����Q\n=S£B.^����T$4D��K�Á=g$&����D��DO5D�LPT��u�Yp5j�'Y\(�b�>D�D▩^ w���6��0�p�B9D���u� j�ʇ�͇o��Y"*=D�p�L�M���wI	48���S&8�O�	���~��Ɇσ�f�@1'£X ��'�EhS9e�j� �#3>�iN>�#�~¬@�@��9�D�|��J�4dA‒=�d0:W��/�$��	a��u���>S� ���9�$=*����!�"�LKpt�s�c���� �<D���5f�=��c2�"ԣ�+K��O��`C����O�@أ���lx)@"ȧ`ͤU��O�����ŒJɖY� ��yq��!�@>�4��m�!�SvNi�A�H�n��0�t_���êqA�'�e E��F��'Ѥ~�.���J��E�6��HMw�H5:e�P�&��QQ��C�,��LY��4}��i��|���K��^'��\2��Q2�V�\�R,�'�3J�����cPꙠ�OŒ\|:5���4+ĳL�T|h���8���%
���Q�P� HB�@���Od�e'#l�P	��	�'�^�c��L�s��#��K���,ľn��Q?���X�x*֌!@��xH��Bg/"������E�
ܱD:8qb�>1b�����(vv���$�';�L� �+ĸ1��,�e��.5F"a��8OF�#Ӊ
]<��BC��'<�R�P��y�ԟ��j&��||�Q��>$�����,d�i���F�7l�D��"1��
�n�R"���A�$�N�=Zq9�/�)zB��F�ŀ�@ӧ��Dx`�Z�J�I���Mh8@�∥�\r�>`4�tj�1O8�1��§p�(�k���l\):��m𕌂���ɵe���W3	~Vp"��חа<%E]�� �p�Ax�y�� �<!����`�A�$xɦ�J!�o´I��u�
;v��z�ɇJ԰BI
�VoB]���>�OFM�b�_�2�m���8IP�-x���;?�Xh�-��~B-�gr����i�m��A�9HQɧ��ʟ2��y��E66\���AF���O�!�Y�_^�ih�O��H���F6%y��V���JU�"TDy`�'��xu�Ii�S�O��	�X�;�1�t,�%5G&X0�O����/�a�.�O�>��s⒂'����OϘi�l��)1D��y����)�y$JT�V�G�.��U�R�˓
g:��`��~8��C�E[
B>��ȓF=� ņ�F�>�[e*L�Z��ȓ~xA,D�!%D��!�6�T��ȓH������N����T� �T��чȓSY���a0W���P"��%��+X8��l�S~d#B�нB+�!�ȓPvN��O�&��ђ��	?-FH��	���+4��->�d�:p��9Xh�ȓA���ȉ��cP,F�_�,���x�#ef�^��'Ɯ.r�0��*}d��;?}�գ�@�f��h��I��+��S}�J�;�H�`�(�ȓh�Di��F��=�a�
|I�ЅȓqW� ���	���UxD�B&(��ȓ:��p�W'Yc������%���A�U(��M�1�`Q!��& B剪;n�$!���2=Jؙ�,��l>D�؃����{���"��Dq-�1;�?D�X�d��Z��d{d"!z=i�H)D�$"��ǚ<�X����U�52����;D�������4xG�9�J�@�ȗs�<���#oߌ��*�ilpyPcBD�<cn�)c�����[)o�>�3�+�H�<�5La�ͫ�Q!
jl�I K�<�c��26qpb+W����Б�FG�<!�g֜N��f�ܙd�	P4	OA�<)����\�Ru!O�1�8�+P�@G�<�o�t|3'�Z}Z�I�u�F�<�%s���ʑ�(Wx$�2��z�<Qï�
�����JH&�����
r�<� �p��2��p�f�:K��M�"O,�1@��P��s��K��ҡ��"Ol��N�o��t�s�!|��b"O��R�AX)f�ؕq!
%��"O
yK�Z*L!F%27;_�2�"O�m�2́)h�hbi�	�j��A"O\�����,�@�]1Ko(�(�"Od��.�Y�֌ �eD�uAd���"O����+��Pw$�&OW�0)`"O�-��G?%y�L�`c�:A4��"O��%O�}=@�C�!0�a(�"OX�S$H�25�`��"�)(ȡ�"O����%� ��U���k��"O���6�aO�h#�[�M&��!"O�T���_-)DxD�Ԭ�!%n�*�"O�ju�W�mKE� #څ����yR��.0oyR%W,'�:��ꃤ�yb >(/�JF,/Xnij6O���y���}6� ����w��&���y�%�)� l�b��)�ċ��ɢ�y�1]��C.A�O�t�%��8�yr�ʫI����k���Q�@[�yB" jDޱ��tݲ�U� ?�y"'Д8Q�2F��n��DY�%��y��E�&4�aJG ^�)"�H�^8�yR�ٿS�&5!c�%�8��2�y"ɖ�~\��@i��x�+�)�y���5�V���۝| @���O�yBɏ+&�ԋ2O��v�,l�K�yR�ԑ޴�x���r0佚�d)�y2掼nR"����]x��2�A�7�yb)�L� l��̋9�D���C�yRgɀ=��<1	"Q���yb�/n�h��%%�l `��y�π�y�r�7'D�y,�ා�2�y���4鰁%Jެsxʝ $�y��E��,B�B�4Y���:LI�y2�Sbd(aR3M/]��i2�o��y���	Y�2�3�à �fpI��9�y���=w-Ra�i�Bm�!-�"�yJ��F[p���ԅc��U�`g��y".��)M2� �ҟc¹�0-P��y�[4����C�g����铏�y�k\�;�|�@�
�
���ؤH� �y���*��10��U�t��8˳e�y�D��:Qbad���z?
!C����ybK�$h���VM֏h���X���y��	K�@9�i�4l���#t!��yo �CFT�2�$E"�����y��(tnpM�ѷ"���R���
�y�,G��ٛ@Z%V���J���yҪ�� �\�V�Y�<99��Q��y-��D:��CN�9�0���yH�l��LN��$=Y$C�2�yr�W�;UѰ��t�H��s�@��=�N��;|�W���N�n4D3�͖��X��	��c��!9>���L�2�6��=iDHtZ@؍���B����M�1x�ȃ�	]!���9wK6�H#I�x:�
t��XyP�K�����	��"|�'2��)�$ׂ5NL� TY ̌0�'�0ژu��� ���$�0}U�� %�����@x8�TY�kU<�:���	O3���&�6LO�L�$'����Y��'�)RЬ ���D�0j0�P��'�4%e�b��<��g����y¤�
b�ꅳ���p�π �I���'+�z�Ç���:��"O"��*��S� %h&��6K�(�0��O�\\+M�X26!?�g~��˰��M��ʠs��;�fʉ�y"j�!*18�f���,}��J:L��ePrᓁ7mα��IN�p�R��}��2� �%|x���D�	<KT�c�B���~2���q�0�S��Ҏd�H=`��С�ya�0W����C��P&��A������'Nְ�m�	��?�:��:��)
E��E�޸��j/D�X��,��I���
E�C��(3_�X�="�>�#Wa!�A%���yI:D�gM
a�<���9��E��K�s~8m3�]i�<I�ر\�z�*��7`t��Zg@�k�<���_m�N}p�A�&�@�;���I�<a�D��2��u�۸X�:��^�<F��<2��)������P�Z��B��z��)1 �Ц���x!��
%�B�	�w�h0���M�#�����%�;`�~���*��+�)+�Odq+�DXTB%��C�?b��Yc���s3H��=�O|���Ⱦ`��MC�o�O��y��"Fc����Z1ex�4�b"O��Fj���jL����Y
��c�i�L]��bV�Hs��(փC��D�#�ڨJ��)�	�$*��2c�lH�I���z�`[�z�H�˲-��<A�HЉrOؙ��K� #�r�ˤA�1@��xW����	�Q>�n���Zfj�0d�("�.C2��H�=q���rt�P�t4�'��l�"�@����-��زp�'y,���$Ș�a{�3?a D��.�8O��i�,�V�X ��� %��ɠf��-2�AW'��G�Z9�4Em��X��۶tg�|hm�{60��ȓ�~}j$��
����0 pm��h�I�C>@�� �L��}P�L��`}�S���~�1R��������ҧl��H�'��(�4��-9	�R��4���Y�$,�"��="D�aU.�4��Y��0��<A�#Į*w� h�l��?��0���W�@j�T�ժ
�%r#~��oF!<�H}Bre�1Z�%p�L�h�b �3o�'P����'w2��d�!5D��H��-��U��C�MO\�qĜ�~��D�P�h�b�aa�'��}aB+�!B�E5�[0�&�8�'���q�@�b�x���+K+%m�!C�4��-0I>�d��%U7ǔ�)dMc�	��T�+
��$i��_�FD3����{k�{�(�4b:��F��(���B�C�F]���%N+&��b@mH<9rm�o ����0rj@�+w��_�'}�D���`(5�~Z�
W�pw�U)�\$�����X�<)t�ô-��X��C�\�2-�R���D��k�.�⥚>E�4-�0_��i���-7�����%ϐ�!�J��e��苄?��]����7��$��
u")�V'���<	B�F�x@�$B���R�]x��h`O$C���"���6<4�x�H!mY[��X�f���їȁUn!�dQ�t����s�ҍ|.K4 ��y�'��L2��@%8�<Z�ޖwt�A���d��=%p�A�CEV���ʦ���y2� p�)а�fA�6a���U��p�1��"F#.h;��+ܸO�' <8�va��'v��`�U�g ���'�q��<T_H$��3u�8�Rr��9hz���Ĳ :�({�����<� 
��[�.5��#V(і�j��{8����
�^� Xs֪��c�:��3f �|��y�2��	�ň�?�!�Ė
Hf��t-.y漈��\�	Y����#�>���қ���!�E�f8(�����!�;
_*�`C���=�rq�e �>��Е>��J L��>�O��b�'!���S�ٖoIb�;�
O�U���^�G[&l��Q�R�6�J�샵k���(4��'�0?*����k��1�
��D��v8�L:�o��e��:𓟔��L�R 8U{P-��{N�p�*O�����AO���R$�/ �Ǖx"�H�4Z
(F�|��d�ߗq���0lK#$�(pN-�yŔ�L&��B����v������$�DL�g�D��z|DM��KM�:֍îY�!��:F��t��,�Y����P�>�!�
*1I�5C��?.b��m�!��̄s|�UG�3z�f� ��0�!�� zM�r�
�����Ƙe2Lk'"O��S&l4;�б���	*�5��"O`��[�Q��́1CT8s���"O.8 tD�	�vH2�HlbD�"O�t��VEӺ�SF�'dN8�"O.�)�h��M��P�#kM�$]zD��"OA�cC+-9b5J�*�* ���"O|H*�E�<
p"_�]u`)Ic"O��L�r�FE���dPl�U"OP5IbCV"r¬�P�C@pP��"O��R1��5�t�u��v�j�I�"O��b�Z�����S^����R"Ot�k5,;v��rF��o�Ԕb$�'����*��x/��2g�yI����O���{�	��j�WN���ٗ2�
\E}2.�!)��a��i�9,��)�9�Cr��TX!�D2k+Z����Lp�"�T�2H�	<�l`k�7��)��3J0)��Q�Hؤ<���  �2�U��!
%!�PΔ��(S
{E��A��V�ɦ�4#f�!�2��Aj�3?�i&���>cG� ��,Q= ��{��-L\�?�#�E�:�[���l�Z���(6c	+7j��U�!HR� �E��c6��J�`��\�S�O1ƹA��]�w����@@�b����]��U�/���pk�D�i�*klv�>�r�N;Y�|���ڱ �Xy'n�<�%��1o�f��"�=,O����Y`.�e�1S6�يT4O4���f�X�Z�۬ID�'�F�jF6Z���[��K�v 䨀*�h�"5sfm0�P z�1�\ *@�� ��(�%�%/E#�G�H"�:RHk� y�"Q�6d��`�, ����^����?��*J�<t�+䨘�n�\x���<�{��|��'�3A���i�_ (�gj2N1h�s `�0�4�{��B�0�=�4�ƺ.jC����)�'	H��5�L�rb���闩KB��'d�y���D?K�F%̓ ��J�fX:�T�>����(L�����ٯC&ȕ��Ƣ<�S�Ra��*/,OBi�S�_��EK�G�}:Z��!0O�����5�n��g� �il��Hw�F�38��P^���Y����[�|���F#"ܽC�&НP�����	Ň��l2�ǟ0X�����h ���}8��m�����BI�G�i>�X�ŤM���q��C�4V�`*��!�5ZZT℩ܟ{>�DT�Ѣb
%(G�!�F�F8<�Z����S���Ij�l�����S[B��"Pa@t����-�2�
2����]���S�O	�0 E�b���"AE�yf��1�'v�ECv��J[�A���r]���N>�šs_���dB7`�������{�蚃A~!�$�(2�D�R���^�,��uA1k�!�D'7=pTKr�����A
�W�!�$�{�tZ� %aɂ@B�V�!�	�"%�wOZ/�0�o��!��6cSB�QA�_6f��Q4��6�!�dE8H{t9��T>a����햤�!��7O�6p���	qgDh�K9:�!����(��&WR�����Y:G�!��a=,�� ص6w��#�#�yM!�DL%�����C�xt��2$��'#!�ė<g�l7� �G3��XP㗘o)!����(�P�H��8���b(�0d!��O0(FA����2:���S�A��!��P�8�B@'�u̔��Ꮛ;�!��?y�Ȭ�$kĉ ���RV �e�!���<{F@�buC�� ���`!'�!�d�L2ޑ;��[�4��� ��S�hq!�51j�P7劔H(����@�
l!�d��P}�E��
�qR��C�N��!�D��2�2��4�Q�	$I��nH3/�!�ϖ}���h���#4�������N�!������bo^S,0Tr[\�!�DE �p��J.>A1w��!�!�$��K,�$qw�y�i���+i�!��Fg>�Y�ׇ.L��LS!�!�� ��dsK�9��F�%h�$�"�"O�󀝶K�L����,���C"Oj���)F�;�Ta�O��v�P1"O�1B�g![��U9Pm�{��л�"O�q�6`"*�X<J��L�h�:<�"O4���.���˧צ\�)�"O��i��Ƌa�@0��HI��.���"O �p��"w�.@�Ԫ$��"O@�1�kL�Je�A��A$�"mc0"OV�b��w\mi�#��
'"�9$D��lA<<����a)Z$Q"p�;Pb�0{��O�SU����2(U�Ah2����4L$ Y՚>�Ƀ�!i�L�|M~�iLeRr��ӏ�-M�.��� RB��_�[��YH��A$�0|b���T |����&Ul�j��|?	�C��6�:p�6}��� �5	Z�iA)��,���J��+<�S��U�@���>E�t�J��S+��Q�d҄ș%1F��j�$>� <�M����.6Mp5�ᓬL-dD����=�����#!9����b$M�-�JK�8�C�~z��)ϵ�n� �J����Q��%8�X���R�V�q��]�>+bDP�S?�F��ɜ[����R*
 IZt�	�I@��?��

�,����e@��)�GҜ-{�L�\%x�	���X�Xp4�2�}�E��p���"�f�[6�K4xB"l���Ǩx�A�>e��@�7�V?1V���L�$��@�"�lT�MNR���P�@��� ԭb�D����t@�~�	&�I�|��)FT|���umn)�1_�4���/txY�۴R�a@�J?֝ݟT�l�a��}��JV/s��!@�J~Ӕ�)!��`j� e��]I�O��Sm��T��	��լx@>�O<AJ�+Y��xn�:�PG��)h�*Tk@�@6>�"@�� l0�	� ���i��Ȏ���d��B��4,�j�N�gBҊ��	�nԛ<�?O��AH�<t��wl_�)o�Z\�|��h~�a��F�"D�E'��t�>ɍ����D�<+�(z��%O���k�����0>��fķGpe9��A�0�,�`i0.kDx�a��+� ��C��S���`E��j=:E%2�ɚA�LU��S�w��eZc��;���bP
F(�O��'� ��Hv˧V�$��o&b$V�V #����F��8;Jr�'�l:���l�����>﨟輨�.۾4�J��b��6i>B7�'��CÍ�*,�ʤa�Ɠ�t"a���ֵ
��t٣�M�h��y�Ҋ����h��}�
�Jf�qP��ˁB�xS6͇�D1xu��?N~Lb��؊lZ����)�d���ujJ(�A2)lZ}�ۍo2Ɇ�����r�˖���P�AS�6u��Lj�
�dV�Wy����
?�D��ȓ^��)c����LW�T8+��C�fD��`q�I��O$�P���	;>/&���OD�@�-�8��d�7�2%��]z����&`M��PîB�Tơ���e+��H �0�kG�!��Ćȓ]��'�7l��Ҷ��gt���>�\�':SeL�F��?^z��ȓUa����Ί�p�H�fE
��@`�ȓ�H�SSi�zP� �P::���C�^�CtH�M�����A]2.8.Y�ȓ���'�ӭz'&X�cҵQ�J9�ȓ \�}��Gεw�ACA�\�p�ȓu#jm!#�1v��DCƇFK(�ȓ	���{Q�Z�3�`4�p��o�,��ȓ]���Al %ˁ#J�%.���p���cI):�n���"R3�d�ȓ���0�ˋ�t�Υ�t%��-��b��]8q��XDpS$�]	�͆�L� '��p�������Xc"��ȓc��,�"�ޞ+�<I1$��,ex��ȓ�e�a�FH}����fV�]jņȓ"�H'�J�Jf���uL�:F����X���)��#(�!�"GW< �&̈́ȓ3��\*�k.���� xp��S�? (�#`:6���ِHƌ.�ͪ"O��vE��A��QBBH@0��i�b"O`�[��PP��eSe�*���d"ON{���a~,H�W�+jd�i�"O�av�)=��V��-�BIx�"Ov5����a��*��w�����"O��a� �`=(���	�.[3�y���r����c	H4�l����y¢�'`��
�ʝt˨1ᓉ��y��@�������aI�U�r�T>�yd��L��H��� B��8Â�̖�y�'[��D��ʒIU�8C��yr�סp^��d�A�@�$��a����y�j��7BPh1��7h�ݛ!l_��yR�҇!�8�0��_�,a�9@鏁�y"^!8�tX�G)���,(�Pn�0�y���IHbY�T�D&z�vؐu�M��yb91�\[�b��ZD�o
�y��>`
Ⱥ����"�L�Ys�ʊ�y��</�Չ�E	.n<pg���y�&r�� A'ȸ_�$�	U�H��y�3s�1��	͔,Y�<����3�y�tb��!�������/]��y2� ��l��	��n�n�94� �yr�}�B�1���f\Ą�I��yrǤdL���K�O8�))`����y��P�鰤��HB'L�h	ڒ.@��y�g��g9X�pK�:���/W�y"*Z" s@X;@�RW-E"�y�OL�p��{��Iw���y��	G�&N�z��|���_+�y2B�h�r�3��=��2&���y�'M�>�2I`�O�3;��P�Iȭ�y�޹Jf
�x�䈧%@���Vg�,�yrj���s�J}�)�����y҄��7��1�!�;�@� Dᘰ�y2�M�D���0M�70�E@���yR���Rd(J�+إ�u.�$�y��K��<� P(T�o+�Up5Ȃ��y�"�k�F9Jq�C�c?j$)ƦO��y��!�viI�⁻*�2�զ���yB���`�|xҠ+hH	E%���yb��{>��H�ۺo3�m��*�yB�o9Ry�cM�9j�H�C!���yB�@_u�U���aݮ��B��y�6x��`�LU�x\	abD�*�yRhӆf2���eӺ6g����dҥ�y�X;����BC#,�(!���\.�y�8m�������e�֬܈�y��:��A���t4����y��O"�R
� �-`�N5�A����y"M�*R�8�x ��
D�Q�1)E!�y�Cբrj��6�Rx��(��y�`%2]�����(�$�I�K�'�y�mN��������Z�qa'J,�yb�6�|s�DX�0��s�̏�y��ܮKN�	@�1�6U:�bP�y�J�^��'�8?�jXB���yҏXK6��(�hC=n�x�Æ�7�y�L%M+�;�/�Z� H �́��yr�It�.� �ũW2���*й�y��\����MKU :�������y��څEl<C&�E#}J��'̔��y�	�R��%��'S8xܔy��	��y
� $b���X��k��[9�ִ1�"O>�iP\A�5k�C-\n�a��"O�R�e��h��䡕���t\��1"O��;P�؎zMĝ�6(K�H �d� "O]�3l��&�zI��ң"O�kS���+|��s���4)��"O��rf'�'LBtɂcfR��U�&"O��(� U�C�Tu�S	��
�"O�qSV�����W��~����"O�����8�P,�6�	��9�"O������%���g���*�I5"O`�4�G���٠�bD�w���5"O�}�5�ٶ[L��y2�)�y�"O��"ca��2l9vaӼ)V)�W"O~���M&R?.����T�z�"OfH)W)N�S��d D������"OU�2%C vm̅����%�^��"OɛN�5H4��3�]�TAn�w"O +r��PJ؅�b�ݭ1�42s"O�q
�扝w;K嫐��Z�"O�`�V�Ӏ7�d�4���*�dL"O�u!��Xh��aM�G��`"Od�B�">
Za�j��b;V���"O�E���  Dz�oL+N4�u�"O*����.'�:���Ͼ3���""Op=��� �9"�m�JR�$C"O���`��b[�,�
K'h�Q6"O:h�U
��W��$�P�̴ 9\�@"O�<����¥�T��RP��S�"O�U�E�Z/T�M�Pb@�5����"O8�"�n��`bZ�q�BX�`9��"O4=�0▐V)2$c���p�8�s"O�d:�BƸw^
���]6[Vvݐc"O�\� ��S ,��E�+p���"O�[�c߄)}Ȩ��c��X0�"O\U��[��	�bB[�8�=X"OP���bOزE�G}ܝӣ"O�����������%΀�}oVB�"Oh<�Eo�$�@��*�3r_(\�5"O$��r C>����@	 
�x�P"O�4`�Jͤd�ء���6�@G"O��``��)A��B7��k5�(�"O��x�ǅ��2ex�L��w����"O^���Z�T�ܤaQ�V�uV��c�"OD��bH�}�r�P1��j=T��P"O�A�ի�1�riQgFC�uG:�"�"O�Ir�lF 1��d�
C+!��i�"O���+ X1������b"O��l����ɶ)U)%�
i�5"OR!g��0:H@�
Ȭo��D�Q"Obe��섳�����]�wκe:u"OT���#�*Yv�����N��x�"Od��gݨ�l}HA��<q��Cq"O�Dz�E!fY���fd��k��y�$"O`�җD��<�\0��ɽd���b�"OHɉ'f
3���t�̡in�� �"O|����׽9��[�ɓ.[�Xp%"O6��F#V<I�j\ң'�/@Wt���"O
�+CK�F%�PF�]�8YS"O���� ��q�"yq(7~Q+�"O����P���F/$�yV"OZ�r��J)&����&��7��D+E"O������|e�4y��pwAk�"O�#�_T�q���˯FEu�Q"O� ��k���qh)����04QXd"Ot5
W	M�(��q�[,#��H1"O�9��є&�vh�&�pe�t�"OTxf�:��	�� 9J��Q"Ox�)A͏�y�赩����"7��W"O� A��Y��
ҋ_	��R�"OV9@,B~���sT�N.��	�"O�ų���:F�1�D!��!��"O �A��̈A
������Q"O�|8��J�i�p�!��O=	�N!Z�"O�RpEPvA`���(*l�܉�"O�=���k�P��凗)>�-�"OrqRf��+: 4����08�iD"O��,M�i��+U
&��6C���y���$j��	��Ӆ*D\1'��y��ռ
EP�R�'l���5��(�y�7f�H�2큼m60��,��yb�^8VVb�b)�0d |�	�b
��y���̚%��Ƹ���O� �y�(�eL�	���Ѩ�3�Q�yB�M�L	�)RL�< h�"��y"�x\��0%�!a>e�!!G��y�̎+�n��c��щ��yRP���H��bW�I��ba�-�yb��ZZ�C0+*FKJ �E�:�yb��6hW��C�DJG1���c#��yr,�:�h�c�B-P$!���8�yb	�*2D�7 ��At �����y���";gT�X#�_�c2��� g�2�y")F:Uľ(P!(�_��R���yҩN�7x<�bo��Q{��( g��yR�N��x�A X+�d�I�,S�y�m�Pز�k��`���X��y�Ό�1&�`j�g��+	��RW�M$�yrD��zNR��!�FaA��yҮ����ӥ��򩂀O�.�y"�C�>���
�$�����,�ybo� ������R���Rb埂�yR�?�Թ2�E�8S���f
G��y�HG    ��   �  i  �    �*  �6  UB  �H  �Q  X  J^  �d  �j  q  Zw  �}  ��  _�  א  1�  s�  ��  ��  <�  �  ��  ?�  ��  ��  �  ��  �  L�  ��  ��  ��   ^   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.�T�DxB�'��PnS�8�2 �f6Q��$��'#j��G  �?�	{7�>� %k�'A�)0�˲e!>�i���%��ə��(Oz�J��_�c�q7(�4GW�ȱ"Oр�Hr�́a6-�E�	f��E{��i�dI�hSm�?�4��Ń�	O!�?�[5)ɂPɌIP��vY!�D+q#b��@^����A�芢
I!�� ���2iR�7�`���R�/PFxe"OP���]���A(�1�4AV"OPձW
�=~�����T�Z�[c"ON!)�fi�	5 �H�4 ��d,�S��:6T�����x�d@�PoxB䉆��i�7�Ʌ4�0�sl."J�"=IǓ�VUP�͎
#nDc���0���ȓu���Т�1�Рxԋ��B�J�<�指�$Ҏ�3�Kh|Y��B�<)��ݧ|@�����E�D��v�<��胹����g��>6X]tg^n�<a�B��m����w)�C�ɟ��b/��C��Y(�r4b�O�����7� ���I��&�PU8�.�x�!�F�3@(�Q�K?<�X�pG+1��	@��̫7�\�Mİ��nW�_UTyKa
-������~¶��k�%^��L �f K"1m�O(<���S��3F��e�h`WGK?i����n�NQ��N��a����$�@=c�C�	�EP
���cJ�z�̀�C��_;J���<��'����O�3�I9Hj)�.@P��5��8<�DC�	� �y�cbN*B�{����M�C�	o�������9��%Bm��Z%�>��)�#Q�����g�^,ц��[!�Q/�$�p1��6a���F���!��1&�̉�"��'�zDBcFM�	!��H��Q��Q�qc�;�$�%7c�'�a|�O$�4��&�Et�2�	/�y�F\�r8bf��st�4�p. �y�G�2:Ѯ�15�a�2,@�I��y!U�p�n��7��3Zcb@c2ب�y�K��*��U�N�`V<������'�ў��ȍ�E�Z(
��2�Pc"O���R(�/(�z���_�{��hB��0L��x��;Y�ȍH�*W��4����y�GO1�DՃ ��2�j�# 3�y"GL5~X�"�<��H��yR%�|����!5��H�숝�y�埕t�\�ƥ�GfU!���y�&֗���9 �O+D'��R�b�y��<s�|y�T
E�?���rʔ0�y���lV(-����%ېP���	�y�f<V��v�T#�����2�y�윖t}HI��/0_|l�e���y2'   ^"���*E#h�RqoI��y� �60 ijQ�>�>���H�yB%�s��h�V���=�V�Rd���y�G�7<0��!�mS(*B�PDB^��y���xQ�D����a��Q�y���9P�Z�����ty�F��y�M�'e�\���R"����w���y2�.+��LyV��~�@`�!B��y�b�2���zb�3.qj���)��y�C�=F�o�#S88Y6�Ƴ�yRE�t/�@��<U@����U�yr�٩,HY9�#I4W ֨�d�ݰ�yrB��Cl��uiO,{����ʑ�yܑ*vp3%'��K��P���	i�fO@LD��0��ƛA(��ȓl���ce�}�ZP pʘ1q�Q�ȓ4 xI���c�,��D���A�ȓ *�m�(�� ���
66m�ԇȓAW^�2e���5A=a!�� ���J��!���l��������S�? H�ق��"c�����s��!�"O
����M��HP�� +t���1"Ot��c��'O��	�B � ��kg"Oa�4G��T���dI�$2�2�"Ol��Q)sN�c����'#�-�t"O k���,b&��5<��t"O���T�#$?bl�g��1��� 6"O� �pa¼�0|Sp��03��Y"O"����|�����V�	���%"O.P�b�ۯ/v�����k��c!�ڂ/ov�AFl����I��+@�6�!��u��x��d.ƘUʏ� �!�dW!=~ �����]%0�(��:�!��C�j�C$)Pa�G	�1�!�D��w�6���p���(���C䉆��x���X�	�ε�b�EV��C�ɷ<}��;0EL�j�	I3(ޗW�C�	�|���v��g��-���APC�ɭ\���C�͊�4����˸ PXB�I�(u"���dDP_|��R�ɋJ&�C䉊5���*���T�DmKJD|� B�I�t�xMz&��8�.ٺ�IA��^C䉡/�n�.6d%*e�@> }���sSD3¥�O�q�/	=z����ȓp�\I�E�P\�сN7n�� �ȓ4�zPP� ,"�|����.]�(��V��VE�$��2�%
!}��`�ȓ�2�36g�"v,��*		W����t-jv�1�2����񎔇ȓk��
�eׂ5�����J��X��Yv���N�w�
���Z�;{X�ȓg�Zx�5�N3�f���#L�%����#�����J�J�b�{�K�3g8���Bq��t�	�=�N|k�H$fK�H�ȓ
�B�Ba�D5r�(e٠$�B��ȓ\}L��Q
K�G^��Xp��#��$���8-Q��جJ��U�¢n'�y��`��@�#�^!v$�7e��(&���K�ɚc� �N\;g,�<a�$����,��Ǡb\�ď��s.���S�u��O��^��=����?q]�݆�!.���U���җ<:U�Іȓ�6���	���R���;y��L���������h��e�tQ�ȓS�H�2�c��Y�!`Za��)�ȓ���)�I4�"7ɔ #��Ԇȓs�~�#�/a��┘U�|�ȓO����Ȓ��)c��>Y.�ȓO��|��]��`q��5�de��k��x��LāG1�LI n�Gp�X��\�V5kd�L�6�:©ݾ='����\�T�؁ŃO��P�$�Y�?�Lx�ȓ���ů�*~Pek�f�6;�D��ȓ1����`^�zt�	[u��(�>��,3,=i�ą�\�*���-�=��G(a�7�ݑ+���2M 0��!�ȓJv���I;�q �ϗ9kx]�ȓ�4hr�"=C��A�Iʑ=͆��N�|�H�j�hD>�����^��ȓ5��{���1(��v�˪d)�ȓ�Pm eƇ���T'$i����y(�13��3\uT�iĤI H��X�ȓp�<E�V�-�0A�MtK6��ȓ�6�A+�T���KW�ü=�~���S�? P�k%H1�輣�+C�B��"OV���U)%�"EhD�Ow�l�'"O����OB�UVE���!�|Q�w"OD%Z��l���&�:k�<tH�"O���0k�����aH ������'���ٟ����	韨�����I,tvɲ�NE�E����'�|�I�`��۟��	柠����	ɟT�ɨ =���V�Î[�`�Ƈ�*N-vd�I֟�	ҟ`��֟���ǟ����X�ɕ#ﴠ�w �4#p��螄p}��ݟ8�	��P���$�I����Iğ���_�
 �t�M!���b�G��]O���I����	���	ϟ�����P��ߟ|��9}B��a7�Q�l$X�����z��$��L���\���8�	����	��I�0P�ea
1� z&�T<}8���ڟ������	럸�����������I�PA�q�ӧa��]+jD,�������	� �����I�������I3�$AQ���-B�m;�W�8 �9���,�	ȟ�I��	П����I(c3�qS��^�B�@��W*�=_'(�����	����������I����I�)u�T)vB<";��fLħ.+RT��ڟ4�Iǟh��䟼���@�I�|�	�w��)�Ɏ6(��1�M�ff���	ן��ş����d�	�h��ϟ���	V���6f��(�,@+12>�	Ο���ן��I����ڟl"ٴ�?9�}D�K�n H� �ON�-�QWT��	y���O,�n%�^L���ܮ*����EK�0�RP�"�%?���i��O�9O����-t<���C$m����EL�d�O�$r�r����$��$�O_�h���4j���RɀF�b0�yB�'��V�O������^�q$V]*B=h_�1A�l�f�s#��4�Ӟ�M�;U�"M����-V0���L* ��P��?љ'-�)��8'y ilZ�<��!�=�e�APht��d��<��'�$A��hO�)�O��Ѣ�АsaZ���v-���0O˓��ji�&�2Ę'������fڶ����"${<�����e}��'��=O,�)9�<���Єum�u�Q��Ar�$�'���,p��,���#��(5�'�F��7gş ��=��L؍cT���]�<�'U��9O�Til�*�~����Y;��q�:O@�l�!x�x�=_��4�F|	�"R.r�����X��-A7O���O��D�>Y~6�(?��O�B�	��|<� ���f���``�[�3}\qI>i(O���O����O��D�O��G� ���[r艎K�~��pį<�0�iG��;�[����S�ߟ�qGJX����Aȓ�c�4�jQ��DLΦ0�4g=�����O��t���<siZ�CZM�d��=8&И�iB����ZX���1BL?�I���R�a1��icr�k�b�=a�d����؟�����@�	՟�SOy"}��	g%�O�a��d5���A��9v>]Y�$�O�yoW�{��	�M�R�i�47��J>�!OE�v���� _
�)C'`�6物9U���̋#���B�<�+H�����VQ8l8!/�6g��1A!�U����Ɵ���֟��Iџ��	s��%�j]#��Z3X��P�Lު6	��y*Oz�����4m>��	��M�M>Y6iAD>*�k�Tx�.�d��'J�6���i��(} �l��<��f�A9��K�5�*�A�^�-����臬rO��D������O���O���6�:����$�A��		�~���OF˓r���PA2���ЖO��� ��P�XsF܀�oD3o޾���O���'~�6�Ҧ� L<�'�Z!'�*?���y��[�1�H�`C�?r��Z%Fݓ�M�R���S�1��D,��ol�J�G}&�Y��1>mV���O��$�O����<�&�i����ƀI04 ��
�U�~(�R�.�&m�'D7m%����$�ަիF(��M~mGte����	��M��i�u���i���O�`b���R�o/?C��4T"���ڻ��-	��|�@�'���'bb�'��'Q哚o�� `�`RV!�9����4���4|9�H:��?�����<����y�R�^d~Y
�Oڔ%�F�:�ʐ8�(7����N<ͧ�r�'%�f b�4�yB.Dh�u������gj�Γ{�����On��K>�,O��d�O��qSa�y��P�����򄬩���O���O��D�<1T�i@�B �'X�'��t1�QN�|1�Ϸu���s��$�^}2�q� �n����]B�)R9�Q�����J�Γ�?IC�
o��Sp�4���
�a��R�F��$m�"x�)֙c3�����N�d�O4��O���2����*�V	XTJ��P�L�*I�vL��?�7�iو���Y�d8�4���y-�K�)�5KJ3Wߪq�ACP/�y��q��LmZ#�M���M��'s����-��'j��<�u�ʁ0M�p�M�-��L>�+O8�$�O��d�O\���O�0	�EȚ'�S�i�I%�h����<���iw~9#A�'T��'���y�C׭���'����yFJ�.n`��?Y�4S8ɧB���br�D<	�c��sօXKE�NP C1AК��A�Q�xQQ��Fk��O|˓˜L��`��U���"fCY�}.��j���?Q��?���|�,O`ql�Y�z=�I4)�x]�w@eY�����4lK�;O|�og�M��	��do�4�Mۢ�s(=f��0��5��y�|L��4�y�B��V�������?mz�8O����he�=� ���^��Ea�M ��8Ѡ:O��d�O����OL�d�O��?��-[+l&�+g�
�\�H���-�Jy��'3&7M A����M�����^�n��$Q���!dW�;�h�~y�'��o$�M���*cI��4�yZw���G��e�H�B�@9l2Y�g!�!Y�x���'�&�|�.O^���O����O���!˦j�n-	�=I�]�Aj�O��d�<�ջi�dh���'��'��>U�|��� Q�i���I���n7��S�ꇱY��P[WCB�u�2X��+�z�~P��H�
em�&ȵ<ͧJ�\��y�ɢk��y��� �Iy�N*�t�	��h��ݟ��)�Qy��Ӭ0��&~�HI�cnG�

�I8CË�a������DF|}�ak�l!@��P�>�J�C����3�A�֦9�ش4k�iߴ�y��'�,�f�Us�,OT	��f � ������5��?Oʓ�?I���?	���?����) ���}�7��շ���m�Y��ij�&�'�2�'��y��l��&4XdрS�8�˄�X'3�mn+�MӴ�x�O���O̬*�it�Č�6�2HXW�T�.����D>>󤃄85ڴy�o�ؒO�ʓ�?	��S���r�.�'E@wc�����?9��?q.OvhnڛFv@�I� �I�	C�5�5��&�%��h��w��I�?�T^���ݴ}���"�>��������'�<�I�"���O(�V(��h��Qͽ<Y�'7���H��?)%,K+Q�$ec�6p`��e�E��?	���?y��?1��i�O&����0o#ȸ�׋M=&�2u\0�$���q���Zyr�d����,=l+A�r�P�1�m�,T=b��ɦ�1ߴ#'����b��=On��Ή�T���O��u؆���]r4�9E��;I\�qs�|rR���	��X��Ο������wg�3��3�T;`�N
$dUyr)i�J��p��O����O��?�R��	�P�Ԑ��%�/?�@�V%���T����4cՉ����O���Z�):>�P���)z0@�&O�(:��Z��E�=xbO�y�Sy��W�.����6f�_�X1�,\�&F��'F��'��O����Mˠ���?��!����Ʃݩ"�����?Ɂ�i��O:��'�¾i�26�$(�ҭI4V�5�l�#�ݣg-��Qw�x�4�	ٟ{d�JZ�dh�~yB�O��
�0�,`��K�\6l`A3E�%�y2�'�2�'L��'���iJ�Y�m Sa��B�N��V@s&����O��䦩�t��Ty�"d��O"];Q�צ�c*R�+�|�XbRu�I<�M�ǳi�����s|��<O���ҵ^��4�6I	�|`�h"*��q"����?�&��<����?y���?Af�^B��A�DW$N:vD�����?�����dXЦuh��쟼�I�`��?���	�=�u"� �I
�!�a"'?��X���ٴ`q�F�%�4��I�;U�A��c��s�n(0��88��G%=
�HCǪ�<��''���+��L:T�2@N��F�F���u��T��?���?��Ş��DĦe0�R�Jo�lV�.+���V�I�,��'��6m7��-��$��is�"��Nh!��)�5h��r�թ�MK�iV�x�e�i��D�O�|D������<1��D�e��3��O�s�꼓4��<y.O����O��d�O��D�O@˧.�TS�*!_���%l�1tHdx��i:p )��'���'W��yr�o���]��CW�S�+F���#{N|m��M�t�x�Ou���O��}�Ѽid�Ĉ=�1�nC"bTڸ`W�~,�d3�(��t%�O
ʓ�?I�WE2�����t���"W�QފI@��?����?),O��oZ$kBܗ'��!��u��u$�$y�u�6J^��O�'��i{�O�apR�˦UHe��@Ct�S=O�$Q�bT99�'�:�@˓����O��Z��%�A�>��L���1u�� '�������㟀�Iş�G�T�'�<��n#
m�ݛ���,!�I��'��6�DS��˓` ���4�P����ݰo� �d�Tk@���8O�o��Ms4�i��ƹi6��O@�`Ҍ���Ŗ2	�m�$N�)�Ht�"�)@���O@��?���?����?a���X�a���^.��	�OibT�)O��m��i�u��͟���A�s�x�1ߧN݈HTO�E0�Ǘ����̦AIݴ	������O;��#[L����+A6(-��٣�Z|F���Y:�� *j�e�'p��&���'`yP��Z�X����@�U��`S��'V�'������W�`r�4a��,Q��s@0�j�.�'2�b,�j������'��'��k����~��	mZR��0���9!�v4��厏]�b�sG)�Φ�͓�?�+�!���釅���䟸��N�R
,J���H�}�7���e'��O����O�i\��'��hy���zv$ȕ�^�.���"�O��d�OB�n��6@��'�6�4�Ď0*^V��u&�Ȳ��$��'��شZ�6�O1Vp*�iO��O�3䥁=�v�hՍP�nn�%�(J,ܣ�'��'�	�t����	<�֝���&m��T��b��p�I����'d\6m�&�E�'���'1�S�?.0ɘ��>n�f �� A�mX�o��I��M�ѷi0�O�	���y�@''�:Ǉ�\��A�5�3٢@i�- t����C��O�UhL>�0j��i^��i��_(Ҧ@������?9��?y��?�|�+O�$nZ)}T�):�/��lahZ�/��9Úcyboe�h�H�Or�nZp��@�ah��c��P�[�����4E6�&O&�v;O��Ē*s�8�Oq�)� ����%�4ֈ%�0��?��\��;OJ˓�?q���?����?)���?iMI�|�:�Vj6��2խ��Fl�E/9a���.O�ܦc>�`�4�?a1.^'Mv�C�@��i28`�"[6⛦c�<$���?M�S`�d-l�<�d�<o���B�.̽	}�����<�V
�/J����H
�����Ov���/��E2�K��Vyps!�.$���D�O��$�O��H��&HҨl���'����o�Ayw�BiE( Շ�^[�O���'S7�Ŧ�H<i���0��e�H�%JЋ6K��<���W���0pa'u��M;(OR�ӄ�?�7��O�I�3��/�Ҹ��b� #�Ƅ"�N�O����O����O��}
��w^p���P f����E�5o`��!ۛ���	W���2�M[��w��0Ư�>�9#ժP%Xp �'\�7M��:�4v�I��4��$�!������jp���/��Րg��
+��"��/�$�<���?���?��?�b�\�lp�pB��,9��Ӗ��$Iæ1��BIџ�I�L�SG��'����?x�F�*� ��0yk���>�%�i+�7��f�i>����?ɪ�A^<����5���Ť{�R���LayR�ߪ�����2��'���$F����D��Q���Ba퇗1z��	ٟ�����i>=�'�6-�#�"�$ݓm�
E1���̚����e�?AfX���	���cڴD�&�#&�˥5i�h���X�v�1�۠�M�'6t4+U�%d�8�'L܆K%�O�4ט� F��tO�VPI���r�f�	ϟ��IɟD�I�����s����AQmR s��� ��C��)���?Q�Z4�v��e3剰�M�M>�".L�l���+5�qk� "M��)��'b�6����ӭM��oZD~REܾ
������V�s
��[>�I�����!P�|�^��	⟰�	�x�U�H�fji�0cK�u�"x;!�Zڟ��Izy¨a�ҡ�b��O����O�˧4�Ҽ�2�-<.��#�X� `��'l����{Ӵ%����?��HI"F��ru`�$	a�Y룪ѭq���U�=W�e�'�������&�|R�
�J^����%*�Բf�@+M�'���'����_��۴m�5�R� ��aL6��q��?1��k���d�F}��hӬ�1��7�	��e	�&�<X�L���޴D���ش�yb�'뺽*����?	�EU�4kv��4~��X���YV��``|�@�'��'���'B�'哈U��KRcX�x���	2ǈ� A��Yش}����?����䧽?Ѵ��yg�K�q�n�C'�G�:G0=�Q��,;�6mKͦ�I<ͧ����)&A�۴�y��G;=vȘÅD�71Ѽ4Y���-�y�̛\j<P��� �'k�Iȟ�	�W�)�b*��y�� �Z"�%��՟�IןĔ'R6���zV����O �d��XA�p@�Zj�"ǀj�lوr�<����Ms��x!�a�Z���m � �!P�@� �y��'�H
۩Mi��*�<����F�	ğ4)���B� �H�aĩx��D�&ߟT�Iğx�	���E���'��PRW�Ʋ�А0� ;2�	+��'�<6�\�_b˓hh�v�4��x�h�g�������"����O�7�E˦I�ߴ�^M��4�y��'��i����?�
d�9BZ4Q�#H�|@H����΄G=�'B�	ϟP��ßP�	۟���1vQ�i�aD	+t#�`5��-��ԗ'��7�4f���O��d5���O|�����a��".�q �$ �G�\}�n�b�l����|*����EL�S��l��+��P�
� ݂,{��wO������0
�����6���O�ʓ^���a�� 
w�E �.��7޵)��?!��?���|�+O\o�U����ɾ�^�ᑍu��e�7e֫D����	�M{��>�g�i7m�ɦ�@��]y��re�`w"� G+Է�,�l�<y��:�z���h����/O������=y��A?W'^(8�c��&���Jt>O���O���O����O>�?��G �'`��	Ck����A�bJ�Οx��ß��4~���)OL�ml��� ��V&�Aī��c��P(I>Q�4ś�OXYt�ih���O �0T�˥,�3r�ؑqK<�0U�ņi�L���$��O���?����?���xt<���x'`�Dʳh�4	���?).O�mZ7Lfl���<��B��8��p5��7f�@٥�����{}��~���l�5���|"��H����s��,	�8�*҄ũ}cE��	!�l�bjR������F���N���O��4�؏}EΩ*L��9����e��O���O���O1��˓,��&�I��r-X����St�s�d��_�%���'҅pӎ��q�O�AoZ<��Y��"��Z��P���W�&�,�A�4_��V�M��'1")V(xab���1^��I�=N��Ӻ%`���3�6�IHy��'r�'7��'�RU>��+s5R�h�%M"Mb����M#��¢�?Y��?�K~Γ[&��w�N��f��]�궧 
=	�@Ӄ�d��1l�����|2�'�ZD䕗�M��'��%A��֚5�,9�j<Q��ؚ'Kl�Z��S?�H>�(O2�d�O���)A�}����G*֕d���'��O"�d�OR�ľ<r�i�t�*��'���'�N�C�"%_~�;d�כZ�*ͫ��D�g}�HzӼ!n%�ēQh�H!�ȅO��0��'�;e���͓�?��_��fa
Ԉ��������iD�D�4@Z�ЀJY�
qx'�֜n����O����O^�d*ڧ�?�Ō;l������N��I��o��?IT�i��I�Y�d��4���y�CG�d���ӧG.H�X5H����yB��Ox6��립��k�ܦy͓�?Y��R�:]��	�M�? ��B�5%�.�@A��P	�y�F�9���<i���?1��?Q���?a�ē(X=���~�:@��X���D�Ħq��$Jhy��'K��e�W��C��]��%�536PT���tyb�'֛��:��O��$�OkҰB��[FH`���V�= ̳Mþq(gU�H�V������*��)-�uГ�IX�P�;��O�=��O\�9m��8$�H�s��ܢ�1D�lx�� $0]Ft�##گ�D����;�	�y��l�	�Lj�����G0W'T�8�j�1��`��K
�nk����e
C 8�di�	���H�'Z�E�RW�٧��3�P�5�U�;1v�A���w�&�ѳ� Ԃ-�@̇-,*H���'�\�a����T�"b�!%]���\�.���c���L��1�Q<�Rxl��Z��r��^��ڱ �!خ�Y�O����O��O����OUʴ��ON9	Bk�2F�m��Eьc5�A�q}��'��'.�*+���I|�CΆ^��̨�CL1|/������iכ��'��'���'����'�� �*9���W��hg@H�m�x�IAy2�OC}���d�
9��HJ��EҲ@́[�&E��Xt��؟H��>�`A�	`�Ip���ǌ�� b���v�l)D�զ��'�T�J�!i�\��?��'sJ�i�%�v��?h���c@N�k�Ҹ#A�r�,���OlI���O��$�O��?��T���:Q���&JМ��DL�~�D6-�&F�nZڟ�	�Ӗ����<I�'��N@*���? :�=����>R
�f(N0xW�'}��'��Oq"�'��F�\33���p��	
E%�=JRE ���	П4�ɸ ��ۯO�ʓ�?I�'�
]p�R>'¤��A�En�3�4�?����?�cBX�~��������۟H��I��	��F64���JR*�dK"o��*%�Ҧ�ē�?�����{�EEX������0Cv�@0�Uo}��Ѓo�[���	��t%?�0��A6�ZE���f�Y-�(Qj���}"�'0�'x2�'*f��%Ҁ=4��j�F��c�]JB]���I���Iuy��˽:>��U�~��ӎљ
Ш���LOK����?�����?���k��K��W?��Hbf��ԃ�㎎ah�u�gR���������~y��Bzx��?Ab&�'e�`�F� 0b��p�S�,���'�	ş`�'�f"�P>]�I�ϸ��s L>,P, � D�'����4�?a���?	���t��W?�	؟\��;>�$`R�jL�C����GI_/t.�9�O���<�@-���	�Ol���?!0F�V�WnR٨1@�CTx@�сs�J���OX�`��Ϧ��'lr�Ox��k$Ǳp�<��"ͭk\-x�#U���Iß`Q5K��I˟t�	Z�cr�C���e*L!i�-\+:�)�4s��Z��i`B�'f�OÖO�)�A��)"�ֺ~�V)�����mڥ)gzh��������h�m��W>���Nj�pił�%{J����ż�M��?�3�ཐ/O��I���# b��``�� =4���#��L�O�������./jQ�J�&I<���+�M�l�H���Gy��~��B�?���Xŀ��aQ�@5w�7��On@����ܟ��'v�C�P~D�!^�C��e� 6F��m�W�D�	����?)��?1��[(Z�$��G��l҄�V)g�4�ۈ�')��h����s"�_6S<�䒧�ϡ�6�������ڟ��?Y��?A���]}򊕘h�>��PbY�>@@%{�Oŧ�ē�?�/O��ŧ4��ʧ�?y�U��p	V�״ k�x���"2��F���O���ւ*� �O� s'��K|��*q,qi�#��I㟀�'` �bc(���O���Ƽ�#Lx�8ę��N�k�=`��x"Y�� #�ӟl'?=�'d�LJ�J�&`भ�7�$ �bL�'#"�U/y�R�'y��'��Z���07�n�S��N;�(x��P�<�`7��O���G�\��b?ɐw�1,�!0�=)8�ȉ'IxӚq3�P���IΟX�I�?��N<�'J݂���_�W't�SCڭN\4����i8H�'P��'R�O��s������+d�̴��h�
_����rΟ�&z0��'�ʼ�2y`0���b� _�ݙ��Fv"
���3W�lx)D������6e5'I�uJ��T�@����vo��2��9K���ŉ���м��g�)�OO/'L�+�䝱?)�l�숎,A��Q2C��Te��[�a���hS�_3<h�皿+� ��.�7������,�5y�#�y0�	�"�0��	ޟD�	ڟ`���ɟ��I�|��dЍ?Sp$���� p��#��\�d�ް��ݟ��%�Q�\�Bp��DV�N�X�f�JQm�����PXt1c��~\��bG@8n����Ǔ<�u�	��M�G�4<�M�0��<V���DbҼby���dZ^��yB�(���n�y_��"�y�b٪@"t2fa�<6��f��y��>9+O6HC�d���M�Iߟ��O�
p�CD�:e�MkƇܥps��▊B�2��'2��_�� �[C�24`�kT�K�$��O�jY��܁t�vi��� �lo�4Î�D�]���Yb
=�6c��;iT�'!NB���)X6ɂš�	@�HGy�a���?���䧡?9b�rV8�y��KL���r����?����9O0��6k@$^АYsV-<(S$`�'�O~]�)�|T��*�?q4�#�<ON�[�Mզ	�I��<�O�X5�'���'��d�Ȇ�d>�٥,�"����H�=�l H��{�^�ԧ��'��O� ����ԭ$ܜ�3�L3E>܃&K[)���:�/�&#��J�O?�H�$R *�q�x��5�	����i"��OZb�"~�	*hu�l�g��}<��,&C�5J��H�����1.}����v�2"<�$�)*G!OV=�+*�����K�<ivG�Q�|DK�G"J�����`�<1�HXc�ԑr2큞8����Y_�<��fW���������kB*��\�<���ڂ4�!�D�iB����D�W�<qfd9qH��R�P��=�F!�L�<��:�P�Gg��S���`��G�<a�G�J� XA@�^�^A����G�<�V$�8iF8u���GCT�`#$�]h�<�GOO?��< �J
�\V +��a�<1��ۀX� @:�.۴e������`�<�6�ҟLt�k#�
e��X`�r�<)DLK0[Q�=�qB�{�RdrQ��j�<�^XS �D-fuz����>u�h�ȓa���z�Ʈ+���	��&\lΡ��u^�d�S�ͧ>6� �Ӌ��~p��0_��*�Eǲe��p��]�5����%��F�3F,^�]¹�ȓ(��cE��,)����1�B':��ȓ'�
)Y�%ٯnL��PB�~$�ȓ�U`�.��<����8�"O�q�F/�X��)P�T�����"O,��Ӄ��F��I�&Ne��9��"O��â˘,<��waA�i����"O���"ۍ	��̉A'�XJ��h�"O �,E���i`�"5y(�i���y�aJ& �� ��`�3% �Cdc��y��W��ճ�>~��E��y�"ݏj2J��0ꋦfFN%�b���yr�'Z3ZQ�gƣfK�@rE �yr��3{�(�JT
�Z�����y��ɑ{�H�{��E�Q�=��ԙ�yg�0H��Òk6D�$��3a���yR�)H�HsS�^�5����w�ؓ�yBf��v<��V#L�`�lI��O�yRN�AK8�����Q=bܺ7mT��yBgR
$p�XQ�fF�P&��ö����y�eŖ�R��s`X-=�0Yj&�R�yi�J��4�P$Ω+'��K! �yb�&���(Z���Ӂ����y����mx�t�%�PC���F]��yH�8�84�-��ҽ��c��y�
�zx+�.�-?F��#f�y"jK8�x���	�2�y�֎�y���w\p�E-ājy
�Z�L� �y@^�6x���"�4��������y��ԑp���Q��%e�@�J�y2�W����-�T�\�3�kD:�yR�A�\}B��3M-�ݙ���y�e��	�g�I�H"���Pl���y��0V��)Qh��>ּ �"��yr���$N=A5ِ0Z:��r�K!�yB"�75P�ȴ��!�@4�2`�7�ybW�W3�u��n�R��R/��'F(SR�2S8ҽD��-�Lx�z���3*�����y�n�)��"� ������k5yl����B��	�]T�"|�'���"o�?�rq��A�  Te��'Ѹ���� �)�ȟ�����Q���uP�1�{��0�>�!���B�AYvIP��p=񷌀�Ж\P.F؟D����Ĉz%.�9-�����.(D�� \�0���<����@�F2
b�S���VD�b�Q��E)i.�}��l���(!$&����d��	XC�<�3��0h�F�"dI�Ϯi��g��~s��rc��򄞾%
>�snm"e�ܙYv�͛�`�Ʈ,�ȓ,Df����ވG��)@'� ���Bl�<L;�z��"��='I '2a�DÞ[I��FG�gX��9օ�`�)+>�� �C���&l�A�N&�y"�]00��ގf��<+�ֺ�HO�\ ����h�V�SR��C���3��B6ȣ�"O����y�~��K]�q��ȁP�iS"��%'�o�S��M����Tas"X�i^�qS��h�<�c&�!WlQ���ܼFx�D��Pv��}���i��Q���V`OR]QC�
��z��R� lOh\C�hI��J'�АRi���/С	A�(�B�Ԧ[%�Y)I��S
�.�$d+j��_�f�hDO)�~T�>QEB�_պ]���P�5�~�����'�j��	:S�t�� ���M�x��	�'�L���t�vT�0�x�\%Kp��$X<BsfW�N���	bӼ`@��Y�)I����^>�$���"�;&R�{Q��[؟8y�CO�P���+e�G�"`��Ytd���1�4P���	R ��Q�k� qf0 S�F�@��!ӷ�8��է'{�Y�S͹��0���QmQ�|x�o��y5Н�����A��ю�O^؈���{��8`��Kݺ�`앭��'�.��)7�J���<i��P�vi""N
j�0�NSW?i��X3Q�9RT#�95��Rs�H?��̙�:�L��ҩ��S���K��!�� �n��>}�Pڒ�&4���&,G:)..�!��b�~�#�DE�(Br����z?A��jZE�/�$wWP���A��s�:���"P�ADj���o_�_�����'=�m cL
(M",H�(�<V8�D:A-�8#L�@q� ʒD��b�gE�3TB�1�$G�"-J� ���E8M>����=h/�R�e�u�S�_v�'�݁���e�*IRb`@7|��d��0�Z�� �X9P^$���M�%�$7�E8kR
� �Iʋ=�XQϓ"���+D��.8���G�2��'�z��q�ɷ�Z�+��H�/��|�O>��צT�'
}f���wdT�1�N�)Uʠ�C�:�JB�ɎN�<L3b� ݢ�{��"q���`��cV�	��%�[?�1b_�&��t�)����g͌f�����:#`drc�x�<Q�I�D��E��;�޹��dE�!K�lٲH����72�I��D��[�)��p�Ç�	���1QF�_v쑆�	t�ʩ��Þ���f�Y�8��_2;w���*A�;6����+)4��S�ăC� U�X�p�O� )�	�{�Rizq�4�']��
���_�f!j�l���q�Z�!P M�j��2 ��l�MlZ+{�
�+R��s�h5*��֒g̾|�e�n#6�I`"O���)Ki�=���&����^�H�T�ɸ05�{B�P�"IV�R�z���K��G�>��(��v\��$F�D?PcW��@�CF@֚a9!�Jr=�=;�]}0)�Ta^:*ב�P�R-�^K�>�t@
9D<�ȅ�T�[�9�);D���sI*P�2�ҤӦi�j�r`�e�.hA�E��������چaD��suo�*-\x-��cV;�y�kM9^L���hrI��Ί���d�x�D��-+B!��F]�V�`	1���Y��u��I9G2n���'$n���@�2�0�aX/.'Θ�'
A�2dA�=y\��#-��r���2��䅩L y��	$?EjH(3�3I��PN�rg!� n2ܱ`�N��ꐓ_���]�{�LX�=E�ܴh�&�ց׌#s|`�%N՝*?�����كN�x_|���ޱ*��(�'<�|���'����׫wO�m�1D�c�����'L2ء��o�l���)��S�'Y�!ÑdP<�$����wm��y��Ip�%;�Q█b`��!�yҮ7�D���J9L� q;��,�y�\LLEZ���K*�pL�/�y�ĈA��rԩ��N@���f)�y�˶Jtd ��M;I��10#0�yR�H&B�&�)��>�^�4�y�]<�
��a��f9`���޳�y
� �(yta�Ml���L#l�m��"O@�ѲaB7AR��BCI]�¡�"O���7Μ7����+խ�t�2V"O�y�.�A3` ۖL���݋s"O,�����	(q�ņ�Ȍ9"OH}z�A����h+�� |�8��"O��`ή1���Y�d�Z� tP�"O�\۳��e̼P��@ج��A��"O��g!��9�RAW��� ��1�"O�����"bBh	�-�
u��a��"Of����� �/a�Nm�"O@d�ꚝm�H0ӥ䋸%z\h��"OVH	T��.'w���D �JF6�Q"ORܢQU�H� �H8���"Oh@��ү~�*%&�-!R���"O��W̋�,o6�Y�,��	d"Ol(�/��Z�tIժL�H�=��"O�ݓ�䔡O+\�D�� �$��y� �����[�6>.8(�KG�yR03��$*����'��[�	ޡ�y⢜�s�`*-���n�0Č,�y���xEK���J̘Ӧ���y"'��w�T���)�$����<�yr��*K�\�H�2i)"o�:�y�ʭN�*���<R)�L]&�y���m�R���>�P��h��y����_> �Y�V
�(чل�y��CKl$I4!�~���4�y<a�y�&�&8�9����y���'���QK(`����U��y"�޵��m����/h^�tٶh[��y�-�|�6�KW늓*�p��P&���yb���Q� ��-��R���'�y䆹-B�yӐ�M .r�(d԰�yG_+6����G��~9 
$�C��y���:c��NH>he���y�f��#�Ip�m�,����y�B��VMīW�C�f�aÀ���yR�$ֈ� K��;ʞD�RB�9�y�n	�ʬr���!=*�#�(_��y"�L�\�`�A�$�fU�D���y��
7(���BQ+{�zQ��:�y�H��[]����]��Xk�=�y�ǀ� ���P'[?$��� q�Q�y�C@+	�5��K-kMZ5�͟%�y2!����)��K�K~������y�&�JV���B]���q����yZP� �D��t!"T)���"C�Ɂb9��xS	G��ݣ�v�$C��64����Λm����s�f��C�I�R�rm{pN�W&��ifi�	<"C�	� �P@�g�D+1`ŋ4�{UC䉦P��С���DYn�?V;�C�	�x��I	6�� TI�u�P�~èC�	#Z��a�M�H7��� ǟ:z��C�f�E:�+�L�!I�_QC�C�	�r �L�`�X<�,(�C��7:82���@�.�F����6zC�I=X�hF@�*h��6�V�j{2C䉍`d怣PjJ�)����G�7^C�I�t�� b©F#�i%F�O��C�I���c��.����DY+ǂC䉋]
�bD�Ǧ[�~Io�3Sw���ȓdl]��&�<&�yg��6f�H��S�? �C�mH�B��{��q"OI��`T�2��Lp�"O�a�'�� �r�ل@�T�V�S$"O�����B��
E^� �"O��ឥ_A`a���P��<��"O�Q"_�M�!����:�&��"Oҩ	g��J�05�P/��h�"O�TU�ا$H�:���l�ĵ��"O�����о3��ſw�\D�"O8Ա�hK5�
�&��L����"O>:w�J�sXr�EɧcX-�"O���eoL�:Pes��Te�C�"O~X����!l�촩f��;F��g"Ot�+�N
�HRm ����Y80Xҗ"O�!�"�O*���sr�R,Na��"OݓTK�BT����˜ �A3�"O>��QKP;<4,��ᒖ�X�"Oh���ÒH/ ��P ��v<ͺ�"O΅X�A�s/.��#NJ�2H���"O�����a<r�,W�5��c"OH��䎣|�(�;�I��0Jh�"O2�j�,_<A�z00�G	cW��p"OH��e�9]ʄ��V��[4R ;�"O�(Ś�eV4�(�Ћ#�Ft��"O�t���*0VY��蕤ɘ �b"O(����҇nl>����X�b�T��"O��(û)|.\	�,��	�j0��"O��A�腰L{�D)UkQ�`�c�"Ol��*�3
��`�	E�T`��"O��SGB�ma��S�G%�U%"O`�X���KP@�����/0x��G"O���p�J�@��FB�]v�"O����dޥ7��ᅌW�ez
�@"OR�el��d`�X�ą(uU�t"O�逕杵t�Nl�"�6qY�s�"Ov��p��r�vpd.ƄlV�] �"Of5�O���}��.�9��"O�{���~�Tl�����q�"O��Wj�/4u8�B��b�K7"O����Ȫ��y�S�g����'"OI��U�n6&� �=u����s"O�)1�ω'A��I���^�0ؓ�"O��Y�d��]{��rn�	�`i�"OVt*�ˋ*�P�mW�Q
�� �"O�s񣃒b/�Ål��Sb�q�"O�����n���Q�LlAn�V"O E�udԞ~2ȀG�w"$D`�"O�����<q�xcDmXsx(�"O�01���6���d��lb�Cw"O�(�#�"e T�`oY7EX��r�"O^����ҖBRHre�I.�0h��"OL���8����E��tk^iKu"O&��Ƈp�m҃�
����"OЁ�p<]l�ԓG��f��9�"O�J� ԟ4��[A�"~ŔXA�"OV�Ar��=;�U��1W
�͋U"O�x�����r̆!���;Ljd��"O��e�	<���AAŸP��E��"O��ۺG���q���6�B�8d"O�$r@�ѻ^��`��Fz�
#"O$�"ed�-~��bD���d~��"OΈC��\ jnh�C'ׁ;��u��"O��V��(i:-��ƀ�|%���`"O��c��O/c��r��;j��Bw"O� *�j�E)��xDS**�ٓ"O�\k��30+�Z��W��h��"Ob ����
ir��Y�6���"O�P��g�*^<�D�=P�p� R"ON�і�߱LAZ�ȕ:\s��y�"O8}EK�U�M(Gk��"O>��6㝸'.�V��HS�H�"Oꀀ�kUM�ipb�rƝC""OX4��r���i�b�(NS�� 	�'�p�� �ʦJ�$Ո���:W[Ą)�'���[�ˎ���1�B�NU�Ir�'p,����_�hse�M�K��@*�'������Q\ ���сm�����'V�i�#�w/��0�L%̴���'bd�aĝ�c�R����Ŏ �U�
�'_�4Yf�o ޥ����.%�e��'���nT�*f`( �� sJ��;�'�aᦩ�� fm���d�✈�'Vt����);�j�H�%����'M�U��a�'.���&iS��4)��'E�H�GHh�q��J���6Eh�'�@s5�ҿ%� ��&N�uZ����'���$�	BJ5Q�h�'�l��'�1c��;�i�V��Cn�ӓ��'��(7C�0:�jٸe�6\!Y
�'�.9�F�,Np���&���P�'�h$�a$CFl�l�7J]�u��(��'���	���$>�B$��,>����	�'������`���N_�NXy�	�'w쐰S�BBԀ��o�.����O�왕��`�$_'uFn���"O��qR́1=.�84dY�\��z�"O��K%5Dv<�EH���� R"O �B���?<ÄHH���v3�=�4"O����$ޮ
�	���Iq24�#�"O�T���S;?��E[ŀM/w0�l�d"O��h�� ������4J�J�"O����<F��ER���]f��"O��u)�%!vq)��F����!"OJ 4HܕC��@(4/H/I�@%��"O8h�6�׉0�(�0�N��y���� "O���΄�N�{f$��B�XX�b"Oި` �u3<pCp�F
�0�a#"O.X�U��(͈�`?
h2���>A
�CPbE��f���e�F��A�r݆ȓ07r�A�)�]���Y�*�	�"\�ȓ'�����	p�)�MJW�V|�ȓ=��uaU��t�#��9��1��;k��GE��H�\���x^Ty��b��Rf��(��u�k`~���7@�,Sd[7������?t��(��P;!a �ǚU�.yDÔ�BF�� ������)���ĉ�t��WRv@gŃ��d{BeQ�'�-�ȓb�KE@���֪q_���y�@�NΈ�!���S�`h���Í�y��ʠ<�
�p�J�A�4����y�F�:/�^\h�ئ©@K/�y��Z�{����@j�|l���yb' N�E��{Ҕ����:�PyR�	&S���R�dn�pƧ\A�<I����!0��?g���XƊt�<�P�L01E��xR��V�����Hr�<i���+��r�KQ�{Zn�"�h�m�<� Zu��� m|�5�ԃ$3��\(�"O��G�� ��]���4^��=��"OM��*K<
x��aU�S�Tq�s"O��C�.(�V�Q�+�����"O���E�z��x!`Ȉ1�t��"OH`
��us��3��tm�� 5"Oqj%Jڛt�l�)�*R�{:�䣧"O�]yw'�":!�\d��/.Yb}�"O�2�->dz�i�4b�l�"OHY7 }�Rm`i�"�����"O�0RG\�Y Z͐�CBJ�m��"O��؅V�yr �r�8;+ᚒ"O<��`]M��` ݫ%^� "O��s6AS ���r��	:�1"O1�E(ѐ�2��$d4��s�"O*��3(ڒ^�B�x��q��_��y¥���L����i|�P�͉�y2
 f�%� ��X�$s�� �yD��(�
pxą
:�X��Y��yR	��*��p
�c[�	�<���yR�)8��1T���+�0%Z�,E�y�(S.ϤdP�'O<veH����]�yb���B ��8�ɀ+qh�� ����yR&U�a�p,˷�͸Ln\/�y�.֎K��b�h1Nؠ#tmԳ�y�."�u��'T�!E�a��5�y�B �QE0��Ą1!��@�;�yBkL<"Җy��F�rT��G���y��Z']���2)����#���y���)���󀀿�D�(�n֝�y�E�J��i�������Y�y� б��(�uC�$�Duy��	��yr���D-a��єLz�ݲ�#(�y�JɎH^,\X!��<��<+����y�EN�3��/Q�-:������4�y��1����dF�3$�}1�<�y�(�]�0�j͡`Z�H35�I �y��)K��U��,Yb�b���y���b�˴��O"�ġ���1�y�	�3C����Ą�J�%�R�Ȱ�y�+�A�<�����::��)ǀ�
�y��̝i�̜�&U�H�����\��y���B��QR���o�؉X E���ybŉ'�
���� 'dĺP����yr��6¼�뇁עW�V(H�a��y"C7By���q��6Y��uK��Ņ�y�S�7�V`Y��A�LISw@I?�y���@1��ȁ�69�	P�HT2�y����Ґ{�eL�vE�?�y"K�_��Y�CK���rqp ����y��S;�~�Pte��w���2�-�
�y��YO���k��R�D� ��&O��yr��{߈  �nR2;?��)����y�Vj��Y�k�3����mĤ�yr`]�a�4��< t 2��y��E�$$�w`�&���I�yҥ	.\�����z�tT���yi�@�S!L��'uܝ��F��yREس�p:JV����I���y2B�m����'�4���$���yr��0/ �{O�j-�8#��9�y" �!n�Q�I�*hT��!��R�y��|����,�M��DjX��y��f
�۳�O�O|�وt� >�y
� ���3'���i�&Zt�$ v"O�m;E`�0g���P�=:��("�"O4�*��d�^���ăRS
�E"OD<�.��8��a�Lt0��T�<AЎD(~.Ź�3@ ��
�Q�<qdnթ�!z0H
/W!������V�<qR�;P����l�g�<A4(G6n�|c�Gӓ�j�u��l�<q%hș��-��ܦ��EQ�Qs�<a�K�Eh��Z�&��k"����W�<����Q�a��D
Q�1d��J�<��c7ms:�K$�("�,1B�JE�<1�"J9*q��j�#(&B�H�l�G�<���6D�48�vjRIܒ���#NF�<a�N��Lsd�H���:h`pQ+��<iE�b���a�lN��K�b�f�<��n��D~Z�(��ŵR�"��A�a�<��-q7&a�DW�d����g�w�<���U�j��B�6�4��F�h�<aT,�W���q�E��5����y�<y��Vn|JE@$iȹj�V����x�<a�-Q?=��k�B�?�,)�d�w�<����(؆���*X<1%N\��l�<I��FTn�XzdJ�8�l�p�@@�<I��Z�JlXI^�b�p�}�<���K/B
�yF�M�,^�u�uÝO�<A�ɛ�LXūQAlJv}�7JXJ�<Y�#j��RPpC��A��G�<ARaD�lQV�!aT�M&�t"�`HE�<�b蓘o\D�+��T��"�&�C�<��[=gˈ�儒35>�f�x�<Y���>*�q�c�':�{�ii�<�tǖ�{(�h;���A���ӭ b�<�6 
 T��@������@m�a�<�4�ɱX����2DԐzf/a�<�.���i���ܞ:d��PG�[�<�᥈>�V�Dg�0���7/�\�<Ia��=;�����\T	��0�(�|�<��֥^)�R��$�؀��Oy�<y#�^*z���d��D88PT��u�<Yuf�8 "l i����$0x��G�<9���n��A�J�8`���^�<�r���=<6�@�B�6d�	�mFW�<Y��-7����˻`�ʉ��]O�<!�� 0Q�U��M�8;f��b��L�<)&$�=�z�ۇ�*u2^4c`#LF�<i�B�q����-K��D äh�D�<i����7g�x�%,׉_����G@�<���۶/Ct��B́�ZQ�Q�7�GW�<	�L*k��m�F/�e��)P�T�<��ӎ�v�aq���Ƭq �v�<!��N�=�����79Φl�.J�<Y�)1����[�y��!QWH�<Q�LG�pM�q�(D�N�_�<��C��J�L�9cNˢ)<����r�<RMF�w������Z�Z��W��r�<�pkE����Lː�BDڥ�Z�<Y6� �<_�����=J�u ��YT�<A�,�� ��P��@Z!"�����eR{�<�!!�`�D��S!�r�<l�d��y�<�ҍ�_r�6��z�ިAF�a�<��l�u�ș�-ōM�E��O�h�<��쐾o=�4� H���S	�M�<�d�6*��H1셅�,�̈́`�<� 0L���ЗZ5��C@C8$�h��"Ou��D��T� ����4��Æ�^�<၌�J�nq`UG�>����_�<A���Ŵ�b �Đ<�*(e�W�<���	z�Yr�-�5h1��h�V�<q再/0P5�G�	X�4q�3��g�<���AϤ����Y��т�f�c�<�q-@�J9{Po��7�����k�<�4/�<CJ�A�a[�n�X���&�g�<����w�nI�CO�IL�*W,	L�<�$KB,H@�D�]4'U��Ba�<Ƀ��97jʰ`%ШTl�B,_H�<�����d��x��$��1��Yy�<)wh)0z�4����	B!ڴ	�)�o�<!r�[c�mR�K�;�ai�"�S�<�2(S%L�KӮ2��w��V�<V�ͫq �)@�N�d�����CH�<ye$Rx�Uk��
8 Z�Hd*Y�<A
oa�/��q����T�A�$q���{ȴ�I�$ˎ���KV�X�n�.M��iֵ𐄐�GJ��7��5U���ȓS;M���I�lTL;��� �:���-�T�PR!;n?����l,K<�,�ȓ\��=IR�^$sF��Wj��LVL�� ��(R戠��q"Š5�q��J\�ej2-�:d��OɁ	�ԇȓjr�(r�%�=�Z򇋇{�H�ȓD��l	�B�0>�ة��L���NL����u�Ѕ�G�, <�������q�R'4� 1	ƫU+0t�-��"�8 ��)9 �u�!��Eb�'>�@��F�S�H��Q@I^|���
�'���Jʝ~�
 a��?hFp`�'P�E�1%�7.F�[�œ9�E�'D6��ec�?\
����K�)�����'!.!j��]'M��Mۧ5
Vp�
�'�(��ѫ� 3�> a4��=6``a
�'��;���}(���ˌDy�ٸ	�'fn�	�&�y"8�JQ+�>�ʘ�	�'3��"��4d\H����ȓP%�-JBER�E���rGE@����]�R�b�"K"�\س�ļM�,܆ȓ"q���Ð(8�u�V��!1�e�ȓ{��u�����T����H氅�}�����żrt��B7>������d�Έ�j�i��]'Fn�ȓd����KN�����iZ�]sH��+��B�,b�@���8���ȓL�@��#!�b0���7h<���\y���A4�����2g@HI��#]��#ϗ.�8��A�(bx���}�����!�9;�%��F��m�H	�ȓ/�ZlRT�ѲZz���C�?���ȓSV`�q�%B�aԈ��EJN�%j��Fh��O���'�P,<��]�ȓ�ؔK��4�D�ӕ�̦|Z�Ԅ��j)�a���	��i�"���h|M���Ԓ!W~A�1��Z�@`�ȓ�(�Yb����T��ȷ_�t`�����cG*G])�C޻E�@8�ȓR(pP]y��(cQT�2ئ$��"O �Ic�I�e�Mh�!�!M�ʹ�f"Oذ�6W�����֋3{�d��\�<A�KJ�3�hi@(�]���J���B�<� n�#e�J#:�^ �i�w��5q�"O��I�`.���w����䐓"O1�m\�cޢ�1'_1d��dQ%"O�Lk�'�59:45jwK@m�"O2����r$���f�� f�h`�"O�9)rN�c�(�:p� {ʥ��"O�a�!�4��šp%�"+`���"Ob��C��Xa���s�7�b���'�(��!�5�Xa`0%T+�J���'��e���#�x�K�Qh���'��+�`�i��2ք��'�|��ubZvA�tX��A!��\��'�`["��xt��D	�ܚ��'f,�ch�7@m�V�(�bT��+��= ��G'H�mA4�	�ȓz�����-ѷ9\2���&����|��@a��>-Tj��w(���i���CX1�Z@��o��@���ȓB="M�s�'&$��`&$�%����ȓI{�@���$�]PC��ä���%��"lڽ1���Ɔ�P^Շȓ,�1!g"̺[�&h� �"O��ȓ>R��W��$r�BA���%#�4H��!�8Ê:v�@��Ս^Ϯ�ȓ2É�Z^��Wg5��a��v,�!!�u��v&�>:��ȓ@����P�ȕ:�~�2��G:p#̵��*�Z`{���W�$��+�4z�"��r���Ru`Fk[xDBh9=�Їȓ3�R4�FBǺ�E��gӴc��̇� 1������7R�5lU%F0���l��̰��@$�"��$`�����oQ�q�d����!uE������D�d����l�j��3 �3e�LՅȓ�2P�u`�	t�|9�)̭iKȘ�ȓ �<�d�^������,(>���e�s�+�1S�Xq�C�)�Ć�QX�Qr�7S��0�B��B����ȓfR �f�W-3ޘ 1�T�=��ԄȓpŊ�0���Z� ��<l��̄ȓh��<XB�5�]2�H�Y9��ȓ,r*i�ghly��] 1�,d���� X�>pH���ǿT������{�,$"!ZR��;/�r=�ȓ��0�K�^�NL3�(ǾM�p��ȓ+_�����i�t��a\?|�m�����B��P�pd:� ��v��نȓ"_�u#��Q�F��\�;�R��	v�������.���� �L]d4�-�;D�}��<D�p�H�eR]B��K';	8�q��/D�P����'ZR�����\7I0����+D�4R���xpnEX�+V�m�9��)$D�D�򢔀4t�
�\� Ai4-/D�lc��LE.��fO^�3�����,D�`�V$'pd+��9,E��Q�?D��D,P�
�ɫ6B*
t� C#c?D���獢1�mф�@,^����<D� �4C�/6��� C߽#�:���9D����LØ2��g&_FP��+D�d�0%��O"�Q�°$�N��D*D����U+&�@�+�ø+D�z�h2D��@!#E	\��9h����D��i�O@�=E���&&K�0�B)��\4�e�R�,n!���[��z#� �y�Æ!;P!�� ��Y�~�<uǚ4pY^��"OtX�V��
7ܞ�a�����"OE(҆�-��Q���ļF}JT�e"O��#�R�3�n�"6|��
�"O�H8�����Xx�MHSqfi[��d�O���Oj�;w��J���HE
^�*��)��'�f���o��'R�;Uo��z���'���vNȝM�f`�A�ϝw>l�B�'��ҍ�~@����}'���'��ybEAV�0���*�v�r��'l�lR���<E<��۠=F�8�'�l1���I���H�� ȄʓB���`u��u�fZ2)�A��ȓ� )�S_ N?2(��н]�bH�ȓ.��-��
Y�*�hѓ"U�I��`��w)��
'.ƕDڬ	�#��}�X\��e��c��ͣ~�$|pփ�)C�����!��!�Q�ld8�b�*H��'����ԔȠ�ϔr< ��"�4؉�EK�"�I��T�Q�Xi��:��o��8�ұ$%�@���v��%�@�L�~�J�z�W5�F���G�Z8�ǩ��_r�
҅	'o�9�ȓy�ع��,q��)�ACT�Н��FN^��$����Kw'�G�ńȓzLnMI���-+���E�T�9�*��ȓ+/ u+A�L�_�̱�MƎ%,B��(�����#ƫLR�1�JF
6�0y�ȓh�ɒCU�3��pѠcɜt|d�ȓ-���!��T�P:|�6��(��`�ȓ����݊a�RZ�KYT�d��ȓ5�d*D�H^d��ɲ�#F�rp��/��Mң���X,yA�X�F�h��!���Gɋ&r@��x!"\08a*Y��af������<Ft�H�c�*nN��ȓR���E�4%Cf ���>K�4���3&hy���	�c���ӀO�;gH���ȓo�X�9S�БOs���զ�7s�4�ȓ�*PbG���OCL ��O�/O�>��[8���5�b ���.t�61�ȓ?N8=�P�S4(�ڔ)���&)� ��-�09�`/R�Zd��OH�Rt�Ȅȓ3�P�Q�`��n[�$r4GҊw��l��V͖�9���%(�pm�.R@���ȓ�(���۳_fB�i�CX�ZR���i�����טPÎU��<�Ե��/֩�Vb��6e԰i2jF�%���,��+0'�'wV&��t��P �8�� >%9��ɿ/�0��M��5�ȓT8��r��';��p���cq�]���r\�`�_1I@H��I܁p��ȓCӰ��rLI;F*�s�&A?yVv=�ȓ�⭃�K%P�Fh3H��(�ȓC�|��$��!h�-��dQoR�!�?9���0|
֠R	3����G.!�H!���d�<����K� x�4Ę�r�DXaHa�<��	1o�4	1�b��*�[�<I�쎀e8�m�T"D�F^bh�L�<1A@�1)����#u���(7�P�<y�*�^������S�
�8��[W�<i����>�|��X�u������m�<��%\�J!�Th�"��� ����g�<��ģ,�, ��l�	2@ +w�]e�<�Ύ�kT�(F�ֶW����BCEd�<� ���ĕ!%@�h��J�q"O pAPf�o�J��P�!s��0��"O�ݻQ	�e����m�x�c"O2P�[6~-6��cϜ-O�� x��$�O���IB�+�
� ƕ�v� �X�aȋqў���I�+(6Qi�E	�:ؙ�l­w]B�IX�D�KEN̋} ��P�E�1"2C�	�K\1�rO��hXN���l�<47C�ɪEEr8�ǃҋq�,* �R�B�ɷ^k���$K*d���J_����$h�P��f�.1 4��$D�)�t��'&)D�(�f=R�|��%��g�(�4n(D���t�:WF,�aw.^�
$�(�E!"D���r�TyG��`�%юyK~@h�B>D��	h����Q5R��K D��2�J/��aJ�P.t�t��g�0D��!�I7s��PǪ1Kz��/.4�x��Z3(�$��9	�����ψ|y��'��83�.i��a�FĔD�FHH>I�
tC�O�z�V�ZP�òY��X�ȓjɖ��p�O�D�4-Rd̗�~ނD���"�z���vp!:A�"Fв$��AIEK��kr�ꏢG�Ω�ȓO�f����?����MJ�!-�=�ȓB���)Q�+B�Eт�	�hh��7<�h��C�>���!$��bٕ'�a~b J(�4�^�����%�K��yb�E�'����,�X��� �!Ƅ�y��FD\q�߃}z�A�'�5�y��Υ���G�6f�\]b#�'�y2�~n��;)U2�� R��5��x�V?z�� �#Z$�("F�V w!򤚧zh`a[�j�-%V�E��MS!�$O"S���e�*h��%`TJZ?!򄞂<6{���8}N��FI>X%!�E�m��L+�  �(�V����A�!�d�-!`T��V�=/ڬ�1��
�!�dD�l2�����X-�\J��n�!�Ę<Z��}����;��S@����!�H�xX��)'�_^*�k�B]>�'a|�!�2�	�B���ta���C�y��firAk�,Y4��`V�3A�����2U���ȈDp��#��2<(�%�ȓV �@e|o2e�b�+NZ����}K����:b0�;���*"݆�Bs��2�2�b���lI?��5E{2�'}Hq���"ŜQB�&ɶ&錐i
�'�r�Y��u9�	Bo�H@��	�'h@�5��7\��A2��F_��I�'�6������^)80�7C�<KHb)a�'�L�G�Cz���V�š7���P�'$b��ˋ*k�"!3����0�ȓ�(���̔�_���Pk@�6!�M���g~"�E0��]����8G2\������y�#��^dɁ�P�A��qS�;�y2���J5(i�H�#���y��č�y2ⓞ)V��3��Уl}̵{D���y���g�\��]�9�S�^�y2�L90���YS��]�b�s�I�!�y� P�f��$IfU�0�7�y��2n$f��*	�����ꘕ�y��N�4U^����*����V�y�e
)W��!*2+$�L
w��5�y2�K$Fh��R�#'�𐖠��y
� <�i�f	�����S��}�"O�ʅ�^\Y ��BjR��ܸ��"Of�1GO��V3*�0G��-t+����"O����l١�(H��Z��"O<āGA�$Қd��C�h��"O�=0�G�x��A�U�Ț��Q�"O�l9��'E��P��n�L��졤"O6�I��);�O�	ƌ��"Oz�ە@O薌I mηP���E"O&H	�
<u� =�a��$4�؁y�"OL��u��>�n
����HC�'��Q��Y�lA&C#�T�C�'����	�+�<h� �ن�p�J�'8�"V��',|���k��?�Y��'�p�iVn��3#�U��c�;}@�r�'�$���ʠDSB,3��i{	�'jN�̏-;9��0�mK((qx$q(O��OZ�}��0�����,h�V	�0�
� �vm��~R>�C�֘[�n��%�E�5��i�ȓ��WH 5���x��4 7 L�ȓb�p�kaF�W~�`A�%6�ؠ�ȓ^�zYi�P�.��$��F9W߈X�ȓ�r�t��Q}¬�U���ȓ@�D��'�S&4�TMIV�ͅy�����|����z��# �|�@IAL�
�<�3�8D�0C�;>�:���� 3LLu"��!D��R��%CW�y�aO�"g��)�&%D���F 9ig����М�,u"��?D�\���ڷF��PY�G�%n�b99+?D�dK��!`�S�MO�3�P�<��Vy��58fFE�2�ҒUݲ���(	�˓���h��d����%�ʎvevP���K3�!�&!�T�� ���Qba괧�&�!���K�>�[�ށ�l�b��R�!򄖉}vޠU�3>�p 
�e�2k�!��R����d-N�5δ��E_:Kp!�$�q'.��E��� �T<c%�H~4�O����|
�O7�H�gl����Okux1�	�'*H|� Ɛ�j(�%�>s��A"
�'8�q�������T���d����	�'qt��e�\�N��Q���Z	�'�������z�3�o P���'�
D+���Xn�a�PH�y��er�'14��G�^;\N��w�FgD��[��'����|:P���<AހI��>'#�0�t�YV�<���4f��kd˼Q��¡)�{�<����96pMb'�ܶ�J��db�a�<��c�gb��(1-b���֍a�<���
�%� �It�S�|{�$Z���E�<���I�Lø�1��V!:�)��\�<a��^+Y��W�&XZ�Ы���X����$2�
S4�'	�*IwA�A)�v����L�H9���ߍ~Tb��v�4I����족�˙',�e��/Hz�u�ȓiU*y����P�b��,��v;Q$/r�A+�.5Qsv��v�`-�2L��1xz��f��<{j	�ȓPa�� @�	<؂�
f/5Hp6��wwr��-� �N�ʑ�J Dx��	{~r/��FF��.֬z�b,�Eg���y��� *)R�["Z�m�}�u��yb�޻#�L5���ߢ<�"���Ԅ�y�h�)��X9 �K	0�@ѣ�T��y�@�L���K+��<��^��y
� T���D]D=�� �r��D"O�r���:R
�q�N�O�8EQ'�P���pO״�8��ݫZVP(U�"D���#@�=5"��P�`	t�*��Ӌ%D���3�I�yn���#�9v�u�1D��x��ޑO� |�F�\�Wn$��e�;D�Xx���'_[�y�CN�q��AIt�.D�,y��L+XB=#�M־�� pv�,D�p�ć&-������T��`�!+D�|�W�S�(��,�rL�+�\\AF*6D��`�D.\��4��H��I���a�9D�\I@e	�B��z5��n��D`F�7D�<R�n]4䜌���D �Ԍ��+D��R����d2Pܨ���#�b��7 &D�䨆�E_E���~R��ĥ$D�XQ�
Y�V�l���I����O�OC��<^�:PR4k�*�@�
\abLʓ�?��_�l�i��J�6�bF�J6s�����;-Dp �kL<6H@�鰦P3v[��ȓ`�|%�E/\���m-X��9�ȓ~��ɢ��Fa�LA ��"\�Ru��%5�łBJ�V<�F(	H�.5�Ɠ|6L��*��n$BD��z9�X�-O���΄k̥��&,�)��r���d��@��g�P��m�4�PCY��j>D��0j��m��p�Z�~�t��i<D��ئM�q�H��$��`)ҥ��.D�� Eǫb�\�.�!�E��c&D�)3Ï7�tA9��x���P�P����
|�i�E� ��`Ѝ��/�B��ȓlt��ࡗ0Wit$z���>K����?����hY ��>ju���|�x��ȓD�t� �N����(c���P��Մȓ%�x��$Vy�4¤h[�e~ƀ��ON��s��ܿ4���)ѦC���d��9\*E� b͌Z�,�	�G�*3$���;2Hy���Ѻ>�lX8�m�K��<�ȓb��h�F�!M�`��fL;I$^��ȓ�T8��M�NV�����P�x,Ԑ�ȓ���b��8��t#S�l\|(��nވ�G*��.���#!S�i��V�qr
ز�L�@�&�n��ȓw��!��C�":瘈�g�U	��ȓ&6����� Z���t��+���2A̽����%�p���<s��J0,`#  W.:� ���$ȦspD��tY��"<�&����8t4��)Z�L�����35���k*l�&u��8bPia(߂?1�ET�/���ȓ)�]Y��CQ��bǂ�@�f��ȓ-ty���¶ckZeK�(6X�l��B-�A�R�Ń} ��f�浆�b�����V�zAƠ��(��9����P�c!�( �<�p�®E����!����J��~R�*E��O5��ȓ?��bQ�ԌZ�푫l}�	��=D�d�"יTg���O<n㸑�Ԇ<D�Tz�G���1:��M#<�X� D�� �J�U�݊0e^�{�6���@3D����НK����U^4,�;D��zTĐ�?�y��[M]���p�<D����fG,F�i���x���:D����@_ �4�����<���,D�T���̃ ��R2*S�z�����'D�� \5b�gZ,��H�!��W��X&"O��jq��kײx	Ȍ<�Eb"O��aW�؈��\
'���`E!�"O���`�kE�Ih�+��f�ni�"O0��&H���B8�d��H�@T�%"O�Y*gؗA_N�[��#q�(��"O��b� �1��3��;����"Oʽkw���4R�J� �F&�"O�M�f��bӾ���	=$#f�:�"O"�A�38�С��)��0����"O =�W@!~)�acwȌ0Q��
�"O  �e�.|�LqP�G�n}ހ�"OĜ�p�[�&���K�M��ڜe"O�`Q�i���R޶	up"Ol��7�H>4��D��ܦP��qxV*O,h����n�ؓBX�[����'K�0P�� �% 2J�K�^)0�3
�'�!���:��@�$O�L���A�'�\EH����x@ C���{��a�'�=�7ˇ5�V�*7�ԅ!E��'��h�ӧ�1A�����o��ɒ8�
�'��0��K8��pHV��&Җ��'�fi��8pB��u�N���9��'Uz����+&�����c<�����'��l+���g`�(Ί�}�`�
�'�� 1K�洂�'� z�j��''�<�vn� l���e
V�>��9#�',�Q5鏕KA�c�[�3��l{�'�r�YG��N���k�ȇ0��
�'�M�$c��7]�(��7��i;
�'ؚ�P�ٌ
z���Bҿ�0y��'b.U`���@���N&u�K�'�r��a�Q�n!�E�į@$���"O�� ��Hq��d AP�F��""O�@�ZR`��8��Im�� r"O�p���E�f�z���N9vɠqx6"O��؃E�Dj"u�U�����"O���GcX��u��&؀|�����"O��0���!�Ba�䐫+|x�!�"O�����Py����7�E�x�FY�W"OV����x)�!�!{��[�"O���W���-� ��0����@I0"O�,��*ޭ*�)�Yp���"Or�Av�?�8��l�-�j��"O���/F�e����V',���.�!��	��hc��.h �� �ϑ?2�!���FC��"�Nꄝ�A��~!�D��tE�,ƥ�;u��aVMV0,i!�d!ݴ�ㄨ~�$�� ��vq!�$a�l%�foR$a���c#$�>5!�Ę�@�\�� �S�>��DIO��!�$B�pU0���g�rYR�']4B�!��-
�x���k���AL�4�!�$2X7����ÓXʰ]��do�!�DF�tT�"��\R��p䋋!�$Q's3�!�hY�RV"�#��Ppg!�C� _�yjflN��񁓠S�-Z!�$~�"H6K�8I'V�!v���A!���0t�z��-�>'�U�r�Z�9'!��DQ��e�G!2�~$8���!�ė�5;A�#�a����!t�!�d^��R��J�NҀ�U��'�!�7k�
1���N�Y�amG�r�!�	��&�9�L�m+������!�� ����APT�,b"D�ar��S"O\�
w��=+ؼ�@@Ǥ8�Y��"O
T�d*�3L��9Ơ�[o�	�'"OP]�q�Yw�l�UF�u˄b�"O&��3 �<�ly+�D�_��P%"O�)��,� C����PW�Yl*ȑF"Ob���")4G��;��zb�"Ol��r	[^u�À]|�: a�"O�ڠ� �{v���Z�{���"O�p�q���������C�"OL��Z3�RܪԢS�Hֈh�"O"����2����'�b*P�� "O�*Q�.w�DY��f�.I�=�"O�{�䁚0A�2�f4<кm "O��be\�4��kA��:�N��$"O�E�C\Khp��@��z�n�g"OI�'�\"��q�" �p�r��"O�<"����5H���-���H%"OPdud��
$�Qɀ�˵>�j4I�"O �3�HЬO1t�a��1m`NT��"O8`ꡈZ,0G
(e�$S.�(�"O�𑬁J�t!oD�"CP��A"O�qREʴc/0�nV���.!�dг<U�eB���F�b�͌�Ar!��4�L��É&�R�X2J	�4t!�dP������#�l�&�"?n!��Û:�:� Њ��z���ɶG�!�ʶ#������9�Nݪ��W�J�!�d+�J, �dG�?�����9�!�dڍ]������#5�I�|ќC�I"�����ŉg�Z�A�41ΞC�ɽ"H���i�-PFDxD,��yP�C�<T���c!�̀<�D Z��̨u8JB�I;x?�Y�K�;m���g�~} B�I%d�x��_9Y�������,B�ɯ�ua��	y��qXE䋳R��C�	U��M���LI]�1�E�՚5�C䉪wU�x�&�M�	%�� �m�(#M�B�	8�t�5(F��X-]P�B�L��K��	.Ek�y
���9d��B�F4�	F�42|��1�jB��,th���z����^�KDB�I\��T�h {��ȆB�I�lݪ�+�-�(b�.�B�C�>��C�	+-�ʩ�Ն�d��8�PkT|��C�ɚ4!����P������L�<B�#E�Q�%]�NR�q"a�1o�B�	�^�HC3������Y�W�p�
�'"���[b��h�こ�L�RU�
�'�6b�![�?��`c�o�(}`
�'�ؐ�tgY�`R��˂�:gI��'��R$�=,���Ɨ4:����'�H���Δ_����"Õ%g}1
�'.l�3BƆ�.�v���l�P�*P3	�'b%�aR�y��i@>'�1��'y���sD4)aLa��QQ0pZ
�'U��R��6c������)�'����4�_�.F�asA��-@{�y�'�����RA]�0��j�6�P�J�'<����X?m���uHU�𲈘�'s<��_�$�z�c�
(��'6j�X���	��d��|�~��'��I�C$[�j I4�;?��k	�'��mȤK]?D|8�� &������� $�F�&� ����p7���c"Ox���|C�\�#�Z p��e"O���1NO�,L��Џ!���"O6D"�ƿw"�A�t`��-�!�s"O�ڰ��IPB�ޤR�`hw���yB�<����i�}��|��K�y zIr��D�ܼy�A+�䓶�y2��bY�!������F,�y�'�<.R��ˑa�,
�R%*����y����d��P��4�����G܁�y"j,1���6��*2�2����ԅ�yR(@6�^��d΋�3:�ٻ��O2�y�H�sP($jsl�#�2���e�yr��/{ )����!v�8�a&X��y�K��N�LMP�΂��	8dJ��y���0:�u�P�E,	o@�ϙ�y���6��2��(w]`Px�R�yR�&����Իpx	��!�y����1�Jv����1���y���y�v�9P/	��\<2�*�3�y�c��x�0�D�ا'��p������y  n��p�SZ#:�$��	R��y�D�&<��qɇ`
�P�V��)�y2.5�ś�G���h�㛵�y���,&"X���ҹK�-ڤ��yb+M�e�j��emw�ޥT�� �y2��rȤq" D4m��v�R6�yƃ�?��8���7���p$�y@�sV ɷ�"6���qť��y��]�v� �!����3���;�F�2�y����m� O����ˤ���yr��i����)
#*�&�Db_6�y�
J53�̸�b�&4����ȅ�y�Mߖ2�L���Z'O��9��]>�y"fX!¡��Τ��Ȣ��yrK��IZIzw�:��l�bJ��yn�@�I`��{�l	�c��y"kC�	a����\VU�vJR��yb�%AY���3N�조ࠋ��y)$���I�<�������yb�D )Լ���������#�yb�u�ƅ�'pq��E�y®�6�tzt�+��� ���y�$A��Y��I�|t�u��bX#�y�d�2 �R�FP�pN��xv%�1�yb�V�o�h�&�e��� K�y¨J��ġ�N?aI�]pS��yR�;A45�J�.��H��E��yB#�u�xpG��[` {�n�"�y�3a�:AY�C��y&�)�	�y��ߖ5����&a�����SsϚ�Py�
�T�#���J?@Z�ώV�<A�Cӊ_Ȩ���<�l�f S�<Aw*�'��C�B
_�i�T�GZ�<��	+,���xRe�2[�j帆��n�<1�Dk�V���o�+���`&Âi�<����*������'t%�� ���N�<�P�^z 4j�l��>?"ٳ�L�L�<y$��H33�Ě
K��1G�@�<�s�ɻBa�3հ!G���%�Js�<1C` 3>&@Bb�ߑg�ج��Gt�<9dKI2)�B	���P������m�<��ǌ=ҡ���D���ف�h�<aD$���B��Q;y�L9�&Qe�<� L�3��֢R���%Η�
IDE؅"O�m8p�N�<8��l��@��Q�"O��2U"Ѥ	|�ja&�T�~��c"O�򓇙�Im|b��w� "O��V��˄�0t*_2|�*��"O9��m��ZEkħF��"O�8�6�ƷJc$���L�D�N�	�"O���E�^jr��&�L��,+!"O��sՎ�q�܄(c �[�N�0�"OZQ��iT�����l�
�zW"O�-Y��9
�&IU��'Q��8�u"O� �Ů�d�[���2ܼ*�"OR��d+ݐ-R�ݲ�o��e�r%��"O��	e�׆\�Pq�`E�-�j�:D"O����e��d�t�p��Ђd2P=�2"O�ZW�P[�j�H�)S�Z.1H#"O���2혇�XE9Ї������"O ����F.���>T�N�yt"Or 9BOS�7�H �D�gODm��"OB4!�F�ґ��B8`>ʹ�s"O�X1�Ŏ�$� �JD��|�`B"O�1�U����f	�:R�`�G"O$�[pkȕFLFHq� 9��5"O���e-�M�,�zfCH�K�8�"O�]a��D/j���DN�+�dՉp"O.���
c��#�⚣2|nثS"Oh��pG,<���7Bd؆7�&D���G�V
��Z�LX���ŉ&D�h�ǧ�P��rT��G�\5�N#D�pQ¢�J�� � ���i�$"D��)�$�2,��9A��M\Ҵj!D��uj�*��؃�ɑ�jH�V�)D��&��>64�HD�.;ht	f�,D��ą6Kn킓�ěl��H7�)D���L��Ҡ��3-X^���!D�@ e߇��Baf�
I���0( D��Q��A�<�+�j�9�q��+D���.R�}ɲ�Q�
H��|�6"$D����9��׀�8W����*"D��ba��+�M���8D�|b'�-D�ԑGc�H�h�X4�7V�q��-D���sR9v��ԁ�`Q*kV�ԈS`*D��P���	X�5�'P4
z��J0&+D���#!Wy؞H�!�_j���'D�8	Aa� E����HL� �P��&�&D���gBf=�P+�.��%������0D�@�w/�>O�a��D#tb�9���0D����P6�T��g�]*j'�d�G�-D�@���\�*��K�k,X�!�i-D�Tf���|��e�4]�py�%D��n��m놵�P̙�GN�b&A#D��@���:UM���T$�2R�� D� X�c#iB��Yf#O;�
���I>D�\�#fS�/�b��F�8򶀙�'>D��H�@ע;�H�qFE�j��ؒJ?D��@V��]A��[1���r��(8�d>D��(���N4��(����,���׮?D���&b��Ea0,�㥚 +��q`�=D�عdMۛV6�� T�>r���EN=D�@[*ǜg� �I�K�fR*m��.:D��B0�V3��h�$�MO�`�,8D�� �#�6
P8x�j��|���0�6D��h7c��5�F�H���L�F���B4D�|3S,�"|`� �D����$7D�� �l s�3�)����za|�XP"O�� �AJ.#>��cd\C��0�"OZ�&�Љ�IZ1��.s9�=�e"O4�8a'V�v�Z��ŭѠ`%
I�0"O^$�%�Q5n��騶��:F,6M�p"O�Y����.5e�5�������"O�m�f���
��j4bf"O�0��H��d��$��l��T#�"O|�z�B��W<a
�dߔNE2�"O� ��'�#?�0�I��=���{�"Of��"S&㎙ѓGA���[4"O�p���F�lL0�Z$�T�gB��SD*O�1�J�6B��h�\��TmC	�'����o>en���M���M�	�'�՚���P/D�ITc�
�����'��LA㤉 �v]Q����xI�	�'v����H`�c�E49��S	�'r�p�b�A
pyF��� �H�!	�'��@%I��q�E��	ML��'\�	����1��t���3l��'��aP�ڹu�u�4�ъ}%��:�'t�-p�ɔ�<�|�n�M�r���'J�8���iz�$���\9���'��tXF�=�А�6k��5;�<�	�'��D qH� D�pt�f$My^� 	�'D��A��-@�}a�c�.E��,��'�|�(��OHL8TK*�\�B�'���8/Aqzļ!�g�-/j��	�'�l�����-V���4>�`�y	�'�H;��:4�H*�P�:hq�'c.@P���]¨������`�,t�
�'t��*��F>?�!gnQ��j�
�'�F��&
�)ف�@]Y�@h
�'֘񐎓7jԠ�-I�]O�]��'/p��`���krmTaj�A�'�H܁ө 6pA��a�I�2���'tx��S
7Z�Y�pk!� i�'ڤbv#ݨSܨ�B�����lQ�'\xQ륉��/�$1�RDΕ|40���'`���2�O�+x�IKrdO�c7�%��'Gt�J�'mrf q��V��<�']\��#���9�a㐿�\���'�h)k��X2,��0ao�v��A��'�P��D�U���KA j��=a�'�:l�T���Y��03�Փi�Qs�'D�9�r�ݘdB�P�NZ�/��(I�'�,PA ��!^�Z�Q�L#.�l��'=�H�,S Q"n�HRA%-���
�'���¤ �;�H��dȮ(��@�
�'�-���L�h�x���A%$0L��'�D��&��'�%�O/�x{�'�D��ĕ�9s��[�iH��RU�
�'}� (��G��aJ����9
�'_PX���U_:Mr�ɔ��i	�'���N�$�q��	*G� �'ւꕏ�=jA|�b��F�#�X�'�(p�Ë�'�XcP˅�+��I�'�N��C#N�.��;n�'��9c
�'*V-�D �vY�A�Ҫ-Y�5�	�'�F\35�� ڢs� ���%��'h���4,%�(�H33�`��'~6lke��+$��pt��W��Q�
�'f%� K2aG�ir��D��
�'�1�L�E�D�) [�Er	��� $D9R���^����cd��H�K�"Ob����V�b|�P��l�^L+�"Op�q�*t�~�p��[�X�����"O ���d�(< ��@�Ə7��"O*@ b��f
�5k�e�:"�C�"Oм	�E�h�X�d��r���@"Os���"[֡j�?Pь0�U"O\�����$ie�F�W3H�F���"Oޜ���=���Xя�2u��`�"O�hQ�B��m���`�K�v�pu"O4&l��y��T9�8~c���"OF�Я�%���K�lL�]_�"O�]�&K7Y�%���&Qhj��A"O����p肶�J^��5"�"O�XZ5lW:sT�ö���	���r�"O�@ NB����C��4�=z"O���ȇ%S8��j3&�75|�(�"O�!F���#s�	��'�3��V"OKB/l����Ť��A�N|���C	�y"�K#�Z,H���=Z�t;vLS
�y"�E��vȩw��0�,��#�y��4;#���!&è�j!ZBOC��y2'M�|��D�A��pp�NP��y��N'̙��W�4����,F.�y҂גt2�K-t��o,�y�$O.��I��GW u-��ꂨ���y�+Ғ2�p��R�یv�J$XŠD��yRHqQfE�RAP��9�CNH��y2�߉T���CK��J��FS��y��P�u�� ƌS>��QT	�7�y"�+D�@�JV�H�j�@�B̈́�yr �@9�F�O�dX�y�	ͽ�y��QA�4���Y�[�\m�wO��y�d"��K&��/T��12����yb�N.l��ty���9�@�i� ��y��>Z�y�N#Y$=��Z��y�Gpa�J�A	�Q3���0�����'��dEGP�(�s�ٶ%�ȉ�'R�܋��.G�&e�EVlk��K	�'1�d[6h�zb@X�A�*f��<��'������(2us'M�9[lʄ�
�'%�<���4aꈙá��`���	�'X�H�!��1_	&XB�j�_c2�R	�'�z\�-��։ipN&Q2�uI�'i���$�n����<J��<�'@밉P�}�d��sĒ B�v ��'f�Ʌ�K%	k�!S`E5f�Qb�'��E"�A���6���](bEZ4X�'�� �)
5d&��{�LP=h+ ��
�' ���&�[�ΘkQ�20\q��'�*@�ۡ;��uh�C?�����'��(㠜��|�"�δ]a X��'�\�qj�< �"lY�ט��'�z5�A�0��*�W�x��
�'$��!��A�/��d���.�x���'F���qd�$W�,�֏N}kt��
�'�X���e\�1T����'�����'�
lva�Gv�@�@3�:�	�'�,d��*[6���!0x�n1�ʓRH���uØ1���$b9?�Ĉ��H	�u�%�:n딴ZfB۹S�Bx�ȓj6���b,N�|�£oV�T����DVN�x�bH@C���n��H��D�ȓn�Tz��D�m� !��=����S�? @ pBa��IB �ajM���52�"Oj�J��!�R���h�5̢M�"Of�P��q��S��N�@��15"O�$@I c���3���>Ԫ�"Oʙb��O,W�	�*]m���"O���a�"C]�H`wV���qa"O}"v�� 1���sa�E��@��P"O�)s�O�e�:i[�
 !q��"O�w˝$Lo��롄G�un���4"O �Zp�2�`�գ��S1V]���Q@�<��M�2eZ�z���[���U
%]��	O�)�?��b��X����j:�PAc�<!D�L�m���a��LFʌ,a�F�C�<�)^�B^x���WP�\8eC�|�<��bҭ&�n��F"����c�y�<y�+�:�ly��/�\��� &��\�<��@��g���
1?�| �e�Y�<�Eg�>��w�V�Y�`�U�<�����D\����� W�����H�<A- ko�4�G�� m$���	P�<���
v��-�P�K�K)-���f�<�E_(X{D)��8�`8�w��m�<!pN�;�ʗ�#�~�A#`m��X�>�f��>~�(��� 5�����)�D�<i���A�T䛧�H<_\	�'�Z~�'�?u�q ��;\���>](���(D��8#R	n��|��4#�:�>���"�0� Ƅ8P����^#V���ȓs0p���%'�J�#/Ou44D��:�jՈD����d�c/X,��4E{b�'�� ���v����!C?']$+
�'X<@2�j�#�n<At�0 �E��'�F�G٤�p�:��#%z�=R�'�.����G�4�TM[��đr�u�
�'Q��B2G�0lZey���&J���'�
0h��ٓf�����aT\"u�H�,��IC�xT����}q(]e�@L,�C�	9R� b��D�G�1 v�D/CC�I�}<: �aΊ�p4u:��ś0H8c����ɐ(|�4�q�Q11gh���	7�C䉬[��]�aN�6c�Zٙ$G(��C�ɻJD]`w��~8�ڴep�d"Oؙ��F�0��
�J��*iY�<����=��,(x�0�K��7�(t��^�<�Ph_�Q{6؁v �	a� ����V�<�r�\�ju��e"�_����-�x�<��o�N�Ը�b�?u��Y��	t�'�?%���)I��M��o�2H��R��7D�P����=@ 岴	��1���2�A1D�@@�K�TVH�����{B`$D�(XS��`8�������E(�=D����H����qS�L�M��ݰU�-�O,�I,Ph�P����6(%��2�bWv�v#=�'��>IBt�=C���酦�n�`�)�O��'ޞ#!E��-�L�(bPc��J
�'�(���C \�A�
K�0l�*O�"=a��5g5~!q�L>��r��@�0C!�D�-3�����cŊ��1Ԥ7<Lў�P��K�M
"�tQ���W:^�b�"OJ���A�ܨ� Z>:�a
P��z�OY�R�X	p1W�.l�(h�'�6��1�E�$�����kK�a��%�'�@�a@�2��A��gָ�^x��'�@�Z�Bž�8Y���0?����� �I��%[q��*�ʇ�H٨��"O���ːf=����G&8J��"O���1��/�"�+�ɜ�>y6,��"O��c�P�Hy"Ƞ�*��8a:�"O��zҢ��u��5�
�R��!�:O@�=E�dI��WJ*�s�l	�d�0m
@��yb�ԴP-ܝ���NmY�A)���y2kT��D{g�?b����p��5�y��ܧ8���pg�Y���P`Eگ�y�⛈�2�౪؍PR�pp( �yr͐��d;D�.CR渒P`'�yr��1p�T�Ö��2@� m˗FD"�y����Yi<a��%3}C��:�y�'�M�1R�KĐ��L�R�yb$��������x2�wLG�yrnI���J�E��aNQ�&E��y�%�\ҔQQDS�^DI�a�Q��y�7l�U���T�aF���pM���y""��(���3��5H����@4�yrfA W�F�2���X�N܁�@��y��_�	���tFK�ebl�p!!F��y�ELhml0B�nͧF��؛PR�y�B�m.IZ�+��=�D�6(U�y���*�Z���+��4+��%i�4�yR.v�� l�&3@4���F��y�H6X4�i� *��Յ�y5L�b1��0�xk��Ǚ�yRD��~$b"$DC�l|�:��\��y��/	�܍�S,U&]��������y"OǜC�\8������P����yR ���K� �>3H �� �y"���2:6����C�#9��r&^�y�BV� j�E*@�[�6kvF���'5.t*��Y�$�-`F�+\��y��'��͑S���g���'`�L���(�'�H:��(GZ�1;���<�<��'�؈�h�� � 
$�A/EU���'E~�����1��`�*����'e�9Q�Α4z޸�VLO�$ê�'~p���ς
��ӕ�$n��	�'�dkAZ�8`�M)��V.�,�Z�'�L�qa-�t�j�r(S)��<��'���Ѥi_�$��`2�<I���#�'l��{�X
7#�-p���?�l2	�'Nlآbu�h9�Ƙ<���y�'r�}�2�L�æ��,�+,Wn���'{�y@e*�G'���ƥ[0$D���'#JM��,ޘR�,�8�dYs�8C�'�>Uq�0@��F�s�((8Q�m!�'W�ŉ�ڨ�@��Lϓ5z(P	�'�А���:!hF�Y�.��,��'@\ݨ���<t�B'� $�<X�'$�<�5&	�#j� ���s�<Qh�'O����]�x�8���N� �`���'G ��aG߃t�i��V� ˒���'�<�#��A�	}�Z��ي��tq�'H>\�UDN'%�(�v�]5xj����'��بp�J�s��`���\t��p[�'���O^H>,	a�Èw��	�'��#�X+�$)��-�0�X�	�'���ˢ��798`kL�%;�Q(�'���òˋ5E��!Z#�� 2����'h�����5Z�U�+���`��'IvA�cM�9~p �`)ڜ6|L���� �!:��@�7H �4��	h��"OdXB@��N�X`�0��J��݉!"O��J�-$n�¨S�៮h��@�"O�ݘpk�P����E���"O���c@�w���P'�S:f"��"O��8�+JF#���5�/h��z�"O�E���E[t�8B� ۱*��� �"O�0�Y�y��]	dbƧz��D�"Ot���%O�JDH��c,� "O<� ��T�h'Z���f�<U����"O,<x�c�# ��5pƜ�|FPd"O���$ 0�С���'xY��"O�a�eJ0L�`(Qe�ޢB`�V"ODЂ�A�y�F�©���l°"O�q�r	�'�05Cc�F�!��I�W"O��Z����� �h��JN��y"A�'z����U�f��}�����yB�+YbY���ϕe���Y��� �y2j_@�hf��g�Q�î�;�y���}�nK T�S�V���,��yҪ�������F@�P�`�!�y�Sl?������g|������'�yb`J����J����O�\���L� �yb(ˎ@�9�#@�B�b��E���yR(��9?ꈡ'��3;������y�Yd�%� Ђ;a�l��m7�yB˘�A��7KP,7I�T�����y���+9v�����+��0B0��y�&F�tb��	Th�VU(�B�O���y"L���I��o˳L;pࡃ��y�:]�q�CX>y�H�z b��y�kޚ��I7`K�x���h��A��yB��#��p�ړ�-�ge;i���`�M��0?ɵ��w��h���N�5@ihqC�r�<a��	o�t���-=B����j�[�<a�-�	�(Y����6����DKl�<�F��Q�B pT꟠��y�m�<�REW�P�@,�G �!#�N�0G&Md�<1D M.��R�[�o� ���c�<) ��S�U����0`�|�R��Z�<�E� F����\2��U�#�Q�<���){`��G/ݯ-�Z�Hu�<1��)G�8��uj��W��Mbd'�o�<a1C&oh�0�`��nE\�Z�fCe�<�eAB2+m"�����'Z��a�z�<A�n��,AȪ�'B�i;Z�֥U]�< ���/߀��g�E_
#%mLg�<i��	�L�f�A%��m��=��ȚH�<�Vd �1ؐ%Z	L�X"��D�<y�I�J�T!!J\�:�@]�GA�<�՗��\��8R��j��K�<�ը�Nutt�"�8� �q0� ^�<�@J�$�xe+��YoܠYe�c�<��f2s�x� �� �c���1�KZ�<y�eN#n>�C�Hv�\�Q�I]�<�R/Q-D>b���WQ�6|�f'w�<�3��#>���`T+~� ݀a$^s�<!D ۙ(&P�"�\.:��aYD��g�<�K�3Eǐ��dl�Z��Ѐ�j{�<iCP*dM�e	�ɝU"�}BC�j�<�g�Y��\*E��2��"�%T�D���ƲM�fT��`�LZ�YQ�2D�����Q�{Ĉ�Ivx��7�.D�<����eْ�����|�\"�f/D�� �t{���4lxw�(�,� Q"O~2�O�@N8��O3T{�D��"O�aY&cݮς�;���)hQ(�"O
HU`�kî�� -ú,D2H�C"O��BW�@�qR �1���9@�5є"O���B/�6�
�)�yF<��"Op0�5�F3E�R�K�ОB��ɰP"Ov`
S�S���Iʗ'�?ky��"O� rc��"�6,�����f���"O�4+��B�Sy&�"F ��]�����"O�`!�aû*B 9�O;k���2�"O��ńG�*7�{R�N�n�(�B"O�\�F��8!ƍ�A�� (`���"O�$���J`��i$B9J"O eG�<w:d��O��`���"O��R�K���eX��J?��ܒ�"O:Lũ^�M�=�F����"OP�����Xul���ڛ@�x�5"O$511��\�tU�2E�O
 A�"Ob1�!7D�Ȱ"���)#"O��8��X�X<"��D��-�F�W"O�!�3�F]E!���1v��5*2"O�9"!�O)���A`��uҜ��"O8A�-M�k�1���k96�"O�j�1S�x�NG�/p��"O��I��H5���с���)��'��P�G�a�S�O�P̛�O��vo���1dK�`Z~��a"OX�b lA �����cV-2�Ĳ��O���>�ny�	�*�f	�d0%h���㇃&�l�E}�IJT�	=|>d�I(�`YcT	"�~Q�w�N�6`��ЁL "E1!�TD<`!��)"]����dR��� �Ԃ��:�X[҂VA62�4ZR1������Ǜ2AK��G\��́]I!���m�(�"��x����~+�,���ۀQ.��ߴy���? �BO�z����O�@�&94�v��&坴2���"��$�O���EV�_#�� ȏ�F�dp�dF�
dÎ��1'!a��y��FMa� ���vz��'�D�@k� �`�5f��Z�l<��P�E����w`��M�!���z9�QH^4U� !��Y:=�����'�DŐ��\`��C�ɵo����`�-	��S �7H��jk��d`�)��CE�K�u�Af�+K�(�`Y|��<�
�p��K16�@�Ѭ͉ �3�"O�|K�K.r�dm� �҉, �T���50��j�W&�2��2"�%X��4�K�p�jM���S( ��x�A 9?�=�V�M0�^���I�F�ੑ��\	5��m#�B��������>zF��p�](©��J$`��c���uY��	�lj$����:A��!�b�;f7�c���.Y~���Q��)�]��
Z����ˁ��`�QC*�o�(�v	��A�"݋f�֟4����I�D�W��.d�4"�aP�~�d|�0dN{;@�B��A�@��M��E�l�'կe������+��� �n��"E��^Dt	(qDGw�'��@铨��l���,����"����P�v�۟,�|�3���C
`ם�"��Fg�-�T��Z�h��&<s����w`�Eu�l"UEa�����yqO���ɡ�U�T:�ɐ�K�oX�Ѷ(,b�~a�����q���Зf��i�4�z������ɱe����g��*C	4��AD���T�D�QlC�&ds�^���7m�
=�uP$��mΆ��@ҖW�I�Pf΅��(��耩k,a��G Za{�Kp��(�"ѤyXǏL�2���Q�6�t�x�{����FO9\�X�Ѧ��@�A������;`�F�H2���:C��)g��Z��F|2\
C�D�TK� �uC�eO P`���	M��" �sU�<B��ʟ��\w��{�ܔ8�X�y��>q �ݘx0!�F��2�đ���<�W��#l���;��h ��6%� 4
7F�=qeL�C@':VEpf Ԓ��6�L�|��g�+
�
�J��'>F�;[Ԗ�ȅn�5w���խI�D
i�$����:4P�K���<��B��eKB�xe"��$`�`�`�nJ�TB$#��_H<�p�X*J�a;�l�8m�qʒ��b�_�$��S��p�gLU	$��.eͻ|��:Bn�!n^�˦.	�%�l���%N��G��Y�`A�� ONj�n�	^��t��k�.n�h�'�6�� C�b�e�&9���h,H����R&�ȸ��I	Y�L�C䗛R�6er&
�%�μ�ߔ=�61���g�!��U
|m�%�p���DkSD��Ola
�H�)$� Њ2�3� � �%�*X���#�! ��͓�"O���d�D�]���#���35��X��Z?J�B����I9��d9�g?ٗ� G<�z�{��('O�U�<q�]�N�Liq�F�K��	u/���?����AdX���[R�*�p��j"&h�㤝#�� 7�Z�&:a|b@�8(Ҹ!�Q�M��q��+�~���ʇ�	'.b���q�ѧM���Lek��ضC�Y�����H��(O��9�,go����ޑ٘O�j�!⟝j?��q�dI�X,�2	�'9��s�B@>=�Ҩ���n��0z��( ��KM�xӧ���aG�b�F$b���E��q�A	"D� !⊂!����)G�"D��"}2����A�鉉h�� �uh��h&����B�|�C�$����O�<,��AJ0G7�C�I�L:`0�!עd�����2c��C䉔W#����a��@�c�Q�C�ɸF�>)��̴X��\KqA�8]�C�ɞ4�������M��Xx�IP�2��B�I t�<�9#���P9���4%�9u�C�ɦpo�D�V(�&�����I1:�B�I0v9�i�V�?7��4���	�mO�B�	\u�%�%��>Mv����>L�C�	������h10L���ǂc�C�	�p��؈��	�ӃEPۤC�	T,�]�Q&$W��%���Q��C䉱Rm�Qb`�
1���2��+.�C�	�*4c�Y6�����!�>*�B�I��\��݊1��̘'��_޲B�Io+|1�a��b�̬P�c� -ԂB�	%��Ш&OBF{�D:�a�I�PC�	�jP�#V�X��$�ӏXwKtB䉅.����n�#��qP��*�B�I/i�u8!�]Tȸ@�cۮ0V�C�	 v��`s��<"+�]�sFU-w�C�ɴ���S��4�pm�Ӭ	dC�	 ��ʀ�׸G�^�b3.N�OA�C�I9ĆT��#�R����}n�C�	�n�(��Uj5�\Ej��W�g� B䉀<7�zU&W�GO���K�Q["B�	�<!>��#��84�eP�d�4B�I0�dE,�!l�t�i��7��B䉳)S&��D�G ~��0*�>)�B�I?g�:������5Bqx�g_�ٲB�I�#�rhkq/&n��JBn�'m�\C�ɑ�B�a�X8M����ca��"�(C�	i��	82c�K����F�+�C䉜��u�Q�	�b ���䇓��C�	�|OZ[!%�=�$�ۦL��}��C��6��	��.�;*�w�0>N�C�	!VY�����GG>���M7(��B䉊<>6�@��O���m�� �:2�$B�,j�j�R��F�D�hj䌷?\��D�.6j� (�OB�N4� dE�aW!�d�G��颖&ģ��[��]�!�]/DS��ȖLL��Fс`ˡHw!�D�5,7�QVL����@����!�֐y�PH`C�H�`�\�A��k�!�e+�<*�p��L*5��@�!���8`-��/F��쵙�#1!�$Y�m/�h�W�'�n� �Q��!��� CU�d0vQ�)��A7M�j�!򤑻h��5� �;+?V	��@;y�!�Ԏ.�@�ŋD�f�J��
j!�d״l8!��*���"q�Nz!�$��tB�y'@� �Y�~!�� �x�@4it$\Z���C��P��"O�uce�T;iN�9s�eյ ��'"O��82#�	K�~t���P�)�"Ot���ŭ���c���L�
�"O���aB�W�	aw5�]*2"O�u1���I�d��4 �7�ڌZ"O�l�fOG� Y�1��A�
?Ѳ��p"O�d��j�;n�)s)�(q��K�"O@�#�W�Q����^>�b=;`"O���tę'ir�es�:0�>-��"O
��ѫ�&s��8�G�[�´S"O.��̛$c(u�"E+3�`5`�"Oް�%��E��J��P.�7"Oܤ"7@.2�"9 ��/C��7"O�L�wΜ:�ٹ�d@.g0���5"O�D ��S�[g���wC�%A)l�; "O�T�&MX��Q7�J�EL��"O����$�1m�+*$&1�\QG�~�<�bK�+��P�5eU=?�1��t�<1$"U��zs���J`��PC�k�<Q�'�	3zB� "��1'B][��3D�� �O��������J=�G0D���7h�$j����(�O�<5���/D�X��`3./�	��&I�/�)�r@ D����U�me����X�frrx+a�>D�4�g�ڿptdI1Mݩ"n���+?D�t[U�&w88�P�[�R�r��/D���wB�+W=*��H̽7Ur��9D�L��ގt�ŉ�
�&�`���1D�@��K�j�@����?ht���("D��9��F�1�p��&�=�|��n.D��X��`b>dI����b=����(D���&�8IF��g	�t��ru +D�8��"��b�"���-���1�)D�@1e�h�����M�8��F�3D�l�&�U~�b-k����dճ��.D�lC�IE��xT��![bO�)SA�(D�<�!)� =|DH!�d�!O�ƅ�bb=D�D�S��&Hb�9jқ{�B$[��:D�jW͞�H�T��`�R�d���t%2D��𒁒#W16����kT��E�4D��$`��e�#ច3�$�À$D�����m��A�I�m�� �"D��[5�� =/��c��ض[/���I%D� SM�C���PQD�6'�p�r-D��K$I�j[��.1�&�(C��
4C!����d ��e��~j��
�Iܫ)C!�ٻNO�ԩUoځE�X��t)!���9­�V#�(��9�m��7!���>O (��ц]�Bz�C��׏=`!�
,���p���bǄ���I&@r!���w�P�o�q�2�1�@�#_!���6\��+�3I��@���&J!�$�f�X�P�`���S�hJ!�đ2,`J����BM�ZXB�g�!T!��
��H-Q"��bؔ�БE�*4.!�J�`��$��l�3�N�)���Y!򄁽o�&�+�H�H���@��#c�!򄒳4S�$����q�*l�UfR$ j!��fu:E�D*`���f#��E�!���Y�%L�\�D;�b��_�!��1a�F�R� Q���J�O�A�!�A�lr���4`TBw�*�gM`!�DM(�4��ūN	h�3\!�� ����G)?B5�F���+��#"O �cgV��м�p��j��\��"O��@G�@�@A�o]M��r"Oƴ��Ũ]�"Xh���<-'�yav"O�qA�W	F�0:%��	Q&ò"O�� �Ŗ1h��iku/������"Ox�� �_� p����� E���F"O"Q��i1��<��J(c�&d0�"O�E�W��8��/+�8ˆ"Op��S�E��:'�pJq
F"O��`�aA"F�����jZ Y}D��"O��0Ğ}�� b0�FO����"O%��L�6X�ʩx�ㄇ2��,	C"O��:'�?�h��њq���`�"ORq�QF������Sȃ�N�"�w"O��1�mΑP��)P�� >h���"O��s� �`�����E��"O8L���;%�b�Y�%ހ���"O�������$I��E��}�2��"O�, p'
]��R��	1�ڭ�"O��*�,C��$#m�025"Ot�vf�����,�)�$-�`"O�|���+i<��jły�"@G"Oh��#��<�%[B(�1:��}��"O���v)ȓ )lQ �gB4,xz!6"O�@�`@ΑD%�6Ǘ+�x��"OR�[���h�p)�E�90�0�{D"O��$&�o3&@  � =L��"Ov�I���W��E)�OKN��9P"Op�����:2B��"�]�;���u"OlZu�^�P�}��X/*I�"O4pA3���(Ы��d�=�U"O����D��r�n$H��A ���i"O�����Q�`��S��t��"O��c%S�p@�3�	Z�vy��"O�m�-�m��Qg��;	q@"OT�P��7��U�2��k�̐�$"O�v�ۑ]d���gԸ\4��U"O��!�أ!�T0�E��]����"OP�䙈uP��# �� ;=�U�w"O�5Q荙�^��Ղ^9Z;��Ң"O~�4 �,,�L�I��2"Oxiu��=~3|�cΞ0;� �"O��)��^
������ >"e.��"OL piУ��<` �O
"B����"O��+7+�F�<���͒�pNBE��"O����x��,��J�1)��0�"O&�Aa�)�����J̻L�h1"O�M�w��:X`��d��<6|��"O�s҄�:5 �B�.4�䱘�"O"M���#��yc��O�f( "O�$s��@>T�0Z�c4[���Bw"O��Y�`�,-8�`b�-h�^}�"O8��8=��ᢌ�_[rMB%"O�P��`��*'�%� �ǉOM&��"O���&����EۚV:Q��"O��##F�U����aM�;�rq@�"Ot(���sL���<��-��"O�}r�����`���&��%YU"ON�[��cD$#Vb��Da0h��"O���5�ʁ$�)��B��C�����"O���RI�hXN1!A�ҫ	�
3"O E��E�S������g'�,�P"O��(6���7�ʔ���R� `���"O� ���Bس1݆���Օt�,���"Or��E��5��%��Ż�"O������(A�gjI�O�P��"O>�"����cƊ2$4��"O �J�V�wU�H�.� �Ț�"OZ4���R&��f��O�#�"O(�� ��A*B��� p8t�r"ON�ё�0T�,�R�Y�d����"O"Aᢍ��U�V1 wI�n��G"Oz�����H4��!�h��Vi~!�"O�0�@WK���S��(ED7"O~���4rw�-âM��H@j�b"O�@8�	��H��͘�/��Ka"O�i��E� �e�wPD x�"Oрb��/����J&j`SA"O��'��(Y��X �G�T\���V"O.�0�Q7��h�	�15���"O��b�.�L@8�C#>&���"OfԠ�*��IJ,� fE&0b�yg"O<tk3��>4��"#	h԰ې"O�P�$���-�@jf-�}>�s"O�4�+��R����A-^;���"O�41��s���ɀ���_&8P�F"O41��wG�p�c
`����"O,��Ƥ�Ada9ǣ�) 
th�S"O���c�Ae \("!ĺ\��"O�q�ă�4�ԢU���b�,%2�"O4���h`�MK�l�:��A.�yr���i8�o�[��A����y��3rq�S�	��M�`!T�_��y�iT�{�x���i��K4.C��y�,�2w��87TX��r��ȶ�y��qx�cVp�"c
��y�gS/wі�Hi�Kc֙3vG�yB�RD<t(��ډi���⩌7�yB�:5<�<ѷΌ�{r|ݢ/ϱ�y�,�v!�p�AE�ioP���$�y�����߉\���s�+�jfh��`����J��f   �?ɸy�ȓ{�~���l���Z��剓!���ȓ~Z���F�)DԶq{�_	[��ȓ-�Ό��ҴEt5�'@W�Y�ȓk*�8a&B�3�����D�{V4��jz��giַͶ�p�An�A�ȓW?^�:֦T)w�����6B{N\�ȓ2�t�@�Ț6|؂2��j%zL�ȓC�H)��k[/��K)8�)�� W��@�G�z��J�
� mȅ��*���tb
$[���
�.e�a�ȓEH��k4� �\:uO֍H��i�ȓl�d�Rj )zp�2h2[�Q�ȓ�.���l� xN$Uy��� �V0�ȓ?�A fb�	8���b�@_F̇ȓ�J���	lB��3c^�}r	��
�H����Rt���FG5(A�����E����%VR�s�E1���ȓ��q�S�II�ʁ��i�)=����{�hs��P&V`�˃�B�PX�U�ȓ���Tk�:b���Q�A�x��ȓ P���"���F�1۶��`F����IR�|Y�����r㩁�x�bІȓ \�(���Ӡ�~"u(�%l��m�ȓ+IT\J�#Ȧ|�9�aS�<V���ȓ3����j�8&���!bm��cm�P��S�? D�&h�&���� �Y/T�w"O�0���D�@1�4`�#7*i��"O䀲jG���@bo�2��s"OL��Ba�,{:ܡ5Ė�~>�I�s"O�L񦣛�^���9�39>��W"O����3(D,$ Kӧ%z��v"O���Y�VP5�ʬY��Z`"O�]�rn�Iۀ�����$
��f"O���1�ݢ"S���,N(t+d͊�"O�ų ��)��T�����`*x�4"O�CIM��V4��#*Dv9��"O��Ibo�)X�tZ#�·a>���"ODP��LH�h� L#�ɋ�S�Z��"O tإ
�
m����Ǉ2u$;�"O脐��=LԹ�ɢ'���B�"O������,Ȧ��
�*g���K�"O��	'i&mVu�D	���5ӆ"ODXJ�+����;�fЦG�4 �"Ohp����Ӡ��e��o�\��"O�u�3�\�*أ���z]��
&"OqQ �,. u���I�P)
"O���Ԩ�6}>9�sϑM��-�"O��(��Ru~��CD�<�I�"O���R��l?��+#�/9�jܘ!"O�� b� v�,�©��eٌ�@g"OfE��'%���au��� Ƙx:�"O4����p�
&]�q@ ��"O��S4oZ*=�|U�f�-RƌK�"OHd�g�]DN�
B<7\Q�"Ob$!6c��^�@4��Z� `���"O��R4B��Q&��֤	�}�t"O$p`#hE�R����mH��6+ "Of��P�&| �O�62x�Z�"O ��^_���`��<Z�L��"O,�ڥ�W<�2���%U��3"O���s���>��#lZ�i�"O���ӤL	��+P��-V����"O�sP-ԊG	։q����O�<P(�"O0�+�N�lF�(���1v�b-)�"O qr��/?����Eй�b`�"O���20gK����R&mn�I1�/��<F�''
8��D�2H1��@BDY<��3�'X�8�@�U��ē!H%,����'��-� m7Ux�+!	� <D��'p0�*
�c�*Q��=�jI>��ν��<�}��m\>@}�rG���]�~hqr��Gyb�]�v�t)�y��)]�d���B+�:���μf��ɷ>l����.�)�,vZ�"֋ .R��AeN�X2��r�Ũb�
�*��T��)��� ��)p�m�qv#C�lRl��q�Ȕ8���6Q�<���v*���Z�"�0���IE������#<ب�"b+���`YdoX<[�<ʓ�Oc~�������mV2R��m�&�Ǹa�R$���Ͻm�d!+����0|b�I
�k�Me�N�uv��:ZR|��4%5����q��;{H-"����~�K|�uJY�P��Ͳn4}�X�֎˕Z���U,����S��M�;j6�Pt	^�1َ�I��٩t=�$i�F3�	�0|2�K�MlY�׎]{f�J�B�Q��P�X�J|j%N��l3�Da�м��D�P��	2ê��?�~��f�,1�U(���:^�2H��TV�<9��=A7��hS����H�{P�BR�<��,ܭl���3%�}�!�Wn�r�<�.ՓO|���&B[n<HU��n�<�r`��	u�0+ �Z�~�v��C��l�<��Q/b��
3鄷#z��3���e�'~ay�*�Hx<��MՋeB������y�F7&,� ��'����FL5�y
� ����$�T=k�iV�y��Mb�"O��1C��7( ���0(���"O	��"�9:��]��m�6$�	�@"ON�)�'6���(�i�'n��0�v"Öq��^z�l�	H�<@����d"ONm���ߓ{��q,J�|d�Q�"O�� �,�#`FH��̗vY�b�"O���S�ƞDj~��ɍ-s<���"O���c���	������y0�Ub"O�TI��U)1XP��9x�@1"Oȸz�Y(�2��)��5Be"O�]b.mjn0ڳmL�0K�H�"ON�
ce�@z2�C��,T/ܬ2�"O� P�'G�8�4"xJ,{"O2y��s/��Jo��&���'"O �q��N>P��MC�" ����"O�Pk��%���P��e��H7"OL�0�(]��9R����E��"O �҉ZU�����
�%
�}��"O
��AEߤ>����
-M�|"OD@��gӼp�¬��J4z��bF"O,��6 ��t|�أ���Hx9K""OB�@��}�^Q8j4��B"O�Lk2���\�s0g],+`P�{�"OV8�քS� ��P��8PL�(�"O�UYUb��U~Ri��'���Q�"O�)P�Z
7�P�M:l͞�8�"ON%q@�"/��J5�>�A)�"O����hM�C��XX����_Fl
�"O�1C�]�S	b�c��B#��K$"O<܉6�B cr@A CdB%�
m�e"O��؂Kώ�6l�K���|5"O�q����_p�(�2a_����36"O:0�5䉻i;>�ɤ"')���q�"OpK���8�D����GQ��yТ"OȐJU B��I`#��|T�"OtL�� ߏt9Z9I�O�D}A�"OL�ySG�&8���q��|�䲄"O�<X$N��]�t�igʀ�{�L���"O�$Y �ØR#`I ʙ�;~x])�"O�5���-�� !B�%>�I��"O��� >:���Q�m�|�uzF"O"�x3,c�P3ƥT��;f"O([�DU�@NA��g��\����"OP�C���<ʄ���L>@m�Ts!"O�qY"�ߕ#"V��ܼP\��`"O����+ S�TpWʝ9.바��"OhE �+ѦZW��(P|�*h�R"O��eRP�=��7�hI!�"O cC��%#�B���eڼ5�����"O,�(�=G��� ���L�(@H�"O�$�2d�h�4dw�r{̅:�"O�x��O�t]�
��* ��y��_=�89QʔS�ڐ� ��yB�K<F ��ʧ*�2OKZ��rͲ�y�m2Yih#)� I��9b`ݶ�y�J<��0�:qb��a�@��y	��k�0��a��,`���Ja���y2F~�F�p���S��AY`�վ�yr�L��� d��a1��q�ӽ�yˢ&u�����C/`�P$� $E��yR�Tbj�!��T0ڄ��,�$�yҭ�P�Y��c�%QP���s�O��y���=8��;��	�8BY0�}�<� <���׊q������JFp4�c"O�,���ŷs�ވ�����3.�5ap*O���e�9Ea�
��\`�'"�����&M���ˌE�@�C�'� ��!Q<r�� Hg��9.m+
�'�p�����7�^�&�?*ݖ`Y�'��=����-ub�	�#�z�����'m�Y��A�k���E��xO-��'8�$qJ���t�vl�4_bΩY�'�J�0�Ł��aBG�W��m`�'dp��FK��Q���H�>�E�'  4����>��Y��(:,\���'�z)1�cȧ��*UJޡ!/Li��'�E�'�§j���HD�^�J2Ʃ��'�fٹS	��,�æ�xa��{�'I�m�u��6����E�o�p+�'\X�7ɇ�ow�9*���`��AS�'�h�K��4���F�A_�d���'rh��.��x���LC%V}8��'�8� �Kګ��!P��G�M����'�REHq �/4P��gX�L��L
�'rn�`oV�ܳ@��H��
�'���b7�ٹ#U�g L�9�|��	�'6���KBt|}p��2��	�
�'�8m�sKB(���4�69N�z�'����1�E�MRp���3�(9�'��d�V��M���E;�}�	�'�N}��
�l^�Y�GL+ Q�t��'�.y��G61u���	�1u��1�'�`P!�R�l�L� �o��k����'i�h��ɍ,�~3�/ݖa�@��'�ny�E�H5*�@fk�l�����'�B�y���5b�K6�ːz���;	�'K��q�jNx����]G��q��'O>!B�l
�M����"��<��`2�'W|���/����5�ʑ4	�(�
�'h<|q&¥@�� Vk�#�f��'�J4��Ǉ*_��3���*`��'tlQ U��-��Lha�1�N�2�'ld�I `ԫ\��S�iY�_�����'� m#d�݊�b��g�5H�p���'W�|��$Ō`]n���I���'S���ǧ ��cM:q� :�'ʦ�qn�3Tea@��
0��)"�'�n=+uL�;#/��bJ�$ݺ��
�'����qe
Or�0���L���ȓS�<��`D�/t�1t��C�Z��ȓK����&\ ���Q�@e�x��X\I:+��s���AQC�=����K�>���C^~x�ۂ蜝}Kꠇ�[C*Sh�� ��X� �K��x�ȓ9O�IRp�2qV�%{�A� 40��L(Jxg��j~lx;eNb;�y��y�0�t�%�P�kE�F�|���ȓm;D���>8�r5�1�O15Be�ȓ��<��bD�o�^�SP�4~.�Y��eH����X �Qs3�-� ��M�r�-�I���� �*�z��$���a�郯9����XBT�A��5�n�EE�'*XD�@'�3������f0I��2/"Y��/Gmp���'G�<Hb�͘^^3#��1I$ʕ�����2�X��X��$��1E��I�ȓS�ư+2a�� ��oC���S�? u�A�ħ+� KO�_j�Z"O�IYB�ߢl<��Dt��tY�"O8�	3�¹h��z�.�.9��]b3"Oz �6A�H]�b�,�ɒ�"O�ظ�n��,ش��Eg��V^�"O����`�3�p�2�(�Vيc"O2H�S`�a��f�LP��e"O�	���e
�� �+�%b��d(!�$��&�Dd���~�:��T�U�R%!�.Ex���֎�'�,���2!�
.u (�#�>R��`P��I2ko!�ބW��\�AѠ��}0��֎!��D�~	,4�������r����P�!�ߓ�n����$u�3��ي?�!�w��Mp����>�* ��� (�!�D�	\w��@f'�=�X�� �!���,�t�B�'�ܽv
�h�!��E:�ج[V�g�M�T�R4�!��T!8��m�r��m��U�7�E�g�!�׉�DI�]�}��(6��Q�!�$�Ixy���t�Z�j�1F�!�%\�f�a�Q�y׊z��L5t�!�DU�0�t�QT��7<]����A$�!�D�H����Лf2̲Sל"�!�d��^�4�6EIv0�7ki*!�$1I"�A�F8F�Ī"-��8!�d��&tv��WgM/E��Ȧ�Py�ءa?�)�M��'&y*d�ڮ�yrf�
���DF�l8�֒�y�B[9viM����H�r��:�y���r�ة8B��6QE�k�E�y������Іޡ2� ��� �yR(�)o�UH���h��@���y�i�-@�(
�*	�j���3C�y�����҃��2��pi ��,�y��K6y�(!t1>�'	���y"V�8|	�S�� �@�뀍�y�<8;�q�Dqm;&��d�!�ߜR�~ٲ���%M�*�'@'�!��5G3^E�G�%�n  �hB�	�!�$֘�ȡ��d��B��mI�Y�!�dJ�!.4��+�?��(;u��SX!���Q��
0��+�����;F!�D�yw�E��̊�yl��H��!�P3slZ��«V -s�e�JJ;S�!�$�:��CS�N�ȤٳC��>�!��:wݎ�*����_HU���sx!򄄯{�����^'BR��%��Qj!�<L�
�+�n)G�(�k��p�!�d�*0GB�{��O�cj�P���6QO!�\�=�6d�C�r�"Q��aV8R�!���X�. �e���X�r�A�&�5!�$�O;^�s�m 5S���9���!�D��2HB��A�_M��; n32!��˰EK�T��ϫ.� �I�ķ	!򄊵I�D�C,�	��b!����!�DL�6���W#��*`��F�U�!�^&V��*�
��]�U` �.L�!�ҏf�fDcK�lYfx�n F!�DA#��%�V@��x��V!��X)
�jIJ'g��?0d�F+��!�䎙�]�CkW�	&h������!�J�+��h��_v��*��E�XV!�DB� ���^)2
_(��"O� �Q�N�r�% C>��`@�"O�t�Ώ{'R]�ph�FHXe��"O�t�$���u���Y���}�"O���A��	g~a�Qχ�"��@
�"O�}`��g�mIԤ�.b�e9�"O�qC#�5�]�2ꆾ�M��8D�|2�
   ��   J    �  Q  �*  �6  'B  yM  W  &a  *j  �t  
�  ߉  <�  ��  ��  A�  ��  ů  �  `�  ��  ��  '�  n�  ��  �  H�  ��  h�  C�  � c � 0 �# !, �3 �9 1@ �E  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h%���븧�O@��1�AE�8�QP��Z�	$��
�'q��&װ-��J�gI�H�'|�仳n޽�j�R���*[�����Z6����C�k\���T�[H~�B��D]HV��
	����2�W;���'�^���d,�'HW�ePU�K�D��!&I�� <��6���$�8x
�Q{�/gY���=��^�б3�)�+("�F/W�4}����ys���Lס8����R�%:������?��.ߥR������'/�F����j�l�L<�@��=l�{�nM%VZ�����i?���S�^
p�Ė='�:���l� C�I�HX���4������ݽ}z�C�I5n(]r�'oϋ%P:ӣ���?��Ob�"~���/Xr(+��ˀ*tv�	s�E��y��]Te(���aE1#ǒH��f)A���F��4�$�͌]a2u�0��@���q��"|OHc������Ţ�\�?� ��>�	�v��yh�5��dY�eݽf&:P*�Aޚ�Px���3:� \I
�<I�y6C.9�֑���>�4�*lO�0�±�
������ڨ����c~�>q-OT�	�F��pa��G�z�qf"O|	�t@1����v�K%H�J���"O�كh��<������47u�HY��',h�O�i���B$;��hu�Qzj�(�p"OheБ������ �_rW�	��HO��/od���
b~t�`��~�B������*� 5�d�h�!�(ǶB�3L���a5���Q��?�RC�IM�R��&l�����G�g�I���?	r䐃]Lx q"̖�G�flpc�C�<���+��XuF�/�}����}�<��){ji��eH�T�H��R��zX������ ���J��ZVvE�$���m���Q"Oظ�AQ�W�4!Z��۶7^*8��x��)��!WI�8�Ȏ< �����)J;JW�C�I9~@ h�)N�̖��臰T$����q��G�y��N H)�ݨ��ב5�b���+\܍8�X�`�J��0l`2�D|2�S/����gN^+z1jE��>�C�	'Gp)��@������;W7nB��+O��Qp�L�*�m�)�~�BB�Iz7�l�E��BMx�{����<6m�����'��\�Aބx�8����ؕ2��H����$�<!aA`}j@�'"m� 2�U�<�4�C>y� �R��ČF�ȅ�ULT�u���O�����@�V�:a���?�X�
�'�` �,�.��ujw��0s�Ԛ�'�V���*�^��s��Ŧ,N-+	�'g.%�$S6*i���Ԥ��]<h�'-�$��WC���R*7Όq��O©B�ɖ�U3�C)G"t!��"O���Tc��t�:���Pέ�s�"Ox�r��f���&���\��8k���u���'C�ؔA��V���RBoشo=�Dn�R������OS9� A ��C.����1�8�<	���O޵C�
n沉ar-8�Ȅ)@"O�iS��#df���Fꂑ$��{��'��	-26pQ5%Jl&��%��ZD�<lO��<��h'��J��[8<�����9D�<���J>{y�R��5�μ�p6D��c∝e�tLڇFK�F��@�.D��S��xj���`"	�{�̹7G9D�d��G�6]��uL�. Xr����5D��s�c�d
D r��z�(P��.D��ؗi�7$��m�� ��0��|3S'2D�TyϘ47���8��B�&����*��j���'U��(!l0&]X4�2c����5�}�%��$W�ژ#��7K����)����`h�3�6M3��<aj����8D�C' ��f�t���C�sQj��/�ON�[
�1�5��
Հ��to-QML=��>De��)4@��"%ȫ|Zͅ�b�:��r�HvD0k��1� �=����D�8&$���i�e꬐���>�y�
�=����`��I����W�R�y��І���Z#FB+X������6�y�n�	h����P�:T�r�/y�����A8�x$Kk �1��P#Ԇ4�����$@-Jy!�#�G&�z����<$�0�T�sYx��C�Y���'�ў�|����#v�ᙑ'j�C�k؞��y��Ω�,�BT2t�my���y��Pb! ���#�<U�!P���'�ў�O�x`��Ku�˦�ϟ�ex�'Q�i�@�M�E6��Q�A�	�4�'V��QDJ;���94L�#9Oʰ��ј']j�3BNߨj�x�G�#��`�'���jP+�-gN��jP�X����cӮ�}bn̊#2�m�ǅT ����Zr�<�a/O(1�ޡR�'�Xy��	V
ָ��D{TO?��ݙ3y��$MN�!�d�C[?S�!�$G�y��qFb��0P��0�F�*����>��M�6
�P�ꒁ�.j���W�Nr�<1����03��ǡVQ.  ��q�<��B�Heb}2����2����To�<Y��+Q����`6XF��F@�n�'��y
� ��!ыe�he�1GC+9m�t�`O��j��0Q���F C�
Q���ج��T8����I�'9�p��e� ����+4�Ot�"�'��l�`�[����s��s�|j��HO$��-�3N\��2���P%"OޘR�CKe�lm��FW����c5O|�=E�t���\#6����/�n�`�N���y�M�fs���7j�:zl�������џȅF�:�(��4gE6��3ED�	���$�<ѧ��1$FH�xd$VNΠ5��a�p�<��A�O�H�2	 �(=��2�kQ�<�1ˁ�r��y�vʽYR6!p5a�M�<����C�\��J�9 L�8sd@��D{��ɗR%�I�e�=V\��O]� r�C䉲#J�Q��G�x�Ԋ��.B����	�7;����~��hOj���L�?}�4���`��K*���'�2 ߳
4b�얏�lՋ!�Y26HoP������� )|!@E�Z��v���
 �0=u�?�(N�Q�Q.�o��ݪ��E�V�,��p?q�F!���{G۸��ؖ�]cX�,�O���E�M�a@j�a�	#\���R"O� ӿ�Z�00��H0ֵԐ|��'��O^b�(#�l܁2P�*s�R�\��ǩ4D�4Y��y���h�Ι&a��0D�|Sf�94�,%��`��w,.D���K�o;�0����> ��b �'�I\kQ��Os`����4$��M_'>&N�P	�'Wf�# S	���8����*�NE�v�:��h��_�#�����n_�AF��0SE;*!����7� =� D�"	�H1R���A�'�a�iZ�UBج��S�Q�� 8���y"��zh��Fo�J�d��@�y���Ql�X�P�4��͂��Y��y�ܩ"Pɩ"�J�5Cd�#��+�y�
�����2��=Wk����:�y�@o��:pH�H���$ �<�yl�aEX�9�o�2H�\\rtB��yrGOWG$�(CfR�sܐ�6�ϋ�y�gJ7.����F�q�Q ��ߘ�yƔ�P��<�1�A=�`MYe)F��yBV0D��t��(�:/�e�"P>�yr�C�[
|�p���#$�4Qd\��y"bϵ>,�]�aW����#0���y��K%Y_l���,O� GNL�B�M��y�8c5:5��	�#�!(g�R��y�^�6�Y &�ӱw*1&		6�y�j��o=�����i���y�F
H7^D���*E�PѱaO�yr��*8�(S`���^8*qL��y�CE�UI����Р�p$�y��D��Cr��4n/�`�Q��y�I�1A~�"��s�p-3`�6�yB**t�yIB8o�q�'nâ�y�9�fȢr@�oa @ʖ�yB��8^Jd�1L�,�rk��ybF�l�8�)+ ��Aqf���yr�?p���1��p1�J��yRĈ%�!�i��"�.
DM)�y⣋��e2 ��	&R��b�A5�y��I5hb@l��ٗ#*�[��R��y�FD"?���-�<���H��y©�Li���-����/��y����e�E�S�U�)Kp�QBY��ybG��N<�PN�n�t���(X��y
� L�����S��z�ŠdrR���"OJ��4���C��5�i�j�5�$"OD��P%�pD�P�b-�蘥 /D�pQA�OY���JN�77�����@?D����Cͯev���R~ְ���O���O��D�O����O��$�O(�$�O��(d�Q��5���� � i�O��O����OP��O����Ox���O��Ѱ�΂�R�@m��,D�RM�O����O����O.�D�O^�D�O����O��@�؛���"7�������O����O����O����O��$�OT�d�O���W�M�Q�ҝ���1X8�tᑻ�M#��?y���?y���?A��?���?����^���P�(��|�"�����?9��?����?���?����?���?�VȄ�|Qth��
�w���ڂ��?���?����?���?����?q��?�5&R'q5�|36lL�)���;�?����?���?!���?a���?	��?qD�>03J}�hL�B�xтB@��?i��?A��?����?	���?����?�DO���[P�\��*e)o΄�?���?����?	��?����?)���?I���JQ�HТM�q�t1����?Q��?����?I���?����?Q��?!�{Iʅ�/���ӱ�P	$x�	˟��	����I����	꟤��۟P���n_\Tq�J�);8��;�G� -p\���ʟl�I���럼�	Ɵ1ݴ�?A�tm�(0�/Z�Z�,�XQ�Q�&� @��V���	Iy���O�mZ
/����ށ�Ր���?9�E���<?Is�i�O�9O��DQ'6�΄C1M_ {0�����n֔�D�O��!Q!g�����$!��4�O���`���'N�8� �J��S�5@�y��'R��O�OZ���_%_�e�Dۢ��x@��i�����d+�� �MϻC��@���_8(��eMR�P��D:��?Q�'��)�S4:d�nZ�<adk�5 ���&��Dr�L
b�E�<a�'�����$�hO��O�1PL�`^�1!�Q(`2v7Of��� �v�M���'�����h䴄���X�܌a2��l}��'��>Ob�V�RMeˏ�~�����K֎>b���'�b���^�H���d����L���'[ܸy�,�
��A��ǡ+��Y�U�X�'���9O��ZC��`�]�F�D�r(�Rv1O$�ozK�j�Bӛ6�4���2`�	e�8
 Եs`&@�E?O6�D�Oj��	�E�P7�(?ɝ�៸H�� �e��L�t��Sk��(��P9������d�$�D�;bk�t&�jS䅭?����M��!�����O��?A����P�V�ç�!�!�����$�ئ��4%����Ox��s�N�J�j������M�6K�T����VZ�����Z�Z�'{�Iky�O%5��p,� �ۄ��-/rх�*�M��_��?i2��J�,�ȥ+T=dy>�Z'���<	��i��O:i�'x2�iN6��N��$8���9��e�Ă�����){�Z�h��%*6�?�'?e��	p�҅����5�T�hQʖ�!���	x����PC�0�Ҭ��4�.Ո#��NyR�'�6�]�p��4�M�H>)�$1Dʴ��N
|%���?���?��|��S��Mc�O���cNf�X�-ˏI7$�Ҏ�3vRfk�$��h'� �'��Oΰp��1lk`)3�E�0|ɖ Xe��M�Š�&��d�O�ʧ:��5Z����#�J�s��U.wЂ��'*��?����S��aͮ[��\�A��Z{* ���I/�T����$Q�o�<ͧ_���^�8P��,��T�G��Rϒ�~����؟��	Ɵ,�)�SLy2r�D���C(~\��������ae�%rY�I��M���* ��̟���&SU���"Fp!�*##x���ݟ��u�����̓�?i��ܙJ����y�]�����g-�24Q�� �'@��y[�@�	ٟ��I���	ҟ@�O�B�0��@��x�+� 8h��Q*r�F�`h�Or�d�O:��v��L���	�l�J3 !=�9C��G�9�^�Iԟ0�K<ͧ�?�'>��Qٴ�y2LلIfd@�K
	���yRFV$/|���� o�'*�)�0�"w�;���B��tK�_E��9ڴy��,O(�d�
��`A� ȁF&U��8Y���O>�$�O �O`2�לLNLQש�)Z&��2���B�Ӌ#��mڕ��F����(* 3�>�c��O2F9�2�.]Ɵ��	�l�	��E�T�'~ء���>w�h�S*�s���v�'�6͚�p����MÈ�wcȉ�SI�$x�A����?jT�i�'��'fb��Uԛ6���1��Z�Uc�i�}޶��*�2x�(�b���m#��O �S�g�<��8{C N�Hst#SF����'	�6�C5l@��?�����*H�\)�@Z�Z�(�IA�F�!�P�
ћ֨b���$�b>	���Ѥ&b���ND�k���*d	pv�lZ����U�I~���'$�'=�	�?��C���V0�#f#�C�x�	������$�i>Q�'��7�@�CN��\<�X1�hSZn�P����^�����Ȧy�?A`U���Iٟ���4�V���kL8P�̚�ّU"�R�!ב�M+�OP� ���0�2������ X<�D��t�͹�J�P8��;O����@pz�P`�3F�:���b m�x��?9�i�N�͟f�nK�	�r||��@� ;�|@q��9��!O<���i��6=�*i)��f�~�6��e$^�Z�"M�c
\�1j<_E���������O����OJ����6��I��\�K3N�`S'W�)2��O��Da��jP���	���OM��"B� ?���H�) iz�O���'���i*0�O�D�O{p�c�fӖa�1['o��:`0��,&���Bu�Y�����|m��f��O"�X�G)�"(�%�T3#.�ebj�O(�d�O"��O1�~���a�5�b�U��r���l���$*��'�RboӀ��q(O6MX�"��(
�i
,4���� [((�m��Mk����M{�'��\t:"��r-�'1x�F'�7cFX8��%�T��'q��n��p �f*[�D�H����MK�M�ciވ���O4�?u*����� �uwЩ��Θ1"�P�3���?Q����S�'Zt�Q�4�y2��M�D��I�3]��`�5�yR��I�5��������O���4�V����C
7�x��n\	(���O��D�Oj�R��-D��y�'���P�Vu����M	(A'���O�H�'��'�'����i,_�.1�G�D/^x�<Q�O]R���Z��7�%�S�&����O��ѤvB Cv��
���b�O��D�O���O8�}j��+%zu� �%0����Ģ�L�nh��'9�n܁5���'�6�)�i����"�z���	[(m�2�����Φ��ش��ش��䍄�y���
��5{E)ПrުiTaJ�&aX:[�?!,O���|���?A��?���"^�<��Лu�|�)��'¾ѣ(O��oZ�-!�4�	ğ@�	z�ğ���	^d�P�jn��XF,�pr���?��fۉ��OGBI�W��5G3&�4�F�2̒�y%��?�JHS�O�%s����?��L&�Ġ<��JQ	>���j/:z��P�\��?���?i���?�'��Ҧ5���ϟ�0S�̧��p��-ב�ʨ���o� �۴��'�
��?Q�d���W�#z\I��l�/#o�����#5�"u�Ҿi:�	�#����E�O�q���.�'&юI�嬅�5�Bt����3w���O`�$�O4�$�O��� ��f�����gǇd".�6�;C�@�'�}�8��s�?��4��1m�1��M2s�&ur0]*(�h�1K>q��?��)��H۴�y�'`��b�Ǔ(�x�XTH�|��!��'i>M�ɊE��'k�i>1�	@��:=DE[�Ή#4����"��+C�������H�'�l7M �����O���|�V��OXm�w(�Mb0�I�`�M~�J�>I���?�4�xʟ�	�]�^�H9�&�V�fC~qҵ���x@�虖��n6�i>��c�'�l�&�ppC�TNf�(���
���"�
I��H��̟d���b>є'-�6M
oh� D�n�(��V�n&��P��<�i��Ox��'>�&�('��h��}�x\p���.��6��٦�����Ц)�'��(��DB�?I��Z�#�d�,/]K�(�>[��k�HH�$%0���#Ҳj�ʽ�!O�@�����&J�*�0G0�6��Zađ5�4&��Y�.��j�����Zo�V���k���j	���ɀ'�@;9Ɋ}�-Z�q��l���O(���d���C���hW&hIB�%�xx���> t+���bb D�S�m�ԥ{�BL^�x��@� 
�@�  ��/&����iEaܼ�����_$/�daPE��`���%:���RRjBI�A!�1.��̪E���
v�����Y�"� 0qS	I�M����?a��
U[���'�����/�8|dv�؀�
�V.ؠ�h�D�G�,�	�'�?!M�/v�,��� ��j�:r�M�r7���'�Z�M�S�蒮Oh��?q�'fNX)Rʹz<��('��
�N�ٴ��4Dh�a��T�'~��'W��K႘�W��=Ic�	�,y�,e�^��V�2h��'���͟h'��X�;1N����
�,ѓ�˞�l�-\e`H>	��?����$Q�pdx�d��b
̈�dJ��-��LZV&YG}2V����z����I�~d���I��5�<HQ���$M4�vO8�	Ɵ���ٟ�'���qP�z>����  @��q�"!�9�rȲCKc��ʓ�?�N>���?9��L��~B� ��䑢�M�Y<-�Wa_�����O��$�O0�&V�	P?q�I���(7�^# ��kpL�J�\�ܴ�?qM>���?9D E��'�f�`��+g3f�3���<�Xa�4�?�����B�X2�Y�O���'(�ġB1`)��W㎙i�$p�
L.-��OP��ON}�Vj%�I{��.��S��mP�ѶUFD��צ�'���Nj����O����NDէ5F�A�H�	��=|wF���xyo����,����?���D�\'*U2�`v'\�d�(l��+��M�`��Fϛ��'��'-�T��>�(OXQ97Ȕ� N�����1W������EΦ����v����O�H�p�q� F�%f8���%.U�7��O����O����Sq}2V����o?yC�d�����-�] `Y�D��a$�d:`!���ħ�?1���?Ʉ��l�!�3kT.8<�C�L����'O���>�,O��d(���ڥ�JY/���ಬ
f8��s�W�Hy3��W�	㟠��ß4�'0���h1�o�袕+��H�x�`T�l�'�B�|B�'�r`�Y�$��kJ�2m��f�(5��@ e�|"�'���'��	X����� �Hx��/K�@� #��02:�x7U�h��ן���{y��'_�"�/�""L%��8
e]�Yl,����;D��?9��?!(O.� �PE��1�����F�9��`s I�[�`���4�?Y����d�Ob�D8V���,��,ׯWb�q�ժ~���z%톊�M���?Q-O�x���
k��s�����X���!�m(3�ӌ(��7-�<Q��?�k�&�?�(������k��eʚ(9��Z�tnH�〈�s���\�l*'\��MC�Z?���?A�O�)HVo'M���2DF24�<�#�i���'|�t�'N��)�|n��h��=�G�V"H� J��^)P\6M��j�����OD��O$�I�<�O�������p�)��E��!{�iӖ!C�π�ZE1O>����̭uL��H
b�z���B�T�ݴ�?���?����*i����T�'��-ԏ�L"AoW�\W�����bl$7��O����O�qFJ�d�T_>���^?9�K��pJvG���֍��+�ݦ!�ɼk��̔'��'��'Y)sb�X�1�@T����
.��Χ>�k�9y.��'��'O�P��q�V�"�h�RŒ6d�h��	EbE3J<����?������O(�ʜP� �qІŤ����B� �C��1p��Oʓ�?���$�O���v�?ݓ�K�Y�\T����,���n�L���O��I⟔�!�] E7���|�n��7!_�*C�X8 ��;�	��d��џ �'�p���(�I�8ϒ|�ӯ���Ƽ��O�oq`�l���Xy�'	�"�UO�~"�F0B��Y�f�fF���¦]�	�d�'�FE��M8���O�������q���)�M��MCm֔r��i6�ܟl��;`E�m�	^��?ט,��=I!�'D��-�����6��<���Cg���~����2����R��
�tŰ����(���£}�����OF��O.�'>�	i��4��jAL��]L(`ZҁE5c�lo�x�Q�۴�?i���?a�'>r���\cn�� �VP�6����:iΎ�3�4>��B���?Q��?��'����5�=۠`[�3����p�H9�M���?��)��i0�x�O��'�<�6�57�� 5�֌Q(l�a�}�����O$�Ĝ�a@t������O��Dȍ,�p!�P%�;]"�����v~�4l��5�K���|���?�+Or!9����<dtD�fU�.��t�u�R���	�T���IWyr�'�B�'\�I�|2Z��c�N;��l0���4a�,m
w�Ń���?����?*O��d�O�yv�H��[g�Ϥ>#&�bEOZ8�$���<���?1.O��D]>{���Sr��M��m�$m�y9�
N�7��O��7�I���I�^+Ě�lcӆ���.��qachL6g<]S�X�t�	ԟl��jy�B��.�
�d|x��K��q���`\���Ŧa�I}�	wy�AF�2QR�~�DjƵ���ɣ��j;�17����u�	ByB�'Tj%+%S>}������s�ie�\�9�6�DG�L4Iz �'��O��$��2a0��T?�Pf�^:�p�*
y0���d��ʓn�T@��i�J꧃?i�' ��	m��ѹ٧C&,Բ�[�9466�<qGM�?����TR>���z�j����Cd ��r��.i�Rmnڙ0�ܭX�4�?���?y��i�Imy� W:���ɍ|[�M�!J7�EY��D�O0���O�?��ɆNp�(PV��X,29еΖ*.�Z��4�?����?�0����Ty��'/���R��x�a6�`4sF�_b���'�"�'�r`���)�O����OhHI 
�O]D|RDҲ!s�d�J�ʦE��$Hd��A�Odʓ�?�+Of���XhY�����m�0b� e�R�b�V���1�y� ��ӟD��ڟ�Iry2Ȏ�Ib�\�)�;IԳ����������>*OZ�$�<��?a�f̆�R�
�NV��& �������<����?!���?����3<>M�'p7r�������#��'1)��mZLy��'��	̟���Ο��`�l���5�0��01�F6t@����hֿ�M���?����?�/O���D#�z�T�'3��p�c�v�j�(�;UU���j}Ӵ���<���?���a��h�O��Ą�1��dYDˊ�X*M�3�v���'�[�`ޢ��	�O�������;%��U�4��W���2��}
a�[x}��'��'h�ʟ����$땕YF,����!�i�g����M�*O��������	ן��I�?��O�]�9ǲ="7�͞v�P�1�^+k�&�'�bM��y"e�~���O��a+�-�x��R�b�]�@�۴���!%�i�r�'d�O\�듿�\!:%�Y�#g�8+ u�S��C���m��:&�����'�����j3ph{�)�D��� 8�p�iM��'�Rg�����O��IW��" �jX�ԓq��r*꓁�@�Ba�i>��	ԟ���p;�P�W�,D�hd��'Y����Jl�*���`5�Q�'��I؟ȗ'�ZcNx���*�vM�EIZN����O��38O����O��D�O4��<q/�(.ܠ�v(Q0MvF����RE!<\A�R�H�'��[�L�I՟��IO4�8��!G-"��P���6�(�c��k���Iʟ������ly��Ǧ
^��V�ht�sj[ 4�T)x��H�a��7ͺ<)������OL���O�E39O�����]ZD�s�̀"�<T*�L���=�	柄����̖'�@d��~�����3nz�a㫉�F|��ـ�B��U�	Gy�'B�'�\��'b�2JT9��	��H��T�Vؑo�џL�	UyR`ݐ%��'�?)����P� ZL���)p)�QR�%�Y^�p5^��������0i��g~�ڟ�)����K� ۄ��]����!�iub�'rN�J#aw�D���O<�D����i�O��g�R�q^]�gK'� A�jX}��'��(@�'�R�'-�Q�i�pvV�4�ڦ9�i����wp�� #8(�7��O"���Op�	�p}�Y�d�#m�$I��CD�1Ҳ8dmN��M3  I�<����"����H��Ͽ[��a�l�	'2���Â�M����?��<!te��P��'�On��u�>q�V�Ai�+�ru8�i�^��P �b��?����?�u��)W ���q7�$����!��'�J���>Y*OL�$�<Q�����.�=�VE��x5�*�s}Bj��y�[���I���'?���g�F,��4���	#��?J��a�Oh��?+Oj��O>��WmT����
$��1!u�M��u��0O����O����O��Ī<�T�W3󩝶
n��t�Co����Q¿Dg��Q����Iy��'���'��,��'V�	��	��1G	4�s2e��M+���?����?�+O,��t�Ec���'$`��'���9����lݺ7����Q�u�&��<���?��e�̓�������ː�qi�ɋ�4���oZʟ��Ixy�k�y���?I��Rs`�(���b�f��Aj�+��K��I��4�	˟p�x���yBٟ\�`Ů_�����s��C�Դ��i��$\p��P�4�?)��?�'b��i�)�V�aƬ�BW#ѣ6�&�p�{�H���Ol��D����'6q��i�#(��3dxTk�G\�=l�Q�i&�8���l�2��O����H��'{��A` ��$�2=8���'_o|�)ش(����?�,O��?]�I�O�t��B �@St	��+^��4c�4�?����?�0���O�	|y��'&�d�[�bM�e��6Q�0���ZF��'��	PU��)���?���[��0� RW���%�D�^�v��ӳiBK<WG�����O�ʓ�?��S�B[�̃�$Z����Ɔ! ��'A^@I�'5��'���'�BS��I6jG
B���	@�]��h�?M�tD;�O���?.O����O>�$ӱgh�B�B3NP��
/�Rt��6O����O��D�O��$�<�q"��`����2z_|���� �oK^��c��ڛ�_���IZy��'���'lΨI�'��(�l����u���^����uӔ���O|��Opʓv
���Y?��i��k��8��ya �+J|'tӠ���<Q���?��iy�����dߴO0�=[U�	 ��U�%�>��f�'�T�T��Mڝ��)�Ot�������8i��hEL�Gp����,\y}��'3�'N.�ӝ'�'���A�i����7�6��� R�0�&]��Ѳ�%�M�"^?��I�?�)�OD���n�^5T�(&�V��n�B�i����lR�<aL>!���-:�X���0����Ҫ�M�
Ee���'���'��$# �D�O`�qڡ��R�k�����f��z�aI���'�"|���J���*c�?��Z�`�� �p��iG��'����&O���O&���@V��S�E�:��ԫ姅<	{T7�*�D��3j��&>���ʟ���c�J)��g�&������<I7��3�4�?ё�Ra;�'���'�ɧ5ƍ�_E�AIЈ\���T��cI����[X�'r�'{BU�|X�F���-��<�ٵ#��%ndQH<���?AJ>	��?)�L�n��%�!e�;h���� >9V��������O��D�O`�(Z�ᡤ3��˅`ܤNR��b�$E�%�TpБx��'Z�'���'κЫ��'�t����T�k]�����>y���?����$Ԧ��%>Ma%��� �4�Q9ॊ�7Oś&�'��'�2�''p�y�'w�Urx��h�5��Rt�l��nٟ0��xyr��9���p���X�Cы�j&r��.��)�"�"-�d�	�@�ɶ����O�	@R��#c�L��,J�gJ�HU'঱�'��P�(b�F �ODr�Oq$�0��\1D�C�/|��1��SU�̱m�ןt���i5��Ix��T�'���� �	
¹�3�C�b���nzq��Pɦ)��ǟh���?�1�}�\�z�NaX$,6���CD�P�2"47m�i����9��;�Sɟ�;��D%()X�+��]�D���.��M#���?��[J�Y����O4��p��i�"��Z��씷M�6�?�dӸ! �?��I럀�	�c��#��P�RN�j��C.o�HB�4�?)�I�)&n�'�B�']ɧ5V�M�yPx�cm/�J�7/F������Rm�<q��?q����$������ǈT~���-F7[����cJ�p��?�H>����?���%	މ˷οPd�\Y�m� bڱ�������O����O�˓a:�`�0�p�y���%H�AY�eݒX!���Z�,��Z�'k�*_�8"�HQ#m6�"�&A0D���T�U�1x87��O����O�$�<��Q":I�On6�E8KZ�2�F�D�`�q�{�4�=��1H�Q���?1�'������
�s�BӐ}����4�?�+O��d
>A�����O���O��ܮE��=�+T�I
�x�cӼ��$�(���s$�݄b��'L=>�J`%Q�<zm�g"=���l�Gy������7�N���'��D�>?W��1�M����/1�˦�	���3-�S�g�B (W�ʇa}L��D��&[)^@l�;��a�ش�?y���?��'0�'.�!� �����eRQ8��'f�a;S�i�􉃈��۟ Gb�7u�P���μa�`�F��	�M����?��'U�P���?	,������ܸ4�=p���0p�U��u�K2��';�8���1�i�O���O��w+J�+9�+�'���P  �O��D=��u�'���h��p��E_N�� ��',p�JW"7d�	�)�<`%��	����	�����:e\9:��M`ti� @�Bn�����矸��Gy��'��'!��O����ݕ,X�ZE��
oy,�JѴi�`H@�O����O���<q`'�`N�	Ă01�d�uj�AH�8B�&�}2��V����~y��'�2�'CVIҙ'`b����	O)�T��#m�����Cpӄ���O���O~�Z^�ej�S?��ɐ��"�@ƲvB\�0��Z�U:۴�?�.O����O��D��WZ�D�|nZ9_��(�/�8��d��&-�6m�Op�D�<!Eد�������	�?=�(ӶD�jU���Y~�0���E4����O8���O����?O��O����
^}�5�Z�Y����$�z6m�<�p�J7C*��'"�'���'�>��i	F�Xԏ=g@�c#LRp�h�o��t�	& h�	L��h�'w^4�#ϙjjڅc��(1��oڼ9U��"�4�?����?��%g��ey"�τ&���b �tR�)�> ��7mݞ�~B�|2�i�ON]��m��w�H���+�O@�+B�撚�����I��@�OH��?��'1JD���U-�`�@��6(4���4���Xx�S��',"ޟ��0��EdN1��br�Ɖ�M;�k 5x�P���'[�[���i���&mہ؎�ҁJ�Y�^@�f#�>�h��<,O��d�O��D�On�D��W�\@���N�:C<��0J�?Op
��"��O��D�O ���OX�O"���O��ǋF��XX�tGC�x�Z��T!�k��ɣ֖�X�	�`�IKyR�E
Q6�1f�=1�IS�����Z�K�6��O:���O��$=�I�f�ޅ��t����ő
gt�p�Ú/{�PU�'%r�'���'D�Dڸ3��k?#��B��T�d �T��F�^٦U��Y�	��P�I*)Դ��V�/��4r�
GK�g#�����C$oW���'��\�0r�$D�����O6��������8�4E�&���`�@ʂ�w}��'���'LޙY�'�b�'�Rן�6�
<�"�^�}-��z �}� ʓ-������i���'���O��Ӻ3�f�?((u����y4�CE���I�`�֬n�l@����8�S{R�13gV��T 6DW1c�`7M��%gDaoZ�,�	��������d�<�B�e��4�Ì<5[���l˩H�&-S�y��'q�	r�'�?�7N�$�j�	�h���B
��3��'��'�V}y���>i,O�����2���?O�qR��)T)q��{�~���<1��U�<�O���'S��1+�6=坈p���*	�U�7M�O�بN
w}"^���IPy2��5F�I�  �X��6l
D�uC�#���Q���*?�!��,ۢ�r�g�`Fās�BD�1R����k�H��DAR���PR�N64z  Ĭ		dLҩ�E�Pџ��!�Q>�Mrb���:u ,�>�2��>�Q2���qĜ���=�0�1�Ǿ4Q�9�޲G���a1N�.���Y�>��]XA�ۤZ\����5dF�H@�Қ+�F��b�MB�	�#G��N�!Ȱ̉�ц͒� �4@��Ac�M���P�������T�sݬQ#RIŐO�
isC�̮t�$�
�2��cdB�\*�I3���[غ)!^8�?I��?9�H��(w> bF-fKX�pC��#g�f�Ӝ+��)�/��
�z �PN� *�$�<!�Ό�P(�-� :����Sn���(�b	�7M�Ayu�� �Б妗� ��<1@)������x��C���9��9,?���'��TI���?���,Y0H��ve�:@3���U��+N<�0��W�22����6���tL��<y�
��r��	��O����'��'P����Ǽ0Y84)�i�0>)��D
 ��t
rCO�j�֧�	+��O�%� �K8
����(>m��P#[�8�n8�#�M��4�O?������	�$�ʸ.B���u��*� !��O��D??%?9'�ܫ %�[����+B�\7��(��<D��Ƭ��^��u��`D#5Ւ|!`�'�P����z�%94�:~Rԙ��P(@�N���?�ӏ��ℂ��?9���?������}�l�� �<|�J	�0m����0�)ߟ��$�Y;<� ��h�E���%L �e���y��3|sR���ri�M��I��.����?�=a�&\���&ϔ��.�r֍�H?��  ������'��ɵ|I�	�d�2$ �:aeU�M�0B�	�2yx���1��s1D��`�:�����?A�'H��P�e�"�j��R�|�d�Aŉ5+�9 A�O��d�O��dF�,���O��S%��xo�ş���I^-0B�Js�I�V��036b5�OܝЪ�>�dN]_F��p%T�jt��W]e8������Ob����(�t�"Tj� �����H��O��d�O���'\Z�E l������`�@�B����o���"đ:w(�E�� 4B��Q��	`yb��#�x��?+�p�0"���"��S�e���� �Մ_����O���H�w��̀Fg�,NyCW���' ���i&�ۃ��
E�׻Gtp�Gyb�Z�5�<|h��>�nk��� �@�G+E���Ɋ��ӑ���F剐k�^�$���������P��с�QF44Ic�Ӌ�yb�'�}���:�:��-�Y�!B3�T��0>�s�xҁ�U�X�x��N"���	3/A2�yr��[��7��O��D�|�%���?����?�#�W(em� s��?6����\7բ5sՆ��"3�MJ �5+MIq+��b>�D��_�z����P2�Vt�ĺ��3A^<h���T� ����'lD�`Q?�d�bXL��Qp�X8�@�-R���E�OFc�"~�I���YR/P�
���q��D�B�?	X�j����J���^��"<	6�)���Ӳ&�T1��N:(���#���?���;��"���?����?9����O�.؜|�r��VT��4qyj�ɫ[���@ԄQ�K���cT!8�y�	b$#{a�m8,ǀH��$蕽z����F�+���1��KF{Ri@r�
	h�_���́�l��~"�@;�?Q�0J�r'��ބ�Ԍ�R�q�ȓ ��s�V�����@�)q;\��)�'_t�X9�isZL���F:U��O�K�����'Rr�'�������'7�)Q�zCb7M�O�ՁR�".��(ӠE�>�4����'V8�C�]��T���-T��V��5��1�9�OЋ��'�2�|o`�rg J# =��#�ri��'�˟�?�O�䘱4�?Li�f�<�����'ۘ���ɉ��h@�`δ(��;�'qb������̦e���`�O�&�0 �%7�졥�\����0�j=��'2��e���T>��d��>*=<1@�U�h�T�k-3�E��	F�t"��'��+���OG�e�]��Ey����?�����s�ȸ��D�>v���6h[�[Z!�$��O_)ö]���2��RRa|�`*�$ߝ9FU���5�M�f��W��fYm���Ir�T�J;�r�'��F�rwtUQUF'	�� xSB
�
y�H4�'d1O�3�C�+�!_D��V�^k���gN�!bzJ�Gx���'�d�� �НmHVqү��=�\5������O�)�J��S�=hc䏴m����"O^���耜27V�ۆm�7�֤�5�	%�HO���OR�f'ͧrZBE�d n�`��O��d�<h^j�F��OF�$�O���R����Ӽ���>����,pϬi��lVd?q���d��`Rۓb���ӡď����ƾj��ke,aӴ(���'y!|�6g������(g�N��5�w��{��<`���ݯY|R�'�f�SEEͽv�L4 �`ʤ$�\�'�BJ�7S>)�.�x���p�߯k[�#=�'���b%5�i����t㟑x�yaK�1^�YB��'t��'��A�d���'(�)اq,	@��C5d�l�"o�4h/��8��P�!7���G*�(�󄚉XF��	"57��9c� I�ұ�tɋOYh�EH���$KNr�'�B��%EG�Qت�H��6w�b�'X�OF�}Γ4�����O �M[��W=Ck(Ȅ�	~�'�@���"�\ȹ&+k��PA�'�t7-�O˓s[\�%�i���'��Ӟg3B��fv�32�� 6),m�Q,ܟ�I�L
���ϟ��<�O��3Gn=G?�Q���#a(����Q���?��ChN�cv��ȗ#�t�"�H,ʓb���I某��؟0�O�U�ǭB�������-F ���'��O?�I!^�T�q� &�����1�6����k�I�bDPI�4ȑ�/ z=�0&��3Y�<dq��4�?�����IϷk�
��J��'��p�C��oϐ� ���
^U�d�3��oT�y�ʅ�f��A�� Ȧ�'��?�cl�(^�m���K�Rܲ�H¤8�������V������ȰO��LF���V�$�+Ѝ|~����,R��^�Y�N�?�y���'�x`�cnEp\����F�IA
�'
*Ʌ� �	ެL�g擇@Z,���Tz���I�$W���j'ƃ'7�|�sI b'����O�,��'�7AW���OL�$�O�x�;�?�;u�j�rV�ͮT2	#
֕s��5�y�5��I�<���䅇c�ݨ���1,Ȩ�	�C���Dί!�I)e��?r��B�DSf��J(���'0f��a$B�`Xƹ��)��uٰ
�'���O�d�U1�パ�f� ӯ7�S�O�1�@`x�$�)��	�[,��R��T(Oa��Bd�O�$�On�d۟ZD0�d�O�瓹x~��F�N�2B���n��5�7XH�tbc3<�D��˓?�H`�UX��a4F��VWL<�s�4_� �N�t�}Z��'�T�a��?� �K�ܕ���	p��(y^�|h�"O%[fi���-z$���@1NQ9�"O�Xc4��5]��̈�P�ϸ$ٷ5O���>�5��+b��F�'��V>��`D�e��*H��nBa�ɢK�$ ��� �	�7�F��IP�S�DG�m����S'Œ*����a��(Oxu���G�M��.�.V�	c��ڢ�<q�-
۟G�\�D2u��W�,�䔿[����ȓ�z"�T15Z`�;���9 �N��	���x� ��IU=?Zx�cA�I7�xy�N�Tó�i'��'��m�������@�	�"����3+�'zs¥3#��A�&��,��|�<��On5�[idD0 ډ(���Մ[J"@Ӌ���O�� ���!�`rTbϔݬ��Ԧ]pd��#�)�矘8e
S!G�4)�b�;,��]��H&D��C�L����Ip�_�7ǀq�� Qꑞ�'mNq�7�U[
���Q�����?Y�n�'��Pz���?����?1+���~5�QFB����#DG��yr�_�(����
	#.��2,�h[*\B��#Db�	*���Gcέ�<�{��*�^��$�S��D=peX�!@������?�����I}�F�w��Y� ��ny��K)d>���pcA�8��AC���0<ى�D�gX�t*��D	� |����6p�jl�$�M+I>���?A�'KD���Lg��Q �3h���bՎ���SSLß@�	蟬�ɝa<T�S� ���5�XA0�DU��䪔#W�� �8#��`?�9���3�O
ya���^��eH�aډ	������<��bhO�<slU�S/PX� Zץ�O���_4H��dc�6ON���J�+_�To����'��?!��b�5y�H,��OǛ-�6e�.(D�`��`
�>��*�'�$y&.)BV矌b�4$�^���GG��Mc���?�.���)ŮB�g�84��-	� ����!�)�2�$�OR�d��1x(�#�|����E��YthH�鞭౭F�'�h����i�93:q���P!;�>!�A�=$Q���C�O����O<�D�|�f�͠]�0��z_$�zg��?y���9O�XP�N�?"�'��t��8��'Ol���l"�$�K�4T`=�A=OV���¦���ǟ��O� m�u�'>b�'�9R�)�6��0�e*CVEZ �b뚹�J�zQ�!�T>i�|�I�5�n9c��3i���C�[kܕ�A/(��*M>E���1g���� ,|�n\x�/���Sf)�?����?������rO�,��a�p/6��{Ƙ�I�����ɥ u��8aホ����5 �0/��#<��)�� X{妈:�+Y�}ʤiq�`E,�?��� �0�2"e��?���?�����Or��/,; ����:y�N��d
�w��l�qͷjϊ}��
��J�ʑ�;�Ē��ޥF���jR"��k��u��� t�8�k�(P�"P�a;VL���0�Afڟ­��U��'^h���6:�Zm�S ��Oz"�(��'�Zm���'a��r��Y������lZ�P&�� 5II%9j����-
L��%E>?�ߓ{��ٕc�$E#L	[��!&�����V��ᖥ�&�M{�S�P>Q$� �M3q披)&��@��O}��'jI�?9���?y�2d��$��� p۴�?I@�^?Mt�l�t�-}��1d�U8���E���E8�Pa�	N�Sn��b�B.dO�hui�&$��
V���dҦ�;a"�%=���#��GT�Y�"nΨ�M�����d�Oz��'�<M���Ş=\]+���4w������?iv�G�Q{&L�C�k�:�K@��<)"��$:=�&Z��#��\��u��'��R>�C /W�h���aw��UE|���ۣur��۟���$r�~�kD�x� =�o�E����z��ulo�*��tI�	?��ͫ&�	�P�}����N���'���T�O(Ԙ2�H
���S��=_&����$|S��k��$�O�ʧ)���rr� C6,]0�f��B
�+��?����?��|ʊ��\�8|��nV�5<y@GϨH�a|&<�^�Z���[��Z&@�yQ&����.(�4�n��T�	w�D����'�� C�F��TR �X٘L��kڈ\�h�,˵w1O�@��/S�e�q�K�:_4 �R���!����a֝*�<h�y���'��D��K�.X0��U�K��]	��j�"�'�2�'�?��A��q@��C8��M��Y�Ly�$�Oz��D� 1��㋧�j�D�عD^������۹�~Ҳ����b�2]��	���O!���'4mS�ή��'�B�'����Ɵ��� ;��8
#,�"}���g�)À�ɣ�N����\F��(�B-�d%9�%c	vC�lK@���^�Y�d�+nT�P d�-0� �3ړy���2aʵ:�y��KNH����\����?�u���,O��d�<� 6	H�'@��@Q���&T=Ԡ��1|O��RC��4�<���Ҧ�� +V��I@ߴ��+Ą��dyB%��eM��]��r�RPk�z���8禈��$M�������ȟ(��B�ǟ����|�e@w��1�*^�!��2"ƕ045���W�śv5�1��$Ӷ��<a�aH�LP�j�$Y�֠:E�ʪR�l�1���p$�FO�1��<!Â˟���ӂ�:g`2t���� "v
��I�'����?��W��@ʸ<�-4 ��ʢ/9D�h;g�7��c��!�Lp��Ba�,��Oʓe��C�i�r�'A��i{��Q+���v��2e�@qR"���,��Ɵ`���;��xjR��K~*�T�s�AZ�X5����5(�tm���	[ �,r𥗔X�PlⓥV��Y0B�ۨ,�*훁�")8Ң<��#��������	c��� I���ڐKBk�"B��K*�2��s�T�q��4w����7� �굨(�OB�'�<
,�����	�!ӛ���U�i��X���Ms���?�-����I�OT���O6�z��?�2x�W��d�$9j�d<g���nF�S���d�b{�5@��;vt��7���*�@�:��1�)��ةSB	dm��H� C�=�Z׉�:$��i�������_��?qD��hiÒ�G���s��<�����>ɳK*G�xѕoU<n��[�`�i�'��#=�+�"`b�G�b�)󇋪!��p`��O"�dЬ.F���%��O����O&�D��{��?!�1yOHIzԅ�2u�Qa��a?A���zx�`��A�3�r)cVf�+0h8I͡��@W�5�Oz����4�h��Cﮱ���O�`���'��{bF�(0�
}0!���M]�#7�F��y2�ٴ;��I��@(A"��r�nUk�`"=E��E�La�7�K�{%�!y�U�Hx ��l�3c��d�O���O���4��O��w>�a"��O���4����ô@����F�5b�|2�հ��� 7�q��F4p��G���)M�|����?��H(��{m٫K�\��D�L�P),,�ȓ~����!KW���Tc���,AlX�ȓ'�K�h�2K��$;��,7<*��u�OșѢhݦ]�I��0�OúȘci�G���V'[�Sv%��޲9�b�'b�Z) ��������|"�+�(� �5�X�M�v<*�+�J�'���,�4GD�D�����^<,a���T��$���(O��[��'{r�'�BY>a;AO˵�
%��j�6��3/�<�?E��')���w�G75�U� 5sp�p*���'�H��hM�
 1r"'�4�P�q�'`@ � p�����Ov�'r�8���?!��|�c%��0d= <�͒�i���I��ũ�?I�y*���#�E�RT���	ŊE
�<jP�?[���Fx���'D�Y*J&�<��0�$9��BD�"(��'���N#|�I!{4��Ǫ����ؒ�<���Ї�I�A��H3r,�%�������DXn"<)`�)�R'D$N�u[��ŝ_�6M�2��?)�jF�mQTd̔�?q��?!�]��n�O����0,�IR��W�!D��a4nE/��$�	j����D��A0%Q� �5s74�#&U��D��3)x���ڸ+��HI3"E;R|�)B
Y�[��$ʚ�b�'��'��'��9;n��d���!��"�̒<��C�	T/�9c�%�9��UZ�<.�����4���ħ<��#�#��fn��1��p2�I�9iX��3� 	����'���'H� yq�'�b8�d�v�����R�f��(x���_�1�$J�#_
���JN_X�@{ᮙ�q�ʀ��Ì�*�"hbo	7ق���\��
��<14(����� �$!��VX��r�M��������h��dJ~�K�*f�6�Z�K�h&ܙ�	�'L�h�U)^jn��e׉�0�[�'j<��hO1�`�1q��0 �V�uDT%���y"Or�#�+��q�E�QYc��42�"O�j���ZyZ��Y�kx*��u"O�u�؇T�ER!!�~G��9�"OFi�N�&�����'U�У�"O>���شI�	��̥v����"OBİq��13��Z��Y���y�)�2Ǫ ���
72� �k�P.�y򡛈v��pi���*�P�$����yR�@3��L*c)X�P�P)���y
� �]`U-�Z�8a_�nօ`�"O8��7 Wei0L�ω�urj�S"O.LpC��X�%�/}��E��"O�h��u��ِD˙�7�qc�"O\�ꖮ�>;t@F	�q��"O�8�C�ݰ��C�n���"O��Q�Hۨ^�
b��+>�8�`"Ox�ޕl���g/��
�B�R�"OЕq��1 ����hUC�"O�av�Ǥ5���i����Lzcf"O������9'����</<���"O��G*�u�,M�՞6@
b"O�q##�59p60���v��|�$"O  �G� L���䠑L��9"�"O�I!d�ԝH��A��eI8�"O�5C�ȲC���ua�w+�x�&"O��$��7�6H9a�R�U�d"O.0cteȸ���Ǝ
@�U�p"Ov�Dע,S�#䌌h��	Si�p�t,�6͑��������j�Έ�p�.�kD�L0�#\�z�bع��n�a��O�aV�M�Vn����ñ���MK� 	�<).O��(e� ;�X\[x�۰�>y3�����$��+͂<h���&�v�pҥ��nH	{�>�K��G�E�xѤO*��ҥ�]"�p��/	�$'�px6��*h�Z �!����!Hv���p<�s��Q]�Dd]�dA�%�6	ۡ{G
 �H���tIlI*Q�̓F���D��e[:�{U)�|��Pk A8�L���)(�����٥7������Mc�E�=��t���0�)�����t����U�~ �3�ȦG� �:��Ї0cNP���'G��n�)
]~�B oƦt"���j�C@f�C�C6,߾M
�O�8B�+�:�A�reC"z��Q1d�d;� ���<����"�:�Y�HI�#�2	�6NY����G.ƶ

@u�oe���lZ�5����A@�[fT���fi��q鞥u����N8x���r�P�XXc�^a�'�����,`9�b��8���*㈘�
�`�X�
�3n������n�1S��YH�2BőQ}�O��\���Y�5P��6a�<9��'��%[~��DMqP ѡ���#f����/��� Y�L�{�.X�<�(�S�S�808m��;1B�����;lq������)W*T)�k����J�.2j��S� �n��!�NZz/b�b�P��0���3Z��9���A5��+s�E,s�̰9�-�9�Dʊq� P\A�̐���'b�R)��Dڪ1n�!RXv�͒���"JB-k�e�:s���c6
ڝoR4�3͕� �:yS#�"+����)U3zS\X	��p���G} �<h��`F<B3�P��W>�yb�)v�`�!0��>|䡂�l� �G���@��@��X3�PEp��M`�
�C'#��`��3G%�O2E@\u�lp�E[> �D��cM��PC`�SԤ�ATB�m9�	 '�6�'pSb��w̌L)��9R�`U�+�_��Y��z�EablZ!u���ZA
ʠS7�z�I� ��Y����O�L�B�R�!�
�B�"m��_zD�`$�	���R�>sV�г��86�VM1�\$]fQ���7o�+}��a�c�4��d��S�:{���G��M�b ���)I°0;�"�~|���p$�\|�� �c���F~�gZ�5z���Vh�,=���� �������vȫr�V�@0�=����9`�Pk�b�ܦ�
��'��4Z���U?\�bы78�iK K��i�N�S��'d�$E��0t/�MC��'�>�q�Y��,,s*�vy"����0ͫ$��ٰB	ï�M#��l695(H�C~.E�0��O<�)��'�5 3��7S�u;ōY�V>`y�$I	`7mK��?�P��%g0]��) �k���a��AC W m��N�/�jT�A]������қ��O�]�ѫ��Ib�E� Ǩ�Za/�7LP4��
�;/c�C�
��i���?1S(ݰs���jE�7���9�hR��#%0l�!�F� W��p6(X^��	,m�j$��n��IB�ā2K�6��F�G�k�F9T���u��7��t`�c�^��g��(�J�xG�\'�v,�`Y1v�x2�8��D)䙉�E��*��c�<բ���D�7*�8������O�8��Z19&6�p��4}P染��>�5Q�����16�$¤�G�9z� �"��d����DG����6M
?>If�E�>C����!ѱE��R��-�%rİ3� ��I�B��V�x�� i�D��g-�L�2% �!�7���yjS�/V�� �(u~��@�!M���Ir'��ɥ�_g�(<�M�r��>Ʀq8V�B��Ĺ^��h�S��J0᤟uAi�S�䚦�)��<�ǳi( ��j�S�� 6m��'x�x"B�F(�I��S�$YѪ��CE=iЀ;�G��U-���RDKLJ~�G�> ��!�I�VK��IhR����*["!�d+~�����߄La��i���7����>9�M����f����剬&K@�z8�dP)�+h�e�� b7f����ɮo�eT!E�Ɍ}�Z!�$�*� ؑiF��F�Bu����1:��y��I?i��<� �RM ��Oۜ]8B��Qy2$K<3��AhWe�3_��	�D��8ò�17'�6��9�'�e�ajFh-*�r�#N�?��O�:���y܀Q�N��i#��`�����8� �pI�vrџ�Xw(Y>޼���O&C���#Х�GU ��ś9m~d3&�OX�9��9O��P�.�9i�l�`�B>�x ��/Eo��$��J�L��T�����U�q�� *�C�a=�E8fJ�<E�R|�ԧQ�s &b��k��I�f1rQ曀AĬ���D�L� �;��_�^��O����G�/��JJS�2� ��Q�� lH0�v<�3G[5|" �b�~�ʸ�Bo�S�>uʹ�Fg߳x�T�#
�F?*��'xt	��J���&8��́4Nb"��O��+diITa�#kXI� * ��(��F��dU�9��'���~ޙY���7Ap29ʱ/B0P\Sb��O~\Q�/��Xs2B��a��x�A*)l$BA�E �:@�V���]��q��O00���r���~Zw�R�J���@�U�6�U=+�,I����;ԡx&@�'�,�Xƣ��T"Z��E�'p���k	�f�R�jaN�Q ���ǉ�uhlx� �d��)�Yܘ�1�ߴW�Rx ����U�DԈ�P��������@F# Ձ���/(tx犗&b��1�ө�4͸'u���Pb��|F |C�˓<4yS�ѯ*m6H�e ʧ=����Kp@��$U�T�N�pcF���)16_FB����+g�vE����V�pA��,E���,�Ԓ1���v���l�5b=B�`�gPYS�Y��hG�ZI�\ �'�v>�Ց7���o���|�Fl�'"w��3&[�8�p��S%(D&y voC�$��o�8~8t��ɤ81d�c+��U��V.0o8L�G-6��IXg�V>I��dB|��y�����$kN"/��;@�ՃLK(݇���xq{��&"0�{��-�vd�ƀ�O i ˪wk|�� kO&͸'>�m��/�F���	FņsJ0qH��
C�`!� 5Fax򈙫 
�T��(0��n�	EP��LQ�6��b�	?L"� �!"�	Q�Ł). 
���g�6���'V�M��
�B�zԹV��n^����O���w��=O<y Aϒ�I1�@�ET�p��-kj�ű1��FZ�35^�+l��2��[��d�������1n�z��$ӸZ�dF!�az13�M�u貌8�)V��2�p\���0收xنP�k�a�;��$ᰬٟJ^���I�e|x�gA?�O���B��o�$Ԃ$�@	"����[x6!PJ�'���J�'��;A˒!a��܊�C7i�d P�HQ�EcVZ�'�f�;��'bp�KW.�zk�P�CoN�݈�C5t�N$y%�	,#�Lce����',������**h��J�B�3b�F��J��P#`D9v.\V#�n��M�a�*u�Fe�g�'�� 颅Ϥ��˓K��b���� M�s�MR�n�b�,܊�i(O�Е�5O�ulvQ(��ҍ(�x�$T�Z]|Ӗ*HP�<i�n��,D���4�=)�j��RDȤqe�R)p�r���dט2.f��̘��=���Yv6���� n�� Rg��
��\Is��uܓz�$Tj��Z�+������<���ZgO�" �ι �+��Op����)�?Y�Ǝ��^�qT��k�-R��H�0%DgƖ	;C�o�%BΑrţ 4H��'!ҴP�%�x"!i��'g@ip+A V([J�R��{v�'7bdh��!t�D�c����ߵd��}���y��	�!��\I�gʗ~Q�9�CHA�'� ��;)�N�9_���qw �EqΜS�~�N��'9�)��9z|��@U-H(R#:�P��h&�E{b�?{�PT	�ĨN�TA)B,��?7���&�Q	������P��&~�z"#!�4��s���*JR�J&�Ū���q� NC��I����<���8G���3�ሴ���I"��O�"<Y�/�x����e��^��d�,J+ɸ'��@���=�`���k�x�8K>�Enۜw��D#@�[�GP�qH�G��d��{�C^,�U�?�F�ԗj����>YrO�}���r�'��;��� �%��ew�=��BG��	���_-�hO@p#8�9{���_8 �z��ϯ.���+$�|"�ߏn���) ��S�DƝ[Uj��?-�����8��b��9I RUx��$�%1�0�єL��!#P�J�����$�����J^:zb�问%mi0�
���8++�
R�@��O䤡(��>iQ�.O�Tq��Z�s&N\rԍ�/(���P>O�t:c��]��
Y�Me�Us�K�7.�O�� g�6/��Hc�ʇ4�c���x�H�O,�s�. ;���mӲW�LY���xr�6)RIK��-h  ,N�+��m�*��P� �q���'.J�O��(�K�{MR�)�JI.J��\�&lبB�5��,��b,��p���(O�$4��PrM9!������o�U���x�n����b	@����Πg�y��G����D�XS�xRH�y�S����� �-�J1��[p�O��*��<����8�.����:x^.��p��az��1�F��S���v��]`��>�	5��(w���	�!����M�iԺ1VkG������L��c���=)�o
�.L���UfQ
l��<Q&�A?��Ȁf����məo�=ڰ�,��j�	�L_���?ُ�IE/H����(�P��"ԈI=҈�`�@؊���[�B���KU>︧�AZI\T8FdFUK��:Fa��V�
�O��8Bi#LO�|�a*p|��ϸS-��j3/�_&��{*��	G! �1'Zɋ�ޟ���!�3��0ҮX��@!�7F��b!:g��/cm��(��O����@$g��?�KR�Q�Onv�s������D!u�t��n��q�ډ+��[��R�I���O�1`��z��8�"eR�!�j�i?yC��7iȑ���	3N�Ʌk]��<� l�:�oJ�d�kwG�}���֎Cz��$��6GqOZ%��O�b"����s�A��]�`�ӳ���d����P?g��y���}�:�H"��)��g�S����_��㢎o���C�٬�Q��8T��y�ᦆ,/-���&���G�/�5r�!ǕXX8��rgB�]��n�S�4gJ�r]���S�n��$\�f�rx3U"!���K�恘YVµ(�$��2 ��H�t���a-L�&Er�T>�'�n�z�%I�&8*d��������P�'ݒ�k��R�KZ�+T�[,%An�x��d��@��D�E�:M��!���2�f�I4ӄ���H?a*((�4irˆn�����4���LB�Z�X� ��PFD����R��1Or�ADR9�yw�8T�V��Q!`MzL:��5w�Aeg=^�` Ҭׄ
�Pa�Ϙ��	�.Zl|0���lA�����	
$`�<��
��|1���:,�c>�wO'1Z�ej�̙�O�
	�'Mª0��u��T>���@���G��<�X4/퉴�K$�`�T*�*0�Tw���K�E���_?�~��D��p �։�>(��3T�@��0�sdH��~e��*�ڄb��c��@g���	C�$�)g�p�)ׄ�H����y\�W�6��H��&AI�Z��%�	'p�iW��D�s��A�7A��zX�)Q�d�Ţ��)}��� ��I4]p�Q�D�E  ��;S�XQ*�-ΐu)��""�����2a��Z�[�J�b�h���|F|���c���H"��)¦�`5�?;�剄g�d(�v��6~���!��H>���D��)�XL��ן8=�U=x
I2��ٞ�h�AG��#n�X�A�������[���:�~�����'D���j��SO�98Cj���#��e����`�az,��Q���~b���;\�8 ���rw�Mb�fm�<	fʓ�L�flÁE1�'��R�mS�q�~��,�[���r �AU&��0L�i�a�� )��,Pm2�s�0#�/�&
Bݰ�k�\�@��cb{2h�d�>��� H����A�bO�|q@�Z>���W-��8V�7G���!��Z�;U�ȉ'HP�!e���+
0��T�U�0h+��?���+�HdY��I�	���%=���[��X"f#�){�\����	m�Dj���� "��!���څ�~��P��,�4(_����äI��0=�'\���'�fm�SaH�N(��� d�S�{b�L��(	2�S�d~Fۖ�F�s�}�c͜�G0\��b��C�S�7)tY �N
<x�5�R�ۈ0sNC��70b,���"�rD �X#Z*|C䉡o^����MǬM�d�����/��B�	��̩c�.�b�hYSŜ�%4�C䉙g,:DY�e�>"��sS"ז'?�C��\?��Bl��!p1��)2pzC��(�]A�(ʭm�E�$�Z.�C䉌8�L]�p�_	:���8en�>B䉕<a̰dMG,3	ReSG�PyXC�	:u�F�A�(�&
*&5�d�Gt� C䉈O�:�"%���� =�W+E�21:B�I"b����F�+ځR(�/P B�	2-�	�U�<@&^� q�Ȑ�C䉨�"l����3l4�{Q�ċS��B��*/8Px�ƍ�� b���cD�K�B�I�<4�	���!(���A����>C�IvU h@G�WU��0E/W/ErB�I7_�}S�@'1����T%�B�	2mwH�P�ث"�t�	\z�C�ɵ&n�]8rl��"3~�S�+ʦ4�C�I2g})U�ȪE芠3�'H�in�C䉝Đ�b	�h�ɂK�Ks�C�I�E��������{e&�A�\���B�I�.�%k���y��Жf?ŖB�	\P�<Ya��y�4��G���tB�I��9�7��G�h!łH�i�B�'@.։0��
������ ��B�	't\�� �@N&pܼ��O�rB�IK;$��
�z��L�U���1�B�!�~	Y�֬$���s�%=BH�B�I�3
6��]�dp� åi���B�I#a�H8��M$$F]�� ��hY�B�	�P�,9��A["�Ih4➣=��B��@��X
�����: ��ێ�hB�ɃN�nc��^�(�█d�C�	!.b��y��J�D�f�w%$Gh�B�)� �)�4J��(�q�U��#w �"O(�;wIDBH�H�.[�)ZV"O�#V�X�=SDt�T�O��D��s"O,t�Uȁ0d3§F�3����3"O ����F�u.F���G�j��eR "O���Єe�Z8�w�G�\�:u��"OH� �ݒV����(��R�)2A"O�ё�΄:j�{0�ۂ���;S"O�����	�A���Ig4�e"O��0���[�|�"�$ܘUTB�"O���6C]\�,��Ϝ�A�v"O^ȑ6O�>�.D�v@	cpM"OD�`/�5P1�1Yf�(YR��9�"O�����7"�`��Q�F� �"Oօ��/�\9��	�: ��� "O %��둡@�1W�3"����"Od��ƇA-fJ�&A�7;���"OR*NF�P�� O�}�؈3�"Oƅ1W�^�7[*�ɰ�>1�\he"OJ��r��9��I��E&8���a�"O舨����>�Hs�LG�#�5��"OP�s�G�r ސ)���;s��0"Oj��a�A�w���;�Ф5n4L0�"O��:Ԇ�,QD����
�mN��K�"OX�2�l�	I>�8�G2mHB9av"O��J��	C�#��E��`�[�<q�D�)%ٖ�0�	�H��I�`��c�<�c#9g����o�
����p!�$(`?��+�&� V%�(î�\�!��!]4�x�@��2!�Y�mH!�:VijQ��H�v����5��>;*�}���`���c�6H��j,�f��k-D�a��5��tB!T�J�	!�*D���N�>�T����:qq��z�n'D���,vN�ubd�9d�"ͫd�%D�����x�<S0
�� *�495%(D���D��$+u�ٻ��W�B�ɘv�2D�X���[
��@Ȅ�ԑJ
>#��5$�X�6a��{�����Qiޥ����y"�ا&偄aP%v��p�A.�yR�1=|�v�Xh�m�����y"��u�T�Y�E&Y$������y2��I:}x�i��J�o_��y2��sp��V�j7��%�T�p=�}rCS�V� ��ȤhE�U2��ɒ�y�D�?� I��	��o����%��y"�)�~\0�c���D|��9�*4qB��ȓ	iH�û)$��M�@C̦8�<��ȓrb�Smɇ;���p�R" 5t(�'(`�Fy��)�$ǈ@&̷��0k�M�"7!���	�|`�e��^��|��A 0!�$�!&�^ rV%�Ib6�k$��M!!�dğ8�Jl�ck�5YHj���f�11!�w��5#ϋS�4�)���Q�x�"?ʓ	��@�`��M(n�%��)V���;�8��Ba^)�X}���̥.<Z ��^r���3���\:�@�S�لȓ���B��Ur�����_hQ��}�ذ1煐��4�F@T��9�ȓM����
 "̽H���#I7B���H�zB��`JD-�]F_7�`������䆒�u����J�8��e�ȓl�|%��f>p2���׀O�g�X�ȓ&>��ҭ��>`;'�ԴT���S�? �����v8��Q�L�MɌ�H$O:�Rʚ�q��`@�</n�U�v�"D�9��\6J���r�
Hx1�t�?D���ܟ�jI	� ՜K�B�Xwg=D�$C��G9n��H�:Mb���(!D��1a��;L7��2D
	I���Q�"��ሟ�����Liȭ*4�7!Z����"O.��E��31�y	 A��h<���s�'[�ɤ2Y�y�1	
[�4@��E�/��B�	�X�a���ߗU���3�C+rm�C�I�YͮxB2�֘|[
�cł�8��C��]�e���XK(T��'�	��C�	;CR,����[336�m����E��C�Ig�<r �+ǒ͛�E����	>'�ɇ�I�	
h�"EIT���ˑM+p����!��m�w�H�cK�Iu ��CIH��q�p=���C��Eif%I�$�|�S��$j��"=y��O~���w�ҵ/� ��!O�D�rI�
�'�H�檜1B:�@pB'7D� Z
�'p)�E.�y"���.U���	�')l x�#G�?A\k��%���X	�'����GOM�S˾�`�>�.�
�'���!&@ŗ ?�e�&�$`�r���'�:�0t%�Q.H���KQ�ZDVL�'�T���cN�9��=K@A�=�]c
�'��e	l�1������
+Hn�j�'����/v�b�&�
- ���b�'g�d;g*ǎ;wʬ�$�D."�89�'}���q�{P���C��k�t�q�'ب�g"�F�B0ӓ�9c�4�y�'�>�#Q�
�l�l0�#��-u
�p
�'�n̰��S�i����
@�q"��'�Ƅrp*��=����5DX.O,�=E� I�-N
�yc#����z O��y�f�<���""�L�xR���"�y���8~�
��wL�{q�m�V#��y���~oF�*vid���e���y�FR�d% �X�Z�ӄO�2�y�@<1Z��
���-A`�dX�k-�y�h�8w]|��b���oN�<YfAJ�yb�>J>�p���eU�[�N�y�%��V蹥�V�)T̫��y���\�	a�C�)5���!+ٓ��=Y�{�/P'n����U+E'2z�C����y2�[)R}V`�)*B�;PMZ�(OX���E#��T�����}�b�Pjp!���*ˇJ���጑$9~��ȓ������� �b��T,�`Ą�Y��JV>56ݪ��B�m��I�ȓj�j�RBN'/p�(3��}�z�%����I�g"D%� ̛^ �Q��B�9�v%��#����̲&�1\��B�I9(��uF�4d��Q:���`�����-�Ě)
��1P�͋�'��0X,�!�d�C��A#�-&�VR�l9c�!�$ŢJ�P�B�ݚY�L��w΀�!��Y"0�U�D�Q&A��dˤ� �7�!��$P�Z�I�m��`�)B�7�͇ē ��B��Z���I��,�|]��	a�:m�]�mN)Es �aGАfȓX2�)!EO�
v� 1��&XT���ȓ.��C��ު�� �'� 1pD���IaܓF͂��Ⴈa�N��� �P=�ȓ'�r� �k��r�Ti3㌪"k�=��S�? ���A�EU��0�`�
;����"O�eba�/+.vEiA��,y�1"OJ=0P�K|q�o8Q"O�	�LK�&�$aA��ҡ�z��"O�{p�X�8�x�R�M?YC����"Oԁ;4���N�^8jD��@)����"O�l���VS2��T�C��b�"O�LkU���G �:G�<N<튵"O�� �]%s�"���M�;g�
� "O����4�X�%#�8r*���q"O<[�KП&�	b�h�r)�}
�"OhР�B��;H�{�g۲+<9v"O4�!�W_>rmAE@�t1��"O
�XB
�|K�XH�Ձ_�,�0"O&�hGgF6��X@��۴D�4���"OX	R��S)�y��S�xPFb�"O�����	9Y���&	�3r�p�"O.)����12&`�_%O��]�"O��a.	8|^8K@��I�J�H�"O�3�M_bb��fD���Y��"ODݢVneOJ�2í��eǮ�'
O�7$\��I2k],��(�K	O!�P�$�T)����.�:9�6̉"3!�d*3?&�I�j�*Srp!�Aċ!�Y ?�N@z�m1j���D�B0�!��_\��zU�
>[c�l���*�!� �L<�c�FR�WH�m2��ϤCX!�dH-o�Jh놅�oC�a9eȅ 2U!�D�|��2P�z94�1�P�$!��M-P�I�ϟL���"�U�/!�Z�#6FE��fͶS��Y��䕃i!�ā�����F�](�4Q���&!��A�#���3���sNԲ���}!�$��~\���ӫX���2��O�!�C/�f�NbvY�D�x�!�D�1p�V�rb��z�.����C��!�d	�Zl�R!��$��X+��A|!�^42�I:��[_ε%͟�=�!�dRW��)AI��W�|��,�av!򄁽L�zA[4H̺jN���L� 6m!�d�%R�0Rcϥ$9�-�-.�!�Ā�xf��#��19��P#�G�H!�Ѷ	���9�K��V�<M��
N)'?!�P.IO,-q0%Y�vhxI�H��z!���-�`"��Ϡz���H�&��9�!�䜕ys ���M�F��4�!��^�$�@�1ϓ&n�e�	�y�!�d�?;�zd�X.����f�-/�!��"�� ��Q�N� #�8]�!���F�D�媛�7�f@��R8_n!��V_�IҴI�$!���"�$��f!��@�o^5aR��"�X��b"7S!�d�95�li���	��P�A�A�IO!�d�(|v͋AG�?�Dt�� ء.,!���F�����h��K���iY�\�!�$ʕ&m�@����a���g�,	Y!���*-���aG�	W}����DW!�d���e�VCT���Mū~G!��)n�0�%3�Q�S-E��!�H:(��`Z������a`�(T�!�d�������L��n��)��AS7}�!�$�y7����^>���%�+�!�DW����EY#D��P�(	�G�!�H�MH:�{��2��a���e�!�� P���o�mlX@�FsvL��"O�����d�[d�Y c�}A�"O�JQ���P��E�\��I�"OX�ֆ�� 6LK�˚,@h�1"OX)� q�Z�$ǬO%Z�"O��zU� �g^Z�8�l��r䐱�"O
���#G(<N�t�+��5��u"O�@Z �Ǹ����'+��i����"O � C��-�p�5x3U@�"O�1�B)6nR-Ξ�b"�ZU"O2�r�*v�<���+�=\�Y�"O��ꢆJ�� ���$�#3��%) "O��xa�¯%k���a�r/Bm"O�-�dȚ-��� ��%-G�e[U"O�l�g�__v�@a��R\���"O��M��'�|1�B%��}��"O2$Ygj�~����E�[�̌��G"O�E{UZJ��V��nƲ�2�"OnhKBD��Q1����O�?��$*�"O�����/2�=��� ��1�"O�(�m	TP�cI e�����"O���b�Z�d V<�"	�)=�J��T"O4|R��"#����C��n� ���"O�L�Q�ٯ}���ٺ,{�Q�"O ��dg
O�d@���co*y0�"Op��r��f�AP�̄�PlA�f"O�(LX�"U��R����Q]HҐ"Ox{������ #l�40���a�"O��p7L͜z���"�\06��\p�'tx`�䇗/�4�u�̧M�:�Q�'(El'T��A`�@��q�
�'����BA���AE��:B�h	�'����H:?{�b$l��5�P8�'8p�eA�hptyCDF˛1��,`�'M4�0���8+��P�/�+Zt�K�'�������0}��U��-z��Ȩ�'�&�Q M;vsS�A�w�(��'�n��n�:r´��eG�%D1��''��HV��F��P7�Y�$��u��'�dP��N2?��=SV$�"����	�'1R|*��<q
���[ !ڜ11	�'ϼmrR��?6h|{Dʺg�'�f�HUN�5����4%R��@�'nR�k��'mt�C��O�n���'�(A
�CUu�2�IU�t����'S�mZ�,H�x(���JC# ќ%�'�
���l͹�p��ƤV��Dy{
�'0J�!���B̍p�"ʰ��'��it ̈~��<�%��/J���'S|�p0X>':٠�� �n�X	�'����F�;c�Xh����i�ޥ	�'�*lc�B���8�`�g�>/���'w [ N5�`�sH����y��'{J �A"o����%��4�#�'��t����|���B�W�2|��Y�'�0�QL�Wl��.��,��'^Э�ek��y���ff�9���'����8�fq�Q���L:�'_�"`�F0j�$���S�|���	�'����_E���R��ݛaS0��"$D�LP�I	d~p�����=�:�ɂ@ D�t�c�C�;PWw3L����{�<y���.0�-t道@�P��ץP}�<�C��G�ĸ[3�N�4��l��{�<� ���g ��T����,�0~Ԗ`��"O�S��,g�C"n���X@4"O��Q�d�.�a�M6U�f���"O\�(Rf��!y�$� F(pu�""OP%� ܕd�ƨ�`^�+��yD"O6$�$�y:ش�S/��w�́�"O�['����pt����8XN��"Op	&�7M��:�ź"Q"M�4"OZ�c��p)��ea�4��$"O��1 f���P�.��]ڠ"Oe�"�k)F�3�!�4��iu"O4���I0�%j��7<�\�)�"Ol��1g���$���C]��"O8��b��e�2�I�;_hÐ"O�u��ξ<��c��]�wU^���"O�\�� 3�	���l�lp�f"Ord�ыϨC�"�P%`���""OL���.G�lT����ѰF���K�"O8c�=���! MS��l�"O�AЈ+
��Y�5�����5"O��:R(0�c�Wc Z�"O�)��"D�b���B�8kL����"O2���Z.�^Q�� Y|@
�ȑ"O�d���K�ޜ+�098�"O� ���~�  :�N=a�B}A""OZ�{Ï��3�NJ�sḘ�3"O��b�|T����<�x��"O�0�Rj
�M��Z�,`I3�"OP8I��i2��7YYl���Wr�<A��F�p3"��N 2�(��6�z�<A�c�V�A��	kj1��f_�<y�mρ`���$K*W�t�r�J[_�<�v��!u�X���%3�R�N�[�<I��-=�9!��B4���f��[�<1 ��7��l�s%���`y����Y�<iSn��d�r ��P<3��H�BYm�<��H 7�����f ����E^�<��m"Ttq�!� ����Y�<1��Ȫb�:��	���}xuO�X�<9��z�b�16���PH'HWS�<�*:��	QDI��$��@�W�<��d�SW�"7. S��ZƣN�<�B�D$sP� �Æ?�T��(�J�<�f�[�|��M!�o^`��&h^\�<���@�	X���%l�\�0e�Z�<1e���(���A��/ =>�9r�,D���0Ɩ�xIҡX�J�����@�6D��K��ïm�R��d���Yg�%y�m6D�t��8�����A�.F�̐��7D��)��Z=1�@����;KJ̀��6D����cL�k`��aD���<�Á/D���rO�X]~���Ň	L�`E�6�'D�����υ>�إ-�O���##D�d҂b�-:s� �E+��J�̃�%>D�p¥(��c���P2�+�H6D��	�V.�x\��"L�4�.v�&D�h[��q�ڐ��F�yJ�Y
��%D���D!�,5Ta�T&�4>��	j��"D�x��d�3�$i���@�~�Q�2m?D��p�G�l>|�Z�ǟ82��A��;D��y$�%q�<�A��ܹYf���o-D�j@�T8���C��8� �|�<u�&Y����&׹2|��p���d�<�D�r�yJǊص	�틅VX�<� ���	K���!�n,݊\�s"O�x�
�g~�(:&��;%�d�IE"O��x��4�:�c��K	<��5�F"O�-W
O��n��U�b�^�+B"O�K@�΂,���EB*t�튧"O
��u�L�6�ɢ^?�*���jJq�<�É��"�@s$�I��q) m�<���A��ف��<u Zlrm�k�<��	r��I:v̐�VI0RPG�g�<�0G�BO���D ���`@$�]�<	�+�'96ыB�F�f��� \�<�Ӳ�A��*A�|0Y5 ���C�I�v�f����6|"�hK�#�+/qZC�I�pފQ�%

:˒(:�a�i�2C�1k=���,CFzT��E��~:\C�	N���B �D�>��5�6m�xB��<R��0��%}�<���N�S�C�	�0?Fxy`FN/�:LX�;K��B�ɮ��|p4��l5(�3�ȼ~B�I1U�r�q�� e�%'��FelB�	5��y�@��]�vQS:puB�Ɏv5�}�&�˫&+�YB��E�L�C�	�~�@9෇��d�s��f}�C䉯��1�!�&" 6��"X8��C�	�� �rA�2��t��U�\C��9=7.����?Bs5PFg�  VpB�ɩ~H���S36��`��\��B�ɘ2�H�Ti��:��r<C�	:g�fm�Bț$��9�B��F9�C�	�d�qD�'6�0"��E��C�Q�P!cp$d<�|�*��?T�B䉧5L���E���c��9a��C��9z��P �JP�$��t����/�~C�I1�4�YQ��,��ࠠ"ǀ@�ZC��fق��B7�İ�PA�u�hC�I:�}�6��tä�AW&R,{E�B�I0av�Y�2@�47@��Z���2ӴB䉅$.uX� ؂�vEs��N�f'�C�P�½S �0�����aɷ/-�C�I!����"Q�b\����z�vB��),�t�����s�1@��R�4C�	�K�����E�M��D��#�t��B�Ɏ(��[1�P�5�������nT�B䉉:l�� j��w�dXy_�Ш��"Ov��s	�:0�D#�Aæ�zM��"O��dUQ���Q��dcnm2p"O�x+���L�T�:�H�efջ"O<��N�6@�P ���p��"O��X��>q��U�i��N*�8"O��dfK$����'=n��#"O�t�ٜ"�^�;�FՄf�h�A�"O�)�T�YHm��+��ye�@�w"O����C<M"p���	D��!�DX&U^�������0�k���5+!�d��pG,�x�b�8|��e���!���;�8�ɷɁ.E��&�@?!�U���$��o��<(��$D�u-!�]R*Eh���j�읢��O
M!��:�@��$	���pd�! H!�D�^e��B1<r`�!�e�%3!�Ϣj,�b���s��ɢ%-!��5S �aroH ь�YE�A�{!�$@BڎDQd8?�ެ�Gݪ.�!�J�Z V��oN�E����%E@�M�!�� n@s�5���Ak\)/@����"OF����"u�Jed��8%�8&"O��2��S
G�b�[cK1c��7"O���@�<@'z����'(�"OF�`OȌN&ʩ�D�_�( ���c"O�HKuMW [�� �cՠE
T�8�"O�0�#OJ�.�����֡x�xc�"O�m�D�+/��t��ƚ�g��p�P"O4�B�J��,�$ �����"OXh�h�4��(�f%�+��H�v"O��$�֏.;���f�$s� ��"O((�#*Т!¸mX�E��6۰"O����N�(�lA�'&�	�!�"O0rS-��[o��Ř�>3�I�"Ob�z G��z��҆��b�
2"O��S,����p�^��t#"OR�ڀ �*q�T8�S��I��8	�"O`���>��Q��/z�\|�"OB�XP�����3%�]i�|��U"Oƹ�"<`{�1!&F�3{ �B"O���C�� �d�:���b�̌�s"OT�)�e�6!�Z��1c9&ĺW"OFe���$���!te�t4d���"O^آ���>���̈́�U(�Q B"Ov���ָ5��d-ȌO+��ٵ"O49+E�3J�MJ;�$p"O���	b����T�^�,d�'"Oa��""��eH��F�!�`"O�@� ��G�n�{�a�4^R$܀�"O��kCAW�Q�����6�H�X"O.0��(sc�0�'](M ,��"O\��K�g>܌���۫5 �(�V"O�xZ�KĢ$wv�+�)О1Ơx�"O�\(�.قj���1�	��{`���"O�P��N*x*p�Q��<)��9"O��Y��]��ӦX�W��"O&��Bϔ)mr�-U��m���	��y�D�i�I*2@B#}30���)�y�
U6��i�m�%ۤ������yRW��y�D�)v����J	��y�/��p0u�b�"W M�͋��y�,=;*DqRI�6t@B� �yRGK�,)~��B�Փ~�<�`�"¦�y�iE����5Y�����ă�2C䉮LP���?*��QQ�%�)R�B�I0f(�B&,h��Z�-[#n{�B䉭z���:Ia�5"����L�pB�ɒ8�̌���G� c���5f%*$B��Q~l������* �F��C��+X�@2��]!�Q��ݷE��C䉬O�#�I�V)^= P噣EܸC䉘5��G,R�|��+�*����C��j���Sw�Х�DK���C��l�T�A�C4q�M(���6U�C�#5� �愬$�89@�EB!#��C�	�CP�8s��3uO�����ޙA�jB�I�8B�HT�T mJ�@�X�.B�Ɍ�
ɳ�m�/S� I����|`(B��s�E
��(<+�[&e�24�PB�I־����+m�L�0�ڐX�C�	.J�Q�F��.�A��8Mr"B�I�mN(�ઐ�ne(��4K�	�B�ɫC��:���7%=άx�oQ8�TB�	�Z�΅I&LMm���9C�$V�C�)� �X�qhY�'��Y�R�jS���"O�-I�Kوu���d
�FC�Y�U"OF�����
�:Q���΃ �Y{�"O.�j�^�1
T�Ȏk��e"O�� �m��5�rȓGD [.@HS�"O�Ѳǎ�3G�N�*V��a`��b"O�L����"�F�2�����H��"O��QqCȸH�N���ŉb��@"O���c�� DϰXB��Л�"O���4%4���s���,��S�"Oz\�"�T�CJ:��L��L�F���"Olʡ��}��5ɱ��o�d`��"O��xb�Ԁ,��V��0_��ţb"O�DZ"��,�֍�����6"O��� h@�l��QS
Y��D1�"O��r�	�6��C�S2H�l�"O0@O�~���sb�o�ҡ"�"O
�%�k�4MH��U��[1"O�i�R�P�O�ʝ�婝+�IH�"O�]{PA���Q��-aR"O���GiG(g��j�fL�.���#�"Of���\�=�k� U-X���H�"O�1)DMø��K[u��`1"O�F�&h��hXe��%nN`	��|"�)�S�M� ����$8�ā'�K,/�(C�	0�j 
�
a���g�V}�BC�	&\؆�{�S�>�ʬk�J��K��B�	��$�#KT�=�j�yTȋ�B�B�ɑrf2+R�V+m����	�C��H�m�D
��J��G.�*D�C�ɲ]񘴫�`��V��`qu�C=�У=�Óo6�Q�CƐ-�6�%DR�[��,��(ʐ��c�-
��%"�Bۄ�F��ȓ�;�+T�6�x bU��^��܆ȓD�,�zA�:$��	�ᐚ5�~Q��o7F�bLIt��+��X?ӅLt�<1b�
9
X)�ع=W�,a1I�o�<� �<r�G@ܶ'`�� �Tp�<Q0蕋1_��F�	��"�o�o�<��I�85��I[G%͒y��
r�g�<�3BL�V%�$yF�b���eb�<����h�����J��F�欛�	c�<��eß9<�,Kpb��*X��B�e�<�T��\�N̺#bZue4��]��B�ɁE��=��@J)�8�S��*	ܰ�ȇ��16�d���J1�(�r�۬XK�C�	6}��Y�2�A�r����'����B��s�¥��/�Z��p�k׼49�B�I�j�BppACEK�ؽIWG�Q-�B�	S�u���� ����J=x[�C�I�\S,	�MV5^�ԫAJO�&_*C�1&/��3!���P0�D��M�5M�Ox���O������逑
_S%���4��*v!�5� 	�Ŏ��P�G#r!�dŜ��u��`��a�zع5���dS!�D�6>�*a��B��k��4!bk�!�QM2j�!��1���6d_�4c!�ů=,�P�"�ͻ )n8�҂�g�!򤛁~$���	H:`
eRp�O�����.j�]A&�.�\e*q(���!�ϡYR�Z�M�Kx>�꤇�T�!��S�hWZD���|L(H٣� �I�!�C�_|�7��F���Ŏ �!����"�^�:# �4��B�;�!�� ��a�Kػc!xɄÑ�=,�c"O����ѹ�z���V�2@�"O��h%�+MlI�@W�G��<Ҵ"O�T�!�Z�m��q�oQ�$����"O0l���N^x��S_�	��"O=�U'��'" XC��Ñ&�h���"O*�	F62�m#q�$ ��	y "O��5�\0a����Jش�&%Bf"O���$�a�� ��1s�����"OJq�S�6+>��u.�S����"OD�K��	�Ș*�㇭u�F�h�"O��BA��5��}�-R�0s�h07"O���KW9�18�!��C�e0�"O� s�FO�N)	r@�?s���*"O�p+����
�8*w�R3�L�
"O�Xp'IG����C(@���"O��u�#�b���Қ�f�=D����K60'��Y��te���:D�P�kX�D�H�f�ͭH�Bd:��2D���3��
pNF�����6� ��Ҫ>D��{h�<R��;qd�|s��Z� D�̱tc�+PT�%� �6�@�j>D��S��Cǆ��`hK�Y����9D��3��^"�u��I�-�蹑 �6D����m�}��E�E͹�ޙ��3D��*���<<��|����bV��#L7D���d* �yp��6䎐��K&h D���à�$ώѱ2��CbQ˳�2D�4���Ɇu���G�Xْ�M5D�� LK�Pp�dB��1tC.�t�3D�Ĉ7�3N~^-�I��#W�2��0D�1�K�3������<�,{��+D��:ōŖ=�~������F���e*D����kԟa�6Q℩�3@�����'D� ر��/��́�Ѥt�jy)�B%D��d/�5bX��Ui[�3	t�Ҍ.D��*C)�6P��(�)>���,D�<����paƉ�e�� u���P�8D�X���ŎD��8�F�2H��A���5D�@�0�޾[v��2/GN�����4D��S��Ѐ��� �2V]�Dʁ7D����Q9xb��u���t@j`4D��b�Ȟ^��aa����+s:Țf�1D�L��B
�ZB���hF�tܺb�%D������/�8uĕ<F�:�hw�%D� ;�I�3_g��j�����q �#D�@yGF��6P@rɘ禱"r� D��J%F(*�E1��m��U��<D�D!�G=Y��\) ɚ�*͚��s�;D�H�u*	#b����R��(�����E:D�4������TH�99�t��"8D�� ǃ�j,:�p#ˁ=�����8D���(�h����p'ER>NuJO6D�@{�ԅ����'�+��8�s�6D��w�W7L���K�++��,���/D���ď�8@���2��$5���1D�p�'�ʰs��py�)	kڝJ�l<D��cb�!<T��"S�rxn\���9D� �RmV�!�� z�f�/1�,��#l9D����߯g�,�A�-K$L�,<0$8D���-H�l��X�?�����M5D�\2�Œ�E��i�(�����0D��J�OMj���:�I� 1��E�` 1D����͉<S�Tp����E�)�e)-D�� �)#U��!5GÔ:�(�Q"O�L1�J�O���@ڐg����"O�0��2LLX��̈́tz:�a"O������a�l����hF8��"O΍�Wg��-҅q���z�ɓ�"O�Hō99�B��Ă�WP�}��"O�#�.�04 ȉp@M�1.=�!"O�8���O�`�:��l�++5r4	�"O����[-xBp$c��B�	"��w"O�0@I��=�~A&�/C�j6"O��Yv(A�H(�i����J�3D"Of��a��B���U��)x�T���"O��x�'����%�#: �'"O�0�fiI3>�^U�W؊6�T�"Oh�s��L,~�DI�D�/sؒ ��"O�Ѥ�
�6�օxS�,�b�;�"Op����@=0���#��t�:"O�mXǆRK8���C�R�8蚑"OU��b�7~���9���� a�"O�9'�T?j^�����;{J䊧"O�H�7J��%����ل)1v0+q"O�C7N��}�@���K�0�!
�"Oؘ�'i�2�٤��1+@���"O�hD) k��p�$B��ɂs"O
P��EޮňA� C�"�y��"O�9aTCH�wg��p��_�y�r��"Oj�����49�
�'��6�B��"O���0Ḷi�>9��Ǧ1�֌Je"ORir�J;P��x��I�>�-ӑ"O��AIW8PH����X�_6� �"O��C1��\�H(+d$S�E��I��"O�1�6�̝~�$Ȱ��B��Q��"O��ꦁL����$ɚ?��0)"O����C��z��PK)ߢds88"O��KSDV')(b���g����lz�'w���"��D�C�
Hvn�	�'��X
TM��.�su�B
R�! 
�'� ��s�Lt���e���&���'�"�!��8�)���-bmи+�'���$��p��z��֎D|��'m�My��EUKH��;h8X��'�f	 n��n���
���3#�1�'4JP�dIA�$�r�AN/$���0�'�~!�Va��G��<�p@ )F�q��'*9�P��ph|��qΈA��U9�'�܉PD!�	r`�"�Iв8bR���'��C���R�<��G��5ز9y�'��aW�[ 际��2\ �M3�':`q�P� ��ړFއX\	
�'�x`%J���ȃb2�I	�'���D���4� -�2�6x숍[�'c��22l̫$Lt,;q��i��
	�'�`=0��P�j����Q�a��i��'^�QY��^T�6���� ��'!^�
j�K���&�:�'�`��0ǒ�*I�k���{α��B#��`��\<ìi[B���j׌�ȓ^�$�>p*������P��c����*�w�����_�{V�p�ȓ]m,��C��P<�����Z�Ra�ȓp��+�$L,IUi��  ]b��ȓ*���[��R%S ���F�p��>x\P���>��IQa(XB��ȓ$�X�E(8�P�G �$h
)��S�? N�{cA��vľl�!�+`��j�"O���C�Ӏ-ɴ��S#��bx��'"O 5��(�,�J����V#�xʀ"O@�h����r�T5P�@#�0,m4D�p�.�r�^�QjN/��(A�N*D�8��H�� K�h�u
��r��(D�;rfҋD�t�#�
�v�>ݰ0&D���SF?<U�4�Qh*c�6E���'D�Ș�E�0WF������d�6���� D�4Q6G��W�@[G��F�AE�?D����ͫz@v���H7k��^�!�$K+�$�@�B^	G�Xr��W�!�$���p�A��ˁ�$8:�-k�!��AX���*��\*JD�ȳ�#��!���6'H 
D�;�� �ԧ�-!���;_z�0p`�@)j�]�bG��:�!�Ă%l��QbU$,˦��%�!��&
n`@����gK2MSR+�P|!���#t�G,B�r� ��,fZ!�d��]ɠ�K��s�p�� C��!W!�C�ը�K�L
P)�02cn!��J������;5�hW��wg!�݄ ���įG�%���o��MJ!��V;b錠��*҄C�����2{�!�$�5�4R�L��9~2��rM��0�!�$Y&]�b���LiG���%�׏#V!��Q���(ƅK�*��rTk�/_$!������K]�'�A��� �Z!��N�����4�ǈ}��dxe��)�!�DH.Y�~(�G	өa�f�)pȭW�!�d7?�x��(��C���V@?�!�$C��6��$�>�\ab`�mb!��8<.Viz��_m�\K��P��!�d^�F��ҧM�r���жJ�!�$ſW�Pt���X�6� '�\'|�!�ē+p�0|����V��:� ڟC!��63�}p�R�(� ;��Ɨoh!��Nm����G5E���)��FK!�D�=0e���H� Ϯ	[��~_!�dY� Yn��V���6Μ�P���|E!�I0�x����� @P�B�m!�$��E=z��M�LӘPA��g�!��L:
TR�Ȅk��M�1��|�!�	�P�|`Q��?���P�)�%�!��]gN�a���.y^�y1fӲ)�!���m�@�����Қt���ٚ�!���6$��$�R"7pV		�P*.I!��6L��M��?	��� �8}W!�Đ�K7�#��B�'���SԌ�%�!���[켈ʔ���>�z]�G�� �!���S�� ㇉\ڬ\J���0�!�	DX6��4��8g�~0��I��t�!�d��������B�6�h'/VUt!�D�D��%��U���#�C87!�F�G�6@��Iy��d�� L�:!��+"h�kCB�z
Eq&�̋BW!��gb��9L<n"M�# .w!���0U <�:��%d����]!�г!��9��W9ul���C�ټc�!򄇨��@�%J Px�so��8!���K*Z4zF!A�S%B���# �!�}�L��Z:n�@��N�Jo!�)-��s�-�a6�k��ҥe!�F�f�ZH��].W�� �o�9�!�� &}��J�/g�l-C��P$⠁�"O2��� ���X�� ?X¨��2"Ov��m�6:�a�FͳS�r"OFG��("/���4�^����&"O4)rC��30���G#K�6��`"O ,����RBċ�\�z�4ɉ5"O�DS�/�.4>�`XP._��`�b"O8U��a�&��$(r/��8��`#�"O�(rQ9?��A��>wk^ٚq"O,@E�4�����G'aZ)��"OD���L'��3�HL�a �"O�Բ�f��[r��Sd�`2��{�"O�%R�@@^x<�DH1u ��٠"O��#����xƐ�6~Q��"O�hw��}&����TS����"O"h�w"X2�m� 
r�d��"Ob1�G,�4� ��<��M��"O��@G�U;B��m���o�l�XP"OЭ�Tj��?�`C��N�l�Pj"O�(��F��)`*F'��-)"O�������� +�N��-���s�"O��qfT�4{�� ̒�&��e0�"O����(L�-CS�U�9{D�#�"O*�R�#�;/X��IN�mrY�"O��Xe�^�=v��1��+h<�!C"O2ܠ�$�/]��Z���6Zn���"O�|�GÑ �nyS4A��eet}�"Oк��8%�p ��ə�G� I�"O| �Ȃ�+�ҔٔJ#'v��"O6p���̱>�VU*�
1N�*��`"O�� �̃_�"�y�Iƻ�&M��"OT����6 ��dR�A�k���Q"O�`�*�&|�Qx���a��x u"O(�c&�J
�!����/*�R�"Ob�H��G�+�l<[$��x���U"Oܼ�s�βb�֙r�lY�ajɻ�"Or5���0 ��l���6ZY+�PT�<A��̹0$����bdiQ��L�<y� 	 -`�qG�K<���nG�<���0<����eHV�A�t��"�C�<�S%��,��+���6��҇/�S�<Q���y"�)��U�1 Ii�/g�<I���8���K4k��ީ[TJ�_�<)F=�d,�c$U9����^�<aCL�Lg��!�	�zĠ�ƭP�<������ �Fl�!~i�<���J�<�3d��'��Y�pD�Ds^����l�<7&�/,.eO �7������~�<9`��2�^�b��T g�I�U(�u�<��	'qy����]N�7i�q�<�ֆ=XOR1��%�5�L�r!� v�<���`(<@%�.\D�9�%M�u�<Y��>T�h�PV�	T� J�Xs�<	�	�#�8�N�$��Z�<	�� `���^+Sd$�Qt�	�<�v��ٌ<�ɂ���E��S�'b@q�S�M?.*��Y"e�l�-��'vH���Ռ2�� #5
C�ZJ�<��'�B]�¸P���SB	}��)	�'���k�C�������!�{6 ѹ�'���)��۴Τ!Rc˴b���8�'�B�C/f� c�-Π�[	�'����D�Z�,i2���+n����'����s/B�\>�!���(�*�H�r�)�� �@AÉ\#=>���p����d �"OR<Qs��6�te0
5L�(;s"O�QXňM�v2����T7@��bf"Op2�L������
F/T���k""O0,�2��To4T���U�{�H� �"O��q@*�?cS|��j?$�H6�#D��r�h׭J.ڠoԐ*�ƭ�p� ��^����^�Rň��z�Z��tM�
��C�	�1�*��@l@�fe�G���.B�I4wB�5F��ip�@<+�B�	�����/I�P���	^�@�
B�I�,�,�Ɗ_�k j5Y�kW�l�C�I�hf�Y@�Ȗ�F}"��:�C�	2~�܉�J�Z�&qRG��2PB�B䉗��� !�7y��(��A�B�	�T��x���S��R�VB�<� @�i�=�J�Ơ��$B�ɍJ�~L�b�˺�8 �~B�ɣW>~����4]�>dKӡ�p:�C�	p`H�a��&��K��6v�B�I\��`���
-��K�A9tr~B��3�B�k���EC��(����c�"B䉫7Ⴂ�X�@�<�r�iX�7�DC�ɤb ��qr�[4dstd����~F�B�	 b>V�SДv�K����@ZB�	�=1���>K�!��3}�B�I��-{���&E���-�(�HB�I!x{ iy�+u��D�S�Ů�:B�ɶy�8�!�K�����M!�B�Ɉ�us��N����CȲ��C�	�j�J��29Q|M�Z��C�I�[��"�@�+�h�����p�B�	?�� P2�K�踗)���RC��5�B�!�Jѥ���p7�I٬Ɇ�>�3v�H�Zw�Н?N�&���	{���	Ⴧ�F�����e��(�@1D��q�e��'���@��W��m0v�0D����2?�t�ѤP&�N5��4D��j�O�A����є\�R#�?D�$R�N4 Zy���p�BXDn?D��c1'Y3'�l�z���8~�&�"?D��CCJ�l۔X�w��X��i+�C�O,�=E����+n�3J�N�-�V.F��!�d� 1�E*D�&�(���T�!�Dʗw|y�'�Yi4�e��!w!��w�ڱ�L�	�@A��' :!��R8v����	�<��-;Q& "!���,��b+��c�&@���'�!�D�yA����^Zh����M;ў���I av�ɑ��H!�$�G�pC�	�����d)V� �$�R��ɕ��C�	4��鲪��Iqz��:�zC�?Q���穒�V��dO͓�jC�I6_�:xj�&P=��$�a�)ҔC�		&��ZsT
c��eĒ#,�8C�	+��P���ĭY�r=g�K�I�B䉶G"�����z�2H%�^2i�B䉉W�����B�hԝ�qj��a��C�ɮ^k��9���US�q!uǅ�C�I"��HV�-W�]���ĵE�|C�
=�<=�T�9rrPB�¾8lJC�ɏ.�rMh��H$%��3�怱3$@C�3�,��VH��M�l$�EJ* �4C�ɺo0��`�Q=~wZ4��΋'��B�)� ��-��^�k�]!0���"OJЋ��Z�h�r��P)�� ލ@"O�	Ǌ�G�d:b������"OJ P��w���ؒ�
�xȖ�X!"O�x#���;2I��"fD)v"O*蹢��p��L����|��S!"Ox�(&!Η�̤�th�=ٲ���"OL����5i�*�D�(o�	�0"O�K�		#�dY�� �_���B"On,���_�|��+�AG6	^�\�t"O�ͪ�F�n��DH����@��;�"O�` ���GҒ��A��1�$�Z�"O�`;d')_4$q�Z�C��(�"O�ұL��x�B(�o 7i�$�"O�,��"�:Q��A��n�f�ȇ"O�]�ŋ#I��E�V7OȌـ"Oh��A'�(�T`D!6 Z�P2"Ob�f��/[�6}���_
Ja��"O��9�a�
B�f�j'��u��T3"OR-���Y qTHr��ς�L	sR"Ol`!����~�
"I�\]>��@"OLHq ��KL�6��zL�4Â"O�1І�:I� ��"苊D1� �A"O���%�����Ef�7+,���"O��zTkۍ*"D�JvEB�
���"OtԊ�AȬI�:e�QBV�y�6,rr"OL��Տ��!��CU��68�p���"O�a��:E	\%h-�)ky�Y�"O
�������Y����?f�5 �"Ox;�C�F2h��OIR`	1"O�d��L��8X�Mbw��X:���%"O�	xu�Q�	D��2�ܺR�$��v"Oh�9 ��,CHlC���oϨ���"O�\AUk�!@�d=s�b�@� tʷ"O��{k�A �[thɵ$����E"O`���
�A���&9�n��"O"��%��
ń�(,
A��"O�xj�%\�{�����@F�|�t�"O��q�b��9�М�� ��%d��3r"O:�2rk��s2p����-R���b"O�H��k��xZ4q �o��3U� ��"OԘ�G�WH	,9�c�2��ju"Oj���@��5��� #�<m����"O�I�w�Nqy��	�n>ha��"Or\�,/�B���,D#(/f�[w"O�����X��U�Sj̇V<H��"O�p�G��z�؅�ai��Y���@"Ob8;ׂ�);^��e��#����"O�!�o��
j"� ���H��9�'"O�����2rw���B�
���@B"OB4h�e�|'��k$S�Xѐ��"O�8Za �3?�X�qa'̢c��xxD"O��� ��`�Di�&��PU2�yR"OJ2d@ߧ=��`(�_��Ux@"O�h��D� ��:T�H���=�' 1y���}�zM����B�\�'�2A�MȳI��	9�n�e�$U�'�z�X����ZIs5/� `|v���'��H���S�9�_�^M���'�@�G��D)h@.X�UW�J�'���6��+sG+H����'QB��Ï6z��A�H���P��'���ّ�s����2E��Z�'.�`!%̨uҮ����8GZmC��� |�!w��/f ��Sp͂ d ZF"OR�Ɇŗ�,��գ`Ꟁ7�f��"OX�AG��q�<���"2��DA�"O�)�C/I����aM$r��c�"ONTI&B&<��17/E�&��x&"O�d���8��UsDm^�a�"O0��@�6�f�JgJ<5���Bc"Ofd�n1'��\��	���X	*�"O��	A�Vԡ�4(d���"Oz�rT�_�'P�( �H�Kb�@r�"O*1(���t5D��gV+���"O2ȨT坸M�С8�*w���"�"O���Э;?$������y���D"O����69�"P�V} �G"O4{�U2{ΐoJQ�q�"O����<a�~��ût�U�7"O("C�Z�z� Q� Җ��у"Oʐȷ��4��`��n� �v1�"Ol�F�V�\Ch����\��F"O��u!�'S�5��ѵ3�*Ј$"O.�Pu���H�Y����/V���3"OJ��E�]����j
�v�X"O� ��/���S&ǹ&@�ʣ"O,9Ҁ�7?�`S��ҾK
��3�"OJ�x6Z5 ���閜	n���"O�$zd�@�� F��F�`�a�"O
P��I��8���X"�4g"O�t)�Ι�6�>р�F�/�R%i"O2}��5�~ث3CC�x�\�"O��s֍^+J�NI�F��9�|d�1"O.ui����ij��q���<�r�I""O2%I��$? ��X�F�b��tX�"O���Y9u2�K9���s�"OlE��/�9h�m �(O/�<@�D"O��[�
��@�tiV�z�E+V"OM14`�$/�(x�gS�&��I@4"O��"�ă,a9�)�%�9֡c""O>��	?|g��Jr��|�D#�"Oftz���T2�a�6��7�6!�"O�I1��3t$�RϱG�X@��"OR	�c&ɵ67b̡%��>�����"O�}��Ô�k����� Dyf"OD�����"*|�����!�.�"OX8��N�M�&�e��U&N���"O�PBh
m�D  Ww���"O���,�B'��hS .S=��"O����6>�EI׎�;d�f��"O^�"bЦ.��hF�ӅA���e"OH�"&��L�W��:>0����y��%E-��3�C+P�j0Ǜ�y���~��a�Հ%���	�Շ�y���Q���'��jdm�2�F��ya_h��a�Dβ�,���(��y��9n�`�$$[�w*����=�y���@�RRT�
�����@���y�o¶C���4P�F��P
H�zU"O��%�ޡ~�����V���a"O�j�F��+�T���Q
H`*R�"Opy�iF�E������_
$��`"O�Њǥ���F�)D�(g�`�[7"O�"��ԡ{��<��L'k�6��"O���ׯZ-z"�x��G���.�3"O¸�k� p� W	u�T�9#��c�<	�"
p���hؠ{�^ܒ"��]�<� �Qt �	�̤��G�6`ΐT�"OFi㣥՜v����-���"Ovi��
��b�T�8m�,1�"O�,��4S��*��8���i"O���2F��p-�BU�|�juQ"Oh�b�&�0+π(i'lĹ:R"�1"O��j��f+A��v�p�"O�Ljשا�R��iѵC��`+"O,h�1��-n\d�c��?q"Bl[�"Of���A 7?`�zb̀28��c�"O�9�d4dUMڱ =(��E"O�{'��C�$8`e
2�l�4"O�-�p���D����E:!�,�A"O2��F��U�
Ͻ9�zYIV"O~��JPK��I�"�����{�"O�Q ��QE(z��Ԯ:q~��"O�!K򤌀9�4@�rb�5.X�{�"O�eA�R&1]I�FaC�P��s1"O2��6CQ�(^*a�3�ً&2��"O,�[�)\�J�v��1�����H�"OV0��.�/!�AZ
���z�hE"Oj���+[�E���fɏ��8G"OQ9��,8�ha([$pP! "O<�+��X�6����Ԧ����d"O� �$��3��	A�@7W���f"OL�8�N�
-�l�Hu�S-	�tM�b"O`�"K�s| �s�F[�i�v��"O��8c�X6vZ�A�W��x~T��"O�D@��˶X9��@v��0Ts�ц"O�m��'��
��t�JKiΛ �#D� �e%F6�l��W�.gp��T#"D�H��*Ѥo��EB�. ��rA?D�t۴��a�ɫ��C�Ss�u<D�|���ܟj{�t�Lr��!��;D�$AS ՠa5���/��l��Pk0#:D�̊Vh�>95���E	��[����A8D�@�s��=�PأF��{gN�)�o7D��0UJ���)B���-CG�9D�8ڣ�ļ`�68�['R\�I���8D�\ìر=�Х9��7.6�qS��:D��'K4�Ҽ�Q��W����*OZ-��jP�_��@s!�:���v"O�I��Ο2�!��?-���"Od�����G���rweϳ=z�#"O�-��)���VY�D��w�ޡ��"O�Qs���~d%�����.�cV"OPI�#F�5"��=	 ĕ<j�i�*O���զ�2�paqA X�\���'�Q����9t4A���Q~&���'
���.U$9��q"�t֩y�Oz��䙙 ����A%�Ur#M�H5a~b]�\�B R( 0�hB흪s�5Y�a&D�4�$�ٵ>�b�K��LxA��	$D�`�7�Һ�Y� !_0Du*aO#D�t 6��(�|��I�� >�p#"�O�˓���r��1^�f-X��36C>L��"�.L{S���#ή,0bI�5Uդ(�ȓLu�L�tF��^��h�I��r�ȓq^.1����P��3�(H�ȓO�'�X�ص��/Y�h ����I\}B�D�>zA���R�K�;�����<�!�Ė�X���'A[�w�\�Õ����h����
$�_"��$��R;?�>""On�y���3VC�A���h}�5¡���﨟� �Y�pc� $�$�ؒ'�0�{�"O������?���7����i�F�O~Ez���K�k�������f?.8č��&r�y���c��1B�2w�x��#hY47Y$�=	�2��0�6���#hjy��(��I=��O��=�G �]�ŢT�{:�z�OP�<�3���	9py� eOXj1FF�G�<q��P*,�^���O;lc� x��C(<�ڴK�   ag��N�|9C���5����;�<��dD;Mp#�g�"Q��ȓ4���⬝;&5�y9Pk�3i,��=Qۓ;v�@qt�+z���(CIΘm&ȕ�OZ�<����F�[p	{��N�Y�P�P�ôV�!��	�lj,�qV�J�h1�Q��>e�!�D�X�B\a� K:\�ı��R�W�!�$�r�P���4�jY���
� �!��X�f���iX�l����.Ϭx!���6d� �t�=��( �͟^^!���42X�"F�����+��ۚS!����T/,WfС#i	M4LS�'����$GJ@ƑX�%޸*�4���Eӯ& a|"�?�D�N溜�e��STʙ����8)yax��5'�tB���$~�\s��H2'��B�	��
T
u&U?Ve,�8��F�G,���hO>��d��'~�I���ƚ ,�Rr$9D���� H�{3VM9R(�Q��6�	`�����A�!5+́X�$Q/y-��3�I�G�x"F��.��)1��i�e�l]��LB�I�~���l\7@i�u/��3�D�ƓBzN�!���?A���AP(	�x��<�>�ד"��ci��+-j5��M��CH~��ȓ3D3�aݢ��A�	(���h��0}���iu�a��?g ��#��/U�N��<����T?m�ҕ�S��K�r��3�
E��O���	ϓO��)��R�)d��d/��KJ�%���'�qOV;%JJ3�����A^4��"O�Q{�&�`���䯋%n�`4�&"O�-+ʝ*tW��A/�q�(t{t"OB�����+��H��@Cg�����|�)�;"�`�wjuf$�b�]�bM�C�I4��� q�Ϡc��ЈUC 4�O���$�G�,��G�>��xH����_��~��W�<iSiúd��Ȓ)ӼV�y��GN]�<Iԋ��$X��[�e�m�# ���'��$^	�(O��!H�צ!�Q�P�<N�T{�	��0=A��I6վ��E��b@@�P@��X���=�S�O���q���'�ȫ���&h�lx���'\�����#<l�r%݋>�<���'0,H��"I+�^�����*�Њ�/�S����G��`�ab�xl�%�˔<�y��>|z&����!}�4����>�y�I��� $��zA>d�q���yR��#<|V��3�O���E�P�N�y��-i���ʦ�%r����Z��y+�/D�L���ow��r�Ƌ�y���.0��:3�Νu�ĺBǞ�hO8�<٬�̈ ��M(B�ma�m�>8�6\0c"O�+a�V-0��� �Mΐ��9��'Pў"~2a��DЄx'�e/� K3HA���?I�'�kP��S뎱�@+H�.ݖ���'
0��M�|�Ѝ�GƵ~]p�'2��D�֐�{g ���r�'jZBu���G��b�rɂU�5D���!O�<�&`'JpgA�s/D�� �,"�)@�^'��!y՛��	z���Iųy�|P��)�/,.���f^�#l!���=x ��Ch�#@"҄Pk|!��7x�nUQ4c��1'rH���/c��Syb�|ʟ��	�,x�J\1	�<y���6rTC�I� 42-�0%�.)��C�%�RɄƓh���bv&�c#��)�h� �p���N?Q -�A�h����#q� ��B�[�<�W(�;뼥�P�ۡT�  �]�'ʛv��p�O��p3֥�f!�=C��(x$I��'����G&���4��+���*Ot��4ESd�d����}�'jQA���P�Гn����'��m���;(���#���<ȋ򤀒�0<�-��In�<AW�~�^��i�A�<�� ��zP�5c�!�BQ�P�KC}bP�$�V���'��Nƶ4����<��`peE0s�~��ȓ����CIܒL��S���4T���)O��Fz��i� T������V��n���̒8I!�d�1���"P��0[�,��U1O�������s�E�AP�{��T�qO���(��y��.0PC��kqF�����o�����"��4a�V�xa���X�US3'�Mk�'A:`;D��p��ŀĖ�TF�mk��~��^�V�ZIP7��(d����H�ybeJQҕ�l���	kv)�(��O��~��$�@��w�fG.y"VǇT�<��O�$�&F�!��
׺\����>�������Gi��bf�aZ��с�S��~��I1V�1O���Ih��������#!0|qtQ��&��㉛jr�$����Zd�2J��O�D�ʸ��O�R�X��6_Ϊ�Y��.�h=Q�'Ma2�W�UӰh(�L�0�J� G�A5�p>	L<�5BK&V�����ٖ�TmŚk�<قeP�A��,��mX�D� 3+�i�'�ўʧ��:5b�e���Z{
1Γ��?�a�Ӊ}��lzG��`מY`"����hO?����1���X)t>$`)b��-x�����2}rj�J� Dz�b��~~��`�S1,�B≞X�(���	���x���u���m�㞸���*i�i���L�U���"��<	r��b��IfE�J���)m�H�er����z�#Ƃ�8p��`��˴UG���"O�IA5b����;q �(��x3�Ixx��X�J�-.�d�C��=F6��Um(D�l�'�Z�5�Fi���/E�(�X�(D��a���$�r�K�y#�A#o;D��p§�/ :60
�/�6
z��c&D�`�v�kdfaNQ+~H���"1D� � ��'���W N7�H��F<D�Hj��W$`����˘
^�L�:«:D�x�%L�u	�C (�HR�/-D�$B�逫?h��T��->t�{À,D�x��B~�.��7�ѓ�(,�V�(D�l8��,����Ρ^�d����9D������7mZ!�AJ�Zlh�J+D���I1D�8D9���?`���%6D�d����&%����ů�	���P�H6D��c��Y:�����-p��#��2D�`�A$��zT��A��"o,�,9��0D�x3�O�4:4�I�A@C����+4D�x��jZF�I������!�?D���a˖�l3JE�3��V�<	�tb=D���5@�@��A.T�K5F!`Ƥ;D��#�I�? �BDK�ȯ)/EH�h'D�� �-{�2x���I�[dD�Z'"O.t��Mϖ ��SFC�Cn�<��*Of�pG$� //͸p)�-����':�4!#�6f<Z��D�'J���'�A���f�nX�����y�	�'��-�
��Tt�)���(O�Ȱ�	�'nX���  ��C`IػoՌ���'�z	�f��_��t��H��V���'��YҨtl���ǀ[d��Q
�'��Pɡ�]�j>$�
T/�#I�r��	�'�B�K��`Et���rP2
�'��9��Nǻ)cdz���	9�	@
�'�T�0�c߼C�@��r��	����'r��aw��;=��<�Q�/ԸH�
�'ﲨ@RK��Dez�:��A�~h,j
�'��yя̀lp�Bp�S#q�v�	�'�L�BlшoȞp)��=����' H|R�'���c�b�%B�\�����
(O���O^s�D�	S��,~�d�x�X�X&�I<��!���!�D́�I��"#�V����r\!��ˬbTpP@F\9��H����> �!�dɔ?��� W �>>�R�X��2G!�d��pS<A�Ī�s��� ��݊:>!�NI���d�υC���P%�Ū6�!�$��&,�7aX}h����)9�!�dxf���2�;�F��5�šA�!�d��3u2������pn���`�!��S�H�|t�C�W>��u�E2�!��vie�s��+��J�F7N!�dS�OEXy�$�>���1)�%w!��ڨ@P��̋$q�����IU� �!�D�I�!�F��R��N(Nl$��')V���K6�]�3�v��`�'<9��C�*0�Հ!Ϳl��q�	�'�"���%��#"�B�j�dh&i��'�*��/�V(�!pOHf�BhQ�'6Z���>&jP��+f���3�'~t	*R@W�+&``�V�[����'/~ ;��BR��kSᆣP���	�'�LP����RLD(H�v�	�'������'U�EQ��W6X�
�'Jޔ����=�� ��"I�A2��
�':�xQ���n��#<0 ��r�'��4�q�N>w��7�EyH*�x�'�j�ٖC�3il�����yM
H��'��Y1ć�t~�,�Q��s�\0��'J�1��mC�QR+<��a�'6Rx�t �
L�E�PeL�%��
�'JQZ��ĶdST̠vPV���
�'���H5�Ën�lA�7N�A
�' z<����,"�i���)�Z
�'
nY�MǠ8�4�F�� B�d�
�'͆��.��t��F�C�lCԼ�	�'���7M�<H��I�]�[<�+�'��њElM�N�J�(Å�2^�t5��'.��Ul�7���z�O�H�
 ��6�܅���5m��ibk&�θ��H�� 7�J�2���;�Y���l�ȓN4����#n�Es�*�Q��ȓ�v9�����s���"@k��l�8���p)FGU�d�hA���j���5J& �@�&i�0!I�E�ĺ�ȓ����Y/a�h��,O�����F6���*��2 �3D��)����S�? (8`J�
0�1�m��
�HV"O�0�#"�<��8aB�$h(�\b6"O\�� O�j���:�Z�L@�;�"O�hK7��CkN��F�n�`k��xrkH�W����I��1���Ǘ	���ܿ2+D���L
S���&��=��f앤o��-��kB'�B�	�]L�Q�����F`�B��-�">��+I�2�I��q�����C�J��!@�*i&�ĺ"O��b��K�l�heo҂ Рx`:O�}�䈗�S�*=HH�"~�e" @���a��Ґt�0�)w�Rf�<� �D�7��/�(!^laFǂ]~���6\Z���,E8�#��KV�T슳0�@<`Sc/�O��g�2~o�m9�L�
?^d
f��-@N���Px�jT5�!#���k�
��&���O^��"gip�#��'pD��a�02��U�7��	-P�	�ȓXĉ���`��3�,B<'N͓)I|iYfM3 �&ҧ���5���-XD�q���n�ZkT"O��C�C�q�й�%�A�|�����#���v� r�'?�i��~�~m	�Q�P���I�p�tx��_[T(���T�:���˗?��݅�{���f�6fav {0	�4D~��62ڲ5��\}&(x�����l"�틡�X���ʈ|\�|ە"O
�:�	D�<���kw�		�"�S�'@Pbbh�O"f�E��/�� hE�a�'��"H:�yb!ѽN!�`sNW;��q�C����TB 4�r����O�1D��O13���3�P��c��P�.��""O�H��X�us���r* Q���A�u���� A���9�BPeX�Dp�R�n����_7�h�'\O81ӗ����L��qa�J� !�deĔY����7�Fa���C.���ʇ�_�`4'��|��V;0� ��d��z���r���^�z���Z�lќ;y~�;���~N��>�C��9�N�@����ul{�ě6?/  �WjX|�3��-6����G.w|�m�fg����ZC/�v��J��ؗktָr��=�'W/��i߷Z��vG<}V���U đޢ)�%�^�a&�~B �<%-D ˖�Kw�ti����(J�V�{��2hS�8)Gi�$K(f��dmż%-ZӖ��v�nA��b��P�+KrP!�iP�[G����cKYx�T9��к_N���!�S�/#�"����&٤�(�ÜjZ�Y�oR�@��`R�[��>ع.O�>Bt�
^Ĕh��N�!	�Ԩ�J$����#���ʅ#C��̀���C��b>�cŎ��E U�!i�RM��R��:���%b"R	���ɟ��3�	,1��0keO���Q�%�.���Bc�0Q��D�1`Y�_����9��"Z�N��hp��愛�,=�d�p 3<:Ȉp �kI���	"��P�']�sBe����C3�x:Ҫ�$r�uQǀU�4!iD�#��T�;tW� 5�@y��^>�y�F�$Xla��W�|" 0��I%\fy�����z.�E���0�D \��<ų�#�r�Z���ӐOƱʑ/��8?,1�[��}�Ư�8{�Lt*T�g�(�a!YJ�If�"� ��k����*��AX8a�΂O�4G��X�1�,�HG<M�1LΣR�%��l���؝E���'
��6Z%2�A��W0zY6��@k)�}j�.��H�|�祃��`0F�#�|�C��W�(Ȁ����h���CA9�!�$�4+��aCX���l��A7.^]�J9>�J�L[� A��*���Gz�{~ �FV�37B��U�ø�p=�%l�R;~	�@n��M�U�v�NuK��D8R��Y��"Z�h��|7$�/��>iV��J����dȅ��Q�� y�N�ؤp& 2�E+)}�
 I�a^�yh^ �O┨����w����㒛"�R�[�'3��2�(�k'���ٝsM44�C�(��<�FBIN}��Y'Ă�l6�"|b�=����@˽7���$(݉�N��"O��bd@�T�B��`���������.C�Z�KD8	uT��-ߊ��i�h�'�.�:�IY�S���s�c�S
T�����^�R~�(���aD9�o�1w��<)ek��&D��X&��TX�|H5i�89>B�m�~��t�5ʓ@�TepE��;< j�H�}����]I�
[:�V��F�Js�Pd"O���HT�[�:eC%[{�a�uO �
�T�腪ҷC�2\��G_\��m�jm�,��`g�"5��GގP�"\�/#�yҌ����i�ҏ�~�ԣ��_��!�0އ+���A��C:�i�����w�zp��' �����\�3�h�l�:?W���� ��t�毒�6�|�����Hu��$F
��!?"�qOJ�@��3?� p�H���t�����T)\-�V�I"hrd�(��Q3v�>A`B�L,^�nQ���	`XJ�a
�%_�����'���:��Q2 �����ǽ����!ϝ�0S��^����|Vo��8��'�j�36�C�G��U��+���%	�'V
ș2���	v�3��20l���'��X���^�䌹1k4�I?	u��'%Z��!�&@�-�������#N�M��	�4B�X��˻8�4zЎ��a�u℩W�.Ţa��-!�ɴ-�Q>˓2.��reA
���S(W�lF{���k�XF���1]
 yP��������y�i�GJ!7X'cY ���*M�y"��*K�Om4��W"���yB�C9��皮F���k)�<�y�*շy��(�G��G������Y/�y���@�!X57���&/�yr��lI"]�r�^�֜blF��yҤD	s�pY"S�8(��WOE�y�$׉�H9���%'�������yB���~�|�D�!WW��ƙ1�yRO�tV�j@�AI�L_1�y�g�9�,`*�OX8\@+�%M��y��2?�5"Q��;$�x&���yB��;�0��D]�Z��8�Gݮ�y��(T0hl� dr��#4�Xr�!򄚀-3$�sFז'�̽JS�L���$�)���W�=���� �\��y��@R�i2�K=k�t��@)V������k�����b4�h�ǩD���S���5��O�\��5�jX�J�I
Ekq
��02��Pū��$�칔�tX����l�Ty��ӳn�%?�L�C@�,L�<(�=�?���S�<�@�S'�O�ku� <i\T)�$bLf�"� �W�qOT�Q��Y� �KV�*@i�/i~Z�a�N`�v�qJ���?�`O�4��)  ,7}���OE���+W$\"fx���C����x��ݼsDQ�4Z6�(M:�I�ZF��AG�fjbeA��ʶ^-��5�t c�O��R���E��HĒ����?)�r�g�B��p�9}ݤ��$(�8�� �>Q@%-���'S^I:����NQ�	��LGh��F���B���Ti�D� OMp���Ho"���P�oG\�Oq��x��$2�8qSAU�R�L��Q$�L�����#ͣM@瓧l�6�* K>�村 ��`���(C��1����W��(i`L��������O<�B%��[��6�)8x��CˍY�t�)�OHՉ`c�^b2�R�ΘZ��>����V�x�yP�Rz�d�s�2=�rdQ�֙&��\��x�Z.z}�EK"�7IVXb!%�Q�������<���'^��(U�ۭ}}�}+�ͶN��dN\HGB�
)֠��a��Q.���6��]�F���y@F�i�G�#
ru���{lL �M4D~�8(��W%t�� �g�&}���f=&@����´��A�+�'c����g�1�"��H����`FM,p\�'Z�&���I.#�lx� ��/eL����R��	�2ZƄ��OF�rMC�  @1u�@o	ڙzc�-�$<K!�O�pk�.�#!��?�Zd3�lA�LcD�I�G��_�<�������a4�O �J�*�`�Vp�$�΅9�`��M�T��49�EK���l�D�J�4O0P
F�B����@5(�Z����]�O+���nƗ�a{�)�2a�����OL�b��O9{A~@�ӁZ���x�"O$M�eA�Щ�̹C�L������1�A����W��ڴ;e��E�n#P�Q';�!��ͦ~l�@��*~���Eky�!��:B���u��s>��A��͐D�!�D�;��]+u��+J/�-�����~�!�D�����
���
�!�G�
�!���M�`x7�J��蜉O��!����t�D��!��]�Tқp�!��Ї�x�w-� �J�(���2el!�d�P8��`�������W�!�d�)�fL�6w��"r�H�P�!��m���X�a(S�"0���!�$�60��c�+�+>ԡ��Zb�!��f�<�B��O;�u�sjQ�L�!��L=�&PJ�ĝ!6ۀ�R�ŏJ�!�� F���A85�����'��"OHE���,=�<�9�Y+YJ2�"O����X=�"�S��F/�5"O4њT�*o�,	w�_7�Ċ"O��p떬u���H��F'�����"O�Ł�_�m�B��׬I��x7"OZ]��tq����߲�� *�"O�ۖ	�;��t�����=��J""O`|�P#B;j�X�9£\)�����"O��brNP�NPH�SG�ܖ׶�"O���ܨZ�r�8r��[$�"Ov�0�O�#\�25���%��� "O��B!�1h��#�O$-~��"O��5�$e����%�9$�`�"OEZd-�/c�2��^�;�V�H�"O�X�v" �A|�Tr�&[���@"O�h�`��4���`�B͛p���q"O���Ǉ8U���� ޫ1� �g"O�L�ĉ[�5x�*��E�DM\��"O�p��eя�U��:}( G"O�Bq��P�����D�qQ�H��"O�|���W
�e96#I�]���"OJ��aK�3vBx�Í�#C�l�"O
I�f(�5��хȜ�F����"O��д�� k��0ˁ��}����v"O$Hc�$�.k��@��Vp$��A"OD��S%[)i��-����v���h&"O<Y�q�[�*Yj�NN�x���"O:(�U��@LR��P삳YWj�T"O���6�7�����K�6�h��"Ol�*7� /��zVꁆO�VQ��"O\ԡ�m�}�6 ��'
�~t��"O"��6��-g���k	�'t|\�"O5!��P��H��ʘ�|2h�0"O0�g	�--�����6
hڽ)�"O���ˌ�'���#��H���Y�"OJM� ��Ȕ_�A�v4f�x�<�P��o�2��Ek�N/�)Pӡ�t�<��e���z�:���6NUڢam�<��ګs��H��$��g/����D�W�<1�B��fyj�eΝ�+)*�����y�<����n`[p�"clJ�� IRx�<q��`����X�KvLفVj�\�<���mw��t̓w�*}�q�S]�<Q��ƆF�uI�@.g�� E�g�<6�;(���p'(G��m���GU�<Q7eV�X=�VnW* ��!a�H�W�<a�BG�A�\(��G�+	�\=YE�JN�<�T���df�U��d�&u��%K�O�<�1-ϐ�Uq�j����b�B�<�T��r�蘛d�T�x��	��IB�<	�؞|N��D�]�`�r��A�~�<�"�h@ԉs��7n߂�sҭB~�<�4�O!,��%��f�%�Y�.]�ȓw�D��ej��B��x�@nƗ'�6���d�`��s��5X܃� P�<A��aƬ )�|x� h��N�S{��ȓ3��Ћ��[���d��D	�=t��ȓ2���k�>�%B��H#5����ȓ$��4��F��nyX�� �E�U�R!�ȓ&�
݀7'�.X����)	���ȓg�f��N*I ��	&cצo�8P�ȓ"�64�2"D�L��M� ����ȓ[��-�e���9m��Is���z����S�? d�ڰ�X%&o��86%��#�h��"OZ�败$A�):�$T9;��"O��EJ�*q�D��B�o-����"Ot��5����ܵ�BU�d��ip"OneA�+V�}u�@�P�&$t0P0�"O�����7�� ���[o|4��"OZ��F)�"�b���JE	PGh��"O����k�ȹ&��HK�e���xbI������	�Ux�\kf(ՒںB�#�??����ϱi\���8$=�@Y̑�3&�8BY梈��'��y���ʈH����r-O���9����m�M!q�����OxY1"f�
[����&*�|��'�f4��-��B���!�z���'� ��iE�ȤO?ED�&
k�؈5�I�-��9�5�1D�a�Y.	?��`��br�ڢ#)?ɑ���%,�̀�'OT���\�tKqm�ZJD-��'���b��8��@���^8
��(A�.��R��A)�T(<��
K�0�ĐDl��Ѐls�mHA�'[P}9҆���e�}��/\7��ҳ%Z'v�ĭq3�MK�<��·�#�����5#��,��L�<)R����7 ��ҧ��^H"dJt���1u�N#k�Ny��"O����(6���x�9�Z�1&���!�ۮ'uV��s�'V:	�7�ZJ� DKȈ��0�M�t�ޮ$�1�P*��=0>�H2I�b��B
�'H� @�-cMD`�)W�L@��$�t�lc��t��h>8��#��i�t\��`���yb�T����&��0�$TP���y�T2BA�,�`	�&hH�3�HD��yҁ�I�젳�%ش��Ι�ybG�,uV��6�G���2��ybD]il��&L��r#'�yR��(-��Ȃ�ӻ?䬑��&�yR��d��i.���bF�F�j(�'�10���ɧ(��8��0�*d��GLMz.l��IM��캀�)]�4B� `WH8DcH|�h���'�Ђő�$���OppR�΅Y~��x�&Ж~0�ȑP���l�4���$���b�`�cS�u��QZ/�!�#aʘ%�����LK�os����x��\��'X.�hi#M�A��1�O^\����=�&k/X��h����ė,oN��?�A��n�h����)\kt�Ҩ(�O�$B+�xf��1m_!;���Kѥ�>&|j����Y����C��Q��[��<E�N	&h����MU"^��ĉ2��O�Y"�J�Z1��酜]�ޙP�=9@�cq�^z�Z�?��`�:}K����'����T�4�z��L���|%A�'Ԫ(�b��U�O1�x1y���,M6��bÙ0�D����� ��f�B*3����Y#���C�b١(�n����Ӟ#��BT��2�eZ%>B�5{��}BF{�X.���O��]Y!�I%a�%��I��� ��~*�$
�%B�.q��ߕ`��ECpo��T���ԫ^��E1&h���|�B-O�>�������lrw"�7c(0a�*��2p��L�u%q#�"3�q��a6��R�u�:|JP�ƙ��I9�a�� Č��g�s�D�ȵ+�b�,�Y�d|Ե�'�8 S5�̫1�0���y�Ol�Ae"ѕr�8 ���K�k˚!*�%$R�U9�OT�:�#,�D)F��A(r�����@(�5��Z�� R����g�l��Ab/\G�2WJ &�C�IM־�+�fF ��B�=k��U��ʿbv�!�'�ԩi�ئe�
�,I��82r*UAx�$&`�"��$RZ�Ȃ�.f�����݋���k?D����4~*��1��>�@��<�䘄=�|zV*\/�ȟ�,a@��/+��e) �17ax��"O����Ky\\��&f��br�-Cʉ
��	�ׅ�h`�m)�35��3ʓ{�Z,C���b|�d� �HS���I%/��r5��d�����H����)�%q��}�d.��4����	8�OF�3���na���$I6�r��	,�J�� �o u��k˴'L2��O?�i�T�C:,��xu�T'�`z	�''$�����$�"��E�'�DE�u����aJ��B,C�ZTRb�T%\&?�� 0x��%w�X6M��a84�$"OR��4�
,L ��FM/�@�Ak��Nb���t 	m�0l8�"L����)$�V�bei���p��X/������D~x����I��%sij�F�Q���A���Q�'�B���ğ�r���ۀ ��E�N����Ԯ:�Z��w$ߌ����!A%4*C�X�D�6eJb�*�"O�u��M�,�qe�<�d���'���R���R��S��?�B�>9�|8�4�J�6�S���}�<�DD� ]@\��R�5d��<{�z?	�
�q��9���9LOdа੓u^��❲ ���9��' T��#Ɲ<5�bJ�ze�!����<b y�g-;D��Ȱ$�tLL�3���cM}+Ъ/�>(6$�!=�'`*!�SN�V���7�D#0�ެ����Z� =o�  ��a̲O`@}�"O�y�g�Ѡ}j���.RX���"O���� 	�X ����z'��I�"O.E�P��>���a�j�d��"O@�ECօV�"$�B����"O�0c�N�"*KԱ��!�h�x��"O*�c���`�y)��F�"Oh�h��� �r�a�!X&/?j���"O�M����!9����*�5H�jlQ�"O y r�SR¨��	� d�x�"O�����,� x�Q�� 
TiS"O,����&}
H�[3b�:d�	C�"O���Q��q� 1��/�+��I�!"O�<���b�h�H5h���y��"O�1���P�B̼���(�w�����"O���`k�s}
E��:i���	4"O��C��#7(ЙR`�.�g�� >6���#��Y�,��^<N��私0Vz�3�!D��A�ʧN��l�w�&8��SՆ&�h�D�L��>9�C��v9�ɘ5"R4h˦��C��T�4ڐ*�qC��O����嚪w/�*7"��*U�۩,]qOZ����Y����=�ָ1���K�T��n �	I�|�Rn�1\Q?aà�Q;�	�b�B8 }^$YI@6�q����px�H �
���[6�Bm�8�	ăd��  �>���1#�D�F���=��K7p��'"���X"��,����&3�	�%Xa�4FB�~�	U�c��iw��
��*�h�-�ZYi6AN�s`�鹰��'�"���5}���NK)q ](f(q��-H��ۡ¸'��a�� u_N��:-N�S5����
�Ӗ%����Ǉ'.��JQ&O'ΐ\9銨���I���O(��#��q��땍Q��C�?8:�1OZ���I�5"&����d����8b Ğ3��%# w�$��q��!V�A3ؿR0a}� �u(N��P�M���M� ��6]�0W��		����'b0]9�@
v"V���ˍ���e�pF�>I�$�C&���,9ZLE���h��0����Tݺ�I:O�(ʕ�,k�X�dJX"(��0�(��_�d��fK>@��=��
�1h��0�Oq��I�J�-K�����7�@�3���[�J*�)����y��<ϲ}�T��A��T�"�FoN>电h̂�i>L�8�>a������6^�����)�+��Q�j\#%��H�勝�{�V�IW�5�D[o�'$���r��`s��ϐ@���+��Z�HJ�|1��O�}���	w'�%0�� [����ؼ$��hhw� *���	�>6û�扬O�Hp��4�'F�fQ�i��f1=,]*i&lOؤ ��äI� ���ZN�@kQeځG�8���|�	�'Q�X�#���Y���>Y�v�;�2K^�}E�@E���c�H��`ۭ+���H�B��y��P�2��P&Z��E,�;�y�-_�i����s�,H��X��S��y��D1��Uk��{*0	u�D�y�/4�q���E�F0�����y�z���"+�qF�����;�yrf��O��Z!RanU�7/H��y�(7|��1rS��b�-���&�y��`E��'Ev�jq�'��?P~B�oP�`a�-M�a�M$C�)� (4����( ����u^�S"O���`�iLHQ�Eg����"ON�%�
ڒ�{SGO-b�Ց6"OΙ)P�8�Z䉔6h�����"OV�WjZ?'��!�2� "�ŏ��y�ŕ�\'��9�MЇ +��:"��#�yb��:ݠH����<���b]��y���4o�)2��<r5ƥc�J�$�yr�N%cqfi��H�=j���������y��<2Q4I;��8c�y�&ҹ�y�Ґ?jtB���;3���1��ؕ�y����7�#5��)Y� �ےɂ�y��F=E�0	U�8i5/Ӝ�y��Ֆ@���"�FѪLM�A#cC	�y���	!@�ąC��m���ߋ�yBE�'H���T!Y#��!R%j
��y"�� }x��{1)ǎV��b(�yR�A�7�W��Lia���yb�}Z�T@V���Y��(�&��yB�Q o��Ћ2B��J�J�2*�y�&�!b"�k�bńtk��#�W��y�c�O0���O\�a��-��f,�yBO��rJ8�q��"4�Q��,�y2c��K���PC,%k�M�5e���y��PV�ajRa�
d�ꥠ��yRj)R���6�l�=��	�"�OTq[�JV$�ڙRsmף@4$� �lU7U��q����-!�$ ���oPplR5[�laA�e]�|��Cs�S�O�D�Z5�ە;��X�O��gP���U2�Y�3��n���)O?��7+���m��ʙ	A�!3�E~�`�a��'���䧘O��E��T8�r�X�L-�)��b�!+��#l�ӟ���ق�~ҥ���0|b�N	�"tx��֬|)��AC������
"�dm���S�N��FK&!z^�cdCA�
&*A��!���@NP���:v%���x\<���MM�O�p��)��̅ᓨk��C�a�8��E�g��"�6Od̈�*ޱAQ���|��|�e鱄׼%��}2�#��?�7nJ�OQ?��r�F�4�� ⃃�(��͊`�E�.6h⟼�ᓌd�DacO�/(�29`�����c���3K1���f�-�{�I��ֽ�숞`�'&�s�E��=�4�D�t���`����M�,gB�k�e�:���W�m�B`1�{���ÄwϬe�L�$8%�+e��
>�����5,����=E�$2���.X�q��j���HO���ᓍ� Ц��"=�L�	&iEOmd� ���)���'qR�AR��3s�a��$�.;��'g�"=�~zAJ��|�湒�!HHz�G&�|؟`��)'��Rp!Y� ��Q�ⅆAs(��>q�����!;,/5HW�I�]��lУ��?��bt�OQ?����/jB9t��b����o��<�B��>�'i��0VJ�%�8=�CΈ?r��=��}򯜿a�����O,r2aX$e�́��xx�cy��'� 9�/�dd?��Y
������Y�)��'�P�p�����.����O|0�	E-G�
=a�����|�At�T%7�(sVd���?YPD�J��3"����?��N}ЕH�i7ؘ+rk	%'�̅�S"O�Pf
��Q����'�1I�h{t"Od�x�S6:P*�CP
ю
<��`$"O�*�� %3�%jӨ�~W��W"O��3����v����G؞BH��v"OP#攥?�洘#Aة?�Z�"O*i22Ń�mL�8�Q@ZC,�"Or4��'�?Κe`��Y��L0P"OP\�V��s��H��c
	Ӏ�jE"O����.V�p�!Z1Pż|��"O<�*E+J >w�u���͏n�v���"Oܰar��,^E����2��UAf"Or�w��23�؂��0p���4"O� ����B�Z����ϑ ��:"O&� P)��{����W�%�Z�"Ob�C"�³!������:}(�I�"O���[*j�q1`��Iv
v"O�ɶ-��Ɲ1��&�H�ѧ"OVA!��(����dm �;���a"O~0藫I��8,)W#X9Z����"O�t�w@�7OW�	#)��S����a"OzD�q͙�E���L+,j�9�"O��(g��� �a�U(%\�4[d"O ���LK�p>Ri�ň<#gt���"O�ڴդx��h�G�4>���"O�M�0��.>�����i:��!"O��Ab�1zy�`C�4PS�{F"O�m�٠roh�q1n�|;2л�"O(!�c��2sTdPP�,0(h�"OX�p �U- �~|�cI�@�u��"OX����^?{����H�^��"O��E��	|�
D%["~d�l��"Obar�$d�΀9ai6;d�a�s"OVEQ���
)���J�>[���"Of�C��C��~�B'������7"O�Ph�͋�1├J�O�]�޼˴"O�lp��Y�e���-C'A� �2�"O�dAw��B��gߠ~�0���"OH�S���L��}�$��uܐ-!��Gz�\0���GF�i�&_E!��=���F�# 2�H
V��y_!��6TL�:�"�u���"��m�!�D�?R�6ᣣ�!'�DbA*�.0�!�$�VHB�SF w�LtC��X�a�!�)n��L`T�$	��l����U_!���#
�h�I���+TM!�U�;Y�m�u��{���I���{8!��[)vS����^}C�[/7!�d�\���H�Nm$1'`I�mz!��օ �lI���<�� ���:mf!��8/�"�)@���#��r�";Y!�W����΋:�aѢ�Č7^!�$L8_JEQ�� �څ�����!�]}�D8Ï�	~����,��!�)$z�����
}�a�1���D�!��]<u�`[�K[���� CΑz�!�D��S��=�צ˶~�J�Z��<V�!��T��bG�p&9�FNޡ69!�d�S����T�D�F�d��<,!�@�\�T�࣎ �Z�C^�!��QDXQ�C�������J�`!��ꂠZ��R��ki�!��,(�V�D%�rE��Q�<�!�d�Aҁ�J9.����% �a!�DX�EM��3��r��!���_`!�ď3t< �91�JDtp�.���Py�lީ'Z���2$� L���'Ĵ�y�#�r�젡e±j�����Έ�y�Kd6��+s�C����8���>�yB�^�9���ku"P�fG�a�S/�y�DKAލ�ŀ�e\}#�
!�y򉛥L܄<(�(����i�@��;�y"��CqҔ
e��y�0�/�y�

�R�ka�0sT�X��!�y*�>_2����Ҿ4	�?�y�ߟ#V�3p�"��l����y���b�`��X8{X(Juf��y
� TM�Ca�XH�AMG�U��@:�"O�d��,{���];�`X�"ON@y�
���Ӵ�S,1ц�+&"O$@�P��@h��˒���Y�B"O(!���ĵz���8'��p�ܐ��"O�ɃT�V*�fK݅��ِU"O�Ď\1jh��%��~�*��s"Oje))X�1�r��VH��{VDQ�"O(0�)&���r��/Z�H��"OFyf�p/.��Ÿ[n�r"O.�+�aG�2^st���P[��b"O���"I2c��F�B�vE�"O��I�ɳL���!"Ƀ-ZqH�*t"O�ykB敾3�Z�ʕ���z��Y "O��r��4u��q��V�\t���"O��(3A�+kܼiL[|���"OdE�T.R�8��)A>5�A"O����`�0S1��:$Q����"O���i�.'R��d�΃fI����"O��S
1[�L\V�GJ&
IC�"O�e;phԆyx	y@͉�-j�"O``���J�cJ�-J�˚$Z�PH� "OH�Ѐʏ!EE3�6m4�h!"O,��V]�i��M�EΈ�_ҹ2w"OZ\�ƍ�7ֱQ#Unn�9#"O��@���gA�x�V��'YW,-;f"O0I�V���cPt���F-�\[�"O�	aT�ׂP���P��߯;2�i� "O�i�'���C��Ȳ�S:w#�aC"O쩀�"�Z?�P�4�4�QjP"O0��po��>�։�3&I/>��"O"53"�A>gi��_�|���"OZ��Q�U+}��rw��Y@���P"O��JBB�"��!���;RJ� "O�P�fe�+}�]���Z7	>��C�"O��jq�9w�"D(��ڰ	
J�$"O求a� {z����<ZZډR"O��{�HKJuA$��TIP-�F�<9`�$j��*��)`�
�q���<��Հ�t�X��F�
'�xyb(�w�<���ٙZ�� xRB]�$
��M�J�<1gͅ�)B�4آ�W%;e��B"@{�<QeF�������$o�q�-��<1Pb�;j�!U@-�<bl�U�<ytAN�a�T �i�K�<l�0��I�<�7�t�);�đ(�����C�<�Q*0v˾�PF�CS�FY�w�\B�<a��N.k�hА���\N�� ��T�<����#54�5D�:B�BN�<!����G��a3�
]�B ��!L�<�v+�9KȮ�+�e�+3�H)��C�<Yt	 �|��՛��@ H"<�c��|�<�׎9��}���xi��!EAQ�<��l�s �D�w��E��*Ef�<ه��]��r�Y�[+|�shJ�<�Aݠ}�����Y
7c<1˴��A�<�w��NR��C�~=��^V�<i�KH�8��$ʃ�6�`�12�z�<  U�`Ǻ-�A���a�5{�E�s�<)��'���3d]1&��`2��Ax�<A���h�f�ڤ,.y>�x�4B�h�<A�( fU+%o��>?"][�N�k�<��GS�>4����W���zpQ|�<�C�#<9h����al>��Fm�<� $زC��n�Hu��˫n���"OL�bW��4_`*uـD9wjB@"Ot��,�B�D��Ǡ�|��d�"O��ScႏwhJ�&�1AxtIR"O��Q�\9��8��$��fYzEؖ"O�p�f.U���A� w��#"O���A��7d�����U�U�4�
F"Ox8*ք��xa�ڠ�Ո}�����"O��01��$B��D��F��%h"���"O��B��D:J�^�����;f\���"O6e0��E�Mը�M­�""O���Bf�tn�|�D(N_� ���"OJ���[�I����A�-<����a"O�Qٰ���O�&�U�B>cZsQ"O�lPc��O���j��^�c�iP�"O$�	�D�K�P�#��(�Ƭ�"O���S��y���SbMO
s��� ""O�]���DF\[�k�*+��1�"O�Cd�N�=x� �/;�h�3@"Oƕ�a5d���^�*DT�g"O���H���-W�����S"O,���G-vQb� 1�y֢<�q"O�Uv�Vb�S��=4����B"OJ)D��(wVt����.1��<(%"O��͍�"��p㶏�w��u!"O���Rk�;,̀�4��),�j%��"O�U�P��KqZ=ʃK�$~�~���"Oҝ�K�4Xh�6��
8/��{"O�I �)T/ ��Ё�b?�|��"O8:�X�i�|���
$By�"O������u�2H��S�"Ox�'�I/8},01��	Nx{p"O���%f��#�b���B��Wv���6"Of`�7j%S����b�V=Z=x#"OP�	cbȭ��D�E�%d5�p�0"O`��A,ѸO\��wc�,
2t���"Ov\����.z��p�![�w9Rȡ%"O��C%.ܠF�l�afAL 9XӦ"O�U�U&\9] Ɛ�杕5A�"O8���Gk6���<P���w�Jl�<Q#G�����=�I��`�<�Ѐ�J�`�ͅW� Y�a�b�<��Ev���jJz�2��\�<��W�]T��@(�S�=b��U�<�I�Q�$ĹrÅ�STj��NN�<�@�3z�$�ih�t�cFA�<)��H	%���G3Ӟ��ЉM~�<a��>�R�QdE��Όx٦�I|�<�D��#i���B X��,my�l�L�<�5!?W+��C���9`���WE�<�D (�~X�&M�G)�}�&FG�<	#�ھ*w|� B|����b��y�/��4����.�dNӎ�y�4VO��x��,:$� Y��]��yBfN f �Җ����D17�ϗ�y"��6> P  ��   E  7  �  �  �+  7  �B  cM  �V  p`  �j  vw  Q  ��  �  k�  ��  �  6�  z�  ��  �  D�  ��  ��  B�  ��  ��  �  ��  ��  ��  @ �	 � � ;  s' �- �3 �8  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r��EQ�( �gVlɦ�M,H"�O��@Pg�9^��@9dr<8�q�"O�Q3c茟u4P�뒤���%��"O��$f�2����� �IY8�(��"�;�g�6��I؀)?D���嘈p�l����J)�4rŭ|���=E��4a^dX�(�7#!���O�iV��p���%����'HN�+���?�|��v��6��lp��~��˙}ּݙ7�I�<.��2���?�`;\O��'�LG$�4[����G '\�Lы�������I~���4��;���5M]��A��D�>���O��u�T�Ѓuk�a�V�ѸC�00�L<�N��E�����̲d��b9���3hY��~r�)ڧI��q�ȗR��z�	Usv�,�b$�j�����d�7JC:�H��B�{�L�I�&J8u!��L$���W�۠T������,!��/��H%,����P��/32d�xR�)ʓF<�<
���J �*��Z�(�5�ȓ,o�x#&�En�҃���h���
A�t 9j��b�F+� ���?��nma��[ a\�0d�N}��X���O��8�AAd�",⑊��~h)�'��	�2�"�J�l2R�z$��}�F$u��'��� P3Ġ��g�D '4��'�@��.��e�5�V� 5�h���)�S��e�l�$� 0�!f1 �b��'�y
� R�Sa-`liV���{a�P���Z�'~�>�I7Bf��S�I
�#{ -�6%�C䉇O`�7��)��(1���~��C�	� Ǿ�ƭX8����ƌuJ.B��>0�հ0�S�{�t��J]�HϰC䉍q3���`	]-��A"�֓B��C�	 �&9�u��UJ�#�4A(C�	�Hl0�n@
R���v�7��B�I.f��U�P����@{0F��,T�#>э�~�F�1i/d���=��ѡF �p8��$� 1��U �T9G��(فB+D�hP�I����rgR3��|*4+D��`e�h�Ŋd'�FS`��Q)�a���OW�`���(��d�$�`����yr&�8��Uh��G�Z���bB��y��U6BT~-��Ѣ`�d@	���*��x"L:yTn�����/5�p!4�P�A�LB�	�faNe"�B�[�<�+�.�$���>�/O��#U�7d���4j��*�2�"O��P�E�碙�5*�6:��#p�|R���F���J�N�t�ل�ơ!�6���;�y҃ύe�8�� $�#������2�?i�)�e��|)�@K<6��XaK<$�,�(
�'xr���N"l�U�/��f��0;I>!	�[�Y[bB�0��e\����!D��9D��%`���U.��\4�@�3D�L ��f��Q-�}H�ՂC�l�3�O �>�k��)C���=�tyZ��V��<�>���/K`8
��Y<m���ऩ�T�<�`�掭	�˜�I$1��EP�<�s+	�el&�(��N�d���`�O�V�<��C�x(0J��
��- �G�S�<��1 d,�H�J�Q���APS��(Odͦ�����gNy��xc I������"O(�9�k�:et���BHJ�Z�8�c�2�]%�"}*�w�$� � �>	����栤0C�\(<��Q,����FJ�90�哑A��O����'���D�ɶM=�}9�n��R��0X"^�%XJ���-�$�t�j�j���1m/Xm���E��j��G{���/@Dg�At�̲�6	˥H���O	mZ[�O����`ΰO������Y�80QK��"R�p�z��DF��(傐ef���	ΛFV�GP�����3tR��#�M��O����X�rܠ][���-_x� Y%�u0�ɤO��'�Ѐ� �'qW�0��n�:r�x�`(-6�$��Iw�=D�y���+3�DyT׏ ȀG~2�����H!!�fpc�@P!M�㞼E{J?Ij& Ӿf<�z! Z��J$�H]��yB�Dr��i��ҜHGvhs�Ѱ<��,1��D���s��V�,4�;���( �B䉐!�<�0d`�ZȜ�&E�{�O8�=�~�f�O��zዱ�͗/bZT"!�MЦe�1�\�&�W�2�H����yOP���	A~B)�o&Z$�&%H�X
\�����y��*Hm��Y�$�W����T���HO:�=�O��(V�>�"	��$B09�D�p�'_���i��5��qpQ�8R��4�hO?7҃c��@IM��w�N����%X!�����cé\�}֋�X}����Ez�reA�9��9P�,�]�!��\�B�x���7,B���'�a�Շ��BTӅ��Ikj�[@�x
�L�ȓI(`�FĔ�R���O	(�>Ɋ����@�3`�02ԡ��e(ô�އ�y
� ]aՍ�13�J��#倻`������F�|�u�ӵP-"����G(����b�<D��"��А�B���9�ĥz��n�^6�9�O����H{�j)�£��4���'�*�zO�|"��74@�fѴsG8\pԡ)D��@_���	���,�aU'�O�qȄ�3k�f�B����Y����ȓ5@y�7��*L� �&���PD|�J7�-��D�[�<l�C
�}`L؇�D�!��CR�y
8r�m��[�,̓h��������X��u",t(�
4F�.܇ȓk�:�BŨ�k?�����{�
4�'�ɼL�PH�?�O�9���/:���&Α'q�0!	���94�Ea/@�F գ�f��5!��)t ��Ȣ�Dg���ƃX�!�$�"K ��`�^��d�U�ĸU�!��	Ғ(	b��SKҸs�$
�,��;����Ob(�W�G':*0#G#2?HQ(d"O^����<A�t剗D�"hD6�3�^�	��'�r٨0�-F3ʠ1B���n��Ó���\�K����"1iI�<T)���JZC�X��k6����O+�ܨ�MÿR�2�G{R�.����N�u��qT"�,���#R4�ybC�O�� �+��j���ML���'p�{�پU~$�(��]��*�ó���x��'#X}���U�s͸�ǟ�3xP���'e�8�_��D@%�
s�|�!�CAX��Gy�o�2sK�A���v�@�$��y��f�r��ǣ����A����y�����FF��zʤ��C#U��y��	h=+u���%n�\�B�y"�Y�0��d�3,zr=�G7�y"�ُ¤���Յ���zu` �yB�%r	JÄ.��=#��p��y��r5ӕƍ2��ҷIϒ�yb�kHX�1S��>� P	����yB�Ef�~l�f쑗	=<53 ��y�(�\j�2d�Q�
�v}pC%��y��4���r�	-@�0�l]��yb�ä*}|Ő�C�t<����R�yBL������DH�d8 �JK<�y�!V�o�Hr��Ô"��3c�?�y2����xӀT�2��1`�9�y�ʘ46�fh^���g�HL�<���Y���m�v��D��a��ΚK�<1�Hr�D*��?gZ�­E�<AchES���5��JM�2a�H�<���R�XHz��,�3d0sQ�E�<	�c
Z-N-����	N��Y�EVC�<	��^�G��eSc�5H�����h�~�<)D��s��� ��4�����Gx�<�"�/r�QY�]�4x�@��w�<�VE�(I���uEl�N�
�a�r�<�V��#*\��p�D�j��B0/�p�<a�'��|D���hU�B��Q�<�A�X�����2<�@�ʗ�R�<i��ā@@И��B� �1��TP�<�g	�/ܕ��Yw��Y3�Tc�<�1��Q	�]����:��l�]�<�C#ޣ[�
Ix$d��*pRHy�\�<�ce��&� ����	R���JS_�<�1-�2T�p0��#�~� ��X�<�a)L�1$gr�}�B�n�<�qc�> 4`�㘎�1��f�<� �8r���s�(��3C��;��(�"O,r�hS0W|.Y�Oҽ)Cb�Hu"O��C���dh�F�@ـQ2�"O��ąC�"J�#��1�\��"On5�@k��f-�g��J��D��'�r�'.2�'���'��'���'	`��mS"�hͩ�'ń�4�a��'H��'e�'�2�'�B�'.r�'n�MH n�?f�0�S�*ƿ7��l2s�'�R�'���'t��'���'���'�h��� P8YG��cd�m���E�'���'\�'\��'�B�'uR�'��|rU뎏C���䧃z{H�b��'�B�'p��'Q2�'�b�'LR�'�ұp�%�RrM�$�C�\�X���'�r�'�'<��'�b�'���'� ����O#
�L�U�Y�!�(2�'s��'d��'L��'E��';R�'a���3&H�\�Q�$��4�p��'P��'I��'Kb�'�R�'4��'/�5S#̨fi�%����k#�'#�'��'�r�'�R�'�B�'��Ӑ�R�YU� ac�.&���c�'b�'*��'���'T��'R�'��ث�n�&��h�Q��N������'���'��'���'F��'S��'�d�J�d�s��:C�fŰ�	��f7��O��$�O��d�O��D�O��d�O��$�K*vPb��
3�� �X*�h�D�O@���O��d�O�d�Otm����	\�<��ތz�:�q��\�1�-O���<�|�'��7�F�>m�E�L�J$� 
#��1��x7���ش�����'2/�>��-U2l�r��ҩ��Uǎ�����?�A�M��Oz�;�bI?=F�@#i��Lc��xs�Eg�?�I�@�'��>q8R��8�N@�'�îj����D�݋�Mۖ��I̓��OY6=�����OWƄ�&�_�.�r�O���n��ԧ�OL�sV�i?�.^�ȭxS;@� � U+5W�}��� P�=�'�?q�*O�1��|��nH�9�
 ����<+O�O��n� x hb����(B��\L�`k@�0���ZS�_� ��IȟL�	�<��O��piݡ1��	cAO9!�8Ð������l��}��$�l�����t�fM�5f�B�v�Τ@�& sU� Gyr\��)��<a���P�����[1��0�S�Q�<���i����OV�l�d��|�o��sV�1�E��V-*t�����<9���?���n,ı�ܴ���v>=��'Q�.��	�7��ms��T1P�n5�b�"��|J*ON����֮ہ⵷f��<6(�a~�'j�F����$)��I�<i�P�kHZ+gX,U"�@�O����OH�B�����I. �j���E2���ru���ku^��֯��Op��~]��
�6�?�9}�gyBB�!�.���JxZŧG�@��X��'��'16�e��P��i� ��H�.ݰ���@X�E����?��<���?���d�+2K�6
�����́����%D��M;�'@�9@�'����`�'<�������$5dD
.9���c�V�-���X&:O����<.O?�F��.o��JW��$4)@E�'扦�M�Q�O~�En�6�OzA�.�~��l��i.� �u���'���'�E�~x�v2O��$�O~ �҂�(kT��N(Oe,8`��G��?ٰf%��|�+O|�$����c߅k.�k��v��$-��զ��3�7�Q��o��+��q��8�M
�!A!���i}��'��3OJ�����*|D�8�v��G�`]��Ds��D(:�p4��8�	�P9�hLl�ɅH!\:0�;��Y����=Y�D�	��Iԟ��)�SAyBbu�P`���j5vP��D�n�YC��:3|j�D�O�9nl��	3�MC��>)�򐄁#ذ;3�+0���$`�ؠKdq��	ʟX	�� $
���]Ky�G1/ߔ���G\�I�E���y�]�L�I����	柨��� �O�8uQ�e�'�<��i�/�(����t�J��<i����?��yw��;S�� [&Yj�g)U9.�6mH��%�N<�'���İ �ٴ�y"���T��X �K	� �v<x6���y�ψ�0��h���g�'��IƟ��ɚ�f\��@�?��Eb&�X�44.��	��������'�6mM�a���D�Oh���̀�@�O#
���F�W�&�$(�d�J}NfӺ1n�ēF�tM��̚�
������ ̓�?���M+5���2�������j�0������z��9K�"M��I�Vo,�����O����O�?�'�?9#ĝ�(5������!j\��3C�:�?Q�i@��2�'({����]�=W�x���>e�B����u�牯�Mӆ�ibF6-ҍ��6�1?13"�9o.��I
!*��:�g��E:hAzqڵ �ZH>a)O�?9 �S&KLlL�3#��x���
f�@g~�$a�,١��O�d�O��?��G䘿�|��N�,�b�zd�����$�O�6��c�)�	L:#��H�撁&���h́n� ���Q F��˓7*��4N�O�L>�,O��ţȢ9��S�F˰e�h%���'i�7�K�J����D _<���Sj_.��t��L������?�2V�P��4,l�FBp�©�g�	 HEi�H�5M�L��%L�7DCX7�9?q+�0a���)��'�� �L ��ޞp'fxS��^�����:O���O4���O���O��?������{�"I���A�Z	���������T��4+�d�'�?���i�'����d(Dl�x3CK"҄Quk!�dĦ	X��|��)�%�M�Ob) a�يa0��"��rc6-AV�|1��P��-�r�O���?���?���u�X���ެb]�,@e�%�v,���?�,O>�o�$@.a�I�4�IJ�D�˚&D��S I�HH�ⓧ����D�t}��t�Htm���S��aA�r4��o�'���R�%KET+����%�Z��-?���x�	?}kh:�4��H`�B�Gɰ����8�I̟��)��Zy�x�rxt
� d�fsD�9d� +�n�D�D�O�n�B���I��M!B�4�Ucr'��(10� ��p �~��� m���I蟴����;G��sy���/k�i+���� ��9�y�V��I՟���˟\�IП�O��L�ALK�|Ä�맩ӊ#�\�Aw�k�(���/�O6���O`�?����ӗ�F��H#�K@��E.]؛6v��$���?y��mh��m��<�p�K+*�@��S�ʁ(Z�����<�b�I7����������O��dS1D0pi�t��y ��g�NwĄ���O����OZ�g���!D�G���()A^6'21!]��읱��S�@�I��Mt�izO�d�4�	&c����4��G��)27O��ݭy�,�z0�_ �fʓ�Z+�O�p���O?N8"D�H"���["i�6*p���?	���?Y���h�0��3Y���%���x ��*ԳC����Ʀ�8�$Ο���+�M���w�$9��[�F���!�L�GF���'��7�Ц�	�4�F�4���Dy���?-���Ćb��@�U���
ߠ�³��-ec�'��X�'d8���O�Uо�I���%��L��Oƕo��B��0�	��L��u�'~\,bG/�>nu�����a8�tڐY���	¦�I>%?� ���q�ji@2�L��Ԉb�)L�t=gI�Tyb��=�6���$-�'��	;NWHAt��*]��x�k�D�T��	ԟ���d�i>�'9p6�Q�[���\�?UF�Z�C��k�r|�Do��aD��$�Φ��?qZ�d�شU,�6y�h��_
���ȣ�P�b����-��y��� ��(+4������UG����) WG[� �l���d�d��M�!	e�`��͟����x�	cy����8y�$�#�$�	=V�C�I��?]��'Fgӂݱ�7�R����%�h�D�°V�4�ꄤ�>O"�E��D&���?���|"��H��M��O<m�Q!�:"n�F+м0�$�y��W0�P���c���O�ʓ�?���?������L�q�[Q�F1C?
����?�-Ojl��J2FE�	쟈��c�J�3겘Jg�7l��%`�� ���r}�~�B�mZ����|���:`�8w�дy�8�X��ƫ=
v�*��I�bQ�r-Ӳ��D���N�T�O��rk�
�6qҷ�Z�h�pD�aO�}n�&�డː����y7�rN�	�(ڟ�I%�Mk�"�>Y2�i6��'(�>xJ��΅Y0p��Ɇ�M��i�2�b�i����(i> RB�O0P�'�rP�R8ĸM #��~T�h�''��X�����9(�kE'�(�����͂��M��aϻ�?���?����hq��.o���S�׾s낑p�gR�H!��n7�M���x����I�	{��<O� �W!�j�d�!�J�|e�y0O�P����?�WF%���<Y��?)1���w�I��ϋ�|l����?���?�����ʦ�b�`ԟ��I�<Q��ݚz�h��� �
m"pYy���b��X���*�Mcw�i(�O0)�u��.Xo��EO/�4D�u���3��˭q�m���t�S+q��I柠�آbuqS
�L�h�h!D��+��*�J��0�
3h��YJ��@��4
D�Xy��?��i��O�NC�-ͮ�(T�2A��]@��� T��˦�S�4v������&���� J� UH�D�&!F�|��Î "�$����=���1cPI�Q!�߫!��,1C�-' aTFE��M���) �lb�`��u��y�f�;M���mZ�wN"�*��6���B�!F�ޙ�v'E�P�je�B�ޥqO|H7��F�|8�ܱ T�	��Vq���t��jx�M��֛n	Fe�7�5W�6� G�ٻ(mIW�Qm�2ICG��V;�)���,6E������+Jp�Y�ve��KX��%X>-��ą�zc>IE�&"m�5���%VHx�A�o�b�&��QX�x�t�XS%�/�t����5Ml&1��i=��'�"�Oƺ�_�<���H7�p�Rl�-&�<�l�ǟ�I�]R���I؟d�IП��}
�+[5��z�!ט#���" ����C�IX˟��	ן���?��'X�ӣ.�@9˥F�!�Uk���O��y��4C�������H�S�O��.��>ɢ� ��J)a̲��EO�	?S�7��O��$y�|��'�O>���|����~-�L�ab�FR�d�-)�D>
.,c��������'�?i���?y��+a	��Fq�x���eɚyH�<Ok�'~r�~���a	���Խ u�]#���:*E4=l�>�U�I�= P�'V��'.R�'��[��t��煦�1JҬȖrl��u^�H�'dr�|��'e�NI�s�耖I�g�$H�@�?V�:t�S�����O�D�O0���O��H���?x0���M �e1`�G�m� ������d�O.�$9�D�O,�d\�#�F ��iR�}FXQ9P��0`i�1�O�$�O����O��$ƍg�����O��d�..�0"9{�ļZ�� =kT�ao�Ɵ�'� ��Ɵ��t�S'(4�O� ��y�+
[`uє�J,j�֑���i�r�'�剨g�Μ�O|�����B���ˤE�!eh���g�R0a��'���'@v����T?e9aХ�x��c���<�qJ��qӮ�_m �aҼiE2�'�b�O�����S� F���kX�G�D	���ۦq��ȟ�%��؟ '� �}��A�E��у&׭�t�x���)��M���M���?���2D_��'�`3�얳bh�KSF#f�@ �Cr���� �Is���?tk�+3�Y�Эh�J8��iކCۛ��'��'�����>-OR�����b��#6f���ĝ5O���"�n:��&ֽ'�������I�k��$!��N�w��M�F�6)UzX2�4�?I�GZ����dy��'8ɧ5��Lcn���`�hOZ�����(���ԎX��O����Ol���<�eET2q9�\Ru�
�lX6Y��ˁ�K(�!S�S�p�'��|��'AN�k��q�OC�7稘X��܊�)�|�'���'��I�k�p�0�O4d�(���g�`1�!ݑ7F5�4��$�O�ʓ�?���?�D8���o��m�GB��� M��d�Oz�D�O@ʓqN��wX?��I������@?Z�t��@��B�`�;�4�?�N>���?����'�hy��d���Єp�.	VN���4�?����N+R��y�Od��'��ӳ$�&]���v�Թ���0]wVO$���O
���$6�	]��$E 4E���;�
�3-����'@�X7~�6���O
�����ק5f���C�$��B,�*�����C�M{���?	����'q��[���bH�����w����i���(5`i�6�d�O��d�!�'��<W��A�X�|���V����I��Md斡��'�����BX��Z�% c�4(�2�HO�nZܟ���Ɵ��ĉ2���<����~��T�O�*��PO5�N����?��'��l��yb�'��'�>I�&�^֜��"�r��(�E������p#�	'���ɟ�Iyy2�7%e@AH�cS�ʫ��D�<en���4�?��J���?,O����O��$�<�dM�%o�R9Ã�� �HYQ����]�ўx��'hB�'y��˟���6-'��@�3�P�3j�:}JX��������'���'"^�l`ԡE����ѡ �~��$)M�B��"�C����O����O�ʓ�?	�7z���UA6\�%'X�e��xr���>B��aj_� ��韰�	Ky�c�O��n��©N�]4��Ua�Bl��ӌ�����	��(�'�R�'�,�R�'�'��,��̭!���B!��3!w�\o�ʟ,�'���wy��ݟ`�	�?�ؽD� ����d�R�qT���Mj�O����<iЃ�w��uǎO%Dbf4����LJ6	�GB�����Oԭ;�)�OF���O:�D�`�Ӻ��O�<m�z��gDAe��x�s�����	ϟ8¢Q�p��c�b?5(����x8��7�<��4�0�{��<��O&���O�D���S���*&��$��bB -��)�)�Ly�7�x����W��S-/I���'f�^�"L��J*V��ڴ�?	���?)tB����?�Ox3�c��3�.	��.#�1l�O�@v2�Ɠ�T�'���'�rX9 G��q�XB�b�|����Mg���$؃`I��$������xyG�|�@�0V�E^"藣]O7M�Ou���OX˓�?Y���?i-O Xa��҆m4=��`ϊ-X��
B��]	�`$���	�����byB�'b�ސM��}C�N�[!�X㫖*j7
�`D�'��I�����'L����͠?%[�9Usҡt���Q�� _���I����@y��'��A�/
�%
�X�f�P���U���V\���?y���?�*O 5JQ⓼-��%a��ݺzfD�0�� d�l)޴�?AO>�*O ����OZ�O)��ۆ�N<�4h����n���4�?������;?�&`'>q�I�?�؂I�P���~=P����D*#*7��<���?!v�E"�?*�����kLZ8Q��h�d�$ �EzR����	�����	���	�	�?��u��]9��)����Q���7@"�M#���?)q�����<�~�Aȟ/��85�ψm]���&��=�� �M���?����"v�x�O���Ң��*�q���@:�����s�n�p���O��d�<�J~Γ�?qP������3ӀU�}��h��웈V���'g��'�v!Q�#�4�X���O�<�Ã�O�"��w]�\��ك�ަ%�	��j�T9��L^��'��'_R�A#?�����xd
h[��/��7��O�yY��A�i>��cy�ڟtHa��4K�@�P�O�[��1*�Z��X�̟p�'!��'h�Y�L֍W�3;d�p��&hm���I�Y�z5#K<����?qN>�*Oҭ�H']D�)�	G�9�Ҁ�FaӫJ����<����?Q���$�B�Χ�Aq"dO�lM �V�F�=��Xnpy�''�I���	��XC��u��R �Z�L<���+A<l䰤��2�M��?���?Q.On�xP�H`�$��5֯۰IEb�FB[�9Gv�s�R�M���d�O �d�O` S"?O�˧�f�)�B�>4�Ik�E^$�:��i��'��!DgܴR������O<��J�s��5����?�Z$y����~�p�'���'��g���y��|ן�q����1��$��d��^�(`Z��iZ�	����4�?���?����i��ɰ
ËV��x��EK�~Լ9��u�T�D�O ��4O����y��� (I�
L� �k$�
�����i��@�i`�J��O���� �'�I&T�a�F\�C��I2����o9����4S,9ϓ�?A-O��?U�I &�lX!�Ȍ	�����?SJ��Voc�R��O��d��`�'3��x�b��l����,~���B�L���l�؟0�	՟�B�'y��'�?����?Q�i�>6�
���oK�j�ĉ�",I���'�= ע�>�,O��ħ<�����jJ�t�b4h�@�_�P�[d �G}2_�y��'2��'R��'��Ɋ8x��'9Y"f�BhW%y�ʸs`)�	����<y�����O(���O,�v���(����r��ei�aC�d�Ol�d�O����O$���]�26��B'��a@����
GܼYv�iX�I�t�'Y"�'�¢V�y�Χl���G!Z٢Q��C.
s�ꓔ?A���?�+O�0�V+�T���'���,پ{%�<�C���L��oh�R�Ħ<����?A�HS�0�>!�Գ}�%����}���au�Ԧ��	�ĕ'�D@Ä�~���?��'ZϪ I�&e�<�Ӡ	�TX�b�T�,�	؟��I�9n�'���?m�\�������T"3�4�5Lf�B˓<պmXԵi���'��Os��Ӻ[F��4 �!Ç18�M�ܘ�M���?�B��<����$,�S!��}`�ɕ�h�<�QT$
s�6M��%-��nZ�4�	����-����<'��,aqĞ<l�6����J|��E��y��'\�I@���?�a��o��36��'e|<Ũ��#kśV�'���'���j�¸>1.O�����,)A��>T�T�#��g���ad�w�(�Ī<El��<�Oh��'Aߥo-��R'n��p�A�ǫ�;/l7��O�`�Ia}BR�l��VyR�5v(\���؄L�O�X��$���M���o"���?���?��?9-OZ�ف�>2r��t�f�����Ǡ7�Э�'d�	ן�'e�']�$�2t��c����6: �S�g�@���'��ퟨ��ϟ8�'�j p�gd>5�E'�H�昪��_��RQ*v��>	���?�O>��?y#n�<���8l�$[�OB:�R�!��#74�i�l�ן���[y�������1�-��w �xb��l��+�ߦ���G�ן��	�g���Q��}�|P%ዛ�p|Iӫ�iw��'��S��⦪��ħ�?��'u��H)�`�xRĒ獃9B�p��ǔx2�'��i]+�yB�|ߟ:��"=�XI6#�6V��� �i��	/L��9��42��ߟ���=���VB	H�[3��"�a�)�V�'j2h��E"��|B�)��R�bI��.Ӕ_�^�s��H-Qv���IU�7��O^�d�O����{�P���"mՀcI�]��_4����0�ip�,#b�'{�'%�0��@4q�X�
�!�>_�Pa�"Enl��oZݟ��I��U�M���'��O�	�c��%j)�ŮT�E�u"t�ir�'�*e�e�<��O��D�O��GOC@���LJ:{O�e�qh���	�_���RO<����?�M>�����v������㍊1���'�lh��'R�ٟP��ɟL�'���C�],Ck�ݣd���D�^}�H�4f�c����]�	����	�N��$�ʗ�g�nٸ�5UČ��S"�\�'���'��Ol޴;&(n>�I�	,'�T���܆s�sE* �D�O,�O^�d�O��iB��O�8�U�ƃH�jI�&K�9Anԁ�F,�T}"�'���'��I�S�f	 O|�� �T�y� @T(l�� lބnP���'��'���'��E���'�p���&��e��'_d���l����py2%I�p0b���d����:�G�}u&��#�G$Ț�؂ia�Iϟ0���ޤ�IE�NJфӓ�Xh�툃V��<2 ��7��<�<?�qӄ0�OJ�O8�.���V	��X/@��!DB�5�'	Ҏ�@��|�����,���nQ�Cv���3��Mk���W�F�';�'E�d�#�4�d酤	�W�`!�� �6���S�ey�#�ɟ���fy����OP�wd�2JW:$i ��p�"A1��䦉�Iş��I"^ٛ�O:��?)�'�>���WA��0�B�$"~�!
�O��l&\��T;��'�jI�W@Wj �ae�H��Xu���k��!
���'��Iޟ4�'�Zc.y	�N��
س��Z�v�"�O:�8#0O�ʓ�?����?Y��?1jkj��(D0r�HDv�da��i"�'���'<�����O��1�fV�vp P���7x]��[O��O���O��$�Oʓ0�@�7�h�1Ǒ5����"Y9vZl�R�in�I؟��'or�'`򍚉�y�&N�Qܤ A�Q�}=~i(D	�	 5�7�O����O|���<a�A��j���ϟ֘�p8�g�-��<�#o��kF7��O�ʓ�?9���?����<����?	��B��:�Oб>�|@��!q����'��W�����������O����$�j���a1`��2c��wUХ�#c}�'���'(��'��\����9<���8'd�}�tJת_�` n�gyb�Q,SP7m�O(���O|�I�j}Zw�DyR���8(PH(�`D9]_\P�۴�?�~,4�ϓ�?����?I���n*R�t1C	��&��²�Ĉ�M#��?�����Ov�'��	(Rnfm ��9��]�Ab�s�6�rݴ'�ؠY�(�H�S�O�����S�4rg6<��ۓ �	>�7�O��D�OB��1�p}r\>��I��D�S�H�Q���q���������a����'t��)p�|"�'PB�'8F� �P��ƞ~,6��SQ>���i��d��I&����O��O,)�O�X��E���B/��l�2��u}B�[��[�O|���ON���<����!]��d2��1g��/v�nDI�␐�ē�?����?9)O�$�O�d���C�B侼�cg��7Ҽ�[�.D;#1O����O����O����F��C�M�AA{jFU��
4v�P�ݴ�?q��?N>y���?��&�5O�n�3Ȑ�S�L{���� �hU�꓾?9���?�*O�$�s�c�4�'Đ�{�&�v�Y�j�s\@ ��j�����OT�t���l�y'��A��!��������m�ßL�	�D�ɨ|Nt�Iן�z�O�*{�ֽs1dT�]{l�k�.Qmn�'���'�*ܑ������i�d���!M�b����6,ϝPh�&�' ��C*v�2�''���D�OkC\;XQ��WP|�[��9O\�����7���;�h����i��FS��r�
c��9$�[q���!�7-�OZ���Ob�)�u}bR>ŚbJT�| ����LW�-i,�#�0�M�"d�z�'����|��'���7d\�\�<��Gʇ%9�(@��,l�"�D�OB�I ^���O�˧�?a�'��	Z'�'(\�H
o�����'�	�6��DKJ~�W������Q�V�L���\P	(��͓X\�B�\�G�Dp�ׂ��w��X�1z|��dƦ(t��ȦL� /�%{��Z%�z�'Hj͔��$���� $�)x��	���h�I�CBt�M"f���o��� ��?-0���&�#l�Zv��D��)r�D"J���/� X����J�B��G"��8���%v��}@��4w0H�9a-�
L=�
�㋜1���D$Z ��Ey�Ǜ<H�Hx�ł�|D�3���?�	��iA��?��O����#��C}��G�	O�������s�ϐ��A�u)�?V�"?qU�ѡ)�p�w��|�~@����>���ZN�W�(t��┊=�|$:cI�e���0;��O���<��aI�q,"%j����Ni���F̓��=)���i��%�"�,\��g�J<�6�ig0؀b���W�\��GG4���˛'O�I�l/�೪O��d�|���B��?A�N�\�.���	����W�L�?���e��<���P8NÈ��A%�>�O����\M��H~)��;%D� B�>�����A$ȴaB&I�.�Q?��!�N	!<� �� &��	� }cA��?���h���d��d�:��g̾t���$�
2�!�$Lc�Lu)��2�����ˁ�ax�E4�"X�(�	Y`��h�I��H��!Z�H����ph��
�L�|T���	ß杌v�����e\-mB����2S��pY�m'_0=��d7r�J���L�g�	}@����G�zm����n�6l�fT�_��I��Pc6��ej'�3�����m����
�qр.U>+4��9?ْ]��S~�'�dQS�QH1�B��C�k��8��'�)rՃܲ8�]�`�$j��9�O��Ezʟ��l ��Ą�2i�Z�Q�ɇnI�<{f�c��(����?	���?�Դ��D�O��S� �h��̎L��5���0d^���i��e��[+4oZ*�'�e��� SFb�yF�R�p nq�R�[���D����k�ȈsX��3$ꙩnH�1���ZŁ�@Eo0.�d�OҒO(��5�s�<�F��.xCH<�M����uHv�$D������T0�b!���B�^ �tc����4�?*O��z���Ԧ��ȟ��T�D.E�D��*Ke��d9̊ן���(4\���	՟��	�e���: #�V��0���M��b�\=J`��]�U�l['�z8����g�;E����oC��h,m�$2�8ٔ�W:�>���N����$�_y���:���OP�"���fr�e;uoġH����Չ�<1����'L`A��& �E�&Z��s�i�)CJAZ����|E��!�'>47�Xw%�|1�.׫T
8�B���0�'�@e��'�0t�gӚ���O�˧W?�a�HV�b�^�C�8��P�D�n�z����:o�%B�"�)�d?~X4���#]�i�4]�O��S'%�"�0D.ӆg�����M H��'���������ٟ)��G�ģ���J�����XΖ��B	&��w����5�)�� �&��3OX�yC~t�s&�&g�C䉹4���`{vfhP� ����$@W�'ն���4^un�а*� �Ȥs�M{�j�$�O���^<n�m���O��d�O��4�8��A�Ћ0k�x:afŭ-[T��Ҡ�f�5qp�c���q�I=L:b>�O�1AQA �D��˰.���"��Q�$y�P�gn�#8��T�� Q�q��'o��hvm�X^��6KH(a�y��H)a��L>� ���N� S���-,��6�_�<�c�3h�Z��so�		���D�^~!�S�O����f��,Z���HK�>5�n8�.^|�R�'���'��֝�<���|��՚K�,��U%`�Dp�!�O%Z=��h��J5��8�R 9���dP�p�'Sq<qu�'
(y���s�.�;��ŝ?ua�	X����*���)z��\5fF�)S-D�� ��&�;v��6́�y�����$^E�	�0L�G�i�B�'�Ԙ��ȈE�Qfe�5\�A`E�'�r��#e]b�'��i �sC|r��b��x�u�ҮY����r蝦�p<��\�[�Z%@4v���Z(szy��I=����<���R(i����BVmI�k�!��=/g��B�	Px�$�Sm��q�!�$�¦�s���m��A�5�/R�@�rWb�|�"u��z۴�?i���	�i����S�H��C5�lks�E`�*�$�O}x��OXb��g~�
�)&z�шOS�)l���ҥ���I7-?"<�r�G�.$���`�V4,��V@�Y�d�/�R��i]6��	���Y�z� �gN)T!�$ÝU}x��Wd��Z��!� ؜9ax2l:ғ1L�,���E�U�����%��^CN9XӼix��'����*C�iZ��'�b�'�wJp�b��&K*IŃ��\i�$3�;�dS�j����|R�ձ{Td�h��N�z:M1�k�g�Ѻ�a�w3$tm�6�M���|r�ɳMt��I���laŇL�
�1O�|a�������A��0Ӕ����̣��I��;�"���F�_��#�C�:��?!�i>$� �vdM�EI�Q+e@H�{��xb��[�oN�R�\����I�t�I$�u��'wR<�0�Y�j��P$��t���#�(�bD�m��YJ��do��p��!<OH�+R@�E1Z���^2!2j�q�N�iaD�Q�eI09b*�Z�E*<OJ�Q%����vi�8		���&6o���'0v�*"]�n��ڇ̌�*������DD<�S�$@^�l"A*�-5���l�ڴ��H�����ia��'|�C�S)C2X��Y�bY�u�'�#S�A���'G�	�2uU�|2�@�g�\prh�8KD����p<I�F�x�|�4�h�a���#��=2W���㉡+{��D)���OL�a5��K�\��Qx�!�d˶s�"��0g;�h�&�+FX!��ɦQ�׌�J @��m�J��[�f(�긅S޴�?Y���)��JC2�dU�)�(�q� _�i�LE�w2L�D�O�M�	��]���Q�EX�����t��R>Ep���"�rYq#���4�m�$}��#3E��b�z ��5�0ʧmn@a�D�-;����LU ���Ot`;��'���t��T��2$���� �n�Bx[#�J$˘'���'������K��b�bB|`�Ó[ۑ��b�ɏ�6�fe��*�*�*HR`���MK���?���V�t��P����?����?��ҿ�3�{!��e&F�S�Oɉ3j=	�O��yaE |1��'����"��Y�@�x���'J�Qo�������Iզ!:'3�q��'(��r�Y%q�8 �F?�p�e�{�~0o�ܟ�AЏa�n:�<)�g-�qk�.˹_n�E���*q7h�2�'��hY�V
��Pc)V�D����O:�Dzb�F?9,O6!7�ʪ[�|1pT��*`���(���*�pBN�O|�d�Ol��j�4�'��i>X�)����_Q�y����g�j�b��N�a~n�?iJ�r%�Hlվ�ba���A�~A@ ���0?i@�Z!PE����U�h �"���ޟ4�	ş �'i�ґ@K�ArL*;4����g�"O�iE+��U`2�{0��e憘 �d�d}Y�HC� �=�MC��?a�ܤW�4����P�5��=� AJ��?��xN�� ���?i�O�������Xf���F�p5���3E��ɢ,	���&��,MhX��?+�����&O$�!�'��'ܠ��ďQ7d��� �)V,-ܢ\��'��z3��z2�(/;�m�S��A<a �i�H���1�n��2ș?It2�ʊy�!DHr0듕?y/�h@b���Ob8�@ճp�v�8%�T�h|،�@��O��dEb0����E@�}���WgT*�M�Om��-ǺE��i9(H2-S%b�L�.�'V�#e�ɐa�:y��&U*\�ƣ|�.�w��g�K����.�E�$\�n$��'�>���!��s��߾z��Yʄ�ڮbK
���=��,*�ۉ]��L�8�$I�቞�HOd�3ģ�<]���AdïI�(��E���1��ޟ�I�?������`��ޟ$�iޡ�Y�w�DL��E'{�rU�u�a�X��ٲ^$ң?���6 ��y�F�U�NhS"�O�̘'���J��O�g�	�d���N�fZz�{O�23�y�	�0��8�D��)�<i�=�L����0q�>�(�K۾h��dp�'���h��ց��� �A �Jsl9�ONTFzb\>��� ޴��ܧ&$��� |��r�X-6���yfb�O����O��D�纻��?��c� "����`��d+s����\;�|Z��A.0I%k�g[џ���|nZH�n\�}����'e
(��aG�	c���pDN�G+�(1CLQ� �\	���:��
�<�B@#`ID,h$�0��u���
�
�D�<�����'� ��*E�BI�@��0z~pej���.ړ��3�4�C��QX���K�����Oz��G���1�4��)�(D`o�؟��IN<���dy��z�J�1V��E����p�"��(�I̟���BU9M�@{��+c�ZQ��e�sn���ǡM9���Q��8 ���H�I-7>H��Z�@��	�ʊ;4Xa�gt�CG��q�6� �����O�����'�F6�\ʦ��	�i����C���'�����^%t�a�'V�H�'�4���ʄ,5�� ʥrJ�-�
On7m��a�̙�'A�
?!���3CL<c�F�o䟈`�4�v�0_���	Ο$�S |>�����Q��,`p*�L���E =/6���ڟ`�c��$7���@�c�$P���)�|1�OV���z0�`��]��*�B�^)��q���Y!D�EP�\B�O��Pk�� !�d;�	M�8i
H��v �O0�d0�'�?��%S-Z�(@����`�
VAb��	�'�5#�Oǅ����� �쀳�ő��I�e
Z9$E�$@��d��m�������O$�$�7~ 5��O����O"�4�S7��W��C"�������(e��!1f˔�C���̳m�c>�ON� �,�<+]�� !� ;��X�	I0��T�%7wRD�p��C�q��',",��d�"2��P��Yd��2��'��ɬ'���4���$&�I�-��tzEY #���f��<C>tC�Iv��$ʉ\��ō6G��lF���'��DY2z}�`�*-����E��2X�\�@S:v����O����Oty���?����?�,+��e��h��IJV����ƟG,����,'�OP�+ҫ^cD���U�W`�4PѢ5� �XT✱a��G��_X�D±�ɐH9��H�H�Ԑ�egͽQH��ě��� ش�?	+O��D!�I83(�1�)� UV�Qf\τ�I[����|���&�I醑��@�JO��ᗃ'�DV��uR�4��,QW@�o矰��':�lJ��Ŗ �h"j�������C]�X��Ɵx�'u���*�Ď|�I�-���pf��)�h�C�Y?d��񤑦&��Y�|��_�e&V��]�-ĭ�EÃ��p<Qe���P�4{���':t���F�b�U0��Y�93eS���	M�S�OB���aΦBN\�C���{�'�86�S�$,2�R �-::�����3zC�<�Tj�4����ДOl�12�',�aK�d��`�+�!���'������ڭ�/L��8`�^�r���	��;�8�r���mj�H��D]�K*��0����M�Q���ʗ!�gZ�����+�!'��I(�"�-!���+��?ZB"��O�}B��<|D���@�,>;Ҡh�J��a%@���'�]#��ЧpD��!�J�r�:��'��"=�(�* �~�Y�nź3T������2���'i��'pz\����UM��'��y�擹�Bh��ip�Xx��?Y>*�O½y����I�Ԓ�1OBLJ�BAY���ʠE"p�DD���8Z���tC�M�9�q��')����5r�e��B�\+h�.q�6Qn�ܟȩ�.�ڟ�>˓�?q�k_���	G�>� tr� ��xB����d~B�'
�4�}��Xm�@�ɤKS$$q��V(F܍�Tcӯm�B�ԟ�z�O|˓�?��'�?Q.OrA�`J�IO6p �-�;��p�P"OP�1)ѱDz��ϗ�5�A�"OdMUv\+�%
c��Ya�!��y2���\�J ����)�Һ�yr��3������N�iۗ���y���4&����� ��xB������1�y�.AD�%s��\�r誑B �	��y��τ7p�`����d�"(#�L��y�FE�K���U�	/_,�{�e�:�yN� V8 
���	N�֭�2����ybƑ�m��$�W���)@rG��y�ʌ�o�I��]�m�q�F�ɮ�yB�ٛO�$C/}F��Y��y�fÑ'�������B�K�o��y�������挚�2��Z��h�ȓJ:չ�A��ל��%�8lb���|� �p��'����ܶkP��9�)i@�\/F;�8g���^E�X��S�? *q��Ñ6@�"7Mѐ�X�b�"O�8��(w��5a,��Bya"O�m���NC�$B�؈=����"O��`�A
�fm3Ђ-[�N�*�"O�L��H/6ƶ������Q"O��cw�[Kb��"t �q���k�"O����'�Ҝ�yF�Ŏj�֑��"OfHʤO��0m��q�Z7vkC"O�L
���eh`}qU(Dz�Y8�"O��b5S6α8v���q%"OdD�!kO-w���S��|�d�'2��pC��,A�T���0z������!jV@��?!@�(�0<iD�tll����4Z���r��f}bkå7\�Є�	v�H��Sa^se�	*�
�sb��[�;|��z�8em<�	�V�h��A5��̐�@���O��Ā� ��~�	�M� hٴp�X] �����a��"�MEz2`Z�6,.F�4��2Dج�D]�y����D�X5t�(�E�O��ё�|�n�|
じ�*h�R�服�U(�L��}b�N�e��Ɍ�3
����!���5f��qw ^>a�4�s�8V�:�'��7ޭ`X��d�	�=����7��'˘��!D���0W�UY�θѭO�%ϕ�:,2�(I�b?-a�o�u�Vu�2d�?��qI�`��T�J�Sc`EoÖ����$�ў8�d!���y7��:T ��$��)�!P$�8���R!A�(X�1��$3�E&��ASg�0,�xb�0/ݫ���>����k0@8V�h= ��IW�A���/M.4���8[qSu-�O���*Ps�	���iD4&j�m�;�z����D�h��%x&��6x�T!oZ�0�Z��%E�DOd���
$��"?�ňO�Gq�=��@�<.g��hT��K��y��5ՠ;W7�� ��G���yR�_/� b�ƾ5����B����P��1|Od<3�'?��£ɫ$J�E)�bZ�[|tѩ��	|z��H��O�b���D{R�?�*�R���3Ï��,��x��憛V�:�>!��^^�O�@��GL�w���������7�I�y Z	�'.�8���A��f��1����j޽B�҈`׎��B�Ҽ�s���N�6��ӧuO����͸A��A
@��>X�m��
S ��ڱ�nӈ�A���-�V`��З��Ѓ��:�>%V.L"I0�t{���i[��'�ɔm���s�!��2��gyX)V�c�C) rR �R	��\���fm/|O0�K�w("�PAȏ"_dY:�%]/g��3�*�/U��"�M��ܑ�8���������R=�
1��E2' -at)g��;Q�9�Ʌ`�>h1ݎ}����G1eV�t���D�+<`f��O>a�I�)]��M2��-5�ݲb}�t�'I,�d�p�S��fI�~�:��f ��f�^�I�� �<Rى���:>@$�^��ų�_f≿�1��)����I�>��[u#�����׃7���O>���'��㋞���અe�NܓB�K�K�E3���r#��b�8��'f	w�G[�Hp�'B�O�E���zC�Y灅y��!���Ķn,l��3��5�Xɓ�"�ax�C]�%|�lpI���Cl^Vmp�Y-f�$�)O�x'����O�qOĠA�M�V���b��[?;=��
Wc0Oꕂ�Ni�	:�ܙ��J_�Wc�%Ba#��c������<i��'Ҏ�ʧ\��x��\�z"�[���70�ЪO,��Uq-��%A���?�s�n�
�S�~��Ӻ���B�@&�3`��g�@T�C�h򉤧?�K�k.,�*l��6�[�'n6�ڔ
Nz]�b�n�p�bK�O�#t��%i��?�zFB� ����Ѡm�`��Γ��Aٵ 	�^�z�Ғ �_���ƃi?Y�e� m�V��˂,7�j�D	�5���%m�������Oܓ���tj5���[�K�WhH���-iC
�������0!p�,|Rt�e"!xZA��+`���츧�ia�Z@��3�%�]�pR�`�1~�
|r`��"�f��+��'���<Y4�� �>8��'h�L���DjC����N��w�x�f�O�:G�D�i�2���X���'&Z��!탕):J�!�%3��H�'R>Y��˱�,�%MT"S����'}J�l�.m��hٴ#zՀ �.b����E�y_��;�O@-X�����Ě6M��|���w�\)�a j�	Ņ 	{:�b�Fѵ"�!c�H��)�0��5���Oڅ����b�K�w���( 	aJ�Q�(�$�Ɏ��uY$��U0���MS��m�P+���>z��TunH=�v�v��18�H�R��!-o�Q)�����s�F��rh_�1z�)b�զc;�:�gTm�d��&�Pl8�k^����T?�Ro��_����%̄<0�����o��2�������C?b2���5ݟ����}��N��M�U@Z#BbaKps��w�L��ʟ4	��%1?�s�O�ZQ�f�<QL0'�7~��%�դ�_�f���1�|�d^(�y'��1	1j���Fd���zq-B���7Xѐ��ՕHi^��'ɀ ��'3JT`�HbLM�%&�D/$"*9Ҁ1�@֨dF��yB�6Ǧ��c͔!�"`��-ti��"[>��bB�0Mv��ͦ?�C��Ҽ)�J(k��!P�8L���(,̙v���np ��3扐f`8@�Ҧ�N��Ð@n`x�iV
Z��JS�WB:�OZ��BC��:���7f�C���s������-p ���8n�1O8�U�:j��a��o�>�+d��6�t�G��S�.;E���l�FG19�؁9��T>]2r�C����.�UтJU��P�\��^)����L���D�,O��#���`0�5�� #��re�5� c���pa���ڨ
"	�.�b��X��92��{U�*f�����ߋ160�cC+޲S���"��)�$Β}�� �Ù�a���gS�Ka�\Z�.߿��ͣ��\^2T��݅uj��iE@�:�b��)�@�>wܴ!`%B���3c��00��x�3��,a�#"��:s9�-c�+Rs�jW�I�W�qO�à�i\:h��1�}���5�]HQfA����F�8��l��⑴i]*ȉb�ZU��AD�ަ]�H�ҭ��h�qO�(d5�y�;5 ��'�%p-�P�&�I�E���Q� 4�|BU�
�<d� j���Y�p�p�ҭ��@Xd���/�V�Nb����'�RN�)7n]�
�M6�4\0s�B%�ĉ8�l?Ebɐ��!`4��M��W�&�O4��E��@&�Q ��,i��%�Q�\'�y��ɟ
,}�Q_���s�ɋH~����
!�l6 ��Fȅu(����w���&#n�ƍY��e8��Oƌ[��%��sC�\�1���ě��)���؅ *j=�s�E� 1O����L�<h,�yb� B>�!� we�98�)O� ���rN�:R�rasS��S��	��T>5������5�Z�X���&@E�ԌI���%y�>��7�,Y'T͓�yG�,Oj��N��DL!��xY��֊(�	�8٨�҂{�uX�F�4RP�b� p�O^�G��H�-HYC�����#�t5:��I���зd(��Y�P�ҳlݼ 3&C��E���SƯI��6�+a;4��	Z�&�%|���Ug��2�Vb����c���Ɛ����!d��c�EH��Te2@��#Y���ۑ�"���#��ٕ��fل��EECdqO���� \>��#����+f���;�R�j�B�?ER�c��S�LB���*Ыd�"��Q�F�E�V���/Ԛ
-�HB$_UqO哭F2�̻Ǝaq"B��e�!}���KPG� P�%[4+VF�	z�#|�'�v@�^k�$�D���{����@�A̓;�����H��]�X�_2	�����?牢w�x,:����{�I���^�~�x�5��r(���O�:��O�x��g��oy���'6Ѻ�2�y����B��W��c�[�jc�Q�#���*�������Is3�4m�!m�l�Z��w���$@>2P�9���(_G�	
���'� 㗆�A�m�3I��)�x���}h��O��)�E^�"�T�'��?'����@"���#*Y�8��q�}��xDCs�nޡ:�'C4|j\��@J��b��Uk9�ɋX�t�X����L�"M��݄I�xvg�+Z�|�9���J�I�4��� ��EG��3A���v���2u��k���
Hh3ˋ�y� Q�	�v_���s0����0}B	M��deZ��d�@-s`���#S�!ZT��*f��6V�Z�"4Y&M�$�Z�-�d������-�<����W#	�`��Z�l`ҁ�=m2<��'��5z��Yg�g�I�F�@��h�(h�S'��#�$*�9poP˓2�AΦ���4̫J�3��D�W|���hA�%O�ei4D�A�=����xA˓(@>�]=�z%�d!�9>���5%�0`8���M�+��Ӳ�+\E[j�S��O�0w�~�R�̟s`�x��'�p2t+��^��U��ד$ј��A-�$,���F�*oN��hÑ\T�M��B��`��6�������S�ڻ��8�� ��3w(:�ʧ��V�t��'n@U�GR!k$b�x���X x<a�U'�~�Cg������W䵫$b�jMt0ˀ�щN�YuMn�آ�L�Lh�&?�xX$�M�I-��3�h�$Z?>������՚ЪcFH�u㒟eҀyZ :O�I�[�-�'&E�$��%O�4�rw�2nҐ�!iB�b�]� ESK��Hؔ)R!A,���4FE�̊e,�'24RDb�Ik�ڌFBs�(S��)�	�9��A���ۀUˢ�F5<�|��f�����K4q���c���E|�!J�C��f	{�`��X(HQ3F�ւ$��r��>�b�@����!O�I��o��,�tn�;BN�5�Ƭγz�3�)��H�#},=3�eô%άxC�Y�FR��{R��u'̽RhڜAg/ޖ[�v	���T2��)�����l�ag��1	�QII|�>9�@�KDM1��œ?Jh%q�煸)ĺ�I�4c^=���G7�N�9�0��Wwr�$�����p�G�)1��q�/ٍP���e�Y
K'z��'_<��"Hߴ���1e��+$x�1���k
�l	�H9��0E��C_,�����<�򏎗cj%�͊�2x�D
� �p=�ı.�	�vy��,S�>>v�²@��
�m�O��d(��ƬWP�!
�G#{����~�v��N~�s冿b:�	�f���T�@Ԍ�\�V"R *�C/��;V$TnMh���Z�F��`��hh�ؠQd�/�ʬ��eժN��Z�v�`���X�g�3ʠI���w �}��
�[���r�X�	5j78{a�R9tiq���2���O�����36|��VPM��BP�[E@!I�E����ŔV���W��S�U��͛��Z' �g��$����
�v����
���Y��Ks�����X���TkZ/$@Np�1O6���MO�Sz v*���e �� �I9PJ�0�<B�#L;bd�Z����C%��B���`�ҕc�@Ǭ!z�h{��'��=@�+<���1C[��Zt�O�^���²n@bp�	�B=~x	�m͠dD�Y:b`[Nb��S�nt<U����-k+�h#S������ǲ<�"�M:th��N~�=�@��qq�:f ��x��[�cG�I$N����#� �&��Oq�(� ׮`X��	΢�b��Ma�m��JW�j<�	��b3�)�O$@�5f^�Mx@�"iڸ$�(���� �剄)c�e��R�� %�Sa'ZX�iز&X�E8Ք'��Q�D�ѥV���i���(��g�'.���m_�\^�B��Cs(L�$ͅ	=�$CA�C3`28�@�W�}R\�҇@�P�.��&�1�j��/OP����+G�h���ؿA#e��ύ'��	�?F	�͏;G��\b� ���O�)$|R�[��\���%��xO�a�wW��������%?�����*��cV�m��cnRL�c��|�`�O�@[��&�̄X�8�e�Y2P}�UM\����ƍS�^�Ð�E��pc$ȂS��5qA�*PE���%-��i���Q*@;�J��xj�����Č5�\@n�fOB�В���h�g�Q2ذ�IR-n���:�D?O@��Ȗ�jp���ǉez`5ӷ5)���*�O��
�rUZf�A���P��GM�B{H�ܴNü�p�?�)�I�|�����<�pP8ve�?��{�Z�t�ڴ?��(��'@q�T��O�>7Ё��a_��A��G�����<��=Y�Q>�f�nAh��ԫzH��c�2�N<�ȓy�l8h�$����eÓ	^}�Dn����{
�}���J@G�lN��ek_�b��ȓ:5"�a��p�Y�}�BŅ�R�h�'�5 ���S�x�.��-�(<��eS,�`�P�� mA���.��2�ɋeN4���<{6D���w�`����A�E9n����ȓ9����D�\�N��V�]Y���ȓu�t���D�m��b��;��ȓ	*��q��!2�8�e*dp4��ȓc�n�kq�B�2�!�&W.��1��i
�qd���%�B�k!�dr8�ȓ� ّ���YŚl�F��]h���Z_�]I����0 ꏱ��`�ȓצ�04��#H�DԪ�+7������������1KB8C4!z®��ȓ�da���Ҙ
�<���,��\o��ȓ>z$����Q��h��n��ȓ^TH�K����5���X�J^�x�2���}��}�dM�
+��HS�9�C�I:���	w!��A�a�	�@~tB�I	a v��u#G�R��� �1P�xB�J�V���-�th��k0�LB�	P�Ѡvn3l�K��-�LB�/hr2�{�m(h.s�Ɛ�tC�i��`����!�@�A���5"O" �@�EWp�l�bOҢ>a ""O�-BB���_:Ȕr�AZ�j�yu"O@���
v�^$�@�Ĥ$�̝"�"OEYbl8'$f=��o<'�E!�"O�Ey'�ȍa-D ۄ.�|]��"O��pO�hW���w�,_�v�"O����͟?Z`�u�A�}ْ�"#"Ox=�"#�JU���`a�%>���"O�My0�)`E���Q ��n
&�8"OL��S#�`��H2���"Ox[6��m���qvI��,�܉#"O6!FA��k�l����XD�"O%��e/w�jWiЕ|`ۣ"O��1#^����YW�I�|G��"O���3�J���r#�,M�P�B"O*廃�#!�Uz2�3D/���yҋ@�7��4@���R��� �aͪ�y2J�7�0;�%ױF&!8�kP��y�o�%[�dxq���pj�:É��y2"߭;&6��N�1��RCD ��y
�  ��b�}������C��|�ȓ�� �bF�$�=�ҠF�+,V���f��(�䎙�7ڞ��ŧ�5n���K�P9F�.��X*dfϳ7�����<��7X�����nA�"�Jl�ȓ-��u���R�Hհ1�%-P�kT�i��$�0b�����`����P�5�4��-���%闥\�Iq���`��!��-=Ȕ0�)�'A��W��A�ȓ#?$I �`_3zk*�p���C2А��,�p���#�7R&-�PPFju��Y`���`ǈY|$�r��җ
2�ȓj:e3@О4|���9�:%��4�*U��C�7�)�f�+۾�ȓ�BU�Gf@��%�zg:i��C:D��a��P�A9�!p� �QI`8@��"D���Ę�7�!�Nr���Cԍ;D��	%WxE��ŋ*:ޒ��i;D��@��W�8�8I0�i׌\5jiYn9D��� %` �bd$@2Bs4;�g7D��K�ֶc\"�P ݳ4��U�)2D�4����1T��Y��AY�M�V��`)<D�D!�eH;~���"eוl�(h�5D?D���e�"`4�|�U��B ZMJ��;D���C˗�h[J��t�CW��thӠC�	j��Pؤ���B�FT�U���8��C�ɀU�(=r�i
�	M&�@�J�'��B�iI�V���zZ����
=7��}�7"O��{�n��u$�7��}��{�"Od�a�KTF)� ÿ1�h���"OnpH�h=5�<-��8Bu0�"O��cO�w��H�c (<� ��'W�I��H8g���4@sE���J �B��+7�NU C��,aG��B�I�d�Bͫd�4x�h�'Y+A��B�	�	��chO�vV�e�QaU�gN`C��t���K�\i^Ĺ�N�i�rC�I$2���C�ʁJ�y�Q�ܿM�V#<��y<�z �E*h)�a0#B3wu����A5b�b!a�4�h �V�
�4ȆȓT�H��������C<%�ȓ83f4�P�ʰc�H�Ij�
�Рm�L�����V�Ld�Jĺ�JP�$�� *B)�y�n�6��eX~�H��H��yrl��F�)�g��*a82�d�yүX)ao�U�VI!~k�ly�O��y�G׀q�,E)�`�fa
�nơ�y��s�&M��i�2R~
(�1�צ�yB�ڂv��aj���0��#����'xў�O��};�#A6-,�(�E�,0��'Ff�
��Ҥj� �%��,����'�Ȃ���.��T�R��v݂h	�'&�@6'�P�bU��`�R��K�<q1O�16응��h$����F�<�T
��n���!�2t�(��u�RA�<	��u��5샰��I��f�<���38&��sB�.,���i��a�<��F̨*��C�.or�KC��C�<��),�,Թ�"�' w�9��A�<f��7g�=v$��J��0��{�<ѱ�̋7�R`��K�70y&(��q�<)�.K� \, ѓ�-*Qn����S�<�Tl��y!�h��ӧ[U�� ER�<	0��E���"�M�'\-P�	�P�<� �D�!k�4
�Lp���+� "OP(�g.��3�D0Yի��wE��P"O8	r��?}�lͨaj
'�!I"O��G&�2]�!j�"��d���P�"O∉ba��rf<
��K$@�H۴"OxUQ�NN�2 r��E�Y���`�>�
���*V��j�sQ�E'���ȓ �L���":l��و��'��هȓl�ı��l�1��ѫ%����ȓCY���u��)�&e��
��=��1�� ]��F��)i@�`��8�ji�ȓBZex�KE70�lg)�i� Շ�j��;�$C�"�F0sMO�pO����%��U�t�>{�  㰧���<=�ȓXJ���I�8P^�u��j-H�ȓPĤD�3�J!3��XA��'��ȓ&�Y�s��r6�y��$mNbą�-�$[���(:"^��'��� $T,��a�"���B:a�ҍ�v(ɹx&\�ExB�)�n��i�<PW*Rq� �i҅^�<q���Z��u��
H	��9��
P�<���D�g��-��i��c'e�I�<����9\@8���Т6�69�tD�<�2�Fg�	9gM��t�[��ID�<Y��Ф:��oB�q�C�k�<铩�Qv�9Z�oM�vaJDQ�\s�<�C*��I����T�WM*�:U$�E�<�!'	��!c#vP�JJ I�<9G���$��@QG�F)]��R��K�<�Gn��o��qҌ׀w�~u��j�Q�<)7�
5�*@R<.�
�-���x�C�F�����Ғt��0�^����hOq������sJ.���T�]i��s!"O��Y���@i0��GnŢ+Pn���"O0���Ꮇw��t8t���?�.�;�"O���F囙D�j�{�~��"O��i� ¢�6X��,3q
���"O�L3Tb�.ۼlJ�K[]W���2��؄�	4OBʀʢk�@�����B2<C�ɻb��c"!^�zQMk#�J-$C�	�)�ՠ��(����cSb�bC�I�N��Dcw�C����z�OD~VC�I5~!K�)�~+�첇E=L/��D=�S�O�T�+F֡FBpBw�"|����"O|5��Ù4g���%I_33
Q
"Ol�)�@�BFp|�f�dZl%3�"O |ñ'�:H��pk��8�p���"Ohr�I$7�2��eً+I�Ū�"Op����PH�7.A�̚�"OT���u��#�m� {�"O��(�@�eR�qmѲ!U���A"O�9���7�f���A��S��uJD"Or �U��1!r�����
4�Iy�0O���N�z�jt�W ��1���Q�!�E8�Q�kP�DB%3.�=�!��K�1PP<k��9.?���6L$��pD����{��iD䄔*[Z N���yON�5d̑5�
ROV�i&����y"�ЙPɤ�z���?4dTLQ���;�y"@:dr��3�@��w9"d됫@��y���u�l2R�L)���+�y��#��g-]�;.��K����3�O^�5��%$Z��:�e?�p"Oj���W4?�%!�kW��(��'Iў"~	� Hq���+KN ��(0���	"O@Ę�����|��I	�}֢�*V"OH�x�W:|��e�
��^�)�"O�آ«�e��9�'�֋����"Or��@�,h�~D���n/
��B"OX̣��"u̮=�U��S4^	R�"Oj� � rR�.��GT���"O­ �!M;d�|kE�޸Aء���	c�OG�qi�*�c~�B�G	����'.�X��`Op��=s��T3�.<c�'k�՘�kƇg�F�Hr�J�I��Lh�'\�mJq&[/��@1e�xp֘��'H蔈�'1W^:0/�<�� ��'	�T���
IP�Bo��7��a�'�����Q�lX"G��4�SL<Y�����3�1Y�Ǉ�i%�=�NY��rG�N؟(�EK�8T�}���n`�!���3\OD� &H5�K,W���:�,@�n`c�j�xv!��g_�و#���Cw(|;�H�2�qOLIʏ������j�ťҳ��]:�e��y�T5P<���йu�������ybkܫYH-aQ�]�p�>l� �-�yR끇a�B- b��pf��W,J��y�Q�KE*�Cd+è|~$ J�[��y��3R����3�ݞx�h��E)�y�*T�ƥ�Ն��l�&\ف&��yd��Z[�y� �P�7E�I�����y��P�U#@ダ����=q����yb⚎}s��E��#�(��=�y�����s��>�n)����y2F� ޢ];CU5�prP
(�y�f�``✁��J�����ဏ�y"$E�6�9�DD!�p!A�
&�yR��
�<��,\  &~q�����yR'֞q)����#�p�pLBH��y�D��]���a�ǌ�s�hs1�S/�yB�A%P�8]c�*�1́9�ʝ�y�C�,�)�`K�~�\�2AIA��y"�
8�hQ����*�����y�M�X���vlY��(9����y⬛�8�K j�Zk��96,S��y⭉���(B�bR�N cB�Ü�y��wN`�1B�:yB��y��E'r��RSL�7���ϛ��y����P�G	�-���*�!��yrD1B���l�4-¾��6L@��y���G-�a�"�? ."��F�Ã�y�G��d�2EI�I)2�X�u����y2���� 12��5z$n���*�y��<9D�U�F��D��l�$����y�e%2�XL��FA*>x�}S�e�.�y�
�=�J��7�R�J����`I��yb��c9�[d/�=B�+en��y���4��|JT`�7;������Z��y"��+�т�/4ĸiYd-W��yAT�}����4���)@��J��y"�nP���LZ�8{��@�<�y",��tl����.�#���E���y�CO�C�I�¿H�.�u#�?�y��W_�qH��Q<*El<U���yr�ZjF�*"�N�1�|�%�K�y�M��IԊ�����!x^liJ,�y��T.i�XU8p��$l$(At���y�ˀ�g��-���^�d�
�j�,̈�y
� (���/V5^v��� .ڄ �����"O�i����f���X�M�3��+U"Ov�3��&
��P�d-"B�p9�G"O���1(��F�-�+_� �Tz"O ��E��_�����)��H�Z�"r"O0�ᗉ>���1"͚u�b�7"O�$��ك2p`@z!A��8%��"O�T����K��H��T�T��"OT�����~:T��Nբ/[	r"O��6�B�IB�N�lR�X�#"Ofѱ������� ��,mD"�Rt"Ols��F,L�(;����3���w"O���Td�4�`	o�!M��y�"O���u!]�`:��� �3�~ 
C"OD�� �ש4w��aWm�7��k"OH���ͳ#�4%�gLc�X��"O�LW!E	�YE�=�~�@�"O|���j#
���is���\�8�ps"OV�K�$�&#���0Ȗ�Eh,�c"O�a��o�al4�C��Sb<��"O�������L�i�Q�͌;w����"Ov(�BN���r4��3^��� "OȀ"T�ɨq]�e�A%�y>
��Q"O���s�Χ ��5�Uc�!:����"O�h��ALV�4�KB���g���+�"OBTSg��bCdA��_�"eɧ"O�l$f�$�6i�F7#�F��T"Oȫ�ҢKL@|�A5V�|`:e"O�	�� �'J�9�l�)B�%��"OJ�ٔ�J�(�6승V�<��"O�(P O4{x�0�*3S#>�rT"O�AB0�07��L��I5*-��s"O⸩���Y|��P�C8T��R"OeB�>8M��j'���(����"O|-z�I�pP��8���?����"O������J�(���AOF��$"O4C�( �fQD��4��{��T�%"O�1���T@��@�3�f�zc"O��is�҆)�(I�]�Qqe�"OZ���hѹ,�>A�"��2U�9��"O�IѰ�E� �X��%o")��"O<{FÁ�o[��G��]�Q��"O��Z��U��=� �*#��9�"Ot��W��,d���Ex��(�"O�u���'�:��f#J�bt��"OF�� �S�R�84җ�H}R�y�"O(�
;=�r�b�`=�p���"O�])F�(`8>m#��Ϋ4�⡻C"O��� �I8��\��0�� "OZ�`W�	�Is�h�jć!1@�{�"O��bl��-�BT�B/%&��0"O�q�J���h���-橢�"O�����?2z���J�zE�*q"OP�hE9
=6P�t�)��ŋ�"Oh%*��l߲,g��	@v��H�"O�Pۣ��am��.d0��"O�����HN�fш�g��,��D["O$ԒRJЌ
�&�9%h�*���r"O�8�sK�|���gFI;=�"O�� L�+�H%S���S`lyІ"Ovܒ��G�S2�lXU��I1�{"O$t��eȐ"�`��*[h.l	z"Ox��fEb�x�+㊑$�$%�a"O~���J�~njA��>u���0R"O� ��͋�3�x�" ����r"O��B�>�Lk� L�6���C"O�]j�@�q$��#��=~��(A�"OpX#��\�clz��FiΊ5F��R"Olᱢ�X�E^�X`��96��R"O�(��-�)YI.�8��S/. �"O �����N=ΐ�«��`�����"O��
1̃v�$� �,��Ub""O�HU�@�^r虱�G�,�Dӡ"OTI�@�
~H�y�A��&ţ�"O̔���Y+
�� ��;��tzD"O�e�f�;I(��o�"x��i�"Oh�A����J��&"�4�zF"Op4hh�*vK���G� �h����"ONH"qhD�[
lxQ���m�f@��"Oj�i���w�����c���"Ox�Hf�Q�`0� Iw�,�V"O�ԈT�J�[��T�Hԥw^*ݘ"Ot�k�\:4�U'�[>Q�d"O���F&0B5
f&)m��"Ot��7L?!���ԅ
�8��"O���b�=� =�F��y��I��"Of��Y3�i���4	�����"O�"@S�q5R���\k��"O@h�r�*)�$����y��"O,�aE�	�}�T�� Ԅt�x���"O��R��V93l��W*X>3$zȈD"OFQ�c��hvHX�Zr̒�"O�mZϋ�tB�a%f�(>h$��R"O\ؚW��@.Hj%vs`ԑ�"O�����m�$�� ^�`� "O�3�AX��1�J]�o�&m��"O>��qkA�V�����U;l�L�"Oh�Я�?�,�!&	JLX�!�"O�*!�4f�,!�@��X0��#�"O���!D4d��e��W0 Q!"O�����(3P|�caTP"����"Or)�GP�^�5r���
����"O�=N�J� Qӓ�ڒ�R��t"OLӑ�:c��Ċͼ���"O��R�$*�Ku��Y>�s�"O5Z��'&N��&�x%4	@"O�Ђ��&4T��䗞��B�"O�zg60֦<q��phS"O�9S��>4�X�VTUJ0"O���0�=sF�CQ,)$^��@D"ODxI%��?ޠA��
U�Hx�*"O�p ���_��Ps���%Wvx�Q"O��xuC��+�|��B_;DgP|C�"O�Z��«[��%�%⊲U�X��c"O�%��I���E0(�L�6�� "O89s$�Xk�Tr�� g��I#�"O�uK� ��('y�\2of�E�W"O�S6���Xުݘ�#��J]8���"OT��)O5xJ���DZ�T
�+�"Ovy���kwr}#�!��02�p��"Ob���-2z;�M�5`�+Uy"O�J��*�`�sR�ٶeBșa"O�$ID-U�ll�Xàj��N9E�""O6M*ƯC�*�PA��I�.�p"Ol�0uH�y���J��X�O�ʌ��"OmF�Ѯxx��U*U��� �"O�K���$4�XZ�
�R�X��"O��`�E�-H���U
]&P�d"O� $(b-��?e�=�'�W�Z"�r!"O�=P�BLC��A$��S���Q"O��Yb��O�͈s�_0Ʊ�7"O�|R��ڔ� ����9w�`��"Ot�p��@��<˵a�~�0�Ȓ"O�2��O���rៀ	{^䠕"O`����\G�@�B���|�l���"OX��5g�d��o�8dv�u�v"O8����+�m�d�@��y�"O����FY�H������H�ܩ�"O<U���K��4���bK+|h�}�'"O����G/=��q���i)�(b�"OD5���ăF�A;��
�6%>}��"O�
�GE�k�Yh�lƍ"(�v"O�a��M�ec���Q<<V0l��"O�hVn�0�B���J/5:| �"Oh% ���S�¹Q,K��y҆ 9>�0k�z��1����yRE�@�.�9��Ҏ._X�Z7K�"�y2I��F���8��4%�*H�6H��yB��yҚ�Rw�^�!"�(� .��yBዌ*�Yy�nwa���y7�QC�'�\����<�(����A�� C�'96���F��Z�6�ig��S�4�	�'��J��#4���f�@�y@���
�'��8�惡'*䀺�F}H$$�	�'`�MP��D��iz�)S u��-i
�''a0��G�mꄰ��i҈i���	�'<D�pT �2HnP�Zc%*a�����'ԉ�F'�$��	ѮghМ	�'�KB,]��y�.�C&�s"��C�<��χf� %�dJJd&���~�<���Ι:���*R	s��)���|�<�A�ݹ~Pfب��^����i|�<�Ќ�=A�z�;d�=%���"'�m�<�!!�
@���
S-A�1�éA�<�a�RB5|����|H\��E��<�kE�	=�t9�A@2�t��Q�]{�<A^��ع���-b�p�	� z�<١���?��� .��e-(����t�<A#�V�IҀ��W�D�j�]�!Bp�<�M.s@jb��v0f��Ddk�<)�+	D�d��ԡѮe���z�	�`�<)�'U=#��Â?M�%I"�\�<!��f��j��C!{}#�AV�<����X+Hò�Ӗ\��	;�e�w�<qƋ�A��Id!�B�xQrm�u�<Q�_K�HeQ։�:z��T��(�p�<A@A+W�9!����c��A)Mx�<a B�Qټ����"�`�hEs�<��l�o1:|K�%��?{����S�<�v�͆r��a����!L�X�MR�<� �6m3n,c��&" ��� h�<a��|�P ���	2�ӀhQc�<�G	�Wr$����.��iK��w�<�U�[  ��X�Á�{P�-�c��t�<�Ua��.����`�*|��U�u�<)R͏&Y�֕8�)�8��X��.r�<���Y=DҾ�B2��PJB��G�<a��Nm�
��JΆ	��t�ԍ�i�<1Ĉ��B�Hm���P`��� u"�g�<�q��:qa�c�.ψ&��+�*}�<�w�J�& X�f�bݨ����Px�<�S,ԿI*6�3G�'e6}s���K�<� �9� ��̅ &�Q�k�N=ɤ"O����#��X�"|�箓j�t���"OB d�V��8�$�ss���"O��UDW��1�b��ccr�"O<}"Ċ�`�C��P:Px�+�"O���ׇO�,�@��J՘<Y�"OlQ��H�kI���âWV���k�"O�	3��A�x�4��&�M�����"O���%�(]n��뗛��))R"O�y{q�p_$���j,^uXڃ"O
��B��)kT��sd
3^Ϻ��V"OJ��m	����t��KZ`�"O���F���Ov�`I�G#8;�Y� "O�e�EG�1�9Q��b0bx�C"O "����
MZ���&^ �"O���B���A��]�D*�U T"O�A��a
,1@�Z` �%!ڌT"O"X�B*^��A��{-b!y�"O���D�\�n��<X���e4,�"O��ȵ"�>A���S�	��r�>��g"O�d�D.*!�jx[�.-8�4��"O�͠�A�Je����Q1v���9�"OL@9�Jѕ6��bv�^�%D���"O
�xT(R��i��F?\��9�"O���"4��<B��)jԽʔ"OrX`�lرBMH�s�o^�5_���"O:�i�#��>��I!�X�J?�٨"O�D�Fe�%$H�GLT�9 r�r�"O��	�aXh��P$b�?�X��"O��၄�0yp��d�K � ��"OشyF���_�B$���<�X�"Oj��c����-Y%�C�uטL�F"O�1b�DΑm�9s��=Ɔ��"OJ�sL�QJ���gᙴ�~�h�"O�׌Ηcm�`�b�Qn�L���"Ox\�I���T���^)S΀0�"O�����)g���P���9H�D���"O�ȂL�8@��T�ݴ�b�K�"O�X�f�l]ԭ��E�pԜCs"O� �b&�Z'��ψU��B4"O��RcC1c�@Jg螡2>'"O�,T*>ta���Q�sA,]��"O0���M/�|P�	E�46`��"O�) �ʑXN0)��)>	1f4ӗ"O����W>w�@���G�3-��H"O�]c�N��)!�AB�g��2&��f"O�hC'ȅ�fW �I�F%�9�u"O5�u�-�V�{G�KB��	�"O�u����]\<����ӏ�4[�"O���A��v��K^֊Q�"O��+Џ�C�Vq�՗73"�XC"O�mY���ic�A	;LN�p"O�-���v�j��#*�"O�pӯ�g,
8���?A�m�"Ob8Q��B@�\X��?)�lA��"O��avhZ�d/pE�G�Ӊ)}�x�v"O��� ��z�@��Ɍ|FDj@"On}��z�%ƞw�	� �;�!�$ɇ(����ܮIj�7M�;n�!���5%�]#ISx ,t�c�X�>^!�d�T
�#Re�`�lQ4JŪBJ!�$;���0�$�/��a��
!�D�p�y�d�5T� �ԏc5!򄗚�hp�6l !"�1ȠcE!�� $�;�A�#M- �G�)�H�PC"O4��R���!t�i�s��5�0�"O�u�Fj��e�^��6��[g,J�"O����D97(��V��zgĐ�"O�\"�ǚ+C{�=a3cC T�<���"Oи��,�+����rçS�:8��"O�M���ۈI{ի'j�$3f40�5"O�%�3d�<�����"J�)�"O6�"�E�R���d̮+@v]�7"O�	2�%������U蚋9�\"Oʹ(c��1���sa��#�t�6"O�dA  �5G��I� ��J�"O�Y���䨐V�Ç=�2"O��u�5E������B����"O&��$��m�ZHb�a ^�v�"O��O�1�B�6���SS>�T"OnA0�E˾��x���#"O,T���Q����۠.Q1/<~�2"O���u�L/?���� �*D%9"O4�B��:lv��'�؈\��!"O�8p��	��:F��%�Ĵ8#"O�Ӈ��/�0�1s��D�ʌ�"O0�M�"�����M����9w"O@
� !!s�p"�g����e�"O��R��Z�I.�yR�֥ ���"O�8-��L�(<9⃍��Es"OtTr��:|v \p�C���mHT"O ��e��)*�P���� �"��"OB�kq�M�y0�%%�Bi�,�"O�TR!��$~�n�X4d�xO|BP"Otݛ�.B�Iy�u)�B�D[
a�7"O䝱���%ikVY!���kE�-�"O�2e�Y��4�R���B*U��"O�	��`��@�Qqj��՛�"O(p�4N�x 5�!fF7i�n���"O����?8��E(~{&e!�"O����ET:=v%�u�^ �6x"G"Oډ 1�K�D���  oѐq��"O��7�̪:� �QG�����c�"On�R	,����u/�7G�@�"O�F�-{�PP��{�^���"OR��p#ɘp\�`
�d���6I`"O�Ƀ��гRDH�/�vLZA"Oh,���?X�\�#� �����"O����Ú�+`Qy�ڰ�"�x"O��Q3�A�9�^,Bp��>���؇"OJ�	�j�9(��(���V�\ �lá"O"�`���:9�x���k�9
"O�P�a��"u�%!�L_�k�Έ)�"O�R��I#S�T�����D"O��!��FҸ��
s���v"O, ��NS5tɈ�Ceo	�����"O�	�! :Z� �薟p�3"O�`j��!v+41���#˺�Xf"O�m��J'Ae��� D%��CQ"O�8�
�y��a"u*K3D}l�36"Oj���H_�0Fb<"��9$`|�ض"Ox4p`"݄o�5;��×Y%��P�"Oj��!ܮo�i{D�%K���C"O���Yi������ێ6ܣ�"OJᅒbς���Y��&`@�"Ox1B�B\�Q��c�h<A�T��"O����Ύ�6%�G�ŧ_ �LYq"O�Ȑh?T�0]�"B�j!J��"O� 5�q��i `i1��Z�&"T	T"Ohl)�� ET訁�I�"5"O�p��w=��1��xb�Hp"O�L7MR0*TX� �i�?S�V��"O�!�aL�]+�Y����m�j�S"OB���Sz��+�.�R-#7"O��)7�W�d��{v�Q-6"@�"O��j(�]��)�M�R|!y�"O��	QE:`��}"'��\t s"O��&�T?<�~mKC�\�"�y"O���� `��Ԋ���t|0a"O��s��ڵmMp��EFq�5;�"ON%ҖC�;J���3B��1\mv��"O����kI�&��0c'֦gN��""O �{��O�]��P �&ݟ~?�i�"O4�@�Z4���&U�((x�7"O������5q$X�A�̡:"�}0"O�օ�F�h��J3C�ri+�"Op!��I������Q0"O�ݹ��?ڦ�p�D��Q�
8	�"O$�p6�Uْ���R�z,��L%�y2+�nt�#%��Gaj��ƌ �ybKJ�WH�{ѧ�6F]�Az�d��y����	��:����lZ%�y�DU?"8R1!Qc�`{�G%�yrBQ+fbN���'��T�n��_&�y��
#m�6/V6���a4�yrĆM2�I
̱K�Т�!��y&�Pq��ht.
�pT#�B�*�y�0c�z8��%H<?����aϭ�y2�64Hk5�ɩ=2x�n��y��a�`2�O�9^�xJ�D�	�yr�Ϸnp=Z!c�/Z4�0{����ybj�K�F�ä�DZ�&��RiO&�y�(��Y�y�sJ��Kx�e�H��y�ƒJ�z�JE8E�~����?�y�.GW�1 G枱n�([G���y�D�t�*�`b��g���d^)�yB�@�P'ШT)ֲd9\������yl�[�f�͝�	iP��!���y�T�.��i�d˝�r���0έ�y�V�@7�u��)Z&d��T�p_�y��O7�v�GiC	I厡+�c�yb�#>`,�FGٮ<BN������y�AĸX)��]�K<e�S�C&�y�!��H�YJu�(��uX4�]��yb�J4-��!����;*��Q{Ӎ��yB*E�$8,
7OR������"�y�)��A۳w��z����y��Yan��͕�t�j�@��y�����(��� ���P�@���y���Z&@�b�f��ր��,V�y���/�N��Ѣ@��zȺa��y�ցc �jQ(|J���p�3�y��N�C���描?�"���f�y�H�h��&G�9�$B��W�y�c�<-��Q�$�L&_?,�P@(U��y�C@-*�1�BR�� �����y�(Z/�T`V�L= �^��ƍ��y2lȚJ���r��1' �x`��\��y"��!"�fH+qH\�n�|yaQ�	��yҊKWuBQ���	m�a0΃�yb�T#ʺ �� ��_�L)(�@I��y�+U�`l���K ��!�G�S�y
� ��"7@�>/�!!�B�I��Pa"O��*��
D�����Wl�!"Od(��D٠P�ޔ�o.?-0��!"OMȣ̃	/��yD�E�{(��("O ���j�1t��g�P�^$̕��"O���3�@LÀ�k�g��j��v"O���V�e$�Y"�-��z%i�"O:p�!Զz������3��e�u"ORsD�QR�	�d���`i�"O�G��3p�]���͚�XA"Of��H�5#��m��]�����'�Ԝ �](�l��.ƈQ:^�1�'��j��B%
���0��^�ԍ�
�'���1���?��q۰ȅ GlN��	�'��tB��LY�fȳu{�x��'������L<���i�M=k�����'?H髕��(rf*`e���:�v\��'IP�o��g-J�Y�795"���'����RL��y�-й6�Vh��'i�8�P87�!�fnȮ=z���'��}qR
�<Z-Z&Β:e" �h�'a������\~��"l�f�x���'R^�@�X�x�B�5I�6�1�'B(��!ʬC�2,�I/#��M��'�jț�U�	��h0���m�Qa�'�D��.J5IDT�� J%d���'ƬuB/�	N�P	�w�\.�|z�'t]�� ��N�F��6��}�<�x�'|�Ěf� K.��w�>C�X��
�'R�� �O[St��G/8?k�
�'�9��*J�\�|䱆ۿfƮ���'L0�ӳ7 d|�E/���Y	�'d���F� 1@A��T-i�'���(��E�~����&�fm1�'Y�r�k��Y�$T�R���J��'��TRMS�V,�+㏨=R!`�'/^�Z�l��u�*��u���7�eq�'D5W+֘�������-��q�'��I��
���f
�""p|h�'Yp9p%�/l�2�����XD`Y�'g��j���4{�@����Ml�	�'�������{2f��a�
��$��'�j��!�+F�0��(ǡe�I�'��(��P(ĪEq�KKo� ��'m�P[�����7�Z�:b0�'O�d l�OT&Qq�N#1����'#��1�(�=iLI`J̌+:���'E�ᰶ�Κ\p^x��T��D1�'F���%H�!h�!�RF �`�'�V�:�O@�5H}���I�� ��'��%��%��c6�;Qu�<�'t8�����s��0S( '��\z�'�D�v/�.��8z�O�MHx�'I���IY��ل� Rv����'K��3T�gUؠ⣌P�J�
�i�'w,y֦0 q�p���H�|I�	�'*
��w�|'|!+ѥ�6C/�4�	�'��<81(ǆ0������
=0�AB	�'J�$�ь��<8����O0�i�'Pd�׌�?}U �1r�9<),m�ȓ?¾t:�\�\�:q����)C]4e�ȓC`��Q�Γ1&��s��&X����ȓ:m����g�:�(������	�ȓS��9��ϓ[�<u�ѪMgx�<��S�? �u[�O؟FTF��F��>z^R�S�"O��QL�7�"[O��J\��"O�����b?��2�(��S�"O���vEǸb��x;��Tk��i�"O��!�A</"����%�h�2"O� x�%��&��H��ė~ҹ+�"OJa�Hێ�z5�A	u*�Ӕ"O����{�L��m�����"O5	��^�O{H�B)���J��4"O|)�C����(YU���Ll,K�"O4���㏌.�"HSE*QL�P�3"Ot�Q�J�P�P$)�.[�ڰ�b3"O���@ 'C"�8��řf��A��"O^��5n߯d&& ²CS ���r"O(�@1Hʭ�	��B E�@ӵ"O��Ѝε|�Bu�AY�obH��'�֔	��E��j�n\#՞t��'>�����L8y��)�+	�T�ʓ3_H��Vl����׌�^�8��x:P%�͗d�j๗h��H��l��%��	�l��%W��ѡ/�*1����WL��P�V�R4��K��
l�ȓ$��x"W ,f^ zW�Il̮<��D�NQ�5.�35�e��z�Lцȓİ��1�d$�Âߏ	�p��ȓO%l8Qa�#n�hɻg�ލ�^u��O:���U-�NL�<����)@����tɂ�CW)�OQ�Ӕ��ȓ�\�u��(cH:��W$Y�?�M�ȓ$h�I��e����e]�t�rx�ȓz��Y
�(��Honqɖo��$�ȓz����$K�;7�`a���& :5�ȓ��4����(<�\)���${V}�ȓcń��LAU��-��)�E��؅ȓp���aƭ��F�L���&O�,��ȓo�Vq�����N"@����4�ȓM�.0+`	��w����K�����ȓL<��G/f�c�H�R��ȓVVl���)U�`���#Y��ȓh��c�Z:nO 8���6� ��ȓM�b᱒�5�l� ��r���ȓ�d�JB�N�U��,B�	zd��t��PX��p	�L� ���d�L���L�`���e�h����rfƱM�����c��Ұ� )D1�[��`��ȓ]&@)t(Ʊ2�*�e��Ȅȓkl��Z�iR�?��<;P�|�n��ȓ/,���	O\��"'eL=@��ȓ5�P}btbJ�,P�b�K�Z���ȓH�lȑb�K�b\��#	V@���sf�4'��^~B��Gڽ. �%��-Az(@j+�j�G��gUb���L�ڽ�&&��|��9I	E��N�������K��V^$e�L#@X��t�Q��IX�l�: ��p}z��;�	(��\���!�G3�a�ȓ]Jș�M,,�Mr���Қ<��76�`��]�!�,
K�T��ȓh�\��$����i�^�<_V��	d��$I��c��9F`ӱ]�y��eHQ2�M�����c�̙�4�>���!s���et��X#j�%��̇�]�݊��Ǚz���p�c�:}���R��,�萈�s+�5��S�? Ұi�G5F[�� L(�ɱt"Ol�p���^b�h茮#ء0"O�e�r�ې4s�T�@e�j-<0W"O"�4嗢B��y"B��$hUB"O2M�m��a~�4����4A#�c�"O�虧@M�hEз�H"�"Oub�D�A�8�I�fF�Nh}8T"OzP�6g�
�t���;K�~9�"O�uk�J$`�e�C$)& �"O��s%]	\|m�!�ԷS��(	�"OF-���\�d�!#���qS#"O*!{Q�G�����C��6a��dy�"O�5慄#$έXR�N������"O a"�އz�r+��{��]�u"Ox�Dǈ�O��ڇ�R�QR�*6"Opm��3S�"�1 �
�D��"O�qk�@��"�E�B�� �dP��"O,�[��9ox�� �\H�~�)'"O���AY�eGTĳ�G@ �"O�);�)˲Z��谔/P,2����0LOZ�#ӍE6t�y`�͇T!а0E"O�Qb�'0Z�Q��O�&��aq"O��yC.�rH�q�C�8��@�a"OfD�"�K�u�y�Ս #A��$�"O.��t�|l���wB�.��e�"O��x3��F���
�AY�c��y!'"O�t	Ө�?U�r,��/�N֌�z��':ў"~j�H_/e^A���~!�Z���<�y���:n�xݱT΀*T6�����yb�+,�A"���)��0!bcC��y�J�v��
��8E��*O��yr�D�Zz���DA
��<�����-�y"�Y�a�ͫ2�L�xU��S�(�y��%%O�1"'�uۚ���e^5�yb��=s�fm�A�	@�Hp�����yB�K��&�;#�#P>U�4�B|��np4gǜ>M�\�H���?آ���h_�`t�4h�$|h� U�ń�A36��V��^���@�M�i�I��D�4SeG§8����m�pFꉅȓ-��`�t�#4l��î��}39�ȓC�Lժ҅I�k�z-���5<zP ��Aݾ�q�C���q�v��1�6��ȓ{xZ�@vl�=�))h
|����ȓ�B�Q�
��yZ�-\c�E��]�Bd��l@7��¦�טN!%��N(nl�T�2]����X�BMLl�ȓ�`��O�sy`���jн`�vŅ��
8�AGج�X��A�L���	�ȓ7c(�2���Չ@�؈�v�]f�<a�a[�Y�T�"kQ�mL�m���GK�<Ԏ8X m�7۠R��eiG.�K�<�i6p|������*�N��L�F�<��ꉄT�^|
� U� %�t���L�<�3�.�eIBX�_��� U���<�oH''��@�@E;���1��G�<���" ��yCiJr��׫�|yb�)ʧL�h��ǠU"���iQ�N� �p�ȓobԤ%���Ev���ځM�D�ȓtJ�Hs�G�Uf�M� 8x��ȓ�^LR���u���A7���ȓ*��L���c:�t�Ei	)p�.Y�ȓ/2�a���e�$��f�)j� ��^ƜL�6�֧���!�@?O��)�'�ў�|� �s�%�!r���'�Z�/�*I#�"O��Cb)޷n���3��$s�څC�"O������
}dx`�5��?�hR"O�l��A�6<��)94&�Q��5�G"O��K2�
q�&#�O�L��a��"O~�b�LA�v��!j-����a"O��!l���0�T�Pp�g�'}ў"~bE
Q��`���3T���&��hOh��O�q.ܑ)k�z*^����!��/g�F���!@9�Kһg��8Z�'�Nd1q�Ӆ�D���*d�0�Y�'ru�튂y��I�ͦW�q��'�����5Q�H� !N�Sz)��',4����S�Έ� ��Lx��:�'�l9�6.�|�@��ુ^�-��'� Y�4�_ ��pP��8H�f� �'����F� NhT���Br���'z�,�w���/����������]�L4�U��#ʘ�P	%�~͆�5&�if�M*�t���:X �ȓ|��M��Q��EζМ�%��D{���ȪM<6�P�쏛V; ��6�?!���'0��k��N�2��hz�o��֠��'cH�!�K�Z𨋴(M<����	�'j�k��N#/�^l8t�E?xk쀀	�'���,L��<�4oE�r4�L(	�'�܌ptlUSv�֎݈S�B͢�'r��	���<C3f�ж�O�bшH>y���iF�n[����6X�x ��)Y�Pg!��K�b�Q��F؃�)�DL�K!�D��-��)jC��$L�F-Ҡ@��2a!�ZLn�`B ��D+�� ��<=!�$èq�8�Zp��v%M�A*!򤓋dG�a#ҀpHq��-S!�D�-6xt풜/���0(R���x��(����p�ːS�R�sh�T���j�"O�H����^U���U�Ҩ]o��9�"O���'Ȏ� �0l�0+tUpH"O����p�d*ݜldd���"O�9� ���2X|���<G��H�"O���v`� {p�����g��}+�"O��r.�����K��s梑�p�'�ў"~:'�x�q)r%
��K⚇�hO@���7i�()�[�J+n� H�6�!��5yT��`יJ@y��"�!򄚩l��٠��ިD:���CY!� )(�ڹ0j@`R\��L�_�!�$���I�6���($�GL (:!򄎖"FZ�"���	|d*���-9Q!�dJ�zX|��L�)��q�U D*1!�$> JJ��Re�.���� ļ
�!�d�*T� ��,,[�5k&Oώ-�!�dD>��M����[�4�yc�Ւ5�!�$�(s4�{Aa7��$a�!��Z�!�$�`�-����v��H2��ۚ6T!�䐯�����] }���mE�:!���0���6�M* ���P�Q\�!�7Gt�Q���c�D\Yn� �!�2"Z�t�S]&�vS��\�!�DY�`fb��e�>��j�	V2+!�$Ғ7�1�D:0����Y�e�!�$\kܨ��'�5l��e-Х=�!�d�!y*�-��>�^��F�)w!���XU.�Cnʅ�Й�����!�� �uPaJ�8\f�!;�͒r���q&"O���ꊧT�������<ի�"Oz4sfH�K��r�����Xi�"O0��B���[��L�f^�@��aS"O��pEY�aȌX��kz����"O���4��cD�D�q���"O�貔OL�@���ã��k�&�	"OX��ƫ_(`��\a��C�qۣ"O�@�qCI7��ua�̞�q�mz'"O�Ig���@z ��K 0	���U"O��S3G5%�|��
PT�}SQ"O����`J�T� 0C�g��|����"O���)��Lߘ�*c�V�)�"O:�1��a���[ ؍U)��6"O�V��4Qʅ�?M�|��Č�B�<�#�9r?J�N:6��r�lVd�<ap��.r<:c$��A?�p�A�Xv�<�%fV6v:J)WB��&%���Y�<�#����p%�K<G�U�]"�B�	�rB,A��,[9M��5��d8�B�[�(fȂ$O��i��x�p"OȰ��� p��3�V�(��!Q�"O��%A�B�yb��?��D�V"O�@�whD��P��Vi�����"O�,�6B��"�P���IK�}�@x��"O�QBWU*�� ��@j���C"O줪q'�4Y(M�4��8dy䝊�"O��{�d�s���+�$H==z�#3"O!��
H&R00=�A�$"n���"O.̲���!o�%�12Z±Ѐ"O���`�wT�a�3+S=?�<�h�"O�����\Բ�H�
jzb�G"O�I�S�_�h��Q� �ōM�����"O�ؘC�9Q��2����#��8Zt"OV�sF�]N)�x�G�<5�^!�"Ov���JSJuf�J���?�@��"O"P���:z!^)�T��,�}�f"O��5��
=��lQAŀ��@\�@"O�<�a�	�dӪH8.�I:�l)�"O�{��@ ��䁀�C�#3 Q��"O� Y%k�_�hDܛ1h�ʠ"O��{u T��x%	�![��ɒ "O�@H��r���M�$\�i`"O�-(���b!ڤAVχ�c�y@"ONH)3j�i�h	��K��K�����"Op���NƦ�(� ժ۴!���"Oؠ��CY4-l8���S=����1"O�`���ۜpl��j3��8��|k�"O�UQ�EH�%@��j6����"O���ܔ-H��f���J����"O`x�#m�	b̬�%�\�F5�"Ov���Lؼ�)��d�Q5"O쑑���ND�՚�F�:X`�x�7"O���e+�;~��EXV�;S_�X�b"OB��f�8���.AVJ1� �y�n܊l�̬�U/��z%�e[�B�2�y�ݢ�
J�'G�x��0��k>�y�;4����k�q"�RF(���y2
ɔY�H"�C�m@�t��ܕ�yR酖J�b���a�
a��b���y"�*Ax�ǥA�()k⪀��y2��8i,�r$Y�p�x����?�y�& ,�Y7,��Q���2�yr!�0i���㩚��jh��ꐘ�y
� �!�!b�/_��S��5!�6|�"O�P�c߽K���t��'�(<��"O�![��Y�M�"u(�L�4K�TM��"O܌���I;L0�13�E�&�z�"On��̕*GpU��ݢh�VШ"O\�5��0^,�|!���[��P�"O�x��T04��l�s�֥yd�f*O�@qq�-8H�+sBM1��UI�'�4�2���#��zGl�!!��mS�'�>�i��9wy�xW ��-����'�(#a�+3oF��Qc��
i�m��r�ӇN�#��ؖ��1X,݇�_.�Բ�l՜�ȁ����t��@��HaɅ;~� � �M8W��A��b�HA�f�ռ�����[
�8��g�u��ب+A��Ԧ0���ʓu�)c�'f�rf�B3W B�ɖ|�PͩC���A<*�gΈ�2B�	)hEDA�s�U93�����M%n��C�ɉ\��BU�ۃ���rB�	�XK�C�	�~}�҈�3* ���4�lC�;H�����;i�ҥnн��C�7l���i���<3�1�A���C�	�v�eY�KI�B1
8�� шu�LC䉵:d�8	u"��)��a�R�8�(C���\1�� B�21�#��nC�/Ma�hC*_e�28!��v��B�ɘ��Ȁĝ�v�ͫ�Q8B��B��" $̤9㣊�*��  �#�jB��!/�J�Y�+?.N�X{���3�TB�I�,2Lr`��<{Ԋ ��Hгu�B��5O��1.]�rQ<uP��Y�C�I��|�`��[ 2=x� ��G[pC��[��Ͳ�"ǀ:_�)#Y�:C�I:GF�ٹdj*ogF��Qj��\B�	�y��S��`6���=R_�B�I%@�ͩҧ�1y"�#r*�fA�C䉮�HY���G��&�P�*ǃE��B�I�w�h���ĳo>M��@	�z}�B�ɝ{hڍ\70E��cH�h`�B�$+�5s��|6I�4IF=�B�I?�"\@%�W�^0]haP�3,B�	�RD ��
7ms$q!3j��h�C�<s` ���Y�Oz�����#n5�C䉴U����6�ҋf�Q��`Q�i��C�	��|��c��m��9��w�C��#UCfq�q�:@��aql�)8�~C�ɑd
c0Ve��tS�1p.bC�I�mg�I���!&\A�J7s�B䉍f:�`Z�ܣa䑷�>h��B�	�l�,q1�!��Y%O�.aЦB�I2=����d�;Ġ�/'`�h	�'��K� dy�s$�l�h2�'�RsuB�#kf��#��N�	�'W2P#����z��1���L�y_�c�'4��1�	4hx*!����w�ڵ��'Mj��ׯN�,����㊃ p�i��'P�c��ڶ$C�jB8`�>)�'���J�_}�t�yq�Gh��X�'�ZX#�P�.����Ց)/f�!�'V8� g;H���î�Ԝ��'* �Y�)�O,������ȉ�'ub:�	O�I,2\���!
m����',�(ID)=p�"���jf��
��� f��cf 5u�~`pt�[�<]�@@�"O��R���$]�X�ˉ}[r��r"O��CA3�0�ѳ˜w>�tcE"O|������k�xD���:LP#"Ot��7i�1e"ްaE#Y�&^�+�"O��p(M�2�҆��<5��"OB1:�ց�\�S�A
0$T��D"OHT�Eu �9#���1L�P|�"Of(����KvVu�##�)�l�p�"O���U�jIp��Ă��[@-�"O΀Q�08��y�bU&�i��"O*d���,�B!lOf�4C�"O�x��%M�Uľ�Rb���\�*�5"Or@��!Q�\��HT�z� �!"O�؋�-��Y-b�bU�O&���"O����@�=蔨�ƙ�4ݒ�W"O���4c�0$���E�ͽ7ɴ��"O �JJ��|��ʨ$���r�"O�IK�+�"�t�X7Ҏ%��"O<����<�+� �M�<-a "OzTr����P�Q%� ivz�"O\,;B/H�=N�H�Q�O�S�"O�+P	W!<�-e J
~�"OxM��"F�@�e�f$ѼQ�^@�"O ��`�>r�,��Ae:z{Vt�a"O`��e��DE�dpO	&�ja�w"Oj���n�:?:͈���	IX��T"O��cW"CQ�T50�cƥO.Q� "O�a�kX�U(����Û��j`�"O��@�i?"��q�| S�ŅI�!�d��.��#�G�Kb��q�V�`"!�D�;[�,pi��E�]��5��dڨt�!��3�lJ�G��Uw�8����-h�!�	¦�� �V��0��(�6y�!�X8Nr5P`�ǃN���#5ǔ#QK!��?�ޡc�$�,����A��y�!򄆑t��-�0�¥Rpp�0pDÌ.�!�d���X9�B䊻nb��	C*�V0!��63���F�LI�{��1 !�D�*����Gjә0;ީ#g�[*!�d����@R"!�W>����Q�I�!�䟇i>6�Q�+ɂo�8�
@�O2F�!����h,��KJ�l�<Q#5�w]!��@��l�R-P
rOt�ۖ��'�!��)���Aēx`�IucI!�!�D
s3�kb�[�X�<�⡍V�!�ʭ#!<�s�ٲ�Ay&j�<!��ϓ[�5q���Bu:r���X1!�D�{t��@�Ek��@�b,h�!�d�[\��"rm^	=@�c�ڇP�!��2A���P���'.`�AGJ�L�axr�=���̓G�è&nI��5��u�ȓD8t�P�W;-�`u���G�nLΓ�?����i��v)n�@�� v�
` ��A�n�!�T�r��GĂ���)�5���K>�
�C�B]���>I2���C�Ij3�B�I����Ğq0��d�-K�`C��z2�K���
A���ᲃ��N�JC�	�T��B�)�0h���$��=�B�ɺQ��@�s�D3 �^� 2&����=!�'^�>��$�t8�WWp�傴��JY�B�I =m�,�"��*��UQe��h�rC䉛p�R���=E8l""�Nh��C�Y��Q�,	0wQR4x���԰B�)� H�����ci�������Jx�0�"O�q�`I��-e  A�ƀ���a�"O�a�'��t��Fn��v`91"O"�xA`��Y=vѹf*Tz� Aj�"Oz�u��\h��jcn�9�"OV��$����"5H4��S����"O��sg� cl$1��-�rS>Y���i��dD�=��� �Ņ�c�<cm!��'�qO�9��ʧ���R�ߦ}Z�<�F�'A!�� 	zN�4Yq�_;0�i;f���D)a{����(`��@-�,^c�y"LLS��XD�$ď2'9�@���'�q��ø'�N"=%?%�Ӭ|-4`P�OI�ZMa��ac�G{���Y�=�h �0dCG�it��C�>�'P���'�����&��6ӄE�7��9����.��{/t���m�w��d#�	@26@�d��4g=�J�6����_�[BE{�Mߨ�L��@Z�o"�|as��/��x`"O�����C&�q $�%2=l	�R<OТ=E�4���4�"��$���8���y�E�A�Q �+��"uZ�2�.�>�HO$��$�?0���r�/\�'>dA$�r !���V�8-�4��u$��s���!�D�xv0���Mت:<�x�)$�<�<	Ǔ5��mz����(��\%'�Նȓc��|JpC�%2$$���ɸy>v���NUJ�b'��3b8����0�Q��x̓w�PF��O������mf�E0Fj�QvD��NQE�'�џ�jc�P�
Sz���L��6�Q���'�jc��i�[�OJN�PR�{��	�����y��خAʵ�e�ҹm�6Yn�9��'�1O:�|R�&�*�J)��	5L$P����}�<A���+�T�Cd^�%���� E�~�b8�P��Q9,�����d�+�O��O|}��ɲ=Kg�ТN��['�x�'1R�A�u�` �'� Q��A��';Hm��S�_ .���d#`s0��'Y�	�gL+��PeGB�n�Յȓc�z�{u"^�PXQ�M+:�I��Ug���	^8��ä��(dX���_��q���8+Z� ��
���I}�'JfX�v���|M�f�C_2uʈ{r�'��)1c���H���P�+H<�����ԸiM��ʒ�@� �,�q��8u��j�'�� Pd`�V_D���(g�����'D���T�˫}�x!e�Ez����'�zT�p���Ov��a���8���+��D*�'ED�!A�S/�8�a��ob�����r`h�F}@��� �K�x��=Qۓ]}n!7��1}8=���[<0�<���M�v��)��<��O�F��q�Lp~�'�0)*uiX�2v�q�"��72�E�
�����<������08���N-䀱���F�<Q�]7U3�q&�Z�B}��3�A�P���O5��g��b�4Y2��5k��1�'�h�c,A���� I,/:���'����.R�c:d���U�-�Z��'����ޮ* =��mG+5<2��	�'8]�+�"b�-!MT�� #�QD{������ťD�`ڡbW��
.� ��-#lO(�H>!v�˳��q��k��{��AL�<���ɑe��Ń�N�8{���AAH�<r'?P����gNQ�S0�9CB�E�<��@�,�v5�OJ%]y��Re��x�<� �Q���˸br��)�!`���@c"O��[/���|�Xe��A
Tm:�'��O���c%��v|XьD�����t"O��PU�>Xn��cӊ��y+��Z���O|��Z��� rU��lB�>nt��'~�����\&��c�U�(�¥c�'�T3a��(9��E�0�W�%DI(�Oң=E�TA��������64\�02ER�y�c� �ȭSD#Λ-�\�tBV5��4�S�O�&D�RfRE�������҄�/�O:�'2Xq��l�,i4�ajB	�5+۴�PxB���Q� �刻D���J�B�"�(O��=�O�YSL��T��6L��v�����>a/O2��$Q;q*�,����X�(;���7=�aR�OX�a�1>C�M�}q�`��"O(��c�>9�ڬA���Z���i�a|B���pƥP:D�:AS �#H�%�d'D����/.����[�MEȁ�U�(��A;�(O��x1S�kT�^κ)q�mH���"O�����UEP)R-ўnS�u��i���d�=�~���O���u����`�!�Di��	��Z�4$F!�FB��UH!�D��wn�Bċ�P-.�8���6u	!��F��(�5(�( 0��x�i�'g�!�$D�{���FS�K �=�ˑ�^n��*W�Q�"|�Gd�IN d�V���$��IW�<��g�}"�a�JJ���f�x�<A'���:}�\(��X�۠�H����i�)�=��'���s�g�$T�`Xp ��/Y��uz�'3�a��O�_�IY���V)"��'B�:P�'�Q+��7>b�����G��Q 	��?y�O��PG�2L�2H ��>x荣��94�TC��B�3:�*4j�	uz~���"LO���q��������֡e:DHi��c�hO?��@�	�l�Ib+R�2�z��៪�Q���剙jUN���]>ڌ�`�COy��C�I& ��9�M:��}2$,�;1y�C�ɭ|W ���<��q�1���B��,n&�KY�!��ؒ�#��B�I)=�ʽ��-ū0�����ݟc��B�Ɍ#�2\P��͕v@@�K����B�	$@;�oR>�,� �I_\�:C�	[�^13d">M{��
�(�<VC�	 J��Y�f	��E�0O͞j�B�I5��0��h ��(v����B�Is�9 a�-]h�T$ƇwTB�ɺM؍�S�[����B rB�
:���S�	�lߜ���ᔟ:�pB�	�;���̹,(��w뜴>�HB�	�$��$�6Þ�g,�yA��ABB�3ʨc�j^(,)�a�g��B�	�w1�ܓG�9�(MP�+F%f@PB�	�qq"�bV�=T���3q��B��<d�����ױ�4	�ɚ=-\B�I�oZ � �gʆK���  �1C�I�U$��B���$
�r��b�C�ɱlW�t�E���
�7/��P�2C�	%��q�W:T�2���
E�BB�I�o02��P.�o��e�( 0�B�!L6��2��
:2�hR����C�ɞPT,*֎�-��`!D�O�zC�Ɋ/���%��-m �0��W�B{^C�/" ��x"�-0�M� �LC�	�p�d��C�l�칡!�Q-`�TB�)� �	'"�����(�nPG���Y"O9��-�5�H��� �!�T��"O�(�׍K6h��Pd�^O��Ke"Oŀ1́�j���`�����W"OH���J]=�@ؚӡ2�x�"O�,b�˝qB�U`k�,iP"O�I1�g�+E���v@�3�H<q�"O��B��U8NO�A(���:2���"O��35H"}����ۛ-�r0��"O�г�N�8�Lə���%M�V�	�"ODTî۷]�^U����(�@1b"Ot �M�B����U�2d�@�"O��C�9�}F��}c ts�"O�q���(4�V�9p���nI45�u"O6��N��3.ؐr�Z�V� T�"O��w�od�e`˷0�:$"OL�WL��b�� 3���-rSR\�"Ot����;~LnTk�҂�x:"O\82�����KAb^;S�N�J#"O�ʤ���৬C�*�R]��"ONA�ƭ�������i];��"O4��&�G�pzU 3"�2+��#�"OVu�&fJ�|�A�#�ɴV�� ��"O�q���H�R���@!U*��"O6���d�S�n١×��j��"O�+��10�l���{ֶ"O (Qv	�.E���3�
� g�X�CR"O��i�%�!b�~��	�����"O�� @m_!ba�U�O=�PȒ"O��{�D =��6�]Tb�Y�"O��x0�B�cJ�8?OE@�y2"Ol�i�ͻ9~�dٕ�3)��e"O� H0`�N!r0��ܒ�`jE"O�4
RkA�*��U��;>��"Oά;��
��}s"M&�z9 "O��BEB�H놸��ރ�b �"Ox,�0N�<���D)���DR"O"���Țg�X�רŒ��`:�"O���W'�iܝY�fì��h�"OJs*	�b�R��ۀ0��=� "O��0O�:M�܉@#�w��}��"O�a�ƚ0&2�jcC�}�̽�W"OZt�M�#����b�ƾ�	�"O��*��	�i爁���>[(���"O�\*��:f
֥IЂH*@ı4"O ��E�w.Z�2��
*���f"O�P�󍈲bxTLs@b�R�ɇ"O$\�C�V�`����T�P($*1�"On��!�*Vl��s��6�8��U"O��!P�>�5ׯ�R�`���"Oa�A�k�zq�rm�.xvF݋�"OP�#A%I�?=F���[�g,�"O�-�l�
A��2��ۈKs`l�"Om�� � �`�����8ΠI�"O$8��	��6p�Zbl\�&Y쑰s"O��a��=-x��1kȌV2�� �"O,n ��x�cdϿ4���"O
�2��ӎ"�hA������R�"OD��刔�6/��a"m23�%�"O���VH���b4��G��Ƙ}cu"O����
fق HD���7���p"Of����$AOx	∎�x�"��r"O@uL�=rFB8��$.��3"O`�ˤ�05�Ԛ�f�>�,�g"O� �<��W5�"��M�9mV��"O:ܡ�̓"�!�E��͹�"Od�:��õ%)���p@��"O������)�: #	�*?�+b"O\�b��jB��
�S^!�@"O��k���3Ԛ��$���Sp�I�"O�;��KS��ŀ��W�L�&"O��c��B?g>V)�t�3t�>D��"O�()׿�����
^T�4�"O�}o�J��	+0M��xr�I�%D�����%E^x[���
��A�/D�ĺW��$xK�)�T��Ţ$8�!�D&.#L��H�Z���Y�@�(}�!���&��KGD�95�ȡ�ϊ�@!�I�k�zx�@%%���h�-�='!�$�k)Z��p-�r�tٳŭ��T�'�pѣ���[�SܧM�<:���F�MZ���?,~��x�ĨR� ���q�I}Dy�W@-���xNm�~&��ٱdU��i����KF�p��'d�-�Tmr�SⓎ$�P)C�
��!f�<��Ԁv����'�U�G��\r�'����Q��!{���J7i�cZ��S	o�I�b^���O��Ӥ�ָM�J�'���2RD��4n�XK����,%���
�'NZ��H�"I"�D�wk ?7z�EL��Z�J1�t����#cg�T�^Q�O��;ӣ��~�ᴎ��,��'�J����R8nx�P�'�$�Ӗ��s�2�I���9=ʮIK���:l���q}�m�V��|"��7m��)��ŌsMd�1�H����	���r��P�{Q?��
)�p�S��)� �Ӷ,>W��"�f�1ʁtX�H�4
H��Ç)��m��U�e�H���'�&���+�vbp��9y���)����H�	����H��æN ǡ�����h� ��X5�@Rc_�v�b���l
�P \��U#��g7�-
'���YϢ�S��*1���*!Yc�u�s�ܷ\|`-��ɪ>�t��vaO<p�p˓g�@	"ɞ�9�^��K H�A������O�L)�$g�g�ɳ%��� '�N$�lۓ�	!|��'�L����ɒA��	j���t�,Y���c'DTI����6P�ig����<V�'�؝�����q:���<k@]:@�ܛ"δ��j�yc�SC�4��5J�h4��gi}"��C]�[�*�9S���P����?�΋A���#��y��kEܠ,4�ӆZ<.�h�(�VR��B�ӿo���'�1�Ȕ;��ͣQi��8�+�G�
eYP�	�6�N�q2�U,3s���|���	@�Z�"��;7b�3֥�{MR�L>9�%Vm���$��,WJq���ޡ%�ڹ	�MT!W�I=�9����k���@ʁ�*��>m���5O��95+ڑ���#��6�T�T�?�O����ሖF�0�[�?!Cd��@�Z�M�|IM��$���#BD�~���'��	��3��CMR�k�%��|��h�S$	�r@��hd��AW���鍯���y��ȋC?]($�J���=���|pn}5fי"$��E�]�';��g病Thn�I��A8X~������j�i�j�^m�FjI=����"O��Kf`V�z��B����(��O� ��K7P�ӕ�	�5`�1 �)ҧ@"��S;H	j&BQ�:��ȓ/�d���e�}Y\�Y�I�(�r)��ˌd�aat*^@r������|R��\ͬ%k�@ݗ&� P�oQ/�p?Q��	(A@f�����:��$	�dؑ4Ԉ\X�)оn���#jLJ�	q3m����<٦��d�'�H�g�P�J�a_*,`Q��qR�� ������q��B�#�0���O3f6r�q��F`�B�~H<�΃9EI��C1F�M(��7�V?A�D\�2�8�i޽|���R�A\#!EԽ8�� �&A1ּy�̍ά� w$�7��x2�Xr�:M"�C�/�H�q���%j��iqg,%a~>��b�T�Jx�֊�s�>E2ַ����xb�2X���s���vp�s�,հ<�Ǌ�V��$��Y��j�pf�����`��͹~ViJ�@S���@AȊe�ҌYr:9;`-,Ov���Q3r� z"�Q����>��̖��1�GMqò8Jn�BH�hQAJ��x�� wlK�n�"|I�B�g|Z��*md��Ɠp& ����U����l̚"���X�`�3Z��IE��?l�ĠA�(�q"$����i���y��H�^��C�h�h,��"`ɂ�Pxr0	�ls��.�`H��' �,�s`	5��ʰ�i���B�=��k"�Fy���06�4�"�#̌����q��
�p<��k��6<r�2R����y2�-� ����Tb��R�A�l->x�G�*o�L�0�/�O@qH`�� f�� ��H�r�-`D�>I��`�8D;`hF)����R��0#O?�[6��C�,��ڇU����$D�бB��)hB!�gVh�"HXDg�.�&��)O�u��!��ܸ����c����o�����5�
��S~�aɁ�\�pΎtජ��2����e�o�)2�Lȇ�>i�f��'\�!4`ζsZ1�`E�hX���Ȁo�r�Q�T�r��N�&L�5ꛏg_FH�ō�<��W�n<�㞢|ڄ
 �+��1��AԲ4Ơq��@�k�5Ĥy�� �k>UYĆ��p y0$ʦ �v�	rD0�DȔOT��3�(O�u�s�
�N�ֈӤw*��c��'��q��A ^`e�P�� �8$��,߹Q���5@f<`��[A��vdC #ώE����x�'� ��$;jA>�|�1e*nK	|JQ��B�G�C䉥^�l�H�k�5;T��d#�I�<�ɒ]�䝹a�����S�O�XC'A4k�`��3Å E�6h�'�l囦��_]��B���en(qW�<���M�H���	�d=��"�7+�lۣ�E�-MT�U W�p?�ŧ�xд`!�nI�m�x +w�җg�X2ѡ�W�����y�byL�<<�Z�4F
K��EG}r���"�\��3鄞Ja�O�1����t9��$-0�	�'!B�Jv�H�^���#r@ܧ̈́�r�'�����8$�U��>E�t�^*܂�㞑�d�Z�BB
�y��K�H�y�qKG�]��鐏U�R�����Z?F��2ML�z�����(Of\h%�Ҋd���&��	DP;��5b�`T�=y`Bڳ@9:��u'\�5J!��ӰdS��0�dP��;�O6�륣S1s��4�#������ 3%�:]=0�̍���$�t�lLR��$Ι����ڛN���*��*[J�a�K�i��{�$��u����>OV� t�W�2,�\�$U�e����`�'�p7mN̂����Wv}r���7'�@��t�8n�#�f�/>�]�bj� &�O��b��+��-O�A��
!��� ^����t,f��sӤS8^�N�lp�OL�H�th	��pzP%0Ix؛ro#8g�$B��V# ^6�,O�!R�ݘO��1BA*Y�x$��#B�o��(ю�Bh����ƣx;!�DA�	B a�g��|"V�
���?_�0� ��4s�5�W�>�ߴ�M�ւ�9d�Hʓ�5v�ȉ(���I��\�K��)�v��;G����U�@߸�#�д�?Q���7/�f�b��X�[���K�<�"�+E+���*?}��T�\b?�k!7��A�g��b�
�A2�I[�@����.N��>��E-O�2�8�h%�H��bmcU`>}�
ԑ	- ����'�<m0��,�(����n�l)s$*�$��R�>A��>��.�(g�pHˤ)��&%(S��V�<�0��<U�-:Aʖ?�pDҶAVğ��eZ"�j���	Q�D��MU3���1�铻RE�C�	�@�t� �%�ArR`�/lˀC�	�}ň��V��>��t.�1_��B�I�.ZZ����ң^G�l"�+F�jB�I��(�Al�>������R��"B䉑'J.�A�l4�Z�����B�	���%*6�3����C�@�C��:�ڝ�E� ���y���>>z�C�	n 6H2c���kӋV�h��C�1C������I�<9hbђ�|C�I�\����B*:I��K�DO>OG"C�	�m�ؽ)���,8��82��
��B�Ir�6Q �dѐS�%y��^�Q��B�	��.Q �M�0��E��V&�TC䉙C1���
�(�b�B(KwBC��713�#',�
gr�2$ҨH5RC�.@����H˝\�\0sa)?/�B�ɩc�.�ð��$X�Vt�5jS4w
�B�	�-b�$��Nݒ��%�!�Y�C�b�4"�U�`p�}!N³r��C�I)����h�e����A�d��C䉕^�����IR4�� sDϔm�C�ɔ�vBk�����%�Փ	afC�)� ��1B���z��g��8�,�"O���9�T@qB�(�%�0"O��It�X+;�<�s!�\W��!7"OF I���$}r&�{��Dl~$�q"Op����t%�����KST&Dx"O�IA2�D�%!�#�V�1[�Yɐ"O��+�4�ָ�N��E6l`qR"ȎJ��Z-�����0H��HQ"OV@�ǓJ�0qcP�H">��B"O���O +�48��q�,��"O��j����(�fQ٧�ڽ?�|���"OJ�I�D��^�5���B�ǶX�!�D<��Y�E�'b6f�r�͂D�!�&_��`���J=�A��%�n�!�پRG�("��W�8�ndS�D�!�$X+3���P�ǃ/oKTb��Sq!�dP;�2E�8� ('�Y�B�!�Dս.��sK3L�Q!��/~!�Ēu]N��ǅRS(���<�!��76K��&���:��}h����-d!�D
9[�.p�ba
"%����g%�&j�!�䝐HdP����S�S�p)q�))<!�䑂.1��E/^'dǨD��ð/!򄌃9��p��*��1�B�qB��!�DH>=e"�jA�y\D���[(R�!�$_��� ��;{)XK�'8�!�D
�0mJYa!�?��T�34�!�$�a.����4E�`�,��+�!�N	4u��`5m�.E蚄�R�=7�!���X�L�S�)	�BAӕaR
�!�DT�>/xPZ4��.�h���F2O�!�Ċ$��E��:^�J�K�&
(�!�dЩSmXE`�����(�7�+~~!��O����"�����W`!���B�Ψ���̗M�&u�nĢ�!��l�2���J-U#��l� YrC��SNV�©�!+����KC$C�ɰ:��C��F�<
.����kB�C�	�X�qAr��*w9�<j�����C䉹#C���&/�?Z#j� �	\�q<C䉫`��a OM9W>^����ݿ��B�	�8%���'^�"�b.*G�B�Ɂg�6���'�!�08`��^[�NB�Ɋ�82�
��z�H��Kں��B�I#w�$}�g�R�v@����#bvB�	%P��p���E5�M��/W��C�	�e�T�3�V��0��]W�C�	�}�p��U� �m��F��qI�B�	/\��������{W���A�7u�B�	�h7x��`k�{t{�F��q�lB��_��Q	E��%0��AXQ���B�I!\?$%�tA�.n�`%�.��B�	1qm��^4���!$)-\�B䉝s� H���,U�IC"�0 �B�	�e���Y@h��dۦ!q`cD=v� B����e�I�6xy+b� NN�C�	:�|ݚ�N�9]�G^<��C䉖`�Ȱ��'Y�c�>I�e
��w��䆥5�T%�v�D.^��ey�˃�[�!�	���]���"G�L�F�K/$�!�$؜a�ʄ /�:gu���TEF!�D�W��8qC>���o�,H!�DB+�� %2Q����d/�"`K!��; x�����ۂg�@{Ԁ0!�� ^d�A�[��h���ñ)�z�$"OJȚ��_'U�E)�F;>܎��D"O����NEo�	h��2&��d`�"O�]�dI9��p*
H�.M��"Oj�����:l�x	��O��I�4"O�yz���=&�2��w��z�I�"O��j��
/��A5-�B�A!D��!��Ŋ�"�6�-���5D�D� 	̬$�桹 K@{�����5D�<�p莜��
��by�ѡ7D�A�DV)�F�K�&�m�.�z��4D�(�Pɜ&p��*w���iZ9�a4D�pȧ(�vq�l(�i�m��P�f0D��#!���i� 0	Ч�if
АQ!/D�$3����V�٣D���iSf�*D��X�'�	 �ش��� ;#�I�#�&D����H�+]D�����.3�݋��*D��:�N�4�X�X�MJ/Ð���n&D��2�M�NRph���3M,��t�8D�t�#/\����tl�0,Z���"�DF0-^���{��ԧUS�$m��&[��L�GD�?�y��_"K����$�,�j�+ׄM�+=�q%��;�$*���ēJ$B�8t��e^�УT�]?{Y%�Գt��>zqO�O%F䈣B\%98�0v��u�9�W�;-�I��#A�������>yz)�R��{sF��1'�>[�'rB��a��?��KЕ_�tĳ3��XCU��- �
 Ju�ܑk�ꥻ>�����Q�$I:��1d�e��� ��
T�r�d��B�q� ˜<Nt�`�>�B���
:���: ���Xg�U8��"c��=^�:������N�@�@�����7&�d�J\����'*Px�(�V�g�I�e�tCt	ƤR��i��d�l�'�4 ��$�"�@�D��l�v�(��U���P�A����<��@0gS�XvU�'�6T�B�kv���&P4��53 �$��� 6o��П�1�� �~d�I#�>Q2ǜq������5"V^��� [y(<�3���1�~Ԑ��'8h����w���{cjƏz��p��!�/R��w+[������� 逘���+�ܡ�KHb��xB�6�`�:ή��$&���)���V��"��*�\�1"��Z~Rj��W0vc?OL�w�ؔu�5����K�0�k�>a`(��}R�d����J��A��v�h�G.���Y���(O,�͇��>1�@A,o�@�shU�V
���v!Z9v�����7-B���I�@�~� �ܵ���@�!K��[��+&�P	`�n�š�$�*`�"�ʊ�=�C�m	��x9�b�/4���ɣ� �Fݘ��q(��)� 2BB3�V$h�ZMC��+x&��D�k�Bq#�l�*��d�c�8IA��!l�yf�?|5��3��
:>�u�<RS�E�¬
�~ɀU�&lP�|Δe��,ޑw�?%���0QȽ���?���[��G�AIޤ3�<�O
0B�$éE�u��B�^Ny��! H:��O2�E9�3}�m��)�>���"M-}ƈU�4����x"��F*�-���7�t���Ӳr���X�b�j�ʼ���.̨��m�d����M6���d��V
|`��<A�n�	G�.)H�ϐ"7s|`�K�a�<ɠ�a���Z���j�����C�j��T�ÁI5���� P0^�:5R#��`�1��"OZL�$!ٹ��ۤ$0���!�"O H�&�^�C�D� `�ڧ���B�"O�)�TH<c6�x`dƏ�_�����"O����Ĝ,(o�)FD:D��"O$��QC(G��:��34 քQ "O���BϹPVLyS���1"Ѐ��"O��y�&�!Y�<�`��K�8+,б�O��`�EЅ\�H���R[*4f�G] U��4�O��D��z�P`qIűf*��Y��'��pB�a�PT�'����e:K����lsơ�	�'!H���ɔw����eAuR	N��Q��
9�BlDI�Of�e�"�|1�ň���L�:��
��� 괈�̐;M�L�b��wW�����ω\���'��E�Gg�P�g�I&T�J1�jS�D�}���$u~B�*O�p@����8�ι{nО[8ne	�C�L��؃M{X�P�ub�%�<�q���]i�
$Ol�P�
i`��'�>Ⴥ\k���Cg��9�"�kA��\�<��!��}z�Ⱥ"�7Uu�E��^���l����B�>:"�0%�b<���@!҄e��\CF�T�<�w�ة)��C��[-�x�`�{}����[��x��z>q��'ق�䃔rS%����c�����'���TO�l���ۈ-u&�RF� "�䵺�-��\v���$ۓ	�`��Bҝp7,�kW+��8:ayD�%9�dL���Dy�L�$bf8�ϛ�%R	b%O@����?n�<@�{���CF��y"�K"_*y�ǩ�/��'^.q���D.�a��fяP�6���/
 $C�lI7�X7�ē J����1�p<%��3Kj	k�
Q�x�|}s‛w��<�T�MȪi�4�=j�4p��>���i�'M�!�ğ�#�l�bRǂ���X����5Q��2�*#<@�7��Ha*H��O�8:�҉)�^�Zo!�D��t���C��2h���E�ݽ>!��֟	�ؤ!��/��)ڧBYv�v�łd2��*���<0��=�ȓ/��j��6�ł���eH:��"Y�H�fK��PԂ=�@�~�?����/H@~xQ�N���H����O��ȋ��F)Y� �y��B�B~ⱘ�])`�
�H�C�$���	�3�e[%J�1&t�����@�>)cNѴS�\�qâ���'dԈ��c,&ɂ�iV)��F����QJ�A)�OV�".�9���V;���R�n�x"�N$��=C�S�"~J0)>�Y�`�m\rHr���w�<I�fHN���
�a�� Gvo�$V�
���0`��73,�g�'r4���Ǜ&x��8�n��`+�(��	�b-� ��B:~���h����P��$'d�n��G���a�܁f��L[��Z;R�C�Eӥ�ybM�5tΪ��'�j�kL��m�IK� j�Өo|���e�[��Q�`��ĝ�v��ɱ�p��iY�!k6d�R��| �����ݳcO��Yl� ���S�O���"��+�0ș�N�R܊5��T6!�Ve:�f�5�h��y���^j0*�M��bȬI��Y�����4G��Va�g��p	�Lئ�B󁞕:�� z"�	���$�Jl�d���7�Ҭ�gbA'u��-r�!
)%�F���7����h�#�x��6CWPmy���#
ڔ�Ud��M���)(E��"4�>)׭6C[@]BŔ!	 �OsZaS!)߫F��aP䃤K�& k�n�@���e���D�_d���r�B�0��e���'^�A��B�|�ئO?	�b,Fv���h�Z�Ψ(�m(�I>0 \Y#��#��>�z�NA�J���]�	x�c�(}��	�*F�'�}����)M.͙��Q7����/��F�Z�>��>���[?rU�tS��_6~.����]�<�qF�%�2Z�.�-��'�!��3$�4B�NVm�,����T�t���+ҭSVf̑��*D��2᪗���d�@N��@�x �6L&D��(���Q�0 � 3zj�I�'"D�BRˋaN���q D�&4H���)>D��	��Ϊ2�(	�J��.2(��:D�$�b�5GSYST��*y8�9 F�8D�<kE�˶E���D�ܺ2��i��6D��+eJ	&+������A.�Cp�3D�4��M��S~�����֤Z���O4D�ԛDI�B
d��$L���pb5D�0�tF�;qA %r�.�&*���� �$D��if#��"��RJ�`�h�X��7D�T�4΃������k��  2D��r&5ck*��ኁhZh��*3D��@�dZ�N"fYT ��u��(1,1D�X��ٽG����e]�x��$Z!�:D��kb�_2~��c/	�Lk�L'D��" �b��S���N�"$� �'D��cW�\�O�����	��.CJ\���$D�� ��k$�U��ᐣ)V�^Н3"O��qR�ފ�H`gIGd(H�"OH4�Kf�DD�
�b�Bt"O��C#IJ�0�s�ˆג��"O[Al�C��q���R>T��٠�"O�-��
�^��q��#l�4"O�:�Dϲz�j�������y��"O����أ�.�C�e�p�H�"OЅZ'�ɥnA��pѤGɌ}y�"O董e#r�9��AE�m�P���"O���ɐ�@V�q �+6����(�y���h��qIQ%	���y�ޘ�y�I�	�f)���%9��`�7�y��!BZ	��t�X遇�K?�yB-=$i4�)wc�a� pyb
��y2%W�(i��b��\(�|�Q�Γ�y�ɛ~�Q��쌙T�� ��b���y�NΣc5>��V$�In�4
BAվ�yBφ�J��@�&ĠO��X)�����$A��<Śr�D�6RO��dd���m����
&����F�Obl+��NNW2̀M��}r�O %�8h�gh��bT�"co�^�c��b>��J�#�ԠB����7�@Y�[~�I��HO>� ތX���I32s��ʥAk�Ȁ���ӷ��})fkH|]֘���0�\6m�x?��E�i~"R��?�AL#���!��^�K$>5��g�"�a� �����b�"~nZ`���f�U$��Y���N7u����Lyr]���v�O_R� ��5*͚�O�(8٦���)��%���vŬx �kUB^�p��"O�x�`�9kf��O�7s�2�:"O��Q).DU��i�[5o��@e"O��։�,b7�HS��!I�(��"O
h��e��V�D aa`ՙ@%�!�"O���p#�4X.�Y���j*��9�"Ol��7�#�L�reՁn����wQ�E{��)ьK>�Q�va�/Z�bP��B�7$�f��47$ɸ��=}"�1����!�sM6`�i�
���Ɇ-n��ӦU��0|b�EG8}��e��+�/:��ȱ��]}r-\ ~���f�M��S_�0AhQ��.FT�k��Q!:Ӿ6�[�,h���?�E���^���M�Fnδ���58�Xdn�5#��'������"�T�&%k����G��-�})rnEn~B�\ �?�'jS�%��H\l�S)(@����`00a6*�5�Ȑ�Ā�-�t#Ð�?���,�,j�l�9b��h҂�Q�{Up0���R τ�+v�柠�G%G]La��᎘e�Vm�d�v�Mh$�QVM5�O�ŋ1%�8i�@�qnɛ*cx���"OV8@��X!tuj�Z%y��YV"O���p��[p���h�"OHc��'`�\����@	#wda��"O��i�"�u�4DjUϑ�Xqt��7"O��Y���J��z�")q��D"O8m�G�ȟ[��R҉ڃ7r�1
�"Ot�Jv,U�d� 1k�)Nir���"O�铕H6w�уH�1fT嘥"O��0� ��H�����&Y�/]z$�c"O�@[�H�{; �q��>5EN�@"O�Y��k�?D$p���nW>��I��"O�1Z�+c���F#O�X��0"OVH�
�>�,`�j Z�f�w"Od�����e��'Ы@԰�hF"O�24A�(.� �+�Ʉr�(��"O��R�Y�
5H�N;%��ҥ"Oށ��K*U�N,;���F���z2"O��*�)'��yD����JtK5"O"H1"����P�«���"O|=bԥut�*G�Z&]H�Q8�"O� �h��MVX%Ɓj��Q�N@n�C"O$��A��l|��9Cl7H/P��b"OԄ�))F������,<��4�"O��Pi����y��K�(���"O�]x��La�2@���,k ��"O<ySa@����RmC/F⸱@"O�`��U�"���k��#p��c�"Ox�G��0W>��*����XW,A�E"O�̃�D_�,["�;-/w��!�"O�u��N�%Ʃ�&7Z��T"OX02u�]>h�tYŋ��]y%"O,����J*��U��
ʮ.� ��4"O؃�ܵo�����#Ũ-"Z�z�"O"���c�; 1�`#.Z3��"O�I�a �%/B��XG"��)7  Y�"O:��S�_=a�l3��:8P]��*OR0��ƙ�)M(�j�$��Xڬ���'�.����	�+V�E8P_�J�H��'�b��WG	/�PQ�B��>k<���'�}p7:����Y�p*�j
�'��#�Q-T̺l��E�tf�i
�'�u��
�6,�~I�@��
q:t��ȓ73�2ŬY�a��E�FA�tȄq��x[��N��r�D���J�K���ȓ#⦍�B�\ks<�1�h�:��͇ȓt.���p#H=�D!���ȓ��i��% w��p`�U"y�p���>�e�v���`.^0� ��)!.��ȓp�x�穇?
��d�X;�d����1�I�6�wʕ�yA����!FJ����4}�*|P�(J3 )��N���@oM'=�� H��E/G�l�ȓ&��r@J��SE*�ȸ��m���(ք�< �����J�L�1���X%��J�!g��ћs@�Z��L��V����': � �����3��p��v��eg �*��E{gg�M�$��ȓ@�., ̅F�Q*���)��5�ȓCP -S�I,FX�x�c��!�� ��L�T�x���D*&�R�͊}� ��6��S���h���m��J,|�ȓ&�Z\qR*�<������!coX�ȓU(�-�S����xuġ`bh�ȓX턐`���"|���㊙r�H5�ȓ2.�h�BK�9BD��b=1 蹆�8��<JV"��5�J�P��Э`	$��ȓ2Јj�!�� Fa�ȓ3��1��	��,a��	0�p���"�PQ#S�Y��R��aB[s�a�ȓ[5�+e㞮*�����*��.�B��ȓ����J/)7f5�'�øW��ȓ��C0����0���1]��p�ȓE*Hpș8R|�(7�H�o����ȓ&Uޙ1W���%�Ա�&Y�Q�
�ȓx��XC�'M<MJ-z���4V�=��V���@o���q+�I�/H.l��LØ��W��p���hʖX�ȓ<�̀�A�A�
����w��>!�ņȓ@�j�A��w�����a��;�.I�ȓ*{R�S��ȕ}8b�i�4n���ȓQ�:� ��nܾ �-4^D���cb��Q��JP�s3�ڸm(��ȓt&.y�ł�_��5�� �*E���p�J����
�CH�#��F$!��l��S�? ��4ht_<�Rn�~,���"OLqp7�J?^�ڝ�K߶,�j);""OV��Sgӓkך���B.�pU 5"OD�"b�(�V�1e�L��b�³"OHҦ�T�>� U�'�Ȩ{�n``"O(����X �,x�t/ēr��8�f"O��{�<>��m^ t���"Ov�pg�b��S1���Ѝ��"OĘ���/
6���L�K"��1F"OlA�Ç��6A�ҧ,
2���"O"��2䊄N��$����9��aK"O����$��a��!�cK�m|��8�"O����$mp�	�C�[|աC"Ot����Qn\e�fb��2�H��&"OL`�Q�<s���� F�@�"A"O�B&�"�f����v���"On�*�f�%N�t�Y�	P(����7"O<�E�D$k�\���ۨ[����"O��5�^�',~$r��.�J�xD"O|K�k3ZV���T�y�pE�4"O��u _�HA%#?9p�y8T"O\�`d�Їv�H@���/	B%��"O�D���6Z�Rʷ�˝GQp���"O<���ⅻZ�hB�L8���"O��0|8�9��C�#�8 "OH�ɗN��M��AX���d�S�"Ođ U�E:p=�}�7b��d�d��"O��I�l��W֬a�D��:PI`�"O����A�o~*,s@��4�m��"O@Xy��
�
������G"Or��q�E&C�� ������)#�"O���si�>(���/�P�Z���"O���2*��΀���3]����"O`�Ʃ�h� (��h�_e���B"O�����$l����(U�ZZr�zP"O"�۶dKg0�h�F�Uj���"ObE�!-	�'��X�aƀL7��I�"Odp�fI�{Vp=��䌮1D$�"O�K�/]8^ib�P�S
sX`"Ob�p���Gѐiv��\�h3"O�dy�)Q�D�b��DI'q��ѐt"Oa#S��uW,c�/̷���w"O�=�'^au��.�c�(�"O���"#�=�����B�d�Y2�"OX#"�S�l�t��v�]��a�"O�<��B��s�`X4��3X�]i&"O���q.�6�+%@ԜK�{"O�L"� ��#�V	�p��%W�Ő$"O�Dp�F�3ٖ(0�N�� )Ԑ��"O ����MQ\��cl$����"O�D��E��"}�M���<n-H��"O��H�c�4���� A�3p!3�"O�O��b�&0h0���Ɛٲ"O�	xtjLw�v�P5�ۃv�*p��"O�Ě��UR�-��NXK�pU��"O�D��+X���RM.�qp"O 92L��|s®�1OȠȑ"Oh(x �_%H��Ҏ�)�"OE#�/�*��u��#�6�@�"O��["�(
�sSHm��3"O�}�%�^r���g A���p5"O���ҧs��w��R�4��5"O:q��49�@uh�l:K"F�)�"O¬JV�V-�щ������R"O� �uyU�בJ�РWKZ&#><��"O���B+O�L@�  ��Su"O �B �#UJD����=x��Y�"O�yGڭ!2LPӥ� 44^���"O� �s/G�yO��"7 C""0@#"O��k6�
���|�­��->���"Oy��l�=n�氻�,a�U9�"O:�X��@����`�ĉ�"O��YA�8����y��"OְJ�(��5��p�@?N����p"O�zS�G,w�fR��F0p�D��"OtM�Ah��TԘ��Kq@�R�"O>�0��N���3���o��P��"O,,)�bJ<a.�� ��G�6�H"OhL�!�p{J���΄�o��!"O2A�roV9�\:��0b"O�l���Y@ܩ����Q�]�W"Ob@(W"+/�1U

�o��[�"Ovm�dA�f5���X&Y�"Oܢ�#H.8�6!q��δ��!�0"O�T�u
����v� �y��"O&d�3 �?�y91Cҳ��!J`"O����d�l� �BM4wɤ|��"ObQ
��D�0��u(U�@M��"O��� GLЎ��DX�Gʲ�9d"O6)�bd X=Ti����#~-AB"O��a�c17��h	�R�5
�D#U"O���7+	�&��Ğ�9�4$1"O0x􀑃$LX '���.��\)�"OV [RfZ(n�*��!^�$�$,1e"OND����`	���ŶP-����"O��s��w\�`�V���`#��A�"Ol8�T��1<R���Չ=,Xa"O��k�ʐ{L��&�H�G^DI�"O�%�V�D�1���+!�X[�|��"O�#��7d`��I�舺,ꢸ�p"O���mԉ>��0D��e�֡)"Oh��~����G�;Er��"O\�����PK�Lb��Y(2U�"O:��1�6{�� Q�cﺄ�q"O���"d��r����~~�2"O��ӣk�ŀ�$$Q!W8Dږ"Oj��S��-����M)x�
�2"Ofɲgd�5F�\M
W��d�(�1�"Od�'fQ�B�lӷD�<z'
I��"O���� bH&ȳ�CU�ij�x� "O�݃�,SB?^Q��b�)b��c"OV�;'   �>�I��@��Nͱ��Sv�Фz�LR��M+��)�?����?K~���qQ��w���[�F�-0�(\S�M
^��	���'�2�|��4޵[��	c�'=��p��_pd��&�(����'�N���!G矤���|�Q��''x�Aw�\���1���\��Ԇቷ�M{q\��?����?��ö<\��{�aѓbd�=*�A'��'�꓌?y����K�A� ��3t|i�m�0��'e�!OG�k2$Z��$�ߟZw�'�a3�fF*��(`�E�W�M�v%ΉLrR�'A��'g���'}��jPJ-k����`���'r'"�}ӐEiP��O�d�%��s�I!�j�b:�(Ӌ�p��dcc�x����D�I(E���o��<���F���֦�?i(r�սV�����@L\xs.�Ɵ ���j�����$�O��'6��'�v��d�t�nٵ�͜qt]3�[�|�۴���VE&�?i�����<f�� $!|�s#�ƨ}�J�����#�������	O�i>��Iş���A��"���1�ꅶG���C�P֤m+�/)?!���'����^����D������g�ښCv�9� mF˲�d�O���O�4���sD�(�evR�Z.r��x+e�K?5.�z��0Z���lӖ⟈ګO��O��Dڀ>�H���-�}
�Kߙ\N��[�ô
2�	�3���O^�'?M�=� �a���V	���0jJ;3=��R�6Oh���O
�D�O8���O�?u���u�^零����l���ǟ�����(�@����j�4��[�BiQ������6�M>	��?ͧo���� @�L~r+Z%-<��A���JW�P$��,�0I�%��p�d�|2S������Iǟ����Z�Ep�����9�a��ޟ0�IQy��nӶ`���O����O�'Ā��ICl�̑�4v4��'����?�����S�Ԯ+,��ԓc��	 ���$�Q�N�a��ź���O��Ա�?9�%=�DK�y�nh�5��5�󧉔i�����Od���O<��<a�i��12�/Bh�	�f��9QJ	+�e����'*�6*�	���D�O� �(�
ξ���N
>sV����O���շ"|ޠ�㖟@�4WP�d�~��L VA�}e�ۍpQh-I���<i-O��d�O���O����Ox�'{������S�� z�
�$���i�XL�A�'�B�'���y" ��n��szX�J��\l��(�.3$���OX�O1��C���.39�DT?tMF���F�Yu�,
E���D�Vm>Ĺ��U�O:��|��+�
��s�\� �7A�s1
�3��?A���?�-O4�o�R6���'
��PJ�K捎<Y}�POŵL��O~��'o��'�'_����	�A.`��D�2)���O^���);Wh7��E�ӭv����O	�4��%W|��桂1I��3�"Ỏ�s��KR�|a�G�0�0@�O��m r���	ǟ���4���y�!��6e><��oY�?�J��T���yR�'��':��sv�)��$X	�"X��O Xi�ֆ=��c��Eyf�Җ�|�S� �I؟����Iޟ�p�f��#�ɛ��tL� %$�[yB,k�`���g�O����O蓟��D̲��Y��O4W�\��W���`�PT�'���'ɧ�O�PaE�A�Q�:����
�b�h���
aU���O`�jFEH��?	�+:�$�<ђH�;Ad��&/I%�(��M׶�?)��?	��?ͧ���������K�ן!"h� �yuƕ!0a0̰��ӟ�y޴�䓢?�]������	9cZ�K��\ :��_�<�!�6��;���y�L���쟄�KJ~�������)m(�|xQF_�!���Γ�?a���?����?Y���O���qW�ۈ	��ؠ���r�2��'d��'4�6�_�(���Oz�mO�	�9�F��W��Sh(��%�Tc���	��t��0<嶥nZ�<���bs��gf�X��Ӂ�Vz��%�o��ud��ݾ�?YPd��<Q/O�������d�O��˗nS`�UjR�\0'��Q;P�P�x�Q�<1�i^H�O���'��$�w�f��`�0=H4�9 ��Q7�생'�΢>����?1H>�'�?����,��$�h�#x�H��)X�@DXׄ�k�"L�'��Ď	Οl��|r�[px=#2,Vq��J�&Mc�B�'�R�'=��TY�D�ܴ�6@�mD\�H��m��J�E���?���r�����b}��'2��Z�ƨrz�+aϚU����'�'��d�d1����O0ݸ����
K?�Bb�X$4���8���p���*��x�H�'r�'���'"�'�哟d��r)�s���ħI�/1�!�4Le(����?a����'�?���y�@ڷ>4ʉ�h[j8�H���/Z�B�'�ɧ�O��,�"�ɯ�y���D�$`C�%ۋ^8n@���yRJ� DH���I�M�'J�	Sy�T�(a0,	�G$$dDu�vm�0�0<�"�ih
�K�'�b�'TZ0�u��9_gV� B`�g|�<@s��FS}r�'�b�|B.��a	��{�B[�H%�a;r�G�����*��T6FY��X���P:�'��G�t_�!���:�t�S�SE0R�'�R�'�b�sޙ[��Y�2�ʵ$Idz���)�����ߴ^ ���?�V�i��'��w� �r�
�1�n'P�\y��Ț'�r�'`���(�"ݚ�O� J������ �T1����Cc�P;U�Ғ Y�L���yB_�`�	�?�I��Iǟ��"� �ul���	�s��Ej��H�R��N�z@�j��'�2�O��4�'��?�>����'`�5� C�v����?����|*���?�Fal��r��?��� ��ѡS�d(��4���ԾQ�V)��'��'�剃�A�Ui�ml���*'6��IП��	�d��3wA�ȕ'��6-׀���T"t ��I�ATY�t��
�P��
�I'������D�O
�4�f�JtD���"�[V	�_�,��gBv�7M|��ɩP������O7�e�'��T�w��٣V�V�/Iz�:���(Ytr�I�'D�IX<5��'���'���ԭQ1~1X��7S4X�T�!'�B�'D�j�IA�d�Ov�� ���%�蠱�݌	��r�*5&�E�p��L�	����ɟ�`Ɠצ�͓�?�A��s�� !���Щq`c�=�J�X�ʮ�x$������y�fW�\�x�u�I2c���a��ը�O|�o�H�p��I͟H��b�dm�~u�]9 dB`N
�&�����AC}"�'r�|ʟ�|*@
��<��5M
��|C�ȧ/�*�ҌZδ��|d��O~9�H>��@ 4l�}�"��.F�&Q�@�?���?���?�|:.Oʅn��)�l�ѐ��+K۠�dH
�~�$B��ܟ��	#�MCH>Q��[������F�% �D��W�ȱ�~P�a��P�	qN�D�QK$?�@�R����Sy
� ڸ#�F�*S��;7mG�?'��I21O���?I���?����?i���)B��T��d�g���Q�b�9}N<l�4<���I��`�	F�s�d����`EN'H!�b�ɮO�j������?�����S�'y]�ɲܴ�y2.�0(ن�#�B�+K�R�)��y�m1$F���?!/OJ��|��F��)���+@2��x�G�_�i��?���?a/O��nZ�{6@t������ɨX(D��Ĝ[�`�$�7Z.��?��Z�4��ğ�'�p�qi_?	"���F�vh�����=?qWo��oٮ5����|�'jئ��ϼ�?��cG8@�����`?&@HB�	��?����?���?)��$jѬt�/Γ$p��`jS�Z ���չe��BnӮ́@�O���ަ���uy���yG%��w�}KM�G�(��֯(�y"�'"b�'���G�i��$�O�Q�t�ޫ�:�.ߘM��Ԁ�C�"4�xg�Y�b�`�O2ʓ�?����?����?��b"�u
�N7C�08��յs]p�/Op$lڈ	����������?������		nJ�ʴ� s�0�:���QR\a�O����Ox�O��O�d�|aT�Ìp���I�	�&=Qt!	1tà�'���
Ԥ�O���|RF|̓���m�lE����<�FD�pKr���$�O
���O����=C��-[�f��L��tH/:14y&��+_��EG@���b��ī<1����������i�	���b[/K4h1(�oӉD�n��<���.�m�Â3��'\���wn��{��4}�KF��Sn�Z�'�r�'��'T��'G�%�BK��C��2�j�3�P�X�'�O|�D�O�xnLo��S̟��ܴ��\!*k��`M�"�@�$���H>!��?ͧg�&���Do~�A�;D�j$CR	��!�5GO�+30�e�Fs?������<����?!���?��P����/S��0���?i����ĦQ����۟��I� �O
 ce�۪7uJA��C6�>�c�O~��'`��'^ɧ���4E�����$;�d|X��P�%��M�Q�>F@26�5?�'%���L�;��l�Ǔ�c9�I� *B�	6�M� D��}p�J�>�ĩS�'�i�����?ё�i��O���'��Vi9j����ԗ$؊Ԛ5m����'��=��H-����xA�e
�~��,O�` �B
0z["Q���ާ)@���4O�ʓ��=�S�-j�9�
�d����1�"�&!�'S��'=�iOæ�ݯl(���a] _V����hj��I���$�b>]���ÎhP�I*OTd+n�"_�(̓%WP�ɱ�v,"��O�O˓�?�� D� �˻\���c4��LG� ���?��?!-OxTm��Z�܉�	����Q�r��E�'U��1
�73ء$�����$�O>�d0��~r�Q2̃i�n��E�F�H*�d�OHhAM�t\`�t�<1��c^p�$��?Č��6*F�y��-1�8d���L�?���?���?�����O��� �83vp� 1�Ϫ<Z�.�Oʡn"v�f���˟|ߴ���y�ۢ0&x�ۇlޏL���iq��!�yb�'���'�"�PV#�"���7,-�0��@a��H6�5
��√����e��O�T?O���|��'�?1���?��jD���F�=
�� ��>0mX.O mڡY�:��'�2�O�D��'��e	�0�+��
�rN�Xw�&���?i�����|���?�rM��^�"�2��H�mc�ƒ88����4���Y\��b���"t�J�˂H\�F�D��$�&\�����p�1�r�-���U��6��h��e$c61B��P�
U��<`I	����jYO���w��	�����֨!ZDU@��8��8
j�   	x��)YQ�����>�8@pa���D���!�@x���E*���1�b:��&3=1�����!ߔ �'�| �asSB5Bv1��Z#x@�(s���]�(��V�z��e"��<{��{���9q�"�R�Hv�Q@�"i���)j'�G/Ԥ���K�(v$�2�T'�M(O��D�<	��?)���P���O���Cg�� e҈ h��I�-�*���Of���O(�D�<Y$�ZtN����Cg���pK�y�f��,=�����ޥ�M������?��K�����{«�D�X)�fER�"f�q�m�9�M���?�-O������b���'tr�Oo�(�Y$6e�1c+,��e��0���O��DB",���'8h���&-�k��$C!ON:�m|y'H�7��O���O���a}ZcD)7��9v\��3%ޛ2?�x�ڴ�?9�H�"m:���׸O�0T��(V�܂�ǂo� �ܴ\��T�i���'�R�OWl�����~����f6�tZb,D!�LYn�����I�	o�'�?�t�ڬH�(�hP��&�Ω���Z��f�'	��'�����Ǳ>a(O2�䫟8��#�&
v���C��j��$�I/�Bb���IƟ$�ɏp���`N��-�|ՓDg��r2�y۴�?�1�ׯ��I]y��'ɧ5��6q(�葶ٸ9���+�%�#���];a�����<Y��?�����d��iP E��K4�p��X�_+⹰�T}�[����^����	LLĜ#��38=�ⷁ�LP*0��y�	�p�I��4�'��T9��`>};��ŉl�z��N���0Tfs��˓�?�L>���?���η�?���=S�D@��5[���0
�F���̟8��ʟ0�'
X���%�~B��S�����T�|�X�FD	��|h�i=��|��'<�&��qO�a��Z��ቄeք&t��y��i���'��I=$�2-pL|J����q�? De�F��^�>0��<XJl�%�i���֟������	d�s��01
��˛y�)�g�7E�\6M�<%-�F(��ɥ~����*������bE�B�t��I���TPp��~�^���O&�$�O ��O���u�ܴ|�R S�RN�`���
��DoڡR&���4�?���?��'hՉ��\c�0H����-\N9����D�A�4�?����?y����Ķ|z/���yfc��H�J��%��-h
v<@��������* /ˡ<�O��=��c�JXhf�)�A�K�2�"�)d���Og�OJ���*_�T<�c���j�$��T�i��cƒc��I���	/�	�W�>h��
 xa�y�i9T���9I<	�!o~��'�"�'���f�[(�(.T�PoGR�@PN����?���?-O��d�?	��۷B���P�ʄs���z�{���$�<����?����D�Fn�p�'r�L��w��yb$��*O�,vʑ�'^"�'z�'_�i>-��"xÌL{!�N�$dL�0� �Q[�O����Or���<���)�O�^�R�兺Ux lB��8W��[0n�:�d/�D�<ͧ�?�K?)C�G�6��(r)��U��X���~Ӑ�$�O"�:�̥�ד���'��\c����T�O�t�Q�Gɞ$��!��4���O��D�O����|�+Ok��\&\  ��6c�h�b!��A��I���bcf�۟����@�	�?���uG WU1 I*%+�?���$&˕�Mc����B�N���4l1 ��$-��p��?w���'�i֞I���' B�'�b�O�): ��S��ç�@���I��ʋ�I�Ɂ��#<�|��J�ޝ�C��xJ�{�ꇲX�n��%�i7�'L��؆qT�O�	�O���9�<�Ek�1 �p��[�B�J@mZ͟��	Wy� �~Γ�?I���?�p�Ά<� Q��\���\�`X5���'��(C��2�4����;��*MϰD�s���Z��"��� D���$���I\�Iȟ��'G����H��u��j����$[(�Z�(���h�?����~�ǂY�P��W�B � �Mk5��d~"�'�b�'��<sR��	�O��l���P `	���Z=�޴��$�O���?���?��C�<�$��n��Q�L8�� ���2���؟��	ҟ��'�h�肉�~b�n���_*w���(�+�W�ؠ��i��_����Ɵt�	�K�����`��<x1�&l]�`�JC㘥 @8m�����ILyL�T�맜?1���b��ǳ<��Zs�[���¥L6 <��ڟ���ן#�9�s���|��;�ȋ�[� �k^�7�imZQy̅ ^\\7m�O����O"��Tk}Zw4ޅ�bffm9(�*�2W�.9��4�?I��b؂�͓��$�O�>}��	�3Y��x�?pv���gd��4+�����ߟ��I�?Ey�O��P��l�1�U�B(����
�fS���ĳi���'�\���
�4�:��gG".��@`ɏd��k�i�"�'�K/b5����OL���y�Ҙ��S�,���CSj� g��6-�O��$R�S���'Bٟ�D�!�ʡ5����483R�qc�i<2͈*S	����D�O4ʓ�?������4�cZ�#F���'T`�'3��'��'x"S�H��<z:��3���*���ͅ c��!��O�ʓ�?�(O��D�O��dZ�RJ�pJs���/Lnp�eθ8>�5O<���O����OL��<AuO�{a�Rqvp%�1b{i�$JcLW�+[��^�\��^y��'3b�'ev5 ��5f�ڣjdXx�jN�-��
�%����$�O��$�O��T��ɩ�U?����jӊ`���%H/��1a��P���ݴ�?),O����Op���5��'ʅc����@X"2'A#j�(+�4�?����dE#�<�O���'���I	�]�S�Y�z�J`X��G�D��?����?���<�����?i�1��"}�4�����]�N��%�w�d�U���B�i���'�"�O�N�ӺÕ�Y�a�����@���K�Ŧ�i�n`�@�	��'#q�Pp9�-y�!�Q�f���ҲiFR��"Io�����O��������'��ɧn���+��mh�t�r/Q{@��ٴJvD���?a+O��?��I�"2�ъ��΁|XMR)B#L7Lts�4�?1���?�!�͉�'�B�'4�$ܸ��
��"n�e{[r��ډ}��'�R�'�¢U��,d�4A���ҩ�a�b6�OV�s0��X��?�*O�����A#�N��*|������ �ER� �p�ZşԔ'ar�'*BS����U�9dH�D�%��)�@
!
a\�K<y���?�L>q��?����y:�r�h�#
B�JC�V�Wt�������O �$�OT˓X�ڑ:R0��48���]3Jɡf��Mn��j1Q���I�(&���	퟈��|��� ��4�n��GE�2��BҼ��D�O����O�˓2l 4��t�= ��P�D'���V��e��7-�O��O���O�q)��(�l	�V���6�y�#���F�'��Q���#,����'�?��'��E��M@�$�)��K%�`{u�x��')rߺ�y|�ڟ��Z�H�8p
�D#��ƛ/Fl�1�iJ�I�1n�$��4C����S���D	�1���A����8Hg�'�&�'7r�!�y2�|��ɕ�wT �ؑ��7	� i3���3�����T6��ON�d�O�)FJ�tT� �C6#p&�!�4�L\I�p��i�R1�'��'����D�^=�P��L�ouz���F]"���l�̟��IΟ��PG�����?Y���~2��qr�k��F �B�׋�M;N>a�`\7ŉOxr�'<Rl܇J�p#�(�>�Tʝ*
�f7��O�$�%G��ҟX�	@�i��Z��_��ڤkC�[|�1hϳ>Yd�U:�?�+Op�D�O0��<��W/ n�B�d��D�:�*G�Y�`�������OғO��$t>ݚ�cS�?��p��1$��y��� �:{4�D�<���?�����䚑	�-ͧvW��\��g�ٗ
!�@'����w�	���	'�T��+�r�LZ�JѲ� Q5+��\��O���O��Ģ<�ƭ�!.��O�\p�EK4��ԣv�y�I��~���6���O��� j�l��>}"G�?CC4�{g�ڿ^G��2����MC���?�/O�i��Ba��\��;C�����6��j�+Z<M�0�I<1��?rƕ/�?�H>i�Or�qQqʗ6D���H��Yݤ1�ߴ��+�즽诟.������'$�h���t�&���S;�����4�?��8+~������ܸOeJ��!2pO܉ ���7����4;젡0�i��'sb�O��c���,�(�\�!�����Iڒn�:�MK�L�?L>ш���'6� �Gf8���_+T<2a���l�\���O���+HSƘ%��Se��ƪ5�B��ź���?W���p�4��'��8�d�O~�D����	p/���� Ab�t�t�Ц���		I��H<ͧ�(O~���CS�m��e3D�[�Cѐx��'/�ן4�	柸�Iʟ|���ڇ2e⍛���R�Η.X���Cr��O��D�O��O:�O�$�� 0
H�O���3q�RD�h��M|Ӹ�R��X������}y�KQo0��S�
�@��R#�8��2��޴듛?���?���A������x��h����Ufr�YC(��IП���ӟ@�I�� mڢ���O��r7��'`���D�+1�:4C�" ̦Y�	Q�	��\�'H�t�H<�6�<{��|9�,
V �#�ɦ���Py��'�v^>���ȟx�S=x�jHQ5�";�fQ��ɟ[t�p�K<�����U>W��]0cN��`%��{y��C��
\�67�<�qm�k���k�~��r���lc�4�rd��@᪡a%�{����&�O�, T�H 1A Ѱp�@����R�i�p) `Lh�^�d�O�����|�>iT�{F)af*+|@��b�6�a�'��R	�}qQۧ�I� aH���~ӄ��O�$��t�l�'�,�	Ο���In<x ��^:�2����S�P�j��>���y��?���?��!T x�v�� *e#�C��L� :�F�'Y\}I%$�$�Op�$$����q;%FɌ&��eZf��1sp"X��Q�\bP6�	�O��a�̐��*	 cn��J��!��F?!^���7�R36}+��U�WT, ��k/]�AX!>��=����:Ni�4F9�Ifx��G�\�9����ϣD��>Qs�׏~ĉۣ�݃g� �T.�sT�KP.�P�r8҄BZ���b�_��:�h��(G<�[@J�',T���+�|��X�� "�
����P�"�ʘ�s��,/��d8E�C�y�`����&#���.L�Y�zG�E�3:��8#�:A�&9V��K����pDDN�F-E�0�����M!�B�����"R��I۟��ɝ'��&	� 	%�W����T�[.��E��y�b=9�)?X�Ȣ<�	b�>�)�(�/b�vaF0G�<)`���7��i�ҵ8�y��2��Fy�����?�����Om0m+bG�8�� Pa�]�
hHx�'u�Ҏ��V�W P�$��%:Є�0>9s�x.�7	J�I�o�{1�g�˳�y��.����?.�*8IWb�O��OJ�P#��B]�C���~�Ӓ��=A��P�Y�H}va�O�h�矔	 ��8�tX�EH����[P�A�(=�<�L��6{���\�"~����t��5�6T�rl�i�1z%�YB�O�П��Iz~J~�N>)��'s/
[d�}U��;�ju�<!D�ǍG	����'/<�b��#<��)��Ά�6�ㆨ�f/����J��?A��y���)!#.�?����?��f��.�O���X�Z� ���U#tSʩ�$N�NL��Ŝ�����	�W��㉪vw��'�f�M╨m�ƴ �'��)���'�Y�Հ)O�\��@ާR�<0y��K/Fa���w�O0�B��'mr�IXyb+�'pV8��̗9�y+B�S��y��1G�ʜbN�wN���#)Q�r#=�O��I*y,�0޴W��ѫE�S���iҎ�<nI���?����?�H�$�?Q�����k͈|�H��Z.��tIӧ�<9�xj��<�R��B�!lO�q�aӑb2������/��XR$�R%HD���_]�]���I2����OHP��[(P)��)�*t,��`a"���OvZ@xD�N���U`]��!�d�	c���qJ�Py�=([����2O�%�'�剕J�p�K�O��d�|�4��p��k��Y�&<�f	I?�zY����?��f�Nd�h�O��(�T��>�O��Q�B���X�e2�Mߎ`� mC��-.�鋳M�~����}� ��5A^�exd�g���3�"��t剈M���O�?��ή_v��T�ʁf"a������	����
ۺ9(: {օJ�&ǎ���L�ID��Q�'�̆ �0�&F�z�z扅	i�d�O4���|�LA��?����?���h#m�P�ۓY��@4�bC���5@\��`�P��Vr�*�2b>�$J/v7��,m�`z���v�&%s��u�L�# D�WO"��S��?AA�
c�	 ��m�d����8C歀�4s�v̭<%?��S[yb�R�Z(�1gی�v��b���y2���j�{�U�i��\ �O�`Dz�i�>!Ǡ�aDh��@�Ha1:��sk�.�?��/��@����?����?q�@��n�O(�$�gI�R��T����ѭ��j�	$�.�0�N�?)��ИR*8�*g�R !�'
bx��C��|���'R�+��.h~�� �A�$��O��
�K��8�<s�J�ex��yq�O�ȁ��'�:6Mڦ�?Q�V?���ӗu;$$i�P�s��䚀�0D��*�c���`q�mL�>U�� �HOf��'7�I���"ݴ`t9y�g�+f=�1c�@�~���?���?Is���?����D���?Q��]�:x�c�H�O��ȐUmԚ�rQ��$f��T�2!k@��(� �c%.��Ɏ0|�D�O:ebMe�}�V�Ƭ X�7"O�Y�)��8�pl�A�n�5b"OVE�&��,�a@�'�r�h
�=O\�>����֛V�'rbX>�5f�Uz���S*�0������Y���I�0���(�f��	I�S�d�V��~��ŭN�|N�=�6Ü�(OB%�$�S3g>mzqe��MB$`�Vi�F�&�<Y�mR�@F��@�&vܔ�i��L�7��`�g!�<�yd\mLi���4XR]r���0>iU�x�@� 
��P��^�To����,�y���/_��7��Oz��|
`NL��?���?�a�%��4��N�#g�������p�������I�j� ����"�F-*S��",���AS`�Y����2La�);'�L�T�����lS�A�T�'�1O?��\�_[d���Q����-a�!���&v�K���`��qHmH�{��҈��?��(��d��軖�W2��(�����I1>qT�B *C؟���ΟT�I��u���y�HN?PH��FO�	{� ��E���~rbH+��>���|��i�3�M�,D�8J�Ɛo?����Ex�T�P�y�x���2�Ԓ�$��ԃ���O*����#A��q���+�����
%{!�d�4:���9`�	&D֌���бd�ȰDz��)΄d�4IoZ�{V����K�Q�LRR��p��Iڟ�������ph�ϟ��I�|j�N՟��ɓi��PY���fP�C��7L����%t�IR�Qfeȅ-�i�խm����D�V�B�'�0���mA����_3KE����'������A-2 ��;Cf� ��'X}�U�ſ��4ꆯ�\� K�'ڢc��h!6�M���?y(����>�{��`\D��$T���d�O��ć����,�|�f鄌~*,������`F�ūp)�s�'�܌���	�1��ғQs��l���0R�Q���O�}w�Kc�"�ǋS�P>�V�i�<�7�I�{����f�#Q~*���\�|sM<���؛yo^%�#��c���� 	A�<!%,48�IԟP�OA�Y��?���8��8�4M�/�c�IK~�,C� �|��y��D����`���C����e�'��s��"S n��.u�D��ܥ���fH�~��~�IQ��mY�gY=Ef�5�f�	�h�t�(Տ�֟D�IJ~J~�����$λq�x��EQ��ejs�X3Z$!�dX�X�L��B��h��Q(I8X/�����?a"�(�
g��q���x���`@⟐��T�~���؟,��ҟ(���u��'��ڹT��Ъ���/Ҿ�*��ء�~�b[���>�c�(�bݢv�U�����r?��mlx�P�g��)��%yN٢knN��v桟P�Ĭ�O���I>k�t� 6�،[�x`P6T9#�!�dH�\���\
x4 ��/�x�Gz���\�o��Pl*	�T8��@�FB����7N�������<ia�Z��	�|Z5�� ����mL�j�p�BH�U���ǂ��3Cx��B�B�ayrꉛ<^p�ăD"p�$��	yE#�J��!�=~����D��B��� 0�L�,Z����Lɑ\����*�O��E��'���I"nX�1!E��w∨�'�����z%��W�$�'����	�Ȥn�˟<��G��K��Z�N�;d�ТJ�"����0JQ"`�e�'��'�P��W�'�1O��h�"u
���'8�5c�
lת�<��+�L�O(�����'k�*�R�H.-6r�ى���,��u;��;GX$~���AiT<{fDB�r
�*���ڢH�૖�e����M{��
Ezjap�ٻ!��;KS�Xb��I�e�~��4�?�����$!S����O�����I�x�i�^9"H��QQH�8QN*5�9O�c��g�'����� ��[8���d78���R��&�(O?�ǫsM0 [��	R"�����F#p�*�d�O���3?�SF��?y�)R�3;x8	��ێF� +���<	���>Qg�ͭaV�i�aL�!rH��%
|�'|B#=�OS�ZT�ԐU,�x"��� B��'a��=
�\]	0�'iR�'��w�!��؟쁔�Q�?�܄s�F��	�ٳvl����'�0�O����(�?gd��E��+N�,�PU�Op��c�'�T%�a�����"gͥM��1��'X`�`���=�El�tPSFl�^2�$r�Pb�<)t�Ͽ&2�3`�Ճ\`Ը1Rn�"=���"|2T�ƳCV��%
�g�l4!f�	�"-�B*�7Y�'k�'L��{#�'��0������'S�c�$>�)��ة{��ƃ�p>1�jHFy��L�Z�������TI��0����p>���|��?����6q�$� �0<*C�	X��5���Q��-i�&��C�ɚ�n �IG �öBG)�����'T��ѧӤ��O˧>�j9b[�N1<���	d��P��H�3�?���?�fn��?Y�y*�
�ۣ8�����h#V��+��,%�¢BD�=
�����apU�hr�'�!c��h�0��FN�?͔	��!3��E�r"O����$�*�0�l ܠ����'|�Oz؂����A� �r%>�����?O��h ,����	�\�O��պ2�'���'բ<��k�me�l�ѤCZ�L@pP���B�T>#<ѵ�Z2�huq
�'��B&	?]�pU����O�C�ܢeȾy1�#�C�����L16���$:�)��LX&JT�F��P�ĵIi���L*D� Pd��i<��٠��\�*}�A(�P\����ĩ�"kB<G
ϻ@�Q��?���í��C���?���?	W���4��X{�A�s�@�v�L{��A�v�O $Rt�'z>R��L)s�A�$}�T��' $���)��E!r*��v2r'2�C�'ZW?�EA�����I�:L0�u+� #	���Ka�vB䉟ߐ�c�,X5�Rኰ*�-�`���SU�~��ش��ċcQ�������G!L� ��?y���?1##Z��?�������?Q��f���7D��Xd\@��������	����JL2���,���A2eܳQr����	�s�N���O��0�	՘l^e2�FBE����"O*5�F� �+��]��$�}+���"O����a�7L���#�����B7O8��>	&cL�N �V�'�_>��慕8u�| ��.�5XX��٠�f�X�����I.5��	z�S�tg�"f��`+�Eò}��a��(OH��4�S�H��`�-Κ=�D�pf�[�1.أ<!��]ϟ�D��e5#��tX$Mġ	�؀��͊��y�/W�BKl�#5c�8��[�m��0>Ǜx�ӗ;D`U���������F��y"J��S�6��Oz��|:p%ԁ�?)���?�a%I�	��S"='
��J���Lt���嘧��I9.tf5�Ŋ�cI��ǉU�*�X�۰�[j�����(n�]H&��;c��!S�/�r��'�1O?��ŵk&\��b���S�z�ף���!�ğ Q�NiseW4]�2� sHM'<*�T���?���/	�<�X=�q�� 0��Ȫ��Hퟀ��5J�<����쟤�	�����u���y��V�v�^*��
8�����~�n]���>�P�� 8��=h�0b3Ãc?92g�Wx�D��c��w�<ʶ����:g���� g�O��� ����*x��)p����
@�yҲ"Oֹ�'M�K^���pJ�5h	�)��Bd���Buh�B�ۦ����A>9�� �T���3���jg������ϟ��	�0����x�'���	��ܘW�M}�t$!u,S�|y��; c3�O|Y �X�x)㡃	t	��0��hjQ�`�0�O�	��'V�gH�"�D5�"��EF%�`��y�G]�L0+�~�>��!J��y2
���)��Ք|���`*�y!�I��L�I�4�?����	G�aF�ۦ+�&[�J�끎S�5>�I��O����Oy  ��ORc�ʧq��q0�� A�cK�8h��Dy�"ő��b<S�
�}�a D�hB��3T�<AEj�d;ڧ��ͩ��^��k螄}���c�2���H�(��e��"ļ7��X��	��ē^[�i8. ,C�Ƞ��S<���̓h�*;Ժih�'�哛_�P���ϟt�	Il�Y�P,߂*A@|
�.��W_0��6��ܟ(�<��O�@	�MުB�@�[�₳_�\5��l�,#<E��aM����I�iC��h�C2S,����?��y���'���R�Ɂ��Pu��.TX	�4��'���Iƙ3��:�HR�����Č@����U�8�T�s��>0v����ڀr���$�O68�T@J�V����O��d�Ot�;�?�;b���r5�!�I*T�4j'�O��3��'�Ԉ�-2�D��L�^�B��'fNI��J�p��� .6a�ee�=����>���o��l[�%!Y��h���j���b%D��)�Щ/��u*���.o|�1�(@'�HO>�Y����MaV4'Ԩs�>]yxY��f�;�?���?Q��+zh�K���?q�O>����?-<H�;5C\�A$�� �u����ɒ���r����c�8U�D�G��^�^��� aTr��O��Q�l��1PHu�	��Ɓ1�"O8ղ �G!b#���
F�v�	@"OI�N˩�H�;��z�N��;OJa�>�s��.RY���'��S>��@	Q�Rm���8�\Y�@(1c���˟ ���.�����[�S�$kC�"�.�I�L$w^�I4�V�(O�@`�S�HH���S [�"[��+�f�!Fo��<Y��H���E���	1Jj���ī�-`��R��yBς6�|�$�/��I�@�3�0>yB�x��ڝcj<*�M�"���v�T��y⦈,ۖ7�Ot��|������?���?o^&q�n��U�~���q��XX�8�3�ޘ���	4x]�P��Nz�v@r��M��@�%c|�����	��
\ј O���}Gl]3�N);��'�1O?���D�z�D\Ҩ��+'!�䒘SK�@:dهk4�B#��}�8	���?�� ��G��h
e�:xA2�����ɑA�g+Ο��	��\�I��u7�yG!͝j��u��D
����EU��~�J'��>y�B��F&�,�&�J�knN@�r�\f?	s��mx��ᥦ�2x��pC���~*���D岟��Ӈ�O����W�&��y��� "(���%"�0`!�D�<�5�OBZb=4�\�~|�uFz��iU;w�m�<w�B���̊,OJ6ay�aF+R�����$�	ҟ���*���L�I�|�W�?��qB��\�F}�)X1*Nw��� �~Uj���'�:� d�ɤ3TL�Qiʡ���)V��3=���jS��K4�*���T�(��p+�7��O�TB��'K�u�XBeR�5��*X�j$ў�D�`*WR��pqC�8<E�!)Q��y�(�2Et���F*_"/�&�[4Ɩ��y�h�>i.OP���K�Ȧ�����O��Ց2��) t�Y�b$A2����� )��'F"�ĕ$��T>�b�h��Im �p0�T$K56����)�:DG�D�˯^`����(S��l: .���(O����'	�>��6/�&h"`���Q�SM�ٱ�;D�ȁ�)�C(n�5"�&	k7�9�O��&�x�է\�?�eʇH +l->�Q3�{�x�rD&�M;��?),���#��O����O� �#}��@r��\9���u� Ym�$?�|Fx��.04~!���*���1�D y��Qc �)������fq{���:r%�AP0k� k
���u�S��?�td@���9Kw�@�(��%�
m�<� D��
�.��t���P1[��ɕ�HO�"�L�)E�Y�hULL
%��?kW����ݟ|+E'L�Y������0���D]w��wR(mI�@J��|0R����ԁ�'C�K�q�ą���\�`��r��o���Ug�p��	�Q��)y0��$\�X`��!1"�	�c6.��+|O���ܜ	�(� Ƨ�.�֙!C"Ol����+-��@B�ӜS���a�.Ye��������ڦ���ΐ�GMFБ�o�Y�`���\� �Iß����=������'z������l��$m%��ô�ʹ@�J���<�O��J�Q�`�"Č' 3z�!H����A�%�OL��'�\�~T��ϲ{b��[����y2I\�}lV1ɤFܗrC�d�ũ�-�y�
�n����/Xke�캖f��yc>���W�x��ߴ�?����	KtAdh��Hν��T�r.�`	�$�O���OB�P���Opb�ʧ`~��s��;B��5K�$�2T� Dy�c��蟄p3��Q��5:'iׄ+^�8z��I�%���0�'1�4Q��'�\A���ǋo�ɇ�5�X$8��լG�z�B7�˃PUX�����ē��,�U�
~^M�E�^RlϓG4�}a�i�B�'哹6X&��	͟|��<�
�K�ցd���%A��d�p���+��<��O�i�U	�pp�)X���kaH��]�n�8"<E���o�������'�A�cLGj���O.�?�y���'-����W$l:��p��.2�� �	�';�|	p��,,�*�.U�Cj��O�pEzʟ21:e%]��9�ѭE�Tz0���O����3��e�b��O�d�OX�����ӼCW)^,о��6)ܬ!�jђ����R�>AC ƷZ�Mb!���#D���g�'	<�01dZ i9:}��B�<c5��(B�ϒ#C�3�5+E�M�S�����d��Yu*�����.���sD�#=P��TT?����hO�˓D�Hj��	�J�C Wj�v��ȓV�mj)��Sm,���G�ve���B�)�/O�����Y2H�16*�ٰ�mH���ہ���T�IܟT�� �>q����Ḑ=�p��I�8�A냑EiH�wFŰ"v�i(6K2�Od��W��CC�5E�Z|듃�(]��,�Gc1�Oz����'�b�ٲ"Q0]�2N��jT�	�N��y2i]}�1�o^�x�.LJV��yb)��\�d��`)¹h���x���:�y�9�I$-|�u`޴�?������[ D�h�gi(��`����[~n��E$�O���O���&a�O�b�ʧ2� �R��M�+p� ���U-�Gy��ݤ��`P��C���"Î� WX�m@�	�h�D#ڧzn�����uԀkчܔ)W,!�� ����`9i�ʤ�`�&XQ�Y��	���+Մб �c�N�b��&|DM͓��L!V_���	\��ƗNR�'6Z*��T�-�48�! Ab��u��I�q�F_�z�cS��)#��O����N	5z� `V���'b��� X�J�B����Q��<h���ן"~���r�ȡ�V��p���eK�(*�'�ɟ�Sش��)����˓��P� ���g�H�w��2l�8�ȓN����A�MG����K�<A2�Dxҧ9�A&�I*{��XpP��gv"�Ac�-�.}�	͟pI��$]�������	ӟ�I]wNB�'�r���U s�K�B�pW�`��'��)j�+}y!�K�=F������!���~}6����?K�Pq���K0�|hg�V���I:BV�#|O0��5$�,n=L�r�捍j�h�"O��2a燖H�y���,CHt�Cj�R���������0�o�|y����'��`:����˟���П��	�u^��	ʟ��'CU��Iɟ�!Bi�VY����F�`|ԋ��.�O��Y��u�ڝ#��נ�4�j��+�On ���'��I-��7C�!ͼL��Q�y��$^�9�G�2M)܀H�K	�y��0?4`b"�H�J�Q� ��"�y��9�OTh�k�Jl6��C)%6�q��"O���$Bہ5P�tb���ߜ��u"O�X�#���l�gꂆTg�a##"O$u�"j�D��%�OjXu��"Ol\��o��z$�!��ț�jv��C"O�  Ը��		0\���v"^�j�r���"ObL����+C���BE�	E��d��"O0)�s�_�1r��Eώ�H�(��""O�e+ǩV`8��M����!"Oh�q�P� "�L�с ,�t`�W"Or� �%B��>�7� 7�����"O������^���;�.��ށJ�"O��`��E/D,������N��6"OzT�LM�0����했Q�`Y!"O�ը�g�,D��`��2s�R�ڠ"O��9�!DE (�����5y��Ҧ"OP%�Eڂ,� ���I�6{�Rle"O޵���;eu%��M�T�
)P"Orݹ�*�L�F���ꚢL�8��"O��XW�\

O�P��H�|��U"�"O�QB�Xp���H��/m@�9�"O��R��׻F�郱,�{��`�"O �ksJ�R�y��jܖd���;�"ON(�7N�.M�B*�h�)!aP5sE"OT��A�0B�x�%���w� ��"O<�Qʌ,>{TT�G�/q��!��"Obh J�|G���3^�2׮a@�"O0���`�:� �P�$ߞ��"OVxF�{.m:Չ7\&$�jE��?�M�LJ�Ū����pq�ݟk,\5T�8"
�F��x!�X�����<o��	�jR�|�=���`�H cg:u��4���q��]�Obtk6%F.c��\7I���B��|e�
	����eL�&�Ac���d�p��I:e�9,�nD��Jm2��g̓S8�A���!���R �L�9QV��3�C9�~R��"a�̋�Z�0(�i�K�{����@(�/�\�ͅza��� Z8Ib���'��]FyJ~�0":}��`	Ѡ���ё�_�I�����S�.�>-��*C��4��h��j�^�!vO�Q� Su�D���O	CǎͱD�=ml�R&�Z4X�j#?9rd�`�>�kg�YU��0Q����}�@��*M&	b��?d��8�B%�'Lt��X�[�L���?Hls������Ů����"��X���Ũ�q}L�5a�������̉�jG,�?�3�ɗ p��M�V��Ƞ!�>�D|	��<	'��(\{l��'~�@1�X�\��԰�)�37� {5Ȱs����a&\-K��3w�'�EyJ~����/�Mz�L�*H��H֊�=(���ɛ$BT@���'w���V�pY�CB�.lMK3��;}pa{ҍ]�)�ʓ"�xl�v+ˀ.�x���+ϪrÄ�aش��<)e�G�e���H�-R6}�1�?V]�ĳd�*4H���!i�P˓n��u?����+$ A���xp%���#?�3}�`�����ܰ�J2D��a��'�$I��C�/pcP�fɋ��T�C�LPy�S�����T� 3�(��TQ����,�
2
j�,X�D�<��nЏkM��%�P�6L�ʓ�0<�M2bB���Aϊ0A�e2�C�v~BᓾU�q�`��:-v�HEy�'v`V5 � �"T#�D=���E��=Q�C�S�d�T��N��H��dp��S�C6x24I5�l��Q�)Bk�\��P���C�!3SX4���ՠ�X9�+�t�k�~⟘!��R��BG A�k��:b����L{իƃX��1�Ne7�E�Z�bLITe�:45��<��@����� i@&Ef������.@�Ox�ɡ8��LCEI 
���Y�`��.[bVXi��Ьwj�캀`yi�T�$n���?y��8�S�3b���鶩���j���9]�b����*��F�7��`�)��?�b��:��E*��C�-�d�3�[Q���>I�̀��a����FǕD,�B�(�����*ܗZQ�����k	X}J�J�1hY�ᘛw�\A)giV�
BfM:�(��X�B��S����I*1V�D|r�_���x�lY1'�*p��(?Z��Q6
�>!�D�#}D���O��`l�s�����󤄁ZiX�R����0���X�B:+�JF|R#+ʰQ0�Yk�X�'��M�3��;/rl1emڝ'6XY&�ɔ}�~q��*�O��{���4gR8hZ���'H
V���Q"�ɓ��Ė|�R��QD�2iΞ%�����&��biT	4�!9��`܊� Үt���Ĳ���I@�%�$�DA?M�|�$�Y�6.nA��B����E{�O�~hzR�����)��w~� ��iɴ?�j�x�*'ԃR~�!�H��JQ
^H�'�J��]1C�����Ka*zĂ�K�T�0�fJD�ʁ'� L)�`*b��;a4�}�'89�2�Z4�e*]K4��2D��O�DhGy�C�r,Z5�a"M7���6L����d�@���tf </�hT���RU1O�*Ц��U�m�\�	�f������?iU=O� :pJ�]�E��G��~���࣬�$���&H���x��,~JQ�P
�$AG���[��2C����F�ֆK�E2�K_�%,1�'H�,�jl��=�O<��4�z��M�PL�\��'�	�Z�RD��^���$��p���Z��-+�B�I�f-B��m�")��c4RN�&4b�X�(�鼻pb��_��qQ+&q�ȵ��i��R96�1��9O.����V0rp�mԬ\����V� �I�3���qz ��\~�)���~)��H���J<�<�3��j�D��
˨��'zD���0T�e�Y����,�cT$�)��X�̆>+eH�� ���1�6&ЭuKl�V�4<O*���+F�[�)9AN��u���·���Qv��Sk��Y�gYe�'�Lp�	G]6N���� \=>Y���':l���M�A8�I,"�.�`ǉ�3g
歑�E|iL� ��"}"!ƫ^x�'N�Y�'�L�]�XpK�F�bT�,8�!4I�ޓO�-:�)	s�b>�${��(�����P�會|�y���u�bH�L>���>�L��ug�yc�#���?'렍�7oϦ�6�b���4I�
�q�*}�l�O\5�cl�q|�����Ć��d2�<�9�+��p;� pe�Ei�jAb[�����S�rI�S�'x��ҎE�)d(������x�TP� �OH�#�	�&��QI�;���*�q"�^�iE���IŘo���c�'��k�j�U��#�]�
�}!�Ɠ�P/.h�Eh�M6�d`�/�<�$A�e�4�ږ�=}�A2}�'�7�<\��g]�2	t軐���b��8�P�(�$M9WE��s���Ku�	S.�.=��d��H���%�p5Vߎv�d	�Ɔp�tSN�@�N���� H<�ڈ%?7���J��j%/�|@����{��I� �ُr���3	Ā�0<љw��@�FbȂ;�f���A+%(�u �Oݳ2W_�Z(C�HSd�bW��\��%��o_+6� +��I-'�p$Q���=-�O/���p��=3U�| 0�N#��(��'w�U����4{`}@��7y0�3'd��d��!��l��҆�!��<�슓u�Irj4}Z��*n�[�H��@ �6��k���P��	��yWxI�j�7R��+�(\���>I�ʗ�_���`M�V�@ AJJ�d,|�$��-�D���8��@�KV�b>93�\?8�����+ϕ�Z�MOL�2��O�����Z�	is�'�󎈆JP%�@dΉ  3�)�,53�I�T�O��J�	s2�P7���ΈO"���e��@��<Zv�C�{1[($?y��Dg�ɠ/��{4�U�f䤟�`!K�2s���Kd�H�; �ت%�621�(1���7	,�tt��]5,��U(�ꆋDF�U�D��G�Dʓ[��R!�3������gDU����/���D��F�8��+9e���r���2y�VQ[��`���<.���t�D5P.����4��6��\�F�9l�4���m�0q�����~
��O�P��J^6���r!#��Xj%��'5x-���+]A|�ғ�d���W��ؘ��f����WZ���u���1|�lYs�t|�2!�.\/:y�/߶ug��Bï�SRQ����^#">4p��D��9U�;po���v�!hP�ϫ.�7�Nb�>50D�@��ɽ1�<�Ԁ�p���!BDħ	NL���ï ��yBL�G}��F'^�u��˞�nM0q����U2aEM�ٱu��I�ހSW�^y��L�A'��9LYSǊĆ{�\1i�m�"Jb������<)ge� N�b����F,Hm�.��W�Y�0�IFLԍ��aR�z�V�0`�f����d��J���}B��F�e3��4 ^'?����֋�C�;����҃�#oneX2ˊ>��t�W�ϟ�S3*�H�	aKZt�6-����
(�"5�=��g�
���'��|��l�`�lM[�jV"(���ߧIJVQ
�Ɣ(f$��	Q,�?�Ϙ'�4��[�_��tl>z0
b�[�``���6,i�@�5!ޱJ��q��J��l��.�O��pH ظ��	�"*@��w<Y84�v-��s���$z�tH�~��)E#���ԋ8ɮ�ӗ��]-�Ź`e"�$Q/;Z�w��$Vz�#/�55z��>�'`�8:o �`kӊS���z�o�u�'����rG�b�Oq� .��|���b��@6�\]�/�/r`B�ɳ"�h
eQ���5_qџ�(�HD�+���R�GX��X` @�"D��v�ԟ��d�����p��� C���DHx�A��_�R�$������NE҄�7�O*���$Q�9�p�u�,6L���=O���'���f��.<]*���\>7����	D����Z6 H�l)�Β��0>Ao[4��ɚ�"��`�׮Tf�7Aߢ4����'�H6z�Ha�S���ȘIz�%z!ȣ��W��S �� X=Gx��'��D��DY��@2�S&!�~5B��0j���)d�:df�GTo:�bH�X�џx@'�̈́}3H�#РG�Af���H�'4"�M�3��:j�����c5��n��Y��%��ύ�鑤i7(��	H�L���*3�1_ B�	�i���o�>����'�$?���z���ˊhy�i��'�)���i�~����/�f��矴3ҜM�*��g �8�g��p=I$�'@���C匼;^����ֿ5:e:"�X��8w�	Y?�!���!蛬3W�����Ɵ���J�0S��1O���Z�NX�}�1O�X�FH�=6�e
7��+y;�x�����'��y�j�!^�5		�\ӊ�� J�g.���)� V��&�n �=:t�d�4���`E+)�x� ���'�CG���i\ yp��CHbiq�O�#&N;A�@,O���y&"OȠK ��m>�,ˁ�� ��-�ƃ�$H���iy0��`�e���C��O�-ɇ	��@K(,��'�\���N�6�	�G�k7f�����'͕[�^u(C�q�j�u�L1�"���P�JY�L���07H�`t��-�4�>����?U���1E�q�����k�n̓1����c�y���P��Y-}����Dp���4F~؜3�Z�i�l��W��jl�"�ݩq㬴�
�Ex�,؀+ɭU�<\��R�w��SXO�6�Itg�o�"ūRh���G�+�x�-Vź�gDm޽�G+Ŋ]?J�:���i����)*D���#11���Y63$Yz!�� ��1PwH ��e2E��7B��sQD�օLA�b�p?-2�.�Tn�$�ia`Ǉb|���D���ѣ]�l�V�Q04�2C��Ӣ#��e/��(�B�"�d�:,86�M�v2��V�I@�'�l ��6�$��%� �<ʍ��ΡX�| ��l�l%��-� H��=��� X���bf�t�@􈶆ʾ~N�p�p�Y�l���I1L����L�?�~-9@��*c���D�
�xD�9���ϢC���0��N�����D�3_~,o�~��_jl QE@Q�lU" AW�@]$C�I�d�1J�|�JӁ��o�`EJ2�3D�Չs�|�'i�ԋw��]Xz!�bf�q��L$D������Ől�B"�OJ42��(I$� �N^+x)X'N�	ܘ�Yb-<��d��$qan��lp����*�Q��(�FѲ*ڜ�� �C:R,H�P�%"�1V2�hN��jZ���$�S�H�R�-R�r��@�|d�rC��u��e�ܞK4`���H�
w�|b.�1:���R%눙e4�-ۇD�4��<��)�+2��[B�˒=�D�Kg&�z���<I�wHP�a��#d�� i%Ɍ*� E�	�'S�x��#�8M���2����7�7
�j@E��;#�.�M�'B(Q�ę?�]
�$e�c�A9P��'Ƅ�W�C��:zs�Pxt�9H�)�!��c�6��3�Gg��Q�L���B(9�b�?=DzB-��^���k1�N2."�ʁ�>�'(�#od����-N�ı&*�#���Y4@�!�$�8UN��L�;��mO��}������j��>Q�� f��Q �&G� :r����1D������=N�U%�c�Z]S�"d�����������vJ�%Ȏ��A�ޭ��i��Ά�y�#\2@��"��ZO� ���Ě ^�h��Ğ���։V.E7`����X��!��H��!�g�I�J���9I�!�d��
�ȹ��ˏWGDh+DI;A!�$�� ����
�;I�<�ႛ�"!��1>�.-)1Y�c���a%0!��ԞE���!�ݑ8L��bA��!�D�X_~�pB*ݮ^�4Q���O��!��c��a��KIE(Ea��d�B䉵H����X3��d�up�C�	r:�07*@�+p�I儏z�C�	�Z�l�٠�E:h|^�! ��5�B�Is4����D[r����5I�\B�ɾ�I��%H�p�N|�� �[�C��3]�I�D�K��S=]�B�ɐ��xb�i-�0�+���#rw�B��5ZN�m؃,�c���LJ
׆B�	�
�mp�Rf� MXc�ƍ5��C�-*PX]J��ٰD�ʬ� �~�TB�	��p,�BRc��-�c?B�ZC�	�D�PY�$� 8�A_(%�C��1.nb���lK$AC���p�ݍB&C�	) T�e"��DLơbc�<$C�+>�
2��~��U!�g�3A�$B�I����2Ɔ�kxE�va�mH.B�9�^�X��ZՅV�K׸B�IS���i���=L�6!ȄK�C�ɼSO��hri
�!�.�	���~[B�ɉ3؜-���C�l�%3��
B�I����s#U�ExܽX�g��>C�ɼ�0����u�������B�C��2�@łq�R�G���ڷ���C�)� �@��%R�d��G͞�@��,*%"O�\����(Ί����\: ��"O�%�!�[�1`�E���Չ8�h|��"O�P����_Fz��`�2���� "O�M��M�S�����D�[%� �"O��"�G'�<�B��6�r&"O��:@��"��<#b���F�9f"O8�е�R㮭Q��cw�i�"ON	7JXpt��o�6]��͓�"OJ�K����h�!D��"OTUS6I^P agg�)����"O$�+�R+*�) T	I?~�,8V"O�8 иIZ��uH3�����"O�I��@?t�)p'A�l��l�a"O\�b���C�b�JE��8p`�h"O��J"Ǵt�bϊ,#�n�S"O�a��	�wR��Ӵ�L=t�~�ڲ"O4�TK\�L-`a`�ϐ78}x���"O:`ӂ��uĸr&iM�Os�q�v"O qA�W�E����9C���}�ȓQ���z�2y?��)�O���D4���2����L0�r�Vc\5,��wx�E��ґC�P���02��!3v Ye`H-]FJ�/�5Q����� �hhB���H����]�|~�Y��J����!�	~�ja�$!*Q}�݄ȓc���I��Ԑj �8��"?�5�ȓH
]�Ĕ�J�t�kWK��)ü���v��\�f� 9,�e㧭����$��NL�p ��E�� 3o��{��}��S����fy�̇^E�Ш�i�3����֭5D��1aW/HO $ӔAô� �2�4D��y"Ė&C�`�5��M>y���.D�\���9�i;���y���ѣ�,D�Ҵ�R9I�P��@�Q�G�]��m,D���w��=*�5T(�?D�d��I&<OV#<����K��!����X�0��'=T����
�k��y*� M�8����6D�x�G�/ �*IkS�H���<j7�'D��������k�NpSP )D��J[ `��1�C_f�l�qDF%D��"�-�(w*�ci9N�48;�Ɓ��hO?�d�
~��CW:.�n��B��k�!�D�O��F�%��J�폠A,��`��iH<9P�C�|���68��Ո���a�<g�ZT��P��jK2^�F����]�<a���J��z��.�ܕ��@�\�>���Ex����B�oSV$�gl�X84ѡ���y"Ɇ�1����>I�Q�2���0=	O��h�'���Rv�ß�>��M�!,�Lԓ
�'Q�]���Ӳ>�p���L�*)�٩	�'��u˶��5#P�!{ .�(��)�ϓ�O��g�'������%���Q�G{��	F"q�j�'HP�bp|Q*�b�L�!�d��oز��p��+�v9a0�]�x�!�d�!�,(���h�����ǎ<����i$x�;�Cߟ1^<b�e�K��۔H/lO➜���:P�I�!������
*D�,{w�H4R��Pe�'&P!�#��^�����h�Z5Zu"�4A��`��%e��C��<<��ꈰ-eD0���rBB��V9�I� :�������%A�>ʓ�M3d�2|Op��`ႋȦQ���~!���'����&'��as�Zmz���v(�5t!��O� �1+T�'�b���
y��P���Ii�O��	��,
f|�M��. v�II>A��9�S�S����kW�Ov�{&*L�K�X�aP�#D�`0A&��Pؐx�+	*�H�iSL#��<���]xRre��� ���w�H�<	p����L�i�|�}�%_z�<��o���}@�)�	P�T!8��s�<y�Б'`���r'��+1K^m�<�Sl�cp� Z+�	NArQ�ri�e�<'�<XA��(�CΊ04t�S"J�5l�J�����V�6SE����P梄��y"�&ֲ��FB"z1�96(�/�y"�T,!�T��K�y�h��ˆ��yr����pC�#9r�0���E3}�"C��9�ژ�aDX�#�f���e�:F��d1�tY�����;P�8"�9df�ȓ*Ep\i� Ͽ+��%j�EW1dw����r?��
�4|A��a%O�Vx�t�ȓL��(t���^<��y`���w���<ߓ[Ī0H�Y��"
+D��i�ȓ����d�72��	  H�S�r��ȓFnd��*S�l�N�97%�>"�Pم�	0Px��ɾ|61���Z�\�G��Tc
l(��%_N�T��!T��C�Ikeh	goW
oPJ�H��V�h��B䉶�����X�fX`HyS�>.�B��;�А�%��w�13��[����LF�9Opd�%_�)��Y�n�^���s�"OP�R�(i��9�c̤������Oأ=E�Ԩ�<gc��a��1e6ph��hā�y2Jc��s��C�P��aZu4�y�a�HN���)Os^|"�ҭ�y��@,h$KDDȲE ��Btbۊ�y¦ϔa��e�8h=r�:5fҐ	!ў"~�B�ֵ8ԣC6�}��E��H��ȓ8OD4JS�Z0-��Ȧ%2���S�i#�������e�P"�X4��A"A!��04x�s3�Xפ�sP�K�\�!�DO�~\"��� �8d/>)���8��=E��'�Y{$�ݲFmJ̙�	�W���'/��4�G+}R�`��I�	���$'O�h@�i�.S�&<	�W5���I�"O~��S�>�� �g��{���#�"O"�ڰ#+$���
����E�"OL�KǺ}���3 eJ88��u�@"O,�A�Ì�A��1�B��|$Jp�"O�A�+C
$,��r�F�ȅ"OʁC��a[��� )��1[`"O��wdQ�!��L��(�0���"O����ùE�la���$#ո1A�"O\|�����[��A�K��5҃"OdM��G�B�$�I��J]R�:�"O"}*��Q�zD\h� oA/M=ΰ�W"O
�A�����P�2`	1]�%""O��í�<fh���rH~�"O�DY�,0J�,���΍j��("�"OX%"C�]�ݜٳ��Q� )FI�`"O�M2��F�S\Լ8wH��9�b�"O�tp�ΊX�A���\ P�"O"�r��R�'-�p�@(�x�s"Ou3�ȦM�@�q�L͹���"O�I���+��9�J�$"t�P��'z�$ғvҘ�p�<+��6_e!�$No�|9�'%_s�Vh(�j =O!�� ���Ƨ�m{��9!�V9!9���$"O!
&��'2���}�5�d/\O��bج�R\�F�@�VJ�b�"Oά��-9�.�qQg�BY��"O��Y��R�.\��'-�)`xnD�2�'��O��"�*]�u���u�Z�f:Q)�"O p��KU/&�`���+��=� "O@t���M]j�2`lL?&n]Z�'f���u��Gh̿hv�8�BD��-�"<iϓn~B�R䄏;���̓�}�P�ȓ>�0�㲦��[� A�Q6*7 �ȓD�p�@;��T�
1[�]���Hd8�)�Cfz[%��i���ȓTA��[ɢ ��x�����=��S4¼b2��.o��x���<L�����B�\���H��$�4�����51`�ȓO����F���H!*!�(f�dE|R�S�K`�W@�鸭�$��{��u��U�;�B�1'�fp[WD�.��H�ȓ2���S#i����b�A@�&m(���}��@��՞qw�SkR;	
X��ȓ�L���#H��0�C���o�0�ȓSy"�{��T�p۔�C*�fxE�ȓY���Z�)6O�:�$��3L�m��O�JP4MO�T8B�ha��Y\���t�~����ƞp`��5�P.r!<��\���$�:S�=p,ڭ!��,�ȓv��i��V�h�N���U+k�4m��C�"�ْ)B4����D'd �ȓQ[�y[%��z�j$�t���f�rѴ�������'ؗ&0�݆ȓ	Vд�T�	Kj�|��n�S0��ȓ$��!�ǂ�Z���C�.ՠ$ڊ]��g�ԙi��>	|I3R��8Βu�ȓ$R՚�`׺&�:HSq,�8��ȓFO�0�`��@ +��n"}��]���i@�X��.e�w�/�ԆȓP���W�X9JSTXW� A�
E���q
�@y�Ы'銝<h�ȓ^���g�H�f�ӂ�ƲJ�|��ȓ%U8�@.��9ᘕ��B�[i,���G"x��'���/]�}Pt�׉����ȓQ�Ib4�\�d��YP�M�1@�������9! 'ƛ1��	�KV,F����kN�����
�*d�6Ɨ<f��i��q�M�+Rp��Bf�K!K�<�ȓ��]j��2	qh��͕ e�\�ȓc���1)�G�Z$	 ���C�����D	�C�7;��a�H���,�ȓ[�T�i�NK�$��H���Zk@���N}�Ͳ��B�d@�Ŋ@�{R�0�ȓ[Z�� �L9T6� ���]*C�$i��Z�z8 R��2 �R�U����=�hؚ���� �n]4G�>a��I�����s��5{ՂM3ANP�ȓ �$�6&�6p4��UO�.Y��ȓQ��L�Q���S�$���cJ�7\[�ȓ3�����G��,�ac,�J��o]Ċ�!^�	�q�I�+^fE��'�hkŦH�+�*�1�dƳN|j������3�*��e�xU!�KN�<�&���f���eb	��x� �O��4IJ��ȓd�T�2���(�l2ӈ'$A�P��n�"t��m�`����d�E$SH8M��S�? ��Ģ�`J�0$�E?���"O��	E뀛e�N�*Qf�Y��-�"OLq�קu�L�VB�5��41�"Ojy�c-�.mҹ�#��u�l�p"O)�)U��H���"&f�"O-YR#����lP�I]�.Q��s"Or��T��.P�I���W�@d�"ObX�q��9 ߢLy��� <�U��"O�9 ���kf����i�/�ё"O�[%��8.�
u�. D��qP"O�)z�bzxHl�q�F�89��"OfCӋ�=�PAHfmN4B)�TR�'�z��#�ɮ6��h��iYx�qC	�'Xt��Kɽ�2����~9�<��'��Q�tK4}��)h���mo�� �'R��I�n�I�y�>g��� �'8��@�%��M�E�ʅv��y3
�'� ċS�"N������j�c�'V��Xt�;Zxd��!&	2'��K�'��R#N�C��IBQ-�6�N(��'l�x��i�����"UC���2�'7	��^(L��Ē���<�$(�'x�����pV0����/���'�f�F��u-Ysa��t/�И�'�>xx@ڀ$}P)� ʎ(q4�)�'&|��q��$E��YÅ�-d��(��'D�l�B�̫t�ȹ!�ھ��%A
�'4!b��}�d���.	g8k	�'���[�ˇCw8XBU��' �T�#S�L.�,��޵f�P���'�6����[8��Ihvh�%��'��`+ �?/��y��gAp��5q�'@8	�����//N]�y�|qQ�'v=������I�<o���'��aI�O�%��� �h��c����'��k ��h�0 k§J���x
�'�<������<z���1a��'�tѥ�ʀw+�=RPŕ�|qJtP�'��h	�#�U8\�7`K�w�Ъ�'I0:�e\�eqz}�g$пv�V�@�'����Dة Ȥ�膡L/{��i��'�v��6��%
y7蓷?��k�'!TI�t^���v.H1����'Jq���I�BX\Z�ܦ%��y�'6�'` g�l�aB��
����
�'����d�0�4�0�����h�'��l*ŏ�,�Z2�`�N�1�'o�T:�/��I,��рe�?���A
�'�raӖ$P��v��-ЂU
�'�.���h� O�� q��������	�'��9ru�[��b�"Um�3���	�'���`�d��~�� ��U�
�V���':�3�%�>��I7K�0	,`�'_ �+��+a0���)D�s�Q��'�D$��ZS�P[����jɒ�0�'|�M[�냋,��h�cύa��q��'�Θ������cD蟅R`��'��`�w)�6N�\k#(Q�V���'���`��� C
V<P[,�	�'A��*�d�N3�oܙW�ʵ(	�'5�5�gB-"c�eЄ�� �*MK�'=��1�*a��$��u \U��'-,�cgb̗{+yj4��u~-S�'��pC�]"%�Q��^$X�q,D�� �mK"�A�:jD��G��b�j@Ȥ"O���v���M�������C�4		�"O���B&3�ݨ@A��!KN���"O����(3޴a���8S+FM�"O�|2Ah��80��#NL�' ���"On8�&��-��� Ն��X� ��4"Ob�ȼ,A�(p�����"O�A"�
���գLJ����"O��#)a�@�T�Y�4����"O�Q�t�S�fX`�$M
]:� �W"O���,
M�D9ࠬS,�\�7"O}1"��*\$Z�B��I�Fl�1"O���R�,9�V90ؓ4��`"Ov��gg����d�6-Z���ٵ"O��H�f�aFę� �
-�:��1"O�1�E�S�& *S�t��(�"O��#6C̅P��
RMB�cyn1ce"O@�+U,�<�hA�G�̂ag�Y��"O��P,F�*�l�X�n��L�"��"O��"�v���5+�$,��A�"Oxxs�$����S={C�k�����y"�G�u省���������u�(D�yQ/<1�:a��"��+���f)D�06ּb����h۝l���锁+D���F�Zi�=�cX2<Ux��"(D�$P�f;z�A[�eT2v�f���%D��C�"P�S܍��G�7	m�1*Ol]�#L�6��p����_Lf�*�"O�P��d��Bq��Z�%EEF�izE"O����"��:e��H
�9*0Lt�%"OD�z%�Ȃ]i� :��F�>;+�"O2�Q�,�(x��� 25�!b"Oz�c��I�&ᐙ"f��	���pe"O,��⪔3-�`���e��V��Qq3"O$X@�g�
���Hs��v)N�:�"O­���&F�"7��a��$��"Oh$0�������@-W����"O���/H���`2`�3^M ���"O.���3jEᡮY3�� B"O����-��#�,k��,I^�ա$"O�Q�PC�@�R�O�:n� Ҧ"O)J�`�D�YzЍBG�����"O�ɲ�Q<0�($�sN�%+H���"O�t0��,�@ݪ@��
A.��S"OF Z�l���H�u�߬4�ͻ�"O| Ca� �{T!��j�B� R"O�����Q�t��2F�8 �w"O�Ճ�f��OO�݀��V�@ *�"O
y2���W�p��f�P;R9��"O�(�BK�_����Hň
$L���"O��sq�B�q�IX��̃`��"O�x�a�E�@�G���&�Qp"O0�+U,�Y�p��Ӌ璕s"O�I���Y*D�Fh �O9?N���"O,Ec���nz��c��9Y����"OI�V���N��aJ��:-��"Ov\ S�7n��Z#��"O;<dx"O�a�Z&ݚ�J"��#q��la"OF�����OW�����%�­
p"O�M �+��B��Z&�)�D"O晐�
z0�
��Ӿ.��ys"O:�(���Q��JuI_�0{6�!2"Ohu;�)��\�'�˱Sq
L`�"O(	Q��Ӗ�X`<(��"O� �i��C9r�a�`������"O�s��W���2����"O`�qa @�2�(�ڂ�7�d�"O$,@Տ�F[؜�F
Ŵi�:�)!"OX�i"�C'/% �Y£J@.�Y8c"O2�&	)��1�t�5���"O �P� ��d�B�#l��UX$"O4Ű�G(_.bDBϧQ�8e�@"O`}�a��0���U
P�V-�U��"O��Y��������c��<��"O^�:�-ΓTt���������B@"O$��AK�*:�T���M5���3�"O<9��Ă�q�r|YEy?�]1�"O���b��[��5Yg�?3!b,)�"OL��L�%�T���	��I�g"O�u��E'�t�
���1+x�"O�(���Q(F�a�w
�|��`"Oq�����H�ǻm���"O��a�߾{���� p��-� �'*!���w�N�������R��'���!�Ծ,C.h��b�k\Ľ9A�X�1�!�d�;q`1hUI�1?�D����+!�d=}�	C�ڳQ�����Z�3�!�$1M�T)��Dy҄D!IK�!�$\#G��ɨ��F+=�����ҽ!��H%3!��_�F��6�\�!��
��)� �ܨ��ݸ۔^!�$P�z��b�䗯'f�a��ܸu	!�V {n��kfT+v,���.�!�ՇY~��Ԉ�#]lz�鏵J�!�	8m/�� �_�$q��F���!��4aF������z�*�#�^s'!�$��XD�u���
Ӫ�z��ʹu	!�D܉TRn�"D�L2����$�!!�$ *9@��`cj��M{f��-!�!�$��X��)C��Y�ב�!��7K��c�LH�$=��C7���&!�D���<�A��F2�B�. �!�33���0o��f�U�A`ݱ
�!�D�<@�Z�`@)͑5 5`,�!��0YE<���Ճ2� @��x��'�ў�>�B��w�
���DQN�@P H�<i	�K���C�$7<v��S)	gl	��3OLA�M]�u�v4{�h2�ʭ����C� [3��
%-R����ȓkQ���p%�����Bú�I�JBf�<a�C���AA��!���B��
|�<��L�$$U�9��;+@�
d�m�<�Ӭס\�T�@C�����"�i�<q���5<~`�Nj�r�c/A�<�d�/�T�ِ�@=>d𤤃~�<��Y�6������΄��u%�E�<BAk�$�KÂK����2��J�<q��G<yՀ�B�	�E�Q��<�7��$|��4�ژ#mTQ���T�<�¡2B�e�#.�,�~i nR�<��h�*C %0�␧�4Rt&PM�<��L�1I>�#���
�p��E�]C�<Ѳ�J?Qui
ҋ�=�"����RC�<�3h��u��Q�SC;�UHS+�|�<��킓z�5��"ǊZ`�B�k�b�<�e�ȴ	�>�	W�P����A*8���{I����k��\�H!X�k]�;D\I��+���{�h>N�y�%W)O_6���S�? �x��V�v���X�E�<�J �&"O�=z��2s��z�D�-�P�2"O���!B�쌲 �I�W�ȅ�"OJd�+և z��u��b��W"O�ɲghМ*�p�6��YZܻC"O�̑�O�$:BH(���)`92�"O�`9s�T�%�r�P��{�|��"O�t�g�j�"d�A4��P�Q"O�d�sb�-n��,1b�D7���"O���jO	�6t��cM�Kx9jg�k�0�'�!(�ڐH�q*���1D�PZT�ˉ^�t1��$c�&LADe:D�|��F3rL�9���RHɁC�6D�4�3dX/^&��7�	r,BeB��5D��b�C�tlUq�N��m ���Ѣ!D�h��戩&Μ:�g/~�TcG�+D�<ЄO�,�i"U�ϒh��X2�+.��Z���,�:~mB�(��X���g@*D�h���{0��I�"��b�$D�qB�ʈcD!� .(���y��5D�P��
!��1��"�)���;E .D����oU�bv)ۓ�^fＵPV�*D���rd[�*:�\��3�{`'*D�C0/J���B� �;�Dp"�(��K���ӐWF��GEӝ ��HZi'W$B�	�n~.��eI=m�@SŢ�(!�.C�I��ܢ��ʸK�~��7���&aC�I�{ ���ulԢ/9��
��E >C��R�6�3�hȼ;GhIq�´d� C�I>(扁2/9f����'�q C�!	�iW��݊X��dȝ��C�	�nZ���w��L�ʅ9v4
��B�	�n���c4+�pyte�bA7X�|��db���dH�� �fCT(_%�� �$D�KčN�{�X�  �Ҭ~A!�F�>D�0�t�_�q� X�@0����7D�@qS@�s�Ar�	R0g�̕��N D�L0�Q9I�Q
��ko���3D���$�V�X:L�GG�#,8��W2D�kwY**fn�j�
��:a���%D�ܙqh�>'0����BJYLLK��"D�@���� O4���T�ItL"D��i��0�ص!t�R(�#�k3D�l�� 4Ѐ@&��_騜�M2D�Ԛfc ��@���>Rk�$C�B&D����b�&x�ei���7S��Y�$4��Sm�*���~ 3��J0�B�I`w@q���cZ,�CV+
�]ʠC�ɨ	�v��e���Rm�is��V&B�+l�Fͳ AA8��b���|B��&~F�� A�'jR=(�#òP'�C�	9'�>�0ń�^�(db˒��C��S����.XF@�9R���hC�	SӲ�3"��9����B��8C�I�S�PRE�X�V�h ;�V*�!�$�;c�>��J����k� wq!��spʌ��J���M0�/�7`U!���s���E䄍3�*��띝I�!��ͬ^T
�+��0 ���aQ��U�!��S&��т���Z6�����k�!�#'22�UL�� �TI>Y�!�$V�T��2"�@���]	V�O)p!�Atf-R���y�"y��	�LU!�d��c�(����{�(L@���HQ!�� (��GF_�"2J�{���0ID"OXp����G@r���6-�x�"O&-�B�E�J �O���lI�"Ov��tC\�P�W�U=P�n�8R"O�1[bf�gz2��wL�?����@"O°Ӕ	�+n���	 P�xU�"O��Dn>a2d��H�R"O�q@��c��$�#,�(�"OA( �&h����мR�"O�h�w���w4��hڜ_����� D� #ZN���I�m�`͜ Q�
?D���4b��tm^��u\�D+��/D����g��`�z�(�Y8Zb�ե.D�@�2a¾R
�a�G�X{�H���(D�@+�,G� 	,��ÊW3v�jB�B�	�.X�I�F[�A(@�@B�5^� B�ɜU��}�q�½|� �.�:I�C䉔j����P��+w�9�&�-q��C�)?�!2�m�\��+��\Z�C䉚�J���˒� aJ/hC�ɰJ<��2�IJ"򢨺s��15ijC�!Cj(9	$�DCc�8�Ԏ��|xRC��� �慬@�P8�$X�<C�I1n��MB�o�7h��i6O��|L,C�	
q��6��T 2�PJjC�I~�(��t@�F��(զ�\BC��+u(�|��BǢ=���is�\�:7�B�� �UH\%u⢘��G�}�LB�I�/�P�{�*�
 >$��#�>Iz�B�	�?W2�!Q<����#O:E��B�	�tZ�H���$�%�*9���"OF�*�D��[ܡ��C�65ƁX"O̤��F:Q��8 5G�)�H�W"O:Ya���r������(�r�)�"O���G�աM���ѳD�M���"O�R'�	�1Hi�gD׊�"a9b"O2D;��D��Di��2L�>��7"O��H�FY�6�`��
�Ah:�B�"O>�L���h��dց����"O��K��>.�T��Ɍ-h$+�"O�ᘁ脽w�Z��cl�)\�����"Oƴc��X�Sp��@�K�6���4"OV)�w�-t���k%
_"B�u�"O:���f�q0�y�s(�
w�>�2!"O���@�2$�(�Y �0�4"O��J.\ ���D����d"O�Z��	{�&�x桅�A��Ԓ�"O���F¡i��4iE�	o{@�I""O���g�6?�x����<^D�t"ONq�`F,2��L�Sl?4O`��"O�ajB(9-J�TC1B��A"O�ȉ'�K�H�򠇺i(���"O�P�$��b1��3���i���K�"O�%qF!�7A�p q�@V�E�%�"O��R�HK�m�<B5��^ϸ�t"O���7l���~�R�n�%����t"O8l:A��;���Ydڥ/��ɢ"OT]b�f@�U��J��PiƄtB0"O�<!aރ=;T}@P�[�j��$�"O������hCF�W�C0��X�"O�t�⍉!{ⶅs3e�5r,����"OLQ�n�;ҹS��U:gtA�"O���f��������C��Ej "O���C�,�@Kk����=16"O� ��I�"F�b��<��
O7E� ��"Or��⨟�2�8�JB��� |���"O�I9u�h,j�ڔkNH� "OLy���5v�L)Q��ښYQ�P�`"O�$�i�-K.tah>yI:���"O�}�	�a�,`�'��$5 ��"OxMa(��y8P#p��3k��t1�"O4����=WCT�[�Ǘ$��e��"O��;#��(4D���N�	�EQ"O�@r�L��`�#�e�SV,8s"O���-��Ou~��֓/#��C"OҘ*�斺6r��	#~<����"O8����ܔ{�Bc���~|���"OFX*��h������r"O�@󣋜;���	3�٨��C"O}� ���l9Վ��J�ZU�R"OX�'Oɖ:�X� ��M�u�j\z "O���Ð<~�	F�� �2�H�"O$�� ��7P��B�R���գC"OL1�f��)B�-�E�4*`�l*�"O���A�$�{rmI�c&dh�e"O�Ԓ��ߡ;m���,B�����"O��� 
T)D��L�����!"O �kR������[��Mr�"OH�Ф�Ά8�D E/
bB
��"OfA
Q�H���E0 =�ِ"O���X�~��� -֠2��"Ot��.�Vߘ�rf��6���u"O���3�Q2%�k����
��+�"Ov��㯀5<[�a�#B%kX�c`"OX����>3a�4h���"O��`aV&G�|!�LU/!��H"O:d�4��2W�d��- �4���"O�%��#A�d�ڠ�%L� ��Q"O���4�L:xL�ĊHJ�J|�"O.��Z�A(���jC=5���Ѐ"O0�����e6�JgDף����D"O�<چ[=D~у��F�]�|� "O�T2P���Vڊ�3�ɻYA⭒!"O���fG��u2p��w�͈]
8A�Q"O�yb�e$&@@�
��M+�"ON�ڷ���y>���(=g���+��'y��ĕ6�HT�$N�+[k���c
�x>!�dLR�T�skT�Z����F/�!���:��EA��D�!�vy(��^'!��U�x�\qFfP*[{Lq1��B�!��\2_���v�[��`.܏f�!�G�$բ`ҶM]�pv�M#7MݯM�!�d�5RUb:#˝�X]�CRI��!�D�,�z5y�n�)H�@c��b�!���`���j��m6�,�$�^�8�!��K�|�����Ct��3��!��0��5�6$G
=�f���-9 	!�$�����5�+k�؀(�n�"~�!�$ܪw^�赮޺H"���ggV�)�!�$ތ?t��o�?)?�U��4n��	v���@p�B�Lh\�X%E� ���c$d%D�d1�A��$M��a\�f|9��!D���AL��dP��pH�P@�Y�%l2D�@+n��.���ѡ�9&�9�.D���s��;��u06)�#S$�Wo+D���V
ÐG�0�@���0x~4�R@d&D����]�338�:a���Ku�03�D#D�� Dd�a���H���l�g	 D�� ��`U�M�⑘Ӊ1*x�9�"O�H�6�R�/�tH��H�t����p"O�	��c3Zc�G�3_w�8"O`�p5�L�k`��H7���3u���e"O�i��I�x�2���Y(Fc�XP"On\b�E
�!6�k�mC�&h��ӑ"ON)h�Zy�0��l���Vt�0"O�yDA� x�`��@-)��YU"O0T)�U�쮘��K�q�NPҐ"Od �a,P`�)Х���A�X̀�"O|);��9b���l߲���p�"O ��	An�B9x�5I����w"O����4W��8�����n�j�CP"Oz�9��Φ8@��X���U!�qY�"O����Վ- |�����8!����"Of�XR�@�v�
 	���;!d���'c���S)j��m� =�|,J�� ��a�ȓ9b�J"�H3]a��KչsȢ���g��]�E�	<���C�
�p�!��'O<�"��)F��Y�$�6f�"<	�'2�l� ���2P�2/�3g�J!
�'A��U�Z:���������
�'�X���K�{t2��ԢP%��p���&O�y����K��Yb	���%B"O�M���4y��x��}�Y�"OZ��3���- ��*��Mz�"O�is�<-@�`���3�r8{VS����I2�N��p��2qnؘ;��ڲ!��B�I�&�2�㉜�(�e��^�m��B�	�v�8��$���^�A�P4����O֒OT�}�k��p�#�Y����G�&�X��l���[�O�$�ȕ��I p�P������8wo�5�ݙ��HJ:���C���4鈉[��L��E
�j�:i�ȓ+j:9����:�Qz���,S�0��\��h��DµA��a��!z|<�怊�|�!�䃌=�m�'#�^u��G�_��!��[=n,�(oO��b�M�8	Z!�?2qft����8��c2�ʥs�!���@��8�ÞC~�SB�
t�!�$V�qDY	��68q:�Ń�{�!�}˨�@Uf��C]��Yǂ!)�R�)�ei��jw�Ϝ'���H '>8��'2>:����y
m0��FʒX�'������Ot�b��`Ņ�cV��'�r;	�z���G +{Y��'���P�d� �Ұ��C�#��Y�'1���W`�:{$	*s��q���
�':Ɣh��>Ms�h�G�
�eI4��
�'xH\�2\�Yf�-�W��&_�X0

�'|���KZY����
���Y��'�Z8�Р��	$,�)eb�� ���'A���`G�/���'��	1i�k�'$ 0ó�(y,����o�%�%h	�'5@,KM�'��^�+Ӣ����ɑ�y��4
��sF��![Z�m�K���y�-p)���u��Iఋ��y��@�zp���,�y��r jܬ�y$�n�>ś#��r^���7�^"�yr��246�;���!<���W%�9�Pyrdގ�8��H�-��8Yv�[�<�!ʚ��杛,
�*�jq���Br�<��}[��re]� �V���g�e�<��C�QHUpE
�Zz�]��LX�<� ��p�ӳ|\��*�B+[��"O��sR(?�d1H$Qq�!Y"O��yG醕21�H�Э�B�d��"O��Q� 
3 �1�+��<����"O������8`���l�����"OBz��W3ݖѲ��W^0�r�"O,���F�k����` SBL��"O����jD`~ܵpa�<}C�"O���  �KGP��4I��;Zt�'"O|A�# �%��a�TH�F=���d"O�Ś����-�uс��H*,�"O�A�a���L�N����L/b�=��"O�P����p��4PGhW�f�ԍxC"O�d�V|�����Cv��؃7"O<�q���GoL ��|�xtK�"O��x&6) h�۔aV"Or���"O�j��˦h��Y��@��ZkL��Q"Oti�b�	5=P0���)kM��C"O.L��z���s oG�>X9��"OPE��M�)��J5~��p�_���'P���P�2o*|;� �N$ܺ�'����JX'vv��R�]�|�H|J�'�lY���>zb(P��w7rI�'��@������>.��1	'����y��؉|�d��'BM�q-�t�6�Y��y��"��Ģb w�@%s��#�y2�'�\a�.O�\���r�c� �y�֧3A��	�.�7Tl����T!�y�I��[��k0Q�z��`aZ�yR��`'Z���F�y���  Č=�y�{�.��7q�� ��酊�y�m$����*�3h;��h����y�d��:�!`,��Y Z%qS���y��ߍ2�R�H�֚K�����?�y# '���R�%N1u:�x "��<�y����[��#5n��m(>�9��X��y2E9�"P�'O��i`(]�UF�$�y҅�=)ӊ}J�,�0?F9P���y��B [�@��]$���B���yR,��Kۦ�)�'F�D�Hh�J4�y�k�
c�N ��" h`v�{�n��y���,/�0(�vU�^"D͐�jѪ�y�挽�XѸ�^:�׀U>�y�Ύ�e�
A�����N�n���P��y�BCz��:zKx@�Ƈ�;�y���|0a��݈mTI��$�y�*�1|�N���{c(��м�yRØ�Q�\��+�+m��S�V�yRd�8� -��g�>p���dZ�y�@A�ivY��l����Q��,�y�"��sr��bd� �����7�yr�/D4��Gu��]҃j��yₖ�s�(�`�N�t����M�:�y�.�� �UFܡf�2�K�N2�yA��� +kD	AC�3j��	�'+����HX5u�2�AE[\��J	�'s�SE���:��p$ڃi�h��'nx�M�5o�p��sC&i�VX�'#�Ѳ��&0�eZ�" �/{��C�'��spᏨUK&5P5)޽&�`J�'��S`�\�f䤑��Av���'!к	�	5|�v��O
�!
�'��@�î�c���`�M�UG��	�'��r��L$�eI��}��2��� �L��$�>M����� d�ژ�U"O�E�&�I*��(l�N�X�"O�њ�B^�(�`u"�6`��#�"O"8�$J	DQ��O��<��"O� -� -��T�b�ݨn��{�"O耰�I�
'�X��G�ކ\�>��"OxH(%Q}��9{SB��JF�"OrB�f�X����dJ_�nԛ&"O ��#g��40�.Z9�b"O&��Ř)BqX����Y܌*�"O��wC#0f
\�pD��gn��� "O�����!+T����"Q�"_V5	�"O�t�3�Y�29.�����KW�x��"O>�S3!��ј��y?j��"OX��2j�������U:�c�"O�`@@D��ՂIa1��c"OZy���W;k��0 �(DE��"Oh1$��SB<[�a�Jt�S"ODX!$ֺ ����vk�+C ��#"O�d��,�RE�M��""O4qX�%�&B�P�"q��8
���t"O�ez1#\l�$��
ӌ�"O�(0�B�:-f�!�K0;X6 r�"O<l�P�fA�\Ah,E�1�G"O�0[�k��5F�yjg��Y�Ty�"O�`x��$������șc��X�<�P뀱/�� �(�:Q��P	���m�<Y�K];u�%jC��S���k����ȓR�J2����YV !S��I�3���'�a~r9D���"�bX����%\�y�`��0�Fd"3DH	0� ��.�y���̴��� �%_���eܕ�y����T\J��U�txV��0�ybg�O��<��&@��t�b���yҮ2JF"���]>"�`�Ȁ�,�yr�!o�A��)�l[���>�y��C* *[c��#R Eyo��y¨	��ڒc�7� L#W���y2#��l�@��٦0IB�	��׷�y��y��e��l�	vfD�s'�J�y��Z���P4%�?�.IY'$���yҢ��	Fxa���/��!��jX�yB%������<(µ�c�#�y �S��0 Џ�&;(� ���y� ��F]��Ib..�B*��y2&Y�I�H s�Wb�$H����y"+R:6A��Α�����疹�ybj�4w��j��^�yV�M�u#��y�H�,�jL���pzB���G��y��̂�e{�a��g�<k��ڟ�y�'E)c(�@:����[�h��5���y�^�-�����M7e��X��>�y�C�9&��Q�a�� ��S�y�J�� ��E���.Wr��v��%�y�& �U�B��޸����6hS�y&]��p(���>}j ���ь�hOl�=�'ne󣇊�;�$]�@D�h�2H��'�f�@0�"b־����/Z�H1��'���#eQ���%�%e�2nԘ�'�V$ �
�~@�e�7�d�
�'TR�QDB�#2X��GR�ሉ�ĩ<1��i�Z� �A���)~`աEO��P!�ƴ{��Is��2(Ǧ�+��_�j�!�7.������Pa��S��M#{>!�� �A���B7#7��ۧF�B�lb`"ONH3��=[�t�����p!�"O�D*�K�<[�����#2�Xˤ"O@h)0���sl6�ᗈ�=*��0���|�P����S:�L�� g�츙���I�VB�I�qUN�:�H�*�l{c��G B�	;c�<��G�/%=���3XC�I(j5�2 ڷ|��H�`�5X��C䉎7��eų3���$�;�8B�I!�.�P��J.C3��lUtB�I�K,���ս	G����ː+L�=)çy�PH7��#�.U��ǒ@d���&m�*�K�4&a3Ҧ�� ~�(	�'=Tp ���~�<��� �:I"�D��'Tdዤ�Q�3��x)�+T�D�X�'��Q�U)J�QP��Y
:Ր
�'��l���=N��LQI�}B���	�'`	z��)*�x�W�@�b�<M���$�<���)��2����F�j�tL�c�70�!��J9H�0���B/�28�P-L��!�R�c
�D ��֋1�ŉѓ2M!��= Xp��
ک��Hp��ؓ!!�d\�k�L���a�8�ܤ��^�Y0!��S�*X#��L�N�˄�FE!!�S�َ��6ᗣm��\3!X�ў�ᓻC��8;���A�L=����9�!�$��%s���b���0�w%T��y"� s�	a�'�]���vAH��y�P%!�Tո@��H�(�s+���y�AAW���#͡B𢁉�D �yb�Q��r��q��Ae��Q����y�ꅆeO ��	�>�	3�/ɣ��'���P�Od3�ɓ�a�T�'T4G'�0�	�'t��h�E�pd�E:�"юFF�<1��16��h���_���"�w�<i�!ܑ-�@
����u-��C Èv�<y)_ +�Pd��MS�b�ct�<!�B6>���)��FR*��!\q�<ѵB8b`0��GllN��Fϓh�<�%-�/����^�, ,�P@�z�<�OT�6 |D�Ç�%en����r�<��PT9���@�j\x��Dn�<�ҨͽBv,�%.ќT�t�����h�<� �G�9�B9� �-j��qQӄ�y�<�d$׃U��CF]a����r�<�"�۶�h�[�M|4]#�Yk�<y�'��K�5:��B�b�6��ф?D��f�=ÐڷIM�CCI0D��ط�1!|�����͟���	-D�$�H�2~��)����uMn=��*D��c��S�
��4^-���t�؅!��U?8d~��@�(F� �̀!�!���!x!z�lC�T9u늖R�!��T5I~|�3�%n#b4��k�Y�!�Č��.��$��1B��z�� S!�$L� َ ����I���ɘM�!�Ĉ%I�vxaրTl5PPЁ��(�!�$A<p�cI�z?�i����N�!�M:i��ؑ�n7r5���1!�DAX����QK͘(�@R���y!�đ�]%�	�g#�Z4�S!��QB!�>!��I� �D�9 �-�v���x�!򄐪z;z�ᤩi�� ��Z�J��
�'�(d�b��V��آA�/P	ޑ�	��� �i��q��EK�1-���C4"O�y�T��8�NXZG'K�0�@);�"O�<�6G!C��maqG�X�*0"OX���"���(����=�V+�"Ov�x�O�Z�,�"&��1[N2��"OV�@�I�Op$��J�&W6�Q3"O�I1�P?CF��f�I�ȷ"O�̱�l><0��%d�t$S�"O���![�b�q�$N>n��A"O�A��#�� KƎ]�Wj&��"Orl�ҥT"�y��lf��Q2"O�D�%h�f%����\,�҃"O"	��]���&X���hQ"O�u��N�-�6� 4���X�"O�9[��_�53��s��"w���#"Oj���d0]�1������T��"OT�f�	�p2vau��#6z�K"O|DД�ޠI��s�-#�w"O��Ru���}�4��#��o�1�"O����G(-x��q�R7wV��A"O�M�Uln �Z�f�,��1;"O@YV��J����Ee<np�q�"O��K�(�35�4��ÓPL�e�"O��Y�P�H$e��	��; N(8�"O�(��nD�ٞ4)�i��"	�`"OĨ��`�n���V E�֩١"O�q�p�ٽy�2q	��o�4Xc�"Op���L.Oj��ߢZ|X\b"O���4��� 1�e["~�Xؔ"O"�B ]1Z̸�Mۄ;a:�1�"O� $
�m����t�	\I��"OJ��sŎ�X��1Ic�U7\ˠ"O�)�Cש�Șh�ʞ0	
��ȓl_ Qhr,�Rp$�)��N���`��7V^��7f0��-�Іَ(`)��Y���K�+�`�v��Q�<���(r�"0!L�}��R!�Ur�<�Q��1������$��@��W�<�ր�4D�A�G(��=���E�Vg�<�"��9�2�$���ƹ0�j�x�<�V�S1R$%s���}���� "o�<�3e"����mߋT�B$�DƀF�<a@߶&�1���Q PKxp�u@�L�<��-	3V��D��������a�<)sD֨+�v�W�°!zR�S��W�<a�R4<�i��ȟ�4Lr��A�K�<qdP1:�\<�U@\���-�fHI�<q�M�s2����^>b�i�D�<�`%)v��1IG���%��́2��J�<)�@��b����P�C,D8ҧ�}�<��]���Ahm�94TJ��H{�<YW�^.K۞�ʐ�̻\�:�9�P`�<Q�HF�@���u��)���-D��c�t�X�; �X/B��m
�J1D����
?E04#s�X(Ǵ��5�<D�xㅙ�o�0$!�WD�<,�[HC�	� 4��p�"����**`�C�ɱJ?<m R��A���zb�*sxB�In���K l�~��i"�ɗ�K�B�I�(�	P�	��SY%R�T{�B䉟L>P�[����8�
#�F�NtB䉝j��{U��0���s��Q)��C��&mH\���Ҕa����,*�C��
5��Ē� $x�8�CJ���C�)� \�#q�ս�p�q2 ߵ&8>�c�"O�8��Ͱt�~e�q�ɓ|/ę��"Ory�����)�m����M�"O��!���g�,x�#�C\u�|�!"O��cnǆr���횔'h����"O����F�J�JT��Ýq��U"O�8�g+	�7J����xVh��"O, 1���Q1�Y���6a�$��"ON�Z�I,C�v9ӷ�Ɩn�
}cS"O�� ��U��Eh@E�\cL ��"O��`sL�V�ӥ�X�s�N�+�"OnLH�e�0�呣\����s"Ob�I�%�1	Z����ND̲�;"OD\X� ـz������5�pI��"O�%�@��,���d�U*y��QA�"O��Å��.D��Q�T��=J��g"O�R��`�Y���̸h(�2"O�ɻ�.ͳYۊ��隝^��T2�"OvP�TNJ2N��I�W�˓.���"O����۟��1�BJ�=F:��4"O���Q��1vL�t"���m.���"O$��ѪE�'�:8k1�A����"O2͘@*�"hغ���P6%�|��"Oxy��)A*��L�d��t%��i7*O໖XE`n����S� �'�Bݲ���}��@��*7�r��'��Q�Şh���[���.�d� �'�Ш�t��629�tC���,�D4��'J�ڴ��LEƐa��9��b�'�4�rc^��^�{Ӥ4�ޑ��'f����`E(d�.y�r��B�bD:�'�@���ㄯ��`P�ɀ�:��41�'������ɛ|�(-�P�͞1}*yp	�'Jh`{��
f̭)�E
�|s]	�'$��wi ./wz	��aY����'�N���eG*t�I(1�R=Ѥ���'y&4�V�F� ����O7>�9�'�����]�R�i"_��P�	�'mK�:h�.�J��'b�~u���I�<�sʂ-4�N�Sa�
*8J����ND�<��e��`��5��t���ZSD�B�<i!A?nN�� ��;��}� ��g�<5L�H�}i��L<(��
��^�<���
�i���#a9U��ɕD^�<QS��Q�Z0�	ǶWaj���Y�<a��I�u  ё��8Sܦ@!�R�<�#B��9��(϶K�B���'�J�<QQ-��>%�����jȚsp`��"ON���F����R��
���k�g�<Y�AU�$.X¡iV�;��@8��KE�<y��_�+^j�9C�vP�@�3gN�B�ɂl��;fi�<�ī���N�jB�	����a$�o�M���r�C䉦_�J��Dµ��E�ص?y�C�I5��� �D޽O��D,[/&/tC�8@؂S��;��萒nڇObC�ɖN2@9@�O<b#:Yrf��H
C�	��L� �l��U�"���_y�B�I�V)��&q<]3�FC�3?�B�!=��Т��V�8��W��n͚B�I�3G~D��a�	����$�N	�pB䉏J��-�����T��f�?+fB�I�D�����D�y����
dB�	44P<QqH�7l�+W��o�LB�)� ��a�f�	b(�c�V%v21`�"OVq�o'+��tc�JȬKX6@�"O@�e�%sq>m#6�OQq�p%"O��c��@8V���)��59$�q�"Of�:��[	y��g^�&�L;�"O�mj�'�C���BWg	:$�8�"O ���珪"Ğ
�G7 �8��#"O(u�'dˢ6�$�ul��U��u��"OH�੕!<��L�����Lr�"O � pkN)C~U9T��`�B0�'��x��V�8'`�?8��0+�'&�١��&#N�1���7`�:T�'����R\0v�e�_ S����'���S�5ZA���%Qɘ��
�'��X�W�UTN%��*Z,A��H:
�'_ �I`J�"v�ι�V�D�?ܚ��	�'���f[$'>V� wg� @�T�`	�'� �xf��9o�\�s�@87Ӿ���'����ʟFQ�i�����-����'���u�W��Jt�ݙ.��Dj
�'� ]D��E�f5��([D�H�	�'�\�Q0�êKTH�Po��O;Xu3	�'h�P��οf�Тđ�BH�(1�'�V*ʙ^qn�p�p���Z�'��cE�Ӫ(
�z�%�:��!:�'Ԭ��Q�N�p�B�D��t�'���Ə��1aq����p!��'���3�ŝ;��-1�I�24L$�'rla
�c˄w��8"́�*{|=2	�'
0xH'MXI��q���ύRxZ+
�'%.�)�˦�xB0�>O�(y
�'�8��E.i3��	e���{�r��	�':4�Jf �?�6���C�&�t�P	�'���Y�L/�6�`�%��MX@T��'�b�1'7M��R���;�L�	�'g�-H'B��"$+a�(��'��,j�ʒ�dG�HZ I<N����''XL:�OG�܅�
R��j�%��y���8'
$��G �M(�a��J��y�F��hx��G�L�	 '���y���>���`�L	19�(��ꔠ�y"��Y���@f�7C�*�نM�6�y�o]�~X��r�,Y�:�\��j˔�y�֋4���	5�=2x�U�?�yb$�)Uň�j̗�e7�(�T��,�yB�oEx��!ɹ#w�-���^� C�ɧ�pb`	_`m�vD�bh�C��|�;�)�(�lвFY ͒C�	���<37�L�_�<X3�ȑ+Ea�C�ɱ7 I:���@�$����m�C�IW�����Tv�:�{aF��rsvC�"i"� '�ʪh��3����V�OD���F�?M@�"��~F�0K&"O��k��bվTJ$�Z�'d��b"O⼩Pg�2���`�0���� �iA��䕹<O\��fe�CV�#P���H�!�d��μ�cg�8.6��	�-C'o�!�]4B-�@�х:-"�!��4�Q�lE{*��#�߮�ڦ��j�j"O�mx)��+��C���bߺ<�tj�X�����O��d�c�7`�>��慦�y�A 9\>b�k�"\m�M��-ؚ�yBGJ�#6�t�N��)]�	آ&�y��[,`\(a.F��:4Q�"��y
� ��1���<	b��/=;�qi�"O^H��F](%ԕ��Y@����|�'P��UM�c=2�0v��n��$�
�����:'g,����
r�z`�.�m`!�D�j��p�*�y�<{1m��A��'1ў�>�HW�G�0@�]xQ�{�j��S�0D��*4��'CP�X��^uA�}��!�	m���
A�_Z-SM�,$\��'�#��3�S���O~��&S�iʮ�@�� u�t�����7LO�)���y����b�؜o�,���Q?��	�Vł��2/i**���Hq!�DZT�dۣ�M�T�"��8`m�1��B�IDg[=NX4i a��>+��ȓ���S4 Qn������m\��'���T�]��5yu
��PEn���������c
@�K�[��ā�j���� ��{��)�i����B�/-#q��C�ဈSU�v�'E�O?7mӷN� �ቀ�Ft��qB!�D�o@���5.A:C
6�R�n�2]'�͓���hO�S
�Α�¾>x��A�4$9J��D��'���*��Z*>��%	:B�\Y:Ó�hO�����Fia�Jٝj`)E"O�0�akT� K�r��ܴ=G�`���PD{���ܚ���b��U�v�d��e�j azr�	q-<\��Kњ�p\d!��$-�AH�;J�h�24� �Id1O��D)�)�5>�2\ �� ?NF�sBE>[��B�ɴb�h�*C��TV�X�"�&])�b�PE{���-��jpl��� �X������y2�?%�.h�f���P����'O��y�k�1f����!1��������y�a�2��L��@ߣ%}���c�Y��y2��)���R�B��D���ް<���d�:�� 9��Ẁ�:�Ӧe�!�DL�ް�+@h�N�	T�K�g�!�D�<1����ɐ�>�H]R�.��!��mv(-�\I� &n�]#�v3�'{*̙s�üϾ�fB�$p�D�z�' 
� ��	�A� Q`a�(� �'�F��m���a�e�.
�d���r�)���	�>�@-̌UӲ h0ȗ�y)��N<I"��2T}N��V���y�#Ud���ӓk} C���N�bB�	#j�D���#��&�̺��4i;��I��y���)U��9!C]&IN�LZ��q�XG{ʟȓO*}�E��@A��!#W=5B��"O2R��߄�JLiĂQ�ܬ� `"O�pv#��"/T��a���>]��"O��j�(����
]��}
�"O�D������JT�����\?�%iT�'�OT,�@a �=԰AB��5 ��e"Oܔ�"O�7f����:R�t��P�����ا����f�-Y��9��h�N�A& �?��'���ص�Q!W�X��e� � �"�i�ָ'�F��v�Åt� ���J���y�'=j�u���
� ����W=�Bԓ��:�S�I��>9��4��* .�u'ݡC8�{����0���ۮ�2Ux��E�rB!��K=)�xu��K��ΰ���X�!���O���qΛ�4��Pz�/��u���iP�~�DX� ��c9TT��)ܑ�ybc˥+�����Փmd�`9�c
�M6jB�ɷj�8�#�M�A�x+��Z�(C�9U ���)�j�P�iЦ58FC���� <:C�T&2�2-��aR�kqn}�"O�����J��88�Wn�5^�y+��'����n7~f����uS�lJ D���b뒵#����Y���'>D�4�!/��$ǌ�Is�V?qSQ��:D�L�P�zv9��$U8����f7D�$��Nr�iʅ@3�vq���/D����[�?�������	bU�b&"D�l�Gi�(cBJ�#+G:I�Ne� f>D��
q�E!%�Qr1`��J��{G& D����T	N��
VAO�3z�h�(*�O���-g+�{���Sa"$�&dKA�lB�������)0����FO$%p�B�I ����t��=v��4�	&�RB��>� �״s���HE*��0-PB�ɼt��[UcF9Xo&�x� "%8B�I�K��I Z����ψ/gB�	�Ҁ�鱁ǻ���3ςc]�C�$��p#£!�t{��K�Xo�C䉉D���C�<=���Y!�ݬgtJB�	c>�u��d�Lꂕȓ��'�0B�	�"*�h��KQ�f�&�b7�B�I���02��<x��1���B�I19Np�)���^~6�ٳkE�b��B䉤1�9h솜-'4�c!j�VB�	x˴�Q�/����P�L� �$B�	�5y����-Mɬ�Z�
�0�TB��>w�� &�\,h���8���=D	H���4}�Ą+{D8���)T'I��Az1ˋ �y
i�bVсv��hʕ�ڨ��O��~Z�ǁ�%��GoP^��i�R�B�'��y��D
WW�ҤL-R^Ҹ	��@��~�xb���}�� N�t���n��j&a���x�炂i���sb��V���d���y"n�"��Ěw�ԧ

��2�P�y2�8��K�9D<�� Z���'A����%4��htoƈ�e�0|�tB≓,�HЀ�MbJ�ڶ�\%�{I>���'�$9c��=�ɑTh��FY�$0��y���	w��`s��Hh�L�3���yrƟ�%"$� ��!;���c;�0<���^3O&���l��D̦�Bff��!�)�����˄Q�^9x�%�1�!�O&j���E���m J��!�X8�4!��]��1t���9�!�D�1��8�G��w��u@p�R�&u!�$�+G�XH��*J�~�2i����:g!�E�ԅ�#��0�͌�e�\d	��x��7�S�'fړ&�%g����*�:��؇ȓ<�����X�����P%��P�ȓ0�l{2�˜]^����R	 �����{?���ɀk�d����":����ŝd�<�1)�#E<&��ၘ`/���Snl�'�?�!�aT��UóaH���HD2D���n+!�,\B��b�^xA`0D�|P�&;�� 8��C�:t bD.D�aHM:�����#��l�#�*D�𚣉Œ6��Y���u����3D���F�0gZ�1��
�9-�`ӵ�5D��J�@L�.PR�7��X�~D�á'D��Z�ć�:/n	k�̛�'gHLS�"D��5�۶�B��W�M�3A�� �$D����X�UtV����L ]�yrើfT$C�n�!�<�#��_=�y
� ��V��Bq�)e�A�L+h�"O@���`��1�bMs�A�Lrd���"OQh��m�t���eV�H��"O� vɇC�b1r��k��U��"OڍɤbJO]��*����5qS"O4;U(D^�rl�d��<{���""O�D�1��-8|���]�.MP|""O�x��@,�<A��Ǎ'-m�Eh"Oֹ���c�<ܰ!!Z^ج�S"OHr����#��س�-�y��׍"�24C�̉���k�#˾�y�K�1rn�3 �ɠǀ�	R�W��yr��w�ޕ`��
!��;lN��y�폘s\��"���ga�ar�)���y���4ʨ��g��n�ND�����y�kN/�T� VaڌiSX� ��ϸ�y��ǓMjƹ
v�
=i�ڬ�!���ybȘ��Y����q�j�2!m��yҫ�4�\Z���S��0C�΀�y����f���C��M��:7d�-�y�n�kr�h��@��@��d3$O��y�e�rNB\8�M�>{̌�Q`��yR�Y�$���E��<aӄ�J�!д��O�c�u�vI�׌[�X�*8�4O�0�pF��Ew�i_�$�%"O*�@�kX!l�H1�vo�2@T(�3"Or1+�iH�{��jc-�V�􉃲*O�`��Ҍ!ל�9�e�M�
���'O�=S�&�"&�)�e�9kJ�h�'B
d�hC�{��X+�O�b���')��	r]�jhe�4e��b�'�$yCR�6f�T�-!7L�C�{�<91�N0K��b �Ì�@=(�n�w�<�G�N�>e:*ciߊs�l���){�<��R�|�B�+&L�GcR�#1ƑJ�<Y'�
:Z��s���O�u�AG�S�<������"ue��^5ER�C�H�<��-��_� K dT�L���ȰB�R�<�@����~Q
���d����	J�<��F�g�ec$@�1Y��(��$_E�<9�lm�*��'LS�(m� :T�J�<9��A�8���V/�e_���#��\�<�� 
� �X�l�*)�����C䉅@h�ȗ/��`5���W+N@�C�%V�|y9��� ,	��
3AU�z�C��&cb�Z ���f��q�;eL�B�	�@���!��)r.����#�JdTC䉙��%�N4찃�Ǯe^�B䉩My�4�u��yF�Pp��B3R�B�	?:���'�1?���V��?L�B�	�m]d��M�9N��A�[��C�ɇo)�c��r�xҌZgC�B��6~���3F5K�P��X�"x>B�	������9� �Qf�W.[w�C�	�g��M�*�����;7�B�ɼ{�B��@k/d9�3V@\.^#�C�ɔ'�0��u���{4��k�t�C�	�{��|"%���e�1��ڟO��C�	�L�(ԀP����ese���"a^C䉋]:���aI8ņA��H) <�C�I
z�P�;@�]�wN �L]-b��B�I�
D���ǓrTp$3���V��B䉍5(� {���H�CJ�P��B�� �=�D$��Ov6�D�S^!�D��?�Uٳl�(#�~��$A�p6!�� �|���cbv9@�lZ%7��"Oz�����&�1�,�(˴<S6"Oޥ��}�:K���^��f"O���1V�i�-1fa�Q��yC"O:���58K٩�J�j0�=@E"O� ��,���29�!f�B2̉��"Ol�P6#H��㗥|�������y��0A~�Ӳ��$���=�y����E�Ai����$��e� �y"�C�,��Q�a�*�I!�߈�y"iX� �J4�,��j��`F�y��k��uHb��<��삅��y��.kCfٙ[�l=� )�V	��t��q�d��6�]kC���F�I�ȓDj 
��Ǽ+��X��?y�z��	�Fnz�ʆ7�]x�Lp��X�����h��0^ђd�
��#�%	6;O\G~�ʖ�Z���D]Q��B��pH��A�/��m
E�m��C�	�q�z�A�b���r���%J������	3nV�l�(��h���
��j��$�'�B����"O� �f\"F����P� ��ȉ@yR�V�+Ob��d�4W��5���X�iB�������~�&G�4�D1�QR=7Xi���)EG�����0�4�;Q�'d^0*wCC�s�������(.g�};���E"q=,XZI�>���� P��r�U�aE�e��F"O0ذ%m�*N� @�EÑ�p~,1��ORe���.����# �<E�t-@ �B9��L��<��o���yB+��(P�N� .}���V�v�9��`TE]jV���U�v��@Y�lH@1ɐ1��bF��If��$K	h��g�3F7F�򒬔;��R�N#z8!KTC4d�b�r��٩��O���[�T9dM
%�7љ0������\*��5C��?��'Cǚ���
w�"�z���? ��V"*��f�V�o��P�>�6yL�ɂ}�lL1���	u��j�+�"Na�˓R("����.��S�'�z�0b	6nI��Ӯ2�x�8�bL�$�h�'�9CȖ�w,���&|�d�!�%3.�h��S$��4D�?��&�˶��Ej�O~�(��0_���3�[�p��ؒԉ�&U����� �x�Cb�d��KW,T9
��4NO����W.^�D�x�C�9�?��g"�b��EK5�Sf۴���l���]T�C�	�E��pP�E�C�d4I ��7|\�I�0V�YČ��oR�c'%�	jV����!dS)hmQۃC��8<��I��☱$	]�V��Q`�D��r��L�w�֓L���C��'J�Qh�	I6~�`5�ቨf �ew��<8�,|DL�@�?�Ɖ\�!��<��M�O(AJىm�p��cHG�g����Q�.*����w�׎�x2㗓c/�U	K�R�LK�h���V$/I`��퉢�y�؊>mdE���L%A�$�q��/E���#J�!�Ă[��z�H�ZDeㅢ��:N(l�F0��� ������YJ~� �;�Ĝ�!.ꡣ�4|��i�KQ�B��9LGV�!t���jXa�KL���9t��@�L���	"v�xw@�T���3
�q����];V}ʊy�nѦB��J�㋸"^Ss���y�-��^��c�����Ai�0=��E�L�z�'��Z�X.��=[̙��pmc�'n����jUfQrE����/N]�1cK>����LX�9kçX�H�BPf�!5/XĂ2掔J|l��T�
pI&.� \m��$�ږL^�xe���	�,������L<!BL�UyTo�?d���:�cIKH<�ES+Nną
4�Z3z�j���iA0#8��D]�CǨ��D��0Y8!��cʘ:�.�}ay2�� ʌc��Py¦��82��hU&\{x�����y2k�<�̚%ʈ/N��x�@\��	�X��� :!Ub�'!�0IB�=j��*"t��-�SqX�&��k��@�j$\P����Z)���U���o�N����O4as���!����KhĠ�]�/���b���>�6qG{ҍR6f�Kǣl�'5�A0�&N ~�T�y�m�C��a�,6`�$�g%�O� �8����}C`��%}��t�$�'6�zAkZ5 �fT�O�d��l����o�\y`�5�tmy��Hd�!X"+\0�y�J�"�q�jLL������
���+2c*��è�'l)��O(����&���T�<��(��<r�R v�/[��}RB�.^�Pu���O��L�`�	.��&�H<jY^��{Rd��-�\c?�$`���B�Y�3�'��<,j(HG{��f��`*�E{�'P��5�G#���K^�]e���V-D��hA�̊M�LRB;r'Bx餮�O̼�P$J&@)x�3O�"~"#ID�w�~�)d4QP���b��y���=G�2�c4;̞�˱g�:��D�:��,C6��|�N�𤋄@���Soƹ	Z�uAP��}ba�R�\(�J x��U��!`����N5/1��G�U؟�j@!����I��K-u���N)ғwHT9��ᔁH�0C��:����/K�K^jFܘѮ��9�"OL�p�˜3xR ܃�
�q�ư�C�i�t�SV��xW�Y�dNٙ�"nZ`�Zt��޻;D0��Y=M3�B��R�0�Ja��\�|�Sc���h�H,9�*/D�	�e*W;1^�	�,�?�=� C�$8�Q`	3(��L�-�K8���rmK7S&0� P�L`28�e��
B���k��d���_Ta~��	?~qb� Mz@�d�O��Z�Fɛ#jкt� �,���|jT��$~�4yC�h"4��9�AS�<��.gǊ�F�_6��u�Tiψ���B��Yk�9#�]5J������9�6�4�XJj� A�]>k蚔�Q"O��RUS ~**�����~�����)Wg6	��B�@���nF��DF3��R9g��#��`@�¶A>���l�T�F�"t(�R�h¦}�5� � �z�"烏X�0D�W \<�}Bj��#1h���!���۳�0��'�����؍Q#00�띖
<�P���i�*ޜ���ֈn��p�!�d��t�Sf��>�00W�]T�Ƙ�M#?o )��A��w��9A�I-§%�4��D(.Y��S�h�@.�:*�B��e�a����>�3Jy��x��$�$�;QaA#<�r��Ǡ�d�I���d�+;�|���R�d0 [7�A�g0�z�Y	�Ƚ0 Q6��0�N[�bx�ґv�R����Ήw��{&�,�a}"�ߜAE9p��*
��0����'�~yH5��t��j�Ȁ�lPH0��S��6C��a�O�%� C-#	DB�@Xi��/�<Cn�	�LTq��I��Ĕ�+���F!�\Ia'����O�0��;0����=$�R4"����sUP0��i��y�!�P#t`QK�!GXPU��i�z$D�	R��$h�Q�AJ��Gy�'���S)��LӌA/�yC�JM���=��ám�P�1�!��x�Hᰴ�ӁY�Nh��n͖z���[��O.5�UkvX�4���=4G�͡�&U5%����R�9��:[�8{�C�{k�l�!�+iM@��U?񪒧Z,*���Bզ��@ӆIZ��*D�0!3��=1���I�`R.L�=(F�<i"�I� �� PMa���F�v$��%d�L\N,� �D�<��	 V`������#9 ��%�.��=�2)#�gy��0wN�iV��!�E���T��yҠ�.@B�e��4O�-�DNE��y"�ɝ	[
����?I�,�Ϗ-�yR��nRz��q�Wh��0Ν�y"b�4U����[�� ��y��G�6�8��M2[Gte!�К�y­48�(���/Y���8�#�%�y�oV0M�B���̈́SUdP���9�yR.�,7rdqj�Ο�Lߪ�ʑ����yBK���|:G-��N���ѡGZ��y"5xdn��#MaP e���yB�P|��e�`*Sa�#�yJR7��d鳡ז'�4 g#�+�y�!M)X9ܑyU��V����ά�y���;��S�k6�������y"�C���V�L�:5j���y2���'E4m9�	ư,�����!�y�#��-��?
��Yō��yL�>d��9C�1P����4�8�y
� ��Q��U|����f���{�"O��1 ��M
�x	��\�\�Q"O�p�c�z�\oIR0�ڀ �"O�9���9�� S��ڠiP"Ot����J)^jp��M�"��ԫ�"O*���B�'p� y&̈�k���g"O�b�]�
r�Qa�l�&G���0�"Ot�1R	�/y��jT����܀�"O��0��+A�F��jkc�x"O<���er*xk0c�vFd�1�"Od�X �Ұܚib��;;�ȶ"O���EeD 0��y(D��I��)�"O�@���H O��`p'k�+��Y""O�̙���L����wj���r�"OuZ�d�Z	��懘�n�p"OA)���w�x�0�fJ6;�	�"O�u���B5PIXU��8>V���"O8E@4�jdz`�V�J�V!~x(c"O��{�,��Y����@K�t/��"O�	�*N�k����4�J5J#�h��"Ot�k��"�P$��-G��P""O�%�g��4h��@"B�/!: ie"O�]�4fE=f*\&jy�(�"O|1x� ږ[z��[6�˶l��!"O*Aò��#*��E��[Yx{v"O�k�.�&d�x"&J�[�l옷"Ob�rJ�Y|h�c�
0�|��"O�P�ed�24����]�`wJpR "OX ����3|/,�� V<��d"O�ax%-�5gV@c�+�.|C<	[�"O����@�g������PPC"O�ё�n�=�܉�2��g�B%: "OL�S�P�c|�E����1a�p)m D���c��'k�H����&8%	�	#D�Dk���Fp��"oFH���?D�ܘs��G?�\�WLۉ�(��6�.D�@32fɏz���W`�,���#�(D��Zr,�K�8UA"C t�{��'D����
;u��Pp��/�2(�bM D��S���h�*}S@�=.��(S�:D�
��D�7w�� �˝�o=�R�6D�pj��K>*1ġar�̔OA*��N4D�,������H@�7�M�b�,�;��)D��V�ۘyJR�c5
I�z�Ƞk`'D�\H�.X4�T`��еk[�  �# D����S�iN���@(CB�]���!D�L ����P��"`Ûdkp=Q�B3D�T���DT^�"�.��#�p�ю1D�ě��LJ����.�k)ڄ�sg-D� 15�_0i>��'��Z��-D�h�h�,��ĩ2��/��`�S�+D�43Ƈ̒��U��y�ڝQ��%D����f�E����F2#ʆ�Y��$D�����nѾtp2�Y�Qr�C��"D���ʌ�X��0ťS�j��x3�c5D��:�k�/ �$|�fM7Xn��t 1D�D���/2O*�A	�p6d��&-D�x�� %9�(�"���N�����*D��%��"VZe� d*��B�+D���b�	=�� v-J�[�ޤ��<D��Y���:�0��f�W' ���h�o;D��Re~��l��	���誷J9D����ξ,J���P-%�jyB��%D�S�'�2�<PyI�D3v5��/D�� ��3�.H& ��I��f*&�((��"OX�&�D�7k�eP�d�C�.���"O���e�*M"��Sc�[V4X�v"O|�:d�L�D��scE��'��;�"O��$�\IA�RB�P&�`"O����Іm|X�'"N�e�J�cA"Oƴ���	9J�p;�Ò�6�1E"OLu��i�Jʞ0	H̴,��]�"O�i�����$�!0߄��0��"O�p"fH�[���F>O��(�"OZa)��^%C/�=��E	�d�@H��"O�Q�ՅwE$�j`��f���7"O���&�H2���.JC~�8�"O2�R���,	ܪ0#���KKz "O�Ѩ6�Mq��ႇ�Ơ����"O��4D��q	D�JA���2lIC"O֭s�)�1H�
VBF��tU �"O��bÅ��6A��!�T7d��"O@���@�Sc��� �3b�cg�'�D��e
� �HEs��=C����C� vȢ�Oʈ�EbC�?�4�*e�2})���,8�!�)W0i��O8�T��5\8��� L��N�Q�'�8�`Ѡgl���ϛ�~�82�'�|�c.}٨)�CV��}���^�K5L�+|(H�S%��h�<��ܪ4�x�:� �?W����M���剃&�L���LW4%��g���@�WjA�Cۼ)!��������&Aa`�m0�ԡ��hTi&z���Rb΀P3�j؟ ��io�A@tN_C��g�*��$����B��Q!L|rc@-И	�" �U~;q�Q�<Y6h��*F�Qj���2_>%+ee�N?!�m�c���R�(���Ӓd�d�y��*Sz��YU���7�B�	&-�I���H-f0"Urai��y��p�)O�Ѹԉ�xH��J?O�h��B��B$�墌�Re�}7f���zi�	��pq���?7��}��d�*Nv�ؓ�\9B&j�K�k[��Oze�$I��W��>�����(��	�l�@/�M��b4�.�Q�vf�fJ���̋%�f1�(S��_ ܉���O�U�5������l��4��@~⧗e�٪���*���!#!͝���4䮌3�,����/3��4�@ҧFhdPd� Z|�QX���&"�ɶCf%�e��g�axBeO8t@P�{1�P�&pv�#�$�&��O�	i��AC�����%��x�ӎ\(m�x�3@J֟P�:K�팈S����7��	t�'�es�M��w��XB��<a�E5,H�9�#�O	��A�2A�R`�����$K3p�YT��#F��牥�y"E(("�!v&��6��.�&tW��dҚam*���`�G�j@zO~�q����E�l1�[֠K����9��Z�{|�⧅�i=�G +��8LTt=t�1ԉ�zZ��Ɏ!�TMwC�A�ax���Fl�a�����^C�u��b���O��&O�t)�J�9Q0MQ ��+b���M���sk��t� �(���� I%*&ƢR�uS`U���<��b�O��m��n�4P)�9+���}��A�e�&�P��"D"�:�j[c�<��k�:��m2De_4��I:����\��D!+������m	䒟���M<a�董j���p�:M��Tz�E�T<i�hѢ�}�E��4��)vK�$'�v����Z���?��)Jr�؀/3W�֨�u�T8�,ٵ"��]�1O.�rU��a�����T�*uԕ!�"O|trwn47��!�g�.��e�3�'���ȓ�W�$�bXɓ�H֢c@��"]�yD!�D�T.E�s��>q=,!���޴B�'<(1��J޵Ca�$,Y�,����!�K%�LYd�E��y�	��s�ҸE��W?���Ǖ�r��<)��>��ⱟ�'�$i��GC Ūh)Ȕ�4��j�'خ0�+�.��@Y�CL_ܬ�d��x����̏Tx��8� �0dF���і��l8��6,O̘3O�+:y�(O���!/��N��d��蛰rI�0k�"O*L��t�йxQ�#7���A�>y�B
HrT��#�E��ř.���π �z�B��z���h���c,: YW�'������c'��4������i�
X�tP�!#����4�3�D��Ռ�ᐦ	3��9�c� �ў��i��`g4�y���E4y撉�푿L��x"��g�Y��n�d����WD%�Ã��{oUɓ��<K����ɲ=:XQ�W&є>��?��$/�!)~>�wY�x����`i$�[9P�dK�	�y�,V�/�`���H�g�|k������ s�1��Y7�@�O�9�SM��	��xzua�S�t���R�!A��}"i� D������G�����6�<�ٗ�Y9B�r�{�육} c?�d��e�v��;���1�K�.f~D{b�پj�-�2H�y�"��a��������G"�͇�U�����d@.n�6����=脤���I̲hk?�S�O�A����H���B�E��1�
�'����$\	#���s5�V7#L)I+O�`�.�X[ք8˓K��	�3\d��#�@�ZpRl��I-9-�HJ5oH�y��MQ��J�t%ȵI%,�
`r��IX1�cE
(צe�=8���D}�B?R�D�$
��s�-�P��Y&Ȍ��H_��yrʌ�\�ʜSG'P�Kl��疼�yBT �P�QM�?��ma ��y"Ȏ�G@���V)`��-{�ר�yh=?��U(�K
7hZ�)*	�yȇ�� y��ّU.@�d	��y���u���Pc /ؠ+D&K��y�惓8���T��^{��#S郆�yBoUs�B�Y�C�^���@9�y횤yԨ�� Ê�Q��\��@��yb��\٢Q�zW�@ya��'�?��m��p���C>y��
a��_�~�	p ĺOa{�߮9�H��OV͠��> �[���Ԉ�"Oz̢P�3d.����n��:�	22���y�
��Ö�~��� ����O�șy��C�m���o/~�(���'�*Yr�Rb`��V��-Y��x�r듓 �"U �'ɺ���+�>��R5�����ȧn� pPI޻s���A"O����A�/��Bւ�.!w���O�]����`H�f/b���:\�蕏@N�'��Y�AB��9����#_�-�דoi b�AIb�6�ć�A��9�g�![�!�r�B�C�:9+��_�6q���L��T�#�%}}(x�R�݁�p��=9�@�u4�H2���O,���A��t� x(��`X�0��-v`]�+�x>U��"O�<뱇ڵ>KLM(�@�4��#��L�q�E˓�'TSϏ2U,�4�2je�u�T� J�^l(�� 'h	�	آ�"D��v���C{E�!�'(tn4�V)C"nϬD�'�%0����Ť�bQ( Fz­�6�6��P���.,A1�F$��=��a�'-�؀�'.���1�'9�����!�$����۝YdU��}X�c�'3���i�%�jf��p��"�I���U0��O��A���i`��x���Rb�R^I����[�l`w"O�s.A�`7�S�~+Љ��|.ĩ��)��DD��pf��(g�K��Nc��8D���ʃ?ʐ`�@!LX�Kѩ�X�>➠���<Q��Q��0�`�g�����i�I�]�<�dH_TU�$J��/��9���T�<�2e=Py�ghƒF��Yq6@�U�<y�l�&=$T;���X�*�r�,_�<�2ß=5��`���I
B�D����l�<���C�8��3�߆0�rx����U�<�W͸W�PMB)U�j|QHP�	V�<A��Êa6
�)�\=���a_u�<y�^�@(b���Ν+.�V!l�<ɐgӝnr�ch�Q{����jGq�<��ᅁ=P|J`HO�	�&qQcIw�<ٕ)
�̵	���Y- �@ҫQZ�<�E'�)~���g!�۠\;d+R�<��(K6d]@˂aZ�i����#E�u�<If'ƥQȆ�`3�^,Z��C Gm�<� ��Dg8�����%f��1��"O6IҳC�%�h�j"��u�! R"Of��w��vڼq���1	��YC`"O�L@G��4'��=�7%��M	R�"O|l;��?'@X(DE�2K0��"O�8����#m�J@�ߜ<
$��@"Ojy*$��teD� ���Uz]AE"O@|"! I�!$1��k�j��В"Ob���H\
l������ߟ'�a9d"OP!01�@ 0�^1犓<�@:�"ON��5B��8 s��Q��!�"O܁#ǀ�"'�*V�=M� ɹ�"ObEI�'*"%��� �A����"Ot���"L���(q,�Rr��2�"O��*Gb�U�t���HyR\@Ɂ"O<���	�\EFd���^0Q_�驐"O�������0r��3'ZT U"O�P�⃑�VKL��*�^4 8�@"O�Ȣh�
^�`u(AH_�Z/4i2"O�ʴ���K�䜁�_�B�dC�"O�Ab�2.Q� SEҖ���e"O"Ժǅ�#خ�"t��9���`"OX8���Z��6i�n ��,�s"OHyK��-��q��Ѯ5�!�"O�(Y���y��6�_3���Z1"Oޅc�'L�~\�1�:�� ��"O� �R�/!L���`�O���P"OL��w ߡg�2�7aU&="2 "O
������CR��u��B����"Or���k����s )�!2�ق�"Oƅ������\�gOԣ\�F��s�I�Wݢ�pS♒,��
tK]+8{��	�x����V�����k&e'�n��~B���ē�>�s�e� ,+����n�����A�OD�I1x�OQ?��5�Ոx�@I�M�)�N]��f��@�G(�)?��6�ԑbnS�Y���gÓ�h�!��B���p�	+k*��e,��C�ў<��ӳ^W6l17�$(�,rnim���y�D!}�����N|!B���,$�cR헆��'%�#=�}�G�#b�ґ�<T|~�:�K8yH牡�yҷiF tO?a��O��'G�L	&�vۦĚe�z��E�vċ`�,�(:^���X5"vnϬ��4`��RĆ�Q�cy�S� �A�Ow�P6���r�����ia��4��'"�p8O�?�&��eqJ�aD@��,1 h�FhV��ēX�l�OQQ�,���0�C���Q��5?�q2O���;}Zw9��SU��	,�	c�Ds��u�s) �yB��0�N�9�4��)�)O(����
'Rc�P�B́AOT����88�VJ,}�����T�r(�0 %���l]�0��)�ynb-)ߴ��uY�O�Ԓ�vݥ��imq�Ɏ(��q2��q�F]𧶸��'��(��O�b>�yt!ÐE�p]���,CXJr��<�e�Ə�����X�(����]҂Tk���i Ԭ� �+�n5�5-5z�̙�'h�P��F�H��\�D�2�K���v�4U8p��K�¡@�=4��`7o�x��� 3��C���'������:�Z:���$�,�	�-�֕H��O�,"ҏ�+%��M�f�d�x���"�󤟄j�CF�� �0|�#�K�hAڴf�H~����K68s�vI[�H��Ȼ�ϴ4T@t��'?H���4Oר^�*q �
@�m����y�D�bD�CVXi�O�����dY`B'��o����
*���լM�O?7��8���X*���g�T�!�O5~��Z�͵?�I{6'ON�!�D�HI�A�c,i�胁9N�!�Ď�b�Ћ���/�t��1+ԘY�!��E�Tc��n5hu"���8oz!�䄓1�r`"wh�
��ؙ�	�8LK!�DW&�<8��E�q�D@Re�ޅS!��]1N yH⊘y~�ؙQJ�2!�� T�����}�2�B �J�)�����"Oȡ�ւ����dȚ�
�����"O�����W�W�R���J2-N���"O.ܳ5I�"x��\����#);rmZ�"O:��e���,k��R��wr��"O����؜z�pd���?S~,C�"OD�r��A�x���A-%MB��f�<�5�V
t�ذ�Ɲ���s��_`�<�T�«�؀�B̓+��A�[�<�!�S6l��䁥b1Hh�-�v�S�<a���;a������ ��5�5�L�<ٷ���W�~p��@�{�)R!��K�<���%nNh��`�<\�h5qw��q�<���Ƚ�b|a6#�:�.���E�p�<ѳƝ�2vds�fء����"-	t�<IL�1��a8�I�!BY��KT�<Y��
���̺�˻�<l��D�<�Q �#p|�:M��<`���@�<1R�Q�)���O�E�3�P@�<�3��6��P�t�DA��P��y�<	Fl�;BnY��@�#R4��E�x�<���w٠��w��`�8#p.�L�<�@Xz���Ir�2M�Ȣ#a�F�<YT�S�;�R�C�G�Z��`��ZH�<a$g@�]-J��!�81e%³��D�<Q�J�,-��B�F=W�\�f�G�<���w�(�N��?~L����m�<9��	0Ds��pQ�;r���Hg�j�<	�.	�L�6$
"iNU)e��f�<ɧ-�$0�K�B�%���`���{�<�cL��'L�#���lQ#2�L|�<��5W�DU��I(d�P�r�JT{�<yt�;�ڣ�#q��1�x�<�� &5�$����# ��2@w�<�@S�;��H"�EW8'�t��l�o�<Id�Q�s�@���m��+}�5q�iRq�<��)T:!��%ұ"V�2�ȓ:k�i�C�膰:��ޣN|�D���D݈'�(���S@аa��X! =��!�(I�( ŏ^�U��M��(�t BKщ*K��2>F�H��qg�ea���2b)���7:.�d�ȓlh,��w��*@�D���W3-�t�ȓa����&�Ч1�)�w���
Q�ȓ%�$��#웍L�LMдj��n'"ȇ�aP�s �W�^!��S���A����e�f�7�؁i��#c�ޛ{�j�ȓ`و�YC�:p��x&�Q�m�v��ȓ�V���,	�gA:�.��yR�[�t9�`82�Y2b�B��aJC��y"�'X�
��0-+T��8�F��y�dP�.�$Y�E`.�30���y�*D�z�&A�R�
�8���S`�/�y��Ȋh�<��O*��;u�M�y$�'!ij:�B�$�ސ�q#A��yb�����!��)�buKD�U*�y�Nѕ8�@�`�H4:V�8��F[�y������t�5��d0�(�#�yk�܈Հ��� �up#Y��y҅Ǵ
���ۡ�VA@����D]?�y��C �,�a��9`p:�����y�S�F��� c3�Z�S���y«RmH���� (�n��7���y����_����6w��CW	�y
� @܁��I�Xp$BMX
V��yH�"O��C��,�L��M���R�"OTY�G�˼j�N�#R� ��Z�� "OX�J�CP\r�Ђ0/X�"�~�;$"Orl�1&=yD5��i�"O䰂#b��n�@��MC.l����"O�����Pݎu�ѡߩX~��A�"O�9�f�B�%����]i���""O�p�d	��#��)Ss��&xZ�Xf"Of��0�U~~ �����O�6i��"O����Ǵ_g*`;��G�`dp�JW"O(���ܟ3�. ���>	V QX�"O��G���~p�̗iULĳ"O�9J�����d&��s��q"O&]�`.
�Z��T/�0Q[���"O�|�3l7O�!kUL�XA8�y�"O̕�����l�KU�j�18�"O�`�ҟiJ�C�i�18�P��"O�4��K�&%Zm(�n�Z��<a"O�2mI;���SG�,DF�,�"O"L"��N��	;��Tބ3�"OH�����T�T�i�/ϫ1y�M�"Ov�����Y� hU/�#{f(`s"O�{c Z�,�8�k������"O�91���--J����HB��"O=#����@.�6OɂJ��(�"O��@�^�b�����T�J�"O����ǂr`�RE�D�V-��"OH����Z+JY*'L�ty2@��"O�]�qi]�S.x哒�T/D`TAs�"O���	��u����.Y�`�"OVAQ�X'a����w�
�nQ���e"O��Jt�6nv��� �9�B-�e"O�`#�=2j�����K =vD���"Oh��'G$a0�I�3��/jN���"O��CS(�:PY@ $*i���W"O��8E	LB2U��)�#3c��he"O>͢ �۳-H�s��=ZO�}"�"On�b6$X?g��zW'�E���1"O�f��)h���PH`YQ"O����H͂}T��"��ʸ;c���"OLXY4�9q�(V��7Y~V�3"O�%h�&pĘɉ�B1(iV��'"O1�UcF��9[ӮJA*���p"O.e�����_d�!x���5��"O.��$�~�*�'n�98�7"Or��Tc_"k��a1�ҤC����"O��[!�
;w��(Zgb��Z
�RB"O�P���t�&ف�g=-��
7"O��vo^<V���z���|�}�"O�8���P�\ 2�L�ZP�"O�ayrl���<�J��[!	�aF"OF@���8\k�` �Σ�u�e"O���g�+0���Q�5x��S"O��9�e_��5I1�ڲp��}Ha"OpC��Q�~ȩҡ�.O�����"OШC��Z�d�hH	�c�*�>��6"Ozuz4g\-~��$XsI��@��"O�zu�D�k��x ��i�I�s"OvD�@��H�4�A�&?3��Ȣ"O��J�˙�[hy:4����R4"O�����Pv�J5*˿~�RY*�"O������=Nҕc%��5,�v���"OHd��n��ҩV�58�(�"O� ��AE�/S��b�ħw8J x�"OBSa�X0=�IK:`E\p�%"O�=*��Maci�⃄E�$$��"O�u#�k	W���8���\5C�"O���E���A��m@,0蒴��)��<�a�(r�a�LD(��U�b��|�<y��*怀���7K�1�HB�<ك�h��A v/*~���Ŧ\d�<���Qg���L�	������w�<a6��
^� �C�Q
�b�r�k�<	�Ɏ�,��	r��
iJ�!k�<�c@�4k�%�孁0��ت�J\h�<Qr�[&%�4u���ғq�Pt��&c�<1d�Ȑ6M�aLn�B����E[�<�%"ۼ �d�0҃@��ݢ�&OU�<��@�2~᮸@�f�"58g.Q�<Q�.^~�C��C=*�X`u�J�<�¤�3x[�92$�\����
���C�<��	�=m.�=Y#́"����&�f�<��nx[�L�rb�?$t8�	��NZ�<�� �@��3�	>uzzX�T�QJ�<Q��`����A(=���D�<I�O��Z���+7劖L��UQ"��[�<I�����훥s��s"Į*��B䉆V{�����M�(t����M`C�ɬa�4��MN�B|
g�O�u~B��<K��)��T
+�8�S�J�=q��C�	�;�p(��/YP��r�Ga�C�	d�b��h�f�"Ys�.
MjC�I��<Ӵ�!�`��{�6C�44��J�h�)H~]�w+��F�C�	kv5��Ȅ�X��1 ��!�$�I�ِ�M�-��x+B�C)�!��^$N��D������]�!��]�!�$1~�T0BH�-�����2>'!�$_�l�zDB����]��6��#�!�$V�*<�y!���.Cl��U��}�!��&y��lY����9�C�*W!�&A��h����'�5cԇ�( 3!�8aP^M���M�9���2g��<,!�D��f?�ղ苼�e��9�!�E�4�1�l5'T:��q���4�!��	?��غf��a���Q��^�c !��po����Ȏ%�2庱L�5@!��%�A	X'c� q��L�5$!��
���=x���!���K� }!�/"W2�Hs�Ĕ9�d�y�'�!Cq!�$@K��s�ϸ}9ƜC�F��]!�DK
\����DC�F/~U�#��kO!��G�T6��ծ~p}(��#4���<!�l�������Se��y2���
e���y���[��՝�yrk7+�r�k�oH,_V@��N;�y�C��F݄e;��@!{ht!YQ+J�yr�])p��]	E��d츐��"�y�K�4|2*�Ѓʆ�O���:�I��yB�=<����-v8��ر#��yO��}T\h�� 9spz�����)�y��;D�H�!ƨ0h�^m�E�ɧ�y��38�����g���k�9�y2@�; P  �P   >
  �  �  !  (  �0  �6  4=  �C  �I  �Q  X  B^  �d  �j  q  Qw  �}  ��   `� u�	����Zv)C�'ll\�0"Ez+�D:�Dl��b=O$���'h4�l-�fdre&ĳQ�-�I� f
|��aBHX���c�HdI���fh�Q
`C��?��O��?!@�K!.�YpNZ%([��ʿ#� �:gkE�"I6I`��٭l�s�	:�u���\��D�'�py��$�=t�tM�e-�[� uI'I�{+�ő@��O  J�(m�A@Mܦ�aG$Eן���៸��ΟH�bl�3v�Zd��� ���8`�����	e3�-#�4��$�O�+� �����r��3�R�E�؈!��9D�'(�O����O����O��i�+�Ou���'�d���w#_�I�p{��վ9Jԝ[��%�OZ��+@ �;%�2`�������'��듬O��2X�|iB�?�0�n٭4�Ft�UA#g��0�L�O����O����O��d�O(���|j�wI4)�0�� h�L��aZ+X|���?�cz��l�MK���?A��T�?���/�?����31�x���d"�����9#���a��Xܓ���;@��0f�E�8�|��U)\�Yҕ�ӎc��!��Ɉ\-�7-���]��4�b��h�4HF]�GRN����{�,}��k�z��3�i�n@kq�$/�(!a�
�>x��*ՅL7��u�Bir�Lm�MK��-���:�'�.G�1�Z�^���ځ�)�F�Rb�i�7���)�0�tI�$X�.��t2"&׶|Т,��(�)�R�*���/�����-ʊ�B�3/5�M�ѵi��6m
�O��dr�
D�2A챫��V3kQ�1V#J�\0�I���M�~���"Qަ鮫��(
�O�"ggf�sQ�0���'��OR���.�R7�p٧[�]�Tc��OR���Iҟdc4�۷�M#ʟбæ-�U��ŉP��	��'��	�x�	�|���>GQ���f�ʟsk ��ɶ<�X���J�k���T�οa\>��ቌe*t��.Z9{��3�GBß��h� �,�tӡ6�9�ro?Op)��'�B �<!BB�c�0���t���Q� Vӟ4�I��@�?�|*�'ئYX�뛬Fv��S�J�9��:���i>�
޴%�x��W��6�$�+�Z�An4t��	�?�ubء��'F�4o>@�x��d�ɂbT��P!.-0/!�d�<_:��0�&!7<U��c��!��R�~�L��e� ,$NT��B�d
!��3Z2"��Ѹs<��7ᜮ�!�$ֳ �4���F��Q<�8��Ғ=�!�ě̤���+X/�5�"�>�2�Ֆ�O?1CD���>�-qP���d�h�Ηd�<	���� դ\��a���d�<���6>����ߜI��8@&��c�<���5����̔0b�TI� +�[�<���I>=(\�[����H��V�<�@E����tcc#�'DK� ����Xy"bR2�p>���Ի9�P@ѭ#d���e�\�<!�%�*E/�T�TD�݈c�I`�<�-+�^0s���3/ҽ�\�<���sP�Rɇ�H�֭��oYY�<QWm\�A�( H[(������`x��p�l*�M��O,���cC)wDp�X��I#M��ʲ�'+���D���|���Lkȁo�?x2��`���赐�M7/�fE2�OL,�B�@Ó T��U-ֲMH��gDfӤD�>*�(�2��phnI�'C�Y�����"��'��7��OڈQ�C5)�T*cH��e�dJ�ƿ<	�����(�H�rh�|WD�b2cL�2�8����O��}��i[�I���Nڼ5�G��L�h�:Oq� �O ��u�A�E8����ٞ�Eh�M�9�� -a��v<��y4��� ���Ə۷ARlH��U�Й���N�~�\c1�5@+ ą���J�<u#@�pu�H�>��ȓRV:����Y�G�h��+�-5�	�ȓH�q 1��*е7cحf�=��4��O���C���?)���?q,O8@����'Z���tk;/,��@[4`Ű��@C�Oā��D�Os�˧�O�9IT-��-��ԏ�R$$v˞�p��p��K�u���Aՠ�n�1��eH�L��~����ٔ��ܭJ�Ő3��2L:��e�<I�.F����|�I�������e��	D�*.�īU�/}/|���I���'є	��C<M���WᄱYL<���?)c�i&66�4���	�<!�f��6���ii�٠���{<6����?1��?9��5�.�O���i>���:�(�O�\z�iېi�s=�C�ɞ'���SM�?�
��Ձk]��b�>��S��.��a�s�ƭQ���� Ȍ0���d�b����#����(�b]/5��X�e8D���'g^�8Q|�
� &�l�!+�d����&��{T�:�M��O����*aܞa06f&l�HX3��'��۟t��ӟ�R�d��T8R!� �?$�С�S�? N��M�'��k�&�|���6�'�l�XԮ�8�Xp��&�,�y��Y�8B���P+.�ͳ$`�0< J������Jo�Թ �ٯLBv���L7D��1��	�`�I�\��ߟ�&?9�<!H� aj��%��u�l�9c�m��,��^٘d*�@V��5 v��YC����By2��FDF7�O\��|"����?���U F�T���yǆ�۲.͹�?���W�Jܱ�����>�s��|S|��#Ŷ4�ʙ��/Ng~ң��O>1[���.V���p��!P��8�O=?	��֟h�I>E�C�7.���H�#)\e�����ym�Z��T	��P�^i�P�D%�O��%g���JT�N`6��1�X X�+�/�M;���?y�Y�n��I��?����?��yl�M�g�	t`��vOZ�1O�5�5�'������0M��8���L�	�R�8�y�EA��0=Q��� � h�	;FP�$��Hׇ��ET�<��e�g�c�F��SNK-r Ȅ���	�J���]��!��R���p�W�O,�ؽڭO�0Gz�O��'��M�� S�,�$�Q��n�,(j�/�*����r�'���'�R`s�m������ɿY������`\�axuN��1��܉5&T9 ��a!�!�d�(�$ރ/xb�
��[�PY���B�շ90�Yዶ *hm0�:0�a.ѻR�&����U�>]1�1�4U��O�d6/��=��OW�(ƢP@��CՌ��	A�	ϟ�&?e�<i�
�8�顡Gހ|8�p w'�gy��'�6��Oʓh�غA�i��'6�ah�^B��ơ!�����'�r��'l2�'�Bƃn���ʔ�>q�w��	��[�2�(��@%����zÓN��18T��9����`ہo����Q}�` ��۸���8P*W1�0<� ݟd�ɹ�M��x�b�R B͍S8ܱW	Q�x��u�)O~��=�i>��<Ʉ��'[X֨�H@3q$�Y H�Oy��'����?3�%�h�CT�R`�5y=�-�I^y>��7��O�?ͻi�+�A�/�b�)�*h�4���'c�ñU��'b��I��|eB���R�K�^�uh֤��a��q����s@������3�h�zp�$ϰ8mL����ҋ8�]ib���S��O��o����ON��2�J,�qH8�f|RG��y� �"��'���'����^��@rG�_�zb��5��j`�=A��@o��uy�>�Z�i�iXr����)�
+.�q��u�8�d�<	�-�:����?����ē%�Z9s@C�41�����>���~8�åzџ�Х[Ǹ�cu @�(�E0���dj��F��&�Mc`��?'��>c���R/�;4B���^ @w�)!4��Ob8n�ȟ��N�l�|�'��011��xU�@ �q�@ɇ�ўPE{B�'0�h�U)W$�X`���<�|0�@�'��g�>/O|��<�
W@��f
_vZ(�0�@�T���E+<b��'��'��	o�'B�Q�Pn	F\D��N�.B����Ϣ;ŤqI��N��`䜆7>LmБK���yK8'*�A��Д-�0p��'rLTZ G�y�P�.�l�v財�?!��~����'W�	ߟ��?!SFҏ���r��0�8C��H��?���d�O��&��8��efB��}����8�ʓ�? Z�8�'Z�� t�|�dn��a3F���XI0�]??Ғa��Oʓ�?A��?�k	8etL���ƭT�I��'f��C��-�ܰ�]�f4Z	Ó{�����d��h���#fG����o�P0�V�Z�6R�-�#���0<�����$�ڴ�?y��m`b!��4XV�2H�(>�rm����?I���?�����'��'��PӰi�t������>6�X�r�i>Q��"'T`�U$X)8���X6K�5����ByBL��06 ��f>el�ßd���+e�q�f���b0#��8�I� "`�2#�43����b�0�zfjo�%��LЗ3^qH].�q�'���82'mkZD�g
ȑ[��#}Z��<Ȳ�q��!�`�'`~�,�	�?��i�7��O�"|�7�ThhP�Q����u�qP�B\�۟���]����b�]���&O�-0�X1�,�hOt��Hᦩ�ߴ��R��D��e�,6��(}I� HC�'��=�G�4�Q��-Lx��u�(��t�D�rTC�	 9 $�Q+͹WX	SA��g�6C�ɟj��PЃ��ؐL��B�`3.C�I�<�h̳���'V���rm� �8C�ɪ/4p�A� �Tk�dh���
E8C䉿x�DJ�i�h��ұN�ʓ~�Zl��I�l6����F%XD$�:���%X�B�)� H�0Ո
���q����*6��"O諗��;P-N!�G�%.�ly��"OV܉���\}F�c.i��t"O(xZc��岬x�b�y��l�A�'A�K�'_�r���(A����QmB4_���'w���5��:m�J�P��!+��-��'��ջS�Z/b��Q��*��2�%��'3�͚4#�$��ū��C(��c�'@�`��m���Œ�! 9?,���'���� I���#ũ�*t�S��� K�Q?ap �>^�U)#��<S8��Մ*D��AR�T��:�gdS�@���;D��+㋘7R���qE�O&g���ئ�9D��#&�?e:�ۦK#1�0k��6D���"�] "ۊq���C/y�&U0T�5D�Ri��F���Kz:��X7M�O8T���)�qo�x��%GGLZ�R��#S�B�'�ⱉ��`���sa�a�tz�'�����@�Y�*hZQ��n�|	�'¼[���0eu���ڭI��A��'�.use�R�K�� ���>�-
�'d�r/�9 ~��F-1�
t�)O~"��'3�3���w����`Y]ux�'qfuh��J�k���ؠ�!@B|� �'��$CqH��O1rE1� ѮF��;�'��T�V�'"i���G�7@�$|��'n�Ħ��/&(�奜 O�\a�0P����p��qB�w����M��i�ȓ|v*1��� �fj�9��l>����:ā��s��8!3&�0�ȓJ��Z�k��^R,!�m�HU�ȓ\沥[���� ���Z�	Àޤ��ȓdR V	�w0�lKE*�,V�������~�a�ۯ\.�@SSJU `�:a[��q�<Q�Ꭴ	7hY�צ� ���oJm�<yV�\��@��"zz��Z�/�q�<i�N�719>�S�̐�1`j	 ��Oq�<��C��HO�!�W�,~-�A�bhp�<ဏ�=Ք�Pu�&�T���$���6�S�O���B�V�=�d�:t��\�8��"O���$O�x|ppv�̤d5�Y3"O"�K���qn���l��nLI�"O����@[�$���K
!��)��"O �h#��\z�h�
4��pY�"O|ܣ��U0;z0����B��@Y�:9�OR�� ��)�T�1'습%F�qg"Of�P����z�0�ǆ7<�*"OJpy�_����o���#�"Ork����>u��j1/��/!�ĕaoR��!ȁ�2�B|ӢΙ2|-�}R!F��~���(�,J�k"_�Z�ڡ����yㅼ��S�?�* ;�����y�Eu�D,���73��أS�@$�y��L{�K�Z43�^903�ӗ�y�J0_���U%Ր�ReO�y��:d�B<�R�������$�M��hO�]�r�S�#K�� C�l<z�0O�M� B�	ZyF��V�@,�juq��ѭ��ȓl�28��ڶh���-L�3Jl���L� -�p ������0����M�<�a+�
%(�
Sϖ�W��*���J�<�d��xc�YG��_��U����ڟ�q�)#�S�O�x<9�O��I~�ś5d�_��l��"O@)�݇Z7f�{�B�%'� 9`�"O� �C�ꀿ]��5��A�;�.�c"O��ZįL�=y��5���h�4�"OR����6yK���tH�H�^Y�"O��QW���m�*�3��))� �{TQ��P#!'�O�(�� ԿP3\�T��Q匬��'��a�e�)J��5	�	�i��D�'�x�2�Dٴ��8��#�+Q�z�b�'�,�* ��]�D���Q�R���'�p�8��;+Ҙ��&�7��[�H�T �4�"eP��=�0Y	N>{p���s#���W!h�����T�[C���ȓ.�(��w���+�|V��9�����_�����4yd��Jd̙Jj��ȓm��d�	�/���Xu�ŒN���R�،���3 6��2�G;L(@D{�n�ɨ�&@1#�P�R��U�p��8~%
F"O��7Jͧ%ELE񤠇.f��c�"O���V�\��p򀏇�`�����"O���4LKe��h3w��d�m
�"O���u��*5:c.�t�0B"O���S�Q��\�(kf�F�O�����)��؝x���2P+&I�x�	�'t\�b2*��qѕ�7G9H$8	�'�z}��mآ,��EQB���@����'�F�cG�/>�z�aV��3�0�I	�'F��)UI�-`��k�C4|�����'������i#<�	�����(OXp��'��T�ơ�.R�T�Q>ek�'� ��wIL��H�$[�/�t�	�'(��P�	/O�.8��M;I���'~<*E�^8 �^�r�1Xl����'���#�휾|r�aab@�8"���A�]d^Q�$��pt gI�T��ڒ��Ԇ�!�h臯�++c��K���!Z���Mo�m���*C����c�@!���sG"yZǯ�	W&&�0��N	I�0<�ȓ �Υ
��רa~��&&C�5����ȓb���4J;&����A>�rmD{BNG������ąO�5LX��#&��~��9 d"Ot����a`����]#k>��"O6�C2���;E���g�lD��qg"O$�ce���M�� d�̨�"O��t��E� ���I�d��˒"O����D�X�|��B�>e��Ta��'0��p����3��4�F�\�#Т<�.Y�� ��4�6��fDٱ](��N�_�����r�"�A�ʋ��CƖ).��ȓ.���rJ['��XBJTF�=�ȓ2PT G# �rZҬ��D	(Kd	��?+x�+�d��[g�]y�ؠ�L�')�`*�8:Zb5�/-*�p���Z���Q0pX�ЌL�"�"��q$D���4��z ���夂-��u
��EI�5�ȓ&89Rk�2R�.`�w��@�d}��(a�ᢒ"D�vNм����M�,؆��2]���2;�,hK�$eݨ����؋p�4C�/1�X��$F���b��#���C�	�K�*�{�0>P�S��d�"B��j� i\�DY� ��/�!z ���'������$
Ҷ�Wc�9w�^�b�'D ܃0�-�DTs���+u_@�ڍ��ȮQ?YA�ܮYs�d���.NKh$[��6D���&���|������.%2d�E� D�<3�e�w%p��0
-lz2Is�=D�� 2��ՈM�,\�]�"���{}�!A"O�రǍvY�� B�|z�b�"O���pn�:j$+Q̎!,o�!)�'����ӹE�v�Qe�T�]��"�K� ����ȓ�P�2�ʕ5z���b�?iU��ȓ):���q�Y 8s�A6�9oT<X�ȓO���b�PD��H�=8�L��ȓ@T�8���37hpI�'��Rʎ����b	
S��P�*E���V�p�'���P�y=�4�`��!
�����L��>܄ȓ�"y��B��B�stiP� ���ȓ ��|��*@'Y۪s�L�<9 �%�ȓ|Ph�	��ɀ.Ǫ=��d�G|A��lʮ;��5k�)�d ��GL08��I+8���I��,+%�~!ǀ��:Ҋ\246D�P��fI�+�,�G��$�v����4D���%O'`h|ڳ+�"��� �&D�LS�m8`���b���2X A��h0D��R��a�y%�\�g����"/D��C��#
|�0��- �A|��E.ړFn�D��̋k�D)�'RkP�1f\��y�#B�>���!&�D�h��T0��J	�yB$Z^�d���BI�yЏ��y҅�,U�0P���IL���ׇ���y�d�n�<u��A�
P&A1�&��yBf$r����ub4$:�Z����?�0dDD����ȑ��� �^�j���B��`8�_HB�ɼ:��z࢚�_&:�E8C�	�?�ty�	#`��YdB�	9-X����A�_c���֮�.6YB�	�xN�C�G*O�e 6oL�u�C�I(A�x\�ah�!<���S�-`� ���z�IÜ�̓@=N�H���O:"���OV�)M�jw*�#�/+K�-�D�ކ����K�l���O��dZ#]8��'�6;f�c�%����w�z��סL���	p����y�">y��d�z(�� Q�1��,j-��(:�K�c�i��ڋY��]"#�	�Dg2�d�O�c>��V�%.4�����_�����<�����(�!^�Gk�Y�H�3;����I���$�K��%��a�|%x�����Q6�Od`y��%�I�?�IC)���תH"�2�aTOX�FB�	�ڀ��',ԇ#�]Z5�T,x�2B�	1O5
H`di�9aN�]�פ��g��B��7T�h�oɪ{+�	��.�lC䉞@���K�ׅyh�U�©W�RC䉿_������E�~��"a�9  �����~���*(��A��7U"�!��fV�y2O��-������I�(y8����y2k����Q F�>�,�	u���y�f�.r�i�:�٠D���y�D��{�F}Ce��0W)�'!�y�ʔ,J��)"4��'3l�dVg��?Y��D]��x�3	�BX����H�C��Y�1D�h3D��?p��L{�oT_�T�Ƭ-D��2�R�0�f��g"�"doV�ɷ�*D���d+�QF����;V�Qa2�-D�X����`3J�Ʌ�3n���F(|O����>��%>.�\�PpFDW�H|�aA�D�<9�^�OR��r A�*#Z���|�<!$M�0[֒(�cJϋg\yђ�z�<`��64�JMQ�O�weنMv�<y��P�0���P���ޕ�ITk�<	 L2Q*��`�ݤJ�(�iBLj��I�vTDxJ?����	�f���J7P�k��32D��b��ܐa��N�Z��A��*D���&C�B���KVɠ3i�����4D�� �	R��1*r�U��C��<f���"O�e��S�9(�R�,V�N� k'"OL�F�Gd����KT�!�b4ZC)[��O֢}�&��y�n��O�B�����'4΀���6$t���8	��5��#�4�|ćȓ^��,�A��'!b=ئY�E��,�ȓl%
s��i��Ka��:V�H��gp�Eys �(n���3s	z���vf���΍�s�NL�TM��P�.��$"��D��R�Y��e���:�d�,t!��P�R�0@O�y��-P��28�!�$�>�.�Z��3(�dL�A`ΆT!�_M�L�〷B<4)��{����'�
e	���c	�Y�#+� A��B��d�f$�!l�_�	�a���ȓႧe2���o�=!#��'�R�'��
!H>��So�Q��H*?O�遟++̜�Dc4T��9����?��pQ`�	�c��l��,Ѣ^��'a����1���4�v�s�0q��1b���` r�'��'��iV�@��cb�5!ќ���"�'/2�'�b[>�Dx�*R�1���F�5g�@�صK����>!BT�$H 4�����i'�XIu��<q�YE���'?�O�Ҕ�`p��K�3���ӷ}�+��O�ax��ɜ��CP�ĵ$�>�@^O�HX��Ҳi��':�u$>Ms��*���1�٣Y%�<9Ъ\-�M��?F�9q�'X�S��?)���?q�'�:�b�A�J@��m�>����`U�*��&�'E�����'��P�r����u�o5�1fuF�I�k�fDjf�@;ž�AV'�O��F�d�
��ݺ���?Y�'�?�'K�uIS���u��#B[V�[q�Ws\,���O8
$�Ox�ɑ-
n�s��N���N�u���"� ��g��
7!�?y��Hߟt���pJ����OJ�I�O`��vʈ��D1X��R�dv<��oHП4���OR����}���h�$�e�?7��-��/�2a�'�J�d"��H	�:��l�<�q����D��>Ur�'�?a���҄� 0���8pv�Äo��t�|y�'a������?�׼�@��x�P��/�?Yoڈ ����k+8,�X�V�ƨQ���ը����Γnnt�I��;u�2���?Y7
Q�_c��!�柈�"��Ȃ�i��DqT:O�@ �'�r�O��1O ��;��`rR��B��@�Z�x���qӜ�xb#�O���?��S�g}R��v����&��/W�P�+A��y2�WV0cȟ�xp���@f� �M����?q/O,���O��$�O���{��Q#70�Qr�ƹ<@�8P�ݦ��ğT�Iӟ��	����ȟ��؟Lj�9���rk�7ot�	2�j	��M#,O��D�<�L~b/O0�iSOC�)N�p*$�U���S�,�ߦ}D{���i�6�r��^(�u�E�0f�����O�����g��C7M�I�$�P��<?!��O,^�TY�8�衐�KM�,&!�$R)RA��Q�� /Rxb,�3�\�!�DEp��8kpNZ���^�!�$N&_�"�%�>6�E��3�!�d�:#gތ�b��5�(�b�ۂ<�!�dT�xl���ۿH$Iqt�ҼJ�!�����%k��UeJ9j�!��P�tp�$��^؎�e��z�!�R�0�^�C��N�r��CB^'�OJ��B�$Ci���&	�o���h5&96|8��G*lf�1�:o����.Kd&�w���X1K�Ǎ�!�� ��<@{����	�xyq)w�����<Q�����a;��
@,R$:"�x�QDZ�d�8�����-5���� e�$1N���L3RSP%'����{�[f��huT5{#��hm!�䒸y����T�Vf:6�k�@\�Rf!�DZ�Cl k���3���.F- s!��+�f) ���?�p-d�!�<GJوd�
hhZ&IQ=q�!�$�Xd��
�(�e����gv!��b��jr-�w�n�W�	!�DC�n��pS�f�B��)�,�B�!��K?" >qHp̉�Ԛ�ѩ6%�!���p]D�h�E֙5���
�S5Aq!���+c���Q��Ǿ�`p*s�V�	U!��uZ�� ��.�P�r�#[!�č�z&�ųC"A�p������mQ!�� <4�e�]�(��C�� BAh�{A"Oz���2@D���7�f��"OP�B���#��%h���xi�- 7"O�ygݪ>݌$�MN����x�"O�ݚ�k8J|V�i���S=�4�"Ot�rD�Z��Ĩ�1b���2P"O�ec#�I��H�,{���E"OZWA�O$���ֆ�7UH����]�<�B�'5Y�A�g�7~���TG�p�<�w�ؑ7v2 �FU�f��heHj�<�䎎UB\�ᦉ�}C� �G_}�<�0 �)��,;ufX�`�!��$�a�<���q��: ԮU"�M�VC�D-(�pv�96�R���� ��B䉮��	�#ԳJN0��]�&�B���a��)�$݈j���g�.B�	(R��8���Q�̊1I�cg�C�ɜ<����`C�ǎ$����L��C��L���Dn�1��(BTF��C�I�R�����-�Iy~��dfѰ)y�C䉞f�(Z�"p�$��&�*7O�C�ɝg=��3%�K0o+$� ���G�vC�I�<xi��)i#����� �6C䉙��U�Í��Y��c���!�C�ɻkE|�S�?|�+0��-�C��#���S���4$JX)c��D0p��C�I�j֘@zL؀j���8B䉍v�z�΋B��dG޹MB�C䉠/�TyK�@ڀÊ�`��>kpB�I�ze+��)�|)`T�V�n�bB䉰~���[��L�@�N](Qc��V <B�;&�1��	��̈�mN(8B�X�l�1�M�qJdH!&4�!�L!=��p5�Ğ T�ٓ�QN�B�I1�����*����1'�)x��B�ɬRm���(�S�ԣU�R):��B�I�dЪ0��OŦL��C���1-�B�ɬ]�Ĝ��e]�b���hԂ͎eW�B�ɸ�d��G�6l�a�ǌ0s�C�I� H���&��9��=�V��T�<C䉡S�ޅ�e�_�2i����_�3�C䉋
HI�e/��.�tI�u�ސ3-�B䉉F��҇��.K��r�+�zB�I��uy��/m��-�sI;M*B�ɌPx��B�ٛ@4�q�d��#lB�	�3IJ��W��w،	a�*"�C�	QdӖ�F�^`�ͶC䉒R��}�rCέ!�Xu�N^p#�C�	�I�(r� � wF�x�n�q�~C�	�4ܚ	sG���PJ�1���$NC�	�;���b���/Ba�)�~�pC�I�/�|̋��S7�Ҕ"AE� W,B�I�#�q�+-ۜ�*���%4B�	�WjN�d�i�0�BŬ@6PB�ɽV%|A�q�C�G�3�,�6R��B�(%�j��pI���HBc[�qhB�	�DdT��g�@�o�ѠamU�?uC�a�Z)��%m��H�6!���B䉈^�fJ�/ֆZ�3K<r��B�ɊY!���sJY9C��RPBB�I:4��U�+Yd�
��E�HB�	�v�C���L,��b�B�4\C���Dk�3�(�G_���B�	eB����^��� h�e�zC�)� �I`&j�>O��@���0-��5�"Ol�P����d�ֆԹ,���"O��#�j��V�4x��>Z�vL��"O,�R�ע(en�贋����!V"O����*'�2UjE�:sr�B�"O9����Nxٻ�L&*p~���"O$���V�f�x#4��_��mQ%"O����x"�iܕΨa"O��i�dG�0�<�e)4)�-"�"O2����)pj�s��"[���"O(U#�*��[�0�ĻR�x�5"O
�A��P�l�A�$o�h���
g"O#'�)K7H�ʲ�Ţtin�p"OJ�t�L9�8D��53x�"O>�҅jZ�t5@XH3BL�'P���"O�%K&-�<r����_�
�l�x�"OVh#��ðN '��n��y�"O��;e �md�X��h���8G"O�ف�%�R�*�A���0O�8���"O�����2?���Tc'$�RRp"O` 6�],P�p s��L��q��"O�4�q�/(:� �!y�T+F"O��ѫ�7�ً�H�Q���f"O�1�/Ĩvq]�o4n�8�j�"O���T62���bS�'��]S"O��S'J%ʸ�H���C��Ń�"O��;C��1}8�����R��d�Pe"O x"lR�{��q'�E�QI���'"O�r��ǌ�ls��Y;�p!�"OZe� Q*g+�DJDH���4�8�'���'h�4c[x�0��Q<�)�'�Z��`��7H�P]hԠ��Ĩ�y�$O�~]��)@`�J΂L 3eC.�y2��=(Ĵ��W�XVG��f��y��Kx��͆?M���̈��yO@0As\��t�	)DL4Qc2���y��QU9s�JK�����6�y�>Kl�
��Jp2!�0O�'�yA3v�$���\ DB&	 ��y�e$X�ò�S�J�1�%��y�'�Xz���V"�,t��J�-���y����-'�a�B�M�ps6G��y�N?�b0a��zrZ5��N��y�#�=7p�,� �X�IB�|��Ͷ�yR+��8�����V	H�1����1�yB���!cJt�F�#J!l@��ٴ�yb�_|-<��$�E/�������'�y2��x5b�����BČ)RC�ɤ1��w#X@��� -`�ZB�	Z�P%#Sb�(*�%P�@C��B��? �D��ڟԶ�öH�0�B�	�F�X*�m�8
��1��+YLC�I-2B�붨�X���Ct���LB�ɞw�R��1��{Z�#�D@�8B�	B��@"�÷@����&@z��ć�|����]�R��e�*5�!�I/&�i�D�Un~	*�����!�$^؄i04�Z8b����.Ģ�!��H�a��
�J5TZԲqO�&0�!�� E���c�';C�a����V�!�D�!��� �.@zY��B�!����8d@@�Č���G�K�!�E�^t,0�8d�n3SFP��Pybk��XnBq��eɈ|��jB����y
� ������K�Vd P�C &�Ő�"O�8#��E4w�L�3/��6=Х"OqpF��+#����J�0"O��Z(��|�t �T��}�VT 6"O������Y	�y:W����qi2"O<P����YdٖC��mq���v"O6�Ivϓ4/�
���kʉ?�6*#D��I�F�;1>�!i�8YjT��t<D��b����S����'�u�c�/D�zթ�:t[6��nE�N�8%��.D����@ DyJ���v	�DL9D���L�|>T|��+�:�<f":D���JCx�p#���0���1@	:D���"�Q�l�������\I���E:D��rc&R�x�@d��i�*D����;D������8P�\q����U���zC�	�g�T��w��g�\�*&+D50׀B�I'J/����Ą�?�v��#]9O�HB�	>9,�9¬['3PŪ�i�	T�C䉼Tў1��h]�L�D��̙�j��C��`���E'Y�##��8�L����C��R?~�*����:�0u�㩈�=pC䉬{Y�|H�I��%�s�9qB�	�)9n=�kؽ��B�E܎;�TB䉿~�<	��i�' ��2��h�^C�	�+�vuc�kS&VMĄ�gn��&^C�I�V���B!tF	J�ə�<�6C��,(�l�G��U�p`��J�+LC�I�	�0dA��#%֤��A�<C�C��e���2.H�z��!�(�~C�	p���۔�[}� ����jC�	�cX����S�T����F�:�ZC�I�_Ll���ψP�Y�	��BC�	>}��53ϊs �d8p�"l=,C�I8��੓�yUL!iA�,5�C�?�`p"f�f�5SA���C�,a�,����~��uxdʟ�C�	��1�NK� ��F���C�I!Je�����(C����ͪrAnC�I4k���M;�x��G��*r(B�	#a�H�2ǇX�ܙ��H,B�	TD���#dB�dQ� ��a B�	�6��9�e��3��i�Xhy���?D�8�T�O�{Pt)��G�� �/2D���gQ2A�9H�O�<'�(���.D�4�Ǣ�r^`9�#ӥ6���ӱo,D�T� �9�j�#��T+R�5��b/D�h�肄wmBE�rO$X�tyq��'D��I'�3Vfr���7
�V�1��0D��; #ӌ|0�1��4	��0��/D�����kb6�g��<a℠��"D��꣤2�*���I_��=���?D�l[�dU�l!`"�
e��� v�=D��җ�C�.�M�G��4�&�A�E:D�X �'�#*}�zO�u� �zu�6D�TKf�l��lCR�(p1���c6D�����-g_F� ������qVl4��J6~8*4N�,��9�0n�e(D�Oʑ�dҽ	�Xh����o%~�9�"O����)ؓ^��8��@�'0X�(a"O�a��)&Z̕xӈƕMGd9	�"OKǘN�*}����&yQ�I*%�P��yr S�FQ�7���{ނ	��O	�y����%��\`�G��%��2�T��yBP#0���K�ɇ�q���ŨG*�y
� ��:��U��!�U,�Z�q�"O*x0���)&"-���3�F<��"OT�HSg�z�,����:��\��"O� ��1���0K�0�K�"O�ԩ&.ܼO�X�ʳ���.�5� "O��##bŞ����ᩝw�x��"O��x$d��|�J��$�Y�qR0��"O�ABPG�)ijQ�]Wp|��"O"Ѥ�l��}0�GNk�<۔"O4�)��O�:"�h�/R�#�Y�4"O�P�����h(8�֮���H)u"O���_}�h�RNCh�@30"O����Z9p<(QM�>P:*Cs"O`��\���z��X
�� "Orl�ēJ��	��Ѧ
4l��"O8X���9S(����+�D���"O��1!�k�������l����"O.͓�M�Ѝ�q�ܜ}c���W"Oj	���	�rd6L�郩V1Rً�"O��$@MC&iv��&y�y e"O��bv�3N$�)��%q=<���"O�����d���!p"Q��<���"O����ǔ1t��u��m�LE` "O�Ys�e_46b��U�Z+r��U`�"O��B6
I>�؀*b�%/��9�"Ov9PA�|�;�JUWV�H�"O���g#J��Z��&��R"O �q�N8����֏�/��"O�([�Gҳu�\��6��t�����"O��8W��8�<{W"Ī���X�"O��D��4p���W@S�R��"O����� �E�F��צ�P䀡Z3"OX���U������9�\�T"On8kk	�t���z��`�6I�"Oz���G��]�B�DP���S"O�xT�� $Z����$|A�"O\ⷩ�6
n��R �Xt�t�2"O�,
��P�~ m�
 ��Hc"OJ�	����Ia慫g�ޤ�t"O�p�b�����P�Ф��L�8a"O��8qj�C�쵛䙏VQ$M��"O��Ǣ]�+`�RT��T�"Ohm��@�j1���X5`���jT"O 1[�
�5ftPD�Ս.�޸s"O��0�6 5�  5ȋ82*`��'"O��c�
Dm+&�1l��R�"O�M����4��$L�,�N��"OY� '�Hh��d�)�R5!"O��q�\�B�v�V�%jQ�R"OR�8���D2���өK�{fhQP�"O����Rڤ�i�.VY��t"O&�
�m�	?u�D"� ��9�"O��֥��ǬA���Z�M,|��"O�t'ϴGڢ J���zo(��D"Ox�:���-^����ڳHg���"OpՐ5D�b�T�O'xIؑ��"O��BY�cz��u��5U�x���"OБH2FU*@�v�J�N�)|�5"O𬰡�6T �fK	6�B��@"O��ڥ%�g��(��G�N�)��"O�({7�CX"��; F	~yQ�"O��q�A:T�^���YL��"OP�bW�םGZ"!Apb	��$-�"O��4IEd��tb$Dܣ��l�u"O� 0���	Pr���t����"O�T���Ԭ]H����j�X�� ju"O�P��^/�|R'�T�g��5�u"Óa�-��K?nu�@'�3z��r"O��z��ܠ��9��e��!�G"O�����P�v�{���:Ԋ"O��+�o@�^�`ݒS�ߴ�B�t"O�Ux@�(Fu�ԡ�z�q "ON=Z�èLђ�� C��iXX�(1"O�d�楘O�P�7s�6(��'ԺxjbM�D�v]A�鏮S�$���'�\9�L],-�� O*I�\�b�'��d�9��A���.|�\qK�'0�Jǋ�q	D���ų<#����'f��`Den\pD�<Y�%��'�5�De�;�Ptd-H2�� ��'x��j� ��a�v<����)��x��'����i��ZoS�+��I�'�F<B"�]Z�dBOU�*���b�'�Le�a�ݑ	��-��Bӏ_�؅�'.��b�
�4�蕃s�T�E
伂�'����'[W�*`��>�l��'�tQ�q�G�d���C*S[�v�h�'vB	�����7*�˂�\�Z�b���'���I��P6OT|X���)w��s
�'����R�p1�5S2Fш+�ܙ��'M�8��nĽ&��s��
]�B��	�'����e_(6�ɓ��(T����i�&�(��*x�v����ۣ[!N�ȓ�n�I��ȪC�rA�t�����h�ȓ �~�)�KB('��I��;6����{bP�$nԶ`h�H�d����&�X����0=� I1Y�*}�c��0>Ǌ��AMTk��آ"�E'z���"+�-\D��W\{���(�xBKN�p.,�I���<h-rU��HO0��!/QW̥IA�D~�''/�\��A�	|@�ƌe� }�ȓ!� �1�L˃o�ZV��=���l�x&�h{�� K
9��O?7-��6Z��e�s
fiSe鄉E!��G�~�h�n�	�RmCg&�?^�|m�8}��0�H@�-h�e��h>#>q�BY()A�M��HJ�ʵ�Eu�P�P�hr��r�$�3���ڠ*���� dD� ��(3�L�Ͱ?��O�_H�����;F�]H�nW`��KI��pÏ<?�i���x��������*#x���3�#\��#"O��R�W�6�aQ"���6DFp��˙u�~�d�	6eҪhhGl�j<�>�I�;Zj$�el	���T�&%P�B�I9e{:��� �z�\��T܆a�*�Qڴva#VG��>ʁ�4�Nź���	d��pge�T&�Cw 0�����ڄ=h��>pHF��J�2?g��aW��, ��:�K-t(�w~����և�UlX���`֚!S*�p%�)�ɴJ�\Hb�J?V�V�cE#��7�?#�O�Dr��oS�
�����6D��`s�?8%�f�������.vw@���)A�*�&�Z�c�1�MG���w��1��F2N�����Q�b�Q`j4D����_����i� 	�4!��`�M��c�!_>� ��$r�l��Lb�o1*Eeڇg��9' _�=��{rNJ�3��D�'`J0+����E��55�Ĭ�$N�!gj`[��Y��YQ�'�d��V+�5B(pi�a@[�U����?I�Z�L�
s�F+P��4ːV�	]��N�{�m�0�֥3����^!�I7@�pD��f�
 \��4凒}��I�w�Q�"̈́i��7�s��k���B�\��w�U���"�+D���*ڎp�ƙӆ��/1����e���D?������3�IuB9����� ��6��4m�>��D���l
�� "��%����{6H��^��  �'��d1��(Z�l�uD�>C����½,�f��M[�81�����n�;&'Pmrb�d[X|�"O� T��E��>(o��0�cX �lQ�q�O�@{7E��^C"�O�>c�!�
$��)*COŁ'K�H�fl'D�̢��=f~"4���z��E�l"�$>u.���	,�L
˿kc$����4�B�I�H;X�q��&A|S��V$��B䉝�4p�-:C���AgGY�C���� QĜ�W�ڐkF�Fi��C�I?uʈ�ᕏ� ��xQmɰby�C�	B����b��l"P�;\�C�	 '��p6�F3�F�(6�9s�DB�Ɍ=):a2`�V��r�3N#�B�	��LX�E�)"&kS�B�Il�
�����
 W����&N^C�	�(ҍ�Tm�N��Ab�CC-��C�I�(���yw/��,C�	�$l�(%��C�I##l+wa�� ��e�'N��hB��+ʅ�e .��-Y!S��q�%D�̺p���̃dC'p�����!D��b�̷,:�ꞆD�pqj3%"D�`k�A�'gf��)�#^+Hq�pX� D�,����2��Zv�ߌN��)�'�/D��h��V���%^� Ji�!0D��"D.T�wU������-?D��@��{Р؆�M�bU��ʅF"D�܁s���p��g�=T)"�;D��۷&�P-�&��r$� �-D�Xj F�{c8�����p�%�%)D�(�,�F�ȥ�Q���V��-[�6D�(Aр��[���9p��/)D��a�@(|
��t
�	�4�1��!D���vO������(L��C�1D��s$
0�i)d�͵a�2���1D���Vl�|{�A*'�kd�	ӧ0D�t�cdʽ7�8E0dǊd����i$D� �Qg��_Y��c�`�qSf%�1 -D�p9/J3lր��)AkM>uB�a)D��t�" ��]�7�EZ��$$D�Bܸ97��c!L��T��B- D�(($�βs���qC�W�Q���`.D�H�wo�8?���5)�{G$<�1c.D�F�ӲHeܬ���
-�  ���&D�`��F��'�J�1 �Z�X�`'D����K�����эǀl�� �`�:D�0 T+�B5J����*���Y�'D��)u�]/U���7��nq#i%D�XP"l�65%t��5lʋA} ��
7D���E	S5qt�{�Ȗ�-��%�?D�0�ᆏ��
�K!���o�@զ=D�|���
b�|��ע\�  �B/7D�,�R� ��a��}�LG5D�D�Db�w$ (�C��04;p�B�/D�$�0��0����7?�J���#D�H!ei�7f�NP�bA�t�0�*Ţ;D�����	��\���X�/.�	�D)&D��+�*atL�Ŋ�%A��գ��!D��qw��%v���,D~�P� 4�4D��k`�ЫOo�cP��>�N��Q1D��	��R�N���!�H�m��S��>D����+u� sy��m��:D�\q��Q�.�z��K'��УA9D���V�P* ``t�S�Fql��׊&�I�v��jG'��8�"�S�ߪ�O��P��*T�2�P@�Ŵ�Ͳ�1D�t@�瘶?�p [��T1 ����$D�,8#�	�@RR�HBV?	Gi�R"D�� �XfM	#,�0��Y-O�<=��"O�3�-I��UJ�'���R�"O��墉�2%��I�� �?%@�f"O��ч�U$?]�Y��%���B�c"O�X(�o�5yض�1��;
��Y�P"O�����.N�z�0�A/x�D�"O�0�"P#M�y�! &_x�ه"O�+V�ԟh�Ȉ�CgN�\Vp�"O�Ha&� W�0!K6��0O��"�"O� �ϕ ��a�	�0�"O����̷(f�����\7���'c�!�կ!w��C+Ia����'��sV��0B`����f�Qq���'P�L�V&W9�.�Y��]�NZ �	�'��Y���S�-N>��L=u��U:	�'~�5:�%U�i�P�EG��#�.�	�'���KflW�*��s��̩`�R	�'n5��G��Ζ��28Q
�'U�А�eI�M�H�$k���V@�
�'Nhm�t��%L�Y�	Õg޴�	�'V���D&O=n>Az&�$U��	�'�F|��ϐ�P>(���J��H�ze1�'= �*վmbxS��_#EX�=�
�'����D��M/��8�(��K��+
�'j��b�$��r��8���*H
���'9:��DA�:h�ČE�X"�̆��� �w\�26�qx��F@���"���S� E�p�r�a<m0�ȓ0m�Չf��:L����͵�����m���C���F�Į`��y��.�x� ��hAz�@��'|�0��+����5�@A<ш��Jt��̅ȓ}S� c�[�HR�y w#������ȓMk	�N�*B�ݫ�U;�,	��I���B�K�.[tt�陎�D$��fZ�̠cJ[�Z��!KF�Z��ȓ�hdS(�&VU��2��<��W'z�0� W�z�B�_1|*��.��ۓ):�
�BQ�Q8A��D��+40`��#.~�ʂ K�X$C��Z��4�IV F$a��U2��C�	g(�U(�] uئ�����&itC�I�E�aH���'>o>t+�)�0�B�	�}���#���*m- `�`�4P��B�ɘjT���"kȁP��@�߂.�xB䉫f̊�RDL	F8�=R��B�W�FB�	/@*�e�?i%ܩJS��]]B�	%4z��+D���d�₨�~@B�	�09V՘a�N�X6Zu�U,�7|p�B�	�u�.��5��)uX��W
�w��B�	�jM*�1�n��>�]y�X�-��C�	��b<B$��;��uJr� ��C�ɕq���˒N=|���0�שM��C�)m����9nĎ��Q ԦR �B䉪j��-`�	�ĘaQ�m�-��B�I�?6�l�#��%\��rPI�U�B�ɧw�z�{��ut�r�%$0�B�	6^V�Qv�)[@!�� ��B�	(@Ǥ��jYO�@z@T&q|B�ɷ�n�CujT+C]�`��R5lRB�ɾ5ЬTF�W�M�(��2A�ZB�I|��|��k�? �؝��L�E�"B�zp�a�F�%.�Q3/͚/
B�	�+��(O�a.�5����B�)� "q��וi��A��a�W�U	�"O��ZQ䍨g2���æTY��H�'"OF����MI��	0 ��>D�q"O����]>rX\YI aÀw>8L�"O̼bfÂ�:�0c�G4G-j%"O\�;�JL�]�n�I��x��T�D"OF|�e���8�TCM�6;�6"O<=��Pql,��ЯR/3Ʃ8B"Ot�P2/^�[��"�݉;�j��"O�X��.�$=J��#[�
j���"O�ݫ�
��(W\����>G��4"O�H ��I�2-�M0,U�����"O�9(�l o��1f+Ea}P@��"Or����M{v�
J�\UҩC@"O"��w@�$s$�a�	�%<��"O�U��qh�ǩ	2.8R��"OƩ�Մ�7��q�s�Db��"O��Xe �?���#�'��WPF@J3"O�Ap��'��+�gT?F�F"O��ՌT�،A9 >|J3"O<9����?
�@�%B�m�t�A�"OV!2"@��G�jm[2K���(�2"O�L[e@�NY�U���̘$����"O	�,��r8!A�+��?��]HP"O�]X,�*<�a�K�
H��e"O����-|c�P"�Í7h�d��t"O��
��o�X���h�
O(z}z#"OR��3��#hJ�"Q'�	Ҷ"O2=��6
��4�F�.;�,���"O4]�n/��:P�ؓf\��w!	Y�<QDB�1?�d�C�>��}�E�HV�<a5�؋��� )� �H��P�<1��C;n�6��Q!A?u����sIe�<��i��@<Q�(��e=�T�
x�<�W`�/�hH�-�G��[J�J�<Y@�[�<��E�&�� EH�<����tk���R�Z bZt`���G�<i�O+Vu��`���9��"v��z�<�N52 �K�a�I, ��n\y�<�2 36]$LoS��`��$�_�<i#�ش3� �A����>�0��F�<����"\���3�e�0js>��� ZF�<�`
�!��AA �D�a�!:�_@�<1vHT����h�x�0��{�<����*��Ϗ� � S�n�f�!�dP�`c�L��#�=Uz��E�!�Ȉe�ޭHR�I�q�]b��΂k�!򤟄v(�����=<�E�Əv!�Ğ����z��ξU�Ph��ƸRq!�H%HH;e�׾b~�K����z�!�D1.�8��w!��-�� �/�!�D��[5�y�Ǘ�f�ԅX�FL8z7!�Dʔ>�h�tf��6� @	��-99ax��I=[������Ð%1�J�C䉼@�(���Дdy���c���C��.<2����G�b����]�B��9}�<�&�M$7�U��H��B�	Dadah"OϚ3��RT�Ƙ)׌C�I�T�	��-�kGv���YB�4��ГO��r���U��$C�����a2�ǖ<K����/�$��B�	:��{7�H�CA�,����w�C�I�o�� aa�Z�� a��6��C��>$�N-pB$$X`�M�3Z�B�)� z-2� T4"�
���%i��"O( �lՒ\0u
�aC�k���3�"O�`�D�J;(��i27 ӵnԠV"O�
!��Fpp�I�E3����"O��A�ۭ��!�cF|\��"O�E�g)�/g���s-ٓ{QȔ� "O+e��)U���&B(m�j�
�"O���b�G�@з�Q�5x`LC�"O�UV)сIB��E䖊x[�E"O����'ɟzA�񠷨[�DvRm#�"O��� ˁ�,�,QA�Y5J�4)�"O�h�q���m
ƕS� �0@b�"O��`�ό4.�����i�"O(E��K5/M����b!��A!"O�U�Ӏ�������N
�^!�"O���@*�.�B����3�,�Q "OļxC���Xut���Y�Nn�HW"O䐠T��P��1�%�!a[����"O���#�9d�>���$5X�u�"OP4�Ń@9����"<E���E"Obe�b��y��9Ц�VD`x�"OD��U�|C"4���9-1 D�"Ov��',�!i�I���	R"Rr�"O�y��H�kw�%r�A�6 ��@"O�� �ΆNG�x%ɘK`��"Ot�����$t�Y�W��%g�r-T"OZe���3�ȁ�!��0T,��q"O^��f�^�E�rqDC-/�|�1"O8��`� �m0���a��<���#"O�����u�Fq�t��J�����"O�m��}���$��8' Y�#k.D���I�<4��h�g׌L+
Yb"�-D��Q&�Y�)d�
�Ls3B���*D�����T�
X�~�H�rq;D��C��qr�֭�� �"�Т+.D��;���bF��Ʃ/A@�ȃ�?D�����%)׾9i�
������6!?D�lCĚ�Y��|Je*��
���<D���l�@nܩ��H�Fђ�I��&D����ĕ3s�9��$�o%P�3��#D�� ��Tުݠѧ]�<�	2$ D��[0L�6p$;���<6� �	B;D�i��3���b��`��)�l7D�l�!/k�v1z��H�45D�RU�6�$q�@��Zg�t�.D� ���Z&.��XRr�Q�6��,;�E&D�zZ�`�� 2 ~zA�ĮW�%!�&�P�tcϞ}j,h``� X�!�d�>z�%��̠.`�rb�Q�!��Ke���� I�s�ozs!�D�J��(���f�m���\
!�J~��v�
�no���#��Pybn/@p@�C�<��)�Ҥ�y�+�26>\{'ٳ,�a�UFM��yr�97]~q�D�u��dH%H�"�yb
�9Tt��X��B�9u5���y�N��hݣ�?-U�<KSc�yb�OR8E���*Z�x�"b��yB'O�%ݔ��b,Δnav��ǣ��yb*_.~%qh��H��7넿�y��R*$��˛es2�@�J=�y�˃�r.����DаR\������y���H9gL�4����r�H*�y�����/���Jw� �y
� 6L�d��jonH�L�![�,���"O��C��E�d�
�:$A�x�b�"Od!�!Z��E��ѥ7�l�#"O�q;���?Z�$4�d�0�
Q"O,|�t��,�][FcF3q��m�f"Od�أ�K8Y�����4Q����"O�(��'�H�b��g�e!��R�"Of9�6nT7�`Hd�_� :2�"O0�H Ō*Z-�QPg
�1w[(�"OLpB�ޤ{���F F�[K<��F"OęP@��O�б��o�3�n���"O����AR5*s��1`��:Z�}93"O�=Vk��S�
8��Z�����"Oj�賊�����Sݨ�"O�h���B�KLb�bD#LM4���"ONe�$GB0.�\BŢ�U�3�"O�0zU�����S@�^���a�"OB���b�].(-����F1\�J�"O�مg�Z�:��'-��=\��"O XQ�Ḑm���8A���W�P�*t"O�M�,]36u��q��Wp�����*O��z4���o�FA �L9{�i�'�ْǠ�^� :�ŗ�-�H
�'�:��o	�7����ƹ+� 3�'��j7$���`Z狊�q��=��'��(��'�3"q&L�nM7q�@�' �8 Q��"���&�b�@��'(��Aā&���E��'�����'A�y��-=��Q�X�J<��'��l0��ރ�������O
BL�'
d���۪G<�D�Þ�s���R�'9e��B1I4A���p�� �'�B<@�& ��90�aĀ���`�'V,(�jU�,��`S���|��'>m04�˗#����� ���'f�Hyu�9{N�2ŧy�< ��'_�9�n��(���խѢ]����'�\�x6�@�^���)J��ы�'��=��б.�S�#ܩ1c~���'t���GO�2b.lc �4*����	�'�"��,ev���薍Sx��:�'�>�$gu����GᎿ ��J
�'\yz��4�D�k�N�C)x�r	�'��$2P�	=������f`���'�aHg�
U�����o$�j�'/@��gJ8��(��
�"�V��'Yt�8ԡ4_"� �R7��4	
�'xL�#GH�;,���g��$u�X�
�'h��`�@1-zFe��!� _�<T�RS��]�Į�<�d��J�<a�'V4m�+�i;R,���G�<�7�7t�Ve!K�:��(��'D�<���/{@��	�%bpp�ӣ�|�<������6I�;>��P��
|�<Y�L�*Q��9Yq���^����h_�<Aw�w�V���߻T�.١� b�<)��
�,�5�ϴ�=��]�<�uG�d<\"eM2;x
D�WY�<	��I�?�u�t�1�x5(�R�<��)P':e�Ó��&�#�Y�<�0�rM��K ����!cs!l�<�W�.]�c��?
fl�4`�k�<��$�	uo�ͻ�I�]��i(2��j�<�s�l���r�e��Q�r	Г�Pj�<� ���1�%��8B�ΐQ�FXX�"O�Y򐇟�Lm���! 8AhF@��"OF�3�FҔt!�x�h܍ ���"O�qԪ	(�~9�!�K�D�6"O�HQrJ2O�p賂�D� s�ɰ�"O��S��7������$S�HS`"OP��N�1r�t���cVINDy�"O*ݱU�Q�?�h<x�ERAe[�"O�I�c
<$}DyyD%�&���3"O��BFӀQW��;S���0d�V"OJ��䏜5i�FHcGȀ�Ym���"O�P���9E�\��
\!Y0J��1"O�H`�c�9=\�I �H�=���:�"OʔpG�̘
���8�!��P�fD�"O�k���?[�l�da|��'"O�!j7O��&�P@Q0�e��ӆ"OB��V�Bhq@86�u��qZd"O���sł2�����,�
d�fa��"O�񺃆�W|�Ȃ!㚽p�"O��	�c��I5��_;h�>%p�"O�eb��E�6N��S�F��Ȕ�b"Ojx�@T���-�գ̤*ގ1ç"O���qHQ6	���OL3vpH�"Oh�����'ݲQNA |B.��W"O^��5�
7n� ����
!E %�"O�!�͑�:����r.K�d⦈""OF@1���)wF^��"�5|��=#u"O�	� N7Ť �(������"O�e@�(̼i�G[�N �"O,�D�M&�&y�����d��9�C"O�̙�'�'��Q�4*Z`��"O�
�g��k^�S� �	�ၱ"O���f�|��(`�̨/@:��0"O��F"O�=3�h)'�=k�"O����CVDԘC����8�`�aA"O"M�6�I�V��p��c��%�Ϭ�yb-ݚ/���Vi�5�2��Q.��ybKO<�ԡC�ɣ88>�Rm���y��
	[Ѝh6�J*3MlT3�dT��y늗 S��e�Z+y@�i��8�y�J��z�Aw��)۰yA#m���y#*~�U6�Y-N8�x�B��y�I�j�	�IL�>����-K<�y���d `�!��&X�x���ݠ�y����#�����լ��,X���0�y��<+$f��DĶr���Ʈ�yb!�H�TsG�N�,��G���y2aB/Ӗ���JD֘M��,�y��Q/Z�A�B�8�Je��K��yҋ�1 P�}0��}��j%���y�/3��xQ/.!�y�Q&X
�y��Y���A�k�l�P��%�y�A؋-g���D�^�j������y���o��a�#BH*��M�פ�(�yf�!z���U�Q�F�ضaA%�yB/ɥ4s<�k��I(	]f���B���y��	
���G� "U��#�yr�)VjB8�q��sQؽJԪ���y�/��^_�8qn	e����y��-Hit)�"���b����"���y�)
GCP��7菶F&�1;R�/�y2Ǆ,HL���"�=�p��am@"�yR��9��Uv ��u����y�Õ6\�RB�9 m��hЊ�y
� �i�ì�Q��<Aըϣ8�bT��"O��q��������%��y�"Ol��C���숡Mh��U�P"O�=1�c_"�����ձf�^=G"O�d�ԣ�'^n���ޥ_��U��"O�5ˤQ&_���A�y�ؤە"O"�CکT���֛j�F�;6"O�� �"]7KW��kϫ"���A"O�1А�H1O�ᐥ�!�A!Q"O�e�q�T.X���+�=#�x�3"Oֽ#q
����؃J�0(���"O����Ξ8J����!��=��X�"O4 �p�S���c�)6(J$"O�*d�H;�,9F)�`
|;V"O.|�Z)�2�84"�0���"O�ESF��(��ɹ�T!^�XZ�"O�b�d��"�=��MC�%wF�B�"OlXÏ�!bE�0o��;�"O����E.Z����`"�IR"�"F"O��)B�_��j�[� W0o��p�"O�,�%���4��01�֊oW��[T"Ot)��P�2ON��G�؆q"\2�"O�hjP�F wS�; ��8L�\���"OvQ��ϳp�8���_�q�nS�"Oڃ"�Oe��� �G\�$er�"O��˦�
�$��(qD�	�,B��"O��p�&I(Vi��8��МO�*��3"Oz�U	�Q�.���Ώ�P����"O��`��c��}����}����"O~t�w�H#!��T�%{LX�"OH�'�S y�j	���4C@6�k�"OXIy�mQ�pt�P�Feݨ&8��s"Oʼ;��u]�ńV40�Af"O��k�h����!�gQ`��"O� �R	�*#<�Y.8eJZ1�"O�Qm޹eF~��a�kW��`"O&����u�R����L�|"O�� �	%��ܣ�$0�L��U"O�5Od�i���\�-�t�a�"O츱u�v*H| ���/R��p"OT��+Uj�JՀ��6$�F`�@"OP��u��Qi�i�Eܐ����r"O� �� (l81�FN6R� F"OI��M��s:l���g3�[�"OTd+ �ȸM����`��V��PS"O�d�����x�O$s�3�"O���D;J�椒o��gV,��t"O�t��c
k���Q!l�u��"O~L�O�8;�0���-��K/��"O��!e�	09�{����j�J���"O�8�s��?N�`@4a�;w��x�"O�%P#f��^5b��CX�Sz�q��"O��ؑ�P>u�\���;B�R���"O�����O+t��� 6����!"O~,�w�40�tS�GS��n(�U"OR�XdA�	0ZH*� ��:�氬t�<1���S�p���?�t\#RɖY�<�b`�-"U�h�4.�z�$�ufBA�<�S�ǻ8��\[��[���Zĩ��<"R�-�VԊ��Dj�J�S�Mx�<�q�\�(}�Qo�-�N܂�����y<@� A�,�&��7��y"�Z�e�Mf�Ig�Ѕ��,˦�y���&oR�J#���^e��bI�y
� ���h�88�y	3ꊉ\�eS"Oha��W��H]bU����ɀ�"O��z���Po����S�<��u"O�Y&BG�bK�mR �
.}��T"Oz���H؎�(�U�0~�T���ޟ̘F#3-���'���^?��#e���
%��/>H�6�
�b�l����?��Ha| ���A� Ў�+����J���g�d>���mǩno�PC�Ƒ���x���%ғD@�M���P+*n���oE�O|�T����6Y\
�8%M�;gg�8�rF�.�Pa� �g�T㞠�P@�Ob=o��M������T򸀥�,Z,���ϏY�y��A�S��?I�L�M�X�t��w��bCM����	"�M3W�iț�	�08�
��[���`Jg&���~�G_�u�ʑ���'�2W>Ś6��ܟ|�	ʦݙŕ|z�U�d(߈Qr4k�H�Q�=�d�5s���ѳ�ɮd�P��?y�O��4�ƈ�1���	N��2/Ǵl$��9�M%�?n�0��I(VG�pщ�s�)��L����5��J�q�v,��hڀp�x���*��M�'��4��6�'Y?7��xn�pXRc�9n����5R?���O
��$�2U��f掽{�ؠѵ��r8Q�T:�4^d�6�|B�O���>�"T��Y?`�D���D�9����۟�B�,6�T)�I���	ퟀ���H7m�21	��A�-�TUZ�Bͪ|���b�&��p],�8X���m��?�c�IW���F�u/p|��ɔO"�i�ק�n xgÊ5G*�0ig$�~B��!#Vp����<q�$h�D�٤	]�wu�e�7�;w�oԙM��|��8q���I��'m\�s'g��?���O&�����'W$�����A��� bX�y<��qe@Ŧ�Yߴ�䓝��'��DR�/:��c�:M�^|ZՅ�=��i��aU0a0���O>�D�O�����O����O�I� �׿
qX<Ҵ�f��\�%��=����-ɦi�E�A�o�Z������$Z4�y5/M3%��Xe��/R�U��-���d��b�a�Z��R�۾Z�ryCwBۇ��'������M["
��=w��еf�:cʚ��B���%��O��DK��֝�|:"�Kt ��!�R4I��ț7&Kv�<	�$��1�&�ã�ιj��PC4�o?���i��6�<�b����'��_?9��(�	j���r5JX!)��sՠ�������?��_A��)S�D�X�vl;6�֖#GTQ�&fy>e���+BL��D�5��@1�2� ��P�0�Ѻ0���xRe�q�ht	CO�3��C@�2�SU�t<+�$Q6$�����{�h��?Y��i��O��桅�#p�L��f�1+m���� �]��.�)*�}baa r\ ��z�����
�p>��i^B6�l��hȠ�_(:{2d
g�,�����~b���7m�O��$�|J�-D��?���MK�R�#�A:�2d���Ꙉ4଱�Aƕ�1�*�:5���B�h�H�-�V�)|����N�:A��c�YŤ%YE�a�r5Zs���_�<��s��/�t=8�M٥5��ʊ���s�e�5*,��ٚafPhײ�t�~�D���'��6X��Io��MnN-I�� sFMFe���� ��v?��?�����O�c?kG�[	o�N�8E__d	�"�7ʓR��i��'h���FR=9V�M���ڲ)�2A���O>Iۓ,�1�  @�?    �    �  *  l!  �'  )   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic�'��}9�n�<Y'��{*�Q놏 $n��V(�u�<����8#¢][G�ÿr�(�@� �Lܓ^�XFDFQ?!�f���E8"	Q��ۚ3���B��#D����bڥa��a	��+s�����ѫJ��\"�v}R%_��7���t+�.�h�@f!����ƓCI���5�y������w
]+��
�p|�#�J/��{��
��n d
�!�'CX��y' � ���Gh_F�00�Da�H�Xx�3'��Z�A`�Ƣ81!�dK���I�$(7%"5p��"��JEh���+D�mK�+�i�Q>E���b����0&A�������;D��p�KSr@��5iA�f�`ɸV�.7к�3!T�h2��+�lc>c��8�Ԛ>:����C�a[�`��"��:��5w5�ZPJq TD_���0Xw�@3q���a�'����D4�Y0&HÕ>���V�6Yџ�bɈ M��q���eS�]Z��%��� �q��ZU9��&4��1㌐� &T��ʏ8&��	A1�<�T��b��!#�p��9!�k��?���	ڍ�%cIS�  �Ch�O�<���f8�˔A�3�:��u���jЊ�c�+���7MB'3�L~zf�|�I\�,T��&N�1ވ,��l���?�AL�T�l}
$�O�^<5��J�67����Ƈ B����C�(thq��'z�T�A�"|�NE�z���`��@�G���iU����'��^� � ��{g�L�;lh=�#呻g�
��84�b���V�ƘJ�Kɯmμ�#��6?1����[�x�C,���x�Q�"�x�OT2$���B%q��yC��*c���z�'�6�(�nV4a��y����U ��qgbC�ofDrF�i�XȎ?��Ϙ'�	�CE'#$�������H�'�V�F	k�.��E)ߋN(�#��S�?���ҭ��䌂]���#�M�z������t���j-lO�Tp׈^V�SC�Cb� :Ђӝy�Z�	6v���ȓw.di3���S�	����/
��>i�˛�/޸���$�'M�=`(��S�|���ۊ�,��ȓ���`B1� (J@f[Ne8U�Q�O6 A�O��Ȍ�Y��sKٲ<�\("�&�8�hf/#D�$"�iFe,4����xi&�[�{�6̊����&�����E%;��P��()�iC�g��{�ʉd�V�n�$9k��U�T�����6cnh�ȓPlH��@�u����l,��ȓY ��6�ּkےHed�i�p��ȓNX���M�ws�q˄k a	����z��e@Ec�
q�ܘв+��*IX<�ȓ.�(�Z��&>V9(�ˀ�<(�ȓUF�%1�OϜ&�iGeC�P��9�ȓ
8B�FG�8[�	���4e~���E��mcgW�U$�UJ�ɓ�SĶH�ȓ.���*�
����+���:0хȓW٬0F�W;��X4.V�6�T`��Pm*�#�Q�����>\��ͅȓ������<[B�ch�=0-d���s�t�{�n�mɤ�	�hN�Y|����Mx ��U3=�� �e�A�����
8@i�$�C�H5A���\�J9�ȓO�x�����*	�qc\�:��ф�Io2`����΀	��Px�ȓ_
v��l��rXhPѲ� I8vd�ȓ%��=2�Y"=o���ŉ�#!�p=�ȓ����!�"E>)�c�?;�ņ��L�p0';��"`h]�z%���[tȕ�U�W�T¾��@BJ�B݅ȓl{���J$t;tu����	����<����4�^�#%Ra�w�ƈ}A�\��n?���R2#�)�!@gM2U��;��*�"fc@M"�e�B)d��ȓ ���`��U%Nz�ً +6�m�ȓ4��\#'$��݉+Կ^�d%�ȓ�� ���C(d����d����(D��a�EI�J~8�3��|���3�`6D��1F�ŘW�������yT�q�UD/D�,"bB�GD���Z�k�}B$.D���TJ�BI(����Y(Q�̐;�+D�x)�ήeP��t���S{�Xb�M$D�H� dޜG�X�)G�O|D��Qa#D�0�F)5C�(���M	M��rs�"D����ȁ@��(��b�����{��+D��idN��+�ݨ�N48t�bDL*D�T0c珓C�HQ���cj6="�-D�P�Ӊ¸<9ܜJ�̝H0�Y%-+D���+��c�ĉr���K�U�a�;D�X`V��c,��P.��t�u��8D�4{B���>�0T+�����"xAq�&D�(PV�Y�h#��#B^&?�ܫ �%D�P0ր� _���z�a��>��<X��"D�H�+.`��H�%lk�4CpN D�����%||�Qu!ޜK�$��*D�1JQ�pm~:��7'���M5D��rh�6Z���
we۬t+2���>D�� ��{!��_��a!�#�+d�P!�V"Ov8��`.!^@K�G�*+��Բ�"O�y���3�̨2��a�$��3"Ot��D៭V{�I�'-L�T� ��"O�1��G�}����r�l"O�Ck̯	l�1���\Z�E��"O"�r���pj8�@!��!G�كe"O����vg*y+c�<C�$��"O�8 �f��.��UE\1r5$@��p.&��fS`X� j�GX�d��0��<���N��y���w��Ĳ�ʃ=�P];��O��y��A�$-"6d��7�� '�W9�y�gI�h��C��y,(TѦ� �y"�èz��4��� �i+Q
G��y"�8~p����D���?�yreJ7>g|��`�ɉr$���&� �yb��qi(Iz�I	�<9���;�y�ҏon>��)��w���rw��y��Dd��n׽u�� f���y2+�h����qDx��EE��y⭀Gb�Y"Nĺ�0�#5����yB"ɦ:��T�����d|%�$MW��y�AA*4��'�
�斐8ĴЄȓm�M �o�r@�pΔj�!����X�h��>��Ҧ,�J�X����p�C�и�ƭ��H�W+,��n�H���@�Q��U{�Q!���C�����P�#14�:�嗄-,.̅ȓ[�|pˢo�Ƹ��sV&@��C�9e���8v�ί<| ��6HQ�o��B�"M��q���s.	��"�B�	w��Ā�,H d����(O(E��B䉞_��� P2'���Y���B�I\$�CB-T$n���
�I�o�&B�ɯŔ5p0�G�RX�"cC�q��C�I�$��ܰ��*>䠙��`��C��E���p���"h��	�JP�}��C�Ɍ>��m� ����Ȩ��-У{��C䉇2��馬ɨ'ФkՊ�}�C�4T.�Hy�E	2�����3ӒC�I ]e�Q��`Җ* N�C��.-�C��������<Epbt�L�9�C�I�e�@��V���$�ġ��4D�vH�����B(�dB��S��!�.Dߢ�Yb��(Q°=��ߜS�!�B�Ff��*�F�����
3�!�0P�4�XscR�Rj���Ԉ) �!��"E�p#��mep1A��L?�!�D	�1�b�C���F�x��ͻ�!��d_��f��*��)�B�Wm!�DǙG�8���Y�?]�I�d���3>!��8g�� �ŋ:Vd��"�!��&`�zz�%̘H6@��ƅ�d�<�բ��	2�����[�'�`��0�]�<I� ��y#4T�G�R���:��b�<i�m��F��D�b��b��Z��w�<)��t�rU�Է9��QB�*�^�<�3�C�z��	4��=(�|uaԪ�Y�<���Q���8��M/%��
XR�<��
[
vx���w"֬n����M�P�<���1>�T�"S'\�!]�� -�L�<����GYI��BK��f�*�`�F�<YUʎ^a�p``�0eQ2�1�E�<�bZ�vg e�3l�4Y`��HYB�<� ��h�#˼~c��Ġ��)�l��r"O�!g~���" �3n�f�Q�"O�M���ϛ,�-��H,g�H��e"O���� w��-I�ak{��
�"O��)��9:�.ik5'_�AZ�qg"Of49b��X7j���'+P'X�`"O�;D�ޤ��!ADa
>�2���"Oč3�U��D�@"S�C�d4��"O���2b��2�����~@H"O2�`a蓲S���a5G0j�LP�"OD�"���պ�I��˦}:�(""OjT��
�����@�W"�̈�"O�AHba�63���A툢[|M�r"OQ�p#�UY�e�K�J
й*�"O�
�`��mbpiV��6G���1"O�����{'��l�
7X�&"O �ǲ���"���5��x����{�<��LW'E���*G#wE@e��D^�<����S{�D��.Ω4�2<Aq�V�<с�^=i8���,�~� ��GK�<�S*�������_$d���m�<��U�Ot�$9�G�&~MR�Ǚk�<�Ǣ����u�<hsjա��Ep�<��
�	���/Ѱg�)�7�m�<DD�\�3�V�I��� W��h�<A �A��H�& E��� d��h�<��08u|	��bـYo:]�%�AN�<�dNU5g�vD���U�2���$�J�<�4�F�e���0�9O�<|;vi�<�e����*�
� T<X }2�J�F�<��a�=^=D���EF��ph�C�UY�<a�I�s��0�'�R#u��b�E�R�<IP�R>h0��AE�j��P�j�<��/�8h��1�+�U�ĠH�d�<�4��:$�����]}c~!�`�{�<y�
^� �ѺWFr���x�<�n���!�MT*"q�Ar�<I�)��
D� tѨa���o�<�r��x�*pQ�I
��Ih�<Q��WX��9�<A�fձ@El�<�e�V7Cu�����	� �|`y&B�f�<��IӔDA�q`a�*& �'�e�<�� �i-ԑ��E�<����I�|�<��a �^�\{r�����K��N�<�&�Њh��Ay�KH�	m`�&��<!�bV�AWE+���/�H�aMy�<��%�"}T��(�)C�N C��Wy�<����sH�H�-�q~��D)�x�<�� �9G��M9@T�'�s�<1sծz{�$�QA��j��ܘ���E�<���B?�����8�^\3��K�<Q��R#]���w���Z�z�('H�C�<5n_�BAB�[FƼk-�s�N�g�<9f��/]+6�ؠIX�2�izw�k�<���
����{�P;U�:�p@��5�察=��C�JՂ �����Y���q�9 ����p�F�Dވ�ȓ%�lHQ҆� Q>ecVg�9 ��ȓY18e��N����+��L�<�0��ȓk�Ђw͝�0\���$^��hl�ȓb5QcD�]pp�"�F_�>I�Ԅȓ��a��4��]��P8U�@��XQ����\���K�no�!�ȓB������?z���F
�3X�A��S�? ���6���z�X;3 �,����"O�%�+��frv�1 _�� `�"OT0���>夘+`�� �����"OԨ��bޗ6��Qf-Ț*��Б�"O<t�l����ҩd����"Od�S�)^�E�J1��,�

�f��u"O�ڃ���0���!l*cb��T"ON	�/�7 ��I�!�;F��"O*X!��M C����O�;.�P�"O\ub�B��#�<W�QpvXK�"O�I1	�f1*�c���0� �g"O��($iT�o�R�q���#�H�"O�I��PAZ���t���n;� D"Ox���,P��`<(�����T��"O�e(�̎?V���AG�*<�=�"O�}�$�н=:�Tc�+Q
%m�0�"O^���`܋-*f�[�k��Z\	��"O@Q��һAd�1A(�85N`"O���5�Ί-;|��ǒ�4�"�#�"O�)�c��5c�|�D��h���d"O8<�����Ȗ�� �%"	2"OЌ��OG�˾1Ƞo�6l��)$"O(����ϵm�V�B $��h�H��"Odmӥ�?D�FV�ԄG� ���"O.�Bf�20)
�$E��h�"Ol3Ԇտal�I�"_�y� �r'"O�x�ң]�pg��˯&�xt[1"O����ӄ'x�$��EF3>\�U"O:�pr��p��I!��<N��M�`"O8�+K�xo�ɳ����*[&"O�8�pΓ�Z�q*�A݁��h�G"OV��V�ˆOPJ%���B�	!��"O��z�G^�A{�E�'Ƽ{��"O\0��	�F��L`R�R�.g"H�E"O��e�Q)ڔs&d9"bܭ��"Odd���LBW|����-f^
�Ac"Ot]����,��	��V�[C.���"OB�c���x��3����"O��V�!E������~����"OF]��E]�kJ�J�%Z���\� "O��
�f�nĜar���5fD[R"O��Y��� �̡@f�H�ZF���"O^�x��Զ��12�jƟ0;*4T"O|X[ �p|��!ꅺh:i '"O�	��i��#��hy
����s"OXS�,�1[Q�zgh�%��A�"OvY��IhT�U����u�"P��"O>���Q&RQ�
��
h�.Xٗ"Oj�"�Xn�2���;6|ap#"OJ��U-�9r�"��`�݄A7��F"O.dQ�K.Y[���@,ʪH��0"O�P'��&�Jg+E1)g
�В"Oq �7~j.�+R�_�vN��C"O�,I��)#9������`e,�xA"Oa��-X3�ȕ:�iM�iJpDc�"O��⒋Vh��Y���u�6{�"O�]SsH�eD�Y���ʹL�d�E"OF���G]�1�*,�eF��_> m�@"O� (b*�#<.Er�'1���g"O���F&l�W�Q�Qj�\	"O`��F�Ow!��`%0]�%"O���V�l ɂsC]�r(J��"O	*��Ԑ�hԍH� �xU"O$�1��2�n@�Ӡ߂	� ��"O� h���Ӏ1~�ڧj	%,��H�"O�d���V,*���B�A+D���"O<@S��H4W[�&0�q`�"O��ДI���꟝1���H�"Oj�s��(,��J�,V"]"O:xV$� �gI[�)� ���"O�ܹ�h�	`v��c�ԻCB�q��"O��S�B�pl�\�6��9��"O�]Z%�n)>Q*��Z���"O��A�H�Y(�#ō����˥"O���5	ޚ&�P6K�<�t�Җ"O�����V~.�X�q$G _�t��"Oҙ@��FR�|��]�%��ܳ�"O����	�  �P   >
  �  y  !  �(  g1  �7  �=  JD  �J  NR  �X  _  Ge  �k  �q  x  T~  b�   `� u�	����Zv)C�'ll\�0�Ez+�D:�DlӨl��>O$���'h4�l�^����Ο�0����S{Ȭe�2l�#K+����!cݑ�6E��?�:����?呀dYL�D��D ]���K�d�W�jEɂǓjU)ՠ(4�HDh�u��l)Q�'�?����V�rt	�[�9���股"�n�# �6R��$PC>���%	�}��6��m����O����O�����Xd�� ��B*)uz}�@AV9M�~��O�Di�(�O���?)�e�?����?auI�z�P��H�8r�GD
�?���p��v�'�"�'���N���'>�$�A�xs�+h�,a`P�K��4OV%+GjڶoՐ�+�*�& ��\�dDxR�O~�P(C���ҷ�y�+[��z�ϸ ���'�r�'PR�'+��'�����SS��;y&�H�g�XU�,��o��<i۴g]�Nr�VTl��q�4`_�li�i%>����'�n��2��טas��I�W�6�0�Q�DA�{bW?��$�ծ?3ĘrG��c��8����"I�<8�#C�se�r�k]��H�4cL�f�O��4�@�D�t�%ޮ8�}�ˑ�Q�2��vg��<<�7�`0̓'j�-Z��@���7X���ݩ~�F�n��M㑽i,�#�Ή�yM�鷭�S~m�U.F���Q�'��~�(6m�����4z+��S��
�}�Z����b���`��M������>�lC񫕈-'�QٵhM�;~���i�z7mɦSc�ةO�ބ{@D�D|���>�R�O�!k��T�d],rdP�ش ��M�'�S�p���K�N*CU>x2���'R��%��a�r!S�]l�u���'��O����O���#����O�t�7�D�4��8��V^:�������D�Oz��n>�hB��%5FV!�E���] �$�
+%�U�f�N��4.�n5�"O�ł0l־R#�E9t��f���Z�����OM�N��\��p]��'�ZP���?!�W����@�(t��1��f4�c�O,�d�Ob�b>M�^�~���3{�}��f��N��?a��4���n�7��k��?l4JTCjLCJ�K۴��',�s������5�T-����O�<p��j@�=D����R� �(L����QЁ��c;D�Bs�J�Xkv]sD.TH�!�u�;D��#��;*H}ؔ��3$��m!�7D��V �5O��8�7�� ��%�7�3D���Ԍ�7Vx�� �,���O���r�)�'V�Б4\>V����tM�5x�'{2��%�ː�r�8���:pn�)1�'ሤ�`���ܬ ��f<�ٛ�'~Ɓf��pA|A��\!3�|5��'c���e��F@���31�r�	�'5X,�8o�<Y��[�-2)OB���'�1c!U~�  ��O��C�'MLP�Y#^� ppc�R ����'&P�@CX�I�F�:��*�B}��'�
I0q�HD���Z�'����'Z.� ���F� 2u��(?��ϓUYp�{��i7��:�V�X�͊�G_���ׇ²}<��D�<����?��Ot�Ɋ����M�@�$)���2��pH�M4����D ͯ3�ax�`�n9(T�ý6��)�TN�}���6�*)�Ƌ\
s�0qa������	��Mk�x�9Ks�]��.���
�/`��,A(Op��2�)�'x��c�Ä�_��I��!���?����h�(l�`,�2�mz^�%Y"�Ԇ5kr�K�4��k���`�S��'����8l��y�Į'H��cr��(1�!��Y:i��R��y�
T��@ w�!�ē�\2y�F���x��ī^�!�D
솰��5�2Q��̎�,r!�dD5 �t`嬀�|���V�Oh!��A�=) \�G#i�`TP6�%�۵~����O��$�O�˓�z��I�:���B�ţZ�����Y4�$���,ؖ�֏���i'_M �+Ԧ�_��$e�˵&Z�T����R�Y��C�a��|S�a�Ļq�b���'���BաR��Z���*ܡ�^pɡ�蓮{,OmHE�'1���'8b���X|�nH#A��-��ă�H��y��(���͘��X
F�>��*�8����O~�l<�M�I>�'�R(O81�
n���+��N|
���\�Y��O��O��Hݺk���?��OQ�0�cA�2�ak� {�.M��'���xϓslL{c�Z9Y�Z\����)��d
�'dLKS	ެ#��L�8WnB����@�?��'#�h[�lT9.�T���$��'	���a��u?8ä�$��J>9S�i7�'�� f�t�x�����ī�W5<u�E��Ih���Zy�'O�'{�!��Y�x6*1	��_�F�� 6)�FO��Ʀ�hr��w'����'��Uk��@)2���y���?Ҟ��g�ǃ.�8Y0�#�0<��l��[�4�?���=��T���!es���£ڶu��4����?���?I���䧡�'�FY�P��#f2�Q��F�?�l0��)�a�^U��E�?lp�p���?A-O`������IßL�O�����'09�IĚ|���⥊>r�(5	��'�R!��:��T>�'��(�f��B��dp�d[�t�ܥ�Ob]���)�' �a���b,�!Rn��,
�'�Pr��>+ɧ��Mۃ��:NVl<XCfM�jw �0r"Oj�VK.t�������]Z�ٴ�	K}��9ғZZX�:��d ��XD�	����im��'�rE1��l#��'���'Gb5����#\5K32�k��=,���A��d
&�azb	
mn�����K'�4 %c�/Ә'���W��(r5��.B��SFT(1����M>�F����|�<�qA�(�$y���
��81]Z�<qb'		� x�H���i�CƬ���t�����|��:o,�`�K<^�䄱V ��>�H��X46�B�')�'g*����$�	ҟV֞ �B�uZ٢$KW�46@�RD�r���G�s��ݘU
�#>T�E��LQ<OG��VnUm�ȝ�0c� ����ĕm�h�8�(U�pH��(z\R��'$T7�En��?�����M�dو�(W�|�*-X���*t�R�|R�'��O�1O�c׏߼:�2i�wIg�h�]�x�	��M3��򄎴*�F�nZٟ��ɬ}m��W)D�δQ��H�2���I�����L؟�I���B�H4lxL`x�O��*v#����w3���B�j��/#O`q�I�� "4� ���7Lq�an�K�j�Pr�D�X{l`'`T�i����ǒkT��'C�7m�O~����]G�Z����8=>��VȨ<���������
�o$ ��B*
J�ƴ	SH�..�	�����k�S�-�Or�r��Q�G:��X�h�1ʬ͑�'d�ɶ.�,��4�?���?I�'9OIc�
����-�qo^�#��'��x���?����*h���|*����h���Ƅ ��5���3<�$D�'e��� Pɧ��Y:�Z�{����l�%�x��'��0�(�OF���O���6�'	�8c�GF�\H『S�B��%���D��b�eL�XH�i���JHT6.8�����X�'c���GLڢhˢ���ɀ�3� %��ljӌ���O��D��=�,�D�O��d�O���y�y��T�p�C$�'l�L�ɣ9,����7�3�-"`�`aV��A)D�'��J�4TDnc>c����D�������Z.�iJ���O���O����Oc>��?!�M��l�#g�	W`2��N�y��� 	6����g
=O�(!��~o�	��HO���Oʓ\�ԕ��oB�O(f����U,
�rH��\9���'�B�'��Ig�8]��x�f�=Fm�`4��
��Ā�SGL�8J�g+~���_5T�^��!���v�EH� <��zd聊-6>�Cd�':6)"&b�wr�a�Z�Ԥ"�#ͳ�?��6>�v�'�I؟��?ɓj�",�R��=����k҉�?����O���&扶ik��. |��� �n(˓�?i�T���'�ѐ�`i����r�L�LR�F=@���w������O��?����?�$䊙bi�0#�ԿY�RX��',���"��G��ס8 ���Ó>�ƥ��d]�
�a
��	b��#��*.&<�s
]�u�h�����0<a!�	ğ<�޴�?���(�\-�cb��ð�����. �~0C��?��?����'b��F��;�,�`�+���8��i>����Y)�Ұztʤc'O�����	qy���I*L6m.�	}>�lߟ\1tb��W�h�+��A81g�a������$=�:p�X�d��S����fM�&<�.�ZA`���?x  `�'�\T#7�1F���a-]���#}"�$?�t@��	\���VdO~b���?i�iF�6��O #|
QdM-h׌LKS�G�De6\��ZA�Iɟ���@����eҦn86�U�2?.%cΘ��hO��D�˦I�ڴ��a�֑`u��RS��@O�j@���)�6�Ў��(OD݋�F�,�<�	��Eq�P%��"O|�f���|N$h�*x�ڭ�"O����JV�G\la��@�<&q�Qc"OV9�%8&����@@�ZTX-8�"O��X�?�>�ق��  l�� �"O^mjL5)�e�$��!jQ((��P�X�a�-�OF�)���b3L�IQ�/7Z�p��"O� h��U@�Q>� ��� h�H�3"O�0+��K(-��Х��8��i��"O��P�gF/nO�Qf�)l�JT	�"O���*�X�L�;Rf@�@����'�>,��'3D��瑐<��HӃ.��#Ur}��'�́sfP�i�f��Н!����'��]��k�`�ฉ��+q���x�'��"�ǣ7P���EꒈW�:���'�.\+��3A*u{ Ȝ�w�`��',���`j�a�ج��˅* �ؕ�����4TQ?i�'%M�B��P�Tj��J�Gf���y�i��dn���Ӭ���D�S��	�yd�X���`%G-�by��#G&�y��¸8ƨ�i�ݥ�l1A��2�y�L�	o�9���عL�H飕���y��k�J��%L�@d0����?A!G�N�������2�$@��l�e�n�j�3�m,D�H��A�snL�3�o�F��d*D�z��Y�/�XZV�P�&vt���'D�0x��N*,�IenI�
�$�
�!D��x���&k-��w��Q`<�!sA+D��:@R�!#�Ɨ��M���<qc�w8�$��� &(��ao�1��n=D���1>n	��mS�k�`YxpH'D�lk�O�v��wM�Xޜ�1�'D�HH�%9=R�Y�&�3E#^C�!9D�����cR��#`F���B�f6�O��2��O2��	[2���c�[��U@�"OH$�s ωJ��y� �ŕ{�|�r�"O|�����-�0+�V6e�R�e"OZ����X�]�b��a�!~b4 ��'����",!�X�A�띙*h��)�'�`��nA�b+\<�v��D��e�'h�<k���@44��q��I�����փY�!���|�z��2bI��<	`�Iȥl�!�D�Wc,��tK)ߊ :rɖ$
�!�D��zl�"�J�f�Y3HQd!�䅡L�e�tʑ+-��!Y� �i!�d�#J|���!�Z�OC(J��v�2����O?�F*�P�Xq�Ȍ<G,�CӏA@�<aĦ��]���G���,�+��}�<����I~���	.�Ȃ@�x�<���ܼ|W����� ���k4�q�<�3MK�& J�3ƂH<���S���n�<饁�.5������g��k�g�hy���p>1�`ڌ8���a#��q��!�Rf�<�F��sn�J�7'%����i�<����CQT�Ǉ�2�2��	e�<�r�D<\?����$#鐽h��X^�<�1��c�9v���	�8�kS�Wx�<��%���b��kְ ��@5(���W#%D��x�
�t�p�hg���Йy4O6D�< �k]�H�� �DhݒM}���'3D�4{�-F�jq��ɱ(��4<���1D��
u�)3�&Q���c�R�H� *D� �s�]7Ȭ��+�'yc��贋=ړ	�aD�D��7'�(��#�V#�4�c�����y"KV��r��PE�e��a�Q� ��y�Iӈn�1p��T�N�^ܺ�)Ϯ�yBĖ�P��(�w�uJ0��qѪ�y�BL�3�ЙA�i�}XQj��y2��\�����6Y�����,�'�?1R'E����r�#q� :\��0#�%c<�-D���ĭI��A��#Z*� �8D�� T�� @�-�`X� dB�)8��"O�����ӻ1�p�c㋔V���"Oڸ�P��� �ĸ14�=b�L�F"Od�:�o �([qD�^�l���P���W�:�O���EA��zCҕb�L��c�^��s"OL�� 
I#B� �2� 5d0�ˑ"O������0N, P���`ﺀ�&"O�;Qe	[�x�$�/�f�c0"O��Q1 �O��H����(���Hc�'Ym��'�@�R#ѩ/�������蝲�'}.���@ڛf�	D�J���k
�'w�);B� `�>�Ҥ`�<5�M��'Y�Ѓe�[�~y�G獮%چTS�'�
H	q�L�!ئ.�'uˎ���'U��S���I�t,HUΌ<mG^*��D�*Q?S�E�{cF����R�dx�c-D���*L��T�F�C�l�[�,D�L@�
�p,�A2��@�`�{t`*D�@���$p<m 1�gZ4(�(D���"d�hb̄�w���k8�ZaK(D��S�#_"E���&�H�[�
�p��OةS�)�|���JʃT��B"�+3d�1	�'V�I`.��8I'���Ѓ�'	��z ���i(Wm���
�'��e��SED�������2��
�'��p��˕7+�`aā�b�,I�'�r�����8�HꆄJ�0���,O���'��=2 ���pa���P�Q��8�'�t�S��\�3n�Y ҨL�Zcj��'����C(�V)�r�l�Dʬi
�' ��E��0`���P@�'>2��a	�'_Zi����N��ȗFȵl%�ݢ��\ ��v#��zUϮ>�6L���zs<i�ȓ�*�c�B(�8�/Ӷ;��i��f�nH��-���>%�SI�-#���ȓ3��9��cSp���UE�14Z��ȓ0�\Y�iX�z�5���҈����&��ө�	e���K�C�LuV�G{a�����(D*�rt��"�V�7�B���"Oެ���.D�H ���,���ҵ"O�U#1	�A�ly��[[�@43�"ON�:�/�sɤ�� n�;d�8��B"OH8�U�(Pb�)A��X�0fl�"OZ����ܵ�c7哟(-�� s�'2� ���;o�d:u�S)r��(�Q��	LH���_쎼�땇P����/d�D�ȓ��5;�	H�b.�!�� RS����Q_|D�S�QJ�p�b0#N�)����{��� k��1�B6|�F�ȓm�,1�b���-0�%�',T�+X@=�'�H=�	�@S�`Xp`پ�pH�@m�' ���
�	�ʋ|	S�}����ȓUI����ρ2wfZ��!C�4��\��S�`�!V^�ZJ΍:�d�P]�ȅ�9�����۵}T<�H�&Ͻ.�����	QaV�I4 �~q���/O40b�B�%,E�B�ɭ|�f��uiV4V���"EūU�B�I� �p��E��;$����>	\LC�	<^�Tx�F	Aj ��+�E�C�	�O�faa_�d��=Yc
��sY�B�%O!>����ߓcV(����K���=i�&�w�O��H�g���;���ˇE��T���'�,�K�"�6'�p�!�ӱy,P�'�]cbM�!V�|y�Ώ j�<���� :t+ �n��Z��V<i�ݳ�"O�[m\�}RHx˰"ۋS�	�"Oz�:f̩7Z$	j�!\/�Uq��'�>a����	ePP$�ōJ r�����oNX�ȓ�z�`6,CE]$\p���j��хȓm>z5��J�4g�`��Y�"ͅ�H,�${U�İ0���[F��<'J���2�8�X�g�xx�� �9�jX�ȓZ�X�;C�J�(T˖�]�'����R����R8(�����/F6^u�хȓrEP;�!�6!��`�A���<N��ȓ:���:��G��:�,'[~���6�1����N ���#&j5 ���P5l�Е`З2cB��Q��;�х��8Dx��=���D��|x��􌂔0��B�	�2æȱb��ZUړ��z>�B�ɸ���P�M�	B$Ԩ�� �BC�I�\/U���߯x|X ��E�!)zC䉹p+D9�����n@걳`Ƀ�L&(B�	�+�r� o��Z,�	��/r��=�	UP�OD~����J?�(��ϹF�dt
�'z��3�	.R��C���1	���
�'�έ*wc�L������x4�
�'�ʽ#W�IB��`,E�l�]	�'�p-R��T�T<�2��=��UJ�'+F���D�"1P���%����#��*�Ex���gK6Me�ʲ^��P��>�C�I��]�"Iȅ?R�Ps@/Q2+��B�I�\Yd�Y�ǂ����L�kӘC�IFŞ��#�&�2|Уe�'cs�C�p/R{D�lh�f��y7tC�ɫ �����њq<@ApT���6�*h�	�Y@�I#GH]�z�]93$�����C�������>u\1 �LW)p:�h���D�	�f1t���ȟ0�I���E�1C!�a�#N�O���P����9`e��AĕC9��@�\�΄���K�:���O�)��#z�n���L��������#E�b�'�1����@�.{�Ȱ[�a�&@`4���Q���	F��ӱI�(9�l{6�	�j��!�O`�'ϰi;ԭrJ̹ᅓ�mG �4\��4�Oן���/L�h�O�N�f�O�rN��%��E���eF���c	��O��k���X�↨/YT��3��O��Q̧4̄��¤�wJ	)0f����Γ#Ҹ	4�P�1C�#҈T4�蟸���HP�n��D��"�t�Ay�8O
y���'b��������D���Y�#±~���ȓz���х Y�b�@��-%�Z�D{�M!�8905�֫ʤkh���o�!���*`��?��"�Ր�+C,�����?��%��n�O���a'�? ��EI�fMuA^與�݀$ hE
�	�!�h�� f�O���oB6I��Q�	ٝ�b�[������2K�?�NeX��ڳT�S-��'�]+4�(�1�G�0a�,�K�O�;2�'�2�I�<1Yk�k؃9Ӓ=(S�(fC�ɒ'�l[6*O�%���H�"/@B�$	O�����'1O��q'��Z��U��
@J�q��'�����ĵz`��$PK���
�=g�]�ȓ?�$iD`��*-6 �+�<a*L��v&,��M��d��(�"!���ȓ=�J��5aƚD���#ݤ&PXŅ�Q�ac�
F�-Ra�ZB��+6|ON�ꢚ>�q��SETE��a����5���_�<a��z�KN3�s SY�B�	*����A�3��O�U�TK
�'hd�9d��%C8�K�/Q���	�'���j����,��Ĉ��]��,2	�'��aWm���H��� '#J�Ј���O�'hB�QA��&x�@bȗ��`��ȓw��3օ�4����HK�q"�y�ȓ7^��ѡ��4�VձF�T=|��S�? 2܃�!ҪD�j�&��-h�PP�q"O)��?7xD��B�E�,�qE"O���5�,_88�H�jʹo�N�:�E%�OB�}�TB���%�J;���"D��O(j���L���B�Ǩ������`�dU��B!�x�"��{M0E��bŀ�С��e�N�r�o
.f���!�@G ^0�@�ȓ�T�a�ٻ3��QY��D?>���fp���(؛!V*]�VL�=%�u��7t|��DF���31"@2pĄ�"b��9=!�$�:746dț�h����j��C䉍�&��TC�-�9��OŖM'JB�m��e{ˀ�<����@�X'T�PB�	�4����b�$E>ݒ��R4]�?YW�D����'�R4��dC �����$*͖P�̓��'�j���'�B�'�t�J�/K10���?y�O��@�#i�N.��@����h!`���R�2�	Q�/�/���`fp�t�K�s	mzW�;\d�G����O�}�v�'yb�g���$|>M�Wǟ�O¹K��� C��.���O����z�']�|'C�96	 �y��?j�b��?i������i�_}2���r��q�J'�~$���V3j��'���'��ɟ4�IZ~����8Eq/�lG���R�L��0<y��X�z���H܎$�
���c�9/�Ov6�1�I���'d�(���I�D�����R��A�iyB@èX��d�w�B�'���';���t�m�L�]�V�z7�ڽt��-:b}���d�*[ �|����?7������5��^O�H�P�4KH�{v@���M�IҟL�����<�YwlB�'���'�$��a��0ē#�ҡ`�o�\F�'|-]���<O�8�۟�^w!�z�*$�c�/�x�6��BkЈ�I38�>���O�t�O��'(��OjB!�s���0,Z�qx��8�z� ���<R�'��y�@�'��w؟�^w6��=.��@Q�lX�ٲ�5H��7M`���M�O���_�~�Sٟ����?(W뙰*�I TnǭrH4Hȑ�G� �BϓD�t ��˟�
Xw�21O��0���46m�A�Hҥ��-!z�P�6���mj���O�扵oR�D�O�X�՟?���ɟ|�t�$<�x�"�k��A&nG�M��۵�yM�>�?���2���y¬������9����P�\����ps�6*H���Q2x�P����ܟb>�l��A�v��K��lz,n�� �ȓ��xf-D�"�����F�NalZڟ���y��'��'�^>�حR��)�J�U��d`�t�h6-�O>�D�O��$�Ot���OX���Ot�D@0%p�0*��p�H��v�LM���lRy��'��T�ByB�Q;O�bгA�F�V[&��3��g��)���2t,��l}��7F�0Fh (��d�>��|��q;�&]k�2u��Aa)xQ�ȓ4i:b@�]Ύ�uJS�H��C�s���`���U�V��0��|��C���؁{af�p���!0)ʣI�<B�I|r�; K�%O0{&���B�	�N���# R<|y��TI�C�I'4@���7Z��Ҵe�%SD.B��^ Fy%��(V��h�,),�B�	�&^R4:1mR�9t�q�� �8B�	�LL��!�B�dR��6J��;�b�t �� 8�<��*��ӌE�!�ح�|`cH"����j
�VJQ.ה?�$mQs	͘;��@��$5�Z��0���8|X0l�">����)؊������"^��!e��K�r�a4�?dA�`�*F��X���L�@*��y|�y��y�9(�y&S�m�0e� N�&r������"�y��ɏG�lY�D�BJ�r�nӜ�y���Px�a�(I� �S��Z��yBaW* ��R����A�H< �@�y���J�FP���D���c�n�?�y�䔴 |�jR�Ƨh:(M+��;�y���50�*��u�̳^즱k�I��y�.V��<��MG�X%��Ȓ,X�y��֖n[�-�ql��d%��A��6�yB��"	v���`��&�Tea�݇�y��6B��0���Bu��,�y� �F]�5+p��p�����yc�L��p�-M�44�J�#�y
� pHUcHY=L`��̆A����r"O�xЄ:��#3�	+e$U�t"O��q���,k����-F�9�V"O8Y��7<Z�z�g >����"O)���գT9��!��%n���"OX飑`û8�>�Q�l�u~HP��"O2[�d�@� �G� 8L,�Hg"O���F#�"{ ��n��k��lI�"O �h3F�vU��T�L�
7r	��"OP�0�X#+x،�.�$y3S"O^�H��T��i����-R��0"O��*b�ɹjz`=� ��X�PS�"O~(�d�_�_m�L�?Z����"OjQ��@U�����" )("O�z�hI�C0���n�^"�0�"O\�3�O!WCB5y%�w*� �"O^�A4CI+�4m�ʌ�{� ��"On�v�Z;B>PZ�&�7@|J�؀"O.��RC3D�<�/a�0�"O�"�n��[��HG�iV��"Od�����C�ޤ�gl �w�j�0"O隐$��f�P�*vjΟBIZ�[�"O�e+�)�5Ԇ�bs,�V<z\QB"OD�a�[� `��e�_�[� y�"O��`d��Q�0\�f�0y�"Ob�����c����7��zq�uiE"Ot���!�2�M�� �Mf���"O�����KOL����� �#S$��"O�	1��ҽy����O �����"O�bB�)ߎ=Ɇ�,U{�SB"O̅CEF#�:E�u�8bt@#"Of�
��L�A��I���W�\Xq��"OV` ��H�bZB��BR�KZu�"Oހ�偐�l��U��&��(9R��"O��`tBW�|͚D�$&��2d��5"O�iṙ�|i�x��EJ�9�� :�"O���N� ��}AE�w�@�+"O@|���.4x�&��{z 1s3"O4���gv9��)��lC3"OTй2�ͽdT^`:2_-	#D�7"O���bD.0|+��Fp�L�"O����cY$\a
y�ҋ�RX�Xy"Od�l�4�6�[�-�4f�-�6"Ob1� @ۣ8�*��'쏝>K:!�p"Ojغ�n��3��a!Q+N�qj*��a"O*x7.�6;�m����YZ�F"O�h$�Ӌ}� �@ǉ�NM܀0A"On��$��Y� ��ufD%8��a"Ov����ܜ^�^T���ĄDȜ�E"Oȕ"׈ �����Dk��Pw"O�i���%n����T¾p��"O��u��%J4�(*#�"`�BH�s"O\`��+��R��ɩc�<9 �"O��S��
�89 =��Ӈ&�tEҕ"O�,��B�Z���䞷E���B"O�x
�"�!���7��-4����"O�t7���L	2��3V-��"O&�Y��F�)n�E+aP�#�XA��"O�A�hp��3nC%(�0q��"O:E��CK���o��]K�"O�t��+[�R=I� �	��;2"O^�C���X>�4c%��_�VLb�"O����)�"F�%Q&
�V���z�"O@@F��:��qiZ����!"O� � q�aʨr�q�v�Q
��]��"Od���o_z ��j�O�����A�"O��	R��)�&@���G xxe�w"Ou���+�R�f����4�6"O.�B$7h$ 0��A,�z!˒"O:��**���#L�7<�,�!"O��rP��,6*�I&�Q����"O�X3�+܌/؎�����=J�peH�"O��0�Θ3"���u��+Q)�q"OR<p1��N��p�Q��3���)"O�܊����T�0���g���p�"O�����V�<�q���� ~�� "O��䀅�^��`'�^�z�bp"O��E�.wo4�p"K�jZ�1�7"O�Ly2ʙ�!pz�3i�98�1�""O�]���CdO �2��,2-~�ʂ"O�����O)W�V����Ԉ.����"O��r�* 4�޽X�#ε-zܨXu"Oj�� ,2bH8���#oq(�F"OP�k�#�Q��(�S�4)����"O@qA���\	|�K��(y���3"O�hb��E�(`�q**r^��e"O�jb�R=�D%XD
�
'gހ
�"O$�����Q!r�q�k��i3l��"O�q�`�Պ.Z:i2#J�3-rp�!"O�hb��|�ZykP�:��"O)XS�)l�XL�S	_�:��l�f"O��6�Ēc�F<C�:�xeH��y2/^*8J  ���MR�Rԡ5�y�"6���=r>Ԭ� �D��y"+�,@�mtA��j~��H��yB��4L�hT��5[�����U4�y�J%�&u����S���q�\8�y2* 2��=@�ɿ8
B(���yb �%y�T��O�aOX�۵�	��y�;�D�$ǅ�YIV�Q$허�y��T�nZ�-@4�7Y��S@���yr�̓8�)��O'�qR���
�y�C���N 11�Go� ����y���?�6С#V.?��)����yҫ�)gG��a�I� ��:�����y����:�0��ՆuG`�!��yb�`��e!�Z8PF!�����yB��b|@�r�D;0��S����yB�OALvMK��^{t����d�/�y�D��9@Z�[D��e�����X�y��:0�媍e`P#����y���*r2�+ժ�c�Z0�M�yB���x��E�Ҙ_Sj��l��yR�ȋ�bI!�`V�NƮp�V.���y(N�/���-I�MUQ&���y�㋵gH`���j �!KZ��� �!�y�Ǖ�B9@d��#ջ �2� �O-�yR#�e~YqLӛ������y��R-;��x��P���X�����y�k�:�XE;!�O�5���܏�y���&=��1��M<!��կ�yb�L�e�����`���@{�`��yR/Z<<�Xԛ�X&r�L@'oK��y��V�#4 ̹gnM�Wf���gŻ�y���v��U���JT��SW�G�y�Ad����d�Y�<B�\P'����y�!�I�u� ��	3��%�F���yb��m�� P�0|q ���+�y
� ��C���-��`�:@�U �"O���u�ېXc�t�4���n1Fi��"OZ�:1�#p ���m��|)|]�q"O���PCT/0�h�b�#�!����"O��aw����n|Z�A	9רe�!"O�x#�U�,V�-zB+�h� 1Q�"O�Q���E N�����Y�����"O���t�#r�ɒ�i��X��D��"Oh��m�aQ���gS� �1(�"OP�)�-P��ɂF�=c���"Oj�c��/�v	u�X�Ko�T��"OL0��(5.q���S�|�&�T"O,UJ��X�+�`�y���	L�EI�"O�r�!��5d���ʸ��Р'"O.���'a
˄e��w�0���"OZ����JE��	ȫ:��G�>D�P��ͣd#@L�e%I��J`�"D��S��G^@��!(F�[��}��F"D�;Ǌ�-}@���$[�)�B�:D��
��

Kd���oB�=@��2	:D�|ifj�*g3^}x��_Y�pق�;D���b��:�QR._%X���� O+D��Q"o��8���D끃tքq4e&D� �֊�z.d�K3�5\��b7D���F#�u��	��P�̘Qq!*D���E�`����82y��B��&D�X��UT��H4�^>�8!��%D�hӰLB�c��Yj����ktLY��%D�w�9���27�G"c@�Rw�"D�Pp%��V�p�x����z\(��%D�k��g�ι��� �t�h��7� D�� 4���L�*� ��ܕi���>D��Ӆ�^L\u(�	�Y�bD��.D�`7�ֳOa���6���9h".D��y�Ƈ�G�
Ղ!�[�!��H-D��R�<@\9�GaZ!��,D���0`ό����')��q
��),D�иSIY�1��z�WY��g%D�4#Ƥ��*�z�D�.w���P� "D�T�嚯)&�9���Q�8��i�t� D��i�$IQ�l����$
���iv :D��ibo͌@S�y!�&T�^�Xe�9D��B���`�j��6��:�~�sV�*D�\��%^#<��$(0��p�B`o3D��ٴJA�m�:�6�λ1����/D���J#�M��Ig����.D���I�rz�PL�sb:A��+D��S�o� T�����;x.A�3i4D��;��I���Sm��&a9��1D��ZF�Մ�f� l[H�d4D�\y�˃�tK�U��Kص�*dB�-D�İ��G�~H��'b�T�6(D��� ��cܖP�&��a+D�Q�0D�x8v`ӹz$,�!�]�g�Zq�<D�@xwM�E�Rqx��)�DI2Dn(D�D��� b��C�L|�j��v�$D����By�*`�J$ygLD�ӄ7f"�h����'���!�]3��O��aGV
�1���;V���d"O�'.΢/ef�h�F	��ybD"O 4�t�Hnd�f(��\�A"O�pzC܉G4@�J�E`(2��""O����h���#שK�\�r0"O��
��m�Q	�%1pX�"OXAa���r-�`��ܾEZ�@"O� Di��@�S� �í�.e(`��1"O���5�A��h1;wFTyF����"O�m(E�K!V�Ę��dI�E�f� "O�٢P�%p�I9������"O ��2��`i�N�H���"O�P�����a�VhC�?�f��"O�HiQ�>10�뷠�#��QA�"O�-�Uas���C��(.��4�g"O: :
�s��,#�B7-����g"O�,��-˾L�L��0C�����"O���a���QRU)���&b�2Xt"Ol��s �7/����ˁ�R4��"O̼iB�<�Ѕ�К`�2iXU"O8���.
��1Äe��)Y�"O�!�g��:] 2' 6���R"Oly�Q���'rT F^!Q:�""O����ݰD�z�I�OԶ3� [�"OJT`�)�=2�h�C�A*���#3"O��IG!B��|�W�KP�j5
"O|��R/?K�LK���g �1"OZ�r���5�tI��Z�T�N�B�"O�4�EB�=���ق���A�b�
W"O|�3am�5ln��bD�%�"Oz����F�,��ЦE�]�b�C"O��b>v�Q�T�0JW�"O���s�=�8�!/�'^M��c"OpY�B�B�l��ˀ(zGlu�""OA�k�.�pU��Jب���"O,5�#�@�#����4iʻ�J�Qb"O  9�#��J-�HZ0Q���r@"OЬ�RF�[��9�D ��� ""O\��E6#v8��n�r��5�"O(���*Y��.(�D�s6"O"�(��9�(m�eM��D��(��"O�<v昼U��K0�5k��)�"O2��vɐ�ɌՋ��ę~x`�9%"O�����D�bh5I��>�l+q"O3��L� �H�8��5�"O�X1@�c%�p�MH�$��#"Ov�c���&|�����5<��\t"O*��3C��>����Vb��-*�Mz�"O�e��ٟ,��(V���$��B"O���U�ێ+K����;�ej�"O2XР���:ԉ������Ps"O-Z��C�F������/�V�Y�"O�%��L�I�ˣ��Ze#�"O�K���>�ja��Z�*�,�(�"O�X���W�-��
4)�`���"O���⎆�{[T��I3	R��""O XS�d���l��Q
IArQ��"OR%�'�؂8�<�35"�1FA��A"O���2��ddH�C�X�~�@�j"O m �ϚxP�X���VƜ��B"O����H�-^Ei�C�4���Q"O�@Q�a�ҽ��c=hw �f"O��*U�&�"�s��,Q��#�"O4y"0&�!��� �+`�4�i6"Oڸ3�W)9�`J���cΦ�2"O� pmP�	B�ih�i��4��(�"O�$pt�X�b*�D P�{�
5�C"O�9�����lP���.I[e"O8�rw��9V�b)��H�;y0E p"O&A���O=0� ix�n�&h��'"O$t�e�q� �e.7"mV�Q$"O� �����QE`|uئ,	�zg�$�"OB\R#�(h�\�!��+0YP[�"O���wbV�q>(u����2�ib�"OP�*1��_.h�R�[(�0�"O4M`�A�:
�X��BV�|(���"O�	�w�ޜ|uR�2!��}p�Œ#"O���L��o2��;�EO*IX`�c"OX�"c�)�dL	�EA�N�Q��"OXܸ�JR]HX��+�^��0��"O�(24/�!S��ʋ�)��b!"O�tHR�.���IV�C� �^�%"O�����v'��4B�j"O�a��ңBģ��X�}�2Y;�"O�ݩ�f��,4��k��v̂�q"O���Y6P8�)�+��_f 8Cf"O�}�r-rȡ@���fY�	B�"O�T��`��)/H��H�{j��w"O~���K��y!-pR�I0"O�8{v":LuEp�nR:w����"O��ԉ�U�\�⦤Ktk��0P"O�Ѣ�ʀ��4�[aD;'N�@0"OH�{�h��j~N�/�f�U��*!�dU�fB64{�ڊN��e3�R�/�!򤏌H��I"` y����U"]3^�!�V��س� )�p���E>�!�Dӆ���@�%�
l$\�m��Y�!�D�1gV��S#КX[(&��
�"O6qT�%8�X��&��@���"�"O�K���2|��(�P(��e�� 5"OLƀK.���EI��!�h�#P"O`��6Q0�,�q�W�Z�tAB"O1�@0p��Tj�E@$�z��x��r
���D��/,5��*�cA U�@A��zGa~�NN�c�\�z�-S8Z�F�"�i�=^�)�omX2B≪p��L+UDD8Z(`�r�O?S�t"=٢KE�璉(&*!m�1�8�!+�{	hh�� D�`��7"O�t)�b6
�H���F�1#��i�� F�V!QI�����>E��4��ub�D F�j��Q�I4t����%��c�ʅ7|/fp�Ҍ<�Sv�i�Z����,.ӚP�cK������	:kd���,d�>h��&�)=a|�I�u�I����uE� ���;z@��
�*?v�QyO���D��uS��)d����t�@
]�O�J��G��d�&-HbH;Ñ~*e�N!2آ1�Gc�+4���]�<QĢ�+������װ:���o=�����d�j�z���S�yx��E��'�������[���@A�;���")D��[���:,@�Y�$/2�� �B��MST�(zK���	R�U��Q��8���� 	L[���T�E��BR">lO��������J�) �2 ���;� �9z�pR3+�9�hv�_�#�"����*�rHc��N>Jr�f�m�nc����J�ʨ=�%�śzy(� nh��S0\���d��%��@��O $�C�	>P�\	M�&1_����H�*S����`Q�i��Y���0�t�OA�:	gL�ps��g��t
Ȓ��>C�	7[��Ua��ֱ*(,r�%�._$p�ٴj,R�8�K����ეຓr�I%/I�a4�<j��@qn�A�����!TgV��Mo��;BĈ�?�`���[e}&�:%JϑcČY��'��`B�p5P�hF*� *��Q�#��4�Ō:aj�(ՄD:��'}_��9�.�94�h�jЍӘG�>C�� D�T�P�B��l�EУ�<k�V��d1t$�^�0n:��<��ȹp �EbK�4a�ȴ�$`�<Yw)�Ut�:��;��Q���֘5剪V��`B�����g��n��U�/Y����@��Q�t���	�a4�2u�~�#D�͡6�Y�*�=�� Q�O�PC�;}��s�#ւ�<Z3�� ]��p�_=<Ntc>9�?v�*���#�b��0��4D�� ��{0k\�EH�tB���g\�O�,@6�����O�>�AcL
�z �YI��32\�* ,D���E�0B��[���S�����l&���1'h��IҴ|����X&��8�FZ�%vC���U�r��$��x���Z�8B�I?�.�+�mȪ-���͙B8B�.P`���9(�H���
)��B�ɠ}���1V�|(>Brf��5�B�	�N{&�A�aܩv&*
�N�}q�C䉪t��%�$G�0yN2�"u \v�jC�	Z��R@�#l�J��L_
=��C�	G�����_�k2��"��.�C䉒���Aࠊ8ƥ�fƝSb�C�ɄS��]:���7-�-�D&�7StC�	������ߠV�v�#"�.T5pC�	�MF�ۣc�=NX�1��S�a8hC�u挽�mS�3,�iR'�bz�C�Ʉu�X�#4!�4e匠b�eƨ�VB�ɽQ�B�
r�W4/ڐ�{��()"�C�I	^��U��ቲU�N�ҥ�:��C䉪v��=��k�LQ`�AF��;��C�/$���� A03P$�I�$D���C�	�4vt<��g]6@0C� �4�C�	)V�ڵ|���"�Cy����'�Э{��K���Y��%�9����'~�A����/0�!��C������'=d 	�z��ң׵}��0�'��E���j�^�z�B�+|0����'�U0���`4`���>~Rb�!�';�)G��G���t
�wf6,j�'D����þIBX!�	��t}0�'��)AaL�4�|��(�/f�Ź	�'�.,)bJ{�rdB�C������'��t�BMO&H��@�䉼=k>9��'��`a$"�4�B3�L<+��y��'��Mq5�î1�L����  �n��	�'�����(Rf��w�SM���'�p�J��޲_p�0ǉD56#�=��'�b���
�V�>�[�i�'&�Dtb�'���� �x/�)9���]r]��'����h[?��,�QJ \	���'x�Ѱ��=�$�"p������
�'��݂��E�ZD�%{c�	
2h<�{	�'�9 -;����b�5tʠ��'����Ñ�2x�er�dO�F&d��'��dm	�}�.���f�=�
�'<���$J���3-N�G $���'|�G��2�x���u�	�'`bC��[��d8�,�B�n �
�'m�ɫ�L�z-����
p�"M�
�'x���LxXX��Q�m0 ���'�� S@� c���@�6�X
�'�v���jE�^�#j,]�<m��'.�&bC*
g��x���c�A3�'��J�aC��x`(�(�$mB"�'���)T%5H>������zK$)�	�'B�8�E)�1F�B��#mďh�ɠ�'�@1 ��n����tj�t(��'p��"�Nw��KT��+g��	��'�X�I�)���J$�6Hp;�'f���T��FoA���C�JC�Op�!U���D뺕�6�ًf��%�t�BgQ�΀���#~%�����#D�h��	�i:\%�0j��AP��k=D���n�b�T��tL��1H=D�� v��L�z�������B���;R"O"����P 20���	���[A"O��b#H�:����K�Xk��Q"O��X�.]*7�K�Z���O�<�yR��[��2�[�*��̔1n
C�I�2d�tcE�]mx���Ɖ$�.C�I6:��M:0	D�&@	Tm��	�B��		ؔ�*�K�5i��|�vіJ� C�I�^Kh��E�F��ƸR����b��B�Iq�pX�e�)C����pO�kX�C�I�!��4B�c�:`5p�M�' xB䉏2�RT�d���B�L]C�� bB�I�l? �[�Юj��Lе��s�VB�	�\�%��:\��H��/�C�	1>,)�4L��&e��Q7�2��C䉴=�:����S�"m��f�W!QPC�	�C��R�[5L����B��&�B��!@��[��H�bD�aj���_��B�ɔ&X���?u�����`�B�	�E�h��DC�%u�@�����B�I3v��Ѱ��9�Hxp��&	��B�ɊCN�=jF���9qF�� ��B�->���s#ʅB���O�K�`B�I.PĜ����J�n��j�k��_PB�eB(Q���W�lq"T��3XxC䉶�N�-M&i9H��M g\pC�	�#�L��ª�5?�:��!zt"B�	#3��l;��%����-�gg�C�Ii��P�dK^"�|k�k�3��C�ɴIC83����ztH�đ/f�lB��-4y��@M��0@P8�g�`B�	�=tY"���%B5�m�3�<��B�	78ɊI�R�/|̩�3&�]��B�ɪaN�8a�i�-��e�LǱY�C�I���ţ�b^�8��XS�H��C�I$:(���$B��T�����5BXB�I�&#N�0VN�n&"�GE��^C�ɻE�Zdt�S�W��y��y?&C��%Q�f�S�7Q�ꈩ�!_�W��B䉁<�$��B·s�����_�_��B�I�W��Б�	�3,!A\B�	�+6���ş�_�9`u�I J�B�I."��3@�q��K��ü4R�C�I3x⠭�w��)Q�p�EBB�S��B䉬4,x�)��ڛ_nL+4���C�gVR���"e��<I�蘘^��C䉤O�m"B�6^O�¦lհh��B䉰(� �	f�y�ѡe"�'EQbB�1V�Y%�����P�ȗ�9VpB�ɗ>�1�gƉC�VAk7�J)B�*F�<9�b��<�)���'�PC�.A�J+�R�Rw�`���ƙK>�C�I�}�hmފ)���+��� �~B�(#h�X8���R4* G��=D�B�ɻ��M`R똫2 �)h'���C� j�R%����;1|��RV �)e|�C�;SA��٠�	#9�h�	Ğ��B��PR�5b�i5�$��/B>Hb�B�	:f�е�P�h�@����,xK�B�ɤ&c���eJ	 g&�R�Y�B�I2{,���V�L�8}:=�1(�l�^C�	)l�1�a�6h��8���E���C�	�=N����ϐ*& �i%32C�Ɍ8�f*s���3��q@N��B�)� Z��6
�:=}�+��UR<��"O���B�:Z'v��"��2GL����"O,ݠ��ZP�R���[�J�:�"O���)�)i~�8�k	92Ȃ��`"O2��eR%������:��uv"O^�����z�r�"�+��G2y��"O.��!c�T�VA�I�' 4��g"O�@���Q��
�"'&����"OP��R���0�`Cóbx���"O�����W'6��U�DD�Ah�ra"O*U)F)P�'�p%��LZ�@*zU�2"OLH¬�.fr,�f�,	!̠�"O�8�Q��� ��E�F�T���"Op��$�͙ *>(�&{���)"O�P��гs|��d��|1�ô"O�����D�e����0��%)�a"O�i����(N�t]�7�]�q��m� "Ot�)�K�D{,�7�	xhtɒ"O�� !��C��2�B��&@<yГ"O��� �DJ�zbP�A#h!�"O�yiwEN�C�Pq[��(:��M��"O� �G�?��t��!��D}�6"O�,y�J�o	�y1aM���4z�"O^)%C8E��U�am�q��i��"OP��'����8	tB�!"O��ؠo٩Dy�́�?c��Z�"O�0x�od���X���(�
�;A!�D��>��1���\H��[�!�Dz	�vNB;U"�Ѡc)[�9�!�$�d�����v4=�u���D�!򄚄`|m� 3m�Z]�Wg�2j!�d���;!��'vbH�*'H/Xa!��F�/v�AB�x��(9w���H,!�Ě(L}Q #��uB�n��	!�DA##1�
b��B�:f�G!�$��gɠ��"+�b58���7�!���<J}b`��eҺ���)p�݇ȓ�0� �V�E�~ +ע�	�bɇ�`�*P!ϒ�5�tP�*NT�D������	�&|f�PTEA�q���hˮaO&]��=�vj�QGT�ȓu^��#�b� W �J��<cרM��V�c$���'�QZ4�	�}��_Đy��	p���r6�S�~�����s)jMzqCF�~�x�!*A$#�%�����lZ�w?ISN�&�RM��C���v���=�	�d�>i��E��5�`]��l:y:�����o�H��/�f8� ϓl�:��F�]}��`�ȓ
o��3B��uIF�@<yC���ȓ,d���Q	.r	�4!�l]�8Rą�M�ǁEGU�wO�)�L�;�X�<qEȔ>L�I�T�Az��2)WW�<�"����]Sr�Z'�f$!#Ej�<9� Y�W�H���Q�S���d	j�<A��<IْI:@�'*uB4��j�<�)�3'�9[��&����ׯ�b�<����mr�C�Q,x^p�����J�<y�抏!�!�b�+jDԙ�B@}�<��EU�NJj6(�&a�v}	��d�<q4�� ��YW)�ks��B�l_�<10�9V/��8'O�W
n�T�_�<q�I�j:8�I�OK�U*�`�5��[�<iW��7��!��%�}A�$X�<� $�Q	A.n�XDr�m��a"O�])�ś�hJ2��� "Db�	A"OtZ5l͛^�9�o֠c��X��"O6�Ї�IK�(@���C#��p"O
;��;<�B
VBh����"O���
�;^�b J*'e���"Oʔ�b��30�v	��d��RH|��F"O�%˶�ӏ a��'Rhy5"O���5@Lp��PG���Z�!���J�h!��ۻp�aQ�K�'r!�\��ra�B�4A���)�;!a!��Q�~ ���w�]��y)��D!�	�i���z�C��s���	�\:%;!�߮D��y�M�A�BXu����$��4��s�Ɵ�7l�d���yRŒ$F�� ��*P͠@�y���NM:xRbdө'eB����6�yr��	7�p+D(�:�ڸ��(���y���*#49B�K�2�5J��ӏ�y�)عV��"&`�HڦI�y��\_���5���.��6�״�y"$�=
�%8 %|8"��Kʤ�y�"� l�|	�.ݴy9x)X�%���yBۿV޵�`��n�b�K��y�B�M�hi��M� 7פ�O���y��0m�jy3��Ų)A �h�L��y��Л5�X��&
�4d�� ��y�Âg�بS��������"䃺�y���C!&�aP�LH*Lx�Ѡ�'�yb�=D�	���ʜR. �{-��y���px��Z�%�Q��X�5��"�y��1u�1W��4���10O�	�y�䟚mE�ܛ'*'2�^l �fU�y�G��yY��*�F� �t�H��J�y���1��1���*:�Q쀰�y�f��¤*�+V��(�s��<�yR�G#Oʮt�p��y��)Ӣį�yBh�-1(����<�d�Y���y�!J|�A�m�2��ʄ��yJVx@� ���*��Y5�	 �y�K����q�/�d]�d�8�y�&�*j
2� qN��s�Ԥ�y@^6mW~���ㆆw��@�d�yb��w���2
�r-K���y�� l��P`�'G3q�����ǎ2�yrJF;j��];@�kkʅ�`�1�y��V�U �Ģq�|��p�<�y"B��/`�3�EЀj�V@աV��y(D�{z�|�QK߀]�vͺ����y� 
�0�E�L�8r!��=�y^H^p����� $v � �T*�y�L=��RE��v�����yr(�&�=�7�KkL8Ѵ%^��y��
��H���K�av�ڄ�Ӈ�yB@F!K��%�L�U�S#�y�"�B���a H�j$0�*
��y�mP�|��ѳ H#98��CG�S��y2�!�
���@�+�\�&��+�yr�&,6(aګr�+v"��y��C���Kd�����yBӢ@Px��!_-�X�+�`^��y�#��E��-p���\ԄX�!�y�&A6~2t�&���ǭ�+�y��Y"E�4�J�	�	&��k�Y��y
� ��9��%N@��%H��P�su"O�$�p!X�
d+��x��"OL���/�43B(Rp�εL��)�q"O�b�%�PfZ� ��I&_���j�"O�yɂCԳT`b�sb����V"O^AT
V)�6�� Y�c��!��"O8�@�d�)�ޙ�ǠW�wz|J"O8@�3BۛsYj�뗏�kJ� 8�"Opq�2&T�r� �v�8q,�	p "OT�3�J�.�|-��lY�K��;6"O�j䆬a+(�CG��8��%ӆ"O8���ZD`򧈆�c��:`"O��@B� R�s�G����t"Ox@b��զ�Ȥa�l؋6)�E�U"O�'b�?�<(�b���k(B$K�"O(	(��ήMX��D%�-W!��YW"O�����	��!�!%�M� ��"O���ZL�F�ꑡ,u��Сp"O�Z6+��&d�4�`.�r��A�"O(P�Oma �g�.g�:P"O\��sf[�A�����Ton:Cu"O���qB�,(\2�2a�Q��a�"Ovd���X���yhf�S��"��S"O�ͫ�o�{��P��@^�@ىu"ORi�ӭI�0�-@r`�/-�Bq�7"O^ � 
6%I.�i��"&����"O�3�F�=a�B��H�T�>4��"Ox�9���rU4���Ș�Bo�	�#"O��6��m�]�%NO8lO���"Oh�zA��95��s�oںh5&��"O"�����g�� iq͕�lr��"Oy��J�m���6��.��y�"OX HA!�-@"6�:v�1tA�X5"OȌ���ԋ}�Np��/�x� c3"O��M2I	��H���H�1"O~�cQB׸@�!j�.�g>�zG"O� �ĕS����!���T�*d"O�%�A�??�����KZ����x"Oz}z��C�HQ8�R�KO�e�
�B"OFP�`�"z�`A���4��8�"O�i����=wBvH���^��$y�"O�i BA�$�4L2b䋪Swޜ#"O�L	e$F�}c����� �@�h(��"O�Y��*f�� 2R�7I���a"O<l`��?&������H�M�
8��"OJ|`W�)&Mrl�P���"O QHT�\�k���@c+�����y�"O��B��wʤ�q䇴�zh�S"O��QPj�~1"u���:�c�"O>LY��(a�l�����?���R�"O�PHp��>m?�ì �~z�4p"O�1����k�"-A�Adi��@�"O�a�(D* a � /gZtAC"O�]�q�^��i��]@<<��"O�@�6Þ�4f��#�*/
��U"O�`5�]�LfYȔ$^�qv�Y'"O�)�R!o�*��l6�=�"OfE�v���e�n`(�,)l��"O��)�/4)1L;c��j����"Ov�b�!��;>Z���W�vh�IP"OZ���՝w�p#e�&d��Ї"O�̀&J\~�#�';_wH1+�"O��B��
� �@p�����N� �@q"OԝyvD������� �;"O� �d���˾y�6$� ���Y���9�"O���E���e�V�4v҄�"O�,���H1aa ���I�BIB�(�"O:����V�d�(RO�����"O���BI[�R�B�I`Ϛ�*]H�:�"O����H5l�R损2U�� "Or����1ۊ�af�\�>*�� �"O�\;"��Nq=p4(H�Q!��0DB��4�fd���`@�^ !��A1��5��ǁO���� ��_�!��I (�~-�p���(�|4���M�!�$��c08!��[13mf)C�/Y�(�!��z ֬r��ͭi:;`K5S�!�D6I����J�"���:ro� �!�D\�h���  �x6\3��K�!�DQ�P��|��Ŏ-msr�Wd�
 &!�(*?�|�����*�,�[�Ԯ.!�K�v��M�'O4H��mS�Q�d�!�Ód�0��"��+J�E���C�K�!�D�sw���5��=��S�H���!�dA V0�#�G��0�$�t(�y�!�D�.3�-u�ָ;��-�'�T�!��6N��ё��b�
HHwT�u�!�D�;~I��C�d�6
�@(36  �+!��^�t��(ył͋�ĤPb�ӂN !���D�4����
�u�^����g!��ǭVL��1���7�(�4�Z:�!�Y=n�蒯�4Br��pb���!��MT�	�!��A(h�z��^�u�!��!Ia�Xs������9�B�� {!�d�jk椡de��M��  	U)
!��,,X�r��ŰE�0����_0?d!�$��~�P�hV��P����Ťc�!��]�xS�D1*=HB��d�!�$@3RW��3G�3o�D;��W.!��ıB�`�FZ��� �fʐ:�!���W�f�p1�K�_J$�+ �P�J!�䞯Y�(LҠ`�����$�ǽe�!�$�&*ǀra@�cn\��Q�X'g�!�D"J`���㥟3O���4hˮ5�!��W�h�W�����`+�!�8s��Iu�#0���Qa��C%!��
(3tF5�q���'��X�͔9!�DA�8��C�N.�@�Z���K!�)N�ZH�3/��9���>#�!��y��b��3X�4ٱ�L�%�!��|Ԁ�pgŦ;��� �H-�!�۷M<"�A0`@�"��� ��Py#�s�YT�Q�9�氡�
���y�F�o���b�?5�e.\<�y�fU�[h�i�k:~����%�y��ǅY.�1��>D�yj!,.�y2�-u>��%ߖSd^p��`Ŝ�yR�0�F])��ֵ��m:�m�"�y�G��hט�yv��H�x	G�L�y�&�Z1�q0�HO�-NZ�s����y+J���q򫆗"X�9��A��y2h+q�tid��=HUy#�c߽�y"�\<)�zs'�3�ċ6I �y"M8�xi�+A=+�N�(����y�l��N�2�ɆÆvā��D�yb�o��s���l����yl�=uL	rR�_���@����y�KK5-&�WY��y+�B ��y
� �4jc� �0���a�o��f`p(��"O>x`흒5_T	�'��fI�U"O���V���"�z)��̇a�9�"O2���C�"7µۅ㓗��Hi�"O�q����>&�����>%�����"O���t�վJ�T9�-��_���R"OT�`��VmA���bP�K�"On���ݯ1�άh& R�+���"O�K�҆a�.U�P!CT).a�G"O&�B��"��ٸ�i*�&���"O����E��a�p��#��(ό1c�"Ojy����&(��!(��_�<H�v"O��V�ҿ"P�Z�$C��"O��d]u>8��4\�.b|��F"OD�(��ʄ��+6f54RD��4"O1��Ğ�iW�M0��љ5FҠjA"Ot��6GM�:F�@�o��"O�u���!
�`�EE�*}��"O $XDH�\�T�aЄK�UF��"O��j���P���3�〼5�\�+�"Op�I�Cb)"�$�*t6"O*́����R�DQ�&+J�<l�"O�R���#e��q�Qr�eC"O�����$V�b܂S
O�D1D"O���ɚ+l��#�'0krzݡ�"O
�26�A�YÆ$�TC2#kb��"O�@T�
?+y>9Cu�I�`M�ljT"OHD�0 ץtO��S%Q`r!"O�0��C��`'T��ǥX�Ls�!3"O����ǶV��c'��ic�9��"Oly�0M�:8ƔF�KAlC�"O� ��M��Z�ذ�7m^Z<.�p"O���䎜�*֤����W��i�"ON<H�C��gxp��V	a'����"O�-�d2@ļ0�ē.���	�'��%��E(.0�2pZ�d	�'�P�D$��؛2�V!t�  �'��������/0<@ӑ�?rX���
�'?fH6H��Ԫ��etz�P
�' v�u���:�py��_�`+����'Y���ȝLd ��Ο Y�2�'� d�!̐�`b$
5��"p-�P��'bX-��y�~���灂f[�=i�'��Q�'D*{�h1Q��*$���',QI��*~z��y aֿ��$�
�'���l
���@'@AT0�KXg�<���#H��05K�Pt���4�}�<���
�u��j��5`)ҴC�I�C�<᢫D8`0L���-R����Q7K�@�<q0��n����� B+1^pA�pg��<yt�ɐb�x��⇨'��uD�S�<��l�����4O�>{��5{G�D�<T`���t,��$M9r�Z��!�ZK�<i6�J	<_���rE�5q�j�4G�L�<��2~4Й�
�g�"-���F�<!���~h��32KR��q�&�B�<�gV-��h��җ9�Ua�Bs�<�'��/�ܻӥ�}������C�<AЂ��o5�IC���,=mʍ�FGJ�<���gv�U�ŏѤp�B�Q��Q�<��C�:{�v���ˢaGF	�#�N�<i��?��$�% X���l�E�<�Ʉ#z-ά;�ǥ2z`�7.m�<1gH�I&>(�� �_9lܪ�jDg�<� �8�e�ȳ8���Ӄ�.+���g"O��Yӂ��_�:1��@4��"O��s���'{�+��է.�&l�1"O6�1Ą�P-��fI�D���#�"O���U�בh|:xK�]kX�Q��<+��X,%ٛ&�'f�TT?1b�$MR�	�՘w%�����H~H���?q���yҢI-r7���[uKDiR�	r>-��

�;x�@�lW�yŀ��u+ғZ7�df��5Ҹ�ӕI'Q��\�"�`7�`0�#ݦ"��L�g�"��#���GQ2㞘S��O�mڕ�M����Ɇ�F�rd�H�'�Ma�ʊ	r@l���k�S��?Q���DD��@veܿ(ra�`#RH��l�I#�M3g�iΛ��0)HV����N0v �&C�~�		�un����'�RR>mxCk��|��ߦa{�럈j��0��E4l���:Wc6_�&�u,K�HP��-A�A[���F-�?m�O������43t��5�j3�Å��l	�i�VTa �P��h�OS֙Qe(�2m�匊W��Ƥ�yAT2ȴ�BL: ����in"�R��MB�Ư`�R��/��i�B��I��pt��2$<r�b����	{X��(V��)C�qׯ�-J��y��0�h����~��Ob��x�	��lN�`��`C���S���p0����?���$e���?����?A��T���玲㭉n�+ԩ>�Z �q�P��X���BB:��S������nD�"<�E�J�a�h�yrd�>pA���̀�q�v�9eK�C�QJ'�����h�Or �P!�ҡ0��̕'6(չ��X8���DJ7&�H�e�O������OX}o0-���<q���d�~:6�kt
6/]\�����[!��:�P4�$��>�摹$�M?L��޴G��Ƒ|�O�tV��З��9����j_ 1��	�Ɲ�H�m�V��ߟ��̟���u2���ҟL�ɸ5-9P'��m��	��.#���АbD*]I `R2�UnLxC�lG�:G���c���&�h`��S�J���S���Y	��"Q�L����o�%u��떠�5�H��D��}�r�iC��SP#F�Or�KE�@��6��	��T�hHd�Ӻ�O�^}9�.ͳB+ʕ��I�NV@��'�(x1!*?� �����,{A��)�'�&7-���'��\J�is�j�d�O����)�C�T�(Rp�)�ّʮi��X�;���'��mӎ4�@u"��;pl��i��=�p��'U>�@��R 0�ه.��&XEz��00sF�X���1�"$J$È�uan$�[w�ܬ[d$^Ni��B��_�b��{�� q6qO�/t�$�O��&>Ul��6��P�-��`��u�F ��(ox�h������9���;���I��0`��M`�F�k����d�ަ��ݴ�M�C��(�P�����]f�ܩ���N?�GE��*W�v�'P>�3c�ڟ(��֦�`L-Z*:�ۑ��dQ�"p䐩	����%��UC=0)�Iۓ��?�O�$��0\`$c?x�b��t	5���S�iߊ�pDɑ7-�Ɓ�e��d������I�\}{R�~���RA7�;C H@�&\�|o| xR�i�����}��dw���)���%�;
�ޕqqċ�Ug�@�B����	ş�àT�'("��s�֕��-әx�4$s͗8tQ��R���M{K>i���bu� )i2�Q� ,	��;���t�`؞l[S�   �   r   Ĵ���	��Z�Rt���/ʜ�cd�<��k٥���qe�H�4��S66<q���\S�f�ث.�"� ��p3��yT��7%�7�T�E)�4Om��;��[yr�O�X��j1L�1dd&�x���+[�� ����,L�=/2}"6͍�N��$Q�샭Ub���

�z��I�xY�&Ԕ���(_�>PHP�N$Ap剁;��	)�d�%��f�	Z��1ɕ[؛&E�!�\Q��*m�yK0B�?�C�'���U�%I���� EHY����Đ7bxY��'����� ;:�8K�b�����Q ��2BaE!�ug[1��4�3̂�G�	�[% ���<J�b̊���<m.�fl�]��'��f���O�I@S����ny��� ��T��K� Pe��J%�����'�pYEx�Iз*�4���K�t\��{B�
�Tf�#<Y�*3Uk��^<����O�j���h���oӀ��O��A��D�Ÿ'3����2�I�@ph� �޴�N"<)�`,�f��!�K�#��Eva�
�Ƀ�h����>	g�%�3���{r5�� �4�2tb�,��On��'C��Ex�o�e��i:~�W"��[��b%�N��D`�(�w,�#<y�n�OR��S搿BE� �o�/:ty�"�ï�Op J<�4ϴ5�~��a�0j{�!�GD?��8�J{�OD	[7�'CX���'Y=�8�ٖ�EI�MQ�4s��X�'��P�h�OxM+GZ���K?�ǻ�H�� �8�j��$ʌ%k��:Ӌ$�I�Nr��I!�>yqeD�$��Q15�\�R���fi�G}�JV�'K^�Fx��N�$��4�vlI����C�5�y�'J/D d  �T3�p+s"ON�����O�8e� B�0 V"O�%R∛7I$XE�'cD"%�mS$"O��%f�Ud"=��]��{�"Oh��b�7xK�k�*?�<�"�"O� &�� �A�Ġ��/ժQ��p"O�LZuk��5^V`�&O��t��MҰ"O~���S����@�\�u��Ṥ"O�ٺ'hί|U����kɻN0�"O��X%�N�&{�(���Ƅm�t�+�"O���D,�? �$��V�Д=� |Q�"O��6� �&����R0u�#7"O.|�L���1C��F����"O2����#f� lʶ#����"O�q%=�q u#_����7"Ox��dG���ԛ`BA2z�d�9V*O�`�ň8W4���(>A��Y�'    f  �  �  �  #  j)  x-   Ĵ���	����Zv�L�\�0R�PΓ���	�q�v�+�`^�#�>��D&	�����S�h谎�lr���ꓘ�H�ō��H�%z���Q-҅M�����Ԅ~T��B6薒�J�Ɗo�H,�s"��N���F�;z|�<5	�/SZy�hɏry��C&�[��Lr�'�=���VD�1nT��Ѵ
�!b��`a� N�v�ð`�+����Ju��h��I�?��h�@�On�D�O��d��K�� 2<��N]3z"0��U�Ҙ	��͈�[����`:�O��
�K&~�49*��W�y���v[���'.<�O�%��=o�Bq�m��-k�-��X��+�O���:��p�ۻ{H��{��
_��B�ɋO�N�i��G2Gp6����{�6mV���ԟ|r�ˁj�LES�L�9�>���O�:SB6��	U��'�"�'� ֝şT���|��NR�\ S�Z.vb}��̀,6�th��4��>QRbm?I���6�ݓ�=�v�CFjH_x��cF��OHL�� �zY��b ��`A��\�<�"�S���r����'�|U�V�<14��"F-�1�C&D�e,nI+wf�Y}R`f�@�O�]�У�̦�������z�C�	��� �c���zV 4m5#_:���ƟT�	 �����l�S���O�~QSr�"|xr����Q�' �����W���qA�w�$u*Ѡ=].ў�؁(�OxuD��%"Y�$����0A���B5
��y����0fH� �24��`i���ɰ>9%��d�!�`h`r�'���0l�"�>���
ZK��'lbY>}���������,tN��I�'ϰ_�j�(���0�@K۴6�(`x5) �I����O*�b�8A�V���"��|$L�� �O⩡ү�31������(bJ�D�k�5:�����\1J���n߸T����?���1����'a?���iG�S��j��R5��H�f�r}��'�ўx�=Q�#=*���c�dA�R�5kFJB����+��d�<�/�`�K�Λ)�����,� 5�Â�����I��x��˦e�0��럌��ӟ	^w�2�Ԕe"(�x4�5N(�ٳQ��|��7m�Ob��%�I1kwz%����\�R3�F5r��Y���L�_�@�8�*�O��R4��~ @���|Fyr� 1���u�S
I!�`H����Gz��l� M�>����~���Y��`sf'��U|4\J������d�O���;���Y�́3��@�~�|xDLQ(�Vœܴ���GyO�~B���$�4Y�@	��F|Ӿ���T2m�L��MIW�<i�Ԑkc�}br���j#�WN�<1��G�D�A1m]r��7�T�<9����~�XU��)2��%��@�y�<����X�j$R��)3�z��B~�<y�Jȴk��ႄg�o6V��Wd�y�<Y�Tu\vq〯N7`-n;R'�v�<���ҟj�t!�+g��+��_t�<!���a�t"wX��}#�a�Y�<�5i^?X�4\(���*`���B�T�<qD3^^@�b��Xt����g�V�<I�+óU&Б�/��CL�+��Z�<�d��Ѯ��@��D%��+�(Ln�<���:K�	Q`I֘C��F�t�<1v�.!��QD�Y���N�f�<i�
1 p,<!t��e��Xi�ϒm�<I���(���u"�
*`�,)C�o�<)�ɉ�֤�Z�d��V�t<���l�<���O�|-�P'�{v����@d�<�!M-�� AlF�,c���MS}�<�T�ôe-�X�vLJ�@3鉢lz�<Qӄ�$A��tr�"�s�lᔅm�<Y$��; �zEA�iW�b2�y�2gMg�<Q�C�f[�}�RÝ
w7��h���g�<1��!���=t��`eH�<	�,�/K1��8f�}��L�ţ�N�<�nũ�f���Oց+�:p��_�<�h����k�gG��D``�]�<�&��'@
�)�tf��\�x�Y�<q�+�<>�Y��$�Z�<	���=q��Qy/ڌ)f�Q`R��Y�<� @0Ô��8��,RL��+68�f"O\(���� �X�bVd��i�"O x{��nr�IC�C�f����"O���re.��Pw)E�P蜝Qe"O����F0Wl9�̄o���;�"O�<
t"V) &bX`�z����"O�SV��3je*���jԳ>،1�"OB�B���.j��\�F��pg>�au"O~��p���5h$Y��I�N[��`�"OT�eD�y!� 8����
- �"O2���aŚ(�v�#��Q2,���D"O�`�����be�uz���H�����"O-�F��.V�",��̈́1b�L@W"O `�	]����˷M����"O����Ƀ�d��v�W-�68Q�"O�Y�N� G�R�IuB��oM���"O��3�KԃnBd	��Z6:��h8�"O\h�1@�R�r�;e
ɕ$��`��"O�T8��Z��t���L�E5�k�"O�2��2�h� ��R/#v���"ON�G�R�T�eQ`I�#���"O�	yW�>�֑p�
Z�>�!�"O��W�K��d}�!��4����U"Ot��8Y�<�PQ� �>���"O2�pA�=n�g�4I �I���$D�\��L�2e��ty�B���r��H$D���sʐ9��fn��(X�A��%D�48�B�`c^4˂%��2��h�q�$D��5��I����$T3�@�$D�`����t��1�'T�wp��r$D�ف$�4����)�R�;"F?D��k��_1C�ްP�D�kF����$1D���T�tyR<`�	g�h�A$?D� Y�ЋP��˶Gܣ1��|�3�7D��{�KV�:1ڬ��.FE���R(D��d�D���÷+�9d�*`�7D� �ߨ}j<�C�#���2�E0D�<��^���{�GÔ7��ᇎ"D��0q,N	#��H$ �	��z� D�`(�h��s�����9^���4�:D�<�!*ٝ{R`����6�LA�r.%D�h�Fb�&w��0��Z+"�5ґ8D�41���4:8V�`ӆ)p�AA��2D��Sa��x���b椗�O�¡9��0D� ��a��e���C�)wu�"vH4D��ze�3^�1�Ƥ"�ڑZ�%4D�pb ���q�(t��
1�e��1D���6g̷V�� ���]���M�ס?D�<	1+=M���ZW@�/R�%{Bi;D���3g�3̠Hr�Ό3~e��`d�-D�L��S�[ʶ;cUΙr�)D�d��Kɵ`1�	j0��Sfd�k��(D�t�������{e͎�:�D@���7D��Jtɀo�,�e)6'l�z�F D�T;�"�?r#���J�5tk��G�,D���"�F>~�"��	;����*D���$"
v��-����]�6a(so&D��q���0$g��G"��(��K�K(D�T0�]Z>�ūǠ%tp5�4D�\!�k��_
��h����&�.}Yp�2D��[7�&]��pA5Abp��;D�L�2��1=��1A���Z;�{�*8D��q&$��dR��VZ����(D� �v�^/_;V]+���![<ֵ�WH"D�� ��A�.Y�|`N4sTo�c�Z��"O��{���%"ڰk&ς?�����"Ot�Hg!I�
�q'�\_�E��"O��:��T6|L|���;(*�%*@"O�1�L��y�.,�ԥ�>U�H1"O��1&��aou�$�ʳF�LcG�'Ԟ4HcR�ܩk�o�H\�%aH�b�%�@�&D�L��E��6�
�#�Ɣ�
���C�%�	�qu�c5-�w�Ogd�ڣO�"vAt J�a�+��8"
�'�Kȹ6jS�e�	#N�pi�	_)Q0��i��p���<��aɒ!�!{C"�?��,�UJ�hh<Y���6*
�ːʈ$D�&9R1hGOx�m����L)�I@��'�`�c��$>�hc�N�yF�9�w�H}P�Κ�<��bw 2Lq�c�S��s�A�&L-�t"O.L(s�Ν�r<�&LǏD$a�>yE��_��J�ƥI�ݻ��W�h�Q�Ԯc3^p�Z�LC�I�)X���#�x�F�Q�(�����;�B��凐7*���2�3�$��^�A`Ώ�s���,�)�!�$��)^�CS�G�i��Źv��b���S���t�z�b�L�+W8�"b�'u��:d�V(M0�@�5ޜ$�`��{5Bh�Z�Qp�%k@Ӝz\\�t
�O���q�
N�H6���ݶ��xr㄀QPH:!I� 벭�� ������ �ɲ��#�J�:%h�#T�����ǝR<]j*��j�@�t����yJ$N����틁y�(x{�KΥG dA���ȰH[�n%/�rȻ��4�#�D*u�� ��([����j�o+��J
5R�D���<
# ]��� nG4�{3�X��Pȡ4
�%x 	�rL#<O��3�菃J=�Y9P�;ZM+��I��*��b�P�sn<Ej1�*cl�%��IзY��!�/=�\��%"و��x�b�k�1����-�!Z@d����BXv�]:�`����Z�*ֺ/L���t��2N_@����:,�d��`ż�y�o�3�KAl�Quؼ�s�R(|&�5럑TD��Q��y�(Ă���y�fƒZ���F��I�L�Y�x�nֲ�QZ�'�
33.\��iH*+N���h�e���27�ҕ-���ӓQ�v�p���:s>X	a�ƇZ=�i��	s?�ʘ�O5z��2�ɮ�H��t��E����E��1}t4�;�'�A��ρ 7-�)��'#>�b�}"�٨O.XAj͞GQ>Uz���4=5]��)�b����D�!D��aDE ;�hL�R'P��8�H��SP�T���t���G����A_L -�T��ǯ��:�Di	�'�L���c�	0gF��R%Ѳ9Z�@ɔ9*�ƜwnĘo��{��J�@n4T��4]�������=���t6� ��'��S�*��Dk�К�ۤ&�����'��);�f֞bI�|��/�:Gej����\-Z�~�b��h
l�gdK+_Q֠+b�QH�<�A�I�o�`�� �է4bE����A�<Iwƚy�ě�� �v�2c'�]�<��ʗ=v؊X���
w�¹��hC�<�GɦJjh��hG-�ν� ��A�<q0GK1@������a����6%	u�<����Q�uK���*"�(�`� �J�<���Q�R1�o�#d�����P�<�T��ȩ;e�?ez|8Y��b�<s���Q�\� ��9<��`��SU�<A�
^��b��dB5j� 0�#z�<���N<;p=�dɌ�=��|��gMt�<�1��-v�ӃO�7cl�!��r�<�uO�(#�Uؑ�ڇ[�`:F�M�<)Am��P9����េ~TF����S�<颋�mV\���Qp��s�&T��8��Qm����LE�3�a�C�*D��س��u�"�ރb���!$��S�<�A Dz"\t�w	�I�L�(�m�<a̅2���if�X����Fa�r�<Yu�͌Z�u	Ι,Rn҂�y
� ��Q��E74�&�S�
J��ȹ""O"HK�H}�=�bjW1E�~�u"OJQ��H T��х��)3��"O� ���D�Z�D@�l��Q�U"O��4�Mc����v蚌���z�"O>���!^�9�vm�oT�o# �k�"O� C� N#�>L��nR�"n.��"O�Fe 0]����ZI7���"O,Kю�p����!���"O }��aٕr��;A��7!����"O�p��ԑ~`�ux�(�2�A��"O��c��:Rj68����M���"O:�+!@ƞy� 	s'��'����"O@�!Jɬf�hI�S��'p��"O`��6��� ��e# ��%b+4���"O���F�JT%b�
�3Nv�EHv"O����`3}݈1�e`O(Z� ��"O�\���	y�(�ᬕy����"O����I����G
01̡� "OF��
�!fh=���65�`-
�"Oj���2
ܑk�C$d6	Z"Oq���3i��0QvC7S�
2�"O$�۔$TJ��Y�C� ���"OX�9��7�r����H2R�TH�G"O&1@��@��Ӆ G�B��Y�"Oh\��K�}N�\c��� ��y%"O��9$Ws�Ƭ�-�<4��3"O��"��<?r�ڰ��	2���"O�=�¬�-���8U�ϼ$t���s"O@����=1b
	� &C��}H�"O�y0�K^�<\3�MJ��0K5"OV!p�吐ZH<4����h5V���"O0t�(*W�pA��>=R80�"O�� ՌD�k9(%ig�%1�ԁ�"O�-�W-�:dxB�C�E��W"O^D��8�X��S�P�$0�"O&�!5�^',A��P�ʼ4�D�A�'x�M9AnN?�0t���:>:x`�0C\�C�I�Y}����	X�]-�P"�m
�4C�ɥ6��@�T�˳R)�izf耷G��B�	�l�2�)��s1�1{�N�1'y��DE�L��!/��c�<Q:Pj�IQ!�Č�kj\��Cσ&�@W_�RJ!�dE�8��@*���v\� ��
/!�$�20�H��-�=\RT��RĐ�w%!�dI*B�.1㭆�,:ޔQ���$q!��O+���)�r�ĴHc�B"G!�D���;F�������"O@yqU�ֹew���f�b��"OuK������r ^�_��1"O�ǃؤ~ �|�T/��5��LI�"ON )QK#o���a�ę5����"O,=���T49d0�� �P��Ji;�"O0�!�B�=;YT��c�4d;���t"O�t�Da�-9!3Đ.v���b"O^�{ �R������=
�` "O�zb�_�%7��i���r��=��"O<��*t$��`K�V�5[�"O !�A�R~�2�Bǌq�`��"O�9����	�d�қ� m��"O��TkB�W�=Ӈ�Q'{�pD�g"O�tB���7��-؆�TS�p�8g"ON�a�:"�:-�R��9 �� )T"O���L])�+pdC�����"O� �X��hD�+Q��0
O@�i�"O�)���yI������*S��{�"O��x@��dd��C-Ou,�ۓ"O2d��-D�b�s�� h����"O��y�m�+m)�$���ّP���"OԐ˕�^�@%��;Lf�	q"O��ꒁ'{\5)ٕk��L��"O��0�ДvXđ�#�,y.Y+R"O8Tb�"�3[%X�
�rY"�C"ODa��9n�HXB*��/�̐��"O��)F24^t��#�KOb1�"OFt�uIݰ$��B� ?8��"O� a�]=d-f���@�cI�%��"OBP�"���t�{��R(*8sE"OX����62% � Sh
/)�h�"O�<�Ɩ0�dg�_/3?���C"O����
�T,�@U�A	�"O�}#�#;��C�+C�/�`�"O !h�)ة��hh���#��Tڴ"O\ðE�KP�� �Q���:"Oj�3�9�`I���1�"��0"O��bqn?P$.		�,�%b��B�"OF]��O�fz�h�s���X.6I�w"O^%Ia""8��-Q�67��s$"O�XZ僗6'�$�O�Ũ��"O&`�� ��`�r�r�D4PDp0G"O��5cNppP���wF T��"Otȉ�F03���u��4Z��c�"O@�,��`���0�n�!MQ��2Q"O�Q���W�m��H"��J�P�&L�q"Ov0�%IT�WfZH��,K�jJ�P"O2�Q���KY�5�k_�yL칑"O���ݍ#�~�p�
�*/H��"O�h��'�-b���p��82t�U"Oʕ�f��A���{7�]+.�Z�"O�X���P�衙FMm><�6"O4y�$L�eR��
�琔��r�"O��s���E��
���8?�]�&"O��J����f��#C2���4"O��k�N$]hI��JA�E� "O"�{�@)z�A	�0_���B"O8q��J�P��Q)ب6XZܩ1"O�����K�QXR�N�E��"ORP۷��4lp����FG/C�)۔"O�$�QJ�F{�,� �i.�� P"Of�g`��4�ȡ�)�]`<��"O���`��>3��y�)�4n��)�"O�d9��� o� �a��/Zt>�c�"O<@S'Nt�����%S�"O^-��@ݢN8�Mip)Bj��kc"Od���*M!$��|��I�a���i�"O���H6��A9#�ʝ:`|X�t"O��8R+�";��1�O2gJ�݁b"O9�S�T�2oV}� i��Y1�ġ�"O|��㣉7�<�b�Q�Q@f�E"O�I��XQ���s��5(���6"O���' �qv�E*s�C�Ov����"O��@	��-�6� �%P�8e@qKc"OQ�ЉCB��%�Y�t��"O�S6%�	 P���k�"O�ps�C#�4`[V� #�F\��"O�yRUnH�:������w�I��"OT�a���5&�f"G�I�XQC�"OP�`o#Qq�0�BшT���ZT"O� �d�դ�"�L�"�d�6�{u"O�4À�D3n����3-�rܰs"Oȝ�5b�rB�#N��!� �i�"O>��� ��Ǯ�����;\��p"O����57x�Ƌ�"3�P)"O|I�t�A�)��b��]*��Rs"O��A`@�'�Z��&i�
R���"O, ��e��S�J�����r���"O0�*�#�.E�lF� �V<ʒ"O�fBҙ^~<e	A+[4!TM�c"O4dq�������"��rxx\��"O�9��R.Ȣ�RT��8gH-�r"Od��t%��~Y7�·vf�l(e"O�%�ɤR��2o!CE��C"O�H2U�[8%�� �$. �v8~}� "O���\�9���Z�N�x/bɈ�"O��Y�1�F�܈R! ��'"O�LJrhբŋV�q
�!*7"O��sZ�u�F���x��cc"OVL�1�J�17�t`�@)7�jh�t"O���R�AD�"��͓g� y�"O���՞�2AXd��6��"O�e`&M4���-�S���"O�Pe��?�b�cKx�+�"O@�bDK�;0$�@dĜ)[��+r"O�������@�����*q���+�剢"�a���:3�������b~��F�K=�y�0K2��3�I�R9�0)���<�?I���%m4I��^�W�6�Y�i`�U�ȓ:-�=�ba�>�$��vb�����'^����F�U/��p���h⅑�n�d�@�'��ȫFA�2'�T�dXj�,i@�'0����� �V�R���7-vxEa�'��!;�"$�l�� ��#3��10�'���0w舦w���XS	��+�6`��'Y�1� )=���d��%Q�A�':*�`an_25瞭�A�٠�0��'�BmX�/מuq��"`��>4x��'��*G��h���S��V�?5`���'�p<�� 84��P�U�8�����'�@�X���PU�T�!!F�i	�'
Ҝ���YÊ�ԏ�������'|}�#H��&�}'mג<|a��'\��v	y�2]�n��R�N��'��%є�W�r�Θ�)�#<��+�'"jMbp<��![� ��0�d�'�pQ���v֦8��E!��!R�'��P��-.v\#mMml��p�'����T%*���Z#f�j)�
�'�P�C�)^��%�"FZ3N�K
�'+�e��j�
�.u9�"�ZfBX�	�'�F�6f��\��9)Mc.}��'���')���n���Mh�
a�'��%ص[��
@���_��9!�'���H���%z��gJ�(Q�~0�
�'O��#w���-�ɛ'\~^�
�'�N����`5Ƶ������	�'�&ػ�w\@���J̆|ݲ���'�%Z�q�ʑ ����|�8Z�'���	���(��������np�'��t�F�����V�
|�P]X�'�0����� l@�Y5
J3qq���'��@�u�?L��1h��c
$��'�*)�cY�v2� X�ιiϼ��	��� ,���1Z�t��Azq�2""O&T" L���2Y� f�/\E��"O&�1KV	Gp�������RZ5"O�@hvj�&x�)�c0�^��%"O����
�70ѳA��k}����"OȌ@3�U;��m��@:�4��"O�T�'n'<<�%/������s"O9����(���L�~�>L* "O���IJ���Y�K�c��!a�"O~��FB�I�2�20�X*A��9�"O:š���eC��ꠋ�R�Px"O��"�.s�~-ȵ��?H��p��"O�)��u�͚�Ȗ4N�B��F"O�q)��N1%��X�ٛ3����A"O�����n��K�fR$%�b��"OX��F@�w��-�Ce��I�f��"O���e��rX�!vD�W?2���"O�m$�Kkn-�0�b�|�B"O8�sCD�7�����O4.��+�"OZ�����^U�A#��U�r��upc"OPeBcIυ8�X	�`� X��m�"O�c���Z�`m�@���"O����EՓ�����O�jg�Dk�"O)���$o�J!x$O�*i?���"O��8	�9yղ�s�Oޒ:P�"OȹV�@=&��$�� =� ���"O&��)�P�9s���$��hD"OR!��Ɓ�@b�(2� ����ð"OppX®�+X�b��d�G#+�AC6D��;'�h�$X��F�]�b��U,6D�D�k�;^\�a�gƄ�zt	6	7D�@�Ri�!wd��ABqaV,���4D��*���6Z,�}�G���00��1D�!p ��em�бa�����1��-D�АB�U$@��E�$-�;Ǭ5���*D�SBI2jn��ȳ���x%��`'&*D����R12�IZ��"-�����)D�����(sO�qh`�=X^ġ �.'D����1�$|��!�T������#D�瘛.{�X����2h�<$�6D�D�&&W*Y���Ԥ�'aPЄ6D�Hڣ.   �P   �
  5  �  L!  )  �1  �7   >  zD  �J  �R  �X  ?_  �e  �k  r  Gx  �~  ��   `� u�	����Zv)C�'ll\�0"Ez+�D:�Dl���q�6O$���'h4�lE� �]��P��v�J�hJz��u�iЛA���!2B�Xu	pݍ �'�?�"��?�[�O��A�� 
"T��'��>+�kJ�+��93�!�eglUٰ/�'�uW�ǒqC�T�'Q�� �cS?H�PU�㫍=d�өɅQzT�4��O$5�'�͓Obf��R��%QS(H��$�I��D����X� LX؂y+����IK! �П���l@��
0!Gey�'��ٲ�O�r�'& pv/@��feQb'��DxZ�:�'�"�'t��'/r�',���u�i���df���
�Q6�x����|p�H�b�%�OX手^^>�e!Z<Z�
��-cP��O<���PV���Е?�q�D�-�ؽX���Gi+ၴ�?1��?���?���?����	dޕr�(q7�`JG�t5��r!�O��L㦩��4h����'&p�ݐVj����4o�\H������CN	�潚��
�3�>����V���y�Q?9��R"[�A8 + �c��R0Ԯ]z@Pj��9�<�rf/[ᦡ��4|��F�O��A�!0d��FR,5��Q�NP�c� ��$sU&7M)iӂ��e�ˋD��d�I/]j���&-�*[�J�lښ�M���i��}2f��pƊ	�Ҧ�;@�<!���H�c�
h��.x7��禕#�4Oؾ���&c���Q�.�3�g�V��M&T&�ɣM��t�"�id��  ��dv�i�7-���ջ�a4#y0�0�.L�4^�y�M�C�ʰ���ijV��	 �ܴcq|=�vh���JEǈ�@Ũ�#�'��O��!pH׽>����C)�=!���Ot�$��֟�y��/�Ms̟�4����%��0IM#(xF��W�'�����	�|r�/�S���Ш�'�4��I><��(�2#S�c��8Dh��gjL��	)�R��e-��{�̼�0Lßt(f� �D���)`N��c�"2O����'!2�<�D,R�q��b�`�Yx4��7�Aޟ��I���?�|��'���嫃)(|QĊK;~p���b�i>�*ߴx�U(A���Rf� bh�1v[b��q�i�O��ȣ�$���?�$E�As�M1���)�����"T�T;�i,�S�������ȗ�<D��b-�G�tY��[k��� 7@-D�Pz֨]0X�L�/[���d�a'D���Bl�2b���ا.4�L�B�&D��[�̇ \�̈d��KB� �T`�O���O?�(�K�a���j���-0
U��F�<���L�+'�X�����*L�<�2*�y �s�K�	�^��b@L�<����6+Rx��$)s��ⓠ�l�<��aϕ�ӪF p� ��c��c���D�Dl M0M�T�P�	0�(=����P��~�'�"�'X���'r�'s��qAc�"�rq��� �/��@2�K�Xk<� r�^��0���%<O�PA1�ץ#\0����-�T	��m�9Z7�Y�bEH�b:ˎ�K�Vi�%6*�ў`��e��h����CG�x.�k K�5(8�H����<��O�CK:R�:UCUh�)�p� ��'�!�����쐘 �@�nfm�C�ԵW���o�����a�4��ȨnFθnZߟ�ϓC����'��a���YT2��	]yR�'_b<�&}x���q"������@��L�,�T�� ��ju��4�ˊO1X����>�jͪ���:7����؍_*��
�ì�b��"LX���q�'R�`(��?�Խi��
��vѳ��M��(��@��-���ڟX�?E���ӭ{F�A:ӈ�3K��tX���(��'�퓻�M[!i�2��3�_/7�0�֏"��v�|���D��0�����䐵�C2s��#0o��JA�(P��yrb�?]������^���)gC��y�͓.n?@���*��_�jtpc����yB��WWN���U�O�J�����ydK'I!�E��`�
�:I{T�T$�yR�+V�n��%وv:���bM�_]���|�'��2���'���'n�	�1쎁�W�ԒZϦ�t�^�m�IգG%����.n"2��F��^���I) hD`��ߥ;�T��)��N_.��&J_2���Fc�"��&$.�V��!��OX����¸��9Bi��Ni�Lp��uӺq�'��u����?q���?i���),�U1�	ƙEi:��6N���<1���ԏ~>�����¨^H�3���G3B�'B6-��'����?�'^�*�,ͻ8ł��7��CFP�5"��%��6M�OD���Odʓ��'��p�d+J�|��w䂺`�P!R�@�-��7�N�M+�2�?�DQ�@O�d�$8�eT%$��@0ǌ8�z$A'�΋X2�ɇ�ɜj=H���	M���Q��n���p}i���O��m�yy��'R�'���'��S��>� �e�?�l����X��8B�	3xR�	j��ѻ1V�(g�H�k�,�O�lo�џ�'vx��#eyӚ�d�O89{�-B��(�:"�����Ob���!y����O��Ӂu�B�D.�)� x�t�^/q�}��A1N4��J`�'��9ʍ�d˸/��j� �y@����P�o?axb�U��?Af�|R
�/:Ӧ 1Cŀ� ����T7�y���
#����+F�eO`���F��?�d�'�D�ْ`�/\?�@@aM�od���J>��kg�&�'�_>ps*�ԟX�vi
51���B���+W��bB�����.]��r������Or�'��*y���xB@-/�h��x�"�{1�q��3z�x�C�ӡ�h�^ è[$|�F%�ЖzCv8a3���R0d�OV�lڐ��O��6�m�gd�!nÞy�m��C��H4�'��'�	 ��S,V l5�E�ƢW���=���;>��vy�9��rv.M5"�X<���R��m���z����O��C!
�(1��l�O����O��fޕ�A(փjjv�@O
,a0P}��'��� ���` J�?��M/.�H�2�]�^�p�,�:|���q�شq��ǔ/ ^-ˏ��y�II�=���Y	�l���Π�?���i����A��Y�����ID�z���df��!#L�x�G{��	������Ù�:��'�?z��`w�П4��'����<a*���$�<P+@}��K+��G�2�[����ib�A��B?�?A���?)�D|�n�O���q>��B�-QX�%���ض��� ()�C�ɼf4E)��'���zDǉ�*���a#e3�X	�#P6`�!Ъ�p�h��2/S :�dAU���ȡ-bߊ�փ��/�р��8D����B�a�tÄ��Eo�H���*�DE��%�8���M����?�"��<w��U��d��>TRI��!�*�?���)ɨ����?�O������'<���&~���.ʷ2�}�	Ó.��aFxr�ٽ;�a㢋C�,�Ό:�(�0<v�֟D�N>�GD��.��Y��b^� �)���`�<�H֊�0�
�C����բ�Z��T���V���ȗZ ��W���|2�U%����f��M���?!+���)���O�@j�7Q6���q��)m��c��O����)����+�|�OP�q�%�q�x�ީly�Ñ�8��2�S�OH�`	�bGbS��ˠ6W�EP�O��:��'��O>�®8/@�<J2m�3=��ÄB9D��z�� >��<�L�4��+��8�-��>U���L;#ߪݩ��$&����	Ŧ��I某�I�)�D�c��ڟ`�	��D��Ӽ�`�5J��h�E�O�9�G�����f�P� D�ER�g�gV��� )6t�^�����3{u�M>1�	[���|�<a5C	=:� !a���'��ҟ@��������䟼�|�'<�.��=�ī[5"�ik��.!����>6Ѹ���fZ`�" �O��C����ٟ��'��*4�E?>�.X
���Y�*���ɩ`�\6��O��d�O�˓��'v��"5�(c�p��Č�C��#�i���b�'��Q��E�:06$IkQ�y^a�+Z1f5ve
�M���9��a;,On��g]�k�\�1��A�-bjH�jE e]��'��6�OB˓�?���B@R���%�P*�>!����%����L�	v�D(�� N_��ͳT��
:��'l� �>�*ON(rU�ڦ�I�<!�I�V�ĉ�Q��[x]��B�ڟl�'!b�'���AD�Tp�ғl7�!�6O�(!��R�<Q�M�H$|?9b��'��a�ai�s�u�� Ow|6�M&CF$p���j���]�Ȑ�Ó������M����?9����F�t�R(,�P\��-�?����?���?!O~z�y�J��HA҅%��"71s���'Lў�ӕ�?���4MHJ�HTj̏(������'΀q���l�J��|�٦��I4>6��&�6Gh�}p@��J�(��I�$���5�~=��.0_l��	r�'NT<I5��#�����,`x(��O΁P4�
H�&�1C�J���dF�D�ğ4�	��#F��ur�Ի��0Z�	��Ms��i1�S�-�t��,H7B.�R;֘cSc&���O���&�S���^$P�	�F�ͨ\y�WI�'�iuӚ�oU�I�I;rY	�Bрl���%���	/jnE�?�g�'T�`&c��a�\,˴`DM�f�`�'m����B��1�D�L#����'�"�z0(�1s�,��n��J	���
�'�0��*X�L���sgC/F/|Db	�'8��@�Ro�a���AdQ��'p�}C@�W�<P>�S6'	�H�6��/O���'ۦ�ѷ�>\������������ �̩g�R�cΙ�Cօ�JA�G"O`�����r��1q�♐�l�`R"O����^u�գP�@�e�$��"O�5�E�Q&)9� �3�k2�r��'��(��'? P�pÀ��bUA�k�'[���'&<�r!@W9+�0A� �P$��'dn�B��"ܗZ�zHä�y��P�7��i���L8A3����y�FE�N�X(� ں�0��U	�,�y¡T9A�h�M��,n����hO��Ӣ�ӹF�T�ƌ�Z��9Y���P8C�ɽj�:����~�5+Ӌ
A�fC�I�2@D@ūS�lwR�㇨QG��C䉹B�:��W�Ǜ�>lR�P
#�C�I#e\�P��Gy�.T�)o+�B��;$�V�04.L/
� @�+F́��?��,G����V����}�@k�J\ol�`m&D�cW���,�N(�C·38���1D�I�GZ��q"'29�����1D��Y��3���6Co�M�T�-D��1AOU!4N�d9�i�7!��S-'D������7�^���$JP���<�f��{8��7!ݤL6>�sE��o2�'�#D� 2u�V�=�*<�
�)ap���?D�� eb^�C6���͋�0�u�c?D�$�,����يS�H9=� �n:D��a�;|E�JKkY��X�5�O]��O�Ͱcf�9�����.(2Ub�"Ob���ʌh�v���.F�4�h"ON�Q���E�a0��ˉC�*��"O���5L֓Y�d��b�����F"O ب�V�Ͱ�9!�P@Ir"O�|��-�jj�����.c��A��ɠD`�~ꅉ�		lbw��F)0�%�IX�<�&+C�}� ��(��q$����H�W�<��	Q�K��X+MH���sS�P�<���H!k[�U !K�I3�h[ ��H�<�c�� ~��Z�.M�;f�1[!�B�<)0D�2i�>D�l�8�T�؟�h1<�S�O�0{`�Hz�=��G4";he��"O���Q��1>�.}(''_k`�ȥ"O���"U�w���	`�p!��"O2���CҚ� ��  �R�R��"O�����^gj�A�&E�1"O��y�ㅍPG��t���g�:�(�S��b0�,�O� �Q�t��N�8
�+�"O�-�AH�:����b�9O�)��"O��DGȋH�Ay�B#5�<\9A"O6bw��W�$,���+FOV8Y"O���#�B�@N�{q�҅^4��r��'�HY��'0bA
%+�M/d|a��[�Z��X�'Ɩu��*�P�Ra[rML��(0�'5��*@��.?��Y1%.�I]�-�'[��)'��!ʮt�tCP�6P��0�'B�a[�L!�
����46���'�Tq���~F*T�U��'z��8���*#Q?=�3,�Or�0����![���0�.D��:1�	8t2Q�a��]L���*D��(�DW�cqTȫ]�?�. +�o)D� �F� �5�:�rt�M O��1�%D�<�� yd��׮�V���b�0D����bT6o8((8�`�W��-��@�O��q�)�Q��Ac� @%���)X�c�Z�C
�'�f1*5�ϫ)$d�Sd\+pF�yx��� ����Ȁ�h�QH�D��D�4�@"O�s��1�5�t�� ��a�"O@�8�A�����?=:(�"Ol* ��dZBI�VE۴b"\]9�]�����%�O����!�~��Ӯ�5&�9�V*OJ�Rä]e������T��r�'� �:p�������A� �̙��'�l�r �P��T��`\�k\��K�'	6D�D��2+���p&�)j�	9�OpԑU�O�}�U!�*6ZQ$�u�\��"OX�q�Ӟ[#�<�� ӥ��}б"O���F�<�J�F�ʘ`j�"O6��EG'�:=j"�>�� �!"O*�R�H�&g�h�Ȕ �N��q��"ORu�㍞;2?$�⒡�&��X)d�I+b�~��F�)x�0U�FԄ/B�J�(Tt�<�VlIz���b�
_���q@�i�<��Ă*��2!K�����qA�k�<Y� ;F���Q� X$��a2��f�<	�D��Hw�@A,��#jjxQ��a�<���U:y� 쒁�./���3��WןXh`�=�S�O�pAM�c�2c���<��X4"O����O��v\����0Ö٣�"O ,2Ui\�4U�e�bͳ9�nT;�"O�x�(u �(�6j��{T"OҽA���;�2�2�� 
��S�"O\�����a!�z�䖐0#�^�x��"�O���@�K��� ��)Y%$0�"O�5�1��I&zXc��U5� �"O�(�#E�c�����x�! "Oz@c �-��pڰ^;EJ2F"O8թwn�3hʸ��NX�{�\R��'�(���'t�����UP5�6�W)L\�q�'!�]�G�Q�}ZȌqv�1�Ĉ�'�.P2���#p�F����|�0�'MR�� K��\;��.wp��
�'X\�&I�?\�`��Y��Y�	�'��j�K|���h!��PPH��Ě�zQ?݉e �?Z�M�b%��7y<�!ҩ$D��b�іeh�BB�c����#$D�T��Ş8�,�H��N; �e/D��gl#A���[E^�w����.!D��цޕYU�5:A�ϳ�X����9D���En�κik#HN:1X��#��O�ͳ�)�	����a��6e�0��E��"O} �V�d!اA�,Q�r��#"O��E*�ҤpT�\�Xm�"O�m2�#7Q��#A/��c�����"OF����дl>��C A����"O��&ED�><y��ݲ[Ԙ=�PU� >�OZ����K7z�ر��($6]J�2d"OF����97�� su�֘KK�`;�"O���Q%�%]dI�3��?�m��"O���3���	���Fϋ?@���"OƠfi�0H:ĚF.,�f�'����'��h#���W��$���ۢ�x�'N�������k6UI̎�VR�1�
�', d��i�I����Tj�1a@ <��'h�IP�E͈I��d ý�L-��'�|�D�Q�S��p�cb��}��|r�'�\�$���D��l�C�)u� ��䉃(�Q?e��
�8�"���I2*&���ӧ'D����Ѭ-cNqba��27q�y��$D����؊}X����됹��) �� D�� R]C�G�B1����KG��X�"O�)��H��n,B��ٯ���2r"Ozq ����$ <j�h�V�'nD�����;;�2D��
��O�}�S
Y�Z�pЇ��P�Dځ`S�)3�[�t(@U��n~0H�Q��w�t�b��/����{tj���LĨ#4�TBtG	!'Ji�ȓ'Nl�0e�1,����B��M����ȓ";�auFE$0����E	�@L�'��m;�*��hZ���hj��*�(<J���H��ɁG|�j$F�"@������[��F�L�^Tв��OE��ȓf$��P��)K:PH�%O+�p���+ �@���.J0VlzS��Co�؇�I�<��I*Bqp�J��i�p���-�E[ B�n�$B��_�ZXf���/3L�C䉽/BȜ���5�@L�ᆐ�Y��C�ɪYҪ��p���w��Gg�C�
q/�ˢ*ƿP���ѕ�W,F�HC�I�@\ָ
��xT`څ��C%F�=�b��h�O�F�y�Ҋ
�ҝb���w���c�'��x�F2a���J7�C����'�S�?HF�q��`F;�|�
�'�p��������h�`ԂJv�#
�'�6��#ػ�)�r�� ��-K	�'>�A���ڄ� b�D�~`8\{���T�Gx���[����L���S�#�^B�ɿ'�6���
$��Tb��E6�LB� ~`d`�A�X�/���ru"�m$FB�I�2\���&ƊX�j�+�E�l
�B䉚Y7��������H-����?tPB�I7Z��	�蝈VY������c}f=�	�Aq�	 Bv6��,^ߢ�a �K^wk��O}��H��m׮�zѳqS\���'˜�Ӷ�'�2�']by�GJ�#}�b|2��]�KZ�	lz>��� �!`�,e�g�G�c��e)�}�8X�
Q���hA��ЎMɴ�v!� tR����!�7m!	�킈L�FXh��DQ�%:��'"1��X�6+���!U+��k4ո�
KAyr�'a|�B\Xm���\�/�֥�q�D��>1�^��ꐫ��&s:�v�?3���Bi�<q%+��?q�ך�?*����+����G�-�b� �J1�����=C���$��iu������]RwN���ʧ��O�T�H�Ds>@�;g̳i���қ'��yŉ7��Eʒ0
��?5i �=�Ta�IL�KFvyI'm��ȣH�O��$1?%?��'���1�� ޠ���̕�TC�ԉ�'M^X�S`9>��h1r�R!:o�I��Ċl�O}��8���4K0,DI�OR'oBP�OW0\$2�'#�lA�Aj���'�?����?9���D��nL �a!��5 :m�q��$\&�@��΃&��0�+G��D'=2���R�7PЁ���_�a��q���	N����P�P rt�Q�e�g`6pF�?�ҏ}���<�Q'���(����!a�����\�t�'kў�͓3�v�I�-Gl���/�����[���P$h�D��r�*��-
=�	��HO�)�O�c��`T�<������K���O�0H7�'Фx�r�ͦ>g	��ZUTT�R�'I�`�#��*�Ԝ(4��c����	�'7�@�oŸY�ìɥ^�Vd��'X`�P��q��{�Qk�,�
�'OR� ,K�M>LU�3i��eǘ�
ߓDl��O�yآ�.�T�X�М=�T���"O��Җ�B#���B2���9�"O�|�Ԃ��^m�CW�,�T�XT"OȌ�EJZ�`2,ٻM9at^Q�"O����3)>�9��шq���"O�؛c�PB����1�=i7�dX��O9�\'$>�fuk�%ly(���'e��!��n9h��։3�5��'^`�r%��{��tمd�1�Re���� ���+F�X��-QFA�LhBX�"OP�H�L�Ԑ�j�l��q�"O�I�初<4�yx���5��@[�)G�O΢}��s��&J_x]��
=j�t)���nTy�GS�I!�eq�A�<$E���ȓ[�E3n��R�D����=n;``��fx=��ꑈ��q�7�_7Z�ޤ��,�"��a����1�EjN	I`���b
�E��_?���F\���	�'����(M�M�W�a�W����B䉿p�ZDE��+6T�5��D�Q��B䉞[�j%��$@v�cr�@� -B�I�k�P����>3=����6lQ�B�I�
�*U�u̶}�䌳�+=tlN�?Q2�ڜ0ڛ��'��9�����+~��C��*6�V����'�",�Q�'^��'�Jh���'1O󩇑>�6�Q��A7\��$���I�8�'b�@I�D�?�� ��ڤ��$G|2�(�?���)� ��bU���J-F�Y�E�(%�!���>9B�����Q�f�(�# eJ{��}�<A���4A�(�W̞;s��*�K�iy��'��[��O�Қ?�'/�%M�x���ǎ`��e�2�%�,��>�(��{L��똜O��3�(�	���$���U��4�1�$��([8ł5������|6��Oe�x�p;u��O����Du�� F#��Q�؀�T)��ꦭґ⛘]ҬlZԟ(PuC��xϓ��M���]�����D�yp��V�H'jQhO
<#���?�u�!��'.�N�O<�$�����d���r�
�ws���D��8xVL@jAɑ-&V��O������O�扜tr�s��n�K�ta[�L	H��E�:�l���G��?QP�����@�f����~�d�O��9Ox8@�B�4� � �Y�5(���şTs��Ot��^�fV>�dv�4� �?7��h��/��B�@R��M��OO�O0$�n�<�2@�ß��I$P��'�?����S*�,]b�#D+��"�Q�m�)y�dtٝ'�TM����?I���p��p�\�g��?nڮ1;��h5�
$s+�)4	�<����s���$r��O�O���E*gs�ST���V�̼z��G���4�P�̧f��l��4V-�U�'�����?����?a�'�:IњO/�<�GQ�a�&� �/�
&Ĥ�ڴ�i����'��韄�)�>���	d���c>[|"4��|�<i/��oJ��s�QF�Rv��i�	ԟh�	Пp�	�D�I�l��56�I�O�͢��Ƕ"Z������M����?����?i���?!��?���?��i�(?ư���� 2\���%Q�m���V�$��fyr�''�gy�X ��D,����q� �y�7� �S��MK��ۢedܝ��b[��>u�a�No}��'v�Z��K -vy��J۱-��!��'`ɪ����4�����%r�`�
�'R}�q艇V�l(�0��>7|��'��eM�J[d� ��2m�,��'I,��,G'c��r��BJ�ea�' E��]"B�*Z��#�%�y�)�""�B�yG�3N�`[�F�y��*9F����"SL0�M��L;�(O0D
�'t�Q���Ҫ,v8J0$E����ȓb��9a��7�H�����>k�Pe�>����3V���E3��Ԣ�#�H�m���Ku�i��.�
+rL����
W�l�[���P���@p��  ��L���0	�6(�>C��a��kݜx����d���:�B�='R�l��MNf�)R��I?����0�0X�藊T<�;�U%7&��S��|��?b|��k�/%#$4��enO�u��B��^�`$�]�"}�l�EϦmRB䉷W��h���HW�X6f�+hB�ɇ`���pt~mI)�H�JB�I�7�����D#$�Xaq�`G>U�>B�?�&��Q��>9�4�[��B�I��ٚ$�H�;g�A!�,`/�C�	=$��ᯓ;JĠ��4; �C䉕#�� ���G�f=�%9�� ��C䉾?�H�Ҷ&�0{G\�]Fr`C��U����Q)}��K\<X`C���V9��b��=����}{�B�Ɉq�,ݛ��&֨Đ��(vp*C�)� �p�O����� �텲9�V���"O�E��K�=�1���4pA�xH�"O�񪃾R6Y�g*V�cP쵂�"Ol�҇'M���I�1��cMj�q�"O��rvO�FȾH��;"N��R"O����e�D�\m �MI�����"O�HbP�h��u��M�U�� "O )���0<Az��b̒�Y
L  "O>���1\Q.�a�� !�@��"O�#Ҙ#���"�>Y<иk�"O�p�
Ѧ,EإKP�T�h�X��5"OF�Q(J�,�D�󄃿]��¦"Ob��#�J�7f��#�#?�a"OʱRO\�r58�E��K+f�Zc"O�"�\90�䨱C��&��ӵ"O����e6|��kc��!{�\j�"O\`�&eȖU�������X�SF"O�xY�)#�`I��C"ߤ�4"O��TD��h�l�@�>#5��+�"O�;�jY��ꕳ���4||�B�"O�T a�-����S�3�^��%"O�q��*��� �e[�}� � �"O&aJŎ�4&6��F��}����"On�Q딻iNl�P��1�$���"OL|�c��o�nh����?|��![�"O4$�'��<��p�թO�V�ic"O�5j'k�@M�lIt�����؄"O�i�;#I�y���Q�lp�3A"O&1�FE1~�6\�7HO�*���"O���O�h�d���P�� )t"O��t�"��Q�aG\Q�����"O"Ȣ��zjA� @�C��x�b"O��K�C�����L�pz��J"O	��!��^���i�9�6T	t"Oh�s��;|�:��G�q�l�T"OĤ����f�ld��F{B�`a"O����hD�D���ӆZ��-h�"O�8��Ņ�|I���QE���NXk�"O8�C�!IJ��G#P�uh�v"O��t-�NP��DB��DB4�"O�P`��.;F��G�\�)c���"O��@J�)H�.�bS@��&o>�u"O��(Dj��i�~����p���$"O�ZAǉs^���)�H��"O"xC����/�y{�I�l�����"O*xC(A�5����+V�JQ"Or�ڇ凊0�\�$%	��� �"O�s�NQ��ZD�6�>L�j�"O^�`b@�l�9�g���00M�B"O	Bwn��r����?�Bق�"Oր�FnV	6Lq��W�^��MP"O(m�ᬍ	��`9�k��E��;!"OhA	�i����5@��G�]5�y8�"O��0 ϯW�8��(L�Ѯ�H�"O��z#J3-�0+DGW�Y�����"O��8P��F��*�[�6d$�"O\t[Eg�D`�A,�j�2��B"O�Ii���15&!��	�@F�X"O�(��K�`CL�z��Ύ0
���"O(T;&�&YX�:���.Y!T��"O�A�G+�k�= `O�Hx�cv"O����&w(��+�\	���s"ObHR�f��6b�P��*{b����"O�x8��Ѕ-+(\[&�B:�1@"O� �T�� �W��L���D$:�X۶"O�x�@͝8J�@��q�7!�M��"OJy��_�2t)x�D�*[┸"�"O�Hi��4.���s��;Z�2a� "O�� I�$�*�qe��+��,�S"OL���; *���Jݗ%��L{ "O@h�`�γ=��(�J	p�ԨS�"O
$�0LA�+nl�ôn��*�i"O.᷄��08�%���>g���y�"O"8�0���5�gΓ!�*���"O����z�ԩz�g�U[Xh2�"O� 7IW={k ��֫ЌF��j�"O&���n�D�|T���=%7����"O�UH��U�X e�{%�kw"O\q�r���Dx���7,����"O��*s�ExM
����!:�4"O�-��M��0��S�(Zu21@C"O,:�Ĝ�!���b�O�rp�s"O���8,3����kY�`@�x"O�8+f��S�.�(pKB63=6"OZ5��bCkHD�F �l(F��$"Or\�����s�|}zq/�F���"O01�$��nr0If�ȼN�D�
6"O���"@�,����)4����"O�	�JL;Ib4t"�eP��f�B"O� �����^8qJ/ǜ]c"ON0���ګ̤�cHB� ��QR�"O���b 1;��T�6�X
S�^8p�"O4�	�NՋkWzka� =�F<R�"Oh�c��x��Y�$Ň,~�� "O���.��e1M1CT�Zh,I3"OL)k�{4��ro6I<M�T"O�8�ѥ�<+�葁�g�/8@`"O̠�6!�K�N�#�=.��4"OBl��䍵=t��W/�%q`x�'"O.Yp��B0K�������'����@1:x,Ro]�
C�i�	�'���!oZ4¥�^+4낭Iw�E�<�B^�?�&'� |�Mѡ��\�<���X�l�M�r�ޚ~������O�<����w9�ըAg�"�w�PN�<Y&	�=�(�"���aT��%�FT�<Q�G��^�\Pd^�p�|�DÖM�<	cjN�F��0PՈD %���`�q�<q��.!.9��Օr�e ��C�<i��9p�MЅAQ�6���DD�~�<yD� v����@. ;t��Go�w�<A��B��M�K� ��5��,�o�<AkMR�` Q�vU|M�7�Wn�<)�^z��D|JA�`��<q6M��pD9�ܽV��(�+�{�<Y��4U2Ҁc��ɺ|�0Hq拆{�<��T��x�Ҥӷm��Xï�y�<�CI8l<����1
�|l8��w�<ٷ/��u.�kuc�*&2��!t�<y�gU]JH��S�[o�i9QF�w�<)���_����C��V�����q�<��u1�R��Ǽ
j@���[p�<�`,ݩ~�Ĉ���X�=K#FD�<IU����qBȞLO~�rc��K�<�m���`�H?+$,�J���p�<�'�z�^�rT)��O�����Gv�<��T�i�<v�w{Dr4��I�<���\g���s�@S�0��i�!�Jn�<� �̀3$��b�����X�����"OJȹJ_���qI��$|���U"OjP�P)�	~.���CP#�l�I�"O�a�4�P+Z-lu������u��"O|�⦀��lX�6L�$B�y�v"Oj��.�Q�R	3��ސKB�J�"Oء�á+9��|(�l�?H|��S"Om��ᓵX�* Q����C0�h��"O��*��΅�yj�ɯ��"�"O�Y�p�6&��*֩Ε}��a�"O @ӧ6��9SI+2���"O������(&�y�(�9Tm<|��"OdR��S
7H0`��$����""O<PsČj�� Z I R���{�"O�Yc  ��%��E�����q�"O��K���5&a�a�>�B)�"O�-�sȗ�\X���.� 
�Դ��"O4�7��C��
��\�i�>Q��"O��S!cP
*J�Ǣ�����"O���c8\���&˘�0�Yq"O(�5(�1g����C�U	^ԋ�"OY��R��L���T'?YRy�7"O��P�(������_Sm��"OPq
�\;K"*�OT�!U<�y"O�l��N8y!�t{�.Y�~\���"O��+�n8xN �@�ѸP��	�"O�lBr��)T� t��d����"O:<��)^@��c�O��H�"O���w��|�\�W�˹�"�+ "O�L�SL�`2`�M�T�2�c7"O���B��$ԁLP���b�"O� ř%T�������Y�"O2%�"�^q�\fㄉ���bd"Op�B��%v3|Q�t��4y�Q��'$���+6�HH#�8E�m9
�'E�$ʴ��=#�����G����'��Q�ą�?m��0�ۗ>�0���'(Ш�5G�N��,���ރ7��@�'N`�:!pH��U��|����'alp*%	s�)R�,:"I:�'��t��оa����#D�z��-C�'��ܺr��'[w�T�E����
�'��(�C�C�Te
�%�[6ke�	�'���cT'ԀI*�YR�nC�1?DX��'�|y�a�YO\��Q�_��^�z	�'�`Y:b-!3�<�P�+.b� 	�'%l8ل O<+=��{����*�LS	�'[j=�@�U��rph3�ŋ6�P	�'ބX*.�u���:v�I�'	T��� V+���b*Y�����'
f��Çe���JJ�`9
�'딤���4{=�I�%�[�<��q�'�~Q������mYj-$m0�'�Y���Y!!���k� Xqp�y�'I����H!�0�EO�=jg��j�'�(��� �)�X��o	.p0�'pѰ���R�\)�Tl }�Yq�{��.$�,������'/����Nɴ�������2qA�J�{���8l�E��[2� ��m܍O`dB�I2ވ�Y�7JR�x�D�/�B�IV2���Ъ߄]�.}�M�33�B䉤P�X�c���E�9���/�~B�I�jǸ�3Vy��CfI�#y`$C䉾,���ɋA[���h��cJC�)� NQ�.�n!9�B>^>���"O�J�C�5E�x�*�#X�p+09��"O��٣�Q�I� �͝R�TU!�"OС�4�7����A����"O&��kҀv�4�!r`]�!�$M�e"O�䢁
�"w�|�䆖' �J1zE"OL5#�HɊ4�L��SƄ��0��B"O"<aQ�U�rt��&�$t���;�"O�<���T�H�s�/Y���E��"O�Њ�/ݾ�b�@���ض"O��J�c�`Dɳ@�Ǆ�4Yy�"ON�8PmֵYD���"�g�=� "O�D�Dٛ#��89�C� ��(�"Ol�,���B#�81kZ�"O���G��g�~��`_":���Q�"O��Q��ft	��'үV9�0�"O�jJ�F����%g	�4���u"O^��"(͸0`�E���� C�"O,�x�aσ`py�떷C�VQ�E"O��e*�f��z���1Ѳ�&"O�i��/ÇD���� Q�>T*R"OHl�P �c!j ���z�r�"O ���.�
��Ɋc�nq~P�'"O�P5ʭH���K ��$Z�����"O�LH�*ڡn��ps⚑�h+"OJ��P�EbU
��]2��9�䞴�yBC� *2D�DF�j��A�X�y���dk!�Q�
f��@�[!�y�ϱB<�P@�Z�h� N�+�yRK�{@ ��K�&%0���y�p��E�>��+D)�/*��Ĳ�'�L�32d{��c���7�L,��'$��&D�/fY"�-d�B3���yr�R �P�
�g�6�M��n
�yB���_�5��B��,�@��3�y��3F���Dݑw��S5Iֽ�y��
i��|�!�@/��d�dĆ��yR��40iʵ��F��Q�`4�yrf	l"��(1�]>6mDɧ�y���/o�T1�,�3)OP8��Fş�y�h�i�p����
�h ��Ա�y��Yo"�yj���&)#�y�'ɕ3g��[��I7�tL3�M��yRd��b�:@R%�$�hq)��yBN�5 �(�*��2a�HYw.�'�ybEM�FD��xפ�T�4d#�d�)�y⯀�p$�6l�Gj�T��	�yR�ԍI%jT�!�؛vʀ#��Q�y����Z�C����D�zd!Fm��yb��n^4hW�ECW�L�FGJz�<���	�(Q���NL=Ei\%�KUB�<���9K�%H"߼fw0�X� H@�<I�˞�B�<��ID�3��<����Q�<	u��^m�X��_�OE�`SBj�<I�̏�4jj� �D9�N��1+o�<ɵ�ƨYh��R�8#/�Ð�i�<V�	D��3 � �@��<����g�<!�HQ�t�d$Y���LFh6d�<I�ꀴX�@(n�I�1X��+5b�c�<A�� �:e앪�ޭ	L����y�<)D&
0����?8?�)�B�_�<�!�A��)b4U6`qe��W�<)���%�F�Wڵ	v���B�p `B�!�����B]�B�)� t�P�@����x���̶*���W"O0��#�R� �*i��I��}2iJ�"O����c�0�T@C�\+R�t"O�X�©�5 K�]Q�a��O�V�B"OҀ+3 7s~`(
�-K~�Qp"O*����Y,l�ZG	�-"D��"O����Έ�A}���D-�::\�s�"O���+�h�b��lJ�q:�"O�ĸp+L#5�nN�\I�G&D�((����7��	)L�� ��kT&1D��{���&-y�,�'1j�,R`�;D�t�!G��zm��kA�k�̸Zh&D� �'"���պEn�04�XL;�$D��2�N$	Ut��Uc�� �>���!D�*�˘'+�=��D�412$�dG/D�:����&߱dt�H�Oe]�B�I�d?�ث�� �`Ț�bI�kZ�C�ɴ
���CB0��Y��WC�I O���"�
~��Qd�U-t�C�	�?�*�f�%mvt�s���-k�C�	3&w�Ĳ��7kEN�ɖF�u��C�	�w�6�k���* U.�"Q_�f�~C�q�%� �Ѷ�̣��ǅq��B䉘����@�0'��k� E�h�~C䉛S�bT�H����\PqH�k�4C�	6VrH�#��!Y�8{3�a2$C�	�Ox���F���z���m@�j� C�	9{��:g��D�� -��C�I�d��B�g�#�nY�`�Y�(-C�I�i=Jᱣ�&9PQi�JǗ���J�B���I�9+��)�)U~�M�QI�Z�!���A��>K��8�g��\t�<Ĝs6��4��<�@j)���G&��~�R,K�*�Z���PC�'�u�5�V A 隵�M�s�T}*�dK��hB�I�#E��3g��BĦȡC��Z�D#=�!�ұb����Rb"�1�J������r=�f�����p�"O�q*@)X�|0bI��̞�tQ�Z�"�B���+��:L�XKm��"~��H���t�ڐYa2��L�K�B�IR 
x���ŕn��2��ƇI�E#�4qֹ�vɝ�&t��4!��|F|r�^3���I���8���U�5�0>@DԈ"�s���k��)�iX6RZ��i'�Q�O��%���˺���Ą#���H�&!�¨����41B�O���"N�)Y��ە����S5�~�@�G'f,����<<�@���Wj�<���hL��jа(�T�񏀏a�`��ɔ
,	��Z�Y�D��;Or���<L�\��cC:�&�p�"O����[��m�%��C`Y�f�ަa3d#H�:�!v \KZL�݈�O�,�nV�sy��@lP�ތ���'��h�ȋ19�[ �7}��SW�Y�ZKJȊ�^�8�0|ѳ�A5e�����A��(��3�y8�w�ON����$Vt:S���4�z���i�,t2,KL�-��t9!��5A�a�]j��gg/�^Q`!8Q��d�	K�<�&�l:�'Br�d+F#$�R�#XD����\�F]!��C�4D&����)B��U��#0><5n�_��"A�I�*^�y �wݥ#��$ޙoh.y[�È�Z��U)�'ʈ}��{�aL�2����3#ι/�
h���;L��3t&ȉfe�(�t�P�v[����Ԙh��,�d\���Ij�U�3�i��Q��&*̴�{�n��� �~b�������"�=���B�`�d�<�&,����g˽fd��&Ϳ�~r�|��4!g���MG��'P���R,K�[�12@��$N��b�'�`�+���Dx^�k&AM6 9@��<yE��$I�6��5��bf�	BMJ��P.(�2`��끑�p?yd섹&��)Bt2L0Ѕ ]3%|� `�q"C�	�$W���댎U�|�+L[F#>���Z�B�~�ӵ�J`�'���J���nء��@�<E����S�? |�KqŒ�{��RTX$%����OD���ć�z@"�O�>(F��j���¨ƙY7H03�<D���5�����F�8P�	��j<�
1 8���ɚ*�Ɖ	�1�X��2�dU��,բ\C'�P'1�j�Y�Z���o[��i珉7 ����& &�؄ȓ>=�5�vː�zd���ܛIDzԄ�a�F������s��סkR(�7"O�������K#�D��k�� U�XY�"O���m��IҨ��S(�+aq��"O��;��ؗ�>�X�OhL"�3t"O�	S1˖6�R,3��e��T��"O�����8�hP�R�H�+}���"O�!�	=Q�r��#^,rP$`#"O�����W.Lx��3R0%X�<b�"O�U�v(��I���O'u@�	u"OB=�q ��tస�Q�<e��p�"O��%+�x8��b�����"O��"�d4\A��㥇�
���"O�l4m�#K#L��B�;u���C"O��A��O�6Y�u�K�G�T{f"O��A� ۝$W�����E�s�b��c"Oz�0D�\�zw<!щ'˄�I�"O8��%E˓Lv� ��#M2��y"ONAS��ˤ�.@��ͷ&��@F"Oؑ���C2X|�2Ph#mo��:F"O���G�N�B�3���b��k""O���ԍS�Lb���ŃXI<yhT"O�(#/��$���Q �A�C
�"O�dB�-@$X��తҹw�n�b�"O*Z5%]&�hRb���庁"O�(p&
ǟ/}"�zt��j8V=��"O���%U��2�FH� H��a�"OFp*#J�N��$EV3r�j!t"O�+@�L.1��)�C�ɍ�~j�"O(� �[�6 �:�QZ�t��"O.D���R7&�TH�%�@QnT�"O mCL�M�q�A�9J���1"O�]��O��Næ�
�C����81"O�<�2��x��;v��2r����"Oȝ�1kӹ}�����l��l<,�"O�@pe��5�<��0,���F��"O� e��[�6��,�T�R1ۤ"O�`��֓窠;�$��3�ZXC"O4 ���I-S���kQ;9p�0�"O2���B�J�qj�a4tq��"O��;#d�
��6�۾\�ˇ�y�C�Ty��p&iIJ�~���L#�yCG��ЉV!7G�j���"�y��R$Y�h� 5��N��HX��6�y� ����i�L��H�L��y2e�?~ �Wg֬i��;�eû�y�M@ p~H��B͒�Qbf� �y�
�r!2��/��˵��y2�ȶ(��Y�p,��	�r���H��yb��.�:���)�(o�����yr�ܠ"�"���H�0�
�*����y�%�d��ܠ�Q���q�V����y2�J1>Z����,a�)y�"	��y���!wZ���C�
 �
��Ѹ�yo�+P�)���.�h
$��θ'M���7X+ށ�EHQ85���YM>aT��k�$倐��i�re�Is�<�ǃ�e^A��I�H�֕
U Rl�<yq�˭4D��(�2ct
*�'�d�<� ��ɴl�(����M�n�T`��"Or=��i'���(��N>�&Xw"ON��F�јFH23�iGJ�@�"O2<X1�2� 4��o�"�К�"O�q����p��H6�?8<L�W"O@ݨf������	�):��!"OĹ#rJN-�� �( �mj"ժ�"Op�0��ɈS����R��+/���"O��E`Z�C�6���-@�-����"Ov��&ƓXϢ��LZ8�T(qt"OU	��A'����A���Z�PQ"O���
Q�a}̸s�޹ �j- �"OL�h�'�L-D����=�c"O��;�ʠk���q��X��l��"O��kf8ܜ�R���!K�i�"O���Se]�(�(r$��:1f|���"O*�2�I N���$��
d�<"O���'�I j��4BXtb�x"�"O��x�(Or�dA���	V�>�r"O���`�
6f(��kY�o�e�s"O��ؗ'Y[�y 7M��p���"O��s�M>(ޡ UM�f(%��"O�)S��.�f���	dZ$��r"O�q�� �(��8����f��"O6�� ��:���3*��6p�#"O��U�]Z�E�ǆF�6� cU"O^53vd��_�lt��K؀7{@1X"O�u�V�)\�r���Rv�&"OfC��݆`�<AI� 9se(�sd"O�l	B+	&��|y@�ϗ2a0i[p"O��ч�֜W��y[qM� V<\��"O���7K*�fe��m܃CN���C"O恀���<76=)�N�g�n��@"O����/Uns����K��.�� ��"O.���'�{B�dA�%8ٌ� �"ON��g�k|pp��WC�"�0�"OF��d��1$� $�T�dHa"O��TgH�aQ�mᕋ�4n5�u"O$��nZd	�y�d쎵e��d�"OPx:�Ǐ@����勞�$�,��"O����n�n��`��r\�U"OX�aԠ��T���W�Y07���E"O��Ѵa�2R����"h�Chd0y�"O�;TT�J��dqHE5fTJ��"O�����e��iR���AE����"O���p��C�T( ���w*()�"O��Q�c[8U��B���78h�Ic"OB5ٖOA���Ro�?a����d"O���Ȁ�U�bTJ��E9,�Z)�"O�j��T'�$ۤ'�4f^�H�"O�yrqo�
S7�Q�#u��a�"O��0��	n�̄H���7HI��"Oi��JEpr"�jUBEz2@��"O�����R����E���˧�[�<yS��6h�r�͸	�#b[�<)""	�[�Dt��m�+��a�$.A�<��m¡� I�P��-�:䫰D�T�<�pjͶ c$�S �ީc�<i��R�<ACnĝ1�]���P?����`K�<��R�E(� hq�E?6,�Q��L�<��
V�u��0��<Kuf$�U�2T���� =6��h��)	��؉�6D��9 �	�:M{b(0V�H��g6D��s�=�ݛ�E�`�`�!'D�� zE�#�R.sՐ�I��N�"��"O�{b� )� 1`��g�h�u"O*,cf���o~l�3�/x� i;�"O�h0V�n͈��nC���Dj"O(E�����0��G�ۘ\ZeH�"OD�Ц�@=E�r��jS���my`"OhDB��Ո,RB�xb�C8f�P��"O�5K�.�\b�)��nԠ*�` 0"On20��A4�#N
�X���Q�"OB�3�\�q���ʤ暟6�H�*%"O��8��ǋ7�y�˒-mu�5�"O&L*WZ:4�q��ꔠG��y�"O:��B�q�Ġ`�L�(T3�I�1"O�(��V�2�q*wl�p��	�t"O��jb�)�Q�b���9���"D�h��E�iV8y��҉>+&sc$D� 0��\2�)C���{S�YW+%D����
y!r�I��Ȩ6��R@�6D��	��ֆgm 9"��4�a���/D�t�,&x��Cl���XJ�B�I5
���Q�C��C�����f�9V�C�	=�L��b�G�Xx件c0s�$B�	�}"5p�QDbD�P#�[g�B�Ɂ
�*�;��30�-q���8�B��?ZA��16��=|-H'�*alzB�I�,�:8�m�A\q�R�ߵp^�C��S��U�w%X����!&^/��C�	2m����'@�$��ց�+�^B�	�p���i4B��$Š�@Э@g~B�	VR`H�	��8�ɉ*�vB�I	-Q�x��&W>b�&�2rcܜ�,C�I9]�dU��5D�N!���T�:C�$1f������SF	1C�Q�*C䉁R��ٶ�� ���W�:R��B�ɔav�bv�S�J�
]{u
ΡZ��B�ɴh�PБ`�e�@T-� j�� "O 3�o� Cn�&UH(ؤ"Oh�H��wB5j��ڣ6�3!"OH��_�/!�ɛ�( �.)��"ON�+u���$�<1!�Ύ T$�4#"O�Q�1ěՀ�j��W���!"O؈CKL�uB>�#%�e40�!"O�U3�-��+u` �nW-����u"Ot5y7)�4DM�I��P���	@"OfH��MJx�y84��:~):�ȃ"Oh�V����O-I�|U���LY�<Ib � _�`��1bŴ���Q�<��
a�J	ZP� If���OXx�<irI_ L_R Cg
�_�0���Dr�<�qjԁ�$�r2d�Bd�@1El�c�<`n�]�����Z�i�r���,�u�<i  ͒}'��ҧKN�I��C���m�<��Ԩ�����˓6eB��t��C��D{�*S+H�0��+ԒΕE���\�C䉴F��H 7�L.������(l��C�ɣ�����[�gܚ�kQ$��V�C�ɅV�1+��{C4��F �H1�B��5l�f��Q
M"wL�)�0�_{��B���ؽX%��o~tIdE��]�B��
M3Da������2�?3�JB�	���	&�3f-���Z�B�ɢt`�Y;�h�-)D�+�H$;GC�I"s%�����(��(�0|��C�ɖӒ��tְ)RX|���ǝv�C�)� `���
#�P�f���T�^)�p"O�}�aؾj�0I��t�0��"O���ț8Z_� $Q�W>�q "O0(��J e��䣠і�Ⱐ�"O��V�A^�re��#�)4"O
��'��]P�y�m�:�2���"O�4띞}���(G�o��b"O��ٓ,ܘ-jv5�A�(k�T�"O���N2���KN
1R�Ԉc"O�� H�b�V�*��g;�9"1"O������	E�t��l��b	cG"O���W������K*9��a "Oę���Gqk��Ӗ`ɛM+���"O����!�%T�� ��#
`]��"O��P�F@`~�0��֞U�p"O\�!TdVP�j�N�!B� �r"OF\� �U.)_ʵ�@���4�*lY0"O��37�μ%Fh4���O�:[�\�ȓTԶ�0A�X�M`2ՊS˄k3N���L��@�aU@�|��ۦY5� ��y8B(�q�Y�\񓠅�C9>�ȓzP���̖&X�z��	[pa��aH�5�Ĝr2�Y��<>�8�ȓb"2ʰ��i,R\	��ϓ|?��ȓ (����,Obth��̩��W�S�Y�ka�`ơ�5����ȓK�|�2��;|L�K�m0b<0��I�dĢr�2S�$��T3%|t���H��Y��Ό�s
��cC[)Y��������I�l���E� u�Nɇȓ�|H��b�'�ͩӪ�|u��ȓn�\��U��a:�	)*@}�XͅȓH�^-���	2��x:�A�*���ȓ\6��� #\6��LJU%Ӥ���7��"�B�"z��·O@,-ɸԆ�T�؀0Љ���E��愩c��M��xiҜ���9Md����Q�|��ȓ`ݘ`����QI<�r* �{3�M��o��9����u?zH*b��(u�ȓK���y���o�6�y�`ڶ_a�ȓ��ѩ���0�T��2���4u2�ȓ#}����K��<��Q���$i���h�h��\�6�"��b�P�7J9��s�}�v%����x�#�;�P��S\�c���<��Y U�G�H��5�ȓ��i�R��,`������lV
!�ȓɨ�X�@B+B�`��Ӂɵ$Ь0�ȓv@͡"iV�qy�w鋧[t�ȓ#�<1ƥۊ���bO̟ L �ȓiu�Q�ej�ΘC�_$V�zY��U�,j�O9n�@󤢕���A��nFX1��f�<X�9�@�MD�����TBÁE�v��i�'��<,�ȓ.�(8�@�4M�hfŇw�
��ȓUȕ�2&��P8���Ϯ�"O�Q�w����)x$��S�U6"O��&Ó�_v�����_��ِ"OX�:�m >��Sr��/��=�#"O,������f�q�oߠ�摳1"Oj�cr��e*"���HC(�%x�"O ��H�?|�y�'��]i"O���N� r(D���,�n �"O@�Z���bմi���G��0���"O|LKF)��f�����a� @'"O� ��33�Н��VC��y[&y�"O��s'MN,1Ρ���:A����"O`�`\�l�J��(%��z�"OL�����:},=)�F"7�@�"Ȏ��n�]����%�˷h���"O�pbv_&�����	���T��"O:X�S��(g�H�qv�T<��@"O*UY�ᕊG�ĉ�&�[�f�N���"O4�C��|�H�
�*a�6�&"O�����?G��yb�D&�x$�3"O��R�2��y�VjS$?Ȥ�ۣ"O�����X���prϟ�A�\��$"O���lJ�<,,i5�âg���[d"O�030G]un\y�.g�h�9�"O���r�Ȯm�`H�!K)x�B�0 "Op=��˦|�̈ˁ���{��m�F"O���	O�Yr6��8kr�q�"O�]�T�20�m�ׇ�2[4N�*�"O���p
�%T�dI�#!�"�Ah1"O�,
VIπ,����`�.#�l�"O-��%ՉO�X]J���ڡ�s"O��QVG4:��X���~T��`"O��[���.s�1z��ؾ��"O�Q��mA|�:p.��tъ��"O.`�ƄƋ�qS�Ӡk.��c�"O���@��\�P4�_�3&� �&"O��i��+��<�di-L]��"OH�;�(�=NM�Ǘ % [�"Ob�ر"�7��a���O	.�9�"Ov�!"�E'y2
�z愔�a�S�"O�(pI���ٲ"��%hH6x'"O&Q&kN�TF��1���af���"Oh)Rs'�Q^���E���HL`�"Ol1:P@��8���`��KJ�C"O�hS��^�M�����t��0�"O,!�T4Dp]Y&+H+uքe0�"O"�k��#�d����[0 ��8�"O�-��cF,$*Y�R����F"O�}a��
=8*D�.��;��0"O��{���
-.�2q��\��"Ov�B�Õ�FV��'E�*1�����"Ol�B������%�6	i�@�"O�	!�N�3;�0`��$�_���"Oȱ�.��1(�Qi��04"O04����J̽��N,Xò=*C"O±��M��
�X���4����""O��ړ͞7Kd��O�$�����"O�y�SOW*t�xE"0�V�� 5��"O*�'�S���m^�p��c�m���y�P�w��#��n�&�0��6�y�C\��̐a7b8R��b��˝�yR���x�i`�;O�n��rC�'�y� N7$&Iy��X�@����VJ���y��E�\���Ɯ*���1�]��yBҗ��T�t�į �i�(��PyRBO�]Di5fQ�z��<Z�\@�<iVE�`9�E9���5D׀1
R�z�<�c~��1�kל'M$l3��u�<��%]&�	�����KQJ9D�TQ��3��  �Ǘb�a��.8D�̈%JI��MbV ��G'ځ�6
5D��2
\=5�������J*��:C(/D�Q��]�`��f�3Z,^�$3D�\Y��)U~Q�]�&� �3%�<D�� �M�������b	�i�(�q "Ot)
5�h%H�!�8p��ct"Oi���(Jv	Sᗥ.�,���"O��0L��N�s0 ^�i.X���"O���'fB:fK$@��(׃#1B"O �8c!\hH��Q��%Ib��"O�����L,�}I�ѐ{�&�H�"OD����O�����O�x�Re8"O��y�GP�`wJ݉�̴g��l�"O�Ũ��.ql�G�~�K���y�g �1����e�%��aH>�yZ�d��D�2<@�3B*���NU:�'8z	�U-ձ	SL(
B&��M�y8�'K�*��E./�u(4-�(K/J@�'
�3��!#F�����I�����'�| P�����#�1���*�'�@��q&�7	�8�`ۀw�@q�'m5��G������E]�tJ@�
�'��Y�!�6L��R�#�7=h4�`	�'� X�@ǦJ��\���%R^8��'+�0����#ɚ���
ʈEI�'xj�;P���fQ��@�K.S�'�h��F+I�l�H,�t@^�_��d��'�f��A&\�9l���a��U��y��'�,���DK,VBt�G�y��e��'�<P`

��6�բR�.�$"O��]���� ��]�JΦlk�"O q��͓P߄��Ӧ\^���"O[��R�=�F<suC��Q���"O考V�ۣA�1؅"R�5���B�"O"�̃�7nh�����c�����"O�u�␄\��i�
J5���r"O
xǉ�b#H��'�Qr"Z�{�"O�Q��26K�?DjnE�`o$�y�jL�<hv����$7\T� �)�y��F�aİX6�˾!s�<�7@�y��G�PǨ�X��V�����֬���y"�P�n9$%�M�~X:�����ybh
}�=��e�g��\i�,�*�y��B���2���s<�U�v���y�>dM��(Ze��Lȳmۖ�y�a�74ʌ��
�t�*�$�yΈkkn��3`lB��2�Ȕ�y��>J���r(\��`08M/�y��K�{h�
����7�@� ���yR�#��Q�C?)�@My��=�y"�:$K�0���ɷD��V���ȓF��E�0�R�Q����gkJ�[��\�������O�3+R�Q�Ң>���ȓ,ϒ���˱f�-�����(��8�ȓ~�����/n<|a��22�Ʉ�i���l	�K����D�e�1��0��c\�&��1@�ܟ\X���P9Ʃ۾mnIi�Q6�x�ȓ)	d�P��95@4�i4F�+��Y��,:�-Q�c�@�^�'�S��ȓ7-��kv��$[j��n�=u����ȓ)R�,�%O�xdc��X�]<���ȓ-�^!;u.�۬���
R�@!��/&�*
�|a�A1$��4pT��ȓ/�B�b%�T�4}\$���h�⽇�B��AаOI3/i����%�� ���r�Q�j�3KY��x���
a�2 ���4-��8:4�X ���af2D�� ����ņs�"Aٶ. �m�� "O��ۡAׯ]�`���"�=!e"O�-��@�?E�\ �M�^Ҝ��"O���פ��:X�uF8I�0yi3"O����0&AbWg�6�p�R�"O� ��c��j�}���a��1�"OX�RC��PH��W�B	�R"OJ�ʐ���k<� ���
 ,,S�"O�I2��%s��R'��@��y�w"O
��Tk�y�r"�۾I�؜�"O��W�	:r�*�B�V��&"OK�N2mc�� ���
D��yr�@�ɨw��$M�k	� �y��72l�CiM�mqX�9����y���f�T�J����V��k��y̘�D�����$<�ʭC���y�J�jR()�����@�UJ�4�y��G� �#�$���	�y��í$�.���4|�H�$���y�䓨J��5�nɥ&>�! �I���y�FS
!�*q����!��mi��©�y��L&
��Q�I"i<H�H��yRO��P�4�Ҏ;Q��ݳ7��$�y�!��E>D���9I������ �y�R�"!�TIR%+IlJT!Ǯ�0�y�F��t����� WkD�2v���yr�Q.��IS�H<fDJ��.�y��!%Cr�؅u�r�ig���y2�X��L�7H� �s�#�'�yR�P�׀[~ChRPgJ��y�\Yc������{:ޔ�gˀ��yrP8X����EXrI(��wA�	�yBc_�����رq�r��Ǭ�/�y	G uz��J��T�J�C7(P�y�/P���0����H��j����y\E��2�/�:F��x�!����y�O?�TY�ؖ;�E��mR��y�B��\;xQ����Gm65�`� �y���jB��hs팙VAtk�A[�y����|�XR�c��˗d��y���E,�X���D5U��Rw�N��y2G_(![d\���#JL�x�����y�A>�F���.�J���0�yR�ЏD���	Rm�G0�qw�'�yR�O� ��m�B��B�8?.��
�'�a���fIe�G���J���	�'����aa�w �iQ��I�
�I�'������T�����{S.��'z� 6H��@��l����F�,���'�>��Y5<b�ȗ΁,x�TQ�;D���v	ۊK�h0Y�K4[���B	:D��Q�A-c�����im�ˇB7D����Ʊt���雺NH�1AI"D�p�`B"1Φ�CD�Z^pzV�!D�����D聢��
,`�S	!D��HA� �)Y�Ԑ���
<ҡM)D��r�D����ئ�+7,qZbh%D��i���9��R� $�$����'D�dY�`�W�S���:w[��J�"'D�$I˔��U��	.���8D���PB�^bR�"dZ� v���p5D��S!��p���v&ؒY����62D�:���>\"���dU#U<�D��1D�0�T�PɴlN�a|���4�<��B�)� v�gI�
\JQ�����y�6Y�S"Opib��\cv`:tΕb��;"O]{��М�M�cH�|�u"O�!	�	�k�4��"`�|��8 �"O�|bg��v��5�EC'9���R��IԟDQ�攊���'��Y?�*��Q�R\(�&�ܝ$^\0S�OS�e�TH��?A��]��=K`��m|��	%!R &0����~>�b��'h���F�~�<�І#.�=��I"l)���a�$~��bB N$� ,��%Z�h3�,+e�}^�� �k2B�T��O@oڳ�M+����	��8��� �h�?+"d��Z�eX���IF�S��?I�W�j�@u��g�BݛtCP��,�	�M;׸i�����9��ɪ��W?l�H\)鐓�~�'Y�e�����'F�Z>E� ʟ�I�����l˽,l�%.�2l�j���䝏s�nX2�Ƃ�d��a�%�8 )yT��?ŖO�d��|�!(ó�v=�o�� < Կis��1�f���+1F=�0�W�]Ss�U�Q�z�����#Ԫ?~X~a����.Kb�	1�i�Xu��՛�jrӂ�d?��qfN�?� �0�)�?���be㨟��	AX�@�e�T"!Y(�s'!
.mH���/3ʓ ܛ��xӀ�O���vݽj�ϛ�� D��A&Mx��ϫ�?1��l�VU�����	�t�I�0r��J7MǶ:��9��4+�����\���`Q5|�m`��D�+n6���G��?�) �/F
��iF)C,[|Az��:�0��W恅f�6@�U�]&%ܳ�~�Vڶ
��=i��<I���h��M��
���IFIS�4}除
���z������ʟ�'�V����h�V�R�f�%6x0;�'/0pD�K `k�"*��������[�4����������lpT�.̈́�1��6
����i֝K����O6�d�O�%SN�O�D�O����T �Fu#+�/`j�����>��0��֙,�HP�����ZKH�����ЕQ؎�(D�T�o$4��ѫ��a]���'|�pfd�")�8yh��j�@a`C�Z߸'�4�1��M� ��Is0qC�0žu�s��bjO��$Ʌ�����|��m�^ۖmc�l�K8(��I	I�<�pMJ���p�#�Ӂe \P!��G?�b�iS&7��<�3�$~�v�'T�Y?��疊���&I�g��X��d��RO������?q��p�p�L,��<�%��e��KT�l>��DG2V6}(���p��)>�a�X�3�%ݰ=����7��	�U����#peP<+��X�2�K�BqA5��35$�a2�{���?)��Q�O,�vL<$��df�P/:�2�d����5�)*�}Z0�q���o{|�Q���83����H����}�N6T�%�j�����3\$���fƮ~���Ÿ}d��n�ڟ���L���P:Ig��'i�fe�n�8�&I�=V�`k���xV��GěW�&h���6\r5�$BĊ��4[>q�����L=E�D�ٚe�&��ExR��9s�L��P�W;�\"G!��*T�3�i�� }��{�ODU���)��E�`�@=iՎ�ʦ�`���O��lZ%�M[������F� }��p��	$]Ό�aBK��~��'R�'\��P�~���*+�]3��$v�
=(�,F�'1���f�B�O��'0�ChL,
��ՙ����×|��'��ј� ��   z   Ĵ���	��Z�JwIJ(ʜ�cd�<��k٥���qe�H�4��S66<���]�f��->(p��o�!9�0��o��gZ7mæ�‫��y���<�a�	M���$a6v|�,/ff��K��J�➨�U�xr ��4�f`�`�i}����!p5�q"�
�8�|B�O&�!q䆨?vt�-O^]ڗg�]��(Oԅ
�IN�����$	�o�Y��Nш4鴰i`��9�<Op��mR�m����|�"��+?��!ywn1D`���)�5OqN�:�L��1 s�ނ"�~�2�O�l�'"��Agc�>�`�%d������@��6����A���&\dx�oИ��DP�X�D�8A]��3�\��Qn�{rt�r�Y.(]S!Ɯ=v��G"�I�D�$hf�X�H���.ڊb�d�BB	 �O�)����ն���	�g��P�g�"n�vI[�$�:?�:�b"<�Dg$�����8p�1�0)>�6���O����$���j����r.����JN� 劶�d��OF�y�Od�r��A3 Z12�� �e3�T�|k5�ɳoR�O�𙥪؂5�P'����Ѐ[�-�ODd�����?�m@Ȋ�B)��H�d��q�~��#<9�/.�$��O��`�������1�ߧa���Od�N<�c_���!�H@��hk5��-9��y7�O��Y��i�J�EG0�?A�CQ?ͧ�~rq���R�H�ؽXTh�u5��gJt�E�d#<��/}B`Q4)��1�s�!A�4 �΁;��d^�Ot�s���	�?e
M�'��,j�\ٻP��K!�d�? �  ��u�r!ʯUi\q�9/��$�O���Oa:���O��$�O^Acc�r��i�a_�T�ԕagJ�)p���Bgo�uZe*� C��s4m��C�Q��/�e¹+wa�:���
�� R^���݉k��#Ӥ���
��#%�9�MɅ� c�9���^�
 f�,�ȸP6�ɪH5���հ�M����$ӼR����]�|��fƇt���Y��ٽo5 E2f�`�'aayR�N�r>�c���f�T�T�ܪ4e����6Iܘ�lɟ!��r�`L��u��'�"�S���;bR��U΅�f���	0%\u(����'�2�'BX�����O�MۦɅ�v�<$�!Bk���@/#�T�s�F9E1|@���@�h�<i��J63��i�r�1sT���&�v��|s!	�< ul�h��,2�֕�B�әM��+Sg���L�1����MC�i��V?i Q0S��ِ�±!�\���e����DY��?��$�"z�x��r�t��Lk O�H8����4_盦�i��$� ��@L+^%c.T8�U��sQ���M+��?�+���8PI�Or�dӖ5(c�A5+m�x�mӒu�a��e�t�В��P5ߦ�P�֭^~�Q��A�R�O��Ա����CE�(��Ȼp����T�iM��GCP�Yo�u�a�.�Ms$!�p|� oL6|w����A�V����C� ^+p"�Aґ�˦��c�O��o���M�������L�:�fU��M��V���b�D��~�'��mX�p���+@�9C �����01��/��M+Ӹi��'��S-��q8��F"_
5��HAT$�����?��P�*~�@���?9���?ه����r�|�k�Ny�����=��X���$%�,�q�j�YJ�[���u�|��S�P�F�іg)�� ����U�c3�P!�H�����C -��1�'#C��X  �ºc|��$.�@s�C0���z�Ƭ��%Ҵe�LA��5*�'������?1�x��'<"U�DJ�G�j-�1ѳA��y@�!R鵟|�Iܟ�'��}*�*Ǳ)?Xj$�|��A�ժ��7�ɦ	%���?��'�8i1a*Ʊ�`�Z�BG�$HX�s�H.;,Y���'l��'[Bϛ���'�d���bu�b���n��1*�W�H~B=�A��2.T����bں}#��X8,���dZ1\�!h�l����S��I�='����K�7-��nZ�2_H4�p �2������#�@�OŢ��'�D��A�.��i�w}\ܓ����>)�7��Or˓�?!��?������������^�{Ș�ygi���yr,-A��k��^n���Ǝ��~"eC)A��7�<Q�N"������O�B���ɒI�U����P)�)s���d�Oz�$؝=��TO3&�	�B��Ri�S���D��0��EH)�D��a�Ș=�t;��#H�t���D!=��	�rCƘ4Ul�+ԉ�g&H��O��R���>�b�`B�8l$��j�@�O�alZ��MS����i�:e-��8��Q�vl�$�bSdˆ]Sߴ��'��#}��Z�٪1�U>>��Lar�1����d���ߴ�M;5���6��&�_�;�~�
�Jq�'��' �O"i��  �   d   Ĵ���	��Z�tI�/ʜ�cd�<��k٥���qe�H�4M��\70<����z@�v*ɾE P4%�M�R]M�Q� �6��Ϧy۴8��$ �Ibybl� \�!����V��XS%�,8@ɲ0�PK9�=a�#?t�7M�dn8,��W*¹
�c�.2���&�ʠ�"��RG�I�Us �j3͔;���<2Jڽ��%W� 9�P&�92���Ej�6*;�v�tTx��/0�H5�V%�?)�'�������%g� $�r���9F�(�fbSA}��{��c˧~f���'�(� >0�kÁ��<�cH�y�p�I֍�I���C�+UC?�� )�Ƹ��Dy�+�	�0����Xg7�	�q:\	j��W�8����J�6��#�ߢi�~�@���δ�O�y��?l�ڠ�ጔ\^8E˳��X�'���Dx��A}���	���ɲ G=r�`��+����ɱz��;��$�/��*�:Fu12�V�+��j�K�'�@�Exbb�2G@�`�+cx���13�� �}��LT�'�pd�'�ر�BD�]Y��H�!� Qhh�k(O�d������'/�� 7�,h5R���#@�u�N<�-�t�'��Fx��˟L@c�ýV���6���@ܙ��/>�I���쉂�xr���%�6�J@�=7"�-�~B��}�'�i%����'��U[���CK8eS�էRub����v�I4���	��iݩ��rD����y+pm���1-Ƹ��%S���'�\%FxҎST���n��N�(Sb�!H�AB�P8�Iv=�x�1�I>H�fak���0����)26ۘB�I?t� �  �7j<C���Ci8,|�)h�E&}r{�'.��=1UI�jR�IJ�!v�V�"2��ʦ݊�ቮ[N�dхĉ� �����I4]q��P��8
$b�TS�I�j��I�5�A� ��܅0�cL�*��� |�#<�`0�	�O�TaAFS���bK�#���t�Ɉ`�X��'�bh	w�N�[�:}X�G��>(ybHJW�'��&�t1�f՗,�<�1�� <dXm�������	(S'�'�����h��OB l,����b���xy��Z@?!�l]?��	��� \w��H�A�
h��'i w�)����;�O���H��b#��KF���Q�6�tD͢>�� �4�"<���5D�ThF�H�_2���A�<)@�� 2  ����C���q�.D�l�#�    �	       m!  �'  .  >3   Ĵ���	����Zv)���P���>��'���qe���OT|#�j�9]ֈ���
�*U��r"O1�4ŋ�/^LPi���0HEfIqJ�O_�����+�\#��i�,IP4�4>z�Qv��:\m6�1�I�Sg�-e��4MD`ri�i�rA���o�B���I�^p8���O�f�Q櫁�d��k�}�"�Xu��s���*_V0d�2#ښ!=���$�89�]ەNL&M^q�&GD���	��	ßభ�:������q�de�1a�v���l\y�)ߍO��q�2�'ˆV:)4��a%t(ՙ�oR.�:m�QE\[08q�ۜ���'F�Ƞ� 	Z���"�����Z���񖂍�)Ŗo�ğ8�A�ڟйܴ)��<����~��W�1���IhV4�vM"�ɳ�y�O�qmV� iT'ޜ�2� �M��qsV���FyL�O�}(W�+C3��C���`;��yռ�����?����?�`��`�d�O��%�z8�[��>Ղԣ�0�� �i�-M����S�߶x=�b����O��k�Fd�|�{!��TB h�@��0k�-;%���@�B Go�bs�3b�jz1h!��B3b��-A$C�6b_� Þ�%�Z6m�æ���yR�')�O��W/X\���It��P�� Y�0B�	�3I��	f�m��)զ؁��(��	zy"���B��7��OB�d�?���/ם^<�4�� >����r�}�6!	��O|�d�Oj�f��P���!mK�w�l�m��F�:%�I�@��:tP�X2�m�'��x�Ah�`t��2/� T~����I`Ս]9N���)	BTH̥ ��	�s��D�OJ�o�꟨��$ �Q+��9s"��p�n� �v����9�i>uGyF?)���r�]1/���
q��M���?y�ʟ�x�'5�p�D�Ɋ�R�bĨ�Y�pYg(�>A�	J9B����'��'��D+G:Yb�'t�� �C�cQ��S�L��-��mj��)a���O���?A/��O2��`��n2x���ؗn��y���'�"4yed�-{�Z��E�ѝ=��?��S,ڕ1#�9���7P����ȅ�H3��OZqo9��T>�Ss�t勳[:��SQ�T�,�����ww����I؟H�}�qjSu��J�r��)3��W��?QZ� �'S�> ������8/:�@����<:-�Ȓڴ�?)�?4p[�����?i���?q��}u�n�O@�F�T�MRRp:s��2L��Ѓ�ڈ^�����3�&���F-�`	��(OD�ٷAԭSv����X2x��`Ps��J|��%XsP��d+	�6�3�]Ĥ�wȌtC� s��~�t�'i�y��?����'�	׫x���q䫎 F܂�����l[!�Ē�tYP �3�Da�hPGm�+7Q�f�4��|���������a�	%Y��`���=D���Rcɒq����O����O�����?����į��DN�ĺ'o�-/��\�����~�P��6�׍Yv���@�Oqxȣ��(�yцh�S��T�y�u%�iK41���D�O� ɤJ۞l"�T��]�p��`"���Od��%�)g�%±fUL�bZ��Ʀ�G{��ɅS\�8q��:zA慹'��m��C�Ix��ztB%/��B�s������'��3��p��J�D�?�Zŀ�F��P���� [�XHvCo�B���H�O��d�ON���	��hI�A�A-h�ԟ�R@C@=_�����A��S�ؙA�ɕZ��`qS-��'4���d��� B��Bi�
���<@�Ņ�hO�=�@�'n�6M�@�'="�	p��'h�9g�ھ0����'�R�'��%ӵ�>R ��+�It���
�Dm�ɟlS&a��iD�k���i�eϥp�j�lc�\B"G�;���V�G�	Ӱ�GzB���=ת�K5B���HjaE*�y��U�֝��A�|-�Tۅד�yBRb9S�B%&��vgͦ�yr#ψ`:���wH@�T�Е�yR�'�	�n�P��)�(��y�b�#�L1v	T">+�e˵ᒱ�y���B)IGa�h4B��	�y"/(5�bh
��O�C�K4E��y2FZ{FhKB([�;��� �"�y"Ƙ�V�B���fP`�H��Tb@�yrI�0�ޕ�JݘNF¨xdh���y"��<B�E��b		^�T ��]"�yb�D<%쾕I�m�:���MC
�Py��8j"�z�F�-*�`��u�<���c�����0b�n�8�]N�<�Ь	$���:�a�&s�h�j�F�<� ��j�H切�0�6Y`�ďC�<ɤo��w5��0�ߵ/Ң𳤘_�<Y�*���9J�À�x�`��B\@�<� �\0#�/dhlh �>SgE��-�3p��C$�Ζ&b��2w�i?>#|J]�<�$�V1��%��L�@�X4
��1D�
rI�14H R���k#$yӮ�2�f�)� ��ɆP-$*�	�]�H�Ђ#Z�̹�"a�qm,�����J�\d��ၨ���cGΎ� ��P ��\)J���x�-�lh�� U؟P�󃅯3�y�Mۼ5�m���3�ɬ?"m���5��;Q��'�47��d�L*Q���ABG(a  UŧJ�y�AE�Q�&��T�]%#�@y�D�BG\�tWi
�o�\T1t���M���?�sS���?Q��O\m�.A'����cYv%��'�v$��Ŷa�l� �7V"U�΂�L�� !�i  �ĮK�j�RYQ�M���Q���H '��%��&�;m����Ì�O�Q�����X gh�$��.�+M�j�	�Ǆ�o�s�
��Ri��0P�X�2�
S-X��@Y+�BS@؟��" ���с�ޟmW���Ic�@��(�~������B#y��i�	L8
@r��W���s���o�� n�p7*[L.�Uq�a D��@�
ߡF�@�h�"��=��<����pkFܸv�2y��f�����O$@�j�*��}-�=��O��Z�)P
Q�&q�6|����'��HP��9���7_��s�ütL�	���ɾ68 xr�����J�`��z��j��7��Onh�@Y�@wP�l\�O8=��$ՇBrK��@J2��
�� ��|+��0,w�����1��BnC�@�S�4>���-(�O(L�#�!@.�=����+�@�����2 �U�':���g�H�PP�"�Oc�ܔz�����6m�Q�4��& "!�'�R7-��:5++D�0@u���������w"#t�@C6��/X�Pm���������x��&t�4u�3B�>�ǅ_1-� ��ȷr���2�]\8�0���� 6��p�SdȽO�~��@dD�g���z ��*)��� �G�/��zĮ��'����o�]�'+F�q֫إz@�1[�B�}R���d?'=�\�l
�5�tpY�#�^k��pT���Î0�Q�J+gC\�h�MPkU��Y3� �O��v-\��#�BRa�<O���q�^q�n�"�(�`�L�t=|�h!�]�S�X�*q[t,Q�Tk�I�4x>B�Ix���׫Oz\t�>`�3"����׫N�hA�Y	pc�S�ft��.i��1*�O���P��M�f��q
B
�4ب��')4٪�M^�N%R�`�\^"ؑH3O2g뾽��*ͺAVJ��'���p$r���+(�R�F~� ��n�L����1H�@uUhЄ�HO&MQ��\�?�w��cຈ+6l�$%Ltj�F�ސ�ʝ"G[PL�wA��vX�t���'�V�J ���iɒ��w"��{W�� cU�D�|X���'gȸu��!�ִK"ğ�I����t��w`�`Ĭ�W���Ö�u M��'�:D�c��
k
��rvDCC�K\F Y����1J9��(ݴH(��� 0+��2D-�����T�H�G�]�q��](�a�.��!��'�O�q{�9�$�mywF��� � "tR`�V�w��6��8����"��tSb�^�W�J`���dSZ̩�e�]?*M䘒�Lӷ/#�h��mԆ^4�Q���G(y-I�p��rDL����#!�d֎z��,�� &T�~4F
�7�V'�%�`�|���i��a���v���
tdU5&��y��'�8�afO݉~]�p�o��\�2r�O��1�/|O\u�ELI�#3��r���)�0��"O���e@�c�@�W�`��"O挻�&M)C�8�!ᇟ<)U�ā"O�,�ǂº6���� �%d���y"��nP��m��.z��������yr�B�d��Q���+!��aѡ쑓�yB`��L�L���,L�e}z%	���yRd��H�ѩ�,<�`����y��_W�X��ƀח���eCG:Y�!�M�[x� gΈ)5W*Җ�@�H�!�d�xLʑ����Lg�@[��� [�!�D�>@�Qp#�U�d��*��!��8��H��V ���f���{�!�$�<��q N�_��A�L�v�!��S%o�S�G��0� *�hS��!��e{
D���Z�S���BC/�!��2t����Vl�m�J���қ6!��L=�T�E!�f��@'� r"!�䔌9�ȴau(Snڠ���T�A!�ǚ<V�P��ˎ.fL���'R#Mh!����\�U��)QM�x�u��G]!�� j�8eX�*9�l�p��$#V.��&"OV�$J�$YU�<�q��4y�P�"O��7��aN���X�j�c0"O��bg�0�p��l?#պ���"O��e`��y�F\+eͮb6vy3S"O�	s�d��ԉ?+"d��"Oz�����]�u�%k�7���آ"O Tb��E�t�`r6*ע	�>��"O�eC�ɒ�z�r�Jw��'REA�"O����&�'y�@K�HԡW&B��"O�q:�mЇI��%P"�Ëf& ���"O%��f
�!�H���>'
)�"O8�ъ=��`DKJ;E�q�"OV :���a���'�}��"O�u:≚6�ލɅ�p�(� 6"OR���_�rqCFћ'Ot@@""O���VjTw����n�
 A���"O��c�� n($|��\�BxQ]6��O*�}�>d�,�UGI�Rx�m1�J�{��t�ȓ{ �Zp,Z��i�Ui�]hL(�EG����'�Ja��f&�Q���[4CA�ד3����@����VANb�l�J[�)�"�%�B�I�#��Q�C
J����*���O�����
Zy�u9Fd�J�O���� o
Ta"�2dEr�	�'�Eâ�#I(�9�鏁\Ӣ0S�BAp��<��j�O��1%���� �D"��T�Ln2�;��߇/�����P�;�J)� �O�P7:����L U н����KR��	q�'�{�²�O���a�p�@�����U��D*�[��Աf���b�C]�2�m���[�y?�B�I9(3�!y����g<b< �-؝Q|�Ox�zD&K�{���(mdo<9F�dg����Rf�H*%�B�0�:�y�.�tg��*Z� �qĉ��mBqHsnQ� ��a�?h��L~�y&�����3F���HY�pR%L��?! .��B���a�@��Y�@�9�.Ep��Y]F> ��J� ��w�'��,u��0��|z�Iul2�b��$ĽB��݀��=�԰ˠ��~�B��CcK����T�ވ���Y1=)L��� 8&� ��yS���h�:
V9�'��L[�R�j(9Z��	pIs�t��WcLI��"��Jt��3�D<��O�
�
���x�����l����� ���`����"jӐl�F+�?��~8�'X�� 7�P�+?�`�	�4���M؀��A;mQ���'�Q�W�,eu��yo��-O9�Dz�B�g�y"�N�p����êb��•L'��Oz��3c[�O+�|�w��r��נ�/a�T�r@�v	R��4��.�TB�ɄlM�1卑����ـ|
�9���a+
�A������ |&�0D��@�h�l�2�uۘM����/�y�$�J�@����:h���S�A�a�P�JX���)���|�<�0��<T�H�ɰ[P:Y��OW�<�D#C^,��Tj��J�����ȃ֦�a`��%4J��P��v���k���AvfM�daI)lOέ§��l�`!�Ӽi�(��q�I�`mjAhe��W�T z�'��-�$A߃_ �A &�e[�{�A��,��f	�h���G@�Z0��H?��u"O���Br�q!�S�dp�d��o8��"�xr�<�g}��ەk���Q�L�c��H�rݮ�y��S�a�.x³�D=3�D����:4B�|{N��d�=yd	�ŎV�V)­q%�-o;�{�*�:Q��I
�)� 62Q�h�4�C�	�;����Ŋ�܁��լ?�$C䉯#�H��ea.	��Hsa�<S/$C�I�- ��7�F�vw�䐶��,i�B�	3��d�Ɔ:K�T���T$)�B�I�6Jvɑ��Iw�d��7|�B�IX�>�B�1@p�3���Ii�B�ɤjD�(�g�:T'&�ޜ.�B�)� �q�s�QO"Ց��^�7 �p�"O`�Bc�U	rʈ�ABg��Qe6i1�"O�s�(�N<ԡF(׶!���+p"O�*�`�	.�����(J>�Bݳ�"O�m�Q��%T� �&� ?�(��"O�\1��%Lx����b38�lR"O�]�f���l��#LU�*M�P"OLē��}#�܀`L\HܺB"O><B�Bч����!@�+kB0!"O�pC�C�,�4�ɑ/�'�<�r%"O�L�b�Q�$� A1daP�R���"Op�0C��M����(3���"O�l��Q�eI��2eG���0"O�*Ó,9!���c�;_B©�p"O �"��43���D'�z����"O:��5�E�j�ti���ӑ$�zh��"O�
��T�Y�|�Rs^M�.�:�"Oʰ�G���ږ��8j� P9�"Ol�0��F�.e���	��qP�"Oq`�FRo�<i6)�?��y�6"Ob��3I�������;����LW�q �[|z  �1O��܆ȓ7�� !'Q#M*�Hu�^
#�I��G3��tn�%"���sSf��1�<�ȓF��i��g�~Ũ��{���ȓ�ެ���Ů2i>�KV�ٚń�]:���-a�x��`DV�pp�� h�h�A�-6��#�h@�S�]���A�U9�rY�7�("��ȓ4�>=I�kI"�dx4	+xǶd��D �أ3�G)y6 0@PO�I����cf���!蓉,�ΐ	s�׭``L���h�8���W�:��R#�^�R�؆ȓn�hؐ��o �Ś�EM�dl�(�ȓ}  �P6C�?���&��#
�6a��ӢP&ݣGR:�iҦV�^� �ȓ?���0�G[�/�����z�숆ȓ<p���5eH:/w�Ys�̉� ��ĆȓC�\H$�0#�r}���/����ȓ�F��aFE�OP��ecʲ3)�@�ȓFo0!�WmFm�x�2L4E~5��wz���#O��0 .[�{�܅�sUB�b�T}"�GJ(2
��g���c`�U�LsƝ�	�N�t���9L�dI��wU
�P���	;�2�ȓ
K�����z������� ���tz�)�%[�W�>E�En�_�Q�ȓ[9��eM��rH v�Ƨ;����ZU@x��dy~-�%�	GHN��'�X���l�<Q��8Cp��
`�tb��ě6=�,EH"�@�(06��aDP�!�Ĕ+ZV��ĭQ�b��Т��Ԛ_}!�	�M�:��$���!����L�e!�$�>����'�I�RQz殈�U%!�DQ� �	�0Jn��y�-ն!�N=�8���6����uk�(N�!��Դ��i8F,֞%��ꃠ�y�!�D�d`)�'�O�$!B\�P�!�A�2�4ړ�	�|1�4��W3!��ƛL�>�tK�&6�*xB*ė%G!�Ċb�8���S�tySW��&-!��*�BQ��/B�qۥ��(!���ՠ��!�Mcr�!�p���4!�ٻ^Y���L�4d�0,V�g�!�L�pLh&J
ZQ������P�!�� �(s�.B蠕��a�lT�!"O�Di!BR�0w��hB➂sT0�1"O*5�F�ژB!VHӔ�F�|fnMb "O��	����@<hs�W LW��J�"On𒖯��hԖ{4aT�s��PV"O�,��cV7
�+�J�<x�<��"OV���. �pp��j@j.+\T��6"O�8F�j��0+!#�8	�& �&"OB���^h�\�â�HV"O��XC$�7�eyE� x���ib"O���ID*@�n��bͧj���"O�����	��� ��D��qI�"O\��a�!il�Y���=�:���"O��2TMJ�|3n�h��ݨ��g"O���G��k��-�ciZ%��tK�"O��C2�ڗqa��)WSʐ��"O4��"�u�f�V�Ѡ)�vӒ"O�`� �c�2��)UXwDɣU"O��ȑ��G����Ygr�#a"O�\�C���Z�� H @|��.�!�DRt?bM#aJ,1��Lx��M�!�$�
t�<K"�S5f�9�FE�?�!�DU�~��r���+8�� ���#=2!��<1�n�P�ŶP�c�E4_7!�D������Z'����!\�!���J��a�fLJ|�>�1U���!�D��f>(�&�� ���q�!���pH�"#���#ӿyO�ȓ%E�`��oJ�����\�[����@���
�lG�g�q[�-W�`z�E�ȓ �Ax�%�Bb};ƧU94_>��ȓnM��jC�2,�ITG�~Zhl�ȓM{�=�PӉ<2���S�1v�ȓl'Xh�U��_�z��ӌ�D�и��J�呥D>b.h;��W=T��̅ȓi̍���I�$�4c�ʷ�B剭9HK	; 2<��M&�Z�f"O"�/�L�Ul x��'@�l�C�Ɂt_8C�l'^زa!1O«FٚC�ɉP��Ѩ��u�!*���f/JC�	98�U{�mU�x�n9rg�+�C��2H�Đ����:V9��%ч��B�I>W(t����f�$��f� �B�	�d�.0��1?^i��
�K4B�	\�^4��)[*e�J!R��(;�C�IV�Bǀ-i3>���NEY�B�nj�A�ʻ#\�x"� �TC䉅iT��%�<� ��r��yNC��\Qn�{�K:E��\����N�B�Ɂ �����\�0�|�g�^�u޸B�	�>�*�h+'�`�B�_�^��B�ɹ��9��h�>f�P�b%k\�&��C�I1<��e���Z�Ia�rE		�HB��,j��uZ��^�?�Ԣ�"�eFB�I5?cD��)U!"*�<�9�nB�I8tJ��ʖ�U�C�T�җe��
�BB�ɗ,�(��E;l.􂄂�j�B�	�^`��!���L��B,?T�C�I"l�bA��m�����QBD�]��C䉱�6�����V#�ZcK]k��B�ɌrZ�P8�@���u�$��|B�		'���i�L��e�`9�vi�(��C�	�w#)�P�:հV	Ç^KB�(��f\r���$�.��C�)� �<�'��!8��9ňA5��#f"OF��pC��4G�M:���f�Y�4"O���P��5|Pܩ�AP�s�� �"OdP�#�Q;Sr$ŨS-WR�@#�"OD�C�����[#��X��mK�"O0�5DF7�Z�r��	�(�����"O~�`"��1L���˧Z9�D��"O@L�F$�61F�Шg�-#<P�b"OV��Q�3����속Q"��'"O��9���SX� !.Z����"O�='��Xe �̋<~h8e"O�E1�)�*f�IR)��~V�D�"O�Z@�\�sx<���fB��s�"O��A��6*��qg��8e9�PXd"O��&��q���1W.Ʊ4z�`�"OfdXC��x<I��=gr���"O���֬ў3��H�2g�W�D�"O��[��+�JU�0'�8E�P� "O�m�RJ�h�!�Խin�j�"O�x:E�:;��sV�ޕk�]��"Ol��ѿn7�@z$��.s���"O&��b��Y�%�T�A�@M*�b"O4�v(Խ#��(�d��?�e"OZ4:�#7!��2-Lip�"O�� �Q$f��T�_�/,F�0��'��'�t�Hg�LP��}�E+L�9~}��'g�}��d�'���	��ʉ�f]��'�l\��L�aZX�QC����	�'��Q�Iy��Kb�Յ;�=#	�'��=(���)����!�_�GJ��'T�͛�dR7W$�<�D�W�;H�'������?C(	��b� ^#���'�H��ѨA��eP��& ~U`�'
����K�x��QMނh���*
�'��=��΋J��F��n����	�'���jց�#S�EaU��t���$��%�OXq:��N vY���E� \����P"O�t���Œ_��h��=F��"O������NHl8+qC��tL^4��"OT�K��G3g�����U�d�F"Oz���]?�P�r��(a�m���	�HO�6p>�H�`�7F8�|�çM%?#�B�I0LQ��JGeS�d��JB.��I��6�%�S��M��AK�a�t�[U�Z�)�����N�<�c�M��Ie�ĩ�"���	K?�F�'��|8��H*N1!�1��9	�'kx0��K>,(�!p�ń-à��ʓ+��� A�9���1f[�QLP��ȓl�"xq��(M$d�P��C�B��X�ȓmw�!`��"���5��5=�,ԆȓE��x�% ���$x��*�-�&��ȓM����$�U��hk7@6	�h�ȓc��=�cH�-Xt$Hm(�ȓ\�`�P�M��pċ�Ӿ��l��/\>�s�0M����e�ws� ��%��1��]�İ��
P)9:Έ�ȓ`�V=:b!�w�Tm:ǐ!nC@���y+j��0⏂z=�8jX�0��5�ȓ�>\�7���&�i�Ɲ�t�@\�ȓ9��B�n�P72����	*��݅���m*'E��2��@S �,�Ԥ��a'6E1wG�=1�E����(\F���74��3�K�1(� }j�F�"J��ȓo����AV|W�Z�d�U52\��S�? �!ʂ�̉;��,SwaA Aj.q�"O(y
��Dg����v	�!5"O�H��Ԭd�iq�"Q��a0"O�=�L!q��`���P�$�0���"O���DV���H`�����;�"O|�!UcZL;ƌ�%#ݝa���"O81kEV:�x�AtAˤ=�x�"�"O�!e�ϝX�$*4�_�f�&�1�"OJ��5苖)�x,9`-�"x��QJ�"O2�b�HC���F �#h����"O���3h۸H���R�J�>R<xv"Op�sq�>J�Z|	��Q#9Q�И@"O>1�J6!�M�4g�K3T�K�"O��(%A�0+�Z�����||ʅ"O씪��T+ M�9r��q�,
�"O��0��^�h#�F�!��"OZY+�Z�	>4Q&�O�a"��"OhAW+P�b�М2iT4e����t"O��d��%2��R���r�	�"OU�҉8!;|qIWgS����"Ol\�g/�"r���+sd�	0Q�"O^�٣b]3~�=!�C�LV��d"Oz,��O�d_&x�(��bKz1�"Ob��rj�8�%D��+�"Oz��4ჍP��A�᪃.,�6��%"ONĂ���k4���O
y�6d�r"Ox���ⓝT���#_=��!��"O6t(2��\萕��	�+!�~��"O��r�)4���i��ޑ_)��2"Orm���KB�U�Q��	B�A��"O����-#�j�z�@�"?2({e"OE!E)�*%�ȍ�յxZE��"O����#4�X32�Ěv]�ɉG"O(b�нJ�rt�r�&O6�*U"O�:�@�U�`���L�=d�T@�"O�܁��Y**�����N3�Ĩ�"O��s%�#������0(Z��D"O<��b+G�VEb���}p�m��"O��K!BJ��$xR��C�E�0"O�Q$�]-Mz����� #�8q �"O�	'H�bL�r�P�n�j�"Ov%h��-�-��o:��6�3D��3!K�3.�^��t��B���d�3D��:ևM�(I8R�ɺa�� ��=D���4�݀��U��+}��h�!:D��
`C\�A�1����=CSg7D�DI�Ւ�م�}�ʹR��0D�p�� A/~�R]A��;_��5�0�*D�p�bj ���y�e�D�y��8��$'D��"�d�;����#GΦ�ʣ($D�@zVM�eR�t3@4u�u� A"D�T Ԃ�)^~t��K�8�Ni5�2D�H���;u���1�
�*=xC�F%D��   �   j   Ĵ���	��Z�tI�.ʜ�cd�<��k٥���qe�H�4M��\70<i���:G�&�����0E�5��y��cA�6-Ħ�q�4x��$"�	}yr��2�p�Y`f�lٖ�&�H�܋'왭e�a�=��,)�=`6�ĺ)Π9Q�$�x��)xׯ;w<�ɋI�q�ǩ�{���(�8YvN �q�	 ��U	"�$q�Pa�� �`����[$��͔9,�%�	�Q��`�d�?q��'�0�%ڱ��E�*ߓU���p/�EdUI��A�����d	*3�i��! @9OT��U.
e,�ɏ]�����b�&�FŉrP�G����d�����Au���t�nY�t�P(H����OF�����BTƕ+u�ҸuG=kՀY�[H�a"@\�Ƹ'0�Gxrk7�YP"F�]�CF�p�p��	�*���a�Z��h�����ڔ�290�x;�6}B&V�'C�X�=�SDZ��`�W�\&0��bb���b�ቮ^���%dV����!�c�(��Z	L�Bc����A(��NFM8�%=o��*E�)v� �'�B"<�d!���2,<��-F�+U�"���*>"4(ቻ��s'�'즥���Gb:}���HW|I��y��y�'�~�'�xa�ժ�r�ϼ@�(@T� <�~���k�'��M$��s�'���Be�1]�X$��*�/F���C�+h�ɄU��	��i�M��Kp�dņ�I�ɠfQ���s�O���'��Fx�
b�DN� n<�2�� C6��d,�I�@��`���I��0���E�W)��a���	dQlC��5>�� �  �&4D��ic�OZ&�g�{K���"�3D��2�g�*�~|���'�Xyw�.D�|Hb�	;_��dy3c��W�@��4,D���n�����[	T�9`���ybO�5V�y L�1&��;T+�(�y�B�2�`�F�_�.H� �#�y� C7)��q'�\�(ke���y�l´uB�5I����X�H�HMJ�y�MZ�E%R�RþP���¦R��J�'������=�\I"�iĞ���Y�'�|�T�K&��I�Q�� ���Z
�'�N�E� �� [�@�H��)	�'��C��W�l,��瑄\�����'U�5A���o�C�F]�i�8py
�'j"��`��%:p(Yǋކw��$��'H:)��ω?��j6���i�4��'ðĠ��M�F�Q�Ի�    �	     (  �!  �'  .  W3   Ĵ���	����Zv)���P���>��'���qe���OT|#�j�9]ֈ���
�*U��r"O1�4ŋ�/^LPi���0HEfIqJ�O_�����+�\#��i�,IP4�4>z�Qv��:\m6�1�I�Sg�-e��4MD`ri�i�rA���o�B���I�^p8���O�f�Q櫁�d��k�}�"�Xu��s���*_V0d�2#ښ!=���$�89�]ەNL&M^q�&GD���	��	ßభ�:������q�de�1a�v���l\y�)ߍO��q�2�'ˆV:)4��a%t(ՙ�oR.�:m�QE\[08q�ۜ���'F�Ƞ� 	Z���"�����Z���񖂍�)Ŗo�ğ8�A�ڟйܴ)��<����~��W�1���IhV4�vM"�ɳ�y�O�qmV� iT'ޜ�2� �M��qsV���FyL�O�}(W�+C3��C���`;��yռ�����?����?�`��`�d�O��%�z8�[��>Ղԣ�0�� �i�-M����S�߶x=�b����O��k�Fd�|�{!��TB h�@��0k�-;%���@�B Go�bs�3b�jz1h!��B3b��-A$C�6b_� Þ�%�Z6m�æ���yR�')�O��W/X\���It��P�� Y�0B�	�3I��	f�m��)զ؁��(��	zy"���B��7��OB�d�?���/ם^<�4�� >����r�}�6!	��O|�d�Oj�f��P���!mK�w�l�m��F�:%�I�@��:tP�X2�m�'��x�Ah�`t��2/� T~����I`Ս]9N���)	BTH̥ ��	�s��D�OJ�o�꟨��$ �Q+��9s"��p�n� �v����9�i>uGyF?)���r�]1/���
q��M���?y�ʟ�x�'5�p�D�Ɋ�R�bĨ�Y�pYg(�>A�	J9B����'��'��D+G:Yb�'t�� �C�cQ��S�L��-��mj��)a���O���?A/��O2��`��n2x���ؗn��y���'�"4yed�-{�Z��E�ѝ=��?��S,ڕ1#�9���7P����ȅ�H3��OZqo9��T>�Ss�t勳[:��SQ�T�,�����ww����I؟H�}�qjSu��J�r��)3��W��?QZ� �'S�> ������8/:�@����<:-�Ȓڴ�?)�?4p[�����?i���?q��}u�n�O@�F�T�MRRp:s��2L��Ѓ�ڈ^�����3�&���F-�`	��(OD�ٷAԭSv����X2x��`Ps��J|��%XsP��d+	�6�3�]Ĥ�wȌtC� s��~�t�'i�y��?����'�	׫x���q䫎 F܂�����l[!�Ē�tYP �3�Da�hPGm�+7Q�f�4��|���������a�	%Y��`���=D���Rcɒq����O����O�����?����į��DN�ĺ'o�-/��\�����~�P��6�׍Yv���@�Oqxȣ��(�yцh�S��T�y�u%�iK41���D�O� ɤJ۞l"�T��]�p��`"���Od��%�)g�%±fUL�bZ��Ʀ�G{��ɅS\�8q��:zA慹'��m��C�Ix��ztB%/��B�s������'��3��p��J�D�?�Zŀ�F��P���� [�XHvCo�B���H�O��d�ON���	��hI�A�A-h�ԟ�R@C@=_�����A��S�ؙA�ɕZ��`qS-��'4���d��� B��Bi�
���<@�Ņ�hO�=�@�'n�6M�@�'="�	p��'h�9g�ھ0����'�R�'��%ӵ�>R ��+�It���
�Dm�ɟlS&a��iD�k���i�eϥp�j�lc�\B"G�;���V�G�	Ӱ�GzB���=ת�K5B���HjaE*�y��U�֝��A�|-�Tۅד�yBRb9S�B%&��vgͦ�yr#ψ`:���wH@�T�Е�yR�'�	�n�P��)�(��y�b�#�L1v	T">+�e˵ᒱ�y���B)IGa�h4B��	�y"/(5�bh
��O�C�K4E��y2FZ{FhKB([�;��� �"�y"Ƙ�V�B���fP`�H��Tb@�yrI�0�ޕ�JݘNF¨xdh���y"��<B�E��b		^�T ��]"�yb�D<%쾕I�m�:���MC
�Py��8j"�z�F�-*�`��u�<���c�����0b�n�8�]N�<�Ь	$���:�a�&s�h�j�F�<� ��j�H切�0�6Y`�ďC�<ɤo��w5��0�ߵ/Ң𳤘_�<Y�*���9J�À�x�`��B\@�<� �\0#�/dhlh �>SgE��-�3p��C$�Ζ&b��2w�i?>#|J]�<�$�V1��%��L�@�X4
��1D�
rI�14H R���k#$yӮ�2�f�)� ��ɆP-$*�	�]�H�Ђ#Z�̹�"a�qm,�����J�\d��ၨ���cGΎ� ��P ��\)J���x�-�lh�� U؟P�󃅯3�y�Mۼ5�m���3�ɬ?"m���5��;Q��'�47��d�L*Q���ABG(a  UŧJ�y�AE�Q�&��T�]%#�@y�D�BG\�tWi
�o�\T1t���M���?�sS���?Q��O\m�.A'����cYv%��'�v$��Ŷa�l� �7V"U�΂�L�� !�i  �ĮK�j�RYQ�M���Q���H '��%��&�;m����Ì�O�Q�����X gh�$��.�+M�j�	�Ǆ�o�s�
��Ri��0P�X�2�
S-X��@Y+�BS@؟��" ���с�ޟmW���Ic�@��(�~������B#y��i�	L8
@r��W���s���o�� n�p7*[L.�Uq�a D��@�
ߡF�@�h�"��=��<����pkFܸv�2y��f�����O$@�j�*��}-�=��O��Z�)P
Q�&q�6|����'��HP��9���7_��s�ütL�	���ɾ68 xr�����J�`��z��j��7��Onh�@Y�@wP�l\�O8=��$ՇBrK��@J2��
�� ��|+��0,w�����1��BnC�@�S�4>���-(�O(L�#�!@.�=����+�@�����2 �U�':���g�H�PP�"�Oc�ܔz�����6m�Q�4��& "!�'�R7-��:5++D�0@u���������w"#t�@C6��/X�Pm���������x��&t�4u�3B�>�ǅ_1-� ��ȷr���2�]\8�0���� 6��p�SdȽO�~��@dD�g���z ��*)��� �G�/��zĮ��'����o�]�'+F�q֫إz@�1[�B�}R���d?'=�\�l
�5�tpY�#�^k��pT���Î0�Q�J+gC\�h�MPkU��Y3� �O��v-\��#�BRa�<O���q�^q�n�"�(�`�L�t=|�h!�]�S�X�*q[t,Q�Tk�I�4x>B�Ix���׫Oz\t�>`�3"����׫N�hA�Y	pc�S�ft��.i��1*�O���P��M�f��q
B
�4ب��')4٪�M^�N%R�`�\^"ؑH3O2g뾽��*ͺAVJ��'���p$r���+(�R�F~� ��n�L����1H�@uUhЄ�HO&MQ��\�?�w��cຈ+6l�$%Ltj�F�ސ�ʝ"G[PL�wA��vX�t���'�V�J ���iɒ��w"��{W�� cU�D�|X���'gȸu��!�ִK"ğ�I����t��w`�`Ĭ�W���Ö�u M��'�:D�c��
k
��rvDCC�K\F Y����1J9��(ݴH(��� 0+��2D-�����T�H�G�]�q��](�a�.��!��'�O�q{�9�$�mywF��� � "tR`�V�w��6��8����"��tSb�^�W�J`���dSZ̩�e�]?*M䘒�Lӷ/#�h��mԆ^4�Q���G(y-I�p��rDL����#!�d֎z��,�� &T�~4F
�7�V'�%�`�|���i��a���v���
tdU5&��y��'�8�afO݉~]�p�o��\�2r�O��1�/|O\u�ELI�#3��r���)�0��"O���e@�c�@�W�`��"O挻�&M)C�8�!ᇟ<)U�ā"O�,�ǂº6���� �%d���y"��nP��m��.z��������yr�B�d��Q���+!��aѡ쑓�yB`��L�L���,L�e}z%	���yRd��H�ѩ�,<�`����y��_W�X��ƀח���eCG:Y�!�M�[x� gΈ)5W*Җ�@�H�!�d�xLʑ����Lg�@[��� [�!�D�>@�Qp#�U�d��*��!��8��H��V ���f���{�!�$�<��q N�_��A�L�v�!��S%o�S�G��0� *�hS��!��e{
D���Z�S���BC/�!��2t����Vl�m�J���қ6!��L=�T�E!�f��@'� r"!�䔌9�ȴau(Snڠ���T�A!�ǚ<V�P��ˎ.fL���'R#Mh!����\�U��)QM�x�u��G]!�� j�8eX�*9�l�p��$#V.��&"OV�$J�$YU�<�q��4y�P�"O��7��aN���X�j�c0"O��bg�0�p��l?#պ���"O��e`��y�F\+eͮb6vy3S"O�	s�d��ԉ?+"d��"Oz�����]�u�%k�7���آ"O Tb��E�t�`r6*ע	�>��"O�eC�ɒ�z�r�Jw��'REA�"O����&�'y�@K�HԡW&B��"O�q:�mЇI��%P"�Ëf& ���"O%��f
�!�H���>'
)�"O8�ъ=��`DKJ;E�q�"OV :���a���'�}��"O�u:≚6�ލɅ�p�(� 6"OR���_�rqCFћ'Ot@@"��.H�$���J#s�Yi4�G�uaN�25M�@�!�$��pD��Q���N/��z4
�J9	Cl�|�	�
�Q>�4���",S90�F� sAN�hͅ�Ax�H�Z�j�v-F�o������DH�dcԥH���&�U��\5���B$'�H����>\O�)��Y�"���'�Hh��VW�	)��&`�$��'�����j�x7�E���Ex��+N�$��e$D�]�S45WT�G��q�p=0CdP��� _�y�g�������mI�k~�x��닝�F�h��Z��$��=��;��L>၎�ͮ@��+�26r~�`�Da<ᅆ�6���8"'� {�1�dpԴ���c�r��o1ɶ��������G B��<)&��J�ax�-M� ��@�Y�pi�T@�o�'��4����D-��{I*Pj�'�քsaI�f�6�E��r)�V�<ic�0�:}"�
"kօqiY�����KjZ5 *�
#JԵ�PQ�v"O�9&"���i��#�tmV �w�α#����%���{<�MB�n0<��O�1O���f�=Qy�$�,����!�'r����|{���v,
+c�����9�q³/��,G��0"*1����D�Y��ؤq:� ���Y�k�џx��j�0������'�`�2J��kǀ��+��zA�M	rGX�pϦ�
�'�2*R�W���ݲ %ִg�Tm�,O2 s��S��P�m��L�U����Of���CӔ��C�-Y�k� �'��0��H������ĉ-s�<u�� :䰛5�_˦9�aƋ�n��OT��O"�)gÂ�C���ڐ�To�YS��'�"�+cˍ�J���Y0E�6i�:b�
K5�	�@b_�E�i�%�����D�,,���&�� TI �&PџX�sdD+,dQ�&
@A�A�&��b�ltX��}�xyC@�E9x����b}�Q��JV	h�S$	�8,:���',Ѫ�@�1�t͑C�j1�Q����
LH�Pg M'>�f �/��(�!��N�q�&�*�c\�Q�M�b�<+p��g�b���1/�T?����y�-����};#��t�I�#@Ƹ�y��ő;w�|I�.�)3��[����M;v�^�o�֤:aN�p=� ƄOO��PA�:FҨ�Ӧ_]؞�zG�X:U����7I|��)E�I�r�8�ض��u�dE;"OR�"R&<��	2&́Z7p c��P�[��3�j1F�>�	@$�3$�TڧME(�,da�l1D����	N�3�@.�<�\sB!ºX�8�1�Rd���^�*���F&�8�xI�q�Z��!��Y�#Ü��D�Q���"�GR:�:6ę������	�3�,���O=�%���Mz:���JJ���_�v|{F�Êr��T9�CCbp��O�P��p���S��e�e�٫l:�����╂D�-XU~ز�a��`�ȓy?�DSFܖZ�Z�*X�p���N�$�[�&ژ ,���)��q��@� �U��?0�x| �㏡^��!�ȓ�bE�k��LQ0g��*���ȓr��0�GB&58�¬��%��S�? cT'�J��X�'C��E#"OR�j�CY&rp|�6����B� �"O���RmK�L�\����'M9�8z�"Obء%`�}��ga��pQ�"O�����09���!swu�"O�yy���JЈ�;D*L=	L�w"O�A���o%�H��+߅l(ԣ�"OJi���m�hd�>�}S�"O4���I�(�DL8�O�.Фݳ@"O8h��N]�0$�16`��|�PU"O|�Ā 7"�iKD�Ć+�Ny�'"O� ��<Y��}aqc�+L�⭩�"O�BǠ�h��1Z��ˈY$:�i1"O}��%�Պt� �,}f�YB"Obe��1\�,)�l��n�⨰"O��jg�R�IZ%���8�f��"O�٨�E Ȝ}y��zR���"O(�@�6b�д���pR�y"O�i�j�X|bF`ե@�0�y@"O`�&��/P&��SM��(m*A��"O�ERí��N��p�0f��N^����"Oڡ���6���'��7d�q"OA�'JI�ڌ��Z�<+<�y�"O�0j���I�vP��,t�,p�"OpZ�%��SW9!�_�JdVyA�"OpYFG�7jhN�j��		8~��B�"O��&FY�,<�qY5��53���0�"O�t�ġ��H̬U:t�W(�r	+�"O L�jA1s�ţa�(�΍��"OV�؅!\�HN08�CQ����V"O�Ăs��r��2 	���891"On����2;� y��K�>[��g"O(	B�K!a�fi���#j�Tx0"O2 J&l���֐�DO7yc`��"O�|���,X'�TX��+.���"O��S&��k�6��0ߝq(�� "Opx���V"'jM��O}"����"O2Ac����#l�P�֥}���8�"O4L����A�b��6a 8�*���"O0`C�U~�]2 ��4���""O��S�蜉&�J��4	ɷa�V�e"OZDH��E�3SިC�*�t� I(�"O�A�pE��w�&�b$I�3����"O���ݾG:��[�iF"z�n�xT"O� ��A�F���� �Fq��"O���F:��Tա8_��!"OR$���ťx����d�:���"O��a��d���z ����1�"O|�1FP�_b�zģG�g`�9�U��[��3>}R<A�ő~j�!�.�Ph��������Y#n(�D�ȓ.��&ۍR�����_+�)�ȓy�� �Wi
dmy�l��A�p�ȓr����Z�GA��Xb�û!ÊՆȓ>u��H�B5=���p�\�;N���0�Mb����[n�P�L�8B�N ��5�бQ@m��c��eAR�¬�ȓ:�F i��[�r���ڒ ӿQ��`�ȓ;jHiB �\>S��pRfl_�@�z8��vR`��W:��ꦪ�11��9��j� !d#P꽙��ԫ��Ԇ�OyP]���B�U\l)x�ʋ�7�t��ȓcN�Ae'#h�Xͣ�ߝ7��X��U�<8��ĸ1�б�琴5����ȓ^=��g��:>vUIv:):���S�? �y0�l�
l\}��d�����"O�$��#�_�D�X� ��o��C "O���d�>A�4��L���Ⴃ"O��X��Ȓ����MWy��I�"O��c`BF�/�6�C�,N�B��(7"Of�[(��\�����T3�ă�"O�01�J�����S���"Oq@�51�sAL��+x��"O�Ȓ!qi������O�֐�p"OV�B��#dr���Q<[���A�"O���Ӌ*o��Z��A-Ra�h0"O����K^�s@���?'w#A"O��IڣD5"踖BR)=ϒ��D"O�| ���ZO ��V'_Pĩ�7"O$��ɉ!bJʐ��ŝM^`�*c"O�u�掅$VŐ��F��ʅ"O�hp����y{�������u**da�"O�1����(t��5���\|�"ODC�*P>�~I2"��K��E:"OʤQ� �c׈XY�j޲'���kT"O\!h�J]L6]J�)�#w��)9�"O�|3�*�c��"�">/m���"Op}�bi\���UƠ�i�"O��K'���C��6m�@�"O&��s��@$��c&�ٖ�`JQ"O8+$���YHv(�!����ؓ"Oތ�F/U2@�J��tcϗ~$Mk�"Oظ	�]����b�Ѐ;J��3F"O(a��M��yv�_�2g��b�"O���7g�69��d���ԝTdp�+ "O��J�D�K(���CkT_E�$�P"ODQɣ��-3��{
��
�5�"O�!���A�zQT������?�\�0"O��w�_�?.<m���\Td�b"O~��C�D�"�����^��B�b"Oz]���kFb����$9��4"O�s�'5x@a󂥘�s+&�"&"O��(����D�T��dB،n�4�%"O,)�vaOHZ���CB��:� �"O0ĩE̓�I���c�=j� (Bg"O�T�6#ެz�4��L�9�|�J6"O�eC��4 ]���+w���3"O�1��D�-�$��5`?[Ui�"O8��-G�r}cs-�$��"OJ�f
� �L�(�ՠ�8�(T"O"�h� �n�NT*���/��,�P"O$�3 U(6S�Ar�Ė,��1 "O�@Y��Z0j�\�X�$g��0�"OĔ���M�%&bY��ڧfZ�!�"O��X���.u(,@� #K�a:b"O�E�`4T=XP8�?.*�q�"O�XY0�ӦaДr�Ò�JT�W"O�Q#ahS/(RzXb�E��TYF"O���˃:��`�`Btcb"O
}A�� n�ܰ��ʃ�.���"Ov)�5 BO�5�R ;t�P"O�J5ɞ�'����.ٜ8k��x"O��J�� +����.u8��c"O�9k �2N�Պ�a�RW��F"O�5P��P�MZT����N4�Qp"O�:�(%'t% �@����"Oʍ{@�L�
 }*@�J&f���"O"xP���Io����ϞL��y�"O�pp�92��Y��Ǿ�
��V"O� ��"��/r#�Q`6���d�@�KQ"O��{�ϔ|%J媧�P�ymei�"OȅK����S���Klj��"O�u���B{W�DP���4l:t@�"O$���&G�b�y���`��"R"O�Th��\�`��|s�b��1Z=ر"O��T�)�TŨ�[,d�Q�"O�+'��]�!�Se�0����"O�d����r��]�f
�?Ld�a"O�X8���"Z�V	S����0�"Of!��*;�1t�Q�z�,9��"O�d:��
6�y���ϳJ�����"O`�2uN	�&k�j�	��9zs"O�\k�b��"��� ���!"Oxt�EI9z�6��؎2��u*S"O��X1g�i�r��4a�0}QS"O��I�+@�c|�mX�� vvT�@"O���WF3F|��n	�p(	�"O�M���D ���V��bSpu�c"OvH�AЗyX�;�c�2���"OjHxg�&�� %��n.��3C"O~	��K¨g�1%M�1X K�"O��aN�8�dp���#.4�"O��D�&i���+rD�=e+h�S&"O*�'�;��j���(T2NQؗ�'��'�4u ��H�(<ja���~p	�'zB8�pjA��A�g�Q�$p�'�b]�Wc��4ѷ��PIf8[�':.�f@��H�V�;�d �HL��B�ay�惊kv^�+�a$'h�ȓl���ro:B�|�c���;$�D0�ȓD�P�����dj�Q��b��M�x��^5z��F+)k�tY��k��20� ��=S^]�qމFԋUa%�H��ȓyT(�!V�&w�̋��#�xć�@�4�bU$L?�����n�����x��'�6yG��[��\�VӌKQ:�h	�'�,h�gȣU%��Q���mF�$��'�t$�7�Ԥs�*9(���e��$��'wtay�I9w8��.�HA�'���/Ң:9ƌr����-�B����Dq����C�8�����6[J� D�3 �!�d�*]������X�\��@��6�)��=����N�8��_S��"#�!D�t����`�ġsa�a���#�����ziΜy�&�;z^�@h !^;{�
m��r�  x��>�^�`a��#9���ʓ}��(IEI
���5P4&��q�|B�ɍW �腵U��9
H�.D�zB��!q�D�g(�$~��Uk7G¿`�:C��<����RG�,�R�Q&6'K�B�VM���
)j&
�0-�8$rC䉘XFZ\y�c[�C�:e(޼g���ȓ�<�b�ȷ?(�1� �Tt���G�t|ai>�1:��W�+-�<�ȓ�hʰb�m�R�������5��?T�zrk 2���ƍ�=)�]�ȓ$&��a I^-t"��w#>\��r���Sn[(zxq�b�TK�V���F��<��ɉ*:V!Ѳ�Cc)�@����%K6d�/����vͅl�29�ȓ5��c� GTU�Ŏ��]��9��Z��Ed
ITU#f�ȓ��$9q�Q�_o���I2���S�? ����)D�H����<��s�"O�HVAǼΆ$b�	�<I*���"O�	G�M�TՆ�(=��:f"O��8B��$/w6\P�D�=~9�$"O�+�8nW����bտ"p�Q"On���-��W�q1Q��4��q�b"O�� *���qe�6��Q"O�X[@����ic� l��M@R"O��"�j�=IA�2eͺn�.�XT"O��ؒg�P<i� Cѐu���G"O��!�ʆ	E�HJ�!��U�`�6"ON�0D�&��9`���~��U�#"O�8���M:y�6�g`��n<3�"O��P�K�ͰL��/\�?19a"O���F��-_��P0�7hj9*"O|�+��$^UL!�D�Q53��H�"O����Z�$+LıW�][���"O�P� 7B:a��/ V��(r�"O$��a�n�8a�����Kn����"O�� %n�W��������m��"O�,ɢj���=IE��˪��S"O�(���©r2�e�]a�"O��ٵ��>�t�����.)�8�*!"O�� LB! �B�;�E�Q�R�"ON@���;YB\��b� V�h��r"O4�0m�ZK��hT��w�����"O�h���{��� �*˴-Nh��p"O�-�O�(��@��.l���v"O�,yCN�V@�H�g���9ΨQ�"O���&�֐��y��fC#�t��"O�J2%5�.� Pe[,�� "OHD9�B�(;H��ƭW���8:�"OV�h$IO?|�Ĕ��Jڸ^��t $"O�5��W/ET���(]R4m[$"O�a��Ԕ&�V�XW��A:nmA&"O�T�-��C�US�`Ϋ<����"O�Ű�*�a�����קF|A��"O�����
�(r�V�3��(w"Obx��J�O�81���~7��[E"Ox�S1G��J��Ƀh�l|��"Oh@�bZ�x���̏h]�9cd"O�\��kĥ~��WkC6`�pق"O�sE�"'?�%�f�ˉe%����"Oĭp�霝A��-����6 "Od�9�H�0:�,�H��k�<�!�d�uTD�j�坊�[r��a%!򄓖J���:ɶ)Dk��+ !�ئ5��*$58�Ƚ���	m�!�dJ q��uZ��_�t� }8w��Q!�$�6Ǩ�1�&����|P��ϫqC!��A>�2U�b [	o�F z.ڭ�!�(D�Rt��a����S�80!��>A.� u'��.�v9�яR06,!�dU�Hg h  �   n   Ĵ���	��Z�Zv�J�(ʜ�cd�<������qe�H�4��S66<��ʄxG�f�َ%� �8�MαmF���򄒻�7����۴ub��=�	Xy�dݰ|N6��#f�%~rN �E^+Wa�:��]9ap	�=���3�l�&6�	o6MhP ��=�r	���G1���Æ��C읏8A�		9�[�H�y�If������`kP��%m�<&���ťR�Y��MN-c�0E��$S��Lj%˱?�I�'�X�06*S�!RHHh�A'$-�$��O1��2r��By��G�FO,�0Fk�O��ϓ&}�|�E���y"�ƭR�#���;>+�!2A �"�~"h0�N����	��I6�ꄹ���5Jv�g\�a�DW��۶O����K&�\�b�H�iu�;�X[�h�a�͊c%���Ϗ�[��y ����O�����^����
^n��U�
�~L>;B�!L��'�f#<Y�D �I�h<ٓ"�� �`i�g�߹�6M���O\���D��
a&%�1 e���RD�ڈ\J`�s����O�!�O���T�	+`�p&��X�����^�����I=vO�O`�E2�.ɰ �I~�U��6�O��;��DI0�?yC�\==���RRHKS�TkDP̓zS#<�T�5��O 4P���\_�A��뛳-�d8�Oʭ�H<��-Z�MK�G��H5�d c�S-pi�ԚG��ßp{�u��
��S��?�2�>���~��d �j/�X��O�UL,�q�d�?�OJ H�x˵˞9���5���*	��μ>ѱ`9}:�#<9���;9�+��ʴw�e)Eȑw�<�qN� 2  ��*�Of��e@�&+�1sN�9U��)��'�� 3w^�yվ�+�h�O�U�#�(-���v�C"�H��"O��S�Vu�tx�e������P�|b���NA��Tm�xun�}�6��_z�{��ѥw|B��@m�J�<�p��D䘲�
�� *V��X*KzIpI�	;.�6M�*W�BI��L>)�f��.6
1tDD����E(<I���5r�Qf�M1(xY�A$���X'O�<�V�������z
� ������9�q%3��I��'�@�b��Q�ka��]
&`�l�҆"M�$:��N�{��������yB�3hv�!s�o����0�����*_Rp3�i�C�y`�$�>EQ-`�D��ț�Iq(9�!?D��QPїo�6�s    �    �    c!  �'  �(   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic�'�C�\���E۠_����p���T�?D��x��=X�`�JTԖ�Q��7�	�e��)�A�Ur�O� 9s�jƅQsp�r�W�U���'z�ٲ�	D�LT��R�m�Eg8S�O�;@e�@]���D1�g~��:FFF5�0��8Pe���׳�y�d�(�R�+���:�P�ѡ͙&�&��E%U���y�7�'��0q���`Pp8WÎ�� �a�A��r2��=/��@��?#� "��71
J�ভ�/c�1@p"Obt��������)W!T��2�x�C���Y�mJ�.8<9��S�5�E�G��*u6���@�%2ǂC�I�ut�1�)�]Z�<�bӥl�YC/_8c2`ڡ�ڃ>�6\�2�1�3��ոkT>�y���	UKD �2�B����d�j�Ը�6nO*�t�Yˣ )Z���C�;*c���EG�%a�=��>��x�!V�U�7�
dJ��+O¹3Z��Ǣλ�2�����A�J��Px�%8rcX�l}v$��.4���C�P�^�XNP�]�����8?���0;:��k	��(��C��O	 ���.�1gb@3L�X���'�RP�+E �ީbF"L�=�LS`&�!9Ruv�
&$��ڷ&�ŘO��', l"bb�Z�(��S�sZ��	�'� m ��>A�l����$t�d@"'�-@0��0���xܬL@�E�!d��y��{$}��5����f����0<�$��5|�; sU<%{��]�? ��1�
�������R�C9�K�J94���r�2'�ތa�d�8]bl�3�5} �v���Bo�1Ў�@�l�{�O�
ycuȓ6��MB�N�F��y��'�](� �(�`�eH*Ġ	��Iϥ2�P�����]P���F� ���G��Q�Y�MY&� ���0w��̆ȓ0��	�LĚ/�Px*B�Պz�����`KD�����b�^����(U�S���4rHoK1#�a{b�Q.)��l+bLB��P;��)Yd�,;UB�8g)�i �k?D���xH�Ix�e	N����1�	=d}B ˓�J��>)2�k\��8`�#�Q����=D�D�!�),��5�a� _���On�"��v�JC~2�	~���D�-I��mO�x
��c�[.eS!�G�CK.ph�"Z�!vd͠b��\�v`�%N-^EI0�'�h��� ��5#�!�?:�k	�M���-OrqR��J<���:D�/?0����"Oq�"�K��P(� �<Q.�1�"Oґ�⛭n��I�4_�0�"O��h�� 7IEftc�O�@iZ@P�"Ouk�>_�D����1oڜ�"O���e�1YvVD��/#X�Aؕ"O�(����(���.P�3�0�R"O�@B
n����E�Z<3vJ���"O����?
�.��3^�\����"O,tc�,�<TI�qNT"��&�+D�t7&%2�x���`d<��H*D�p�qB_)G}�)�.^UHl�*��=D���c��(��(�``�)u/,���$>D����&6WB`���s�Rx`�.D�4@��E 9�z���N�0��1"'D���̭� � 2��B��@�$D��B Z�#�L�`pmV���I�%!$D��a�Ć ��G,	���ԣ D�dk�l̊W �:���7r��ū�d-D�u�M�T��a@�	<��A6�(D�  ��<ܩyr/=�L\��*(D��+$��hY,\��l�y�લ-,D����m������*�$9�.D����B�:�
�D?�d��a"D�(``�:c�]7���:�i3#�<D�,1c�0U��#�dA�[*vLAG�-D�Jt��|��8 �Dw�( s �,D�h�.%Z��E��i ]0Ѝ�Ţ?D��cfNV/%ֈ@��' �Z�r׃?D��ĸ-&� 4	�%"

���<D�$��΍/dZD#vf.� ip?D���T�˩r�~��Y4 bj-ЗJ7D�����;l�x�%� �\�K��*D��kP��qr�ʄ�Jo$�q7	=D�8QqD���A
%I�6xq��R6m0D�x�g 
u��zC�Ӂ�0��:D�Ԁt'ǉ���qc$"�H�#�8D�tju왉N�҅�'ˎm�H�7B9D���c-�f�`���9�"���%D�4rC��(�O��.^P��(D�,�AJ�=T����n&���E6D����l+>��z�Y/����&D�̉�޼4%��zT�T�P�x|�#D��G��e�@�{�JS�=�<��%d D��!�Ȓ�Ix�@��'R�J����3D��Cp͎��0��&��F�@�3A'D�� +��:&d;�%]
=���R��*D�� �>4���=Xc�Y�/7D��j�)I���9Q-�@Rp���!D�0`�K0?،����[��\�,D�� �A��#�Z�j���ڝy��Q�V"O��P��\�RM|4��2 ��W"O �aa�9]�̰!t��"BFV�xw"O``�"�L�I�$uAg
Q��v�"Oޜ�b�])!�����菸�0��"O6�vAD�!��M��I�+e&���"O�x�Q��o<K�)\�W!��"Ole.�
-ሑ�a�F�	�|�R�"O*1�q��Ci��z)�1�8�	Š�9��!8�xX�dKE\*Rd��e��(\L$P�!D�HQ5�
�~��Bd&@9P=D�����9H�PU�c�]&?�i��B<D�D��A�%Ю\���M�em:D�8�rg�
E���e3�Ѱ5�7D��J�,W�y��P��QZ� D���)�=CL��OT�VQJWi?D�X�P��0$�j���l5r��@(0D��s ��%`1��6�-H�xQ�/D�|�FnF/T8)��i�f�Y�#2D�t���`h" �Wf\.FQ��0D�$�ua?<��Qs�.ڜh Nݻ��9D��SG�'��"�+S`�n����7D����D.xs~qP��P�T��$�! 0D�8���U<0^�����>k�Pix�1D�P���A�,�{��H�9��D<D��35��T����wI�o���Z�=D��A�[15κ]����(l9���$�?D�d"r O� ��3��"c��H��<D�� Sü`e �Y�H �hv�����8D�T�B�.���J�I�'N�{�3D��80#N1'�4�����P5��%2D����[�$n@�ᠡͮny��I��<D���Ƣ۲0�e�̚-�`�+RN8D���w�U�������S�&i���2D�t����PdY�*ǋv:�١�*D�8��'��e� �@���#�a0�2D��R�E3iTN,ڥ�H�fl���(+D�����s�%ZWnL�L��&�>D����+Rq�p���]$�r3  D�4c���1�x��g�Z��(cf�(D��#��V*g���B�be��J��%D�x+!@]�lM�i����n�C�.D�l"%&�{�t:e��)G�8%�c,D�t 
�!/�p�󩇳I�
�s��=D����� '�h�	��қHF&�a��;D�����W�?���fc3��'��q�<i�#H�f�6����s�����gYR�<)F.E@��v�.{�L����C�<���C+"9bS	ީ%���h�h�<y��@��Reh�V�q��H�<�fmI%^����JT-W�1Ӌ��<���N�Z�f�ޖZk%R��B�<�O�Ab���b�a^�9Td�e�<��N
�@P앂�ŕ*q8���Eh�<���Y�  �|�OXw�^��c�<��I&gd0�BbeB�k�Hڀ�Sz�<�&�KI��5rmծR\XD3i[j�<��LG� �-ba��-<@�Z�$R�<�2_�}Fq�JS=qU� ���J�<q�(��4���`�#���:�AE�<y�i9	��< �Oߣj ���ь�~�<�!B�gG�]{��!=A�9j��Ty�<Q���>6sD��eMĞ~ d9A�s�<�SK
>0�2�C BN�..����#�l�<� >���.;Xp�f\��Z ""Op����ɠc욜���38��p�"O������\��) kD:	��"O@`
!�O�|-��ٰ� ��s�"O@P@%/I����r��,v�Xu�q"OH��QM�XֶȒ��+%%�u�"O� �q�)��Y E�;
����"O�4c�D�{r�����$9�"O�8s%Ҏ7u ��-�|l�6"OPP�JT6&d�)� ��f�����"O�BU���4�捐��H��x��"O��M
�ZO�-p1��<p�����"O�mL�i�n����<]v�XQ"O%�g�%k�	��\?Zp��"O�����P�}�x���сL��r�"O�<�W�?tтqÈ�x��%�"O���`NΦ)�T�E%E=��ɐ"OdM��ٖ"
 ���?^���D"O� ��v�|=K�ذm�.���"O��� ��������ױ-�|��@"OԵ0�Q�+��@c�]5�����"O40��킠.� +#KQ�l��@� "O0Ar��1��A�䩈�"��Pb"O L�S!ˁ�dc����Z�"OH�z%	׬P�ĹB���azG"O��!%�	�\�f����KR�Z�"O���0BD S��x!�
�FLU"Oa��1]����#�m!,�8�"O*���D��e�dⅡ1#h!�!"O��Q@��!�d: @J)g�T��"O`�i%���u$�%�i�j�"Ou�����8R�2i8��"O�iVȁ1���Ҏ �Ln�m�0"O(����>&`�g�C� xb�"O��BO
z!ҽi���Pm�P�p"OiK�lXV�`i��h�Qxt��"O0$� ��\� G�n�af"O��ѡ�SgC
��Q�M$Yx]k�"O�|E	3~D�f�ͳ2>J�C�"Oa��fB#ז����h��	�"O�`�u��_x��x�����A"O��{�CS�~b��B

�(�FPe"O��Y��W�6��b%��o�$T�$"O�iH���K��-�j��q"OF���T�| ��!��h��R�"Ol1����j�}Z���R�j1
0"O<Ԫ�+[��`KDj�ٰ���"O|��
S�R�~����_�jqK"O�Ȫ�L��p8�X��,�8�R���"O<`A�'ð���`2F���"O�$�ٯ���!R�]=���"O�x�@��5�JM��I�O/�,�@"O���v'ģ~��G;	�X}��"O
�g҃0~X(ö�yIf]��"O-p��w:�x4G� B!���"Op书KŅ�Q0V�?d���P�"O�a
Ul�Px�����j�8�9S"ON�1�3 Z�}9�hR4Tp��y�"O���T��$9A��-�,@�"O�5`ㄹ-�q�2�� f2�ۄ"Of�ZP��
O��ëƱp�����"O �2��L��% M~�"H�"O��1'៰DY6�n kâ�"O@1 �B
��v��v�(X�X�Q�"O� *EX3B��H��}�w����"�"O���,ҹ;,a˲I�>�h}c�"O&d�7-X#9�mYa�Ҳ-_]�U"O���@�ؤiݖ͉W��"_ �!�"O�;N+r�(���	ƞjAn��r"Ov4���.C��Y:��҈1����"O�ܪt���fQ�]	Ř<|�Q�e"OH��4gI]�~e���416e�U"Ot��A��1g�|��vO��Hl��"O�8����N�eR��M"�p�У"O6P���B8�<�'�*l�^p��"O�hR��N�7��l�u̗�^��t�s"OD�Z���}�z!Z�M�=fv�Ȫ"OZX�F�[�&5��
��D1����"O`�Cu���B$@𲗊K Ojh�³"O�A9ݞ.:D��0jʋz�Lh�"O�X1���L󦴙`C�-(�,{D"O�� �+�M��ܓ�A�';�
`""O<\� CP/�p�"��3?�5�"O�,Z�U ����ܭ&��p�T"OD�ȏ��p��ga��~��m��"O�0��화�����8�jq$"O�u:gD\6 ;�@�U#��2�����"O�<!!�	=�Fa;EɃ�ؘ��"O:"�(٥����J�+�٪�"OPC&R/�ĉ��ł%}r���&"O~jai�3�HI��٤uU�i�1"O>!Ȓ ]#0s�h���2Sp �g"O�|@�� \lH1�t$�e��F"O�P��(׮cYZ���,��_��"O>�Ke���@�٥�	2eH8��T"O���A�xz��q��D�G���"O��3��Q/6��!sƭ��=���v"O���ťl`�t����A��Y�@"O�p�Hϋ%"���vH��"O�$o�ٶ��¤K�}� ��"O إ!G��Eq�C� ��h�"O��*p틎+�ԱH׃	�F�,�b"O�ER�n�R�S�?Zӄa�"O�s���>殡#Ǉ���Mjr"Oԥ�$��)jƃU==x�"O�Ő�E5j�R͓�䗜/�ȸd"O�hA�bv��UAQ�-.�E��"OEz��Zg`mi�j�34?ZP�V"O<�����Vu�ӊ�e/jeB"O�h��ǅ(dH�1Xg	V*E�|��"O�({g�٥s�9�'c	o�V]33"O�3�	U���=�A�-�h�3"O�(Q�#��L���+e�
�5����"O�U�� �ZW���'���nԘ�"O���`Y�4��H�,V1��K�"O(|����pA�$�� olS�"O�p�7+ GW��2�)ϰjaԔ��"OVpCFc��N����1L�Q@"O��O�C��'εKݐ�i"O>�$M�4*Jy��2o$>�Z�"O$�hS��Lh`���I�6h��jR"O�i���N�,�Z��!�N�7"O��k�IO7���+Y{�IR�"O���wK��k� �l_:.@C"Onp���%f����6K\5r6l�"OX\��N�1Vᚁ��&��P6"O����C�<	I��׷d�t�'"O0�РhE�5\:�G�rq�};�"O� �M�dKڜl��9����-{Q�1��"O���e�>`��+��23���"OZ@��^FԸk�g3���U"Ox����;�n�[U�g�@�P"O�H��� ��M�W��%a�5�"O��jY�1@�e`��O�1A���"O�A)�
��p{�͔x0�:7"Ol8�Z���� ��u�@�"O~�G�8IS���J�\
ViS"O,���"��~I	Ā#�8]2"O| �Lk��b4CSA��(�"O��ؗ�F-0~ c!�>���{w"O�Ç$�#n��(��@Z�UJ�	jF"O��!��  �   p   Ĵ���	��Z�JwIJ(ʜ�cd�<��k٥���qe�H�4��S66<���EO�f b����Ɗ_)2$���Ϙ^86�����I"�y��D�<!ĊɠH�hp"� Y&:�`�<W�0��D�c�㞤IR�ɼ4��˒*W6�����;qz� �m�=���V�(�`[���D:vVuR���d��(4�ġ��$F�ar�L&[�B!�!a���M[T�Ĕ0�����(�Sߟڝ�aa�!RЁg�\}���G�bU	4����e�cc�!�O�p\9��u~��o�|�R!8����q%�,r^R(�u �!0�m�R�O2� ��<�y��]��3�gÉG�
��Ł~}b�+S���ӨU�j�Qv"�&Gdh��g��>�rq�=IG�8�<��Gj��נ-	4���,h����c
��[�S�x���س.H#!Z)28 SPa!}��K�'-���=Aw����4]�Q�G�VX�v����b�	"Y��\@ԤWDxF�b��f�lyh��� Z*b�|j�ቌO�I1`,��E+_F��6��2X��˓i��#<�0M*�I6���ņ�h��k��7GD♀�����r��'�2���)L/���ˎ�ZH1�y2�NV�'��$&�4�rĕ�N����k ��5�V������I1C�'*v���cbpiTh_�@��Ct�r@�m��Ss��y��YR��'�8�-O뮼�h�_c��Ya�%�8wJ�ko߄|��y���]>�O�3H�(�4� �D8z��cn�!�nt��&�>9�8�;Ǆ#<���L�]�M���;J#� 1B�d�<��h�= 2  �"���oH�w�L�R�SC6Y�ȓS-$�K�ʈ�x�P<�3 \ �"���f�`T(�� tX����"�h=����k��EAd)E�m#"퍟D8���!̪d��<Ԯ�btGA�Mآ�ȓ!���Pe&���f/¬	�"h�ȓz��iҡI[���Y�͒#e�Դ���R��ī=;VX��oWH�@l�ȓ.�|i�2o��R���a�&97�хȓq��з	7_�u9;Et���'���wnƕ����V1B@�ȓc�8Eǘ�<N�� �$ձ\�~8��L)�I��)�f4�ɐ��*|l��ȓf<�mԤH
da�p�j�t�&)��� S�LEB��'�8�L �-�
4���� %J��X�'�\��¦�v�:ɬ�'q�Hs�.�4���[e"��H�(���� ,�� y*zX �"O� \m2�-�5��\�Aˍp��Ȼ �U��,�a3*H���)��<��*�?`�����W �6��l�E�<!�͊6 �t�� ��.��)�����<yC�M�Dy�­=\O�����9�
�`vm�y��	��'�����O;3�ra�E YjN��'�K�f�^0��y�"@�lQXt���T���`�!�4�O8��f℃\Ӭ����)�3d��c
�w��Hq! ҠZ!��77L��r�8k3�I� �*X <@�C՚*�`��N�"~Γ^
T�
�W/7:��yqJ�i�Q��9������Ϙ ThY�p t��I�y|��i�'B��$��F����
�J��ez���a|��
#Ḑ�e�ӣD�d��k�d�5	�F2p�a��'׮���AQ�W��-��������䟁?��u������(�8PI�Z7 �h g�]�>m(q9"O2h*B�\�^��m0F��7o�@Г& �Ĺ�uH^���)��<�Q O/OK���8*����\p�<�B�Sx}� ��]l��t����l?�3`E�-��h�e���G�EU��� Wb����	��"1��'��r��>FP"��'��P�<��'�l���%�	N��Cw�I*���'��mV�B8'����JJ?���S	�'�d�"J�"h���8V癈Bh��'�~(�����<�P�됞w+bɲ���^;�>9(��W����S��0d�]�oK�!�$��P_x�T]�d��!�n2p�]��A'O���hQF�S�R('��O����6Kv��(.�~��7"OD�8�P��%��x H���@@��9�s��Y[JT�'�T/{��I�^�Ԉ��;M�� "pD�8l�
��d��E��9�m (���Q�F��"O��`c��)c�Ԥ�sB�`���'�ea��JSB���AMGG�ȓ�}��2 ���K�e��( D���79�O��b3�_��$�k��D�2Vz͙	�'�L�
�͂0Jz�p��@�(^��ao�+�<(�$癀�A�����7
�,�I.�\�șw��К���P+Rh�Ј5q�X	�']�L��;�7��i�����!ʗK3N�p§<D'�u��-L�T�d��'~2�k$�ݗ��	=l���Sႆ$"�KfD��4�4��d��9s2���}��!�L�$S� �i��%����T�\�1Кt ��H��B�J�K�I��q
�'�M��`\��� .� |���B�y2N��~�����7h�4��h�-��wȏ)7�e��[�I�a�$O��CBڇ#�Y��'/���P!�z�b���J*�0R��Έ�T�'O~�ҙ�AB�#-�����|�l���j�(� z�w����5F�h}� �G�ۡ�i	�'����Ռɍc��X"w�Y~��e����Q�0��H&t��e��j�_x��H�,�a��pz�
�y��M��O$��%HBaJ��׌Ϝp�D�	�v�<1��]�\;rAS�B���%C�+'H1I£�.C���b�ه^4�͂"�$>��bĬ�+S֔u��	�;�6|b�˔1n"ɚ�����RjȘل+וO
�eKpi��L�r���J�nu������� �ѱH�y[c���N��AcJ�sH��'�� c�؏wZ"�&#���s��06Z�� w�D�@mօA"�9��(+EtP:�Ɲ% �䑛wo�U�A�'X-(���V0$�~�K��5j�}���C; ��q�РxP`1R�M�^�$�c�A�@�1��E�"6����O�r�(Ѿ,��'��)��Y*6�����[�:��э��d��2s�O�iC�hj�DV+pB |{
V�t��4��2;�:æ��6v�b˓>���`,;,O��[��LUߊ=9!�E,����V�t���W��+�nK�#��1��ն`LL�>i��'�M^�0���i��(D���Ñ\��	1��t�M;�-�H7�������s'N5 �l����c7�>���I�F*B+�? ��K�*P<�3$]�|���H!� "ZM ��UJ�<T����w�^	W 4�����X���۰<�D(�2zz���g��n#s!�J8����j��x�2h�L�A)8���@-?���`5B��7�е� �"O�5�6
Ͻr��m �B��$� �Ap��S�I��h n��Py�#}�k `t ��������
B�<	D �8i��xK�i��;��ġíѡE���v+w��b�����H���G3�Y$F;Yy!��H���j ��n'���f�F�W��	���,���Vb)|Oi�DꄖVy�\��3a[�j�'n�2�ٕ �V)��i����NS�R�~dpG�(�6��	��� "�zv!���Ԉ"�O�rU41����)�Tҷ�Ա�h"}���0@|��70x�y�@Q�<A�jTXP@�`��3$g�`ƬZ7�RE��EU�dC�I�k4Q>˓��8;��8�����[�&����ȓS0R|����l�F�rQ�R� K^�l��u�rm[�T+n����O�]C�:�d��qmH�y�{r�֝۞T��g��������TO �ք�`l��+D���
W>Z�^-qg7p&��@�+�I$V�Y��蔯~��>E�	��}��KH8RP@d"�L)D�����P�����K�_&n Q4-�;}_�"����	N��~Bi�)H�M�1�[�nɚ�dņ�y�k��(JDO�Y�X�"P%ƍ�ybI�#F�=���'eĂ��-
�� Ϗq��x�?L�9��q�$��P7Qф0�W-�7=� 9��-D��p3̝���,��/[� ̼s'�&D�$����r��8�X?�)��"D��:�,�
1�����?zٔ@
C�>D��Hǝ3^μa�`�fN�ɛd�>D��h4(W�s�� �Q�Jt����+D����$f|��f!M:L�6'D�l� �$kVӃ��.��ܙ���� I��eta|Riؕx30q	AK D<�u.�0>)�`�.A�xa��L\�{��4S)����ۢR�\Ʉȓ=�B��� zg^9�4���`�|������	�g�O6�#i�|�ӌ�i�:���k���y ���G$!B]B�nSL��3+-i��5��Q�FĮ8Ѷ���=�Ъ�ZL��~�� �u�+@�؊��U�U��K$U�.�H�㉒V�R�3s,�Uܶ�sPJ�<�h̀6m3~`p�A�V�W��X�!�'��`#��`���I�$�N1�
�+���@�+���W$��W ��V.��+0^�' \i��8|�B=K�N۔Q~�H��^= �7��!��]G0-��&R�}��ɂP�ڠ(ƴt�DҁXa6��G��-@����X@:%��O�"�+���M7g�q�r�U(:� �  �J�5�az�j�A�X̓^j��h�DηE/���d�Q�0�~iI�״SC�|;��N
�`�ח�?)uϵF+����!����'���t�է,��"�h�Z���L>)��CX������@RU�2'ت�2ԐթK���	�'��<��Q���l� j��G6�?��l��$4q�FI�G��y2�9��xV��j�Yv�J�T&%Ё�ì�1U�L�1�H��b�'2b���<���iÌ  �tR�R�z�rP��	\�2K��j6$C�ɽT�.� �GD�wdA:\XK��ζi~<����dB������r��d�V!��? Pp��z?1Ǉ��=�9X$�O�(�x2�݆Y�=�`"$,O^�0��S��<kܴ
i��T\- 	� �0��K����^}��ѳx	,e��Oqy��W
A����Lr�I�0a*W������5�8Od=ڥK��`e8�4E���˷��G�b��� M 'X�]�I�(��H��1��dQ��K�:�Gr���
�FY����آ;� |�b�A�\Y��E�Ơ���K�O����N�R3d$���S�|�Hَ\N@ �vb����?�Px���o�2�90��4��"�+1hn��iқ���.�,��f�n�>�) �n�D��|�n�7\�
��Q�R0[�4XE%FjX� �c�$c�
�y�Z���
Z*:���.�-��)��Dl�^Q{�4q�ص�M�"~nڮ/,� {Ce	,���@�
x�O��!���z���	Wed #�UNJ��#KY'��I�l��lj��\X��y���K��ģ���en�(X�ě6k-���=a�u�'UN�u���?K�`c�Θ	9�<���9D\�%��'�MԋόO�����,L��C����h�~����]�tY�� E�%n��!�CA"�!��ŗd�`T!wj�( �sR�A$D�!����`�pP�
�����NS!�#�ڝ��I�O�
�����%!� w�y�$�.Oٔ"t�)P!�dӃZZBa*QkRC����c X�m	!���+z1�(I&r��d�q�@�K!�$�φ�H$h�03�� ��34�!���~�0��6.ǁj��\��n�>}�!��
Y�XXcCY�f���@�^�!��O5��e��H��S�Ʌ�e�!��Q�Pd�O� t�,�!�� �P�c�P4"i�Տ�mX	�"O�%8�mR�#���0D�٣[�T�4"O����BOS$�q@!4��"Ot���B�*�3R��K�Q��"O<�����H?��� ��Z"O���K�#b��S`�C�p�L*"O,}ᔯ�N"&���Y0X�hٵ"O6���(��:�c7cP�P�XP�"O` r�F�M��2�m��~��4"O�i�ӌY4̖�a6>�%lO��y��ا[�����Je��f�A��y҉&0���0�(�NW�����'�yBL�=�f��̩~e���b$*�yr'S�I�v�C ��8`�ĝ��y҇G-"B�D�E� v��yF����y��{��er��}b���(:�y�Cԛ3ʘ����t�i;�H�y�䞁,<���˜�\�*�:!�R"�yB	�t���Q�"��U�>i�`���y�%�u	<k�њ������D��y2�/'N�,rC Ս�&��Rh ��y��I6O��2���3}�e:3���y���7ܮ%���
5��(٢ �:�yҀ�j^��CP� ����=�y��`��aϾ�����&5D�p���70��d�68��-3@l5D�hj�藇:�%�Y�^��c7E<D�p�bF��\v���f�U3��L=D�L{b,ښ,h�
�'F}�)ju�=D�8f�66t�k� �[�4�91F;D���2��y�ұ� �U>4��#6D�Ъv]�K��Spd_�jt�27D�D�2�Ջ@(�1�?�ѐV�3D�x�1)�h�EJ�C�	��a�#:D�����6W��+"ݍi����%<D��3�IǢK1�\8�iO/� ��(9D���ᄝ�nM�A� �>�ꠘB�4D�ԋ�^W�����	Z����S�2D�3�N
h�N��`�K?v����2E3D�8��4�>���"ǖ{r-
�#1D��(��&Tg��9��ѿ7��(��.D����dE�xAK��6�zܠa*D��!!��DX�X3���8�T�r��5D�8sB�'A�$T�C�^�^sD3D�����ɣP��l�q��.���Z��1D�أ�hK�WX.3��D=D�� 	T�"D���a�v���y��^?Q��QBn5D��	�Kфej����Oe����$D���M�\�x`�R�(�j)�c#D�h����nn���e�!^��1Po2D�Tf�alHU{��+*.=��3D��I��3s(�ّ�E;7P	��.D���𤘋+	Rܱ�dB�y4F����.D�$1��Þ*��ذ��/�:��d�1D��{w@�C���� 1T�e!�5D��qnO�e��&� �Xc�'D���N�9Ʊ�P�S�<^�`���0D��١�.�R���]�~zu�WC*D�8����&OC�i�O۪|i@�o+D��x6��	"Q<�i���6�HA��c&D��&$%=T��Y����0��Q�3D���A�G�7k���*
2����!2D�`�І�F��XЂi_+���ڤ�'D��h��߅>����%�ڷ-{�)׏(D�� �I�F�"�S�]�xK�0��'��)@ �$*CI�&g�H�@��������rd"D�h[5鍽{�ޔ1f��<Fl�\���"�K� |sei=�H�(���n1(��q���$�ʅ��"O��� 6��Irp��H����oذ}g|Y����)��<�qN�xd-��/� w;��T�Mx�<��%A0��k5\6����U�<q���)���a�%3\O����#ˬE����F<�)�C�'�,���X/�L����fA�A�*W ~e 		�	� �y����:ij�l�6l4� ��OM�@����&�(��Ă$	B
d�^�13��0A��S�"OY��� ��!�f��()��Z�Qf��`�H_#��)��<� ��1��E�$�~5"(��G�<iW�^�x�<��w���e�����`��<�g,CzXr�`&J=\Op�z���i�C�?	X��q��' �U�r���!�� �C��"�����m0Bԓq-��y"BʒY�H
�k��b}�q����Oꤢ�� /����$Xk�@iU�4#2p�R �Y�!�X	�����L$T���ψ1(����Ѐ��*ږ��L�"~�|�����U P�j,$�@�ye�]�ȓ_Q��X3�ʀH��L˲(H2f�h�ITP7��Ű=�`���&����!ȝd���
ҥFX���5��	B�E&,���L1hQ��,�$�y��؟z3�]����3�����ą�y��,ݔ���'Q9#,��C��y"fɨQb�:ƂAA���p�dѥ�y�Nʊ��6�M6.P�@�K� �yԀ)��MΫ_�`�Wƌ�y�EM��J�ΑLHμ���A���'Iʴ���R�S�'9
�*�̜<?6�H�HD~�Є�"�R�ʔjR.��cA����FQ�o�m�ɱ�LE��Oq)�%ά0���Ɖp�IjdO�t�&B�ry�s�,�6d�!�#�Jg,���_���>�0@'6Z����i�NR��rA��wX����RM����R�h�Ԣ�=E 49�a�0u�i%�-D���ǤK
��[�	ξW!�PL*�S~!� "�Aؕ�M��B4�c?����t|�9Q�B�#x0X(��+D��dM>Q����F���~�᥎I���+۾Bjn諁H�[�vb?%�Odhk�a�0c��x�5
'd�HO^tЖ�&]�򙛣LA0m�SÁ�n�tQ���߸8�P q��<0l��I�� �ʀ�ߒW�(|`j�"F!��D�>&�lm�� ��D�J$1c��$/�=��"�Pn���Ԑ� |��\s<�󌅠>�f�34��k�(T	�%8�\ ��-����Y�L��:U�ܴ��D���%8t�	���%	��n_�T�t��-�S�r��B��!�D߄V��;�lK�(ؽȥ��/��!y�� �θ��`�	YTX���o��% � e^@U9�NE/,�^p��O�������y�<H�E�-�H��I[wZ�)��]�r�hR�̣i&t��Ռ�iq2��$�'3r��C��^����v��	aO�eb�'�;1)���2/����:�i��Ǻ:R��.8L��M���h��ǉ``�(��ďi߈i��.�|�h�o^��ZQ��N�-e�bL�a`֩
�ꥨ�'St: ����UA���d����V������^eo��za�W{Sv@�O=��]Y�F��|���w�N�x@Ư~a&މ|"�=���h�@�@$F�d�b}	�'�Y�]�և��QKz�+��gv��eˑE�I�fr���%�1��S�~����e
/���[q��*=�џ(��"�/��aҖ/�2|�������@cœj�>�����$�h5���|��]$�l1��I3+������<r:0�E囚g�\˓C��`L�j`��#u��j�|#}�K�P��u`�"^-vl41y�<q�H^4{H�r�)R=Fp�	��E���yy�G�)6�"�sTg_�)Xȭ'?�ԛb��)zc$���lڨ�`c�)7�Ћ")�kh�IW�#3��U��ʝ��=��!Vv� $S�e��P97#Q�F���	Y@��ݰ�O.OA���fw�3cF��y2�g>�3ǓQ�F���A	��y/�q�^u$_*1Ķ�X7-Y8��'�n��6l|�G��됇@��8�Ԧ�4,�Y)6��5�y���-b���y�m�.[�`�V+H�+B�B6l�����:PQ>�S�? 4i���2u�Y���S(~��M��"OHI넀�) <)��,P8.�>4�4L|�R	� ��ă�|��qArخ��r�z�"ܷ.q�C��c�X]�� ւA4���	��y�ꝌG�P���/?k@�ywa���'"����N�P�t$��Ӿɪ񙗨�f`�8P �I�C�I-+�.���O+Q�paF�5N��͊m�X����*O:�K��Y�TA5b¨]�s�Eܹ[� ��!/D�Ќ׀TZ]A���1�lӘ�2��@(,$��J!�'���5S!`Z@ڥ�9$���
ߓ\_T�S��^-(�
6�M�cOZl+f�4t	���� X�Be!�d�t[�����P�S��[ i�O�m; aL(�R����0�`�F�uY�2��2o!�ċ�ٰ��jVH��C뙉'�̋��J�b��OL�}��9�xd��M�હ���,�� ��$B�䓼r��K�F�MB��ϓ|B6����>��=�B�CJ��yI���N%fmb���C8����Ʌ�F�d]��Z���n�=Є�G��,2�!��=w�A��@��!Su�ǅj�!����ad�@�G�T��b���!�Ę�}`^��ŝ�D�{G�~�!��L�cU8a��O㪬�T@D��!�""�I2bo�7٪L�m��\�!�F!L|ꅩJT�i�aPSU#|�!�DN�!].@V������Y�K�>X����VP�0��\��@Ӗ]3�0�$stم�0o�*����̟��gJl��%냯K�l���Ǐ,D�P��/����$q�M���4��O q)`�ϒ�~�eϡR����G��A�O�B�QG�j�)�)��n<Q��"OHi�dI�0�$0�%gG�e0��7�O�@i@sJ�Yw~�Q�'Q��Pb��h��Sq�{�+
�TXђ�,ON�����`�*z��05	�`�E�5,�M
pj�aB�$	 �&�?I�Y��N�)v�/lO~ęU�(d�#��	/s��a[��r@��\�����ȍ=���0�����)�Ŏ^3j���[wb����s�,"�
4v(h�'۸��@k��`pC��P6z\6AX��
�.���F�U]}��eaנ��+C�|J��y[8Yp�w?ęz�^!6F)ф�v�p�(ӓ��`R�*f���A�U1~�~m�b�Q;��QwkI(�q��ו)n��î�p�����'{�nu�Bf�
>���<a�c��98������i���Aov�h���/Q��P���N;O�!�֌@
�Q3���*Bl]���J27زP�s�^+-`M���x��8K���$?��]�
�8�hy5�?ZA�b%��pf�8�S��M��ȂX�<Q N�Gx��r�����
R��h�g/>k��,<�y��E��CL^�1�
O�%��HD�RV� J��J:�L� o�m�T�J��ȠO��{A��#���ʖ�ĬQT���z?�o��A(~K��M��8:�F8��l��F.,O��IԨ��v6��48�]�ʲ�����[��0�$k�K�S!�K�I��= Q�Mcy2�E�+�8�� �a�~����V03�@���oFwVO���e	�<����4k��=�e,��R�:�q��t��}q��n��
���S5Z�j�@��S�\��e���I$�'^:h*��A� \t��#�Kuh�� �B'`i��@�z=�ԉ4�W��h�0�ӼYa�ѻjP�6��m��_��ć1�A�fAV5���u�B-v�ب�E�$b4Pc|��b@g�z[I+���V4��'���S�*�t�@SN��*]3u.�9@Z���:-I�Jܶ��V=9l �$�Kc���!!M1Λf�G�	��� Hg�ӧ������o#�#d�����R�@������z����0|J��ǺC�l����}�̭+���^}r���7����4.Qx����S�}��9"�)��;�M0��P�{�qO$�p��@	���S���\J�@�{� %��i�`�B�	't�`	T���qKʘbC����">)��N-�ȣ|T�<(��S&/��?hpP�,RP�<����7 ���)��w������E�<�e1)�2�+�$S�R�١�%�}�<�a��F��KvC�K2�a2��}�<��JC����j��MG�%��a�b�<���Y�FE6��dɚP�P�
Z�<��k�$��$C�ޛ0��@e�P�<��8y��@�<��UX�+Q�<� �10W�'%jl����ш,Z�`�"O�"�S2�|�2�S�6� �i�"Oޠ���n0��a�T/��Aiu"O�����ОMU�-�BgM �X	�C"O���nV�>�y�#HA�,��"OpP��İ*:�X��S�1�65!!"O�#AF�1vq��"�����"O��J�DL�ð��ʆ��I��"O�\Ba���B`Bn �?�luӴ*Od�Kg�[��=���27�8�	�'��]�df�/;Y �*F�%�"��	�'�EG�D�i����/,l��@�'Ǟ)Q�(���L��ō"e�f�#
�'mx /�fz.��@�>^�0�p�'�
�p/4
��p�G\!y>�8	�'��i��W�� ��g���49ڽ��'0f�	.$r)L��e>Y����'�(���fϨ��i�Dȣ;���'��ar@Z�,� ���5ː`��'�t�����]�T(�A�.[w�Mp	�'��,	��R-Zwba1�W_����'�j%0�ƈ�3R@� O�W����'à����/�8�d�E)�)��'u�x��"ε��*P
M�:"��'m$�Z�Yuj�R��F�2�6���'����cH�,���fX2%$ٺ�'�6T37Jͦi4"Թ��(:f�'�~-���$(�F��$C U�&���':a[�$��n���\ �����'�~i�e�֓M���1허)����'��k��>E|�a�`���_�4��'@ �*�͂c��tBӥ֟C]��a�'����`��7���z��;�8I�'�L�鷈:w�ā��$֪S���
�'4���V�^<�%� �I3��˲#)i:��Ë�1-����|Oȝҁ@�Up,M����<u?�]��e'
�y�헰+�����������L���fɊ�ohy��,�D5��ȓ<�p0C7HY�{@�T�Hr@�ȓP��%��^� ���F�e����M�����G3V%�-�"NQ��b|�ȓ*T�ƭP���ӧ�	����<�ÇGI���O���J�)V�@Er�Dd��
&��'�`7��؍�'���B^w� �3?�')�d�$�4J�f<���V\���kFA��E�,OrE���O=L��W%]�,(�hT�g�B1B��T�|T�	U���(1��	�fǓ0��	�M�d�8 ���@}rh�6i@!�֡@���	Ll�OE�Ub�H��%v�u��h^B�HSd�V���Rr�7��%���O�?�yPƋ4%�А�œN�	�1Ad�L[�@I�A\8�'���	ׂl}@��"l�,xԜY�)�ZQr)��'�,Ô���Mx^Ԃ
ç)�R��G��jѨw,S�R�x��Ż�~B�=c�P����+����O� J��p��cyp%%�����8=|E�X^M%�����۞r��d9�����d��K�UD��!7(�<a�kFy��IZ�a�J����w
L����تΦ����,��	�'�8<'?-8I~�6#�20eb� �q�$�6"
�h2И�0#�V�m�;a"��}n:�+	�{Q��B���=�4��/O�V������������|xX���S�{��@�b�*wU�  BF� @�h���OV��'@�2S�W�?����j�|_�<еJ�xg(%�@K}"��.U[��3S	I%���Z �\ �+ZGjX 5l�	C�D�$�����x�f�E�~�>q(7���>sPF]JY�@��`��S�p�^3�ݠ��Tb�ѩ��\:�!�$-]��J�O 7.5ry@p��
%�!��/1�X��AӑL��(c�'�;e�!� 
g"�9��L�S�Z���O�i�!�d�>.(*yJR(�8φ(K#��2!�� ��S0��?iT���J��p��E��"O�)pE�ڸ��q
���7����"O��!���o�T�ZB���8k"O>�`%o��%���($���mrX��"O�I��ŨN�@"q��M���ɐ"O�h��K��P���	��=A���"O�;��Έ@r�� ���0/2F"O�%�`����	�b�:"W�c�!�ٳBl⸒7/��>i�	�v�ͧN�!�_�S��`��-4hf��nE	2�!��4d!�Հ�m���P�L�!�FY�<=�;U6����"�!���I#���'��I�pxQ�B�[�!�P�R��A{U@V�H�P�����&&�!�dUz�>�o"Z�&H� ��!�DX%=��b��&Z܈c�.Sk�!��-_$*w[�byI��"!�=~�,���@e>NEZ$��'p!�^�@�Z�0��L����-z!��2�`�"�F�SH�!#g�<r!��3WO��j���a>��B#&�:gp!��w`�t%R=r{7JB-S!�*W�|{���-�T���F!�%)�����_�m{�@�fA�$)!���{���;rT$d ����>Yj!򤌆@�T�3b����E���]K!��[�R��!S o�w���(r��y�!��-?���J>|���T%�?F�!�d�.���g#R�tx�U	��aK!�D��_a(��ԁ̏P�ĹQ)B�#F!�כ[� �k��(��	1����m�!�D����4#P ��0Z� T�A"[�!�W�y��q����O�@�	㉈�!�L:o�.Q�q��6�D9� ND �!��0-PZ���ʅ
����Т�!�ĕ�GjLfB�Ut��qɅ�!�$=xޑ�a�: �r��6)���!�d�&@E��
Ԣ�F*h��P탄b�!�D�>|�t��$�Ux��<�!�d�F������'���ǂ���!�$)3��c��-Y4Re)G�N�/�!�]%o����ʰ*w6h`�R�y�!�$�?����ӛjZl}��`	J�!��͒Lŋ�̃{���@" ��8.!��LJV�P�b*��e��rr�̇%!�DÁZBJݲ�	�r���3��|�!�o���`$Z�t�0#� �!��4E@0�#���4#�aD�!�
'��4��([c`��+VN�a!򄛙R�&�3&�8nC�11�lS6rP!��VG;Pp��M�P*Z}��J1%�!��Ǟx	�B�3��*�jѵF�!�D[>Y��ģ���0FըQ��O�!�dNcs�HA`��� ���*�!�d %-���1&a  �0�RW��*U�!�Z�4�& ��LSX���g�<q�!�d:9<�5q��4v��y��Z?\�!�č��b{�M��	�R��фW%�!���}P� �`߇�4M(���G!򄀃=F$`%FP�d�8����ZIV!�A��� Ʈw�y �\%SS!�$������-�-a��7L����R�5�r�!mڹ�lI��y��֬P��D�!��}ɦ�9&ڗ�y
� �D�g�ʁgF` ���!j.�#�"O����Z�<M��$�UW��Y�"O�a����"'K� �C�<o6pI��"Of8{�C�>�j&�<`%pE�7"Oj��b�Ēx{�HE�]�5�Ekc"O�)���\&0�@8����2�`"Oz���ߋ�2��v��	� �r"O:����
)��|Z�#	Q�ؘU"O��q��#ҭ��E%Җh�2"O,���/�`����#�+)$ʬ�C"O���D� �TK���d`p�"O�)sW)��Z��#\K�l�"Oʴ�P�&�>�I��k�`���"OΉ+��ԇX���X�^]�~@BW"O��D�ϯU�����KW3v�� ¡"O����n7����٢#��	b&"Or`z _�
�xE�s��r��a"O���&-L���A��_1R%09"Ob<�'gq�0&j�1��I��"O5�$�B�E]�e*ѹK�}��"O&�xD
N�0i5d�xS��i�"Op�P"i_�1��0��P�'<L�5"OJ��t�V�H�� �%[��§"O�|ђi�"rHhׇ��pҐX�"Oа��C�$���ǔ$��u�0"O<���gÈP����2&�-�x�W"O����
�HO�Ar��W
)��iB"O*���ܧ|X��{��Ü)�X��"O��R%́�#��cg-��#�V�iD"O��qv��B�Ѻ�픛"�d�S"O
d�d&�6��X�M�d.�qW"O5rc�7>l5!���Ѵ(�"OH Z� ˕)��`+2%��[�t�"O��`��8��ph�a�z�Q
d"O������(���OR����"O*��uAH8^�~9��d	�\�R�"ON�"(�;��	t)�._�,5�"Oެ���3�j��'y�.�C3"O|��n�r~���`��;m`Z�@�"OB�+pD�>ڌh9�k^�r�z�""OD�[�N�7'��y��a�t�"O��*���k���U�/b	I6"OȰ!�f�,J�COQ_���V"ONI�S�ޟSs ����g��%"O8���K�{�������|�� �"O0TZ��H�sm����K����"O�%���()���F� 9�(d	P"Or(���f��]��Z�7�P�q"ON`��c�d�YC�k���*V"O]���H$"#j$��l�E�z"O8���ӎ{���I!0�d�a1"O�l�kȗcGb����kYr�qC"O֥�U"���Ait�X?�ũ�"O��{��ѯ2�@,	��̵P�0�"O�;���a�U�� ԛ=A� A@"O$XV�v�� 7�1|���	�"O�`�ǟvg�t�U �V��e1�"O������4C�,��(Ȱ	5�u��"O���#�X�{�����@�&y�D��"Oy#畑 ���'�D� \{ "O.Q�C�Q3
�� �wE�]1֕��"O�9 D_�"����]5x����"On\�g���p�L��N
��"O�FI
�phQ���
Ҥ��4"O� l!pa��	�d ����/��9�"O>�"�[:J�0�"��s��A�"Ox 4
�:|��1uDFb"O8�1�˞I���&��d�)�"O�n�*��Dh3I�����OժD�!��Ƞ@:ݙ�l�j���0��!��Je4���J55�Bu��D�!�ć�?Qr,�g��*�	`d�!�D��V�@кA��"*�j��D�!�dD���1,�!�F��UÁ�_�!�{G��6AN�/^Xj�!�H�!����@�Bd"\�f)`���4�!��V�j��M��-��`p�E/�!�$�L�Pq��C���=;�D�F�!�d��Y� ���
-'��I���P'Oޡ�d�$5�
�p��:}J�`Z�A��y��� i��S��O�]k��i Lӊ�y�Cݽ|#�K�,C�H�ɛ��V0�y(C�nhct䔤R�tH!d��)�y��]1�̀a�ڟ���
����y�%����9�ԥu����D �yb��r�ŋ�'o(D�5��-�y"'S���p�sJ|H���d7�yB�NFP��e�)<m��(�	�yRlZ�r�B6E���!�ϵ��4��'���@eD�1=�A+&Ɛ+lX���'�4��̗�xO޸be'�	r���'�^�J�V�9�rk�/�+�:Uq�'���QmѢG] �td�3
z��'�*B�@"�@�3JC%����'w���fȀP2<�B�+U��(�r�'t�����W�������Y��)q
�'^u;fE�9}�0�K"A�����'��	�n�?w����B��<C,�J�'����a�Т�F�5����'3���@�1��`"6��,&e4p��'��ԁ�Ɍh U��X3�Xx1�'ǾMA&���S�X!*����h
�'֌����+U8Ȑ�tO(u \0
�'�����.Km�D0�	^<t�X�	�'Bh%7��w�pT��9 �D��'p"����X&���#]&Q�;	�':�`E��q�<P6��C�
�
�'Ѹu`Qfխ	e�l��4�\�	�'a�})΄1l��A���W���\�	�'ox9��j�T|ma�\�_���'�x,���	
 W���b�� Pm��'J���e杹��,bả�f��i�'$�����6^����C&'���R�'{�E�biB�{�0��#���P�
�'�B\��c�%#� ujG�H4���@
�'�Ι*�@Z+L%�D!��-#�JiB	�'�xe����b�~l��-ƍ!�P��'"����L�e�h��2l�
eI�':Z��aش"*���e��j	�'l�idA�O���A�0$�i��'��4�P�	��+�F�#@*�@�'�D���Kj�^�"��Dh5��a�'JhH����L�Re[W⑴p����'Lb�"�	qF�]����#��Gy�<aw�'\��UrU'\-p���AFPt�<� ]�L��@��E���m�<�4��0�6i��[0ޘ��#�	f�<�2�����dE��)Nq��hM�<�+w�   �   �  ,  �  �  ,*  u1  	8  "?  eE  �K  �Q  /X  r^  �d  k  _q  �w  ~  W�  ��  ې  �  c�  ��  �  '�  ��  /�  ��  [�  �  J�  ��  A�  ��  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C�>����鞿6�!d��x�^��I��~�!��
�l����v���:�9a��:uZ!�L�,Ƞ�#g��UԀ�e��t�!��v.qc�ʁA�P{U�C-h�!�DD�x>B��cG;c�lK�,��"�ayR�	� Q2���F��u�t��� �/��C�I�Ld֘8����D��T�U�#�fO��=�~bh(e������M?��m���Tg�<� �������T�����R�g��dR"O���ѣi�A	�͖<|l��"O�ȁ�N��SO��µ'�#{u�L�"Oҕ�sGY�>u�0@�'B>]ԕ�b�'I�O 5j����)ɲV�л�"O"}��J]�P#JLa�׊R�Q�֓|��S���O��Ḡ/��l"�88�n�:!�D�	�'X���P��u�҅� D�l7�<��'{���6f-虡4��	.�<�R�'L�Q8�C d� ��욯zA��'a�l�3�F!C����4},0|ϓ�O�4 6g�'���z�h�!�P�R�"O�$Kue��Vrl��MΈӲX�S"O�!X$�ZD��z%��B����C"O:0���b�V�a@���VĪH��I8�\��׆pT����Y)i3	=D�$�&���;�#!a��9��H7D�|��BP���x� 脖~g�T�#5D�H��
�Kh��Fo�Z�s#�'D��)F�^��$H�/ǐ'��(#D�8�\�.V>���bYO�9�4m%D��3"�Pq�f�2P.p���(B��$K
~%x�b1Fb�la�CN�.��C䉮T��[#A�$I����(��AC�C��H�XtN)qH�!!��A��C�IHh,����s�6C K�R�jB�	����#塕��Z����}�B�ɥ~�� 2
?<�[�"��nZ�B�I)&�ĝ[uj	�%��a��;�hC�	�f�-� ���=��d�E۸a� B��;}�܉�e�1(��1��ġ=JB�I�!�\3�oԾ�p��C2h�C�	FxXz�g��dp�Հ	c�C䉇>�6���a9yVa�W�vdlC�	�!2,ҧ�?U�*�����5�0C� XwZp''�q�1c̀�ThfB�I(wM��+����k�I�@�ӽ	LB䉆���F^�=*Q�@GB�	�4�ܵ�!�� (Yv	`s��7�B�	?s�r��d����hj��I(8�C�	�g��d,�(M>�h�h��q��C�	�TTx�5��<�� ��&��C䉿[.� �� �a�P��/ԌV�tC�	3F�!wFY�b �'NV��C�	>=F�m�FǵxZ8U�ց�	tLC�ɦ:�p�n[�u�ҴY�!ӣd�BC�+;���U&�<b��T�@�����C�	<+A����Ǜ �R�I�.ݻs�C䉂Ԫc��T/T.nL���ܴS�B�	->�N�9�N��T]@xËZ�a��B�I�E�Ĭ1� ̮j��� A��'�B�I8[�2�r ͫ���TP�]`tB�$�0C$�!O�偷ƛpuNB��]EdP�o�4'��m
D�ُ9.2B�4$�t(*d�8X�}cRd�+DB䉷L�T���k�2n�i�CE�[SB�ISQji��6��{@��/'�C�	�sϴ�;u
�?�X�:b
��~/�C�I�F!*t��N�:�0�h�-	NzB��<�C��3}"%���CW@B��&`H�ܸ�Ζ)��p��+� .fC�	'�n�x�$t���2�I8�^C䉟2�F�@�╧Nt��q�ŪXtB�I15D�"� 0h},�H���yA�B�)� ��aF�H=�`z�aN�'b��v*O��xc���2�~�0����}��'���� 0����
Wl��*
�'��ԁH>pxcG�o�����'\za�2mF�3��H��ˀ%o�����?)��?����?���?���?Q�=�q���-xpB�ѧ�B�j��9��?i���?���?9��?a���?i�vD�U����;�Pĥ��?P����?A���?���?���?���?q��S�x�+��� &�h	���#OVlI���?���?���?���?���?��j�$X�գ���l�o�d����?a���?���?����?A���?��(b���[tu��+�B�h�J�2��?���?����?���?����?a�I$>�K�m�����Bl����?��?	��?���?i��?��,�lyGm�1��x����n��,���?��?���?���?����?��g�x˷EǂP�C���'�
�C��?����?I���?���?���?�7ⴹW)>��
A�������?	��?����?i��?����?��s��A�N &)*�n_�a ��0��?��?1���?I���?����?a����*��)[�|��� ��r�J��?Y��?���?���?y���?Q�z�(��P��
^CB�ve��A�Z)[��?	���?1��?)��?�c�iC��'�:�i�ƩQ+x��r-dԙt��<A�����0�4)�f����s�P�p��&�:�S�C{~��nӘ��s����9��S�Z�A�u�_�ƚ-��՟�R�(����'Z�	P�?�����uc2&MD+0�ѯs�du�����Of��h�d�Uk�19�A�v�R�q�2�a�����#1!#��L�'Ad��w1���G�[	7��%�ECN��xM9�'$�?O��S�')����4�yR���B�@T@��)T����pM��y�9O�����ў�ş�%�dȌ��#QV5���%`�L�'�'67��-�1O�0�vg��k��Lץ
�ؑ��/�����d�O���u���'|��Gw��Ȃu B�}{�O4�DK�1
>	���I.�?��H�O\�p�n߲iM�:Q�F�Bc�m ��<Y(O���s���$ޑ6��$ѳMyE��uOv�`�ٴX�t-�'f�7-+�i>�ꖉ Q2�8��Q�'�a���o� ��ß@�	�ED�n�q~�=�,��&c�<hJ��~KL,�&ş)���#�|V����p��џ�	џ�Rp�N
W,
��IV�LH*3��oy�u�mIB��Ot���O̓��d^��%D�8Gr��i���Hb�Ʃ<����M��'L�>���O�;5($s �� �h��MM�Kx�S� �>��@jhy`�ьO�ؖ'c(`�C� ��,��D�	H��'/��'�����S��ݴ`� 	�@F��	�/􁻂�D3`.d	�Z�����g}r�i� 	l��tK#�^�p� �G7Y~���D�Uo��m�^~�닥�ܠ��w�'ojk�3=� !e��!'2<)�+�T���O����O���O��$9��b�.Iy�$:?F ���>/�(���՟���9�M�$)Y���dNߦ�'����M��d�di6�ώBb�(CUFN:�ēM���Fu��	]YD�6�7?!g����(� 
����s���?�Jx�$��E�F�$������4���$�OX�$R)�e�5ᛧaU�l�FnUd�$�O�˓Z>��.M�\��'erZ>�05#�+$�����LDA�=�l)?�_���4 ��v
&�?]SGKE!F�:�tB��@¸��4u T0h�I3���|��`�ONd9L>9����IF��Q.2�Ψg�ކ�?a���?����?�|"*O�$o��Zm�U��h�r����L_!h��I�������I��Mc��B�<�4w���E픧��=9� S{$��sǿi��7mC0H+�7�??Ae힧����3��[�j�x���,Ү��qe\
�y�P�L��ܟ���˟(����ܕOΰ5���m��eg��$��XXmq�(x��-�O��d�O����dD٦睈B]�a���q#~-�
ӈh%ډ�	��
O<�|z��0�Ms�'�ص 7���NcHLp���A#��؟'��)�4Ǆş�$�|rW��S��k���FTn��"��6%�Rw�\�������	hy2�{�T�*�OF���O��.���P�C��Ii�r�Э8�����D�O�7��]�'e�:D�P�1R���i�d�	ǟ$#����2U#B|~��O2P��	�x���0'��(e�(ј	h4&ז�"�' �'E�����"�!�3����^�qo6`x3�C���4.G~�S.OBl�l�Ӽ#����Is�y	V�A<e�L��E�]�<���?��i0�a�ia�$�O���WJ���!*�v'z���n�4���2#�F�RUp�O���|����?����?����>4��D�5����LN2,.� )O�o��+�m��ȟ���X�Sȟ��G/�-?�н�d��Y�b�*�(C����I妹��4Sg�����O���H�3U8�UY�� Q�YggI*Ly EY��d�*\�n����*h��Of�(2��2�K�4�X�d��蚘���?	���?���|�+OzUm�
INL�ɺ/?� IRa�8:x(�cC+��H��	6�M#�2$�>��?׵i�\��R�*1ՎQ�G�N��Q3#7��:O`�d>Bf�Z��Vb�	�?��=� vmS��A%1TCV:l5t0s�4O���O6�D�O$���OZ�?ᘡ�.n�Ȉ�ɇ8�Z�#"��Ny��'_F6��+5�)�Or nW�	&P(vă����j�*@M<	���?�'hҰaش��d(<	��E�ϢiR�|
��G{J�#�C*�?�&�,�d�<ͧ�?a��?�U�O�"ߘ8{V�5i���Y�	�?!����������ٟ��I�� �Oh�I���.�J�*��6�&��Oܘ�'R�i��O�S'Y��YA`�<1B,�!!���t�Dy�eo�()ں�s�:?ͧZP��DH���bd��q!�M��1��ɮ�	���?i��?y�Ş��d�ͦ5q���$u��j���v_����+^5A�X��'��7�>�	���pӄ�b��;L��6ʍ[=���EOH��P�4*;r�4��$��X;~���'��5��]�5ɂC�5{��W"���Iuy��'�R�'���'��[>uP�Ɠ�e���QBOϫ�j���gۀ�M�Q�?a���?�H~j�v}��w�"𠱩�
,��(�EC�g�ԵSv�b�v�l��<ɪO1�0�1�}��ɡv�j����W�Jq�偄�qUd�	�js~q��'6H�&�����')n���J�X�����V.TEK��'��'m�Q��"�4h`Bs��?���'�N BT�O9z�*q��@V���i�B&�>Au�i��7�WC�ɤi��9:R�II!b��2
F���*�#ϟ�t�D�|�c��O�D��0��#�d@(5�pBvI�(]�
�c��?1��?���h���$Λ<�f��S�[�8s�Ao҉H���Ϧ�P�B��D��:�Mk��w�t�d��3[˸p�WlI��`�'F�6m�צ5�4}��`�ܴ��Y L�6 ��z�v-c���m��!�@�~���cB7�Ľ<ͧ�?a���?9��?���1]lM)eeA�S3���r�U���dW��M"q�ןX�	ڟ�&?�I2de<��4�E_@�y���إ
��IY.O~�Dr�>]$���[�Ş_4�ځ��o�(M�wӄ#��!���\����B��f�	cy�
�nH����K$t��Y@��f���'zR�'��OL�ɪ�?AE����@g�ż'�� Y��'g�@H  ϟ�a�4��'����?���fk�QθZ�K[vhrYyA-V�2�h��iH��e�X����O�q�d�N�& S�b�ײ�0�����Z>��O&�d�O����OP�d1��R�L0B��7�^	���->t2��'$�ix������?�j�4��7����N�.6�6�`F���\0�x��'��O �Ҥ�i��I	T�{��&L&�`��ǌo�� �p�ؿvn2"Lf�	y�Ob�'�Ɍ�J�4�A()8[P�ԗ���')�ɮ�M{����?A��?9-���(��Ģ|.��S�D�	���8ѐ���/Ot�$g�\$&�ʧ�"�c�X�n-�HA��:G�2�#��D�$�N���"}~�OT��I#z(�'���3V��VT�[r�ϊsjV��V�'sR�'�����O��	��M�1%KmȾ� #Z/��
�!��zF���.OT�l�`��/�Iݟ�w��	[��ٛ!ǆ�}�\E
\🸠�43�pڴ����H��Ÿ����+Z>�$��2�r�U�1�D�	my2�'���'���'��X>�WDF3Ӕ$��,%s@]A����MK����?���?�K~�F!��w�h9c�[	T�V��W!�_wZ����'�2)%��)��+��6k�� ���M�p�!�'аC��б�$r�����#|B�H]�\y�O��Dؼ�p���f��سQ�Y�4��'���'3剸�M���I��?���?�sd��l<dK�C��L�2`C�����'��ꓬ?I��H��'V�Hq*��Z�,ʳ��)+:(	(�O4�ٖ��(J P:`�IN��?`��OF)x$$�3���Ԥ�<�l�`&��O����O*�D�O6�}:��4&Te*��4k�t��0FS!{GR�(��K��f�ɸB�'�J6m3�i޵����u;����$þ���i�j��������;ش�R1޴����(oȤ�'|�8��6?��H���9$i��*v�7���<ͧ�?���?���?���=|&�u�aE�L��%9uFY����Ӧ�1
	�,�	���'?牝T�d-��!V1b(�3���>�P�S�O:�mZ1�M��x��t���k�$	׆��l?�0Y%ˀ��T�aH����Q0�����!"ؒO��.Ɋpk�@��#J�����|���H���?����?��|�/O�oq@v|�I�E
j�!�J�� �VA��ɺ�M3���>����?���i'H����?U�zh!π�(�S2aWd������lA�S!������ld�Beǡ�썣+��H�B4Ot���Op���O�d�O��?���E�`�8����U�3
d��b�Gϟl�I�d�ٴfy ��'�?��i[�'&黳��-������
�i2O�W웦�q��\|6�+?q�ȆD�ШB���3#7�#�윀r���H�O�9;J>�-O��O��d�OĽ `�����)��� ��E�g��OJ�ĩ<�'�i���<��柠�Oz��(�	�H�Ĥ� d�zX��O���'k|6MS��i�S��du�|B�I�Z��"�F6Q��	V'uSB�RS_!��4�P����ָ'?2�h��M�8�h�A�.x��	�'�^Dt�/ƺڂ� ?tI�	�S�~�-Дh"q�A��Q=�P
�e��5<��@�쟃�С��B�ncn���@NR�iX@���HvgĐd<��6错;� Q3�O�R�\� ��e��oP�yh�͹pT<"�̟E�V�Q�'��0��̛���4/���H�B ��A!"��*��Ap�,�8���f��[���,o��kf"O��g�F8�(0_XeX��S���pT&I�c��'v��f�7��ݫd�L�y �E8F�F��q�Ȳ ��k�� ��D�F�[�|��`�`�����N"r��4���Ŭ<a>�F��e�A�!��F|-�FDN&aI?:<z8H!E�bXlaH���-H(5*��.$���%"�K$�� �c�O\uP��� >�6q"D�K�9C6�9Å�O��d�O�,�@:Jy�nW���y[�IG��������X��#E�k���Jg��)�(O�<s��*�� �	�Y�"+$�r���T<E ���9P��a�'Ot�'r�D����?�O~����t�z�c^���´c�:��$K�����?E��'��	�-��`8��`��,�>`����'�'�����
Roâ:�&����O���D��P䊦o�m�R Y`+'4!��թ	<��!�1Bz<�ꡨǽ4!�C&��A��;W Q�pHߋz�!�$�2��|�Df��| ��J�AH�Z�!�d9�Z=K���bg��%��br!�$g��e��m�� L�9�4BƃXh!�$Y�f�T-�5���B�XZt�@�y�!��i���`1�Q�T��
C���,y!�T�{V��%/���P]PP��H!�D�7Ul�@���h����Lև!!�䕘6��B��Q�چс�AJ�r�!��4 Vl�$J(P�x;6�)=�!�ě�a�H�8P�%�9��$�x?!�d�/&�b�F���l��S7@�!��+ێ�(�NA�+"*Q�� �2r�!�d�Q��"U#H�a:(PoZ:9!�$D6~=�UJE�N% Q��՟;!�6NS*���	� �'�n�!�$T�r�p�ra@A���u�<&!�DQ�.o
��'�Z#'���׉�2�!��� �@��A
B9��-Q��|�!�$D<��y	d"F�b�^1"�m՘x�!򤃪q54����YXX��l��r!�ĝ�[�6��GBY��{�K b!�DZ%�X��_�8�x@�%��uK!���*N����(����cӶ28!�"z��Lyˎ��jd��O�_L!��?-h�D� [5G���V!�䃠��(z�SN
}S�f)R!�ď�{��S�'߳7J���Q�T M!�&>�$����
n*�U��O[d!��s�<�)��?t�l�ir��RL!�){z���n�;u�>��Z~�!�$M�17[Q��E��yұ�л�!��g�A��{��I�V�z 衇ȓL��air�O�E���Ƃ�4`�괆ȓJ=�!�*w�x)�JB�d��"O��bR!JZ��݁B%��g}t�KT"Ov����&��)���)���z�"Oh�wM�0�p!��u���(r"OL!	R@>R��a��f١��R�"OvL�7K�e0�����ߘXՊ�s�"O��%� =hV��U�nӪ�2�"O�}x���ј�cW�W�N�V��$"OR�ă��3`ٰ��W�N]�a"O�Ps��ϻT
�#
6`��m�V"O:ԃ0-� &���cJ���[�"Obm��a������#��BGJ�k4!�D��N;��h���)eF��b�>!�d�#"^ �B�B�B �͠���EG!�l���k��W�H̢I�'d�>?!�D��Ji`��Q\�,�QB�?.�!��C7'�8.)v`m�7IM6 ������ i!C$µu�p�n�30���"O��A�a[�F,,l�-C&�nyx"OB�0d��2HL�x3���eې�"O&M f�G0
8���.I�bl�q"O�xcGE�X$A��+�|�"O�ѣ�FG����Q�N-SC�q�"O�B"��@=�H!W#�+vEp"O~���X61���g_�"l��T"O�8I2�й_Z ���'˥����"O��Zu�h�挠��� LN-J"O:��чѧD�9�4i�#7�t��g"O>��C	}_26'Y�<%R�94"O��B��������ܪR��A�"OL���"�=p',ac�Ϗw.c�"O��!��8M�H��/#����"OR,ٗ�qIr��:E~0U��"O�+��"���bg�'5{�LJ�"O����n�S��qq�JE�MD��T"O��
'� 
�Xx)C%'�UI�"O�p���*3`�9Վ��.�Pl��"OD8���܇pI�`9�&��T��*�"O��Y�,���N��e/�g"O�yg"�/v�$�H�#]�*,d��"O|��p�Z�1!i�R��A>�y�"O(	榓�]3&�+rb82�"O��sVk� j�M��K^�K�j��u"O��!��r'��:3Ii����"O���Ǘz�A��s�^(�"O����o"*469 G�HXŪ��C"Oĭj�DI+!����'+�=�S"O���0��zڂ�Y��Y`�y"O�!���>^��)UD�_\]P�"Ob]��HV�+�\y�RC�]�։)"O
�fE$ }B�Ŧe���"�"O���5�V�?�,����Xئ�	 "O��2��������#��9��"O$)ht+�0Vs!���'=���A"OVy@oϦb$ ����A���"O�E�N�`� BfݿK�zE �"OP�A�'8Z�����	�$;PLB�"Oބ2��ԌPW�p8������"O��� �]�%�X�* (V!�@��D"OLb׹�V�ز@��*_�P��t�<A%���}{�ms����"i�4�]G�<9�/�2q���K_=b)x �fQo�<1�4a����ڒ!|�4��Q�<�LT�P,h�!bU�P�:�[��q�<	�	.XP�S��ňb�y�"��q�<a��ݒr�&)X��
�d��f�[l�<�I�7 :fa�k�8���ʑA�<���6N��Q�g��V}�`�+�{}�Rx��	���)a��FF�_�����%8�O������<�N�LѤ0�&mj+1�o�<qS�D�;	�-�DI�D@h(0�KZC�'�rHi�0�k�uc2�1*=
��� �2���O�����G��d$}�ek�.����N�i��O?�ɝDB%�� I(�:X�R�2"�JC�r�($K����
�2#/�0J�$��I�D;�@��$��#��lx��b�ߣRt�Ň�&v<�p���A	��$�\4 ���O���b�(@)*�!�92A�Ѹ'�J�D>�Hr�'IH��'��Ip�/Y!*��E��Oƃ��<ȶC �@=��D\��yr˔;1l`5��D�zH���jS�W7L��&�ņR/>�ZmE#)�M-F��é��9�����S�? ���Q��
/3j80�(�7 rg�i�JX�mV-ǰ>���(�$ً��:O���x�@K؞�Q�aǵR/p ��$��z����Dd~)b����w/v���S����c
�(�b��iH8EDx�	׃H&�����T�9�lyU �4;Sn�b��E�T!�䄑(�� ���L�H��+�l�N��b�/ �' �>���8�pv��~��(�c��*Z�zB�ɜ+~J���Ϩ]�]�Q��(BP6�_�`zZ��R�lCP`\2H�8���I@��%q�$?lO"1K ��d���~h}�1��0��q����7�^��ȓ�$�s��JzX)� -2B���?�AN�Z��H��I֜4�ԑ7'Z�M��L!�Cě�!�d�%/ND�,�$�l��C������թH��b�"~nZ��ҴB6��a�
	+�n�vC�	��`��=%^� ��j�L�@��+��'��xb��U6W�B�`��IM��u1�D\�d0OD���64����*5���r"O�-��/�;l�����!4�)��	�dm���):>@\�a�܄0��IBᏑOb!���u�<�&��?A���z��׬]�����p�=E��4�p�C�\H�I:��N:;�&��s/�x�ph	�K�E�G@]�#�U�'��[D!��=�0�ӗ:=zr�- ;���c�JX������u��6m�p�\��E.k~X��K��^�!��,&I<tXf뚾H��@�d�Iq��H�Ee�D��>���!��Rq�TKc��D�e�*D�<�U�76���ӵ�!.l�`a��tӪ���
LK�S��MKCE�4cBᲖ�l��)Q�Cg�<��Ы-�E #�^�^	�`�g�WN}r$(a6���d��U2QТM�8X@=z���)~4a}��3<��I.���e�Q� ����G;6B�<3ꜰ0&EG	:�i{�Oq�"=�!L�)�?�"�D�.@1C[�t֒��<D��I��J�5�<��Z�G�8T�C�d�4\����w�S��Ms�F	����B�_.Q�Xm���[�<I���-Sr��{ �. ��f�Uy2��p>yA�\�V<��KթH'9bA`D�PN�<iDh�c���#��L0lJ�UN�<A�nX�����*	(�}���J�<yG���'Lx�D�E|�lp@�_E�<�5bz����!b��{�����[�<����m�V)*hj(�S��S�<�Qn��6����'ԦN��Kf��L�<y�Ē�7��r�*�96�飰��l�<�`�ƨ!��I�愜��A�Ġi�<Ap���/�:���J\��xp��l�<�ҦȂ[F����	-[<�ي1̇e�<��f�l͚l8c���j¦?�B�	�nw���#�Y4U�2aCj�i��B�I3&�I$,
�-P���_�`&�C��8c2R��E��x���T!�C��0,-��ȿ4i�ZV�Y0`zC�Aih�@�G��BU���=@C�ɑ*`(�j>>Lr��?��B�I� p���+9�d�x�N�a�B�I��h�;��E<� ��&L��Y�6C�ɷ������( �I�C�	*n͸���e�	^&3C䉁?�b�r�o<!���� 7)לC�	�Yޚy�FK3e�l�h��`��B�I�i8��W�5=���;��B�I�U��Y�v�?A���HԤ��L�\B��`���JgIka4�Ǒ_!X"/$D��� �ϠVbR�gL@%Yܼ���/D��  ��nR5W$V�b��b.Љ��"O���a17U4 �0́�S%�	��"OPi��jY�W�<�d,�?~ZI�Q"O�`�-Ϟ �R��g+�5�@��"Ob4z�,I�U��4
�)Z�3@"OXM�1��X%Z��6� K�l�s�"O��ƒ3>�
���a��I�:��'"Ov$ ��2j���f(s���R�"O��Y�,ʙ�
,1�%�YkX�F"O ��'/̀���CϩR~i�#"O�Yڄ�ޘ\&�\Ygτ' ��sP"O&ܰ�
5Y]\��c"0�&@J*O�S������sV�1�`S�'��񩠄�3�1U���K��XJ�'A��0�*W<@� ���ِ@ 4�
�'ۆ�RO�1`����OH;᎘r
�'BYʴ���V������I,8�ƝS�'�^գr�[�k��Ea��ڢ&@��'�ڙ�D�2<���ϳ~2�!��'����F֟N�,�AY���K�'�R�!B��YD�k�i8~�V�C�'5�y���΂2��ᓢ�Vs1z���'[zDZ*��z49��4l��@P�'چ��g�#+VX�q�[�d����'m
�A�#�~Y�P��,1��`�'W���OA�J|h"��<�x��'͒�R�f 6'Yb��`Ç ���'%��IEOQ������V&��'Ȣ��g �4b8�	�	��}Q<���'8�����'�� J� ��@��X�'#�]s���|��Q�eEm�X=k�'�h̹!a�ڎ�C$�� TT�':���ʃ��,z�i�)i&���'�8��w	�>lܴ�C���̴��'�P\�e-JBg&�h�]:!����
�'�z%�S-S�H����s�ܸ
�'�2�Fn��'�&9�v� .�ab�'-�)S�N�Q�;A��-l�έ��'-´Ҷ�N.@�q`#�ؘ\��\3�'�q+���S�9+��T"?3\���'+n��iNb����8��(C�')�xpi_H�\�h�JP�/a ec�'
,� gV3A{&����(�$�Q�'5���˖8�vDQe�-ml��Y�'�8���"L�``Q�
�����'��2&�Y�2��{B�]�;p��'o���@�6!iQ����*���y	�'���b�# ,M�I0�����I	�'4Zy�AOP*L!z�C��N+9æ��'<�:6�TE u�&��
i�	�':�(g�B! ���R)�]!Ԣ	�'�"I����첢k�,�F���'ў��f�46A�[�&���j
�'A�8*gC�Vݦu
�ψ4#�<z
�',)��	(%)�(���t�9�	�'��XC��O�>	zU�O�X�`S�'$��23H�x��q�����v�����'�xY �#�+�"itO�$�@	��'V�]3�EE���������'���{��& �������"�A:�'�v�9r�
c`�0K����;�' p�AAǌM$��06G�=Z�'����`�pE��b�ŋ�'���	�'$e˓�S�i��%*�iZ���}���� I�F��&v�"�R�P#
�[�"Oj��nC��X�Q-D,u6Mp�"O��V�&���;����"O��R�l�b� ���#h����P"OԚTm�)=�@��bQ������"OP\��&�	]������L�$�D"OV="u��BRx��qC� �����"O ���aֵ���K!�Y�?��Ԛ�"O�@� �ʍRQ��yCAʎ�ĸ�"O�5Xp��_���Q͕�K��ՙ2"O�8��&ڋ��	P���cܤ`��"OJ���gUHD��p��Ы}��X��"O\���])X��-��c�F*a$"O����7
NLm* �_�/�(p1�"O:�!�'vH���l�(V,�4"O,���ۈ	5�pr�˅Mv,��B"O6�K�ʚ20[�l�-ɚG^�l:"O
@1�LD
J��h�U�R�ոd"O�9B��O��KӬ�&8Jص"O�=���L6D�B�"�N5����"Oܘ�@ ��P�N�"F�S"O�l�0N�"��9����I�1��"O$�s�@9jEBT�@�r!^���"OD�r%(T!Cv`u��hs����"O���H�r���P&�V1'�fi�&"O�a�Q��!zZLD��ǈ�A߾��"O|$��K8=�d���۔a���"O�	�#F�h׋�iqL��G"O���piX�R2�I�kÂ>il�0�"O$)Iq���!�/�CGt�JV"O�%#ծM�mBdXc��Qb����"OFk��N�WP� I`�/O�̊�"O��;p'�r�0(ʣ�
 ?@�p�"O��@L�"Q2�[�14��p"O�;3L��(�����:@�y�!"O(x�b��!%��l��0�y�r"O@�5圐i�<���L�;:VFA�P"O"��Sn��`((m	;<h, �"O���af�g�Эj��J�Y"l�"�"O�hT�\10Ą�ɂ��+#"O�l��0W$I�E��P2�"O��t��@�R�3���(��J"O���jLo-������74�,C�"OF(�UGaJX�!Ƣ�C�]r"O��YR�F6�
�i��B(�fd��"OB���cT4(��e9��9æ�w"O�Y.�1%��b"%D�N�Ľv"O���Ǝe�����CM'��H;P"O�i@��Ff��$BɳC�����"ON��ો�V��a2���T�Bh@�"Ot؄��W�yC������"OB�[�d�0 ;�92 �D�g�%��"O�2ri�I��i���oؔ�""O�i
�_��+��@� �|�jW"O
�{&�P1����V��
�0��"O�M	6#�*�N`0��2;�,�!"OtQ�Z/�6����
�Ŗ� �"O&�`1"��.i�gh6�fe) "ON��e�F'U�.�7�¨B��P�6"O������X͊5
C*Řw�40xP"Om9��+�Ui0�_�R�8��s"Of9SV(���-�!� |�"O��*d���P����qm�r��s"O�����4Pz,�r�oΌ��"O� �H���[�^��R�ΎF�!3W"O��Ѧ�;&�
�ٳ�(�����"O�́���P�����b�$�i4"OZd  ���&�9�����F"O��Z5t� ��۵62���"O~���'�uN�� Ê2M0�)�t�'��D��(��h�$ �O�r�=�ȓ;�$	aTd�V�4�PR�6��	��y�Z!�ܬ#R��R��?4"�}�ȓA�ָ-9 a���]�H����aJ4D��u%;\E:��CA]��-c�*O A�T���X�n���n�{���D"O��#6A�JNԥ�$`	�Iѐ��r"O��@���1��(q"�;V'��ا"Oj�:" �>e"͐�A�u
� ��"O�l�r#ʴ<�L1b�<_�	�"Oh	�I:6<f-i㠎�;��u�"O�-�T�Oo�i�f�Y����S"O|ܢ�ˌ5�~��u�ژf�e""O
pA���T�p ���6"O�����K�AA���dR�0g"O�����.���#�N]��r0�W"OFU���&�~�K�B�~Э��"O`T� �B�q �C�CK�"O�T+3)��|�U"M8[��-Y�"ON����.EcDq�
B��d��"O�0儋�R�TÁe�p�ޭS�"O� ;���f�$� ���c���X�"O$H�C��A��U�BM��/N�T�"OJ91$ܤ	��X�ۿD8�x�"O4P9'k�G�������MJN�`"O�IiFg�;D��d�`G�}��"O��@��Ne�%"ǡU
M�*D�Q"O����B����a�����w"O��" = L�Kp/E20��"OVԓ�I�|P�=�)_�Q��"O����Ίd�� TB
:fni�"Oֵ����@�^̸g�@��h"O���CBT�M� �����"O�!�MX-P�fPr�^]�k�"O���D-2rc�V��T��"O��k\/���
�k �5Kd"O��a$��>ܡ���%T��"O�q��b�b�nm�w�[B�4��"ODmQ
������� Q
�I�"Oڬ��@V.`���
T�9�I�@"O��9��\[&@��R�T�D"O^�y�]�+@��A�;Y�0�B"O($�#շqæt���܇��y��"O2aԩ9� 8��BÑ �~���"O���a��Da:�h�n~���D"OxB2��!@������"nl,y�"O� ��n'A|&�BP��P_\�rS"O��>y�bG_>S"��"O*@q"I�l3���#��?I�#"O���R���`��	�m�F��"O��	��̑�nА�핳M5*$�"O����ڦR@m��˕Y n��"O8��`I/M����*��jT@$"O�1�E��d	�
4�J,W�H�+3"Op�P�ˬ�ܘh&��&>�(��"OP�Zq	�Sb;�抣e6&�U"On��g�K�j�BE�P��7��J"O&��螂(�J@/���p���"O� �s���v�F��4�i�<�cD"O�I�$�!0��Q�#G݄}�&�#"OQP#֑��y;�^��:�h"O��[���d}Ԕ��>,$��5"OB):_2L�!��_!:>�0i�]��yr�4͈U����(�l�w�Z?�y��@ld��0拷�쩓VjP�y`����Ҽo��정��$3��	�ȓ"B���R�%"�H���L���ȓ,{r`�3����t`X��_8��ȓ��@cA� �X�w��;�l��ȓdx]p%�C�uH 8�I�b�х� ߆0;AGQ�t�:t҂*R�B����5Z'AV�&d����K7Ji�ȓ˰!�IW��l�Qj7�^Ɇ�b�D�l�!((�֤\
��ȓc��U@�G�t����T�$���m�(!��$C �L��%��(�9�ȓ.�T������`)������ȓ��S�gU9��H�&��[�x�ȓ6̨�cង���Q7-�k}4���POZW�6)F ���F)xp"O���D)BtH��aID�� �q�"O����k�Z	��u)�#j稬82"OR�y�F%S����t� ���"O��p�=c1���ǈ�^����"O޼��-*�� ҡ���\���"OZ���ָU�^�� �ȟ(��͊�"O䰊$j@.K� �ׅ�$�|��"OD�Dm��U��d�#�0�w"O\�`'L��{H�Y�գ�?�Q�"On�Q��؂Y$<�h���;:mA�"Oq�3����}��- �"O~�	@����Lb G�*e~l��3"O���rd�D �{@�P�� P"O*A��OȥoX:�"Q3���C�"O�J�r�X�2�O�����"O$$c��_9>T@��:��4��"O�=��qk������ 8/L�Z"OF��Q�.~�6�!WԌ9(ܼ:a"O&%!����|M"lJD�ۦ$P�T"OjĩE$.A���ظL��|�@"OT|��9MR�b"c��E=L�+�"O�H�񮓯6��H��E;̹B"O�@1�ޚ(��9@,�S'N5��"O���e�9F�ܤS�JX"^�ٻa*O�Y1T	�Kba
���}��y)	�'w�Tѣ�D?8]ڭ�S��<�ޑ��'f"�Ig/њtb-1$E�np\m�
�'&��s ��#w(�f�S�_���	�'d���cԋA��j60T7	C	�'.�C֕B٢������FrB		�'����.�2�r�dK.>���Q�'����6Nͮw�x���S%v��2�'b �����)A��a�NIG�)��'ly�%�ͅs줼S�n�	b�8�'����*)����+�$K	z@��'���H�+�.��8 TI��B6!q�'��@�+<7\��-%A(,E{�'���q�œ?BG����8����'���#��ݵ{�H=+p�X�B���x�'���@�u)���@΃DJ�q�'�j�!C�yG�a[�셞B�ȩ��'���@�ɢL�QcQ\B���S��� �E�$D�yj`�Bc��(xx��{T"OX��a��=3>�)��R!No(��"O@�x��2������MW�@��"O��[�Cѡ}@Uk�$n>T�"O�l@�O��P�����vak "OH��V�c,�c��h��y�"O�CP��c��4�;#���`�"OD���R9"nB��w떈Y|:8�&"O�b�������Z` x�e"O�a2���Y�T�CҨ�!ET��3"O����\����-h1��b�"O�d��	�.�dd�m�
�*p"O�`����tۤ-&�C
�����"O�}���8<pAx ��F�D�6"O440��]3C� GD��3�|�5"O�����DIP��`��d"O��YW��l�a�T�.�xYې"O�����T	�e�3��&\Tlp¥"O4��ꃪn��@�B�F����"O�-�r�W�4������K	1^��z�"O|(�fm��V�6AW�0%4�%"O�R3������!ǰxӈE�c"O������
�z�ՠ�&�F�#"Oj�bs� U�x��o�~��x��"O,�"���>@�$����� ~~e+"O�9�^:(�b�Va3zY��#�"Ob 3eτ�	� a�t�<K$(qQ"O���p K7Z��H�5C��2DT"O��� �E�_R���X6{���X4"OP�+�j]3X*
�`��3��4��"Oh�i]�M���WFP�q�d��"O��B*�)�\�H�l�hH�"O��fhϮ*>,p� <am�5p�"OʱӅ�V'i��J�O�_V�T �"O����2Z|�K � �[�@ �""O2�SƬ�I��`��O�O����7"OfL�UB�%Q�:@1�b@�+����s"O�	*�MVj�q��׋j�޴�@"O�=�e� b��1���_����"O�=��,�%�
�C͂�_��1c"Ot�@`�H���Dk�
�Y""O!12��{����I�y�8��"Or�b�F'uK��qۓh s4��ȓk�����7x���9dN�r
&$�ȓ@)��pm�;���%�г.;~��ȓjhm9�HU�D��Ap�/T��8��ȓr<���ä��F��Y�`e�zهȓ/0��sa�Ia�Qn;ꅇ�&4��(7&M@�	qe�M2*$ҽ��|��}�G��&�z)���O�*��ȓ����9-�)�RŖ=E�r�ȓi�J����o�й�A� �g$��ȓ<$��b��3?`ģ���2#EDՄȓN�B�[��+"��}SU�׬��ȓCe�[G�:]]6�9�_�c\|����BcO�>etT9j���!UVh��#3UA�#�63^<4�H��ȓj��<��@7/8��i��Zk�����a����1LB�m�#$��-f�`������2���`k�9����Ĥ��z"���.а*u���AB������W�L�z�MĆ\ڂ))�-P<Gt��ȓ�����Ȝ�7D�u���� ��@rL3�O	�)�,����Z�D����S�? �4�El^%��1�5�K�
���e"Ojt�7A�3W�<��!�;z�Ѳ"OJ��'B\��i11*�2K��"&"O6�k(^��lC�iY�wH��y��E�D���K�V�"�1D�·�y2N_�B�L(�í[G�,ȓ�'�yR�0�p���DU.	|d&A���yR���P�z�z&�S"}�r�b堆�y".�v��Hۧ�ֺa�]sD@G]�<�al2�ꈚ���.)�]ҥ�}�<�h̰/A��/��p׊��W��a�<���U��h�G�	�t���5��t�<�j�=~J\,�A�Ğ�j4�Wlp�<�d瞽"��#R�v`���p�<�Uf�.>0�B�6^܉�NS�<)`L���z`�Γ[(L�+�Q�<a��	��lɷ%�n0���`NO�<y3�M�i��h塌����eEO�<!�Ay��8���?M�;a!s�<!S!eȆ3���2u�EH�<q#�'LCT�PSU�|�l9��N@�<�VO��ZTȄc�~8Șb��u�<�E�j�����z��0t��t�<᳉S�W��D���]�B=���m�<PB�']Vii�eƉ)�d��c�<Q%1Z����^�t�����A	E�<�w� )�x�	���`*�H�d��e�<�&S2��8ɐkK��4hRi^�<��@��N�t�Cϖ�f4(A�$S�<yeK�Jn6e�o��a�N5��*�t�<�sg�=c�`�'��c�=a�o�<�%�3y�*-�Dτ�6����#��l�<��-C�>Q�JX�n��]�3 �s�<�ӌ�#�P� ��I�tlj�kHU�<a�Ӽp�ذ+��@�1�萫Ӂ�M�<A���O���DD^�v���e�o�<��i%~.�`�ǋ�4{bPk���g�<�v�G8ze:�b���h_^�(�_I�<I���8Z!�ѤX�`+n8xdF�<�P�Q��2����M/��1��-VI�<�nƌ&����큈G� @�Z}�<�7���`9��ˡfQ0+ʰS%B�{�<�1o�D�U�s���P9�9{�k�v�<A�I��8hZh�$��X̮���)WX�<1RK��l���Z2�K�̈���Q�<�⋕{����U��c�:9���U�<y҄�=th�!j�fW��F�`4D�O�<�W�P$b$ք^����aV�^I�<�7�G�*�<0a)�)pnY�BO�D�<��I�6j8t��3J�2�����@�<�3�Bj�zͲ����*M��Dh�~�<)6�" �V��"-ON�!�À|�<YSN�>�V��	ؐ`5>�q�kSz�<��(X�Kyl��ve�"�F�+��vx���'LD+1B���a2U��i��d%O���u�~R�"�ܞ����"O ���A[>��X`�DK�{�La��"O�A7C��}�D���D	U�� ��"Ol��� o|����B�R�|T@�"OВ���3ZJ�h���7x�x��"O&��m��c&Nb�� �"O� 8��� (j�|Ç䒽pC�d(�"O�P)�l\��J��7ߠf���8S"O�,���!���a��3 �LI�"O� ��*w`з,�Ā:�D}�
���"O����Nɼl�������E��S0"O��b OԿ4���a��܆&��9��"O��p� �w[�`��fҼS��=��"O����I��$	h%�랖D~���%"O|�X� ΰZ�� �C
jN؂7"O�9�
S=k����d*�Ch�|P�"On�y���3B�P�Hu��}(��"O~���)œx�.q[�	E�m�"OY8��	,J��PfߋX�e��"O�u��H�(��a�ܳ��("O(�!�&�6�3$�0i�؀��"O����$\���t���;�"O8�ã�+|�L�*���g�2�
�"O@a�vHc|�dC3��|�h�S "O���6![�g삡�$�&���"O���'D_� �WD0A!��z�"OD8�1�Q�!,�TB�$<�L��"O,��^�K��L8�&O�B�09"O~i0D�"�ZX�ͬ%��$�w"Oj�R�k_�
]y��X�U��0�"O��R��9x�t���mI!I���U"ONA[%iEo��t����F�0e�t"O��4��uD��	8*�Ќ+�"O8xp�G�^��uږ�\#�*�J�"O�<kQ�ǒ&����A.^����"O��@4�Z41F��p@R P ]� "O�0J�$��f*T�ϓ.Cab�S"Oz�P��� wΪ��mΝ����"O����ʰ;2�ē��I�߼�1�"O
0��D�5��������c0`��"O���g�dNԴ	0��F'D|�"O��C'��su"�B�Ȑ>E�}���D(LO�YQ#@�	R`���OL�~��pI2"O����\3$I�yXh�f"O>�86��L��xKfΔ�_Z ��"O��p��||<���9iC~�S�"O4��I��"$��l�>O*��� "O21�P(8�rt�LҰ5z�A"O��A"�Y�T��@ ��-qX@Qw"O����홻%�Α)�(�̄$#"O�	� � �BZ�g��d%
�"O�Y�
�8b`XR�o����!��"Oꉺ���BC:IN���uH��|�!�$���`u����={B�h:���!��ğ��q�.T".�=��'_vz�y��'�1O��p�� /�U�5�?pQ���"O,�**��l# �85�I�(J�k'"O�d�D�m7p�����O=D�)g"ODLi��ЗA��UJ�8_�ԡ �"O􈈆!�@�V�����y��"O�LS��J]b���f�lp��I�"O�Jq	�.i�r�`��n=�I矰�	çrwR�Z�!�i[���G"Ht�ȓ]T���\�"�T%#�E]�^h��*�~%��H1DD�q�Ӌ���ȓ?���TJ(
�.�Ag��+�ʐ�ȓI&���C+|���x�$ɉ�p��ȓC@`R��}�"�
 �̯J`��ȓIW��7�LY-��{SL�@�0��NNl�j��2G��	q!I �t��Wԍ���?ٴ4`�%��!��ȓt��k�cUv���OU0�z���}oj�"�拍��S��Lc/Ć�S�? l��5�\?�!J`HYgܽ�"O>% �b|���  IN��"O.���п7҄�SL[8 />�q&"Ox%A�#κ'e�]��N.X&�m�"O0GD�.�t}hւ,X�+�"O< �s�W)�جw��k`b��'"Ou2�o[�\�D)�gU
\U�� "O�Hx�ϋ!V�N�B2G^�{��v"O� R�c��{��P��&U4��"OƝ٠"U,I@ �PB1n+���s"O�����	/6�;�B	_"|��"O��U��,�	إ��9�T�0"O`�S �Bs8���DJA(�"O�e���B�m��|��@�y�n��w"O:�����
.����!J�ē5"O�TA���$�|�*BׄAН�"O��ub�R0�};�@C'�b��"Ov`"�,C�h���@���Je��T"O�<If���%0$X,W�`�)�"O�y{�/�Nr��A<y��t��"OTH���=�l�ʦ8���z`"O�����%�Z� >9ҒU�g"O>�Z�Ǝ�W��@���:�B�2B"O�q�5�[
~�l�o��a�i�"O�P�ii�J��-�t��I��"O2�b��]t��X���M�W"O�6�P�k���z� � h�~���"O�d(	??aDٳ�P>Y�>a��"O��X���(�lh��،s����"O&�vI`; ���"ĥy>�m�"O\����[��<��!ޮN/0��%"Ot�4�/}t�z�� W�HI�4"Ota�s@͔=R�	Ǭ˨#�$�j�"O:�q�횋P�E�ԋO�S5V���"O�t�����Q8�%`*O b���"O��kM��0���2S��0la�|��"O�9J	޷T�
���ac�i��"O
��e��G�ةq���2va\T�"O�Lx�N%t�D0#�֚"�(�"O�,�C�0����b�,I���"O<�āU�A'0�:Adçy�`��p"O2�aɂ�^��[f۷NYf�i�"OȰ��$O�<ĔAS���-��u�g"O�,�B�)�2R#�.��hiw"O�������)�7�U5-��Å\�T�IK�S�O��\@� dB��qgX@+.%`�'���`��оRi�8Х,�=�2uK�'6�=b Nؒh�E��O@��;�'C��bBN�T����\i�'����,�Z����#M��6ܢ�'5����A�.7ɰycE h�|8�'�RAGӏނ	�2�ŚtQ��Z/O@��)�)ʧ�B���ΧYT�\���]1�\��`�L�¢
*(�)��#!�\����Ar&K>C�f0Ɂ��8a��ȓ2�(9w�D3mvI�]�UxL��ȓ7��X�e�.����3O�J�d��ȓ 醨��))}�� b�#4�ȓ|d
2�ġ:L\d�t#�$t��a�����1Vz�@ �I�g;�|�� ���j����Z�.�#���)���0��I�5C�T�S���i�l���.�X@�򇉅n�N��e��%je"T��\����:�� ��"byj%��S�? �y0��]�N���Y��3jq����"O��p��p��pJTA)k@����"Oa�	[�L����t�� \949`'"O%�C21Ը�Ue�8s���"O昀� �i�`h���!H
�"O��i6!)ekL�F�Ն)��
�"O$}�512��C�X�x�"O0	g�<~n���`������'o^��Rl	�<�݈��Z�ER$�'Ђ�Z2�� %��T���U';Ҭ|�
�'�t�ä���P@^�9�
��g�2�:�'�6�P��W������oM�S���'5j\: '�6[\��q@�$��Q
�'8��*EC�#��ps�,��t�U0
�'d�esv#�R*
�1/��a����	�'� 0�	�<Q��a�0h:	{
�'Gb��U����|%i�	ۦg�e�	�'X��+X�jy)��C�k���G��`�<�q&��|�d��̄/ar��w�`�<��0��@��,EK�q��I�Y�<&B��6EtM:3��#u�X}�֭�O�<ɗ��8V��BL��}*ZQ �g�<I4˕�>�`� V�V9�eA�^�<�e-td�(�7��^R~$��+b�<!�9�J���R/k����/�u�<q�gȣg��Z��7��{�TG�<!$M� )J��7�LZ8�q�Jh�<Y��m���郞��u��m�< dY
.���՛v��"���`�<���T�k��xVd�C=h�z���[�<Q5�
6-~B�&����dB5�DP�<	�L���p���_@��r'&
u�<Y"O��'�p��ǖ@�䙥��i�<q���VQ��C!7�v�Y�UJ�<��U�j��J���b�(؋#@I�<���P]�ڔ*��ܲEQh\e�Nx��'?,�(A0�P����L�t��	�'�:(!�*1�^]���L�3 ^H*�'d��j�%�	-�d��p �~���'� ����\�ntc��_6�L�
�'�@�!�d��	�4�i'�F8.�F���'t��%�A!~�J�f*�= >��	�'{���,Y�?�P��2m����t�	���'q�}��-U�{�Z� �jQ��:	�'e<	����%>��������'���R�ѺH�r٣R���߂���'$�+���"K���pO�#un`��'��쁣��
K�2Q����!V����'p�y��B�3d�-��%�* "�xi�'�%Y'h�(@���kR����бr����F&L���qf˚M@l�b	�I�!�d�>w/.�㔦J�tD6�"�d�L�!�@e�Y���8�1��
�g�!�d�Q �%������g�&_[!�$[�9t���_8i�V	��b� 1!�qt�4:TW�U}^�
�AG,# !�<, Q%@�@l�����F�]k!�A!��	�a��wX�m$ �`!�d�SH��3�o�)BFpcc�݌Q!�d0g�QX��@�E�Y��o�?H�!�$�#"�2�ISbB�u�,8�h�%T�!�W�A/�=��مg�j��:&�!�i�jYZ�D�� ����B5�!��Օwa6��2�C�V�z䇔�5�!�� �᳗b��5ߒ0!��	�HQb�"O�-�C��;J^Y��	�6uԴ��|��'`az2݋v,�(j`L#S)p��"`��yr�Q�:���H���`�1�F���ybg�L��Q`��]��0�@�yB�."q�[��A-���k�i��y�ᗃz�%D��y��Q�:�y�ʂ8621��J�=qo�)������OT"~b2���K���"e�,v7LP8RC�K���0=�di�:Pڈ	�"פO�HX�g�G�<q���^4�� ��"���P�B�<�!I�P�8���5x����z�<����r�`�u�H�H�@Tq�<�M˕R1�9C�냒QK��v�R�<q�,:(l�h� �3��0p��IJ��?�	�'6��ɰ��B 56\�^�VA�u�ȓ��h)�EX�k���k��H:l����Q��ab&g�HR<�9@@�l{PU��z�P��J�W�8��c�<@�z���J%`������(����|���ȓA2ĉQ�>&�pR��2�:9��a̓2�B��n��^`�Y�Bl��s���G"�S

��4�֛�Nu��!0ԨC��4A��bG<k?}S��Ò;��C�Ʉ����hU�`�1�6�O��JB��<U���Zf#��)JDK E��
�FB�I�zx�} ��(5v�hn	�c�0B�ɸP�$i���@4A@�j3�\W�ȣ?q��)Zݶ5`��� xr��v&�"�ў\��	�h��@��"��e��Y��H�C�I �ιc�E�K&�� �K7 TLC�I/�␙EH 7L��U�E,N91 C�I8g�ʀ�+n8�%JᏜ�C��2A����w+��G<��iwꎲL$C�I <>�� ��ɿ]R��gE�����d*�)wHh #(��#�8}�"���4B��H !&�����4#�@'��F{���G��U�
e�DBG�������yr��L%��j�W�y�t`���ybAA�.���9C,6�x���OX7�y"�@0\$4������&FB�Q��y�&@j������JG�$B��S��yRf]�l��j��F�@# 9䎏��y�)F-(E�Wh�9d�RC˝0�y2��m`�i��s��1�@ŜpI!����Х2��P�V�����I1!�Ğ0L���A��޼>��qR��#00!��&:b�Kdș�l�8,r�&ײ*!���]U�u���� 
u2L���; q!򤟦j�F)�4k	�+c��g#I�:�!��P�pi�a!�*U^�ab�*�!�DǑP��(qb��o:������~x!�$ԭA�R�z���@1��ի�rh!�D
�\�D�!��*�Ä�
]!�d��aͨ9�����F�I�Ĥ�(p!�d�=�vթ��d' ���eD!�D��=���#���rg�}�g�!�$�'s�ࠃ-H8v�%���!�
*&�4��k��a�@�;!�$#p��0hС,w\���b�5�!�$؈��D[R)��|S��^!�D�^FҥJ�Ê*"T��.� .�!�$X�t�L���iǷR"dU��ݖ{!��DRm �h��jb�\R�� t�!�� F��eG�]��+r�P�BߺQ1�|r�)��;9C|eb����}Ė1B�N�=Pq�B䉡;L~�Kw�Ʌ$����&U�b�rC䉍>�4ɑ�b�h�A�D�h8>C�.6ta@�8W(��2.TD�JB䉳OW0a��O۩b�I��b��H}�C䉬,�%���_ݞ��Ev�C�	�
�n��%#%W��sD����B�	�>�~ɓT���,����H*B�	;��4��1QɢȰaKD�2�bC�	�@|d8b���M�dI� ��B�I���Ű��@�i�((�%!��_HC��> ��`c`�v�(|��e�?@�dC�Ɉ>2|�A���-W�8S��G,Z C�	�1W�0$퍫]]D�d�<;hC�I�_��8UK'Z9\!�w쑝Q��B䉒,M:����O�Y-D�d�B��� ɝ���E(�p�!�"O ܓ2��,Nɮ�	�f���Ca"O������6�L�#��o�ʵ�T"O�:� L�s���9Ab��v�"O`���e(Ǣ ���Y�#%���"O*�����p<x Y���!��`"O��CM�R�.mbBBW~826"O�Up�(��
1 ų�(zYj�٧"O��!��q������qQ��'"O�#��J(lb�j�)?=x@"Oj��GhO����J�wN�Y�"O�d ���+��ݪ���vM��h3"O�%hf���5�6D��M_�>���Kf"O�YKV�-4�Z|a@ύ(%���`#"O�Z�Æ5�pq �����L��y�N�&n��hs�Y�5@00���!�yR%o�U����.��h�Ȕ��yb F���P�X/Q�*�RC���yR�O�ѣߵ7m���n	�?��ȓj�l�۶�?z��}k&ÒGP��ȓ�|��$��5V�I��N�P-�܅ȓ7�*��(�i��튑˓3+¸��ȓsن8��׆G����E΃-�<5�ȓ�|�)�#�R�"!д�]�f�4��ȓ4��3�-�B�}1�ȜHVDH���t���A],�$=c�ѠS�Ņȓ#��Y���I�NRTc����fQN-�ȓ^�b�	�lQ%<�"��p��E�d�ȓE ��
��XP'V�q2� 9x5�����l_&=a�t�ӱn�0ͅȓn{����C��$C�
!���ȓ�T{�瑒2�l��.60\�ȓjt|�gP5
�����pS�p�ȓ)��P����]3�@nRY�ȓ��@���;J�0;#��/hB��ȓ4ƜeK����/�4��Ƣڭf}!�d�20:�k�F�[����E��/!�B�kq"5*����(�@yZ�KM�!򄈱�$�JP�ݯhu�al�	!�d�9mԖ;oO��eHG*	16�!���.-�m�L�$& ��)_�*�!���=,qn�����{|��G�ڟi!�$ܫ,u8�:b�Ѿ���P"�,-!�ǌ�
I�7��<|�4��Вtm!�,:�*qm٧/�|��ʞc!�ɇ;�ҕ+"� B�8Hҩ�<a!��(V�BŨS��X��C��!�� �Ũ�kɚ+b���6�Ӡ8M<MYW"O@-�Eh��GKv9�rG�2נ���"O��i�A�~H�po�����U"O�	���U�� [�+��<��#"OJ���B�x���j�
v�,a3"O�@�D@؎h��p��RchP�@�"O��w�Eb�xDk�K��;^raH�"O9�S��TՖus�HB�~'�u;s"O��kpH�(<8�ၰ�]�I!�I�&"O8-�嬅d_&I"�e��8���Q"O�,[%	� �!�V���H�x�"ON�c�	�vt�aI�0F�p�4"Or�#v�ӸVa�h��4-��P"O��ÀFO7j�qJa��C"`��6"O�\��I�5�~�� H#C�d �"OD5)�(C#a�J�Z�'��{IV1a"O(Y�Ƣ�5b"�e(� `���"OZ�SKX�Z�L�a��Wۖ"O��Վ��!.�"v��=~��Y#"O���G���X*w�3n7\��T"O��B���72h�]��)��J��k"O��ӲSt�&	��(
�cb"O �Y����L�"I�3�^�S�d�QQ"OBM�Ph���)r�ֳ%-|�P$"O���Q��r0Ec��� �|@"O��p�o�!F��Q��["d��"O��sda��%5~�`U,iV��z�"O:	�Ɗ�8�dI�#f����("O
�	���PW
�2a�2��$"OH�J��
3����hI7O����"O�m��LtP�Q�Ι�Ol,�&"O*@� *��@��y��5�"O&�#���u��Y��?�:��"OސZ�I�8=�ԐR1S�c��I�"OJ-r�䇓HV��S�(����[�"OL9�J	�<���sG�$�0x�"OV�@�d��4p�#���hն��D"OPq֬B�G
��T��I-�	Y�"OF�"� �5r�b���fܬӷ"OĴ+$F�f�*B�T�M��z�"OzyX�遛b��+u�����"O�T{�O� ����G1Wt0�"OzH(`�'xl)��_�n>��#"Od��!�3�0�� g��u*��[S"OhI"� #D�p91���h�1ZW"On���V�r�d��hȝ(�vT�"O�]�4��X�,���fٝ~�Dܘ�"O��y��ٿ#.t|ʧˊ;*T:�:"OL�C��,�LT�mְgO��"O��4d���M��,Ǻ2O\Y��"O����W ,D��
C�s���+�"O� ��,DE\d���JT����"O���dE� p ��V��3r5��'U����H�\"8�W焊G.�"�'��;զ� qu.��Z�j�6a��']�E�#�I�h�<qc�� ?\M��'�v�wr��[�a�-B��e��'�V�)�咇�L�iT8<*�Ը�'$f�A򨃤y׬EA��1-��L��'H*�k�j�2Cl8�ʐl��+����'����P N!�00�*Y�[	�'!��8��
/`��2�� :M���'匕�. ����-"R.��"O¨r�'8b@�y��Ǒ
o)�e"O�  �8���a��m�fm��&Er���"O����e�z���8>jZR"O�P��k��t��cf׉G�x��"O$ �g,E5/N���E� ax�"O�Ay"�B�gߞ�sd��RE�@A"O����J��<�h�JtC0JC�Hk "O�T�`E�S�4�b��S>H3a"O�}�� T�D��騐����M���"D��C�`2K������`���3D��ƏZ��H���G�����*3D��4AŏJ�"P�H��K
�Qx4�2D�����/�
Q������B��/D�|����P��e�Z-@g��h �/D��e.ڵh��LcF�� G�4i�f�-D�(y�OZ8<�zq�U#�$��1D���� 12�\�k�`Q(���e,D�$���8z���a�S
����(D���l�|3fK��l[�Hj��!D�����R^¶���%> �����#D���qkA�ل�C�(M1�$����7D�@�#�8q��,
7��:M�����/9D� �5���]���pǆah��9�j7D������%"�̹7�Q]xHqAIb�<�C��4KO����	ژh��嘥�IX�<�dK��d,��tǜQT�MТ�K�<��"Q�l��8fbN�{ɂ��cŖI�<Ag��������ܾ!O�aA1dC�<��fJ9����*��I� !@�A�<���3�xx���]��]� ��t�<��KM�=n	(��X4�셁D��m�<���A?p���8�������`�FA�<��)N�V�nY( ��;H�`Q	�A|�<��סFDv��@!�Y�||q�)t�<���#$WH�PԎZ7w"�9�t��m�<�1d��[z��33��3 ��1��Z_�<i"�Ȗx�bݢ�hX�'>� ��^�<	4N�n.���[�0�3��Z�<y�[58�p0��_�:��SG�Z�<釉*k��ɓH��8\AYcG�X�<1�@~,ze{�Q�Dw �j5�X�<���ԪNS�0� ��&,��i*p�RQ�<���9Ąl��`	";2���b�<���-�*ɂ��8�(��Da�<���V:v�N"���\���`�r�<Q��U�=@!�R/�G1T<��cIo�<�SfX1_�t��$�!��aE-Hl�<yA��2"�h]�Sh���ܙз�A�<A($E�JT�6���9>�Ҩ�t�<9�!�0Ĭ���}%�蔌Ae�<p$�(taPo�WR�YHԯ�c�<q�j��?]d�!@��8�#��Ut�<QuCM/xn�:����B׸ZrBنȓ4A�¯T�$E��Gɝ���ц�=�����m����F�%*��݇�i��A��HE����b�j}��S�������HT�֖�<�ȓ�X}ÄK�.��V�ۑ ����ȓa�B���i	�z��ro��\&���ȓ��\@�ΐK��岷�P����ȓ@�~-��%P��Ja�R%�"���J+ � �\�6��cI 3x ń�L����L�#�&� ֹb�&�ȓm���Q(�7y��<�Ңa!2kKG�<!���ް���ܸa�rQ
��<� L�3��\�N�6�0���
@�*���"O�\	��T!'wv=�6�S�-甬��"O���T<B���$I;ֲ��"O�qQ����.�4 �Ï�K�=C"O��S a]�`}�QJ������"O�}�qg��H��t�#m^5k�F�Q"Oh�86C+%B��*BϳYE<0��"O`hHa�F+M��G��� >rX"O��y�,rI�.�'6,�B�"OPu��G&��{�C����"O�8R��< ���C /��&�T�`""O��JtL�QJ���sC�i�B��"O���F!DV��1)�!A3i��
�"O\�`5䔉S��d�b��A�t�Z"O`D�s�  �<�#Qg*��"O�}���C�OϞ���AF
\T�aP�"O�:iƲi��˳.[�L��\Z�"O,����
U_�di D,�άZ0"O41{7��=h��\�v��+M�����"O����'ބX*:l�R@7nLMB�"O���P�#"�pCD.O�@�az�"Ok�*�T ���,�(`� �"O�0S�쀑*���l�)!��3F"O@}:�����(�j�"�X��"OZ�{n
'?�D��3�:���z"On��T�X�M��<�2�H*�ZA� "O\T(&��OA��îP�sr��8""O��	P�Ln"J\���> ~�L�!"O��j�WfT4 �/�Cw���"O��	h�d�d��\q@��"Ov�{�l��б��o´e"O���)X�G,d��&�ΟCC�i	�"O� :RO�@_,q�Ǌ)d#*�Ї"Ojh��Ę��M�G�;��ӕ"O��r��l6��@O,�� �"O
LP��e�<D@��O�I:6�"O45Ѕ,g�	�1@\! ��� "O�@yU&
=�H�6	C%-�ŉ�"O�P�M�8 (�k��L�G����yB 	�{��k&n�>i�ⳇ���yL:Q�V�X�M)`�@����8�y��\+%�\���]A�q9Gj΍�y�/���>4`#.�V�����n�'�y�aĘx�����B�K^b}���y�MG<l��ٺ����7 ���ì�yB.S�"`~m�2�A�'^h(B��y�c�Jp �V�ܣ@�)�w`Q�y�˓X�|�`*i囶D\�y2+����`kC�HfB(�	?�y�cͷSF���$B�\�������y"hZs��86G�4Qh�$(6��y���2%1ܵYV��Q��p���y�D�PY��1q�F:r0���ǋ ��yr��pv�`�G�ΘcH�j���y�n�+����_�	�V�CF�Ȱ�y��4y\!��/�t 􀸶�ِ�y��V!+,���M(�j�UHO��yR�2�ޙ����M��0(O��yr�ɥn0�2 �ģ%6 �CJ�y�I��P�yO��V�@�P��y�ؖ6�je����V�V�IQ��?�yr�S%{�x���Fz̈��C��8�y"F'F<�d��	ۛx��+�Ɛ��yBoW��ָj ��s��Њ��[��y
� �9A���lm(�"R�75�V"O���b�
\�e!���/2���"O P�2��3������y0 ��D"O�J��U>/N���2,T��c"OB0"|P�8�I�$�����"O.�#%L9y쑢�a�x�� p�"O"u�"	�W��qb�5f���""O �Y)P</�\���}`U�B"OT�p$Ӯ$T���Hp]�I�7"OB�2U(�/3	t�1g(��L�j"OĄp�GN%���7�˟i�(�"O�dQ�\�D�P$8���&DX�0"ON`���ȈR�l%���q��� "Oੁ���%'���jg-��z~�s"O�{Ť�.+bR���KN	�\�
�"O���`�ܠ���{Ɗ��z�|�;g"O��C��;a���ĩT��8�"O��ZNV�IE�u�%�{{4�@"O����!��K���7@Y�0��"Ot��gM���9cK�J����"Or�#��V$��8;q�V�}��0�"O��&�Ӫ}5��@C����"O�qɢ+��f��t��*x�Q�"O:ɚ��W*o&�!8!�Nr^� "O&��1���&�����4�>��"Ot�A���BA"�3�6A�P�"O�嫓A�[�������s�T�a!"O�$v`P�Fm�`.������"ONi��j˧y�Vŉ0(�Q��p�"OҔ�1?hd��'H�&v�>��"Oր�F��Z�z�S�蝰0���C�"O�)���eu��*��|�bT"O^��1�[>Z�X���*P���Ec`"O�`���JL�� 8n��L a"O�<�F���F���j�3�(�!"O���AG^�Wc�ˡIǊ6�h	�2"O&AP��
.mP�9 k^�t�5��"O�%�����[;~490����z-�g"O��cqA�p$�8'`�=,����P"O��`�T�=~~�#�nWC�DP�"Ox"�Ƴ&�RkI� ��U�7"O|H��	�	:�t�8SJ<~|yb�"O�p��4,Y(,@�	���is�"O^��6�I-�b��k�}��	� "ObyQ-S2�$M�$
S,���0"OD����u�Р 	� Y����"O�@Q�NݮQ�ҡ��D�B��<�"O$��ڸ|}�Y	Ą�	c�p
�"Ovc�Z�l~�	w�E�Z��"O��fa׺n\��P� 
4O�a��"Ob!K�����\4�y$y��"O>��W�(6P-0�ȊA#x�f"O��z5O��[�����Q�D+S"O��b��w�y1�/� �@���"OH� э~��Y�Go�?^@���"O�!Aō�O↼��]�r��"O"{��&�`���];(7�՘�"O�A�@��s�j� �_A�yj�"O���򥗦#��Q�DH�[2�]+�"OΨ`A��!%��1BÒ�*x��5"O�!���#J�	�C�
����"OV)FL�0��8CU���V^�:�"O8�Yp-߰� ���r��P�"O�-�T�:���m��b����5"O� �HqQ(�9k0�qZ��	:�i�"O0���MW�t>�JCM�c��MXV"O�T�b��(7>�k1�,	�h���"Oҵ��ӅFO�(
�㕋\�} "OjD�r���h7��եL�"�@u�a"O"i�'(�6ڪ��n[3qў���"OV}sv��;Nn�ڱ��:�0�{ "O�,�iب%\�x �g�?,���"OD��iG�$`kw��W�PH�E"O�9�B�^�&!A�A�n�Ka"O�� �@C�$���o�RO��"O�i����0Ce����hs�h�+2"O2��(R�~�Aᐭ�7ۜ`h�"O�A�� �Q��{b���(��"OT:�ё'���b�k�;y�0��"OP	D�Gˎ�h7J��pLu��"Oz��fI�B�L����Q �}��"O�I���c�� �bIV�:�Y�"O>\[Q��`�~1�*G�V��tڤ"O���҉DN��3�*K`aZ	��"O4ub��ǡH&�E�C�ܿ(�
y�"O.��5/ ,:��S�³T�|�zU"O�ɲ �T�]��K3Q��"O,� ���BG�:UdM��㛝M�!��Q�e�)��2<r����!����,bqgI�V"�9�UA@�)�!�@�z�����."�<�QV�\�fF!�"sr0	WE�e��A���&,!򤜎T�,$k��#LlZM�$D�h!�DTi�ɻҨ-u0t@�c	�o!�d���F%�G�!~�(p-�u�!�:��I㋚�$��ݘ
�!��A6x4,�td��tm����2U�!�DK(\1���1�����	J�!�ė*U 	��ᕗ^Ķ8���e�!�D�&�2- '�C�0f%��i��=�!�$��UL!Pc�{�|��)���PyR(�2hX�Ls���oVZt[b��y�K�-Ҥ8���� ^����� ��yҌ�/KW��Ӂ�#Y1Q�R���yBۭ�jԙ1#���^yyb����y�o�(x�F�TjW0��bsB�y	�=P���&��7b�R�U>�y�BϏ3�>Գ��.�@�����3�y��G�^�����J�z1�ᐅ�y�N0
0ir�Q�t�0�
�����y¥A-G_�e�Ǔ�@jU"����yR���Mn]�蕊����m�y�	�n�nDj��T�xϪt�&����y�D,K n0��_��iㅅ���C�ɳ;6+o]J"����=М��'����,��;Q(pk0���a<�-��'~�y���[= ( R�l�V9�
�'V�=J�a���5c�
QǬ8��'��i���0�����J�n{�'�:��@4I�5�ț1�3
�'�̜ia ʔa�j�3%A>�L83	�'�� �/3����`K?Nꈫ�'�j�b�ǚ�a"� ���=X���
�'X��j�>��P)�$��|h����'� �çh(}�|���ʿ��9�'��X�Gc�"<� �@Ջ,%@��6�\,0��
v{R�{WFMx�t���A�S.Ze������
9Tԅ�S�? ��� P03�V�Y�ʥ~ȢD"O�]Y�>Cf�="ֆ�,��9q"O�U�d�'4Z����W��aI�"O~�fiH�A�����?4V$�aG"O|qiT��~l�Y�D��)@v�&"O�(�F�2*��lY���
GL
��*O�Е��h�\�2!�����
�' t�Ϙ�Bb�R�G���{�'�F5���TG+���Wn�D��EH�'@h�ȝ2�}�PKM�oԎu��'�㍐�j���V���a�L@�'t��S���0�^/X�ੇ�=�z܉A��_�� 9�)̓\8���ȓe�ĳ��ݑl�<J7�&k}� ��H��} Ǭ�?+�.4HS��1$���JO�(ɥE�a���a! �B�)��{�kƎ��@��F(��v� �ȓ:7I�D)?Ρ�lV�3���N���9�+� +�6\ G�
ݜ���7}���O	�AA,�Ud!��@$��H��|�ׯ�*���`�ް�B�É�h-@�={��ȓz�� ��2N��ȓ4�K�7,�i�ȓ'>�X��&�.��P�7�(I�ȓ/�,�:6ףg���#w,ӈD��H��#;�8�V�ɲA�sá�WFE�ȓ$���FB��>~l�ȓ%�RE�wk��t����@&ي4 F�ȓ#\ �#/T�� ��ʚ�=�޸��M��Sv�- #���Eك&�0��ȓ2�b����]�Hf@�k�ޣ:'t-��TT��2���@�"mN�ϪلȓdN��'e�6)D��B`��n�<�ȓV�Py2�@%њ��Z�&X�ȓV���H䀅'��⡦Bv�&��ȓ@&��e�
�E��D�ԅ�i�b̈́ȓ���[��U�vפy+D��a��M��wܱ����	x�����	�lhD-�ȓ6��zRh�i&P�
)���ȓ����ȉ�>�d�'AZ�!��l�ȓq������7�PAx�aF �q�ȓo���qM�4i`�mȥU�VT�ȓs�FH�ŬC�[��҃�|�p��PU�U����%�ԉ�K�(�ȓ{EN��Bo�%����b�ԅ<�@�ȓ?��p��/�aB
09!� �:����z^e���pNl�(G�P�V��ȓq�0 #Տע4�����]�@���$����
�$�3�mQ�6�����7,.�P gC�:� � �f	�Wo���:Z�x;�� "
�@1@��ދJ��I��t��a%�{�8 `�/e���ȓK��1����>�\ccL�S����,�Ry����9j\�����[X�L��x����#��<1ؔ�#B�ftZy��g6��glD�&�����iiL��ȓL��-��I$;�2��ӧ�1H�8<�ȓ8��,�&m]9Y��{7鋖Tr�<�ȓ�|#��=R~�!��̝'��)��&x��&kϛ�n	i���7��ņ�jb(W�q��_`���ȓD�\�����	KO��	�J��XXY�ȓ|A�X�&
(	r�
DK�+TH��g���c��d���"�)NC�)� H�Cdin���ʇ@ƚa"���"OxM�E&Z���ŠL y�]�"O�|�7��.z�`�`�C���"O�4� \�s��Rn���"O�M���źdp*����>/YĒ"O(L@�o%r*TYc��.K��j"O���w)w� �	��ݕvWʬS�"O��	��6z�Ljn,(3Rp��"O��4�_0}yJ�X�M�]�"Op��ԨV�7�6 ��
���K�"Oxx���ʤ��"C�<d��d�v"O�XS� /;r��t�RHan�b�"O��0�zD@����8b�����"Oha�7ʀr��Q��c�5�Ї"O��3p)�	>��V��	v6�2A"O�y豍ƓEk"���HT�kKr<k"O
��玨~Z2&� K,�%�"O:\ZB��	={$��"&�D� "O̫�Gk1P���n�"1l��'"Ov� Í�}2���  y�^��"O
E�I\�p�|�R�"�2p��"O�0�@D���u�P�z|B�"Od�����#���`�\�
���1"O������%ML���-�f�D�0"O�����\�f`C�e
�Ph}3v"O��a�!�5[�$5�%���d�K"O���E�B�\8:�8�ҮO�!��� �zQT�V�mN�ř��%$�!��6i�5`%ɔ*Lڑ�"��M!�dC-!6h`�2�*���nĊP�!�$Y�5�x���VϜ|㴇��^$!���(<"���`�8
�E��G�T!�H*o�j� Ì^�;��<��Ǖ�b!�7O�h��bV��zi�A�p"!�D��]�p!�H����$�s!�d�#=��;EF��U�8�p��K8	!��?%J�ɷ&��tg���虄n�!򤁯7-��!c�X���>�!�D�hC��#���4 �y/Z�(�!�$�	��k���s�t�I�!򄍧.0�Ei�A�cj�� ��^�!�$�2]��C�MV2HR��s�σ1�!�� �aN"��$GW?�퓐CE��!�dI�H��!��ܣqB�I�#�g�!򤅧\��тӮ0W��%¡��+8�!�dMH&�2'�
�Z2U� L�n~!��֋	xt�b�C�ww��(p�$2w!�dC����PWIi�X� �H�,w!�$I�"�z�x�	 R�X-�al!���Ȥl��#����'[H!�䝬=��q�m72�P�0�O��x-!�$��j3���B�� B��j�<��N��k�ŉ�f�:��.���ȓu�������r1��+~�*�ȓ%[.C��(�D�"� *-�`���th8�J�˘�f:�*��@?9C���A��=+�F�9ڎ���7T�B5��@�R�����Vd$�+pV����dUf0���9�0L����N�ܥ��-�d�t�ӇWv��ۤ@X��2-�� �@@�gI�L�J�I*�LV��ȓ ~J��R7U^�9䞼����a�L1�`�-���r�ݠe�\��
��j �øG���j�"^��Ȇ�S�? �=���� w��\��:��(�"Ol� ��;gj��#Oэ�&�P�"O�"UA���r�C��|���"OPD���� 6)2���U�4�A2�"OD��@/]"<�"��6�ˏ1 �ʴ"OH�yA�L�$��f#��B2 !�"Ol96(}�2���#M�� 
�"OZqɠeF�9��[�,ܪ#�jK�"O��d����h7&^9!U�
�"O��"���ifB������K`�rS"O2�$K^'1����}B^��"O���G&@=����±)b !�"Oz�
r��x<��q��f	l`��"O�bk@�^�na����,*��9�#"O��ؑ��d)�B����t��f"Of��5�Y��`���#*yXa���?D�h�@A�$*�h�3i�.-� K*D�\���5�p'ҝ)�6��'�&D��R��EN=���c�ì�(��!D� �Ѕ�g���BGhB5����!�>D��:gA�OLT�DdV�U���
P�;D� ��	�&gP�C�O<B�\M���9D��Z�/�ѸT;� �<�~�h@�8D�:��ߣP�^�q"��*v�p��G<D� ��IC�s��$("����<���$D��+�AE� t��(ǥh��z�f8D��s���S���s�:Fx�p�#<D����L�S5AH�o��&����9D�<2'$�D��D�����b%D��i2�H^%���G� �ɤ���7D�H3R����V ��L� px]�0�4D�ء�ر�6m�#I�>f9�w�0D�P��G k 0�	F������;D�����y]�ah�1V���$.D���Ȃ�Nd:|��aA>�d[!� D���C�� k�@q�dA�ckhQ$T��r@�Ymmh�9�-Q��8�a�"O�]��m�C�*�@&�E<�0���"O�<�o�&L�B�KS%˹8c,��'�(]"�b�-V��a#�P'iL �����!����-�4>htER�H !�!�D�3/�DC��|G0A26#�1�!��V�^&Д[�͟mMLu �i�){!�G�����z$vx�&�H�!�1 ɡbә�4��!�DK0~9N��A�ث6-��A����!�D��
,+wl�,SPa����9�!���k�"urF�	�L	�d��6*!��XlN�SQ!c�h(i��W!��6庵�d!F�p�^�z��Y,d�!�dS
��[rW<���H�H�+�!�䚥N�z�'$?G|$�A�Q�!�D�?C��C�,Ɲ!�����a��!�d�-#:����-(ʮd��C�:+�!��$An�ȃ [1{�����Q/Za!��W�/B00n m����!nİv�!����=D*�"��7(�����!���z��9yu���������5�!�$FzN�M2q�I.W4%y�ϑ�
L!�ė-'�.)����AD!��	�'�����ԬM"�p�"a��R �3�'�����"v��e�"k�U5����'pԁG:=���AG�ZM$�ϓ<��ag�V��D&y���$	�e'��Q
�qs!�d�?0�����=s�ء�j_�1��'x�\���?	`��� ¤��.�b��tp�f�{�2�Yr"Oڸ�j�((4�
��t��SPbͺ)�B�,�(�9�`$�3��ۗ{2QU�?MH��A��T�E�!���y��2�PR�x�yeÉ�A|Z�:˚� �5�XX��(")�4�HX��G!F��ط�(�l�ttᥓ�A]�)��jb7Ÿ;��@�0�2. }x�!p�<9Dh4`h`����`�sy�ᙇwPh�#'���i\
���(���sM�x��9�!��8yg�`X�kA801�EC��(u� ���
���3#޵Wq
�:�Y>�<�Q���ű@��+��Lkc�UHX����F�0F�ɓ	�6�]%
֣�x�Z�I[���0[@y9E�Vc8�:F��� �n{��!��Q�$�q`P�3|4��Q`D*it�=�Q ����ƅ�m�}��K�+�aҴ�y�X��z5:Ƨ�
���!3���I�"`{T�	1	Q=Lxu r�l��ygA�h�(y��צ�~Ma�.�yb�Fo���*�e�}����BX+�|���kX*AP��W��2$��Z��o���Fy�D_P��\k K�pǾM9ҀS���=GL�'.�7$��U�:A����v2Z��Р�bt���]ݮMr ��a8�	�g��ed���tn�uK�����;�I�Rq�U{�F�����3	�j��0;5G�?�°"�m�:I��ƑP�qҮ<D�4J ��p���I�MK!>�ٳAi\����bg�C֪(��iѾ��-j ������@ߙHY䵰"�=4$Q�4�w�<!�.Ҫ�q�#j׉(���g�֮$�6����P>�h�����-{�r�"�Nҫ|��<YքR-xh y&��z�Z�*���i��L�QC�������M�P|+��c@��'�Q�]�p���4U�"\s���:�p>��	7�8�RM��-:2�ã�b�ũaϐ�H��6	U�o�"X�a��I�qQV0I���6y�W���!�$�1\���C�e�,�p�E�H��<�%�^�SU|��2�M�qU�U��0��O�*��;�Z�����8����ɞ:
8D�ȓ|���Y��Cf�\�RaB:q�,1�7)I��* �)�.0�K��ӡ|���aP�"ʓj� qK��ͥYIH�yb��9b+�!���j�|��.��c���JTMA0m~�����<C�(h��
f� �vN�-ւ!��"\X���6nA:�I����	�=�h��K�<�r�F�v�m3� N���謟FAY�R$���@g�6#���D"Opzt�})�!�0+O8�a��v�|  �'��)��D�0@�P�J'§�V��MXa�c�#d�n�(p���6L^C��-�h=�#$��$�nM��4��l�R��=E�s�5-�֘`n�ٺ���N�.:V����#'	P��ӟ��{� ��wj2�9�M�,9��D.� !=�A��@��.A��c��,A�	
�� l ���(��Aѩǒ8Kh	Ex2�-#�hɑ"����Xgh�����ah��oOЄ�B"OH��&j�>���Q��V�{OF�T��)m�2��͍���S��?tR�5�Y[G�\�VM���Kv�<�R��98�N� �EXr��f�p�<9�*ÈJ��X��A��\1AM�q�<3�ސ[�����QQ�t�E�n�<��k=\��)�i�?�`��RC�o�<IM]���yqh���e�A%�d�<��+7~��W&�*8���Dz�<y�	;m��*%a��e�E��`�v�<i����j��+V�!xvB�P��]l�<��Y$n�: a2M�"X��U�� �D�<1ǌ�'ǘ��T	�=��9�	_A�<A�L��:�F�R��W��ܼ�F�B�<S�ױt!��0r ��4�L��M�{�<�Ģ��d�!�Αei>�C7/JL�<�CG�*F1��޽r�4"� O�<q���6eFua����%˕@�l�<��\5?���WI���T[���T�<9�+��d�0�`ې'��H����<9@�ǈg�(�b�ě�88E  ��m�<ѵ$��t�)�:F��DX#��j�<	3���Nu���7�B0MZ ��De�<	�f��$���� �,.�n��i�D�<� �LsE��L����_$~E�T�"O�(Bp�ߡ}��;uF�"x>��HT"O�,)����r�`[�f;7��@��"OS�%�7임 �ޯ*����"O�ڲ�!H�<٧ٕ(�� !�"O.�f�A`�
A��#�R��Pq"Ol�b��9:�c����SV��"OB���N�3�hX�!\�.F����"O�Yє�P�_r�Y:�[�i� �"O�EZeH�3~� U²�4@G��92"O�@��·W���B��A����"Op�ۢ͑(`�,U��ѓ\���"O4|�r��$?,�1׫�3d����"Od�I2j��c�RA�F�D���U�G"OT$��
k皔 @�PZ�0Y��"OLU��ɉ1�$�YBW.(`ڒ"O2�[G�܁`�H�(�s���e"Onњ���b�CF�ߠ��D�U"O�U�����ؚE�<1����"O�$3�ț����yb�5�mk@"O�P�ԯ�'���!�G��d4�@� "O2,���8�}k�� �"��"O�Rab�,C"���1�
��F"OX��Ī$:>D��d�=gPI��"O|l�w���Lu�����ˉqH��;�"O���M�:5�Z�{� Y8O�ܰR"O������>Yu����τ�s4d��"O��yc�A�[(1*M��f?��T"OԠ��9K����퐮z� "O�<��"]3\�j�P5LK.�IY�"ORLr�Z��Y��k�#1^`���"Oh���"3hȹ�)!p>zź "O,Mkp��.%�V��F9Ctp��"OJ�R� �v�����G�ok��3"Oƅ�.7DQ���Z=�0xg"O ����?10�V�J�L"�["O�t ���[�$���&חV���"O�TYюW2*h6YJL[��"O~���Ht����#*�=	�:��F��'w٪�ڍ�	�Kd�)c	;D��1�HٲJ!�d�=j�����˵ l*p��ԁ24@ѻ��I?��gl�|�'�$!Ă�V�`˅EA]3���'@tB�eV�X_��4�I:W���b2j�E\n5��刡LA����	�`���!�9yYDT�%�խZ���d�*r񺜀D� *Y��ۖ L�.�![��P�4���0�l��*���!��ېI$
���F��f�'�$�G��	<"ђG��3t4�F��)Pu��h�+��nO<�Ò��1�yBh�X�vq�F*��t��1�&�U�x��8�厗�n�t�CG���i6P����L>��n�Mc��i�%�v5D"�(<i��n�|P��B�p�9g���Sa���&��pҘ�`T·�q%���G1�������!,�!��Φ/�axR�ߦ<� �(�mX�z~$])��a� �`�T��h���� �̵!�Orh6Ι	\͜-JT眄wU¬�Ɲ�<C�N8澨9��H��!���s���xAAaKG�]0��IH�~x`݆ȓu�HCu@Ŋ-�b�&�Qq�A:7K�7R@�ಯ֟[k��(�G�f�'��.Gf���EW$B\F5y���KV��.Dn���*݌?�n1�`�S�6���X�����C� =(5QC	��<���(D�`��ƥC�u`tp�Bs�$�F�6*��kC#��w*��ʳ'��w�u�%�]�
�ڡ��-��\�Ɠi�0�#f�\��%���R4cS���'���cDMZ�m;D!�m^]dΜ ���L�`��� ������	4�!�$�T���x��`�
t��(q�dG�Q��!��0LƠXLC1�ĒO�`��iP�l(��u�$=�0
O4]�$"��v��9�J'�%��^�8
�c�N���0=� �PB0��=`��ls ��6��@���'���
�A9��T�sF-����4�Aa!�;{V\[�H�I�<��g��&�h�Rp�7
-$��M�ɃoR\v%[�}����$^m�Ojd�d攈c���6L:f�����'�(9�Ĩ	��`��Mv�6*ҒEJ�b������ � ���ē� ��슰(�@�"^sBh�Ɠ�*y��	��.u���ՐEi�y���R�yԒ0
щ��
�Z��䒠pL��/�I%z3v�zr�z�#�	�Y����<�g+R�X��<AR� ~HiR!��Z�<� 
:>��T ���,��g@J��@�c!�v��d�!(�B\8��^�y��.�>�I�)Cy�~5`��ѻ_y���ȓw�@��"{���×0*k\ ��_��c�"�$h�"��%l��<�ȓR5B�+�)n�+-"n�`�Q�"O��rA�I&��óLs˜u:&"O�ѡ��՗r�`Q豮[�w����"O����D�?C�Z�;6�]<��m�T"O(��q�Uk8�R%�
2����"O�)�'f��lF��&*B�*�,1�d"O2p� �(�X��P���w�1�P"O��%�47�`1C�,B
M
2,��"O�tt�2T����A��q�	
v"O �Y&k�<������&h�Q"O�)3a�)Q6`	aC/�zeb=��"O4%����302�{�,�#zEΉ�q"OdS�l�s$r)c녂G���kG"O�p�����*zpu�j�8st��[ "O�}Y7Q��R��d�Ot֥�W"O�̓���o0~e�`�!P�D���"Or�C�ʁ)M��l�� ��p�Cp"O�q1�
�z᎜c�H� dy�xr"O��8hB�о����/fb��"O�a��SC�F�pǫۏXfN<��"Oΰ��a�;%���bQD���� ��"O����C�h�:T+vĞ�[�z%�V"O��r�N�0��X�	Q�a��8�F"O,��r`�#k����ȗ~���f"O�u�VC�;pF���7a^}��"O 9���t�Q��V	)g�ċ�"O2|�2%�Z�8k�)��at����"O�EPT�D�MZ�И�'6P�{�"O*�s#�V�O�u��ѯd����"O�,Z�M�:\�,p�Z8iT^Lq "Oԉ�c�����r�.��N_Z4��"OvuZq� wƴ�'��%ʐF"O��!ਛ/n6\X��ſP �q�"O�]�Q �4	N�� �M�[���4"O|�
GEU�lf�8�ϳy |T"O���I�W���J�&ů\QFy
A"Oh���zҥ�g�[=*�b�"OP)CD�B�iu�\�a/y*�$��"O�cg���>���J�oT
P��"O���P�Φ0��уM�7
�4��"O JN҉�6�Q��D��.�"O^�8�V�Z( @8t��ag���g"Of�7`�*�`�)���W���4*O6����ܱv���
�V�s��1�'e���C�	���cϝ	�f�S�'E��1A`ʐy;Z��1fye����'�Lِ�cwJ��PPѱ$���z�'�81j��p��m G�A;���'��cƊ	#JR�0:'@";�$�H�'|~�DI*%R2��fG?�h4I	��� R�Jt*R�|.DT0&�,)c!y7"O�)�k��v=5��C�?ri�t��'<=��׿��	%I�.IC1�O	6xձ��� C�I=7 ��R_"�8M42[�O@�ib��jg�t��Ef*�0�g��p�y�o��g?�B䉺�Tͩ�)�?H<|9� iU�(}��Cq.U\~�a�+W�T�}&��W(��'���"�1g�h`��+����Ø+}N�H4�>H�Z��a&y�h����GE���K��Eʂ]$t�վ��b�&�w�@Ah"�Ō��]�J�q
g��V���o�J�E���W�<Av��8sD�!�w��*��d�Jgy����dL���"�>,�����	�;|:%q�Ƃ+H4�`�C�f�!�����[d���o=�с��D�I�t=apAڸD��p����{�Z��]>�<aa-��u��Y��)V�8;�Xh�KsX�H��D�5d(�y���G@�F!�g̍.k��s#,-X�`xxU�|��`��	� F���+�e���p�.֊YJ�<١%T�&J�ۥ�c���(T�����O��	�@�&�����6VX���'���w��9\���-�8ĩ(��x�ց[���1%vd�q�I��E��w�rd[G�hW����Z[(�B�'��lĄP��* ��/��u�h�BI��A �#I��R˟4���o�'�Fi��#Z@���j\�t_TX��n��Y
W%D�n�PE�+�!l����@a��q��i��d��%j��^�I���P����&�]�Ipu�fb�f���D�l3�v�c���8^�:܂��51�l�SSY�@�C�^�(�V�%\}�PC�I$	��`��b�K�耺t�F !<U�`om�"A�F&S{^a¢���.Y���4�sޅb0�U�Z�b����u�j�#'=D��hB�+�G�4���$LV�a[^�8ⴍ�t#�/�J�z�cF&G���0��J8 �Kt�X%�@����5���d�9,Wfܢ���6 H6��t���c��y��̒�{�Թ�L7nH��Cv��5Y�$!��I"c�(��F�Q��q�%W�DB㞰����'�-���j?L�j�L�)���0�O*��R�Y�8Ć��k�?T��yC�'�8�"4��mA�XId�<P�zlƩҪDL ��$�B��kE���a�0��~��x���T��sƞ��vg��F�D�b �,D���-̸v�]����(0��A%i�t���;'�i��\Ӳ��Q�����9r�Q���'�~<�
f�XC��b�7\O�	A�%r�����D�thVH� g�iؤ�8��^)d�,�AFĦy��-�K8���q�_�jQr!���U�Sjmke�#�	(����`�f��}�����dȨ�k�t�]�E����ȋ���@a�
�yҬǙZ��BF��Fw.`['*5p�t���.��`͸5P'��v�:M;���k���-�!��
$qiJ��nD�M�!��G�E-D��3�%Ji�A#A+E�3�v�S���<�@L����5�Z����D|�EA�JZ�#%AC�Q���rPEX���=	U͟/S�����AKx�Y�͔.J�x�t���WZ���	�N��	a@v@;��Qfѣ�I�+id�#<i�;.ƈ��F�Sy�O��Q��{�>4��f�!FX�];�'��!q҄٩dH"���Y'7�F��qO]&O��Z�Rz�)�矼
��%�����_�q��\��$D��+��<,��9GK�h�
ݛQ�"D�P!���s�v��@�eF�89�� D����&Ǽ_v@��n"tMR)� ?D�\#�FݏB,�u�p�q$}�cd?D���E��:�\-�fC�S���ڷI1D�xB�ٰJ�=�[��40��L�!�$�PMz�Q�Lϔg�MjA����!�dJ�Oc�)(e�ǝ	�����x�!�dӪ}G
8�D�=*Y>ݐ���*De!򄏛[ǆ�p����x@���&�#?a!�$2�	����7DT��(�84U!򄜫YP�@! 6�������:G!�ĝ3��Q�m��<����-�I!�$<vpƱ�5J�7)R}�흽P�!�YGB�뵁9?�@�\%�!�H�Bx�A��� f���oB��!�^X�u
�@�N�>՛�?V�!�� H�8#�Ϩ.�������H��"O<�YS���@6`�2��<���"OHU�A��_`��,*	�}S!"O��#L*RL����!��n���[u"O�YA.��U���ˁ,전�"Ovyc��ppSS�I49��"O�x�/�t:�h��%/�Y��"O�AbU��eD��
Ts��,e"O�)�V��/)�(b�j�3��J'"O�aCP�2�2H1		��!S"O��0�ǻ�P(r�h3�a�R"O�3 (D�/,
9�ѧ�M��@JB"Ore���L�D0 -8�������"O0DR�����|�*�G��w����"O�����$��xYW&A�T����"O&)�e��x���%�����"O���ូ�Q�O��g�d�q"O�<�P.�DX��J!a����"O4��B��}*8y-ȈD�����"O��FYp���B�M�)
@}Y�"O�i3��$+,PP�6&�p�\}��"O�u�b�ށBl��)��J�
��!�"Oz(c�_�}P�Z�gU�_StJ�"OĘ8@��T$��D��@���*W"O>�s�cI�1R��PD�rQ�X�"O��P*8&�,��Gʞ		@�qA4"O����ZTX��2G*���"O�T8ң��/�QF���]�D"O�,)��		~Z�$SV�F��rA��"Oĉ�J��^��c��X�A�p�&"OR��R�!Z���Ыk� �I�"O��"�ŽT�^�:dM�/r�6(ʒ"O�	bu�R��J�.N_UR�h5"O���Vc#����l��s312"O\m#�L�6m|<(ؔs#f r��>D���,�w�	j�&Gu� ��"�:D�X �/���Ƭ8��?
y��ɶ�?D�8� ��#~[1�2>K���(D�䛃�[�^(��y�R�F�����) D�9d*��/,���BM/~HD��s�;D� �a�Z�H��5���)L�f�2�9D�xa`��b��[@\5B|<i��:D��ۖ�nz�8	d�� i.H؋b?D��I�eĜi� [��W!FdLB�N/D��b�ؽL�V��'l�lE*D����.F��Za!�d��F�z��&D�hI� I�6�J�k�*L�
�����$D�x�����T���3rf̂,D��3EߏN����K�B���� D�$�A��2-��zW���8��<D�xs1 鶴�5&ݝD�
����6D�4ĂT�-�-�]��0��8B�	�z��L�k:@�J e۶)FB�I���p�W�eB� x�W�$:B�s��$q&���8�p@��9SB�	�H�vE�C �Q`�����Q&C�I�� I�bذ�d�b`f��C�	1ne�zs�é�����`�=�B�I�q�D�1l�96eHAk��A�O܀C䉩��L3S͜L�N5�C��m�~C��f��LD��~���&�6QMjC�zZT
�3M%���o��bgvC䉟s��3�-^3k�U�@�	/~W�C�/?L�H�c:&�X�с�8�<C�)� ���T´C�uC�m̊��l�C"Op��3�;v�;Cl�{��љ�"O��Bu�ҏ_o� �,�p���S�"O�]��MތH/tS�!n�x"O�����,
�Y;7l�a/�ę1"O��hW��(F��Cu���[!"O\���C.v�I�'*<���"O��#�P����"�$6.�2�"OI'$D�z�x�x5!D�h����"O8k�@<DZ�$����<k�"Oz�J��;|C��r��{G�!"O~)	��F9k��|���SJՋ�"O<)��G���6a����aZJ	Y�"O��B2�;1�A�a��"���
�"O��{`@�)�\��/iwԜ��"OVؚ�+�b# %P� ���2"O :D�4K�tض���9kBi��"O��jo�������4m\2�ڇ"O,ܰ`Ʌ��89�����9ؔ�"O!���?^�ҁr�(�Z��<3"O`@�C��6}�l��B"5���@"OF���2 ���K"�A�!���j�"O��ѱ*�+g(8��oB��� �P"O�}��͈���bcy�"O�0ʷ�3�:�b,	#(_\�HA"O@-y!O	a�)4="D�[�"O4X���}�RHt��'�]ʢ"O������Lɘ��ۋ�I��"O��Y�A�|�*�8D�� #��Mb�"O�\:U��+��m��'�(�� 4"O�]����`�ҥt�ɉ�X��4"O^�Kd`�,��m!0e�F�V���"O��"񥆉|��,P��FPt�xA"O��' �:�Zm��E%29���"O��A!IQ�����4]-r90"O��V��'�\����w0�{"OVɋb�-���c*�j�$*�"Oh9�Ř>*�����
�z�����"O�ZÐS����rE~�\��"OL�y��Q
��ue ]�`�D"O��4͵EO��aD
 0��k�"O&�$R1=t.��֗S5��� "O$Y�a��6xA���1<�
�"O�E9���$(�9�nO$_>.<h�"O��8g���M����a*ļGJ���"O�E���Lrb�8��U;D� Y��"O�x6�ҜX��a㗢��� �2O2���ٵy&$��1���$�1 ��ɫ*ϒ����,@�X�$�V�f0B�I�.�BMjs�_&?�����('3ZB�o�n�x��=*}�����L�h�C�	��� o\��Z-)��Ȗ����(?q��U�~}�5��M��`�<1ԌˊX��-q��UQ�H�1U�
w�<�a�¢��@` "�k���S&)�l�<�*j.g�=�.Ԫ��_e�<ɶ疼KpxH2'UM�ܐ��J\�<�rُNHcƝ=S$pZ�bRX�<�g,֢?%v���G WE�	��nJj�<���7h�� ��DP��	d��b�<rDث��E�2�r�,^j���E{�G(�����"	�2��x����u��<q�����'v���yU�C�2LP<����&WQ��9�V�4I��ا(��$A�أx�}z��Z��76O�9�'
1��?y�>0nԐK: ���E��E�f^��D	�����?� ���Ԉ;?.�Ivcէm���Z���H�'
v��i�'`��p�A�&��Ua�.��Oڹ��i>��\�`y��S�/ت�����!pz��%�P{7��o�S�.PX�g�ݺ>��S���'�%�'���a���ӟcԘ����! �x|S`�ٿZ�>����(O?1�WDϺd�	�	��ł�"ac�<��?3mZ��kMe�2]
4*^�<Ys�  ���'eV
K��,jEq�<�%[�M̆���d��#u�� ��v�<Q�O q���A(��(�6��G�u�<��d��*��=�t�zA�^p�<U�K�N�0��q�5JӁ�v�<���%(�p�ڇ�w�p�³#�r�<A�čA�Mh/	s$��+��s�<�0�\�P�2��@�߂��!BIW�<�� Й-�0�c��,+5�CQ�<�AI b��e�,j�x��&h�<�r�S��Hf
�*�T�#ĬNb�<�p�O��t���n�"t�ƽ����C�<!4�TPj�!]:�����=T��J�M׊GP�[��(1`��,D�$��h�4���CF�0_?��;�+D����n�?U��P�a��t)�	��(D�v�i�ê���j,�+^Rܘ��'c�0�����8�ʹ匊+j��x��'�\	/Cd'���Tˉ8_(rt��'[D��@�1~t��3����2��'��Ĳ7�ù^�003��%Py�i��'z`a�� ����oV�xXҁ"O�Q��R��m2���e{�"O~���
Ւg|��f�OV�8m��"O��{�jP%H���S�|x�0`b"O��"��t[r:�o#O�\"OT��c�޼G�D����G��};"O<� "Q�Ԁb�G�K��9��"OF,KՇU>�\tq��2\{�"O�Dį��@�y�i�6)�NܢT"O�3�Z�i�D�V��D�aW"Oz��S�L� �q�����p<�"O*Ⱥg�?}�x�Zu%VT�\y�"Ox�Z �I3"\���� ,:̪w"O�$U*.�:�c�@�#m���@Ot�<���4\ܦ�S��R �e �iF�<�0�<QLxPc��X���t�C�<i���q4�rD�O�S$BY��|�<���W|�qhEF�	(�\��NJp�<��-�8vA\�����f3�4��YV�<IuaN��{&b�*�n!s��\h�<���:H
fLЙ�4���Ίm�<��@'NO�E�D
H<�!�:�	���S?�b��v�C�!�d�;�Ԑ˄HG�a�Tat(��=�!�d�)U:,hF���p����>�!���f�p}�$+̀{�d�<D�!��;�p��C�� n��i�cܓn!�1y�J�" ��J�����4x!���+�ΐˑiBS����T�'
!�B�=^�yжK��+�>i	��I�X!���(}���#T�2]*6�1a͌!�σ.2 ��ߒy���cj<'!���x5f�s�)^�+׊ZD�C�{�!�$�|O
͡P#�M�E���	>�!���
�3qO��e���1%�ՐF�!�� �,��l�0���!"�M�!�� �4�se˥H�N�s�)��aQ*��"O�ɘg�ωS��E�O�{1Δ�@"O<4BfIE!g��0���DЀ#�"ObT8��Mӄ�x��>�@��"O~��@��Jy����(��+�"O�ܱP�GC�0��0[ɪ1�"O.��"i�&E��ð�>�.�k�"O@з��&/6��j��LĲ�"OX�C�jB
8��i�>��9;@"O�ҥ�%HcV�۰g��i�DQ "O��`Q��6Yd��(��[�B�Q�"O�lySǅ\��j����\���p7"O&��`�M:����83��ɉr"O¬�0�)[�X��W �F"F1��"O̙��A�"_ܲ��ɪ��/E�yrN)
Ll�����	�~�� ��yG�L<b��d�BVI�`������y�
ڀe�$Qum+c�<ēE%Ԍ�y�X"�YG�C-^Ȇ�B%O*�y«��l���b%l�;f���8 +@�ybM�2<�LAbq�-
^�,��
�y�i�d���r�9|�´3G`�?�yr�7|���8�h�KB�K:�4�ȓ_nq�1�ѷ	N$萦�+O���ȓh0�"�����['Z�9[�̈́�~s��b��!�r,a$EB�2�:Ʉ�,,x2V
����i����%�0نȓ �%8�mX*���V�R�5����!!g	7~u�����ޒ
��-��{��T�&̂��ʔ�We�)-�l���$�.y�p�֨Czm�f)�r�L��t�RI !��+;�4�F��ni�݆�7V�m�"��Q�F��e�%���|g�� 瞹+�A�SI��j �i�ȓ?�*	A%r�lx�Ğ�_v�����s�K�����E���i�`���-��1 !��R��72)h͇ȓP�Ј��ŕpf�u�i�	hE���(yy�B��WQ�|�'���8�ȓj�"�Y��XZ�P�(�*n깄�~�*����	�y���TBD<XSd�ȓ*q^��m��h!<0�&��k���ȓ���1���{��)��ί>M(X�ȓf��" Z�h�b�[�wX���G����׋E�7���$Ҽ~�怇ȓx\t�h`-��7P$�s6"\"h��@�.��b��	=�|�U&�5��}�ȓ7b� �I��T}��	WKP�r�J�����QCːx8�6�3A��9��b�� ϞY�at���捅ȓyŎX�s�R�q�X�x��A�5����^�bd�d�@ ��bBi��<�F���elv��S,�gꌨ*��� �Ą�a7�$
���T�,l�րB�4���qr|˂̀[w��!����y�ȓ	>ژ:�I�es���.�(Y���ȓ_nD���M�8�%�P�ը�2�����cGGD�J�, �Rl�ka*M�ȓNX�z��߁	_$��jӔR�\���0���g�TE�4��c%��sC��ȓ_=4�RDwfe��KW+E���ȓVs�T[��?/����R/T��0��G�r�J�
aĐe��@�7rp��;��Y!	�01�A���S4de��S�? ���O�>+�TMc��	3LY"O~��#cP�Qy�tP�h�
N4Y2�"OJY���N� ��8�i@�dhm�"O�e#�AYN	��&ޮh슑�#"O0�a�k4m�~�c(ҳ
s�}��"O,2��D1,a3L�:;�Q� "O�u�L�� D��e�"Qƭ��"Oޭ[��/�>�D��RW
̊A"OX| f��&q�8r�M|<\�P�"Ol%�r�-%�uʢ�!4-"�z"O��pʍ1m��M�D�A � C"Oބ�IJ�,a��Cm޲|z��"O>�+�(Ē_d���'LJFRF49g"O�8�FJ�{A���*�<1�=�u*O<e�#���KO�M���f���
�'=�Q��#�o���D�r�ؕK�'*|H���M�5vјU!�>�&P��'��%� �!z$t�����G��k�'��G��%�����a��P_�eq�'�����	Ю6u�� ���I�H�0�'���Bl�=���1� ҕx^��z�'njQ�#�!=�TE�F(H�;�xd�	�'�0�ڲ R�,\�+#��?3���A�'��[�l�;ޔt钣%1�XZ�'}d=q�OT(+l.������(Bd���'H60���̅
�;�!V7%:&���'�jh�C���&<0Hpd��(��k�'&F�;�Ζ�5������$���#�'8
0��j�c�m��5p����'�,	#���d
d}8��ye�a��'�ӄA �"G>���mϚ{��IB�' �����C��V8��d	@�G[@�<�&�t����7P��A��x�<�b������(�i��8��ae/F~�<a�fG�`Ɇʧ��
7�N��ZA�<ԅ:S�6}��A�npj���g�s�<A�o1p�u�0
8�l$au�Pl�<��N1Rm켁`!�%V�p��	B�<Yq�D�06U�a)N�q�v�#*ST�<�E
�
A�]hP�L+"pP���P�<��ŋW���	��I�x���+�g�q�<7b�'Z���he H��b��Øm�<9ԅ��K�\T�F�ucd�`��!�yI.~�8�I�G_
���
��y"�,7Cz���^?B� tH�hܒ�y��7C�\����F�"ȑ�V��y�%SA.���J2Bi� � �D��y��b�)��CR�:����ǆ2�y��D+v�^���AL;�ptYrb��y���	�@ب��S�d��ac�B�y"	��j�Bd�T�^�`J�J񫑈�yRf�.j�1F�G�j2 ��֪�y"Ɏ�=�e���K%��M�u���y�fD=���S�H*O˒���I��y��$����hKS��� �0�y���[����$Ets�ّ����yR/�=��Ҥ�O.W2�4�_��yRf�D�n}��K�op �	��y�j�)5�n��FJa8��K�AR��y�Ȁ/I<�0eŔ�{�`��P�y����f1� ��M�k�hI��ˋ�y�oA'!>������dq��T�
��yR��zGJ�B��n��1����yb�?%�R �7.������y
� ���ЂE�'�X�+�.;��2"O0z'�T�[��U�K���6�"�"O�dxV��	�^A��*ɡe��I�"O�A�VgV�m��u��	�$DB$� "O�=��E�#���
--�\ �T"O���biQ4j��-�t� V�z�1�"Oaa�bU*�RP;6�� ��٦"O��X��ǆe=@
�k�=� P��"O�I��6l� A�0�
, �JQ�"O
a�� �Z����g�'g� AI�"OĀ�f:M�T-3�
�[�\�"O�����Ǫ?��^�D���4"O��x�
   ��     [  �  �  �*  �6  �B  \N  	Z  �e  0q  �|  ��  ~�  ��  *�  ��  ��  U�  ��  ��   �  b�  ��  �  m�  ��  Z�  ��  ��  � - p M #  �& �4 �B XJ MX �e �n u \{ �� =�  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����O��=���Y�+�F���eIq���JK\�<1!( )�%p@�ř'#�ܙ�TW�'w|��I�E�J�����{�)"�/�F��B�IX��-Iӯ�7�ة5�Jba�u�	�'XJXw�
P��-��I[� �l��
��� ��{�*\">d 0� o9f�:�"O8����e����!(�"R �R"O
=�kZ�t�:f�C(kA@B2"O���1aT�l��yj'&�8l��u��"O�"3�	K�,@A�˽\u���%�'�剁IQ,h�A� 
��T@* �L���'!`5MV�+�z�i�ݕ.G�P"��HO���Q��cD������z-�"O�܂���u�0"
]�8�Z���	��0<��	XX���0��r;�}k�c�F�<	E/�����b��B���t��E�<��NʭZ� �被�������j�<�R�)����ɀr����F�e�<IcY�n��,��%�T$IUF�M�<QCK�@�������Ip��EB�<�e'��%�!A�*Q�)�THX�@�<Y�!]2yΈ��� �I/�P����p�<٤H�<��y��фk���Bn�<�1�D|L��a��=�m0�yB�E�`+X����I��A��y���':�kQ��h����y�+�F,|��Z�0�i���Z��yRE�!���h2ԋ+
����y"��;(?�h��c�!T��	i���yB��/4�M(���M��9�����yb��>��| �Gd����X6�y�]<�B%�]�9F���FOR	�y�O�n�Ε{T I� mVt���y���$j�(薫�%+'��#"\�y�
8Q�����'�/��H�r+M��y"nƜ����6�X'"�v���g��y2$ɏz�6�t�V|(�#B��y��$`�]s�Ș�{`<��A"���yB E�P�t�*��5�&$�O:�y-��>Aa�'����rB�y2��5�P� e%�a��ID��y"�B?`Ȏ�*�C�d��A�@��yr��u�6JCf_�Vb��p��5�y�h\3A�bP�T'2�,�$#݈�y"Z =�<��홢
<�t�s/U��y2���0Բ��e���8��M� �y� �mz�ʒY�3�Ɛ�y"��n�Hո�$�9;
˦�,�y2H�4 �	C��$I���v���y�G55�4�u&R�&� �y2Q��^Y�Ga�S�&�2��E��yB��2j9�a�V�OPJ���@ԋ�y�B&o Q��#�K���x,��y�І//�P[��ϬH�Tt*���y
�pBMIA,)>���y�EY��y"�Ԍo6\����m��}H�F�3�y�ѥ}LHS�O�uj�-h���,�y�oGn]��{磜s\�ʣ�ţ�y"b�d��-�F�m��H�Ē��y�8����o�&RzZU�1�A��y���:3�R�`�c��IY�Ԋ��׶�y

�}��9"w#<L;\���5�yb �o�rq�' K5�Hs#�(�y2L� ���� 1�9��뒋�y���y��Q��Ϗ*��� ��yR��v�iq/_�B4,�n0�y"��d����f!�o�!�y�9X�A�Dd��m�	�΂�y���C�h��m!�0��p�1�y
� Dd)��5%�Z&@ń�$�jW"O�D8ԌE�Vv� �n��nϊ�1�"O��H�C�Zt�-ȵ���W"OX���W\��B�ʙ&.Д�Je"OԼd�2!#�1�e�y�1�W"$!�$��2r�e("CY��9$
�!�^ 0!���6-�@x|0�S�ʣwT!����@�f�8n<+ ��f0J!�|a ��H�X��i�GFb�qC"O�EVȕ�}O�)ȗ�N?;气)3"O
�P�W'/a��� oB�e��ۇ"O�l�g��5o���5�Z�hd�X�"OVPcE��-[L"f�ԋ�N��q"O�<� L�2/�>mzD��*$<z�B�"Ot���&��Q?Ψ� -Z� D��"O,9�ā "�J��!_�(� "O�p�b�3(1~�C�GV�P����"O�tx���a����b�/)\� �"O�m�Q ڂ,� �
�l�p%���%"O �Zp�_�i�B�g
\�@"O��`�&ȴq� )ISIW�\|h�v"O���eCʙE�U�eK�]#�]ٶ"O���F��J��U$�{�a��"O�`�M� .�=$�أ�i#"Ol!����	.��`�#5�<��"O�i��
.�p\���ۛ{���2"O$�Q�>�܌[�J� y�L٥"O�5�5����*�Hüo�h+s"O��q��j��\[B�ԣV'\q�"O ��7-C�4�2r%��N�]�#"O��*�
�,p��w�E'J�����"O�=��j��o����	(&�NPh�"O���n˱v�&mp���)�j�%"O�5��JG 6��3E�,��"O@d�ˡW�`�p�)l�J9��"O���fN�Oߘ��
�) |KE"O��T/�&j���	�W�	U"OL�ˆ����	>)���"ODEC�P3c����C�	~;��
7"O���`B�M&6p"��eׂ)k�"Ota"ĬT)�!�@�U�V��� �"O�P��BQ��2��D9pf�	�"O�|�G.�7t�s���e�] �"O����J�'ajH��J�lfd8�"OU�V�M��Hq��K!Xd���g"O�0K2�̳��1��U_�i�"O�Y��+^�.lZD�\	E`���"O�\��J���ԏN�JVh�"O���D��U0m���YBtl�"Of��A�r~be�E�M�L<�x�&*O���� 20����!̯li����'�.�����4`���:BM\!a��B�'��t���;p�T���
L�.(y�'�� q���k�h��H��A� ���'wbQ0 ��`H�E3�	��f�]�'�L%��,Yb�(��J1l��
�'<rq�����"�����3Ggd`��'����i�&B��5h��ӜA�T	K�'K�m��	�r�.�{'�¾<��B�'N]:ǡv��)' ]�H�X�t�<�i�:0�8L#���ir�����Q�<�㭄2	�01eK�Bl�5�2d�<��g�&H�@�Ň�#D^��F_�<��aW�Pd���*=��h��F�<� �Ѱ�NC;�4�xi�"�� �"OR����PJf�+P'}j�Ѻ�"Oz��D�'&���sAg_�qP(�"O�ݣ��	0*�X�DlS�%"O8$���¨c�h�GC1w���P�'�r�'["�'2��'b�'}��'�ʀ1#�ޏ�vة$Ş�8}|\B�'�r�'�r�'��'�B�'w��'�^��%ȠI�	���"Vk�H1W�'b��'d��'"r�'���'a��'l���*ĸ]�V���
���'���'���'���'�2�'���'������Д
c$���́mҒ�r�'���'�r�' R�'��'���'�-34m���$q�h�r��{��'�2�'���'���'���'���'���"�CD6;>&���/_�)�Nț4�'9�'$��'P��'���'[2�' 谊��Vn�3�k�s1����'��'���'92�'���'�B�'�W� ,����e..�M�`�'�b�'C2�'�b�'=r�'��'��h��BM�{͑8�(\P��'9��'�B�'��'w��'��'ǖЂDE�;���#�!~���'w��' B�'<"�'���'+�'y�D��N�Nb�0�ǃJ�d}�A���'��''��'��'t��'w�' �H3��,q���1ܪ�I%�'�"�'T��'���'��i�8�d�O�$C�MB��(�RmO�%"4Jiry��'�)�3?97�iy&�X�c�(UB���g6������D�����?��<	��Jm��s�hНD�yxN�:!<pH����?�4�Z��M��O��8�I?1�S$�f[�,��뀱��94����'{�>kڀ_����� �d��\j�S;�M�!
q���O��7=��5x!�@�y r,��I�D�!�'�O���e��է�O��(��io�D�&62~�
����1@B��x[�df�����$�=ͧ�?!"�ަ"�!��-����s4��<�(OP�Od�l��bRFc��!uC�:�P-�v�=a����J]�o�	�,���<��OPLҁ�\%�������8���H�I(g8��8$�'�S�g92�Gʟ�A&�	�`ɜp�3�E�Ҡ��_y�U���)��<	�#���V<9D+�
BrVmAek
�<1��i�R)R�O@�l�I��|JǯM" ǖyC�! ��XeaU���<��?q�lH��ݴ��Dd>٩�'6���!�K�����9᪋#�ic�i(��|�/O���L8�mu^aX#���a0���4$N���<q��D�.��[�������.�J�ꓷ?��yR����'��F1#���
cIQ ���`��G��x�������	�+�8*G��OvŹL��Y�l�pi��u�N�	�E�?K-�l;��Ɵ|�'���F�	��M��I�<��˃t�#���~�ę0���<AF�i%�O�9Ox�d�O��/+4�%IV��=7yAI���
("�p�j�I�(��ɑ_W��ܟ2���*���1r��y���) �0��Oi]��̓�?	*O��S�O��=��l�d��<��f^��K�yb�|��|������ڴ��"<LIg"�*O&��%�6�~Q��'$�I����Işh�VΖ���?A��Mz��1�v�R$���@�A�d��O��i��4����?� I!tE�Eb�J�;��x�6-C�<IO>ᇼi)�� �y2]>�� ��M��9�G�f��Ԁ��8?y�^�������Γ��'�?!�D�,���B��	s�|y�Ɓ��?	�(��X�R��'5B�ğ��q�|RD�C
"�ٲ�B�%Fq�L${2�'%��'���tS��	�4c蜵caLV�!j����HˁR�҄q��
;�?�l��f�$_b}�c�d`��@��$�z���~�*u9%f��M�Ʌ1��n�<��}�=
t�nn���'�,� 
�B��@锯���'%�I埀�I��h��ޟ���y�4"�Rr�dsb� e0��j�2S�7MP%aaJ�D�OB�$�i�OMlz�͒Ģ?Z�x��0��=���s%���M��i��D�>�|"�iϜ�M��'�|�f.�U^��`��4&8��'��se���<��c��|2S������� �8x7T�j#Α��^@��_ş������Jy�h}Ӽy���OP���Oҍ+W�O �T|c&�<E���6I=�ɷ��ğᦩ��4�yb[�H�R�����3�Y�h��ī��x���03e���־ �F�:?y�'#���h]wצ��ڨ $���`��T��D��a����O �D�O��Ľ|��D�j��'�|!�@/*D��	jn����''�6MQ�NBV���Oj�m�H�Ӽ��B�T����\�ȭ�L�#S��DΦ�k�4�yB�9�MÞ'��n�b�ٺe*D+d��=��ł�cZr5����j��)��|�_��ǟ������	�L�R�E+g\�]ya Mt<ʱ��UKy��f�bm8E��OP���O���R��dbx /V�8��2+ط;�zY��>�P�i3�7mr��&>��������G���c�K07��|�1�YJ��{�;?�F�����0_w�P�O0�wb���2K{&YB�H�z[fQH��?A���?Y��|�.O��l�T(*���� r�B�f��zQ�Z���=�I(�M�����@n�ʟ�l�ҟp `�>K�LC�.�9U5�H�P
�*�n��<ɶ*Gq"�7 £>��S�?��;u��8� XyIw��l-Z��4욧h^x)
�<O
�$�O���O$�$�O&�?�z6��"|�̠ن�R/-��t�1i�4�	؟P
ڴb���'�?I��i��'v�͡F��/���j�]�%J��47O^�O�V�|Ӗ�DV�$[�7���+ׄӞl��j�Ҹ��`3���9񺈚 �R�wQ�k�,K�%��4����Or���,R!,�(� �eɢ��E�KO~���Ojʓ9�F��"�'Y�U>mISD4xޜZ���(�%SE�:?1�Y��ݴ]a�F=O0����јK\��#��{�LQJ��w�x��EYV��������Ӽ1�,e�;t��'eDa���Ɲ���Fb&]l̓�'Mb�'"��O`�ɒ�Ms���v�*��ղ+�"q�3�,'j�mp��?��it�O���'��6MTc��c��ƴd�r�@�����plZԟĺ��������?	�ϋҲ��l~�
ê*�(JaM��$x���ې�y�]�4�	ퟜ�I��h����OBX�b���61#�]H�T�� 8S��f� � 2&�OL��O���N�$���1D��=i��˵Ŋ�Y�i�w�T�	ܴw�&=O��|��'�?Ǣ��Mӝ'AJ(��
�q��1�%*�s�'¨p��I!����|�T��Sߟ�b����HC�B�+�}����S����������iy@q��q�O@���OrsPs����*0��u;��'�I���D�OB7�a�8�'������ ���`��Q�.}��'��(T���������X��ku�:�#����5H�32�eZ���6
j��!���?1��?����h�����NQ�8�+�?`�fԂ�B����\Ǧ%j�e[̟��1�M3��w��m)r/�N0d���ִ%Mxtȝ'"7��Φ��IlʖEoZ�<����<�ӣA�X�����J6|��iIE�մa"�]R�iԣ����4���$�O��D�O��� @����w.��Q�00���3��ʓse��`HT�'U��'��OW�!�w�h� "C.Zb��k�@�M8r�	�&$j���N�O��t���h
Mr�A�R1ʼ�eHJ�I�|\X�Or�yӋ��?��"-���<�E� ?�
0�7*�J�nUj$�%�?Q���?����?ͧ���禕Jƣ���ؤɜo{0�r+ġk�,���ϟxy޴��'�˓�?�ܴ�?%'� 3����DD]�$�`AhǫN��Sܴ����*u���'�O���X1C(0v�׮N�ڝj�oL�������d����L�I埔��z��LUX� `�Фm�p���Ȑ�{�i����?��I��v����'��7m3�$��-�*����p����t�ۄh��In}��l��Dlz>M�s��Ӧ�'l�D�@7(�rL	��کe�԰�ִw�h�	�p��'��i>�������T�6�U�>6֞�r�l:}ަ5�Iݟ4�'��7�ڇe��ʓ�?	�'���j�1wj�D6��9��F��k~2n�>��ipT7M]Z�i>����ZN1;4+���a��U��Z ���S{4�(�]Ay��O�D��	8tE�'�ld�Ĥ�?�9�6)E�%��G�'{��'�����O�剶�M�t��f��i�B��.ੂ�����p$x���?9�iy�OL��'ۛV��GL��	 %ɲX��E@%͙Ah�7��Ԧ�F�����Γ�?"�ʀ9L������J��
	�
�%-��="�.�wg�İ<���?A���?��?I*�0i"��(F��pK�Ƣl��5��V���-�Zyr�'���Y>�����Mϻ'�L\1���% �ı����Vd{�i�7��b�i>a�S�?%�q�%�L��S@�n��q�k�V(I��`��f�OZ�aO>�(O����ODa�잵-w XP��C"VN����O��d�Op��<�׼i�\�أ�'���'���¤͜3��h³�Ȱ1�8�e�'M�'>��vn�V�jӞ%��B�ߚ2?x���+(�4�ws�P���aP�P�Y腙�Oy��Otl�ݴ;����� V��bQcO:2d~]a���Zi*��O����O���=ڧ�?��D�4|���2F�:(BP� �����?�&�i��yX'�'�#kӬ��5�4���#gش?�������Cʖ��b3O\o��Mct�i;dpBc�ib���Or]z��"#��A�� � .��$��؆�0�D�<9���?����?I��?9qh����B�[�[���ó����Đ��=��*�ޟ���͟���m�4�'ip�r7-� �4:5L��I�(`y��>4�ic�7��E�i>��S�?��/߰?p��eď5�T*]04c�Z�?Pі'�J�ӦLڟ@E�|�V��i� >L�Y�G��
Hδ"rf�ԟL�	˟0�	���Py"�a��!��O~� B&B�q�05���˨b�#1��Oxl�p%�t��O8�nZ0�Mӱ�i��P�D��@x�E�a/ʆKZl�v�� k��9O��䍭k�(	��'�rʓ���;]:8�s� :S���ċ:F��q͓�?!���?����?�����O�dc�+�*v�L��Q�o�&���'���'�N7-V0b]��O.�l�n�ɨ=���	�L��&V�J�E�{�����y��l���)G������?Y�I�O:l+Ă^�<͒���u������O��M>9(O�i�O����O�� N؂7Dd���<�dr��O&���<�йig�]�'���'1�S:���x�ɏ�-����ȍ(��%K���l�<AJ|���po�����}Tt�D-M�b��U��&P�}��X�@@s~��O� ���f��'���`/ŭD1��5�&����'���' ����O'�I<�M�5h�+2�!�BD��ܔyV�(_P ����?qоi��|�>�A�iȰ�1n�;^@���W�)�x�At
lӰ�dB�|��7mh�`�I���9%�OŦ�S�? �u�j�"欐Pҫ��M/
�IT>O���?����?����?A�����Cܙ���U(�I��=D�l�	zﺱ���H�	�?��O���|����u�F܁b�
'sjX�H\3��mڸ�MK�'�i>u���h�!,Z���̓P����� �;����%FRO�e�ӲU*�_x���g�IQy�O�R�o�(����T[���"H
��'���'�剻�M;����?���?�EN�����@G*j6D !����?!I>)�P����4>�6=O�NȞy�wƗ�:�%B$���A�cgj� "h	"5�zq��@}ZwH�ђv��@�y�D�/�����8���	�Kܟp�Iӟ@�Iӟ�E��w�☹��\>V��ܺψt���'��7�;pv����O��mZx�Ӽs�eF2W�xu���Z/$��[���?i��MK��E!���۴�~2	[�!�����h�$S��	� v�h��O64X�]c��[���mj�i>�����d��ן��Ɂ`���)ގ#�b�(&E�?%�ٔ'�6-�R)"���O��$'���O� �`�7T�x)��N�E���H�LT}�Op�n$o�Q�i>u��ן(��҃zk� �&C�+��)�7S�C!v���,?&�&�Z�d������\Q.-��b�,yAvI��[�N��O����OL�4�@˓EE��b 8R�����a���iQgL�I���˃e��O��o����r�OT�m6�Ms�3Y����^D����SP���$�M#�'y"b�_Q���:�����۝ep�ٕƐt��IٗE�cJ���ON�$�O�D�O\��7���P8����>a� }���A�$)r���۟���<�M�#LN��Mz��Ohx�d�հ/\������ k|��gf��'?6�ZȦ��ɚU-p�n�<��^�SAǵr;��c�I�8~�  �
D6"z�D;����4�����O���?2��A��R��c��E�e,���O�� .�ƩE 42�'ubR>�!`�/�ܠ��	�ut�(��$?�@\��M��id��8��(ZG��A�
�T��i�tb��:54���h>:�tI�I:?ͧd`�d����Bp���7�X0kb^m2	��10���?���?��S�'��D�ڦ�C���I��B��7D���&电H/��I�����4��'����F�?[:��e!��fθ �B�NW�7���QB7a�Q��?Y�I��,��1��D�-v�`����<�����v�D�<���?���?A���?	(��\u.������(��4�U��+�E�ś����	���%?��I��Mϻ*Fx�(�9����)�4F�@Q��i7�$�4�Z�I�O~����~ӈ扥txH��F R$W��*X�5�N�ɻk&�B��'V�1'�����$�'�Ԍ�AG!̾e�g%��k.� ��'@�'bU���4T�(O@�$��I��t��kG�@C�A-}:�H�%�dCV},k�6el��<ѪOԨhfl�]��!;v-�	\�E�W8O$�����1��^�h����?1C��'�*���2&���	�hΰ5�����1+}�IԟX�	ޟL�I|��y��a�|�9厃e`�lɈGb�tӼ4+�l�O��dE릉�?�;M�>�p�O3R#�=���QL���7N���d�|��95\�7Me��� !�DZ��O�t �0������D�Ӻkє�� LR��{y�O��'�2�'�C꼁e��r��0�e�+4U�	��M��,����O�����dA1'��%R�'ͼ ���a
 JTT�'	�7��Φ��ħ����r*�5K�%C�/��L��e]��-2�e��KYbD�'
8�P-K��d��|B]������uy���`�L�"��$P#��������̟��Cy��k�����OB�Qb��(��9g]�<�D}y��O�il�B�p
�ɢ�M��i&2�GkW��H�Eҝ8�Pp���V�ܹɅ�i��d�Oղ�*^��z����ӱ�5v�W�+�b�i�)�0-_����O��y��'���'�r�'���	�*B(�	�]9��YQ�mG,������?��Pƛf���iW⦑&���� �"iTذ KG[L�
t.��<9*O��p��UzK
7-)?5/,���B#�D \5Ҽzab̩b�b3���O�M>!)O���O
���O���a���T�L��C�A�l�����O����<�`�ie����'1��'3哋'm��i�W[B��P�0�T�>�I�Msd�i}ɧ�� �����U �H�<չg��8���r/��1V�9����;4o)�g�	C'�\Y$l�3*�&�Q�������Iٟ���ڟ��)��Vy��s���c��2�OȊ;�*t���A=/F�lXD�'��`�6�Ī�OL9mZ�셺���2(�4�!� ����ش�?���@��M�'���^�V���S�����,^���D�G8HW^�Yw�G��Ĭ<q���?���?q��?�/��*勛|��d��[�,P�ԌN�q�JZٟ���Ɵl%?����Mϻ�dP���3��1 Hr�^�Aɠ"}��`$���?����m��mZ�<�6	H�D�Hx��H�=��xp����<	Ĉ�9�����������O��D�0����@��#w>\Z�a'R�<�D�O`���O��vr���;$b�'bA�&5����X�.�di����:�?YS_�dy�4Wě�*6񤄣)�D�!"�*G���"/�6�~"�'B��)r��f����CV�(�ә	3�Gɟ���	� Y�����<?e�9���ǟ��Iԟ�	ߟHD��w�m@ֆ�R�D�@+яAva�B�'GN6mƮ"l���OR(o�P�ӼK��PB�,����0�dՉv�W�<!b�i�&6�Oᦕ#���̓�?aSH�y�d�	SH�? DP�����vb�`��TtҥI,�ħ<���?���?���?��L�c��)�G˃re��9�f���$����vL�H����'?M���t��A�D7\��[�
�4�t�ȯOx�n���Må�x�O��d�O��؃@Ə�^3=J֭_,-ZZ��aO
R���j%W�Hi!��W'⪕L�Iuyr��=�x��n�&#D^��7f�"6�b�'���'P�O��M��[��?	$�Xu��ٓ5%B}�<u�E%��?9F�i���|b��>�@�iV�6�P����uOB+rD�$jg�ʞ���c�)�M��l��<!��mb�������A.O�����l-Yѫ^�Z�zQ�S&%� 2O����O����O����O��?q�cc��v�j���M'"�8�y4n��������ڴ}]�	�'�?yF�i��'پ9�@��_�8\��EݲF:�2�=O^�n�&�l�*���/�.6Mh���I�oB.���c׼C6ly�,H3o��D
#
6���w�Icy�O*r�'�b)�``%�ͧo��#��:���'s�ɸ�MW�N�?����?Q.�t����s�z�k5,�}1�E�P��p��O�Ul�&�MK�'��O��d�$3c�<�iJ	9O$T�%�Ԡ[8I9���|��O`�)K��?)!�)��T�̪e��d(Vg*`�`JM<�����OP���O���<Y$�i�m�B��V�~�PrF��๨T&I$��'^@6m5�����Ҧ���Q�sl� �Pd�"�X97�ђ�M#�:�v%p�4�y��'
�](s�B�?�b�O,-�%Z�������/(��t��:O���?���?i���?����i?|)<`����xX���!�́���o�)p,��	��	|�S�����sB���H����U1E���e��'A�iVv�O�d�O|�t���g;��5OTHAU,��Ez�HJ��L� r()s�3O����%�?� �:���<����?!!΃O�ؐaGB�,�, j�@���?����?�������Mf��ޟ|����H�r���Xa�N�,��AE��1��	��M���ie�O�ИV��A�܍�EZzs4�a=OZ�D�J[`��Y�X���T��OXc�eIl�S��?qTx�TI� 8�tY��?����?���h���8�D5�O��v��|����_�(�đ���2���ڟ�I�Mc��w���4���jܖ ;����t��'�6��Ӧ�"޴�����4�y��'���H�+��?��$��ZT��[e��H�����62�'���̟���ޟ��	ןL��9)��A�p�]�S�=��@�T˶Ȗ'+x7�«\���?!H~���e
�q���c�h��LL8�^�Q�Q���4)ś�A5�4���I�6m2`I'#+Ա9�a%"}h]���=CI�u²c�<�u�6z���Ȏ�����P�w�Σ-���#c�#z,b��OB�d�O��4�2ʓ:ߛ�E����P�zĪ�Ö44$����� ��e�~�<�)O��diӞ�$�>i+�eРa��F�(��C���`(0�!l��ϟx�u΀�|���C#?��'�k����"�
�<c��]�lN���O����O����O��$2���/Q������|^��u��5$��'�B�t�(q�c<�h��^Ȧ9%�P�al@
#��kc�"���S ���A���y�����%%�6d���	���޲��x	$�k�"��C�Z�H�G�Iy��'N"�' ��Ҿ@Zp�Kը��� ThDkґ1B��'��&�MS�� �?)���?�-��p��B֫8O�ۅ"�+o��ך�L��O�l��M�Śxʟ|QT��,A2�Ҫ��ԋrG�Q>1�� A�/�h��|��h�O���O>�'$�!c�,��.�FH�;�N��?Y��?	��?�|J-O�em�g.���K0�I�1�����ˣ'�����Mۏ�ŧ>��iI8iz�G�X��d�4^�	��i
��s��$oZ�w|Eo�@~"'�Y��X�ӗ	��	�I�<�T�J>h�6iJ&�3U<��	cy��'���'�2�'�bX>-:`�Y�]Ԣ!"P�Ϟ}��,8�@^)�M�� 4����O����D���ݝD�3D�&�֤ �H�xr����4�!�4���)��ҤK� qӒ�ɤ!}k5@�tӼ���i�?�~�ɲV�b��'�v�&��'�"�'��R���p B���Ǟ�����'�䦽�IyB�uӒ���O����O���\��A`�I(\(s�K�O��OjY�'_�6HѦ!���Ƙyv�ɱ�V~����+�}���O��a�GL�G�j��6��0�:��o@�<! �	�.�V��dNQ�@�����t�	˟��	П�F���'�M�t�9O.�{�/t���'@�7͎q�f���OJxoZR�Ӽ����*S��¶��|)��ˇ
Y�<1W�i��6��O�Ur�Et�v�{)~�Ӷ���z�j��(��"���(�4�d	W����4���$�O>���O����
M�\$qEIt�h@�6ꆫ)Q��$�Ə�6Q4��'"r�O5�ޟ|�҂Ӊ[�t�S�$�#�9Hⅆ/���BҦ� ڴ�y��T�O^�n� {�~а]�H>�-;b�=+�v0�!����ĕ#W&�X���O$˓'J����j{�8G�}8�L��?����?���|�-O=mZ�YZ�0�ɋj
�)�#c
�`n}�d��H�ʵ�ɹ�Mˉb,�>���i&7M�O�8C�KL
:�>@�G� 6Y��c������7q���I�pLRi��OW0��ü�>�@�&�-h!C[�2� �s<O����O����Op���O��?1چLNuF�}$.'��4��h��(��䟰�ڴ:]��'�?�%�in�'F�*B���1���CѮ?(_��1O,��?��|�b�^�M��O>�RC� f
����<��
���F\��F� �?�BN,��<ͧ�?Q��?���AP��@�dǐبwN��?����?���!3�lH�?����?I������dD!AYY�6�厓7��$�vyR�'ٛv��O|��Y�>�b�Q��Ck�d�� �[v������^�p���O�����?�pI-��³���jX�&�V�p��w�v���O����OL���<�A�i���UgK�}� �\0��!�-@�]f��'� 6�&��3������3ԅ�9;'����N� �rY�Piѽ�M#�5��Iߴ�yb�'�윻v.��?���O�]�6���n (٤E��5�����7OH˓�?����?A���?����	W6v�Y�h dY#��8I�Ē�ћE��$��ߟ�����y�
J(A8(�
d�b�C�Oh�6-�¦�Γ��4�*�i�O&)Q��c��6Z�nx˶��y��Ax�Ꙇ[0 牵l[j����'��m$�����d�'~h�֬��H��s��)+�f�?	��?�����q+��Exy"�'1Zei����!���
uhα��$�}y"�'���5O��o=�R�kEN��cU@��"A�ϓ�?��v�6��d�}~��O�q�	"{�"C��z͡�%�%r؈C����&�'jr�'�r�sލ T/
6��86aS^A��r$I�ʟ�k�4vw�hJ���? �i��O󎅩8�$����ʓ+��i��==��D��U3ڴ�?�1�Ӱ�M��'�����'�����R{�`pg!-	�����ޫ$�f�R��|�T��П$�	ǟ|�I˟oQt03��f)����]����6�*�"�'6��4�'  $�AO̡%x�8����<!rȸ�>��i��7�n�$>]�͟ ��"	Eg�	�P�ؖv�jܰs�A�V��R�$8?�ag�%�(��L��䓧�՗G��5���X�A��� ʹ\p����O�d�OP�4�0˓r�.��8����g����4�R(j�(�`W�](,�B�i����OPEnZ��M��:�(X�Y�H�ls�,Hw�Z�h���*�MK�'�lY8F�y����$��ฯ1*$2��g�-]�" ��
B�Ę��?y���?���?����O�~]X"��(�(��!׊|�h���' B�'7D7���S�M�I>�P�]y)B�Ӏ��r�ؐ ����y�R����4 ܛ�O#(Iʦ�i/�	�"�� ��E�R��g�ǟXD��wE_b��.\��Gy�O:�'ZR�-��%��d�
o��*�1G���'�!�M[,��?����?Q-�:U����4�!�R Ң&j�4ƕ��¨O$mZ��McM>ͧ��w�������R��aaPe�u,4i����}�v��'����Q0 G�|b�P�F[��"�ڹi�"@��� ���'V��'����^����4v���B�3/�Z��c��(�0#�c�*�?��U/�6�d�Oy�i���+���U�XH�(Z�r�%"1�iӂ��{�X6�g�@�	L�n����O�Z�8�$�EFȉj���Q i@Y�� ���d�O����O��D�O����|��!	��t���$��H	��	U��HLt�b�'R�O�S��`���KS�Z�<HV����yf�`�Mt���h�F�O��6���w:6ma�4�$*�%�Z��Rl��
���Bt�t��Q�E�,���\o��vy�O��G��wҊ]+�FHQ �@�v��L#B�'5b�'��.�M+4��(�?����?y��>�t��FO�I5��%�� ��'���ٛ�+l�$�O�9 ���U$��V�����}��5O"��W
T��A�l�'%O���?%aC�'}�<�����pO�:V�j��������럔�	Ꟁ��[��yGˈ�F�\Rc�?Wҕ9�+�2�i��.cU��'��6�8�i�Q�E�L4���L[�y�"�q�'e�l��4s��	~Ӑ�1$f��ڟ4��lUq��サ F��sG�#$l�;���=��Y&�̗'���'�r�',2�'�|�H��X�"� p�aT�E
�Ц]��[�4?J8��?������?	� ��v�h����(P���e��5�M�4�i�JO���J�ɒ�L̚�8$�E�<�dUH!e�#���igf�L��ʓi7��+�F�O�{I>9/O$;J�;�B�#wD޺u��T��"�O$���O����O�ɻ<��i%HQ�'�Xx�!(��V�U�@�Z�T�Xa���'��7�*���������!ݴ�yB'�G��!���>$ˮY�,B�t�JiH�4��I25z�)�'�O�7LaB�lk�	�v��0���y2�'���'���'n"��K�Y�@`�f���:��֍C����d�OL���1@�>����M�I>���Pq�ʉ��U$S���G�����4Z�6�e�L��T�6-e�`���~�yh�p�ƴ���$n,0 k���l{�	Vy�O��'tH�i�I:S�E�g����wѻB�2�'I�I��?��D�ɟ<�I�̖O������hs�&lX�-�\a��O�t�'yN7MѦ�$����?�9�aC <G�jJ	���[�-�e2�c�6�����AG�OB	+I>��!�z�K�JâT����f���?���?q���?�|*,O|Lm��Z��D�6�0�*�K�I�E�D�8�H՟\�I��M#�B.�<y�4
�"�)��X&L-`T`FcߙH�����i|��ΰf�v7O(��ɪ^�^���'fg�	�^c��h�*`2��l�w/��	Oy��'���'2�'Rr\>]�'��!}�80!EǞ�e�ES�\>�M;��T�?���?��'��)�O�imz�E��؆9��d��o�$��Rk\��M۵�iXɧ���ON��پXY�6?O� ��9ҮJY�pp��l!�W=O��H�@���?A��6�$�<ͧ�?�`e16�V���S|t1-��?����?������æm�k[�����ȟ�l��n��U�M�g`��#Da��Bd���MS5�iLO�|�D�@�{�
��#	*g$x:F5O��G*.`hD�Ǘ�lDl���@-�O���S��@	�W�H)CϤٌ����?Y��?���h�n�DJ�=4
$A�K�c<������
}���Ԧi�T��ߟ��ɜ�M[���UÃ�M���$��{=ځJ�a�<�ܴ����'�@A�i��	{��R��O��`�F�L�"��׎��֎���][�@y�O���'6�'XB#��p�в(�2=����uCF�d�I)�M���I��?y��?L~r�:'mb���}q�h��)	Ǽ�rS��۴t�F1Oh�����O�|�Al,����sM�-39n�qǃ��p�z�"Q���
#��� y�_yb%�-<�����&j�4��K2Lt��'���'�O���Mc3MY��?a��=�ܱ�f�\�(H�����?)Ѳi4�O��'�7V�)��M�x�B�V��Bl3�M�3��	�%̈ͦ��'s�H��'�?��}ʂ��
�2��	z�S� ѣ!�00``6O����Oj���Op�d�O��?�s��^�W�T��F�Yfi����� �IƟ�Iݴ=U���O4^7-�O��
�N�����e��hS�ߪM�����x� jӢ}oZ�?�����ަ�̓�?��Q(L����,�j9
|Hs�C�Z| `�%��O�i�L>�-O*���O����O[u��D 1���~%ޥ����O��D�<	&�i���3��'d��'��^��0rF���L�w�݀E�
5��8�M#��i�O�i�Ţ'�-8V�J�&���	tgX,n�L��E�;}`˓�2��O��O>�4,��d��l�N��|;����?y��?q���?�|j(O~aoZ��B��F�/��T��#�5f��zt���	.�M����>���i��j'E��Cݨ=�(������qӬ$mڙY�@�l�B~�%��B������I5�,�Ydh `��H3GO@�Z:T��]y2�'��'B��'��_>�W�	.�(�Ekʮb��Y�
�M�F�^��?����?	H~��1��w��M��~7�-���Q �N�ڇE}Ӡnڌ��Ş��yڴ�y�뚰{�
�0�F�; �(�  ͅ��yҮ�2Hޅ����'I�I䟬�����ݨ�-B;5(V�
�$�X��	ٟ��	���'J�6��*����O~��
�l�dRA��<Xt���n�c��⟨��O�tnZ�M{�'�ɲ2U�u��)W����b�5���W�D�A�#V�Aj6M�|R���OpMQ�`G�t�")J��F�S�M��,����?���?Y��h���P�D���"�k_�&�8ݫ�b��_���[������$�ɩ�M���w�R��7�K(M�|qf�Di��p�'#�6-���I�D́m�y~���DJ����0{�<qC6(�-.�DY:#�\A�D�i��|2W�����p��ȟ���ar���@��d��_b�a���Iy�/e�<�sm�OL��O���H�D+Pir! 3!�� @�Tr�̂�rѶ��'�07���E��H��d�b@ì0RY�FFǨ:0ܒ@��2S���"��@�%���e�Fb��Uy2 ԑy�x�*�(���X����/M ��'�r�'��O��I��M�W��&�?5��8;��pge����u�!�?٢�i��O�(�'�87G��IH�ʀO׈:�Պ1��0\���B֦��'@x� ��?m�}�`�ƌ��Eg�$���*��0w;Or���O�D�O���O��?�ѡ���5a���ˉ(T6h{��ޟ���ӟ�X�4}#��ͧ�?Ӿi0�'��*�.����
�J�� ��/�y�P�P�4L2��O$�P�i�I;vH��%D1�p����[�vp-q���;V�_�Ay�O@b�'WBd� �1��	~ךM�`�A3f	2�'P�	��Mv&��?����?	+����f��X
�q� <�ɢF����*Ob�d`�(�IT�'@,�Zb�זn�񨣩�8O
��B��J+e�"�Y@AK~�O�Y�I0t�'�^x( �X5U�� �`�A������O��D�O4���O1���T4���Ao���$a�/yQ�h����G�����'�j���t�OlnZ�mg\t ���%'�]�eL�@b8���4�?a�A7�MS�O$���K�*O?�G� 9$���3d� �j-h�Dc���'���',B�'��'X�4J����`�@9(۷n��Z���{�4h�����?�����'�?�Q��y�Z�&�T���	�vS�dp�Ϋy���a���XyJ~�g)�M�'9Hahǣ]a�d���ޣb�6L��'4�%�o����*��|�_��Sǟ�j� ����thpl�8e�l��"Ú��l��ԟ��ZyR�c�V"&��<���^q��X�NՀ*��G��?�(ċ��b�>Yоi��7M�$�'�"�`shB8P�2'�O��2�O�Z�K�k�T�#e� �?9d��O�Dx�o�B���( #�!�۷B�ON�D�O��$�<E���'Z:d�%�@'*�Pɡ��t��eJ`�'�>6��#8R���O�4l�Ӽ��
�B������%7�t��7��<)��i��6-�On��A�y�X�0����/�V��֢��O)"eϚu��Q������4���$�ON�$�O,�$%b���P�eAX☲�%�w/�˓^�EE�,z�'���$�',]9�҆	*�Y��Q�*�i�wð>Iv�i_7�}�F��	��� �4�;N\���lP�5Bd)� Q��	�1��c��'�&�$���'���bD�ƟU 2ds'�ǝP5j����'	��'a����TT�<!ٴe�T�I�s��� �-��Zr<�I��}e��!��6ɛ���Iv}�s�v�m���d����#eS2�r��؅@�:AS�
�<>|amZb~�M�(z���\�',Qk,��8��=kB��"_"I(�o;e2�d�O����O����O�$)�Ӥ�F|rv䁕U挔�P�ҫP�0@�	�h�	�M���R�|���;����|�ܬnD�����B-�h9+4�ʚj�<����Mϧ>*R���4����9�%��OV�`%0�Ď$wn�*���?).6���<�'�?����?	�A��� ōפJ�My$S�?����$T����� 
ޟ��I�,�Ol=�o֍&۶�R�!P� J��i�O�-�'��6M��ϓ��O���cEǉ=�<�$��n9���V�^ �a����4��x��'���O�ff�=iQ"E��!��j�L ƫ�On��O����O1�P�Q���j�c���4H
;�NL
�Z�Z�@�8��'���fӶ㟸;�O�lڗ>�P�YG��a�� % �7�D���4�?�օ��MK�OଣR�0�
I?!�� ��g�v��"̈-�Դ�2�s���'"��'"�'32�'��ӛO����MԼ�|�v��g�L!�4@���/O��d,�I�O�}oz�=zTc[�[�,�Z5��=8��d�ǋ�MW�i��d�>�|��b��Ms�'jbd�A�
�rݠ�j���A(�'\���̟�谟|\��SΟȻ���=7�����}�(�K�蟐�������my��n�|�Ó�Oh���O6�x�d�+��`� ]�t��9�!�3��3��d������4�y�Y��iW���hxx�	�Y�AR�*?���_ep-c��Q�'t~����?)�΀zQ�����I0���C_�?9��?��?���)�OH)s3m�-t�8��s�̼,�|����O´nRs���ϟ�޴���yWnš9� �q�C1B&��hui�$�y��i��ylZȟ�v��Ϧ��')��cEP�?��M�	:鼗Eh�A�͝$&6���N>I(O�i�O��d�O0���O>y��=dFj�"ŏ/Y"6 ��<��i�j���'�B�'��O��!�	&��� Ά?1n��s�K�0?��5��
x�r��r�O��u9�G�&�hѩGwk�kď̀{�4-��O�m��[�?A��;��<�/׬f}8�� ;. *#����?1��?���?ͧ��D
Ȧ�r`�Ɵ��m �8�B�����8��{@K���d�4��'8�ʓ�?Y�4�?����) ����DȌF� �g��3/��\R�4��d�%^�<���'�O����"��8����2HH��.K��ʟ��Iן���ݟ���[�'<�]["f
#�����@�$Tl�L���?Q��?��\����'gh7-/���X�ΰ@c"�(L�r%z�hč~\��K}��q���lz>�'�LҦ��'��I&��J)�X��l	~�,y3B4 Lp�I=j��'�i>�����������
��-�'�K�.��)�I��l�'��6M�)p�����O���|�s�� ���Y����0b��u~��>1G�i�J7-g���~�� �/�N��:��E�giW�<��bŃ�z�<����������|���#���%�T�C	�%��`V�O-�'���'*���U�\��4x$�` �KG�;�����!~1,T��jK��?i�~a�V��[\}�uӠAH�)����q@�	�e��聧ŦY��Ŧn|~��N�X�><�z����O=��i� cz��q�+�pz�<9���?Y��?a���?�-�(5@�	��Iy���a��Ix�y�G�Ŧ	����	�t&?��I��Mϻc�D�{4�# xY�-Q4w���9Ŀi��6-h�Lק�OSb�V�i}��"0� ��2E]Q̄0B��� �
M��4�N�O��|
��q��ʔ�[t�4-nS��`����矔��UyRhw���+���O����O4���^]�ԥ�ࢎ�rKjM�R'2�	���$�OZ6Mn��'�����iϐ(\Ƞ"�b	:۠���O��ASb�>]:.@��)Ӿ�?���O��I	�$h}�P�N7hF���OT��O����O�}���'�̱�P��*W捌KF��~��&��C�R�'nJ7m&�i޹�熘 hJ�q��%�Nt)&(b����4͛6�'H�#1�i���%\L�1V�OM�c+�)B���.��O[D<�)�q��_y�O���'5B�'�2ÿ^6" � \�+�� }����M����?I���?iH~B��J�"��D�t���<E��u�X�$�ߴ���8O#}��Ð=�}�@H�?%��T*WK�:YjܱW �s~Ү��'V���ɼg�'W�I)t`v��w�74m ��@M�U˲��I��T�	ٟ��i>��'J6��	dXL�d �on|!bV �� dz顡 �?U��d���?��X�������I�)L�*�H���Ƹ�a�*�X��B�Y٦I�'�\ia	��?��}���rك��28M�$�uŃ�`�<в?O��$�O��$�O��$�OZ�?-X�''s�D�A��*x� 7L|�I��$yڴNo���'�?�W�i@�'�)M	�R:����w� |��1O��Nj��Fb��Y�:��7�$?���!(�����iJ�'8�*�#��O���I>�+O�I�O��D�OH������8�U!4X[f��O����<�i_f����'V��'-��![� @�LPL�����ĄU�����ɤ�M;@�i�D1�3� ����V�a��8�l8���䋸.�ఠFk���i>Ii1�'!��'�,�1N�=�0���Y9/g�db�aFƟ���ǟ�����b>ݖ'eF6�ԲB�90��N��삀f�9K��1�!�O2���ꦅ�?y�[��4"BI��HV�� � �OHP �!�iV��ێ#ʛV��xA�+�#wh��~jA��P\t9��T�w�	�@�3!z}X�ĕ�v�v�i1朕�����׊{t$�˖�Q� O��Y��=5RB�P�툹&}�h��֠ sQ�&C�V(ʒƊ͠�� �7YfْU胯2UԘɶ�������pĕ�T����"�5X~����f�섋�-#>Xs�dո$|����IL�A�>�ɀs�Z$H<ԓ�$[�
<�� �_�e/��V�K��Em�X�|�95��(jnX�Zԫ[��}�dHQ�IwT|B'S�_�bq��n�D�,Uy��G;�-+��� Xp��eG�&5I�A��%�7�O���O��	@c�i>� ��Eр���g�=)�Z ��	��M�_~�X��'?�ğ�Z� ��=�J��@MT����Ͼ�M��?i�[,f����x�O��O�EY�JHz���B�-N*MȚ�\�ԗ'�(�z�y"�'��'�R���ߐI8����j1l�H��b�w�F�#{��`'��Sҟ�Ily��0����H��9_tCrl~� 6M�O�h���d�O��d�O��|&jmx�)o%��YƏ"{y�m�p-���'���'$�'��ɥ	� {b �W�I���/<�9�@#�I�p������'�@d&x>�H��F3JFRE�"�[gהIwb�>!��?�N>)*O���[����L�f�T8׊����[.a����?y���?.O�MIb��o�2I�:��2
�3f4CT�-;lՒ�4�?�O>�-O�=�����+M{:MX�N�;7�B!"�DH'�&�'��V������'�?�������wc�C�f
@{v��(�p�Ty#�	����S�=�ڨ3  ߇ �8�Z��x�V7��<�D��
EÛ�h�~������fD%&�}�d�!lN��r��ʓ`3����i(��i�Z$�@��F�A4
��"������de+�Mc���?����"Ҙx�Oc��q�Ї"�����\���遦dӸ]�搟��'���y"�'����K�����d��#e���#d����O���J¦�$��Sş@�w#
H�g�<]�T�A�k͌5�VL�'_�	|��c��	۟��	iB���l�$z�~!�EE��n �ߴ�?�j�/����4�'#�'n>$�!�߰4�P����������>�gk��?a���?�-Oę�զ�O�.q����O�@�pnվwlz�$�������$���'���Z7�ρI� كRc��Pn~Dy3) ���'E��'9�Y�x8�����BA��ʤ)�`J�p��O����O�O��	|(�'7��ȕnD�C ��(C�� (�()�O��O��Ĩ<���;if�O2ri�7��#Ƭ��sa�c�x���"tӦ��8�ĥ<�# YM�' 8�ӴɿW[��(d�O2'bP�o��p�Iry2��t����d��kL[�kp��C'ƈbͬ�HA*)Ӊ'��	�,�V"|j�O���8D.� �L�*�H��޴����~(�MnZ��)�O0�� d~�NP[}ۇ�ϖ"�*�U폅�M#(OR9	6���'��禙鷤ܾE�(�a�ǎZ�pUzw"u� �:��Ŧ��I����	�?�H<�'0�h�"a�4�Q���T����3��i:<��Oʓ���<I��^r�@
M%.樚A �y�����iR�'6�Û�2��i>���ןd�A?��-��&( �K�gH�-�T���D@:��U&>���ş��^�"��4(�yk�h��0LԑmZ柤;�`�dy2�'���'�qO�� O�?t*\�flҚ/��z�_������l(��?q�����O��
��XY^��;1�^�,�V�5ɸ=��˓�?A���?9���'F���*��3j)�%�g�4Q��[�hV\�q�O^���O�ʓ�?��������6[ �iۤ�S�r�Z�� �M���?����'��շ�t�@ܴs�b��1뗷|����C
qE���'���'L�	�<�3��|��'������iцl�� �b�j�(Bw��$8���H��P<k�tO���Q��]��D��!�h9���i#�Y�D�ɜ''PؔO?"�'{�t���Rn
U�Ѐ � Z.�� ��(�c�D��Z��EңN<�~����GJ��� o�RP;c�[}��'�j��'�bW���CyZwKlI�#H�k��q[gb��[�Za�Oʓ:H�HExJ|ʄkR*�dЊ�T�&�:��ۦY"Ŋ]ß�	�$���?q�����'�bDC�m�0&]��h��b	� 3'`Ӧ5)�DԬo�1O>y���99��%(�<!%������D��U��4�?����?��5��4�^���O(��5LJ�u
§m�D/Yuv8���Y�PE��	����'���O�I��4E�=��̈wX�5�i�"$I8'��I��ȟl�=qwʍ&.S��JL�.y9��ҭ	A}�%a��40�O���O(��?1��D�F0H�e�K�6<�|P%ϑ�|��0(O��d�O0��"�I�x�3�N8�+Gg�ΰ�6.ć<�Jm�k<?���?Y-O��� !<����T4��B�-s�a�V�<�t7��ON�D�O��L�	3e�N�)R
zӖ̑Jɷ"pL�B �E�d;:��\����ϟ�'�R�?]	������EF�q�rp	�n�8���A�i׷�M���'�
�9*�Q�H<� �t9T�Igv1������Q��i�BQ�`�I%W��Oj�I�?]���؟(��L�v*�#)I�� ����'���B�W�\Yi�y��*H���,e��aa��3Z� [�d�ɜp.��������	ԟ���MyZw/�t����$)Z9��(�?K�(���O&���?Tk��z�S��` 5Ɖ�/9�d�3	ˤyn�#K�İ�IПd�����S_y�O�b�&��x��-.�j�b&�ަr�7MӸ�B�4���;�O� &`&Qk �F��Θ1���M����?��{�$�(O��O.�d���"%lL'3��ф��>Id�V�P���''�H�4�ħ�?I��~���g���U�G"}�I�",P�M3�it��,O���O��1�	�th�� �����0�MFOX�&6�<q��_y~b�'S�T�8�	�ZU�`�竂�A��Q� �B�8��\蠪Ory��'lb�'��O����T4Ĩ�5���N�$�h0��N7�0ƥS�#l�	֟l��vy2�'h��Aןra4-܄5 %#��O� p0�[��i�R�'����O�����c���	E36�L�i�� V\��a�B:����O8�d�<a���t,�����i]\y���WA0�+L�
Si4�l��@�?q�QU9A�O�I=�T`�$�#�����N<�7M�O:ʓ�?C�����I�O��d�����w�S@��'0�qvo^M��?�0���"��<�OXNa�"�>㺼Y��79d�O��$�O^ ���O�˓��(O��?|`x!q�T�(�$3���:�IɟdY�C[�{K*b�b?�j!F�%٠|r��2I�ݸbD|�HxCC��O����O����>��|:��&
zP�ݤ'�.q:u@=(h֨Y��i���[�	���������/�脁�ٹ.�=��&�P�nȟ���Xb2�Qny�O�r�'��
�jL�cEc\��ԘKQ��v�^m�<��.=	/�O
r�'D��;%�Tp�n�,qX�}YMIm���'^��5_�L��ҟ���x�@��6���2rmpa�ɯ;͸D�'��zч\�����O*�d�O�ʓ3��ӣ'�$�p*G߽+�X�Kw@�1Ay�'R��'��'S��'���J_H^����c7V�P�	]���'�B�'�R�'��'�hS g}�f�K �R7;9HP/ޙ �T���`�}�	��$���I�h�`ȟ�V����	4&��"�^ac���Ms��?����?�(O��A�B�Q�$�'OXP�(08���$I��*&Z���c���$�<9��?A���Yϓ�?a�'�r�5�)� ]��$�Aߴ�?������# ��OB�' �T�ՍPqLq	7g��=&d�V�A���?I��?	F&�<�+Ov��dO�?�O�(`F܋���
t����`��˓^i�4��i���'aR�Oy��Ӻk� ߲e�h�@e��]��T���Ԧ��IퟰrrD~����~y��)�G�vI�!�6\+���b=>:���\�iς6��O����O���P}�U��
�j��!�<�t�ÁC����Ǌ�&�M�c���<!���*���$"�P�(��Dj�,ͳ,b�!�©�Mc���?9��IGHP��i��'�"�'OZw�B$���ڧ>�\*0�$V��!�4�?�,O��d0O�S�l�Iԟ �l�"V�&lHtcA��'��M��9��((W�i�b�'�"�'�
ꧤ~��h  y�'ϧN�PV�ǀ���N?l&�$�<	��?����-+ݞ����
14U$šu��N��� ��y}�Y� �	Iy��'���'\L���a�W��`�cFJ�C8��8����y��'d��1L$B�'��ɳt�2�OY�l2�6�9(�*�;� ܴ����O*��?��?�GC�<�dYDڦ(�Ѣ�4A�8��k,\�	<i�ƙ�	���'�jQH�~���D���g�<"&��Z�'�d�YŹi�rU�����d��Μ�	����_� f�25��@�/
V,��n�ʟ���uy���
��?����Zc�̟Cl֔ኍ�� 	�!^���Iȟ��	ПS�jg��$���'$v��`reʹD�v]�����=n�[y�(R7M�O��D�O���j}Zw���uhI�ҕj��R�^ٴ�?	�g-<��e ���6W,��}�3b��8pl-�´�>C�gT�(	��!ǉ87�O@��O��)�b}�Z�L�rm��n������;�"�XfAX�M;���<QO>i��t�'�}��Q�:��d� hhD�M~���d�O����g�@��'��I������	�'��"p "���%7b�=l�����'�X���	�O���O�	pd���Z �=��bN�E�lP:��ɦ1�I#t�\,2�O���?�,O����p9
�o�3倥ڵL	�k�T��R�x6'v�L�	Ɵ`��ʟ���ty�bX��)�uo��S���^Y�eF�>9+O����<1��?���m����g@��)�#�k�"0]�,Sc��<���?����?Q�����ʄ�̧S}���� _7H����CK�L���l�py��'I�����	ڟ\R&�~�Pf��<��ڤ��(>[2<�5�Ǧ�����$��ӟD�'�5�D-�~��pބ�3ak�')�r���Iϳ`���#�iGT���	ޟ�I-��	̟��I�$�Zpb3n,q�jj� �[o����B�Ƛ�	`yb���it���?���b��'U�|�V��D���2�&N��	�� �Iԟ쨠�??I,O>��u��AW3M�h���ɢ
�7Ͳ<IA��qO�&�'�B�'�����>��s㒹v��ly�A�'Hlּ�l��əo���6��9O��>� 2�ib�\�T�~$������L���i|b��FG{Ӟ���Oj���e�'-�I++Xpc �/*�BS!Gð[ ŻݴT@1Gx��	�O�18a��E2�h�����X㴯��Y��ӟ��	�X��U�O�ʓ�?1�'��M3��Ğm/8@K���7�e�4�?�+O�i��9O�S������H3��B�,^1�U�>g�t*a�,�M��nŞ� Мx��'��|Zc�\L���`G8y��O�aؠX��OA�3��Oh��?�����1�@��t�Ҵ7	���v�;F�1��'�b�'r�'�r�'	�]�&��+3��X�6j��n�*E�pȇ�@#�'�2�' \�XS�������7r8�Ĳ��'o@`c�Eܺ����O��$�<����?��c��'BRt��HW>X�ҌX��ڊi�6(��O����Od�d�<I���e�O\&�rMQ��}�e�C;<�� �"a�l�$>���On�Ā�#��D'}b�Qg�0z��N1L�;��5�M���?!.OD��@Th�����Q�Rb)�<q�z���Øt��\�M<���?�lB�?�O>��O��L#
�/pJ����uVji`�4��ă�m�|�o��	�O�Ɉz~2�ԯi��`h�OSd$ �%�O�M����?�֭���?qK>��dJO0<p�&�5B�s�]��M��J�Q֛��'��'����:��O��s��,ba�����> ���Ʀu�an��&�����>����a��F�@���N�( �(Q�i��'�aҊ%�fb����p?bJr`��bǑ��H��ʦY%��SA�U6��'�?���?�R��7]�~�sc���	�$8�Ç�-����'~�A���5��ǟ�'��Xpж�q6��)&ER9��(mi>�-�m�����OX��O�P�D���GRXQɉ��5X��^� =�'��'P�ʟ��⟰���ÂY0\���#���*v�ėeYD�eyr�'kR��̍�����K0@�����\���ו jh��?	����$�O���O
9`�Of�:���)&����<�D���[k}��'Lr�'���#fː0�H|����$�F�&��9�\��@ۛz����'��I֟��	ڟ�*���\�i�e1�D\��"�� A�`+����hp����O&ʓ}(�����'���E)zh�,��iD�o�5�V�Ȟ_��O����O]9aI�O6�ON�qO.哴F�Z3BM���7@��T���"���M{.�����XA�'@a�7��h�����F���Y�ڴ�?��VB������ݸO�ݙSFZ�dU�]�L)Ǣ��44�Lˢ�iR�'��O��O��$n�f�!�k�"���a�ƞ:O�Z�#�4?��9�B�I�Oh�t��u��=��J<x7��2L�٦E�	��H�I�E!�	 K<���?��'�v�P�cS/-���-�&!�H���M�I>��%O�qG�OB"�'��C�1�yC��M�;��rA�y~6�O��ۣa�W�i>UFy"��	��@#'�Į,�;�����̕S���<���?������-ۚ� L=������.7�D�࣭P�Ɵ�G{"�Oxđ
L�=(NZ�p���i�b�'dR�'�r�'��5NHH��	�`���	�Mv�c�)��@n�(����<%�,�������U�7�6m@�`Wz,���oҾQBBIT�M��	����Iڟh�'� �kq#:�i�vI��y���?Z����Q��< ڞn�ȟ���p����~"v�B�R�S'��33�(Ջ��I�u�	��I埼�"��}��'���O�p��ޙX��ȷ�Y$�
5 �1�D�O����E= -���T?�K׫�@�\ @��-�E�a�x�T  hq&�i��?��'��ɐ	⅛7�Y�=�n��SM6�O��DH�PZ�b?1�t�����ҁ�� �t= �c�>Ȃ���i�	�����?�JN<��S.�3��dP:̉�J��k��t��ixEj����`�R��q�hM�2A PX&������M���?y��Z�\1ش�x��'���OF��$L�dBV�ia�U&�d1�d�?m1O��d�O����0UJN�x5��tF��B�U��Hnɟ������?9������!�Q�T����1 �M��U���]}���7��'�r�'��_���E)Ů9�@�Y��ҟh��C���7�P�K<����?�J>���?���޶,�j�0BC�q�{c,޺Pk�M�<y���?�����䚖R꒠�'�(L "N^z�&%	tE���'�"�'��'�2�'/ht�O*`� �b���c�fy��$X�|�Iʟ��'B�J,��)�O(@�vسh�̽�U�ч�����ۦ���u�	WyҧZ%
p��H<��)�K@���1�B`�j�զ����8�'�|��1�	�O��)�-��'Oq�� ����h	��$�P�'��)Z��$�?5ba(I��x=1B-��`vd �`�h��u�R��i���?���2��*U�~E����o����F��\@`6m�<᦮ g���O��ă2��	��Ʌ�%
�p,�شg(��Ǳi:R�'I��O
>O�������*�'m��҇`S=	̈�o�9?~#<E���'���*D�ա��s1i�$����Ӷ�$�O"��6m!��'�H��㟐��{bB��BgBjF��脬?GX��>AdnL̓�?����?�� Du��ɂ+x$��II�M�6݃��i�b�E�c	8O����O2�OkL�\N��D��7d�P)�L��i����N$@c�������	ay�L��M�l����[Z�Tҁ��x=���4& �d�O��d.�D+}��D�I1|E"Ch�v/�lS ��
��'��'�Y���r�װ����+1�4��B�i��9�� �����O���;��<�0��G}B���Yh�g�%u���`����O��D�O��3�(�����f�J��$آb]�}q�BT5="�7-�Ot�OF��d^ �� B�fЬ4�wh16����'�\�HYG	*�ħ�?�'(�q�Pp�j�b�fE5+,���x��'��@�\�_���2�앣i�����4��v�l@o�+����O*���t~��ŲX\v�P��*z��a����MS�'�: �Q��"fSrt�6� ,����4[b$�J�i�'+b�OјOP�Ę�Y *;d�TZ�^��᫔�A����	�#��7P��r�J�W���M����?q��<�$x��x��'�O��VhC�&8Y�,��ɴՐA�'��'}��g�$I�af].ft�P����T��7�O!��̬<e^?��I]�.IJlM����7]q=a�h_�aI2���Ox�����Lq�<�U#'擝2���Ifd�&I�d ����&�dC䉶p>b|��(�?,kT�h�K�e�l�>��c7>���"D�@�(��&�T�z+Np��Vw�꩐��1D���[ �(T��&+�c�fA���t`�"��][�Z��%�+p�(@���6h��E�\�F����9,*^����R�[��՘�f��f�b�#bC��� �0-ԗ"���H2O��#ʟ�m�t�V�Q0$J�#�.V	 ��+^64�A�I����	��
�:Ј�/'�1*Uۇ: ���Aݟ��S�!� Hb�K�t�>��創y�$ "�Â���E�_	t�ڬ�7K�;G8\iA ��g�9��剱0�x�$�O��?�j �N4K�a�U�>e~�*��x�H����V���x��˙cLR՚aᕶ
�P��D	s�I"P���K�Խ<;,� e�#9�~��0���˯O����|�"��%�?!���?1��#��"p.ֵR����%��[��K�/"5�"}���j�*�
b>�D[0(M�
�����_Hā�D�lD�� �A�\�D&�ş"~�ɪ_+B��㧊�^��k��N<x�"T����w~J~zO>�Oґ��գ�e�/�b�a�S�<!&�?)��sSN@ˀ�0gj�P�'�"=�O0�ph�b	0��4Q1�F	�T�aT�' �G��nP���'8��'nb�vݩ�	ʟ` �*��$��A�Ձ�2�l�ᢡ���?�0�Wos��`l�{
�3ړ�jT@t��+������F�pN�0��'�$m�-�>�(@SF{r��n�	�&��*1��!�ت�~b(��?���hO�˓20x X�I�v�~��4�0t}�ȓ4�� X'�'aj���s*̂^����)�.O��s5�MݦaH��Í7��+��".2yy�`E6��O����O�Q1Q �OX�d>U���$%�<xa�\+GA�Y��R�(h85���$�1�Rlx�tx�&B��ܩF�:�}3�ݕh�\�B�M;X����P�nx��Z�M�O�����߆E�(���xb�=��������� ��M�Xm�!2�#rz!�d�j��}��ԮXL��H:pw��X}�[�xӓc݁��$�O�ʧc�D�sH�^r�ɋF��jU;d^��?����?)&$�)t�8ŸN��l \A���e��S	 �x��(�<w��$�I)�h�<icȘ=l�Ă��U�!e��[�I�I����%���@�N�W�Q��bk�O�oڀ��OclM�#���4�j1Q�'�
���h�'T��'D@9p$��g(Ƒ8F�Ћl	�s	�}z�'cJ�h�U�|(�9�šӜ6��ḟ'��"~�<���O��'Hi�Ղ��?�J�"��ҫ��/x!a��uĊ #ČL ؞����߉��T>!�|�ɉI6�d 6/��G��!�1̝�6DG�P���Q DU~���'Ǣ��4��%I�Ż��װ�P�wlکNeB�q���n�G��9�j��a�A�v��A	E���M��?Q�t+d���"�R��kÀ�7_d"�Exd3�Udd�I��ϴ��ӈ�.�>��B'?Vg~HI��?y�`ܐ����?����?�RW?�I�	�
u�YI�����58�$Γv�F�ᡁ�2m�ɒ �C�'}��!�c:����CM��_\��I�a�F~�Р,� ���Uև�����OmT�r�Rh�DHr�� �D�,!WV�����t�'m�Z���́U�N8k�A� *�u�Ԡ&D�|)a����ԤP6�з� �(�M(�HO����'Q�I!O\�\!YwsU���J�6Fz� dh�%>r�X���'Fr�'�"d�;Zt��'g�)̽1R�'RB$���0Z�z�D�1^�1!�D��ٖ'�n�
���5(x�����%2��{H��	�� |Ⱥ�叝f��`[.�>��m'���O:��'�)b�i���x\� �Y�]c�CTv�<�G ;�\�"Ck�`Pdb⃆�<�U��'� p��Ϋ>�����)��~g�kՍ�C+<�����,kV" "p�OR���Ok$W=��H�+/-���)W>��iJ^�vhv"�E����6B� &�Q��G�i�6	eD�E�j`��?��C�U�f�z��`B%J���A�*�w���I'�M���)̨s*��3j�c�UJ��\4 ��O���dK5Sۀ+�L� Y�5�W�D�"a|�G.�d\Bz�����;(?��j (�H��K�M(=�'�^>9 ���ҟd���C�g�w����L�F�e�pO�5UH]y���X���kU]=�?�O01���@����b lA�05��3�݌h?�X2��55��k���t<4���O�ٛ`��0"@0��	q�1��_<������y,O�O��\��HŇ�
��0c!/;~��T��8D���ƥ�=���
��ǰGjĒc������HOZl؟��.�;^�z42��Ǘol�k�AUEh<i	�"�i���$F=D�B�f�<���=6,@u0��٢Jc���IHb�<aF�U@�P0����8ovI� i�<Q%N�F<	1�1M�LA
&M�e�<�Ăя[��ј���/b�nh1T�_�<`a�/	ZXxG	W�l���ՂMD�<9�e\�h"�1�6m��{���W�<���X�t����J�	OF�UȜQ�<��#bH@=�ȓ	�:9�5�d�<� �Ծ}��@�B��oJ�my�^\�<QQF��,O��P��=�x�At�[X�<	���a�y����U��wR�<I�!ԙFM8d(�IF�Y��I�<ia��Z�IS$��i���&�l�<���F�_�8m��@��c�d�����g�<��0=<� B1��lr�LӓHd�<Y@�R�ZU|�A`lMv0B0S!BJ�<��G��
��M���ǭ(�|�:`�D�<�⥘�4��@`�$l-ޜ�1�i�<!�cT^�����5;ءe�~�<�B�&sP�i���2禼{W��p�<IP��6c8F��ě�_�ڀ���j�<�g�
�Z������Nc��aAo�e�<����X��H���~�>x�b��a�<�T��$2���)\	C��[1��^�<�Ѧ�/���Y�܂$q�#��V�<9�F�.$F�P��W�G
6(x2,�V�<���+�
v���`��BJ�<�B��F'L��"�M��:S�!D��`��)��YB̕?s���( � D��GDC�0���
��8
|Ey��(D��I�%,"� �s��!-�2���#D�� ��[7�Hs��hbD� n7D�PkL��J���)�eJ%?�"��,"D��[�J�? �Zc�I�4�"Q�2}���F�Dh�A�E>���"T~2u��AL�Q�d���/D�,�"�/N=�TAn�  �Ă���j���' ���&��Ϙ'���S�G2	�r�ׇs�XP��'*��Q�`�37��Ș �� �,h�l%�~�Cμ ����iT�4���ݗ|�f���C+@'��(Q��U"�zR�.3Max�NW��։P���r��I�`B5��.'f���f�5�:�{*l}�	���7�:؁q�'��̺%����<�:�*�A��h �O x�q
D�O
���D��<���94.	�J#���A'�S�8kE܊i����UӂO8��'iD� Xb���(�\��Қ;F˓$ �r3d�j+nH'��?9F�S�։λ_Uȁ@S�O�U�<�#.�/b9�؆���Ȁ��fly[SM@�H��xQ���ON� �e�����<ݳb� ;�lxY/��I�/�ȵ�G��N�@�D�
\��𤅦��(4/�e�`*�<Y� �6g��\!��H�]��ٰoE���i0���'f�
��aF���<9'��%2U�Yr��y��1�MDs~��Ts*��g���&g\�@��.��@���]n:�kpBȅ�� ��I��	V��CW�L�||&���$4� #��n���RC*ܽXp��0R��8�g�udB܊cW�%�  ��#1F��ӝ���4i����e^-d�����U:��1�%����m+@�� $V+�*h���*>��q� ��. �Cê��z�:��u`7k�@��,FTl*i%��h��@|�%+�N��u/ O��W$I�4
`�z�K88�F5�R
մ/�]��	?@���4*��@��L����N=1�(��-c���d��;0Ȅ���D�9j�`XV'�.��I�L��iô�^(����v�4W.���K�$hCz�����O�`��BJ8m�l����]��* bҹ��x2�0c�Ъ�ÓnHy��Hʧz>�7N�2 ;d��5�~r��Q�����'w$��2��B߼Â�ˉ3��ݰWB�$<���*��Sc<����)g�A�M�'%�Vl��׾0��MS���j�9�kQ"F���/
<(۱jK�<�5(��M[�*��l1���,"���+h��ao�#S�v0{BnOP>D�@C
�=	m������K ��p�N[C
��T�Y�oq�a� 
M�����I펕��}�O�"���L�4nd�2FD3qp����O���Gm��"j�i���J�RU�kΜ.x��D�>Q����r��P�Ċ3r҉㌉�?i��ќ
��O?���*ץ?8V��`d�q83� �_+r\��k�)H�!Y㠟��'��l�GL J�w�@��� \�LY'큔+�pQ+�O��N�AX�� �cL�Fm��P�9	Ԙ�sY={ה��;����+ʊ5hw�^�~ȀJ���O���"�Y��y9�Ҭ`�L��Kۭ!�|L�8Ofrh�Zn��kʀhE��Ga�1u�F���\��l�Q�6��QcԽAh���1�݆Y5�d�19V��>ͧb�|]�W!B���4�&VT�ĦO�k �}=ɢ�,F)>.ɩ)�h�A����� �1��1c H�.����lU0	��� C�$0�T�R W��+���< |�	#u(tv-��Bh8�ȇ X$�)����d��˞>ߠ�(�d�+�^�y2�aq��'r6�;!Z|y�\r#�ôi��3!oØS �'�>Mi���)߹�1OU��\�s� ����N����V�'Ejh)ƠJ.�����J�7nN����	Q6O慊bǖ�k2퓰lA�m�Pm�a�IȚ���z�O$,j��O�˨4�
�8=Ely �'H�܊�*[5e�TP���O?%�z�Q�'O̱�2 CR|�t��$Q����'�0ؤ��a]VUx4�Ώ~���'z�ՙ�E�*F<5��dX=4P�'�*"��'�B$�r���N����'���'
|�n��P��1#v���'��j���2
�
͘�*�#'[�%�
�'` �b�n�o@n�����N��u�
�'��lJ%JˋZd$��S��7NQ6 �	�'���!��9oђ����^B�	�' �<k�Lɴ<�r]�F�O4PI�4�'�zL#�	�B 0�v�ُRXu��'���X�o�R�[�N��p)��'�ʠz#�+��s@Ǚ%"$�X�'���˂���te�����Kr�S�'��@�6����`$�$�e$%��'e�@q�/ުMKja����b�(�M<���έ+�TqHt��,��5iHo� /V����
Et�$戩Dr���ȓ-0 D�D� �F�� [�f�����A�J�p(d�H+5	��+VO�[�g�	:"/�ِB�13C:Q�C��r�jB��	FǼ�p�Z�c��dA��#)"�A��ǰ�xf�L@"pҢ:,O������v�&�yW@D�KX|���'�Lm�s���=�����67;�hq �E&7� {��\�is���5Ɗ��x�͈P��P�#����ӑ څ�� 7�'# �g�9��
�Nt�a�~:w!�$�$b��C8��墓Y�<AV��mV�`xK۪&���bU`]||��%������"�k&FU�~&�bF���k��XW�Q�`J�(%!��Q���.B^���#|ܴ�C��*T�T�
��Ăp��GM>��<�&U�0i;�*/��kS�CX�@���QV�{V����#��7I=֬K�\�M�� iG
YHB�I3�|BE���h"M���y�(Odڂ�(K��q(& ��G�X���)�r�pY�Mʭe�T��#D�_!���)Ѳi:�F�8�D%{���z�ڒ-��GddM��HU�2���W��x��YƖ��'N5�P0)����x�`��XD�U����%Al�T�&A�0N�I��D\�yRDFIh� DK�S�? �.�0v%�q����T�Z:��'�Z䣔iP)n���j�LX�ek�ap�k��Y�>X3�l�,ZrHY���x����u��Z�,P.�`���$�ē4T���+�M��TQ2�U�Wc�%�~M��5D�Q��<⬭2�nDf�<I�� P�|�Цc9M;�b@JP�P� @��i2汓4#�(�u�~&��������,�'"Fv�*-S�$$��y��Ӄi�H[�mJ�}��x1ѩH2�*�V��QѶ��W�����d��A]`�����*�6�! ��-&ay��5]4M*� ��_D4l���? ���`��3[�e�Ó-��C
�'M�`�%%D�w�^�yCi[6^,��iJ<is�Ӵh�HS�����un�I�'c�|�� [�sa[-[)4Ʉȓ"T�sd��m����s�.~Q�$i�E�2C�ꀙF�Y,8������OP�g≢Fd�&/>n6��"g�\B�	����K�g!s$�
C��!hb˄���P��O�pd	�b)���z��P&K5 _�]2k�>ay��M�nH�(��dךt��¯ݪT9����$
j�A�O��
�'_2d���Ad�����cA9FM�سJ<�'�ƀv������J�h��hl�[�Ӻ�U���V���UV=H1C[}�<�"��j��(2��w��x�W&(�� 覭_�&k��8w�?�yp���y�M�HP:�u�O���@�J���O���	K�9�~��|n"��e�T��.n��eӚ)ܤOL�j���1[�i���Z�(�:��P�d �g�x�y���(�NM1	�!��V�3��R��v�i����9�aj�c�\8 ���4�x��2�\�/)�)��Ʉ&��A����/����I XЀ�?Nn�H7$?Sݸ�{:�I5j�p);�Ǳ���<��B�B�1p��	S��w�ZVˆ��	�a˚5��B$U�,H��ȼ��䊄L���U�i�<hɂ&ϕ3�|шyʟ"�[`�V'L�kL��u�Q)u藄(bUA7�\L8�H�3 .��҈�ܴA��]3#�F�&ܐq���Y�@,$� ���0l�2���onT��P�:��S�43�J�83��bAZ;{X��I17�t�s)^(��Ӻ�'�����W�0����Q�b)��蟖Q�<Ͱ�(!/3��Y�*��9��IYۓ#�@keE7��-A1�H�
>@'��b��l�`�dl����� 2�i݅[F(� �>��P*
�A�6D�Ĳso��@8���I0 ��[aLW.?��IJ#�l�d C�yʟ��7켣���*<8���D�f/@�ر��^H<�$*R!F��0�]*'C�a�lM�]n�'F���&#٘Z��djD(ؠ3V��}�Ł"�(���0s��4jl8y˓�¥���`��0r
�	L.ȋu�T5@���B⍿|X`�S샾\ZuC��-*,�؇퉞x�f�I&E^�J�����
�.KC�ə)ov�ҡ�i ��уE�#�C�I<Y��\��A=qSt��h�/��B�ɹ�}hu��4�F��j��Z��B�I1R�r1���dSP��5J�"oLB䉗�8H��	�,��}H��QC�B�Ɉ�؈k��B�1ұK��	 �hB�	_�<�3,U�1�t�Ҕ��)%C�	�f�)� }�f���P�/ǜB�ɗd�~�J��҆M��(��
��"O�����?�Xu1��ش?�qg"O��Ԁ�w�LI�K��X)�"O8��2��1���i�l9�c$
�y"�Q>��� ��7V���L��yr��64��&�0*`�ћfgL��y"��*����Uc�,%֐�PGڊ�ybo
q���%��S��\Y��F�y���!49f���JY6��7�6�y2�����p��Ĉo;d�Q�@:�y��R����g�R1c,6Ͳ� ��yr� 1W����f�n:2	�$�"�y��� jGԘ��A�d�dmy�Z*�yң.Q�����H%Kx��CC@7�y�&
bz��`��4Ő�E���yR��<:��%�u`��2>V�ˡEӓ�yB٤=��0�� ��̰q��y�lňOOF���\���Y��a��y
� ː�9"�TJ��� `��q�"O���e.˹I�j�H�6I.�:�"O���G�39\���C�S7�l�"O�Dc���'A_<Z4�	O)�TP"Op�	�$�;USB⁆`�v r�"O~!j�B�BHlX� a��M��̣�"Oz��\_��$KO<O��BG�n�<)ժ��yE�H���ϻ� ]rq�A�<���/��0##�7o��h� �t�<�K^<����&'J\
�T̆e�<��KM?Ύ=�F~�2���{�<����?  �! L�sT�ɣ�Q�<A��@`�Ġr�X�H���q-ZJ�<�P��i��|�S��1RB�!��ȌF�<�QH�����K�B� o،gLH�<i�č�D��J��Ĩ2#6�Z�C�^�<D��},�2���>�ŒWWX�<������dAe�`�J��`�Nl�<ٖ+U�3�~q{6�V]^� �(�d�<�u-�o�:0re��c,��A�
X�<�R��)*l,�g��b����C��k�<��ƃ�`�1C�@d��+v��e�<�RF_�����f���>���a�<fgU6��9/H�fqE'/Iq�<�׋�?S�"�*�QS�Go�<i� ��K �KV'[:ʒݙЧ�i�<y��a�]�����)��
h�<!���*´�:���Y|���f̀c�<)d?T`�|��! ` �9p�aZv�<!Q�0�bm8�n�Bp<�3��v�<i!+�	��5��)W��A��k�<Q�b����;P�L(�P-'�Wn�<��G��w~�QG٢O��]	���E�<�!./H/v�:�n�Lm9��F�<A�D��j�y���'@��2�h�<Y�ڑl�y��ͿM�U�EY^�<�&�V'N��@�W�7ʀ�F��[�<������@��R1h� ��'�s�<�1g	#N��	�1χ`{֥��y�<��JU���J3I���t�˔�r�<��D�3i�R�H�ǝ:��T'�E�<�f�]x��t!��F0��#��J�<1�!	�6�F�z%��%!�#��C�<Q��%M����͐!P�&�k�o�|�<I5)�Q�J���+�
�C��q�<y�-W�a������-]"�����p�<�㚜$#B�a��5AT�CgD�<y����m��x4F̰g�ŉ0��C�<!�#�:]�M�cc�n(�1�@�<y��U�1j.M��/ɉH�fP�W��W�<i���\<|�'�JlX��h�T�<!�Y��Y⃠�w�P� �w�<��R!sk4e82�H*�~hs"�Ks�<!S _r�����Ӑo>��1P&�c�<ᤀ�����F��O�ޅ���EG�<��
]��r���]�0��(��x�<�CĈ�(�z8SŊ�5��I��(�v�<9b��T��r���1)�̉r�<�֊�
SH"��W�7ל)%l�<	��(�.��#�?��4jv i�<Y�CNS_$ ��>��C���ybA�/'�yae��|٬xK�`�
�y2�N�*6�ip���mX<5��n�1�y򎓄zHy�Ë��(h�b� �y
� r��+.�09�WO�5AO�� a"Or����29Sb�SV��nm
r"Op�!�"�6|nt�C��g�TDJ"O�|�2��'kHp�v�²rA>`�G"O`D��\�	Ӭ$�V�Y*C�"Oލ���ã^D��
�*ͶHn���"OГ �<�e����p
��y"CЎG�6�'K)<�2�aUƆ�y2�S(Tza��m�8�mY"lP&�yOS����L�0)pdr�5�~��'�ᨳIQ�g�$I�U��"m\R���'�eb�0kv���T�C�j=2�0�'2>�#HA�l�8�yu�N`�&mC���O"~����spDm��L[�"��1¡�\�<iK�.���W�,8�qz� R��p=ٕ�$ ��Y�VL+q�q x�<ae\�Vk�A��醜B
I�6�Vz}�<�Ol0ؗ�)L��Uɡņ�.0d�"O� �c�ƪ`�xX
wk�2#.<Q��"O����@�I���%�X�YK�*�"O�I��hĨ0��1�4JZ�s2��{t"O4�������%�s)�=�p@a"O� �NL�?�,P��._�*$��'�1O*I�v�+��E0�n� z_0�Q�"O�a���0\�����\�'�u("OR�
1�� "�0m�#J��!"O��qu#
��x�b��L	��J"OH9;&�2�p,	�L[ )�$�U"Oh��G��EB�u���%4�Pmyc"O����"T!K�|��0lV�y��9�`"O�bg���9�PjPA�̩*�"O�г"�+j�v��e�Ie���7"O����bm��;���8�*"ORJl29�f̚Q	ߵ:�����"O������Cx���A�N�c���]���I,N �1���'l�$q��k"�C�Ie��y�H�b	A�k�8�C�I�5�T�Z�(�	�	 ���Rj�<َ�T>�;%���fu�!a)ۈ~c��+�>D���1%W+�:�u�W7hp�y)Q�7D�x��d��bX*�(�]��=� 5D�H�q��9:��)v`Wj�p�Z`3D��"Ď�b���JN����"n/D�D(%_�9Bj�B䣅8+����b":D�b OK�1���+Tg�bX� K�l3D�0�ҩ�����sj�4hnT`T�#D� �+�	���k���B�04���!D������}�(�T,R/>z�R�>D�L"���i�&�� ��$}̱@�I=D�J&���i !'��{;���Ă5D����D�	OX>��5��	6��tL3D���@��4�s`/�":b�KDg1D�T	2i�� �� #�a��/�	���.D��F#��($ԝ�RF\6��p`�0D��Ѥ?��x0d�x�g1D�X�����k`n�b�E֙j�v	�G�*D�h�&����)��D�!\�N�Q�(D�� �f����5��%�0�XfJ%D��q`�5d���$A����5�w�!D���޳k0��p�̀�O��u*��4D� ���ӧ~Tl��� )�ti�2D� ��T%P����w�!j�[&.D���A�H�`�Ȅ�SAR��P�@�i-D�db���(�\AX� �\�Fix��,D�� �=����=�r-���6h��pa"O,@9ccS�JP�IW���m�W"O�|��(؝*�~Qr��(*n4�"O�|3��ԅU������1-�LCA"OjT���	e6I��&E�u��"O�\{�g��$݂@vU� �@�ۗ"O0�# ڼ�\Л��&N��"O6@j��Ð3{�@ò�w�TpR"Oi
�ψSa��hA�
��^���"O�Lc�(���"U�j��@��%چ"O h�ELIOjD�s��en��9�"O����_+)�fH��I^'f=`P�"O2�C�*� (��M!P��7���"O�KϬh�PлQ���.Z��"O��Ɖ�+3�b%�DңF�tx��"O��Re�F9`p��A%��=��"OHqr�Y�ޢ 2O��$���
V"O� �aB�E�>�(���e�jp�2�''ў"~2Q�X�)4���DI���.��u蘶�y�)ЂIP����/�(ue��^#�y�C�ȝr6N	%����G�y��K2�I�HRsyV� ĭP�y��H�\��[���^�6�$g�7�y��(��� ���^6�1�2@��yjT�m���V{�eRϗ��yR)�9���K��9QtԌ(� �y�BՈV��qC�+xfT��!�ɜ�y��I��I�셵|- ,�.�yR����� e�� u��E�5K=�B�ɦ!�r `�ނ���*J�,k.C�	mU<��/�a�  "(J8��B�I�;��6i��0�6Q� !ʬ$��B�ɻM"l�"�I�X:�yU�R�CT`C�	<K���%�Ԑ)��d��l�6P\C�I� C�]hFN���H�����<C�I�ts�A��Ȑ�V�R�X&/�C��6B'nL���!�\"s-��&C��`Py�TEBh1l]���k�C��!7r�	R�/M V�%���B�I :����0�P�h�hr�By]�C�	�] �4�?�޵�u�S�~�6B��V"�B ひ}�	�� EB�.A���`�����x̌=f6B�
.�Ri���[�6���C��G�B�	!K
]`l]�k�8�ɕo��B�9�F=aef&�.�YA⇝��B�	:��[ІvN
��I�tC�.�F�0� ��9�:��"S�VC�	�`��Qz`A؜&�ؽ�B�8,�B�ɜ����eRYB�l��씝&��C�	�~VҌQ`�8��	�bQ�2\C�ɒ}��x0!��.�ꉱ'%ΕJ�C�Ip�=9B��w	����֧-�C�I$['���QW|�� ��S ��C�ɵS��,�'�L�ȅ0��+2�>C�	 vB�����>خ����ݻ8�C�I+��J1�2x��q��LP<n8FC�I�wNt����A7@(��L���B��?H�X���R�0A�&U�I&�C�I
O���;b� �>]��c�Sm̨C�,$E��c�n��W�᠁%E�f��B�	��<��$/��At�ۧ+�U�~B�ɯ�;�$:v�@Y���onB�I�Ru�J�`��:�n�Ix�B�)� ��t�j�D����ӮbJ"�"�"O �r�E	�Zl�3�&B:�����"O0�2g�c�Vt�T�S0W���
U"O�x��%ܢH�	� ]��yE"O��&�ԒQ�,��4�݈Y����W"O�8�g�K$I;�X�A��M�@y;�"OR�16��*6��$pu�S�2}J��d"O�+b�̢�Ld ����}�5"O�����	.2x�!a��4ֵ�"O~���OQ+�@a���_lB�Cp"O�2�����@�2NT�	�"O��H�������#A� %��D"O��0R�kxڍ!"[��&��!"O4�*�?G����+��`�"OV�ڑM�~�`ѡ�;4i$�8f"O
$��'@������ �LT(u�W"O���
&�B�#f�G���r�"O���ǭ_(���T�fi"�3V"O�1�k̥E �ґLA���2"O�y���.2 17��E�d́�"O�)@��K �l-Y�K��\t�4"O��KF�[�6�bY��ƀ?j�"O�P�'�L
����Ç�m^�t#B"Op9y����|c����"E�'Z����"O�I�J3� �C��BQ2iД"O���Y�>�*X�ۆ<<8�1� "O:��ݫ�a���'?LP��"O$�@�N�1)�.��%�Ŏx���u"O�X��9�sWT�O����"O��r��@F_z�i"̇^ݠR"O쥩�&L�R
�x!qŤ9��պ�"O�M�ѦG�M���j�4!����F"OP�eAܹ��a`��E87RtP`"O\`+B+��c�2�#�h[+i���5"O��Jg�~01��!֎��"O�m�0�ï.�n��A��$��"O�I���!*�8��A��:�ha	�"O���\z���z"�2D�����"O\��CE�K��x� �A��<�1"O��s�fʴp9L�`S�)M���B"O���`��_|����Yz����"Ot5o�8�e�j�e�B�8&"O�E���>�����%FPy�"O��I�΄���a��+F�6����"O��ؒ��/SS��c��C�u<��P�"O��c#L����ec7{L�`��"O�I{���)-Lt,ےB��rG�="ORyQѭ�,R��i�&�w<��a"O<��vH�9�$IX
����yB�Y�heT�0�,P�@K�&�yR��l��[D+C�*n�x������y�I�)#�j9���!�<��pjA��yr	�^�,�Hʛ��Q
q"�y����6)�'�<Z�)bW�+�y�Zo������A�1�Ʀҟ�y����|m�"�2o�,a�F	�y����+��(�#H �P af���yrAݪ���ȐA��R�!��_6�y�`}�X���t�r��լ	�y2�](����&�I�eo y����y��Q	;��qMZ:^�:��e�9�y��&�zp[1��6,C%a���y��44?zrQn��[�@�'ŷ�y2�Ϋ?�	�����W]T���m��y
� D���o�hj��SJJ1{m���"O�e���3Q 8!��ehp �"O�y��AHH�&L�H�*zM6it"OK�
a�B��V V�A�qK���	�y���e}fu�4\�j����bc:�yRC�-�4��W%�?b�z��I���yb�K/!>�{�O���k2��y�Mʐ��SSE3tE� �1���yBJǳM>�����l��}H���yR���,nX�ѓ�
<aS\Ѻ���+�yOA/���QƢ,n�ԋ��B_�<!�i�^v0�:5���K��0�2��w�<y��LEl䉲O]�V���KFv�<� 엧(X������匝���YM�<I�b��K��q�FM�2c����HJ�<�C ȅU�ʨ;��ܮ82�L�I�<��(c�>�9EB�RDH�AT��M�<� ��PȴC6j�	�����Q�<��fH�p���A�"*�:D�AN�<Q�y��#E5���AIU�<	d��q��#���Z\D��G�T�<���ɮv�.�R��0t7���R�<�$"�a��hT�E�e��YPg]K�<A���:de���1_�$��D�O�<!� �.}K(9� �+O�*�ۄ�M�<�f�	�T�p�Q�ä-��T3pɔ}�<ႮS�*�������e5�lr��v�<����5�`��\j��%zPTY�<�QH���&
پ|��x���	~�<�5��M"(�8Ej�-:B�H}�<�mM8N5�0V#[�W�X��q�^{�<q0���Z���V�S�Q�p����x�<�Ӆ��[T�h�#8+����i�<)��ӗyʶey��2/-JA���b�<��ʕ�)�9�3�i"�3`��]�<ɠ�� L�α�ҁ�$W�|Z!�D�a�$���p��yq4F��mK!���)�Hp��o��!P�/!�d�T��-��� ��~���L#!��QI�̺%�#(�nxi�i�ml!�ݖ| �q�H!G��*W�UZ!�$�4�d��e�X�q��䰥��4Hc!�d=��Sw&H-M*�)�B��=}!��e�UpR��6dI�ʴ��u!򄉉 ��`3���! 3X�Z�AW%'=!�DB�8��P��^�z�0�s�O!U'!�R3�(yf��2��Ia��%!��qq@�3��`�,��`
�V!��*^*y9&��W���H΂.^!�d$]p����6iŀ퐢P�i�!�d�#bUl����B�2��UᗈX�g�!�Ă2@^�v�
	c�$;��Ӳi�!�d�P_$�1I</�ĵ�WŒ�a��d�cĠ�Æ��IP�����.�y�iD6nk�� ��=V��2pN>�y�i��x=�C'^P ��0JM��y��H&Lil��I6&`�+�!�y�K�>_�t*�I$
dX`��V2�yr)�j;�*�C�%2��]_ʚC�i[�\�W��&dB�1����vC�ɰY�� GC/�(��ȓ+c�2B�ɤ&��r��6@O�T���w�<C�ɍ�x<᥃�3T0Rtŧ�%`V C�	�fΒl���˒+e"��@��t	�B�)� �i��-U��ƹ( ��&^f���"O�(e*�����gO�Y"��[�"OR���L 4��L��핐	��cf"O�E�Wȕ+|�<`�lH&��P"O&�#1H0f���.M�D,����"O�u���ïN;6�Ǽ7Dd�C�T�<��	�	&r̼8��o����U	X�<�B�Ja�̬B'h�a�p���z�<�%bV$~1T`��Rd���U�Hw�<	g�\"� �9�%Y�Y,��p�Mt�<!Ga�-�a8�+Q�㊍�@�I�<%��:ߐi�֯[B���x*	H�<Y�O��s�4xD*P0{��EkǦ	F�<�fHZ��B�R�!P7c��7ǁE�<��K���8G/εF�\��IGB�< N��e�p�`ɟ�`@�L�4N�@�<�"\*^^��!�*�r!1OOR�<�!ν
�ʅ臮ۤ�٨Sm�G�<��s$�-x��!�HdX�_�<yuѯ"���
�2?n���[\�<!��=�%@��2pR�j��Wt�<�v
�K�v庶����j�A਍p�<Q$ē�L	۵'�3g�m���F�<�ㄓR|d�AV���+7J����]�<��F/P����f��D���R�<!����`I�f�Wn�}y�&�M�<�	�?6��JW3�� ��G�<i��ح��X�v8�R��C�<�ZE�tX��L�mL��tքV�!�DR�S��sb��rGN��M��\�!�D�,`�:փ�."�iz�]4&@!�ݐBR�ţG�)@�N��LΩ&/!�$EV:��Eh\+��5)�KL)!�$ړ
�R�+g�I�!�H2�E!򄎉"�Rh2���z���Z�G/M�!��W��(�)a
�/w�He�ۃ
�!�d^�G5 �Y��fƚy9�DɕD�!�Ĕ$44X����y�p���D!�dEN��B��� ��	���>'c!�D�JJA*3$��p��0WD�vZ!�Dϣ)��a�,˂�<��ԍ��I!򤛜Hu�Ux���5��0�d���*,!�$Z(q5F�w`���� �$!��z/ix���+\.R��vIܽ9!��T8|st���.��-<y���9"�!��0�)���o��xg�<(�!�d��K$,I�w`ƾVgJ���3~!�� �
 ��j�!p�1Z���!�d��pV����.\[0Y��^!�D� c��C3�A�VN|�TA�>\8!�V �~��� J�:J
!C�.*j9!���Y�t���Ѻ.�^iK�.�!�
������H	n�P�sǅ\�!�䔰���g�	J�z��Gk�-�!�d��*X��E�=r�@2��)!���j���Ή? ^,Cr&\�
!��ߝ!>�9�f²;�5���b�!���n�I5#�0�\�XQ�Ɩt|!�D�d�n-���S��ڝ�Vc�(z!��*P�r9(C`L�
,��@����'$d�Z�EY�L?*8R�.I|@��P�'�y�����A091��K��G�<	�,�V-�]&��^$��]E�<i�/�'"lZ�ca��/R���c �B�<� Z�"M�V�v�3P��5t4�hXE"Ofy��(�/�Hx�dE2��� "OB����%�k�b �.�J�"O&Q��*@*]j�CӠ߷K��Д"O,�6.�?.<9:偒*�z�0f"O���p+ �%Є�c�!4�X��s"O���T"�#&�rAJ�6Z�x��"OY��̑{'��%O*�n��$"O�Ȼ�Q�mp�Ġ��4w���"O|]xp��b\�DZ�ɂhib}��"O�X���V+Ǆ����^vX.Љf"O��Hè;�p��JƊ5Zvqq�"O<�s))L�b4����@h"�"O����˂:Z�2�i�X�|d��"Obp�Pٸ`������j��#�"O�@9�Æ�;e��S�ƞ�g`�0�`"O��q�K�j�h-��G?L~� u"O�)��'�= \��(hԝ{�!�"Oȹ
��k���@���!#�;2"O�챰��5pm�(Cf「W�� 5"O6&��;��8���Z�-'D��`-D��y�ڎ'4���׍�N"`��/8D���P�� ��w�4����!D����0_��5�m���'�!D�,�WL�c��-qP��4QY?D�T��'.]Pu��-Ķ��t�t�<D����a9d�\*$�ȌŌ<D�����;��x'/Z���X��h8D�x#�ą�h���p��wv>�!a�4D�H��	�R�vA��̀�1M6u���0D���q.E XB�`'/�vy����.D��0pe��f���@&���l���&D��c�"�>(
d;g,"M.�4Ye�%D�`zD� ���� �[(�Uyv�(D���'����aŠ̢�\��.&D�d�A`Z�KQ��
�%�=>�Lu���%D���ӄ�8M,!��`�P�J�2h$D�$��KԞH�  w$Cg8V��R�6D��q%1&1��3`%�B�4�jQj3D� �Ī�פ��VZ�Cp��E�2D��5 �����0�T&J�I�//D��E8tg8� qOޛU�8Q ��+D��CF�7P��ȁp#��-��g*D�
��Y�`�8���d�������&D�`w��.jҦ=�B��Ho�8��"#D���EN&�Âc�&JټعAo D� �w��|E�	K �#ǺQ�A D�L��L	!�%��f"��P�!���R>��6�s�й�Q�@�!�$ҦBF����'ɚ������yR.P,7�T�Ȇ7��4h�e��y��7ׂXSt��'��r�
���y��kn��G��8ed(sP������0>��c�	Z��a�+���v!LG�<�m�K�qQ�l��.�6h��J@�<�a��x1�Q�oN�H	���)Y�<�q.�#`�%� �[�[e$ũ�� |�<i6Լw�x��PC�&	tIy���q�<�P�ô��u�˙+�΄�E�\G����X�ll!�	�#\�gT�U7���?��R*� �Q��*�$�`U$8�>=�ȓ�R�⡪�!]Va�Cl���~��'AV��9Ap��W+�xx�ȓ=Z�=87�	�7lL�4 N'[�>���S�? �ڇ�
.���[��\�L%�f"O��c_�Qk��s��G梉 4�~�D#2j�+��x�*Bm��"��O����O���O���qO��c�C��".pi�u)�>�>�Y"O4�#1���$R�ʓmܫi���"O�:����P8�i���=y�;�"O��Qu"ߙ��#ԡU�(j����"O��H�+W2�a2j�Q���B"O��F>Ѐ �1 �.<�N�t"OI:T�Ir$�pb�9�F�Xc"O�E�����=z>X�� [�7׾��'"O�5�Z)|�J�-�(���"ON��a�R�|��KКy~b�"OR�(�3iD����Nf�y�"O��� +9A)3��@�\ܝk�"O�Sf��_�00�i
�0@ hb�"O�O�-��gh�:_z1��"O
�S�Z�%�h���ӞF1�A�"OF��Ǝ�36q4Mk�͈��y��"O��Vjģغ}��.n�p��"O�0�@I�$]H��1p�F�l�B�"�"O\�Svl�e(�K���0R|l{B"O��@�̇�gc�i���̋�~��"O,�5A�J���#��۱�D�J]��G{��I�8{jڵ���)pMk���D�!��-��ux�H4\>����4�!�D\o::PҐ-�i��`�e�`!�Z�&�T�3N$H��9�nX5�!�V � ���j�Z��ruh�v�!�dW5>�1��c�i�ZAx���=�!�dްwXbѤe��s��á0lm�Y�'�А��U�H�!ucR?����+D�(j���
�RT(ҢD�dū�&D�X�C�8���4&�@�8��Q &D�P����(���eJN*dc"=�U�1D��pEަM�����J�� A�d-0D�,i��ՇgV�`�aC�Vf��(0D��f㝊~�,�#�E���U����<��,�+�źf��k�]�@��!\(� ʞ*t�����ԕ �F�ȓ-�6�H����[�QҳGZ�g9�H�ȓ1|I
�I˓1J
�×R<��ȓX@��d=��1��� �l�ȓ;���#6-Z.<̨C�I*{�2 ��C�ȣǬ�m�l5i�D�?I�zT�Im���0<	Ro^?:8�̂��ǅv!n��d	@J�<ASǓ�H}P��%ј��G�BE�<�����'7��۲O�$ �h�QE�I�<Q�N� \��hEg*";*��0.}�<1vB+��7F�2{�Э�Fɟ��y��ɩ3F��p� �n�8��Eӱ�y�L�=��q�5B
Dj��%���䓪hOq��ea2��+������ O���"O`�D�Ę/ph"'ǡ��1��"O���瘶]����U&G_��T�@"O�]y�(:P�L�
Ǯ�A���"O=�*УvB	�R�W(0���k�"O^��cY��=1v�֕4��02"O��0`K�-s��"B^�K�*�Y�"O�M�bW�Z�����$%�n|�G"Oj�²��Q"ݸw�A(
���"O(P{�b�=}r|Q���P0��PD"O̔�S�Ξsr�z�(��T��Iñ"O�Y���� �H(Y�i5W����E"O� b8{���J�z�F�%?i.��"O�$$�L�j�؅�N^ּ$_�,G{��	��| ���
u_4�ȗV6�!���gS���(Ӑj-�Y*�I�:|!�^��b̪�Kع5,�3�G�c!�D&�����B�t����MY!�dϫ;��D�2F[�g��-0�D'6Q!�M�x���8%�VE�G���!��^8;���x���j���'�!�d@x�ڱ�Q%^(�x�huQ�F!��A�m^�1��$� ��'Ѹk6!��q0@�9 ��<3��\Iaqx!�dN� ���u�M�(���+��oW!򄗐P�a�,.J<)�5ߊ0A!�]�/�� ��S	q��p�dL&�!�d�_tb=[`-Ʀm��#�D��G�!����e��.I�;G`���J�p�!�21�Tq����M��ba
>Q�!򄚯_�^�1� �Y�p�(P��3}!�d�J�bP�%gT�Rc8I��/ݏK^!�H�0�a!sĳB|�]�V��]Z!�O�U�БإLC=t�ĸ����w�!�/�(
���,b�8��� #�!��T�&L�Pώ�P|��t.˪�!�$�/����<T��H�+Ѡ+�!�dY��i[�aV/0�������!���F����$)�ۀ�2`R'=�!�d�:H�����T�U�(4aF��ɴ"O�3$Ɛ�UJٴ2��d��"OnU�QK�*��M�H�#;u���"O�`�f��'���P�@O�'_���"O*�	с�;�����/�2Bf�8e"O|�p���,:������A��8 F"O�)��G����i��	DR	�)*D�����-Y��YT���,�,��  (D���F�� En%YFc�5EjkT&D�Pڤ@�e:���&��#b���1D�|됩[#*�Tm��-�?C$���,D���§�=�p{���;�U�g*D��s!a�#��1�1�˖?d,��"�(D�3�������.ɣfc6ċ�D!D�T�PH'��%� m�.�  �3�2D���_y�Up"� F�Zf�<D�4�$�ŻK0 aҦ��5�#�,0D��R�R	w2���g�*M	�m{S	;D�8�F�
�2U��x0o���#�H=D�G�/q<X�S�dH ��h�F=D��
��]��`�!&�S�jj�I�"0D�`����OI+�'LN�������y������#��Ș@d�	8bS��y�)[�9�\u�uiD�aP��[��y2�mƔ�Y1�&����A�B� ��к�.$0�	Ѣ�P�'��Q� 0�����K6z
h���'B��Z�j�I�����ЗC%�qY��D7O���L�.`�����?�h��e"O��'ň[��3���0㲵�"O�Г"�\�_��Q��N�:u�l�7"O��! -G'e�2��F���Dl �aT"O�@鳧±\L2��Հڸ|��D��"O���_ l�$�)V��3	��}�'"O��CĭFT�v�����Q�ϔ�[!�"NY���B�^�l
���tq��'�'D�V>�&?eQ��@�o�X+6���P�d����W�<� �!�%	м���E��DW��0"O��X��E�~����ƅL��#2"O�0B 釷dg y� /	bc2tB"O��!��Y�zn֌P�)"O���@�=�P�3K�3llf�j�"O��q����$�ك��	k����'�ўL�I{��Si���w�A�/p���M0-x>$��'=������{��Њ�&$0�`�'zd�Cv�ߢE@����G5	k�'Q��"�υ��~a���R�B���'-��c��B��� Ԯ��K���a�'r�����M�S�fI�Ц�>�,�0�'�ySեB�n�Q0&�>/�����"�)�Ԋ^	��l��1t�"	�+���=�y�핱{�Q%V�s:������y�P�Q,AA�>���Tş�y�H]���J��73�.�@��_��yrǝ�A{�q��kJ9S�Ή�`��y2�Enզ�S4,�\���"�����ybe0Zn�	�E�K�%m������/�yb�]4>(J�8�ߗo�6��R��yBI4z���kӲf�����)B��y�Q(t�bX�F �_�"QqJ��y2�
����'k	)S�r�!�Ԓ�y���C�Q1�L��!%�Tb�$���1H^�A�c�=J��ѨƘh�p�ȓz����%ŵ>�R���B�4��%���	V����7ɏ 
8���š�:%~(��L+D�
����
�/dz�����X��C�ɧ.[����+� x�S�Bߘ2C�]�.��ŮT5��4�"m��3p2C䉯P�iD���ux��3�\B�I6Rٳ��=P��´I	<��B�	3fh-��c[#Gv}���
Z��ʓ�0?�%[�b��H��ߨ4����G��^�<�w��+�n�B�eI�1�(���[�<�åݯ(f��j�- 2�� ��Z�<�  ބ"۠�AP�Ϣ��`�X�<YD/���`�J,?ZX�`%�@Q�<ɃRp� �5��'4�B��q��x�<�-X�"�����F�=Z���k�ڟF{��)</2
����.�t�	a㍜-q����O�$&�O���Q�5n����&Q�A�"O�@(ж>td�i�@�{k^��"Or�ۢj�DG�*��?l����"O:H@E��+P�u��"ܽI�!�"O��Rԧ�-Z�, I��!)Š1�r�D<LO�]��M�<Qj��eW��hq��\�0D{ʟh��@i��6 ��mٲBP�Q|~uF{�'�0I0�&6��"7�<A�Ȝ��'�f�#�gĢ3J��
D�_11��
�'8xq��9��s�ü(
~QJ�'�� 톥n�����N*�'� ș�l�+I��mӒϑ�M9(!8�'�`�0�y�4����8W(�B�<q5�\;>EN�"���)Q��s��Ju�<Fn��a��� &w+� ��D�j������'��p�'I��,!�$[�v\��H�%�*p�����v\����"��"؅ȓ)⼉k.O�䃠��&\��ȓjJ]K�C�܍#� ������i��2#�Q�!n��X��Fʸ��<6\�3��P���С+�͇ȓR��D
ށ���#���vٖ',ў�|� 굓2&�� 9��H�NR:&�|͐�"OT4��lKw��8�M�<~Vt0�"O��:!��&K%�1�%I#yf�-�"O����� N����~Vn�:V"O��R�HGYb�y:���g_.8��|�)�B�Ū1�ȌD��S�b�"BzC�I�*�ִQ��\>B^<��	H%�VC��G�h@: �P J �ƥ.�B�mB9�s/�Z�y��F�D��B�I�#]��8�@%.��XK6H�:"C�44��p�7�����LE(_'�B�ɗsVg�I�%6t�)@�P$X�*��(�:9�s�7c���k5U�O�¬�'�ў�|�&ȋ�\¼�X���52"�A��v�<�6j�+��qDB�|� �Y��	i�<�v�֦r���gB.Z��Ѩc�<�fo�,��U!lȦ4I�	Q7�^�<�5U�'cj����,�|��f��r�<q�R-_^�p�!Ce���gZk�<1&^\�v�2w�e�
��̄]�<���;�np��cؚ$���B^U�<q�)��D�q�qۓe��x��a�g�<qS�Y�U�싃n�<ͮ�sfk�z�<�ł_*h�q �N�TR|�����m�<�b��x�`�3�\�z�R���"�h�<BW+GoD���$�R8(��ebNyB�)ʧ/�օ0�KX�K^����\+����v=����qV�*!v�N�%�8�Iry��6��"��)@�"@R��3C�I�q��ԡ�دv�����z�$C�	-8����GDX�M�DI2gĥ=��B�Im�J���+ލ?�2�br���lB�I~%�����/���Q�E0h�RB�I(YvH�!d>�ҝ�3�יHB�I�n4*�kQj!��"S��2:l��Ot�=�}�����_D�PKݻ��1���D�<��P0z��P�HJ�Y{��yt"L�<I"`P�}�����K�3vW��p��^H�<�oQ�L�B�)g�V�w�=�G�^�<Y�Eܖop����A�P�@�!��Vx��Dx �4�ġ�`&Z�v�6�YUGC���D �S�O�]�B1�� � RX�q�'�0��BL�ꍠ�)�:<�J���'ʎ�yq�%��c#�B�����'Lp ��a8Q#�rRZxy�'YJԚЬG�p-z��C�Ķp�`���'u��Aa H017"1�eĒd[pY��'wظ#5E�|�@}y�!�^J-x�'�\�����]lk`���\۪Y�
�'(���L+R�h�{���MRM�	�'��A��1wM� KG�J�B�T3	�'��-P�h�vsx}c�g&7����'�Z���F9^M�e�U��^x�C�'z,��@�8\ ��X�1V	����'^�e���%Ym�(*��7V��M�	�'z6��
�r��B@�GY���'Z¤h�%� L�����=3|���'�U�ҬI.��@k��ʰY��'g��� ;T�I +ʓw�Qr�'�N��CLA�ǀ�J����E��'-�z��-����/΀W�mk
�'C^<����99jY�OM�J�*��	�'�� x�jm̌��@㍔E^�E�	�'1`ɫ�gɟ�V��׈ 4
E.(���� ��#s�ͧ*���A���@�y)!"OT�˗B�9)��m�`��Z6-r�"O���#A)pXh�5-�KN����"O���a�-U�2}᳅�R��"�R�lG{��i��r�����hu8]���X�1!�Ƒ"��h�M��a����I%Y�!�d��x(���OP>��ks���i�!�����zVK�)3��A7e���!��"z\L����
,C���%+�;�!���5+6���g��.��P�dʚ#0�!򄁝P�����bW7@�歙�㚽H�'�ў�>U�T�Ӽz`
Qx��Y�5pUص�&D���C��<���L�-��̙)?D��P�ƶXTf�hg&�b��|+�j<D��� ��J��4�q�6��� �E/D�d���M�Ɂ�-"Q)L�â�*D�8K���kz$r�@��rT�i'D���`���@�g�����q�$�$'�S�'0:d�3�� �r�A�d��_����[wJ�q�^���x1/��w��ȓz����B�4<���(�e!�>���*"̘��\�27��@q'K+&b��ȓkt�	e͌F�H���5m����dj��f*.x��IHm�
z]�	%�L��Zy���*,?� ���LL�Y�e٢j��B�I�\���/ħf���!Ł��fC��*� C!˗H�pI{娀$j���O����¥F���' �R�����:�!���6C�Z���`C�
��@2���k�!�N���9B&e���@�옽a�!��!2B�@�`�F!^��8��"�'ў�>Ut�9x>z�beBIpo �"�,D��9���^	tE�&��w�$�"-+D��0r)ؤR��=�p�;HP`@:F*O* �b�ǰSH�yE
�0+>D�"O�UU,��W�HѱgnEu|m��"O����*O��z�P�3�X��"O
T*����m=��A���}#F�'��	�<�B�֣N���#��: ���'C�<�)H�?	q���"W��%��s��ܗ'��$�����Ό8!������>kC��gy��'�axr꒿'�z� �ז��Eʊ�y"ɜ�d� �P�+��R�@M��y�H�P��d̍�VW攣w�բ�y��ZiI*�����J7�A��g���>Y,O
���F!2c^�Ц�mܢi�!k�<9��� e��Y�*��@�%XvV�'��{�?O�B�lиA���hw�ҿD$��S�"O���ѭ�'��)���$Af"O�E��$��N�P0�S�� �TY�C"O앛eQ*P�(w�A T�(	q�"O����M��}?.���NR?0����O���f�0~��j��[�R�z�$/D��0�	�x ��qt�U�hV$��t� D��x��Ғ>Ƣai��ބe;p�0 �<���?A�I�D���0+>�Jw���� �ȓ`�g �=��"5/E�)��K+��1���	��y
��H�o֝�ȓU�ڵ:�I��
G"���4E����	Ο@$��G��'�B`d	=~�Ɉܴ:�����"O*��iD=!��e� ���=�B*0"O�8R�.\�z��)��-���'�ў"~����><��EV�ފ>��y�A"?�yə1�fU�!�8g�XT�����y
� �uI�M۔(S��W�%�x�p�"O���!���. KbꀚL�h(U��$�G��8Om%�޶�6���)\-~��8S�'��D޴_:�� �oߛQ�ʹ+U.,ў��?��y��Э"�*�C ?� l�����y�ՁV*����߼NY����Ȗ��y����qM�,�s��x�X�37���yR,��"�уgQ�EW8=���_��y¥�+�
Ī�Ũ���vi�?!����h�X��F%hѠ��4=d�<�f-�1��C�	'0��Xi4�N"m7����@Z+fH�C�	� ��x�P �K߮���V!jhC�I�"��H��	����MR�$�fC�Iئ#T�S�o��h�Q�ϿJ"DC�	�$���{��R� 2D^C�<n$|��%������f�`|C�I=nT�kT哢
֝��[D>�C�I#GxY�V �=a�`|a�%M%.B�4.bI�`./nAZ����E���'��Z5���'��L C()&�����>D��hU.J�\�"	S��Kwq|4��:D��sΔv��}��NޙM,�@�`;D�h��cא0M.����Z rA�<i�B�&ekD�:V�6�8@� 4N��y�.	H��U�S�����0wy$X��p� 9�GA��U���Q��n�v0�IQ�jy��L�L��d 3���#�م�4��W�&D���h
�nE0qJ;]�8��1D���6(�=R+<pA�֗"��9��-D�Њw��q>ū�1$�4�D-�Iȟ���@�S��.��g?���Ջ]�\5Z�s%�S�<���;{�DKW��J'�5�7�Kh<Á�*[�D��/��]�DȆ����'Taz҃<7T�LhЈ��ks6*�G��yңI��I[��ʹd�����G��ybM�}z %#����rP),߼�y�τ��=ぅ��|�	�&���'}��?�� ���в���;��BS�=D�������,*�@q& B����m;<O��ı<Y�'Z�$�cEA�v�ԉp���7Z�����-O�dɐ�??>թ�-�$Y�*}�""Of����ӓE�>l�sG��.� �@�"O��0��6nb`� ��s��

z�!�W&t����4ǌfTi��c��[���Ɵ��II���SR��	�4(�/vj�,A�oƏk�ޓO��=�}"��L�q?�t�Ō-$_r���iT}�<!_h,X��ɾ>�@�r���6���	f�Iyy��L� +���q,�2k�!-��B�/6D��࡞ab�������9&�7D��䫀4$�L�rЈ�$�z��4D�t��B�|/x<�+�s�,����?D����
\�
T���L7^� �QR.=D�İwG��w2���S�	5��`�A�>���Ox��>U���8Z�	��%�9Pl�,¥$;D��1jR6����튮h^��vg3D�,���-\Șș&"T(|u&I��/D�l��:k�
��ĠR~��TSqE3D�����ǟz��3�����$�+D� 3���5[�0�t�*d�rR�(D���u'�%���r��	R � �g&��"�Sܧ|�͋��̅j�~�(� ٴ���DB��Tl|i0	ȃ9��	3r`Z7MB�ɫR�¹)c֎/�*����k8�C�	�Qv�s��T�/�H��G ��C�)� n�p�ӿy��`z��۞s����"O��SQ
V���`��2l�>i�'"O�T[�ǂ��� ]=
�ū��$+�S�鑹X�P���A^{����/�	��OrY���K�� �^7T|11�"O�,�#@]��ʸa��P8�iD"OT�aD�)�&x*���EL�!�"Ol�a����H��!���K9�\��"O,H�l�'R�Y�萬	SĈ�"O!��O�l�by�&�#�J,��"O:h� �Q.Dj6��AK8&,Ĝ�"OQb�g�9���3��U#Ju9�"O��:qA2�ЃWA��*E"O&�aWn�6�p��~k8@�"OX�R��S�F���6dM�����"O�8 e<ud��C��0�"O��d�ߋd0�)����]� !q"O��B�۱g�*��oS�J����"O䕢��E=8��K��2���y�B0��D ��l�h��,�yR�A2!����*�9�f!+R�U��yBH�4�-�f���[���b�(�y�)�<�dl�̫"�d% �[,�y�]�l����/�Rq�$p7�Z��y"*,Q�h�1�еH��b�(���y��D�[ �0rCRjn䃁j��y�(O�<����)L!1d�2	�y�F�6��yVo�ul���p�]��y�h�����`+�7y�������y��+j@��A�����U���yB�J�o��C��M!�&%r�ɛ �y"K �]	>U�P΁fψ�"tc���y�h0e��|�eQ�l�t ��C��yb'
K�`b��f�D�w�D�y2,ԃoK�;���;[�֬ �oݼ�yR��z�Ѫ�A��T��LH�H��y2+b:��ZUC� O9����y��] �������0����y�I#m��< ����[�i�D���y���(���՘Y�	sUj#�y�K-dB�Q�7%B�fx���7�]��y-��RJ��k���<P�`Θ�y�ƎI� ���K[T��sOȢ�y�/��t��A�X�y�DQ(�y�P+�\ÔNU
�q�1A�1�y��,H�l��"��:� Y�$բ�ye"0�|tr��j�~EA��y2��E��3v�ڞb�fqbZ�y���T���'��[w>h!�$ʿ�y���t�r��UB�N�JPCPIT��y�`]�o�(�J"��G���uń �y�B6P��5Z�b�G�~M�TD��y��K2���d��C�����y�	6E�@������6����3�y���i��MZ?9�>uH����yأza��m�/P�1r����yR/ü#�|x��f�� e�u#A&3�y��\h
(tC����M�� ��y2�4��8hqo����Ȁ`.�y��C�v��Q� �
����*6�y����&iX�,�?U��I�G[5�y�,�0r���	e��I�
L)�mM��yRέ\�D�D�k�dq�q�O��yN�n��IFP8\_��"Qm��y
� ��I��@/c����� I�s�"O"�Z�`��u)�Q��D�<q�`�"OĘ���߀K��J1�͞p���b�"OJa�g�+TRXC%��\�y�"O�����G�䈉���*cd���"O�$AC��!�<�!u.{�FU ш6D�D������sҁ�� �T����3D�$B��$,.��PL�b����<D��Cu+�M�B�g]�'�D�F�9D��C��U�=��\�C�)m<��%�!D���O�q�
�}L$Y�'-D�`� "<��P�
Ʋ{Bڥ()D��s@g��C|,iԨ�0u-nQ�C�+D��8Ц�&p>r�!��9��Q��"5D����$�y��d�sִ��8��&D����&X�#p�P�� ��V<z�B5h&D��Av����#4���P:"}!�!D�(0�LA�Vs��N..���%J?D�h�Ł?
D�A���͵k��(���=D��A'і
�l�!�jǼY�Q��/=D��QB)�&�T��v#�-�Yj��0D����i���q�Ϛ3,ƹ���!D�8�q)�%=�Z)�"$�%ׄ0�>D��!�lZ�u@���N
�J��c=D�HۇJ�xM: ���2U��1e�5D���"D'�Lp�3�?T�ĥa �3D�8��A�;�Xh��]�o��@a1f1D��y1��8- ZMPF��Q��\�2h<D� 2QB�c.$1��W��x;VM:D��&��6o��`V���n)X��6�6D��C~�LD��z���'�5D��V+Ԑ�����P�'��|��`1D�P���0pƕSv�к"��`� �-D����6/��T�-N�Pl�a�J1D��2��=�p�ӷ�L $վ9F�:D���j��xK��q�*94`��e�6D��-Yi�0cI�-/�R�+gN�qN!���+�lx���A�nؒ%&��9A!�$�2/��)�M��w�M��D+S!�dܜ{��[LV��0Ah�T�>3!�	V�&V��Pq|����V&k��ȓFq��x&-�#B3��F+$F�xP�ȓC�� xFE��������w�B��ȓwH´��o�;�|+ K�}Z�T��,�EAs!�X��5��>�d���.�d�:B�W6@d�	+��M3zC�)�ȓsx�#B��W�,�2�gR1\TɄȓ_7�p���D�'I�M���R�Az��ȓYh��@��=v��pz'"L,_�l��2��PO ��!Э�*�t��$��Z����Ab]�n��ȓ ��A%��.��-��nٹ��ȓx��X��<\2 ��G*$mJ��ȓL�v�se`�G�F)E��$88�$�ȓK��K�I_�<� �..B��ȓCn�A�M�(v�f�S$vRx��ȓ����]�^�� GM�~��ȓ��8P��3Cͪ���[Nh��d�i �DJ�1�B��@R�dd��ȓz�@u$�,VqX�`�_s��ȓT$l	�4�H�!r@�;�C�&*~���c=�剢�H8��ᥣӬI0�؄ȓU�>X�@��>��2K�'z݅�jn���hٺZ���#�Θ!I��5��S�? P�yw��ʒ(:�L~:q�"O�₁�+=�@��Gm��|ı�`"O^��C"קQa$�k��*t\a�""Oȉ)Fc^'y�ސ� ,O[�	A"O�j�n�&#p8�DU'a=i�"OȑxS��<y�������T(�hn2D��gņ�(Հ�R�m�8V�hy�<D���t�������	ԋ7���X�E4D��ӆEH0k��fC�:Q��M�@�2D�܈��� ��C�[����%D��p4	_���z0@�#1[LUc�&D�����-Z����0ECE�(D��bD�^�P��m&+�<AE9D�(�gI�Fzh�EIS�<^xYB�5D��aBII�-�`��A=Pzc ?D���D)V\�Z���!.���;D����'�0y��g��	q�J�07f8D�t�$��&�\�`��)
�!��5D��	��C)r��P�w��*�x\��@5D�$2��OR\��зP%����4D�T�E!Yh�8��^�x�GK2D��Qs�N�R�Y ��xXy8�.D���m����"��Y|��:A*�X�<���( �����%h�=:s��i�<��"��Tl��3JWRZBm���Gq�<!���5=g��srJ�c�UI�b�u�<�"���&V��eE_%c�fl�1-�n�<y⃘�&�	!!F$�:�3Ei�<B�Ld*�X���I�8���!i�<����X����A�?Gn���e[�<AĬ(>�M�b�#G~MZ�g�^�<qu�Y;OA��AN�p�Z9���AF�<�2U5Z��PI�
I@�� ���<QT��_(�3�+v����{�<i�A�u��%jaII�.���kb\s�<!1��"�uѮݤmd(ۦ�f�<� (F�1�ʙ�D��H�*d�a.�y�<i�B�sM���� N�jx>p٥J�P�<т�'5��M{�l[Z�]�f��N�<Q�ño��@3EC�P������U�<�q��=��E��%���ʍ\�<)׬��S�@�	�-B#���Y}�<��oK��\Z'��e~"� �c�<��Hםg���椁�O肕gVW�<1!����T�&o�_�\B�aMP�<Y�Ȗ�c�0Q�U�*�%��H�<Y$Ր��${a-A��L����C�<C���[M:�S� +@�:�*RbD�<�2��2H~�ӣ��Q�,J2�C�<��*I>8�q�'��b�h��s~�<��jl6�1" ]G�r4���_�<�W�<oμ�w�ƖaM,	��ˀD�<�3h�+����b��F@^�Xv�@�<�%��#c��hAD��S�(� D��D�<�&^�qDj:4�]WX�@� �~�<��dT`B�z�@���}@�y�<�!��{�ezp��{\0�8q�r�<����7n�i8��J�m 	w�<��ܴњ�YpHU�M�J��`q�<Yr�N�V��
sˎ��qIR^o�<q�%͛_�$��5���k�<��rk����'�bo��s4-GA�<a�G.4�"f�	�=+�+ {�<9U#�\�½	GҚvjtے��s�<� ��3ᓹ@j�iP ��f��MHb"O�6������E
|�Q��*6D�H���ֻ�>�Y��,#��g�<���E	���IK �*�Z[�<�V
�kH��e�`�V��*GW�<�5�L>�lq-^SY��(�T�<���MOfz$�q"
�@�r���[g�<���aDJ9qc�تz�<Q���f�<���+W�~�
/�)*9b�0c�Ld�<�K4�؇fM:	u@��5�TX쓧hO�O���ԥF�v����`���R
�'����+�'�V=1� �@� 
�'�~������cu,��oRP�	�'�2⅑,�x�*�;NK��t�/�M[���s�*D$DT< �JHAG*"J����"O�:��;�vȂ�B��D5�y�E˞��A3b�%�j�rO��yb�\�A4��j3��yx�������yr��LF�e{�m��vQ|��ǝ��MK��D�k�'��M�p��߰ !��G��*)ك"O��%�d��Jg�����"O���to��)~L�3@<w� 9�"OZ a1G��#�����hR��Q��y���e�l�'X�1b�rw�\+�<���!,�x�*T%0T�-:��:{�!�=YD% ��O\m�@'�<Z!�Y
l�4Q����e� ����!@W!�F)BVM��A��t	��{U�V�`p��p��=yC����d����8R���Alf���I>��/'(�P����T!%�qːCL�'����i45���B�	�� WkB�(�pE{ʟ4�u-��7V�I`�HZ��^=��&o�8�$���)�g~2���)�v��1`η9^���t�V$�ēyX�<�~�Vd�v��;���R�oAKy�'���D�j�.�����,����@D7�?��4�yRU��C�����H82nT�^�0�a%�n�ȹ"�6O�"<!6j�:d���@��<��+�e�������<�J� G}r�;
�.��䎒<�*�P�V��hO6c� ����!'��Js��� �&j� ,Q�"O�|��D�%�Jh�A@GZ74����,'��>�p�9iވѶ)߃�X�p�@%D��R��وT����ĊO<�bB0�OĒOh��&D���2!'ǔb�jmP�'hqO*%�ӄC�N��TƔ�E��h ���[�OH�xG��Q�~�R�ٙAv�q��'�0���*�F&�L`e.�<:z�Z�{��)�iב`�̙�� �$�6���J6Oax2�ɭHέ�O /�����MVPC䉅E�i:R�I��mbNMo�.C䉴>�5pE�_Y `Q��,�4��B�ɂ;~�@rFI�r<�����G,H��B�I�6@|pA��\t��+���e/\"?���ے��s���;s�hT��LD��d{�H�>E���E  ��s�%P�E��)+�	��y�Γuc�X���R(���ڑ�E��yB��2*�h�H�-�P�ao
��?��'q�Ip��ݔJX��p	�"LL��'���×��hI�����ppLK�'��	�j����Ac&�D" }��'�2I���F	|<y*���J��$�}B�irayB�"�tM�u+A�"%<�e�3�y�.˾%�24E��ql������y���*q"qo�*> ΔzU냨��D�:�?9�'��I�u�q����+j��XsRhh��yA�"O� ��ے�L�l�^�I�'ۼpX���"Ov�[&��[�`��Vō�U)�q� "O��c��K'�����䙌T���:u"O�l��kF��a `�J&H~�2�"O��%��p��E쏰VK �"O���� �N�I�zeh��B"O�!!rO8'��arW��MN�ܡ�"Ot�9�̜�E����##m&q�"OV��∌�l�X�C"#2T�B��'q����!��tv����A�A���ȓ' ��%�4`�L��]�;"��ȓY0l���+�<���dg;��ȓy{�����_X��"�͸]VQ%�HG|�_�����J���WmՉ)���*`C�.N�|ĳw�ѕD@hE)eʞ�7c��G{J|�@�T��A�@F�'P&���T&Nb����'�h����ջA�,��Gl|t�۴�?�����iڼL�&*#Pa(ƪ�1w:0� �'tdVGM�6�$1�/O�"�R]	�'r%�#��)��=�G�F�M��`@�'7�P To������	S$h���Q'!D��h�̈́�-PD���S�6>
IA�B>D�B��V�D����mN�g��d�=D�@X��
 ft Iw��eg�A"=D��ŗ:[yru�!ȉ� ����f@<D��i�Պ�08J��C�CP�0ې$:D���J����jS%�;j[�X��l��=E�ܴ^2P��/��r��T ��X�f��ȓ���b���:H$f�Z��k�����Em�����.A���æ��ix�Ez��~�F,ӆ+p��(�8o�ژ�F��O�<����+��j��G�-��H�%�N��hO1��P�t�˅�"���J����6"OH�@��P8@���[2v��A3��i����|bO?7��v��}�G�Gz�
0��5z !򄋲;��!��_vtK�-�*�!�$�T�`���db��cM�%W�az2���7O��U�ΐ42@j%Ӈ��>�!�DD�>���AJ1@��*1��~�!���,��$K4bȘOʭ�& [+!��G�x���#�׽Oe"|�d%0}�F��QD��M#��þ|�dp�T���~�*�`�D�<I�OM3'�4ɒ�8/���Ja�e�<aF��.�,X�@���R�*�/Av�<A$b8>>���¯Q#u�j�%Qq�'��xb�W4O��YtL�&#��t@�ƞ�yr��
yuƸ0t�e�����~"4O ��D�	���x�@.����Ҧx���L�D�}�O���� ��,ò��7]��qG�4}��2>Ov%Y�I�#(�����M>!����&?)���3f��r��W��M)��ұa��0G{ʟ�����	A��5�%	֐Y���1OҢ=E����N��(;�-	�R���@�/���y�ݶgv\�3�.II�4,�Vj�5�M;�O����Xj#dh)sQ��D���Iw��/}ʟ��*�'k�dѴ&��Q����gX��� �3D�����6U���w��AF�;�	a���'<k,j�)L�]��� �	'���8L��&,ii���+�j�����;`�Js�l�b?i��+���c�
��v�k�2D�	��ʶ7bJ�j�cM7A�"�)�+2D��c��I�_��l�IL~4T�CG2}��|*sG����Fb�4d����3b^4".�-�3%/D�z H�"0~�� �ܤ�,�	�1�I��p=� �H  �͸}@�c9LZ�X�5Obm�	q�I��Gl.[fB��x�֒OL��ē1��A
��]�B ��w���A�ax�a�'��=Q�[%M��$0#灸CV��X�'�Fm DÏ�^Z�X2��-=Fx��'J�ГT�ҥ>wԱ#ʒ+k�_G�<� ��O��Ă2'�Vcӆ�{�<��b�45��Y���H���x���t�<Q� =7N�s��׵-��IJm�<��C͢dp�3�.A^x��!L�_�<q���UO*H٤�ά��,�^�<��lA+c������"jH�};6�_Y�<� �W#�b��0#�.s�,��T�<�C�ǐ-l©��
Y���L�Fa�O�<q��O.<@\�䤓�,}!c��L�<��A�` ȣ`�XI^�4i�Eo�<�rK�<��p"�',���$�h�<A�/�5�Ф6��iTJ�<���08x��f-͉a���J�MK�<�ь	
R�p"Do� zn-���ON�<y�TQHi�B�݆1�y��OT�<q�#
���9a��-�B��W��z�<�&V��,�`���~�"\)��o�<�W���u/ѓ���@"��n�<a iT� ԫM�վ�� LLE�<�U���>	 e\�m�@T5�m�<���҂�p4ᱭI5���)S$Va�<ّ�Β<<� #f�6�x�a��s�<��&vI�T���2:��i���Bf�<�W��_l�p@�E�k�~��d�<GHH�К�aW��o��Q'�TZ�<2�V-0",iBM����8��cYV�<)�@^�p�� ���B��2@�U�<�L��ժrK�<�iZ�R�<q��3s����2lɁh2�q��i�<�Q{���'�ܻs�x���O�i�<�@M�@��,
��^5)E����d�<�-�}��- ��;_�&����\�<���W�n�Sr/��J��!���C�<qg莲< 1�H7iY���bf�E�<ɶ����P�s��&�\	�&�h�<���W��=k�d�7m~тRf�<A��
�u����� �~"�\j����S4�< G��C��<ɲ(��Z���H�I�(e,QY"d'D����	X)N�Y#�����u�G#D� ��rz];D�G�1r�1�tN?D�t�1�X�bd�y�C9�}�r+?D�,��2���"��X�uI�1D��8U�C%Z�X<�A�h�n�r�,D����Ɲ��XR�MH�kF�1ئN(D��X� E�����Pn�(`�yy��%D���.�N���8���"8���E"D�ȱ�O��:s�`���ëI�I�' D��b�'#���U&	��}h��?D�����N~<��i�i3�q�#o>D� �O&-����@�;S�v��#+D�(8��̒g�J��L@�L�^a��&D�1�[3k⬓�#��Ku!�!D����s]�%@��)h�+D��Ҥ/��dP�9C%�6� x1p�5D�,�Άg�j,B�ě�Y9lA��5D�LibD�
�}XeJ�9u�ؐ8ө1D�)�F��(��8UD��
�g*D��!���0M��Lq�R7+���V�+��7*����{��� 0�S��@$���W5<���"OιPK��U��
1�R4�\��4��"l��Vc(�3�V�_3d�1�H	e�l�r�͛�;�~�BY�xݸ�;(h�y �b�H����I�����V�ē�5H��%ғq��SO�2�p%�����D{" �Fb��3��C7[L���#�d����f�X�a>���0�C�y~�٩�
�d"�	�]_��z��0��SoL�C���o�^61 Y#w����h�0y������%A�����;PtБ
j�Bl�w��,[ªa�ȓ���4���b�V���.�	b1�M L��f��>_Ċ��ڣ���4�l���u,���!λ=d��Q��bcHb���c�zy��O+���e)�6��LCp�϶8�ZQˣ�߅Eu��K"�P���d���4<���ٺ&De��N4<�VEӋ}�)O�(a��3��cј��_��O4�낡S^[�t��DB�, �0�A�ӿ��5��+efYS��W@��d�ҌX
o���F70Bn�8�Mͦ�p=As����AI�J��z��� �44��pѿ|� W�;LE-M��� gㄽ{S�R�k@��\i �i�nX�U�X�U��b	��Xk$����<D����0�"A�BĎ,,\*)Kc'U*u8�3��Ҧ*L�����&+O���r�S02{H�݀F]���w@D0?����bf\���4V�8S3��(ނ��V�Mn[|e�r���4��r�lS�H঵iRd`Z&#2KZ-�q�Ը��$%F&��+�B#�1f���&ψ��\Fx�C�H^r�J���9g�Z%��9ĝ����aN�PWF��'#D�2u
�^�X�ڄ��pn�,�"�Q�^0�̕*��	
]�D�x��?Uy�E�g?b���D#�� �pAX�1VCǾ{D�b��0
YY���c7r��gd�������^�us�D���K3��
��7~��)�V��<�JЗ���N~�<�UK��H4����*\YQ��L"[�|��4�ݜ8�
1���c!���k�	K3��ɓ�/Nyi�B�#Y�|���֦ T�S�I�0S�Tr��r�bqzQ�1=�џD�)��v�rm���*���2���<=���l�?5�z )�,b�F䓃 �o��3�A+ ���Zv�<<�=�f�O\���Ε�m�A0@\ˢ�1�,����.U��R�Y f�1FH�"��	N�FI��&E+�j	�Q���_�,2DJe@���)�28Z���N@�F�
u�aFD(�v9��T]� *d
PgD�#�ǅ�u&ܣ��љ)�Q7�d���h�N�yQ�,"�  ��`7�	� x��E�5^�=j.�wa��!�C9a���NŞ"��,�ҭ��8b���$��p�w0���8�{b��p��8\^buO�.��m��rM�#?TH0���)���ɂЪ	��E!W�B���ye�$��\�Ojʸ���@�U�`�;S��.����M:
�
"?�4�^iN�TYV�H<sW����̐�{�����!�2Ҋ�K��˝y����Ȉ+I�c�mI�sP���w��(~������]1ؘ�G�J���<`����o�\��d�!%4܋����	�"<����T�L� ��B=Iz���#CD�j�2���2&��u�Fc�ߦ����S�%_Z�y��>�M�Rǎ�s�m���ʉ7�G�ی)v��x�(ݚ8��T+�������KW�ص�Ci��4 �8��@�.�M{�
�;6{"uɖ� 6 ��U����;CMɋ]C��RhΆԤ�����Ւ���_*��t�1��^T>�r���YJ���	Ѩ%�UU���Uo1P#��(���âl0�7-o�L�b���JMX��ƿ_R�#?(\��o�R�>�V������+���)&݅���v��R̜rQ�c0�Y��)��k�8�7�>�`���}�0	�Y.<jq)��.DBd�dFm������B"�̹��$E4MIj�-޿Xr4,R1�\(*NXX���h���õ�B�	�)�P�l��1� �H
d���ܳ&���'���@;aVt;�ݿg�逍�McW,�p@1R$S0\� ��ٝt�\܊P
�%F0��a��Q��į�r@9rD�0B�pq �q�D����0������$�
��Eގ<�| �1L2l���2��]����0����	ȭ'���u���?�l$��l3�8 IT�Կ���"��K�h5+��ÐA�T͓akA-�ı�I���.!��U����B��
N�p�D�0�����(�s���\�����I��P�ɑ����c�4����A�тs��+��]����)C��>p���뛲��q�6�,Loj�s� �k��	�q�5j�8�d�G�u��'֮���K����%@0ɕ�?/lU2␠ �:�ᕡ��R��s��'F+!Z�S�[�]9�IU�=,fIr\�1H7鎭Ӣ�DJ\�3�M�s�@���H��Cb����E٠+���'n�Mybkg���#��N���8O�����Y�+A�/��ǈ7>�T%��ă���������uv�H�slU-G&i�X�&�+�'�7=�N��CӼ3&-� ~��<3�@ַNz��W'Ǧa	��^ec�����<�0L����Op���GO�eߤ$�en��w[ ��T-H�`dU�_�(h	g����T���
ǄQ��@�5�Ôt\��
�-I�j|HŪHY��/�4萙$�!C�b�i ����?��ϚO��*�J��b�\�woŷ	���+��@�n�QPM�}�D\���P.�E��W1(uv�EɅx��jqN�{�j=��g�tU�hЗ�,䠓O�l���Q��X1c#`�n\)BE�jXx�X��U�� Ǌ3��gƵ-�j a���l�p�CJ�*|L�+t����CEjǆ�x��Y&*DH��2i�0;X�����H	v��x�%��pm�<V�Di��Ӱf�F �`�(�s5),�:5�06�B�	�N�=T�Ny��,R0g�B0s�M��c�.�ݼh�h1֍��F�~�*���1kW�">���/��	�C�0��eO�aҀ��G�k�8X�2���ue��Z�N����m��SDΓ^�ܑ)U��
�be�P��"7�ڈ��Jݙ�?��)��X:lQA��`����y}�A+}�n8��y��F*E;�	�9-�n��@i^:6�:X��E�!>ӄ8q`� aP���L�&٬#{�AVb �@�ўl��ʓ�@N,�����#*�"D���#BH"��1��!
:��D؄�.R$��	�$-�Ё⟖e��j]*2�A��5]"4=h4�N
^N�$����UI���$ߜ� ��՜Nx����6{@��!� �t�F���H�edD�4���iU�Ls�Ĳ!�4�~�5hv��voF�9h�r��ϰ>�D�!�J���J"V¬h�bD7Ay����,~�����4d&^XK$GX.1���H� ���`w���+O� ���tz�����Y*J��鉗=�v���mD�;S�@8���(�]��-��Y�m�$Ov�r���t�1$���vH��	96��%e�.�<ɑ���!G�7�������[$>^�[D�Z�ua�b���KU�i��O��2���x��x��IΘMҼjd66k���I(mn�$p'�U.���� ��=v���2	A�x�~��fO�}F���:/�\���o�䁊0�E=q����� ~�d����w�0%h��߮w:����#n�л���=Z�:1@�$�/v8牣o� ���hRC����V�����
Ԍ��c/�ĳԊ�hL�PΜ/F�,yvB�=I�셙�đ/���BT��Q���� ���S�� ��5(�X�Ί1_��q�qe]�?Yp#҉�(�U+Y�����F�=$�x��ܽ<ьq���GE�@H�+��(0���#�6?�J$υW�ʅ��'O���5,ǽ7��QHTo��>K@ш�_�|�sc�Or�9B�G�#�v�:���E�>�A֟���D�\��5P	F����lR�>ZB���'����l�;PVАe��N� �d+�:�t�ʲ��'cLv����1I���K��(.��h*�D�;K�4$��;�z���+�`Kz���(��.;�#Ek��bVJE����&00�Ox�dV�QI׊W�cƮ�ӁLchPx���{�����͇N���*v�R o|���	����X�4螭` ,�޴1�:��#!���u�@%���T���i������
�`*J��q�� ���_0!������q �O���k�+a*H��1?���� �Q�̩k�WTv����
S�����9 ��805Ň)��O���R�/	�ؠS���	°�8���}�$����=��؀̛�2����'h,��ȣNLͮ�@Siκz����E���4�0e�dMR�{]l� �j	]�<��Z$T��b��?�>��f��{ܥ2ġ�&J½�c!�o� 1���*B��I<L����@�sΉ��^��{!AE�/F���R,�_����j�k��l�"��3,[���������� ����B�h����@�R��V�t��J�Q>�@�"@���"~�M��y�k֡[�6���'[�xɄ�y�0+W�^�&�1�)�&X�l��Y'o��O�p�;+Fh!cQ���/x���vK�c!��������-m-�D#`����OY;���BΛ3_������	c�qc��9����I�c=� fH5"��=�S(��"��	d����r����3i��(�C����p9���2eͬ9�� �0p
 ��E\?WGX��a��A��4�iY���P%d՜H�AS�i2b��7M���u׊�%�9ʔ'��ʧb��L�v �	����	$"�
}$���$�����B3K{,h�
ǃAh�2d�G�2 /{��c��D�!�.p�gՁ'u����iʹ��e�� K��n�<E��4+\Z%�q� 
��UIq�Cl2��b��O���h��x�IDfR�.VJ9�A��|��FPO��+!����GL��dB�M��	6���'ܐ,axrE<w�t� �%��x`4��*p&��+� Ζ����iɆG�N�:�B[=t�\��h�Z��{��:}
9���ےP�zUY�i��0 , !A�'���2`�-lt�b�6V|`K2���F����%"�A����`�[f��@�'��5�$NV��XBc� ~u�M<�f����s�JV����B"��Da��qpD�vacp��7;j���&�i�5OM&7�!��Aݤ��W/AB"Ĺ�ό-	�	-�:�0D���~��𺠊`��vE}�T�ߘXN睅AF�a��:lp��7B�q�.C�ɑC�V}Y$���b|hf�n7,8��Gdb���jG�e&�&#�:�Z]�f��p\�=��& V���)
3Y&VL�#oay�B̦LV��*��j@�RVcN�F;�xj�����.$^��"ԭE3��u�{�v�Z��'��9�J�6}6\��$�g,PM>�椅d<$U)J��]y��ÇkGD�!��CV��=�d�E�`6�0��Çe <�@L��y�dFv�92#N�2A�Q@��Nh�XW��2��(sPā��H��d��t�=�O��Б3��	Zq@SJi�ʵN���ؽ!�OTH*�%�$�2a�,(ބ����X!��l�1/�/@pĊ�mH:_	�	QB�̤�.�T�>�Ĕ�H�R�V�X<i��!%�7d� rC5�b�MR�f�ٚY�#�1UB�]����gzщ� �3WΜ��%��8�TH�@�J�1c�칟���Ƃ���Xr��>��f���"背'�6!1뗉kP��'Mn}r*�-߰X��L�W_i��$֧&�h�!�
��?1ï�,�M;׍ $����P���?)`@�5q�ji	����/p���
�<d�L!���'b���Rg��/�&�k��N�pKqz&��s��	��u'�\�@���Ӛw�
�h�'L�\���ꉝ9�$3U������bUH���vIXi��{b��EԞ]��55ߐh1@j�6�,<ӣM�8�~X[�-I���)��ñ>܌u�#膷1ל| ��3�4�C�Y�?v �)BU�-�X���֬+�Z��P� gT#=)�

u:x�W�	�F����px��k0h�NZ�"ʖF5�qQ'��:��\yA�D9%�b=Ad�ww����NL@�s�
v�n��'zŬɡ!�'��9�h�$Vh`��'M"9*�,�O�����Oش#1&,�1$S�5��dj��y;�GR�lY�-R���=g��To<|&���eؠ�,��ӆ_(M� �S�'H��yb��%8���+�(��H���J6~��t�Cȟ>!��m�b�	�)|�h��)Φ>����͟(��\�B����ygn�5@�jܙ"�E�$�<�6��)�HƟ,)BP!�����Fyr۴s��sF	+j���o�J?�+6gɸ7`���v-��.�X��_�g{��+�&��n���"���O8�+v'94nЉ�� J-��J�u�q2��/1��Ay e)�P�|�EOһp�Q
S B.5��uA�cJ�L��{i.R�]�'���R2����N9��պ�E��}6RRi��K�dI�¿ ���9E�h�b�[�7�.ՊS�� O�ollE����E�H�hA�	PM�VfקYyعB����w�<�@g���6 ��//r�Ј�}�13�R�f�R͢�g� 
�~(�P����h�g�V�e��i���\#��V��f�C�O��H��IPk5r?pM�Ǎ�a�����Z3-�y� �����ɜa�@!��.DF����ˏM��YVkU�?m�5����o��.3�LV���џsg�{���X3���T�0^�Q�F�=u_���#�K�P�E�qc�s��a�Ũ�'�#R� H��ȕzZ�8RC�͒	T��zD�)ɚD���/�Gh��A�ʼX�j\�`��+���[�"Q��|�����.��0�>'/�0�-G�Km��RPm���B��b���Fد��'���7IQ������B/�`d�=y1��g107�}��ajM,b!؂�����%�"C��B3f���)�Kr]Rb��P+1j����\K��	��Y����jT���Eq�8����:��%�M�d��(J�T ��O+P2f8S��	�(S������=�]�7�� 9T�:�_!�R��j�'~�0��H{$ /�P�'A�zw�T����O ��MA�?�g�̵K*�� �G̷C:hCa��:7��1A ���`s���7`�S*_S����QeM�7A�W��+ ���(����'#�Sg�M)l>�)BlV1�ҍ�)r�]�d��
A0�"O c�D�ZhƜ�B��;W���G��7N~4���̨/ֺ�ԧ���
4>��Я߬�8i$&�"�!��ѕ,^��I"�ͩd�a'e�d�d�8lH)3u����0=aU���!?�Yb�AʪU�DaчÃlx�d٧��Vԛf�NechH$AÆ�P�	�y�`۾K��M���B�f�RD��y�A�Q��uR�ϒ?�ްZ�B[-�y�G�)J�UH����~��lJafָ�yb�O� �8��}$n`�i��y2EK�2��o+m�#���yR��N_~��I�d4�U������y��
:���+fE[�KZUI��F*�y�M���܂d抃�~�zנϯ�y�kՌQ��XQN�c�8ӆ-Y��y�$��%��1��8(�*�SӉ�y��X:[Ĥ���t�����̑�y"Y��ЫrH�u���� �yB�@�!�����A��0��z�L,�y2��-R�k�@E- >!�F^.�yb��b�0�s��$/�6�S�O��y�/�=A�F;��P�'L���nڝ�y(��D�T��eXM�2Q��y�HS�q,�Q�T���b��W�y"�Z`TU D��o���
2�L$�yr�ܙb'2�I��>XthQ�M1�y"遰��k�B��]�N0�"O^��y2�]�x�� 3���H_����~�C�ɟ/�&ppg"�;Ss��G�)|V"C��7MX�h��Ut�����4|�C��!����虿g��l��L��Bk-D�|Р�WX���C�R$^��vA(D��Je$�='`�i�S(��g�p�{��4D�<�k_5��ѳC3{ X���A5D�@hǀV^��#G:�|16�&D�Dy �_-�Ke
�Q&y� �)D� )�'�,x�DB���
)*ܔ;u�0D�8�t��'{p�q�G�X���S�-D�����ʅ!?2$j�Ʒ1��|[��,D�$��i�<�|����/@a@�B+D�zī#|"q�Ƌ�.�H9�$�/D�8gnp# ��A,@��@p(*D�pCUhVUxsZ�_��d��a5D����叢=v82�Zm+�J�!.D�l�"AN/x$t<"�ٌn ��p�(D����'T��Y���Ԗ�X�.*D����)��<�x�1Ɓm���2�(D� �A��'�(ԩ�c�
�Q�)D��ዧ;�V� ��ފ�I��$D�Л�H�\G6��P�kǌpXd 4D���!Y/4_�� �5B@��#d3D�����D�M|�1�M��� �.1D��)��F����g̭N|4�u!(D�� �kPK'v�����%���Y2"OB́�/ӫM�%R$� �#���"Ov�[p�A�%C�,�7d	����"O(�uM�>M�4���#Q:�|r��|��;�x�=�}r�*��A�	
�M��<%C�hTq�<1g ��A��!��hB�t� 	c����r��O"	������i��c��S�4��0Kβ]�Z���=V���.û"4�*��Ptl�1SL]D	:�2#� clOpP$�HO�1K�o�/d�>蠐aU�]AZHt�w��ċ��=&xh�闐S�ӷ�X�Y7�D��a��u�|���t0%Q`�!�O���q.�$���I�n�	-޴Z��i5��b��ޞ<O�Mq!��U��	)����Q��ˈ/ԤB���T�$%<���R��/��sr"Oĵ��ɍ�xd�G�r9��Ui]����Y }>2GC�<Y�ȡ���y§� q1ԫ�9����*R�|��1%X�#Z2�`D�'��x�T�#y���p�)WQx�3Eƒ$n� R�E� ��b�EF?Pe.�	�!!RhH�k�+RXh�u���?�\ :�e�.b���U�T�h����Q��&v
���
�[�6!��K�(����z���PM�<]�ӢHЁ|� Ⴗ	�ߐ퓥@=,��zҏ��D �@�O'N� q{�^�9������"��\���4QM�5���E�jO�J�k�Ԓ~M�6�OR;<��ϒ{���"�J)$�r%��SD����/S�F9v�a�`�i�Z�j �j�h�g-|c��r��e*l�H��ݼC&�·xo�Ś��4*q��/T�X�C(G}%�/�*4���m�J��V�[�:����T��2LCĹö�dӨd#'�|��p9V��;q҆�@])�J�%�D8Cl1Z+Ĝ["iV���X�$(�J����晏d�@�qS.V#E���\�`��`Vπ�G�^IXG�2���>,�L�6�Z�� �ק$ې�Q�C���NKK@�)��P�AgF�L*��rgBОeҠT"��P&e{~X�4�/s.�ifM��S�aB�g��H#�����aԨT�	�C�@��Q��})$#Q����)T+�<��ŐF$��|�<i�C߸ez��$;J:��uEղ%?��sF���J�Ʊ���ϋYZN#"��9gp��+�9O0���U�'9��;���7�>���Ф)e���P��`��k�p>џH��T�&�R��-�&�n<��
w �fdZ+��YJqI�]���!�"@�fM��a阧�b<ۥ��w!�R�D�i?��:˔0 �˘��p1B�$�(O�D:S��;9̚((��X���x)D��&7ZZ�ã*�-�dd���C�-�f��C��b����1�Ƨ:�8�2L�
>.ȴV*���jx��,C ,�`��s���c�������-?�fݪ���5l�Z�S4#\0�M��'�-Y���ƍ�+p�d��N]�_tL�ό�o��:��F9a��M����<�`p��AP��z���ܕ'EF��{�� מ9�q�$�>�f|����
&��hs����@,����"Pț��n ,�F�#��SJO�鶠Ñk<h�H����MSӂH 8y�@���*/��b�H4"Vd�C��������-�G!�	�� �>���A.��1��<F|/Z�����/��A����Gw`�ѵ �	� ق ��Kb�k�'�_����(-�$%sG	�"
�<\rk�;U�#<q��]�SR�aF��Fq��V�u��K%&Dv�����^N3.��$��L�uQDGɘo����CC?Hf.´�i�� YsMY=�nH��i�D�"��"���5�jqɵl� 2�B�(�ռO�!@%�V�_Ä$zCJ�
f8R���i�`���+ؑGhH�R!�F�y�8s Jׯ+�@Q���N٥FA!]p,8�(ԥ�9��U�^n���C�W�Vy�`-�?���� Yy8ʓ;���2�ŋ�
�K�*)4�̒F�\ݦ�ΓY\p�C5��_�B���-wW�0���A���p�[*qr���dI�����c�nR��\�n� 5�-\;�`8f�Ơ4��9�FLc���Cn&�2m�'@ɤK��I$^:�H�ܽX�U1��[1v(�P�%��j���[�e�`U�5#�I%]=�`�VKܼS�uy�1t/0IA���ŀe��EP z��ӕDm*@��H��I�.& ����2O�F�̧A�6�ā]ˊyy$cK�gR`�'��.�
<��LX�C:�PJ^��pG�-�4�EYG4�TZ�v}�����A�X��a3��XR�Sr*س2��h!��U1 ��5a:#��k3H��?#��[\�k꘲3��d�U5<��IU$7&�!��&��%)�} ��Z��RIj��yfL�2"�Z� ��[iԦ2+��&D.'*�e@a����?�D��
���U-}��\�����?���
 _��N�O�^��4��� �E(�-}��P����M0\��A��dX��2R(l��1�H4X��p*�:��	s�W>ɞ`�p!E(	�剈^�d8;���dZ�Ę2�����KN�{�^|�+�'v�@�a�/H���ǌą-��Tzwo0��g돨|�J\�ϥp���s�c�;U�D� 	�9;S�9�t@�R0�c�*Oy�Hk�F�( ��J�0�I ��L&-J�����C�z�1A���%`д�ЁI :	9�]�'@�&��hb��J� ��#�y�.ā@VR��"�L�̔9��_>"���
Z.���Q�3��)�a,��{��E\���HJ�lj����:cp�U��ީ����p�IƘs���n6��갈�kf��$�M�av�q�6����0ȋ�Z�2���C8b���d�<��O&��@*��:<�RW5	�Jt�pN�/��1I�¡-`X�[�^�u�=2��s��ІE?�� 'Y!V&^i�k��gH�1H?�D��eL���U�4p�h)�$pu�� ϙz�ZAr��J�rdRׇ�	�������6u�|�m�&t}��)��y�Lq�M���<���ȍ�}6�(� G��-��j�R,=����D�X���㎟M�H�(A�p/����P;���$΅�D������Z��`u�N�M�@�P�K�r,�D>=qx%Ѥ�Wܐ𺆥� M�a|��״.:M��bޜ<;ͪuk]�y)0�8���o��E��i�b��SŦ��޻	�|�K�;>�Xt"��?t�@��ODM	pc�?U�>�Q5+�W��җ�I�|�HQI�c�=Q�2�iE�\�T���lU�=Ʉ�ԍ<�%j5	@�[˨��󋀒No@���"V����l�:9�8��&4�Wd2JC�Ұ��騥E�8p�sUf��6 ;���^R�x��?Sl"1�@����e��?�cu�`�? �]zp�%\V����T	
^쩣�$�0\ҥ�'���Rg+�,$MN)���;}OPI3W��,p�f�"�K}��7$�6��tk�$JB9�D��9xFDa�Sz�$���n5JOx����ɾ+�>= �*�A&�T�M�]�+��1[���͗�M��(�ֽi�8%�aE�d�r=��^���,�i.�I�B�|�z�A�~��D��+� a��"=��� B4N	��g<rw4`����3KD 
4㑉��<҄��sC�!�E�D�BK��0n#�p?T��*w<���Ʃ}��!��Ӧ5��B:�@U��;.a�Ѱ^� �cP�Q���iP%&�9�p��9f�8�b�6M�M�&�Z���>��59>�9 ��+Nu��{�S�T��P�l�	8F�����:3 �Z� p���ࣄ^�Ov��s`ӪP��)8Wي>K��I�	�E�ׁH
|�̍��'7mQ�|b�	�Q����<�A
&3d��� @Ӏ>�� J�!"f��43J�dN&)��kI!c�����ȅgJ !��I�a�2�hK1��	� lFDjF�@�f2�A�ȓx�����e��k0��5�B@;"kV`:��� l&�s�}��3���>��@ǪN�uMr�� ��">��X³ʞ�t��p��.t�<��+O�ГEC�	+٘	b IO� R\k$�'6&���m��8�"��!%f��a)�m��4�E(,�	/Tx����N��
��W坌#���b�g(<O���'���*5�H����IE�&h:a�1���!��X)@
���\�i�fS�V�%1����ܰ�i�%h4}�Ae"��@ �J7@�����ڌtEބ2�OT��⟌��/j�Lű�DV�쌸�'(�(!�V���H�[�uQ��+VA;3Iā[Ύ�CA�5�­9�B4�M3@kY~!�|�V�1!R��.Op��c��*��Ёr
�03�䉲d�.>>ԕ�2��-Ϯ��'Ip��Cc\;+���-���Ï)Kt��1:n�ݣ�A2MB8�ĤN�J̰u��K�=��@ŰLA�鴬���O@��� M+f��q[c����wFC�P-�8X�j�(|� �ĩ��~c0��bO5������M��������W"�8F\ [Dҡ���6�����a�g�	��n�AqaႳ"شS�O�Wy"�)`��e���
"Վ ��i�GB�Y�'"T�0b�Pw>�a�Qd��ODR�C�i�Q:�B�+_�U�~�R��*��QB���G�R5$�`��$?z���0��蟬U�Pϑq�<�%�ۘmLR�xc욕	��@��	X+�����O?�I"!��������v�8����$ ~�)2��YZ��"Giy��T2�'ۣ#����M~
��{�};&��H��]��nA���д������{�L�Q�ɎO�$|GF�24xD�������J=i�#Sg�o)J�``�J�m��KM26}PѦ��O���fʾ�Zc.۱�VM:#!��@�ph��K���]�ePt�C�&Z����ELdM �;�����:o��r�D D���.P��i�:Э�&<�֠q��T>�Z��P*�$���M��4���-�����:��e�+v� ��7(�I�La�.�_�ԄB��P6H� 9�#��c����N�~5|7�҂!�~��",=�r�S��M�&g�8鰁QIP;R)Ve�a�_�ox���[� ��BT�Q�g���'UzLȗ9������8��i�BmܥK�
5��Y����I�5p�(�:��'�4 �MS�pP�x�F�:b@��D̓U�<=G���Rc���fT�(F�0em� u\��0V�@9"& �k��,�o!,�̐hF��
���r��'Z؍Q��l��e��D_�9����_�,����-�8���i�O�N���o�{�����'����6h�@��(Y�f3E��H<A�f'b�IQ�@s�A 0(�!b�@���fy7�7?/�e���^h�(�$! �~'!�F*u��]�&�1VX���p��Y|�:��_le�s��)D�����(q��Q�.�$PH�FWż�����ԙ�#,�8s���g��@H<apT�b��ฒ��c�<|���*�R�6iN�)� 9i�o�] ��R�Կf����"�R��'
�M�'R7+x�!kG[	�:5�nT��{V���9�URb΁�1�Q���U[���`���� �.�q7��2e%�	!���	דp�HӢā$0����`��9h��%��� ��`#F�M: M�eA� R�WJfDh���bƐ#�D�9�Bh؎-��� ��G��B�I8\�4HB���3q4��[ǅ�Rfܜ�ժ�6�j4W�N=w[Jc�&:X�>XRØ?�rfJ�ڼEe_!ٶ���L^� �>t�2j�UH<ѷ�]1'�$�1uI�&LwLA����$|J�%���R�8q�T�T�y�Y�פ]�%�.�%�g��	�aI�	Ӥ�*d/$G�ͧT�H2�%Ű��O���4��4�\ѫb���2�[ѭ_�x�5���͜#��� r��e��53᧙Hn��!r�	��~���>�Lj��NQ��O��5�e�'_FL�F�R4L��(}B7A/�I��E�o��*�j�-&,tԂ�KP~���"���hxl��*ŗ� �k�L��D��G�~�XhiQH�~y���H�H@lȹ5��.R��mK�HG� �Ä$ƝY`p�E˙�E�r�b0A�3KG`�ė�K��Q��X̻�Z��@j��_g���D,Y�R0��OV�"�,V�a��x��|�=�1
�
r�p��� �l�H�"7��dyQW����
��6�ԭpV����Qv�d�xP�A�h�B�G�Y�ay!�KW�`uH�x�-�Gٞ��#ږw5��J&G	ؑ����)��i�t���-�9�V9ӳ�E#�V��5@�3����!e.6�PfǛ %��i�C3��� /�3d|�)h�@�MB֟&�����	;�y� �
5mЙX������o�2�[qU��1x�灹j�x�&���G"d(�ɟ?0��X��V.�	��"��;I�;!�\�63xͪ��8&8�����1Q>�8L����Q�ևk�xe�"�E�)����4ib]�&/�5+�F��",_�J�����!�j�xm�r-E�,���ݰK��)7(
|Q����V���4l�s�����e�*�1u.��Q��D��xZ�p���	�BQ�.�^����E����*T�?��M�U�ݝrL�(���H}£n�&\����g�}'x��KD-p@B�%��D���b�� �Q����,tIV�ص�� A�0�G�&� ���S��A|N�3��X�bl����:��Qd�U�u�ͨp	F�^����S�Z�C{N�g�h`��OD�%ce%�*F���[�Orr�:L� �a��l����H�?f���U@I�{�m�f	���s2/�*;��x��\+6�V4���!2K�!�3K�5Aԙ����
�dۢ9���?e�O�\AH!�"��Vx����v�\�(�#KŖ�9`A�E�t	��E	#� ��3ag Ly�9�U ��p Y @��b[Ȉ�qE�`.���gц�hIf��P�N8ړa,J�	��W>���c	�B80uS!Q�f�3G�>��jR5%L�!�o�<{�ؐi�����
UcP�;5��8����#-��85�V*�K�a,�}08�y�eC3��	9�ꅠq��H��	'�$��֋�a�tZ��YfO�`:`�B�h��a�H� ��F����:���k̘c��'��`���\�]��P#��P��=�rCӏ)�7�68_ġ�u�41Pjp�A�����h{%�ıA��D�!hX*-q
��q��U�^8KDj�&����bg������5�g}R��1�6([%J�3N���oС��D(0o�4�s��?A���
���T#|���RSѮ�J�BRDzdj��)n�,�E�)  0m	$�ƠU���{�'���9����r��%�󮚆Oܔ��3�n:���O�m���	��>�u�d�����JԒzVƠ[!n�+�4ܺ ���L!�w�'?ȘP�3e�����������C��T��2|Ȓ}P#�&�e�`��	8�
��'ұ�4B�IL�IAw���|D�r��C��0Д�ٕvF|�wA����s� H�`�)v4h=��z�I���-D�d;'D�4Uqڄ�\�aq���&	��$�b��M����'6���Ie)ؙY7N�0�J̸�0�NĨw�kӢ�9�-,��(:u��;\dX���"OBه��:J�Ą��̚7U0�*"OlB�GR�q��}��l�$�e"O��[6���1�1�ӐzT��"O�)�3��iNa0�O�0_�ܝ��"O�e��〸j ��Y�-Xv62�i�"O����"Q#m#j8��.Y4.�8z#"Od]�1,R\�H�-T7v�x���"O�E��g��R4�ê/�����"O��:G�9ֈ���<��"OHT�t��95P(�S;!K��Ӧ"O4��`�d��+��FgV.h��"O6�[Re1FuT$�ŏu(ف "Od�Q��_�8����#��Y�"O,4�p�с ����̔s(D�p"O ����T8�4��6(E2^&�1� "O�᫄���m�%�6��-С�p"O(I; ���`4�8qs��l�d\QE"Op\���N�!ݖ��A�YQ�,5Sg"O� n�x�r��A�-.�ŃV"O")R��E� \a4��%8.�%"ObU wEN�CJ�!�Q%�"&"O��K6�W�в Z"�#d~	�1"O�\��⒝ru����+�V���"O�y QmҫW8ؤ⥩ub��s�"OD���SՒa�VhV!
^̢"O�t[dd����� Ƨ����8"ON��DD��e��D�;�~4*s"O��11�D�^>���.�T�8٩"OF�b��#<Ľ��,U5g�d$��"O`�ʓ�R(���"���5�4�ɐ��+;�4���I�2��mY�j�<qg��`R�.e��"t�Sd?�K�wت,oڬBf>AzG���h�v���� �d ;�a^�A��(	7Fǟy�8	��hf�6��#(�%�������
l����B�.m��J���`pz�ЦJ*/&���&+$Kl��O�����V �*Kk 9�3��+�Lc�N(2P���F ҃�0|��(��-0.�
�n��Kb�]����j�p=�Â*@�t\�4�+zL���=Vְط��;�Pp��F!���ku-[ }����I�G
nz!	*�L!���
r J�G�&�jÃk����@�w1 ���q�uX���u>eXuo+(1@�n��X�h����O��R�t�䬂E��F}��鐐tr8��Y��)�
ʻq�XA7�Cj���rǞ�C4�d���:� lH�F7D�,P7��7=���(�׈��� D����ƶGZy�Cf��,D�c<D����Q;�d� Bܻ2���q�>D�� ���a^	}���	��U�@��	�"O �z�*	>qi� (E��c��E��"O���u�B�_�f@`u舻1Rh���"O�%�O�T�����f) ��a�e"O�e����%P��4�r��)~����"O����\�6�@�A4}4�\I$"O�a��Nl��t�%��(@� s"O<����S IO�Ѱa��`)2�;�"Ozx��! &1܊��G�T�b�<a�"O ��B>�\��]�r�h��"O��p�Ւ�(Y� a�)y�l�"O�*��S�Zu�A ݃<p� �"O�%�7OK�s!�{t��>h�y�"O�̚�k#R7F]��gB�{\"A��"O�|[ �n�r�	ĸ	C~Ly�"Ozu���9�Z� ��Q:xl� "O�բ���C����`Ŷtd y "O�5��D��� �ѮA�c�|Mc�"O�HI5H�#Y��7�\dH��"O�Ę�iE�l�"��Ϸ9IjYѵ"O���+4.�jh���AZ�9�"Oڬ�rl�bm�uLSu;nYR�"O@X7�L;D�Yj�+P�L9�H"O!��b�gx�=A]�""�A1�"OF��B3]�ѳ��V�@$"O:e�tc�h����N��H��"O̩e*�0ԪHQt�1x&�s�"O�-6nA�)�`u	�N_1O{
�)�"O4�� �=dҽ�k�o�`c"O!�ǑR>��R��\vDA�!"O&�(5.���e����,;[�Y�"O!1d¨3|�U���<e ���E"O��Ո�"E��kL��05t�k�"O�L�w���Q$֌�QL�:,��=��"OVp�ï>�-Xp넳=����&"O�
���Cй��o�+�Ԛ�"O��S���/���$N��b���I�"OV%÷��?0��)�ΈcĄxx�"O�0�a.	�6��d�NX��4�1�"O�ё�
U)�޸�����%vy��"ON���V��, Sdځ ha"Op��m�(�f|��GN�6��e"O��qP�5-����[�%��1c�"O��bq��Aɼ�����z�M�"Of}�c�$#M�ax��<�6�g"O~�*q㙨dpȁT)�7��Z4"O4�R�`�
~,�`gǔ&��� "O8ܣƂ�x3<P!q,� 0����"O@� aiۃ&{��:�e�U`�XA"OB�����%�f�²aY/���"OR��e�!8N�I�c �2a劰!"O,�C�ÑҠ%�vn��|��#�"O�ԙ�D>��܊�,N�\2ȩF"O��k�lZ�2,Be+!�ͦt�2&"O����P��Es7(Z����Q"O,Ps%DR5N�j�{ I�p8ސ��"Ov�R'(+^>p�V(�=R���"O�q�� �,u�h�8s��%\B�T+ "O2A[�߉Y?n���%/PE:t�W"O<E�u��N����3ꎩj�dl!"O��"R#�
4�pF��s��;�"O��TL�91�J��w����"OPh4��bKRI�T�<����E"Of��GfϜTy� �q#�5����"O� �{@���v�p�7x �Bs"O�iUn؍C�ĵ�Q�u �c�"O���T7?��Y8V�R�P���"O�)�R��.'��2�[|�����"O��@�yUF	ҧ�S�Fd�'"O�m!���4U�4�
Ϝ٘�;�"OH�4�I�(�Jv�Ys�"O�8��Ҫ;+
��`ޏiH�{�"O��bBE#F��t��iЁ��"OH;�N\35����u"܉UQ���"O� ��ʊ�{���B` :+=p���"O~PS��V�Mp�p�3�؃ML���"OZ°���BdZ�8�L4bE��
b"ObįT	T���1��MTE�5j�"O��� ��:{.Ȉ#ג;A �yq"O��@R��C�+)>_�Δ���Ep�<��ϋ"j� �p$ٽ�j`� �E�<a��_�|;����6CE�læ�_x�<I� e�8�7
O3Ai]��m~�<����A�T���O�0t,�(1@y�<Q��Q�e����CgǴ	��ZR�r�<�K��S�j$@�:��R�*�D�<�� �$#�(M��g�i� �w-x�<y�*�׮q� ���B$��)q-�i�<A'ċ�<d8��
߄#r��*ńMm�<iGk�6���F'@�^���g�<A��g�,���ˀd�4X2�`Em�<A��Y��mAw�4.�jX��Dr�<1R�A."�X�aÀ_r��:���k�<�WH���]��i͜^:P�R�%�c�<�ra��.\�����2ad�:G�_�<!w�F%O����N/E�!����Z�<9��'{p�Z��G�J0HX���U�< MX6~S�{$C#?z�Q��T�<! +	/u$���Ci�U�(!Q�bN�<I�j$X��T��KB�Z�^����
H�<)wC�S�&!��G�-4-�Q��F�<���L;��]CQ�S6%Nf�d��i�<v��5�
��!-���*���e�<9�
�g%V���(ÅK��]����J�<�w�����U�U�'���bcF�<���,9�g��9��ᣤJW�<��e������Wn�\ADi�S�<�f�ů1:؝�GdS\R8����Q�<q7&	Mh��Ӗ9r�P2KK�<�֊U6a)���d�@��#�@r�<�T�Ә6�h�S��[
P�!Q�F�<A�C\A�t G�ƴ#�Li�JGC�<�@�
C������F�ب�A�<�6�D���1���L�px�c|�<11���ŀH�(gܽ�p�{�<���6X�I�I
�M �Ld!O�<yI6_�*�+#������ "�C�<q���<4��!�	P�NA� ��u�<!5cJ����a�L>v��$a�M{�<�f�V%���5��#rdZd�n>T��R��Ҝ)U����QUnD!җC D�D"o�#t�P� d�.2$"+D�|���D�.qQ`�ڄR����t�4D�|�"��&j(!aB��I�G�&D���-�;�D�u��R�����%D�9 HH��ZIIQL���q�VL D��R��hl@0�&	W��y���>D� dc݊!�l�)1�Q�5� ��<D�� ̱(��Z�aT�|��hF�Zu��w"O�4��c�*he��H�%Ӕ}�>H҇"O\���(@��� �B\�YK"O8Fh�	춬S��^i,"O�q�d�
�A2�!{� ܘv���u"O�M2w�3>�z]#�`
��e�s"O�Y��ѸP����E���х"O�0#梙wa�@���C���I"O(���dԫ7A�r�œ4v�=�"O��SȂ3l��]�����!�"O���p�Ӕe�̓����D�F�Xa"O���4gF�b[4Z�.�}u��x�"O�D���ї1��ęU�	^h��8�"O��CE�0���؇�����"O�A�2��/��=����w�bq��"Oqѧ���V:C/��a�ȀQf"O"lX$˒?<<��.��H�J�"O��E�!,���|ɫ�(ý�yr���.m� i�a�=)$��O��y�٦eu��PĆR�9��}�����y�&^����r#��#(s�5�唠�y� |� azu���� ������y��4(,����Ӕl����y2	D��e9r�q���eF�yRh׽#^�M�e���n��HaciT�y���Z�����"Rv������y���?s��{$�Z�:!Z������y�j��J�@9&+\b���@�Ʃ�y΋�.PSC+ΠW<<0�� ��y�fX*k��9FmXA�,�'M_�yR�R(lb�NM�6R6�K�N3�y�؁��8"@~��i���K<�ybCݶ
��Gn�
��`҇�ybf�@p��"�V8��E�E����y���T> �+wD�+��i�g��y�L��][�҃M�KJ�YP�`��y�ᄅ�l=�SLگy�ؕk�y�&�.�pDJA��l�|h��G��y�B^�8��#�E-a0U����yş�2X@ĢV m"�,��y���TK|ٲC��">"T�r䋕%�y��^�Fj6�5a/R���!
�y"E?,��pJ�&�����kܟ�ybb�'	Ѡ ���U��X!�����yb�S3>
e[�'���Ag	��yB��0+������r
���Qݱ�y��j��bGVT�C��y2�� �.����8�F-�!�R��y⨜�4֘���7�h<q4O�=�yR$N0�`�]�jf��C�	�y"�B�Q6f��¢,j��	"C��y"�M�d�*4��ȝ�Ţ�����y��_�Vk*%!SO��},���E��y��?Jь��nW-<	U�*�y�F�e�B૝�[L��"��M+�y��υb�6�zt-͕Q���z��8�y�f�L_uhS��H���o@�y� \��pa(����=�2,��AB��y@ x��f�ńf2���.�%�y"�#)m�$����Y�^� ����y�����^�����M��4����y"*��
ܸY���7�H-9T��<�yR��+���(��:*�P�9����y����T� ���_# s�o�=�y
�  ��)�\� W�7Bx{�"O���`�Ҩ����$�L�/@�p�#"O� �pޥ+\����@(3�l{�"Ol��i�>�S��M."�Z�"O�H�Gz ��,�&z�S`"O؅�O�p,�; K%Bf���S"O"��C BF�I�f�<'_\ H�"O��Ь^8�� ��I,nC(���"O��q��I�l}���L0�]h�"O��E�̕f�0J���k�!�'"O��`�g�J�)!e�4c4"O��H
?��Q�!IV�"� �$"O2�c��٢oYDX��ȶzz��D"Oz@�O�g����gOF�X�"O��p�m.+�na�@�:���"O�i�6c�q�"��u�,^,$�r"OL�c   �y�& "̀6��[��'#�Dc(?���M2�5���3,�4IEm�֦��I��0Jr�Aڟ%���}z��Ǭ����hV%ۤ)a1��Цm+��^��M����?!�����x�O
f���S�a �*A��&�L$�`�s�x!1M�Oj�d�O�uF��':q�΀��
�I�M�</-$���pӪ��O���W�/Rn&����эU'y�ħ=�bY�Ʌ,"u�֙|��/Q{������O��D�	L|>r��J�ہ� +��m�ǟ`
��T���|ʎ���#A !�#%�#��`5`êb�6�'�"���'��	� ��ʟ\�'Rh� �Es�cH1��
׬N�;�F4#8�'b��韰�P��=����gnۃw%��� �.yƴ���}y"�'�b�'���'Pp�۟ ���!7\�9�c�ة!�(c1�i��	şd$���Iş���$�4�6-\�]�f��1�2\�2]�pj+�������	ß\�'W��Z%�~��[�R���ܫ$P�(&�>b����V�i��'��O%ڠ��ڠ��@�ЦZ7�uHDhX%JQ�f�'qB�'�R�H A5�Sly��O'��6l�VR>y����Fk�̲l&��O���47�x0�"�T?��gA��@ �	�
l�\��w���d�O�Q�M�O����<��'�?�����
��b��$���t�XT���Y�	̟�� �45?b�b?]��95`	��ɸ0����"ii�j���R���	�x�I�?u1�O˧n�$��k�& ��(�H\�]�G�i*(7�D򟂒O���/e^J8!�oˀ\�h�ڑ��=����O����OH�h�<�*���䡟�Z7�L�:�c"��8M��١h���'�:L�Q�:�i�O���O����k��=u
4)c��-*�H��@��ʦ�I�,3n�'�T�'�?�L>�.D]�lt�ʜ�
`�',9v�	�"	�Aг������4�Icy"-/y�́P���./Zœ0����禼>����?a���?��Ț�?m��30�O7k�DU�P(�+f$rY�A�|��'��'�b�'���kf�'e�� �W*�ZP�d�/�����x��˓�?�I>���?iB��!@9�mmZ�U��90W��I
�2����%�l˓���M�Xx4:çKT��w�[����!���c*���ȓBN)��NL�#��{Q.��Z����JcV��v� �*&��"/����w�e���ǉ��t.6�RC�M�G��"AA؎V���C`ƋK��ؤ�^%$x\]�6o�#:�L�
@�{�0���Fאb�L� ˑg�X�&��$*���7"Tp�y��%^>ap��F^<�@2!Z%Oh�d�Ab�
��Ⅾ:��f�O����O��9TBS#qC�HCd�"�>�80mKtQ�c4\�$	45)q+ΐ�dH�O�1��gG1'n�ݐ脩d]`��¦<wy֨�q�W)�"��3)��k��ɭR��pn
2V.����9a����%����c�IP���䙓��	�X��'��+����FX� @	d��<)@0�ȓ[n��P�E�U��Y�Ě�k�Fx�"=�S���#��9�
�vQ9QNנ��'��1�U��"�'��'�v���H���g�ԑ��h	o�^$@���R��PB��C�4���g) �P���?�=ٓ�S�Iy�0��(_?}��-��
^�B��.u��=J�@i�g�'��qKҁB<X���xf�E�t�0K�'��B��?Y����<�Q�	''��zg�/v�����	�Z�<1���
��`�[*l�D���㙓|������$�< �o�J����"5XX�/G�uY~����t�	ğ4{���Ο��I�|�1�	)@�>T���Y5g�"m�@ł�V����,�VT�z�_���<a&�K1/8|K��7�$YWIv�7��>)�t����-?N0��	�)����O�@�'xcB��D��"��`�7ړ��O� y�Ȥi�0���$ V͙�"O<4�� <5 h1��޺�Y�9O�=�'�I�55��s�4�?������8�
|�7�ԙ���;-c,H��-�O��D�OP��!�z������S0~���|*h{~MK3͂(~�� �W�'b�CnCC~mb ����9)dN�ﰴq��-��i��݀K���C!\R�'�%��Z��gl�"�D�|�$�KW���C��ͷF��02��?1���9O�iP�ۉ&�ڵ҂K�8Ln����'�O�\��G�kf���)����K�6O�rv�Φ���⟰�O$�D�'�b�'HT����g?����l��F:����XJ"�xd5�T>��|�IS*�M�vA:9���gƍ�BV$��dP�X��D�J>E���x���õꂵ+".(� ��	�rԋ�	��?����?������Ҋ]�{�UP NK  ���Pҡ��y�'��}���9k_"�b�Ǽ0�d)�/��O�Dz�^>��B�$�i  �x�����ß��K/��������Iݟ��	'�u��'4҈�v	r`�B(�b]������~�f�u������ɝcFB���	>v����ʐ>$���ńpw��I��&H���K�@<���ˁl�꤂q�N�N�ָ���ƃ$��Ռ;w��mӪ9l�V��a�S,,�楙q#ŀHRj��`h��izC䉥u�H��� �|H��3V������Ē}�Q��6��'�M� ���	:���� �Sn��Ā��?���?��t��8���?)�O=6x9�,�>�͙4��.��(��ҍ'�6��(X�~��X���'�����UIӰ|y�"Ğ3?$�#N�oTDB�.ֆK�$H EB�	������dJ�AiR�'����E,K�b��ѹ1� ��'K�O�}Γ3k�sʟ����K�ŕ?tTQ�ȓ�$KgC�<X��ӤK�>�L�����qy#U�N�7��O@��|RgOF��+f��89��[���	F�5@���?���=�`}�c������ �|Z����HA�@̕=�}�S�	6y |J$ڧD}li�B�n��a��c�<#�R�Dyr�Չ�?ɋ��@�s����Ƨ �h�0�g�13�!�!_
���:��('۔�a|��;�R���X�ģ	�M�xDJ��T��H�p�TnΟ���k�T�ؘE0"�'��
�	G� ��R��7�4��w��+`��Hi���'�ia��M9H1LqK5ͭ~"���;*����@��:���GEеUTn���9/c���Ŏ�I#��փ���>��'��tم��<M\���,�Cϐ|�Ai�O���"?�[��?��Ժ3P�Eʢ(˕'�^H�3#��<y����>1w��tF��;GH�z jR��A�'��#=ͧ�?�Cއx���:��Јn�@�Q�&@&�?���J	�\i���?I���?)��j���Hy������M:AfQ]d�ré�����*�"�4yaE��p<��b��*��sD�ɦ�\JaY]?!R�?@o��fg^
t��x����B:�j�#��Z#�� `�: *�Ð�Fx��'n����O��arX{�/L��YA>���ȓr7$� f�``$$
R�N'O7V�Ҁ��}�$[��P�o\:�M��	�6�xep�f�3[����#Ā��?q��?1���������?��O�Jh��O����ƚ�}^�� �Ɨ�Z&E�EXY v�ٖ`��0<I o�7$�:t3���('*��@N�d\�����$Pl
=ˢރDjP��	�-&���֦���E�/���`�,��D�"$��M˻�M���/3��<A�He�t�a��"���#��HP�<����?tH��Q�i>|�cr���<���i0[�(Q����M����?�*���#$�K�>Iq�%�p،�2�±9���D�O�����$*�|�&�7n`��eם$���ٷ�r�'(���ӳ8���d/��k슁H��)0�T�<!�N���IF�S�pƧ>sx���0%W4ef��T������?E��'�`|���%|�5�[g�R1��^#�'��d�gڤ(�A5�������'!^���{�����OF�'0�R�����?���p(��ڤ)R��t��u_�1!
�o6��'�>{h��Ȧ�'���?	dl@�t�)!BldQx|ˑ�_�@�� y��U	�:5�E�",U"%G���r ���\��qyg.4F�|�1��?yC�i���'(�O���',�A�D䠱��U� *sF�ֲJ"�'a�}b�S(�4��'�Q=K��U�uŒ��OP�Ezr��>I�MF[�ji�f
K#CؼY�BNݗ��xB�=9�d�)D�i���펛�yb��2r����Ψ`&�� "+͡�y�l9BvyB��U^���E*�yr��W�Z���@�	
򭨑��y��m���d�C' �N�pj'�y��*����F(�0Dڄ� @��yB�� 	�)b�k��R�t�1"���y�#T8a�� #P�4N��b�
&�yb�ϠW�̪F&��x��T�G��?�ybjS�\gj�5.��l�֠���ʄ�yb��fR��3�	�f���+���y��?g4��A"O�Y/���K��yB�_�#-dtZ��@�Q�l��bO��yb��.8e$U)���V�D��"K��y�g�]�.����	\0)���yr��8�&8�'J�$�s���y��@t�D+���%r/<��1���yBbM,i�Ldǎ�9l�Ұ
���y2G'w�,8�F�_k�8�P��y2 �g�*�BrbH�h�RYć���y��>��S �[8]��ICc)��y��F^R���*�9`>����@�y�a��.,F�p��6\\ޱar��4�y"��]��Xs��T1V�ٱ�o�ybh�
�R��2�$ Įţ����yr�	�w	�m]1
*P '�y2�1H���x�cB��,S'�ͱ�yb�%ź	h��M" gF��D���y� @l��#��w�� ��y�J�#J%���Vn"�9��>�y
� ��[S�ݴe�psj�g�\ls"ON�P�ʚ�
)n,����\�$�A�"OZB�[ E���	�K�fc "O�0��,��z�N8p��A�t��"Ofa�h"�������#�,� F�>QGAW+kǦX(��`�"~�#����1)��Ց�l�Q�*G�,���Ol�S�"W�?����r^K��x��˚8z�@�.M�mc��H�C�s�<��U�8l2�»d�T�2K|*�eĥ7I��長u��JE�H:l�(��#��HAP,�℈�4�����z2�Љղ�O�KGo�E�H [֌_D�60��%.&F�RP��xCrb#n���`dj��� ZԈWd�60$�����״"�Ʊ1��X3�(@D��?+oQ�L��$�-���<Aʐ*��'�"����6�>���A��D!��!�>n� iq�*y�h�5F$�|B63轢9�AB2V0��v�=����8
F�7B����фQ��IG�e�e^���eI𮼢!"ضn���ɨZ.PAф��)^��L�Zw��x�7��+�4��v�>��IC���S.܃}94M8g
���3�c	��?ٓO˴n`�%>�y�/��-���"�[�T�(E�'�[Qyjm􂓷N�\#��C�9����Ɩ �8x���UP�'��e�O)A�ltKGO�c�Z`�ۯ?H`�Qb�^�4�xb6*�Ev�ܸG9a��T
�K�"#�ɏ�`�Sv��p�8j���0�ƨ�V
"o��IF}���&ؠIeb��e�!�p�'�ּ�@dN�*�!�ς�l)4��`݉M����%j0jx<Y��jq���Dl^�]�� �O��睭I���AJ�p��PХ�ơt;|�T!|��G��#)���3���h�F-A���^��]�`K�:��a�Dk��<�E��7�����A
<�Ub�jP8�mc|�'��!�<[J��;�c�h���Z�� ������'�ƨ�����ħ;G��)]-s�j<�P�U��y �T,�(��(C4$!Z�-��G�~�C�ʜ".	2EA���Y�5��S��	Ued(zZ��$(0����(�区�<��I�B#�'r�=����)��u9g!�8Yr(����	�1�<�6�,���#�Z,ml�%�K>�?A#b^�*�]Y��;y�*%y�-Ou�.���{�F�?嫂NԜ@纀д�Vc����cKְ�=�L�H�ˎ�!��8y��D7P��ϐ�l�rʆ�g��iI�c�n����1�6�����#���=���1�uw��-_^�a�1.ʆ3��>�<qvRc�H���.>��1�o�#� Ton�y3��/z�L��̩?� �y�DR\���Qc�!Wszx9A��8;�@5"���Y�p1���S$H���I�NvX�Z�A#>s0-�'�x��4�`���EZ��o�%�b��?Eb�� �T6ݸ�lA9,���Xq�_ư=)��U����1n�b�� �A~�0�֩��|����(֙q9�]y�,�e�O ��O,Z��XI!s��;1��bs�͏ɘ(� �	3e� ��F7�u��P�_����L8!%��W�R�P��P=B�T�#�Ĕ3�~���o������቟~vŉ���n�9[�a�,M8���shG�(��
����Ѐ뺟�����AkL	�K�F^r�23��yYph�΄ 1<�~�a�-g�&���l�}@�jA"�&���p�'; ��"D+R��1�O���杻��X+����E�
|s�&U�*"��䋳v)zU��ͯ?̾�[�� �~�|Dk3��s�$U���K�Ez�!g�H�O���"҇��(�&�%?����\�d��1ۑ�N3�aإ	*ʓ�����L�$�0ٕ�^R��`��?�˅Hv7�z"읬+���!!�4����gB��x�jZ]���g�'�
�ZG,݄0o����B0{I�y�JX�H
����5D����ְYҸ�+Qm�yü�h��
Z�n�!�ۚRU����"_�qK��'=�n�r�f	�Uo (���D��ʓe V��O8�q+�+vK�wF@��͉70�*�k�ḿ2�2���'�.���%��a��QfC*9<����ҭ��ɦ�y`%��O��S5$J�w
�$9Щ�h%�I���V6D���'㠔z�/7'�Y��O�<�"ŕ�8۶�	���!<	C� �m�\�͓ �n iʃd�����O���Ȟ���Q"ak.j�����$�@��oW\���~�g?��# �~��e�B�b�̅#�NE����C�L��~R��P���a�(F0s=<�s�ȴ5��	�S���T߱bS�Γ?��,��l����](�B�9rY��@�C���S��:�\*���PU���@%`�\��"��"��	�e	E�K
Ur�E`�I�Ou��/D�M��x�t��!�E
Z++4\��$�1o�; �HAia��\qB9e �u{��}�Iz�+��^��������G,���?ёH>i��L4S�h8���k�q��X~R#@��-᠍/q풕�bB
-'5�g}Z9n���#��r���㉖1&��Qc��\x��z�⛋66b&jÐ0x& a��ߎ'���jg+1 "6	�o0&��ֽ<��py2�؈k,��HT�=�y8�՜1
�CC�'���J`%֠N�� Kޣy��0�g�+�b�h�<a�ˈyh��K:�<���|��w�R�����HӖ�뱆�'�0<��֮r�Va�2LO�q�.����ۂ�����b�@ƿ�<�p���y� �d|u=��W�d��:̔���W%hy&�'��(�/��X�mR��ۣ4�t"T�O���� %�$a��
SL	6(�I�uH��7� ���O�J���� b8q�@�5H��qHyT*���-�1s9���ŪYG�C�b9s�P�u�H�	X19�:��T5��Y��!Cx�|���p�h�O�X��	�q�p�s��J0Э�!Ǘ.V��HPw��x	c�A�~��h��܁��P9o�,�K>*�.1,���.Cet*6lY�$H9��PdȒ�y�-�%7����᠝�M��� E:Y�E1�`�S&ph�`�I�~��<"�G@4�f`9a
�O���'��ܩ�J�_X��J�ƿ{L��0�ڽz-��N��p��g�ŭ���WB�%�y��D�] <e�BFm&�\���A4�B�M O<Kw��Ș�M�5I����.��v�0�(��PDX�M�"l�O��$��#8�D�ƻ�` T��'/4N W͡,N  sÓQy�u
ؘ*�ds��@ ���Ow��$qB���pr�ăV�U�;�t�0�f^0c�:K��^(�^�G/�hOv�bW�N35���0��Ī-WP�%��̓ebQ�ۮ��CƎl*�k�N�>].�1��e5t��4S%@qCKF�094�(��7���2Q
T1w4dE���+b�TmҕB�o"���!L�o*.� RF��d���(;L�T�&��	&mDL��O�A���U��.?q/�*�.f��e�����4�!�$1���[��܃Laq����QC~�D�q6�X��T}r�6`��e�ѠB&�����߈��D��pN�]#�H�d�%��*TiLax��
��%�� &!�Ia&LUg\FI��*\�7$ �����C�m
Gm��K'�D;�
A�;&�[5�'���H����fn��͔�FB����O�e1�-�E�	���WI�Փ��\G�����MC�n��.Ġh(���i���xBaJ
F��\J�@�Ow�Q��-u���"��م$ U��G���D���鞜sj��!6�<Ս��n�`Id��lS�c�O<��X�h�QD �02��T��K��C��y��A����L�$�+p��	`D���'��K����wˎܘ7�ƽ� ��ÓL�����מ���"�_$��[H� 6�̥z����&�{A��U�`�L�K�|C�aR���<YA�3��0F�T2ig�$��XA~b���$Zލ�*ƓF����e.K��y"�ܺd�r)�'B�(д;�F�ʄ�Χl�<�ȓ�jM�5-��VJhѢ��M,�N]����&S��j�
��Ń2�Շ���<�6���S3�ܶ��ԉ� ��m`L�$%\c<Q7�̖?7������q�D��dfH�q�0D��M�.��sú�9�):Oڭ��+D%D���N� :D<�@��j�'vX (�2��cf�Q'r��A�u�����8D��!Y2��eZ�>� [6���y'H�D�;#�+x����v���D
p��(V����`�|�<�����n�`���CD�a���x�t,vS!�"�����Vq��O虚5�^lh0Q�B�ۃ`��A�����tÂ�O�<:��5��O�:mQ7��?Fhh*`�4�y&��65h�a����b��M�3��pԧy�K�R
8�RA��]8���)ڼ��~9�P�B�=%n�$?qHg�C�9-��N�B�P�LK1��`˧J�Vz���$/eJ���"�<*�c���O��zc"�/���ŷ'&H�NɈs�RA�'G\�h/���L˧x��sŪ��y�ݳN6YU�εv�*Uhe��$��	�+m"T���X�	.��y�a2�O�T8`CO?.aĩ�rfƚp�r�����>�ԣ�F�8*o�$�E�X=�%��tj�P{7k]"��L��5q�X!(m��Ze̓�J���Gi���{"�yӐ4�VNΈN,8� ��	�4G���'IbpȒO�$z�h�Kg�:Nh�C=O��o�2t0Z���%7�����W���ݴ;}0w�}�$�g�40Z�穠|��iw:�D��U���CE%{��rs�Si8�<���ݟ�pA�*v����dg]F�l��F(+S�D� S�Hv�cPŗ�(���
�HO2�c7�yH1��C��7�RE�0�D�;)"M�i�ihq��̶a�Mr��ԬW� r��;���&cr0Q�W=O��	�S�l0"%;Uԭ S�x��Z }X$ B�#�0�I ���t��҃Mt�剄���}�  w+�Q�����?�R"��f ��C IցEa����J\�E��Ծ2� �8� �sP���Ƀ6M��sCK�!�x�%��7E*<j��y�ρ��\ JЁ�����?���U�󮏳%�� �d�C�;�Ȅ1%�O)�9Y�Ny� ΄~ͤU�� ��Ń�
D��U@���x�M�5	C+��B�f]%$��Q��6Z� �����<8�
��y����|�&M�.s�p8�&����'p9�"��4c�	z��9O�VJUh^��@�Ɗ���B4k�D��f%�H	���(VZ����Z<Fi ��Hq�dޘpe���� P3>���J�lΫ6��SZ*�ʓy/�ɬ�<�R(Azl��0d�i*�o=���N1w�dTK���M����3�:�+⦌�*�@�RǓ3��`̓�9�T� �!�*HL�8:�a�KV�	�t+ 0��P>�����^�N+$@G�S)�H���㏹n��D��%\� �F�f� ����~�c��WJ�i�`+�,1@I�u�F|$󤬞�H6�Ē!n�y)���h��!Ēxm�y*���'��x(���$|�i���O�YPA��Z�j�ㆀ;��[��Ɋ>S,�$G��D4�uK�}���4"�X�p�o��t*�I�j@J'
>��Y�B���'�$ݹ��Kv
8�O"~�Jc��;Avt�ï�&�����i��x#��_����,ˡ9��xRf�/D�N�*@aL>kVI
��oeV�@ �����"i�d `��Rޟx�3�)� �P*v�]V�``�Y)r6DA��FEH<q���_h�ix�CЛj@�Y8��V�<i� nC�\+BD�0�nq��A�M�<�5'��v�Y�#(T�CVf=3GM�d�<�ao
}ۘ��r�Z/\f�`��h�D�<�BA�4hJ�����4<ۦ����}�<񓮇� �ʔJE��}�H@�Qo�<9�;]����p�9�pU���e�<���C��Yxq�Θf�}���j�<�r�Z�>���W<xz���� �g�<��@��Mh�C׫�5-�h���`�<�q�ˉ8�0���5BxH�!q^�<�g傗K�Lz��޲so��I5(X�<Y���(jc�pp����=��9�5�PU�<�R�v�y@֥%+�XI�O�<��	]���F`)%�tb��c�<ٖ�ˀA��y��[�v�V}���Ew�<��	
1�^��Q�J���0�
�s�<i�2a��ꗁӇZ�$�!s�<�� �
r�� ���Q��,�Q�Ap�<�&�u�l�!+��Zx=I!�Xk�<�A(��p?�A���H�� �Ae�<�&k��j����P�oA\�R�^�<9�I�(_�l�:d$�&;�
�ŝ]�<���&x��	�Pg�gk$BT	Xq�<y%cO?&U�ժ��x�Ybab�j�<qu�+��I��ޅ|��5�\e�<���Ӄ_���e��"eq���b�<q�S6!��	K�¿�qn`�<9�.ȞV�$�
>�����_�<�n܀ZJ8:ak�.z��MI �UZ�<��lT�c����Y�]Kz	Q�A�n�<A��7[���Ă.7�t	�'��P�<�g�Q�'N|�2UGS�2$T��d�R�<��B�>�㤩�&0��)j&,L�<)%�/#B��'o֢2T�Q��F�<Qgj�S=�����ŊEv�ق�B�<���\�:���2WjUA�j_�<$j�zk�@���\�MjHI�� b�<�g&��H�D�<Z���Ї�`�<q"Ś/f�E(�.V��X܈do\t�<�/��}Ψ�´ǎ<LN��Xp$�I�<�qɎIRz�C���8���0��H�<QS ���!�D �,����E�<�R�%&���҆�%h+���g��B�<� Ӭ��VK� z�nq�(�h�<i�B͟S�LUz4j��BXۗMj�<�!-ӻ:f��� A�����f�<��脾s,�He�ɧ-���vl�e�<A�Ί�C� h0��$�J�w�F�<���1uF��6�ߝm3�H1�o�w�<q!"���܍�tiqkxP�CH��<��AM](���J�S���Tdt�<�3%PPpF�{šDؖ&)���s�<���֍�������p�T��,�r�<��El�����><�]���p�<��v�b7��� ��q�
y4PC�I�dڈ�p�/	/Q�ܝQvd�>$�C�ɛ"�J�Yc��5{��9в��6!��G>p�l	��H�P��@ku��
e�!�ě�a�ȫ�@�/*��`3�ZT�!�d=TX�uh��pd��k��!��'KF�C�ʒ�yf��*-Ɔ��ȓq�T��Cm�YJt\��`�U*����S�? ��$i0�83�i��w��p�F"OT�A�K�9s&��+���Y�"ON �C�ϰ8, ܈�+���1�"O���'��t��|𒥌%�J�1`"O&���D!y:^a)%/�0�����"O2L㑁��7F�|��P2R*f�B"O$��٩7W��A���B�^���"Opy�`��g/�A�կY���A"On�h媃.w�T��D��rc��"Ob!�7@�^^T���i��x�8TA�"O��s!�"}Fұh�i�3��`"O�$���'`�ȵcb��_���r"Oڬ␇ַ0s�\c����z��8��"O����X�m�Mq��]�ت�"O0��)�:<M���(�b�s"O� 룍��(ơ�㉈�N`i�$"O�$���A�lV�akW���a:��'*Oh�;�`'�j�{B���,���'�����L�d���Ҷ	�|Q`�'O��"�*6ɪ]����:��
�'^n���1i6.\�@C8t��c
�'t�ݸ5˗9f�Y�f�C�*b0
�'5���S�UrB�Bu+����	�'���ZW)M��e�O/�2r	�'��8R"וk�V|�t�_V�r�':�k�@m��	�J-wbQ�"O����9I}hPegP6_N|`�"O�a���ևH���kί^X� "O���"���8���ӊ�)*�J���|��)DҠ'��]q"	��	B��C�Iu���X�.K�/R���4`
��C䉾:9<��셤e�XD	TC�;P�C�I?_���;�i�/qyp[E�s�\C��+u�~�)V�L'l��5�Gi�"'��C��,R�بS�69���s��H��C��/��5�9Zgd����د~�VC�I��n��f/K�2�NYH��'G�B�I;q�b鋔oWf��TI�� *�B�	�&>|�S@�*\����5��a��Oj�=�}Ҵ�[%`&np��O
@��*XY�<ّ��Wx�Ӭ��_;�(h���U�<��lHN�Z�H�:T8�SWF�T�<Q1O.c����K:O:�k��TO�<Q��*��<��!"&�$"��N�<�k%-��+�MΤ*���1�  F�<QS�[�k������+t���AlTB�<	�ȖcH�t��o�f6,��1(\F�<i��A�����'J�}.L�<�����=�G�*-Wza�㋟E�<��pB i�䥃D��AQ�SW�<)�,[�x�F|{r@�."�2@F�T�<�7i�G��a��O�&2	�r#M�<YcX�>N��+U#fT�eR�FH<��ǵGs�[p��?o8��U��1!�L�M��!
�g��d�E��O5@d!�S>�ʔ��:=�`�b�#C!�d�0`j(����$<��V�H!��
?j��C�i�!�h���*ռn6!�R4`�r��g���m�6%�S$��J�!�$���[�,� ��T*�c�U�!�D�������L��}�U��7!�dS50BН����_��	3�E3!�$����rb"�8*��dp%"�
�!򄘺eq�a�������[3 �!�� >�����Bp��E�#0zH"�"OԘ;�+՛:����ӫV0XJP�
�"OD������4�;��C�sܖ��"O��vN�5�J\��nل���� "O�5oV!}=Ɲ�r.�4��Y�g�'h�I;v
� 7�<j���#��:`B��,M��yz�'G2�΍��K8NG�C�I2����4�E>i�e9��_c B�I�A4Up�j�=]~�z�ğ�`����0?9��X�S��av	ʩ�^p��eTL�<YM��7ft9jw�Dp�eTJ�<v�̲:E�(
q+C�$k�n�IV���O8�y�Ȍ{�	�0�4Y���{
�'Ⲙ9�T"NQ.z�K�.|j��
�'��$�Egݱ@Uha�a(��	=���	�'�����B�jK�}\hE+�'v��W�u�@�0%��?oа����'T��rI�	O�f,)�Fޘmg��8�'Nj�c�j�(��8 ��b�:� �'z�̳�c��n]ҹ ��a��i�'j�"�U�~7�X���[x���'�|���
�5�r�H���i��]��'�JH�2AWA��y�@��b�����'�@]��ݑh�8���(���tp��'�R���b�0Ext�*���?6Q���'L��bD�Ih� Dj�5- ��'$�I8Gh��<S��u⋛b�r��'���/��'����ϽB�d��'D&i
�n�3��(b�߶&�VM�
�'�Zț���3[�Pɑ�I�%�����'ou�j�&+D�g���p"K\�<��Ǎ�40��"S�لL��eȂC�s�<�S�U!5�B�9!��FW�� �G[�<a���P���	%(U�<���QS�<Y�@��	5���%�RB{�<���!{��b�C�s��ʵ��b�<�R��|Lҝ�5L
# >�@�ZZ�<��!��Y���N a�%���m�<�Ӌ�W���#�@S�����-�j�<�4-��2�����-1��ȳS!�P�d3�O9��"�(6T2a(��-}� U�'Z�]�-���#�
ND�m)� � 5!�ē�=K�8�$G IԊ=����2.!�D�V��I�0M�d�z��ac�,#!���TL�Z�"H�\Y�X9����?!�� "�L��t��AG�i�훗M�!򄛬��-;IE�8�X�+R���S0!򄈖@�� �EK���0h�q�Z?H!�r���\���5��-�����'4�|[��F=0�+��F��08��'sF���'J�l�)�E�)EHP���'�~Eړ�F2�6���F� A!`L��'�`{t��yE�pS�bY:)��H�'�b�ɗl��G�
p�s�Zs�:��
�'�ވK5b_�A�^��u,�,i�2	��'bd�
 h�'�+��ēe�0K
�'������20n!�c��+~���	�'�N0�t&J)=t���B��:����'�88U
9t�xc恧8.v\��'�����	CZ1��M1NA+�'��Y����+�>E2ଡ଼�[�|�����X�L�, �f�P�Pe�k�!�!�dK�*�D��iɇk������:���Gy"�@r��5\{@�:�) .�6)��"D�� p��`�|��B���!:��z�"O��D#\�m�X�����F�(���"Ov�����}DtE�%�  *<"Ds�"O�A�'˧J�,@,�Y��!RT"O*A��e�,HF��k�dѐ�"OH<{�F�S=`\B�e�o�u2�"O�Q�t��#g�}��.��p��"O�냇P& O�<2$��< fy1"O�y@`L/������F&0��"O�A��GY�^c�A�\=(���"O��ի�.L[��a��*5S���F"O�l����'v"VxӇb��"(�"O�AC%ԇu,�t�O[m32��"O�\�pE��&�(��D�{H�M� "O�\��MWse��ѐn* �"O�T��jY�P2<|�m��	$�S�"O^���G�K>v��3��K��1�p"O�!��H�;V=pˁ�Z�2�[�"O|�i֢�7ٜe�����֔��"O�%#R �L� ��"/�%q���"O.���J�-Z�h���4Ih��"O�<a�N���36m[S	Α2�"Oֽ)�'##�D�{��S�O:�qE"OtYv(�5e�\�'oL�b�\��"O�8Q٤z1�s5�'4j�t"O~�H�Μ�s��@��U�4"O~U�2�ʜ;�^q�����^��#"Oj̠�Yr�0b�)ڎ��"O.��w��m��)��N!�ZuA�"Oht�-�\��9ڴ��%�>hا"Ot��3
�2�C0N�:���C"O:U��MO>�1`�BB/#�8���"O �5�Š#��CL	�f�N�9�"O|xp���HuS���r�.���"O,ar�$4C��a����i��WT�<�#c�-3�Aۦ`T#zrH�7�e�<Y����m騙�u����B�&��y�a��3��l�@�_B4�9�$H$�y�e��vŮ	�R� �0]�  t���yBjo}�5��lK�q�Ty�E���ybd��Z�|��HC���h�뇓�yRj�W��Q1)�4?��qy�H�9�y��E �J�h�L�ijФ�S�y�Ø�8�n4��q������K��yB'ܥ{p�Y�Ѡ��a~�!F��&�yr��*.*�"��	�X��9��
��y�D�_�T	�ҬMX�F18��y�j���slΈhZU�B�%�yb�DWv̛ %W�k2��)����yҮH�Z��l���.1��y�bB'�ybnK��]�3nݒ/��T٦	ѩ�yb�@~�<�'H� ?@y�Ȓ�y��R?J��HC��ܬ8�6�rt���y�WQ��()��5M�9A���,�y2�@.��8+�+�8B�`��3�=�y��0Zp�����q`�%�����yr*�X�~ ���Z�4H��`ܓ�y� _�p0P! D��]q�逹�y�ȝKp^My�ǅHpf)�g�Z�y�P;x��:#��9����I���y"��v+�%�DHþGό=��\��yO�G���ed@������4�yrm��a��[6�:6¾$����y��(y����'��SU����y
� ֘ڗ�М�`�ش� �(��"O�T�$�����u�S�^�hI�"O`(��B߉X��Mv�B �p���"OF����#�"Z	0H A��_�<q�ٗ1c�1 ��IPD�2���`�<�B$�,��HXd��;Rt2`o�c�<�ƮX" p��̧	*�)��b�<��拖#����9 �\`@�L]�<�'a��R�`@�[7CN��
S�<����W3��Qr�0SgH��TO�<a�gԂ3��@��#��A2# 	M�<ё'�L�|D�B�
f\H@���`�<a�M�zU��R���gYq�<!��F>:"�i���(
jT��/�n�<�bFG]=��/�0b<����T�<Ѷ��I��b���cw�8k�o�U�<��蔖x�L#Ɔ Hj"���)�l�<	Ă@
&�9;��ٌ1Ƹ�ϟr�<���UM���K����`]�J�k�<�� YH"���ٽ�(Y�Zi�<y��1E"�viG�����c�f�<�4K�c|�-#��՚g�hH�4c�<Aq��Ii� 2��>l�ډ�pE�[�<駤H)Hp8ySi�#UV�-�Ԇ�r�<ɲ�3\�����cW(k�b�[p��e�<�V�P�
rD��E�,>3���CLF�<1i �
���qъ�+7xۄ'Jg�<���� ��M1O�>�鵬�X�<Q�Ӎ`�|"�mʃ;2Rm�DB@`�<	bMO?6�J�P�ƿgg:�rgj�Z�<Ap����(Lb��6g4�%��~�<��#ݚSj�Q�rJK�pr$��1�P{�<!�S�X\~��C�K��P(z�̂N�<A���AF�H�abZ r@�^q�<1�*��l-�!��	CO����[n�<)�jP�P����Y��Ѝف��A�<���
<��0�w�ʜ �$@}�<��A�:h��9ՋY�U�\�$B|�<����� �D�B�^�J0��F�Py���%Xu8�:Fe�q|^ur�e��y�d��u�h��,ӉS�n%#��y��L5!�f��G�I��x	�GA5�yb؈��v��"u�� �ˏ,�y���7h9d�ȼmO@�1!���y(5pZ1����OLC#GV��y�A
���,i3F�`��Bo���y"���O�FL��K!Pqؑ��y�gH��b��a(���9�"#�&�y�HJc?0���]�qzHQ�\��yR�Ƌ4���9GO������ߪ�y��X�}4p$�j�0k&�#�o���y�C+֩q���%/~�MIs����y�
W�k(����ϯu9�i2�oʽ�y!F]z6a7��6 :�C(��ybd�:x�tJ�kP#*P9�����y��#AL�±-
�w�8��`D�y�b��e�,�*1�6f���K1�R��y��ݚn�Xw�>Z��(��yB'�-G�$�c����8
���y�J] F�l�#���
Cݜ$0��K��y2EH24�"�0��Q�H)8da���yB�&X;���5'��V$����T�yb�Pl��,9�kXLH&�y���yrK��o�pʒ��SѲ�v�_�y
� �*�,��"G6��G��Oł��`"O*����X����
\cZPW"O�9iEա*
�M	Q����x�<�耹(~ ���HQ'u�^I!�B~�<9�,R�6� g�U�d�P@�Ey�<Y!� 7a`A�3 ��h{6�%�^�<qf�ܻrz��O4U��ɷ"G@�<�ႌ�
�E` ݅d~�U�[{�<���H�y�b���<2�<��r�<�_/Z���A��'�y!n�B�<�՟[��<� \�����|�<�V��/> ا�ݷ[�8hdJDA�<9�f[	Ha��L������C�y�<'-G�C�ּ��-$B����}�<q5Α#�D�3�m�.r�lȐ��_�<�r��_�Z�c!��2�.@T��Y�<I���I�B��q䈿gM[��Y�<Y�cD0#,E�@J=7�.�r���}�<Q.о'���Ea�1�*�*3�T@�<�w�,x�|Ҕ��#8~4��|�<���480R��	�}�����y�<I7jG3 cnEC@��4��Z���s�<�"nY:L�ƨ��L��|l#��q�<1*�9H��MP����b��_n�<�Ϛ�S!�}j7n��?}��z�+�j�<���ǁO�PEY�H0$���uA�^�<Y���\4�Y3 �3I�Ƙy��F�<Y㩕y�,�	�ǅ\�"��@�<��=vzٺ����&� ��A�	w�<	������p��U撨�F��u�<��F��ѨMK���0y\i0�̈́l�<�f(�2�(,y�Q!s����%[l�<��2Pe�Q�­\���� f�<IaMP�r�n���B����(Kf�K�<QEJA�;������ܢKA"f�l�<���>vŊ��Q4 ϴ�b7�p�<��i�N�&��`BJ%v���E�c�<q��X�P��
�Ȅ3�,���o�^�<�ů����&BO�Z�4h'K�X�<ɲ���Nu�H�e�L�H�#2!T}�<QS&C.�&J5��Y����S�<A��a2$�d�IlH8�D�[�<y�@cI�<��>�d�1��JX�<�ѡÒw��=$L�\ t�qC�[W�<٥'ΕF�$0	�GM
D�IJfG�T�<����ߎ��d���l'D�4O�P�<	�Ɂm'H��"�
�h4z�
f�<�w��cZx��L�gcܨ�V�R_�<�P�Ӱ=���X���<|���uU]�<�1-��%%��уh˶LV�rj[U�<��K��5I�؄��9,�a"$i�H�<��%ݼs���H�,��hኍ"���E�<�G�O�"?�[�Ȅ�)��܁ao��<���� �>��\�ac[e�<��a��*�x�fػC4�% �_�<�t�K�>����ܲ��0�Š]�<�v@7:����'&!X؝�g[p�<�B@;�p�cn��$���䇝k�<W}, e�F�	�C0�Ph�<1Do�(Ì���U�3�!xE��m�<�� ;Q5,|㯊�>�~U�!MMR�<IP�	/6�м�1nPR�*�� ÑJ�<A�N�R��a0M�A��(ΗB�<	C�
�U�T#F��Ӷ��U�<�  ��ަ�l����+�V0Cf"O �gg\�b�<��`�%'8��p"O���%kE&1Y��WÇ����!�"OD�@�틃>m:��#�w��\��"O�y�Ɗ�n���!"�}��13"Ox���A���MZbA��qx��R�"OV��b<7$�H!" ���a��"O����H�� !��U�J��"O�(�����,TT ޠ4w2��6"O0��#�Ǭ'��}xu�Wk��"O4�*�[�
�x��M\1Qa0F"O:ujc����U����B^����"O��ٷ��n�0�`�ݭ>��1�c"O6�jU)W(�X���G�<8���hp"O�9�ăD-tl�4g�~|Ψ�Q"Ol�ydo��M�He
�#�����"OxWI�:�H�!�r�(��"O9(��^� a����6n*�8"O���hQzOف,V��r7"OL�;ŏPf�)X��V3I0���g"ON�9��Dz�����A͝��c"O��e�&3>��°�4!	����"O�)gK� d
�,C��3���Q"ObD0��1fz^�J�o��h��"O�Mrr��&C�Z�;��w�@�"�"O��a���Te���7�*#�@��`"Ov�;��G�6���p5.����"O���0�`��B�ML�"Oj8�rj�4z*�YA�bP�^�����"Oh��6�A3 �a��%RU�=� "O���@�vrfMȱb��3�l�4"O��%',���7!��W^�홐"O2���+c�2=R���{ft�"Ob����2W�� � DƘ��"O�q��◇K�y
�o��;�V�j�"OҨ�"��*j@�Ԋ�F=\|���t"O�l�d�ߐb �i0o�ǮLQD"O�YQ�
�u �+�p�l3�"O��1�O^l�y��_4��!�T"OF�H�k�*�25�,�@u�s"O"\A��-��,z�&��:�yb8Ǝd �GN��Ҁ$^�yҁP�Fa�I�)A�q����P��yB�M�Z
�*�+H�"�
����yb��fv.@s�
U�>���G/G5�yRCK�A�:��S�
#o�4];��ȓwa���r��Z����`�ѳ&��Ň�5\��_�6�$��Z�� �ȓsc��Yw�^�K��X�ǉ5!�
4�ȓ������=F �t(�� HF��ȓG��DI$֫\�tXw(ݓ�0�ȓ%��ꕄ�U�VP��U�z`bć�b80<�0�>bu��[���D����ȓ	yTQ��E��]�!ÕW�|��j9Td�V#�.I�{�����݆ȓ^<���ъ:�*mJ$�"rxe��bpT�t�UJM�d�;j��I�ȓv�4]�e��w^�D��7$�l)�ȓgnH�� N�xl
E��N^*U�����9�k
G��U$�|Rل�3}Z5�T"��g*�#C��w�b@�ȓF�@�C�ÍX�~pc���1n�݄�A ��%%޷-�|h�䣟�2 Ԅȓ�`1�6O�4zt�!�ǧER����S�? "dy��Ѐs�v� ˗$! ;�"O�T��'��h��)��2$PPr"OT��W��(N�,�lB�0�
 "OZI��(+b���+����K*0��"O��Qe�ˉ�����Q+j^��"O�ۖ���$�0�!ي:jR4��"O�5���W+d\����rR�:d"OfT�$���%<d\A��P�]�"Of��!^W���C(ك
Q�8�`"O��u.(����F�EV�1�"O��۱�LI�Ā���]�8>�T��"O D���Ҟ ��eQ�IO14@x�"O�m`G�Z%G�� ��73�UY�"O�!nFWsvd���8J02Q�C"O��:��ݽ6�^� �mD=&}�2"O��C��0�d0��JZ0j�5��"O ���	�19���@�гR>�b�"ON���'��2����H�)
!�dS
V�B=�����L�d�$t�!�P�c	�|�h���$K���!򤞷?a���)6�Nyz�J��!�$H>4Z����	6.d0D��!�D^��� ��J^;6��%�J/!�dX,=� M1�NU&( M���7 !�$�("���R	�b)�����|!��<p�H3����d<�5�5	�!�$�35�v=��B����h��.#*!�#��ŦT�~A��h�>�V�t"O͓���;#n�DQs-��Q��"O�0�R��+��B���%d�B�!�"O|)���Z"���qǔN��TBe"O�A��B���ʌ�� �~�bI�"O����h�G{�i�W�Д]��H$"OU�p٠W �Yb �"o�r�:�"O,IH���:�8am�!X��`3t"O|�
���>x��<)���a@^YZ&"O�r�Dɓ�>51��܀��05"O,�P��z�\��,��0]\�CP"OШ�n�9��3n�1&�R��"Of\zhE0d0��&��:8�8��"O�[�"I5Xċe���A0����"O΅�U�N����χ~*X9��"O���woC*r�6Ɗ,7�D��"OTe:����Z$� ;׈ʉ	�A��"O�R&�އ.� �a(��#(���"O�A��	\D��%s�	�w
�š2"O,���J�<��@�O�pũV"O��L*T��)��H�N���t"O��:�,�Q�l%� 쏛qVĔ��"O��2G+��[�H1�3kS�D@n�J�"Or�(E�12`5qvJ�X3�t� "O�\뵉Z_���I#{���a"O�9��)P��abj�2 ��s�"O�׏֪s`Jh�t.ė �X�Y�"O�4v�?,�p��e�$�P�i*O"��5j�%!�(
",�Yz�'#��9d���% �F˖�$I�'Ͱ�@��в'�
=  L�Hm��'e�\�0��]�j
� ɬ�z
�'� ���eѬ|��YSC%M!���	�'������rv��A���9%�@�'I@�nϓ!� `�R��.��h�'8�ш��3C ��6�U�x}
!��'JjH�t-�1b�iW����� h$r -I4'�(
�産*��}��"O����W<ws�	:�ŕ�V��"Oj�{Q�؄}�Z@�;[h����"O�|��Y'zm�է^MHF=s�"O*��
�}���s��I��y��"O�5�E�)�<��F,�� ��8�"Ot�� o( i���(l�E{�"OJ�b��ע3�Ɛ(�%[c����"O���MT$���C% p鎸qP"O�$:���e��A3�܈*���"O�9I�R.R��F�gu��9�"O��p��)rǠ����\M�XR"O����I,%��+��`e�=��"O�Y3�C�,�(5���9Z��"Ov�{�Q�R�:�k�"�*�
=@�"O��8�"P�,�(oO��]>H�B"Om[�Ò�i��@ փ8�m�D"O�a��
m��y�W���3�^��d"O�0s`f�R��XZ�ٙ �8(kp"O���Lɒ&�ɉ�L'��H"O���_	U��A�e�E=A9�"O����+>�MH`�&V,x�t"O�1�W��ND����ɩ�@T�v"O
��j��vόX���.��\��y�Dz�x	I�Dk�p�T�-�y���:}h$����?ؒP0#��yB�=v<&��6��/ٸ48b#�yr�ŋ=� y	B��/��걩
?�y2��K��;��߳f�J�Pv%R�y")��f�D e�z����y�B�Z�PԱ4o�-RQ��+���y"�)Du��%������jH��y�� Q�:9�3FU*Lϸq)u��y���H��(_�3�����y2č�>�j�_Z\ȴ�"ː�y�GUj�*%��E_�M1���d��yRI$S�2�!�؍O�nE�6��PyBΛ���PF�	vRR�a'�\�<�gH�e��݋��%�B<���|�<�"o��s��D�
'qt>y���o�<9�ٗCW�1��T!K�
=CT��O�<�T�Gf�GEՠ���V��_�<!��F���������B�l�Y�<y��?Ǝ���u�abei�R�<���V;:X�4*�i�*@�sD�<'燝U�����1frFp�r	@�<iW$�
2����#�J�z`:�(}�<�aLN�e�HE���D &�ER�fWu�<J�L����FB�.�0B�o�<�$�íf�*�r�ºA�����@Hi�<���[�$n�q����y�T���]f�<���*7�E��f��n�p�b�&�`�<9")�$	<0`I�ςtP���l�Z�<��F�3<��Is��=T��y�m�V�<	p��K�$%��
()	0�pE�R�<�`eM�!���2�%+��-�D�M�<���qd�u�&A�)6�IJ ��n�<E�^�H��}�,@%Si����Mr�<�q�$Q4f}x�)� Ɋ| GGr�<�G�ծ�Lcu�@ ��Ԁ�y�<��A(��3%
^Tg����+�|�<Qd�{]�(��G��y���@d�<	b�ؙh�kP�@� A�S�]�<q! /O�HPK!�,�qQJ]�<� �����D
Xe�s��tLҼ��"O��馆4E��0�1�P�b��i��"Ox���D(�l��ڭL���� "O��ȡ���	I�P��b��3��*�"O��B���9� ����M��]��"Ot�8�^�	��j�J�i�ĉ�"OҌul�l{ pM��*�jMh�"O((�EjV%D� Q �F;_�dqt"OVXd$�t���{��;��Q�d"OJ�0��6Q�X�d�w�ެ�C"O��&fۦW��h*��4|�|�[�"O��& �1�F�k2��#0�2�"O�X��Θ-�0��A��x\A�"O��i����XW��3�aD�B��Yʴ"Obu�WB��L���q�t��"OV��0��'"F��q�6Xl��Ku"O>�PB(�A�0�`b$g.bU�"OHuSBD3%�L:sޒ�Ś�"Oڜ�u-�?jc~(����`6-2D�0�2
�u��M��"֥W� A&i.D�h!ʳ.� ���oI4w_&��&�1D�dp啑>�4��r�9@	�P��$0D��V��aղ�3ׄI"�|Ċg�,D���q�H����UH�1�8-s#=D����
5
�:R&��Y'���:D���ul@%b�z��4�j�e
7D�|:�c����3M,�$ �2D���*m����.Qخ���/D��W��z���ZՃ�_�`	�G�.D�L�1g�2Vx�3a׻7r>�h$�'D��a�ؑ8�N�JpmV+����D'D� ��K�,A��|J%�S�x�>i9T�$D��BS+j�
Ur��R)[���j&�!D�`#�L�|�����>����!D�,(T`ڰ;�yW�Ut,���=D����I�es*��Vm 1�0��P�1D��ȗ�K)����C�v����q�-D�H���2�,���M�pڕ3w"*D�@���!C>��ƸD��MR!-$D�P�FAW����c�"�Vf����N,D�p���*]4)2��?mi|��L*D�����p�r��" R�M�*XB� ;D�H�@���xvN�B�Eʍ$��D�p�9D��T@Ɩu�l!�ƴ!�hyf�7D��x�
#*�q(�,_]VxiE6D��AC�	�lR��d �4t��4D�Lz�`���x���)D�2�p@)1D�4:�K,��h�e,.H{N�v@$D�dJp�W6r���p҇1�r��)"D�����E3!q�e��C�d�:@!��?D�@���2�Nt�5��X�R%)�j<D�Rs�
=/��l���,c����5D�,ɂ����5Y��9F24�k��1D�0�eG�0~�,���
8�Vt��+D�D�6�Ѿ�1�Q��6~cnx+&�.D�8	#��J�򱳦��Gފ���E7D�ذ��ȳ`��t@�Ҙ<@Z89��)D��rר�E���o�7fDP�06�#D��zDh��:E�a@�0
��I��6D��Rw�^�P����2)W�.+�M�5�6D�, ��#<�I[%l_47�\� ��*D�����,Dx��ް=��xjB�'D�<��/�50ݨ��F��,�����`&D� ���?,<H!�*~�ܪ��)D�� `��
;P��ꔌ�#M��r"O���q�%G����2K�76�Zd"OB T&��Qf�9���=z*�X��"OV�G�N��N$Y���2��s"O�QYӊՏ��@B�[-?�|�@5"O��I%�(<�0p���
CT�)�"O���eY�r������	�"3h@�#"O��	��&P01� �X��)b"O�h�/,\`�Aք@|�YC"O: ��E,W���0$�K�$��"O8�"�H22��irEY�W\��3"O����\�b.�U1"��"3����z�![�eHs�`��ôk�Y�ȓlV
9��U8g�V�1j95SH�� 4�l��*�$|���hf��*-ܜ@��XHx���P�P,��FX�ȓ8I�����M�x�Tx��H��W\<���,�r n2xI0��۲B%�]�ȓ!�,����؀v|�P�r���z�4ͅ�&���?���Wŝ�I����ȓ8�X�p QgdlC�@�$|@:��Cz	B��ζK�Ή���D���ȓ��})����2A{�݂2"����4�tsd��XU����3]���ȓ�p�i1+H;�0��  D`z��ȓ,ѤX3w!,eªQi�d�6R�h��̨Q�s��PoF��M�;F���8k��j�D,��X8d�NX�lE�ȓ	��1ѧ��o��Y���� ���ȓi@��Ĥ�D����#	�PS���� er�p���ͺIXpG٩u�RC剓Ci �ir��&n�M����J'�B��;U`xmY��e�Z�!S�Z�B�	t x$���;q��)�d.ϯX��B�Ʌr>6��	� �P���K�&ׄB�	�Z����Ġ�4��%I�Jx�B�	�]��kt�s!���*�~���%D���V	[�>�*���iP9y�B��".D��(6�؟y�]���3n���O,D�D(�� 6c� I�f�!����D+D���sH!J~ 4MK,v��ѠB)D�P�ᅂu�H�"�G�\�NZ$�;D�@�V�����1q�b.eu0��5�9D�|��B,-b69("��.,Y�07�5D��2��Pu�*�B�G�{���go&D�� 5
Y�I4��5W���0D�)�ɍ6�$�0����X�@�j)D��R�O850K$�L�ʶy(c�(D�T(�
�z��΄�z����Ш&D��)��%l��� �_�Ԑ���"D�(��O�:34hRr�T�����6D���`/�g�L��r�H۵�9D���U�J�V:��C�W�3)��0B�;D��!��eD����т48�	1�:D��� ��I8"�SĎ4:9��R�9D�,� ���zb���4�߀%��Yj4
4D�����Ps���9*��#p�8�T�-D�$�E(��iW��B�O�\G��cF�,D�tY!LVm���\+�:�sV�%D�p�`Uh���q�l��z���׫?D�x�b�5�|0�E0��U0%�<D�X�aR4��rs�lv�!3�#=D��2EHI)p�
P)�`Ď}�f�2Sj9D���RM�s���Y�(F�e�Z2@�2D�� *鰵��+���`B�<(�Ȩ�"O��S��F1C�e×3&�"#"O�`�4o�3B���I�.P�&�D!#"O. 9Q�K ��ͳp�ϡQ��{�"OZ��&�H�6�4��k��[
�P�G"O"� �3r`80�)L�6H!"O����\�w� 4�v�ƙO�1��"O�@��)Ҽ|�W�כ2�b"O��{�#8�>�c�i_y�|�Z�"O Qbf3���U	K�'�@�R"O��ɇc�0��=����{Ղ�X�"O��F��a�޽�Fg^!�Ђ"O�yY!��6Q�^�AF�*	��)�"Op�S���=v��mR�>I$|T�6"O�$;���P��):Qwh8@"O���%J�3��X�B��au�8ȅ"Oj�Y㇈�2D��i��R	��e*�"O�y���ѣ#�=r�?? ��"O�"�d�Z��d T0J�8��"Or� 1W ���8
�j�"O8��H�5Q~�pA�����k�"O��#�}ʥ��M�=,���u"O�(Ⰵ�)
���� O;�-
s"Or�֪�8�8�R��m	w"O�`��"ڿ�XQ��&�
�X�"O6}�w �;��κ<?�$��"O
�"��?\	�VŃ�C\�X#"O�M0�i_�1~�qR&%�v�R�"O�@C�F�M�M�"%�<mP�D8�"O��&_\H���T��H�"Oµ�FLЇ"x i@���*<��"O|�����4T?�� �+KcQ"O~Y�G�[-t��e��Ն5���g"O.�0�Ր]��Q�Ї�.e�d(�&"O�-�4-�n|�l*�	-B� 4e"OD��	���� ���P�r�[�"Oݑ� ��(,�ʐ"@�h�T8�b"O�pᥣ�6�HQڣ��}���F"O������b�
�[`̐v�Ш��"Oȥ`aK�������1?��"O
q����6E���y�C��x�F�R"Od�S"Jb�V��CT?����R"O�4I�1N�85B�b��mh�i�G"O��3A^�Z�LP���^�aT���@"O��bP�2`�Q��G�!;ju��"O��f�ha����f֧	�Qh"O��#��Z�.5zƧ�5|^ d��"O�la��D65����B�7LDy�"OF��k��diA�Ģ9�u@"O.؃�MV�N*ء�	<$���"O����E�0Y�~�p��O�/&У"O�a)�A�)|д2�Q\ȼ	�C"O�M1�j�6Y��L�+5��I{5"O,IZ0hȧHN�����1!��۳"O�U��	l��a+�� Z�r�s0"O��ŤN�'��1�U�>��QP�"O\� ���ݨ��X�g�8�$"O�(��׋�jh���S�f��`�"O$���+t� �G$f�l�S"O�q�ț#�f�2`"�$.h(li"O�9!d k�Xs W0!�����"O&4{���o�n�qT��0g~�P�"O��eǁ�4�P���g|ĭ��"O8caD�?F��T�5��5M�� 7"O� *��&j��`��T��M�=M��A�g"O�вs�X0h$���L�;Ό9�7"O�����}��8�cl�����"OV}�`C�b��Ċ�đ�o���z"O"!��.�/&���h��ڠ(�+��O�<9��ʬ�Iق�Ȼ+�����G�<��B�;w��ъ$슻j��}	V��]�<9U��(5V R��:4����E��\�<a���# p�3���Q(��Z�<��DL4��%`Įn�jyഀ�K�<)��r��4���̤O�	�FƋF�<)����hlI�$/C�z����Þ\�<��n(k�TI��(S�q\bEX��Gp�<y �Oc����$M�6�Y ��h�<��Ѷ �:h�gD�p~P�5��N�<qGf�<g F�A�X�:�`�X��L�<�`�� K��aDc�<( ��G�<	��A�mHa;�癣d��p@���C�<	4�@�Kh��D��~\��F�S�<�b��
�HаQMpu�牌L�<	2�^�'E8����)�ư��`�H�<i�'�A�v8�F�;���k�n{�<�E,��4���$&��%5, �"�y�<2�ȄQ-�bE`U�L�,��E�_]�<aSj��5�d�Ł�i]>�uG�q�<1'��� ��U��`1ፂB�<�p�_�K�BQ[֠�e�9��FG�<��B�%]Zd��C©D�ޅ �`�A�<Y3��p�����.[�MJ �,_��C�I���hSj\O�x����0.8�C�	5��J ��-pfY���7.�B�	2!��]:R�^��$��d�)2f�C�ɴy�v����%I���!)�7i!dC�	B+J���Ɣn�@�1�a-&C�I8"PaP.�#.X��$
=*�^B�	�j��1�"bڶjW���ʄR�XB䉯��U����X����]�DB�	��@���Br�((5O�,��C��*_�n�R��`� �����[ZB� gf2T@WKΐ[��T8�́�.�dC��9U�"��0#¼z���MA�h�C�3K��\��q�>���ޞ�$C�=�j�#��*�E���v~ZB�I������BRY����.dC*B䉰:�����O�U��х����.B��+�H�zs!а3.�5���)��C�	�$b�]����(\��袩��y_�C�ɛo����H�uv�s�@�++�.C�I�k.��0"�٤fw��c�靨/�B�.SiB��Ϸv�Ф��h<CA�B䉧!#� 8f�<IE��(���'E�B�	 ��@̀8w���T�R��B�	����'�K F �����jǚB��'<���Н,�0���IҾ'r�B�	�[��V���`u�1�΄lGVB�	3	|%����7P\�0C��<H�.B�I�j.�8g�-<�f5+ǌ#:��C�	Ur��c�2A@>q�'J�v�C�I+G�}�,��y�2٢�(]��C�ɾo�p��AK?X�0튅,�&"[ B�I5]�yТ��Q����! 'k�B�ɰZ'�� 
��d�xx1,R {�bB�I;�\1��	�M����am-K�>B�	�Ь�Bg��/l]��@w&ڗbw
B�)� �%hDL�20�l-�p�Y�*�R:1"Ox��6���D&]1�� �j	HE"O�q4���H��L��*R�3�(i�A"O2u�O"�drJ��]�22�"OfUy
�+4G�M��&�&HȆ��"O�t��j		+� Pa%Y*��͋"O�iq�!C�L,�rPE�
��R�"Or �'�^�<-KW%�2� S�"O�eYpi:��[F��^�څa�"O�l���� ;�uz��"Od=��B�oږ`r�
D#:WH��yr�^7$��iĕO��Ġ�eȬ�yR���Is�� � _�U��͖�y�ᅥP3>ТE�E�(%�-���V��yrT,�X�����7/DĀ�k�y��0.�@D��R&/N��$�$�y��D��"Qk�
�0��@jU%Q�y�K��h�z#	�'\���������y�k�2,�`�@:�l9x4Ş��y���e�T�∬q�x��>�y���7:2ht�ԥ�%e( �2��.D�da��Y6e�H� �I aE�9�R'D��)B�ǧX�F	KF,�,�h�PE�!D�P����MN@���ʄ5g�����F<D� �C�h�H����Q�
V�6D���#+�~��T��Č�j�1��4D��T�ȝe�j��A�Sc*�;t�3D���G�^_zd2�)]"X6�S�5D��!!��(_P��9x�y*�4D�4I��	8>̅�rm�~���J0D��K�#*�~�@���"�~x�%,D��*��r�~xp蝭$�F�O?D�(�c�N>T��gG��a�$��4�=D�ܢ`	KdAP�fC�3�Nd� �6D�<p��O�!���u�@�;��)�6D�tӴ�5~ĻF�Ea~b"+3D����;d.�ʃ\�l܀�"2D���B��7%\�xt�5*-!��*D�t
�K&	Ά%)B��9��H
��5D��9�a�'<ڐA�װP �AzF�(D��� Ϙ��|��b԰;��Q��4D�l���.Z�(0� �,$E�}�'2D��#�*ǽf�v���O��Z�K��:D�ȃe�(�	�L�n�4{�*#D�4*�➀B�J�c ��pa�U#!D��R!�D<}ך	�׏�� �DY�p
;D��:�k�1�D��d�X9�Py��4D��vH��D����X/Y�����3D��B�jĶ(,��GדJ��	���0D��閭� {�0	*�$<��$�,D�؃3��(�(q"D���I�l��&h%D�\��)V�`,9�@N$P�B2�8D�kFe��'�䉲�Qa`W�!�d4O�"g�U�Oe\(jV%�|�!�$�k���ؗI��X>��ʤ%!�D&'h� *W�4ѧE�;!��,���ۗ�/>�4x�DdV�i�!��mF��Ҏ�so��{עB�*�!��D�tY"V*��F�D���5�!򄐐
�v` ��),$$�D�8&�!�4)q�`2�ۗ� #�,�,W�!��w'���	��8y�]�!���N��QB�$�L0��߫v�!�d�;H��5	{L��@�.}Q!�� � �aK� ~�˶����b"O�����/1�EA0\�* @�"O0h��]�$�ʣ�VYd�Y�"O9��@�`�<���lF��Q"Ođ�&�ձ)� �J�'X$/���U"Ovq��E���a��C����x3"Oj,����B.꼺��ԏM��D �"O�(B4�Gܖ\!ϙ��p�ٱ"O�eK%��>1`��-��c*�2�"O4H���W'
�&��e�΃pp�Y�"Ox�r+�bn��GG�7�Fx	�"Ov$O��@Q�8��G �ܱ�`"O�"���c
0���J<�2"OƔ�Ʃ_�J}�#BZ�*�ً�"O�c7K�������ٗ^��1��"O0|�$��;���
%��VЮpha"O��qU'��Y�L�E�F�M��80"O�d���/6�����:6�*�� "O���п:��X��"�/8��P��"O�� ��^�d�	�̍_ ���"OQr���0���Ə(u��	�v"Oz��P�EJ�u�p�	VWPi��"O�bF�LP6��O���-B�"Or����$��tC�F�Z�)R"O1����<h���"�Q�A�PB�"O�l���(m�h���^9���C�"O��I&�����$2�߽��X9�"Ol!�U*$�@�aռ4�.��"O
|#j=<� JC��I��ɧ"O����%�)Q̸Qr� ;sU��QR"O|U�gͺC<\Y�dO�p���@""O��y�"��-`��x�G�3;(�(�"O���3�¼���I���(RC4H�'"O M g��3>3�b�.ٷ�.�k#"O���  R�E��<�G�Y'8�^�%"OhL����]� -�q��2�|�"O�����w�h��#ޒk�,�(T"O^���;=rc�1���c�"Oԣc�yI��S� ���P��՚�y�
W�D�|b�狞t�T,s�BJ'�y�E(2� ����t9x0u�X��y��
D:ܜ�
Qh���4�<�y�˒�v8Yʷ��Vy�1z�c��y2F�yjX#@��cȖ	��L��y��U��*��-λr�(ɘbO	�y�늴AJ��b����	S͌��y�C96H��e��2zP:�92O�y�����A�r��%	�y7@֬�ya�
�]� _�G�4&h��yr��8s�.�	���CF<�(�,��y� �� g�-�R��<!
}@�mA'�yB�U�o�P�@!�0��h��C�
�yr��3x���� 3-����t�W��y��	�$/r�2!h�+2����V��y���:v�� �`��$��i�����y�o����C ��:!@kd�ԑ�yB,�,�x�teH�zn�S���yB�9�ZA���:��Urc�%�y��<�ލI�F�S���Р�"�y��T�M�ir eJ/���G����y2�\�{�.M���ǰ
~�Ё�	�y,5�F�aլ?z h�I�C�y��EC�N	y�c���E�ЀƑ�y�&Ȣp�X��S�[�*,Y���y
� �ѫ#�5A��
���.`Eh�"ǪA����3B�(#-]k�Y��"Oh�����u��H%���!Ӯp81"O*��b��쵠��J�P�"Oތ�7�7fP��̉6�\�!q"O���`�µP��Aq���-/N�Y@"OE��ʷM���ˑ�G�8��E
7"Oإ��Bܮt��(#�ޑ�"O�x)�IJ;ș�a���8�5"O�D{��pJ��a�*O��,+1"OT��"ƕ�`f�t��b@#*M��"O��Vf6B��-
d�.���"O��QsiY�xخd0�d��T�ڃ"O�Ś`Ɔ�9�aJu��8@ `�"O���f�ݛ�#P�&��(�"O�2E�M�4�d� �OW(d"O�,����k�(�K���H��H&"O|=��-ه[��Ap���z�>`�"Oܔ�$��bmtiG	ɸ�M`u"O���W�J�Ѹ �Ùa�Ʌ"OT �B�>���(L�)��Y�"O\dv�Q�<&�b�_v�X+w"O$����rϜ���gY�.��W"O���(�C�p´$�8-����G"O|�r�#�3s�鱀$�%r���S�"O��ͥ;.$�K��P<w�Z�#�"O���@�$D���!�J�U��3"O�t+dG��� ����EtDj�"O�T�P��`Dj�0�$x���q�"O�h:�(�1o�.p!f*�#D��$�w"O.����73널��OȻ�F��q"OXmxE�Z!oO��³�9�lyҖ"Oʤ�$k��e#���!zf���"O���4�.J�� �c��<M�T�"O�D9t�ʪ:d�!��("�Z6"O�11ǎI�ix�p.��a� �"O2���O�8d�
���rpx�"O@M�&���{�D9�,��$��pH6"O�x+'�ɵrQ�@B�D6N�D	A�"O�ykW���n��R�S(zƾ|��"O�M��#u�����,w�<Q"O�p��'��-�9*���"�"O0�1AÚ��i�* 3-@��r"O�D*W&��!
�	@ɝ�pw��ۅ"O�(�6�IXdY�g��\��!"OA[$ ٘��ԣ��N�E�h4h5"O�i�F����3w*�s�h(3�"O�����E�<�E����L��*"Oҩs��� S� z��I��z b"O֝k�,]�H�����,�7�PЉ"OވЕ�!t8�)���ȗK����"OX��`K�i���r��y��t�"O�|"�C<'0�<�d�V<Q�Ne�"O`q�r�
 ���q��@��B"O��r�cԚ
J���\�4b]�"O�5+�,F�<����hS�H��"O�����.FR�I� �o�ޕ��"O��3�i�d����@n�C�2 2�"O꓃M��R���E���"O��YG 	
;�`{楝�Z�0"O���P�m:DX�7P��  S"O��B��Q�'CB>g�@�s"O��H"��	{R@#@TF��"Op��ѠʭZ[�툥/O���H�"O� X��@����$���/0,�	�V"O�p�UG�!y���6�Xh"Ot-��]�%��Q��
�u\���"O��8�c��?J��)D��*��1�$"Ot��b�_�x��@B��A�a "O*�Y�K	��,a�T�3�U(�"Ox�� #9!����{Vnm��"OX;�*gрj,�F`dZ2"OĉHB뇔$SjI�H�O�����"O��b��RY�*�5E��/�LY�"Op�"���d���p3�T2�nȚC"OT�R���e�*D"���(*�*E"O�'$�w���C(W켌"6"Oz��r����@bT�Y�b�A�"O�����CQ��h�)D��1�"OlLy�AܷfV�(37!�<B�"x��"Ol��0
U�u��O]a�0���"O���R���B��1� ƃ]�N�"O��i�-2�� �m��<1��"O������&nɌ`����-k�XE	�"O��9�KI�"dġ�)��A�9b"O@rPh����!�ʥDuF��"Oz�i��]�3�,����ԐOw��0 "O*����ѬP|����!eؐ�V"O6���K[%Kvt�Fn��z|�k0"O��9EΕ�,xpal[���q"O�Y�s���0��8�FB˭	��r"O��H�� $:�H�(U�Eq.�)"�"O����d��P� ��1,3( zQ���s���	�[>�ɢ��'��)�q�J�-�O�<
 ��8! �P �&���"Od���5z����s�)��9rO��d�l�C� �"{&�P�KT�,�!� 4z8T`��5 Y�vҫ	�8݆�U�ʽJ�T������M�މ�ȓa�P�&"^�I(��Ă�Ŗ�ȓ�@��@����B���-1���'��5�$���~$���_���a������	�Z�X#K(6 j�	Cnŵt��B�	%ST�sУÈJiXA�֪H~C䉢* Qr)N2�B�����29��(*	�',H-�QhY�ž���$Յ{�eX
�'��!�l׼Q�p���O�0r�ΐc	�'�p�ӈ�%Ai,mY0� �5]a	�'f�Ye.�q ��w$�"v�I��'n�P�ug�2)�]FM�u���C�'b���=m��6_��p���O2˓�~��$F�T�y�d��ԁA#9����3�ɩ�y�o�?+�ܭ��U4s���N]>��'��' >ի��5�=K��1a��� *LOH�'L�$�O�:�B�� �qw^$i��84��܄㉼XN
�X��A�ZIڴbi͢yW2�>���Iب`���X Kэ^RZИF�+!�䝤-�nd;�I5q���1%�<6��$.}��>%>O ��&������f��9G���'1�	7f���2��&���P�����6mw�y	�������>r(�ug��{�����@�S��`��W��|�DcF�%w����*� �Q�t��P�ȷSl`+��������d��x1���Ҕ=�����!�$O�|3����&β���R�!�d��O.��B���ɂ��y!�R�e@��x�&��z��J��<j!�d�+g=���%�K��5qg��"gi!�� ��e�H�{r1�a�9!d4�"O�qAC���7*���Wc7��Y�"OF�!��H�q�a���0I4��"O�HP��P�g���7��@A2� �"O\a@�c�cD9s���zEh��"O�qh�nI��,�y�ދy9\Zw"O ��!B�*�����/v�@"O^(�w�$k��ě�i�J��1O
�=E��cæN � :�&_3K��SѪ���y,N�,1Ԭ1ը^�+.NuA ���yJ��S��!��E���H�g��>�<���D�1Att����&J��1�f���Kb!�ߦ2�>�CZ9��Y ��_��|��i����gG��s~0 �%C�V!X��I��X�Iܟ,�E^	1z&����ӥ#���s� '����{B�)�	g����CI5���k4c�7>�!�d���#�I0�֝�"G-R�!򤖨7E -�D��(�LDsfB.N�!�سa�bu�*�.�ZQOU�!��_X�� ���{�"t�B��\�!�@1 ��S��E�;�@��O�$;G!��	3�R���EƝ�ԉ���TB�I����;LO���C�S�z��lح8�PiV"Or��Dœ���-��-E�"�R3"O �C^	�(�ċK�M�� K�D����Ӛq������8^�["�ݰ4�>B䉴j��!*��l+�МV�B�I rtI��N����r!�J:��c��D{J|JG��q	2�*b��#H@i1rc8�~��'�FM�0+�u	�l�b��$����'	 	J҈ϗ5��UkR�Jjbz�'Wb&O�qY2)����&T���͋�֘'$r�$!��B(]0��#I�1$L��K#�!���{'��cc�0w�qz��΃�!��R]������hj U���˓X�!�������Cmצ\|ZE2E�ݝLC�J�����7te�1D�B��vB�ɡ'� � �H��_-?�:B�	�B;$��!�@�p�ȄB��G�H?b�d���`����UCN8V�8��Eۚx��C�I=uB%8��|l�d��V<ܪC�I3i@�E�Ւx�v�F� h��C�k>쨨Dd_#|yv0�ᑲ9�C䉀 �H2��L�x!R��M�)�ƨ�`�)��<їd��p4���#��xSh�	�H�y�<Y�N<�ht"ga�P�AB�s~��'N]��?-�̭�ҀѪOJ4I�'��,+eA��Jd�P�)��X\�	�'�ṭ�U�V���;AΘ~�f̫듸�=>=Z4�N$$�2(("+�%�C�ɩob|h[�)E(a� t�&E>�|C�	9Fv���L<U�q�V��C�>������B�==Pp{���?gZ؄F{���ʓ�~"�'�v�hN�iNp�@Ϟ]�Ε�rO�ubr��uy�!��j��,���
���;�S�Iٖ/�8����fn�-JъE�a~�^�(��B5W!L��� xO�� �1ғ�p<�!�ۺ.�|<q�ʙB���6	�U�<����*Q�I��ᙙ (UCW�B˦Yz�,�(�����3NcX���
�46�����'��)F��-3J��#j_�YŮX`�	5$�T�uCC�2�j�T/ǔb��¤�.�R�R�񄇓��@bE�O�})q�lɊ0j!��]�Bk0q��
�9�^��Q+"p!�� �`� 3k҄��G_�����"O�|P׋٫B����c%\'io��;'"O���)9r�#��D5?n��{�Z����T�'�Xq2Ԍ5*��$��18h���'T�l;�d]�`f��ZE�W&.^�y�O��=E�TnM�G+t��$[��0�!����'�~ ���������Y�O�3S���+B���y��Or�"~b�(R�	ì)K�m���!0t�WG�<�d���8���an��;���F��<�ϓ� �p�U�^���*йNO����	�<��(y̜#F�ӥ'�r�BT鐰��x"�־f�q�B@�BtBkt͍���On���iԘ	��С�cI�N��Qy��ܟT�1Oh�=�O����A���A�*?�j��E^��!��b� t9���^�m�C&��2�!��"L˞|�#��5wP��Ґ���(�� Y�8*7�1o$���W(��il��'���iy|�^��C"�:}����Dk�);�L,D�L�m�7pexE�E��>t+��)D�ܚw爢 %���!i24d;%�3D��Y�JL;g�uhq�ug|�F��<��5�ڤi����4i!�;Nz���s�'�����H
�j��As�#�����'/v`��*+Ql���e/����'�����G����D�)d��'h���E��6�ͪW@ۆ%@�š�"O���fμn]fq�Aώ1P�d��"O�ԙ���D����2-c$1J�"O��H"���WY�/]�:sz ��"O��*E�<g{��I��ӿnm�b%"Op�Ǜ�XP��u��2rT�@��"OB�hMU
����J˕e_(U��"O��³�
�c��,xf(R�Ub3�"OF-�H:h�8)�@�L?8Ha�"O��ŏʰ#�dŚ�B��1�,��3"O� +�c:]�� 5]�"��\��"O(<i4�F��f@��@�V�<pc"O�ZA�-`��d*IfSjԺE"O,����5�L!W���Z8 �!�d�D0t�Y�D�hp���W<)�!�[�q(R��C��'Hc����#C�!��w�p��)I�7��I� _�w�!��_4n�l� `\�p��Tk��c�!��ٓ0n���焠K���D�7*�!�D�g�(�F �"6i4��gfܶP!�$Jx@t�� O5\b@���J�!k!�$ tm����(^� �<1q��?Oj!�䇴G'�u�$LR�i�B*a�Cy!�D�
�pLR���@�$�+��ξdv!���7Cr��Zv�R�#���8���8Y!�$^�+��1�F��e�`1��"�:�!��j��𡋊�Sj�`3q'C�>7!�$��(���M�m?H�2Q�Q0{ !�Εs).5��&F�I&�J�k_�q�!��͚1V��_�};�h;��1D�!�D�iȼ$�)ׅ$
��QkE%F�!�ִ ��d�򏋫V�nP�֧ø!�!�U�6�ŠCY)_�u�'�%�!�B=�Zm!χ�O������fy!�DB�#�0��qI�>�������J^!��0� ��]�	�s��AE!��L�\d�hj���X�Dd��.�fP�X��H%Qa~2��
�ׇ,���z�E��y��Da����CN�&�֌Z�� �y
� �m�fjԻ[�H�6i֒3�*�z�"O�E2%,H,z�d�x�q�F���"O �4Ԣ{������V)�.e�"O�kBi[Kh���.[>W^� �7"Onq�D	5�`�0s̀<P6�M�"OZ��b�.v1�� ��E�j��3�"O
����Y�?�\̓U�vVL%Y#"O�[��%ԦγmLF}�Ԉ0D������<�#� �r��a/D�D�e%Ә*��p��ř��y �%1D�����f�D�w�V�>ﶉ��.D��+�a1:�!�"�U�X�U�6N-D�D�o�7hp��Ff�
\ق)ؔ�+T�H:��\X_ư��m�x��Q��"O���+�ТB؜�B�[�"O�ȈQ&�����ЛIW��B"O��R���|C^��տY@.}1�"O��9'�&o~ BtfߛGjl��"Olu@R
�V���(������V��^��y#�'	��zCh�ZN5X��D)`�bq��@��6�D��	�F�rv�ә=��b7%Q?�Rlp��ˡ��	����O���)g�;(���'�蝈������Yg/W����"��~�L��gbʐF"T�Ū?��$�a	��^It╠\�"�J�����`@oՐE&�	h�'/�D��	E�e�h�)&��	�qF{҉K$�>yZa�*i���;f��ɄB�x�ʗcجXc���k\�B$d��}8�Dإ_��� ��L>1���;�J!PR��!	�pQRP[���h�c�O��Da,N�@s��(�\�XWAQ%G�P,����:=,�P��	'u2�� z�����Yb�ȁ�	�w��Ș��4�t	c1WܔDPw)L��y#h�|±M�v����!@�4�n);�Q���"6\�z$
�jR*R-lO����)I��!��@�.�h(pG[�	�t�t��K���A��� {��p� &J��%�$i1h���Ol�D�>�TBO"'��u�P1j�L��`�P;!�2-bR��A�	; �81"���_>5��hս��+bHS�?���A��v�1���b�Rx��%��o�iР Gߟ49�Ʌ�oQH�ӄp�)��Ǔb��e|� ��e��n{bK�%0��Y�ǌ�zV�4�񡇳#��% �CYa{�,������0iŌ����q����0�B�)�S�b��-�<�t2A�ï���D�bH���$Iż5�*Ih���}����cS�&�N��/��T-��o]J9"y��)��mD �l�//�8Y� �F� A�����Y����B��e?�N*sJ�w���49��i�:XS6Y`l��	!�pGH�[��`���^1̀�����s�t����ʔ_�1���(�0'�G���TϘ�eGBLсJ�?.��$���F�(|��)�����ҩ�Ry҅�&7Sp�zS'@b�@��$XdhR��OPv�F��)�Ш������%�oN��b! �XS���,Pt �DK��1B`�4���w�p$�E�2wք�ۇ�¸I|�ثQnBW&+�->x4�����z4�e�2vԀ�ӗ��Ky�̃��C�`T�5)Ȓ�2) �1SpHu���F�[��Qp��%~9s��ն[�l�dɑ�*p�bV1Rq哴6�`4R�kL;o�$%�5�Q�6h`y3Ǣv�ʠ��k ]= 3f55�n(n�v�t}"4�¢ l�Ъ��݌JD�)�"��e�V�����;L����ٳ. �
��x�acՌKE�s�Hh��D�Q;>5,֎�|����2 y�F/�3o&|� x�0$@�4m����"���L�wk3#i��I2l't�x�˗�L\6�U�A!+�Ji;%߁.f5�%8R`�'�T��D�K�Z�9�H�-WМe�' ��d�a��1tF��T�U�"��p�e��
& ;��^NHFQy��J5\\x�1�C�rK��$��ֺ�bM�O| �p֋M&��dC�L�@CSE/�Ms���%1�`���Țmc�L�u!P-�Pzɇ�?����KX�:aaH�0�ʐ�ei�0=)�X%G59�k���]�R��B\T]jx�SA�����U2;"�%u�����T�QNc��Qd��85Т/ |i�d�GsT: � -�8��G�Hh��	��@$  �����~
U�d*"o"v�yqE��R�p�	�6��=�B�OVQjp߂U�� 3J�b��O��8s��lH����>���`���`:p\h�`U� �.����[� |�:�#G�d
B�1�
B?���X Ǜ#e6f|8@���tl��
���W�<_y8�k���L�z��0���&b9�A� ͜�!����I_)�P2 L�!�8P뷏]�4�*fĔ Ŕ�92+ô~�ҝ+��Q/gKV�Y���$�"`�Ϝ�:�z�'A�̓D�֔�8	���+f���1D&�>A�)�wrR%�'� 0
�Q��+��R���0ׇ�2fu�4B# �榱��E
��Ի��&Afi��!�{�F���h˾��Pr� �6\ �-���iуZ�vu�'v��P��XH^(uKC*�+jxx�A�@[�ɜ=�4%S�2�R�¶�W�r��a,X�LT<Y�j�)mvd�)W�ۍ1��ec���"~�V�j�-F�L׌�)K>a�m� MԊ�9c);ғK۶%�����T���2sC_6*���4Ȍ�+���*39�u��k�+I���P�HV����^�,�����荂,�|� k���Ũ��� ��q!IF����E~��<1�q�N	L8,p��M��Z솔2AU�D?^�KY&�u&��qCN���j��+Ƶp�Đ XaH�"G�(
�<8B<�\<
 �PbL��Pb�g���(˵�߇T�0ii�	C$��ǲ]��] �%]f�Fm�C��u:����&N\�qHF씧8A Xx' �	��y�nѭN�ı�&�4i�0���) ��M��)T:s���Ɇm�3<	u("Z�P�s7��hтiS!��Q��%��)�V�4�0�R��ޑ& �E�!�� >�j�"����c;�DU�Ҏ��	��9*��\�"?���nՄ-�:���J]�#���)�c̼ �TIВ>�!�D�U���b |I��Z �'K��zp�5��أ�D�0/��2�a�3x0�EK�?�N���	�-�&aj1._�B��7�(�2">	��ڥN(��/Z�F���X(~�6�b-����!*�&E�^
�R�j��[�����O��������Or���A�v�b��@'-8^� �'A���ԫ|<e���ǹ8bpA1��N9N��|���)������@'u�$HZ�G9?:��'��A��n��Ϙ'8�5a�̑xm���Ø�,m#փ�5����J-Cz4��!j����A<��1�i�tHK�"��yqB���+�����Pg`C;E��G�D�>��{B�yq�IA�n���t�L$�Bq(���W�
� `�6"�*|y�T� 
�Uq��P���2[��3�u��X�ZH(�(�.R�W���E1��On-��B�L=N��#�U��Qq����Du�K�S�"��cI#0���1��P似E
��8��$:�n?1�eE�Q�D��Q����	�I�����G�>�t��N'��D��:T�	0�|}.ٻ$� &B�H�qC[<ܑGǓ?ND" �% ��I��F�?Y�8�5_���I��'mP���Eȡ_i��:Ȝ� ���̚��$Q<\01V�"y����m_.\�eJ��f�������ٲ��إS9V$�̣z���XA�^�]�����8(68A��t�~�@�ܺ*j:$���C�0=�SΝ1��X���BN�Yr"I��M��Np��xd$\� -�L�H�{���(WI��AH��];0n����0�]B���3H�;Wjl�熊��'hd�3���	� ���Idb\(9����	Z!B�zr�Ũ4N�0F��.A~�J-�N�r��_�e;JȲ��cR�����M�������h/�l"ٴ����*�ViI!��,^F��̌6M��FA�D@/ZHl=�o��8��*0jTK�.3��ܣG�I
LG��!����/�r�cQ"$���Ȅ�YA*8��G</t%)"/ڈHO��L>!2oZ�IL����fL/v�ů� H�j�t���f����Z�T�Z0����N��� �M,q�9CE��I�z)��a�)c�([����Or0�M�2#�m���W�b���D'����ɯa�aE	�D4�uh6���L�x�*&��p��EA�'c�*١Qb�
��4m���&�T��83H��aT�"���S�*�N�뮎��x8%�H�p�\�Rդ_�mnB��d/�X�rl���dӘ��m	1�����V�I�t���
	>2�Иx3�_^?�G��-QE���#ޖ �<�����(AGXXz��ȻX2�EYp	�ڄ2$d�����C�*MpB�T����4B^�?hQ�
�5е ~qR�P����%ȕ ���M��n�E12!a0��Q#c�9{�2�ґD�!���;e(@�R��&�!#f6M�tn\�V���4|a�t$'*�ĝ��*0?��hA�Œ�w�L��!��!@���M$Ru��C�����m�������T
%G	�S����A��"tѠ�ͧT~��k�-M�
�-!���+D
�ig�
&6���������}�b�0?	�CÚ$)N����#6��d�d���s7.�!��Ը+nVWi,d�b�L%5D��bݖ0�\q�f"W�+i�\Js�K�[.�AY�Եi-�&�'1N�0���|�(������a���#j����k�2"�yp�J� ���J?�	��ә��A´�N#k����S�i=.h�v���dU��a����wa4��Ї�38EF��ቘ4=3|AwƓ���'c���@(Op��`���§�!��@`#�5tnDy �f��/{@�h2ឌ;|+O��H�䂼|<�v���N�7a��n$������h3B<��lD�{�xR��p���`�G�JŢR*H1|Xup�Ñ9��88q�U�/�� ���4H<�۴! �µeU `〉 ��%yRMY@���@" s=j�ґ�Ĩ��u ��6E�a�!�F�n�c�UA��d�\8"� �/@��۳��HA
p1K^  �2��8=<<٤����`�?���CLH%�'�>L�qߠG�@ �</3��p���O�%�䏶p쳲C^��,d�Yvyx"�ڀ��t��@6��r��9e��׈VgzT:���*���F��j3r�`e�ǥB�����	(��@�e����-肇^\��ի�"ۊ"T|0�(r�Y��X�+��P�eF0��	�g~���Ҁ">��� �¤�.Ų %G�e��|2������I�lX��Ӭ��xx�#�-[�7m�����88ʸQ�GG�Ш9Q��O�o]����%|q�kqm4h��8"������ҔF�|-R�٫0ܬ�0B��oܓnTb	'&�l��$Jd+�U�J���EG�qbv�i�Ӕ(V�ِ���F�:�ATF[�w�<A�r%�XUit��O��a�O�҈��b��,2����;tBR�~6d�����	�@��M:�Oƍǖ�s"�=G�-,01���`�
�9�-�!v�֝ɺ�u�H ���8T��78Lu%YЀ$)��M�AR�����R��@�U��|2t�ʘ
22X05k���!ci�KϺ���n�Y�"P4����D�ʣ)^�-ѶN@�5'�9CI������ؓo�yS�1�襉�gT�d�wT�Th��ۚk}�xů֡|�p��E�Bٶ����!�	!l��X�� T0��m��IߛT��d)`FҊx�Zy�-�$O��)��� b(���ʔ6��}�ԩ_�Q��XA���~�&��A898�����e����a�b��#��D{r�&gG�tc�&'n��Ĉ�ܞ1� d@�U�QL(���+R=Fl��Ysȃ#�L�iE�SN�0�3d�~�Vʏ+#��|�ٟ�*�A���8YP�R=$�����P�IS8(��d�Z�T`ܺ1,qh��@e�+I9�!�'|`����ø+X�p �ō)�|a��[-t&��R�XАr�m������/J*(�"���m���!� ���`F9 G �8���gOS/T0�qQ��uh�[��	�|�&զ��0��G��u�Kן2=���U�_�GXu�@冏K�n�a	^�����Yx���KV�hO2d ���o��U����%z�X�Ă�g����7-��a`�F�BF8pXF�l��]���݅ r�a�R��ۆy��_�<�V/�!��"�&C6�d#>9�D�E�䙨CDS�S!��P�Զ�x�8E惈K~���Ό|TMa��Vl"��$[�����O�D�Rc!��?���h7F�?��YC��ܓՖ�����n;��CG�|��A�o9��k�ܴn�1�0m�>�p�&[�<q�FN"�=X�(�2����B�c���yRoрQ��� �.�,�H��Ξ!�)HՈ3ɸ���胏g���m�-	����C�x��ؠ�O�E����� ϩ;��W��	���,�.�Q��}�������F�⥉2���D��LзCB9gͼ!�g��ul�oZ��b``g�5A�� {g.L�w���� ��� t�q!�I�dCZX��m�P��}RA�[�����I�9Ԓ�x,ݧ~�u)O�|k�c����b3� .���)v�P�6���4E����X��O�b�b<H�#G3Ƞe�UHT�-�0vͅ��Mj4�L�@���a�1�X��a�$@���c$� >J�=�Q=��yrtO�<@��t�2�V��1�AU.s�@�5 T%�'#O���� �� �8�P�#pdԃH�6������!��t���GcB8t�������ysT���.�#{=4�;��xa駇*�(<���C;q���ࠖ{v^���N��y8��ۄCp�$��+%'����Đ5ڪa����L�V�Z��:DaP�M�HPʄ�D)!+�͠��1ӸA�j�Z�1�%�=6�)X�K�/��͛e�͑2ZV��1�� A����"*��[�b�Ġr�?_���w�ȾW�P!Q�������ޏyG��{��#u �k���(������I=P�H	2��?����x�� �Rɚ?ҙ�vJ�3���0/����p󤍰.��ɋ���
o��]�࣏=�����-�K���P�J��n��E��К ΋�1���`���|��q����<+��U�V��G�OjM�W�!/i,�<�`;r���P&��ɚ
����C��+@�?���pd��xF�P�1,ȇclT��3��@n��lܵ7������ײk��L�57�V`��R{x%(OQ>�ᰲ�(z�E�kK�y�#űN�D01� sRxݺ��Y�c5L<�����t(	B��,iN�%1vC�2H�n��g�ƅ{����j=hZA�A�]BpqN��
\)��"���'����J1g��R��S5��IXtaJ.T���|J��nځ@��
%�R��4��/���(��r�IH�{Ϯ!��*B+"��ePᬐ���'(�
uRd��q0�ԆSM����y�y���	�1���@1.Xn s���Lq�CZ�)�8�F3E?xE��^0*�V� Ë�HR�|�iؼ�y2�1��)��E����7n�1(�R���IW�\A`�?x��%���D.Jl`���z �GD�j���PĂ$�O:��֠�-t�7���s�4������i
�t�0G�;w�$�����l �$��F	pp.�cW����.�Rf6����Z�ko�}0*��3�a~���X��j��׸-dD9J���/�I�G�Q�`��b�աc�Ȱ�.Z|pu�@�V:)lH-b�L .�����Ă�oïE(\���` ?���@4�X�y�5(�:��8�cG;X�Χ-�`��B�2�F��!�8PV���ƍ<%�pa�(E��Se`T꺋���-m�$��%�Z' !8@*��������-+�4!HAS�_z�I ��6�4����8ˀ�Įk�M�፝�Q0,3��/\h��BJQ��e	�\Ip��D���fPy�ő�,�D�h?)��*.�hL�E)�/'0PyJ���W9�����F]��]�eP�9�f�VN���©ŀ���D mϪs��C�� �Dْ���z�+�%�0�����+M�q`/.u�&mY�oC����>����	[�oV�c��{��l�?q,U?XF�ݺF�9��сf8-�R���H�{FI�1w9`�4W��qÛt�>�zf�?�=a��@�o����ǉ�l�Ғ�J���t��{�OCy���q�%ǂcW��"e�0�j9�e�,` &%N��p?iR�؃������]'n�I(�._�'~����@�.w� H�)[�S�VX!��ǥ8�`R� 7[��B�I8�H�����o�y1b��=����*(�`p���!b�ի駈�Hq��/S/7@(�bP��<I�%*3D�T���qߐ`�G�ڵJ]>Q�auy�a�%h� a�倆���	�)lrXH� W��@I��G�h������z��ѱ�Xs�,���85(�g�N:9�(��'��a+�NϠk4l��s�����ƭaD<9���įݨp����n!�*���@��y��W�N�x�Ț:r=�D��� �yB$P�u�^����it���N�6�yB��b����%
oAHt�N��y�K���TzǬ;e�b��e���y��0�P�$ΐ	YI�MA�Ζ�y�%{bV��R��&̪̔&��y2���TV�i�&��*�WJ˳�y"߰fU��_[�8Ƭ�
�y�=+E�]0�߬[D���	��y/޿Q��(���J�m��D��y��M7|���JA�FI��#v/6�y�E�E=��3.J�6v�B6�Q��y���;r�=@+�|�8�
 /�5�yREI��̰9�ʏ?g�8ݒ��3�yR�::�T�"��*^����$ �ye���6*��Ie8y�D����y�`�-(&t����A��)����;�yBfQ!1q�KƭD�q�>���@��y�B&EV�a&�S��#�K�y���A؀�p%�-C}
�ȇ.W��y�I�L��$8,@)<h���E��y*�4]a�t�wl�X�^� ����yBr��ѧO\Դ�6�y
� P�3�7kZ4�z��U1$zP���"O�8G��2tc�9`��� ^h��"O:�3�<zn$A��+aKb���"O�Uà\���YД/��Z>^i)t"O	s�gҡ� �"VLܥ3?|q�"O���KD1z��;�L
;Ij�S"O�}���-mV�sa-��x���e"OZ�X�쟶W�j�6�ڪ.�"��U"O��˷C��H[��G%ؘ�e�"O�G���'�\]2"�ŰoA�<x3"O��`�ҒvIR�+�Jܑ?���"O�Œ�J�����ɄS�p���"OF-��DW(O��� iP#ir:�T"OX͋�S�@4�
b	ٽK��#P"O$�[VA��`�:Q"\�(�ԤB�"O96�ʁr�V�7��g͢�xw"O�q�%fd��� ����v]�U��"O0���R�;�������w���j"O�B�n�m��c}��D��"O��#�Փ,�hL�"�weT��"OȲ�h,w<���K]���P�"O<�� ��O.f�Y�m�N}�%Ҷ"OP�x��	8h$��0��;ή(����f�j
ç�j13CZ�^��c���h��	A��326�����\�؅ǘ�	�N�cڟp��`9����>�fY�O��E�EJ������'�J1Js��,)�[5�[,`�� Y�%I�|;�h�6:LhT]!!�0-��W-xJd3@�D@�K�mz���'�6�Ilܧ)t�z'�R�WB��c]�	[p�D{�"� ��ţ$bՑl���pG�].�)U�.HB�
q�НjX	K(\y+��0!5��D(Q�@@z��L>���X K�	�2g(3a+�9�6�ؠJ��b�)0f�䐡g o^�F���X! W�y����0����j�C~FA1噥o3\�0���p��Q���(L��W����B�Ȕp�* ��rӂ��Q��,0�X瓁)J��`�m����*C�U؟t�_dM���q#F�!�݁k.�O��#��=�ؗW�&B\� M� 9SZ]��-;!b]B�BE'����T\2,���▤+����8R�'K)�(��6+/pl��ރL�R,+a&Q�s�n�OP$1�Q	w�zE�rFK��	�*3e�i�)9^�K�*䰴��'.IܬZ1�D?v�z�D��*'�Q�B4�\�[ǎG+簰�J�4  \|ě6˖7[%�b��ANpHb�F?l�~Y��/�^$9d@�E���ug��$J���P�پ%�t���@�e�_���S2`�
&�P�<:�ω��'h��	�������cb�`궎��U��1��)�)X60Y`�oWc�O�|%�v�i�����7^����L$�QГ P���@�vbP��o"��i�´���އ8��@e�=(�4p��EE��a�kF5]�.���k5teVyt�i�p|�eB�.�&\SG�D���Z.E�M�5oT![2��`H� �#ª �Y�V5�E������+ �v��WnM<8ڇH��mɆ�
�I�����w�M\.�1���ڗ�,YSv�H�}̨�Ebق�u�1,��a����7'�Y%��q���&}���pQ���<5.TyA��]�`��E(ɗg:��S�T�L}�W�[��`I�Ú�5,PqQ�\�j���i�p�@��8�\5a1��@�6�1�mN�Qaك���^�Cdm�7��p�=�D��:B�2��O>dJ7��W#�,(q��/pJ�*�c�'v6H�[ebJ n(�R�$ޡ38xrGCd݉�R ������M� ���KR.��1W�!��C-����%> ��5�]�0����P��C*��J.t�h`ѢH;wW�`)C���&'T:1�A�8�F��#%˖3�R���$�0���8]�DQ��D�?Q*i1:�H��c��6�ƥ�0Lˢp�*�Y�M�>��a���ɤ0"��<��%�t"08��(�:
mP|��|y�%����ZbՈ^_�9H�H�P,�#��̯$�T��]$�9 �,�0G�i�H��Zwd	��{.-S�ʌ�(﮴��X3�M�7�i�X�QFE��(S+���<J�L�dY�})��0'�t8ð!a�N%xS��7/�Ɣ��aЍQ���I')� 2�.U���ͻ�0uIq�� (��+��GD=Tq�F�d���F��Gh�h��YѲ��ӟ��Q��~���f��/��If)B>L݈����l��e�rېd�(�K�쁾J�V�1㉆�c�����r����?�dC�0R�b`"T��f�3?)D���g��Zg�����E������q\�b���.-"t TH��y\�(qGE+s	���R�F����agĈyH�j���>�m���ܣU.�������Y�È���5��I:D`���ϡ@{����F��s�t��'�?	�iJ�皯_k��׬�;{L<���k�%v�тU&ټu�`���$S=����,��H&���`Ȍ���H��	Ez-�YxK焳b���[�M wݒ �ش,]V<6 �֑��A
3�rE�b�d
�i�Q`��-��8Mty�釁so�\�b�4��t"G#<����"�����jL��M{���QD�k B�^5F�1s�ŌCr6`��87(��U#T�5�\�P���Bh��PŃ�DJ��5�N�4�2�OH����/5�6I#���V�@Wp؁�'�=��	���z9�rh,��	C�8���W�D_`ġ��7��q�B�k�5O�@A��:@ ��O#(=Jl@��K��p=�㨊�� �©ՕC
�$�ХZ@L�)���F@aAT�Ͳ_�]���3�"EX��TG�0��e��CK�='�� �HqQ�N�E��	�S�ܞod�I���6|��`�G�!D���1�70߮�Q��J�`�%ÂnѢz �*�.�����9�H�.�9�w��+ 늄ȡ�'ޞ�x�ޡ.��9�*ݧ
;���4M�T��7�J����!3�1Q����B_*89C��:Np:S�[�Nhg��c�i!�䃀m��۳"O@5��!i�4��K�U�-��oԣi�P
�f,i���%Y3Z�D=�����!k�$��J�]�1��?�,qЊQ�4{�����;S>qqW�'R:}Q����I�Al�$^�-�G��Ỉ*��ǂL��	�E�t����<>Ȇ��NR�H[b#>)���L�-��gY�A�0)�,#����I"m�
Ȓ�G�W����ͅ�?���L���7��� �PjP�����~{3�C;c����>�~��ī �Cd`��4.h���W�˘OX4���7F�c_�3�r�+��c�䆾Wdb��g����l�@���KhHٲ�E������:X�~ex�,+Z�}I�����*X�7�5�`%�h[�$vls��^?GDȨs(3S���``B'|Op9+�h[�	��D�7/�'ZK�����L�_B����ȵ��d��$ܾN��̓�E�(
��P���;�/*1����)���9*%J��`�L/}"��E��ईhb�77q�����iB����E�)9�Ex��M�6������,_\���t��p"C�Y��T���'�&�Cņ�z�P�ҟ����#m�����>�$��V�y�O�K=�!����"2��$ZwHN�3����#_ [�bO q�,�7*��CJl4ң*�e�z @!�|�����#?�,P�놂 �$�'*=ғ2*<�$d>5OBh�U&H���z3!1KI�3C���\j�#�H+0 ,�t�Q�7JHh�%&	� ���C1 *�xJ�`�*��	y��@+YI��XbB% ����'�T8	!œ	C�<�g�[�bR�F�ůdC6�p���uݨ-P�f�klL�
��C�D�,�#M���{! ���M[ڴE�&�0!�:y�2dj��1;,�`�d#�$�1:(�h�'����wjB%@3J(ۃa�0B,�X�(	�^,4F���3��5r�2J9Z&��J4�:�Xtg�W�d�����*��- �)R�n7M�)`+-Ѵወ  B�d@�m|����i�0h)�D��$��QMNU�L02r�IN�bb�����q�,;	p��&h�~F��G��7�n���A׿m�t �w�Dzn�m����~��N>���v�Ib�X{�q1�D�n4�M�-��#�Bm�E'\�>X��F�^݂�9�o_s�YP��8o?�eQA�"�@E*g�6-1��lì��9��B��tL�r@ѳ��� L�<8�e��d��q�e��6&>^��NC�9����m���X@v�P=ii��oڼ;Z�I��B��L���:zz(��#�Z�((뮂2��e�Ξ�J�� ���A9gxU����k�6B 3Z4�
g�n�� ��+'
(�E �*v8���o��mQ���(WBmKP����x�d�@� �
�P���yA(�6]Fr�q�� *QI�V  =(ő&ˉ5���	�FwAMK�=̀���,2j5+'��м�s�L要���.a�����'s8�a�ʐ�[c2�rfHO�]"eɕE6��E��	�/18h�ՂД_\�ioZ�)��(Q���N�R�⛟dI��K�	�|�x�E(�9�A#L��� ��-S��x�2ϐ�m�	��d�)
h��J5�+�5���X�L���@FˬQ��`�2o*d��� ��2oM��ۢ�I��j�@	��I�?d*EL��ֽ36�sSz,�s��SĠ��b9������ʍ�
`����&J�=����lK�>�J+b��#�OȤ��D�?O �p�+^`�����l����,���r� Q���~Cx��ɬZ�0� a��Wp���$�m���ݴ"`�sr-�=$h �j�C�j��M �Y; �t�î"3h��Ξv����]�Ȩ���{�	�B��ŀ����!bg���.�,�y��َL���i1�Y#s�8��k�C��F�)Xpŗ�8�$9#�$��e]����`�/&�t@��	�O(HA�E+O���q�"�X��Ŏ>+��H�T�_�juh�b_�n��ē �H�˵�ֆu/��-SzHAA�Q*w�����<�8��Ӓf9��:G�S^�lMEC5#<R�!�dP���%0���3Q�G�$�|(2LƔD"RyX�R��{J�m��1�5���1� [�E�A���L�@%XuH�'R	��C�j����DP$+9��1C�K�W���Cw�\�r�I��c	6�8(�.]=p��IgK&.2��aӀ� U����s�Y�#ٱ<W�XSf��Z�H7�V�c�=�刄0g�P��`ʹq�n�2�V/���A
 ��r�C�ޢ-P��*k
|q� �8*8$����V.��fA��A>���b����+%���|��J�o��Qn�4�O�}8��)�d�?�Z)jP	H"N�𰕠��8����!�	҈8��j��_���K�91�؀�#M���5�Ϙ<����q#I���*8Ƣh� `�J�8����Շ7�f��q��C~��� f�K��pdI��(�*��G�\a�h���S���0��;-��Yqv� �:1h��:����g�j�˟ԉ��]_٪0�u��x����7NCȝ� EG/]YȜJ�i��Xؖ�H81����
�U�d�p)M�l������\���)�����B��#'V5]Â��Ɇ%>�dL�/<whE�U�On@�q`�CÎ�5\���#�i�$�DS�/�bd5%^:��V�Y�*�����T$Eҥ#Y�h ���ϓ�.��$A��_9��f Y�8��2I6r.j�	���)T.fq. �Z��7q*f�1�'�(W)hmڴ��F�u��$�uξ�KQ)G(��c����ӈ����I��l���Ѻ!�I��m��;�4�1IG���K��5Ӗȸ7S?��-��:��uA�,ـ:��1�Lʳ>��e�s��W�']<�`�"|��R��7z�8�`�AЩ\��a%��;U��+�aC��%��Q���k�%ܾg$�'Pw��§m��+����L;������[��	 r)X%Gj�'�0"�!N5J0����JM_��%@�i!A`����ze�y"Ý�e��PiĆ�P������";ʹFI��El��%��=������OP�:�-�*b����-�ta���Pb���'o 6��]�B�]\�(uF
x�|0�.�ri���� ��W�-V���a�(9zj�Z�l�W�RHS4N��[���s/@�`�EHķC�Ҁ��ŉ��hOL$����L��D�RM�#��=h�$��-g����)�|�	2��1AF0�r�8O��L���&���'0:����+Ϋd�I���9�j��Q�[X��Rf�I#H|���DG�,w4bt�qK\�$��%A3��SꙈ��G�l���bIߐ5s�8{%���>``4��)�~���Y��F�q�#7J��	�tg��-�Dy�$ɺ((Z��c�r�()^��5�3Hr,\����E���B	^8z�	%�� "I����e}"uP0�W`;�����(�6�V�rI8��Z-*Q�+�d~(m���f0�����RŦ����%tN��X3�\�qt����S��@z���4���S�AF�l�H� �(M$wF����]8rt��ƎD�T��4*���7��P�����h`�Ł��uF��Ɯ��AЏJq� ���[e�O
=��ȉ*�2���dC�J� �a������B̟,!텋^h��ψ	����*VPh�OZdi�C��%x��3�ӻ1@��oݕ?i�Yx "�+��'�(00�+UZ�ЭI�N�|��i3O�j
4����[�$4�&_��8ٰ��Ӽ58���j��i��r>ᛰ !X�"4����7�,Ř֠ܞ+�i����murըE&�#�剘��ɉգ�l�LK� E\z�m�78�f�j����i��t)� S�y �2�4\r��X�y�/�w8IQlB�`U6��%� U�
i��0�>HZ�e�Z6�G�v�p��Q�
L�Iw��p�n�2��_`��Dېv�tTg�/p�f���E�#D�Q��ǔt�|�rG�˰>�܀W�&��S6LE:x���+A�y&�pB�>a�@��K�?���<!'˱;�Ԝ+RJ+2>��  N�r��Ke�̺ ��Y�"����;��^�T��K��^,="��� =q�����:'�^���i�*x����.ڕW�n͑��D?[���׍1�	?Z���w퐌O�i�I��L ^�E闝a0~,� ȃ6R�"�RF�/&�r�6C��*\K�M�)%b>�J��`1r ��H4W�>�Jƣ���ǘ�a�l�qM!�2���ʭ�~Bˍ3o�pGIY8Zp!���2|�д	��P�s��e��e��;���Go,j<�q��S*�p4�Cf�5{������f�4�:0�;gY��(��9��kQ}�!���YS8I�j�0>� ]����#@���еe��1���SKP�~��!*�*Ɏ]Y.-!c:�l퐒�@��H c6a&~"�V���m�J�8t�5�s�� $F�/Xd��	3=�<���G�$��EC�R�W�d)�'=�8i�i�.�J%i�8�*���eǟ&���I����@j³y��9���E�E�̭#�ß��$��k%A��b��� ��-�̽7(���5�0XN;0ƿ���j�A��  ��D�Xz��n-u�HI��=h�M��"��+*PKء�2�I$h/�(�qÆ7��=Z�(¿n�A���O),D(��"�(� fصL{rDӸ`�8;�̖�O��E��;��?I���8.�j�լE�]^��·� M$��/��_�P��Ee�/x1��r��+�z%��̅>XV��gc���P� �p�r9ځ�Q�0^���MB���c��A.��b�B�0j���!�$j.]�E���*T(�#�c��{"��FҴ\d��¥C�5`���aSH*�'��Mٴ�8�����O;pQ����Y�+���J��A 4����	�.K�)bN�`�4oFVb�u8u�L�Om �dIH�t�1�晅Ulܐ��>)�Dǁ��TX�Kc7\�:��B?1w&B�]��8�a�W|HJ?I)6ů�pP䆂Z��X��W7+$�e�+?�Ɖ�� �mz��D��p��}��m�7m���a�D=0�,g�O��<ej@O�5
�ҵR&a��sQȤ�c�F$��H�;&�u� �S�`�r�S(>����bD���Gԓ+�� ����� ���WyJ%��*I�:�5��NM�1���q�甒)���}ΓQ	&xU�T�z��xEg��4\�GB��-Rj콊g�U]�S-)���0�ڗf����G	�d0�����i"TӲ,U=���wF{£U�VXޤY�<$	�y�Ԩ��I�yJ��"�ԟ��X �T��ޝ�%,�(+r@ r�vcđ�7V�[ʼ��'�O$� �M��b�P�C��(�d0�퉮H6�t�o�3�툇��4� h�#)T���3w-�y�*��/.�0P�, �f�C�,�?�¢��<j���18���)�/i�yJ� ڀtAʥIGŅ
(@:(*�'���b���
j�a�FNߔ���C�X��J�	[�VXT�GO1Fx��A�x�D�P����e8VX�gi\�p?7�Q���%���-%j�� W9p������N��C��${��,�aj�9Bz�Z�	��6MF�?	�h�,��b?�r�.\����J�9Y���3�4T����D�D�֔�[�}ބ��"O$p�,t9�`7�	X$��"O��"��ʙ��!G�eM��A�"O���f'���!BE��A"��"O���ҧZ�h��l���!6
�C�"O��RS,O�&8Q����*DQR"O��Q&�[�Ew�����3$ �!�'�����)3>A��IK(2X��'�����+�;p^8���A�n�,@�'2 ]₋�D�@B��Ρ�2i��'��������@eH^&	�>��'�u顧G�ZE��6�di�'�~�q��<e㞙s�NΥ C�|��'Y�-��&Q�+�>��ҋw[ q��'��,���ūGr=p��A�78� r�'_ �(�E[�`��ds���\��I��'�N�2��Q2	�N�� ���`�|2�'�	rs �����H�ilPQ��'�v�iB�a��9#�׼_/��R��� F٠u�X7�X(����@1"OE���,�nak�E��q~�#�"O�h�!R�
~��PVc�PP�8�"O�y�Phέv+�呀25M��"O�����Ux������6P{"O5�����X�T�L�z��p�g� �Q�1�ɵID�@��؍�~r��,�A����nJa�0!K�0��7�!�d�,����	6L����R��$ ��Q󏍎#SO\	Z��_��M�ᓸr�C,M!
�<e��S����4�*8���f�pOQ>%�l�]@<�ḟ�G��"(�䘏�(O���Xd'�����B�֤ۆMq�\��`����h�q�|�-8Ց �A�{<�R�e
��M���E':����Sⓔ�e�;b�R���C�C�lM8���=�z}�I
�����+{���ç ���[W��,B4��D֕@fH�"I>�y2d�Jb�Ij>["? �䐤&�:��8��S��b�Ik��C9>���$>���ǘoox�rD��gN`�`'cX0�~���G��?q�$��v3�х�Ӫ\���!M�q�w�EE������j?:��Z�y\YK1�ؕ�`��_��m1��(�����=?�r$Y�/Q* �%C/��41�X#Z3J�;�� ,�5r��OՒA⟹o��h���}��LR�0�\)��Գ#�ȩ�%C:Z�&Q#�UBXH93�'3���Z�[>Y���c�0c㖰^�d,��ڥ-8�J317l�uk�"OI���	�[��[��7%Mh%�L��L���9��J;u�x[¤�����۟Q�֝8�*��a+ <(��s��,@.��'�T"�'/���	��1.��겠@��z�3N�5/��~2G�H�)�'O��I E�`t�I�*��=2�	�~�+�V�i�@��Sp��X"ŉ�
���|��A��i�:�A6?��'e~Z`�FF<mpD�@+�%R]��n�t���'�Jq���O_��gE(8������S�F뼥�免q~���'\����7��ɴN�ڴ0�'LK�3�����O��ض�Y��M3s�J���>�"#��eVT��V2l~� BoS�ovHl��f�R\Q`�˹vӦ�8�ď#@�X���Є�S؊H�ve�pO\Q_B<�ȓL]� `Ջ�::�h,8�J�x�b���:U>P��o��|��ȡ�u��@�ȓ5 ��ׂ��+N�ԃ���K���� ���iV�γe���!V-׸����ȓu
�L���$Dr�@�a�R�"I�܇ȓ�ܬ��/�'\��\*��7wj8��/@)�vG�R\�8��l�1������a$��3rx�v.D>����ȓr��;s��0]:�D�7��zdt���Zb�tۄ�ʺK(Ke�,ZlC�dQpͪc�EP�d������s"O��!K�f���J����f�1�"O�$�٪KԔ�Q���#�Jh��"OtآE��	�dtX�ζSyl�"Oh�P�׀@���y�+U�~�+�"O�=�P�ۄqK�m#�ݿ[���D"O|��uA� ɮ�9`�4.���$"O�t�҂R6Q���eة
�9#7"O4��΅�.Z��B
�M""O`A+���o>,1IDa�Q���W"On\p��)(L,4��	��1���"O<Y0�.#RX��j)Ht ���"O����M�T�B%Ѕ/��*��|#�"O0�`�	I���c:)�	�>Xspm���0d�ղTy�|JG��e��-��MJX���s�ǨE��q�,^�yb��.=�RyKb�^9+�$��K+�y��J=w.8����%J,@ڰ"ŏ�y�F�;-�n�ʐ'�M$�e�Z�yr�J`H�@���|��bý�yb��20���Llk��P5�	��y��O$���2Kb$����3�y
� ��iT�D@�럨=���"OzXCda�.aƔ8d)�Ezl�@"OV��wE�����È�am��"O�#���>��k�슩+E��s1"O���m��2�n��s�K�!�p"O�ࢱDMQ�����AK�1���z�"O�q�+؏X�V Җ&L!`�2lJw"O�0�sOaq��q�0rBE�"O�����Q��ځ�#�|f�ɕ"Oz�W��'#����*;I �s�"O�p�"f�~	�i�uյJVl��"Oqp2�7akj��I��m�x�c�"O�ib�$)bK�2�B�Q�0�`�"O���<� Ā�w��H0"O
�Б!��O��(�r�$%� �!�"OJQ����#���@���1�R�R�"O*#� �W�D +�C�|���2"OFI� 9^�x5Ʉ�	veN��1"O��`ͅwz�١ǚ�,[�0"OF囔�0���С�_�I<�0D"O�uؐ �%`�V�#���!'N�!"O��$��(���s�H18t�CU"O2��$��Xe�L����*!R�k�"O`��ٞ��mc%�^���"Oh���I�(4b"�fU�L�R�"Oʭ��&�eBT����h=40y�"O��!�'���A�#%����"Of���K��҄�WE.�8��"O��J�e^�@���7�.���!"O ��i�X�A�$�	\��z�"OZ��B��C�xH�bDT�X�@�X�"O��K�2H��PgË52{���t"O�`����*GuL�H�+�zy��"O�Z�N��D��(GH�xi�L� "O�)���ŧ`��`�eL>yU��{W"O��+D�u��R#���#�UkC"O5���M�~,�� �O�x R�"Od�R��l�*��#��}��d"O�@C`k§'�I�桀��r۴"O�THe`Ј,1������C�T�[�"ObT�@˞-,gR�x���Di�"OL�`b+��2�MZ'c�-^�B��C"O�tm=VD��L�	���"O����q�l�@K�:H�p(;�"Ob��J٘
�J%5,���R"O|�[��m�$����Z�"Y"O�9�	�G"8�֦\���"O�Q	g�A*e<����2�vu0"Oک���ʸP��uA���N����"O�)c"G�l���a�=xu�X�"O�,8rM�����%��D��"O!T��0D{0\�%G{�N�15"OT����Љ�6�K����J�"O(�jn�!��y��IڒQX#"Ox�n
Xi���AbZŚ�Ip"O���M��c_fTi��J�R���j�"O0<	�L��:��M��i��e�lLx"Ov�B�@�#�A!����T� "O���E�܃>6���	�� s"On)�B�p�<�
�(Ђ���"O|�9��8H�H&�4� ���"O� ߫�(%$G�_�d�B���N!�J))Һ`����"�&�"�OE�[7!�Dɻ��c�"��VÕN�j!!�� ���E��;��0��]�D��I��"OnD�O�0t�|����ؘ(#"Ov|*��[(��\Ñ�+�n��"O9H�n�B�Н�և
,A(�!�"O�ɪ��I���;ֆ̔5,ȑ�R"O,\1Wȅ�~�4x)uEޯq�IG"O~ #�
�yhИZ�.äU��I�ȓf�� 5��J~�S&��VTH���Yޮ(kp��iG01i��LU: ��:�v����.4ː��bc�*)�ʀ��|�)��O�R5PdQQ��#Ofe��:��P���h�1���!K[���ȓjϲY%�A�g�$� �,$� i�ȓ8cJ���Hҟ�j`Eᆔ?��`��}�Z�e��W�u��ᛑ+�%��5z����I^�2T��#��M�Fۆ�ȓ{�<i@eX,p؀�)b)�G|����c�L���e�o�e�"��?wxp�ȓ�����S�=g��l�P��H:"O*)�!ɉ2h���+O2�p���"O�JQ�)�k��-��i�5"Ofu[@��.T~e���m��x�2"OdMKC-B�P��1�Č�*S�h��"O��c� �a�l�3�Οp#l�Z�"O(l��͆,-�P�ڑ�\�\4#S"O���dJ����ST��`�(��"OvMP���2=�
,ȥ̅c���"O2]��gڽ~%X��(�+*��R"O�a�"�	�U�w�eN-��"O�%(��J�e��<�̍C]N�{�"ON(i�����p��K�!�0��"O�Ը�f��(R4b�
�;]��:w"O��K�K9�h�P�H.��|��"OFt ��ZRJ������*�<4"�"Ovi:QD
�3�ܴ)�CЯȠ�Y�"Ot}��^;�P�Iu�<T��|K�"O��LX*��E��I�e�l}P�"O�-���0s*�J��4y�<xY"O����/�M ��	v��F� �XU"O�w�OO���YQ���:�h�"O�kUoєrN�K'�Dg�]�"On���?�*ɀ�i��ShK�<Y��WK���@!5� I��KC�<Y1��>�r\e��a� 9�fD~�<iGZ?6W���U��h��k��y�<�AeB�:M�sb�=l<�c�x�<�ShG��B�$X�;Aw�<)����/��eB��΃����Tp�<y۝s��̊ zG�Xa��B�<AE䎂k�e�fCQ�����&�B�<S�A�U�$Ҧ��HzHz��w�<ylE39��)w钵�	RS��I�<&��8R'�x1U�bD�ia�H�<���Z�8���b�%� <^�Y�BA�Y�<�%"���r�Ȣf\�{�(L��G�Q�<q7HP�FI�p3UMO�K���d�<YqM�	�^Lkj�'Z�xK'�x�<�fNR�O#����)��Et�$C0��r�<��+k@�H���O�:kؙ ��Zl�<A�,��W����.��B�`��j�<aF��4>�PRecĚvμ��ц]c�<A�-v8d���\=��ș%�Pk�<)�N[�m�،	"�W�]�&��a-f�<9EI�%gP(�ɍ��yD+�J�<� ~��d�E�y+7�ȟ=T��x�"Ox�Z ��1�n(#S�MR@�"O�9�3D��#��@`�i
��K""O�m���պq�Z�
�mȗ}�i��"O$��UP�[� d9R'��-�|yH�"Ol�s�*ٚ~���f�!�i�4"O�����X�Q�I�$
�"O�<p�n��pni"1jG�O��]�@"Ol0�ǀ+&��=0b�T��ed���y"��F8(4�3��59�,u����y
_
t�@���8�� :a*Ź�y2&��]���b� y㤄�sE�y2➂m8e�X7`!C��
�y��ƽ��`�D�	"b��	c��yb��$��Yô��l��!Ó�� �y�I�=G�H�c��^��̀����y"J��'��(�fآ\V�<B���y�j�0a4�uJB�}z4iQ�̱�y�7j��\� ��w��������y�ǎp2h�`�#P"r"5�¡N��y"	U8�Ra녓6R�l�r,��y�o[=L;¬y�$YZ�pܡ�bX��y�
�4LD<�C��5Y���cn�H�<I���!�"H9�.�y+>iz�	^w�<���W�T�C���%5`�e�J�<yF�O�W��� ��"A?0)�0BAC�<�Γ�=N�!�2�B�؋FlIE�<��D��t��eGK�t9iP��v�<���D�_)���%K�b����)�s�<y&*� m�!�D�Y8�rYs�<y��U�0g�|��x���R�G�y�<��_�N\�T�%BS�{��(�!B�r�<�IL9W��D[����B��f�<aG�É?�N�w얺psjy���_�<�P�
�B�J����ó�����]�<Q�`   ��     �  d  �  �+  �6  nB  �M  �W  `  l  �v  �|  .�  ��    �  G�  ��  ˨  �  U�  ��  ��  8�  {�  ��   �  ��  ��  �  ��  � � �  �/ l9 @ \F �L �M  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�	�� R��g� �t��B��1�s�Ee� "<E��'�����?l�i�|����y2�6�Şw}��̞�� `�d�ǁ���a����dE�D��p�i^�;>��S��%+�|�L3}2jN,m��+�lRu��iT�y���>�����Q�g�عQ� ��Mˌ��%��|ph�9IV��1�!�;qu��UA؞X$�>�XR��V�ԎPԜa�g��:]&���d(8a�МA��řcYx�h�G��%ڧ\�ƠB�!3]��`��G�44��^�Ȅ�-J�S�d�Ӱ%�'
<�'Bў��$��Fa�,ʕ0�i�9j.!�$�!i�;��@�f�I�Iſ+� �牰D�-�Dk�;�Q���c�C�	;<�4Qd �
����'�4��'��Bm_�K;�HاA�H5���|�����Hȸ-&�tbr�Žp#��v�/�yb(Ͱ6��9�L��o�(��^��~�!�S�Oaƙ�gh�[8|`c��e��e�'% �;?ʡ��� J���
�'��s0i�3y�Bd˖��Vy~9�	�'�F��A�^_8@�D_�M}F��'����7�[�Y��:C��JF���'�*ex��N�d�B��9;� b�''��SѪԮ4	�#"K��7cL�8�'����d �el�0J�g#����'�HS��Q��*�р�	����'a�|@0l�9�0�p�A|�`<��'/x2���93�]���:%���`�'W��P��҈4�����)뎨2�'R2K����y(J�0�D�Z"m��'�~���j�$)ԡIg�0����G��O����^�E�� �9rdx05$?��{rɚ��I�m#��Q��Lm��$*Ǹu��ʉyr�'q�x��H��t��ѯ���r�H0ND$��=�3U����"��M�霂���.�69���ȓAR�L��/�B��ǭ��-����=���?Q��Ӟ6 ʝ)��^�%x"T�&��~�<Y���7?=f` ���4~D|9qM{�<����J�Fa@o�`Ѡ�sS�Q�<�[y|�d[� r:���`n�EB�`�'F�|�ڮe��)҅��F��b�O���	^���O(���b�>�bI����O��p�	�'eF�Js��#y��L�Ǆ�U�
yK�}�x�鉷4��9{�ɐkL����N4Z�rB�IlZ6�+l�	<�ؽ���Pdֵ����'] �cV�`����jG�%��9�'jX-���_�"�ba던�Da	�'�bY��R&��l�� ���$��˓�(O��5,��N�R$�7/T�j�~�J#"O�BS�]9af�K��G�Y;b�s���=lO�A��ydVEk��ה:0��"Oȑd<$�X���$Υ|����"O���t.R9ǎM�1���S
nj`"O�:AJ���,������eh�ha�"O\�!��שn=Ҍ��$�	'�<Y
�"O��#@E�U��C��W�9���"O�؀�J��}:5��k
:�P��"O�D�G@فE5ZA�Cj`D����7O���df��	Y0i؀}�~��)I�5,�,���'���ɉi����AE\���z�&I����5�I�|9������?& �S &�T|�B�	���0p#� ��� �<}��B�I�Jz��5B�% dY��T�A�6�F������ ��A��ƛRTV�BpH�>���6"OL�ke�I�Z t�A��V)(��2dU�p���h��Q#w��
T�� s!�F�H�ZC�I,A:� Iv�CQ��2�iħX+`B�8P��(��_�!�l�s�H�3
R>B�I�T=dX�!��N�ZAz���._B�	,$��rVk[	l��-q-�)
B�I�e|Lru���Z%��� $��>r�C�	0����ThW]jP��-B�6Z��#��c%O�>�ȉ0�F.`�����4�O��$�QԅƪuJ�AK����>���0ƈ3D���� 	F��AƂ�5�a �M2扃5���?�|b���b�c��$��iIGhd�<�0�� T�4+	I����a�`�'O�yB	Q�$�� ��>;L@�cc/_1�y��%&�&aYF.đ-�E �Ј�y�C���v�Pg:��P�7J<�y�n 'Ǻӑ%�0�؍qbC��y�ώ?~�Pt,(t������	�?����v\8���,�H�Pu��!i|���ȓ@��-Ӥ@+n�P�Sd݃B�v,	��O�����!3��q9�(��D���fcҖ^����)"?��,�;�2%��۷�����(�f�<���H��z�eZ�j�
1I�<��l����v����¡К3^lm��	�!n��M{�O��e�k�!�"��"bN؜�"O$Iǣ�W�$�����w���S��D�O��s�{����P=j��1���{�|x{V�D˟̄U24�K4�ҔT�X��CDP�(��:g(I�&�ݱ*�������>�rԇ�,�*I�K�J��f�3��!�ȓ%�M�adT/J�������n4�ȓ�Jt�0o�zB]��j�b���^=�P������[Ôpc���ȓSܐ�bɇ,�����ODN�ȓ&��MJ�� m=j�%)F@�م� �]Y�Fѫp'T�C��J�[@�ȓ?�,�B&@�����1FTl��b3�Y��N��z�	d�.n�B�ȓ9����[��䪧(Ų!xPl�ȓI�@��Q�(]�r�I�Z<��O6�dұk������@�]�(��׈��H $��<1ѧԗk����n�hU�ݢh"69YŨ�<�\�ȓ[�p�Q��L�r��a��_p&ȇȓq_Mb�o˗%�@$�+�# �����<_p�+3
�h�F@�3$����@ua���7���9�'A.S�\�ȓ:����<%�.��P)��(����|��6�Ѯ#���ޠg��=�ȓ-�E�� '��ߓ4�� �ȓ"cr�@�0!{�	�fΈ�
@�T�ȓu+�,J�$��P	�)+vN6Utz��0܅�P/ٮr�\��v!�h��x�ȓ^��`�$5)x,�N8�f�ȓz� 8��O�]1l�RT"�39���ȓ{/������-��$~(�ȓi<ش!ĭ�_<"c/ק!а�ȓi�Y�&T�w�^��n�%4P��ȓ*�f�K�JB�$
��R�ĩ�ȓx?�W� ❩3 �.��\��`�Y Th.���)˯vD�ȓM��R��+�:v�Փ"6E�ȓz #U�$ut�A��7-�4q��S�? ���*E��t��Ś���(&"O�"&H�8��U��e)���u"OnQ�A��r<x�D+^�@:8�W"O�h��&Y���k��N+/���"Ob�p����U ro[�[Ά�[��'��'��'��'&R�'�R�'Ӡ���J<OT���ʗ/p�4���'���'t��'�"�'A"�'�"�'�4�Q*J�$BLc񧆈aR��!��'�"�'HR�'��'42�' b�'���D��'�� �1�u�3�'��'���'���'���'���'h�v��k��<"#��>2\�E�$�'���'���'vB�'R�'E��'�Dm٣��"D*����Y�r<�f�'���'���'>r�'���'��'&����
���`}�&�ȐF.Jp��'/��'���'e�'1��'��'"�����5`�P� �R�F�RC�'Z��'{B�'>��'ub�'�r�'@����k5c@�A�*�-5������'���'�r�'e��'or�'���'��)�ը���e��Ȓ?'�=�F�'�B�'�2�'#B�'7��'���'_dQWhV gg�0S�M��˂�'���'%��'��'Q��'"�'���AЂ��t��!�,�W�'{��'�B�'���'���'+��'u�� coK==�vlz���f�R�*s�'���'��'���'R�a�����O�Ձ��	{����rrgjm(*O��D�<�|�'*7�Z�-	�&z����g�8�Y8W��D9�4�����'�	�"�� 5_OՒ8S�	|���'��U;f�i��I�|��OO�A�&�ۧ�U=��d�aM�?�6i�<�����D?ڧ��;"n��d��PE�,T�+�i����y��i�ʦ��4uu�i�����Kt)۱��
}gJM���Γ���I�k�\6Mm����&���@Ad�p�t��q�q�PΓE�Hx�����'���`��\�#�l%@��Y�F>rU�'��	n�$�M� HKZ�2�i�Ǭ�?�B �B��}*�2�>��M����y�R���V��ctK�����0�GH>?A��Ǩ�I�PO̧ƪ��P��?�gM�i�J���ì��q{�D�+OP��?E��'l�����R�\$�U�g���Dl�c�'�D7��7C��ɽ�M���O몬��.�j��m)'N��-�'���'�R+�>�f���ϧb���"�#e�ɴj�:"��
�.��^�z�%������'��'�r�' ��;����"�cg&�"{T�i�Q��3�44�ݳ*O�d7���O8"�)�f��dAb
1VH�U���D}B�kӠo�1���|�'�ZT��CY|١��C�~0��/�J�9ї%$��ҿp*<y���t�Oʓh��مϋ�!�x�b�H���񉒎M�����?aPB�9S?�-ၩ�3H�0�5�?���i9�OV��''�6�_��50�4���Y'� wh� �gjފ�^��Ğ
�M��'�b�Ӝ *$������?�\c��|;��� y�ڈ�Ai���`ј']b�'�"�'�B�'��OKra�	�
����G4�l�-�Q��'��nӀ�2:����O��O=*R�O?'�ে�8�8�i����O�xlڶ�M��'L�xݴ�yb�'�͸����w0Z|�F�b�uq��øG��z'�E�m�rP���i����?����?yCP? ��K�/G&⌈uI�!�?����?���_�ၣ?�?1��?��i(�TM�q״��I�o �f�)�yr�T.��|·6O���b�0m�;m���|���U� ���Mdld"��,PVX؈Tɞ�4F�TP�U~��O@���+��'�d��\K��u8��V�ʩ��'�B�'�����O�剠�M{� �c}�M*GB�9T;�U�ڄ?`+��?���i��OH��'��6�� /���DY)l�`�#���+T�l��M5c��M��'���$�@]��&<D�	Y<P��q	�2oN��$"�,���	oy��'4"�'�B�'��R>1ZuK����T,�2-��$zSˎ1�M�$�Ӛ�?y���?QL~r�	���w	
M`��G#T�� fJ�0�h�,p���l���|Z�������M�;g��M1RL�(6�����$S�u���'��r�
�O�[M>y*OT�$�O��21f�W0��T	̙t�-#�D�O(�D�O����<�i�1�T�'�b�'g���vHژ2ȠD��r*�2�'��'��֛&�`Ӡ}'���A�'Y:k������Rmz���ɠFi*5�A6+�8��'������T� �'� �W�݀g)�����T��j�'�D�eZ�Fa���� š�O<�oZ�\1<%�I,j޴���y'�U2j�r�@�ؚ[R�j�ѿ�y2�w�o��MWo��Mۘ'D�A��W����5j`�p�5�Q.p���O�T�
@�ג|�Y�����d�	�l�Iş�Jpm=Z�FM��aW$����@k{y��|�xz���O����O�ʧ�?A��)���#��yJA�ͅ.���殮�ش��9�I矼����+��p�Mb�F�2�)х����R��x!�	�u�u���'�B�%�d�'�h��6�I�>���;e�PVd�4#�N��FL޸b��߱2�A"ᦂ�E�h���FbBJj����(�O��l�M�i��a!Q�{�|����0��A3�(XYr��3OR���=F�Y��3�0˓�bU���  %!��G8*mhl�cd�4sn�J8OzB��6#��8�5��i:�i���O�3�|ʓ�?�Բi��M�ΟJme�	�ƅ��Q�vx�Tb����I<�#�i��7-��Pq��g�������$\IZ��Q+J�/N\��,�z����4�'��0&���'���'4B�'\`�[#��#���Ѡ# b�����'��^��
ߴ_^Z����?�����	A9L[���6�ۤ.l�YiӤձK��������	�4x����O�� X�� �.@���1�����I�$��ӓ傓?P���?Y �'P�@$�8 F�C�Έ��'X�l��m��EA��Iǟ��	ן�����	yyB�f��Yk�����;�뚙+��2�n��d��$�O��0�d�O�˓e����9.Bܣޝ[�f������qv�6�Ȧ����QΓ e�q! "�|���	�?�S�o�H8�nO�(�f�QH�d�7-Y�����O��d�O\�d�O��D�|��p��$�%U%���)Dd�@��igL����'gB�'��Of2!q��J�0<p�[dҎ}-~ 
DU�M:`to��M���x���Đ/�V?O��	�g�Pn���5A��[!D�v3O&	AĦި�?I]��'�����T�	=_'�1��Q�l��UA�fDll��'���'qrS��[�4g����+Ov�$�*Q�qFo�'V��Q�T+<?\��ЩOm�*�MF�xB�ց�H��dK�c�J�j��y��'�� 6F�
� �QU�<�S�>b�Fşp���_mQт��[�d�"�K'DϟL�I�<���D���'~�U�C�W:�pj��8��'7T6��<<oD�$�O�n�ϟ�&��(msh)�^��*�#T�P�X�:�M�@�i��6m]<rհ7mo�d��*3F�#��Omh�S4�L,5� \8�F�QE
�!Jl�Cy��ѬxÛ�:�͈-�B�� B��j9,����<�� ɉ�r�%�A��gn 9��=D��&�MsöiD�O�����IǬk��-����~4���A �73�t�#�ԢNR˓[xĨ��o�ֱ��&�	Δ�qR#J5 ����k���Fݜd?:���G�����*�2e@���6"@�BeP�1O�G�Z���ІPW�K��H)�|0�T,�(ކx�3ɉ�jÀD���Y�,�9�O��3���r�-K��M;�_�:�����QîY�a�;�J��\q��PR2 �q�u:�̍��tx��M./(<�,R�	���Z�ʊ��\0��E����C˂�/����aK4�,0)q��D9`��#N4*���J�S�x�T�Տ5&�Ā�eO'ސ�(b� v\���E�	?Y��kڴ	E�Ю�pg�����|�B�JC�M�	ş�&�H�Iş���!�>Q$�
;M�(h(d>)���]o}"�'���'��I�$o mM|����(p�q תډT��P�q��2G���'��Z�<�IğLq�� ��8��ݙS�2^2��B+�'k�ߴ�?1���DΠE�>�%>u���?�؏k�V|s���i����/	�7�<A���?����ş�?Y��ae���4A�US��K'&	��u��_,�E�i�P�'�?1��%��� �nU�4�3���e�B7��O��DZ27p��|���&� � �߽�&�	I�bX�=��ArӀ9�����I֟`�	�?!�L<ͧ,�>]���R�KK�`�S86Ҵp���igt]�gY����ş@�3�	ϟ����ng�*�Xڱc�]3�p�۴�?���?�,�Z}����'�b�[*T����S"	�]\@�j�!����?������<���?a��U�X �뙎`h� ��SY��s��i�2.���6O�I�O��Ĵ<	��Ka�x��ꖓ=	����CUt��6�'���x�y��'�R�'R�:ߢ��4چ4�>��&[�wT�����?9��?�(OV���O���w��M�yy���q���!NT2^1O����O��<b��8%�󉁀[7fT�#��$z�
3c�-!���ݟ$��؟�'v��'6������)�/�B|����k�i �\���I�d�Iyyr��/w��i���4��%��E@)S%v��l����	q�Fyb����O&,ҲHG�*�pu��,ك`�Q�ݴ�?�����ܲ5�d%>-���?�أ
��T���
�8S��D-p7�<���?A��^�'�?y��e���4	F����Z�����&yӼ˓O���i=�맢?9�'eR�I�W�S��;��p�F��6m�OP�N,�S���ē@0�PϘ:�@ L��N+�1m��Xz�I�4�?Y���?��'Gꉧ�4��!�Izm-W~����,E�6]&@L���?9����<q���Ω�tʜ�X?JMP���eȚ���?���?���T鉧�$�'*��Ԯfޒ1�BȘ37P��.����?���&��a�<����?��'��eX�`ҹO�8�Y�M H^q��O�Y��<���?1����'Ɔ����|h���m�z:���Ob�����d���\��ty��')tDk�lQ�k>N�e���Q��̛
#���ן��	�8�?	���z�@�����-C�K�t$,ixi��d�'���'�I��#j�s���qTJɠ6i�(1P5��ܦ���蟨�	a���?���$�x	nڊvW��Y2�ŦgΠ�1F\����?a������O�y�,�|���)�j��B¢G_�4���@P�d9�p�iW����O�$:s. �|��'��[$K�{�tu����$�
�۴�?i)O��$ڦ$���'�?����ڷ�E$3��%��3�����Ί�D�>���x����c�M�S�Ĵ<�@���t�4Ś����'I��T3)���'���'+�$X��=� �)@5� ���eŘ+
�ڑB�Q� �	6Բ�!a+�)�n�v]���D�J۔L{�j�$��7M�%5��d�ON�$�O��i�<�'�?���P[�]��n9D�����+1՛��ڕo�&وy����O�mq���'-��*��H	:r	h�o������|yd�5|��i>�	ȟ���m�t�Pn�& ��ip�O_$�`Y a󤓟rꞤ'>U�I����rȠ����R���r�H�dIo����8##�ty��'�B�'�qO0L3�m�,�2��F�Od0�]���NY�j�,��?�����$�O�db���	"4�2�k�$���d��.<����?��?1�R�'e���DG�\2PZ�d�v@5�R,ֻY���OX�$�O,��?�f.W��d�߃)����HM!S�:�X�KD!�M3���?!����'����!z�d�4ZFP9Cĩܱf��Q��Ԛ	9,��'���'��I꟔�	�B���'��- ��{6����&N�yBv���nm�R��$�	꟔*�ǝ%G�O*����M����%���B�tb���'��	��\ j�w���'�r�O�zͰиKB��SEȠ*�v���*�	ly���O��isLY���U8-> �LC%ZZ�	ޟ�[�B@ڟ`������	�?ᕧu7ɺr���f��*�̹p�"���ķ<�#�y��ħO<Xc��=Db�1�J �7���l��'����I��,��ݟH��Yy�O2���~���P%^��=ð�E�Nv,�Ox�Ex����'�~,+P�V��L!c����� �s���D�O|������|���?	�'7L�3˂=66�A�4�Ӄ,+�	<Hp(L|Z��?A�'Θ��#+n;�a��cHI��@��O@�0�/�<����?	����'��0k@0z�D�!K�>��	�O�!i�M�&��������Vy2�'L*�K�D��?q� )s�����)�J*]������4�?q�r��hc�Ϥ�@��D%/�M���
I)A�'qr�'��Iҟx��JLR"�J>+�
��p�GGp�tZ e��u����p�	[���?A�L�.tj�lZ,δ�A��Mk����đ.J��?)���d�O"���I�|:�'!�a���EԖ�Y��C�?�~<�ܴ�?1�B�'�N �W�V1��]c�p+u�O��0C��B�~ H�m�ߟ(�'���91E�ӟD���?Q᦮A�b�J�e�̶a�*�!����'u�IV6�t4ъy���$*eT�Fb���˟�X�Z�
'Y�0��+���������	�X��{yZw����"��+t�ur+��ҫO*�]Iz��;��i��^�B��b����0QFFS�����Zd�'�R�'��TW����D����_,��[!C�j�z1�����M`O�� Ԛ��<E�d�'�~�P�*�X�P�����l_��7�h���$�O����#y���|���?��'�n`@�K\�� T�pæ9�ɱ8��8I|����?9�'�U ���J�I26o�)Y$� ܴ�?�X��,OH���O��d2�I�&
-��C�&�d@F�@&\��;�ti7��M~��'B�Z�P���>��P��N�<��8q���s�T�Є�Nqyr�'J��'��O����zp��1C�"Ԩ���ᎷG^�8�aF�l��	֟d�I]yR�'�LHk�ҟN���Nh^��5! q�T�t�i�B�'�"���O�u$b2,C����>+	8�sS�z|�h��#���D�O���<���:�0��)���d�z� �x��7!\8(��y&	mZ؟��?�bR>�W��Q�If�����;1���`� 0j6M�OF��?q6'K���	�<��';���	K�,�,C�K>B������O���Wˁ�S�1O��9�`aS%WC�����f��3���?I@Ö��?���?����B)O�n�*zb.q�5��
��	;�~��	�,�G�� j>c�b?IkU�� <���"D�dIV-��{Ӵ���O���O�D矨��|��-�|)"F���Bua�1C�����i2����M������$��QH���G�P⺑Y�\7_,,oݟ��	��@٤�EEy�O��'����-oT�k5Ø$/L2��F��<OD��<ɦ.8C��Oq��'���"H�I�'�U�Tb��2F�"g��	����'��'q��D�&:�ۢ��N�|�R�N[���I�> ��l*?���?�)O����W��˰���#v�<�		��ȵ��(�<����?)����'�bL�6}楪j�/�� ògX
��j ������O �ĺ<���U��X�OpI@�hE���ۂ�#"���2޴�?!���?�"�',ht�%ǣ�M��Q�	�>��GNό)�� ҃�l}�'(�Z�0�ɓ���O=R(�}()r��ȭ&$luG�@�%*<7m�O����I��lK"�#�d0�4�@�ǉQ����,T蛶�'V��ޟp�*�L���'~B�O"�1y�����-h��޼7�F� ��<�I韤HC,5T��c��']�����43�l�*���U���'�2�?���'K��'��t[���$w�����}����$/Ui8��?���ڮV��<�~���R�}��u��՟
��p�sN���q@�
�M;���?����Q�t�'�� �Zؼ6%ޗe���Aר�5�6��]����Z����櫛�A.&�bՁoL|���i���'@rL�oɒ�����O��)� <��de�2yR�B�J
眑��i�2_��B��v��?	��?�dŎ�uP��g��?245)԰>6�f�'#�u�c��>�+O����<���[AB#hc��J�1M@���Q}bKG��yr�'2�'��'&剶��2��,M��؀@�ܙ۾lI���yk�����O�ʓ�?����?A���5<m�a�Fx�ڴ�$Y�-&��<����?����dRL8ʹ̧q�:���Q\6z���~�L�lZay��'|�	����ޟđa~���Ƃt��hC1
�@n�p�T��MK���?9��?�,O�t��`���'ҽ���W6fV�����c8J92�t�����<���?��bJl�' �$�K���f��2ZF9�gH�F6���'�rQ� O�4����O�����T,�!Ck�F�u��H��X*��t}"�'�"�'��c�Oh˓�����b|X���/'w�y�C���Mk.Ol�1σȦ=�I�\���?��O��I�@K��3S�:
����C����'gB���y2P����Dܧ~��ըW���+���l��A�m� �h��޴�?���?��'���ny�F.Yʲ�A#*�1
�.8�W��]w~6͑�-�=�$9��ӟ���Ǘ'��
�9&�+���M{��?9��`�vS� �'I��O0���MV7faL�Z'O�1��-+ķiq�'l�ڟ��I�O��$�O�|S��.�D�u�W6X��]�b�ۦ���<!���4�?���?��*���R?Ʌ�J1s��qڱo	/"a	c�UR}r�V��y��'���'3��'��9x�J �0BD=Zº���b,���.��ı<Q������O4�d}�X�`$2�Pxrj	�t2R��#Ρ&i��<i��?����򄘆"02�'^�J�ɆjȳI�Bu���2#�,<mZky�'4�	��I���Lt��⣮�e>P��ģ�r��Ie�V�M����?����?a+O:�A��y�t��5�cM�o��g(4k�Z u��=�M����D�O��$�ON���9O
�'j���t!�d�#v
��C֌�r۴�?)���ǖO�`�O�r�'��Tj�((YnȲ����#�i8P�h��?���?��D�<�O>	�Oz��h`	�I!�qaV��9f���4��Z>:^��m����Iҟ�� ���� 0���'���tB�
j^�E�A�i�2�'�`Tə'3�'�q��P놀�"|8�2��sn�l�T�iTz�Pt�b�����O ���~T�'��I9L@HhۣZ�4`@p0-2X�޴Rfb�ϓ�?.O&�?��Iͦa��	3��mX�ED����i���'j�e��d�>1+Or���`0Sힰ�H�[D��i}��s~Ӯ��<)�O�<�O-�'�B�ޢq-����?8��-�u��,,�7��O�us��x}�Q�0��My��5��~��,�#ƅ�g�eP��?����#h���O����O����O>ʓ/�V|���L��l̘ n�"j2}hM��#�	Fy��'T�IƟ�I��[�h�,�H�Q�	e~�GM�h���?���?�����$��k�I�'�\$tI�C���ܿ&|l�Iy��'���ɟ,��۟ a#Ag���?%_�e�@$O	$iݒ���/y|6��OF���Op��<QńN�@��ğ�� �����)#H�!��M�K�N��?a/O~��O �$��* �d'}/��m48�����!X�5ӽ�f�'�R^�x@
�����O����Lm�pe�->@�M	�,Ա+��V
�g��I��Iڟ ;��a�'�0��.f���+�'I��J���aZ�o�Ly��U'^6-�Ot��O��K}Zw �U
A�ٳU�"	�U/X(eV���4�?q��WԂd�V��s��}j�-;cr�=Yc��-i����gB���wl��M{���?�����T�@�'�ؙ��a?.���@�i ���$1sld���
67O<�O>�?��I�YE�-��KV4VP��)�7�8�4�?���?y��o�Ity��'��D��U5 ء�&

�i�IF���'��I���)j���?��U58�A�$Ej4��a!�<+T�P��i3���0�*���d�O�˓�?�1�J�iV�O?4�15��6��ml�ޟP"��m��I��p�I��L�IayRIK}��j�^-A�X�"�K�9�`��±>�(O��d�<����?a�P���A�¦�4"�"�SI��c����<Y��?��?�����@�@�5ͧ!��� �Y�[�Fkd
�b�%��IP���	�:��	xb���B�5f�P��8���OX���ON�d�<I3jŒt��O��@R!T$fu�`�7a�nl{@�~�H��&���OJ�D�L�O�=rv��v.Va��כ�i�W�i�R�'��ɏ.�� J|.�M��'oGh�@f�e��K��}`q
�x��'�B�Z	���|ڟ��,�.Tc�I�!��)6�i��I*+�drش}�֟$�S�����$��X3�Hl���^�a{�iI��'y�H��'J�'�q��uBM�K��Q!闆Qkеˇ�i�8�[CB}���D�O���䟸�'����j��2�K��`,�q(M�%��)�4F�������I�<y�z�<�QwHWa�p�Dn�&�:���i���'���@)vb�0�	N?������	1 ISPE�q�T!f��<����?��� #�`�K3|c�m�HR��ŵih��.bO��$�O�Okl��0,lY�e�Ճ}��k���"S�	P�'����П��	KyAY�ܓ��ݰ/����@mO�6�:����!�����%�T�����p� �Mq��N�&�PQYtkSm"�:��H�<a*O����O,���,�2���|�a�T`�@ ㊊D��ѡ�F}��'5�|��'4R
�yR��>�Zq�Y9$���+%��q,ꓠ?���?I(On�H��[�St|��j싈C�0=:*�
߆l ش�?�I>���?��߹�?!K���qaJkLXj�ኩ3p ؁Q�a�R�D�O2ʓ1�n�����'s�t`�?f#����BQ�p�tjp	�3Q��O����O�L$��a��HkS.4�#�ɪ���5L�:�M�*O�<�@�Qӭ������ ��'mzIV&�;�Ν�A�X@{��ش�?��S�N������O����B��:w[��31���>�P�b�4�Ԕ�Ҿi�2�'���O��O�Cx,����=����G�q��oZ�:g2����l�����䜑f���g�=��/i� �ӗ({Ӯ��O���B�6���O��'�?A�'k���0�܇��b�)	����%��#;
b�0��ß@��#R(nBQ:V�g�V�I�Kٴ�?�S�٪��dXJ��'��'K�<z�H��(9���R�8M�$�`�C�>᥌�%�:��'���'k�X�ؒP��,�[u��g�j	��K!� ��O����O
�d�O��4���-0�xl�iA�j���a��{.4�&���I֟d�����	�%�� �I.0�X��
zp`
5�+>�"d�޴�?����?�M>���?Q�cS&�LoZ5���9��x�!�NH"Z��?����?��?I���?��?1p`��E��	+��H[��8���H����'��'���'��x���ēx\�	�#��}@��.!,Vx��x���O�˓5��1&V?��I˟L���0d4��h����D���0qݴ��'��������k���W�� ��zk4�r�ɯ(����'B�S���'�"�'���]��-x�&�6��L�풐\�$��7��Od�dDn7,}d��ɘn�^	�悅�:���Q�ĶC���%U�a��'1��'����'0�O�,Y�'�U�fp@���-M3�X�r�Ql�qw1O>q�	$V1���c�F8a8�(�$-	 ���4�?���?�oȴ~��O������
�I�]�LU(�,�D]�p�/�ɤwǌb���	��I�&���tn�	tL^I��e��ش�?��g�+щ'$r�'9ɧ5�+��&Y�����`����Ьͷ���D�H1O����OB�$�<��́�BG���h�:JUp8�v�.[ ���C�x��'��|��'��&9�*��C$��.��q�GRg^��q�yb�'B�'E��'A�)x�՟��B�,�E��hwC�7����Ƴi���'�җ|��'�R��$��D5NG��;�U9+�Aj�mF�^�I=O�2͉�
UJ�0C�e��K���b��b�b	��t<�fPS,!�Ͼk)�D�tiڱy�
ي��� ;����JІ٣&��Z��0�qg��T�9
D�:d�T��[��{/}R�̈��!��*�μX�ءrg�ŗ>��S$iӿ|� *�1A*r,IS�;K��kw�Ūt�h���g:A�y��e�a��&k@8:cn����::HX���]��`r�d	�4/���Ȃ;,��'xb���Xff{/F)(����e͊��@]�&a����\끍�<�O�1��Z�K�&�q�ʐ!2�@`m�%t�4q�'j��'�*�p�%�<E��9!�0���L�s�(@-ژ�#b	��?�U�iB��?�G���B�VEJí��sڎ��5�M.,�}ϓ�?!�kl�hj�l��f���R��*̡ExҌ=��|��P�T�Rf	R),p ٪MH���?q�cJ�j�Z���?���?9p��4�d�Obe�3�H�K�<iEk2[��Ѓ�������ދa�����ɀ�x_����8X�-I�^i�$�
)U��I���z�)���%iX)�Ac�?�=A��K�1�����#Xr���/f?qE�N��	K�'*�ɱ=/,M��G"j,I��g˖|v&C�I�Q�LݑTg��W�Zpjf��3����?��'�9 �kd��x��Az�.,�s([���Tg�Oz��O�$�4u����O���:/0U0P��YR$!4�3
�z9�fb��e���	t�欆�	�:�<�r�Sd��X�1��/D���g�1w�t�б���)�T ��ɰv�4���O0YK��'t����@�"��y��#5���O�!�5υ5pء�"�F�"�8�Y�"O��dka��i�D�E`i�1O��'w�m�~9�OV���|zC��_��Q�@�	"��`�U�g�Ƒr��?!���U0��!`ʜ0��ƍ%�*����B��e6E"��N�U��)���u.Ri�A��-��Cv'��U��E0��Qr(�fՔTf~ИPb��x�,�Z��)$�2�D�O�?���e���"e��*��ayzI��@w����g�$]�q �%�� S�S	�n��$�g�I���;��7G/�[d%�.!�I�M�Pms�O,�$�|�[=�?!���?���\�	�&�=!��d�U�>0qf��&�(G	��:���kB*��c>�DHh[`T��ֵB@Z4��U�D��"��Ⱦ�*� �8vj�ZE�ċ[/�"|��0�Q�)F*46t�&�Y}�1#n�l��[~J~�J>�W�+O�)p��L�|�G)T�� �؂ӫ
0�;@D�1r�I��HO��@̂�`#�H3�P���`���N���ßD��@�0����ş�I🀺_w�r�'��<I��f��03��ӻ9�1R�'(���@�:��i�b�=O6�Q�/*�n�� �űB^����O���-(AB���d�\8�\zu�Yk���h����o�b|y4���DD�O�d-ړ��DٛWuh�Av�B�o*�d��U�#P!��B�&���j�����ЙFzʟ�ʓ(p���i�����+�+:�bU�۠s���i0�'���'�2g��r�'�)�;C�7��O��g)�%L��� �'8�����'>FdI�U� C�	Z�)f8��W�ޝD�0Py�"�O-�p�'4R6��k�}Cq�
Y�`4�f�@��lZ���'����?Iْ�E�JJ�	qn���}8��+D�p`��,s����VW$հTEv�;�O����)�f�i#��'�d���1Q��+ˌ�3V�	����Wd�ޟT�	ៀ�	̈́M*bx�<�O=�2
IC@���4^/MD�6�I�����8�'&��Br�]#0ƴ0Bp�D=5QGyB���?Qd�i��7-�O@�'k�����L��r�Q���8i�d��������$�>q�ar����#u�]�' �a|B5�dT�!HZ�Rag
�Z$�C���1�d��|5��m�@��c����4-�r�'�B� �D�� Rq4���m��&��,i�bb��g�';P����D�:�Dȩ4�1X�r�s�c��k���"~�I�L��9jЅ�dN:ܹe�%�Fф,�Ɵ���W~�'����@$'� P�YN|ڴ�	�yr�'"�}���0k�r7�Քu����׾�OEzʟЀ*���f�N1���8`u��,�Od��]�y��1$��O����O���C�����?a�N�v�t�V�X/%]���1�T?�qa��r�����ɝ~�fZPhӨ}��2�^�97���u��mCe�.|O�i�˂�����c<�2���O ��J�O���O�Y�l�	ky�c	:=y����`��Ph�Q81����y"�E�|�E� �P��qZ0B�Q͠#=Y��J>�?A*O�,�N�˺�AcErx�!)ak�/bv����X$�?Y��?��z�bD���?A�O4���,�%Q�6��D{����F�mS�p��d��p>�����k:~,��40IT��Å>@�n=�ND�I�l��I��<��Ҧ����M�9���JG�Z�R ��S�K��M�����$�O~��'|�>�Q�NV�0T;Ǡ��d�ȓR�]8$��WLu�pJ�k���%��Igy�Sp�7��O��d�|���/,�#�JD�
���F��%f������?���bW���@��&ul�2�M�u>\R�W?c	 ���1�q��EN*=�$ʓN��bP.9%�$�Sr��q=��s����Ol��Hܷ	LY)G�	r4����ߦ�޴�?-�8�jg��=0���ǘ�S,��4�O��"~�S��8�E.��������/->4��I��ēz�� ��Fۿf�\選y����'Q(|�d�+<b�'�"�O�0�b�'/R�'6M�DcO�xq:��c�Z������]0����:C�@�C��ق�^_�����>��X���W�r���J�ݬW���c@�lo<�P���-f�ih^2�&ܘV��A�pIӶX>��
I�����l�\$�i�>�l���I)�S��?9��J�e��Ё4W�?נ��7j�]�<I�!%Q|p���l�$-�'!�b�' �#=�'�?���3�L=��#��p`Ze��͑!�?9��:wuHiK�?���?)��ta��O����	o:X��F�7j��%2��8|h��t���=lO\5��I�G�(VV�=v�� ��O<��ѩL9z����@���&=?�5��f�|H����?q`n���Ӧ��t�'tRT�t�WD�<nB��pǮnt��d/&D�,9�	��q���a�_�9�<�(�� -�HO��'������oګX�B�Cq"��z��!�4�#� ��	���	���� �����|�R�im�T��4^��ĉSw��Ci��? p��ɴ$��l��Φ�I�S��ZH���-ŵY��)6�O�5��'��6���~�]��j˻6�5�s�c�*l���<�'r��?�{��AưaR�߃-�P��*.D��agkNm9� �@h.��(���k��+�Opʓs&h�FR���	A��g�^�LxQ�E]�ɂP�L*d����'���'L��`M3m:T����4Q.�T>��5�ZT�h��
�	S��ӣ�1�����"Vpa ����3S(9B���?Q�AMKh ά��Z$����!`+���I��M����R�X�v��s��	1/S�]F��O����/2�<����<�l4Afx	a|�L6�� nX�U@��Pǐ���H ��n�P�>Ot�!1̦�Iğ��O��<s��'Tr�'�!#��2�R��3kLin<S�C����"ط�� ���3hF��'�ϿSC�V�s�:H�1��u�PH1��15״�ZԨG�/���R��#�J�/B�:�rX*���fV"EO`Pq6�ד$Jpl�bF ��?��O����O�8` �<D�ų���?]L,t��:Ot�$3�O���\)������O<0lж��9�HOʧkRD���GŐ���ڏt���2���?���+RN� ��?����?�ƻ�����O�p�@�WN+|���
������O����GvN%	f�']�L*�+�^2Ҙ����9��3�'�F=� A�~L�ϓ\b�J&��04��;W�ʷ<4�`���a�����et�V�f��Y�@�I_y�� ��� ���"}���Hӌ�y�nΟakT\�`�/K<�B�*�#=�/��O�.;6��@�O�\V�8[��І!򄜡g�~�K�
�� �F�hS*s	�
�'u �� *@ +2�Q��1��=�	�'���۳��)* 5�͚w�ba"
�'�x��D�� ̔e�@�Сk��a�'�0���Ц&_j���$@�ykP��'��LAh�#<���X�o���'�z�:�EzN~����)e�$��'�>x"�AU��HdN0ML����'�H�Xti�V�-Z3��/=)�|��'�|�¢@�J�dP��@��1c}K�'M��r��s����s|��	�'l8%��d�\������B-zȸS�'��pU���Lͤ��`�
w��"�'�N`7b��~y���8�X���'�� �Q��D��T+��`2�'�tY1��,D� D�6fȠp�X��'$^�W˄*th�$�g�X9Ԏ9��'7�)��tb�g����	�'At��`�Ћu'���SkZ�x0�'#�����fÊ���M/NGP�2�'��	���G- T��B�ބH�>a��'��l��aG+Z��ǢPG�T�
�'K�aE]�0Z��%�=Et0��
�'$쌢�H�j�ܙ�D��&��R
�']~��&μKZ:��&%�t��Y��'�d���F�P�qv	W�Y	*u��'�� ��Ը��$A5�T�{6:�:�'������ "�q e/�ׂٳ�'7P�H6 xp y��\�|��e��'�J��Qa�;�T�S痖��<!�'�b*҃\�Z���PwD�R  ���'t�m!W�X�s�Ե�f�K��x�'܄(�¶tE�a�f�� 9��(��'$R9�U�_M2Hآ�D>1 �	X	�'��)� ŔB>���ҹe@�d���R�RM+��?`�ɧ�S�3K�!+20��y�U��_�Ҹ+�H�}؂Us�O�x�Q�H;f\E�7��K��06"�,
d�dXedT����gϜ�(}fq�?)��C�azX��JG
p�5E�m����J�%ւ9P�+V�i�l��:X$.űGo���0����6�N��A�B<;tf�X�l��0JB��:~J��"�O�(���Vk>?��M�*�X8hg������P�_�<����rVj�a�'>����7����d�j�8"�ȇȓH��sE��;���B�/ϸ<���L*�a�@�$Th͓~�q)�z�%��jG���; �%��a�tEP�fުB�!���O�V�i�B	�?/.U���@�Oפ�n;O���s�S�^����E�Y�F�+gJ�{�>�\Ѳd�EP'�A++[�ĪE�.O��B#$�e�JX�&,G~��I6��4X~�� i[&/�٘v���m�a�@�J�d���*|Ov-J6��֕�#C/v�\�����)�O� ��}�viA�=QG�ƘV�t�ɵk�6���:O���@�φ�JOx�hZ�=��B�	�WHxkČÜU�<��v�`��Qx��wÄӾ9,ű��d����|���A*�ͻ\�2��+��B��(v��	�0Y��,�gt@����$G��d�Y�+�V�✡�i��;���qGם1����;��P���|2����F�6��K�H�ؘț�� BT��"�n����=��%��-T%ΨO�q�2H�!�.Ӈ�K"]Rt�`�ȇH��=�Ν"=��1򷍟FԞ]�@�̑jb�(з��O�xc@�ɅL���"��~ʟ�i�o�"OFu;�hĖv;a0㕟��r���mmv!�d�m������؊*���Vf���i>RA|+��ês�6�ڤ�ݥIF�!їb�<�8�b���~���O�a ��3T���0�
9Dw�ۂ�&��<A1�Z*ø��i6��	$~r�9V �P���ZÅ�.>?��ɹ#�2B��q������	\�rع�jJ�?���!��-`;�8Z�)}�K=@vms��4��@U��צ)"�K�y4dT��(ܠU��M���b.Q���CKV�x�XA�Ʉi����OTrphF��F��M02-]$�"<a�2��ĠP�O�L�'����@-W�B�V)G1m�|�2�AF�"Z���a*x$�
v�SQ*��=�Ә*}��O�w�h����Q$.�(��{��;�'"�d\�J>��/͛4~��I�x�D �!�p(Q	�/�䜡��	�����Re�c��=���h��6(<�y�#�Yt>��I�vojL�F��5xb�dC#��>NC��ˤi�F�%B��H�D�`�%<}2B4�S��@�t�"7-W�lF�xP��=S,���*zNrɊ���AE���7�B�>���w�*�[Ն��:´��@1�0�E�$���y��ߨ2�,��:�?��'�JvV���
SͺU+Di�6v3���6f	O~R�¨-lfE��e�2^?b�I���'/p:�O�C\�����Җ�y��y��6���ɳ�?9�G�ܦ����¶��>�c,Q�km�m�dY8NmڼP �=zF�͓h����H>����V�'V� ��)#?��b��
<6pD+�'�z�0v��R ���dWT8�L �c֠�|��%�64��i��$�f�eŗ;������@�l˺+�I_������\kd�)��R=����w�se�SI�|l1V�x��B�x2j�D���ɳe�<P*��~�˖7RG����CT�C�<�b�X=A�򼲢*G=�0<1��@���5����%�ׁ<T �#�مx~l�sF�Ɣ@x)�>j�}�g�x��*@��5�ǟ�6NH٦OL�NM�r�r���9IB���>A�h]7l󒅐���@���CN��%gN|��+X�d9�}#�I-j�Z	�;��I���"�Р�%O<���.����m)�P���2V�i5�����mB�%*�FJx"/O��y�$ث-f@��&ƋQ���2�A̛\˂��aX0�ʈ	M��;A\"���M�q/�I$1��OԜ�	�+�睔j��(��ҧn�����H�.m���B��-�V%�y�.P1c$ˋ羉15���Q�йo�
&剹Y$<���!���3��ժ3_ę�A�>�������� �ҳ7{H�ٔ Y{�'m�<�uM�b�2	����>R�6$BҦƣ{׾9Ce��)�`�#�0n��;5�����'�� �r��N[X�\�B�^�9�T��1?��9��,:?q����#��q��I��h]��'�A?�e��S��*�H%��x��%S��Xp�W"�y���7o#.�@l[;��<BtŒ�?N}�2��I6��1O��������,���w����ႌ �Xz>��N��!�D](@b��kgk�d�ru1CL��]TT�"
�<����vP�|�<!0*��--�aE���lm�=�b	3#M��J:���Ҏʣl��1E�DlL�i~F�"W䕟.��B ��x���z�k�2�����ާ�Qn�grN8V��yU���$�\�Pe�is"#��0�S-�82�i�G2�(y���Y2�f���gb�&d�֙� *X�T�:Q��$A�Hс/s��0�Ƅb�Q+��1���
�>A"�R)H�d�H���,pȘHaF�SDb���B@��@������O0�/%nn@��n�?Fy�A/\��O�)����݂0��?������ic�C�C&h��D�גJ��87gƈf�:`��8+d�,�"�H����kg�S@�'�h �G�6+>�$�Ϟ�Gr0�����<8@�fK]tq��8 ���yB�k��%�ǎ����������9��(u�R)��ȂF<(�Aդ��7���Qq�'���@��W>>��S�B}"iX ��/�yb�y�~�cP/��A`x�C��w~���U�)&�2I�wm���c�Ej,Cs�+u��-q�c�X�!So��r�^�;d�=/^�%��jҏx��m� BI��f����S"9���E�܆(`��o޼$��b¯8t�l�JY�GHf�C��Z,���A�J�J�u�L�'5�� �\��|�.ɗV��-ʟ'�P�)�2����#N�{�,ZB%ږe��˓x)Z��	�(ۖD��\�i���?i��	�/�YR����T[U�ԆZ�1�V�q�01u�O��LlΓo��XP�	�U�U���AA�o)f�tb�@�"\X�a��� 4t��pg�_&�)��	�_`�S���!8��:3#�0/`�P��{�<�g��7;�(��Ư�(���O^��觿kc� -�������v���x�	�x�����	HH֔s�	��==;�ġA�֤3�A�Gޘ��Pc��P�.��xbH��)��o��=���T�Z���h��M��ݒ���8�!��	D�b�I"��s \��/�O�"�ɛ`zp��IL:R �<٣�
k�Dy1�5�7"���Ӈ�Ґ %��>MՐ��<�Ѕ��Ew�"��U��xƭY�N��)�G�0�a@O�'\�D̓�� �
�8���ߕq`ǟ�&�l�BF�%.sJ1ө]9G��8k���$��P�6���Ҧ,��4|p�+�z�������!pv�]�E��<���;]\=B�o�w?��k2 !4�@�m�^�1��aۇI`��	J-��<��i˧h��I�Jo�? �}�ARF�ԁ8r�:�v���΅E��D�cW�I��:i�B�?Y�GaW?j`�]ZP���Y�9"�E�OR�}�� ���@�t	�/-��3�(�&3��D� �T�d�6iM�@�-����C����06�a�R�6;R2��EI]D�(���i�<Yn�UV�s�)J�X6���aV�[�i�W��r��Р%sʹZ��9�>����$�T؅*��]Fd�S��S� ��pH&�^� b���L>�?YUcV2R��TM,mKf�NɆ�f$!��݁UD�вl.za�m�'�?�O|�	�0�׎ �l],3YD kA/%�8��#d�.Y@�yB'EF8���w XiR���Wp-��'�;dZm���o��sq�'�ҽ!D��}HIu��Sp,������$�&	�e&ЙL��hЦ�O ��ɂL��\�s<�a�|�d�O$f�*La�g�%Ia�-N>
&�E ��6R�fyp�,<P��E��_�|��A>=�L� �LQ�15pD��7+����7�D- JWW�aأ}b�'(��HcÁ�G	~4(��&|D�a��J�t��y�V�6��LP�O>�џ �F�3&�,h��ޤF8�����)T�0a����?��Lh��P�8�>�u?�Oa���h�bO��pH�Q����"KC�(�K��	/G�xB�M�.��$&m޹��̓\$������=Y @8V���m^<�A�O���	ґ"]�L�f�,^�ISF�.���D28�Z�J�j��%@^ұOp��ϕJ���Tbу�(���'�d"+ ���gS�D�p��'�)��� V��8^ $��;^8���I�<ɡI�so�\rC�':��8R��\��2�n���|��u ��F���OU�N�{��a�9Se���Q�źc�A��6��4M@���?A�-ީD���0R�ޅ8b�U��-G[�,2�l+r�R<q^*�⒫p���S��SP��B�gźl6]�`��0~t��m$��xrE��6K�d���i��e��J<r����3q�k��R��~B?O��i�hH�="˓b zʟ. ���� i��hъL�n�`)�h����'��4�e)ҕB�H��T	v1�82��~b#��>Už|b�t,��p"�"v���Q�OXU��D�+��T��1��B�'��9J�j����,6��ʅ`�#~`��P�I5<� �Ú���]3��I����O�'�_�	-Q&� ����*�p���o{��(e��yA�8�ÓU[N�S�A?!�.͈��ԙ5��yZ��DE��Q��îL�\���O��'J:}ڑa��7c��rV:� 2nL�r��}R�JJ�}"�$T����� �y� �Z���3�U�y.�YAg������i/��q��
xc�A
���b>���`F�2�����=[r�a��0۱O�%�"�Ք]m�����KPld���=�4�de�z�/O� �"���عQ.� ]�ώ��*m>�x�'_�`"�$���-L�Y��_�f�rȂ��ՁcI�U�չ��t*�%��^b>Uj�Zs�C�'�����B6�� 7i��R~8Ey���?Z��aQ��Q-2v���I�L���KD�(Ց�`�+:�d�@��`�C?����V� {����}��&V &H<`�	[�ѹ2��`��IA�Y������=2t�I���j��9˅�P��$Ɋ{��H��$Ο��O���M�CNí%�>%ZeW�M�M���V��Op�p��M7�]��`Y��6�	0'���8<|��h`+�
.�m�CS��;}"/��J��i��ȣ�ۊ[�}@ 3D@9z0�k�	Z�Y X�4 ��sS��4���e�gy�O�xQa��v��L���Ƹj�<��5��d�=D��T	��,O�見Ic`l�F�R�>�"(��$^�n:��0�+�.��U��gyI�>	����Xyn��V��R��l�����P���@�&���dO���;B�εYd�S�K�	¼!�2.^?!7�0��cT�)��i��-� Ew>�p�$��H��%"O�U���Z�$,9Y���S��%�p"O�8p�
ʂ6�� �SBO+.�f@�""OE�!�� +Dc���5mѠw"Oh�Q!KF�D��f�[WH1��"OX]���G�9��Y��.��&[r��"O�0��O�l��P4K��+M̠��"O~0#&���(��P�Xl-��"O�X'ͮ/�(�ZT��:t�6"O<<����Q� � e�G�"d(؁�"O��#���Y�L�r&��tcnq�""O�� *B��9��I]�/_8P�"O�`�ӣ��<����H_�EI�� �"O�xfgH=8ْ�		��H�K?D����"�3�8��j�\隭�/?D��A!O8f�V8�H	�zf*��A�'D��y`*	�7s��K�����D��	'D�8�G�
��Ͳ�`�#��A
ǌ&D��P�߰6W.��.]7f��)p�%D���F�^K�@��Y<rP@��	#D��
p����t��!�J�Xp��&D�� ���jO�gbHUr!�H.(�dj�"O%R�ñkz�U1'n܉
��	W"O�	P��F&�p �$¨�W"O��V ��bj򅑲���2�"OPQ"6�W�������#�� �p"O���w*��R=
4`A�A�$�x�"O"��bc�`a�P�X�(p�"O,ss�
m�@}StA�'i�A�"Oxt�3�]C���T�ܦ9M�	�U"O�4P�0'����R�խ#�Hp��"O�ԫ�,�3U����Ǟ�&Z�l3�"O6�t��$s�0��fNV�^�b&"ORX����'��j�A��Jm)�"O�*d��8��Z���L}� �&"Oa�B����!j��Mo(�`�"Oveq�iԴ��M���S&L�2�"OgÆ�ِ��F$ c4"O�D��ĒY-�iSR�V0i'J(B"O $�)j2ZQ� �ȕ
���""O���0�%[5n���!,zd�J"Ob�s���S�v��4Ć/8�V�'"O�����,̰m��"�t�� Z�"OȜⶬI8C0Q�����2��u�g"Ot=˓�ϖ6�hi �fɓ	��L��"O��R��NZ\,CF:�t(2�"ObyѲ��q(��坒*�PY�"OJ1$�^�\��q�B�xup��"OxA�p�=!��5q'�&>f`x��"O�LiRǌ@���*rDU1oj�ds�"O0С�̃k�ܓ��.�ٸ�"O49��L>��jĨE6@�mɢ"OPme�3 $�k���!�<��"O�����A��tH��z�Is"Oqjc��(KU�,�t�·m�z�3"O��9��ܻjD�
�Ϳ$�D�F"O 0	`D�:*���&h���ޕ�"O
��b�:y��#'�_�����"O��!��X9")�B��,B��"Oz��VK�#iN��W�A@@�"Ov�����%>�U	"F�k��Y��"O.!���Y�cˬ!�r�߻!p	�2"O��{@cH�`���Q�@I�:fH,05"Od�`%
:�C�O��P��"OT;�Ę�l��D�c�U�p	R"O�����,PD"v��#�U�"OT� ̙X��=`a^w�p�"Ox-�����;}n�@��C�UZ�"OD1��R m��h��R�   "O����D
aN�E2vf�l�M"O�����$ô�J#H�1O����"Oh����7�X� b'_�)�浺�"Ob�c��?$Lh;���P(��1�"O�,[�'�4�fQ��%Miv�Z�"O��P���@��qK!cӋ �E�Q"O�,#�I[��e��b( ,���"O�����>d#B(��gQ/�Y��"O�t�GI�,e\3e�s�x�x�"O ��T!nI���)y�@�J%"O"AZ.��Hp> c�����` ��"O�h�(�,Z4b��'��-���`"O�Pà*�Z,J��ch�#X�>iX�"O�d	TT�I="5T�k�R��u"ONY @C�(ȱ'� [���q�"O�eH@��a�`9�2��.'�$�aR"O� �xy厉1nBڵ3f���Z��bD"O�ux"dԥO�hub'��7S���f"O����	фL3\)�6��*�f�h�"O�q�e�e'��v�	-�u"OT�j�)[:f����ѡH:\���K�"OH�s���!��-�+K�H؁�"O�DA�.�B���J݊:��*"O0$�W*��j�Y���'u&ժ�"O�����S�G�\��X9I��"O�XsQ�!w8�#c)�
Ֆ��"O�5�M�a���d�@5�v�	l��!%EҶL8DI�d��?O���5�3$���DI���� E7=��L��B�,�yƳ1�=Q�C�2KL�c�Y8�yR
� �
d��P+�&h��$Ø�yBk�e��*j��q�lt�H�9�'�ўb>�h��E}�\�R #(� ��#�;D���QI+�ycC��?R��T�k9D�8c�-�I7\��%EЩU4�ԉ�k8D�x�6ˇ����r��)=�"#��4D��PF�$_����F�F��Ĥ2D��X��K�W3��	s�H2WM
���/�Iq���u� ��@l�&��*g�MI�|��9�~�8EX�b��)�ƀ֖l+�P��Q��y�@�F���s!��2&�}�ȓ7�vdp6K��|RU��j��o�"%�ȓM��Up���:���N�>@X��%:�0��Qa~�p�\�"�J؅�U��b��S2L��&@��f�ȓ�ttȕc��1pVusb�Ǆbꔩ���g}���0��Y��F<hx�`"Ucύ�y�G��-6��ҳ	I�/?X�:�) ���'��$�����<��E<v\��R�]�}����"O�Tؗ`�=D�S�v�@�8�"�S��y��j_f�Z���jD��"���yK_�g�TI!�Խ{�(�����y�"ڂh��9Jq�F�nn���aMA��?i�'\��r�3e�����5��' <�(r��y0��l�ij���'Y����CA8W��+0�˥�pɲ
�'�.lb�� b�53b���!��k	�'V�\Bs��8V,F�r��vl4��'��,hD��[�~0@1�>n�Z,{�'�z��$ȍ
0X�pl7>�+�'��]yT�*�@�
q.6ꮙ�
�'�" ��K�ipa�(�OP�B�'�h܋f#��Q�:�i�j^S����	�'�������.s9T��mD�NV����'1d�ąJ WP�x6� �xH�0��y�iڄ1���s#��-�������'��{�B� jY����"�fl�B%	�y�/[�3�L��\��8��Ɨ�y�ꆄ8��و��©[�����Җ�y��@M� �ьX�"<�d��y��)�j����,�l�w/Ǆ�yRjBr��e剴�|��8�y2�L�.PT�j��]�k���GC"�y�e���ju���R���I
*�y"I�"�I2�υ.¬�&^��y��&f�����o�|P�h�=�y��![$*q #��j��Հw���y	S'9^��{�H.y/�MK���yO�V�ƍ�1�Z�]�Љ�!�
�y��N��`�!0�@�!ﰼ0��
7�y
� �ZDg��LyF��F�pE��"O�U���qx�sD��-�$̚�"O h�!��kn�`0c�?U.>Qӑ"O��*F�M���T�� <A!ca"O��c��(������C7�Jh�"O�D��& 9���!��A����"O�cAl×��xd	�� ����"OzT�!
Y ����ũC���"O@�!�\�j�"(��n:b��hy4*O�eې�B?��v�K� ��O������l
ve�2�J�<���sh��!�O8 �H�Y�|�; ,��6w��"O9+5�&a4�z�	�Pԁe"OB����X�1UPT�B�H�o�n]�'"O��/[9z{�u
3/L�^U�*O�3c��Z,�F��'ڼd��'6�H#���$W���ɡ�ɱ�:U�'z|"� �D߾њf(_i,\��'b���k�#Uʘ(� �^�P��0�'�,ɡS�T�t\a�E ��ڽ��'_}�Ƨ�@���N���)��'��� 'C��h֣�/K����'Z�cGK9��jt� ���"�'�"y��U&|���0��"�'U�Th߈9�8K���<�2"OnIs�7)�����Q������q�O��]�G��D8���l�:R� !��'���8�iX�~w��P����A��'W
�(v�Gb���Ƽ��'\:� AK�-)���aՉE2=��'�y��ũ�2Ai�6Ob~��'��Qz�/O;jMBѪ�JƝ2�����'�Ɲ0��u��p�Ů�/$��Y��'��m�aӞ�>��N=#)B� �'�b�bȐ�i`D�IG.nlɪ�'���ru���>��ŒƧ\�j�x�9�'�ڵcD�x܄�IQ�a$�Y�Op4Z�C�*3~h�#0K�! ��}z4�d.\O����;����!��"g"O���M�9d}!�L.,�xa�%"O(el�m@*����O7!朱q"Oj0�4�G�l��R�m(�॑|b�)�Ӝ=$��q���7���'�4	�B�	u��4J�葃h.\��&@�Z+�C�	��rL�� �`k*Yhpd�� �C�?&�p�����0b�����-rC�I�aH������5g�\`3��3�\C�əvmXD����4*��8�$�Q
^��C�	'C�`x�G�g��M�2Ώh�C��2RB������+6L"���J��B�	�51FA��P	>��P��E98�B�2Qj ����H���RT���B�	���	� G/�y2��V�V�fB䉫L���rɇ>FѲ�)�J|F^B�	�6K�)�W��D~��Ga :Q��B�I8��x�2��\$P�����x�B�	�E��-P���J� ���P�B9�B����A���ҟrʶ �Em�5��C�,/�Ȱc�+m��XR�^�9|�C�	�-����çP!��0��� BB�I$/D��5K�(j�✩��B�	<<(6��d��.8u.�![#Ay�B�	<@���:BHа>r�{��b��B䉰&Fh���`���J\�:+�B�)� x��ƫ�%�ڑ	 唗AՎ�ے"O����&?�R��'�A[�q�G"O.��E�ڧYm���°a[jaH"O����8vN���M�u5�<��"O�!�A�%}2��JQ/1н��"O���腯M�d���	� ��"O0 x��C�i�Q��M��@���0�"O�e���;��i`�N�Bܠ�##"O����N1!�ִh4@	!�6X
�"O�q�pcȫ6�h����.�X[C"O��������ꆏ�z׮ȳs"O���䁍F\H8�H�!�
�+W"O\���CO��*��ȯX���P"OD<*�mB!Ͼ5�P��#�8|��"OL��m�o�Ԥ˵�� cǢ�*�"O�E���.D�L�  "��,`1"OҘ�/̑A��YK�Z�e>A�g"O<Zr�	? "<Z���>^��zb"O�T� &�.ː���6Or�C"Or���#>_"���)Ȁ�B93"O����s��asÕ26��=�D"O�ѳ@�ϔ/~40
q#ƮBFT�+�"O��YO�]����0-��	:�D�!"O�K��e3�X��w3����"Oj�����Z�cƮU�$!���p"Oph!"K�d��������֜²"O�
G�)|!�Ƒ�F,��"O0U� ,���dP��!@��P�"O*Hi�L�[�r��p��b��B�"O��	!)�5}?��b�J�"/��x�A"O�ܓ�A[31Y�B"I�Va�E"O�0���M�=s�U���(�"O����
+��Ѡ�̈��"P"O�@����4�h�[�O�B��u"O
��M(_/Xp���(X"O���ꙊxӾ)�#�;=�l�rW"O\�#U�ā�j�)�H9C�C'"O�t�b�?H,�JVkI	9��m�"O`h�e�w��@٥K[7Tnv�S"O��1uIP1-�h'M*alt�hs"O�M����I�\���޿W.�x�"O���ӗ)�)?��Xq'ۦwG!���i��BL���*@���/[�!��E��-"��X1�,x��Fp!�D�+�\9�̳5����6lO�V!���#�nвP,�-�B��3j^,�!�ڜ.H�XbF�|m���S�F�W�!�D�Hذч� C�p9���đy�!�Ă�EA�D3�cW�w�8�t��g�!��+J��4��;QDr���nЙa!�,��0⬛#d��0�pT!��G���TY�˴U^*�H��a!�Dª���#�ė�iPx)�5Ξ�GT!�$�	*����N]�AA��3�͇$X!�D_:װ9��)��j��b����8�!�$�L��l��kG���H슂
4!�D��ߦp���8f�l�%�"t"!�W�
^Nm�蟩o�pM�kց!!�$C�����P+P'WK:T:B >j\!�D��9�6����"d��W��7>!�$އ6R�%���(<X���+�1>!�D��A�۪�PF_��k�ϸ
'!�$�_i�� W��x(x���D�-!�$<	�<�iG/�g�tQba��!�� ���V�ق"J��3������T"OX�je��jr�رpGݨ$؂���'t.QK��8$켉����M�]��'
f���$m�s�C�:	�X��'n(X��K- �vD�s�ȏ �*�d�<��")F�z=P���j>ms��N�<1�M��L����u�O�L)�� e�<���X5��Z�[
e+����@Z�<�D�3g
԰��_�Fm���O[�<Qt�2UP�@R���%t�A�`�M�<�w�oO���Q�I[TMB2hAD�<��͓�'�I���� ��S�W}�<�G��+fD�xvn±P��x��j	b�<!$i�
i�I�#�x砐�@��C��5*n���ՏoT���d��E*C�I"U"�|P��\�T�j`�1�ŁB��B�ɬh�8�
'�&"�r�r�O�$#"B�	2�.���J ��j����+u�<B�X��������)�T!��C�qj|C��<���b����`t��(mx$C�ɦ_|��C��P-3�4L�W��O��B�I"<�q;U
>�RHSIU
Kk�B�� b ����c�6\I�ťr?�B��;zd]��	W.���Dxq�B�I��|����YL���M�?�rB�	:w����@��N�(���j-\B䉥}��j�O$�"'
Q �,B�>'s�L��$x0D$�[ �B��=v�*�q�`�:[(� w�Y�q�C�O������(r�d ��\��B�I> �XA(��&1�;�m l��B�IXk(4��ۦ<�mj��Ԛ@�nB�9?O�$�b��`�NQ�.H�m�B�I:Ov=�� >���7��=tǀB��0N*y�/�eM���"� 2�vB��"d��!��
�tQ�b��f?$B�	�p��5`Ə�\��*��K�u �C䉩:����=���@�Յw�C�	���<��EF8{����0$S>w�C�I�	�5)q.ה3L�:6�Զ��B��6}�j��fI�٪�Q��2T�C�	���1rbG�N�v-r!��?LC�C��2ri��s�����*���.�pC䉆v1fa�h^(Y�<=Å&�u�<C�I���4���DO�.���H�	q%C�I�Mt"X����Y���!���B�	3\��Dh�	�m�5�ad Y��B�I�v8p�"�(
=&/X�C�
;��B�iif��\/�)y'��5���R"Oإ�u�6�bQj�F�OPn-y"O�$����+Rvx����!��y��"O�D��	B�|�.H�NL�w�,�"O��Q��
j`�� 4Lt�W"O���*2?�)Sc��V��t��"O:�` ��+C��8w*��R�"O@C���*VTXi�C�����KA�<�G���S�D13�Klh���@S�<�K'[�<|�v���^`N���#KM�<!@�[o/r�u�=4�R9�˅G�<��.E�$�F;�%Ϡi�x�)�B�<i��Z�Ct�� ��]��u���@�<1��=~a\�ڐg
-xV�a�k{�<qu�L6m>��P)] `��M�<Ĥ����wLW��(+1��O�<� ~]Y@N����P��C��P
"O��s��0�(Г'H��k�|YB"O�"�#�>*���Fl��SA"O��A��Ƃ��%�����R"OA" FU"
.�1dɍ�?��i�B"O��;���R�$�+SIQ�5�\pc@"O\0�A,V��|��h�1eE���"O@t�C���&��V�Z�r�"O����h�� i �жٚFў�p�"Ol]��� �Fe���Q*��p"O �3DtZL��B��K�4 "O 	;vχm��\��'W�(�H�"O�Ir�4]�Iu�ށ%Ƶ� "O����6~���ȵ�P������"O2X���P�;�vA!�M�>�\y "OZxAbaJ/��y�U�&��i�"O\��"<N����b�?AGv�b�"O�1��@��z��A`��@.��"Or�f�d`z��d.�>F��5"OjH0WI�+�j�┬��w!�e;�"O�E9R�ǆe�(!B�yf�s�"O�8�ƢA�Nрeȡp�*���"O���L�*�X��C�B�]��c`"O�<�M����l`G�� ���!�"Oj��d咜*�2t;C��6�(�v"O��fA���0�	��ŕ�6���"O�\[���:b|�`��L�!%��L��"O.���Β�P����E=s(8�"ON pÄ1E-*�Eɱ_�B���"O<�
����T+u�+��H�"O��#�XO��)I�̥>�
4`F"O\���j5`�2���#�o�P�"Oˤ��MT���"�3���� "O©�bᝆ/ �b�׻�dXQ!"O�" #Ļ>hR�f�
"�(D�r"O�`HÍ�0o�~��Q��*߼5!�"O��C0/S�w���ڔn�v��"O�s2K��y��l���A�A>�D�R"O��C�54���q��"$,fQ�Q"O|�����?��(D��T ��"O�@9֌>a��U��IP�hŀ"Oj���/Y�����RX��`"OVU�e	S-p��;�愗6'��"OJh�n�#tP�KP�O�8X�3�"OX�ѫ��e�� G�ebN�yB"O�yg��%Y��US�&P�Z�
=��"O�m#�bBn~y:��κ`�ԉr"O����#�t��Q��*�:G�x���"O*�a�űa��c�gH���#�"O�lxe�;�p����07�mC"O�|Y��#ӰI�Qe��\J���"O����:'PFhRFٟH�X��2"O���E�u��aJ�C�1`p� u"O�#�E�+�h�V�ӃQ2�X�"Op�s d�q��ӣ��	��y"O��8THC;E�J)Cd,H�M��6"O��p�a��H�q��� ��"O6��슨q�0	�h+O����"OHi�A�0Q�ĭ`a�V)xT#!"O�y�fH�>qt��x�G҇�|� "OtIR�@�2���ɱ%��X)�q"O��R�ѹ]f���� �"O�還��<��#֡Z7����"O���5D�1Qe�&.0��W"O� B�
��[�b����ղn�+�"OJ�35��&M���S B�g��p6"O
� �B['R�E�b�
�OU>�0	�'�0��%/�� h@P�3Z( ��'�DHb��4j�8@�g��a 	�'c<-P�UD�����+B S��Y:�'B���!�)a>� ��3C	p��'�*(�e��T
LӳE҉z4���'B�a*��G<M�u�W�9H6Y��'��u�ͫp)��Y'my[p�z�'�$·��>C��1���+ *��8�'��1H�m��5�|��Vo�7�a��'�hi����� �RY[��@5e`��A�'����Ge^�i&�)pHǤ+�}
�'������E�M!�T�e���+5v��	�'z�k����~覨0$��vI*�'M��[��%QKl;3O&$�<�
�'�=Zai�	 pB�I����(�
�'��@�J4]�~\�a��ݦ��	�'4�\0Q	,q�4�KQ��=t���'*2$�d aU�*�H8����'��T	˖�4]�uÉe��I��'���Q'�
�`W
���ȟa�dՊ�')" 6o	�gO�<As�J;Rb��'��Y�R_�0�(������'���š¡���r �n̨K�'$�tIt-ȟ+~P��-B.^/0��'�t%�0LJ*D�8�hV�J����'+�]q0B	�Z��D�(<J�X��'p<
���1�1����D-Ɯ�'J����k�`�^�?��a �'9r���T&bP�V��6�z}��'�(�aG��N}��9���7N
�8�'o��&��E���+�mϥ2'����'K�<�%I��e��{�C�.���'l��Y��:o�٫c�\��	�'OZd+"�<M`�ۗ�TE���'Y,a��J�4q�x*7IN&�~��'|��Q���9W�>�{���..����'٢�����V�E �
�8	�P 
�'�t	�I\"&��qG?p6��	�'d��^�~5�� *<����p�<q�Р�R�fM��*Ӯ�0-5D����E���h��t��3��q*�#2D��k-�O=��	 %Ρ,4��V�/D�0�H�^�M����!>�Z��1D�@��g�#t犱B�	KL��'�3D�d���Ԣ�i#&M�OF� ��2D�D���$ܜ��l	-��b��1D�`���~x(�����/U����@f1D��Q7 ��8 ���X����2�-D����M�����pV�p�D3��*D��ⰋD�S�  	���؜"�I%D�R�A�b���MНd�=�w�5D�Ȁb�F$Q�,�$H�>04��C��/D�H��(��I��u3&��x�4�+"D�\�FOK�7<�aN'��x ��<D���f�S(Ᾱ���
=��P�>D�T�U,S3_��A��2��%iю=D��:D�Ӝ$��@%Aț�e��b8D�P/�L(�%c��>%�l ��٠"fC�	���T"���d�$Q����TC��
�\���f�-��l4�Вwp�C䉏=�h�2(I��0��Z�&��C�)� @�Ȃ) ɐт��	�4`�0p�"O$�%C	 ��}�P�G���)R"O|������@�h#���N��""O�t�dG�aOb������ɣ"O�0S�N�c��hr�M5@��Cg"Od}ʐM*o��$is�T0ԅi�"O��7H3�T�:�jq����"Ot���(=�����T�\� y�A"O�l2e�a0摢�GМ/�ꌂ�"O"��)JA���QU斪%�驤"O��k#9k,t�eЅd9�Mx"Or��	�.m�q�����m8�١"O�ZA-6������N#�q1g"O�	IF �
Q��	"M� �d��"OVfD���#1kA;rB�3�"OX�d�$R�]ұ� H��"O�J�B	�l04��'�/AK�	�"O8
� 2;�a�ŭ��6Ke�"O�����+�d:E-Ц}��]�#"O��!&�ۇzX�y�,�
��"O��`ЦS(B�AbeÄ�H�c�"O��	��v�Ve��cÑLƦ�"O�h!�!�X�%�B������"O8��4h�)�<Ի@ѻ3��"O���C�����A"a �h�9�"OJ�8�Sak"L��ƴk�|͋"Ob%�.�\�����0x�ɛT"O��yPᕓ ��)�Q/J���S�"O��5�߹n�.	yt��9��9Ce"O�BDL�%�
����R�vN����"O�����>x�"k=$�
�"O�t�"�Hݞ�2�J�, (HHPE"O~u��@A0*ڔS�邥cu�ك"O���֤9�^�)G��?���S�"O�cv%�}���ӷf��ё�"Oa�wm/0�z!�-2��a��"O� b�lۻDֽ��%
�P�p�q"Or詵(N+-@��Ǥ�7�f��"O^Ё�K�<~���%2)�Z�"O�1ҡ�\&0̼�[�d����x�"O�ejU���\�fՁ1F=�(lhS"O�p�@�X�lp���b��`�  ��"Ov �@:^$l Ă�(0�$��"O:hX�	
�\؞t{�G+|ؐ0�e"O��S5i��x� ;%�
�V��l��"O��P�J�)�|����ۍ-�%a"O.pX@�#�pܘ��B�<ʤ)�"O@2"+�a��@��K�_��Ѻ�"O�����ᆹ4a�p�<!6"O�Jኋ��:yң%�'S�<�
�"O�D��<�c��D�gPذZ�"O��آ�Z7v(��"�d$��"O���a��#m���#a^�l�bg"O:԰3�w=&��.��
�޾�ybI�y#����K�?Ǥ��6��$�yB)�;4~�ň�hU�/�B�4�y�	�����ᇶp(�i[0���yBmO7<�t
!
�z��x7����y�������h�����)��yr��"K���V��B����4�y��L�?��IhT�0�E�u�އ�yB�ڛ���%ÁiW�x��1�y��C+�ZEQ��_c ������yB�Swyl���#�P� ]�%d�y
� p�V�v�5�	H���"O�+F�p喝Zק�V{>d2"O��"ō����H0�O�2oy0m0�"OTH�E��:f�1���K�5�Q"O(�9��14<D,A����y�n�sW"O����@�:u�B��ѩj�}X�"OZ�$']	,��q0ᗽ_r����"O�e�V�� E�b@^�7"O ��%^;q>�(FFGb�E(�"O����fWoX�\�w*X�"ΑpV"O��1��t�>01��P#(p�a�"O��{�d��+6��$E���"O�-�#5V�<Lcĩ
�Q�zM�"O0�EB֤	f�@9GH~�$4A�"O&H{��C�PO\|*�GH3�
���"O�a(�Þ�x�&�&�o���"O��S�Ťd��`$�R4�|Ȕ"OJ��F��y�&lcգM
*1p$ c"O,c4�PdH��fE˵l�N��1"O��pb.R��=a�dT8T��8�U"O@a���^D:eAm�(1I`"OR�(��dQ���A�����yr�M�@�F|��gۅ&]�؀���y"��)I���H��C� ���� ��/�y���]�P�&G�� �����ybe�����p-�x$JЎҴp!�d*�HAPD$d�0����:S!� �n,�"爤���r���B"O������,����(��nu�u"O<���T�Qzn��,T�e����"O\���ÍM�0L#���=�t 2"O�()�)��I��1ԇ\5S�"OD�A2+J�7��S�N�p�T"O�0�F�={lX��@�+���r"Op��еK|��j�EǺi 
�y�"O����<D��⢊�F�LE�"O��{th�E����A���X"On$�r��43��d#��9"�M�V"O��g�С��4�7n���<2`"OV�z������R��R�(fiB�"O�u��)OZ�ĥa��4NU�yӁ"O�hX Er��I*��@�G�>q٣"O^�i4c̄V�xȻ�J 2t���"O���$ئCi�M�D�\���"Ob�p!��;נI8�*�4�i�D"Oh�9V+_�'��{�D�"+�f�	"O���5�;,5�0��T�@�E"O��Z���2E��j�:4�ʕ(C"OF���m�,)�4�tj4�Ä"OF���(R�i@��a��E2d"OF(�B׮8 K"O'jhC&%"�y�� 
-n��6��=p�Ҵ1f�Q�y���W�0��i�#l���"�E8�yRDگe��H�k�^9L�)�[�y�)ǧo���p��?��A7���y�X0}�x}�䏙�K�(@��y2�
�U"8��� H+`�2u�V�y��%W0E@WE�P����?�y�hI,?��j��\����4�yb+t� Eq�B�>O$4��LV?�y���A��AthG�|���+DB���yB���$�>I��]7},���c��y!��F7�E���q��Tjc�]��y�������"�A�W�F¥��y
� �90���"�9DjH�
K0�)�"O̜�%hJ?����5^8�3"Oh��L��΂\��\�ri�F"O\�S�!X�3�rx����*�<���"O�����4%�}�wh��Q�\�"O�aH�N�Ԡ�A�DV%�h	d"O�A(�C)`6r]iʓ!J�I%"O^ ���) ��4dhŹ`�C"ONp[��=fV�l�'�����&"O�!�I* 5�+q%�<R�h9�"Ox�r� F�,� ���N'N��P"O�,xp`�XD�ۂ�Gn�x�Yg"O&<��Y�<�v��R�������"O�M"�b�צ�"��mHX��"O����-
e�P[��/; 	yu"Oj,X�����t���c 0lp[E"O �Q��)��zAB��{�5%"O�ez�L�u疽3d_8��4B�"O�H��ᔍ�8[�b�fu�h6"O�JBG�1��\��
K�ib��B�"O�%��	�rB�{��޹@��(y�"OXB��߿#WXT�6�c��Y�"O�ib��MgN��#�AHv�:`"O�qUG���db��
pV� �"Oв� �BtA'��Â�C�G!��!s1�͏m���" 
֒�!�Յx�\�*�G)hb�yʰ��<[�!�D��E�h��C�Ui`�xa��p�!�� �84癹r^Pp��ED�0k!��Ax�t� ��B�ƌS�C�
�!�d�?Frʑ��N�	4�j�ۀ-m!�¦1�%A�o�'>���AE�Wi!�d�.3�(���[c,��S���F�!���t*B���%N~�|���V�h�!�$Wd�lQv�U�v,,Q�É�!�E:�n:W�Mb�x�u�30�!�6P�dX6�)><`̪�A�,M�!���;�Ph�E�֕G�����<m�!�$A����"���k��R�L�C�	�.rb�x�iZ.N �Bb�K>T^�B�	.h��Ԣk�"yf����mH�
��B�	84�&C&��,�n��kȕ,Z|C�I�Fkv	BWI��z�:)�F�ŧ|&B�ɕh�N�CG��0,��RiC$�C�I"��e��T�60�S̈́6���IP����l����[{r(�b�iS�`���A�5D��P�#w�xx�f�Q9Iʠ1` 5D��"�b&P�h��O�(Qb����3D�йF�!i\�t���L�HNLy�*O@��Ej�Iuҕ{U��)�] "O���V��$~���B�,`Z��"O�I��@$�0m��D�x0ؼ�q"O��0MR;&��݊��={M�D�3"OvL��O݋AE\E2A�<v�P�"b"O2\���À_���SkX��|� "Ont"�kS'�ʽ�r/G�t�ȹ`v"O���ǀD��Zh���T��E��"Onlb�(Y�6�A��؀n��"O؈���?I>��2�ds���"O�pяY/ZF�����O���1"O|�� ��tt��#!ΝM�4�"O�!� �,Q���JG�^>p��Pp"OZ5p�@�OE����"�:�	"O����2H�&����[7"�4Q¤"O� ���F-M�8��I�8v�y�%"O@
�gL'������D�n[�l�"O�I�/��A�Z�Y,i���r�"Op��28�3��|�nX�p"O�u� �G	νY!�T�M�rHSP"O^A�V�˘u0zY��,��rY�@n"O�}�"hɃfsv�{�!C�#�<��w"Oh��� ȉ(a�R���"s.܅k�O� *F(��\q�s�+]BL�J��O*B��=>����_�Cx����,�B�ɸNo�X�$�E�@v(Rơ��|��B�I�}� �W(-j0�$�ƈRcpB�	�c�����%s孲W�9c\�	�'��C&HB� �$�ևD�T~�-��'F����N>d�\h�փ�Y��!�'a��� ��=97�� ��^��~�S�'�D�� G[�gEL}�e+�$J����'�X�C�+�7k�Z}�u��;yO��;�'���17�.~6^�,�u�:�2
�'�N����S>���F�-q΢t�'W�x� (}k��Z&fb� ��'�ũ�ȃ���<1e���a�<��'���*&F�3<\ �k�W�Q
�'6N��g^�l�/�N���b�'`���#O�;Wh�����B!:zf<�
�'�F4R1�.�d��r��7m�x:
�'&m�$��J��P�G�S�&�H(k
�'&!+�.�������vux	�'Ͷ����׎{��Ѹ7�X�t����'�E���[�$BǁJ1I��!��'�6(�7�<��VIG�1�'�������2�͊a���2�'����\R��M�'��']�l��'����V�A�`��x·�"	L��	�'�"d
3ȃ�;KP�bW5DX s	�'B��VE $Fռ����@	z��l��'WA
�\ 3�f��#;`M܈@D"O(�ȗ,
�|@d-��$@*�w"O葲����L���bɢO>�C5"ONH��C�;��� $ζ#.8h"O<]�n�
?���v�U��̘�"O�At�X�k�4h ��)-�n��7"O���O�2FA�䓷��%{t�"O�)�R
�/d��Tj��es�uzG�' ��ȟ�G{J?�[�nV�q3�(Y1"�C����&b=D�<��hW�A7�|x��3*{D}Ba�5D��u<�vea,�/2���5D�T��*���1f#4aU6�c�'D�ظG�H>w�"���♼y���ǀ0D���bh�>(2�4:�eE�8�H�@"-D�(���LO�r��b-*�zh�	 D��ڢJJ/�ra�~���f��y���*'��L�t���jK�1����y�f�/%��U����Pi 1��F��y��D���A��M�>�pt��y���7%P�iц��Bw�r���y�,o�����ڨ7�"hH$�y�$S�s��X�-�pY�����yb�.�UQfe�3!��a��`���y�阚Q�f}#��� �舳��W��y"d�p�%흗z>i0`
��yB��?)zƕ`�b��6�p{F��y�
Z�����	Yt.)�._��y"-�NH I�Pā�'E"l�%���y
� �Qf�	�]����2�HIr "O�}ȱ��"~���XWE��Sڌ�҇"O����Y]{�Ր���;����"O���%ѭ����F�׊h�h�w"Oԍ���I� ������Af@�R "O �@��*��F/@	;j���"O2���f�Ѳ�o��_�պ""O�t��[��d��c� 6P�h"O���O�B�X�bD�F'$P���|��i>h�ʍ֟�&ě$c���AVb��z+��ʅm�s�<�瀼/fn�[��!�.�z�+�n�<��!Z=)����1N�"EE@J`)�s�<���*�p0���I'��F�o�<��m�.7��Q�G%һT�hiD�e�<�q���\Ҭ��n:}��q�A{�<�)ұx��"V�E6��hƬ�x��~���O���3q�SX�plC���U�Z�'�$�(	"���%�Y:����'2�{�`�%}�j�J�L�9�
�'��ysE�Y(���cD
�DBЀ��'16��w%��A�#Iwh�Bf	r�<QǪC�Z�@�M�5n��s/[S�<��,6;H���Ԇ[�\���F]I�<Q'�Ėb*�!�F�G��B�m�<q7K���Բ��τ���a��e�<��Y�[M�`RbF�:�qᨆd�<�3GQj��a;ѭS�"iY�E�<!�+�+����	
�����W�<�Ө[�2�:Hs�c�k0��Pŋ}�<���D�I����塈�i���iK}�<a�i�~�T���#� x�T`�Rn�<A�厄ka��ZF)J�LȖu
B�l�<��
,&]8hCĥZ��ȹ�s�a�<�rN��BK�)��	��$N�p�u�ȓg#�qAD�;���{�iR�x-�U��#�!�V��DE�y;������$Z2���� ��c��χT^� �ȓb�%��ꔣVB|cd��* "��ȓ:  K�:*�jDcD�%+���ȓ~�X�a`��� { ꀍV��T�ȓ8B��a���#��-����S��E�ȓY�B� ��FjJ��ǃ�/�:=�ȓX
�("c��&�n(���ٺi�V�ȓ,r�ѳ�EP���!_9K��!�ȓ=�*�;��������4�� �ȓjM`@�S�N�c�e�\�!�ȓ7��5R���<��ĭ�-n*~U��D��.�=��$�G�V,RT.ф�utp���N�;��A���! !�$B x?ƴR��w6����'?!�'Iei�Ҁo2}4#U5!�Իh�@�b@À�t�1��f3!�L�S��s�$�Y&�E�-!�DLW�m�E��� ����&Z0�!�$B�~�p�(ą��2?H#e$��H�!�Ȟ<�Lٲm�7�*5�7c�5g�!�҉>���B�mF���:�B���Py2�U�H���Ǌ�=�:T�!��y"Ń�Ī#��2vD��QR��y����J���ra�s�БV�J��yH��3�Ƽ����y)�8!�
�yb,E8<�X,�ŭ�bF����y�j�>
����	š##�]������yR�Ġ""��&C�
R:�@h4�N��y
� �D��� ?|�+��Ӑg�z���"O~��AW	\M���"X��Ř"O�yW�@-p��E�G��h3�"O\h  �6eW>X���V[���"OlY��
�"�e�_(*C��$"Of�A�]�i���K�3?l���"O�)��Bˍ+Ƹ�0��	2<-��"O��ce
(�;�D��%�U�1"Ox�B�р[]�È)c����"O	p�H��$�p莾-�b$k�"Od�cA��# :�1V�
h��	"OF��C��%*=3�e������@"O�ա� �x]��DKi�xY�"O��8r��)|��r�̗2�Pc"Oz��LA�D"v⛤�P`�"Op�����Q1��b�@L9�(�CG"O�D02�ߨm�N�`��Czv8r"O���s)��A�ub�:��,Z5"O:@@;����� <kf���"OT�:��H'~6����iS?f�@��"O$�3���:�.tS��q~�(��"O�E��!�I�M0ˑ�'��mS�"O�;�Ȏ(>�A���=��ɺ"O�,6A�����S��M,ֈ-��"Oy����(vg"��س.`l;�"O�e�Ι*3�<0�	�!\���"O��`��B6b.b}�ӈ�z�\�ѐ"O쑁�	>2op�h�ᗅ5��#"O�0iWB�d�!3O�Xq�r"ON�J4�ێ@����!�G g�4"OHp"�Z"���K��ɿO���i"O�L!bBJ>~���Uΐ�j���
�"O�xr���^t�h��O4]�c"O�ɲ���=�����጗5xf�yE"OFD�R1J��`?�9�%"O6"�L�=e�(3m�%> �ۅ"O��)K�)r<cu��$*��"O6q�F�!��,��3pH�"O��Est(��L�
���"O�q�C����J K�H��;�"Od���A9q��@����;�>��"O�;s�1z��(�ЊJVXJ�"O�Ƀ�N]m�j��V�[*�
G"O��z!��<<�-ST#T���f"O&���hʴ
v�������C"O$��&��%*Ȃ ��l��]�f���"O	��m²Ll�*Є����"O���e�͏f���TI���L�R"O^��!��!&���$�#��		�"ONac�g�$u�˵K�h���"O��@�Ǝv���#祓I L�s"O^�P�N]�\�͓sE=(.�uxg"O���`+��7E^��E�X8����"O6hP�$~��� �z�V�y�"O
yam�N���$_�\s���"O���� ��L����E�d\x0��"O�hrOGq�}��-[*^?f��"O��AE ++����clN�?L�b"O,)���B�x�@�%�[4��"O~IHf�ÝpR����7%x
2"Oj��5�6;��ӂ��<$�م"OXu�-��`��iB����+�)��"O�X{�%��3!Z���gD^����"O�LCE� 4�;�F�T{���S�? �a�A��F]�y3�&A��a6"O6�0%˕5+@ȓ���(4!�!W"OvE�C�3��l*��˂I	�d�"O|[�"�=.�&�Z�[$	�L��"Oj�V��2!� �飦�%v���"OD
�J�#��\�����%�q"Ov��3"�(q�]`�S��4"OrذRM�U�ΝR�H��@^9�"Of�{A����xq���A�B=Rj!�S�3�X(���J�Ydf܍iU!��O2N����)���)Vf-S-!�D�N�L��G��f�{e��0!�ğ�6�l�2�&<��<��j�>^|!��K	0B�bA��q����<)N!��%	�ի����z#�eh��M<!��T)
/|�Ps�J$
P@�5��V(!�$<YxyK�Ub��yFf�.1!��4n*�:����Jh����߬
!�$�d�puA��P!����ĢE�!��X6ez��-��(Y�C/�@!򤐉4����W�f�s��ӺH!�
�D�H��6I������л�!�K����ڱ��8��E�cόr!�$�x��h:a R�c�f����	�+!��B"CIt�{ED�$�����m(l�!��ܥq��i�RJ
k���JVl->�!��]e"�S�T7g��-�w�ۭ4�!�d[�s��QA#F����]q�I�!��2D��0rD@ �<�F����DP!�So-�QuH�"i0�!D�?!��K%�Q�,J�{p�K D��%�!�7g_��{w�T>f�s�b�	�!��8loޖ
03�r`"ˊ|9���'5�Q[c��>N�܁@��|f� ��'y��6n�[5���H�r�t] �'?��Ҷ$�-�jT���X�r��PJ�'�P�I� 
�䬐����x5��'[�X�1i�g7���̈́M�L��'��m��卶n�
 � d�
@ʂ�`�'/�4P5&�aDy����4�>� �';.\ ��9`>�9���ٵ.��I�'�.0z�������fS�W� qs�'��&"/HŰ�$P�8�
��'���n$V�0�Ι8A/����'/����n�(d͜�RJ�";�Rp
�'�μsT�%��0�a�Η`?ܸ��'ytYv&׌3��I)A(�k�|��'��q���+M��x�p�4y��1�'���R�-P3T���I��L�n;�,��'J-)���
�]𷃍k�1�'Q�=*$��xnU���j�+6D����/F�H�����m�Xq"8D�`�j6P�b�IC�L�Q2pM#D��c)ϡ6	���M��@Y��� D�l8�hO�bo�pH�33
���&?D���҅B
��8�S�H2_�P�A)(D�ģ��ͣj��\��.E,ss4ġ&D�8gHP"<��hR���3D���0D��j%�״z��=S�[-4����J.D����C<k4D���ivP[�k D���-�i�&�·�٘R�l�#4�"D�XI#GJRN.�yw�����a�a�>D��r�kCT|ذ�ˬ@;�5���7D��*V��p�8ApB��2���!D�� ��� o�6l�䘣�G	},��"O�L
2�ػ�l��H�&�\�W"O�LZS�[�k0�\	6�A�,i!�"OX�6��R�^�va�"+$dab"O&��狒!.��qQ�� 	�,�pt"O�]�'��F7D�j��3(�(���"O
��R�3�4���1l��x0$"OP���B�P�,����2]O|C2"O��#
�&}�$�S�6֠Uzw"O<M�Q�p��Z�#Y�x&��"O܅��f�u���jrW�r��dZC"O�8z�/��gt���C�@6��uA"OBSi9%�Ȅ"�<9}Jt��"O��
0�߈������@�"O��BF�V�M�h􇇗^���*O.͘ e��� r�`d��'��X�ǚ�c$��k�F��i�L�
�'ص�ؤ_�nӥ�U�fp��	�'9X-`�E%&:t��%ռ`�J�"�'��D��+Յ]�R�����9&	LyQ�'� 	���-q��}����	g
�0�' �� �MQ9(bn<{$蒺+��R�'��Zf�H�v�͚��\&m��,B�'�d|;�0|:ܨ�S�R<1�L�
�'�N,[A��-P^���F7H,��'��b�<��83�"�t��')�UR Ǖ�v�^������Q�'��q�qR�tR�t�=�J�h	�'�t�`��
|2��R����0�j�'�@u���p���ݠy66 ��'R����R* �&�q��'�
�z��Q�;����4�޹�'A\��G%#��+q�Ȝ
h�S�'[d��A(Y�C����q��8��
�'��x��3N��}�F⎜hƩ�'m ��Pl%u�#V�\-Tyq��'ߖͣj�}�X���M�6<5�ɲ�'���(�(�'#�6@��ߴGN�,{�'8U��h�<�7�h}(�r�'Ő|j�-ʙ3� ��閝����'S�����[+X�DԺAMI2�=�
�'�|��w�[+V��䂵s@Ȉ
�'��*���8;br���/wP���'�,��tL�4��!�l�l���		�'������+4��#P���'h��F���ta�B\i�	�'}�P�-S�8�� ��DF��8�'�L��,�*'�8�hpB�IK�$��'c�4B��όD�!! ���t���'GLL�G#��P�1ǉی
0�i�'6
D�t��A�V͠U�3Vup���'��t��#Ҍ�0q��ѩK����'�Ν� e
�wR$���EWc�-Y�'�pMajD�:��Bh�7nR���'�)'�:h���s��&,����'��y�Á�?��d��Y��q�'�HV��l�	��D��=�D���*D��H��
(����H��[~��GG+D�0��ǌ[�\�1dE��)��j<D�|���@&R3DQ��b�n�zV)/D�,`2fޕ/c�h���]�|+6%%�,D�X�Ɖd�*|�@�+9���!�I/D�t�v�R���w�X,,9|�hq#/D����[A��z��:c�zQ���8D�� ���q1G�p�a��#�ȹ��"O�k�j�-O�LIf�è�����"O>�r��a�a �(�+eR֔��"O���E&\�V&LzA��Ok��&"O
�JuQ�z�����l8l8"O����Q������ ~ �I!"O��7�+S�<q3��R:8/�6"O��R��(�Z8�C	�U-R�I'"O�'Fw>� ���CrH"OJy��f�\z��RS�_Ȱ8�"O�M�婔�"!8�qЙf"O�h��+e]~�rGo]� #�l�S"O��m��\U�;��̯y0!*"O&��F���$-|��(j�"OJd���x50��*�7��uR�"O��r��@��TR�HF%0�2���"O��s�oo�R���)���9""O����D�� HI* ���yS"O �7$^K.�,P����"��(y"O��� )@�|~���WC.|H�"Ot���V"c_"��oܡ:,ti�"Ox����	/>�*8C����/�4�P"O�����U�9 �`&��#/�Lj"O�uH��(�VPY���>)��U�"O���͖p���R�6�8��D"OH2Fo99�䅻7k�.�jl�7"O�M�#�4�TX�'�X3$5f݋�"Od������9,xp�
-���#"OB$�M�>>�Z	��``dt}�"O~  �V�b��m٣Ҿ��d�c"O�Yǎ+� ���L�GgH�"O���j�)��|RG/S(g�v��s"Oz���9�J����FD��#"OZ�k�:Uy�h��n�9*-���P"O~�@�`�^�x�P��0�ѹ�"O|�!D��M�~i�3�o���XW"Otl�5�A�]��}��ϛ�u���7"O�Mjw��k`XD!ʮug`@�`"Ot�kĹA�d����Jq����"O*`)!�M�f�:P��?��%A1"O�����t��Q9�9����"O�l("c˒~J����U�?��U�$"OF!�g�U3Tc��C��L�`�"O�Q;����~Y���Y��D�"O�0ё��/x�Lu�T T�l�BQkr"O^!�I^>w=�-�V�Qz;\!`U"OH���Q3AV�U�%�U�n0����"O�9�õ�Dq	��א.f�S"O�x��-�U�y G^1�l]��'�.䩵+@�C�dhd-"�ڹ3�'jҝ�@g�w6,�D�ܓ�|ɹ�'�v�3���0�Đ�ΐ�h��R�'�6��Ή�d)l0#��dl ��'��c�.8v��!�=_]�h�'e�Y��K�C���XB
c�.���'��@r
ُ@�-bV�B�S�h��'����󧊿3��Bu�M��A��B�<	@l�%3 ��(�L��b��0�D�@�<)bQ'�$�x����;��E���Yd�<��.�	D��q �����ċ�f�<Y��D�#E  *���ogL�6/Em�<qF瞈�|l����ZO�AF��q�<���{���c@dΝ]4��ûw�<�&K�.�D$;#՘BS�9A�L�<� �	��g�=hvҁ�
�`*�U�R"O�pp�M�6����S��bL�"O$P1�����Ç��3�,BB"O��K��>q�e�Ԁ#%CN��0"O�$�X� ��}��@@k��i�'"ONYP��OR��q!a]7�h]�2"Oz��6 6���+dKS�L�Ll�D"O� b5`�!rmƘ�j[�bU�9��D0��)�'S�X)���]C���4���ȓqO��ѧ@S�-�<��L�@@X��%�tec*�`6�d�[y*Z}��v��5�o��`4��+q�S:b��=�ȓI2�\34�B�c�DI��f�x+�y�ȓHQ�����A򈆄���ȓ,+ �6%H�Pb�[�������ȓ]:T� g�0�L
e�#*��ȓ����hR~F$��]�
����Y�.ay��"{� �B�9,`Ї��G�'�L��fP�a D��i��a(�'n��k�w���Fh�2����O�x$Ў"��)1�P������"Oz�Q,�+w�(]0��V��@!��D#|O��KD��8�ȓ���f�08���]x��k@�4�ڨ����.,PD�*D��@��+�Vj\*/PI-$���$0?�-ٖ(��IǪ^�oX�(*V�c��E{bM���c�
�� i!qKW��y�b$4�e��(�tyP���y®���̐�or� <�J�-��'0�	r�O��ɩLE',80!V��l'���fh֣�yB!�l,� �k�9x�,P�@���y��)��-����h�eJ�
o��<I�,D�	�!�OFq���Ŋk�����%���f��L*�`�3]:iSe���B��H��&6�O��j��)# !	�.B���bhU�$O�L�� ��ؘp ш(��dH#*��G�* �OV�Dz�Oo�Ie&�'�S{�h[�'�?D6�͓��	p���q�=2@A$"�U@d�9SO-�I: �Z��$�!��8�`+àR����@� ���$�_�x��W� �J�n}كl �ഊ��9}��Y��4�0Ǖ�P �����<���Ĝ�O`�q*C1dsbd��� 2�$``"O$e؀���M����0`���Ւx�BLl��(��5�$MP�F��F�p�0`�"O�)p��1:�M	�G�vU2���"O
�ta߆���jd��6�,���"O��a���4�l�� �e��AQ�'3b�=���(OX!8��E�Z�%#���0XF���u�'��c���< ��@�@�!��Y�"	�'7!�dN#"Լ�֠��N��x��	�����D�De�.Z"�O�vmA�-�y��.,O���"ۗwJ^L���@3��=xr"Oze�bf�{(�=0��Ԟ80�*OЅJ�+_5���k���=���	�'�rLY��Y�&���oOe�	�'`QG.S 3{�$��ÖV�F���'8�11�����h��Ğ��ı�'��p@��a�"M)�J�7���I�'J�žp��@�a��'� )�ķiLfu����-�q�'1��5�����q�J� OA����B�)�4��D��"�(~6u2De�#�y�cH�M��D�O�o����b �)�ybaͳ[�U0�kQ 1[d�qL,�Mcu+�0�?	/O��G��t�? d�J*P<  ��Z�=?| "Oh20h]#
l�;&��*#�d��"O�M`�ᐤV�	�R�ޓu��T[�"O$b��J�T��@�Ǉ�@�����hO���3W|С9��Y�Eab�`GF�=5�!�$�`�Y�P��|h�/�=H?!���:��e �F�,��4�g�;�!��-_�$ �č-BL��%��!��5H,t(S���[��Ay�mS+y���⟠Җ�D1ʓ������Z�g.6�!��Z&��ȓ��ɧ.B��jLiV��{�̕Ex��)B��N�V��hB�W0��Ls�+�X�<RB�4_X ���=�( [�N�<Q�n�"&��!��O%2�f�ga�'�?��b哶*��ȶ��6����m�ԇ�	�oSdU���VL��� �P�T6�C�In�z� �>n�ǮN�x�DC�	:@�@XZӇ�*)@� "��oV~��{}Ҙx�Y�4$��ݖ������H�$aj�b�[�C�	�s�3���MqLɣ6�η\����`؟ܸ�eA%=sK[zv"e�3�H>OBџ�D����4e���w��7- �f�h�J	�'�}�m�b3"�F�"�X�O�z-O�ҧH�M��˧uD��3f @�"O��Z��̞P\�@䄓�{3��3��B���I�9��wFط[���vOұ;!�D3<lD@6m��l�P�(O��=E����V}pp��7�0Q3%���y�BǇ!�TU���-?��������y��|2�'�*� q�#�^����U0<|  ���Mh�d�ju�!��h�HH�T�w�!��	=��+���$Ep(Te��֒>Y��<%>c��ْ�2S�U��"�|��s�>D���b@5D��H�+\�H;�,B��<ɏ��&u�V����ٛpv��H̟8�nC�I8�djs.� (k��!ň"AL7-[���?Y��8P4n@�GIѕE��X�5��c�'C�'�r��|�D ,5
���m7 ��yD�b�<�s�
(�t9ⶌ�1�V(zU��_؞`�=��b˶>H*�X@�z�����/�[�<1�i�p�@�x��� (��`a	W�<��!
�HA�9���P�P܂L #�M�<Y�� d��,��-D	5bJ(�"MVJ�	]8� ȅ����.XHFj����9A��#D��͖C�
D��
��o�����!D���h�D��`��A����r�s����0�)��]y4I�d2Vu+��@�N��"��1D���&��C4��#��Y0kkp,���+D�8�7�ؼl�
��2�C&�TH�2�+�OԒO�D�"�����r�Źd~��E���b�'U�����7:p�c�&��x�h(I����	"w��9be�Q�_�T�h�l �v��C�	������
?���Y4�\���O�˓��S����Bӎz���@�ېc:����u�0���7J�D���
[�b���h��t��)�tK��#�Ǝxhj)FzR�' ��j2�\�+�>�2C�\�߲�YCO�x:7��;Jεz��*���:1"OF�r�HϦV1�;�ޛeN�\�O��Y\H<��bˁ�:,,T�B�Id����'���� �GBG�$aP� EGD|r`"O�ܪ�[�VQ��5 D�a��"O�p��n�Q��p���aJF Q �D,���$�	+�`��Z�g�i�c�ƛ&&!�� Ԙ���C�찹�&W��]���	ix���2�E�7hy��(@3i���B;D�|�e�շ%��M����qM��Z�3D��Ӄ�V�2!F�Z��R0����0D�Hs$gԑqzLj ��Y\�Ha�.D�h��-��U4h4fL7	������/D��J�ܘ$b���J�rT�R�a;D�pi���p��yꁇ��./\(���5D�8مl� t�@��&��i����&D��`܍f�]k�b�8O���SE(D��3s��J���f��rz9{Џ:D��v�Xot��&� (�PpRa&D��AT�r�J��&N��ZMyB@9D�l
QC�r_D��p�ͨ�V5���5D��D�*�Z�����8�$݉�#0D�h	�K�!|bحh#��.�$Aj�I8D�Dɂ���8t�U��&=HB�/5D�xc�e�v�Z�Чf�$)���+4�4D�H�R��h����%&�R21D��0e*-+n�K���/�R+�O+D��)��P�~eʧ���1֐����'D���uP�:�t�w�	/FŲ�s�e*D���aI��a��(0%�L�ؔ�=D��£@�8�&d�5eF~�Y��n<D�\sWNQ�Qæ���C�:XZu�R�;D�#��ȼg����ݞJ�\b�o:D�H�ˎ�S���@GK�\f�聃�"D���f�4sp���[�Zkʐ�%�?D�|!��#%v6����Y�<��H���>D�4�GD�L�����
�Բ��8D��DB�v�BM���6�����;D��Ȣ�ճ7|��DÚ'/�*�3$ ;D�X�2�QG�q[0ᗈmW��g7D��	'nT7��8(�J֢v��� ��3D�)��)��$6`�6��@���<D���QFG�ZN� ���F�U�7D���ӥ�@�����MX>�8�0�"9D�����!�r�h��
4  �"�+D��ʧb��U#�eK���[..D�L�%��&��A
�IK�erB'�O,=AQ���f�@$`�X�&L�u�-��:�"O��E��?b�#"G��h�s0"O�	rPF��	��Pb�_�i�z�"Ox��F���DJ�@K>t�^b"O�1a�ѥW�j0C��J��J�"O� v���,=�n۹E���Y#"O���U��AbЬ�͆���]�!"O�����@13,^i����j�"O��#IV�� $��x���2�"O��1i	-%��P`������"O�Z�	םkA���Dھ.�0��"O� xG��F*� BdO�k���9E"O�=!g��-+�\H�t$ �o��c"Oꌠ���F ����h�^� B"O�e�b��}c�P���"�\X�"O��vOs� � R@�<��uj�"O�p�r N�(�e�&$þ AʝkS"O�	�c��e�F�Q�ؕDMnśD"O��#IS�;�( t�ԩ
q�0"O�U�Gʚ;�Ĳ���	�@��R"O�Y��I� f�Hj�b������"O����d	=���0E���%-���|cz���%+���,���C�V�O��U��8	hB�əe�\�ƪ8��al��vR,���̪��0H��A��S�? &����@�4ja,ъP��� �'�,�U��%B��L���G?mY �/�
I��xJ|����4��ZR�H�b��x��7
�<Y�ǀ������ �1��$�Ɂ�\�zEy��5nxz�7E�?�!�D����Η�T���H���Q9��O�U�l�E�E�<�)��0�6���|o�H�ěv����`>D�(F'�����!��U�P���߁cu�e	AI��|6�`I}���3�ur��sY9L����@L6zS ����b�X(��4O�h�W�j���I�/Z)8��RU�ǵrm�xТ�
|ܶ�� ݮ�p?� �Q;+&�|/i�܄s'�acB��{��'�͸�M̌�	�
�۲���d�!�<j7٥Dd�8�iC'g�v;����y�C
>mV!{�`E=f���_7r>���S&T1  D�#���+K��y#���5y�^�c�NE�珻����	%�~�Y�mлn��ڣ�.�	�A�^��q�)P�U|z��#�n�2 .����F�+H)@��(O���a�ߒT��I	ՉD�v��fh#?�aP�̇-oǪi��S�4�"	�%�_�C�z��V�:����A�t��֌��-M6�Z�M�X��bt�F�k�X����A���� H��mk�aψ6���?�:=�M�%	���\Iɒ�R�dx:!,/���{aU��8�zEJG&1��r�ٽHaJ��ӭV�nh*џ���I�n9A閌Yی� Bg�#3���H�K�nnA`���0|�Ǝ�.\���
W8��y�*	m���(�"+���PE�IR���̧\��XQ3��9�I�l���"���Q3�؀��Z5*���ŗ�.����e�Ȓс̯+�Zl.�+�1���a��=z����F�K�?����'�Ħ+���Hn�m6�l���>x5Dp��+�U����V����/_�<��+rr�@`��dJJXK�aU7���Y0I�$4
��p�$5��$�?�� pv#��ހ}p�� uw\�c�̓c?���BƐ'�l�d��A{�����,A(`Q�l
C������O��2�b����D�_tz�u7H��B4\���3EPn�am���p1���7*;����E��l�.�d�#æf�����y��E�<�@HD'�0_O�	AT�F��X6�G���sF��;'���@��|�#Av�r!W��<-束%������:tnF�;����*���	+�r��ջe�<)��{>�ʠh�8qb\�CL�*���Bx������7���H�7M���\݊Q�ؚ|�a(�I�?>�(O��������"@��V�=��*!���<]ܙ�� G�up��ci!�$ǐp~���)��h7��r� �C,Ru6��#��7R�"ػr��z��ݻf�(8�nYEH}yb�ڴ �������� b���!�&ryvT�QhB4�<��fh��DyGƷ�0c�i���������HJ�j\;��cbK�C���yg�@w�
isBď�&�,��l^�r��Ig(��?E��';��c3��`J��2�K��ʔa�ãI?2[*}`�dX�P��H#a�%>:��ScB��Z%��6��A�w�4@%f�>Qc�83�� Kfl��'9�*#Ę�M hrU̓N* (҃Bj��2����y��(��4�؜Y�c�f��G(�g8x���̛6��Q��`���6f4[��^ C4���3(4p�s!�³#��#� ��'��(�c�:!z��CF?�<k����&<�%�SeߚpePk��̷M.�Y�%Z�O\�!fE1�����K��`H:���D���R<�3�>sɲlkSυ�+
`D�9�X�S'lJ43�J`�A��D���<p̴h���s�B-��g��0qJr�HF.�ϟ��B.؜p���>E���+<���QΔ, �u����-*�r#ɹ�T�" �Y1�lx �O=���.���Y�ec��~��ϭ7�npQEF�t}��2a�A-��ɮ#��)u����%��^D���X�k�F��2�&���b�S��I�v���*��}@lޚ&�	p	Y��Oh�r�ǹ(��ہk�Wn���D+3hma1C��O4�q���Z�,�Z��V�?`p�DI̟zH�!���/a{����V%��ܑ�d�B���j�U��I������0��/uINU)�ۓAz�0�q�[;t�n��+�}c(O;rAW ̼�Q ]�9cL�i��[�Va�C"��J�<Q�/0z�� �۝}c���rS�,<����!���'�Ȋ-y��Q��C�y�<���ڟyj����gI��?qF�V
D���r���|F�H�˂Z���c��<�Z��a�1~�B��'�K�~utE�@A��l��öh�{�L��gVFP��N�h����*Qў��K����T� kA:�� �C(�Ɏ;�� ��/��裁m�����c��<\�0�R�J�<�V���[�Q��!��
5r񤹚�JD)*�������s&AUn纝���U�����	�`L��[8[�z+��ظ�����h묵�+F2U��;VzР�O�*�@�b�WK�مȓ�h$�O�iv�`�N�u��|�@J�;�e��Ǎ���HW
��b8��/Єo`� q-��q��H鐺i�\����N�j�2���<TH82���j�����V��5<P@ 2�~�dK�U���Q�](R@#���v�����~Aq�Áo��	1��pϮ�S���f�&,���&$���	4=�&��q�K>aWRH���ߞ?�vL�3H�F��FE*���n��8�2��$��e_Np�2�=�bd��HS7`ʐ����&�L��g�<&.@kvlX	���x���FK"����ށ�!f��_}� 9䎎8]�L��`�΁q��=�LE����ŎL�8P�I�#]~��(�u����AH�"iC�+O-th�w���(`Rx�1,7]XN�OPp�q���^_@MȤ�7y��ѣB���\i�Ņ��O/p�^�*�i��W��e('ϒ�UcF�R�'�Xa��u��y�ɐ�b�"�Y�N�T��iw���}oZ�J��A�rK�D��i�5��
t���*�)��d	$)�4^�-y@�FI��M�B�F��}�e@�	rذ�Z)�F���# �|*�$k�W8]Y$���E;5x��"�e	h��EÊ*�V�Gy�.'+�0�F�_�X��B��:3�b�M!�v��5j��z5	'��(��#%d�
��P���xp�I
0R�xaA��	>ށ��⚈Wo�	�V�N6�Ո��		:ҡ�G��Rc�9���O��� v�������P�ORF��t�D,����$z�IJR�>E�Oڰ Q�NSr��7I"t{�`b��
sv��s�IK�3���$����!�H<ɇ�PNJ	+�a�y�&]�����y��$�T1`��g�Z��8ajܴI}���S�ρ��YXQ�i$N��&i�|r`�a �R8"إ���9k����g�� .��=լ�p�e]�P)BU���w�����-ۍ0P�:��!RO�l3_�����ǚ-� 8@*�(&o��t/i�f`E]�pњ�X��ͅ4#�%	U#]�mY�-� ��D`ےQ7�%D}�E�L��i�GG	�Β�k�6.�H���&{q�0J�̩<�¥&r���i"H�3$�6�[�yT�l�4�ʜ�.���K3�p�Ƒ
/�ay�K^�e0t�&��R�q����� �:4���cA���XK���A΃�G��͈�N�2�������;�"�Jĭ��[��
^D����.C�A�xq�7��~�����(K�p�nOV9Ss�QR���Z��-�R�C��3xM!�Ο,B����/;��q�f,�G����� M��F��M���(O��pMNK���!��6m�j��<� g��h��&(�|��"�X�!f� ���L���)�L��p��e��8�
$-�l��RM�8	X�!Q*�1r���D�(���PQ��)CwJ�D^lٱ�	^x�,de��mS
�~.0 q��CRP����7r� �هC�`q6q(�O�Y[j��?��BQZ���D%Hb����C���m;�&�k��D�����W��5+Sc$-$�a 38CE�"�tA��G"�
�.�
2�F�P2�F��?�!OX 0許sK�� �z,E�F���9i���-M:h�'�ֆK|�!�$c"�%?�x�Q�ȡ}߀E)��>h�0P��l�'�8�M��J,�'�ϏXr�Q[.hJTm	�y21':D����.�p��ܟ�qO|]y+ҺmW����OP�4��D�W�v�.����� �IS�̄!�~Y�;H�M���þB~��#a�<]R��*Ǟ�O���i��4|ST���.A�fx�I�4��d?�M�'e��	�0��I�c��}�E,��28��)e�*'���b�L���)�B��ðl�6�V	��ؘ:��UKu6o��j@a�LF5
��S���,h��,�p=��"�63	^�����l���M]�OTDX�s��"w��aV�
����4�At*)��ď76�!���~�����#-N�ҺoD�Y(tE��q�@��g��P��}�'Q�.��&DS�G��$���>H3R�P���{*]D�L�04�t�U�'���@�B���0Ó�J0P�H�iH�x �Dݽ`dTq�� g ,�Ѓ8���h�n���	H?�����΅`�����p�jᧄ#:�^min=g���kǭvZ��h���3殜�r�~�*���;K�Ls0�ɯ/�Ā�.K�3u,���ʀ5Ē��2O����X��úI� DS`,�-+�ШCq�1p"��T���91�Y��$B�`K��
�ѓ��.�x��D�4Gcn�xʏ6^�c�abNx+��Ѫ� ��8Gn�(�@D�Dd~�0�Mˌ7^�$A��g�.	o�6�qq��h9�]�t ��ha|�%>����b�T k�C��t � �r^���E0v>7m�",nҐ��m,�Pf�F X��Bע��i���O Lqe^7~IZ�
0�U�"%��	$%=L Є��?k���� ��Vm�DH'��!ƁӇih�)aLV�Q�(=X�.��d$I�F���|�K/ C�V�q!D�'�J̐�/�}u⨋� ק���+`̄�Z�e����9Nf]����8�^��Oڅ~}�����z���S���_��A�i�Dp@5��
HE��8c�؆T��MX$�'�X�
x��䣓#��2�2@@ѩ@�v��ā��?>Z�3���hbߴ9���Ǉk�M� 2��k�i ����lN967�i'�'q̥�ả�W�ށ��X�q��#\�
l�v�C�I�,�ŇݑTQ8�����k� ��$A]t�5����_�x����O҆�6v�|�d�K� Bp��@�Y%�O�9��L�h�l�j`���H��z��N����.� f�j�)v��p�t�c J�@�>16M��dM�AKLF�?�TK�+`��lh�	b"�x��O�?�����玆WIJ�`�"
�<�`Ż��ݾ*t�H(�䔈`'�X�3�V=9����(!��ՙ�!^�L�{&	G�2�sg��*��ڤ�'~�0 ��� j��D�$$��S&�Ac�
�N!�f��OB��#%�3t� X ��"m��p��dʹW.�y�w�d��*��f�V|�t�P�(`
�Cof<���H�8�-�2f�q�%۶c�7*�L�hŁ)l�!Jg�Ѳm9�H��+ċu�B4�R�� r��#�5.�F�P�Oƭ#B�!5L�I��愝���.q�qO����e�waJ|�&ɳJ�ʼ�Ө�
Pd��Ƅ�,�BU9w��)X����o��jn`��B*U�w�.���̌4�-��&6�/�V	Y�!�D���	�#�r�ɳ	W�!��
=pl�lzbh��9�d)r��X�%�H�3�F�& �f��c���$ʘ�Sf�����}���Ĭ6�v���׼d�Q��������B�J�,ZyR��l���k5�A��s�+�y�`����8P0�0���V��8J�獗i�Ґ[e���
�� Cu�!�y�nȯ��͚@N��.VB�g!�I��a���q딕@�N(ҧv@t��CC�;��!��B�QyM�g�ڿ<9B=(��� �ig��|ܠ���#U6��yq
Tse��-����g�	i�!%�X�=�X�k!�W�|�����'�����\	]���M4���r����
�΅�_���"b
��Y����K	����qED��𠕯	/5,��H/�RN ��*����'2�"����~�"H�7Vx��-Y2Z^L�'h�*$�Ay#%�%}ь��d>�*�HQ3_l�'-�VF`駈]>k̩x��+"�$ꗽ.�����܋ٴL�=i3NE�hS�tq! �'U��y�ׇ߇7��s@��">�+�	�%~��1��P����π3u�ڗ�����_�Tѭ�e� ��\��0���^�D����"U�\ 1� �aD�\��O���	��r9{B��X�~Uh��ѫj+��h ��?��K��|��B���ii����m�p�W��+T�N���&A�G ��f�x�����Uja ���$Ëe�d��47��&*V�:�Z��ɗ�,w���A��b�f��*�o�`���ǈ]%+�U�BD����>L���`E��#�2	��X!�~�K���6��$2�O�z��mI���8`2<<*
 '�>��y"JJ�$�*#����M欙���1	n��'�ͲV�`�W�����	s Wz��$c)@�O����!Iۺ����!3�Fq Y�WXJ�s���	����Q 7��1!%�վu^�c�49ue�<qT�QS1@^+K[X��YW�4�"C"�p�Hel��AI�(PI�!�ݱ4��
'�, qD<��Ч��Ke`� ZB�� x4pvcì_�%�Gn��6�eʖ^��� ��>vrh%�q-�7v8,�1AW�	��k7������>��<!q�_�c��x׍��n#L�ѳ+�I�r�`�r�\���D>��09A�ߩb��H�mT�m&D��ûie�������� '�
'N�P�&O(Ҏ��) (~�(�pŉ g��U�|"�E�F���e˵��t�M�.�Zs�*VL�l�`��$��rA �#1mX�:e��4��l�=9��C��2���k{@@ǥV�X�M�,Q�p(��gD�wTA�ˀ����jGkzBhEхT� Xᭀ/T�`���&�A�~M�5�P	��#N�9KdL%9T�7�IRJ��eɖ�FԂF�⨃�nS#)���C`�WԾ��G	�/jϘ� ��>�`ae��8�t�l�*�ם8QLq�B.����$$�R=��o��.X�x�DD�/�v�'\����H�g]X钴Dҫc��ApaE
k���h.�$�!�'Z|xT�C-�Aiu� y�Y����B7����W4&#}��wZ�h�4
�j���P���R�H�o�D�`�d�T���zu7�� �U0V��eF�{��,M3�ă7�ܥ^z��BF��v�8��d�=z��I��Gn>#>����Dj���"���
�0�2��&
���@ߤL`����:��y�H¯F
y���H6bH �-ǜWx\�1��P(Y��LxPCFs�p���`а�\&�� P��Վ�������%b[�������5B�3@��D-�)c��t���Az�V�cv�Ǿ��OL+���	���?��%U�w�r���{m�u���ޣ�yB+9���� �K�C$��MY!��/69������)�'\N�ѷ-[#l��5j�QBć�798PK�O�+TB4
�)Ӭ$���=ф)֒Y����$#B��	�	N(><����8�!�
I|��2�=ut%�q�=z�!�ď�>��a��M�#���;��֐�!�Һj��թd��Y�*��W�A�3�!�$H�'/�P��NԊ/��VT-R����ȓr��e�A�D�D�V�� n�21�츆�oN��R���NND�:�G�2ߒ��ȓ$�(5��F��U�,Hwg֧| ��ȓX�P5��b]<hMP�S�8SD݄�=�����U�U�r�ӵ��-�����Ԡ�>@u e3�Я "쁄ȓ/%0�h#�F�!��Ĳri�*8���I��"d,B%K���FǕ�P�*p�ȓ!fn�0��0�4�0�W����H�|��cX.'�<�H&�_������>US��K�\����R�K����H�=�$l�)���`F�M�U3��ȓ0L�'�>A���W�D�T�2��ȓAF�QCi[�v(������ņ�[4p8Q�ڈH�xh� !Q.�:��ȓ�*T8�͌�H�4X�!� b-��5o�8ӫ�X�]�U�51&H��	�|���=C�L�pGΔ	bڠ�ȓs��8��'��`�Z"�DI�]�ȓ��}C�ܼ| N`����E���ȓnF �J��,9�LP QGR�p�����v�J��ʄ�y����p� ��TW���5�b��2v�/K�R�@�"O�lc�[�H�MҥOE�J�̼�`"O�)�d��$I�ҙ�a�٭8`z�U"O���fEC�$E:A-E:>�4!�w"O��vG�rD���J�*R���f"OZ1 G+ZaJ�K��C(?X�+7"O�%�A�,��X+Gg"7U��b1"O�Y�V�.;@^ ��f�02�Jdɤ"OV���lC]e��1��X�u�,�q"O���bCD?_$�p�WJ��C��(��"Ox��fʞ�.;b)�V�Y!*���"O�m�$�ƖK�6XZ1H�"���!�"O�� ��J!A�&�qŇA-=�� ��"OŠ�щs�h���e?[�b��"O�)hSl;K�9a�a�[�<��G"O4��R�"ǼL�Bϗ�>��"O@�!AfB�d�n���,k�jl{7"O����JC6J�^�ǁ�9�E�""O� P��nGP'|��2��_�6�D"O���#'T�%�� ��dXs�O=�Bm	�!���O�>(E�
$C�����Ě7;�(��3D�xfK�h�����x����<Y2�Wp�U��0<i������e^�8��I�ƕpX����ͪc(����,z0p,k��2
Lb��Ų�'M@�!���H[��`g&�B�ȍ�	]IJ��m[�K]��@G!��_�-�$��H� � ��C�4S�!�䊕c�� ��	������UA�'��P!�k�!<�y	`
]�Z�9�)�矨KX����ӂ�n���q*z|!��2�V�҅�P�h�8�K�@��1)J�-_mUY�����`0�<���b�@�-%�m�C�@Vci)�e1��2�B���+3����hՉ �����Ȁ�.�m�f/�/���2Ŏ(+��
��v�Xhw��8�ddb�bZ}�V��ɅwŌ���.�&(�����]�, � N�w9���@Et�da�#=C @t���g�~�;T���!�]�d�ޭ���L�Р��`�>h��Yaf�\�I�d��(��rTj�4���S�.�8j�ʒP���	�l���X��@�zz֡:#�XM�㞘�rl	�f����{�i�{�҉`��5b�(�٧�Q��������M�f�S�;�`�cBuɺd����"<	S��j�����\�J�Q�'A$F�����Z�N+ȓO���c Z�J#��Q �$}PRt-�=8�հ$�F�Sw��iT&Ɨn(BMx$��.C�~D%��[��� [�-�V��H?y���w.|h������AL�'	z0 Qٸ
g�����t2�˄�ފ����B|��8��y��F2��)a�N�U|t5�t�M��~�		s����k��!l���ӌi�"�I�I��A�K2dȈf`�+0E�d�t�@�9Nܙt#f>�:��I4M�4��aH6fĈv��-2Lh�a��E05��>GJ�z���$�1h	>, ~�-xn-��?I��ˁ~���e h.}k��ͺOO��e���"N��F�g�ڠۤd�![�&tIpb�m"}c���:LH��%N�qf�51<��ӂB�d���P��z(8dBc�.-\	�)O���	6������ow>T"G�����(/7Wݲ�r����6i`��ɥA<`c�m�����̓�'ʘ���6T٠�"QmТ�&qH�<O��7p��A@6;��aKN�&K8��30' �NP��虴`�d��4x�@��� mu�Ο�nM�IF���W�N�`������PnZ� 5�Œ	�.���'���$��\�65���V�ND�; @�kmXM�\�z�� �	��7ӎрt
�� Mbh�p]�|z#͘I�D��D�� �%C�� 92��!�R�ȿ����g�R��	oZ�GW.���?V+���JU;dl�cTU������(P抅���n �Y�՝/�@Dj���5J���ٶ`�X�5K���& �`H��ҩD%�`H����h h�s�E�V|�����ąu�6�E��9�J�P��_jy�CT�Q_�Xs�#Ԝ{�n�*a��'޺y7R@���Z��y)��M�Uq乫��&( >I�(��Q}�@hu�;���x$r��T�?�]��mÇĘ!L��Q��^47"^��A!7xA�1�D�����A�)��<�â	0뀴�Co�;A�-[��M"=+� !�	8;�"�+$��3$�0��'芨����G����1dmΨ��C7O���B�a�\?yCƍ�o�Y��ǖP�b�P��'�	\�<��E��o�����iR0!��oZ�9A�@m�1�*ejf��2|�tؓ�J g�Q�O6X���Iɤ9��A�5���Y�,~&㔣޼��Éy�Þ=�
����#-��Q�B'�2K5�����dz�b^�4A�GB�z�<�0���C(���o3��ŃE�Z,�+ߧ)�J�>��R���Z幱�1R�Ҽ�A�?,�"#��Tw4s�N�(~Kʕt��hdj��9��2��y��ѻЮ�$��|ƒ�b�@N��?!!�jKt��G9}���D&Y, q��W�k^�b��T<G�PQ�!�#�`��^�j��U>C�J��&�t��v��FP�+��Of�0��
_	�Sf�*\��YRw�>��LT�c�֝V���$�U�K�A��n��d�&��@ HK����<�"f,ӏ�4��K�|�u�C���j~�bC�� �p:	ށdv�㞘�4o 38ˊAhs#י�d, V��M�8�c,��324]�c ӊc����P밬�p-R;:�(�ؔ�˅�J
xJ����\)Ҏ��M��Xค�g���e֡j�	/�M�7k�
�Bq�M9R"���wp�5�����] �E"b���'O��H6�N�Yu��W�fԩ)5��c��̉e'�d"����UO��`F��\����&
l��A��'VqY�H�p;�)�AΝ�)�	�@ð���݀��ʠ]5�eq�� ��B��K)-�����Z�L(��.�,A����r逝Y<�I��D��`)~M�GJv�L�+�K�8�1OH���=�ެS6�5r��)7�?��x�s)�:f$��c�N^Vq����_$a���2f�>3���IU'
IX������Rs٨c��A��hQ%썎z���C�Ǒ9��YD(Q�����ɟ<T|��Ӏ�E��lAumޥ" �'.��x#���d��H %+&D�""#��w��Yed

i�¸B'�@#%<X�wlћU@�����+u^*rÔ�r��1�$�j�̘���M� �4?�ii@��]� 9ksЅ�jA����D�х�36Q�0[?1�U�,@�����Z��р���0xPY���v�0�2b��<=@G�':a�q9���$[R��A`��HOB�{ƨڠ3Dfxc��3�!��A9g��	2cF�7��=�0!� _V�#f(Z�0@p\##�0�5�%E�c��d �.��h	LQ��q��!�b
�v�V��Ơ�u�'��ya�F�9^��ka%�sㆀ�0��Vڴ�%ѰZ�x���`$Q��Y %�ů�_��4D.��)#K�b��=�p�ܑ1�TX �^.5@�ZAG�]��y9Ę|RE_��WŢ"���g��^�a�ץj[=B!8,D��U�]���T�a�P&!p���d�^�����/O��Uj2�ƛ,F��J�=��@�Q�"b��r�� ��S��Pm��x�#VQ�0�0*]?e�&�%<8r�!�oB���cрДl��l�S�V�S�<� Jܽ8���-t���3bB�6�dX��n^�'�=!"�t�@N�q	4�Ȇ�5�l
�XEi�l��Tb "�~1��(�S��i����"I*�5H�V���x�	ڴh�1����Ob	�0hA�T�&��ND1H���J� o�^mi7�R�2�N�t(=�I���
 `�i�FA	�Ɠ�4℁k���[&��u̘���T(Q�����%�/XÀ)SQm�� ̎�U8�E�X���th�Y�Ĭ�0%h��~�^�CG+Z�0}����x��5i�I$�����o	r�|i��G��L!J��1��СC�<X�L�C�,_'�m��4;j��gkX)<�t���kĹIv��!��{����>X�D�I7� ��c*38TA�!��1�eè<<���Xs�@1��`#Z2���
��64|	���8��.�"pt�x&��� 
�2�Q�W+�;���Ч��J��1#��>��YҘ���KF����͕-���YP�ɘn�t,��_��bֆ �#i��⑤G?:f���R�����ݱ�`H��&�Kd,�r�ӧİ<��	͏9��tpUJ��I�Ε[f \"0�0DP̒<=w<��!nͼy�)��BB�8�3��ȋ��#1�*|(��'q6����?~�B�))j�P�BزF}�X��D�d��'��d���Z����s����@L,��.�������Q(`@t�zx���L�sd��V@]�MS��,w����	�x���PH_���J'ϙX̓�T#��'2����r�F=  K77�fIB�ʂ$:<�rǪ� �D���%7�� XB��q�H!��~)V��ਚ
R�F4��+°7�h��Ǣ�	���x�NE�n�$��I/��Ę� �%3
6Y��f�$I���Ɍ	6���$�J3�����Yȇ�F� ��,�M������`��\�v3��Ueσ/�ɐ�.AN��Ժ�gaA��qj ��12�Դ��ݱy�m� �ŷO�T$;�N�*�	�G���^@�4�а�`�O0a���ڥR"��i�.QPf]��_��Q�0�I�} qO*|��D�?Ld�Ғ�Ì�f���8NV�`d��*�4s���Y�����%,RL8��@j���'�L!Ѡ�*�����<D,qO�d�R �}SdI�&l>=he�6/ �p���6F��h���S�Wu�`�� Yf<8��Q�"�l�����ݼc�G?�A�z�Y��Y�e����C�4�9dʇU�MJ��/O����LP-o200���B��_�|��a�=�@��{�NYx�����C��0O^(�h��� �3]�8� ��U�M7��:��
�8��a������0��˞������rH�e�a��S���!�iT�8�v�H�k3<p6ʑ? ��G��n����wzL�m_�R�\��fb.XƖɱ	�XĒũ�灅--&��ǨS�U�Ɛ�CʰW�\Y!�Ӊy�*
��9?7�Kաɔ%4���� Q�ʄ�cJ0V�Da�'"^���"��4d���>~���{��$^���E{��O��W�=hl�1���9e \[P@�h\���1d>�cfA�D�@�ƴs��9&ႁ:b|G|�"�`�n��c+��fV�� ͖�!)�iN�:��TQ!T��vJ�]a�j��+͖cB��pm�##.�EXV*R�z�TlYlM2)�4�8��)�6�7�ŗ4��}�ô'b�0ȡe��4�� j�# `+��K�_�m��mS���Tab5$j�����(ɋ�*�7�yg�ۋs�Y�$̎�Zd���OQ�0>�kL|��(`d�D�~$t�v��ڥ� �kXrt���h$���A���c�ʍ)�Z����*\�c�a��>ޤȀB�'^��C��ęH9��`�N:���Ey(
(V��5��M3��R��O�������[�WA<Y��.��T/ ��hVL�I_쑣!l�	&�1J���N$����y�'���%�	{8LX��F@��~��Y���WcŦod���M�w�ؐumшx0Xt�&恘	�j4i.H\��e���!WNU�e#��ܰ��C(�4�^�	R�'V!q�C�-]B�lSU��?PMȢ�Б7&���D��P���!U-^ ش\�����J@z ��05��X`R�V<(� �b&i�l��c�'y�tSLV�%s6AT�(dv|Uc�&x�^)3�M� �BVg��uQ�e�ɔ�Ԋp��*a}fa���{�X=0�RGA�hT$H��� �������O^}Ѣ�π!ڰd�g�'H��ˁ�T�+
�8`bM\�O�ꅐ��BELt!*��4I����M:�DD֣v�pm�4@ݎI���zƯ�m�|T�6�ȝ1,T���@�f� �v��'lٞ�Y�B�:i��:�O�o�rt�7'@�dP����(Z^؈�\�haj`yv%�?����	*V��Isf
�` ��+2� ���i�c�K�m>��rIR�|�¤�6��X��c�$�L�5���Y�U~�@�� �$Gw���3�'�����	~n� �*z�~����A�Opt<2�`�d��G��	���A	,A�^�ˇ��Y��CQ���dr��(*�%��Ÿ_b�\'� �I$F(�� �&/�@9�@gȷq9���$Ӻ\�e����!İ�&��\�����9x^Z�Z�A��l?6���M �.*�G}��.:��5���+�c���C!��
�?��q!��ua���đ>���q��*� [��	N�
_�qx��,��A`��@�q1�!�L���BiJ�"�,O�y�ԁZVmʔ�&Z�-����YM��&�+*c���2IH��U�d�Rk���F�/��,Kq>�j�!a�W�ƜQ�Ɣ��ͪ�S��
C�APmy������-9!�}�͝C����h^� ��[̄�gs��9KJ!x��C���`�F\B��E��8�Gȟ��
�f�O���O�n���q��gr�,3�L������r��%��f�+�����^��@��^�?a���w�΋R�z�al\2a��
�ɖ8倠`�놞U���k�^���K�pEZ��E�j��|��#�̏OW��ʂL�nׄ���')�Ԩ�e�./M���M�{^@�!2��ٚ�MjЎՠ�'$%����E>oJPq��m=����ߧ6P�;�D�u~➘PS�@>5>\��/��4�8���	5ߌ� � �8N:,���O�Y5̚�I�5b9�#!\������@�x֜VZ X��0�?=<l���"+�ti��̾�qq�͔�qb|�KE*�>�-K�j���{3��(VHq߄ݲ,�&�Y������0I\HBb�C���!%�I�^��*�D@�%'�p T���SӐh�%O�(sLx�"�G���q�M$X����`�ఒ��­ F����i���@W��)=�&�Pd��/���k��r���� !	�D)��4Y�v���生�� B�ǥ�	+�h����W���K|_v���!K� \�1�Kأ=�V �GH̓<�\<�E"P����F�$_�
�dԷr�^r���+;m�A�U ^�gEXA[�� U����s�Z&]��P����Ԥ9�
Q�C�D'8��`CWwo�M��<,D`���$�>*TD�C��3�`�YǦ��<�U�7J�<�%��&Œ��:�0�c��J2L��`S�
{Ҹ���?R��!aD��>�Ҡ:�:�K�h�ݒux����%I:�j�F��%�8qRIձ?���`�l�*�	�A�!�V-#`��~B�Գ:K�uO81�W��]�0XT����\gD� z?L�`E��F��ّ0��tL0%�'cX�<p$�i�L��֎[[�M`�"��Fd^!�,��o�����A$LDT�D��?	�VȲ�M�A���*��QEb�'�/l�ąQ�se�0� ~��͐rfA�EV��GQ�Fh�=��Hʆ!:hA�@M J쑭�`����FP�X� xS��za��Y�j�c5��I6�x,�7fg����F	U�LȒMV8x�
��$�ܙK���;�]�)�v��7-����'��A+��qb&��t�`�U/_�4=��y��uL���EN�;��YS��v��@�˨[������u���&&�-�rʖy���D'e�09pF��0`|`��U$["��I/`�����ȶEY�����R$���B���-���'8#�$�e�d�p���!@�x���#Xa�q��3��	*4�W��H�V�	'��)��E�?OR1q���xڴ��;p��(#���yӱ����q��
�"S��Ph Ӎ�9rȓ-a/0��q�A:�Ȁ�L!�6�3�(�S��J�}�p�I��DБ��{?A�o�h��h�&�"��'����-L�,�3�*wZ����$k-N��q���2�D<a�%<lO�=I�	$f �;5�*|<QSd�`Xe��;Q���jH>��;P���b����EW�O� 8�0���mK�8���4F��ڼ9�#`��fF�V��`	[4��r҉L�;��8��&o*���ø7/⠒j�0��і'�ڴ��*�(|2��OQ>��p�^dW(,��ĨC��}Q�B2D�+�M� 	,h҆�l|Yp�1�ɀ6�(���'�!��8l	�qҠd��^���
�'�����O p���0�^U����'(*���E��K�-��LA8O����'�xt�c�׏ (���Ǒl�z �
�'Ja1��8>k.]ؖ���ۢ�X
�'ivQxc-��̛`FV�n0�	�'��Jr��i¨˹LZ�L7�yR�^a���;���|Ұ�Y��yRh��^�r�6+
\7t�!�-в�y�I��B�b�@�Q/�)�@EF��y�*��+�)��M0E]��)�e���y2�
�O�T��u��0���l¶�y���6k`���0:����y"ͅ�L���d�P�-�j�����ȓ��m���Ʌ肤i�D°:_���:���!'T�&4h)�N*)z�8��s�� �ǜ��#���WH�����){����}B�����'p��`�ȓq�X��C��<��C�ov���s�����F�71#��s�Iğ�4���o�N� �e+p��#���{����=\�	���ԜL�]�Ð~K@�ȓ#{6�ʑ�M�:>@�C�g�����0H�<��	� (h����덄zN�u�ȓk�H�a'd�<f��N�!�>���	P�a۵��8��m�Hw�NY�׍�������`��ĵ �O��@��#���'P�����Ab8F���[�`{ �P��ʦ��h�C�x#�O����6��o�8�P1��;x�n��LI�����T�+�r��<�a�4�sը�z�GD1bC��A�X�xt9G�
+7�'�a����`����3�I�Y�V���_� ���v�>1�4�O�O�j�	w%�7|�4Y���c����J<�0�?�S�'j�j���K�J�R�wl*{�'c�PFy��iHj�*H���l&L�3CK�k.�VE��ȟ,ȡp�O)I�2��.�L��x���
�����3}��!� �I�`��˒[����}�p��%�D0���<�(��9Za��.Њ
�Z���٪�Ƅ�|� ���k�X�P��-:lqO��V�[f�+���vE�=+I��un�=`Ĺ� ���oV��S�O4�� �(�P8����M��0EQS�I�B�0Y	���d���s��i%��ٷ��(�>�`�#Iy�eX��p��m��,t ��/��O�'%ɢ5,MxP�m ���Y�}" �`~a���+� [��R�5����&��S�1��6OR�Z�.2�g�? �	��FS7w>BT�T�u�*��O���'m�O�Su�8]��ie�
3�$��(�/�����OV��M<E�D�D��xV.٢/W�TH��B7�y��A�$nha�4�S1M����b��$w���D7^2:O�<�4�zc�b>M�"#A�u�|1���!/��"R�5?id+d��p�y��)�:0���a���6r#ʹs�mT�7���Mޟh+'��S.O2�I�h1#0�L�ƙ�B$V�����˓�y
çzĬ���C��F�C1B2DC��W�O?� ��$��?]�d͟��)�?�DǮi����� �x��1{��0�!�D�3e>z�YЯѧx���I�/M�!�$�!p��!,������!�ɮ��0����I�n!�(�i!򄎫A
��9'�T������$!��إpM��"�/ ��B�"|!�F3>\^�i���#F�0yTC\,�!�$س"<�+�Kܕ̦xR�L	�0�!�$��r9R,x��ܪ&� �b�m�8q�!��zfr�b�G�<A��x0lV�!�dZJ,���.���%ք/!�dW�eQ��+��e ������Z�!��FF�vC�;[��Ac�3mx!�D������2�"S�ӵ�D�-�!�D�-��Ԓ-@2j����K�mQ!�d̏+�Δ���D�o�Fia�n�-OO!�ޮp�ȉ�̉=��d� MK�Q!�$ �	S���f!!�F�Wf�Qz!�D	�k5�S�Ԃi~@i�U�ͫq!�$H7!a�<�AŞ�L�Q�nU<xc!��9�\*@���qP���A�!�ĉ%,��d$M�	���6<�!�O�H6��A�/J�L6C�σ=~h!�d��O�bL��!�n�K�v��t��'w�5�AL�zxt�'gB���	�'��r�ƦQ3V�Ń;k��)��'�q�pJ�}/y�3d��l�$��'($����	�i|>)���ٶMd�U��'�lP���b$�(n�BF���'�1� �+TѸ�� h��|���'��H�s�C�df*�@��^��t��
�'C��� �H�EJrG'U� n�)�
�'N|RF(��~���F���'�ֱ�'��,�Q
)}H�V�Uht���
�'Rt���K�H�H�Ћ[~�Q��'
����Y,J���ӌ� N2����'�`�'�#x��9:�+% b��	�'�LI#uLR'e��L��)�%���	�'�"����8�V�&S$���:�'��KW7W,`,���u�]"�'�ȴ��GIBjVG��PV�Y��'�0D����$ JH���GܜIB�'��m�#bZ	s̺A�t��(�f�+�'�v�0��>[P�9��#:��)�'��U{Q�X�~0��;��ݰHn\P��'H�(�`�@�Q]\��lV(@ZR���'���s�H�8��92�O�8*ϒl��'��(��î\�P8#@d҆�"����U�MO�k�L�G�Y70����?D�h; Šw�a�6�(L,T$>D���TʛV�j9�T�՛=�,�Vd=D�h���H�$� )֕-,����d/D���'��I6F�;T!�e&-p�n/D����E�,�a@�(_�TP$��% D�����ߦe����e�;ܕ��?D�� �2N��0���FO�����>D�� ��c7C2=^2����g���
�"O�UyrC�qx8!��F^��e��"O49"�$����OW�x��"O��2#��!`��ဘ�Hy��9�"Om��̘&d?L����w$���"O��Sc�
9��@ӧ���S�"O0�b$��J��a�V���5p� ��"O����?Ttss��&8謀6"O��r4� �d�$Ч���M�I��"OJD�գyL~4�v'��.:" @�"O����,[V"���ĎD^�S"O�P[7�S�cR �g�<x��T"O2����׸x��Z3U$���"O*��# 5P`( ㍐3�=��"Ob�H7J_�WDx���@k�H�<Ap�ܢ\��YA2`
kP�xI�&D�<��A�_��O�L��$N_y�<avAC�cEĐ���W>7��4 �ŏq�<�s�Y4�6A��eV�]�EqB��n�<�F@CS�̡�ViՁf�bYYuiKr�<��*ǣ,ь��̏�3vx���o�<�����wo���4kM��}b���l�<�ŉS)~!Pʶ��\��8�Ch�s�<��aѥo����D��:�,=�w��x�<eeW�Q�t���Ju�"M O�h�<�Eb~VՑ�� PF x@"KY�<��bHm�~���һ�HtH� �N�<	 @L�Bf�X"���
T\�æ�C�<ƤH
h��H��l̄N)p��!D��PG@4r6�\�U��F�~��@!D�tQR +c�����^�D4c � D���u/��$�S�	�r$�:�4D����È,�JD2cʅ'�I��-D��#�K�8^R��k�IǇ���2�G(D�����@u�*$�Qr�%�e$D�d �f� ^�10�aQ,g~n�	Y�!�ۘD�T��#K�OF��g�M!!��ā
�|�����|O������3!�d�c�1�����iH��XU �RF!�DJ����0�C[��9��.��^A!�!>�.Es�eƱ![��@�mJ�q�!��� DH���˔AO�r���!�ݱD�V��'DQ��Y�Lĵ�!��]*NI��5/�̢��5=�!�ē5hZP�4O���faވ�!�dϋ)Ը�77�I"�#P!��=z����BL�3V��R��!�D �X���J��!5~�b2�)Ai!�d�y~�e�A
N��q���ʿV�!�$X�_>�8��F�����T.�!�D	"j��Po@�B����f��!�ąaK>1&� g^�:D�#�!�č7-��]{0��R\�5h����!�dC��&�y�����%�)���!�D�;SD!����c��8���B{�!��;r�����&��k����A>N!����K�7vP3Waֽ:E!��,U���s���0r�&^�O2!��-\�|z���0{�r��Ug�� *!��5z�P��A2~�R<�0@)P!��@�CE���EN�	I�(�j1m�B!�d�J���3i��\�Y1,M�G!�d�t�v(p篎�uݸ�r��&,�!�A�7A��f� ���ȗG !��  ��fo�^UH���\j'"Oк�c��Sܤ�s)A��4܀�"O"\�BBד^�bQZ�h	�\ך�i�"O\��dMD8����H3o�xQ!"O�)�hHu,�"�Ƚf�$%2S"O����H�v��bÅ"g�x�r�"O�< e��c@�P�Ď�t����d"O��b'�&Q
�ԃ�oӘ6�0p"O�<Z�iY]��ه���h'�L��"Oxd�B%ϩ@���B�'%��c�"O<S7�<�"=C��E�r�,4q"O �����"_���*pb-1��y�"O8Z'IS{6�!��x�J�s�"Oހ �!�h��xs�/ǬǾ���"O�Ti4��X���4P�x%�7"O0��U$B
X�� &Ώ}0P��b"OzDU� �cxP���u"�(�"O�1 $S� �M���S�`Az"O��W�ܻh��ҋ׵H�H�"O��q�C;�~-����$t�Z(�"O�L�r�ˌ\?Ld�C釈����v"O�l{FV$k ���͉�T��	��"O�4��AD�0쨡�4������B"OZ� E�8H�@�Ѫ�W�HEa7"Oh��# �/�V���jCU�}aq"O�D�5c^[r
|�Jˊv��@�"OxI�w�P2{�б@���cV9��"O�4C�L�m>h�X㧟%&W���d"O�����C�eTXx�G�(��y�p"O�����X�?��)�t��1O�J���x����*���P�1I����ȓeDf]SB-^e�d���q'^H�ȓX�Ґ�VF�%y�z���E�'v���HJ���e�G��,�D�_�~B���^\cf��x`�A��%Cr��ȓV7tH1��YL�ZY��%@��-�ȓ"��!�D�T�4j��J&MR =�B�ȓ:��q�e�u`mJ�/��o��5�:�+e���*����D}+tm����3���]�>} 3�N��4��>b~��e�ٱ)�P�����M�`D�ȓx�f���lsP��cž@�0���|�@��V�ߊZi�j���D�xĆ�w(��5Lׇ;���k�f٩38^ �ȓKJH��`��ʦ䚗m��-2��ȓ
�+��
�. I�!��z�"O湛T��/0��-z��,7���"O��h�.��e��][�hM>�Qse"O4��!H��n3Z4��f�� ��Չt"O�2���kf���dR;M�d�У"O�}�KM�!�D��۫`����"O���PIW*J��I�hȳ9l����"O ��f�	�����/e�a+�"OVyK���9�ܵ�B�Km�~�H"O6��/
�,\L���E0'�`5�6"OMS�DV)�ʸ[goF�*�xhr�"O6��XB4L��H�tᐌ�(N#�yB�2zR="�肄#��uz�L�9�y�L��E2VKޥ0�� {���2�yh�WĪL����2,*�sBK �y�h��h���B�</`&<���!�ykW�.U��L& �F��5F�%�yr�6���B
�h�<�r)��y!�C� ��(X��C�ɵ�y
� ��Wk_!�
ҊR�:�� #"O*0˶�ơ,=ZIJ3J�A. �"O�@
�Ǹ*6��a$dZ.U��;�"O�)��9!���2hT�8dPV"O�|���F��Jh𑧀#2�0��"OV�i�i�(W�%�D�ׇB�@Q"OƵC���"$��|� �?���7"OQ�Q�Ӛ)��Uz���7���J�"On����ӊ,��a3A�	 }�,P�"O���d�T�IgH=�sD�(׼���"O�!����`s"��#�X(Y	�"O�r�.F:d�
L1�\2SW����"O^L�wL�t�x0�T}R�Q"OR�   ��   )  �  ?  �  �*  �6  �A  �I  ]U  sa  �g  n  bt  �z  �  *�  m�  ��  ��  7�  z�  ��   �  C�  ��  ��  V�  �  ��  ��  ��  3�  �
 � �$ m, �2 �8 i<  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��Y�1/l	aCڷUClM��%ɘ��n8UZ�&]�KR�P��,%T��<A����!Ez��F��\���i�L�/Bl!�S�t�3�a[��~��	9"O��"��IvH�	��EL6j�"�"O�aY���VAv,84jٟ.��"Or�{��+Q���A	L}>q�e����D,��ʆJ��t(T��43 �B%�!��/@��*e��-�tF�Q���hO񟶙��$ڸj7�7�B�Z�X�,D�|�7�g�Z���\� �~���|\�S����M�o�|P�L�"��uȨ�Z�'�L �r�ϓR�<H��Q/_��e���$*<O249��G�/{@ыR�%2��Se�'F�,���s��P5�!�s��5E~���b��ex���*x��ᐦO��HO�����`h%���a���
T�V"O��X"�@57�R�6#�^vʸ��"O0d�7@ 4i�8![���Z[�݊�"OaZ��R�,�"�;��T�xD�9X�"O�#�EMd@R�+F
]�� *��'Z�̈́	�dlqi۹&�ͻ���z���$=�����"	t1�.r��'�a}�c'
�ǓE�T�8c��Ұ<)W�>�O�����mF���& q��I!���F{���(aDQ�p�"Ǵ���-�2�1O��̓�4@�2�3�  ��B�G�ecʜ�R�.���"Od���/Ƽ2�K�Ȗ6nƲ��3�O�=E�TV*�\�b�Z,�T�k �N��y�J�v 
8��&�b��,��y2�
/B�R�x�k��1����jD���>��O~l��M�Vk��8ċ�4$��1�"O����B�)G�"8ȡ*�8U(Aӵ"O�l�E+Y�U>�48�Jӡ/�����"O�-r@�C�\ ����$z�t�R1"O�����'6��]?Y��R"O��³C�&���	¨|����"O^�{��G�
�d{�"hh *O�M�5g¤%�-ۃʗ1)}2�H�'��Xp-�� �\t��m�kJ���'ڴ���"F�<�b��$����'Hٲt�S#����!�
k�ܒ�8.*�6ڰJ獀�6vP9I4e�'@���m�|yZC�%x]��N�����Dz��~���IX�Չ��^k0NXǎUd�<���F'W1�%I O��՛"�Ҧ?�"=E��D��I���5yb �`%U;S�؝��B�z;�Hņc�6�����d�,T�'_a~���T_���+��X�<�j��L��?a����8������(c��BS�9+q�|��]fI�����ht4tZ$
v�X0�'�a~���[K� �	��C����᠂��y�A �f�\�iS�n�*����y��K"��0ՙj2�䫓bR��hO%��)��8�4={�I	
kƞ�v`[:*�!��·|&�!B��� "�� �ռ7�!�J�`�����<�R����t�!�A�_�t,��-�'!��;���|�!�dӗg"%pEhތ�2���jȓ�!�ɲDEz���$��o�ӉĔ=r��x�㉳	xR���7`�bAj�O��
��dh����i˹2s
��)���&#D�`X0�Db�����ᗘm-z�j��?D���"*��Ae̍�C׺r�0�鱤(D�\E�Ґ +��)i����㤟�D{���H%��1� @Yh&�A� =!�$^�yUVxi�V9eǒ�Sr/ފ6�Ѱ>�a!�[}���U����k��A����'g���r�Np��d�{�l�X�'���:�/��{()q�R�v����v��E{�'99�\B���T�]h� ��z}
���9�TPh��/f��PL.s?6ɒ��9$�t[D��
K�,���(�X�Т�#LO\�@�"J�O	<�PSe$*^���a5D���Q$_%&|غ�)�5.�;�G4D�d�Ǝ�D�Ea��k�d�)�O1D���$ޠ�����H<P8�H�ƭ<�$�:�S�O8*���~'L6��*��i�"O�$�LUaa�q�ƦN8eLy��$^�<Y�~�R�� �-I��{Ώ�"`���	J�	l�@b�j%N�

��n@�8#�'k��4	ҏu8Ԥ�TCֶ6�L��˓�(O��#�1d�����BS`!1"O��@���.�HU�1GR�eEޙ��>��)>�S�'~|mc��ǃ>@>m1��@�]Td�ȓs�\��Eő�2��Ɇ���̇ȓDz�8`�Z�(�8=���B7�0�ȓw�.��!�U$��Z4E�}DD܄�`�0��2Þ0�쉁ōT�(�ȓ' @����	$Vd�T��	�v���S�? B!(d�ʑ�xǁ��W<�D�xb(/���%��1��[&H�8a�"N>4�F���i?�p�ҒR7�m`�
VUԵ�EK�<���+���p.C[qK+���D_�Q��7�eq���H�)�ȓR@Q0���*���� 6D���ȓN��U�@�ƈu[Q1��ο"�:%��@��Ϟ�D�fq�(�or�ȓL 0�	AS�8�DI�F~��ȓ;����g�ӱM��0�i��;�m��}�|��GMQ5
�-X���&T�(��n�Z��@U�]d=���д��\�ȓ_��e���΅S��!��.'n�@��	c}���.A	��0�!P���z@
��M����s���C��5!�m���	 h	�"OjiBCN��l��B�]�!�f�)�R�̅�	,��"�j
�>Q�P�����~V2B�IKO�
�F^�%v��%ƅ�>SDB�ɞ|��D�g���d`�h��+B�I6
P�S5�(��!h���\��B��ӟ��'L��$(J���-܅+/��P /*ʓǰ<�� �Tx@�1c�D�+ƭk�'g�I�h��h��Ͷ	F�B���(�MD"O�}��%�, ���U����{I�<I����b׌ѓ�"ڰatz��[��C�	5�]I ��D��=� ��;�V�=yÓR����G��<��M�`,(�����?7E	2(�V�ì{��=��Y�<�A�We��}�֪��5��=(�ZT�<aWob��r�LN�3����FS�<yfɝ7�*�:��Ͷt �h$Rt�<���؜9�Q��	�5��9b)�o�<1A+U�����F��!шP��j�n�<�U!�2���boӱuH�]a׭	g�<��n�9���I��-����/_�<		�7.�����f5�dx# Yv�<�w�
�������*� 8G�o�<I�i	#�Y�^�,R(YQ�"�E�<�t��!Dk��X%����t����y�<Y3&H|�6p��i�D�0@��r�<QT	�Z��r��+�0%!!Ak�<��&G�k����� ��'�	h�<i��$`�zH��b"x6�Qc�k�<�a�]T�t�tMU4R0�a��Ap�<��E�&F�����
8`���u�<i�I҅D�����e�!21,�Q5��n�<�GN<����F��_��#��a�<a�c�(��q)��\1JM�Qx��^^�<�E�|����挭.�&�P�Ht�<9�%9\����$G���q�p�<�r��1��u����R5�ea�<Q�щh���Z%K��2��MD-TZ�<)F��~��Tc�#�m	�}��V�<�W
�w^콂 ���d́'EIN�<i��ع"zB��@�cs�:��H�<�WMӟk`"-�S��j��
�Z�<�V��(gDT��@�=u�B}��b�W�<��΢<˜�����`2Q��}�<13埦ZN`��N/D޸�p�O{�<闇_�F��,�o�vG��R��B�<��2u��8#�E�_K���"E�D�<�Wʄ���-I�ਂ�&G�(B��1"&~H'\�W9��!���QBC�!Kz�$��,L��,!'d˰ �C�)� �����E\�k!��$SH�"OtM��imƴ"@N7 OV��v"O�٪��`�;r�[93�@�"Oܔ
5#ԙg���W%O/\��@"O� �tl@�~r XפM>$�$���'�2�'r��'2��'KB�'6�'�@�A�E(uYT�+���(22 �!�'�B�'���'pB�'�'8"�'�H�"�Ȃ�V ղp	�A�\�r��'���'���'��'	r���isB�	ߌ5j���F����o����O���OJ��O�$�O��$�O^����Oq	aP㚂��!CcA��$���O����O��D�O���O��$�O�d�s-J(�w ߲���+	"��D�O��$�O>���O$�D�O���O�dJi�\q2P��)������{�V���O����O����OD��O��D�OB���<~�ܻ��� iԙ� �7���O,���Ol�$�O���O����O��m�Z�[K\"� � ��8dZ����Or�$�O���O��D�O����O��_�Q��8l��5�i���@�����O����O���O����O����O��d_��8���M8�����'ɘ�d�O��d�OD�d�OL�D�O����O�����܉��U</b��k�;8����Ob��O����O��D�O��D�O���0+��e8��
 ��s'�A�����MK���?Q��?���?�׿i���'Z����Cʗp�~S���;�K����������$[��qA�	1 0
�Ěs?='D0Y�-)?�E�i��O�9O�D߇o�V��� �a��8Rt# -t���O^)ا
o�����Td���O�"�cӬؘ~τ55��7*�mc�y"�'+�	s�O�6L3��4'g���'��+xI��N`� �#��>��1�MϻI���u��<O�ܸ�Jt� ����?Y�'��)擽0y��o��<iΈ�R��U�p&įN����A��<I�'f@��hO��O�i�FU3�
�a��ȱ+$��#�;OV���XԛV�۞ט'��=�R��;QɁ���<0����	f}R�'�;O4�9�$��D�25pyp�	�	��d�' �h�>00]����H���X�4�'H�� R)��T745a�Kڒw�x�T�ؔ'���9O�Yʓg��9���[�DU a�:�Ӗ<O0-o1%������4�L�:ńL�v�^��d�;���#=OH���O��dÀk�b7�1?Q�O���eF޴�D��:	%�Ā$C�2ah���CC�r�l곤C�}&�|�F��T$4K�+ĭ$R�9�A�8u@�8+�@D8t2��镤��*#������d3(����D�d=�x���%u�����-@Z$��� �a:�
"ݓy	ZI��i��hf+��S����U�b��{DТ;����V)&sŹ�OK�y\,}��ݥ9�E�sDV����14�f�����jj4�� ��}���H�OVriK�O>bb
ȸ�,���$���^2�TCg%��Q���YqJ�[n��d��
�h����O�s��@22�	OgTu1ì�'2<�Rg@�|���'g�'��`8?)�+��x��uyw�F�g4��2!V٦a�	��ԅ�����	ßH���?����]�D�G�zT��ڒ�b����u�i����jӊ���Ox�D��fQ%���,
1e�����F���	��� 1�4%Q�4v�(�z*O�d�O���d�O�H���U")�J�����.Ly�I��ܦ)�	�X���(!�՚K<ͧ�?���E��}s��U�n�E:��N�����V�p�I�@"�?�I� ���<i�
����K��5�$�r���MK��uz����x�O�ғ|Zwi����� b�&���A΁M ��O�A���O,���O�R)�i ɝ-}^���M�_�P�ڀ쐚r1�'���'��U����֟H�Sk��7�.�h�6���'J�\66c�p���(��ay�"��YDt�S* �����H��p�G��>n��?	��?�)O
��O���'P?�Ȏ$:jSFإ)VX��u�>���?a���d��e+'>�C阌;Q���ȇVֆ�i$���M���?�(O�D�ON=��I�"';DI�0��;@ubw����f�',�Q�h�$G�)�ħ�?��� A�kn��Y�+]U<*��q
ئm�'�B�'x[��Iꟛd�l]��G�(�b""� �M)O�D�P��Ӧ��������*1�'��ՠ�+�/:�&I�m� ��4�?Y�j\��(O�S�?Oҭ�4E�0(�jj��Z9β��P�i�hf�w��$�O(������&��ӭ)�ƌI�lԀq�B�$�ǡ�<���40��=(O�$�O����On$���q`)Q��$="�0Xq \���I�h�	�# PN<ͧ�?Q��~����K�7I�	C4")\�zl(2\�L���|���.�����ğl�����R*�� �G?4`���4�?AsB%�����'
�_�H�#��6h�ف/�]�r@�Mk��r۠�<!���?Q�����~x��a�PA��c�ٌen��!\W���������'�r�'*\ !���4*���\0�r��Ø'q��'�����K��Y`Z��~>�P%-���l�{ҫ@��	� ��I���?Y��#}>��l�2��܁�`��,ˎ���f�+K���?�������OB���E�|�'a�M1��F�FƊu@U� �ډC�4�?ɋ2�'p:a3%�ējI¹y'��+E�r�	G�lZ����'��($���ڟ,�I�?�s3��V�V���*�A�K²��'�� ]/s�X��y��� @ePլLU�5�F瓈媜h"V�����x�F���՟��I�H�[yZw(�p���}!�yX���i3V��O��Q� 5��`F�����n� ɘDh�W.^f�O%Uۛ��,� ��?Q��?�����4�V�d�y�F$3���'-,��7i�0[s�o��� �Sj:�)�'�?ɐ�	2R�m �@�9���ŇT7����'B�'�&E��W��ܟ���[?9£%�f�[dF�K�feV
WL1O�}���k�S��0�IV?�p��#�
u�c��H�ĉU�@�]�If�\�'��',r��K>dӸ�/��V�)�!��*��ɥF۲�K�.?9���?q/O��� 9_69R�/�'B�\���!�&p��8�E�<9���?Q���'�E 8c*��ZC�\�e949�U@H5O�<�qT���d�O����<���.�@}�O����cד��,�ՠ)�I��4�?a��?����'�>�֦��M�%�S�A�����Σ~��Ԯ�}}�'R�\�|�ɽQJԕO�©	v�)ygl�?!��i���n7��O��|�I�h�x#�H"��%��%��)z�!ZT,F�6��F�'��⟨�S��G���'�"�O©���N�uƌ�+�AF8f��I0�&2�I�����#��E(b��'	�0l0��˓�1��f�.l��'_���62�'���?��:���P�LiNQ+���Z�b�>���X��Hm�S�'HVP}�c�$G"�A��)s��m�G���� �'��D]�����r)%E���¢C�!��lS��M�p "��5�<E���'�ݲ`��Y��@J�H�GN��bb�l���O�䑝zx��|z��?a�'���{�#O�_�d�� *֡��R%d7,U�O�'i��ُ;��bf�� 1.��� ƔJQ�6�'N-4W�p��ݟ���Xܓ'���5j*�J1)�+&��Q&�h��E(?��?Q+O��ė�:�)�j� ~r��J�D�D���<���?����'���S�c6�Z��t,�V�L�*j������d�O*���<�:�$���O�ͨtN�l=��	�
�}\����4�?���?����'���h���M[��b&dc�*ݚT�,�S�Qi}r�'�T�p��.�\��O�BaGA�<��QG΁=Ԙ�;�i�)S� 7��O��0��gl����;�$�/^J���r��;o�6�m����f�'d��П(�B�Wo�t]��+%�Be����G�zi˓�H�^E�d`�}��'�85e�1՘��)�.C,RQIaĔ`\�i��
���	ʟi���՟���㟬���?��u7b���y`�K�(Z��B�IC(����ON��s�ʭ1�1O��XUr�F�*s�m�R`#E�U���СU�2�'e��' ��\��ʟ�Y#
�I>�D�"`Ԙ������M��Hh}��<E���' &��G��2w@-)��6y�v��OzӜ���O8�D�z����|����?��'�8@[�BZ�ge�QYB@�	7��I�e<��5,=�1�M|����?��'꾹�1n\�	R��Q��I��HS�O"�;���<Q���?�����'Srȣ��ޯk�<l�@i�i��x�O��:V�D�5l�	�����Yy��'��(�!��]��Q� �BE��)���#��������?Y��K�ˊ�������A�DDh#��`@4�W& ?���?Y.O��$�����5a�*�I֢Q�%�X����=�*6-�O\�$�O\� �I�9�TP��g��)k����ّ&J��r�0e��P���	埌�'���ɥ;���$J7�I<F( �L�sH��!�U��M����'1��ЗL+0�jM<YU`N8y�j'ǚ'�HQ�S�����NyR�'Jx# W>}�����Әp�L�9�Ŕ'hn���b�~��}��'�$�S�������	��!��zۮA���T-��	��Q *�ҟp��Ɵ���?m��u�L�4.���fIԴeXD�z������O�I�V��;�1O��F�[��.PRF��6+B��0鰴i^�ӕ�'���'B�O��i>q�I)x����"�|ik���~	05��4/�)9�+NP�S�O�r��W=p;���7߆���;V6��Oj��Ob��p�<�'�?����~�bR��]��l�$|�ܠ��F.o��b�Р�)����'�?���~R��5c0\	��H�} I
G����M��=o:-O����O6�6�I�cr��K�
�Y4�2o�N���#�p�0U�In~��'t�^�����UW�ZRJ+6I=˷��(��c&��eyb�'���'��O���s3l(���mv�����Z<K�豪E&Y�1N�	����Ify�'@�cVߟ�1ݹ�E����h9�����M{��?Y���'��$�t���ܴ��m� �8�Q�l�o���'���'��I����T@�`���'�6�����)Y���SG�U�A!�~�p��:�IΟD�d�آOĪO��oB.o2�zE�ï8A��鲾i��V����6�~i�O�R�'��,8~{]+ed��&�r,��H$"��b�|��$�8��B+�~j��L42�s��H��`�"��G}����9PJ��'��'���U��ݖS�5R��Dh ��%�t�<��?�ħ֠#�]�<�~*�홨}	Bd۲&�>2`���˦�j��ğ4�	ğ��I�?�����'�D�R��U3x�<9yB�ݖzC��{Fdӎ0�$�@�X�1O>1��+׀ �8��%x� l!��M�$X�=�&�iz��'b�(Y'g��i>��	��h�H},I�b�q+�@3� �9nq<a��F0扬(�@�0H|R���?���K�dd8��2&.�u�	\Nh�z�iF��,N:�����ORʓ�?�1]A%���x�ā�Qcֵ=/�5�'&uZ�'���'2��'�[��0�L�N��3���R'�$"�k��Ȅ�O�ʓ�?�-O���O��D,)���x!�\h�Ԃt� x :��<O��D�O��y���O&��<Q����:$�iO�G�"�2U�L�Yh�'M�Ni�FX����GyR�'���'�l���'�Y
U'����,�f�l���A3�`����&Z$d��O$˓(�֕ppY?i���` ����Ņ�Ш���۝dTn�8ݴ�?�)O����O �D�z��|nZq�aQ'�������	�>Hy
6M�O��d�<!�̅L����|��?��F莚Z�PH�m���U��L�TyR�'B�'L���'�s�@��8�q#Ji$ y��k"�oZgy�l ,��6M�O*�$j��I]}Zw7�=k]T�c�MҊ=.��'���9��ꟸ��A`�X����,�R"2����А�iF"�X �*I�7m�5ӂ�mZ������<�S���$�<Ѷ�K�XH�ɖ8Z���(���6D�1�y��'���N���?Y���!x��x�&-J�0rt%K V
�&�'��5O  D%�>y/O��䨟T�T��8y7�t��D�IT��"�'���7Gf��?i��?!G��	^�+��;Q\|R(ں\�61OHp���>�-O��$�<���+wo�$v*���F�	�`A[%�Uj}���yb[�H��ȟ��my�(F���bmU�E��uB
�F31n�>�-O���<���?Y��N)��3��?y�ޝP�	�-'��r��<����?	���?y���d˱n�tΧqW*�Wɖ?X(�W�۰���m�gy��'����$�	ӟ�j���~�iH9JZ>�y�M$���2`�U[}b�''b�'���p����N�DH�w���`�sմ�v�ݱ"3��n�����'�2�'��J��y�^>7M�DXaRU$U=.\�9�g돮r��&�'��U��RW� �����O���0	 ���!�Z�C��8E
5ʥ\}��'FB�'��Қ'$��9Fj���-��lHVM��g{��@
Q���m�[y�Bտ�V6m�O��d~��)J}Zw�PU!��j�� 䇹�X���4�?��K�
E�}��s���}�$�G�>����˩<��M����h`:�M���?�����pX��'�q�1�j�襹��*9%��Z$�s�й�8OH���OZ�� ���?-�m�8A�9�$���k�&�����M���?Y�'P��FX�8�']�O�h�IG-!p`㊟���AָiJ�U��y�/l���?���?a�iJ3s�Q:B��3pG�H�Ʉ�t��v>O&�p���>	/OL�d�<����ˎ(�L�����!��@�1)b}�d��yR�'["�'R�'t�	�mgJ��)�?[��Ċ�#�<u|<D���Ĕ��D�<����d�O��$�Oހ d�˪�F�'��	0rJ���:2��d�O��K�^�6��OT�E{t}��>�Ҕ�r,�*�m��ረ�V�"^�<�����$�8�����σ՟L9�lɑ,�n�H4���`-z�������O����O�ʓxw��cF��D$�0��\r"�[Z����4a�6��On�Op���O����j�Oz�'�8��c�D�t�6H��*���sߴ�?	����$A��&>Y�I�?M�E���);4i!1N�a�1�4�ē�?���l�Z��������H'r�Xj�\�t`�PZ>�M�,O�,�#ZǦ�b��$���Rx�'�XLJ͒"(�4�!1�S��,���4�?Y�upd1������O4h(�Y�yYZ���\fp2ݴgی=�i���'���OZ�c�x(!��$ܥFY
l^�Rd׳i��5nڡHT�-�I`��d���?�����T��� �%k�H��a铍R뛦�'�"�'��`��=���O�����|ёM�>�,8��? �x�fӸ�O�pg�M�S۟����`�I�YsvU[��_">P씙��/�M����&������O���?�1@h��,ʂI.���ᯋ{��'P捺��'^�	��	ɟ|�'V2�qD��)��8�B�*H����G�VO^�$�O��O\��O�p��;�6 HG�S�T"�a�����l��<���?q�����6k��qͧHa��SJ�P�}4�@5�:��'���'�'���'�Z����'c��k$Kс>J�;�,R�X����J�>a��?Y����D�4L�@H&>�RT�16�DM
V�J�;�� zR&Y=�M+����?!�/�z�������&��闍9~�{�J�to6�Oz��<�')Lx��O���O݊7�@qE ��B�\*i�2E �$�O��� ���(�T?���%Q`�!Aj��K��h�pӒ˓I��Y*c�i�맪?��Nu�	��ܺr�#?��Yb்*+�67��O���[,���0��0�'/Բ��@�+
d@Y���	�W$�7-	��EnZПl�Iɟ������|��&SǮ��@L�%A����U$O��?��Aʛ�?9���?1��)�O2��FҜ=�|��bH$:���f�����ҟ�I�q�L�N<�'��I,I�ؼ�c�Ű�x1�ǀ7�t7�:�I��&>��	��T��8612�%�(�lx�ħX�� h��4�?����[����t�ɀD�p�m2��y�@D�%�l7M�O.0���Obʓ�?9��?�)OV�� 4XsA�>)� �xb�D:�Ig��5cw�'���I꟰���˄l�,�ۤ���TH��A�3'�6��ly��'���'��'�,���'B���^sU� �^H�����rӊ�$�O0�+��O2��E�&��Ǹi�j��׏c�hX`׎�&z��AZ�O`���O�$�<���\�������D5����I�uvZ�B槉�M����?��������O"Tu� X>2�6��U��9\7�\��4�?���?9�k����?Q���?���&���Z�'iPAb7��LD�D�x��'����\$\�0�y�����!	BD���gܝnF����'��-;��'=��'���Q��X'xn������4 <Es4&� 7��Ox�d���8ك���U�*�`(3t
A`�T�2�J�o��ŅesH7-�O����O��i�i}"U>��kT�"MriqDm �f�n�	��ݻ�M�Ď����'���|b�'�$���N+"O.��V��T��y"i���D�O���F��f���O��'�?�'.������;��d �k�>.˔�&�I�d7�AK|����?q��v�t�z�/�9C��]aR����m���i�b��*+^��'��꧳?qJ>q��_6�<	�'h�ay��n�/F�|z"5��8�I����py�hH���"�?}���jA�V��쉤Ǩ>���?���?	�����o�.�A@�<E��$�V�:hvX�t�|"�'R��'R�'\���֟��3�?f,��&�Ȍ���1"�ir��'�r�|��'�R1����4i���r��>uڦ��#�"V��9�'�.�R逩.����O(Ω{��m�`���:8t���'�����,U+.6D�e�
�1��p�'�Xyh��h^���&��Q�ұ������j�$[�KA�{���f۾�����D�����cd���lY�Jܢ�B�J�1�����ǼR�NEʇ���&����3���W<"|KtiR�|�d�C)F3�HD0׭��R�ʁ2�nǚz�Rd
O��@����m���2%�^E����O���;d� U	"�V�,~�a�h �I ��:�*��r�]h�������$:9 ��'ۘϿ+gb��"�b%\���y�fԡrv����ϧa�PT��oĝ@	F�3\fV\���2Cf�,/�G�M�<3�l�2$ $3�l�rҬ�$5TҘ�C�'q�����x�O����Y+�"�����-/t�"O���D���Y�$�\�֝ۡ�	�HO��@�����,Yͪ	[4��b'�i�I͟��s��NNa�Iʟx�	�[Xw���'G����&I���p��:h��,��b�O�3��g 딍�
����č!-Yl�PrH� �>m���#9t�9�#C� i���?�=Y�)c�@�pƾd^ք�u�K?a5JUɟ���c�'�剣'�tXF@�.��9S�%C�rdB�	#K�Y�#�#l�q��+ )-�^�I���?ŕ'�(��b�:9!�"��o��ᰱ�S�C*q�Ѣ�O����O��6e-8��O��Stf��"�@
"g(u���0��
ܱ/Zj�!?=@|����%y���Ó&-0����
0����É�;]���x4�5��	�P���O6����Y.S�
	��.�	���5E%ړ��O���:,V��RD�V�z����"O\� F��h�v�b�fو��6O2��'��I�ndDPݴ�?a���ن��9��� jVr�:��.Z�ˆ)�O2�$�O���E٣|� ���O8\?ne��|:Р��W��H�D�Bo}����J�'3ni��Ϋk��h�W/Xޠ��V�cl,ꓪS�z+|�ᬓ���5V(�B�'� )���)�֌y�N�D�|2с�%s�Xದ��L�${錳�?q���9O�`9���5R��Sꞯ/�`�p1�'�OT<����C��Ĺe���� D:OМ�4O
ܦ��ǟ��O!� 1��'3��'�Hpd��9�2��S�OU4Y�.�v$`�k��/�T>E�|�	$�V ��UIU�pkq���=�R�P,��,�U�O>E��pr|�Q��=cEF��� u�6�7�Ǚ�?a���?Y�����'wJ�X�m_�B�B�� �y��'��}�*�-,�� 5n�sbT�1�	<�OX�Fz"T>	�'	v�8%���']�T���Ȍß��	L᨝�`@�ʟ��	џ`�ɥ�ug�'5r�V!T�$I{��MC��9sK��~,V�* ��j�"J�m��x��	�4и�R�Ҳ�Dx�aɦ{�~��k�H]�t�O��Ybu�'k�Ua�*F1ug&`� �Z<���'6��3�Z՛�-l��� ��f`��LQ�>��D�2��0 )�"Oni볥ֶ۰�`Ҁ� �fII�'�����M't�~mo�OF\D{6��+�lĈB�G�d��I�������E�ϟ����|��Ό�&5$A�g�L,/Ҽ̂RIV�"Mc0cܔL6�|�q�E���<�%�zZ���r��1"��&@X�)
�[!�X����5V`�Ѧ^d�'�&D+��?	�e��v�5Q��;@��5hՒ�?ɏR�s����
*��:�X�&�����$D�|�e恢D2��m�z(2mh�x��)�O$�)��T�s�iLB�'&�R�8 B�j�#m�f��'�Q�JEd�� �����П��0
 ���<�π "�"8�q㛴|zl�v剫V[����(ڧu�P���=4{
M�"/�LC�<FyB�ˣ�?q��)����[��Ջ2�����Ty!��0(D���vÍjwԝS���ZTa|R#���13=���H]�d� D� S�Q�$*$�±oş��	G�$�W`R�'Fb#ʇ><j��OB9f~d�)�b׳&&&��p%��%��s�XY��"��~���;xU��'Zt�`Q��Ǽ\�t؀waN4h�����b�|Hz&-ɗO;�>�n^�s�,	�$�C+Z~@tMO�x$�(���O�$$?��d��?9�ع3����ߘ�)� ��<y���>i���/�V�H���:+1�`�w�@D�'	�"=�'�?�ER�	@����H'.�� ��C��?���r>�c����?����?��*���ܟ�A�6M6�(�DЫkؚ؉�｟$[C�I�6Ѱ�R��ί�p<q��4�Nu���#��8��Zp?��LN;5�F���BUW��x�E��X�Aj�e�6�*���	]r�]�2�'�����O���l%�(��a����+�����ȓ4U��p�*I���/��j	�YR��d�|�*O��ɂ�զaX���:c�>� �T�?c�%#�Vş���ƟD�I�g+he�	���' FYu�ҝV��ع%��xH=�$R<�~�H4�k?��8�F�Z����lK�?�����`�C�Ig!�U%�A�Äݕ%��b��D`X����&�үd��"�lÈN�*����Ֆ-^L#aJ�Q�?�C�s��U���D��4N���)��f0D�ta��ҹ,5�Ɍ�hp�6jn�`��4�?�+O�r��)�Iԟ�O�|ܰQ�P	]������Œ�d��O0���'��	��y��T>�`#�4_�r, Ҽ@���z�H:�v�D���&�F�Z�K�z~�"7N�0�Q��S��OX��(���O�\(7�O�
� &ߧ\A �TD�O��"~�8�4T�)F��mq5A�-n���I�ēUDZl������k��Շ{�4�r�Y0�i��'��Ӓv�܁���,��#(��Iї�ưu��+f#��(��}P�N鴐Zf�!P��遾��I8��O޼C�˿S㾕���˔|� � �/>�vd:�(W�<�Z�Ȇ�?�Q?��Hb�����U���ck�,׎L)���O��m�X�IS��T�IҟS��%�z,��.R�BM�JL�@��Yx��� L@�����0����*}�Ǫ(���|C�O^ls�"��@�W�Y2y~�u��b74��92톊ܦ6�P���9f`WP�<���2:}8A��R|dq�q�<�%%�,�������B�BIg�<yd��-L�z����(_V����O�<�խ4O<0	TO��x�]I�<a�MH  ��A�˖J��+�� T���d�[נY�TD�?�ȵ�si6D�<24��{Ah���� 'G+NO��y�ƈ{�p1��Z�dfp �Va��y���k;̩���Y�r]�%�B�yR�J:nN���A#]:�xţB��y�NN�w��$�ÒV&ne��i��'�n���͘ %x�\��5C{zq[�',���kz�*5HR�V�<{DhP�'|��K4��Z�k73��R�'�d(����L��!餤�22?%��'�N�����޺���-��3��u��'&� �E�ۡa\�,�JN7+b����'�Ji���
��jx�)�#h*�I�'�Yfm�'3 x��@�=JYVl1�';:�C$�P�h\��X%'O�G��h�'d� (%�ԛD����50���'hN��E*BvT��$�;���'e�A��X�2�6piPÎ�[l�[�'��e���M�x��t+�� 
�I	�']x� 
Ӊ,BJ���?y�h���'S"ՠ�]�D��!�'%�r��'��q�tb7:ώ��q�ֺ԰��']J��W;}�QD(6bD��c�'�BY�uD����0��5+b�5���� .u"g ���P{v�5
=�;3"O�{�M��z�ys�7
,��"O\�$�-;�"=I�m?'d�[�"O��;6���v��s", )�lV"O
T������X������4 ՞>����gX32-�U����<�
p���&R�}:�8R�̱�|� Z����@ 7*�c&�ȇ�ē��1�@���Z ӕh�ȴy��nt�PH�=I6�sƈ\{�S+$��m���O�z�a.K~�tc�!��)%�����P�9����/Z6�bؚV�ɩy�
�G}Ƒ>k`�DefM�"�L�7k�k���^4�V�(��3���ri\� �dbE����5k/�@W����Tj�f4����'V�
�s���
*eFl"�XJ�|aӦ�O�QkB�E0Cq��ABaA<#�(��q�	�f$^1O�<d��16��k�S�4�r�]ґ���Qa�;3�R/r8"���/?yqjV�:,`e����+�2p����nj@�ۻZ;�Q�@���C�`ϓ|���5
�	����,y�1��*gz�B2}�GG$䅹'�ԪW�&u)1N�"�t�rBNF���cJ�r+��N|Z��״
mF	Y�Ş<vb��F/;L h��g��zb���%ǚ.|b�� ���9Fha�#.�*�O����.X��Q3��'�z�.��`@��<�6�R5��G:����%& ��샧e��; ���<A��<|R��;勄!H�4(+�@�:dl �c���O��"G��f´�J�O�6B�6�Dߔ_	�T(��^��
����L�( "i�����$���̓� �P �����ɼ;3`
V(��3#ƚ�W�v}��DH~bJ�Co�����p��Mb��	*�5��c��@;�c��(�dْ�'3&!Y���w1v�&Egݩ��,¬	��p��Ml���;������<~�Pq���Œo��0���աh:��K�-�`���':n����K�J�'��K�d\�0C\!�:ષ�^�{��a�C�5L��t��:�脹����o��x�o��7��C�.��| Hۄ����&zQeSh�X��$�dC/�ug�x�)�!Ej��kb�R��.��GBD}R��A|��#p$]�l/y��',tL��O1 �R,� �A:8
�3�{�(&\�qO4I�'0�X��a���:���n�+�65� ��?��U��li6(Y �����@��Xg��zI������Y�^��I�ܥ�SÏ=Gz2 ��{�ώ}��nǫ;c0�q����j�'����e2��!6ləx+ڜ����N@�X"�'C������9�	�՟��<���w��P'��N����(E�;h�(r���!5�N0���L`R��䂖O+�3��۵*�D8���'�.i��
X �M�R�(3�O�>�S��9+ ��"��]�.e�l	!�CZ؞�	ѭ��m�$ט=0�2���L��
"Ȕ�)��mH ����	�<h��'���H���`�O$ C�����=9�,"7��*��$B�(I��'�FPyv�I&���O�ظX �P1����]�rcv�J���k?�uE��OnZ���Gz���$�F���U��z��1��DQ<:�r��dL��̡�c��H�ġ�O���ɋ.[��j��'3!�0�G�dϐ��-���p?����D���� Tgp X��Qn�ȑ��(��8��*Dzӧ��O���2!�M1��4+�=�$A�8a|��Ij�Ń�h��4`*��\���I!l��{utK �R���� 9w����O�����{����F�#�h� p�U`�Hܑ]�X����I�;�F�!�`�8@��Tb�@̱X��@���\�y�`ȐJ^��8���:\��`�����˪#?�3�Q�*1Q��:���1D�ĊK��p�<1@�Ԫ4�qq�3��g~�(�����Z4a�hR(�P�$B��u����}b�f:m�Ϡ,�0����
/[FhAc��æ.��Ik<l�'�d����?ͻWnI� ���j�buR�-�i/r��/ZQ�t��3:�Hx@��8;�>i�6�U���1��|���'n�rbH�:I��O<Y�H��6�*XX'��1|�.�����u�di�4F�x��s�����?E��@Ip��%'�(!�Q�X	��	�D��Zv
��P��g�')��� ,)�%Q`�lj<(��OR)I6��|Y�yR�-5���$`��б-�tJ�)N�p�[�y9�fD��p?�g,~,P��b
S��0�ɏ�N�f��,OLDJ&��.:�?Kn��������$�����7�޽  ��m���wO�%��.�,����FI�L���A�n�*B���NP���0F-��OT��?Q�Q��J�QI�.�8�q(C� O*��B-��$��P���B�fՃҮ����K�5{M�0~"���O�=*v(�>���O��(*���1x�*a"��'��´�0���Z�J$��a]?b��;�B$P����	�0�;A@pF��fʕZD��&��[ff�Wx��!��2Y:~�#��� ~�`L	�e�<�P-���BX��sִ0ږ׽<��`y��U�v��΅�AvP�:C.\��j/��?I�#\S&� 1��*Vq�HKgD��a��2a*2��1A���n� o�����\!"7J�LTH�is'��;0y��	��&A��J]���D���-.���N�Ge|�J��+`���0��<yP�W�t� � �C�Ax���n�1��T.ш<�$�A��'?��L�U�h�"-uȬ�������/�$x(��7����1l
�k������H?Q��e���� H9��,w��adk�Rβ!����eF��0��]=6�$�Y�H8��7���i�'N� ��0�,|ZQ�M�2-�DH�E4�H�O,}XU�D�S��3�b�q���*�)�X�xu�
3#��X��,.��0$�U��1q4j�5���O��V��q��qYR'�#A*R��՘>ᶬ^�T� S�a��'&j���8�@T4=
,j�Hvf�݉�mE$�굑g��� f�bcNʽZVE�d�N;9�����v�`��W�Y��3�j`���b����ě��<G��`@�ˍ,2uAS��g�b>mJp�޺Zq�$3���W��E���F��lJtÎ}�N-�W�V|�ڨ0�jG1��ɐ���0y�z����}��P�*?*�'UFP슥E]z����K�I�K0,�YW��J�p�H0.L�!��ɸf�Dʟ\���1!��%�%�ׁ$Z��bᖤ5�l0S2�[��`�Q0i]z(�tC�:0��(��%0�V)\���� K� Ic�֓v�%�'��i���gm&I�"�+����h�4d���8Vf�`$B7-95H�$�N*�L��DԮs("�Q��P!1�a~�F�X<X��fa�;�|I �� ���a^,ZQ���*F�4��ŀ|ٓ0-����I`pb4�t흵�ƙ��̆vj��:$O���p�L�X@x s��Hp�$�W�-��tȅ�4ϐA�'7�L�p�R`�<�;[��8T�O8���Ը-����nX�?�<�A�'$�l��� 6C��#��(*M�4! [�"���àI �:�Ύ�]�a�&��.-�ӊo�y�c��v����D�%8`\��f���$��`�����&C2v��u��Q��*0����4Ji�l`֥ݳB���F-qL�u��'UZ@�R�ʔ)���{��L\*�Jѭ&h��M���Y�W�ܴ��Oq��x�+�C�8����Xh�xo��h�VH�,E�!���2�=�r?|��S�֓[�f9�Eر,/ P�q�O��H3�Q�lB�d{��[>H�+G�|"@jp����39��� ����X-.��8;*��@Ex�����
��((�G�΅g&���W,H�K.p��$��;��]zb*;<O(uєA��a�@�h��;jm�3���:�(��3\�8��n2��5$i��yC��7�`扬V�(]�Fo00Ĕ�2NM�B�B�	�f�����"-6ܐ����n:,�x�Ι���!�		H9�0�&�O�s�0�"�c�Ճ4�C�#�bqE���<o!�ԁ0�Ӿ58"lۆ(��H%)'�?-��#ôi���I��h�t�'t��UI O;*��Pg�=+����I'�
� x�ՁM�~�x�`� ��?��"u�N�� �� i�ܡ��i 0�(�� )ܠ��a� ��c�V����E j��9�ZJ~A��@��i�w��T  �quT>c�Pʄ�� "w���E,M�Ԑ r�&1�	2.�%��A��ѓ��H����'�$oƆGD��:�K\8>\1�DJ���U����?F�oܓ�xb>�R.O3=Z�*#��6�B�q�,%`�5ѧ�K�r���c'"�<7HQ��#i�qr� n�0��
�69^O\  �C�b������G�r�̧.U��U���W3 ��S��8p�V�9��HX{1�}�����?i& ��{c������Y�"�9j�����䜱MD2,��	bQ�β3Fr�]5 ���[��^���Ê���'���p'�5;�45k�����>A��^	��qr��L${a†V&�U�p-�#_��S��0姚�+	��fh�N����O��5hݘN�p�
�ڤI���+�7O֌�p '�Ɉ�M�� F�t�l�0a��B���1�+Jz��)���j{)X�G�/JL1O(Z�O��p<������'!G�-_h��0CNQ}� w�b4�r�ǛL��5���=L(�#)W���I�)��B�"�i�Y�TIP��  X�j�S� aS��`;��{��z��!(j!,4K2ˈ�����s�>P2��S�|z���&rS�Ic�]�N���4lB����X2)��6��֯8�s�l���S-�<J���@L�tKS^�|�pU"͡@���<�!�/���� �LOܙ����<V���unKB����ɍ�(�X��gm�<i�Ǻϓxޖ����0 P�?�B,TL�0嫄:%}r� �̦����_&|�R��_�B�����IC>II�Y(!|Q� Z�):K�a��Γ����%�6Y�:@��&!��	ܢ(Y��
�wH9��!��k���f��5_����S8�����5.V|Tx���ß��@��4y+e�=r����@ 2�2��(\�R���d�� w�H�@����ˆ�Q"�y��4�"S�
�5U��lyס�6ؘ'7�m{ө����JW�9OP��%��j�dȁ�ˊD����\�:@��K���	)G8�t�ҥ�.}�bX� RC�䚐-z, 񃬊�G����L�3߮ۦ�2H��r�}��<����	�=ᑆMe�S	�v��ɪ���4
�9J%F�MC��O5Rq�B	Gi���Ǔ6��1k���I�J�cTE�G"��k7��v��I5)����V>����D��v C�A�Rb4�k�H���8c�1�H�� ��b]ve��t�7.�c�ā����x��AW1=c��[5�K<h��T��
/�y'�;D��#V�Щ\�F�m����'jF �e��GB��A���O-�ˉ�>(" �Q�Ƅ_aA��	���LW?T����uk�O���P������D~� H�y��a�8�䚸]���'���;.��w����O�V�9��Hf^��-I)M�X����i������ux�$+��+[Y�x��G�g�nX�0a�
/�6ТoY�d|Ex��5�&��bjq��I�ٟ�y�3�)� ~� �)�#'���E�AT�����mH<1�1��u ��@�T)�Û�y�cS<+��`�#O]a��0�!�(�yB��4)�� �b�:\��kW$֮�y�C��'\�\ԡ�ce~�sQNE��y-�<?���M�EMd�pֈC��y"�6�DA�n�DV�դœ�y�e�;f��i�V�.g7� ���P��y�'X3;/�![cU�fW��B�B�<�agD�^��	$o�IQL	Y�u�<�ԀR�'<$lQ1c�-RR�I�p�<Q�Ii�p���+<@ u�7��`�<�����y��nH����0 ]s�<��F�+�����~�>����<T�P��eK�w1���HG�`o�L�� D��r焮�B\�c�6"ߎ@��;D��C�N�(Hֵ;d��1#�r�F#D��i~m}
����^=\,�e�!D�� �ӺI������$�:L�� D�L*U�1
�J��O�`<z�vN>D��!��G�z8򯃶Ail�{�f0D������7`"T)�h�=�p��p�/D�āFʟq���E�YX�#WO;D����!�"L(X�t����`0��O:D�$ˑa��~v
�Q	[��1Wi7D�@�HٳA��L�A�2&�zq�T�/D���ŀװ���@1@��0��+D���#)I}Q�Pr�D�  ��ɶo*D����˻ }�a�r�]1��)i�*D��"�� g{��$�!޼�1`A;D��JD���k-p���B*}g�4sO9D��ke�G�E�.,�c�M���B�e8D��0!@�-a�����ބG��Pwo6D�X�t��;^P�uc�`����3D������S=&e"'χ�*|]P6�.D�P���8N� $	�=�Ti�Uf"D�H
4�^#mK@\E��2x�B��e"D�J��ۺ$bRp��D*0�E0�"D��0�ϣ���Y��_����?D��dG�'6M�V 0(�%���>D��k��E��liP`d^�/��e�"k7D��2$��,�RȚek��s�j�B��3D��j���FX���gJ�L&^�A�1D��o�<(vV������P�n�C�<yGK,NT�J�G�#�4��� �}�<aE� =��� ��^�����^z�<�n�>�����⍠��*�s�<q�i�ZBV)�A�j!#^y�<ɵ�U!Zx}��U�]�����_�<i%��w<f�s��%s����]�<a�a�O�fՂCV��HE��`�<�w)	_2�5�.�\���Я^�<9���p�(8�e/؈]���!��r�<�g�/Y"t�9����d�7n�v�<t�U�%�z�� �q��@c��s�<�"OE1+$x��Ŕ+�bų�h�<)�G)��8�b�Zx>����c�<QH���=[�S�XJ�e�	�y�<4�	��<Xq��ѵp.�e��s�<	���œ�*3^ v��EV�<Y#쒅[t�e0~hTTC��Bl�<�B�F�G����V*.�����L�_�<�� H�	l(4s���֌���^�<�"��i$m#�C�(f�dA�Y�<� ��$d
;Z@ك�R4
UD��"O��!���Yf]�c,�;G�Y�"Oz�ۢ�����,֓G|�3"O�륬ۄ��e�RK��.�b"O>(����E���� �ә	���a"O��a�b�3ъ`���˽K�V�@"O.}2�ቚa�^�Z�A]nN܁"O�=�	޿{f�a@�~�8��"Oz]���Z�*	l[1(UW�ཻd"O���H� �pT`07cs�u�%"Op�c"�"3 ��2��#u��"O�<����-Dj��#Lǿ4t�k�"O�C
�~�pLJ����?� `��"O�i�Hր2�
�7+��g�8���"O�Ȳ��P1y��M��ꎞ�<���"O��BGx4`�G7w��$�"OJ���V5pX:��fJ7���a�"O��N�40��!��a�,ˡ"O�D��r�����%&{��t"Oj`x-�S�b�[��B�,]̘��"O�hU�=ok��HgN� ��,�"O��C&
MGA��K�Lk�r�xc"O��k!�۱x�i���EQL!1�"O�Y����r�H�6FO��01&"O�M3GМ���{t�F�)�*��@O8�%aB�-��Lj�`Ǉ*}JIH�f5D�Hct��'�p�֪ʦ[j*�J�L7D�p�%C�&q�( �&��Z��T��5D��� LB�i� 9�d��u �S�� ��5�Sܧ
+2pi�o�P2��3�K93��u��
�0�{��z��@B"ܷ$%^ ��H&�ha��ږ��TP�ʐ(U�֥�ȓ^�:@�����,0��`"Te���ȓpU�*��9`����/K)	�ڜ��8w$�`)V4ʚ�RAb�9 �ȓ|�V��1�կeRĄzr�����ȓL$~��A	�$����cO�W����Mr���d_2$���NʄPn2��ȓtv$vE�
y��8�ҷ��y%��E{����P�~Ix��E	��e�J%#�B��y���l�"@��N�ꬁ����y�戙hy$Y����V�YPK�y���>u,� G��(�.��g��y�(P>T�|��d`[%):(m��yb��1sRu�T	6�޸Y����y��v���F�+
��݊ ���y"H�;�6 �!�3�ީ�w/P��yB�]�!�d��H['qE��H��y2�'p!�`���� &c�����#�yb,�'3~���l�8���[P�Dk�<i�R.��|C�]�?Q�=K�mDt�<iUE3{f|ݣD��U��jq�o�<��c��o��!j� |N�{cpH<��	���a��y��W$�< !��2�PTȱ��\�*���[�!�d4�
�A� �Y�̈�"�!򤗠k�L�[��~L�
f�	�=á��Y/.�J�@����C��؅�yB�*��i@雜U�v�r�e��y��J"f(��ZCFΓ]0<T����y�,�7C�L@E
�Z� Z�D��y��q�dc�%�&M[!D ��y"�S�%<�Y�t�ڔn�}A񨂅�yr/Q�`pug�$�
B������ Hxq0�7�e���.I�F#u"OƐ� ��q2�G75ڌ�2�"O����^�o�,��IV"�f��"O I�D�5�J�N�����'"O�����I��z$� -�N�F��!�'���-{���#5NZ�XT ۅ��?�TC��?1��P��NFr8Ȣ�8H��C�ɡ4���7��{�0Ȇ���B�	�P�n��Pg�4��m[� ��q���0?1�(Y�~�:l�長{�8+3�E�<a$�:4~��я5L� t�d�f�<I��{�|,�W�Ȱ&F�y��`��m���O4�<��E���A䈷!ؼe��'���:6� L�ll8�,�p���i�'ND��W��=~��d!�&L�`4��c�'���2q�S�,x��ͣP>�M�
�'9��ro@�&4��L�K<�ۓɸ'0ܰ��T1o�����J���K�'_|%�Ҡ����I�r'�7JH�Q�'/v���H�E�<�Z���,L��	�'�j	�"*��p��ҥM_�9n,�z�'���!�.��Q�|���э1x҈�'`\�:b��}ښ ����>�P���'�>C��U)z�0�:�'@�dS�m��'���v� �+H��c�E�]��k�';���d@E�o�8�cO�ln��K�'�
1iK> @'�^#f#�c�'�xX�g(=v���C>Z���j�'��Y���G�8�nH�K�u��'s��k��.X֖͙T�Ůp5����'ct�C����3�0��AbS�h�Nuh�'���h�V�H�L�eB����'���Cb'�4=>�(�o8�B��'���X�L�a�\e��Ó�iFP@�'ab���N�7�,�
A��"x �'=6�Z门ep@�p���%j�%3�'=�ؒs���M2�R��%	�t��'#�\�W��+��!3�նI�:���'��X�Sg�X�,�Yr��A*�P�'T�Mɡ�и\Je�a!�>�Ĺ�K�|���=XH�S�#'�����D;����f�`��c_ <�p����~N��8�$D�,��	D9!~���e��)r:�k�� D�PZ�`O=;vxk�`Y�!�J�S�=D���F�0<��q�i�-ll
]��:D��Q(�c�X(�cjW�p�.�ڒ�3D�pE�F�C����!�(���2D�\S��-4��8s,S&\3�9��.D���`�Z�'����D�� �ه*+D��+�O�hT��;4	Ζ}��h��)D��J���6�`�r$i<a��%3b'D���ю���S挤Sx�iKc*O�AX%���t_@´�Z�,�=K�"O �b��(@�L8vˎ�!$"Ota!��O���#t��!ńp9"OH�$I	�O��|�7�9j��
�"O��z��O�VŃ�E��8���i�"Of���+͕sHܼ�R�0n �{�"O@���@ݦO�<\r�c��F4Z���"O��;���/Բ�����0 "��P"OZ p��I:m����6���I�Tٱ��'���$#v9��K��vǐ���D�/UTB�ɵR#�!(�A�D��q�G.u�N\ˎ�*�g?�CMJ��)���%y$ܐ`��SM�<� �\` /�CbH̐�'T!,Dx�"O�U[�&�h"���H�-s%n��w"O0yѮ��[w�Ȧ	��-�"O�H���C8E��bq�K�p:X���"OH�� '�=d�Ld��4D����"O�I`��/��c���6H�.��V"Oz4�D���#t��;|v%�"Oͺ��A��ԓw�%f���!"O��%A
�ib*ŽAlX���"O4��w��@$��[�H̠Z\|�V"O(�{Fh�0�N�kW@W��Т"O��&��9t���0 ��V;`t�"OJ��coܞ���X�o$����"Oi@���""Q i��nCV�#"O�@��aIg��M.�$3A"ORh�툎a�*\QaK�^(ʑB�"O�t�!��:2j�m�&�7l�Jѹg"Ob��'�
�=> ��o�D���2�"O����O�D��hI��ܨ0I�B"O`�Cbk���%�g�E&VՒ�"O�� Vω�zh-PQ�݅ b�A�"O���E%@g\��B��I�hm�"OB������UJ֊J�l��"O(�I�z{��J
�4�2!�0"OJỲ��;;
mQ��Y2d��x"O �f��<�D]��Nz�f�0!"O�uI�[�:$@�!�)ψ.�L�i6"OE�����&��P��1W�t
#"O��S-K�/�)9�%;�"�ۡ"O�ً�Ο�R���5� �M0BD�"O���ڞA_��)P�\�.��)�"O^�b���~
��c��Êj0��G"O"35Ā:,��ꌐ?�}��"O�݈�E�7y�@ I�
 �y[�H�"O��E,C+Z���#I�M�Xi�"O�����(&A��xBry�R"OL��U�W۲������(�����"O���w�#X�8��$�X��u"O*љ���O��ЋԺ�,��$"O�#Q&��NUc���i��K "O�i+����4��JS�̱�BU"�"O��`��%*�����@�B�x<�"O���� (�(����[�i�0%�"ObL��IQ�J�I�g��4n^� "O�Q#,�%GtaB��=�b �"O.�Ae�Ib�^m��D�~�cb"O��$�T����V�G�wނq�"O�����7H"�RSU'O%ZX:A"O�Ld�S&h�	�t��y{<��"O��2�]���	R��
3x���"O$���Ɂ�;%�Ac�ZBb����"Oޙ�M>y
� ���:��G"OHi�&!C�}N�]P��J�;�`X��"Ohu�A펕mT��C䆹Q,�\��"O� [�\X-���3���&�S�"Op�ꇎ�mƈ4zqg�1/�43W"O�q�C��D�>�K2�B*7�.��"OtԠ�΄!,D��[7�"O�ݱ���"�-K��^�2�J�j�"O@�:�f͌�@���5}i`0�"O�P���ϲu1��o�6X2x��"O `#�$�����[�D��(Ir!P�"O0Z�،ـ ��	�p0�b"O��A�{G���E6%'�I��"O� `�Hq��Z:)с\;���"O�ڎ[i���� �4)#��0T"O����^�
4���iuN��"O��vbـD�Ă�Ζ�Un\�@"O�l¥hG|vV+�nT�LŮl%"OpB���ԺI� �O�p�R�"O�M����|�=��Ĕ��`��"O�*5�Ɗ8r�e�ήu�fI �"O�iP��<d}���d��43�"O��S!Y�ܡ��,ީ�r�*@"On���\�L4�`�l�/9�ָ5"O��!�o��+����}"l|J�"O�
b��x��}9&k��"���"O�*׉j3��"i�6漃�"O�H�a��E�|1Ag���#�"Oz	�kTo{�
�&��(����*O��s�DJ
F�@���:` 	�'������!��dI�	��h"���'�����M�F�~�8t�^7�X�
�'V�k��9H̹�f�3Y�"��
�'n��ə=�"� J�M�F]
�'`R����i{�a@�/�|����	�'�l�y�H�:�-4z�i�
�'n��2t�-a�HuG���x�H��
�'�89wh��X
��Pf��3q�|�	�' ��W�}�D�B	��[�l�Z
�'��4r�_{�Fm!�N
&x��	�'Ҏ�Iu���^30�Rq �1 ��d@�'\-� ��)څx����NuP<H�'�$PiӉ�?7����$bR2Gr�,�
�'��T���_�'�( �c�K�M�*<�	�'���Qw��9����	Iv)�'�X���X� @���P�k
�'�B�Q�M؇s��]����N���	�'� ظPk��u4J��A�� `���'d��#C�s�����NEP�r�'��P�鈏{������I1��'���cu���s4�ZQk���6U+�'������� EZ&�#���
�'�aSA&�y"�:V� >���'� � 4T�\�Nݘ!�y��I*u��<���Z[y��H)�y�I�/rBޝ��	C�O�4�!�+@7�y����lyys��xX����@��y��q�",�CݻZu��K��y�o]�[IT�T#\	~��Ie�R��yrJ�*R�ʌ���H���q���yb�Q��v����ݑ~��@Á�
�yB�2(��
�$�=`7�X�a����y�
��4��QT��E:��z���6�y� �o��i �ȳ;��"C���y��Z�]��p���+_�������y2��uR0Y`�bU>
���$J��Py"�]��ܑ����)6���x���X�<�f$��3����B$PK`�H��HW�<���6]��ձuOT�~��,�l�R�<���*U��Ic�ᑗFߪ�0�)H�<i5�^:y�*u��f@���|� M^h�<�B�O6 i�r�ND;fl�i�l�\�<`A�V�`��.X/F{����GTY�<�+B�r�%�fݴ@Q���X�<I ��]�2u�0a��{�Ah�̒~�<�p��=��\JG���\2��[�.�t�<�QC�~1\paю0
�m����s�<� \���L�$m��3�߄O��8t"O��(ӳ���v��?�Z�"O.ố�!/ܜ�v�ԝRG�=!W"O��B�(��{c��(h)��g"Op8��5�
��̚�04rACu"O:�Sjy	�\��@~5�uH�"O��1�!�D��0��o��y2�Q�E"Ol��*N0(�r�@M��"z�(�g"OP�5O������G�Cb�9�v"OFA`�OZ�*�� r)0cAtQ�P"OR�BA�?B��"��*ŮY(�"Ozm����jH.\RgN�q���"ON�qA7h*�jS ���P�S"O|��7bD:R-�����(��qD"O�a(BK���2g�F8	.TJ�"O����	PQ6���e@2�� �"O^e�"Ƒ�!�2�G$]�n���"O*9A���Tu�IsF�J�\�݈�"OT)A���s��Ԙ"P�p
�,�""ODTq���6z!�r��.[���#"O6�آ�H�5>M�q/I5��h"O(̩f�
�s�x6L��.��&"O���œ>uQ^����p��5�"O0 � ���xŘ�<��[#"O��ȅ�W�9�@�҉��7���h�"O�xˢ���j{0�9I��P ��;�'���p�%�%d�A��Fε|Kh(�'��-	+�0a�|��6��+)$D�x	�'d蝨3�غY��!7g;)�:�@	�'�l�`����'N]���D��'ڄP�G�ˍ��	z'I1�mp�'�R�0��C'\LI��!p~���'$�UB��V�%�lQ�I�:fz���'�~�k�J�T�j5yaI	]��;
�'�$D�A�ɒX� ��W�zeP	�'_�=;T��!�|����Z T�(I	�'Yz� @��9�v�,����'���P1e�[�ݱ�hנ"����'��V[\$� u�.�k�'L�Pԁϧ=�% ��f��3�'E�D�Iެ�:̱��g�@�c�'6
x6��-f��IU�ѥX�`q�'���I	3����k��Y@�}��'6�X�����R�k A	�R�2��'��Mʂ�����5��$��)p	�'O $c�ğ�[2n�Q��I��p��'��3��I�u�jG�� HM�mI�'B��u�B��DJ���i�|h��'��MY4���$d�H�(��e��!��'���3e+y?�����2K:AZ�':�]�P���r&N1{�nۥ5M�J�'�U;��n�����͛&�ޠ:�'��� @���C"��;	�'�h����L�y�E�&H�
8�Y�'v�}�6�	�}'2�0F��d�ҵ��'i��!!�ˉVR�eC��R%Lt���'�,|�da�z�hxG��M߶9Y�'NU;��#4d��8Wj[/tK2�'>\pI6F�k������	p�4 �'�8�Z�l�qb� �(ҖURH��'��= ��
e���&�������'e\�
Q'$ ��ᝧ�h���'P�0���W�l����Iԩ y��#�'i�a��D���-P	�{���S��� ��8�m��?Ϛ��H��d���"O���gHyX|���T� �"O\�pD��)�%�f�q��M�U"O@��ZސTzr늏���"O���aߐ��|����
o��Q�"Ovx��C\�rH ��W��-}�Y"OJ%����m�hT��뛘d�  T"Ol�@ -Q�081�I�8���!q"O��9��;�Z�����640�e"Oֈ@�@�^�¤r�C�6��!"O�
u���a�����
&�lИ"O^�y���9�@�'%����"OF�#�`���݂��H�h}Q�"O��k���:��g�]�`��b"O�D��#_�H��\�����_�V�z�"O�4*
/� Qe�1@`�2s"O@!��g/#X	�N�2�0{�"O0�+� �X�FA�����\��a"O����cW*>{�e	 *߇"�|9S�"O<��6M�,bϮ� �D�p�:��"OT\{��=/�,�sl�"9x��R�"O����Ťw\��2à'h�J@��"O��PD���;L�S�_)gK� 0#"OƀA� E" 0����#��Y-�9��"O4�I��@�zZ���^�աC"Ob�Gᓲ;���� d�ޭ�q"O��ƞ⾜������"O�q�-X�+�0H�'i�&.��l�"O��`eK�w�*�+��Ǫ0Bq(�"O.u����DF,�ЅΥ8&��9&"O޸CS�E�&f�A��[*׃B�<����X �XRG�fdT��q�E�<9���aj>\D>A	N)�#�}�<���4m(�`� 	8.A�DЖC}�<)d���O��1c �\�pnڨ����q�<9�j�:*�i�+�m��E�iVS�<)¦�k��i�˜���L[�YJ�<!3����<a�,]#BNɲe@�<��D#0�$�#	:ySP���a�y�<�1WOF��R-!'@��Q��^�<��*̽P�q@��+kT:A��b�F�<awkZ8�-h6�/�^]�l�i�<y"A��O�|%qu#��@OPi�<�G᎜�=RQ�ȊgtDcE�Xg�<YP:	la��μ\->�fe `�<���ڿ=��I'ݰn�&= ��B�<)"���B`B��K�1� ����f�<9�៭k{�U���	H�؛�hi�<) ��#F`t��i���Z)�!�$�e����
�".��C�L�#�!�$1\q�p �d�#�5{Q.5v�!��Љ|�#�ы^H��vKd !��H��၅���x�%�r�!��3��M�2`=�0���!��Z�`�J��F�D%��+�f�M	!�d�4~�T�Gn��n�b�$�/�!�M�u$��A��+��	���
�!�d�$�*�"��,"�p25a5p�!򤓗c����H�3rhx �	;7�!��&q2P��k�h��2�>h�!򤆊8�~�8V�h~����J%b�!�D��a|����X.p�����M�!�䐴[�6iӱG�_�����C�!�d��e������ɻ(� �5d�oz!�� *�s'�I���r�;G;%"OT��0N��4��)�kP�,#��B"O�a`�N�E��9�s��
h��%�w"Oz��CM��ZG�5i�D��q"OheS�a�h�;��ѝO����3"O&��vL]�S���]���	�'�Lt�Ucɫ�͠�⃶�$�
�'0}X�l_'�<A� KI=39�A[�'��IƪW�yh�:�.ڲ-"�'k�H�3NS�3j�Ip��',>l�'X��٠��As�xZ���/%�:I)�'���G�>(�pK�O�T���'Wxdf�@�ÆJ�
v��'��5���"/��h��X���x��'w�͂���&*y�|A�BN���x�'�
i�8cƤ�4$�x�X�#�'S�|+$B۷e~�@C#Dv�"���' ҝ�n�$0ļ���
VbWf���'Z����*B�6iF)a���^t\�z�'G81r��;F�z8���'�x9��'�>� �(C�V���Q���3�a��'����5��L�FaZ�-����
�'�V�Xc�m�l��g����
�'� �b�5DG�O��ʴ��'�Qaw�:�0�R6-Y�B�ص{�'C�Ic���N(D�RT��5K�he�
�'猹b"M�Z�mZ�a�Ffjx��'��X���|��xbA�%;��q��'a>l3#,��t6j������8�|��'�&b%��$0N ��J>G'p
�'�us Lʌ3�t�2 [�,����	�'�ZpHS��H�Dp'��/�,�

�'������[�(�+��� �Nt	�'�f	y&�O>mi�	R!O�-�0�	�'U^�X�8��$֦�#�A	�'Ƙsc�	�v_r��e/y^<y�'��dK�cц�ps�m�4j	�'b�-mD�Iv���sd�%R��2	�'E��[w��)��ᗍчl\���'�$]�Ώ,4�6�aP���٩�'^� :�IP�R�\H�V/J�o���`�' �K@��'���q�^{�P�9
�'�6pr��'����9l�%�	�',4 )3!C�*�8WM�1uK�1��'�P�8�f�6+��$�3kŞfTH��'y&HZb#�]80��i*coL�i�'�.���ŕy+h�0���.Vj��'� �9E���vԑ�"h,�>�:�'P�}�"�Q3������x��!
�'����)Rn��1�IQ�> p�'�8��j@'VYM�%�/	�r���'��QxW�\�4��aq�̞o�hy�'x�x��lU�p�r%���E�/�#�'&�(��5۬h�%F�)m��T��'"�l�� �=�J P\�$!�'���U�I���5#'���
�'�2�{�MCb�e Ux]+	�'
�s�	�6r�2�4� �⥋�'���C�R="�^%���U^�	�'L���J/s�nY�#dD����'�>X�s��j:`�#�&/(�� �
�'��A�(Θi�4I��_ L,H���'�lXxV�N�_~��+�QI���	�'�rp�$IH`�����!B�TM�	��� �x���[@Ru���0�N�`�"Ov�Ң� �q���C/�>����"OZ��#Jw�� �(�/�X郓"On�×'ʪz�V�b��LmPAp&"OV%z�M��:�T��P+����"ON:C~I a䉛)-���"O�吅$�;]APؘ�'�����"OL�cbC�g.��K���'P����"O�0�n�}ԞЉ�m�c��|�"Or��S����$���M�<��9�v"O��(�[�|Pɢ��u��!8�"O�P���G
�,��*�<��@"O���5�V�(���jU{���3�"O<��"ȉ_��D�f A j6���"O��p֪?9�}0U��<,c���g"O���C퉩�,R�LN5f܍�5"O�d�&�ΗG^h�FKByv���"O8�1$�xu����t�7"O0�k��V�lPd((/q�hcU"O���آ ">A���>���� "O>���$ؕ��YfgÞY�*5s"O�4��K�:�c�"q-�Pi�"O"�6�Qrv�b�g�(s�Ҕ"O���faR1��(1AY�!�6�8g"O�Y3Dk٤4jl<"��)R�t� "O���S�C8�4�1$NyL58�"O�Q�R�ٯ�S��v�<K�"O��)'���4�	��9L�th��"O�]�!�Ej��EH�|}��"OfѤӭ��q`��wPh0�"O����T:�|���m^�Si.m�S"O4�E��x����̋�_J�0"OX�RU��(C�jg+�;G��4"O����Nå!����f��t.�j5"O&X�O��eM>	PqC�=jT�%"OpU�c��;�����>%2j�"OD ��E2ZU`C"܋ �a��"O�<Hӭ�$t |�[ ���ȸ�"OB�Q@(O��0�H��O5�QA�"O�����G�{�]@�K�!0e"O�t#A��}�Vh��h�%$�*��"Ob[ ��?"� ��%*F!*C�M۴"O�9	tc�\&-yg��6Ӯ@r�"O��	�eݸG�0�c�H%c�8�"O�X�\��� Pa��+�>Y�R"O>]��*�:ԩ���G�4����q"O�FжJ"�	7����"O�h�"KH(�<����r�&q�7"O�$:a�4�H���@+`��Ac"O(ɩ�U��ݳ�
�?��Ԣ'"O`�j��NvL8�bI.�L���"O���c����Ua�� �����"OB��ć�vN�A�R8x� ��"O0DR�ҤM-X<�3�	�/$�{w"O0�@�摴8׬�� �]�,��d"O�:Q��N
Q*�_�yjv"O4�*�H�)0����:_��L�"O�9B6�;B@5��rV��4"OĜضIU }�2�3�pm�%�"OJ��D�
bP�)�K޼5S�U�b"OvŻV��8�
�	�݆q2j�SB"Od����ʤA..�*G�`%�()�"OzA(B���0̲К$@[�(vpR�"Or|��b��B0��*q�Om���"O� \�C��k���:cQ�7iD9��"O��A�E�
�)�o�l���"OPQY��ǵQvμ�c$��b���"O`!��uI4��6�.H�:�"O�h����Z7��w�ņ~��̈"O�0#"��G�n��W�-\�h�"O\d����!{>nQ`İ�"�(+�!�Mm�r��� x�^�����M�!�C�rʼX2�
2?Դ@��"r!�ċ@܄�p5oI$g5T2�%��Q�!�$�JZh�㶧[.(}P#��3�!����\:��S�ŚH����7.�!�$_$dj�Y�OW)i@����\��!�$OW�x|9eb}��i��3�!��!��h���D^�Kp�
%�!�Ď���d�U�܄fMyҥ�!�D2*p�aH�@?W84y��ݪV&!�d�4���Pb�q:�!��ٱi{!��dNX}�Eb�(IRPcw��
!򤕫j�KVE��a
2,���&!�$;Ԝr�k��T�Q��Z0Q�!�\�25���Jha����P�!�P�*~-Bv�O�}S�\ QK��w`!��X�Rq�N�`2PY��Q�9!�$/NPl��W�K�^��03c]�wu!�DǷ/���d,�O�"����/m!�$�e��u!3I��K�rL:e�T�d!򤂎#�QCׂC#�Vѩ� �`!�d�+h;�B$�Ԣ����v`�@�!�Y9*A�Ң��=�^A��)�!�[$3�n�JG&%&��,�a̅3�!��Wd�(�%��\��m��T�[�!�$ѽO��=���٣a�@ēb+̋B�!�B4#_:���/0�����K�{p!��@���� w�+�5F���jc!�Z���m�8��A�o�!��'Z����ŝ(H���%�K1g�!��r��iZ&�[=Y�~���
;�!�D��.:�p� �ՌL3�KU�@�!�]"�0��[�R�f<��L��C�!�$Cy@�drD�N�H����,��>z!�&lg�b�@��r��P��j�$ie!���9n���1�ď^��i�Dɑ�o�!�DA.*��0ϔ`P(��55�!�=�}�+�u4����1�!���-f�6lq��	�\-J=���Ɂ$B!�d"��i��H��NF��cf�*2�!��.����,
 .Y�Ñ�M�+�!��]�&�`E�RuK���C�B=�!�'
�t�ĤaG$�����!��܉_�ޑP�-^2߈����T�u}!�d̼rڰ�h�Viـ�Q'Ȫ_W!�d�?5 "!��ˈB��@���ch!�$��J�h�`@��[�R1����/@4!�'��}"�	z����2��^�<�cF-�B	���l�����X\�<�ԭZ�=`1�/�8Fln!��U�<�D�f4𥳥�7_9��/�S�<�˂H�J�pG�����D�P�<�'XL�����PK|�RV�R�<��3[�qz�&]�E꓎�F�<�r��;/hIȦD D�pY�qnC�<飧�9B��"+�#�����N]v�<1�,O�jXp�̉-D�=5a�n�<� Dc3L�b���Sv��!�E"O.���I�+��[ԭ��"��"Oqct��$.fH�Xc�ۡ�xE�"OR�[�d��j���sĥ�
F���%"O���A��	4�4�dS�,��y��"O�4�f���@Aμ!ЩZ&!~ڸ�b"O	za�2$�r��Ǎ
���C�"ORqJS��(���T��c���""O��a��s�R���/8��-��"O(i9�fӯ	4(�0E$�$ �N�A�"O�d�Ң�1b�r8���6,���"O��&���fo:�s
��P�4��T"O����gIO:^�z����a����"O �C�_�Oy���$�[�*8`H
 "O��c�j�ł6	^0/3���"O֤ F�(&װH���m-p �"O����eP�K	��ӄ^�z��D�B"O���wC��tMXyid��Bf��[R"O�J��K��$��E�lc�dqW"O�Q�f��KZhh���0c�iPc"OX�cWgܩ<�{e�F}����`"O2��2JQ�	�
D�PH,C�r���"OE�O�N�0�*P�T��̻"Oޔ����!�fR(9	�a*�����y��Oexȇ��-4�N��O���yb̯g��-� U��A)"�R;�y"�4�l�7*T6�~`)����y�CA�D�c��(���տ�yB�X���X���"K������y��K��iX�́Dz�X�AK��yB@ �v%yV	 �:2Ir�";�y�lͬ_Ϭ9#AŁ�0v�,{p�@��y���=���넭!>�F��L��yB���u�����AP
4-t4��,φ�y2N�7u;n-q�c��+.��!�F���yB�D�K˰Mڃ@�*%`�qcH��y�c�-()�b�9�2�A��y��O�V��X�A��	��22l�<�y҆@�<P�bH �A���ξ�y�ȑ�Q�L�KQh�3�ҹQN3�y��ڙ%&Q�q�Z�)`@�&튤�y���1��eGͭ�5I��
�y��Y�H+����P�.�8تgk���y�i�',.j��V��R>Ap���y� �D�E�D(*�0�	@��y��X9��I5/��?�@�C��:�y���g�����
�L��H���Py���v�9����*� ��I�<I���KA���7�/P���A��<�B�
A0��J�|Dk���~�<Q5�ۧ>� �X6ˎ�]���&�Sz�<���K�jZ��iƌ��%�EHx�<Y��1eZъ��ސ|Oؼ�0�q�<������(`���N!���T�<�닔~v����I)�Pq�j�<�$-W9#�P`�A
G���ҋPc�<9q&�:Jd�cQ�_pC(D����b�<�d�M`�8� +A��*��'�^�<q��h?�Hc.��IW���3FR�<�w�Fi��mq6�[�*�:ّ6�z�<y�^�Y�-(2� �qDg�w�<�'Ԋs$6�r3D[�:�ʤ�e��w�<�敞TXJe�g퀵c�.@I�<a#��~B%P@�5�0��\]�<� ��A��$��Ԫ���'�����"OF�� 훍b�z�����C9�y�p"O�<�Î�2c�L��C��M
<8V"O�$��mӋF5�P t$Q ['JE�"Ol�aD&ʵjL)㣢t��1c"O���b�8Dr�HB�kʹS�"i�F"O :�@��&�x�U�L{̤s�"Oޘ��*�vA��Dп
0��4"O�1�`�M�jq�	0�<��"OH ����V]	�@,W�H��"Oި���T�q�R-"@&C><�
y��"ON��@܇ �p�dEY�"��9K�"O�M����/�H�X���{t�Rq"O��ʂ��-l�|�0Š�$,�Fp*�"OLM3'� ��8�/�<~�բF"O�����5m$n�2D�jrPQ�"O��1�G0e�`�D�1>S�T9�"OPe���Z<E�Y����!L|�b3"O�IUR�!�K�+@0�-�"OF�*v��8O7��;@�A�yOx��"O�;$EZN	<�㓫�=v�P�"O��T'�H���[aʘ'>�Ij'"Op��!���q�@#�3h� �"O��b"#7y��!���3,<�"O�(�LD@�2d̒�f�q+�"O�#Gӯ
N�u&��l�t8ذ"O8Z��Y�6A�;���f
yd"OvP��ńr�pE:2h�+Z�&("O�QJ��Ov�$����T;$�Z<٣"O��kW�,C0��7'HW�8;!"Op�EG�=�nA���Ԅn'P��"O���6�3
���ط��}����"O�(Q@aU:-i(�Qֶ5�:�%"O��b[7h��"�Ɖv`��(@"Oшs���ز���PQ���"O,Yy�ㄔ��ܢl�5-�x"O��c�nC=�$��s,٣1B��)A"O���C�We�0��*��W)n��"OL���� 1(Ȥ�A% Y�pj LJ�"O�œE!!$Nё6�QaG���E"Oh�"e�G4	?z���M~]�"O�-XԊ	�)�D���W�1ʰ"ORE�V�خG]���!K�����V"O�Ÿ�bѐH� 	 *��o���S�"O
a� ǦU�$���Pd��#"OFm;gi��)�%��Ѩ]�ĵ
""O�@'���D������"�"Od��5�d�P��.�`���"Oz�y�i��SQ���R_*`)�Y��"O�}9�\�j��#��}x�Z"O��4�̆�~��)ԔY���"O�Qم!�
�� (�<�2,�"O�I!n��:��89ņ
�v��"O^��eр8P&m���3C
���"O�y2E�I1E�KP�ע6<(S"O�U�Ү�Gh���E� G2�8��"Oʵ#��Gn���/R�f)\Y3"O�r7mI�;W$xH�'N�|��Cb"O�Y	A �s�e�C��	���3S"O���7�}|�y����̑y�"O�9�r�%7qR� �DÎ��@�v"O����8XY
��%��U�}�"O���`�˂*bؕKԤY2H(�;�"O�@ۑg
�= P\�I_�Z#�\�"O� ��B7*�,@z�������4y1"OȚf�B1!Ǹ�����a �e�"O�{%˒"�M��sW�[6"O$4��F���ɰ��_�`9�V"O�ؤB��N�\����@�o D�+s"OXqZ�,~�:�ja,E�d�YP"O�\���T���GaS,0l��Y�"O�� BH�;>e%!A,$�!��"OpY[��r:����Ņ<wr�i�"O4�C�++c�� ��-�u�$��"O�$@��O>h�>��"LTxs�"O<�&�	��K+�*b$@"OЙ!DE��q��e�s�=r\(#R"OL0�S�N2md�s,ai~�`"O2�!t��5)��R���yW��KD"Op�Ԡ�M��`�M�F�a�"O��)��}���F܌HR2���yRLS #j� r��G�@�J������y�͎���yz©�� P� �Ѡ�y"#
�0�.}�t�#�r�
����y��Z? ��Ui�d�$1w��d�D��yB���(�pM�cg�/p&�*��X��y�_,4Q�HG����#(!�y�?6||ztW���h�c�%�yB�Zz�&�A@R�o!,�Ї ��y��T7N��ܸ%�>S:f�;��P��yC7f\�h�ˉ� j00�eH��y��U�3�P�RDf��!���y�>Z[R��7�Z�I�l�@���yr�I'y
:|!A\�I,�shE�y"@�4!|�D0���Fl)��]�y��ҕrN�	t T9M�Dz.�:�yB�ۼd\� �c%��
�mpKқ�yB�,P����˗Y���%*���yb��(9�&(����K^�h�uo��yB��$�� �r JT&R�!D�G��yR�P)n�b��R���F��yb�B-��`CƴAczp�&��y��I:+�`2�%[�H�� ��
��yr @�6���k(LC�ԡf�J�y�ĲF��$y�#�����z�� ^�<�v�@�. �a��uB"�P�<��ՙETd����!�)��)P�<1 ��F�	�@�8�����K�<�7l�:{|$y*AK�HY�u��E�<���.y���IV,�C��J �}�<Q��,y8��!ߣL^��*f D�<U!ɽB��aC�ҚNST�B���[�<�gƘ�O]/,lh��R�~�$�ȓ&���c�L�&5�Lq����꜅��|��H`�Ĺ�t����[3W�(X�ȓ�2�j� �D1� �A,o%��VDJRg�&���`�#ߥ/�湄ȓC6lܪ�푸(_8���B#up@e��&\���q �5�� �AJ��ln����k�L\�VFW9FZ�U�6���n�耆ȓO�
�*�m(�L ����*�<��ȓ;{R-:�M�]4�0��H�,��ȓQ`x����|޼����g]ȑ�ȓL
�2�+ͷ /P����O)#�I�ȓ5�V���(2�Ρ0'$^C]H\��,H�1��B��vܙ���-K ��ȓ.ȩ�b�X�H1p�J֖/Y�9��Ig4q���T�nLR�K�B۔9�� ��S�? ���'`�4Ri&���A��Bf"O��S��ք	��1�n��(�"O�i�nI$	a�d{�A M�"902"O��(��L3c�X�a�N�VL�Xh�"O^<	��N�Y �%:�L��Y<P�A�"O�t1��Nت|����,c'�x�7"O�-���D�d�Ҥ���m���;�"O����W&_���0K[�o���1G"O�,zL^�J�F93P�)7Bi�"O�h�'d�1|�TR7	�T�� E"O�q2� �J�y�hG�v���@"O�ِ��;H���K���\�F��"O����e߯pne�d�O�z��L�"O�\"g
�Br242E�w��5z!�ݿCI:���+
m7��Zc�ŝ
�!�$����B�4N� q{�c�!�D�V!U�o�4 w4�{�"G&}
!�-2����w�ә]dq� đ�V�!�$Z"!T�Sg�gJ����m��C#!��#ӠՊQ�_$� rLX�\0!�$&
x �x��AF`<҂J�bA!�dJ�j@�8� �HtL�=���Dv�!�DԳ &\͠7hH�q74��C�Sg�!�Ā��(� ��X'4#�q��$(�!��K�����M�'D��1�VƆ�E�!�Ā�l ��Z�J۝9�\��3!�D/&��҂��2,���	�c�oW!��R	! ���Ռޥ@�1WLW�-F!�d��_����J�O��*P2VB!�d�61|����3��R2#�Q>!�DZ���@ U�+������^�!�D�46Dt��B9��yk�� �!�䇥K���G-0	�tI㫊�P�!��tD��-i�<�c�Om2!�w´㤎N��*�*v!�d
�;r�<i��G���3��T9d!���?�Խ�bj̄��ۢM�(p,!�ɺo"@� �	���0AC#P0`!���:O|,�����5U��9�Vh�\�!�~�sD��?���uA[�5�!�d 3�^���08��/���!��L#-��%:2�R;	(>)�l9:�!�D߃z�J���bK)Lj��sd���!�D�"��� t", �\ɳc�mP!�d~H��AI�<��p�)��J!�D�9i�wEٔ����2a/!�$�
h��I	���Q�04��֢C�!�Ē1*�*0k A�!�d�$g�<l%!���%8� H
f$�+�!�BH�!�dKm�`�+��7`��%2���[�!�	���W��"U�$q
1GD 	�!�D'C�u�#.w�����}�!�dQ��8�AO�z�6�)w�&5�!���lD2�ç��ab�0Af!�$�ޥ���3�J�o�3ޞ�Y�'�&!�,�:��"!2�p�
�'x$1�ᮕ>>#d�PFW�D� p;
�'G�2��Ų��y@nԱg��[�'B����ǲM����7G�h���x�'�V(�eK��l'6aӦfV�NbhA��'y�����-Z(�P��Ţ=m�Q��'��{P瑮y'jQ��鏸2�Z�x�'��a��Ǟ�K���f�+2��(1�'/dM
�P�a����/��R
��� �5�/�$�,�s��Y	ZZ�Y��"O�0x�'
;?T� ���4�L�5"OtA����QumӏK��F"OD���ȭV��bl��O`PA��"O�	3� ղ��釛mo8�"O�Lb�g�:X��A1
�643T��F"O�⑫F�J���ah�/�젒"O�!��&
xJ��@�{%�D("O�˔�<���PsF��
�:7"O�,�&�,h�A��
�ͺp�b"O<u�'�5��1P���r��4��"OT�%�8Kl)�ÁW� ��8�d"O ,a]"$���A���j7"O��ȡи�`���(���c"O�)4F�0D�����)Q�L��A"O�Dy1.]40�~�)A+ �R���"O����΍!k�ػ`�� d� "O�p!d� $��P�\�;Y���""O`a�SJ��Tc��bHFY�"O�Ijp��lh���T>V��%��"Oh�^	�4R2�Ë ހ 	S�<y6�Ae8� 9��x�h����y�<)���k�t�� �مPM�lҠv�<�B@�6���&�RY�Z���@Z�<9V�-1SFIa�&��{-��QcE�X�<�S�6���g��U��}q��T�<i���7M�61��A�� ���BM�<��D4�x`��1���Pg�<��`�i���_�`�/I@�<���t<`�� ��E�r�����y�<	1�17����B�傄�s�<�4B\��>��x�̝��P��pC�;1�VɁ&N�����kK1�JC䉹G<�
�昏'�@{��˯M�C�	�[��\#�Pj��C�l��v[�B�	#F<,���@(S�����G\ �B�I
>�)EeW.=�`��ˇ��B�I���A����I��t��L��C䉂~#<�J�a��I���f����C�I!d&Phc�2�p;�ܿP��C�	�Q#8���e�\V��Hr�=f�C�	23% I� �:G�����X��C�I�v����f�4^�	07��j.�C��#�0����JcN� �B�$�B�	�ke�� F&�lv)����v��B��6m+�\�Ƈ^�,y: �q)dC�	�E�!���ѱA����Z9>��C�I0^��3���:���C���"s|C�	$](и"'Y�5.X�a��O,[P C�.�\m0�#� ?t�BuIےZ�(B䉨)�H4�s��
F$a8燕)1&B�I�8]�� �̌��8*Q�֑N�\C䉺B���)���l༰��Q.3u`B䉰Jk��3�A�(W;r��d9?�B�I7jd�[��Ȟe@Q���m��B�	�de�\C�h ��dŘA��Q��B䉴Pޔ�#gė�0A�����(hzB�I�HdV@af)��4�,�9��ڷo>>B�IZ>�1�I�eU]���X.�jB�I&�48rP��z��<��׭<ȊB�	�-�4x�4��X���r2��a�tB䉬*�IH�K@�Q�℩�R�'VXB�ɰ�6�ӗ"�7��dK�N5!�DB�I�q&�`�"FT�?v��Y��D3(�ZB�)� Э[�j* ����(�dA�T"O�ш�b0�q�Уԑ5��i[�"OƘ��ΌA�j@R	�٠а"O�<q6,�����R�H�E����"O��h"�+;��1��
!�l��t"O����ۜ$����4c���3`"ON�`A]�[W0�!X_������b�<	�O�*F�8@a�5��ڳ'�f�<%œ�{	�UA���=^�Ų��\n�<I4EJ�}�9ѣOA���j§Ph�<Qt��vf����ō~��M��d�<��O\*4_h�Yr/���<aĘX�<��,�< ���ȼ��&F�P�<1FOW=|��Ԩ�'��/�Z��)�K�<Q�)�-�����V-�N�z1�O�<	��[_��U�%�M�Ȉ%�J�<A��;=WD!�unZ'�B�d�^l�<yC�@�NLr��!���pĉ�i�<��Cyʎ�Q�� @���8kJ`�<�Հ��l��,�l q�������R�<!V�;|Ɔ��C�tU�y�U�R�<��Ⱥ!�h�`��W3+���2��s�<���b��!���zxB����p�<��IR���N�<+N�K	�R�<�G��SP���$H�u#��S�!Ht�<�2O����F��
~n^)�f�q�<I@�]e�Q"FZ��U�Aj�d�<����,.�V��%We4�ҁ3D� ��
0~��Q����ö�-D�l�௔s I��)Y+4CF}c�6D��j�@
<�H�r�� ��S�C5D�PQ6���^m�C�oV-v���Z��5D��9ANG�X|�+���� O�X��,3D�T�������B	ݮDKWd2D��
׋�`mR���8��ʖC/D��YDъF�d@y��K�`9�1��d,D�d�h�";L(`�%�O�r18�>D��s��L�(`@T��˔z�&�2�!D������`�:̀ࣔ�W���5#D�tiw,��RS�!�n�&#���K D����ǉ1������Qi��B 0D��¤��@;Xʇ�O�9s���#D�D�I҄"�ʥ�uQ�f����H!D�  ?�vU����p��,a�(!D��wgԜ��; A[�I�F}�I3T�D�0*C�Y(��.$'6z�"O��R��"�����
F
M:"O�\�gKT�i��?U#�|!"O`HtfƏU(���0��%<.x���';챙f�J
$jp�fL��@�h�'PJ��WB1Ld�e�J$ ����'!�Z����hp�1+�{^���'��(S`i��
S�`��m���*	�'�`�{�#� ��A��N�k!����'R��BbAA0\(���e9(}��'� 3�Y'!
��V��
\��ē�'�9SPE�:����H�6$/(e��'�05'��k.Ԓ�o�_ބ��'i\�8��)pB�n%��A��'[dg�T�� ��'!��`�'�P*��R���4�`��6z�9�
�']\x� �B�՚P1ao�YzV�{
�'F���cb^�Vc�+�O�O
8�	�'
�K%o�828L�WeF�v����	��� [4� $�5�s��1"�c�"Or���ə"X��e�c-S75�d�1�"O�����y������c�p��"OF�K�d�4��ɘ�D�V�h��G"O�CI ,�4r�Cնd}��r1"Ot�)���MJG�Q:0n���"O�a[��9oR�;1a�3O��S"O�Pp���	ĄX����WG�DB%"OƩ;�b������=%�
�z&"O� 0���x~��	��=_�:�2"O��s���j2r�bA$)|
A��"O��Cc'�BeT�!3LɾI	؜y�"OHH2&�~���sWKO2�����"OlX��F�
�HH�QJN�v�by��"OF����/!x��g���&ЩA"O�r��4B�:�F	|l�ͳ1"Ol�����qV��Vlm��"O�4[�A��^�lȨ�Î�"jn��"O葂�R�&7ؼ!���N,�sU"O��ʑ�l���	���2L��=G"O�#�E�p , {�U�^zR�˶"OHy��l�8Ƈ�`C�<�Q"O�@�%R�[�hU��G6�q"O������=V� Ug��)[���"O<)SPb�gtm�2g�X��g"O
7�;J��KGWr�H��%"Oh�Y���>/���Bv�@�K�~Tx@"O���A�!L�qU䑊{����"O�M2e'�<�R=��e��� 3%��|���	�C�x�d �8[<;u
)���)�O ����6	���:feG4@�6�Qp"O���P �&fA��Ë�x{�O^��HMo~�  &�tܒL0�'*Z!�D՛<֎1Z���#=ZȲ����/�@��ȓa�� ���V&��8�G�!�~���7 t*1�H�w�r�$� G-�l�ȓ�4��e�T1�hYWO��<,�8��~�AN�R��a�SjԉRSh���	�Gz�	�bײ���+G̜�A�  }��B�ɚGg��A���.�H6�%,P�B��-��c�j,�Vl��@��lP	�'P"��!KØ=� L�b�9#�'R�qRDE,f�y��K�Y���
�'���j�Κ�g^L����S{�u��'����W3H�#2o�P����'������2
�*�@<JLP�'���;m>��÷FUv���O˓�~��ƟLF�4`���[@(^Ě�S����yb���
F�`�q�ǷO�9�S!���'M�'7>9�B*�#E�J��d��{��I
�,LO �'t�d�f��x��.�h�@;T�>I������0�0�8�g�O�5J��Y :أ>i���է+9���6'М2�.���H><�!�$��a=2 �6� 
m�DM&�J�v��+}��>%>O���!�xİX�P�,:�Y��'I�I�^�q��ǃ4Rv�A�mW�c�T7ms�X��>9�$q�%�T���ֆ7k�Ї�	M��\n(p2��}nu�4%��:t�����rFH�.�� �so�(�$��������󤋵.	0�B��nT��oP�=�!�$βq��@��͇�h�aV$?U!�$�8��"5�#a�T�#ω��!��=`t4���E��uڌ�oY�I9!��H�q�Dц�΀��բϝ<}!�� �l�'a�#O��1��Ӡ=�l=j`"O"l���G�:0� ���	H�>-Kv"OQ9���h�����*Tuب��"Ovh[���H��Ƙ�g�`"Oڅq��Cz�^�8PF�$:X�e� "O��§ �����fW�K�H	;�"O>�q�2<X�0�Bc�?nԮ�S"O$�*�-$�꒢֐(���>O��=E��o��C��	������7�y� ͪy������ƀy�&�ɦ���yr�;fc��+��Y �"��F�C3��<q��9^P2���^<R@��(��D�!�P@pت"/!,��pDݐjV!��9HbPBB��#�%0�O�ay2�'.��'��-�e��� �eK�:��)������G{J~�H�%*�N9��%��<jDl���U�<iVC��9�r��#NS�n2(�4oUP�<�G&��%��dr��� �ʍ�f��J�<�ACX2X�0U�D<xB��H�<i���F�@P�DN��,pR*�O�<�p� �}K�a���;��-��fI�<1f�4V`x"���qlb��V�TAy�>I�~S�@�r��3��K3`�7�8ȇȓ,�8yK`�j��D���4DVЅȓ|��X1�ּ+��Iץ�����>��'^a��!F�E�����X$;j���h���y�Ӳ.�"{�퉾f��	6bW4�yR`��oQ��Ŝ0^���d͚���'�ў�����}��:UO('�4Ī�b�� ��ɩΐ�C�V1��)!F#P��$B�	�vFh����>Gܹ���XO��C�������_���9D�E�JݚgN-�I��4�?�N~u^3����G5PE�D�Z�<��O�"��)-�k(��Ӥ��R�<!@M�R�@i1�@7DU�i�� CP�<�g*�� �L5r �F��B]K@[��xr��N[�I*���X00IB���
	�'���Xq/�"�Pɠ�אLj&hC�'�Mۗ��?m�y��ͣ�ź�y2�'�Raؑ��Qb����?W���'�r	bJ��A.����I�`,B�'����p!�m�d��`�D�$la�'<��wA �UWȴ��N@�\q��'���� ���������QS/WPg��<E��'�"��wd9/���w�9S<R�'yj�"��P�:eI�-R��y�O6��$�.0�y�Эf��=5Ě�w�!�D�&0Z�G��(4�x�#�H<!��8Y�f�PA^g�RM�F �I�a}��>�5f�Uu��9 0`PE���x�<��J�{�|�sd�4v���A���y�<A��&\0c�j��K�l�ԧ�t�<�uѮ	�U�fa>R�$�G`׭�hO�gy"�O��$�/�$�
�I�d��*1#ʽ��C�	0q>�%{ՂJqar��FR"p�HG{J|�(H	Ul4q��%�a�`��B$�O˓t�NU�׹GU� ��)Q6v Ez��'B��5�ѨM'������H��
�'X:HpE&�.7�^��dJTNdP�4(����%~^>т�	BV�D��|*!��6"OL���g�s�6�JlH�h01��qމh@Y,��c�Y/@�D!DxR*^`8�tI��;$��e��|E���1E D���f�S51¼=�bkk�)���3D��  �*E�np�	�H �U�BP*""O�P㫝}5�9	����$���"O�2�-ʻ_:¤�7� Jèe�dY���A��o�'O��a��/{�z�ВPTR@y:	�'�ؕ�V���F�xmq�(8I^� ��O
�=E�tI?��0!��	0N���Т��'k�`V����A2���V���K�<���cџ�yR�O��"~Z,�2��#O\�9s�yi� ^z�<Y�@BR��Y������hO���<��nX�A�X' �Bh|�������<9�;������Z�pLxtf�;��x�_�"G��%_V���I�+��O2 h��IGh�BՊ�*� W��APLP�p�1O~�=�O��$�=�$�E �'�>)P�l�9�!�d�$<��� �"�`y:`I��l�!��@�]�T軂#ި �����(�<�!��+x�;�L�{���WW&:��IEy�\��$��'�� ��χ���y�� ?�E��'S�T�2MF�+�����R+L����';��3"�@���5����݌pi�'%|�q��]� \����|P|��-O���Xm�4ب�X1w%�T��@�%�ay��	�L>�sF�%,�@,��J# �C�0M	��H"/�SZ���@� w=�B䉸[���E�({Ȕ���mK�T�tC�ɂ9���D\��v�P,˴�B�	3�t�
�@��$n�h��Ό .B䉀~��a���F�S�Jp��c��L�B�u������yx�VnХ*~�B�I[]HԘ1mɏm�R�!6���aoTB�	..Ez聵%� G�õ�%�8B�I&`؝
p�K���A���hB�	45�*,�qoB� ������`Y�C��U�xK*�=88�[r	̻1�|C��#3d�r�`]�p��Ș���}�,B�	�G�Zy#�
�
3 �754C�Ibw~��
*��6��]�@B��'g��=R1Mȅq�:9�DU$M6B�I�56=Xk��U��*uh�0D�4B�	rN���1e�4�B�c�*̛7�C�4v��<Ѡ'�'[<���/�~�C�I�AL-�R��38%#˂9�C�IC0�����,7L8��`�f/�B�	�-zL���!�R�Aa�L�jC�	�H��६�D=N��'��s�B��������[H��(��B�Ɉ������oa�P��M��fтB�5�jL���©$��#�`�34�C�	�<��xHV)�<~�@�P�*:B�I=Ptp���ظ`��<z'��}�XC�	�q8s-֋$3@�0��H�o�VC�ɪ6�ʥ���S#f���A ǅ\oHC�	.Z4@s��!���K�!�C�	�i��B��>���[����.�B�II���R��N�nmp���f�B�Iiؚ��Ed9N�R���D+:�B�ɲrNN�";�(��t�6wbC�	,<�� ���شU���� �B�	<Y�*��䂗�@��Q�(�0w�B䉦s��Y f���\����J�B�	�Z.�� �{�h
E#��t�8B��y��jnO$�lHb5히;!��釫�)a�����L���,�=�,�Q0f�?|���
�'�0u�v4�ě�@��s�\ �
��� ��1MX�h,�IFW�Z�fy9�"O��3uoҤzwb0��.��	�p)�F"O�4�	R�\�dpj�䍉*^LZd"OP���aS�)��+e�D4h�$!�"O&��T�ɴW�⥲b"�r}l�!�"O޵�P�@8�Ԙ� ­6N��S�"O�h����9u� ��OF�/NN�i�"O~���↼5��,2�5]BTH�"O����js!R��el6+�0
�"OR�2&�`�j�a���$��II"Oҡ��L��{�����˪:�H)�"O���C��=�Z�����&Q�J�sB"O<8ac��lX��e
f1z�"O*��
��xv��1H��%z�"OLi�"��n|���c%�A�b}��"On���,�j}:��re��l#PH+b"O�p��h�QL&l;GAˎ|�e�2"On���֍S�s�n	���Ahw"Ovx�t���*�iڄ�X�%�"8h7���c���'9܌�z��O��(���L1?�Tm��툭Fs$��	�sG2H@��+�@Q��+`�l Gd���I;W>��OgZ@5�B6Q�X��'�����7J�6��N�o�҉��t�.ճ�X?��B��V9':�ʷ��;a������O�ff9�s�ê~�p�;&JL?��Iܧ&閝K� ڍ\���1����E{��:d�,�F�ע@!v��)g@�IԽ2�IF�g���v�/u�J�ˀ�S�P���5B�v����L>�� Լ,���:B��: �=
WN˦���%�\�J\�7���C�کZQk���(����L4v8a[����胈#��d��46<X���9��,�t���wҭ�䏙�Ryˣi� M�&\b ��I�����v��	��1g"ӼacJ}`dM�Oy��l�8���W�]j٢��'�p�	���ąѱl	�ip��	
H4����'�J\���Yab���Ø:|pv����l�I�L2���O?1�0�h-�В�%�w�:��g�:qT؂ƒ|r��vD��fBO/=TFMGR�|� ��1�O�Q���2�����k����dA�Kw$�8��'����Ȼ���炍3�����@��:k�حۀ/�m.>���nă1�|�������z|�v�
o�Xx��ֻi���?��;u��Q鞟\s l� -J�b�Z�!��c��ɑ����
ը� Fɕ1��d֞ @'?�[!Ϝ�^�D	'Oŧ<Ht3QC�;���z��Ζu�NH���5>>#|�b�&p*��$
�,$ 4��z^���F�I��ؒ�O�}ȳO)'3<�$>7m�>��� bS��K��!�d���
�F����=q��ű��+�����*	��+7�[�(�|���?i� ^�Nʘ@�w.�"yp�r��= �|���2�W�T����2'S�S�	����+v��y��+=���#�
�2�� ԯ	�����<��T��LA����� ��=�� ���K&6��(ďZ��?���I�F��ƨ���Q�O[U͜�T�ԉn��\���6h��u	u�H K�@����O��U�6��WȖ�4��9E����5)ѴB�x��r�w툄k�)X� e��ǉ-/�i1�.�8�?���зD�l��BB�T�D�-^^xq4b�����5C"�x���eWD&��2��Z=��x"
֬]Y��H7P"|%�kƲ@Fɂ�+�4߅�j�5�\�i��!p#׶\i@���^����f^�<fM��y�G�<{��ص��H \7��q�(�
�b;{�YC�s`� aw�B,%%���7�I$@8�&�s� ���Z�y�yф�(7��h'��kp� p��٣[�%那�sZ�ܢ&W�\8�$K�9?�I��뛟 ��;v(ք�~b��P`�@�w��^YY$J�#��y��M�x���8���aI��k.�Pc�t�7I���xu�d �R2�9*A��8p�*FL@Ȧ�3w���J�Y
�g��YϚ)0Ac��2D@&u�,=�c�@�g����]�z���a��^�d�K�b.'���'��8^h �U�F?D,���jA
~���FX�|�b��%���"lF�e�N��C!bح\!H���.R�ࠐ��;,��5��j
\�R�����#���,_&F ����m��DK ?�y�QV(�f�� �Q��?��#ܖ�r]��LG	�3?��,G���R�٧9�0��?5P��,��,��mʃ�����U�/�J��"�&?�4�#���;?F��l�*,����"��wC�B�ɗb<Qbٙz#b�KwD�a����,ЋO���8��ȓX���C���F�0�o�
l� -h�h�6QD�adA@��f���ˑ�c��)�%�C�X�Gi�0V(��ڠ���-��1�
;H̼��ǃ����-S�UJ�:��z%C��	}�����&b�z��S��+P=��Ɛ 8>�H��kݼC,����}`9�C���K4�ۂ* �/O6����	l�d8�T?Kd?@c>8q���"t��1eC��C��]�t������z8�D
�Ck,!���>L�a�3gE) fGs���s�ʊ�8��P�0��J��>��`�P�HO��EI8C� ���ѣ ���v�A�\Q���JQ<,�b�H jSl�%��F�
���oѡ%��$���4XY��#Dd@"n��9���p-j�o<HF)���XԔ�����z �ij��	�Mǐe!$aR����hQ�ҥ^"����B �z�kΎ� I��B(H͂Et�����X�xbڨ��T�矜Oj9���ؤ�HO.k���Fh���cO�$����&̒�1�@M��@�'#,|�0�HL��,�x��ӛ	�m�bG�!�ΰ�1���<as�n|����AN�K"�]֦mʁ @�+���� {M����Φ��Ri@�����$�;-o�h�����/��6	���8I,���S�? h䒱��<ULLp���:*�0$���ƮJ^�S��A�옄�2-�l삑�<TIPHѮ�8.� 8�8�����V">Dl��A"�~��C�'�x����1oH�5�Q�@Wqzy�s�Ҹ+�.�������I�D�|�p�-��c�����m�([u�">!�h��K���6Tu��E��3���2&�|OH���OX]�1�a�S`�I4��rs��i>n���H!�Y$Sv�#�eG�:��
`�$ŀ�c�-8T!�l߷l�t��l��O>����5KZpABb���qS�� @��D(Z0�-�����X��LRUQ2n9�]`d�[�ة�+��W`1�փZF08|�u���#Z�G2:6��8�ri�7B�98�Z%�w��\՘%�A��'|&���c�5|O�t�'B���t�d%M��w
�;$��k�ͦ#OxH����/z�ޡ; �;��`�DG��ިv����Pٺ�@�/wJ�c��Y�?ດ��I�x��1h�@�c]�
�4P���(�ZQZGC��1�1r�(�E�,I���U�v0xS�i��e�h�J�'�,��1��H�1{۟ظK�>]4a���$��ۤY����ӟ4�Y$�_$HeH��#eԝ+� �!�.�A�a��9W�|�%�^�=Ӯh"�#��wmL5�e�_����
& ?|�0w�աET�t�5�>ғV�4M����^��E3b�7D�hY8��&n����k[�$��A;ԩT�>]�V+�=\��E�5A�vaX�mR&AG�}Xt�_ ���p���eEI�^A/�8��'��0b��C�z����RU�Q���V/:��꧈j�zq�E���z��CA�/}����n�Ӻs6)�5�M��4|�!	��G.B(�1c���4\�<AaJ(���4]�8Ei�'�x�b� sPy�k� ��a!OƍV
�l��>��0�Вcwf� �I'iJ,,�B��(i�`�(%�i�"�`@�C>n�5�N���V��0*pY����`>�}H����.��4J������;f$d�p��mN���j�!�r��f�7"zq��A��(�(
�,ϐM��ܴ$~\h�#���Ѣ�٦;J�y#b��E��$�|+B�F�D���ƭ8[3������-w#bM��Pi���˥��i���r'bVR���-�;_=���N�r+veh��k�,t�ď�.b���ʃMyQ�CJ�*]��AVp��ׇ)��Y��%-cIQ�IO")xe�2ɟ&�Q���,*J�8��"?7� h} ��U�ɟ�b\�Ć�I�%�vg�?�u���<p8�Ah�v�i��"ǆ����ӀB�AԾi�V�� �֣�YZ��@�k���B�l	"�h��`STn��l �Z��h��U&K4�T��m�(5H�a`Z,]g�TKq�?H��:q�i�P���͔n!���G)�D�.�"	|���Źkȡ�&�x��@�9-�\�oں����4Ü�8M�XE��u�4�c��M?��:7ʐ7@�͡�6����e���w|�$IS$YܦŐ��p�B(���%h��1.�r��L)B0}� χ8� ("�䚵>�^���R��b����!3O�M�s�Q<}� �G�
�:*�$�6;�R�0��5��K�n�#�\�A#�"�H�[�E>V��4"𙟔���Kx���9ԠR)3/rh����"� �W�\�y�����샹HR��0���X��4��I��l�(����ɍ������{�𕊦�OT��p`*P?^���	�cZ��*ģ�����["p�j5#n��d#�DX6��j{h�*E�3(Dn9�A�bJb��FG�/�MkfE��Z�����!yJ&t*Q�ɵz` �KN8�7����x�7A ���
�Z�:�]��H6-� E:\�ɕ=&E���҉a�!4��4K�R�3�$���2�Pf�>��$I�BqJ񌚣u�ҙ���l��}�0��?�*�ag���x["��H��� g�.p�r�T&
%��=!qf��1��D�5'�Gn�x:�aP1(þi���2�H�L�	�"�)oʅ����?%�U U:�6��7g� \$�5Y�N#'h�u��A)r%�Ep/O�F�+��B����0W1a�EW�4�ʣ�}#��C��g]z=i�ϙ#9p|��g�߯�j��7��1�+O��P�ᆛ�T�+����k��c�EK�'~��Aʔ�ո��戚05^�� raG��D��j>{åK
!X��6�S�V��lX�R�9z���n�05q�iJU�*!��� ��p<��E7%^�P��� 9y�C<VhcrAD�'n)����t�@�����������<�)X?�9�c�L<�����FE�N��䃞k�z�
׍sv�!��땯L�je�>La�#�۳�PݚpD�"P�@�ۑ ��=p�9��K�	E�8"�딼Fi�'���b��/3��3�P�NE�*���'�&tyEH�� �r�� �U�d� ��
�V��p����HB"�!J�pE[��z(�@�Ǎ�$0V�D/��$ɐן&���{��!�GB���uG(@?v��\�T��=KD02#���M���I�����I	Cj��� ��{�ZY���:1��H$&��u��>d��ōO����7���
��0���k�Z����ڈ|��H�4:l��;����w�2�� ��'�4H�m��V38%(��;���P �B��0�#ӃR����H���2@�'V1<)0��ށ:�����C:��Q�}P�E�W��Y��lk��3@��g�ٕ{28�EhQ 0���{�� ���H�I"'������_�3a�<"�"ҁ�f�" �� �<a��{2 � %��!�_ �C��9:�HS�'Oꄈ�g�nM`0 c��W�:�X��.ړ:%.ЉĚ�����!L�t�� �L,X�R�qJ	��PN������Ȕ;���  O@����D�ڡu�
��Tj�2R����΍VK�p��L���O�x�Ӭ6��x�e���X(�4?��aa��?�J�ů;V,y�c�3G�t0�`�+1�F�����5=��(s���	�ʜ��+����f�X!Z1U�d6�h%��gP0a̸�E�1^y�adV�Or�H�&̚l^��H�aT�Ix9��'0�&ªM2��"���2Y�zqV Y�1Ut\��1\V$���Ɠa�yJ��&X<ys%D0\�n4E{'	i���K�(Κ�De��GK�
~���o�=1���1���'ys�,�@��n���c�h��VM��W?m���$�A�Ē�
Ť���F���e���Д��O�PJ5|�.� �`�;OT���K=z�����_,�h�A�m��!��㆛�j9�%�4u�S$7��kȯs��� N6S�l��C��+"�X'�ݗ�"q'��P�]�(e�m8'��: bӈs�Y��8O`��1���~͑sB��C��9��2_\a��֞=*@�t�ٓм�QEԄ�z��BՋF�����0T�F�l6R��e�}ƠA���=�4����{^P��,�66j�1cр��>(���sv͚:�hT��4k�@A �/	B�0`b�ƒX�>��޴n+���A�F�� �2����!���E ���G`X�2��4��=;c>���#
x	�mS��"�����=.1���wP����O�	��i�r�? �DZ�"��)�$�Y+"敳�Í'$vY��Arܓ�*�����r�J5����i6	8�HU�R��s��m�Xi �P�E��a��*��v���8���k�!Вm�X0!����^�5F��4��uY���c����Ô0��$�?�A2��ӌWȆ��EL�}X�7m��N�x���ٰ4�(�Y 
=lgƕ�H��i�^��EQ	���Ff�8/�`���*�"76P`!ՠ>i`̝�2(�,k�T :��E�S���7o
��Ø5[�����-�z4#��2�I��
��E�4�!Hǂ1d�J�Y7_���SD��/�hh@^�B.f��	��I\P�g
�I�"F}��պ�!�9{2�`! ޅC-`b��xq��G?�QV(��q�F����fPe��`��u'�N��� �U6}5�aR�v�^��t��e�#ۧa��u�G�]3֢@���>>�Gk]5zc�%{A�Dݵ{f�+�K�N|b٫ @u��A�g�͑w
^- �KK�L�p�îm@�a� հ���Do��6��F�wXk��ʞN�`�0�O��Cd.�3�%���D�:L`�e�s?y�	'/.���J�e؆j��ś��l�`��.��j����w9DD�#�3<�ұ�CwJ��i�_9�1������T�$�)0�t�S�O��p�@ ��R)B
?1���#C,E{�Yx�a�4�"���ɉV5&�r��Z�ZQ��<9��H��KF�ҟ+��)�JE P.<��,��e(�'�T`b���ʘ�yr�٫I�:|��D���(���P�z�%ƶ@�P��^��
Ӧi��E��P�
X�j�Ox$H6j�%�!C���4x�A�D��e���X��L�C�1*V��� m�X���Lt�e�5�����`c��� ,�����^�<�#a�ʹ@4��[@�۩8�dE���a�la�a��V/��!D��y"�Ɛ�J�q�`��c�h�SW*��A�����"���%5]P!�P-��T�IH�E)t]�IJ�%5�O�A� oY�&���c�F�|I��ە	���K��9?F�I�L��u��ؼ"�����K�H;��49A�.�f��2b�<( =Ss�'���	��Hv*�ȅ���q���� � �y��ͨ"�F�k���xt#@O�VzԬb"�8��a�П���
��@�C q�:�0"oAbj#>QA Bz\X��YC�!���|��Ϙ)H��1FK�Lih����}����t�e�L�$כo�@!���O��y�B�^w��+�e�(_S x�s�O�����_�*+T٢bA[�Bf��O_@��E�5?����#�zM��%`'��ࢋ]�TI �p?!��R��`hb�ʄ@a�H ��
�(Q��sU "ӆB�t�T�x��C
b?.<i���3o*�P�e�Y`��](��8��� Ԝ3"
!�OF)���]��.�A0�Z4L
&T�@D��K ��1-&�m�t�6N4�2�D ?�$�Y�:�s������*�4���ۿ^��h3��<��=����O�o�x�d�ݐ� �RLĢ/v��
q�1�Mҁ�C_�� 4�O<_)��3ړ`RB���	�j�.%S�H��9���O^YZ�Bъ۸����֝[J�!ò�\�>!Jva݆��@��=
�u�%O�e�~B�\:s����B=S�I��hOp��.��)I&��0O���'6k|)�.�c�88��*�ŭ2D�\���N�2Bxl*3���Q� �b���O��1c$G'1T��2�lЯ�~���Nwf�����jdj܂"��$P��C�I�\]`T���6wv�C�,f�a�'w�����F�'��18ϟ�PK@K��!�l�R�ðUhT��w�7�O���uM��()��bF&�%gx�%�A$��W�`�ۯ�x��E�M���^���]��V4��OLQ�
'��OX�	3S)�Y�^��v�@�D���P�'�D����r�\��U�a� � �'�(|��hP�4gB�,��	��I1�'~��#�=\�@%�di���'�C�,�1|ΐl���݋f���'"�XCK��dCd$�K�X\��'hV89����Z)q�9�t�'����G^�S�!s��� |"�j�'?nl#���?=�Ț�$y�H���'� �УF�K����!DؑD{�(Q�'j��8qM�ۚ����i�̙�
�'�R�����}Hd`yL�d�d�	�'ɌU�b��s������^Ȕla�'� �[��٨t���
 %��M�*`��'�KG � `|����ٌ
g���'�
M�%�ޞ-֚M���O� j|(:�'rD�f�5����b�����'�f*6f؍TΘ:�
G5h� p��'PNl�cl��j��)�I٩?��mk�'}�� �a����MR0�XpB�'w��ȕၼ}ގ�t��;*	`���'��\Q�G!o�ԩ�th�m	�'�Z�"� �@iy&��ynR�a�'��LG��ˮ�B�,��e���� ��ԥ# j�q�aK]����"O<`A&���S~�%;�Ƒu����"OLu�c�uE�@�$��&ꈭ"O�����ܱ���)�1�t"O���`�%Dlf�:�d��M��%��"O��0��W4ڡZ�b:�I��"O��Bc�و��D���&�0e�w"O8u
V�=~,�(SG Q0�\4Ip"O��9���_Z)r��T�$�i�"Od�'jA�'�<����!8�N�"O��h�O��R*i C�\�X����7"OxS!k]8W~��c�B'z���"O(����5l8|Hg�*�z�!�"O���!�#DN���r�K�4�x��"O"\y#�Q3I��X$O٭$�<�bC"O�h��ޫ8p��C휭s�x<�u"O<k�.�1P<���įs��p��"O���¢PJ�L���·�(�( �"O�����V3/Ԅ4{g�S'����"Ov�{u�5�;�L�E�mp�"O���-�(-�\X[�-��4�@p�"O���h�;���[��L�B��� �"Odm%$,B~��I�Kԕ~�$�A���
?g��$��'��� �)�\�� �b���>��1��A�Є��	IR����5<C����Ȗ.����dE����-^$ �O���Rl�%D�<|�'g���}"���v,O�I��ܢ��4�l�)�j�5�,��!��F���@�
($�Duqn�+}y���˪�jrϔ6��	cܧ&*�auƒ�	��Y���ūVu�D{�	�)F^�����uQ (J�*��A �)�����`�
!s0�� *K�Y@̵���]��D_�Q]x�:��L>�[1ǔD�R�X����Ԩ^���X�
S �p"Q�r�
�o�<BXG�D��0R^��c'I[�b���4ŏ0:΄��<r���/�\����kp|��Z�A��5J���� ̚f���XK��#��� ���S-jvp�%�>G��5"p����(�$�D~n=�a΄7��H�!�O�|r&��<){��,7ָs'��P�q��������s�ѡ�坵.r�	��`/:�+QQ�'\x8�cw��@IS3��#��=ғO��� �9����'Q��pi��K�`x�I�N�\5�b�7*��-W������͔z"R���-�b=�8�^=�'�6*��J����^�|�����H��IY`�N�>5��h���/���IY����S��O�'�uOׅ7��S%E�V�<`ɗ��Wmducˏ9SY�!a�.C~,��`�V�`ѷ�;��'p�1�&����̴�+�	�
�ig���n�
h8A��z�d��A��[�O����i��-Z#�
'
\!��~'��0�J�0�Ċ)Y�d��MP�s�`)���4ML-;`Ѡ<H%i!�F�b�R�fHH�a�)�� ��~�(v3k��hH�iQ#:Z1���`�P�S�I���l��(��c�9]���$M�G�v�1 NҽQ>�	�p�%��gA�O�R٘T+�%w"U;G��?�A �P�w>�%��3�p=�� �z� g�]��4�Q�Z��I g�t4���H��r)���ߍ���Cv΁�Bg�	3�a�f��H�ܘxć�/~t ��[a����O��Cwʉ�RGF�0�u��ƚ����s��6j�
�䅋\Z�0q��bn7	�B�H��E-�䡊u����?���T� #H�r�
_h�$�
�g�d sW���z!6 �c߰e���Qm�3u�� �B�u8�KF	�d�j��)������xɌU�B���iA�T��� 'E	�z2�\�xI�f$���?A����#9�A��&��9O��PgEG�_��%Y�.�.W��@���"}�uAn�=J��b�H}�j0�7�����.��P�L��"|�a)��J��:�
�2qpq�,\$�(e� ��#@�^s�ֆ3��˓K��R,�[�,gg��K�(ȗ'q��:��/4a���I��6�r�gJ(d���RF^?�`dQp..Rv��:6(ڬ5e��べ�����-��9�GB�1U	���1hG�x��x��t�J�(�r<��6P�-�z��	`�dIc�m��k@+"�X����S>8P�:�ģ �i�Oҥ-�"ɣ #T�F�F8 !͒`�*I��'1D�Z�O��A�o�?�℣<]�q��v;&p:d��O�8a@�-�)#C�@�ъT�
*y��B��r38LZ�+�B@ߥ_b�o�M�~��"�M$/��i�U����?لlW�-��l��M�$^`�3?��$_a���EƎ�~;��Q�?y���u"�Xl���GcѸ{T᳇IK�P!Z�еf��{3���}���Y�bĈXc��Q��B�RF��B�z �I�'aR:H`�O8��p���e�e�p�3����&A��s��=���Zq�8���
k�\j��\��J���G1	�����
&v���p�O�AhDn�\�h�r��5�U)���C�'m 7F�,qX�E���s͸<�����M3Ư��m�T��2a�BR�k �^f��e��T�,V	R$��>r�1�' �`xu�х�ı�O��RP�� �u3K#vѪhS�4P	�Ḣ��6Hm|�:d.��n":C��,H�u��F��B�}���R�mr�>�� Y�p�>�)�B9�٤q�8�1�Y���O���P��OȔ9r��E�t(������(q�4�#cV�q���+��Ѝ҄MϘ-2Afs%� ��4PCg�����EC��R'�p ���u�^Pד6J�+@!\"Qh]�!��5j�A2b_�����-�݌I�&[�%'�勡oJ,R�~uȡ-�7o�yB�~�)� "���^�2��ebYQ��p��5)@@@�Oʆ��
�,F(o{�I�BAĆB�:��կ��h��#��L�xÏ���*�/R�}����4<O:��p�� �� HGKȞ+���׵i*��rdT�|-��T�>��x�Ł�(BR���V�<TF)�CϋY,�J�F��"I�."��a�(D��c+�D�����G�2��i)G�;���Z��/\�v�zS�ޔqvh�CkL+D����eJG�6��Iw�f��@a.�_���	amģN��*�`#�O�2��Ï����^{���'��>W�D�W�À/h����O \�ZbA�})h�����M���G|�I@�_N&<��ōx��I1w���e�E%D�ԉ�m��A��@!q�^�8�r!�)���Y�Q�aI��:����dQ ����J���д'��0�$,P�.Ѩ�ݝqr1��$;3�ܾi=�xh�-Ԉ_jVLؕ	�2��	��Ҡ��K3�3�I��j����*rL���iȡ	a\`��
�		ฉrG�.{���@f%��/y��n��/4T�bҬS=?�F$����)6�9Qw@Ȓ$�0��.b��(Y��S�R!b�4=��и���u�J0˴cR%�T�#i�(g�$bO�2N? �yA�<��Ԭ;:�����O�N�G"�yj����џp(0�߈8�鑴�w~dl���1���Se��3m�0�G�$z�[�
ɸT$,=�&�â��i�G���~B�6R�+����=��P%�1(B�ABs��:��[.�	S��s�T�NXy��e�<qe�� ;�^����ŗ��$fn�[+DmJ3I��[Oƽz1#ʪk�N܈�b�Oa����)9���V��Z*D#=��O�&T�8*bi(E����'g��lEu�$�L�*�ˎ{}di��'V�2	2��F���������fABs��O&X`�'$jht	 hͻ1ky��BE7]paz���6����ƛ� ��T��M}Ш�q�ڍyk���a
��O�:Y�T'�8>�ɠ�ƚ��쭻H�<�۴�M��ft��Pǖ�"��PQDȯ<��O�T	q�/�ybg� }xiA�J��"1Cڐ
{�y��l^�*�x�p�ϽA�ȉ0�%
��m��nK$��#�	ܦ��T�xӤ��b	Ç=�5�'�0�.6��5oL�(r�a��FD�]Wiδwj�P�ִi�0�U�I�m�4���̛mӂ|94�V���󶮓m�°�F͈/Cކ9JD(X��qa�)s��:-�wB�����I�0)��
�Gֈ-jO>��G��FՀY	�`JJ2�؉�$D4L� }��U�7����Ȟ}BRx�D,R�=X}ys�KM:���wD��M�0U��AT6�xa����`�tc0�C
X����R`"�K6��	�+�B(��.b
HixQkP�bXFX�R�ăw����fB�&a:@���JF�nڗs�B�����k��C��
P�JYqwm�L-�n��Bq���B�9RT�A��&D��R���K�$H4RV�x�ڌ���r>v�ڄ�ǣE����)	h.N�H7��l?���KdP(i�!�)`��)���"0�t������2X�ћ�J	b@2H��
�&�Y!yTN	���K��I%5knp����S��{�ឞX��p�FN�d�+u.^�����Im���Iԯ���c'��<?�h��ƌ5N�i�b��/X�i+���}�<�#��U�%(��m�2l��q��Q�}|�ڣ��(@�N_���(%�@	 �����Kp���BU���!X��V:�|1�]�s)@}1O[�Ft5�ӏ֣.y�={W����=h�Ė�lYf!�#�ؖ{�u#�ՐbaJ�����<`��!�ʀ"C�
/Cs�0��ϝ7kjt�"�ͫ4֪��Ī/�^`�,�4l��x�TM�mZ��R��{˼}_�P�ĭ��hH����埮Y���ȤI�^�̓�H��5�è�~���O�)[q�� +�[�(�걬�?Y���ҵ[��\䛅����t���)Zr�G�\(����⍾3*� �@G�,�HͲ�!��s#
0}�������ፎ��O;Z Ա�-O,@�C��	J��� ΋�W,�d(���:���� ��<嶐Ubd(L�K�hY1*��	�.L��gV�5W�A-_PR
D	�v˥E�s�І�ɨ*싅�V�[�}i�Q1���0%-H,>c�)#��s�9#QKۍRԎ��SFa���2.�e"jeӑJ�^p��#怩�q�ܖ&�đ�A�X����+f�'�~�����;+@. ٳe2��="Wϖ�J-Լ��cM�&K���|%�P�VGw2Ұi2ᐱu
0�BΗn~�0W�'�����~"�t��W��bed��*�J�/�=~�r� `MĨWC�q�˓,����.���H�*�6�8�z�O��|P��UN��9���+X^��y���"o�N��Iߘ7�ԥ��%Ȝ��-�f�T�>��x��Ɠr�f��WC��5t��3H�hYf$�.:z8��H���8��`���Fs�h��W�K2f��C8O��		 <���48V��BE��p>I����N�V���� JBωڶ�����1��qI�
�#'-䰘q͊�Kb��)3�����8b�B�Ҥ��T�I3��i��y.ꈀU �/DZE'.I2.@&����.�I!��K1�ĭ$`arj�:tC�YI�a��qT�` D!`D �P���)�����U�WD
F$���Г��'Z����?Ad�`�q��
g�Aٔ��$p�4������f�~��X��@v�l��c��Rߔ��i�	 O�PW��0<�S�h�i�;D�nu%ƒmf`�5�8m��{tkV6Rf&}���F����&q#��|ڦ �_���a���Wo@�(��0d���5&����	�)w� �1b�A@j�k3�]/�±
wO���� T�V>4%��� )��r���\J|H`D䕼VĈ�*�������$�DBP�S%l-�����?�Ɉ{�����/�+�������'�PT0�f
�w����1阽CPu��1n�9��Y+������"�PhXc��~��ߋu����!��6?i�s2Ê/W��`WJۛ�hO~�Q%������R�Էy"ґ@�����"mGl��t���F G@�#�����W�I/B��0H�~��е&��A*�ҟ�@ �םmj�� �{����P��z���R��Hl�����V�d�O�.�I�'�~�$�A��pu��Qt��`mVdC@Pd���S�D�
�Gݒ���`��F*���T�>�����%�2fߓ,��a"��q�N��)�0/j�!�k�#�`�i�Ś��-�����s�
4>y �.b ���*��ي�!�  �D����~2�R��.~d!@�픘�hO��Y��Z�0��OŤ[�}@�d���Q����E%^�Q0d$p�h���ŉ#)�@hnx�4�G�M�z��Vn�dx��⃘�RHbP���i�r#>9�l� uVrk0�I�k�,��уZ��*��9s��R�ǒ+���eJ����S��-)j�OTf� ��9Iz� ��I�z�d䱃
ǲ2��<C�%\�X�@yf�|�ܽY�PQ6��9�v �O�1!T����A��<��� �����܈
�Ä�@w�}R�oY�i�X��`�̫9@�1dG�'"��f�T�	�֐J �E�F|�YB/�ɦE���*CՄ��F��<(v�]�"YB�
4��0)%`8�Q��f��Y:�%T+@ݐ4۲�G � 6�&%UXi�����* =!5�:������[��E��&#�T� � ���X����Q+�O������2��U���ٓ<)��X��">�`Bs�֟ �#��Re�)�#n�"���N
l;@���Oj�E�Vo�Hٴ�x�ˌ3|R��;�n�>�������'~lҦņ_a�����\3Dw�d���ȕ��c��Ƶc��IFbN$c�T�q
��wcph���؛c-� ��h>��f4b��!��ρ#o�H�Q�ʮ}&z�÷#�uz>	JD�� ��I�����(ɖ��+ދZ���l��?�jacYz]d�SA�#���zTNA�O��U�3Qiݎ*�o*D� l��
�9�Q��m  �εjD��M��A�c��k؄7�>8�Լ�G(&b�	�GM�mΊ�ۣx��}��P!O� ��X�>���h��g���$��iƘ�Co	�n�buq�-�/Gx���#G�0����
֗��j��	y6f�Y���o�dy�<Q[����
��)�2�HQ��Ja"�s!�L�Ύ��(�	�F����=�d*�LX�/�(�8�ͅ�Lj0�K1�쟌���W�6�eY�F4r&�s	�<
�j�)Îٗ7�nb��9�.�3�xpK�B�"7���z��
�F�Ze���>�p(p��!K�hp$����n �$�tO
G�Vi� h�;�l(�j��<���F��D���Z�Y�t��U��~���oѢ�zt��-Eu���c��Q$��f,C�f�z4�ϼ>���` �{c
p0� ˕B�F��B��	@�'�@�H4͔.z"0M��(���WƅC�`\0�%Y/y�`X�ᬚ<vhJ0x�#Y���g釧ˢ�[�愃@�j\��Y�}�vl.�yGm��jA%��SwZ2@�2��]��̧O�l�L�Q�1��$�S�����ML�{�8(�@�
Tj�p��I1[����'L�>Y�f�5�M��ˍ�}� =HF �Pm�`�6T��S��L=u��9k4��*��DSB�o���[�$��B!ۿb������ߙm@������[�� `�:D0 #�\F1����1EM�*֬=�]�U`Ւ{ڊ[���q����Po]�HxTgCK%J����Ɲ�Qdw<�t�t��r������KrHQ��
�M�b�P7�	�;�4�ҮB��+P!�&a▴�@؟��FPݥ�$���@����xxShůGN(I�A��p���`�2�L�T�����7ON��.L$+�P������<q�ǳi�a~҃��ri0q�%�2'��C� �d���LX�|YH s"i@>#^�Cπe��E�#��k��ĉe��	��l�^�	S0�!�.gQV���N<�-��A� i$�⵬
�[ڍ�'l� �1�	�
�Bl��	І;���f	Pq���`iE�O�A���@���dG�(*�B0g[�/�(x�a�$���ւ;��8!E�	U,��"��"���h�A%tk��)�XPƀ��q���G���"-�����	�L\J��:$Tb$�0H�/�л���e?�2C�C��iq5�^t.:�!��/;�](�o�V��]G��u���T�X�R!��Iط�����=�&9����VS�I��KZ�~sv���(I�[��[e�68����g�+M�����k;WQ��>�2_%B�Z�J�*�t��m�<Y�?�+و*2�����#��P�h[ީ����d8(x�F�[A��޴��I ,��
��T��(�?�=9��V��F����%:餅��c�U;Jv�M�{�O��ꁊ��P����Ǌ�n'��@��#����$�m	�3��7�p?��H*�! �U/	T@��I[��Ōʪ#�D�s Ъ\��v���ڔnHش��E 0z�07"O�1c�Z�u�t����+ZD��;��'���x� ��]~V��u��{?E��Ur[8-{�gϨ}`����U�Zz!�d�}���rI ��O�-mT˓'E�5)d��>�����Oz����� )�@�ꆶ_������'��=񵢞7y[�}��Ԃr�|�2�a���^9���G<��L�o�`$4(ب)�$�
���a�'s�Œ�@�`�'3p�lp��N-+�
�~�=��aVtCBތFg*�rq��_*(5�ȓ��!���AU� 5I��(�t�ȓ50�]�w!�D��c�J�IU��ȓ-l�q�RӵcpF���+���
��ȓo ��k�m��ȷ�+�VU�ȓF�L��A#�5z��)x���s��,�ʓyp,J0�����{W�;	)�B�I�Ba"�ش��3rYw�ݒ)�B��R��=���R�[Un��V�\��$G{��U���v��É�y�!�d�u�Iq�W72��%�c���!��Ǥ#PĶ��I_uV�H���?�!�A�JP*A�Yw�)ࡈF!�!�)n����u�@�Hb�� �J�w�!��G�r�E��8P�.�3�Z�z�!�dǞu�>�C���np����	�!�䇆I9ve[�ԅ#�ʜ��nõ�!�DV�dc0:�"@ _���c����\r!�Ău����g��?ᜑ!@�R�:!�� �!���ջo�(���'�<5���;�"O��K5f؟h�^%	�fƑm��!�"OX�!�A�{qX�ct�["T�fu+0"O$���ہ0���0�N֚��"O.�u��0��d��p���"O�X�#�G:m5��P�hJ�s*F�b�N�;}`����	�%���3�B���~�䁿i��0��4(��r���$J6�?��E8:7���� z�$]��.QaT볣OF�O���G�M��k�JY#$���d CgS���Hfvt��!lӠOQ>�KV"ȚeEP�#E�j4]Z"�,�d���(O��B�r�
�*�9�ք�S��ij�W��P�韞McҞ|�&c^�"���)U�z�ť^*�M�C��Z%��l�S�=T_�u����z�' ,��QґA� [i.��I/���A��Xh�'Va���CoY�v�f*��:��j���y�O�!r��m>1��c��j��t:t��h� ��Hӟ���I'CF�I�`��$>	2 �9wS8�JVʟM&@�0�ĂQ��{'�C/�?�t"�3{B(�����]2�+Z�&�pĊD�@?�5�a���c�ܴ��J�G�J�c?�l��&  �bt��(	�A!��q�&?�@�`�@��%�"�`� х�9�؍������0���OR�1�N�<V託���}bVAKMѺq�'��]�$yt,	�f����[�|�؝'Ɛd��&X>1d�ةcx������8ibZ�U�@7��2��N�O�M��� uxR���	(_��9��O�_�f=-�J�t�I�_��1��_�d9	��A���i��K2n�F����H�X����v�K~��~b�+�z01��y���a��
:ʼ�Q�S����'u�}%��|R�, +�B��T��*y�P�m���:�'�T�#��֝5#>�1֌ �{�VyY���#p�Έ�w�C�c�
6͘�/���0|B��Ѣe��xP�����q�e�Ħ9R��W~"��=a��ΑA#�l1�b����j|���'�,Z�iq���)�%A$		���@��T��1��d /�J��4I1�; �S<D~� q���9��ܐ$ �<e���H�t�<� ��'2���lѱ#28R /NY�<9&�=Nne�FFF1?�9����S�<��섶���R�n*6��C���W�<	u���n��d&�*/���v�]j�<AT�[�,�z�)1�, ����Ac�<a�N?9�<xb�\.+�i���D�<QЇ�2Z�qb�B�( mjL۴)�i�<1�U�y�NԘ�Eݠvx��7�Aj�<����&f8���c��q��u�h�<���1���.X.{g��Sa[H�<���L� ���@^fњG�@�<��K����6n�Ⴊ��9�!���D�~HP ��m�9�f�Q�!�ضB:Z�hr��ag�1!s�O�v�!��Կ.� �0&��\��3ƣ��OO!��w�� �kE >n��A�ݻ\!�Ę�i��ڔA_�p#Ե�� �	r0!�֛zݘ�R�LB�Q��B��ќR�!���^0��Q[�}���ʁ/*�!�D�Ukl2F��	� ���ϓ)!�DH"OH��H�냀�	cT6!�X�0q���L�-|p�q�b�"D!�͘D�~!AeɊXe��;�!�S�!��	t|2谐�G:j���hv.��'�!�߸.�t0s��;~���(sM�<'�!�͔DФu� B5��xIe,�7P!�W�%�X�`�J�Z��1 CL_7`!�d��X�e�-���k��0K!��)J�>H�a��^$�*�i_�A�!�d���!s5o�h�S����!��6!��z�e�saZ��ǧ?H�!�d�/�,="���C\xS7�Իo�!�DEq��X�&�Q'jL��` �l�!��� S�6x�)bHVH��P��!�� �@
!e �(��ㆵi3���v"O�|{ׁ]  ��!Yp@@9,�s"O�Ѓ6�a�L!�/��_��]�7"O�Y:��7^�&�iP.F'v� HJ�"O�[�C�<:|ِP͎�&�R��"O����P�Ph*7DW�Y��Ir�1D�xq����__:u
`�SI��k�-D���f�*H�VI��S�=�EKj+D� zb$X�m���(����Dt\=I�-+D����݊k4� ��Vx�`m#G�6D�
wc�E��"�eՋv��DB��5D�8� ��gs�3C�*U=P���)D����j�"?�`� p	3+�*�"Vj'D�dA�&ݩ><P[ .U��!�U+%D����E�tG6xR�z���dn0D���1%O"*]�؛���3�)���1D���E � :�(un��d�$��g@.D�Tz� �0R�2��U��LA�+)D�,�q�S��+\�ZL$�hC��X�<�w�P�`��@�c	���k�Z�<��&F ;�`��N~�<=�Qe�K�<���&88
�������#n�R�<qG��4"�"S���Nd���c�<�6K��4)�D�����=�L���Rd�<1$B�&耉��Ԫg.`,B�N�^�<���.�9bKmX�=S!�A�<1�b >J<��"�_p��rD˗}�<1���>P�t倥���8����q�<�͘�D\mHA-	\ptrW�@g�<) ���M��d	��G��` Aa�<�_�(�|���P���\1�%Rt�<�$�_!Q0#�D	�&NzD�	e�<q�^�Pn4�
���^�a��b�<)��ߠ)2��C
��v�8T��G�<1��Ƭ
������1(�^8�r�FF�<�r��/4��T@�.'
.v!����~�<�����i�S�s���aa�|�<y���!l����Lb5�`BLa�<	b��:�h��/
9?��)�d�XR�<��@� |�b$�,�E��d����P�<�qC��9�^��̒)"'���RE�<� X&��i� �j+� HD�^V�<aEE[	�a`��{ضQ�G�WT�<��d�4>�4@�jE7Ҷ�g�
F�<	b��`���t������b(h�<iW�E��D�"�"ӊ�� �d�<�G��l�d�i�N͈M�0Eg�^�<A�d��lZ�D� ��xA��,^�<i5iߎ]������6k"H��D~�<a��
*yN���2]�0%��N�O�<A�K{�\ԉ�͝$��YꑈAw�<�4O�)Lt�ɺu�,y�x���J�t�<��� KMٿX�J��FFk�<��K��4���!ֻ�60���Je�<��V����P��X�|T�'�_�<�G��4���x \� �SU�<��ǂr;�阣���=�]y�%�R�<�����9�1��+N[����bO�<I�A9S������R��`���f�<�R�N, {=3�f���unk�<�tFѦ8�ĳa��F�����~�<�W�n/�̰���/�ll	#�\Q�<Y��"m���f#I_G
|�e�T�<i#��&f��s/��(�0u3�`EO�<� \���⟉d�
�J���P�0I�"O�5���rO2=0U
ݓk���h"Oq���L[����?#��!�&*O ��E#�+���i#B��H���'HC����p	 �ꓳ�v�h�'U��ZW�A`�.Y�b�R�yH���'���b!��,JڑI�d��H�T��'� xcd.� $�Vuh��3t� �'��Q��έ7����*x ]�'W�h� ��� \7A�8>FH
�'�b��CD[줵����fUB
�'ҒXx㣘�;r3 i�3{���'�9��A�5�h�2柵q���h�'t�s��O&G�zm����#S����'o�������)��Pv�M�T8��'+b!�)KC��ҵL�I���'�@�cB�� [�J�zh�Fs�P��'xT�����	��RtIK�0A䘇�n�&<F��:skh��tO�,*[~��#IX�!"�y���fR�5a�ȓI��#�|��q�T��� \V`�ȓ8C<d��R?+ L��Ţf�$]���~y�vd@8�ȁ�	� G�:��ȓG54�uD	0�t03�x���ȓ�Ȑ;͔v>�lPF��9d���X���	�D��_n^�+�bN1
� ����t@�4��FLb��P��8M�bчȓx�� K��΍U ����/�1<��%�ȓ9zL(r��tztm�nB� �̈́ȓvG�E�r!�]f
�3f���"�n���q>�J��Z�p��5[�Ҫ,v"�ȓD�ң :e5<��wj'Q�`���P�"0�
֗:�.h�.̉,�a�ȓ�����N��T�t�  Cڅ ]��ȓ5'�"��?��jd�ê�p��ȓlU�C��_�@p���3��.h��e ��`6.��Q!�;�iÍn: �ȓ\㔼�	y��,q�5&�Z���5�uZA��?����f�0cr����qQrpYW	�*3ڼ�8��˫[��ȓ�^�h�]�z�d����&'_����,_L8�V�
v��I����W����>|T� �����h�O����̆ȓ|�F�{e(F�Y���9���A�\��ȓ.L�=�wJ^�ZБtLR�G�z��Ί4�l��6�w��?4�����fL���j�!\�堊�y	�e�ȓ[/��`�#wBФ8VKˎ*n�0��bޚ\P��;{���;�hǠ��b��=
  �	�0L��C0�%�ȓU�yAo���[w�Y>hʈ�ȓx��!��_v�1�'�"9T��CE�u1� J��P�umK�;�hІ� ���Vd��Ɣ*�jׁm�v`�ȓe�e��H̶R��]�O�T�ȓ��0"&�^�bo�}���R�-�l��%o�YA��{���[f�\�>�ƕ��|��܁_���H��-�0\䝆�&�:���E��=
�kC�
�A�%�ȓ:�������	���Q�􆘄ȓ4�%� FS�r ��_b@�\��-$�4�s`T�Z�b ����`���}�FI��#��r��9�UN�2����{�4���¾!`|x�&�2-��S�? ��bWk�8ע������UqA"OV��瞪;vDYrfˋj�lrc"O�� ���7d���T�)`��"OJ,꓇_�n	T�cGő5EE�Ĩ�"OV]ReW�?޶��RD*>A�@��"O��9����Ë�U�n�� "OF���OUs�d"ƢŤ-�j<{�"Of�㑅]98�����!D� X"O�eҁd�"E�8ɂd�@�Xx@"O�]"E߬c�$�Q䁍���"O�T�B�|��c��;�b�+�"OF�#��J�D������H-D���1"O���J�T!(�cƩ�	P��� "O�%ڑ�דg�y#�?^e� y!"O��S����d��� �NG����"O�qB7����@y�1,F?FP�`"O�QK��#;r����k�4�0h"O�aV�ŭz=fk1��<��W"O^8A���*)sV��s M�+�@�"OHZN��D�&�������6"Ot(V�O�]a�йE��2��@K�"Op��F�+d���� dY�'�����"O&�KC�X�X���ŅnoX�S"O���T���@X*��2���{�'c�Ȫ#�Cp��DꋴCb
���'b��!B�.C'�� �l�GTr,��'^�)�-ėyU�i��\�Ff�c�'Nu�$t3���F=�-��'��2�hB�ct�CP
:9�,`�'��4 �-FT������ni�'������p�	3�����q�'��%Iq�V뼔)�j�O�(�'�T	���>��1A\9�fX:�(2D���0�E�BDݡ�Ғ�b|q&D��p�B׿��9��N��U3Q�"D�S��   ��   O    r  n  +  a6  \A  �J  �S  Q\  h  Kr  �x    k�  ��  �  5�  w�  ��  ��  I�  ��  н  3�  v�  ��  ��  ��  T�  ��  ��  ��   �	 b _ Z  �& �, `.  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,͓�hO?�zP'���|��6E%V�ၖN'D��At��j��KC !sx��rh8D�@+�-�65b��@��B��`8D��S�;���!%�*��u���6򓑨�E�3#νw;@R$��Kv��U�'މ'<�m��.[&�9�BM�3�ڴ��'@�X1/�U��yk�H�+Y�8仈��?�S�T�ݚ���t��e/��� �(O��d��%۰��w��
K����d�ҢB�䛿�X⟢}�wi٪M,�Ad`�,M�<Xq��N�<I-�� �J��	f[p�Ё.D/����#�HOP��x0��0*��`�2准N��A�!8�O��hG��:�޽`�y�fC�<f���?��� �S��H�eB��B�2Q��!̟C��0E���3W\��"j^.ܤ�r�S���ĉ�t�f\:%m�8/���J�#��xb�Ob�>7M1?�cɓ�%��H��k�a���ç �\�<�2��*�L��(� �&�cg(^�<q��(4`�l\���`�e�Rx��Gx��
	N�`
a��j� ��5ㆳ��'^(�EyJ?�ІI͂X*q{ C�5,2@���'D�p���;a�h��A�&3d�ͩ3G2D����iZ27R�1��e�'����.D��(W�Ϩ��A!���(A4�IqE���`��	b}��K�kD��i��̠:�D���eգ�p=ٴ��C�:a�T�\*͂��D�CB����	�'��rF�U���j@	�[$�� �{��']�O�Oe�A��M�G�&��ӳ����'�ў�}� �0�FF'����k��W�L!��O~c�h�㉄�\���@��}2u#����k���'�a}Re�"~"��@K�J��A�W$bU����ɾ���m::MbGh �Szn�c�S�azR�D[�ux�%DYT zQBgeQ;aY!�d�>@��xt�[<0�a�I�u�����'����`F�;֢	*��E�ՂA,D���O\6���n��e��,rgJ?D��!#C��f\ک0��0JR�l��2$��SF�]"'�ZE��Y��)3cݨ�yↈ%O�BIzv�[J����ع�y�[�V�P1K�*B�%��5�&OO��y2m��p������]6 ����Eo��'+ўb>ّ0���%.E��)69MR��I6D����#�
T�^Mj��H��&���2D�p��(k�d�ree	�� 0� 3D�܈SB�#5s�#��G1sư�ٗ�2D�x,���Xf�p|�����I>����+�Yվ� 	��b�� oI*��B��+w��9�P.(�4��&p��b� E{J|:���J�i��!��/�r��W�<��]�V�L*SLU�.^-�T�S�<��E�E�̝
�B�/YY��()M�<�Ơ#q'~Pv˨V��H��
OH<���֑.�*ԀR�\U#&��S��%��{R��Y2�[g�R:�}j��	�>a{b�'(��R�k��'w[(�kÎ;) 2`���\1�cg] _�	@���3J/��G}�ŕj�O�� ���Y��A,^o�`k��d?O�4��O ,�ظO�"Z��h�u^��F{Zw5�O̔��"R�.((Ԩݭ4�93�"O�y�+�_���Z��ع"�!4T������9��xFz���7�����m� T����?��D֏&˖�G	ؐЮM�TNON�<qwo�;8T���l�O��ts��G�<a�y$��!U��#L��רM��y"�ށ)�J��K���W�Q��yBF��v��TIU)�1I_ ��!�3�?I	�'p����I�;��1�H^�d�L�+ÓJ���35�4#�SJ J(y�'O6D�8S�&O��d�$R� 	];��3?��)§8�����֫=eH��� Qf��|��&0&	#c�!j|�`��M��VV���hO�>�� &��A�D(%�"�i$"D��$�I�^�F����5�`<hu <D� �1���;�(��
Æjv���q�:D��	�j��o �H�� ��'`:4��l-D���@�7َ��4�ʒ��x�Nl�p��ɋ3����N�(W{� ��K"X���Dv�"o �A�D�[��F2F���[+yh<�c,A0 =���"���.��d�D�<Y�a%�!�ËYzպtZ7�Bx�<1��I<i�i�7@�����qx�|�'�\̀dW�E�����(�¸��'���C�]7`�r@�$�s��̓�'N�H�j�0
�fd)�kxTh��'u�s@M�4q�z���=n���'"LQh��/@�$�*ci	N y��'���)W��L�jS����W����D#�O,$��k�61��!����5@D0qr�'��D�E!�?`����%Ќ7.j�&#*D��Kr�&t��m�6!س�Z ���-D��F釋r-�XY����t�9t�%D�8R]jD�6h�@N� �	�$�0��)� 2����A ��)$)2+ �H�"O\3�ɕ�v��eqVH���;�"O���*I�N�,pڐHX�~� d�@"O���h@� w8��&�'���s�"O
	X�o�9�H����ڤ��'��Dy��)_�a�R��R��/&��a� ,,OТ<yu��2t�pie�J2+9�D�"�	X�<�O|(�G�T�]�<����LSGv�r��d`�<�>ͧO.�	�\qh-�G��~�@�a�6�j���'Ԝ��N6p���'�Ÿ}���{�\�4G{�'Y>\�ǫ�;�>p���6�@݇�#n�t��O;�A�$ь�6��=9�4�O�O��iQw�ό2���t.��4�I�'�����5Z�F�RD��4>!�PY��-O�9 !��i���)c�74a×"O�E��dƄ`��4¦�=r�ڴ*�"O�}p�ю#R�0E��i�J���"O�$��^�p��!�Ժq"H���"O�h��ЩNZ���a�/�֭�R"O�41W��)A���� �?b���z�"Ov8)��V(<M����F�!x��P��>	�$��	�׸>%|���R��p)��	Xy"m�.��ܚ��afN�z�$��y�Ǘ`
��ۂ��UK��˄K[��yr�	.��v�F�S�
YiA�2D�dC�������6��d�(�a�$D�DS���3?^lm�E-]TƐ,C@$D�,��/IVy��Kچ��3��"D���f�P+o���eM��o��<�%;D�l��[�+��A �S>��S�+#D��h׬'�J܀pi,IE����5D��0�F��A	�ϰ���7�2D�@a$̒�(Q��`�*��f����h,D�hg#�ʞ��G��N��k��*D��4Lܢ@̢-25��Eeʸ�s�&D��7-�9]䠸q'CX& �0�DA%D��૆#a�RD	���>]�V@y!"D�`����<x�ajw�W�8-�p�m>D��1��N�x��v�փ;7ꔱ(;D�d:��ڮCU�AB㇖g��<�Ҡ9D�(�UJ�1 Hp���3��#� 9D�l��'ȤP�~�!a�S�q!����9D���ϰW��()V�����r�8D��q�ŀ8���bm�	�*��c�*D�y֪��@�Y�a�I!5�2Qivf'D��P�c�|���Z&R�N�/%D���Ʀ
�@:����@�1Mbd%yF*Op���݁�8 ��]���0��"O�I��ī.�>-ȗ!��6�$YK�"O�� �O�,G ��U�]���K�"OFaa˚+"�
V�[zte��*O$�ʢ���Z���L��I�A�'vtH�AU0U��Th�� 5,cl���'�-�t�%o�~�@Q.�l���'�J��h!1N�Y���!N��S�'R�kW�̣n��(Z��O#}eJEp�'M<ƕ�B��ƛ�E���'� %u�%}"i`�Z<�"t�	�'΀� QHU8�U�4�8�	�'��TBЋA$D�
QJ$E� (�����'l=
��?N��\
$g�'�nԓ�'���Q��X-�:�`@-\��R�'n��� �1Q:���C�-n$59�'#�-C$J0_�d��2�_��d
��� �Xʆ�D�L�"-�D�q��,��? \�
�'I-0$!!ATvńȓOHX��F���n��X����Fώ��"@@���	��`K�=Ilv���c�nY��� v>�X&�Q�@����ןt�I�0�I�h�Iϟ��	ԟ���{��` ��
4xJi!VK�s����ǟ��	֟����� �	ǟ��I��	��>�s��� f�8ԀP����I�����۟�����������ӟ�	5Yg<�k�FE��r ����+�d �I쟰���<��۟��	ӟ��ߟ�	�6�!��;((�2������<�IʟD�	�������������Iǟ��Ɂ&Ⱦ|��X6{=���B��<~����ҟ��I�	��������I�����:V<���A�tV�2�J�1�F���П��	�����џl�Iʟ ��şX���	�F 3B
�1t�8�Q�|�%�	�X������	����I蟬������ɱ,:�SD��U?(yr�,_!������X�	�4��ӟ���������d���i����#AqB^��^�f�����$�	Ɵ��	�����ПT�	ݟ��	;0ӈ�8g�[ht̤��$�*鸩����������I����ܟ|�	ҟ��	+�TԚ��+�`�Aq��|�����$�Iٟ$���������������	�����*�#H����4��iʑ�����IßL������I̟$��4�?)��<$d,K�@�-�t�(�E�T��i�UR�L�	Wy���O$�m,keH���A�(R�B��7���|��f�$?I�i9�O�9O��d�0K�~����>6\�P�L�=9��D�O���wGt�����ԡ�(�O[l��F���9��r�*�=6��y�y��'�IA�O�(' |�d���_�.���1Phh���8�D6�S��M�;J��LY����"�h�ئ&>I\^أ���?��'h�)�S�pR}l��<��b��RJ̩���#c���5
Q�<I�'<�D�/�hO��O���Fhŗ�8��G�k���(U5OTʓ���FD���'Č�a�5�@���H̘J~*hjR��NJ}��'��9OV�Ũ
T,�}��ͨ`�.��<�'�bR�>��1��d+ן�1g�'$$~�ؤ�3�Ig.��2k��i%�ly"�����dT"�V��p�����F�5H��Sʦ��Q�7?Q�i��O�	�� ���'/�h����+��D�O��O��I7�m�*������ �k�mV*�.	x�@�0��`j5����4���D�O^���O�$N;'�A �R%ԕ;�\<�L�Sg�&�R��B�'�r���'�n}��(\V�%����)��yj�o�>�ݦi��d�)�Ӟ=����Q p j��!��U�|�<�"���S�O�y�N>�+ODP
pj�D褥�2fA'h�.Hz��'=�7���L��k}� U�A�e躁�!+΢����XϦ�?iP�t�I�����J���֩ߟJN5�ȕ%N�rplA~�4WX��ӭ69�O� G;&ȴyV�O�DT���,˓�y��'���'�r�'���Ƀ7|��P*�bt�	`��1"q4���O�Ҧ]a.�i��'|�yB�߆�x �rC��1|Zp:�|r�'��O��a�������<<���
Y�U�ѪG9IPT������V�&��\�������O
���O|�Ĉ,{ �����r���2K�-f�.5G��O�����=��'	�O}W�����i�D�0kӀ��j�y��'b
듥?)��O�2'3�z)�`��AnݔBA����L�:��=x�U� �Ӥ2t��D�	 |x^��f�SI� <�4&V#q�\�I���I���)r��?��Ė���@��"2%ɗ�]�Y��8Rk�/�<�'[(7m�O|��?�0[�����y,����*���`��a�t�Iԟ�
q�Tڦ���?!-V~�i��$S�t�.�`⌢a��r�#W�Ģ<����?A���?���?Y.�:H6i�"٨I�&O�kL��n֦MH������	��D$?�I��Mϻf)���&T:l-��:p���j��?AI>�|�uG�8u��Qϓ-X�xW�''ux�l��o֤��w�pB��O��N>	*O�S.pTEҕ[,(�1�r��[�F�����E������	���� ��e��'�qڂ|�v�C����ş���R�	�n�B,[�GM2|�T��snB~`��e����Z�ԈL~��I�O��R�|ٰ�P��>u��p�(R����?���?����h���ĞR���%�{~X��#d#Q6���ݦ%y���ky�OlӺ���E��]��,˷�����l��t�f��ş|�Iݟ<��f��E�*�:��Mj����L���_�R6��TE�v�<ة���
������D*�MK@kL��jB�ʍS���M��D@�?q���?���D.O�r��8�V�ǵ�k��9t���?i���S�'_����K�?P_�����8��0�M��^�옴��W{�$4��<�𠝠B0�XC��D	q���u�S7�?����?I��?�'���_�QZ���ş�*���&9�r(�f
]A���bhW�|r�4��'����?��Ӽ3��.�Bb`��>P��m���0E+|t�b.{~b���a����ӪBD�O�� : ��]�8A�N�oX&%��:O.�D�OF�d�O����O�?e�+0��H[�zCfMZ�C��X�����ݴY�l�,O��o�n�c8���!��,���s��H6�$���	����K���jP�&?�a�D�j� C*��Tn�����E'Y���1�/�O�YCM>9,O���O��$�O�� Ƅ�LU�!9%� �j5�7G�OD�ķ<t�i�hj�'���'�哚(ϫ��*P���R�:xbE*�O&��'��'rɧ��,0�tt�@�	���Q#�&ѯ?q���2	�)kn�Z��	S��~�� 87��
� �zZ.�(V�L!�v��	����	ןx�)��CyRCgӊː�B��P��*\1q�*��q�ѭ#�(�r�����]q}��'�l��߀k�č��\�{�j��a�O@�D�y?�1������0nW;1��ԟ~��� ��1�A� �l�Q����<))O��OZ��O����O>�'�Ƅ8QOѡ6B p�tiI�.��` �i�Q3�V�D�	L�S�P9���;#��7&�H����w	��jތ�?a���S�'��M��j��<Y�'m���E'X
d�Ѧ���<نa�>X,�מ����4�B�DN�|�&xr��Z�3�������I��$�OZ���O0ʓԛ�/ȔU���'D��]�\D^Aq׮ �N�ks%=r�'�R*�>!���?9L>)7}����D�7��`pA���<���4J��S�
�j-O���ø�?y��O%0��
5��k�n�ia�\:�"Od���ծF7�,˄�_,}F� ����O4�oZ6�r��	ܟ�2�4���yGd�C` LY��؃W��iF����y�'H��'[&���i��ɂ" ��a�ޟ,! �= �Z&J�S�J�a5
)�d�<I��?!��?���?I���Z�h�Y��_�=�t���9���-"D�X��t�I�(%?�I�UÔ�H��اIy��u�Ԕx��1��O����O��O1�t��� �$$��{�#��j�j�!i����9Ҕ�ЪQA��a-���s�	Syr�
?O�^,�΁7Ƕ�����0>��i�z}�$�'DTcWB�	&Ď��el��7b����' �6�8�I
����O��D�O�t�v����y����d2:A
��5b3H7�<?�)�8����s���-`�^�Ҕ:�d2 9jՓ�s���	�|�	��p�Iџ�&?���n���B�ys��$=�p��oI��)�<^���O!m��"��'��6��OZʓ	5�UJ�*� B6�Xe.�d���<Y��?��X.2q0�4�y��'j�4��[����ѢI�k{���^�x8�I*d�'��IY��.�EzRfE�W������hlHGxr.h�b�i�O0�d�O��'l���P�g�
�����Jm����'���?����S��_�yv�Ö��
p��aA�e݆S������֔Bq*�H$[�據[T�"�~��)(��\��J��pI�P�L-!����<��ɟd�)��]yIc��U0�-��!4i{PF�.�p�R�Lؤʓb���ćW}��'���Kߖ�xQ�"ˤ]�"^����	�5+́�2I:?���͋t��)3�4c�Id �Mtu�ȱE�:�y"P����ԟ���̟ ��џȔO���юB�^��a��DX"4`�D�pӪ�«�O����Op����d�ɦ�]�N����G&;����!����H��?�L>�|�6 �; `͓Oظ%��}��Y�Od�H�C��y�	n�`Q[CI�(N�T��NU�\_f%�E��?(�$i�O�U���taX���O��Wy�=��䑆z$�Wלe����g#�:�M鵄ZX6��Dy"��
,�
 �`�1M�� �ţD����˵~�<����W��R��G	�K7MP/ V���Дo����*z��#�Ȼ.�:�T�Z9Q|d��n*d�hlJ1)ܢ�@E���4F�>��6
š��}Z׍Q/}$��˷�ǥ	�x�RE)�]� -Q�r�R:@b�d� A���6��q�Ĩ��<<\9�!-v����OU�tBA&n���Ȣ1�Ĳm�Φ-�	|y��'���'WB�ZsT>�cu�UРZ����k]��7�Ҧu�	��'f��#��~����?q�'e���S�I]�B�
���֛H��ʄ�xR�'2"ˎ�E��O4�&,/δ���I�i��|�b�*Ɣ7ͥ<agL�'kP�&�'*��'D��a�>�1x~��1�	a|y�ք�6EO��n����I�(�:X�?����ɏ3x�#�-�>%�P&��+�M;��F�����'-��'�����>A)O��%藊zr�x��M]ql�A%����	�u�ߟ&�������7�(��B]��4k���Y���'U��'E���G�>�*O������D�q����q�wl���	|��Oi���x�������蟔)���;q���F�6%�hS%(��M{��W�Z���V�Ĕ'.��|ZcU��#T��K�X��a	7D҅H�O`|�$�O��$�O�˓`	�q��I�3A.l�"��h~���[7N_��Ny��'��'���'*����͞�Jzv��'�ߛBhQ�T��9�BQ���I��IEy#G
Kv�-aT���(�_����f@:~l7��<������?���,H��'���3'OǕ}���C�}�d@ȯO���O��$�<�c��V��Sş�3�!�A�`x���&^���`ߛ�Ms�����?y�||F�"����	_T����!Vt$��߽|�"7��O���<��!�/^��ԟ����?�A�	�&��QݱJ�K.�%���ݟ��ẘ���d��^�j�!�
�p��Ӆ��MK-O��Z�KHߦ�������T�姀 $Ii`�ƇwW��c$�	#pI6��A�i��'���'���$�|n�:�=�U�H�!,�i���:Q�B6m�	-�m@����L����|���ŗ]��b`J���L�@	ǝ���'}��'�R�L��y��'U� �T�؀sF��۳�"L �	�n�X���O����
 ��%��S՟��Ic�(���_�`���cWI��!�&3�4�?A����Y��V>Q��M�C*U"S�&Ip��Y+]*Dڰ�M���ɠ8^=�'w�'��'�AH�Ç�ʈ�hM�:!1��%I�1Ox�$�<��7]�HIV
Y�[�vqr(U�}��K�����O��=�	�����j�>l�A�	@��IցQ��ȹm8R����?!���?�*O(��R�A�|�'Ɨ&4�|�[2��8+�补�Z}��'m2�',�	�ORI�|��9����R���˴�ڠ.-���?����?a)O촲A�KU���vb�J@U�Q�\`��V-c�	ڴ�?�J>*O���O0�O��[��4LN���ɐ�_�2��4�?�����$,��&>��I�?ט��^�i3��p���阯 �@6M�<���?q���?�L~��CU`+[����J�1[+ԝ�æ��'�ڌS��tӨ1�O���O�N�S�0�I���*b���y�Fؼ �@nZƟ��	�����ɭ<.�����F�����냱*�^����8�M{𮛟�?���?q����(O��F0F!#֦�%� �#b���4���#�O�����)�'sĄ��T��_c6؁���!a,P�f�i�R�'<"E@�*��)�H�(	գ�B|:��e�� 1�ZIF-�O�4'>�������	�j�`�BA�"[6� �C"��,�ܴ�?�Vˁ&a���4�'��S��BA�����9+D-�4ߦ�M)O���<	���?�����dǬ�N��U�8c��ixU`G�"t�҃��|�IΟ�	S�	NyZwA(8"j�&E�1p�\��Ԃڴ�?�M>I������OzAW��?}��Cְ �:�B��n�(��j�H��O����	qy����M��N�� Șb�9 ^���ZL}��'B�'��	� .�:����d��T��N�a&�t�� Gw���l�؟d�'8��'cr)��y��>�v��&Bʰ�g��#9�4�S�����	����'%�}2D-�~
���?��'��x���rB<\0�K�&Aᰠ)�Z����ɟ�	�L�X�	����'����4+>�quB�FVd�������vU�(�o��M����?y��r�[��7e��E��	R�R �pd��B'�6�O2��A�{��DT��'�q��|��#�I��0s!�΍E��TI�icD!1�ct����O��d퟊��'�剂�HC�*��dxd��Ei�>�b$�ܴ5��̓��$�O��?��� e�����ެ-(� ��ċ�"�(#ܴ�?����?Q��M���ly��'!�Ā�4>QSC
ʌWvy*��B�����'k�	�Z}��)���?q�OJb�X�r�Ǟ���{B �9{u���'�����>�/O��$�<����5	�2�4�p�ǘ�uE�R#Z��50�	ݟ�Iܟ���Z��'��hK�1}�N�X�H�����0��%d����D�O��?����?�E��-�\p�P/��;c�@Ã�٧%9����?����?���?�(O�m�i��|����tBH�dK"����ԎZǦՕ':T�������I"0��牝���Cb�0�-���J�`z�� ش�?���?����Dڝ>�F��O>"I#�$;P.�.A猬Hv���4]�7-�O���?���?IG���<�/OB= ��� ~����!���R���������'�R��t�~���?�������dT�6P�\s�]��<8�Z���I؟���%wQ���'?�DP�r�@<f����� Z)t�L�n�Hy�ċ�L7��OV���O2��Pi}Zw��I(,��j��U�Ks(`s�4�?��Ԩ�ϓ�?!(OF�>iQ���v�ht���8(�X!�&g��x��ͦI�I������?ᣩO��!p�*� �7���cW�w�2��im8���'c�^��b� 
�{��0~�r!� �s�h��p�i�B�'�rX>�H�����O��	�-�t�U
+#&�slӱG�D6��O˓W����S�d�'�b�'��k��*_ ^ �6J�`�0uGb���ٶD$�,�I(%���&�����P+JD񭏧0+*�M�ĸ�<���?9����V�H�b�+߈CQr�f*H&S��ࠏ�j��?i.Op��O��df$|�C� 	Sg�H��k_�;�օP�b�O��?���?)(O���co��|�a��}8��]>�n��c*�B}��'�b�|��'�B�_�~�dH�Y}6T)A#�?s �6)˷(��ꓘ?a��?A-O80ɷ`A�S�a<�7�6c8���9�-�ߴ�?�K>Q��?�"+�<	J��R�[*nCX\���֩=�N�BB�oӊ�D�O�ʓ|j�q�Н���'��T�[�O.�!3F��p�P�V%��2b�xb�'�"�O��>=����e�"Ll��5;�6M�<	3���6ʪ~����g��P��Z�,H��B�*���bW�mӢ���O�$o�D"�D%�S���5�u�ЦZ�D�3̛ R�6M��%�Bn�����՟(�S��ē�?Y�N�6w4<�i��i��sƬW;)��V�_��yB�|����O������	p-�@��JԾj~z!��馩��ן��I�89:�}��'��� ��%���X�29X5	��%��ٛ�i��'Q,��$�/��O��D�Oh�xW���K$%B�ZF`]&*�ڦ�	Iئ�3M<1���?�O>��2�d�Я*gMMBdJ��O�D��'��%s��'���������'�l�9���69&��Vnc|�̙ԁ@
d�O����O�O����OX���_����&TP@�Qo܀��d�<��?�����@
4� �'n�����A2�X����}2�$����e�I럈�'w}��ɣ?���&��/Ԇ�҂oǱ;M�ۨO0���O���<����+Y�O��y��A� 7F���GB�[����}����*�$�O������J��<}P$>� @M�6wU��0� ϟ�Mk���?�.O��,�$>��	�?�%�*O��*�],�i;2���ē�?���c��[������EG�J���L,�q���\�Mc*O�,�O�Ϧ�Ю�V�d�4��'Wj ��Q���P�� ;r��4�?���>��i������O��\�#�L!q�^T����kc
"�4T���y�i���'��O��c�D��Z t>̈2һP�xP6!��MK����?QO>���'4�IJqIQ7!��bԊ��ujΔp�d�l���OX�DF�4��>���~�b�n?��y��\@l,�چό�M�K>�T�Җ5�O\��'t��Y#�Ӌ�,)�Όp���K�$6M�OJ�q7�
Y�i>�Gy��rM����Q������?Y(O����O��D�<A�'�1C��U���O�(9����T�*s3�x��'dў��hHXu!REZ�7�,e��H�4x5��o�埔�'K��'�B�'�"�K�����uB|��6�R�<�Z����Dݛ��'���'A�'��Q�!�t������;>��1"�,�l)At]�����X�IbyB�V�F,��b5��Ĝ��S��I�$�X�j1G��	ٟ4�?qf�O�'d(<(r�b��&Z؄����!$�o���X�I۟����$1Pp������I�����Epm[ x�J��ќ8>ܱ�M<����d�����!Dc6$э�z�&ZEFW�)�N��?s&���?���?��������d�J�hrh�S��)sաQ�M�����Fqr����e+F�Ә�b*k02y�f�iе�5z�����O��$���L'�\�	,[s��`-ƫ �:�UnB�d�����?Q�,��p���������J��`��&�'��'� 䊓C7�	�����q>��ǪGE�Q��EA�>��Ն������x��g"$,Xl�!͑�#enѺF��Mc��Y%�=2E�x��'�R�|Zcy�0kd���w�.p	S�_M
@��O�쒦�$�O,���O��"��(&��A�T!��"����J����'-��'-�',��'�BH�QAؑ4%�$[�AĘh�F@rt�L+��']��cׁ,�2�HCӮ;iv��'��b4�	�ݔ<f�0e�!2�:Q�ɲ	)�щ!��~<��@��>:gp:�%��O.�5hʢx1\� "8��ǮUX�*
n�C���X�a9��G�/��\a�a�;z��0(ի�*}�(���_���B&Ԯ2ݜ���'2�9P%����]��J�<$ |K��П{H
՛Ђ�=�L��2��{�ʌȴ�� �]A��V/��y�/΍B١�ҙaK�MS��M����G��� t,��h�!�	?(�|}�e��+oY�����Ρ�D���ϟ�rdCԢi����SKM���)j�E��?�Oc$۴�J�,��v�Ե%ݶ�H�̲`�[�\kd�
��@�R�
��eǋ#����M?��W P&,$���¯�p|Q�!}2ə��?i��h������0�p��%�5S,4a*b��,!�D� X�r5�t͟	2d�8�GaxbD>�74�q�%nU� {�<��C�?�D{C[�X��䟬�����T���ID��ޟ��=,�J� 楎�GG�U�7EȲS��e�W?��(6D![��>�3��ם$��4�H��FĹS_�[q�EH#�Ř��$���d���L>	�/�' ��E�a�]�4Shq`����?��O������d�I#s�:A�� ֽ5�d���w�C�	�{�0�sc���I����!���P� l���'��D�/4���$�T>
��}k���E#
<���,2j���O����O���;�?i�����B(�8�P�*N�aS�H(��(hw���?�Nm��2lO.��6�]��*؃ 'g�ŋ���*z��
pl��.����!T�8�E��3��+���L�-HD�O.�d,ړ��'9�e��C	9kV%3!��x3z�K�'xT�䍀!�1�'�� ��y�ȥ>!(O��v�k}"�'��3�ju-b�{G ��tW4����'�R�ńwr�'��i�O���y��?R&�-��2��#ElQ�G��d�T9���	%r��}C����C���'�lx�E�ߝM4���a
�'c{XU�
�|t6M�	�$�'"jmS��&+v}�d�[�Љ�y��'��H�mT�U�`m8u�TV�>���'^z7-fJ-��B�8�\�Z!+8i��<�5@
+`�Iꟼ�O������G\6�t��c�~a k%͂�i�b�'-6DA��ݪF����	_}*���'2u�W�Z(.$��K�Ʉ�B,X��O�zbI�02S@�z�π 6����	O�$4{G����LsQ�>QƎ���h�IJ�O�I;+iڵ�#燵�)��[�y���#�X31�����/�0<�鉾�L*�D��(������Y���ҭOT���O�p9�DM�����O ���O�n�3)`&�j�i�3�H�.� v4��@������c�t�XA'�3��'���7�ݘO��`�
M���ٲ�_, ]��=y�!�W��|"�y����0��dL�!���m��7Mwy�!�?�'����DL`p�9�nD}*��"���yRT=��Q$�� Mi��	��D��'E*���D�*�$S��k3�q�$ۢ����`��i
���O��D�OF �;�?�������h�|ՈQ�˿E������?!(L�E+ڔ�l4r(Ô�0=��G/GҺq��KQ�HU�d�i�W$�Xs�kX�����CCk�����2cG���V�G�b<��F$kW��D�x�4��'�b?���'..���l����pk�E,D��8�K�}�R�ېBҳNh�d�0�	����<aaO��c�&�'B+_{~\Đ�ɦH��"d`�����'����4�'�:��x�D�'��'�*Y�cN�y5l�3�
9}���>E�?٥.��scFd��\�:@=�%�m8��9���O(�Of�`�A�9�4a�'�Z+M�I��"O�t)d�J%J ��K��׳i>a�O�n�?"�~���N�9+F8���yX>b�t2O�*�M���?�.��y���O������"�R4�7!�T��#��O��$��Mz�D1�|�'�@p@�D/Vq\4)P�C�a~"��O���&8�S�'-f���u#��)}>)�"�W����>}�g�"�?��y����$Ĩ�����L_yc�,W��y�ћ�F���=Hܢ�Y�
X��0<���ɗdT�	0H�#t��PΗ�6�BxA�4�?9��?ф�U�?I֩����?��?ͻ7�%�ӎ��M����0NгW_Z�q�yB�ݨ��<����q��ڡd#D���Cց�_ܓz&���I� W*}�##�]��e`�b�T�<!%����L>1��A<�1qcLVZ�HE�R�<�A��&>�L��"��`8���E~Ҫ!�S�O���`�fӖ%��	00<�PԠ��L4�Z��'R�'��Fsݑ��ǟ�'1o&E�tk�%BH�����;��ǫ_m<����n�p�)���7���k��J�q��!��m�pH*�!��v�� i�$,�<� n�埌��	 +�zQ���6n~̠sPI��LX�B�I�*�XՄϰit����11�db��}r� �,�7��O\�� K��	hqn�*�Z�B�
�34�$�O�1e��O��D>���ON�O����I�68̽�'�����&�'�P�b�X!�d�8�-A7G�ʨ ���-�p<�a���$&����5�X8r�78�e��h5D��[D"�/��|`t � 'J�1�>�H�۴>�8L!�ϏPѮ-)L�/p3nM�<�`蓮p2�f�'�Y>�d�ݟ�auF��)i�H�Łˍ@��T�KUߟ��� xs`L�	e�S��O���G�K�,��D�h����>a��EP���O^�-�B#M=d���b(D��9��ɳ=_��:�)���M�"$������X`��ʽ4<B�	��h%�'���H؂��S���F������B�'�.u@�K��(�1��h߬L���̲>q��?�0�)E��!����?Q���?�; @��˜9�F�FJL�4@Rb�E&y�I��Nk��xa@�U?��|b%U56�Pia�&�4�Z�22W�N9��+�,.�l�e4xQ����|r��9Y6�t�w�D�w�p��H�)�"����W�O�i�O��P�t!Łp|K&)�JdQs-D� ��F#h�H8��MѦP����`*?���)
-O�Q��Z3<�P��@]]��}j�A@:2�1yd-�O����O$������?1�O��x�wąB����&�ط ־�c� ʛ�x�ɞdc��c5 @�d�)���eS��k�'d��[B�͉+tS�	A/3�2����¢�?�
�@�����cH@�Hb@͆ �@Ņ�k4�0���4=�����P�y%��<Y`�K�4��'���"Y�.�2fE�D<�m��8"�'#D�S��'�R6��i���I&���Q"��ē���i�zTYu$[�x�*<
�Z,�p<qc#�Z�����
�X�dʣ@���I� ��R]�*R�-b���C<R�'z�)� b� P
h��snÌT��X����O����(��A��&p�P��M͡q�!�AצIDEF$y���c�Z�z'��� oo� �'q���Q�c�2�d�OB�'j����A��]h��&*�쉩�+G��TA���?!�/���?y�y*����[��$��GG���`x�aH-<��'n������)�� ��4�S=!/j$80�;;�yF^���H�S�'TG�Ի�I>TZT��0���ȓ6�dn��~�<�׷x�l��	��HO��ť��0(����r^��p+N����П��I${���hC�Ο<����i���,�*G�d�3f�^	,Tt8��@̓5���$�O~D��Ll�<PQ�eɚt�qO.,I	�	W~�hG�e��� �֪�������ҭUm����?��9��G��"����l��y��'�D��p�����ɂ"� Z���OʸDzʟVʓA�|��ԇ��a����*0�̥J4��\��	���?����?�ķ����O��)4^\"Cɢȴ��s�A�`�c)�@[�a�`FС���y�4�Y�i�a��B�	b��'�E�ʝ��ӣA�����h�O����J�8�
�`B�AvTԈ'HȹC}!�D�66@r��ղSU�Ȃ��z1OM�>y��^�B���Ο@1�I�.�84��.˹"�ބsd΋ş��I�y���I���ͧ����'��R��ώs�R��VMW:H��Q)M�:H���#�p<�У'��h���I2P�����k;00h�Ԧ~S|���&@� W���D�|?A������d�0%��(K�_��x�6�V�X]1O����dA~�9��_�H��Y@�D(W!��j�DK.8��з�z��[�\9�ĵ<D���o����'�b[>9�$�՟X��bʻj��Ā�!�kҠ(aT$�Ɵ<�I	o��uK�R�S��O�y�f��3C$t[��ȠW�����>��!I�w���?�
���o:���f�
0��� "}���<�?����䧔�'?]�SU�IZֹS��(q�<1����<���J���F`W��`��$+]}� ȏ�Ø��X�5�N*4�*1r� �V�:��'��'IXiyG��ND"�'����y瀈�O�����gٍ|��U:�_-z`D��6+S$y6\Y�D�^�v$m���i�~�dC�fߨ��$d���7Ā@��j�)����K�N�����y'��f�D
%��})�(D%Yx4CR�E(���*?Q��Hß�q�'^��i��)�|���ĩ$��0�'���Apˈ�����q��f�����O�Dzʟ˓S�n�+Q���"4�Eo�06z�)
A�,>�v�p���?����?!A�����O��Ӕ5�$��`�@�>m0 ��O��t@�
O`��$�U���q�F� 4Ҩ�r`f��PxR���xZmR+N�	td��4B�*pJ����?�H>������~�e��4�M'k��-PЊ�N�F�<�ਜ਼
(:��3Z-&�!��|̓%��IIyb�PZI�7-�O��ّ@�ʽ�$2D����W,����OR ����O�$}>�aV��O��O��p�kz4�W���3�TW	q8��e�-�I!�X���g��2R�(ԺN���G�1��|���t�l���
�	��yr�N�>�b0��sK�#`N���x�q�H�ZbZO7��	���$��(w��E�*���'�bV>y��^꟰q�IW�PR�(4#ڊT:D�[؟��I�c\|I�f�:�hapԭZ��?�O哋!�VtPE���]�So�D$��'u���ES3����2��Xv�>���S�9�86	�mJ*@dk$}�?Y��i�l#}"�'CAB����F�J��`9橛b����'�v���	�Ԥ�E�6b����������ķA\26�����:~��F�'i��';be���@��B�'x��'��#,��Y[�߷[�t���'�4�<��~x��ST��&2����&j�t����1�ɛb����_(c��IP'*T�J��D���w��c���D�Oq��'K�a�1JJ6z*f�0w*�Z�ȸ�'^Z"&נz�����-�i0�O@�Ez���Ƽm����"�Ch�Ia�A�&e�D� J:B-
���O�lZ؟ ����a>U�Sm��rҔ�"�J9=C��2A�Hu��2�O��+��0
��(!U� \l��0\lE���(�h#t�('� ܰ�m�ş��IΟ���ay��')�O� F��� ^?UN��4]�Y��@�"O�S�D�	3�i�F�i��AAA�~}W��[��ÿ�Ms���? �Bj�9�����`��q��鞵�?!��9jt�R���?�OSH������B(<�y����P�$�Kv#�PH���	�-���H�ViB��tE�����A�K,Ot��U�'n�'�z��A$� �N-
G䀖��Y
�':az��[�9���6���>��	�'��6-�{�������#
��Th��)�1O�I��E�	�I�� �OH�4�'"�ܚ�b�#9���`X�P����'ObI��mi�T>�O����c�'=�L+�jٶ7]F��OF���)��3 �`�����U�8mvB���&�'��q������O�:�Zg����=��o�SRF�'�6���E�~�����I��<��HiÓё�� ��3��� b�P�h8#�,D��!���_�z�8cՈx��S�0D���"�[���Qoئ�rUz<D���%6-o m��LL �J��-;D�겎M�[�\�#U�y� LӇ#$D�tٴ�R�#�)S�Q�U@���#D�4#׍ȻA.ni(�@�4 �����L D�\"g�ř6l�����ƠL�-(�G>D��Y�gG0��$B@_�l�����0D��*��v$�3r�^�.��� w�/D������O��Ix�5Kn�kWJ,D��K@a�"c}~��V�9)jD*�d)D���A���|3"�8I�b�xi'D�`C�G݌[GL�i�HU�
�L|�t%D�0����	u�J�ؐ���f�H��M(D��rk�&��yp�Z�h�@��&D�tTB�rGء@ę�IR~���#D��
�.k��u���$�|$�a
!D�p"�l�$:φ��Ud��!l�t�c�?D�$3���4L�H�
�b�l�8q�>D�Dy'��#�X�^���awm2D�\����A�*�W!��'"�iR�*D��'ͩuŞ��ӈ�l�ֈ2��%D�H����z���2�ْ@�h�*)D���v �0i��B⍖�1�Rjr�'D��+5�sĞ�@V5&="a0�8D��5�K�L���=3߮�P�6D�T�R�ĪTe����Q��@Y��6D�0��f��)��	��ʑ�@98	�c-4��A���#������'���$�<m�:�B��Z�D�00�I��<��C$[�D8E�#ct|��,�\�'Pz�����E��B��rx�!9�O$,XP
f�������?�W��W.�:<8�Ņ�#y�i ��OmDr��§ӣ3�\i8��'�B�8�!�I�z���B�(>��� ���%�)�'y`�}B"�µE��%����f}4ݐN�d�ax�'�-LTp4����	�3��|�Q��в;6N�I��?}�`GA�'��%q�G�Q�0LkG�
�"~��9�FǗl��q�P�$�,\$U�4�j,����@;]���<�TD��N#,���H?r��!ȡ@�v�'Z6S`��(K?0=և�:�r)�'�B�x�H�/���3�28�P���'ԮG
Ġ��9}3\!���O����OW���+��NbDɜj���y�^=��h���h�rAO�g��E}��eh�a�Ft��iZ�a� #!���6�(O�>�kT���`V��	%U������zHb�1!L�8���4�J1�r_ɼ�B�L>X۴%�D�V�N80�F��@=��=�ÆܪcfB���-a�������'��T[F��G<� �DE�w����I� 	���{J�|8a�ڥJ�\�3��*<O�}:e�ʅ
9\�1���0Hhd�ՠ­(���ȇ�"k: ��ɭ>�3Vtl[�	���2�hT�Ft�'�BY��/� u��#�ʒ��<T)��D��j�����O����{���*GnR�b'�*O��I0A��3X��p��OT���|�9K0C'	� ���U�$ք�6/��D�tp�� �	/�\tiD��օ�2'e�=�iX�:
`�VF�V Ś4a2��!eN�*��B�]�* ����P����2mH(����O�;2T��q b�ɱm*?q��ȴ(b��īK�*1�Ą�Wy"����'��$�/�i`��;LĦ� ���R)1���i�I�o���q#�I	o�1���v��Ba:w�ax���N�����)Z�O� " g����I��?@�6)+�����G6�>��JqΕ}j��R�+�:A/����@�Tg�}�Hc�7��UE:�`9Lp���13*ISQ��@��� �?��?��?q���>��������ѐ���	��b���'��`��dD��Sm�K�`,¢��E�8c�h#�O�����F�=�,ԁ� �O��'@���gAy���ip,V�9�^�9�'Zɹ��FGbԛW��C������%���k@��<�l�S��*�SV��F�h���F!11>���(O��Ҁ1�pm���ӑ$�:p�%
)��'\h��G�������R��=���ȆG�:�bh�C�/;R���'�p�Ey���)޼��?��,H��;n
L�3G��y��]���ޢ\a����O�
M�7O��S��&l��!
�����`&��Y�$ߥ��	�O��Ez� Ҟy�zIإ
)Y�8��D��'�����EQ�}s���C62-���?�I��9RP��X0:@�"�̃f�����*���D|�4nB�=jңX,D��[��7�Xi�� P�
sFX�1���8W����Qìp焴��w-�O�h�cL8Z�)����:?-�(2��H���'
L! Va�]`h�x���v�C�b��d�[�A*V�V+"F��1� ֹȖp��0�I/$�8��?���$`R B�W	6T$�*�$�=��M "�4�z�b���7M;�'�xaÖ条g켪���$J�� U�,���u��˟L��Rkoy����a�\ m���f� �Dy��K�Q���~��+�>Q����_�iB@h�0�[�m�F�~р���O�)�@���l>x� ��u����aM]ش`d��w�dӺ�O�Q7v�X�� Ns$Mj���`�ʍ�P.�$e�*�
�D�ğ��̈Le�IP2��@�뮉��hO��c�Γ!��
ާ^�>���|�2O>��$� z��=�!�1O�����އd��D2`��b��X�f���|J�?LO,U��w�- ��̽:�L�ޞv%�KƎ�"0��ݩ������k�2ݟ02����`i�m�X7�<B���iĆ����Q���q��1D��]i��
p�~�ᇮZ
�>A�`˵&�0���׬Q�~騡��џh���V$M�+E�&Ww��+$��?�A9S�mpI>��O�!�S@�;fn4]�R�O���k�(>m~���Ȏ�Z��N#��D{j0���hO��"2P�[����/˸2qx�{�V�l�ɽ(����q�:9?����7�s����p,�+My���g�0X�0��P�ϛMG��А�?O`���"S��svƄ-Պ r, uΤ	���,g�`M�V��!bGb��2q��p�����d�R`�E�'o�?n��5eˌB7�����	pC"�3�Q���aN���ä��<O
ꡯ�RU�@�m�Q��� �^z�Z���JT��
U���C�9{�����ꈳY�Ь�Q�ig��j����cNf4@�jV�X��D�YPb���v���=�ܐSu�қi�%�թ�O���O8�I��C)pS����'��y��ٍzF� S@&�=�̤h������� 6����?QD.�}e̥j_�M#c�QcG@�!E͆�3�J:�F!�� ��<yc�_��y���3��5��nX"s�jћBa�5��'�(���u�TT%?��XH`�NA�:H]�P�R���Dz"��+�$�y�(\=d�Q*��Z	���!p�:����@.�$�+�!X0+n æ�HNe�OVݤO�U���� ����mA�iU�O?��17,Ҥ'�*6��mh<����0uf�D��LM%���� S4A�$!��Y�Z�%�Ĥ�O0D�O��IB�Y"�����'�d��w��] �-`�@ v��r�AV�=w����C�����t{,�a�'�I��.ծW��AA1�>&���K��Q=~kR�D|�b�h���X��q,3Go�Y dJJ�к �1`0�DZ�VP�!ʱ`�2�>���� ��a���#]�u�Uf]o�'=b!�'�$q���X7!�n�[�'K:T#&�?D|���]�=H	���S"�>���A�e~bS>��$��MoB��EB�?e�&��U�<���5pp4⢋�O�i[���#lL`�In:(d��>��n~bE�8H�P;U��N�|�s0h=�?�����갪���G&ѡdM�l*S�%�	@'>�ˡ$G7x]µ+�è��a pꃞ\�ru�'#f����x�M	]�F���W2@��ñV��yK�玧@x�1�+S t�8iA玗4��y�����ywo
�	��m�p
��r�f�y�A�9C����4��6� �j3�i>�;c��6\�V���O�ӄ�vA����NwB	i�cT�x�8DD��B��ɈPy�P�j�&�����!����u+
�=g��c�P[��aX��x~_?A&��7���w�\^�E8�>q`2�<s�ԋF�r�d���I�4-���'�?�7OY�(� �MҠl���)��3hP��pN�8<v< �	�B��0���#���g��,%��g�;�L�t��Y��B���vF�x��,�p�!�� 4�H kc,��{L�p�	��M�|ڱ�۰"�$�S׈��t�Z5�a$�'"�)FAR5X(H��'i�q���T���b˕�F	
`���^:gj�}BA!��?i������R>Sl���?)É��g2�qYt��Qk���,A<)ǁ��C�0�MP�VӶ��h�M�
8���zQb���uk1e� ]�\� ��?�J�-'E~ٰUj҇j��=a�3O�9+�Ö�>U����Gp$ؒ� �(����E�e�SOƓR?��ҕ�'o��)UlI&xud=+�L��)�*��O�I� �gް �ˏ7[�h	�A�>aEF�?/6h����I�d����;��Y� ��BI�w¥7�@)x�hѫ6C	����u/L:1�
���I�1),�j�B��$���B/�Lc�$���R1oJ���&_ �D��|2��O�<I��胪f�dJ�	)H���'<H�U�B�~� �ފZ�(�a��is�6m�?t�������J��{��?7��b;�T��mSN������P��t����'
q�GWo�pŎ�igL�MA<0�k��vMjAS�|?	�葡[T�iVb>��.�F��R��%��nޡ�9� ٦}����'�"�q�PR��|�Ɇ=e��)qH�����#�T�d��m�o=x	0��O:N��BaA���=�'Y�)��Xp'դ7��h�W��x̓w �i��<␤�V�ܠE�RL��M����D��!�� +2��	<-~C���CD�:��Z�nHK�䕉>��M�dM�O���eN��T�^���#̤
V$�I�fh'?�8���Fw@����[�xaDؕ,�����&V?��x��	g
��t�:���:.� `S�8]n�AS�-N���i vU�`����|F|҈A!hJP棑7���@���~RJ�_4�S�:[�(�� I��s��2�Lßl�p�J:+��P�яP�g�<���ٶOw������ڰ>��N!�x�"[�C�\��z5��O�ĉ4l��<��^U*x�&K\��:���gV�#�\�VF_++K܉��'n�퉐�?|� ��DL������h�j۴#َ�)�ЈB�ҙ��
�����RP�*`'����D��,� �X�B-7 .QSL��4�<��d  Y+2A��Ѕ@�
�P����� ��j�\|�8���I�
�"4	Чhö����'��q� �P |�24��9��d#D~��Ѭ�*e�E�Ӆ/��G�a�HԢB�=�\�na���0������K�^�a ��v<m�ƣݸ8u\� ���][(<cC��/�ڌ�W�%�O�a3����s���`�J�A�a�)�G,��M3$m�P���L�O�x&>��w���^(�Pƌ��,�
f��p?9G��vİPb�DIu�8�0fhR�Sv� �ԭ%6DQE��CƦe:g�x���L�p�0�����"8)�O�3f%�dō,E�`���<aǈ��`�%Wr�(��F[#��4�V�J$ry4�#7�7o|Pxr�>1Cf�//^,�����YJP�@&�F��8�.���	Đ�pcCG%`��ئO��aƇ�* r4�ĵ`0<0�&��[�l� $O3��\
�0eY��2�ժV��@���C�R��	Q�-�1\�h��'�l�إ�H�����v�#��޼=�L�������C��"��֬�̩�>�ݚI��Q	�"��-B��.t�*C�ɦd��c���n�@Ys�Ťu-`z`�B+|��<���A�����	kZ%��(�>sVu",RzC��+��Z)q���&�-O�-���ݕ+%� f�v��	�`C��0n��v��'�A1uJG�?	G�,7| ! 4't�bK�N�'j�m�����vNp��Y&�ȂI����)F2L�Kݔ7�1sЦ�)��� L������U�D��$�ڊr�@�{w/��o*p[��'	�T4��V����Mʜdz��^�s*(c��;O\�� �Xd�'����2�ҭ��Hx��`��T�PQG
O�I��m�_|��:%͚;�ڬ���
Tf�Dx���X?�AqZ�u���[c�5�~b^�KPd8���D�m������а<1�a΋���8).�2uC��.�{C,�Tn����O4�+���wD��C�� �0q�I �l���ı% �W���	&��䓂RGf���ON%7f&��PP#b�bDj�M_	�` u�S-jX��f!V�F]���� 9,��qSq��N�- ��*���,X�I#�)��Q�����V0|���`f�)N.�C�Ɋ9�,��1i_()h�S�*�����=I�O�ر��'o`*V��'>mª�����
�'�tP6M$b��p����l\��6,I'%S�A���=!�@	�͆�;ϖTS��M1���Ė�{O�c��;���o읣�$��%~0h�7D�8س�/d�lQE��:>�6+9D��"r)�ɨvET5�6�F�7D�$a��M�t�(R���8 �,�A(D��Pd�����̲:��aB�8D�(Ю��mG�Hsu(�:�٠�,D�@;�N3��\�'A�!��{� 8D�x�1%Q�&@�4+2Z�+���jm5D�L
փI��(��K̪D���c�3D�|YC̾Kw輹C��R궱�7D�8Ctkz,���
.�@	�� 6D�L#6V�P����2V5*�`�#2D�t���<'�α`""��dm�%qGh0D�� �i(�Ŏ@�r��2����8��"O.���Bĳ]|�pJE�I߶�"O��ge�:}�����4SĜ5�"O�x�Wf�5tx c
��_TNC�"O^�9tLr�I��nɍuk�B"O=z�l� O�@�,Q~���Y�"O��qd#���(M(���$p��uZ�"OB ��
��b�u��	�(���"Ob��^�i��b�ׁ%ʥ��"O�а���ְ���A�a8� �"O��愝&lnxa�́>��� "O��H�(%�q:$�]&9��7"O�Há�^-	��H��ݺc�.��"O~�2�ŚeV�0�� �v�j�"O�˧CW�za�Q� �͒�%D�T��#V���9q!���HF*DH�j(D��c��	�"9��、='p �B�!D�tv���&X���-_���c4D�Ȳ��[o�>��6�D�y���E�1D����"t�壵急VE �w:D�܂KצB� �Ġُh=���c�:D��1@���;��h��X�u^H�둨9D�hSe�N�O �T��DW�*�y���7D���tL�{�:��)��	��"D��	��Nl�����X*�Ua�L#D����)�SH"�b��ޡ�n�q6`!D���C#�U��,
��� d~�� # D���ՠ@+�̹K"��	�P�( �>D�d�W�I�F	`H�A�"<PH$R�f!D�<�AW
FX]��eS�xkx8c�<D��Q��Ţ.	b�����4	߂%�Qe%D�t�fd�[��ɚdȐ>��p�$D�(�D�G�I�>�ɁkN&��U�� $D� XA)�R*$��GA�(+�0�@� D�08Sf��?]v�br��$���!�
#D�4+��_2 
����:y����=D��b�'ډ~N��CVm� v|d���:D�8���0�]J�]�3�c�!���+")�u�Ѭ�Je*АE`:�!��SC����#�Q���z�.P��!�$@�i�5yo�w� �$L_6�!�$N�Z�*@ �� ����$�{�!���l����.V��uhp�>Y�!�d7SԞ@3%S<�d���&
>:"!�M�i�eی?D�%Rˑb�!�Em�e����	*���Ū� !�OQ��׃� �=zI��V!��:,��<0ƪ�-�� ��;ء��@1��#H
5� ��1JL/l(^B�	�JYJ�k�հ"�Ha��K�*B�I'��@ජ�/}VdS�e�n��C�?k��d.�<$&:�CĎ�U��C�IF�����A���)��C�	��Ė�A�FIHE�ϋI�p
�"OI3F�^2G9La�� x�p�e�'�ў"~"�Ӕ�8V�� hY�G ttB�Ia�>�𱄐b��k���-igf��$h�9q���U��`����g�yҌ�8_WB ��C�%w'δY�@��yr��1�aO���TEO��Px��i�$51�P�H<���r�]�a�.���'4"Mba�A�F>�)�*Y�,�:��2�S���J�Fl ��.���,�����)�y���K��cC'EA����"��P���π ���e���i�X8��A�X�$�a�"O��Ʃ_�c� �d�H���ב|R�'��}���ٳp]:���%Z�@,i��'kN�h��ܸv�e�v
ȳI�ڜ'yў"~*pEZ7�F� �dQ.)����N�<�Fԓ)�@:p�Q�Q�%����s�<�AH�0JJ�s�)\�L���R�HF{��i�#Ŋ}��i)H�.I��m�C�$s�F�2��H+�5�7�Ԙ�C�I�)�V�7�ܝR��D��:�8C�	�OZF��ǭ� 7�2p9%�@4xL2C�	�Z�"L��-	�\B
�9�+��I�0��hO�>U�%�"@��0;���d�T$#d�3D�Z�޺4� �͜�Gd<��2o1��6�O�q)��ÍE����� ?~`bh{0"O~勔MM�{: ����ގ,W�q��'E��X怅)@(�/�ًu�L�y�!�dܵg��k�eХ/�����+g!����ykq/D�jsc�;wR�F{ʟ0Y:��ա'�.���៛V��"O$�R/��$k�D-'���8Z�<���'��9i��׼O�dkF냩Vt�����$\�%�h���ű)'~���D�/&!��=v��@��+q
i�$$�8G!�%B,�;�E�8
<�.	��U`�'��|XB���)#E	�E��>Tp�'����#�l� �[�`M����'ȼ�S0��l���1�" �zX�B�'5��tה*%~ŉ�SHX��'�5"bٿ+�+�usTUk�'+$R�B6NNȀ�,�>|l�	�'�J	��V2� ��-�j(B
�'�y�E*ˢPl�!�J<� ��'5r\�@��2Kezy�P$P#����'��	�jM/Q��Q��3�6Ѐ�'{H��Z7�.��S  =(
މ��'vt�`TMNX�t� ئT6�H��'f��1�(�P4���R�U:�������OOe��M�b!R�M%�H��gh�Т�-h��UB6�T-r7�,�ȓuxPb�/��!F��+iݖ`��hC�P+�R"���פb�>F{��'�a�E��v�����R;/���2�'�����*S�#��%YUI�"W�Uq�'(.lkV�T�`��]���!u*�Qx���'J�(#!X�F_Z��c	��*kh�	�'\�q�جE+^iqs���)���')���ƿ{�34bPB�6)C≝F8���a��d�z��j�n٠B�	? �~)XV枎K�N���PS�B�I�C��Bd� T@�FR$V�C�I8tĨd�׋M:]��)ϓ��B䉀/�}�A"��	��*��B�	:fjyHw���/��$�a˚s�P#?�����T���pF��+T≡�2�!���,'[�H��ː�N;�0�p�O 	�!�#(�ؤ�s��'9X:��	0K!�d�O��� ���R�|0:�)�H���[��'`ў �q��/I�$4ʱ.M$za�2&�OP�	�$��cr�I*\���yU�@ bB䉝@�45���*2 �Fcɛxd.B�4C����tg@�o��&��'�C�_@�,�T/�9X���w�NX&�C�?*LD]�Vxx`�K�\��B�)� :h��/� j8&�s��',N&�+E"O e	q@̂Q���	��y9Tq�B"O.�Q�ʝ
M&DNH {e"O�@�Pc	�(�M�'jStE�D"O�d���2w,P(h�ڵ|�:(��"OU���+8��jv�T�u@\� �"O���Ǫ�9bq���2�4 $Z�"O��Ƃ)(�a�B+�� ��rR"OhY1� B6���k��,@��"O��2t[6?T6���U��k�"OP��u�J/Yv��$�Q6�&�8�"O8) 7��*E_�� �q�T��"OXe)Rhޟ>V���L>B�ȼ��"O�[R	���%�Ǝ[Ep�uk�'
2Hɠ�5f�$��3c�)B�8��'�T%��[g���b�ʞ'�d���'uf8�b�V�I2��Z���좍}��)�)<5��m`e�ʹ71��bW#]1�!�$6�\���j\�t��A�Uc���!� �G0"E�rl~�yC��ŝ3�a}��>�Uē�>xF��+��ET�]�Ga	b�<yG�l<\�S)B��H��VJH�<sg^�.����1�ér?P�A��Sk�<!��ʰFXus���+&Y6�AD�R?����S�dR>���됷J/�(a��޶o�fB��+N���srJ5 <��AE^�(B�	�XH<�	���P�(a�ri�iT�C�	, ��4�T
ɾh���"q"��#��C�-�����c��c;�5�C�0K�jB�	�H�ểW&6H�5��DR�.>$C�����+�&�3y�jek �Q.p�B���@a1F%�24c(M�B�O�8!�B�I�<���I &��TՀ����B�I�i�,!�D�i	,U�g*�1{��C�ɿ6�����R�*��#��o�!�Đ����˰nVdӰY��ˋ�����	�T~�u�2+]"92T�&۳z
6B�	�~H�J�	M.x�VP��ډvhC�ɓ"�j�����bxhd��r'�C�I�nI��x2�^�-�L��F#w�C�ɛ���0tkW9���H`����C�8sJP��U@rFv�Aa��!� B�	�j�.�`�Ȧqe��ŝ���C�	����B�� )����[�O[�C�I!,D>tV�E+
�n�����C�I4�2p2%��9 9B�c̽��C�ɶ0�1	�	ȝ=k�HvA�� C��J%�#��7:�A�����i5 C䉪bVNh�#��c��M۰�ߏZ��B�I�&4ѣ���)z�h��S� :�B�	�h^h#R2&q2e� H\p�C�I�lZ@�҆�qD��׫� J��C�	�IYz��-�(�LӅ㗳FX�B�	#�����jJ ll���-��+��B�	%h&��(��̋#��E�c�V3=$2B�	�PҎ��i�fε��ּme&B�	��>���,�P�|}ؕb o"B�I���)c��*�N��b��V;B�ɜi�0�� l�:�`��^VC�q�8H���:hY���,F�B��*uV�1I��.b���+�Ç��C�I�&I*xP�ҏu^찰&f'��C�ɌK �qR��6B�̨�g�^�JψC�	"D:���be�5!��8�C�9M�B�)� JD��O�={&��u��X,*���"O��+��ϣ	m�!a��FrF۔"O�e8Ĉ[4��eJ���*>g���"O��!-C7D@ �+�t0�"O�� B��mQ����
�} ��"O� ��m�TY��2�+�!0\�a5"O�R�mڔ\' ����R���@�"OV�!�~�0܀P!�#�L�ba"Oj5HRh��+�TԐDʋ����S`"O����6%fQ�I�5M}l�"OV�(��j����D�!e˦x�1"OB�㥇����2h�J����"O� !�-�� ,^̀��x!����Nx!򄂾�t1aG�#g��gZ�j!�D=����R�:STy�E	�5h!���N�p!ё��V�F��31Ns!��N���gζD�Z��M�p!�N���i�jMG��l�B�A�}g!�A;PƠd1�O�K��A%	^�UI!�dP�5�\���e�r�ZH�Q#!�QR`y9g刪xp�<�#ǾU!�d�'*Ɏ(��.l�@$r�(5�!�Dء8G$iy�0 ��=�ԋ_9A�!�ُ��LK��!x?
 #�M�z!�d#(_�⢎�9.�ԩ���	%ij!��̣E�rq䕮?���� �@D�!�[�f9�|*�=8OLa�tKZ�"�!�-&���g�#D�a�$kJW!��%}�����X(r�(�ů"�!�d�s{���h����1fȚQ�!�J,�����1&2�����f!�oMl�1A-�1����#A�q=!�> g8P�H
�n˦(�A�^"[!�$֥5����'Hb��(�6A��H!�X{6��a¤߿Lú������!����&�)��0�Z���!R�H�!�$��������c�TiT�IE�!�$�9�l�J'Ø�]�\0�'.�!�$�"4na2�g *`��<�!�D@>>�p3���
�����7�!�D �{3`��	\��E�H��&�!��S�5?�y�@�W�hq�$��w�!�$W�HŞ�"�&	 Q� �@��ƌQ�!�Dϵ��#n}@m��,G� C�ɑcXhl�s��'Ob0*�b�z�B��<Wl�`�����ar0<��	A�w��C�I�w��a'ܗ5BzT��z�C�ɺDP�1i!�7:�X�3hE ]��B�I�6��H#���8�k!��86~~B�ɒI^�c��[6�aa�DIh�C�Ik���ҁ /$��y��G!w�B�ɏ'e��ZSg�g?�q`"�.Q(�B䉑k�R�r��ʕ��E�2)A�ɆB�A
�`��N@�� �o]<�hB�	�<l�x��e��)z�CAV&#�B�I 4�ָ8���j�ڒ���;�B�ɳw��$��/;0!�Q����C�ɥ2`h� �
=*];gH׳4��C�	�T���5�]�<�cB��9/�B�	y�Tl��	�r�q���B�ɼp��2��9��(s�
4h�B䉬1����˅�y�����E�j�B䉗V�4�p�Hm�4�ؓ��'WZ�B�8+��{$���&P�˙�
�B�)� ���$h�p�RQ���a�
)�"O��G�O�
���gՂ�"�	&"O� ҀגO~�T:dG�<-�dQ��"O:y�d���؋r%�r�N�$"O��J�N�?��<��*	�^k�,�r"O�,y��ä�$e
��\�؄��"O^�cb�I�k��q5(K�"��J�"O ,��$ͻ?z����Us��� �"O\Qq!c
d{4X�e�� #BX#�"O�E��iA
w��X/�\y��u�!�D*Z���&ְY<h�	'�Z�!��/#�N�E��+)7|�A��N�kf!���*5�r.�"%V����M'J!��4e�Ш���X�R	p�ڲ�w/!�d�a� �a�)-rX��
�E{!�I1>um �M��A�ZeQ��Q
H]!�DH�6c�J��u�P�ϼJJ!�^<N��IxU�K�P��@�#D?!�$�9Z�\�I�b���L��`�?E!�Dߵ[~@JE�1(8�җ!�$�7\��`(��ϸT������'�!���d|���)�)WJ
�#���!t�!�$�mY�\h��Q�I%đQ'�އ$�!�D�d�z]Ip����Q�8j�!�D�6J�hܲM<*e#Vd�!���$B�����L�bqڌr���!��O�#����dA:Lk@��'W=t�!�d��X�����ā�)S4��6N��!�ě>v��-��Z��Ҵ,3H_!��ӑ���z�$�>Zp�&� $�!�D��w�"II%哷 �����$/�!�dI�Lvԁ# Ȃ�T���#g�@ �!�V9Qn����k�I!�g!�D�	l����Ȅ=Va\[cB�`!�$�7w�~0�P���y#�mX�o�!��[�[�t�˧�H3
����m�Q�!�Dϗ"���q�&ӹ0�PJ�/a~!��ʨw[d��IO�mޔ���
�rj!��|��<��ΏP0�f�G�^/!�D��A��o·-�Xԑ�*̳Gq!�䓣n�L����8o�
9%+=Xo!�M=��e���7QH1�D�ʂ9k!��ԍ-��`sG8'b$ӫ�a!�� a�Z�s��^���ܱVkŰ)�!�̪k��X$�.�� [�*l�!��%;R���F̶1����@j!򄊮@�m���½g�"��t#�jE!�$͕���WM�j�r��٨@!��)K	NEz�E�`:|r0�58!��`46Ļ�c�=dY~,&Ač)!�D7]y҄�0 Qf!�@��!��]�+B8h��#����(��g�!�R�~�=�b W:��i����-H�!���Z�.��3I�4��I�֠�=�!���T�0`)F����xA���v�!�DG�VBֵ97`EA�b�Rf�, !�ٻ[L2�ȉ�b �����ٴ>!�$ �e������92~���A�m�!�D81���/W#FL4r���	P�!�d�5'�J��劰;�����K�7&V!���5�ms��]�C��|����Py��g~��r0��m^d��aϔ��y#ַ	�3�nU)`̦a�񀇣�y"�$CB�EPr���VW��[A��y
� 0�F�G;E�s	ѨT-�y"O���Q̒�1)
=ks"�5����"O�iP�M��F|h`��FL�7�!؂"Op�؆,�d�9�N�aH�}��"O�	9�mK?w��㔃	 aH,��"O��i�Ǒ��-�!\0��t"OF���O=9������R;(���5"O�+T"( �t�	�)��'��Yg"O����̓t4ftx'	��K��T��"OPt[��}`�YrAgN(_��x��"Oty�V��<�����*_�`��"OL�AG
��D���F!�Υ��"O�H�X��ӸhH"���-�!5!���Yx�q c�-&����H���V-�v�p&�A<����M��ybٿPv��H�哹dq�,a���9�y�P�k",�P��/d���&��y�в^�T���$��T?�����#�y�ID?T`~���g� 6k$�17&��y��U"�����5�� �Lޝ�yR�[�24Ș9FI�-�����㎛�y�Q�hl��M�$�0�r�f2�y���*S��k�Q���Ԫ�&۾�y�1��ȩQ��bBl���[�y�MV�k� X���B 6 ��U�W:�yR��{�2p�d��*�ܼ�$!	8�y��\��3%���S��E����+�y�kY4F!�q:MD�Z������6�y�L�%n�zȳ�D*��		�T��y��(Z�^�	�-U%AEz�� �D&�y��IV��$�$˶"��3����y �E��4���� g���
���yb�]�>���2fVl=�́��0�yRB +�x˱�)h��$�C��y��S7{������c�	ek�;�yHUTQ�p�.Z�)��E��y2�[�*�d��W-O}4@qe�y2fJmު���#��5G�bR�M��yb�0J���G�"*m�������y��ݯ(��P1�ߖ%:R 1@;�y���9��š�C��G1���Ѕ��yBfR����k]�*�(|ۧQ��y�o��Hcj�*b��(r���D.�y�����$�"�>I ��8�C�I�f=���'�u���U�JC�I'��!��29���o�x"\B�I���E�^j���H��G���0e>D��g��6&*6�`w�K��x�1�1D��˲ȯ5��]�g��C�� p3a5D�1�C=v��`	����2�D2D��#Ŀo�XQq�/E+0�D"¨1D�hڇ�H?1�����϶[��Q���0D����� S�𝢖 @�=,�:B�I'?�*�RC�$1讕S��ڙ[#�C�ɫS�9Ŏ!Y�PUB��^(#WdC�	>9B�Ӈa�0"��`/T�8C䉗;F�d1"j��.�M�2��2/@C�	.a:8`��ݘJ��P�0 �D�x��0?FH�K����  ���ū��]m�<�wfF|���� !�U�qg��j�<q�C!�-�re�}h��WL�<Y'�U$2I�(�V��GJTE�<�t�ƯC�n�5��P3vy���C�<م"�y�B��#G�j��y��Z}�<� ��5d�r�x0
�*i�L�@"ONmx3J_�mN�)���/����"O��"�n��E8xd{�0-��U#D"O�dN�D5�X�v�F�Ov����"OP�H�;c0݁�-�*a�O<�y���fy�̸%�C�YX���Z"�y�EƬw�����m,��Y oQ,�yB��
XY��6@����c=�yB�U�T"8�����< "�@�!�yOՋ���!!�A<���a��S��y�bH�;
���$7G�m��yR�WuD�	Üw>�i���y2�K�g�1`5�9XcX���ޫ�yrg�!	ۼT�2��IjF�I�C��y��@��$ZRh�42A���/=�y��[#�i�s/D%+ ���%L�y�o�))��|:7$@3&j�T�ŀ���y"�RJ�T�S��$�ZM���"�y2�C?R��i�ꏣ劑x���y'̉#����D*A�~;^=K��Z=�yBA 
ryα�fU�o�9������y���?VMc��
k����"ض�yb��T�����O,X-����$��Py�Dݤn|��pD X�+y���RU�<	���:��d�'�,Hc�e\�<��I�<E`���")�95�B�NS�<i�����
C٣���ц�W�<9�K���L��u'^%KJHr2K�T�<Y��X�Qyg�ܞ�L�	�Ex�<@�P�)���P)�<�y�&��<�%�
�9j� �"VL��Nq�<�a"Jj4��cI	�-�s��e�<afa�	7��y:eeI8~�s�dx�<���˖*�jt����OE�0�b^_�<��/�,Z"��S��{��P�g�Z�<@^�j�Hp �B�$t��N�K�<��eə-�BpJ4�&dfzЛ�"K�<I2U�v:�1���N��@�H�<���ֈc� �ae��7��P��k�<�d�E �0�;�4j��<!���c�<Y�^���54g(��c�<��fA��0���H�c(�:R��t�<��A^�x�
�{#)�
*I�]RC.�l�<�����!k���"CI�$��q�<��j��U����T�� LZ�X���l�<A����yl�Qs#�<A$UX���i�<��i�K�D]ȳ���=[�ݫ`�i�<Yg��;/���(P�
?M���3�(}�<�6o��R��#T�����C��]�<Q4k$^�ᓁ��F��؀INA�<a�Jعp&(q��^1v�N�`amd�<�5��)jߦ�0D���'�`� ��YZ�<�������,��ǔզ-��a�<�`���ɫgE̚QH }���^�<��%��=�SFeΏAB.�G�R�<am�>Rb��������i�n�D�<��^�>����v.TA�HA�<�$AZ�9�<��= _�yAF�}�<1u���:`�+�� ��1�S��z�<I����\��CK�P��,����x�<�ޔWRm����s6ڭI��?�y�B��B�f�A3n�	hۦ9��-�yT�S�~�b��bcb��1���y��l�\ rf�O�S��Hb��?�y
� ���$U�
%.���ڍ[.�Q�T"O�h���]!%t���	ҹ?8>�i�"OČ��0�EI0�Ч"O�`���CL���nV>0��p"O�@��˳&L�$[�Ku�P���"O�[��>5.J�"�H�O`¤/!�d�k`Rђ�!��͹�eQw!��ViV␒TI �|��Sc�X�!��G�@��KG.+2���� �!�䂅M��h�׌�6b>j�h�M=7�!�dG�)��yʥ��~�X���J�!�^�o/�ٳC"ֶ%�M�0���!��߷3�)��G�5"����i3(�!��7T��y6K�6�FpGf^�xn!�¿-޴����)�`<3�g�J�!�� 9lvD���lۼ�zЀ�0"�!��J6AJ&���
����E�#�!�ܓ���㍲;<+)�Ꝇ�Y���y���7S��E��t_^�ȓy�|�E��>]5ި) $T�V�ȓNFPAFO:a�Lɷd�fI6u��4��l�5	ʖ!��� ր%�ȓo1L8҆�,Go�7����y�
�'����P( �������.�(���'Pa9���o�~TI�$�3-R�h�' 5r�+��}���(��	�'�d���넥P��P/��ٔ���'# �J�[���+A�d<K�'%V�3�-F7}��-�&W�Q2q��'x4y�	�=��K���W/4�'y�,Z&Y�z���c[�WCJe	�'����v��Ÿ4�җM�U��"O~=҂�ݳG'R�A�&�&P7���r"O��)g�ۥg�	�V旺3)�a[�"O�A
q���9~PႆC��#7"Oty�d�Hg�M	q���Y)�"Ov�
gϓs@�3�5;(�a"O9��B]�� #5i\	�:�a�"O  �ˍb����ITX�"0�!"O`Iˁ"5-��]X]���@I�l�<�0 S�1u�|�7�чG��R�H a�<)G���߆�����-�P̲7hD�<�#I�x��s�"�[���j�A�<#g�d�D�R ���[��@��jD�<��a�0%O@M Q""|9bvnB�<A����{O��jƚ5��ip��S�<��2m�"�Q�X�|ji�2��M�<ǋ�m.�4�#O��E�%p�G�<�CXw&��#2/ˡ:���D�@�<�\伤# ���l�s"�z�<� �T�<��1d��|�Pc��s�<A4�7�A��B�*������f�<�DI�1^\��O)	��E2�Db�<)RK��6�Xi��Թ;ʄ��׋�S�<!�'ݺo�.��G���p3�pId�S�<!�$ߗ.�d����0g|]��`�M�<��"՝	���Jâ-�.y룏�R�<yPⅆ"mdL�!�ȧC���X���Z�<a�N�T��E#Sˋ&!�|�w�X�<Qw�ʇ���h��=b��
0b�[�<i?��]�gjҩM���	 �X�<���"jNqS`���<q1��{�<�ѡwS�P��sajTQv�x�<i%�=��I���.)XH�&�D~�<� ���ff~�TE�d��=�� J�"O�dZ��א9�} ���M{Rț@"ORT(��OR4dX��lΗ`o4���"O��q#o�9V�e���/$i�@+"O����gV����2�ͣ+7t��G"O���ݶU�l`G�:H��Kt"OV�bF�S�Rhb�����jd쫢"O�P��$��L� U���"O��YBԼv�f�6�0d!rT�A"O��H�/וe̌ B��&{JY��"O� ��ޮF������I1}�,��"O��+�f��`�HX�޶Z˾��"OȊS�3N$8�㬘:q�P|�"O��kEF�2ּ<�k�=���T"O1�c��J�d�u+EiqLdv"Olp�J����x��,[_x�
""O8O]%7GFd!6��! �,��"O���"��
G��F�h� �"OJ%�D(��f�&�H  P��"O�[�4	�D�X��IZ��}[�"Ov�Dɇe�����R�?� �[G"O�=�Q	$l�f�bF2����@"Op���C_�ՎL�e��}��H "Od��4��� �c�,�}b"Od�x�"׾�ֈ#
x���CB"OX̹d�!4e��H�#2I�6Q:!"O��[�]�X[��hF�ҪP����""O�+��)nV�c��2n
P���"O*e��f*N"���#��-��z�"O`MqF_�X����J�8њ,�A"O��T�J�P��:%J�-(�L�ҥ"O $��F�=w��I�FÒ�f�ZŃB"O~�`q��
��� �3gR0 &"Ol
�l�z�p��M�X#�*�*O�H �Ni�PR�
��qh	�'#��sg�3�2��pG[�<e2��'i�����ɲiL��
�NС6JF�3�'l����*�X���*���p
�'�v� Sb	4N4(�x�A1%%��'\�Dɰb�)�nu�YØ�	�'Ć[����,��*_1���{�'͸5��y��ժDf<
��
�'<�g�/�K�8z!@�a�f�<��C�H�9fCO2Q,.�3vDn�<�C�Q�t�B(X1=���9C�
l�<I�ҺH�s��V/N��I����R�<�Q��D���,nqw��I�<�I��W�:���)�~t��8抐l�<�2 O���!���H|�hM�$�_O�<���!n��-��ʀFj=H�IO�<A4j�6L+��
:t�8�e�J�<�gN߅I ��*�X q�`p '��L�<�!�Z`��A�Q"�|5`��F�<��)1+�T���3.V4\Xs*�~�<�	S;[�3o��\���x�<q��3��	��++0^�2-y�<y@F�;$ʤk�� ��X!T�Gw�<q��-S�
M!,���(��
h�<y��$H�	����jL�� 'e�<�ȏ6-�̠�f�Ҫp_8���`�<Q�*nb�q
��% #�t ���Q�<y2@ϙҼ�J�(;͠�6�_J�<A���>D��-�9_��b�}�<���*�8���c-8j�U��D�<� �9�J��(�K�h�J��q�"O��i�O�n�����Q	��q"O�=���.���EU����`"O<���n9�&)�*��U���+e"O�D)# �0+7BL3t'Ɯ`3�!a�"On����W�$�4�T��z�5�!"O�i�`%�aN����'���a"OJ�A�6]���3dĹ5�BA�"O��󈚡���q%��R��h�"O$E"�g�4�D�Dg�
IUnY!��'������G�w�.��3ϊv�(�B!8D���$�ݳ7"��`:qz|�ʔ,7D����OnYk��8�T���8D��(�(�w\�x곁��)���-2D�8���!BY�e��D��=I�1D�X҃��)`�$A�$�‵0��9D�ܹ�*Y�
�I�I ��n%�p�"D�,IW�� J�L��g�@�p�+D���bMeբb�$ɟ&��6h-D����e��D���m�.���j��-D���c �I�~L���Ůhf̐2�.D��*�O�?\��  6h����0D�)�B��gb6����ϕ���"k*D���I�3Z�0�c�F�?Kbz��j'D����ϙ0�L�	W�ȱ~ �=���#D�$C6mȍZ�8�ZT4|��?D�d������[�J)o��BE<D�d��M�S��0��A�6�Bp,9D���!�\%:vY+��s!�ݹ~�xC�%#�Z�q��	:����<=:C�ɢR���g+E�8 @�8e��f��B�1x�$a.IB89�b�xٞB�	]H���O�o�` �*N�5B6B��6���2ec��l�PD��ڱx��B��I,Lu��F;?8*�p�%�?�B��k�N��$g�=oiD6fѮ4VB�	��q�w�>'m��C!~�XB�	�:pT����F
Df��R��$RLB�I�&�|���R�|��W��&{�B䉛 3�x���_�M�T�a�	�\��B�ɥBT����52�8(�DS�|��B䉘VpP\�ӒAГ�U	"4�B��=Y�t�"�N-s��i���T�D�B��+:�<���A�&�^���-ѡ�d�9WQl@���$,&d�2&;M5�y�
-�lqK���'0�����Ԛ
�B䉽"�)�*f%H��g��X�nB�ɒ<�T4o�&C����g'04B��>\���A��:
 , B�0L�^C�Y98��Dm�@ۡ Ѯ&�C�ɪ2ҠܘU��9`�έb�̋^vC�	�TӚY)@�Kf{���w�L(@*B�I�N��̫t����!�4ΈD��D�O J#�6���p�d;L ,�Q�4D�|av(��`.Hxp�Ćq�4Ġ��?D�t�1/1r�(�I��ǺgCZ���>D�,Kt!BJX��*@B�e!�Y�c�<D�p�ři�`��� ����CS/;D���"R4CF ��w(Y�_�>��eH:D�|Ys�>B�`�"A�Y ���$4�(zA�{�EI�E_S��H�ek�B�<� �DN��n��J���3j�W�<���1k��1#��p�"H���J�<���V؀�(���s�`\�DSD�<� �A�C�܁R�41��&F�`��"Ov���b�-|�n�QRF�MV���"O|�)�h�	9W����O�N� �(�"O `HU�W�̢�0�DK�M��� �"O�1z�j�#w'�-�$iW�5�e"O②�������Ǥ@�xځ"O�AHtN\AlP�x��n�,�r"Oz1��cj%��R�l�Z�"O��"BeLw�����\	[ɘ�q�"O:1Ǯ@�>���A�D��θ "O�4�E�A�1��C�f�hHk4"Oȓ�ǒ�R�>�`"�70�J\��"O�Aqd@%n>��"A�J��ju"O�L�R��"<�v)!gO�j>`6"O�Ń��=5�p��@��4o\2d��"O81`DE��""l:UkESx�&"OHIR��6o�Ȇ������`"O0�ᣌ�d��5��X�����"Oޥ�6�^�Q0"��j��~�°"O�p ��X�W�L����|�`�k�"O`19�c��4
 ����7!��C�"O`���D�=Q�d�L�����"OAR3�K�j\��`C #\�yBa%W��h0��Ww�p�*�kD��y"�Őo;��i�.�5$hR	[�Џ�y��H�Nl�!
�+9�� K��y���4C'~���,	��z��[��yR�p�r�C)�du��ER>}I>�*	�'v|Aҷ%G:��'�G6bxH�1�'��m�b�J5Q"��g�F�`f�Lj�'�R@g�p �����ф)d��k
�'A^t�!����b���ux�Ű	�'[5@��
�]%Z��Q扲>�l���'>�t@��ݿX9ЄK!�66*�	�'��@�B���4`!B��T$-��t	�'� �10�T��#rl�(.�my�'�|u���)�>!���+�!�
�'�] F �,w��D��+��G�B��'��`�!�8��⇄�5P(���'�H�����?Q�0��i�>�p��'��ۆ�H�A��2lڞ݄���'kf���>]{�����B�~�zq`	�'�T����gKެ��T�r�t��'` qir�:-���d�q څY�';���1KƞlV�����1q��	�'����b�c��8��K<���'/T�2S����9@��۝.�� ��'�����[����3�\:"�>��'�p�p§�EMfpÍ���՚�'N�5j$N��صs-G��^���'���F�F9'�fȈdmƖN�Ij�'�T�P&�U�,�ZʓH��8�
�'#�E��d�N�s��D�R��
�'
��持G�(��FjH���̰
�'��HO[�|+��ƂD(P����	�'=<LhVb���@�Y��ֵ^�L�	�'� �īX8fr�*&d��[y�8�	�'�&�b$J#V�Q(�'Q�ZJh;�'�
����H�J��%JI�W9`h�
�'�P��f��g=�����C�=n�qc�'��X�S�ۧF# !%��5&��	�'~�\���*<s�9�T&�ZT4��']�0���?`�M���	(Ω	�'T��p
L.e8�x1a�P(|���� \��$�=pvH����$!����v"O.�+�$D�F��*�2,.5�q"O��80,�:��� H?<d�RE"O�!qL��uU���q�֜L�����"O��A�C�=��XQ^d���c�"O�݈���E�h��Y5z�ు"O<� EE�]���R�I)m�+�"O$��P
͑e�A��P�C�a��"O�PapĒ1.��;P� `U�,�"O$RTE�>�<�a�L�GC�\K�"O&����ar�D����	&(��(�"O���F@+2V�{l�v��C"O��!�I����D�K�C�ur%"O<	���$)q��R��V�|:f"OD0x7f��lx��DFЮl��ȹ"O�aYƢ�"?��,y�ߛ��p�v"Ob� ���3��Ya�CX��6$��"O��S��JhEء�Q�er�"O�l�3��S���Q ���Km��3""O
<2�"ʏV�`]����^-��"O�}�6M��$��D���nY�Q��"O�ݘ���S��9�5�YQdxѤ"O%0�i�c>d��
�
pc��pQ"O����I�,�|�U��U����"OLPR&�7�����" �%Z�"O��3-B&&������*-)"O�"�^@b�����*#�Ƞ�d"O��Sף�*�����/�2QZ6"O�0&�B���,	�DE.��`��"O�4B�J�8	/b�;�$KEņ$�"Or�'��%��<�DM�N��Q"O��(�Ň�f傦�L3W����"O�=p ��\6T�ô�?�Ԙ	�"O����$G n��C�A�+8����"O~��EG�"$Ȱ�K5c�ޘ��"O�,Cpa��o�:țV��nD��"O��S̉5r�T��Ƌ-}�;R"ORu�v�J�d���Fd�.}�1�"O��1ר�?K}X5;�$�>'`��"O��@ԈA-$NLI��I�ް�3"O)��Sd5$ ��E����i�D"O��:�V�7C0�)!�J�p]Â"O�*���E=0�xP��3� �y�"O��k�ǎM��DoV�R���h�"Oj�����b� �����ɠ"Ohݫ�j�-�� �.J�ge 4h�"O��8�*�(���:��8To��2"O����)^�
RF�ƍ*���"O�a��`�'J"|�K�a�T��@��"OzL#�eO�IE�t�� ��h5R0"Ozty�řEt$t �����a"O�}� Δ��B���.ب�����"O^h����JG�1���;�N��3"Or@
�O�<p�޵%˂A���P�"O�s�JR�U+�����i���"b"O^�����'\����J��@�"OB\�%�;��l�DU+��=H0"Oڵ�5��h��qd��{���E"O��i��&+�2��ƀ�"e�A	#"OP�K�aQ� }��@O_ 8�"O�쒁)��Ws��2f�Ur��`s"O:���H�	�dтn�2}�<H@"O�
���kp���B^�e�D��A"O�CᏛ'N��SF �da��"O� L IA�g�(�(!FZ������"O�L�!�>3(����eK�1�Ԁ�"O�Q�1�ʏE�ll�'ע7u昁�"O�R%�K�"������,a�Z "O�1#���
�
��QFߙRI���"O4�����-��@Hp��;�&�"OΤ aѢ:͊什�A� ��QX�"O搉��¡6��<s�,�p}*Ux�"O�U��L	�?j ���ڹ�`�6"O�� S�k��HKf�(a�肣"O�\���
T��(!�
T��� �b"O�I�wFJ�u%�@bA�(
��;�"O�m��h�7Ah���"��%G�
��q"O�]���Vo����FV f�2�Ѵ"O��Z��?u��x�bO�c��	��"O�M�fB��������&E���'��'��)�3}��O�jz�hE㏸�Փdf��y�y���*HV�lsS� �F���Q�'i�I���3(BY*c�E�U���`�'IR���G"o�Ʊ��-@ L����
�'=�|�ҍ�1Ch�YJ�Du�
�'X�`�r�(+�x��f!�5{|\��'�l�����-<#��ic��w#(d)-O�˓�0=!��DuC�ѫ����:�� Pe�]�<��	-Hy��� �R����P�<q� c�F�0��	:�ZP	�F�<)ѩW�ys�e�GME�7�� d�A�<���(��C�@��e��C���<�` �xR���[�i�X��d�V�<�e��>?�X��.I���E���V��p=y�'��H�F��w$��Ժ�a�4D�l�!�v�PQ��)�kf��6�1D�����Cl�Z�I�:Oj4ղ1;D��p )�("�t���W v�\"U�9D���S�H����	r����Om�<)P�E:vD��$��nj��υ]�<y`%ӲBhX�i��_S®6�N��?qJ>	/O1��R4j��F�4�B�k&LݛI~9�ȓPj4q� �χ> xA �Ř'�.ńȓ�F�j��ں3{�К�ƁP~ ؇�nU�t���Oޮ̢s��1ymF@�ȓBr��9VfΜ*��yé�~? $�ȓIN5"!��.��01�R�<$��ȓ�VLK���j݆��芏8��e�?�ӓ:��}1$*&ހ��GA.�$U��abL����7"�Q���^ԁ��Co�Dc�ùz��9��͇6X�D���8;�]X�K�8R�H.C0K���ȓi�A��G8��4j�H�5b���ȓL��8�@�mֈ�p�(M}�܇�*A^m�U"Y��t��1h��?��Q%���'�ax��q����'"�"~\8Y4O���y"�K�4�����A=,��]hԦ��y���Y�ɰw�N�����E�y�P.(�=#a�K::4�Ҕ�H��y�J.ZAn̈P��n�x�P�	��y��8$��y�e�U76���2�y��7z��S6�߱z%�xҗ���y��^H��Ew�*����/�yr�
,"4����EN6�b�d�3�y���'ZRyB�ǆ+�.U�&폏�yr��3�D�੍�#kƄ�"��3�yR���c�����)��S��y����E�,�Z���'��Ųa,O��y
� ls'��Eh6ؐ�Aԫ	����3"Od�9��E"`�0�Ѣ��D��"O�陖/�"LY����ϛ�V��ѵ"O4�ҧ�Bx�p�A��25w>��"O4�A�� Hn�P���d����*O�|�vυ(X3��S�n51�T��	�'� 9w�L6A��d�6N�(����'��qf�*B��L"6��$_���'�J�1ש��'���#���b`���'t�{�  `�r4�gʍ�n��x�'�Ĺ�
ٵoB����̂���'���2��Ҁ,6��#r E3�`��	�'U�P($c@�AJ�Ժ��U�{���'���JV�Ѝe#쬒 )YkpE
�'�6yy�D�N��+`�E�}q��
�'��}	Ө@�?*�"�` �� �
�'$@%z��V��X�s�'��iA
�'f�)�_���$��e�<&���	�'�0�F�[�%b�X�͎6�Bej�'�*M��L�^A��9��R $0,Б�'�qf�G���WC�.���'�(H�CŰ
6*��6OȆ}M�M�'��XBp�Z�&`j��2�&v�����'�$�q/�f!�¤A:_�,qk�'���#�[- -�6e �S TX��'d�i���ʔ;��s�DAԠ��',e�k� �S�l�j�:���'5���`D�/j�$Lː�Q�d���b�'��Q�M�6t��A{%��0^^��p�'.ZL���>"�N���~9�
�'��e�e�\U%X�:���8���'���S�W7 ,�ȲEV/34ݓ�'"t]j1V/8	���D)ո��1�'~z}0K&_� ���&���p�'�*���e��L�^�����k#��
�'�Fa1�KGz\t�Q�E�\�,UH
�'`` �*�\Z𪗒y����'���"*|��PbeP���y�C�'M��tatjةx�(q"@[;�y���O7B���!�&d�K���&�y�-��md��+��u���X �G��yB�<H)��'mh3ز��A��y���0�(x��/(=�h�t�T�y��D� Ȝ���ǁ�Cp�뀆H��y@$T�J=�q��/?��hC�̨�y�#� ��`q� '8�T�rW�U��y��_�� yEA��(��yxV��y�F:N��xs��/<���Fm��y�)�-~Ȯ\�Ba� "9�)�e_�y��O�(�`��+1�5Qi��y2ɘ��j9���
�8��QG��y�?�B9��̓.a\��P���y�;.ܱ���D
{ڤ1�I �yR�H/} ��B�ˋs�����,"�y��-����g�f} 'f��yb��h81`�ő��T�!��y�l�d�X�惇�X�j�x�@�yR
݅Ki6�s��
�I�^�Sь�y`�<4u����j!v1	$gT6�y�n[��&D��/.l��tT �*�yF�Q%@��qkbT�*�J�y�iA
j�(PYD�/H��s�S��y2Â�Q؞��h�}z��ڰ�y"�ۊ:N��� �f�6L
��y
� J�땪/v��t�Փ1=�6"OPx*�#�0OR��v�0V�0 "O�!%�	��N����� $�l:"O��Ҧ�w�~���g�/7���F"O�7L�$R�C�B|��""O�MW��.4ʕ�f�öGf�͉R"O�-`D�G:�����lZ�cT�"OFr�aȞqK��Ic��2Q"��2"Ofm���U�Wbf(�ǯ_-Q�a("O�m����mբUB�.ՙ0� pc"O>��ue˔u�½kw#,_�t"O��vO�dz�S��H� D�d"O]�ݥv2�%b� �6Ry�V"Ot١� 0��1�!k��X@�"OB�( ���(�0�D�(oۘ��W"OX�C��#��y�'��/gR��"O��Pq���%(�Pe���Z�U94"O,�B��)-^x0��ЖSl�]��"O�9�.����2�FO4w")��"O��ǔ,d1����� w6�%"O(x���1KHݐ�N��A|@�[�"O4�+��-:��g�V�7[:���"O��Ѓ��*��h`W������"O���3���
�h��,��w��-�a"OP�:BW�C���(BFǆ "te��"OĨa�eғ5|�����T�D��I"ON��'�E>Q}|��A�	j^�!�"Op,�QǛ4|�-
��݊Dn�T{�"O�A��9~&<̘�.=[�j13&"O�=	����Z�"1�V�N1ȶ"O�0sm��f��Y��߲x~V\"O��`�IG,&\ �Y$lJ�vtTHe"O���+�%\ a�L�:+Z��c"O�Tz����yX"�R�A�%�U(�"O4���Ƴ}�8єJ\>d��=2�"O|��E*E�	���bp�^���"Ol1���(8�Af�� �|��"O���F&v�Q�� >�\}85"ONE��Z)E���Į��t���"OjS�A_u�)��cU�`
ԣR"O��Ys�żN�"A[8HM�p�"O��cuh+Jb`)B�P�<�$��"O����`D�+����nϺls��*�"O�mbs��Y4�x��Y�'[�ۑ"Ox��#IΪb�2�c�!J���P"O�ث�/4$ӄc���#�JA3"O���&�?"\��7��v�t=�'"OV�`F�h����!�ء�.�D"OV\0p��	~e���� ��$3v"O>0�0�гV˺�#�"���D5��"O ����"%������b�Mb�"O���$�ɒLd����:<�5 �"O��33��2�qb�ʕ�E�<�Q�"OJ��$��qpx�RDQ�Z�9"$"O����DX�"@��It"O0�Cq�Q�$H�!T֒�d��y"cN*`�8�� >�4ȖL��yB�C�{3P�e���2������^��yڌm���@G%�"^ RC˘�!�_=o��iƪ��^� �RHZ�U�!����b�:���y>@Y�΅�!�DQ�����*uZ�]"�����!�d��fn�+�l��uK�	ZE��2!򤝘G�\4rC��RB�u/�zN!�� ���֗_Ʀ���D�e�RTx�"O�]�h�(l2�D��+ɸА�"OJ�%C�7����s�D,���"O]�%�%-ߘ*@�F��f %D�hӤ#�!z���k�oۄ%;+��!D����c�6I��NZ3d�x-[VB?D��dA�>i��#��+5���>D��$�
Rdj�ɣO�*�Q:Ï>D� �&nA)-�.X�F�J����Ջ D�P�Dӡj.�����Sﺠ*� D�q NW1%���CN�i3�X��B>D�(��)����Pr� �#Rr"�җ*>D���	�I΂#��F�,�ˢ�=D� @�h�԰a� ��*�$�qe<D�$BU�θn�le6*�;-�gJ7D��Ue�r�-��n�c5a��f)D�1K���4�ŠW+�ʕq��9D�4�w��J U�1U��M�j9D�(���� j��@N�b/l���A7D�P���
�`�!�"m�!�*7D���E-��Ś}��뢼���5D���ӰxPb��CVc�Ջ�*Ot���A_S��m�,Ԫ���"O��v
9@��`YsM�\�����"O��� ׄ�
�B&�/��љ�"O4j�o�(�hͫ"_3k�)��"O�a"����h��\7\0 )�"OX�;���	�$Äቸ	r@Z3"O�Z@T�l6��[�����&�ybӝ(�������q��Xw����yrf� R�M���	�b�ALB��y"��&���٤��_�:U饍�(�yR&���]Q�^G�ׯ�y�J�n���C�W(Q�+ˈ|&C�	�O��ѱ�_�PD��ǅ'[��B�I�8�*������9�<=z�"��F��B�I�m�r��"gY%$`Łň�B��B�ɰ_��Q�E�
 �zBI�%'�C�*f\��c�đZ��hj�DTm�B�	�a��eQ䓔r�мR�h�<E��C�	&C%���䂈2���T�
,��B�	^�ەȇ�`�,��
0j�B�I�nF���	;A��b'�7��B�I�BT�@Pjش�� G�ˡ�DŦ3e������-�Rص,�{H!�$ ��p���� ��Ȓ�6T7!�D

�`hV��8���j��I�!�d��L��u9U.O3G�*�oMj!�D,Ow�sU��:m�ݳ��Ãt,!��ݽh��dz"M�E���P�Z�!���2wf�<S�:Y2<U3bbڇ%!�d�"��QAգ� &>�����mH!��L��p�`3~9��	V�[0!�\;f�\�
���(ΐ�ըO�y�!�d�<j�xsHS(!��S�Z:I�!�d��m��yw=�脠b��!�̷xθi���ҎY��HA�H#!��Z�p5$�� �I�A�V�{#S4p)!�d	[*
�ǼFo��5n]J�!�d7�"-�7���3Qe;n�Z!��Z.���h�GџMY(	�#� -!�d�4Ť��3��Jt%1�j�!�Ĝ8mv�S��'@&�:� U�A!���5[��<;���'%d|2�TD�!�� r)S���?)IR��n�=ܰ���"O��G�L��t{��.4�P���"O���b�B7�DK�`��j����"O�IT�R�H��a�ک�F"OJU������ԉ����
Z&8Tڧ"Od��#�<_N��@ĈQ�&�!�	[�O�fc����#x���DE�'��8��'�\��g�8(�]��X�2��'�~8��ė=�3��S"G�������*�' ��Q�.	kv����H
I#xX�ȓ:��Y� �Qd�r�b
P�)���ढEE�Th��Ĉ>Ivt�ȓG��4
5� �la�8�8"#��=�
����ĀU9v��Ǯ۲%��p��M� 'W�V$zt�[�Z���BFq�<Q���$t�I���w�|�4�Pp�<YT��`�5���J�w�@��d��w�<AV�$kW�	�K�������Xw�<�0mF �*��S#ցITBG�Rv�<	4h�-SP*8ؔF�N�y�c�p���<R�[8����G
?�aI)�b�<QSH�=F];u��&y$
T��U���O�4y��:>^���\���.�y��ǔA��,R�`�2�R`ŗ,��d-�O��f�U>��l	S%J7|�i��'��	l����t��>�F��k_�"�lC�ɲ[�,,�h��t�p�ȃ�,b�<����:����2q4-��$'HJRh'��*�`B�I�v04-�P+��E�n��C�=,)Bb�$��p<Y��4aζ��֪��W�l\�'��x�'>�?QQ�b�4���P���|-�� �l>D�H+G��1��ʴ��e�$���E=LO���&�D�����S�z�� �釀~��^��H���K2䛂�Ez�$b�����	a�Oㄕ�Lk�>�!ꇳ>$Z��H<1
ߓs@$0*#���,�H�+J�\r�Yưi(�𤖝3�F�Cc�.��D+��K�Q���(�|�S宔�:�N!r���"`������2\O4@��+X�G{Eʑd��6��<�C�i�Fy���i��,"��D�p�\)��&[zJ�4P$�)��<�  W�un�rEŖ:.6,iS��b�<����%c�� �+_�{զ�<�	�]����%��f�����ǟ�n�����hO?��r&Z�T��dr*J�e���+D�p�bd�I|Yd�T�wv�H�K>?����=�7��&�8�h!��((�P�+w"^w�<��\	�Z����S�3㨸��v~��'���� c��QҲh�O*�	�'�X`⍄=딁��K@�|����'<"L�cLL2�P,����
L�Z	�'ݞ�K�!?���c��3:�5B�'O�H["��6:~!*�ć�,>q�ߴ�hO?7�W:+�D�3HA�~��ӬNW!��#:H����L8�b����]7\!�D�]�^M��oW
@���؇+B�%&� D�H#97�pS.�/v,��`O��yrF��t��x��+K��c"��y
�?�$ s���Q3����,��y�K_)Q���	�E%���˴J#�䓾0>a�#F.S��:�+��z������`�<ɓfːG޸�c�ؿk�ұ���Be�<��h�t�"� 7n~e6��"�F��E{"NT��M�iA�D�ivL�V/!���Ms�|8Ci�.L̹ ̛�,���hO>� ^����TSpR �q��;l���c�"O���s'ź^���� �O<\�Y�"O$-�u@F�y6���$�+�lHC0"On)�� �,[��RB"��c$�m�"O�9p#%Smfm�� ܱK!�=��O�=E�D��.6�vM�K��	9�MkP% ��y*�}��<�d,�/| �S�Æ�y��iό��=�����'��X��I�d
�"E5^�nT��"O`�a'��5�Z<�#��:.Q�e\��D{��I�;#�8E�5ĚO�Tju����!��
n|q�b�C�����FLÞk��'���$͘
vt�1��:d<�+��?��h��(�@����A�l)�ˠ&�jhKt"O�t�RD���h鐨�P���������E��ȁ��
�G1;@�q�"^�y2��(��S�"Ҕg�b��s�"��OT#J�Ȇ5�F�dK p�,�`�Br�<р͟K-4\��L��,�'"AC�<�!HT58��$��3Q>�Bl�{�'4ў�p����A���͠ ��6�E��H��Y��
ޒKCĭȰ�@�K����S����,h ң��k^��	���-Ğ���j3D�p+�KԹ�p)���j��� �;D�,��lX����Ȕ3f4(pZ`�7D���u`���P5������B#D�B���?y��K%�J�M2���'D�t��h�1A)�=���bPHS��$D�L
��<�t�6o�!f��=� #D�<�֫����s3��9{�Y���<D� �X��}h%"�*��GE�<0�O �=%>�yS
L���!�NO�,( f�9D� ����Q��#��ҊFe`H+��#D����ƫe���z�$��d���3*#D���B	�_�0��e*ɤd��P+�!D���'�K�)�����	�#^��3� D�8���8`2�D
=PZ�Y��&=D���` ֙oɜ��R�
1^�y�n:D�� %,�;T?Ν ͽY,y�V�5D�������,���A2Y41�w�1D�d��.�%��GA?�8��*D� 2�_�E\�3��^17=��:gh*D�i��Ĥ)�He�[/�|�-#D�л��W��B��!W�%��AR��,D�`ae�Z�->J ��aڇ�r���
*D�4����8��q&*�
�\E�7E)D�H0"��r?�� D�+Ft�t�3D�<AwjIr�+��@ʤ�$���hO��hm���]T|q*��D�kZq��"O�a(�� n�-鳡�E0��c�IG�'
�I�4h�+�G׀w\�1@c#��C�ɡ\��Ђ��K/�E�7M3��N<�/O��=ͧC�Y��bH�����j�t� 4�ȓVe�lt(
,44�sF������ȓ�����"\^�h����J�����I e���$KZ���'��U�(�6)��k�NB�ɰ4�$�4��%����?+�#=��|<��݆.�vj�O�X+R�ee�JN!�$�d}��Q ��F��g��r��O�=�� q��!TM
��DD6]�`#�"O||"��� fѰ�n��*t���+�S��y����V^�	�g i8�J��yO�@�xlj��*����iF�yr�͐
(�k4u�x�(�+�yRow<:Q�*_g�LDkB�@&�y
� ��)E�3|bL��C��++�\�Q"O̱�h��W|쵭/
�A@��y�<	�D* �Ta�P呠2  u�w}¬7�O2]krŜ�n;L�2gɣA�`1�U"OPq0҈��fh�3���"O&0ȕ!ܔ �A�)$g�,����4�S�S�����LI1tx�f��Q�,C�d;�0`��K���I�4��2M�=Q�V����O1)�ส�!ڂ3�h�ȓY�X�WD.V������rĥ�'�&�c%_!��C~�ԡ	�'�(I�2,L�@��1���
ļ�	�'u�s�O�%����W={͸a��'�x�!����(�H-"+7�t��'�t�Dkʨb�u�u�����
�'>�P��3g�<�����9^rpR
�'x���H��v�M@n�C4"��'(�9���iv(!���¡;P��c�'��!ĈPZ��O��~˶���'YʈX���}Uށ�w���s'��R�'zm�*�{m�� ��p���:�'�$�a �14�}��do��'`�Yc��ǲ!(��3��|� ���'�N�����9DQ^h6���hvb�'��-@�!��N�R<(�����'�4	@A�����A���<t�]��'���Z���8ږ�Z���s�tMh�'�m�B�TYE����тqll���'�%���ì#��tRB�5p�H�j�'X�@��d�+ ����%ѕdYAy�'�J�a��_+{�M���κ��'5 �;1gLX�4��cK�=𲱉�'�xyYӎ�:�F��V�k`-�
�'�n:EG�|��tb!,7�x
�'x�����<pN�9��C�{�f���' �R��Zp u24��:c=|y�'P|Ap�k�t=.��#��-�'(N����n?2�����
LVe��'�B-Ç��f�������00�'J:���
�}� 2T�`�'��]�Q�vD����	$�K�'誵ʗR��4���6HE��qN�({&n�Y苰"T�ӓQ����M�'6���[CKQs���N�^13'�@) ]{C�ݕ}}���Rf�)�K�-���z�*�_�.��g���QE	E�i8�O�����ȓl���؅Ԩ j�pG�q�1�ȓj�����L!ޔ�P�D�D���8�#��5l� �S�m��P��b&�}�T��&��xrc���p�P�ȓ|	�)��`R�F'2�qDȑ�[t���6�qoB& ���3	גfa���ȓk�j�B4E��[d�(��
�$�$��ȓ<�@Ph�`JS����-��D��d�\�zPdߗ����2�ϬM|1��W�Μ�����Sŀ)^ӢЅ�s�z<ra�2Me�%��g�Q�i���fśs �I9���C%(�HM��o9�4c�m��<���B��,y�u��DF����0<�`ѱ�������xM���=� �'Ö��vB��:k�,�2s��3Q�L�s�R
7��B�-'��Y�H�6B]� Qd$Q�C䉷��P;�C���M:��Q�Q��C�)� ��17��v�0Qrn���4"O��`�24�b����P�1"O��)�/:!ȁH��_�"�x��"On��r�U�(W��UH	d)>���"O�\4��N�P%���
66�k�"O��)��9P6����049�"OpI��ʑ�%ٔ}�F��*�Z8�f"O��O 7%��89��;F����"OJ��A���g�a�����h���w"O(T�A�IDl�oB� ֪���"O��#��_�V���I$.��]���K$"O��HG���&����P;�ȅy�"O��Q�C
�e&za��Fl��0�V"O�x����+��iA!��N >�a"OбC$�@*(vys��C����([��P�䋯4��1�On�ȓ� �r��:�p�i�g� �H��ȓ}��Xxf��V�,�QE�̂0fơ��\I�@h��meLhq7fO|���
B*�rf(Eز�A#DY&X���ȓDV���~U���g�8L����\��kȕ�p���7s�y�ȓhY�t���7E��kg�L�a����ȓg�PhB�N �&8����9��h��\�:�!J�*!F��J������CiKSh��mؾeuu��r}^)CrT�$��p����4=b���*���q��O�Ψ+F���ȓhb�H#�H<j��,�9��Y������7�͎;C�1�7�]WW��ȓ"py�^�A�e�T&P�z�`І�}:���"�;� ��V�ӪB\�ȓH�%��V�R�`=���%5d���!�)8�g҆;�� H٪N����?Q��>~@
�[���'YPL����n�as�@�z�!�B�|�xR��	q�,���F#q�" �w �&GZ�'�#}�'���2B��V(���D�BWvQ�'RfɢD�«5��ɰr�U�5�Ѐs%E�HB �bS��)X���5i��P!�F']P����j��z�@�64Uiရ�֛VÜ7O�X{�cȲH���B��y"��L�����=BN� I`�
���'U�8���o�b|���ӓ
dB�����38���j\W��C�IV`jA���N6�z3k%%=� �&ח|wN��,O����Y��i2(�
[��؁F��@qƥ�Ǭ*D��ru�ȋ;Ć�	�N
�1IN�{�X	Rb�'�Â>lOXb�,�D
�DBH�8�h(���'��C�"�f�CU�i0��k�Β� l��"$S7>��� �҇R��d�G��g��C��㑡z���rnP�ڸ'�zQ	Gȇ�=�*g�:
i��i��O&B����a�E/i�N���F��7*�'�J#}�'d�<��$Skd���א]��"K��Q"��>�&�)��	ՔQ�'����/���z,c�3U�́��j] ����AG��0>�����b�P��!�Ah�4tG@�ޟ8�JŨ���q���@P�y"I�l� \Z'�P�|*�,�n�ij�����dBQ�GV�<�H�'z��@�&@6��t�dc�
�Xe���ui2���H:^��`�g���yW��!ΐqxs�ۆp_d a3J*�y2�@�g��4�r�Z�q,����j\8	y8	&�-}�5*�B�O���f������E�A`��y��A�eO����\�N�{Ҥ\�����A�Ҧ���m٭X���`P$CQ��tc�oޫ[ܘ��N��@6���ݨ�P)��������%Ը��O��"���W?��B��(4��	��J�r��ӿ5>�p��8�zH���˟nLB�	�,$�mj4��y6x��冗4����ߥ@�fm���X^d`q�0.&��?�ϻ%Ҷ�E�ӥ8�����Y�<����9)B�	�,��Տ�8P�u  iY�"`X� p̓]����?1	"�%�-�
��q�P0e'xa���6f�E��I]p[&�%,��� �%k5,�#Z��"��~�T���'��)��nX����ڴ6ِؒ%(?V}8g�,�复�U�O5�h����s����ɩ����C�EP"O�=��O�,n-b�s���4g��i������������O쥉7	��w1L��'l]XL@��"O�0qO� d���fIQ"�5�=Obf�츧������]0t!���$���Zg"O����ϗW�TD�N�Y0t�0V��CQeӻ<bń�	<[݀���bQ,X�Y"��G�?�����Uy`��n�EČZ�=���jË�l�����''b��U�K<P�āiu���b�Z��գ9V�zV����O���O4):�ܓեL�,K�%��'����VEO��D���
;&'�A�۴Pդ��#���Pӧ���k4@���A��[|�\2�@z=�����Z~�T:�O��3'�ݱt�B����$v(�x�U��f�6Q��<�c�'�&��3`�j<���'�??�����y�g��=����a���ނ�ݏ]N�Q�E%8|(pC�Ыn�U酆�
��x�ƌL�X8��W�H������fd��4�%}�K ���1i	d'��'(��,��$��{
�3R'� AK�B�Ir
:��T��	$r���PI�7[�:� ǀ��O�d�Xb�����I2����.�s�L9HFQ�Jl��-�c<x
��'n��e��f6p�'�n���л7��ă�'I�>-*O��C�*�&��dƛE4��i2��1X����S��\R�,�t�+5��m��V5!�$FE4^��Շk���t �$UZ��$"Oʡ$�&u���c.��CA�9A#}�2�3}2�A�8��t�>E(ع�d�)\jx����34��@b@
�l�0 U��(�a�(& �HA���a}�ù4�dq�S�H,8-�1-÷��<�s ��K+65�mC7�y��� E�F���i�?<����f�lC�	D$�Eb���T9�d@�*m��1֕|�D��(h����ʢ� 5D�����-0x�h�(��-<-0�+U9�y��L�\�Nd�K�<��bN?|���JD��Pd��M(����L<Q$��.D3l����7(j��q��\xH<��Бy�ah�Ë���@GAR����%�0�p��9�p=�C�7E���5�̤D+�59FRW8����-0���V��,KXr� �M�J�֡k�+˵5�X��DeF9!!��ݢ1H�0H�p�I��φ��`������
�!leZaàY7#|�Mk�th+�'�7`A��q�\�<�'��!B@���)Ǫ?"���C��y	5rtU~�t��#A�	;Ľ�|�K>1��a��(�C'ӡB(r}�s	}<9 b�@"�=��H�n�L��^v���ƨ�!�
|8d���\/�d���{x��[�"?���mF�>��QKU�7�v��+�k5��D��M�;[�\�РnE�pZ6p#!l�+g`�ē�FْP��D�Y_�D��jZ��Ț�세c��I�T���%EW.a+�!e�[�+J�QC���ǱR��X�56�"���x!�$�2I�����˛n����)�Vmj��m�(���ٶ�!	���:e�~r��u�	c��*��;d�|��"��_Ê���ױ!�qs󠓶;���b�`T�Xqr҂��2*M�c�,pR����&,�y����k��h؃�؞{�1��N���O���ˏ�;����߁$�`�Ii{�Ç��P�ǎ�x&*pɒG!$�8 q��#2��iXAe��z.��(���ٕ- �K�O"BK�x���[�<��~��L�
ݪ�l�k�T)ȑa�J�<��$]��x���� 4:��hB�U���$|1ё�A�6��ܤ�z��c!�d4�Ȑ�X�,nNt�4g�!5�~B�ȌzĐ��R#R`|� CX�c=��y�F�^�"-u&�
3C�UA�^UjaybB��t3XAI��tF栣�H�,�O�bWc�g|Jhi7�N�(���r��@,wY��� ��odnDbw�/�la��9$�,�EH�r�ʬ��ߛ@F8 �G��>Qt��.r��*�=����dջAc^��~2�d�SKt���DK`b��EkUg�<Y��R'. =��͇ "⌘rfDG%$�(y����)�p"�)fGp\&?2�x�J���Z$�0��	WD��G���y"*�?Z���-��*��`AVH
��?-H ��m�(��pQF�'�$aKR ��o�ژzAG���T\��DQ	V� iC��T�YU�P�C?ym���a���y
� X)"P�c��zӠ[+��0�`"O�ٰA��T�X�HQ7<9#�"O��Sf�+�D����{�!@"O@�ѷ	U��ؤG�&Ci����"Oi������E�Z*q��"O�yB2B�WG"�;ҏ�#dP<��"OpRǫ ��)2��?�"�"O:���޹>36����ǳ|s����"OƠ�P��Jzpx�TfX��ٰ�"O�}���];B�q0b�rn(���"O���&�\�Q[���ЈC�"9%��"OB(4]nZ�BD��r� `�"O���Ğy�%1��A�<�B5"O�T1��#[*z-���}�mhg"O�Yu �?ID�7L٭qh0aS"O����喃.�tH�CkιP��*�"O�(s��4�ʴ9��x���g�J�<�T@j���em,jL@�#ɏD�<��R�K06tYBL�M�4嫢BX]�<�#)	�.mU�@�z	�]�VDF[�<a�#Y1:O4���&F�e��Hs4�T�<����va�ŪG�M
K%�ٕ@�N�<��]�ZTt���R ���0�C�<�cN��qz���_Zv���O�}�<q�A8TJN��\<a�Z`z%m�t�<Ѱ��[m����>&@�BFx�<YR�ٳs�QR4�&�"$���A�<�6��L]�M��+��;d�=����~�<��of���ўo��A-Z% L!�D_��N���N�C,ess- �!�D�+|�q� S��#D�Tl!򄌲 E 4��.{	>��pB}C!��j.Z�I#*� �.����3�!��X6v�h�)L�)��Y�d`�	U�!�D�6t��� م�G�6�!��ű0��;a&

����,�x�!�$]5l�ȕ�$�_�v T�᥋TLV!�H	8��Ӈ)��@��t� K,{S!�Ј4( �q��;ژ�X ��h�!�$ױy},McuK�9;���G���%�!��� t2��q��dϰ(�����-!��zB@�q�
y�1�P�#2.!��BNH<T/,W"4ӑFϯ�!�$�w��4���0M��q"�L�A!�DP` 40�	ÚO��p�@T�|�!��( ��p��%O�RL$�1�!��_�Q*͒��ԙn<ĳ�lXV�!�Dԕs�8��e�\�}r���"!֫q�!�Ě4\�X�ŭW+sP��"C��<!�H�@�r,2��lT�lQ?(!��ǭr-¸�6/�8s�}� �T)Q!��!o�U
��]�9t�ST�k\!򤛁".�bզ-xzq��N0A�!��7r�@���9l�v����k`!�Ą*^���*^��IR����a9!�D�(h����S>4�����f��v!�ď"9u���eϓ�{�a�7OΙiy!�ʉL���d&թEk��3a*x!��'}x�S��	S�m)V�L"k!��a��s@B�d�8(HӍ�0!!�D>9��l{1��{�d��˷e/!򤚣�������+ngv���(!�d�$�`!��_�������p!򄆞:��Aa�*K�a��T����)�!�� i@����bڎ�c���5W�X�"OJ�$�ӒB	\}�'B�*	�	!�"OJ|zǦE
/�9AbE�`:)��"Ob�e� ��$�獈�a�"OА0�^5p,�`c��12�V1r3"O���T����Pl�֮D*�"O�l���<�v����!_`"@�r"O��u��#i��U1�S&m[D�"O��p�m�Z�Er�[� 3����"O���sm�,�  L� ���"OXi�@I�i=n������)s�"O�
��n]���,ܜ;Mҭ�"O�0֨I�*qL��᫉ 0���R"O(��s��3kb�SVLޞs˞u�3"Oh�1e��1��ɴ.��x���c�"O����ŭ:,��LɉT3 P��"O�����Ԍ~pZp�'jBl4X��F"O��0�. -0n�H�`@Ts�\%��"O�d�%I�f����1QR�s�"Ol)P7�փۊĘaK�*��豀"O�� ���5��бl��G
P� T"O.%Ѧ��xu�j9p�6��"O\�X�/��5�М*�
U�����"O.���#Ú�c�H�<HT�9��"O��[����U��G	������"OPT�h2]\�5�R�� .��u�w"O�p�'�-cH�1e�>0��8�&"O���RI@�jst�P%���$��"O^�����q��Q�&\9�
��`"O��������hU���*=:�"O���%WrQ����?���R"OR�K8ER���Oj��E�B"ON �M��bapE�R8'�1�`"O9��&V1}��ʓ*_	̩��"Ox4��D{
�%�u��jmHe��"O�	A�G<V��ʄ`L4�\�1"O�)K�C3
�X��R�|�"OY�%��J�2�q%N�>r���Q��ޜU=�(�Fk:�a�"�t�#[���CJ�]u���ȓhE��PE��!mش败�8P������W�V(J��3��Y��
��V/n�d��-$ݸ�#��)D�4󖫉{D��6�t��q˥`F�o������8ju:(C�ƀ�b e
=o�X����t�N���	���Iy�l�W"XoZ�]���#�g�F}-�p
T?�C�	zSt��rAQ�S�Ȉ�c�νF�z�Й1�_ I1���ңMU�O�D@��#$.�Q�V��`�	�'7L|��;�-��_����C	��`��<qW�'�gy�L�)�r`�,���akǽ�y���sB�6�q�C!'U�8EסE3iO�шA'!lOL����� ���b��1(��F�' (�؄#��D�	ѿi�����k���ۀB�$"� ��reG�d���f���KV�H9���jp���'EZ!��O�(�� 3��Ӕ1 ���Ra���Цx��\1S�ވ|�'��"}�'޵�E�Tq� `쓗ꊿTL�hP�bVPM�Q�O�4�}���
�UO��ɏFSr40f���1����A�_\�`�ǂ`at 3��1�O��{VO�Fnx1���� �'�p	{D�"��@��[f/w�x����� 41��ѥdήh��ϐJ�V��T"Op`��JOQ!��z��]>1Rx	�FG�	��X!E"���;Sņ�&gd|���imޭ�\K+�8q��?[f�[��-D�l[�¬3`�Yx�he"�oR��Ń�z0��0bC[�?u���C�'{��G��1N�p�hQ��^ܑ�Y��8�mD�J~7�3z�I��F��m��q�3��+� ��Ǚ7a0t��'��",��p�C+o�;��Qq�`vJ����G/\��5U�pA�@����i��15Bˑ3��t����
�y
� �\�Ҏ7���`�&�$6GƉ���)� p!KΟLr#�\:یH����{�혅m@ ���YTޙC���%"7D����	�1vޝ���_&^AN���aY:���0�\�8�u�'��I�	2~Q��I�*��8��<�@�Cb^����+|O�`D�+���A�4=)��S�Ŀ
x@�AF�*_�8���<�H����'���Ԡ�?+u��ِ��O�H���d�)s�\��!�'S4Kf��t̓s��h�P�ȓA��5�����Rƙ#��΋1�q*ܓh�.�=E���!�����|������[ */�D�ȓg.�R��mͬ�a�gQ5�Z�ϓ wZ5���*�)�<�@�4��/��1r)�贅ȓ^ ��HF�9_+�e2h��;�<�'�x��ƭȡaz���2+�\Z� �gU|��'�%��>��^�II�Y{s���v��1$�x�H}0-��r4B㉧k״�pC/G�(��� Y�P�4"=��ӷnPD��a�7�S�}��$ۥlX�'����e���C�P�E�� �0a���b�5*�7M�0+� �q��S���)�禅�lԇA���,
�Mg���� 8\O�9��-S���̥]`���b^_7�y�S;|�������q�
�"��y��O:{��p牿�6�;���$՘'�2�� �%T[q��	y��)+v�%p�Lۜ7`�a)��%��Jǌ��xr�'.�I!�+�S�n���\�6piʂ�=}��W�*n��d�9*�v�'W�条U8	�$ϿP�
8C��K��B㉇x�YW�J�!�q��QPi�t�ǁ�7w�pN���I;n��q�v�<�s�������ɳG ȋ2NI�G�'��㇠Ɉ5DA�'��lpt�_�0��:g(��()�)O� fHܠ^FH��On
���U��&[��)s��'/��'��y�"�$*����~�։� ?;�)��Ҽ(6Hq�%�����K�b�^�<����Fs\혗 �-,�t���mQ�Y�d4A�>��A[�����ɮ�<9k��d*n��5 1xT�B�I�O�XDc����iBt%K�[\H۔��63��)zP�'�N��T�X�_�P��SbF�ClMH�_�Z��#��2An�:�Q!"�'4$�Y7j���ȓ6�H`t͘5����U-IV��<�u�D�}L^�`��I�9���{a�%
f�QI�(P�!�6Z����
eWF<�c�"\�L`�E�$���(��ɵ�൒��qǸ��KR/�$C�I%w*F$yu���)��d��U�yn�B�ɑ@��4�q�<NX������v|�B�I?n���e���d=�P���&<r�B�	&	 �haF&_(u3�r��4��B䉳'0|pz&k�ь�B�n�#jw�B�	f��p� ȫIYZɰ�۳s>jB�Il���w�-h8����,)�BB��;���p�!��q��Q�[rnB�I�u���R)I��| ��	R
@�?��
٤%w.b?�"$0 	��Ď�Id4�:T0�!�D�P��y��I-Wݢ1��R���-I`�r�VM�)ҧ�f�QO�^�yi���a��Ȅ�NBD�+�$Xl�i���F��T��XC �zc̋�W�-��*�Ԇ�W̓n��a��Q�h��`�eY�l^����	h9��'�ɔD2���L�5_!���L�Y��Ti3O6Q�E"��J����䆈0:H��qBRGz<"�)C�#�Q�� ��U�+0yX��'�6 	�F�3?4`	!�0b$���m����CVH<a&
�*F8ac�^;]��=�/s?!��[u���ꇯ�O�!#�&���!��D�<1@a��G�~ æ�Z �yҮ����&
� ���pjچ�?A��K8m��
b��	������RF&�%��Q�
7*4�a�Ad�H��/�O����/şS|�|�GY�PE�uA�Ж5ܔ�Bg�6�?D��E� �-,Ol��H[.ZnU���W�
Q�@ؐ�	?`����!$m2EȅUt�C�W�eS`h� f�`�p�r����Y���p��@��*�#Ohz �'�ڐ�-T��D��|�8��)���O��� �C�=�F��fhK" �b\��'�U�F��`�,|i�KNEFQ!��i& $8F/B�d���qD���'f��O� ��he�&n�tC0��1�]�P@�ȓ:p"ɥ@��<�HÁ�%�'���Q�����y�K�%,���r�n�$$]XĊ�p?	�"X.t����f���n^v��e1j��pc0D� ��S5�2��F�J�$�{��1D��ŭ��B�n A �H�.�8Ċp	/D�ȹ7!\$��a�gㆥ�����h9D��۠-L.y����	܄��3D��"�ڍ=DT4���� ��3�)$D��P$��9&ʝ�Fj�)jpn&D�ȁE+�e���EyH��#e�2D��"�
�5�vKƍ��GȰ����7D���PbI�^��|�s�;,`d/>D���t���J[r�@.Mf@	C:D���'��w�|�2��@�Q2��7 9D���FbBA� ��۔>� �2�d6D�r0� 	(D�{A�/o�8�:T�2D���0bI�b� 8���$��-Y1�/D����Ձ!�`js���y�D%��7D����b	# �iv����#P��yB߽o�A��h�8�c`��y2�Ͱ�v�����ݢ�F\��y���]�|��! Aj�t{��J��y��<C��B�-˟Dݘ`�휨�ybm&�P�Fʀ�1g��`�@�3�y���{�p0�q��!����W���y�J��β$C ��t��'�0�y�c��b����A�RT��CN�%�y«�7tn"��@�[6����Gȿ�y��7Q��#��h��vh˒�y��^��N��&�3�)�E�(�y�F�X�d]�A��k��3N� �y
�S�v�(�JW��Rd�f�Ѧ�y�*�x!���ɒ�L�8��.�yr+P!!��M��H=mLp���yr��(J�`�	W�2pڊU�f�2�y"i�&ߨ���(����= �@K	�yRX;��-0tmo�D���*L��y�(��gP$\���W�2��\��'ٞ�y*� �6��E��F햙��g?�yR�1��ᬚ96�X�sWA��y�D�U/.m�+�*����N4�yoR�n�Y�l�	EFO�e�X�R�' �����іI�������3
�'�ZD�R&�9{%�9���ׇznX���'�
Þ�J�x\)�.��{Z"�:�' ���܃&`��).E�t�L���'��I����/"D8qF9��5��'�,I�@%���F�*;s�4q�'$�ya��Q8F�0�5I�"ff`��"qT�4��V�����SB��	/A��y���*� ����U
N�:T|EFx����1i���x�f��Y]�5��H�H�!�䆲y�^��ɘH6�,��d��g/��%�S�O^`�se�@�b�@��1$d���'�0<�!uf�P��eD5C�>!��IÉ��9�5�*^������L&D�4��O�ӧ���L�閱(Q���.�-R1Ξ���A������ݻćٸ*��`EW8>=#Ճ��e���#�'Pv����O�)�\�"}���J�xI�˝�?�l��7ʂ/atܨ�O���v����?ӧ�)�)Y�lU%���=P\ �O�&s����<��߶�y2��m�OA���B�N6~e��0c�ߥp��`�Ĺ<�2���y��:�g?�����N��	�V(�;��(�O�t~�p���=�O�剱舘b�k�jEq��$;���ɩ�D7�3�)�'�a��h:.k2!8�X 2K0$�qkQ���뢖x�O���G�� �x{0C�xȄ� ���:omԉ�����0/�p}�f݈M@a��@���4��'Ǡ/ۜpp��!A�=�Z�x���Ó,�&>	֧�i�����֭lcJ$:Să�gy�듿~���3��E��'�{�Γ�>%S��"�3�'�>�����%	�t�h��9!�/^�J*�ĉBj������D��R��񢴂(����0|���ޡ3F$�
tɈ%;��lх�A-_j�2sd2?Ѳ+��0|��i1;Vi0�KA�q�4ܑb심K���CՆ�M�%.�;S�y�ç3�b] &cC�`N�u�'I�$f�h�2�	���M���;N�&͘�LP���Tl�F�Oܤu��OE�Y8�-K%�$3W�9��m�~�V`��c�2TC�E:cߓ�~��I�Sm,	p�P�\q��re�K��v��# �O�?�("K[�>��m���K�A��ݠ���"���Dכ��	V�,[�{%"��9�!��0� x{�Z,=B��3o��#�!�dM71���&Mn&u�G-�'|�!�$��q6�l�!g�2v<�L�1I�:�!��:����"P"4A�
S�O|!�p%�yG([4p����f�-_!�$M
-�������B�U
b�}��"O`]����a�L��3LE��W"O���L٤_�.m!�+A
[2� B�"O��A��n�.AYGJ�8dya��"Oȝ��ξl�<`:S�J�>i��cf"O쀨f�0D��`i���iM6��"O̥bC�M5��	e<5R"(T"O���&˂Pbia�x)*-�"O��3��=Tnd����Zj�Pkg"O �"��F�^ł�@�lK����"Oj�Q�$ѐw�(�8�"�iK���"O�ȵ/�4C3���a�'	=fh�"OlF�=N8�a��ю|~��"OZ�+q�Z�)�&,�2_d�9V"Ox�ÑÍ�j�Bc��4{:J�kF"O:刁ɘ;8,���*�8.Xd�g"Oѣ��^�fq�p��	^]HM��"OE��9�T��&�Z�unD �"O�KRB�$w�jh���ڴS�|��c"OZ�K����{�8�'�,%�ػ�"O��
��l!�s�עt8�p"OP����͉&��rR�Ξl� ��"ORHñ�߷JŨ�5Ér�&@�$"O�9�`Ӫ�ʁ�s���q1�"OԽ�f���L��QQ0�� Rč��"O�Q*�%pJ����� �BP"O@�j��M�r��i�.V�%v��"O��q�a  2�vĊ`�M�2SPm� "O��BCQ��8�V@]�&�*�г"O:���A�/��
wE�{vظ�"O�-8��[�[�����hR� a ]��"O6�Y�f��B�@�;BN�\�p�G"OPk����b��
��%�"O�چ�U�*�����&��=�R"O�Ȋ����^N�18u�V'M��`"O��K�oK����Z!c�'Z���"O����� O��bV�U�E"Od�r�x�����L�I��l�c"O�L�t�߀`�Āh���p� l�E"Od��Q��V&PCB�?��X�e"O�z��:I�l�C�J�UAV�zv"O�4��+I�;��ĥ��u>b43"O��1�O�{Ylu���U?`��"O��rI�h��Y��A�K7��:�"On��*����;K�	eSP\��"O��˞�jO��T)	"
;�ɂU"O ��d�"qrNH�C��-�H��e"O� `D���R�A)�A���Y�"OLMːN��qARɠ"� �9]耹�"O�l��	�7mRp�u�Y�GD�5��"OBE���6�����'8B��iv"O��K���G��Q�3HJ�C�%�S"ON�ò�>P����D'O'l��["O~�@�DI�E4�GC�@��4Y&"O~�D�Ρ:`Ѐ	��R��h��"OЁ�҄Yz�%���J�]C�$�G"O�� W��]0+��0+��b"O��z� ݫ%(��4�_4\N�B"O&	���J����C皭�!�"O�a��T�Vt�G��$�x��"O5[�h��65�u�� :T�
�"OP��pj6�\qA��ȸT���q"O�	�:�X�*V�F�U�����"O���#��(+g0���F���ģ"O�l2F�+H�(9" \?��t"O���vD-��Ts���)�d�C�"O6�!�@���FDg4���"Oz�#���υ�A��ɓ��'O!�Y�D�����H��H�s����!�H r����Ո1����c �;=�!���3\K��[�Eot��(�
"!��B��q2�Ot�l�3�eS�!�$�$/J.ͩ���/�N���%	!��.mL��b���E�Ā�4�!�[&]��I��o�;I�z���.ہ?�!��F� �gkC�laf���,ݰ�!򄂑o����'�F�d'�Q��K�*_k!�$_�w- �׫|�>�[�j	�^�!�U"Zw.����߭b��!:���&�!�d�)��P�B��e��L�]�!�$V�
+j�a�|4�D�'K�!��>F�r8��֟/o�%!s�S�p�!��(:&X�SE@%[���$Ι1�!�$' CԡgulN0���?L�!��Q"��"W'fQ�4q"JBK�!���������j9P��U�	�cs!�d�%�&h��#�o)p�
�B�6!�Z>J��uc���/=�ȫŌ��R1!��X�� ǥ	*��a�X0.!�ďM� yZ���Z-�SeѾ*!�D�GP��x��W�O�(Uy�dX�g�!�D��Q����j�=�Zz�i��	�!���$7~��'�/:�=K�E^6n�!��w8��GJ�L
m�EF��!�ڭh*R�#�ǊZ�P��
�!��*D4z��A�C+��c�\�Z�!�䖬_���6�ؾ`�nUAw��n!�$B��� Jve��w>R8��
;!�i�2���D��8'8�C��4!��Kg���P�Hq)���C�<�Pyr�-�{�.���x���]:�y���#,&��t�sj_)���'q(��&�^h���BfA.e�u��'��-�5JϚ��EЕ�a :���'y�,s&)
�r� ����ӌ���'*�#&Oȉb� �JӢ��D����'������P�l�0����N�Q!�'�tC����4#pBwy��z�'TƤ��"	�+~�����l}�ժ�'^��C2��U�)�ի�6?�e��'�h��iW+'&VyXT�F겸���� �`x����$-�=	��1�p"O�D���H��T���~b��""O@���ψ�S�% we��mk�|�"O��竑'���Z�@�
�$`�0"O��	p%ى�xzuC
�SS*���"O�(�V�L:xS�q5�A66�p"OD�ca���J���Eoɺ2RՓ$"O��e@V�g>`놏!nC>�a"O�j��Y�8��XNK*(8"��2"O�maem޽|vP@쎳'��D"Ob�"�A�`��z��֐�"O�E��:WJ1��	ݮA@"OH(�� A_����� ���3"O^!Ja<_�Ly��HH�l�(a�B"O~��gQ�漹�̗(�
���"OƔySj��m��:�	!�n��5"O 肂��g\A��^	�δ��"O �J�%��x{*RDS:	��'"O�E��c�	R��8k��Ƣ�4M(�"O�Aɷ�e5�5�u ·.���Z�"O��� �R?��Iwo�m�*��"O��H!�ݷ_�XK���
��5"Oz��4L�:J�D�C�M�<4&|0۴"O�Mcŋ�4cѾYG� (_�$iU"O0��J�Ex�� !L�x .剗"O.��v�K�>o>y��T�� ��"O�5D�5Y�b]qJGw�H��u"O��0���0DDK���e5~��"Of�C��  �&�kD�ʒ (���r"O6�R-�8j�d�;���r�"O�d겉�sJ4���R kK�\�"O�Ik��&?��ȳV��q���#"Od5Z�*C>J�����7E`P5�B"OPC�`q���BFA@���"O��K�N�_�,FS-U�"O� BQ�B�,ct��E��##"�!�"O��gB�2�2	����;#4���"O٣���,�4��FØ�v���{�'fX0PTmcY�}�Q� �g����'@����J�A�P��9-F
�ʓnHpV(�Wp�p&�94zԅȓw�Ղ3���h�Sp�X�(�t�ȓ	������}�ҹ��j��.�R �ȓ{z�Y+@���[�J
���W����ȓ��Ѹe��*AϚ)��o�A�� �ȓ~�a��:+�TE���L�0��X����'G�=1*�s�LW	#o(pa4D�x�7"�!Ҟ#�Δ�V� D���,D� rEH/`��]�5%Ѡt�mk#*D��!.-Ʃ��&�8�v\�p'&D��hש|�r$��,�o�yرe)D���e���/X*�4�I�l���c�%D���C+��Q3.!�6჏WA��(a�$D��R��ϰ)�,41B�α�p��$D����
�2Ek�Xi#l�7'H�L<D�@��pm�tS7��!;tY�A�4D�T���Ϡ_&�Q�
�%x�AhT�2D���Dd�
�=S`-J�D����3D�@)�"h=��%Up�4Bu�;D�(2�e2m��F&��5K�,D��J%�G�[��JFe�6�
}z�-*D��"�D�2�dY
Y�e�0a<D�t@ K�b��#�Hؓvx�z�<D�<����
�"�"�=FL���,-D�� 6��f��0���˲i׊��5"O�L��G�>zܪU��.Α#i0��U"O���A�,<��dR7q2�h�"O$���+K%>�[��g����@"O�$���Ġ-��QrA�f�J�x5"O�-x'ܺ,�PI��gD44yd���"O`)�LG�1�&�as��ah�U�2"Orm� ��8
~�0Zá��[�"OF�i���8$��IRAO(TP���"O"dĦ	�|��/�"<-��"O���e@�!>^�X-�"8�A"f"O�L� ��!eln�"Gl�k �X�#"O����g�3��`�u��=�*��P"O�!(����]P���T 9L�0�"O���cH>w+͌K)8��d@O�<A�   ��   K  �  w  �  <+  �6  A  0J  FS  �\  -i  �q  �w  [~  ��  �  *�  n�  ��  �  ;�  ��  ̶  �  a�  ��  ��  5�  	�  ��  ��  l�  8�  { �	 � Y � �% �+  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,͓�hO?�zP'���|��6E%V�ၖN'D��At��j��KC !sx��rh8D�@+�-�65b��@��B��`8D��S�;���!%�*��u���6򓑨�E�3#νw;@R$��Kv��U�'މ'<�m��.[&�9�BM�3�ڴ��'@�X1/�U��yk�H�+Y�8仈��?�S�T�ݚ���t��e/��� �(O��d��%۰��w��
K����d�ҢB�䛿�X⟢}�wi٪M,�Ad`�,M�<Xq��N�<I-�� �J��	f[p�Ё.D/����#�HOP��x0��0*��`�2准N��A�!8�O��hG��:�޽`�y�fC�<f���?��� �S��H�eB��B�2Q��!̟C��0E���3W\��"j^.ܤ�r�S���ĉ�t�f\:%m�8/���J�#��xb�Ob�>7M1?�cɓ�%��H��k�a���ç �\�<�2��*�L��(� �&�cg(^�<q��(4`�l\���`�e�Rx��Gx��
	N�`
a��j� ��5ㆳ��'^(�EyJ?�ІI͂X*q{ C�5,2@���'D�p���;a�h��A�&3d�ͩ3G2D����iZ27R�1��e�'����.D��(W�Ϩ��A!���(A4�IqE���`��	b}��K�kD��i��̠:�D���eգ�p=ٴ��C�:a�T�\*͂��D�CB����	�'��rF�U���j@	�[$�� �{��']�O�Oe�A��M�G�&��ӳ����'�ў�}� �0�FF'����k��W�L!��O~c�h�㉄�\���@��}2u#����k���'�a}Re�"~"��@K�J��A�W$bU����ɾ���m::MbGh �Szn�c�S�azR�D[�ux�%DYT zQBgeQ;aY!�d�>@��xt�[<0�a�I�u�����'����`F�;֢	*��E�ՂA,D���O\6���n��e��,rgJ?D��!#C��f\ک0��0JR�l��2$��SF�]"'�ZE��Y��)3cݨ�yↈ%O�BIzv�[J����ع�y�[�V�P1K�*B�%��5�&OO��y2m��p������]6 ����Eo��'+ўb>ّ0���%.E��)69MR��I6D����#�
T�^Mj��H��&���2D�p��(k�d�ree	�� 0� 3D�܈SB�#5s�#��G1sư�ٗ�2D�x,���Xf�p|�����I>����+�Yվ� 	��b�� oI*��B��+w��9�P.(�4��&p��b� E{J|:���J�i��!��/�r��W�<��]�V�L*SLU�.^-�T�S�<��E�E�̝
�B�/YY��()M�<�Ơ#q'~Pv˨V��H��
OH<���֑.�*ԀR�\U#&��S��%��{R��Y2�[g�R:�}j��	�>a{b�'(��R�k��'w[(�kÎ;) 2`���\1�cg] _�	@���3J/��G}�ŕj�O�� ���Y��A,^o�`k��d?O�4��O ,�ظO�"Z��h�u^��F{Zw5�O̔��"R�.((Ԩݭ4�93�"O�y�+�_���Z��ع"�!4T������9��xFz���7�����m� T����?��D֏&˖�G	ؐЮM�TNON�<qwo�;8T���l�O��ts��G�<a�y$��!U��#L��רM��y"�ށ)�J��K���W�Q��yBF��v��TIU)�1I_ ��!�3�?I	�'p����I�;��1�H^�d�L�+ÓJ���35�4#�SJ J(y�'O6D�8S�&O��d�$R� 	];��3?��)§8�����֫=eH��� Qf��|��&0&	#c�!j|�`��M��VV���hO�>�� &��A�D(%�"�i$"D��$�I�^�F����5�`<hu <D� �1���;�(��
Æjv���q�:D��	�j��o �H�� ��'`:4��l-D���@�7َ��4�ʒ��x�Nl�p��ɋ3����N�(W{� ��K"X���Dv�"o �A�D�[��F2F���[+yh<�c,A0 =���"���.��d�D�<Y�a%�!�ËYzպtZ7�Bx�<1��I<i�i�7@�����qx�|�'�\̀dW�E�����(�¸��'���C�]7`�r@�$�s��̓�'N�H�j�0
�fd)�kxTh��'u�s@M�4q�z���=n���'"LQh��/@�$�*ci	N y��'���)W��L�jS����W����D#�O,$��k�61��!����5@D0qr�'��D�E!�?`����%Ќ7.j�&#*D��Kr�&t��m�6!س�Z ���-D��F釋r-�XY����t�9t�%D�8R]jD�6h�@N� �	�$�0��)� 2����A ��)$)2+ �H�"O\3�ɕ�v��eqVH���;�"O���*I�N�,pڐHX�~� d�@"O���h@� w8��&�'���s�"O
	X�o�9�H����ڤ��'��Dy��)_�a�R��R��/&��a� ,,OТ<yu��2t�pie�J2+9�D�"�	X�<�O|(�G�T�]�<����LSGv�r��d`�<�>ͧO.�	�\qh-�G��~�@�a�6�j���'Ԝ��N6p���'�Ÿ}���{�\�4G{�'Y>\�ǫ�;�>p���6�@݇�#n�t��O;�A�$ь�6��=9�4�O�O��iQw�ό2���t.��4�I�'�����5Z�F�RD��4>!�PY��-O�9 !��i���)c�74a×��_���O�l�S#N��k ��`��S�	�t���'4R=�B�I	\�r8��j.Nl����",O4����@e1��k1��:-��82"O`��A��I�*$C�E=e�htqs"O��A��&a��CT%��88�F"OX��=W�f<If�ّ�0�Y��>I	�d� �[fM��(0���S�P�����py"�Y�`�{���2f�� �&/^��y� ݤ:��A#��S��<B�R��y�d��g�Bs`�}v�9�
�y�k  <�B�!�L��8[�%в�y��E�w{��@�	#qJ]�T-�-�y�Ǌ$�N���*���� D��<�yB�LTn�P�I�H�q��Bĳ�yb`p$Fu�B�G�;�<@����/�y��O�6�ԧǈ,���R�E2�y"�Q-ntt����Qu^�:B�Q��y�
�(мu�Q�БG��y�Q !�yn[6�& P�m�?��Y�����y�̿BL����[)g�P0�r!�'T4�����7C�=��&��F�A�
�'TH�pB�/��@"�l����<��gӲv�
|H��և[} uI�O�<YG鄊}���z��G\����T�<y&+3j�I�,��|0���q��f�<�a���jŇD�K;�l�3�]�<YQ
�|�f<!䪀~1���Ä@Z�<�&�G15��hD�ėo^�.'T���d��"u�44"��I2R_Π���,D�p���^��R&!�3%vR��)D�0�.R3n�>�x��C�&w�#t.(D��97�eZ,$���L��0�R*D����/�����c�%
�C.���:D� *�&�څ?.n�I2�Z�is�C�I�,1��8��9cf���p&�C��(C!6q��'���c�TC�IVڝ�BEpE�V6��#�"Ojt���mTh� b����!��"O<�;�"\�� `���r�~��"OF�3a?9+�	�P�+j�HM	�"O����$������J	D���"OD�5�i�"�1t�ܱ(nHt"Op�[����th���$�gꢄv"O>m����(�h��e��?b2tP�"O�� !$9p�3c8{�T4��"O�!�#��/b������
��}C""O���QA����12���2�"Ol�CkŅ �'+�!��A	3"O�1S���(7:Id ���>Y{�"O� �!bq�F�&(������j�ӥ"O~�y�۵*D���4n�
����"O�P`7�?_��\y@�E
��� "O��Qf���@����\24^8��"O(t�vnÖhPJ�b���$8 �8��'���'1��'6b�'o��'U��'��4)6o	(<@�R�o��Ix���'���'��'���'���'���'�h!�UA�(n ��r�g/�P��' �'*B�'3B�';��'a��'-&!��-��BIZ��� cwf!��'��'w��'Y��'�R�'jR�'��L)���d��LɁ���y���RQ�'�B�'J��'q2�'���'���'�H�r%M^1D���ځfÍ��%�S�'��'<�'i��'��'�2�'� ��'~� ���d	
�'���'��'��'g��'���'�v�s�\|ݒ|Y��]S�]�s�'���'���'N�'���'"�'�\c���2����ō�/@$HE���'��'�B�'���'@��'���'D��2ō�c������H���$�'���'Ur�'ub�'u��'���'��݊C�]�:>j��AI�� -�!�'2�'+��'e��'b�'���'��*� ~'$�b3b
)a�� %�' ��'8�'�R�'1R�'���'.�;���	q�M*�š5,��8��'��'b��'R�'�b*e�����O�-!��rP@���״&��H���Ry�'��)�3?�C�i���늣s�~��u��)gU�5`U�'���ʦQ�?��<)�)�@�9QM�/�x	��+���Ȓ��?a��Ǡ�M�O|擰��J?͹4��>R���E��:Di�B6����'��>i��ƚ=}bI)�`76�q���
�Msv.@a̓��O6=�6��t���CIHak�e��L�U�vh�O��$v� ֧�O����'�i��$�;,�ˑ�T\F)	��\W��Dc�B� �ȣ=�'�?��Ҝ*�4�0�ϒRu�my�N�<�*OH�OʸnZ
G�b����[�7K4C��Ɠ���	u@Q���I�4���<1�O��F�����A�"�j�	ӗ����<Z�4�+擼["�K�@��h^��B��3w��AQ�DTy"P���)��<�M�?�战$�<0Ѽ�4e��<y�i��؉�O(qn�S��|r�a�C-T����M�u�h�bR&��<9��?��j[>��ٴ��D~>��'qԎLs���;E�2E�7��P����O�A��1OX��|j�'�?����?���h
����(Ĳ4�h|��h�.{4��,O��oZ2h�t��	���	�?���zy�L.T�C���>]!�!N�f����?)����|����?�3"�q��Z��U��P�'�W=g�l@����f~�O��z�D��I�Mj�'��I�r�� ��%F��l�yL�7����d�禍���K��4X ��A�$1 �j�Wb#VCf9��8�MK�Rk�>Y��?a��0�!��^�hLk���g�D<�%h^��M��O�q�������>�	��H���7x���0��$&�J�c5O����Ov���O����O��?��BIҘq� �;���6sv$`��Nퟀ�����ڴxX<��O��6� �$�'u��P%ĄJ�4��/��B���O��$�O󉂅4 T7--?�;X�Fܡ�A'.f�#£ö \(}��mF��?!�B/��<���?q��?���,E�u;祙p��|��ڲdΔ0����	צ
OV�t���������ec��0���+J��V�p0�5w���	�����Or����)�	7�9��nےq0T� �I�_����ě�y���'����ӟ�ç�|ro̅ǀMj�)ʅ�h8�U] �"�'��'�ʟ�B��<16�i��
GL)Xn̩:�A��U�x�
f
J?p���'�d6m�ON˓�?� P���ɡ��{��ֽ6�r�bB�T�;��I��L��OO�Γ�?Y���~o��)T��򄂮0b�����#ZM2Z�`�۟'��	��y�� ֟�I��t��ß�ӡG�lD(�C.�-�&i��]1��ݴy[hu����?�����'�����;[�b�i� �&=��t26a��q�Z0�I��H&��SџT��/��dm��<�f�Rpn����L�.|R��A�<	�捍Hz��d�����?�P`�ݑ���� ���@��DkM$O�<lZEa�H������I�tĶ���-D,z���v� BP�?�6T�4�I���'�"�Z�q�GV<i�R���Gy��y�ܥH�����0�J~����O�0���>L}#r%Z�*�yX�T�5 �?����?Q��?H~�pj���?��J����6����OS|�,��j���P�r�'�|R�yG�(��-�U啉K��mz�)T;vr�'���'%F�J#�ir��Ozk���(vk�Y�\-R����0
�R�@j�alX��O>Q)O�?��(\�E͋>J�,e�u��S~r�|�H,����OF���Oz�?�+�`8�\�ڥ&��b�!t�[)��$�O���/��ɞ o�pY��C\�R��i�v�!%,d���x�8��'9>( L?O>(O���ڟTQb���\�RR��O����O����O�)�<���iu|l ��'=��qL&4ޞ؂�䔚eUx���'��6M;�I3��$�O����O$��#��4A�����B��������3,X6�;?��+�C���	�?��ɿ� r�*�A\'I�p0�I�c�X,�0O��D�O8���O��D�On��&���V(!yE`�f
(��$9�� �
�O>��ΦQsv�_y�,`�h�O���� ��U�ƁٴF�y�<б%+�D�OT���O��ڂ�nӐ�ǟ@1U��U�0a�ej��hЧ	,�R��'\P��I�nw���jy�O_���'��J̪zG����&�W�Ԁ{C�8(���'=�I��M{����?���?9)��k�T4�De�����3OJ�D�U}��'Қ|�OIr��M�H�Ҧ:D�A�(��8pش��Xy�[�Op��ԇ�?A�*�O��x&>O�cv�Bv���s�ܸT��8��O��D�O���O��OpY�%�<!6�i�4�b
�`�B*Ef�4����vE
�/����M+L>��4���͟��s�Q�?=T� )��^򽲃a��H�ɺ��o��<�N�&����'[�|����P���N6yf<��'�	���
#�ş��	ԟD�����ӭH����V�.̱C�y��
�4Z2��4���?���*���?�����wC�=��)�L���Ųq<�7�'�|�O���'��M�g�i��d�.�4�QB"D�"��=�7̟�t��dS?$Z�
�~���O\��|J��dY�^�k��R�Y�ԭ����?����?q,O��l�J~ȍ�	���I�,�c���	[���p�P�G�f�%���I�����ON��?��S'p*�uh�R�NqSSJ��P	�$�Or!��K�)v��Y���<��'j���$�
�?YH��F��`�m�2?�;�(�k�<�E
��2�ܭ���V�?рM��mP��?��i��"��'Tb.|Ө��]��rP`�a���c�l,��؟��	��p1`M���i�'�D�Yv'[@n��/��	I�ˑh���;wc����6���Hp�Q�̓C�(i�a�C ���'�\7�"6��Ob�D0���+،8�����{LX�"mJ[�Ԑ�O����O��O1�P�A�a�F�B����$<lV��K�8Vā9�(�<I�+@,><����"����dL�D \�x���(M�h��]�ma|�D}Ӻ$����O�Y�f�S�G]r�C�{.��+�O�qm�l�I���\����L�UG@N��a�����Y��{j�%lY~�g��?Gx��'��)���Vī-��,�#τ>r�b�I�,f�x�z��+�X�a�%H��9����1݂��̃0ZX)"tK��U��\�sDT�~�v	���#r^���Iv��d�S$T�k�[��P�@ΘDc�l�PLǁe�!A��Z"�\�u�����WMc�e�aCɒPK����NI��A`qNP R��Q� 
��%���ڤl�<U��	�X��s+��S���!�LUN��p�	��1��H�%��4��%Ad*ǰ0�������E&R��˔�������<�I�8_t�ɯO���?i�'��j�I��i���tL�BٴD�ݴ��Ca�x�H>���?y��k@O�(�lx�`��'�mAԫ�m���/B�x�O ˓�?�K>��2��Z"��jh"�Y�EO:4H���'�J��0�|��'�r�'{剃S�h���NV�u�!��d#(Q�D�F����<�����?mdӲɳ���1���!t���
e@�W��O����O���<���UX���4p��PQ�Q�}�|�S��ן;�V^���Iz��ʟ��	�|*�I�u����ƃT�dk���N�#H�R�ةOj���OZ���<)��#��̟��g�-�ޑ
C��U&���V�ҍ�M������?��=�p�����gz��2�%	�J���	���\�7m�O���<�wM�3IB����,�	�?i	R	�yo�� ����0�r��lƛ�ē�?9�1���Ex�֟�����	�c�$�&ɖ(8��ұi�剡0����4�?���?1���i���G#�2r�V(
��y��z�}�j���O�����O~�O��>U@�.WJ|A�E燥Sɤ��v�y�Hx0�J_撚�I��	�?��O�˓r�M��@k���p@��;Q��ɩV�if �{r�D$�S���P�ℹJ�R�P��xy��t!	��M���?���r�� ��T�̔'dr�O���C�4<�̪�#�P�d�s�i��'a���e&��O����O�-�3hZ�t:,��L
r�]�悙��I��%(��Z�O���?IL>�1;5Pe"C le��BS�í)��'τ9냖|��'�b�'�	6f��+��$qJ���N;���7�H�ē�?1���?�,O���?���� &�j����1���1�Ai�N�Ļ<!��?������G�%ͧ:���ȣɔ�(�Dȗ��xb��'���'�S����C���'�fx�X�M�JTJ���
}ڞqI�h�>	��?������#`(y$>� &˚�`�V��W	^�xo( 1�#E��M���?A(O0�D�|*����S	�.� ���NB�(���=D/6��O�˓�?��@@��	�Ob���k,��Hw
ݓ3�>n��h��01�'�"V��A�!�Ӻ��L$kE�d"v��R@�TB}��'p-�p�'��'��O��i��:�ϋ� �*�e-G�1��}�Z�D�<��hW^��ħ"� ��o��q��� ��|�2�o�U���*��6��O4�韶%��s��Y�Ƒ/#.�a�X"����F|Ӵ���O����O����9O��$P��YS���>ۂ����1kO��m����П�k3�I����|���~R"�mҪ�M��aǦ�C�j�8�M�����f8�s��������m�*a0��ۚ?���$Y�a�t\�޴�?�B�7I������'�Y�d0� ,� �MD�j�& VK"��3�i��	����'���'��V�в�������1�Z(%�*I<	��?!�����O��S�Y��d+%�ڎE�bܣ�>�F7m�O>ʓ�?Y�����O�H��ÿ?Y0֨�%�8p°�Y��EjZ�M����?Q�"�'k剄A�r6�D_ y҄[�t��hQ����U��'�BX�$��'!���O��苁9l�a����z�@5�bA�$ �6�%�Iȟ��'&��[M<)����v�
�H�BF�g�.�f���=��ҟ̔'�*@�S-;��O�������#,V��-% �⤻i5�	����`��\�s��X
%aP����H�t��/��47�<q!
��L�~���j����8�O��+�6��$Ԁ[��+��~����O����Oj��O��	f�ܴ>$4�BNN4���H�"_�xdo�4aw�=��Ɵ��Iɟ��Syʟ46JE�vX�D`���k߸hz㋚q}�ݤ�O1���M�<ĬЉЄ��/��j����̑զ5�	͟,���Iː٩�Oxʓ�?)�'EhmytU$/��4bB��0^L��c۴��g�T!�S�D�'��'Z3CE�/j�$�1G�0�1��`Ӫ�d]��-�'d��|�'eZc0�� �hCr���ũ`����O��X�?OF���O�$�O��D�<�1�B�x���d�(�Ra�fl�~�@��W�d�'j�\�`������I�]jt{��0nN���P�U��-	"�f������	ß��yR�T�s���%4u�BA"LC��3g�6ͣ<y������O*���O�� Q;O,h����7k:y���
W^��#�L{}B�'���'e�I�ڝY�������X��Y�R�B�׼�X�J�>^�Yo��'��'��	����Mcc#�]縸)G���{l��a������ßP�'e@鸑l�~����?i���z�h�F���B�a
�h��I��Z��I�D�ɾz�Db>�E*k��1c T)��N-,����ꦉ�'_�-c�"m�&�D�O"��柪�էu��G�{��1�fD�v�رF��M���?A����<���d$��K��!�����Ol�7-�(�N�o���\�I۟�ӗ���<��O�y�d툱@ %zLqɰAN㛶�J��y��'�	|���?�eiN4n�聕��/`m�}3Ń_jǛ��'��'ζ�b�>�-O^�䧟�E�x��]Xd� 
�8H%�wӤʓ�?��#�<�O/2�' �E�	&�2H �o�~�0��h�4Z�D7�O"�����R}�Y����{y���5�'�(T��(s�z�ص�����\�Ÿ'q�'�S� IQ�<�٢rOށ@Jʄ���I3��P۫O��?9.O��OZ�$� ��Lz4ʛ5�؝qSH?�Q�;O����OV�d�O��<ѴI�+2�B�<UH�9�Ж=Hh�`%���W�h�IBy�'��'a�|8�'r�������]��S�Ȗ
���
 $z�R�$�O����O������RT?-�	��p#5n�+t|p&�YR8*�޴�?9*Ox���M���d̓��iyr�!�hS�2������IA*�Bݴ�?����dٵ	8%>����?�!���a��50$��:��)�	�OZ���O�!����A�*�3��5�2�Z���P��T���'�<<	�z�.��O��OX��Bh�eK� <��C�Y�(8�nȟ���?�:<��G�Ib���OZ��j��f���D&-Ω�R�i���"�w�����O�������&�|���U�L�	����K.�X��&�W�	�}����t��^���?!FΫK��j�Kì&A�E��+@G���'���'�J)x��(��Od�$��x�N�e�H7��[�:��@Jl�ғO�a�4O��ş|�I៸�1��	(U� h2����N �!,�5�M�2�=Xxb�'y��|Zc �L����dI"G�ľk���Y�O�́q���OV���O�˓qꜹ��̕��<lȕl�����5�ԫϱO��'���O��
���1�SR8u�x��3������ ;O.��?9��?�,O�5;2*R�|ZV/�	?(b��D����N}�'y2�|�'x�n�yb�D*����NY�F
�Jծ��H��?����?�.O�u��H\A�S�0S�4H0��)��(�w�����A�4�?�M>)���?i��Y��?�H�����I�j�뤣�"D�="�Igӆ�D�OvʓJm�E�Ԕ��'���Ɖ�i:}�#E[�*��Q�%�>Q�rO��d�Ov�Ik�O��O>�� 8Qf�
G#ۮ3ل$yH
7BZv6�<�V�+)Q��d�~����R%��sԏ�:��E��'R  �jPJ"d���D�OJt� G�OF�O��>9;eo�;���ے�P��<�a��1�g���e���@�	�?UB�}o�'�8p�Ǜ&�HY����V6$D�~��"�<�ԟ`S�#V��W	��5�IӣK��Ms��?��]-he�@�d�O��BP@����s� {ǥ�G �7m#�ăy�B�'>���ȟ$�I5��B�A�${���n��v����4�?� ��d=�O��$;����h����v�@"��:�H��\�x:�	Mҟ��'
��'WW����Ĉ5k��T�!�@�  Q-W����N<���?�I>����?��ѭD=�d2��I.��x�o ��}C����O@�d�OʓS&�1P:�����ud�8G�\�4�[�xb�'��'�r�'`�d"��'vz�  �B�iB1*�a����;�p� QX���I��X�IHy� ^l��Riz A����š�L� -*2��~y���'��'���'�� h��'A�`B�A�ǠˌZcH|�+
kVl���IIyb��!&�����kLL������-�*� c�J�-�O���?�ZwN��fN͕b���ϛ�V���4��~F�l������O��iII~�I�/��`X��P�.�LT�@M�>��$�<q�����')	�TaR"Y�63�M	w%�`}0�lZ!l�Jt�	������4��sy�Z>��"�׋e@dH�Cl��yڊx�*�����ա��b>e�	�e�.���KJo���S��K�f���4�?���?��,$�����'Xr�W�v��TCv���H�ř�LJ���c��Ɗ$�I��p�	��������׫�&�4�j6b����"5\���O���?�M>	S� �슂�����
�R�'�؍��O�D�O���?�-;���K[=���e 3z������?�+O*��%��O(�I�^; E��a�]e�1���2�P6���"�Oj���O��$�<��U+󩙘\���.QB̩�΋l��	����Iy�I����=97�Q.U�I ����o�
d���i}B�'���'1�	�ERP�J|b��BC
9�D�QK�p����7?�v�'��'nb�	�$�L�9v��s�F��"��;�6��O��$�<�@l&��ϵ޴��e��p��Q[��CsF��Qhѻω'%��'�6�ˉ�T?�:�1j��e㖆@?d��h��t�X�:�T%+��ivN��?���~���*W3ąZ��l�!�Ei�A�7M�O���֑;��b?)a+R"��\�uo�V��8�Ӎ�8�4��		�_�~H��� +�*x�R(��d�W�T|Q ��Kw�Ѥ<�<1��U ��Ձ.D����IŚ_BJ`�BCA��ԫ�d�|��%�" <4�!�OR��0�wK��Kj�H�@F6��U��p�,�K1f�#����7NL�H��E�Fd�r�*�0�P�E6}\�
�d��`�shP�CHD�F��
_^�1df�ti(�@wEZ�*n�wo��`�DD����ʟ���֟��I��u��'s�3�"���S�$�'�'>7��q���~�"�0�ML:dP̫�eT���E~���H+6	k�6Mgrj��Y�6
D$�8qG\A�g�
���v�:|D�#=bOܰb��IK'������	M���	���E{�]�p,���}�,�rAŊ�^)!����hT��5=J�@��޵HD1O�\�'��I�Pf�l��4�?���h|2a� o�~�0�DK��H� ���?�wً�?y���t@�?aI>�7���w�Hś$=@"�" �J8�,Z��>V>0ٳEZ~����6��|+P��$Ri�|Zp��6DH��Ȍ�Ix�)#�'���1�Q�R5�p�u��	N̍p
�'kd7��D�t Q$3��yY��Ә*1O�}QS��x}B�'���T��I=C�4Z�F�>u->�R�ꑖ412��I����%dM�b�^�x�
!t���|�*�NܓF�Ą.��Q�恷��Ӛ>�Q ��XMx�6��L�Q?eP��� '@j�J�G�*Cv�h0&�2}�d���?A���h�>�$؛.G�=��=wk����
ν2k!�D�1g�y1Nՠs����B��ax�"4ғ�� ���|`��E�77���Q�S�|�	� )Hɰ���	����	֟�2>� H�x����.1�:�� �I�c_��;B�Z�q�c9�3�D�W�Ҵ��F7[0T��0:H{t	�����H�}|ZI!��L>!t�m((�J��Q�8�a_�?A�O�d+ ������b�"#�&��RE�_5;�B�'$�=�V���=4q��F� � ����'��D��D�leqU�N m���@�5W�A�g��)u����O���One���?a�����,�fyC(l��чE��|°����pV$$�!�!lO�ɺpa�"Zj����>D��q���(~�!ScJ-k�e��� 3d΁Qj5j��ѡ�߂���C��OB�d;ړ��'v���LC�c��|�3�+[���"�'�ٸ�*��?j�A˳�WN�.᪏yB%�>�/O�t�c�p}2�'�xb`r@b�A��zpT��'��#0��'��)֍E�~�sȲLi4l~ӄEb� ��a�"|����'T���pf�L�.墷@�'W囖�c�p�k �ޘ�C5b]��p<	P�A���xڴe��ɷV�t�5�� +aR�Vp�b�@��Gx�D9�h�$�hAѓ��s�(�8V�8���ߴ���%��b�bIӰ�S;6���Γ��D�2	�\T�'MbY>����Ɵ`q�Njj����X�x֙�bO����)�R�*p�ё
/����<�Og�&Rxĳ�m�z�N�z�C	���'�!C�
2}��gL��h��s3*	~R8�臭,�̵�a�>!�'ڟ8p�4�>��!T���*T�w���F�+T���S�? D-��AK�.�J�W�� d�'��#=!u�]�!��B�A4
8�iK����R���'@��'/���G��pI��'t��'�0�]1w�a� �D��P3LT(���<i��YMx�@�$ʐ�H��Є�Ȍ��a���7�r�x��$�/*���m�$&�/&��Y��Ę��L>!�e��i���o˥ ��@�J�`�<�Ӧ��B`�V!`> =P��`~r/=�S�O�|�Y���=ʬ{��ը����6+� `�'���'��~�i�����̧Ax��(M]�bYǩ�C�ܡ(T-�n<�0� 'k����p��>u� X�i��5�~����h��!`�숗O�pU3P�2jH��Q��ßT��I2?���;BM\�z(�T�C��90JB��H�3��GiR��e��"MjBb�XX�}��́/�6-�O4�$G�->cbO��F�����ſb����O�г��OH��d>	���O��OD"�i׶> �cqHΖ}�U ��'�$�!�b�@�	��	1�gAQ$�� տ�p<9f�Tޟt%��w E6V�$�,i�.�9u�{�<�6��+2A� .قZ�����M<	��iU�a�`��~䊩A��w@�yEvB6��O����|�*ސ�?�ІׅA���
ʅ@�d�'E�'�?�@�~�9�����Dj��@����3i�N�#��0}bj�O���H/A�3���U!N����+v�>aW�BݟP�<��T��B�p<r4�>.t�����H�<��jPs����2�߫j2]��KFA�d���E�W���B�к���GǇ�,�R0m�ԟ��Iҟ(���fԮH���t�����1f�:�@�욇\|)�gLD$���<ɕ�IZx�(���	,���x7����piaL:H0p����,�h��DSR�_�aZ��$�DY�a��L>����.���" �R��Rƣz�<�KS*!3e��dQ
����a�y~""6�S�O|`,�s���%�Z@+q�M�B��.�4�H\[��'���'�b��~�������q�F�9�隌���3kM��x��m@(�JY��ɣ5^���B�G�vB�EZ�1�'lG�`��X�2�'L�a���T�����~b4A U�?����?������O~�h١(�T�ڠ!�bˊ\��)�i(D�L*��1�L�!͝�� ��!�ɹ��$�<!���=z��I��\`�h��%���K�	ǅ^��$H�C^ϟ���.P`pl�	��t�'�0Uc� C�m�J�aF�5�&02Ǎ�<vdx�1C
7<�t�{��:O~p�A2�<<��HͬQ� �"dM��O|$x��������F��p<ɡ�Uʟ`��By"�B�=���nL�~�8�e�2�'k��'z�IT�ǋB�Ԕ+c�#D"��1�'��6-[7v0p����.6P��2CG��i�$�<�����)ߛ&�'bP>���,����W�p�y	�Ɔ�[7A�G�I��@��C���Id�S��Ob�B��$]�P ��e�1і>��`Zb���O=���RG�;2u���6��/�ajJ�da���ONc��?�c�h,�����hӎ0i�(D���B �1!鸄�Ȁ��Q�l)O�qFzB���`�L��ai_�o�h)�ɽbvj��?��v��X���X��?����?��Ӽ�Ҡ]&�IA�
?C��IÇj�'k��@ah��p^6�&P����u�|2�]�:���jU�%��)4O�U,�x�
_Śqlڗ�8Y����|��,$D����ñ&�~���LD�E����:��O�)�O��ș�S�k5��2dF(�ʽh�/D�������3p02嘇��K�H,?���)�-O��"�!ЇD� 0�:*��#0�G�iI@y�GD�O����O^��ǺK��?a�OVx�@ ��`�� �S?s��"" 
�xrĘ*d�x�sA��?���;�".v4�0�'c�x���}'���'$�	2�� �?���k��A$��72���фNE o�����l�E��]:��"@0 3�h�<A���P?	�R�o�џ��I���e����j<�S��:���Iҟh`�ɓ����	�|��i��'��� ��-z݃��R���Q��G9O0l����J�dT�x�D��&�i�OH���xr�ݒ�?�����d���E��'
�4!(���/��d�O���2�)�'ʂ9T`�uƍt���R���l5�� t�p���)>��q� HD,��,f2O,�TF�R��i1"�'��Ӓ%5L��I�.Si��
V�g�A8�*?����ޟ�B�Iݟ��<����Y!z=Q/�@v�1d���E��(�4�Gx��d �4x�� W� =[t������	<Bz��4�)�S)�\����_��P�mS�*&�B䉢oi�Tz��˫`=x R��/Ж��DT�'t����ٙK�Ġ�@dL 7p��J�a�>���?�5^����C��?!���?ͻ81JMaB���x"Cʼmf|a�p�P�8-�R,ğ!bz�� .����	���7eO� .~��4
]'Qd��#L��E?.�c�$ڧM��9��R�g�	V�!� ����U��������g~B,����C�'>v��(�1$��J�
��39�C䉘�diF�w�̽jS���\�Z�f���'��$L�&� �(���lx�Z�h��Lȏ>����O&���O$����?)����$삨������"
�a;�oƵ%=�T�Bb��*��Š��Hq�7m�0A@�
ƥZ\�����'���(T���Z�!G�D����?������?�����'H*<�2��.7G\��V�F+J��b�'�>x��A�����D�G�J�"���y�O�>-O�%iDI�p}��'R��z�CC�^���gH�=3ʶP��',M/|���'I�/Y�jҰ�wī[o�xql@�J�(���ͭ%C�u���4��I�����h�O�'e&L9��&>�T��>Z��p��=	KR������O����'��S����,@�v����a�j49V�9�Ij��  �S�
�M	K-;f~��'
7���ߴR �H����0F!M��S�DU͓���1|^N�o��P��f����*��%_�W�f�5,Z	)w�(�b�SQ�'�$�'!1O�3?���I�'� � �E]�H�%bQ~�DD��(O�cW`\�L[�t"�o��.�`zǞ>�d��x��p�S|��"	��8R싥FE�"��J��c�d�	Yx�����B*'i�р�Z--�	�8O��Fz��׊.����8f� ��þUj~7��O��$�O�y6�n]�d�O��D�O�NP�&�F�X���ٹ�-� ~r�c���U�6<O�����=%,��p���N�"��C�$�<U��y��H�)���1�/�K�y�K�.3B1Oi�S�����(E�(adK�1���͝�c�Թ�ȓ+�<���*L���Jg<���'g�"=E��m� l��iÆ7��`����b��;��(K�"�'���'�]�|���|��	����PHq�
x�6�,<�vUPPN�,��I���<A���<l`� ���#Ha񫆲/-�e�� \#��0����<�� �l��h3��9j�f@ukĲA��	2�M�p�i�O\�~�A��	PdxU���-|*m�@��`�<�f�װ v�� nI�b��TH�OF]��InyB!_�$86M�O��d\�i�T%���r�~D�uϋ&e�J�D�O(؛���O���x>9���Oj�O�4j�/w�<�Qpk�<��	���'�Ӌң�>7�P���l��i���C�"Z��p<y���\&�|��W-(����/S�����5D�$��-d��$�	�<��u���3��;ܴG�8�g��L44hֱ ��q�<9BO< ����'RS>eZ�����H0H�A�X�`�	�\NƤ��N�ǟ����-wV\��cJ�S��O|� ��&5j�����%eNʰ�>9��K
y|�O񟢬��$�M�ʁ�q$��a�t���>	����I۟ �Ix��W��0WF٬6x�q�֤Զ�(��<�����<�s
<e��:��3�QQ��L������g[Ή�Ѕ��*ЧP4�m��<�����rB�.~8����������_�5Y�� "�BX;K��2|���<�͕Ux���"ݠ��t�B ����y�h&A�t��۱LmP�A�MiЈ̱qI�<3�c�Бq��Oq��'ItS� ݃]�����ճ��'�!�� :���1r���|lb�OȄDz��i�#&���de��ޭ]،X"O�)�Bl!+��T8���#$FZa*�"OJ���	V�2-$�Y%��i(0�x!"O��1�@�?@���)�E�>O� l(6"O
��"�s�"=�����e��"O�h�S���1�ER%'B�=����C"O� .���E�%z)D��=G�<p�1"OZ�*�hW5r�P0�!5Y���"Of�7�I#.VZ�۠nߨxThȨt"OfH�q�����f#R>T"��"Oĭå�P$Q���c�|��z�"O��s�_�bKl)ؖ��c����"O �*�kѫ;�����N�	�
Q��"O�D�S�H4/dސ� CЛx�V	ؕ"O`�1R��c� �.WH���"O��'�]�XW:Xp��8�||	�"O�Y� b|8�N�<��pA�"O�����iD�AT� `�x��"O�,;�DA�������_p H"OfHr��a�2l�%-�q��@�"O�SCk@�C?<��v��F!�Ua�"O��Q�Y��}ےF0�ܚW"O���6'9MA�8a����A�Ы"Oar�kԂ2q�!`��ْ�Cq"O�����N��� ��EǾ���"Oޭ�WC�$�D+�w�r�i$"O�<	�>�x �OZ�y9f"O���qB�?/%x0���A�tl3�"O�4 ��T�v`=8�	�/|�� SP���� >�<��
\a?I��$]#B���&P$1�<�(�,[�iO�8�D�'���e\�Az�%����D�����逮���(�ɘ|�g$��]�L)h6�ӵ~�t�J#�J�~���DG�t������]�_�S�c�3� d���Q.Y�|���c1}�mC�'��d�~-0�@ל �С�6��X^�dt�P�yw<��>!Pj�=O��@��4Jbx˗����9O8�0AE�f;�h�Dݴ3:R!�v���LQ��ɮp�6PA3圮���I,I�L�r�n���@k t6DÖ,ڤn�X@�a�:A4q#��?�<��)	��˥�F�s�y����0s��ސ�l�8�)��^�1b�	I Q��h؍]������2��t���	��?�a�.�S�O8�q���SӾ�#�d*!뵉SQG��Db��06��P���g޽RÈ�a�*�#%��$YH���)}BB�S؞0�J�*�������\�f8Q�#�0�ا�+� DQ�6I(�*���a�O��'�,��F�W�Q8���%<@�2	ϓ?��P:���|�@�0���M*��D1|𐘑�횃w�0Hp��˄rJ��9	Y�8z��d8����+��Bd��d*��>�R/$"�e(���a������!	qqO�}�䏜:rM�@C7\e���'	~Ȩ��(�T��ͻj�� �� L,D!�;�i�12A�-�R"�<���@�ّC�"=�;#�[�w�v�ٖ�}&4�!�* ����dK0d�"<ѥg�=p=`b�P�?��QW�A�'aJ�!�C߬�:�x��Z�`����*On�hCgˮ�p˱��%�m2Go�<y�%���O��*�e�:|���͆.L�� �"T/%0���V
v�l���� !�B� U
��P�l�b��''��Y#�D��c N��gK�x#N<Y�'O���B�Ը{���"�`~�[���y�oI�P���&��X�`�|x�X��)B*ͻ+���Ce%O�=�pɁ�H�b$ҽ�f����GzZw�z����{��
sw�H�m� 9�9��Ej�'�����¾i���2A51����C��=�}����9���3 �40�����?�s�(��&�
K d��'߃Ƽ���X $K�v�'��<��o� 0�(��.�IbxM*e�ԥ,|�arH�=���� �Ǆ�J\���Q?f�����?�<���\�1�ˁ�F���ǂ��c�h㵨T�%�6ep5�o��OrMѶ���\xı���G1f0��*���ʁ�)�J-��|�B�`sC�@NY��?`���&�.v�h��$��?Y������
�ub*��-J�8q��(��$r�j��'�ֈ��r[��&�O*��; �A�i�c��c�h
�,��l�n��),�p���O��'�TKG��r��q���0/p���'�̑��	�h�| ��
.XTI���0.�z$��6�%�1E+!I*��J����k��N�Y�ıl��Q��)B1[]Cd���?I�SG�O))�O��IZ�HElt#$����'���k��B��xI����x�D���G�f�,�c �U�Kl�'�JѬ��(�W[h�tcS+6t��BC)1
}r��F��6�D{Ҋ?!��Ҝwh��kb� ����ʠ �� �O�p�3h����I�1���"NB#�(��Ŝ ��e �	�H�����ӫA3�aY�n�$m����� ��6����I�{���
6�&hY�$���� �Őy4� l�9� ��$WJ����V���j�}*��Q⇘*�����F�p Y���	�\��E���!�\���U}2'B?� +�*L��u���349�"<���ި)�0��'M�/WLr<�r�Ni��<�t�^-�쌘��O��p�'m��̓f:^�)we��\!�R���T1�tj�녺2����	ۓ�yW O�Ѫ"�IC�e�:*�0 ��-�j�`��I.V@��P �����a�B��uN�V��+����o~<erπ_�'g�akAf����OUB���bZe�q��B��7�rH�W!o�UQ$����S��'�`�z7��a�]x%L������}f���FE52P�����flD���t�����/�I*uHA��#"��o�9%�P,�A���hr������;�O�E�����'�
���	(������M�ִ���&/�IH�Cϧ$O��dی�$%_=ReK�u-$奟>��u��9�'؂��h��+<&�p3㋣N��,:�'�xM��>�tE+��h�8�B
=�@�H�JO�"����֮�$�"s	��@������ g��_�/ӊ	r����Z`�(!D��#�'ŷ)E��g���#ͧ�Z�Y�JH�"P{��ǅJ7�i�ơ̯a�(�$���
g��%�.U�5G�?Æ#�6 H�aW/�A��AU�m�p%���rl��4���(*�3��'�kE�G`C�(���Z�<yQ$����3`.�y�h�S(�lcM���g�@$���'?O��
�o*0���^uƘeJ�*h��mZ�D��#��l���@�i��I�\j�0ɐb��ݍ)�EJ�-U�{�|Aq%��
)�ܚ��J�4^R��㉌f��I8�w�$)B2J[�C�2ubN1}jxh�J�2�4�8�'���Q���o$(@6B�~�����d@!W� `gQ����ɍ+ўT�еm����K�f�p@p�BԡaE�]r!A@+*���bÒ>f'���Kw҄���cɨK���Ln�+z��jt� ��t(Y2q�x��B�
/;w��k��
��MK"��P�(\�a�5�4Yt�@Ҧ��_D�\�c���Y�'�N��i��G�t�#�L�#
����H�@��Áo�	��g�	�o�x��1)�ȽxB��j.� ��B��W�.�`�ԛ�-����~�Od^=#�aW�k�iP�5�4��+�:t��^�h��,M*��4��N8�Px�] �y��@9=�XatB�<�@�@0��Ck��ҁJi�0�!�d�|�2�ڟ��$C|�0^ce���� %:�8�w��q����%ғ&�Hqi�=�@��ژN�ZIh���f ꤘF'S%B#�@ "�D�.;��Q�V�	��uc�����S�4�hd�Fl\5H�$���mW8y*��Z�3k��A���<��u��
0�nI>Y�ܹ��1O�`��J�s��G̕�\_Nt��V��Ö��+��Pf�G�e�X���ޟ̲G�/e�h�BH��qz��Ò��?)qC��:��$�H�,M{ L�A'��� �q��X��M��m�i|h$�4�"}Zw� M�E/��U�1�ℎg�Ԍi�ň&h��qP+��8+N�z�AݸfތiP��>��O�[�wy�e����y�""�� �&���oN	:�'��Ls+ߞd S�O�X���$m�VL�3j�����]�@\NM��5�)E8�@�@?��bÄ3���$Ʊ]��كR��;hʄ��"u�b�q`�?,�� ��O�ʧǐ�CW.̀O���O��Y(�1x� y�f
�dO:��'F���U�tZ��GMb@�)f�qH�Ә)7�X"iũ4yN� �C}�X ��ӟ�H���+0�8�sP�%rИ<#a�~2�}�Ɗ�2���+�F�;����MS�N?�Ή�fo�OB��e�5e�P�S�}��nI��u��/Bڨcn��[H��A�O-m"GN�f`h��L_$�Մ�	�Tw`�i�C�X���H�ȷTZ�Kq־� t�eLͦ�r�Zk���>��?	�dB4hN$#w�ʼ-�=��c��$�V�P�f���"�������dfɺ�Ȁ3�I�uao����V�fȸ�ؠ3����?�2�I�>���a\�q�J��'�.O�����V(`j�YQJy�L��,�_kJ��B���]���ǹC���D I��7��k�0�:s�J**?�3����ɶ��:�ʤ`FC�u���j�Kń�"Y��;gI��`YV���|�'��m2�P;�"ؑ��;`NQB���ch ��e ��]��{��^1b�z���^p*Dƃ^	�D�+V�w�h1�qW��`=�Y�����w0�X�`F�J^Y�Ԫ���Q�
�'��Y��h�;H�V��'��I����]���I
:2��Ц��=p���'(�>������ 2&.�6��t� 'OFm2���'p�zGZ�%dL����^'�I����7��Dքx��(�q�$���@���'��A���-q��;d`ЬB��`��O��s�Ѐ������u�a��?D�� Ctَj���w�޾�z [@B��2�?'�{�#�-d��ӫ�7/?��J��E���'���H��g����F� x=Zx�.����Gm$��f��5T����ƾ	`$u����$�"�GOS���b�-w�9XR'�П�2q� O���p�a��e��	�S�'b���p'��,C���m��VJ�b`�t�pL#Pd�vyb�G�H�4uj�&S.���`�ܔQ|���''vm0�jJ�H��L�O4�����֨	u.O�P%��k�A�(��I�!J��$�0U��0%?�$����t� 1U���捱G� ���V�f�S�� ��~�\7*ď�>��A���T�ũ�|��e0�y�LX���?ႝw<��H���7\��\y��Q~��	�S���W����+�J˟t�z��dG]!TS�t̓F���	�4t�)�bZ��?����{a����|jeaؘ*���G��4��Q�4��qJ�HD|RMɹap�╎*v�اF=�?
� �L����-y��e��.V1;6$�2�ܔ8/rO�kb�gK��o�����(O���&�ͣ��5l��X12?O:���J�0X�R�5cs���"����yBjS�%zn��tÒ� �U��I�o$6X��V�
�,���I�`�@�P��/t�(h �)v;�B�*Uj扢Fr#<��yG�(I�
T`�!�6/d��i���0?�t˛E@H`䪗�K���z�N֗+�`\kQ,l�'Er���W<r#��5���=�MZ����)V����	v��e
��5������iE {ڜbS�M�@�^L�	�WW��c��
�F��4dH
}{P�'P�k$��4Vz��B��Z�4�4]C��d�����g�h躵j�(��	�+F�qc�*2��A�DP0z�^!�� -��u�j`!�F�&�6��g��Jv:9Y��6B�i@Dam��غ�
=��QFc�2��g���K) @�7�1\�T sf+B�x>����J	H�Ft���c4Ldr��9[!��Z+�5�Wiۆ:?��ui�?5.:( d�Y!��O6���g�k��s�IO
ة�-��w�d�K�Iݨ~���g���0<q��L
bV��ND�|3����ݛ7T�����,m@ř���K�<�'Z��7�?zx�Z1||���D�^��|�G�\�v��#��3`h�əNe�8x�O��'@�	�у �OtH���Ƌ���|\k�=c	lxW�F�jz��A6����c�'��	K�m:&�PT�V�Jp�� �Ǐ�Z&�aU5-ո�A��N�'h4�E2�N����E�� �b��fRrQ�ON��uc��@ZL���B	�XPl��N�3_���I��$�0y	����2,1&�ڲˍ*'>��^%X��$������På�f�xbj��R�&,�K�:4��S�xxE�`�(U*`��"7��H��B"(b �B�Bv)p�ыӈ'�[]��#U�^Az5����2m�%%��*��)���G�)z��`�J��նW�M�"��MC0m ��_�^� &�˔n2Q��[* �IDB܅E�YQ�	��P�d�OQ���&#����dC�y	H����O�OaR��P�X�a�r��n	#_8$�'p\F�5}�d�ҡl��+�n8���5��~&�2�j�9�L@�@ψ�;�2���%9$�� ��46��$r�O�  >�˧��Ha��'4>ak�K��PGh�S�gجu��Z�+!��x�J?�$�KJR�A��[;B
�-��M'�!�D	�j��t%�	^ܵ��	���'�ܴ�����P�#EB�)S�0I��"Ph?=�!�d�	�<��K�E�A�󡗞x�!�d��K�A0%)	]A�<iSCP�F�!��I(R?:q�+#���DR,2x!�_�|������x�F�fƝ.Ij!�D�12�yk��RB̼�3�:Q!�$�	}�`p�J�G��h!�@Ѿ+�!�D�*)v����@��\q'i!�!�DV�C�h��P�mS+̭C X���'��aC�T>$,��Q	!9'�E��'�
M�w�I2&k��;�E�77�Ԭy�'�D\K�ǅ�V �7�Z.z����'�ԉb"H��.�̐���=|����	�'d�H`�O�
].T��"s�VA��'c� !�
�U��̀������'��P�I7|�ܑ�"ꑑqrp4��'�ZMɁ�U:W��X e� 0r+�!��'���i�;1S�#�+�jM �	�'�h��
�m����P<T���	�'��`�eEE�g�����a�;K��(�'����c((5\l	v��J)�I��'�RTsƚ.w3h�0���?;�Az�'|�U�Cb[������g�10-P�H�'D0dcB낮m8*���^�SbJ-y�'���ЬĦ+�ew˕���'r��Jp �Ee��J�>
���#�'E�x��C�?��X!��"�|}��'�hD���
(8��X �S�*�V� 
�'	d�b�4c�x0%@��\�I��'�v�q0�L8O;�`5,�#�.$"�'�6��Oנj���C���C�=A�'��T`�N� خ���ݱ:���R��� �Tj��?=r�����BKT"O���WcߒP��U:T�\3	|3�"Oဵ͂a�ܙ���
���0F"O��RwCF1e������Km���"O�7O)M�L�r�P�@X|��"O(a�'! 6���bCc�5Pd�m"@"O�b�+�C���`b������"Ox	�#�:�@۷�1�z-��"Od=`u��	��q"C�֩MN��u"O���#=}B��q��6-j
{S"O�0����8��7V�1�`��"Ot�p�H-
֔i`�f¾bq:�	�"O\�a��q�A3� �WZ�,�4"O�ي���(8� �w�MSr��7"Ob��Tk�$Ynl�`�� g`����"Oδ���A�x���T��"O��1T._�H��y�ŃuO\�F"O(��̜#TJ�R7�HD���"O6��� 
5(n �s*	�\7&�c"Ol�����)*�t�q)�}���"O4�2v�i�<�5iO�ؠ��"OHВvל�ހ:�R�R{V틷"O���)��d�h�'#yf�@:2"O�đej�D}dq��&��"��("O�𪰩��$֎�q!��K��-�F"O.HBC��3&DaC��*vԀ���"O�,�^7C�N�3!AU����"O �X�m@�~@ֽ� ���C�, w"O�P�7�=gB7@�0vo�� ��'��*D�3r�>tC�Ğ���<Zu*.D�HY�G�%#>�|)����#q\m�F�-D�l�s�� =*� Y�,���
��,D�8�%��Znpi0̓�o����=D���P�S	yXDpw�ªJ$~L���:D�آ�Ĉ�C�V�1�( �&�)���6D��1u�E1e`��f�8G������<A�1�x0[��:���bKٶu��Q�ȓ99dPa���a%t��4���X��|F"�S(�t}�G�TB��L�&X�@zC�	�tG\��@,٤lK��'
��^�hC�I8v�P�0�a�5?E�18� �E����$;�u��ԉ��T�(�+�K
&H`R���R[��ݖ�IXĴkNQ���1���s�	AB����I���gO�u�t�/D���+Ħ� ��6Տi�:	K�I2�	n؞���AX
qz� 2ѦԮ
�2pJ3�O��	Y�*iKWj]%	�|̓W/'I��B�	�ٶ!Yb�ſpFl�yfj�s��B䉈o�|�(@ό)(6@����l�����>ٓ���'튄�G�@�Yx��@�{�<�qn���0E+G#F j����k�u�<Q�A�U����"�!^�q�Lyb�'�Z5��b�ug�,!dI�� �艠	�'�0-B�ӥ{�j�I�⎦`'7"O�iH��쑢5fZ�O�}h�"OPI�Da\-�,(�G[#B[4��"O:,+E�E8n����0�����x"�'�
���7������6Ś���y��UP�N!��ݗ/><���п�y��ŷ1�"��l��(�z��R�y��Z��r,�C�Y'^z�k�����'5ў�OO��"���S�$�ba���&x��'��� ʻI�4J����$(U��'���g�6�����ƣg��r'�)��<� �-R�-���y��@
>�^@82�'���'�eŁ�<�1H��%I I��'a���Ŏ�eE���ME�Q��ӈ��&�'
/^X[���#u��$H��F!f!~Y�ȓo�>��)]��+�H�y�����,�1���tR��oR�E��U��!7P�`���9
�=j����t����Y[�qr���"�4"6-�:k+���ȓOO�l��'�>!94�Q$��4tOFt��c�Z�Ђ-G8;�4�����P���0�@���Z-�@H&�ӽ �=��W亸Zѭ�a��((&		x[�ȓ@R��J$k�s������7!����eq�XI��1f�X�j�`Z���Մ�Id�u��<�ڐR��ּY�-�ȓxB�RmFTD� ͔�)ЖЇȓR��ר�W �hR5|i�u�ȓ#� ��FX	'|�(F�U�F�v��ȓ����x�����,S�h��ȓ6ؘ="P���Z����b�*��|�ȓ��E�q���|1V@CPI�>jxM�ȓss�t(��1a�P��Ap�}�ȓ
�̬
���'4\�ʃi~.0��Iy<Q"i�!n9np����>&�X2���z�<Id
Q"cC.0�};XE��p�<q�.�)#�}kQ�� �fy�e�h�'�a��C��=� )�@@���_ �y�ǲXz� �r�ϤY�
D$�'�p=��}2n�8vR��E���g�b4�����y� $_�l��#�I�ju �� ?�y�L1{D,J��U9��"h_$�y� 6��h�@/Ǆ+��h��Z��y��=^~��Պ��$d��hĂQ��yBH)U�]� ��+IDbA��b�5�yR�Čd��D�@PL���a����*�S�Ozf4C��+@�����U9pQ��'�uC!,U=T�:	��ǴT � ��'8���DjL�U��� : ���hO�a;"�ŲRx��!W�C�Z�=��"OF	�7��׬�9ũ� Ec7��a�O���	��ܛi�l9�T��$r.�ES
�'�zɕ 6z��1a�ꛧ4��1Y�'��9�"
PY�Q��TT�͡�'�Йs倀& ׸%�q�E? �y�'xdW�E� h 7;�A��'�80%�+�>� p'��tl��'�Z��d�K�Y�6p�WLZ��,�j�'�*DruI�>	�8@�OU����:�'���c�T�r��¾'�l�*�'Ò�A�LU�b1IPAH�"B1X�'�E��o]Z��Հ ��6qe�� �'������MD����e]"��t9�'�P#�G?��4c�D �v����'���K&E��I�ǅ��d-��'6����_0��S4K�l:
�'��m;0�"Y��r̚�Z`F��	�'�d!�W�	$%����>O��x@�'�T]
ȱ`p��X`��A.�)�'�zQ"U�[N=��G�N�h�De��'�vȊ$k�=G���׈H�8�\\i�'�r1��윁S�D�8��$����'e���N�9�V�ˇA���m���d-O�4@� �H�F؃퍽'����"O��+mW�x_V�׬�;�Ab�"O� Hyy�L+n	���̛6w�.�I�V���	Ǌ;���u%��P�CJ��.!���u����反��;p.�=!��*Eg���F��%P�t�E ��lb!�W;��8a�Y��I�.\O铜�>���IA���p����3R�l˵S�<��G�b�����!z"%��lL�<1�O�i�T�@���30�@�'iLE�<A��ә0
}��bL>s7J$
�.�zh<Q ��Jx�jɠ7k~ٺ�A�$H(|C��7�<�6�ȺQ�X�YD�o�C�	�7��@�Q������c�Q)F\�B�I�<1���U-�&9�vA�v���f��B�	�R=:3/�,��0*^�hQ�B�
T��-s��[$�޸Pg� z�B�&W��@�N*ꀁJ!kZ�V0B�=M�Q��7B�lу���n��1�ƓH֞�p��RS�`�^�VO�$��E��=��kW�������|�B��ȓ9�fPHu�Ɗ��	2G�-V�lЄȓf���D�U���( ��#���ȓ2��q2c�/��1�Q(ذ[m�l��M������$� ћ�%-=ĭ�ȓ������F������,��ؠ��q�Y�Fᆇq�E�	��d�ȓ(T�#aр_�~e�Ԭ��5!e��h6\���`Q3y� ��O�
0�*����}1�(,�|Us�"w
4��[j<|ۧ�J+j
<�3 �5;B�h�ȓO�j$�Sd�x� {+��ިD�ȓbќ9j����F�J�`J8k�  �ȓK�N�+�!��ع	�퉷2�J��i�"�c���z�t��H5/9(��ȓa?t�#(�(o@B��7�U�<� �ȓ}������͠z���̑A�P���!Rv��qg��x�YA�`v22=�ȓ5HVu�BJ�&���� ��l��QSha�ĚJL�2��]~�̄ȓ�2�� ӿ3��=��ǚ�y���v@��Ɗ�*�0��� )>7�i��s���bۣ�X���$'a�~T�ȓ:Xf�P%��*r$!�lǩz)ȝ�ȓEWLP���:;�:u�L˽3A=�ȓU��T{IܶImR��E��a(]�ȓ5�\��e�JBy�"�<H�D@��-�I�t��%��S!W�SO$ ��|���c0Y�"��@`���6U�")��/�\�fÌ�f�N% ���4����L'(�B i���Z!` -@�L�
y��_Q���0eT�]�>@�PCS�I~����:E-�%F�j\��{�A�FH��'�R�kELȏ��s�l��B� XA�'��� &�Ȯw�,0�k:3bQ�'E@$���y��elΦ7�8�{�'Wf��Q���/�n�c��09"8�'��(�t���o!�٨��͛#
8U��'�p]ҲKْIV����$J���'���ˆ��q���K���H�'�v��eEd@�mK �)vcB%��'��0 ˗,�Ht1g��0o����'\H1+N��l��Kf(R�h�b�[�'.Lç�I�T�j�:�,\N���'`��˶�F�voD�[��܎P'�C�'jn��# �5�U����LO�$���� �(�Q!ϴ4��c`��a~��ر"O�c'�ǭ� Y�g�B?q���1v"OT�
@�n2�E04�Z(n��"O6�Bg�(LeMKC�Sio��I"O��@VH#Xe�BꟂ"�q�'"Ob����aH,
�$#��Ac�"O.m���Q�<I|y��Vr�ҹA�"O��8ϑ1r��H���D�r+��[�"O�� �*l��r��g8��"OF�S��xa�Q�l�/f��4"O"y[��]�	�f\���۹%֬�W"O4Q��뒼PP�́�ϐ*Bt�E*O���A�D/]���2�``��'�����/�4�JS�X*x0�'��S��1f/�\j�A�3����'`lA�!m6*�����a�*���:�'�Ұ��N�*R�Z��I:�n�B�'����d�x|VS3B"���'V�p块lv�����${(�c�'kN�+�ɓ�A�:IJ�,l�P��'���b�Cظ 
�Ш�=\���'�x��%�W�E|�p��*�S�<��#	 ����	б��)��[R�<1�# �g-��h՘[�tQ�uo�Q�<i��ԴQ5�<�qEB�p�*s��E�<�BZ�J����A+��k�
a�$�Wf�<�D̦?����PmY�F8�w��K�<a�Ds����V��%G��1ɞa�<��
;N5�b�@ޙtP@��M�`�<�m��)�Ԉiw���U2���I
R�<y��ZMێ`�#�پ9b�|rӯWt�<v͎ <R��*���ʅ2��As�<	�B�>��(�k�,jؘw�p�<i�!Hh��\i &� Lv�h��XU�<�D�^5VFe�ʖ�+�r�b�J�<!a�	�}S.�� hE�m��B��A^�<ٖ#B͂�  	#=.Ʃ:PMX�<Y�jۇf��	#��*-_�a���S�<Y�jX?�bX4"E�(�/��ftB�ɿ}:�A�MU3q�*Pӊz�@B�IcƢ{��Z�f�f����ϗ;]B���X5#�a�A�f<��4�(B�ɈDo�=�i��`MN`y��<��C��)1����AhS�O�$i׏�eِB�	�30�(r1�Ud�P�[D��K�B�	Y�6d�`�@�訨��vQXB��,�:aBQk�<��|��J�]�DB䉩{-H��J�� �� ���-TPB��/:�.@)�ػq��	�FK?�.B��lɒ);����tE[s�^�D$B�ɦu�<P��1�^��BFʼZ��C�I:�*��8-+2�F�/u��C�I�y�Y8�`
P0Y9
5k��C�'��b'�Ȗ.�+. 3(� �'�	3,ƞR�ș�	�U<�e��'o��A@d�?���ʓj�T�\���'��M��: x\2G��P��'Eȼ�4"��5t�x S>s��r�'�Ldc��֩4K,`���d��X��'*؉Ȁ�D�4���'�^���	�''�聓��4�Й�T�H1>�S�'*�U��+�T���� Y�-�`���'θi1g?ntL��+ĝMe�<��'6��p�I3�LUD�&@����� ݓpG�\�(���i�"O�u[����t����.YBXq�"O�щ`jZ<'���rQ���@VVmZ�"OL��d�$ �}r�le_V|JS"O:�#`���y����+;�� u"On�cV����13�h:mx�"O�!#c��:��Dy��ѹ~�6&"O�a#/K��V�(�#Ě�#�"O>��R�ܦ4��Y�u'C�2Ӳ��"O�p�2l�<!=h��4' ɲE�"O���V�S�4��I���F0´q��"O��ĝ#��E�A�4GK��:"O�d�E7P"��pR��#N@�ْ�"Ỏ�7	G4Qj�M�� �rE��� "O��Zv+�;,��ز�ϖQ��"O��3 +�:K�X��PdK�m��"OԹw��$�T�5���6H�=�#"O6(���:��)��I�i�h5"O5h���߸��nTG
Iq4"O�e�r@[��6��QC��y�"O�,���ԴT�:Pn߳pU��'"OQ(ҜO���צǪ=��mR'"Ox)�D��q��5h��2"kh�""O��I��5�t�sD)MS$�r"O��rn,Ai�A�c;)6�P�"O�ڣ�C�z�F��F	�8����"Onp4IBs���fa�8���"O�����s�D��p�&�ʣ"Oh���7E�]��F�&[l��9a"O�+F*(�F�۠��+(����6"OPe;bn��?�*��%cժf��h��"O Lx�F$Zʐ	"ʍ	�d! "OF ����(�����a?U��$�"Ov���ҵH���#�ТF�>p�"O���II��AhJzD�E"O�\p�82��<3�@��7n��i"O������*Cۘ��&DP�9�"O8�$`I�r�8b.�:f�$��"O�{ƢԧS��!QqE�X��i	""O��J��˹�B� SE�y��L��"Oj�k!�QKA��!��[1����0"Oj��D�)5b�HH�,	l�*��b"O�Y+@OB.^E�}A���.�2��b*O�\Y1��0wI=�Eݹtk����+rP�*g�F<J�8��㏅8l9Z��ȓ��%�ɒE���㡎	7n��ȅ�Wf�(�bW~Z6���0
�R؄�.��L�R ��]��hB"Bo��E��|�E8t�&��d�sMAإ�ȓ�h1Ï�}1F���O^?ZX���*�>���	U#{N�R�&��Nt�ȓ^o�L��({3��C#�7`������� ��ʑN��93�$�
9^�͆ȓX�Jm��U�p�*I�`�W�Nihd�ȓ�qB���%�F�H�I������!!,]�6f��<�A�!I�c�|�ȓtW4��@N�Iǚ!���6�\��ȓ�YS[�}� @��p��;�Q����/2�-�5�C.�(�ȓ��I;%"�h��m@�*E��ȓr�tdX Ʌr�J|�_�lvlh�ȓzCF�1�$��qW�!��o�ui���<l�!Z��\p�n�/�dцȓq�|1`5�ݧ� �ʲI�,��l��S�? .4:��S�F.Hi��Ȱ9(�bp"O]p5�΍F��M���+QE)�"O��S@J
YhP�Po̯TA<(�P"O�81diκds�,���ţ "OP��͎F�0x��8q�Pn$D�|ġA ��l#6�:$x�@I%�;D�0� �8$>�`�m�gt�P�&B9D�h���B�q�bѱC �?���j'�"D�����mA��	P��=���²I#D�$��$�
F��!Ɩ�n:�܋1e?D�l�5�˷&��j4U*)�*1m<D�����
/rgz��pf� Sm~0Fk:D�x:Q
*A�����<H6g%D�8��j��,�JXQ ��q��%D��JT�÷R�b�#qb>�i�c+#D����::�Ha�NٗRծ�p�6D��k���*e�x��]�܁	��4D�L �χ6Ud���B��Sr�B�4D����ˌ�|>\��i�W=f1�8D��t�Q�G�4v*D�TL"i�;D�D`���������3��c0�:D�h�s��%�v�#j8�~%��);D�;q�
U�v1AV�[���y��:D�P�'+����b��Y3`2�Ь8D���e���4B����F)��
8D��r�h�3JX`���7����Ю6D�����9-�.�ui�R����1D�4��Κ	+�5p���n�@� �3D���%ö��ht��:`A(�"��/D��!���F�z�E$�/g,(p�R�+D���E�ҸB���r���&� D��J+D��ä�(N
��u�֎o�iX�&(D���p���w�^�Ci7X�0���8D����
M�XT�jcK�b�$��6D����!�c�D)�ÀG�J�Q*D���C�(�M��蚄-�Q�F�z�<Q��>)z� r$A��I�EOu�<�c�	g��H�R͡o���*�c\X�<�����ҋ����j�{�<�B�9f2���99���E�WR�<I6�m�0�Ñ#�j���X�<�a�ih�Q�	J�6�hG��x�<����>R�:4XEeˠi�r� I�s�<A�jB<:��]��mѱ�8u�@R{�<�d�ݜ�D�*E,fPH�gZzx�\�'ynb&��3!��9�t��p�8�'R��r�ٯt��{�C	d6̔��'>j���ꕤd+F��C��WZ���'���5$��;�`��Q�f$i�'�zܳ"*�H��#�,H�K[����'[0��t�Ϻv+ش�`�%BH^�#�'�P���-�w���AP�@�MO�]C�'�@hڕ��(���4�<j��9�ȓZT�:$�Y�=�(I�U���.��)��7 FhX�W�m:��h���%$����cXf�1�#�4�����(�<1��/�ԃb$�9:Z4�"�'�`���ȓ
�D����>��p2bۋ'D�q�ȓU�Fmp$����4�%��9ʈɆ�],��� ۗLH���`��Kd��ȓ`q��˔F��$��a۰�[}�X��ȓ^*cІ�1z��3ӥc���ȓVT�x�w�Q�%��6�F9Z��ޠd@J �-�~��P�ɚ�^���S�? �|��	��d	'��Ds��
Q"O�q�G�(;�\9�2���:��$"O:Y)�L��l�,��3�+�ܭr"O*���W^];0��	8x7"OT{F�
��9�C�q��$Z"O�}!NT�!o��P��ɝa5^A�"O���G&1���`��PDb��7"O�Q�ʗ!4�:�V�,| @�"O����u���#s%�%��"O� iAj)Hn���6eە>���g"O�)A�Ofp�y#D�1��2"OT|��jÿ$��u1���>��x�"O�5уl	C�`P�僇$;#���"Ov1p �ԈcטT w�A5`o�=�Q"O*�F��!H��e��u�e��"O��`$V96�j��e�H����"O��*g������S�e�\�Z4"O�Ԁ׍{��;`�\e鶩��"O�Ӓ
��f�֐�+A��zq�"O��ag��R�sce׀n�
��"O��wY?P��բ4.س?�@"�"OJ��s���轠4�V�m��aQ#"O�a��ϴ?�:� 
�N��g"O�!4�
$m	~\��<f���"O.�z�$�,���� �ObL���"O:
A��T
YC�.�-� P`"Ol��ƌ�\n����
z�����"Ouа(�59��c�bø~��0R�"O�	k�J��:�� ��%)�N8 W"O�y ��9|r�xBX�3��t#�"O � U�ͷc``�p�ǀ!K�5��"O�pR����4�$���NZ����"Od\���2GI���4C��<��""Oe`7�ZzV	�`��*K:���"O`�C��ғ��&��(A�]k"O2ȳ�ށl~� �K�73�y��"O&����tfLaY���!QD���Q"O8QP�Ꙓ;wp��nH:D�4Q�"O��B�Q�
��A��[G��"c"O
ثv�ca����{�<��dD�*�!�Ď.o�L	�MX.$��:�a�#�!�$�F��Q��D�b�L�Ғ�Á}!��u�~|��!���T̺w@�{�!�D��C<������%Y�d�)q���!�,�`��M$q�X�*u��O�!�Q+6th:A�_�-r��\�6-!�ׁ~�$�
�iHE����D49 !��@2%�aŤ =B�0-��|���'v���J��Z���f� ��'�2TiD�WF�p)3b�h�����'o� ���C(>���뗯,p*�[�'�4�	��|%Ҝ��/�?Rڴ��'�A��c�4@q�)3 žC���S�')�0إD�i��#^8etK	�'�n$2r�W�?#L��$)x�	�'8fQ#���,Q�-���κ ����'�V���+�8jR�������'���ņCy�P�DM���h��'�zؐ�À�+5��Yv�U�H�<�a�'� u� `�n@���G�Pm@�'T�(H���m�` kV*�(�|��'� X�7#��0k��ɠ�h��
�'B�[q�؀!��yt��zhx2	�'���c�HhF 8�*�(lߚ�@���  ��`e@�}�PDy�e�q�L��"O��@�*͉%�i*�!n���k"Ov����	�&B�9��h�7;���""O4�0�CE;���æ�ق��h�!"O��J�>$��g��-�>�+�"O��)2O�;6F�(��(Ѻ,�#"O<%Y�䓶-a(THɞ�l��V"O0$��Ô\���ذG�x*%"O����Z�j��}3Ђ�	f��%Yc"Op�ժҲ�`��Ql��:�rp"O��"���<R���WR	��"O ���n�[�ŀF�	5�	�5"O�Y2�H \��գ�@ �8E�"O~���	�"�ԑJ!�D���"O���2� gԔ���� ��su"O��CȌ\"���&O
=TJ��2"OĈK��Y�*=�r�D>tGh�i7"O�]��-�2n�L�4��-�8�"O\y(��	;<A�����w�b�Ps"OD��W!ARf����J�9[>�X��"On��#'Z�T@����dWq$R��&"OX́�%�?(�Ys�)G�	RN"D�H�F�U<�йWN߆=���[�i D��)���3W'��{3�+K�9���<D��H�oLhr@��%�}k�*��;D����(W���2U�Z	CF��ڑ�;D���cK�|��	��b�?u��͐�D/D�<s�ï��LKX��Zɡe�.D�с�_8~?"�����Z�v�1�h D�@Ҕ���/��hQ�����x��=D������0k�,b2g��CX�p(�N:D�P�*.*i!Dʑ"I���9D� ��W�c�0�yt̱O<<�t�,D�\�5��?\�t2C$�;2����*D�D#g�~,��Yg��pL���6!5D��` H�P�
��i�v�(P��0D�\��I)ܹ{�E�g�P�%�"D�pc�͋��"�����A�L,h�/ D� ��I�g���e��S�&���/>D���+�0Zx�b�,O4D�<a� N;D�t8�c�*:�F�z#��G�01y�.9D��(񌁠nu�� �סMc�TA��7D�<8����+1z�y��I�tQ���*D�lx$��v	�|rb'�~�����<D�$yWTIv�8F�8*�}�P.D��ȱ킲\����`��B���B�I�����S�Iy�HT%C��B�6|Dfm�m��p�
��Y�Qw�C�&[v��A��(g���K�npC�ɾ�dI@���/T��h��'*B䉃y��q�0����y��e�P$*B�IG)X�)�$�'Zѩ�,�%8C�E�����O�kXV!Je�PHB�I�q���眷)�ൌY.�
B�ɂg�=�ՊS2���Hw�)t:C�	�A!��0a/�
>���#�?y$�B�ɯL	|D�a��
w 1Tƚ���B�I~�� ��'D���,�9X�B�	V�v1��L�	{|� ɡ1[jC�I�P�x�CgMW�%eR��c�\�|B�9&��(�#�B<*g�x��ٌn�jB�	��"��֩�&͠=ba��<�HB�ɽi�ЎU�JQ2�Т��
B�I�]��8��۾���� ��C�)� �xz2ᅏ��0M-&���"O������"n��!�LQS3�Q8"OP���/!EN �B1L�"����"OBԸŇƬ~�ڂKN	)-���f"O*s���j"d���5	4��"O���'��:
`���W�Z�X�
�"O��*.�=_bz �W�,�)�!�$��l����T'FD�iᨚ5!�DE�g�j�ⵇZ-��#�<!�D����xg�Y����6��_!�1n&R9����\�|
��o�!��(D�K��@�@D`c��2�!�Ā-3��9�v���O�&XJc��YZ!��3�zl������|	���F!򄋤j<0���.��m�feC�86!����8`I�$ӝ#�`�H��_�
6!���k��iB������w��9!�!�ݑ9����jJ�n�6� 2Iݡ1P!��1`� �`�2�`��إW!�d��?�~-ʖd�j��V��EQ!��L�d� ��O�&x�&��?}B!�N7��UӦh�h��Pc(�B"Oh�	ݿ8������r��c"O^a)NB	&k̀C���<R��-:D"Of����*F��1fi��C7��z�"ON C��x�Jsf�+A �lK�"O��1Á�7�,I���C�J���3"O�!��
�"��V�Z�u�԰8�"O"t C@�[�Ny�g
�%V�h@Xg"Oԩ��Х:GZ-
���Y2�0`"O~���`� ���A��X*�N4��"O��k��C�F_�7'���"O�iHS�Zo��=",6sT�2�"Od ´�ٸ4����+�3 \р�"O���q	�k��pRQ@^�FȖPsv"O�Z1�ȶΰ�y�� ��f��d"O��;�"]�;���X-q^2q��"O8,�Ќ��;���a�J�85A"O�i� �!�|:3��^|��1R"O�8�*�!��X��N@vP��5"O|h�<����d@���2"O�z�AmCΐS��-)��j�"ONQIABھpKV #�W�u�q�"O�,�Q���.a΍�T.�[��yX"O`-�W�C�I.�X��ԷP�X}P"O�$�Cؔc[�(�aI�Fjy�r"O�,A��߳c�����T/_� �"O&4bwj��F �v��"�PU@�"O��2Ҡ
�uK
5�RF��-��b�"O&�)V���(�$���њ#��`D"Of��⎁#4j� )��!Ύ�$"O�A���̋z���UeP�V咹"O�A�4�����X��B53��I�%"O����ɝ9@~<����2���"O> ��o�Ml�8���V�|B�)�S��i	�'2\���TO�B䉂~*�YZ���Jh95NQ��C�1*Qı#AD��Z�,Щ��͉Q�B��JO{p�=^t�}R�̬z�B�I.K��"uO�wF�����K|�pB��:A��a2W�P�T��
G�ɼ�TB�ɽQQ~���A�d� ��D	w^:B�	"1B� �K��l�A�ψq�4B��8)?	Id�ցIk]x�(��nL4B�)� �uk׀�'_�b�KA<5k�ig"O$ i3��2�����FO$j@�"O&;r��*7c�}�q�&y����"O��S!%��\Z��aD@�n����"O�e�0��/-�T��elO> �J�qf"O�-9R��=P�])Pb�5r�(Y:W"O��A�Q�x⡪#7�T @"ORH��/��G�F�8`��=��X��"OL]�����>E1$�lT� �"O�h[�kْ,��HЭmQ��1"O�\�s��+S��p�u��m0"O`��#J�y��dG��-8�Z�P"O�O�)K��(���Q@v�e84"O
��抃! ��8aƬA�l�f!� "O���v��/��9a�h�Fr��P�"OTp�J.oH��J�I�"O�p�ȇ
�LddN>����"O��2d�v�*�5-ǝ �8c"O�Ua�R.J�����鏖芀�!"O�C�,ڸm��� ��@}ٶ��"O�T[Ѐ�]��u[塘�OԚ��"O��R���f�!���7����"O�ATnN0d��,1b����%h�"O�@�Q$MI0�SC��T"�!�"O$]��Ht��R��7@l+�"Ǒ���/^��ɢ��$�R\ip�|"�)�(oG2\���Y[��%k@Q67�nB�S/���I�+k����O
%�`B�I�ɉ�N�M��UJ�(fL~C�I0(<p�U��8�z���֤�|C��9�5	v-�c���1*�'�<C䉋]�:4�#gɍ0N���`jؔ@*�B�=P��%0��	5Tx<�Pm6�B�I�U i�F�	*�MP�(]~���?�����L�2�"��I��)�ER���[�"O�%���G8@
��[����"Oڥ���O��Tq��+^�"O(0��4<`�#'F	Sl��"O�����j�qD[1)mr��"Oġ�R	B�� ��BL?N�4��"O8��r�S��IQaҰ�|dp�'q��J�
K5QA�G LG�f�)G�'D���sn�U���B�\M$0�!D��aM��RZv�b���
gRı8��>D��i`�� �FI��,Z b��ec��/D� PU�B*M
�Ќ���@w/D�H鱡M9��� # �����*O�4Ia��l�.q�2
�-_��;5"O�ab'�s���2��;zдz7"O����8el �Hp�O�Qj�9ڥ"O�M���\@ĕ����XW��"OT��Eb��C�~����
)�n�r�'C:��`�K"�ؓ��'DCRL*�'�z)�J!�t�b�f�@�D��'|
}���ʶ����[�7���0�'=j�M�!P� 5$�ߣ4�|Tb�'��\��o=Q\ �R��"`?����'(���lO7z�z(��L�Vİ�
�'�^�{���0-��'�A�#�D��'��(��,�![):�#�.( �R��
�'g�Ms�&фK���P ��i
�'Ü�sO�.B�"�NY/f�0�'RX,U:Q�u ��c��H�@�Ow�<�����H�
��e*KAdH=a�ǉo�<� h�k�LW�"/�,�"��O���"O���W�05��wa��d���"O8��i�B����.v�(+3"O~��Qc�G|H���M�,���"O�xa�ҝ6��`�V�,֠x�5"O0�
2�?*D`��#��1�$}�P"OpXöƘ�>L�ؑ�-]�A=�,��"O����s
����E6�a�"OpH�� I�T*}Ӓ�˨,��"OB��!�YH9[��\��<r��*D�Ta�kI
A!�!�ٚ��MY�k)D��QED��o�=�q�V$6@H	I�*=D�(yu��4/s�ar�T=+@TT���-D�$�A�w��4��Jm�L���?D�TC��T ��|6lLGx�(��:D��ч�B?b@��8�dگl�͈T 8D��
��ٺe)XH�H�'n D������s+ ��3���=W|eh�9D��3�9K��ɂ�E �h�r���l#D��2�	�TÊh�`d�vzFU�U�4D��0%�JY�fg_��8ez2�2D��1���
��Qⱦ�md&��j1D� d�9%���!/P(3E�{�0D����22��ݣĩ Ә��H"D�d�w��nnƩQB�P!t��BQ/"D�\
��Zm�����ۀa�&�Z��?D����3���Д瘷��шfC?D�*QH ~(�hC��j�vrG�!D�X@f)C�N�*p�ѯ�41�Fdx7�>D���q4EP��3i�HIzx�S�9D�xB�x�HУǏ�\l�+��*D� 0+E��Ѕ��	ϩ0Z2�<D� za�JQ��c�͘3C�䠒o&D�$������T��dX�TZ�((
!�$�<)��������u�x���(~�!��� R������Qf����G0T�!�D�.~o���!�jH�cQ��K�!��%(��s0��)2*� ��Bl_!�>X�]k��7(���S���!�H?.Fd�A���r��tc�3m!��$]8��Bu�ɔ B�a���4�!�$@�<ڈh���{�Q�Wi[.,�!�K	t�r8jv�@�R��h
�0tl!�$�w�X\���Z5�4�2�HG,|!��T-� �/ɝ1�����D<zs!�Ą�yw�71��xѲ`F�^q!��k��RsKZ6��ib�O��_V!�dK����p�D\���X�"A!��Ȫ��2vިW8X�5�!*!��̱b�L�p#Pq\n��vKQ	hB!���E���ƩX^�YJ�J�!�ĉ�\�P�hUH�:d�����߰�!��5?�}k�o�;X�I�j��C�!�̡+ǂy醣��}��(R�� ��!�ƃ<N�k�&"&��u���%�!�dY�y0�1.ǈH�� �ć,�!��$g��XprZP8pʆ̾L�!�$�8
�q��/	д%KB@�!��M2H�}1�-Ǡ)˅��1Sh!�$K�n���J�=^�H��3Q!�d��sM�}���s��P�KK$ k!��Uڎ`��N�: _��x��21�!�d4r1� ����(NrD�E�É_?!�ԮM%D�'N�t�p�y��Ͻ�!�� 8�Z&'R�8�*�Gߨ�
w"O&���^]{��b��]�nYA4"O����@&������ƥ95p���"O���	��%������Κ/��"O��pl��I�:��w�2n��j�"O�Y���ns�9s�ɹ�|݈�"O�a�їtxr<�Íӿ]��9
�"O��[e��>"ܪ4��*>�N �$"O���%Յo��Ը��Q0/��y��"O����`�,;�$2 ]����"O�9+�"nr>iSD�/[`Ƹ�"OYڔK�� ��xqt�Ԟ>'�Ms"Odh����-:����Q쌢4�4��$"Ofe��듫|��U�r�(��"O�T��U6e�����X�W�I��"Ol8k������J�3�>�:�"O���d��e�p�l?����5"O28 R!f����zQ /�u�<���	W���w��,��]�үF�<�u�D�H��R"��j�A�<�T�x�����Ѝd�|�2��}�<��"��Uda.Wt��+�O�<Y�e�9w����GѼCsl��o�I�<�GED�D������ <���,�D�<����)$��p��`�T�q�i�<�d^�8U�t�%
8r;"���WOy"�'��U[â�;m�$��V�C�,Q�	�'��Cv`�^���"ր13��Y	�'&`�Ja���1��Ų��Xc�%�	�'�Eq��)��U�T�3W,@l#�'�IZfo�5O�.���ץe:~�+�'�����¯{� �lY,n�'^0x��� ��J��5a����'ﲬ[�K:'.��tʀ�+Q8q�
�'�P�W,�^#��Y�E� )�q��'m���B.��rx�)
*�+7(A��;�:a8��$?RT4�D��%"�t�ȓ3:��p*O�1eb�YG�թb�.�ȓv�~��g(R,�r��aN�E�Ȇȓ*DHprJ�2Nb"g�,C���ȓ��@�3�['e�:��N%(X��ȓ 㺌�"CCIX*PQ���3�%�ȓz^0D��L��;5$V�t�`���b��	�d��d��q�A��&Nr��?��m��cٯB��;�"��o'�ȓq�kQJ�:=1�Y`R��$y¥��D��LI��1_��ՂPŚ�>)f��?���3?� 
���$r�۫#(~10&N�N�<I���?7)����+i��a6T�(��/Ȫ��C�B��b{̵���$D������$�Π�FΦl���n#D����'�D��0:7#�c{F{7�4D�p��b��� �� �7x�j��U�3D�����z�e�7,J�z�R���O6��)�	g�'�� �� 1�j4��ab�|`�'Ӹ����F��YAH�Y<� �'=�!i'�C6R@Ep�bAe��؉�'0M���H�Z;6��(��pŨy�
�'� h�E��*���q��l/r�
�'VX��`��M�&-���٠Y�Z��
�'n|m8Q&A6Mք
0��K��%��'�j٨5�&u(����
\h�'�JT@d,]Q�A�N�a=>�	�'c*y�t!K1xrR���h�W�>P*��� *1��B.&C��ه�Ґ_��:�"O���0�ך:P���/��=���#"O�%�����C=�A��A���Q�"O΅���#^�J];uϟ�w�~X(�"O�e@GíX�`�s��)M�q�s"O�A⁓6NǼ}bANH�14JM��"O��ST���U� ^����"O4�X��R.?F��2FF	�o�H*�"O�Y��.
CJ�����η5��"O^���n�"2��䑺6�bI�C"O�YS#�	�A��Ԃ�n�	s"Ol5����ik��n�G܌��"O��Z"OZB8}됣�'<��!zr"O�5%��<z��B�'�F� ��"O�刐��;�l	G�2'Y��"O숊t��7�����F�4XZ��"O&�+r�Zג"�˨3��ѣ��*�y�N�"���6��*=�v*%����)�O���� }B���gѡ��A�"Oh�xq$��Y%z5J�%��>z�I�"O��!���	�E[�D�q<d�"�"OL�Ј	��c�'6.�1 "O.��#�âG� B� �v>T��"O���VA�N*|��"T�o� H��"O���(���Ή�������$"O��2!͏O��􇒖t{���"O�QB@E�yk���CЄ0k�L��"OH����-��u`K�juk�"O�x	`�_#��}�6�� �X�E"O%[��	�D3�B�G�<���ȗ"O�Y#q�� dEb�fL0�x�Yp"OrTs���$�L�`TCW�k�88Rg"O�Q	��ƥ�mi���5:�h�s"O���Ǌ=�l���	!?��<@�"O�Y��Ŝ;������V���"OB`�Qc@�D~q:#��`��R"O������<�p#4$�E����W"O`2�JE�����>O;�p��"OD�%��(gS�Y3�@=xTA@�"O�wGq��%���2[_F,["O@����ǊS�`�a+�6K�cc"O(���؟(}�$S'!��ML4��t"ORH�vDY�/.D���NGK8��D"O�TC2��L���p��MJh��5"OM�L�9/���m�<��R"O�����#p1���I�
g��1�"O��C"��+#�I�+
���� "O����J�]"ir�iZ"|U�"O:�8��YY�̓�J��K��qF"Ot�ve�3S
q/�� "O����;F̋#�+$B���"O.��7�A6+�Ɛ�4!��	��"O�����+B���@���d�ҥ"O�aQOP�r��)�7��
��"O�Hc�Ȏ�sY��3�� � v����"OL�҈;j�VHs�jO�CIB�"O����N;8�Y*V*K!@�4�%"O�P���ќ?;Ȉäi�~��1P"O��C�6V�3�.� �3�"O�{�PC1���1���p��\{"O`��'���]���8�"O���˜@�B���2=Ǫ���"On�(�d��4�:�����X=s�"O.� !��'=~v�ѱ�f���"O�  u"��ۯ"��83�Ąs�f1��"O���cM�~1��H�A˃Ad�-p6"O�����*������M�zNP�0f"Ot�Ua��M��`z��JH\c�"O��h�G��ݔȓ��ՌR4��h"O�L
p-��k�%���Z;>d�%"O�� �j'I��9��)=��ɫ�"O��IP���D*��+պ%N���"O��eb�Ri2(x����Y�dP��"Of��!�J`���Y8��)H"O
$Д(�
M��SM�jS�#"Ox2AV3gmN;�.���� c�"OP�	�Дrj��aw��/i�p�J�"O"5�"�5.b�`X�lċv�6�JA"Od=I��M(n���P��,y�H�:d"O�,��o�"z�"QA
U-�����y�Âa\�U:�/V)BDXI!�gE��ybA�L먱���4:L;��C��y"h�����j,}��)S���y�⋳8	����,m�pUZ�K$�y�/�-A�[�L��l>���(���ybϜ�0p$h@I"j��#�A+�y�m�UL��R�j�d��$�y���yO*]���R�_�l5I򂌎�ybI�XJ�9�E �3�z ��f��y���`u�ă6`��z�� ����yb�ʿ�. *0$��F4Ԭk����y�F��.��x��l]?V���r���y�L���	a���:7D� ՎB��y���(b��2uo�,�	�tm��y�� K1�DJĆ]�#s��o!�yH�9p2d	'�L�x;�G��yR��?&�N���S3����Ri���yb�P�kF�����Ѧ-�0٥�C?�y�C��#D�`�/= ��(0b'�y��<C�5��fZlJ.�Q�ל�y��p5�	���N�\?��b�Kߒ�y2���0�"dzqO&	��cV���yrF�x;b�E L4D\�p���y�)� ��i��̗ Vh	�$��$�y"ì�v؋�σ�
�q�1n�+�y2�E�bY豥�}_ �Q�˜��y��ѹ/��J�EI�o�m0qH��yb!�_��d��`ئ|:���p���yrc�2J���&�q%Q!�A3�y�D�2;/�g��f���n�/�y�B��|��P�++fN4"֧���yb�t�(yp+���ӥa��y�æ2���Z0.�J�`�L�$�y2�!�����LQ	dHb�#��y"c�7j� ɱI��~�
1K��:�y�l�x����i\n��(���X#�y�ʀ�@����Ł�.|C�F?�y���$�`��E��%�&�H)���yr�Z/Q��dl�3\֘����y/]�eW�ŘȂ��8�.W#�y�	��x�Ҥ�߸]K���Ȏ�yB�ۍ_Uj%�B�9M.�9#D�:�y  �y�Fy�t�HQ�UASd��y�H�5�<y����y�uX����yR.S�T�6`�t��t�:�R�(�y��uLt��J
Uw�d��?�y�)�
g0Z�2��'���a��ó�y�kWG. Xs�D�-���z����y
� ��I@O��q��Hv�;Ԏ���"O�|@�Ǝ;����d��H���k2"O����޴b7*p�3�Z�M:�"O��*pN8dQ���'F,��((�"Orh���M�}4A�'�0�H�"0"O�qH�B�*$\#�&�mڰ�Ӵ"O��b�/7��p����j�B�S`"O0i�!M�X�n ���-7����"O�%Xd�>M�ܥ� j˓:�D�C"O�yj����1�5��LH"Oj]�1�S�)~�3G����"O�8H�,Ȋ�:\��,]�9i��V"OH�K�d^��\9��מgWB;�"O��r�΁�k��Xwa�U���k"O���jí$��: ����"D��"O��t��)�>T�4�ՇOi�1k�"O�܀v
�*|U���cǆ^��@�"O �ᷯF:w�f �DF�o���b"O� ԍ !|��r��C�(5��"O�H���R7%�U0��K*O����"O1Ȅ+��0`0��hWo2���B"O<�����^�j���!(hh:d"O@�D��[��Ɖ�}"<��"Oĸ󁄛;��9$���#�m�"O�m!�9p#���D�J�@��"O���lʙR��]�M��HD�<����%�ʡ)@��
�N��E�<�E�9p4$�'�-/o��P��y�<�ѣ��9 蒬'��@cn~�<��Q,e�tdj��B,i����'�`�<aqϊ&B� ��\�
n�,[W��B�<A0hE�f6@�ӕ� ���yB��~�<��� ] �4�J$
D�"5K�x�<9�#�kD�z#��$6``Hrơ�u�<��?_ˊl���B�IR�Eb1��f�<�U�
(S��Zs��%Gl�K��Oy�<�4.���x���3�S-�~�<�)�7@Ӧ(��P���iaj |�<�!I\�a`��K�(�%� ��E�m�<�e+�47��H�PDd=ɵ"�r�<i�!F�`T.����k�v�+@��f�<��M�
0O>���E�EY�;���`�<����t�b5 Ek�3���b޸�y�슑%���ZcȨ{���@�KD�yR��t�� x��r�tiDϜ��y�Ę�!@���*p_���PaN�yR��.%TLc�Aň3!\��P��y��� O|�����/�T�7F��y"B�a����:WV��(E��y���0EhV��!��:3�б({B�����ْ��%<,��Ԣ��LlF؅ȓm�dpy�h��D�&��VO	�;-�؅ȓs�PD��@^!=Z$���Np{�a�ȓ{d���.��r i��M�a���9-.ћC�ѭ+$ЬxA��6m�9��Sq�U`�&ƉxH�����X)I���ȓ3�>���
�N ��31,�(u�2��O$�Y��ψc����'.�(؅�c�X�sΘl��hܡS�@�ȓ7�؀�g�<k=@-0¦òT{���b��iӒ)P�j^Dä�M5���ȓn>F��e��F�����G���t�ȓ]�򘚗G>�6!�WJ���d��=��0�Os�d�2�ؼw6��S�? )��
��X
�8i8�c%"O8�$N7v�	��BL��"OD����љ#e��s�'�dhBiX"O�<�%J�Q\́Ғ��}��)�0"O@k"��`���&��4��T�%"O\�At
^)��X �W���z�"OP�A����~���"0,\=]	|� �"O���lh�hDk˨h��8��"O��R�_4I�Ps j��Q:�("O�U�5�ˀ�H�H����"O i��fK�>@x�W&)�t�W"O�`�E��R�p�jk��v� �"O<���7BL����ҁ�"Of|�"�C2VȄ�T�8
q�c�"OB��w��(J��Hp��/�l��"OX�9��`U�&Ʊfs1"O� �A�����#"��0�1t"O:]�# �����e�S#���"OD��ǈP�[�z��O��d�=�s"O5hh������n�/C�xP"OH��A-A}*0�P�LP�$�(y�"O�Y W��B�)�!%" S�"OH�µ�R�~����Lw
��c"Ot@TS�
�� ��p�ȕ��"O�,٠
�>����q�ɗaq��c�"O¥*"Ǝ;�	AU�S�jh"O:-�l��h QA��c��9�C"ObT��
I�2$Z�� �T�m�8s�"O�hөU�M�v�qၘ�PӾ�@"OL!`��!u�3�\ l�����'�����Q�{-f�� c��`���z�'�A��U�]��WLV�Vgf�3	�'Ѹ-�sJ(�tt��ǆ�L�N1i�'=t���a>������E�����'�,��#������;`��9	�[�'h��Q!JşpJd�7G�6�la��'����j_%�}��i	0y`���'�.K�N�f�b@ҕ!���&�J�'�"ѡ� �y�L!(Ua�j�"�k�'���R`��bWB��,��/&,
�'��ԣРݠ+`��v�U!����'F�@�Qe�MPD��E�ړ�����oq��dA�m�tM0�͛!@|���
�D�q�T80�y���5�j1�ȓ��K�a�0�X�C��iJ�(U�t�<��Q1-���Ӳ�9;7~�u�<�î��<�X]CU1	��	���Ot�<i�&T�f�8����-+���J�<��NC��¡�JȤ<9�!q�<	r�F&?��x�)�2O,���y�<�0#�:E���%#0�@<�d�vy2�)�'5:H05'S��x��fi9r��Y�ʓR��M �o�[�D"S�:�\C�I,U�x@���=;v�{�$�v�z��hO�>9��ϑ\X�(�)����7D�t��'��
~���儝�@C�,2�2D��a�B	�R7BV s��"sͭ$���p�`A+d�ˀT���ᷥ_ 5��%"OF� �X+��K.��<��E���'Ց�,
�.�!	X�I�o<@.�;��"D��J2�A�.b�4����z�^h�$D� s���2/��cʤae��k�"D���&�"U��Ac暛�X��Uk>D�@�ׇ�8�2ujQ�[�G3y�;D�� ���
�2���J���,�l!H��d:�S��V�6u#��5�2${&�M!���@J�����?� ���M��].�O
���v������}n�U�B�CI�}R��:���Q�fM�ʍ!s��x�� &D�� ֪Z R�Q��9jR�DJ�&ړ�0|�	X��XɆĞ�6{B��s�GX���O|��B�<���#`�!3�j���鉂�hO�i�?�������D �r�Z��!��O��h H2M�f�s�1�,��i��Y'�vqiq�G��C�֊���!�S�O͊T[������qŌ�*�L��'��a��΃�.`zt��X�X=�y�'��O1�Z���c 28�������#O���ŕxb�'+B�z#�P�5��b��2ͤP	�'ўb?��c����pnǘp�l�ѳR�K�,��I���=ٖ�Z�*3��`�CژWpN�H�#I�<�Q��'�()��
I*`�>�	"%�y?�'6�OQ>��$ [�ʵ��T�x5"��.���y�D̴"���Qc��s�>�������Ą���>1cO�$@2��K��4'��<a��1x8�I�Ɂ
���Xa�L,�옇�IT�	.=�Z숕���<n�ţaŒ�h��C�2���riކTB��M������>�!�K���
Vȉ� �z�;P��u����I䟰7Ǎ��jx�r�_E@�����8D�p��g�:Z�{Em^&]�+�P�a~RW����ՙ3� ��j]�5Fp �RF7D�@��c��1��L�T<K@p<���'D�D����	vbn]⯁�k� �C��)D�����!۰���o
�0y�ƨ*D�$�&mЃ��KCn�4\(\v�+D�PSs�G�  �"b.ƷJ�+�b�>)��Z����tHs��<��ϕ�)P���)τmq�d�8���"5L�G��A��bﺁ�e�݄w�Jc N�Ti�1̓�hO?�3
��?
�@�[�$Ѡ�:D�d�a	�d	��K�'~� E@4D���p�W�Z��)15�_�=�<��1�/�OZ�	�>��z�N�����Ip�Кl�"B��?h3��9����P�8CWKP�w��C�	�Zx(�0qI�2��6�O<�C��.�~�JӀO[Щ��ͶT�t��hO>):�	+r��,Bt�[<fn��G2LO��9!��:!��UH�)9P��I0�v���{K�	2P�yQ�/%ULq�ժ-D��@����pK�,i�D� ��,D���%��6h�@a02k	:A(	:G6D���C.+�(��aD��.*iؒ�5D�( ��ǞW�j\�4�CH�:�d4}��'�ܐ:!��u��!�"/�z��㓱ybT�t�Gn֧j�4����t�4��!�<����'�Dxr��1-�Ȉ�%���l2T�35�=D��@����`!�1� �G�+�Ju�>��(�O�!��D�>��;`�����25�'�F�����5�%@)J>x�G�B�p�!�D\\L0�cmC�B>�d�_���'Na|�'��]���{�-��-~�Ԅ�.�y"!D�-����D�@��d����{Ӓ#<E�͙� �ճ� �7�� �G��y&� |!��qUbʌ2��T���~��)�')�^�q'�[=J��I�J4>�ȓ(�܌�B��9��,�,�!#<p�ȓ\� �9E`�A5��zQ�y 5����s�� �4���1)B��iD�1H��H5"O�����-��$P�"[0v��W����I�sb�y ��Px�a��_�C�ɻY�Tb%A�+ lV�a���LB��l��UBJ>Mi�}cac�S,B�	9]�� �j�&;��q� �{9�C�Ɋ?'���8������0wU�C��&G�f���o,��P1�&]%}�C��9ah�h*e#C�UG\0"�ܻSVDB�	�����eJ�/�>$8g�[�~[FB�ɑE�T��B�۠\+�D�b6,"=ǓN���1��6��`��m��1���ȓ쒅yUb�.~p�jBT�e�ȓp����G�54�`����H���|��6��yC (~�R�Nӓ�d��O���#��.��4�e��	ʘԅȓS�~M�CE��Q%4�c7�'nⅅ�=x����ʀ~'�M÷�)#x�,��}�9ka��Fo��R$��(b7�ĄȓD�N	�H֦D�vJ#5L,�ȓ���q"�+Y��,ڤ�_˖��u��y���9&��ɗ���4L��}?�-��	�R/�hy�(طA��ԇȓ\���#��{���oQ2'A�Շ�D�I�la�f�d�0%8d����0�p�g��[%��&�3?Ў��ȓ��h��
��9s
�����_z0��2E0�P���7-�ȍ�#LM6����>1�jI��ȱ� f��m��]I��)�'�|��c�6�ȸҡWOh�(�ܴ�(O~�=ͧ3
�"��)�|�΃9@Ȯh��	x�ßd:c��01\��FLݱ�<)��{��F{��	�4�b-^�-�4��>�!��(�P�z�g�`��ȉm�S�!��?<"�I:`ŉ�:�h\k��7j�ў����S�y�D�9�Ry�.��/��C�ɇy�����%M3�Y� T.-��7MC�	1�~���ig�Epa��1h@j	:$M�FX��r�'Z�gͲu`( �C��9�	@��D9O��sEI؟�l*��rY4�
5"O���3,��ŢԂ�FU� E���';O���>K*D�!�ޡxT:���ď48�!��-�R����p���)�!��U�&lǄ_�R@��b�@�r!��şi�4̰2�"I����]d!��_�f6��Ǉ�<-����n#C^!�L�6�U	��Qx�a�.��@a}�6?YR�K��ı���)��,ے��t�<�5��eU��s/�L���%�r�<� ��Bj �gi?5��dsRq�<ae㔕T�\�PfA,J$�b0�ND�'�x"'��^����-|M�p���y2B߹U�" +ƈ�?J�9釩)�?a�'��<B$�M�y[R�2u�ڔ(5�:�'�>L���[�V[|eK3`K�`\��'R�]Z��5.���s�ƏDu�D�
�'��$����~�ʜ���<�Z��'�A�e�����zg�:�^u�
�'�4���"�zs��Ѥ�ڃ?�r���9���j�S����!��-�� �ȓJ�^��J�|ݑ�#E	+���D
�)pT�Ҥ[u���=Q^4��d$ biX@.<5A6JI-��ȓ֘��Ӯ� ML��G�S��Ʊ��S�? :9�R�&y���X�O�5�Ɓ��"OٓX*,t��0I�:`�@�"O:H�璟�<ћ�ꁰ&����"OX�J��ߋd� ��I��m�Sw"O����nӺZ��b��N�rdx�"O��ǩ�ܔ�%�A8��)�"O�-`��ג%�'%��8�A�3"ONQo��2f�Z<ba
�W ڨ��"O���#�
a��-z��4;{`1U"O��ffک�Vtke�[�lf¨G"O����I�?
d�;�ϔF�J\�"Oh����+P=.s�	9T�Za"Od�`��$o�N�;wE
&M|���"ON�j��W[�@�1E6l�6��p"O`��šΐ?�i�jU>�*`�p"O6��4GQR����J6h��a��"OFIqB�(X��X��J��*H�"O�=��%f��X���D �2�"O6m�2��=,uz�.�& ���"OA���C�й��
�=H���"OD|Q"d�'%�Xss�W��͚E"O�h�I�.=�Vx+��C�V;x]�G"O���W�۵~3 �p��({#N�q"O&y����e�<�*�y)⼉"O�Zw�	��� 	�/h]��"Ope��J�/o��2�i^�&С�"O�h	W��='�~])�h�M��L[V"OH���F�_����d���9�"O��`�n�|:�u��$�]�"O�\j��W�M{b{l�%"O����aB:k�*�8�nV�}Yth3"Oҍ��'�4ʶ%B��\	|j�""OK�Zl���Gh)e�Z	Z��	��yrM�x�\���f����'�yb�D=no������:XK����Ԍ�y�_�h�T�(����+D"���A���y�m�;w��8���
/�dy�q'R"�yn]?/Y��QA��.T�4�z�����y"��.[�^!!uD��BC��0�	�yB^�+,�H) i�MܒI;A"F�y2N!'�hL3��%v���I��@�y�,�(>�My��/uz��m ��y�H 5�(��Tū}N����yR"�<e�P�"�9gŦlse��:�y� K�E��I� o�����׶�y���K-l��F�J&fո8�����y"�E:ypX�F�� [ �+G���yb�O�F��x0�L���D��y��Λfg�[�`ը8:���p���y�B:;Y �&�L�i��a����y�g��XḄ[��n= p�N��y��+8Fx�*1@ҲW��!���3�y��M�dے�y�!O1����kǛ�y�m�{eeA7�C2�¨$�$�ybMǧp� �D���s@t%��D��y� �H��"���U(�R!�yr��N��ЮҺ�Z�G���yB"���1e+���쩁�����yb�R��|�K��ɚ�ǃ��y"��J�Fd��;pw p�!��y��0N��l!Bk�l��1s�-��y��в#k��� �,a4�ٛE��y���!�j���,M�f��:再��y���5i8�1@�Q�c��ͲԮ��y
� "	Z��Qb�^�CfkK���=�"O0�S��%�A:�9fݒe�"O�|�b�	�r,�glǹx�XM�`"O�4٢�\�.H顴�[./ɚ!c!"O��ƕ3Z�d�D��D�"O腂,�6]�����*�^,D�4"O����_��ɲ/�h-8�"O�A���\��墁M��,al ��"O��۲ꒀ�����NW���"O�t2�

_rx��p�٪WA�E{0"O�`r��_�
	՘���|L���"O��w��;SY�̳cA�n3L�
p"O&}*�o��@�&|��B �=��j�"O�9�da�=Q	�R�A^�6p\r"Oژc,XD(as1B�rvL�'��1�6�U�|2����̾L똈�Ι&� ���3D���g�R"s`���Ή�1y�]�G�p�.Tj�N-�k�(|O^Q�����"�ʍ�"쀲Q�H��	�s&��̆&�ZUlZ�'mf� ��gXF�!��s=��'����FW�r�y �H�-����{"$Z�c��]�e�͞6��>�8G�;�x��Wfd�p� ,D��y���]��;T�A"b#�u���H�a�$m�U�й��+�(���zKFH�NM�4��=pP@�-�vB�	7H(���j�2PC��`ꙶ�Dp��"�
Z�~c�����=Y�+�?Rm��ր׿+��Q�0�Ca��<ȅ��z�2�� �E��õ	�+�,}[�Lܹcg6�4���3��DE��x��d:h6�J�h)�$bQ�A/��'I��Q��8�,8���iO?��Ū2C:LOĩ��B�����D,*2Ԭˌy��,+0ШGz2�>��q��E�jx���a/�'#E��x��eYX�H��֝�<��Q�%E�h{���q�Ok̕^"���\>�����0����K%=��L���'��L��P$ @j1�D����4)��#aJD�H*N���c��p����2��8�BP���[8 ��9��E�T qøe 6A��!�t��'0!0��ox�����\��.e9��8�%P{8XnE��P�H֣΍!eju�A���9Oj8�hҩ�y�h�8vx���V�. ���yA̐�0?)#H�F�ʑ�eHK�P��z���[t�h(0��X���bu.N $L�O��?����.GRR�Gg0#�r�PꎑJ�� �S��h�&�D|R�Y/D�y�)\� vpb���&C��.p���Q�
.H�
�<*j>��Rg�+��I�"�O:й�LJk�&yA@�K�R}���'ɠ�ƈ�� ���TԅO�"������?qi0�M�Fa��9�2��F�!�\3�ǎgƀ�"O.,+����0x���n`hE�����G���p0�������֕,k>4��O�6h��kkpu�6���(��6nYH!�1u���l�Tx����{(S�J��-B ��B-8p��F� ��S "��:Ȫ#�'n�%9@�0'V)Dx��1[/���Ц�f��L�ԥ:�hO���!,։`j0��*(0&]�Ί��u7jӸ'��is�MVA��S'���MׄV�o�a*����ڦHX�zP��A���bC(��	-l����aԞZ�)q���;���ʶ؟����1��T��;p�<�U��1	0��H�R�!�l��%"��r-�C�JR+^���FΏZ'H�2��N8�6���/���K�Y\$����q����L����M��ɤ��U�E%��NA�L� DܻP���X7��\RN!��dM�Hʥ#EJH����I�vO�Ղć�6w e�Dk0�^�
 ��H�_�촘�&N�.�l��h�����G*[P��wEM�h�V���e�*\O���+��&��� ї�؜�g7O` rbo؏2 ]9�jM(zr����D��(zs�����7T���#�%K���PHMkS!�
/�TS `âQ6MX�'\�FN��0�b��(�ᓅf~�YY�$��(�L{ @#}�i�){�E��*r�8 �
��%�}[�~"�d��<��I!�Z=����b���_��ja��{B�8N�4�+&�:b>7� �x	Da�6��!B.L p�d����C j��c9RQb �'��S(4nm�Wb��\�j��HI�&���
�*��FO���D.!�%03O�5���q��3?Y�!��=-Z8c?�K� I�dY4G�"�j��V
�*����JWq��D�/1�� ��Џ� =�3��8I�~�.o`�8~��d�-7��(�@�0}bipމ@��E:�Uas
[.T�e@/4��U��'V^�1��.�?>�<����ڡQ@pj�݀,�>��K� ���		���|nڞv�j)S�K��5��Ȇ0^�Z����6�4���1��� V���gS�6 ��&L�zt�ÓQ���P� �7f���#�'-e�Kt���Be..� ͲL>���,(�8劄"0�S�C�lMBqh�a�2,���8UT8��f���-�(�ȓ�:�0�T�r�&�0&���� �B���aI~u#c��v��=�;-tEjr�}�Z�EOc�j��ƓIq(�b��5�ԁ��H�|ӂ(JEg�/@�h�h=�O�p�5Ȇ7uPX��hŚ^D(\G�'X@�(D�ZB T�'�B4 �.˃9�d�2#G'.z��'�dUД�I��1Z �B�F�:O>Q4��A�H�օ͈������L=(�X�b�
=�2��"O5��Gϯn>�kԣLd](�,�Y��O*�W�3?��FЛ:�������`����Uz�<�6�ZCv�(��ŔSy���Ү�0o"���$�L��@S�G�=BJ�]�%잭+
D���9D�H�D�[�4�|x+��>ͰѤ5D�غTB�g�2��R���?'H�+�,D�8�Q UM*�	�':(DV�8"�*D���s�z1lIKDC�.��)�b)D���j��C���y5�S��4+$D�(�F�#b9 �K�9�.��@/D��BGኌ �0�V����m���8D�l����9rH�,��CY�J�*MP�=D����捙js�����	p.>�Q��<P�NS%�㞢|�&6\̻`�$9�����AG}�<9T@h�Go�lBy�g�yS�O��Bo^5����W�:<�9EL������-��7��~���\>��P(�X��ͫC*�)��Au��	��t��R�E�O/LO�i�2ɘ�] ")[�E M�����	&)��Q�� �W]�Y[��}��ȪVเ�`ٟ[Mt@p�@ȉ��B�4Erx`F/�$+LP�A�J�9?����x.2iB��HWL�!>2,�ǲ��Oz�ac�Ls9;�BCv����'&�IC��L7`��$Pqhі2��q0���TSF���
QI��Z��S-&�PБ �:B�����E�� �!�q 6�Ob���F�*.^���ϿP7���Dɖv �M�E�
�?%��I��DQW�>,O��`֯���I�Ə3zξ	���d����Q�nb�L[�^���0�o�]�Mہ��
���)��!��_�ΙJ��J�*���wg�����uV�M��?9�:�D�.@�T�0�E���O_XY��׳=���(R)�)`���'���$cضe(�Bl%q��X���M6�MF���,�hD:m�5��'!_��$�X�`�^�Th�(�OE��q�&�OjP�@�T�n��Y-��x�x tEG�z��] �'(ы�㘡(?Ї��hݼ�p���8'-zx)�N#'������OS�T��� �b �͑�	U�+��tt(F B�I.h��	��*�xZH��؍<��>��jl� "|Z���d;p5(��o.��*�h�y�<�K(v�&�@�fŁ[bR�hKz�<I�ßM�@�!�D�U&��I��v�<1��_�`F�V/:.�4)ԭ�yr��(�e(���;6D���L���y� NN0T�t���#���j��y"�6AU���ǖ���[#���y2�C�"�2�!#~H��C��M��y�m_�ar�xfA
)]��e�*�yR�٣cV�pk�j��V<���`��6�y�M\�[:� �AE���r���y��B!�#�F�*�,�G��y�%O�w�� S`Q�`X�k7%���y���+|��1x܉ք�	�y���|Ռ��v��q���󣑖�y���y�#� Y�z���lT��y�Έ���q���2���ˍ�y��|�h���ٓY�|pJ	�y+�i����a�9����y�! U$�Wn]�p���"��y
� �T�!�WV�I�
۾��6"O�D�W&ԛRg2�J���~���C"O0�jT�;��IU�L�	�U"Oތb�A�b.�$Q3�QUn�e	�"O�!�Ҥ�-꜔R"�O9*�L��3"O�s�$��))t� �#W4'���"O���ՙf$�q���/g�t�2�"O��ӕ�7f�����Aݞ#� y�"O0hK��X>Z��@�$^8��"O� H��ގ���yth�#��s"O@ՂD%��g�&���I�j����"O4i��L.>=�Ȫ�m^����"O m�d�P�V���[ k�@�@�Ȗ"O4$�D�j֪�2E*[�3T��V"OJ������i�|�(�>Z�JD��"O �IŃY-Q_v�R�Y

���Aa"O��c�ާ,;8M��cъ���)�"Or�sU"��b/�|�#�3����"O�i�Am�V�Apԁ�M�ɸ�"O��z��:,F�Aa�6���2"Ou��b�K: |(����$�"OV=���.���%��{פ("O�̸B�D�n��AJR�q�c"Oj��hA���M��X��v=�V"O����%M(�P���	��E�7"OF]CQ��)N�8�0�Ʌ6�q t"O
E�.Ğr�05��#���@�"O"h���%>)S L�u�yw"Ol<�����@)a1��?-� ْ"O����f�'\�feΎ
�m��"O:[&Ì�u<ܝ��� 6���@4"O ��R�T��}A�hXn9 �"O"؉֏F~��՛`���-[�A��"O�I��W;D~�u�0G���V"O����G
wi���(e�*�y$"O� ����9(�
�{ �4n}� @�"O2�-�-	��0 ̹Fv��	!"O���ևӞGK��u�	���`�>D���b��7"0�(��x���H�+D�l06��Oܮ�q��?��H���'D����@�?B�0��0 ��~�@"�C"D���@�*
�+d>�Zg�
�y���`g��g�q�105o܅�yR�љ;��yHeO����������y2KlX�ƒ.z�](1�� �y�.N�_&��K����~�0��&] �yʍ<9yr�/W<p��0�"�y�����%Pq�ְwjN��uC9�yri\*ne���iֈSz���ecI�y�e��*'<-�0l��OLѸ%����yB$� S�%#c�� m�yȅ�*�y��ٱ;����u%K�g�F�A$�yB��;۞`y5��N���;�#��y"�ʶ�0ē `�@��]�`e��y
So#@�@� A�:Q�f����ybN�$h��Q���U��pv-���y��:U��ZWo�A&-��N��y���4�hr�+9��hX� ^��y�MN��}HĮ�I|$ɠ�
��yr`�r�\|���;B�j���R��y�!XzbY��'0����� ]��y� �|�f��TMY�{�x� W�ص�yB�F`3Pb���h༰!i�(�y�p��z�� �p2� ���y
� ����D/�lt��b��*�~�P�"O�$�Qo5�"Кf
ΐa�6� �"O����$�b�u R膙b��x{�"O4}�d��=6]
��$���'y��sd"O������h��C�Q=Ch8M�B"O��:��1}�r��w�-Ze��B "O�,!�/������;;��e�"O�����$k��\x��S�\�l��S"OlJ���|W�K�m��6K�"Oʩ1��T@��%���J��}p"O2} �I֔% ���@ *uxHX�"O�h$�F#V�0y��n�3`ԕ�3"O�Y�D�V.=ERչB��Mr`�j�"O��{4ɝ�x
r\"2'JR}��"O*��&N��8�0��J�� J�-2"O�1���v���D�
�@��Q"Orܨ��;1�yE@�]�n��B"O(��b慌\N	��>ry�(�e"OXI�S`�y�]Cw xP�}2��4:b����|������8|�F�v������!D��:��yc�d��
[��p��o|��`sόn�C��,�R����O E�̣G#;\O0I�s倐*�����Lx�ԉ$ժvN��W�C%D�q�"O��"���|����$AJ�$!�d&��D�#["}a�,4P8��^t�$�HᤜT�<A7�E�z�����ƈa7V}b�C�q�B��
��.��	�9Q>˓Nb��k禝8&�|� �E�dy
X��z[���#�(�3FE�.h|�j����J�:aa{r�S/^K��h6,�-:\��b���p=�"k��/�����E�<�M{@�S$XP򯁝r'�!���T�<qg��*d����$����h4NFd�T�vJ�c9n�D1��Ɇ$��h����]OVD�UȔ+D�h�@aB^O��h��ē�g�����`;�Ȇ��:#�0�!f�z؄�'�`G�,O��`�a	E�zH��B>cnC�i�><��H_(��|"$�
V�]p��<ڨu�e�MS�*�=	+tU��`{�(r
�4���Z�ݦi+�ő����m�71d�@j�+��q�4Ig -��=�0ʓsت�'8�V���MF�h���V(D���hА��t4Od XU/I(���9���ئ���,N`z!��.Yq\4z�"O��ya[���fi�Y}��"4)]����1� b�2�	�@��!���R�u�~첑G��G��X�3�-|O �I��
7;{� B�4,xT*V�ۡ!Qv�;�cь =���E�g�-Jbŗ{��c�U����#�C=,�E�&�Ig�|�p o%/ E�5[�b,6+��|��(ź7��Qz�O���Qp ���y2/e�yx�@5��� �%vN�2!$U��$ʺsVp��.��O�m����&��n{�E����E!��3°q�DAv�|��\�V�� [ql�Oi�1�l؟�{��O��m��቞]P����M�s�d��D��0Y����<N�~ �uꁟ�M���S�8�Q�����iZ���'B��q�U��h�zp��	XL�է��n/tu�DH�3�����#&ո��9�B�Ov}�d���	�<c"�0A�.��!�%]j�!�d�	m����d�^�;������ޤ��f�O��O?�	8>V�=а�D6;l����R?,6�C�	�F�����:�ƼJ�NB,�D�������$�'8��z%�%d|}��I�Y��$)�'TZ�sa�NJ��	!�愆i���r�O��bM��p=��&��1��Q�G���@F�dx�� 拥KoV�`�B� l��e��ա�N-q0��[�<	��-r�x���"g�D@���_X�'��A�F�l8��E�d�[�O^�3��]Y�<ٷ�.�����3-@�y��ئ�1 Z'1�� W�>E�ܴu۞�	wf�z��b�D��9R�����p�Z�$U%��ɪY��F��%��y� ���&B[�djN�,�'��}6�Kv�'a�m�r��'��w+ݹ yTIcH�%T�(�b04�� 
 V�׾���iĢ��z`�1v
@cG|�Ob�vJ�gIf��p�8}"Lt���4��Z�\H�眽dzŻu�54������<xd�����3��,k�+/H��s�;*xF((K�����s^�b>7�Vt]dt��P\�D��a�$Fa�y�I�X�l���d}�(+z]DT�w�КM5��H5�ȼ����<I��p����*��<q��g�t$�v�X�fb�ƭ�U��!av����Kq��EÆAʊ&��MOٰ9�ǧC�@^��؁�=D�ȧF�o�%�,_�'��ݐ��z`j��N���QK������3�i��rc��U!Hi���t `)[�O#4� �6&�h{")܂��̺ �ؼbFtX�@7%�a}2B��3��y���4}�~���\��<��G�6x�j��Q�>iE���y\�����|U�h���Q�<��B$_*%3��"-Θ���C[R�I",˔����`�?ek��A�*�J�r3D�|�6hH��:D�<�'��
^\���%��1W�"Mtv'��!�?�g~���&c���1m�+� 0��hS	�yj�1M#ZD;E�[�!�-�����m�����4�0?��C�y-dA(�-
4_��d��K�<ǌ��}U�,2L*chh@�{�<��[(�:�l
�R��\b`��x�<��k��R,RTؑ+U"+e��Za^a�<�5 ?4� %�c��_|b,p�Gk�<-E5dQ�GfښXA�P���ۇf5�C�I�����&%�E��$stȘ�J�C��+�8A#��A>��#`�1 vB�	LAt�Z��e�@�K��fk0B�I�D8*�s�S��@�cF�2��˓LW8@B#)/�)ʧ VP�8��W�R2T�K�87e�ȓP/tx�d�b�hs!��7qBX%����F�wk怄�	�XD59R��6^.ŠP!��B����$V0|)�Ɂa�t���E?>�L)˅���@�'-��9F
n��K��D	I>�� �J S_-���7�8B��1�����2Y�rc����s]\+��턤�A�|�F���5-R|�$�G$[�����G�W2��09,�b�dF}:.�/�Y*�����OY�������� �2�h������'fqq�B�a�ƭ�O	4S�F<,�Ji�)q�Ȭ �` 2��S8W��%�TI�����%�Z!Y�.��?�O����4FC��Kmhv:���Ɇt"H����?�6G	g�D�g",O.��f�@mD�x��.xw"����:j���QtFU�E�R�Ү+U0�������(A%�&(��i��$Fd���H�~-k�o�7B�Ĺ��)9����}q�	ZU.Ϳ*ZN��]�W����[ ��O2�M e�+m� ҫ��K�h@��'� �PpB�} ���C˭KP��#X!�wAû8�Ȓ��A��ħs5x|%�|��%ԑ�rzvN)X\1Ia� �O
t��e�e�%���a�� F�>A4��'�<y8���3�����#hI�D���ŕK����T�����ʪN�Uk�ƔW���� �q[��H3&E4W�hB�	-W�(��j
>tA�`ϝ"�f�>�W��x��"|�`l�%�N�꧉ͅ[�@=�0�ZS�<iVA	�m���q��^�29| �uh�t�<w��$/;�Us����6�����u�<)#��<���6F�/올�ENv�<Ѧ�ah���P�}�$hk'�Qs�<q�f���:z8��뤈��2�HC��00��Ո����cl�B�օ�:C��TGt��F�lQ��R�W�]}C�ɷz(�p��	/}?F� $��j�B�I=HCl�`�Ύ!dz$ٕNJ"�<C�I�Cj��c�C�Gq"pS��ˌ'5�B�	��$ c��QS��yv���g��B�	3}�PT�!N4-��!9����C"O�����A�i`�(A΂�pT��"O�����RtձF�;q�$�d"ON����<8D2�M��qH�#�"O� �]�c*9$Vq��-/bsv��c"O��j� �>�6��@�N�PV��y�"OLax%��Y��pI���-^ ��c"O�1���� ��da����xuha"OF�
�)Bռ�2 ��p�I�"O
1 ҅/�����ED�f��?D�����H<Q{��P-Z#����&!D�����ڔ> 4�k#��0�0X� <D�X7A�?T���
��a���s$*O",R1'ܳ'����B�q�x�U"Od�!�M�$�bݩ� �8e���Z"O�����v�����A�i��J%"O�acoͺp�2=0s/��+W�8�"O@I@�R0�1J' �*zI�=A�"O��f�W*C�x�\#D��"O�`�$
P@0�ae˘�y�@0""O�a� ΀B貜 d���w��$��"O��a�nݲJx4�1a/����"O8u2�-/x�В쑝G���
�"O��:v�L�_����ƋD�A��"O^�R�g�;-,$�$͐�V�� "O5�aa�S ia�lÖI\D��"O�98aƪ2��A�CŃ�$B��"O
�B��-�8�DޝG h��"O���wN�-����E�ɤ[�2L�4"O0�0AO/n$�(b�o�� QA"O �c��Ú~otq��A�R��0�"O�]�r�%װ��BG��FM��c"O�b$`պJp�ٓPf��9b�h"O|���H�~�r��Q�EłU��"Oր����3#�Պ��$JM�`��ɣ�~��iY!`{<HW��4_n%C!D%qV1Ol!K1�'��LQ2��#1<r�S��Bs��[
�';t9��֖A�a�?bZ��O���dΞR=N�LH:3+*U)��@}��G�*�q�V�N�m>8`�hB[:��'�铺0|�!<��R؆6�q$�M?�I�D{2��<���N=/5�4�'eX�YDAR�+X�	,�y��i��С��P�O��,x��*KG�0Ӕ�C+A^ܴ�Z�\2Ҧ�f?y�.�?�J�g}�U>a@��)_O\0�O' �t9��tl�������TJR%���2��߂>��X�#�Y�
�&�	�S���f�(��i�|Q�P��H�&d���7@��~ꛆ�0��$�?�F�I~�S���D�(��_�x2�FA���'��	�{K�?M24fP�Tl�q[2jA��8	�(?�D�¦Q�=�'�zX��5i�H 蘪�o�
�h��q�T���)���H<�O
�O��Lz�k�	-�ȼK�a���������$W�T�lZw�<��'~a���gF(�
TU� 0,��!1n:Hyv��)@$�D�>E����a�%k����$��ض�81����[� ��(�����$!���v���xa�ܲPa˩�H{cb�����-�d`+Q��	aw�m�O|��cMJ?Uy(X���1n���:צ�[��µ]l�姨��I3������`�?P��b��#�PR��� �??1J~
u��4˭T��d�M�CɈ����2��B��6A��	�E]^�ᓉĂ���͛�`� qb�>/�:��P�� )R�q!t���#���Bp�I;�.X��	5,��P�Y����ʶO�eQ@Ʋ�0|��A��1B��#�~hۖ�����Q V��"}��37�v��"'�bu`�����c�<	��H3d�<Ak�k�#��R `�<������ڗ���L3<M�@IT�<�&�"lJb|S��o!���5�h�<	"C�,c���7/J�woҍ��~�<�eF8t����vȇ�Nݶ耳N�w�<����B�tkG�Q�M�.|h�ML�<��z���I` ������ TR�<!���?����F�Q�1�K�<� h�:�H�4"D����J" ��)�"O��r& ��~�~ �M�L��2"O��C�تX��ao[*=��Q$"O$���E�h*�q��G�;<���"O�� R�7��`#� ��v�R"O�)[�$�!k��Xx�n�53j���"O:0��Q�P�y:�Q:h�`#"OlQP3�D�	�
Ysǅ�s�Dв"O����e'x=�E
y�贉�"O0A�"LX�%`t���-��]�P"O��"0�G1�ܠ��$Ƈ#�L9@"O �ȶd(�@��,o���y�"OhX;Gm�9^%�3���h-P��"On��'�;<9�-�<&Ȍ�[e"O>��� �`�,a(���"O�PS���
j����d��:d"O&�ȆA׎8i��!	�^,��"O����Ԯ0�8���Μ#jڮ�"1"O�	P��^&p�eYn�	n8AJ�"Ou�R)Rx?���>M��pp"O�K2�!�N�@�_"K�D	�d"O�rE�!�P�Ј�P}����"Ol���
�,�N��h]2#n����"O���\>q��T��mW"�"O�@0T���M>�|hƈ>"&��"O^y�S&�����1�R��"O p�r�H�|�< ���r��� "O=�l����pi�� �r��"O1'�	/_�`�E
�3pܒr"O��B ػu���aS�D�S�Z"O6�"�T2�1���3%A�i9Q"O.1�P��kPb��fJR�
^�H"Opqwh(!ht�ںHָ�;7"O���B�*Q8	iץ��dpt"O��3�(��͙��ĪU�-��"O�-3C�� �VIj`G���d�T"O���I�����ďΩ��E1�"O��֡��q�� ��뒘Y�����"O<���@r>�E��I���@q�"O29��h�:	�x�jti��6�Y(�"O̍ӪP�H�1��k��I{"Oj��&�*>��l���)�Ƽ"�"O蠹�<8@lcWM����ʷ"O��I6ef����+����i"O�	�A��c�na���%��"O�j�(�>ݩI�c�xr#"O4�b!X9rڤ�bh�IP\��"O��d썂H-:4"%��>X;ʙ��"O�e��*�)錍k�׼e*$�b�"O��!0 ���!�*U>�@:"O�(���*i�����͵'�ԓt"O �"v�FU�������
��"OAPTŘVh��X�iؾ ���"Oj	sj�
M�tpZ�*^�A�lu�f"O�y�#F]s�WJ6db�8t"O��Gi�<}�-%(�s؛"One�U�ѡj�x��(M:3YL]8s"O6���O������Ŕ(FD��"OD�a�Q�N�Nx��ŐN	���"O>,y� N�HR�)�t�͝f l"�"O6�!b��ql��Y #����"Oԙ��e��Q4B�y%��= VТ�"OH%ʆƐ�M�X$ˣ��"y4��"O�A�����s���:s�i@�"O� �����8O�� `A
�u�q�D"O!Q� P���yX���"b�"O00�tHR ��(֮����AX2"O�� �Z���Q��'�D3�"Ođ��C#eo�8Bgڮc�<;v"OX�Y�G��a�A+��f�H�v"O�Y���]�«��Dȶ!�6"O�Y:4D(H�B09�!J�!���15"OhըEV3y�����?:Ĳ�s�"OJ}9g$�6%9!Ś!Z�|��$"O2l��`��TV�iRF�'��̲Q"O:}+PFбk���{�Hԗ�x�B�"O.H�Ĉ:K���Q(�
>���� "Od�d�ҟx����!� �,:V"O�M��<z�ܡ�a\�Xi��"O�iA��4�<d;U�!Pip�v"Ot��O�'�t-��P�Da��"O��CeɍX�� &���&���b"O�q��f�'<��R��åb9��b"O��
f�U?,.8:&�W"k%"O2�!�
��e`��H�SN��0�"O�5�PlǑe�L؊�bZ$�T3�"O�d�B3Vހ!#��E#3x�m�T"OX��2��/��ƩN���"O8�	z�.���Ea�V5��"Ot���a�_�n����+}��4�6"O:� g���g��}��횙&���b�"O����M��^�	Lo�6�A�"O��!n����J�."�nUc7"O�cf�5ܔ��1 �c�(�k�"O���-I#<�8�E�5o��tx$"O����L�XwN�3�Z���B"O�фi�8&�]V'��tބ	�&"O͡�)%��S�' + ��k�"OV����2���1CFH�\-i�"Oha��)�n^�ZA�?q@, �"OͪA╁$��M��hE�q/�X"O&��Å���.@����# &�8�"OT��%��<���Au� *$1�s"O:,���U��
E 7����"O�"P]���7n�'��l�6"O�������kzPMs����b��d"Ob��7l\�qv<D���<�<<2c"O����P5[��Y�!&�-d|�u�s"O�Q�F�E0�0ğ�gj*�1�"O�}���bg`��"�'<�@1"O"��$��)���خ#b���"O�$��*����5㕈�>�G"OztA�	[5�i��g�,i��):4"O����N/����AG̞3nX���"O����-����LRa1�0�3"OZ���PG=T��
�1Cr�(H7"O�٢4e�>RN��J�	K_X`'"O| W�U-��\H��<2���"O,X)�FT�%n���MP�{Ll�"O�0s�B�eG-�vkƓ#Q��R�"O��)sㄬ�X���
�N8��"O��C�J��Y�Xc�ށj"�$�"O
�:�cL9 �aB��F9�pT"O8������,��Ǡƫr�$�"O�	�N�
�݋6�"I�j1;g"O"����\56I�H/(e�����"O@% 2��NR�PЮ!G��0�6"Oh����>���dMS*=o
��"O� ���!G].9����N�H^�싄"O dqs	��W��<�d����؃�"O��p`��5�C�H&<��a�d"O���Ra]H� Qf�(� "O�#E��[��s�l1bG�Q�p"O�DF<�t��@�C5�LA�S"OF���Cؑ��a��P�Z�T1{�"O ���@�T�T�
R&~�T�$"O �5��4'���dS�3�4��b"O��9b� ����{���
E�@�"O(����I�C%,�����X�n�QD"O�ya����P�)4!� ���"OXջPC�7_�u`7b�]�|�1"O.�)���{I�`�"I�z�%b�"O8|X��B1�U(�'2Ԉ1�u"O�(����B�L��К0�Te�5"O ��U�&� iG�CԼ��&"O\�6"�(t�����%�14��e�s"O��1���di���DA�O��q&"O�9�ḣ'ک����K�ļ��"O��aleo.���BU�~�Dy�b"O���#���~x��҃S�n &a�"O�}���D"Z����!��e�� Z "O�qM%R_�R jT�v�*dk�"O4�"����dړ��­ �"O�|B��	~ς�@��Un&� %"O�@`F�2	�P\�7)�n��T��"O���2�R�C�t!(GaE�x�	c"O�ۧ)�n�{�m��q_����"Ozqg,^�Dо1[g�I�0NJ��@"O��R�6z`�"C1VZ��A"O�Ya�.N����(��ko0��"O�[�a]��Z��[�PN�) �"O"]NjG&��		C���C"O�3�J����lE$r4��"ORT�w)K���j����`�*�"O4�si��]���B��O�f1v=��"O�*�e�
R���p�O�����j"O��r#��9�F=��n\�,a6"O1�V����0����ZR��1"O��7�C�p�}ɕ��W��xAB"Oh���h�J�J���D�&��u"OE���Q|ȩ�lY���h�b"O,��ƎN/j�����Ϫ9���"O�S�NH�X�$�*��Ǜ��Pc
�'f��X�e��4��A�Z�z���' .��#y���7�P=U�����'$j%AjֈUPp�$̞�]/&���',Ա�>1�<J�P�Q��	�'~��	��f��bǮZ�I^`}��'E`�aDℽf�I`���:���'�f\�P#G}�hǀ�:�����'��q�`��t����%=+*M�
�'2���������테V��e)
�'��(A@ªv�n8��+_5Sd�=

�'���6�_G���CBN�1R����	�'�X!`v��~v��dC�N�B��'�¸{S+�S�l� B8F�D1A	�'R�1aG�~TI�u�
FN~]��'Bt�z  ���   �  C  �  �  �*  G6  �A  �M  JY  d  |o  �z  7�  ��  ��  $�  z�  �  l�  ��  ��  @�  ��  ��  X�  ��  �  e�  ��  R�  � $	 h � � b# ?* �4 e= �C 9L �T �[ �a 2h rl  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+a��6 \��	�<4�d5h��'�B�'���'	�'/�'�B�'��I2w��5Kk����e��U�D܃��'�b�'A��'���'}��'��'�>��5�\ h4tIR �>���'l��'��'���'2�'���'b�Iz�k�fVЂG�[�x.(���'���'/2�'��'"�'"�'�^�qs�S%V��c߁Lb>ıf�'��'@r�'���' ��'h��'J����b���@�3MTV<q�'�B�'�'���'���'^��'��`�$�͡9Ql�#[�=�"���?i��?����?!��?9���?A���?P�Σ9<�x�
�&�+K[�Jъ���O<���O��D�O����O���O��DLw�eȴ���ŢW�2(�'��O0��O���O"���O�d�O&���O,���ƏX���K�8�n͊���OP�$�O��D�O����O����Oz���OL,���0�"&�:3�f�j���O����OD���O����O����Or���Oؕ����JT�
�G�Oݨ��Ԣ�OT��OF�$�O���O����O����OH�0t�ʰ[O�XbQd|�^4�G��OP�d�O@�D�O����O���Lئ��iީ�ć/TF�U�ՁN�:�Z�34�ڂ����O��S�g~�h���%k�2�8�!#$>=�B��PX
`���*�M���y�' $HBR��,�O�o�b-��'�2P�&�����dΧ)����~�D��	[�\�2f$�*�B�Yé�]��?Q+On�}�2aX�n�<�ah��nY>jE��+�V�R?��'P���nzޑ�R��
ks8D贀E*b����!	ٟ��	�<��O1�XYل&mӐ�I�&]��T�c�>@�0`�n�L���<1��'��F{�O�bH_18���T��t���b���yr\�8$�x2޴n�>��<!�&	��TME�>`t�9r�����'�듰?���y*���Q�(��Bu�X80�̈́51�9����I��Z$Zch9�S�rhY��H"��^'*�L�"��>L�b��dyX�H�)��<�����m# +$:�!�PE�<�c�i|8�k�Ot=m�_��|2��-!����ӥW*;]S�#S�<���?��
�p��4���m>����L���  �U�v�KE�D�^�4���@*��<ͧ�?y���?q���?�2阊x�n�  iX�r���r�>��$����d%�Ty��'���A��:� #�B�%j��0j��n}�h{�4n����|��'��N� d@�܈#S)w!t�8p��/9�X��d���?!b�� v��n���ug.�dPy�&�1?�n䠢�ƅ~C �5�_YS2�'���'j�O����M�"��,�?�ELW�E����ɐ;d6���Q���<)��i^�O!�'Hb6M���:޴6����B�V|�0��%N05��\��O��M��'Ѱ�	��P�+y|yxc�:Z�B�OO����w}�
�	R�}`<�jФ�<]�"��'���'��'%b�'8�<��� +�� o�xAVDa��O���O`�mږGi.y�'N�7M6��O>��lK��E�H���0Í7r���'�n���M��'vk�Y�ٴ�y��'|�Q�d4TL��V'�dI��K:XTT�	O��	)�M�*O���O��d�O��Je��1�� �S"��h�O��d�<��i������')2�' 哿0�[0'���q�Z�	��M�I,�M��i�O�� �`��A��g��(i��=?56�h��3?�Izv�=?��������V��Ӽ�d��S�(�0�C (�4p� "�?����?���?�|j+O��n��^$�-X��O.?d@
�P¨�^By�lh���<
�OԈm�<$A,D�e�F��6$0�)F�$K��Kڴ����L��;Od�$�/37��x��K1��E/��r�g�Q�P������8P�Y�4����O,�D�O�$�O���|��ē�kԄB���M��@�'r���VP���'yB���'76=�
�CU����tψ�W>h�Y�Ɗ�E�B�'��O1�vHju�o��$�J���b�u�$�KSʁd ��ix��P'�'���''�7�<ͧ�?i�+$���uʃ�;��}�0
�;�?���?����$Ǧ5�Se�Py��'N	2�@`|�c��):��ع��d^}��'��d=�7�Jd3���Ea����f��.T��O��Fӆ���R���	]w�4h�I�j\B���=>�ɋ��7S�൰���3Rb�'���''�S>]�0"+:�J��<�2���r��@ܹ�<��� ��f�B�創�Mc��w����#���2�b��C�ӟd[^ ��'M�&f��|n~�HynZ�<y�2�^${���D���,_/lF�-��	ӳF��5ӂd!����=�����'��'b�'ޕ���σYe`�� Q�f{�1�RT��@ܴU�1�+O���,�әr��7�,b]S���=L���8�O`=lڕ�M���x�O����O�x��&�Z�ff����b�&��t�������c�O��iD���?	��<��i�I�eS Y�FgT�n���D�@�y����͟��	��i>��'�Z���5#wr*Cˌ��/�<(L�&T��yR�h���3*O*�t�JIl��r�@p��A@,:�,�#O;-�|��A)�����?����l���@~Rjk���=� B$ے�NG@�j��~���f2O����O����Ov��O��?%���]�?5���ShA$,| �D�F����ڟ0��4R����'�?	��i�'� } ��֓G�����_�)`.�鷟|�fӸDl���L����	�+���h��]{��`��Q�$�P�&�_?��K��Oʦ'�\".O����O��d�O@�Rkb�xR�_��B�(�O��ĭ<�ƻi!���V�'k�'��	?��U�����E �c��[�;���#�Iğ��Id�)�Q,?�d�+�L?Q���;��U�b��sc�x����TƆ�3�|�%�t�у��4��'hѾE���'uR�'����T�ߴHi:8�D����(-J�j�Ku�ʓ����y�?�X�$�	�Ne�ň��E���ܰE�3^��q��ٟ�'�ʦ���?�)��p���_i~R�9Z�N�scl��!4�]��鐟�yb_���I�,������	ȟ��OƆ$��@/��(���Q��y�io�؜r�e�O����O������Iܦ�]�m�S��Ȋ_26�P��R��.T�� �Io�����pB�nq�:�ɎJ����"V�>��ysďw�0��+<�b��S�'N��%���'r��'a�	"��I$4|r�gO	O`((��'Wb9���'m2W�ȳ[wUzqz�V�T������Ar�oVJ8��S�h& �?�0]�R�4X��x�K�2�X�{��7��09�e3�yr�'��xsnͳBAf�gT����>7�¬�ßP1�ɖ�z�jӡ�Q	i� e&RП��I��(�I՟�E�4�'�Hȑ&��@0X��"MF'���K��'�,7��_Y��d�O��l�r�ӼCG�M#nF,�G*  D�u[��D�<�@�i9L��h��5ey��F�t��a��4���G1!zD�*'N>(�3�?�䓎�$�OH���O����O>�D$/�,Y`�+V0[�V�h�꓊7��t��61W���'�R�Ʌ�d�����Z#|���0����ؐ�'V��'ɧ���'B�EJ�Ҥ`GG�1T��!��$�Q��imx�&�8xHP ���%�0�'0��bJ1|��EIW01A�@�P�'�b�'�2���t^��ڴ-DrH���_6�8�	�-�D�R��ۗ=�������M|}��';�w4��I�� r�qIdm;0��8��Z�PV6O�d�pVv�s�O��	�?����Fu82l'Kp�<��ɫ>)��	ǟ��I��`�������t�''_��r�)~O�m�#�IF�c*O��� ¦���?�մi�'��(eI��qD��(B��$Nې�|B�'�B�'H��0w�i����O^͛R���G>��a!��&
\�A�T�lR����O���|����?q�yfr�i3!P�`~h9��L�5�����?i,O�ToZ�]��`�������?��ӊ��pr&��i��Tٷ�X�_��N��I矬�	f�i>	���_�<�ȶ���x,��Ƀ�7�J��e�C"yv�x� �"?���L���υ���Q���ؑD�>X��k��a���?���?��S�'��d�ʦ�Ʈ
3���@ů�J�H�@�M�<僧�	̟���4��'=(�8{����	/�m���=�z%t��2�7M��y������?Y�n¿y}��ɘ���D�h���xǃ�6��<C�gX��<����?����?���?9+�P��p 4>��}j��� @q.X�`%����]��h�	ǟ�$?a�I�M�;`��$�}R�]k��Й=�>� 1�iR��*�4���	���t���k�p�	�L�l��"��;6��7 ��<����7��풓�'�%���'F��'w2�B�+�QNa�f��%��T�'���'w�[���4 ���+Ot��6��D�V���aN��SD΢!#���H�OLnZ-�?�O<�"i،T�)%㟩o�����c~J�SGx���#ƨ�O\r��	�PR��UD��7&�9�2}Ɂ�O��B�'B�'���S�����e��ni�׆P�0�<B�%������&
��'��7m%�i�M�#.��i�e�fE�<A�(��G{���������:B�>�n�<���z��)�B���%�G,�A #$�B�0J�]���1����4�t�D�O����O����dj�h)���Ȭ�Gڛi���v����8�"�'z���'>ƭ�6+ �������T�x��E��'�>���i�L7MRt�i>����?�Zr�a�^!���N�����HV�8@,���%?!%��,
r��䘋����I�<D]��@9T�B�8�`Q#����OX���O��4�.˓'�e\(H�L�1fh d��aŴY\���C��B`�8��+�d@}�'o�"`�	�]ZV����}�2-�	]>|�`đ,`�nZ�<y���p�L㟔��.O�i��TD��GSf�#��_�=��B�3Ox���O����O���O��?�rz�HBF�"j�4��&B៰�I�Pcߴ,�@̧�?���i��'�*1�Ǹ^�N�jC\= ��阷!1�$|�,�o��?m�E���Γ�?��hE�,�d��B��K��x��9�"`#2��O`��N>*O���O.���O�� sj̻V `a��"��B������O����<9ŷi�8�1�'�"�'�哲:'lIц
�N��r{�h�1��	����	v����)޼b�@��T�&V������x���kr)�VĦ`�qͲ<a��q2F�Dǵ�'�
MPa��$�����ɑ��0[���?���?!�Ş��DW������P�r�y ,]صA�!,������$�K�O���'�6mM�9��ta�cĵ~��U:��)[���nZ��MքG��Mk�'�"��%:���S;��� ��a��k_��B� ���0:O��?Q���?!��?�����<tD�Ӂ�>R�H}��lF�g}�,o��P8��I���	D�s��9���cЗ R����d�1qj��� kF �lj�(5%����?�S%e}��lZ�<aQMʉ#t�0�m�7)�����
�<1"�.ؘ���!�䓯�4� �D��1��KBK�c�0`�p�@d�p�d�O����O>�A���#w&��'���E��F��vi�%j�8���BN�h��O���'dr�'��'_t���׬hOfӒ+!"r���'C2f%-,N�P�eY���$�z�*�����d 8��͑'�(R���4�Ѐ\�����O��d�Oz�d2ڧ�?��CNu�<��� ��4�C�9�?�u�i��*Q�'R�g�f��ݜyB��w�
�P0�[U�T�B]X��P�	�<��Ц	�u���(B_����{��@x�Ye\Z7;,��Oʓ�?����?����?��G�*�Sv��>[�<9Ҍʞk^-.Oޥl�8x}�L�����l�S��b��]5�)я�;
Q�Q�����O ��(�4�����O2� �g��k:0\2vh� X0@4a��K=Xd6mTy2��wU��������$^�cR���
�36��h�r��]L��d�Ol�d�O�4�$�	"��"ʤ&���Ҟ����`�Q�g����&�Ѐx��m���(j�O��D�O�NG��tHG-�.8�Di�kœL��vHkӪ�I��xr�_�*��)�<������h�'0N��� �^=�x����<q��?9��?���?���Z4{ F�rK� ;H�9�g,*�B�'���{����V�<��i�'����7e�W�l=jt�ب��*a��'wd7�V�M���w��io�<���g���{3��h��LA���$a
.wGXՁ6�'n��%�ؕ����'��'�.���X�9$�D�  X(r&�(��'[�W��X�4$������?I�����"��q���7U��;7�������������Z�4dމ��)�=L*%ppL:T���eK�&}H��d�!��Q����,E���Z��4@%�9��%6�ε�U�U$T/��I���I⟈�)��oy�w�xL���5pkȨ�����NiK�@��4ʓ =�V�d�O}B�'��ĸe��i��	�fl�(W�*�Q��'���V��2O��^��vA;�'T��	�b)8!_OY���q"��M�v�	By��' ��'�'�"P>�g��N4���:c�����`�Ms��?I��?AJ~����w��"�#�$(V02B-i:
D��']"�|�Oo��'� �aǰi#�D\"y�`AQ'��y�H@�ꜷ8��D]2�L����̓O���|�����|;��&/�`x�"/V�0J��?Q��?�,ORl��{h�	��	%*Ol,��DψGҵ�)ԅ,�`�?�S����П�$���'���_���@�1��ِ�x�\�	Q�Qj3'R yԊ�����O���$�,�*����
�H[b�V�*T����?Q��?����h���$ 
�d���YU���H��&u��DŦ!��V]y2I`����$uF,z3��!!�>���"J�x�<��
�M{3�i��7�[0Ed46Mt���	�n�� ���OF"p$N�;g�4�Ђ�+m�"�ëa�	ky�O��'���'��.]/F���lE!y�ǫ��I��Mk�m���?���?N~�0G��Xs"��~�z�B�:x	neQT�tk�49���o!�4������]k�⍡'����U�&��b��3��*"��d1uE�g�D�@��IyrFY֌��.�!�x%"V�(1A�'���'U�O��	(�M�����?��	W�8	.�9C�~ �	�#*�<���id�O�$�'#�i�<7��<w�qy��E;$֨�PI�L�l���b}Ӱ��ϟ<C#@U�^~�T*;?Q�'ƿKu���y�`�uH�f&�����<q��?���?����?!��!�%R��Ax&��g�D��N����'��Ns�vtk��<E�i��'KҘku�\�0M��j�*L4EM���d-��	ئ�j��?���ݦ��'OҸiEi��p��S�7����sf*@��$��+9��'��I��T�	ȟp��!
^����ʟyI$\���4K*����'�l6-̬.�L���O��ĺ|:��S�Ҡ��QoH�pP�UyGƖ[~b�>y`�ig6�:�?m2A�>7()���Q�BY:EB��'<Jղ�B�[�4����jBȟ�{@�|"NI�7�}��-�M~�����Y���'�2�'8��$P���4yk�ԁab�{��4R,�#Y�� p6��?����$p}�&x�|\�qŗ?!w�Љ�.~ׂ�c��V����ߴa�T�#�4�y��'��)��$��?ͻ�X�h��,�{��p�cZ!����2�~��'�r�'���'�'�y+l����]%���@^�: ��Q޴I,D�����?������<�w��yG㕾Ȏs���(A>h���	���'�ɧ�$�'��oVX��;OX���@�Xx�����V�
�Y�2O�
����?9� ���<�'�?9��P�H��X 3m�����̀�?i���?1�����˦�⁬�����	��p�H^�s�@ؚ��T:^^m���f��l��I����z�ɠ5�$M@�[�9q�Ar�7b��	ן(��!Q��ڄoڿ��$��)��'��kN6:(�Q�#s3X8Pg9y���'i��'Ib�sޅi҅��O��p���3��A��oڟ�8�4Rl��+OF<m�I�Ӽ#�K(&|ࣔ�L4 �c"�V�<����?	��0j�]"�4�yBџ��2��?� �]�@�~�T��ه�$��l7�$�<����?9��?���?ɠ�M�FH���J�:(Ov��'�0���妡�#!N����	���:�h_2N��d�S�_�BX�ޡR�����|�	`�i>U���xz���4h�+�	�o�����%Ա,��HnZ��d��aY�'��'��I�
����i6rx�E�*Q�p��؟��	����i>)�'�r7m:NL�D�6B�Ёi�טo�<���E�nK0�$�ئ��?V����4G؛){�J�1��D.@��	i�ɛ5"�DE�#��_�6M#?9�s�I1���A�Ȉ�^�f�ZiX�X7E�y2�'�'
��'���i��>&��YE
�1H�@ؠ�Y��O��d�O�)o-n4��'R�7M>��I�q��y``�J*g�h�6�� ��&����4!��OҬ��S�i����O����Ei�f�3' ۰zs|S�	MC�j��v��Ob��|R��?)�] (�3�5.�hE�)R�c��?a*O�m)D�Y��ҟ���J���Y? ڞ];#�  �"������d�j}�+|Ӵ9�Is�i>y��R&�9�H5b�J��!iS�	$ԩ*媁�`=�A"V�Xy��O����2)�'�<��D��Kuf�9A+5\���R��'rb�'����O���0�MK�W6}�p)^I�hTނ7"���O�������?�bP��;�4ilؑ�d�W7���ApK��{�R�Ӷi�(6툶E~�6mu����%
7����O}T��'���[&�aK�x����
7*���'��I�x�����	ן4�IO��L���X�P��+0.h����	Y��6�
��D�O���9�	�O2Tlz�E��Y�2��@���֔�D�R�M��'���t�O���dK�#�F1O�X	� �;R*��H� �'Y�!�1Oj�c�"��?	�E4���<��?�ǂʔ"ᤤa�bN:[4ACl���?	���?�����G��咠̟����\�3K,P�p���\)qrr�Z�́T��~��	̟���i�aش����Y&.�A �i�)��	�X�d\&p\l� ����&�K�'�"c��D�b����R��rŦ]eR�'D��'I��͟TG��3yJ$�3$ą=t���b��XR޴DMԀ���?�4�i��O��̆?���O.e�����DO2p��=Γ�?���?��Z��M��'���B�w���SrjXdk�N��w��|����%>�q$�h�'�'�"�'�R�' ]����U�E�ȕ�:^u#T�PIߴ{�N�I��?	����O��p���,\5J(�ā�+1�R|ӂ��>���?�O>ͧ�?��_���S�&Y�̒3��14�J���M۠_�����'�d6�Ĩ<9R
\:9f�AH@�=�h������?���?y��?ͧ����妑�n]џ����4_�2�c�2�V��|�t��4��'�|��?���?�f3"S4��]�N�=���^��sش�y2�'���F)��?A �OF�I��AZ����"�����!D�_|� =O��O��$�O��D�O�?�Y�L]T��h�/�.!��I��!ݟ���̟���4ud�`�+O��m�x��^*��k���Z(q
��-G||$����ԟ���"4�$�n��<�����0�"0j��<�nO!*<�Ŋ �!
(��$̓����4���D�O^�D���ӀF "�({�gw���D�OD�$���G�r�'�V>AS�l�Ӧȸ�"E.ȨԨ&?�S[�H�	ܟ�&��n!nlR@�V)-x�8�3�%���&<�.���'�C~�On�I�ɘ|�'�-��O�[7�9�'/�?'�ؐ��'���'�2�O�剖�M5�����/�8r̍yEIܲ}n���)OTml�i�t��֟�J1A��r�0}C3�O>^�^��!Lğ�I�"��n�k~B��5L�Ҙ�St�IS8�$%�"�{T���a�t���<Y���?q��?Y���?y*��L��CI"w�@�)��)<�	���ꦉ����؟8���8%?�	��MϻP��\*��س�ꬋ(Ԁ*��	���?yH>�'�?��=��u�ش�yR�45����P���"���c��A�y"i���	;f��'��i>A�ɑ4���{���w�\�p�Cś��E�����	�'�n6�_,z/�$�O4�dM�(��sW"M<�h� T%U���$)�D�e}��x� )n2�ēHS���M�O$�у@�����̓�?�E��*�p� -m~B�ON����8Z����7?4z�ˇ͜Z}Ip�N:�'���'���ß�P	�1�$���+!dL��!^ʟX�ڴ��k-O��n�W�Ӽ�aL�A� �rR��nfZ�b�nS�<��i�H7�٦��\ئ��'���PU��?��Cg�'rY�4I���)p�%��_u�'�i>���|��ҟ��I�(��4`ѩ+��k�N�H�2 �'��6�ΤD�N���O��������<�Dm������.�*�\�Hை�h������nZ ���?q�S�?�6��A~ K�c\e���_�H����7?q�iE�m���$�������8b*�b�&őn-ب������D�O~���Ol�4��қ�j��z�r ���場�Ǔp8���6�y��~��⟰��O�yl��M{#�i�\T"���8���jÞFd<�A�N?��?O����|�൐�'4p�I�?��]B6��aף�^VP�qG�?���Iݟ��	����Iן���X�'U1� ���&8�7a��J��?���:���"�Z����M�K>�%�A=y�H:�K4�� � -[��'��7-Pæ瓝}2T�np~�K���� �������RݡPɂ��|CRJ�)�?��	5�$�<ͧ�?���?�c�X���	�D&s� �p�?���?i�_��|R��Y��?�+��!oz>�a�!��c^~x��摴��!�G�4?�T_����4!N�&�8�4����3o����F��+��N��J��0+�Ô:��p����� (r��P^�80�j���(����q��∙4Ӛ������I��)�by�k���r��]R���ɭ%�SDG�&ʓ��V���m}��c�6����q�	�'(��T<L��I�	�شr�X���4�y��'�4,���P�?��`U�4�ś�=� � '~b����$r��'���'ER�'N��'a�S�YB�\bu���
� �G4&�B���}"@����	Ɵ%?�I��M�;=: �Qt�ܛ_�T�i�,��?ިЄ�ij��$4�4���i����� e��	j� �q0oϣr������Ρm/���{�H'�'�8'�X�'�r�'8��C���#�\{��J�$�k��'�B�'��Z��s�4p	��3���?���K��ڔρEy�V�"A�T��2�3�	���d�����ē�P�s2�ʵH@���T�B�8Mϓ�?��9>��Fj����d�����NR��MVc��IM%I|�!ys�[�q����O��$�O��.�缓�Ɉ?zD�᠕2���8g���?�r�i@f��'�ooӴ��]�i�00�vɿ{������+1L�	�����x��K��eΓ���_+3��B�dI�'��%c[�0�b (H���O���?��?A���?a��]q�Ѡ��;:���&)$j.M9-OZtoZ�W�"	������]��$� Aߟv��)fc�$��2�ɂ����O@�$0�4�\���O�1�dj�	#B�i�������I���0��7MTzy��͙Dh
���䓵���v׊��6L�dm�MS�����N��O|�$�O��4��x��Q�����,�r�3.^��!���)P�Rlg����)O���g�l��&��+Ck�	Jёe-G�>w.U��O�)Γ�?Yևݥ=N(���B~��Oa�&�D�&U2Ft���aC��y��'+"�'TB�'�R��'���k�]�������(�$�O��D����:c�}>��I �M�M>���X��J�(T�s�d�2�+�3z\�'g�7���/l�r�nk~���l��4	�";{�MIB̯}wB���ҟ ���|"X��ڟ����)vn��Gh��%��-��*BJԟ\��dy��o�rm���O.���OD�'��9:��H'k=��4Bų�8��'�~�C��f�p�9%���?���� *f�SEd�"euv�dę�=�z���'UN���@��O�YL>Ԉ�P�P�ޑca���BW1�?���?A��?�|�/O��n��`�4\R�Ά>b�AC���X2Kקw(��O�mS��&h���MK�"�Nxɫ0d�p.��D�0M(�F�i�xMl�D�I�`rB ���i4?ѣ�^����@��m�$PK��<1(O����OL�D�O����O��'�V<��τ�?n^�IK  XXE�2�i<�=���'m��'�Y>����Mϻ&e��ۗ)Ĕ<w0e����`ъ�k���?�K>�'�?�L ���4�yb�Ę>�|��e��!Gdq1�J �yr�G�\�(��������Of��^NR��]� PLx�� /n�^�d�Oj�d�O��I|�n�(�'���O�qΌ̡�텈iGjĻ��D�F�Oz��'���'D�'^@e0��1�����0�p�'����q�~H@�io,��B���|��\�&h�#✥=i����#k3� �	����I؟��IZ�O1��vV��37�M͖mh2�F�(Gb�y�V�H�)�Ob�ā�=�?ͻd*Z�kÇ"��I��hw��̓2��fq�hn.��n��<���$�@&���D�sV,�>O3j!��)VzLMp��Ԍ������OX�D�O4���Oh���F�(|b# �5�* ዟo!�ʓ8�V��[��'Ғ��'0�u�2@N�w�Ӆ�ľv�v��#ǻ>)��i�H�$7�4��������a�#��&Q[p$�g�^��L�n`�,Aq�<Y���kQ����)����5Ct��)�� ��8��:�z���O*���O\�4���r�&�ܝX�r*��6H�oL�(�+���j�*�g�F���F}b�s�VL�����h�J�.
�d�o
2m�8m0瀕�Q��aor~���!V(Ѕ�S�$��O4&�J�|�A񉅯� ��D���yR�'���'��'�2�iK�xx�Ze%V�yD��zd/�Uw��d�Op����E� ��Vy2�a��O*%kN�/�ؒq�B
�͂��2���O��d�O*M��JmӬ�Ix��%�\)3pgG[#b�I��FT��I�'r�'���ܟ���˟D�	�'�*���A/1�"h�(N%x����۟�'̐7-
:�����O���|��	����h�dG6ѡ-�M~"g�<���?!H>�S�?щ&`R&1`������k\����ƍh�&}���0X6�x�'3�4,Nɟ��r�|%
�U�b|�ae��N�p��b��2�'x�'J���X� H۴Iq�ٛ��T��|�CcÔd��dٽ�?Y��42�F�dL}2�'�ʇCA]�
�A �2/�La��'⧒*a�F>O���]������թ��"I�2��Л��X��y[�X���`������	����O�X�Z���C����ˍ<\��5kҌr�X)xg��Ox�d�O"�)�|�]�wtrp�"�[�~�Qc�8Z�$qxAcg�֬m�����|����:&�A��Ms��� ��[�b�8<�DSU�o��̂�<O�7B�i�BM�Z�	^y�O�ү��8���ZZr-"��ׅu���'2�'�I0�MӅkD-�?����?��*)h`���
�ehCh�7��'!�9j�F�q�j�%�䡡�
�-�X�w�{"0�k�8��)}�<�Y�.����OF����?���Ov!B��ߙK�<H�B�j�P�{�&�O��D�O�D�OH�}��/�\x�g�,�D�O�d�R����H���E���'�7M�O�O�|���EAāoq��`�fSMJ��P��*ش"6��M� _�0O�����KiI���y��-�Bg�`�2�h�fTMr�)f�<�$�<�'�?��?��?��)6"д�o�1Vz�B�����d[�	YdϔRy�'���`[ҧU)M'���a�ު?G֭�%ʄv}�'5�|�O�b�'jq���S�O�x�/�=B#�P�>��O��4f���?i�#�Ġ<��S�"#xI�����+�D��?i��?���?ͧ���	ɦy�3���4� E<!��a�D���q��o�ӟ��4��'����?��Ӽ�THT ^��XQ��e��M[�k�)LP8ܰ޴�y�'r�0�h-O$����T�+s�P�v�8�{��ݑ;��d:�7O���O����O8���OT�?m�Uj�G�X�&�);.�	�����������sڴSKf��.O�Io�����'��Z�AV�f�ʤ�D�1u�\�u�|B�'���'8P{E�i�?�[t��2���(
I��A�"�7 ͊H��������O����O��׶TIS�c�`Ӥ�S9�a{���?y)O�lڈr6*<��ʟL�IK�t��K���gN�i���(p��-���Z}r�'�r�|�ORj�"�LԱ��#X���zfB*^�fy*�4oA�#�<�'��	p�
J<�ݺD��?6:$B"hT"9^��I�������,�)�ey2�u���HW(4���\�� �6�	�b���O��lZ��C ��3�M�C�ц���8��${���E�^�_��֠~��p�1ks���΅� 埒�O�PU���0Z�����*�)6��"�'����D�������0�I^�D�NMH�
S�թ&}X;���58��7-Ġ]`����O��$2�9O<oz�]pP���& �ǧHk��"��M{!�'����O����iA�d�uXL+3.WΈ��Ś�	��D��v�H�	��WX>�O@��?���4xL�y�ِzh:�$���Yj�4:���?����?�/O��oچg���I����I;�l�ah%Y�*L/�l���?�]���I�&�`�6Y�H@$��� ���{d�`� �I�H�rb�G�A�'m���ʟ�"��'h�-�t^�)��FC�}�T-���'���''��'&�>���vp�yv��*VM�u%�_Ξq�	��M3$���?A��
�6�4��a�թ�V���o\,���"2O��n��M�7�i�ؑ+b�i��d�O��r%����!�^�`V�߼eI�oޚz �O���?����?q���?���ho9��'l� 0k�
#4Ԥ�,O�nZ�:��I埴��w�s���P/�&c��Ĭ֡������O/����O��>�4�Z�D�OD-r�`�)�(%�fcPt���t�W�lrԀ�"��9���*V�2EHe�Ijy������sB#D+��pV�
-L��'q��'��O��I�?Y6fKן��ׅ�'��I*#g��!�f�ʴ�i�@�ٴ��'�x��?����?���+ei&A˃☉X�l��O�:����ݴ�y��'���q��?e��O����lXjd�ϑc[@���t��j�2O��d�O4��O���O��?��A'\����wK!	�p��&�ޟ`����h�4N
�@̧�?Iտi��'����ND[�5�l,,�,� �|��'Ib�'�H�҅�i��?rKU7mk.�P����vW�E�ĝ�v�V}�����$�O���O0�$ԛ\��i��)
�Rm�Ö�!���d�O6˓w�K��I��'��[>�1a�C�
%�0M�xp���W+#?Y4Q���	���%��ȟ�{�I4S��T2�i�:Xd�0�$��w�T\�A�B8S�t��2�#�O0�ZO>�C- �c��1$iC�Dp����ӿ�?����?��?�|*(OZ�o�a�,����{i��k�m��EH�)���ß�ɪ�Mۊ���>Q��?d<����}!g�@AB�j���?�4$���M˜'�	���ry ݰN��<b�A_�%��� -�=�y�X�@�I��P���4��˟�Oy��9�$U"R娽,J@�O͎F �6M%P�����O���/�9Op�mz��1V A[S�p`�-�b�Af��͟4��G�i>Y��ϟT��VƦ��~w�a`thL�}bĉ��$��D\�5̓G���7�� '�З'���'bf(!pb�/-��@��'4E ���'w�'(2T����4N�Ta��?Q��{�590�I�BNR|�!����E����&��I��0�	l�@r�r�h�bѐԣݢ_'B����8��#�P%�����Qy��OJ���	�#LV��͸�!EznZ5N��}��'^B�'�b��Ο$�T�+41�EB ET%4:$�@%�П؃ڴ~�������?Y��i��O�N�+5��w+�=f�X�!�C�7��ަ�K�46�V���F;OB��	\r�',5(�{bdA�@��%XS^�꒮;�$�<����?���?	��?AG�Ԃ1`�����:��������DŦ!�s��EyB�'9�O�r�	�_��P`��B(u��l�w�[����&�OO1��y[r� ���E�.+�j�CA@ƈ~舜�@@�)���#��"��O�l[I>�*O����oZ�W��ġ�[�M�>H�f.�O��$�O��d�O�	�<��i�X�;�'��]hS���q�E��.;(�aV�'��6�5�	�����O��4��Ѳ���WBl��󣍿Ef���>4'86m8?��:v�(����ߩ S�����Hr�$Ed�ڝ
u�n�,���X���$��ߟ���֥#0F)�@MW�w�0��A���?���?��i��0]�H��4�� HleC�Kэr|8���/�9$��mJ>���?ͧ-�X��ܴ����ek����W�E�f� hg0���ِs����z�xy��'���'��#�"](�(��+9Tn���(ǘ��':�ɵ�M�qkL��?����?i,�����Nj�Y�c�_�H�
���8��O��d�Ol�O�S�L�8�DJ�]CbxêQ�Q��(ʴ�S5�zdn���4��e��'�'v�� p���]5~@
�D�����'���'�2���O��ɋ�M��NAK��x��n]?C����"�9g�� �,O�an�V��F�����MK���$@,�ѫVf����'��t���e�V�i�b�F.��cf�����O���� ��;X(���+	AI�'�	�p�I��x�Işt�	C�t�8y�ڴC��JA�xb'#W�_�7�D���D�Or�d6�	�O���w��la��D�DD�-8�r����5dl�Иl��S�'p>���4�y���s?�ap��T�oFE�g@I��y��� 'SL9��&x�'P�i>y�	?�.�Qǭ�B�y�Sa�4Y^���ٟ��	��h�'?�7m�62����O���KG [ӳ��� ���yw����O��nZ'�M@�xBd�(����LۦB���i��y��'�(ď[4���A�O����7�?���OdQ:�-��e&DI�E �0��]����O����O@�D�O$�}��� %�-)T�_�&VT8Ҥ
�F`Uk�hM�V�
E�ɀ�M��w����'� Mjjd�� ނ;H%1�'22�',"�ۻ<��7O��d�-1^�b����yȳ����N�)a���8!��>���<ͧ�?1���?��?9�ួ�*q�`���Sm՗���Ӧ����ޟ��ȟ�$?牫� ��qFT*�:�2*�}�ΰ[�O���O�O���O���K�~mh�ݼz��a�''Z�f��X��ǆ��ɴ@�*!�d�'إ'�4�'�|A�Y�}$ �U��I�Z@��v���
B�K�B�v����
&rtq�b�"��m���hr�O��$�OB�D�~)��T�5>����G��2�TI�$a�^���Ȩs��?�'?��ݑcq�h�J
+�\ +C������@�� ��
�Q�DQ.W���2�ӟX�	ҟ��ܴDf�4�OP6<���B$���^I�H�
�U�̓O���O��6��6m!?��u$���ȑ!v�𪱧ԦCm��G`ڎ�~�|b]�|�?A��A �Q!T
�����S�';�6�(KG�$�O:�d�|�bL*�bᱶ�H�(��e�R~B)�>	���?�J>�OPX=�tb!J�p]P�m]0��1�U8J<�!J��i+&��|�QN��h'�t�B>��"bL�21�"L�o#���4a㐔�+U5�P(��Ȅm. <��-��?A�w)�����J}��'��P�V��jh�r�(�7|n؊'�'�J΅����֝�jj��'��D	h��];S*R�6gJ(���U��ľ<!	�q`�3tė�h�b�/(>� \ۅ�i��\���'nR�'��|�nz�a�D�<���jFG3*��PE�Ɵ�In�)�8-�(�nZ�<y�+��uxk#�8w����EO�<!QG��3Cj��|�Xy"_�����t�N@�6��z4Q�N>OL@ow��}��՟4�I9�be�H�2b
< �b�@ޑ�?)!X�d���0$�p�A!\�������6���d�)?)rA��p38Uy�4g�O�dx���?1cC4[X`)��nP=��(3l�p�<��G �_xd�ie��5~8h��-]�?9�i��&�'P2Io����]-+����g)�PM����+�j�	ҟ��Iݟ���JϦA�u'�A���iїX�UC �ܥ��d�����O�ʓ��O�y��a�0��]��Ć�n i�ǟ�dz�4'� ���?Q����O�%�U�Z&;���r&b��0K�>���?�H>�|����<m�=�Ĉ�w��R��	�~&����44�I7!��;q�O��O�˓,�X��VNU(:�X��J��o�F����M;uH���?iu�Ȇw=0�3�!�\���
�	��?!��i�O���'8�'�B�ߚk� 4���)/d��gNB�f|Pw�i��ɟ9-��֟����əG� 5�",�Q��:T�$2�OB��A��t�E��-L��ꗤ�O���O(=n�<KԐ�'_�V�|���wI�k̨&J�����'F�����)^0�ƚ�֝�wA����P)f�e��@+x_�Q!�YA?�N>q*O��H�ߌY�,�ӠIL�1[h}!�5����b��~7��'l�U>e��.��hd �a	� l��8� ?&S�$�I���%��g�? �Ȇw�h�����$8�*a�V�P>����g�PQ����N�v?�N>i�crѺ:PD�U�0k$d�P<�D�i�ig��#%O̔*��&��D�6�ݜq���'��7�5��!��d�Oΰؔ�_�[�A�O_5P�x́f��O��M��6%?��l�E	�Ot�n�� �I��h휝Sh]	(�d�I@yb�'aB�'EB�'��P>5�$A\���)֧1�e�����M��
U��?��?!H~��m���w�<H�Iڽ\����bA.5�L�[7`�r@�	Y�)擶T�X,m��<6�#��ɻ�*�,� �r���<q�J�<e����ý����D�O�$��*#Hl{#N�SrR=I�GM����O����O,ʓ����9��'Qrl��~��Am�/�b|�  S1R��O�l�'>�7�R̟�$����J,*�FMI'J
�Π�4�4?��N�% �9�K	��' >�dJ��?��A�a�X�Hr'�f،��q% .�?q��?	��?��	�O`8���.��a�4o����(�O4nڌ x6��I���a�4���yW�T_�j9��BŪ�N����C0�y��'K��'�.�0Q�i?�i��r��pRV�'CW���u@�$���)U�����D�O����O���O��$�IW���tAΥ5Հ8c��ٿ��ʓ���^m���'O�����'�Y(�̩I �͋&�_K�a���>��?AJ>�|Z %�:V�8���%�,6�,c�E��p%���4{P��+.,�#1�O2�O��p��`$L#x'��0�E�$_���ɧ�M3&d��?�A�)I��,�#�W� �c��ز�?Ɇ�i}�O6i�'���'pr�ͅo#n�J�	A4I��0g�!'$�x��i��I�f��sSџ�����n�<�$�#��j�A�ԬŸ,3�d"�O�T� n�Q�"�	r��Gǐ����O"��Oz�l�
5�)}�ƛ|� ��Z��=ůDv;�h�����'[����9o�֖���Z�,KcZ�%���QBcI�V>A��p?�O>Y.O��іF9o�`��<�z�q��#����������u�4���&��k�J�`%<��A�Þ�	�����O��$)��?�a��+E��se�{�\Y0���&&<a�R�Hۦ��+O�I��~�|bGQ1��,��d��A?��(^��x�Bv� �B��_2H��)�@ ZE0f� 6 _�`����O4=l�L�l�	ޟ�I�*���ҋ��p�i��F ����Ɇ ���m�^~Zw��9��۟$ʓE��E�;EXl��&�ے�����O����O����O��D�|��� [>NI)�@1a���焰e���g�)G�'-���'c�6=���0�(�	�"}a�+_�Vt�!�L�OR��2����%dX6�i�$��ɂ	/tz�	T�`}}���z����DG$7�r��G��dy�O ��%`���䝨C�H�T,��`��'��'��I�M�#���?���?�DH��]<� hfiz���T����'�Nꓝ?i���}�}�7���3�~���1��d�'et�S�m�:p�������L�������'Avr	�9�ҙ�"�g�2����'���'p�'�>�	�9�l�xrBn�M�MK&�8�	��M�1�^����Aܦ��?ͻa���b@Ҋ0�ΝRr"6����?	��?��DZ��M��O����������J`Y"��}�,@��C�/jΒO(��|����?����?y��{\�,A��-���Ճ�d�`�y-O�Tl�;pt(��럼��C�s���6�L�:Κpڴ��t<+ `
�����O~�d9���P#^a��q*�w#N�⁚�)0i���&��5]R8��'7L@%�0�'�Z���@�h���P���\r��A�'r�'�����T����48�~$��m�ޙs�)�6@Ap*Ύ	q�p����D�f}��'���'���ǮO�R�
����]r������Zv�F�����*q��4���窱���e����b�JP�:OR��O���O�$�O��?��7eA24;K�Ɯ�(�0f��8�I�HشAz�-OW������+ƶX˺%��!�F���I>����?ͧl�>�S�4���F�Dr�$ |0�J"'@W[h�ɰ�9�?�G 3���<ͧ�?I���?��
��`a�G�ۗ^��`�H ��?����Z��3-�ݟ��I�8�O��s1��`��Xh�%	?."���OvY�'�2�'�ɧ��'�lX�R�@�Y y����n����6G2��5���i2kRC�I�z�r���Q�l�<[�iK�R��I��ޟ(�	�� �)��`y¨y�D=;3A@6J�ʰ����!ᬼ�eF� ʓ1f�F�$Y}"�'�,u҉ɽ{(�4Q�n|���'��oޤjp�6��lbr��8H�$�~�U��#S���3!k@�f>a$��
hP�kFm�8�>d�`P>� ����x�|s�iE�z,N񡥂�|3 )��柚O�p��	]9&�&X �*�,&Xd��6����2� f�J�h×
P,��Qb*Z�=�L���	;+�-��Fܢ]c`�f*����O������0��� P.�dK@�Fޕ�@�m0�hU	D�#�*�[QU�X�:{�a(C�a��Ô��*E��/q���/M�1Z�B���B�H���1f!r���<�� �W�z�B	@�@Fo1�RԪ9��-�U�?��\iDKq����O����$�>s І6($�CJГ(����p.�?�����K���֟`A	� ���rlK���2��UK�2m���i`r�'�b��0-[�O���O���
(z.%��ą c��(K�+�-U�c�X:��;�	����I�����˗q޼�j�^V��5�Ď��M���`�(ԫ��x��'AR�|ZcJ�	�/ն>#��[���w���b�O���B��O��D�O��q�~������f�։��$�P�:�!��)܉'���'r�'��	!Ȱ�E �
�8���#�;R����@&������ǟl�'����r>�����:-�R��w���2k��>����?YJ>�,Oj�iX�xx���
I'Ǒ'  �h��ʧ>���?�����u�45&>!õ#N�E��dj2�ͫ+[�MrS"Z�M��������1>a�O^���A�bdX�c�1W��X�i���'
�I'jWјH|2���������Ȗ3!��R1
�&��S���'��l;ȟ�i>7�[(Z�l.e�����뺩�ڴ�����T�lZ&����O��I�K~,�5A��,�O#_��I�'��=�M�.O�ё3�)�� �D��6(N�H�Z�`��A+�7�ЍHպ(n��$��˟��S����?i%�E�P��T�у/�$U8�Ξ�`ܛf�O>��	%`�̀s�XmR@��n�.~H���4�?a��?�aoE	[��O`�Ĳ�4X�,� R�D�BC��� �7�I�whb���	�X�	�/LN��Q�� $ŚYB��NjH���ݴ�?�73/+�'�2�'~ɧ56�D:"U;��=h�mz�G�%��O��D�O��D�<i��\Y�3H���[��X�Jqƛx��'0�|��>�ʅ���p���E�5(ɀRBDm��?���?Q+O.�zUB��|�%�R�$	�T����hR�t�")���M�'��|r�'B�G�^n��@�fθ�BeAA="��Z4��	�d��̟Ԕ'00��&�~��f����&ƛdJY�d�\ p!��i���|R�'��hP�/qO�I�@�O��x����l����Ӿi_��'��	�1�ݻ��~��O�����HB��!3>\����4 ��x'�x�I��U.�U������cB.��o���E�뜻�M{(O<	"����������?}ȬOk�*1�� h��+؄��ӧ	(Л6�'�L�!txR�|B��D
U�qe�#W���S(J6Ǜ��J��6��O����Op���U}V��R�G�	��i��=:Q�����M���
%�?J>)����'x�y�"�;��u��A�[%<�z��a�j���O���.h1�'��	�\� �T��SM�%k�p�QӁR/4����>7G���?���?Y�
	�y\���I;z6��W%D5e�&�'G �[�+�>�(O���3���:�{p\��Ř�ȏ�EPB�;�R�t@���ޟ�'?��'(�_�\��O�".�.���'I+;T�њ�)Te t	��OP��?	K>����?���,U|��%b�=}u�huiP�#�&Y�����D�O�D�O����y�:���[���t�zq�����-�$�i��IԟP$���	ԟ��A���Ba��æ�� E�0I&˒N�����O&���O<�[����!V?i�Ɉ+qRs!�r�ny�"��4-+��ߴ�?�M>	��?Ya�M8��'^��"A��!���R!3,�,[�4�?����dL�p/�X�O���'{��J�L��� �ޚ'x `�ɸ*t6O*��O(�ze/��]:T��>%���[��E�e̒Y�ч��Y�'�UjF�z�`X�O���O���(\|Ai�C�Ʀq��dD`�a۴����Ov��[��w�s�N�����NG�j���a���qԴi�,E�Ѓh�D�D�O�$���%��S�F�>��U�Qy��+~r2�
�4%������?i-O�����O�����/{���Kd��|�d�	঩�	��x��B��L<�'�?1�'�ɸ!"�*^иi���7a|	��4�?Y-O�|�ČF��'B��'-2�>8XXL�R/Q'a��Ȃ�K�`@6-�O:IV#QR�i>u��b�i�ո׍@R R�b�)�ڣ΢>1���?H>����d�Oja���΅A�P4��'
<���cAU��ʓ�?�����'s��'�T3��>Y��Q�A�v�ЅcP�\�.�ҁ�yR�'��	ɟ̣e�eb�N��{r�a'O�(n=>d�aNF����ßL�?y��?1D�K�ffYl�-I�TɆ�
�TBJi G�j�TO��D�<A�x	f�*�.�$ �ŀ6A��}|�;D!D+gp�ne���?���w�	��z≞I�}�w�ǜ3� ���ߤkS7��O���?�a��$���O��d�k솉wz�D��O&��}(#��m�''B�'��Ly��+����	�+� =�v�N�B=�c���Ca������͙П�Iӟ4�I�?��u''�/d���Y�X&h
���U��M����?����'=F�L�<�~2c<��}��P$u�z	)ר�٦�Xg��M;��?������x�O��;�V>cܥJ6mΏ0?r��a�lӊ4sR��O��ħ<�J~�'`�A��-F&�C��I;�h�h�v���O���ďF��S�T�>�����YA���i�&��US��Gw1O&Iz�B�c�S���	��5��-Ȱ8E�4{������M��"��e���x�O2�|rgKM��:ą�d����@� h���z�j-J����?).O��ęW�? �TK�d+ư5b.R��`���5��D�On�$?�����ɠ,*��q o�$s\�ax�a!w��ACjΡxHc���Iuy��'�d!�֟4(����%�JX*�@�W�,���i���'��O����O����Y�r5��`\K��1q�� �a�ʱAۃ����O��$�O�2Ul@����Bl���������aW:-��7��O��O���6�p�����LJTA^,L��
$�S/2�|7M�O���<�T*F
x`�O����5FdA	��� .]Q�!2a�������sB�d"�i�?�J�f�,+R�����u���W.s��ʓ O�ݦ�ʬ�R�$�x��'mu�6f�!���"R�N�}�T(j�4�򤞷0,���T[�m�s�rQ��N"3!�$��BC:�pPK�iwfUJ��'"�'[��OZ�)��N a��!�������x��+W��N4��+�y��i�O�13r!؍JiL�iCb&����KԦ���������~���OL˓�?��'s@=��*�,. ̕�S�Ed��H�4��ew���S���'���'&4P��*N�Bu�&�έu�@��n�B�Č:$�t��'9������'8Zc��I�B��H�`L�}���X�Of혀�����ʟ �	��p�'�>P���y/���`J��tH�!�Z�8&����d�Ojʓ�?I��?a#	�/{mj��ǂ��<XBP��rѼD���$�O���OJ�x��i =��9i�x�lA�J*]��T�ļie�I⟤�'d�'�B��7�y��0�ʹ�EC0F�2��>-�$6m�O����Oj���<���MW������*G��5n�"pn�<H�t��Ɠ��M�����O����O��>O<�$����/֙Z��a��=0���k5{�p���O"�y�ꌳ [?e�I������X f�Cb�0��uE��52B��O����O���&K�d�O�ʓ��tO�����J
�!���"$��M)O� �'�֦a��ʟ��I�?UڪO�n�P��V�П=B�u��n�.���'��n�����<���T�?xJN�i fI�^`8#�7�M�냉k�6�'���'�����>q.O��{d@�(fJ�%��16�yh�ȑ�=�AH`�'�$���fSa��U~�v#�Cª[Q2P���iB�'�B�j�2�����Ov�	�H�����77z� 3,�']�6-�O ʓ>���S���'PR�'���5v�J,��I�d���lӴ�d�:/�Ȥ�'���ܕ'Zc�l���s�fX�@Y'3`�A�O����5O��$�OD�D�O��d�<�퀍ao$d��(�;��D�פ���V���'}�R���������,����L�q�N�{` H:")j��7La����������H�INy"N�瓻%!88�s�I��E�Z8��7M�<!����d�O����OrA�e7OPp�r��z�A:�ۓl��]B@������������'�I���~z��C[҅+��^
��3Ċ(Ac,ɫйi$S��	ş��I! ���	a��[�B��Հ�/\H�;�f�����'��U�����R�����O��������T2���ƉE�=���Vb}��'-��'E��O^ʓ���N\��L���Ԑ.?�@s�W��M�,OYP�%Aئm�	�H���?��O�NN(�Z�P��@7D'v��6�R ����'��nG��y2�'�r�'�q�"�`d����UTf��C�i�65x@/`��d�O��D��'���h[z����.	X�Jd��V��*ڴU�Bm�����O��+ �Uе�@6��8i�j,oZş������hq�_3��d�<���~����t��qV�]4=4�I��o �M[��?a��'"&�S���'|��'��E#��� )�����H�H�@Hw�f�$ǌv�.5�'��	֟�'�Zcgj�
m@�	K�pa	#o�l��O��T>O���O���Or��<��a�>�x��CxL�sfgP�644%�q\���'�R�����4�I)���Qs�Й)�\ġ�/�>5�2��a�a���'���'\V��
C5���N��(V>���i_�[N0��J��M�(O ��<����?��z�^͓QF9&DՍvWDqF��}IVY�V�i�B�'��'��I�:�8������cf��S��YE�I��N
�2Ul���x�'S��'��-��y�>�*�7H���
�)�2G�P�G
���	П��'���~���?Q�������^�N�"�Y ^�.x_���I�����Z~#<�O�:X-`��ׄS p�Иp5���M�*O���Q�m��ן��	�?�q�O��=y�ܻu�T�3� ��,�+oq�6�'��H����D�<!���-M)n�(T��fB#TSν�C�M#s�U�<��f�'��'��(�>y-O:q�G�U7�\�č>���Z�ʜΦA�W`��$������uݐ�HV헃5.��z��.7�> "�i�2�'nb���D\Dꓵ���O��I4g�%�M�-W��*@Ǘ�0�(6-�O��[e�I�S��'���'��2��E������d/	`���`(b���d(U�ha�'��ȟ��'�Zc�|���B�${�:a����"�X�X�4�?����<-O:�d�O8�d�<��g[�-E�P6A%"�>���I�s�aeT�0�'�[�4��͟��/}��d�Q(��F�|�ƄO:�B�p�On���'B�'�Z�H�ķ��T�2G`'I[?6A��7���M.O8���<	��?��-���'����Q�_��ۧjJq��1޴�?����?q����Sg��OgZ� ���@�KTM
��Pn�:%����i}�[��������	&5В�I_�ď����	�t�^eD�	أ �?8�&7��O����<	���0�O��O��9�0!Ʃx@��c�)t���;!2���OT��Z�_$��/�d�?y�"�,����.a ��y�nn�&��3v�i���'�?��'T�	�*i���V�ظ,�Xe�#(ɬ7@�6�O��d@�F9�D(��0�*� �P OH>���ʊ'xݢ6���<Rm�꟬�I��T�S4���?�ᎶX.�p�/��Oo �2q�F5\$��ˎ>/|���O<y�FĀ�a#����]��uФJNݦU�	����ɕk�V)��}b�'���)����o�kZ�E���޿V���|"�ڟM�2P�H��Ο��i��
�$O&~$|iUa��Z,!�tӐ�����%�4����'pZc:��I���=��Tɠ��=?
䝈�O�����O���?���?�/OJ+ ���X�k�肻T�&�	��K� "��>�����?����"�!�숄冀p���-lT��$��<�(O���Oz�ģ<�iZ�;��	'�D�DH����#V�2{�������s�����	�s�z�	y�>Y��K�c��S7nO7u�A�O���O��Ĩ<i�.��N|�`叓p$�^�V����.W�Aƛ�'��'��'�`U�'����

pW�e���O.j�]n�̟@�	|y�� �������.���:� �޹e�p!��_�����IE^fm�	F�e�c��	O08�V
�B#�SD����'V�)|�9�Ob�O���k84�
��:b���IZ:��5n�柘��	��M��v�	[�'#�E�P'�.Zsl����bt"-n�=TP� �ݴ�?1��?��'x��O�E@�KH%�ty��!�2��G�	XQ�v��'�����3�F�S�ꅬ�
 Z�m[ +jX�� �i~�'�b��Q�BOT���O��I:y�(��aH�An�K��Įy6m<�$'T�.4$>������9-���0�ؽ+����u�BE쭓ߴ�?�'U�H��O��0���x9*���2*����J�58�l�^��;��C��ԕ'���'�BW�t v$ �8K�DiM.{�0�p o�h �K<����hOx�	�q&�,�c/\�!�ۣ��_�n7�O�˓�?����?!/O�T��K�|����q�hy7�R�x$�}��N}R�'�ў\�'��a	:yHp1rcH�|�顧��:p��?����?y��?�����I�O ���C�*�A���ԨA b�æ���r����'��asK<Qf͆P;�4;"EC�P|\�C�Jզ��I؟l�'adp��-'�I�O�Ʉ�N�̂w��	%z���	�vV�mU�O�6LD����Mk7�D(�,]�����2������֦������	ҟ��	ȟH�I�?i��5&	B2;92|h��b^�Ը����MC���D+���f�-Ȯa�Lє$��m���#o?��a��LM�7M�O����O��p}�_���R�J*p{��`G-�ܥ�퓦�M+�BU�<�I>Q���'��i�J^&F�|k�-�7�x�r#v�����O��$��E[���'��	ڟp��8j����D�"t���p�R2t���oן,�I�t�d�~��?Q��?�B�ʉ?���&zE��eNߛ��'�Hp���>)O���<	������ ��'���a�x5[ w}��;�y��'�r�'���'�剉5*�0� �x��!�BM.ob�����=���<!����$�Op���O&U��	8�$r�L>����M>>��؟��ݟ��Dyr`�l����A?��S��[�}]�!zG[=R�7�<�������O����OL��]�ȣF�F,L�xx�'�c�y�Iy�
���O����O:�����$^?Y�i�%�	���(` B��N��iv�����<����?���0Ӵt���ihj ,Q2[eN��	��f�ܴ�?)���$�7*�8�O���'!�����*͂ �/�JJi,�F$���>����?��e���̓��9O��ӬTKV� 2/�	�~(��dO&Q>�7M�<��Xx�6�'A"�'���d�>�;:5� �E��^�D�1���g�P4oן��	�f��Iȟx��ʟ$�}Z��G�ָ"�fv��"ꦕi�-]��Mk��?I���j�Z���'�Ђ�n�Z��_�{pڠ�bw�D�18O��D�<����'ഀd��f����vJ��J:x�P�~���D�OL�D��2˾�'���ҟ0�xZ�p7i݈���
��#�9o韨�I�<qfDi��'�?���?a���gK꽳�KW(T����wmL>���'����>�+O�d�<����� C���A�45�s	���)����$�I����֟L�O`�ć�ܪ֕�=0(Р��!D���I����I���_�	��R�^)�A�P>Z��=�ElQq���m�˶��?����?),O���	��|*��D�B�2�G1n��%	�jJq}"�']��'R�OJ��f[?��Rg��{Ж�z��ւ-[z�#�k�>����?y���?��<F�<A(�p�$Δ%��qb� >�(d���#�^qmğ�%���IDy��L��ēZ�q���W�+O�� c��&`�>\B&���'��>�I�Ag
9�f�:�%�d�O�b�C�	/r�<C2h	j���Q�KL�E�6�Bp�	2 ���vm���;7��*
k�P���z��!q����m�f\��,� �HӦ投�,�r�ɟg*5�&�)WF�h�����rL�� _f�x�%���,"L(�2?����	�#C6�01���i^�`@����C�h�+\j����͗:KX$p�iR`�b
ť�O��d�O�$Ϻ#DO7/�xH9���e�ҭ{��5u��P�!ʎ4����'U �+��4�0}��@�]Ҭy3@@�t9R��U�c��4ʃ�m�9��#((�};���.��(�v�	�I	`q1Ge
(���7E�$Og�)��[~b���?ͧ�hO�(EE�F|�8�`R�Q#�"O"�HGo�'0Ŏm��"T%z� y���� ���?�'�ƄD˅I�i��'X����A���t�����'kr�'�b{�9��ޟ�ϧNu:]@O̞�|L�
A��0qH�ͅ�#��PHj�,v�a{r��Z�u����Ref]/K�Fe���78�zyS�ڔCa{r�P�4�b�퉚�)P �N�t�"yq��?I���!��t��h��P&�ΰÎM3^�B䉕Q��EB�#�	M��R�o�
p��b� ��O�ʓ@�*IPRU���	�'+��Y'η뎌z�-Ǳ
N���ܟ��e��\�I�|�Յ��hx�pK􏎭4k��_�oՈ�4�X�6	���#ܛ��x���5W��cm�@���"M����(Q���r��1�R���D�[���'��	�{o�@����/l�h�;$.�<v�b���	�B�
h��O�x�,���Q�Z�&B��2�M�j�H�A� g�p}"�%M�<I,OLD���Lw}��'�#`�b��I�~�p���o�u�7f���J��	ߟ@ �N���I���|�*�2�����L��u*6�w��4`�>i���-�^	XæE�Q?��e��P����)���"��:}BJ��?I��h�`��#M�-8�"�
��i0��� YW!�H�KM\]���i��1�V
=g?ax=�V�L7�ƿ�\��� ��N��a]����ԟ��EG��v����	��������y��	al.	��c�l�}cY��L� �4Y������ UN�g�	,R��� 2m��9�C�0b��|�"�9���J��kQ�Z��.�3�Ā�1nĜ����h���0Dh�xPh�*?Q��؟�SX�'Q@Đ+V+��eK�*�'R��	
�'�|��mÒK,�	
eΕ(0��O��Dzʟ4ʓ!�^�´/�]�l"DK�x/����'&T а���?���?ᦷ�t���O���-���"@ɜ5��C��EK6����a��%fԜpP�]� 5�(�W�'�H$HgKon@� ́(��&�qQh|��0�΀�gLN8�X����n�\�4B^	ލ)�@��[Jb�d����`�4��'6Xb?�J#�O10�*Ł��,��M�n'D��qI�$~��P�Y���?��)��Ľ<�w ^�q̛��'�򩚛^��L�EƏ�vB�Y���Q	D�2�'�Ldi��'RR�'�P���JIV7LYzv��r��H�.��-Y��L+z�n�����p<I5Ù�˨af�f>��3� E?&���Q�G�.P�� Zs��7q>���	:=����OV�o���Y4-]�_�(�h��
/f�<����_y��'��O>�Z'�C�dW=��,I�(�y���Rk�����Xo"����U���[#��'L�:(6 �Id�'�ў��R+�}�z�y7Ί0ef1@�@"D��1�NT,#��!9B�X�VnR{�'Ӱiz�.N�A�]C��;`36�z�'Q���FfO�54A��%=+�2p��'iXM�A�5ʎ��"N^���'B)�!M�C5��Í!<�A��'c�}JD�(�eS��֗	�����'\T��)�LR��a�^N���B�'��|�1J��C�½�Ѩ��G!2M��'ÌQ�D��'iB0���H�+h��'�H�Bq���y`�	ăC�v��2�'M��V�X+�ZH�Cb۫ aZh
�'�F<c ̑�)�u��J��,قp(
�'e��㡣H4<�])bfC/A2��	�'@�+q1vH�	F�+t$�	�'��	;6΀�i�2	[�B�18�s	�'P�H���<p���i+ŜWENT		�'�L�P��XH��2d��L�h5��'��d���)��c�
m�9��'����t�E�kzpػ�g�l��!��'��)+�e[BT��C�)�Z�pq�'�P���=D �2�)U�@,q��� �0v�J���C@����"O�ũ�� ��r�_�eoL!x�"O��7.M !��m�b��+ISޑIt"O�t��ڃ^L�FN==Cm�&"O�����ߔ+hHC1n
�|<�1�A"O�M�蓌)�zm�f�;5�PP�"Oz�x�慦j���Wo܎C���ˁ"Obѫ���*7��y�-�;<�p���"Ob���D�z(�h���1�@�k�"O������w��P�Ѹ^
0yA"O�e{҂�7�V�&�Kg`��s�"O@|ZR�D)�r��gԬ^�`�"O�D�@�� 	�ݨ�!"r��}��"O�H4�ڽm��0 Gʚ�KQ"Ovm���+��9+%��(�z�AR"O��'�'Tcl-9D��6��lX�"O|�f�G�P}�pd�ҖAZ*�q4"O�a�E�z,
9+�*
s2�P5"O�8�#��8J0� P�k�����"O�HCr�ʕK�� �D6@*c"O �	U@�&_$�00J',�!��"O��/\����Ԡҝe�����"O��ă\3B�~��gBʘč�$"O�L���ʯ`]Ҥ8��'��q8B"O�1!���2ƌīR�5/�Xp3"O =�f%�ل����!o�pe"O��`ü���B-Ĩc4���y���'m��2b�
>�����:�y��FNJqq�k�7�xlIv�Q��y2��2C�&���V �k�CY�y�I�W�\�ƵE���T�ћ�y�jM�}U�,z�"Q#o�h���*���y�`��y����wY�_�@2����y"A�"��c�ީ'$��dǎ%�y�!J�a��tmT�%ܴA�!��yr"�W-(����!k��2L��yAR ��؊�	(*�~�g���y�I0&���jD��+O��p�+��ybd	�h<�����^V�};ƀ��y��U�+8 ����E4�\Ce�М�y2���%���i�㈁I�AB��yB��#<�|3�&��������y����5y�M���H,
��0`�S��y�1*J���� 0�ț�H�yⅉ��⍃��'���# <�yI߻�ȱa&��2��X�dM��ylߩE�V�k��D�1�L8�Y!�yRm��*�,�q%<,`y�ȃ*�y�BW%����&	�7h�Qq$��y�&�,-c�b#҈d0R������y�DJ7st�#��ПD�<��t�X&kF�Ts���;�g?IC�Ycb�0�Ye[$4�$�t�<��CXm��;7\�&���v ^*9a}�d
�+���mͬtގm�3P��=	g�ٴ9+�X��$2��
�N(+����U��'��}
��["i�j�*��:e*#�ҧM'fP��E��/�Ո����!�"l!���z�<��CDANY���D8	�O[?I��W��h���zeL���b4H�*5>��"OD:i;�� �6(��*��>�%�-��=�%Q�
H��c����Y01��G��,�ca�Ԧ}�&���=ٱ� �2�K�o%D���F٧c�ʹ�t*Ax�� ���;Ka�]z��=?A�&½�~ʟƹ����ӓ�X�aH:�h�N?"����z�<� �4��7���p͛.q�F-	��N!(��Ʌ��$ݘ_�7�����S�D�Z-/ 24:P)W�0�a��J��0=I����v������<7�C�C��17$x�mCq�pл��
D�13cQ��'��'����F�I&ƀ�e�B��ڍy��F�КŁ[����yZw?�T������S�@���Y�'��r���	UA����%2���X��H�<�@Ѭ^;A�yb�HI���8~���|
��@�\�ݰB��K)���0/A�$���t�;\00���8���Q"�	��(�05Y(4�S��.k9 ua����<Q��Z\U�鱐(}ʟ}�PBYB��!A����6Aj�'쀀�eT�]�0�H�'�e���G��Tl��a���<�#CH���ɦF�֟��u������lH�H�IZ�n���zg�U�E����<9�T�A��̓dK�O���6��ڨ-���%��A��i@�cJ�B���@XR��$\O�`޻l��`I�L�rCܘ[��3��V���q7��?��ң�DK@*�ȕ�eNjd�	�Mb��YB��?A!�L�#	!�$�s&B8�v�a��%��!��*�2q�"��o�< S"�G�؂m�D"�"����4$�Dc>�#0$��X8��zkϪIAlJ� 6LOz�5gԦ$	&"�;O\�#��?�.��D�)Y$z|�d�]
p ���
��M3!�\�/Pl�>�O���>S�Ht9�� s)Dٷ��"w!T8�7�K2E�Q>�^�C�xS^nH��Ab@�5`�8-�'P`��(F,�p=)�DZ���a!���@�(ɋ��MX����NJ#A�P���?z�؁K�L�U��[q��d��&��y"L�9����u`���0���!��w��`q��[R��*1���(��d�����7ԙ�!�Y4cK�`��"OH顲`'l<9�@�4���P��.J�Fp!����y�� O���(Į� �!T�q"�[A!\u'���R�"��Ս_K����j>&&��+bӺ�g�I�^ތ�דG�И�����x�"4K�:ʞ)���L�j)y��	֦I����c|�����`���8��,D�`B���8\x�Ra��t�#�(D���PcJ25�ҭ�f(����"D� �B�RBq� *L��9:1$,D�H����r��J�0��Q��*D�(��̙3v�>!�Q�GN�����y�Nڇ�T(u��I���Z�@���yR���4cԙ1���<V� �`����yr��-6u2�+�M��ap���2�yb&X->xU��̞3[�0D��@7�y�ϡR ���G�%B������y�څ�X�C�!�F���B��y��֣*�\Q�#ܷ�L �D���y���8J���f؈Q>%��P�y�Hۍk�H�&�R$��Z�Ȭ�yb�U Y(use�E.[�8	ă�,�y�lعg+�Dc�G���C&e�-�y� T�;h�Z`��3L��l�@+L �y"�¦�b	����J�Dle��~�KI�^v��$�5��y�D�1J'�E��i@(4N�|��ߤ�����_��A��Xб���E�C��$�՚g�ґ^��!Ѡ���r�<)�*� �Q?��R�̞ �����"o�>����)D��"AO2"�a �Tr]Q��H),�a����O�ZvaG9Z�P�A�H)Z���"OV�yG�A�?BlK�D�'&1�$�R��Q�#9�O@ʤ���[��-h��m.�$�'"O�<zP�+�8�Ec� {n0x3"O��J0ː ;���ʉl����"Ox�A�S�(l���gʰ�F�C�Q���V#%�S�O�0}B��H�`�.	���^&]�e�'��P�![�M7��
�"�2IU��O>IV"�0�0=���`��Ԑ�M�,fdpf�	_�����L��I�E�sn�z���s�m��G��e�uNGQnez)M	4��F	�;e>Őc-ӧ8eR�[�$��7u�����1D����٠��)ԥ���T���B�<��Q����(�� 2P���هV�yp����:�pIV"Oba��$'���0��K�2�p%ȡ�|�J�6�az2�t��<��8��h]8�p>�cJ�q頬���w� `��7\�T2aO�C�bB�	/F�Q@A�Sb� 1�,̳$�<��B-B�#~2"��7����ѡē�z�B�c�^�<95�C�14fU�F�H*!�E�ѵS;(�[�cWG�S��?�B$؀*K� 3 ��RQ|���
�K�<�%��<�zx���n[���̌q?U�ZK�`��$،n����
B�1$FP���~Y�|�A���E�w�@�jc�3R]������g�z`��!��!����s/�%pfD�v�Dy�`%��F�D�۞��U˒�$�U�3��8�y��1#�x�ʰ(�}E��l��h��9s��F������R&Rb ��QG�yL������y�����\����u��y��L��~bʌV8���1&�xcŁ?������Y�l���$�>�(͓\�n�҆��5$ʹAӑ
V�-�f��HJѬ])wp@�4�o���ȓxP.��g+`7�)[W��2�|��oU�q��d�.>t8�5ߡT\�x�ȓ��[�eœ����s�ܨYY� ���Dp2��
mk��$æ!�ȓpEVݺ��#A�����lw|�ȓV��e�� ����S��l=�3"O�����4$#���֜P��1p�"O2-��,E�7g�!����/l�H�) "O�`yƉ֦}��d�5�V)Ku"O�%�Uҩ7j�!�T
�Si9t"O��$!�'<�aˠE�*PT�V"O�!J�!/�Xp��]T�@H�"O�5Ru���/G������,P$��"O��'HF�F��pí�?(� <0"O�}��������3f��4�*\`Q"O��z���r�l{���),䶆"O��
0��$.�V����ε4z���"O4�I����m�t�Y�-�+I%ش"O@�:�B�2e8����Ŀ;���	"OJ�wN�#�d�j�+���}�"O2�Ė�p9���Q�b����"O�-� ] %�.�x�	V7U��Yx�"O�p�!��x�e�1�Em���u"O�Q !��<L�"
�*�.��$"O�\j��
��h:�������"OV� T��^���A��2�h"O����J+ӈhH�V/l���"O���B�u>�y�ȥeԆh�&"OLĹ��a~l�bJ¹<�<5�"O(dj�A1:�4���^�^��"O���"�V)+Gp��l�;_ʶɘ�"O�)����p���2�X�QƝS"Ov�H�A�^�a�ơ Ej�e�"O��1��ާUf�Ҥ�S�W A�$"O
�!�.HN��K҅Y悕�"O0](��؄%�@j�+ؙ�ҐHv"O����(M482H����H�n�  "O>d+cA�&9D�vO�>��E)F"Odx�d$�
a�F��.C"��"O�8�Q�r�n�#7K F�PKf"OB@�BPep���k3Q֐���"O�$����|�H�y�ʐ�St��s"O�s1a;��Yc Ģ6j���f"Ob�*cŞ�C��I�d\\��x�"Ot<�A Tk��t�F��UX��,�y
� h�YW搷[|�%k���1�"O���v�G�y �m��j������"O�� �%Q_��9sO�$p{paie"O��@�˟�8�&PY�6
��ۡ"O��(!&٥|X�ɢPjŜ/��$	�"OH��s��ѹ�^~�`��"Or|
���>2謹0h�{	��0T"O��*E$(j`���W�*(�"O�r4n�7���Y�
�%��s#"O2%�b�͌H�F|�VJʦ{
ڰ�"Of����;Z���f\�^� 8�"O6� �D�"��@�\:�N$0�"O,@#0�J-vg�:3KE�p����$,\O�9�Рӳ(�J�*R
JWZ�[0"O�a9�n�	=�F����]�&;
x3"O��ktn/>���۱��--5D��"O����Z� Q��Z�l�0# �h��"ORة��%2Ơ�aj̜��a"O��rD��,��Y�W�n�0f"O9xt#Ɉ3ha�.Ҭ�w"Ob��QGI�6�^\�@.�fEP'"O�0S� �M�p��`��Q�x�"O�djֆ@�(�l  Qn�G����"OR�� �_?Ӗh���D*Y:|�"O�jW�C�E����,P�X@B�"O(yT��Y&�𰠋�n�n1QB"O�y��O/]t6���l���� 5"Ox�5�� g�Dʐ�ǡ{��i*�"ODd�vl.R�����k҄�6aX�"O�)�f��D�X����mb���"O0�K�f\唰���EpO���u"O4<�@$Z%���ZЈ�`�
5��"O�x3�)��H�0Y�FH�I���"O&Tz�B
_����Bvv(��|��'lfA��<^��.�0*�Q0�'y���a�ۇ$;�	��J�*n���'=Z��F�ܰ/q�C#D?�0�
�'D�dső&�|5#M֖Q�=�	�'=\ĪfL�zz�a�cQ�b�N)�
�'���8��8�Ux6��D�$�8�'_����%�$ c�EEL���'����4V�8�^��Q��!4�|��'�l+�q�l�� hk�X���M���R�Yc�j  �F�Z���"O�ЕB-x� �r�O=C�:���"O��ʄ�S�,�����#��{#"O<��6�K*I)�s�B�Q�J���"O*�s��c�$q���G�C9��h�"O���)Ǿ�P< ��+��<�F"O�<��$�z���I��9/���1�"O��ip��_,���S�\��"O,)E�ݢ��Q�ńПR��B"O@�V&
�nyK���kh����"O|L�c.���x��ā�u+\��"O�8�Ƈ�;^��@�\}���w"O�)ǥV  ���F,��8�S"ObQ���mXצH\{D��q"O��K��$x<J����Wy�0`�"O�E��e�?|�̢7oԣ����"Ori���\�|�*k���t).�h�"O Qsao��\R�Q0"�Y�$��cV"Otɘ%`�5Vd0��b+T
[�I �P�\G{��)X,n@J�[6��Z�D!3U�,�!�$D,<K�Jw	��Ll��	$���%�!�� �����ô^�dL��[�V�zC"O����J3%క
TnU#��u��"O�Ӣ�L"�t���b���	�"Or0!2�� Bb �5-��fo�YJA"O��9�
���(��˒WV¤J�"Ol�`��ˁ�:  %��.8B\Z�"O���Wώ4+,�1��zĴ)9�"O6�N�?x��(C��P;L��l��"OP̪��H]��K��ͨ�E"O���!����Q�&ZbD��A"O��)�鈳0��D�BA�W�H�!"O�*$N2c���@�ɛf�<��r"O\�Fn�V��LS���!n岗"O`i;Uc��jx��ǧ�� v��"Olu����S������Ȣi�T��"O��Z�Ɛw[�ĳB�9d�u�U"Oy;fL�nd�8Ea� .����"O���t�߈Z갡��	~E�%�0�'m�dE�P
���Ѫv��`�DCR�O�!�D��M."�K���Dꊬ����,C!�d�7j:�jd��=�3.**!���Nb"ܒ�j�'d�!
����!#!���#M��sa��~J�P@X�7!򤋁py���"�/A-&y8į�4!�%@�b��'T���y-!�$������q4r��3B�!�D*9�rq�
��} �����<u�!�$�����h�6���5'��!��A����쎴D�詆���!�dD]�XԢ�NR���F�V5E!�sy؅�S���\���5��s�!�'Y+��"�$݉D�T�dL�n�!�$P�x�A$G �
G�)�G�2- !�DUq$��$��&��i��� s�!����]B ��-����B;U!�DڡA�Ƹ3Ge�L���B��%7!�$��G�,]��C�%j���LDG.!�D%2T�X�j��\�I��Ȥb�!��4�`��
G�#V����ݹ�!�P��
���F
A.��p�M�y!�_5�j�˲�
�%&#�o��$ !��Ck�Ꝼ�NY#qR�T�!��صL�T��3#G�ETj8�0�x�!�7�j �""�"E��p3*Y�t�!�$��,�P%4}��mjd	E�a�!�DE7R��yX�D��p��p��'�!�K0��a��δg�l�s��PrU!���W�(��B D�X�&j��Z$K!�D�4h� �o�<&p�UQ&R�F2!��3�  d#�%�����Gu,!�d�X�ڝ��a .�d��$+!��Ȼ9�T�`��5c6�}#�=E%!��ψe=`ڵf�)C4]Y`J& !�	�"C�`��,j����t�7}!�!wL(I�N�U|"�����kc!�^�G����B� ev���	F!�DZD�$���pp4��&#�!�䀓K"���l%=�4�jI�V%!��[�6O�`i��� H�b��w�!���&��`yrm��J!�$�7�p����3���lMqJ!������ �[�Z��	ِK�j5!��Q61��(W�@�>��j�F�!��t��5+��Y|�l����~t!�� �)qhM$	7񀅫Ҥ���r�"O���r�S4j%���I��c�`�r"O�}�fc?6�z|YF��Xl���"O����ā7<?T��Ei�y�J��yR�W.7YP��Wn�{��� r"ˉ�y�G��&�~�{��� �:�[!	Bs�<�3�B�
��ܫaHM8ـL��[U�'Ta�t��(K����=5�� 0p���y�합m"�uQ���*��1�l���y��;sth�BS75���M� �yrN)����D���L��4�y���2����-���3v�Q��y�候%�����ɼVn�A+��0��-�O~ + e�% ��b��]!�"OИ�G�:�`q�a�Ɋ7��%"O�ZG�ҭO�0m�0�ߒb넉���IwX��I���;d2	0��Y�-C���3�>D��J��<�r`�2iY:;���Ã!1D�P�S���-�0��p��vAx���a.D�����/�����3ih!��C+D���fA�$w�.��$cյQҀ@h�h$D����D�/!�g./2>R�)/$D�|����_��M)Ư��`u:��$D�X�H�5p��r��M-0
x1���!D�4�3d�Tň�����<���M>D������ 
���hi(:� �<D����B�"�*Dc��ǾR4U��m5D�4z��'t2�J7!nz�s�,2D��sAeʰ;��P��V+s�D��.D��K�U5[@ (,���z�-D�8��A��6��J�5�(PW.D��#uȳI^�A�.�{��\���(D��rӠ^�w�J�y��جWV��3�9D�T���.���+����XpE��B*D� �ʗ�B��[�)]:|5
%[Wg)D�D�_=T�(�s���٠%3D�<�G�ل%צʕiC1;$��	�+D��n�!vM\� ��kɆ���7D�H��MBxU����>?�2�`7D��Q���+8�)R��l�n��"D�����2<)�WnO`��d !D�p)Р΋��hF�|YX�?D�@��D^,�����B�1��+D� ��휪)�<q+w$Υ_�,1A�i?D�XY���� K4c��8�8�7D����
G���`��.��s����3D�,�E�8sO�|�6!S��l鳇&D��0���)<���`��f�t��R�8D�(��Ä\d�
X*B��0���1D�@��f��<�L�J O�zXk�/D�<�š��}��`�S�͛B�tls��.D�pC��v)��&�>n�Zhc#'7D�����//���-�8��C��3D��� ���C8�l����[�����&T��p�H�3�:{&֔X��)��"O�,��BF23�ZX�B ّ\���	�"O�����,/���a��(�� Q"O\��i�
��y���.�F�:"O�@P�E�[il)��'3Fkf���"OR�:u�]�)�y4hG�TK�d��"O�i�5%�!p� :s���:���s"O41�` �5�:���O`Y��)�"Oر����;l�����^�)ߊ`�"O�Q�g��iҌ53�DռGh���"O�  �#�N2)���cO�co�d{"O�7�K.�;��
.Q|T��"O�����;l<H04`��#{0�s�"O��i���4�x�1�� ^r`m "O�l����4�>�D�F8\e���"O��[Q��J/�]x����>*�$9"O��Ò�Ƈ�Xic��yq�|�s"O�D���@�Ф�p�=M�\le"O�AC���)6N�����$Ja"O@L�a��0��  �� �LiC�"O�T�'�=j��� �a�+T٤�p7"O��cUG�3a_��1N� Mm�Бc"O4�2�΍�-�\�"�_�xXx�21"O:� �J�~��w���x;D�� "Oj��&�p2��aR��1)^aS"O.Q��/Q���A�D�-N�Ҁ��"Ol)�� !�`]+�HAה�B"O,��d��H��)8�C5.��"O�|(Q T�z�Zm�^�[Ղh:�"O.��#���"y+�Μ3u����S"O`��RlV�������X$�"O�*�K.m�y!������"O�M����54((��.�L��yJG"O �y��ݽ����֮�g�&�P"O�x1#�?j���u5�� [�"O�%�v�:/�9z�"��1R�"O�<:�	5?U8�P1�:�!��"O�Q#�%=
,�Q��(|����"O����Q�@<"E�F�5�����"O.1�U瑁��p��eid܁�"O0!z�C�;�����خ	VޑA"O�Y��Z'���#`��'��T	"Or�a��[�FjZ9�r���\�{�"O��[u,X7?dDtcq��H����Q"OL�Z4��	� ��p�@!�����"OVē �Yh,��
��8kC"O�|H����L>���$J�n���"O�t���)9}(��Rr�� �"O���kZJf�@� ;M��D0"O΀�G��n3�pk�K�I�hX�"O�9R�M+{v���XEC$aC�"O~x��ޯ1�&��4�	;+V�I`�"O�B��X��铱��!M�n�:a"Oj�`�CH5w��p�+�g�r@)C"O<�"i�3�-!#�)ʶ���q"Ox%��H�c�$Q�C'�!C�4b1"O�9x�d��7-v�a��<�,=�"OR�3�a.������#tD���"O���Dƀ{�� P ��;n�A��"O����
��KM����kʁ�y2J�?LJTp�O��t�TX�e��y�jI�P�p���	l]���!��(�yB��9PpjXE�Ҿ\;�+��y��ޱ!�E� ���~�*��ɐ��y⡙� Ҏ��Ì�e�z�"����y�%�jx8a�ʟL�`D:F�+�yr� #.y�bK�>�� ���y�G>i�l�D��v^-�w'A��y,[�X�6 �#��*f 	����y�n�e��������,�����	�y��<�rIR�#�80� �&��/�yB�׻pb,���"�D�(	+�y"O�!o��Q��m�(�~D҄
]&�y�)_A��5���ݯ
c�9%�U4�y
� �)����08��+��ւ/�|@�"O:x��-�.(�}�#�L-)t�"Ox��o߶�|H9mũ)�P���"O�P�#	�B�ܰj�+٫nʮ���"Ox��l�NG��qM]!%�2��"Ou��C&��R��Ƴwgz�Ӓ"O,��*�B�\ ����&TcЁ��"O:�@��9*x�4q*�*j�T�� "O��`qDF�{z������5��h��"O�E���]�^T {Vnݰ�F�@"O�0��Z�E)���2M��W��|�"O��b	-�,i8�Ič/��"O,2w�H!"ǖ ��)*��"O���!��"�F��	�h��� �"O���n�d�2�C��5!�*��"O�\���B����["�X� %"O�jW
A�q����"_a����d"O�,K��y�� �ЫD���s"OH�g%�%#z�œ��U���}R"Oz�HN"qI6 ��f�-u� �ȱ"ON��1[�SNa���8ozR4��"O��Adj�� f舁�؜NL�a20"O0�2�ѓum�d�H��:`����"O �@e-��2���b���n~�:"OT�zF�1_�R�TK>5a�ɢ�"O��Z� ]R���j2h2OV��r"OH(����/՚�;�l�CH&	р"O�)�"�ӨA��-r%S'!>�	�"OԜ!�N_Z�4W�I,5���"O���i�$6�^qҕ�H��.�"O��KR#ׯ&$�O2k3�"O(��mI*Z�C2n�6S�t�@"Ot�zR�I�	���v.���3�"O칋�f׈f)S!-�,r��Ӕ"O��ф��)f�����TXi.���"O>l��6}�����d��@�ʇ"O����D�)Q8uy�aC�h�6��"O�L!�NF�T8.܀d���`�'�.�ˡ B3��%��!�!{�@���'�v�(��8p.�*�dؾ����'|^�aRI��ZLT�&�Q04�`�1�'�
XA�/���P�G�"0����'ǲXۅ�Z"=���0��QJZ�h�'��͒���p��9b�U=�Z���'_X��`�@v�9T���U��'�Ę#CCW�����"�M��'v�Aq��]�f}�T/��|1����'��i�b��x-���Dd�_���'g>�:l���P��̜L����
�'��D�$��- �Lu����(F?lH�'ъ�0%E�*]����.F7��Ur�'�PR�D��>`�!��X�$q�'�Fu*nѱ�����2O�R��'���ӗn�e����]$J*�(�'zP��Û�R,JQkG��9W� 	9	�'.�}�W�54��IR"BH�1�'&B�KT?�A3�h;>��q	�'x����mƈ��H����3�p��'�:Q��MΈ9@�0u�� '�I�,Of���L�A�JD	�l�X�Yp��
�!��D��fͰ��ظwD�Qg��tq!���f��4(Q�	1T�
�@'!��H�s�j������$���;E�!�U�Y�&�D-f༭#�����!�O� �)�s�[�-���x���cD"OxuJ��]�#��4��Gӈ$��i�Z�P��N��X�lؖ%�@ɢ&�5]-𴀅c�<q��0>A�FM�NT��ӻ�H���^�<qB��3�����h
�3Z�僗$�O�<���*	0�d�W�E�	��$�H�<���Z|�M��"Ǆ{��CL�jyb�'�0�P�J͚q���9h�a�����'�*�b GU�#�D%���6a�4`K>i���(�I�P���C(�&�,%�~��ʓ�0?9����A^�;�RE��V�<�0O�/_^���7n¤])B��M�<-,�X��h^ �����Q�Մ�5�h����=!rmٌ`rx�'ja~2� ;(�x����&��zT�P���<�����'�tIK[qSR�B띃?@�Њ�'��H��cP�{餑"���	3�X���'���{��I�]ٺ<r�M
�
�'�������%P�yHIʞ���'p����Ξ9-:� Q�?{�(���'�h�$"����E�m�h��'~�	@mג#z�x�v�Jl�<DA	��'�kՃΊ|�\��O�mʩ	�'�q	��J��\K׋�5bHQ�'80�1ӥJ�^�h�[���X���P
�'E:=B�����s����B)t���r����E_T���dΞd!Z��ȓs,�8�w�G+�p���F�����7s�� ���:2+�!хͭb���ȓg���1��7! Mկ)n����ȓ�vtJfh�}8�d�d��(#�=��b�N�qu�֡;��Y@��
ȴ��ȓd�����/Ղ�~)�"��Zh��ȓ��;&��c�x3�@QC ���Dg8��2�KW��[Rn, ����ȓ�,i����,!2EN��%��KԖ!w�ǲ|%���'m
t��ȓO��y`a��RF�4Q��:���ȓ?!LtCU �j�eBI�fz����N�H�Å���g6!�� ?M����ft��Ca�$��E;<h����
l�q��������R�2Rh��4�t��A�.H'L�Sd��>����ᄠY���H���CD���>��D{r��o\�0ƥeu��Q L�f�X4�ȓP)�aqE�[��e��/B��h��{����	�EO�a�*[ p��J�n�B1��+2�l�u��%
	�����r��9" ��P�M�Y"���>���P.�=}Xf��sl�-��@��e��[v�W/<g.�p���j�$��{,��X�	��qojt� />�ԓ��x��W���g�2��c�,�>�y�G��2�1��׃|4e�M��y@�=ezn�A�,��x�-F��y҄ǯqk�l#wa��&`���Ć�yb�۶ T��p#ٙ�VE`��O���6�S�O1�a��މ8Ӽ����`f�D��'̺X�6LL�z�
�#�l��ZѠ5+�'0�� ��{>���C0Z�4i8�'M�����\����ri��Q;�H�
�'��`�,.A��e�R ��Y�H���'�,���#� �.��
Kh��'@��+0g�Mϒ��0d��o�<�x��� ������5�>�ڠ��C�P�y2"O�mi2�������To�N��P"OP �� �>
��A(vډb=�(�"O��A��6�Utl�p�
]� S�<�L�B����ːp FKAM�<	�L��4�C���i��(��KM�<Y��"p�L�'͘�$l���CS~�'�a��!����H�f�"���A�Ș�y��y��A3� �({�h��Wmƍ�yB����@�I�m��)�'���y"eۄT=��{"�B;drl�iW��Py*S�՞C�
/)6��2�m�<A4�#$�H��M�)n�F�:R%j�<��,L�!�Vt�#)�;�����d��hO�'n
5�f�R���a���0R��� |��y2n��X�<�1��$����z���Z=D^��4"�S�m9WD#D��ivŗ4�&�{pÇ�.�T��!D���q��#,�܈R���1��<:�	%D����7|�i��<=���C6D���$	�c���j�E�:=e�1b��2D������rH:���#��m�h$�O���-UV���HZ\G�$	v�O������s��$��!�2�1s��`C!�D%`%:��",�j�>�S�.Z1!�@�QF���.�]�|�8��T'!�=��c��6�\��D��]�!��+M"�점kܥD�n��� TY !�ֲ'�dh�MZ���G��B��ӭs��M
�9(a�&ܞ~�Hʓ�0?�2L��M�.��bAG{FL]{���D�<���""^q�1�^�j�[�fk�<�� ���4\rB㟋tRX��A�m�<���������Ѓ3Ԭ�5��U�<�ѭ�%MF,�A+�8+f{�<92͆�U��Ȓ;�B�R��M�<I�+�&$8�q��䐌q��0	G�<6�[�Dު��0����q��ȓ@�<YW
J�{�,!��ΠW� ����<q$l�U�uAt쐙d��W
�}�<Iҍ��on���3u�aY�GD�<	�Ɲ==8��0�L�8$��F�GX��4�Iq~�l,��b�%�����?�yB&��2P��3�S�h?���P�yB���3T�mxGWv��31��yJJ�`�T�X�`?i��R��	�yBh(O�IT	ޠQCvQ��"�=�y"!ߣ!@�$Lƕ:��<����y�B_�IbJ�9��A���=�yr L�L>D���
Ֆ$L�� �=�y�U�R{�]CjW,�j Z�c���y���+)�0��2��@��V- �y�A�/���+e޷Z^�e��Ɲ$�y�#���%a"�Xj��ɻp��)�y2	�uh����fD_˦i 0h���x"(;���]$J���H�n_�q�!�d�}�dlSeό�l�HirMиT�!� ;7��r�Y02����tm��_!��U?ϔ�#�H�V�@��%��wZ!�� 0p�r��&��)e�^���I�?!�D��$d��A�)�6��D��dO!��A;B�'���ӊ�6=!��̻Z��T�7�ُclH8B�K�NJ!�$�Y ٵ-o��4��T9!�� DIB���R�z)
��Ǐ}��Z"O�m��� �bXa�KkH;�"O�h%��M�j|p�N�-T��C"O�����0#"�@�c�]�����"O�X�$.,$y�Ƣ:x�t��B"Op6��V�\��O�h�R [U"O�hC�?F״D�6��6�8 S"Ov���E�F��铥(y��U�"O<m!���j�-rS��	<�(Y*"O*�!�D�Gb\c1�%k�b%!"O*���C%B&�Trq���q���"O���E��=+�!t��25��R"O�xٕ	S�cX�a� oV�q=�"O$S�$I	Xqr)0ahM�y��c�"OrrM�VA�4�v��2����b"Op�h�%����8�̡�N��y+̪�&lA�/ )L�%k���yR,E�Mn�Ap5�,����n�*�yro�� ���B�O2[�䣴�
��y���H` %��l`� :�$B/�y�Y�>caj��]гg΅��d7�O�y�D��{Hj� %#�wc��xV"O~�Ѱ�
?�m�⋓)�֜��"O����AŌ��4��=�p�ID"O\ ;�Ԕ2mX��¨��=~�ܛ"O��ϑ�&���R��By�ږ"O\����;$����kG�fR2)b�O�����@x���:(�ҁ��ù<����&�I�{�^�ad��e���"�C�'4$B�	�/NBh�!�7N;T(�%'i2C�	�8�zY��
�H�+3F��2�\C�)��L��I�N�>p�(^Ex�C�I+#��9�G'��?L\q�M��bC��@�����͉�(��^�2sFC�I�
��P�Z(Y]�d��E\�6�����bx�h�<���fYH���+҂�f�
3��z�<�M��-K�qJ ��"�
�Ԩ�K�<����@� m�Q�,��xф H�<�@ŎV�$qej#Y�X���E�<QS
"s���3�DR�
�u�p�TC��( � ��%퟊^�Tйa�,c2�C�I�Z�����JK��m�/%��C䉮k�y06k�.E��Q��+�7%)�C䉧]%�<٦,î��� �iߏwq6C�I�I`�i$�ԭs��M�A�[�C�	�� x�s����J�IV�L�C��,U��)tcY�@q
��Â�6 �B�I�nB�(���6o;	��F�1Q��C�9��1���|�i�!��c��D-�Iu��~��mV<�8Vn��8��b��5��d(�Ox��Rf��Ys.`#է�4G�%�"O@4��oX@�=�t&�"fR<  "O~�[NU-p�ְj���>�<�"O�ձ�/N>vivEBD��`�%"OV� d��2�Y	2�K=�~42v"O*�ye�)pS��P ��

ޡp���Z���D�3W�%ZD���Q+�
?D����U8x���i�=�;!�=D���ȺI��p�D�`�0�$%:D�����E#31���ũ�6C�����2D�����T^vvP+V甓\�$���*D�����3Q1Q{��R�TZ�I,D�x�1g��Z��(i��U��ړ�,D�ؚ��	�:ka�R*�462=PC'%D�� �5�áG�*#��ڳ��W2dQ�v"OV����J�|���ۧaƶ7�E��"Ohq��/�4[���p��	'���"O4y.��f��[��߫}����"O�����&�>mI�ݷx�D�Y�"O�!�@�
(�j�!�̀
y�H�[A"Oʁ��Ya�||��m���|���"LOVK��B�v��,߮K�H�ie"O�ȴ�ںȥ�IV�$Y�!�-�y�	Z�l��Թ�-L�E��	9����y���@Sf�\�3Ѷ �&k��y�e�:f�^QS�ء+�����)�y�͇;|P��`h��!�4��f��?��'\r�R%쉺'�X]�bB�@T���
�'k<��6�Ӧ)2h���U�1����'���B*����9QlP#�ۦ�y"�P �T���b��A��aP�ٗ�y��I&�����ِL��AIǋ�yR�ѵ]�б�t#�@�~�BWg���y�� 3�T����+{Θ9����>��O�x ���G�� JI�{e "O�i�#O�>!Vn��	," �ц"O�5�CJ��GϤ�&��
��V"O����Ul��D(aȎ
�|,d�'��Cu>�4�$�N��F�ɻl��� �~�Z�%XM�@�I�&�Bq�ȓK�v�G��LZ�h��ݰ8���ȓSҶP�Ƌ�i�Za�D���"\��:P�ۂ(!T�j�d
m��h��gT���W�P;'��`��	�Ec���ȓ#,�ɢ�։`�rq�h ���I�t�]<�d%�␐?�"�J�r�<���"50�[8\px�ڇ�]l����<a��{��Y!	@4L�Gl�<��5:檝�'�0	n��Qp�<a�*݇hD>��Ʊq��U��-���y�4Y�0�TXE��PĎ8�y��ՅI�T����clE8u ���y���Z��U�ʋF��jDc���y�g@&MQ��"�/��D�8m�s��y��R5�����E��;�QѢ��	�y�`��!z�iS�k �V�IRjN&�y"�S�T�+���S�>�i�!ս�y"�l��%�A�D��+��Y��y��sq6M$��6,�\|)1���y�/�l"B}A�,� ���w�
6��'�ў�OP�Ds�+� <Ƅ@t �$0���'�>���&9)ְ�K �#j�0�',��0�J(ѐ�B�Ԯ)��C
�'����SJ�{�x�¢�S5ޅ�	�'v��ł[4vXɢ$G��R@�'fj�AA��E�`I�B�H&hmS�'�h�*e�T��)`�0}��q�|�U������ �j�
dĹ�RȎ�\q C�	�W"���O�J�أ�ά=�JB�I'f�$T�q� -�jM�RiL�&$B�	"WAʔ8��
f�R�b�"
�!qB�	BC,X��@�#�"������ C�I	_z�4s�P��FdA��\h<yUA���=97�!u��R��K�<9�'�;x]17aEgߌ�4M}�<!W�I��n���Լx��@����c�<���^�;p9`��:��˅�Sa�<9�KH��j�[�I( �H����	a�<� ��)��\�;}��
S�@О,�"O>�ء�܆6��|	�HZ�3��a"O�4[Ү�:�a`d�Jx:B"O=��M�&=xJ��Ԝy�"O��c��O�r�6P��0}>}+���p�O��)�V��e�Hõ�U�M
(�	�'� �:��T#G�-�a�,��<��'d��{�$
-C{�	�M	3(g�W�<�R�Z�(�6]�)�8	CrȰ�,�i��@�<��S;7%�	6�J�4<`�ȃ_M�<	�C�t<�X��דzа���H�<iu�G�\�!a�l��\�0 ��
B�<�p��*ĸ
�.U88�P ��}�<g+���[�C3;t��[Gɕn�<�7F\�My����ְp���BO�<�V�>f¬�M�2m�0��
I�<��R5�>�I��\4=4�)�e�Zn�<I`�]�3)0�!ФM<�
�g�<���J�,(���f��P�%_�<1���=[����}L��e�47O!�!�"�hI '��è]7@!�@-L,MR4`�5#Z<�AI��!�D�z��f$9���$�X�_g!�W%r�;�'D�l��b,�T=!��;9F�-��+ESL~t�2H�I)ў�����ahh��d?Juq+�6B�I�Y�<XA3���I�!0� �*i<lC䉵*P4�lK';���FV�2'rB�>B�D���	(^�] ��/B-TB�I�J���C��*a�|E)ь�sA,B�	p���bG�X�"
Y��M�5"OLT1�kJ���]r�&�~q�B�"O^X!$H�lAZ���ڡ t�ъ�"Or�I$��."�Hqp��M#s��`�"O��;q�[t ���yQāHv"O2��VG�yL.%X��%IZ&Żq"ON� )����"��,��s�'>��f��@HG�[�	�"���$�/[nB��/X�҉ �,�QTA��i�O B剡�`�&��	�Z��gَ4�!�$��YL��	�*ӆ���;�gU%�!�DC�e�!C�@�8Y1V�˕��	X�!�7��1���9 �A��b!!��k����[
\���"�;f�}����P�e�8b���!��[�G�:��Ԅ!D�X �睁I,�bS`�*$7� �� =D�#vh�lܺ��B#��S9֜���<D�h���$��,Yc��$C����" D����.THD�hW ҂�0e��� D��q�f�8��9e��'w�Ε��;D�8��d�J�Fr �������.D�|���2E^�����5]|t��-,D��9f,ԑa玅Y�M\=vb��c7D�T2��;6�$MJ�Ě��R-��5D����L
e���S`W��
�f.D����Ҙ� �Y/`�ċǄ-D����ݯI�llic�V�^˼�i�)-D�t�TDL�������!Y�|�!D���(ȩ z8�A�iNpt��4D�\��L�-5ĪMC�߿�>����$D�(���/x���7N�,Q�ލ�BJ!D�`���)!$Q���M�Yw�	��>D���d�U:cY4TKSh�d�i��n<D��2ТԖWZP�2&���F����0D�� L%�p�C8;��)���F��q""O$ !j�<���mY�8��$��T� �'�ў�OH��[��׷~:��愔Y�IS	�'�4�`c�D�d��&��$La4ȫ�'��S�c�w\�B��_�q��((	�'˒m���տV��	�eLK�g����xgU���̙`/�Q�BY�V�� �y��t�!H�c�"����	��y��qp�4
��"ȂHau��y�X><h6�PנF#d؜��(�y��R{�YYaA� h,e�Ǐ��y��Q�� ����o�43�+���'�ў�ON"1H8M���h9+�v�2	�'_�� �C&��a��"4HN�j�'k���@��<�U���(�N�)���*�u�dsV#,p��*�"Oq>.I�ȓ!�1���TD�1�A���T��X�\թpgƹ+��`#R&ca�Ԅ�2��X '�F��R�#H�-��q�͚�57�*�0& H� R`q�ȓls�cN�֞A�"�R��ȓ-E:��m��Y�I�~����Z�'�C�ɬTz��a��S()�����'ޝK׎M�K�I�QZ�U���'=�9S��4�r�j�Aa����'c."�#$c�$��a��Q2��	�'�j��.Q��Y+���?Q*��
�'�h��Lc~i�ș#D��	�'RȈ�B�w����k��-*	�'�d9%��L��v�F�Y���y���d=�Sܧq��P�]�.�KW��(?
!�ȓ?Ĥ��dǊ�*�^ �Guh��kD,�R`�:q�@��`a0D�	!#�&f�r� �  ք�S!�)D�`b)�P;rx�S^�L�H5N;D�ph�*ы~;��b�N�ERL�rDk:ړ��$5§�lYa�ǝ�بAF�� bd��ӟ�����U�\-m�U�~�T��`��b@B�I�s�H0A��n�P��A�VB䉔X_����6Y~=�uG�A�fB�	�%�~�����v�LA�f�Y�,B�I.7�n%�V��WN�a��։�C�3�8KcKσ.�&���������&?�R (�\�	$N7Fp]G{��'��hT�^����:��<gq�']�`��
�36�|5�S�׾c؄���'L�M⳧�y0|��K�W���s�'���E6D1�VKW�K<S	�'����ּkm����-WUȝ�	�'�Z���JE�Wъz�
�`�����'>�uPp�Фs��ԩEH�����'����!u5�����qh�Q��'�ܼ�@�2H�@e�c�ĉ��'i:�*5M�����Ɗ/F�|��'��2w�Ģ'���*pŚu��	�
�'��,���כas,AЧ@̬D����
�'�Й�%�G�j�b-�WF�C:����@���^&P�\E�@�H7Gm>|�ȓ&��P5EȩO��\H�����T�ȓ܄i�dM.s��x���/;�~�ȓ�3��w��DҰG
�,�Pe�ȓ ��N7z$²�Q�,,�t��(�|�p��s˖@��ė�#X�ȓ:��&�A��p�{�n��%Y�ل�S�? R����lv&,��+�"�0a�|b�)�� mK��c��L$�q��+��B�ɨE��k� ^�'� �i%I�)��B�ɠ%� 8c!ˑ�M��)c.�J|�B�I5*�V�QQ1d��D�P��;��B䉍�0���S�h�)�b���B䉬V��`8bo�`[�I���ݗD%�B��8*�Fh2"��j��U�ড়
�B�I�j����&�!g:����� �PB��|�6��fU�*��YA��;s�Z��d7?���Nf��*�
�Z)p �Ci�<�IL<�0�&!�$!�ȫ#��@�<��k�3<�l��	�bxx����Q�<)���W�
Պ�M�.r`��AFV�<�Ti
��)���x�z��@P���I^�S�OLpD��K�*0��u��_�T^>,R�"O�I�6���(�"���SG��Z@�'ў"~�!#��;(��T�Ez�!󁨑��y2�#!� �!&͊g�ܤ���
�y����Z<�Lu�d��C��7�yrE��h��<a�؊b;�Tj�d�$�y���Q��Y{�*�,+g6���P��hO�Obʓ�?9�f�-4v�6��"0Ra���ۓ��x�G-)].`q�P�M��D/ŉ���1�	矌�E�ȓ�� ����4U~Z��ȓrǲ�1&�аW�6�h�L3�\�ȓU�VxQ�Н-���IP�/"Ɇ�:fVehv"Kdl@,jV
 z��,�ȓQ4��T�+2��i�*Ŗ/�杇�I�\��mL�PYJ}��E,,a�$�'L�=X�
ԟZV��H�_6*i��Xg��)LOL��'����,t��ː9E�Iz�"O�Yq0c��K&�9#mߚ'���g"O8 X��X�B��I�T4R�)J"O��V%Ԭ.�t��� PL��"On���^�VӠ��PIY�aE�Kc�'h��'c%��`fi��i_�؉�BY�f?!��!=# �����ppH�r�A�"EG�Oz�����tI�!���B1�wMX�T�!�d�4e�\y�k������;s�!�D׻,�J@g@��'��H�&L3�!�DK_����C F��f9*�*A�)�!�$K� -��X��H��Г�(��!򤃝8��0�C�x�RY�ʓ-a�!�d�Fu��h���V��ԣ���!�((Qp��Q���m��EF��!�D�2c'~=�b�0p^"@
��
j�!�dH�h����V��Kʩ�R��=C!�l��l�1-6�ɰ�<)!��-u~p�V�"r���!j�;!�D�?X�pP�! KH�B���S<1[�{���ޜ.��5�e�Z����Qr�9,!�$�7�Y)b"T#hP)a#d�g)!��<��"\�To�}���U _!�Ϟj%(��ǩ�Yv
� �»m!�$��bؼԩ�*M�e��i%�!�D��A(��!���+}DKd�B�y!�$ ?�}���
b6��DN�L�}����0h�=W&F�#���}�Ă"D���e)��Z&}�'A� Q�u�Ql5D�@�$�Gk���� �E4dТ�ɷ9D��9W�C^��6d�<,.c�Lg�<A��8Qհ-�d��gFL�ZE�}�<١� }?f�ҷ�W	*�Ƞ��Qq�<� 2��۵�����#Żh�� "O֍s�5G��@����.=����b"O�X0ҁ�'�`!:�+���U��"O�`��zL��"B�קj����"OȈSn��,<�XH!�HY:���"O�źsF��� �Bc �)b���"OqI�)�8-�<@���Zu(X�"O��A!$L���@f=(�#g�'21O�BT�������?n���"O����� e���0̈U�, "OD��T�1��t�U�Ns�I�"O֕��g�Ly6�;E�G�on��p�"Of�SG�$h�Oր%�\1�"O��s�+�����e9��܀�"O��r��++y*���)K� i��'�ɊM%� ����,u�U�;��B�	�5w����(�+ޮ�� ��5h�C䉓B��Yҧ$D�4�Q�+�6�hC�	�1β���dD�y��ճ�*C��%G�JQ3�eE�1^x(��ӯ#}�B�IvGDa���	Oa�<��퐠{�B�	,lA^䰑FS{و0YC�ϲ$����$�O��ɀR���'�^�;(�L���kf@ʓ��<��O:�yqeݳU@�#��~�����"O���G��i�$PϣA1���s"O�ë�t��++I@�t@7"OftZ�&ٯ.^I�� ]B��"O6�p��1B��i9��';��V"OT��C� Җ8�b��G4T���'���X]���qCΗx&A�F�8f��'>a~� �q4��N��Am�XQj��D&�O��)���-�~eTfX�ƍi""O�h$��0tL
تpdE�6��d"O��bG,T8aQhHZ�K�_Ւ�w"On�p�RH)�g�M ҆e;"OL���TY:X��
������V��d�O7�]����\��<��58��#��'�2�'��Մ�^B<� ��,Bs������?�	�(�=
G�a��X3b�d�6X�ȓZ�l!�����j�8����_�*(��
�|���� s��]�5��?Z�p��d��3�k��V�^
�nC�	�c�P@A�H�yS�H�v�F�)Gv�FR�'>u('�	����ͯIJ�)���O���d%?A�땻I�H1�r�s5.i��(�ޟ����^WD���Փ3!����!(�ޕ���f�`�j�;<���əi����ȓT����M�}�Uf%�@%��'���
s�$I�uNZ7�\��ȓ<5z�2�P3 N��w�t�Ih�'��IDy�U�n�.q3qo�|h>���c��D�!�� SG4I؂σ�KZ��@ݓQ�!�Ƭ`���F�&`�"q`7�Y�y�!�d!qH�x��>ax^��MF0-!�d�&�����29e�!qP�ĸ%!�-Jhu�2f�/)J�|;DD�c�}���(�d@��
���;7*��T`��j%|Ob���&o	�Y���H4AN���5H#D��x`�.}��F�H?5���H#D�̲ �X�C��ak�JLByF&D�P0',�c���F(�$б#(D�� B��#F����,sNtp�i&D�
`F�F��`FD�y�0���d#|O2b���!�	V|]y��ߩGv
<iO#D�� &��k�FF���ߩaG��0G�'��B������TN{(��`Ƚ!�_�� 5�7��\���7@��!��݈+	�B��!���s#��V:!�$~������Dm��(��չq9!�d:?���ڢI@�&l�K�/ !��G�N2�@A%�x~�����~.!���@K�͐:j6��U%.!��Vd�H��f��Mal=�A��72!�d�&�!s��\�7���Cf�.!��� f�bi�Wp�R��!����
d��@ ���'G�M����L�!�)Tq�b�ʘ���hϔcT!��	!v4�1heNɺ.o>(!'A2?!���*�t\P���#P�H�V&�-!�$��5U��2CCJ�u�j��g뇘S|!�D��Q�p	�7*g�NX7��"�!�$C,�D|�c���,Eh1���!�!�D
8р��f b�fd��.�>ek!�D�/�*	���'"gٱ� _.<�!�DՄQ\d
�a��HRމ�n��!�dM=z�`㯖wI�T�v$�"zD!�$�̈-d�Ӯ3i��E�ظb>!�DЦm�pMZ�eo�@*���W&!��,,*�"e�Ȧ��a �\$7�!��K�[ٺ��n��p^8A��?�!��J�
�Ip��.RD�JFސM�!��;bt� �[/U�~%�s��<�!�$�9��j�I�!C("h���!(�!�d�+�KA�<�6u*���"G$ T��'Ȣ���º!�S�N�On�E�	�'Ȁ�J����m�+C<��x�'�l��%�8b�z��7'W2gݲ��'F�T��G�rMF�����5f�L,"
�'�h���
��]�rǃ�S;�*�'1X��,O�W3��t㙇J\M	�'�
���$�w�
Q�A�Q5� P��'fm�Uoԋ0�#6FƏ2l���'���0���=G���0�t�&�	�'�6Ȃ7�R�#�	�	i�����'ht�� ��\�����6e���
�'@0�H�j��I&���^H0	�'����L.J#�t9�K^1\J�M�	�'�j|Yt�kB)�e�UD��
�'�> Y��הi�b@���8���:�'׈Y�*�0j�.�g`59 ���'e����f�;�Az��V�298,�	�'�q3���80��w� �=!	�'�"q�OI8XrwG�7e��i�'�j1@ �������O2x%�t��'U�шA%�,*�H� f%U�v:x5��'��A�$	�)��mإ�Wg	�'^��rc���`�����\���	
�'?bXꇇ[.�h��C0Z8��	�'Rtb�"��y��a�D�M�Kw��	�'�Qk�#OCLqѣ���B[8��	�'|V\H�)�1Y4(rjU7= ��	�'��crH�`�$�ZA���G��9
�'K�JP�,#bhR��X����	�'�4-������n���!�N��'dJpY�,�%v�N�`�gM2M��� �'ⲬCf�@"����f�X�N`ځ�'�X(���"@�XBG��YU`�
�'6:�� �� ���ЄVo�Q"��� b��+L�fb4-��K�l�X��"OV��'��."�;�J0��h��"O��`���W;8�NIc�Z�: "O������w��x�W�Φ���P"OV}�r��m�a�f�S�%+~�"O�9p��0� �Q�A�~l� �"O�ĲD�+ǈbC��.Hl$�"O����ؽaM��2�,�v���*4"O@@ؔ��6mXp�˰!M�]�zQi"O�-��,;FR"��A��x`@0�"ON�	ţ�)0�mi�J�>Q�p�w"On�	BD�*�9��	�O�j��"Oڌh�$�|��̺!jՍ�"��r"Of�ӗL܁�
����X��V,�4"O��iu̎�m"�Ā3 \��eB�"O������"����Œ%`��"O�e��c�,�䨂���U��"O�pYc'�j��k�2�$ k""O�tHҌ�"m�׉Ģg�0=R�"O� �t,�=C�^�Ӓ(�Q�~��"OZ��Aʑ!mP�RA���m�l�
�"Opq���U9D�⑫`NE�L�V�:%"O�P����GL���P u�\�Kt"O�݈�� <0���/�8+�\`��"O�H�]�� �����zb�H�"O��j�ϲ-�$q��B�$V�x�"O� ��+YK�dA
��"4m����"O85󁭋���I� ;�t��c"OJ� �i@9-��=��ŏ$QJ R�"Ox�4��mNp���A�=�JI��"O�A#�	�P��ɫs�ټ����"O��x��!U�vnV)!��T�R"OZ�c�Ȇ?s�ݹ֫A�p�}��"O�@�!��{����ӖG���"O&Q��#�ox���9ry�S"O��P<ZqhX����&<�Ǆ#D�Đ1Ϟ�@�0|ړ�=@����q�6D�h���J%;��0+����T�����i6D����_+�lA�M�M�xْC7D�`A�땲G KH�8�蚲�3D��q��:2�������%Y��$�-D�d��NK	s����a΅)��� �/D��z���&�*�K"j�66�ʽ�v�.D����R#��`"�ʃ�X p$�)D��`�e�S�<��ȶ �~ &D������=��y�gұ]`�I��"D�ljAkF= Ԅ;�IP���i3D��C��X6���q��3�~H*&�;D�XB6Xc\N��p��k��5�ƃ;D�t� ���GU�(�*X�0�l��CI;D��PtkR��B�����-�<퐁�<D��aN�3n#Th��D<Q�qG�:D�<�Th�sS��iǅY%M͔M*�9D��a急X󌘒�۴�����#5D����"�'F�iA4�2QM��1D��q��93��flNzΐ��¨/D�����l0()9q"��`��,D��J	#2XV�����M��jP�+D�����	{/�P27Iݶ6p���+D��9!(Ӳ&d���o�x��0�*D���b�sI�m��Ę%n����@N)D���7
R):���c�L#��ic`H-D�lb@D�/�H`�EOI�!�iK/-D����8.�h,2p�(9>��R$b)D�� �5i@�Y�:���ȕ<$��m�t"OTx@�%ˇMɊ�(SN�R�a"O�oB+6Tz�ᇈ�m�p���"O���`�Iל@h�HߛM��!�"Oj�p�$� ~�@yŧ)m�N��#"O IP*ИZ�$��s�(o��PX"Oƴ�BK���m��ߦr)�("OB4ȴ�B P���p�ŶFl�3"ON�!�dA��̰Ŋ��p.�)""O��p���"[9Α��C�;6��u"O @xČ�s���!c�Ҿ��p"OF�*�(L�XD� ��c��&"O�%O~ 4Rg�%.�tx��"O�|AUi̬Pc�������b"O܀cq"/�l�!Um��]�(�"O�9�����y9��ӿM+@q�"OLҧK��gnn���N��x'��8�"O ����c��imO� hh�"O�AIE.H�.|K6@?GWv`��"O��C�D�y��Y2�U�"�"�Y""OB��h�M�[�BN�N���Z�"O0x���t޶X�F����>$��"O���l�#S;.$cە�*��v"O
��_%��RW�	]tl�B�V]�<	�+	8�iq���Kb�scNId�<i���\�ȣG�[���c-�\�<��c��?r�����?m�H�U�<i2�J�.�]���0C<(��	�N�<�i����42`��,N/�A�K�<IV�ӱhx��a�;uAI�<q突�f3|�
'ܽw6R(�0OB�<qQ&�.6��qZ�a��_4K�)|�<)�O�;>z�)E/��\�r�rR�w�<�dD@69*���5H�N��ҫn�<y��9vuKpEW0
|�BRm�<Y���2 k��13�C$�4(����M~�d��<y�y�����P���'N�}H��Y��M�*3!�F	?��q+���qA�(I!��
�'ıO��P
�������/��� 0,�NZ!�"f&P�3��Vt�Lp�'���I$>I1d�l<a��L��v�.^x^k��\y8�`��4��'�T��H>,,l	B�S�Z��Q�'���"ѩȩ
����#��Wr��IO�l������-��3S�����Ӡj�1�!��ЋE��1O�e��E�� 2v�qO>����6R����jJ?u� �se�@|��}r����b��*���!B�+a&Ɲ��1D�X�D�֦Q�u���2i�=�1*ړ�0|�u��,���x��
����BQ�<���.�Vl�U��!X�N��e�s����?�c-�Q�TT+�Ah�~I��3T��S��Hj0���e��yLe{F�1�	X}R��c��QN��F�&}���2D�(��KD*M��}a�&ãe*J�&2D�����&�T��:w�u�Q�0D���a�����,H�j�&A�a�/D���'�ݜ^V,\�3Aπ\7�yt+D��;��{�TS�'�0D���eH(D� zg	(%�N�JaIwR�B�*OF	"Ьʋ�4E�R$<�59�"O�0(q�V3s��%��ȺQT��"O��!t�?׬��'�"��e�A"O�ْ��G8{�d�s4�R�y��P:�"O&)��@ՇP��L��lN*f�zi�r"O� 0Yrj��6$���մYlz�"O�9���7Zk��i�*�88P�E��"O�pt��l�V��RJ��uQ�ف"O�y���$<� �B�؈[�� "O0��d�Od�=Ґ��s����"O�$Ak_"�aH���Pv؜K'"O&�RF� <j�Xs@"��)�y)�"O�y	 CզG�1�G��#�	�2"OdY�G��	R'�Pg��T%s�"O�M����>EU��%D�0�*ͺ�"O��
[���hg%��hgh��##��(O?�I�y�RMi2��~��k�(*&nB�ɕD#&�QD�2p*���A�L-,C�I<6^��閭&: �x��ފK[�C� "\ �f�<���a��'�C�Iz��z��Ó4��J��;%vJ�<��T>�b .M�W�zx�Rg:Tl9�b7D�:e	� phL�*uG�b]�"�7D����Zy��ya�@�!+���0D�����(j��؟Y�R����-D���"I
��@��3��|0=��B-�O�˓nR(!pցM6P����	��&|^���-�<�'��
b&>ԡ���V͜@��(n9��Z�e�揁+�\��q��	*�D	�`"X9��ġ1�8��{�,�h�Û�x(� )��U�+kv��W4�	7J"lA�G�2t�p�'%B6T�C�	 .�\�P`��3�pD��J���<A��T>�R���n�ȓ*B�n2�7D����$�K	�`�2��=1�h�b�9�(Or�}�+�a�a�8�$��f�!9�TF}���6$��p���1$*�eL� XV�p�a~��ҥs��Q�EA�Y�r���형���&��|j�|���)�����ɮB!�$aE�ސ�y",�J�f��0�XU�|�w�@����~7O�c��'kR��Bg����L����;Xt���DU`�K��&fj�d)ӇѴZB� ��g��h���&a��h����Hn��c�k���ay���N�qB����߳X�zIqG��)Q�=�N<1�N�>E��'�{�(^kXm��T5FY����'�,����!;�9��E>��@���'ay"/T�ΌL�ҥ�,�RT���A����HO�l�@�|")�HT�ȫ�-X�xS�Ԃӧ�y����hG�:x��xqc'����y��4�SJ�c�TC�}9w�>�<B�ɭ2�T]��f޸�J��)��?)�C�I�z^��(6��%N#�<Q�W�3�����\�q���xz��̭'a
|���K�yB:�8R5��=�O|b���Y�Z��wF '�r�iU�	5F��O���:W����Rɝ-r�t��+28�2C��<E��1��ب2P"�8Ǩ�m7�4�@?�Ob��Mkc���o�ڭ�u�ơ>���1bE�<1�̥D�<����E&[$�Kg�N�<I���������'@�X+N���̜y�,IQ"O����@ڗZ�*��f����uY��d"|O���Nۍ&d)1k�m�t��R0O�����.K���7F�z�ơxAF$��z"�^h̓O[ܫ�	YU�@Z!��~3���	@���H�d#W���8`e2*�>IJ�(D�āX''Vdc �A���J"*¿�y��-tJRBh^  (�P��I=��D=�S�OD�I�P���6�	���<�����' L�C��Ui8�,���ڎ��{�'m��)ɉ}��]*�&)������� �aܬ]h�z��RD�0�k"O^���[�:��t8���I�~�%O��Ⱥ<K (Y�%�7m���Q�+���Z�'�1O�3p	T���˅�N9(�a
�֢���}��~��	�t�Z���l�-��$����z�f�	��p?�q�ƨ��� �{�\����R?��g����'����.�~p��)Rd�?\}F���'�O8y	�O&�+�<?��u�ö0���)�S��y2nQ��4���@?
����+N��(O��)ů2�':�^}o!,J��x+�Aӄ;�LQ��x�Z�l��:��$����d�ȓCev��&�0B�Nu����bE꽅�2�D�N� 5�!r3C4CZ���>q�����lJ�LT�ZQ��-�����S��y�&E1@��cp�̮Zv~��Q�ϼ�HO��T�>�R'���S�(U�t#ϴ!!�d�,��Pr'�0'�z�s��[�!��P>8l��H��uZ�����N�Q�,D{*����M��$���Vg�
��r��3�-�O\�#�nH�_��Z���5vޠ�zȅb��H�:�	i_r��*f�v Z���;?B��6�̙��!z���c�T[!�$�'ўp�G-wb�� hƳO��(I�eA�<��_,H�D��tK̬[=�u0"��@}��|�C �g}�mW*]	�T�5�Q, t�1e
ߥ�yR�P�2Ƽ�h��X�t��IMX��P�)l��w#�"K")U>D� �#/͔5�7�у4�<9vi0D��h����*[�1v�Д`nV�Q��-D��a��E�U�6��@�(�@S�6D�x!w,��5�^��y,���a5D�,Ӣ+K�S.Ĩ�%��nF$�!��>�L��==蜹ca�ϗ&�,uB����Љ�Ɠg2��J!%�!�DR�O@>e9@����K��/|"1����� ���:\s�܅�#��� N?=,m���0K���ȓh���함V'�lQ)��!�T�<���\+v�:#���MF� \Q�<ѵ�Z
.d8|S�lј1	d�`�K�<i �IM0�q�ԩ�J|�Y���
}�<9w�]) [��ÀɊ3*��Y2�"]}�<q	�o6�IAMɯq�K@�`$B�	=V膕8��F�`�d��B�Z;(B������V�y,D��sၻ��B�I�
	�0�� ��wjjY�ƍ� ��B䉕r㎭ҡ�#�
Y$)��l��B�I�Nf�0�V��,e���W��5B�ɯ<�&�,� X��Pa���-�&B䉅zD��m��-�p�R�%	�O��C�	�/NH�@R$�"yz�h�k�kۘC䉛p� RB���A5������	1��C�	$Z_$�*�̝q���v�,/��B�I�#��-bdK�3.���㊝F��B�I�z��h�@̰�(��R�F'�"O�,����P�`���_)GSXm�"O�䀵�_3(���/:58�@�"O@��䘳n��@�.Q/Ք|q�"OfM	��M�U�@IM,l��(s6"O�m��T�"��,)�
M�|h�"Of�ց�.��<�g(ɒ�D�!"O�)�qAS`^ij��OS���"O�XI++|r]���X�D�%)%"O�؀�*�b���@�
Z=�Uà"On���A6}c�	���++D~�"O� ��r�Q�wl��qƝ�E� �"O�hg�m�r]@ф$"���q�"O�4k�]2e�����,�q�P� %"O���K�}����G���P��Q"O�A�qLի%��d���	�l���"O�KQ�'y)��_�婦���l�1O���VJWk��!3�ڤ~&��s��77�T�s\�7H̃p[C�	�Q ��ŗ���$áȳ?pXB�	)T1˰���~ a�N�PC�	�K�>Y�f
��9�J��/��2C�@`�y��X�%���ˎ�4wC�ɴ�D�����I0����:��B�I�du`;S�ڙFq��^0Gq�B��>��*�����v���A��S�'��a�୅�+�4dң ń��
�'�.�JY�?[4�R�& �X�`�'���Krb�bab�2p` z?���1|:�3�"O�nj�В��C�s��ņȓ(Fp�fm�w� -أj�(09�ȓ*�D�[��>oT8�� -	�DH�ȓ2��(0`�&fz��g
ȥrb�ȓ��}P֨�4�����5qwR	�ȓ~2}1� ǐ9)T�����2,���V-�-Q�"�p���Z���,]T��!P��`�M�@����e���`���&yO�u�i�`�%c����P�f�p���$G�2q��Qu�܄�)�<����վ2�vщ�i�H(�e�ȓ-*bd�B*N=l%�]y1F׽
/d5�ȓ[�̓�́*C��$Yc�P�zu`�ȓ���ʡ���x^0�H��];bH�P��s^R0�.	9�������9�>��56�������  %�0�ȓA�`�9s��(d��d�G�'�F�ȓ�ɞV�d'��lʈ�=�g��6����'��aK����He�=`h�ȓ@�TTk "
�E� ��c♼m��2D	%�I�K_#|�'�^\�uOA: H96/Сzs����'FxF�u����4ĝ<u��$����bn����	�>� �l��SPe胊��b����-�$�aM�H�A��'P?�bB-���WM:D�x1���f��5f6OV����e9�ɶL\������IH ��jČ o��ABY-!�d(e�-c�ȁ�3Z�d�F�H?AF��B�{r_����	�/lƔU�ޫ!�(i%��2�FB䉇3��1��*�=��`P�]H�y(�h�3��?�G�S St�heAԷ,����A�BD8� ғ��}}�!�s,�$� �RQ���:�ܘ�y"�G�#��(KPK�J�������OT�a���稟|P�����
S�\ 	WXS"Oh]z����{�4���V*:��r�����գ�{��9O��֎�Gyұ�4�ƥ~!���g"O@�P�+��yR�S�/�A�c<Oƥ�!�P��p>�dV�JK�ur��Y�Y]dR�Zg��҂� k��D��D��ҧ��Jqgi�!�ƖجQ��ʢ[f4jD�Gi&��@P-�/Q?[�ҥ���3R��3 �h�*�c!D���Ø���"��S4	� �"�G�=.:�E�����'���	��G�"q�/�P���B�'В̈U��$c�%#����i=D�D0v��]�bX����*��H��'D��RUN�5O�J᪐�E�H$�,���+D��
�����ɈB�^�xB�s�-D�@0&`�*)�Ȫb�_�2�%�i1D�� �t�1!�~��dg����
"O2����0���{��|���:b"O4���^/*붡a��C��@�s"O$ �EC���:9V��q"O�Ջ�^ {�^E`үF�z!� ��"O�I�vO�
��PZB+Ž}f�ұ��^��P�Hm"�4�%[���:����͊�b���ȓ5��5H1Z-N䱒���Bg��s�(�A��'��x��D���c�X`�$#W-FܙU�'4��׏M�]�v$�����F����{��h�5��"O̆�ɪ@�	atJ	$.�~�	fYi\��	%-�j�Y�NZmX��$�|#Q#Q6g�6����ӕry:C�	 ^Q��y�3$��Ĺbd[�*�O�Ё��]�2)�EE*�d刺(�BQΧp)R�� ZqD���	�T�H<�ȓQ��!�����Z 4Mi����-.�����lAtyҌˊ2b@��DOs����f��]�kPzkG��H�ތ9f��?XvC��/}��I� �������%V�|�L�j�����K��O]����#�xFLh��ʸ.�x%�F1<OB\X!�K�+�l�Nq��Rp�A�$n���C�J�;]���.D�QP��WB���\�\t�D3�,���^r�Xsm̑'�#~R�o�� ��P�L�{���wCFT�<�ᮇ�4+����œ���ɨ��p\h��)}BO����I#��I��E�f�4:���]m�B�	�F�a�Sjޢ
s�ID�J�`$`چ8��!��y2@�8��%�?ɓ���x�h����}� p�3�M\�<�T+��}LUÓ�L�O���<�����=�̈/�����1\��T���M/"� ��ƙ&�a{R�� ;CT����b�j5�I�8��
�P(g�U{D�Ch<�� ���1�&��3��Ħ�y��[}R.0?� ]����:��!��Ʌ�%L��
��Ѧ��l�5��z" �5*��$�'�d�P�O�4�ڸr�EG�H�f`�7
b��{C�*eMR��K��(��	Y��(3` %Rf��c�&���	A БQa�����4D(�lK;H�`���c�L������6���ô�+i>%��I����2+׀;W����@�9I?�I�+�S :S��0P&��D�Y�5���M+4i*�3�,�PA���Px��ì`�t2����6Ԙd�4j���<�Z̀��?ac�	�H���¯`�t��2��Om�"ɝ����B\	7�b|�ד!��;�-?Q'އQ*zHh�@ן@��eN;|�Qxe"F�sd�!Tn�9Q���2�O���M�Cdj�#ak	����J��5~�V�?7_
�����+P�7I�`�R� �f՚!ɷ�:�a��7)�8i��W.|�`��X��>p
��A�Cg�]���R��������,[�D�dA<mt6-ٱC���tb�!m�98f�݊{�&i8�!8.�����тa�����- �2�R��S:7>A�$,z�� m��8�0�NB��w��.�.�
`H�; 66y�Ĕ�x��|���EIH.8^Lx�wCN>%����^u���4o�yB��#π�vT+�,�["\p���o�58�g ��������Ӳj�-x'�u���@N��	F��<��έS޼WX9���#=#��2EM�s��M���ЉE����bO/V�ʧA%�B�Y
�N9s����^w�Us��΢>݆� ��1b^u���4d��$�K<�$+ϻj�P�����$$��2�n�)d��-�ˋKH��1 !�*v괌ֈX�?��Tdۘ���
*�u���.(y���0
'���3F� �P,�g�-���D ��;�|�]T�
 L@ v��gD�}���+D)��2���zM�|���\�C��*@��~�5��{���d9����#��4��JO����:bͲ_;(�1�OF�Z�V(8�~LR�*I4�|ِ���uĬ{v�I*u��x�S�=��C!�L�dR��j����'O>~���*wމ'EXa '�O���s��CY��ߴM��	Ѻy�L(�`��}쒀��O�����Z>�;�� /(<��	=DѤ}��AU?gF�M{�B��~ٚ�kD횦hR�cv��'k\�s.Or��Gdx���g(_>� YR�lF�~H��'��z���+�'P��I�z���	��a"eL�	xEr�G�0 R��H��6͸�T7�ɳ/���?�Ox�E��'1&�z� @N3Q߸��G A�Z3�+��43�-K�{ ��ŧ0"�`7� d��y��~���^E�z��_��@��e�eX�(��W�Iʩ��NKYr�V�5�b�H�l�	Mia�FձHb�K#
V4��đd@5ی�L>!��B�8d��a@��J �0��Nc�K"� � �"�*�D��K�H��1B�mJj#��Y�� \9�Ҵ� A߬܅��aڎ��S[7N(H]Q�N�nh�,8�MH;8$�'i��߮A:��Kt��i4��(��R(.Q:�!`�H�J�<B�	'[�虆���.1ƨ`�I�}��$�h����B�0D�l��<}��� �l�ǖe[��ƏE���K�"O~![�*"]����tH�!�l�얳7��B ��RG9�3����x��c� i~��+�쒯PqO�RV�׉����͋��Ii�Z�m��}>�5zCb£]���F�!�0?1�i#Y��f(�,	�jq�����q��9�M>��!�C����AnY�F�>I��ǩ!�#q�V)��"(Bh<1�"�vЦi���*j.�7e�(+�uYw��?M�����1}Q��>�;���R� ѱ�����(�57<O$���
��8��O^̸�'�W�����f0^6�5�%"O�� Œc�xYYq�T�z�:kW�|R���"!;'+�{�Oed܈bL�/?���!�ћP�\`��'��X� iVd�8�(�K�L�v��S�7�b�'�J�(���>٤D�:z��;��ڬv^�T���lh<A'��9U����YRH����_�P�fT�ȃN_��lZ8V����:O�i�K���'�Z<�t��i$�$�t�C�VM����h ��ԥB�UI�6�Ӌe�����iD�p�� !��%�<x����)�D6M�%�a��6LO&QS���5,r���	�`޺�J�|��I�cٴ�zA!R5��=k���B�t��,(	ys�W7;irQ{r*��U��1x0Z���'��x`��
����$� �jv��� e48s�4�������is���6c��8��_>�a�{���'͒W��Qа%�,|���j@�:D�DH /E�|����v�d-��i�.�Dh��=M�XW��1.��E@ M�/D�~�I�O�	�0��l��f�*y�Q1�(&kP����Y3����u ٬zw.�(Ebwu"A�!o�
^�ٺWGB�W(�!'��Tx�� f�&4ܬ ��!Z9Dl�7"�y��X�BLk�}���2���݂{U<�b�C��0��b�/�Y����!��;6��y��a���ӕE��I�pE�=�'�[�MU9�'則*�Y:���in��7ȟ�94����(�yr"Һqp�UB�*I�8�(���-?% �3w�Y&"����-�"���K?!�1�;�Ҽ#�����
�%Ff~a13{�}b2~*�Z����L�0�>P�G;�1�(_�*Ɇ!s*� l�#�!<O���>U\� �o9��CG鉺8�`2����p�ߴ��{7�^C��Q��dJ��&M5&/�I+�=4�lJ��űHO2�3ү��2(0�Eh�:�h���}L�m�w�O�dj�a��JM0b?�� B�2�qj�E��ӕkB mDC�	=���i�7�b-��D�x��� h����ױ?�N���O�N�a���c!#�,e�$�+�딓jZX�k�)�O��`gl]�x p80�D)*��z���%T(ȁ�҉!H!�$N���m0�,�)wp�hQ�c���`GSj�.0AƠ4�S�	�����̈�,��0ˤ�K�<�~C��>$���{��ρAрT�`�B�0����D�4H��H���)�'s5�	W��)h����QJ )��`�'e��J+���#�g2d�,O�#c�C3�y�� �\ w�^7hO~��Ad¨P�
���	(b���@�<�Lʱ�_ c5
�7�im���8��thg,��4�`��#B�h�F}��̇w�6�E���34���k0 Q4���y�zu*1��H�Y r#���y���,}'���*����1gX-�yr�"Xi�č��0�RA�E��ybDՈվ�h`#d��`F7-+!�ą�F����f:O�@�Y��&!�DW�

�b4�7i��l(5fD!���B� ������x��!�"-,M!�E�\-
8Z�I�brtT�$k�u&!�<k���ւ�M�d�ۢ�Z!!� M6���NѾQ�� I&ݚ.!�!��A�+��2�vq�X�b�!�$�&DҔ��۲h�r���D�!�JT�pS�NL.���2pH�i�!�d��][��ʱ��,Ыq`���' �9��&\�]j�%F�`�N�c�'،%�'�3J�C$��.5B�1`�'���SD�]�\�F��v�Î(TJ��'X��U�^���e��y䎉�	��� ����&d�r(�(M��]�6"OL��g�9t����Ũ](R����"O���`�٤��p���(ɖ=z�"OX�i�oO�_nQ#v�!>Ύ|Q�"O��q0mO�+Y\�1�6��uȇ"O=@�W^9���#� �YC"OZ�YFn�,,mQk����Q�8xe"O��h2�A2rq> h�e�7�fAq�"O��a�,\�G�F"΁e�Djv"O���C���li
���D��i��"O,ܸ0bL?#�LA�Ǐ�0_w��c"O̙8�딾l�q��I��_۶�:p"OTjS䛏/\ i��n�@m�%�@"Of("�M�Y���RM�	F0B�h�"O�k�
M��%�Ϭ�Mر�'�yRM��!�V���j����QR�y򍛪D��X�!!  9b4A�OƉ�y�[ў�����?x��l�f���yR���=Ɋ!Z�E�F ���d�'�y2��9U� x��J�R�)P&��y���'�f�s��M��� 7Iˊ�ybNA�N
aZ���.Q��h9� �y����nl�DΰY�be�A-��y�jY�zoH�+�U�pF��y2N�Y�  R�c�;;���ش�
�y�`U�1;�5C�X>E�0�-�yR�4	���C��@$��c��#�y�b>I���OĠ~�c#���yb4!�1DADۂ����y��$2�@@����t�`�+EmM��y"$
�x����gF9+*�P�
�y���3Hv�Q@�(1��8�䄅�y����z�e�.P�|�q \/�y2i����46�^'���j���y290�	J�Z;	v"m(�O�*�yC"����%�K
B+'�Ħ�y��Y�}26l:������a��K�.�yBnT�BL�yzW�E�Ҁ�����y�-�'g�2���i{FT���Z�y�&�[��܊�,Sx���Ӆ�yr�I
82�PJ��H�S�d��Ao��y�Νu
096a�MưƥϚ�y�B�����
)�!p���2�y��\��)���U`����4�y隮H�q���J�Fu8db��y�Q0NI
H�t)٧��!2�d���*�}�d#� %0��A�]#HhNi��>�\��G͜4*�R��4m
����ȓ<���9���(D�D%�"�Y?��p��W�15�R9M��}yu�,z��ȓ'�TEi������0F�C�tQ��ȓgXH�5��TLp�w�\6�4��ȓD��PP@M�[�PXa2�҈�XP�ȓ$��}��j�b�\����츅�F��d)ho��`��<n�"e�ȓxÔ B�k�$2XY�E,*V�ȓ'M����R%U�(,�$�;y ����6h�����R�8�+M�[V����j5�����?v�q �ج4�:�ȓlH�a"d�Q�w�R����T0.Z<��+�=��	R&4o�i�,X�ȓ)�X���2[W��@ՌH��-��V�by!p��8�R��ʋ	�����������to�Ui�n8h��S�? N�b��P�@F���p.L�=���i�"O|��G^��r�Pb�&W�-R2"O�!�.��cs��C$AX>���A�"O�%2��r����n�(P��$"O^G$T0v�V=�'��'=F!�M�F��ܹs U�!ߎɱF�&?M!��J�l:i[���$5�Vl�(W�!��9Vl�r���]����8aݼC䉎s	F�#D��P~T����8��C䉓,v��btf�p�q���=30.㞌�g���`E���<nq��9�ܸ>쌙����y���S{
�q&�H�ay�m��bD0k<T���PZ��E�b�>�ho@��r��d*z���� ����Ɠ@�|�C����OR�	��]�s.�!Z�ܙ2��`� ���2H���q �4^�*�K��H.����D�5]�>�t�I,���	�<ux�Id�\=Hs��j � �=��B�I=R�	�E�Y޴㄄[�Ŝ�Oڠ�$Z�Ʉ���8�cC���A�C�!���0%mŲ]fZd��f���(�	Ų5����xxDV銎7�Z$�'��-����>�aU�<:������s�ISM�Eh<s�
v[��땣ͬZ*$X0��S�xr�8w�J�X3�غ�
r��sGHZ�/�z��s�A�7����ɣ-�j������
1��ϓ!�.�R/�ov����Ɏrf��ȓAxv�k&�(Q}� ��B~ !'��PC�"Ay=+�'y�O�T��uM������<��y��';��:w��b-��D�0�� 壞,q�L�O���3?�7��:#�>��v�W*� �����^�<	3h��/��y�H��X�d��0�P�r	`�a}�W�1�"�Yd�r�
 � �M��y�/�7unBiІ�v 2�2ՄÇ�yb$�>R?�%�5�W�k��UI����y2#���Ԙ����g��0��h���y�����E�!a�  �pSQ+�y2��/��}��3*x������y�g	���2�O�++�Y"C�	�
�A�t�Q���M��+תa���*�@�lޤw%���J:�Ʉ�&nl��\'�0��_<S����c�v@1��^�8����\3:�n�ȓ� �T�Ӛ!���*�Mp���	 �p�$����6�Q$� �~�`p��
�t]u*R�)
d��IS��p<�ȓ+Z}����t�/Ö
���D⡞<�&��x�!�!Z��QK�x򾥺�޻W�F�EOh�5\�A���FO�|=VI!]�b��@�x֌�O:�(	n����2%����3p�8H��ȶ~n�K�O>%C7�ȶ/躭�0��&"W<H���2uQ�d��ۺ
g�l"b���S�˓o� �I�i�TL�TI�D)Z�I�I��B'��Ɇ�	�M�$H�§ Kޥ�u�(l���huE #CG�i���^�o}PL�����D�x�����1��O�8�"5:�z����!�
(A��>Q�iK�@3Rx��ѓ�N�Æ'���ʧEM�c�DƓ9�<vF�
,|t�*Ԯ�,0C|��a/�O~��D
N�X�δ��	Y��V.e@�ءT��GV�X�Қ��+{,�k�EQ�:�N �'Jhy��J�+1(���V'�v�X
O�YA�
�gK���ө�5��a�>#�xQd�8��Xk�a�![��#*O�D��-��k�bM�O��p���tt}(3�����akq�'6`́5A�?`
��G�m"��a�̣PxQ��*�!L>�"��[/pt�4�'�(���դj���E~�fE���xj�~;NP���/��ɉ�b�����Y�������LJҀp�_>�r�b�
�����35��Qg���<O���a��L5��آ�� }�hT�r �>T��h�!ώ/��G��.T��O��ȊQ�D)k6�Kc��1��Y`Acu`�R�f� �Fd#�%:�	��1R6~�i���4!��(s �X~�'CЩa���9 �� |���P�ߤ��\�$�ͯ2���ҿK~i��	�[c6$��r�|B��/���C��(L��hG�Kg��\�R�z���L>aCE��z��a�TMź����J�	LǾ����5Q��F�d�Ho�? �}�q*ϋLՂ��w&�"��ac�ڴ���t�'O�Rc,�?�F��敨��@����7�&�'�D��O����J^2�N��'�(IC	��?�]��*V�t.I@�'ڪ�;�(�7i���`ƢY������t�&��S ~������I}� ��y0 ߾k_��r���TM�m��_:(�+��¥.�v��p*	m�����B|��T1�J�C��L>�f	�5 ��<�BEM2{�t�xT�[LܓS�Z4��&�K���4lDA�h�ŀV�t��%A�O�H8D�6�O�IPBKA.3t�1��X�E�l;��'��Od@]?u��͘W�V)�O6��$�/k 	(�N�q�$���O�DH�c�L�:!z�i� �F��;(��	�"G�Q�����O1*<�'�:�2��s)�{����;�>���i�x��c�ܙ� d��IB"��1�`@�ȓ: T�����'�J�aSJ[��9&��I#
Z� �%�#�*e��l���1;T�4��d��-�C�I�3�~��愕5Lo�4�pi�<h1D([3�	��I {�v���O��A��HP���c�C��ɃO��q"��"��<���_��S6�$�XP�� ڛ��w���ϓH~qQ"`;�I QQ�wC�1el(�t
`g����	2mx ����M�� 6�`Q�6�@��|ȥ��oz��H󊖕�M�W�� �|}�
�6�&��'��xA$EG$ןH��$�@�K��psoR<z`��g�5qEp��$jЊ5�,�#lT$U��&�S$��F*W���x��7���$!85�~JD��zi��i�,�B�T�G��� �,j*A	�	�|�� ż����?p6��#�+Z.�	ХG�<a�l4n�����T��څd�6\;`f*����`s�A`�,�4 l���S���_c���f�H�U�lx����ɛ]d�4�u��(D窴�c*³3t 2��X��jT�
*:�: [��G!��<Yvɠ)زdvfA0NȴȡReRe�'��|�R�ٚ �2)�rgʗO��u{b(�U�Z0�R#�:�H����ܶE��B�<@�z�3bJ:6j~I��%�J�\˓(�Ԉ���B�{(.[UO.4֐���)�|.e��e�0C2������!�d��Y 9�S�X#�$��,�:-���UB:��1LR�[�\���~bD�d�:蘘����5=��Ș'״����DڇX��a����,�&��#6,×dI�u⤠!��2k�t���S2M��󄓰[��8k�c\�0  �odў��t,ּ.���7`�Ʀ�Z1�B�1��ɲ7昢?�z�Y�C�(��A?=b��Doc\5Y0(�'��bd˸�yFՒ�fQ�0n�o?��63��$��4F 8H~�S���8��)TFJlY!�D�N=���"��hՔ!�@٦?V�˪>!��і��C�e֧A��v�y�ka�@5O*\�b����L����|���Q='�r8Y��D۠��'B��2�XZ�O8��a�����X�׀X�Sx��C!�	�L%k(����P�~
�N���2��Κ�jn�Hiq�Yw�<�p͈$@���Ce��U�l\A���ğ@"�쀾8^��x��>E�$��`�28v�R	ܼ��O�*!�d��/��A;�ț-.0XK�F؂ �"n���X��`
ay2GS�d,	�ʅ�8`B4�C��9�0?)Cb�;;�B-�a@_�X��fϘd�v�ɵ��	��xB�J.F�h���ݓ_a��c�����O��r4�F���~e˧����U�Qd:FgrRd"Ox��ט�V<�5��&V�X0�"O���f쇕7'�B�ˁ{^@�3b"O��QEf�@�b)�p�Ik1��"O�蘶�.I�Q�iG *��!��"OnĊ���N��@���\�=�v	ٴ"O�������qF�֭W��J"O�U[֮��T�<0B��O�%B�,��"O��A�Y2 �,�2UG�=U��`"Obi�r�9;�8(xv��i\v��a"OJ1`��)uH��;~1"}�"O C�I25��tI�%'3l�"O IA�L�k�$<���ݹj
���b"O��A�'ϼ,Nxp�I\$a_�E��"Ovh9��̷(^�Uq���8 X2�HT"O� f� $� �^p�q/��,HX��"O�l �.�	OfUF�G� ��c�"O
�A�!�1S�X2��u'Ь;�"O�ѧ�Y�w���0�˄Jp���"O,�s�E�.)���X"�L6Lp�"O���!�)8Ą��Y�X� ][G"O���2o�-}�Q$OU1I�p#c"O�K�KY�Ui��¥��|�|買"O�\	�.�P)�\�RaC�]n�% "O��vG�,�����i�����"O���3Eڌ!�p�B� 
 B��U�"O褰�AS�c�H���a�4U��c�"O@,ʗ�\�$�̭Jao���U"O8t����HM>EX�Ś?��DI���8��x1Am�$~���$�RW1O�I� ��X��QBc%�"��Ű "O��␉[�w=⸰�S$B�4��0"O,��Y(j �aB"F��w\�[c"O�1���\��2�F�]<���F"O�h�E��&9\ZP0�%�C5���S"OF�!��ˀt��E�(-̝�"O�tU� *`z �q��C}~ ɇ"O����ԁ,��x�J�;���S"O����R�g�~,#WI��W�@�s�"O�h�"n+"��5����b��IPP��Z����t�L��VL/0�,�82F�	1e�mI���:h��㞢굮��mr�I����?$����4^�X��O��3�Ł��0|b�*2g����TH�0k<�`�bEI���6a�zP�F�F
�0|��lX�'&E1��Q��`���J}"	�,�@0��7�哧g*0)1����]�,�rce��#�^�$ӒSZ���u�"���sӈ��P���D���+c����nZ��t��*�����N(]"��EM~]�Є�G]ƀqdA�E��aGC'�F��ȓU�@E�S�p�{%��A�zȄȓ��e�%@��%��j>�rĄ� �r؉#@`&p1�d��p:����$�V��%2�v9��ˑ W�}��X�ʡ���"j�q�D��B��k�'ў�!����/��0��e�S�?�|ɇ�[y�8B�X0N�U��W8L8V���0vPay�Z�~d6���^�+��-�ȓ�q@3&�.?d��d�R0)�X�ȓ+��L��;v��f�1R\��-8�|1.׌v)^}��Ң,o����� �P��͋.ÜД�߹�����;�X�
ա�<q����$�7���ȓ���!�K�2���QH���ȓR � ��-� �c4��!�����*�J�%IŲ�h
 �����0ziS�H5P�	���+7Ш�� �E��ǰ-���T�+0 P�ȓż��fOP�-��C�HH$Ȇ�2A$�Qg�Z2D,�xd�P�#%`a��T�d�a��!�Z	��\?��ȓ�4]jB��.��|;�DҒ*���ȓWUj�X���/.�5k�Ċ�ф�-j�rq�K=>�����:A�>M�ȓ�X ;��S�NV�sDͲ����ȓ#�ז�8�# 	N-[v��ȓ-f�jCB�y4�4���v����P�<�ɢ����AoN2*PB�I�|lj�V*E�
�֩�B�G��6B�>!�H��+��!K��Q�%7�fB�ɷ�,�xf����xA�ĀXW�VB�ɤL�a�v�I�J8V�$ �2�B�)� F�A��@/IX�0ñ�?8���"O�Drԋ׋0$�K�&)��,s"O�5s7�\�T9�x!�Ϙ�e�� H&"O�$C� 	���2@�4��(�"O�%i��X�#v��`C�0~� �W"O���6�Ĝ)��"Tg�]|�Eh�"O� Z�������	El9��g�@�<qC�I3*1Y�O��v��u����t�<%eC�0�\PF�֖jz�)�+v�<��	k�3A-�	v������TZ�<�䕣n͈�C�ZȸL��FS�<)���"\�r����.3�  $��t�<Y!�B!D�t33���FX �Y�<Y���[V� `�6zuXS�<��䗕4�8�i֥�'"�b(�-SO�<�Sğ�n��̫�	P'@��cd`E�<a�ꀂov��;��*4��#�i�<�@�?�L���㜕�:�����d�<ɄR[I�,س�L�,��q�W�J[�<�SÄ:Ծ��nυI�� �/]o�<IueA�(�A2�-̓_��q�vQS�<�ԭ%"[�|��X�oUn Z��h�<a������EV#i��(QAo�B��hg��C�	�7��(�d�_�C��>
�;���	y��c F9SC䉴&]B�����<��鵢�:\��B�	�x����Õ-yxpq��ɥn��B��#߰�����.�%qVo�5#��B�	�G����jF�;����D6?�~C�I�>��e(�Iͬ$	vE�"j/bC��[�KG������+[5v_�C��&�@��G��æ��cnF%�zC�	�`����a:$�<c�FO��BC�I�EG���3	ɡ����W)	�S�<C�I�e��`0d[,}���ډ.�B䉅�, �D�+<���"�L�u�B䉔gj��X���#Ŋ(
���	wxFC�Ƀ�u�nѾd�j�ۧ뙺#�0C�I�%,���d�Q Wt2�����-�C�	�r�@��`͍{� h��g�@wC�I$p�h�D�Ӹ3��`p@N1TO�B�I�71D��UB��u狦PD~C�	,��B���	5�"eA�U�t��B�ɆJ���B��c_ͨS*�B��B�"���B#O�_i����LP�6�<B�I&`w,Dz�%rotݰ���qi0B�	�9Q�ם^nf-ђn�L&B�	�2�T��2燡"�8��k��[�*B�I�4<I��-e; Y+m� yc�B�I�y�@UIQA�/�7*��]��B�.X���B��<GBj�E���B��9I�H+�/+���
�5�(B�I�VY��N�*1h37�	'B�	$u�:��Ȁ��<@P�~��C���P��+	��`ء��)A�C��	1��JnE)E�"a7�(O�C�	�=6z���A�eo�����9:B�	�+�U;C��#E��@�C�Q�!0B�I:*�UPtf�4C�d�J���^C�2{iP��7g�/(t��%��6ʄB�I�]sr,���+;,LXRE'�|B�	Dh�0��ꍋA2���hT�\B�	�E=���,&(0rxp$!�=Q`B�Ʉb�JX��R^R	 SK�4"��S�? �4$g�=3��-�4l�&|����"O>ᚶ��&��}�7,0���W"O��y3o/q��Y*S���o�~8Y�"O�$����C�֩�4�ǿ�r�Z�"O2)�'�϶9V���׊O�<�W"O�X GF�t�&��fʌ���`�"O�|jw��v�q���Rhg��2u"O�lAd�%[�!��͟��e�R"O��7��\���H3/F��f�B6"OD�`��*lI���-�����"O�%��bǤQ��i$M^�j �Ic"On�Zׁ�J�P\��)]�U�YP"O6��#
,=ڦ��h�r^��w"O���a$�"���b�hѠ�"O�U(2��p��:!M�L^,R�"On���n޼|��̲5F��Qp"O��Ig���VȚh����Y@l�rC"O������=gk4���
!u5�Z�"O��C/��#8����R��$���"ONys�bՌF"R��Ӑ��J4"O�!)�C��t�.�S�*� DXp��u"O��s�_]�,�ɖ�5�z�u"O��@�O�4��q�T%+�v<�E"O�\j�MT-&��( @C<Hj^�Ó"O��B'�c���࡮��JHثV"O@|3d�L����"���3*���"O�|@���"&)�p�
n\ kC"O�5j 
�\Ō�f�X�)UT���"O3�ȟ;>8���m�/>z�,�yrd�s��X�R臤h�z��6����yfJ/<ER�XCg��/7��ti��y���Ɩ���d�$2����ME�y��_�v��X���>�<��Q��+�yBC��h\�'Ȅ���+�ƒ,�y��L�*���f��b� �Y@$0�Py�j�'{�&�b�G�k
����D�M�<ᱩ�>C�lm�՗UL�"B�IJ�<��	Y��(�IN�_��0�BmQB�<	���`h�ݻ�כ��(�a�X�<�qk�A��IRI�-�����^�<��*�=M$��G�)Q��CEjN�<a���t�f�r#����z�H�^�<�� K{�P��[⺐��F�\�<9�dܵ%���v��x^ �"�k�\�<qeO�r�t��ʖ4e6~4!��^�<ɗa�'{�|8��bճ|���g*�Y�<�&�̌:�DhӋ\�\��]���]�<	$�Ǘ5��HC�YB=���W�<�C�)F:��$��B��`�[W�<�R���n��B� =w"٘�D_�<�CQ,~]��XR�ų��qaO�Y�<���Z�@(X" &�d�p�Hq�<I/T�1�tu���bZD�-Vq�<Q�`9քd��A�q���s��6T� �)�HYf�f)�,t�����'D�`�Մ�W;�Q1У��g7B�aW�)D������09��Ĉ�mҥ�3c)D�ph3��5=4(��F�D)`�q�E'D�ت�le����Q%�,���o1D���pȏ�p��C�C���a���3D�X�u��0�Xq�ún�M ��2D�49UR�G���TLW�GgJ�r��.D��y�&ځ�&�H2
л��p��+D��h��I�N�\�����;��Kc+(D�� ��ZS'33���#eT�3�r��s"O��s����V��iF��%"QF��4"O�u�EÊCg�[׃�<HKF�!"O
��td�r7�b4��3���C"O&��O�)��HYL�1u�`��"O��*��30�"1��*AqW�ġ�"O.��WKU'@�f�.Y�ܡ��(��y��A=�j� �#���(�2G�4�y�����lS�L��U�]��y�IdY�栉$n�5�$E��y򀐱 ��(�U�#�ZM�䏟
�y"j�&�|5K"!%�#�4�yoʁ��se%Ĕ|8����E��y2�_<Ju�1�A̖2��ujC�=�y�[�_��@%�Y�xX�S���y�i�*z$�QS&EG�rM3���y�´T��|#Tܧs�ny9����y��zE*EBņ�=�DK��@�y� ��nd�K���+MZ{A�P�y2j����Q�F�̘O�	�7����yH�(&x���?K���	'(��y��1�R̓@�9T�eS��C�yF�	)�
�8b�!{��͂�H��y�,�4����v��^����K��y���g~&�h�T���yud ��y@2I~��Ə�VzdB��yB%�W�M���$�Pa��S��y��)RE��C���,��Y��鋨�yr�P�~��ڶ�^�vd)C
���y	TML�]+�J�˼�Ñ����y"��[��M+��Y)4pv|SQ� ,�y��	�,ZLh�䕆?E��W�L��y��ߚ2��@�1��n.
��&��?�y��J�]}����eOPHG��yb-\?�n��0nO�H��Qve-�y��'K�8�ׅײ�E;6�
��y�Ʉ�a�ۄHӮw�j% ���<�y�A�FV8rP�n@��y��*�yMH� jt���
����B��y�%15	Np[p�֎���;ե���y�T#!����.Z�:Ѐ�`� �y2���O��`	���h�6o�#�y�O�w����S�;v����)�yҬ�$ @  ��]��e\2�
�DcTs�<�4��@ px0ϛ�+>�y���T�<)�U&Q��#�V+j�8 �J�O�<��*2Rt�Fd��"��'��@�<Y��$ia~�C��V#]�B�x$�E�<��d�<� }c�S![ڸu�0��D�<��-ݿ'���"�*����g�I�<��D�~5ѥ,;��@ `��{�<QAH�k�젡Ѫ�Uа��F�x�<ᖅ�/���
R�R���A��\�<�R#W�~B������{�Q@�Ls�<���V��]�	����!��k�<�)ب~$^�ȕ�� � y��h�<!�L��K��"3��(<E�̠��Tl�<�qG�e"�`anD%Qs�i�`	h�<�A	�<ѨՓ���|]�����c�<����p�"����jA/_�<��KO/jԁ�EN�o�.LR�VB�<�.]"7�(�pwH�	k�|��#Wz�<yg��m $$���ɺ;_�����N�<��ī#�4!�/ K���`�e�<��`\���<�Q	�'�r����[�<U��v�ȳ���+�R���b�<�w$,X,B��eg$�����`�<a6�	(*8<��^w���Ob�<�A�uR��bc�={���b�c�^�<��7I�)���R�E��$ip�LO�<�F�0K�D0�Ve���M�s&E�<!	��\|��]ú0y���~�<d��.�u���	neDiK!��x�<��
f&� ���P>k�BT;�.�v�<� @ȳ?3��mɃ/G����w"O^Q@,
��¦�D�5��0�S"O��a�gĲSe����mQ�Μ�"O� 8���<�� ��L݁f�8���"O�Y��� J!"AQ@��$���!�"ODj�D]�*�<9!����� "OXL�2��G��`�%��.���yu"O�5d���I�SaA/u���҄"O�99����3Vh�!A�6P{L\�"O�5�B�<U:�Ej4����<@�v"O8�1�NH��Е�5Ϙ;�x��"Oн����"b��X��M��a�,�'"O�<�B≛n~����Ѽ2Ym�"O|k"�V [��	��ȧnG`�IR"Oj!X�G=ƅEo�Q����f�!�F�$�0s��p�����֭=�!��R�q�<�@�T#���Y`��J�!�Ưa�Z�B4jH.lGr���.�(�!���sy�d��br� ���=�Py��<�J���{#4L���
�yrOϖe/��udȔ\s>��� ��yR��/���D�?j^lZ�ݸ�y�a��y�>tqL�<��4�Һ�y�)��[&h9�#݀7f(�$�߬�yB L�B���C�m�85t��$��&�yf9jX�J���'�Ʊ[gm�/�y/�b25�d��' \���y��%_EB���L��Ip�W��ybe�2�B����f�ADĜ�y��H�`x�ЄZ1U��2����y2��*��������p�ai[!�y��G4ά��y�RE���y�Nϻ�\%1�D���gʟQ<�a��1�J&#�At٪�L"�2��x|��*0��@Nv��&��J�Ѕ�]�=�E	�#y+�򥤟�rzP4�ȓr�ҒOr�| k4��	�T��f0:A�5'·.����i��Y��`3�4��탮d�leRqQ�m��f=��v��	�tz�i���d��$�p�׏�/k��%��-?���ȓ�,T�n�?G8�г%
[&!Q|ԇ��>�a�K�-�j��U��%.��	�ȓ#�X�@�O��~P>dS�f	�B��{�<a:? �t[�s,� �c�v�<�0n��i��|�a(T{��P�&�v�<!P$N$F�f�[�'�w����.�s�<	7�Y
���Qe�CI�!�Sr�<���ى@�A�a �?Bg��Yd��p�<��F�-@!�	Z�(�?��;�"�i�<i�@�<��T�@�N�v	�ELd�<���F���E�,�X2D�\�<1Ў�&><$1�E�+3LP�iU(Z�<�ԃ%!<�R�*�)dqfѱ��U�<	'�Ҕ44������:r��P�<�}޼�b���� .8��3�O�<�AI���}ӡ,7CJt��⢁K�<q@ʂc�pgF�(FXdL��l�J�<���ѤsH���%�� dm�E�<QQj���� ,Y�cf|�U,�C�<��IJ�?����Ǟ&5��V	�A�<i#Ϗ+��Ģ��Z0�y��\@�<)uD�g��z�NB�xzd���[V�<A���@��Ё��D0&����	�R�<� ���N�T�#�aO=�vAw"O����b�&Y1h��@��EmL�"O����(��p�4��e��BĶu�"OD�����`(C�Q�A�,@�'"Ot(� +I,���s�\a8,QV"O��f�K�y��4z��G�l3�ɱt"OZ��M�5���ê��N�8��B"O��zE��/n�R"��;^\��A"O��a�M����(I pY����"O0��� �$7KZK߱�P��"O�M�:!��Q�]L]�"OB��1��IN�(Q�!�f�8��"O����ŚW1�rP��6W�2�"Op�g@y���K�*��"O�S.�,p��1ʘm�"O���@HHtŤI��i�S����c"O(���) >�X��Ņ�9��h�0"On�j�V
X�Ve�`�	w����"O^!!"*��sV ʔd���"OD�:T�Χ3wJd�r�_7?PL�ۀ"O�5�2&	�4k�Uk���(]N��;�"OX���-U(�TI����VU�H["O.�I��Qj��P�ޕBG���7"O�=�І��4�dh�b��#>X�#�"O����^=J�I�w��j0�HkD"O���5Ώ��b�Y%J^44�acT"O~�j�Lߒ8A�0AHә:m��J�"O
u�G'�F���@A_d�&"O��7��O����؅0^��ڂ"O�Iɥ�F� .DJ6��Od� �"O�ѕ��{��Т�ũE/��R�"O��ч�p�9�fL��E�����"OС�H
�I�B�r4J����"O,���7x�A2�j��"m��6"O�$!�&�� ��1 �HL�DNL�sQ"O.��*ËQT��b�ը4/&�"OFL��#K=Z� }X6�O�f.�$�"O�@4�\bȶ�Dn��{�u�P"O�ź2(�j��pM*n�T�j"OԙѠ "Z�P�W�����*ODa�U�
�2�n�r�ꕱj?r�[
�'N�D"ƌĲ(Ĝz6o×cD8�
�'�4�Ia�`�vu;'��$b�H=��'5��A�(�m�n���&U¢�{�'��r�/ަ'pDp��O*��	�'�v�%��=9|�10QA[QX��'}&�ꃏۊm\H;�ؿ�NI��'��I�cɍ5id�b�H]�nnT�����?��T]>�ۢC[�(�,�{��3���#�YJ�<9�iV�c5.���_&H�0�@��B�<��jO5b��`h\$ U*Y2���z�<ׅ	.h����J�k��TB��y�<�g��6���E� "?��[�a[r�<�Ӥ?5ΚA��o�F�@�sbbl�<9�ǥJ��Ă�%Ղr��4�i�<��
ҡ	~LS�)� ��4���c�<i�b̪JZ�st�N<��%a�cN_�<	�-�R�� �8G���bBRQ�<I�	�u`�i����/�|��g^N�<����$Udb��0�ЖG��+6�H�<��I�^ �� �3���A-�E�<Yj�5&��q��Fz
�#�f��xG{���%_A�р��ڝ
q%) m\=uAC�	?S��A�V��9�C��	ʾB�)� :%��.�-!g@?�` 0"Ope�!��!l�dy8�e�%6��P�"OJ@X�d9>;$E1���=BQQx!"OA
�(�8~�-�C��D�l�P�"O�����ho���,V�W?������O����OpL5��-A;�B�%�Εb{��	�'"��&�=Ebh�1�"�=`���
�'-6���`���H�^"mꨈC
�',��LD�#y���qJ�0����'
<h �<^)L$Q�32=�eI�'�&�u��vi���Q�� U*����'q��e�ME��Ia2��#z����'�]3g��O���1m�g�����'�p ��B�F(푶LԮ	���
�'V�d���Uc�-�)l�8p
�'�R���ͩ���Ӷ/����
�'Q�`�C�O�ж�ۊ�J�	�'��u����� �v�}x	�'�4��S,,�D��叕�+�y��'�� $b��W�`� ķn��D�
�'��I�녕~Q��!�Q�BLT{�'T& 8C���l���,	5t
���'�8�ue�8v}EQ�k4� ���'>�K Ր%ج3VfS(xP��'�e�A������ 'i�$R�'���H�!��ܥ �ƙ]%@��'t�0SQG&�zĈ� Q��M*�'��e��!��F
(4�oE\O��3
�'�z`��M[�a#@�#~v�� 	�''B�EE5F��ivM �}��k�'���c��� �T�Uf�v:�@Z�'�1*�
�I}��넅ݥn��MR�'����\FH��F�YD���'|������+m�1:oΛٸl��'n>5 ��U0j:���ÝFt`�'PH��$C�1i�Ƒ`0��������'�B���8�Du� �	�K�z%1	�'	����l�;��p ��!B���`�'vB}�ōØT0�Y�׋�=�2u��'��(A@V3,��"�
�Ah�0�'$e �
���r�K7mBu��'�,�A9]T�E�P���"6�K�',��S�D1^� ��G�^��@x��'T0h���٢l�z0�ģ��dq��'����F��
0�d����
���'���c2�� s�|�a��/L��$B�'c����,Όjs��XD#�P�<��'��P�[�����_E6~I+�'Y��Eޡ`e�	�?%,���'������U"<�ʡ��]7����'��Y��*I���E��*+�A�<�dnݠ0�.�x�F0 ���"�|�<�����񰃡��>v�ip��z�<��h�04��M��	X�}K*@�3%[t��?�çe1����KY6D5�`%�P =yb\��&�����=@�ݸC-;U5����g��(�������s�6wLdهȓ{�V�Y��ш~H�����9Z2 �ȓ1�����HG��D9H�mӹ\���ȓD�m�dHT�v��-#p�ȓ+�rv戗U�L�F��b�,����r�q�L�B����d�I�,�zL�ȓ�� ��Q:Sa�����h$�T�ȓK�ƹAD��X�z�cWm�3Ę��S�? ����a�E������K$��Q�"O���&MOa)�}C�� �:��C�"O�es6��<�J0x���;?�l��"O��`��\�po��@#�s��������O�����b� �a�J�ooR5ѫ^)7�ў���	*S\��S:β����,̒B�I/l�d[Si�~BlxI'^�ZhB�I�&�xH���a �\6wRB��;�j`��&]2p52�fމ	�B�"��TC'C�F�d��f�9����$|�����	�X�F����P$�&�D�7D����
�5N:qiO�7�<I&k6D���g�	�����ͅA���Yn!D�@۶,6]~� �g�ˠ$���iF�>D�l�3�K�x.=P���#�Լ�u�<D��he"�\���i�:���6�,D�]5�0�	 N�@�h+�a��xFn��sj�:yt�[q��.9�	l��� ȁ7*�֐�A��O�Y�2�(��0�ObI��sP13�dR��<��"OĽ��U�2��q��b��3"O���F�so�E�bCɠ{�j���"O�4���ƍ#�L�:5+6�q"O W/�+oj|�3�*^�q2h��"O,<��`ͻjF��	 @�c悥Ґ"Ob��g*�Ӕ�Y�>E��d��P� ��ɂ��3�/��f�}��&2FA�C�	 j�bȚ��H�F�"@�$��%9�"On�0� �%*U<! �N;s��t2"OҬ�������EC�:��2"O�I�t�âku��ҁO� |aXd `Ov��t����ْ�ɘ,��бUI/D�l��G��f Y���IuK�T� �+D������2ps=XtG�?i�LI�!�*D���qᒗ%���CF��� �)D�,��،V+pA�4��1��Iɓ�(D�d�C<��У.��Mb��x�,%D����×�r��WA�	s����"D���"�7���;��3��qГ�+D�p[Q��:�|qّ-�a6���%��9�O�8Ȇ����b(�� Ưi>�y�"O0�q#N̽L��2�T�܎i��"OF�ʵ�ݿqވ8*S'�,0�B(��"O���¤R%���i�Ƃ7O�J��"O�XU�ơ(�@��$	1%�z}��"OB≃�;Vj$y$Ⓚ�4zE�B�0��G2k�v�a���*��,�g�#D�X@�쑚
rN��CdVV,�D�g�#D�H���g*�� �RK�`���.D�4�B�>#��Q.��`4@ D�0��bT!rڑ��@~��D�:D�d�Va�"Kfa��Q�Y���3�J9D��ꅫ�QI���G��\��Q�we7�O��¸ �BAZ}�&e*g��<Z ��Qz�,#ˋ���3�R�j�܇ȓ�l%�t��=;�\
�@6t��ćȓN�1Ir����L��	�aW�ɇ�CpF8�"F�6�l�	�C&'rZ��ȓ�!3A�6�aa����7�TE��
������	2�𐠂�53�0�ȓ!l�]PU%�r�(�2D�SL�ȓi���-�I�����耆ȓu�N����3g��8�H�sᨴ�ȓA��5Q��H�@\8<��	[�ơ��S�? ��j�
@<dSZ���* �c�"OΘ�D
|^tY�H�,�,�j0"O4A#$ă6�� B'D�M����"OJ�󲤈85T��z��0�2���"O<��r�\� �؀ oD�Ȃ��"O���2�ֺQ蘤JE��>7T�y��"O:	c�+B�&'4A�  \� h�"OL���.((�����!Y(œ�"ON��+NV@.4�S([P�[�"O4오��m����eݢ[m9�$"O�����F�̔8�d�����X6"O��A��Ɔ):�-Ag��݈l9g"Of���l�X'r����8]�|"O��%IB+1D2=�!�6 ��K`"O`�y��T#��C�f�IƠp�"O-��,Z�d�.l.L(��X�	!�$I!Rh�tS���:"w�L{���I��O��s��~��$X8�H_''���+0�H��y����C���[�Mуn�6qQ Ѷ�y¦�d����ҏ� ����)҆�y�S� iޠѴ!D��US��^,�y�E�V��p&E-z:�uR�!�	�y��CL��E��@��$B ���Ȗ�yB� �pM8��T.�Ή�D����?q���S��l���0�֡����_���C�]��"C�/����|�����`_��I�ȃ7���X��V�1M���ȓ�����I�[�ݠ���n����*���`ͽK�n�0�MF|��_���R	*4b$%+�X;x�-�?.O�#~�vm��s�!H��1��+�B\y��|��<� ��D��r���v�A�o&D�XhT��]E�IHrcA.	>%�%#D��[D��N�L,�d�/>�Ę�t�!D��� �M&b���P�^rrа���!D�x����,�v�!J�0\^@X��?D�T��[E�4�!��%)�"�K�<��Hy�^�d�O��	*ߠ�22�Q�Q�T u/T5�!�[�������}�A_j�!��U�h��0���D� ��K�;]!�$�*G_v�˗�۷.x�bu�-me!�0}`���C��]���腤)e!�$�1<��B֌i�Y��$~V!��ӲG�xI��Aӕ:D���7$
�T��O�ʓ��|�O�©!-%ͬ� "k�I
���'���Q��ˠDp{�엘?�v�q
�'�|d++I�!��߀?���y	�'	n�X�� ��q� L4�2�:	�'�*�Q%�-vn�(�E99�b�;�'a�qUd q0��W��!a����'��Y�@�f��f	�6f6V�C�r_��F�D΂�"5Х%P�jjL���B��y� ۖ:;4!�S��cXM���޼�y���-+�(���M*f{���&�
.�y��SM>�d��G�R9�U
ܠ�y�m��1t��p��B�l�9�G��y2��>!��Y��Ù/������$D���A�ID�hQjC�w)��5D�T��K_�q��Aץ=�8���4�O��m`���v�QF�j��"
�E� ��`K�u��A#� D���E�\]*̅�6��0` @�+��B�S�d=�ȓTR�[��'/�X�B���p��ȓC>�c��N��H����N%r�ه�S�? h���!��}z�|��cE�K�����"OL��BV� S�a���
pjt��Q�x�W�Qf�fC^�4�a!D�dk�ƻL��x�@C�*��9y1,!D�D�&��*Z=�&��T���S��4D� [�d�S&Y��c6�B��t�3D���h��<�N��с@,)l0��4D�\ ��� V�31¥~�����F0D�X�E:{�d!���z F!��.D���íյq���×�۲�l���-D� �ӡ�m3̡�A�ݒ�4���G*D� r���5"��f�@($T:tk�b3D��8���Z��r)ܤkf 3�;D����ȿ)��$3�N�;[P(�'D�h�)��80��"sF�
&����g'T��ʰ�C9|tIR'Z_j|@W�'
!��P�m{�L����Z���to�5�˟t��I�"��V�גXP�P� u�JC�I��\�q�+U�����- '$C�I1>����o��dn$L���ԟ* C����p�Ws���j,K�&C�	R��H"�
��O��pZ���Jg.B�0`�0��+^j��9����T�=�'�a~�L�$f�[QJ��)�N��H��$,�O��S @��*
�����U�M+��j�"OF�A@�?t�S�eB�o�X�!"O���a �$��Z�gAp�P�"O6<@�"S2f�Uc�%c�4�'"O��D��U=�E2��V&q��@"�'����Pm� �;nV(,`�W��!��V�qx̃Q��~�B�r"ڧ�O�����F�~���1�j}BQ@	1!�.��2g�5r��ĩ'χ0KT!�0S�pI�W�'��P�2�ËKE!�ąW�>h��F�v�*��L�,^'!�� �M���j�8$���w��(Wk!��\>|	�8���;�0С@��O!򤞢<� ͫ⣈�p��CT�V+RB!��RLŬ�XC#�?E��5X5靭e�!��8y�cuł��!��I�!�˳X����hE�x�~�P��W�d�!�$�;���
��Ңa����S,@}!��Б
�ҕ�$�Ƀ8#aaŎ�Zo!�D.z�2(H���6
2�JBE��	n!��ɖn�:����H;L브+cE�KY!�$S��p�P[�':ȍrg$�c�!�$���![�CÇʈ����%)�!��{��	H�-J(ds�d�M:a�!��[3k��!@$瀇xj���P��;>�!��*`��d���Fw�p�o��?�!�d�=�(�-�4MD��'�Ҵ�!�$E�k��'+�'8D6�3�K��!��1`��"/��J0:��I�sE!���FD��fL5�QCÄ�7~=!��[�B��6�R�{'��!C��(!��(c\Z]��nC�g$�q$� !���j��҆h\�&���O�!�D�(�8YG!���4�2	�+OB!�D���q��#A]�@L 榐�&!�dO:΂�pd��U�L��`Ɩ�p�!�(
��@������-�F%�S�!�D\s���c�^*K��M��j�p}!�X���=���>l�"|I�ۮ�!�P^���atOU�5|��ٗbm!�� Z�%]�D�$�Ae��	��H
�"O ���ʐhf�Q�0�3X �z�"O�5���b�L\��L?OVVTkT"O�հ@+G�.����_�w�\I�"O��9F ��Ȯ�0��+�
�s�"O���2��t���bAL6[�^���"O��D�	mD�3��6d��X�"O(X�Ag�3)�"<�Э�+۾�P�"O��Jw���4� �L�vg�C7"O����`�ͺU+�
ۜ �^P�"O��r \�r $��.j�N�P"O ��#�L,|��B ��T�3"O�h�'���f��䛙���3"O�x۞�����;Β�)ɦw!�D�cXp\hBN8�� �(�=�!�d�(|���Dfƻy�`y�D�t�!�&%�)H � �&��IP0�$�!�$��(�^	�6� �*�$#H�p�!�d�	.��aԧ5r ��Ţ+p!��rY���	2b��Q�o���!�d���L��c��m����[�Vj!��4$b`�S�K]�t�B"h!�$V=t���hEe�u�b[1O	�V7!��m+�̙Pwo�BŊh8	�o!����e���:�ٴԷt!� ��@ A7e�����+U!�d��lh2�F�;�b{���56E!�d'~�x�W3?���0q�	�U!�-�h%q�LӶ:}p�R�f��3$!�$�%`�,���?ǔH2�V:!�ЫV<*SH�4'��Y.a2���	�'����AN>Ә�e��i����'(��� ψF;�ah5� �n����'H,H8t蝍z�<���G(:%(Q�'���yUρ�\+:4k�C[�8I��C	�'� Q��H�,b��@�2D7�6��'�V�xAÚ�["��d��Rrq
�'���@w�^�^pܤ�4+K�
v��	�'x���' �D� M`g�I���(��'<�1��8}���S�"�+C���'����ۖ(��@R���)[0f�y�'#n�Qb�CO���ѕ��5>� ��'>��5$Ӌ,x��Q�=QΡ8�'}.�%kո	�"X�3��-u^���'�61a�*�O��a�5�7q���'r��P�@�(�Rd�[�f~E��'���u���Xc�6,J,���'�����'	.X M��	�v���'&��i�QC��Q�@��j��'�PԓWa�1l�j,����2uHT�'r@)5D�A�<��>���
�'h�Ds�"׭
��EJ�g��5�l8�
�'SZ�`dJ?b�jsf�-"h�
�'g0}�%�k~�t�R��o�
h�	�'l)��eB��HeG٤��H�'�HǣW� ��1��;$pY��'��]C����eܶI�6&�=g���
�'8��P!�O&LI*Ȩ�`�dj���yR���T���B�4�D�p�Ш�yb�'j��L�! �9&����H
�y2��7ąR֨��5[V�Z#�y�)��?����a��"2Ț�����yb �QM\�{�l�`� ���߱�y��K�Gj捉p	�
Y����fվ�y
� ����e5m�m�RB��v\����"O�d����Mw ��`Oy%@Qh�"Obph�^2v&|`/\0n~Q��"O��b"-��t��#X,dk.er@"O���߬7�p��!Z=hb��2"O���&��?r�(�g}]$�	�"O���6�?jt�4�:A�"O�\S��@�u&$�j�;6���"O�d��oO$v��)棎~銀�5"O0�H���4fXl�Z!�#]*�u0g"O
��O	l>�$��j�tD��"O8��w��uL��9������l�"Ox�F �%c�Qe$��J����5"O,U;c*ĶE�0I�S��#5.��g"Oa��k��3�^E���4l(�8�"O��m���p�/�&7x���"O"��F��O~Lyf�0�H� �"O���f���|?�	I���*�a�"OL��w���_����,@�S؀�i�"O���a��H��M �ˮ�Hi��"O̥s�C��7q
���L���"O�8ss�O48���HR�&�x��"O� �IPr��Y�D�
*h��S"O���+Q�^���P�Qm^)+"O�AAwES�!���P˼wW��r�"O�*���`�<�ҩ�+hZbu"O>(2��%R
v�XfoӖ=f�i��"O���рȣw���@�.�9dڽP�"O�m�PB4p|Ԕk�\�"4:��"Of��G�0�� K@0M�Y��"O����-�0�ZL�96"O`Ĉ�g���\\R0�T�Q7�)x"O ����E*%:���$��� @��R"O|m!e��Q�� ��� F *��"O�}�#ٴgb7n��`.&��"�%D���G @�$;���'L,e�� �*#D�`#���!o~f�0�gHo�Ĉ$�+D� Sp���
�dŤ()H2�N'D�LqmI� @����k�ր�ë$D��	�0-��x���Q��Y�&� D��p��J�cz�`���ډg��쳰�>D����O{d��`�$�(5� �g7D�����T` y��ϳ1n�+�*O��qP�'��T!��$-�X�(�"O�r��Fht�#%N�s�v6�?D��	&�M�{h^��`�/s�XQ�>D�H@��h:`؋@���!UF�� D� ��AR�"���R�l�-�@���+D���ǦP)���}6DLâ�'D�D!���ce !�.�#K� �E$1D���T��!x*��s��Ă<C*���!D����J�	W�v�� ��7k7b�x��>D�4����[��C�BrO^� �7D���FE$G��e;�.�4$-�X�7D�,cR2Y�`���L�L�)"�3D�P"�ˉ2y�MX6�HFȔBSb3D���J��m�Pԫ��5F���K'D��3���" �"��\
ؑ����/!�$S�)�Y`�	�[��x$!_!��U����t��/_>u[@E(�!�
>���:U��Uv�˲oO0(!�ރ"i<��Z�KD
��RH\��!�D��Z�c�b"5/X���a� 2�!�dF2(��m����E~p�S�s!�� ؅IrOB�Q�j��3o@�; J��T"O�h���
q�����B=_��Y5"O8IB��^o�L��0�T���*�"Ojy��NI9X�H�̋4�
X3"O X�Wjܔ2�P�
*54��"O|l9��w�x1�^~b9;&"OY{�K�7A輁�jO�#{��a"OR��2I�
^��9)d鉙7����"O�0�V#X>�p=PaiWX5Ӥ"O���#�
,������4^�̃"O�TYP I$4+,A�r�N�l�:X��"O��t�X�x�l��PNO6\�"��$"Of�C�<Jy	3���T�q"OR�:BO݋#H�*��2a��	�"O2�CԂ$�J]Õ�Kp����"O84p"jR�D�ي& �(R]X"O�LCT�\�u��aEY�%b��"O�xP���3Bf�gM���]2u"Ob� ��[
G4%�:N��v"O&�S��:k�<ıc���LG�A)�"O���$����p'MC�v\b�"O���S�M&z�j�b%��R5^�
"O\���9��85'K�3 �p�"OJ���#Ĳa����f؍8�X��"O�y V���[q�� ����2�$��"O�(s���1|y��ʟ%k�~�`�"OH�S�Å9�0AR0��	��q��"O������9Z����dI��Iw�=��"O�!��̠<�E�F	�k��`"O��fg�BcNE{�H+8bv�I2"OB��%�1TC��s�]~��#�"O6L [��i�&@1i`�� �"O����# @��p�D�����!��7���P?7�Bl�̑{�!�d�G/���¨A+8hp%�{I!��gil�3����+b�Q�:9!�$@,'�cO�F�lE
��2�!������D��Y����Ɩ>�!�$D�4(�!���V�?��c�Kޢ �!�F/q�� � -
x��� �!��ȸ:��t���_�y ���L�y�!�DK_ǬX�-@'I��sKD%�!���'��4S���AH,��ͽ�!򄑔<� ��E��D��#R�� �!�d�9}.��u$�0P�b� 6|���&�b�уў��섊�y��d�d�s�T�:��ْ!i\"�y�ˑ,�J2��҆��-[A�@�yB.�6o��I`��.�tii@���y⥉��P�o�
[�$C�˓��y2,�5C��\�d�̤1 9���Ȫ�yb��ԾL��S�}&�9I�F��y�ₕD��0ڠ��l�ֽ�"*���y��0bD���0�� KrmI��y�aH�E��"C�[+Ǯ`1���y"��<- r�h�MC D��!�V&�y��р!���am�:0#�uaaJ��y���q�*}�ƢZ1x%vb ��6�y�	�=6HfcV��o2�A�'�y�E�~%�����~+�J�o٪�ye���*3AS&t�l��P���y�����B�<��T�pf��y���`(h����/��E)�yR%�A@4��_�U�ZYr�D>�y
� th8�Ի}���)G,^  F"O�{V,ڎ4��]JE���D��"OLi���8�B�P=?�P�"OV�`�Y�d��3��T$��Ust"O6Q`j�!�@�9�H��O�KЧ�y�CM�b�@����<Nd��Bg�-�y2E�h�6Lh�o_Iv��vjR��y"��98Gj�[�o��E�Eb���y"�� n���";�䝠k�yBWR��3w�]$P�
��yBfH� ��rA-Æ^	�����I��y�`��m��@ⓤ����n�w�<��:��9��_
+8�8�$)N�<aG��V�!fk�ݚ�Q1��M�<�"���{&Y�_�d	�����PT�<��M�0?_�!�������W�<YqN�#f�s�g3�,ui��}�<a�F76=Ƙ(�j�L�@�I'�Ho�<!�!ďgn� �L',ܽ�f�Am�<��߶�(�S��"@���Ph�<�р�D����.S�U��<�"��~�<�blI�u%R�s��G�#I��@	Dq�<�� �7DJ��Wl�%o�:-괃GH�<����$O�$)!�6?[��i��A{�<��dNh!*���۲�\���a�y�<�@]��L�)R��z���"x�<�a(�0=�0�{S�2 ,��r�<B��:�HUŁ�)�b�l�<�V�������D'y����uH��yEz; ���
��yF���y���Ib^]P���`{ �_�yRƼ^�D����	���A@bƂ�y�	�b�@��˪��*ݐ�y"��F�.�3���{�����I��y�)_�P}R���,��x��,
D���y27;gp��D�t���sI��y��\�P�r�J4e4AU��yBȉ�y��B�hp>!"�j>bƱy����y���.N i��!j�Rt`BE��y2�!2tx��B.qG�]��bއ�y"��x���c�*ʡdc8�CQI>�y�!W�w�ġS�F;d�z-����y�釿*���T�l��^ �y��Q;2�\ ��	�R485$U6�y⢇�k�<�y��9)�r�8�)F	�y̏�]�����i<J�J�Hr�B �y�n�8;� ���ՊC<@�e�y��	����#��-�h�C�O��y�]�y��e0�B�{ѧF��y��4��5��`u���"��y�͍";o���R�S����0�yeQ(�}��h��Y������$�y��ӊ+Y h��φQ�6����+�y�X����e�N�^�r��ݎ�yr�^� ���P���ءb2E�=�y/\�; B=����a�*�h��Hj�<!#"ٓ
��"��5�px��B�<�i�J�F����&\����(�@�<�eφ�p~D�����[�y �|�<�!�G;IΩ�e�+2kn�a7� }�<��/�����3�@�v��R�Xw�<ёAX�erN�1rQ�E�p�h���r�<�5@�t��s��A�~͈��l�<��oҧD� Q` �d�xy���g�<�  ��6��1'�əo�S(�P�"OaX��ޑ@��H6m��B 1�E"O��YņZ�)�l�p�(����"O�-��0t�mE�s��4)�"Oġr�Y rC��;4�ͿuCD%ې"O
�q����A�\9F�B9J y�"OD�[�[�f깲b!BU:ei�"O��%ߖ7�V	�� ��$7D	Ƞ"O%i��ߗ���S�n�P�"OH���,
3`"�0I��Y�V��#v"Oā����[g�5��l@�Q��LA"O�!�L�?f�0�R�F=��5"O��x��K����2 �'���a�"O��[5 �n�|	R�!�K���9�"Ox8*��ɼh7���ekɦO�&��"OZ���|�6̓6�|$�i"O����FE�<5����uoD�&"O@e�r�$|4�2#O �,ek"OT�IG% :������EbdӴ"O:���S�NRU(��ݟ}U�$9"O�%ȁ��"�h���]�z�a'"O��sF�;`��D`CV����"O�m�&�U�t�9�Q*!���"O6� ����a*ed���J�"O&q$��8tF1笂����ط"O]���	�V�>d�TK�9u�Ԣ"OԈ�.�n���V�/�R\� "OP��ĩӑ7�0-�`�)0s(EK"O�}sn
�w�K����F^Ԑ�"O,$�!V���E�y�FTr�"O����Z�B�Q�P�ٸ=��D��"Oh̫��X?i��C5���~2,�"O8h��� ��Y��D�"B�+�"Oh�S�ۓk{�mX�F&�P��"O^���/+Fz������HyV"O�B�B� 1�\$;x��� "O:�"T�fo�D�fcʙj>��*�"OС��ގ ��kB�L��-��"O~��Qo,l*�-
� �2Au���"OĬ���WG�X��#\X�`BA"O��'��vk�Cc�8�إѕ"O��4��>jX|H�r-C)m���S�"O�}����<�ʁ�˃.R~�3�"O�p��ޔEJDxZ�i��H�#s"O|����ǷLC�A�3��T ����"O�`�bޢ2k�܊���/ �p,�&"OnM�2G\�W6ntc@�A�_=��y�"OBI�儫�mq�G�.#.��AC"OV��l��c�f��FH/J�2�"O2u����K1��;G�آ58�l"O����{eb��"�+h/�u��"O1(�,��03��%r(4��"OP@���CE�8�/�;.�ـ"OD��M�I>(�'�)h����"O�\���#u�ш�戍}ml���"O�$�p쁻.�Ԙ�Tfћ>���Ӷ"O��r��4-- �+��#(v�1x�"O�|���D1*�+�KQ�lt~}�"OL��tdQ�T���#_�O���g"O*E0*�'Kz�]�a�g��"O��3��ļ.�B��vo�*�	'"O$Yc�
�e��j�J���"O�
i�/��<: �CK
,jG"O��8�K�p̈T��/T-]0P�'"O� ��R�d#�|�"���K��:�"O�P)��B�Uˈ��
��Z�r`�"OvЫ�j�S"�bV��6��-#�"O̛��� }Bl��fLL.n����"O���B�;p�<=2e�W�"2���"O���ơ\).�<�u�ʢX>RL;�"O�TpC)��(-B��
3( ����"O��	�NIq����e.a��"Of9��/�T E)�}�P��e"O�a��Z�^�>	��AҾk]J��'"O��KQ�%q�7��P���d"O�``E����3r�÷K(��"O�僧e��f�!�3��)g.i˒"O�����W�E[*�-^��%"O��C�Q���j�)Ǐj"5� "O��b��=iH,�E��h���"O���v��K������&K�U�$"O�db���$A̕c2�: H��["O��i�ǜ�P�*xs�,IB�*Ob��+�3�̴��S�(Q�p�'�Hyt�	Z�:	9�㕑j.��:	�'�p���&�<Mf	�qrBEQ�'Ǯ�s%ޒ&���b��Ҩf�Z���'����>4������+d`� �'���3Gꀺ^����˫{m$I�ȓht�9�w�]�V��m`�	�f�D���~��PYӠ�+��m25��
��\�ȓI�P �V*'e�pc���>N����Ɲ#$M5�(�q*;/�F���+nq1'�"�t��&�X:0`q��
�h9$�ӂ����g��d;����Lr�}A$��#+m�9�� �M�n	�ȓO(����To��!���_�8���?��Z-L"���x ��cЂ\�ȓ�\��h�3ON��G�(8�ڈ��a�JYC�k� ���SbW&q?d��ȓq=LI*�)�(��z�jڢHK�l��!-8Q��Q3ܩ�0f�39�m�� w^�k *�&hY�UA��+,�B͇ȓ �D���B =急�"��2=�(�ȓh�nr&돕>�\Y��L�pYj�ȓ|���*6Đ"=�)Y�B�k��e�ȓ)�U9`�C�q��,����D�h���XalY�$b��.��s�RwR6��ȓw@v�R�퉞�vӔ�J�7v��f�f�S@	�6�~9
CAX�WP��ȓfl���@#M0^���Q��W3��a��h��qlJNY��9'�C�x+t����T��7�BL�`���,��Q�ȓ*nH�eD@��R�#�
�U�Jt�ȓw�.��B����H �G�+\XV��0<��{sF��s��)I{��5��zilxX��N/P0y1힉b.JȄ�o��@Ā�-�
���k�-L̘ɅȓJᬍ��C�xPx�ad"P-e�ц�'�"����tU*i��+s���ȓr�I1��V�B~mQ�&R)czȓ$q4`��ϫ ،�ǯ�!�r ��b����NT�)"�}Yk�E �$��:��ٳQ*��I�ܸ���ז?�T���`�lC�P���$��$�.7`���W�M�M ��<1��5_Ҳ��ȓHo�0	�H��J �d`�ċ� J<��Qp��)0F�.B5rah�!%uR�Q��S�? ��xv��hz�R�bW��A"O�D�C'�3Xnt�"!b�d8�K�"ON�1�cY�O�J�ʃA��j�(525"O��"�	�	o�B������fǟ��y��C�4�R	"�ϪX�Fxa�S��y�+ܚ �N,0�0}�tظ ʟ�y⊗!@� ۔!M�p�V�PՊ��yb�Mr��x��f�n�9�g�>�y����Xh���%W��P�!B��y�#�B��d��cHe�: .���yB�]�z��	w`�v�x(����4"���S���G�9�,�k#��=r����h2�yR�ݧR\���
n�~��!���y2BؘI� �q@$	�c�F��dɭ�y�E 6�����LD1���Apd��yRI��>]����+
K�H�@�8�yr���7��iwe�Vh�U@'���y�����pd� �����d#�yҭ�M�~!�	���MJ����yB�,7f���U#��
a�N��yB�� (��Xp��͞�ƀ<�ybi	W������_i�����yR&�D9Ĝ
p��3�|=�4�p=�}�WP$q{�@Xm`]��gȑ�y�P�q�$�$@��O^�h�b˛�ڈO���A�7b���+2c�)\�blQ�� l�<90͢U!�-����#"Qt	�p*�|}��'�45�!�Q�6��ӫ��j- �'J�c��.�TX۲*��V$���')��p�c����!���(�<���d;O>$0Q�]j�� �[2&��s"O��p3�Z#���vL�j���&"Ox�8e�1rx���ul p����"O�(䁊�8�RH`�*�O\.er�"O&�8G$Qm�𠐩ũpД�b"O��PAB�6�X�6�ĵ#B�(S�>�;Șy����@r����քbT]���<�;�jђZj�A��P=m��|r�0��"� u� q���M�a1�=�>�דPN���\S!
�b1��(OG�h�ȓ^μ�؁ϝ�"ix\���#WbM�ȓ w�ȃ6�)eR��j��̖. �t��c��
a��6���R�K�@Z�5�'~�$$|Oj���:w��$*Ɯ@=���4"O�k��B�T0�1�Z/Թ9�"O�y��B�*,�p�ҕa�)�0�"O����$ݽC�:Y9�Q
�n"r�	M�O�m��&̡1�z�:w��"�Fip�'���Âl޻!7xq�v��-�]�<yU�ڞ�)k�2M�8yذ��_�<1b僸?5�qZ��I�8��07J�Y�<�2,���$kz8�k���U����W �y뇏��[��P����z�Fz��O$�}��P!2�����^�T���"��eX���O����X�$�����̌	�B�jd"O�	qDƲWZ�م�U1{�J���Q��Dz"�Ӌ8�`VE
l`��1jF����'�h��dޕw"0�{�T @������?�hO���Ч_�&�h��Y�9M�48DI���yB�G+KD%rsiB�}R!yT��ɨO�"mB�~۰E�`. �rZ] �Y[�<����H� |�E#A�@��J��<���ٷ���ÓT����P��}�<�ciHFB��`��)�l �˔U�<� 2�(�!��Ae)�*�@dQ�"O�!�ыS�'�LC�7��i�"O��@�O���2h�nХ"�"O�hs��B-R��`�M�f$��"OVq$E=M@���T�4aHa)�;O~�=E�ܣX{�e!b.�]DvX�*���y�!Q�=r��R���6;���$E��y�m�\���fRq� ���jÃ�y��U(*V�*& I2~�:eH�N�6�yrGDY��zF��EUH0���%�y��Ɗ|��1f�|����k���y�e�76��Ly���c	6�B����y�P/����͆k.~�(S����y�Z�f9�%���b�>)s`����!�$Y>2�,(B�E�@�
��FD�)3�!�d�,��a�
�}��	���%O!�&!��\��֎>�XYP�g�!�D(Td�*�B�"I�h�g��y�!�DJ�]=P�jE
Z�ػ֠OO�!��X�;�8I�f��0HYcT�]"C;!����&�����疥 �tr��f&!�$ӴS��\J$�l�l�nv�!�$@=^�ڝ��E�?�0� g�S5�!��p
B*J����#i>M�!��^�B�Z��A�H^�&|` �"O����/G�t�H|`�GK��X�ʇ"O��b4��6�x dG�4�Xu��"O�$���1)Ep�C� �5��hp�"O:��Q���h{@��eM����"O�9�EE91�ٚQ�ĜD�1#�"OZ���#=��������`�:�"Ov�rӇ�0r����F(�p���"O�)��"�=t$A�R����HF"Oli�& �*5���h��9���)T"Ol)��-�&Y���ڐ�B�E)�H�'"OB����C&M��0kF�� {
~TH$"Op|�c@#t5�B��͌4�N�a�"O�M����P���cIM/A�؄q�"O"q��G�(B�X�V�&m� %q"O��RL'=�Pr"-�Q��T�&"O����<$p%cqi�M��-`�"OX�ZS�3�(��E��N��Aq�"O��n�i" q4%Z#���"Oh����=q�f�#�d����+�*O@�KW�R�},��P�8�I9	�'�.�ɕ�'���  3qBP�b�'ܐ* �N�u
=P'�C�t��1��'�D!�%eW�Y�nP d��=�&xa�'s�\�7�����x�痺�i��'̀�)����D� 6�� tjԙ�';*M1��L�k�� Ye�~F�m�'*�U�Y�Q�m�t`
�z��X��'��)����8g�x ��k��1��'�j���Ϝ	M�E��Ȣ$d:ْ�'ND}�ph� ��P��΁��ƅ��'�p�	�M'140��!�	��a�
�'��):���O*D�R�E��|���	�':x���!�6b�N�p$}�����'a�@����b�����Ilz��{�'q�����zu2��'+�4_��r	�'t��9�ɀ�d[����@H)]߮03�'�e
����u���`�*G!2R���'��1R�!I��Ya kB6��q
�'�T���!m*=�G(���`
��� ��q	�6 0�T�r��+Jl��"O"1�C��:Z���B�dΆFj�*�*O�u��	@{Qi��}�z�
�'�H�+1�Q=Ѩ�xA�ͤ?�"̡
�'�"�͇�-}j�Ɲ�fΩ�	�'p�ȃ�N��H��ĝ��:�	�'Yf9K��c�B�a�*#��*�'A���&%�0���[��9�
�'��c2�+&��2(΅&�� 
�'��ʀLW�y�z,�qal�0���'�h�	gkA�@�&��0L	6322p��'�#'�	<`�����/o�8��'���	���Gd�-0��,��}��'@pغU��$�
!Y6���M	��!�'��xЂ��3<\@�H<|XjU��'�]�Bl�s�tq٧v*�ɫ�'����υ�֥��iNa����'K�	A�
�!��ŁS(�2[�0��'����GO�	*I������No�ի�'��`�_ z��єaH�H�D[�'X>D�2�$0�xKaCu��k�'�a�u��;5�{��k˜=��'����Rj��#&�	0�_��r�'�ZG�V�I߾��g "W�X�
�'�򄳡Ȓ�}�A�҅�Z/H��
�'���Z�IM7�\q���W�����'�T���ME��:a�_	V�8��	�'�z|R�Γ)+�B�cF)6�	�'	\�[����]4Й�s#�Z���'��Y�2J̠�	惛<��'Q`��`���5yޑz�cC�tO"�J�'�JLP��ζZTx ��͉@� ���'�^@��� ��aIr69��,	ħgu.%p
�N�ԑ�C�]�^l͸@l>����ȓU-���o�(i%������!r��ȓ|�jm�CH!*��k­I
9@��ȓ2\�=�F��}R��K&��[k��tR���K�mZ�9AD��L����ȓ��4�V͒�Uu\�P��a	~4�ȓ_�ƹIB�Q�_6���Sɋ;CŰ�ȓ#(�"�k?O��Ljd,�0P�8 �ȓ/���O� y�R�J�E�|�|��ȓ;.& ��T�8�X��+2bZ\���l���4o���B��ƍ�� <��n�:1ȑ'�4)d0�5L�D�(h�ȓ[|	� l ?�6�i��R�X ���ƕ�A���F�q9�I��p�d��ȓRY�tRtJ�e�>$!�c��,ܴ��ȓT�ʂ�
	�~�PR��htb���?],�+�ˠ)]��X�Β��0�ȓ^%� ǥ�1�^�p��	U�^���b#p�&�$/Ѡd�� ��l9�ȓX���h��D<� ���Xў}��x 4��iŽV�BhP���yц�� �����EaL�!)Y�9�ƌ��"��,#��[9Rm%�է-NP���;�h�8∗�{�Ή�dM��;�T!��56�4�pNТQ�Cc&^
�|a��j��o��>�耱-W�*�.���|�R]�tn�|�n���&�1�"��m�"]ر�8GN,��G"����X��m�Ð6�PSA��4��ȓi�hՙ��ܟy���ٯ{��ȓ!zM�F�^-|�#ǢW&4<=��S�? �ݺp-^�]xy�����8���v"O��XG�R���eW�V����"O�)��`ز�50e�F�Ƭ��C"O:��EAV	-��͟2g�T�ɠ"O��3�Z2�|-(�[�����"O>42��L�g����ū�44�n0�F"O6ZF��J\��1J��sEl�b"O۶ _�|j���( :��[�"O�ղ��77%N�b�胟Z3R��e"O���I!Gw��:���e-L�{�"O��աH�7C�4��v"O��T"F�1 N���
ɻ2�.�Z4"O� ��Z3Tt��K6�K�g(�S"O��+vk�8Z��"�.{Z�9u*O��W�W���CЀM�����'�z\�@���i^��bR9n�'�$�K�a�x�u���Y��-�
�'���a�VtAv@ Dy

�'�6�ҶCO�,)Ĕ �J�M�4��'��|��	����\�Tb��E�(���' 1E�(3ɶ`��F[�A��'ֲ��3��]����B 	��1��'^�7�S<h��`��j�s�'�4�e�<P������c��B�'Q ����{,
�LaÈA��'ҹ� C@dh�0rl�VY`YH�12�	T�6�)�1|Q�E/?2��D!)	I�Z��
�'�hy+iUl�D�S�eO=��Y1�'��h��^�.y~��I�x����#Ƙ����C�%��s�h�>�w�?9c��$�?]WF%y���	�R^F�a�	Al�.tɔGG��x2c��$���V��rb~��(���?1a��l�A0����d��!��mZ=��O'T̒E����jb0i���ߑz!�V�|��#�l�eɶ�ۇGET`%����?A˼�Y�4z��$R��?�+�Kg;��O���-�..?��b7(X�e�5ZD2�O�$�@,�����Ff�3.�yłٲKgʤq��D&p0N4aa�T+�����d�@h�'��0�YR�֌�bE�0fp��Љ�$�> ��g�ba"J֛^��#F,O�08��w�5�v��pOذ\čCh�: ���IOb��񨒬k�)��
�Ay��5m�.�&��A��,�|�;ħ� ^�v̊A�Ӯo�=��*�~��w{h 0�J9"Њ-�L2���'7�P�'G�(w5�dC�[�^��ӣa�=��h�$��3������8N�È�eJ�$3+O,�B��Q�����OV�R���'~��bt�@�6�u�%�Z>5EL��c��k��m�#�,"j�k3d�8�x���ݕK3��
��V|�'�4���g�&k�~8b�aɫd	P��}�JY�|��D��������(]�!��0� W�He��o��\sn�z���K�h�I'-��[��͇�I!�����N7s�$)�Dɗ�()��8�(ȓ.��L[.�O�vu�"�K�'��$����q�"-�'U��1*R�j�%܊�4V�qr��D}&�U��>�a�	�[�� &P��q�cE��U�%�	e1�a-܅9Q>�]�q^rpi� �GJhHgQ�0 �hJ�#T$L�CV�8Bu�k����к@GqO�1=EQBh�.)��#�
�px�E½��%���0r�����3W2�Q�_2���	@��\�rJJ�J@êČz*D�e8�H�ƕ��X���S�mUXa�H iP����8�(mQ�/�Ȱ�V��[S�,�V����d9��7QoJ�g���4��Q[�$T,j�TAx���&h��1a��71AT��ViZF}�F�ޑ0��qcӄT�k�V�'Y��n���9 C@ˣ;���� �� 3���BC���gQ>}2��
�u.fR�Ŗ�n�6� G��&Q�8J��#T|	��(Rv���݆*�ܡإ@]F�5�O�-:��D�IJ�V��$��,"�1ON0��@�0��)��]
��Ņu�ք��%��yY����54B�)"�T�iT��K�'�+��q��#�L��d�C���:b��5�X��$;�Eh��`�	�Jq:�H���8_K���ϐ��FIN�!
�3rIr�2����U"T�x�+��#�!�_Q�dhT�ص8~�Tk� 	-A���)eA��@�i�S�I7E��
�k��P�lxD��4�w�IQ �[9]�ha�O~�ҭpa4D����R���iT��y�t��a x�*x	EH�C"���{,��2
_@Zf�0�I�~EVy;
[�(����-�*x����Ҟ<ֶ���:A�����בh�H˳�%�:�"��W�+�|	ᡦ*�O��a�^�N�f�sD��Y�Z}	r�䕫-D�t�SF��A�$�AfH��g�? hʤ����	��t�ڱ��"ON(Dc��zS,p$$~��"���@1J���SC%�U�w��0,S�>�	�*������G�j|s��ϫ~B䉳1|����);zu�K6$K(<���_)(����)T�pc��s�'��VE�L�Q'`��(~�����`���P��Ka�%M��C��:��Ő�b�F�P��93��"�M� �lL���J�\���Gy�ɸ80��9bn��nH�|�2��c��ɋ���s��Y(-B�<1���\M�=f�k9z�G͙_0�D��'�+�e�(��)�y�c� @bi��O.;�ap�'���Q4�Q���!�'	��8�t�O��K�oR�paz򯃏g}7Dиq5B͸N� �y�kA��$刕(��M�.NFX:�'E����H�$��� ��&��X*�'
̼h ��p�R�f��1�ݫ�'4���T�%7������'�Pq����;��X��L��Z�'L�O��<	���sB�-	S$hH	�'�Q��LA
l�n̲ЪT�8��'WP	t�(0���
����8Q�	�'m��"2��:_��l�D/��r��0	�'�$�B��@��zdi�?\����'����G�>�Q��W�B�5�'�����L������8d��'c^�1�k"�H�5'�:�R�'.�j�OOR+��Ζs:0�ʓbw6���i��C�=��BӸz�D�ȓsd��;&MF�c6P]�r�ͳX��q�ȓt�
Ux��-�ȱa�.�4:�rx��OV@i��VD��H`o��9�*�ȓ[o���S/E�X�鈁"K�a�}�ȓBx2M��ϫ'
%���/�Ɇȓg��x����$�W�c�v�j�'�:��&�ŴR�:|ГKڔR�lI��'}X���./3�h��k-B
���'M��6!�7&��%I�> $�:�'0������Zqi�7��Wp����'�4�3��<��!����AǆX�'w��� 
�
�R��03��0��'�(d����HQ\P�)�-��'�pHqE�]P��)f�P=#ڼ��'�2ْC���	Vڍh��ێf�K�'�����35�FYɇ�U�(�T���'"��扳HJ���	�*N6m8�'��Ʌ�^�r=Ĭ�A��2P|�5�	�'1|�Z@��Nтъ `[�\a� ��'�$�3�(|*E��E�+[�r�'1��Y�&���駨�#a���'��0@��($�(A�3�X&!����'�
�uױ4լ�+4�ɒ
.
p��'�x�#�%$�j�U�0��0�'D�����CFX�G�^.� �''�<9�/U
`;th�wOQ��ѹ
�'�ah��w ��f�{���z
�'M8@S
Ծ)���|چ�i	�'�p5
��ڔZ�ϭ~\P0�'6F4��O��ji�I�$�1h�����'�xԋ��Xg��%r��ܑ>���'l����9-�N@�󠅴�H���'+�Jա8N���#�/��В
�'�ʁ`����z�
�k�;�ހ��'Azy���abԹ��ӯ>=��2�'��Q0!�I�X�Ѱd��4U��'e��^��}�&�ʕe������ ��;���7���J�In���"O���«�^�؃�@�&qa�"Ot���Sl���a�F��5��Q��"O═p	^�t�(p1��$O۠,Yc"O�	w��1	4z������:�0"Odq+rd](�	��%:�(P9"O&��Ǩ�+�N�0��8��Բ�y�B�{2 	W@L*��$�ц�ybn��\���B�>F������<�y�K*~x(r菢O�ɑ@썊�yRS�Y�%Z�+��R�ܻ�M
��y"���Ρz��:Q�l����y��"�.J&�X%R�����ä�yr��f��J�/��&��Л��yR�<I��y��I�e���@�H�y�̐\>Z��l�Q�H\``L0�y��K�-��ī �ГS�PH����y�cD�J�͹a
_g�iс�S�y�T�����hD�\8 �z��I��y���2�\�r#J�,|L\��O��y�ü\b�QS�C�v���Sp\��yb�Q�x:�����y�2i8gNƦ�yR��2X`T{�dz�	��ω�y�# b0-I�(io���$Y�y���?o��Lj���	>԰ȫ����yBfߚi��*���3�>%D�P:�y�	�6jx��#N�%CU��y�n��%ը` ��_���y#ج�y"l�q���a��+hB�ړ꛺�y�Ó$]��X��M�g�P����ȶ�yR��-(A�8�`H\S�=h��"�y2���:]��GAX'�i��Ņ�y�F"!A������&1��0HB�y2ȕ�c�4����W�,sg
X��yBF]`�L� $�H??Jm3��گ�y��ލ|���9L�� �C3�N�y"a�8A�nM�&j|T8�-P��y���B޴�r�E){��3�m���yR�ޙ]æ�:�eI� 7�Y�[��y2BG�r��0h���&Z��0�Aӝ�y��J��(#��2�R����y�(\ ��q B�T�'�-A��*�yRf2J���b�8"49�+�@�<��֩W���)6�<]�D��P���<�� U�������D�j(� B_�<q���BK�\+��9<�����F_�<�q`�VC����l����9s�]U�<�S�P�����1j㒑B�dL^�<A��� Ԍ��_�~`´��X�<'⟄eZ����h�Z�`�A�s�<�'���Xr$"C�9Q��A��^n�<I&�ճo8��)�J�/0��g�s�<����m�X�(�!7�`�P�i�h�<��"��T-��D,_�V����BF�h�<!@쀲oJ2)x�eԤ'�N�"vnCe�<iES�\P��Ê
�����u�<飬��S���б. ppȣ�%�^�<I2�+z�p��J�ԑ{��W�<1g���h�ȭ��ދL��i���K�<I���<�Xfʀz���A&�O�<�a�V#VG<�K�G��:@���@�<2��c ����@��I ��EG�<���V|����D��� G��2 �y�<�6͐"|^Ly�D�:���S�̒t�<� �Ź�@��
G���E ,͡�"O*� *����Z��ȕRT���"Ol-�T-_%y[��rP��C�$+�"O�}���]�M�@����s�<5��"O���Vm��aQ�3@��0�"O2I�U"ݫ{
NP�f���V�T���"OZ @�8,��9���O#KaP-�0"O�("���?o1�m��K��{ʹ1�6"O�MX���t��)ITI���.��"O����m
O�n�JS�[8~�~���"O��:���Fr����"��O�ε�"O.�8�%�<cI��Su���^�FИ"OF�Sd�S�1�����w=��K�"O�!A�F˸"�����6 �a�"O� �t�"V�������1����"Ol0*���2_����u%V�,4�s"OԌ��G��z�����2���bq"O�����V��� �D� ^_��"T"O��RC��9wd�Q�cӼ|�f�Z�"O�y���+z\p`"��~�h�r"OM�P�2���a��&�W"O�|0��-=i���ߍm0�A"O����͌-�>ٹ ��s[&�q7"O���$tq�tj�
Wx���"O�pHiV�s�Jd)�I�7o��Q�"Oz}vh��3�a��O�,z�9�1"O&�z��s�ġz&�;*f��Y�"O<��K��i�N8�pL�&]�� "O
��s��%%�U�0� 627i3�"O�P_$�`:@��Z	B�"O����d
�NxQCr�ޘaJM��"O"�&�S?r��u:�Y=u���X�"Ox�p�[+jUJ0M�9K�<}�"O�	R�	O8]��8 �*����"OR����g(����(� �Sc"O<��H�@[��V��e�Ƅ�"O�PY_x�� �C��46w �(U"O��(Ԏ')��F�Dxj��"O|�!�]�Q��F`��Vm&�S�"O@MBcI��p�.�W� 8o��"O1+���9d[� +ǩ�
9��K�"O��s��/,˜5�0h�;sZ�C5"O8̠��f�-� ��n[�݉�"Oޭh�M��g�Fh:E�	�����"O��T�_�;����	�^Ɗ�(�"O��7J��0�[7�F_��Z�"O.Z"k ��%�(O
>~���"O��H�nO	1/�3b&C�pTle��"O���e�F:�p�p�_O`���"O�vo��|]C�B[�L\$5��"O�a�%�O�4궀I�jHZ���"Oƽ{T�Y9?�Vuk�O�@t�"�"O<t� G�fA�u��{���#"O^Y���]ᮍS��C"�H�iU"OP�y�!P�ck��I'IZe�lJ�"O�y�M� �r�#T�@B�05�v"ON���H��u�7ALa�(Y��"Oj�#�E�]zf��"`YsҶ��"O���ͧc�2E2��Lͨ��"O\x�e��%]��(!a�N�6	i�"O�pgdD�A{�5�E�Gn�(M��"ON���f%M���n��V��DÑ"O���'��f� 
��X�hT!��]"D��_U�1�"�!'H!�� ��r%�YZ��� �TTc�"O�pU���r�|�tE� ����"O�\�%ÌI��)���ͣm�fA��"Oԩ)b�E�j�*�$�-d|49C"O"d;�ǄS�e�¬��`oh�"O\0ʠE�_�v�iQJ�EP�@�B"O8�kq��j�|P1�W9l�>4��"O�8FEޏ��34��3j��� �"O �TET�a�HXJ�dI�Y�Ԝ""O�j�]C��z�#���M��"Ohha`�������s�)`&"O�ar�e�I[f�C�!E6��h��"Oh��J��y��jX�w�&�St"Orp{u�!�X�bp� ��x9B"OB8*�#=&��҇�(���*6"O��:3��ub�1�,͓~ڬ���"Ofl�4�×"瀉kaLA�O)�i�"O��cc��:/:Js�BC�p��!"O����R�E���S2|�Pb"O����,ū"g*�JwŅu!��Җ"O��+��ӯ�\ʣE�("��
P"O@��s�C).(���F
.8F!�'"O�5���W�p��ǐ��1��"OT�Uk��Y7�E��C� uI3"Oh��qLV�}��T�2'D�v�J�(@"OX��ѿt�4��e�	c��� �"O��hM4y�&p�E�0�lmC�"ON�ƭ^-<&>�wG�L�ʀ�"O���vN��U#Fu�B%_!T-,�4"O\�J��'MERx�veR�/j	:�"O����� d�-�%Ś�k��XA"O@��4E��xt"�kڝ1�d��"O�9桂"L�a��:���x5"O0�)� ��h~u���	�b�X5u"O,Q!ÁK��Jb���u�,t�"O��@��v�A���ρH�0۴"OY�#��d >d[s#��z3j���"O �����"�p�Ď�P��`"O�!�ū_?8*D�bOs��Y"Ojxkgo����E3׊�F��}BP"O��0׉T�m��U��H�s,]Ӆ"O�a:��U�|����j4���"OFx[��� �52+�	SeF�J�"O\@!`�7�bhs�J��5^��*"Oֈ�#�¦/J���	T*1
%[W"O��5�� ђ�(��K�x^@s7"O�j�!	<D�E��m�~!��"O�����^�1��64��b"Oj��sU�~6%��Y7RY��"O�] 7�7.-��b��ئ�t���"O��2��Y�oм���)ꮀ3R"OF�	 ,L�N�0�#����@-{t"O��:�J7��F$48��z�"OXe�)6�tm�AC_;L���"O���G�u� jt�&r�n�*�"O����aػ\�"H4 b�P
�K�o�<��`0L�x@�QFU7A�R�i�`�<��o�Hp�S'�V���˓�i�<�Ch�mψE��g/U�n�$d�<	bJ	�-D@���o��ns8���'�f�<Yt�Ҟe]�p��@!? ek���d�<�' �I@�DZt��!tRZ�2ց�O�<A�I���MP1�a�M2�-�H�<�"��s(���㊚.&YJ�
�I�<� ���AP:���l��-�`D`�"O��A�۠Th��f%�$p(�{!"O��%��!~0,��꒲*xt%�A"O�SQ�C�J�C��Uv5�E"ON�I팂h �1�wA؁v��P""O�h����8|�9w*�;(ɖ��"O,��_� h[��1���s"O�Ԋ��;^&�)&j
[c
�"O��y�a�,z����a*�^�>#!"OܠT+J�z�h��qlN�~��(��"O�Њ�Ꜫvn�L�ТB z#Y�"O�|��i2X�A�aF|X��"O� �l�9�,�1�?Z�Rd�$"O��R�f/6��$kۖa� )Ѡ"O���&���Xѐ�U2!���:W"Oة�#GاG��h"�|���ق"O��)�ޥ ���B���c�Ba�"OdXاό�$�ā�	��*�ԩ�p"O��5-�9�|E(�ƚ
YJ� �c"OB��3T\
 ��$K,h5���%"O����&�9��9��#�9C"8dq�"O2I���Is��s̴P"OԨ鲃������"���x$"O��r��;, H��c�DU�ă"OK�a*Zq�#/n���� ]��y�i�n/�DZ�S7'ڑY��Y �y��:k����k�3ޠH f�P��y2F�f��;	G��H�O���yR�э!�D1�qnQH���P�*��yB�Q(7*`5����=RI��O��y�Ńh��,2�ٞ0��E�`×�yro�5D�&�Ht�ɂ3�n�;��Z��yr��8"��;���,����0A�,�y�e�8zn�P+��$�vQ����yBQ����+��+h4a��!�y���"�$��0-�2 ;����/�y2.�����U�L�Nd8���-�yb�U4pZ�h�e�,2�.06�X#�y��݀`�$% tK���@I�����y��Z'���a"��e1�4CUi,�y�
�p�,!����`��\A��M���p���0?�6H(�(9�
*oҎ�[FX�<٦N�7�B�ՈO,7@�:���[�<)��.D����ǝ[���ɷ��p�<I+�Rv��q�J�
q�3T�^�O���a�L�T�1Oq����b�7E����n+Y�hUS�x2׃[:U�b��|����c�F�
S��3pHrhx0$ʟ41N�-0T�b��~��*W!(r�kAl�'=q���c�{�p�W>�?�W����Y�wj��"���}�j2�'�UpG��)L��ǩV�CzyX�ޟ|"}�D
P�"�t�c���$a_�a
pd�2I��!�mG;�H�Z& FT)�ᓡ}�. Z�ǝY2\q��^�<2���"e~ލ؀��'����3C*��|)�a̞� ��/ߛٲ���n�r��Q.бJ���+����~rK|R" ni�1iŇ1��:���'�- ��Đ��#��s��nځ'�hQ��B���Sf�[�p�BC+�%[c�n}P��4&�����P� -��2�J|"d�+&�v�yp��0W:�P0��K�;a�v(�?�~�u�ؔb�^4���T�T���u�n�<9�.�b�x�(��O*�AvkE�<!�� C(�8��N��� R���<���s@b໗��5+��q�sn�w�<	�,�Y�m�d.X�%�0'��|�<�7׻!}���"���)06n�{�'�ayҥ�&L��qB�".�<�`�F�yR��#v`i��O�����&U��y
� "���o��/xc�O����p"O��2�[�t*��0���"ª�� "O�D2�	;Q
թd���dИ4"O$�/�
�̑��/ζ1�v� �"O|q�g#]0_[�:�]��)"O��!�(F"W���k�Z4��Aw"O0đfI+ؖE�L��-���	�';ܸyb��~m8!g $
�Z0�
�'�d�rp'�=	e4�Q%ƺ5�f=�	�'����ԃ� �pd]0x��	�'��ȪT/�<�D�G'�&E*dy�'M ��!=�.9j@
AVt` �'�P(���=z���,[�;��Y��':�"���2�&߃�f���'�j��A�RX"`��� i��h��'O\ &BY���cv��_ٖ�j�'Ӧ��Ă�F�
�{�+�6']8��'�0�c�gە:���1b/�Hl*�',�C���8�.e3�Q�n��\�
�'���`�  |*���I�gC����'��x+�+n´s�ūe�Ly��'����D4
�$9ҭ�d^����'%�(�)E�fg%h��*R(03�'��q�Q ����12���U��x	�'tl�)e��r\�IZ�焒<�X��'�R���I�=����Td��&XZ]��'��
֣H1���#.�q� �8�'!��
G		�p�2��V,�?p�BU#�'���E��'<�ZR�/˚k���
�'�is�
:$�آl�v�(u�'JDC*۞(��ic�G�=K��I�'R�%���Β)�K��F).F���'�ܝ�r΋�Mb��̅�TRL��'SD .�+_�u��ʘ"���s�'����΅od: \%��� �'mZY��τ�}Ku�ׁVJ��TZ	�'7"��c㓕gK�`�%��1����'#6esW��+�)�(9 j���'����e� �
9�#�A=eRܨ�'*�e�tˀ�
�|سm���s�'�`<Z��8���hАY�l�X�'l4��Fd[��X��cD��>	����'>&�(�eN+G�*܋$��2u��B�'?$��UF�$\�����"̖1��'�BYز������Oθ_����'\&�0��,<��+�(̇c�h���'v��D���I��R�Ckx +�'����bΑ�_���R��<��]��'pl�����K�h9�2�����'A��PEB]:>\�1l��,V��Q�'�ι�Bƾy1�諁E�(��l8�'Ed�2 ���hJ��+1A��!�L��'v.�B���>(>J��&¦���"Oxp���ʦA�IbKA]����"Ot��C�A�1�<�I���u���"O�xђ&�+k�%a&i�g�B��&"O�a3��7���I�!F���;t"OI�ĉ�*�jl9t��:��l "Oځ�B,٦�A���n$>%c�"O܁�%��qn��5I<7��"O�TY&Ꜻ4��d���˂F��y�e"O�xxv���6ێ�k2k�=*��E�#"O��Hv�K6�>\��N�c�,p�"O����P�z~�A5���M��dj�"O� 4�"��[�i�4�&�. l�"OP8hDd�?�9�O�5_��`�"O�Da��8Ը�C��Hw��#"O�I�N@�t����kȐo��y3�"O�E�����H|��*ڠ � �"OV���
��s�,ATI�g�`�S�"O���S�%��h�gѤ{Z>00�"O��y��o�����>@EXk�"O�E�s"]�([��ɡ� "qc*O��s_ W�����"؍����'�0%8���` �H�܋6�i��'a���Eg�4I4z��&�>�a��'y�h�a _DsB-*�_ 0)T�A�'�ν���f�p��*�"3��[�'^F���ɻg�Y�	�(JvH��
�'S�iJV�S�gs���wE;-��	�'^U���k�Ʃf��,���'�V�RD�7>tHh��N%2����'�J���Hh����e�[>��QY�'�yRu�J�U|0ar(�g~�*�'T��B ��7gw���NS���x�	�'��QK �˜��}P��)B���'v�PYgb%R�����P��ZQ+�'>z���-�'Q(�� ���)�$M�'B�3'W�:1�������$@u��'4�Tk`ᒾ;�VD��͑���'iHB�J&&\ִ�qŉ;Zp���'��\	1�J�7.�iP�۷@5|���'�d-k�c�J�|���Ꮑ$�j�	�'@ 1p@Y#Z�tE*2)07�H�'DD��"L3k��c\)�\�#�'2P���L�Y����P�k�H\�'�\\��Haq�pR����O��)1�'�Ra�FK5V�@��U*S&TX4�Z�'C:LB�a�6��8��Ҙth�{
�'�0,2�b[^h���#J9f��@��'V@0��^�w�UIr��>_��x�'8��u
��ʝQ�X;%~P-a�'`F�K�..-<� �JR����'K�!����i%�ɐ��
G \��']�E�M F�)agNs��H�'�&�!b	5��u�.	,.�=h	�'��f�P`R �+��׈��P�'t�غ'4x45��_�t�(��'�*\�qM\7Z.�$���_H@�X�'��bF��t��#��4p�  �'�(�!��yΈ�C3g:1��
�'P�hQ�ES#�$����a�S
�'|����΅�H��c��X��B
�'���x��#3�� K��-S�Xc	�'(4usD��i�hLJr�ʩP���1	�'����$ O�\/�R��K�~�0	�'%ح�uFYY��0��`��q�1	�'�,�C�7ѢX�Ѡ��y� ��'� ��)�#V�<,jBJ���P�'���"�^��N$�� ]� Dy�'�)��&�tuAL�T�"�P�'J�ȉdEؑ4�Zp���Y�PX�(r
�'�ie-���0�I"�D�' ~���a)y�AAR��<Y�t��'b��$��0!f��
�1��P��'��%X'îD�2�b 
<��C�'��m��?0�.Y�4�P1$���'�<�{�U���%E#�p���� ة�)+�hHh�hZR�,���"Ox [��;:���n��#����"Ȏi�	�4rz4�4 P6G�DA'"O��6��>iܙkV/̙{��=�c"O���Ǐ��9I�eYc�]1*����"Oj����_!:������O�8�b�B%"O]�V�04Y�fs�8�h�"O�%!Re��9=x|����B�L��"O��CD͝Mm,*EHn��C�"O��Q�'Y-F�r�#�v��aT"O&�Q�H�'?dJ�Ȑb 0R�A�T"O�l�d�4��S��&T�4hA�"OP=!��̱a�b���/ܒ|���H"O�4�����V�ǉ"w��A"O@���G^�X�ˬ-QT%�S"O�m�	�=��`����?D;r�Q�"O<Y�KQ��sd�a
&a>D�$����%ݚ ʠ@�[��U���<D�HS��
+�؁bÌ�#"\Q*PK0D�ЉC,�5aBP�#K�Q���"��1D��`1Ĝ�;XIJw.Ԣ\�:y���/D�("uAM�rD�JR3b{
qQ�1D�TX��Ю ^E3C��/:M�3��1D��b��/���e+��E��yC�0D�0:��eh���C�W$p��Z��!D�8Ƀ�ȇL�ΈD�V4|����W�,D�0H� q��J��
H���q�&D� A0�d�q�a���:r*&D�q��-?Vձ���?1JX|b2�)D�k�Ê�1^��r�W
F�R�	D�%D���2���p�q�wb�q�bm��1D���v��r)�yp�X�^��ƃ4D���EbP.����l�=FԬ	�=D�L+��/*�ۖ ��`��ɘ�):D��NǦV�Rԃ���7�p=� l8D����Q���P !����1D�4��͝18$�a��):�����-D��"���/b�y�q�KD�ΐz��+D�<��E�u��i�T�Ţ;�I�,D�py�K=Y�� ��ĕ|�l�Sn D�����|�0BO	,ۨ�� )D�|���	tOʌ˷� 1-�`�Xѩ<D��r.��t,����fB��b��s�<D��1������@:��@k��:D�����$:�$�0L�7nd�6�:D�P����,v|^�3u��r+,�K 9D�@��o�)q�����W��4�"�d!D���!mɂ	����'%
$0q� D�4��ݡ`�V	�`�Ӝ}�8%�!D� �2�	�d|Tإ�*��n?D��0�(�1keT,Ҳ`B�>a+=D�����$&���Z�Ϛ@"��H;D��KK9T�Yp�H��pr�!��i;D�����>k?ܘ�˃j��A'/D�$*FD����x5fBNd)�g-D��ZL-����u@U^LV����/D��3�+4u���@cK�j��� �a#D��� ԱS�Fe�GΉG��hp`#D� qc�j���p�J��Ĥ��!D�ԃ!"�R"|��I,윤!��;D�"�O�>5�\�C�H�n�j�9�D?D�TJ�k�T���Z��D�T$�l�J?D� iP
G�+KޭZ��Fk�䨈d=D�2g�ZQ����I27 ���`�<D�� 8�t↵=��4�]=D#��Ї"OpMZg�K3?�<� ߖU8�$�"O�����AQ"�$�Y�|��͘V"O���F(d�f`b"��eZth*�"O2��e@
�VJ��u��0*�Xu"O� �Ï��|�m�v��4ta�"O�L�%	   �*ot��R�Tږ���'�n��-��Y!a9>�T!�G��6U�@�Is�t�b%
 e}��xk�j45.�y7lW!_� �'
6T���}��neV���q�vPp����'�pDHFM�2���ֆU��*�	wLg>�YS���k��X	��7f�����C b�p�	��&n]#V�Ϩx4��D��K��� � R�-� ��K�'�-ꄎ�7 2=�B�o�ԠY��,��'��M�R�h#��-1`X���Ҹ�|�B�36I�à� � 0��*j��`�JP�lWj���7�����e�庆e�:Ҵ9�ъ/a��pJѮi]x��S`̙6��'c氐���վ��!-"ِM��$\O@�/�tE�����m1`�;8�6�S�e�*<�����5���3.B�_�Y��N�-�|3@+��{r��40閁�V���g��AlY���'r�� �����i�LTu��
����T	�+˪����V�r� �#���N�@��aLۍZT~� wM"\OhMK��8�XR0 ��$\ikb��5jz�c ���?�"���H([A$J#hDFł��i��4۷��-���A Zk�Շ�C�I[D�1�i�1�n��	�ɴDV��� �6�E�J[J�UcT�~���vC"�i���T:W�D=;�z}�'.��"�/��M�g�a�$�e����ޤxg(�7Wp�ч@\�\�pKM�v�bEW��c?O-�ߙ2~��ë���h�Of�:V�ы*�%�4��?|�*ѹU��ac���nY�HER��ۓ'q]�0�S	R���s�X�\����		Q���/��_���i�i�0���)�\�p��><����',*��W�ܶ����m��Y�$��y�-M�\�0��"¨{��>���k�d8�pNN�|j�`$D�<�EE� ��a��R�>���Qb��[W�@��1}���E���$A(	;�hA��4� Pq҆ſ6�!� ':��*��	U>�8 2��A��CʭL����;��HCևF�6�*d�%[<C�I�-?�(�CH�+��
C��Br�B��)5TT<B��̋V�Z�a�+֗v��B䉐{&xM���J(Z�>���;0�B�1O��AP.��4��Ԁ�;.�\B�I�ҁ��խ_ 9�p.�#N
hB䉟��Q�e�]�R�����FŞB�ɐ"���sP��+��}�Q'�$.%XB�I>y]�A��"�9uW����޴`�VB�1hՀ��d�� ��Q��<@!B��&����*��v$����!�j��C䉺^f�Q0�	��φ��6_�C䉅�H�3P'�t`R�M�l��C䉰']������#��(: ��4i��B�u�q��P�2���
�̰B�	:,���O����r5`��r�B�ɂ6������X�8�����e��B�I
m�2��p��)A���4e�5)�4C䉞%7�R@H7p��tˢ�ʛo�<C��=�f�H��т3t� �����C䉭H|���Z#D(I��֡*�C�ɴi`pYy��U�(r�Jվ`DC�;�(�Dϑ� [N0s�V>9C䉍,p��K��H�T0�Ei��<1�B�8����� �:lB/�C�I7
=Jq�Ƌ)98�es���7BC�	;k�0Tw�5s�9P�fB�g�^C�ə����qb؄q�j-c��=hRC�2l��`ҕO^������:�tC�	;��@{
�	�-�ţ\1\ZC�	�P ����*)ät��A�x� C�[rX)���4 [�0"H��/zB�	�`�n�����Wܸ!�"�,"��C�	:Xdi1u�G�h{���F���:��C�)� ����S.n�dH�G�,Vh�s�"Oa��E=� �q���=OX+$"O�ي#dG�AC�tѐ&�7���Ȅ"Or�x����W-�س&��I�$��F"O܉�P#
�8n��!�Z�!�洲"Ox�����.a#��9㌇^^�09�"Of�`�Sڌ�(��,'iz��f"O��VO�8d�����M�}U,��Q"O����������-JiK���"O�����Y>S����	��0Ry3"O�487)�[ �r4o�;��8`"O�aЮ�.#D53���x7�'�ڦE ;P
�]���a j.W1�A�� ���;减�Q�qO�>1���^���7����j1�E$���� +y�c?���*Ս��t�P
ro�8��'�<��i��UGα�Ì>,OPH�Wd��tܐ(�q�ڮF}ƥH�D4~G �`���3c��b�4��b?1��E�%-��ↄ)QA(U�U7,�����*2(mL����QVx���f@5lJ���+j�*Q�Cŗ:k hI��;i�n��F�%<Pv���� 6lF���'�,�ͧ���/�@���*��?%b��	 "��	Zq.myD�x6 �2���Q�)y(ؓ���b|�ىuJί3�r���
H؄8�'px�D���l�౉.Ӈ%���pʌ�{�ƴ�OP8�A��.�A�R>3;�A����s�O*�R��gFR�Ņ��/�Eb��'���S$�<^V���X%G*џHB6�Ew�b���-�0!
`�a�A�&`�T�9�KW�=�`,3����%�b>	�@�!�x��DU`z��g���8j��
��7�daE�|\�=)�$�Wav��S�X�p���2_Є��SJ�
=��A��<������?����s�X�Z�p�#)Z��*X�?�(�
ݥ(Ty4�E:��tDv�X��!F�XL���>���$�����#�7:���B�b�8^�NQ@A `���f�vղ%��B�A�	m����\�?�O���	��"�~4�,y�,l9�.]b� �(�'n�R��e##?�1��/K�Α8����4G�L2�fx��3��K>w�3�!�kN�	C�Y$s��o�7`�0d��m��g�2�d.A�l#JF?����q�s�6ʌ�i����#H3�.P�%Mr���̈́l����c	2�<x��]>�cr˛�u���%Z�"�(�
۽���y5�`�t(K�[�Ψ��a*�S�n*^�~�4x8\�����4i�z�zQ+�_o��E	2���C8v���o�,1�bT��Em����[��B�hǇ-�L��֠A<r����[D�@:�i�ym��E�ٙT�\	�e�H%P�`�wN2[���A�O(��D B�6{�����+@��r$H8E�b�u�۲{`��
@6��6-�a�]���[zD	�f⑑r��(��7d��8��G�h.9i�Q�FIz ��C��xr��)w�Fbƨa�O�̳�eL;�TZ��M�':�}�qO�<8_̜��iģ0a�&8`��ed��O8�X9%�NI�tr#8_B^����LP5�T�T��&$0v�����
N8�L��Op�H��F9]ADt�AD����"C9-�e�3AE;H��AQ,*4�Ò��:N`��!D���b"�/�Y��9��K�+�������M�W��$�]�7�詢0��+	ڜ���L'��+S+_�����y��-^66���ɛX�&�+.O"\���O�]��"�@��]k+�t�����|/��q��^��ft,@Z�3��,�|e�r�91.��s���Afj�jn�)��;ӂ;?��@ܭV(37������*��8����W�ŧ��e��f��J����Y~ITp*@h^me��� �:����'�ĥ��m�fFZ!J���kXcq ��#	D0�W n!@�+�>i2=�D��w\?5R��D{ ȱ�"E?aw4���#t��U3�4,~�qBD=L�B2'�۷6bju�R'�-N��tiĢu��m{3�'t�q���I�R��Am2Dj���*g�Q$O�
���'���"D���6(: Ǆ�� !K-O��nâ t�����P�>���c�]�u���t�2���S�]<��	�l@���I_�i�^�����C�s�浹ơ��U�A�	3p�(a��n�$� !&;�{��u���hu\��F�&�ʍϻz���K��H2`�]�"I�e��o�t� 0�L�HT,EС�'������P2 ��`�"�P�{q ؼ�~bh� �p��\������K�*��yP2(c$Ѕp�_�;��H�@Q��b��Ђ`�ɉ��'2D.�#�
 ��k֕jdh�"^gr���H��(~6�ҠE�!!�A!F���:����r'B/	RfAIR�U�	/P`MQbb��Dٱ��M��Ph�d1R�lOr���&H d�V�r�C�*?�^��@aVj�0`Ɗ�/%3@�
��ćPr�к��P�7���^�$�ZXXu�M�:�1OX\HU�,��'�TT������;!�(����D�6:����N?1,�R�(
K�ZH�q#����s�R)�����w0�u�fAϕ'Ժœ�/����'���jD�.&P�p�も7�lH��!ЫG?*����2*$pS�|�Z�#R�#
F�8p�5�d\ᇁ��,���M9s)\��
W�N���c1,OP,��k,<�� #	��GW���ϋ�_JH�����Xrm�VF˜|����ę�Z͓�@w���G��.q�$�"´Y��\�|Q`��O/����~W@�wON�O8�12l۵8R����A6{�� ʔA�4+���EEQ3(`8U� �gsdA��
*ܰ?�T��/��dy��ֿU�B$��c˩N� �ʂ늖}�_D�?�'aǭ�8x�.��v#�.z#:M9�'���Zv�V<2�kV� 0pːh1i��f�b��sc��g�L	���z&6?6yݕ����`D�Σ+�6���.H�K���뉯L�t�"�R0$f�����hx��%�7n��P6bBl��V�׈;RDq��9O$��1�z��K��g�? �@���:��y���φfD�̳���H�x����Z�w���Ba�ȂD�WmA�?a:��G��N��$mQ,	Yf��ϊ&2�t@ !J��L�˓�h���O�aXqÕ�Xv
i�7����X����0PU�gP��p�s�+�e�}ҝw���S�!��LRc��o�h�4@v�pBR$�JlQ���!<Oh r�ay�"�@�<�PW���Y �C^'M���$�P��0���T<�e�$N�?J���G�:�;��Z�����EH^�9�-Г�{���Î:i��)q�ըof Y�ۀ!E��7B�b��y��&ѷU��-X�d�!z'�E�Z
e�.Ԡi�8Q�h��%�֡�E�Pm���4�@ru��	�J�S4 ?��?S�-�)R�g��У�Զo*r�so��<�	�	�Ӟ�H�;��_�j�X���j_�~B���l�=5���̓|��m�����B�í���߼�"t��RC�I[��M���[��ʪG���r�d�7 a��� �ɹլ�
$K�/QD�]s�&�����k��K�h	���pNW:p���ף�b�Z�����`��G
�5�1&�	�c�^����i�t��E��
4�@m���N#I��A��.ZM&�(�L'��(-��V�d��UDC1�^]�!	�I��I�i�&4Aw�S�`c���4D��P̊�	�S�YS6M`��L�+��6��k�RAH���Bʩi�e]�x���h&KR�9A,-i�=w]ة��o�a�0�����w���[_w���#梘.Mj�$� �&y��Q1N��p|F�@��T�����Ś���a����T��a�Î�iI��B�ݝJ �+��T�p6�H�f�^/u�ݩPH�:mnB���~�f�Ч�ȃ� Æ&(0�����};�(����idT�J�!��}��q�t}�k_[���¨A<�D���ז.��m��	:'��YDc
��dY��4�0}I�а �fH�ЏQ�/Ws��\�$ |cH�hĺ��"��16��Yb@C%	0�����H~�@�Hj8y'�ؕRt �&�3�d��=7�P� g]-7����ÞM���c��ŏr���RS�_<4�?3�F�p�۟�ؐ�Oͥ>����\�K)B�U�z��� �T�"P"�+w�օ�t���Xڑ#Ʌ)%v�n97������}:-F�@����Ō�+LȈ��S"Z`�l �R��	���R��si��2W6-۩[��r$ͫ�E�
�V�Z���#D?D,ѣH�!3��X3��++B(jD�E�:��$Z�iJ6T�P�����A6Z���� 2�����gI�|mb����Q3[P��Øp��7�*h
��%�O2��@G�yfz��f�0?����=�ӥ�3�$� �F�J$�B�\�8_0�AHS	wc�X�T�C �)����&� �&	K>�� �0=V�����{w����8�LȂb9Oz��G�� K����I��hON�E���Q���__69�-��Du�u�QAy��	"W� �HP\/�vL�#��?����@�>�	W�F�9X�ݳ7Ȝ�m���Пs�0�#Ҩ�:�V,��o� ��O.x0$�ٔ�<�Y�_�~I�'��DؐQ�Pm��BW��i�K�ą\?pBIk��_0:H~�#��v�q,�����؜'���3i��u�k��jܓrD �!�\�r��l#��8;wh�S�����x�K7g�����vC��'r��tsv*;9vd�o��"��a�50*:�˕�[�y��T��(�RTL+�S>]���䑢<�yvD%y���)�0�\�a�Y�a@.�!��K�r%�KA�y
&�"pШtI2�x��D%dJ@�*�A=]�Nu��+̷D�(-��'���z��
�Ym���i�" �~��0�@
9�TQ��0I��x�f�y�������D�d��7o�=�����<�|!�ıH�)\{����ƭZ�!��J�N�F�*q��'�@��i��%��A,Y�9��J�K�R�Xq��
�t�ڻR_Z0&��.;�* ��nX?t���3�ŀ`�6�S˂��0=e�GN8�6%�]%����-U.�M� $D"kT����"�#gl�"%��EL<�;$ur� 2h��]�B�xG��E�PXK/҈T�ij¨�V�X�Rm�5%� ��Q��'��Ec��O�RP["��U�hD�ŻK�/o���c�h1V�u$]�j��)?2��9�pa�TC�ѓV��m���#sH_�F�C��i4>�)�$�?Z�ؐ�B�ZcF�:w�CJt��͹!/�c����k�8#*�E�e�T�u;"�Q���1D��xB	$E4vi��h֬4�l�	%"��h�� a�X(�6mʳB��prR?�I�jU�B�ED�L�ؙ���`2Lz#EO~�a4@b%ϾZP���j�:WDh�@6��5W��{���@Q��4�/FGb��D�F
YhUT�B� �R�ֈHAf�����5AU��;�Bo��B�X�
Iy�Ι�w]�(��Z���|S�@1r���s�eK|�� ��4c$	wY�sU��gNZ:���X���B��FIz���D�d�RŨ���%]�H��|�H `f*T�~7�x�ug�&EAj<�7��'�@|����	(<9���!p'�̠�섖+���`B�Rf� z�"���t�uRR
MC�F��a˙�*X
�&	L)�F��HG�~��sՉ�d��>�R�������3ғlㆡ�DH��IzJ���
A\BM8Ej%z�%�s�E="�� D�W�<Xr��0=|N��"K�G^�?����
�	�b�K�Gx�ȑB���{�j����<@����򮐜 z����._| �{��R�k����4��	�%F�=-w,]�Q/(u,t{ ��_l4��ҥb�����?�
s	��>�4�@sA��h�����M@�;X�!�2���~b�o������"Xf�� ��[Y�ՀV -�x	ⅆ�
kIS�I� �J�ꡨ@'k�YT�M7b��r̔��P��A��CO�@{�Ȯ&�T����%��k �G%�`�~!21'	P2��� }^��c�V q��Pe8n
��ge�:b�jJY+.(t�����v�#� װ>���Dg�.�qC�-_�W j9��9K~V%ɂ�\w�'	�}S�M_2U��d��X@��VEl��}(��i��s1˃Qٺ����4	̂%q���%A�~U��2`Jހ^�:�pQ;Ѣ"#�����V��㟰`�*�<3v���B�&ANPQg�O��p�c�G�<��Q� KZ/1D�:'#F8"�X���K�����d�(u:~�KB	��9��7�׶:Tv�P5FrC>��g� >k#K)%�l�����o��q0b�04�Ήj��^�ٶlN�(.8+��+�?�5n�i��4YP��	6�X��M#gb��"�O?���� b�{��Q0?3�YQv�^�]ϐX8���(Qf
%�cU�I�b!\	I$�VI��/(h V��gBV�m�fc����	�\�R�,�+:��(����+�a&P�y �
DY�����n�PXH����D� 4%؟'@��E���'�@����P5�`��ѕvL���N��tL�P6�N6S3Ui�D ��$K�@��`.�\{��rA�����J�X���P2Q	�% ����<�J�SSb؅�|U�<Ys��n}R�n3$=�3�U�7&�U��h�$$�|5y���(T��2(0���֐P!lС��D�L<�R��d`~)A��G�y�89S��D3*0���Q"��8�JK�@���zc�%}ȥJV��7���i��1[�h�����f5��(�ꋚD�����J'yƹz�̏2�� (��Q!�6Rָ�႗{'�x�B� As��M
~(p�Wb�.2�D6PԼ��"�D�b��ǡ�O� 2�������FxFi���Oܕ�'�`��g�T'I�4c��z����AZ�o�4�bb��#��-ه�-I���_^I��d�'�t��<�5�<$�`���iT72���)�LT��f&��]�tSP�#|��)�d�og����oV� m�qB�IR��vf[9_�l!#��џ&v�e[$.J'?�T�Ca-V�{�`}1f�;�	�z�jaq���4C�@���9�ry��M�c��usT.������bv��ra�z[nр[�?�y�0�Of��B�H�E۞��I��':/������J�ظQ攨-��I�c�H�i$�5��@K�l^��Rk��{�C[
d�>�R_d	��w�`pH��3����G�2U��ٴ�5�c�0�)�禭�����=~��TmӟZ>�H1�E~t��s��2H�6��� ӈ�^���'ǋ8u�<��-R�_*�AE�|vl˧��).m�0�w(P�$��1*�>LO�d(��q�!��oZ<A4rɂ��8,!(<����c�tXt��/���"�/l��y�nB�bղ�����>Af���\�4�"��wn�YCU{̓vd��h�bK�ըC9"瘅ig0�T�k�@ 1�PUH�j��U
n�1�� �N\�K��f�� ��Na{2�C�C̈�yQ��"!�iKm�h+(,`��V	Bb^�UѠ��^w %��SN���mT6, ��� �Р'��T*q�Q������+#XC��I��)S�`��o�L�26���}<l؁tKX3 �����D�d}�'��L��!  �j�\�v�Q�|>n�ӻ[��aA��ĖG|�� ��Q�]����.F�0oG�f)�w����n��b@�Ce��j��]�6�P�"0�G�(�%!dF�,5t�E8c�4��{b��4�ðo�>0DV)���G��'��Lѷ�O�p���ᐠ]F��r��)GK��8o�E��f�v����q�4��#��cUIg ?\O2}� V� ��S��+Ѥ�z�BӶsj���m������|��'÷
��|��M�,����\�Mf�@���
��hH��B�I*68���rI�$s�\|�b�X-v�6�H�.��A"�&+��:�Ҩ20���R�i�&�����
A!8-�f��*u2�j	�p>�ĉ��$1��	)rO�Sf%,��h�KY�k� �rWdM3a��A���'��%�f
1�3�dD$�L�	��@�X��eAC���d�&rƴ��G�
1�*�kg�33B�IB�L�;r$�(�/����=���>@�ոChƯ,�ܠ���Bx�Шs膮/�Ҽ)�da��&	̢"r���A��M��]8BM���y���)J=�2	��9hn*�OG��'ij 
��q^hU���ӨJV�l��bW�M��p�P��S��C�ɝZ��LY#K��N� �!I�M��ѱ�i�4���'���G�,O��)���V���p�FS�iB ³"O��Q2m�D�<�s�Nߢf����'�D Q4��{X����֦Tx(#�X�}��8ەA4D�h�t��Q ,\ˢmٱH�L�g�>D�pK���[��q*�J�]���1D��ہ�Y���,I�h�"� �.D�8K�T�5wZ}h"G]F7�j`O*D��a�쒌��Ȓ���  �����(D��1��"1`m*BM��V�~9b$k'D��𡔅�j`��Ǔ2�TUt�9D��{0͐�
�P3pjN�S�\��/4D���ԁǺ.�t��Qf/�
���@7D�D���G�݈��ˁwKX�i�i7D��YC��m*���ߴS�@$#A2D��16�#��	Y��X�@ �0
3D�੆BT�u��M�9Z+^T��0D�H�`G"N�}pЈ��F����.D�T�Ŕ'�D`	�C��Ql,D����Y���C��Z�Ĥ��f*D�H��oK�t��,�f�����B�4D��Cp��0f�*�v����M��4D���d�h���C��K(IF��*7N3D����#K����a���S�n0q��%D��JUh�
BZib��!��A��4D��	Q,T�f�.\!&��'[�D�y��4D���Ro��x�j��Qˀ9�@�c�0D�d�e�;s�P��f	Iv�=�(�ɎNy��@(T��K�T�6a�b� �戏b�4 �CG��,�bQ��.4}b�ΒX�����=���8b������tD���
p���H�W����0bM�)�'Vp��ծ�^w��ʅcçDH>��w%�.\�H$�e�)���/����u(V)Q�����$҅:w�5󢉞�^�`���?yN�Fǎx>�rp�@�!4���I�mK�����ڭ��b ����M�V�PX��3� ��BӏǆG�nQ���@I^�s��4�zhp�OnB⢈�0|c�2N3�u�c]�y֌���S�1w���ȉ��F�$�P����!�"L�=J�ٷ�C�75�$ɗav��A�>]8�%��?��v��*_���kFFD,	�ɤ������j1�$jI<E�$�՚`�܅k��W�C�ly��%\rZ���8Hz !���"��	(�m �Wo���MǧBʜ�*������d��0|���+@�Z�:��޿B��U��@��
D�E-s���3 D�^4�����ӶP��&Ծeo��j� ˚z}�u�!MKxn@�S��)�?��'?������yOP����%�\��5��	k\Bd��$���HX"��	^�a���RQ�&���M�X֭���n�,uKҘ[�� ��@��a�j��ç�ȹ"wd��b"~p"�ūr�� �1�|{F�� 6�G�~R֟�8�a�IU
��4�x���D�"c�VQ萐x�ɄE�a�䬑�`.T؈".:����ۂaω'u@���#J6�a�d�$)�1MЍ�
<X�E	LN��'6j�"�@�%92O�OO������*`m+!������4MҲ��a�O*\�oM/�~
ç��в���Ʈt�`�w�čϓ-��M�p̪��35n<���4�ܯ#,���-\��-YsnY�@���2�'��q�S>�Y����$)�F֧����`!e=�	��~�����<�Oe��c�f=I�d�#r�pU�s��� v!��ِb���RL�k� Q���	�6I!�$ڤ�P�F�4i�ڤ�ͮH�!��'t�^�8�K�,Nڈ�7�:z!�D(1���h�O5PAPm�3F�?o!�J.@�)O9H�|�f��'kc!�d�<���y!NX���p83�R�_�!�DC<���2��3
�,9[t�L�u3!�$�<q��A�/��=ߨ�����5K2!�D�*��bbET:��PΐG�!�d��1�F4�P�@�%�B<�s�K72�!��ZP�@C�e8x�!H�&��#�!�d�s�HD
�mK*e��[qf�'�!򄞻_f��L�?+YQ�״"!� e�2�(��6���c�N!�E�P<)�c�D�@�^��Ǟ:!�_�cbų�M��:�T�@�!���!���Y=��Q��&az\H�G)
�!�DѮ{�����z.��.��c\!�d�Bv�P ߀i����Ԃ N!�Ė72�"D�u��,~qA�H)�!�䚼O�,aɐ��
wb����	'j!�T�j���'%j���c0.�O!��E���mΜf�����hU�C�:B�ɫp��!s6-���W��hB�I9D�40���s�H ����TB�I�M�����Z$f�x���"�rB�I8p� �]j<e��*ɕ3�jB�	3�$�[�'�'���шF!	�(C�	�?X���Eҧ^�c��5V�B��)V�48�� ��L�a�*��B�I�Q�>u�H��HV�̳ma�B�	L~���F�x|�&Kw6�B�	�NĐ��%�1H�X �%ƛ-\:C䉋'�!ȖG�W���� -���tC�ɸ!��D��+f��r3 B�8k��E��ĘY�u�-Ha��C�	�F%	jdm@%��Q�  �;y��C䉋qi�02v����Z�V�xB�	X�v� �C�5Mp����WRB�I��I	�A�'<<�C���$��B�I,h3�4������=��J����B�	�Q��q+`˗�f������ 2 C�I�B?�������Y�����tC�I�}�l�0�ƃI*h�� Ɖ~��C�	�z$YS	[%I#�{@ L" @�C�)� ��!5t���>a�8�"O�][�iwv�x�΋�PU���"O�<��"�?l(��]�GF�(ad"O���Q��t��]��K�1F��H"O�0��&Ӄz�8���ʏ�I�@���"O~Q!�b�E�P1CD�`�$��"O8�rԈ�x�N�+bjD��S"O�0�=[ ��L�xƠ�"Ot!󀌪y�f����̹!ݢ��v"O8ݒt,�0`9�p�A�M[�.�9�"O�9�s"� (��5Q�НD��-I�"O2] #��#��������f��"O�s6�<���sf�ԭv��xp�"O���A�E�tZHD
\�4���"OV��ġɔ#�$��MP�c~�|��"O�EpЌ��mHtA� LĄ x��3"O�T���6�j�YB,�S�.�1G"Ot����K�U|�P�*<i<�Q��"O04ۤ�ƟA��(�oHGT� ""O�II��^�K2Bm�N?D��"O�p�G��`���IW�Ky-|8�"ON�s�BC�e4ҥ��Ù�"F| "O���G�ޏ6)��IA�=�8q�"On�[c��&IUH�Co�'2a90"OT� ��;V�X�q!��m�1a�"O��E�I$ބ`'N@76 &"O��3��=Hs���wLαy�L�2B"O�L3WL�2E����Iu޸��"O����!��c�M`cH��9w6��`"Ol5��$�7�-cr̎� N	ړ"O0�Y��߳J'lZ/R ]��"OT�5�<6�;S�/e�M�!"O�	Y��A�$k�j�)U�L�F"Oxu���5,��)93��;S< ""O�Y���M�i�FE�'��;EX؈"O�<�cF�o�`E��&A'E�XA"O�8H��J�!��t���65$ތ��"OD40�%
?x3�)��I��(� "O��s���:�C���г�"O�ȸ7��xzൊ D�)]�FH
F"O����E�h�n I�c_�0��B"O0���jROy�Y���� �%�r"O��@×p^b����E�@��e"OrUj��Ԓ,j�-a���"~�0�B3"O�x&�Q�aX9͹J�bT�G"O���C��~�
`��o)o�ٚ�"O�4IB�;LB��P�%.qZ�{P"O8�
D��tUtx ��V7"Cʌ�4"O���v��n\���&���_���!G"OT�@d
��X�"��Y�k:T"f"Ob@���œ2���:a��#���"OX���]5;��0+��X�]\��P�"O� �d�p-��Q/���3A"O�����եuLp����sԔ�s5"O�L���S�H����恅|�ܨ90"O�d�w��Ff�3� �<�!"Ov�`īN <\8�B�P���	�&"O��j��ۅ=���Ibb�1$g����"O܅����o^���0��fPD1�"O�%xB!�.,�(�2dR�.Bn�a"O��c0�v�L �J�wN@�"O�͛��Y
%�R⨈3l�bX��"O�E�s+�)a.��1h���S"O,9���>>��ɴK)s����"O� �]IA�գp�~��q�{��9��"O(x���n$���E	/?�BM0�"O�`��Í_���r�dF2|uj"O }� ��N~��Zv�B={�	"O��HG�H�uN�<Bs�g����"O��EV�y�d0"�N�/i��7"OH�Ӗ�*;��;�F"2X)"Oह�&VW@ 9
w������+D�D�4��-R��qzr�μ��� 4D����̄�ZQ~5�2�߻- ���)%D��0��֙{Ȥ@��A�1R�L�"a!D��9ul��`gV�j�'�P��9��"D��y�T�".��(ۤ#n�q��?D�@��ȃ� Wn}���/�����(D��b�CL<�2�ە�
�?�q�(D�t���ǯ-�~��Q
3K�Yk�1D��3����jyl�؅�F�v$�i*��-D�dCqK��q�hI��~��@ D�4S�I*_���d�}�p�2�?D�h�E�A-|����C�	ez$���0D��X�B>���Z�lB& z|�B�+D���F�ԥ�����Z�(@pP
t	7D��	7�8L�x�b���34��c6D�P)�k�"�p��W�D,j�� D���d�˥?zP�iR+h><�9p� D��Ӗ!�_= 8���3N$���<D�\9��.,�>t�MP<zb�{#�;D�,�� W�Z�Qֈ�J�>�b�%D�h�!<ޖ�G
�+A ܛ��"D��1UF�[�>Er� X�p:�i���;D��Xd۬(C�� 1�Ȋ���,D��Nʮ	v�P�e�C�Xm���8D��0���S��P 5�UE݊:� 1D�x3�a��f��*�ҹ!�6�7d4D�`P�L�TX ��N�3�� �"-D�h[q^k�N�$-�N�����7D��C���	w�j1Z�B�w��d96$;D���c# p��xS��9Q���ul#D�,I �	"�(1W+OF���C�<D�x6O�>?e�����H���
�7D��i�C�K��9�WB�7_X�!�E5D����D��H�4e�b�4���G1D�����)	%�=�0 T�r�8(Pl$D�|���ˉE�����O�(�W� D��9ry�d@1��=P���@+,D��z����ؤ��Q'���ұ�&D���5f�f�ĊS�ц.�,ee?D�h 4I=]�6��a�N�"��`)�#=D�؊5�кp�^X�T)�&?l�� �<D��
 0�`��	!D�P��2�=D�p;"�`m�5gO�E:D�T�&J�<�:=��T
-����+D�<[G�D�9Ÿ�82MH�O�ze8Qk-D��R%H\�(.f��F�p�zi���+D�Ȋ!�S7{�>�bũI�p<(���<D��ZC�!���k��1��C�*<D��zD���+ﺜ8�.����(�7D�Tc�g��)9�V�m�X�{�5D��Q:XsH�A�-j�8�{u�5D�<3֤�X��hyAAӃ�(���j1D�� R�Y0mGd���{��	��A.D�4a� �;Ԕ	j�؝E�v��E-D���R� �
�������f�Y��,D����c�+$n�Bf�߄|Bɢ2�)D�� �Q	ui��F�P<I5���b��ak"O�2��������n0|��"O��1��a� ��@
 nYH�"O�@2��5Ɏm�%'Y2�x��"O�	P�Qr�v���	��Lzy "O������nx��c)[����%�Py�NΕ]n��k��Wp|����X��yr"P2\�$��@n�la�аa�I!�y��N k.�O�	fBz�Y�̠�y���/0w��b���H�J�fJк�y2*J$y�V)5)�Fu�(�MJ��y"�B�w����'�n��(���ynڱa`�1*�.�<2���E����y����(�&�Y�9>�yDf݃�yR�X>	b������0��D�R��y�ƅ2e6�uA7��h*���c���y�(/:H>\K��ٰb3`q�q"��y��HƝIB.�^�~QRԆE�y"���U�D��(V�f�i�-�ybF���x��n�a�@�*7�L6�y)F�
�ʅA�f�3$��������y�Q�Z�\{��ėQ�҉�p����y�J�
h��L������yA����Ex5�[O�:��gG�y2�I2 @  ��     �  d  �  �+  �6  �B  �M  �W  /`  l  rv  �|  �  m�  ��  �  4�  t�  ��  ��  E�  ��  ��  (�  j�  ��  ��  ��  ��  ��  ��  � � &! �/ �9 X@ �F �L /N  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�	�� R��g� �t��B��1�s�Ee� "<E��'�����?l�i�|����y2�6�Şw}��̞�� `�d�ǁ���a����dE�D��p�i^�;>��S��%+�|�L3}2jN,m��+�lRu��iT�y���>�����Q�g�عQ� ��Mˌ��%��|ph�9IV��1�!�;qu��UA؞X$�>�XR��V�ԎPԜa�g��:]&���d(8a�МA��řcYx�h�G��%ڧ\�ƠB�!3]��`��G�44��^�Ȅ�-J�S�d�Ӱ%�'
<�'Bў��$��Fa�,ʕ0�i�9j.!�$�!i�;��@�f�I�Iſ+� �牰D�-�Dk�;�Q���c�C�	;<�4Qd �
����'�4��'��Bm_�K;�HاA�H5���|�����Hȸ-&�tbr�Žp#��v�/�yb(Ͱ6��9�L��o�(��^��~�!�S�Oaƙ�gh�[8|`c��e��e�'% �;?ʡ��� J���
�'��s0i�3y�Bd˖��Vy~9�	�'�F��A�^_8@�D_�M}F��'����7�[�Y��:C��JF���'�*ex��N�d�B��9;� b�''��SѪԮ4	�#"K��7cL�8�'����d �el�0J�g#����'�HS��Q��*�р�	����'a�|@0l�9�0�p�A|�`<��'/x2���93�]���:%���`�'W��P��҈4�����)뎨2�'R2K����y(J�0�D�Z"m��'�~���j�$)ԡIg�0����G��O����^�E�� �9rdx05$?��{rɚ��I�m#��Q��Lm��$*Ǹu��ʉyr�'q�x��H��t��ѯ���r�H0ND$��=�3U����"��M�霂���.�69���ȓAR�L��/�B��ǭ��-����=���?Q��Ӟ6 ʝ)��^�%x"T�&��~�<Y���7?=f` ���4~D|9qM{�<����J�Fa@o�`Ѡ�sS�Q�<�[y|�d[� r:���`n�EB�`�'F�|�ڮe��)҅��F��b�O���	^���O(���b�>�bI����O��p�	�'eF�Js��#y��L�Ǆ�U�
yK�}�x�鉷4��9{�ɐkL����N4Z�rB�IlZ6�+l�	<�ؽ���Pdֵ����'] �cV�`����jG�%��9�'jX-���_�"�ba던�Da	�'�bY��R&��l�� ���$��˓�(O��5,��N�R$�7/T�j�~�J#"O�BS�]9af�K��G�Y;b�s���=lO�A��ydVEk��ה:0��"Oȑd<$�X���$Υ|����"O���t.R9ǎM�1���S
nj`"O�:AJ���,������eh�ha�"O\�!��שn=Ҍ��$�	'�<Y
�"O��#@E�U��C��W�9���"O�؀�J��}:5��k
:�P��"O�D�G@فE5ZA�Cj`D����7O���df��	Y0i؀}�~��)I�5,�,���'���ɉi����AE\���z�&I����5�I�|9������?& �S &�T|�B�	���0p#� ��� �<}��B�I�Jz��5B�% dY��T�A�6�F������ ��A��ƛRTV�BpH�>���6"OL�ke�I�Z t�A��V)(��2dU�p���h��Q#w��
T�� s!�F�H�ZC�I,A:� Iv�CQ��2�iħX+`B�8P��(��_�!�l�s�H�3
R>B�I�T=dX�!��N�ZAz���._B�	,$��rVk[	l��-q-�)
B�I�e|Lru���Z%��� $��>r�C�	0����ThW]jP��-B�6Z��#��c%O�>�ȉ0�F.`�����4�O��$�QԅƪuJ�AK����>���0ƈ3D���� 	F��AƂ�5�a �M2扃5���?�|b���b�c��$��iIGhd�<�0�� T�4+	I����a�`�'O�yB	Q�$�� ��>;L@�cc/_1�y��%&�&aYF.đ-�E �Ј�y�C���v�Pg:��P�7J<�y�n 'Ǻӑ%�0�؍qbC��y�ώ?~�Pt,(t������	�?����v\8���,�H�Pu��!i|���ȓ@��-Ӥ@+n�P�Sd݃B�v,	��O�����!3��q9�(��D���fcҖ^����)"?��,�;�2%��۷�����(�f�<���H��z�eZ�j�
1I�<��l����v����¡К3^lm��	�!n��M{�O��e�k�!�"��"bN؜�"O$Iǣ�W�$�����w���S��D�O��s�{����P=j��1���{�|x{V�D˟̄U24�K4�ҔT�X��CDP�(��:g(I�&�ݱ*�������>�rԇ�,�*I�K�J��f�3��!�ȓ%�M�adT/J�������n4�ȓ�Jt�0o�zB]��j�b���^=�P������[Ôpc���ȓSܐ�bɇ,�����ODN�ȓ&��MJ�� m=j�%)F@�م� �]Y�Fѫp'T�C��J�[@�ȓ?�,�B&@�����1FTl��b3�Y��N��z�	d�.n�B�ȓ9����[��䪧(Ų!xPl�ȓI�@��Q�(]�r�I�Z<��O6�dұk������@�]�(��׈��H $��<1ѧԗk����n�hU�ݢh"69YŨ�<�\�ȓ[�p�Q��L�r��a��_p&ȇȓq_Mb�o˗%�@$�+�# �����<_p�+3
�h�F@�3$����@ua���7���9�'A.S�\�ȓ:����<%�.��P)��(����|��6�Ѯ#���ޠg��=�ȓ-�E�� '��ߓ4�� �ȓ"cr�@�0!{�	�fΈ�
@�T�ȓu+�,J�$��P	�)+vN6Utz��0܅�P/ٮr�\��v!�h��x�ȓ^��`�$5)x,�N8�f�ȓz� 8��O�]1l�RT"�39���ȓ{/������-��$~(�ȓi<ش!ĭ�_<"c/ק!а�ȓi�Y�&T�w�^��n�%4P��ȓ*�f�K�JB�$
��R�ĩ�ȓx?�W� ❩3 �.��\��`�Y Th.���)˯vD�ȓM��R��+�:v�Փ"6E�ȓz #U�$ut�A��7-�4q��S�? ���*E��t��Ś���(&"O�"&H�8��U��e)���u"OnQ�A��r<x�D+^�@:8�W"O�h��&Y���k��N+/���"Ob�p����U ro[�[Ά�[��'��'��'��'&R�'�R�'Ӡ���J<OT���ʗ/p�4���'���'t��'�"�'A"�'�"�'�4�Q*J�$BLc񧆈aR��!��'�"�'HR�'��'42�' b�'���D��'�� �1�u�3�'��'���'���'���'���'h�v��k��<"#��>2\�E�$�'���'���'vB�'R�'E��'�Dm٣��"D*����Y�r<�f�'���'���'>r�'���'��'&����
���`}�&�ȐF.Jp��'/��'���'e�'1��'��'"�����5`�P� �R�F�RC�'Z��'{B�'>��'ub�'�r�'@����k5c@�A�*�-5������'���'�r�'e��'or�'���'��)�ը���e��Ȓ?'�=�F�'�B�'�2�'#B�'7��'���'_dQWhV gg�0S�M��˂�'���'%��'��'Q��'"�'���AЂ��t��!�,�W�'{��'�B�'���'���'+��'u�� coK==�vlz���f�R�*s�'���'��'���'R�a�����O�Ձ��	{����rrgjm(*O��D�<�|�'dv7��%{�l�ƀ�M�hX6�	W�~����d�ܴ�����'���FnM2]i���5�T���*G;��'�:���i5�	�|*��O��>et@2`�h6�IC��s@��<A���$)�'~K\�9���[Uz�	6iǃfc���&�iW6�J�y��	����]2T����l <Px�G[�s�$�I���ϓ���i��6�d�����	P^j�p��?6���S�lc��̓"I�~�����'����J*�h��q�
�#�Z���'~�q򉗤Mw��N�	�|��(_-��h�c>����>���?��'M�I�F'Uc�M�7h�X��E�ԢQe���?��۰Y�Ȝ�|���Oʜ`�z�:��/F	������G�&Ѫ/O˓�?E��'�bi��	Us�ZȊ�#�O�xi�'�b7m��r�I �M���O�P�Î�3x��Ǭ�Gঁۛ'�"�'��$
��v��T�'h���O?Z��B�{��	B1"��;e��'����$�'z"�'���'N4��� B�U�ȑa@)?�9IW����4e���)O�� �	�O��R��T�Ttʓ�̽6}60 ��M}�*s���oڇ���|��'��2o�S�]QsF�Z$"5i" �6 #�հ@OS��� H�Θ �B=֒O�� r5�E6��#'mF�:f���	��M�ЄV0�?�$Ѡw5 ��6��&�"���I�!�?y�i��O���'�7�_�i��4r��(H#��aU��*��Y�4ǔ���b���MS�'�"㘥8���S>p���?��_cpv����P�����%�z�����'M��'��'7��'��O��1;�'�0X��f5V��].3��=��'��Af�˖�3��I�T�	Uy�AѠ)�8�J�,�1��B�#7Xg}¦|ӎDl��?�x��Gɦ%��?���^h�P󐥂�Z��U�ԡ3P�wn	�Y�������O�n�?���ߟ4�� ):0 C��up�1��]�N+�heN��Ok��ɤ\�"4�CM )UC8���џl�	�M#��&<,��X;(G�s�`V�y0��ϓ4���_��yB�'"�f��	Q��]k���OP�i��W�Q��s�i L����f�G`,�xW�8��d쟒x*�D0�O��R�K�J���prCT��2uc�D�O���O��D�O1�
�l��J�l>��#�/Y��ԑ��A�/������'���o�,�R�O2XoZ%�t"���-���Kŉ��SX�)r�4P���MS�IN�f7O��$�!0T(%��'A6�I�<D�3=Ƥ��plԅGfJ}���D�OZ���O���O`�$�|�̏�Tl�x0��ڿD�⑑�É-^Л�dT�d��'>r����'�X7=��P��ǇK֩CEOۢ�f�Bh���شw鉧���O��Ԭ��s���>O�	��-���T��Ân�bpw7O�Щ�-	4�?,.��<����?a�兎l%*ёP��'��i3wl��?���?�����Ϧ�*��S��t��ƟL��(M�h΢�3gCQKG� �����'����O�ToZ�MKR�xr,�'Y��(v�$^����Υ�y��'�N��0�(\l�$:eX�h��r��!�i�bҦ��c�_6N�X[�J0D���'"I9 �Xa6/۞RTD�(�e���$��4�a����?9R�i��O�N�xC�!��ك���?4��\��۴U��v��s���2O�D^=&iX�3�'wC������.���.iW�`(r�&�d�<����?y��?a��?aD
\���	0��.{��d��?��$����FMЂ*���	�?���PyB�� RL��s)˨Y�h��[�d]��5�M��i`�7�K���?��S�n��0�'�%m�TC�'�/:���ք����N>dvčA�y��O�˓l��L�ER��tnV.j�ƈ��I.�M�ej�?1��@�a!Є���Z}L�����?C�i�O���'U�6��H�4x�r;���,x8b�N(V@����'�MÞ'�2�
�7�>��S Y����?��\� R�;��x1dn�	6��B�6OZ��$��(=���цܭDϠ�#�)
c��d�O��D���e�� J"�i��'��ęf�ŧ
d*�A�	�7H�D�G�*�̦��4��g�M�'��ʈhBF�2E�x� 4(�lA�=*���&�����|V���	�����ҟCcٗ^����r�=:�ؼ�㈚����	xy�,m����O���O�˧k��5��$��lА��k�z��'���[��v�p��&���?�g�X�L�h�c�	$1t��Sg�qΌyZ#�V�tE�'\���Mǟd��|b�= 4m�06�$ ZIO�?�b���O.�D�Oz�4������I_B�S��ր�lZ��e�ײFٶ���D�o�8!ȆU�(�IB����$�'-07�B!v�
�t��[S���Ѧ�	%�nڰ�M�&�E��M;�'�
�37�N�_���H��'"����ύ>):��DmM=��lb ��d������ϟ���^�4�t����6�ش�����3`�ܙ��i&d���'7��'P�O6��~��.��Jpn�W� e��J�ɏ�7q�yo�5�M���x��$��5qƛ�1O�D*�&�2.�j�ЯՈL��%(�0O-�S�-�?9t�2�Ģ<����?Y�a��wʄW�:3GD��c�?Y���?����d]��eR�/PyB�'Ъ���[�SgƌB�F�; �a�����Y}҆{��mZ���[��4��ԖP&�\��lG�^�`p��?�d"I5sYt�1�΅����q���n����j�Z�c�`Vb�@��Ѕ��H����O$�D�O���(ڧ�?aTk�"Gǖ�2*�0*_\�:��?�?y�i���f�'�d�\�;�4��@�b	6�`3�Ԇ��x�<OVpoZ�MS��iw�͡��iE���OXa���&���K�;��хe��k�c�0�O�˓��O��� �8|R�Ȼ���1��D�P��`Y�4X	:8����?����OZ��@c�_3k T�K&iHC-���w�>��i2�6ͅR�i>����?	Ǫ�����='j���/D;��b ��Myb���	K�=9�͎o�Q���b���ܖ��A��sdyk���5N��1��8j�X��L�4m�#e�Y��<�&��__��*G��&>	�f�&*}�)5�^�}N�<iu �a�Y��.Ò/�����Y
-��R�=P��B����ɒ+B"c��t�_/It�0���S��}s�a�3�`�7�L��h�Z4/�2-
Ψ�S���r��$��
���j�2ag�Ѱ	K��C�#��x�)u�aF&�dh��2��. ��i�5pH
9����"/򽢀�ty�ǃ$���R�F�*�����J��x��#��t�!��r�d��O&��<��O$�$�#]���J}8����pc��r_��T��>����?Q����,�y'>��@��X���i�(e����r%X�Ms��?-OX���O��� �,W�.48��Z��VӳϏ,!$��oZʟ���jy���>d����D�k��Y���B�	�^�1��G�6[�4�	Ο�P�h)�Ο4�s�N�3�"�PH�E%h��A�iy�ɰ_o*�I�4��S����!��D@�en. �C�1�Icq�J�@u���'s2���x-�i>��	�?O�<	��ܥEYl�H��M�Z<�E�i+\ŲTEk��d�Oj�d��ze%�擪%FznmC��M�MGz�R���M��JS3��D�O*���1O~��W�8}F(�v��zO&	�T��)5$ml�ß����*d�����|2��?q��y_�,j�
�;}k�� ��
;�	����ɰ@�Nb�D���0�ɼ/^�I� �,�����.����#�4�?�֫
R�����'�S�Ln��]���z�Ǎ�q��
�K��M���=����<����?����D�N��9q�E�"Ih�M{e�ۄi��J��ES�����	˟l�'�r�'qH�	���*U����0�P1dT,��'���'�BU�(i�mD*��4��1\@p�s��^a2 �������OB�D�O^��?��Y���O��-j��̤@�N�3O�D�n�Y�Or��Ot��<�@Ɠ	��O�ژV�2R�*�u�әZ�ޘ`6�gӊ�d>�D�<��s�'���K���5��&�ӖFČ�lZꟜ�Izy�&�G��0����k�G�+"���A8ig~�wD��G�&P�L�����I�2���4�s�� �q���J5 ��qF��Z� �i7�&A����޴%���h������<T�U ǯ�+GdB��e�Y���'�ҁP
5"�)b�g�	�kk.�
�fީO/b�d-	<R�6-��u ��o�ޟ\�Iԟ�����|ri܅��u"G
Ʀ�2�~h���??@��ٟ��I�?c�\�I�}$�ՋD
�^(����.r�P��۴�?)���?��Y�v�����'	"*��;�8�S�պ9-�X{b͛���?y��F���<���?��'�ڡK�&�j��h1�Zut�Pش�?���З���O��$�O��ܺ
;~&p����8�Q��>y�JF/?{�=�'���'j�I˟�*���{��f��-8H��і�i��t�'���'����O]R�s�j��1e�ac�k&��А�����ԗ'I�М_��IJ�`�X)Ec)W��lK�K�e����'���'9�O��DU2HSj�ie�i)^YQ�ǐk옼+Ђ��U.JT�O��d�Olʓ�?�hR���O��Y`jY�^���I� xѰ��%oݦ���O���?���]�.��$��@AÔ�u����t�^�^d���v���D�<)�;�B��)�|�d�O<����'��	H�oʃyS�x`,S�?����>��[r2��ώA�S�T%�-"����dV6ũ �����D�O2����O��$�O�$�J�Ӻ� T�c�� |��ː)Y*a�#P��I�b��5y��<�)��3
6Mr2(�)m1���Q�'��7���IO��$�O���O����<�'�?!��C6!]\|9��B����s���:��(کآ�s�y��)�O
tRGFO�����"Xy���%�æY�	؟4�����`�����'��O��F��s9�J��~��@Zwe�n̓M��u����t�'��O(��t`�(+C�ub��*��p�r�i�b��"P�՟x��� �=�eج�� �R��i6]+U$B[}"J)n�����O����OZ��?�n3n�Ti�B�Т]A�H�G+V�5k.Od���O���;��۟x��薍I��l���p�����Á�u��%c��7?��?y/O��č0 ���Rע1�����W8hp�"L�Q�7��O�$�O|�`�I�2�����Nk�pa�DJ����]���8a%^����ş��'�a�;V�S�@"��R�<����Dߕ����5�M#����'%�N��E����O<����2&��!Q��@�4�Ȥ�Ʀ-�Iry��'Ɋ ��]>9�'i��L��S���@)ȵ�(��&X�R���<i��x��u'�:@_���)���T�`����$�O4Ha��O��$�O��D���Ӻ����uQ�	¨}N�{%�Tx}�^�`Q �/�S��>Y�=�WnbqF��Ge��s�7��J�z���O�ʓ�b-O��O�3�㍶�f �����2lQ`�l�q}����O1��$�6$j�MS1��)\'l��6-E�R��n�����'A ��V���͟��	\?!�k�"3�"5#�M �8����MD1O�]�-�]�S˟��IS?Qr���Jp�FP��(;�J����I�(r�L�'3��',2���E�.mZ��&T���(2F�`�I��R]Y 9?!���?+O��dP1	"p�� �+�h�����m%p�0 �<���?����'X��Ͷ��4�5	H�RK���3�5V�� d������O��Į<Q��m#��Oc�� C�:D��cL��)�۴�?a���?��'����W�'�M��C-"$T0Q3�b�3�U]}R�'@RX�|��� j��O�¡V
|�pL)R+�/2�(��P�Q�6M�OJ㟌���n�dYW�=�d/h`5`�@���S�� ��F�'5�ݟ�з#�W���'��ONШ���V�K�(�᪂??@���=��ϟ,���G�%��b��}�Z� h��i��G\2�R �'j�g��>���'$��'���[���Ky��D6A��X0��\�B�tꓷ?�v�F�y���<�~�U7Р#'�Yb��袀��Ǧ��F՟<��ן��I�?�����'<�bt�X
	�F�y��=I��aӆ5:G��E�1O>���
b��`��(W��ܴ��6v)�|��4�?����?�ˊ��4���$�O<�ɴi���@!��)�`�h���*��`�y��*�~���O����mJ� 
���y%�G�m6��OR1x�C�<!��?A���'p�kӬǚN�P FK� eҝҨOL"1�G�%��I�H�I^yb�'���*����:#f�'u5ʁS)/B��Iޟ��	����?���<��h���U�no��kgC�p�F�y҅�=D��H�'���'��	����7j�S��IŖ�j�04'��<"�KA�	ۦ��	쟀�I@���?� "� X���m��"	Dͺ�m�_>xa���n��?	�����O���«|R�'��h��H�6t~6�ڠ�ZhcLd�ݴ�?Y���'�Ȍ��\�����hօ��"%�w���`�H1o���'l�$R�[��柼���?=k��̊��gB�-�=CR�α��'�B�2�̅��y���A�i\�p4��a�� 4��Gp}��'��$�'sP����@yZwF�P@@]+=�`��ٵB�HS�OX�$��W�P�a����I*&&� ;��V��3��&x���f�`���'{"�'�T[��S���1QH�K$�aQw�o)��6	�/�Mk��N�S�`�<E��'.5BD͇
QpT�Ά3gyL�a�jӈ��O��$۞\;���|r��?��'Hl ��H/r3�A3�ɽ�`�t+9扼6,� K|���?��'a��a�H9B�P�6�����4�?A�,Z����O\�$�O����;Q�����\�4�j�	gH�>�Q�+�Y�'���'��� [rD@3GF��[�]!uI�䳕���vGp�'���'���D�O<2��G�`���g�]�1-	:!٦M�������ԟ�'5�@�iH�iץ.����%q���c���&zțF�'�2�'��O��	
W�� ��iW����\�w�b{�CT�7E�� �O��d�O&ʓ�?i!�,���O�L6GߓV�㓊�\zƱyq(JΦm��N��?)g�Ů��&��P��[�(�S� K1]Tr��S!c���İ<���P�Ȭ )��$�O��)F�]E��c��H�Ƣ�'I>v��>!�7�f�����p�S��!��|;v���dɣu�p|��N����O�}Y���O��d�Op�D����Ӻ#�/�2�쑪���3}xrU�O}r�'��`�/L����O��uiӏ-&,vu�i�H�"��4����i�B�'�B�O�����L]n��0���<.����Ҝ}��$mZn2\#<q����'�H�K#hF��V�%.� �F!��Af�R���O��$������'��	���S�? ©G�x:$TX��0����i�_�T��@f��?���?G�٬ǆx;�G�"/Aޙ �� ���'OX�QdJ�>�(O\���<�����h��|a��E[�:�H�}����y��'���'o��'��Ɏd�䐀T�d�����0<D|I`j���D�<�����d�O��D�O�d%,ܡ
pR<���V]��E)�b۵�1O����O���<�H����J4'̺�H8>�9 $��0ěS�t��dy�'���'��D
�'6N41�o��T�v�� �>�@ [Emx����OX�d�O�˓Lj��7Y?u�I�A��̺tN�b����
Vz���4�?Y-OV���O���D��[?1�㘨	�&����
>����¦��I͟\�'�����"�~����?���k�6��$�y_��2��m�.O���O6�����IXyRݟVt���Y0��Pp*?�bR�i���{�V�R޴�?����?��'#��i��A�L��dXIU��P�XREzӚ���O���d<Ox��?1���U?t�xE�G
���@ɵ�V�Mc�cR�/����'X��'��t*�>�*O����'J�'��T�]0�
)R����U�Bl��'�H����;U>X�B�ۥa���k�ɧL��ݛ�iz��',�0{�$����O���2'��80$NI|7&�b��=��6�6�䄖2K�?9�������-0w�����wL�=C���WN�A��4�?��cϰ��v�'&2�'yrb�~��'\b\R���)rT���'vR�O6I��;O���O����O���<�	�2�0JOR���<��d�0z%���S�L�'��\�H�I֟PΓ]~�}�B����~]`�mB;w�aQ� u�h�'���'^�U��;�����EL�pm��'�2}d����M�.OR�Ĳ<����?A��-���n᚝#�4b$�x%	у���U�ia��'�2�'��	']�p���~��Ɛ�sg�L�S'�I�4�	�i�zu�w�i�B[�H����8�ɑ)Z�Iu��<`	�!�`��F^��+@���AG�&�'T�X�ȳ,
����O�D���%��(Ggr�I����'r&��Ћ�u}b�'�"�'�RQ��'��'7��2pڬQ9�Q"�lջQ�3>��^�����=�M����?1���zP_����ZM(p �!�Xs��	�:7�O�dœ`��>� �S5G���Qd!�F	D(XGMS�P�(7M+)��ioZȟp�	��H�S�����<��'^Nk��J�-��?��(҅�yB�'��N���?�ॏ&p���ш�	U�!�kC�L���'9��'�а��>�)O��D���#��O�r48����
�S�6�Oj�Kbr��S�T�'���'k��Y2ɑ�-{��A����囕T�&�'S@IW��>	)Od�Ĩ<��{`�D�q���Y��R�V!�@Y���T}�K��yB�'.��'�2�'E�I���e`(0��˶@�#X d��۷��$�<�����O�$�O��e�X+yH��!_�^ä��SHL��������Iӟ��Iiy��B�,�5
,Zp�N-lHaR���
�Z7��<i����O����O�t�2OkV�>5Xf`�?K�&8C@�&/��V�'���'��U�t��˟�����Ok,�	��]Z�N�It���b���)��6�'��	՟H��؟t��+g�@�O�%k4���s���p�kƕ!2���"�i�b�'o�ɉQ�����D�O��ӴL~�ċ��ڥC���@�lP4p�'���'ҁ��y"�|�џ6�+vn�@��)z׌Sl���
 �i��'�h޴�?a��?���|��i�UP�#�������?=�T`�t�r�$�Ol�Yb7O\���y��	B��X�8ք�Qz� a�
6E��Ĉ?d�6M�OV�d�O���SS}R�`xgAʟ?��X�$n(l����/�M['�<�K>��t�'6�TRU�B�X�0�J��R�w�r-���n���D�O�������'��	���������`׭	S����N���QnZ�'���ٟ��i�O����O�q��7�ы���4N�]�AȦ��	�Ʋ���O
ʓ�?i)O���8���N_N��˃-A�w�}E�iI���y��'���'��'(剗&�@p�ݩojfxaf�I8��-PP���Ī<Q�����O��d�O���*§xnD�gh��0!��NY��D�O"���OF���OV�@Ԅ��d4���&�E /�6L��:.^�+7�xb�'e�'_r�'�.���'�d��sĖ�Q�`�9W(߂ h$8��>)���?�����)���'>���n��(	�6rT� K"�8�Mk�����?a�B*A�>9�脍$�+ �.2D�j�a��ʟt�'vLA��&���O��醍V~Z�i�m��b��Ÿvn�\&����˟���˟�&���'op������\�Ҝq����ml�PyB)�C�6��F���'��K/?1�ŝ6P�*jǖW���;Aj ٦��Iʟh¤��$���}��&�`�@A�ã�io� 4Cͦ�fꒄ�M{���?1��R�x2�'��<����J{�i��3l���2�M;��<yM>i*�V˓�?�p��,�rdr�CE�R�u:�#yٛ��'��'��	k�@;����l�"���Ŋ�0x�h!�F����>	֫|��?Q���?�2�Ɍ�V�G�`N��r�b����'�����)��O��$%����0� K1b	�e!�c�Q��\�q]��xdŏq�IƟ��	����'�b}�c��%0$q��c;�(�pcZ=?N�b�@��W���D��ǀ Vl�p!ȑ��R)�t�fuSQ+P�<!(OX�$�O������M��|�S�T' `�'MΞ	�7�TB}"�'B�|2�'�H��yB�s�0s�L��E�}�b��;0	�OH���O��d�<ѥ�נ[\�O�\�b����3�-	$	R<Z*`�"�$#�$�O �$Q�Aټ�d!}�՛=۠�3�36�9�D��M����?q.Od����^�۟(�ӟ=����A[��Yk�(+z��J<����?���^���'k�	T�hz� �4+�:�}��Kh�]����̓��MK�V?Y���?���OD�)G�@�	��v<�~�K��?��`�������OӪ�#�[�$�ҷ)�#M\rEi�4g�pu�i���'S��O�:O���=���ƁV�cL�-�
֤jŴ�l�˴��I�Ė��*��_�$�4y�dl=3�"F<M���l����	��d�c�����h���'���U�pH���f�.e���s��U��Oxa��d�O���O����G���0%��d#� R��A}��A�(k�	zy��'{�'?j��4��`b�IՁ�>`�
9pű>	�/q���'�2�'��X�#�_�	��X�e�0P�2�;����.���C�O����Ot���Of��
�Ƿh��u��IH7H����ri	 +$@'����ԟ��	��p��6���I�h�J�""E�+v�"XD����h	aڴ����O�O\���Oe���,ڛ�˯S��|ru�W%lKls׬(����On���OB���O�P����O����Ov�zSf�ɀ�ֱF�pY�M���d�Iڟ���.B-�!G �$��I*�,�7eP�>�bu���ԛ�'��W��c�Ϟ����O$���f��'��~����!�%7۪Uz�����?qRl�"��'��\c���!�`Ͳx���S���F�ZQ�ie��'������'�'�b�O��i��2��
l��!"C����/yӄ���O��z7�C�<1O�����M+f�d(��A�ibr����'�R�'5"�Oo��4��n�\Q�!G-{Ŵ���Ɉ1l��6�F�8�S�������r%A\8�J�ʅ�'�0�r�V��M���?��"K��Je���Or�I,��$��	 J8p _(oc���+0��ݟ���ӟ��ȇ�u�$�˱f�'�¤�C�_1�M��Y��h1S�xr�'�R�|Zc��)�#�0a�mqP��l�F] �O
�R���O����O&�)M��r )�#+�D�p rr�	�I({��'?�'��'>�'��80����Q� r�k��0ܐK����'N��'�R�'��H*D��	�� c2U�E%Ǜq�2]z�h�(���'�"�'��'�2�'4��:�O�E�`鏭b٢����/>;�P��:��K)u�N� cn��<��e�g�+���4+v�W4ct��thR�7��C"O��b�[8jJ�p��d�
]
��O�@c���@X� ��hiw, �Ӭ�>2Rh�D�p�n��E '�X��;f�I2O;m��P�c�0Dn ���9i��@2��85O>�"'�%*@�s�I!Y�t032f�&h"���b�H�(l�5�G�-c	��ˍ �����RDĀ4��%� |B(���ų(�HC��'sR�'��H �c�2SȔ��;P�N}�ǝ@J����nQ=���S����'���gMT{NTW��I�@D3�A�O�d�ж��)GJ$�S��?)�L�6��6�s9�wfћr���G������ڴb����"|��WL��4��o����s�@��̇��5.v�iW/ƅr��pA��1#<���i>]�ɀ{;ލ`4�V4
�(�!�,Db:a��ٟl2P�XY7B$�	ʟ����!YwX��'u(�f��a�1��)[�% �	+�a�O�ܹ�G��]�~�1�Ө����$��*ot��S*0ehep����Н�?yq!��l��@�����3ړUN�ҍ��JC�Q�����D��|�m�d���˟�F{�[�t���M#�Z2,!��q���%D�4p�Ԍ8"��uf:~ԝB�	���HO��Ny�\7mD	��KabN�5���2���ef���O����Oh���@�O:��d>�K���6)-���?2T�A��G"}4�цL�@��t����Dx����k܁w�Z�2
54��Ё7�C%e�p|�!�AZHj�"PO�Dx�`�!��O���Y\6��@�.~��m B���-:(�=���3U24����0f����^�;!�$̧v��sw"H�t(��Lƚ;��@}�Y�lB�
���O
ʧ1�ม ۟d��k��άGc$@fN�?����?�4�9U��a@��^�.�����i��L4�X�̇�R��4�4�˙�(O ��#�t��+f�,4�' 9&:Ţ#��R�`=ză�3Xt�Ѣ�(O�,#�'����Ł+��hl^*'n�ԲC���I���Q���
3a�_d�C �Ⱥ\�6�3p
=�O(%� ���Q)Z��U�WK�zt���y�P@�J�����O�˧:�da)���?��^���դ��,kv|�"�>j$U�`�4k"ع�`õ��E���	+��O���k�b�NL�A"܇!��4��	�TZ�I
l�yQ��
@�:@�Pl%���q���I8�=���¦KK�۲��x����Iߟ���'��h�V�	�hJ�|h��@lH�2|x��S�? �4b�%\J�Hd!ߟ~���I�ቭ�HO�8�t���˛�u�l(�F�%T^v���2��¥d�>�	�� ���<�Zw���'��H�5�P�@�􁰍=g+.�R�'֜�k6fZj�R�o;O։�q��^d<�ӔcQ"���%�OXI�p���(x�Yv8��H���emܟ>gJ��E�����=g�r�'TўH�'B�h���M�'�F�;BA)�nu��'�d�2T�%;|ΰ��L�� gX"f�)�S�TV��{"	��MSu�Rи�"����p�P���?���?���b��Px��?��O�`�bu�i�B�A7?�Tk��L����F�L/�p>y�!W��dΰ@��)���פ_ݳ���%A�|b�
'�?9$�i�:H5!�yC�l�2��6������s�"��<	�������'u|���b+�IQZ��
�!���;n�a��)>~1*�0 �̕1Z���I}�Q� ɂB�M����?1*�X���;� �F�K(8X`�J4+8���Oz�DCPOZ�ڒ?�|���-r�n�����
?iRe���Yb�'�F�c�E��h��500�*H.��Kbb�6�������:��J��b�4�?�*�:L�ӎ�6(�!��a-�]H���O �"~Γt-�tåw0eXg*�D�,��	���X�s�����l�i7%�R�� ��+!�i���'	�%xNʀ�	��͓O�f )0&�>���`�L@�Dy�.)�6m?�|Fx�,B�L���sg)�� %���I'yϤԳG�2�)�矼�D�ta��eM�#����B-«_C�Y�	ǟ�*���'���6jͲ��4k��E�8a�౟'���'� � �h �x*b*va���Q�����:~PD���ڂx�(��ߕ>����O:Iɂ�
4B��$�O����O,�;�?!�!��P1��̨G���"a�I.G>P��� 	��e �T����sdU�P���z�(((� Y��FJ�#a�����?𾤁�R F��h�'�*�B�$˚xq����O��ԟ�	�<�'�:MGJ�g��A ���
�����';�y��<��A�I�4��B#�瀅	���dͤXf������Pu#��?��i8��4ܚ����?����?I�b�-�?A�����4I6ܻ��i�м@���cm<�p�UR�����vO�=�횫�M��B$oj�	1���MnVU���{8��QU��O`�lڷg.�F+��QḆ�a`���� �4�?1(OL�� �)��M�M�@es���x8X+��j�<I�	���Q��Ȕ"�Bآ��<A�Q��'`�A"Oc�R���O2�'j[�$j� �5���@���`z��!�V��?1���?����z����D���ݮu�І�<_�S�\����@ 6����>zv:�<��^͢#��$���gQ6f�(i�O��di5`�� �#wY�@����$��Qs�%m�T	n͟�OL�0JAdΜt�� �3M�,	��'i�O?��i��)��aI�Z*���E%'cP���O�I�sf�LX���(-�4���E�=�2�I:�D��RN���L��H��4!���t�I����1a���R�����f�&ų�B�"F��(�)�3Z1�hQ��&:��i+���0т��5�rxy㕙%��4<���s��uVz�����2=,L۰/�<-����EE�*�*���)!J,wި���:e1l)�猒A��qDx���'�j�s�G�qu�cI�)��%s�'05	�$6I�áN+��b����F�����'�l�6fF��`�v�BG^0��'BrO�cO a"��'�2�'��"l����� c��׎����]�=i�,:S㥟��O=�Zx���&�ȓפ� wV�t.�OA���/?X���n|؞X�6Wt�3�O�Ƅ ��V���$�=3�t�'�r^�x��I�LZ8�)�*�~\��%�+D����J�0X�4y�IX7Ű�H�Ȓ�HOT�'�򄝆+Yx}o�%N����9y�e0"��V��<�	���Ip�����I�|" aU<B���4le�)��CւW���
�Q*t`����*}���0
����5���v���Q� U*�:�OP���'
n7m�B��`�Qhӳ1�J\9UF=cƵmߟ<�':��?��Њ��>���dF��ER�JbO$D��94�i�H��!Ϛ,#����a��j�O�˓����R���	}���H�!�y������A�$�jb�'#��'��˳���7�b��?0���T>mhq�!��a(WQ�`�e�=�x� �iX��(�7+L�3atX��c���離&`v��3�W��2M���H��Q�8Ѐ,�O��m���O�`t���>e��T�K!vl���'��'��a����g+��AD�N�qz���-���� ځȓ%�7M��u�$���}118O�m��o���	��O#6eH��'���'�<tr��>FD�A�+@_��#�	�w���y�b�b�0�ņ֐�������Ͽr#Ͽ'5!�EEn�%��M?]����iDW��� �Q��������X0q��4�Ͽ+�S>���ںx�(Z��D�2���s���?Y�O�$��O��ð�F2h�`����Eh��9O|�$(�O�Ұ@�0.�W�H8&�	��HO˧}.My򧜓vJ�@��D\	dtR��?�GI�&�*���?y��?�Ĵ��d�O�|h�,	e!<Mz���?yl�3��O��O_�$�,�@�'|:1���K hKU�AjW�}X�x�'܈*!n�B�hR	��:���$$̥ ��@F�REZ��H:��I��~��Y�L�	by^#z��=c!�c;(�b& /�y�iR�+P�l`��-]4���6���3`�"=),���O�N̲���ã��2�ЊU�W�u!�$,�JaY�D�/��Y�ċ�'��Ј�ݭz����@�L>�	�'r�ՠ�d�'�$Cv�,HX����'9�[��ۻ7tҴ��A¦�r�'t�R�Gٿ'�����ɪ��L��'�HL�#��X�R�8c�_yZT%"�'��,豧L�p�4$S�b@z��#�'˪��u���!�s3.@�EM�9�'@ͻ�Cǃ{�j�s�W��HE��'�2�h�*z��r��	_��i"�'y�*Ǭq+��
��^z"I�'eL4ä�yy�L�ыТV�����'$�4(%�L2�)�F��i;�'@ް�g!H�~'
��9<6���'ʰP)�$���,�'��/�Ƹ��'ib�ˡO��v\ 7���/Ɗ���'f�=5jSpK
���V#��L��'���X�+$$ykF�0��d��':F�ir�S�$�H(%�ʏ�de�
�'���a N�:7�����"� R��
�'�<p��IŜp���;�
��B�ډ
�'}�P`Q�1����'� 8��	�'��pz�OYP��7��,ZN %��'��b�U>5�6�E�Pr}c�'T�!贩��@H��3V��Nш�'�b)��V��E� Jb��'��P�Ǎ�@���a�ȭy�p���'��:lˊ&�(	�1k@
�,R�'�YeZ�Q>�A�ں�H!��'�Be����LA$�À��qO��h�'sL��CC�+)v�0�>
yR�'R����L�;H��w�3/����'�֝!��۲U�4���oOK��*�'쌡��a$k9�D�1���K��	�'g�u�e�1o�=
6���mR\$v�C����*�� �"�E�@�6�~*4o�$W��ݛ-ʺ�b6�E3u�T=��Cɯ�B�ɻmJ:������h[�Aa��	�wi�ۯx��ic�X�r��E�G�p�
��b�"l���D>_T�6`�%g��b4g BKax"�ʔaˬ88b`�y�`YD.�a�|Q���A*
hʜ�EH1}<�A�5Y����܉>��{B˾;6MJIH45�ҝ˕i����(꺄x'�N xA��lߖ	��B�392,�������rR@<�"咱��;��  �"O�!�!�1+�yr+�:NiQ� �*f�BZ�n��c?�mࣰi�$XG(Sj��g=A/���wl�B"�/Sv\A	U� 5�TA
�'�l�@E��58L�����-���6H�(�?�A@�('ΘӴ��-ԭ����\���u�d�+d�y:s�S&%�p!`���Maxr�é[U��S�3?���k��*v�����oK5l6$�!DI�X�$�y"�ܭyu�u��nSZ��{���5�f$1�GPT����4��(��䟀@h*�eQ-5��pA��®`��)H"I�2��A.�"mԍR�%@����I�����*�"O �1JL�����Ɋp���x��|cD�i��A�{�(A���3&!�5B�|�&�P�޹λj.�b����*���c�5+�����x��R�^{�X{����+lCD���ڿ��GT
�݃GK]9x(��S�ӎ9��d�$��<<Ĥ��x�:�D]����K\
=p� "��T� -�n��F��:oTɻv)���O����N)4꬀�J��W���ԫ��^�KQĝF��Tp�&�
k��h�Q��P�@�k�@�O2������Z����~ʟ�y�f!'@���jM�L��r&���;�"�>kX�� �@NO�e�� ��%����FNd$�ӭi�bZF��M:N��GB�W�^ݘ�'ց%�X�ڠ딿8���s�D�R�עE��=K����<z��dI$JU�,Y2#ƃT�.� �Q��c�|ҖO?}����u�uI�
8V���`G �y2�KD���
OfpF}� ��Xb`��I>'�2F�\�B$���M��!��\TQ2b���R�J��>ͧ!�-���i�|`#4��(ZPi��6y�0Q#�V�'��i��M�6=�`��b�k�@pg��S7
�(���Z�\��"<i����lá�O�)̧ �esn�>@���3���<6`�	p��J����9��U�`۵"�����0�%��8��O6����G�4�����d�� q�'�I1�J��$	�[��b�D�����g>}r'����G�V�
	�U:#�¡i��+1���b�}Z�O���B(��y���) ����R��O4 �6c�+�ܼ FCO��O���j��?V !{�J��zY�i顉��
��Su���'V�:T[��i�N����@��>�[#-Κu���p��H�'��)�ÞuR�[�񧿫THW�t^��筙^����e�'p
�ϓF����s�Ox`�I�!��Бd��w��鷧�|�p���n� ��$y��r���"� 3��|}���=y��%�T��H�(�NY
$j�YIz�IH����'����2O�*ap E�2',I���vh_ g:����_�Xd� V:/�批N���&�p��/-�l��׼\o���RCYZfe�+�p̉q�H9k�0e��m&O�-@�h��(�ޜ�E��S!*���"$�ى��ݩT�	F�O� 5��fp��:sBϪgޱ�P�R����fb��s��~�;}R(�q	�ML��jǚh+P0L<!/ĮuQ�D[+>�g?Y���i�|�jφ�\<��#H7;�l Yp�YH�:�ꑄ]����cآ+LB��cK�
U�F|cq�	(8XQP������5?���I<Q����/�n9�JJ��'[�5�͂9#���%�����J����C�+t�@T��m�>�X2�h4�	>GSv�#�i��3hjhF��X�l�B�:���6 �,1�!�'�����#�����D�yشS���p���3!�}І��o�P,���<�$.�	YWʤ���G�
L�z�R>
b"B�I�D����ɝ�$,�d#�G^�m��I "H ��?��'��$�K��5U��;�*��I���\'ga}��ۙ��ᣢBO�pW�h{%H�/J�T��b�y�������:a�u��B�0yޔy���5}���P^��"�vqx�j�K��hO�%@c$�7E㰄��M< Z�Ђ�O8�(	/b�e�+i�t�8����p�1�)֐I�ƽ��A�hX��y��*9b@d�2�J4*��M/?ɰm��N�hUr���uO��C!Oh�T>�Y�f�K9l5j�Nɣl��Cc,D���eY"���#��,L��|�p�V�hٖ�#v��+x�x�䧘Oش���Nͼ��	]Ė,r��Yn�����[J�<&�(%V���+�"0��NN!�P�-O����@�y�1�1O&E� `L%|�F���A�r�
��mR�M��U�CdD+���"#�_?M���,h���sL�1<�^|"�)[b\Hˆ�~G$��	S"�j���"2�\����H5E*a�5-��V��, ��9�U�T�"�&����,Ox�	���	UW\�x'Q�#�kS�'	�\e�H�J<��W#Z�RZ��p`��=��a`�G����'��A 47O�t)��;J����&����W�'픰��G�e��z��,Ą������p��(c���PK<���$F�m���~��s�%$@�L��E��<%���G�A @h�4|�D8��J�?>���E{��2LHl	���L
��� A�i��!"G�մ��� �
x�e��'�Hm���+�����O������0�1h1�׫c;�h��+��&�,�/�OJ�C�A�xn��W�3>��s �T����:l�d��C8�ɭ|
��qp睫R�`�7O�
𼋵f��:���M�u�4 P�D�Dҩ[�Bڧ:��a{���:|
�y� +��a��H�Po�,϶0Y�G�/�d�7�Q̱;�(�"_AL�Y‏8?@�"<��2|'��#�@�A���0���<��*��&oT4�L�g�;V�|X�L�O�=Hs�'x�ћ�읪܀�a�dJ�HN��2(2�l�iA�H�D˦����)2 ����̎�I�4O��6 Hsl�kE�O'!�u!� X���)d;�aے'�;_�R@Zj���@��'�"#�<�P:��˺
K�����yr��g3���0����~bLI~�����`�0� D�Q%�|��s',?�O���2��9eqP:�d�	j6�Q6A1�^���T'�&����O������^���DQT&���ˆ8�����j܎Q�<eK�(Z>{s�D�cg�/u ��	��ĚY+xȒ`a���O�-B�-	y�Dri�:a��8��E�O�m��� :.YIʷ,�|�#�V�V��%�$��J�@��3�e�+�� ��JY+2�4	���<�R��X��%��ZQ?�4GV%� ��Ӏx�Ĉ�9elAq`hELBX�;4�'X�W�t�'dA��,T�:�F$�vɏ
�<��I��y2jU0)��x���ہ�~�_}�'��@p �M=�4�K�)B�Z����$G�y�! &\J��"�&À D<�C�#v�������Y�pE�y��Y�p����'�(q Dξ?a��G��N�T�áU*\��=b�Aѳ1���R8@��P H�P��;D���cr ڱ%E��!RZƊ����Ǿpx����A:�"���ٙ�h�i�/_L�����<�vL�xJPQ@�F��e�@D�4#�-GT삣%$�tHZ�T���ي�9�
���_�d�'�X�^����x�H�������: �
�?� ��3~BX�a�V�Z�v�a�B_��X8�/��X6l��!e��]�*�ϧ�?�O3|tcKP��a�׆�p|��X�N��*d��a��>��y�F��j��ҝw%�9��%6s�CBگNN�S���\�Ra1�'������d;-��q%4w�A��dƘ� ܪv-ш=bt%���O@��0���<A�Q�J�Q���H 
�|�B�.C(�(�v`�2��5X�� ���p ʛ.�6(�$N�EɈF��P���` �B5��Qc']/�H{A��y��(P��<u��T� ��W.�}��'ʔ��0�ԃ�#��8E(Z1�LY�M#H<z�I�8uz���NJџ c�&�o��XFN̙F�д�Vi�0��f[�%dĝk�I�(K��]z?�O+$s��T�dvn��΄;i����s��;gl�Ke�!jn�xB�ߩ��&e�咀EL�Q.��G��_����(^I�����O��P��� qbi���W�,p����/�i��X��k�Qq��P��;ѱO4U�%�^��
}`��B��Fă�J3��J�5����m��)�B�ծ�4m���Z'���OR6�ؖ&��*Hъ�<Q4䆣3����U�n�9�� �2�n98��	@ZD�2ȏ^��,E��O �Ka'S�%���j�	ְP�À
R�T�2dY��[�6`	�G�L( �?��d��`H���9���s���#/͖	����j̰0����G��<���~��$�p���MzI�T/K$	T��{��]%9i>��C�l4q��爠2�k �(VK@��b�4Iq����B���n�H�G�/p��'ڌ�"�?�� ��9'���Ks�!+^@��t*�AȱO<�@d�?o��xg'ܫ�yu�#�T޶%���5,�`���A��e�lY&��4���D��	�*Cr,��Ot�I'�$�B��-���f$�dgr%rIX�k�z� Ti�:.�r=Br&'�U?���йV�ՙp���ӣ�$����+^����1<<�FR;`k���dI�F��9rV"��oy��Iǀ�9��uh���#�rI�O�0����Ӻ�I	��H�� 1���A(T�D��2ʝ@�UX��U�b���$@�.���3Q�I)@�x���/,y�����6}���I����#��d��'̴��\"E��秘O0������e�k���4<�ڕ�jCV�6%|����%F�� ���Ȕ2R�EhK?ٛ�j�H-���d��3�p9�㗝)/��'��"v��|����V�t{J>au���:�0���WA	 1Xq�,w:��B9�l�S �U����|��O�T��&x!C���lb�x e�?%T��e�4؎�"��' �&�����sU���h5A�#Fxv��g��b�e��� �O�T� n��	��DpMJ�qt��D�
(��-�B�4��f
)��%�:Y�L�*!1�ё�S�6C�������I>��4H�
�?��>���&,�E����#�"�^`I�k��4:~c��X�!��@H@3lZ�0�Iy�-�N��{���1�� )f�EB�(�M���D<�s�@���	���'ڞ��կ� *�dApH�>f���噎}:��C@��eK����ԟd��D�%8����Ї9v��A�
��ɧ~��ʵk�l8������O�TI�p��|q��M�_��� D��H�����<����]}"��=� Y��ɄSw$�3�w��̇�ɉ{���������%kL�;oNV�Tx��
��~Bϑ8�r�'�.�S�s�((����U����S�ǎI�Tj�F9D��+���<Gi�Ea"ǐ�hC�@9'�$D��2����#s�! ����֭"D��J�a _Vn8
'���;�Z�3�H!D�D��́� [�hB�G�&�PTzfI)D����� �|��aÓO�$y���3�H3D�D���W=}��ء�*�m���{�!6D�8H�*�dT�I�B�� d���5D�$���f �i�1�6>"U��B3D��zb-���G$ֽk5D����=D�\1DB�7A��0���֨k��S��8D���p!M %f0%�U!p�$+�+6D�� eD�i���sl"^,
yP�.D��29HB8X�h��
���q��*D�\a�Ȟ�~�"�����L��f�>D��Ö,��h|��b��R������;D�0Ic�Ǖ�@JD�Ҹ\�<����'D�T�2>�Z��+�d�"�ԋ'D�0��@��>�X�!�3 T%P�%D�h�ĕ� �� �eM�[oм�G�=D�`��0h�4��A
2粄J�A;D�� FU&�QZ�\��eɋtW��"�"O�Y���X�y�*ɒ�FҰ�q�T"O|���![�=����6E>~� ""OlD9"E�|8�+�#�p��Փ�"OΡ� ڙH��%�爖3
���#"O���n�*U�ąsM��y���"O�L�uK��.��-�j�d��R�"O�$�n��	�H�l�4�"O��K5n�T����kP���<�"O<�iU*$&��!���F�y.d��c"Ob|S5�������ؠ/#Rl�t"O*!TE�)+}bl� �x��c"O�`��F]�f��c�O�Mt�t��"O�H8qaB�xG �a�?!tl��5"O�tg�	Cl��Q���2Uz�"OZa��!�L��@�ћW�r��d"O$�bs� �����vyZ$�"O4��B�I

��:�EC5�u0d"O���5͜�k.p{�B�[���"OFIٶ�]�V&J�2Q�ֻ�(@h "O�-�@�0��բ�8��#C"O�9�(Dp�
�ip��4YmʀY�"O��h7�u��Ta��ݐ;g�qV"O
��'˪P�$8���Ī&`�� "OX���c�\�~U�	ԥk�ȡ�"O�Xhh���P��ʵ
�t���"O2	��d@�,��BP�I�;� *�"O�Р��̆ � ��c�3/((�T"O�h ��;7~���K�8:�0V"O(,���)#n<����u�'"O�1��A#N����KJ���4"O8�e熞�܉��n�<E���s"O&,"���]N@C���ВE��"O�X$M�?H$���:�3%"O�@��.�Tj��_�J��q��"O�\��A�A�Z�'h��p�d"O0j�	�#+��f(v���K�"O~���mD�\���SA'p�h��V"O�8��-��4�����F�	� с"Op�p� �\ �h``U{n"`�U"OB��ɦs�.TC�ɂ�V����"O���I:rqV�Z`�T�87��ҕ"O.�ɑ��~Ѫq�I,$��%"O�H��H:�| �kP�v^p�"O���Zd�و��t!���E"Ol�s���9
9~h���+i�T�S"O����˖����q�D�U�b�q"O��[pG�7��}���[����"O�E��׶..0�$�D�X���"O����A@Z����4 X�ӊ T�@ ��G�����F��	:f��psB(D�Ȃb�_�U(����`,�*��2D��a�BÄ)�V�b/��ee^]��%D���� U?x����ԍm� �*O�����.]���QR(#�^l��"O�xy4N�B~��!0���x'"O}�ra�e4���`��xV�,�Q"ObIZ��s��t�X�j���@q"OJ�1��F�����ԥiyN��Q"O��Zc�lC���hH�DL�D"O�p꓈�50y�Vǔ�:��s�"O6��3�&TJv��� �"O�q�d��;M�0ՙ�$B+7&|�(�"O�Z�`�?P�B�b �?��� "O� v=������>���� ���{�"O6ȸ� L*�f�Jw-'��@�"O歐�iP;2�h'�:^R��"O4,�!N�mQv�ad�<�X�"O.x�� ,�6�D#��@"O������b����[�.�:�h�"O Pa�Щv<�h�A�;���"O��4�6�`a�����e2b"O��� #�%NuxXYe㐨��la�"O䩢b�]b-\��wO݂D$�Q��"O�p`��J���H��I6L�3�	y��$x�2�y6���W�Y�f9$���0���{�D ��T{�ڶJM�y�E�6����(�
Gֆ�MC-�y�";���I܏M��L�%��6�y�$�=|v%�1BʟKT�`%�G"��',ўb>mcB��j��8BUm(W���� D� � G*��0�K��4���F D�tˣk֭"�����o�gȔ<pwL?D�H��
j���z��|fpRР!D� Q�IB���0����y{8 ��=D��(�b���I@$�Qur�#&<�Ir���'zA"�ᗄ�
�\�3���f��\��y��0g��Q�`��F��i\ ��y	*h;qG�<d�e�Pț�@�ȓaƆ��Eϋ�^aV�*P�"l�|��s��M�gg6NeP�����Nu�i��~�whN%L7*A���DsE��������Q�)M�I�t'�<����H���R���`�A��A�������b}���,hjn����Q<h|%��o��y"�ģ������
�x�B�@���'���ډ�����s̍�#xr�(��O�oE�iv"Op})V &�cr* 6���z�b8�S��y"��_���C��Y��#I�&�yr	��0�\M�%�Ʋ���IB���yb�[h����JJ7#\ɒȏ��?1�'4�ږGC�Y�ސ� o5N�>x�'�Z�Js@�;�b��WkT 7�Z	��'��%2$�\. �廣iJ-EGN\�	�'M�Ab�Eڸ�P0��ʦG�T�q
�'2M2҉�&$Bp���6:C�4��'�(���OG
� QʤE�4��,��'p��&�(Mj~Bs�-,:�T1�'��5��WDm�x�'�S?+���"�'ԑrDJ/ ����V�Ȏxc�;�'٬���-!�v�*���0C���
�'��-�Vn)/��h�E/.}N���'��1Rh[%P�^\�`� =4P����yb�D�K�|�	D���w�8�S�b[���'��{rFڐ�d�,��i�ZQ�@
,�y�H*�D�AJIgY�]���� �y�F�"+�]�fc��Q��ŀ��g�<�͊��0:�X=D��̈b�N�<��&U�L���dƼ�U��h�p�<i�i�&"�����V�{^&�ZG�p�<)f�5m �*���}���[�%h�<�p��p����7Cn��@n@Z�<�a�M���,�} ���4MZn�<Q$�ĜNc@���� `��A�f�<a�V�{�+b�N�fX��A��a�<��/]�N@|Zү12N(�Dn�^�<���F�'L)��Ӱ|[�����@W�<�RX������Y0B��M�dh�i�<� ~�e
�(�:a��Y�}D����"O|�5k�� �\��H��U�}S�"O(h���.�4��F��6պu�"OT0ÔZ�	�@�+�l�l� �"O�x����;n]T�8W��8h���'"O�Qr�@�]&x�P�;� �`"O��:��[����[�I��k��`�"O���E�4��Ti���S��E�"O�x���#_ےu#5oQ�4���"Ox9Ʌ�Mb�����JM$��2�����ɫc�:�����iŤ��3�ED����-��ñ��Q#_��b8�W+B�<L!�$K�j� k�^�(?��PCː
w!�dI^JraQP!�"U& \[ظ~]B�ɻ>,$� �
;��� �'g��C䉛)��is��	 ��Ur$�M.@�C䉴;)�]�A�0)H֩��aF3+!�C�ɓ M��)>^X3�k��9��C�:>h��Ơ�9! 4�"�o�bo�C�	�:�m	X� ��r���`ש#D�Dq�i��ʌ�tO�[l�"�e7D��SS�Kf�ɻ��
+Zb��Ӄi!D�w�:B���S�1Vn��a=D�T��^;a1�e�r'Q2}q�҈&D�`��k�>X�40�a ЄRR:���%D�|�բĔ��i2P���E������/⓷蟊08�JP?EЅ�s�RqF"O����?F�̑Q�I��.�ɶ"O����o��dH����-Z�"O\���ו: Z���@�hձ�"O�h�F�O�c/&d(��t{[���'H�k@
45�D���!�-�H�[
�'V�=S!�>3)�aRuc#T�I��'�.�Y6�$|��X�sJ���i�'Q����*O�.I�����Gh8�'�\�pd/�:8�2��# :�{�';����x�,8YU��Hy0��O�eҲ� V �Yu�L�Q.��"�:\O���SkW�>��K�	վH!B(1"OJ�ZVD[ .�"e�c#ƥ"4|I6"OD�k�nA�.L��hEn�F*OF¢n�,*����M�|�pp0L>����߹a4�R���Dv�@�f�Tf!�D�	��H�ªN"yp�؃I@�"g!�D��-Dx"f�/+�ndـ�<\!��$���]�{�hp���vG!�DC4�A���	{�*��'>6�!��!j�=c�\�f�>]yCa"~�!���H=�ɘ6���"��i�%R�A�!�� RF(�r��<JP�8���h�!���>G�.�i�M^��S���^.!�D��p��Y�����V$�#J�6
!�L�_�0m����y�����&^�!�$�+�`)�A�6m�A��
	�!��L;$�d���I�W��j7� !�D/��m�G��E���<!�$�#4b��H� n�L�N�/.!�D�(v��1*�%$X�a١�R%+p!�D;r��� ��A�c��	��Q�fY!�dP� ^�8��L"R�� ��� pT!�):�m#�F%nǾD���ɑBT!�$%ր�%�Ѕ.6DI�o��V�!�D, �L A!ď8��A�7^�!򤉶_7^�J�ɣ$�Db��7!�� T��C��<I�L�Fo]S0hܐw"O>@;��Q��έ��˴,�-q1"O@hs���|�����%�=@洼q3"O�X ��� ��#����\�)�"O�[��[�"V���
��e��"ON�HU�Y)��THЅ���V��"O�@���6&��:�D����"O�� Đ ���kC�;5<��e"O�ěe��L��A�k�5>� "O�Ƀ��V6(Y�p2� �~0Z�"O�CH��ڹ[���5��A�"O��a��0yy��2��%�d\�"O�5@TlV�MJ	�4�
����"Ol0Y�`˥|{zL���4e��;2"O6�UA@$p���V.Y1O���"OF��2ɘ7,nPl�<3���"Oҙ��J߻цS��J�'}��"O�2�s��1'I�c9��"Op�A�QA+��%ܞ!L>��"Op������I������`�V�y�"O�� �!"M^��R'UɊ�P�"O�	+�U
*�I����![%���G"O
����"VD��Z1Nȿ|�T��"O���p�C& Ѣ!z�m_bl��"O z6-��> ��B�R
)8@��"O8hQU�޹f���;Ao!Q ��0'"O��gk�$w9�-+B�D�欥�G"O,IX��<�h����N�r0"O��#G"ԧ��Űb�T;޸��"O؍��cFj$�ъ��I�ꀓ�"O\A����3S�f����ơ)����"Ox,�UiX � ��֮-%l��"Or���O.���*U¶Em�"O�9H�F�h9F�c P�H�FxY�"O$M� ��	��ur�@���c�"O�0��'źP*�8���8E�,2"O�$�4�̒A�jD[�@������r"O�ر��}n��2E ԍA����"O�}�ޒWe���& V>0��S�"O����K�faT	�j~,���"O`�ĥY�X� ����-OO��"O�h��+R��ft���t�B��"O�u���{��@�7���~���A�"O�l0�ˎ5�Qa@�1jg���b"O� �� �!Զ�S0��)X^=Õ"OvyꉐG.����A.T`�E"O%�q!,K]>���C@�w�.�W"O<P��$�m���Ӣ�U�x�d"O������hb���z�X��"O
!3�'Bh� H�(��a�"O�`�ѕhv�Q ��Z�d��X�"O�X!���`���(�D�#[w��R�"O"�@�.��ݶ��ʺys0�:�"O2Y��#ح�bPyg�D���d��"O��	"��dy0���	~�C"O��Q�q����d�E??p���P"O��#��%gP�<�!"ڸV��!�"O<`#&M�Y*Z�X�+���ԑї"Oج�7�3���ь˖k\�!�"O�!��п[沈)��H8v��"O�d�T��JԸ-h-kaB�[ P;!���ge��Xu��9�8P#ÖE!�D��qpv���\=O�����"�P�!�]��:ġR,o�ĠT�#�!�� �@�`ڬ|'�$Ё��I�n���"O����ޘM!
��0L�>z�Fؙ!"O��g�� '�T�DB�
�
h��"O@���I�O;T��i!Kk��""O�����B�cȄ��Ađ���"O��� ���|���@�.4���"O:�zE̜#�*l�S�F|���"O��	tiO:%�p�cn:�d(�"Ob�����D��U�$AF�b"O��rӌ�b�h���,^mZ�\��"O�`r�63��U��63> ��2"OT��r}3jq�j\�i���c"O�ixtNG���J�Iɣ'��I�f"O�=�F�9_�(1Ί1rz�+�"O�Ѩw�ǩ2Ϣ��NA
0��@g"O�5�3�w�����G����"Oȝː`�|�hĊs��ܘt8"O&uA�%f��x�NJ/RqĬ��"O�\�sMÃ�dB%΋�m���"O��׬�0%A�l�jpF���"O�sr��lc~X�P� EdN�"O=;I�)/,�����,# �Y*"O�(j��O�l�+���	�'��P ֠B�a��!�gD�k�����'��m����B'�����	jX���'*�$X��V�h{ (�7�8\��	�'BZh�Ǆ�!|�"I����[����'�ʹ��` �!:�`v��M�����'Dh$iԎ�^�^�U� �[ ��`�'�f�
�l̑>��U�T!%d]�X��'�v9�(ͯe��0\��!AF��y2BP�"yY��PBV�L�S%�1�y�[�,�*�g�7P�p�9DD�1�y�E���&�t)�Ӟ��Cd��y�PE5��������� ���y
��Ԙ��i����pUL�y��T�x<�����wRz|ՁӅ�y��	e��肓�]�޶�H��_��yBbT�k�,PK����E"�t#�"*�yҩ�d��l�26~��A���y��K&e����k�>4�V�
�E��y�-�
���B�ɀ�)���a��y�Nڣ��E[�S�q����yr�K��	#�E^�����׋��yR֞$��Ó�"h� K.�ybkR;E$ʉ��	�9SZ4`#`ś��y�l�$,U��1�mȍG�3rO���y��Y�	�4*���;
*������y���$Tl�`�D�06��z�B�6�y�Z�r��c�)6qn��4�K��y���/6b�#���Y���sM�y2���jd|��ςIqf9��)?�yR�WW�	�veQ�*��3!�6�y�i�&c�)a$pEXgʕ;�yR�S�	ɫ2B��7I���,�y�E�"�@�JF�4�uk��y���kR!�*̾ 
,�KӉ݉�yr%%T{z-�r� t9�(do�(�y"���
S25���'؂u������*�3b���j&��thH4�8P��3xYbn[0kv:Ѣ�ojh�T��3�hř�L�t| �AAA�B�d��ȓ�tQ��$)�pk�T5:ҝ�ȓ,�XyS��B�8��5)1���S�? �H[�#��,�m�C�T�(��
$"O��)�N�n��X��âH�|��a"O|UY�#�)=5�̒a-ǡrK��� "O��ZwÆ#OJ9[�␇W�db"OР�׎ِ6�0��s��&U
�"O8��C)ۤ��E�a�턘��"O\���NK\�Nak���ky�,��"O*Bq�{�pȢ��5j�!��"Oꉲ֮�#-t`�XZU���P"O�l�0�N(P���K�D�A;̡�e"O�ahe֞�8��%J�p'����"Oaу�<>vL�Eb����"O`�kM�M�
�̍g$� �p"O�	i��ݙi#qҦDC�u0B�h�"Ofy
�N Hy��F.�ry����"O��@�˛\���a���#:P
�"O��3�^G��\@Q,C/+�r��"O&<��υ|�N8Y�k��T��`"O�d�gD��>z��4쀷A���aQ"O�s6�S�
��AZ�4*CNt��"OF�I�+�.S|D��wD$>�W"O����J�\0#Û�"S�)R�"O��b��Јy�lҪ7��L���2D������e���P1a��C��4X'�1D�A@0.�ɊP��b�r���:D��)�$ҞA��$���6f�+g7D�$���T�CĔP*P�K�_J,0	`4D���Ă��c��P�aD�P�$�8'�6D� ��1S6BT8�N�>D�2`n5D��� �B�W� ���$��hqh.D��{G*��1zc�Ҧ�$��T..D�� �)=T~�xC�N�O$�M0D�d8�$��{9~Bf�t�c�a-D�h��ʛ�w������G�Ҭ���5D�0�W�J�n�$���:��rW>D�D����#8L���# �`�C�D=D��L�-Y�� �Q@!G0*\�r�>D�Ћq�&o=>0��ˎ�)�^`pu	=D� �����LI�KN/h��0c��7D���G�q#~�����{��0W7D��q�Թ=ϼ��D�K%t[� 3�c5D�8�QZ�H�ᣡʛC
�t���'D�����7b����͚�	n��`�%D�Dj�'�VH �
ܝ,p�` �k(D��ڐ��B=�Ex���=Nr���h!T��S��,�v�*���}XN堡"O��r�`��N�Z6MHN�cc"O�hH�(��LQ�F�Q��"O��E	�?���
D�	
/6x$h�"Ot3�+�i2�qK�N�1 (���"O�xɒF����#m��F���G"O()��l"���W�\�U��"O\�W捰�s�*��講�"O$|��ab�<���1���%"O��;r+^~�D�bX1q�v83s"O Y�qo�H��p# ��"O���`*R+c,F$���K+=^a[�"O���f�"M����I,�i��"OP,���W�l)��� �]�xb�jF"O��ҥdʽKX��b�4o���b�"O�ꖅ˷"S�i�0��K���;f"OM*��*1D�#�!J�q*1B�"O�"E�=���c�*�/�iC"O�c� �9���P7bfuy"O� xm�R�ϽN�!��#��e>@u"O��sEьMܤԨR>I(��"O1����0"d'���"O�UqnW�x����6sF\3�"O�Ti'�%L��{C�7c��l1"O�a )D�_m.<pGÇfʹ�1�"OT5�
�	FA(2h�M!�AW"O�8�-Eb��uJ���g!�9�yR (O~(C�_z	�)?A ��Y�pp肎]�d�Ӈ�'�q�ȓHXL�3c �<T��k!��:M����ȓ(���J��t`��  /�Ф�ȓ,�=aƏ��J�q��=�bp�ȓhti0��L9�ڄh`�@NV0��j���8e��&i�������:)�I�ȓQs*$	�i��jn��,�
6nN���9��)��R�*L�q ���1��e��9����2'�H�L�y�`�k0��>��XH��{Vj+U��6�h�ȓ`�`$��_va#gL�<��ȓd��y@BC�XM��r�~���en4����[|�����id��g$<��#�'B�h0A٬ ���ȓZuD)ذCZ�غl�ƥ#Z��ȓ]�1[sDW�jC��)$C�si��ȓHW��n�0��5��-+xE���ȓb�2��Z�6I�󮑪0\⠆ȓ{��=�$ڞ`c���j�%^��0��^Z�jD �j�T�Ɯl���ȓ"�Aiɠpq:��R�%��q�ȓ�������`�T��� &��ȓP*i��/<&��w��$c+8D���FѺ
y��P��F٨���'D����g�%����ϓ�#v%�s)$D� �be �+R"��e�V0^E8�(D��BPC� 	��|�7��\Q� k9D�(;G@�f읻�'X�Gx@]C7�8D�P��7q����&.B>L�t��e*D�����@SHn�a_�N�~Isub#D�
�ǟ+g]l%P2�GL���D"D��e��;*�L|��+�}6K#H D�� ��T6-u�htQ��3�2B�	%3�a�a2[$�X&���j�hB�	���rV���Z���`tKA�2zDB�I�j��E��q܌+���s B�	��x�j�N�C��hU�U%C��C�/HV�P0j�6c�PÂ�7w�C�	-6��!f�WrR&�"�gM1i�C�	� ��i��MuZP��Ǌ�Rr!�䕯F��p�g�5)>`XÁ�K5F	!��*j`6��wΒ��´;6�Y>!��
�	Wʽ#��N;[�d���J�d�!�ی�#�M��D\�'�I�!��n~������q��p��!G�!�LRα�vG�/�ȍ�w�^�#x!�dT�j|23+±#�m��EE#a!�Ę�?��ت� ��Z�C2�� 4!�$'+����eJջy�n�`DR�!�#
$�=P�Cة ��@��+T�!�(TNp�نG��=�Iw �2v!�D�?e�-�E�^!$��%�ńʢn!�K2�4�0�פ/��$K�D�MW!�d�ZWLI����+\�c��&et!�L1�>��̮<��4���*a!�� ܠ[qi�M$x뉵6���"Or|��C�UU(9�R�Q(HPIU"Or�i�-H��ٵ�^�D�����"O���W��x�z�E!�(��p"O���b,�R������ݠ "O�u��O�%@��J��,b��}�"Oj��w��;l|ށA�mC&�x5"@"O��0}H�\��� pu��"O ۇ�1yz����Pm�H��%"O������mi�<;�!*�|�R�"O�``/ɇy���C&`��-v@9:�"O>x����,�%z�n��Hp蘀""O�ʖ��vh#��cP,�f"O��r��(T*�sg�M�b�qh�"O���gH�1n`az�C�2G�R| �"O.h`�@J�*�XAl� 4���'"OЈÒk �%�Z��e�P�xf��	%"O&�J�+B$Lk��	�hd>��!"O����F�#�j�P5*[=f�`C"Ol4�P+=<^��Qd�"}�^U��"O��z��,s�4��"\�z�8R�"Omk�7�TuA��4A��	Bq"O�ٙ��R�|������O[>1�"O��@�K �l )T@�6=2Ԕ+�"O��ƭ��S�<�Q'&D=Bb�"O(�0G6zE�X�� eJ!��"OB�tz�LDQk �Ax�� �"O��X"�J�%4�U��*�kaE �"O�|�p��s�Ω�I1Q�	�"O�1���Yh�H��j3��*w"O������U"@�X���h.�=z"O��Ȥ� 29��y�M���"O�{�@Z d�x��ƤA��"B"Ot� &��z��#�AB�#0~d�"O�P�ui[@��6��3��D��"O2 P!��Q�՘��?`�8�c"O��K6�Y_ր=+��+~��]�P"Ot����ҰC�W'�@T4�D"O<e*TD�X�t�%�#�eX�"O@���LM�j��ݠ!�4�"O��H�/���;� �>�B:�"O �����2-QP�O c@L�#�"O5�f䕑C��A1A�W$���p"Oh\��L�e�l�L�(��+$"OH1�6`����r,ċ-1^��C"O��#���(/����g,�r>�Be"O��	��K4*���ؔ+!e���#"OZp���%�nP�Q*�*j��B"O�9���p,�%�Z�p�2��"O�����gH���A��
@(�"O�9���H�V0g��
�`��"Ol���HA�Dd����U:#�́��"O��)��/+����[f��e� "O,m	H��6��x!�"^�{�����"O,DB�C�0B���RH�!'}�"OJ�a�J�u	:2$��?�%�"O�I���<��J�]�6��"O��'mM#BT� 2���8���p@"O4ɠ�6�*qq �҂G��T�4"O���$@ &7V��h�+%��"O�]���j�I2�'ӕ\$xy�"OtHx2��;l��s)&�,xG"O��R���↺t2�p5,��y��hB��Ȓq�LA�D ҄�y
� D(
��R�U��@���J>(���p"O||�	۬M��!
W>�)��"OZ������b%I���/ ���"O�\���	�8�&\:�Jǜ �ه"O� �V��(h64ԀE��FwP�"O��
#��\�⸻��#A2`zf"Oa�F��+�Y��J4X\
L�"O̽rІ��-~Ԉ��B�'U�]QC"O t����#	�TH`���T=�q�"Ol��#+X�vgnx�u�́5C���"O���"C-���Շ��|B�"Oeb�bԼc�#�ʓ%��Ke"OD$ v�R�Q��:�-ˍTTA0"Oz��&�r���cf�Z([V��@"Oe,��EJt�1��Z�lX�Hc"O����L�Q?聴f��t?|<�d"O��	�*+�=��F�{<l\B�"OT��	���P0z%��D��1"O�|�v�D�b��	���9;�Qۅ"OjeѲ��p���k�#V�L'	Ya"O
\��%T�%���P�L�'LL�"O�9A"Ì�1N�C�t�d��"O��Em½;������I��R�"O�p��L�3'�)7 ���"O���`�&��d�& Y;4B<Ҧ"O�ȓ�ψ-#�N�Ғ�Y�T �г"OT(�7��h�e)���c*>��b"O(�p"��1#�a�N�:#��@�"ONq�6���
D�4,�0Ph4Лu"O���R��:!8��pJ\-&R���"O�� +S��F $>� *1"O<�8�R
	� ��Ś�`F�Y�"O��Z�I޴Y@V��$.!�����"OZx�RFѠrt�N,7D�t"ON�uBшy@2��B�0IH���"OP52���1���� �~�hhy��I�<Yce�	_S�:B��t��� �G�<�ƈ�;Z8<p O@�Vj�a�m�<���K�M`�S�Jܟ#�6+��_b�<�+o*�Lم�B�YI�5h3��a�<�2gU+<=��`�c�l�S���D�<	'��RG��x�BP�).44�A�<YQ�U �BUPp�q6����Ji�<y��ܹ88�sIP2�cejLd�<A�I�9�"��g�X][���/�u�<��)�	_
]�4kH�	�l��`SI�<�&�&B<\!��LBvH*���J�<����3GD���f�-ЈA2���^�<�ǡ�<XZ�Y���O�B,r�ŔE�<���%�L,~��#��K; B�ɡ	ZR Y�+(��iEm�740C�I#u��0�e�,;�����j�RC�I�j��T'L=qP���CD�#T�C�ɿ9���+RG�� UH��F#"s�TB�ɚU��m`��G��0|"b�!�hC䉽S����w��?FJI��T�
B�I.�h� �n��+f�YuEߵ^x�C�I�D�50R��r	�`a��$�`C�ɟ`��)3�H*"s�-ha�\�ZpC䉇ac�ۄF�n�he�H�JC��zT6�Ȓ��EL� �W3�8C��?�0���7!�ʗ6	�B�	"NP��$f�� pR	5ttB�	�k��9����[* �� ܦ�4B�)� ����ʖ1���C ����hV"Oh�@�NۆF�ɐ�$��%�* 0!"OP��䇚�c"�2��ShЌm��"O⠐��-0�}#�(/���Q"Ol��eM1��2&��3F�*���"OЩ�QG:4�l% 1�?d�F�	U"Or�U�^�ҝ��LU�Y��D�g"OP�QT=P8� ���1�ֵ��"O��MŧD��4C�jM�K�x��"O��g�^TF2MzSCK�}�x|kU"O6�UL��d�0�	�k�X�B�"O8U�p�	8�:��NV\�["O�Y���fw�[-A:kh"��B"O�\qGP#9]]{��'gD��v"O�}��D0A�,6��;Y<F1�"O,�a����X�!�F �~Y��"O�}� �X�ب�Sd�0%���`"O��	��<?Kv�Ȯq~���E"O���F�	�W$Q�҂��0D� �"O�H�6.��cιz�B\e��HF"Oh}���Ex�S*
lbR�h6"Ox=cĀL�Q����V\p����"Oީ#���oꮜ���Zp�]�'"Om�R�/T���g�#=���8�"Oxh��Ps4��/�^q @"R"O�(476��$c5��,s��`�"Ot��)o@t��-��|xeZ7"O�MaRL�~���٩(\���r"OZ��0�ՠ*���Рb�>���8�"ORx���eJ)ো!@fB{D"O(q ��@�Cܼp@���#+�)S"O�:g�I�0�@�����,�8�"O0�{C�	���HFCϗ�<�PF"O���"@4{�t=Q�O0jϰ +�"O4͑@�ikTZ�$Q�=�t��"O~x�W��u6��:�\Q�ޑ+�"O�c1L�_o��qEB	:4�"O���4���8u��	g�j}	"Opٲ��W?K�r���ו@����F"O����b�6B�N4�iĄey4�Aw"OЕ��X5q����W��k��k�"Or��AG��_�����> ���"O�@2��ڪ;,���ϊN��ib""O������v�Zl#�M�Cά`c�O��@���C���!�Z:`5x��O��=E��h^�^��RW
�?6��Щ 嘠r!�D��^�D���B��;��l:Vĝ.&�!�$�I)�p0q#�d���%��`�!�	��<3�'I�q���	�3:CrC�IpL��!G�	"\gz4B�'ϦbrPC�	.|�af�vǞ`K��
�P[VB�I�O�� ��9vo�`�dȚc@B䉺L�9H�G�8X�α�*H�@��C�I�jRm��L2Ҿ-ZT���} �B�I�	l8�GiN+, ��) eO�ۤB䉄3�*�0Ō�vl�AsB�L��FB�	�o8�x��}q�-Z�˖EB�I;#%�h wgP�y�\3���:1�B�ɤN���el̥U����GI�`�jB䉻D>��ir�E�2��i� ��d�zB�	�D�r��Q�mB�(B� C��&���(@�M�F!�i�,y�B�	6p���M�	�Ţp�ǒA��C�ɷ,TІ�Y�R%Hh�QjC�>-~C�)� 8$��-A8��})$�<W��h1"O�a�� \O<ģ��IoQ yK�"O���פ�F���bK�%��˶"O��1�[2k�P����s^�(��"O�U�Z$^��J�&y�IQ"O�A��d�2��Q%1l4dI�"OHᩳ�_�\�� ��3n0�	��"O0%`�*��B���+$b�O��zS�D���L���n�z0�OC�ɦKцDLC2S�, ��3�C�	�$x$Bf�,�t����s0�C�Ix�̸�J+&�m�u`ݟevHB�
���ڧ��^+�0C�nΟQ��C����mc�O*h�����?R8�C�(P_x��IB�6��H;�bݳ3PC䉝47"9j���S�Z(����"fC�I�)'ڑ[�d�#h�:�c��[(q�"B�q��`�/Kb<dL:` �B�	>vXv�P�	AX<��d&�2,~B䉊u�|,bS� 6W/��i%Kg�C�;[a�92�piة;%�@0.�C��<e�$����-j?���Ff]�B䉜QQ���	c��M��I`ŮB�	]#D����ހ�8��D/�B�ɒ�T�nĢa�*d�p#�=s�C�əF��,��!�⬅���L���B�	�C	R�A5������F#��C�ɼ/�6�st�O/t*�e�G.�-O��C��,�@zeň�8qn��v)���C�	"M؊a�@a֌?�2%2#N�:g�C�I.���7ɖ�\�u�䑥V��C�-kyI�NȦz)�`��	�*iG�B�?�69H�
�[�@�Ѓ�F��B�	��H�a���
���v�H�0רB�	{���§g��w��)�AELg�C�I��8e���6�q��&P�Ou�C�ɇw��Wd*d���ǁ��:���"Onq[�(����k1&I`|��JE"OV�7�/s� tb%Ċl^�Q�"O�癎hh���Tg�*Uء(�"O����,��Gz�Ձ����2`��`"O�xA�/׉]r���LY���6"O�0�Aq �)q�a��{G�Y*"O�ݠ'/�>:�T���H�~6*��'w�	ß�F{J?�i����n� ��j�,��cg�!D�T�� f�:6��8Z;���3>D��e�4fL����uz�z�;D�l�0�Ӹ@���W���Cp�f ,D�4��EA����-e�J	JAl*D�p��"�7x�#�IL0%� j*D���B�-�<�ءa˝`�%ID�(D����,�(s����
�V
�Őv�'D�,��]#p#�48����7���i D����+*�A� E3i�@0Щ!D���d	+�`x�+j�Fp�£2D�8hB�:�Z�{ !G[/��K��6D��ju��q�(!�D c���Y�6D�x�`F� n��8��A�T�f��M2D������B8����A�4�H�E 5D��x����~�CF)C0L�f��e�5D�\ꓮ[�[u�0��+-�e�ҧ0D�����T�UF�A���&7H����k0D�hp���uOȵy��G�#��a1D�L�:D8��`9i$.�e!;D�� �@;��X~�ђa!x���"OΌ��/\ _��`�Gv1X�"O�����(k�L���/T=��"ODȻ��\�y J�Q�A��0AB�"O���
�M��D"
3,{�4rS"O�ĉ#�M����*Ƌ��
��X�<��%A~&�i�r�� T���)y�<�`�@�z#R\y#e�'.x�!��E\x�<V$(X j�:$��[ʀ�BN�������FJ🜖�(OFX:(�I�΁iA/Y���u��"O�9鱢�6:g�����Gq���"OJ-U�T4B���#Nu�!b"O�e�̗��`ș�'WҠ2"O��H�NY?�8Ě�CJ�b�� �u"O�� F�e��Z2���w@�8!�"O��XBV�&���S-�9Ƥ�u"O
E�6�z�B6Cƍa�R��T"Oj�v���~nZ�Aw���H�t"O�i��X��ۓ��#R�l��"OZĂwč�1_�E M�uO4m*�"O ��r8��%/>�d�U"O~�@tǖ�OKJsUY�@m�)��"O�M���( ކ��lB6$V.5z�"O6Y�6ֺxn���@�ڎ��!h�"OB5���" �hm:�*��#�bh2#"OZ}��	�Bt�cu�(M �[�"OL9��

7rD�8%j]�7H�8�"O��fF�1�HQX�J��I@Հ�"O4�E�(�N�0��T>f1$H��"O������ZNe+ �±6&�غ�"O|�Y���.g�شz�K��Xi�"O"��"eT������%0u'�2	�'G$P���6V����쟒;P)J�'e|p�e���pBd��tS�'�jYr�O<>�< �s'�'H� B�'X�"�J�(r��K�%ح=�j��'�����ڋH�ru��m��4�e�	�'�`}��6 �����:H��t�ȓY`^���O׿���q��M�[ ��ȓJ�ڈ�0E8L_P����Gh<�ȓH]�U��<I��-h"��*掅��O�Ԅ$�5��q���X
����xh(����!R�m�0>�ćȓOq�`�Έ�S$(局)S�^vPل�e��m��/+q6Ĺ��޶>�2!�ȓ!���q�l�6c�2�괣Up�L��m,8誄�:"n��R��0���ȓ� �;����0͂���(Q�a�ȓ"�*=�eHVx|���S�$$�@��ȓ���Ñi�'��P��X���`��-h0��ʗ�� ����ȓ�Ȫp�W��$�'a�F�z����걡��̀��E`G��#�y�� x�����D6'��@�_=�y2�CTpQ�Є>56�yG*��yr��F�x@)CÁ�zFD�2F�܍�y���im&9��A�:��4�"D*�y��0l4�T�(٤���x@ʱ�y��6�\4`p)����rl��y��S�%5~Q3"�آ�ؠ�fGG��y�OU�6jb
ط}�l��ڄ�y��=f
�i�H��}�v»�y"���852�*J,�- а	�-�yr'��*���ie��v�2!��ɉ�y
� ~�J�fF�rդ\*f�E� (m�p"O i#�j�9i:��s�Ԁ	l�k�"OH���fJ�B`�Q8�fյo�a
�"O��9��ÂD���i�T��!�U"O(e�g��;�.5��cһD���k�"OE�2I@A���α@����"OXQ*#��޺��B��<yq"O�F(�Ll��D���
"O�Tۦ���De�|�&�Ȓ��$"O�l��GJ69�L�3k!?�Z@�b"O` rs_-6`������6��CG"OQy���_�NpPs�՜Y����"O<My�ↅ6:tH�6�ķi@�d�V"O��3��W�5���tOl��"O����ۜV��yR$�\��`�"O4�Y4��Yhb"b &���"O�x+ n�W���Wf }t�)*�"O��ړ,[�:v��pdօ=frp��"O$EO_�'��R�J`�t�`"OV%�e��T8��K4HPb1h�"O���%�8u����+Z �<���"O���o�����@J�m���E"O<���<Q���w���,��|��"O�\3�O
?/�)0��G�@|�t"O��%T���3F�R�wA�4"O�	�P"秃�0	�����17!���<rH�Z���m��	q5ρB�!��[,e����?U�b�#��g�!��uO�z����y���W�N�`�!���^Q61��I�y
)@1�R�6�!򄏓S����a�M� �q�9 �!�ִ]a"iJ�X">ʍ��F�v�!��S��Ҝ��h����K��!��{�|���J&m�
�d�8J�!�Œ_����' � J�ޤb0#D�Ar!�D�hX�H���  ��0f��MC!�@�X`&k�,� �{s�U*s?!�7[ ���M�R�$��a�;!�d@���0	Y�WL�(����%V!��ٳrt���U��"q����47!�I����7l�?1����5w!�D�y-����
��)h&�Zlh!�DL�]˴(�b/�2�ƅ��B�&"Oƴ� kC�JH�@z\$<�u"O��(�Q�d��`�� �`�"O��C6�B�ݐ��=�$]�@"O��@2"K�/5*���K����J�"O�%�fm�4{����k�d���r�"O:a�	��@b�[���c��2�"Oz�3��z������C��${u"OB�Ѓ�]�8�Z *M���C&"O��)u�ݷFd�YIR���=�!"Oh����))��+&h�)�0���"O�\ȇm��W���hdɿ��YJ�"O���I�?^&^,����R��3�"O H�V��;K��|�t��"O��X��F1e�pe3�'ݜ;�Xir&"OҌS���/!>%�0F5_�� ��"O>�2�=�r���BZ�K��)!�"O$ ��ϕw����0 ��?�<�I�"O�륅_�t8�,H�n]2t���E"O�If�~��!W��y�:\1�"O�y��bK�@�����A1q��|
�"O(�+�i2C�\��"A��$�
�32"O� ��� ��G�Τ��"J�Q!*�x�"O��[��!M!h<����c4��P"O�a���g�t�$�'%�P)�"O�-��C^�`���Ġw۞�8�"O���1��j����N�	��Y�"Or a���N�X�ʢ͍�_OҜ�R"O��� ��|�@���.FV|4��"O,�����z2�@�>a27��A!��Ў����d�/e�0�øm !�$N
}����!�� ���箞?2�!�P*y��(��ȏ�o��!u��J�!�$��e����K;j����J^�j!�D�!{�����.ʹbb}��hEA�!�ޞL�T��1"�W�lbN�T�!���9Z�4��՞X�`�`&�7|!���7������sm�����,Fa!�Du�dGS1[\���KR�$a!�dN%h�0;V��)3s���֠�?;D!�$�)i�޼�SM�|y.9�4���j&!�$��t��DƀM���@G��!�d۟.N�y�ň�.`��)� C�3!�䊉��T��ڸU8X@ѯA�V-!��"��Eڲ�[)b����
	y�!�� yByy�i��);R��6�._�!�ĉ�ac�	BF����Z��T�!�43�
qA��B� ���!���!�DV�;	$��o�6��|Q R�!�1�h���&]���yJ�L
�%�!�@�sjt�y�a��+�6����!��W�&�±�K�Z4 ��M'3�!�$ _xpx�j��i���y��߭'�!�E�PPa��W�Z�`5���8'�!��ö_�<P	��):~V�R-ڸ`�!�
w���PsE �zt����Lխo�!��ٜg��E�e��;]u���ťP�!�$�3`�9F�C�8��Axe c�!��ք"�04걤���x(�!�$�)q�ac �h�(�c�����!���"��	��	�)S ����[n�!�^*NTtZ�@ �>�����N�!�U����7�M1��PJ�8T�!�$S2���se��A���(T(W=I�!�DŇ5|x�qwM�.��t �f̽q!򄅲\��ڤPol��&�'qY!����Z!����pT|�p�d��+��� "V,�d.� x��dNO��y�)d_֝P���`�\刡`ҳ�y�O\n��
�_�<i�5�y����!�t��&/A !v��IE$�&�y2 	[��e���Ɠ�������yb��12-�b�N�q0!�HA�y"�Ä?�jyݴ2%�u��*!�d�:���� *ܰ����"�!�$�n"��<wѤ���f!TO!�d�)5Ka:�b�<}�0a"�U�E!���� ���U9IȁH�$Q�Q�!��h�aqpbR�pD�92��e�!��N��ؤJ̰�H�fGp!� �+�$�XÆ��޸pt ąXU!�$����2�P�*�µ���¨>!�D�8�ys�g��9eL��HK�l�!�$A%ٮ���Y(X�Y��G"M!�䊌'`ÕS������Q�!�"��1q��1A�a�r�B�!�� �X�*��4Ӭ������n�\��"O>��`�N<f��t�-������"O�@k�*�q�2�8�,��6��A T"OX��ჴdS 1˞�Gd�Ӥ"O���D$�TYhRj�I5r� r"Oj���`׫X���؀)]K80�$"Op����-�����M2&��"O�u(�dS1djTD���ͭu!���W"O�u@OC���J�R�j8hb"O���ƀC�y�,IbBnN�vr��%"OJep$�0S�"!m�-VX� ӷ"O�,0s�ĶU�@#q�ȰL9�E[�"O~EU�@z���q�ɛ87*F0�"O���C�L� �f!
G�N14��E"O���2��l�
���W�-�LR�"O��{��͵/�
�(&#�$�ъE"ON��n\����Dc�E�<�w"O�ejN =��Q((t0���"Oj=qf�@@�(˵�-6"��X�"Oҥ�&�N)&+�À�������"O��p&',���� F]�c��u8�"O�`�����1� �=�L���"O��H�	����F-R�8�q7"Ol7!�U
�t@!KR8;�pS�"O^�0��("�5� ��5-6RC�"O���u&��/f�M[ǩ�9�H\14"O�:��R9S��&�ܓ/�x�u"O��p�쟑k�z)���
�7@Es�"O*�r�2�6,AbI�9|Q&Ep�"O�Ԑ��0MV�PA+�<1�`$��"OD	i�䌣	V����?�p�8�"O@!U��2A3B��A�λoq���F"Oʭ: ?��mR��˕hmD�"O�X�넪q>���q�A�U�#"O����N�0_�$̑��I�ҕ�c"O��5�W>���#gLP/V�� "O�x�@i��Z `R� �9ZG@uR!"O��6d w��8�7o� t�tY�1"O�AoL�.P���㈜�m˴���"O�I��"�bcgՑ�Ft�"O�ix���
Z��7�E�4� e0b"O�֎ �#�L�Y$F�Z��ñ"Of����+��8��E-���&"O��W�P��:q\���Z�"OLa��a$��1��b�%�"O��X5/[l��8C��-w��-��"O�/��a��L4/�:��S���!�I [d�r���X�:�-Z�V�!��,D�dE�J� oJ�Cv	i�!�Ćt����əgk.��_�!�DΗU�8iS"��'F�J͘Ӏ��K'!�d������I��_?-C S�'!�$?�F��Ǎ��aO
�'�V>U!��ɁX����g6�:����9�!��+�(�aU�ǾL�'�ͬ0�!�ĖW�!Q�i�>}��8q��,�!�����t��g��T��M�bÅ�{4!�d]
���.F%�����"6C!���
fcI��ڸv�u����M=!�D�t�x��3�Y�.����5!!�u�� @V:���,Ay;<��"On�p��K����]�@�J$�_��yr�ˊ%���``�L���8��b��y��FB4.<�`FRj�������y
� �<�r��{vbT�&�7�z�"ON2V�֐U�֨Bb`̏��SP"O�]��B_i�v�bp.Q�i�x""O�Y�a�>3n�����<&N�YP�"OB�۲�T�+�`dz&		��<P� "O:蹲L�}_�飀� X"l0�"O:�	�J��0#��y�f¥#����"O��dL!H&
�E�F�(]9�"OƱ���
��Hu��V(#��{�"O�Չ��P3Hp<��@�n��ؘ�"O�hDCز~v�<bjӓ^��d��"O��s�a̮KiP�RI�$k�b�H�"O�h�GR���]��	�b"OZ}���S��(s�J�"��i "O�Eᓈ[*�ʘX4(ޟ}�(��P"O������3�bm(�g�����"Ol��N�M���V�̍r��"O^���j 1�x afS+QT�}�v"O�uq ��b���#����x&�0p�"O\�9R.�3'D��j��$=i�"Oz�*��*M ��3j�4t@ܸ�D"O"���GI�">�ćX�v�2$��"O<]���g�.�6G[�r2a��"O��r m�>B�+�g�+Y�h�"O
<���ǨGJR<���'E�|Y�"O*�P��[\�`���^���A�"OP�k��L�p��y��Y���r�"O�apD���xiN��떦_�z�P5"O���a�¯xЬ�鏼�U�E"O��Hk�m��I�@Gԓf�ԥ:�"O��b�֟-������$��"O��"/�=x/v5�o�5o�����"O�S�"�(��qh���)Ȧ� "OV��&o�k6������}����d"O�I�H�<F����U!���"O��h��ա+w���dK׫�v���"O�Q�q%бr�H�%+�P��trQ"O�e�tj��.��@D�S6m��BQ"O�p"���+*^<�bh�Mΐ��F"O������vN�)&hޔ@�.%*�"O@�b +�8Sd���"�2�C "O��5I
$\�Ha��/[V��i�"Oݓ4��-�X�9�CZ�X�~���"O�d�@��z��U(�Dy��ye"O�}�^<6 ��B���gpp���"O�J��20���ir�4iY�����~��s��F�&&�9�E
Tp�!��Dkm�+P-L�n�Q7	�H�І�}�Y�V%�|�R�ǧ>U�A�ȓ)�ڕ��,c�ar�/�4لȓ0�D�D��+*�X�y�FЍ0X݄�>V����:��퐄*�%@W�<��3�\�z���O�J�!� �%��qҠ�MˉPlI��L�'�ȓ0��1UP*!��A!�?/:���%��	��*���8&+����h��B`.����G���1)�y�����&�j�% ��ՙ��5R2�p�ȓZԎ%�g�!�y�5*/ \U��v��z����B2��b��;_F��ȓl_���+�+f����")�Q�ȓF�JH����T�v��#�>�@L���<�cAbJ�i�z���m֮fK(8�ȓx|}���L=l�d)]`� ��S�? �t���Q�vtIѶd�I�I��"O��� L�꼃".���p�"O�8ȁhيD<�U�d�D�j�TP�"Oh�rhW�#R� �'�=qL�t��"O a��rcNU��H.���"OX(aA�� ��0���S�0~���"OhVJ��(P���!`F%����4"O�L����u����������Ԝ�@*T�)�'C��A��ǁ$6�����n�1i���ȓ"�^�چ�R9j+�8s�b��H��|�ȓ{��Y5�&db����kș����ȓ:����!��&X��B�)X����%;T@>��B�\�F�ȓm��ܨ��
��ȫ�݁"	"q�ȓ4K\d2%^|Ȥ+c�OA
���l����Q&2Ga���D�� �ȓ�5ꒂH"A�S��R�`�$��}C�����3{�ĩ�7@�(����r�'u�ֆ.B��|2uH^�wcv!�'��2f��	��f)1y��j��O6��'VAZ�� ��*} D"O:��V�ðO�y	���H�nM����?|O��Kf��
>���Ь,T�T2��IFx��8w.���da�Bi/+Ӳ|�`c-D��%��)^��C$�Q�!��ajSE.�O��5���`M��Df0���ϝ�D��u���J�';|u�e�H :|���$ߕc��
�'�����Je8	�)`@�E�	�'PYꕉQ+;ܜ�9���&\70��}B^��F��c��^��y�c��r���0���6X����'�@a֎�=*�t���=^�@|3�'�ў�>	�g8O\�Cr��|y($8�$E_�R��&"O��ˤb��بƣ�%WF��W������WL��`����>Y~�� �K���$?!��V����J�D�0�n�S,E�<��M�%x�4D�AF�1b��]
��K�Ą]���t���3���.n��Ƨ���t��C�<�I�����vQ4]�a	GG|q򥊓&a�4�"a!<O: �����xK�-K�US��3
O~��R��!Z�,�w�S�bn����.]��O�'�Q>�TC��٦5�qZ-N`��Va1O�eӌ�#Z�>��QJX.��4�t�%+K!�( fXa�d喵,���"�^4VF�'b>��=	��I�(E��L���"-# �q�,Y�E!�W�D�VIq�D�jJ<q��]	�!���c����&��ָ��T0"�!��3.�t1����J�B���KܶO"�&�Ӻ���s�dp���B�G����+
&a{B�<�I�R��B`B%�4�0r)��%#B�I<0�H��a��h>��T�<s�"?��	ٻWg6��(A+n&��\�@��4O�c�Є�xy^}'AMU��!�`��\4JC� F�q��W�Z`����U�pC�I�:�tB�=�J�L�3Q�B�I�Y=��"�X�������=��B�� �V]"a�]K�xX"��$�B����m�q�;]�̚�Ӣr+C�I��9AN4#^�y&����<C�	f��SN�-*V ��� �2C�ɨD���o��"�
�H�C�I�� p��³D<Ri��A'@��⟠E{J?��� 00(�AWMS&
��bgC6D��I4+g�$�0:ّ��xg�������Sg��{
r��r�I6i�*�n�8=��IVy�L7��� ���sɘ'~O��gnH� �0�"O���G5�4x�Ǜ%2�R��Q"O�A���ɽn�)��4��i�"O|���(��b�v+d�B�+"�Ɇ�hO��C�sd���4����oY;�!���3#Cr=�u�Qfet|YQO��vl!��S�;���R,1eZ辉Pq"O����� �`q�TQ�ե(Ŧ���"Ob蓧d/}�	�`��-Y�R�:eQ�|�	�qO��<9�hJ�
�d ሒ-|��8CX�<)oBzN�s��+�<�ÁS�'Nў��Z�i��L'1�~� w��=<��Ԅȓl��%�fd�W��8uo�:���ȓE�pP#�iQ `�:���nN9"��F|��ӛI����Qm�K�^�j���i{��IT��P���ػh�ԘP�b�6f@̨ 6D��˕#��wD� �U惣V����5D�$K� &ɒ=�D��}��s��h�4�'��' �	H�i���Y5$��X�!��$���c��"D��{�d�>'vT���M�I�$�֥�������E�fE���&s*^�У�#���?a��IL+[��j�	ɐ����R!�$iO.D�q�V+��7��8����c���l��kZ)� KV>�~�i&��!� C�I�W�Bh���F�&�fX�]��4"<ɍ��?Ej�`ǯ4PJ2tB��78�5�%4D��	Y�oF���F*S@N�� �)�<��哛!f80S
A%���#[��B�(G��h��ز$T�|���� v���Y�IVx�l+�I-3�m�$M�??�8����+�O�r��P�v
X���q`���N��ȓO2���"E�/$���G'�Q�^�mE�������yR-L�#�<��W��=w�eAa�yrON�{R,\X��JG�vd+4'Ђ��D"�S��ͪ�\9?�f�a�m\x� Y�"O�@j���p/���5̐?P��=��i�P���IG�� �S�̴���lH�r�F"=YN<���-��Y�h�@�o.xL�PbW/��Z�*B�$�ͳЪǗ	���z�c�=1����?�	�B��y"���"�� ��	i�B�(Z��B�J�9f~p03��^��B��15�,���
4'��H�>��B�I:J	�a�nCV��R�*G�02�Ol��$��'+�u����22�%	B(�t�!�Նh�^��l��Y�ظ�IFR�!�x����ؘL��80�hKA����'��O?7	>-m�R��^6���&�M�V�!�Ϯ�������{yPyJƦ�*�!�dʡD�y�t���<��S�ʎMa|R�|�h�2W~��Ȍ�;�
��cO������p>)%ۭaJ|AD)�THr�j���1�OV���gQ;<ul,���2{�c�"O^y���=y�9��E�V�Z�E�xbS�$'�b?��n�_�P��,A�]�0m�6$D�l¦��&Gd�`��+L8I���"D�I�AB�;��K7!ʩ_����%h2��p<�AJ�3-�m�G
��Z�.����x��P�)w��JLjE�C�
�y��
��Ļ2�@˪���熛�x��'�$	S�
�78{̸���H(G@��B����>A��$̘41�j�:� ��Z%����y�l?�|�����%�0�x�N�yr�9�h4���?�T���א��'�ўD�'S@�B��ߒV���Cl�5~0h
��� �<��f(/�9&'�
����G�Iox�d7@#��xC�@�Bf���c'D��Q��T�<̈́�h��_y�e�$�#D�X�a)�9>$r]ru�IoP�)���5D�L�@̣,4^�a�LF�+m�ca3D��3���	-h� [u�E
ʐ-��l1D���g/A).�����'z�����.D�0zQd�'=� ���@�8>�����1D��tk�o.HcĬ8thf���A.D���D�I�XVC�"��)��o+D�(jFJʗ!�D���͖�f�d�)D���!�Y,p+\�W͒�$��k)D����Ѣl+�@����J�{DM(D�,H�n�@����˺.�%���&D�"-�� ?Z@�Wh�c��pH��1D�l�M��h��6sɫ$@#D��[G
Y�b,�h�r���^޼�tk>D�,
�g�;yX)��OJQ����1D�@�+�Ġ#��҇��
�0D�t%�H�6��\���3C̩c#D�,@�hֵd�|��֎]�pp�eHE?D��cPoի2={d���@ Lm	�(*D��а%V�d�*5�a�p�I;�/+D��j&jOl�r�J�,��g�(D���g�W.0U�����3��@���1D�\СNðr�ޠ��Vek�|!�k/D�D���^��ʵ�E�̼�'�?D�8��F�*Q8�k��M{XS� <D��)��H�N/9�ʓP��)�U�:D�8!������IqP�Ǘ|Ct��W�8D���/�g�p���8m��@Q�8D�(���o�z`X��C%4|��9!7D�l����ma�1���
M���n5D�\���8
�QѦb��nйwL!D�蛃N��l2!���Q��8Sg�4D�D����`�N�B$�Ͻ?���z�L7D��H�
�`��E�E�Y�wҜR�!"D������q��<Z��Z|x��"D����$��]�p�m��`�Z��u(+D���) �
P�#��D�5�qL-�O��@V��#I$iyHQk�4<c�*/_z�sq"O�) �A8?q$��3�ݞVz�I"O�p�f8X:��FH�"v"O�X��l���JH�I=��	��"O A��KT�{qP�Q��;|a�z�"O��REbP7'�� �a\Ba�4�1"O�ݢ�C	\9��"�Nto(���"O@\ ��B)�h�c4���6U���"ON�ѥ�7-�|D2P(D�Jn�1�"O�[��ݪt���a�A��;8�y[�"OjS�M�MHaP� W�-�x��"O����p_?8$H)�G�
pν�ȓ�P	j�ĉ�fF)ۢe�%M�nȇȓ`����"޲(��XCt�Ŝ"�Y�ȓ,OI��&�/=|��r�M�3A~�ȓ�}�æ+S��� b�3i�=�ȓS�x�1�L�1������*<�L��e4��ө7b��i�I�N�4��Ku�A�S)3	���k>���wL�R�J�-R,�� �lW��`h��1BZ�6}�hD����~��Q��&��I3��3Q1�L`�Ȥ]�q��E�����&B���S�O�	C`��.J녁оFT4�p�'w��Xf�Ǵb Y5@�8��5�-OTp�1�(x�;�H6O� �1xP+	#����ǌ"C��6�'D�X1���
`�AW�I��rN�;��c��v��t��I-2�Q����n"�}ᓀ� -S �<�e@�/ <�i�Dl&�u�K|
���,��3��N,? H�x&�t�<��,e�H+i
%f��|���1/#��b�̀�V��p"�JφȎG��'��I ׆	�/�D����B��&��'	���*Q�I	�8R�+wSj�0� H;������!@D��"��׊a	��G}�`T�C���b�E�5���BP�+ڨODA)�H��(gX�CsJ�)���E UFS>���UH�:��A=y|ȕ�ZMX���I�Xb�`���2	�,@$��=�4�VWS��2�`H" @����C�zSx��%[�7�8`�?���B$1�|h��e%��unU}�<��☨P���a�n�~80�BA�4o,��Ju)���w��.��U�O��h��D��z�8�O�(+`�R)e�,�Y%�N����b��h�a��6��'_D�d�%�ـy�te�`LѮ�uz��)Y���������z ��&�~t��;_\��h��p��<�CX�f�(�$�.:�`��
J�1�'�f�)�
K�{9�)ZFIDHf��M��w���B�X�.���g�bU�5���,���R�?�I�^[�CgJ�'(�����E�Rf�&%+��;2�;����F޴+`�I�>'K��c�^�%c�u��&$ !��/@����y(�" V�)�#4Z-y�*Q�~����Nt�����W��D���D���y�h��/e&�;�d�\��y�Jʚ@�l1�r�ED���k>�a���1+o0�c$D_��YYt��AĜ�B"LYD|Q�i�M��8t��`�b"K�I3ȕ(r��`���-�,�`���>�A6���J%�G铟f�d�XT�,au��j,Ց{�&�9��F`�fg�+�T��)�<a$Ƒ�c|���r�� ����#��e���.Mj(x�L����Ϡ���q dUȈS���Q��ŭ+Ed<�!ۊ#�����3]e��� �)C��(�
�IT�-�FX:�?9��{љ�ń&-���C}�֝�����m��иU�\&�<��SÒHE-���Ϗ^]�� ��Қ>��4�D��o��ذ͟�N�'=����Z�H����)�%l԰yn�s_Phs��y,ݩ����TN�iD.IJ�O�?��]ϻpc4)�ȄHĦ���Lwl,uK���Ҟt��,�N���1���|:���Lξ���h�pl0IK��A#Pt�y��ek���!�|$��nZ.0�qЖ�P80eJs/��_N���^�����ͿId�r+�"[6yS�'�^��Qm�+�,��S6auFP���о��!jR�%W.MC�'E_
��1mK��"�IR�(��U���i���Gh�'� �hX7Nl%�'�R ���� d���Z�|��1cID�KE�4����0�1
ԯu_�����o$���HkڰZ5\�ŇI8 �X�P��w�ܟ H��&b����>-l
��L��WJ�r��>k�@�R��N��u"1%��"a4��fi�?/h$?�ݻszI�XY���ҒU���P��34��ԑ��]�R�$1�%��?C��]R�-yeK�]���
`ĔD�-7Ct��eI3 �m�P��B���R��X��(30��?:�GV�%�r��$G��dx�&�A� �0��А�:�0�Ů*��I�=	 -�7�J��b�E��l����%��3�ҕ�#��O����r�[�]�`�gX�<�Mⴊ�,s���e�6u����-��H�������U�P���Y�9������M��%�􈗁6W�,Р$Z�y��A´j:�d�4�������5E��"����L�!���k�[�@��
¿� ��t�[+K���ňU>6�6�ې�C-Jݢ��T���]�T�Cê?���weL��OE7zӆ4��i����(�Px��AL�DA	kdN���)ʥQ�N)����?P� !4��h�ir%���
�f�+��P�A��qʶ��L!��.G>T�	I�i[&m��\�'����OZ;{���pa����6w�x�"�i�u!QaB����'d�N��|���#n�Dbv�.*����$'�	bL�`�J��,K�H�Q�L!!D�=b����ʃemI(�A&7�,��P�ʈ"�̑���^. [3CH�8
8��x��I48qpB�$�Rұ��#Lf��4#��p?�R`�=�� �'��	c�LL�͆,����"��h�H���rаڴXqx�Y�o1���"cZ�y�͘�QbfX�p/ۭY�v�8]@0���[r��"쑃=��E#�HKN"]����/�1���شR����d![z�����8��ecU�
K4i��p>�����0��Ί�"1�Q��I�n�ǥC�:����H��#�C�w���,F_t����	�28(.T��g�E�t���͏L�%G{�K�`��!�4'�?�֠��.��'�д���̬"��YV�#Ktb���(L=����Qf��x���]�tS��� M Q	A�%|��ak�,�O����I�@�X�G	
��"@��:L�@j�Ġ~��tK��6V3����d$G�@ ��)�� H3�3�B�;r�y���P��U!`���1�"O���˔�n#��읜L����oI(Y�L��F��m���$������u�<k.�5��\N��1��Q�%��)^�`�UL��H�ԙ�Bn]5Y�~��%�K�YǠ-��l�9)��U�����FM�`��mq7���S:�kc��.4��� MN ?�����13N2�"��
��(�c��p�8�D�m�'#���a������ˋ_V��"�)�l��
،ؼ�ȥ!�>)�)�����A-�	[\��_�-�L�AÂ�;<�|� ��``J���lŚ1&�`��/�~�`()�2�L�A�I�8u!aݾE�e`ح_����A
U8��-[�Y����A܎K�lZ8ͪ]�&�A�Y�(��Q�Ɂ{>qȑn��*���H�iH⬴)I>A�	�J䢨���Б���6�؜�DnJy<yؑ,�$L5��*]�{)XTJ��޹��u�q��8����w�ĦB�𭛀l� F-����y-^Db�韻��7M�0J��\�d犟}���$Eخ0=)�J�7N~�ؙ�/�)NW��z#CP1I��T�$G����T��.1>�T��}q�!�e		A�j14�A
=�H4��g^\��0T�BK���hĂyy�<��'��kZ��ab�\��80RE�9ZS�D��U)JM��΀%X������aL���TZ����Z:[_�|{P�#d8�Ԡ0��x��9nJ�-:qᆂI��<�� �1
�
��b	;hA�Z�� ��#Sώ6�J���B">�ۇ�=5��L����Z�|Q34b��[��4�T5��+״@$.��
<6��(��I�Ҩ��ꐇ>�v݂Ēx�O��ub���)D�#_ �
� �0�F1� ��^�VtyR��,[��Xr"�E[ у�Q��\ɪݴJP�q�ˤ{sf9�5B\*]�J�;1����S�]!��	:j���C$T��x� 	̷xOn�ˆ���8KXu�q �$	��Xۇ9o�����6�P���̷zFz�N�L-��-�0\��ધ�5n4��t˕0(� ��+�/xI�P��f�Y�'�Zi�b��k~�J�3k1��+��)H�����"�j�|
�H�B��|���z���qÀ+di��iʤ�$:CP^R`Y2��'>�-x���"'���꤄�h_()a(��f�� 1$���{x�8р�W�^�*)��Gj�a�@��L5I%ĩa���D�6sl�P! �R�P$P0ؐ"r�E��ΎLL"�bA/0�����d�e�ߢ �)K�1�p��1��Y$�b�`��x�P5��%��!�j4[�ś�Qի���貭@�m4��(h��V
X+��v�9�	*j,f��ҨW���;���=ҁ�Fb)�be���8p�������i*n��R��'��sghX�>��N
C2����ٱ_f)BC��b����P$+< �1�`W 7�����r;ʝ��&� JO\吰ף��	���i�1�tD�
[jbA`r>�����"NEJ��شA-D#�G8a�H�[
��
��'-��h���IQPɻ�)�6b�9��B݉.�}��Qc�1 ��#���r)P�[��IQ�sx�̓(�y�u�O�3��ŉSDd�T���6^��ԅ�	�@4J��@nqON(
�)N!4\`�9P�E�-��E�$��"P��zc%G��ə�!ڂ/��L �ჷ9��3�l}�2H'�8�N�vu�y��`�,qO`�1� X#jN�}��%�&exvl�7#�"�)��d�|Z�hR�GG&}0b୻`��)I�!7�����I�̼�w��ZcrX���]�1���%P}�~��e�Ǵ\�		�(Y�S ���<��:�bX2Ҍ!���yV2���ՠv�������	��yӀ ��xT6�!`�*Y�:)�E�:TGfH0(����%���p=�$�C��f�tbB6����eb|�A�� -2@��Ȁ<_�7m.b7&����Dl>��c�1��&Â�]�B�8ز��a�������a�)��}�!O�(�&���͊?V�a��C?�α���.���`T2�"X�/��{�N�2��:N�1�=�̵��mD/��A�W����D�K�b��58��:yّ������*{eFP�t�3i� �����=m����,E&�V�9rc�=X�8�c���g�T�0rjD 1Nգ�o�9BtNA��E	��O��;F�@=A�P�{��=��Yy��O�bG�#4��?�Q�Iܖaf��v��=C�^�3��9��MQ�=gN���b�o��l�D'O0J���S$�%�����-�OJH��L��	� ;��O�7|hu�VŇK�=���35g��j�7mAZPؤLP� +���(1wz]��4�%,Ž!�h�j�f��cc���'�hf{�l����,d������F����a�&�rs,��[.6-��gH(�A�l��S`��kRo���a!V$C�1�fe5F�O��bো�&jX+P�K�A��)hV�ɺ��De�N�d;Z�����a�p�Pl�U	��"�A��d򕫂�)�
%��J�z(n�yM$Z�2����X���ׂF\�'�!:3mJ�]�6�Kl
Լ�2�`Z#0۲X��B<�� �mJ�%�c
6^�"�#���ܨ�J@� 5(ݨ2"�8=��mj�G����I�v!�/+��˓�'�����_�1�*��Կr����$)�x��Q3��4H�7(��N�����4Ko�Q�qfêz�	C9�8��,� 6�
]J�Nq�fuV�' ~�3���2TC�TV���F���`1hE�G�NST� ̈́
3��$a�Wvr
���E���\�`��c4nQ!W�H^�h�%4�L�JUmߓPFfd�FGո�O�2�)�Ncz� %꛼#���`�Ϩu�}�􆁯6�XLh��1��#2lU���3h��0uN1cѨγ'�Fuip� �0��PyU���ؙ�'�3r�v�d&O�V�d%p�	�,t�cnֳKl�t9%
�����R���t�b�	(U�8E��ѻW56`�5�
7̞Q�e�)D�kE�'SR�ѝE��ɒ�3X�aC�� �%�
�9��/ar�!Å5#Y @��ПB����FV�7P�y{�w�NRF����aH�� +'Lə	�L���E�7��}��b��~�PP Co����5ƴ[ �I���U*ĩf�XJtd땂\}��t �@k�����O"�Jb -jxU�4oL,2v�(x� �iܓ;m�` i��bEàK��}kr��sf@��\❏-�����<y��yȔ̆�B'�٨PY	Y���7j�O�j@"��$��n�{� Y! ��R��Z'5h>��Ӎ�6��2��wn�Q#���<�r�s �"��j�fZ%0c$��c��5��}:���jB\�:���)�҄�o\g�'.Ѐvd-apP�bZ�8�A�Z1�Z� ��W�y@⣌ ��%���Z��A%݄#<����۳�V���R�YB�m��I�/�s 
5���2!N�"�<!�$�8Ƙ 5L��%u"}����-(?�1�F'
�r�q��]�5lj4�"#�"r�`h�������cf,5�zǮǥ�h�)1��1dd�	�' ��)��:��8R�mH5l(ȀBb���~r���nD�A�6��"�ǟOJ����6gDan�l�Z$a�"�N=��	�$>g�I���b%
���T&U�#&_�hڱOKR?
֤�*�'Qc�M1a��hAh��O�Wv�p�]��T�Ѷd>t��ӏa�qq�JE�kHx�s!��R~%�+Ť_ܶa��)�&�Pzd�3b�^X��-[f�\,&ϥM�1I�#"�\bt(3c�X��4C��xb| k"b�`�� �
�J:"��G�N�rT�٢,,@����	6��qi�E�����/p<���)B�|���㆙�0�ʀp񅝀��D^�5�l�鄦�*� �$a�>s���Y�lW�JgB��	E�Iy0H�
�^mr�C�#�ܖ-{��h�$��x�*��N�Jj����E@@p�w�S�p�,�4�@-��l�[�|��'ꆕ]X̴�A(̿pKN�*W�{�hH��E����{gd�?�5
/)m�� Ħ�:&��rUK@�WH���Ϛ4dX�fÏ�6y��@E?j��e���ԣm<��03�QB��<!���[X��?V�)�+Avj�B�pG��Z珂�E�������GE>Hp���(u�<L	�
.Et�;	�	�ªܽ��qSMC1nIqẻ�jhX�Ia�_�@�$�H!�6�	4A�(� �×�R̎x�����a[$G:��xr�Ƅ/�6��MO�}z�����ud\�B��S����qA�����@&�,�&�!эxp��� 0�k0�ˇWR�U`E�f ��5P����
P�"S��Y-��!(`�B)
��b0� �R�� "Ā���� @�*0�E*H�@8�dr M:|f�0Hj��_��DhT#ʧ"���K A�"$�5ʈ�C=�h2�i��э@�r�4���!ɥy/�U9D`�� �	�8|�h���F�Ӧt�<<�T�D>/��&�e��,���ىt�r�{�m��1Sh�y�#Y���(�n;3� ,A����d��4�=��#M�^KVt �BՅ�n��6�Ug@�RRd�P(^M`p�o+L��$A) MZ`����l���b��eF�RB��U�ʍ��gۡ=c�M�"�@��x��]:+v�	�[�b���hsV�\�@b�;�J�*'n�=;Q�P g�FU����N�..I>�ۣ7wb�qtň��������9R��}K|uaB
»8��Ӧˢ�t�5�l$�2(�� �F�'j��P���C�Ҥ�ٕ}�zm��ُ`\ɘ)������\�z�X���V�`s����n���GJՈ9d�I�V�V��#}�w��9��96[�D",�:b���+�Kq�Pt��I���,��M�~*fi���y��I�P�����ߙN����K�H>�l�!��i����`�]� ��ψO�q �m�4c��4cV�[�����q���ٳ؄Ƞ�̟���s��a�Y�t��y���=h�)F�� N��q�`�*m~،�����=Y��3r���O;�@���P'>��P֏�+���{�/$��V�*���s�ı~)
q&?�م��b��낦Ѭ.�Q���(���+�G�6�`}�O?!Р�0��v��$9�~��C'D��0�>d��Ha�6�3�j�<�I�P�
���,}��	�4'��ؐJ�K0����@	Dr!�d�q�>h�5B0��tÖ�I�qO�e[�d�
�0<Y��T�C.���'
��S& Rp�<q�n��c��E�6���?��L#R*�r�<��/Gvs6����y�)�J�m�<���ՅdAV�����6$.8+D��d�<90
�q�LВb��:�E�f�c�<�-O�T��.��=/2���#t�<�B`�!��	EA�VF�+�#p�<��h��!���p��S�))(�vG]m�<yS��3J�|��eS�FE�T �@�S�<pL�eF*0�+2G~
��㧅I�<���	�EP8���T�]�LACE �J�<醇=2"~�0�)��P�a;���^�<)TK�-O�v��$Ϊe�����Y�<y�50��ȩ�铩\��&b�P�<�Wj�h��<����'1$�����g�<Q���NRbi��4ɂ�Q�a�T�<��ձ.�-[Tc�|ih)qPK�I�<���,#�̰`%ώn_�bd��@�<CO��Gz��W�ӉY��@�1�F�<�de@(?�`��!��_֕	�C�A�<ArkI�*YH��r�K0II� '�t�<1��Y�yvE�����T��~�<AB+�k�~p�!�>�RL)�L�s�<٠�A���Y0��2O�ݳw͝h�<�'�ZqX@�!/��L����gMk�<��Z@,�
f����2 �x�<�'�V<I
p�RR�V�j��T#�O�u�<�$�W��r���F@��Y��v�<y3��;M$�[�LF�}Vty��Bn�<y�%9g��	�$�*3vP�L�<Ar�E�(��U��J���X�I�<�â2��4!pf��V��t��k�@�<I0�C�/�̉᧨����)FB�U�<)�R%i�݈a�	���{&?D��"`�p���s)�6@�X�4�<D�����L={�>��3̈��lD�B�8D��a
Rr�h��7j$,�� �6D���	�xxD� t��?���2�2D�t��j�@\9V`��J���huM:D���A`X�;d5��+J�f��܋T";D���$Gj��1X�a��Q#�KRG$D�3!��-w4(jҫ��-}8q��+"D�<ÂB]�74�00�F*��e�7D����V�D��r� TT!,�9�&5D�J"�>���R�ԗ�{�A6D�� 4`Z�'��%H>w\���"OΈ�eI[�u���R'�	Jn�x��O��ˤ�: Nr�O�>����<����"՟m�V�b�)'D��Q#i
*�fp����G>|�2®<��!ʶOK�(�	K��0<��' y��P�@�i�b1�/cX��r 
�D:i�k�s��d(���5�r�"'Dӻ%���+�';�9BG�J
k���>G����ߟo?�2�9L s��;��ra�J�7;��c�L��Cg!�ěM����!e�yPf��7mȼAɔ�Z-Z69Їe׾Z��򧈟�� h"��q%a�):���tD�?�y�\��K�0/����HH'{���`$�~(��BO�)��\�G���|F|�B0GL]���,1��XB��*��O( c�����y��$7������C�B�64�Bb��`ࢱ�X�#3���OB�)!0���oXt9�� +ClL���G�D��ŗ����F��M[S#^	;�<���BP3\�İ4�3b��Z�M��p��͞����I�!�yBI�u����%����Bá�� V��b�ΊX^ɘQ� �5�5��N�����lp��p����ㆫ��}ȃ,W5
�$�"#�ɚD� ��)��G8L|0I��F�ΤrgÖ�4Ḵ�� ǧD�Qc�4T�j̊f�P�А��I�i���Ex"m�?3��X�Ƚ<5�<�%g�V�5�!��Dӎ�'�<�alY @۞��#�΢Zp�V�M���H�!l�x5�M��39"����W-O_(�P��VBڢm�?!b([5ObxPZe'�/��)/�N�Y�%Q�k����\�\����O�qQ͸ F؟o��ٕ��(+�Z�	'e�
l���џ�O�k�����6S���LZ��V�|����-L	m�h�
�'EЖ��7-� r��}1�CJ�c�$�Z$�~��0"��q0��b��|��!v��QQw�g�,�B$-I�#�����%�Bh�ЄɈ�<���b
�z?Qs�ON,řE%����'�8-��'�RK^ag�֡{c�I`�R/h���o��x�b	��Q�$�فbֻ8�����KV�{b�IR�y��{�p-����> �����V%
��	�pg^/E%��C"o	a��Ix��`�H?#t�A��B�qC2й���1����paD�I�lɒ�J�i���`��F��$l֭�d�ƇJ�����	M�z��@j �jz��i�Q�Ė0U�"���+�yC�]9bLC� KjkhS�~���ʷ��"ěd	�`�I
7��_��s��0�*�qҢ���I]�Y�,�GK���M� �Z5X$��k�b�j7=��A�BJ�v.h�S�l��y'EO�2��x��Q�!���"*X�)Pb���MbB!N�*�����O��l9@�P$'三�*,Z�k�P5&`EQ�F��'�2A w��M���,(�丂��$���#/٠i<J�w�2����?b���`5 �,�>Qb�	�U%�K@4R��rH>A5�E�Q��"���%�Dye�1V^\c��\�x� ��^�%�H�0�4�`�2@�t��9�(O~����A�=�M�wlÈ'�>���c��zΎ-	ŉ_�5˴����	��x��Wl�V��q��H��[�[���Do�d[��w��x6Hp�"XkLH�|z�o_ e��EQ�k÷R�~��4�������[����%�]>o�̤�f�0<��ŉE��
Y�����(��ksT=��/�����U�ܼj�֐򶧕28���ɣ ���05���n�8���ɶh���D�k�BU3G�N4+K�I��yb��(C�y�D��]F�IY"�N��Bq�eN&p� �`�D[� �����^�@@B�ÎeJ�iJ�����]�̚d�b�J�M$tY��ʌ	��10׮�h��������j��В�@���@���w�R��F��I�d ���v�������CH�a���
Q�x�Lΐ
�>E"�<8q�dl����Y_$0`�I&�j}�Dg&y�N%�E�� 熬0�,�N~|\�lԢ_T0 Ү�����w49Ku�A9Q�> �֮�e�����T%���o��ҧ��R]+F� ),l���7F����̜6d\ �q"Å:���r3d��\����� -&p�s͍.2K���%�O�����X�:�Q�뒯Xf���>��W%^� b��}{�*��͎�0�<
f�:Ov&�1N�W(dk��
#g�����'��@��!C�cT�$j��I�!6�p ���6R���"ޏ>���c!oU����A�N�ƈ�A�׿�n�a�E���F�:�NR!jb�^�r�h����7GF���	�  :w �?4�Ź�װ_�bM�P�w�A��#^{f9���W��MԎ�)uzȻ#AN/a�ɺ�wD�ɰ�)ʴ/�d�S�ٙe��+�'{�=�sjK� 6�8S��Nb	�vg =��\PK34K�E���2j{�-�j
�<�#$��Kv%���'��z�77�,��b�,rw��BӓQ@pqEO׻=�f���Ա=��IsJ�-ӛu�X;b���AҸ$gX��"�Z:K��&��s,�SR퉂t�T-#�i�?W3���%��3�Db���Aŋ�6�^ 	԰a�H�3�#,X�cE r�N}(��o�ִ@�I�E��L �f�����͋��>�u	��bX���$��Bg��`c�P_�،QV�YIx�i��
1N��	�dU�%DFo��hCD�߼���G���D���A ;�H��X�<!�
1�V�3f���& ا �%_���
�9cJ��h�|�P)%�	5�@0����,<�kA#R���*l+�@� ������#K��Җ 
	�b�B��������)��T:5�G��,N��k�Z,�����a�a1����#���
�)мWg.�P� �e�r�R�	�.��Gz)�$ٲ��%
��iV��X�I�6I:���^�fԂFŐ/|.����$L,�}+�+U_ݰ$�u/D1�0��st�M9g�OQ~ȋ�Ϟ;?Y�Z�g�y��4�I�(<��Ҽu{�d䎏�.%�q!��ٲa�0i�ǎ�7k�T$adB�ք�7~�T�n�@(�e9شc̎A���l�ȥP�D�/ X=!&D:Stf%:U ^�-�$��В|B`��/�(���b�aE(�5��Q ���B�B�	.\91d�ɲ�� �]���Co�
2��� L�?"��!��;7���@3A�ʺ��p"����#�؈6��m:� ��Y�G�9h�d���ȼT� T�A��at��N�����{�oC&W�i�'�i�n�@H�=V�,P�!dx6+$'ȄS���F�H"b�¨ �JðDy�lx�Icp�<F+��:k�')�Fx2,+�	�%H�`&�1xLIx��14�0�1�AEqn�-�!�f <4iҝ!T� ���OPqhv�3������p�"���M,z�>�;��@��
��c�Q��#V)�$dt�[7��2aTx��ͽy��;3+ ������T(���.��6��E �
.l1�>~��<KëY�!����f�P ��Ӈ�� '�T�G�ɴ	:8����$�ēh~lx���,O��{4�X ��ٖ!FE]*�ڔ�K�BFz�+��͏zz~��b]�S�ԈĎ�����/�F�sA
\���ъ�*����R1?���A�OᡄI�/+���b�lߨ�,P�M���*ab,'N�f�KL�����."��z"�iڨ���w��݉�J��~,`T��@�Ff~�S�
��K��bǧX]xt�8�£>�Djޭz��i���-�zS��%������ta����^�,�7�1Fa����/J;Ǜ�g	�j�36Kȑ^�f	�BcC`�i8�H!��<6%F� ɖ���PD_r%Ybk�&"��U;
�ldB䧈
��=���C_Τ�� ƦC|��0�\�'8����'�fxD'ɍ������H���z%�<5�,�Hs'R0H'�'k�Ib���e�Z�S��4�*�ϕ�6�>��S�K"��ɔ��H�2p�� �-ұ�V�7YAynڇ�PA��O��V+��J�LI�P�ɀ'Zb���R��O5ޅ���{�ܠ�!$Ũ,퐡��c\�%��Wk͈LL��2�x9�an��E �ۥƅ�".,0z�j��vȗ aElZ0������h�j!X��'R�y�($h4�L���� w�̵� ˋ('�Q�fK~��)27	܊����q�_�j1�P�׌�"r�¡l�W<J��d�D��9�G_=<�����e�4������$�۱C��'��OPF����B;~�$��п)E���$���G�� k�MRD���'P�h�����t��!�X��@�A��$.ކ$(r�҈��'B�`�D
K��rt�"y�D�
�B�� �-{�J8j��^��rQ�#�|����7�i�~O�-Z�^5��B�)ܸ'n�� � O�tBf-��UH�ˊ �MȄ�G�f��hSeA�1o��]�}4i��Y4;�\MX l�����Ɠm̢��2b�%C���:�h,�
�-'�U:���! _���dRɒ�rK	77���R�H�I�ZN��A%���]�dx�é�?�Ŵi�����	Jry8����ebF�1\vL4
'I��i�0��kf��L /Ś0Nn��*�;G����7e1�����,�!���K��_�yR�6Ɠ}��A�>v���Sq��!c0y��G�ywm��f֤�AL��4>�v����>	V�Q�=�@�Z��!LM�����R��:@!/!�&(�T�ɋ�,I��m� �<�"���IA���Aj�8Xa����y���#������!���z���HO�]X�G�A�B���Qvw|���u~�q��J.y��T� ��`��9h��\g����ˊ_f8毙�r��9@��Kl�'ef0�fL�L��\Z3�K �>�HTFր2k���d�
$6k�4
�O��Amh(�&LN��x
��
"�4�`$f6���r���nx<���h�"��z�/c� ����'af9P�E��,H�զA#`Xu���W T�mؑ���\mL(B��ij%h@%�&@��f �&iLY��w8D��ًctT\S��P�� Gx����6y�D 
3 ]pb�̪Gdb`�$��J��iMȩeH͏j�^d*���j0h�p�]W����V	')�b�+��P立 u`��V�"�O�}ki�8]> c����$X'�_5@�\`��� ��C�U�XͲ��.k�.ts!�C�:�J���J�_��$�F胶>�=9DL@�qp؝2�h�-u"�s��ĢB�XX�眪���
����B�Vb�L�ssҁr@��s/�34N�E�p��&��^h.`J��	)yv�zehA�?`�!��F¦��>qAf׉4��Âɟx�ڈb�L�&ih�8�ʀ�*��б�)fɠa2���ʦ��%��=�f�L���y���L�x�"���#������0>�u��\�n�"4 �<�θz&-J�Rg�./�fe�Ï�+f׬�ɀ�Q�r?XԊZ,͉���o\�L uhл%zY����ܟd��&�J4���#��a��,1,Y�=���8<2�D�'�MD�2��#N�иև�O��H�gǼYh.�ґc�fs&���J�0qf����-1F�Qv�Q�'��T�F	X�V��*�L�c*,:��Ll���;*\�w��z6b@�F��H�&�8U��1B�a������xg����ȝ$ϒd�G9ndܺ'�}�a~�O�90���$��3/�p��q��/���C�!�
L���B.����Q�"/��5ର��0)�dԐ��'�yw/�-g\��d�#�|�aaV8�p>��i�[�>��+�|yB|@c�5�V��HK�S�^�g��!:P�q΄����pE��<~L`xrc�7�B,��苊��D�O����h�uF�����0,6]�=I�%ؖ�$l�d�D�F�����6 T�Y� 郥Nܐl��c۬b�f�'�=���ɴ;0��z6�{��)I�ِ��O�D�C^�$�p�����i"�dω$��Y�
8\\X�V���J���ߒ#�`��u 5j%�J�Ď
"��9i�L�s����"��=T)���`#�l��D}�J�;/W��k�	�7��)x�0��A�7H�L��Ė�2��� nHۄ!H&+�FX��jS�}����6I�@�����$睨k����%Ƃf�r�Sr�ľ^#�˓	��1�	 �p�h�:�'PԚ��g�Ux~�*�����I��h�}��a�'�2}��1q��y�*���nߛSuh�rs'̜��a�W�����0�v��u7��c���7�2Ty����q%�ؚ��ͧxmp���J�P_��IQ� �S���	�5
��q�b��,f�Zl�WJ���@�����(�2����{��Y@	Lt�/GD:�-Q>L��ݳ�!�3F��J�F�	5 ͓�*ٿ~=Ctj �!R~8��3����a���B��R%��9�Ӵ*ɕ�� :$�)AuDݲ�d��@��H!"B��DptF�%jX9�ʗ�&��< �D�G�6�5O�GZ @8�#Lv��9kR^�FA*d��%l8ʴ�˞�&��O�CR0`xrR�N|��a�ӎZ�>Hc���oG2��q�E=����Opq�I� ��1ň��L��@A�6!������?u�`-�c��9�(��9�4TҔጓ$F<XP6�@�c�4�3/�N�4!��Cg��i&( :� x�DAM�!N2Lx޴
,�q��#�-�p�����}5D��`bڶ9t��_�2����Ux¡@�D�F�
t�L<��}8q�:� `L��Vt��T��#S�?�ܺWc�Y�f� 'k�'>5&a���.~?th�e�O�<~t��H��`�q��n,Lb7�8^My�-�%~�99��@$q�p�c���e� q�'��-�]0�Nd��5#���qV��2������-Z��|XR+b-�U1��ܞ`+�qas�M<;�xĊ�(�&��ɩ�%ӇIzU�Rf�q6ع�%/ZV*MX��+mv�Zc*Z�Y���Ffm����t>ԥ�E��S ]�VdP������!^�c�TXr��A}�ߖ�J9k��J�@3bh�E[�M���Գ`/*=�Ot�"��Xg��h6��#8��X�EѮw� �������UH��.۴]a��D�!f�1�#��Y�2���G���%тp���tn�=g��I%-*U5(�!��I�2좓�R�����?I����32���Y�#�!���k$� �A�Ɨ;��X�!]0@����2|X�H^P'�1�%aCT���`mE8h�-�o�/f��;de���[1��z ��� ��6�e�e���%��`>m��A3O^<Zd#�Λ1	D��p�^�Ș@OISp1�ई�T+2�i�}�c�NV׍��L�d�1	E��p�lM4#�Yd Jh���{SOR�1��d�`�јD�ЈF/
�5�*�X�,m݅ �fpɓa���	Ѳb�L�C�jG$)��ǟ)��	֊DJ��O?R%B��f�h���͉&&8���O�Y��1t���D_&�KT.�$L^�T)S��/M�iQ�!1E�>!�;�Ȣg"~�R�/I-�Flxp�i�ȭx#�N#P ��eSɦc?!��)DƼ�У�k�ʷ � V��/�>>Y����[�$B5���"�(��g�'�����!ZW@�P�A��J�aY��~""�;,
8�� �C�9O<`������W�P'��2k��ȒF�F�%�U?Ua{"+۹f�.��v �p���"�L0f.�@�e/h ��1��M�I�h��!���-`� ;H~�d�+]u|@ NN�BU��j�h�'�\劣@C�sw����~�7+�
"�I*ċ�i��r��	A�<1�$�3M�GQ
b�1C�ty"�_�D*��B�Ll��S�z�1��C=(	�9R�kÓV��B�	�L7�e�H�Ղ�`\�r1��DIn�9Xax��ٕ|P0G��U�
��7�G��y�e�8ohmP�ήJQ�ZրY6�yb� 3:��� �=s���9�$���y�-�5.5��7^��jb-Z��y���
��h�#�!X�М��`F�y2ㆄP��I1E�G����'��-�y��M��m �G\�;�x�X�ǒ��y,Z�g���!��Z��в�-��y��0?� �V&eޔu#�,���y�d��	WR��'��X!��(����y�f��o(��*rOW�P��T�$���y�O!M�\�A2f��8�l���	1�y2�<'��h��T2��u�A��y"8�s2�2'��	d�΂�yR��k��h��+̠�À��yr��7��B�W�t4� ���ȝ�y2A�-���3��=�,��pNM��y�NʅK�n��_�8H��� ��y2��8���qw��	�L�k�/A�y���[����doؓ�j}�C-�&�yRDȯb |��m �p[��#Æ��yr)�"MB�a�^#{�h�s��#�y��A Z�P���d܇&y�!{ C���yB�͖b~0��-'蕃�I�y�H_	f�s����X�2I��0?�T�C��t���&A��2����{��R�GܓR[-�Q��w��1R-�1Uq��ٰ�
�	�� .G�a��$J� ��ı�4A��  �D�����$N���т������h

�H�4%R�c"5��Pm!�d�A����:T��KȚ+S�8a�NV�8�Љ#}Ҫ=�%��蝔1���3�*T�@�p�������'��&�)�IƗ2�qe��M���t*ܞ]��'$�LGy��d�B�y�TA3D�T
n�H�t"'��$ڡ�(O�>͢!�ԀLO�D��o�h�����bӦ������J�%+��,	�e�>sR@���^)lP�*��>�v�O�$�k!��U�2�I%��..���@�k�9��USs������0|��DB5�n���)B�5Ub	y�!�{O&�X�8O �RC�����Op>0�֌]]�� E��Q���C#h����ŪQ�P�)�'R�H�P�耮qP�%���E��4(�����O8�a����d��.h��Tz�DΗ>���2�,�zw슖;O�6�R[G�KE�~֧�S�P����KD"��
SDC�A��`�>��@���0|�$���u����~I���bN�~H����'N����3� Z��Ȏ!#r}�3��+Q����O��'�FO��a�S2Lf�����+:��T�T�C�%�t�OZչL<E�4g�%l;Də7f4��Չ��y��v��S�|�a���$}�"5���H������Ҟe.�OpE�ߴKz�c�b>� �$�KJ���h�pe;b�3?�)qӢ�ʍy��)�<k@�ӱ!�K���@�ƾX��$�������56����d]`Þ�$'�>O,R�xL���y
�'��0���2p.���N��: (��
JS?yQ-w��	��?UH�LY���C��?��W$ N��a���y?�)��?,�!�y?J�X�܀ܑ�*D|!�DI+u.�:�	CJ'��*���!�d0s���c��~�x".ϊ�!��F��@ڴ��[�(�B�g!򄍯|�1����
��@��(��W�!� I�>$�V��|��e(Ua���!�D��9:`q���ɯkm�]2� ��^�!�®9����h 26.Ec��BC�!��R�v����,d�f8#��Y� �!�d��>"�Y� $1&V�C��Ճ5�!򤜯
*X۳��#K����Sn^��!���%B�t+��>�Й��l��g�!��S�7�z�ݝF�P=�U�ѩq�!�D>d���	(Ԅ�*&�499!�d�ti�eKɹu�&���YK+!��[,Q�d�g�2@������<m{!�d	,J����#�`�(�,Uo!��'��ňE�_�qe*�������!�d�:M*��T<	�T<0 � �l�!�$>}�	�C��*g�a`#ň�`�!�d�/&��Yba�5w�j(�)H8!!���-��QX�!Q;)��A1� ad!�$Ö`z���j�3���v�Ʊg_!�D�:l
��U�0Gl����^aN!��u�jʖ�R�cX��P O�Ge!���#"�f�����HF$Mz�����!�$ �AG ���S�:�\���3t�!�� �J�`b�ϯ1�.u�Kߓ�!�R�rW`��6 W�{2P@�ˈ�L�!�6K]�V�z<��K
�!��w:��R�DU�W�\(([Q!��	EG�E���	Cܔ�
�A��!��$:���Aճk����c�"!��8Bք\��T�`&/!Y!�D��2��D�c�ZN�� xU�I%�!�$GiC���&��u#��;�"K�8�!�D	�T+,�` ��d�����x!�&4��p�#�	G�`d��nžl�!� *� 
Q	�(<H�%�՛'�!�Dطt[\\(��(K-�������l�!��9���!�ʎLy���ܡ@!�D�'N�0$�?Ll�A
��_)!��y�� ��?*�y8�ǃ0a!�d�"&�ڦJ��\B���C'}�!�d�5ta�gM`*��(C"�hz!�d�6:�´�ׅى�(|��N>�!�$A�V~�,B�JϗO��	���w�!��3vf�8�A��yvp	P���0c�!�����S1M�)F���B�aW�l!��F:k��(1e�P�4�"4[!�M�pM!�$���IP�F	}�\)Ҁ�C�!��b���i�l�(L�~���g�>�!��#F���I0�	�4Y��2(�"V�!�D��z���eoݡ��Vd�'�!�dE��tJ�b)���!eb2*�!�� Xlu�>B��s��B �i"O�e��BQ�|�h5T�ͅZ�`�"O�:���=/��r�B?P_�-�a"O(��íW�d9d�#5���ib"O�8��Lj��*0������"O���f[	��I�7�TbZ򤺂"O,CT��g
@(�#[="	�"O����cP�o�(���%J$#�� �"Ofu�b�X3V"�`QS*Up���"O���/�8dr�5�U��+� *�"O�t�b�йtPB5�T�+	�mI"O�M��C�d<f�+�4�8X�q"O�L(`,�(f��KN�}�JՃq"O��zb^�o�pP[�*�$P����"OV�۲Nʏ��  �)�Q� ��"Of�rĝ0A�0�r�°�^l�w"O��H�E�xA�i=.R���"O� :�l�6��x�i�1�റu"O�HV+C��00��QE�� 3"O^ah�E�yU8u�'��`?z��0"O� 93��kh&�8�F��)�<ؔ"O�M�WBM�W$2(��/E��蠤"O���%(�e��k�n8��Yٴ"O6]3"֎�N�sH3㔡h�"O�%�sCõ+]��`�(�^� F"O Pbș^έ�`��[Į|Q�"OPzs��k�A(�M�AS�"ON`P.�;8)�f��Y�V��"Ov��S�X�"U,	;��8�t `�"O4���.Ο3|����"�(�"O�{F��ry��+��ȞK��XB�"Ob5g�	�L[��X�6�
�#g"OFpA5��eʤ�g4�����"O ��4'�(j���Xæ�K��a�d"Obu�c�� ����gڶ^�z��*O2YЖ�Ӛ<)�E���+]1ޅ��'������"m>���	K
@�6!�
�'��A��`]q���D��7�% �'߬s�M�֘�(݈;�r� �'H���ƍ��%�E	 b���'�؈b�\'W2	#��� .t=��'A8a�!g<Kb�Di�r�	�'2�@`��v��	`ǝ�#��!#	�'	���6��3[CD�;�L- +�I��bN�Ű�a�a ��άH9XI�"O�����5R����d��֝"O������J�R�Xc_�Y,a9�"O�C���P�J��!I2"�ʄ��"O�-H��
:	�.��f��h>h��r"O8-�u&Y�O�x,0r`�����c"O��zWG"��a �bx���4"OJ���>C��	Z�E7QA^؀�"O$$�3K[P�AF΁	�A01"O��0Q)�M�J��r�R?vSz�Ӡ"OX���P肝���	L5���"O ��&�{��H�F�X)5X��"O ����9.���z�c1PP�i "OF)3u/� J�(@�oR,J0["O��)`*G�����-02�٫"Op��(PL[F0�-:��4(�"O\D@�E�9x%�kl�T츍J�"OJ����6?�$�	(�FX�5"Of��B�W���æ��t�N�"OT�r�]1�|�c�dV�v]�	�"O� .�j2Ȃ"�z�`b�>�՚�"O��#Ӆ��l��U+��!Hx��"O��q���2(���@�>5/����"O��+�������%o[� .��g"O��S�O;lY�8b�=_����"OX���BRv�n$�k�+*(-�"O������8H��e�B낈�L��"OL��EĘ�H=�	�'��e	&�E"O��B��],N�\9h��$h�t@h7"OHՁ��r�܁`�T�A�>�Hc"OXA
�$�=����c(��A� �)�"O2ث#��7/(0ِ�2��z�"Otq�h� *�L�U�@h'�La�"O)X�+���qRN،���q"OpUP�.ҝ9���Ҳ,\�r�(���"O4剂nΏN�~�I6)R��:��"Od����ޭ%����(M:D��,�&"O,L�̝=�������\��K�"O�
#���V!�"���"O�x:Cj��a��낄V�B�� ��"O:�[G��Q@��0*@bX݉�"OLpR��d��8��H-_7̘�4"O�8S� �&�#���r$ftA�"Od�X!	C����A3�ۡ!$:�H"O:@�6@C"�}a6ƞ���"Oވk�/	�GkB ���7w��B�"O�����@�	�x`�T鏟?$q`t"O6���gV~;ɚEc!�LE�"O�,��˺�<m��\�*�L@�"Oބ���R���D1g��<�B�qv"O*if�B�pVx@��cF�4�sB"O����B(�c���|q��"Ol1*�(�m��m(��� ��h�G"O�ٻN!4��[�dG9�� r"O��6eӊ?����)�� ��Xф"O��WGV�(OD���a���aY�"O��jբ9 Z�ʀǋ;�$d�'"OH�(wc�"���FG�O�(�'"O���3�\1a5Rac���SC�Yb"O�e�u荗L΀@S�^%V:�Z"O��P�#��v���c�F2*�H)�"O�-A��ʈT�:��G�t� ��"OB�cb�k@�D��y��+"O���=V��Eȶ坦#;X��S"O��戲�
�	c*tѱm��P�!���1\�`� )���Ye�-~!�Ğ���:V*-+��
��ـD!�ā/������B�f�r����%�!��O�x���a�b�Z�S�^�%�!�$Q19G��(`!��@�~�ɕ�J7�!�d�*B!�\�!M�lP��G�ǃ'!�d :<��Y12N�F��*��}$!�D߭�����(�R@�p&�<`!��!t���gH=q��pѥ�28�!�̙-�	W���
a��K�8�!�6-(��]�T9�!��$˪,�!�D�8,i��)Ӡ�X/⁸R�@�*!�F$���󠪎���0��Ⓓ[!�d��@@G_�O��9�U�f�!��̚s���ذ���5�@��'��!���0~
���V�R#w�,���A=L�!�#a�Ћ�bP�S�X�nU��!���f������F����k�(!s!�ę�d�6�AE�K?-R� E,��5Y!�� �1!FFI-<`Lm��çPϖ��"O�lj��ϊy!�
X<,��0p�"Ol����M�ڐY�J�3�^��4"O���+X�_j� g�Z�Y�<���"O�1y�l!:f���CB@�1�"OhTrB����L��aT�j��@��"Or\rU�ˑGp����N��ز�"OT��pn�J�4�+dDű:@D�R2"O��r��.��ys��!V2@iʐ"O���Q��o��ܡ2"��*����"O4��.)|&&�E1�� "O�(��T�ҸMc�HB�Xa�A"O0���`� Ґ�qЍ�2V�2"O��2   ��   �  F  �  �  �*  �6  fB  M  0U  >\  �b  �h  o  Uu  �{  ہ  2�  ��  I�  ��  ̡  �  Q�  ��  ٺ  �  e�  ��  �  ��  ��  ��  �  �  V O	 � �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R��I^>�Z�l�)N�HI��S�6�CJ.D�Lh!Nġ ٳ�fݒ!�҉��,��T�I̓L��@|� ]	r"O<��w�R9{&m�7 �)Aj��P䘟�F{��i.[�����N�&�6��Х�}�!��U��0C�/��10.�`��s����<��-�|����G�� 3�iC�ą�IH��?�������O�3: � � D�<�%L���.�����%*4�U����h���� ��#��]C��5'�.��"O�у1mF�1�dIU��'i艂��O>�=E��܆5�>=��ҡtN�pH���y�mX�~�vu�g��G491ŮK��yR"�0A��٧�K�E9(ʡCI��yb��!G��p�$��i�^����P�y�eɯ0�<Y�(LO0P�3��P�y2,ئ ȷ�ɼE.x9u�yB�G�6�vy�*˰Q����	٨�y���TN>aJ�������"�!�y2+�e��[����,�ű�hV&�Py��G3h  i"��yD�RAXv�<AU��{1��s�-�P(�A�t�<�4 �xA�!A���O�hH�V �n�<�6J_�\~������Q�W��t�<1@�]�)p�bI؈k�FE�F+r�<Y�[.i�T�9Q%@+||����.�U�<�1��i4�T-�dym����v�<�`b�� �����*�K�y�<0��7qz��ekM y�p�#�N�K�<��:g�����+J#^��)�a.[F�<���ׁR��!�jI�\H4!x�<Qb�ݟ]z��۠�ۙ	H�P��w�<���f[�%!j�?���cl�<����E��iH�
�(fU��Ti�<	�!]�hRU����, ;�N
J�<��ÿ[�F�:a�#u.�G�D�<Y�l�&w��J"ٝL�H���A�~�<��M��(P�\�*�1&����/ZT�<)�����L
!*5c��q��N�<�S�]9�Xt��+F�yFiSH�<��E��y�t�׆*	Y(L�É�M�<1RB�VrȲ�.]�L,�`��N�<�Iƽ2����C�#�^Q�H�M�<��jr�, ش��uX|<�)�]�<��#,�<��嬌�roܵ�u%�Z�<Y��V�-5�i��Z�Ҳl	BœV�<q��2 �d�k���T���[��O�<	�+��>e#f	ڽ��z�L�<\�"C�|�AE��5�F�n�<Q0�|���`��T�*�����@h�<9�.K$.0�hV �BW�1ؔ�m�<��L�*������Y(i��j�<�A�s�"ء�ɐodA0��d�<� ��*c� m����T��+�I�j�<��m6$�4���6�F(�vȔM�<Ʉ�ɃRԀ��DO�����j�p�<�U�ǣ0����Y\!T�����b�<�6E�)b��m��$��H�#_x�<!�Ə/Y��j��@2`f��2D�v�<�F���PD'�-?��dX�
w�<	���%&TKw�Z2G5�Y���s�<y�Ņ;ra�i���­-,�*Ԍ�E�<� ���vcV*w�Mkf�G�<:eY "OXU�B����4\�ǭ�M 
}��"O�T;UaN�I��q� �R�D�B��r"Ox,BKW��X��
M(����"O�쒅D������!�����"O�YAd%ϥ^ jY;IGJt: K"OlDx�Ҍ[�<�8e�M�@\# "O� ���@*`���I�?UM��8�"O�E+��	7z�y��K�>M�A2"O�ڠ��>t5>l�4FȲY1
dx�"OVT���H�p���#� �I���"O�!�"�~��)[U$����C�"O0���Р0��ϟ
��:E"OF-�c��p\�娥�=R��(��"OH85�N�n"���&�Lk>�A�"OlmP�j��i@�d��*d^�j6"O����(G��@����.R��2�"O�qKeđ,����n4��`�"O8dbElًf��0���N	0�Ā�"O�ubQA�7��}؇˔�_/X]�!"O�쳲��@�D�/)�4�*"-��yR�ùF-,x@@�!7�,������y������1Q*a{��4�y�MS��H����V�~Ё�1�y�i��+<!��\��|q�/P�y҆� V��(�r����ƙ��ѽ�yR��q;���B�܄��͉AѴ�y�珳Y�H�Ҁ-E
�B-xQ�7�yb���p��U��\�9&�{���!�y�O��r�:vj˕ 1"!��j��yr���P��F�F�yA�-�gV �y�#S=V��a[��9r@:��g%�$�y"���!�֔��ϫ6����	�>�y���k���״0����K-�y2	]���`Ɗ]�T�2�A�m��yB��4�4�;�ǊNhy��8�y���>^}��8�[B��ųt���y�l	S��ئ�McꚀ$���yBb���8��۪W�؊t���yBʇ]h<e��K�0@9��+E�W�y��
<��=���C'_�yB�֡3��ȗ6��T�CQ�yBB]�=İ��ܢK�^������y�I*OM�$����H��-P��J��y�4R4P;c��1��}�a�5�y��=������|E}I��V��y¨�X�U06D�iEr-�Q��y�)Й3��|x�K�6g���p�I�9�y�k͗)q���qgU.1�F� ����y���Ȁ�"�R>7*&y��%/�yrCƆ}'`��M�,v������y"�L�jd��C��;!�q��a�<�yrLͯL������BQ0��0'�3�yR��zPY��Ҕ@=z]٠JԀ�y�*�/j*p�+#5�jP�[�y2Ȝ'��Y�.P�(�TI�F��y�aQD"`<*��7LF�̢����y�Et 2�lU�D\�Z���y�'��d�,����]�@9]+ʍ�yrD��~��Ň�:$"�֍���y2"܈e^��Rߍ9j
��Vg�y�/����s��1"pP����yb��;Sr��CA�$Ѷ}�$�ś�yB���1F�.1Ȁ�x�*YI����S�? ��r�/�;.�8m���
��lZ"Oj����e@�9B����X��v"O��ȶ�J�DVb�x���ABx�zP"Oư�e%��2�T�O��J;�dC�"O�ð��%'
�:�A]=#���T�'���ş���ܟ��I��h�Iʟ��	,#6��B��gb�9��n@$�����8��ݟ��Iܟ��I����	؟��	>,D:����8�;�N8>Am���,�I����	ן��	П`����D�	� ���0j��F9
X8Q��	 ���	��Iß���П��	� ���8��,@��Pb�OG�Y�&U��`ƌyf��������۟���ޟ�����h��ߟ0��9��S�e�(���)2MO�+�44�����	ʟd������ퟔ��՟�I-j�J�C��)��p�b%%� ��ߟ<��韔�����	џ���ڟ(�I�d�ڐ�S�I���J@"=ؐ-��Ο��	�0�	ӟ���˟������I�egpa����knA� b�X�N����H��ʟ����I����I؟��I*]��)�T`�Q�U�s�[h�ځ�I����ß ���@������џ��ɦB;�QAέq���JE�@<�Nx�Iן(�I㟀�IƟ`�I�� ��۟P�ɔR�*x�E�8r���j��_80����I���������	����������3,X0�;s�, �0�G�M�{�2x���<���P�I֟�	ß�ߴ�?���"������Y�_(��7��'/�W�jy��'��)�3?aG�ii:�����x��Qi�+2���Q�Ǉ�������?��<���U��X��ڎ3x>�KTe�%�2�Y��?���W��M#�O$����L?� v��5P@���f6���ä*��ҟ�'�>Q�g@�8வ��-m�Xke���M�%�u̓��O�L7=��<#7�f<Ѐ�1J@iٵ
�O���b�ק�O�xC�iW��֯$=�hĔT��\Z 	�<|��$j�LI���=ͧ�?�q�x���*Ō�3����M��<�/O6�OnuoZ�7�c��� �C�p�|�q�7�<���Cl��l�I韜�I�<��O��Y!�N���9U�������	(O�34�5��(N"�U⟔Z%'HjpB��ҜJ�"�X��iy�[���)��<�u�:�pP�'��h�bb���<Qұi����O>�m�R��|:ѪR'B���#�;ym�4�+�<q���?9�N
���ٴ��d}>��'JI���Ti��p�	ӎ�$��Pӄ/���<ͧ�?a���?I���?�wi�\�u#��J����A���Ħ�jp��I���&?��I�GٶPJK����5� �r@!�O8Hn�2�Mk��iQ
#}bDL��E�nˠa�U�~���]I�p��4/�~bc
W@F����'7p`�O���-O�q�pd�?�(8[�-��3���O���O ���O�i�<1V�i� pA�'휤qU�IK4Z�:�O3�X���'�6�$�I���OT6mӦ!�b/T6X,̤��%� rø��PM�_w�9o�f~������3h�O����7��&#��w��ʃuez��T�	ݟ��	ߟ���]��U��Q8��&Rw���ȑK���x��?I��i���D_��T�'��6�:�ĒI���kEK*F=!4cL�i(E��}}2(iӆ\mz>m��
��Y�'�$8�N�
up��EW/
�)�PH�X�.����~�'��Iş��	���I0Pɴ�s����}��a�6P�P�I��'�7,U[*�d�O���|���
svT��h]�N6�P���z~⊰>�¼i��7�\ݟ�~��&:h�����=� I�8i�h��jC%`P�Y2*O�˪�?�gi!���"o�� h���k�
��A�v���O��$�O���i�<QҺi¾5;7��x=ĔУ���@�L�%�+s���'��6�4��-��DV�=�E@A�SN�Q�H�3U����;�M�@�i���h�iw��RWJXq��OK��'�X`���`Y���/C>��ə'����(�	����	П<��I����]�J�{�bH9G�h��h���6m�K�P�d�O��<�	�OH�nz�5H� ���D�v6"�	*E@��M��i����>�|���M�'���P��m5ԉ"���B<��'�z�����8(4�|�Q���󟘫�"X���A�ɛ6��=a�����Id��UyR�b��|���O��D�Ob�0FϼBT,ɘ4-G�Z��i�6��)�����ٺٴV�V�T�qh�#�Np�5� ���aVd/?���1	8ʼ:�lˡ��=����!�?�3�19�*�S4�͸Xb�㱩��?q��?���?i����O8��τ�B[@ԁx禁P ��Or�lZ�>� �����Đߴ���y'�\&0舰��� f�J�P��H��y�Bh�:n��0 � ���q�'�J�r'�H�,Ǌ��	R�L�U:'
�(v�<K'���#��T�ܕ����'��'���'ZHL10	U�
�ԀG��/ Dn��T�h�4>7~1���?��"�'�?)�4n&�Q�!�h���T�����SDV����4<���"t��E�d����j"�[<v8��hf钸A�0o�X3�I�KE<����'�b�%���'�)��!< ��T��I�
�n=���'��'�����S��+�4x�@C��#�d��F�1Z�]IC��+k*Y2�yj����[X}�Jh�,�m�П�#�L[�!�`�3����q��˸tN�5l�o~b�	�,�
e�E%BBܧp�k� ��#O[1����J�1YV�-�R3O����OV���O��d�O��?�6ޢ/�L��j wA���B� ���I�4qZ��̧�?qd�iB�'® �J��4

��Իh!R�� ��O��l���e���_:`>�6�+?Qv틹f�ˊ.�Z����әr���%���Z
���{�Iyy��'C�'���97/����D��F�� ������'h�	��M���қ�?Y���?�/�Jl�P�օ=tZ�q�Ö	 d�Ǖ� ثO yoZ)�M��'x���L��;B@�����
2o�@@e�4��DK�C&*��i>]������v�|��(�ԅ1�,�*T�!��	1(�"�'���'s��4]���4R���s��E+U�L�[1�ݏP�8@�FG�?�?��;śf�'��i>��Ox�mR�d:��k�ą3�Q= j���4K��&o@
Y{���t*u�m��ԦmyRm̀b��9�7`-nb���"��y�_����Ο��������ݟ8�Ob^�;���U�`PӇG;IX4�*@a�`���
�O���OԒ����N���:$�(9!��D�f��!s�CQ"Y�	�4gM��8O�S�']{n�Rݴ�y�(�9�=���WA�w�6�t�|���TAɶq��x�kQ�	vy�O�2��� (���m2ت��Q�B�'�b�'m剠�M��ʂ6�?a��?��J�-}����F�5Zwڼ8Q@���'
�]{�m�b�IC}rl�('@��V��^,���Q���Y�q�*��٫F�1�P� V!y��2��;ڔ�1�b�;ADBŲ�'��p=̉.�M+��?����?�J~����?���h��B!%�7b�x5s�ɓP5*��5u��+L/f,��'��6�-�4��n��R�|i��
,���ӸI�$L֦�h�4-��v ��&֛&��D��-w������1p�-��l����}�����'f��Oyz�4���T�I�\�I:7�Qc!�	Q( ��I�!Rq�=�'a:6�1�
���O��埀��=���I�fB� k�j�.���jl\'���'���i�6��p�OȾ�۳��8�Vl�A;F7<� 5��C�>�iDX���p��\&�q�wyKK�L���ʱ9d���C����'���'��O?剃�Mӗ@��?0�}+Vű��Z�y����+D=�?��i��O��'sd7D�	�ش�6��/HT�9%
�.�X�E˱�M�O���.���r��*�i��s���4�F��J�=P� UC�h��<A���?���?i���?	���'E���B o����GV�dl2�'-�%k�V��<����AʦM%��+�ܫ6���vDF1�~MX�W<�?a+O���e���
+Gw�6�9?�W��83��Q���CE	�2o�.�,c2+�Ol(SN>q*O����Or��Od�O��%s�lw�؜LB>�V���O��vћv�
(�"�'��Z>��Ъ˲^R����4��2Ģ+?q�Q���42��L�O>b?z&_�V�lx�2f�Y��#ܣw<����1O�����JПDі�|2+�*H�!F��4�0$�
�2�'+��'Q���[��3�4$ؤ��@^U�@m �NH@]ޙ�����?I�r�f�$�{}B�aӨ	Zp��j��9�cn	WT*��q���9#ڴ]nv�
�4���D��)��'XT��O�F�,U��ݫ�[���Y*�`�\�'8b�'�r�'���'�哎^��%ô��-m˂A�[J-���ܴT������?����OT>7=�Р���!�2Q�P)�)ւX���ۦ]�ڴMW�Q�b>��ŖڦQ̓`�ұ�BK��+��c��N��<�+� �3H�O�đM>�+Of��O�Ż���x��肤q6�=�ׇ�O���OL��<AҲig��[D�'�B�'y��`�&:�P!ӢL(�����TC}��a�&�m���M;�P����挲c:��d/�	Fҝ(��:?�C)��u��[P����'b���$��?)ţ9Y1���jB�`�ԝCO]�?����?)���?	��I�OTHq@�r��pi 1Mw�*���O�0m�1{|,��ן��4���y��`e����	ۢl2�j�Ʉ��~��'ݛCo�Z-�%k~�z�z⽹%����e�>F�V �KJ�p���H>	-O>��OF���O��d�On�)�œ�l�\a2FJ\Q�2�+dŲ<A��in:3��'�2�'��O��Ƈ�*(藁I�r�D	pw�Ł#@j�LH���t�j��	M�OT��0q���6Q��)����P97l��)�0��Q��C%	\:S�")T��zyB"��{D0@C�m�NdYcȐ	��'��'��Oi���M��C�?Q����6*rC*.ǈ�k�ჾ�?���iD�Ox��'<�7��Ǧ�jߴ?�Q��P�J�1R�9z�ī�ǐ�M��Ot�1���J��=����[q�_Ҏu`�H�oF8ȫ&�F�<Y��?����?y���?A��>|C��U ʄ0���í	%R�'Bjo�J8�&1����֦�&�HC@��1�. �U̕*?�P����?�ODEmZ��M�'L����4�yB�'��yg��f!dKu*]�&C�+v��/p�ĉ�I�T��'��������쟄���oL(��e ��{2*l��ʛ6U���០��P}��j��g/*	��ʟ���$�M�'H�
�+BI�$���b6M_�@]�|�'e˓�?�ݴ#������Oy�fKY�/J`���͒�(1�$D@�l��!��g��Uv��?ISf�'XV�$�RW��,C*�Ȗ�RpE�e����ퟐ��şD�Iߟb>Ŕ'��7��<iVƑ:��!EWn�2��	*']���u��O�����?�Z�t0�4��A�{���X"����yV�i��7m	#t"�6M`��@o��nT�|�'�O����?� ���ũR?xr�#��XY���g�i�2]�' �'`b�'�'e��%���9#@[�n�E��IIOHYb�4?v�l���?����'�?�Q��yg��='K��6���&�:A�a��95&&6m���E8���4�0�iꟜXs��v�,�3���%x9x�r��;Nh�	/1,��w�' ZT$���'�'1�)�`�P]�!a��[,F�Ne�@�'$��'��\����4P�V4"��?��	;
,zPJ�1
(u 2k�9�hͣ��E�>y�i�66M���'�:P�`'öٸ�o�2���c�O�mSS�"Fq@M��8�I�#�?io�O���.O 8�Z��F�*h�m�CG�O��$�O����O��}���d����*!,i) ��[�Z�!�f��A�-B�'��7�&�i�1��+�0FCPQ2�Ŭ�� �V�j�A�4
"��b��+� o�Z�\�eA�m�JEA�$��	��P�4KʡH$u��IX������O|�D�O|���O���R:�����Ȍ�(�z�j1:Vl����Ζ<�'�r��$�'_ܹ�7�
�TTb1dE$H�� ��>���i�\6��韐G�d��s��4�#�I�?�q�P�^�	n��gϴG��I�z�"A��'��&��'@F�C��6XҰA�s�5|�pU���'�r�'�����4\����49�lq#�~�t�#G���	�uX\���-y����\y��']��/`ӄiy��^� ��`vmB�?'�7M"?����u^��	�;��'`[k�e3~�{�`�`�8�����^���O��$�O����O"��<���쓔@NDUisfI�
�I���I�M�%H�|�����6�|��]�H��`�\4��t9u
����İ>�Q�iG� �'g5��4��$ԻD��p�'0D�X��U�b�$TD`N��?�$�(�$�<)���?����?��䘊F�ތ���i�L-Z���<�?������ަYBjE�P����0�O](8#���<nv�	(��*��D!�O���'Q�6�Ħe;���O	�[�+'mv�p�M�#X�s��$,��Be�	Y��i>��`�'9da'�P���#�(21�ԕM�D4 �mGٟ��	��	ʟb>��'�7��?j��8��3j���h�U;�����O��DKϦe�?�cS����4|:.)�����8���A')uPM��i�7�P�=�7-,?��,��iB'��d^y�T�� H��W`
Gc��r���<���?����?���?i,�F՛��ܶI�12%F�%3j��$�����X^���	Ο�&?��	��M�;N�f�͙�&��p� �p�t��e�i��7mAɟ ԧ�O�~��iC�^5)�!	���o%r����H9U�D�~ڤ���B�O�˓�?���L�8:���Ϯ4�� ^I�,!����?a���?�-O�,m5`4��I����kTu9&τyr��`5l-a�F��?ɔ\��ܴy�����O��a��9�1��G5�CEХSd���'�j� �(�P������4���|�$�'�a����qr�9���S�Y��'���'���'��>��	e�BT�Rƚ=8�ʽB��#r�D��%�Mf��?y����6�4�P8���Q�uL��m�>����A�O`��jӂ�l�\��Tl�]~�rFv��s�y�*BW|:d�1�\4i�X�Su��	����d�O ���O����O�dnQҵb�_^\�EO�}�V��PU�d@شu����?1����Ou�آ�n�004�)�U�-��ڀ%�>���i5�7���@E�D�G�W}6ԁ֊B�0�\��U�7��R0d���I?H��J��'uX�&��'�B�Qb@&2���@B N�{�l����',��'+�����P���ڴf&����vԄG�Tw ��dЂ8M@�s�`����A}"�h�"%m��MCa�̝�l}����.�Э��I4gD��Aٴ��Dъ	� �J�'T���Tܮ1)ASt��-  ��2N��u̓�?���?a��?�����O���[��Q͞�fc@b������'N�'|H6�]���O�m\�1�dT�A*j>bx(esv����������|j�X�Mk�O���H q�0�T��;ȑ �o���`��GeғO���?����?��?(^q ��E�u�P�s)M�&D�����?I.O�m�:T�����R�N'QZ��'�^�pM�X�ɲ����y��'v��E�O�c?���'D�� ��&+ǵn���`�N F�"��n��m��������*f�|d	�6:�eR�a�?M���qb��\Tb�'	b�'z���\�`۴N���2��b�����I�T�`�D�?!�-T�V���W}��w�4E�.	�n�(X���9R�X7I֦1��5�oZ~~S�O(.-Q�	�V����D�̑����aB2�/�:.��<����?����?���?�)�ح"�Js��p�FBYk>�y�pI㦉�F)ӟ,�������W��y�_�X��Hȕc��6J.)��T.�7�զ�����	��6�j� ��n͔AD�Cw�[-qIDePf�}�x$��2u�r�FF�ry�O#�{�����ǡ+���%� t���'���'5�&�MS�ϐ��?���?a%�4d: SQ�G_�~j#���'@R�``��,x�b�oZ��D�4F��9P`�Vh�<ZP.O6��	�#�D"a�T�r2l'?�B!�'l2l�	<o�p(A�K���4GF��GT�l��Ο8������u�O�R��*<=H��FL�BJR5B��I(8�g`Ӡ)	Q��O���ߦ��?ͻuO�A( �1�Q�1�G1p�n�̓A��6�b�z n�5hT�nZ^~RИc���S� �Pxr`	��ܬ�A�çA�X��#���<����?I��?Y��?a����7Ht1� �3`���EP��� ˦x���ퟠ��Ɵ�¢�M,M��q����A�:�����M㴼i�D�8ҧ8\>`��.($,dċ��n��h!D�I��q�-O������?���?���<9�M�9�ఔC�-F��QF�?����?���?ͧ��¦I������l@vE;${0�(V�^�֤����Ɵ0�4��'��H����v�0,oZ�
��P�O�G�DA�q��f<��`ئ�'6D��� �?����tD`�1��@.cU�=��,�0�n���p���I؟���矬��埠��aA�6\��Rv��c�a���}���?9�*D�V�U#����'�7�*��կL=�<�D��8t6<� �X#W�^���Cy��'���O�>�*��i��I�_�~#� ./�����dOY��]���` R��N�{y��'~�'��bV�Ҝ)���7���WVR�'�剁�M���O��?a���?Q*����*@��2#%\�A9И���O�m���M��'���v�P�H�56*-UE� ���ZsaV�ؤ��ۢ^����|2���OF��M>�&�Ԥ����S&/���2�듾�?q��?I���?�|Z+O.n�|��%JT�\j|����7_��K��x�ɯ�M��"I�>!��iĝ���?8( ЭQ��iJ��|�2Pl���rӖ���� ���ݘ*O<��Ш@�_����go��> ű�8O��?	���?���?������)f92�z�昽6P��� Q�q�nZTL��	��IA���r�����a��Z�q`B�Gx�T�জ=�L���I^}���N^��:O\-3F��*i�z�r�B�]����>O
�rD����?)���O^˓���Or��P�e��	�į�t�Z��v)P�`�Z�d�O��D�O\˓Z���R�n���'�g{Qr-���/s�ԉ� _�N|�'�bm�>���in*6���]��O�-I�#՝&}$c�l�":�d�×�d
�ʙ�&:(���n�S� .r�����+�+PU�A��j\BónO���� �	��8G�$�'���Ï�E�9�׎��F��<@��'p�6��6�����O�Eo^�ӼC�N&BSB����Lp�h�A���<!e�i�^6M\ꦙ�s�O����'�R�����?��܉#�\	WeQ�k;������]�'9�	ן��IߟT�I̟��ɨR���rD拻�;���o��=�'�X6��5lǘ��Of��<�i�O,i����3���06�Ҕ5���)�lWT}ed�jYmږ�?����<�|�/ȸ{����`;w��Qȱ��n ʓ=�d9���O� J>�.O~T��m_� Q�i	��O��XH�L�O��d�O��d�O�ɺ<�`�iK2(Z��'��tj�+�[��yBi��tOnxS��'��6�+�ɬ����립��4O}�F���1�.P��x� �C���0Rq�iZ�	��0���OaL�&?��[c�~q+��,;֑x�k��z�֨)�'hR�'���'�b�'��%�ENݏ@T���eR�X���<9��+�*�.����'�7'���GT�3a/H���!���T^p�I~}BbhӪ<nz>IYp��Ц��'%>H{`��(���o�C�p0��Ǆ�3��y�I�x��'��	쟰��ԟ��ɾh��Ae����hR��ðK]nL�	ҟ��'�`7mC�d���$�O.�$�|Ba���4����: ����t~m�>�Խi��6������~�F,ae.�1���6��ԠB�En�ɂ�h;.��+O�Iâ�?�sl&���� �s��; �<)ĉ0�����O@�d�O��I�<�1�i����f��~�P!��C����&#K"@mr�'��6�3�	4��D^צ��b�!�Lp blU�e��<�B��M��i�Ҝx��i���� �H� ��O���'���[�SXi��$+�!�'��	��h�	�0��Ο���@�Tဟ���E�̢8�H�Ra�GS@6���@�D�OV��#�i�O�mz�=Xen�j���*W�����2Ѓ�?��4Z�BR���д��"���	/*�ة�q��*�R@�*�扈+XU��'+ P�IoyB]�T�����Ćȡ7O�z��:-��u�S#�՟���� ��ly�i��5��A�Oj���OpU��(�&Z�@Y*.~���5��3��$G禽��4���l�>Q�.Nb}�0i WpBⶪf~Ra�Ӣ��h�42��O��@�I32�RB~a�0A�o�{�ఄ�\�(	��'�"�'���Sȟ���8P�+�㐖>^ժ��:�4\�����?AG�i��O�m��Q�fo�-l��J��I40*�Ħy�4*��������f��p�UI��jn�DLQ�]�:�z�Ȼ1�� ��	�Am�&���'�2�'�R�'�B�'=&�:X�F[�,�t�(��RAG����Šu'�ԟ\�I��0&?Q���F=p� �O��)	J� �����(l3�O|Ym��M���'��>B��B)"ka��#Q�CT���"��#R'Uyb�o�V\�ɚ8�'�剢+��\r�哪ZQ����V
�ڑ�	����� �i>�'A�6���U��$U�Z+h�r�.�Rq�x ��t�T��R�Q�?�%[���ش^���nӢ����:L�٣�E\W��$��hςe�6�<?1��Q�|����P���i�k���[srebPK� [4���鎋aQ��O��d�O����O.�d?�S3� s&҇�Ɯ�blSa�j$�	ɟH��(�M��,M�$Cb�B�Ob!�J2��VBA&]{��hAa�� �'�87mΦ�#:���nZv~���� ��( �Mu���*r�e���\;���`ܓ���'/��Pʘ�?�dH�#!B�k���B5�}A��h�<����79`�W�1F\��>),1Q#@��2vf�q�$T��t2�#ԒbIB1��!Ө�KPB�!P��G��)0��
X�.��SJ_H�7��YIT `�k��x�Fb�{�"�qU�l����AsέP��9smVLkUFL�~]�q�:p��$B�b��o,@Y�"�/%��T�dDܴD�6��OT���O|�IO������ߴ'��a�@ě@N�	'����ȟ�(�
ԟ�'����sQ! �JȻ/�ȅa�iP�4�U�ش���_�`�x�mZ��i�O��HZ~�.H����! G�68r����ġ�Mc��?�/?�?	L>q��Tf��<�rtS��=?�p2�
�#�MӠfHa��'���'z��F,�Ɇ<2F�ф-�@f^	��ݔeR<(�4l}0Ő)O��D�OΒ�����O�h�@ɟ��й����~Ǟ`0��䦁�������;C㚀����O�Ӈ
�JHɡg���N���MP�S�yR�ͲQ������O���^	u$&Ac����is��qO�_��`�'U>���'�U���	�$h����ѢǞS��@ZVo�up���O��q���	˟��	ܟ��	ٟt��dвc�Aʇ�»
$b����W�Ce�I䟬���P�Ir��T��YV]����a0l�cb9�\�����Q2��?����?	��?��ы�?Is �q��c�g>:�=؆k��s[���'R�'��'B�'�,z���!�M+��.T�>�PA�̹d�j��w}b�'sB�'|�ɍb-�0"O|2�+�O����36�������ݛ��'�' ��'X̙��}R��	ш��c�^�����!�M���?���?��
����O������c�v����n�%�6��3���&�����0���1<��c��F,j!��q0���'n�nZß����8�r���Ɵ �'����'Zc.���<Z-@`e��+J���ܴ�?���������M�S�*���C��2�`@�cP��6 n�(vD�	ǟ�'��4�'"X�$ねL�h�|��4�"]r�q��^��MsBڴDg�l�<E��'����#�	�B��ű#�Q%M�Jy���'<��'3��'(��c���	m?qtJ�:�3�(��B�y����p}��'<R��%#H��ǟ���Ο��{�nAh0H�Ũ<)������n�Yy"E�|�)�[�a��N�D�p�h�F�.�"Lj�Y�x�pM���$��?a��?�*O8�cKN�S��Tg��prx�6% �4y'���I�d&��'7n��S'�"`�`X*��b�E�ͱ��'��E������ݺ<?���#�8½�d@��y�)��U}Zh�e@�J��C�$��'9ީyƠL����⊬����2e��m!!�n]-n|�WaH�M$\���E'�Vl���R$q	�d�������ò��Bҵ��gE�%5Լb�J9&����_>*��Ȓ��e)��)7d<0�S��)�@P���Ԝ��r$ϭ�"@��.��EAN5p��
� �2��z;��;4 �k�d|���ĜS�������?1v.Jkc�LI���=FTA:��Z���i�Df�@q��R �$#��"��V%��Ɍx4ĝ�F�^�Zy 0�R.����S@҈F娅�Oހ��暧7�"��.1`LJ�X b�O"�lZ�H�6�)���X�iG1A(����Vl*�B�	�r��c�χ+�FxcE+UJd����g�'��xsR [���b�o�-��rej���O����?���I��O��D�O���WԺ�FfǜorT9� ���bfHY �	]6�E��>��3�h���L>��J�(���QjQ&�t�A3K��p�a�/�&�9�J�ȴ�}r##�Ty�f-��Ȑ�v�0�Pe�+�x%�	{~Z`L��S����	���cA��7-�jJ�(��i�ȸ��~h<�q��-T��h����,&n�Q҆�a~҈4ғ��	�<�ń �m�vѫhh�t-y��E��dT�	��?���?��h����O ��p>}�.S�c�mR��r�*}�"���<R����?U��l�>|R���w�I�m���,�zȆ(���^�iE��)P�X��&����æa�6�D,w��b��T#���K>q���(�Y1����]I�F�B���#�M�Q�iTBV�D��F��[�$���)�����cH ��U��U�B�ؗa<A����B��K���<�#M���$���N|*G�>u����\)/2�|3��O�<	f&05��d+�(N�GLār$��K�<�I�2�8$@	�X[�u�Bc�~�<9�-������.π`�Pف' R}�<��F�>���Z��˔<͒�)�kB�<a�%�NJ�I'MD�ka��C��|�<�5oثrĸ]����(�8(jU�|�<���U�3b��� Ȍ��pLB7l�u�<i�$��M��&Ԅ��T�%�y�d�	h}L�J�΀,2�r��W;�yB��)z�R|�1�2Ft|��0N��y�B�X%v�����J`^U����y
� ��Y_�gt����T,��}r'"O�L�òA'00ZA&ؔ0��}"Ov�����f!�Ef�(8�%�"O:89&@�`��=Hv���7� �V"Opr�a�j;8����ۏ$��"O@D�@+�P�t�0��~b� b"OT��dN9Y�	{u�1��"O�q���8�H3@ڍ3�^qq"O,��āB�aXX����ȞHN�"O,`h��*����#��)��"OJx��;%Ŭ����8N�x�"Op�#��ըB�Z�B���	k>��f"O���Nk��8rp�\��
u�"OB�2/�
�XSAҍXK5H"OL z0"A�&(A���:K�0"Om�`̈�D
2q��@ۨSH���"O�=0o��:���SVo=���t"O�� �+qެ�G��)B�S�"O��"��:�~��Q�Jlȣ"O�������g̈́�z��"Oh�P���<�X鳔V�e��"O��1��e��  KA��zI[�"O�񺰋�<���I� � gܞp��"OVh
���d�I�@n�	:ܤPq "O�8ڃ,Ĝh2�m�����k���"Oj�B7��3�n��6�1|^m��"O$ ��U�\M��R`�f�4��"O�SeD��	��D+t�X�t�1"O��@��^�(t��@^��"O��R�18' ���dK�WI,��Q"O<���Q+�d�Be�HdfAyf"O����&�D���cR'pVXHf"O\$
��XR���dF�h�p�r"OL��!Ȑ4�ĩE&�zaF��"O�,�U57@&�"2�R�)�LM��O��2�$�Oԍk�%M�4zɻ`��q��L�7�'�ƨ07����	$v��c��-N��P"�?D����Z#SĒ����+{�%"�+�^q���)+�ar n�t�	�a�U�Rg�C�	�~[*�b��	t���J��Ҵy��0鳭B	v�1Oģ}�4��	2Fl0Z6�q¢I;
zZ5��)��Y���d�fi�s�A:��)K<ў't��W.U5v�Xڄ��L�|�J��1e�'"������<�,U���b�����|I,��ԋL�XpG ��v�Y�7F
C��Pː��!7��I�d���=�����/j�đ�h�;C��×�4r��'����2G����		ָ1H����Wnp�i�� k}�%V%��DB䉔�ʴ1#���	��LK"/�I���\;Q��h�xN�%�'�Z��O|�`�Q�A���/0NHP�Cѭ{ vĻ�N?D�X 7��8rz�X3�@ X���kD�%�?�!�_����A����4
�����j�P�M�sɎGY�ѱ�+�o�
8��Iz�p�C�%M!'>��+��+2�!���8MdV��5��:`?-��.C9B�̌�Bj�^���h�#��t����tb刐 7�	��"%����t���a`�?�7-_�dy�5�_&A~�h��ʟ5<���钑�!��<���ę .�����F&�\��1O+L��*\n��Uc2��%�0Q���yW+kpP�[Ӫ�WD�( L��y��8;�����MN��81����l��ADR?^-^���#�3�<�+^w`��҃O�w�qO�8�Q���`D��(� B=JTh
��'�A�Ca�*vXsV�@0Z͔�z���
o,X�{5�eK`��D��G�ب���݈7��zR��l(�A������G�ֻ��'>�Ъ��O90�hJ�D������:/~��'۞z�=�t-Ŧo��yx�%<}�C剹|��bI7�JY�`�U3OI����g�v�r7���j�4����=��aM~�<���z',U#m\���
kPR��'��@K�c
�:?�1j�G_9 5��U�����@.��	p�a�r3l�S����
�1b�0�8"1�>�I��-q�P�VY��� Ԉ�<	F�X�M��,s�	;~V[������ �0��H<,\9TL,7������)���q�ʅ� E��q�.�8��O�G�<��`�Uu�=l�4����K�gp� ����G�I�3�I�䁀�@W�t��}�iɾ@�2�"O� H��݃t�"ق�͆��\$��/�$<�6�F��O�a�%# W���ͻb�(A�fmǓj��5b֧j�jl���0�f|���ֆ"H(@0�L�=`����'bN.}X��G[�	�<���ïv���"���>@b���q��W �l�%靲#Y^���7��+RW �`��޵u. ��`C�%ǲ�?��%cC�J��+�`�},B��co4D��B'���@V^ ���ʢ�&"��4��	`�"l	�-xtf� �����C%F�-^�b�zFE2UȨk@��r�<�V�H;z{"Ay�c�3-�~Њ���4(��	�W�68�����M�S:�"�<�,,h$�ϙ72��%( ��R��ô$Q!=��
�R�<q8����%���(��Cm�f��/�{�\��	�*eh@4h{�ʠ��"؆ȓ ���[_-����A,P`��ȓ�@+Qa��w	Z��t��?^Pq��w�&ؒdE^����[��6$��	�h���*=J� KN�"0��ȓS5N$'ϙ9|�8�6�@/`M$!�ȓ0UF���ŎH��@�/w\�@�ȓ�����Ûpil���U>U���ȓ.���{0��<���i��<	L ���h#s�ƺ6���©��{��ȓ\d:8 ��˥hc��!Ū�	ܩ��{���xӁ�+BvD`"���Ze��ȓC�\�K�e(PtǁE|���mUԙb�E�Q����Df�+rjՄȓx5�Y8!���/r���*�
8ھ݅�vA��Dg\�e}�M�P��xd����	`d���dڲ[�F�Zr�74x��{�|e�gg۴��yr��ع3�깅ȓk0*�K��]�>�:Ub�a��q�ȓ �-� ���c���6�Ӊ"�����T����<BGRi�&��+�l���k�|��	�%}��J������C|VL�G��	^���q��əE,<������7�Ƈy)�� k؞��-��-������N��܁Q (��)��s����S�DliQ�Q�gaɆȓ4�2�![d��@WL��j��@�ȓD< �S%6%�p���//����ȓ#|PWʆ�|U<���S.|�Q�ȓz\M��m�*-��P� �F,�J��ȓy� �'둑B�e�w)
)t7Щ�ȓ��Qփ2/�n#u�D�/���� �&����Y�'V>�B [� ���ȓO�����HE Hi����P�ڰ�ȓ7���qN��VN�I{�iH*p����U���&��D�(ň��G:�0�ȓV���2,�:�^����\$1K֭�ȓU�[ê�N�قI�$�� �ȓ��˵	EgB���ˡ6�9�ȓzL4Ng{2���$^!�t���P��rF�&vb\���kѪ��ȓFpZ1����*ܮ��򬜴!x~�ȓz��	�`̎X�q�0�D�A��S�|����ͥ"2%rW�̌t�걅ȓ�n��p��3H!e��	�����9�$���J��o�xء�H�>9C�͆�`r��'�M�R4�4��7\��͆�D��PPG��c� #E��)vU�ȓF���R4�Y�V,
�YF$)��
\�0aiI�H�(A���T�̅ȓZ����Q�h�RE�ʑL^�A��S�? ����MR6��j`�9B^�"O|͸mRyW�YHEIV��r%"O�@��NZ�DRh�!��'@,|Ԩ"Oƌɷd[{�j)���F�T��%"O���茬F��E!�L�HU{"O��˴c�s$���B����xh�"Oj�b�G�0��M�U��G�A['"O��ٲ��ej�I��!S�άd"O�������ʃgݎj�\�ɥ"O ��Ao[�hh}�f�/� P��"O���rD��S��s�#H�#�fc�"O��+6-�>X ��@M�8=F2��Q"O���[���JD̊M�J��$"O8���-З߰1�
&@���V"O�#�\~��R��/l���A�"OJQJ����f	D1'(�G}��!"O|E�2����JxSǦ�rn�ٕ"O�\��B9�d��M��hc"O�KQ��59��0ze�Ֆ!4i��"O��`f��=�踨f�M�a%"O�Tk�l��X8����[�]J�K"O�P���K�o�2%P��XR,�%"O�L��O�R��m�JǇ:W. �"O���Aʶ,ʬ�hjOtdhQH�"O4x�u&
�=���yԨ��n\u�"OpX���#�*�Ӷ���n��X 6"O\5)p��#G���p����qe"O�	�a	kQ8�)G�H-~�y��"O�#�
2S�"�r�(P�R�"O����A�/:+ʈ!�^$!�\Ah"O�ٹ�gǸ',��ñ�ѣw��AH"Oh�*h�q��P��(t�@"O �ơ�D��t��kB 	�~�('"Olhy��6:`J�HU�J�t�"k�"OP1a��c�t�Rj!��"O``�&g�{\Հu��C�b�"Oy@䂥u�쁨f�_U�t��"O�M�-���*�p�GV$CF��"O�:2�%��PP�_�i&
]�"O �0��\'R���
_">hh�U"O�qS��Q�(�Wi��L(�"O������s)t$xPHW�_��I��"O�|���(_��d���S삜��"O��sV$O�}ƒ��"�&|� ��"O�h��
��zd마v�r��""O����i^�f��L��A��X�"O�����D[6Nс=��={#"O��D���8K���������Ye"O��{Z�K�.��.B.	�c"O>����G��葶��$>H�"Od$C�IEq����!�6$����"O��k���h⬄�fKV�R��3"O���PK�8 ޥA�
떵�"O�`�I�Lh`5��R���+�"OP��7@�)�dEK��Ė�l��"O��B+�-2�l�a/R�6�8p"O0aկK�����B�<�T�G"ORl��Ҁd�
�͘$j��EXu"O�H@��,my�@��NRSF�8 �"O��ce� �,��D.�j��HU"OHE���\9���kY)y���U"O	��&��a��!X��FN�X�*�"O�t����7�`,�h�C�:g�!�$Ԗ3�̒`��;Q7�偒i'�!�� ��رE��\�3��7{Pu��"Op+W��uI�u��%��$U&$"T"O�p��k���z�E�$C88T:�"O<�c�) �p@���O<�M�T"O�:�
W;j��FD3j�@��"O���«�#X��"�c�#h�(a�"O�]s�Q.B:t�ѡb�Gߞ�JA"OP�jG'�;)]�H0 "]�K����!"O�`PeB_�C٘51��_�x(x@"O��jGAZO�>�S&\�H��"O�1i�
��� P%޹	)��b�"O�]a��X%(��|a��I�8Jp�"O܈j�É�4MK�>KL�e��y�\�"7�m��ΏI���uh���y��"ꈒ�"°�f1�䄗)�yi0����
Y�x"�mD	�y�%ˁ2Q�l
4F��Y޲��S�Q/�y�ہh�N�+t/YQFnqV���yr���9�,7JLKm�L�5eI��y��S�]�Xe0� �2�~-Y4mJ��y��̗G(����H��%�ӫε�y�mG-)� Q��t�
d�c�ŭ�yB�-l�\e!��pG�x2�ⓝ�y�"v%@`wǗ�9X��;⍈��y2dR�$������+���;T@�y��L�\��� ��q�{f�Y��yB*K�n�6�r�����!�ܘ�yrH��|������ԛ&��p2`��y�Fl�䬸�d�~\|�sF����y2CH�$�@ju�ɳ@!�8�թ��yb'�o�Le�+��2��UFP�y������Eлz�Z�G@K5�yb���7�=Ӷ��q�
 ��B��yb��i58 f� :>H�%)��y���J����]�,xN鉵���yR�#hv�x��� 3������M�yBG!�.�J�$(��=��ۉ�y��M����+�)V6��� ���y҄8v�4��`�T�X<s5��y���u��!i�}
D͛�cD>�ybZ�V�KBIzl�*C��y"��
T^��PCa��	�ԔY�f�	�y��WXfL�
�����k���y��&:]�d %�9y�x��4BȔ�yEϢZ�zĀ�u���˱�э�yR��7��������,� M#�yB�X kx�8�%�\?v�6���I��y�j�9<.�Kf�­?��űe�˘�y�EX>��ڒfʿ��䱳���y"��N 22���
�����W�yR��
���Aj�64 I�)���y2�R�QY^�[�̑G`�RT���yB��&�u����=f��4�c�K��yr
Ӷ�4qva��YH"�1@����y��ȃ|�uكf�z��[@�Ӹ�y���+;*�ၣ�?	�`Iٗh��y����Ab�������|�,� �C%�y�G���yq�EJ|���1w���y��[2>D��P��&l6�G(�y�`˭X���4	ıS�fl�v戛�~��)ڧnU��[�LߦUj0���կ�8P�ȓ�搃F�N�k�L�
�)Ozy��iІI ����h���%�TY��me��Ӣ�?�f�#��D�mu|���S�? ��yTA�+C��H�L�C���zיx�.�D���O?�Tq�(" ���puk�2Oj�͘�'|~�;4l�av��	ÑF|��a�'���zsϒ�-#�$�@m��E��TB�'���,�,��( 픥I>*X��'�콱wƋ�LX��-<X^���'pd�B�s��0)�@S�~$B��'��l� 3x3:�
�R�x�pZ�'���@AԀ
��]��@�
G�q�
�'f�pC�;j�V�e�͡C��uk�'Į��Vo��]d��Iը6��1r�'�!cg����L!̩2�p�9�'.i�nA�B���K(tyԩ�'#��s%�/jqԴ��aA�����'��9ҩS7P���P�R�xY�	�'5� h�A��#y��&�ׅ.����'a@����*�~�x��/}n�U��'d��Z�@���]�?���k�'�X,Y�E h`Z',Ėf+<�'g�l�c"ڧQ\���A�,�f�+�'؄,�rLՠ,�lz��
{C�d{�'�B̪w
O�I=:��#�ĩcqŸ�'���y,P$<"E�SmĪn���'0~A7%��ze|tɢ@�Q��'U�{��=tK���QbI�"A+�'���Ae��P�X�y�n
	H��'W��(��ϚB�� �%G�3]:I��'0���!�a2 i��^�(~P��'��x!EϯY��\@���.Nt�
�'��T�Aӳ=��4�Q��Q�ث
�'ZB<�U�$bྉ�	Br���'����-N�'�F�h@韾P~B�B
�'�Rm��E\�H�h�P�a��I$��r	�'�$�`���n�tK����d�	�'� z#AI�Ma��I��B6$��E��'F�$���^<Y\���̽+|���'ִa��+p�](��I�!��R�'�A�5�*3�=s�Wy� B�'?d1j�<��=I��K���'QD��+",��ű�+I)jچ���'	2H�o�m���!U9\�m��'@�s��:�}��e@�K�'�ԼBB�W�Z9��~��1)�'U�8Y��%�ɜ	x2���'-����ٳ*�Ő�c��Z!�'�\�R	ۙG�Nq(%���jx!�'��ڋ8'&�3�f  D�	�'L읭(U�ְ �K�&� ̫�6D�z�� j@X��(��!73D��a�ń:>N��C�/�6H��a�1E2D�,�Ec�V���.�>��|�%�3D��	!�ye�S�ܸf0Hz�a1D��y��ߘ:�Y0�BN�$p@��<D�4����
T�@��T�+Aʹ�R�'D�y��JT��)�O-q��-i� 1D��Q`,�4��1A"����0D�0��Ɛ���E�v̵1�k.D�pa�XÖc&�*����-D������Y6�lڔmϊZN��A?D�� �eX�Z�D��cLVjIC�=D�|��)�*B��P�Yx���?D�0ir1��=Q��"�p�C�#D��s�aH�tY�1d��4V,���<D� 5�
�CHv�CA+B�F�Ց��'D�� ���2@
j�dTR3���xqp�)�"O��P�'
lƢ�S���h�"�"O� ��"aiQrB 0#;���"O�!+A�Q���Q��S�c"D��&"OJY#�Ƈ1I���O»U��R�"O���+V6**��2�$ab"OdܫPh��h>t��d��E��h�"O�4r��S�����I��T���"OQi2ȉ�n2�	Ua�j�t<�"O��s�L͙j"�Ep��ˠ:���`@"O^���K�@�P�@�M���U"O�������y�j���M�y�� �"OLu��n�;�4���
�ra��T"O����R6k��PBgJ�wx��� "O��g.[�{���c@�ur�`�"O�xj�0�Z���3P�9�"O���dK����j�/O��"O}A��/5�p {� ���4�;u"O�3��1k��@�-K~�u�s"O<�yN�x�77��EZe��c8!��Zo߾Ĳ �M,( h4-�1
!��Y8}T��G��m�@��,
C�!�$Y�|�x�jT&Xy�����!�dZ�\��i1��O�-,��ˊR�!��˜n"M��ѼY>��fh��e^!��&8ZW�ɝG�H�Q��TS!�ă�?1Xc3�C�4�&�B��S�.J!��D"��M[��I�ld�fB/
=!�Đ�%ļY��jLq@G�!��z��M�B��h�>\{�ċ�Qd!�䑡^�@�@� ��P�a�!��r
�c"Y�;���x��M� �!�]�k�H,dI#�n83��?G�!�DD�t����+d�dM[P�V�ny!�UC���k�5fܢ��({^!򤒶"�~�$EWyxl�y��;%6!�D�7F�p�ۢ*3�<����_q/!��4zu�x�&�U�u�ܐ`�煶p�!�dUj�Nա�i�4Uܬ%�Sg��?�!�$�-F�� � Ή���RťS�-�!�$!��q���J;f���S��r�'V�����y�2���Gŀg��C�'�xAA�ňKI���©�<[#�T;�'�T��!��bHJ�Rg�\�XJ
�'
r�@��ԬX�b,b�!S4Ym�lr	�'��@	�T��CG
U�tl��'�6,I� �1buI$h�2_=�p�'�@I
���)Ed�QaT�B"�N�1�'�6�g��;?��[�oF	�jm��'�8�����8�\�1ő�φ��'ި��`f �K���+R�H,��'*�{נO��f��P����k�'�&��p��6ļt#�e�w� �j�'�l�37�FD��0w��F��%@	�'�l���"1VͰ�����6E��#	�'޶}�MkS�L��e�9r 2�'���C�T$NN�Bɑ�.V�z�'���H.AN���C�Z~)�'��T���W�t�T���G^R��e��'V���Cl�^�nh�#�s": ��' ����v��*����h����'P�푥l5!i�|���T�M�8D��'��-)�EY#$����A�xx"T�
�' :Y�'Ԟx����
kk
Ph
��� - abZL�%��c�=2���c"Ot`1�dư	'�͗)Y/��Ȇ"Oj��&��+Tɫ�k�WD\Q��"Ok ��"ř�ʁ
4b-�5"O&̘�FH� ����C�TX�b"O�9��n 8PX8I�"#'�p  "O�y9!NB���ć��5���H�"O���띊E���zw��<8^��s"ON�"ĆP�"��#��!B/X��"OBl3oܔ%�dⶁ�e����%"O�]��I�&��I���~4��"Op�����&P�6U�WA�x��,;�"Oཱི�A!F��qcM^��Ve��"O��b��Z{��˽&��k'"O� s����R��S �
1�$"O���5�A�Q`����Ò"F��Pj"O���].T�XM�BH������"OP���h5�ٓ2-�%w(�k7"O��q�aC�Vd@\@�!u}�
Յ�@�<D+7�<��!�� 4h�"�O�~�<a�ÄZ�� ң�&�B��!K�}�<q�553�q%�<E3,�s˒e�<!��ϊw��W��R A����G�<)šW4O��mؕ˔ u���2�OB�<у��E�ZM� o!��s͂d�<�ѩQ{؆��DX"$� �c�<ЕIt����0fб�%�^�<��匝+4�g��h��}c�&�q�<�v.���<5'�
?��9�Kx�<��"xP�3"$�L��F��z�<��/p_ԙB��zơQW��v�<��j�J���Q�lԞp�&�D�[h�<	b��c\>q�h�6��{%�|�<1a�W�,".y��Ά����t�y�<�פ�.x r�I�L��!�VP�<1��+Q��"�
4��У6EYJ�<�dG5_Lx\3�#�G�i#��Qb�<�'P�=d�SC`�g(����c�<�W� 8�i�;2��T ��a�<�t ��$`x 	<"��!�g�<�׌�"~@b]4��:)�x�i�!Ba�<���,nR�1���(��!2W�M^�<I��=!�9��Js�� jE�VP�<�1aK�Nc��q�X�E�ܨ�#.O�<���Օ)A���N��9�LK�<��hO�yr�dmێ#*�ق��q�<�0&�!_��X��0z��x�̕y�<I-��{aѣU�,<�5P���r�<	'@��x��ţۦ�:�C"\m�<�bј(��
�&Z�<'r@�1hm�<A6d+�=�a��<]�!P�ă@�<�fL��N���f�8H p�lh�<���"@<4�S��57��<yU)�]�<I�a��\L];EŖ-2�H\k��D�<aRm�3 ��R��+Gd��R�%A�<�t�1l�j"�F+Tm���F'�@�<	�lL
?��u�VJ_'Xp��𶣞{�<�W��1
��R�_V�$$������:\� ����&�H !�+�Xg�l�ȓ/8F=�Ae_4����BeݷF�4�ȓ\Š����Ӝ&T�ċA�ɵKR��ȓ�|%�U@�otX�Ԭ��
ْd��2����.;l)P� K%Z���U����$ˋ&TZ��!�8�~$��S�? ~|�B`�7�Y@4��:F�y�"O�	yk g��	�7��)�.tڇ"OL�r�g�oЦ�����%��DB�"Op��@���s�M���:�"O����AR>Q�(���摼R(�)�"Olث��K�&Ʉ�5��5{[4(a"O�X"Q�
=咠Rp��&h�����"OL� 0_v����<X�B��"O��h`��Č�� 
� ���9�"O����hN!2������'�΍�%"O���j֡|���
e������7"Oơ�RoAV�Vp�NWu���@"O�tIթ�tҥQ��Sj�Ъ"O�@�m+uX:eHsc�)gl9�R"O"EI���ډB���u�rq�e"O���ǓX  @�C�%�fbw"O�A���w���6�(��4v"O�h���Z*.TȦ�		eX"O�{RL�3�|If�6Nʼ��"O�E�F:("6<cӀD/r8h!"O캃iL$?�y�5������"O�e���)��刀eM� �|���"O"�A
U�)-��r��D'�d-��"O�Ӷ�m�"��!bN*K�p��"O~h�Qg�+��c�ʟ��~ ��"O ���E$Ay`�G��9�MA"O��i�Ϝ)bb��R�-VH"�J""O����D��o��(���.5�p��P"O�M��;��KV!G9��y��"O^�[%�Ԛ~�&���!My�Q��"O�a�g��ل��P�@9pV1�"Ov����K7+\t��,�''�(`�T"O���#fC�^�����%��/��1"O���� ;�KĪ����rE"O�l��i��i"�����z��)�"On!h��yMP���^a��U"Oj��) �/	�"#(�9?,� �"O��k4��)~:�𶦃�-vc�"O�� s�Y;-2 �4喃RD��"O�m1eKP�c4�B�51��P"O�<�6f��LW��&�%lV(A�"Od�Z�ї`�!C/��:�a"O�t��o�}f�1��ğ�j� Ёu"O�i�Þ #\�TÃ�F�H� �"OX���9��Z��PN�+�!�D�@k����d�� �rH�C&�!�dIv�M�����}��d,[;P�!�$Ե	�����p �E�y!���
����F�R�A��bI7J!��D
Qê���	C���!�ۤ�!�D�$`f����+>h���^t!���6��"N�GGl<r'��^!�˘f�`(q��_)X�)�VcZ?!��<6m��p��/�j���Ò4�!���P�Ag��t��	�!F�=�!�ʶ<�0�!J����� Ł�m�!�Űu!�	h�gZ�~c��CO!�䙵<h�Q
�f�i����܆�!�d�$?���!���cTl�(N�!��N 
�h$8P�Ɋz�UX�M\�;�!�䃆*��أ @ྐ4&��>K!�4@>u�d�hk��@r���!�U"j�U��$�L��
"	L�!���.N�`���X�L���\�{�!�� �`��Hk@�x���[�Z�"O����-�q׈�:gJ�-�Ԅ�S"O^�v�̂&5�R��ͩ-���"O�\RR�OXRQ��ܧh���Kg"O>%]�?���3A�Q�/��U`�"Ob-�4��XT�y�	ڢ6�0	 "Oz��G�0"Qh6O�39ߺ�$"O���B�͛T�����n�&͎uBu"Oz������y�:ّ��'	�T�kp"OV���ͥvb�C���f�����"O�]�tZPy� ��%W!�)����$ړ����_1����{R�Ц�o��'|a|�BA�(��كE�+2�@e���y���k촄Ig�l`���B��yr��.\�*�:D��)^Jp("���;�y��/a�:� 3��Y鰄�O��y"��̐��ȀR/����H��y�.����-J@�I�?56p���S�y�b�	o�J}b��S=B?l�t���?��'�Q�g	X�`9 �l	�4���c�'� <�f�:N�҄���
'��1�'v�3��'v)��XC|I1��_�<AAIȲ6!<${%/C�9�|,[t�v�<9��11j���[�� �hS�^�<d㍘?��<+�]5�: �G�u�<�ҥ��(��E�U�ӠXr.œ��A]��0=a�FO�;�t<� ���p�˒E^�<	F*�-O�. ��� ����X�<�0#�.�������H� <ӳ�H�<I�%2z���PcgU#1�����A�<� %�(���b�c�e�n�p4"�B�<��!��/���W�b���05M~�<�u�� _ ��)��V�{ ��3�eHQ�<���'�p��c
\N�#�K�<IA��0)����&�!�1��_�<I�o$���3�V�6[ʉ^�<��oW 5�*]��_|<���@P�<���^] ,tX �Ur�6�J�RQ�<ACLQ/l�.�gD	U�����L�<Qq떷���� JQhj���f�Q�<	u���3dIat	V�Z>ʨ�`�[K�<���B4o{\;�
 �F����FA�_�<	EV�$8�����xk��]`�<q �V?�̽##f�>I���˲�f�<�@K#3��	�W!��v|@Ѳ��G�<��Κ?|~�y��óP`��hpc@�<iWBȼfXa�U�줰�^���'&a|�H�	�Ԭ�3%�wp���)�y��N�$��a _�@��Y��
��y�S"&��E�ʹ~�X�.�%�y�솴1	B
(�l��P���y"��l
�t�MO�+���7  �y­ϖr�H+��XF�{O_��y2M�	'�\���W06�{a���y��� �b�0�]�G碹�!V�y�O��U��4*x�(�w�E�y�9���7�БKr���/��yrM��M��EU�-���JY#�y�nK%ZCD���I�9BV���Mڲ�yR/ߘa�Ԁ3�l\IŲ�9��y�$6��"6%8I��U�u���y����v��X�8�"�φ:�y��3f��I�f)B�����K�y�`��{�P,��D_�C)�I[�͐�y
� $����/]dՁ!��J�I�7"O�������s�F�$=����"O�ez��B_�1����$ui��'C!�ªEA����y�JhQs)�)c�!�D�.sZ�A�B'G6lc�T��W�g�!��T�Hɱ��X�-D�H�'0�!�d�B�e� F�)����f�Q�!򄆭��q�%@�ycT�
W��9:�!�䓿)�$�0Q�[<;��%.K!�D��k��C HO"&G�9;BƊ�-i�O����$�`σ]dГaC�2A����
�'�|l�"�.c""�˰NV4(�d��
�'�lpc�^�@��D���&/Z�	�'�6�����^���Kc5��M��'7�\@ ��6�E��2�:��'�P���,_�1 i����S~��'h�#��ײ(2b1K�mҗaj���'F�<`��El�R�y�O�*���#�'Yܰw�Y6/�ꌳ&kB�'�&�
�'(遥��T(<bVBG��&U�	�'����^.v�zI���ܝ=0��2	�'���a&� :z���6֐��'�젩�ʗ"��<B#�^+;���a
�'��\p1���h��Mӳ3o�=�	�'�4�p��ck��p�L&Y(&$i	�'�jɨ�''�xaV5X
�+	�'�.%�^A��)�J��E&�5�	�'�riq/F:.�
���X�R��e�	�'(���wb��Ii�02���G�8 ��'g��*��}@��ݫC� � �'�qpc޶-�
��R�J�0l*�3��x�ѹ[����I:� y�=�y�Y0^	T��pOG���&��y�P��9��P!T�P`E(���y���jٸe�qc��{\�	ɔ���y��W(5h��r�bR0{�"�����yҤD�n:�<��:w����W,���$.����'��p@����	W� =�6A��'�z}�g	~��\3�K�'9����
�'^m#���Ńb`�2 ��!
�'��-3���l�n�HY�)�(m��'	���ʌWn�|��8;��)�'������5�[�0���iR
�'��b!˚�򀴀0�WX�Ԩ	�'��tc�'@�c�jLn��H��	�'�T�"�A>(�t�XW#�{n�Y�'�@���,�?eS*�����|�r
�'���pM�uY�f�J �d�	�'s�13,44� � B[<��'�<4�2!(#E�sB�q32�'��ʦ�O>e=(y����iCZu؎��9OvM�%�������!P̼%jW�D�Od�D�O.�$�O��'<�N$�Z�^�9�&���e"O��H5+�$�Ne�f��9�� "O��IC�4>�d�+���U)v� �"O��1��<9v����;\���"OXhx�#�tD��j�
�pz�"O&�@��ǋatPUŉ 7^����"O�lӡ�» �Xy�g�G?$u��P����ڟ��	ğ��I�\�IG����=1������F07�d�����y�.�1*<n˓爉c�h�����yB�T�w��鰆�b> x���yr� mZT����lߜ�s��+�y�mqUD�O�.b	d�C���y
� L��bX��>�`�K��rU��qq"O�=�M�<l�AK�2%�u�7�|r�'b�'�"�'�?�7#�(B�yz�kU0]Y$4kG�%D�\�d� T�h� ���B�R�$D��󰁌4�����@:g<�QE�7D��F��_��M�R�\�"�4D�p�'�֬x�T`�N�	F�֭(Ҋ7D����ߚ=9��gˆ;T�U@D)"D�t����e|�1�B'�.�ЂL ���Ox���OR���Op��4�D��Q.�dk���9�h2,��<��Ð.|�xx�k�wդ��0��p�<Q�K�`���p�N�@Y����GXj�<��"
}8FjZ��n��v	AN�<i��#�A��^: �9x�b�F�<�'Zx,�(w�܊R`*ы �	yh<y��� [�,ar���7p�
7�_����?����?	��?�����)�5�F4�5HH�B��Q�ѡQ�!���}	@���J�@���ƪI5�!�ɥ�nݸQ��2$�q�K�,V�!�d�;>gz-��d%��(��&l��'q���bF{Z\(C�K��w�p���'��*��eR��ql^�i�p���'��T���U�s��2��$B����L>����?���?9���?1ΟxQ��S9HO�u�pǞ�_�ٙ&"O�����D�K�e��c����"O���4�X�� JE�><�J��"O
5cFN֙%��8��	�.�X�!6"O��E���zP���0!��	v"OH��gB����:!M=P(B|�P"O�eQ�/~�]3�䄋$�|�'Tr�'�b�'��?	���B�|��V*K;Y�졊0�#D� �0���*~��	���?���a��!D�|��-�~�@8���9*�\%9l!D�����U�/��e��n�s��ץ�y")B*J|z���pg�M���y���M�L4�T�� �N��#@Ҩ�y����v	�,ׁq�p��թ�y�V��f�/q�pt�u�X�<�`$�#�젲CZ+g��ڠ�[A�<)t���X<p( ����/q�$��j�\z5ϊ.kX�e�eS �:4�ȓN�v #q���V���$$C���T 0�Z��4���G'$�Ԅ�F��CJ֧Bdn��g)�%��0�ȓ<&�10!�9,hI�艕B��m��-�>��S��?���ʤ"���q�ȓN�M
צT<QD�K���6s�`��R���0S �f�R ��hʎr,Єȓb����u�ݒ<����h��<�n���o_B�6ȝ�!.�!�O�o���'�џ��<�W��$��p��M����wn�ٟ������w�[1����M�^b��ȓUa�j�G��yBG(�����*R��?` �����p"Odi�"�^�b�Nu�d��dB�X�"O �r��8%��p�eK�7(�`��"O.II�"�?	2U�L=?!XD��"O6)�V��;K>�k
^�{��-+C"Oj(�K�� yEC��0�> 
"OT�[�IC.,ɐ�Y��A5[b�}Q�"O��)�΋�0a��(��utJe3�"O�aC��ܲa�A����"Ch^3�"Oℛ���G������<���{�"O>��f�-�<�&�N�f	��:"O� �B$w�� '�=(�dH� "O�8�-:�N�a��S��T"O�@��'���~�kq�9U�D` v"OHM�Ly����2K�����"O��r$��<H�xٳPn�����"O$!�a,��ED
�0���c�L��"O41��']Y>������w�\�!�"Oֹ"6��s�씫��<��B�"O�Śh
>�x]a`��tL��"O�yq�% s��:�OF�!��dp0"O�|���D�r�D�CR�ޝC)0��"ON<�$�@�j���إ0����"O�I�Fl^s�f���./uT�F"ORT���ЀQ���Y�s ��"OJ|9V��-±�glQƺ �W"O�QRq&~��p
�ʐ�g���4"Oz��E��M ,�8�ʞ/
��I!"OP�ۄ�N(���� k����"O���Q�;$qI����$���X�"Of�`�͇$g��r�:��yI�"O�C����w�\I
P"K2v,���"O�Tr�I�ZqfUϕ�L\(R�"Oč(��^-T�P
E�\SM,t��"O�8�qk8[}l BnU6=��"O*dBu��4x_�P+�R�tdS�"OU��(��rZ��0���H8�"OxT*�ŕ�K>P��'�J�O����"O©A���2#R�x����(�"�"O��P7u��Ö[�Fovha�"OX�26�	�`#p�P�LF�,A�x[B"O�����	 �\A�W�Т:��h�"O�hy��V�S4�C4�Ƌ}<�[&"Oڝ���@�`b��8x)��"O�]��!bN�Y��9r��y�a"Ob)�2���Z��K��m�l-��"O�!ie��K7<$�5�j�5y�"O��r�[)Bw�٢���4�2"O�(h���4%�H���r��,��"OƝ��L���YqN� /�n8��"ODE�$�E�O��c.�(Y��UA�"O�Y��~\�-�4A0�P�"O�M��$(T.h@!�P�
��a�p"O���!�I���;3�� MD
���"O���!�
��Ttd�B�� c"O� W��J�X��W䎽T7���"O��X�@C�w�l��Ë�<�pUz�"O"�q���)5G�2&�("��t؃"Ot)��ӊ$�NP¦�\26��4K�"O�� ֮��]�\�@��B.̄��w"O�A�4�����(8Y�v�s"O�L�@�(@�����<�R�0�"O�	�,ȿZ���J�)f��}"O��$F�8a5hѨi�,Er��"OJ�3��֒dt�����?��(�"O\P���'^5�UIc1@����"O��i�`Y<�s╶q����"O4 X$H]�\�0�K��˒ko�d�"O^֠ �-˰�x�bЯ;Y���"OPu�;Eh���|F�A#"O�%[���ǎ�@6�!I�"OVɱ ��$��2'�?%�	z�"OB��%6dB@�:<��@�"O��Y��2G�Z(�1�6����"Oj�B������F��&<R�sc"O� \T`�HS.>X҄�Va77x�V"O� b��v�@J8.+Ra`t"O:}��/?��pcB��".��F"OD8sn�3E�p�)<�:ѯW�<ђΚB����*�-ext9�Mm�<yf X�s9S���B�,�2 Q_�<I�(E�A�x��ʩj^<�H4��W�<����<� jSiN�2~����o�<)V#�p^\0o�9E"�-����a�<I���#��}�*
5 /�i3��v�<q!��T�NQc���/'�Ӵ��yr�O`d�s��áYۂ;�"�y"���|�F-#�j�=O�pS��H��y��C�|����)P�E�}i��/�yZؕ���ɄB�lڳj
9d^��	�'��A,Q�Dʲ�ѶK��e�	�'�@��!ͨ��E��'vBܓ
�'Z�zӁö^s �3VEC�ͫ"OlI)����R&���r�ޅg@z�bR"O�#l��rYqr��5:�"O������9!$�9�d�2p!"O*�qEY.r�8a�b�J*�ن"O�Y0ԧ	���#SA�)v�eH�"O:]�2Mk -�5�J	��(w"O�t3�ο)Yt�;&&3zLN��"O@���"N�/�"��R8j�9`�"O�ժC�&o���B��H��"O ��S��+~>�ys��1��̳�"O�!��t���H�OZ�nm�p"Of��.#-2iz����9����R"O�UY� ��-p�qq��,�\��"O�Px�M��SV�jԨ��&�1Q"Ob��%��V<DY�m�
u���I�"O<QHY?]C����DXNx��"O���K&Lzm��A�S�"O��v��;Ո�ô��kX�"O����(��'Q�h��kas� ��"O��"�ϙ�.tIҪC�6_�QD"ON��b&��Lx������+%t�23"O<QH�fy�Q�A[�AW&���e���y��+R��)b+H+0��y��W�y�%�%5̦1�)@0"Ӥ�	���y���M��s��ڬ�g��y�Yz��h���� �I�'�џ�y2(��pM@����Ȟ�������yB!�!�T�Z�'B��#����y����HŻ�pL�" ����yb�*�@%��T6�(�Р�Έ�ybbʎv \��ֵ~r������y�L'P��eY�lW$��>���ї"O�5(rKS'd_,�
S�	�=�(!�"O��#��	-Fȳ��S�K�����"Ob�[�D�-�A����\zB���"Ox�����k�<;�VY���kB"O�(�s��:s��K���O㖅��"ORy(t��>\�PD�c��	�8�*�"O8�cn��(�XЫBN�2kԨ�p"On �gG�hK���#@�Q`��X�"O!�#�\�[]�廗C��=�L��"O��R�j�O����ռ�͙"O��uNKK��YS@��q�R-��"O�U4�&YUȑ &OԴp�H�0�"O�E�'	�wH<���Y��(Ja"O ċ��
�o��YXvL��ݘ"O� ��q��628��rRk5@�j#"O���aG�>�ΌB�*� ���� "O�1Q��~�����(�}�"Oe�V�Ɉ��1�M�O��w"O����72�ԩC���B�p���"O� dd�b�|1��x�xA��'.�੡f��9��Q�U�O����'�D�s�jIwC���ț�C(*���'^0�@A_�QJ�m�#ى>�q��'8���T�s��`���"Lh�C�'v��; �T>g���捻����'Tj�bR"ǽ���肢M=S"�(�'4x��"��13��9�'��D���'ܒ���N4�f��Ү�,�X��'��!�l)��}T��	�'�^��s@׿��P����1G�I�
�'��9��?u(0�DR1��'jp��1I_:���$c�x1L���'-� 0�	� ����&/U�pp��Y�'���Q���#�!���1#N���"O��b�gO%l��� F��/��3�"O��P��T��=��g �},�!"O���Q��&p�`x2r�R;Q�i��"O�Mc�	�Usn=0o߉6�P�`S"O�d�T�[Ot��d��4��ڳ"O��p!��2o8��
A悪!�4P�"Oܰ;q�B�l{6aq�E^�T�c�"Oh��HJ�}�J4�&�לM�Hِ"O4=kË?�$%�'��5�:�5"O�0�)[�4�<�&Lɐ{=Z��%"OT!@����u:lJr��w6&�YP"O�(R��<G�=��$/���F"Ovx*�#�/c��`p+M�2n�"ON�[��%�*(�Ϗ�;���ۖ"O �P�"^�D�酥B��D�t"Ov������(��2��aE��V"O@�ٱ
P:k�YY�*D;�l8Q"O��#�eI[t])3�Ȧo�vMzD"O�L�0(Ԡ�z��	IX��2"Opi�Qf�.W`�m�� Ut����"O>�+����	���#�a�"O�9$����h��D�eX�]3�"O����(�,p$у�¿QKFtcd"O�`G锗&�I˵M�ZIp!˒"O0�H�Ұ!Yr�� �
�=4n�F"O��I�BL'm*f9 bKW��T"O�9����Uy�q����&
�x�"Oz��� _�zg�<�BoЩc���k�"On �V�<���ӳgP��tq��"O�蹔h# i��'��X�$�(#"O���(VGjV`�oԐ �hD��"O9#�r���P�n�nU�ib�"O�=��d���DB��֙L�rs"O��P�T��)���+,*�)r"O��qP��*b��@@v�H�T��`��"O愰'EE�06f,QĮ'��`�"OB�Iw�)5��B@�H;@�^��"Of1I��P�'�P���v�|i8�"O�r�L��|��x����:crn��6"O�h��ʄ5�01���:I_�y�"O�L����<��P�BLA�XG���"O�m��Q�����%�653��y1"O�M��ݏS,�T��0A!��"On�����rGD krn�>u�� �"O� $qC�I��}���ږo r>|�2"O��aI�T{�hҒ��K�&�#"OtmY�U4�<��ؒ9���y�"O��$��y� d�7�
�^� ���"O^�٦`�1%:@���JߦȚ�"ONܠ�O�v6����S?K�Dq�"O������(����U�{���8 "O�QK��1�n]q����D��"On!�E��@m����B=�"O��q*�'"8f%8J�
J��
 "O�Pc㪙-*S���$��#)�F"O���`
Sd��XP�R�,�Lĳ"O�ħ؏c'�y�@��>}B*�+T"O��G��F��%,1iHX�眬�y2���J�8�&o�n<:��Q"�y�I�_��[g�!l��ջ���y��)Tq��E:�V��A��y��H�~9��"��",��`�JV��y"+�>�P��T�*g�X�@�^��y���5T���c�J""��(wiB��y�/�|G�y�B�K��-Z<�y2,�
#)	��?��1�VDǛ�y�À5��Q��ؠG�|u:S�д�y�R�N�*hkc�	�I�
i���yB�?h�@�!È�@T{�	D5�y��R�	�ց)��V�f�z�S&�D�y�kB`���\�/��2Ɲ,�y�h�2�!3�g� z"�)��W.�y"���n�x���.s�,��q%��y2�%l��v���m����P���ybF�Md�L E-׮[)�ف��y�*�CT�#Q��aĜ�
1jɸ�y�/M�Ru�Y�W���`��ya�(��1h�z�>3������^�z0�؆�%���I@W]8Zs̆�b��<��[��@#�,]d!���:N�\��ȓO�tX�$��J���b�d�4['���ȓS���D"E�F����Vc�+$P����~� MU�+A�5�,��-Ĵ���qd�I���H�
+��SC�ݪd�ʝ��)�������(�:ܓ���Y�^M��x]RP�R�_`d�3��[=�Ѕȓ���g�՟Y-$��`	?VO܀�ȓfx *$,��$(��� 8᪁��1�^R��V-��0[%m��rȆȓ���IBޯ~�P�%�R|���ȓt���)G�^��� 8S��,|�f�ȓc���eLŴ)���r��Q.L���#����e�W_ްqE^�@X��<T�-�%W�*,�Q�	�'0߶i�ȓyJ<IG'C"N�����8�ȓ.�0ׁ�5W'~豬�d�L�ȓpȈ���ݮO�0��$ ڔ.TlՇȓW�^8#��;�I*��	p�>��ȓp�E(Wcň"o�!�bG�t������
a��� y���9�K�w�R��ȓ*���I��W���A�{�f�9D���!O�	L�-ˆJ�y.��06D��kUk�%*�ٓ��"MR�r�3D�s�nYJ��0زI7h�Wo%D��s���UF�h�E��ґ�-D�[ʋ�`�fĊը��Ӝ�P��9D��Q�ƃ�n9L9���1`Ә� �8D��������y3�, �e�aD*D�� ��r���+Y�8�0�� -�p�js"Ox�����)t�̕�d�Us׶XD"OB�
͢u�6�1�^�d"b"O	����OH���Y�Ă�"O�*�n9N��P��U��|�R"O,�b���5��uj�A��S� �"O�4zbk
�&]�T�`����"Opj�.�O��X*U��4�~@��"O 2�'��]O��9�iƎy��X�""O}4&��DP�$"4c�!%b�9"O�����)h[� ���Ň$��"O1�%�\9�vݪ��;?�@�v"O9(6�MuR�������&"O��8��&|����CE �6�꤀�"O� ��NV�j�H�CR�Ytb�q�"O����\��t���A��aY "Ot��em�	^�)0���H	Z�"O�ͳ�B��v욇b�>:R9yp"O��J�&G?\\�{� @ 21��"O����؉$��F��Q4nš1"OV�a��1�R�Z3��#O~xs"O�����(���#F�/7~h0"Oꠘ�ǿ!��S��3y4H��"O"��!�ǜ`(}Z��?b�@y��"O�(8�
J�
�����T�Pĥ�"O��#s��s�"\)��	�d��"O�p�Т�bk|9"(�H��h "O4�ѱ�ι*w��#wg�>7�	R�"O�}��狫1r�hh�K�� ��"O0�LA��n���_�:�jV"O m�2��;�ܡ�&
�9\�=a�"O���l�"�4�dϽO�va �"OZ�0�٦6Hj�ru�]�7�V%YT"O
�b�:�"!�@�X<f���0"O��[v��J���9�0-��"O\Q���	�d\Ȃk�:_�F�(G"O����՞��|��G�t���"O����bϪ7�F��J�$&����A"Oz���*�Ti�`��0B0�)W"O\D�ᯜ�#L��)�1c����"ON��"�^���0#���0Xt�AG"Or�y&�j�PZԡ�_��"Op���AƏO@�q׉�%:��e�'"OD`5d�j)2���$K�p$"O�p(�t�E�$�=��p"O�)�b��	0��×"Ԫ	z�P�"O̩�D�
6-�sSaWb".���"O��`��ٿM��5y�O�Dr��r"O�h��I���\)֡o����"O��r������V�G%UR����"O�l��X�
đ"��$7����"OX5*��֦v����g�;%�}�"Oh���.B�`�\)���J�E|�� "Ob!��E.l1�K�Ay�!��"Od����WWv��Y�h0�(%"O�)��M�p%*A�7�ɩ��;""O��yE�I4{�h@a��]�jpg"O���A��H	da��<s�j��t"On� W�
�U4��Zu����t��"O��1�D���y�7��_���3"O��V���=��M�&�2P����"O�ȣ�
���T@`��q<�F"O�� @���I�&l#k2y�""O�4�2�� >�<LI�J�4)a�EC�"O� ������`LD:4��`�IP"O��vN��D0�w�O��X�
C"O���Vl],�&����T�bդ)�D"O4D����ܙ�ӧ��x@�"OP�d$�%¤qA�B=z.%(�"Opm���C,h�����dM6z�hrp"O\`9C��'O<�;fC"���qD"OP��!�F��8t�7`G	roe*p"Ob�K���p��a�s��ɼ=õ"O�p�F��v!3⇒O�z=�R"O6�Z׊�m舼5a2&yz4��"OZ���j�y
�X�Ѩ����"O4�����Xq�c��m��A`�"O��a���p���CU�"VA� "O~� ���Y[�P�¢Y)A���"6"O`k%�6�\�r�^�A|Ƹ�""O�dK�fغ��=ӡ�!M�Y�B"O�!hqĕ&��£`҅1� ��"OH�q��;���ӎL�e���kd"Oh����	�P�`�<L��@�"Oj@�CM߅D}�w�ȁ+��4"OPa� @=9"Na{�ΐ��ѹ5"O�e�S���V��(�P�.� a��"OR�Sa���vQ&�ۗ兩C+�1z1"OzEY�LX�E�����A�����"ON�:`�Y�5��ջV�F�"O���EޥM�x[�-G����b"O�xcq�ˏ8ِt[ cΒP�lы�"O����g�''7N$bBƠH� 4#g"O�Px4có$dh��f�|��`�"O�|�ag� ��\�1�\�S�"O 3�∳/�l=X�
ӵeF%�$"O���u$��5��si�5UHa�D"OX�i��!"z�U0�,6�$�� "O4�����3l{^	�s
��E�9Җ"OΤ۲l_�`��#	A�Ro����"O�I�.�'��j�蜆�� �"OrJ��"��
3H�.QZ�"O��%�xT8IE�,Z�e!�"O��C��	3b��D��jҢ$q
���"O���"�,'4@QƩ¿Z]@�"O8�Sa�BD�l��.�?Y��4K�"O�e����8s����+�(C����"OȐ�G�''�F�7��?��9�`"O"1�FP�nh��b�F�B�"Oz8a�L*�n�" b��L�jW"O����`F\�i[b��O{�Y:d"OLiaR������}pl��"Od�aÇ-Y,�x&�::ilQh�"OJ *� �;H"�)����#TBP��"O쵈%DC�_��a!�Q,@�NX*C"OҘ���4����(Z�^BD "O�4ь�<`�0�g��L.��"O��Iaę�{d~�05&K�%��ڇ"O�i�$�-s��A����/|Г"Oе��k��|B�Y �P�Y u�"ONP�R�T�)�BՁB5*��:�"O��BR��$�:\CS�	����"O�Pj�X�%=`��Aߥ�NY�"O>1�s�D�
F�x�e �#{|��w"Oΐ�#Ulġ`���'`�%��"Oz  V E<L����6O�0KU���"Ou`��P#H��:����X=@�W"O�u�NX�=X|��P�D�$nXs�"O� J����V��hY�4��1"O@�g�[�@�vh2�ē+��;1"O��0O�̑S��=͎�"O��9R+�-R����e��@�F���"O�a�҈<U�)Q����)�"O�I8����I[t8�0�䍲v"OB��g�3$_"�:Ƣ�9W�L�"O��zw�ΊPˮb˟���x��"O�q����/�V���X(5�pQ�$"OR�P�� �a�r�b�v��"O6����@�^(����[X�1Z1"OI �'G4�V��|F�h"O����IH"8�TL�Ag�wP��!�"O����NЫ6� ��&�3]f��"OR��A���`����_�z��4�"O�4���ߨA�R�pw$
+�¬ d"O.�hC@�VƲȨ2ɇ;��6"Oؙ31�L<Wt��I�MY�X���"Oꨱ��L4�*=a7zؔ��E"O(D�B�G��Uf�u��0�"O�h�w�[����� �I:䬸G"O�����tK��s��+\3tQr�"O*%��+�1(D�JP�D{���"O���o�"��l�aE��&"O����/�5$�D�#l�P$�L "O�|��P�j��q+%	�D
��'"O��H�+=�!�bK�`�*p"Ol��u�ѱzPDժ̛=i���"O���"��#Ħl2�jC�5��xI�"O�pP���q���hK�|JL��"O"�B���P�
��#��j�l���"O�� ��װHWv��"��H�&�y�"OZ��T�(g��ĳ�d�<�h��"O�XRd��>�0�s�;Ȅ�["O�q�r���0f�̚��H�QerȂ"O���E�X�W��8�柃[
$J "O9P�_J�@�Z���,@�-�"O�Y���'p�iZ�,��g�.;�!�d�Ms��;S���6J���e�C�Yu!��'@PIfCY�6����2FO�5i!�ֆ�qbV�1��� Ug�Y !��V#x��-����~���E�b�!��E�09���-vF����ɑ!��R�}ʝ3��Z[��0��H!���X��e����gp��)���P�!�$Zy�9@g�P� �,�"/K�{�!�';�8l���56�t����!�DS�a�F��ޞc؊9�����Lr!�)S���aI-s��,r"oӎF�!�䌃$+��CУ߱E�B)�T�U"�!���O�>��E,{T��9��X%�!�$�A��{'�'YH.��!
�B�!�$�({�r���.H0Һ��p%��!���;#��Kv�E���p��-!�$D{��$Q�ǀ4	Ÿ��a� !�!�D��]�Qp�G�[����bG0S!�U=&�Nkׂ��y� �!DD!�$�i���qR�+N�8	�@�a$!�DN�g9
��Vi��jq��'�!�dh*�����z�D,a%/��c�!��R��\�̉0 "��d�k�!�$�f�X�P���5c5�|�T��%�!�7!{�!ɯ'44�V��7�!�]	~�|ى1n�<x@~�)#B��!�� z\����s�S>D����"O����,�w�d�
wn�(����"O����C`F
�렇%��P9�"O��2����]h� ƹ�Ф�"O���@
=x���C�
�^g^��B"O�(Z�̟>K�v{bD-r�\�f"O��i�5\����͇b�\�xq"O' �,T�tT��6��5j$"O~9�� @�
z��S�"�xA"O���
�ii�r���-����&"OH*uGR���<%�9i��s"O<h S�SV�H,�¨	�� q�"O����"o��=��I�(��tqG"O���H��LQveR�JU�`wNU�"O���3n��#>�P��[�o:�	�"O�D��C *B��[VĜR:���d"O��K���&�	ғ"^�Y5@�13"O%��(ğw�E���)����"O���F�?���� Z0}���F"OȄ�Y�fU��S��AKg"O��Q5@\�A�ܜ8�$�r�\��"O�]
GI��8��`�*�;B�"O>|Z���/F��9ei�7~Ӥ��"Op}S��]ULH�r�^'[&��A"Oʕ��B� ˂	�"�$�&"OD��gk�v�ީ3sV��48{%"O���'�;R�Y�A��\�04K�"O6l�1DB!��1��E��'��I�6"O�P ���R�8�q$	�2x�"O����0�M��D@ {�Ҩ��"O4,Aw�ӿA>L
�ep��s�"O̐x0'��Z%��q$�<�@١"O����2MX��7B>$���"OĘ�C)��q]���¨�\B"Oj���nt�<���JHXh�"O(�Tٲu����AV�&:���"O���$`\]{��CO� �u)2"O�܀����Uъ|���pu���"O�k ��dx5���j�5b"O�3r��9o �]xB�W,��b"O�0K�l�1do�(Ksᑩu	Π��"OH܁cb[�
b�y�`��L��)��"O,��@�n�>h3g���(���"O�$����^��ȡ�m�8B�ܽ��"O��#��	#���C��
0"i�F"O�q��*,@8<ZQ�#�D��"O*̉w��)�H-�J���"O$J���1Q���5"�E�Fu�x"[���<�~:��=����  �L������f�<�RB�z m�1�ֱ/��M+$g�_�<�U*� "��僑�����)V�<I�a��.lL��ǉ+��d+��U�<����*�da׋�0�"��4��T�<i'@�3]Z���Mv>�Ä�=T��i6��[5qՉ�c�v�a_<!���6P�U����*|�.��R��\#!��ԧu���
t�E����vAW"U!��_5g��AwH�=zL;��?!��'z��h[��/v���Wk�!��F��	ےEX���;v���!�䂂;�<Q�AGت�~x�IPA�!�$�4k�����ȱn�NE��GV�s�!�$�4h����I�F��`8����!��Q��%/�,ovT�s�&0�l���� ��2D��T��=�e)D(H�J}(C�'���>z�1�� �)���@��W�X0		�'�d��_?�~0)��$VP
xˋ{��O
�}��hl� 3FY�pGLtZ�耠*� ��P}.�YыP�KZH �Q!�3��9�ȓYz&ؐpJX�x�%�`k�+Jޔ��Vmb1��nä!�p�҃J�T�ȓ���ڑ	�M�s�ܮ"�X���`�&� �	+d�I��͒�@�ȓ��d��a�z��uB�5Kb.]��	\�$� ^�2e���.�ahQ,ãJ1!�D��$��r�/����7��}-!�d��z^���3�[8L���B�N�}Ҝ��%�S)pTL���#�Ch!C�#%D�h*F�[�~tp�'m�`���%D�T���68��2&Ԁ�VQ���a��Cተ|	�Eb�^�*���KmҪwTB�I5I��L�6�/.nڵY@��8�C䉪CT�P��͡L�f��D��/N"C�	�r<� ��4wL	6��<D��B䉏!BB퉆��~��y`ELWMU�6M'�S��M�AKJ*W�B�b���S^L�2�
XQ�<9\�J�R+	�4)�$2���N�<���o�����ƍ6_�f��fMJ�<�u�v�� 1�P5�
�@�G�<Q��M\�[�"�u��Y�Oj�<��,�
�T���^�̤0/M��D�<	 o�q\ƕi& Q�Z
��T�ğ �!��Z����y�k��3ؼ͢S��~�|b��L��Θ�>m���YQ�TY�L>�yB��8ZT\J���;���hc�.�y�
4^XA�  �2�6 ����y�ă�	6�M�0 ���d�8�y�LE&rB�h5�W�(�Aw��y2툀x�:�
���J{ m�G
��y" <uh�aqf�F1�%�v@���y���`�<�F��'0t8���;�y�N �9�&���Φ3�� ���D�yǘcѶ9���Y:[}�5	pgݖ�y�N�L�\��C܇W�j�Sp�Y��yB
�,��a�‴M���Ԍ��yR�@��`�`E�(1WI��ʜ��y�E��8�T��2���<8
��#���y�D�5n5ڸ`�&԰�����	�y"���<�PĒ7S�>�˲�?�yҠ�1$FƄ���H�Qаn��yB�Y�L�}:��&)�[� ���y��"ytPU�ui��4���N��y�Ŝ?{c���ce����צ_��yrG:A���"�K��~����F�V�yCs�Z�2@,��I�M+�ʖ�y2
�(�X4`��2tT8�'��y��ϡ�����$1��*�@���yr�b�JuX�!1�6�*Ѡ�#�y��]92��b4����q�W�y������
0� �J4�u���y¨	�r٦9*��J�fW,"r��ybE��]K��;Y{hi�A��7�ybG�O�䀀�H}� �����yB��{�� S�����BN��yb�H�&x.Y�S��p
�)K����yR��O�4��bM�l��Iz��H�y���9"�p�6`��+�%���y�c��A^��i��F�nT��;U�8�y
� ���5,�9j�k�̧I��a��"O ��f�5�� �S�����y�*O��Thö��t#�悅/�����'=8�*q�R?UUD�rN_%�H�'�jy�g)���䂫!���a�'�Z�[uJ�)� #�-��=�x �'.��q�*�: �%�^)~�����'���@#�ܦk^��^4^y�UI�'�Z�Rf.�8U&�)�����	��m�,)S��F,'Mb��"%�]<h���&�P��=F�A���۴D�]�ȓ`�Ī���9���+�Ă:E�5�ȓ��l�7�Ĉ~J2 [���m�؁�ȓ.�L� F$*h��I**���l��xp���`��@[�K�#���ȓ��u�
3Ԃ�ʴ��#N:؇ȓ.�d��2��?3�lIu��*I70��ȓC�t��Q�K�8t�*��.t��)��L�d��$N��أ���(y�r��ȓQp�+v��,k(L�b@
��{jV��ȓA=:d���-	b�N��T�Q�ȓQB��Xw��O0B\ф�O"$a�ȓV9�Aɓ��

��m�Q>B���(�P�:�.�F��Ԓ6	�F�Ą�t��a`���0xAf�츄ȓO�����Z5y4��q|,��ȓ����0/�IkJ�pȞ�9�n���s|e���<$�M��@�/���ȓ &q��ۣo^zc��.P9�ȓrX<�R̟�~`���	�7��]�D0�Νx��]b�FF.^#����*@��"�)�hJ��֬8K���ȓ,f~Y[#�J�洁�Ș�8�PU��ZY P����9c��7��i�ȓ2,����[%(h��f�`����ȓ���H��oa")76�LH�ň�b�<y�E6]�\���6 J���5�Y�<)�N��!R��7��봁�y�<�7�� C�6�X  V�L3e�&�<�2J��U0�+E��0^�R2I�d�<q"�	�N��,Ђ.Uе��x�<���A*��	ֵ�k=l*�)P�<�d�L
~��S�3t�z�)4��g�<预>N�	��C��$)LYdI�o�<��'V�!���"�b�)#\����j�<A��ڭ-Q�`����N0�!�a���<ag��;zv�3�49�xG�J�<A�D�2{[�y��؎'Ȥ��Bi�w�<�v��w�`��a5�IS���N�<�DQl D%�B8D��P�`n�M�<93���!��4d�ƈ����m�<	f����Y�)S�y �K��f�<�u��� I�����+:?j��ˍx�<����
���0E��n��Wn��<A�X8h*� iOs�a�T��|�<� Q�uq2JU=f^zc�A�<)�`�Q��Uqv���V� �/�s�<9�X�-S�4���*9
�90oMr�<Aҹr�y�&�X�X0ţ�7B�!�ʌ*�q�b�U�d�^в��<�!�$��p�N��@���Nۈ@�W�-:�!�$	.]�x�φ���AA��S��!� *w�d�R�OM>Ӏ�y�AL��!�Ԡ��=��
�^z��GK�!�� n䈱n��HX��ޙ+m��S�"O��Y'J�)]*���
�3�.	��"O�0���Xl�����B84P���"O�)ɣ�ML��w�:Tm:�"O򬹣c�_�3�˛�~���"O((�"�FK�f��l��g� B3"O$L�3G\��y�-ͷj؎=ʗ"O�\��I?&���*V�T�U�� �"O���"���J��8&U�"O6��6ͣ�FL��it��"O*a2�R-(o|u�R�H 3��833"Of�N�/\�QG��
����"Ot�xv�H�ue��`@ǟ�%n*虧"Oj�����%jlX���W��,�f"O�-9r�=<���Aɐ�L�ݻT"O�ᯔ�s��Mh�ِ7A8]5�'�8�;s�	'�����]�xk�8��BӋ5Z
�P���O�8Ei�'���s�E�
����u\d
�'�vmHEoɈl�Xq8GFZ�ZP
�'~�)U�oCb���!�]�I��'I�%2��A� �~�R�3Qǒ(J�'L*b�P1���ɂL	J�����'i���E��Z�B�G:9��ݹ�'s\��� /=����-V�>��%��'���7�z��{��ܲ�����'�ʍ�pk�m������ $�z�H�'p,�Cr���]s�Y�q$�
�"O���P�bӆ0�懘
�m� "O$ݒ���V�z�h�f��5���´"O��KC���]�M!'\�*M���"OH )#$�
e ����E��(�>M��"OH��ʅ�_�*��v$�2t�R�"O�����ˈ{�ڰ�W��3]�H@:1"O6!�eF�1����@�ʽO��6. D�����R= <��"n	��HU+�$<D�d�4��wPb�	�P�K�=��;D��y҃�@���`
L�V�@�B7D����1^���d��(c�x��j#D������:'��11��7/�F�{�!D�8�Ba�z��Ĉd8s=Ne�r� D��A��8)tx����~���/=D�t��B���81��.T�}��@(�f>D�lY�ĄlʴuC/!TɈ��"J!D���t`�5a8UDK�MT��p�(D���E��,����j�a�h0� 3D���G��pڑ�B,�%C��g/D���F�Xr���([�EveI%A!D���!�D��H9bd� ׌�V�>D�4:j�px��@1�[$ y
�!� =D��vN��$�P����E,u�2 �� ;D���	F�"Y@�8���7&��c
8D���Gɿ�	h�e,V���SI*D�H�� ٬:� Y�8B ��jp�/D�ؚ�e��^2n�����&M]��3%,D���#b\0��Ĺ�"ڱlC��d� D���&BؖS�Y;�/č%yHA8�a3D��sH[0|��C�j��}�:�Qr�7D���iϽ|�J�����1)<��Ǫ3D�@��B[�a���&S*RT�$2D��t�@�:\�k����qz�Ƞ�1D�(k�C&�<4h1嗌f���'."���d����j�v�b�eBި�ڵ�J��,�<ѕ�ʈ��].q��K�?aI ͘�^8��J��� i8��V䌿�ƹ���Mm(<I��B�<W�IfᕸH0��$o\9v*�����Q���Ȧ{���kP��(��<��j���d����� 2��A>����!�Z#/T0lpO�)k���H9cG��m[n4�L�f��=rѬ�25|����F�m�Z�C��Ӟ�b&�Oڲ�X�O��%K�"ӪtC��� K$����'G�M�&J��@t�	�3�t� E���]��1h�*��By8 �Ҡ�W��`�u�i^y��N�EY�����",N� 9�yh'��k�h XrM�,8�OX�xd�_~����0�M��N�ם���!��B�R� 5$\�-��"Ц��l��
uӀ��*O���WcM�U�f�
���ѨZ�Vx�'�T�(l��a%*rK���)�OHѳ2A�*Yr�RG�Q(X�BH�爕=*d��aE��M�1La���B&Ɩ4�ȳ�k���P��&ʈ,`j|i �I<z�t��$�S؀��򩊐izd�#��S�?��	9u�I�)���W<w�:)�C���M�1�Ҕ"����7�'Ev,q[2
Z��꤉r�-	�4X��	���T��`X�ز@L_�P�R4�'��ɒl�H%6��*�{5���c�A1;˛6iE�WB���5}L90v�ػ�Np`Yw�|ɛ���P	���NC�W���P��JC��3���Sհ�%�Xs7��
<��us��'�m*3�4u2��S67�u��'�����OzW���3�R�~5nD���+���w%^(:�"����G���"!��'7���1%X�RLb�W:33"����~�"I�؍y����?݈2I�,B+,�4�ܚ����X(� �E���D�y�!ӭ�rt���Y��ad)�U4Ն�	=^����N�� m33�!5!F���<��	�{��y��_�b��yH�B��W������Q�&��V�R�;����d��wU�a�W��%',C�I�0���f�_�et��z/ѫQ���Z��^�or��CG�s��ju���5��&��jWҼ�Wc؊{�A�E�M�p��q ���w�<�u�ʹ[H���t!{�0���Z/[봼�E$�I����O�����e���XO���$aK������"
Q�F��c�+���	�So����E=�~d34�	e���U�E p�<���-g� �@O,ZkD(R�+S;���$�&1,�Y`o�n����
aj�e����d��vX|0#��S���G��5H�ص9�%�20�8�iA�S1�܈ ��Q��M;��|�ayZ�p��͋f�O8sAbʹOQ"�)k�8#�.�ŭԁt+�d����� ����3Y�V9��̷IU*�1��<�t��S܅pcmS�Q����?|L~�Pb�U�.ߺO���$�*S[�}��U����oIH.��۷
$��"˝7i.,xᓣF(�,M"U��3.��I��BB8;f6-^%K��0fֺl�Dh�b��	Q�'�<+��r4CÎ8ɼ�b�@�`X�S 5; ��L�(S�4�H�t> ��i�A+EJ�f�l�ƯO�K9:%*ED�cV���lb����4�R QBNA F�'���9��P�	�D�C�	M��H�#��%��)��4��hɔ�	&};��mڢd6�aF�-�j��O��>.�&�
(o�)c0L��j,��a]��<A��(I*�pʡC�O�D9#�39j���.�v ��ze��8�8pc�F��M���D�[�x��2���nnؠ�'�Nԛ5J��*t�Y�f ͈����8���Z��H<�@�_���HV�?)���-|"��'of�!��A�aH�U#3`͠>�h
E�߂X6|�s 	�52���!�?�E�G>��I M�?�l
�{R,�^�2)�F��&�nݸ���3�"d���'�!�׏=}ưkSl��]�*�� ��uWcΞ3�^c���	tC_?�V,dV�(d�mP��A4���S��@Cd��� 3�����߾|�)��ɭA�|1#�
I���;Q�Q�'Ӑ�:�� �6��l>!�js[�X���F2O�xfH�YFr��pÉ�QخE���'Gv�� c��P��䛀2��.�=Y{R�Y!��.	&� �Ё�(������B�0��T 1GX�|�f��.,Ѹ�bfh29Hg�f̓fj61XG�<�d��6���M�&s��!�2ĸ#*�*C�yz������[�P!�VI�4�ڒ�:z}L�E���%h^���~r�B��U%�@�0fȢ5mM�*a!���P|�ᒒ!��P�)��؎-S!�G=@U��HS,��;<e*���23!�$�I��h teňo�$m�G�|9!��_9�y����/*�(�AE�'!���k��%R��u��s3DT	o!��@�Z���� �0I"����!�Y�α+�������ɲTp!��3W�R�R2nL�#d�@X��	_h!�
k*H豴�Ք8L;r���!�DKH�D���{j�yr*[p!��""*� ����4X�{�jE *�!�D+F'��s�O�� �n�k2)V#!��
0���7�T�p�~"C���<�!�$�#^��
B��
���BӢ��!�D�FV��2�*D=M0�,�g�v6!��:Jv���-?ZXV�gr!���-!�
Hi����2���3"O�]pf��34���R���2�"Ov�rʋdѺ�x	y�l��"O6e�%~4B��_,+$I"O��1��U��i{��e�Ð"O� VȂU���U����*['`~�d��"O�D�u�7|�TY� _�FSFq�"O�P���\�� {%�3?E<e�a"O��X�IT-�����^2����"O,,�q��I&�LzdK��\��"OP���!Y�3�V�B#�$B��q;�"O�h��	**���G�9�"OT����V-s�hu�eO�  Ny��"O�
Mn�B4cđ��QSS/D;m!�6R;E�aGK�n��pS1��"r!�d�
���sӴ�,��m!��֏|Ӽ�X ��K�j4���3�!��Q�~Y8�v �d�"̺��6-j!�R0|-�$�R&�?�@�IvÀ�MI!��?�����I�E#�ɹ��H�B�!���Cl��C�g,
`Y��S�!򄛥fqH��]:)�5�h �!�Da�>�AECޛhͰ��!�!��P2)��h�oΥ�t�?y�!�
�I�a1�Ŋ�^<|ò��(�!�$H�{���`�܀1����ߑZ�!�+R���T��,5n��Bo�v�!��U<9�X��934��3��)�!�D�#��HH���W� uar��/�!��H�z���S�X5�����!�D��:nH�f��	r`���
{�!�ߕ�A�.�?�Z����M�!����.�����ȋ-}�!�G�/��@�`�ɨo�葹�i"�!�?^�B��̈)Ƙ�XRS�|�!��o�:H���L�=/���>+!�ڟa�1��EԪ,�QTo!�!��G3p�~�!��1X�5т�9@c!� �����6_������-x!�dL�+�)�O���w#C�$X!��8&Y��0$��-���V���!�"&(r����S
zM��^~'!�DY�qF��c�˅$����!� !��WsA��
�*��m t��P!B��!�D "H9j�Łub��s�� �!�]�RC�8�ₓ�n�f̓���Z�!�d�.�M�%Aڎ\�5�SC[ t�!�,8�ғÀ!�
�g�
�!�D� ���;P�:/��2A`��L�!�d��yE� ��j�[���+5Y*G�!��n�`i0���Rժ��KV�R�!�X=S�M��M1?�-�6KB={�!�$E�y&꨸��O���h�2�PyB�TL"=C� >BV�ƙ:�y"�|����ƥ��GPr�Bӭƻ�yrH̅c�AK[E�0�놋&#�B�I#iL a#��T@�V	x�A�n�B��e�v���i�8�>}��KzB�5+�paAɛ��ԔC3	��@� B�RƜ�B@Z;~��S�`L8,�DC䉴n�����.��AI4` @�M�-j^C�ɱ:1*s'H�l�v�'�K�
$C�Ɉ7zʼ��ɛ�|�8l@C�8��c�HȮuC��`�呲BZC�ɡX���9u�
1H:HL��o��C䉯0�v|���J:�9��׵)�*B�� &8�<�'ꖌ= �9G�Q�ErB�IFb��r3�N���WHȑ/�JB�ɝզ�A� #��9�A�?�
B�)� ����@Ur%���̴<����0"O@0�bM��$�
�s��� ���"OX$���S\��(!�>*��R"O�� O�H�))6m�Bjl3d"OP�X %�C���c��r&؄�`"O؝ŉ�%+���,
�^�^t�"ODp"S
��&�%�*�L��A"O^���Ĝ�)��`i^4K�)�*O�DYEl��9H�4��A�#�'�pp��j,u��s�e�B%�
�'͔��iƜTJ��K<XLj�
�'�:<B��]�\�H���#�^9�m�	�'�X3g	?�B- v Q���	�'�vM[�/Ir�|u��O�U�x)3�'a�勱�� ?²УጘO,�[�'�J	�炱@�D��2��>;���'�}3�aƱj�zX��>+*�z�'�܉��,TMJT���P�]��'���eZ'8"I�MŪP<\K
�'����� ��l��૛?O- �a
�'q}1&��{zH��Èx�@0�'����quN@���w� !�'�=���ݼyk�,�2 \�[���'@~���^�h�D� ��Ӑ���'�\�����m�n sb�i�T�R
�'Ԙ@ �V�&w��ZscO f4�@	�'s��h0�
*q|y겈@Q<lAA	�'�n=WdC�jFP���H�4J�Jq��'=��y����Z�,�.C�0�0	�'�m��'��(r`�Z4(>4���'D�-�Ӣ�a3\)@��ҀY���h�'�0�����m�Ri�!.��_A01��'J������P�:��1ꃢQ��x+�'8x}��J�'�<a@�D�Kh�@	�'/�i�9��]��ܘ~l�iZ�+&D�Pa�"��/TY�P�4Q�Y���$D�xp!(�s�|���Y�f�HL�e.D�pz�̔4"�	Y�│+� Kw�0D���A�RFz4�;V�1Z!�$D�h�R	����:tדC�hU��n/D���&��]�9�Vi�;e�^��� +D�h��Ǒ�#��L{��F�{	<��u�&D��a\&8�U�uH��ux���'D� ذ�޾_�D�8s���4��D���"D�|$FDH��
Q"Z��<0�i#D�`�Ƕ��;��qqn���'4D��3$E�jf%+r��7iC�2D�$�M��X�`\Hd�?�aðG-D�0r�@�yۮ e��nUu+��+D����$Q ?˦	�@	M�X!�,QÄ:D�\�4�F��<)��	F:�<���8D�8��S<\G҉���a�O6D�THF���*�Ĺk$ R.PB<X3��+D�dY�_+yy�LX/ 7Ԣ�6A4D������<� ��#��"~NH��.5D�����Cl~�x�9^�p�9�7D�h
'�/;���%N�8BryW�5D�xi�)�=]�t�)@(�4YJp12D�8x��E#F��!5(�*C��@1�<D���1H� ���j׸C3�ŊL8D�|H$Wz�@�A�&׈��d�*D�T8!
]��r��L�*K��W�>D�|i�ІPt�(��<a5!{e?D�8���_H�8钖��(���"6�+D�� ����=iSLD�3a��"��H$�|"!�#�����	96H|sV�0Z�Fʔ�"c�4J�J�
��	9F
T�؟.M�pgF|1b��U�i�MQ�ƫ��)��1���q*�2�n���� 4�� ��î���(d���ٟZ|�(� �j�B�Bv�O}����� �����!hF�-{ȃ�qP� !O�1�qI5dGT0����#w�9r�>#�H{6d2h$jyr2�� 0r���iӂ�p��OF���Ol�A3ճ^5��Ȃf�OM�!*��'�b��1EL4p��L�	�:n�}��A�r��T�ǭ"`2v|�%A�^d�
׼i��	��ǍJ�,�ቐ��kd&͙=�f��`)	4`*Oٸ�ASn�@ �c�Ys�Q�[(��2�,��,L��!$W.G"�U��W2$Ѫ���@v���1n�
	l�xxs� 6�",���П��fʆ�0�`{���1o�,iӎ��o�|h[s��6�<�ݻG�H	��f��`u~�.M���C≵P�}s���;�n����  <�9� [4Q�zd�#��#}�>s����!ڨI?��Q�'M�-` 	L3ݦ�p��#�J�؄�[%
��Tx�l�mX����	�Orщ��'慃��81�Q��X��l$��"C�H��f�4�t�bXG�ZpHvI��tj�Aa��I�L&@�8�-]:\m���۸.!O� ��6r[H,����s�KP���	Ģ>�F�*�ʋ	H���E�HC�q�����P����A�n\���	)L���J�it�Y3�烊�R��ᴟL�o�?T���O���c� �8�)�#AZ.�n��,���&�rTc��!򄓕8>�MBd*r�" @�]x8Q�ã_���Dсx��вsi���	"�n������Q%/����ݡ7�^�w}cw"O0!�d�Y/_~�Qv�\P�i�
��M����%�>��5�gyrE �*�����H�{8�Yz����yr�1'96�#�5i���rژI�[���jX��W~�|�1
��#�p�P	��Q扄�I�$� |R�m��{ �$�-e�0)-Q�Ul���m۞q�!���;u�(��2�ĝ&W ���
A��Cg����DI/\H0"�G];��	\�� ���Э��K�9%H���E��-=����%�'I��C�,<��Dռ\�F�+��N-�ѨA��3�IE�G��r�fh!3�� �L���?���L@<@�}z�Y)Z<�����$�$�3P�v\	!�	�?ᡧ�=L(�-e��R��e*ف�>�yG �q��q��"���X0O��r
�AWj�q�@�K�f`������*��h(W큦��Ot\��"	^I4��V �Y��,;�Ň� F7m	�u��2'���@u,�;��	1��98B�I�!Ȯ,a��ڈ��q��� }�j�K Q����rc��yr'�"pɛ$J7�2�i><J�kt�Y�#@��VMQ�N�>���ՀJh!���'��a�玘�6�����c߾�pM)"�DQC'T22|n���2���i�N�����p���QA^�<!"��X%�)� D*Βh��� r�V9���iB�fF2�9 p��c�Һ�0��98,�^1ܖ$k�lG�H��i0V�W���-ɲg�t��$ <����S�l� ��H���c��O���VI�-k���Ƞ+�����ؓ�ؙn��[!#16��;w�NTKE�ʳw�>T����J(�����~�{��B�:��G!��t`c闺D���)D�`�qPK��5�t�C�4>�dq�7
n�Q쩈P���Y�Gl�'pf���$�r�&���@���XW�1;���C�D���͆� �Jţ5%_�d(D��:�`�B�'Y����^��ѻ�cתc~�X��y�#W�b|�\�'l`<kg��O�2�2T�  �'W�w��iڵN���Ӊ��Px�"����ٸ�%Ҿ̴�S@���O3u�@�~��!���tܺ�5�ƕ17�SB�<y���/(u@�e@�5�$O�Q�<��+�5BXkG��(Cd�C��A�<�V�׶���O_�>���d�d�<��G?J���fJ�p�s7cFI�<��H�>?�|���
��I�؜ʐ@�E�< �ڞ=��C7��-��;�)^�<vNÞmuj`[���HR� ��K�_�<�V@E��R9`u	X#l�h�)��C}�<�F囗^.��Y`i���	�B�A�<���M&.iZUAӛ&#,5p*�V�<�F��07��r ��(�| ЦIV�<��"�	X�$%��J�>hj��B�V�<!���S#�<�`��-\���A�F�<�/�>�V���*o5��*g~�<ɡQB�I�f^+4���iԦ�u�<��a�4>PvܻэF"~Ǩ����v�<���RI�DA1.���(6�
r�<� �􀓥��^Pqˁ&��(g"O~�;p
(�x�k7j	j2�L�E"Oܼ��J�'���B+�S�@�"Od�I��މ��CT%�3���p"Of ������c�4C�"O��9w��'�е��̀Ƣ�á"Or�d)�!�I
��ڹVB��S1"OxAbe�+xlT�pо�Le�"O^P�t�� ]dN�n��ȸ�)P"Od�����@��	WB�$p��e��"O�X1R��:p�Bg����L8�"OxN�eO>|��H��,���"OFT��
ˢv���C��=W�Z��&"Ot�#�
^�i�zq��%�Vm� "O`�+��M3z%�y#�R��pyU"OV�2�)�83Jy������u�4"O����H�/i�����ԺE�e�7"O�u�-̙n���Y�V�
e*"Oġ�ÑF��d���ա*��lQ2"O�AB���$/^����]pCw"O�xC�,�_�@�y ��Q��"O�4+6HK;jf�tLp����B"Ov@2T�^4Ddqm�0�����"OĘ���0Pj�e�`-	��P�5"O��X����ry�=H
�[��,�"OdM:��ߓ.!�mȑ�ȝGr8��"OJ��D��4�l�� - v`��"OX����<A(ٱ�o�4|,z"O�XIm��	b�Ы�(�gT��"O�Q���	
6)�6�V1>@I�"Om�� �X[R%A�Ȅ*.tS�"O��!F�`m ���g�4�Ɲ�!"OJ���l�B{�X
�݌7N����"O��P����ъz�(Wa�`�K�"OlYÓM�)}b���d��ݒ�� "O���QZ�%�H衷��E���1"O��{��@�Q��\�X�b"O>�`�m�E�Rm#E)�,�i�"OЕ;��A-!�`$��5����P"O��s����"��`s ��"Ox���
�a��5��"�>x��ɻ�"O���2�MR�}�PC�-mĚ�S�"O��pwAE2*��jw�ǭ*�����"O����m��W�� �B����"O�AK�X+ ���K(b�0��V"OX�r֠F�uk�d��@��
�|��"O���6n��z��p�Uۍ^��R�"O�@"Ec�/\R\���Q��(�"Oj8�1�IIi�`�WK^�r4iy�"O�Y�/�-_}�eDX�M��� �'�4	�eҐ� ��((2M�'�T�[���1A�<�J�@Q#D�L�c�'�f��&�F(�U`ajзl���'� :棕q��ܰP�ׄYP�Y��'�D����˫;<t�a�K1HC�Ip�n-Ӏ(+�2�c�lC:�BC�����\#n	2Y'�$�B�ۤ�Z�-�/*|1�m��`.C�ɇO���� ��*��4@څQ��C�	@�@Iz���3���Z���n��C����|*dI7;��t(�cY{��C�8B�@P��7$w��[��5��C�	w�"� �.3[�th�F
R��C䉣V��2kI�w�m�F��}�C�)� F �dV�a��H��L�z^�!k�"O��"*C�O������?51ڤ"Oj���E^�
4�|����=��:�"O!��1xU�� ��rZ.%"*O� ��ᅛ&�tZ�)W�J:���'+*Dc��^%k
�h���/B.���'�@� PKU��$d��Y<���'jrc��Þ|�J0�F�)"y��'���3(�
���h!%�ZE.���'r�h+D���;1V� 5��r ��
�'���SՈ�f�"�"��
iFA�'���zP�Q2X�m���AP�Q�'�ܫS��B��i�D^�I_>���'��
�ˏ�|P�J���S>����',�գDJϠu�(���!LAx	��'�U�@-S�VĵP��$;�XiK�'���p���\�b8��l ܬ��'Yt<�"	ډ7���օ �w5��*�':�dr'�z��(VL�)y$*�p�'�B	"�(
�\}�h˝瞑�
�'W6ѹ����@y���ӡ���B	�'���	)��b�����/{Kv)k	�'-�p�B�l��Y"����iE���'GlaGM�C-(�U�i��U��T(�1�7L�4�C��ҥ~���K`�	K������4� @����<�$C�73:�y@A��c�d]�������ԹM�4eS��Ύx��y�>���g��ħ=H\�P5��LrU[#�	jN�'�ࢦf.���|rre�S��$y��6����j�P�ʩb4�dl��L��%�ܪFR^UH��O��-���ԤV Y��J�T`ʳ院�NI"q�@U�bt��蟈�įK�	�咦��j�����L��0� ��i�����0|ZV@�C��h�sc��_7���q��e�-9�+�f?�,�{nd��)V X������vH����%S�F�`nZ���]��.	���`B¨8�LȲ�g��9ᶂ-t��x���� ,*��yF�ߓn*��JW;Oa�t��YA^*�ňD�\ � G�8h�%��%?Ia�q�a��ח;��4�g���|u�gƎ��yDU�)g�@���U��<(��ڮ�y�O�r �Qزc(h���#��y�DB�-T�$��ι
�^�����y��<rT�!�܏x�~��!����y�C��F8��8E�6��+����9�S�O����@I@23d!@:[_|���'3���i��B�$�$�G��
q��'�4	�)�@[@@
�,+�BJ�'Fl�)T��p����eG����0�'=��𧩌�e����C�3�!��'k�q"$a�Q��a1'�!�5�'�f�����%�	� �
�2��Q�'�&e��n^2hĨ�:U�'��y�'����υM$ƈ�G���r�'��x�L͛-t�]�1O�%<i�'��	����11^:`)��Z� ]���'�v=���633fq�dK��'��� ��'����7o �PBR��	�'�,��*�t�zw�W�0��	�'�Ȁ#��7Tf@�SmL)1�΁�	�'��t�4�K�P!m��툩q�����'9����a6�2�11�ɐV�Z���'��A1�J`y^ ����T�V���'��i!4o$tzJ�0 	F؎���'��v��$;��U�'�ѧDo��P�'|d] ���6+� �C�+����'��I3��cIf\`u+�3�X)�
�'�vup��2.�R�2������  �!ਈ�/3艻�c�]DF%k"O�,Ҕ�J����QC� 53����"O< �HǂlX���Ѡը[)��`�"OX�ѣ�k*xx����yY�"O�d9'�ܚw�"�B�,A���"O��U͞[�<1뀱5����1"ONE�5� �xT	ny�I
F"O����a�v�PH$ȅ%=��ȃ�"OY�bN�-M;�511��&S�H,�"OH��˒�d+��`��\���D*"O���s*V$9ܼ��D�I�X�ʉ`"O�Xyӆ@�yJ���B?�N�J�"On ���#r������r�6�Y"O�Ɂ��sNN(@�H�ݰ��7"O��3-�3@��#��I�y��\��"Oj�r	F��q/� h��`�&"Of�H��ʑ33���.�=X{m�4"O�p�'/]�]^�m�R��J B"O�]"��� ��A��l�8yg2;�"O����?�V����6L93"ObD�c�� vµ���ֵ@�] "O6"��Y�{B�e��AI�qr|w"Oz�hlZRȢ!�e@-k��k�"O$=@�.#�8r��  "�Y"O�z`��{�贫�̀�g�J���"O��ѣ.��3gf@����"OhJe!Z$tr��c��!�hq�"Oؕ���#5�IL�!���"O��y���8XY(P�P��2����"ON�9'�K�V��,`R&�<N�=�"O� ����gr��j�'m��k��!��~�����nhQ���ѦtN��ȓ[��yA傆0���S!�&�����_�����"�����S��p��A0��%'_:P�ER���#���`�Zg቉V���Q�i��p�x��A2����J+V�v聳I�K.0���gl�ٰ��%g>�cg̔GI���h�:�Έ�G�VA�b���I��w���e�*fId1"§�:&U�5��N�n�3� �&a�2ɢ���[����Q��b�Q���I�o�<y�ȓ]=�� ȗBa�	q�$V�9����ȓJ��;�&��N����^�@��]�ep��a�Ȁ�]�j��a��FVH�%(�>`�X8�64�n,�ȓ|B)b�K�&�<�IU��X�D5��W�f�A.N�f�)�6?�4Y����L�x.Ե���0n��ȇ�b���Sn�?Ch�ԈW�cy�]�ȓP�;3��&�h9j�֧)A^L�ȓf��P��F�a��t��5�T�ȓXzx�h�J+���a(U������!X�Ur�d�u����~�L��8<`#uċh�*j۴
�j���\����6$ρg4M�$%�J�ꁆȓVSh r"U� �V���N�V�8��ȓnRj�KrEٺ�8���Z �ȓo�,Y�s��9ǒ�ˁ��>n�H���]���֢H�j�����lɽP�ڼ�ȓ?�e���g��)�ֳ\��T�ȓQT��!�J�n���S�^P��K�t(�pEͷW��1 �!H�$E�x�ȓRc��(�N�;$`���^�jх�S�? ���gdkw�2�P�tTD͙�"O>�I#��YpwG|8L0��"O�p��#�xtk0���{1ҁa�"O�hTNM���hD�SN`s"O��a��Ϡ#����C�=��e��"Ont�0 �D8� "ƒD����5"O��[4n��"�F�P�H�4u &"Ott�K�/F����ʛ�h,˦"O�����[:^n*�	M�@�=��"O�M�ᇛ�A��|3���
�^�� "O�!��C1V[�X�H�/g�ݸB"Ohy;Rc�h@L���FQ� af��"O�H4�I�_�F*�N�=`.A"Of�ڣ��Rb.k��@lG.i�%"OX;�N0��- ӄY��B"O�]�2(]��Тd֣A�4�
�"O��˱�N,���!����,��7"O�Y�Q��֤�b%�$�L��"O�����Q�9�ҡ�� �X��"O��1Pc̦.�lkAT%7iNA��"OZ ��ݸ0�����'RKf�xV"O���jU11����T/��A0�x�"O�h�p�02�&L�#ɖ$<8�&"O:uP��o�m�.	�x�(�"O�;f
 �/��]�c�Go�rt"�"Oޭ�`LM7}�lC�JE?��m 5"Oeڐ!_	dzi�`i��B�x�w"Oj�:R(W&k�f�H�(G�AhV�!d"OFYzE�-t�d�g�;DQ��G"O���r�F=zh�"lG#=ܫV"OX�� ��*\cP�5� C|I"O���GN�$���u(�|�8"O��J��H(j �c�οs��%��"O��i���+v�XE�N���AW"O��gä6K��ڠ,;�.�#"OHXs�h]=^:���#iۿ��xR"O4L�a��(���Ć\�F�s�"O^�)�/�#$�,U��/�2B��ؑ�"OJI�1�B6^INܑ�m=!��;C"OD�j�e��s�f|{�L�G|�$�"OL�R5n��0� ��3|��bW"O�԰�8l$ ��B!a�.��"O<�C�+Ux�a����<F�D�z$"O����T>� �ҥ˕�yo�,+�"Od *��R�6A��´PnA9�"O��a�����8�R��٩qV�E��"OV�
��q�^��3h��Z���q"O$� ���c��G�y��x3�"O��U�ĵb,^�U��(2�T�s�"O�cjɼ|8l���՗W�dhv"O�8��V,g��I5�Otq�s�"Oq'F�6Mh�1���C�r���"O�@ 5��:p`��ц&P��X�"O�,*�B�792��1��بF.��#'"O��{��Jzs(K�n��yplAq`"O�A�CJͯ �;�nZ3FF���"OZ�a�E��9n\���deZA
�"OX��gM�He�	 �=n��"O���w�Q,�Yғ)�\� �#Q"O�0
&�<=�X�UiH�X�t�p"Oju�C�n����HD;?#F��"O�)��H�+2���ȼk 
��"Ohj[�.|����3)���"O>���].5��2�.40튑"O� �ŉ���1yw�� #O(j�"O�@��@؜M"(��.H�'0i)U"O���6b�~,��r ��.v�kW"O.dR���R-;u/Ph�T"O2��7/B&U�1�t�\9r���jF"O쁣`�
�L9�E���
oz���"OP�W��0����4o��Td�ՠ�"O�t���͍0�A�dl&+QraZ""O⽉���mT �t̂�=B��D"O���EA}>��&��	{��܆�_w8��uj�=�q����<A���ȓM<�0à'�k}f��Ө@�>y�ȓ5��p��� g�*|�uI��N�ȓa�6u��n¶Ƕ�3���F�,�ȓU�8t�d�-,^�K��E��^���6qЭ�򄗷<�p��a�6�&�����L�#� #�mc����/�i�ʓH� G@�%`��� ���+dC�ɗk���FN�+J�����U^\C�I�@�& BJ��D��q���#r�XC�	�V(�ck�x��m����U��C�I�DeD	e�#YI�ips@ScY�C�Ih\�X��^�X�ဲLQ.�jB�9d��(�SFR% ��iT�.)��C�,vO�,�V�
�fS�)�7r&B��??l8uG�#q��U��AX��DC�	>�L��N� �U�!��u�TC�&;dB-������e����p�C�		Q��٪���V�<Es�k�� C�IAv��L��I�:Q�bc �B�	$<h��#T�
�Om`ѹ6eY�-�B�	�[c�U��׆]�$E��?�B� DD�c��D��-�
M�K�"O���C�w���S,�7��� "O���	ί3ΰU��ζd���"O8��D�B�#*�Es�KR$*���S"O`��$��T!�UpD
��<�&��"OR4cc��y�´sg'̤i�p���"O���wH��n�n5A%J�O���3$"O4%!��O�l9� ��A�3d��1i�"O�:�.�z��:��_/��h0 "O��KZ�x4�Өs7*��"O�|3�=�,��!���m;�"OP�"���:7>qpH]�����"O>�X�D3p��$*7	϶f�,���"O1ɡ熖y|R��P�b����"O(����̂9&��a�$���"O$���˙�FV���e��5>�M�2"Od��pĎ���$��K� ����"O�ͫ��+�hI��� e��"O$q+%g�$Ƽ�^-��mk5"Oz ��NYs�@�h��"J�;F"O$l��,/^��[*�S"O��S   �