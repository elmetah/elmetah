MPQ    ��    h�  h                                                                                 #�J=Bʁ���7qt.@�ր��U��s�<����OGu}FJ�3�S��
��)���.��/Q,��ݭl�Nj��*L�Lr �WJ8�C\e��P��(�;�*�d�����u��~1��� D�%s��|�F��[Hj��R�hpR,@"��B$���7��/M���H�$�xfq��C�}o����p��uQu�ݭY�=J�����BIrq8Ǚ�Y\ǆ�!���<6�Bڧ8�� �}lw�Fra0ݮ�_z]	^�{�ʠ�B~�S��(�E�$_��
��q�}yii��P�^I��n~I�I1�(�@������Xw���Y2q݇!!U(�����Js�����5�NS����6��K�� ����kt��I���A��c�6ߦ���q!k���w�w�Y2��]|�h8+�W���0��-���+�"��^N��ᆓ+��c�;��L`K��r�Ԅ�C��4!H�[�3;�]} m�;S�{�����yO�
�1k���@ӝ�/aU��,��"+�r%	���6��U��S��z!;&��U�i��'q�#I�`v����@����"o��G���o��T'� .	�g���4v�� [e�GH݋����w��G� �ػۉ�j��uf�Z�����b���lѹ�ɘ���k\�����zpz�{y�G�T��w?��1��tU)=� w��d�=[�#�g��WNH�
'�|~��V���j��	M�`P��\yԾ�kl~�~�ա�����9Ԗ�{0Rv7����H�Y_��N��L������х$�ɍK�7/w2��D�(���0m�4��V�-3Q%�D�8���406£��KP8y`�|�)ˌnD9�*�YY�+o��JޯC��s��$�CŠ��d�)����/e7�J�!Z���n�/E�c��`�����ȀgТ,��{�&�Y �OQТ~s���F
�6ph17�϶R�5��i����1�xQ�gGz��n�=+���L�f2�n���(Jg;�:�s�[��:S����){S9i�1�;�)H�Kj�س��Q�	ۙ٧Հ�_/��A�F9�d*7P�?m�k��_r'����?�
"AeF���O�z�vXK����2Q�ozG���-+�d�	�fȢv#������.������/�71��[1�<�1(�a��|u�v��*�
�B���{E�D�#��?�#{<�s�E���˔[�:���Ώ��O�+��!΋"6�"��:�	W+��;�t�Vi��� �c����+M�K2�6�gɈ�ݪ��)%��h��E+&���%]�M]p/�l:�T�N�ع�|��n�ӏ�P�q�Db�"֑��/b���L�iɣ	\G�جJ4���%�v��J��?XU��G	��VU�}�����
�8��5�H��D!qv��)���w��"8�~_E�:l4i�������f�*����4�[K�����T�R���3uf���Tj����3�U?�as����!3f ��mi��~aǓ��U�VU&�A�����L��CeyU`��sH��Nw���Պ.5M�Y�6:B3V~�Z-���K�`�|���.n��	�E"c��OA�o�9���[`�q.S܃�Չ�Zͬ�6$�o�Q�Fi��&g`�'CO� ����%��R�4{#��gVud\���#a$[*
6�/�p�je��	;��(�t�ok23��Y/�=��5�H����G�e)'����8��'V�b��^A�鎧���>K.:��F�G����3�� ������C�9�hc��|u�&V_����f��_�=���g�ژ����:��_��N���]���%tkw��S��@�~<��G���c�fm��.�|��Q���(D���xD��|�|r0��~�?S�?�_�w��l��8*�)VV5�ƪ�i >OY�w�j�C�۽������q��c�E�4�X�ЌT2�C�ġU�噮T޻;�"��fJJ	]�y�?�ϩ#��DTD;���+察�o/��' �Yz�l��?�e�?H���ٻ1�O#��0n��,Q�|�=��y��Sq~���Tlf���"�>Q����8i���'�*՞c�N���x��g'�]	n����R�A����,=�[w�ѓ�D��{\��x��s?��Qǌ�IV�k�c>�ٚ��:�)��yǷ7UyRa�O��PZp��_�P��5e���+*hcf�i���O3���k�{��L�I��6Sܦ3�KI��)��!6��C�s$���z��b�>HW�i�9\Lj����HA�71���?(ɗj��<7"��>Af�-z�kC�5ԥ�Ը�=��U�#[DYQ������a�謁��1�w���/!S�ct�
�� |p�ǈ9mBM��4O����;���|�'��3�X���}����M��S�t��٭�C����cOƧ����#�45{Od�k���+j|R�����dE��Ž�=�_z�{��v��oJ�eh}�� ��rUGR>h��dcJ�Ӗ���
>�Y��t%\��ܵZƞh�X�a'7�q��b>�T�!�	�:�
u�a��$�7q���wƍ�^u�"�U]ˬa�- C@�<�L����on�Wj�o�.vKZ�2���a�� ��������3C,��~�\�I��g�d��m��p�bY�˞��=M���k �]���L�a^ɢ�	��4a��>Y�S{r5>N���
�9�K��Xn[��q��Z縀���on�P���E4CM�vUo:;/v��%u��C��l{�B9݉F�� �gY4[,��9Q �1��S}�H&,4�Ѱ����&9g�A�I�"���3XݚG,�ۥNZ���ۿ�b�%�VN�c%�4�n�Sւ�Z�yȘ��Γn3n&Ώr	5��+��T�|�Ⱥ9���7Sw��e�?Dy�!�M[�1�0���)�}���c�䗜��|@&"G��l�0��+�ٍ3�u���=f\�6��R��T=0�������js����_��L���b������'���/�UX����go�D���1�E�e������ ���e�Tx���t�h�	����4չ|*���%��p�nj�C��V�7d����G�d)3A�r�^ϕ2-�0����G�I����ւ����-٣΍��G��=�u�P�>L33Żc�P�t�B���C���˛B�mq33;E��AF�4��<�	A��bY�s�j��M}g�@'�r���x�]��7{����}Ł� 4(�G�$�]-���q�i���+��^�T9-[I����M���:�)}A+����Y���"&�U#D��Gt@J.$��5l��S��c�����!� �g?�H�#k/�xI��A$T�cf�C6��}��!��� e�w�^|Y&���/�hN�WGߵ��K-� φ��"H�^i�\�Z+w�4c�
�����6T��2�C���!c7:l}�;�֤����n��vR՗�L	O�Dm1+���x�T@���/= ��|�h�|��;b�i��6��z�S3�jI;O����Ű�LK�~���5��1���]���7k\����o��3'Y��	8� B�Q��;�,e5R݆O��ғx$+���S|��d��X/u��B�%�k�����	�F�ݾ�mz��v��G����2��L��t�:�����@E�=��l�b:Ws���� ��\��[�ӳg�����Mb�`K�F\Ԛ�&�k��nu�s�]á����r�R�{����?�|j�i�3L� ~Ȯ45�N����d�FZ</�NA��1@��=mk?Ջr��h@%;�8�)�4�}7��fړyۀI�H�nQ1*��RY�>�����������! $H\٠i��db폖/e2�\9�nZAD���YE��|c�ţ���V�cv��K�J�{R�PY;��QKQrso&6FE����12����� �i���+x,�g����h:	=&�jߧ�@2��+n����;�sL<~Քq�����s�S�ݢ1H�)ä�K���ړ�D	�nȧ0�__���A�=1��.P���?�K��Ilv"O~���
���F�j#���u�K�K���͂��j���ߵ�+�z	�ygC�#]'-����$���I�W%�7�)P-Ϭ���(��M�]�u2�C�%�����D�6q�0�9��)V���#P��B=�ƌ���HPhQ����4F��y��ƾ*���y�5�W�-��7��q�c��9� ��S���M#څ�1x{g$*d��w��̍��2P�� ��ݟ	]WG�p*;ul���	?q���"�Z���jx���hb^�q��{�/�� ��OɾC�\ĝ؇wM�Iq�%F��Ec�?�w�w&�qz�}r�`�[��sp�5�*�H��6D|���˖�����������-~�#�:��i���%\�!?���4o�k�r+ڟ����"ua��JUJjtj��U�E�s����l�h 
Nk����i�a��_����V�����A�J�BFP�Ch�ypzg���eC�wݸ��%�M����Z�B��N~�-
E�K鑵��(��a�`��`S�a��cg)nA��9:��[;l.��f�p�=U�ط��omʭQ����fG�``W�O3L>�6~�%���Ǐ �p;�V�� bg#<��[e@�����	&�`��;A��ȕ�!�3�
'�p��1���0u�����G���)B]!�n"8c�Z'����O2(���h�>>���z.U���D�����3���;D����g��#�u�����g�M�ޡ	���`V��gGW�ٙ��t�~��n���I�]p4�� �w�K5ʋӳ"h%�)u����/��bm�e8�)%|v�U����C��a���S���_jr�y�� �A?���7��3�Zl����k��d��5��d	�O��#�%!u��h����dO�㞕�E5��XŤbT�`���z_�p�ؙ)�#���
LJ���y��:�dmu��ŜD��
��_R��[�ʂx��5�'{��zǏ�ӫTe/σ׼>�l�P���0i��,�{�����y��xq��ϓ��Cf���"�% Q��	�hϧ����EK����GۇXH)���]9��I�Rq�����=��X[R���B�.�N������Ws��7Q⤸Iњk��t>)���m�)����x�a�R���]p�_�Ah�C)�5`�y� �(*#0f�W�U#3գk xF��'���-I�
fKS)'_ !��fC���_��^i ��	�Wr��9w��E(NHT
7l�9�����$-��hKݑ�>��6��`M�CS���_M��Yδ8��#]�t����s�r�X��?�W@4�T�w(�U/� @轤��O W�E��m��`�/=���9ڞt@�+F�@����:���}1�H�H�=�wX��/p��!�ш�p�\� ��%�Xp�/�UO���N<���qc|ͳ���Pt�l�E6�ڽ��j_��5�hp�I��b��D����U�Vh��d����Q$g�%Zթ����O���0G�ZaP��Se�'^���ǀ��}E T����䔿E��~q���7̺ʊ:�ƨ��u���0B����|-�ʒ@�&�<'ݫ{g���ҁ��j�Js?v��2r�Va�����I���:�T,ukɨ7������qm�0����b�����M8��kۋ��`\\*b�~|dz���Wa�p�Y��{M�zN䘨
�ز9���׳�ڏ��sq�*jՓ���1o�l��p�pE/����Q:��Fv�K%��iC�y-{��$Pq�]p��5s[���9l'1��QSXE&J�a�E����j-�ge4I�l��<sX��Gga4��9J��˿����9�N��e����I�?Sfn��Ӵȓ[$�)�3)j�7	�h+k������Ԙ�2�k�)�l?�E!�X`��u@0`NF-#�}j4#�^ė�2��њ�&,G�w&��}+/l��Mi��h��Das�n�m����A��'d�-!��jy�~��_�΋�@�}���$_��f���I5U�4h�-�oyH�ˤ,�`a��G����
fU�ae�Ux�StȬ���*�����$ۨ����j>Qf�ҁ7�gO�J�v�b��d�c��M�Q��mv-��ͥ���G=�����d֝��� ��x�ۂ��=��P��DL�ܻ�C���>�'	Y����1DB�q.���P"�����O�<,θУ���&��P}b�l]r�;�ⱔ]��{�����,��o�(�i�$������q,�i_��^�ƿ���I���t!����ՁD��k�[���jݽJ5U���+�J�̆/�X5�[Sg�G��&z큱8 ��#��b�k꿉I�hKA���cA�6U���{�!��A�[rwxQYA���SyhW����fS-�M��j"G^�J_ף-+R�kc<nł���8�:�2C\fj!~�@��;�o��hp�q�t�q�J�XOB��1F���cS@��/x�|�Z�����(x��$� 6�m��2�E8�;��������摡�����5�2�^�6|lϮu昑 ���	���+oA�2'��	SD���ם,�Ov�2e��݁*�w&��N�EF����\�?���C�u�k���'���WƂ��<eɎ4G�!r��F�jz;˹�q;�G@Ui��V��g�tK�C����{F�=��͵]M�WΤC��G��Z-�ֹ��B���=M��&`F��\/�(����W]��B�|Q���R�����G��ϸ#��~LXyȉ{�����ZRx�A��/-�Ղ��[�'T�m���M��ãm�%���8��4��:�s�|����yVn��n���*%�Y�qe�UO��������-$Ô��DP㏟a2�*Ae-�J�qZ����olE�l�c`�V�h�����l���{�YV[�Q�rsJ�/F�V��I�1-�m�l����i� ��D�x��g�"��&�=!@9���2F�n)E��1;{�s��t�/ȃ����k�S�rd13t|)>TEK��iN�o�.�W	�c3���)_��AU��Z��P��?�Ю����y�
�vdF�l��E�@HK���hZ�epr�:��+Y��	g0��w#8���#�s�����|���:\7��H�T�2]�(�&��u�1�� �ޏ�1��(K~7�uP��
 #��[��M��xŔ�k?���8�E������{ӊX�9�0�^W�����U�{���� ��|�FT�M��1�,��g뵺SdH��L��W������r�]�`�p%��l���Ķ��:N���O�EȦ�k�b����+/�'�¹Y�ٝ
\�a3�bĖǄYT%�5i�@F�?�����Ό�}��6�NӮc]5C��H�6�D�+糆����Kq�m$ի�]�~�!4:��i�|�W����⏡.�4�8��My��ʫJ���)u\A���j/6��9�U5_sy�ʫL*Y�� �ƿ�P�Hi���a�w�s}�V�40S�-A|$�ߝ_����y����I�@�bw����_M����C�"B��K~�ȴ-��2Kċ��]��������9��kc"��A�J9���[�.�<~��<P#���8oo(��Q�` ��`;�)On�C��0@%������+��V�T���\#��[��^�e����̻�7;��;je��3�����O��.A�+L�C�WGZ��)]�ؼ�/�8>Pb'�`���%G��<f����� m.pZ�<���q��3Vl�֢ʨ�����k�|��9�i���t���܋��*����g��k��$ҟ6����I%��1�]i9��wP7�F��=r����i���+w�mO'�$��|��j����^���,)�.tȶ��rf�#��y?	&��� �N��ly��[�jן��54�#�_2�O*P��t*�4p��[�?M]��NAE���X��TT���ùY���<�'���ǳ��J?�2y�drx�H�ט��f-D1J��v���+ke9Z����'�`�z��N��7e�>������EY�p0d@[,p���y�y�[&qt-,���+f6�q" ��Q�����ާq��`y�Y�c���Ї�8���y]�#���O�R,MЎ��=��[-�}�}�l�� G8.L8s��&Q�܋IL�Ak�K�>dƔ��$)���m):˰�a�ui�=mp�_Ss��ag5[���{��*�fmf�e�&#3��k[��͂���D{�\ �K� )BX�!,�qCj�"�!M��w��ܟ�*�W-��9��+���H��h7�c�'O��k�Z�_�i+>����#�l;O�CA���#D^�����$m#ѿ��eX�q�M?��1Ī�A��Xw�$�/��7�Ϥ =� 2 U=�mx���*K��A\��Y�W��LŻ:���=z/Q�}�" �C�ٌ�P��s�㜨����7�B��k��Ա*]LO�a	����ׄ|H���t�����aEѧ'���V_0��#����[1��h��$o_U}��h�{d����@�������*c��k��Z�!��Nj7'�_�߂����l�T�'п>����2�ٕ{K7'�4��ך����u;q�G"�"��-6r�@���<h!�6W������w7�%#�v��y2̢azV��_ѕ�W��U�N,�V �X�.c2��tm�aQ&A�b�n���k9M��Kk��S�(" �~�z����h�a/�Yk�{(wgNe+
&,�9��Y����V�q�,P`��m�o�C��lHE*G��,�:��Bv�ߖ%k�WCi��{6��ݿy�C�2�[�~�9��1)1S3��&���F��+���T�g G�I�ܷ֮�^X�v-G�Y���9v��w�;�����N�m�*�$��SLi!��>�Ȏ�Ąn?3�G��	+J�+F;��򬼺onI�-E\���n?��{!��m�'�0;�Jh<�}u��Yo��R'���&G.o���9��+j@��i����/	��B&.��鈛��Jf`a���hP����x�y�m_K��\[D��rI���L����5�{U��u���foqͼ�+�{8���P�˱S��eJBjx~��tjGq�=���r>ۃoz��h�j٨A���[7_��{�};kd���([���%-�h����G��嚈puָ���DT���f۽Mq=3�P��L�s�ٙ������������y�l��B�q)k��{�ǷSߩjvC<�L���h��M���}]|;ǳ$r�5���
�]zs4{_�L��$ި(���$p@Ɠ;WsqG�giڌ����
^�X:c�|I����� �q�t�_��70��6Z�ϩ�X�#U����DJ�k��J�5bucSB�[�1��a� �����dMk��I�mJA��cԜ6�`򳕏!�Tg����w3��Y\�A���Jh��W�u��ټ-�R��<ZV"���^�%�R�+-�2cw7���Hؽ8ԕ3CU{!��obp�;_(�.=���l�D���hO��1að�n8�@di\/��΍� ,��꧃Q��ߊU6�	��IR� G�;ń��&����s�4�����M#P���h��ӆg�m�O��%o�#R'���	n�h��TS���lek���|%�Ҁ�	��aH�I]���O�u7ގ��?�ے,����
���	�w��,ᾁ��z֨M�l��G�k���BtƌY�H�߶g�=,
G�X�bW)�1�;�6��x��Q�ӳ���x.!MP��`Aܪ\���˜����`��i�s�Wh�7�>RG��|����׊���r]L~���d���7���<��/��i�u�{�B3�ma���(ܘ�޺�%q�?8}4Al��.�y��NCy�{盺�Pn��9*�CmY�����ݯt����k#$>�e�����V���e(��N*Z�5I��gEy.c;�y�L������� ټ{�=Yq�fQA~s%��F�ϾA�1(;r��KC�f�i�D�~�x�a3g���Ş1�=�C�]N52#�nD�/�w	;V�s�:?��>��!}��eSj'
1N��)�#+K�F	�"�ɖ�	�x��=�_`T�A&�����P�w�?v��F�]��}�
SAFюY��qpyUK@^M��r�`�����+W	3t�9T*#���^r��Z��w;p'7b�Oc�¬�X�(��vL�-uh�p�ÏSu��(!fa=���� +#ƎɅDu����l?t�5������7����_�<W0��a2�+�cW<zbl��4鄍�� [Gv�;$MYW5�'�g���q���{�(���Q�Sd�]���p �lK���N����Pfu� ܛ�"i�b��p���k/s�n�}܇���\uu�=1ǿa�%RE�;IT?iW�x�Χ$�}h�����v:5��H�8D2�/�A�����w��� )~@":=eai�s�v_�����I%4e�а(���$�R!IuW�� �jꄪ�TE�U��sT����^�7ۿ  K�!ΐ���i�a�܃NA�Vts��Aw��������y���]�k��wS-Z�[�)M{H���Bd�L~	��- �.K����-�����{`���?c��A#��90��[�չ.���`�K~e�G�o㵷Q(�\� `O���l�%����E˔�<V��aX��#��[��� T<��ܛ��;���8�F��Z3�v2
SV�g��&����{G+)x9��dq�8�'�6��9���ß����oR$.�åݷ=C�L�43��q!ݨ�XV���9�T��|�O���.��0��
��g��UO	F�ހ�t�q$���l��]��s��%w��X�YMX��0�ӯ�WO/�m��̀k[|,��@��y���W�n�	<Ŷ-�Ar�q����?dB�����i�l�|,�61���`�5�'T�Z{Oj�����c�,؍���kl�(4Ek�2X��bTCg��tX���6��2�̐�K�kJ�?�y�C��l8��`���'D�.��Q'��P' ���iP'1J�z=���	�?en!���ػ�.��x0_�k,b�ٛn�y��[q���Q#fq�b"�^�Q�>��I��,
�{���s�t���H��8�]�.���R�X��O=��$[�K�������T���xspzQ5GI�1hkj�>������)� .���{�|3a���p���_T��y��5Vc���y*��hfۓwO3�Żk��n����{�ܷKz��)]q�!���CEwa�heҔ�	��#�OlW�O9��(�;H�!�7�d��¬��&��!tSa�>Юp힑kqgC|폥�H�ziŴ�i#�B��?����(���|����	��w���/R�RR��{�� x�x�(m}��%yL��IU����k;�6��`�jϻ}gh��>~q�-i�������7g�~���m�Xw��FQ�%!_Ou���y���]�|�&o�O"K�u�Elì���_�������b ����C,��_�U��h
RUdt���Ǎ��[�v���2Ӟ�{Z�ՉI�\'$x�= ����T3�К�y��ԕ�ڕkW7�y����b��+�u~����kz�]B-�9�@�| <�;'������v8У �Pv�[D2���au܋�����G�p�0,kb#��҆�i9F�5�m������b����^�M.Fk��&�c8�������#��a-�Y~i{HNZQb
���9����ia�I�q5�7�L �H	o;ͦJxE%���ɴ:l#v�z%��CD�{q��Z��7��xN�[]& 9���1���Sɫ&�����/�s� �^g�ylIau�2��X��G�q��YZ��߿�YTV��N5c>������sS��(�+ɳȉ���83��Pz	���+!N�-��
dw�(�H��^�?u�6!�΂����0*��u�}��a�T�֗��,�G8�&bd��m�����9+�������}n�Na���飼�Ūj<�9֣�D�;���t��_�A��,��~@�^%�D��p޵U)X�����o�A1�A�.��/��=+�ˌ>P�i�e�NYxy4Xt��U�:���0{z��:�^D�!قjt ՙ�7^7uܮ����ј�d�$���(�FD)-�xۥ��G�ɛ�C���\#� t�_�}���m=���P}�LD4���ŵ��#���6��e���QB�7lq$7�L�h�r
����<"�l�����$?�S��}X"*�rMw����]��{:�г.["�l�(��$����#$qbN2iUt�����^5����I�=��*���,9�z
��b���r
g����U�"�X��J_N��e=�5��S���l���0� �P!�Y�Bk`{xI�A�M~c���6�3��N�I!��h��w��&Yw�}�I
	h�v!W�S5��~i-ث�ϗ��"y.�^� /�@�+�c� Ÿ�"ظBT���C�c0!�����;:�i1Dʧ���g�֗ X8O��}1|����,5@?��/��M�J���J�����6�[�đ��uu; �^�����{¬�	Lu�h���,q=�Be���A-��j�o�r�'�+�	�H���b��ך���e&��w@�-�`��iU|����}���Vz�u�pP��3�68���G)�%��Ʉ�������zq�٩g}�G����c���fytAC{������=�rصS%!W�{��������̜���R�z�M�|�`<#�\孒�Wsͩ��� ��2鎖rAR�I[���e�E�B���L�f��?i8���*���7�2/�c��0韾]2�m܆��z�(�%�48x��4�4�鏛��8�yL����~Gn0Z*[ÎY�7L��\�/�1��@�$�eޠ�?��H��`�Ae#�JL�Zr�v���IE��hc�����4D��[{�5yY��)Q��s `�F�hܪ�1#��"�~�!݌i-���׼x��Ng3K�9]�=^�߸�O2�ln_'�-;1JZs����e�����!S%��1i,�)4}Ks%��ܒ�d��	ǭ}�A�_��AA�I�PT[P��?Y;B�Rﷷ/}/
,�F��p�;�oT��K{.D���C�[捼��A+�{a	N��$�#�fG��M	��#*�r�Sh�R7��~��(t([����um��g������g���dK�k���~V�#�˅�+����/����L��:��;��p���wSA���b�&��W�P�'�F�����n 6�?�BM�E��"^�g5���ɝ�z���gñF���vm](��p�)l��P�:S�/y=���&����]�Lb/uԑ�#H/�K��8����\��b�������%�t1�6l�?Ğa�3�j�©�}��˛����$�k5y�ZH��D�fس�@ʑ,��c�W���~K~�:�ji��]O��R��d�04���u��@��푀uR)�[��j��@�o�VU+s/�6�²OҶ� ���|���Ɣ�i1�vaY��)%�VAӊ�^�Ar8M�S�}�t�vy���1����7w����4kMv-���B�Q~$�z-{��Kz��h(��2���v��rB4c���A>x^9��g[̺�.?I�A�cF�ŷ��o��"Q&����h�`�PO�J��%%�Ǡ�z��V����i�#�O�[�W�������P�q�e;r�S�+[�3w\E�����!����x>G��G)�׿��ҏ8�Q�'B��� m-��j�Oq<�*��.�L��2���'ܠ3̺���G����x>�T2�o���t
*���R����q��ygX�?
qk>S����(���Qr]A2F��Fw�ʼK�s�е���ӊ��rm��,�>�|�$U�=��ɔ1@�ҽ���#�h�+r�����5|?����K�Zل�2l�`��k�O�5j�|�U�RO�)�V|!�G*H�
|2����O!�E��X���T� �/w�����z���y����Ju˷y�B�.K�ϕ
,�		'D'3��,�z��)��&��3!'�S�z����$��e���h���O�0ZJ�,����)��y��qjB��r;+f��g"V+UQ���&]��T<���@OY)�O�K�	y���E�]�Y��ZD�R��#�	�==[�j����F �s+|1Q3��IB�zkEJ>�2_�>�<)���#�=Ah1a+��~��pz�_��E�3�5Q�
�1��*T4f���)�3fk�,͸r��ғ�MK5��)x��!"SlC cp�Q�/���Ɵ��$W���9��̶�&H���7ב�]fV��]���ys>������PC�j��YmH�u!+�Is�#G�9�9 �	�A���M"i�(���}�w9��/J�m7K��-� �d��m�w�� ����Vs��>��;ű�>ャ��m�}�V�9������`ۈ��-���&��ZvƓ��)� �O�T�H�@|>��*���P){E�i��9�_�岙]�����Qzۻp��͜U�,�h̊d�o�ӂr.�vn����� ۞�EZ2%��D��'oB��o����T�}]�uR���sh�r�{�7݈h�k�N��}u�Ep���˘"�-l!q@�Wj<v���B ��C���5���Qv7Gc2CQ�ap��|�zX����,�2��m{��/����m�#�A�bE���rUM���kl����-D��қuL���aH�Y��{�8QN�]M
\3�9�����Gڏ�]qP��FY��#��oZR��AI E �C���6:'@�v+h�%avxC�{�i��,��^�ӊ0[�&9�\�1	N�S麗&� d�|c��۰�{Vg��PI�ܭw:X���G�w�����	����s�NP��� ���S�σ��swȄ�:�:ɐ3Z��:��	!1,+� ,�h)���y��#�1�:G�?0�u!�9���|0����a};V%�Ow
����	&}�7��� +��]�����x�������������@��\��ƒ��o�E_���d��Ϊ���jd���X�U����Vo'֥���5��F᭸%��g�]�He�{�xt��t �Z��r��K}��h�v�99��\i�j� ���7��>�{�Qѳ�
d�>��zρ߀-U{&��?0GN߱������4����:��3z�=il'Px�L�t!�O5���`����d[5��еBPgq#.�2|�-�<���R<�~�a&7�_� ��}S�&}�yrن�3Y]p�a{%�i" Z~(��$&�ߓ��q}�di�{9����^p���~I��9煆��簿��y/-���}aEDvݎx�U����JQ�����5X�xS�F����R A �3:���wk	VI"ؠA6�cң66'���*�!�F�lZ�w�(Y����=�hW3R:�7D-�$��j�"4�q^�;�H��+�Sqc�)��Sس���K�C���!ϏEX�1;���E��B<�bΤ�[F�Osk1����dA@�/)���P�$��9d��U��62�!�?�:��";;���\��� ���^(E�����x`<��I�q�������oR��'E�G	����X��|�'}e�m��r{2����OC�b��?���1W��wum#�����m��@u���v�����az�]�bN�GQ�����ٸt���gt��,
=b���N��Wߖ�{u��G����2����eM�p�`7��\@����˩�š_���兖��R}� ����X��� /��պ'Lt��o�:6+O��2�'/> ���ȾxQ�mW�Ћ�_k�T�%��8s��4��ࣤB��B�y��5�p{nnk�*�bhY��Y�f������5g$4�"���y�P��� �ez=�ifZ-����Eo��c�P���T�όg�/.�I�{>�9Y�\�Q7K�s�]}F1"�w��1��}Z�ܻ�i'�'��P�x��gnR�Ԩ=�k*2w�Lnz�����;��s8�P� �����|��S��1���)�";KN$�����`	�]���_�3�A\Zb�ˮ�Pc��?� ����w�����
�6�F30���/�K�o�9���V�5�K�+��	i�;/�#�f���HҲ���maH�:�7����3W���(6�_¶=u�:~���	���"`���a��w�Y��#<�a�zd�����"�e<��U��ٶ�h�K��βo�)�˹!�!W�F��~e������D ���i�M�TE�@*g��뺄�>�8^�.dÌ�s�ɨ!]�m�p/�l5�����JH�F�d�ֿs����b�YБݛ�/)�]��P�*l�\k����j��5��%��)�1��?A���m	��N.}^3ݛ�J�_��5U�H� �D�3᳷��G���~��i�~��Z:s��i��DhGc����Q4[tf��",�{����"�uM��"bj`�{����U�+&s
Lu��&Ym�� ���J���iiL*)a~͈�)V|Rv$�7Amr߮kM�/;5y�LVS���>�w�!�Ց%Mq2 �T,�BڿZ~?ީ-���KU9����+���q����IcSTPAY��9&/�[��/.z���܏�A���ǾoY!�QA���R	d`�V�O9L��]%�v8����\��V��CNU�#���[QY��6/G���� =;-C�nT�;]3Rb~�������T��G��)���ZT�8��'}e�������1ǟ�'���.���ݭ���8�3����~
��\/��9� �鍋���ލ�X�fGj� =�g��)���#���jj:��~��>?]�ư��wa)��w^w�PZ�k��ey@���m �C�1�|�v*��[^ɯ���M�^�+����ir7d����G?��ٟKl����v��P]5���Pm�O �բ0c�bU���
���;�:�E�7X�4�T��0��3��4�T򻂂����[Jw�y�a��IX�Pԛ�$
�D�Wf�o(��X6��N'�|�z�"ж?��e�,$�Cx3�X��*��0U� ,���y�_q����MECf���"��Q�_���̧�����_��^�*[чD���n��]�r���@R]�3�$��=}j![�eؓ.w���)^?ls��LQNEvI�Hyk >�r��޼)��=�~��s�aF������pU�m_�F���?5L�s׌�`*�KfP�[+3Ag k�g�Sv��Iz�m��K��)�!��[C�nOKW��cT��şOW^��9�`[�1��H�o$7Xi���?���kZ�ɰ>��픖�JC�ǥ��!�p�,��J�#��S���)�4�ʉ��>����w��T/ȗ(�<��q�1 ��c���mI���5Q�R��ڊ�,��,���^��+�}�S��4Е���F�?�4���t����hh�ΊJ����	�O+؃:79�4��|���t���E�Z_���_AƟ�T�m����N��Ӥ�լyUN�(h fd*I��=w���
�l�˻/Ӟ0Z�Vˉ?9'�߳����AT	�J�P��1�e1���C78�2�&�^��.ut�����"X-)�@�Rp<y�q�g萉��7�lf���vrR�2�×akHu�p��5�♦[�,a�-��(���E��k��m��l7�|b B�)��M$S�kGc}��%dȌb�.��'���*Pac)�Yt��{�INNЉ�
��t9����NZ��k�qk�%�����`4o�����g�E�'�=�:✏vF\z%��C�T�{�Mݐ�z𓑦�.�o[��Q9�;1�S�̓&6n��X'�c��֊mgQ?YI8���(�*XaMrGS��U�J�\�L���p�Nk�7��c���S�23�a>�Pĕ�I3�cUp]	��E+�z�����@������Ot?�8!�Ŵ�oS0̅�H�}�� �J+Z�c@�U&�0��cL��w��+m��:�h�sLU���_ǚ��^}ồc�O���q���j<_\4I�����f��?�m���U_�n����o��·�@��}T�3@��B�zA�e��xo��t{��=U�f������N����j�o$��m�7+��6P#��d�e��:@ϼ�,-�I����G�(�����	-��w�d��n@�=��PsCL��8�
}8���ёcE�?qk���B�zq/��/���a���<���<�&�����v�}N�v�v�r�Z(�N�*]�j{�qI��	���l(1�$����l2q�v�iK�(�r��^��b4�I~����^��Hk��N�'��?`�AM�)U
��I�J�s؆��5�M�Sӳ���	��/� �6�,�kֶwI==�A�>:c���6A:H�F!�^ ���wd:�Y�2��?�IhZ�rWnp���)�-νJ�M#"�u^�v�]�+���c(S;��cخ��Ԧc�CH�!���̽;���y������]����TO.E]1����uG@�T-/d����4��秔�D�Y�6M�O�p(�3�;v������ӬE�G�4%��xU�"�>;V��&�>���j�o�qp' �	��R��m��A�b}Se<�L�m�!�O��:Uu����۫�m�0\u�[��������CI`�[��z"��/�2��z�ک]?�G��p�����l t7��B:<�g��=��C�I}�W:һ�l"��f������g�)s�M!��`2�\�Z��Ͷ�� <Ρ���� M��&�R'�����4׻����L�����֕�u�5�8w�-��/��'��X����vmҫ-���lÏbA%B`�8nq�4R­�_K��l7yBd_�K��n��M*�"�Y}}#�����J�K�$��3���������+�e�� ��Z�����E꺢c�Ã���6�j"��x��B{��}Y�G�Q���s�{�Fl�{��1)�إՇ���iB���v�axs\�g��F�o�=���n)�22`?n��"
�X;��ss��՛b��������S�T1�d^)*ReK)C�:��ښ�S	�w���Q_�ӮAw��F)6P>u�?�%&�P�t	O@����
�aF"���1bs
TiK�.έԸ�Qܙ����+E�B	�[%�%#����d�+	��h7��7�->��}�(�|���u9(���X�dV���+#���a*^�4"�#w��}��h
�}�N���pČ�1�_�&������Ll���WM]��`H��΄�'g �JC�2��M*�Q�B�g�0��?WY�Sb{�����g����]^�p��l\��۰ը�e7M��}.ӱ�w�� Ibe^d��3�/�Z���EF�\�C��7��p:)%#4ڝ,[?z7��{���s}ٛ���Ӛp�5�/�H}.�DC!J�rRs�bLg�Y2��D)k~�Z�:�Gi��'�_��ȱ����{4�rð��(��,�#�7uH�lfxj1Z��w�U!uks��c�8��g �62� �<��ig�#a�aу�LwV��5�K�Ah�9�	�����y��Q��[���w�S�,�VMlWp���B�h~Z%a-q�jK0�O��r��hz�l���(~c/#At�9���[��.�}��wWk<O��X�o��Q\�����`�&�OZ��=;l%��-�V;g�#V���`�#�%�[�/!������o��'��;��GQ��3-�|����8�,�������GFߑ)�sG���
8��`'�Q`�V4���������.ܾ.�(���ݳ�3B�Z�B]%�|��._�/$��3�����z��ԩ������2g����>\����p����L ]w{��D]w�p�2�B�ڋ��8��@�� �m���D@|=�?�"��������S�����r��l����?u�s��b%ٺfKl�F���I-׋��5����K�O{���)�}�@� �9������s�E<��X��5TT��å��TM�]����J�By۠��g���ϱ?+AD�;��B���S�SR��'�'B�5zn�öZ�-ex�ǃ�H��4��rb0Pԅ,s�7���y,x-q`��(okf"]�"�$qQ׾z�ZE\�]J��A�E���0��9R�	#]����;R䇎?�{=���[�喓i��U���^x�a{s���Qi��I8dk�6^>P��t,5)�ÿ���A���aaBg�t�$p0��_�h�J�5Gg����~*ʁ3f,ޚ���3��kGEr��4�����0K�[)�|�!l�C֚�����e�}�G!�`��WV�9�Đ̬m~HcFC7����9>��?��&���>!<D�ɰ��SC-� ����k�ʴ�A #����H�����2��Òު^����w���/���a�잨 ���)�m��)�Ý�����E�<xŧ�d�9��
�}8���/)"�>r^����O����L����	t�_X�-@O�{��E��O��|4����L����dE=֌���a_���1B�"v�GCS��WE��*U���h�
d�BE���ұ�Ư����˖^��W:�Zh�z�:��'%1��n���I&T�r��+�I�l�k��k��#7�����/��u���w���CQ-�P�@�m2<�Jw�"�E����9c��"Dv�}�2yVDaf.��˦÷��r���G,�D�~��|:��m�e��©b���D��M�	�k"� �gXc�����+#߃T��a~gDY�{�z�N�?
��19�N�zt��z]#q��<���<�o��2�w�E�g�]�:�vap�%W�IC��{"���+`i��nj�c�[�݀9�:&1��'S���&q�t�l�گ12�g҅IS��ܣ��X<*�G�z���wW�π��p��wN��`��U�
�S8�6��(��zQA��b3�*�p0�	�K+�F8��%��������wv?��!(p�~60�c�T�}q���E�ŗ����x�&�Ơ�ޥ��R�+Vٍ��t�n��_|���ߛ�68R���TME���e��_���H�>�c����7�(�!�U��\���6o�^��rCP���O��z/�|�|Y�e�4�xj�rtք��k(:����^k_��Ʈ��kjEG���8�7�����8��/�d6�����u,-��D��KGj��t���$E����[���c۩&=��Pn�DLUUл����J���޳�1�X�;B�!�q[.]i�ǣ�*��n<�R%��Ƨ�ӄ$��}I�3M�r~���i�D]f��{��=��8�س(z�$܅y�'J�q�:i�ꃋM�z^���AaIy�n�;�ȟ] �˷�#�`��!o�^8����Ut��i��J��5����5N+>S�@���o�_� �Y��j��k���IX�AgJc��6|m�@�!�L��"��w�VYȢ���h5�CW����m/@-�v�Ϩ�"�y�^ң>+�O�cc�4ŉ�AةnQ�gvCP(!��N�u;�K����x���XL���(O�>s1��T�Z��@�8/�[_�{��8�������ݒ6h���5���M;�m@���ǰ�ʖ��Gg}D5��g�Б�E濛̢�6W��#o!'��N	ھ����s&���]e�\��hQ�>*���z���Q�5�vۆ1���u�襈�8�G�/����v�����q�hX)�mn)zB_N�XP�Gs��A��Pt�&)� Eߢ,�=�l�DYW�-*�'�D�91ٕ=a䳉4��d{M��X`-�D\���ˈ�;��U�1��<�#�@R��S�䄱�k�v����Lj��н����)aB�(�/����a�$���mM���c~��/�%�Ԥ8iy4�ɚ�ف��y��4�&�LnႼ*,DYxP��]�`�8�0��$*�����Ƒ1�1v�e��[#Z��X�+�bEeޡc�Vg�8���ؖ��Fl:{��FY�R�Q-'s���F����C1K��3Y�R�Vi]�����xNE�g����
�x=���� 2�	�n�j���`;¥s����6Y������2�+SV:�1�0[)���K��u���5]�	���RO_L��A��+���uP_%?
K���W	�n�@;�
?�ZF=W���Gw���K,_a�o��L���+ �	���%V�#�2�J�`�ƫk�c-�y�7N� ������(�|	8#u�5l�J-��6P�,�-����P���#�J��5�����ج��P���٬���T�(��_0E�E�W��bXb��YU�y�� �6}�m	M�ѵ�d�gF�p���W�n�K�]��B�V�?mf]���p�:l�-��k�Y��F!�<p�ӌ#����b �����/���i���`@X\aU5ة$�ǫ %��B�'��?���d���}T$d�}Zr���5J*rHx|�D�.�-^�}����la~��c:�;�i���g������Q�4Q�,��޵��V����uCu�l�.j��ܦ�tU���s�]�so��	 �F��G���ATi�,fatf����V��Z��AcF��d�����^y%�I�.����w?����	Mg�\�
�iBPy~u��-�#�KM�H�����g����c�)A��9:E[])f.�] �?7*P���o��QwR�H��`��O��K�؍S%���Ǳ�mҿ�V2��D�f#^��[�%4�l�2���X̂!l;�Z��Z
��3�
��9�ӹc����
KIG�)�qǼP��8���'�]օ��+��ߟ`�<�[Y�.���ݣ�f��O�3}�ʕ�[��w�x����l������z�7������VIgi��;h�Y��`�3����Xy]PN��Rw�!���1Ąe�&����;PVmV��w�|�{��n�)����C�u�ٶ�rm����s?�ww�|ˠ���3lxʅ�<6����5;�ǭF��O�s����rޘɍ{�ϫ�"J� ��E�\X�<�T��2�`�v��ҙgb�8�(�7�JF.�y��?�x���ǱZl:D� ]��6��<`l�셒Q�'�/�z),��u��e�k׃��N�ή[`4K0KɆ,�W�Z�yG��q��/���f]��"'Q�Q�~2���Ɖ�C��ܘ�$m����夬Y]���k�vR� �Zw=skN[t�����������n�v<s\^�Q��EI��:kց>������)��=�4+�r�Ca|;��pp�_@�X��\�5BS��Bg=*�X�fG����3��Ek�1͉��ગ��#�eKf� )��!�(C��}��� ����؟��{W�B,9I.�'u�H>=R7��~�.S���!�?�~><�E���8mCh�N�*���f	�ZY�#x�-�h�zD��B��zg���M����wJ0�/>�����g�� y�Sd��m'��qƇ?� )�9l�"���,�VC}Ӿ�*����
���f��j��j�I�~���D}n��H5�q�O�>��t]�j��|����E:�hE�q�{_��U�����=g/��W�����K˯U��"h��Sd�[�ӳ���Ǣ�bU/�q����d�Z��5c�'�u��)���T�������9�̕k�7�v'��]��J4Nuj���R?��I�~-=��@ʨ�</弫ݓ>�,���bz,�lr5v�ȸ2	�aa4��&l?��Jg��K�,W��Y���U���Ȃm�6�Vbv�_k<M�k���O���}s�F��>���a���Yj�D{o�XNFBG
-�&9�|��պ��5o,q�4�>���8�oX���E����:X��v|�%�<TC��e{]2P��)���k�����[I�9Z�1z��SzP�&�h�M���X����gǄ�In� � X'�G�����bٿcB�@N�wQ��tek��SsY���3��u��K��3��8��	�{=+��f���vz���ԇK��?a#K!C;)���%0�a���}� �@�M���3�&�|��Y��-��+�դ�p3��i����A�zI������>�֏C��ѝ�`=_�h���-������\�(U����Jao8S�-�c�Lӭ)�!��%��>�eQ�xe��t1�)�&3C��C3��������!j�>T��#�7�Eo�[��}Wd�&�o��2q�-&C��[G_�4�/ԥ�?}W�.,�˙;��,�=:u�Pi%lL��绀�˙1�ˑ	P��������\B!Z�q���4w�^%���|<$����������}D���C�r9������]��`{���8�+�R(uՄ$7����q�miARK�(F/^!�j��It1C�3��΁�#�li�}#���7�_ƴU ����JK���e�5�(�S�푋X�	�#�� �����P�kLr�Isg�A��&ccKv6�����!�Z�}b�w��Y�2�5�:hW��U�-�O���u"e}	^&M0��+t��c���$e|ؤ��\��C��m! b���Y;��UB]����S�w�l��O�XM1�r��>�@�<�/��Ս���r��JpY���\6�����Ggq�;��s�-�l���լ��8tI�Ԧ��p����0��ts����(oc��'vV	�Ќ�}��N+r؝�er��c�4�$LҰ����T��?��a�Bg!u>�ǈ�k���!��'ёͪ�p�>�C����$�z�ܺ�S��GbW��O���	�t-]{��%����=3U�?U4W�8���"�T�s���ֳd�<��MW`(A\Q�h�Cz^�Vn��В�Þ�K�^��RN���i���1�1�&�L�<ȫĳ��b�kǍ#E�/O�Q�HY��nym�P��o���%xi�8d�4����#!xy8���2n{_*�FYsC��w]ݯfÑKթ$����f��������eT���Z^��F�E�!�c�	��s�V�����j���q{oD�Y�}�Q��osl�F�4H�1�/ώ,���ixũ�l}�x)N�gMťKz=��$;2��pn�k� �;�Y�s����oX��r;���S��1��) �K��9�K��ޢ	��㧭��_s�A���<~AP�hh?E�Z��D6�.9����
��FX_�'M'���Kg�(�
H��GR��\�W+��4	��P���#Z&����%�an��^CO�Z�7	'ꛂ�"�(Ǉs��uoc��+��7=�S#����W�O��m�#턜�KΦ���U�3� m� ᦀ��'������c����3V��W���Z�.�$�� � �B�﨟TM`@r���g����:��ʃ��$��b��z��]��Pp�8l�N�&%��u}���f�g���I;�b��T����/:��$j��{Z�\ܲ�؄1A��jL%Ysc�"8?0���~�.�T}��ٛX���y5�D*Hs�GD�[<��㬑�ӉO�n����~7��:D�di���y�>Y"��,�4�ϡ�o�ҟ,��Y�Ou>y|�L�j�����xUhzs�Q��C�>e� �������oi���a��F����V-�1��ZA^��߿���`��y-����m�b#wz�i�b;#Mb��e��B�~�h-g�OK�˃T=f垓��bo��?Hc�D5A��g9��[8�I.+^P�FS2%��wOo��xQ���ê�`]&`O��I�s %�h��&���-VM%���,#9{Q[<��h���q�����;^#��G�;3�3)1�$�n��Y��e&�G�Ll)��o�˘68`� '.� ��{���FE���g�+6.����-��s3���xzc�rҧ��C�@ɦ�ۜ	���w�}��>9(�7�&���g�=��O*t���Q�k�����]�D���3�wr_�ʨVE�N絆3���Ov�
m�bـ��|�-+�)�u� F���_��Pg�Tvrd�����?+U��7T����l�mj�}O��H~5��ЭA�)O1|ܢBA޳�Y��uq�a�)�;F�Er�"X��NT
($�2��-!ޙ��ܻ]�rJ�9cy�~��)ρ�u�{D����J�w�@!߅���'��*z��V�� *en;S��TD�	I	��0F�,)�v�5yb�aqV�ԓ�"�f��E"�Q�^���ۧӿ��fd;/Ƙ�9���y��?dH]�E��ƭ�R�o��u��=��[OE��H���*�*AP�]s?�Q�͉I.��k��2>Ƌe��')�%�Ǐ�F-WRa���j�p��_{Zܽ�U�5=_Vם�*@O�fbZ�v��3�I`k�ݣ�$A��n��~f[K!?�)���!�C�R���Lқo��k��W�O�94�3̢��HTQ7	�`�Ɍ��|��5>W:����]��C�����?>�aA۴��:#3�q1b1���o��9�$������w���/�@������ T�C���m���?ˇc̬ڻaT�~ŝO;���.�&G}n���%;/����L*�م���i�YR���^���*��bO<"Gk�e�ܗ|*vh��^n�<:Es-���5�_R�P���7�Xx'�=�������
	U�h���d;�/�nE��y�����L\�ͮ�Z��A�0(\'��j��n �:��Tz�[���Ͽ�>���ŕ���7IR�W�g�eZu���-˄��-��U@��<��B���{�Gxx�����G�vv#4(2��%a\Z���Q�fۿ���4,�{��4���Hw�<�m�'eHÃb15ўz��M�ֳk�T���I��& ���y1�ʾEa�C�Y��{J<fN��
��S9���0![���q�j�2�i��T�oF��ͭ��ES��N` :s�v��%M�C�I�{����a����f�?�.[M�9)��1��SU��&������̻s���tg�WKI��/ܙmX�ChG�U�&ט��]u*�)NN��
�-AFz�S�:�2^��p-�Ħ��3F�9��	+h�T�{������(�?��!^&g�	� 0]7�s}��$�;�t�����&�R��Ը���+̹$��5�d���ن�G�*B��,���	���B���[�G_m�����:�-���Оn���'U0`��߿o�gy��b{��ޭ�O����3�C�e�m�x`4�t����]p����T��ۥL��H�j{V���.p7<���g0��d7��J:��m�(-��å��vG�t˚��Z��|�裦d��S*=�b�PdƏL��;�[�L3U���5��rn���B��Cq� �|���R<�}����K,�Za�}?���Y%r������P]\�M{�u��U��J(p�a$�蓓��q�"@i��~���^\f U$Io����w���φ�v�?��XE�1�J���3U�����QJ�\��?�5DF�Sd�Ƌ�`��^ ���� �k�uI�,�A��c>�+6�3y�UՖ!ۈV��O�w��Y��C�K�h��5W�׵��R-�H��^c" ��^A��4�F+O˯cَ�ſ�؟ֆԷ�XCy�W!;��DIj;�-�֥ʮ�W�NJ6��?�O_��1���Pӝ@�`O/z �Th��� ��	��AG
6�RJ�+�yB@9;'���Ȓ������V����a���#���c��5�w��k����o�߯'11�	&��m�)P ^e̄�^�X�>��k&� �+ �<��}2u�-��܄�Rr�t��Ѭ�b�����.n���zxz�N��G����
+�$�t�����K���=�]�:qWKD窝֤�o�6�3���?�/���`M�~�`#fz\�M���m�q7��K��y�����R�b����ď{���'�A˝L`<,Ȇ몷&e���#���/������mCӍ�J���@*I%�8_��4c8գ�Ma�>�y�l�ܮ�nW�6*b! YnV���ϝ��#��fJP$ �.�A���<��gk�e
2�`Z
9�apQE[�dc]�~�����;���P"�I{*dY�pQ#E�sG��FGn�M.1
���	��vgi�����v�xw*gZ`^�@�=�Xq�$2c��n挞{2U;x-�s$6e�l����|��=�S��1�(�)��lK�_z�_��k��	�����_�r�A�vԷX�Pϒ�?���!Q��Ο��Y
��SFs����r��r{K�$���!�B�.����+v��	�b�#5����u?��P%�Yy�/P�7į�Ta���`(��s��u
�:��+ˏuW��O�T���Z��C@#(���_��l%��#�(�����٢@M�� oΞ $��W��SoW^`��ŉ�I+<�o�� }na��FtM�Ά�	�g��u�p]��.$�
���8����{]/�kp#�lm���|ȹ��a�2���B妄�Zb6,��ɻ�/����L�ɖ�v\W0�_^��!3,%�B<���?�
X��d.�I#�}J��3��K�O5��Hnx�DT�ų��_����ë�Q�~r�=:�f�i�K��hl���3��')4G.#�J��glh����u9�."�{jL�Φ�ɥU�Dsv�O��7��� ��C�1�mUOi���aj�s�pxiVh�m��AY����L�yH}�?/�=:6w�������M]�����SBƾ�~���-��K�ࠃ�R��9P[�]`��9��c?tA��9Ŋ[].f~��Hn[-@��i��oEx8Q�,��>˻`8V,O&����%�N7�g˚HA�Vh��:C�#VQ[=r���e���"��8��;�����U�3���l���	k��L��!qGw��)�?�F�8;�'i�ޅ'OC�����R���.-�@ݙ(A�n��3�.'����m�2�?���E>�����y)�q��y�U��- ����g���Wd��h�V4]F����3<]HYL���w���c�|�8�a��,S� �m��Ѐ=�|N ���R�9���+�D����r�N��+?�R������G�ln1;�X���<֍5qIҭ<�UO�����>���A�q��<���v�EzX��Te{����I�H�������[����J|eZy������<;��ND�)��s~ ��U���)���'Sbuz�������e�*;��3*�D���0A�,�����wOy}�q�&���Df�L�"]
�Q�^v�k�˧�����Q��[��nɇ0J���;�]��!جRI�����=i�[*%��$R�&S�����s�?�Q��I���k�w�>rI�E�n)̆.������a�����j-p���_�K��n58�/����*�e�f}H'�`�3�*+k���Ϳğ�em��<K��)��c!�Cg��7�]�6^�-\�q�kWJ|9O����H�@7D�6�d�����K����>r��� �8��C޼&�`x�\�M���#���L���p�Jy�t��/=�����w V/�S��.�]�� /����m�<*�-���y��v��o,��È���*�d�}	�%� ���O���>٠z��`(��4��ƺ��0
8�YO�%s&2�"�|���q�R�w��E	f�{�a_���@�X�s�g���A�e���i6U�M}h��d��t�)�����z�Xt�'��Z9]Y�+j'6^5ߟ~�U�T��yм3����o�V���m7����sƀ�u`���}˿cu-s��@�~�<�y�S���bU�X[#�"rv^��2J�ZaW����VW�!�|���,MGT�Tԗ��C��cIm{8���0b�p$����M��k�:���4����W<�J����a��dY`u;{%�#N�zr
c��9���׋�ۏ��q��b�w��j�\o����H"�E�P��:�Ov�l[%��Cf0�{ӖY���Ş욘n[��&9D��1pZ�S0T%&"��j8��*�B�g=J�I�=����X̀G?�O�����辿�����N������!b�S��9�ͨ��k�=�\�3��0	���+C����\�����
����}?�*n!y1���i(08�,m�}B�`�6;���Ms��&I��Or9��g�+�X��*�_��p��K��E#����^F=���ݞ�V��_șy,V�Ug���Z����қU�����T*o��£"��8�r��ˮّ-ie�:nx[�
t�BT㜨���g��ϻ�ۀ�8��*j�d��Y�7�:��"��:w�d|g��%z0Ϩ�$-\hG���nG*�u��uMb�����O;�Z��=ppLP_��Lf����ko�g������	'[BW+�q��n+?���^�'��<'k��*ǧ����DL}:=D�pr��W���B]�Z�{\a�����ad�(k��$�I�X��qG{i7���Sh^��G�:Ij�`�L���B���1�3��lvrݕ�JU�;��zf�J�>&�:�5��qS?�+�����Y�� ���{�Ck­�I�'Aw�Cc[16-�1���a!�ր�3]%wP]Y���+�h�'WWZ)!�> �-�a
ϹD�"��^\�a�{+*�gc8��Z�9ؚ�K�1�C4\�!V����;\��ˊ��I��I�0�"��O�M1��ˇ�@a��/P9?����F� ����+�6��妮/�;bl��c���9Ȭ����3~�
U��P�����p�k��L����o�'�+�	+Ug�s'��N>�e���Y�8Oy��&��T��������7ut������X�#�/�����f���ȸ��z8|�IC�GXz�Ŵ��?�ot#*D���Sз=i�;�5��W��5�X����!��E@�����aM�`m�\4�˹�?�� ��Ƌ�T����õR�ae�՚��Sק�\��Lۓ��a2��a��2��_6/�{���ξ�̜m�u�%��{W�%��m8ZQ4��"�K�[�YUYy.Z���Kn��A*�`rYi���-b������߾$��o�b�w���2e0�l�Z�r��|�E�(c8ϲ��G�ָ����}��{��Y.4dQ�%s"3AFX�<~��1���D3����i�Q�b��x߿fg��#��&=�� ��b�2ǲn���A;S!�s_����
��?�C�+S���1U�)PGK���&���B�	����c�z_}�
A���2S}P��?�zߝ�}X����Qn
pLF������vg�KݯS�@WC�=H��s�+1�6	�O���`#F������SF�T���e97p� ,(�
�(}�P�Uu����L��З��ɚ_#J�Mr�9<#c����_0��X��3�t��ܼb���������m�0� �
W����'}�dě��Y� X��hM�}����gWvȺ+J����,�����/4����]ʭ�p�o�lȒ�ۜ��3α����)���3bѰ����@/����O�ɱ�\���:���\@%�2͝ޭ?�L㒕�!�dhW}�})���ӆ}y5�"Hi&SD���^�v��L߉E@����~��X:z,bi�Č/����ɡCs4¬��%h���uO����u4��}�j,>���U�9sQ���$Lt|Y �^���(�iӟ�a���KV��}+�*ATtd�u�|��RLycYP��0��9w�O՘��MX+
�B�B���~Ɓ�-]�dK�چ�ʇ���,��X�a����c���A��\9��/[.�����({w�ċ�o ^<Q��A�P`�HOFqB��E%�T�����V����}#�P�[x�%�=�X���=̓��;��J�S2=,�3�_�[�¤��q��=�G2:�)5,8���8Wa'�Bq��B#���şq7��.�.H#�����I�<3.����h��T�������L�޴w�m�Q���ugzV�l��l��6�!4B�	�m]㍯���w(�����C�|�0Ӭ)��m'�����e|���P��6���p��3r�ʜ�r>Y8�Ӊ(?�o����k�&'^l���3���w�5�˭7�}O�춢��i�����٫��㱘E�Z�X���T���Ñϩ�cmm�|sU�Ɏ}��pJ��y�ܤP!�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�&ڜ4�z^�27лXo��R�|n�?S4��{2�в��3�i��R����@��r����>x�<%Vֱ)#�׳��'Z[�Ϲ,@"����4����Z��mg�U�f��Go�����X"�q���D4�y���O|�:�G��oT.�t�U���8 N+[II��
U�v|#r!��HQ�I1���7 �dI -/�,.y��1#r�.$�����S�����ڮs�
օ8�9� ���q� :n��Hm�"���z;/��Dt����L�w���;V�ȶH�Y�m?�ڈ?�9
���̗�������2A���5�]�d7�p�Ƣ��D�� dS��\�������E���RUA}�ŀ����6����d�\F&��n�Ou�m��VЎT����ɍ��J�I��rLA�P��R;�v�Vd�;�r�h������x���f/�{�h�ҩPwd(��nիf-�ab�|�1�vB��� ����6�w�c�b��K磘$��޳�s��
*��s���]
F���_�zy1&�i4�=T�A��	�Z�r���S��O�-au�������;\#��	e@��r���ڞ܄��6#(���g�g�C<b��;��5uJ��P��w�YZM����qNO^x_�=�"�&m�������f=�t��kl���_�s� �t�p�&����o�8v��W���IS!\�s��/�*����؄gM�����#�g�ťZn��q��|�׻�_�Mk�I� }6B�`]�'�/èf�1�T�?��%춐���{Q4�!WUP�C't�,�{y�!5��1O���Ć4���B����J���~��w9���p���Ft�[4R<�-�k��(��4�}s�f*�Sf=�-`� �6� R�Jo`�I-1�1�iݵ��`�.��&t�V�zD=��9�%B�'�#�z �E[z2E�����!������Bp�٧{4TL��<��6^��U-�}��2�l��?� cgiC*2 ��};A���.�G�����v�W5�Ji��ˮ)�A;��@��?�C�VSD&������	�9��4'(�HPh$:�T�CP�ȗ��짲T�y}��^�fPV�lu#����>A��S9勫��6MX��PZ���j��I3�Q�rxs�Ъ�;t{�QM�[�ˣp�%��i��=���Y�IT�`�C����h�����x�@�{�S�L��uE�F^/C�����<�3�����"E�h�$dQ��E�^KpzC���p^ԡ��4R��nY��T�=$0���N�}���p���c�t���0ݯeBJBU�VWsgh��+�I�Î�J7ęW|q�Vmu_SI��в�[8w�7<$�Y��g*l�oM��_�֦d�z�74��>9M�����l�`q�ו���C�k��|�'6y+9�~�V��Pr�q>2�2P��^���g�ڏZ؋�r�l�> G����m�)K��¨e�A�$�L��e.&� m�E�jY���L�_z�T'[O������>}�sA�QD�����H@��zb��ߴ2Ō��1+�y��d�b����9��uu��JtXTps���bQ!�Ԗ�cytr�f_�(E���.6��ާ��� �syD��<{c�|� �."�kta@)(V_����^�)��{{�  |R;"h��N�UU�XSU��5+�C��̘y32(�ݞ�|נU.>��`�'ۦy&�V$/�Q��N�7�=�_G��P��+���<�>�]r:/-�4l*2�N�=��<g	X�$�;��<Ιn�0:�jF�����ḏ��1�	��N�B�ۘ�DZS㠔�䟅喵��{k$�6غ�q����Gؑ����qIIh��j5:����s� P����-�s���߂�����JA��+M8��d������A�jLؗ����[�J�L���:�\Ƿ����sNZ��y��<*g���D�Ϥ(%��q?2�|ͤu��I-��62�߸�����_�\q��L�C(�*n�K�g�Lֹ8��k{��?��a�/�l1X]&5��N�Kc�W��lD�%-�\?�%f�^f~9XӶ�}A�#���gI�Jٲ�ؓ���%YSw�Z���c���O��������D�އ���c������-�t&�� �*Q%~0�5��"$O�`<�(�1��ã^}��f�*��w�Jى^�Ȍ��'Lm*����#|��|]�f,�K�f�x�d��6�D�D��a�?P�Į�8^������;��;�zΏf����s�� �RG�F�fX��=�MR���_���^Cb�g��7�K:p%�v0�,�e��M�ZtBގ�ssg���l�eԹ8J'��e�A�B)��Yt ��@Ś���_΃�./�4A�GƆ꤇�hB��Or��<���9�����@uH(�C-���̠\�EmLm�,@�*��y^6�6(�M"M*gd��r�-���ec^�+�C�Ժ��f�ؒ�W��ϋ3BP������~�k����3���Q� �o�ψ��ԥ��!�ӏ`� ��:�jE�)�����n6�TMj�^6����l3��z��|4T{v���4�f鋄s6cMk�V�H�V>g��c�51�k���Y����ՇQ���VW]6Z���+��1׵���"��3���)�.j:���]�!�"�Y/pCW.܅�7�g<�&���44O���<�ۛB��Dу�e�Zn7�-e<�:���0���P�_�nDs�k�����]W�xԸ�ʉ��  �:�rV۽��q?b�~��/���%"�&>���_Ұ	��ϥ����$�����9lp���=3�*� ��[w��_����ӭ����|�I5�R��3��	��t����wI&��Le�� ��R�?��ߎd2�t�|��.�͸cr��Q�b�,���0�Uy�6;:�r��JG$Q���>ih�I@�g��y�<��9�K���ʔC�Si�<Tv��Z%�����c7 ZO`B�q%1S�J������N��d��V-�	n�r4`@I�Oί�oQ�fݺ�\`�_Rt-l*��e��D��4�-ĺ���}x�8�"̗�Ek��q ?�5�����iMfY� ��0�E{��@ ��S���Ʀ*ee��އn��Y��x��4�&�ﲳ��2��.���L�n�W�S����pj��_.�Y�iu��;--@�1�ڎ�́>_��4֫0��?�}�;�-Z0��&�"9@�i�Y��Z��Bg��hf	e�oq,����"�~�� � 4m���y?|�TI��O|o�1t��a�)�g ȹ�I�
O��|I�P!|d\��C3�����7z^�Iڤ��&��Th��=G #,U�$�W���h�.@y�alg��0����lU#=�.���u��4����k��>��	0��mU�)%����!=����k��D���"�-���M�r�B�X�����y�8����Q�;l\k�.��rW��Gq�ŝ�)�|�h�챱0��r)��p�1��:hv��5U�a>��t��?�瑩���{�cE�:�����k�I��>��f#7<P_A�o�A'�؝�9ε�����y�@pb��L&eQƦ`ҏ�����d�`*XW;���ou�P  e��O*/<7�7�6?��|����s&W�L�h]���tL��m���?�1�D�*� �J�xK��R�sW�L����}�D��P�٦�
���Lu�^^���G�j��S��o&ۦ�kk�9Ѹ̏���] @=��"B����x�dEū=�ͦ�c�� �9%��j�!M���jZ3��;�f����Β��,I��&Cڧ5��(��Z�����P1l��!�<ʴ���Ֆ3流��+��Έ8yu��J�B.���Y	?F�F�%����/o�s.�jg(ƽ�-S��҂�a[�s\������O� ���?T��h	�C[�e����g��l�H'5l��v�ѿh���MT��ZY du�f��!85o�t�X~�o9�>�W<[�$�¦['�P��"�gs�?��bl=��NZa��m��
��X��X�m��O�mfG��Z���v
��;;��e�.�|��1=:Ϸ���׌�30v�b[�����ާN�^��q��â��H�#W'�����3`޷o��{�i��bU���n*
�25���R�b#�o�Kn���w�{���U�*2�p�z�y<(�}ەz�������wy3|����
�ʫ8QFK$���n��)B��������e,�?�Q�M{�R_�#pO��D�+;��,��9�h��@���e�ލ8�ٿ�#+Ԫư\b�}N��<�27G��F
/q8l��]���7L)=�H��<s���+��]��r}1�3 ���,�`';�-����3��$rC��,��I�\�%��(�դ�1�ep�H��!>z��
�ŉ���~�6�]��F1=��<@�꾒�D��@H
�$����A�i}�F���+a5�X�;w���=#Aԕ��u�k+���E��Pom\�/���(�{�r���2��������pۢ1�m��2�6?j��>cG[�Ȧ7����_�s_��JT�eu(GPZ�L\��AS��ڏ�!q���w<�T�B��:����>����l[X�%l!�Yf����ecrT�E�)����H��X���Ь��ݙ%����XӖ�����i�+M�Vj
+��pb����-_.�����+b��xCq�Մw�"vP��`%�lOG�<c0�'�bt����7t���M���*��d	S��ߴR��~I@��JbM���p8a_�>N���-���'�w�f�Ž��yӶ[iW�`_�c�q�d�sl-���7�(�\JG��p�;ZM�c��p�;t��$=��~��pꅦ�;�o
�)a�c����۫�[d=bM�V}�R�1|.�(Ԙ3�aʿ��/��ܝGZ{�$�-EH?S�S�H�i8���!��[}����$l�h��w�ȣ1�E��~3@0߅�@�Z��6�S�Þ�B��n��[$̼0�~o��cb
�
}!�����Sq{y������\P6��\`�E�ץ<ާ���I�W��6Jj�-Wɶ��2˻�� ��K>j� w��ve,�O߾ "&�2{a3���D��[㡿K�ڙ�-z��6���s���l�[cYy����L���1��Z@�� ��F�G~{]Y`b8�n=+�����g�3:�Q4cˊ���B�����]�@;<)� Y3[�������O>D~�N6b@ �eD�H�,�1-ij���{ĳLm��n�ߧV�	 p�'Fh�t��{��|MU�x#�K�f���k��?���+��͙9ﮙx<aE��ǂ����
���lچ�[N(e2�N��{�����������&I��#�yuNƛ�3�q�`U�g醨�<:I�+��,� ��V����F�uW�8�(y_�Xz�p�:���s���`�u��z:���GϨ�F��O"���N"�B�g��)��$���6\Ȃ�}�8O�ƌT���r��,�z)>��k[\@�Q����m����%���}�)���n#�����z�=�}"� �b�&�SF��"7T���PZE�~��n��1[U����O�i��oP�5�����j,�j�ߺKu9�7�1�6#f�f�𮢑|�3��8�ϊjM8���|���t�G���"��� z����	f�NH�N��qF>R�q�i)i��DV�>�5���+p�}�`f�%�*c<�H�.��kFҪl�w�����0`�dO�}zx�]��l�kxm���i!v|#�E2���]M�x'p���
�;i0��xQ�u�EE�
���n��������;���7�����iz,7��M�D^\R$I9�qɈ#�]v
�Nh/��$,A(��i�'��`ߝ]UA�L'B�m��՜�>�����MJ��,�C��\����k$Rh��8�&3��8�b�7���@�JX^�%��=䏜n��T�J+���)�r����f�,:|���찭� �rv2�_G~�0���v�Z�\:�*�>޺Ln���.씖(H�K�U��4�O��ٜ�g���a�C�"����9��&�t�L�o�1BO讐aҦz�
3+)����;)�<38��4�� +~�HP�b�;��;ҙ��1��{ L����VR[H���m�T��+�9E��2��|�w(ڵ�/��G���N���p�΢�g5�Cn�S ,�e�����$����8�A�w"�NH��Yx��u�}�?fe�B�
��"m�,�V3���K�ɰ2���ϛ�Œ�Sa�B�a�y��V���;�\h����+����?7Q��'��F(K��������}Bf��t�[�%q�����Bu��#�
Ӗ[���}�B�fUO$e�N�JW��|���
�R	o?,��s��\d��ƅ4��WޖN\������n2�1��I�OԆdgՌ	W������xו���&��1���v��f�� ��	��_-0��J�C����е���PϠ6��E�����]w
��-h�'D&�g�=�� �n`�	�B�r&�[S�����Q��:���Wi��)
��%@U	�r����jY�>�L#u�`�T�G��FP��������P�G�$n�Z��;����qۖ�^���=��r&�ޘ���Kn�����kYS��쒪s��tVL>&>N3s�8#�	W���6�w!��rs&�����'�R6���M}�َ	��Tb���	�8m�q����"9��eM�L%��#�(혶'��_�3�c���	? &8�c�Gm�4t<�U�'�'���,�K�yJ뙸�(M2o��T��4t���Q��&���e��U^S���A��Fd_S�Hr�Rɏ��.������s��F� ��z�\��Љ����w.M`vZ�-���ɗ,�B���{�T� ��zq;��~TBe�#�e�ő'z'��=���:��aj���B�ʧ��T��$��,����Y<���>۔�p;�M�o pu�i�IA*�r�}��A4�..���T��@�WBЦi�O��v�.;��Ⱥ�]C��D�F��t�=���N��'u�lPU�����C9�Z�d㦕YvIT��x��^^�nPC�nu�nD�k�Aݢ��$f��3����I!���p�aA�~�Cx@%êhDS�.���$ [<�z�%F$)�#$y���I���P�.ќ�ޒ��e�;�R��y��u�N^����
���{�s���w�k"�cQ�QT�i��^�ϥC�#Xp�"����;�Y����j��0�+������暈|ưG����<�J4��#�����8��p7�J���Wi��V��4_����n�d�w�$t_��^"�lr�@��[_��d��̱�(�О9�
O�#�8l�"}M��J�����gmx'Cw�9�ֈ~������z��P=�k���J-�8Μ��i� 4���
�]���e l�$�Ĕ�2}.s�{ �E9!�n��~zW�[)��m���.뗿`w[��7@��YH��z���$u�Y��+�"R�Q�l�n�	�f3s�B�����XaG��1b��/ԃ2Ty��f��E�.�bW��L�v��Mt3sf$h��{4_	|��=.�nx��@�r�_�!��,)�{ڐ �z��+���5�U��k����q|���gE���y �>�J��ÉzEU�B I� 'Ȋ&3�M/��ڰ�?��fG
	:��PA��:�<���]��/0��49�X���2��Y	�#ʈO�<���%�=���]s��N@�I	��N �Nۅ~�Z�#U�;��l�ϖ"�{x�5��P�ǾA��ҟё��P�h~��5���౽�%��G8Q�`���!� x=�PbJ���+Zܽ����R珟ӗ���$���B"J����P\tG�e
v�`}�W�ŗiȡ��2����(2kq�+�2��R�bR�I���6_������i��_���q1h�b�PC^0�#��K׿�L���%����D^a�/��XJ,W�wEK��МGf��a�\Lh%��fZ�5X�Y }��#���gI��۲�&��	�%�^�͑-����+�������
��P���qĩgpcH1���/-t�'�UQvTtQ�	ŐB���>4��u�z�~��NK��L{}j�Zf�҈Ǆ���6�H�[�c�*�C�P��I�5f�IK���xN9���76�1N�aLqE��8+���x��k���=����� ��oRC��D]����J�a�â�R8X�_���^��g���L�A���,OQ˚O�t/i;� �g,��l��.�������oA]�?�S9tH�3�p�qK嘄/��=�/�X�A��7 S�-y�l�:&�`J��|���ૃf��ͬ(��ɐ��Ü�)��m��?,M���-�<6�[�(�LM�C�������Y�x�jckF������F��.S���.ϸ~�P����x�:�삔d��3]��>�����ϵz�rƴ!)�`�� �Z��j�9����f��;nc�uM7��6\և������N��}�{c]��8�����6�n�ڥ�Hy��gK��P��1Ey������􏻔�b�]���1A��~�>�S"&�:�P���X���y]��"]��/]��.iG7����IW��Ы#'�)O�H����vRӖ��V�i2PV�|�5���n�GE����r�hc)6K��'ks��l���J�����0��O�(x~f0�gkLp����+���l|�}E����i�xL��5�
�ti��k��%³�?E�"
>�o[P2$0��Z���5P7��I�N���,$�,M�"�/�$�.q6�ʰjR����Ӻ]�T,.������,ͤ�*G���R�����Wr>夵��g0Jh9�Ӭ���)
�}ۅk1�9���4�s@E�%uÁ�v:�mƴX+�E%�<�䜯��t�S��T��i�#�r߅��3=:���~�oҁrh}��P
~�?ʇ�V�'��:!ʘ�Kk�L����2󔃶/���.��6��	�	��3XaI�4"Xהu7�9+��&�����t
�O��
a�댦ǿ"3�@����;V��< �u� �S�A�� �[�>�ZH=9��ȽU;��8��
O�}��L�2>z��V�w8H��rm���X<�9ڛ��\=���Ew]w�������\���4�p��t�|U=b��ʲSm���Rї�X��Q����%AM✀[ ��2e����,?��ρَ��mw�AV�oW���M�]I1�R��;s�P�o�7�F�1V4��;�=�he�x}���R�Q=$� ��(���xmش��[}�6���q��!��k��BB�o��0�
@u��#zS}�5�BJ�O�N��(Wس� 
HNdoLt�6${�_Ud��ۅ� VW�E\y�� <�{X214�S��dT\�	�C������E�t�;"��Ɖ1s�v�{��~����2����E[��Y��b��"W:�a[�!��r1����8]�y֊[���&T����=8�e����	wu�r�J�S��-凭���&��RĶU�ĿG�*@"��r�T���Aw��%#�XP�A�1�]�l�4�3��"�$�rP�<�у�Z�Z���.�qhi\^Ҽ�=�+&G�h�����]FkF%��y�Rs�}t#s(&�Nb��8���W=�ɀ#�!v'DsS���Ĕ~ſS��wM*�A�Vl��An�t��e(�qm	��V]-�e�M�~9r�ai^z_�'�t�� q�.�?k�󀋔)4a��Uj+�'��,�f4y�_��+�߲�¡k�4�V�\���SX�2cΎ��p��D��Z�F��5�RV,�[ރܹ�U4s�S����g�Ǡ����F�:<+ۤ:�`C�}-���Ъ����ȬE� �&!��z�$��ӌ�B�M6#�[�rI?z�� ���� ��(�O��BJ	�����T���֑���歕���v��yK�ـ }�i\�$*̃Ĝjt�A�^�.E]9Q����JWO��iS���E�;�$���C5&�D�I�����#r���'�P�PB�5�n��Cf��1cɕ��T���%�}^�D6P0Q*u=�l�G��A���-�=��}����▼���u������x�}���\�O���gD[�1G��%�}�P�H�r�_I.�%�]�Q�I=]�fCR'ᩕn���g�u�0U^	sѿ1�(�9F�k�d\�"_���~��6�L^%�C�{�p�=�,�V����Y����	z0������켗�ʽ���������Ɂ�Jaᅩ��AF��EkۅKtJ��WV�}V��_����;U��s�w�J�$!�	ë��l_�č/�i_:��d�������9��<�pJ�l��a��w�a�����'P��9n~8���9܊�B�8��^��ؘ�����U��� !��'|9k)�^/Oe�A�$�G���a�.��� �ɷE�b������zĎ"[6�|��@�{bQ�M�C�k�4���H�J�z<���!p��:+>� �>�����&Ǔ`'��e�KXn�@�t-2b�8��pͲy��f�fEL��.�3�����#a���sS\��'�{aF�|soU.��.��@�(_Q����4)���{J�" ��n͘~�&3Uen��X8�^�n�2E�#�y�t��4�Ö(|U��,�`�'���&��/ c�������Gt��[e�@�~<�k(]8:>/]�04aH�(�����	��k�ծ�<� �r)�j��*�Q���]��%	I�Nm0��rd�Z4������9����.{�]y��4k��G�"���=��B$hK��5I
� @ɽZf������M�y?��MG�c�J�+g84�e�� �����Q��v��Qm�gt�Jcx����U\!B���ZV�M�������Q��l���[5/(?��q_��20L�OIFIG�6���y�=�֚�_�Rhq����ZC�b°7K�Lp����E���T�,/60%X7]��a�K����imD��@�\Y5%��f�;X�'�}[z��&�IjE���4����%���Ӆ��\���G�i�U��j��
{�V��c�oj}��-�g�?�C��Q�?�O��|�&���gG)�K�J��b}7�4fb&�ǑOs��b2���*��}s��@�f��K�W"x�x3��l�-�a�-��`�8��_[�!�T�����) ��||%�i�Rp�@����2�=�W���p�?R��+_��b^]D,gD����J	a��z,�����{]t㕍_OgY�fl�08�h��>A
?�5}ut�P�U\4��e���]?�/��AY�]��&q����:g�d-���+�&I�X�/���(v2��������m&9�,Z2�ڣ;6|�(�v�MD�Z�):v�S�����cx�z�����_cjǲ�|�q���崗P����������)73���+;����;��%��??�!�M`��ѩ��j�P=������gn��%MN6Ʌ��қ��>�l���{P����9���A��}6=;J���H&#�gU\
�=,1���1ãe��ayk�zP]��5�~O��k�o���^"S#�b�������];b�"��/J,.�"7�D<��@���ϠO+����ޛ��*D�|`e�nx7�ı<f�≉� � v�u`m���!DM��hW�q�
�Q֞��v�+R��V��db�v뉍쩛מ ���忰c���?ON�t]��h����:pC8�=g��Cŵ�|Q"��ې��� ��wR��A3	s��HK��d~�Qd���H�xF7 or(Rl7b����d���
���6��S�EE%��J����U0�yRG:����$ւ���~	�(�E>�9�G<cqY�Aɞ���+�V몇��3��!4�	i�വ� �d�u����H@9>�C�3ٴF����s�D̾5���Nt�C@�eӇҪYH1kcɚ��{�5S�\��OW�ߥgz��0=��o�h����3��@��~@��5�q�i���@�N��O���T�4�ɬ���2�ٽ�Zs���Db*"�L�P�Z���g�Ӗf��o����"�;���N4�)�ӗ7|�P�_��ol*%t������ f��Ia=
m��|'��!S�܍�aH���z~73VI8H�DB2`J��:#��i$�����w
���Q�RR#0��8чR#�f����u��4�(���_�>�x0��U6��\��![����wk.�z�� ·P��C��#+נ�eX�'���5��p���;��B� r�^��%�1���^)�+h�w����BrG���N�_�.�Sv[��U0p�>v��� �ޱM���3�A1s�-O��gNu>r�J#�=�P�o�gܘ��?9l�8���p�:�`�e�c+�~6��l}ҽ�*��1��Y��M�^��>e�w>*2�7��6���?�f��� �@W�;�cs��UL���m(�(?O�qD:����9��Jo,�.ڑuL������l�n�-�����x��O^9�'��'�jD������aq�e
ɋ��*^����` V���!��ʈx���E�a��uS�Q��Ϊ �0%?*+��V��|�Z>e;]�x��s�
#���Xϧ���(��Zi;T���l�������T�4���d� _h�qe:8���9pBL�z���Y��F��%^?�Go��2�ȫ��ہ S���� .)[v%\$�����Ք ��?r�"h��R	���[?'��-l8�Ela�5��yv��h{SJ�����C�Y>�U�D�ݣ���5�q��v �=�Y�D����9�;��' y�Ԁ�{sjk.�=�X����7{auN����@�H5�v��e���l��.�;dfv�	�٫3�-��.��`�?:m{��O�*V�v��[[.CƈU�T�l�d�<��q�&e� u5Hr��0ԉ0�g���ĳЪ�W�	KbbPr�12*�yN�&��bA��o��n]��wF-���2�*	��m<���۳���j�ݥ�}�wk�W|�E�蔭h�Q��l��LdѽW:�3NHR �%`Z~�A�bӦq��y^	[s=��T&>ʼ��n^���WޥuHk�P��<=s)��t:�"&�]��nr8�r�Wԗʀ���!�(ss����GsŶi���teM�9���9�����������q���Mz�� �M|��	�)��.�'0/Z�r��%,�?� ����+�[4�ɭU�ao'�,��ay��Y�� �w��8Ǥ4j%iٳ/�ƊL�I�ю�!��͵���,FH�ӬG�R��ےm���|��Ss����dI9�^J��q���������`Z��-������+��_�@�w �x�z�A���P^B���#��ٵ)*5zc�҇.�e9��Q��fsOBAWi�l��T]P��m0&�gd½=N��,�㋶�.N Tىi*�*c���lMAf�.|O&hf����W&��i
T��Z2�;�1����Cl_1Dשe��[F��3
��'Y�gP��:�ũ�C�Yv�H�9��Y=T�e^�F^B2P�ޭu�b�~IjA�M)�$,)��WG8d�-���E��i�D�⺯x$t���o�e��b��[ ��g$I%*v��Jc����I%0*�4	�� V}��r0�Ij��߫���u�S$^ ����u,�ߪ��c���"��]��r�M&�^g�C��2po�M��|�p��Yj�7��3]0�
���C�n*��+CƔ���F��� (dJ�R��z8���ey���Jh��W���V��_�Zg�R[��w�+$��O�B�l֩x��A�_q�d�t��/t���o9^�B�d�l \�1=Z��	h����˸�''/�9%��~�L��yoG�4����O�˦�؜����N� �H��~��p?˘u�+e��b$w�8�y'.W	 V�+Es��!���u�z�S[(�Ѡ����@��-�U;H��z3�nߥlD��'�+��Ե�G�R�B��	��&��\�rXEB�+�Yb�<���Chy�if� SEc�(.��ϣ֡ڔ��1��s�Y��~g:{�}]|��.��\�A@:#B_�^��/b^)3{�� �	�͏f��U����Q��������L�y���#��m��U?;�- ',,�&�B/7oi�������G�(��m���Y<�l]��/�K�4��,�u7	i���l�<�6�	"Ρ�-�A�T�� ���se	 h?N�$�鋃Z��j�1���P�;��9�{\ǝ�G�Ǣ�-�6Ѿ��T��k�hb(�5[H�אɽ���+q���f#����R�z[J��+>p�� ��/7�M����#�~�JZ��� �\�;�I����^�;�)��N����q�R\h(��qD�2�#��I��6�C6��t����_p?~q��q�F��CyC7���K;�L�����z���(��h�/�UnX�5�[H�K���Ѐ�D��|�\0��%wuf>!X$�m}���]�I����[S�~5�%j\��F��JCl��j�Iɐ�lO���'ϓ�4�c,���R-X��v�'ZQ����&���3/��r��;㱢C�T�k}N�[fY~��h�ٚ���1�x +*����{�-�f�HK��Cx�q|�g|���/fa04�U��8��Rl"����LPu���'��J�n!�R�u�����)��.���'#9R�U_��^�cdg{ ���l�A}�g��,����~��t��A���g��l���	�?���A�S��(>te�.C�V̌�|+��T��/�H�A�,�y���P����D�5����������q��(�^��t��'?���m�,1����!6�K(3*�M���`���gB�܉ecO"�T�.����)0?��	��i�P��'�ܓP�ol[�� �3A�ܢ������!R�V��!��(`����Q6jv��\,Q��on��M�6�1���Ǝ������{��m�����!�ʽ^64�a��H�o`g�?䐴cB1)7��h��|]��X3&��rb]G��m��T�7m�"�:��4`p���R�߉�]�<i"A8�/�fv.M�7.����e����O���MU��s��D"h�eMɜ7ja<}	���_.��#p,�JҐK�D�4a�O*�֨�K�)�4��o���K5}V�;��ibY����F��5'��d9��`^�����{��ݴ�M�X�y�pZ�
=K0����l�u�2��D���#�����NR���3༳���V��,)����A )��N# ���Rc)q�в�dC3+p����)G�|�U�� ����0��%y	Z�:����r5Q#�>��&��q��g�ԓy�9�"`nK֊ ���S� UT'�+�`�;p��=71!n`�m�|S;�ب�C���dz�-�{n*��`�������,�Q1����U�P[-}<&�%)��?tq��������o�N�)Ol̨Z�k(��q/D5vz�V@M��Y��h����V���G�d�H���g��Z�n���Ҥ��E��&�Ƴ�h2"�⛼�� nΊ^S�A(������?Ȫ�i�d���x
@g�Q�V�r,������^�Ȑ���@Z�| ���"
�81Z�j"�Z�̂g'��fz�iozx�2�"�t���f�4~k�Ӫ�{|@�ǝ2��o�'t���� ���IH
���|�E!�>��B���t���9�7k��I�T%�WO��`���I#��9$D�v��yy���r��6 302Mm�ZP#��4����u��~4���|��>���0 q�U	���!�[Ċ��%k�Z���!��ʷ��~�~ξ����9�X1�Ȋun�)�Ԝ�.;��d��_�v�X���v��)�9$h�C!�A�rZ�$������v��U��>i퀟s��� ]��ZՃ��F���F
����>e&�#P�Ppx%o�ZJ�)�k9?��?>4c��𩜳�]eb�즑���ߕj�ծ�*�1�t���@�c�A��e���*E�%7F��6s��?�������umW҈y�k���ZL/��m�U�?���D�y%��ٚ�i�k��ڤ��LY 5�h�ޟ�@�hʦt��칧�n�^L��3L�j���?��� S�X0�p����̸��<H �&����� [�xB�E��=��lͷ���vC /��%#�����j��Z��;r�����/�p�}�S��t;��-�(~C�Z\*���ҿl�V��� �N���Fߧ~󬓞[�d��8jX���_B_fY�`��Yz2�F!��%��v�oԷ��{)�o���(C ;��� ���<�	&`HD?-����>"��'@�MM�%�(�A=z�����B/{/#�='�Wt:zQ\���s��|J�=pTJ�B�����NT����[Τ������<����p�_�� ±niA*Qu����_A��J.��iV�R�IW�>�i8��H�m;���g�C���DŪ���zv�h(>�[�'G�jPg[��3%jC�B��6��kF@TD�
r^0U�PUr�u�⬀A�j����
�uV��$���z��>N�@�x�|�z�;�d���%�[� T%�3�����w1�Iӆ9��5��.���rgwG��Z���%�u䚕^��\0����q+���_"$�ϫ�ᠬ;{�^�Y�C�p�菱!a�~[Y؞ӫ��r0�m���F����ۅ��/Ƃ"2���ݎ��J�]������o����r~JVEW{ �VL�_�}�@�<vr�w;A$+�0al��$����_��Ed��Y���d�9�)����l�-*�Dh���6�⮌�y��'�=9Sg*~��oɬ+�P���";��}]�9C�������� F�����c��
�cA]e2��$�����.E� �
E�$`�O�*�:�zi�Y[{����f� ��rJ`�0m�ǃ9�H��z����r��;�+Í��clT��U����`��i
�_X��ΡY��bp�ԕ��ySyfʛEQ�.�R��=p�E��Csx͋��P{{Ɣ�|x�6.�P3���@h!_�"�ݣ�)q|�{��� ���=ϑ�]�AUJI�w#u��	E����I�wy����\Z����Um���'�	�&��/ep����⼎xG\Â�@U����A<�0R]���/�4P��w<��EA	�(@�Z�M<�,�wѧ��&h�/��`��U*�	.��N���ۗ�vZ���_���>	��4�i{���u�>ǐ���村e c�0��hP�?5����Ec?�?���H�r��|]��=��hȰJ���+�Ч�J]͂�cq���c�I�Y���dllJqů�k\���7�$�r��ũE0��qd�q�� (�7�qDN�2�s��ta�I�66��~'��{=b_�I�q��&�4��C'_��u�KiM�LuW��7��:���u/���X\���ggK"��n9s����\�(%�f,�+X�>�} v��`\IoF^��:����%��u��!���!�}���wr��Z���`d=���;��c x�IR-�ڣ���JH\�Q�j��T!�a"�l�]�l^���}<y�f��������L��&�*b����;ӴCf�/�K��x�륗U<��C��a�򼳃��8��V Q��fE6�z�ή��������"GRդ���׶���U9=R
��_�;^"�g�}&踏�����t,�Y��lj�tAށ�R�g��l��湷1��=A�b� �t�:����l�jj��B/?��A>ڱ�	���[��-B�^2�'Ύ�O�k�;�=��_��(����`U���ۼmˁ,��d����6�>j(��M	#����1��܂�Mc�~�������d��]��6��J��P�`[������VH��X3/L��P���N_!�G�x�D&�!;t`�l����jd2x�
���i�n���M	�x6n"b�ͮ�#��(){ub����%]���^q6��,��H�qgڧ�b�$1�Rƃ��j8����G�m]ud��Pː��`��r"�{�"S���M:2] ��"/�</oh�.�J]7\�ܸ�0~��oOV0`�{a,�ae.D�7�e�� 7A�=<k��.V��e��Z#i�~�Dr�~�}Q��[G����I4��_#yݱV�����Cibǐ�����*Ҟ��B�\I��H�����R�����g�G�'pH�=��@�_��Ś� �XF���<��ҊQz����RA��3N�^�-bb����v�M���|��G� t��R&Y�>EvdqV��<�͗1n���_��S񑔏06��y7��:	솬I�Q�ʄ>(A��:����g��y>]��b>K����s�_S(4T�����w!��71``A{<P@�Si��ؖKx���Gd�R�-0��n�=`?�(�.X3�Z�dQ�j�D�����W-��y�U���7�����|��O ���U�5��rk�)�75��4�[�)�Yep��vQ�ᄦp�ԍ��s�����_���nP@��@���s�&�1����2�A*�љH��0dn|�S�ƀ:g��P��X�$iT|���}�@U�"Y<��J3�5�r�����>a����Z�ρ�Ş1"��;�����\�Z�L�g�mf���o0�� �"X̇_�G4��Ә=�|�T��Q�o���t~����� '��IB�
nC�|H(�![���6��W|�{z�7�&�Iye�E�SHr�'1#�0,$2��֏�;�����
$��0���Ȼ;#��ި���uT�4I~���m�>��0���Uw��½��!�hx���[k�Z���/0¸�.�,)��,#���X�y�#���(8��a;�t��-,j��׆_��d��)\��hG`��o��rHڧ�o�ΉoE�v��U�%B>]���.U��X��bY@��ti����r>	�#~��P��-o�f[��f�9��s�m�"�hݿ�E�!�oe�W7��*���C� *��b�1��TDӯO�eü�*3�|7��6��r?C4����^W@k�������L݆�mi��?�#-D��ɑ����X#�dڒ8 L�2��_��̈́����ۦ"w0Z�G�:j^:���ۭj�,��m������ ��$6�����S ?`���Q�Nܵx0�iE�Ohj���*���� ���%��̒�z+�X�Z�<�;�/�� �=�`�+������JN(l Z
KL�X	�l�ZU��v����uߧI�ꬁo@��8���TBM���?DY�}�FOa%�_��y>oB
�����[TS����a��[�>#\�v�j�-�l� �(r?s-h��	�΀[���O���k�l"�U5���v��\h��#�,���Y�c���J����5���w5:�
G�9��;��R��%!�'�(�a%s����h=�z�SP����a�\�HLm���w˔��Y�L?��@OV���v��-ך7���}.�@*�0�8:���ðuī� v=;j[����6$��m*�]�Pq�[k�aRH��D����Js�����&W��xg�H�Nb�������*�D��2E���bB��o�@�n�2�w��i�x��*��Ə�כ<g��۴��w����w��|^oZɉ�n)��Q��@��m��)!D����J���d?c�Q�ci�q=�# �j&+�o,"�Zހ��ß~s��x��kN8�ٞ<+���f}�lW<�ں�]�F)k�8kG�]Ց�����)�"ǒ���s��Y���|�J�q�k�/[ߨ7�`�����5��AH��v�C�&���'1;�^ߵ�Z�t6�1m+�pymK��B�z������e,~s�]I�?F�
���T�)��c�?D�
��%��ٯ�m�F4�L+���X!�Lw�[�<��A��ݓ4��1��h����gm�0��F;�z����g�2f�i5�¸�c�mV:12'�P?iM3>��G�B�E�����_�v�=�i�lT�=�uVlG�"L��l��r��9�L!���▟�T�	T�����Fŷ̔��D$�!�#�f��J��pr3������^�]�W�?�P�*���H��Z���5�7X��E�p���Mt��d�s� ��Z��!-><�__����b= Cb<0��?c�A�ç�c��K����!�0T�b��:�b[�t��l�ؼ)Y��C۲�غ9��ri��]@j����o�J��ּÑ�a>'FNf5�-��m���w\�X�b�Θ�([�?hcv@d%)L����P��(��G���p�zE,3�c���e���B�tLu�=E�~�D�p�S�.g�aO���v�>�2�=�^̏%���y�M�Θ�G��>��/>3��'a{���$�QE�|�>X(i�YW�
e��,���	$k/X��yV�������~�"S��տ�	�6ۙ�Ý�XB�C����[n1~c�+ِI�į����R
'y��˸ZRP���ܤ�U�{���Ҧ��H��f^j�Q��UZY2J�Zs����6zj�q�w�ЭvD��Rl ���2��C�D������� ȭ������.m��Z9;9Y����6�����1�/�Q���H��=�4G�G�Y�����k�+�Ū�K�3��4#��a��ˡ���6>b|�@:/��ds3W9�c�\�6��Dm��Q��NU �@�Ze#B���U1����{{#M��h��0ہߦg���0f�?thYY�%����զ���GK�����߄��IL�t��9n6Px����E>���	+K�K騆9�e�0�N9q��E�;�����щ�9���H��jNEA�3��S`�˒�b���zI�ԛ뤂 b��������5u��ĶGQe�W�:�Oy�:�Ɇ����AOf�C�8uٓv:lAG�5F�aMO����� ��� g��/�M���N\�| }�rO^<RT+%�������)C{��@\ɮ0F��2O�oX�����~�)���nB5����z�U�<65�Z䶘%���5��a�� 3�Y�Y�]A�-���ƁU=ǀN��K��٠��5�Т�G�	�jd��K��vX��U�z�eu����=����8,�8j�d��\[�|R�7l��F���ٷWp@�Q�F	��H��^��]R�p��h��i��Vm�5~_.�u�f��OF�Dmdc;<���5k��l��\G��o0��'O�ړx�^����k޴��Ž�A|f��Eq.҆|Y x& W��a/
h��iψ����w��DyE�V�
�pm,Gv��t�ʠ�N#�G��7E'��G60��Ӭ,6oM޲���u$�qH����1��Y?�/�2,@e��Hj ���������W��Y�]�>�\���OJ�-��>������F�k�uT�LL��E�H�74�������X��%�2�����G�pF��?uS8rq��˛:�Q�E�]�.Gr:K%�ؔ~�ɥ�e+5���:3m���L�Ȧ뼲���0��*�Ї�����S��Ca��"*G�����9}q�&�ǒ�a�/iOG}�aJ������3*=��ֶ6;��<�c�2��ӓ� j�A~HO���;�����9���zL�]CA�Vq�5H�$ma6��J�9�|�n8ă%�S�~��Թ[����H2�ƄQp�z���Bf񥴂D*S?���d���@[�����d��A_�����oɘ>��-
�>W{�!�ގ�FxmI��V�@��߳�尿��j��E�cӫ�f����VF]�;c�h�냇J?w��N5Q��磒�(�v��" �OHz}�x����а$սP3BԎc��=K
R��u�}L�B�o�O#�*N��W�/؅�
Z�o�/��I	�1W�d�c��5�W�N�\K������EP1�%/�n;df �	6���R������M���� 1iv������_#������K�ɴ�����1z��D6�	չs�~&~��C;]��i(�f�R&&��_6=����-T	I�r���S6���^�Y���߶��Q���Y@���r��;�F)��}xR#�\�S����)�ġ�6��P^�?�c�Z������q��^dy�=Vzv&Y��`��������nkX���F4s�F�t�s&�i�e��8b��W�}�5Z!��es�-Q��Go��`�pO`M�c@�(8U�S�'�ƛ�:�q?n-�h\��fF�MW��D2�"�̙y'����҇��@�f?_~>�pԋfY�4s��U���'`,h/�y�B{�^pYq�]�sM4s�ٮ0v��l��Ŏ��W�H�X���F���G GR�ݜ��܋3� �s5�۠?�!������É�>H�6�{`��-TD�(�D��W�������cs��z0��٥B���#i)��z�~���xІ`fU��X�!��B\����ΝT8���M���8F#�i����n���ht �Vwi�V8*��K�|<�A)	.�q�#������W���i�+ ���;�ބ��CǬ=D�����k��uG�\�'��qPT;����C�ѻ�n.��T�TQĂ�t�^}h�PB� u�47����A|\ת?����"f�h� ����d���=�Xx�r��@�຿�==}[[���%%����C6�D�I@절�H4�ۄ��8}d�ǩ�d��8(�u�!^��i Ѻ��y��v�}"�嫫���a�^7��C&}�pJHd��%c��Ye�g�)��0bО�?��7��\[��#f��V�J�����ʍSI��΅�Z�J�XWh�V�ɒ_?+����h9wH�^$�Q�}\�lq����_���d[��#m�����99��B��l�/,��	0�ݯ���('�{M9 g(~
�-�K��ݖ'ʘ����c��F>��w-l�ذg 3�3�y��˻8�0�He�� $��q�a.�v� �E�|��y�z�=u[�U%�}��M�c�_������ǰޓH�zN�E� �����x+w�Pi�Mơ�%��H�w�nX�ε��Eb��Ԃ�,y�&�fK)�E'^."1��J�'��rI�l&pse;�y;{��q|EL�.Li�*�@��_#�ʍ)��2{ܚ� oS�ͪ玌j��U��� ��p�­��v�ry��:�ɏg���aU�h�'�-�&�^/�C����)�jGic����q��&<���]��/�JT4�ց:�\��o	D':ʧl�<�x������k��X��-/�bD	�G�N?�ۄ�,Z�s<�
���ʖ�QM{���"d��ݼt��~��:�]�h�R5&^o�R�н���fb��_&�aO���a��5r�J-�z+�!߽����+���Ь�ָ����)9�qJuqϯ!��\��;���*�_	S�6���(Pz�>���m (��q�z�26!�amsI�v�6p�KH��w1_��hqp�����wC4��*K��\LB���l�G����/~�XIe��Vk�KOM��;T��i\��%RT�fy;�X�!^}��긲7I<ޣ� ������%E?������H��
:�����'3(�0ZJR�����cg���f#-S���Ѷ��Q�)�����h���Wy|��c�����}	�_ft�&����u��4���g�*�*�D���f5�K(5x� 8����0�@a+de��`=8���ms��s���'�S��+���"��i�ZR%{���UD����ƍ�RWeN_�6�^��}g��腒\Z���,��;˹"t.�9��+wg��l[Y��$���!� A����mt QTl����7g��ot�/L_�A�c�V����K�D����[]��R4�x���$_����(����o@�����m8R,�m��lI�6�ӷ(���M�?���X=�D^����c���/�s�1m���9Y��F��wE�PTQF���;�ꮲ����3|��=qL�����t(m��
!�<#`� ����j��e��I���bn"�Mօ�6�fD�$�٩��8��P{b-��E�R΄�Ʀ6O�95H�rg'.(�O1$�����7��s>��T�]"2�P�m�}�S�2��"��܁�~�����ZC�]�%�"|< /\��.H"7��:����y Oc�'�(�웮��D�^�eH�&7ns$<8>���+��rst���eD_�z�J����C��3��&z�p8���3�n�6�/R��X��� gqKY��Ѕj����\u�?%\>f�f�XI�}w܊��I�������ã�%O�Y�6Z��o���ԉ���k�q���Pwa��Vc�R���-���i�_2Q�t8�kܼ��.��jR�g���_}SF�f�6�ǭs��`�~̈́����*������2	�f���K�׵x��6��c����a�[س�Q8������=��1�j�ES��3'�3�R����UP�;1�sa�خR�6�_'1�^y*�g��&���才�#7,������t��V���0g�Mpl�ir��ą��.�A�2Q�t��&�����@�!���w�/�:A�������D���4�I�f΅@j�B��������(5��94��2	��'m�)�,v6��v+"68�o(XU�M`]ݺ�/O�������c��9N�{:	�N��ƍ�Bρ�jP��Â��e����h3�R������g��~���[��!2��`��쩣�`j��~܁V����In,"@M <�6e�ח�ݩڄ��2}�{�I)��[ȃ\����&�6�wbЩH���gq�^��7	1�8��v��.���Ԕ��],�G���A������"�@Y�93�����$24]���"��/���.V�7�>6��mꌠ�O-��24��U-DG;�e~7x�i<�F��%=�<�����D�\��Wk�`��.6��@";�6ǧ0%�V5(I�;U4b�4�%����P��엃3ݍ����[�z������~h�p_�Y=��Z�6q%�Q��m���&
R	����S����'R8��3%#���䊀8}��n�!��hH ��]R0B���d(wX�0ݬ6jY�����B���񈥂0+My��:�m��� Q�>_�S��G��gy�Nt����K���ʙ�S_�-T,���>���u��V�7� '`�=��Q�S��bح���
�d�7�-�U�n�o�`��C��з�xQ6��;����~-b�y�r��d�c�j�W���`����n�I̍Mk��f��5;.��l�aLY\���M���;{���?����H�� p%��HInG�H�(a�*��&�D޳*�l2�U��9���ns�S�9/�ʜܟ�
��π}i��5�1d @lG%P[�̷������a1ȵ���q��Z�	��r�"��v�
�OM�ZET�gLff?A�og���7�T"Ow�6��4c���/�+|e���{o�t�����^ ���I���
�W|�0v!��4R�������r�7��IоR������ǚs�8#"z#$I�ֆ�)�d�a�Wa�{�0W ��+#3<˨�+uK9U4 7r�aA�>��0%��U�3/����!�&̊�+'k�������O}�ϣM�΃�&�8��X6�يo?�n�%��á;"P��'$)+׽Ļ�{�,)S�h�A�&�Qr�����߉���v���U�X_>� ���;��D���>���8Up(r��\���NA>
��#U�cPUu�oe�f�N�9�%�97ݶD̜���eG����٘�@���O*N,�y�����ӆY�ez�*ʍ�7km68�a?z�u���=�Ut&W\�^_����LT\<m�C�?�2D�삑v��Ю0��l�)b�L~��JK���Y�7Q1w�kԺ^Ѿ�X��j�~y��%�w�������ϸ�G��� �ʆ�X~h���xG.E�`A��͜R�w T݂%��֒�y�o=$Z��;���ͷ����%��\+x�+�S(���Z'w�/dTl��W���sƳ���4������O��	i�8�^ށ�Z�B�����AY?�rF�a�%�fu�c�o3�`��s�SH�ҸHY[�X\��qa���|  �3�?
|h�#8	�D[׬�Ťܭ�c7l���5bY�v��yh�ፃj�P��Y�ߔ�� �Wy�5e
��EJ���*TM�������'�'�g���s����D=I�����ρ�a⎠���N"֪ɢ�a'����w�Q���v����q�\�ŏ!.��K����:&���7��!v4Vm[�y�������Q�qQ�Ø��H�:��8�!ŝ��K�m��B�����b�}F���*�m�hzz��>�b�k�oa	n���w�r���+�*�����<��K;���e�5�'wD|u#�ɀ�' ��Q<c��'ӄ�c)xm��Bb�ar ���?:ݩQ����(#ws����+1��,9�8�w6{�vb����o��8������+������}ĸ
<���=��F�G�8ⶏ],�~�#)�r����`s�F����ZH����i���ߧ�`� :������O��*CnQ��q�M��
��9���1d�LpP�S����z�ͧ�;�̑��d~���]`g�F�y��r������ir��υ
��?�Y+F+��+���X���wI������A
��k�y�D��_���
mR�9����4��(02�[7�����?���~�mю2�Oa?�mQ>N��GQ�j�\��8_��y��� � TQ��u^�WGF�L5����C��9!g�@�-[cT8��p�9��i2��{���{��!��f]_�eq=r�ra��e�u�+�N/ȓ'v��ua[ߓd=K���#��||���MkC{;�Y��R`�
sq��-�C��!��C�b
�C9�V�z�Z��좧G�Ʀ�K�2�10k	wbꭃ�9��t�������*ݚۙ�� ��{�@A ��>�Jp�:�Aa��wN��/-�O��k6w3:�����/L�[��%ږ�Zc���d<�+���'�](�,�GN�[pR��h(c��`��Lw��'t#~~=�h$~W߹p`A!�q�A ?Aaf���m���	�=XI�cя$Pg|��/��|��5��/�$ܓ�l{u�}$`EGI^�o��i�8���"��Q���r�Y$ⱺ�)K	��������~��߻z��PI�6r�u��B|,˶$��r�~��c���� і�x���ɚ�y�PQ���P��{���{R��2�T�i+�ؿ���d�j�"��lR�2A�NJ�/���Xj]�jwfo�v�0�Ejd ��2�g�PD���W�̌�E5�cT��W܄E�_�QB�`Yo�<=�ٌ�.;1.k�P�������4��G�V�YV�ߞ$��+7$��� 30�4���X��x����m��@���|13Q���zR�-ȦDD���N쎊@��ez���"(Y1� ���CJ{��c�(���5�0��?v�v6h6b�� t����n��K�?�.[r���S��X9ei xrj�����w��Z�����Q��e�qN0�x�n��˨�G}��.�\�B�es�/e�N<� 3�&)`K&��n�I �s�"� yD����|}uM���ީ���\�ͦS>:��Ιɞ"8�L���u�|,:�k�GEFT�~O4)�X��g��?���l��\>�}}�EO��TB?���M��b�)����!�0\x�m�U��,�͆�K����`;)���n�)*�b�5z(�\sw���c�����������p��`���dl��UU49�%4E���A~�5C萢t �lj[v�K��s�-���h�ܑD�ءL�)�8Cşj����3�8|	G���Ľ���X뭷�͖�h�h	܏JH�_�g~4R<����&�i�_*V��<5��Bwj=ϲ�.8��K6c����dx�k<��l�o�Sܕ��I0VaHO�`�x���ԇk���&c��%�|=��E(����rx���O�
�@gi�(���k@��FVE;�J
�W��rͣJ�Cu��&�>K7���9�AN[,�<�M5/���$��&q?Ͻ�����D$u��	",���џM^��'��(���X����>N%��q�Jxc�u���ņ��kZ˘�����{w�mNo�6��XW%�_���3B���^�U�A�,��kSr���U�:�Zk��r�=[I�~1I������=:*��t!�Ldv��S�(ڵ��'���C����8��a��"�Rs��!	9Ծ%&������}�O��a�b�0V�3�BG�-k�;�(<�7P�)���j�� !��3�_����B��Ā Y/i,{��ߦ{���$w�E>� ��&MiEd��X���粩��$��5� M趕����0~@�"�2����6�/B�+KNB
��ˍL�);�~|�cd��W��k^��y�`K����P��9i$9��ӥ�j�p�֣���{kj���#:2؍P��j����j��=w}*�v�N�G� ��*2�𦗑^}D W��P��'(�Zy5������WPi)�Y�|�trd�81%��'�V�p����O�G+�`Y�⠞[��++g.�� q3fk4Ѓ���t��o��D��J�?@�@Ჶ�3(g�1�?���D���_	N#&5@�aeq�����1�[���v{q�]�H���C�4Ճ�6Pt�M}�h�l��x(�)�/�ŗ�K�d��E'?�l,����B��9�hx�\��S ��������`���w�(�:e�7N�Qa����"Q<~Ҿ��H_S0���`Z��ۮN�ϵ3@'h`�53T����I��eE 0���� ��u�Y��밨���͝�*:��H�����9`��ou�Y�:��8G\�FKFO���л��ONkg2u��AB��Q \U��}��Ol��T�х�7���B)Q�x�X��\��T~����=�2�Bl�)	'n� �y��zS?J��m��&ȫ� *�o����r�������;�<��=�U�����Y�x��m�5:}���J��zj���K"��݄2��#����
b��=� 8�:jZ�Ϫ�P|`�)�u���V��O���e��f	sc�H:�Q���\Rsh����i�	V{j�5L��~�����]���S�c��M�[)k{:lc:���1�0�DO��Dx��Ќ�k���|�7�v��|��E���Jx��%�F��
v�]i���҅�U�"�E�Dz
�3�����iX��;��5���a�7��s�UR��xqY,��]M,���)$�oaq֌U�
�|�����sO,�jiі!���z9�ʨކY��lP��"��>��wˈ�8JS��Lڨ�ɀ̆�kё��Z�o��z'�d0��0X˒?%���<9p��M���C�Ter���W:�x��榭0�r��r�~(9.�s���oD:�����4�L������#�f�x}B������uj٩SK��a�l�"�fߔ��9˼�&�|�����`�O���aX)�g��3�ϲ$p%;���<�V�������6( x9��<H��/�h78;��j��l��$JL5|)jV?��HCH�m�������9z����rf�s/=��ڢ���Y����K����pU���+H��E����Sop��vT5����o��2�3A�Ws��)Tɦ���b��̄�o{:��Pm��V@���-����FO��0�W!� a�][��[�V�O�;b��h����p�d�`Q�A����7(��.��Ѵ��}�tU�ac��F��zEB�ạ��
�j      Ĵ���	��Z�JvIJ(�Ȱs��G}"�ײK*<ac�ʄ��	Z+t�\x�kg�t�D��B-4�+0&��|��(��
�w8Hm��M�Զis(��7�IE�i�e03"WU����L�%LxE�� ]��O�3��м�M��	Q)�t�S��,(��| N@���DB�`���yݴ|���<yU*}".��j����
�Yd.����q�F�q������#����O�#��1�(D!X�K��� h{�#<��0}|^�I�_W���_�<�6�H�K&!h&�O�̰���
��_jb]yRн,U�6��r72��XU�"<AK5�'���S���DSB^i�d�	mk��RR���
Ѽ��qӧ��np��$:}R@�n�'#
��=��
T0-����B�z�`ꦡp��	4��t�v-ڵY �͂��4m�����M��R��c����I)��	t2��Ӄo*qyVqɷ㕱N�`�F�:"<9��*��Ob|��ń8U9���W�N8$����I�ra�k��'Sz� �߸.k��:�*� XP��yR%I�'���&�`3$�ʥLJR��s���\2uH����Qb�	3�Q�p��.�y�+��F�P 1R�-�O��'�t�(�j��H�L����(4���&װ>;2�3j]	J��tEቡN\�A� �
�R% �S���Kx ��'��hExZ��FxB���5�8, ǪٰPm��9�^�y��T  d  � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                P   ,	  �  J  �  
$  �+  <2  }8  �>  E  ]K  �Q  �W  ;^  ~d  �j  q  Fw  �}   `� u�	����Zv)C�'ll\�0"Ez+⟈m �6�I�J���D<c����N�3TJU�� �LO>49�jޅ��еB�%���1���q{&1��<1x� ��=�b��xQ��ȅb�R�F���Ipҙ��"�f�)pUiQ�N�xs��'+h���F}BF#��(�dI4K�Q��pLꐆQ`�jV��-����Iq������~t�ڴ$��;��?���?��Y(ԛ���9%���0 4!��u��?��iWz�{AP�������Q����X�I�Gپ}���1 �(T�A�Y�/����\�	՟4��Hy�⟋�M3�'"�_�4�bXSթV�T���oC Z�r0Oh�i��	/�N��W�M6:�6$*5]�h͓�(O�ԫ���}i�I�Y�I�7)�a�,"�����O���OT���O��D�O��'�y�쑱)ydQ�q� �n�D̓r#H7�?�&�'M����OZ6��O��m:�M�V�i]��'K�I�$?�<Y��EύrJ�8p��	*���@X�HQ�o�}nՊ
�B�k��
e	f��v�1�"��`mt��XmZ��M�������4��-K�LE�{�X�&m	�w���J�Õ��?��B�5aQh��Sî ,����3��]��W����od�Uoګ;|�s�c@�h檼B�͝�. �X�L0Y,�ka�ʡ�M�i7-Ź��G�.�uwge�uK[w��-Q�i�:!h,-�' �@�����ݵ�N޹OK�l*�Má�i�bXR'C� %�L��D5�0�["a��-&���_�_���a�Ö+y6MV�bV��F�@�0p�����h�����'�Ѝ��P�Bچ�i�h����\���' �O�(�d�&����	�tU˲m�c�ԡ�G��]!�D�F�.@�c����������<�!���B|�i\�Sm�@#���G�!�C0bż���	�]��%�6ć�"a!����3[d�S�P�:�⣣ی^!��W���"��+F���Z�ўH"h8�z�:��!��%���p�I���`��+�}r��A3[wP���A_�~A��F��	���'�t�2#H�b�ꍆȓ1�F<��k��M�JQ/��<1��_J�<�5̫2���O�t�H����L�<A��C����z�8c��)S�a���V�V#<E�T K[�ĳa�ۥ~��8{���!�� &�������.{��%y�eN8F�!���;w�0I�@�Ń}���v%[<&m!��6n���C$/ҿ"jF$@ʅ\!�2Co�e�a�Н]콛�'�%[!��1#�xQc�`�xH�h!Cg�$]E�	<.���)B��[G���[�8b�ۖ&!���1:Z$r�n[24�,�u�/ck!��U,}Ub�
tFޙ'�v��$~h!�dKd�40vmJm�9��̀�3�!��>L��5���}Zx]p�c��y����y������hI�g. ;Q��
t�r���<O$�S��cR�8R��[9�����"�zL�p�-�Qt��2��T.����R�(O��ӪƎxn�i�1#L DmX�1�&+4e�];b�/\�1v Άb�x Crb֮�(Ob隱�'X6��ܦ=��7�z��FC-P�z�Q9-�.��	�D�����IF�m��
���N����$��9I��l��	��?�3kȓ,ph�*7�Z4Ic�����ǟ(�<��4p����}��ǼSd͐�I�fx(��Ӫ~J�Cc��}�<��ҴR�6���f�>g���ۡn�@�<�$%�n�*�Q9nq����<��"����h;��S4N��CS|�<1���9���X�N�wo|�
q.�\�<iR͂	3f�����{,���ڟd˔)%�S�O&������̀h`hՎH���E"ORd��G�8��pM~6�r"O�M2�b�>C��d�K�V�����"O�Հ�AȚ8��<�5�ɾ{�MIA"Od��DY�Jq�}ӆh4�̊�OR��'�ЅJ�X��F J#A��r��C���4�O����^�V��0�)|O�pXG�K�L�!�dZh�tM:n�-����5VR���Oz]:S�ʡ $�5�t�Z|՚���(��O>e��P�8ثd��!N�dh�"OZ�z!kV�I��,���8� b��|Ly��=i��t?q�$��E��Z7C�?���F�N�<� ʤ �jظ8��	���("�81�"O�T��'^��䋐�^Ф�H�"O
�"��ʊd� N��j�"Od� g��t���և�=��0�"OE��f�ͮh�`Ȝh��$k퉳;nʢ~B�.O&5� ���/N21x(�êF�<�0!O�P�<x1֌^40���bBS~�<��h�z�8&M^�Lc$����Y{�<���6]�.�K�b�,���
5t�<��@��q�|�DFP��8�fHK�<�r�E:-q�{TH1"]��)�J�X(��'�S�O�$e !� AU��'���9^�-ړ"OL��N[�Tf��(�@/N����"O���R@�%I��+��¶`K�l�V"O���ӯ�]g�d� /��]��ã"O������(>�{`��\�8�@ "O���@˚+hF6(7ߴv��DzS��"�O#�OH�sF؛vTpR3�!s��"OZ�kD�IM� �1��ϛ<Y�	x#"O��F䞲w��G��>!L�I�t"OJ|�1�X�(��ْ�ܳ7.�Ux�"O ��1��8��᠅	m�;�'����'�d���プW1�`�R�U�N2�'Vdh
g��hz�t��3��qx�'L�i+@$��ĺ$l�8yd�Q�'�
y2�&Es�����խ��1b�'��d��n��,,K-�2&��Y�'��Mb6�S�TZB�S�B������	lQ?}�я�]R�E 3.��#�$x�C7D�@b0���i��bdA�5�5�3D�ၥF�j%R��G8t�����1D�d���A�\ (ez��%51�=���/D��鵦܍L�$�"ڷx2�;��8D��Qr(߫%ՎE��,s�e���O@���)�|��3�A\�H�zt�����P����'��Z�� 56���4�	v`�'�lM��ES+���DnB*%˲�q�'�r�0��+���(�m �n�!�
�'ߐ ��8��x0�["]H0�
�'�T�uo��R�Bd�bFX �(O杰��'i��1��@��u��X�`��9H�'"LI�d�H?]PԪCm��KX��@�'=�I�'�(xn��r!�F��8��'�i"�d&�Tq±��C�x��'��+����r^ܓa	�46�Q�K���^[����㉵"\(�@�+�Y�ȓ{8�8��#� }���t�?�je�ȓF�X����1bw��K�(ٽQߊ���`�4X7�P\Q�T�"�"I-4D�ȓ�r9�T�@�@�B�m� �Ćȓu+h��6)�uv��r�˾96PD{�������	#g+��Bɴ=Quş��(y#e"O֝bt�ݩf��$�D
?8�����"O$� ����2G���r��T߀y��"O\ N�O�Tј GAgҪ`�b"OH�)�e��hg�̪t�j�A"O,�eJ	7������ j0P���'Y��k���O,������;&
�h�l�g6���ȓ6�h� ��.�j���L�e�d�ȓ{j
��H2 �Z�wG�Y�FI��Gr�Ī�O�>|��eJ�m���j���(L�~14�#Ri�;�6Ѕ�nW� �$LɈ2��{ߺj�'��5��]/`�9�˖ݰ�Q��ϟb)�Ѕ�S�? v���N��2u��nZ�h�"O~��䂬6�T�`��P�:�Qt"O����鄞������$.�Z��"O"x�M�->�$J�jI<J�z����'X�eK�'��mb�'C<VK�ǂ�@@ ��'���!�`ʍ.�isנA]D[�'M� �����t~xm�AkI���M��'`�)�H�.'ͺ]Z�jN7	 ��'���#���fQ�,iE"�� . �'l�����:0�5�·|;ZL��D�$T�Q?!��P:4z��)��U� ���0D�<ˡL*7�~���" e�"�$�-D�!E�D)�D]�eO�I����*-D��񡧑F���V�	�1�,@�=D���$lo٨`ru$�8k%���B�5D���L:������_D� ӕ	�O>Y(��)�'0F��Sd��(��|�3iE$�j�C�''�	σ�"�� كZ1{�'��5@��ƍu� Ƀ�a ��'z��*�;�Y�A��qV�!�
�'a|!M!:Dft�B��f'.���'�tM[㝰m�@=`�âKL�`�-OHL��'�VM-O�
����[�E4��q�'_��p�F7��-Ѡǔ*&X��'��:g�Z�6G� {�CG%dH�'��m�g'U"�T�` F�Jw@��'�n��x[���d/ �@�����?d.��W��.B�|��S�Kf�0���(䒁2ǆˬ@H����F�E��̅ȓ}ъP�Ø���#nSA��=��t��
�ں?$.�����kj�9�ȓ`�Z�I�A�
+�~�@��lֺ�ȓL�(�x2�U�M���p�`���`E{r�L�����2lU8H%#�n�	$�x�'"OXm�"@��?���@�\�:���"OԨ�&�ܓ1�^q3@Lָ"O���C�6-�$��$I�;Cʐ�"O���OY�|�`�أI�	;7Z<�"O��#ҋ��%�i J��UD��ˁ�'B6e����S�x��+�ɿ�n%UO@��ȓ/bPM�HA�B%ˑ6�Ta��)� 1� �F�am�
2HN��68MPV�U�L
A �@ �6Lꘆ�_�5rdi���8hP��$^,d�ȓH/��a���DJ%A�5Őɕ'Ө���`l]t�D�%Q���� �7����ȓ[t�2��t����W! 5#�`��ȓ�lYrשFz���RE�0D,���@c�4i����	��rO�	��h�ȓ`� �*vʐ#A!��� L�Z�����tF��Ɂ@�Rpp�cX����@U��15�C䉒y�`�!�H�A����HIv=�B����%� ��k�e���2UV�B�	-�!�%���N0����`D0Tw�C��OMN`#�����"Đ�� 4��C�IH���Q���x��#Bh�6I��=���W�O�a0�Q�d�2��W�5�a3�'eҜ3w� ']�U�2C�^�����'26Y�E��C��Ȳ���^Ѩ�'���G�� w.� ���C�,az�'V�pФE΃�h-�����(P�3�'#ʐ��oJ���1����Q��a��$X�Gx���V',D�$9��̰;F,�3�ߨ��B�	�4H^8 D�4y��D�&$B�)� j|��͓�u�XQ�.�:�t��"OS��6�BI�wdZ
Dg
@��"O|eI�Y�\w��J�?^��B"O��)��)�V��e��`�8�xu]���d)�O(dɲ+դ.ŀ�'�>y���@"O�,p���Uܸ]�B
YR���"O`С �3S��E���IA��"O�d�������G��
\��J"O��q��J�Kj���d�mP¨���'�<U�'.܅z$'��wCv�bL�GJ�@�'�VUj�@R�N�!%��k���	�'д�!��8�z�y� �`r\B	�'��D���@�~޼(�NYYH	�'�dlcm��|"uq(���]����t����*h6�щe^IG{Ң��̨��1�H�o���06��#���"O�s��xH��@��E�C��`��"Of��&�ߺf�N�:��ï*^H���"O(ؑ�`�C`fmi�%�2Lҵp�"Or���A�J�`�2��<3:lSD"O�|(V���4�������b�'�T�P���S�X�x9qdſ+����ݠw���ȓi��	���>5"PP�OT��ȓ\��H�	W�㜈�$a��aH��ȓ\ڜ��¥�=D�*�ȵ"YaH���ȓpL��U�]g+�9P�C҆��ȓF:�РƢ\8&ٛ��
���'t�c�js Y����3�dPi�Ζ)E���
X�Z�Jܞh���ᢓ�@�p�ȓ F�$�0����!�٨NІ� ׸���I�g�2M�pFTNJ"��ȓ?>���B�B+�*�Iv�݌#�,���	3\1��Ʌ&w:<�`
`{��A.і*`"C�I�

p�@�3DJ�t�T��(`�LB�ɟ,Ԙ��΃!b���F)N5�,B�	3����� n��D��`G�&?B䉰n���3i�"o�Ă���,QG�C�ɂdV�hpt��Y�!2�c��=A�Fj�O�"�p6�"_D0�v�=u,J��'y�)��C�!�(���,[3qgr�	�'T��Pσ09���r ��S���'~D��0�ö@\ G:F��1�'�ޘE�
"���w!=�$���'�l9ʂ%�?s5�@�fCږp3���S�lDx��)�c��\�5��0jJt-�e��hB�Iu_JȀ��2pnl][�EW�AC�ɫZ�,a����"u~R�	š�UxC�I�-@�_�V%��덈�B䉇]W���5H�: �,ى,9��B䉊l��L�!�]�8V�����B��	����ɍ~Q�@£�JK`��̶�C�	+���+���4v$��6��֖C�	i���J2lɣI
�I����s��C��|d��f#/j\��5��Q��C�	+k���0rN	Un2u��e��U����J*�$O PX�i#�B6h+�,�Gk �!�>!��Ȥ�10�|0���2�!��:9`�!ʵ�G5[���a��
T�!�$T�{�]�`��B��E�F-�?�!� ��$i5B�����
6I�!򤜈em��#q)WEd\��\��ў��Ѝ&�|C����	%�,�il�:����ȓ&��E�VAS+l=jP��o	�,$�U��;��0H���B�O�{�전�S�? �H�Ӡ�IV�������>�!U"Ov�w�؀R��T�(:�@�	�"O�I�%2��r�n�ń,�G�'� �ٌ��S�yw��i�f_&s���k��',Q����{@����_��$k��Ej�<��͇@�jUr���c�.Ci�<9�j��P�P=�@-�fDr�A��`�<a�&Em��i�@�\4s�Pyԯ�^�<y��3R>���7�daR� ]y%���p>� `K?�z���d�"��4�_�<9/�@�ZDY���:(H6A�`�X�<Q���9B�qHU�3��h��j�<�B�ť,3�0	$�98Ҵ��$Pb�<	
W�#�`��mL�h�J	Jx���#����!��_�$d ��Şs5ԅj�,%D�pS@��z�Z���E�`�dEѦ
$D�2�Wk�6����
_��}`��"D�HA�FˇX�6RֈF�l�D&D�l9r Ƈ ���A�M�{�t�9D�� ��%/��(PK	z@��$7�#¶�G�TIńu��ˢ�Ѹ��� �yR �"�����ҫh��M��_��yRnB&
10�"���f;�TbV�
��y��ʺF-��:�	�&a�D0[ц1�yR�]lE�d� ����D��y�Te�r90�M^�-d��K�ꊫ�?�A�H|����������eC��"6xz�2D�4ʰ.�&ps����R!t�C�-D���"�Gʴ<��ȊcE0D�|q�AUw�T$
���:A�`��3D���̖&C|��g �t$�|y�14�ܺG΄�;p^pa7I}Ůq$��_���I9k�xi���m84�Z 7$Q�t����`����I���3H��`k��� K��q����|J�cґ
ir�c&�[j�HP�c�[�'���C��@�L��XS�Y}�S�{�Ё���_3Py��f	�7N�t#>1EY��8�	q�'�~<��4_��âGQ5�$T�'���'��y�L
����&�܊9D5�F��	�Mu�Ӌ�qN�E�"+�)�(㟼�RM�p�����b�B�%#Vl���!S����ȓ�yKA����Y�@%Y��Ԇȓo4H�E�C��1�L#��m��|�Լ3#��ILFh����TZ܅ȓ�.4(��_�8E�`o\�>P����,�N����k���eޘv��x:;?ٗ#۵0���Ov�'��IؼKF�T)�<B�Iۙ2YX�� 'XT�-���}�P!HP�>P���O����kH�x��q�Z/L�IC$"A$.�H����MW4#�v�?#<�J^�tPj)�&	N�� JD�J~2-�?����?ُ�1�r��c�X)>j8X�/�\{�	u"O��T�A�N����L�K�֠���'Z�"=�'�?A�yҩV;�>���G1mЎ��Ə��?I�Ld���s3��8~\Tz %:��,��x�<��L�]:�(z5g3�$��)N�<�'�g�<e�@�/b���
�K�H�<�V���[v�P�[az����^q*B�I�)��l���>v���ާQ������70~�>�JHH�б�dK3w0]� �Rx�<1S,�<d	6	��ƈ._�H�y���\�<Y5'�2�@ �f���:�2tkC�<��B&(�s�G�).���7�@�<�KL L�;�k ��P���|�<� k��FVQ9��B�R`(XiAϐC��T��ExJ?�B���n�́�� �94IC!�3D�$�U#ږn����F`�
f���s��1D��� �.�$��tE�]͆u9�m0D�� �M  �L=j���BꃽS�=#�"O$�)�L�e��'�_lq)�"OL�����Xވ-p�-E-XO�}Y!"��O��}�!�2�(R��Y�\��fR8]���ȓW�Q��@4�D�� ��y�Ն�x����%b� �Rt��7�܆ȓ+E��C!�M�|��8Rw#�8&����C�B�dO.{b*�(�6{��)�ȓW�*���k��0��l��&�4	ɞE�	��?�O�}3Q	�d�r��u��+*��J�"O��`Ao�U=����̑
`<C"O����.K.i��Ȣ�Z+"��f"O�dag�{�����K*q� "OXY"ԉȫz-�£�J�s"R)'��=V���	X�'2ꒈB�Ï�Fh.T��
�b<v�E|rC�	h2�0��A�:�,�YҪK2�'DڽfP�Ek�$x�U���[-|Fy���7XKV���4
բ��N�hH����f�@�l�C��H������'_ Dy"� �?��i2�7-�Ot��*:�&�{�H+[̚��]'^�D�O���<!-��"<���v�h�1@�9Ex�=���Kx�� -O��+@,�F���b�+!48�����4�?��L<)A��(9�l;���+&C#��2hGax���0r��(w"�w}�-8�)
z�V�P�R/!�3��{�n���H�.=����fgX���F*f��S��'���s#�6 �<"蘋M|�шcO8��I1��	,M���'�@��$�h�k����r'��ZM�p��	"��I��~��s� ʡ�G�#2�
�HJ�$Az)�ր���'L��'#�80K�L���D�9w�V�	��z�U<�r�'�f�N�d!�&��kR(��,G�NM����-
������8�p�OHզO0a�>�P�iu��C++��!���V� %�|�(O�@w�>�S�ӪkĚ��!��9d��b1��TN?��iNz�T>�Ip!��&�y�'�_�d��� Ϙ� >��RA9}"៱��ߟ�H���¢��@E��y5nؓf��yQ��'x����r͜<��9O ����Oz�ʵꐇ$�ن�I���,�g�'�%��	3m�j6膘R��x��͕C��B��Ac ��bC<��=Y׋M-8�6M�OZ�Or��Ϙ���4v$��q�ÙV��;s�?��@�'�~b@:pX�� ���m��������y�a��x�hz�n׽DUsq�£�yL�t��L��F;�FC�ʫ�yr>?p��&� }��C��y���">E,�����x������^�yb��_��A0�b�i�>y; ���yb��E�0�Vx����y�$��l!z�0v��(�U@���;�yZ�8��!��Z��G�߻)bFm��&~H}:ެ��qS�Pg߈���'2|]2"�1L�Rh��X��
�'��bᅗ 2RlH��=A��P
�'� 4��)�O�F,�!G�0��5ʊF��D\�](�g�,r���؀L�'uLY��܂(j��+#c��s�T�r�_��z͋c��8&�I��B�!sԥz2/ڧT�j�e��G���z��P�-�-����N|4P��K�Pqp∿RĔ�ADB*�@Y��3�T�򃁢!5�HQ��ĉy���0�%�U�@�t"�:T-�ש��[&!�Kibb�ã�T5���
*v!�$W����(�9@h�"*�/bg!��C��*��1_z�4o\�B<!�D�,7'�p�S�&S(\���">)!�޼=A����/C�y���Q�G"S�!�$�\�3a��65�(��2$�!�d��G<q�gdS"v^0ʴEڜ}�!��;ت-���B�,$��d��!�!������ˢ,R�CR�qJe�GM�!��VK�&�C����'L~�0q�ݡ5<!�Dކ1kj�)��I�4C��
*�!��1UF �H�. rEڲ�__�!�� �H*�/Z���Uy�j�cbj���"O�p�d��(o06�*Q��5V��%"OV�!󆅎~>s'�T��<��"O���%�#B谐*�W�8H��"O�y)���*�)�p'T(s�d�6"Oΐ����P��iåQy��h��"O�(C!T�	�ʼ�\�e��:�"Oex��Qoh�0��#��)i�"O ��W,������'k�̙�$"O���+o����ħ�z�J��T"O t�5,��z�d�d�� ]���3"O�I� '��
��ǃ#[F�mS�"O����F�>pGf�j�E�2�H:"O�����L�( z
T�G?�D�KV"O���_-+><A0���R�ޜZ�"OxYF�	�6���-3�&$�"O���Ba� �&u7�\#�+�"Ol�9�MC�Fq�ܸ$H�^�\Tj@"OF�Fk�3	V�=�Ӧ-��4�s"O��9�,ϒY��rv�N���"Oj�`O1Ch�ӦF�dv>L�a"O��k񏆫,�R@(�%ֳ`K�a�a"O��*e�'|ժix ŝ�D0JU�B"O�U�@MH�![�{Ãɞ#��""O�-���ucT]��#ϓg!�l"V"ON-S���-�-d�C�A�&��s "O�� wИZ�($S��K��b���"O5��������r��=���QG"OĊ�Tk���O���#u"O�lA��	B�\����F���"O���LӌAr�l^��<�Cs"O6����9Q����PiG��l��"O�%[�]1,*�ۓ 9�	P7"O�(k&�ձb`��j��guZ%"O�S���e�@�Y4.R#�0�1�"O��Rr]�H9�*���#b�}��"Oܸ(�k�.]��!D��(��;D"O���f�؄Ri���7�ҫP*�좁"O0�jd(Ь0���H�4�9��"O:D�6�Z�V����`�'b�<�3S"O���AHZ�(�p��v�Y(y� ̰�"O�Q�A ��Z�R��S��%#�\��"O8C6�U4)�0��F��U	�'��x҄$N$gN�)�b˟s���z�'�Rmzجd53�B�}>��q"O��R#�
���#�2kR�@1"O�D����G`T4�vϐ?=���JB"O.��5b�� �߾d6�s�"Ov�jC;89L	X�$��qD�p 1"O�yChM�}��St� S"O���ToԲ~<>��7�
|�L�á"Or�x� AF@x��"�	&Ễ"OP}��9aZ��#�˙x�����"O ����̩1�����q�h�8�"O���%	B�5�����ᒄ���"OZ���$F����I�ج��"ORl{ `׿M!� h�"I���0x"O��#��]'0lF���FB3Y�nM%"O0q1,^fx��;���"}�VI	�"O��� �&s�Bd��'�0qg�! "O�a�ЇM�%G�䃣�?CRI[B"O��i�G�32Z��b(�2 ;�}�U"O�E���v>,Р��SeS>��&"O���虪=��a�G
J:v���"O� <zC�D�U�R��R ձ76�q�"O<-QũU_J�i��N�e����"O�����q�)�D��*�n��"O�}*�A¬n�ց��B_.���U"O:�Z�-O:W���p��C"'�r1"O �n�z-�%��eܴ T"O�����iIb��5o���3�"O^ё�b�ONнqP	v��1S�*Ot�0 C@� �"5���K�<�B�y�'�{��-i��Ȭ D���n!�y��%�F=���W"ed�i�t�L!�y"O�z�0j��Y�b�lPH�`�5�yB��;���ץ�F�t�S	g��B��;v����'Q(tk��t�,r�C��U��1�¯�,��p�'�G�6�C䉇K+�!HqMM�")�h	�&Z>m;6B�I�n�n�qJG o��+CV�?�B��0]�4�����$F��dhA�U�DC�	<����Ȋ2)�h���d�B�	�Dv4i:(K�t^*<R�e �|�B�"c�ȘI⍗)u$�Q�7.�.1C�ɪy���3qfP<2Ƕ"��]6#��B�I0s*D$��W��(�qK�		�B�Iӂ�3�h-+�h8w�ڋ~?�C�I�HjHH�N^>7Ռ��#Ǚ�dNB䉓1`�W���O�H���J˨��C�ɢ`��#p삫��h�`̳6�B�I�',����A�2��-�u�Ⱥj�RC��\��xrH��F���� ��_�"C�	X�]��m'h����Ǥ(B��v������(a�zQ{ c�5^�C�	/Vp|�%�1n��1b����C��$>�V���D�)s&9
b.�~pC�I����"�-���<Z� 5@� C�I�94�YW�04~�*c\�fr�B�	�B�H@��x��⊛�8��B�	�o�@�%6.��da�bD3��C�]I(��0��?Vφ�Ej�V�&B䉯N��s'�K�f��1�3���~�B�ɝKd�h���W� %Ys�I1�PC�IU-���d%��m��I���C�I8/O���s�:T%��q4�y�B䉑s{����.��?�r�STNٮ[�C䉠J���.r�A�K�d,B�I�h!0��!B>hWj�PsR�jC䉗\��0f,N|�zFhǞ[LC�ɐD.͘��=t�8T��B�.Щ����(��ѹ|XB�ɪ|�)ɓm�&[�j�*��
xB�I�-l��KF��-{����*R5FUB䉨K��C5n�?Ξp��fBr��C䉬�J@��m� h��
�_���C�I
3�,+��)�|ӑ��<�PC�	y�vCu��%*7�$)V�)w�rB�I7�ԣ� �)T2�Ɂ"Q�4B�I�^V��k��Y�l�ՓD�1$�C�I�c^iy�	�T�J�b1M��C䉧N�{�!Բ/
�8G��E)B�Ik�h��o!Q�� �cD3ʡ�F>W�͘��$ C�P3.�o�!򤂭od�Ya��DJ����U!�$���!6�+W.��q��G!�@�P�,����B�`+f ��!��H5'Z�i:��H(k��Úy�!�� Ɖ�e�E~X�R��&[�F�9�"O���t �78P� �4l2~��0"O�rעڤ} 5z�aI<Q�p�q"O2�S�NZMq�Gۓ�r!"O��Po��#�,yR�d������6"O��jp�� ���F+x��	#�"O��� ��3[(Jy3�K=v�npxu"O�s�X|��:��@:5��y� "OF�Zt.L�:dmyďB�e�
P�"O�e���j'>:�o�
Sb~t2s"O:4i�I'Qe���rH�x��"O2�g�?$3�Z�#;8*U�""O���¦����(�H�HDVP��"OX� p$ӻ$fЁ���� 0�1�"O�X����)\S�|�eы2IxI�"O�1c�03)� �%�ٛL٠��s"Ox��&�Ci�D�� V����"O�p[p�!�����3��p��"O��R��W���0�`B-Ú|h�"O�8p.�z��Q"P
�2��bt"O@i�Ή�5h����-Y��q�"O���m̢*7�9�ዜ.8#z�A�"OflP�ݖCV]�"bn�\U"O^I���[�r�~�� �] ���Х"O?!���ct ��x�D���`Y�h�!�DG�I�:���cR�p�.���N�,h	!��X`[�Đ��Mui��@��N��!�$�!`��C�+5��e��O��!�DB.����N�n�!,#@!�$��Bw6|�`�݌0�&�0D\�#&!�ڿW~Ƶ���bz1�� g!�O$QQ�eI�L�g]B����5�!���ePٛ��Մ[�$�Ee�f�!�Dşh�9�w���Ta��)t�D�S�!�d��A���fd�p�<�!���C�!��c���� �15�������Q�!��?.O6��(K�H�j��U�]�!��!��1kׄ��g�8tQw/ҢE�!�dB(#�D�xSJ�k�j���m��@�!�	:"J�d���W���9��+N�F�!�d�,@��'�۬RB^(�h�<=!�dR�Ҭ�(�<x>H����1p,!�d��e"�T�2dL)_'f��HۀdC!��VA �����}���f	(M*!�şw�l�8S����p��叴�!�d/ �����)�D ��u�!�D��u�5��=ut"șԊ�	H�!�dZ�]U��z��S6KĪIɧ�+|�!򤜧%�(L��K%j�RЫ����N�!�d�;*�H�+ނ��YҡO
Y�!� tAZ\! �һ'�����S J!�$	$�)�v��a�
��Z�>�!��� ���4���R��#��ÛE�!�$�:i/0�q�I��y҃�*/!򤙰_<T�"�]�`�R8�5�D�gH!�$K��JA�1��g�D�Ba�!�d
Pp@�8s��nܮ����W��qO�u��/I�\��͉K��u�t�|�Db��(�W$,~ `Tö���yR*��[n���l�&Dd��ѹ�y�B_��$�8�D�v�2-kq�G��y�G�8����$���j/r�� ����y�+�%N6n]1�冺X�H��얦�y��L',ZLy�C�
h�L�GG���y��7��cE�Ӈ�0��+�y
� D��d�S�8P�9��3$^�h �"O���̞�O-��$l�"Po��v"O$l� ��4���S�p�v"O�q���p��H��� �>�"y��"O¥���S,%��n=�6���"O:�3"��da �X4ho�����"O�QZ�!W�}�À���s7"O�CNR�V4�E#c�_�>A�0Q�"O���M�,^�����E�&�U"O�P٦�	� }�<��D4$�$yR"ON�a@A�m2(�V�3y�$ q"O�Uh���QNL���ȧfr��"OL5�R̉�H����$��n�^��D"OJ�h�@�S���Xt��hy�|j�"O�$��-�+)�&�qw*�c�V��B"O��D,#���2Q"[��@2"O<$�胾O ���&ϟ~.��b�"O��Um�"���0���<,�l��'��эS9\���"ڵ�� �'��=�Qڒ�R��&�1�$x��'4p@PC#���S6F&%���!�'$l�8t��&f�� X�,�
k9Ա��'�	s�`J7eI�R�C(�t���'�4Ah!�1%��aWc��.���'���)Q�(���;��8b�l��'�FHұ��ɜ(GϬ�.XH�'��R#Jݏ=�PA2V�
O@�C�'q&u�/�5�a6dC��'XH�3�$����l\�	n�9�'��!J�eQ�nT����	?��h��'��I���z� ���5���'�^����V,V����N��(��'p�mp�.X;0�{W�>� ��'Դ�bo�&�h�P7�H;�N\!	�'���{EC4���مG�&=����'#��1B�I�	�B�R1��'�D��C&� �� ��b�c�'��ɖ��l`��
�(� 8�'E��c�'��r=��c�"V��
�'�B�9�!_'�.�Z&�^�N��aX	�'<
(��]>t����r�Д@"PH��'���!��+�RYCa���$m��'tbex�jڝ�y0���.�'[
1�G��i ٢�N�=�2)Z	�'�jmP�¸u`��� �fl��'�,�@@��zv.��J̙Y�:�'��1�g�8bW�P�@,R2M �R�'����a�^�B�"Ql�~n.`�'d�
�.�4��T�H��s.n�@�'��YagO�����j4^��'.�!�tE��-�����Iͫj:�h�'��I���> �*�P#o��b���'���Qd���x���&�?m:��	�'î1r�hߑ)(��BN�A�d ��'�z<����l��v쏩|A�@�	�'"H!k�H��`T�k��x�<[�'c>Ũ��ǈb�Xl���!A��;�'��*VҴk��93s��1_�t��'�t1��1XV2��<����yR��{ǘ��e�PA>� �h߮�y��S3/�����G*[�8�����yrKƂd�X͛!�P���ħї�y��M\m)櫋�D
��;V"���y�`F�O������Mt�x��[��y
� h�1�*N�:d���
-	��9B"O��CӅ_8�(D�#ɔ�&p�"O<�cPI��Bt`!YC�&@�"O<1;��٠�8�`��'4{���"O,9�eY3��!9enOCz���"O��HҎX�J�/ѳ$h� ��"OX����;"���MO(rJH��5"OJ�@FԅyR��ٸGAl�a�"O�`���j��A�"�v�@�E"O���vO�L�@��^(�!�"O�
2kV6V�h����c�� �"O8�ë/bg{���&��;Ѥń�P�8���e� zT|�`��Y�  �ȓ[y.�����N��M*��'=����X�0-j��F
�8!�b����ȓ^��x�B;^ZL�`b���\���ȓ-��Y�Aػ^д@ ,���dх�z�֎��,�,�SD l�B剫 v$Q��͗3�\ۂ�J8z�B�IAJ�R�ʃl֮��V`W�NP�B�əZf�A�R�i��@�2AV�2�C�	�xm �	�	�N3�H���Rs�nB䉣�r�
�B�7Aw��r�Վ7��C��<m�h����ĜL���
vзm�C�ɯ
�JE�GO>�X���(ނv�C䉌��%�P�K�j0��) ���C��=e�q�fOE=[���˶f�^��C�I	phu��ɇ\u�8Q��r)�C䉮g.�X����o	��r#.߬^WrB�I�q�qP�������K�R�vB�ɂ��c��2�n��W�Qn��C�	�S.A��i�\�y�b"��=�pB�I%ӒUC��9�2}`c�߁'Y0B�	�*��*�MۓH"-Ul�k8B�	*dd�g��S	H��b6B��=G`���f�_(���ŏ*��B�Ƀ+T��̈�O)<Ż@���C�	.�����U+h�\�K��5K��C䉓yiZ4#�@����m�	>�B�	,T��U�3f@:$��ɏ7)ېB�C�F��5a-kkHYYD�� zC�I$5A��b�'\�
r�H�ޜ�C�	�c<����̑�$(�v�]dXB�I���u�p�^�aX5� �F�* �C�I�Gxn�̖
QN^Qk��@�p�`B��:Eg���ŧ#���[Т�}�TB�	5M q ��Թ~�I���'llC�ɽ[���G��Y�(���K҃^a2C�	�di�]B�M_���akr�${�C��>C~�$H���#A��q
�C�ɏMkH!��D(B�����'�l�C�I����M[8ʺ�*�A�D�8C�ɓ)�<U䃒3�v���Ab*C�I�j8�EH8Zacs!2e�C�ɶJkĸ1���2a)f���kO�C䉄S�V �v�� Y:�R���<;�nB�	%:wz]�A(%���Q-aPB�	$p�|�2˄�=N�i���'J,B�	6!�X���Qnj%
A��d$���'O��:��R�<� ���b��[�2�'0����S4?M*��BeQ�����'}	T%R;k2�� E���&#��3�'����u,J�9�l�� 7%5F��''x�	�cN$0٤�1��Q�|Bx���� ���臏f����+O�|� "OĘ���>Ga�ex j��C�
�F"O����X �@��v��!΢�І"O�����3jJ��,O�J\�&"O��a6���XT��mǻMu��ْ"O1(C`��+��:�Å8Z�}�`"O��P�G�{�(B��#�p�	a"O,-�&,����"ٍV�m�'"O�܈v틚V�F�f�?O��Xh"O"4�4�̇Y�|��&Z�@��Xv"Opͳ�L&��(#��{���hE"O�ͨ31��]�FdțV�F\!u"O:e�o,i��,�'�٣U��ʲ"O���N

\K蠂�K��.�tB6"O���$EJ�`@�Z�*3X�"O@�1�>g��P$N�ZP({�"O�x
��߮D�
�AZ8@� 7"O���&��x~da�V#��pT"Ot�c�: @�[C̣T{E�T"O\5��H�eG0G.&}d��Q�"O�5(A��4#YX2CN�'2a��"OĠ;B�S�+4��l֚0vY�U"O�ă�� ��u���͉Z�+f"Ox� �Җ��\+��1��1�"O���pl(�|u!"�hxk@"O��r�'�1%�.���'X�\���Z"O�����9$R���¡R�cɰ�""O�<�Ģŧ,2�ɂ�A��0�"O0p�ٔT�dQ�bN�xXD�B�� D���?[Zybo6G� ���� D� k6�U�6��񒀎�}(�j�#D��1w��d+�e[�(Ϳ�J���/D�t	 �9Z�Hb�BM~�,T�#�+D��Z5�����h0�N&e����&)D���EH���rp�Q-P5a���Ԃ3D����杢e�Lq�d�۽5L4%�PA>D�l��B�X���1%i�I0402�1D�t���4>Ap)N�}-4��>D���[+I�e� ���_��:��;D�4�e|���qe'��R��.0�!�ؔ�{r�C-V��e��A"O��Qg��+ʢM���Zw�i{s"O�a�Ɂ���Hu�U8fj���"O`�¥#G	z����R�.,�4�R"O4482���m{u慐�<Qj�"O8È�U�����K�#����"O~�pA�(m����N/�b�Kb"O� �=���ӯ[�Ĕ���"O�y�IѣB�a����P4l�!"O�l��,� ��*�&}�V�}�<93/�"u�Ɣ� /�6qN���* y�<y�V#0`�H�L$d�����x�<��gQ洙��,��Hѳg��v�<�4Rg[��I3c�8�~�ե\G�<y$g�>z���rm� h��4m!�䌅"�8��aRJ[2�$A�	f!��)�a�Ǧ�
��1��N�	!��Ҿ7�8	�.\&#O^8��Ζ;!�\��h�E�$dQ�Q1N\"$!�$��m��x��mҺ1@xJ�.I�!�;)B�����|���� ,E�qO�q��O5��HFT�\�w�|� ��>�� 㦧��6� �c#h]�yB!�2��<�Q��2-����h���y�
	�k]n���"��x��k"Ș �y
� �a9 gY�-V��_��r!"O>�S�U:EG�Q��Ě7�2:�"OD�K6�3V�iypm0/�0�J@"OV��$�����q����""Or���d��>.2,j2���Y� �""O�D�D����5d�*1g�|1�"O�yƯ��k\R���C yUTJ�"O�tX��%w-�D�qC�<OL0�"O���C!_3����"�0;M�M�'"Oj�sa��Q�U3`"H*4�8�"O� I0�@m �I	n���E"O������T��'K�S�>�d"Od�U�4N�ꜳ$&M�E���"O@#�!�)\_�ː��A�`�K�"O�D�����!6�]C#HJ���qR"Oj�@l�y�v��lݣ�"O�Ea3���a0z��Ɖ��*��J�"O4��2J;]jK�Lq�4���"O0�X�U�DJa�U��2�d���"O��:���M������c�Fи�"O�X��B��L��2q*�8!!"ON��葯d���zw�FA�e�A"O<��R�םB0�H�I�"!�u*�"O$�"\Fj�HQ���%��xP"O-(�ĭO�F�zfM�9E}
�ȳ"Oؑ?�` �$�c�M��"O����*5��@��-�lN���"OYisC��Z�!��\�xFn�Z""O�y���)>�^H`�D	5E I*�"O�]��;K�
�?�d���"O`pzfO�����z#�߼ʤm�r"Olx�v+�
{�0tQ��E5>�"R"O��C��͇iB���`_>��e�$"O8�2���!	�H,K�I�}�0�%"O��B��ʈ[����R��|�Z�k�"O�Y�SF�(dbL�Q�&ĭ^� @s�"O�`��G7YD�
V+��2�"O�$��CI�L����� `�"O`�`&kÏV&�\�&�
�Q:$	F"O�8��d �����2�h8"O 0���ؒ��1����@�Ĺۗ"O�Q��>e�-�!B�BD���f"O$r����#�J7�_F����"O�e�Hts)%!�����"O���3�ײ"��!&�͔���"O��i�'N�i��H��]1"O\{GĆ�:�h#���$�)
�"O~|dAH�[ڜҖ��#LxYq"OX��̃?<�)��A�C7PI+�"O�u�C �a.��8�aP�p&�y�"O��)��l�$��4r����,8�!�N�QA
V�~"���w��)'T!�^;@��aS
�
pzG��^>!��7,t%C��ƽZ�n=�'AE3~&!��Z�BZlxi֭T�b�T�AǙ�`>!���/�Yr��ț$���GT�N�!���$M2�s7ݗS�4�l�b�!�䌐b���U��f"݈��T�!�D�&4d�Jr �
���A ��L�!�DN%Qb�K�Ǧ, d�b�L���!�dN�e7̈��Äu�P��weєg�!��B�rLU�W���7��"4�ڸ�!�߰�|�P8T�lۂ$�8C�!�%X�N]�rA݉y�@�:�(نk!�� D��R��Y��T�U�^�29"O*�+@/)����t��9GǬ=��"O�`c�N�sEzL���^B1a�"O��Z�V'u��6/��(�k�"O��D�W�X�d�	r@��Z����"O��Rʵk�lh��##���a�"OD@�GL�?2JT�U�� m��(v"O��C�_�P|�AP���p9�f"O� '���(��]�WdԻLPΡ�"O�uA��O�;d�#1eDC�R<av"O��Ya̎=~�-��DӗM�Nʓ"OZ�0d��g��Ւ�B�t�n��q"OJ�
��&]c�A�|�`2"O^PS�o�4QJ���G�bh���"O�P"#�*d��Q�G�&HJ� �"O^Q��ݦ@����oS�\� "O �Z�� \�b5kE+(`s��c"O�ɣ�FJ\0�����&d�I9S"O4�� ���y��RQ�&�P���"O�8Q��-n ��VcR�p�4��s"O8�S��6!hP��̭6����"O��ҋE�_�j��տ*tج� "O�	�u-��9�B��S�G�_�M��"O2XYP��4�$��� ^>H+�]��"O4�C��7s�<�`b�
e4�J�"O:8؀i��p�L���d�Ô"O�(��� �0"��� �S�4�"Ov& W`q� �./1�� J"O�}���[(^g�T�w,ݻQ�Ա"O�xJF��16��PA1l�!QB��q�"O䵃A��� x��+�-H?����"O�!�6�д@Ux����n�J�#2"O��A� G7΍H��Ɵ<i�%�`"O�T��	Va��.�!1�%D"O4m0���>y�)IE��C0�tن"O$���O�[�6�*S�~�,��"OL���ELX����$hY'oJ� "O�1��]���]�G��6w�i��"O��A�P-y:6TauB?Z^�J�C�ɧ;NT�k��8:xi�a��Dq�B䉏>���|!�Xb蝬Xd�B�p��%k%�V0[��!Vf0^��B�I�"�r��ޟ"_�T��#E&<C䉾?t�#tA�Ay���K!.�6C�I��YH�]�A��m��I�B�I�@H�rA˔�\�ȍj���.]�!�ƞ"����]��ʯ�!�d�	�a�閑Y6j�(�`5�!�dUv�bR�O��ёjM�K�!�䇬Ӟ՘B��-�D��e/�-)!��3C%���D��N�dU��Y3)!���O|yZ@��,&)���1eY�+:�H��"O��8��[7����   �Z�ɓ"O��8���0!ƨ
R �j�$ �"OPF ���8���0"6 ��v"O�$��W1}"4A�ċ[-9�2E"O�8iT��=�D����	?���!"O԰���|B}۷�I.a֭�"O�!!�!�<�PpA�9�Ep$"Olѫ���y�0у�`���`��"O�-������@�.�)m~��8q"O��B��:c��7uad���"O�P�,��W�d�:��H�'`2��"O�l�k��v��er�
��{\8��"O� ����-O�鳃��S�� 
g"O��2�E0��I3&(ם
#�h�#"O�i�Ej�j�@��(SZ��"O�e�EkD�J���"��F>XА"O<!�'	F����W�(|�:ە"O�x�S(P���[��)M��Š�"O�P�ì�[�ةzD��5o��@"OL�2@�I�N����8�^50"O@1B�_- ��Z3$H؞��r"Oֹ)dꞺZv"|2��H�#6x���"Orl�q��B�� c��Ϙj#�H��"O8��@��M(*2@��"O256�ְ>��ԓ��U5O6��E"O�땇�̘��P
2�I`"O�M:��P1lK���LK8�
x�$"O�eH��n�U����T� �r"Oh�K򉊻p(���� ��+�L)�"O� �d��d͡%�� }����"O��QToFJ�P�V�`���X�"O.$(��0m�艒%�"��1�W"O�Q��8W ��C�����A"O�px��;��	�b��	}�"O��- k�`��W-��1�"O��a��F�V�v��5Ԭi�a	�"O�q#���wXJ�L
�"Y��"O��ĮM*q*p�N 1���ڇ"O�t��@�=Wwf��B���X�4�""O�}���<���k7�A����s�"OLtP�cM�j�D��r#uJ���1"OvŪgH�$Y2�	b���*4���"O�E��a�"�r��քn*4��"OB����T �%R!jc�y��"O���q	YŹG(M$I�8�"O� ���"V(EQ!H԰*ז�hp"O�TAŃ�e�R�i��
���"Onm�B�E3R<82���#b4�'"O��U!+@9�P�JE:�Q�"O��!�K�@��i؅z�,� �"O�<8b߿8@u"�(�P��X�"O��)���MH6�P�iW�D+~)�R"OeS�#H�V%�Ej"�F}�-��"O��1a����YZv ��*l�-1�"OE��
^�h�T�
�ή����"ORఴ�5A,��e�I^�Tp�"OH��cρ�*�UG�%�l�`"O��aSnٷRA��p��A�4xiq"O@�z�Уv����ETC��MkE"O�EB!���G���f?P�"U"Ojiq�뎝!F&�*��5_���"Oȱ�V�
�.��3/�<LW\�q�"O� ��th��m�J"Ovp�@.Y�N��dԁH�vlz�)"O.X����_�}�2ӜIdP�z�"O�x��ą ns��`e 0M�p�h"O�pZ�L7F���q�" ���K�"O�yQEE�S=��2C�ވ��Iy�"O�����X (��pe���t*OŐ���lU�q�E��!��B�'��x�/��QX$���M%P����'�b4�Ꮤ�p ��EI�@zm��'�v��b�10�ڜ�,�" ���
�'�jp@&��''��@�4�E4
�%p�'�8��	�bU\)ڳf�50��'"0�(�H�H�x³*�St�9K	��� �YJ�L�8����P�.H�P`�G"Oz,QU��/8WH(h')����"O&�����@ޒ�B�ѻ�(��0"O6���;9l�Q��ĐK��!f"O�\��E��@��k��D�46�"Ot�Su�%���r��v#��
�"O�`"�S�jo��i�C0��"O�a�"��"�j�h��de|HT"O�l+Vό��qSf�V;FLB1"O��0EcH)�x��j�+nBN]��"OT�aS��6j��{�](0��"O5`�jS1*Ҙ&�ߦ)��2"O<�Jt�W�y������hx�"Ox���M7!��K�
!���A�"O�ܰ��X�1���DG-����"Oz2$C�o� 8$��n�N���"O��Aq`� q5��A4.9�0�d"O���b��p��a�a\f�ؐ�"OZ@PmН=^5�� 	�_�d�J�"O�� �A�YT�I�nȔt�k@"O\�qP'��	ؠQTMݮh�h�xr"OX�K�a�U�z��憉<� mF"O�"6gO%8P�SF�V�r�Q8�"OB�XW��2@ ��C�8[��Ѥ"O��Ð%�m�(t�DƖ%���"ObX#��� (�=�'��y���Z"O2�[�+<�ݰ4G���@�"O��:��Mn{9��IJ���"Q"O����F�c����i��}D�`�"O6Y"Bk��,9X�h&6�eR"O&Ց�MJ�T����@�h�%"O�`�sb��qю|�1
��"����*Od���N��,r~���$)k@�x�'q�}�b�4aܩP���/úT��'-X��P9�<|���*!Y4�H�'�0�d�Q�9X�ڷ�W�O�N(��'4���"�"@	��A/07�<��'U���'M;C��ܐRHB!$�̅#�'�ͩ3��7h��*Ń`D���'b�P�MP'-ȸ���T��`�'��;t+� �	v�a �Ǐ�y��ξHO,����[H&]��*��y"J5q$��!(��|��L�����yR�,-����ς�rM`�j�ϟ��y^�3�V��D� dh�@����y�g/V>hs�J֞��� �9�yb����r����ڇ�A7�y��c��ၐJ<�<���Y��y�焄7�r�)���*~���/���y҆U�xjh9Rjţb~�b����y�dȃM杀Ɍ�.�=AW�Z��y���,_R����.Af�Y7Dř�y�����@�2�Y%"[��8��.�y�EͷT�:(��@�U)ga� �y�OV��5a��Բ��aZ�y�JV� �P�q��ny�P���W
�y�'@w�Zg,*8ψ��(:�y�L;_6�󧭋 Dh��f䓮�y�	��v���4�FF}*X�R�݇�y�,�o1֙���ؒg�q�o�6�y���`&д����.N�$�a	˚�y�c_3<�h��cowaihׅpۆB�ɰ:8�f�-][��jEH�Z�pB�	�L�x�`G!N�Ne��b&l|�B�)� r�j�,۳Z��5�r�Τ��ū�"O�\i�D�>��ܛԏ��Pxn��C"OHԹ7�6r:�+��Cx �W"O�xW�۵E*V��U��:(ތ��"Oh��Ԯ�B��$�i�(RF��R"O*�h$�!���M.LmNX�"O2$�w`̵Z��zFH�O�>3W"O<-i�*4N^J��P�%�"9%"Ob��#�d�b	zEO�xlNP�"O�	�ԋC�t7-a���=qc`�"O�ZF��-=d:��.
P_���"OD�����$�8P+�Lmn��#�"OM��Nv.)aN��J;X}[a"Or�i�A\y[qp�R a�,A�*Of��1M��;���V%�1�|U*�'�z)�q�3��aa��	@�J1��'�~��b�0���p���0���+�'N�b V@K��
b��1}��'��!���5
���#B3SC";�'�h��!^)D��PG�&I�����'g`���b��d("5pI��:w��2�'�b|�u��
&Fa�� I�<d��'N�����(ij�%�p L�T�$��''��+Ӄ�.`�޽@sd��N��,�'���A�+��0�gYr���'��%���a���K_�\e�'T�����0�d�� d�2(f!��'���SkS ��5�4k�j���'8���%$m@| ��'y�څc�'���Ƣ��9�bŨa��k云��'d4���OH�4	�lЎu4�!�'D�-��ϔ i�Z�"Uɘm� x�'E6�Q��� b�)�ԁ��g�$A�'�1&��VD���@O:jA����':����Cیz$�Ȇ���W��)�'Q��կ2 9�9a7.�L�<9Q�'N�]A��J�b�(�JP�д���'`���Sϐ�� |t+8vZ�<�	�'�(��)\��\@�<c,���'>s�H.C��93�,.����'��5,G�zO�H��TH�L��'e�	PW� =!j�K��NKed1��'Ծ,�cY:�`ݫ�SN�Y��'�vH
�'�{"VIQ��P�����'͢x��ezX���v#ߡO��\�
�'暕��O@��2���b��C�'� �	PK��l].�a��X�D8�p��'��B�!:�i�t��ewz!��'X��{�(U�|v��)C Z�ܘP
�'����"K��̜Pҡ��T��Q#
�'��4�5JI(�Z*�'�#T���k	�'�R<7j�F�hYpA!G.Q���)	�'\̻�$�\{�h�g�������'d93&-7�X�h&�D,4�L�	�'��1�G�)&�=x�.R�7�s	�'�00G̎�#\,����߼�	�'�ӷ́�08h`0���47AF���'wh�Ц�7@L(Q`�M�[�zR	�'�b��2���9��q��n��%�X�B	�'�T��mHN���A��T�g�N���'X �R��}6�Y���b���I�'<^��fV,��)t����d��':�\��gT}<�4bȾ]�0	�'�^��V�0�8S��9N=
�K��� n��,QY�޸��e,=�0�[5"O�|idY:��}�'e;�2�
�"OD��h�E��u���G�Q�)��"O&�kqNؓ7���m]>R�^�;�"O&�PFg�3:1`�b��B��r�"O2��/��i������/UȤ�B"OꙑZ�dJ%�ً�XT�"O8�P�+��!tB�r��q�>x�"Ob$����	Pu���7���LĐ�A"O P#��=J���*� C�v�@8a"O�a�!DsX�IQ�X!]�xٕ"O֐ !��"t��=�Ai��Xz��P"O����N�*Z�a+t*Qs%��K�"O��J�/�"$ ����3
!,x��"O��G�ԫ'��h1�� v�+v"O��*��.AW�e�1��9^`܅��"O�miV�C.���2�nA<;S�%��"O��9���>�r�I��^!o3�q��"O�l� �0L�B@�$%�,�Ly4"O���cjU�4��5�pn�03�쐑"O2=��L��V�Y�&ҫH��-��"OZ���#C���G��qs� ��"O�)K��I�7��]`���x�Ҩ��"OĹ(����@B�e�e+[/}���"O��Ѯ2%�,i	 @�}��2�"O$I�����\�"�bZ��C"O.M�e�B7x_Ju��!uE�Q�"O����$9~��`�<FD�"O,�X�e��LM3E`��1JG"O��X�gR�@���PO�&:/�X��"O�T�D�(+�8��C/��Xxj�"O��ѓ'߼f�(�ICDr.ai�"O�,kVDD ���>Φ�X�"O��U
E}*hd��օ%�>��e"O��˰��3U�}�Ѣ<2��!��"O��𢌵l`N@Q�'C!�� j�"O��s��yg
���N!���"O:��7�����Pfȃ��*�`c"O�3.M:]*"_��|`"O�TɤM�9N�z]� @��x,h"O����"��y�s�����"O^L2 �2b�$���_�W����"Ou���'.���2C̑�(ʹ�� "O8����-?z ��ôe��@�P"OFp�D� 27T�����8�t]:2"O"��@A'O�4л�'�6*�(�"O���2cQ�4���ELEE�1qC"OV��W��{��
�e2-�q*c"O���$ġ#2`	� $ê7�8z�"Oܝr�^�Q�W�]*]��Lz4"O�����з@[\��F��o�����"O�=��F��T��8�lA�R�T�j�"O����h�1	�nU��F=s"��Q"O��(��_.O�6yKbl�,v���"O"�h4�7�<=:kHdz�"O�y�O D�j�	�G��)�"Of��@f�sU���јR����s"O �PC�j��q�����t�"O�b7H��K���1��_7?����"O�)�e�s���C@E�mIr��"O��'R�jx`�d�1Oj[�"O�ѸD�4WU�B���Aߒi��"OL�@c�S����)ߵ	�<�"�"OK ����y����>,��"O� j)(&5&b@ 1L�#w���[e"O
E&��� �0�w���c�����"O��PR+���)y�J��3�X-"C"O0(�!!N �ڕ{��� r���a"O�|��L�N����I	شY��ڟ|��Nٙv����I�%<B��Q��w�����: 5qOV�$ݔ.��1��� �<z׆���ٚOf�@�G�*��t�3c�}�"ĸ��dN��e"g�ǎn�Q�2Jħqe�zp �r�~�Q�E�m2ܥi1O>Q?bi��Z���'��B���?Q��i��S?-+꜆N��yK�kG kx����˲�?),O��S������+1Te�6�؜
&8�$�N�W2V��Iئ�Rٴ�M���L�G�y�c%��&xj�J9"�۪,E���蟈�)/�DӨ ���h�+�/��9/HLB4�*2���rH�i�P��'ĝ27�q����w�hа�+B� B@��w�)E�jM��4;Į��FF�`� T�޴n�����1��b?��;gߺ=�4I<r�ط�C O��6��g��'_47��O�#~n��KͰ��'���8��P8AN�/x������'\ay��3Q���Hqk�r��l���HO7��Q�*_w�@#¢Ӂq�����D�Nt�Q���<�1��;���'x���͂Apv��a��%@P�gڷL���A��\����z����O�u�wJ�g��\����3OWf�C�P:@�H �i�kg��B�� ��#{��B�y�^�x\��Vi:.HA/^����B�^#��'��OJ���O&�r�8	x�K������
�$�T(W�)�矈��΃Go|q�do�=w�N�Ȑ�����m�.�O���Z˓T��̡�Ci�<Ј׉I)�Ĝ�6�Q%�]hp�'1�-HeN"���4��bgH��
My�B֊+�CJ�f|h!jA#v<�"?Q�$	+���4�ާ-�-�O��{�����R�i\6��C��O\�TMI�V����p��O�7���a�t툥M��nb�\)�`��Q��XN<���?1��O��*����1p �5 B�@����y�	�cl����EG'�ua��A��~��f��<l�ly��/ �|���'D��2,E8=*iU%��A�ν�=���M���鉐V)��x�&�֌ݛ�(h>2��Х�P�����e�"-;��%�N\�!��V�^O��a޴Q�"�r�!*E�Mp�k״x��v� w>H) #�&ғi7&t�I�(+ݴ�?��l����:=�,Q�(*ddք ɖ��'��)��LjB��L-�-(F�#fl��@f/�O27P٦=mZ�VP��jΗF�� d��)���O���%�~}�S����s�����nG1z�<Q�%/ƶ���27�2_���ڤ�z����bo/I�b�}����-��`y��)'G�	H�Iȅ�{��S*�'�"Hq�mӢ���/	d]���\c��!����-Bڝ�@��c���ݴ=6(��şy�4�?Y���iE�����cmNi���ѕan�8�'r2�$,ғt��̡E��ՠձb�(d�*�Dy�Nm� �m�Q����GB�4҇C<+��a4�܍hf�O���䞴X� 8  �      Ĵ���	��Z�JvI�/�Ȱs��G}"�ײK*<ac�ʄ��	Z+t�\x�kg�t�D�7��ĸ�/^ �2��6���n��|lZ��M�#�i����(��]�ɂ��['��,t���gJ<��,�֡!�z��#<�D�e�f�c�#�%<�!J4E��	�xzpf�<��ZQQ�7퐅��9O�D�H�$�'e�:N̔�u��"��	k�Hp�+�>�O<Q�,�l���y��7%]�x@��>{^����	�X'���4O�r0�=4��!C6�ɱJh��XW�|��	N�'7��&�H�����p��aC�MYx<�mf���ቀS��p�C:0ޘz�~���+`f�)�O2�Ȋ�D_&����"�Y��Ȍ>#�����>Pp�f}�#<��L0��/RK8Xi�������4�A�v��6���O����Ȗ%�*����u��,q���>'���&�$�=�O�J�Op��Vˆ6]'����ƒB\| xdP�`c6�Il3�O����\�
�yCWE��v<D9ȶ�� �Oh���-�?ѳ��$-y=�UΛ�S��و�-�R�,�
"<)�&�ڙ ?�㢮�!Pb�<B�$ ��O����\~bђ��V�bh�T+ͭp�>�t��I9�LG��h�O��@bW�`L������yR��dÇ�Opl O���r��Sԡ�e�@�'�2���>a��* �*"<q�	�+qȾ�)���%�q���E�<�s.�
 2  ��H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �   G   Ĵ���	��Z�Jv��&�Ȱs��G}"�ײK*<ac�ʄ��	�*t�Xx�ae���$E#vw�mɶo�8c�i���.�xn�2�M���i��5�IU�A	�A��.����ڱˇ�Z�@�@'|}�#<��Op�r}��LƮO4�E��B� �\)	�X��{"�ӗD��u��<�D��k]b8��Y}R��ԁ�C��v��u]�s�t��F]��a������y�c@�HZڴ�;*��9O�E�AW`6x��d��h�d}���<DL,�J'�����վt�= �,��I�?lR)����5���B�4�K�b��O�Z���h���'@ZtGx�t��6�Z������#�@zF��&���	�Y��H���� i��0ʆ4t:̭1c�.4!��Њ�ě>�O.y+�O��x6���(�%\ K�m�Ɣ>�V�4y��➜�`c�?g7Pl�0��i��y�5�tӒm ���\2�O0��An��5T�S@�&�}�@I�;l��O�Qj��̹��dK�d��k�K��7ԥ���u��	5��HR�$q��q���=�(I����g�L���d���O`���k;���MɿDy|!Z��(���<��0;4NO<|8`�X�E�ޜ��&�'m�M��O$-���D�$�ē6��� ht�d�� Y�Y��˵pZ��(}��O�����>��'����G%
;�B	'<X��B�Z�|��'�I��� m�'6,�O(�9�* /��c��6�,Q��W��J�ɫP6�L���J��,��ұk�xE�n:D�K1�   �O�q0�� T{�E�wIN$%�"�KT��O:�@�f\'���۴�^�*#���Sߟ�?�����>�Ɓ���� ��@!�M��S������o�9
P��u�.�ȑ�2����ȓvz\�s�ʒW�$��."����ȓ4����ݻ>	t���%��BX:��ȓn�ܜ���ź)I���$ip���1;�(4)�8<��qG�pyE{�1˨�*�cf�"��,�hX�#�H��"O�1y&L\(���!Dl�,��E��"Ou�Y�Y�(�+��b�|�"O� �WA�fj:���gNj��8�"O������h����ȣ$8hy"OʼA��6��|Ja��s�<�[c�'K$�ȏ���k6p��6�`���5dV��*��]ZX�R�L�uQ���p+ػ(+����(R>5�S�ʏFT �s�B� 
��P   
  e  �  ~  m'  e/  �5  �;  EB  �H  �N  "U  f[  �a  �g  .n  pt  �z  ]�   `� u�	����Zv)C�'ll\�0�Ez+⟈m�(w��I�J���D<c��.T�I���L��qK�%ߟC��r&c��\-����+8�:W��z��� ��4!SuA�
!���K��	�fbM�7��Y��#Sj���/��{*tMAt
����iQ���cG���R��;�r�J� ��1�0k�\�#8��F�V+t?��A �'~4(��mi�H� �~�,�!c�O,���O��Oh�S��� *9�h1B@E4:�HQ��O��?iܞl�uy�'v���O���'�"0B�I� �4C�-��pf�'B�U���Iqyb�ԝ�Mc�'�2��RV5QRˀ�3�0-i���8O���S)�E��y ���|���3X�<�'�qODQ�@@�x�lՕ'����tƛ�u%�i�cf��bĢ�����?���?1��?����?Y+���t���p��T,,6�Aŏ�~�Z�$Φ�Pݴ#��hj����ΦA+ݴb�f�k���$ŒM��%�u%��xܨ�z���A��=q�D3�'��p�co� [�͡R��i��:���%��hy7-��޴3$�F"i�,�	b>��2�.���A��3Eظ�s
E"�����K��?QVh�+4$�%�E��I��4�-�30�B��"k����t�b|o��}��]��'Y�AJY3�A�z�;�-�Gl��9����M��i�6�׶4��H�B��u�Eb�E�^w������ISF�tm�4��Iæ�P��M���%�F��Ei۴R0Ҕ���|��M�v+��`߬�K`��\�z �`,�L>�S�ʏ	�����`���Q��p�2m�$�8	p���̪hΨ���Ԗ:��H�9����*�	���$�t�Ԩ�?Yctg~(��Q��1+�4��.,D�Dyׁ��4=��C�&K���rBn)D�L��cI�N�����S�����(D�<b�/ˈg�H�A�E.\c �B�:D���Ĩue�ȲcH�ȭУ�6D�X"�!�:(l$��r�����B�J:ړiv�G�4�F�7ZBD@N:{�����'�:�yR��4��9�'㚇tº� ���y"�A#	*@���/h�Z�2���yR���Sk�I����䣢�Ӑ�y���mr��bi�V�~ r���y��= x�E���Qw�ٱ���?��n�B���� ���$8*�t ��Ƴ5� =YE�+D�!E&�=&`�Y��CU���b(D���D�]��٩�.@H���H"�'D�T�c!� �h6@��Gw°9�/$D�l�牑�*w����L1)E�,[�/D���&E9hA���G�+�F����<���^8��i�m0ac�0�)��V%	:�$,D�Pt(�/Y���S�ۂ;��\�G�(D� �P�سv�,�#��9wm>1�e�'D�4��f�!��Y�t���qRD���9D��ҥ�]�Yh1%ӏYBP,!al3<O�IB5�Ϧ��I�� �*NQh�@��D�3Z���������	��N�	ܟ�ϧx	����<(v�'8����n�>X�$��Sk33�r�k
Ó\�2	C'a�J�JI�V�Q� �<m�ԁC1A��Kt�Z"s+��8$��{iʢ>���럌�I�<�I3_�j�s���X��-�UH���T��'b��S�gϐ�гy=X0���7�����HSQ��*h���&A|��p��O�ʓ[.>0H1�iZ��'��1v�N=�	�:HD� ���K5OV�tI��؟����b�pPVJ�7V�5p�\ 7��� JA�~4��tB��j=�  䍑X~BMJ�r��( `��Hp���Ƽc���K*񉌌[Q��e(RQy�ݛ�O�
g�	��T�D�O��b>��U�Hg���#�(â4���9�c+�$�O���Ē�b�D���R=a��9Zџ�����.�8!P�d�2 �Bi��!�%dAp7M�O"�d�O*�آ��'����O,���O��*����Vk�q� ��&�|�rDĦ\�i��!�8\bX�C1�%�S#�ē*:`ɂ�ʍ"�"p��A@-���̍�xd!"�;L<I���J̧*"<���V�|��/a$9٢f[=���d�O>�;xJ%��D���Iß$;AR7A^́��l��cS@	�ԍ�F�<�TES�K�"���ϳ� bZ�,��������'#���I�>	b.����].o�.�2!���y��'�Ҍ�g"�4W#(��ci^,h��b�OC��x��/eIF�8�jC�eR&Tj�hƼ,�x�'NN�⡞�%��5(2h�*i�Y;AE��?	�'���r�A�Ð'��?)����'e8����U-{� BW쎧"65�M>���i�'Q&��'��
FP�c�ٔM��I��+`���P�|�N�����#�&�Y0OG�>D� "YYčD����uA�,1���ᅏ��U������C��7f	5�^ഋӔl�D�ʄZ,)�M�¯�2��(0v�X�\�~u3��7�B�d�amZ���"�	y��<s%$�>`%&��ë���0������IܟT'?��<i@ �G�>��l��Rr���.^X��x���R�$�h�
�>=j��萎O/&��x��Ly"o����6M�OV�ĺ|�2�M��?91	�Y��Z�I�[<��V��?���ߞ���f�X� �$�B�^d�y�"��?��OJP0bد4?ܥy%�:��X��O�lR@�K/u��`	N4d�[ 
�4ݸ�&>1HPGQ�7�L�7���b���CF;?�6o�����	q��m̧/Yj���͑0�z��sH'�L�	@������	�6I��;��ܞ
~���$��Y��>u3��8\ļݡ�o��4��(�&C����I�X���M�F�3 	M��$��֟8��Ǽ��ʸ
)���j׃a�@Ģ5��?�8�S���2���q�l�6l֚��|
t�xR@ٝO�� gn[�N��lz�˴zc��з��E������>[������4
 >b�r�\9n�y�-�$3"zᒗ=@�r4�	Z~2o��?������?�3�2dY�H��)�$0���2#�L�y�'˴����8E��J�+����k)O�4Ez�OHbW���Ԋ�h��T� ���	ђ�I�3���
4�N��T��۟�	���	�O���O)�h�E&��|`��g"d�$�FΞ+L7\=۳�'��a���͇+�܉�0��0���G���xۚ��1�"3�R�R��L�Kݲ�D}��	�8�\]�ĮR4{.q�!HB
s�j�b��?Q��i>^����d�t}28��9,v|8�F� ;m���L>��.����wh`05H�%ϼUJ�&����4�?�/O��n^t}��'p��kE�,C���3ՔB7LP�!�'t�T09���'b�i�4r���X���I)},f�:�Iì/�"A�G448f����h�})w'�/TI`�r���&߸�ÓJ�
�Ƥ8��	���2�����O� �0�'���'2ǖ0Hޜ}0хO-H��h�Ǧ?G��џ��?E�t"�$w�u��Q�I�F�<��?���'��8p�Ǎ�|�.eh�+�J<�b�����?��W|��<i�w���ZB�5.:��0�и�&���'�$��k�WXfi���@��$��'n�)��#&8]+@�A�GPՈ
�'В�(s�QFh`�iGś4UV��	�'Ch- "�Fj���v�Y#9��i�
�'��
�I�6o��0��:)�|��g
�Dx��)��X����RC�:!���ҕm�"9$&C�	��l��`Y�Q�T�x����#C�	u��5+�ʅ�"�Z�ΐ6.�B�I���D��lY Tr,����O�pC��25�\9@�Rx&�B�Ϥl��C�	�zf�)kTE<=� lh�-M$hŊ˓
���I�j�@Ŋ-����3.�FY.B�I�4>`)S�E�+sD�X�F�|8"B�	ݚ�
C�7L,��aAB�d�C�	Q�^��v'R�-}P�{5��?�C�	�h���l�;���bc�B�:����=^��	e�Xu���V��\ G�M�!�Dٙ`|Yb�Lx�L��KW
=�!�$R���{�BH9��0�K�=w!�)^6<��z}``�fI�=���ȓB뮬�!/�0,#n�"q!X�jC����Z��\�s�Ue2<S��M-
�T�G{ra��Ϩ�\��M��d�B5`%�8\����q"O\�DK͒x���j�i\�C�"O��㳂�4O�<&ʕ�'�,H�g"O�Pp�N$��g��g´Ś7"O��i�鍘mѐ�㓋|��\8`"O��CL�%���ɓ㒐 �p���';ڝ������~d9�#�1e��[cM5�x���*�L5�W�rͲ�뗠�������Z(%2u��7p�Z@1��D�<� 撟m�Vൃ�*7�D!a�-�E�<at��6�����Bӱ'p�c�X�<y5��x갯�12��hIm\Py�E�p>Y�S3��*r���]m:U� O�N�<� ���/����`���#=@�+�"O����Q4w�H��6�[�z��g"OpYp�e�W#��S�!W�Z�.U�F"O�E��h�Sͮd"�`[�@Ŭ00T�':R���'�d 4E��4Av���DA�ZO���'q�l��/�G��L�w��
Q�x�{	�'�:� C�ìt,�J$��	F�j9��7�d�i!�G5-x�h[�`Z!J�b���\Y�8����5���	�/ (��3�� !ßpm�e0W�=@2�F{�%����$}`B�I6�9�͞	� 4¤"O�}	��Z�/����$L��I��U�2"O�[�� �:�4�
�	ٺ���
"O.�$�۫N>fA����c��ٻ�"O�����.qNrQ�d��L�H���"O���A#xgx9�Y�W�@��'���y���FkdI�Ü95�DA�N�yN���ȓf!�IHuE�9F6,�A�(l�ه��dY S��%)�0�`Gf@$gr��ȓ޸uص&T�l	� �&��B����&�09�l�!ɪ�P�C�(M��E�(2UL�7K�4a� ��j�>��'!��(�q��p$⅐Z�N-M�/�.,��+t�Ď��d�@}����5O�����$��1��
�#n
��G��/ɐ	�� ���B��R^�,BEL��#�X����Њ��U���L��O*?������@
��i��p��0<B*�ψ:d�B�	�����ӊ/l)F�Ԡ��rl�B�ZBD��T�B*n��YrKڐ{H`C�%���)`�C�#���z�N�`�(C䉈H><DKD��8�m� �9KZC�I�y������ӏ0K|�@��E�%�H�=٢��_�O�F(b#��)P��p�˪��<p�'�  r�& �(�@+�!Xh$,[�'-���U5jW.���ؙW�l��'*4X�	�8[E`t�!������'�BD��qX�WI��ϊM��'a��*��[&91�jF�V��h�}�F�Ex��� !D�P����)5�La���Jw,<B�I�0�-ӑF�,jH9� h�'�&B䉻i�XQ���
����+� 
n�C�I/\"�:�HP7���֥ٓo��C��9:�bF=�ƍ�A��u��C��4q��82�-<���w#��v/��EK���I++� G
�="����A�ئ556C�IQg��Fb�^ᶍ�E
�nC�,'���p�lM�q�Fy  �%[�TC�I^M�B��4!.�I�����C�I/�2�pN���)���E`����:���[c��*��&Mj�r�LI7R�!�dG8 ��S%�%t#�M!3lDK�!򄊔w�1�F��.���Ӹ0�!���_h� K�kt�ޔђI�5!��ɾH = 6��#����Z	"'!�$�*ka����{�!D�ՠy�ўL0P%%�'U�Zd�c�	�/\b�!VIA�R�n����b�2��P$%�����'
���ȓpi���c��~S�5�v�; ����=@z��b��E�����7(����8�R�	G�ނg+^|22�J/iZ~�ȓ(���m	�]�|*���^�2��ɞ'$h#<E�D��.=�Μ�b/<^�&�a��Ȼ#�!�d����P�$��"�ȝDz!�� ���1�5i4v-�a��s�|��C"Oi��FG� ��b
A� o��3�"Ov�qa[:��ɋf�޵\o�$�"O�Ћ�d�-b�p8�f/H9N	�eS��8�#�O.�����7�LrD�A82���"O J����KdQ�$��}%�<k�"O�s �(}0�P#�%ʦX=Duaw"OؐfÑ�W�L�)R;��	�"O�1KcƜ*D?���!pEZ����'��A9�'*eA¢�}��t���XTHy�'�zXR�	�%9�v�Qh��y1��	�'��8��5fֈ����ɩ=^�I�';�dek٤����X�+��I
�'�*�� ��^��!�$�x�0�'ǌt�\�!������t�K����\"Q?�Ì��N�`6ҎH>x��M7D�L��*�2Gb��d'<�*���(D���/��h'
�(f$�2.iFD#�'D����n�|�jI��W�=����)D���D:4 ���"#U�9� �%#D�8��,�!oH�Bm@�"�:X�Q �O��	q�)���#���i���7K�4	��;�'nVP�Pmʭp��(�W]�fdQ
�'F��y��*�<T(6��uP8A
�'�0�F,�k$�@�.o��u�	�'�9c��D�q*�VHA��'�2UZ%GȊQ��U��E^?(�.O�DQ��'@vM�ffПW��PC7�ZX�R���'�� @�'F-���&��1T[}��'"t�!L��=l���MDJ٣
�'6-�a�:3�D� �Ӕn�ZВ
�'��:�-B�F�2�	�
��bxm ����m�����gW�`8#���/���ȓ;v�@q��9s���b�5�|-�ȓ9u��r�C�>A���6J��!O��ȓ=vn���j�2V7���b��E"$�4Cb�B����Q>Y�ȓv/������� ]��`׀	4��D{�L4ը��hY�@]�;�d�#0Ɩ/f��Yp�"OF��"oT�x>^$u�?�$�z "O\��&O�,O*�K5D�;�`�!`"O5鷥�f�r��1��[ ��"OT2�1/j��$��*3��"Ob0 V�@�;!��Ѫ޽G,.����'
�C���S�'�ł��ݢD�bͳ@	χ$@���j�ve�2�V�x��Ђ����X�ȓ1��iCQ(��%���h���z\�Մ�S"ty�Ζ���:�"�i�",��W#B��u��Lp�A�!J�\�؅ȓ-�}A��#LER(��N�=@S��'s���=.�e����%s�xsw���-����)g.�IF&�$Zz�6�V4I�rE�ȓP\T0pތI9��J��J/�܅�,�M��:K�d1���. �2y�ȓqZ�	�J	�%Ј��V
��,R��IxӬ��O�>�k#䁮`��̑��<P��C��$�����7��%��(G�4B�I�z��(q�j��H<8C䉶	{FŃ)�/��`�"� i(C�IW%��#���|��#��`$C䉐X�1��)ÄɄ`�`�Y����=	�K�i�O�Pر���P��
�a�(]���B��z��j��8|Z�Tջ��B�	'�r�E�xf��h%`�*�hB�)� r5+�KV�+� �2T@I8E)n��t"O�z��!�.|R�ݎS*�Qs"O\	C�"�H2S�N9Q���V�'���ۍ���jB�A�U��e*�����G���ȓ@cT"q�ċJ ,��3�W���A�ȓ|���.cX��� �<Ā-�ȓ^J$ѐ���=i�t:Ħ5kXm��ZA��ZccG�ph)ZCʔ3/f�+D�x9`';;�(���!������<Y���d8���!-�O0�t9� $ �D�.D����`a��X�d�{�t���M.D�Hj1G�l5�]�rG�ݚ�y��+D�H��#�:^��uQ�pPU3&D�x�gbC��������Y�z���G&�O�@Q�O0eF�**׸X�Ĉ	�����"OF�qE��!b>��Fj�=���Cs"Ox���K�Z.zPis�M�-��<�U"O�����N\}\�;6� 6p��l��"O<�Bu�B,@�
T�"	Qke$a�"O􀨔���A�8+�(P {T L��ɋB�Ԣ~����1Z�L��;���a �Pg�<y7ݤG�:�x��W�8��V�l�<a0�S"MW��S@ߦ�jP30�k�<��o�J�n)����;r<H��d�{�<����A0̸
UNT�@l��N�x�<�T��8O*Bx9�.�L%���*Z��pS�;�S�O�蚇�C�0�(�I�Iĕ�d"On�4hߢ����c��5EcG"Or���ؗB����o.\0��4"O�����N�'6��� N�+@�(�"Ohpȃ��%H7-O�F��H�FO�ibb�-&@wNY+R
)+��O��'�X�'dȠ	��R>L���?)$�3\�<ͱ�g7k4��xЍ� �?�Q�̜�?1���?����,LI�aQ�SZ"��|
�E�2gbH�b��E�Ҭ�!��]�'1h�5%A�6���Q�6񩌘hI�x2h�<\�HCAL;W��	��Ob��-�=V���w�^� Ī������/����0?��N�%���6��d�R�SC�Rx�R,O�Dpu��Hd4`Ԃ�B�h�ȠS�$�3j��M+�d�9�?�(�J�EH��f���,0�������6�}� ��
���ʏm��@��\_�Y�O�b̧$c2�1q�ٛG?�qdJ&�N}�;�r ��:#g<��"^�"~��F�}A�`a �A�FŴQ�`���<�'��ߟ���i~J~��O|��@^�~�hq�O�_z�<k�"O�]������! R�$}zȺ�3�ȟȋ׮Ҙv�be����(�#tL�d�O��L�n�.0�Eg�O��$�O���ۺ;�m1��ӄ��6R*�a�"�=Bf��v��$z���
ΆX[�E����	�Y��z�k�R���I�W����'B���9���"0�m@�1FxR3;�iH&��Nl�Q%I������&��'�"�$}>9�%�5��ZP�M �^���5D������	=��<K�L�����O�aGz�fӎ���<A��՜������ .[^���ʈK=�y,�>Y2�a���?9��C��n�O8��t>�	p�:Yښ�S�E��:���V8e�ny[�A�9��y�0\\��5�:�$�8hG�8aq���֝j��Ի�-@Qc�m�$X�-�,���*�\������O�H�I'�`����W��`�T�O��=��D��,V�� �W)H|�h�e�s�!�č�gi9�Y�nz, ��*Y�剅�M{���'����I?}k��*2��=7�J�K�z�3�-'D�D��+�ho�Jb�#Fr�[��:D�00D��U{����&T�&@x 8D�	7�̏r?B��ԧ.s��Mz��1D�da�45Ai����-2D����.�&G��9H���jl��i�"$���E��#<����!f�&�`�c,�"2c~�3"O2P� �B#4�t
�'U-Q�"O$�"5��#��[E ��S5���'"O� X��&\	I�H�d��}2"�1!"O�-��fɞ2��A�i��Q!3-1D�<+��
�v�<����y�(�HB�-U��E��'�:D3i��!M�dɢM[��R�'r�������� ��C�It�:�'	���� n#���sA�?�R�s�'���7���|0����ȍ/&z	�'-�H�U�P�u�~]A3+��*|�8�'�̅åa�Sp���c��:B���#����	��`B�捀9c��	�hR,&C��3^y�Q��nժR��t��o�C�	�4�pl$��C���&O�B�is�5{�Nِ6D���{*��7����ah�A)��"�m��ut�D��Q,=7m�O��`>��q!B�\�H��(P�(J��0�	�O��{R��O"���O�� BG�%�h-����#�l1�.Ճ�u���z����Amc���� �ԈO�����(l�����K $+�d��:�8��$`[�@��]A"�+/�=�IP�'�`����?�I~���&7���g�3�T��iW��?���������pBȒ�e1�Ks�M�t[��w�1�O�'S�|JTc1{N������&^؍r.O����O��$1�S~R�F$0ap�*�ѩ!{��
Q��+�0<����2�*T@2.4�}+'��6T��On��v�x��	�+�4%����?Q� @ٵ�D+-��ɻ�~"�����|Γzz2��&&�S%�qا�G�Pb�E�(���k�d]�0^�OB��4,Ռ]U�a��g�ܘ�f�^���O?ю�9O25A�癡-�0�X+;#�R�r	�T��t_�f��L�O���O[*�Sb��>���m
�!��'���OtK����g@�Sl^�+]���&���v0���>��'��'x�t�L��4,"~P@C��n���H3�ɖ'��3H�Hы���Ϫ�ab.�0����/�zY��u�y�O�s� ��f0?q���D�
��`���{Ap����� CD*�'�����O����V��0h� ș8a�$�(qC��(�R�Bl?9�!�I~ʟ�G�=P���, �σ�uC��BX$u���T؟�5�̴/v��F%�B�J����*D��)�a�##Z��!�DIcHR�+Îj�(��*�dU��O��禽�ւ���L��K�ec$I GC�>iM>�)O\�|�D� T?�T�ā�>7]���V��N�<)��7Lâ���%�8��TaQA�L�<	��Ӂ���k7"�1H�:�W�A�<���81��϶F�f����~�<Y�N��p!�&��R,�ƫ�s�<��圯~��ͱ�(ъ~��X�o�<!�J�ڶx�oA�Q��ԭ
G�<�� R�Y�*��\����C�<Q�_�dP��� p�J���Zt�<��*	z����e�,iN ��� n�<����%lBl���];#n���PC�<YC_i���r #޹p�mK�I�E�<���&#����*;k����
�V��_@T��6IL6�C-T�~�n�[E�!e(13N��NH��ȶ1Q�R4G=�\hI� ��<�S�:s��p�K��zt0>�X�ڐB?y�А@ʈ�p���f��VI�I�C��eXp��1	�)e�P��Ue�3���2e�Z%�M�E蛁d/P����|"���2X��[�ް~;0�-"��܄ȓY���{a
Qop�3%gC*zw���1�Na�&�@�6��b�#rZ<�ȓH��p�ըn�|axOI�_�����"���"�*fL��kP!I�t*p��I�dC�g�A��|sw ��xņȓ$1�q�
S���Z����h�ȓ,��Es���]1��Z!���8.��?p�D���U>pSAM�8���� �u�{~��o���!�ȓwd��k�'q���#���@_fE��"��� \�)��t3�0G��݅�5YD�Xp�B!|��A���).Vh��S�? �|{����A�BV�� �p�!�"O0���D R�H�BP�L��]�B"OH-�#Α��:��f��N�b<"�"Orq�N�;ٔ!A���!�8�چ"O`���U�{:����J�Z{8��"O�p#s��#j6���P��\�Ⱥ�"O�X��I�� ��5J�(mD0�"Ox9®��m	 � �nQ�w"O:=I��!������o�.��S"O�X۶�2�2M`p��M�jx)c"O ���C��U�!p5�:1*O�A�kQ���G�+<PZ�'�D�0�JW���V!� 5�����' �h�m�1Z�|]b��уd�4���'l��cUT�P����Y�csR�
�'�$��`�=6��b���c`2��
�'��閡�.IX>M�"I��[p&y��'�"#�P.g��8�̪{8�y�'��壖�R�T�����tr`�j�'���#���u�+o��.ndar(=D���Å�X�c�*Ŀ>Ul����-D�$�'M͊_��!�qUV�I#�(D����`a��C����sc��U�'D�l�)K%%�,|9�(K'pxx��)D���Č2 ��ቼ�H-�#A'D�����z��P!D�==�&�Ge0D�T#$ϕ�6���B-�H���E�-D�ؐ�!Wb�r��Q��ȡ#'D�<k���GdԹ�C�|G�5xD"&D���Q�J�"h,00��.?��E�`#D�d���Uc �?U1��V- D��ꑅ�9_dj]� �;_Tx��'J3D�\�Fk]����*��ْX�dzu�3D�� �وr��y�*�:	�`�%D��C@�ӞaT2A�7xX��ja�!D�HՍ�
]�6�c���)�v��g�!D��b��[�y��@� �ȖuR,y��2D��GdD�H�8���	��b�/$D��S`-_IP�0�X�M����B=D��Y�+G�/�r����P��е�?D���ǀ�ݚ�c�p�:����<D�(��
"{�d��f�<t�P��H(D�����҇W��h��N�+k��9D�4�\�xo�y9e"��pg�7D���F�87�t�5V�Y5�11�) D�H�#N�:�|�7�Ѐ���)�*D�t�!̌\�4%���S1G�hg)(D��"".��@<;uaS�<��L�j2D�D17�T�;���dj�����i�C>D���e
C W���30&�0�x�7�&D�<Z�HQ�!�LPSa���N<�D*D�HѴI�^��
#F"1D��(D��+UH�i�.HZ6���B��	��h'D���.�l�j���8�\�3'$D�ph�5q�y�6�]�'N�Se"D��/Y�Rh�&�X�K��١ �,D����́>�H0CF.[�G�ZD�A)D��AĆ��p�$$2y��a��L4D�L4�H�(�ŏT���5��0D�4k ��1��8��]�#y|č1D����,��T������:b����<D�@y#�R�'>\���@�%nQh��� ;T�(�"�+g̐ �J����[�"Ol@������	��\a�"O� 
�3����̀�_�4�]�Q"Ov��m|����g�66ɢ)�3"OV�t�@>@T�xA�4��P��"OpA)!��"���&bS5=��� "Ov(��H�j;�c��	-����"O��)BD� 3���@�xـ|�"O��2�L�0hbA*��ϼ}�q"O�ؓ�V�@�ji��H�%����"O
��A��~��'����X!�4"O������!O�T)뱋�<GވHp�"O(���_�6�jq떊o=�m�Q"Oȍ�挕1�>%�sd�6�� �"O.-a����q�V�Cd�B�.�̌��"O�D�E�����b�Q:<u �	"O`T�6!96��V�:pb�!"Ory���1*��D��s��a"O$�h/�#�hS�LK�:S��R�"O��A�p�L�P�)W�x�8��"OF�H��ۅbΊ�(d�OT�v�!%"OT4�wi_5-�j�(�L���2 p�"O�0�$��]s��I�Ӵ0�l��7"O�X�����Hh�jY�P�HH�"O�P�;2���� 56s�"O|��a�M=H,RR�` ��"O�BSՂQ�<0h��۳��F"O��:B �
[������`�4�"O�0ق�8�ґR�

4T.Ɋ"O*q��bN�f0Aa��zC�-C "O9�f�%����SA]+:Y�r"O���C�`�#�O�Z1��K�"O<QQ��#mTZ� R FɔTۓ"O��tNN�}��2��e&��y�"Oy��ѳ�����M#% �Y�"O@�&ɂ�������]��"O�y�7��V���PNL+~P�"O�!�]JU ��F�K�jb���"O�20�
v�A����x�w"O(�@�OY|�IPAN}�c�"O ��@T-3��|p��1�
�r�"O6MJ�m�$n�:Eʒ��/v����S"Ol�롢�
J�����	/�X@g"OJQ��()�a�a.�&f�P�h�"O����Tk�2䣄zڒc�"O����l,B�c�"!��
v"O p���L�_�R}�7��<+���	�"Or�
R��4���r��,I�����"Od�[c-�WP��q�Ӗ8�L��G"OZؘHͅX����'(�H�p"O�!�r��?��Hd��mkJ|��"O(��Ί�E=za:d͌�%L�U��"O��׋t�\�@��kj�Y�"O���t@C;)N��"w��(>�y�T"Ox� @��"L� �q"����r"O^�&
�3X�+�a�/�&�ӓ"O쨻�A���Ab+ɞ\�J�R5"Op��&�Ў&�H�P�	 �db�"O�lSn\�E���@�Z�ܩ�"O�xS�lY6M���Z��r�"OVz�$�3��hR"KI�$�^��"O����ɻ�J���+�;�����"O���F�>>��0�Dj�x{&̪""O�1ؐlޱE�X�ɐy_�86"O�dc�$0��Ԣ[�&]й�v"O�a҆E ]��T� +=\h���"O� z)��-��Ē\�� �vU.�"O�� �@Hd�)\�qG6���"O�E��l��m��I���Ø+I4���"O~p�e�9w���@'�ձp.��"O"� ��Lj�8sKU�jK��p�"O&�������Ͳ�J�>��'"O@���=>C:a�����t+ؑ	u"O�,xC
�"M�p�DCQ�)�� "O|�9�HͼoZ9I�Þ�D!��0u"O*x�a+��yȈ^:�e�&"O�\B0b�P� `p���\?��$"O��5�sTlA�"�|�A	Q"Or�I�JV�r��أ�+_n�9��"O�1�T쀱n&�4����D^$�"OQ9S�׾=��$!�*��gV��1u"O�3��;�����
wD�~�<��^�pz��;��P9Ǆ�b�<I��E�D���'��8pzT#�o�G�<I7���h̊'��&=��B�@�H�<95��LPZ\��*�
S��x"b��<Yu�A�Gz±���O�n����`�<��ㄞ/,^\Jb-QG��19w, [�<AaY2{
��� E?�vu��n�r�<�᫅�����FF�(� a۴�w�<���R�o	��P0A��p�03��t�<Q�ȗ�w~~��&i	�1aTz�<Q�W�i�(���#D��ȫ�DB�<����%_�����H{��$@p"|�<qJ�L٦�@�̕kjuX�g�v�<��AJ�S^�"vJ�G�v��t�NW�<)!�H���HBv�Ƥ���]�<Q�D�,�� �.O��7@C�<�u/�8eZHi���W�X�L@�e�<���Q��\��^8D8R��EMWm�<�q�G�a���SI�*$p�x��Q�<����z  M{��K�Tb�Xg�O�<� �?}B��V$��8�6qhO�<�-B�[�6��`Ǝ�E8��ڔls�<�$�	u�e�2E�q~� ��m�<��]?X����d��%��4QSxB�>G_�w��D}�9*3dq<B�I��u�rD,9jNH�5l�9�<C�	c��2gH�j- ��n�PdrB���D}HBШ2f�܁#+�5_|B䉘r�`ॉ�=��$�t#-�ZB�I�b{�$XP%w��HI�'�
�XB�	.$�u�@B��Oq�d�4�!B�tC�&p(�bǀ>�|�J��d4>C�I�
D�(��"n� ��Ӈ�?0C��2\�X{ �݃ ��P��,ԋq��C�ɟ_ն�Ѣ���]6Ҹ �MV�a'�C�	�+n����(��rAC�kԦC�	
K�l�`�ŕ'q���#�ǿa�PC�	"h�s�45��B�-FhC�ɼ���3jr!� :�a->�ZC�I�B�R��r��%O�F���ߩ]3fC�I�{�!�D��~� YBW�If��➠*� �m?j���Q4*�����:�d�.�T��T�Z���c��0$!!�$N=xٺ��������pf�7U!�D�2Q,���⎌r�pX�%�*M!�W4s��aa�-)�8���E?�!򄃞���XW��=o�9�W�Q�k�!򄄨�V0뇫|3r�HuL��d�!��-�8�+��Q�8(�+�I�l�!�� t����m����=_����"OQ�fhU.8�P�I�ܙ(�tض"O@�[D��PT9�(�d5V`#�"O�`I	ܵ).���(W��Q�"O��pJ�&G�8�K��;Y-ps"O�=zf��8#hLa@�H"��l��"O\Pm�����dѠ|�h��"O�|!a��X�x]a ��y,��*�"O��B�hA�I֤haAW�r�y�"O�Y"�JW�)3�tz'B�H�h�"OҌ	`�.F�fX�qB_���*7"O���P�6�O޶��ʇf�<9��Q�)^����M�[g�krM�j�<�UJٚs����
�,�cq&�O�<!/�1����FcE���1;�&J�<� ,��Hj0�c��(x|��`a�<!gςRDʍ�2˔%M��G�<Aх8t[:|����&ȶ��j�@�<9D��qv����Q�S��}�Rn�V�<�O��!� �:��2(���o�<	�˘iȑ�����Q�~�A��o�<�Q��-�y�ǁM�1X����Vn�<IR�ʺu޸�a���4,G�� $��k�<���H<0��B� 1^��+�!M�<��� d�|��sH�+N�p�6�E�<90�������A@o�xP#�j�<�D%1e^8�G5�,�S���N�<���r.�	�b��-l+�*CG�<�g+�_���SQa�4@P$K���z�<I��ɏ!L�BE-W�{��l�t	O�<�A�*
ީ�w�B�O႔aA��H�<� �C"p�@�B��U�����VH�<Iׂ�:K\�[�o �%�r)r���G�<9��P1)��M��6����~�<)�D�<���8!��l��l��N�p�<!R��xN��
���L��ð��M�<VfS*R��� A���K�L�<�CA��f���4�E���Y�E�o�<i���iZ����­��X�!�h�<Q��
:���K���3�쁃6��j�<�T���p�x[eh�Y7�ѫ�ȉ�<�ӧَDq�,�D!�p�Z���B`�<ir%Q9��!��jݵr���[C�<��l�A�]F��T��HN^�<)���i��Qrf�	t�&�q�[�<�%����F���0�H}�<�UL�]�P���G��u��n�a�<I3j�i&�t(���8�L���a�<��Ԙ{f ��r��-eG0Q@g�]e�<Q'(K?j�­ a҄xk�p+"G�l�<Y%��5l�Hw�ārX-���Vh�<���R1Pd�fE� ����A�Z^�<��
��8����10�
1�KZ�<A���VB��!٧U�����]�<�*� U��aT�ۼ>������Z�<��e�h_L��D�3�v���+V�<�å�vC��	B �!�b�8g	R�<���2�ȴ���(r�����h�e�<�Pa��A� �Q	m�@HCi�W�<�1�^e,=�v��SE���CV�<�1��/I�mz���0DD��Y$�(D��U*��Kĕ���^���ડ�5D��3W�
�2G6A��Bۯ6`�v�2D� �D!��$���8��-=D�� :]����:>
5*�	��$�8�"O8U�c��(>�|AF�*2��(�"O�a��
=����儹M�<��`"O,DcDf
>q�����Ec@�h��"O�p�0lՒ!.��F��,"I��"O���4o�^�*�
��Y�ܚ� D��K@)^"zԆ��̈�>NTH��,D��"��[�r� d�eÄT�F�Q@�(D��h�KԲl=-x�d@�bda!��7D��#�	��Z2�T=���HU�5D�,ÈN�)DQ�Bcr� 9ѰL3D��K�a��"�PѲG�ѣV�ʴ��1D�Tà��!�X)��*X>v��0%>D��J��
�T��P	��R.gN���� <D����l�7_���m�n�)��,D��8DJ�C<؈2r�B�|� �p�g8D��
U/��H��z5�C&T��<�$D�<�g"�=�=�₞>:�|�ơ%D��H��?W�>q@�
A9I���#D�ʤ-�-|�4<�����?���� D��
�v��A��/�IE��[��2D�|��#I�)1���"(�1�Y���:D��	BE��-�|�Ć	"WDl���'D��q��5<�ެ*�.J/f�FIS��8D�ĩfbN>9��� "��"k �ZPg&D�`Z�'_�:���Å�"t?40qB D��S3C�g~���)S:�6Q�
9D��1���>�r�hi�	2&Vݫ��'D�����P�����Ts�U��L(D�\Y��;�\�ˋ�P�0���,D��� 4
v�MIF-�*E&��r�+D�0�e@� ��BI�� � )D�,�Kd��9����jg0�R��5D� �� ;B:ZAq2�[5L�]؁�8D����fO�?�R���LZ�!���w�<D�ԈP�A{d���gG#$��,�D�>D����bH�Zݰ��ui�*�lq��K;D���V�ի2ClaYs�ǫkn�|�f�8D�H2�K�D��+�Ī[�<����2D�0A�k-�(�q�,u)Hɠ�a3D�ؘ'
�7���A�Bnl8��0D��z���mP��N��^�XT�!D��"�ɥv٨�bQ덫>e�5�!D������'~���u��!Ge.h��F D�qJ�|Sɐ��$C�dU���/D�\�G���#��PUL�z���2�y�̀�zWYP
Ϋ{�V��b���y2�6zc�9�)ʻq|�tB6g\��y*̇P�����ͱ�<W�1WM�C�L9����.LO.4�s�P&d1�C�I�t�JT���̭8���ss#2K��B�I�t�a�d��%�nd �I�g��B�ɣȤRk��`�cD�	)G�lC�I!7��:��G�HD�9y���FfC䉠b(VY��4i�-4�Y�<YRC䉌hٮ AT���=K���foƑNS<C�"�����"�:�f\ ���5b2C�	��z,9FFѪu�|+�捌$�C�ɠn�!�����\N-�5�ʾ0��C�x:��礒 5)�BҢ��B�I�\欳A+���p%�, ��B�����
��x����ۨv��C�	�Fm�\20�(i�x�Fa=)lC�	2x�b����Ԧ	K�\���O�s!�� ��7G�b'ԁ�@���=1�x�a"O����Θy�Yb��J-x$fQ�"O&�*�[8h��ʒ�Qz���*"Ot]�C�P����&I�H�*h�"O��:��i톙iuF4-$�+�"Oz�y �˪+P�"T�۪"�9��"O�-�����TY�e�Uj��Pаx�"O: ���@�M�0*�Hr��1u"O��p��	2�(a�Z*u@� ��"O�a`�Z�2��n�=S�l��Q"O�M�#��Q>
���#ϊ���"O	P��N)wF���#�C��`"O���RQ�hX>�#d��e�p�ӧ"Oi�3��Ki�P��&J-���#t"O@����#��-�@2�^�ӵ"O&���
>��`�D�R윌3"OJ�Y3�Q�c���v�H9�"O���Q"L�.����Pb۷m�i$"O�q��<����b�M��@�K�"O��B���'�R�*0'�1r�!c"O$U��D�	R/�|
��/x`��"O���e��N�����ڄV*��v"O ��&-�34�-"��W>��� W�<���[.�~�	�I�EQ����m�X�<ik{��M)���?B*!�P`JI�<1aւ(�f�A&Z�0]�����@�<yR% F��m(D���j�I^�<����2}���0��_�u�B񚒉�c�<	t�S+�p�kw퟈ ��R�&�U�<��ߥ_^&���C�[cҬ*��X�<��s�Hp拖
j�R��O�<���?@����ʮx'��[��Pe�<!G�ߏs���B7�W����+�c�<��`�d��Q�Mϸf�x�q�IFc�<Y�k0b���E� ]|�c2O?D�H2 ��U��Y�ӥ�<O�Z�ӄO*D��U �-e%H#Tɚ4�TzW;D�,!��<��i���!7	Ӥ�'D�j�%�+$�(�f��  �5z*%D�<���5Cx��7���i��;f�"D����'�o-$�p� A/+]6���<D��y�(B!M���vBSC~� ��(6D���W�1%��HȲ��`��;��/D����8���e-V�� Y��8D��#AC�=Rhh3W�T �����(1D� 2�%�P|җ�ڠ�f�?D���Z"u\Xx
��P�a6�rs/<D�,{�m�]�R���Q�w��;&�5D������_��`��?RL���F�4D�������;t-��ƀ�3� D�0"0/M�B��y�F�\81�,�BO D���b��\9P���?n��P�/D�8�GY�U���df��g�|P�.D��0�i��B+$��S
��7�x%��(D�H@СD+}�.�hW'G.NtuBƂ6D�l!�"�&r�Ұ�� O�i��*4D�0�"螞H�B�Se��&y_4�"�%D�\h����1;n��BŁ�ig"���'D���b�W-;��a3$�U�p�q�%D�T�g�F��d������!˷-%D������/k���3F1y��!���"�,Y�Myc�ǕE�)YQ�\���O(!�g�*�x4 R.�(��"O�4hn�]z�uIbL��/_(r�"O�K�A�0����+�>9J�\;E"O� ��r"�l���b�j��*��a��"O��Rt�S�b^ڭ�5���c���{"O�`1�H��bh)D�M����u"O�dX�KF�>�)�jP�4
�"O�,sp-9EhԂr	V�<�TD(W"O�'�@
4����%Wq�I`�"O��(V����,Mq�m�/pf��1"O�L��#C:\��Ջ��S7�"���"Oⱹ�(�� �G�V��"O���,R�+Y�%��/J/Sa�aI�"O:M�AI���ps��9:S��B"O�L�+� q����#NH=b�"O��Q7	�3,X�H���,Y�R��a"O���C��h�Y�\Ҋ�"O`���M���@�8&Ұ�"O�UC�ꊊ d�y2�OsȾ�0"Oz��H�&A�0��vN�8�~Ts�"O���e�X4TCfC�1g0�3S"O����L$��pa�`�-ÀY2A"O&5K���#C�BqA��2�1"O:A3�#��b��i�n�@�āg"OЍBE��3��ճ�K�6�J	Q�"Ot�SW͂��V��H.�8�@�"O����2[^D�v���M��l[�"OR�j�,8��m������V"O|�+�M8�V�A�G/OPU!"O�H��t?��HA
�3�J0�u"O.�rʖ�2x0jV�]���P�"O�(#L��|1�
�R�ָ��"OP��`䒌fl�X�v��Rڞ��"O�i��'�$��$Y���
n�L)�"O�E��̓�gMΜ��A��r��(�"OB�R��ޚ=�"���ޯL�D|V"Oz=�&�ŧZ@�ʁ�� Af"ap"O���K@6~�tУ�*� �,D.�y҃�5�D��1���Q�D��'oB�y�BF2=��40a
ԋ1��uY�D ��yB���h�.��ăԦ!��ܻ���yɄ��|���G�5zab`�Ժ�y��"�v�Z��N*�,��W½�y�o�	�lrjǈ �\%XWG��y��ݶ ��� ��p�$�Rǭ��y�lW�"��ò�ݜwd�� �9�y���b���Ʉ���h��H+F'���yB��cXFM��R����*s�G��y2j�#v����gW�6l��a芎�yR#� x;L|��g�Ԗ�q�M�&�yr�S�X��4�vE��F ��`�&�y�	��"t����}����OZ�y�B�4XҸ2��\��r8S�)P
�yr��*]�tx	����5�� �y��ޑr{�h�
�L��ꄉ���yb��&^\���ַ?�qR����y"̋,`�|Wޫ4���ʐ6�y⫙�?��'��/��I�c���yB��"F�N��c��$-���F��y�G�*���7e����h�AY��y�)�X�PQ��"3��������yڇr�.�`�!\�wV��b�	�y2�ø-�±�F�'w|2#A�yRo� &4L����r:N�;�I�8�yBg�d��݉�[* � ���g-�yr��=~����Z�wҬ��2�0�yB�$2v�8`��=�Z�����y
� 2i��h̉>q|�@�-?3f���"O�A����}����-&2}�D"O� p�%̼���jRF~���"O��S�i�I�<��G��.~q�E"O,L���Ţ*8L��6@٩J�n)�V"O��ju��=t�Z�SOǁ?��TF*O��*�a5`R�����{DAY
�'>��2 �'~�
��U����mR�'8<�iS�ۦ����ӡ�5��'�\�x�P2�L��GL�p��'�dĠ�AX#l,(ta��1�P�#�'1$`�$�
�N:���c�L6&�fp	�'���M+��`��� �u9�'��(�Hڹ/Z�����)K���a�'@�eB�,Ŀ!@rMiw�S�I�dz�'K�@`��+X�"����ʢ,cR���'|�zQ�'_?Ɛ���N(��h�'��8X��,:|�(��]+�\IH�'���w)\U2�r��P�O3` �'=y�'l$�P%��a^M��1Q	�'Lz����Q<X����s��	5^�*
�'�>�Ӂm�,0 �
��!4V��	�'|"��!�Ͷ~�Y�fU	'�� r	�'��� �&��V2�e��C
�����'��L�K����p��a.���'��E��#�4/��}��
bL%��'��q)$
��p|B��6
�
��'
��ږ�P�3`� 4����'su�A��D�����-�nPJ�'�}��m�#Zvj�Pl�)hb���'&�PAeO8�$���h�%C)p�'�2��`NH�#�& ɤ�۠m�
�'�~h�!��M5��!��|�
�'��i��G��ړ���}��y��m�01�'�l�J�S��@��yb��+/�� 6']4p���:��5�yrn�&�䤚���j�=Q�P��y��K@�1�e��_��ՑѣJ�yrl�W�&���h�Z��H��y��%�&ݳ@�%f61K6��0�yB��,%�l\q��Z#t���FLˊ�y���6e4LP�j�CdtE*NG��y�`4k�1�V�`69��H�y¯��G�����	%V�X��y�R�jon+5@�(���ہB��y"Y}.��C"�ly�GS��yb$��-�e�U� 5a *)3	2D���ҩ{���Y�m��!�F/D�L�Ǡ$R~�iAQ�Z������+D�p��$-b;�M��Rrq�t�*D�L���8�LMxՂO-��H�5c(D�4#�
�#!LPm3���\U��#:D���F��^R���fͳ b�Q6�+D���-R�nJ6�uǗ%g .���.(D�����Ĳn�d��Q/;�6Y���'D��I�i4�Bbv	9��l!!J'D��
��]9͞1�ƏҺK
|��n8D�ȁC"5��	��R�� )�a8D�l�$�@�i��	�����V��9�e4D����\**�x=tcD�]p��H�4D�̪��6�X��q����Fp�v�0D��ye��J�ĽP� �c$x��1D��[P��[�♒���-+��x��0D���� �Bq�t�Q�E=4�ԭ�wf0�I~��� ���TD�%R���itbR4�44!�"O�����h�����/
*g+Fp��"O���*7W�y�L�H"�Ҕ"O~����t�rx�Ek�9�UAE"Od��O^���s󪌼9�|""O4��
��!%��i%��%^�4+�"O��r�Fg���0aF�6�<pt"O�����7_�@�`�;tH�"OD�R��,r�`�Sr�8��0"O`��5HC��ڕ�+�L�%"O�-Am8Cv���C1v�pu	�"O��@`NF�f�������)g�BU"O�yƒ��:����'D���PP"O�%��ò���'b@H�8�"O���v�Q�"(Z)C�L�J5V�C�"O2�@�i[�#�@,8��U�K��|ڥ"OH�7� 4*L���+o���V"O�X[1���8ʠ�@�[
j��*OF2���J2�Pą +�^��'�.�kS�Ӹk������U�l�Z
�'� H0Ƙ
@Eԕ��+ÍN�d�' �#`��	!�U����z�,+�'o
�#�Ο��,
AKF�aM�%��'���*ĚOj+W�R4g����'O�Ԡ׌�:p�D1vި,��a��'v��j3Jˋ(�:,��,�p�e�	�'�4JL�Kvx�%.��c�-��'%80��[8w�RqqF� ��X�'���
G6ڌa�iʩ1&���ȓPP�B��
J=i1,��[A�1�ȓgp)���M�q�^�X!k@�<&^Y��0���;����A����1K� @k�u�ȓv�<P7��!��d�P�\,�&1�ȓ
ޞ�p�$���զ�=*�V@�ȓYp.TʶA�f��@X�#
�T��q�p��G�0�^���Q�W*���ȓ.;qm׫Z3��qK�����K7j0Hu�r7J)A� �r,0�ȓEي�ࣙ%��%!g�
�{�l�ȓ.W)`% +-�2���+����,_j��f)3h0z���I	>r�ZŇ�I�bŠ��U--��C�;O0\}�ȓ�8$�	�!oH]hc!ȴUp5�ȓxT�E����<����a��t6�؆ȓ\@�끯D�L�8��A�?���&瘈��"&����7����ȓo�rX��b�h8�|U �,���ȓ9�^������"��u� !�'v���y�IZL�c�D�F��~�fɄȓ�Hp� �ӹU��)ǌ�U����{�dPC�#�$C�)�#�J+���xbB��bBH�#��z���6�L��'l����_>c@�U��3> ͅȓ-�4l#Un�F�*�;�!�*TM���ȓM|�𰬆�b�����������ȓq��`��T��R��G�9G��� ۖY�f����9�V�܎�i�ȓ0�u��ŝUӸٙ�M��iM���ȓE_���d���t<X�.W�g�Յȓ�d�(�aE,$N�ÁB��r��}�ȓ2�Lh3b�Gj�v 1"�G^�4�ȓ}���"B��J�F��;dr��ȓOt�]I�B��YTZ��o�1(�ȓddT8��O�*Z'�Y��j_ޭ��S�? ��ㆌ�jJ�1� �����""O:h�ggSH�`�!`�"q�>��P"O<�c5�� �@�#CO�+�ʡ�"O�D G/
�W���{1.�,G)F= �"O\��o% �^xFo��4��y�"OJ�Q)ޘKF�t�7�B4d,���"O���[�/��@�M�;WP(p�"O8|SD�O�%����(CCvI��"O���a�[�!����
��2⦑!"O�<���с�V}a���1\0�d��"OҹR ��+��UB�E8:
"�V"O�����
�XD��dΪG�1"O܀a�@Z�an�6��,e��K"O�aY�_�/.AX�/Z�|N�T"OF`� ��?�,`�rϑ�Q�֭�0"OFI��M�V�� y`/5|�� �"O����L*H�(� ��zЌ�Ѡ"O�ea�F30Z�sto�H��F"O�p�m	b�Q�����,I,�r2"O�݀W�����L�6=ܠ�c"O�p�4��"?��I22ٸi��q�q"OprҤ؃B�#FX�x��@�"Op���ə�*�l�F��Fv��J�"O�@ꔆJ�+����V��rny2T"O�Z�B�mg�q�e��)[�Md"O���*��~���ӧO�o�1��"O���O
'��yS �'U����"OT�8�EC�i��0@$\KԹ)�"Od0k��ˠ(��0` [��d�V"O��xbh�uSv�2F`ϼ8�"��"O@��2�ܛF�P�/ݠxv95"O�3�I��0���HS���jp"O �IƯͻ-�I��b�+/���۲"O6Q���G"YoB,&�T��"O���w��a����7�#lؔ"O�<�B��`I��c�M�xB� �"O�=j���z�$p��,$M��"O,XJF�H�>h,�榖8lm�d"OΤ*v�ӂp�`��&�3ya*��"O��h`:>����$�*���R"Oh|�UÂ+&�v �B�	�9@��"OD�b�^�f,�� �<;z5�"O�\)�ϋ+��#�nHؼ#Q"O�ċ�o�
��P�]Ҝ�PW"O`�₋B/-�9aM�76��H�"O�ɔ�åsc��J��6����"OlMs��L~���qDm������"O`�`@��k������S"O6y`$ �77���E�q�@�j3"O�9����a�D�:I1�s$"O�9��/| �B#�H4��<r�"O 4���G� y�sslIWx�L[F"O�`�/�u�֐����ɓd"Ob6&�(@P� $�
���i�8D��k�8E�ʄ��\�4ڀY��)D� :A�>41<�H����{s�e�vN&D�l�2�
���C�'ޙ�&D����ȍ�5 +��xp�F"D��(ū�'5Ǫ�rG� �2),q�!򄓑}p�M�2cڰ#�%0D�M�C�!�d�'H� �J�%��B"��"O���4,��b텖	�"O�]�DF_�$;�d:��$����"O pC@��Y�4!���xC 0�2"O� |̡�끙I>x����М!6%�`"O��X7M�����0�t��"O�]�!Ț�xyg��ta��r`"O8��dn�nFܘ�@���pfD�S"O���-��z'�����,<�h�ٶ"Ok��!/��Ƞ���=i����"O |�/�-�X���LP�.�ԥ#v*O6<�BG�A����� �g#�T��'��@'N)]�V����K�f���Q�'h^�@b�!#f�r�'��[iB�`
�'v>Ɉt-�?I��hEO'[1���'͞��l�7:��]C��3j	x k�'���ҲϘ{�d�B Bȹb���
�'�<� ����I��<����/j=��3�'V(\�0$��Wzph���J�T�^�	
�'�$�`ņ�*R����I�X�#	�'C=�f�I�%��juT1?��h�'��˶Ȁ�s��T5/�>�	�'�j0�AD��Q�@���%Y7
��'ɰ�iv��iǺ���C3X�!�'�d�F1;�Ҙc�jӼ5��<��'38��%OOꖙ�a
�)��`s�'���i`�e�̸x�*!�^ɲ�'�HyK3�Υx�tu���p��'*��3ũ�>]i�!u�k��;�'rR��aǍ�+�^���AT6�2���'b��S1���+`r�&Zw�b���'�D9��'@v:l����"~r�!�'9&����6mKBUZW���Q��'��@����>�8Z����4��'W܁IQ،jD��rV�� �v���'�B��.���,aW�4J�yz	�'ve�H^�>�4)���5�	�'�|��P�-z��)
W�1(���P	�'Qޙp�S3��(ƫ�;T4���'�p�#@�c���a��D��\��'i��(3Ri�.8�%��T�����' ¨�%^]O���&EB�ETY��'��ī�,N�@:sJ\,K�t��'�R�jH���3�\6���[�'t��� �>/��%��
����'�l��EՈ)�&my�儮n�j��'A���۔T:LT#A�­�H:�'Bl1��N�=#�]�ʋv*(8�'�by"�HC�.���k �ԏ��,
�'vXU�Iσy�	�gK�jo&� 
�'6X�:�)�n��`����*s�]�	�'<\*��I$.نQh�D����'K�����ߊ-iv<Zu��czL�'>��@So
�z�	pd��[q&���'܍aE`��Rx,=q�"J�-u���x٪�����$�9�H���M�ȓ�Ľ���@��b6�Z�K�N���4�dP��@��k,�H�Ъ�
-h��ȓ`�${�T{�x��4�@
�Ƙ�ȓb͆X�g��"����g��Bvx���i���+�U�qʹ��[���v�����d��_ %&�=��W��|�&O�+"TqS$��r�t��ȓ=�h!�F*�0�e�Rs�|����P��D;�~�RU�ӉPP����d�A�c��q�|�#����m��f��dˡP�y˲ly�D׾F:"مȓW<>����Q �x��Gj�#��!��S�? ��H�dܤ2�v����0FC"O�DbP�J�fܐ����&��,�G"OH= ���
�I���HhS0"O��X6��)Q/X�2��͘*e(@a�"OL)�!�Y0" �SH� l�1"O�(j���	����"��DL�4"O�i82�W�Ɣe��x�"�"O�aPAE%L)�Zv��Y��Y4"O�����-l���5�/G��"O4t*�2O꼜aeC�{-��p"On�#`�Y@�P`%)m���"OJ1{�	G�>1��� ą�`"O*PE�1R^ ���
�-���I�"O�=�aۆZL��3Q�7a���k"O�D`��ܫ@��R�A1`�;�"Oʈ�"ċ^T|I��ě��Ƀ"O�L��oZ�d��T)Ʃ�'�δ�c"OTq;LT�n�Υ)��9ׄ��f"O,���K3�6՘p@F�4�X�"O��Αt<�ɤ��6��Y"OvЂ@���8k�4��%W .�\�9"O41I�e��@�P��R�ST�Q�V"O�{�0,0@fQ-P��A���M�!��!p�d��MB�qH�eҎJ�!��@�A�BT`�O��.�z䮃�_�!�d ��i����Zbp H��F	�!��p�0M��kYj�F��!���dO 	�#%��1OL���ҭY�!�$�;^���S6Dd ��Yn�!�W1 O)R2�����+!��4M!�䖸O����D";�l�I.y7!�+��Yc�#*��3��I	�!�û����F�)@�R�J�.ӌF�!��B1[`�A@%��y�(ܫW!�D��V29��'�T³h��+k!���.�x�����u`��ۨ$W!�:��=!D�^װ8cf�%h)!�d��V�R�"�*dj��!�+!�D֯RA�hC����&`���#�!����d�9I%���p��K��P�!��ֵ#x|�T��T����T��!�dQ�-TV�S�Yfwr�`�R��!�d�v6�a�G
�k�r���/�!�$�&��5�%�Ta���aI�!R!�d��Wf<@�aBP�����# !�DD�$q৫P�vx�%(��N!��X�\����� .�)@E愛T!���>��e ڻ=��+�j���!�D���9`��W�s����#�!�$t��+YH�����;q,|!�"O���+���(v���\I �#""O���m��s� թ�R�:pT�"ON���M[t�0��g�X�fA�'}�t��a��n�̨;È @��'cTܘ�nX�4�4 p%,�&#����'�FC�噺���޳F����'b���w�M�CC�J�ZXx�';��
3�M&����HмU�'p�\zf��z�,�)�HE B�
h��'�``�$�S~̘�m�6Op��'e $d��K�X�yG�P/'��z�'��K���<Rm>a�7�W�"׬a1�'�1�X5]�9�aW�D�&u��'�:=cGdȎ?�tP���:Ax>+��� �̺Ĥ�$B�L����85t��	�"O����DV7���1� ߴǤ��"Ojy˂$Z�q�f����L�Q���"O��M�"D�f1�O��=FT�q"O~�h0+
�:�˅nˎ@=��e��� ��v��E�ZC�I��ߌjެ,Rƃ�5J�qO���5gA�x�./��В��\+�~�c�O��A�N�7A��P����,����d�r�\ 3��=j6j`�̇,j.DX�hšr�D1٤�F3`����4��DGz�dZ9�?���D[�OٛF	ٵ]���2"L�!��
�JZ���=�)�S}�6�l�v�v��a�A~�������q��4�M���5;`��R�:CI�ř�eY}?Y�"ғ/���'a�)BJ<1�ѝe�P���;'%l�[��5s�	@�mL��Mcf ȕJ���&�ι��O0��;.̊�cᣂ8,}�=kt%�_�Lo�BE��1�G��w�l8S��'(J�Ăɞ���5gY�ۆ�p&꓃fg��y"̛5�Mccğ��0���OB>7�U�����jͿ[^���[	d����?a���=�I!+��c�h��?e�H�� I�|�<is�ibR6�%��κ��!;pv��i�O�
��(U�[�I�c1d�kܴư<A��0�Y󀏙A�n�k.���$S�JT�h2P������@��OĚ�Gx�$��H�R���4�Zp:uK�C���	0E�n���6c�
���Y?�Sw��ؘ'��7�Ht�F̪5J��_RP@r���O�pI��O���$��Y�x�	L}�	ϫ<�t���1E�	�BA����O������}��oc�p�!�i*�fLӂb����dʓw(@�-��t+��f��:J}�T�kY�R����?����?���?��?�O�b�$�*D���G�d���+��NV����VV�E�2�}�,����-�V<����(kJR�+r��uZ�,t��;(F|�µ�K"����	�r:��|Ӷx5��v��x6灳s|d0sRc�i�	� ��j�S�d+��K�=�4�a7%	�p6�������}�(��0l)�J�#J���7��n?aw�i��W�|c�d���)����mӅ��B�ژȥ R�R�qON��8`�v�iv��.��G �7� ({�O�����^�V��3F�6xV��x���ϸA�LaE(_�YD7M�+x",A	go7�l̙"��4Ɉ �s��o^YB���R�wr�'(�7-�ON�'2K��+r��6Ե�&c[�H�T� ��'s�O?am�\"���D�@��`�)�)���d�ۦ���4�M���Z'4��p�Ǯ�JG�XD?I�%&��f�'�"V>�b������˦�x��P�K�1m�����y�$��̭*ׇ�0�h�`�N|,�	�S/�?9�O������\0��;\~Y�pg�"\hApP�iS$)!"�486,jP�ŷ4�a���"^b?�k}��qB��ol�1ugE2hq�6���tR�'T�6-�O�#~n)`ml��7H��	�W�A�Z��	�� ����ؖ'���)ܿ K��h��ܝd�]+�%�}AQ��
ߴ/N��|"�O���J�V�P�(L�J�C�&�''��%���	�m$ p   �   G   Ĵ���	��Z�Jv��&�Ȱs��G}"�ײK*<ac�ʄ��	�*t�Xx�ae���$E#vw�mɶo�8c�i���.�xn�2�M���i��5�IU�A	�A��.����ڱˇ�Z�@�@'|}�#<��Op�r}��LƮO4�E��B� �\)	�X��{"�ӗD��u��<�D��k]b8��Y}R��ԁ�C��v��u]�s�t��F]��a������y�c@�HZڴ�;*��9O�E�AW`6x��d��h�d}���<DL,�J'�����վt�= �,��I�?lR)����5���B�4�K�b��O�Z���h���'@ZtGx�t��6�Z������#�@zF��&���	�Y��H���� i��0ʆ4t:̭1c�.4!��Њ�ě>�O.y+�O��x6���(�%\ K�m�Ɣ>�V�4y��➜�`c�?g7Pl�0��i��y�5�tӒm ���\2�O0��An��5T�S@�&�}�@I�;l��O�Qj��̹��dK�d��k�K��7ԥ���u��	5��HR�$q��q���=�(I����g�L���d���O`���k;���MɿDy|!Z��(���<��0;4NO<|8`�X�E�ޜ��&�'m�M��O$-���D�$�ē6��� ht�d�� Y�Y��˵pZ��(}��O�����>��'����G%
;�B	'<X��B�Z�|��'�I��� m�'6,�O(�9�* /��c��6�,Q��W��J�ɫP6�L���J��,��ұk�xE�n:D�K1�   ��F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# �P   
  ^  �  t  e'  H/  �5  �;  )B  mH  �N  U  K[  �a  �g  n  Yt  �z  J�   `� u�	����Zv)C�'ll\�0�Ez+⟈m�(w��I�J���D<c���(�6ta�!gE�r�4aE+
�"t���¶c���ů��debͬ;q�E��'8,M���in�h�A0�����9e�$�`���B�H��!	1/.QqUGȱ�,�{Ŀ�:@�E����dAA�����|�RP@���|}[4B��p�~�Aa'�O� pg:�E�P�٦Y:QO_П�I�����(�CͲa����GC_"=>bի5�W���� �
�	lyR�'6���g�'��'�"�%��>�z���C�P2��'<R[�|��_y�D��M�'~�_9{+������zfeI�.ӏz��0O�a�V3Q��C�z��x�Z��F|�c��A�<�M�<,���@LT�d/	�#�ϟ��I����I؟��	����IG��3�̀c�D�u����Fo�+vm1��'�X6-Ҧ�۴U���'7^6��Ѧ�۴ ����'W���S~|�)+��˼N�`-K6�"�?Y ��2nP��ht�<S'��	�t�ģ%��B� seڦ`ٴ{�V�OT�IZ�O(}H�nD7n���bڙF�0=rS.B�on/k0�`j��ў7m
T���F�n0�ݺ�$F`7��¦]��4|�&�
�d�g�\�B��	]�5�g��0��U�c��/��&�aӾ�mZ�s�������|X�n���3a�� �p�*k�zՁa�� �ɇ�P�
G����F�>6���)ܴ!�|]SuLw:>�(V�N>h7$Tx7ՒL,�!x	@8o\.hIf
�H<��e��< g��-�|<+���)%Q����)NW*S��5*\��t��"O!(��"��ğ�%���ƻ?���E��+��x���H�Z�9Q� D����,'� =CG��W��bh<D�hE�U,vh�z�Ʌi"�([A
/D�LP �A��#��Yg�L㰫.D���/B)L�0����K����D$'D��
��T��e3F�
)(~��'7�#K��G�� Vrf��BL 1:D9��$ń�y�D߸}��ā�(�t��R'�y"���>?�ڔ ��#����1�[��y��;�%	��W����K��y��_P��A��i� �:��@a��y�s�y�B��,T8��U	�?ɀ�Ox������*'��Tk�س��=Yp���D>D��+�!Tx�x�k�A��D�6D�<f���V�D�G�҂[�� �bI2D�8�aoȬP�h,3D	۔5 �M�0#3D��KG��:�Q���C�`yH�0D��� )̽�Q�>fb�hrE�<� M�f8��qT�g��{�"�%���������yBH��i�����O�l�iB���&�yB�%Jڵ�DJ�:c4���Z�yb+��P� ��ôwl�I�#���y�i	4p�*l��N�j.��C������<�Tk^j/���'_RJ�7Tx�$��'ҬTΐ����.D���'�-I%�'��>�4����}�Np�I���7
�<�p�Ǣ�7f��5p�l<O>a��$��!����t��S��F�T3uWΘ���܁t���:\Ř嚌��̩N���'zB�'_*Y3�a^A�pQ�jL�6�6҅]���	a�S�O�Qr���\zΙ��aS�Y�iZ�h����Y�t2� L'm~�ᵡ
�?�+O.mC�b�Ǧ���ş��OE�-B��'$��P�Xm��]h�S�v�|�hA�'�.����D	��2��e��)TW���'��I�[�,e`6��wo�t�%�H$����*�\�eL� �m�X��,s�C�ħ i��&)]w�����J��P�'�Z98��?QH~����j$$8I�r�,Jp
��$K����?A�{����AG�%���_`]I��q�'|
�}J�I�9g��tQ��ƲNr�rvaЯ�M��?1�T����"���?Q���?����y�ё �
��̈0ϲMW����p��+��\AO��G�:YQ���5�ÉK=�MiW�I.$h�d�@�C�T�'%�B�V��@�?j��� ?� �'���e�A�J@VNGW��!��O��5��T��i��|�I� ˠ�h�٥J �%Wm1d�d�<���6
���� %6��D��lUy$��|�����$��L����֊�sE���Wj�29od w;O����P�m��`�D�׊�&�p�F��73�0�Op��a�M��h6�E�Z((g�=J�!���I���R�L�8s���%|�@��'V!�$��q� E[V%�&jZ ���յ^d!���]��+��k����W���dX�'N*6�,�$�=���-?��d�# uT��SV��`���H�L���h͊4� ����Z�.=� �$!�$*F@CB��nC$m)@��&����'4��� �F]c��(%�8��Y�Aכ(J��d+�?&%��!�O]�5Y�(��䚀'�kv�Z`m���t�2��>@�uQ�㒻���(֫�ş�Iџ���ȟP$?��<�N7J��	9��	��� �X[��H���P8��&w���w`9$���By�W��7M�O$���|b����?� >@,eR@�:㎜�vd!�?��f�!��HDl!�1��L$',���ļ?a�O�N�s�zbF� �Ja��t�O@X��Z�� M�b��D �X3ЩAv��$>]J�κYl�����Y�p�[�a ?!�E럘�IG�̧c�.\�온�۶�-&����r��������y�*d#��aGΨ��0�%��>�7D�)�XD�8K>�H�+�ަ9����I.r	�]*ea�֟������߼cT"N_뼁�2��'�fX�' Hur��v�3#�Y�
J�Hgd��|b �xR����I���C�T�b*�@�0���H��F�!�&(H����������!�P.��3�{���IK~�'��?������?y�����d%F0|�����zn�B�'�VI{�ǃ
�.����YhtX�.O�EDz�O�rY����+<+��9�g��U�ė�TJ����N�iz����O���O���O���'�P(����R�<�k�ʊ�@w�(�t���v��g)ޡ�p>�P9"6"�n\�5���
�
�!X�]�#�9r�5S�
2,��/Z�Q��@� �G"O�]��[��oڦ�'\R�z�V�$�<�����'\��k�D��Htx�Q�k�P���S�|��'���Ru
ǌU~�R)��
���H>qŸi��V� ��A���d�O�-��-${���(r&@c1�a�e.�O���L�^g��O��ӰK�,V�=hU�O�l���
W��E��`��`}چ�']�0��+Z,4�Xzm�,F)�t`dK�x�"� ƭ�+C�q���3u)^pE}"R��?��?Y��|T�L�B�T0X��� �:vN��I/Od��"�)�'����u�.�c�Ɲ,�ԸSN;�OJ�	�!���i��?k�0K�K�&X��'�d�O�����9OZ杚zW6Ѱ暬B��7��E�@������
$F�=|��CO�k���ȓ$�T�١-�>4F�A:�O�I��<�ȓd&���#^�y��A��0����ȓ0fPS�� O��	'�<��a�ȓlQt��#ե0cL1�E*Y����I'~��"<E�$教 A�Չ��H�r O��!�����CgN�.��1���!��	\`ś ž:�����O�|�!�DA�%��\s��D$E�`|���߮N�!��K�F[�ᣢ˛��
@���|!���}�.�3c���S���iE��Rs�I�	e���$�^���GI�GW�D�`��`!�䜒A���D�ξNR�T��]�Q!!�A�o����1*��Y4Pd0v/��R!��;M����6̈M��m؝Z]!�d
�H��Ԑ���+�>����ǻSK�}2#�~b��0	?�Zs"�
Q�P	��"�y�n��W�����	ʘN1K�(}���ȓ!���BDj���~2��F�:��ȓGfTc��Ļ>�
X��댛qf0�ȓFQ`�b����G@��3������K����A��YC C�-�d�G{�!����TP�D%t���`�f�Ot�- "O��R
Ui�����:��p+1"O�Y�m]�)eB�(v�ۀK��8�V"O�yt�V8S<�&HU�We�x"O�0�͖s��u3��=cD�Q�"O0����\$]�oˌ�8E���'..����S�/���§Cɓ{h=A��'u�ą�k@T�+��BX�س�#����ȓ�4���Q�f� Z�<t����6�"qC� �;lW�q�S��bt���ȓ{n	�B]�,sz����/o	��Vy�M+�
`6QAqo�#�(	�'�|"��$�鐠uwxH	�M
!E��݄�S�? �}*Tk�
A���ã�nG��J�"O\�PDeݘW�ƀ�T�L��p"O�	P��Z��`��*ڣ|���"O2�K�,�Yas	�)$ش�W�'�&I�'�z��1��z�lыī��v4�I��'����+��<����2�Sb�d���'@���[ aZ� #J�og�a �'�~�x`�P"}�rS�V�l� �'�4��6�A,�p��
n;��h�'�.�(�#UB���a`�hq��$4Q?1
�FP�&�� �:\2DI� $D���K�,�q�!��EJ|�wH/D�8��j)��=*Ŋ����!�*D�!�C.m��`s�F�%�T�$+-D�ٰ�Y��9�Rh���B9D���$CW7R?�����N��� :O����)�']Ԝ��b��3~RCQEϊ�i��'~Ԅ�u$�xz$��g�����
�'Ťp�B�YT�s'�¼�lLC�'?P	���N'b	�䙲�~�
�'���Q66�8�����/Vb�<)UI0�La��`�1iaz�(2��dyr��<�p>٠�[0
�8\[��M�!���d�<��&�3�:C@
�,�B<�`�W�<��һ<V�H"6�U�dl����W_�<as��1�rI�qNW<,�����q�<��ː,
�q�6��65��<�0/�kx��0���� ��b��	~D�(T,�9+�>�x��4T�\�U,��
�R���(fT�z�"OY��R�vBR]cM�B}�c"OޕpӦV<d7\EBBU6&�s0"OB��C�T�7,�b�����y��"O� ��̙9��@�t C�X�M��D�ޢ~����p��
"�ͥAc~1T�Vk�<��.��&Z�����g�f��ġ�]�<Q�O�>0}ոr!�%-P�D�Bd�X�<�q#G�(Լ���@H(� ,1��P�<Q��H����N/d��uy$���nRB�	�X���Z�+�]T�hA�W�>Q6��*F�"~ڃ�
b�p���BH�E�n�����ybcY��� �T�˜=!ġ��m[$�y�%K��pU���18T���ϫ�y�+�R�zx�&�>W�H8 FJ���y
q^����I�Z�q#���yr%G$b�ƥ�U'U���v�ϑ���+b�|�O�$'D�����7x@pE�%!� �y"J�h*<�X���<�p	�EF���y���2�\�yeK+2Y��J���yRH�+hO�9�G�+)ܩJ5�[��y��%l-,�z H�����`�f©��>�S�V?I7���;���@�Vo.X�� �g�<����i�*iUM�u!�qT��i�<	�!̌N$\��M�;#���EbPi�<����B�����:U2d 4*�p�<!r� ���B� �K��t��oSo�<1�E�t��c�֐A�)�6��e�'ir����#Ba�� '�]���ɸr�Z� j!�Ď�!n� W��X��4Y,ͫ=Q!���(
�Bird��`[a�cD�=G1!���!p.��k�윿@�t���?jG!�D
qbp��|�r�
T̄T!�$��8�BF�$c�zD�3�U�>��aܒ�O?�����K��u$؞|�0ѻt�Pv�<���F��U�� 'ݦ�J/�s�<� <|�Pm�4kF~P���Ϥ��c"O�t8�L^*t��f�8�%!�"O��0!O�R�4����B)*�a�"O� ��-Q*cV��q�lE�W���BsZ��b�(&�OL���_�l�&�IG��AB��"O��i#bT
7x�p��"+V�(a"Oh���H6Rն��G��3!5st"O�u;fo�/�e��{a6�Z�!�$ŜH+����Jü5� r��R��}�a�,�~�<NR�#A癦D�@m
�L���y���7�|��3j�	��Q�L�y2hP�k��m6_N�`"���ybgƸ\22D�%�J�~�`��S�y�N�u�V��������b��K��yb58�|�c�;��k��6�hO�%z��;R��`�'~O��2�cժ:�C�I�Q���0�����:���NՋ<�zC�I�Ǿ���"�9��H"��-�,B�.��x���]�+a�ո2,׀Q"B�	$NM��J�Sp��s��S/6e@C�'S����Aс�B%��;k*6����"~:�P:F������5^���䣒�yr���  �\�E�]�M�Ĝ:�㜀�y"]=%��qKsMڑA��	h�O�=�y⍑�	h
xiЪE�1�������6�y���x�21���ڬ2)�b�"܏�y"A;״�k!��p�{sL����D�;#��|�(B���c���T9z���y�BH}քlc����S�5n���y�N�W\�UȆ�u�8yU��y�M�y��HY b�	)���Ai�!�y2k̉T������ɍ#�9rR�����>��hNP?I ��^u��E�&��(�`P�<���R�9�AXC�����')��G�!򄜆2(jq�יW\��6�I�C!�?wRQ1!+W3..У��� !�$��� 4�|��]8׌T�,�!�$ ڶ�� -�d���D�ў�q�9�'Z���ZQ��49J�Q�H�W�L,�ȓc�����F�?��I�%/4 	v�ȓ}�p�T�Ŋ��@ֶV��r"O���"
*Hcj��#-�|�13V"O
 �Ԇ҇Ue�����!F�>���"O��2Ɖ:L��BG (>VA���'�buZ����kF]�b�q"���aʢ\s��ȓ5D��skH��v4qa��I�6��^��ۑA�9j�nmK6I��h����݂�f�.�x�1dF)䶡���
M�F�99P�I���U,!�t���c��Q�����h��d��@�ht�'�\P��|��@����HA�M���ȓzV�	z��_`���G�ӄ)�ȇȓ�X��-�B�D5��ψ�bz�ȓS�H1���?��ѣ	PT�Ʉ���Ig��3�(�j�k��sJ\��I,���I�*!
��"N! �69Re̚P�C䉂j*|�׍؉-��K��C'�C�I:���*ÅۯeyxLpnA��B�		oV�<9��)����'P��C��9H�E���	�K*�<���q�C�;5��5f��P:��x&(�2�
�=��M�Oa���Ώ�!y�L0��=��	��'j�s�ׄhC2P9č�
;��X��'j ��m��Q�ѩ"���2��)��� .�X5��+b�ɂ'�&1���"O�Y��?m����t�����V"O����Núj� ,(�Շ	����B�'�QP���ӻ9����B),"������ym֙�ȓt�p�#��Te���#�/ܲe��o�(y[�i	�u�����ݔb2��ȓ>M�U�s�@<��ݵX��ȓb�.,XD�Oi6*�r�ޱ>#Z%�ȓC�hջ��K���,����'Z�A@�b�<�XS�S��p�rː�[��؇�@�J0S�f��N@�m��+�	FJd�����'d�*?�X�n�C���|x��2�[=;����k�=k+���#�֡���O$�R�KR	
??PHH��ɀ@���	�p���)d��? y����
��H�B�I�26�[B,�y�P���dփE��B䉄^���yP�£R��� 	V/Dl���N�'���B�LjhdD��!�d�+�ґ�䅇1&�r��I�Au!�Ē�eN:(�SO�=0��lT+g��=a��M�OL��;3�Ԓ$�������4&t��'i���V2��[�@�>�*X��'�(�[SH�27�
�P�b�� a(&D�|xb�ݜ-Ĉm��C�EK~9Ӗ"D���,و!��[�!��l�^1 ,?D��	7dB�55���P���`���Oة���)�	��	#n��M5 �aGJ��/��y�'R �I�h� �Ѕ�F �3�Θ��'i6-�'�1'�b�xC���)�r��'.��Ͻ{�X�wH����H��'d�!b$n��cY�|W�ƣ���#�'�<B�$H#T�-CN$&5�6�'��c���I��T���B9������J�S&,&pے�7o�mb!����DxGmB���������@�f�ꑮZ� �i>��-ߴ<n"08�W�Zv2P�K9�k�ZA�u��5'�e;E��h��lV$x�0g���1��̈O����'$��+I|@��F�cY2��UB�9��v���QL�/>$�#�����0o2�O�q�'|�L(W�͌g�X�XVπ�R�FL�,O�%��@��m)��E񟐖OC<��D�O�R�RHR鉡Ϛ���9�Љ\ q�%_�"�rh�/��*�aԧ�)2�#:�*��K$'z��5枖r5��	9EMn��Ŗ1@.,� �O?���H��3�H�b�L+�C2�r�!�O���7?%?)�'��dd�2:8A�EeTC���h�'���x�� �u��T�њA�B�����W�On��󦁴�ZDX�M���k��C��'�J�:̌zB���'���'�֝ӟ�����'1r��jV+��;Q�.-���k�O��$�C�� u�P��O��bjU��b���'�&�R��% �3_ψ�D�`��ٲ|l�3F(T���$Bkr���gהwD$�'���b���?�����'-�I�'��dJ�ɍf}�@
�b��!�$���E��j&}���P��?z�!�G����'!�4N�<3���YKs�{���ل�ƞ���b���0��ٟ�[w���'l�iٹ ����T���C��ș
(��&�d�pz7(� TdD�2F�F�'9V-iPC�3v+P��G�u粨0��ő'b$���Qg<�%��7�"?)��`���ֶo�f����y�0����ğ<E{������B/˔�8`S �+��C�I>M=8��H�&W��9�����M��˓re���'��O�iq�~z���2��z�冄S���CE�x�<1$�G��LS�e��cU[�<9���������>h%ڡ�OW�<9�bW�%Ȱ�b�ͅ: ���i#��h�<A��N+)G(0B��bN�)���c�<�s�]8H�B���v4HEcщ�_���LExJ?yC��4U$���A�~�qs&.3D�(p$N	����/@�,�����5D���ॖ�:����.�5�8H��.D�� ��r׃¸R��D�K]�!44؋"O��V
�*��ph�H�>C�-��"O�pC*�,� \Rb�C�>Njd3#���O��}�s}n����v�@i�! NFhI�ȓM�J��EH��C�(��������ȓ#xh����<4u 	tMƄT�rC�I�%�����O�E�c�@�vX�C�Ʉ6Y����/�4��	���^�RvB�	&P�x:���^�K�}��2�'��`�	��/����%X�3��!D`�l��%��g��T�c$��Q�� �@�i����ȓGB�����TLj�\ �F�]�$y�ȓ9Gn���L�f2b}+��B�g=ṙȓ�6���U.���0R|8Eb���%~V��?��O�~"���'b��PJ�)uװ�c�n�N�(��?Q�n�{f�ZaI�H���G���S������K3����p
�c��#>�R��A�8��a�Z�fr��Z-���Y�F0B��*���С��I�0+����Olc>m9r�ޒr�xhF�]�ob�p�	�<���0>��:7>�5AqGͽe:�"T�Gx�4�+O��8vg-bt�`�ȍE�>�[���I��M������?��O2my���2���PQh�o�b I3�'~ў+B�sr$�w��z�h*�	�=4�Oc?����O�i�6�{֏˗Dt^����3?i��OL��@�>��y���6(}���ǡ���\�:�CR��|������rI�ꗯ }):�i@>X�T@�K6|)�<�w!Q5��{J����'��>��$9Eb�	�S���KP���[d�P�C�9}%}��\���I���ɇ�mk�@��n��5�%"_.`��N���Z#��Z�&.�&��qǕs���Sfܕ�?قN�V���C�D�W��s���Ņ�l8\}���u�T�X��Н��$���*v�?��4���O�dKc��� ��M��~DZ����|��`��'L,�[Ǉ_�*uN��A	�=P�ҴL�z��Rd>�	�x^�>U�Ǆ��(�# �O�L�+�k�O�	�'~�xZ�O�s���G䷟h�l�"��0@�z����W�O�	�z�E�7�X-l��L1�j�g"��ȓ\���4��u��f�.�n�(&�
����Z��4n���:�m��'��!1ǣ�9ͤ��'��'\�Ix�O�
 B �+���hf�W,}e��[�'�����Í0%fZ����%J$��'�lxaZ(nu�S��8s�le�
�'z�ʀfĬQDZA{Ҡ�lQ�	�'�b̺UM:-�9h�j+(�
	�'Y�0�w/ͦj�a1W#��S{�t��!P�"Gm�:x8����?*F�|�ȓD�|�/ 0e�xe*�e�&���ȓz[Թ��jI3(<LZ���Wr�m�ȓw�T�c�B�a�� �O��Mo��+L(E���(�� �/�,�̄�:5VQ�u��'aޜc���H(���\�8ժsN���sd�%;�~�?�D�ݮ ��Q����7�5�Ʃ��@`��� J T�|���,@xa��a����N����%x(L��*$Z�2����:k� 1A�/T�JB婐>@I�L1�������0Ŕ�3.����	>�� �+Gd�[0�ǚ&�l00��T>�T]�9��%(<��!O�S@�X բ�>�!�ɇuZ2e�R�X�j�����E�q�!�$ȧ�Bqxɀ��\��#���!��S�uLl��5%��l݋��1�!��K[��nOI�^�D�p��&B�I���Xy�Y6���*p C�	�o�J�A�-�~��#8�$C�ɼ~�*\��Ǒ�V	�a	B��C�	�G6tAR��)}�~�H�̋�B�I�O`����ԼA�Ś��� 3�
B�I�E&��C@����yr�ם׺B�I :�>P��ɤ�iۆ��s^��$O�j֢-"�L��j^�8��?7!�� ��d"՞(O�4[�<az�XQ"O`�f��Vj�����:v��`#f"O�܃1'˶#� �Gmӛ;n��	"OH3�/ ��3�#_T��E"O!22�L'���s*�g���p1"O0$"Q���@���#	ݻQ���"O�p:TMV�D�dd�Ʀ�"xQA�"O�x�n�*WF`a�!,2XR	�"Ox�CF��[-��0+C&-��s"O�LJ7��;�ΘW*P�P�8���"O6	�4�W)�@qR@F"28�b"O�	f$��vt�#��E쬡�"O��QV�s%�u��7o6bUA�"OҴ�T� �[Sj�0�%9hz�B�"O�0HG`ʹB ��a�%�m#2"OD����R:�t�Ee�9tz��@"O�,"�Y)��0*@? ��"O���E���Ȱ���+ ���"O�A��?tT4��ֶ5Z�"V"O���u$��Ґ��$�X�"O����E�s��0x �&dP��b"O�T�6�������G�"O�ma�CT���c\%>)nX�"O��Jd�!Z0�Ǣ�"�i�P"O|��3;l��u������F"Of�q�S*]�!��
�F��a"O���bOZ?�R���Y����"Ov�s"%ֿp� ���@X5�"OF�k��±;�<�����|:�<�"O���5!O�e�x\ۃ�^{~ތy"OL�!����k�@���C�UI�p�p"O��V�-~b%QlK� 4F��6"O �3������$�6!"�2�"O�����z��T�0���aH�,�yr�Ȥ�L����~R�����6�yrB?��t�*�1{�ά��G̗�y�$�.bl��o� ~�:�H���yO��4`0���t�+�((�y���i�$9�mS)&�1R���y򥜿t^��0��Z��1[Шǋ�yR����;1�N6UCN�:L�-�yRF�� ƸP:��?�-��k>�y2ʍ%����*P4|ܨ0�[�y"M57�8��D�yW������y2M�3-/޹��+��e�|���C&�y�,&�!�����%�|���M3�y�!q�5�'��I�,scJ�2�y�˛y��%C	�v��$�X��y͔�	(�����-w�d��=�y���6��H���)?��1A���y��:�]��g�0�4�z@eא�yRl
�8�1����&��ih�k���y2�m�H���]�x@��nU��y�K�;h��=P���l&Ҝ;�@�&�y�
�~(",`�Ɂ?z��hAbOX�yR�[X�̬�Rb� mK�i�#C(�y��U�3y����]�_iDt:6팙�y�G<��吤��;~��T̊�y«ͦZ,֥�Q�R3���t"��yb쐨7�x(vBޯ{�V�3�NW��y��`�e��F_IF�*$F��y�,ЎE���"C Vv�y� �G��y�	�aYy�tG�4&b!�'i��yra׼6��@�S&^�1�V��y
� b,��b\�I�PC�J�v�"H9�"O���&�_�2�a�a��r�"O��*�O���bd��T���T"O�$a���/	�bc�CI~��]2�"Oд9%I�p��y�X�r�P0!"O�y�'�؎*R�T ��)�J�A1"O����Ef^B%BB�Ύ���h$"O��r�T�)�`)��k�~` 3"O��q�L�6@�0� ���r�"4p�"OnMꃋ\75�0T���æq����b"OP�1UB4~��2�n̓K��Xrp"O�,����Xr���ĘX��2e"O~�)4�E��Z銅MB�,{l��D"O����e;� kK�YM*%c"O��� �8��Tc��4!�x"OX傅��,�R2w�/$,����"O
�dMFȪW �&��b"O�X��\jb�x`���i�P��"Ot<`�e!zv����9i�:��!"Ob��G�K8�,1����D?��	%"O\̛�	�18�04C&����J�"O����޹;�1�Uf�9j<(��"O��z� Üt��3DC��h��"�"O�0@0�O05��J�! yHmJ�"O�]�'�5��h3%���GX4dX�"O����
6�9r�Z<�Z�"OҜ	'�I�pf�C�lR�S'h4"O����ѝ%آhˁ�:��!��"O�y`5��TX:��#",�uzf"O�]���X�x�p�ס��d�Y"O� ��J
J�~������0(�"Op��J+'��C ݪ��!�"O�]�WmC�`�ΈwN��?��B"O�xaUjÍbǔ�P�X�(��5�"O$%��5S�$`%	�u����"OH�Q�JZ>�|-�R/V?^���;p"ON���
�@�J(IVW)�h�P@"O<�+V�Սm�|�E�G'>1���"O�����6�>�"2n݇!|���"O~i�7@W��VJN��up���G"O�arw�T�u��Z�o�"s\�a�"O`P˷��v�24����k<|2"O��%��=F�����VJ��!"O��D�n	�+H
DJ�QX�"O�3#�ٴ@��PHG�A���"O~A��	D�=��1#�-#M7ڐ2"OT<���,c�̅s�劃���B"O2	1R�Tq��Q�Αk�|�J�"O.�G ��K��8CnE�~�z�
"O���B�B�I2aؠ*�f����"O1 tY��m�5H�!�T0��"O��`�iL/TE!���Q�"O�YĪ��BC�5�s��8�M;G"Oj��qe��`vo݁-~���"O$j� qА�!��6@��"�"O��1�?G�ɘ��$X;��g"O^���|�<��D/F0'>LJ�"O<�aA��QT�B��&��Ӕ"Opx�i�3�vX2����i&��hu"O�aؓ@�����
�E\��"O+b�,h.Y��@�{g�k��Y�<�� Y+X���g�=c"�3m�n�<����b�0 �pj�98" ��Ij�<3"�=y�|�:R�յQ�����)�h�<� `T8��	0�T]�c��:�"��"O2�"�/��� \Y��˘N�9'"Oެ���A4�ہ]+b"O֤r�B��Cg�y���P�Yx�"OpQ1H@�y��*ԲW4�J�"Oq�"���^]r�t	X�6/���U"O����̢U�&�QcC�rd)�"Oht�<�8���3�>�:e�r�<��)\e[�Aņ$�Ƞb��]w�<I�`��qX�`�$�B"L�[� �w�<���#HqF�����la�6 �H�<����#I����q`�c��e�w#VC�<�/��7���Aǅ�K�.h"r��@�<i�L.\��cS���R+����Y|�<i�[$&*.h�Re�;u�.a"��v�<�����b�Ջ,��g�w�<1W+��/�QR��	p��ܹ5�s�<��
QE�tГ� B�� �%�I�<I�ؘ^��E���c	2�KFz�<Y�AR$�U9��C�
"�-E�n�<��JA�y���#  s��t�R�Pg�<qw��9CP�"�X�L�6T�v�[g�<9�=?��X<:Px;��WL�<� �T���G�l	u�N�f�C�ɯ^vtP�n
7,�Jx2�
�Y�B�I��Dxd�V *�N
F���K!ZB䉰�z�ٖ�+Y�Ѫ�3BB䉭hhA��J6D>E��o�b��B䉦C>�I���M�r��Ƈ}��B�I!y�\@�g+�/ Y>5)���}rpC�ɯ���Ǡ,I�2���Y�C�5a>�-�0.�mW����`M�OМC�pR2h�v�C�a$����O�1�DB��8[�����ʠ'�^у��j�>B�ɥ!�D�:S�Q�N�F��WF�)y:B�I1��uqP�ƠIy���§{C�C�ɨ:������f��<8w� 5 }�C�I7�Q��X	;��m3%�B�O:B�ɒZH]��b�w��]��ͯ+� B�	 ��p�gM�|�5*4,�xmXB�"^4μg��K��S5�Le�$B�@�2� CI� ʨ�!C�
�{��C�ɘ=D�-s�E?X|�KЂ�<�C�I�<�8��$E̬sf�)	�]/B�I02� �7΄�oP���I	P�B�I���5Iֹp��S��E�^�B�I�=��(V��J��0�Tb �=�(B䉪f�=��H� ��L�ҧ����B�I+py�It�̯'",S�ʼ�B�	/��p�PG �04�l"v���o��C��("�I�Bb�/X�!�h>P�C�I*i=��ڶ �; XҜ�a-�h��B�ɤ6lМ��m��_�9��6k6ZB�I:T��x�Wş�v2��d��#e� B�Ʉ[~<XJ�o�:I*��@�!Y1>�B��*Ap���K���+C"O��!��[�{��PP�K4�~�hb���`1qO�40�JT�8�B�2����R����|���T�|�p��q�R��y�j� ��Dic�l�^\c����y2j�8x�-٥���[������y"�K��Q��MVQ(��a�M�
�y­�(]�@8�v���Gj8����y�I��v$*�I��z��D�alB�yE�as���J^P��p#H%�y
� �!b������P)�miz�1�"OJ:3���y�͕ZJ�(V"Or��UHA	U�2�c�o�?��`��"O~��6��	��	�3�F>�Vt��"O�(�c&�6Q��79�J80!"O��R�	�2�<0��YIeL r�"O�4�"$	�w��|Z���,��"O��:4�Р��02w㊶6���"O$<�j�i��{҂�K���2�"O$��AN@=��pث]�VБ�"Op����m�2��ݷO��R6"O���L�� DyvK�/��9�6"OR(@HQ?s��!pkK�G�DI�"O��Ł_�y@VlC0%��
�j� "O��˱��l,n|�Ν�U$��r"O�i�3�S 4�haM�wd�H�e"O�������$E.����"~I��"O�q�ѫӦZX}+��կ,�="'"O>���*VlTѵ(�*Ď2q"O4��%�J�Q��)B(�+�(���"O��7A�Ԕct!ʴ;ƌ��"O���!���V���ᙫ$L+�"O��t�B�r��t:���A3��"O�)�m�p.p�s7��1:`��"O"	8� ՝�\8�i�"�ݑ`"Oڱ[1�ݚm��$���:���ؤ"OP$�J
�2ha��+W+p@y�"O$�b���3������� ~ �L��"O�4����3j����jZ1��"O(��%(�	"j�a$�0rTX�"O�6��� �����KH�N�Y""OnЂvaٱ&\�s�S��L�"ON��4�Ӑs=ԁ�֌Ro,��"O��p� ��U�#ħ+�-��"Ol���4�f��!D'|j��"O���Z�
���ŧK4Ru���P"O�{#��i�L��t��`�5!2"O0�۶
�"[6�bEW�RH�b�"O���ąʁfV`X�����I �8P"O����B��L�q >{��@c3"O�5*2&�1)�|)�kۉ@�^���"OX��c鏤?JH��`�ɟʥ�""O\�1�FձMmfT#�+I�w�1�"O~h�s�@�:����^X{6=�2"O��h���!�ub7d�*[ot2"OԠ{dē
�ؑCq�{c�%0�"O qRAGQ�Q��(�HAR̘��"OP$@��Ƽ������A�[��E�b"O��21����Rsh]?l{  @f"Oh�K0F�>.]na�b�I����9e"Ol{�ρ�X� !��=T(r�"O֍�m�\�V! u�́DN-Qp"O��P�k_�o�����"��ao��B�"O.��fb�ԑ�5�H�AW��p�"O�5��.�s��4�����"O� SE�#l��x{���l��q&"O�ke�%]d=i��ĸL��d�v"O�,���G;MaxX�'ł`��Hj"O<��,A�5J�<X��:��q"O��8d�Z<��ԣ1�_8vͣ"O�K��Ķ��x�׸I�E#R"O��ǂ�w���r��H����"O��Q�Ŕ�s�"CϜ�J�"O�\��ƺ^�Qx��K�Z� K�"O� v9r ���,��ѡ%��n#6��"O�i�t-�#+g���~q��Q"O���Fk@�(���nKRh�9�"O���q�!4r��B��F�TKl�q�"O�m� �п1a\г��
�8Sfz�"OX$sc�[Îx��+��z�����y2'\2��y���O��\�G���y"�3H�Ʌ�N"wl�'���y �@��xY#����H�ߏ�y�a�
?�bu����G�B�g�'�yB,��>��)��l�p5D��/H:�y���1�6@���$6�X��7
��y"� ��1�R ˣ&��i׌�ybE	z�
�ZB#�*(�p๥��	�yҤW�U}���D�ҁO/r�Q�Y�yB��?wh��Ԁ1�������y�d�2����um�d�G _;�yb�ٳN؃B�Ҵ�v=Hfhԣ�y"�ۜQ%� �Y�-�9� ӌ�yroɎF|�1 MG�"�EAr�3�y«�*Ya��D�o�$�;�
\��y��ǅhܮ���.��i�\A� ��yr���I�2�6Ĩ�.��' ���y�l�g�L��qj-*�\�!ǃD0�y򆘙J<���F^���i����y����L^�d��\�����ŵ�y2*R
Gk��0'� $E��O�yBȗw���3C�'p���"`F��y�)W����/�o�dL%晫�y2�*��P!ϿWj����в�y"	�
{|���*����E����y"��4aMv�3�H� 
�p����y�������چ-�&i �C� �y"N� qtL�{���:�L�y�L\*HX��� 4;��E�
Z�y��NQz�a����,�I�V��y �3Z���F��^+N�2��O�yGA@݆�3o�4*� �,ź�y����Q�1`HQ[�D����s�<1�cWs�z,�f���M	��c�<y�iU�$~�#���7"�a*�Y}�<�!�ۣ!�� �B^�o����@f�v�<���.
�\
���0��T����\�<I4���X!�a�VGM�B�
�Z�<Q�������r���Z����%�X�<��-�6J��$r��
`�6,j�iXN�<AF�[�B�䴘l�pyv�K��PT�<�sL&�BH����'��x��$D�X�E����Q��� &6�yAo$D�d:&�M�������M����$�!D�P���\�=vM�"C�&l�1#!D�Q�ȉ0T���T�H���[�o-D�+r��<bވ� ��Q2 �( �a+D��b6GުT��d����+na$��u(>D��sI	�0N+���-s�H�Q �;D�<+T%3��Ik���6�ukeM/D�$Ct�
2�`Lc��f�x��GB.D�4��M��K��hx"B۰�@��,D��!ՠ��`	���Q{�\9�%D��Ehd����E�-92�P��8D��!a�K�p�ܘ�C@uT@m &D�\����,~	&�1£Q>�,:�*"D�l��+�%R�BC8q��誒C=D���agT�,)L�E����Lʧ/D�� ʱ)�҆{�t"���n���!Q"O��b���=�����Sm���3"O��gXԙA%F
Lt<rf"OJ�����G,�L�/@UI$"O�E�A%�9nrH��S)�4��T"O��U)W�<v䭱c�~ �l�"OX0ab�*>� (����jP[�"O��z"�&%�2�����_�t�A�"O$�)s���mY�U{@�
R��a�6"O�ț�@*�hIЇP1���"OxU*�� F:fH��� O��i�T"O�d�M���Fyi ��)s�0�"O���h4N��r����:9 V"OX�q���+]��ІE,,���#"Otq�b�Q&q:Y1'�J�7��maq"O�+��*��B�z��usW�C/~R!�$�=%�IQ�nO�{�jt�1��'%D!��@Y�hua�X*�@���,
'�!򄎄 �`DR�#�����bA�!�d�7w%�c���|4˔��G�!򤊁(�n4�rGαLSn��sM� !�D�Ҹ��ኇ9O�8�ȣ}{!�DN2X	D�*3�`�(8
W� �!�dR�0���y\���$N��Z!�䜹sx�Y;��.�ѠB�#p{!�d��%��������4?�dA%��7l!�\	؎��r��/�M� ��3pY!��ۍs���B�ͼ3�^A���b�!�T&}�T��B��v����VvF!�dE�!,�z��B<nϒH��"��A^!�� b�BYG��2>VpXWB/y!�d�-.>e����$i�4U��j)@+!�$ʭZ�P�P��c�ҽP��'N!�d���Ya�L­,-��Ϗ�!�D�=7�4� D�=���2�@�)�!��!�dU� �Ϋ!�$'ɛs�!��Ǡo-H�ѷٙ[H���'e^��!�	�]��	
�#ض��C4)\6H�!�A�:�6,�S3�&y�R�N�\�!���Tf��¢��q�AW˖�;!��Ƽ��QCcX�GДqJ�i�3!�Ĉ�=q���D�;�Z�k�-�[�!�ˁ�x���Л@̏?v�!�D��c���sǉ#Fܺ1����a�!��Z��Y�o�)?V谣��L:!���B�[��H�I���ק�["!�Ē�M�hX8p+[9m7t�' �9�Py���3���u�$ HH;d�K��y���W���[���
Ge�!�"O�a-.�Bt��B�0O���A"O�\ ���2<<*��:����"O���양9�&�)�J�k��Y�"Ox|���=�R���i�0�܄��"O�\Y�KѫO#��j��#�m�t"O���Э��n3���̞�C���"O���]&h�r�8��8=NQ��"O����c�3h�������`~��B"O�V޺%����Õ4	*��k�<����K��U1���h/"Ar���g�<��(J$��!���ʎ<!�M�d�<1�X������&P���E�J~��^�#g!�)0w����J� ��5$�HJ%�GrRe dƜ�T��d���7D�x;�#�:r0E8��	7�:��H5D�L@���?��qZb ��4�BN4D��  �a�)]/o������&TH��"O����!p�̓�_
UQ�P�d"O�ȷ��3�:�c���yGT��U"O�|��""���^}����"O����"M	Ll[�ݮ"��pAR"OX�kq��i[j)st���P�Sv"O�E
5 ��J �`iCmY�j�z	�"O�Jv��M���e75�ip�"OƬ�D%êr�z Ŕ'��a�"O��M+(Y�)X�	�`�r���"OX�S�� 4˒��&���?��c�"O�m �N2:��E I<���"O�a��aC0K���E��s����"OT�Q��Qϼ4����rr���"O|�ӆ�ӠrY��բU/X\��p"O�q��OөIf�<s�bĆD>\�A"O��Aā�;��AU�B8{�N�9�"Ov}7Ŕ#ҠEQ���/v�1�"O�4G�ݠM�b�㖉E��С"O�R�O�3Zp��tL�13��}�F"O6��m=䨜!�ΞM<p�!�"O�X���s�>��
 �91� c"O�u�4DK\��C2q�l�;�"O�(�Ŭ�q��@y�!F�;�~�HB"OZԸ�bN�O��mh#D3s����"OE�B�^qJp�
7��]��ir"O�3M���� �T��*j�"O~(���5k:��Vˈ�l�&��"O4�0��`��ɨ��בY;!�R"O��aa�7~g�%!g�G9.@B&"O���A�*���1��֠J���"OP�Q(=���1C���A���g"O��Bbۙr�X����IZ�r�"Oшu�Q�v��h��ǂ�,Lܐ"O����'ޚ)�g<C/�]K�"O0��#��B���M{r���"O��R0���;�,\�Ӆ��.]��"OV0�GF�>�z��@cPsx~�	U"O֡ ��"��3�c�!Wx�!Xd"O�L� �?.ج��#�U�uP�}��"O0Y��Cg�$5�WD7W1B,��"OT��,l)�%1)��D.�ѐ"O�1z@� �pC�8
#��8�d"Op1���=&�48Jt�D�)����"O��R�J׎j���҇��~�4��r"O�ء�M�q��+� T<���'"O٢��'���iS��*\�AaE"O� 1�?9(n���B�.m�X�s"O�	ѐcʞ"{����Ƨx-#@!�O-M�~M`��97n4��D؝'!�$6;.��JƤ0.�����ӹF�!�d�1wD�SE�;\"�*bI�N�!�=m�20,24�z��M�S�!��X=4�A�w��k�y��h�z�!�DF?Jʱ	S��\5R��O�$�!�$NZ3��S�C��,�ʈ���Փ�!��QkJ�4�B�܊�j���˩&�!��Ӭ�61Ę�9�H�[�!�D��8����M�e	��C�!�dPK�9K�jV::J��V	P# |!�D�;@1��1d�@�"U�uK��I�n_!�$��}�l!U��hI����8T !�D8���r�Ԑ��F�.�!��̯W�n T�O= Z �&��m�!�� .�hl��.�,Mʵ���d� 쪢"O�� ���]צ�S�/��J���"O�d	C��~���10NE. ���
�"O�1���sՔqE�sT��ƀ�_�<�r(H�n�0`���0{����Ȕ\�<��团�Y��$��mB���W�<)�L�4|�p�R8z.4�s��T�<!#��m���;�i�@��U#��^P�<��IU�x�B�����g���PդGf�<�3�Ƿh�0��q��W�~!�eD\�<���M�TC4�j/ݏ�Jx�w�YT�<��-{���0W#�)T��i�m�N�<�Őz���у��?+�9y"�FN�<Qe)B.Iv2��R�]�O��0I�
Sd�<9#��/�T���>8o�Q��Θc�<�F�
�z9@-06-X$6��<y4@[`�<IUH��쵓0j v	�p��KU�<��$�
f���8�JX�h�|�K@�Q�<I7)�{�|���# �6F\���Q�<٥�^��.��p!�J*�V!�DNmHA�C�2��t!D_�G!���1�E��@I�_b���S�^�I�!�$A�s^9�i�?�v�
�g�"�!��[t2��QR� ��Lh�+FD�!�Ę���أ�*]Q��
�A�=5�!�R<Z͌�8�IH5/�,*�&S��!�=���`��ġg���뱀�!�䌾wTMr��9\���&�OWm!�լ�*�kJݩSv��_�z!��W�<1u�-{ހp�ħ�E!��Y�&Ā&όX�쨑�)~
!�F:�� g$R��>�R�'�'Q�!�P��X�%�'�&9��*C�!�DH���-�"d�;T�h�	�R�G�!�Ą)n6�l�d-xY�uc�ԋ:�!��B�-����w�mM�p��a�)P�!�֛H�X\�&��I6l1%��F�!�D�(\��`
�Y�Ȣ���?"!��$.ZN�K$��H�ʐ��@!�J�4��)٣ݮ$|�Qn��4	!�֤k�МJr�I ���צ��[�!�Ѽ=��L �Y�D���"�!�!򤅟,����􀃓��ly�f�,4�!�D�U��Ʌ��7�<�!�d�0@�􆖰<u�Zӧ�Z�!�$�,sh���I4���+w�'Z�!�dO$`	��p(і}^Q�t�ǈ#!�$_�~��x3J�V}Cpe�M!��LN(��@ت*�\ �wcʴ�!�$ϫo���bc� O�^�p�a �!�2�ByJBlY,-��ţU�E7!�Y
^��y�XO����&�!���Q���2��F�T��@al� ^!��4
▔K6�ipu�ŕ(lW!�D��7�Ha¥@�g�"xh�ҟi=!�DS#]Df!0ҌV�ZS�8���+E:!�䅈L�1wF�hO<Pj!֒f!�C��I���L>��ٕaޢ\��$n�^����/.�"%��H+N��"Ov��@�[�A�6rh¬h~�
�"OJ�؄m̿nؑ��!$Ve�"O4T3�F��W�(:u�I}����"O�er�_"|B�ԃ�L�&��Q"O�Q�Y>1�>�XE��e���w"O� ��A���CB�4�#�S�"��-�w"O��Ң�X�X��p��n�q� `��"O�T���М{F�8 �Y5 T��"Od1��F�7:��(��z����"O�J� _6%���2BӼv�N��"O�ipU��B�lLBe�E73���#�"O�4��� D�\���N�
b��$8"OD�w�V�l����X�~����G"OLH��*��ft�yi��Iw�Xmat"O�M�5O_��X����t���X�"O���%!$ �l�d!h=�Jg�<�#͢w�:��N���DyV	j�<a�#R'o����Ea� �ԨBg�<��ɞ4dr��6��#u�♀���k�<wMĭ[i�m�3�6�l� 7K�c�<	%��-L���xd$�[G�ę�ʚ\�<�qΕ��"h�!�S6H�^�s�N�<��D�GeΝ(C*��z����r��L�<��H�)�м�1��.^��PEJ�<Qa��as~ч�4p�12%�I�<�&��a�3��ƈ)���+\�<!���$Ex9;�g+D"$Xp�Do�<�7 ����:���{���g�<��N�K�"x����3d��CJ|�<q��׼Z��##�>PD�<����L�<٦�A��(���@��#3Br�G�<y����z�j�&P�H��g�W�<�U�ƤL�$���c0R���AMR�<��:$�H�ybUyF1�cE�<i%�E$m��q�P��W͌`��"D�<�sk��Y$td.�N�d�6a�U�<�����>Հ��n�Pt�C�R�<�f�-W
�"�h��Z�&��s�_W�<�2(׹at��DM
5L��MڐLO�<Q�@N��} �չ: ��чiXG�<���ܵ�\h���͚+nt!r���@�<�,�n�Ĭ���
 ҢJ	~�<��\�s̰9���@�0�L8���v�<��E2*�Ƞ��n�&��5���It�<��FK^�*���@ܟkW���5T�8��D)~�� 1�f�8-İ���o*D�x��dK#��9�bJ�S�1�fB&D�Hrh?�Du0di�Y��[��"D�pj�eٶ/2`A�3^6zÈI���<D�h��4(\b��)�7�2I��5D���1�%e;>���F�Y�d@z�)5D�,R��H�t/���`��2m�Z(cH D���!�Z����u#��08�$+?D������4���n��
X
dc1D�<��㓬���!.V!aTF, 6.D��a��<g��Ap��/<0D!��+D��Y�kN?<ajv�կ-�p�#�5D�Ȣ�$Պ29 ����f����F�!D�,���-KET3��>T����5D� b�,E���;�F[�'�s�4D�\9r"� t�&�Ӄ�ˈlf�\X�,D�0��Hق�>�H7<l�bg+D��2U䙵`L4�J���{��t�&D�h�PI�0	4	!A׵B��p  �%D��V��S�hj6/�4�z�q�9D�Hʥ��y)����D� ����g+D�(��YIJ�҂�T�M�*��$(D� �,�&M` �Qg 5#�H9��&D�����>����#��}���)`G#D�� �Y�e`�l�uJ���!p�*�{�"O4���(�}����AX�ynH�u"OeBAM�\
�W�.?_v�� "O@U�]({2�E!��o]h��7"O�U���j��X� LG�٧"O����ቹ}�B�
, ��"O�8C�ʟb���������6"O:�+&�C).�\Ag��Tc���"Oά��IЕF$�+`Ɇ�jE���R*Oް 	l��Ū��U5��8
�'K�IHv�Y�B��ٳ��=@��'(lq�C	0Y���yc%�4G��18
�'��	G�z:M oKR9�	�'��9
�B��){�l�=���`�'�B�S`!\�l��u�Ί�;�'������*6ќl�t��>5��8��'��}��)	J���GIr�y
�'�4d�1��<rXbcj���L`�'9;�*I��mcAI�8v�<J�'lp�av�I i���@�'}�%��ɜ�p�+��U.����'���%�Z `a �(��%}�ʄ�' �(C �	�`(FØu3�P�'ުl��m�!X�����L��k�f�
�'�� �aJ�>%B�3��Ӹ�h���'[4!*�*B~���Bd���.� �'>y�,�$:x���#��
6����'���Q$��s	�jS-��QZ��"�'s���i�#i�g��`�x1�'��8�S�'��i2���Z?�U�'Ϯ�i��#W����a^�����'�f��c%�wr���f��yc
�'�XP�NI�
<xHBVȺu��0�'�i��"�,($�i��o��Py	�'���3�	I�v(��U�h��5	�'ތ\�b��rU��+M�l*���'�T������ сIĂ#K2�'c�A���ۘAg�e�Ç1���
�'�&���-Q����̫�`H
�'V����D�6y� ߋ+a
�'���2R��=L��A�*
�����	�'{`4��G�/��i���{x1R�'�
%�@d7%(��p*��v\��"�'I����m@�xAX�����En:P��'�d��3��#Vh�&LP9���'�>Ա!c�m�Ƅ��BF�2^�xX�'r"��7��^wRXbp��!"�Mq�'bM��B I�:]���^^^�
�'ɦ� c���sV�}'�ʹ��d�	�'29za� ��i�G�Ƥ.����'f�hz��<�5!_�'氠�'��}���l�R ���I���
�'�\P;�(�s��@K$�YDCP5��'�P��-��P��<�V"WBR��'� )q`&G%^�eyU�<�vu0�'�t3���,谐��@<c�Ѣ�'�R�H�N��f�el�.� ��'��BdK��R�(e3�Ó�9^���
�'�^�slZ�VW�j���:��	�'ĲPIrgYB�i�BN(&��}�	�'�\�)W�!�jAFj���$!�	�'=,<+!c�8h�� �ᆧa-�|H	�'��,�抟�Q*� �t��a��%��'eйzgd\>=��$"ˌ\R����� ��ЃI� �r�a�_�JQ�"O`I8F�Ϛq�V�PE�@]�{ "O�ȃrIC�V%�A%�~ͦ��"O�}�a&��f���$�Q� (�"O�ձdkF/?L��jJ� �`��"O8�BઆF�=h҃(HлQ"O���)�y��؂AO�!8I�s"Od�x�G
8`n�@�_!\�1�"O����K!N���Щ(�3"ON�9`�}���BV쏖t��Գ"Oz�C��3~��� k�_�L9��"O� :E%ء_�`%()�l��"O� �7dO<b�^x١hh�D��"O�=q$�ȥ"���B'(3>w���"O, �0�P��	� Ȅ�fpj��A"Ou� ��0(��h�O�E��"O�	s�)��z�>Y�V�E�L-~��"OHM�U�X!��I�&-�R ����"Oh/Kz(�FF��g��PC�"O��	#�҆�"��`��!�^���"O�Q!Nw��x�*�7I�U+�"Oι�v��!%>H��M����U"O�!k5ʊ>r6@�%$�'�F�v"O\�C��	�(
�9Q����>�6:�"OTe���Th��$����%���0�y���:GN�p�7�^�V��\�ԫž�y��,�\bG��������y"L�8�2!�t�R��}�ӡڽ�yRnVuNP���^@�ӷ���yB�X2xĬH�����?Ĝ8kT��yB�::�@�@���d�l�y��9�y�Р �����:pY��!�y�3|v�=�+�#m  �!-Z��y2,�n��epԦ
5d�M�AB���y�R:����lC�_)����V��y�Ŋc�X�X�JC#& �0/N��yC�i8q@V̑�"��rP&T��y�,��0|� ��(M�+d|%��Ɠ�y�@�h������x��mYPŒ�yr���A�����5q�ܙ�&I@��y"�ߒ1N�
"r�К�2_��d��-lta���+f�r���QL<��D�:���YT�����
nT�X��~�� @�ui��zv��o�`���I�hSN�b�A Z&�)��
��\�,�6F0�̏R�R���P:*��P�.3�|�5 T�Ee���ȓebT����$�0�?W?X$���V8;�C�:����$�����a@�b�%*V����B2مȓ9��2��� ���j' N�q����~��q��Zl��ؓ3G^![x�ȓ�8(�OPlb���/��j�ʜ��W�3�.>@h����^�R��S��`"�
I0P�a!��+(��ȇ�@T1G웸Q~�e��ɏ�'B�ф� G`��t���H�MM�
 ��ȓ@�b��#@�\46����%K଄ȓ$HqE�)`AZ��V�^�9_���ȓi�r�⇅H.A8���d����ȓWt�� ���u^�`�0�R�z/���ȓ4���9��4D�5Rh� �.ч�'���C�@�;z�uQTN��*��ȓ	�����cc�$q�/�^d)��S�? ��#�3#2�+C֎%x���*Ol�B �?;z��sk����|�	�'jN�"wB_.g\��Ask 5����'gxՁ¾��ٲ�Č4ez�j�'tR��+\�Zwj�+F���L�v�	�'Y�Xy����I�A�`ĐUIdm��'"�H��[�����I��L�!)�'3��a6��/>��G���|5��'������T<�12�>�؈ 
�'���a�-�1�
�qᦀ38��I�'���� ��B�}q2h�GZY*�'>��Ót���k�ʓ�B@6Q!�'HXpk�� p11tl�h��P�'YP(0c�� ���&e�(��h�'�X`��ɲ�T�KA�KC>$�
�'h�@���/В�I���;�V!�	�'��)[g�B�$���@� �
:�h
�'�{Wo�4���(�7���'�PTE��l�+Ӯ�&j� �	�'��9s�I�X}���XV,z�	�'m|0*UH��V�$�p�a�O�"��'%>q#g�ܚ;;��a2��qy��[�'��P��D-F~l����'n�9�'u|�0�A�+�M���[$U��'\t��Dk�@�2�S:~�̹�'l�|�Q덭mLf)���:o!$J�'N��#�Q5,�y��*n�4��'��|jSF��3���ze��t0��y�'�.�	7M��s,
���Oǜl�\y�'��)wK�	^���f�_����'�����]���4o�I8�aJ�'�  @TW�p2b����r���':�,�`*�0)�J�Q����.��'v^H	���#ئ��p%%U��d�'1�q봈��s�~���~7��
�'�|#F�Ÿ;� PS �?u����
�'_� [���F���rfE'WCH���'���'N>T?ްQ�G�U&|� �'�f��5�ŷg�|I{rL#Ki��r�'�|:�<���aG:�6ձ
�'R,�sB✎Yn��CQ�@a��	�'x`=#d��7}�|���*��TZ�'Z�Ɱ?U<�1vA�(#����'f�E`�)�).Ere:���[����'�l#����D�7��u�Q3�'�Mq��I'T���C'���z��'��m�%Ã�����e��B�E)�'�J�q�
��f��,��bL4J���'Fi�I�/R�}k���

e��'�PͲ�Lܿ%[*a ���+Hĺ�'��QvKP�4��g��&��y
�'!D����ҭp��z�����Ձ�'HX���
�&F4!�X���	��'��i;r�+Q��볥ߖ܌Q	�'�^
4� C�� ��������'-��*fd�i9Æ@=EI�$�
�'��5(�ߤW���&BNb��:
�'H�L[A��j�H����xޭ��'����u�ץd���`�(_5w���k�'KvUB�D�.{P���G�,p4��Z�'��z���O/"`:��(��	��'�lD��� �v<bp΂$� ���'��%�7��P��9�q��h��'�Z��D G[���3��@t������� R�2L��s��i���tG��[S"O �sjO�~�Kw���1���"O�,b���r^��0D��'�⌣�"OR�'�ۯb�X�3d"���.�y"OrA�!%F	�t���_���Yr�	���ޙ7����Q!3͒��NJx��]X���]�qO,��>b��5hfJdD:v)�l��Q3�O�\�1�G8+���E�_��`���dӾB����2�����/Hn�S�-A�=!������:��UC��G�6�bIFz"��?��e�O'�FhR�|� Й����c��堄�L�X��D"�)�}�ɫ4�B��0�Kô9*��Q_�R��D��y�޴�Ms�A���%+C**��"a�Н�n�ɗ&wpY��4�?9)O�SI�	7`�3$D 1�]Ф��jT���Q��8/��o�/�ᳱk�Q�x�}�����Q��?t$L���f���ki��3���y9^!�
Ҡ�?�uE�'4��~��i�:XC�x�`��^+*�%mj����O�ї���i#0,x�=KZ�pgąk��=��'���F�!����^[H @�/G�HEy��kӘoz���u�DW/]	��pq��*o_��0e? N��&.J͡�i�aykJl|	I�L�zi
����Ғ$�x���]c�$8�f�*M$�(K�
@��ϱD1�m��Q'��]y�兿	������Xm�%�2��W8�l
�[?y nƘ'qQe_�L:�����2 }�%l�O�ä�O��Q7��Y���	f}�K��&{���J�:��P�C�L�B��(��Aq�F�,�氃Ê�H�6Mm���m�V��?��SJyR�7S:�s�-X`� �2��ɑ�r���.w��'��'6�9q��'�B�'��(
4eg�N��!D�%b��u�63&�<��D�+0'������V��F~�mQ��8�JQ���#��+e�ȭ5��,�r� d|�abm�(I��D�b�Ir�H��e��X��Ά#X+ft�6�T̌-�M�k��ݟ��h�S�TJ��1(�#�L�ml&�b�o��~�!�S�O�,�1e���HV���rmY#��u9�'c�7��O�˓a2��:\�$'>a���MBL��L��C��iI3&=�០)��^=P���`۽V��;�� ��&ix��Qg��3qp�h'��9瑞�X���<�.$��dU¦�$T����u��)j�j=���Lwd���*Jߑ�T���O���N����	h�m�N�hx	��̅abT,��N�eО�$�)�'�M3doV�1�"�7mԣn�.9Y�n8� C�4s0�F�it�p���\���H��(�)%�h4��'�<�Z�Gs� �d�O��'JI\1����?��4Y�L�ꇮ )m�
�A"�c���e�ζO���҇k��le�%��c��P��������ט=o�V5H#�B{�-k$�e��6���7[�D95nK�Q�dLa1��A��k��@����(�"e?f��� �M��l����P���O*�$ ܦ��	a��M����l��'O�$��9SK�c?���?����O�c?Q���`�Yb$)����&L1ʓٛ��oӈ�O��)oݩ��
*M~�#�J��:�d�g��
�䓣�=�R�9   �   C   Ĵ���	��Z�Jv���+�Ȱs��G}"�ײK*<ac�ʄ��	�*t�Xx�aeӀ�$�3@�##��Q�D�TʌVڄo��M� �i���$&��p�	3g�D�1�n	�/9���啥;SH0��;1@"<�6�y�$ŁV���S���1!P�Z��Yx�Q���bC_B7��ҶB�<q��ĈXgt�f��N}"��5�R���J�/��Id@H�[�Zx�0,E��1aӥ��y↊�'����D�9O���� �t2@;t�Y<%�r����X�:�"��b����Җ]���;gI���	�o>��	��5L���� ��%)n&!�W,^N��'�&�Ex�*[�	�.�`�Hb�-_�Рh��W�)�&�I�$i�<If�	�'�$����w$.P!%��Ay��H���P��O�2�O�h33N��y��X�#L*D���)p�>I�8U)~� �U��="� ���Xj�!���q�48Z��Ĉ��O~)�
)Bq(	т�L �:�!�s �O�i����	��������kg(	6Eo~�'��%Id�I�$'�H�c�d��8����R�_)Q�x)�7́�'�r��	��O`!��s��JQ�]zP�����M�f��<a�c+� ,�OtXNC�<���ս0Z�
R�O<*��䑧�ē-���Ϝ	L❫�ϑ(m-��X$�I'V�2�!}R�O 1� �>A�' ם�>R@�*�h<׆�!��^�i2��=�D�!}��'{�Yp���D��D9����&�c�OV$���$�
�Of�IQe�?@��t!`��P��a2"O�T�T�  ��OJ���O�	 D��M�П �IW?I���()�$�!-/(�$��oͦ�&���7�_:�ħ�?A��?�%�+���cl�0��U��,z)��'��Fo2���Oj��<���\ ���D�k�q
k�8cJ��S��	�����'R�'�2\���4���(C�	`��z���N��jy�J<���?yH>����?�0��Wt5*Fl�x�"\X�F�)W��������O���O�˓WȘ2�>�������#P,�c*Śhk@�T����� '������R�A���A���Yf�J5�s�����m�����O��D�O��9h��rT���E�!Ru����,��L�*�,=��7-)����O��'�p�aڇ|��4pa�3��4�?I����!R��5$>Y���?Yp��K3jNTZb�ڽ9.��s�g��Mc*O����O�y�p�?�n�$*�R�nO����t�<7m�<��L��>�ϳ~B��*t�� ������p�gN^�����r��D�O�d2M1�	�?O��� mN/6@�%fP�2����'���RE�iX����W���p��Ô�8�Fy�w1D���q��L��m� ��m�c���.�-!ۑ�rA����6,h�l ��X���I���q+t=#B��:;�Ef!�Z��' D�'�R�i�fE�k�Pad�;zjd��P�lZ>$Z�#�r�læ#C�;�"5)fd@�*�e`P��&5���p�l�+4�zh	�);a��ȉ��]ȟ���ş���&�u�'�r7�$��0l�K^�9�1�	A�ٸ�*�?v������?VZ�Xg琍A�DF~�j�0Gf�%�C�
�P?∺�*utXX�t�^���"�òlɢq�A��s	0#=q�)�=
���ō�:$�Ȓ�K�C�n���ӟhG{���3r��1[q��J-Խ�%�#�!�$O�#<���q*P�d	pOB3Q�1O���'a��
�0��O���X�+t��Br �|����}� ���O"M6��O�~>�;1�V#��4���~��D S�( *��Y�~���r�!�p<!�.�8Q���iԟ	�Di���`T�,[�v�(��~��x��Q9�?I���W0@Mb��O&*��x��m�#�1O����3 tEɥ#�<M��-����,1!��̦M9Rk�CԄ��-G�a�D|�Q�~���'�(�;�	�>�����¶F������bX� ��F��0�B6���=����OL4��(2S#�D�҅��T>=�OE�Ě�E݋1�ICA�}�|�O�`��OGیa���D訟DX�9-���Ц�2����Ք>I5�����	D�O$��׿{[D
$)�e)6<"�D]��y��6:}p �D,K��}�"'���0<Q'�	�Y��сh�j�\��^���O"��Ol����H��d�O���O�$?gr�kW$ҺT�n�[Տ�����[&����Df�y��|��TGU�B�vg��6��	3�5�c�m}��*-Ґ�}&�<Z�_;�@�R�Z �<�rb�F�|�'	xyz��|Z����7)D� &�@�t���Q ��d%!�D�:|��Yv��'>¨u(!ć9/����HO�Ny�(�t�qH�H�D�4" �K� )��T���'�R�'u��]�|�I�|��"�1�4A�l0	}F8���5�&�h N�[�\����']9s���^�B(ފ/�b��&��c�����G��$� ���5͐� ���N�,��E����=���'R��d��MU����1z܎1�`ET�-��ȓn��m;��M�Z�(�͘�B�i�<Y�R��'��@��u��d�O����ER4uưt� "���� V��O�X3t"
�$�O*�d� A�d�Bg^�/��I�Z�sGA��L��Ѱ&n����2�l�Pԓs�X Pc
?&�N �0(���b�KӤ���Z0B#�	��O�l�q�'5�eӀ�Q.��E#3�M]��*��_%nS��?������'�lV��=�dp"����?t8!
�'2^7MZD���Ag��=��Q���̋-4�D�<�������'�B\>ՙ֪�ş �1�ˡ+Y����#S��h�eWៜ��=?P�h��O��}��Ox�K�)j��@s�[	#%�����>1B@�)���򏙓B �E�� �0��M�13�}B�o72��!p�>��_��t�I�M����O�f�+���4E�ܑ3���u��]��y2�'��y��٦p�ҙ�d�w0<x�6!θ܈OT������ߴ��'9!�I��ɟN��:Ek��m�H��'��}��(R�����Z�iD�a-H��y�jϧ%'�z�C�P �4a$� �y�j�?V�[�J�{P,آ��y"X.ܬd��μ)Pp���	��yRMO�2���idn<����QK��y�N�c�p}���:�@�G׫�y�#�s)������J�P$�p�X�yRiC�_?�����<Z�Zq�P��y�K�+�H�p�ÎC@��Y��*�y��O0	~^�7.>��׉Q�yrꎘ�ā�G�jz
Q��,�yb덚,�����d�x���g�y�Gԃ�� ���Z}�,�%j�"�y��J|��M�K&W�8 �v ��yJ��Y�bE0���=F��yv닀�yR+׉]�t�"�3J��ɴΈ��y�"O8�����	¬� ����y���0rR&��J�(a���y&�9`�`k��	%2}�aI��yBӄy%N\�*Lq�^�	��yn�:'��h�V�g�Ɉ�ج�y� @�tf��V�Q'J}�U �ڥ�y�%� ^Z\������:.=ZgT �y��?.L�T��Ն
p����y��: �~�AH�#�R���H�yrF�1T�@y�g(��� c�8�yrM���e�²�4 �7C_��y2��?4�,.9�E��
?b�����Φ�PW��Y��;�-��n�Tu�ȓ8ܠ9��C$�<����;<ƴ��*�ʒF�
e���Lءi[����m](Erl�FsJ4Q��X<�@�ȓ����v�б��̈�ȏ�a�^M��@/x�d��%�T7쌆}�L��ȓD�����]�B�+G���x�q��v�m�*߾=W1�)24�2��ȓ0{bYr%�[o��,SS*��o�*���@�tD`��\�5s���%�]�f�0U��cn��P���o��ɒw��"?�r|�ȓ)V��t��5���tB
Pl��V ��d��`W0=ApA�^-B��;��a��%:��y#RρX�d]��*^t${���,��U؟�P��
�ʙ�cdI��yy�o�PE(фȓp�� ��8<�.���[(F(u��SH���ܫW��0	 �S�>x�ȓ�T`�uR� �qbP#�fא�ʓ ��%������(Z#/��uB�I�%�%(�M�����'�[�Z��C�b�ę��I�2=��]��ؐLzC�	�t�r���iۦk���r�Z�{�TC�I�z����a�J5R'(4YC�$,0~B�ɕn���x`_�O�@i��ģo��B�*m��� .��;F��PND�A}�B�1 ��	�`��� q���!>�8B�Ir�F�Rk�43�@o�HC�	��dS5��[�dj���8,�C䉥/� �z�dYv$T`��\5X�6B���h�B��[n`uTL,p:B��4.g�L���^/o�.����^�| B�)� ���,S�(d<�Z3��{����@"O(����F�y�Ft��U����(�"O���G�Ñ|Y"% w��b���@"OD��u)ĸ�hm�7@ޅ)&��h�"OJ 	��֔BG�e��,��8���"Ol��#	�x�<�{w�5���A"Of�J#�֢5�����!1Sي!+!"Ob��J�#-�1ɱ��,_�T��`"O�h�u#�r�ZC!X�o��cs"O�8��f�WۢP��Y���"6"O>�Buɜ$]�M�b� �!�,�"�"O@d�)��c��xI��oY��4"Ox�A�O�'h�Yab!Vn!��"Ov��!@#C�| �·bL�i��"Oș8�ꂁM�)�rH'.;��!�"OI��# n��9��2J>��K�"O�u���&�Ԧ�-xh��"O��C��i�2U��K�Y���"O�Ly����K}��R������W"Oy���*&3섫%"�7G�h)�D"O��Mחg$jѠ���"e��"O���&�q�DC� �:D�mxA"O�)���Ȇ4\�ZC��H�>��w"O��ʀ�C��qtHHp���R3"O0=HFG҅Qv���A�kO��;'"O�����r����(<z�0p"O� @s.�>%/�T���L�0��C"O� 0Ē*���@#.w�m(���}�<���!Q�Ҩ��9��0�e�<i�	�UCz)`��m����n�W�<A$�K>'Tx���Dɹ2老����\(<�D%��1V[��]��H�*R�
yX�'[Z��b� 7O
�@#�.C�M�	�
Ǔ�,	��}�"S�g	F)�nʈ9|MS����yr#F�M�q�P�C��n���8��?�
C%a��� �e�;3	�	`��M�<1��>?���2EZ?"A�굫Wtܓ$}@՚����;s�`n�iB�� H(��x��M�Q��$%����H,E²�(�Ҷ��xd�SN �s�8L+l$:s�؈�y�N�G�\�1�a�?�	����
�y�CH^TB��Wi�=m��ҡO���y���4z�q��Ԍs]�Pq�X��yr�<���ͨV� l���yb!����D�gl],d.�9	S�Y1�yb�Z�s��R�o�d����l�%ƨT;ShI
�����Bd!A�p sJ1k%ӱI܌�yҪW�8����Q�Zx�K�ې�?q�S:i��ۥ�'\�"`/�_��&+��D�ZJ�VRd$� L����d�?���e�Y�\�b�J�[�!��ˣMϜHbL����Ls�Lͼ4��O\5Q7'ݞo6<q����:@��}Ae��E��s*+��C䉀1:�r6HB(qN��y3닥8&
���'$��OLF��OP�XF]t��CF�ij,@f"O���Y��� =e��3�iӼ`:'�Δ |� ��I�MI��R䟯d�� �QJ	<x-(��$Ii�~�PN+
66�T?|X���eZS]��P�MY
H�\Ճ_��?��C�	k��ѬJ&��3f̓
�&��7	 �Y�LH3 )��r���L~���[��b�*_�g���KTd�<a���6Gh�G�q�u"ԣ>v(N!hw��=�����B�?E�D�W�yb�N -K��؇ʝ>g��k$�K<�yB���u��%����10�x◡��j�YMO�y[����>Ѻ��G���5Pў�҇L4#��5��W)H�fh=LO�͘T�ϋT��X1�&��^��L����/
�FՈsl�*�Ii�B��H��Fg,�O� �zT�ցYS�P��6�$H���5vw$I��Ȑ��n�3�-p�PbuC�|b1NU� `�ᑣU��`C�oi�<1��/N����E^l\
��r-Ec{���!�n�d����؊��T1���ەT��B�u�b��� �zT�c�T�O��xBC��θ'k@���F��48#cE=f�F@
���1��D��
Q�s�V�a"`� �.���V�[(Q�8�p�?^���˰ң)�d��D�/}a�C[1O:@C�i��`�0A�?G�N�p��ӻV/��S�H�)��$�D'��h�.D^�����&7ذ=��DD�Ec`�a�m�mV�'��:G��&,[�u���gS��d�S�(lo�?�ՃN�v˂�(�'���j�e�*���Y�N5�߂>� �bD#�����Eq��,�W�&$�0��q͛N~b��A7V"��1t��d�I<�hљ�Ǥc>��	&i\���=�$�V\��؄#^�c�vC�oN.��͓��D;g� 49f%�$�F(b��Fy�g��t�PAI6���!�����#- 4��=I2�4D�#��'���I�ϖ+x	��1�C$�a���&O=츀��K:#�T���Bw2~h���9z��Sf��1Oz���n�B *5r#뗦o�>�!���/9mv��Ob
h�%̺%�����lV*+�<��'��0$e�<�h�1I��P�5Ӆ�,����K�[�(��]�(�������[>{�l��`������X�B����m�f�6,rdB��.v�re�~&�Ha���^G��P�� Wx���/4�| "�F�C���٧A�Y����wnV?`�h�8�;�Oj-��C�.V�(���IV�՛�"O �+��S�t���ޛL�f�Z3"O�40��ǢYe8��AM�p�`��7"O�����v�h ��O<>` ȂA�*>2xp*�}��M��D7#Alɉ�AY5#�`9B��!�P e��y{aΑ��|(���9���	/x���E��'�q��Y�T�4�����N�72r����'{��Q����{c���^^��:cI\7c'h�""�/<H1��I�TeڀI���0*ְ����9G�ڢ<14�L�Pmʢ|�	�W}��R����Z��X`.�?�Ȁ:�'Ŷ GE� �E@b텣HȾ �4`踀�����? �Ē�4���3%�Y#2j��Th!1!򄒃u$� �"@	7?@L[v&ǌq�j&n�؎���+�1����&I���%-��yB��}�	rЇ�����d����'���˓x�Z	��N�?��W&I���&D���	6J"���OƦ����1b7D��cd@�	e����C)>�%�Ү)D�����
�c�>���� ���Q�'D�<�4�XiyF��G�,���1rM&D��0-˯=��kī��A��j%D��CPnF�hטia`�� T2�&D�P1���oAԀ����(��q���(D���e �^���A�	ݺ*z�ys�(D��A�)��r�%��Nb�AR�'D� q�f�~H�dAf.�lf��Y�,(D�$� �'$ԵRW�ƒ�2#D��07�6�H+wă�T6�d�v#D��8�*�+X`���V^T�B?D�@�ʁ@lɋ����ةդ1D�ѕB��m�`�3�8R�,@3��;D���t�ˍc�8�T�ۤd��`"BD9D�P2w%6f
=3-Q$��h�H7D� RcM�%ph$kBۚd���	5D�t�"�=)Ԛ��M�"*���0D���F;�X��/$C��A��,D��i��,|t��&�Q�7��p�C�.D�i�B	l���I
�k_ڴX�
,D�����U�H"�Q1TAA�\]^�9�/&D�l۔#	W���ف$ߎn�H$KSL6D�� �Bܣ��2poѶ>��5D�H���Y�����N+Nz��!��)D�웓��-U�z��K+���pwj5D�� &	���D�.��CД'��i�"O��H�`�Z|����	]�zK�"O 9�F!�8 <����+�X9�"O� t��D����X�g>�QW"OZ8�	QC�c��K�\pzR"OȘ�������)b�+S���t"O%��	НC�2I9����\(�"Ox ee���v��@MA]��\�"Ox��dF�*��xa�k�u�R #�"O�y+U�!wALa�I؛���k�"O�0�P+Ÿ�p�sGI�T-(f"O�ۇ�<�`�Eg��G4����"OTİ�)�!Nm<�*2��X'���"O�a�tc�)��{� W!�e�"OjE�E�]*tJ��w&FUH͹�"O���'�֠;�]"98�I R"O�yEm�3rv���G�*|�is"O���L�f�g��.��X�F"OՀ�,�����6 ��-  "O���b�-��}���R6ƹ�"O�0u��!�,d���)��TA�"O��x���4h��-��Q�H��B"O��&�lq����]����"OD��s�pĔ�y�a¤@��
�"O�X�ǉ��`�8( $V#��p@"O�p�h�>|�2���D�ɢ"OzS����1�*�;於T'�\��"O�u�7bف�f��vo�h](4"O��
�&;Ca�	���ˆT��P��"O�`�עV����pb�S�Hا"O�p�⩏ 	"e��Ϟl�8��"O`a���)iat<�g����x�s"O����9��8	�)^�
�2"O���ghD�_\� S�W?b��4��"O2�SpF�
?�)y��^�<D���"OR��m_!�R���!I:'7J��r"Obț6)��[N�y&.��34��k "O�U�r�L��I��g/H$�u"Ox�j�M��2�B�N8ڑӕ"OT��g�����[��u"O�T��<�����vyd�-�f�Cd"O|���[�`���1���H�8���"O��4��&��i���
��Ju"O
���L0� ��$�"�2q"O&$
K��&��!�c��7��9Z'"O��Fn�H���K�%��-p"O����M(J��ڱL�	g}��8�"OB�3�E�2�vX���č�"O֔�4(@�rH��hě��)�C"Oı��L� {������
?��b�"O�l@�M����2F	Y���"O���O5S���8A
C5PC`��"O�]�!��6 $8:�֎k��Q"O0����>	h�i�� ���"O|�)�K�ސ��&	N y`x�j�"OT�;v���X��r���F��-I�"O\���(ĚѬ���^m��P"O&����>-�$�:_��]��"O�}��oV���Ԓ#���T"Oh	"@E�[��A���Q�� c7"O$D$�����E��l����P"O�ͣ ,ʹ8��q��K;�`]��"O$�BG"��4�.�'��,y�"O�l���Ǌ*{�,���m��|Z�"O� P�q����� ׁ�<��� "ObA��Ĵv'��i��O�%���x�)�`��t0DA����ՈB�V��C��4����I�+oƒ� K�C�C�Ʉe ���͇..
Ɓ�Ӈ�аC䉶D�ru��� �����zdrC�I7\4"��ˇs\1�떩7�.B�*>��i,%!��Ɖ��zd"O��4�HJ�.�҂�L�/@����"O"�x�l%r|��2��R ��ـ�"O���.���Х�fĤ, X��"OV���n��.�*!(�.w[|}"a"OP 	���<ȡ�3��&Hf8�T"OPI���T�����#5_%tp��"OJ���	=]��A�S�"O�%���E
���n�H�"OT�p�h�+>7���o	l�0��"O^P�f�ǭA� uA�P�\��}��"OB�9�J��Y���M�/QnL,�C"O�Bé������kB�YĜ�`Ò�D{��	V��v���/	p������0!���o&j`�Bh �@e�1���!�� ja�$�ƫ�Դ� �K�@��	m����$�I�C�CkW��P`�r"O�M�bᜅ+r(�aj��u�� �'"OjP�g�V�Ej�ڎ	2A��"O�,A���W���ÆG2�lJ"OB�I���
��I�˄*�J!kA"O��0'H>C�\˦ �2�^�`�"O�,���M?/�9H5�&z��a�"O2��҃�>+=x	4@F/@��X	T"O��!���g��$�7��`�xE���7�S�.��R5��Oq �Y���1YyB��]T�)r���S�X�Fo��7��C�	-��-p�jí�b��4�QeY�C�ɭ`���y��N6E�6�K�,/4h�C�[KZ�j��D8cYn�y#�ʾh9�=9çsMV0sF��$U�j�p�ƙ.��͇ȓl�Z�: ��y<����DÍ]�l�ȓu����F[a;���GJ�|k�L��Į�������6�:w���1[�,�ȓN� s�ܲkʰ��内I�=��{@���Ud�&�f��r/�=?Y�y�ȓa�V����P{��6I\��L���-��rB2��0#��6@B,�ȓ?�:]�e�J�j�`�#�@�]�`�ȓQ��y8v	I�r�Ak�K�$r �� �4�s�y��1��&����|�ȓY�8���$J|4��P�NP���ȓ^����ǯ��G�N�X�;z��o8�� o�
D8�
éQ��Յ�E<�Pe+T$��@����%CL��ȓ<�#�E�r��!�cY�D��ȓ#�QVj�v��iB�eDt�Q�ȓShL��T�o��,�e% �g'�\��6U:��DPd�b���!��@��8�	y"!H�'�遳��r��e��~�F��q��.��ᡔ.��(j���'&u�D)�Չv��3����S�)��%^�Xe��I��2}[�D�ȓJ����$�q$����V.f�ń�m���e��
	T��CR��3�� �ȓ	��thU�ҌjpV�ۀ�ڕv�i�ȓ~f���7$K%K~A��ߒL�x��S�? .�;aj�m7<Q#ܻM���X�"OD�a�݈}�>)ጪ���R2"Op,�3.��u�:l;V �z��"�"OF�P&�YZ�	���"Ԉ�"ODX��D�H�H����58�
���"O2왰�2RD|���ϝ����w"O<�K	��ki��J��Ɠ?(�U�F"OX�v-�8Mk�3��,z,�p"O��Y�oE�M�>���(�g0"O�@��F��`y��K�d�z`"O��Z���["rL�2���>Ԧ�(�"O^h�UB�S;l��bL�4���{�"O
�F	S���j�_10�ĥ��OLQ��_��|���F݆JW>�[5Bv�<A"JEĭQ�����m����|�<)ٔ[0��5E�:h��[�Vy�<��lB�)��8��ԳuS����x�<Yd'� L����2*�@v�<1$"���$��dÈ+X8�� au�<!�H��L3΅� ����Չ��z�<����(E�^M��
?���槚t�<�1͆1����c��{��Dyeh�<i�候��P�,Ѣs���*�m�<Q��W���w	۵V������C�<�����f��xx��	�L
 �
Bk	k�<�vFL,1ò�i���	�.���,e�<��Eĉ	�Tc�iο�4�[&��w�<�ԇ݀NxV�@��! 5Bt���l�<Y��F9 c�(�Хã\����D�g�<)��9#m�S	�9v�
O�<	2k5n�3�� -��dۑ��B�<�a��6X������M���KY�<�u,N8A���3��Y�-h@{)�j�<��";���@%̘S������e�<y�@[���#Fo���̋�I`�<�%J���b�TD4�D�QX8�LGzb�X�0�0��H� �4�R�bN��y�n�2��� K�{� ��B+��y�Z�Q�2LA�ꆏo����y��:O��pp���x�ز��L��y�'��V�	�G<֘�Q���y"(S�-�09A��~�"a�C��y��G^����5L�|P+��A��y����Mis�/C��� ��ybl��<�Nqx��q�du*�a �y�O�,X����lGc���c���2�yaX����'-�+"L�d��y����pd ���'��Ū���yR�"<Nl��
�`h��`P��y�cI
GC���U
�=� e�F��y�eD�UB����vtޑ�$C��yRf֩pϢ){���k���ʣ(A��y'�q��8RR�tØ9�Rn��y��T����,��s�����F��y���*�fزQ�/u��$�@"0��ȓ:�f�Y� :�zͫ��
����G9%�/~&bx#�S�X�9��S@�aQ�Ӷ�ٓ��ʶ6��ȓ9r-7�4��V��:3�n�e�Ce�<9�O�1���e뇟o�؅��y�<�E
̎-bua(՜0G���"Hu�<���Mr`�Y�3�Ab�����Ai�<��I�Cz2mС��FPj���AP�<�7�ӵ+,\R��8���Ԫ�C�<� ��bPa�v��	6-Z<<��M�"O���6#�R���Q�]$�N��W"O����ޅL��d�3�?4A\��q"O�8Y�Nޮ|v��b��g$�:�"O���F��+���G��I�};&"Ov��@��	_���G�p�Z�!"O���쟅y�V��b%�� ҊY�5"O�؀���.p�[0��F����"O~=jd��.�0A����6u�xAȄ"O8�
���O�NAp�9^r��"O6lxU���(>8l�����K�vmcp"Ol��#$�\��`�I�79���""O����ʟ\`�!G��4��B"ON��JЧ�<
�[�^��tɢ"O� ���Wd[
aq̒#qx� �"O��Z .W8Qxhi��I�i^��%"O��S�@>\� ����2h�y �"O�,q���ygpCK�w�Q:�"O
L3fc��L��S�RZ!��"OD�7�!QX��B
)Q>pC�"O�QP�O+Krxi�j;+4l��v"O
9�rG٥L���g�̴o�Q"�"O��R� �([Ԋ�Ň�M>	��"O�����^�`0�3K��P�"OjY V&�0�|�ѧ%M9{��U"Of�Ԃ�P��}b�k�@T@�"O(��S�ל|�m��c�2)`�QV"O*����N՘�U�ٓt���"OP���d]([>��@W��8-܈��'"O��"eU&)C�`�@�>��e9f"OP�����BQ�UK���6P�(�Q"O���@��;[P@�Gˡ� I��"O��pشa����9a��
G"OT���&׻ǈ0�F5wB�-C"O�����)G�(���͆&)dms&"O��J`��'[��D��Rf�0�"O�M�f��6���ҦE,yu"O��S�M!b"�Se�z��`q"O�a�V�&b�@JX(�6�q"O\! F��!H���"*�B�� ��"O
U���J�蠤	�����я½�y�^\'�q!�R�I�}	d���y�&	,+��6��8D�0d/���y�d8l���a��j�4}4iM��y��D�F� � �a(	s A��y��ճ)����vK�c�" /��y�cP�ģ�ױX�њ��U��y2��Zf~Ur��̕��B�Ú2�yr��)JtB�ɔ�����͵�y��өv$8Wo��j����L�yBΐ�=R ��C��PS�aɎ�y򀐶o����P�r�(����y��G1k��02mA�l���FȔ�y�	F�m� �a�n��k:����C�yb�Y�(�����6\��� %œ�yb�_,�x�+��=48�C�)�>�y(E�&7N�O��-������)�y���
9��E�S�@�x�b���o�y2Ǖ�{�zP�0.1q�ĥrvf�&�y��C9w�$CQo�p�.a
����yBB�rI���R��!^ TI�p��$�yb��@6�
%�H[�@QR�'ȑ�y�a8`X\��a�('�Z��ǃJ��y�	7P6�l7i&���q���y
� v[�aA�4�(ղ���6FK�lе"O6��G)[<n$�0�G�FG$,�'"Od��VɏFn"X���E+
D�Ĳw"O�"�:I� \�"���z'��C"OX�Uf�y ,��"��;�(�"Oa�B�'�f	�g��O��A�"Oh}��͓�9��)�����8 D"O�0�'��k�j|��
� }N�k�"OnA(UJX�8�~<AS��hz|,�"O��.�E�^ �4�\!oV��"OU���ɓ�Tኖ��G�����"O�� �
+��܋�d�Q�"O���\1v2DQ�s��q�%�o�<�Ǯ�TpT�J��I�m���N	o�<!�%�e~А�U`	�a	hmB"΍F�<iD����F�VZ%"�.A�<����z3��jO��q��GVz�<aF��|����<=�ݪ�$^�<)s*Uo\�-B�H� K���N�N�<I�
�6l��i{�懂bQ��)�K�<ٲ�I�U��A̋�e���e�H�<A�g	�C�8�#��B5	�T�Bc_E�<�b�;8�!�r�+6􎨒1,�}�<1al[�};p���Ş2f�$�wa�T�<QkY^�-:�����4����N�<�
Z|:�ݺ�MQ?Q���ƆV�<9q�^�\�S��ťv�� ��X�<i��0[O�q�"�$)1޴HO	J�<+� G  �1��*hd�����^G�<є��_� ���*�%}�H�Z��BA�<I��J�{q"��o�q^��Z�MCW�<��h��(��=+L�s�O�<)��Z� 혦a[�
��Qۡ&�g�<����/��eh��ǡJ`<󰠆_�<���)V܄2p�I�a�fKp��B�<)�L�
�B}�ď@�]��"���T�<q�)��/����f���҂�KV�<�sd'k�(�y u�LJbJ{�<���!#��؀�J��Iu�Y�0Ix�<�eC�y	�`�"Z;+:�9@K�_�<�#O�:�Y�Po�C7J�˅�T�<��B�c�(��p�&D��3g��k�<yPfQ�g"�=RcáB�P;��h�<A��޷t���p��₅�O�<,D�k;^�1�Q
�x]���_J�<aP��V*x��`߉�\���n�<��KU��Y���I1#��!cLg�<A`BX���:�Ɉ��E�6��{�<A�t�@��	�����V�zC䉇�P���@����!�^DC�		d(b�݅_���7���K.C�/Qut���J��~������BC�	'OM��г��(EZƇJ#4nB䉼l�����%�J�K@�Ӧ�4B�&Q�`�D'[�\$�dF�E�C�I\a���[7�&D+�@�Z�B�ɢ"���[ƈD&Y=�X�*Ҝ�C��58�8{U
�Z!@0�IћD�C�	�!���y���%p�.LI��`��d|�2�4��h5�@P�CO=R!�I$;�]x3�\�vF�;����JO!�K�$���`G��`���wJ!��6@�$00�K�z��yVj�9<C!�$V����Q�oʤ
u�H�"O� ~�$��8�е�֊4�� �"OZ0�D�\�:�T�3iX�����"O��h5�Ϧ5������O.H� ��w"O�l�Pb�l.>X�LA�
���"O�a����2$�4�B�?G~� ��"O$�Ӧ"1w2 S�H{n���'v1O�"�턗�������]ڴ"O�L"4��<�4"�!���{#"Ol�9B@G�ٜA���	w�j�r!"Ov�r$(�`����7��4��l)F"O.=�̗��%J�:�}Qf"٦�y���>2D2���T�VTІ옋�y�"ߧW	�T3�"&=R	!���,�䓁�$2O� 0�C�-[Ǣ��#fG�)T��0�'q!��]�`}&�/Q�a�ҍU&P]!�$75AF��#�.3j$��-�C!�Ϟ{�r�sl_���Y�5̍K�!�4G�V�qH��Ep"-#de΍8!�D�,r�����T.`U @A���2!�D�-=E�Ԡw�I,<��!ħ_���N���
�A��c�1��XzT�P+<D���$b�7Z�d�5�� D���^�$(���gK6(���*<D����D�0�p4H˓3^�¸ja#<D��5�Ȯ�"k^>�����8D�X*B�	��a���z�<ԁ�1D�L���
a<|���LNqb��c�+D��Y3g���9�LF�G*�hQRf+D��%�i|N�c� ��+�(��%D��cBc֣I�`�G&nY���SI#D�p�ՃHp�`�"&�j	E4�C�	�o��Q�Sk����˾�l�	�'�,
qc�0����#(��Q�'p�i
��
r����,��$����'�A�6��8�r(���Ԧ~Ni���2OB�� ��[�vdQ�N��z��r"O�rWJ]E6z�K��N:s���{w"O� qlP�C�
����|�d�B�"O�c!���J����%�T��9�"O����e�32�DK"��Gk���"O��IF	K����y`���rP�E{��I�IZq:g�:'Z�MS%.Q=�"�)�$�α'K @h�bK�6ax`�{���hO?���G�(al@Q�ۧ<{�jԪ�^�<є�ur�(�OO�֬R�ŋW�<���D���H��A�� ��!� Aȥ�c��l(�)�GӋj�!�DE,4��B�T�C
�熄�[��'Qџ,�'~L�sR$C�9*r!b�AϨ6ǄMA
�'���� �n��`Q� qDu0�2�'@�1��n��*��T�DW:A�L�)
�'����I���Z c��M�h)H	�'x$�Xqk��bw�H W�H9�'���Q&ĀyHTY�q)%I4Q����'��;�Q
D 51��x��4Q�'�:�03O�!�UI�땰'��aB�'��+���7$<0 ���Ћ���)�tm� ;z(|�Ì��[�Ď�yR+C�[�:���}�`���7�yr��:�U�c,G9e�j݃���y���J��9��IZ�`��=HaT ��xr��	�����]�Q�^Lr��4Y!�D�C�^����S� ���B'�֜�O�=��*�m	�%���jA� j�� ����Of�=�g�? P�pA�&���2��	�x`��{�"Ofe �X�NhQ@!�TY�H�"O�̳ed�(2��Pv�Rb)^�*�"On��+�VV(��R���e��&"O�rFbɍ~crtYtl�5&b�7� D�`S�^�9nX����f�Yȶ�=��5���
�RL)��$S�@!a5�	�T�!��ϫ/�*��NC�j���X'ro!��'4m��S� .:�*�E�U!�DM!4�"�a� ��B����8!�D�����3-�C�80)6V)�y��ɁD�@�jT	��3`��U@�7<b:B�2|N@�.	a2.e"G���B)"B�I�UÈ�@���2���b�C�vNJ�O���1LO�1JU�ҕ+�M�6E�'}ȴ"O�Pa ����Z��� =k��7"Od�d	��ku�lX�L	x@	b "OL�Q���?���ե7�J��|��)�D3���%l f>4���%D�_|B�I�F0w��c	�%��&�/f �C�I 5O�M[�+�)?�"c3�3
ԎC��c<*�Ң��$�Q#F��>9�^C��>:��|�U��&d<2(�p�1[{$C�ɍV��@�B�A'(���)�	�B�Ib޼kÉԯr�	;D"�#��B�I�s�]2ƓlȺ�5/<�dB��H?���� �*�MtdȊz�<B�I�f�=E	� �I 1�ۅ� B�"����E$�P��ٚC�	5Pc*���)�̨���7v��C䉙8�5pӆ޿>���R�#U4XC�	r����5��[^�YC)�q�˓���h��$>��SҌŮD$����n�!��1��qs�^�C'�x��V+��'-a|���N�H��)�/�jI���,�hOn�����ʥȡ!B�Q��1�3�*b�!��к�J�� ��(�1 ��ūE�!򤞝d5c���fa�� ��,Bv!���L��� Hj>)�p@[�m��}������@����1��_���A4D�t����1��eXwΌ� ����E�14�<��b�-ƚ\���6���b�<9P�Cx�c��Ҟ��ItFv�<Y�ǎ@2�����UM^t�<�E%�o���c�Z�r�`���\D{���
*N�f�1�\3�4�:���O#vC�ɪ��U2A�X�?�Y��FF�H�RC�	�Oـ�*2K��,
aeã3tL��0?��)�����X5��<h -�ey��'�v,0��U$p��IIbJ_�8��Q�'�4`��2SyFۑ��8	pyz�'<���E�D���$V8�D	8�BOk�'�a�\u6dhJp�ƴ;y�Sk�+6DC�	9 ��q��R,.+�emW	iڣ?��)Q4~rj}£ T�� kb��aA!��KрXP���N��A+͢ 2!�F�$�S�=kc����j�b!򤊊1n�U}��jCҝl�!�dآ	��A))Ǧ>�~9�S+�!�� /��;�'� l��)dD�!�䒄�|�
���V��)3���o3!�D̎j�y8"d��~cGo�b�!��U�C5�@mH�J_��bcG_�5�!��&�<��Èξ=�Z���@� �!�� � �Re��	ږ�r�^	n�ҝ"O̼�N��o�XQ��N:�!�"Oܭ��-����H07�zb"O<�R0��f��h�EX�w�����"O:���`��2bTDk7�Y�OT���W"O� ��N�[ɠ��;})B$"O�<:c�F�=H8��t�d�h�"O0m�'�:B�>!�#��K�.�1"OX�
�F� k�ySG�(M��P"O>������C���0#IR���"O0�A�@[�k��4cCΐzT:�"O,��F��.u�d���)��4H�"O�CD���&i�c���Z숷"O�|�lQ*��lrC-��;ɂ��F"O`�����ЅA�oW��x��R%"*!�DW!.���ገ0�RTjƏ[�Q�!�D*e�Z5�F�R��-�]b�q`
�'D"�Z��I�
�bЃ= �u+
�'�d ��S99����1j� �P�'
���a:2~��Km�1��M��'|5�R��*FlC$��"'ݸL�'��A�5��=n�pbP�S%xH��''�\A�ĬC�٦m�R�! �'�Pxh�c��D@��W��& ����'Ӕu���_�t��|���ne;ߓ��'�L���3p�c���([;.��'n(UZSK��Iv���e�2�'��uqr!��p_p�K�Iݺ]�8 ��'"n3r�� ����AB�]~J@8�'�� �E&B6P(]�P"�V�lX{
�'�6��7�)*^&�Y��G�.ݙ�'wVR&&�C?�T�4Γ�}��'�����ހR|r����ֿ"����'D��6�тZ
��a�����JD+�'O�)��W]�t�1�a�&�*Y�'l*hR�N�m�v H���" c��R	�'D�5RW*J�I������%��ī�'=�uhr���3<~ī4���F=��'H@̘tg	H���ѣD��c���
�'0���%Ę�O<:��&(K."�|�����:�S���FS!)��u	ƯW��F4�Id<!�ѳH�*m�*��b2$Q/�M�<��쑣r�@�[�KY�	��y�UJ�<1�H�%��K�0��HZA�WD�<�2�I�a�(�r��b��HjC�HB�<هI�6#v�Mi�l�"1�$ ��}�<�N��֑:GbG%��QU�q�<f�D�HL����I�#  ���x�'�ax�K�4-p�*�D�:6� e#%���y���%Yޘz�/�=<.�YPך�y���c�^�x� C�1�Pa �*�y`� ���Tk��0hU��,Z��y�I�7c �hB双tu��k�"�yb/Ե$�`e�� ����ȑb[��y�`��t��|ʗ�(��5�Of�G�ۄ~��ds�A���)Y$"O���,O")X� ��3�ڡk�"O��Ţ�d�$}`u�i��T�"O���R!~`��!d��-�T�Q�*O����醩p���U����'j���玃^X�A�Q��]m���?y�O���Ɠ ��!C���b�H7"OR�T�V�r����S6b ���"O��P�!� <�E�����
��`�"O� �)�O�0rfn̊�` &2�.�B#"OƸ��	T�P�^=� M?,�.�z�"OPe�FC�PR)C�/w�0$
P"O!��be��Ő�N�	��d�q"Ol܊��E�T���2�]�@��h"O6��s�ީz}�p���ܟJ�];P"O�����\�)�A�X���%�e"O@�˗�=H�\mi�	WaSVE"Oޥ� ,A�IH�{碍(�2"O�%��J$V�e0��ØC��슓"O��F�2<$����W�zlCt"O�����C=X��,��	�lt,�"O���"�?J�9$�v���"O~�����L�dY�"��8p>���"O��f���>ET�s�-W�z"O�Ya��N�s�&�!5Ğ0�*O"�ȥ�U7���*ۋB����'s>�CGJ�jE�Q��#
=��H
�'�����׵��d+vw��[D�<�o� r����kF=h���shB�<� �]��Q���sK�,rG�c�<�%���&�h�
^?,�4�A2BFb�<q+֊ ���S���72t���۟���s��h���&)]R930e�Kཇ�{����Ud�s��:ȅS���I�<I3 Ɯ9��}�σ&v�C$M�`�<I�iJ~������n�z�ɤ��w�<I ̃�$F���!AI(u^��7t�<�&Ā�"�p� ԮV 0Ժ��o�<��!Ѻ:<��92�ܥh{��k5�_�<a��Hm��� bX�qR^�˅��W�<�ӲAlDȑ���f)�CT��y��E�8yrBƔe���H��E��y�ꚷH\6�ڔ	��[�ܘ�`��5�y���vP4�q!f�X`�(���ydA�,?�52p M:U�2xx�*��yB��:qgliw�[S9h�䗅�yB�չ	l�a.��w5`d������y"M�R<�h�L[7j�P��Տ��yb���}���)ac	�ȱ����y�	��B�z�hƆ@����(�=�ybcP0&09���;{��Ga���yr H ��@h�KX�)W�c�O�#�y��J*	�L�#$)�H�VF��Py2A��L `���!��D�1�
j�<	Њ�fE�y��a��j=s��Jc�<�!��$��Y�	P&9�����T�<���C~�ZB-E��^}�A��Z�<Y���3�iab� +����UV�<�N�;V�K�,]|�偖(FV�<aQbP6{�T�$.H���a�n_R�<q��X�Rr��q.!ڰ���'�v�<IR$Y�EB]8a�Oe����d�Q\�'"ax��y<�E F*���VtX�&��yR!F (}�@O��p��4;v*B��y2+޲��\�V+ ���D*6G��y�.H�P�2A�Sl�HG���yr,�C,�
�@�9~�m�cV�yr��]�R����׈_���b�5�y��&��12�JZ�R��e@��y�͖�q򼅛�Tf�΍qT�ƀ��'�O� �4V�V�P� ��Dxz]��Ȑ|�<��@�rű�D4RB*VdߋD�!���&_�H)B=V�qRUnM"!�� jLh�+�9n�$�{f��mx�	�"O�q�CD��,�} ��
_�,!�"O��c4M%�:�i�����j` �"O��RJݽ?5 �v�� {�@u�`"O�*GaVq��
B��;�a;�"O��E���
���١R����"ON��Vh ̡Ce�t�-9�"O���	{�X�"�?��QF"O�"R��N�������&~|�"O����i/~.�`H�+�/�e�CO|Ep叵Wq!v�ׇ�H�⥭<D�,jR�-	#��#��U���;D��c��4��X�@K�<���h&D�`)Vو<��{��M�nPt��.D�� ��C�S��$n�2>�NQ1�9D� 
b���a�|�ZBF:Ea�W�2D���DkN�r���ԁ�(�u ��$D�x�ң�4a��%�t��<#��<D�����<[�ʈQ$�FmH�!��H<D��p�
K�g���Ԅ�N�l)g�:D��{���6|� I� dB� d�,&D�$�eNS%G~E�V/�0# �2�8D�t���կ�MA�&�C!ޑ9c,*D�ЫC� 7`�-1` B��k�k)D���d^.m���3��/%���w��O�C��!c���`�-�?Z�0+Ǉ�/��C��%��!�e��{�*�n��C�I>Ms��ð�W�$��;p�/dR2B�Ɂm'�Y��ʓ�{ ��Z��V��&B�I�ld����H�8�4�Z'�W.k!B��6!SH�[�j�%OrT�r���T���,�S�O$�и0��Ӧ�A��+H��E#R"O�ؒH�Mp
�Kw�R'X�P(�G"O -�*(Y`��0ۦb��$Y"O������,�"57��l�1"Ov�H���	��L�S�F���"O�(�f(��uw�p��eQH��+�"O�Ȃ͖9�Pp`�jΕC�@�d�'�ў"~�6A�lRR� }��y��/
��y�g�f+o�>�>�i��$�y��?������"H���y�N�7���b&�t��i����y2�#0����ݲʄ�pB�\&�y­�.��Ų
ؽ$�F�_�y�<)V�zsk��0HA���=��y��<�fH��m�Y���� �O/�yl��m����W�^�d9K�K(�y�+_����s��[�Cd�#�L��y�N�%S)>�C�<K�i)�-W��ybd������?R션��@���'�az�f�^����A�2R�p����y�����j7�S$,��x�7%��'�az�!�WYF ����t��`���T�yrD��4�6 r����$�6���y���<�^A�F�K�`�J8�%��7�yrE�F�`f�`O5i0B���x�*�3g��f*�i�,x��H��%!�Đ���x2���T�8YJ�'�)+Y!�֫G[B�ZUF��������O�!�dR�GY�)c�`Q#~2�b��]�C�!�D�J�X�I��� zݦ@����?c!�$�W�Y�D�)ɠ����La!��*SŶ�*a䈜]��t���2j!���fz� hAe�7��Y��˾3g!�� jtK���B#�jA*�+
0l�E"OlM�F�/h���IIf�6�P�|��)�l�f|�T&�5x�,Pl�p�B�I� ��(2Q=x1��i�I�	�'2����K�nŖa�%Ɍ�$V�٠	�'��e�%bJ���h딋@**f�]�	�Ø'l��c�l�
L
@Q�ѭ'�>���'2�C�(��c1B|;�,я&���2�'��%"M�RN�	��! *^�
�'�`d�ē{�T����{08��'+2�IB�,?ڼ���W��)@�'4<�$�J�f�c�j�����
�'��BueF.7�Vi��jٻ�j)�'�f�y&%̈R��U�1�ڏO� (�'^�ڑ�=���pM��D D��'�a �cH�LC#(�p��|�
�'Ot�u�^�1V��KH:lLԑ��'h9J`+ D�(�a�Ôc���1�'�Vm�Ђ�'^���0ƞ�\��Ts�'
����챒0�ޕY�(	�	�'����Q�"Y���-���$�R�'�9���%�\`�ĩ���C�'�Hd���>+�|���ŉ �����'�D b��x���yY8�A�'�!�F'�8~��reLY�i��E��'$b�3bчvk�="�"Y+M;���
�'�`��cԒ3�����3��1�
�'���0�݊~��I$� |V��
�'A|d���Y�z&�!�Q�����'4&P�7��!kh{cl������'��Ԛ`����xSN���l�@�'��k0ϏrK�YB��C*�` �'jzZ�@��
8���󀅵(�؅�
�'���y�.���6����ߥN�@UP�'D���B�($J��)��ʪ����x"M�&<��<G�&0���0�g��yR&�[�Y�wC��~�)hT��	�y�Ɨbٶ�i`M�>q���+���y�ۇ}��p�R q|Q֕�y"��c@@����&LR�_)�y"!e�k�D�H�B�j���yB­Z�@tI�l�~�P4�3���yOL&f�1� �H�%�Z�b��^��y�N]�>�s�/Ikk"iJsd���yҋ�/ �#*C0����n*�yB!�s�D� �)���@��P��y�$��`�@4
�J�!��MjC���y�/D�R|��m�$�����[��y�*�S!��91L˺H"�b���yP� ʐ�Z�ʂ�FT���Ќ�yB'X.X91���������!��y$I3]�� ��+\ �,q G/�y"�G�x2�l�>]Ȑ2G@��y�B /��I�"���z��X&�y+H(JHMq��^"Rn"$��"�yB*_� u���L]�A*�AQe�^��yb��9z|JkdN�5F���D�N��yrv�!ar#��z� ��׍P6;<C�	� ^�h��j�"�ݑpHή�.C� ��8[�HN>cM�X�&!��5�C�	u�0
FJ� l[¸���%{}�C�9�T�u��-T���B��Q��C䉿Z�
)��S�l�t��q� P����=q�'���H�kD�h�J�Q6
3xX���� i��*�P
��ڔU=J@�r"O��&�0><��rQfӐ1�*�E"OH�2ӊ��;��6*����"O�|PAX��L��N!on��PR"O���b�B�8>���a\wQp���"OX"��dPt{3�ǢC`z�a��D'�$$b�4���j�,pD��ǡ�=xD��ȓ�Ne�I]�}�h@a�BІA҆�ȓOK��7C��<T~@��'ʩvJهȓd+Ist��.r�`"�Y�!ֲ-�ȓ=Cք��͘Q%�P��ɥ8�.X�ʓ5q�ݺ㨓!���#�Aۤ/ TB�>w�*tzuÑ$�v)	 �2@"B�I	NЋQ�Q�h��1:�+Og����1;�N���S�[���)Sƌ�cF<C�I�o��4���8M
��c��
�z��C��!�R�Hf煑HF�8��HEj�,B䉄!��k��ڀ:��aL^�C�B�	�|�d-�"�5 ���g�!)�B��/\�J�ivnS�M5@����=Ah|�Ɠ�LzR˜�0� dó��`��
�'�lw�Ĺ!�t*À��#$&��	�'$p�����32�4���c0h1	�'�@�S���!c2�q��\�fQ� B�'���$\ .�D��:HL��'���ڡ�k]PX�eX�~H�b�'���rF79m��(Q�ˑw��0a
�'߸ђ�׬��7�� oӚ�Y�'��*��ܪe�d���d[�nz-���xB̟l���ё��;fqjH�����yB� ��pz��Yp��Ǣ�:�yҋ��qf�1N]�P� �r�e=�yr�R34X"d��̝�D?na���2�yr��Xf^�[6K��5���!����=1���d��t���g冦8c��۷�Z67�!�䁒Ew�`�mE>;�M���2�!�$���˒=7���r�W%�!�Dr�
�2 ��ڥc�B�@�!�d�6�� h�M�7;���7��}�!�K�D�̭�BW�
�.��V"�	C/��7OTa��R�M���Ӈ	�E�P�#<OP"<��K�n�� $�՗hoJ`�-�By2�'8�'[�\wѱ@���J�:G���p�'�f���1Й�t�M�$Y�'�bt�&���B����D�M�V����'�����i�4�r%�T鞍P�ݺ	�'Ҵi; �1�fik�_1xvM{�'��d�0��=򽻶�b�)��'��
է!6�� a��-TA4<��'��8A��C<m�$�ҕ�Z8Ba���'���pf瘼q��z�!�
LT8��'3����_��<I�9����"O 8��!ju+�O<K��|h�"O��E����BM�R���	ny��Ӯ'�*չ��ڒGo8�C��}����d1^%�S��ٻu�>qC7�[0F�
��ȓk��$@��\�氈�p�ٯ*����=7H���HQ/J�}����beL�w�<٢���&j1a���((_�Y�B�M�<Y�IH�
��#!4�8�DB�ɳn�zX ��� >��x@^�E�2⟘F{J?A`�d�e4~٤��SϾ�06+�O���><O�b�ɘ��L]=��xg`����dA��H�[�&�<5:�
�y[����S�? l`z�M]8[���A���2�T��"O�ˤ%��<�D�caN�8=9Z�˳"OM��k_"d���6K��o2�H��"O��Bp@�	�HZ��G=H$���'4�ɹ)4p�+�l�"G(F@S%�2$���>���awט���)��FNx��ʓ6^4�P�ܝ$��<Iƀ��C䉤/�⦧�8T�^؁B'-K��B�	����S�4y"j�����^y�B�ItƽpO�&R"9˖��%"O�
�bn$���9�R��0���O������$Adi�m��Tl�j!�ژdl�'xў�t~�ͽk�,y���M�,ݣ���-�y��Αl���{� �!B���&o"�yb�� �N��0˕k@��[�i�y2O�y�0Ur!��_�HXeGL�yҥK�� ��r =T� B���y2huB�ģ�T��C�&L��<ٌ�d��fi�"���s?Z	����5c0ў��ᓡs#�d�	P1�)�-�a�@B�	?7&B�˔���.��g�t� C�� C��l�W�@��c�TsA�B�>9�x��t���*�EQ@�S<B���0,}��iӢno"X��Ff!򄄺G��=#F��{�����H�i�!��aN�l��ڦ"{�xr�Ş�K�O<�Y"�%hC���d�U0.mf�"ONXR�H
P0�Sŏ�2;tJ��"O���%��z��EIY�a�"O���v��
G �Q㖻F?n��"O�y�LǡB��YE�ǢM=~l��"O��U �'`�P�Т�`=B���"O&�Jw��'_������Z+ܐ��"O.���ٞt��Qʓ�� �U�"O���V�B�Vjh:��E��$��"O��8a�U�((��� '�ƍ�"O���fk>$p�p�^�L�҅;�"O�k aX�l*�㱯����c�"Or�[�o�
 �������.�:�"O����*KF����b�%/�J�b�"O�����|�VQP�,J�b]�F]�܆�	p� ��3H��uxjqzC�ɐ%Jr�!���"_�r�ZCON(�C�ɊpU QgI_^�N����N�(��B�I�^*�j�a<Gh @�<4�C�ɤh$R]h��[2k�D��n��y�>��-�ɽ6A=�5��F#ҙz�*F�n~B�T��ەA�C�}xs!PS�NB�	�a�tI�7wI^�I�`I�
-�C�I�F�"�;b��=�T��.H�*��C䉀NM���F&]u�T0�+��%��C�IO��u�F/R�xq��� �I=�C�IƤ@IB�R$?��5Ӷ���j�����a/J4��7O�Z�skD6}�!��~5���dd���<���� :�!�¤64�sb��i�����H�J�!�D�bZ����R-n��Q����-T�!��Ñ�2@A�j #��Q8Dˊ�5%!��35@�Y0�K�0vԠ�� b�dC�I>hNp���	T���3Ս�W�@C䉇\p45�e�T��h"Eb��v�LC�ɏY�%�E�^�H3�h��R�2㟠��ɒc(8@D`Ǽuo���WoQ�_P
C�V��"C͟$D�Vp����7��B�)� � {ס�$�~�hE�ٴ ��0�"O$�9�°I�<��O�:	����"O.���eT�a�"!+Wn\57	����"O^���UAP�x�&՘P� �"O�QX4�p;XA
SE+�nՁ"O�5�%&�q��y��C]
(Ǩ�"Or�� � DR ����S� ��p"Or�{���+D�L�a͌q�� )�"O\����c]��A�]���"O()�@M�/Hi�
�N�����"On���%E�o��u�d��h�l�;R"O�!�S珒N��-R�f,�d"O<�A���Vq�M����:����"O*l���Ƈ;��ɡ'E�5����"OJ�Z ��t�:��&�6"���"OD�jB��ZDp��Z�G���$"O� )aC���X�s$˺c`2L�"O$��v�W.Z�2�×Y[�ag"Oz�� ��O�P���Ed��ĩ�"O�H��K��` @��C-��"��C�"O0���s����i�?�N8{�"O��z�@�?2�jEq�O^�cRV�0�"O�8�׆@
R���C8G
qZ�"Oz�	�,�\.Z����	EqX�"OJ�#�dRRx�h	���mM�Q��"O�MB�D��{����$;/�5��"O���ှ1�����J��Ip�EC"O@#`����	`�U)7V.DrC"O ��U,��d�XЁ0+O\9�h��"O�Y@N�1W�,�E�2O�0�#"O�q�����s�*��蠙R�"OZ��dѦX2h<H�/��$�hU�"O�����R�d0z�l �F��r"O��1�
86�����nѼU���4"O��ȵk.uQ
h����BD�+O!��ɇj���sS Й�~P�tm��;I!�$��$Q"I�����x���>JG!�䕤|��Đ��H�ggl���E�a@!�$������V>t9:m����"!��; :Ұ���X=�aP����|!�$E�\Ԟ5�S�XE/`�� �O�r!�D�;��4Ѓ��pI����Iǿn�!�Dҗ	Fd��b�,zcp�b�gJA�!��W�E�d�:��($�����53�!��\�CP/ �L(չ��ϴ�!��䎩�Ӥ��j:~��g�<y!�dv؋g ��	źa%�Oz�,�ȓ??�����V�{��f蜕�D���Hc�q*�T�UB0,��D��m���d��%�A
��_ ��ȓ��p��P�k��B�B�_�C剖a`"p�W(F�U��hE�%�C䉓7��P�P�V�u�|��D9<��B䉶&(6��g,Ϩ^=�8Z�ÕJ��B�	,D8���w���T�si�B�!(���C�,Λ�DSa�S��B��/?{��4�Q�0E���H�=�B�	����R�'��2�
)B�萙YX:C�3/�ܔ@�Q+S:D$�
[�h��C䉪xd��Եj�~\2���#D�X�`�#K'΍����V�t�!��6D��BP�ǚA��#�	��s~�8R�4D�ó���p%~pjd'�(l�ԣ�3D�03�E��EU�3&��5���A�M/D�� ��(����>���&$�D��x�"OZ`ZW�a@R��UD�z�� �"O
�ٓÕ�3����P�C1/^����`sT��.T�葐��N�.�
�ȓ"&TIw)ȴ8	������:�q�ȓRfޙ[�A��R,eK0���[�^�ȓS.�͙&I"T���Xs$��8���(q�k�I0 � �ml�ȓ3yVe�7
~Bػ�B�$gp<L�ȓ��*
��yDŝ#2�"�X&d*D��:�ʖ�w���Tf�/54�
g+D�����54h�Eq����g/�L�#D��n�f��HS�ܽ^� �*"D�dē5,�&u�7�E�k��8��=D� @�JM�_����x&��I��%D��s� TM��V���hqa�����y��*mtZi�7��14��$Js'<�y"��aV6h	vb�w���2�y"�K�
�,HjQ�LpM�����
�yR��Rb��4�b8��q�,� �y"@Mp�P��5�P�kVL�����y��"r�-R�̀O���i`�ݭ�y��&\�Z���F\�6�H@0���y�B�>Y�A8.��h�Rf�G%�y��"n8	�[���D�Ԡ�)�yB��)�\<xW�	�@r�#ަ�y�+��"\�;��O?P����O�'�y�X}���!�"H>j�Xr@B��yr0@wF�J��GS�a���ڂ�y���(t#\m�Q�V��X���(֭�y���� �~5Ip�
�X0��V�yb�ݚO��ͱ��ү\��"L%�y��=j��['�-���Hf!���y��kK��5��(h ؘmU�yr! ?���ï:�=�3*��y��Ɩz6�j��?~a�c���y�*��j�v��� ��b�P��y/�)QK4�z�͉����b$ع�yB��N�&�sS@:H�Q���y2�� �p��) �f�z� ^��y"ᔭr��Pe�I3{�>�  �O��y��	7SXv�b
���ؐn��y�h��LX��"O>Gy�G���y�G�}q�E�CNƕ:��!WG���y�߸sx�)BS/�9A�fl�&�U �y�M��,��L�rI׭9��� �J��y҄H
L<U1�I�4*O�B!��yb��NKH]���N�"����fY��yҤ�;�UR&Ж�j���C�e^B�ɟ>Ѕ����3"h��ۂ*�!w�,B�	�|��`'���;������f�<B�I!�Rю�!��C+P�L1�"O�)����fa*� )�Q �M�#"O�j��
�*A���3(.�I�d"O
 ��De�8rdg]��`�;R"Of���Lǧ5}����Q"�!�"O�
�胶^+p��*0m�f�:�"O �p�6Sb$(Sk��(L 3"O�4C MD�&�YS���j�"O��S��S?z��a��S�<��l�#"O��"�<���WAݰz�X�b�"O`wH���Jf�>���&"O�)�%KM�)�z=K���C��ŃW"O���3ˇ�'�,8�hM.yve�"O� �C�m�e���0Ԩ��<�Mb�"O¸zu�� �(��A�YӰ]37"Ov���R�7no�4��"On�"��:DrM�E���9gr�{!"O,���cC+?�~�AOL+�b�K�"O��r �"���bCwn�P�"O� Ԁ.[����k� 
���F"O�u	E���J �����?��X*�"OͱG��#/q~ �*՝E��,��"O��� 
�"|�B2�\/�F��"O�|+�KJ�+���rw
��n�T$��"O�DR�@�%d �q4�
)~H��ڐ"OL��ՃK�1֔-c��!/���`"O���*��/l�Q�O��UZ�"O,EC��_? en��X9� �GY�<�A�#���b�aS�T���×O�z�<qG�E't���D�|Hm��Gk�<qE�/1"dx4��F�`�uYj�<��!�)T��*��{E��T�fU�ȓ)�0k�`�C��!QĘ�z^5�ȓ$!���&�W
Zt��@6�M�l�����y��ܺ )��'R��I��V6����P�nĘ��^�z�����Y>-!P�ȓ,����+��dE�i�$9����ȓ@c<q�����aj%�҉�7
�Q��h��� �cc������a=�Յ�e}d:F���{d�p�Z�r��}��5�l!B�ޡr������ `�ȓt�"�!Ǥ!R�zdD�>e&0ɆȓpV�3eک{5t�����]�d��ȓH,B�!�LR;nX$Z���p���i���Ä� �9Gڅ����T����ȓB҈�&�<
�0�;��ʵIk Q��W:�!2e#nV�	�pD��t�	�ȓ	�l81�-�9o@$I�ˉ+L�D���f���F�'B(����2H:h���3F@ix��eE�2��s;�a�ȓ)*����-ښE0��I��5��d\0-y�ї]�nf�.�6U��7�D�*p>���j�(ł6H��Q�x�Ii��C2��A�d�:0�ȓ>�r����oq�A��Q�|@6��ȓ ^�z��ֲ���	A˗<7��͆ȓw@��*^(%&���!&�����S2�)�fjȘ* ���1�țA�<4�ȓ!�V��5C���tQa�$�L��n�葐1�E�Z<>Ĩ�c�*#*�ɇ�u�t��k�X����Ύ���4��p�h���{�X�q �}�(4��n�������A�ȝ@�����-B�%�$&�Z'�IZ/L(��ȓZ����?W��u��_��"O"h�s��-��,5d[.��T"O^X0F怗fB�*ǬN�jVZ�"O" ��K��!*�ꍲ'�4��"O�S@Ԝ5:�4b�����bd"O|y�!b�
*T�����D��P"O>)���	jঌ�������9"Odų���|$2�h�4�~��"O�4��̐K~�:���נ��"O���ڐ?�Pt�"
�i�`q�d"O����O�`�W�F���]�`"OZE�Ѥǆa4k�~�:M�0"O>"�"��v;��^�ȝ��"O� � ��� QL��+ �K�:��`"OLPCCE9�r�� �Ԣ=�h��"Or�EI�%_�j,��N% �q�3�H���)˦�:�P�Igk�W���!��/ɖ� �C1W��hE��^7!�dS/�\�F�L/C�rh��G(/8!����upAH���vѮ�Z���d��'�
#=�~z��ǆ?^� ��4Lp�	�v�<ѳK�85�lX��B�"R��@�G[i�Q7�zr
�lP�EA�.B&�u�,[��'�ў��8����(�����2T���I�x�<A�%T=bV�,Q1 �j�l�uy��)�'	
 � ���/a1��Qd���]�Ɠa!��͎
cv$��a�Q���'�������J6�2UCA�I"X�@��OPL����T�h-z�Iwxz���*Oس��JG���RE3m����'@���HZ�F��S�]�=�~�  $2$�k�F&$\���f�<G��q�<D���Emڟ.�B�R�ˊ,��uz�6D�����U|�.P�a.���!1�'D��ʓ$N�S}:��ƫ�"�qt�$LO������L
$L�Aգlhl��э!��m�������,W���	U��du ��!�b�I}�Oj��0�Y�!��S�$`Z ꟼ�y2 V�@n=�#�MO��x%���?i�}E8��@�h@j\ .�9g�2d�����'��q���Wۼ�{3c�W��;���?�"�	��X-Xԫ��;��{`�S�C�hB�IN�N���3j��2��N�b���>1Rfݻ���S�aKh�����_�<��J��=���gL��I��
�dH<�'�)R��� $
�:�}��$��q!��PC��3b��?\r�qd�Ki!�D� S��A�o��m�1�W�R!�D�=66�}�g��\�P;Ձ��?!��H�YMʰ��΄(
�}� A�w�!��-BH��c#�G%|����( �!���l��V���;ģ��p.��ȓ/�F}�acĈM�Yk%fF2U7
 ��
x�UXtb�'wp��BC�A-:�� ��3�BY�. !O.!�� ��X,t��r4y�%H�>��S�`�-;m
$���y��ϑ!6�#O��sΔ�ȓ�: ��,�T�i�fM�����-�������霧oν{1-ݦ�<��ȓ6����H1	f]�Ɩ3d�}�'eў"}:��ZM��qp���t��X�<��2!��\s1d�SN\995"���?��'"�|2GY�~YhDS�mRl���A��yB\��EP��B�b���R
��y2�Eu(L2d��F���Gg ���>IN<�R�H�`4�$"����>��pZ�.=D�l�Sl��&PZ�H�䌇�z��0A��F{����6'L��@bj�<�̽C��
�!�QZ�Z ��ו�|��P�˥?��d�j���/�)�"2�5BU�K�0r��9�"�0^,���Ih~B��D�Yط�=��r�G�.���/�OzP�7�A�r���p��Ѻ :�mc��'��IP~҈Y�&*��������������yO�D�YKIT���<ڡN���y��)�1݀�1�!�(D<ݓ��H
rI��D���׋w
��B@�rx̅�'X�bx���D1D氚o��$�ܔ�sI(��(On�� �1�3.)\���R&LP�j]��a"Ox��e��i�^����V0#�hI�S���	]��h��\���"�P���M0���0"O� Q�K� �x��������ې�����	�8䰝!���:�^X�Wkڇ(�C�I2���� �`�lH��C6E4�˓�hOQ>}�t�?�� �0jC"*�04j�h=D��+6��-rM"�	"+
�:����<D��+�M� Z:v�fT�%C*�!l&�Ia�D6�'W�����C�d��urch��D��(�ȓ�Va�R��=RhbD�?�F�	+O�=E�@��i0`�0e�@��q��f	�yR����t�D& -a���)��Ðǘ'��{�iȰqk�в�j� i�J�{�M��y�b�s]J�#W��=7��=XG!�&�yRg�*%،!��y�~�����0>�'���I"��LQ���}����XB�IH0P�"� �x�2��׋]>#<��'Ϡ�~b3k�J�Ԍ:�'5�2Y3i@^�<�&�&o)l9Aj�;�|����G{���iX��2!̮9 ���_C�	�'���B�){����㙺U�΁��'�\Y��@_�`���$_�Pw�9P	ۓ�'��u��͑C�~)Z�;1k�K�'���ӂ��	Z���ʶ#G��
��'N�(�FD��:�h��e�I�
P���'������fk<�+ ��f�A
�'ξF)��f�|Ț��͋3�A��'� �]�E� �2�������
�'��ز���&G��Bv� (S��	���	�M4��A�lQ�;R@ؙv�^B�����6a�?T
��Ċ�).TO����d:�',�Z #��s�,HF/��"�̰�ȓz�2hJ@�^�v�*}`�=A՜�Fyr�|R�
�*H����AX���A�Gf��D{��K�XPʥ�t)�6o����[��y"!�B�^Aw�.�zmnѤ�y��J��1"' ( �	)��y����C+�Պ����h�&�[�yR�J�=F�� ��Ȇ�(9�6I��y��Yf8����_��
5��kց�y��4@7f5!c�טr�����yR�%7/|P���iFV�PuDZ,�y�*�cORE����c�Uia�5�yҤ �1�V�q�"\����Cc���y�%G�U�������Y����r�X7�y��؁4��j�Ά�c�|�򑌍��hO�����|�4��C�"ҙ{B�S!�Li"�c��^�y�%�MF!��
=)�,3�U�4��8C��`�!��	2d8���Z�[�$�y����ɴ-��}R��4Y�D|����6l Uz0���y��h�|Qr���.}� @ ����'��{@�F]�$��2rĐ���V��p?��O.y��f�Z��A�[Y���$"O`�#��W?���CдC�֨	�	ɦqF�*]�$�@U�6Kǋmĸ�5� ��y�E��K�u�@�^� �W$7AT9��1�(��І!*P��Q�%gN��ȓ:!(qs�hҫI�.4Ӏ��!�Y�ȓ@N&�O�2]�lq���,yx��ȓ*��a��CQ��(Ӎ_�H�ȓ�%�*].K� D���.K���ȓn%���$U$��֪#∄�S�? &�i��T�EZ8�p��X�+�d�y�"O�y86���ZV��ȣ"�� 3�"OX����՞ ���u�6�"O��Z7�
C4L��
��lJ&"O�I���7�;A�V���"O8��P
�43��2���W�!� "O�� 7KT�l|�ȣ7�F�F�-��"O�% 6E$Np�q��^��2���"O����O_#�x r� 7Y�<�3s"O<��g'��0�4<���	�r�Fhbr"OTT����l�h�.L	-f8<��"Oh�a�٧-7��I��PMi�"O�=�!JeC��K��<m�ԩC�"O�){�U<6~Z3�*ډÒ-�0"O�U�������0��y��"O�`)i�q^�� �1�ډHR"O�!����;%����(���d{�"O$VV�E1C!��2��t��"Or$�B�@3�2iۓ`J�h��W"O�X�#l��'6x ����d�9a"Oa��)M"�(��U��+H��x*�"OB� 񅆀9d�⫇��)d"OܵcFZ]	�� �k#�� 
�"O��y �ƕE�9�F��T*�*p"O6���E-k�Դ)F�2_��"Oڑٱ�\0Z�F� �쐕[�d�'"O^U*��ؗK	P���*:W̋�"O~�ئ�H�Cn !����x��"O�r�j�1[�5Y�䕌t���ӕ"O�d��1;���+�"˽'o&���"O��RG뚊g��hj�띺}X�Jr"O 	�ԁ;����L�,`�@���QJV��([�J�z&�'f��@�IG�_��4��A���^ъ�'���H�Eݰ�j��s��)֨R�'��yU�ok´�FØ�}M��	�'G�g�E?6��m��ʝ<Q��	�'�D����.H  ��c�3H��X	�'�U�2�$D���C�g�lxz�'k�sÍH��F��2�T!M�D���',v�1D�E��\C- �E� 5x�'�<%D� x0Ʌ�H���
�'Զl�^,T[�U�t�Hx�8t3
�'oD�X�L؅F��p���`?���	�'B��pSj�b�$���oJ���'U��d�����I�Ô�q�ɰ�'OV�0��>S�� xvGӜsfJ�H�'�D���h��~a��DK#�!�[*2@�[va"=��p0wC�2
�!��C �p%zF$V��	��-ѡx�!�$��dhX�/z�Ze�I�%<�!�䆕�&��G�W� ˸���	?Z!��ў����'�%!<��74!��޺i-^XP�����xۢD�o5!��T-i��]I����%F�C�I>Q�B��a	�F���9�B�I.,0����\�l��л�"O@L�F+U�$a���T���h�"O�Q@˟A��@�"��v$�v"OQ�	�sb҉�'p�"O4�����Hh��!'�	Ad�"O񛖥�U4\,��)��-���!�L��xP����7�B��v���!��)z���Q+Pj��S)�\�!�$E�= ���S�\�q�iS"S*S�!�� ������)k�9&d�9sl<�+�"O��C���q�QS��N�B�= "O�iA��|���PK��tܴlcb"O^����� O�f�8ы���#"Op��3�
c1BܰU�)d2FX��"OҤ@P
W!9<
�IA.� )~�Q�"O�)s8Ce�� M���S"O\t�[�f~ܩ�!�9Cc� �F"OF"�"F6d#�T�Xp�"O�)�k09ْɔ��K1@	�$"O���4�#�ՠ���t5���s"O�H4�Y�Ǌ)�+H0<W앹B"OU�WhY������V�j�U"O�I����-
���E��]��Mb�"O8�����7P�(��C�|L:6"O
�a�� �*�)b@�͋J��	��"O~���΋�L��x�V�E'V����$"O�,
E�� i$���ɪW#r��"O�D��$�(%��N�n�V"ON����qy A)�Ά9W����"Ob�B��og���#-Ð��H�2"O�i�� \f�:����)/�N8�Q"O:]�׊0��ѓ���TU�-��"ON���Q�'ѓ��XtA$�B"O�,�
��z����+uC��!"O���E�g�F�:cU�+�L�"O�
c��?:"����V�s"O�e�ɬ>����F�M�V?�e��"O`dH���)w�4��H��%���J�"O�QY�+��y�v���G�)wTƥ{�"O2������96,,q�Ƈ:�*�"O>8R���!G�4+�F7\�=�p"O !�6 �E�P`:���<m��"O�Y��lL�/?^���@��0\�9�"OĴCr��*�t`3bD�g2��2t"O�<����3Rb��!���D�x�"O�I���=r�@0A�[��As2"O��rkK�ng�)�'"p�Ĝ��"O<m�5+φ �����.���"O�m�g��D`���T�NT��'{V)+q�K�<��N��)���8�f�V�S�0<r�"Oj�6�G<��)؟$�t[S�Ɏao��2�-�O�O!�W�F0!�j};�#��E-f�
�'�"|�ч�j��c�Ű*�>�2�Bz�����OZ���S�����j]nț�J� �,)�˛�Vj��j_f�+�M<D�	�A�P�0�,Q0�\�kt �~�0 �'*�b�R"���LFbz�z����4H�BZ�g�-0s ��U��u��HD� U�ӣ\<sd��ƣ�"�?I$HЕ8?����T�i��H�6Y�LA���S�� �tuc��2n]XqJ![�8+�iV5Q�d�V�?��U�	SXflxb�e.R�B1D���%��3�\�!��4�$L��C<X��Y�ʁ@H}{�oC�i0����|2�͍?�ݰ�w��ě%�Y���L[�q��
� ������M�(��� h��ȳ����#�Ԥ��  �M�h �M̽��R̘. Ɍ��L�ݸ._�q����@�)�џ ��z���#K͝"�pw�S�]T6m��l(7EP,�%g]���p��h�α"#�ER��S���4Hb�a̓X�V��ɶ<��G6
t�
��J&X��cE��]pU�@��S(�P��O�@�B&��ԥ IĦt�)���l9�#���Fj��r�.��(��0�:�r$9df/#�� ʃ?
�f1�O�����"+	�����vA�����Zȣca�4G�!�$��X� B�>nQ���l�/:����B!D
'{D�o�C��Ś��R�Z$�A$��ئ"<����DqF���-P�U�DG8��Qt �%��H�GIH�W4��G�[�k@1V*��v
Ԉ�u��,B	�y�VDP�`�^�x��'Q�e)Ь�N�Q\�-��lÈ�D�\��z���F�ʁ��j�v
`)b��C�ĥ(Y�hZժ�[�<� ��j"���N�Z��R�]�0�.\���Of}�ꍖD�j�)$��.�F#*f'�	4C��+'DY Z�aY�AIu�<��I� ^�`�@cፆc���jO_����a�U��g�C��U��W�@A���ǆ%t�(��I^���'��e(�L�t�H #�1���SpG
n8t`
f����GI¹zփ� ,�"���Ȩ3Ш}�'YUgJ�Pf�U릈	�U�vpK$Pq�z�O��tjQep�`���]�aY �
'T�t��ɐd����Q����l�װ���*2F��T!� \|�|){P��H��iJ(�v�S��قh_��m<p�9�.�%U�^���"[�*�j��ɮo:`��75f��7��O^�-+���=~i0dyC�N|�^�ĵ���ih��O�t,
X��l����ӠV�ܜX`B< ��-��HDȣ?a#�������K�#KL A�H56�6Y�W������K&��5n@�h��|֎}���e!HL����d�2Qد��Ob�k�f��f���i2![nֽ�2]��
r��k�=p��
���ɓl��h5�!B�/ΰ.�����3 �X$I�A/b��c��J�8-*4��	Ac`؆I��m&>s`�^H6� df��k��a�6��\���c��Aap�機�i.*1s��_�O>��]<�.��b��OUBL� �˳�R��dU?�:xr,H�>l(� ��C�9툸��I ʄ6m����t@�g�S�|1A�Y�t�H��L� u���\JyvĎ $���2O��G�̹Ak�LF��.,�
`Ito��ѼQG	�!%J0�&]+`������`[�%AA�zkҽ"�+K�4@&����J4��杪c����:�8eQ�m��`]��&e4?�v'�; *8�EmJ(X���#�j�7�]�ВfŔ�GR�m�g��)G�ܽ�/��z� DZE���b�"4�\
|��M�^���ȧ��e1�8�s&��f�z�D[�}����C@�0\�@�b�D<���F�7^)��k��Ѐ�i��<�3�E�L�!�W"ORUq���{�Ź�턕|��mT� G�͓��Q�n�V`�@�}�\AQ��:�Ӱx��D�l�T}ag��#f�����nK,!��*"�����7�& Q���[�Z��ڝ^.tS�Ps6���@� ����B ���=[*�;���H���
ʜo���D�3��Ҳ'[>��H��*�� "r�G�!���R��+�
Q q�L"&ap4B�'"\�q��:c������<*�s�{�K��% �JΊc��=[Ԉ�1���Y a��:s��5M���v#�-[plFy�<���ǯ+�h<�Ei��v�&����1^<v�r�ƢZ�9#g-�9L9�գGo�G��n���]��럢X�F�r.E�X�!�đ�<�\��KC5R��� CjcE�����(�0P3u 	7T���O=�T���	Bs�@5S=A�(��%�������Y'���!13�K5i�.��O@�v��} �J1 ���Ď�&���P-�3KŞHyw�߀a��0�@�h��M���:���e���1�-�*�b��t,S�O��i�ȓq=��M��`&�p��(6m�<P�'���P�ʣܼE�`IO�O����*)+����DH��wb8e9�'��H ���B@�x��թc�0}
EH���ɫRžm�$��|2C�0dp2�Ƣ�mk�8�P�݂��x�,� �2�c͝������KO�	���Ao؟�!��ON�%`�7�zҤ'D�ĺ��Y(U��G
��V�Ѧ!D�T���[�>դ�3c#H�7�4� D��Ȧ`�	�����;	�!�i?T���C�Bb>��'ؿ�``AA"Ot04傡F'@��&�f�:�+�"OF�����jﲈJ��g��8�"Ol1�S�]�BЪnBӊ��e"O2	��R�Y"~ �fD��^�F�R"OX��fo״cy w&� $�� "O~H8"�G\R<���˲%!��3�"OIdF�x�)���#��5"O8��QW�t=4��T?h��i�"OV��4(��1�¢ı]���q"O�5+2C�n8m���)Qϒ���"O�	�GB�������S s���k�"O�!�NY�N�W�"t�"O�%+vǖ������M��:��"O��R -�� �z�Bя�.,��=�@"O,�A�.$RKzh�4����a"OR��E�Y44��b
�~9��Y"OP�h�`��6����*uʠ"O� bh����c�T�BAȑ'�F)A"O8��ޫ<��RK�D�1 	�'��P)D�ǌ"��гհtk:�*�'�d6���c(F��f�.���
�'{ ���IAb����K҈���[�'}����×�I��P:#&E��t�:
�'�fAj�&I[������Ѭ}=�	�'8 ���O\����_,m{	�'���@!�U�2���
�7�[�'����+�>��`�%Ff�*�'\�`���A��AWbհH��'���c�ݚA����ǝz>X��'J�Q�Q@�j���c'"�v���'�\rS�:��2��	�#Af�<�r�@�Y��E����;,����@Gj�<� ���V� ���J4d)^�{'��`�<������
3��9l�G
^�<����a ��5�X+t��k�d�b�<1��#H�����	��Wp����u�<Qg�.�x� C�Řv�8����h�<y'�2.�P��c��7��Uh4H2D��h�iZ!~aF:��	a����,D�|�f�V�	��Xq��9$�xe+D�� C�v�X��$$IJ9��+D�Dse�8{�$��g��4	,<�P:D�\��윹5��"6��,f�Qs$9D���	��(�c�D�'04!V�9D�p��a9DZ,�bPJ��.E�ٺs.7D��`B����	 �dR�:��Րu�7D��b�'�lDh�ӅP�� �$4D��"��N�Hs�jN�~U!�M>D�<�����hU0���!$Ԡ�z=D�����ԻI���V�*r`�3�=D�d �fS,W�1�v"�Z�&�7�;D��Ӓ���ʘe%�Yt���"D��'��oX��vC�L,�x[�$"D�А�ܿ[6��w��&��|bW�#D�Ty��-)�y����1��P��5D�XraoΝPv����	 ����cA&D�t���޸Ea�dj �	m�\0�4�&D�4��� � ���k���}�e�;D��6��Sd���bW�x���4�8D���׉��Ÿ�n?8:1J2D�H���%��}R�d�?-=� H�I/D�X��-#?�;��I�B	�0��/D���BA��H{\E���s��)�+D� r���(l! ���9`NC�4D�L���S�T�P��� �&�^%��!D�D�b��L���B!�o��k�=D���@�܉Y����-��f���#d4D���M`��,��BЮI��W�2D�L*3���1���r��S�4�qg3D�1�#X#�4��+���䠰�/D��+r�E�z�r�h��ƛdu��ᇇ+D�(�2���t�f8hp��a��ۇ'D�Tq��B����c��n��8D�\��Z:[�X�u��	�\�:W�5D�<����m�Nu[e+W�� ��2D��1����)��b�O�9�� 5D��X���?2���7�e��5D�C3�W'I]T|�''�� yFXSB3D��: +LM�n�j��J�CvN����*D��*qE��Y�pjqnW�4��@zc�<D���� �1q2�#�T�J�b	��D!D�� �1)FȐ?;@L!�)F%^L����"O�퉦.�w�Vm�G��2���R�"O��P���	����o�F��H"O���RF�OԘYR$O��vjbA"O�T��޲�X��֎�?S��R�"OFY��R(}V����MlT9�"O�k)ϯ_������%�)S�"O�$#t--|�t]��Q�t�"OJ%*��	r�� '��0��"OZ�@��Y�l����_ V���p"Obt E"�K�FŁ\q���gK�W�<It�\�1nsuMA�0��D���M�<�A%I=sR>�i��v��FLFw�<a%jI=�rHQ&*�:��qP�p�<�C嗩{�1�#�
2�����r�<�4�	,�8!� �ݵ&㮄��bAl�<�R�Ń>���cO1d`X��kL�<1�D�3�t�� V�5& �5j�O�<�O�S���M��k�\ s#f�H�<Y�N�yא%��@E�H���Ȅ}�<��J�-��1킽'��œ�\G�<�g��Q����fa��iVЖ��<�pȀ�}��Z#��92�z���IP�<!���9��=!4n�1jV)�B�WQ�<9� ۊD��P���S�8���� b�L�<AQ�v�H��� V%}wluI�'Za�<����Sڔ�ȁlשa���8ס]�<1�*� y�Ll_'82"�hT�P�<����l��� �/�.X g��Z�<�p��$�$@y�$_(*D���F]�<9�Г!�y�҈Z�*�,I���^�<�QkB7 g6�:��ՏTZAcT+LZ�<y�0Xo�����e<���0%	[�<ɥM�NJ):�g P"�����P�<A�6���Ia�=A�!Z��D�<Q���u���Pΐ h<귋Pn�<aA�V%(d�h��� <S����(k�<�d�	'�4#P�Z2yz�I��n�<�d�!c^}@&�*	�B�l�	�y�\?- V� �@R�=d���0���y���>3k���J.1�P�ê���yB��/X�8(���*��tHT�Z�y��_2P{������+��Xpj֝�y�%������$r����у�p>���F�� �R,c�L��@���q�dB�7R/h`�'j�l�"��w.Ք5�v"<����m�V�Ȉ���%A��n[2���O�rH!��P���F�T�
��v-��4�DM�q%_�hN����j��[S��|�g�l�8d�n3� �*��x�'��n���S��ׅ ���jƁ56��mH���G:p}XB��e�����d��`P�'W #�lȴA�џ`B@��PY8`�Ű'����M
��ٕb���$ N�%��9zc�'��U9�ΘNX� K���,c	d�bS�A�n��� P��<�aKM�î���B��<ϊA�`�x>Q{�)n'P���*��ucO<|� 80p�/{H�)�ȓBr�t9�GT��@0�@°�ԴJ�N�qP�0HԀp4(�@Aw�p�O�9���80���,���a�Ʉ�G���(�h���	- ��-A�,p�$�5i�|{�f_�� �r�AO�E��,x�FM�uk�I�/u�cRnİH>��hZ$�,3d�'���X��lޠo�P�B�,���#A%+��9�C��cM",��%�d�zE�B�7j,)�5M*q:�f�#�\�cO�x����oy"��w��BMǼ
�� ����Бg��(�t���;�6l{t���UOI;I�X� �"O��P����8�MȳY�t�薨�	&�,��͂Gܔ4���Ǝk���x�X>A��V�7�9�;KJ��,��6���(����IB���Ȑ��ke��-zŬ�E@�o�0���i�H��/Y6x��2s�#���� h�{�hµu�P�
2a�>��ɗ�'��iR�kH�P���҇���	���i��8�e�	�[D)��+�v��6��pX�Y��	�~�T��C�����r��X#:��>���); 80�ݬE��%��ٟd� 5A-Q�Ac�n��*Q�*"O�+�c�|��I�3B1���$�O`�c��86��9���\&`��#RE�Ǌ:�+�ȱ�|�6�Wl�<��(���(ԫ�4[���C#mĨ22�	�h��w�[
��g�%b:���(V�8;@Y3�GH.E͇�	�Y���u�'�tY�I�����/��]Ou�@`In=���ڿ��1��	��`���F'^�x�W�`b�N���/��V1�� �S�1����-��O|<�i	&x|�Q"
���2Y��'������9a�TI�Q�G��N��V/Y�|j�+&���|�9�/���'�r���>����
��)sǝ�����GY�����Ϗ�చbeӋ`����
F��y�	��+T>���Йz_$��0��O�5Avn�U|�s�%Ծ���I9G�e�!���B�L���bJ��k�M׫4�&X`,b�l{�!]�'�p���'3�4s��CŤ ɐ�1`,�q�'	�B�BsÊ�ඍ�&�}K���9{ۚ=�S�5�B���i���fC��t��mh&
F�}&�b��NYQ�i\�`�x�c�gB�c#l���@T���SğܒS��sQ��#�D�t�:׺�I��^���Q1�I���j �V�TD�A�~�!�*�ͺ��m��1�ܴcF ��+��(O@Q��X�BA��K�j����	=]nM3uI/,!�%:���DУ�c�H���e�W�d� e�WZ<�� �i��{^���ɤ~��c.��B�ɑ��Ōoɞ�;'�0�s�ߐ5����"a{��}Ӟ���Ďl͚�S�ښp�*�i�$l;���T?hB�	4�,e�A�&����Q���H��Җ:3�`�������-��7�(�O;Nq�ӯZɼ�̈�(V�<�g�� ���)�!E^�<��F�3s�h`sU
5ZW�}���'-fZcG,�v�D_��(��	9W,���C�(a���ᡆ���C�I�C'��J$��qz����$�+$��B��!��8�Ov��� q�]�t$O�+������'�4���!h����G���c�
S�H`��#�9$���u�xh�ŪTKb�E�H�%�=)r��%���K�c;�J����@��7h�e�%��i�H��D�iiq&�zlX���.3��at�Зe0�O��E��O��Q�IfjT�CΑ F��a"O@}*��5�&�"2��;j��0���'�t�I#-�kX��Xa�ռH�.��ReٟC��(��f*D�H7	� �����#���`,(D�8��eZ8����@*�.�~�5N+D�P8NP�Z�>�۴�҂:�1l(D�@Qㄅ�Ua�@�(\$<ACr�&D��3g^�r<�r�E0>MɁ�'D��!`�2:ʺ�Z3bÛ@��'�>D��FSG")�e^�Qe�̠��?D�d�s^;O�~fnڑQh`��.D�(ˑ�Y>���a����[� D�tZ����r��0���[3H?D���!��Y;@��deX�*̬ұ� D��a�Йw��ti7��5��h���!D�����T6Y`�|��OS�6�`0�#D��J2(�#h���J�O�E��Q�E<D�,;c+�/mX�H6J�Hd�p�=D�`��Dƚ �X��nM����&D�0�UN��VB�����׬H��E'D���e��� �$g�	W��0�k'D���4%�M�6��eQ�'[�P+��$D�ddD�wv��&��jn�p#D�|�*U���Q 
�L ��%D� ���]�,� ���8X�,Ț��&D����ݑ@���J��d{��t�;D��:�M�!�`E�d�ʿD����U*O"lI'�Z�K��9A"�Ʒ7WR��"OB��Ƌ-)V6��/W%,�~��t"O� �Uc႒׎�p�һ8�@�K&"O���T4i�&�P��wɌ�@"O:�� 	\�W���c
�B����4"Oԭ�GmǍ,�����S%���"O�Y��G&M,�i0�� ��"O�H�ǅ�D� p0&� H�j�!"O��'+؊*7�Q#�-6G6��"OP��p旃a�"MQ����!�� S�"O��]�0�,��1b��hv���#"O��0���S1��2a!�=h&yq"O~�BF�$#o���qM6j��II7"O
���Y�:�1��k�:}�"O2q�UE�^?�<h��)�����"O�P�c�Ճ<����#:���`"O�Z�
�R����M�o,�U"O�1A+�	��]� KǛd�=:�"OXl���S�`P���>n�~�p�"O��r��7��
��O�6>� �"O^="֩T�lu�b�ߞ%�X�"O�{f�Кn�4с ��@���"O�1(�ͅ:�d�s`"�,`����"O�)��@�i(��P!`��i2Q��"O�H #�>+��P��M$>��)�"Oj��T'P��9p�����C�"O�µJ��H�~��R���6r,��"O�0��W�<cBE�@f�td$}8""Od��2$ӨvT��[#��p�ܽ�!"O�l`!��\C���:VD� "O�J��
ST�ܲA!�!e��Y�"O�y�m_�x������8�ܸ`a"O&��J^�TvP ��N��:u"O����FMuC�ݫ4��i�(�Y�"OJuP�F%2�p��>P����"O��`��Ʌd�N�z �ϰ]B�)C�"O�E�1�5L��YdN�r ^x�u"O���-
C���"��H� @�"ONt*���*o �k' .�(	�"Oڼ �C13���i�k�2��ru"O��g�<W�\��%���Hn��	U"O����E�=��e�Щ��U6�ԩ�Y�@8��l����#�'n�Ȱ�4����;G�8��	�'*8�sEĘ@�h����E���	�'��+���)�^REO��D�r\
	�'��]:��$z�\��8�:=I�'��@�6�$0S$��34�heR
�'�����M�$��@��V�U,�t�
�'�2�+Z�H &O�N�J@(��3�y�H��a֚��N�NjNIq�(�y"�g�XS��ןY���7�y��7R��qِ)�=p�`Ҕ��y���Y�b�Z��H�D�X����yrkǥ"r�J ڎA�F%����y2�g*zY�@Ɨ8�D���ۛ�yb��;_����+��,���!ԛ�~�l�^�a�=E���)YBe�c�.+��M $Lc�ܙ�5 F�S���F�'�6 *s���6���*4�,X�KC 2&���OR��E!�@��lX(8�q��Ù;P�^dT-?τ��ޅ��� ����>r;�e��/J�C^xL1� [�<ƈ�+�'P ��Cʉ��9V�O�,��צpՒlH�'���0��|iG�$yp�������~���C� QwFA9�t�EK͆l?<�i@AO�uf�#�O4����?m1�A�?)E�`��2܂ ��b�<��7�ȡ������F!�=@dm�d��X�.p��)��y�GE�@w^�!&U�$��Ј�-�y�,��N2|�ˢ"�%H,q{��y
� <���LI%�a��
���b=� "O�r`S'Y�la�接](q"O��/YX�����|���"Oz�"��p	`�dR�<��uC�"O ����_�>M�aM;;3R8*�*On���94W���p�î$���'��ls��Np��:��7�B|��'?�E dA�"d��|����"(lj���'H���3�F�U�^�P!
?'f�"�'�l���m��������i��'F����C�-�/J�o����'�X$ô��R��ٹv&;;ʠ�
�'_�qi�D�,P��lr��$��A�
�'jH�ۗE>�!xe"��J��
�'��	����d~����d�	%Hm�
�'���Z���>^��!K��с~�ԉa	�'�}��ѵk��-�3 �9_�nT{�'m���EeT�w���߂I��@��'�x����MNfԐC�ɬK�4��
�'�]�t�_3:#��bS M�Dj"	"�'-��2�m�)G��	�J�*���@�'�t��sLD+~2&k��L#W�0U��'켍���N;=��4�1͐�Gv|��'}�!$�O�%���#R'�(k;��I�'��8�0)ǿ�>D0�Fί�i"�'a�����2[��� EվMU�!��'�6)���ʷ$:�3�&H����'(D`�ȍ���d`�%T�<�tDq�'��Q�E��H���,�;41:�;�'@t	c���~����4#I�]� �K�'Ej�+E��4O�p\`ğYo ��'u�0��l�,r]9��?Thh9c�'�J�x�(LKX��1"�T�8� �
�'�8��0扅VG���.X�5|��
�'s(�{�c��[뀸��E�+$Yr�'�ZQ��{�b=rtNE)���c�'���Rʔ!6z �p4#9�}��'wJ���lO�.��0�n��b��EA�'����@�B,~���qC�Yk�Н1�'�^A9f�@�Yrr#Y����'%&�[$l�D�>�`���\~6��'���9�#�[���!��j$­p
�'r&�EB);aֈ!�[�g�̩k
�'�|Xb�#"�RYCP`�/q�+
�']������{B>��D�:%�䩨	�'�\�K�@�r43��,��R'�y$N�H4 �sE�ڒ=g<�1oD�y�Ǒ�c҂�٢���j��XQ�����y2.y�z]�r�M�e82��Z��y҇��T������a�q��b��y�R>A|:����	b4r�>�yr�\>)��ܒ�̿/b
��؃�ybD�����@/u�L�h��y���XWP�rt$E�-���r֭.�y�+K	�I9����pD��Ƣ��yҠV$t>���K!]B���a�)�y�n˝r���S�e�Tʍ�֍��y"�Y�3h)�&A�LD���E��0�yB�B9-�\�3��H����I��y��G�]� Ѐ���V<d����y��R�/�ƨ�6'�#f2,8���A%�y"��u�h|(bmթt%�}R�D��y"�
.>�@�T K�=U4d8��ձ�yB^�w��%IN �5�i�5����y
� .hZR�Z�lj�EQ旴]L\i�S"O|�ЧMZ���k��0�xH�"O��#&�	�|�Ѐ��4$
���"O<IYB�
3pT�����;�PM��"O��sVEW��� ��o�����"O�X(C!�I�j�c���)I��`�"OTa�S�\@ɨq���Ǩe�xyA"O��b�F�";7Xȑ'���t�H�0"O��u�*1%V0����#f@U��"Od6��)^6�c���'"(r"O�<���H�t\�-X$l�,L���&"O.=j`�0���j��qAr�i"O��iƣ�"^��x�l�EJ&�v"O�}�a�OK�����G(w<�q{�"O��b��:D���*R<*r)��"Oh��K��m ��#"�C�"O�q�e.N�3P�A�c��0K"O���d G�!a�� W�C�y�X���"O)�'R
#޸��-��'���X�"O�)��ġQ�������P|pp#�"Od,�r���Z���q!偹g�0�;�"OI���X:���$�5�5��"O�`X�p����|�S"Ob4[*M�JÊ=�MV;d�>졃"O�!�ĤË}.�`�"��4�4Y(t"O�0
( �V���)�iU�8|�U��"O6��w�ئn����@C�/���S"O�!*7G:AU�P���9I��}�`"O�y�Ȓ*h[�u��}~�Ȑ�"O<�@��GY��
�e�3vn�2`"O���P�._����[ff���"Ol��@@�!w������|k6&,D��h�A(YI `��o<CŲ�	7�'D���Seޓ$+hh��"�rM+'E"D��3jƾH@݃@�hnfa�C�?D�L��\�E�3a��9%�YX�H3D��Ie�ތ�.�b��:��y�&�-D� �`�c�
���JF�eT���6D�LbD�$j^���C�ɬu#�?D����	W8@X�PkR)������=D�xjӄD.:*���͔g_�u9�I=D��!��7"n,ehT�%+g80>D��{F�y�B�,A���I���<D��	�훊^ԒE,ʮk��1�"�?D��R� � O�x���C�R���Qe�=D���&��p� ���A"z�|T�!>D�l�)��%|�z�ڳO��y��<D�PKTK�������W)�,�K�.D����G�5���S��� C�.D�P@�f_� ����%������6D���R+X�m��S�ˋ:��U�,3D�lR�&>a���A�ԍ�q�0D��i�KO�3�	�穏���y1B�3D�X0��ޠeZ�P�2g�Z���HFe3D�8
�[�2�^�@�P7i �A%*0D�,8�"ҥjZ��e��"����//D��$�S.11�X��)C�#fz�p�;D�q�lK�?pн9Ă�	�`!q��;D��1�'��8X�-�kKVy��:D� ��,�H*\K�eOG8%���-D���N�@��I(���5tO챑bF*D����&[��՛]�%�� (D�ě�!��Z���W�Snٱ5"D��(��E##Xفd#�
�D�V�?D�� $�X��T3A��H�l�1o�\`��"Oʸ@ƞ%*�A{ @�y�8�"Op�Ʉ� �}��P%!�,�Z"O]	�m��_gJ3�o��=�f�$"O��p��
5?\�B�.H�Uq�2�"O��t��T�|� ��ŷ}|���"O�M��o\��aF�m"U�6"O00�k[�G�X\�E!XgR��"O�<��2��[�@�8?�eh�"OBD��^��%8w�r�|�ҷ"O\�3��H+�p�m���j%��"OD��f�_�$��<@B'Ŗ(r�,��"O�Qᴏʙy����1&�$���"O2i���ˀac�� � E�-3�"O�Qv�Q�Fp �� �7<ʙ�"OT�:dG)!Zѯ6m��1$"OZ��4J�c�bUEZ�W�б"O����b(H9`�*u�;,
���w"OB=)U΅�d�xm�g�NT�����"O�b��K[E������l,ې"Oqh�M�:H�$��F�K:��	b�"O�1� �*�Qi {�>mH�"OTa܀n��]1&bX�/�x�F"O8I�fH��(�<���o�(1cl�G"OTphE"F�nY�mr��ßH�X�"O�;�`҂a$�as�5I7Ȑ��"OQ���>8�n��E�;ZLUi�"Oh�k�D��H ���9�d"Ol(��ˎ[E0���㍧8xs�"O�!K�g�J��`��!ȤԦ}@�"O�p�1���5�2l���P&N��p��"O�qԎG�>�F�t����0"O�T�cYx1�1�fF�P��$bE"O.%�4
��0�p��P�\�8��,�"O>8����*)4�Jd�3=ʬx�r"O�y�%�k"���*+D���+7"Oj�J�d�D�ӦKǱe�����"OjY �n��a���k�/�<aG"O��맪��+��`��#��D�xL��"Oh0c���:
�P�A���4�{�"Of��q�Ѷ*��1B�)�T��u"O,ѥ��:e���A�E�]Δ1�"O<�t�(��Ȓ����R�"O�"]�{ݜ�)g�K�2��Y�C"OPX�3��K3�%H�j�~N��a�"Oژa�F��W/����Z 2D�"O.�(�	�7x�̡��!mQ��"OL\��'A7u>hX��Y�h�h$"O����K��^`�A���;��qɇ"O���X�j>����R7y�]k�"OL���D� xZ��i�:���"O�`vA�6^$f ��t.�@%"O܋F�ܨo�
th�e�h	Y"OT�)���o��y��7g��6,2D��+6&�DP�(Q�k�d=�b�1D���	4I�\��"`���-D�XR�$(a��Y�'�41IW�?D���쉺l9
i�& ō'^��
")8D��s�ՖUo� �'	� �0�� D�`�'��Af��GAL&J���@r�*D��[q��Nk���I���q�&D����� ]0�qr/�=Rx�i6F$D��B�c�P� �{�;"�F��!D���%@F�NS^pK`#��E*4'?D�� h��l�6#`aC%��`��(P�"O ��0�V�3��`��&��Uܾ�"O1��þU˾=��X�s��l:"O�ܲ��81 ��J�I�F�aQ"O���""B1!���#��
4�:�Z�"O� 2�   ��   �  g    �  B*  �5  A  cL  (U  \  �g  �n  u  w{    �  S�  ϔ  4�  ��  ͧ  �  Q�  ��  ��  �  X�  ��  ��  ��  @�  ��  r�  ��  � � � 8 |" R'  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	��BE��Nx��T�q��RS^���h!4D�,����3�J�2�%��dj�p/]\�<�a���j=ɩE��?v���.�L�<I�C21Z.ݛW,:?��@�1ʎ@�<Qp���P��-�ŀ�>�8�r~�<�"m��+�f�s�j�
P�Pb�Q|�<����&b���F+x�*��`y�)ʧu��E��#Z88T����d]����d�2Y��)�1r�qT��#x��\$���	�>�j�a��K�)а,X� &���$>}R2ONx�U,܃8� �dj�>j8E�v"O�QXP��D�L؃��[�C���
�'wў��a��-ʞ�%����̵Y0I?D��[�ÿx�Ix��A�� 
�>D�lXCMM�~JL���\�p�H	O D� �@J�%y�⍠��_�~\�GO)T���7J�,��p���;'d5����'��z�J��Q�3�B�u�΄3vԓ(�(��ȓg�]+�ɭd�s3~.�<��X$T���,^�s�$q��"E7lp���I���?�U�j'�L���K��\h�jEr�<Q�mN�R4�i2����w���NVI�<�2˔����� ��CF�F?!	��e���Z���R��M6�߶-t���=��n:�k�e��r"@́�"	�W������M��a��Tw���'+В%ȸ�ò�	s�<9��Lz@@�$E�1����u��n8�|Gz�Ō������b��*bL�(N^��y��65 �7�� �A�#M��yNX*�鰆�<��-��@��y"!�چ4�%¦~��ͻ�ꟊ�p?ن�Ot1�2#M)�,�.��R~()1"On���X
I%X�&B+pW�1!���g�?mڶ��:�u�p��������-�O.�	(Q�xy�t@� >}�UȦ�ü��TP����­B�]��t;�%�^��1 PM�����S���O�j< ���&W'|} �KT%δaJ��� �ؖ�ɚS�9�s��_���2LO�œ��Z�T�U�S�-��T��"O~��~*�9��e�$Q�R�|���L�Tx�E��Aߡ~D����C�:���?�A�(z^��@�ؼg��9jnQ�i4b���	�g��P"�S�����O�k��O`�'���!ҧc�F�0eܵ6�>@P3��, �Z��<I�4�0=���,���s�E:{w䤙����\�qO?ј��J�z��2¢�{~9	�A�I��	�<��E2Rذ�#�W�jX� Yh�<q5��M����b�
??ɼe����c�'M\���䵟��']F|���C�JX�3�;�f}�ȓH����]�)���圁z�R��'��v�)ҧA6�����^m
ę�ɝ2(�n����T�����Wv� 	+�L�Ê��s�kwI�<e����ްo[`|;&�;���Ʌu�t[b���k[��0���\B�Ir؟a3�,{���	���bQĳ)2ʓ�hO�9R�aRtm����6��

5�B�IL$�p�"�O!*)�µ��`x�B�Ih�8�SJ{ `���nC��6��-�c 6^�EH E��<U�C�~ ��7��Ŧ1SKٔ*���$)?�w�� �ƸJ0
3>��`�Qq�<���l�f�r%T��H%��CS<���X���J��$_8�b��K"Q8��,�����_hd�楝rVu��v�'m��zeE��j�i%,� @�my�'J��@�� ���8�KZ�Bޥ��'&(91O��%��`���31d  X�'��#�Α�{���������@��'�"��ͳ&��Eg���⬡�'����#8u��j�ϣF���
�'�R���!N),)!�*��Q�41�'��As�7L��<��M
�=+�'�
�;G���M_�<"�큂q�&͢�'z\*q B"-]�ؠ1GF�hPJYi�'���e� �Xw"��s�1c�6�`�'x��9q��f��D�kYj�	�'�T�s��s�"9�BeǫU�3
�'V���S�V Ǫɒť[�D"�X�'��I�H�Eͨd ��(��{�'��0j�
8"r�D��(�<"�.���'VV��"�ƸZv���`	9`\��'��8HE�[�!�z���JC�P��'���q��X�?NLiBጌ X�1	�'$Ԣ��F�H��q.���ⴱ�'�(��߅n9|��~ 8͒	�'(�Z#�L&74���
'HD1	�'��1���CB�����L�����'�"	@��F�>�T�����D�v���'����B�t���I��}:�'��aZ�c�/
�Vy�����'J�)��N�Z�=` QG�\�"�'�XpC�OM;|�����
�I���
�'������g�����3v\R�'������00WfA/$(ȝ�'��� K� 6Z`�&o�����'���0蒃x�b!�6-� A�T�H�'G.RCM^�4!r�8�8=��$��'(�)�-V����nݬ:x|��
�'�D�ѣЦ&6���L�]_�L�
�'
4$y��F�ڥ��"�TJ�q�	�'򪌉Ą��E�2��Go�K��	����  6�œb
$yq �v�l-��"OBp�S·�q� �P���r����"O�a���5\��&�:7��p�"Op�3g�����U���"O�J��A�:�!e�H�!��6�'��'R�'���'��'���'���&ذ����❂�:e���'a�'r�'���'�R�'���'�Ia�!���x1G�)�^�s��'R�'��'�B�'���'�r�'"�yc�Y
T-��P��)I����'q��'d��'K��'g��'q��'3N� ���8��`�A-H&X;���'��'�R�'���'���'{��'��h����ZP����mĸ"]����'B�'�"�'c�'\R�'NR�' *��V��!
�<��0��	�:�:��'1R�'���'P��'���'���'W�a���S�h;|����,��S�'�b�'0"�'R�'-��'���'�d}�cۣV/��"@$E(;j��`�'�"�'���'��'�"�'`��'���ۅDbIb�K[��|��'W��'�"�'�"�'t��'���'YY�󌈬d,�gh�+�T!���'���'�r�'�R�'$�'��'���SD��%T$5Ӫ�6
�vtC��'���'�b�'���'��'�B�'��AK��T�,� zvdX�s�"m���'v��'<R�'�2�'��Ox�`���OhyjCD�7�@uI�e�$!D�f��gy��'��)�3?a��i���#B��1�~���)�O28� �[���D���9�?��<��'?��:r*�>p�fU�p�
�"�����?q��MK�O��� ��J?�����s�f��4rDl�e-�I��h�'c�>� r"J�z0[�HF<:��<3 ��M�fE�@̓��O?X6=��T9T�U�J�.���S�7q�U�$F�O��Dp�\ק�O岙�i��d�q0ɻ�e��'��0 G��>N�r�lp��pv�=�'�?!��9!f��[fg�D|r�F���<*O�O"�lڶji�b�2�A6$�1Sd"E�o,dqC��`���I�0�	�<�O|�;�HM�D�)H�F&#�����	�c��Z
1�)c�
�ϟl����2���̬G[�Y:�ŎFy�V�\�)��<q���wH�#�ᇕ�.5��E��<2�i4t���O|�m�P��|j�'� M���UKݵ/�H��䢝�<���?Q��!���2ݴ���h>�`�' ����`Q��G���f	�;�$�<ͧ�?)���?1���?��ʉ<&E
8�4���BT�1;��B������u�u�Yɟ��	П|&?�	�o@�U�&*�+E�	�IB$?ٖ@��O��D�O*�O1�bL;7�=A���S��~qD���k6��C��������'�"(�B�Ity���7-���C�iֶV�9p���z��'�R�'t�O���%�Mc6H�?����?�V�9PA�'((��r���<��i�Od �'T��'�j^8lr�H�O։KF� �`��:
ڦ\!E�iH�	Z�(�G�O4q�Z���`V4qQ�D��<l���ܜ^�d�Or�$�O��$�O>�D!�Ӻ)b2��f�L����3�At�̡��ڟ(�I��M+A�ٹ��$FɦA$�$��
U?�L�_��Z�^`�	ɟ��i>9#��DǦ��'�����L/Wа���dO�fi@�]�u�������4�2���O�䉤?��G�R/,����S��Kt��D�O�;P��O�[���'�bR>ŋ��G?bV��RP�T�9��!k�F-?R���I��'��'(�9���0RPJ��q�\�x:�Պ���4ݺ�[�j~�Ob�e�I)T1�'!�`i���Zzx.�� �P���'���'�����O����M�J��{���[�[|:2Y��G��9l�/O
@lL��z:����x@b��<����K&=�*x�@j������U4lle~Zw�Ѩ��O�*X�'B��@���CF���T7|PZ�'��Iԟ��	ן��	֟��I@��`��P��E��H��cg`@�'n�8o]n7��S����O��� �9O$�lz�I2q�K>y�L�ХRe��=�R
�̟d��M�)��X7�yoZ�<q��I2�&Ah㮗 4���f��<�0j�>�p��L0�䓼�?=���*{���y�Bٻo�����k,O��nڡL{���'B��O�&Ch��3ˍ�a����޺�O�x�'�2�'��'��2W��M�����F��U2�OL���"P&0�tB)�Ɂ��?�tb�Oh�P��Ѳy$�E�
T-L��P!�O<���O��d�ON�}���b��B�Á��:U��S r:�B�hy��i�)
��'Ӑ6M;�i�eS�X�,=.��G���,xt(s�$�I����:sE<)nZQ~2넲,��[��z6h�3s�$��'.æe�p@�M>�/O�	�O��D�O���O�	��M�4x�|�@]/�����ƪ<���i�����'Q2�'K��y�%#��  �C�	���У��%����?����S�'+5��!������gY� `��R����'��2 �����5�|BX�� d�ݟ ���"��(e⍺4	ş$���,�	��STy��q������O��2܊e�.I2F��!	�N�%��O8lg�v+�	���۟��Ŋ�=.�L�3bM�6�L�G#6��)n�I~"�\�b���~�'ֿ� ޡr���;C�fW&� C��y�<ON��D�L|�$��J�_cv��!N�F�>���O��D��eaM3Ĳii�'z4�I�T::�����2+.�Ä�|�'��O<�e���i8��M:R���nQo~�:#�A+`��kՁ��[���9�$�<a��?���?�2�[�X}h����e��T�e���?����Ȧy��������Oh��q�́���J�lַH�Ѣ�O���'(��'�ɧ��B%
u&�[5煜l�Y�r�б{=*T"R��`N�șf���s�@�'�l4&��F��1r�Y��{9�(�f�����̟��	՟b>��'��7]�8�y@1��&ZD\�2�^�!`�#l�O���[����?yq]�@�	�$t"��w���wV\9��Y�,�������DK�æ=�uר��vQ�d�Y`yrC��u���S��?1(���%O��y�Y�����t�I��H�	ٟ`�O�:�j'ٴ/���s�ˍ�M�.D��(k���H�E�Ox�D�O����$NϦ�	-1��ւ@	=�`$Z�OǞd<���ꟴ$�b>�(�f���	�º�Q#͇�.��"l��Γ5� �qኲ�$�������'�^��2@�T��q��@;P�\{`�'3�'�T��1޴�������?i�C
5��S�p��Bn�c2rIЉb�>����?�J>��Wl�����ӌFX�YP����� �G�i�1����'��A-kR�g/i�|$���N R�'^��'����ʟ���	|�ʅa�x�q䪔ϟH�ڴ	W\H�(O��mZV�Ӽ�q�,p��ΗnU���fe�<����?���U2ySݴ��d[P��]���N$�둉ȳ:	|E
���k�:�`vl"�$�<ͧ�?���?����?�CM�iy���#�4V�y�gA(��Uަ1	����|�����'?�	?F�\��rJ�A� �!E��U'10�OH��O��O1�&q���>n琉�"�ŃfN�l���N�.�,�f�<��>2ϴ�����䓰��	^�{�%���V�hF�ߣ j��d�O����O��4��ʓZj�6hΎ5��ğI���B!�܋t��c�+
=K��n� �h�O����O��M�,�A�W��mCF�:r�B=���c�6�蔹{֠?�'�CҪQ7M�T� �L�t�4��%`�<���?���?����?��t�i�M�GF�{��%[�
���'h"�cӒ� A�<��i��'■� �
�E��e�
S������|��'��O�
��s�it�ɸ%:�8�)C�5�4�1CAیr���C��N�Y�	Iy�Oz"�'m�ɋ�cR�eC`(��c� MC�	�?���'���2�M��쐱�?����?�,�|!�sI^1Ԅ�:L�
+������8�O����O��O�S5ENhuH��O1\�Vt�UGA#@ ]SD���J���µLUEy�O.��I0U\�'�$���!r. i���ݔx3�M�&�'3��'t��Oi��(�M��&�M��!ӹA�^p�"hŹmy�e"��?�s�iV�O5�'{�)�4J�|�g�3;�X�˶Ï0c9R�'��8��iX�i��'���?��6W�0��(?�nh��) �]kzIpEgx���'���'*��'<R�'4�:����@��u� @_D����e�im�mY��'R�'��O�'r��΀�Z�2�.n�t��@Ɍ����O�O1���$y�<�	��dh��\3Y�&H"^�~&:�ɆVS�u�%�'+�%�d�'A��'?.�2�@��e̤��br�Yd�'\R�'p�R�8�ڴxJJY���?���>��e�f�̈́����1�ܻDJ�艋��>����?�I>a���&:����߄Fn��wk�z~�[�	+B0{��V�5��O9F,�ɨ5���үB�H<��Q�k�BmQ7̉ ���'Y��'����Tb7����Ā�B��D����4siBT;���?)c�i9�O��ȧ&.�с��1��pv�"���Oj��O��!��d�^�t6����៎�p�_)B�l��"k�j�J0�V��䓍�4���$�O���O�� �|d*�z2a�+P�� j±t4ʓx��L��P��'����'��,�"�X�3,.����3I>:,�P��>a��?�I>�|���ɏb���{�	{�z ���8\�B��^~r/�+T6r��ɿ=n�'5�	�bjv1���Y2HS gԣg�t�	������X�i>u�'՜6�B~���� V��)cU��.
���  ��;����]�?A�\�h�I�����
>:��:T�Ӿm������%B�ցە���}�'�5Z����?��}z��:�̃���v&���'�c�dϓ�?���?���?9���OK�}��dK1y����"�0T=���'L��'y�6MD����O�lZ_�	5�:A�$��x��`A'�޲���$����ڟ� a �lx~Zw�:�@�[���6�()D(���
Sˊ\��Ky2�'��'$L�4��児(�d���>>W"�'M���M�I&�?A���?�)�� �>6�Z'bƵ+�8c4��ts�O���OؓO��<N�Vl�`��0� ��s�R�\Dv��oE9w��H���|��.�O4E�M>�l@)$�0h�v�_="B�k�Ě��?���?i��?�|�+Ob9n�l��BH�� ��Yp%OƱg/�p��{y��pӚ�lp�O8���+Nc�x��d����1GR� 
����O��Tjh���Ӻ�����1G�<� P�AS�a��䀔�R3���9O>˓�?Q���?���?����	�:9,��0@�j�'i���nZ�-��	⟬�	f�S�@�����0�\�:�X��GIW���`/"�?�����S�'I}�Jݴ�yr�L�6���t�ׇ���镤@��y���;Nj|q�����4����ߴu�1�p�يo]$I@ˈ�YȮ�$�O����O�ʓițZ;.J��'����2�8	Q�$-<I�ONq��O`�'�R�$Y�.�;�'N�Sd� @�BR�O{�	�p��`�䏎L��&?A��'��!��7�:x²�>���=m��E9�.�O���O�$�O��}λ/$4�A�D���]P"��!F�8�?q�ipCZ��r�4���yGa˷f��[R�J�!�6���i��y�'��	�]l�nS~"lS�X�����f+����"V�x	��X�=i �|�Y���IşD�I�`��֟d�"'O��%sD��a*���%^cy��d������O���O���D�`������D�f���R
C�(�'o2�'�ɧ�O��!����$QތD(<����%�s�d�O��V-	��?�4� ��<��;R�����[.i��ɢ�P��?���?y���?�'��WѦ���O͟��sG�"C|(���B��px�k�xr�4��'n���?���?���	-�<|z��]<&����7>~���4��$^ߎ$c�O��OR�*ϖI�h���7%V��R1�yB�'s�1�Q�L�b��oN(Z�P�e�'���'�n6��'�����MKM>yr��/-z� �
;-��}J]��4%�h�Iʟ�ӥ0�`lZ[~��+_��H ���y �X��PN L�q��E?IK>�-O����O����ONm��O��.a�ő���.}��� ��O��d�<��i9�0���'���'H�:?٪0��'?~����`�8�����ٟ �	A�)��[�k��řFh[�;�8a0�	�.\�5{��	�M��O�i���~b�|��#���Cۻm��1A@&6���'��'��T[����4[)��D��r���Ȃ3�l�3u�����S����?q�_��I�U�~D���22���m�;u|��I՟iD��ͦ��'W,c����?U����C�̘�b�&)���=ܢٙ�0O�˓�?����?a��?!���	��1��I-m�Y��l��1mڝpN8�'+R��ڦ��#LS���D�"^1
��K�K���ş�$�b>�#�g@֦	�=i6D#UO�!u5������9�,�S�T�G��O�q�K>�/O���OF`�ӫ� �vd��X<B<ڵ�o�O �d�O��<�r�i�]���'���'�bl ��7H�q���������}�'�R�|��P�#�$aR��+&��0#Y����IV�����V�^ē�����^V��_��`œ!e3(1����`�$kDP��O����O^��<�'�?��g1�:��݉f)z���oG��?�Q�i*��2�\����4���y�&��^q�XSЭX 0t�HR�O�y�'}"�'X|Jñi<�i݅Iŏ�?��U�K,.f���C$�r����
���'��I��ğL��ğ��J�Ãt�Np�SN��L��}�'X7��8X����O��(��|L�s啑	�:`E�5�쒮OL��O��O1�d������qT��Q�`�4�'�C�Y؈KW��<a� ���h�d\5����M1UְP4F܏T��J��W5+���$�O��D�O:�4���Ǜ��jn�ī_*ܭ���zj��&a̱P��x��⟄p�O�D�O����h�"��j�2Ų-�&�^%Pp!2�r�T�zA��uO:ʧݿK7�΢e��y���'e0�c��<Q��?���?���?A��T%�%;�l;�oL�-¬��J&2V��'�RIrӔ�U6�6�dAҦA&�<p���%�8�
l�\�Ht;2��A�	�t�i>���k���'�-����2[�,xSC��(\/~P� i�*"��=�	55��'��i>M�	��|�ɔ7�R9��G�#�,����<[��	ߟ�'�z6-�!_��ʓ�?y-�f�gn�tG�Ah�ٽ���xr���ЩO�d�O��O���DBN�D���cP!��(ۊ{O\Hd焝C��,��&%?�'<�H�dL����� p��J,&�D�0" в;���k��?����?	�Ş���	馽��˃�=�E�,��U0��q�	ܵJ�>�����
�4��'FV��?!0�ƭ������ʌR@����?	��d����޴���>P�Ƭ��O>�I�Ѳ�+;�0�i$Z��my"�'s�'��'�T>=�GD2ܖ4��!1�
� �B�M7L���?��?YJ~�[>��wj�]����)���GF�~��';Ғ|���ʑ�w��7OK�9�^��q(��}|E��e׊�y�镌��9Ԇ�1(�y9$`@���}ɂO��Iq����#��I.^�ya����mѫFK���­.S��8(�LZ����F 8�^�s�Hƒ �J"=��dR�*q*ԣ��ҭ~4��DQyB��2J�\��`��8H� ᔉ��y\b���KJ2_��j�
�7X�� cK�Io�A� ��Q�(�����<:��	0^B �&� (��L�}pᠣ��}���32T�	�c��u���o]4v��M�D\6�T��Ĩ_��:���*=8e(&o��M����?I� N�~�.�*푖����pJ�.~���'f�'��'��u*�}򧃈aRX(`p�J�9q��Un��Mk��?�/OfE3�Ap��'�2�O�� x���#�� ���y��&g�B�3��x��'�R�F��O���9,G`����
2h{�+f��Q=�7ͨ<�5�1!d���'B��'����>�17�\5E��9̸�[æF;� o�러�I�W����?���4e�|��W�ͷ��(Da��M�'b��/���'.��'��tI�>Y)O
�RM4]-{#�؉ ����
��3@b����Of�za#�ͮO}=���J��AB!MӰ�$�O���d)4��'|�IП���l��˱J�05�4�s#&��p��>���V?���?���?�so iP��U�
2,�|݉&��f�6�'�<<H��>A.O��d6������c͟)+b�x�A߁G���k�X��se�̟��'F��'i�^�j���{o,yr%��86n�3���
�Xݪ�Oʓ�?�,O��O��$O0C�L���'�ta2�@$Z`T� ׭4���O ���O>�{Jڅb3�z��eK؞Yl	H@��T�0=��i��	�(&���I�$@��To?9&(^�F���bH�b���ѓo�Q}r�'|��'�ɉ>u I��,�^Ģ��Tj36ɔ� ��αO���lԟ '�T�Iԟ�:BǜSܓE�8ٓ�Áh���X��.!��$lZ̟���yy�J�4G���?)���
ᄆ�R���7�ݺOȘ���ÉK$�'
��'��hJ����?�C���89:���"V���b��`��l>�����iC��';��Oٔ��ˢ��
>zy�e���Ý-�F�'�B�R�/y�O(�>�+&�5O��pb��

��s3�|�Dui�)���u��ß����?E �Oʓ)����g�	"�nL 1�S�$���Bǿi���1�$<���X�M��^�6�BL�	���*���M3��?1��X���^���'0�O�(����f��F!��/[�7�d��l�����	w?Q���#���VFȄI}��`N˦����I���'�X꧋�'�K3d��g�q(�h@;��4ؤ�#��?	�1O��Ĩ<��� 4�^��4��nG�j*j]��J���$�O��"�	�D��<����FW1?����L֫u���n�� c���	iy��'�(9¤ԟ�j��+ �i������t	йiw�'5�O����<�'�ߦ�s��I�BK8�[%�Q�{3��E�/��O��?pꐪ����O�=) �K�`~��+CD�Qy��1�Sئq�?������.��'��d�C�B�pD����O��{�`=�ڴ�?I.O>��ȚPx0�'�?�����1UiJ���@ͰY�����@�l
Ό$�x��ty�e� �O�NW�%r���cH(Q�谁k�� ���ܟ��a�ݟ��Iɟ����?ٕ�uǋ( �Y5��%q_�M�	�M���Mw��Ҽ�Cg�O���t���f𙃻i�T����w�L��O��d矪�&��:u|���,ָT���b�Lƞ2�L�1ݴ�?a��?����D�|�+�6y:U�����cf��%�D]�%hYЦ���ڟ,��*�)���i=}2��q��U�3)Ԝ5t� ��A<j�0"<q��)�O`�Ɉ^mv���9:�N�í�!x�H6��O\TǴ<�ER?�?a���c׸E*q�^�S͢��"�p�'Xd���O����O����<���5eb����-�!(�/Ɵ��td�xb�'P�'�����D��$�"�JQ�: j�<���I$+�0�oZϟԖ'L��'y�IٟP5�_F���E?�@@����3fԂ5�����Ք'��OB��<�[pLoZ�u�XpU�γ0Q&!�fC�$�h��?y���?.O���&d�1�xli��G�t����
��I�4�?���d�O6ʧ�?!)�24���"=``�I�41�% q�Ʀ)�Iџ�'�!Y�`1�I�O����lX��c�f49`���	�����i��I�D�	����IJ�4Q��؝P�96
3�R}b���T��7ͽ<ArgT�h��6N�~:��ʁ��@���`6�� �]Y��y	��w��$�O����O��&>�Ih�ܴ%���E@K2Ȑ{��ޯEkb�nZ R���ڴ�?���?��'Q���\c+R�b�G
�c�����N��Ԃܴ�?I��?�����|��?���[�_k4�P,Ot�sC��R��^A���'� S�+\
듊���O���.a��F�|�84�d�lx	�O:ʓ�����'��'` �����u�$��(qǐ�`r�yӜ�ٿ/���'��IꟄ�'�ZcK�E��*X96�u���Ǵb��er�O^]A@��`�	�\�IڟH�'��tB�	/���e��(z>��ɒ�S�`�����O�ʓ�?����?�4��*#�>���`�"O�ֈ��)�(����'���'R�'��-8FC�O�b=*���F�ޘ4�H!�ش����O���?���?����<	T��%+�� ֧ �z T���I����	ßؔ'� 5)"l�~���+��P�T�}zdђ��# �y�c�i��S���ߟ���'|�h�	P��4qoTu�Qc��z\ڔ3�[�� o��� �	[yb@�)7B<꧳?�����!A�j:	� d�c�d�3K�eQ�	ş��ݟ8@��u�X��y�ܟH�җ�Ѷ��V��gN*}���i��>�
�iڴ�?���?��'KN�i�]A�-���x�喻s�"-P�fӪ�$�O&��&:O���O���i�R1�8RJc;ʤqb(G�A��։ێ'�L7��O��D�O��	Ci}�T�p�	� T�2#�"4����#�T�&���i�N�K�'�'P��Ì#��F�{��$K����{U�mZܟ���ڟ�7�J ����<���~2�[�&����'q�����B�M#����[�-+�?��I�D�	 ������\�"1�Բ1U���ߴ�?�F�('��jyr�'C����$9��,٦�S�({PD�$6w ��y3�Y͓�?	���?���?!*OH���5�6)��L�Bt^m�Hȳ%��\�'n��ȟ0�'o��'"�DMK�D�#�hw��@2�X4w�u	�'��IΟ��I���' T$z�	|>��+�28~�t�W�&����d�l��?y(On�$�O��D�c[�$V�r/4��;�y�W��'N�HL�'�b�'&RR��+�Bژ����O4q!H]���0�!vh�Bt��-�IXy"�'���'�z9�ȟ����j#t��1�C��!��Lٲje���D�O��IƄP[�[?�������]�ބ�F!�?�~1ە��"с�O����Oj���Th�D�O�˓���&�>�"����y� �1o�M�/O����ΦY������I�?]©O�
���S͉�=��B�M�1��'B䕼�yR�|���Y�bd`A5�Aظ�%N�z��/� 6m�Oj�$�O8���D}�[��#�ݍT�1��G�X0�Q���M�r��<���&��џ�y�#@ތ�q�^ ċ�@#�M���?���H�����[� �'�r�OJ��v!,.>��6�֓$5� {&�i��'�j�����	�ON�d�O�]F돗g� �����;_h�m�,æ��	4��bO<����?1M>�1~��eI9<����k
@��'<8� �'U�՟���P�';�ؑ�9!F�-hJ(,�2�����D�O��O��d�Oĉ32��uq�(����p�3V��<	��?Y���Hр0�'n\��T`4rud|1�>C`��'2�'��'"�'$ty �'�� ���	H���HV&�c��w˳>����?����D��c��%>�+6
� Nf� 5%� dd�95��6�M����?�;l�J����	��y����Pɀ��B��+��7m�O���<qFʞ	щOPb�O��2�`݋$O�c��A�*�<V�8���?��GINup��������.T��\���z@������M�-O��g�����9����D퟼��'$���r���2���E,��o��?���q�Y �����O�ִZG@����@N��p���i�L��5�k�R�D�O$���V}�>I��9d�FD(���98�* �d �"؛��߇�R�|��)�O��]�mÂ{ԆP4B� !V�����	��ɘ:jێ}"�'��$W�[e���`��pB�Sɛ�|�)���yʟz���O:��V���`g��ɲ7��H��n���["O��ē�?��������D�F���0��"�p}���MB}��h��[���I�L�	oyB&�2���fJ&u *I�kY�X\�Q"�D1�Iϟp%���	ϟ|�q�W�n�e��ɼE4!z�!��4h4M�Igy��'���'��	�5C�Q�O���WĎ7Td~�ЂD�M�J��O��$�O`�O���O�[�ONܻ�o�)]7���f�dLU�p^}��'���'q�	�u�.�9J|*u��$<$�0�"f�S���Wi�Qt���'F�'���'�8��s�'��8>�a0�G��a+����"��8o�����SyrAA�<6���柈a�e��%#0�S�Z"���I��o���� ���6�$�	g�Y���0$�M���ſ+t����Ֆ'1�p� �k�Vy�O���OZ��;�R�5�9~DB!*!��Z�oꟸ�I�TԒ��IJ�	hܧfF:t!�g�_򭙄I��i��o%�4��4�?Y��?A��23������=<6L�n^;x���C2^C��?����'*6�CbP_�P��$ꚱED��� �j�����OL���C�Y%���I�� �I@d��$%�&���0���� ���I�}�j�'rr�'6"䒚u����%���ZL���.�1B�7��OD�HE�\i���������5�э8�ECǊJ<>~EA�c�+��$��y8qO
t���" �0�w�7�4FU+o�����t�HP	 �g�<�G�Ay8�h��O�|�z1w��i�'fx�'�b���֓t,Њ��2JvL��D,J`BXpta5�<����	Pd,p�E�� M~ ���&�,aA:f��1�g	3MV�cb��q����R��|;IF�2�5`Γ�@n�xJ�숽z�Jd��a]$
���n��[ :\8�@&�14���j7 =Tr��R��S��d(N�<~Ӱ�%*Wܟ8�Iޟ�cŋU'g�2}�Q�Ԋc�\Ο�I���G�FLd5����V�N����~�Q���dꊷql���SEU�`��T"J�IҘ|�$�-#�(*�.+-a����d�g�Q�|a6.�O��d#§C7>%���hT<z��G�k҆�r��� �!�_s����J�0Y��9�ť4�Ox4%���E���)b墀9�r��1t�Hŭآ����O�'G����?��X���P�(ٳN�:!�G'�,�,E��N����W!���S����'�py`B*v��3f$�;BC� �s
ˌ=��c6°E'�9֧����6`�~(P�O�(���@�-��l6�'�򛟒��O�}pF�rp��3�׸|��"O� 
!��k��0R��q�\Y+��I��HO�Sw��(2f$X��x(V��ל��Iß�8GO�%W�����ß��ʟ|(Zw���'�L!G�_�TNH��EGyn�X;�'��M遄\��z��6,O���g9_miX��A�q�P0��'�)#���
3j���g�5OlɸEjP���-��!��OT�( �'�B�|yb��p���q�"�x8ŒD��y�/I�r��8:��_�Ϯ��@�-hl#=�O���*Mi"�K޴!�pd�c
�B��MY�cu�a���?���?y�I�?������T���`A
%^���"M"/n���I>�4��
"lO�hq%
����xF,V�-tժ�M�4�{UA���a���3r�d���OY@mߤI�(|o��1��7ړ��O>�y�&�K#8�xc�T^:4��"Oz��TJL868�SC�3M �
�>O^	�'��	�eƠ��O��$�|Z�.�4>n
���?��M��a	�"Lk���?��bLH0R��ϼB$�"�>�OڞAӱ_�!?^�*�� \D�y؎�W�W�@��@�S^�a�}�r@��$^D9�^:J�
Q�y�'�8�����?���$�2<9�d�L�n�E����y�'����Gm\�%q8@!B��13�O��'�2e�G7b2��UFƉd����Q)q�����S�Mc��?Y.�8�$��O`�d�O���L#I�>�����#�.(���;,�,��3�|Fx�`ޱ�(�D�-�8=X� �2*h����)��4@�Ԙ y�0��O-~6�����K�7�@���q�S��?� �#@)>��5@A+4�p�֩�j�<��o
 A^���� ؽw����"�^�')�#=�O��K$�������D�KV����';rN���ܹd�'�"�'��$t�)�i�)[��KȞ����E�gGVD�(� CJ�dx�L0�oR9W �<h�M�;{C0���
�<i��E�6�8<3��O1^��LD��S'����uK��o�4��a@$x©J�]�"�'96ݟ������'���
��;���r���4�(��	�'��-ٱ J�~:`��S4+�����y��MmZ_y��)�<	��Ċs���o��l�;A�,iBjX����r�'"�'S����'��6���A���%7���J ��u�#��_���KK��p>!�-4p�ɓQ�����ǲ?	d�C��4ɺ��$�O'�'���IDn�6E#�&�.<ʾ�3��|��'����?!z�˄�d��
u$�kv�dq�� D�PajX�))�Ɂ�Ꮋ�� �f�i��b�OR˓F�x!�պiqR�'��= �����������Ƥ\�H�v�	ܟ��I��BQ�x�K>�O@��%�N4uW�4�ǃ5��A��D��s2NA�i ҧ\�������hZPSw��(&J FyB�dA��?����?�*�$��S݄MӢ�H�I%�@��A�O��"~�p[|��O�f��3r"Q8Q�ņ�I.�ēH��P{�^;�U��	7'���̓p&I�S�p��q�D܍JhB�'�r$�=��\�w�S�B�
���͸W�-y�Am)�5if���,��T>�|��$v�Єq�ȶ?c�4؁Rk �H���P����0�-��]��S��?�4�Շ'""�cD��&�z��R�J�Z}x��?��O�O�'g�4#�o_�OǋFX��*�!w�<��"7�9�g!U5��GGK�'�#=�O֨���K�4˂��"��
��Q��O.�K Mԑ=�С��	��T�H�"Oh(y��ʥ:6��o�)
�|�c"O�)�!CB0�L��C�ܸi���c"OȀ 3���H�hw-�x�kA"O��$��2�������`��Ka"O�0�,��5�ڼ3�2e��4�c"O�Z���V�FD��.��W�����"O���FA*=kD�~�c�"O�+����n��\ˑ"�iˎA��"O�}0���h�mK�����U�3"O�Y��6W��1�OT��:�y�"O.��2,ݘ_u�<��Z�\e��	@"ON� ��_9*��J�
ɕ)Y���7"OB��D�.kl�,MU��#"O�yB��*(��ʢφ�!�
��"O�4r$��)׮����.:�D�x�"O� �@�˗(q�yX2A�_�� `"O	�4�L-a�<D�#�R%~��p�"O������3 ��Y�� �^E@�*Or!;�� 8-�l�u��0'�I��'d��"��؅y���RBɃ'���'����JME>�J1�l�ļ�'��|(�ǩ0�
y�a��f;x���'�������(r���Z�ͥ���	�'�l ��eB�tAؼ(���z%�X�'��)1�gYF }�Шc�F@
�'z ���K&/�8mp%\2X���`�'GhI�[�"?�وG��1G�l��'����gN
&~4��	�����'$H9�#�(n����Z<4"&�2�'QB���߱,tT3 F ~B����'���W�C�
24K���z�T���'m0x�P'C�t� �&dQo�$��
�'�h ���E*9
)BA�W>��'7��#5a_�O&Y��m��L����'���l��v�y0���&$�\��'����W�u��ij��M'�$и�'�vKvL�8�h�va�!#e��i�')�U�k�1;Hp�ȥ�"ZJ�:
�'�~9q!A��Xr���P��ز�y���b)kd]�(2V\���Y�y" �+�h�3b�8�D����yr�_�:~��w��+MT��2�yҎ
?t������Q�j�Z5/���y��U�d���BR����&�p�^��yb(��'`��Ԫ�5r�{'��y��&Y�1��ݠ#�|�;# ��yb��>=�4�z���8�M03�E��yR$N;�����͑��U�2�X�y�õ(6�iX�N� w[��@�ؒ�y2��tB�;�&��j�����X?�y�9bTyk���7Ab��O��y�#XʂR��2���  �ybh""��u����������y���K�V�Q0�Q�u�&!�Vj�y2/��1o����λy[l�q�"�y�b@�Y;��ّ�_����;$H��y¦Y-�d��V��?J�x�#H6�yb��	;�rmqG��m,��9`�T��yB`՟K�x�C�Ib��ؒ��ٴ�y�I��?�d=�'ҹF=�[4��yr��+it�"#@ )�F��s�I��y"��&ب��7i̷r�mq�K�+�y��J�UI����)LW��)*�T�yR�!Z�	�/�T��dp�����O��퓋TЉg"^)9�0��� ��C�ɧf���隀T���7bȗQ��	;��?E��Ə#$��GEH�cL�U�ЍX��y���f�0	�Bc�,��9t�Ƿ����6���s�oX�Tɂ,�l�n���e�2DTjQI9�O*����Z6$i�t�6�(U�H�yb�	��	`t�^gH<�2k�{ݺ���MN00zD�wC\S�'�fl�e�K������!P�]LP�ˋr��!�+D�yFKj<a�`�Kּz��O�y��&,�q� h݋���-F���������� mR0C㉡�xeB��0u�@�{g�"A���o��y�f3o�C �B3>�p"?� A�2)5qVozA>]��k�Y��K5���:[��	����̉[�(�:Ṕq�̤{��0�⥉�~?����87~�M��Bx�ؠa��!D�����MA���'| ��D�,�b	��@|�lѲ�y���� �*<t�4�p��
7J��"O� �4�d��zV�H�,خB@���F_3Vlѩc�'Avh��y��H�D:��[���8i�S�ͣ�p?q��>b%��"��,��y1��h#��d+�{����&��"l/�x3���&(���'Sz�8��P�u�44A���+O��Ɏ�dZ�VG>����f(���p�ٽzY�;�<	6��W���Z�iL�K�*�A$ڳ �ʀz�ډ5�U���2�w�r�q�R;v~���ɨ-���;ٳ�K؎W�FjU�9
�F{RB��>~����Ȏ0j+��1�Z)��^?��?�`#� y|Tx&I��8̑	5ˬK��
��W��p<1C.�l3�.��7�����HJ�,;�F�ua~��OiĽ�'�� ��Y�0@-oz���cyF{@'^�� ��i�^�#��&�~�	r��j�X����OԬrm�$�?�Q�ݳ$ �0,& �b�8OrT�hS^�`ct$�	��t�EM4B~�@���O2ՂZ�T�A!�O�)1zaap�	m�4��ݧ`�h���ۅWG:��B(^`��|r蚖=|�\:�8��'/��G5D�x�J�H�ɵi��j�AzPKĨw��~�FZ8O�F��@��_5�P`�۟~촤��o5��T�'E����[ca<l�. \�Ρ�sHņW����&2lO����ɽx^�A��kM,60$ h�D���#�Εߦ���<.,�M��aK��\5Z���Bn\X��e�� ��8h�k�cɔ��4�VE,�	�{͢Th�@����e�N1�W,�>9s�S�(��G*0>*rSoTϟ���B�:$2 �J�wuF�:w�#�'7"Ȣ���s�Q���Ӻ�pv+�j|,�:���	q��5�'��Qf�A�2��UYe(�?d��3�!L1%�����O���`�j�&�PHV�����`�Xd�_cό]���ۜl�*wg̃S�vicՏ8lO�{tb�-,���ˁ^���F�ҝ%��03�ݟ$�
�D{�G3A���po~LL�C�/Y��~��s����a�$��hGR��d�jCB6I�> 3c��	��(�=�5�	2$K|�/8��EK�R^<n�3$Ȗ��[p4ja��4[$�y�c"�7�¨����'F�u��?n ��y'"���.x`��K'Y�a{R�W b is�O�0�* �ř"<e~""�5e��0�Lx�D��6`���.E��p>����T��A�c+��"�O��11��Y�FΙ5p���2-�bE��s�<�pd�J$\�n�uB[$t��怴dC�Dy2�!'n�qJKV�t����(F9<��(V�/AD�q�V�h̉'߂�X� �Q�P� ��bĈ�}B
�7M��@	�K0
����Hʧr��|� ��p9d���ܞ�}(C���aD�G�7rXތ:�J�^p*ND0=�x!��݈�=�v�N��F�뀌�e��9�7�N�*����v���s`�Cc�d�b%k�i��O����q^���4�<���2��G-t1+&@�-
����&EɲA�T�!����ǲY�]��@�_�F�s
�-�~-I��̕Xp��qdĮ{'���"�ְ0��>ūSc
ZDԡ���0��l�#�*��m��ɰ�iKpQ�&��M<1�`x��Wu2({���ȖlJ��On�1�+�O ��dنQ`z�����ˤ��g̓J�2�1����V��Q*��?L��"<��'x��0�P(����Ӽ
'�� i�k�*} >�ͩt�Z�@�����5@P����L,���I�+U���d��'�<6�� 0�q�}�牧u哊̛f�����,v�(4gC:wn$��F�C*ͅ�	�[I.���O�!���R"^��EhǊt��ѠF�X��$����	v�J���e�ݵd��81#V>Q!p��=Đ�`B|�\�i�&�8ݤ�SRH;�	�.R�(+�%��<a�
\�wI��ԟ�1�D�ֆw/���f�҇%� }���^��M�����X�����Z�)��T�Mo^��Ő�O˾@$�|:���G��Y�Bn�r�ۇ#�M�u�'P�$(�V�,�]��O��.O�v�!�` �>TS�¾yn1d�N�p��A�[e1��q�'�1��Z�
�0"'/ �.��0"��,ɺ4��2r�S�sӂ!�H���1� �Q#�2�9�Qn��E�Z@�4��I����$O4m�Ҍ7%��\�2&H=.6l|�����
�ɔ5I�Q�e�O��*�I���&�Hлi6��a�d$=��(�SNļn������T-D��?*~1OD��j�D����>��xH�JĎ
� ѯ��"ecܨ[�֡����)�"��9rvF���k:?Ih�p�4%�U;C�֘7��A�+���ԥOT	���Y�P��[���5Y8�paG� 8ڞ$;��U�N X����%Oa��Z5��T>Hӌ��Dpe{��Є:�`։\�tM(�[EO�g�L�5� ��ͻ7�gB+���`��1%�����#�35����y���`��_"O�+$5���h�?���c�T	#rt#>y����`�l��@=�\�(e�ƛfc��$�@�%��rE�C�?i�L�(�b�Y G����O"@Q����a�e��<V��<+v���i���`j�A;�QT�L)�`$��	�5ȟ2`��9�F�<%?]񖨛�/]���vD�'y���c�c�<I���1Q�б����I׼$��[���}�+h[8�!j��~�85�%"���8����C; ʓL^f�gyrC�<�oT)!�@���"y+���%f}�Ҝ��YÓ<�Q�.8}1�(���&���V���Br��o���*n4����']d��s� �X*C�H<)@X�'��;⒱�A�I9:ƚ�K�Q,�`���.j�,6m�j<�KA ȧx�r�@��܋IlF�٤�#�O*��@h�,o*`�sǼP0C\��[��Q���F��
�8�(;}ʟ��%@� ,:��ܴ@R���"O�	�5��/T�L���̊����2��0ӈ���}�FTH��i��b>���d:is� -\l�����ΡSD��^h!�"W�	DH3h`@�7�I�#�@����pӘ �g�>9� �I(C@X|�'<0��Q$��s9�$���0�B	Óbɔ��e. �d�i�Z�TA��V�Zp*]�a1�q�����đ���'~��j���3SYv�!Հ�,#᢭�H�̠Ǣ�]N�'NLd���D#F;��ɮO,�c�RS��C�Q�A*��"OD�!FΆ$X��QK���K.h�2�x�.ŉ{L�:a�
��O�L�x��p>�S�,�����������S�/D��p����olv
R ��)�����(c0�I��O�4�@YW�g�Ix��!c��ܽf<�uPc��BH�C�#7��0A!�w(�;/�bN�sp��+S��A;?�O�Ex6��m쒴��k4&��
e�'l������^ V�ےd�H`���=N!���{���#g)�@��J���!�O����V+#�R��R�GB�!��C�`4[� �2)#��:lv�!��.�.�(b�!0Q iK�e�!�d����z�)�[�TE`��ȱ<!�ܱ+�M��+A%'��@yQ��,U!򤈈p�^!I&CΓ$�hLrG �:<�!���m/��mC�~nԱQ�EK��!�d�~
�ek0d�Ak$��6��+�!��ȣ�����GQ9�;U-o�!�dԡl1ȼˆ�@�g,	�b��	6!�[O: hũ��Y*i)E�ڎ<K!���+c�
-�c���I�Ga�4&!��٭1غ�珣������!!�$J�-#�9*�hD�=��Udn�%m!�d�a~x��S/̸E��42��*Bf!�D�)�( vE��o���K�-�4}K!���6�jD#1�ͯ�f�8 ��FI!�$\�F�q��VO��+U�Ίr�!�dɔq�T�#L�E��CfS;�!���"�ΌP�"�q�蕣��K(O�!�d͏:�z7D�*r�X��ИX�!�d��R%h_k�k�M�'d��x
�'�b��j�b�����T�0�	�'L���S��*_|��{7��Y@�D��'����1����	1{��y�'��i���0�`(��kׅmGT�`�'D�Q������ƀ-_��#�'�V���i�m
4�%D�* pps�'�ʩ��E�lφ}!�K�;'V<�z�'�8�)���4@�=��I�NG�UK�'�B�'��P�|�1�g؅@b� �
�'�B��F�֑
��8�#P�Gbձ	�'q��R�
=4�����
M<����'Tޘ�&N z
�!�(S 2 F���' �]�G҃8ԝ3��z\��H�'@��A��%#�>���'d]"�'nD�8��S��� ��)a�(���'�,�z�I>i;ڠ�ւjZA)�'���Q�I4{F$"�H�iFv0"�',��HB�ݎB��18�iZ+
@�;�'�4Y�6���0e�1EIoJ�|��' P
�I�79r������f�}�'p)
0��Nʆ�4 Ɗe
���'zn�p���Pَ� t��5���0�'�Ty���A�)öŘ$D�!>S0�!��� �$�'%ģ�B8�r�J�OD�	��"O� @�)3ҙ�fĊY5vp�"OX@`���L���r�O#w8��"O�6� 3Wz��3&�O�ڀ{�"O(,A��	0K�!YeO6(��+B"O�H�!&�T��dQ�V0�C�"OJd���-i�l��-K8K�<W"Of ����F�V�l>I���"O*e���-����k@'?����"O,|F$Q>�x��f��U*4�g"O����ŗj�pkf��8���:�"O�p�Ԋ�F���i�Զ �1�A"OZ�Au.,�&F�,n���R"OPH���2����f��T�6�9�"O�� �'éC��qae�o�@m�q"OȖ{�IbR�) �i�Ͱ�yҍ
�ci@�9aI�'�6�� ܰ�y�-P��.��
V&�T���P��yR
B�+�J�@�eǝ%\)�d*D&�y�ƈ!o�|���ԋ5���y2a���d2��I�fE8F���y��M�e�z�D��u��y�̍54���/�wj��ѴLO��y2��bj���'prxj����y�eX�9��Ȳ�L?l��
���y�?�L @w��>4��#j��y�@ĵ8�nizSfA'I��cG#�y�:��Gk=�]����yBM�6c�`�B&�	/� ���y��2(^���!M�L�b�����y�i�:P<x��Z7�< �2�Q�y���k�ҀSc�ۦM,��$�A��yBV�*=�V5�-�D�n����ȓ,�r�:���3B�����씊^��a�ȓ>��@�E/FE��#���H���ȓ<����4�@��Uxߤ��G���� 	��!��s��K�F���KOv�В�GI�#嬈-w)�	��X��3#)��*hdb@�B��z����j1�����I�q�*z� y��"O*����{�,�'
��g研��"O
]�ɖ>G�	��(U߲DB "O<�c��XNh����<Ј�zV"O�ɩp�N�m�"�*�C�.q� ٙS"Om[�� _n���+>���13"O�D1V��20���*
�w�JL�A�i�ў"~nZ���=�E��j	�R�+[>B��>��2�
ϐ��%�Ҝ3dB�I�]�D��%/A�>�r��p.D�+C�I�E�p|��d��,r�1� 

5�B�	�f�(���S��$�3�?6�B�	h��-�%:fVXH@��AtB�I�%��q�ѧo�D�3 �*y��C�e$(��hJ���N:�nC�I�]��s�I(6u"�Ù7�DC�ɵ������6>&�+э��EpHB�I��m���v8>�1�Ɠ$�C�b��L9sA��D*0���KB�	<V!gE
�l�qs���'f��C�x  ��])M�k��B�X��C�I5`0�<X�.A.���#5�U=@�C�I)CF�%P�B!.k�;CFR}�B�3��|�2�ɔ'��}�񏏩y�B�*-�����!�2q��=�qiLG�TPG{��9O� ���̪mB��P!lTzZ(�"O�'ϋ� BDa�t�
�H��"O@��ai�"�L��i��-��##4�S��y2��f�����
M���d���y��9�:H8�Q,H���S�إ�y�̼���$��.<�N��c�Ԩ�y L�YVT��s��8dV�Ad�@��Py�D8g���Y�/$J�yՠCi�<�e�.8`�aG��g&���d#n�<�4��2b^r�˵\-��ɑ�i�<!#���
�+� �f,�%-K�<��l�1�*H�b�$xx���C}��)ҧ$<Z�i"ɆNM��	q�Ε�F	��N܂��DlW$�L�9Q+�{��݇ȓ]h0��9)F`Y�#A��Շ�z��n[���I%iگ
��P�ȓu?�8����s��`�晴:����s~������:��X�#1}�q�ȓ
�v���ݍ]�D<KDI .ר؅�"��,������޹��ǲ
;�ȓO0� ��M=U�� [��:*�i�ȓ>G�T��,N�Z̾`CǭK;ir�C����hǤQ�O�p�9�#�&!��B�	.)j��Ɛ
Ab2q�'Lܡv��B�ɀ�D���_/��h�T���.)�B�	%)��] �� j����u+Y�P��B�'	9Z��r�$s�DE��`�XR�B�ə�p5�K�!j�E�d�*�"<	���?u@�$�1=��ِ�Lз�j�"�N*D�욥�V9 ��A��P/?Vlðh)D��W�]
),�
U	\�"�R��;D�K��U�W�2� D��03�T�:D������'ZM�Pё�[�DȀzB�8D�ЫP�!&E��G@E�|Aa�<D�\8�NvV�x��?e`� f-?D�̈��N$�Ʉ�M�pLP��*D�8)�i�"n�:œ�
�  e���>D�@r` C�<�J`L_�@Z�4��<D�X�C)�Q6LmR�hI�D�I�J9D��c���l��l���x	l����)D��W�M�i)`�I�'u-si)D�<���E p8��2��Y��q��$D�8B"�>yG�HBr�T	%P�k2*$D�x6���	�� R�^�l�s#D�L�"BC�m�@�����LI�+D�����;^�:C$ɺnǺ�si*D�L��*@ ��}����d����U�)D�\'$W$�bjÿ[V����E%D��jB߼X|	{F�|���srL-D�|Z����J�rPQe�'�t2L(lO �p�F
�!d�Ȗo]�P,k%�8D�����̏-h`�3�,d˵L5��X����F�l`���І\���PF��e��C�ɮcޢx���7��y g	A��=��'=m� ���+M��·˵nc� �ȓO"jd�M�B���WN�]W���B��>2��O�� 3xІ��"�C��Z�"�ʱ�e锑a�J�ȓ%�h[fD�9'�ȼy�f^�7M�u���\��/8f�|��B�R�tm�ȓO���@�c�.��x%���1�����5��#.M=:sǫɚQ`�؆ȓ9kJ��V,��I�&<k� i��y��i	���ua·RSH-���֚
ZI��S�? n�"�.�Ajxs�^�K,���V"Oj��s���9{��
�L�^@�D"O�Eڃ$�=�|�\q����6M�I�<Y���5kU+@L1T+8`CCF�<Y�ٓO(�	�C)j�fs�M�<�a[ 81P�o�(T�
D�uBIS�<q%BG`©�'�'fsHАUQT�<��K�MA������rl@�i@z�<aQc�=�j8�!�S�hq�fMSs�<qB�r���	��@�&��[T�s�<	!� +U���㭇�L:L�5�o�<�PL �uN��:D�����ii��j����?�Ө-�J����Tn ��ϛg�<1Ea�8Wv!��m[},�(��m�<��M���`��aL�PjNx���g�<��N [��1rG޲&�q��jn�'�ўʧ��ikf*�P̠��G_�0b݆ȓ)L� !-����/�:?=��ݚ�	B'Y�Q�xA3��� �*X�ȓ2�����*�nȺ ������ȓ'��X�d`�����H�z̃um=D��q!�v�:����I�v��) D�챧nږ[��=bb5\"�Y�<D������!,3���%W�j.�m�:D�Pѓ��z���(��תT����V�7D�HB���,�����U�P�T �T�?D�21�˘F�|	�D&�1
�8��;D���K[=/��k�̜Tx �!��?D���īG X��z��J�"� ����"D��p�h� ^��@�O=�IP&#"D�@�π&&j�MT6=):���'-D��
�C�]�j�q��b@9�f)D���V�R=!`��Ze�؀q�'D�0��Ĕ�A�"�s�딭y�Ȭ`�9D�p�r�B�L�n\I�j�~��,��N9D�P�� V7�]a���n��H9�*D�����tx����4^���J(D�`unG�y���p$MJ3��1��*D���-��v��]y��I�K찑��,D���Rd�R)!6�BMx�ہ�&D��k�gO >IT������M&D��ᖳCY"�XV��DՁ�m#D�@@Jɼ}m���G�<nH,�h'D� I'�߬bb��B�%	Z6��"*"D�lDN bW�(�e�֡��� ��;D���=},0���{���(d;D�$���Ǹ��P� W�1� )�u�7D�X��N�/(�d��E�ׇMF	Ibk7D�L�p"Z�OT
��0�������)2D����5��A{�b�c���ǥ1D��1
�-e0��5��5�F<D�8��G����s7Z���qӢ"8D�Db�F��^s^���L1(�	��3D�P(b�
�)�����׼�J�h��5D��0#M�œC�W��:�{�7D��a�KB�<K�X*rXt�Aw�+D�h�Y�R@ҬX�*IgL�g�6D�@��TT�z�3d "V��G(6D�,
��V$B�T3A�6x��d4D���3іp�޼�*ΐu��0R#�5D�d:�%Y�F���ڠiQ�a��h��>D�:2��	��|P��zu�(&�=D��@ f�<H��,�S/GU����!!D��a"� ��J b	�,�`�ȱ�>D�� T�� �
�U���d�ո�@S�"O��#CL�7��SՈ�K�$i�"O�=�V��kk`�b�a�`D	�"O��u�^#^f�`b�^(NÊɘD"ObM8���:t��1Jh�\��"OtM��t��H�OT6~���
�"OY�逪f � �()����"O�l�V�Ԏ2����% �ZqV�b�"O�!*a*�8An�s�ɟ�W�bp��"O�!P�h�_�t ��Hwg�*�"O�U)LO�4(�&�k �Y��"O�m ㉔�s��\pŗ�P�"O���3K�<F�YR�;/�8�c"O(mc���`��� G�ʖ�ĝj"O��� ���"���0O���KB"O4�p��6C��8�@�g��q{"O�a�VCD�H�����JJ�P| "Oh� �F��+cVC`�A8r�0�ѥ"O��$��hr��SK�� ��i�"OL���Շ>0Ѓw��9+x�̈V"O�@��`��|��sɄ�LJqH�"O�m�F/@�(f=�Ç@�O�b|�4"O����hӕrB@e��&�(�
�{0"O��*��*��{UOX�O�P8�"Oh�
�$݆����%MX�a7�%8u"Oޠ¡�3Xk汁��6yO( �q"O�u�t*�"h�\X	7��'O��;"O���)�%m��Ÿ��J?���"Oȑ�&'�RXqG�.s��5@s"O���([�Έ��̐b��M�1"Op�kbLO"�B�X�F֞xBE��"O�Ds�gO�38���'�d�"O4g�W7Pd���^!�Б*�"O���g͸4mm��=Ɯ��"O��:��2X���K�=&�P��F"O
9���9\?)�'�*�"Oܝ��9=P�9 �E72��Lg"Or�j KѦ, ���n͒jm̐��"OT�!&GȖHD0�p����C[��2�"OX	�SCٖ8�<����BYW0@
�"O��B �A+M�8��ޥD;P�h5"O�5�f螜IT�s���?6� "OJ���-G.*J{�I#����"O.�X��׾:4���(h�XЙ�"Oj�y���n�<*''�
:j����"O���B��IT!HRL�S�rP��"O��BU�P<h��,: � Of0��5"O]�1�\3�.$X��F���l�d"O�p�*�!f��=�C˃<PR��"OF@Y�a��0�"����^�2�d:U"O��3� >�Zp-�湋�CV>:!��[�i~�!���@���-� �!�d�2��l����DX���:�!�$ߨ+�TA��̕Q#Bݨ�^>!��L0�:�b�[�,d�5"u�!򄊸qӸ�B� �0���G��G�!�d����9hFBu9%&��!���O8K����V�P]jV��$!�!���<3B����TtPq��,^�!�$�����9�L�?a2�r�ӻ8�!�A�`(+��D�� t��O׶3�!�d�5k��)�,����w���	�'K�IFP"*������oV�	�'�ڡa� �� jeEF�_���� �����57vu��\�@@lQQQ"O���+\�	`j|Q�_�"*�zV"O����� X���B�7�9��"O6��`�d�F��1a��2�Z� V"O�D�d�I�8~�y���\'1�$� R"O84���J�FQ��Gt~�! �"O���c�F �ڍ�3)aN�Bt"O4�㧞���Bř�|Z�"O8�p�**oE|@��Û�ղ��"ORr�GF*�t`�s�C C���"Oĉ�#FL! *���D��ZzH�K�"Od|K�j�Q�5)'E���z�"O�pp�뇭~�Lʳ�M(x^(��"O
h�ለ�&p`P�#����0�"O$��8nƤ��������"OYSK���
Q+e���X�"ON�	��<^�`�������Z""O��j�����2�DJ7y�q"O�arb�V����B�/=;�j�"O(����C���%C��Ħ��`"O�e��b�(����E�F/|��R�*O]�!��!X��� �5T�)��'����FD�?Jlx�g�J�!�'xZ�rC"��u`l���*��P�'�v�c�l¯ZW��#A�F� �'K�u� �&�5�JO�z-�`�'mT)ؕ��`Ւ�Ŋət�@hH�'F�@��/g��8��'X,�i�'��8w�Ԣ<"]Bx��2d�<Q�I�p-VȀ)D�EJ6����b�<��0Hس���g	���V��i�<�P�_�Do�j���9:��Cb�<��R+U�	��o�!��8��^�<�Dᔢ�h�bV�I+K�̸oS�<��L��.X����S�NV.�@�Fg�<	�ʁ섍�$�ڝjz��c�m�<1�F���( 1�$,M���Q��p�<A2'�S����K�Bخ�rS�b�<Y�X¶`B�a�+�F�?0�C��5`�x�kpϦoO����H#C/�B�	�#�4a�@C�P�z��T9A[�B�Ɉ1�\�Ґ��0mX�˦eQ�g�C䉜`��9�!f¾|��ZS�B�&i�C�	�L0ؘ�D��N��,st�ި[��B䉯6����� 8�j̲W�ڇ"֎B�	�K�@�0���50���`BU�%0B�	a ,jD���m�Ƥ8��>;XB�ɏ�e�r�H�WB��2���"��C�I�c����@����$����!(C�*i���(ցM:���kZD4�?����<&���Rʚ��P«�C!��N;��˅gC�Ve��ʁ i!�7
����E�^�pti�"s!�D��Z�T�B�b� �Jϭ(R!�d��]E��	΃�Q���"�!��H�yD�|y�£[Ў� �&T'o"!��X ��&�+1�`�B��X#�R���I�<a��ڋ@�|��W��x�@��!	�`�<���� ��EK�.�<6����\�<�w�ӊq@�E���/Z�؝���_�<���z1�؅狴ikx�[�T�<qU�G�s�#F)��i�"�#7�P�<�S㍃:P��M�`Y�����Jh<p�ū�^d�E�TҦ��A�̻�y
� @��$N�"/2°�C�x�P{ "OR�0@1���;�e��X���y�"Op���-X��ɪ���sL�;�"O�;Řm��m��cR>D8���"O�y%eGhI���O�x0\Li�"Oإ��5�z����^�o��&"Odx զ�
7
\��`�2� �"Ol��үѥ*�(T��b(�ɤ"O�= ��ɫ&�@m�h�;��ix�"O�Y��Q8=ƥ�e떑9�"O��;@NĒ��*�Λ�|̲å"O�́��^ȗd�Pԫ�ŏ�yr�J��ٳ�d Yb�zE�[��yB��Y��|�voW�R����H��y�28�`�H���c��O.�'�L��}�<�"�e�q����fJ=9NC�I}Dм��Ϙ ��Qp�ϰLA�B�Imǚ�YW�̈́h��A�bF�lC�	�[�=3�KU�$�d	�U�M�?�XC��%%�FS+�>�q%F�u�!��U,q��1j��{�Fp�q��\�ў�����Hp��V�6����ۥ>�f⟔���)3p �9d��Bbn��mC�C��⟨���L�M�!J��}���+ūG`�B�I�/�ܤjP�Y)!,���&D�L 8C䉤GBYBn�)|:�"��EC�	������ �i)�lR�$˸B�	R�=�į�$"�
���V��$1��O�l���cD�[P�I({̂!"�"O��#N<ZQ��x�&�?�¡W�̅���D>4P'���OZ�xpG̔,H2B� x��|�v	L/g�R�j2�"�BC�	�>m�(�wA�(!`~-�V��9(dC�	>Ū`U#N�xh󋔞Nܢ?I��	�"�D@ `�<�V���f��;S!򤞌_��)��l�$���%�pI!򄓢j��48#�A�&���I�cȟU�k��(��*�@�i���\��S%�#&m!�d_(l�'B�%'��9���/bJ!���<��I3��5��|s�K�;!򤓚81'�`!��6��}җ��*��Ö�hy��[�mW����2D�X!����rCI�S���M�<Q���S/X�,���B�0�	vh�[�ʓ�?1����D$4��9�0*ד��L�G؏4�!��2^�B�	h��H �%!����
<
���j�"�DՌS�!�$ɬ#މ�7e�0I��q+��!��I��&r������h���>k!�DV�D�:�Át�2{�*��9x���Z�'yve�.����!�I�=#0���'��Yr��A<K����l7�  H�'�Dp�l�V����$i0(�[�']8��d�'�RaC4��g��'L�i���7 ٚ%Y��R�2��@��$8�H�2�M_�#�t{�C'j�$z�"OT#T�7�,�+ ��.�^ �"OrLS�V�SDXI��!vE��j�����^��x˖����
u-�:k5��#O1D�F������EE�&T p,	0D��x�F�4�����E7h�82E�-D���VD��P�FESS�Pp��OH�=E�$��/u`i����DR ���)E!���#�fypc��+46!�� z`i��	AΈ�4��w/���"Ob�瀹4�f(�Ɔ+*0��"O^%�G��W�$��c��x���"OF���Ϸ ��Y��
�"�tؙ"O���mO"P��z$
O�u�]K�"O2]�&A��`c���U���4"ON�k6["l�]����A!�@c"OA�#a�  }��GHF:}�TP"O�L��_�� y%�pZ���"O~�Q$�.Qԉ2T��g� ��"OF	H�*ț%� ��̗5��9"O�,Hr�� �;�"]^*t�� �|V�<�ቫ5�����N���B9.2C䉜9�Hj���6����v�Û����%��W�Zκ@�f��I�|1�+��:�SܧZC�$��Dr^h�b%[4:J܅��_���+�RR��%"��{�d�ȓ��@�5�I)9&�Q��Q�b6t��ȓjL���T��*AL�;2E�8)Lp���[�'DXM�2�H\#N����(Z��z�'�f\x'<b��uذ�j��i���Dޑ@|Ј��'J-;ÂāG�!�$�,�L��7�C��>I[�A>\�!�D�`����5'ԫy8�B7�0>�!�d 
x��F�E&� `�ԩQ��O����ۧq�A��	:e<���l��v�!�d�yB��z&%�}?�uP#�������uܒ�T�cL(!G��|_�C�	�$�6�ɗ�5%�$ f��q̆�X�&�c�F4C�lB�!Q2t�i��C��<�1뉎thܘʗ�ޕeۘ5�ȓv�B(�GIet��E�r|'�tG{���m�( ,�tIRn�iA8��튈�y��[�DEŢ$�eqzY��ӿ��'!ў�OA�P� 3p��4+��������	�'f}9R�C�J`��S��F,��'��J��O��~ԑ�Lݐ�jYj�'Grl���^7Y�\ȡ�Ñ wv���'����B�� eЭв�X�v���X�'��`�g�U� ��1J�D��4��'٠qC�jƂ|ٰ����=^>t3�'�ΰR�d�5])U{v��6<�p��'^)����5���
v&�(sp�i�'�zȓE�
�����!'jк�'�<�{�C�g�\=+D(ڌ%06YX�'2��cg��(���`C� il��'N��!0�#>�ؓ1/�L�c�'���Ё�rZi����bGz���'u��PH�
op���=tݛ�'�&�r�gŷ[pLx$"�>j����'�l�k�9��y{���<%�1(�'!`��ɚ4��y���%� �
�';���cGC�\��⥀þe��
�'��s�S�T���#आR�b��'I2hx7���~&�2�.z���j�'=����ĤK���rAW(���
�'�PQrT���@���sQ�2X�Z	�'���H��+���ਆ��K�'��zD��`	ƍ�',ń�r���'�R��E-ܠzp��Gf��q;v�'�����å	�>��V��-[��\r�'��lQ��5�j�3F�ҫ?�D���'��I�2�Y�CB$PpA��/���'oz٣�['\�[ ��>������ U���#|8y��������"O|��O��P�4a��j-[x�"O�@�s��^�r�'�:7�>��7"OFi#Ԁ΂:��=�lxC~��-,D�(FJM]�J�I'�$:YL�1F'���� m�#f����*�����{ �$D���U�%j7�}X�T�m����r "D�(f�
<Mt�p� ��?��K�@!D�$���CT4\d����e`@���3D���N��T2M`�	Q�x4p���1D��"��5@TL��Z
(��=�!�$Բn�x����8a���2c�Z�c�!��0����W�R�|�*����!�Y9H��]s�}δ1�'I�4�!򤇩XP0(����CkHs�G١%�!��N�@�`��lĈ��G_�^�!�I\����K�F�ʅ�1&�!��bv���E��(�\����̕x~!�$��M���{ N�y��ҤhM*}j!�����P!S:���� A�z.�Oޢ=�'�y��2'�"���Ȼ1@rB�됽�y��J>�0@ei�[g8iK�����yB�_�\7��+����ND��%K	��y��
�PC��&��C�V�5&�y���6T���K�L�񫔅A$�y2�&%O�q�b���I���y�Ϡ�y ��ș��GH7v�C����y������g�x�>��`m ����0>у�~�X�J�%ffH P'My�<�Hȟ5��xQԋH'�p��r%�`�<�)�1p��	�T�͈����^W�<����H��K��ƿW������U�<y�j�"а@�G�
� O�!��VX�<�����J���X�"Z1.��B��~h<)��&4����D�.��Ԣ �y2��0�}�"�#lv��􎜾�yb+�02�	kd��1���#�NǞ�y��I�B4 �'vz�)cNL�y�,�x�ޔ�Q	�.^�i�B��y���?)�d� ���s����`#ǫ�y���;d��a��̰im�4�ЌɌ��O��$§D��
�E
�VTs2���e;	�ȓi�a􃙦8�蠁�웏K�x��	��A���$���
��'H��:N֨�G��-��RS�ܸ�ȓ�D��R�h�
�Ah�)f��h���b��ۥu7��Z���?A��ȓ:eT�⍏<@K���%�P�������A V�R�e�-.�zE��Y�ժ���E�!�F�"x@��� ���`j��H��[H�T�ȓmXFx �:��M�h�n��ȓ^t�C���gH���<1�g�^�<Yq
H/�:ҷo�6Ƥ	���KZ�<i6�=b���c�a��b4�q U�HQ�<y�-��,M2\:2C�Y�1li��ȓ?����E�MA�H�1nB�w
"D�ȓT��p�E�V-Wu�l��)�ȓU����WΘ�yİ(k7/�i��ȓ љ3[G�~<����30�<�ȓ���lH� �PY5�4!,\�ȓ1NI�nY1��I����6`�Y�ȓTk��p��H#QϦ �oB7a�4��
t���v�׸y3bE�Ĕ6F�5��S�?  ��������ٿk��!ٴ"O��@S��xTP���j��>�3��'���U�|���T�e:<���ЫG !�䜤L�fݪ�a�%O�	1w:�!�$	��j���$�='E&�h��N!�!�.&ֵ��d��XTK�
 ��!��H�VFJ��3%íe�����};!�d�<d�q2/����@A��O!�D@?EO`���G
�q���0c��:-C!�D�k��q��XR�x��w��1!�DχA�,0�E�\�n��6�;z/!��/wƬ-k���L��Yw�k,!���kX��e/�m�J��4{�!�$��9��nG�_
�YV��"\!�dK�'B�}�2���	����̒'Q!���)��=y�jهPy��C�J�gT!�̦+5>��� ˠ@�X�CV�s!��ȭB�7��6F�Ȥ)���3�!��[�9��P�p������Q	�3�!�A->�2�b��,K���ҳE	��!�DţFd�}��'�"��\ґ��K\!�$��v�A��=m2�Gd@�'+!�[� �P��#���ݹ�#W"!�d_�
���i�̛%j�ĩ����'!�Ds�2��s�J�vnD*���9
`!�Rb@F�K���dZH��$�,<!��@�r���(����=Z��!�C��k!��_��%¥�8]I���3�$w�!�dA�M8�`s-@	/h�[B��1|1!�dTN��e�ԵO��t��� 3!�$����P��ݬ��^;�J�@S"OD�u�P`�nX��B�)O�~="O8�&d�_Q�DH1���~�lSd"O�y`������.T�b�`�"5"O��6+ &�q�M�?��1{�"O�И��"ʔ)��<��)��"O��  h�-D�0u�����ԛ�"O�L��,CS���W�e�|E t"Oz�� �
�Z�$D�v�Y� 4����"O��N�hAF��*F�'N�;�"O�C����!�D�Dq����"O0� ���ԍDA�@k��P"O���F��b��VZ-^w��D"O�HJuG�����A�]�1\�%��"O`�(oA�(DV�C��$Y��a�"OJ�z��C�3ƈ-뒁F�d�S"Oąy3k�
6��M��/^ i�:5��"O�x*�f�	fD4���?L�]`�"O�e���_�"��K�b72�9�"O���VD��h~ ����{�a�1"O�!O��M�
��(�34���V"O�\�U����!�'��r)�W"Ofm+7gՂ�<��TZ-]�t�"ON��霖\f���h��Y���"O��{�G��?2di2&�$%��B�"O��@��
�
MS� �:�XZ"O��S��G-M� ��w����"O���2�X�(�d�q#`@m��pK&"O 0���N	N��|J�/G z��p
�"O
y�T�8Cy�b�N��`��"Or��T�&���-T&G��4�A"Od��6�"Ҙ���ބ�4�[ "O�aY��v�N��&��"�d�	�"Ox,��ٖwh�u����3�%a�"O� �	X�m��Aվ��2�={9�=8�"O6Hҁ�<?�vĻ����+J4	ړ"O�� � 0z�1PD'}B�ғ"O�$ؑ-�ɖ��2�H� X�$"Od��#���FK>�t捭G@$ũ�"O|4��gތn��i6��T?n�1"O4�	Ө�9��<��EC!?�<�e"O�I!�J�{�����O��P3��!�"O(yb���0��b%.R�@���"O"�����>	h�]�4h�h�"O��"� ���"ə6��K�\�&"O=+��^���@�X(�ʰ��"O���Q��1p��d��J��8���"O��Cw��k?4L�C�����h'"Orl�v�H�\�T*0���wv��@"O�1k�e`�v�I����v �0�"O�i0F�Y�u�R0P���t�>��P"O�0�ΉP��:P�I���K�"O��;U��O*���d`Y���z%"O�:��ۅ�4� e�9�@��u"O,���g6��x�O�=G�D*�"O�� 5��\��<��$�D�؃"O|`s��5Yw:�k7mYh����"O&q �f�
H=0�lSv��-ʲ"O�`s�R�A���اa� 0��T�E"O�<���*z�0x��4�J%:�"O\4�r����x�b/͸8e����"OJ� ߸u�^�XV��W�*��"O2��VG�`��g[6\p�ͫ�"O�xh`��N),�sB@�/MpL"OB�+Q6Z�� WN�p"�14"O6��5�$r����I����s�"Ov!��˙6u�1�o�x$�!�"O���W�Z�l2�l��n̓e�0�$"OH��Ȝ�u(�	e��Mw�Q �"O������^n(��	�"�012q"O��%_'b�����S����H"O����o��ppӇ�D+rЬ,Z�"O\�¢ș�o�}A5j��sȬ]�`"OB�j�:iAT��/�B���r@"O��!��z��eF�d��KC"Ox�7�D/L��T�%D�gr�UR%"Oҩ�
�,I�|m�r�E Y�	��"O�$+���  ~� "�Ş9)�)�@"O,���f�	`�6Q�E�Ϥ����"O`�Ks�fXRa(c�<��Es""O2�P�&V�4�j��7�-���Q'"O�uxd  &�8YQ�	=i$Hc�"O���!�V�vAV`�NەvJ���"O�Uj`�$�aЭ 7���"O��U"d�@$�e�͚R
�Eˠ"O�L��o�P�T4 �K��r'^��q"O~ �U��Mk����I�O'���B"Oj���;h���طD! ���"Od�肃ͭy!ƴ{@>CN��$"O�x���=���
ub�p�QV"OZ	8���3-�yC��Uⶊ�Y�"OrHZ�#��-�r#���$M�"O8���h�Z�s�$Ű���j"O"�c���^�tY���|�*�"O���uk��6_� ��FM?T���C"O҅yd��$Fp,�����s?� 2 "O�A��
	]0�H�,3@�T"Oha�L�X~*��,Q>o�A�'"O� NQ����0����tl���%yc"O�����	7il���+#�P��&"O�R��?1��.�8��"ON���͘9@7`XЅ���ܽ�"O9��H>�(� �vL�T�"Oİ��kZ<mbJ���#ԌZH���"O~\
�dZ;Mj���6��>;�(k�"Oh�y�I��>	��
�/2fܩ�"OZmP� ��3b�1ڶ,Y6av��`U"O����"�/�pa��͎G4��"O��p�C�)0%k��_�d#�YK"O�� ��Q�;&.ؘ�B@�����G"O�!J�j��	Z�%b���X�"O�5���Ƅq��D7fn�
�"O�u@�:HijV �`(�@�"OP�(�*��G��Q�fϊg��p�"O�8�7�ˮݦ��&��`�[�"O0!0�O�)N�	�?
&"%P"O
I3eo�5����"̾��"O�d��DO0��Pے�?� <�C"O��Ս͚�ʕxT���$Z\��C"Or)r�W9o��̣%Mjޮ�`�"O�q��Vt��2E۾a�4��"O��*K�閹�F�F%��}�"Oڥ(a���X&�l2��'��x��"O���%��  �R�1_�b���"O�=�GX�~x-&JŏP���1"O��!�Z�2-�xCI��o� ���"O�`���͝{7�h��Z�yp��"Ol�S%�\0
��d�[�O�:{�"Ot-�aŘ�E�ĥ��N��J�B�0"O�����Ȉi��a���Z�bB"O���5G��l��(L�j��l��"O��J��c%�24�	6#� ��ȚB�<A�A�dd��0�債>*5��Rd�<��@��JKc�D�X܂]�jL*!�dT!8�cժ�+=�,���gҋ�!��w��yH҉��H���zg�0�!�Q�}�D�RT�最�BH�x�!���_3���B�מ6�\4��խ&�!�$��eݶtk�FG&@y���'���S�!��%���h�+|vdL)�J�;6�!�N�Q�,�;0�Be�t�"���!�$Z=-	Xul�I$P�L̪*J!���+g�� B�
�Qx�F�
�!��վ}����R�H&֮��ĥF0b�!�dgd4��ga�0|��&Дv!�2*q�HrU(M�>��Q�#�C�!��44�>	��%�	6(X�%��"H�!�d�� ��I���,�4x��. A!�Ę�����[:s⎨pI�7*!�$�^��Z��O> +(�����3�!�$ai�(�
����`LH�H+� ��'��ȥʏ�(Ċ᪈�;����'��Ca��� �0���	F�.Y���'0�d+�D�\H��	�)w���	�'�J9Pè,}���r��ZX��'��ܘ�.��-!)���S
$�M��'�����f^D��3�!Q�,A>1��'��b�M�Vd��StƓ�N��c�'��P
�nN��d�co��GB���'��c�`ʫn��JTF�h�&�b	�'5Z4@��B_����ӫɒYp�y��'>�� ��$9�\좑�I�ֺpy��� �Y"7�W5ty�1�B�<|��1`q"O��7mR�H�����]�$ ��"O��83ꁗj՘QP�C�q,�0�"O�C1��!Q}��c[�{#P��`"O����쑐߆]��V�"~�HB"O@R�Ŋj�`�Ta�n]f�pt"O"\YƥO%h��9*�BM�onrU��"O���O-���!Vg���"O\в�S�:L� �0A���<�"OL�vCG�.���I�_�j�B"O�btl�v�9�����vaK�"O0��k�Lp�0�Ĵ_�4��'"O��kv �?w��(���M���Ʌ"OK�3����,��pߒ�(����y���g���iHf���Y9Q�3D�<����$(T!�'��%�ȅ;�d7D�X��\�(t�� ^'���{T�3D� �r�H�A�}CE�G��|�GO7D�����e�H� ���/!RIF�?D���eꗎ����;2"օ���=D�� a�@�4��q��޹(p��ra�;D�䚃(_5�n��d�#+��1K�*8D��Q�^%q�4i�fn�.����J7D���'�'WB�y����J�Y��K D�< g ׶5�^�I��C$Ǣ�1�?D�����~R�0�	p%x��PC8D�dx�)��x#��5W���� �7D��HdL;'�@,���W����V�*D��iUnZZ��Pe��-E���.)D�t`��\I9z��U],Q�i�Ƌ&D��T
^�e&��(2均���� l%D�x�9��%[)����w#D�$;t�nhB��^gv�ڂ�,D���3+b¡� %Ȇ8lE�$*D��2A��IL��#�`�AD�'D�����V�A��Рц�]�.�bSK$D���H�	2(����R:�c'�4D�H�q��-h�!/o��$���3D���I]�-k�IGM������3D��z�#B�s���f� �lH�t�q�0D�x� �-�
�G�7p��1���,D����.ŭD�E"T���OMNՉ .%D��+�n��=tu7K �����!D�p�\Q�IÅ�-?�d�٣���y���i�2�B��j��Q�HK��y¦60а��iU�d��{BhF��y�@�*L��y�gdڃd@���6	+�yhV׊�F-�j���y��Z�y҃��\��5P��I!1HxQ��N$�y�8R����1lWZ�dst!��y��I~�j +M�;ͩ� ��y��@�r��̘�l�a�Y9�+�9�y���NT�A�s���� ,�y�j[�	󒴣����W�
8��E��y���ph�*C�>O6�UtHc]C��,�"1c�"O825B�S.Q��� ���	ӎ3�X��֤�
`�!��/!��IdXD�Z�kw��!�D^I�3�.�PzFt�Uc�!�$͠h�:��q ǓcU���2,ӭ	!�D�aHl�AB�!G��a�e_}`!���7QF(��EM -;���"B3o�!��Kl0�3D���2%L�qcAL�t�!�dQc~܌�"�N
�`$A�!�� |�8���Uġ��d)�5��"O:�"4�U�d���ņC��p��"O�,��逇4D��!"����"O�]��� �D����P4@"O��*��wLm�ᩆ�Y� �"ODqy��-r�@��B�*�{w"O:ъ�iG�x��`!���n�F-�#"O��b�Ԁ3@�5{7�ҏCX���"Ob�3��%[��D�i
�T��"O�uZ���2vhq
6%�!R��"O�+3�Zr��0�X.Fh��4"O������v�$Ѹ��O�G����"O��r�U�L��B(�	e�Z��"Op%ӫqt�Q"���9�H�@"OĬYR�J�%8��h�%¨�^<��"O���MWqn ��ޟ
�0��"O�3�.��M���c�i�*D@ "O��y�-ֶT5��0�B��mu��P�"O�|�2OD�qev�P��m\a��"OZ1���I�Q�4�Wc|ћ"Od)��ö缀;��V]��)�"O��s���t��H���'>@ z�"O����H�/���ʱ.��Yf�p"O��[Ԏ�!���B���B�?h$!�$�"3���`"KQ
F 9�iG�!�gz@\W)A4 ���i
��!򄟞;�(x����t���#fG�>|�!�ү96� r��I��i�CƋ�G�!��:@t�8��Hf�z-�%�ۓp�!��-7�0�j��0�$��CE�5H!�6�R{u�G�D@��!i�!��8� "�Nk��w`D�;�!�D� \��"�ե:�H��7O�"a�!�dܛG\���J>8:fL���?`�!�	�X�広lT�	.\�5�D��!�$�0�&]`��1,*�����Y�N.!���0�4=�fK*H�Q�X�/!�DΦ���U��/))�Xۤb�	X#!�Ke$P@�AD�"�t*Ё��B!���9�2X�&��~%V�As"߂2�!��0V�h�j���!�p��A�?'�!��(q3��Z�D����(j���t�!���P=��HW!�50����ĭ
�!�$R�$x�hb��1�~x2Q�@"Y!��4S��ջW��9 ӎ{t+G0=!!��s�����"�H��0��i�
6!���+�nA��l�WG��C�aa�'*p��^$��*��o����'ٚ}X�/^�A��hye�_FP!�'EN@��\3:"�� ²�XE!���y"��nrr$iS����⳥L!�y��S�&@V��Ò}���Θ��yb`ҡp6���,��n�@}����yR#�1�`��p�?[6�v���yRLM�I� ����L�ʰY5B�y�)���@K'-�=��urON�y�D��^�B裯R�^B�	�GN�y�Ƒ��D�Z�,Q%U P�IS���yrd���x�(ϡM�8�`ҏ߂�y�(؏EѠ��ukS�F�,�!!i�
�y�Cy� *sh�=	CV����.�y��U�>��cTeޑ�X�:"�E��y�,��6�p9C����ę��H�yb�au���,^#���@*V5�y
� Ԥ7�/z�e���V4f���"O���Ɣu�B<2w"��Mn�s "O8�Y 敃T[�EsV���u�<�"O�];�_S���V�;��K�"O���LދM�ܒ!"$�L5�"O.<2� %M��d�WƗ(T���'"O����R�J�$EH��D.M�|Js"O��2D�J�>��1*&��1��IK�"O� �p�ަ�zs`nюW�r�##"O��xCa *�8d-�:^X[�"O��svM[�d����B#q҂��"O4k�hHTk
lV��"3S��p"O�A��^�P��0%ÊL�AB�"O�=ʆ��74��)R�]\��q	"Oj���M^�Z��i/1H�c"OD�)@�5R"~(�b�f�Ȉ[`"O�uY�� ��mi��bט�Ф"OƝC�1p(��� 5L2�(�F"OQ�ae����A���A#�p1�"O�)��%9�^�E˖x�(�Q"O~1%MJ�e������67���"Oι`�;_K��x%�d)���"O���S��%ah�Y+���R"O��g��7j.��ʕ��9!�d(�"O�=Z7� zN-a��Hb"O�����G��i!��¦V�L��"O�%��lZ���t��W�t� �	U"O���敍eA.���I���V"O�pH�K�HR�Yb��.�q"O�0����|�J��V;���"O�uI#C^P��)��;�"��U"O��8`�@2v@����)%9� Y�D"O(��a��)8m&���(�w�ƍ:�"O2��Bf[-w���"��d�g"O�Ey�>�q"�ƞ*���Ñ"O�@rD�A8RK_Z���"Oҍҥ�[\|��JP��� �"O2,���ܳ¾,��^�E��;�"Od�1�J�+P���dŗ�)+L�1�"O�|�"-Š\q�$�̪Bo�UZ�"O4�AA�@�n� �s
�T�P��e"O�|��N,\�n=���Y�_kI"O��S#*�q0����3����"O$}y��F4���r�������"O�9�U�:x�i���*V�����"O��"�^�nA� �!W<W"OҘ�U�L�)ȝZ��s�2
H�bC!� �%��01P��=u`� ���8@!�d��W�Q�FU�dA����G�9!���80C�y�Δp$&�z%!�䃋
p`
`�S$�bI`�<-!��V M �� R�U���D -v!��,�|�D!\�Z)\P��б	�!�dÜ���0"�G"t9�f��v!�dցL|��Y�Q����Qn!��b�}�Wa�&M��z�C�7Q!�D^�x��m�WH�x�x� �,��M!��\*tnDYq0�̨Q���a6�Q"B!��G?��R�kJ|n-��.��84!�ǽ�~$���ʺL��	�jFn!��2Q����*��(P�3�IQ�!�D��B�Bɠ
b�����X3�!�d��.���)�$t���7+�K�!�L&%�ΰ�=�Tm�CÂ�|�!�� ���Q?�<h��ځ`�aA"O�(�b��D{7KQ
4��1�"OVH@A��8`�幁��/!�̈"OL���eF�Q�~B�.��,����"O���P+W�k�t��n�op���"O���Bn-LFXCvlF���9�"O�Q�3�\N��2%돖G��ݠ%"O^�b2�Y�����)H*�đ;�"OJM�$��4&��(����b���K�"O�A����8U;����T�~.ʉ؀"OZ�#��1F�I�u��c|���"O�XP(�?phAf{!u��4!�D-X�$�f���xA��J�1!�D��WV�Q�W>e�D@��/�
/�!�і5�ciתN�2����M�!����c�`���\�&y;EM�%9x!�DP(:�Z��#	*bk&��SEH
!�Ȩr��tZ��êBM�M+�cԬ!�DU�D�&��R	��p�bW�w�!�(�J|X�J (w���BQ����!�dZ6$z fc�;JJb�p�O\�
�!���)X�}	0�)f1`�$�G�qD!�$�����j�-I.�CB���!�$�)8��4�C�D{$ԙdk�O�!�dU�p�<;��D� ~P��)ݧ�!��̵6|� F�2\la���GBP!���~��X��M(�腋`%��i_!�� #@ ��f*��k��!%Ym]!�$G��-��I;lT��m� >W!���D�فA�i��&ݡ:@!��g������Qs����b��["!�d��f����Q�v��� Zwt!��/9�Ca�_<`�z��	ز*�!򤋛%@T\�����L�A�N!��U�C<bl��T�g*D+���!�M:!h(K�[�"
��3m�~�<�I)
ڴ��u	�w�4=CE|�<Q"A�����d��)2d(���z�<�Fƅ3W�x�zv"Q�=ʘ�*~�<9�
�%bX��R �w�H�J�y�<��!D��^ĭ2��$����	�!�$%5��@�
:�*�� $�	-�!򤛏T��ZL�"�d	��Q�W�!����t,8Dk��%\��T˲�Fc�!��X	+-��%f��8�v�X1 � E!��+yv��̄# ͚ЙO�5^6!�Z�7bI� *@��q����5!�N�D���� �3s��ap�)��!򤍳-UZ�h5,� P�����<�!�$�)N|9�HuXI��lĄ!�D�H������_OPs8	!�$�,A�`���H<s]n��*.�!�d��yǲ��Wɓ%R|*R�QU�!�D�#m��q�ҬԔ7�P�a�75v!�̈́R�rĸr+D�^
�q4g�*9!�$[7.2��!H��F�!�$ޢF�ؕI�(ҍ�dyw�դ-!��٪%����b:\�Y#�-t!��C�w�l��HڵR�H@b��S!�5��:tΚ�jf�b�#��}K!��^,GdR�д���9<���(!�d�Pȼ}	�(Eh-ʰP���!-!��$<�z��r�_�:	��H#�E�`>!�[�W���Ae��		���w�	�+!�� <�!����l@ޠ�E�S)^����"O��9��_�]��LD(	E�-��"O�1t�]�H|Z]Ѫ$=;�m��'w@z���5���"���%�v��
�'" 4x��6��]�b�1!P`�	�'~@aѠ���� �!@
�� ��'=D�PW푁J0H(g�H#-���c�'��@5��g�Z�w���S4��a
�'x\\��,K�'���c&J�5M�1�	�'�֩˅
� (I&M�łɰ5Ǝ�
��UV����C���fm�x�$�2D�l*�EH�eh���G
68����4D���vEU�4ȕ��F�?�,4�$�1D��SW��^���:o�1|��9:v�,D����a��zs���6Nۯ,d�ti�F*D�<�3�ޱP����`Vbe|�k�(D� E!c�|��ri��N|�S&#9D�l��)ݴ�p1�w�D�7���"��5D�@����W�p��2jHD�Rs9D����Ƌ�\ǆ��$^��b�i �)D���Ǭ�R���#o��9�� �m"D�TC��-�q m�UN�h��K%D�hH�c� ՀG�B=�1�b$/D����e\�[�*��F�A0IiD\��(D��r�^� :����ñ���Dk:D�@
@��+_g������*nVD0�A$D�8��N�"����-���'�%D��k��D9}4-��$h�d(׫"D���k�H$��@�ጯT��!��/=D��kE��)m��\�Ј�$FVt8fo<D�h1#˞/u�@a�QaE��(��I<D�L���"pɊq �%V�$�C�9D�l�G��%�IRg��|ø�c 7D��P�F�
�D����'^F����4D�8p4��:w��9c�ݱbeVd
�#0D��Kҍ�-WtD*�؄ZJ<!F�,D��+4 7x��9k��� ;��s��+D��H�j3	��5keǗ�j����'D�x��X��Va�b�ӟ4��Q�)*D�d���,��@��")�pp�Ԉ-D�X"Ǥא CJ��-��L\[��*D���'��"���Į�K+H0�;D�Z##�;�L`��O��RnPaC(&D��kդ-T) jm��Z��2 &D��KV/��[�񧆀��N�s� D���0��^ߪ ����,5]���D�<D��ˇC�A����vQ�����:��$�S�L�z]����1#��u��HV�c��P�ȓ2!����데U��`�㊏�G՘������@��[�l�Z&)���,��|v.�*v*̺
w�9Hх�6|�l��HO?7���*�� â�٬&���񃟂!�Ҿn�{���>#�n�X�"�N�Df���%/-=4�H��31VF�[���<���4����.?!)F�2�z��i�(���@b�r�<��)��a�|�e+A�c%"	��Ag�'�ax��ڷ(NQ0s�ҸBX�)%�ۗ��>��Ot�9��L%J�\8�B@_��F<�"O�5��월s���`�Tsz��j���[>����6�z�*�;���R1D�<A��q���ҵO�	��Ka�3�O��g�hr%���Bj�.)-�T�P�0D����è���zVL��0��YWM,D���A��uW`Y���Ј(����.+D�� �s	���"7��3�$pH�"OHi;�M��pM�V΀��"����IK�OX"8��A�v�J�s#���I�b�,O����T(8�E.�$oFX��t���{�$1�d�<%?��O$.���H�@�|%��f�;?z���'�>�K� ėd���Q�ʗ�w���N<�1�'c�O��>�F�OJmF@q�o�3~,"���Wh<�R̓c���Ѳ!K6)�������'��z"�A��8���a�`6��EFV�<���U/��h�%���I��I�a@͏��x��,��%����l|HB����y2�Kr������חj(������>AJ��)�E��A>�Q��]�C�x��$D��Ie�D�~=u$��;*"y	 �(D����:_��}0��ײ����E%D�\�!n�;;��+��a��U[� D�\9��r��ҳ��1��Ai)D�t`�[�H֜�Ɔ֭w�D��G&D�D+E�,f�x�Q�4"�c�.D��X0 įi��!Q�)=G��SV,+D�Pbb���Ba�4Aa�P�6np���'D�@Js��5I5����0t��9҆�$D��Ig�]:jH�Ð�\hu (D�Dy�HH��R�
 �ܶu]�H*3F$D�lX�$0���S�ܑUU����"�	M���Oc��z ��	`��nٽ/<@�S�'������}2�rq|�)Î��)O��a.��$l D�4S�� �V�',r�'S�`c#P�` ��� ���~�Xt�޴�Px��Y(K�p��;u�ȑ�
�yR�CoAr�kw��-�f�@��!�y�#�Y�����0'���!����<y���-jF,��� 	�d�` ;т�c�!�d(�Ԩ�m �<Ţ��V���I��eʣ�I��\0ҽ�9T�C�!n��x�O�:��9��*�Ȥ��'�'�ayb�Y�s�	QG��4�0۶�9��<I�"�ƌl%0	 q(�P���^�!���Y�¡+anZ4n&.����ڊ�ў`�'�>����K:*ZA��ª��L�e�.D��@)�,�8�`��[��h!�+.���<�Ν-I$�H"���<�� ��T�<���4#��Z�`�;u�a(�O���$�O$�	%k�*b��0��1���2��<���'`�tY[4dI)?���@ ��-t���ȓM� x�o׃�,�W`��<lZOܓZ�6<D��O�����k$D���M��`D"Opȵ␴��0���Z�1`֨�b�*4����v`B��*G���tp�M;D�ڦfK cu�E�1DR�B:ړ�0<�"@�g?���M�JƄ%��S�<���1/]X��&��5����WO�<	��U\�	J���<��B6,��<9N���O?]2���y�@� PB\�{eR]˧-"�Oz˓j6�a�%.>��z%��������s�����Gʹ�`A�X�{2� D���㟅h� �Ó�]Bԋ4mt����		!xl�P�ȄBh-�L��
�C䉓�F��
v��b��:��B䉀����� ������h�����h��!�{"ON1A�rS��_g �hTF��yr�V#�$b#)P�N�f���A ���}��q�{���@�"�����j�9l�C��ҫ~1!�D]�a�����_H$2��A*��O���� P�V�={�4�#���j	lD��"Obh�c$z�H3M�k�:01"O�ԫ�ׅ(�d ��P�(�L,;���L�OH6$3�	�]��8���4k*2�(�'/
��W�[W?z��ǕyH,�Q�'(N)�����M�����	A����
�'L�R�E)z�fm�H�&8�~L1
�'���UI@|`�-8`,�F�
�'n�]1�A�4���oZ4xJUY
�'3x�
�疻���E"��<��	��(O\#��S�`D�jf��+M�p� "O����f�1UYY����]�"����d*?!���i.�Q`�ƝB��{�d"zAq�'�zms���c�][2'^	Ug��K�hG{���I�}�^�K���I��y!I�O�=�O��ܲ`Z!��H' \�b��|x�'7
1{���l��[�M6�@�#�'L��Q�ܿw<��j�67-�! �'5�M�ḥ2��l�/�&5i�	�'}p�"���6�J��6I�1�x�@�'k�=�B
�?�|Ɋ3�0.@~���'���S� $|��Í.�\�A�'�@�:��әq��$�0@ڪe�e�
�'#�a�2o@i0l�2g�"$��s�'���o��S�Q���
�i�'>h�"�<���c���-"Ƽp�'6�u�H��`�Q#�h#���N>����i|y��8���*��)Ẇ�t�!��ב1��b��yԽR�A�2�!��9� ���]�ʰ�N�N�!���|���yf�	�#V��W�M1[H�t��'��`h�|��a�.I Z\�Y	�'�h��%��5N�\��>S`d��'g�"G=m���;UkL'Hw%�N��p=)�}Bh	�*Ϩ�+VM߷3�
� ����yB��&�\)��J�]s6Z��	"�ē�M���ɞ�L�Z�م̍�2E��C��ʳy�!�$��t5qbaɂN;X�rC(W�NO!�d�4I�у�C
R6���s��8!�>UW�mbwJ"��e�Aj!�$�)~��0.�}�j�!_�af!�$�,i���b"��"՛U �!Ex6�ȓl|��c�˯#�V��4Xp�]�ȓo�R:���g�yc�ɘ�}�b5��LX�%�#愶[{$�c���	1H��ȓd�������>����eF`Vԅȓ0,5�Tj?�<0��&g!����*��#f%>�(x"c��&��ą�Ny�0�e�7
�j���h�~��h�ȓfol�@a�
�>�g� G�<��!mz@9��ي6�v����2��U�ȓ)e ����B�PjƇ�	�b��J~<PM-q��$Z� 	,`摇�[�h*�Ě*S�r�It�Q�&Pܹ�ȓ^���$
�`�YD��C�
M��9�@���w X�	�bܕ!?���G\�ْy6�$���;���ȓo �����]�D��G���Z!��14�i㋟��4	���d-���ȓ�˒h�1NM���V���L���b$�&[��a�6��P\�ȓ+4  ��ώX'<�6�P1 Q��
�ࠣ�0~$ur'��e�^�ȓ0s��`�O��=ޠ�3ԍY qٰ���S�? ll�L ?�B�����"O ����ʓvV�$X���<n���0"O��a��u�z�r%�U�H�೗"O��!r�
E�bM��lk��y�"Ove3��:Y�|D���24�f�q�"O�̫f@�����eJ�y�&u{"O�Ic�K�y@��[Æ�3Q
92R"O��µL*J�p5��EC�Gc^��"O��tD��\�����E�BA�5�"O�*���4.~�1�eC#ݬ�E"O�4hq�E�Y���´���I����"O���$��G8��"S� m+���KPxD�t�'����`�{��cRȉ�qbi��'�*���BUS�I���NElXi�'Yp%r�Ȍ����nC3EZzݛ�'�� `WC�T
ͣ�*C�>���'���0ƔS����*�:����'�ȸ���GT��K�h��-�ڙH�'�l ����V��JP+�p�'���ۃ�À~�0�.@̹��'�"�BW�R�[l���l�O���'�2 ��`�U!.���25��(�'F��*$qwĝ�A���g�Х!�'�E8�0}h�I¥H[6(�2�' h���V@��衤�H9D�0J�'������٢7��Z(~>bѩ�'^�=��%��T�0l)0eJ'w�^�z�'����‡f��q�r��4c�f5 
�'zt��4���?8��� Q&9
�'��#���}F 53�'^�3bk�>2{�9���A/"
����'�� c!愓i1������#c�R�'R����m����''���	
�'3蹫����ɪX�BY�O���
�'CJJa�V�9vJ�k��P�B,,��
�'j�P*V�\�f`h�#���y��!Xl䒕ŝ�( h�hpÌ�y�Fl�t���Bd�g�V��y�OV�o��L�d	���ypo��y�g������	��,���,���yB�$��ă�O�2����[�y/�,�x��e#�#_�֜�Q0�y�.d�Ek�'ӎSeYk�%��y��Ιz�j��J�l�ť�+�y���;i��ڦD�M�捰�h�yBES�IR�!K	F�X�"���y*҂�J�$��4i�{2,�yRd�)0�0,!�B
�*�:1���y��֮x�\�S*H8JFa��1�yR�W�;��`p�/Z��y@�
$�y�  XN�e�`��%��J�o���y��=!ڕH"��%ո �S)M+�y	-:p��9�EΒ%Q��y���y�D�=y߼�q�E�&@�x�#�l��Py�f�)z꬀F'X�+N�p���_�<�g`�hV��!J1��<%C�Y�<y�`WG���6��[�Tq�p��h�<Q�D�P�Xt�C��aQb�P�/g�<��D�$-=R%��"m�zY��k�c�<��Eن9
�ᘃ����H�jWX�<�p�۫�%���ȸF�H3m�W�<�wڛ>c�5�Z��>7�{�<ᶎ�= Ҭ� ̲8�
�; �p�<���H�&�zvm��v#��ۤ�[p�<� �,2Ӯ[�*$5cS��&]8�{1"Of��X�W� hCU�ͱh�  w"Oe�4	��n�mjF��g�j��"O� c&�ش����@{f�sU"O�Yc�&�|5V!ԢJ23�B�"OxM� jʆ{L޴���#zr��"O�܉��V(k��I�C�P����"OJ\3 �=ɞ-�e#���A	�"O8��lP�p�*��c�T�Oߘ�A""O�� ������P���"Oα�G�ǔ5: �� l��!�e"O4	Ał�uk��yK�1UQ* �W"O���@��҂i���W9X7� ��"O\x��C�p�s�GK�j&�HA�"O֬���A���RK�B*@P��"O
�y��ѱ,�,��ŉ7t0+\�y�k	ry�m#��9?�vx���E��y�Bѵ�tt�a���(��iK��y� 2@3�H)Eb��d�)�yR��?4��F�!���@�fZ>�p<G��W�Jb��C ���<�RS�&\����0;D��R3�DӘ�r���3Ӥ�#�M6?�ŀ�c�A�O>E�dbݦ";䨐ƃo�Ј��J�'�y"�L6�i�*�y�YS�&@�����7�F�Ѱ�6uZ��hOd� 2�4Qq(�%ՙ�� S�'��dP$�x�`0ɀH� ��
�#�&b�<Q+T*̩�	02�<�O�Q�6��	w���������V�d��Cդ��2����4�	����DM��k�����;!t����KH�ir�i����aH<Q��-H�����Y�@��h���('������Z��5p�L7숮�<�(��C�����5֣J1=�<d�u�]WF�+� .�y2D�U�((
�M�R���{�  !=Fp8Z%O� dE� p���?Q8���T�& j6�̃T����O��j�
۞F�R��!)�(�R����'����ɔ�a��:Dʈ�R9��5�E:Z垴QfI�#͘�i���0\�V��5��`�����'
2{�@N�i�4��L�s"0(��B�� �TX6耟��u���X��Htx@�f��HU�Ú%m�)x3ؐҼ��*JRW!��=s��4��O��0���H�G��s'��/��l�1�� y/��)�A�q���bL�5���Ctfӳa���j�$]�a�9	"M^�<�ԪZ}�TR�E�-)�x
���?I*0q�kE�"�Y5��r���D�a�N��.(?��ꈷ'Yhd�`I�.x��p[���V�ĳ�&�G��tp5�a���pIɡ;���L�/z���R�!
��,��#OK����'��n��9�Ҏ��ћ�J��y�<���(�)��)��R���ыŪ��$����� �&�� �ls�j! ;���CAƪ\C�ɾF��Zm �um�=С˙ z����L��7�%p�ĕ+jx�c��4�	{B��'�|����e�T��Py¬�<�$�%,ں^2�p��j,�������]����5�'���F�,O�k���PG�I���@.bdQd"O�u�Íڳ1A���g�Yu�����i{�EC��	1Y��%{
�T����_�;J�-�tE�=Y��Dy�řV���	�:H�%��>U���`���jVo�]�yic낁B�����"O�Rů
�t�:��$�M�U�� W����an.#K��h�.Q[�,�/�J�)#	�(x\c�>�HV��6z�Q���3Y>��y�'P���U�g��"/���g���x�XE�!�s#| ��}S��)U�`��Cp����kԼ���X��q�1��t�4��D6�Xh���o�$�cθa6�
�(��P
��9��F@S�c��&�O��#Ϻb <�"�hɁ�ēF��<��oJ�O�RD��&�81B� �?w�Hb��-A�ş-�d��rm'p`�4I�O�J���aԇ#o�aB��h�
��4pV<�� D��.G�'�ѡ�p<�%,C�ޱ �B�6GP\s����^�&D1��܊`,q0���6b��&>-fH�h�x	��,�N�3d��2,������.`�^Acu�}(<A7&�5̀��3"���\�6�	(qd�qs�L=-2$��O˔oj���&�53̘���"�	��@��&��y;��ۡ!�� c��.fT�h^f��X�b�\��}�%[ J�
��dh��S��Y{p�L1�N��DQ�L�J�s�I�4��1��;N�������Gm��	Ky�$$|F����C7@�q+���'2j���.�K�����i*��'��x����@�p��bm�&3O�����Z��d4̇�(�2AjC���*�ݲ�m-��E�a�MM�GO���se�0���qDA�T��,p�DX;R<d!#��M�C�����A�.xP����� �`�ъ�,3�Q�#`X�l�^���M�������}��PKC��x�rmՕ �����$lA��J�/�\uI�@[�p�9��� ��֝�TU�̻��ڡ��*�p!���͸�h��ȓ9}�va �G�D}	C��\�1��!j���6�^]#��Xb�I�),k���VR���u���x�Dş�Q�&Up�0�O�,�b֚\̼q�j�/$ �6��<���cu,[6b����f_���/��W�џ�� �5n�n-�A͔)���&5��}���0�F��AL�MlJ���џ]s��C^�oĔ�d�8V>��u��H����pbF�o�t �FɰF�|D���x����6M�!ʷ�9��A`�c�5l=�d@�D8���:|zfb�lU�kG�� 5w!��,�H̲����C.�J�/ܹN�Y��E.>#,�q�R��ʕ����#Ȥ\��!��� d(Q�QPD"	6ChD��	� �ĸr��Ŝg>��˂E�D�KPmY;�X��'&C*����Կ֒����0� (�B��]����؎���˖>\���P��:f�pQN@ r����p��� ܲ�ɷ�D/�B�I���!6�4t��$��M�uĎb�<c�0!D^��&�����}�^Np!�a�%!�l��4��N�<� ����T	�P�C�<!'�2	�.��L�B:�1d�O��}���¼���G1o�)aO\_����6�(�hM11�M��)�h�Din���
.&���dʝ	�"���c��x�Q�ʱR��}B�1R���m*(�+)e'����ݦv��B�
\L=�'Ǻx�����Ǽ�B�	�5�,�)D��x�� ?�C�i!@2���R��b�����!D�P��,Ǚ4���A*�����Vn!D�D��囐 Dh�u��i�%x7K0D����AJ�td�i¬��}n�ź��*D�8���;d�:�(�"&�lg�-D���Pg�;7d!B�G� Ԫ�9�%D�hJю�
?����X| Θ�tN"D��b3�R�;�1�g�Ү!��̐ �$D�TX͖!d��	ѫ]m���PL>D��p�oZ,y���:`�N�A2��$�#D����iŤ��H�͊]S�gJ3D����&��]ΰMi�	&�����.D����,o��M#`��[
��d�*D�$ �N/%@��4&�W1�-2s�+D�\!X����n̚rȢȲNڒNv�B�	J����'Z�#���jf�^3HB�I!�z�.
4ra+V4`�V���'� d���:.�ܪ6*�PR�]��'2 k/��qYAh�N�J�k�'sf�RD��2��}�РQ�O��e��'z��r���>|=�X�A&.��dx�'��A�Rn�M6EȡK�/w�\�	�'�q9F�E�&"��6�B���9��'�����21�)�0�h$X��'X��J�*�-4�� � �V��x��'9�6#G�8�����ߍ�RX��'M��R%�*:�j<� �V�~v^���'�,�r���<Hа���K/a6:�q
�'��d2�hV;�Ja�g��ݬy�2B䉥I������7��񘱌X*�B�Rmk�	R�6��aS�
}C�	�k�P"tL�6��y��KQ��B�	$2�%3$���A�v%��,�4d>�B��=$�$ċ#��h�r�BQ*��B�/5P-�r�J�(�~4���@�}�B�	#i�-��nɲMSrx� (�>��B�I�|4R�3t��޺�YD����B��>R��H�-��68̴k�%>B�IZ,�u�T�Y=2DB}XP��
�!��ǺtH�X��#��[g��� @�!�� &JFk�QC��D&ھ"�j'"ON��w/ݝ������<D�hHh"O�$8�.×�x�!e��c|�(1�"Oj	��~� ͪ��Q�%A��w"O��K ���?CMi�Ɇ�>@@�"OD b�2�$=�v(��ɂ�J�"O.u��*Ȥ`���i#�����3�"OH5���R ?[�ԡ6�ܮy�*�Ҁ"OL�x�N	#rF0��m�p"OU�J9Y3�t�0�C'!�A�"O�z�]P����]-��	h�"O�Q��`�]�X7h�;t���"O�H0�ل3��D2�(��H̰'"O�@�t�/\�`��K�u��Ջ`"O�@�BEM�Q���a��G"OD��&�ßO���y�+u�J�'"O1p 6���3��?1��"O� R1e�5�XA"�\=ʁc�"O3t �/H�jqb֢5)1��"O�5�'OQ�0�0�i��[�5��"Ol�./ �!fgܝ!	6� �"O$,Y�i��<�
T��$9<
 �s"O��:A뗏o���`���]��k�"O��ɑ�Q�7@���5B��b��3q"O����!
V~Z�ɵC^;"� dZ�"O��I0��#��`U)9t��h6"O�ĉ��P�8(���1�L�l�4�`"O2� ��8��rr��__`E)g"O�t��fA�ܘ���X� �W"O�A�Ј�:���r�[�?<�#'"O�E�Uh�|Y�E��-^��"O�aH� ]�Qtj#k�0B"OXX�4�֬m߲-���S��+�"O�Z��6�2e
����x�"O�a�ubW=hQNaõ�C�O��)�&"O�*�HґQ��1����G��s�"O��p�E>G�]y4!��<�"�"O>XD��u������/k�: ��"O�eضNHW�HE!e)�a p�F"O�I��KɂoHD�	� gh�k�"O�=�2�^"�b��@'ģ6�zq�"O<�;��[�u6P�#��?z��	��"O���b��V�pP��~d��Qf"O�J���q���C�G�*o��a�"O8݃���.@�<��n�;),�qc"OP�I�퀅Ks�,R�Pzu)�"O�t��ʘF�fe��I?���"O��{``ėU���)��} >ax'"O8\��+ ���jf3S���I�"O�4� ��c��Շ҇z�P�t"O�Y�� ��E*� �FM�����"O%SJ^5'�$����rR�x�0"OF��G�[�t��%NI��i��"O>SS"�539z�	�-��$�{�"O��@�+�VG")��o� pԌ�z�"O�d)ᧈ� @�0p �a�ƕ'"O�|��&��x<�T@�ܯ��8C"O8�s������((C���>]�!��t��L�̄7��hs��.|�!�[+3�X��`�ڠ���U"n!��KV3�5� ��4�l�p$��0-�!�dF�{&�P*`�� E��kr��'�!��3e�T,�Ҭ&D����7]Y�!���wqLa���>ў���J�!�� �m��-�!r�e;g,�s�@<��"O�b��E��H��@�Y ��4�"O.��7��6m���p���K�Bِ"Op���ѐ(D��[+� I��"O^�a m�2�V5��EYlJD��"Oreʴ�͸*`�!㗅��)Sꜻ�"O^I�0�ѬA�*�X�ś�Z�nxF"O�(�.A�="�Bã����H$"O�e��!T>��B��/���"O6���@�.	y�Ô��yr��S ��q�E�Q ,�p���yH��ڄ0���Nd�51Ł�!�y2�O�w=B�j��>�@�D�բ�y��*h���,�2,��J�	eT݅ȓl��q;w����z�m�8`��(�n�!񉛹^��:5��f����Jm��*�	0y����"�p��<��[p�Ƞl
��ucŖ�2D�ȓml㖫�$6rrQ���x�����4��J�.8ǼEJ��v5�X��=dP��񬝬?��L��ה4�����ĉ�7U�F�89Z�ɍ�;v�p��,3j����%0�@"��;v��ŅȓE0d�ꆠ�4���qJ2pμ��I�3t�p���d̤0�@=���A�L2!H!��5W!�DΦ$f,Pd��U9���ӠI�h��I3�x ���S�)§X$�pr� !l즁���$4P5��?B���G0��ݣr C�G����3�'}�Y�[=+>�Ad�	[F{Ꞔ3?���M��~ �tb ��0>	�'[�iH	!�OC$.�����	��%eL�� T
H���*8Ja�̝���(R�,2v BU�G���'�����ř8&L���$�\c��'*��q��6>S,�2f�!�D��d��B��00��m�"Ŧ7�B���j�>P�3S,_$4 FD*�����U�%�1���L��L��?�1d&$ �ጅ+-%#eL :���x�D�����6��EO�"Wj�X��	Լ���C٭\�$e�O�?�����:�����a~r���3�J�NϼiqtU��=��,AxH] �*��p�3�_�nθXk���z�k
�?G���6���V�bqzA�ȡ�0<a��
�1��_�;�᳄,�W�}��m����L[��?Lq�)���,��hz!�0���\���	rǃ�%8��	�'#V�Y:a�����~Ғ�+p�U�$;��C� ���6�ѧmؿ+Z"�#�9g
��(���:*�� 5��?b�<02�솾w6VC�	*� �C�"
@`�@�=yP�y�2n �<�����A�+ZЃW����#
ݣ	F|�b�%?� ��/gҰ�7CH�9�|pPj�z����k�P��U8���y�	k�ڕG� �1�䝻C�ź���@7�uA��FCʙ$�7O�M� ү��բU��_� ����I���E �@R���݊%�Y�4����
r�7�M\��S�h����'�y�!�d�-���1҂��lZ����o�1z�qO�L귉��D�z��$���h`�}���O�=��C�%ߔ<�:5�Q�a�<�$���Q�ҕt�����LU�1A��43�*UY��'�,ED�,O��aeF�F5|D�&CX>N�d0(b"O��C+L(f���J�<���i�d��5�r!�1e!lO|��#܇t�N���E�c{�|P���x����'�J�����fw�L �o�ߺ�Q���5��5�"�Ǜn�<)#���S��ĨG���c�PLI��
<2�]N�z������&ڼ�{���Q江��Wh����� 6�*@�#�O�!�d/e�d`�Rh�-~����ᕌ#1*�b+�\�җM�iR� b�O�`t�"�l��f�(�-(7�¬!d��_h���I@�J �Q�W��n�p��K�gF lp��U �܋1C���|8���5=R�	
ߓd�%�e��<=�49��9*����?)��=��s@ ��@sb$	��rV6���O�HP���5oZ�u���ΐR�͊	�';�U3`�� �(;�.Y:f34Y���7y��0��1@��������h�R��6�x��nD�5�� ;ӭ�%tnC�I�)O� ׍7+���s�+8X���N�r�RHòj��v����U����4-���cO<)!탺�1�� x\��sQ�Qf��8��e�9�
}
m{�?  ����0�DSUbח%!t�q�3!~e!c�i�N��℄�#�xr̓�!<��G���F���%��1��'�`A
�Z8F|`�O���,��#J�bϢe�C@A�mIl:�M�'Ԯ�a��n�PˆO�Ѐ�*_�x�!KM�%��3j��<��勷�܀r")����6m ^�X�f6λ��e�pC֮*�ehh�/"�ܑ�� �^��";��u�#�.�"��')|�#�k�?���B�n~Z�Ý�X�8�i7?I�-�.M�J��ɾ���T�B\�<�B#�*�U)w���l��`Z�]�� �rӰ�� �0<a`�V�^�`4@�8�F�bP[���+�ƀ
]���zS���^ӄ���XAиK�b,5!�D�����L-~��Ш �Ѵ�Q�h�1K �Ť����IY�mf\��A��<l�Y���/z�!���b�4iaM�?�
�� �ݡ(����
m�a7����)�'�~9kG'�0Bi"m��D��v���ȓ=|�I��&-Z����.d�Zi'��AG�Q0_�N��� VI�d"'>$�I����l�l��� WK��C╒q8��R�\v�B��C���x�l��
6��G�_>D��# ΁��y�eã�@��Q5� ���y�ԗ	Ӝq���'%OM�%&˝�yB��l	�����E�*I��y2抸}��#�m]#��u�`�L��yk:ms������vH��G�Ҳ�y��	x��i�,_�s0��fЭ�y���d�r�Q�M�1n�2i����y2'0?�c��� g(pEK�M ��y")
�C�( �*A�_��*��X$�y�'>0=�HP���OFP�Sf$�yb�m�0�hP?/f�2�F�$�y2`��L!ԁ�77�R�c����y"��>߶��2(�/>l"q�K�yۋI�cC"��h��й�y�C�]aP� ��^%�������y":fB���%D�(�]S�#Ю�y�hX�n�4�Id���5T6�%��yՃ:�(�; m<t 4���>�yf��c2�}�rKaG�t��	��y��ɕjt����+7�l-{4��+�yr�ѯ,����$�͒4���s�#�y2�ɥ4��y��ڤ0)����yL�O�����O0	B
1���y���cF�I`Q��Z�2�{`���y���2C����V����0�d,N2�y��7`0n�`#��4��i{�
��ye׀�cG-�:]zBӪ�yR���)�!܋r�ܘ��M(�y�JЋm�l�b���v��:��҇�y"H�feh�k�*�?��� �T��yҨ�8k�Pq��.N�H{,ڪ�yb�0D;��
� 44�CI��yr��OP����AW�L�pRS�R��yҌ�Oy ���\�.>�*��F�yB͊>T���"���9��u�$��y� j䔋QT��b�O��yb�+Ww�iA,Y�
f���Y��y-��@�@eA�����0�r/H
�yb��]�>\ �@�y����D��yb�	'v�^�[䦆 |��pR��&�yBA�u4Ȓh�5M��&AV �yR�ҁ&��;���8� ��-�y��C�PL���,f�����2�yB�#do�(����-��99�����yB�#o�Ơ��P&~2�p�u͚1�y�ݺd�IR�D<t;.��� T�y
� � iUc��z+��a��<��b�"O�,Jto:l0�c[��*�c"O���P퓔P��+a'i��j�"O��ˑc�G+`H�F��
E:$��%"OY��	�Uf�@��P�h8�K�"O���1��0YCĥ�"B��i�N���"O\I���S�8h1���FI��"O�8b5�4Z�%���L{���b"Olxb�W1����Nϐ`�p�
�"Otty����6�$�Ӯq^q+s"O�@N�#T����m�4~���3"OxD�&��[����D,ۨJhX��"O����J^ތ�b,M�{��x��'�"\�U�~��x�勼W��X�'�
�q�ރ�$�Y�d0FPB��
�'j2��D��prt[��(:� 
�'vԕ�G�3L��|J��-��h�'�~�1�KQ�E���
6
���'�=#�,�)���ƛ�[_&��
�'+���I�rH�tK�ИP
.�aG�H*o��P�3;�h	I��"�+VY���T;65�Ђ ��(�-˪qg 5��o��T45�4U��d����ȓ�a)�΃Y�59���F����ȓ9o��q�-η8���.R�d��|��`P�a��Fj6�0f���;-�5G|�O�U�O����n:(�B�q*W>:���R��ώu7������-��6�A�Q(��xa��	P�p"cLW���r�$D�ө̱MM^�k��釗/�p��wIG�cO*��1l!h�|6�Y�s�,�e�	�>�i+-�O�O�H��3oG�l̘�Pb�Y�S���/:�t��֬I�%ǜ1�����4��,��䉁C���������UA5H�2-L�0ԝ���J0��A3���#���B �ƈX�Z�i%�Y$1�I�r�@�j*�����K�\�rI�-�&&Zlz�����$��MM,��L<E��%�- ��nr�Dx!AXB�L�'����6�
cO�>x0ϖZ�d��aЃQ�$��g��$�n=�5l�1O�?m��bKn��8�FD�:DE3k�+.�`�	(�D�Ʀ�~B i"r��J�B���AUÚ����\�ç0zPY`2Hγ@R�k5e�{��p�>f������u�On]*�G�\��A߰p���jR�x2$"�S�'E�d�`�^Ґ���(S���	�Y &�G{��)C�d��}���@")CΥ)dC_s���|� �"���8:�O7�8G�㟴C��U�h���$��9 ≱S�Y�.^1i`�ƏJ�����<��<�~
���J H�D��*|�����d}`��*]V��=E�����Z\���Td��җ���M�e� �p?)bEU(P����c��>3��3�\T�<U��
$�(������e�P��h�<�nQ4t��Ί� ���d�<Rg�$q���!#�:(D����J�<A���&��M�,
��s�o
D�<1��L�M�$-����(I�f�c��Z�<��,[�wUځ˰�� b�N��w�@�<�u�Ǟs��Yk6�U�6E�����R�<ib@��v�rs�V�J8� �X�<�6�G�
u
�[Rh�+}��/Dh�<�0`H��h(DF%j
����(Y�<����� b�g�8�a�̔]�<��	v"çܗ�΁0$�R�<9҈��'���J�؁w��Q�<�%օgB�C�']� ��$�q�@F�<��"X� ��KRoPB����@�<ak¥Z/��e'ɂU�Ѕ�D�D@�<qe��4�̤pC��[�U��/G�<���6B�^�PFȕ\@�A��X�<	�fK'�v`on�L�ȃf�*�y
� ���U�4"5~L�-��krms"OH�$�ɚt��0S��E
;�Ș�v"O�\�C��<��I�X%`��a�"O*�2�7<��1�nR�tH�8��"O�8B@�1���b�ѐ9�J	�'"Ox|�`�7G�<�K���0i��:@"Od�"E�u��d$Ö?�����"OV���]�x2��W�V�+C�R"OJ����ҿ^B4�x�O�c�ZmAb"Oxx{Ċ��L���G�SR�IQS"O���Ǫ�5D�LțU���n=�x��"O�U�&!��y�Qʎ0^2:d�"OJd{ai�?GL��p
<&��!�"O��[-I�>i���S�rPh#"O���(�d8�TQ!�C/`ؘ��D"Ovs��1g���9��7l�>M��"O���lϪ;��
bj�'8$��f"OVm"����1��ĩ��N4$�H%xA"O� �� E
ڙ�"�M�0�
�"O�ٸ���MD��Ha��5��sb"O|�B5�1n�j�P�lB%��h�"O��a	�	4B��H��-"O���s�1TQ�1q�٩G���b1"O)#b��t�Rs�̒�4�r�"O �"vm&�� ��]ZbZ�w"Ot�5L�8l^�@#ڇ[|Ȍ�"O�\
�(�dF��c�^�"ܐ�"O�L�WiH�/4x�2,-2� %�f"O�yd'ƸfY��`e v��R"Oԑ ��~͔1@D�f�}�"OB�y�a&!:r )��y̤ [U"O.���mՒ4F0�y���Ԁ���"O��D�¶���AT���N�>�q"O���DLX�E5��2c�Ǭr��:S"Oz�I 0e�py����Hl�i�"O�P��AO뜈
tM�KF�X�"O�ґA�<�yz��_(C��!"O������^S���#�S�hB�8�"O��A+��^��b�.P\�1��"O<����7
ΰ����`�3!���DIa5��:�-���< !��C�t`��>jty��ϝ;{!��[�E�BI�#G��y��mi��6e�!��pA���RDݫ9��CA�t�!�����p7CG��t�N��M:!�ސ9��B>�~q��RK!�DP$+f�\K�Z$7� ܫ�Fȯa!�D<� �i��צq��`;s�Z� !���!*`Y�e���pt������!򤇱x�4��-F�^;� �Cۮg?!�ăcJ�{A$��CF`�[�#�:!�ц�����G��s+�9`iΰ]5!���ڣ%ؘQ&��"��Bm;!�T�|;� �A�2(Q�cGF�F&!��.Q44�5��H�1�UGפr�!�D�\��Y���
�Bp1��h\;,!��}	���'���j֯.c!���4���dM��]��D)!��`��B]f���
ը�a�!�$�� �6t�Ҥ�.6�`�3#(K7<�!��'�NHQV�4s�DiǦ��:!�dKS'�����ك�X���e���!�d��w�U���X!��M��JV*>�!�d\���IO�����ؐ/�!�� �`٤jU ?����Z�6I�c�"Oh�as�J>*lpW)��/�@�d"O0�EɌ�F���d���)��Bp"O�<s0�Q�xy�!���'6��LQ�"O����e�}<鵪Z;v�c�"O�	!���/E�h �w�OY2B�K�"On�Ũ\ o� 搚~$�"O�<2㍐	�6�!�����"OP�S�	 �E��M��b5D�"O�娣�ΆR2� ���bTzl��"OB�b�[�M��䱢�F<	�"O؅��S*ژ� S/�\aG"O�� �I�(�r�y�4&���"O�ar ��h�P�C,	2~�J��"Ov-R��%���� K�k�pe;q"O<Q����b~�)���"L�b"O�"���t�B�%@�AC "OHu��O6�z����
�^}��"O�EAs� 1
^�*0��o�� �%"O��Zw�9��8�uM�JW ���"O�Dr��$Z�;�͌�"SH�@"O�f�~P2�87旬,�!�$	�C���!m�0K��p�R;�!�䀹��������!���� m!��<U�q��.$�(���Fr!����v]��B��J���1tMT�Oi!�䓼:��y�K�F..� &H�~_!�DԮ�����n4{n"�5e�Qq!�D�K��t�.�-,�x]�dCm!�Ą� �
<S�.8R��U��Bǹe!�D�3h~�pS�E�7o���0�8F8!�dH}�CU�-���!c�-"!�$���
yr +�iz|A�gͥO5!�D	4�>,��	�p�`�c�P3!�䛸0�H�b5H<��e�iו8�!�d��='���H�v�C���,W�!�D�Y:%;1i�^�^\`��͠]�!�$ǲ[�tM����$��Ux���X�!򄁊1�T1c�N�4"_<�"s)��ao!�!A�4-z��X�\���gə:n!�Ċ)S�TY��4z�� C��d�!��P�O)L����C�x�[�ǘ��!�d%�Z�I���6�� ��P�!�Ċ7JT�4j����9�Ō�:�!��"t�le���6
pÖ�ۍ;�!��"2�H�0v��?F��L37�V:v!�d�)�:y:�j�'�Е��!G(b!���	b��HS	ӜfD�!r��(`P!��@�U1�٨�L�u8:�3+�;.�!��?KUzc�ͺV4 ��iRM�!�$O1H���W."��j��1�!�$�2c.l[pfČR2�)zí�1b�!�䊆]�� P/0�b\9-B!��Y�v�c�'<_�>�qD�W��!��ʑ:�4m[�*G'�hDJ�mX8�!�I#>|���BJ�K�.���L�+�!��Z�Ѡ�e��Fz�B�ז`�!�4+,��aM6B�
�@���j�!�d �5yFЂi��)��$�	?&�!���K�Zq3�*]�bC���0��52�!�dHf�|X�J�M��� �A�!�A�\��K�f��yBU�N�N�!��҆9	Ĵ�铩q����թȹg�!��P4a�1ypަQu�(Y0�X�I�!�� �"7+V(%��"B�Q`R"O�i�Ǧ��F�
@�ހ�$"O�� �� >d�QmS�ۄ�C""O�Q e"9h�)���o&Y��"OP��Q��?EF�8�+��EX�w"O��i�˟����"쎳%DNDRE"O&)�A�#@U�ASCd9£"O���aQ�e�!��U�F5���"OЬ�����5*�J w�Pxa"O�4�q�[Z�c`� H��"Oxd�v��6N�2�c�ň6�j��f"O>D��E�=C��(5�ʌO�,��"O�`�%��mzld*C4=I� �"O��ڤ��!6���C��Q ���"O	j�-�-�L���B�{�4�"O}��I/>��t�� �;(�壔"O�l+��"���3o�)j^=�!"On�ٗE�)6�ac����X�V"O����Y�-��qbA-ǭZ�^��"O.TC��ƓK`��	C���ڰ�"Ol(��G�)��p[�g3��0�"O��&J�I���j0-A�,���k2"OtY:�	P�/�=���?�Ȣ�"Or�f*�`�!�2�9��˷"OR��%@�O�Z��F��2�cF"O����	3<�\JG�X�\e�R"O6��$�\0A�༊�H�n��i�"O�p��hʶ(�VEC��+>F޴� "O��2Ң�-$8��d�ѥ>ШC�"O�ᚴA��}]<5� d�#b1��Bs"Oh����كWp8�(G��A-:Q�"Or�A��vh�A��S`����"O���!������W΁�;�fك"ONa�f��(d��S`�-~���`"OP4i�mԉi8�5Qv"^{���e"O���@Î-qN�k���
> M�T"O�IgI*y��	�&%D�9�a"O>I*��Ԁj���YAF�
r2�h�c"O�[Cb��f$ʀ�A�	>��pT"OR���
K	nކ9��z�Q��,D��bM��}2P���F5��T��6D�����̀X��A@����z�9�щ8D�����%�9Ht�ߥ����!5D�@0 ���q��	�e��$#6�1D�p	e�ܨ3� �q�#�Q?�q�/D�`�c _���Dj�N�4ɐySU�/D��У�Hv��!Ᏻ|���r�+!D���R�U�FtԤ5��k`�P�wA?D�L R�:x:\c�JTYު�H�%>D�4bԆ   �P   
  `  �  z  h'  b/  �5  �;  DB  �H  �N  &U  i[  �a  �g  5n  yt  �z  c�   `� u�	����Zv)C�'ll\�0�Ez+⟈m�(w��I�J���D<c��.T�I���L��qK�%ߟC��r&c��\-����+8�:W��z��� ��4!SuA�
!���K��	�fbM�7��Y��#Sj���/��{*tMAt
����iQ���cG���R��;�r�J� ��1�0k�\�#8��F�V+t?��A �'~4(��mi�H� �~�,�!c�O,���O��Oh�S��� *9�h1B@E4:�HQ��O��?iܞl�uy�'v���O���'�<�'�*l�R��࢞����k�'�BY����xy�ƚ�M��'�"O^c�؄a��T̱#
��X��=O�4�u�P�qhD�!�%�t*�4*��	L}��ЈoCb�"�O�fy�+�+U�$#Bm�#pI~ �ԅK�?���?���?	���?�����yޕ��Fϡk`:���X�$�i�(�O�1nZ��M;b�i�6m�O�<n:�M+F�i��6-�Od���\��t�7���QSk7�]k~"JƁ��(���8qI�u.,�
���&x��AK�:�V��f�½�M�2�i��6��f��6�,�ś�jp�QЅl��+����b
�
0��DХ"�F�A��S�@\���q� p�lL�Q��m6�M+ӿi��Q��Z&>1Y��A
Q$^�9!�,!P$�Sh��_4�6��릩�شd}���b�/ ��]>�u�$h�]k���f��as��	�&`�T�W�� �*͕#M�Enڎ�M+��i�D`c�J�&�h=��m͠B�]���%(�A2
N�`)p�8s?$7�ܠ<If�����+�<jw���d*�I�I�&<[$�� ��X2��W��P���S���?yI>�&��uJUGǮv�AR�`��p���[�<1�@�,,���2��] /.�}0�X�<��$U/)]�-����\�N��,KQ�<�S-��|v��{�fE�*�BH����N�<�U�d�����-N��4�a�<qeO�*D���O/$��5)�Z�'��$����/n�*gi��HFڽ�cL5�!�D�^Y0I1F�/J;x���V�y�!��˂H��'$ݍ3/��y]�����'M�R��6Մx�㋗I6R@��'�H�1��9t6E83��US�ě�'6l�Kt�<q�A;�B�Nq� ��;h�<Dx��)Q�@�XX(�� YȊ��1gm�PC�	�*q6р�`��g�bA�t S��DC�	s�P4hG�
�X#B�'c�2$.C�. R��F�D,>6Q��G3C�	+2l���rg	(����L��B�	-\��9 �G���,���w��ʓ`����I.umrJ5/�%Rb��V�\%�C��.DY� $5����R\C�	�3��pH�� ܚ\ئ/Y� ��B�I�T�ʭpуǆ1 X�y��X����$�I��l�g�A+:��Tl��y�&
��6�O��d	R��'�s:i�Bi�+P����O� a6'�O��Dq>A��Gf ��)�> O�����s�H�����g�^���сk+.�@4�S'葷�%�4%# �15�x�
��>[0����	����O>�D�O$��s!�6�fx��F��`G��<�����(��I
�k�<"`<�x7��:*xά��'�l�DX�V=�j\����V��]���L>�M����?,�,�y� �On�2���<�HL�#�^-sZ���F�O��F�>e��9%�$Sk̞<��m�ϟ�5��;6D�Q�5�'TS�ĳ���
�Q�|ڦT��ΫP��,`��E#�"�O|B�d�s~��Ûi����N�@~�C�?	��䧶�OA�D
� ��$�~䠃���2��L>!���0=�5��8�8��!�ٜET�I�MW�'��}�fb��zޠ��E��E4n�)ƨ�M���?��9��|p� ڬ�?���?��y�*	~��z#�!�9A��2�$��
Q� U��X���	'������T?�X.�,����^,I�qx�b��[�7��1X,M�e�M�FfD�1m;擫4F����O�E��:�|�2gN�/%���9��'y�I^J6��6��O"�d�O^Ze�ʓVL��奀�5�Ҭ�K6D�\��#I�6bV����]�w�l��h�<�v�i>��	cy�
�!�8�ťR�2�	0O�>���1�'Wa|����"��I�.^�4��p�g.Ru!�
�'�0��u�!A����H�x���RvH���xE!CoN)8��iP�5�I7)��͓�x��ўw��#�A8Y~��3����y2-��W�m9c��X��h���}a�&�|����y��� �\,n�ȹ�`�U�<�� E+OL����%-'40�䣙9@�4� ,1ڒM6r��x`g�E�\��Q�m�=�Jт�������%�ɺo>P�iS���5f`k�2H3@B[���ҖLR
qD�A���]Q��{� (o�� ����<I;`1i��m,�"#��l�	՟���ɟ�&?��<�TG�Tʦ9���y(��&��b�����.��U�G�rX0U��)'J���~y��m��6m�O����|��)Z)�?q�@��΀:�"�
7J�;5B��?���Kk�$i�����C�"�9C͟���d�?I�խH�4ܬQ�k9����:?I�	&��&.D��h����v�ё�4�Ӊ^J�1�aw5���U����C �2�'��O�1�J�����)L�1�G��1V�pS�|B�'�azb,�
dܼ�;�h�9	�!"F�G��On�D�.٠~Q$����A����S�%䛖�'g��'�L��QjǏA���'e�'M�n�*�� �Vd#���uJɖ15: ���%:�e।�*n�L��P�ISq�I�L}&�2�d\��"@��Lcn��U�1!�ذF��w����6�S�8wx=�O ���\E�����F� ڮ9PS�'��I�OA�d5��O�d�Oby�
P����ԍ�,D��1D��7C\&$h��8!��Q�'E�<1 �i>��PyRP�?� H���+)i���(<&���S$��O���'�b�'�"ꧣ?���+�HxE���Z���0V�U.\��g��%`�D��W8����yi`%["F�/����^�Y�@0�f�Z�E����I14�8��I�i,9��[D�2QY�*D�3 �C��ON�$Dզ���ey�'9�ON9�q�^��P	v�V��E�@=��5�O��00�\Q-��
`��FzҬ���|�N`�f�d�<�-F����X�Ck�W��\)�b�>(�쩥�Lퟀ�ɳ�v���ݟT�'~�n�R����'
�ew�'tJ<aP�AU`�J��:��iz���� �2��ۭ9�p1� �@s�J��Q�A�GRp8��ˮ9���>9��D��������I���Ĳ�G *}�v��WԵ�'"��S/os�$�!U<i?Q�Q�M	C N���П,���V�����,����sk�O��O���T!1��Dr�=��ՆD���"�j�F���[�e/D��i.B�mX�)"'U -���B��.D���e�� M�VГ' R��	G�-D��:P�s���D	T2���h��>D�����2]ܐ�,�^�Bt)k>D�L�%K@2$d�9a�D��M8�	7��O�ٸ��)�'��Ep����mHT�٥!S�.��;�'YT�������B�L>z���+�'3�ݪá߂��1Q�[+@��Z�'�
��d�q��;��?0y���
�'�\|�%��$Yqt��ϝ&�
x
�''����c0��jG�% ��*O>a�5�'�>�#���)[� X� ʿrg� 	�'�T�Q����X���G��?8���'�bp �)
 �H�4P :�'T������4(����b].2�j4��'q�h�ˍq���g�E�*N��U�Q��N��"p�� ��,��O� �@M��%��\��� +�����P5J<�ʓ:��� �N��(�:�%@�n��C��:Y�л��4°�s���B�C�ɔ}��XJ@���l�?�M��"Of��E�`�*TQ����&�Z��g�If���~j���1<�Z�Z�ΏhB,| �͚j�<1�
�wIX�	�L�"q`�@�P�<N�	UY,��VIFR�h��#��H�<�A�ʥ$Q2�S�K�^R�p�Ӊ�E�<!�q��h�&�nePB-7tk�ȅ�>Ÿ�;��0KĤx1ALO�~��@�"<E�D��S�8<ɤ�	���Ԛs!�$K�8�d�SÛ�"x�@kF�Yt!�DK�ekvti"Iqet���
$�!�dS�q��E��"�h��q��!�d�-'b����T/Ί���  �PyRƗ8,zT��.�`f�Š�hW���D�[��|�Ko��b��o y��გ�y
� �Qp�����y������k�"O�Y�������ݷ��� "O��W�H#R�܉��l �,*< U"O�dP��?`��]�M��/��q��'�-��'�h5�gJ+RD[�mY��pmj�'f�d�4��IՐ�i�+V.}L�P��'B�	��"@�!�1��+S�]=�[�'$H3��Φ[,�=��H�@D�	�
�'����dV��,��Q�ӿ����
�'n�R2�޵�Hݫ��ئtX ����d:$XQ?mȶ" �#;�PUý,oq��O*D��y��&�>p��B�1�Lx�d'D�Ta5� [���j)b�t�zw�2D�h���Q9T�P�2���Pk��h�2D��v-#	�2P��-�	�Tp�/D���t(α0[��S�IF�P����O��D�)�8F�9 �D��x�b�&�Cɴ�	�'���w�]�ƭ�RT;h� �	�'��HPKP^x.M	�A�,��%	�'��=#4o�`Ř��K,2�z�'�X�`]P0��Qu$8r��1	�'��x�u�� � ��J�UtN�
+O��{��'���R��W�\�Y�XF˨���'�ep�a�i�@�aQo��(ق
�'ậz� �(�fd��;^�\�4�;D���my5�dA���I�JI%D���gԜr�|�D�����h>�O�u� �O��EJ��{��(��,��!�E0"O���U��/��jB˚3N.�A�"O�ȁ��=7��d�Dg��/6vx�0"On�9 牳`�.T�0�P7R'B��"O�<[�(Y'i2��!�U%z�p��"O�ا�!KQ"�J�F�p��C�ɞU��~ZS�@�x�U��N�J�T#��[�<	f��ua( �p� (� p;��HU�<іE�7S���Ӊ�4ił�J$mI{�<IB��p��� c_(9���Jb�t�<a���/X`
<����j��UbRo�<Y��S@�@�qiC�Xrpb!K������>�S�OI�@�$H
�(T�@�u� "�"Or�b�T�}�]�uFd�s�"O����^�Kf����i��D��"O���G'�=j�R|���5��0*�"O�@�`���
2�w�:W��}r�"O�q�Ȼ:�L�	b-m�zd8T���v�7�O���@\%b7tpdC�#�
0""OJ���U("���!GjۃJ��8#"O��)��S����ȡHJ �V]�`"O�����7t:���� �R���"O�Qp"#�,X�%����0}f-��'���s�'�\�����$?��`p��@9C�V�:�'MԼ���Xy�$���[�ntH��'�@$�B�]�C��%�!���	�
�'����7iְ4u� ؀�ǵx礼��'E�Dk���;_�QB�
��i2Z�@�'�*�(r&�2r�2l��DQ�n���5�Q?Ղ��Q��и��ʿpK�9Z�4D��!0tYL��
�8�R��J1D���bΞT{L���� \Ըa�#D�4�T�X���	 #s%t�� �y�뙤9�LUZ�ņ*K������y���'@��\�F�6YL��'���?�SdZ���� q�������Z!aJy��z1,!D����e�L2�1j�Iۭ,^��#��=D�� �y0듹R������V�-a�e��"O�,���H, JA��L�dv���T"O�Y2&F�E��ʄ�2vX:!"O�H)��ʵW�|}�G�	u@XCQ�D� �O`	ɲL
�X�l�AP�@�s��Ыt"Oօ��
��f�vi�H���$uj�"O ���!��B��N���l�"O^�ء�$=�E��ǰs����"O
�f�oW�0㔮
�D�lI@T�')����'�*��P`�:�`̚&��:UI�'ɀ���T�4���y'�0u�ez�'�|i!H,B��X���!�~%��'���Cc��#�i��<��'^�Tz��%6u3��6hU;
�')�}"��H'c�J����;'0
�@��䞵`Q?1��[)C2܂7d�')`��Q# D�ؙ�� >ߜ,�e�W�|,��+=D��e�Լj���X��
� jv�9D���A,@�0
v$�[[��t	8D�L� �_D���84hF6�����L5D�{⅒h�rdF�[/��@�d�O�tzv�)�'J�*��Ǐ�^FJ����-�@9!�':d��D�� ���Kѓu��)�'�>�z��̆��b��j��Ђ�'U^u`G��l@��j�n��P�'G�9H��$3T�����d0�5�'U�X9a-�Vk���#��"U<x+O�P
��']W�	eQ
4�SGZ�C��\�	�'��Js%Әw�Dt��
ۘ3�"���'b�K�oǿA�� ���VA��r	�'�v�a�K)97đ"��F�cM���'���k�Y2e&��k�`�`��l�:���Y�����%���Yg�N�`�������	>R4�dH:�<�ȓ~h4���hܖp�X��u�L�0}t��ȓKb����ȭ2ܐ�A�.�+�B��ȓ6j�:%�[�L#��IͰ��ȓ(�lX��y�����FݠI�v�E{�ɕ�䨟�i!�J�]*ܙ@�U*C��l�C"O�A2�Ȕ9�:M��I�X�p"O>����d����l��H�"O�� 𫇫\byw�%㢀@"O��Q���d�>%jP���G׊�+"O"��4�l~X�����4�J��'�"�:���Ӝ ��G��m#.<`7l�9b����'�me��w{Ԩ�"(��Z<��ȓ
��@��	(Zl*�P�P�?�����I��Rч�b�hD*f�."�H�ȓ�n5��@.����e�ӿ2�"��i���j �>{���#Ŕ����'��D�p=�d��!2�ׄH�D�r��ȓ@U��0�M�!0֒��֌J΀A�ȓ4��QKZQ���� ��6:�$���"O���ER"�2����+}�ZLh�"Of£�O�kLP0!rK�(�H�Y'�'m���')��3CK�55.��$"�����'t�%���Ћ*I�I�S�:�����'�QYR�Z6J�H�B�L�$.����'M�l�m��[�L]��L,Y&С	�'^`�S� � 6�3W�֬:�6���'����!$	.��떇��+d�������CQ?9;QJ�7d& %y-�A����A?D�l��X�]XR����DK����I=D�d�G&�Es@��Ti�z�h��0N<D�� |5q�D�kv@KF�0�Z�Y�"O�|��Ȃn{������v1�1"O\�A�	O�\��M؊Y�X:0�'KdM
���-#d����"3-Y�c�#�*L~
��ȓLr����$Ï�$�dJS��$���6aq%T<DzՁ��i�0��ȓu,��s�����k�S9��9�ȓ%B>�y��[	8�8���.7 ȓr�l@�F�4]��;F$вs"�,�'/�@)�=T��؃ �H�T3s"�-|�Ь��#0�S3Q�D<+D�
�6�ȓo�` �b��&�{$��N^M�ȓ'�
Y�ʊ�q�l$��_Q�݆�v$���f�Ћbx� U��	"ʍ���?v�4�	�e�|�Iю�7w�0��аN�<C䉵|YX�I�`�\�
�S��0�RC�I�D��k�,!y&=���EC�I.n��aQ�5*f��@&J�j��B�I��I0�D'&y��{���s+�B�I����#�J>��R�g�֢=�d	�D�O�1���V		��������'-R�3aA*Ur� bc.uT͡
�'%��r��̥
�X�Ҭ3�a�
�'o�#1���D2`�p(	�|C2���'s>=�tǃlw��կ�(wQ�X��'{PL`�fUyt�u����o�T����9��Fx���ѐO���!�OL40(p@�K�� A.C�	�D�@h0d1xn�+���8��B� t?l�˶ꎸ�u懌>��B�I�h�6��]7��uХ�C�4��B��8|�Ի�B�e���UR�rB�ɘ�Y���J>PEZ�$��l��1��J�D�a~"��`�<���'(4h��G�<���	��
�<USf�'�R) !�'���'��#���ia�/G]}�O����m��/,��w���Qb�c��d؈6~U0��T��'>�Cg�`,��(�⏢6�%i�#>D��d�IS�'q�HP��G�h$�YSq.^ҽ�'a~"��;���� ��a�D�
B����>�Y��ٷ�ʂ	�8;��{��� �*�<	�ׅX-���؎*�BQ>�8�`�?��I�`9���ǈB
7',	�@���X��H�I�W�� 	��<<��\�ʧ��Oƨ�Hcű�t�T�s>Zq#�'`�̢2F�z� �1��>E��c�:
���'[��27���y��@��?!������� ���FqBp��A���%�A�;D���d��(��J"�3!xqC`;���?���DS�f�^P"7)[�
� !HGi��|��Ꟑ�&�4el�<��̟��	��(@_w��cL%#%��a��]��NQ ��;0�
�����Oz���m0"�1K�?#<�ӥ��a�KȮ;.a��,*]T��#��/�`P�0�ֽ���O(��`��X��F!*��{Û��( ��O����O$�`ϧq!�U���/`n�Cq�S6KW�}�ȓ+Oh�FFC,�µ��<.x���HObAoZş��'��\`��6�R{օG�R�}�g".�f�b���gb�'�ҏn����ݟ��' �PP�@�I�T(|�5Ɩ�,��5C�`�92�ԐCG��o,y��)o���p塑r�T��h�r������,H١P*ۼz��Y@diÀ�y��$΅R��ݼ(��r�Bϡ"�0C���*���	c�'{���a�T�ެ��KJV�"٣�'���Co��֪l�b��JO��.O��l�֟l�?)��Bv�闱��Q��ڴn�܅�T(M<�!��L5$��%ؖ*
�BF�a@�ښ;�!��k�\K#i�9�Pt��&].HF!�Q=7��B�I�&�4MP��v>!��[�)r���.�%O��m����z�ȓw��I�CI9�6�-i�aҡ<�I���#<��6(����l� ��$�5kw��iG"O���h�@��xB���y��"O��9� C^:���ɧ)u�qJ�"O� (ѫ�gY.g~��!��P�A�"ORs��,M�3����'�����"O0Ւ��0y4ܨ���K�)��В�茒�O�}��l�pm#d�|�$�ȇOKj1��� �-0(��>?��1�ʅ�X�"��ȓ4�N�v�D..��Rf�P�\ԇ�&�j@§&T��D�b�FR)�&h�ȓ����㠛6D7`��"nԧ"�����t�PiCQK� R�D���\^m�I�kJ���DذWC�e���W)�q*捀V�!�B�x�0�b�J�2^���$C,�!�d��A]\��dȑ�q <�C��J�F�!�D4-��-3�
�F �2�I�!��	l7@��D
|�F 0�@�\xџ��p둂�M����?��OY,9�C%��0�A�Č�sT=��J������?��3Ƶ�7N�8s�%�B��T�{`�)�R���	�hL��������g�?�D �y�fG�:.t���H�P*���1E�D0�g0�r��0�Mmب3���G����OҒ�&(i��]�C����cY5*�D��/�O��D/�)�w��l��ɋ�K��m��#ޜb5�	�|��I'.��!�c�T�r\�Cd� 
^�"˓�?1���?���T��H ��00�:�
�&�zfJ��,O��=�dͅ�A�jd�� �:���Af��X��5�.�%���~Rp֜7X�̓f���a�}i6�\U~ͮ�Xa&b#}*��$
+O�I7���}�z@�b�"t<3�#*?�F�>�2{��n�2}�$�a)V�~O�`wj� A���(#�>���O��}Γ%
�p���1#�^�۠�̿m6�`����H��_��-9�]�4a	l�$mՕGL̨K3jWA6�D�-A-��nD�d�/R��`C ��N�icG�>_���H���I���ɩ  �'�6�d��o�����Iu:�/O.4�×>��ӈ%J�	����N�^01G��2o��(�'`2t�K���<a�\m~BB�4d)L�H#kE�@���f�	H��L�O6��U���X1�S�&�1���=c�E`GA�TU`�� �~��C;���?�I�G���	�5�0��'C�ޅ�(�=����^���?ѧ�ȯ\�)ɠ�5��)A�jWh�<qǀ�(,�b�J��B�~u~�P�������O�	�����ܔ�Ms����GC:�rd�E��V�x Sc}B�|bY�\D����a��Z&|��D��y2*��o��`Ti��#���vN6�y�"�@e`���	E�_�!(&Ȉ�yB' R^]*2H������U(�y2���\���
���C��Ԑ�y��3��ɠ�  ���i��ק�y�D#����t�[W��P�F��yR�F�N9��E �O#������ybA"P�X�5C	u�H�PQ=�y��B~��a	��xT���J��yBK�?6�ïZ3#�9�CG�y2�X%(�ͻ6��ml:P ���y�!,����	�E�}35���'�B��a'�8FQ0=K!��t>�|[6��?j���TDA�4���4*�\��`(Ē1TLD�#�E�
!i��	P욜� BJ� ��`��,�`tF@��/ˌ<�䪠Hp������ 	t �Z} ��7kX*�q2 f�
�v	P��@�jy��K�9=ʒO��S 	̺� %��7��9��"ON�PcI2}eFx�4(�*2m\t!T"Or���.� jD�0!��ta0Y	@"O�H����[�"a��N�z[|l�"O���2�:snj!.�chJ1RV"O~���*�?O[�L�~X��b�"O����k�l
�i3u�YL�3�"O��Q�M��-{q��.bFtc�"OL��&�uI���"��YP�>�y�
�.Z�Tx)aKR;' �����#�y(Q� ���P�%�2&�
`Ҡ��+�yB#��"�F�Z���0lW�͠��@��y��:?|���	%i-��l��y
� �����؎Z�ч��&�H��b"O�H�A
qB��`OS�i �̠�"O�ɴ��@2�ib)#�P`!"O��J�7k����&�9m~
`5"One#6�ry��`�l11g�Aa"O��h �K�L�*pl�){V@p�"O�a��J����I��e�9[���"Od�c/
�F8����E���"O���EL�T�-��"B�h�pq�"O6��5D�X��Q���8��R�"OƙP�Jψi�IR3���O�d�@B"O����0R�j������
�4dQ�"OT�y���$������<A�
�i�"O�HU�S��EmF��j�"OH%��i��jP�옳�7�"�� "O�̡'��v^�� �^�2�R���"O�T�UIS1QX֌����(K�&M� "O� �
�?
xr�k��T���"O0ZD⋍]�����>9׺%��"O�hP���Y�
�jA�/81,�X�"O�@��]�Ag���@BX0"OVu��Þ}kRh[�*��2!� �t"O�(;CJ�K��3lG�A��0v"O�}#E;9�� `�,�*S&�xU"O��J�/�(5|v�B�+d|�#�"O�՛��<o�B{���NQ&��q"O�䨶(˵1r�� o�*E���"ORhBP�M:2+� ʷM̮@`��"O.CD:���2�Ϡy��	qD"OI�!e��#�@�f镞is���"O0Xۗ%�1_�j���j&,R�j�"OX�IƋ�hY�Hs�ɑ�=���ˠ"O�Ż�J
e�r�1	ώl��i&"O��2�7@3�eq���=�����"O��&(K�?��Â�0O�h�[�"O$�⒈)+�e�B�[�4ʦ��!"OB$[�`�5^	���H��<CG"O��h�mݗH(���BkT2c���"OЉ�Єݺt���pZy��"O�\�0�¼z8�D��<cil��"Ol! �I&ẍ܃!�Y�'QM� "O��x�J���!���H�t�p*O����C����)���"D8�'�� �U.�X���VdS�W�2�s�'����/1.OD��$�%W���'h�9#�[
 �}����?V��I�'�d��"��a^*x�ŏ���h��'�ų3m�IqH���*|��8��'f, H'N�4=��A��EN>�2�'0����7B�����FC*e��'���񯄫 � P�DJ:,8Z���'�8 {��ņ���)��[!<f�L�'����l����w���("���'�>�aPlBI.P�7`��2��!�'���5]�P𷆆�	90���'F�@����A����w�ï0����'�<9�3�)\t�LQ��yU>���'j�D�@AŲ|��kg�սr�����'���C��N=U��c��Ȼq m��'�vT�r�U���l1`n@
L���'�^Xb�K�Q2���d�U6uH�2�'��&��)��0��z=�|��'zhE�0)�|��t�c�R!E҉��'޼y�l	&�����u1����� ��&խk�*쳥��!c�X�B�"O���*=Q���&�	���&"O	3�OR�K ��35,���}�"OTXc�E�&�2�K�J/d��d�"O�@%	��}��;�(�a{���"O^T#������f��8@��q �"O��P1b�;b�ݲq�B�v��1P"O¹R�S�m�Q�B	A�@�� 3"O�d��	�7*(T���-�鐕y�"OΑP��J+	dI��-J�F�"OH��$N�I�0+�+�N��&"O~��ūC@f�˵M��x+\a�G"OBU�@��_om`�n�!V�HT"O���D��z�|��͘`�6"Ol�����J,��B5얛:��Y�p"OfZEI��vj|26$C/v|���"O@��@-��t���~n8X0"O� ��;w��]���8*��p"O4<�B�5tyta�$&4vNYB�"OD�!޾U�3dU�7��`U"O�!��6!��y�t�Gs?b=1S"O�]����L���x�c��:zMڡ"O�9���YLV���넛K�
D�"O���Wj\�
�xa�f�[%L�HC"O
h���9o�Pagh�<�D�R"O䥃 i8���)��\2��4��"O���������bRV�Ir"O�C�C�H	�u0g(/���B"O����
�,�($j#ݳM��0�"O��C��7�����DlP(�"O
E�A�-j���K��l���0"O\(���R�0���b��N���F"O�L�)I0���Pq�� .����@"O����AF��^!S�_��xq"O^=@��[.T.�T��6	�,�x�"O`yypJD0Y��@cȄ��i*f"O��!a �^�ġ(m���L9'"O4|���yx b�,�fpK�"OR�B�BѨ	�}����i�lb�"O���@*	�c�͒�iž/w�yC"O.��pLS�X��X�.�3)� �� "O�L�H�Pbd�\�-����"O~p`�=��x��� >�*�ig"O�Q�ݱJL)�,�$��E"O❡d����@�d�R�(�<@�Q"On�s����9k*|A��71���"Ojh��Ɂ 
�(��)F�׆y�0"O�%� ���ڬ�!��'�&� "O�hse�ٽ9�8d"D D�4�HV"Obh�  vbD�@ tZ��D"O�����p_�e	 ��.2��jխ/D�48Ti	`pId��C��TR�k,D��6kJ`_rM��	IcrD1��)&D�T����9�ba�\`A$�!�%D�`�`�۾/���Ӱ�*��la�i!D�H����7�,�{�C9+7�PˆN,D�D���Ӭw�*�S�B'�ء�(D��HEd�1���P�Ա��1�(D��a�A��,����U����P%D���Q�ÀcE.����c�	�$D�$Z���cA qp�-�������,D��!CI�.oʰ�dI�w�b5�*-D�T��W
m�� �]z��F-,D��c�n\Y�8ِ��UW:$22)*D�� ��d�v�45�V��g
,�$"OLT�d�I6D���E�<���3"O���7���K|y7a#P<��(w"OdQ��'|�5hE��J	4qp�"O��xA�uP�Ţ`��6@ry��"OP���.iJ-H�� 6�v�X�"O����V�01�@N*2�t�*C"O��y��9��S�ܛS͚�9�"O�4��� �nk(�ô�ϔ*��q2�"O" �j�
a�8"C��1ߠT3a"O��S5�^�u~̩�J�{�.M"�"O�X(ք��l��X4�����y"��-ax!!���b@ �U!ִ�y���KLLʠ�ʒH^>%J�b�(�y�h��0��0��G؈њw��yR��h�թ��G�=���8W��-�yc�*^*̡�˷5&�se��)�y��$z��-i$@1B4C����y�A��E�\�s'�M�e�ri�q U��yCA�K�������pY�C��y2W�]�H(�TC��X�꧍�
�y2�fL-	��)}��*�f�9�ybl
:N͐Ⱥv�l�-�&�U;�yR�^oϰ�K#Cх^Iua�I��y�̀�v&>0J6%MC̸�B����y��3�� �g��;7�F�I�� ?�y��A�y.&lr �۹1Eޥ�V��y��޸rMD5#�J˾�@�!aK\��yR�@=��<�`ދ�B�@P�۹�ybkU�n��`*�#x&B=hg)D��y�E,5@P�$�i���"�y�.T�A�j�c&F̜�P�iX8�yb��\��<��b�	'	�٤���yR��[I��ۅD��%��r�.T?�y��2`�*�(��P� Z�y�&��y���eL�l��� *B#��4�yr�Ɯ&�>b�Oͻ߲� ���yf !S��/R���,��EN��yR
�\��I���V�ը�(A��y¤J;�fi���U28����$��y�nN-0�Rxc����O����3���ybiߨ% PA��]�JỖN���y"������ܛqC���⁏4{�!�d��z�~а�+��C��u+��;�!�D�*H�P�L
���8�M��aI!��+ߔ�RF�:4:JM�g[�2@!��/u\��f�ҢVJ8��
7_!�d؝q�-J�ة@�P�8���hA!�d�� /Zh�5��7�:hQr���l5!�$S��P9Z�mU5�������Ly!�+6n	��ݸ�H2�]�Q�!������i�<AYf�J�h!��Q2!�����C�W/8�G"�!�Z�^�J�DY�\%���e�b!�D� 5{@2`č7�T��e�!��-Hƈ`��ݛv���h�$�!��xp�b���o��]JQ��$1�qO��)PC�G����a�3l��}���|2f�
SBh`�J�I0��#��y� ��kQ>|�Ι3&��Ӓ /�y2�&l!NuY�*"[T�H#I!�y"GN4CɈ�i!�I�	��A*����yBaN
{
�ᐅ.������[%�y�Z[�Xѐ�� ���U���y�D�,6�,� E�nz��sHF��y
� B� W�I6�I�u핍g��`&"O���VT k�@�"s͜0XTܬ`C"Op���'�x�`؈iA���"O�|�6n>}���g� ���R"O(eb���7��m��h�b�*�1�"O���!J85�E�BI�1�H���"O�!QT*Vdp6��(Օ�
hXb"O� �l����,ʐY��"O�U��Y5_=D��G-ԮYNLK�"OrHkE�
�m	-Q?�\iU"Or��(�r@��B��-hv�D
�"O赫���)��h �A#����F"O�x:P��%��k7
�,�t�v"O��{�L�~s�
%`D�*�؀�"O ͓G�+\�b�k���*�XP"O���p.�4@Ʀ�rSf�&%����"O�q��4Qn����4͊���"O�q�͒#�$9���H(qP|}�q"O�X�%��&���b��ΖiF�Ļ�"OJ�Cg�%~}qEʂ�N�^��"O��C�NR�4D�Ļ�ߤd��0�"O��ʡh)�A�s*��c"O $��h@��81�V��j�"O�	2����\`���:t���"O��3$$I �@�SVhݗYs� ��"O�]�Q
��HZX1Rp���<M(��B"O~�`����%���`�P%]1 �"Ozi��'P�gq�,a��P�7�(d��"Oh�!�Q�P[�a�GmƭJ�A#"O6�:���"8��"�ϊz�v�)q"O�p��+��*R���F]3}u���"Ox:bA�#����;�&�z'"Ol �!�Y��	eR�>�&���"O���߷�I�%��U���3"O2��#Œ,]��MGŉ�.�$ B5"O~e!�`��4@���b�=*w~0"O�x���ֱsd��@��-ZHaRg"O���g��m"�ye`��%F>�9"O��)%"Q ���r�蓰��h�"O�9`�@�"Fڜ�!AO�Q��xYE"OX���{�Fys�g�����7"O�h9s�"����E��F͛�"O�5������#V�T:-�|pKf"O�I��)O=(U� �p���r"O���B
3��Q��GO�W��h;a"O��3�� �lU��Kn�h��"Oh��B#�A��萓%N0M�����"O��
��+J����ϥ�(k�"ODݲ�@��f�*�j[�w%�"O|�����a�iHe I�'"O�`�T�a���4(�����"O�D�s�^�Sݬ�鶎ށ*pF5�"Ox$�ƒ�	���P/;`LeR�"O�MJ��)zD�N��x[�9Qf"Of�kwP?/L,d3E�8ga��Qq"O|�
PeC�Z��<����1F��I%"O��� ��|�[0��7d@t4�S"O��ɥ��*I!�0sf�-y�	d�<i"�
::��`&͖^���6̀�<�����q�F؋$��@7�`3��@�<���<H DQ�	-q�*�
�S�<F��Q)�Y����cx����Zh�<	�M��g�<�#ծ�'"��(W�g�<Q�V�#B�x��$�!$O\9�ue�`�<� �!`c��y>n ��a�%q�Pg"O<)���ۓH�ވ�gGKf����4"O2h)Vi,cH<���ś~QJ9��"O:�t�ɭ�58�K�"J�ő�"Oޠ��KV� 	�� ،>�8d"O`�j�$S&r��T@�0�$X�V"O��J�+.�����˒R�X�e"O�D��H<<̜���?�$�{""O��S�.�k��I��+sS�P"O:9;ň?Bp��a�ߞ|nK���y�(�.���%O�r��Áf[��y�i_�QN��H��9�J����y��Ι*ꮰ󥡛~�|P�*F	�yr ĂZOih$cC-x�H�˘�y��'	�� zc��
v��}SU��ymVz�X�b�Y�j�B����y��ʵ<ʲ�� L�`V��H�X)�y���5Y���A���r�y�
FX�}"��KmX%h���y"ř�+֨Ջql�7g��5J+.�y��լ=u��c���b�[�'��y­��eT���!�1U�� H1�y�e�(" ���G���$bU�P��y��)P�NY��mI=uL�Kv�1�y�*S9&�L��҈n	a�Ɣ7�y���� �� N��Q�R��y���d|���g������ND��y�$ߡm�Fݲ4�ރ ����')�y��H%.˲�
��ԡ#���ХC��y��G�W��.� �9nʯ�V���'�rWm��=�f��	,�y�'��A�8Hv�	a��
2����'�ʄ����)�H�cmT,:��AP�'/�]]��1r.�,�Xȳ�E��y�J\'?��C���s�>pkW�T��yBΎ-"�L8W�^뺬�Ū�yr�� *�Q��@Yْ 2▉�y"śH�09$��#;��Q6Ι��y�iV)=�PUI��\+�P�����y"�B,m����LW�p�K��yF|� �T�V�|�PPZ:�y`W%%���WU���0.���y�D(n>���'�/P�� C� �+�y"ė�B�\��"#��H`$!�3Cޢ�y�
L�x���2��h���y�`'d��PSj[�h�c$��y�JI�ZV�k�A)K,�X"�n���y�P>
�r��]�����ܔ�y�E� b�u3��5�lIاNW��yRK[���<���*ftl�gL¨�yrC�>��(�Rg֧�]P(T�y�I5d&,�a�F��x9����y�����咠�V�Z�*���y�C�$C��M���=(� Y<�y�m�
�(�����7�B��a��=�yr�C5�!
�<r�a��U�yR��f��� #	�|�,�����yBI�u�fPH�x�xp ����y2�TA���$�� r�N�j�-$�y¬U<y_|X�%ڊl�"�9æ��yB�ȈX�0������l�ybh��y�6�bp�kO E��;q����y�L��T��d����0�X󨒺�yoE��@0p�##����ck��y
� ��
g�X? �v�ct��?Rx�QF"O^E���X9>ԩ�3����jr"O��9�F�.�D�zFL׌V�8��"Ox|��� bX,,�H�52��,��"O���#6^��!X�� ~�*ْ�"O�,��d΄wT����MT�a�p90U"OhXro@=hf
�1T��_��|�c"O�!� �E�JEj6E��.����"Oj���:IMj���۳���s"O��c��]f�^�A��.z�|̨�"O�5F�Q4������Լ8C��V"O�dyuoәig��[�o��'�v �V"O�ahe޹iL8��p!�O@ �"OXɸb��L��|R2��4R�Y�1"O�P*��Y!t�2�Q��S��ۆ"O�=�/1uMf8�G��Dp�]r"O�X����:2!�D�=��y�"Oph������i ��[��Rw"O���R�_�*��Re�U�	�n��"O��je���0�(۷F����"O�5�cCҖʞ���%�� QcV"O�kY�i�i@�T���"OH����4����eO
�:��T"O�1�rb�%�]!��upЙ�"O�i:e��F�)���h�@cE"OYp� �!'�@���@>ON�A"OF��&�>��F��9 �R�"O�Ei��An�q�fr,mSa"O�pAɒ�vnް��>x��a�"OJ�B���p�e��L��|�^,��"O|�)ac� G\�Lh��8��\Ӓ"O�h���+���"t�T�p�T"O��1�@�׀|ZG���A���"O$Q��0?�hf#�UK"X�"O�I��a�zS�r6�ƀV��0e"O^`ja�F�n� �;�ֽ���"Op�J�<]
8ɰ�ز:�ȱA"O�QI���"oM���@�\~� �"O2�h�H@��+�ҝ\|L�"O��jT��@鴉�a��X|�ա3"OL�"	���dz��
(l682�"Omh �+4
�R'��c`@p"O�Q0���!ކ��h��-���q"Oz� .�6b��C��13�N)@s"O艻��Ǔ|<&�H@�]���ٗ"O��w�
] sb�0o� ݂�"Oޡ����J�kO�%�Ƶ�@"O�}�2-Q�,��@�(�,{�<���"Ox��Ckзf=�pBU�7$���g"O�u��U�A��8���H�r>,�"O�Њ�Ⱥ{KN����1vt���"Oh�����2��K�䅧A��U"O�D�%� G
���PK��X��Q��"O�`��**y����Ä�S�&-Q�"O��q�'�-0ɺd��#$�A�"O�a�0+MuqY@Ϧ8BB"O��	D�	�4�V�@��	�3�l�:$"Oj�IQ &b�`�c� \#w�@�"O���S�ՐLk��E,VʅRW"O2y �	Q:iQ�$G4A_�!��"O$�����n���3v]
[�@)q���# �9"퇅<�np2g)����'�@p+�EE*�:%p$��u=y��'��3�.ߔ���i��>r���`�'㈁3OFj-����^�\������ ��`�nx[@S�A�,�`�"O����˰,��Y�f؆&@��"O�v��:��}�V��)R7�xX�"O���A�������P�>װ)�"O�|y�C�n�۴#�;g6�e��"Oj:�M+�i#,hM,hs"O��+ЍZ>u	���AkF�)W��Z�"OJ�[�T�!j~�kpП��9�"O�� ï� G0��c���-��j�"O0�b�E�(I�Fb�.?|���"O���5D�*"�BDP36���g"OEhQ��)$d�����+����e"O �	�#X��1Apb��U~Ρi""Ot���#^6*J�����W�b�
�"Ov�¦D�N�P9反M�)0�"O���R�i��=��X�dR��"Oz��#9\Q
��4Ml1(7"O
���ȷ!n|��B�jR��ô"O���'[�n���c��ѓ+���!"Ol��c#W��H�f&܉%�j���"OL�P��T�;V,�gc��� 9+r"ONd���k���p��=#�d4r�"O|�;�E&2�ᅄC�Q�L��G"OL@��l�e 5�٢AK���"O���mּ%�^�զEZ\��"O��A��W�`}pĩbh��
$�"O8�`%�L:8�XUHL q���U"OvM3�&K-M/$Yӵ�E ]�U;�"O�,�f)�0�=q��/@�l9p�"Ob�xB��\`:�:udɐ<���"O¤���^�]�u냌��o���d"O��0��<(PZw*í�� h�"ORh1Ѐ��;�� �����h���"OT�P��@�w���1Kɚ
�r�3"OȰ`�<xB��s���I�"O����l]<�¡��w^,��"Ou�fß"f �f��e 8�3"O����CTP5dP; #|��"O�B"n�;N2<�kb��7k@` "O�!r�M0�\�#L@�TZ��"OzT���WJL!��Ҍ"`�ɱ�"OJPbCK��]&�k@@ dh<��t"O� �噉���<� C�l!��o�Z���m��^�)��<Dl!����8!	ء^X��Еg ��!��&a�.5�r
�a*�E�b�!���	p��#G��)IB�.�7 !�<yE6���:Ep�RƍXC!��		�̄:��M�(�0]�X�@!�	���]z��+��1"���B�!�ć9^>+"AͿ5zi�2

jw!�d�=l<�8iQ�,���{4ɂ�:E!��LgFB��fe[�p9�)@v�U� G!�Ě'KV&�ǆƫ�hDS��P8W:!�䗛E��u�G�F��.	�W�!�@�OX�����+E��P��o�!�DI�|����{�H�P
 
�!�D7SD��##Ő�P���$�!��C���iܼV��eY��� ���*Sz��(��L^F��G��yr��d�̐�GK�!`$�ٙ�y�j�UL��BĝJYK����y�/��ql�M t�ǭ9z0�i
 �yBB<B\��X.��2���
A�\��y
� 䌩a�>���1"eԠ,Li��"O�Lɕ�	Z�t�7��?Q
���4"O|�"�~�E�gQ�H�b7"O�AWkIv���C�R�Gb�s�"O^���R��$�s��8<���"O^�z�HK�iF�:�K+\rT"O����I<=Ϊm�4��\l�`�"ORI9c��32��AB�-�fH'o���� 2�I��&��8���4�yb��[
���߉�$XR�jс�yb�J�-�Q1�
��!�S�R�y�C��q���&N����
��y�!�C֐��|tt��g��y�I�O��ۑLso�,��b���yR���-�4���+ڃe�|���֊�yO@8�R-\�o���Ʈ�3�yB@D�B2�{!�%=F� �qᇳ�y�#�*1� )�$,J.�����'?�y� пT����k_�9��`AT�M��y�aI/�P$�e�ļ6��x"H��y"$ tX
l0��3UN��1���ybD!aN<A���Z�;.ti ϟ��yr��%w������Xh(�r�9�y���/:}� �!dѸ|��$��y��@&&��1�c땪xh�$P4e�y�ɜ{�(p+�̐7�������y2oذ�H�9dg�	"�]Bŕ�y�J�3%�e���4O	�Ћ F;�y�ɂ!P�z�: �\���K��yB�J2�0�(�V�|錩���y2���VВ� ��x�NX	v�E�y�U�<1\0 f�i�h컵��6�y��V��$p�5k._���@��y���zE,�v̖&V.D��AlO1�y�}la��Cd0���	�yB@�8/�b4�/PR � O��yB�Ln�X A��A���C�̇�yr�	9��!�E&/�zՠ����yIY����b*J�S�yඥ_�yrmY	f����	�;v 0�#�R��y�+7�lay�"�>!J�麶=�y��]�[18�#��,g͎�	樍 �yR�D�[��hW��n����&���y�:B�ԓ0cA&2�T��bN��yB��<��QPsD��/+��a�i��y���U�f�3�,�&9J�B.���y2n�3}.<���̄*܌t��C��y®�+SR��GN����+�]�y��+t�4��HD�ek��G��yB�Η?C���� �m|�|b7���y¡��h��8�K��^g"�����y�
_)#�޽q���\؜�j���?�y��Z�PJ�$\�f�Pvk�y"j9)�Q�1m֜R�e�F���y򣀫�X���aE9Q���YH���y�hPu@�����!2�`4+eN�$�y����2x�"[ '���S$D[��y2$�I�� �QI�:V���;��Y��y��<X��H䌇�#���9�/J��yj�r��HH�Ċ1H��3d� 5�y��ދ\{���@� J�	��_��yↄ7.��XvH�3Έ�6&��yb��)�@d�W#��<� �K0�y��\���A1�"�0���#�A�%��'��z
� v���̛�51��\���"OF cF�6��Q�Ȑm��f"Oh����'U�����f�D\�t�e"Oj��d�Ǘr8%AfeҤCO��1"O�q ����W��1�*Qm��M�"O&@4I�S�����o�7va�p3"O�e��/���d��4$���'"O́��X>����[�,�h��"O0��lV5*��p��b9!_����"O,�V��nC6%��G�HZ2Ei5"O����+il�I3��(`F�I�"O���"!�:Z.��a�b�1x�|!�3"Of��F�0F�؈疬?�<���"O�gC ��@�(qKI�j��\�"On�a�aA�f��҅DJ�jvd	�"O6aJ�C�Z<���x�xq)���yRԸ���)Ý{� �q�@	�yK�6 8�Y ��[���V�y��*?	��C�P;B�&mSET?�y2��D��%�o�?5�>��w���y2��]5t�ɧȀ;^���)g��y2)#_���1D+�P����y�f�.{~n;�OG�3v�(�I���yr+��.U<�Q���Pɖ�	�yR�'-�P��̤x�!�H�0�y��0���2̓*ǎ�r�G��y�*7`���,s��+n�y�)~薩��^�e(���#Ƙ%�y��'~O����i��^_*�*�Ǆ��yZi�I�p�ټvFD}k��,P1�C�I�j˶��kT�K��),f�C�I�w���z�A_'��3�A2��C�+�&�
�lʐ� ƚ�z�C�ɉO����B������wi�!!hfC�I�I@�!ebH�E�����K	)(C�;i���EB�bzz�$K%TiC�-*� �VĖ�B|m����ۤC�t�N�H� �t\�A2�D�UuZC�ɟ]k^@(���NH9҃�͌t*C�	�R�0!@1�9#O����e�vC�	�? ��W.$�����,�C䉏y��k�"C���8#�3=��B�I
	�J�'O�_3�-Q��]=�B�I ���R�Ȟ'8~	��� ^��C�I�!m��*Q`��>#��̽H�C�	D��݁"jŪBfr�`���eu�B�I9�`p1�l�D��"�
(l��B�)8O�Ԩ���!�((�U�w�~B�	�t� ��A�X5�i�A-*vB�d�"��A <��AF���tHB�ɐXK\����N�`�����>X��B��~������PFr��B�W�B7�B�I���u	Ԃ�m�"qq6)�ͨB�	�c���� '�Gհۄj^;�BB�əO�ru"v���$[�Ab ��qC�C�ɏ���ض��n�D�� Y7�C�	7l���F�0���S�-�la�C�I�}~l@�udɉ3�2���=y�C�I�_=`�S�F�2�"a��bEpzC�	9�؄���ǐ��y�j�3;ӦB�I(H7.�bM���(u��) c�B�I�A�T6/��#����`���N�nB�IJ��t�_F�dЃs���0�^B�I,�
!°"�HJ���p-Y�3�JB�)� �h��鑁;�l���HQ+ RPU��"O�8R�	t��}""��-�v�P�"O��бoǉ,@}:��΁r�,r�"O�L�+:�V�S�ʰ[v� �"Op��뜓x^i�g�C/��0yp"O$��PG�;j��� C����8z�"O�����|�H�P"�
#?�HP�!"O4��"G'({��#� �� �L�c"O��'Aދp��l��/�?0�6�2"O��˟23\�(��nVY�H@"O<����R
�����;G��mx�"O*e؃�	_��M��K1v&lI�"O���b���0�W�\�<uJ8��"O"PPߣ<z��BJ��[Y�A�2"O�}�%�S��,ʑ捑@A5�q"O%�/
Jb|�`\.��S"O؍5k��tȱə� �08'"O�!���~Ҩ]��o(O�(0�"O,�&G6=v�Ö(�!%xX ��"O^�8�	�&n�F��(��I�U�%"Ol|rrB�%9Rn�Ȣҟ'}h,�r"O�x􅃏A�����	Dp@�Q"O�d��8�
�gț�6���"On�k�i��0.l}���x����"Ob���j�::�Ys��_a�D#�"O�}�5�ӫP%*J Ŝ� c|�� "O�p�g �?,��`��GC��8�"O���WB�&I���1C��+2biz�"O^p��썂!N`�%�T#V���"O�5��fH�V�ldRb�?JP��7"O�̈���Z��@� �h�Ԍ;�"O��c�-C$l/�Ղ�@�<%�
q��"O<�D��$c��4���2(��}�"OF���.��.-��Z&�Q69��"OΉ@���YVl���%G����"OJ�q�(̮|�&U&)� �԰�"O�{DlB�~�|��Wh_�S��c�"O�yj��Z�@��X�����y����X�h@R"�i�t��fg���y�U��d��Ɖ�eԬ�2W�L��ybde�z��O��^ �{U+Q��yRIh����W���W��y�-W��yҋ��L�Ri�JR�L�R�XiU�C�I1a�͋% ֏VWN��J2n�B�	�>�ի�N�d��cB�2 �C䉏S��e!VI��s���yC��xNfB�I�J�P!�F������*oXB�}�:��3/��Z�g�hG|C�	�ML3rNʅo$db7N�5W�C�	�@�D V�֖J�.��G��.C�	��dm���W������aͱ2�C�.J����ҏX+K����A�&t�C�	�u�z&�p�*pMªtCvC�	2Ap0MRDj	s5��CV�bPB�	��*�3v�G�C�e�vC�I�,��|�]�r���@�-G�C�	:��cꟚ5*$!��b��](�B��,��|������$�'#$(HB�	#���zԁ�j���&�D3�zC�	�5*���^14:�1E¢LDC�I�HlT��-l����A/}.C�	�s���M �
�2�aI\�~NC�	��H�&@�7��a����LT�B�I5�ހ���:������!A�B�)� ��qsM�j$ ҵ`V�n\݊"Oz�h��M.H��y�$�\rU����"O`�a���
dh����V),U�X�"O���g��
&0h�\�B6�[�"O���s�F�R����mP�zD"O�\9uj�O��i�n�&�r'"OJ����?`�6%�Gf&@�8T�3"O`,����8Gf��5�D`u���"O��3�=)��Z�/ޞ7j��"Oxm�S˥�
ҴΉK`A��"OP)��k��"4:D��e+8E��"O���X��b�FcO<M ��{"O�th��d���\;w���""OJ��/ך�6��
4l� ���"O�j5�:�x{&ɉ�\���$"O�9t!�!;���)"�\�X�uC�"Oj�j׭
�~ p0q�_}�L!�""O��3։��}�����/e�
1�%"O�ly�C#U���o�#�B)�"O.�BWE̩(��xc�A�A�<)�"Oys./�2Q�@c��@/@��"O��ťV�C{^��="-���"O�ٻ�!��|)Q��-#{����"O��j�O9g�� $�X�a�n"OpIpmI=53��I��J�ѫF"OB1K0��<�ȥ�߽d;�a8�"OqtnK��ġ��h>&&�T!d"O��ɀ�B:5�j�@�F�`�X�""Ov��@��+W	ͅ�q��"O����B��V	L%qʁ8=�"<"Od�X��_%AqB�Ys��Q�1a�"O9c��Ef�"�L�{�9B"O �k�ᑂ[Ir=k��A*,�g"O�1B�@�)W��,���T�e���"OV I�kU?���3u��9PT�YW"O� i�ʑW?��@s�
L�D�"OXK���> ����G��|ɣ"Obap��2`����al� �J�1�"O��b�wRژ�`��*�Y�"O��4��D�e�g)�&q��j"O�-a2�Z4{'hib5	��q��Ѹb"Ot�`gΟ�W�ٓ�۫b��#�"Or�A�˜07�l���eۥW���1A"Ojӌ_�HC\=�ႇ
sU��be"O,� 6m�$z�|7!��`Q�08"Om������sU� @� �Ɂ�BE�<A��	$p��)�cz�H5��I~�<1�A߅R�����R&J��he�T}�<�DJ'|�t�T�J�Oj*�(��{�<��bn�E��D�d������EB�<�GnٵN��p�� �=n|���@�<�b�]cc��ǌLB���kV�<�o\�Y��[���a��#��x�<9��R�h��bޅM�NQ)�%�[�<�����\�$���C�jt*B�^o�<�'�͙@�6h�K�K���*��o�<�4+2@D�3�L�#.hFM2V�n�<Y�m� l��I#���s\^�:5#�j�<��ꜥ(���$�@8�` �l�[�<��3.�Ԑ��_4�P���Z�<�@l��LM��#X�T=����o�P�<����RT�|鷄�_����,�a�<YF�"�@z�+�M8� ���B�<)�lԶ3����^c����C��z�<� 
\��L�@	ȫS@V�_W�Pb"O�lȣiکL���v.KX ^���'k�eB��_V���q�E4vÖ���'�(�)ҫI�U�TPS��d( ��'j��(��$KVjӔM�bd�'��ɣ��ҐfT��T%Ƹis0D�:�aR8��L	�� ���ps�.D�hzq�
4VQ��O��d���f'D�tb��R	��� �F!D8�%�ĭ9D�L�$NΝ�2e�!ƢR�����7D���M"kf�����E��nmA�./D����eQ
��(�.���é?D��Sé��c6`�E �p9�)	D?D��Q'԰��My��Y�N�~�1�2D�$hP���B�Y�D�\�x|m�A�=D��U��y�������
vI	Um;D���{[1�v�W�u,Q�c;D����DU8q���CG�(^ف��8D���ua�5u�������5S~ޤJ�d7D���e��3�rk�D�R" �s4D��%��n�-��.l���X�1D���N٤S�8�q.�0X�uxs�.D���	�7f���O�2[m�s/:D�$��O�:8���h�k����h�u9D�h8�����9���H"�v���n5D���R�̓y�Jũ�%L4"�0J2D����%��
������+$��./D��y�mC�(�C"'K� >�
�j.D�`����A��d0��	4D�]�pm1D�`�2��m��i�7.O����/;D�|CC�u�ٜ|�l��$?D�0h��:V���9�׹B m��N8D��ɰ,�-��sP�T"-X򬒶� D�3��5ɉ3-X
�Ę���>D�`xr�U;2#��G��n�|�o9D� B㉓^F6����>NX�T@��7D��'C٪�`�M
UT�5b�5D�����~�%��V���b&8D�Ljp��TÚ��Ղ��aSr�@�'5D��c�8So�$��.S�v��Hâ(D�|����#L@p��� A$6�x��)D��J��iva�"�ҖL��[r�&D��7��<7������S��P�*(D�P��lY��D����nLH�q�K&D�(2 B\e����&
%���qe.D����/_�.2zL�v�S,朥���9D� �FF^{�4��p�Q O�dmxҁ5T�4�3NJ�BM�k���D��X��"O����e�����j�n�"�"Of(�Ecǒ�Z�2�E�S�����"O��3�.*�fY��l��k��"Q"O>��%�Ґ#�J�i���)1b@���'4��6��(���ʴ�"���
�'�0Ai:Y����" �c<�	�	�'�����L�*Bʲ��@B��S'���'W�M��'
�t:<�����E���9�'�J}��f��s��B�f�h�'x�Ȟ�i=���O�bU3	�'R�X�R�&@�E",ڍ�|��'��mq�a,vY
 ��͞�'v�hR��O�K��2*�bi)�'p��)�M�����g�S#�%�OH�<����wZ<�bUkþG<{�fCA�<�b$I�2O�y�
��\$�@���� �x� �Ox���E�'�N\�5"O����߾G����«{b�}Y�"O�|�QB
&�i1�,LG����"Ot�_�b���Y����f�bE��"O�zs'cn���W�Y�4�\e���	�P���	OΛ����L�Lǯ%
����͑;jqON������s��8n}�թ��/\` �O��)Y�2���` ���*Њ�Ĉ�N�
�{�*̄\���#̍	e��А7��4X��'��}�����aA�E��x82"�O���R�̦�M�8:`�"W�]�DB�闤
��?���Ԙxf�a���cRc_+o��i���B��p>�0�i66-~�\"v��	Z8�ё�/0R�)��O.��R͎���lyʟ�O(Ĺ`fD��~yx�Ý7	Pi ��*�8�R�y�:��5'��j ���!�S�?��گZx����ꚨw����NDU�fBKV��k�G�e?�I(k�,�	D8�s�9X�A5 A�Y:�k� (�(�iu� 0�6�'BM�<�S@��MC�"	=X��t��RRv53�I�b?i��hO�b��@E�:68��+p��IK3�*�Kf�&n`���?�@]���̏J{��aC/-��	�U��3�A�M��_'��i҄�J�҂�̯0𜻆����pq`4-��|:S%�"_&���\�'�fY�d����KP��vu��(�o��5��`��5�dP$G���){���<�@f'��q�u��V���cևer]�[���'~d}�����O��}7�qʡR�i{4N�(����7O�3�?#
�z�Ϫ*t��a��i����h�Vc�������l��p@�f3n�{%$:�D�,�'X0S���?���?i�O��?���?� 9D�h����U7v���eM�Aft��I�?v�=��!�3m�$R� -�I.�h�*�4�9���Ʀ6șе���u0؜����l�ғjehD4�I� lb��t��cbǏ���be�
�.)����`����c�S��]6y�MX�D�'��H	��\��~�$"�S�O�l�Rc�:R<��q
0
*���'��7��OHʓ �n���_�H$>I�!d�>7��j�F��T��	�:��'���G$]T��1��y�8�p�Y5[�*xΧE�tY9cK/#r�e�a���PJ1Dzr��t� ����ڋ���G��$9��Y�Z`;p"�Ih<�xYУϿDڀ�Gz,��?A�(v���'���t��*Z�_������Q������������7-.I�Y���iV����]�<�|"
h�z�m�ڦ�@�[0�Y+ab
�
���C�������M���?�)���+��O<��n��m���ɡ~?|)8�a�~nB��wo�21M^��\Od���S�҆+$Y�$ʋPZ(���iy�}
sc�bwh��T� �`7�T�u{��(KcK%'�
šB�B	_ˮ�Z� K��<�~��Xc�"���Ux�;Q�ȓy,oZ�#B��D�ONUmޟ�E��4A�|A�䮊%t��������?���?�.O���6�S�J��ȲfDU�QrxU��m08%��<y�i5j7m:�$�(םQ�|A�'�8T�)�� ���٨N>qۓQb�D �  @�?y�n��3��x�$)_r;dH�7�_��y�́/b���qɝ�p#�ݘ�%�	��$M��y"�� w�J�����d���bK��ըC�(ۺ����P���@�ϧGjON��p<��m 'M�qb�ԙC�4�e�Bg؟Lџ' n�Ir�@5t�H�NJE/����'��8�a��9^�c#ɂ<�)���,�'%94FJ
�[��"R�͞I����� �JI��e(W�t�2�/�/U/T��=\���}j�ϑw���rCT����
'!L}�<Y�V
"�DPG�^�|W�I�"�v�<�o�v��� ��`���U�Jz�<Y`����5��9	P����z�<�#�.�D0�(&X~�B�s�<Yba�!t��S�t��c�e�h�<�����!Ѯ$�L99-^c�<�-�!R��K5ӊ�Ц\^�<i�D��L���d��1�ֱe��B�l�`�F�V#0�D�<a����<���O�Ɂ��A�-��H���,0�!��>=B�I�gɕ?�R�z3�,0Bў��ᓿg�Ș� �o��);���KtB�	�C��}�	c4�m�#�BPXB"O�9@wD�|���nѱUjH��"OR��v��9P]
BCAVd
��qY�p���R��b`&�~�FԨ�* � F�B�	�]��r�F^�DxQ0J�/L��C�I7<�m���3i�t��Ϻ��C�I�oSV����A.}+��S�΂e��C�ɇP�A��%X�������,L�C��5�̻R���p�
F�+Z��B�I�� }�M�*=�lH	ԭJ�9B�)� �=��(0�}�W)/eF8i���'��	��^ Juƕ�yDcE�:epB�	�_��8� �I�&�q�G'Rt6HB�ɁOO��)Ro���1�ӄ$�RB�I�X�<�p�� f5���6�%$��C�	�Q�Jl��(�XL��o�'�*B�	;HPA��e]�nӲ��"����C����0Q����|� �<ނx�ȓx`�X� *�"M�y�7-�JX�ȓ!W�P�����e�k�ԉd"Ov�1��٢+4`��4.��{RTZ"O�M�UM� t#�kP�D�Nl�=xW"OTl�$.ʘ,t�n�"D(="O8ly��	�$����/(.��"O���c7v3:eC͙�)� ��"O���E���U��p[��E�n5�""O��F�("���o�w��$�q"O(��H7'pqC�-�/n��P"O��b�MV/QsEh#���n* "O���a�(z�@" J�]4��"O)	�G�kH��Sk_7"ع�"O��Q�!�Y���[�LC�'�d�Zp"O�P0��@Ů<�E˃�'�T�a"OFA�e�X�#L���SE;3�"OZ9[��N/`⺥�A���MCx��"Oh�k��1mS
eSZ�!"O�!)���	6et0F�+Pz�@"O�t1��� �F}ӏ�7Y:�PPQ"O�tɇ/�5{�v�u/I�Z|֘��"O���7�E�w(�I�`%#�"O.�C�@\�M���y�E�'3��1�"O����`ԧ�Y	3F�*	�ƹ�0"OJ�`��U�l��f�.x�Rs"O�!�� I�'��j��K�7_��آ"O�S�� J�۰P�3�>���"Oq��[��ސpQ��W�4�w"O�̩��2J��#��5.����"O�ã	�?$����N�C�L D"O`p��A	7��]��L 0U@���"OV�(qEX�mH��0,$p��)�4"O��B-�-h���v�
�fg�-Ȅ"Ol�I����Ok��5*�\�r"O)$f�!f�kW�&k�qP"O��1�4LY���B��,k��xrR"O����0g��
+ѹ1|~$7"O�`�Դ�zp���'d�e�"O ���$Xh>��� O��#�"O�0#3�ʠmKt0rʗ,<�Q"�"O�2�Y�w�tR��3If�P"O�9��[,�� ��J���'R��y�-ʕN2 ��Vn�1�U��;�yDVtH�k&��F���G�M!�y�E�ux��ቆ�E�H�7cN9�y�,�cw�<[�d�6����2�yB(�8��h ��=00��P���;�y�vڤ	ʅC�8+tР`#���y��Q#0]~ �1K�/*Ґ��� �y�$�16[H��2 �	&0<L;@�Y2�y��	NSR���
��>|�����yR��(|,��������[����y�Ɠa�ʰ*����UR����yR�|��Ě�]w*��ra�>1�!��H�&!D���tD <0cF�(&b!�T2
�C瀐E%��x��.!�� ��D���br��(A��c�"O��e��k�&T���N�,��"O�H��'R�lZ9� �m�A��"O����N$}N�:PoF(U���5"O���Ӕd`dRF됫QH$p+��'r�'���'���'|��'B�'���O�\	4��-�$'�mb��'�B�'�"�'�B�'b�'-2�'�b@aE��$cdzMƻZ��T�'{��'�"�'R��'Ub�'��'���F��*��CH��sIڄ�'[R�'���'���'"�'"�'U��Z��J�:��b��L�ܓ��'���'s��'���'���'F��' Ph��S�X#Ī �-��dЖ�'6"�'l��'="�'��'�2�'������)r�����7%�P5���'A�'���'�b�'D��'�b�'�j��6�:{�Z���M9��銣�'l�'�"�'���'���'��'bFM�2�Ǭ,�Mڡ��S,���'���'q��'"�'���'���'mƍqd�C$/4<<*���	�.,�#�'(��'���'z��'�"�'b�'��гj�ar�Ҭ��?(���U�'�����ߴ�?���?����?���?Ѥ�D�}�"}��B%�2 y%��?!���?���?����?A��rٴ�?��u"в�I�V�W�j���s��OR��O �D�O����O&��H����I˟��l�&.��K�G��z$� � ����Of�S�g~��~�,��ƭѢW����R���E��^�u��O�mm�p��|��?q�O)ش8K3�	O�V��&�>�?��h��Hݴ���b>��'��#"�h��/c}5h� /�c�0��Gyb��]W���#B	�KmA���O.*�p�`ܴR�L,�<Q��t�k���Clq�v�
�9t����̙7�����O���O}���ͧ_��1O���BR�[\s��4p��5O<牵�?�A 7��|J��wo���`�\<x�E�=>xl̓���)��JΦ����!��z��%F�/1 ��pH�9@���?A�X�������͓��d�
%|�B�� ZS�@!iU#b4�	��c̛�FŢc>��s�'Ģ��I?9�Z�j���x�z,Y�Ə>|��'��ϟ"~�f��e��E���9򁏚=
��̓8m��'���D����?ͧ:f�J��HjxTꃇ��J�R(ϓ�?���?	�#��M�O��.��Q�ËC:x��"6�u����1g�:�O��|J���?���?A�%���c��i%h���q<��*O*Ml�*AQ����ԟ���v�s��)�A�8=X�F��P+���¤*���ܦ���41V�����O.���D�}Рԣ�H�h&,D��Ǝ��ӎ˱h���¶p|l�*���1��.�w�		���D�b��:r�B]~���Ё�"�>�$�O����Ob�4��˓Q՛��Ýr$%G�g;����������6�y��j����O�QmZ��M���V9��s�I�#�6����"[����9�M#���� [|����<l�)J?y��wTi:�	Ʌc�b)�3�W�!,6�ӛ'���'�B�'�'��!X��R:���{��8*Ѹ ��O*�d�OhToZ&$��H��|B�����s��#x�>�����;{�'<����T�׹C%�V��xvBǻR�ȫ��(ro�M�n�.�S`�'�̄�'��6�<ͧ�?���?��n�d�*W�Q2{�}W����?!����������tc����������Oܪ� ��ܞ;s@=3Ʃ��[�,��O:��'���'�ɧ��<�NH�L�m�x�S�(.+��1`��ε:�p���LkXw}���ɶ0��i�IQ�F�3l�Ƥ:"	�8	���'Gٟ\���|�Iݟb>�'�6��<E�L<[���658p1U�ݲQ
,ʥ��O���զ��?��U�(n`	<���,��:7�]�h�64TZa	޴�?���.�Ms�O������ZL?��B��V�R@�{A�_g���4���O��D�O��D�OT�D�|�� >8\���E�����{SÕM9���Lv��'c��)�Ӧ�]�o�Ӷ��^�ʱ��
/������M�yJ~���8�M;�'S.��wJ׼Wp�!�3��b�t!�'�v{���(�P���ݴ��4����,a+t����`j���G���P�����O����O��<k���ļ5w��'��I
#�H�A�֎B��I�Q�V�T��Ov��'�'��'���ڵ��2�
��]�f�Uh�O�e�h=��	������\wp��IT�b��(@��%1�+<��lxC.��"�'���'��S����yR:��%��$���KB�(�4d�"ԉ,O��l�N�Ӽ�X�!	(Y��80��[&A*d�	��n���0�֦��'q�fi��?}h䃅�4��R�B@�ڵq6D͋?副�M�.O��O��D�O6���Ov��udƷ(|<�d�B�i��r�<ɓ�i~P�['�'���':�O��¹}A: �ec�jCj�i ѳW16��?����S�'~�,�'�/O��+q��NRN5�U�D"XrLe�'��Lj�� ȟ���Y�p��4��U�R͜]�E��3%P�%��>?N,���O����O��4���8���mP�'�¯�I-�hPEg�5V�H(8��J�2��j��⟄�O����O��� ab0!��Y�����5đ2,����n���GJ��xw���O������� D����7A��"uM2m-��1$2O���O����O>���O>�?u���T�]1&�±d��V`�A��BƟ��	韜�ܴG�]�'�?92�i��'ep�n�"
e��+3����Sp&7�d@�]"��|R����M�O���#`-N�����ڻ3��Ava�n�ܪ��>�O���?��?��x^� ��!q&��,̺�L���?A������5g ˟��I؟p�OX`�aٞKg�	���R�h�{�Oi�'.j7W��IN<�O~l� ҀfDeK���E��1;��= >6��&�7`�i>��t�'�X�$��	�C=d4�3��Ã'�5���T֟��	����I�b>��'5�7�Ɠo!Ju{��������g��*�,P�"�OJ��Vʦ�?�"R�X��4.��������J�"<R���3���@�i��6�y�6m0?�妔�E�0�	����Ya\5��ղ;�Z,��f�>}N�D�<a��?����?Y���?�,�>*$TV�%) l�3:�d���[� ��������X&?��	�Mϻs�Й�4�1�p��[!F�`:���?H>�|�Ta�/�M�'��M���4<z115GK@o�M�'�As�ҟ� �|2S����a��Ҋ~H�ȁcS6.��\#V��՟l�	ԟ��I}y�eyӰ!(�I�<���6|�Q�u��6:�(��Ui�S�`AJ��ľ>���?�M>�B��
Иy)��Z	I� ��e�C~Bl���:u���K��O�8e��uZ�ΔJ���+�@�4B��6���'���'�������,Pʮ1����CZ�Z1F؟��4v�\�b+O�o�}�Ӽ3!;3���Ah�$-1J��<1��?����,�cߴ��dJ�Y�����q줡Ñ��1ED09�难f}V���n:�$�<�'�?y��?����?q��#���y��{����8���Ѧ�@x����ӟ $?�	�o����j�N�lx�Z)@
�Y��O��d�O\�O1��p�D	Z$���+�Ľ>;育�nݑ�ܴ��d�.��T��'k�'U�ɫUHʕ��`��Ռ���OZ��m����	�x�i>M�'�\6�Q�f�Z��-�*]����G׈��ŮH/E����a�?�tY��ݴB���Liӄ A2mXpxܲ!,M08��f��7�>?�t,.A���>�s�k\�,;�Y�S$,�*��U;+m�D�O0���O��d�Of�D8���v\Xf�Z�Sg"� �_*G��(�I�� ���M@���d릉%�\C�˓+i��q��h��D q�I��ē}қ�d�󉚸-��63?����'���A�ܦN>���'��(�x1��O�m�N>a)O����Ob���O��׮�&V�ȰYagFR,<���Oz��<ɂ�i��)c��'|��'��57�H ˙) yR�ssB�$K�ɷ�M��iO�l#�#���!7�r�F�� ?n!��N�5l�$s��sy�O�*��	=.��'��%�7^tȪQ ��J;w�8�;�'�R�'9r���Ov�ɲ�M��FûkKf���M��s��+��̀f�f�����?!��i��OT��'��7S�_��Q#1kB�0�0Ы$m�O��mڸ�Mc��	��M��O�Uc7��&��$m�<�v�H�7[�ڔĄ6W�0��F�<a+OV���O ���O���O��'��3]�43��KN�TP����M3�����?���?�H~���}!��w�=
��X5��Kƭ��"���
���O�7-Vp�)�醬
�7�l�T�W �#�օ��gV�K�ɪ5*p�P9�f�t��~��y��'(�!��qS���$O���5��?Z��'�b�'��I�M�Pc�'����O��Đ%Ě�4��4��M:�I!�����LЦ5*�4>b�'�e�dV|f1�!ճ.���O�""�W&$+�H��+�锦�?9���O\\����vfZ�k��!��ڥ��O����O��D�O0�}J�HC�����F>�,	!@W�a4T��a��V.%#��M3��w�2ˏ�4����`n�[8��'0�6M�Ҧ���4i�`qݴ�y2�'���e���?Y2�NF�XX��٬ ��]��T��'��i>��	��	��h���;4TP��جp���� M��0�B�'��7-_�i����O�D6�9Ov����B��@q��I�Ti�7�Zm}R�e�:�m����ŞM��a�T-��Ck)����.$l>�y�읐c�]�'L،@#����d�`�|_�Hhbd͋
���J�n�.��@Z��ß��⟐����SMy2a�ě���O��#s�>�*uȋ�^纵)��O�oF��4����M���iN�7�G�p_|�9���l9 
VT�XQ@m���z(�!�� I~��;Ma*��I�B��́�ꁘ$��ϓ�?����?���?����O�4ur/�ܰ�h�5VA�$�F�'���'κ7-�0P����M{N>q.ɩ%�<Qe$��"~8Z�j�V��'�F6m����4�o�k~�*\�SWNT�W��!Qx����9TH���������|�T�d��ϟ���՟P���� 3qQ���
�"U�O���p��]y"�yӦ,	S�O��d�O��'A$�� U	�����Y��O:aP�5�'�V�AR�&�d�LQ&��^�d�A�ϛb��bl]6E���%KO�j>ҥ�d���4��� �9b��O�H� �M�nvޥ��K$q�8�f��O����O�$�O1�"ʓ$�F�,<ժ1�eh���4c��^�7\4��'�R iӒ⟬�O8�Dѭu���7'
�S$�\�����e��d�OD+gfc���Ӻ+5��;�Ҡ��<�  hd�]-,Ъu���ݎL���6O�˓�?)��?1���?!���	 \���fd�&]�B|��5S��n�(X����ɟT�Im�ɟ؀���S��">.��	�Þ/(ߎ@@����?�����S�'�D��4�y�	8�8�JD�ֺRq�Ջb�B��y2���DRj��ɿ(��'P���H��08��A�vm�4�h����[�p&u�	ן4��ٟ��'�7-N	q5��D�O��$�1[��%{�N�f&	Rm�IUz�t��OT�D�O"�O܁U���n߂�Bq�4�1қ��%+_
�{��i�^b����x�Ԯ{)8�8䪞��T��t/
ş��I������D���'���K#��m�	�@�(��4���'�7- @C���M+��w�B%r���&���S�
�:V2tҝ'���'���T/f��������HD��iM;
,p##��tD��@��g�ԒO���|���?9��?1��S��8��H�L�h&�>^��-O��m��8����?Y��A&7���ǣ^#0("�0w�W?(�R��?A����|����?�e�ψ`[f�G�u����G�}����ܴ��$X4��k�'u�'��I;*J�H��r�����'$�t��	ޟ����4�i>��'�6��$z�����C]�<[p
�	KJbe9"�&�<���9%�T�	���$�O���Of��qmI/3պ��M�~#�W�X��`��i0�ɼjYb����Ol�U$?����<����ƀM����Z���<�0��ٟ�I����I�8��O�'|cqrȖ�7GұZ�o]��������?�%ϛ�C�?��I �McJ>II�*�$�S��;�؃r��䓛?���|��LS��M+�O�Ar���:���c�(��P�n�	6��'W��<��s��O���|����?���� F�$��d��C�l�8����?�*O<Un�:\����ԟD�	t������0 �B��qtXᢣK5���XJ}��'@�|�OZ҄ܡK���pA�T:pW@�҉U	-�ͺ���)
H�+�O��H>�?IW�*�DH�`,\h�N��f�nE�$�Nj����O��$�O���ɰ<)p�ivB� �N=S�D��&n�;��s��T�0\�	 �M���n�>�B�iY�U�V�����BC��+� a���Um�,�^�mr~R��*�����|�)K,\�f�ZN�y]XcB$�#���<I��?���?���?1/�$����:+��T!t"�rAJ��g��֦��T��ڟ��I�D$?��ɒ�Mϻg�jP��zM0a`t���V&�y���?�O>�|��&���M�'�����]��t��j_�x�����'�؅9�j�ΟL�G�|�Z���qT�+l�,!�t�V��]�5M�����d��wyB�}Ӿ�#�H�O����O��p��B�1�찻`S%;��	�v�:�I�����Ol�2�d�7d�(�q��Hu����J��B�I1��Ѐ��!��c>����'�ډ���R���;L�����0-�I����	���IE�O\b��%��م��j+n�*ĵ;���~Ӱ��S-�<AҹiY�O��\�s�D�Ԭ@�i]��is+�Kl�d�Ԧ���4&u��
U"�f�� ��ֵ���aN
/+F�xq�֗\�t�g	��~A��$�|���D�'B�'�"�'�zP�W�H7x�Hh���b��$�2Y��ٴ5�����?A���'�?����u��uР��T�J)��Y���ޟL��J�)�.%
&���o�^`���E+S�JE"@�%[�<ȕ'�L�*H����|R\�L{�S�Gm2p�B�q��B6ƌ��D�I������AyR�z��9s&�O��@&��aW���U�?ZL��?O�Mm�A�X�	��Mc�iv~6���w��k�
����*�7\�ta`��d�*�^��������>i��/qy����@�@�e4Yg��Iڟx��ٟp�I����IR�'C���B@a�*ج�Jp��XD�͓�?	�#1�V��"������9%��8��E�s���>֌�x�$�J����i>���BZ�i�'"�$(r�` <is�O��i!�ԅU�|������4�R���O��� ?R�������4�u�N P/��d�O�ʓ7���y��'l�W>�h'oJDH�d�5(Fj�Q�8?��Y����ߟ\&��D�v���f؜:��y1nΦb�\�R��Z�줙ش��4�*��'��'[�i�V͂�'����׍�rp�!j��'��'���O��	��M����Y��Q�� ?+Kۘ[D�]h�����I'�M{�2g�>��}�<93�x�֤�6I� VX���?iU	�	�M;�O���r���	� ��d�6|E|l�BѨ@Z\ظv�H���<y���?y��?!���?Y(���E�f,����2-32XIQk����ԯ����	ş`'?��ɽ�M�;wNT���hAB�0�K�	�wL6�r���?1L>�|ꂏP��M�'�q�1���^O�p ���	
�'�`��Ɵ�P��|�U����͟�c"	��>I;�E�/W�����R���8��Ryb�a���G�O���Op(�#ґq�ޕ�a��SI��8F�'�	��$VѦ=;۴{��'3��Ǡ�9K岄�˙� `(|0�O�eI'�-5?P�0f/��G��?�0F�OB�I��Rj@Ka�b�V��f��O���Oj���Oޢ}�� \�0�I M���3���� �p���-���ʆ�s""�'�V6m*�iީ��fT��>��iG�� 9q��f�Ĩٴ��v�aӈj0xӌ���6q��f4� ���I�75Ll����0֮��C�3�$�<���?����?y��?�a��U^��;��CD[d4[W�����Ϧ��������'?�	���x+Q��Hc���U g�
8��O`��O�O1� �JE��:�a��(	�U��l�u��}"��s����`���R��t��^y�n�=4()T�ng�X�G7{���'���'f�O���M3�ݽ�?����7���s�hT)ec��e��?a��iO�O� �'��'x"L��80g �wl��g`T�	:�Xa�i�ɁQ)&t��Oq����S�0�D���Ƶe����d�O���O^���O ��!���V�h�g�Hp������MD��	ڟ�����M[�ƈv~bis��O,@c�

6k`�x˷������7�#���O��4���z��c�\�
Д��6g�3QP�3���$WriB��%~r���i�~y�O-�'����6e�H���kǞS�x��ճqA��'��I��MK�$�r~B�'�S�MG�Ł�e��o4���nv���	�����^�)Z@��͆P�VE�1�h  �C�!���s���M�O�)��~��|ү߭M�ʰA��+ ʌ���67��'�2�'M��P��Z޴e�P8��W����@��0�r���&������ߦ��?�@W�\K۴z�@�S�GD#}��`���G��%���iH�6�G:M �6�'?a�G]#r��)����d��dz�̄e����0�ڇ,��<q��?q��?����?Q/��Y:F�^�^�Es�K1ux|`P�覑��+p�h��͟P'?�	��M�;Q��%;���,\�ZdNl����?	H>�|�U^�MK�'�"���;�fI��ǩp�67Or��a�,�~�|�Z����<)2��$���W"�#�������������	Uy��o�6Q8�;O��D�O���i�'7$�c�i��;�(��$�.�����d�Od�3�d<WsZ��t�E�u$.�+�M֭5�����H��d����|��	����I�-��(2�&^"(n�)sKO�B��x����I֟8�	V�Oc�惈#8eP�dS�`/<ģ����)`�Fu�&����<D�id�O�nόhYL�&Q��0DY$��$H��O����O���&a�x�	ʟD��K֝yM��-K)t�D����

d\z�C®1Ud�&�L���t�'��'���'\TU��G�N��@��%F�3=�aV�؛ڴBH̘����?����'�?ї�!GP��Ո�0�*̒v�M/
��	�� ��v�)�*G$$�`֧�7	�У�"]�c�,Ufw �E�H,J�D�O�@�N>a/O�Щ`�ϥB9��'�	�ZղQ��C�O��$�O����O�	�<�!�iv�����'3R��!��)�:Uk�iW?R;T��'p
6�0��'��$�OP6�ʦi���,w���G39|:*���?R�o�f~�*D����Xܧ���G,$����&C�K����l�<I���?����?���?����V*b�l��"2$�Z�X�%U���',rjc�\*�J�<q��i��'/j\�dP-9�QR�̭,��H��&��ئ%a��|�l�M{�OV�X5�Po���#B�+B�5����1f82����20 �O6��|����?1�J̔2Ԅ�1�:趨��.�R����?�)O4n�HWH}��̟@��V���  ƚ,Z'��z
 Zp�Л�y��'���?�����S�t/�*DbQs�ޡ5|����!��Sa 81��5��W��S� �r�M�	� ��H'� q���3��^�9l���ߟ����P�)�wy2�f�)f�wZLQ&̚9j;Tl(5�_{�8���D�y}��'�|\��J�m0iA+���� ���'�Û��T��f��L�Ԗ~��7&%�8�f���+� �p�$��<I*O����O~�$�O<���O
�'(��k��K�)E�t���:iT��p�ie�t��'3��'Q��y��k��.O��`D��PA3-�8���lZ;�M3Ґx���!�}W�67O��*�É7aā��Tc���78O0���_��?�F�<���<ͧ�?�#�.�n�0B��<_(H�PC��?y��?)���������@^�d�����f�9c��
�j�O�����%�Y��)��	џ�	C�I����c�h��J�R2�F��P��
���A�,~+�(JI~Ra��O�(�v��\0���#6B��סT�Jz�����?���?a��h�����!Q^���3�T����i���-$ab��Aʤ�QUy"�q�.��]( ���������+]=aq��ßL�	��걩����ug.]8`v���)-~h�6�غ��`r�lG��$�x�'3��'���'�'
�[cH�v��m����(�~�Z�S�$��4bͬ@��?y����<I�b�{:Ҙ�#�M6�lУ/ُs!�I����I\�)��4��@$��2	1�9��F�E.B4�VN�զM�'`!	���x?QN>q/Oj���5	ǐ����8��r��O2���O��d�O�I�<�e�i�f�1�'h�K�OٸR��馡�5��s&�'�7�*�I<��D�O��4�d\X��҂b���4n�"Jl|����,:�7�0?�1N3�i���䧛��P�2�����̉1���bO��<)��?a��?����?y���ɑ�r�� ���b��Ň���'�r�k���:�`�<�c�i%�'3葲!l��W�p]s�&���x��w�>���Ц����|�$��M[�On��`� �X9A�A6Mt�kaBG0x����u	̕�?qD(���<ͧ�?���?�e���!@.L�(��1+W��?!����O�]��&�ɟ��	�ДO�N�2�τ9Jd���Q�J��$?�[�\��4����$�?*�M���S7�׭a�J�ӕ��r��t�4'u���|ti�O&`�M>F���L3���	[ѐ��?�?����?)��?�|r,O�lڤHCVH9�Ɂ�.��ؼQ��@�F�UyrLm��㟤�O�(l�F�V�)��A�=�����C�nqy�42D��������!��<��D�Cy�o^ ENI�嫝(M��X7 ���ybT�0�	͟H�IܟH��ޟ��OH��cb_(�((�gb1B�da� g��A�"�OF���O���@��NΦ��k.��k�#�+m��� � ( �0��4#��j;��	ۖ@Y@6Mp�DQ'�]g]���Sm��R�� g�f��qV)��?�rE[]�IZyB�'i2������&�T�9�,�!���9`�b�'�b�'��I8�Ms���?9��?Y�c�4���=�N5�Wi)��'<� 6��+w��0&��r)ߦ:��$p��
V��qM ?i�(��i�XqC�9��d���ڹ�?���;x�	"���	cp����?����?Q���?���I�O���4�� %2��U �0|��Ͱ���Oh�l��]�(�I�����4���yg#F<��-b���w�V�#d����y��'���'���jB�i��ɯ��h��O�X��.�!k�8%+gOZ�)�ڐ�2�Y�IHy�O���'6r�'p�ckq"ebU�_,t���p�=�MS��E,�?����?�M~�����%iZ�$� ��w�ODW��^�$�	ޟ &�b>�[!j	�q-ȭ�T@E:)&���J�U�@=w" ?y5�V����E ����H�X �����fj�G�Q����O����O��4��˓q��fϐ$L@��_x�hC���w���`���y�im� ���O���O��d�/ �����]d�6-���X	�a*�-h�P�7�%x���j4;M~�����A̚ Wl�Q+�+���|���?����?A���?9���O]��G��Op�j܂l��3��'~2�'}�7�c���O��n�]�	�]�܌I҈�3S<�|��m�9���'�������:�<le~Zw�����M,H�-ɖ%4$h�G>��H�@��Hy2�'��'="G��a6���Z!fܹ�f�e!��',�	��M�4h�0�?y��?I+�H��̞�6�. >!#r��22O���@y�'����+�T>m� �@�����S�1`t�A�7���g����������ߟ�ڃ�|�
�`F��ѭ� b&��Q9s���'�B�'v���V��3�4k@ʕ@�͌�+,!�$A��a�!sf�	��OƦ%�?m�>qp�i���D�<=�(�1�ۉV��U���pӚ�mX�VPmR~�d�=	���L��ѢX"�W���jRc�[���D�<����?����?����?)/���x�G�4�,��*��)#��*1�Ŧ)h��䟴��ҟ '?��	*�M�;	%8�J@��*rӊ����jtd1�E�i�J7͜t�)�Ә>TumZ�<��ĝ�u�PQ+����Q"��<yG�X��p������d�O����p�6@�TlX�ZPXsWLЮ,��D�O��$�O|˓6&�v��-��'��P�8ޖ8���G�Q!�%
����1�OD�'��6-Ϧ�(N<�aǋ�;���2�Ć�r�Z�b�m�{~"��?�8@UD��z�O�>4�ɘ32�̹�Hq)6"�J0~�;v�O�|R"�'��'����ٟ��*�L
�Z	9�nm�0LA���0ش	�r��?1��i%�O��0��Q;hr������9����O�7-�Φi��������'evHxf���?�P/��eհШ�e�2��u�!t��'�I�	ߟ���ٟ4�	2){�jF��C�-b�!�>	[���'�b7�U<x��D�O�D?�)�O��B��R-��q3n�T��Em}��'s��|���B�*t��0�I�YU�D�	I�C��\��oُa���&$���'5�m&�Ж'RdH�u�.c��#C57޺���'Mr�'������Q�t3�4��@���k9�����s`�iR-M��)��QW��|B�'}�ꓻ?���?�p��*qP �Q�Zz�1�gM-�Vb�4����y �'�䒟,��3Ae��IX�6��'�1n��O����O����O���2���D��4PV���G��UP0N�D]`h��ß��	�M�%�M�|2��6��&�|�D�5s�����	�=ޔ�S�
L�'����$!7E�晟�]#sZLu3���J�r�p3���t��Ǆ���ث��|�T� ����ԟ�z2,^��z|H�M8[C��CDk��� ��Ry��w��P���O����O�˧�:��i%w��,� ��s8`ϓ�?��_������$%��'�RL!Ӌ�9^,1�1!'9��R�mΔ N t�ӁS��4��0��Kiv�O�|K�@�U_Z�S���1�x�%��O����O���O1�������z�Yj���+Ui��ťRP�P�W�$ܴ��''��M3����zlF� r/M�\V��h2�V!c��m�2����fӼ�zm>��b/쟌�O �8Ѓ��l����Jӝ]�F���';��P�	ӟ�������`��[��^m���6A��{�,�D��7� �,<�D�O���<�9OH�oz�aP
�&N�<���(w%�6���?�����ŞTQޱ��4�y
� ���C@̄B<&�H�e��5n8
�6O�L����~b�|S������S�ЇVhS��<�x�Gb�ԟ �I����@y�`sӲy��3O
�d�O��!u�F(1Y(9! CT�a��}aB�*�	����O(�$5�D͊�>9Z�GO C"2�
B(���I�@�D�)w(ܦ��|JB.�����eaJ�'�z��L�ā�|����ןd�	�$�IU�Oh�ʐo�-(b�4*��q#�W�/��{Ӏ��V��i�4���yw��~dځ�˔���`���Ǆ�yB�'0��'�Q�i�	�(��4�Qџ]�,e�R�� /Qb#�� !�O��|r��?����?a�!tf1z���1t2i�E�Ax�S(OHmZ�B���i56M�Oޒ�����9נO�`GF���B<N�U�'�2�'ɧ�OrL��M�vt�dD���:��]>e�P6T����̆vj�!�B�IFy"�>V��i��O�Lu��ȃ9�r�'��'��Oh�+�M[�ɇ�?�aF@�t�����܎z�]��͐�?Q�i��O��'���'8��؈h\<)�@�C���ˤW�*�Hl�¿i��	
\w�� F�OEJ%?���)cIZ�s��M�X��T����������柀�I����`��!2dCt!",�\��M�]�D�x)O������Y2If>)����M�M>� �k��r#L#2r1��N����?���|�C���MC�O뮘�]\���Wc��O�ڵP@��8r���j�%�O�)�N>y-O����OT�D�O ��ԥ�0N�2��ѡ��zo��S���O`�d�<�Q�i����B�'W��'r�S�K�l�!WH�7X(hd���� a.���������_�)���C��$� h?t�"�*���9Y�����F��d -O�Ɍ��?�!=�D�0Z��gY������O�4m8���O����O"���<�G�i6��5�M����RlǓ4LȲ�Y�QA��	�M��l�>q��i6�	�(�8���m�{�@Q��Hc�!lZ%V=�-m�D~��:��v�)�k�|�C�Å �b�.X��~�[�<����������IğL�O3b�Y����E��(E��)jE��E�`�fԘ�#�ON��Oj��^�D�ڦ�1�&u;ae��B�xl��h��e���۴.&���0��iZ��67-s�� �#U��/9ܠ����FO�d�*������R-��O���?��Y�� �6ɛ�A�p%ې�_FP���?����?a/O�nZ
�����������X*��s��Xܨ�|�IП��Opm���Mr�x��FJ�%��"�`�r �����/$E<B �X�B�Γ�40
�@�\�$�62⬈�i]:,�\Sm]�|�����O��d�O���4�'�?9VI��UEj�hH�7�����O��?A7�id����'Q��s����ݷud0(9�� s70���=rъ�ʟ����`��Ǧ��u��8s���'V!�*�d��4����%��yk�U'��'���'�B�'��'Έ���� ��V�ŞxqzJF_���ݴF�������?����<Q��U��9b�dW��sk�'��I�Pm�2��S��t����%�G}~��d`]�5�+�X}d��O����۱�?��-�D�<	��U ��$�rBZ�%��}���׌�?q��?����?ͧ��ć���H���H�vfP!��,�g��|��8����K�4��'���?q���?Q�-�&/���4���g����� �Y�ݴ���;>Jy����O��&��O�*�Ը>
����=�y�'��'���'���)ԱO��x r�ܯ{�L\�ba��5�D�$�O��L��9��Phy��v�O��!
�3'�J0�j�D��D�*�d�O&�4�~-R�wӜ�,n`�j� Ƙy��L��*�}�#�%� j���4����4�����O����"�����q
�xa %[�;�j���O��O��aY����'uR�?���.'G�ݓ�ƼJC�pI�X�O����OԓO��(����#�,5c��gc�ɞ��"ɧn�ȱP�fiy�O����ɘq��'��h�$�](ۚthD�C}��R�'fr�'8��O}�/�M�����m��YU�Y�czA�� ����]y)OJ�m�\��ez�I��M+����9��!�$�	9�LY!�D���v�w��-BԠ}�f�9�� Y4�d�OA�,�$�_8Ш�`�5�D�''��ş�	��h�Iߟ���n�$Av������ ��z����|6����d�OF�d?�9O��mz��ٓ�	3׈����Z>/�5s!+���M#G�ijnO1�R�6�m���	�w�]�s��Z�n5�&KJ����>�*��5�'���%������'�Hw��%�<u������C�'���';�^����4m>Dϓ�?��(]X-������S7O:�tL���i�>����?	O>��J�g-RA+��Э
�4)��`~b˸[�F��@�if1��
�'��M�.���ZC
�l�@�B�^��'*�'���S��ٗ��j���!t�A�o�5�R'�ӟ�ߴCwj5�'��7�%�iޡZ�c�;)�fe�s �<�XP���v���I�\�I�P� )l�W~B)O/wnt�'	�8q��(��p�U�D�L�wCZ��H>�,O�)�O���O��d�Ov<1ťI�p�ܸ���͆m��f)�<I��i��e[�'B�'k��y���9C�DXrR��?�i2�T�,듊?1����S�'	@�� �asÕ/MÆD���ԋ+���EeӤ�R/b���ϼ��&�ė'�R5 ,�&@�~�"��s-$��B�'���'D����]��޴,VT���޵���8kx��X:�q̓P��6��j}�Om� �l���M�a�;{��H�%>�؅����-R���ڴ��d�x�T\���˸O2��^H�]"��,"�$��'ה�y��'���'W2�'`��)�����4@ tB2f�24"^��'<��'&�6M�����M#I>9Ug��N^x�뵠Q��͓d����?���|r@�I/�Mc�OH�i�ۇ��s�F�;��� �-�-d�yH�'1�'��i>)�����ɴ������ �z
�]�jٔ�f!����'�7�=\Bl�d�O����|:����!�=���19f��)a#b~Ba�>)���?yI>�O4�hsp#�"�DH���϶?�>��c� ��AD�Z1�i>=kp�'j�%����
��΀x�CU6~F���h��@�	۟$�	��b>I�'��6퐵q���T���~��L#��XqF-�G�O<������?2]���61pm���Z�Xp�hA�R����I֟� �GF즹�uw�~]�thAvy�ё]��k��8c@�m�f���y�U��I۟��	ş�����O8�
) xy2A�0�ˀ����BEe�JuK��O ���O,�����ݨO�\i�feI��1��.�,�R����l$�b>������1͓$�t1bRo��+�r��U$F���i�'��)b��Ovt`K>*O����O��!Q��;o��]�&������k2+�O��O���<i��i,Hh��'x�'YB%���zc�d�H�Cm��B��d�Q}��'ҕ|��xg�\�#V6"���"�V���dG�l���6as�tb>����O�����$S.�#��.;��p�S�I*4���O����OD��0�'�?�v`^0*mL""�
C�<�����	�?���ipb�I�Oj0l�D�ӼSv�m0��1A�o;��t+�<����?��<�} ۴����Ct@�:�O
И����-e��T�U�a�Ba��|2Y��S������8��ҟ\�g@�Cڡ�5dѷLE�Ty�(�|y�q�֩9�4O����OR���9���DY�&R��e�?KΤ��'
��'cɧ�O�r����L9bLĈ�� �	���y�+ՁV2�������E&T��)�D�<)�ʗ�2 Vͫ@m�T�(89��(�?��?���?ͧ��$��� `T���Y�+3Ј���lށW���P3mQߟ<i�4��'���s���lm���m��b�!�f������
��z*���Ae�I�'���Ä��?����t�w�8��#Q�W �kT�G�}	1�'?B�'`b�'WB�':�n\��+� ;'�50uǌz#Z]�Ǫ�O�$�O@PmZ��Zݔ';6-$�<j�\P��}�4��ůL8[�(�'��ݴB���O�Lت�i�	xh0�hd��1p���	��=|X*� #��F��ώ^�	Hy�O���'`�E�$m��iv"M�e�@-��ꂴIH��'0�I��M��F��?����?q-���1�\�8�PɁ�J�>D������ɫO$���OȓO��/WfN�!/X-rZ�i��O>b
�r��D�Rhm W Iy�O�N%��dm�'������A-;,��j5[�ˌ)Q��'=��'����O�I3�M#v.������Y#s�v�r��D;0�����?)�i��O֩�'�)�~&��Cs�0EѺ$����1B�'��`��iT�iݹB3D�?�ET�0jE,޿�.�Sì�?@	Ra{��'�B�'���'���'��<W��u���^-2�,P��E�p��ܴ|��ً��?������?���y7�ٶ�H��N���d@�K#�7͛��aN<�|�r��1�M��' ^��j�Wm�]�4N�Lَ`�'���r�z�7-S&�䓹�$�O�D�
z�v��#�ܣ)�mC���v����O����ONʓ-țf�����������5C�P�A��ߢ@"V��&��\�F����M;��i� O��x� R�v�(#a���΄����J��v�LYw$F�w�"$Uԟt ��T�81m��F
-�r防�2D�@��?\��{��K�<�X��Q�P���rܴ3��yi���?�i��O�.����S�qϴ\х��T�l�(6O~�D�O�� X6�,?�;y�D���A�p=x �F�)��j��݂�Нõ#>��<���d]z�h���D�d����RA!����M�*�?I���?y��F�:N���ѥۋ���@pd��B��?�����ŞQ�|tJs"L�1�R�
W͊�m�N���Ƀ+m'� X)O���/I��?	@,�D�<a�H�����BA�&�8���j�(�ݴ-7L�B��� ks�\0`�j��Q9r�h((�G�&��E}��wӈnځ�M��hO'r�V}�Ū�_<$�+ ��?�~��4��$T 5��'W����.�.��`<a�ȗ�C=�|Y�N@�q��$&�O`HSF�݄y ��֋1ߊl餄�Oj���O�elZ?a���'�6�|"�8��Q�qe���>L9�G;"��O�tlZ��M�'f��4���V3Xp��
!�>/j��@⎷�܁ FdJ.�?���/��<���?a��?�Љ4a�vх^����v���?Y���$R�� w*ʟ��I�D�O͒��4/�Y�����L=r �X��O�`�'���'�ɧ�� B�gœNN��Fd�L�B�[� ��{p,@Y��Zl��i>u���'�B	%��pw�Y�7�AZ$i�"p,��1�*�ޟ,�������ןb>1�'z�7�T�'�5ڇ�c? ��l��δ���<��i��O8��'��A/)��B���V$51�mm���'�d@��i��	#B�+�OG�5���O�$����*��"�ƨ͓����O��O|�D�Oj�Ĭ|j0�Hk|�ҫٍ<l�w�%��f�M!P��'����'87=�\I0�Zwx~� �"�|��q���O���6��i_��v7�u��Ŭ�?���`%P���)��k��x�@�A	+N\�yy�O��jG���dKC�ؖ��s��&��'�2�'��ɥ�MK�A��?���?9Q�̋=�l��J#H��<�������'����?����#>,�rnp�b"�I'\t�'���1�h��:������)�ڟ��g�'�$$��U'o&��#��u����'(�'���'��>����.��e�WI	Ie�����A6��	��M�����?�� V���4� �A��"�dC"	0Sܴ��>O��D�O����?J�h7M??�;S�����4��x͜+7�ʈ[b*��aI����-5�d�<A���?y��?����?a!�$M�b�GǗ�*��g&�+ON	mZ��:-�	ٟ\�Ix�ٟ@�xq(4P�˴h�@��t�������O&�&��Ɉ52Yv�	��z���$��7��@�U��ʓ�jHhW��OB5jI>y/O��'I?�L�(L!(��b�O8���O����O�ɪ<�1�i̢=`�'�4Z���G��(`�"_2ī�'��7�4��	����O���O�Q����+%��ӑ���f&���%����6-.?ٖ�� mV>�	���'���B ���ϟ�3��E��g��������	����I�T�ZuV��vp��^�Rj�q�#����d�O�qmZ�dϚ��ğ`��4��n����r��|��D×)�2J���N>���?ͧ�J� �4����N��1�
͈Um�:J͔��A�� ��YY��G�\}:�k��(J�	�.��+p�]�tKעe�.�+㇇�>׊�	�hϸgS&A;���&��P��X��.<�u��-찉�AQC�U��M�,@�qb���5Vr�I�\�������T��K�'.�����[�\��h�1O	��,L��HËo��i�̌� 
!J�/?�\l��[�H��l0���s�!�G�X�~�����+�u6A�$'�EH`uK�M�JԪ��'��Gn��ąS�R�� .�aV��V�wf��eR�-x�+GΊ
G��!h��ؤeP�QQ��M���y��x��$�O��� Ӡ�NudX����=�C�R�my��O�S+��)X5�ϤX�NX�0��(�j6M�<�J����~���֞�*�n�<g�>� Ԣ�4䆔	��j���h�Dx���'C�>� � F:&@�9��c��4&�4E�2�i���'���O��O���C�4[}�Ă����L�6$ҌZv\qnZ

Xv"<E���'�>`�R���q�č�'n� ��f���$�O��$ B��$�t�I쟘��`������R�ԡ)�Ƌ�iS���>����[��?���?��T >����o^<��y*�-C�w����'����G.5��O���8�����2��H{P�D���݇7�h<p4Q��0��(��Ɵ����'&Є9 ��j�f/�6B�d�	��b�X��b��EyK E��}�H�;=u���V� Z.�Q3�y��'��'��IVFj�O��L�faS"$gf��bj	��j[w�����vy�X��S�i�~��mB�k����;7�����s}��'���'e�I�y��aO|�.2|�z\���:�ʖeֺaԛ��'��'��I�;.Fb��0u��7\�t��i��<�{b�y��d�O6�}~N}�K|J���PǑ)L��#V��6K�`��7����'��`�P#<�OY����/ˆT�l� ��`��ڴ��D�g�oZ:��I�Ot��Sp~�k\7X,킡�ܬ :����)Κ�M�(O����)���(�`Ya��"?�"���O|�7m60-�mZ�(��ߟ�ӏ�ē�?�@���󑋀c��,IUCҼT�a��'
P�f�	5E�L(�FSc/���t&jӞ�$�O���
m�^I%����͟<�D���BN
�RD>(jӡ�Y:�H��	ҟ��	՟�ہeR�k���㈍��������$�)emh����OH�O]S�J�eVn6��v��&O7�ēX���'���'�R�'�"�����2F�ޘ!���=)`9�Q���'HҐ|��'I��I;a���Y�̞�kI�Y��N����M/��D�O����OT���O*p�Ao�?Q���̂r�D����	a8��o~Ӱ��?�H>�������5g�6'�"?4T�ѳF�'6$l {Sh������O���O�d�O�z1��O��D��TI%�E�CuM�"m�{�Ґ�t�l�f��,���Od˓��%$�P�c$xO|�q� �����n�����O�ʓe1���6X?I�	��l��@3�yG�h����Q-�$`à�ZK<y��?���2��'����2�D�G
�>f>�B��Y�vR����@W�����ȟ��	�?���5f%�*z���+Z:َT�3�ŕ�M���?������O�,���EͿ!�r8����!H�U�ٴ#���i1��'�r�O�ꓞ����V��C㗎.�V���	�1\qlڣ�H��?A����'m�� �3b"S�LPD�Ñ���|`US��iS��'9�ʋ(j"�����O�Ƀ?��ǯG.=~4���͚)|c��"Rj�K�ӟ��	ڟȳ���b������ Xup��B+���M���Z�X6[���'���|ZcR�0����ԛD�<9?�a�UY�t���QV�	��ş̕'\����F�I<�L ����Y�P���Jҍ�듖��O�O����O@hل�u�s�_�sh�I�@Úy>���'5���OD��O��X�E�C:�p��Vo(f	�WgƐ@�P�i��ޟ�&�D��ޟ��$�X?��
+�|�y�(�1&�$(��TY}��'���'�剻����F�$
�BXÀ�c��������Im�\'��I�l1��Wܓ-��E A�<.� !Պ�6W�lIlZ���IRyb�JP$ꧦ?i����)l*��V�#���qRM�

������ӟ��.EU��O,�SJ#�ӆb	�j\N`��<_��6M�<�F��\����'&��'����>�1@ ��S�ҡ2������5dzqmZ��T�I�n����?Q���`ې��C�$��`��׫�M5F]�By���'��'���D�>�(O�`W*�?cz�I���n�TLz�`�ߦ�7.����%����� ���sg���R�Xy�1��`z��i��'�����LG����$�O��I�^�����
7�b�����=B�6M$��",��%>��	����ɗ 
byz�&݄4*�T����k���޴�?�G��d�O>�D�O,�Ok�^~*}��	R��\h�ˉ
3���O�8�&���	ϟ��	Cy�N�ފ��Uk�)��I�gos�!
eQ�ޟ��IM��^yr�ڿs+����	ȫ�~M�`D�?A��ث��'M�	џ��I��0�'�� l>Ir��1aѸ�mT}�d����>���?�M>+O8P�6G�O�i�%_Gڈ	�"����X��3Dz}b�'B�'!�	%o���L|�ׅ�I���s�ԛ[���P�߮ t�6�'u�'@�	��d��L�I�?1�i��
ζ �6��E�C̛��'��������X���'���5���&d��T�a疭�rT[���ē�?��{�#s��a�S���V�_���w�N�|-H+��߹��D�Oz��P��O����O���:�Ӻ��I��	�@����d"x�:�@�ŦM�Iޟ�@ΰ%��c�b?���j�h`P��Ɛ!�6=p�"`��ޒj���'��2O��Z��nwp5JF��p&��1���,k�`�'����Nw�S�O��<��B70ź�*����yP��}��D�Oz�	��2�S���>񗀛�rš��O�_�1h�ȣ �1O*���\�ߟp�	�t��EBv�I��Ծ^��K�d��M��:������x�O5�'��I�E �-)7㍚I�9" hӋgQ9K�4�?y�W0�?(O�)�O�˓�?Yp�˄e���@ O޹]����
��HP.OB�D�O��,�	ڟx`q,�<:x�a$�ʧ\b��h#��5X�t;Tl8?����?������L��|�Χ8��IÄN�`h�S�әQkf��'v�'��'w��5ry�t�ɾ2e"ݸ�O���#�OH�U�f鱬O����O��d�<��&Р��O3��VΖ
��|�0�M�z�
,)#�p�����Odʓ�?)��0�2y�����%n�~=8UB�Ӥ�Ic���:��4�?i���$ �k���&>Q�I�?��f�ja�i]�v4���@�G,�O4�e�R����䧗���B�V�s�L�Pa��C7�M�(O&�A���E"����d���a�'����w���TH�J�&5��4��$��t��T]�{�s����`�0�n@�!H9
���4�i��h�Mp�����O2�D��l&�擾݊����̐M�*+s��;+DF��4b��qy��?y/O����D�Od��S͜%b�xp�aPP;l(x�.�Ϧ��Iϟ��	+��E�I<�'�?��'�(eI��~p��a��y8:]�ٴ�?�)O�@�.�L��'^b�'���:��=����hv��I
�H^6�O|���N�i>��	�ɺtVB��$˫G��� �� aI��O�h�GH�OZ��?����?a)OF{c��hF��4e^9�8ؒ�g�&�t����'�p�'�@1ĦF�5yNĠc�ת<328K�/B)P@"U�$���D��Ty��O�u$�i��9E��YB�S����6m�<���D�OJ�D�O�M�0OT��d�U�	$xHc�#�3q<vı���{}��'8��'��I#�~j��L��U5����/C�sT���KS��o��(�'Y"�'��bI�yU�t�d��8�f��T �5PcXI#`Q#�M+���?�.Oy��ˁ\���'�B�O��ᢁR�q��*�ߙe��vh�>����?��N�ƌ̓�?�(O�S�^x��c��X/q(t����&>r�6-�<iU`ݶC�vD�~���������O�F>��(�J/X!2�I�l�����O80��O��OP�>�/w�.0Ӥ�_ 8�)��m�}D�ƯǔfD27��O����O8���f������ŵ6��ڴ˘��L�x��4fNz�
�b���Oҵ�G�7c�.mˆK\'����˦��埌�	qڀh�}�'1���|���`3)ڪzy��fB3+H���|�ED��yʟ`�D�O�S��Y9�e�7�0T{���M�B7��Ox1�T@�F��?YH>�1r0 a�2�ze85 2.E�:��'f�)�'��I�������'N� �a�A�	JI>��r�Z.W$ta%�Q`�'���'��'���'x��j%��s�JuB5���EH��i���"�yB^�4�	ǟ��Iyy�IV�L�:[����!�3��)���\��>��?A��䓎?I��|�"��Tǎ��5��/Vm��MS�Q�`q!�Z�(������Iyy��;M\��~�`W�!>Hy!�Ҷ_1T������e��C�	ɟ`�I�N7Y�IK��O�HzBę���@%L�`a$����6�'�X�𪁃J��ħ�?���@zr�[R��{{���@�w6��x��'�҄�	�yb�|R[?�@�b��5	ƀ�QJK/`4i�D�i)��,xA �4m���۟L�����I:�Q:sOf��e��/�-��6�'f���|��I�~4��ǅH�X�����e�����6M�O8���O6�IW����#Pj��K��N�T)�d�B�'�M�E��?H>�����'KB���&��� pѮ�Ґ�īi���d�O�d0w��8%���ܟP��I��(��;Gi<�IFD�)� ��>y������?����?I��ՁI��y"�ݾO��������&�'�6��w�)���X'�֘0`�4�C��F��f\Cb�	.8��U��Y���$�On�d�O��?��!ӆZ%eڡ��̏8+>:�"gˍ2{�O
�d&���O�DO�v�A�&mLh�ĂUuM�ء3O�ʓ�?I���?+O�`���|�fn�r/�a��$�-iz�r�}R�'h|B�'iro� �yri��d6)`b�2J`Q�VB�<Jg�듐?���?1+O��2fF�l��Mk
pƘ�?�������I	E	ߴ�?yL>���?1�M�c� H½�TĀp	ܩA�#�M�UoZ����{yR\�B�=���O:�)޻h���1
L�D� �m[l���$������X������'��i�5��E/0�R�%���D�m�zy�f�@Z�6F[���'��$)?a�fS:j%��;���[��Q��V}��'�0|��'�ɧ�O��hA0#ɢ2�,dJ��+*��
ڴ	�� ���?Y��?������|Ҁ`�%H
!��ɏ�D���p���O5�f���
�y��	�O6 Yv�Ԛg/.A�![>^���+���Ϧ���şt���]�rq�I<�'�?y��vkN���Lض\0Ɋ��O�F#b�����_�1O����O:�$N�) �ۗ(��j�X�'J8���'!�%�pR�8�'@r�|RH�� �����#V��(Z�d��3՞�Rc�E~��'{�'���*��D�eJ�V��`%��?2PqZC�H*���?������?���u�^�Q%���>=Jw�Q�$��X  N̓�?���?�(O�XH�c��|Z��W.(Em`�H7M��e W�GL}��'�Ҟ|��'�b�]���'6R<x�aV�K����@P? E����,�	ԟ�'�T�"�G5�\���x���]�ƨ;	��u���l���%�0���0"�8���9H�p")#Ȯ�x ��B76��O��$�<9��P��O�r�OX��'����(W��+.��Bu�+��O��d��v��P��Kmȝq�쏘/�.���
4�MmZyyr�(lP6m�T���'��Di%?!�I�X�ʰ�DO��zƏ�Ҧ��	ٟ\'�&ԸOv�I� C-Sb<A
��_���a�4Q�<d8R�i���'q"�O�Lc�L�6ɇ�Y��"��O`�(K�M3�n�'�����,q�0�`��t xp���	hE��m���$����|�����ē�?���~N@�8ɂ��ô	��`�R
H���'|`�+�y2�'b2�'hnhV�כ6j�����1?Z�a�f���DO0��'����Ɵd$��� ��u��EˬKx��"5�a"�N#b��<���?���?i��x8t���
�x�Ri�@[;�����(�?����?���?�M>����~j ?D�����Ǔ&����N��Mpǜk~��'��'b�*-��R�O5�}j�df�Q2фK�Y���6����O��$�O����I\?�b-�[��M�U�HDn��Q��w}r�'���'��'���#��'���'c�T��Ջqh�Qv�ãe A��/v�>�/���O<�L���$���Ш�+`t�l�g�L���A��LyR�'3����X>y��ן��S�^	9���F+
�ؖ&H��z1�M<����$�b��֝�KN@���ڧ�튗��@7m�<a�<&��v�~����U���!7$��GqH19�C��T,��S�sӄ��OVp�B��Oܧ;��(�ҬK��>���G~���P���Ll��r�i����?�>i����m��@C�_���)�a�_�<��+�ؼ�KBI I����K�e�
�A@Lȸ*�,�0tmZ���-�.���\�JUÎE�I�q�ZXI���!0��:�k�0����L����L�C�_��^\�@���\��1�̫'"�Qzh�>0�	QN�����"��:L:�q[a-��l���Q`��!Sᡎ��?a���?��M��N�O���o>a3ŋD�&?v����J/����$�'U�񁊅*�f��a�]l8�]��D�5�<Es���rTعe��9.�� ��61�Dqj�g�o���C�뀛p���r@�=^$�РSX��\�L�
�)M�O^�d.���'�i�vgI�uk�	w2��'�����V���H�ZV���y��>�-O�Ј҉�k}���� :�*^�X�><X�ͅ�A�Z����O���¸l�~���O��So��0��/
�Q���G���IqC����c$Y( ��9
�J-O�}%��t�L�
��25+�6��$�j�`fc������hJ�x���?������w���A�̀~ɰ'�W'21O����ubn�����9�����((/!��B���H��= ��t���A��+DGf���'��0:ծ�>�����\s0h�D��5��D��Bl��`� T��$���O ����A,��( lN2�����|-�\���W�L|`H�4چ	[�� �>��X.:}��Ѵ���|��D��Ɇ�?錉{�f��dɰ@�Y�;~�ʒ�����D��'n �����~����䁞
�x!h�'gU��(��$L	��⟣XY���8��t�`�:��I�nã�.Q�6dK&�M+���?���F(�+Q��?A���?)�Ӽ�E�T>4��+��/����h����/KH�SNW���OH;c�*?�.�`!���E[ ��<������i2Qأ�P�q��'�F p4�ն�0,��K�C[��P�'k\7m�Oj�c��Oq������2
�)�vUÌ�r(�j��K���$�{@�;u�l0Ud��$���׮6?!��i�b�|RP>�'0d�k� X�	�v�Q�a�;m�Z�A�V8��5���'+2�'�� h�5��Ο�ΧshА����d5i��mr��ל:w����	=-��ϓP�Q���:u��xF�G�3]�T"e�ԁb�Nb���Q���a�N����KBap &, �N���MҟH�IJ�'*�O��D����Ϟv�\���"O\t+!�պs(���.1,n��s���N}bS�@����(�M��?� l/-b��)�*��q<.)�!�^��?Q��vYV�C���?��O%dTH����/�2����4^ѐd�0�@T;�?O܁�����8���/�5uβ�1C��C�x�����?�J>�Q��H�1�j[�[k��� NNx�<9�U�q�ܸ�e��$X}�u)���y<��i.DH��[�	<Ѻ��>�<h3�y����3�>7��O>��|Z�
9�?�0��&J[B-��\�RĐwH�>�?!��-�l�놫HN����#O�<j*��˧F/x�;Tf˘H�IH&A�S=l�OX��J�ȶ����	B�"}*Eo�
��m3���%C�M `*�g��IjOb���  )���RC�+!NQ�!�G�\>m�P"�:s�`d����ax�$�5IXp`�� #_hJw�-L���p��i���'��M�&"|��`�'L��'�w%A�ՠG,DD,����`���rF��B�V��y�m��]��2��t448%�I�׸']�,3	ϓd��qJ���C��У6���(�yB����?�}&�|��   {��
]��a�#�.D�� g��#F���� �y�g,?�u�)�')�k�IQD@���ܒt���`1
��@V٘���?Y��?I��0�d�O���� �����}ufL�bʇ�)���P�!��^�
�pyK$��DԖ�1#��C(�*1O~iKT�'D,� ���0.�f�H3�2���'� ����>9M���#,6'�p
�'�h̫���RJ��"��ɝE��Ū�yBG6�	�O�����4�?Q��G>�Ŝ�[��� �mZ:k��?�����?������!���?�N>A1bR&2xظ�����Ҙ�SgPn8�T��e>�	i�.��)���<c��j�&��ܧ@�|�B\�^����nҰ8מ�X�`���yb�G��:���R:^N�$�g!H2�x�/x���b��`F8�h����`mZ�����t��'�I rc�&q~0�b��>LW��`  (G=��'��P�7�'1O�3?�%�-42�M�f�	Ą�Z��R'	���?����=,��Yj���:g�8({�o-}�,���?��y����ǭ~�
Ə�	3����э
�yr �3z�r�2�A�-���{�I�0<9a�I+@�*�B)FH�j7�W�6��Ź޴�?���?y�ώ����q��?q���?�;i����`Ϯ�y�(�L�x���y�̊��<��-�v�^Iq! �.�^�a���Jܓ[@&���	+�8mR�ሞ�����߿�R��<�A�����>�O����nM�pV� ���;;���a"O�`�䠞�hT�D;��Q��di���r���ӆ:2l�(�␋#b*��Z'2��T��h�)�
��I��p�Iџ� ]w$��'��	ι�� ��YR!ǫq^|�a��^�m��y�f�&�� ���%tP�x�%t�{�`V���C�ɸ't>y�wI� ��y)G!Z�'��4�#b�On���[/|����P"�p�O�9!���&�� ��/ʯ5�u�I�D$1O���>!5�� =���'b��5D �C�tX�jaG
6 �B�'�@�S��'|B?���ʀ�'	�'��(��ņ/����I�y��D��4tf@�?����c��@�G�.��1r@�T8���W��O��Oy�``B:Cx�0�'V6v�9r%"O���"`�;8Z��",�� pv��O,n�<�&-����1�`q�3�G	 s.b�l�vm@��M��?a/�:|�W!�On](CN�s�d��	N.Е��B�O ��
�yZ�$=�|�'.�`�/rb�:3@�x��II��2G�(�S�'#�`x�,a����5��)PB�On��W�'���'����]����w�:�}I�C:31O6�D,<O���Vg��� ��ЕF}��3�'Hd#=ɥɁ�XX��^�6Θ��셫V���'���'����!b���'�'�W�N�E���A�ݶZ�x�F�:hd1O����'���င+p�#`,��p�mC�{����<yW�-!'e���_&0�i  ι��'��I�S�g�U�T\�qFG�0O61K#�����C�I' ��n�Tw m�eaF<5u��cV��"|����(�����D+gY�2�Y�<�bI(�F�����Sk�ũp�|�<�ԫ��(rD�aB@�8RRP``�v�<�Z�Z)�\��ݪj� �0�a�}�<�����J�k�K@)����Q}�<��L�v9
���+g&@����m�<)�`�L�|�9&�F̼e���r�<�!D�Nn�ݚ�ǁ2PV��a�p�<y�MAC�EJ��K6�-�c��b�<�`N\iJ5P�)H�b�l�b�_�<��Z��at
�*�>�S%��E�<��Hq$H����w'VX�<)���bw�0��
--�Ԑ��V�<��dw/���B�v=����z�<ɇ�ʂ��y��+�~�@	� Ɍ`�<�'	�p�R�*E(�(広o�^�<q��&Vf���u�M�5=�0�^�<i��Z�Fl}�B�t�)j�WY�<�[?ND|	�+Z�k9
|BG�T�<!�I�4W��Q��K�;<Z�NNU�<�7eܷ+� �&	}�Tx��GU�<9&L�
�l`�s�����pYA+�|�<�c�ɤ
��jQ��L���DO]�<���DK�|��S��z�,$�S�e�<!V�v�pr ��c��Ҵ�`�<9���4�8W��:W�W�<!VmL8au��ۢa�9�Z���G�<a5�F�N���2��HԠD,�B�<a"����E��+��s�f=�g��v�<���*q8��4+���)Kt�<�@f6(��4�`��Mإ�6��T�<y��C����z����~� 0��d�<��/�{���&���oÄ����x�<YC��*X��¢�\��J�N�<�AF�#^��)+BHHY �7��H�<��䊳s�TX�&�t�Bp qe�Z��\���q)(���al���f(	 K�-�T67�zb,D��ZE�U2��]�b�V(��+�I�f�F���qY"~
���"l�V
 =O2=X�O�<I�ř�@��A"�2�jɋ��ۖPT��J�Lf~���������=L���ӨY�>�� �85ӖB�I�O���
�-��H'�6i6^�p�I�o�q���*�O� �p�D,�<5D�1E8�وA�'�ܸ�"�B�|�`�'��p�@�@,�)Z�ڄ=cB��'���3BV,~����P	H��y�yb�QL��$9�ꑬ����-�Ӧ��Gh��4�C�]��	�"O6x���	N�@�ʅ�S��|
A`�5l�X��������!�	0v'B����q�<{
Bq�j��uV}.�e  D�����ǘ�s��T�i��x@�\O��@Z�93p\7M
=o�h�i�
8��)��A���h@cP��H���0�az�(C�e,�q�C
��yB�Q��`p1ᩂ�g�E(��X�|��x57S�0y�>�G��}����=̰��D�D/WL�<�ĬE+_l3d)�e�O|�ɃeB�6B� 	�Z���#�R�ɁaJ�K �6�'��x�Aŋ������B�EաɈD���O ˄���F �
$B�E�d�����e�REl'@���eh�<�1��=&A���A %�������n�#�d�
pn��3w��@k��?��S�ӤI}b6@ӿrJ��0��=�*C�	�a唅�$$�3L>���S�.�^!RFI8¢ЦO��D��O�Q��CMlt�E'�����'|�	q0/�=���U�O��JVf� sܬ�	3�F�z���O�I��d��U��tRK�@�#`BH6-� � � !�	�l����*"BȔ�,�L �E�Q�N���<8x�r��̘�jN�p�!��A�[4�	�a�.ÔA��߶v���uAD&�m�WR���F��~7>i��I{ލդ�
l��S��ֶ:q� aw'9D��r�n��� �◲Nr�a�r�wA�`��D_/d�n	��4,خ��S=,Ԑ��D$�ɋT:^�ö�;&��u�QfV�f�����6�Bt�D��6#_%0I���(�\�K��< ��U
ñD�hi�דJ���yw��f��X��kA)/͞���	�Ĭx𱨄�&��U��f�8���p$�w�uA �8��B�	3�XP�N�d���H��QR^�b��J��A.��1�C��!uhQ>�{�*E�1���&�[�/F�y�f�*D��
�� &��X�2o�I��l�`��$h8A�D�$'�>� �"ɢ �  �>���5F�Q��Z�\${�Ȅb�I�� RX��M���U�W���*B���N�"���×xTYQ��/ܑG*���azB��.I���aAD*����@�h��ۛ��L��Ŧ�yRM7`�ib4�>f�.x�����'Z.y�'�)Yu�u�F�O:�Ej���g��I�"��J	�'�\���C�?�,h�@�o�ȫ��D�_�0��v?��MNO����U,1�Ѳ���UD��n�w�!��7�aE��0�	�!l��l�p��
��8�
'���p=)��{?�C��B�0���Xd�X֎�B@$B�m�8���4d((�����sy���!���
�-� �	�b��!�B-E�.E�5钭Mƨd2૙�� �P��B4.��`�ZC>ɧ�Sk�\�A�i�k��Rr�xs�֢yl*B�	]�������)(�p��ʃ�F��O��7l�'kHă����w��1:�ċ24% l�҂��|��k@��f�az�hO]�4�@h�"ޔ�+uH�YQ���(�:��x$
�=Wd��M~"����J̓��:"���µ��&qOD��ǏA!S����RbD��s\���n��b����l) ��wA0B�I�|[2d C�C�M�b ʻ*p��@��`Dg�4C��$�vܧ7��̻z�Z��A�ԉ:���)�c���*-��7����(�	4�r�$m�0A�)��W$h����k�l�g�.�b�R���7A�Z!��M8^T��鉀9-��lZئ�0ōC���D2䭐2EF@U��E/f'ԭ�@�\^
(Q`Du8��� ��o\�"��"���!�!��6b����%�Y�I��Y�@�ab��S�ĈǶN�H
t헍{�!;�j�<��C�9�yK[�x����\���a��w0$a����g?��IK�z:�.H�<��g%��8B�	J7!���M�
�
�[d���N���үH `h0ݳ#M֯.o4۴�
�}� ��dL���K�Q�f�|��%I�az�W�~��(ܰe����3��#�.#�a��5J���ឺ{SX3���"�VȄ�	��!j��n�\kwd�[��c�\hqh�&;}x�����f�� /��]isl�6=�I��AgT(Á+�8�p��*S�K
!�� �m�~`�MS������@�]\�!� �6�2�'F���`�V�'c��p�;PR���/͟]���Շ�<VB��S�? 8�*U���	�b�1�E@!oy���҆�rUȚ�'(3���'p�T3$�� lulՓTQ/|Q"mP��� q���d�"5����'���B�\Q$��d�*<p�`�'.�@�e��s^Y��ꆬo5�,��𤖫%5�)����?-�B���]H�OI;����O"D�BP	
jN؁���T�h�@��d� ����,��핧�����@-k�D� NN�Q�K��!�D�;� ��dUC���#�3m�����$2�"N:x�2=�R�'�䘊 ��$Dp�� %8?�j�	�hy��R+(?�\d��@��c���Œ�U�H= ��޸��)9
�-�yz��z�"��gH�tN���?��ƙ10ڸ�p�.N}�D��ǀ��˧2	�L����0B�(a#	T�#����	����+J�m]z�aF]]ӂ����A�?<���ҭǩP��d�15O>!�wz�A$/�Y34��
����'����-αcR�m2� �C|t�1g�{�9"��C��!8�O�<�u�+T��HOı�҆�_��6B�,W���P�'[F)���q�
�a3�]8DӐ� �7x��IR*�v���O��hJp�"�O�L)T���{(X� S�(ڑ���D��6$t=�6�@2�b��\1R *�ճ4��$NȔ0b�ߎ�U�"Or�H�O(1#��Q�J>����� W�P�9$����#}�:O��;P��;ٴA��+%y+����"O�آ�D9m���R�>f�D���ZM��ђ��!j�*�a��QQ����	�K
X�tkǎu�<]��$�>&4̓O,}�G$�|��/s�%�C�� ���P��(p�����O�
����M�l� �ψ8����ݤF>T�2�p)C��HB���$ąbW�(�?���>!���9T�B)��+7I�	̾��'�^�zĘ�IE�tq�n �:[JF{���S�N$q&j3��?5���͞�x�pP	�M�����K�[W쨉#�0^��p
�;=�"|λA����Gm����c�߽5Q�I�d�n���Y���S�O���� Ǣ':.<���C%<�X�F�	J`-x��ӱ+�<U�W��,D�	׀c�����X�]��Jѭ�����Y��<��*D�V��Bf�DI�@܍�s�՟xG���D\�)B����ן\����
�<٢$HX�џ�B�($tV�F^�q&�Hr!ӣfƴ��Ś���'Q�y�1Ȝ�>c8M*��X9irvP�P��+�TQ!3B�ў�k�N���"�3���,OSA\���C�l�u���?K�Us�̔ڦU&�"~Γx���C #p	�zrp� 0��< :BPA آ��S�O��К'/�6O��(f��~r�@�O�X@S(Ts8���U�E�c�
h�'M m\�@d�2?�O�DҨ8�	ϓc�Π���vh��{6�SL⍅�ɚg�ހ�D�T�5 ���
��J�b-`�X���x�'�oIƙ�3���v��e�V�ު��O�Y��Z�'z��}�@��.;�HB!������by�萏"]�B!�Єޫ"҉�'�d�J�"�)ʧr���w�KF�Z��н�r���W�<�!�Fb@v���?ڸ��Q��7ʘ��u(�j�ߊl�ѓE�J�4��I1}8�bd�S�p%�q�2�շ.6Q�5	�1��x�oI�vy����i9����@7��O4-�eFt�����`�^�[�*�9�ȓ �Z�BfBA�<-��o^�_���'	F0�4D�}�S�O��Lk�Tn� �� B[b����'.,p�B�
�@E�3�T�@�N>���\���$$(�% B��+K�=�O\�l.�b"& h�K��ӬȂ��ѣ� ��Q���yH<Q�B�a��`ԄN�S��A���^�'얭�	QQ�G���0gϱ=��34�C�[�J���_+�� �M�dX�`��p�j�Uy�,��,3�)�'0�2��JѾm^���"��\هȓT\�Sb���Ud�+�&�|M��<iE&�xEayBn�.+.´��I��`�<hf"��y"'�rĠt"vL;L��ѐ$����yҍ��@$�,����D���ҡT��yRA�/zN�C���z��P�.܄�y��ʎ0}���"`�;�$��LN%�y��O�=�f�G吺,���Ekϊ�y
� ��i��KB)�P�v��?��YB�"O�-��ִc��0�w��#1u֤��"O�3E�F)����.X�(d��"O|����'T�~��n����"Ol�[�b\>���2C�i��"OQ�eV!H�d�+��� �ݺ "OX<�͍4r��W4ߺP�"O�9�%Mas*�k��Dc�X��"O���f�C��I�w�[�/����"O�EZrEC�Tx��톚m�hUXa"O0iҧ�	i�@	:�K��<r��+�"O���sHO �D����X�OgL��d"Ox�"�c��we��a��*N�h��"On��&��,"(��zTM��]��F"O�$c%�2gn��7́
�p؊�"O��(aA���� c�14��H�"O��*.�v�K�!�(4��s"OhIy��D�\l�	�Gv�
 "Oʩ� lQ=}c��A@��znXy�"O�§��!6�y*p���!a�`p�"O��q��W�����j�,&�x�J`"O��s�	�O�&�õ���Th�"O��x�_�����IAwͺm�"O��I��9	 ��6n�v�V` "O��b*ˤ^X-��d�*�#U"O�x���ږT�$iZ��i`p�C"OZ�j�ݓf~�d�UO� pg@A�"OքƃQ?E��HcF��{>�j�"Ot��׏WꐱE�x���K�"O���E��X��p��|jVT"�"O
4H'�ռPw�gB��$an9��"O�Y�@�t*|��gXGDF�!"O2��� �"���cg��7
�k�"O�Qy�FX.0G:X���*|�Q�"O��c7�L�bj���g灌*�J���"O<�� K�|]���!!˹3� E8�"O^������d
�z ��W�bm�"O�19 e�*μqi2�M+G��uy0"O����BT����R+�N�x�{4"O؍/).QwK�Db��� U��ybn��P�Pi�㞇COP �6/��yr�ńf��ҳ�J>��bQ+J<�y�#9�,d�'��:�t��ӆ���yB��0H��
�ɇ*���N$�yR� �'}���� #�����E���yn�*c_�t��Q�Fp�U"�� �yB��9;���fȮ;[��8%F=�y�0m�<�[eD��G�����$���yb���4Όm��)_�-�B�@p�,�y�Ξ�C�~� �޻RD\��W��y#V
+8p�P�_.J$�؇I�?�y��j��+�9W�EЀ'�S=�B�I����h��ـNnD��c�:�B�	_�B��cdٟsK*8�e�]% ��C䉾�F4�E��r��#��H�N�C�I<le������$D�$	!�ŏ!�C�I�p�h���f��/�~Dy�)�%��C䉱p�Z�(�-� /F��� D�J��Ć�'�T�C�h�Sm�y�����!�!�䉴.���01�ƑJ���[ե��M�!��?b����T*~�T谐/L�3u!�d�k"�qrˣr���n]!t!�$��!{j�P���*htI�M� U�!�Z�*��pP�E�'yL� ��^}�!�� \�`(�.vIK�d�-*$��"O$%�2���ʬq��(J�aI""OԈbMۯ3���s#���&��"ORك��i�ܠ3��,�<�""O�aZ�F݂gu4p���2F���q"O��+�K���J�����.J���"O��SDAΘS�4�QwhЫͤ=�"O�Vj�$�|�������1"O*� V9x����G�q����6"O��y�d�>�ܵS����e�A"O�ɪ���r(jy�B�I?\�.Q:7"O�%�/�19p ��Q�8�*�"O���@'
H�r�A�x����!"Or��E؆Q�|x�w��;'y�A"OF�r��tݺ�+��Dw0�`v"O d�$�V$R,)`"�>p��1( "O��)F#� �d�2A�k��zW"O���qhX>|Đ8G�O�>��`��"ODy��|��E�����z1"O��Z�k ����1��	D�<)B�"O܁���.s_p=Ł�2k} ����'j.,u oӲ�I�Z�1gMG�8��Ԙ��M�wl B�(D����V ����Is@W3EKΣ<���|�v#~RD�J���*��m���t&{�<QG��P��T�K$eD�@�r�D���D{��I�o��Dmy$�}!#f[�R�� ���E�2���4"RRq�I$c�o�<�Wl&C0��G6C�t A��i�<�R��D�F�0d&	2l.Z����b�<��ꗒUW�6�+���x�<ٵ뉥^ �j�nS*D��h; �Z�<�d+� XV0�K�#t���QIWL�<��(a8�p���ƃ����t��K�<���A�)o�)ГЀpT�!�Vd�G�<Yu�������iѦ{�"��Ga�G�<QsF�62����\�J���A��\�<��ŵfo:�zu�ܼL��-\�<��ݹ	���`r��63�M���X�<��iA�1Q��q��/8&(\�T�m�<���t����L�2+����!l�<Q�m�7#���(�Lհ2�L��'jZ\�<!G�H(� l�)�<u��A�<)*T� �@��M�\�t(�a�<�s�� $�pv�C�H� QDIA"O��"�5pHF!��¸[D��g"Ol��DP�h� Q"gӰY�*�p�"O��e
�:^��<�0�@�YÂ@B6"OH��"n� E3RtxpHZ$�l��P"O�22���E���(egҢd�Dq "OP�0R�j�I�6�ׅV��a"OVD�����i���qo�*�H���"OZD�ҶdD�SVo;��ѹV"O\���Dٚay�K��I<�!"O�����A��QV�{'�p�#"Ot�BO�Yr6A��NV��"OJ�d�\lbp���� �D<#b"O��z��R�!�*1�c&�s�:��"O
ł�q�>4��o��U@�"O��A򆁐d�b�ꢁ���L��"OE��@�a����M>"�04��"O���2f��
o�P���>�¸�"O� [��f�؋�/ǻt�R�A�"Oh�W"�k~Fi�d�R��Vd""O\��Ư��<s�}�LQ�+y�"O� ��rr�s���Xt��!BEp6"O���pY�d��e�Wa��v��#�"O*�ÐI�05�\�Q�AJ�<q��"On�1 K $���j�Lߜ;b��"O�#W��Q����w�S�gj8,�"OH���g�/����
�`VHq�5"O"W�q�pQ��(-�l�`���~�<	�&H<n8��H�G�-A@�9�� ~�<�f*���m��+Ŧ0%�]�RL}�<I��;Kpt�P-�9r�ƴ U�^q�<���e��4�cc�-ƦE��i�d�<�&b�"mN�P%��#.�����c	{�<aI�0v��eǓ�
x����v�<��GS4Cn�}�ц�h>�Ȇ@�^�<9G�ݎGN������G&��P�Gb�<�6B�>���� ��@ۜ���RG8�h'�H�Dr vYb����Lor�iS�.D��gC[��a�0��(*�`Ш�.D�P��F�2{rdX��\�_n��9��*D�pr�U��L��S@��|Lv�@C��>�|Z)�"I,inWT90�Q"O�]�WeO�
�ܐ 	êqa.A"O��P����4ZZ��ś7<�D0��"OF%a�)Tb� �@����1MN�y���#A���&ͧqV(�����y�$G(2YĤ��\�>q�a����y�#�Ty��
A�7B���U'�y���#D����@��m3 `=�y��ǂ]�ȍV�Y�k�&�" K���y���X>6��seg"D)�D��y�DJ�rЕ��"I1c� a)d!�y2-Ȉz�j�P�$��+� pP�'�n��UcrG<�I�j�'P�(2	�'��I㢡=4~�Y�j�X�
�'�
x�bG�C�`����1z'���	�'����n+a:��$ȝf��A	�'��-� A�+@`~���Y�iM���';+	�X�K��
�����|��E{��	���ʵ#���-��0��u-!򄈵%��c�膷�8P�A��u(!�OLp{���1R� |��̌o1!�(����!a��QC$��P"!�DZ�r��ə���1�͸��η	 !�Q2���f�5|�}���
!�D��F9�E���G�� ХD7P!�$7_�f�P��>�v�b+[�B!�D6)� <i� y�*4(���h4!�D��F��Ȣf(���zv��?
!�dO�x����˗>þIH���!�Φ<�D, ��]�	�� A����n�!�ě�8$���u�� I�u{��E"Q�!��&ݠ�C��N�c��'D�1�!�$��,�2�hI�Q

$A�b�V Q�<D{*�2�VgK�zMd�(�7&"��J�"O���-xmŸR�SMʈ��'��HӊĶm�,��D�l;�x��'�TpGƆMծ�()@h_���'� X)W"coF}z7苧f`���'�n��&�8s��%*���/Z����'���s��`6����S$QD����'L��!
��s1R9�#�8r9���'D����ߔ@9(]  �$��
���'�B� �u$b�w
ߋ9~��'�����/|嶠�c#W�Ү����� t�9���+ ���ZD�\ ��Ӑ"OH��w��"}�|��#!тI�("O Y£�İ!�x0�p/�z�U��"O��{����
�)�H�8|i#"O�Y�fE�f�>غ��NNƬ�V"O��������4���=�a;�"O\��s��8*�q)S*��3��f"O�t���F	)�:p�S�E�:���j�"O8��q΀�|��Hx��!����"O6�2��A�VB�J�!��^H)f"O09�a�:wu�!
RA�!-�܁6"O""7*�B%ڴ	QcŰÖ��"O����j#l�0�sh�z�(�u"Op��J�VC����T�@"O���0'
G�D`���?����"O�}��
[�/\r%eV�er����"OT1�"��iŞ@;V�גz[~D�"O*T���[-M��L�'��
S���a�"O���q ?<��.L�Pz�)�>&�!���"F�<8��k҇�lT�Ro��!���5%��!��%�7$�Y�mD�a[!�+M�y�k��:�d���DER!�@*\��(F���Rhr�<r�!��Ѐ�����nA4W�z�[g���!���UF�p�RN�<5�Ru�� E.�!�dZ,h�l�GB:p:H��O�)6�!�D�������Z*Z��7H�S�!�˜=\*��Q"�
%��
5�!�D^�B֜��(
*] D�R#Э^�!� l�Ȓ��$Q�Yڧ�W�T�!�$�U8���^O�y�m	;�!�D0�X��h�9<�̈Ul��~�!�D�5�R\qUh.y4�9�Ʃ�=�!�� $�֑j&HW�0!�$��ɚ��!�D�����*G~���Ł�z#.��ȓ'����T�]�&'�yؓF�rᆴ�ȓ#���/�+~�4 t��6����&���ƧxO�HdK�^�\�ȓ0����)�kk\A[��G�S� ��ȓ<(%Y�&Ʉ}f���M�2�����A�,�Q/Y=_|٩��oYH�ȓK�U	Ei�W��Y�D�H���ȓg\��"���G"|$�Eꗏ/��9��,�X�
E�ZE�0��.�w�4	����܈�	!}�bΊ�W��x��@��p��H�5y+�u��� ��$���x��F� <�Z��%�E�Cî�ȓfc��rs�PI(	�M��5&���ȓU�I�MT\.l෈�@u͇ȓ;��űҡU$}4u���O�G�Bȇȓf�|� )F�)7��[�'������%^,䉅ć@�
F��R�P�� �j,����j*�2�ɋK��ȓ>����*�<x��a2d)��B��T�ȓgRa�q�Y�y�� ���3\�P�ȓ'�h��o�)n�(�`ԭ �v�ȓ=v"��M�+e
$2�m*pòɆ�0�ʡif�/=
š#LE�g��a�ȓE,hMY�)���D���yrXd�ȓ>%֕���?��H�4A��ȓX)`\��D�!@#�I�!�W�)��ȓO�nqh��V	<�J�p��Q���ȓP��Gh�>c#2��@W�?,�,��E׎����2��jgK�6�݅�S�? Bك�¨˘��S���f9ʅ"O�0�����(S�v��#5"Of��*K�>���q7F�$9�b��u"O��� -�$̙�JF!c��0S"O����EQ�=���X� �*�a�"O�����u��x@�N-L%bB"Op�I���M,�̣3���.��`��"Oz�h�.�&��y�	\0U���ig"O�iw,�Y�]  gH� ;�� #"OL�8$n�G�j�ӷFQ8c�@"OB0�W���@�ΡɆeˠ�t�c�"O��@��'�B�D��K���"O4��Ռ�(&0B��
��E ��J`"O��@�O�#>wƈ����2Fd%��"O\�z�o�~^�t�C|tB�"O��X07af�a����q8i�"*OZ�(�͕�^��S�E  �r���'f��tDż�bM�2�˟w�ݻ�'Ol4�R$
>Jh�q�rE�k�|Y�'�V����90��1i��,4�&�S�'JT�Z�f�0��Y���Y���A�'
�����A3��st�:L���
�'v��i�'P~�p�D;>ab�'�L�!f�����"7�8|�
�'ZF,��MPK������cX\�'��1��,¬�%�X�n��a	�'�0� �U�GVT�%莢}���'J�A4Ƥ�I�b�8q��k�'���6N�Y<�'D�<gfM��'xh!"J��F��=�fĥ;E����� ��@Y%;�-�Md���ȓt��A��j@-SI�mIQ`�-�Nd�ȓ<��\6႟%b�IĦoʴ���he�!��nX�����x��ɇ�~x�vL�&j*s��=Q�t��[�dE�W���Jj���΄.3N�Y��n��+`CH�̔�Q.1ޚ,��_d�94�p!�b�نȓyc i���+�L���epa(�ȓ*M@�q��t[�tx���& RR}��z�T�jAoʒ@��!�2���=4����K�"t�CeǩzIX��aj�kv^	��= �	"�^Pm(Mԅ��P҈,�ȓ\˰HY�m�Q����Ú �~�ȓd�(�6Eˑs�|�#T�ڇ?����~2ް*�쏤#$"t;�K� ��х�f�`��&.)���a�~Xi�ȓ7�P(��,����>dN*4�ȓY��mb�@^�Xd��S`/�x����2)���b�6_H(��n !d����R�~e�r�@"���;�E�L����ȓS�Ճ4g� �t��P�-H���ȓ+R��c�;V�<� J�3Z�T���rfLE%D�/���蚷1Q��ȓRi����_4T���(�Lńȓ}F��1��pYd�q�C
BH�D�ȓz��	��B
7(�jԡ��R+J��ȓx�y� t��%s���Mڎ���u�r<X�*M�aP�u�Wքj�8��`�~P��HB
5���!G0
ńȓԐ��J�0Y"�]:�W�p����q6���+F�dzpRGH$�@�ȓw:\��(>#^�pj�A�]
�8�ȓ|�P��a�
�R|�0gM� I��S�? ��@wJͤU�%pUkG�E�:p��"OX�s�I����@��A�}PV�#"ODH�I]�f���B��F��|�I"OR10�AV)FLN�x7g�H���y�"O
.¬$WJH��y�tX 0"OZ�x� 0Nϔ4yr`�%6>B�@�"O$XAC��?���#!�S'�<��"OI��KE�aS��k'�%g z��"O�����-G�]#X�%��@"O>`�pI_!
x���B��a���"O�ua�ߊ3y��;��v �{S"O��[u��
E"������,��"Ot�c�/���QVd 58�\��"O�q$���f%����%R�A0�Q{"O�R`�O�\ b�B�rV,x�"O����mV�>D�q��(M�^�!�"O�Z��U<+�=� �Y�(
�%��"OtM5$LX�+U�Ѭ��u"O�8 �-O<F���2\#m�$	��"O�AZQ�D��6�BQn�-P�H!1"O~���I% ��h��#B.�aw"Ol��B��9|�f��E������""O�1TM�Q�l ����2V�i�"OԴ"���k�<�Q��I5� �!3"OV��B��]Xn��C��M�<QxF"O���d�Χ���F�ҕ �� B�'�!�$6K{���	�ZF0�q\dv!�DY()��� �oZ�RT��'�[��!�:�d�W�	�?K
�K�Kԃ+�!�$��\z`�����|�(�C4*�c�!�߶��!#*����P&�i��}����K	^0m����$یs����(=D�|���1/|�x�iX$4갑' �<9
�K����R�Q�w`#Acƕ6%tt��<�0h"��n�� ��-b�4���KU!��h���=	�:�0��6D����+k��t��`M:;�֩Y�	3D�l*���{
f����
W7�q1��2D���p���2=ؽ��'C?ti��d%D��5LF3,��hp���K xT��%D�yE�אFg!�3`��C�b,Z�e$D������<f�9�K�2rvd�э"D��e҇ ��@�I�l4H-k%h;D��"���|Aqg�e<���.8D��4"��([b

��z b�@9D��j�C
`�9�@��hlJ(��3D�x���B5~����L�� 4 ���3D���J��(�wg^�`�@�XAK=D��A�f�Y���߮	�X�p"�/D�T�1�FO�U�b^.��1�u�)D�h �[r|1�_ߖ��0�'D��fG�2+!¹���5+����t�Oأ=E�$�	"��}H3�ɲr	�P-ۡ�!��4Q�2A�%lL���a ,�A!��lx,`2�&����W�4�!�䖙U&n���- �Z2�p��ч6n!�D�ǌ�bjĀV� �3��2X!��X�/_�yc��4L�rd���D�I�!���V�(��'�)�lDR��ؙ.�ў0��I14���a��Q�,	 X�"c&C�ɤW@]���n�U���W�[/�B�KfHE����c�<��	UP��B䉟m �U��5`��M���{q�C�tU���v&�K|�]8�&ҁQ�C�)� �@+���9g���S��/w��h�"O��cE�L��H� ��6\Z x�F"O89"�-F?WTB� 'f%7媙�"O���s		�3��1�X;�x��|r�'��h�F��3�JDbӇT�}��'x�'�s���bB�A9|N	�'��� q��l��ךt��MA�'U��q�<Eh��)g@ڤI�'Ǵ("qI�'v�!�5-S��@A�
�'>̊��wH��ď�4ИӉ��'O���<!�`l`WΟ�1��M��"O���뚋9o�48u��+%����"Oeb�e�u��`�����"O�� gn1=i.�y�IY	�*Aې"O�����R0�^��(I� ��`�"OF�+!l�"�t�!��Y'��@��"O�x%���p�$�Bc�=�6TRO�԰a�֡l,\Y��Q�MH"-���/D�d��mF�+�ꨒ��'vy2��"D�I�*R'ܞ�:�G΋K��[a� D��x(�7/n�Y#F��o.Ph8W�8D���3�R�s�$p�l�~�|�bN9D�8D��%A9d̀P�E�y��+8��0|�`�pc"	:�HQ����@
�l�<qUȖ7yt�x�D,K�e�S�Xӟ���m �ԩ� 0-p�E(��5�ȓ�"Py��h^Txx�JU&n{Ȝ�ȓ� �RJ��*R�x(F�O�4~f`��O�V I�Ăd���ɒ(�7V=2݄� �0� ��/r^�6g�2A
�ȓA�&x! �L	R ������.^wU��$��Ti����k�i:��'�a~"
���@quG0Eӆ8�S'P�y�����x��6���7[�|b���yªJ���#	��Fdy�E��ybKǬRm�(a"���9Q����y"�WI\[��ĉ�2�� ����<ю�V/z�4i�\�MM�#� �-e�!��3I
�1���7�@b�MT!�d@1K�0����;$@D ���ǻ!!��o�V�Vb��H/6�ݒ_�!��V>" u����#�+E!�$�2	�q	��B,�@���A�!򄅨�a�L�*�D�wŉ�a�џt$���OIr���j��/B�؇�H	&t�8�'�h �f��>��3�ąa|2��O�$抑2PG�� D=s���`�"O�� w�Ian�{�/X�G���3F"O��Q虦5�ڨ�7���RԆQG"O����/¦Y�M��V3r���"O½�B�H�4�d�6͌NԹ
B��J>y� ?�Jm���ל}�bX��"D����Ț:m A�C���D�ڀ <OD���ON�U��X˗E��NJ���׋Z�i�B��h����A�k�B����%y����J�`dYU�
�xɂ�͞��� $�R1a��h�p��3�KuI؄ȓ?�2I����O���x��D攄�\�����ZE`@��)��Y�����jԒb�C�|�Eh��ÕvH���L��F��q暖n B�Q����-�ȓ��!h'�S� `8̀�%S�REFl��bpN����PN�@�� R��ȓ`Ζ�+c��pB��z�O:E�D���S�? �zG�L��5�p+\�D!���|��)��"�b�pU`�'!\Ց�˛>CJB��3E3j� WB��O�D%i� [.�B�� 4����B +h�����>p B�	+y0F�Ʌ�D
|��u�e+��X�C�&2�T4��{j�E�w�>g�C䉯2��=��P�Vw�E�B P 7|�B�I;h���3��ɼ�~��I�=H�B�=;��!�ր�J�x�񁦈�j̦��7�<�'�U�c�e��#�/�Z|YP�&D��נ��g�a�(�#J��%�0D��+Q�	�rETpiW���I�����;D�$�-U�(h�#�甾e�u�@�:D��d$�n�@Hfc�Q��8D�H��L��'a���jO6^q�UK��#4����A2 �d�u� O	�H�`��ßh��^�HqC��A�d����pN�2y��'���l�)�O���ԭ� j�hM�"(��c�fa��"O����O'���:P�L�5�$�Q�"O��a� M>KJ�q %ا���c"O��ڂ-J#u�)���/}��D�S"Oʰ���J&`"��W�
�ww�L�&"OL��'����]�aKD�Qu|�\���� ����7�<�*��%+t��-�kx��Dx��ؐw����6�ܚC�f�q�ʙ��y���`�x0�D*i�(A�눗�yb�Ӳm;օ�%�G;Z� |I��	�yrO �3\!rD%F�VD<�c��X�y���=7�Z�w�T�ۤ�п�y"18�ؑ��鈩J FZw����y�CO9ے��!�͆E@޴#C͒�?9�'"�% e�ܥ��+�"��f]��(�'&���N�B��G� �X��j�'�ŋ��%	ʸ��	��z`2��	�'�dD�0 �44���2ƅԘ��E�	�'�]1���.lV�@�p�-u�)	�'�(�c�gѭMY��P�ꖗ'��!�Ę��� r�@�m��ڄ��?2�!�����	G� �.0�Z,+�!��Ҧ7�|��M��jDAp����!�� y�\ ;�J�	\V���2MƼY�!��Լ�-E�@�%�"�?s�!�dzт2l��Z��h�3jC}!�d֙ ����p���#	�j!�d��2����'GX�t|i��z!��#xE�!��	U@Ҳ��ŕ�s!�dV�W簴�0��6!��򳅁�pV!�$�<]WL�]�t@��o�u��ȓx�l�ᵎ�.{��[����z�^@��G���?�����rx� �e���*Z�%�T�S&�B�ɿ[ݨD���.b�A��Οk(��D-�S�OT�ʗ�ڔZ�,	���G�4;"OdU���4U:0�X��_:U�32"O(-��@�> ���:�AG=,��Y�"Of�*� 6~��˚y|��R"OL�Tգs�K�n
gCΡJ�"O���'��e�4]*C0N �$"O��S��)$`������nc����'�ў"~�F��<��Q�&��%
�C1G��y�gS�Lt$Ѵʖ�k�%B�ϒ��yL˫59�\
�>:�ⓍF.�y������Rc�}!��r���y�-D�b�@�Hv˞�cz�$��	:�y�P-xbt��Mǌ\X�1Q���y
� ���! �0
}f4�cJ͂D��D"OZ�ɂ��f���*ӏ[$:�K"O$(�#�1�uz���D�(tZ�"O�yᤂE-M?TY�u��*<$�<�g"O�P�0��f�*��3�.���*d"O��IuN�7�4��$3�f	��"O��O��e.h�Av��,�`��"O��b�j۩e6��S�� W�T]�"On)�ڿl|�����HԺ�"Ov��T�:�Ph�ɛpoPT�1"O*���Y�.�z�Y�hHK_֤1"Od��$Z?�`��OT��B"OX��/a��1+$���+H$<��"On��1����b�&�=FpP{W"O:�G�Ԙ~����5f��  !��=�S��N�V����b@�,Lt�X�]�[�!�dR�z�n�YG�0Q�=����(v!��I,�|}p2m�[��P7 ^�vV!�$V'Y�aH"�T�2��LB���/�!�䔥
���A��VY1�P�t�!�̱h��#��сJH�z���Y!�@	!(�e�W��� Eh]#��T�K��'B����b�8�zW�E�A��􂵆��6	!�dŉ6��g@�5�4��1oŰ�!��_�jU��z�ds�`�?/k!�DT�)���	�̀)'p�5�`Ɗ�?t!��Es��X���Z�
#/3l!�d�zar\��cåW��K2��W!��&�tQ���~A͹�6!��5�e�u%��`I'-J�1!��M�P!��cS�Aw�s�bP�R!�d 6�x�1A��Mc�uD�N$o�!�	Y�$��;J��ha�2w�!���c�㯟��	�`Ώ�Q}!򤂢W��xuKO�O�̔z�̏i!�	@��p,�s�(�x�S��Op���5���{b�3����ɗ�!����q�Qa�NTf��䨝�:�!�$�R)|��AѺ��ԱQ�Y�E3!�L-dj H���|���Z	H!�ě�mN����[g��2�h»8]��$�/;��q�&�aT�Y�+�rTC��/èŰǂ�S>PP�pn�"�r�O�ʓ�0<��.��Z�~���N��δi�
Dj�<�X!G� Q�6������n�<��j�&<@>�A���H=�(i��j�<!��@M4q�u͓�N�q���<a�nźy���;s�*�Z��t}�<���W�$��u��&�#M��(fK�u�<A�mZ2�:��
6A��]�l	M�'pa��&��uJ����J3hXr2*
��y�$�278캦"�O�����O�y��5q�8�K��ϴJ�z킖':�ybTwT��(��=6��s��y�i3z���4��Ds��������x�N˚���J�E�%h����B�JG!�D�%Dyb�2�U$\Q��s���{9!��1���ϴ9��PӆbD�H'!��WnB"��t����Pg�7t!��UHn$Y�ز���+L54
!�P��M��@Ʌ��L��*U�)
!��M�P��i���\����8x��">O��re��9��4���X� b<@�"Ol虂�)�E ��b��A�D=LO� f 9�oM�Hq�5 s�(q�&�y�"OZ�җ�ʱc�H�ԩ�-*J�4g"Ox�`K׆DY@Y#3ȍ-_. ��"O�b2�g���#�ٮ[d,�J�"O��ru)S&l�y�(ؖ��:�"Of�Ug�3!�"@U��X嚘A�"O" �F�Iu��8 �E�h�t�"Ovt�AR7(�(@`Di�&A�6 �"OP��APi���Ј:M�4�"Od`
gf�z�.���'l�((B�"O��(gZ�=E�a� �U&~�R,�1"OT���.J�S�t�X�����8�"�"O��ʢ]����f,?81�m�7"O�)�#�p�ڬ��!(R��#"O&�8���+5��P�����D"O�b��۷9Β�+���"f����#"O5�d���kU6)����h:���"O�)ʥ-3xH �'�,����"O���@)�5)l�8x�%6B��-��"O������*Onm�s$�o�
5�F"O��q4ɖ5���C��t.hDZS�|B�'U� ��K�%!¤(���61�8A	�'��l��:Z8�)��!~��`J	�'�4�a�K�.U
�%�!|R< 	�'����%  �q�-Ӫn&ʅ��'��Lf�C9z	�:Vn�j��	�'���j��P�j��zp�ŭ\��ц�!�q�A.�=]�ܭ��ԬS��&�܄�I���8 <�ɳ�J>K�~�b�!��Q����aEE�)ZO4��@��PK!�F{CVH"U��,0�I�@πZ2!�d�!�8"B/�	��Z�/-!�$K�Q��6K��i�8<�@&�W�!�D@�|@�����4l"[�d�-+\!��L�Q������F�J��Ѥ�4U!�D܋
�q������ؖN�-T!�͸�����h��()Sm�#�!�/o�b��քս1��!p+֨y�!�d��7⠥���ߩ(�&�R҉R�I	!��4O���5�>�P��P��!���X\��ٱ��02gj��wM!b!���g �i�QA�#x���K
L�	O��(�$`Վa��I[�ݞ+=b@2Q"OF�8�E��1_ʤցQ;�i�"O<06D��)��x�ӯ۱!���"O�%pC"��6/��[r�B*+�Th�"O�Qrk�)ɶ�c��A�L�a�"O�%�@�<,��@	]�:���bv"O֍(0�P^H���瘖n��I���6LO���5��	������5Q$�5"OT�AgL;��8��_#�,�ZT"O������a�M42;¸��"O��
P�6Z>��!�|�J�Y	�'8�T�UJ[�V��H��B�E�V0J�'Ap|�`.]�2�tlH��ԟ@3����'�����6*�I��"�=/�!����'G��9p�	�c)���@jP.y���	�'4�iKA�Qjp������4�R�'�2鋃E�m�<Xc��؇F� ��'|ν��I�i+��E��\;�'p����F�~
�8(�D�%�Z�"�'�R4��~^�����|���'_�����:��DHυ~�xMa+ON���S�3��is/�"AsH��T!�� "��W��2f.�TV�Îc"J�0G"O���w�_�p��#�o�&r&\"F"O��2��	�B~T��&,	�S��7"OhYK%*.w�N�ӗ��9d2(-I�"OLI���>�Ω�B�M%/|9�w"O�h��Cݭ;L��2f��ky��1@^�|�IA�'81O���� xb��O�tw8``�"O����*;&��l�4ZQH��"O��j���.}RѰ���/[Α��"Od�{�/M:�^<�S��m鶰 �"O�!�w��:�x!�S.�E�4tAT"O�xJvaZ�N.�X����}��D�r"OX��?X���BKz���Y\�0�'��'0��:��18������[>��b�;T�LCGǃo.ddW����lS�"O�	 �HP9>Tl�2��>}��Ґ"O԰Q ^4d�p��-=B��"O
���"��"�I�mڐ�J���"Oh-q�OK��{!Վ�� Т"O��Rd	89���'K@0
 ��6"O�<`0,ܰ��jU
�9眅�w"O�<�7�U3J�q�a�G9^���+
�'gnyA㩎,��)�SB��^���3�'�� `Q@�h�3�!)FX��'u(���FV2���˱J�G ���hO?e��ƕs��i��/Otv���E�<Q�GЂl��ȯf�:�I�@�}�<q��&���U�C�W499�Lv�<�a�ʘN �I�0h@#^2
���.�o�uy"�O��5ZW�=�:�#�e)O���'e�Ƀ�K�����*���$�b�'ol��&�5;�Mc���O��Q�
�'l4ib�3(�1��W�T���	�'}(�����)2T��e�����A	�'�TaH�8&�����o�$Z2�k�'8��1o֑Yy�4"��N%H����,Oң=E��ƅB1�}���
mFM1	���y��T�$���0L��+�k�y"V	A�؄yp	^2�^�K�����.�S�OW�%Q�ΐ4���a��2<�
�'�.�Xqk_�W����ǳT��
�'Ćq��^	#��}!&i� �Pc
�'�0��!�:j��=H�.	�}w4mr	�'C�q$�!U�ő�����M	�'k*�qV��6/��QsbI��	"�'�v���Cv��yRƊ�k. �	�'�ip�E#w>�A�pM������'��95C�qKd1*�h�i�Ȁ�'��,�� � 2]*�bT$"lx�
�'G��*��J2>HZ�MݦuG��
�'{�A�
M4����ޚo���	�'̮�3@A�.%�����%X�d��	�'�T���ӭ��\���Z�Yɾ��O>����	�0+ߌ$���q�:!`	�1�!��_N��}JoIz�8UBC�M�V�!�ć%-ƚ�0
�;G���7,�>3�!�]k�@���O�/���� �9Y�!�˩6�н� �E
zep��.�>hQ!�(f(tw�L;q_dX�7M��=]!��na*EhJ����'D��`��T���	L�S�Oc^��A��.A\�p�M=1�J=8
�'>�eⅎH�N"Bp��5�x`�
ߓ��'�$�+�&��2=Dd�7��i��	�'�FdzAHLSs��B��	wPp�
��� �5�r"�Th`QS�ȅy�R�rp"O �RFA��PXC��%D�X@�"O�I¥ΰb�8���f��A�D�'��D3�L�7/�č�5GЅL%l�2q��<َ���h=�(ak��=�*̊���Y�*��D"?���T.�z�!�L
 �T��!e�\�<�/�Q2�8.����s�R�0$�Y��]
(�iRv_<��`Z ��̅ȓ}����c� `�t��ԍK#7D�X��G�-H�Тhv�əs XQu�ȓ�E��%�����ǘ� ���ȓy��AčJ;N@�-�JȈ[F�ȓ>Ht�Xs�;5b�-���P���ȓ,7���0��6�"y ᝀK|���ȓL9��G%C�$���R�!6y�ȓhi�i�qM/t��Aa�$M�`L����m�(*#ȅ(Fѕgs���\��lʡ�P U�:�i��J2&�B�ɠ|}�����@�u�d�"Ǉ�lb����$?�4�T�$��le(�>/W�Ys#�v�<a��UR�q��&:$�9;��_H�<a���[�	b�8��r-�G�<�/��p\�e��˯.���2Q��w�<ɴ
����"$�ÖeoV��e�v�<�d�6~v|Uq1�+��s�Lx�<�䔠S��h�R�}���"��Ox�Ȕ'��ɻ7 2`K����d�:1UI�F�RB�kcv ;2�T?B�����̚D��C�	�+�8��D ��r
�8�iͦ>e�C䉱�蔠WGF�,�*�!��f��B�	Vz��C���c�4(Z�J�,Q���$�<1�'��,3�	J�Uv�52g�	�5��A�'�8��@�@�b��E��,{fM�)O�O������Q��.�L��wͫ r!�$����o�xN��/4�u��"O�D(�(�>(4���޺lp��"O&|A Lt�Щ�Y�oP��Pu"O<9���+2�L�!�Z��F�@��'��O�8BFĿQ<��2�j59`���)!D��X3Ɠ(f"Sԇ�skJ��!"D��� 醣u��p3�V�VbJ��W>D��xuh�7���� �:]�b𒐦6D����UB�鐵��4K4L"�0D�����T�nXQIu���N���-D�d �2W������~�P��	-|O�b����ܩ2�$}["��2&&��G�?�O<� ;@1鄉[�6 l���
D?C*8C䉦[Y�蹤�]VMH �Sc	M�C�I�Q�$�� ӆG�2 ����9��<E�t�<�MHR��,Ps
8	�JO�JB䉞5�ru`��C2I`�9�6�BB䉯�Й8� ��2���cp�\'��E�t)�>�T���D�hXԲuW���=�S�O�@��n�cI��M�NJ>LK�'p=@n��5����D"�S�����'�<mI��ϙI ��.ѝNZ�� �'�a�4`Y)�ĬS��Q�GƎف�'1�Ļ���o����G��Gx)��'��Q��l�g���i�܄7�.Ey�'���k��Ĵs԰�хj�)˘-�/O��=E� �"�*�����4\���)��Ț��=1�y��l]4�h5�U�[���ȇB���y��Iiޜ�s?&B��.¿�y�)M$q+̵XW��$H0brkƳ�y
� ��Hⅆ�K�̀Yr�<��[&"O�[���,�ɛ�i�;Gl|Aћ|bQ�ؔ'�>�I僑$J8	`F��^z$���(�OL�g]��S��E�_�4-ko�;^�L���	�<�'��������q�\�S�Eu�P�'���Ѳ��*�h�iH���$3�'=T��L:(�FH�"�za�'o�s�T�еx����b"O�ABD�N�f�ŦG�!e�љ��'C���`a�P���#��/J�p���7<O�ʓ����=X��Qb�ؠjT�閤Z�0�!�'�� P.��A�X3��*�!�ױ6Ȫ�q�K�w�l����+m�!���^D8�l�+CXp���E�	�!�+c8��c��G*��I7臣�!��"?w�%9��ܜ�����FG��!�$H�Wc6Tk$ezAN�s��J;�!���p�0���ɗ�+� ����	"n�!���'�:�k��Ś����q�J�!��P�{�e�=�BQ�����!�Q"f�6 /Y"q'	�<��'8�}B�k�<R�dp�W�ɳ-z��'0(F�3>��1��ȳYޔq�'��1����Y�  uJ�^R)�')\T�ؠL#Աu�
~>�1�'FZ��řY?q@/�2E��`��'�^��v�W$RP�'�<�����'8 �3�f��	ob�CV���.���	�'��׎��sq����E�%��y��'֢-C� ��1�T��˚�i����ߓ�?	��y"�:^�֦BJr֌�UL[�yҎ�>=0�GC�Am�"�A;�y!E�/"6����f�(�DҚ��d?�O���F#+�"��E���(F@�"Op`K�(�%���!ȿ&�3�"O���@]h*�<2�o��%!�C"OnH��̹`8Jm��/U��!@��'��	�<�@�jNI��+D�����
c�'�a���
;as�43�l�?g>��GO��y2M��ȱL�9M�j� �Mȶ�yGf�Ό �068���*L��y�H�?8�T2!�͜+������1�y2�M,>��	B�#)`��#ã�y"4���"�D
��%1!/��=����?�'�b��b* O:�Au&F��#���1��a��"��&=���w�[/D�$Q�&"O�,P0+�T�L���ʟa��J�"O|��M 0A�!*VK�`�h���"ON-�C@����r�*�-n�����"O��i0��;|�X���N+����"O"����=��M0�Z�%�Aw"Oބ�f������5�?���"OKթyv{p�̹N)�5jW�ފ��'�ў�Oj�T��C�M���鑰hp���'�z٣�\�	��Q��EV`
x*�'V�Y�J�8p�E�Ñ�U����'�b��e�)K��k�H�P=Թ��'кc1'�]����`�� F$x5��'��J �Q[�d�Y`@�����'�D�� F\�$��m��*��؀���)���ù���3
��e{�� �*�3�y�N[l�� Ȅ�O�bu���&�yBEيVOzx�֡@>
W������y�� AR@�[ ��1�1�ׁ�y
� ��(v�R:C�^}�ொ.G(<�2P"O�Q��M�>?�z8.Pj��=�e"OԑP5�Z)3dyA�"|§�|��'*b�Os^c�0XhV���X'����'9�aZa)��3?�=���x��"O���ьŌ~ð���b!W�Tl &"O��+&bB=πIX��.v�4yP"OV�)v(�!j���q�j���"Onh+��� gP��Sԣ�7S�����"O�Pw�(iDę�,�l~f�IՒ|2�'u�'�?U��V"6�VDK!�Z�[��Tx�#�OZ�ɡ[�p��ʋ�i�褓G�J:H
B䉦o��ӥ�T�B=�+�-H���C�I<xH$|�S�ҥP�(!�bZ�Kz�C�	D�����͊$���k�dX�
&C�	�`�^t�?]ҾI��.�<c����!�5P��"&�2y}���J&F��ȓ5�H�y�b��!70��E?�b؄ȓZ{T��A�?b)8�e;E�u�?i�B|*DӶ^����q.��C���ȓ<֠a8�ʤ1�2 &c�����=HZ=�jJ��T�B��긄��p`Zn�O-h�!�@�e��؅ȓ2� �"+��%���P+� ,D��r���)�����]�hX��)|O�c��K%I�45�|�+�	(��4��L9D������FDZ���q�3D��[@��-��lz��ٚj��2A�%D�`���w�D��a�-�PmCE@#D�tC�M[<5&��$f��!Y89)�3D��*u�Z�"��� OR�&S���0D��-�l�$�q�P���T�Ĭ/<O����OH�/��}x�ߚs�ݩfD�����u��m�%cD۴����;#��ч�h3��g�=��d�j^�%�ȓ1�~预D�=����w-[㢅��H��I!P���'�y+2��1$HЅ�hm&�:�E�=z�.d� ��B�꜅ȓ�&)cF��W|��;�#GR�d|��Ib̓U�(+�a� nI�hcìH��?s.(ac�'���S��[��A��|v��AjĳAo��Gi�e)��ȓp�4!�A��J��VCVTe��KJA�n�': ��,�? �Ԅ�k���h׀M~�3@z5�`��?2ܫF,Ҟu�l�Aժ�!:l���ȓK�6<k6K���*�R`*�@�l!��/����J��-��AѲ�P�\�X���!,�CUlP��xk��X/�l<�ȓ�n�BF��o�����}TB-��h�^Ys4U$f̼�1p���[�ry��O��`�oL"��|��ґH�ĥ��m� U�u��B�
4��w�H%�ȓE�͉�i=J?b@&�C �9��%3Z��CK�x�D(+%Å<���ȓ'������%pF�)�G��(��ȓWY�@��ER�s�JP	���vz܆ȓF��M˔�!��؃J�?mm��Hz���GU�<�a�',\2Ժ0�ȓh�&ՠ
�xp��/g׌��ȓ�>dJ��Xt1<�@���-�*��3r�2��>}�M�oޔm}�X�ȓ�X�6�
�\~f�&��T�\��P
FHv ��%S¬C7��m����S�? dY�i��{�5i���M(BPٰ"OJ�cgɉKR\U���ٳy�S"O8����S�#7����IQ��P��5"O���6��7`�0�kň��`M:�"O�uA�
4U��19�&͖@����'�h�.ދy�H�Rn����	�'0x�Rw���ID�E@<��'rH93U��]�(� �E�7��'D���vJ	*�A�O���o+D� 2sA�= �{b�ɨ̉AB&D�b �V�4��Q0"씗�ژ���#D�\��$޸vF$|p4!/��$�,D����e|�̨P@�
k�4I��J)D���b_<,��<X�b\<��PJ(D��C�)�
*� 0�B�z�t�f8D�(�� �6���!*N(<0!��7D�4�p*�g�ddK`I�-'��]k��8D�@���%?�>���ŉp��ܛ!�6D���ָ7���q��:��0�b
3D�p�c�	>1f�����4Y���5�$D������tXE�ɤ&``*�!D��;�d��/�mx���w_.a���:D��K��	rF����=eZ�9D��g��*@H����9ƕ�07D�́.�=d�:[���_��	P��'D��×�>� �HAM�37|�i�&�$D�\�D���Cfh ��dǗ���E�?D� �dA��4i���!'P�P(b��2D���"�HQ�q��w�"D�@�%D���5����̊�p���yd�C�	�MS��!L!D�j5��#�.T�B�Ʌe���R�eZ�L�I��&�@X�C�ɽh�� ��b A�8d�-fB�I�I�����M�4 ��uY�EF�WH8C䉑,���06lL�.w�!�c�5p�B�ɍ"���z7)	� ��i�
�~��B䉰��t���V$Rm�|y K��5�(C��O�8������B1(q^C�		��Y�%>Ln���)b{@C�	�:h�*��˧D��@
"��C䉩dbi	7�Ƚn�ܡ!.�C�I&F̞�Pe��e��Tps�J�C�	�:M��Auh��%x\�˥��&39C��5"80��>H;
��C�O<C���	��ݺJ��\j�_=!��B�I�C̖� �f��z����ۙ �C�	v��Bu+��Vf����>AB�I1(a �1bI |�a؄�e <C�(w��&��bV��a%쓕m=�B䉒~\x�UN8d��l� �sV�B�	��\,�2��	1X@6��^��B�	((mz鋇3]O���@i � U�B�ɴ<\�����ޡF��Yh4����B�ɟr�|�-�
at���[�B^�B��<!Ĳi.ە�P�����C��B�ɔ,d�@�d9\n0]�AkU=I!�;Fe��-n�9�	 �C�!�䏎&���4���TlhAG��5C!��1!�n� ßYČ�!��/A!�$�(H<5�K[-g�"��!B�L2!�4pL����'���hg_�;!�D�Esb]�ӡ���y�/��O!�Nj:���hZ\وH
�N�V�!�K T�H�{�*��B�~� r����!�� hi�F��Od�]�0�_/�6YS"O�!:Zp fk	1���3"O�,�`B���F ���v�dm�#"Ol�k2�ʵf
(p� X�5jn%��"O�ؒ$�=�z��Q6hWlq�"O�Uyগ�~��N�	P��P�"O��a�&j�Q���C�	��"O(9c��}P��T�["Rܪ�f"O����(�0p#U)�f`p"O&)p�s���Hā����=g"O�}��+��Ĭ0��J�2'�J�Д"O�A�Ղ�:)�fe)6/^	���i&"Òz$���R~F�y��ӿvMp��"O^`��6u�x�	A��yHܼ(�"O�!oW� ��ͨ�V��L1e"OB��$��xrQ�%
��B��<BQ"O�h�bE*\(6�rK�!+�t"�"OT��ff�����"<R��"OZ��A������+?��{@*O��r�J�%����UmՓN��"�'������G��`���Jȸ�����'C:!���V(Z�[�KI�-�}��' k�/�lYg�8}X�̳�'	|���u˼�'Z�n^�)j�'y.�K���b��F���g-n�(�'��7��������f����'��=Ak��Ap&��l�!=�U!�'�i����F��E4�H+Nab9H�'��@�w�Ͽv����NGB�
H��'�6=PG�=q x���3ib���'?����@=��P���0mf���'UȀL�����M�7 '�Q)�'�ʔ�r�;3h���w���tX
�'���1�JQ3c�����>�.$�	�'�hh�J�V,azd� B��``	�'u*E��˗"���I��4�XR	�'�廀�@*e�Y[�	߆.F����'������q �8@��Ðu܀k	�'Z�b��X�Z-���U��'���Xg�EF*��VA��Ezk�'�8Z4�KB��ԃS��=���@�'ʒ�y�m�b=`�C�j��/�h@{�'F����f�>)��D�!��,�n���'ݰ����8?�	�v��'xܕ�
�'T8�Fk���ک;�F�FZx	�'&�m[w`�V��R�K�~�J���'�$`�FH�`I�Θx�<Ap�'T��e�;"��T!�k��(��'+���I^�RG�Q�J��\� ��'���Q�@��yR��� �*1:	�'��	���+e��R�	������'���̌�sB8�&�@�Z%�!�'��Hw��M8��զM?pu�	�'{�)[�M�7[�!��N�I�H��	�'E� ��ؗEx<��[�4݌ 	�'��%f͟|�<U: '�=��'�~�ځ�WYf �����'?�X��f�4l�f�Zň�,��0�'�K�YL�aP��Ȫ6�Ĕ!�J�R�<ɑD�`?�A�Q'ѡGk��r�UO�<)5)F�huęQ�aŷ׺uهK�q�<ق �),�!q��37��u���b�<��FÁc��U��.�-�
�3検W�<����Ev�L��c�17���h2L~�<�  C�ίS�Z��RfŖB����"O|��6[�ֵ��#jr�"O*�-�90 �ʡ`N�r�<H�"O*�j�c/?p��hU/�`RJ�@"O8|05�B�q��"'n�HK@�� "O``	�@]�#�x��L D��(�"Opdo�wyZe��nN�#G��i
�'+`+U/ 7��J��ָ0����'i�C�Y%J.f��b�J�Z�
Ժ�'����a�JG>����O���@�'"qZ2`QJ�|�`-�8K|0A
�'f��F��Z�񗩆�:~t�'��lq��3�e
 (�D�29�	�'yx�D |.,Y�",��5 �0	�'w������~��R�L�0+�H����O��Eh� @�G$,)C%V�.x�u!�'��jS��D�4�3(�������'@�0Pg޴_�KM>}�U��'-Ш��R-3ƞ�B�e�"ͫ�'j����c��a�G�4�����}͚������d�uOV�*tƛk]�n��T�!��3^����ԆT}�q���q�.���)��@���
"P����O�c���!�0D���T' �;0�f
M��͐�+��8��	�fS`�������d	�<����x� �e^�lm��k��`�ˍ%���L8P��C�I�%���04��t�V쒦�K�r���	�OD�@���=��O�d�"J|�iI��h�5*s"O�@ࡌ�9~,
��e-�7K6���i%��h���%w@�1j�	����R�D=Yw!�
���Cs�ԒqE$�֠�TE�$r� ��	;)�
TKVeZ� ~T�S�m@e�V����O��$�>U�e�N5��a]�s\ĩ��4�hO?7�P	e�:1C6ū���#�/6!��`�h��AD�6��С�;L��|؟��E�O!#Z�����E��c"O
tp +D�L� DC�"_��"O���K�OƲaC�OE~֌� �"O�9#��Gf���P/�����"���G{���BYCr�
'(��C�P��b����	x���@c�Lx#H����T������:D��� ��>�T�c%Y�N׮���ɢ<�	�!�B�qG	�|����҇IY09��IQ~R�U}��x@�O�5����!�y��Q�l��T�r��'� ����P��y̟ �h8��Y�%�0���y2 $��XшI���C�Û�y�`\�Bmxз)W:pqF4�k�9�yR�֎x������h���S��ŵ�y2�@2�\@�s���ٲ��y���9<Q�S7I�>0�0�x�*
>�yb�W�v�:XD�5���É.�y��	0�j1��7��b�� �~��)ڧp-�5���S��ԬΕf |��ȓ}SN)� �Dw�U	!�Z4�݅�	A�'�։�4��Pƅ��P�"�f�J�'_x�S �^ h�#\�
&���'�R��F�;4h�@5��<&i0�'������8��_.����'��ArnOw�t�8�o[!\�^%��'�(u ��N�~F( �A�=I*�OL�=E��>V��h��G� q�0j����yҡ�����@�Olh��q��y�)^~ϒ�㔪�:Bl�pѣ�y
� ����G��7{�Y���r���%�'�ў����݀g����A�^�1+ى*#D� d�ش`m�����Z��ذ%� D�t�U��~��<�س��L	��0D����$��	В��<����B;D�,s��� ��Q�C�
Z�J�B�e9�O��	�/��s!gZ�c�f�jG'&�����<A�Gu\�Yuf��7D ��)�U�'.?�;qA�8S�HR䫘?{�<(�<D�8Bq�L�05����[_BH��f�<D����ή/b`@�C� �;qmz�X�$���Y�3P�۱J��h�$��ZA�� %���D K��>��5qB�V�)హ��"O� ��*�:6YDK�OU����iTў�'�~�\�\�d˴e[�[�G�	*�	��K=D�`��O�7]pLJG�A�?�h�E���y����Oz�Y��C���0�A�^��8 �"O� 
F.K�%��.��mٴ8�S��o^}��'!`)���5�.��elGr��D���hO�U:���i�&t�@��(1Ŋ,v�'��0g�(�s��W�e��T��-���u����I��+��)������Ʉvu:Ekr"O��WÑFP�m�T�P�bD@�"On0X�,T�+�P,����W��"O��S�ʗa��K�L� ڀX���>a�%4��u_�X��$u�@3��؄ȓ��03bىl���M��I�ҙ��?N̩K��t�ÈNJ�U�Ix�����Iw��C���r�I)U�f��!C4D��d�^8D��a����b܀���<y�^��@г�Y��aՇ�#@��ȓq�n83%Z�Z�b�aփH*b��ԅȓC ��Q��ZJ=!��'F�����w�z-�7
�=]�i�hQ�i��ȓ8�P5·0r� �`�̣�\	��w�\A��#�1�.�+�J���t�'��CfgޖA���J`�ʲTrUҍ�D=O�1��E		� ��F�-D�U�7"O2���A�4}d]�W��R6H±��,\OƘ1�����y���,��4��3lO�!{FBnx�%�H�HD.y��
OH7��q��Yq�g�	V��FX�!�A=  ��׫ĔS�V��EO^9d�!��	����S�LL�,ɮ]�ŭ��k��IIx��1�+���v�:�z�^�36J&}��)�ӭ.r�dg��|h������z*��.{�Q��GzҤO�RT2��ǩ�vK�(y�B�I�lR�u��8A܃���D���DQ6�%�t�Ӊl^
8b���B�v�x�"Ox�RWG�<@�� ��ڢg���z��H�Q?�ˤ�K0M�ɰd���(^��8D�hVD�(C}�!S�P�G6$Ġd�4?yB�?�S�O�l�)@H�!/����.��!7z� ���'�,��ƤҹP�xA�]�u�ر�'�W\?�W�0�<�O�谚��?"��mB�!�6�
�'��`��-O�]fh�A� m)$�m޿"�$�=�Ok� 	�FR�%2�q&Z*XC��pS�$D�h0�ҝ:^�! 5�֙8��<jR"D����O3 �����8p��m>}�)��&$���gHEÇ�Z��C�ɛE�{��ѪH	:ձ��D M�D{������B����" Ã�]Y ���(D�@!��70�uC�e�4\s(�F/(��ē��'f���Cǧy�9��ݮQ�:���HO� @�YTa�}oHłv��:^#Z�X��	F8�|�uƒ�A�<��@U.�7;D��ҁ�	�s�u�G^�;g򅊳a<D���_������:9����5�IW؞P�B�5�����N�.s�@(9D�|�ԩH ޸�Zseطuz�h--��p<�\7n� F+�"R�*A(2��A�<i$�U�)��a��QW�n$�d�ɦ%��sGP)Y!ÅDE8�����׾@�ȓ%iP����W,A\��!�Փu���ȓS��s@5/a`�WǤUO�݇ȓ��D��n� � �(�c��l{�'�Ԙ�QcA*��H��\�eq(|���'���d��^F��GK#3Et{�'�������<I�l{�A+2�d�
�' �q��� L�@t�_i���v�=D�i�M�i"�	]:w:pfa<D�8�T/�mǌU;gg {!�)$�8D���b�f[�Ă��M L�f7D����ޥ?� d����c&�p���"D��W�|gP��#�\�"��Q���$T��!�-��}�.����v�P"O��Ӧ �3���&�:�H"O����
1��ke���<��0"O��@�F�
/ taq� G����N�t�<��o?�*�Ӱ�>�Z�T�X�<����!c�ؑ7쀸pmL� ��P�<qm�H�bI�'����^K�<q��O�YZ<1�I� X�R}�E�SQ�<Q"Ky��\�׀A�q3���B��J�<a�"��@QL�9�b[�T�V��chC�<�7=J���+ O����ӧ*B�<aTeHD)�,x"	��W=H	�%�c�<I�ѣ6����g��"D1~�:"�[�<���F�|m��kCG
R; hR�M�]�<9�� �4#0���B�M��B�<����
c�����o����5���L�<� lB�dT���,�F z%g	|�<iS�\'�d�S���#Zf�ٔ�c�<�����\��Y&��k�By�íS_�<Q�K��S�"����� )Ȗ�*3/ _�<ae*J�±�è����څHIs�<IeN�+8��qy��y6ƅJ͊r�<	���IB�C���(��TB���q�<���63�~ݰ��*��I�Oo�<a#Cڃ)�f ��DX�lV(�ѕjp�<���-<��M�,R��8�j�!p�<�֧��;����J�I��uIP�<�pM� {����T�b���SU�<�L	8����Ɔ�1��*���S�<Y�C��z,Y���7<�x��S�<���� �(y��J�ɜA0��u�<��EK�mF�|��l�1kNq��v�<� _'�-c�
�B�Lx�`�k�<�r���*���E��<̮h���d�<���!L���3�.`\�9A� Yg�<�T툕6V�E @�	�z���P��\�<��ӈdh��r�A�;@.���/T�<�jߗ4��]s��A2D-Z�Q�P�<9��`:�ճ���y���20"�K�<�a��H�K�B����a�Q6$B�ɌA���2CΆJU�TKt�G5��C䉌mV\�ӕ��T���q�/��L�B�ɗ����FɩIܙ���/��B�)� �[�m"��]�"c�%LA"OJ���L��/������F�|p�
d"O�l*�瀿K�$�w"��~i<Jg"O�{S킶O	�LS�ġ%�޴�#"O���E�������X�O��ȓ�"O.A���E4�f`���޶{�8��"OdDx�iΣ}4� ��ܕ=��"�"O*�0���, }v��$�M_�ʘ�d"O�����/���Q�֧%)�"O�]K�-�[=���UC[d�Xe8E"O� [�LF(p�����8	���"O�
" �,Z���e@�%S����R"O�2@�g��ЀE�B�P
�"On���P����`ƅQ�B��J1"O��ώ*�j(���L�O� ��g"O�`�E�W�2�Խ��b�d��"Ob�j���$/���ěG�X��"OuHF�:�$������HQ"OZ}��N;g��+�)O��X�t"OP�;H¶w	�E`��ƃ��H��"OF�K�C H�����҂����c"Ol�	���z �]飤��dq�A�"OH�,��l��L�A�-��"�"O�����]Eƅ˖g/Li\�S$�D�U���$Y e"�=dTp��2C݈S�Ab�"O��� �G�s�-9�"�	�P&߻ qO X��Y�lX� D����C�A';��aB(D�;��_@v�i@���9n��CM�1I�iP�8�O0`a���/�j���_�'���'B>E��
�F~��'sݰ8*UIȌ���v�\��y��@	d."���Ss�#F(���'B�9{4�F>���9b)N���L��H��N=D����֭[��x�u�E[�`8y�g]�-un�4���<���\�*��]�V&J�3�����B�u�<I�h	�3��xfGP[�����'���%�1F�]��\@"��r�F�`�C� ���d�!D����!HTy
�Ѥ�'Q���;D��)���}��8j񡝑S%$��V"D�� @�; �	
t��'��!�#�"D�� �'�?ٌA� Kԁ)(�]9�b7D�� �j]�p�) 
�W���*g�2D�Py�G����!Y�ԲN�h�b 1D� �! ҏo�p�R� ��U!N�r`,D����.](]�
A��	1 �VJ&D��:���>2_质�e̓7�P���$!D�(¡�g'�4B�\K��I�l+D�xCE.��`6�x��<P����N#D�8 ��Q�%{���T'z���j�,D����A&�,��g�23b��J��1D�*�JY,$�L9SaJ�B�x��)D�&_3��e@OO�mQz	�2D��@�c����6Ɍ?IdR;60D��h&EֈE����K��nE�'�.D��r��p����@��ұ��*,D�DBeԛ�K�C�|ݰ�-��JS��D�?P��u��J�`psfđ��OV� ��&�Cr��b2	;��M2^^)@&"O�9rc���
%����&J<��I�1O��� �8Oo��O?1@��C�`�l����1D:u�1�!D�����!0�����gD��D5S���<yǋ��8�;�l),OL�R� ��a!��ց��6�D�²�'�L����/
,rs�8M�)�v�Ģ�HZV+@bH<I��ظp�2p��ń{�z$�"�q�'��x��ݡ	��t�~Z��R$[�n�E��Q瘘Qu"Zz�<� R$�����{���F�V}P����'@���-l�d�O4��eO�>\�1�4�X��D�b(y�C�/K�`�r�&lOr��U�ԬSM�ݨ��[��4�ĦQ4;��A �(���6�&��q�R^�P	˓S���#��΍.�@-p��	�<���<y���&=���i�<h��gJ:���&A�Hx��`h7n�����F�)<�<��$�.��x2�9y��D9��95��IU/Sr6��W�����[SύU�>�9_���w������{�܀�;0�f�/�t�y�^�,���t�xh<�����z�h�'��`�S�Hj@�i��Q��q:��H�;��9�� ���J��^&��p%�8���_�-G8tbu�\k_P�rd�<,O�x��J8;ޮ��e(ڸetr�S��OgM2�Hݭ$V�B���V�|���'u���bB�o��x�Qi�[���B�훟L�̑uN!�$7=�>-س� 
;:�� ���_B�U�3i >��5� ���$��0)P:d�WjE�|� "O*Tq��
n���j�q��5�×b+��F`X�#�i`���[�2d!vBQJ�d�v�ϻv��v�N�hb�`�>2���ZLR��}lT�R�� ��9B���$�ڨч�-/�00��'��(�-x`L8��}�fJ@�R�q5ݚ	�R�6���p<AF��wc2�*���� �����0xô@�i�:4���܏/�A`�� 5J����3��=aNT���P�Dn5n��1�
E_��h��i3Z�L��.նh �H��.�7j�Qъş��'����h!gַ"8�es��`�<���- �&����ǟ3�"=�
��mP�jP��]�r�	3��A��l���Dm����e�\��w8a�! :�!���W]���0�'�6Ԩuf�������O,W�5�5��Zdj��^<^���2ŏP2]�Ƙ�f����<I�):h䈁��R%\'$Ls�	_8��36�@�I�b�Ȁ� $t�`b�N��"͒BV�j���A��]�U���X�Ă3GX�P`p��5%�26��A��4�d�,�$�1���)≁�i��&ġ��O�&Y�6n��Tgzh��W@�bA 
�'٠���cV,h<���n����
_6v���>Њ���@8����@������g��L�ԪO� GY�Ɠ<@8�0(<���oɥR뀠�0�%�����/��P"ӓ �	�Bݷr�rL���Ѫlut�牷s�t\���+np~���G�͸@�D�G����eƪ�~����Z ��?:>�� ��. �1�<�0��!�!�A�����|*r� �5�0p���XLzV��j�<Q&Έ�Y�zMaU�S�4d�	��
�$d�$�e�WW�8�YS6O�DF��O�$d�?4h
�"�DK��3�"O"�Hү϶:+���Չ����3O�h��Q0.�T� �i��p<1gi�/sH��F�":� �qw)�H��XZf\$�4 �3�E�����D,,w^x�z6�C�;R!�DX"t����Ɠk����D՗q0Q�,b7I�wp$���I�0v�g��.(�����@y-!���.�tj�CK����'�7R��*$zh�D�N=��)�' ;��)H< 4�#��F�,#�E��� �@��P6p�n�!�GјH0�I�	[a�H�q
��� �S��d��u�)it��>4b��IT�M :�~2�F�O���������Y�7��̈��S]��� @��
�Mq����3p���x�<�b��0X��59EeP!-�Qr��9"��$�U�ޒQQ
	��b�&8��� �����_ ���s`�!��Gx"�S?t`	���ED�OHX��$ 	=�܍��_��ԝh�'H� ���.�2���9!&�l2��Ӽ1�TIgއbR�i��LE7.���3���w��e �<i���O����AJ\�"B�*V8z�%AXcF-@�d�
  ����#e\���'�<��*&b��L2�-֫pը ���-��Ar�O&F�n����F0N��)��i9�ՒnD�Z�� �S���VAP�^9����lN�=:s�P���(��|ܾJ:0)�p*X()����ʏO�8�j��K4z<N7�]�ݸ�#��	
c�M �ŀE��O�:��+$"�x�4#|�V��)4��"�O�?:�I���gܓG�(��Ф�?�@����I˻Ga�JV!�)*��Eҡ�R���+�Ɵ�b��b]�F��'W�����C�D�A�#��={24s�K6�`��<��l5�gy⊈>7�rѩ���d�z�cCU��?a���/q��h8�0=��l?Z�j!��K8��M�Ä�ѦI���fPx9��ɇ9��Q��dUoϠ�B�6�|��`��&%�
ɀt����=ф�!�*��'���� �y�4�b�܍Dґ����:p�\u ���&��m�~2�s@�ÔeݫQ��Ah �`�<�c�����H���iP1�I!��)"��̙���>E��3��%Af/C?\�옑�)ȳYc(Ն�S�? ��G�T�H�.e �FH���3�T� ��1)\�9F�'�F��MH�9EbU�B�0Ln4L)�6��c���'v1����.�}"�����(-F![G��>�F��G��44��0�&�P3��R��%:�μF|���#�$:�@�vܧQ&p�E���[��ɺt �������6�Op䩶��Cx,�Q�ʊ�.~8Rd=O��	$G3��\�J��OQ��@�Q�<���4k��*�(���%`�I�<y�W$�:���X-5O�YxŲ��'r� ��8�XlK N	���'(��ӡzs�@w�!$uh@"/[jt �����8� ɣݯ1���{�!��a_��k��]%Nt��*��?tqOz�E���2n���0�N�"�6��@�HIn,G}��߸	&�49��I
�{E
��sEJnm��A�\���p��9B
�ba�я�>���M��D�'�h���f�S��$�'Xw����NTq$�<�>\1��=$!�Ċ�7:����ʹ#��]*��;�!��S�t�PV���m�H)����@�!�+E�p���c���p��.e�!�$��3�N�Z,Ԓ[��pF���k�!�ւ2�F�2D�
	_�:�s�%�%Ee!�E�C�ΰ��E�C��8&"��'X!�W�a!RU���!Z�6@�q ��U�!�_
y4mq�F�k�l:AnW�s�!���=Mp�j$�m��C.���!��@�;�H��"m
�^U�¤�
b�!�d�6�AS��G0jD���"U!�DϢ=0���i��1/l�9��(;a!�dK>#�xh�k81�X�`$кj�!�FZ�*	h�����FD��s�!��E!1shi*g��>1���zT�؃!���3�.a֧�5Q�<��!߳+�!�䜭UV$�b�l�'[,���<O!��|� �Q�F6l0�\~�!�$�-��85+ ��ё�<t�!�D��p嫑���Y����ݎl�!��;�����H�S��ѳJ;!�$KIP��a	9�\jh>�!��X�MD���F��J���Q���k�!�Ď�G�j�tiY�u�@�0Ak�x�!�D�Q��d�c؎B�ȣt�L�`!���0������D���Cd�W~!�֧{MX�X0�B._��P��U!�$��2��҇���"k�Q�PB�0Y!�$U�w�*ϟ{K��a�B��&8!���1ORTK�<&,�{��?>!�DI&=�
e8��'kx��9A��/"!�d�e:�\�G�	&D�8�[Uʑ�!�d�����"�n���(�GX0L�!�$	<�Tp��!ٜ=��c%�3[�!�C["��Su@�]#>�qa� !�Dɨ)9l5��NA�O�b}�6�	�^�!�$O%,���!D\A������&De!���h� �8'���bTpR��'r!��Y�P]�YI�ߔK����U�#7I!�dϮ'`p0["O�[��l���}.!�dݟk@�U0��Z�P����s9!�$�N�Q�g'@0Nchez8�!���f���٫PP	�O��A�!�ȫK�^���A�(E���p%M$5�!�dK�}f�,�
�_K^��,ݓV�!�Y&>F�#Q�Ǻ75����8 �!�DG�w�
9���$ìeI��!�!�$U�$fЕ��j
�Y��i�V� x�!�Ě�,er�G��n�ޱ�v�ڼ}g!��M�f�p�1 �J,]�\��C\^�!�� <Q@ӀӾhP�i:#�H�d$���"OF�
���
[:��iS�[�5��"O���D� Д��cNF�<	�"OJL��eY�xh�`a�Ti��#�"O
�K����ƁR��������"O��:���_����ԢĸA�4�+�"O��:�% -m#���1@��`���"7"O� ���W�n�|�����4A�z�!�"OȨѶa���꤂ ���LL��"Oz�`�!�-n��;@위n��(�7"Orm��G�!v���0���Y����"OBРѯ۔S<�XSu�؍b�z�"O�j�D�z��!��
�7R����"O���e��M�" X1�P{�Z Zb"O�=�D��t('�Z`0 �"O��y��R 0�v�R�7P�1;���y�<!�Ĥd	��G���,�PI�WJ{�<�e�_�RX�-���sO��s�@�u�<yQ���p��%��Z�B��n�<9�oH�.�XB�7]�\����h�<93a�&z
 ��.�0g�m��a�H�<�$��3{捩V�)j����B�o�<���<y�2Yk$�ɧL���N�<D�F�*0tYb�޸N��*�,�a�<qӯ��y���rVHƻi��.t^ �ȓ��o^pڤ0"E�$|���ȓ%�����++-�������)�ȓk1Ҥ���Μ?ֈň��ݥA (��ȓTm[B� YhV@�Ԅۦ|s(���r	���O��*YV٩rh��O�r݅�WƢ��F��$����kŭVQ���!8^��*υD6�+E�]kD� ��v�<�*�oNR�����x�=��0I�֭ȄC
h�S�EQ@�ĄȓoXx�ʔE�M:�ӡ��{�8��ȓ.�Vp'攣N����	jKn���m1�i��o�O�a�B��bڠ��[@4sP*ȋ����	Mɇ�	҈��`MB�kEN�����}�ȓ4���]�Dy�bd�"��\��47d �`��{9r�P���	�-��k�XM"nE� ���,ޗr)�Ԅ�j"6��w!S�@l��ʀ��d�� ��ts�,!'FZ�%j֤2���!��ȓA�jp�������C/-�ņ�s�fq��_,k2:X�T��J֊���:*8Q%$)N,I�!�ۑKP�5�ȓixs�����Yh6hD^:p<�ȓ:u1W �'$�᳴%�&�
T�ȓ4�:(B��M�+#�6|�ȓ������(��A��h��=I���ȓk�ܪG���k�r�����r�ΰ�ȓ��U�����1|J�� %��0�h��͸(Y���"��ey�Ǒ�u��m��n��"�P!������K����.��Q�4|Jdar.�3TH�@�ȓe�r�R*bRT��g�˷ �p�ȓs7yz�H8R^z�BR�[֮��ȓ~'��aQ�I�lD��+����]֞�[ H�4���s��mK$�G}r�ɼ��F��A��xa�d� I@��jį��y����Y;ABT*)�@AS3ʏ2�y�O�4!N��B�|���ǔ Qށ��c\ �Y��6vi!��A�ZgdK#�_�f3.=9��_H�ɐ(�р�$@A/ay
� �9�	�8��	A@C%r�}��'�e�f�m�����;Ddxp��Dk�)Q��QH<مf�S�^����59���B
�t�'�|��[+�J���I�|�^�#Ql�f'0H�F���!�$�C��b��[��A��*�t��I� S$������T��=E|�"u2�C��Z)]|~���Z۪�g��25=<���g��I&�-��c���A!�:AY"	�f�����8��5OE6+]�ȅ�ɯx.�M���1Q�Ԓc�R�"�قUZ�����cL,��xAļc�rq#ҀC�i�|h`��
���i�x`p�)�;0J��ʗ� :b?M�s�ͩ$��%�gg[�� )4�-D��ғ� �0!��ݹ`�
��˕*>!�[�S2?ڙ��@0,�Vc?O��	&�>�h��!�_3���C
O��0Ñ8p�	��H�a��L�eKD5��1�ǞŐ\!�N4�0=��脾y���"
(NN�#��b8����'*%�(�GnI1	��=nZ�b/��&k������	\�[�
��#�dq�)ʭzU*��J�0AZ���O�@(���g��<᥄�-G2#}�/�2r2��6FT
1D��& ^s�<Y����Pt	�ҭ�X���J�@�$��nD�c� �z ,�)<l����V|&�$�w��-@'�;�~����)Za{R�S=�[G�%늕���
�v��+]�n��-AU�ƫ,����s�؝��U԰��(�=Wj��4�\-��U�>9'��>~Zy�掟�
�L�)c�S.w�<ܓwa���\�G�-X�I��Z�g��AC!"O��2Pn��:������0�nm[Sd���İC�J_ԅ2�*74E��"@��м��牃)�:�pM^�j (B3	u�<a�Q�[�8cEo�@�b"X4t�-�u+@�S��I�O��)#�Q�;Fz���ؓP��L�"��ƼI� ���a{ �2b
�i2��&��i�@���n%#��~4�������ɘ�ֲ�>fhț	�b:GiI�,���i�p��~6� F,5�>�Y��)2��B���ю�@�8D�4{V�нu�~�(��̪U�D=j��3f��{��'�)��<�'C?=9�ٚ$MT�2I�E�j�<��8J.K��]�?���!2��B�<)�`�{OjTk�ƙ�h���]x�<!���=��	ie��J��t�#&�c�<�'��l��H���dRi�u�<���+;�Jm�����0�4�PD�Z�<!�Y�#�du0S�ܱ;��ҥ�Wy̭r�B��=E��₡D�N���g�x��'# �y"f�-����1&�R�k�Ώ	�ēbN6��n��p<�r��6T�٪�$��1�NW���Ö�
 �>Q�A�O���d�Hl�l�r*S4E!��i�Pt�����9�I���Q���	ĕt<�!����V\�p�CƗ,��y��f�
�!��J�LJ���k��@i�"�2�����(m���
*��)�'$,4��n��a0�YZM&����ȓ:C�\c����5O�q��G�V L�O5ȼ=[�ަ/v�`�@t�����`a��1�뉄W�dP�P=��~r/�7#"��I��P/]�~f�@��h#w��Ay��uO�b����$Vl��i�o���"PF�m<I�Ua;q�Bu�w�I- c� �p��ZJ�+�ɔ{��خ�0���U���L8`� � Dx�C��d\�W�HV�Ot�cDd[�H4(ъ��G@����'�>Q�1i��W:2�UN:?�)��S3j�4�P���!��\�`-�nr�=�&�C�v���p,�<)���O�is��y��X`�������ܒ0;pp˷j�Fj��	�����'Q04�󥈞H3����i�2$�iA��9[��ٔc?+�J<S��$�O�|�U�X �����g�)9<�{ub[[Ѐ�a2�K�sȈ����̩;$���څXՄ��W��,GTm[���#��A�-:\O�SH�4yH@����J0r$��r���r�F_�LlJU3s��(il�� �ћ�#|�l8���lTL�#�.�@�'��17-�>es̩���i:~���r�l�#}��X�ΐd�켳w�-qƂ �P�F��'ƌ��E��|86� �:}��K,��]#p�C�<���1�gy�H͊\�T�`��qm���
 �?�%�Us@��IW����0=��g�'Y.t�F�ڲj�N�Q� ٦��D��L��@KF�	2k�B�i��Ș8x�|j6
ם.�.����v樹�!��=���N4U2򚧀 ��q�R��%f��j�ɣ��I:x\0��C�$ +�C��dh���"�BBЧP^�8����y��|��A��M+��2(Rj|ҙ��
]G�n���"�P}���']d� ��@�?u�]�Ӂ/��'�^(kTC�:���
҄ h",{�Opt���	�TH�N����(�)j8x8�Qe�>eH����	�&|�@��̔2]D�9�cß=���&�ơ}Q�T�
O�=�����d���#o[�*J�c%�;e�@d�VL�3Uaq�bxcC��_���hG�Pj!�"Ov|IA��{���"qg��j�Uka?O>-��		)}���N�"~r�/ϋjZ*����$"ry(&(�y�<��ВKw(�[ԅ��|���#F�\~�(�-�dE�'�^8��U��<^v���"!j��Ҷ�-�O^a�-Y���!ŋ
\����&�~��yrCj��PxBɔ�`�Z�b�i�-���'ߤ��ONQ)��+��b?�cw�@dEଳ���oxlh�,D�H���V�[�@`)�ƛ9�Nta�>�%B˱'2��"}�fa�7FN�"��ɒYp�;�'g��G�$B$��0�C�R��z�'�Ec�mp���(���?oD�@�'!쵊a�#_�U��2���'ܐAK�!1��`S�7>��',�18��ȍR4�+���1U�\�	�'���5��1àti�'��^hX�y
�'�4LQ6$Q�^@l (��f6t�)	�'�Q6 |W:q9���U�
|#�'�\�wݝX��pw��Aj�d��'�R�`!�/��Zv�.;�0�1�'o���Ft�hz�+3�����'��	
R�*H�5�vL��?��,��'�LD�aE� �8��(�
Q�
�'�t�i���#�t;EA	�0�p�
�'�����k�- L�oԼz���Z	�'��T�&cJ�\{�̲�;m��,��+`��q���&-�Q=k4XԆ�NT�����X�u6��s�M^=F�ą�`(0�K2% =^l ;�A�d"a�ȓ�4������U'H>i��q��w��}� �׹m|��pX�|�ȓ7���1�k�-���;�%��h`�ȓc&�h��#R�,e$�[��W#\����7��|��`�Hs,�A"M��~ }��g�4!��8����&+G	G/�,��7D�����JP��@��hҐ=��0�6��0
F,
Pp�unU�
Op��LV�h�ӊ��)W�Ż�(�5�^�ȓ'ht�W,�Z�����5f��ȓ�tA��흊]��Bd'��5�M��"��9x�/[-���Z�NS�j�x�����qW�]0O�|j�g�Q����}^��ծ��(s*A���S}&���ȓi6���)�p8`f��a�t��ȓV{z|��_�y�X���o͵\��d�ȓ���d��>i�̜kwnR�=��n�`��Z�^�����U��Q�ȓJ���C��p�D]SB���m�ȓN��K�Jؓ( CUs m��:��<����&T<)�Ǝ$=H���ȓ8���n��]�����m��8a�M��l����Ġl�\@��־�p]��~w
3��ǃ}k}B�+�7/ 4��ȓ'V�U�׼m���g�)>/��sr@�Ydx����ʀY[V{���	T	���9|���{R�\>�0|Ҁ�߳uS�%`�:�~�ك(Pe�ɔ:�|�ѓe>� ���ɼ2�P��"��kG�9gX� JA�ʌ�%��|:@	�'B���"!��h�z@��	ǟx*�k��S�H$��~����?d6�, �nX�8��$b�`���Kv��B��N>� �+M�]s����ʞ�wa�x$`G� �������=r&OGt���݄.�`e[D"S�>���e��A%b(6E%0�3�^�>[T}D�Of�+Ů���Y����$݂l	�A�;R�Ţ�u;��	@>ɸ�*N.b�*�K��r;��G�����*v��>�~�-X�B�a�T�M	b��}A.�X�]
֥�,Ddܐ(	��Ċ��0.�f%�ᓓ�䄡�BQ�@M9UiR���F?Y!�PRLQ�T�nq��M�OT��!2q�"�I1 ��q҃�B \+*�+����\�=�,ҧ���1Z&
�E�t���F�n���cX#e�UQ�o�km6�S>-�2��fC��s�5)�4�Y�Ǉ�("�=a&��y�F������'
�`��J<{�س�OO�	����P�@V�D�R��y�g�)���f�h��v�ܥ! �B�	5y�KB<��DS���S��OP�U�,\�b�hiR��<��V��B�)ҧv��`�JxTpj�L�c��5�ȓc���)D$p	�YgW�^0<��bnv�[�!o�T��i��v���ȓs���GR�����C��H�%�ȓ�Z�QG�Qt0���#O�g2�-��o� U�T�8VXm�@T��A�ȓsv>��c�U���!��
�?+�(���{"\X��k�0�XĲO_%�C䉝z�L�-9f28L25L+K�B�I�e����g_�_�&��"�:C�I�"�% ����/�X͠C@�wC�ɠ<f����"\F��Ǖ�Y��B䉈D����
��-<J�8��G0bo�B�Ɋ	B�A �l��?92�85AF�r&BC䉔��R���P�jq��ʄ�]�B�IYҴ����N�@���&�2 PnB�? �SR�??}�d����;mjB��-�6�P�A�d-�U�W�U :`B�	1�`��i��:�ĐB$@��C�I�u�Ё�#dF)GL�t�#m^2
#�C�I�>6�ܻ��C5<�h�+#?(��C�a���Z'�A;t�^Ȳ4(!��C��8X� YC��]gV�91�
.uJ�C�	mV���#М=�B�xk�k�C�	�<�ڑ"B�L4]Fx�9f��VxC�	V�Z���ݘ`g�Њ��f�6C�ɾ�ԡר�/�:y����v�C�I�r\�c'�]\F�� ���d��C�	��Y#M͖]g�th���1�ZC�ɮq7F�#�߮Uͤ�W��Za�C�	\Q|!�f�Z��0:�T	J"TC�	*g�.��E5Z�<a'BN��LC䉬�Xp���B�J�A�� �l�C�	zf�#��]�B�R�` ��B�ɚɸ53�D֍8d��q�y�lC�I
_Iz'�N�C�&d�Gl�,eBC�I�7kF[iӺ}~�2�ܔg�C�I��X� mI<n�}Q��k��B�	�)܈4!���T���W�٠x�:C�	>�`�b&Ʒ)�I���}'C�	�R�hy0Q�Ͻ����
���C�	�>T�1�'3\n-�b�"N)�C��+�d�VkA�r&��դ�)�hC�ɫ9�����G�<��Iy"��DzB�	=|�D�y�(�c)��S���>
�B�I�uph���6]�VQ��[�C�-8&*�q3N�@�P���ք�xC�	&�B`*�DԨ/PD���?pRC�I:~K
�[�!C�8��4�)4��B�)� 4�J�D�U��ڃn!F��"O����Q�ecٲ��͈
�쪤"O��֠��\� 3��ލ����"O����K��ݣF��4<��PC"O�9�5OD�mE,� �"&�f��Q"O�y�2+ 
�5c4(\�X�hz�"O��Y��U�qbTl,X]("O�=s���4�$
�*B*��2"O��r�C&s����p����"O(���	.^��T@T����R "Ol���̙����KwB�qp��A�"O"e�4��ꬺ#Q,l*=�$"O����!&g`M����Xh�i�"O*e�EB�f��@�5Ɓ�\T��j�"O�tx$0H�!��Ge��b�"O
� QG�`}�7�����'$�H��� T�3'��=vA�u 
�'{4Ѡ6+I"%$`a���R�q�2s	�'��5�qb��SDq�픡f���	�'��`#�)~T����'	`X�y�'}��tO�;{>R���݂)�~!a�'�=S$�69����ddL�$ɺA�	�'L�ˣdY�L�(�t��P&R��'�`8y"��#��X��K��l�K�'b�-��ā��M�d�T�_�t��'}`�j�π#�p����O�>dD��'ydt�#f�y	&y��Q�Ƹ��'G.h0S�G�F)tL�"Sٔ��'�Ni��GU"h�b�5�$�)�'�F@EA �<.�|�6�Q�0���'9�H���=-�hzv���1�h��'$����Xr	�uڀGD�3�e+�'_�0;�C�5EZ���Ѡ8s��C�'h�����$Q�oD�"�!)�'XA��q��s�H��.�H=k�'fp��J�7\:�s�ݮZ�~,��'�z�b��ިr��!�)��P�BXQ	�'�&��QD�1M�ք�b�I�J�]s�'��1�'Յ->���H*5�5{�',Y3��L�}�B\�v�$+[�)��'f�(��>�Ru�Z%�\���'� $���\2�����3g�0K�'���$�@��bP ��$b
k�<�"�fi��`�*�>�3��[A�<�ǭ3D]��Zw��*�<��v�\b�<��`@3f��W�P�4^�A��Z�<�W Z��p$�8�X����x��B�s�|iYb\�00� d��0�B�ɵ3r��
�!*�*Ð�Iy��C�3�$�(E���9k�+8<�B� 3/�����*)���Ue�.5�2B䉖\�]�Q��'�ޔ)�����FB�	�]�搊���4�b��"f��~8B�)M\0y{B ��"Ո��(��QM�B䉬`���q�4`��B %�/J\PC��&��b0nI�UZ���ou�@C��D�L�v��he��� ���.C�	[>-9��j�����g�k�\C�	�o��;�"�4;t�1��Aԙm��B�ən�f1��S��aك!��Z�C��)^���#������nC�	/B��0f�G0Z�0D��{|C�I�m��@3��=k'$��q�
\C�I�1h�J�O�:}T)�Ȝ�q�DC�)� �	�Bk�&[p�֨�W԰���"O�l�Ջ���֘h��%vEC�"O2�`F�� 0]B�F!ilt�0�"OL�8���(e��0B%I�nb�`Z@"Oha1��o��ðMU2K��"Oƭ
�Mͣ&`0�W�27���u"O�;Ud\�IV�$@׊�0;�<P"O�A��	�@�I�u ہ>8�2�"O L�&	���J�ϋ/Y�ڔ��"O�|���Z���3OK�X����d"OR��D
G-�I�w��%�<�i�"Ol�0u皦S7L�Q0���"�r�U"O��k�g̯-Ւ(˝Wg���"O��A&�O�X�������ɷ"O���ծ�2IJ�)�I�FX��3"O��Q0�V5B�b4��VFH���"O�I��
���T�ҖJt�v�0�"O�!k�$�:[I��c�<���C0"O�Z��D+,��q�ݚ(ܤs�"On�It� %�p1X�V.%���
�"OBթ�T�	n�!��DH�@̊w"OD���$V���� M*�"�"O�-˥���}���Yh=�"O���)RZ�۰%�;F���a"O&�8��~T�HR$��yX���"O@�r�T��@�[eiO)��"O��I���㖈]yt��[�"O�P0�a
2  �r��Y����%"O�D+��γQ�4��pg��7�B�2p"O��h��M�\��k�F�=m��)�T"OT��W��*�Dqj��žu�$�A"O��iW�-:dd1(�E�Y ���"OT�1@�	�>`�E���HZ	�u"O~���Ƃ�p*Dl�@9_n� �"O¤�Ձ�SS*IcG �%r�LSr"O``�6�]�R���k	CXePf"O~��m8�ڨ��E �'�ű�"O����B��)�,H���~���"Oj(xc�B�[��׎$�JW"O|m�2%â�u�fO�� �:5"O&���MW	D��d��M�@DI:�"O�!y��K>VM84�ڝA@��"OLXy�
�g�,��[�a�"OBtsf$��<+���|*���"OP��T$�;а1@ƃ�?�24"ODz"�
a���7�ɘ:Ҳ�:Q"O�X��"��rIKAKݛkts�"O�t��.�b�"�iV>fT�DK0"O8qY�^0��IA�Ǘ7�5h"O�E��U6i_z�0T�2`Ȧ%�1"O�mа�N��[3 Ū""�����8D��c�\&Byr�[��t��	��;D����JS*k���0`�y倅{��9D�P�f��vU�\�G&+N�ڠC2D��;�L��qG���j{�l`�%/D�p��L"Z���/�*U՚us�2D��@6�A�K�6`8POK3y@Ѓƌ3D��cc�!�:�*�䕹~j�Q )1D���%�ݹ@�fe��<�!�,D�`Є%Im9�D�" �m5|���=D���$]R�!+�)O�
"^Xr�a6D�8�U���H��u��7�x��2D��`Z3p��W~G�)���.D�y�$�>8����%X��E"D�� м�k��W���i�h��)��"O.rpa)Lߞ��ҩj��:�"O�5zt�u�Q���z�R�"OJ�($�rV�����"�:��4"O0|j��R���p�L�$��P"O~��nR[��i[��p61{�"O�T���z��`�֧e�leZ�"Ob1��.�$]�"��0�W�����"O>��&i�7I[
t����"O����%�9
$�ؒ�'�)B'dU��"O��C�E��Y��q����)>�E"O�]�5�C5 _��2��rT=��"O`��N\?3�|(e��s~��:�"OE���um��y�=[ц-�G"O������T��(�ܧ1�"M�"O�x1bei��pѩ
�A�p�"O�����WK�5[�'�S5|ܨ�"O�����C�V���K~;n@:�"O�%b�Hʃ�&1R�E
%#/$Ti�"OLA��$��b`���g���"O�裓��)%ܭ�rg�,5�٤"OH�U���[P��QD��u �	!�"O�91��o����bŞo�l�w"O���    ��   �  $  m  �  *  �2  9  #@  gF  �L  �R  1Y  r_  �e  l  Wr  �x    f�  ��  ��  <�  �  ��  �  G�  ��  E�  }�  �  ��  �  b�  ��  )�  o�  O�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#����$$�S�FL�#���<�R@�S���L��B�)�  IÉf�4k�@�3l�Q�3"O� [P�GQ�šQ`�e4ݳ�"OlkQ��?UD�J�%\ lVh*�"O5�Q �$��<f�8F[d��"OP���$*�(m�Q��=[T �+a"O�Icw��#&��9!�`�.F�EJ�"O����Wc"p:D�ϳ8*�5� "O4`1SIL�x�!8&Y< ��v"Ou�a)͋-^8y&m�=cX��"Oj.��P�G�u�h�BT�T>z� ��jD�qɖ#��M���ib� �<ȅ�ɯ��'L���E(Ϸ(�*�����?0��=��'���r!G.x[�i	$̃ ���r	�'Ǫ���!���X�d���v���'hI�P)D
ZZ-���ߦ|L xj	�'j���5%ɽMd�(��[	 &)C�'Wf9;����3a�8vϒ!��'��q#W�r�T�����g !�
�'��}��ҿ�m9�\�p��
�'
|{b��k��|3�>^=j�
�'�x�dg�-^��d�ǛL>��1�'	��!�+*�l� J�@ ���'
��F#�"��88���,m��;�'�v<�0��(5��u(  G-mp�%j�'� 	��K
k�U��H(l�> H�'�X��t�P�.�9��y	�'V6�[e��O�&�x�L�\�����';L(�h>z���Cbh]�Mx����'��-�&�;+�*	�@�D�5ŘU��'=�dC我oĆ<�wA�>:��+�'���&�d@@8G@�;,j�P8�'�ιS呥
ݨ��3�,Î���'b̂���z�r�P��*!Ш���'6�(�JH�ÞA���)�d��'���F�W�uoֹ�u-�r$
�'�ՈÏ�=Y�Z�e�[�:�������@i`�ل:'x�2C��#�y���>y�4i�@a��-���a'܋�y��D�',�i�pD�0,��Ta6�0�yB+� #xj�B�)<!nu�#�*�y"� W���4���������y�K�ZVv��U�׀}�L�j�bݳ�y� �QX��A��{�4I��y��/S�,c���.��@���y�b��΀�ꡋB,i�|�9�ɗ��y�#�!7)���X$��O-.؆�wv�$q&`��_Ȋ<Z"n��9�ȓDR��JW�R�a��7fA�Y>�h�ȓ#��i¥�F�l�q�ƴJj����<q�F�є�r�y�3a"���R6� �-����)#�"E#��0D�Lb��0z���qc�1_����$�-D���&�A�3�$傦�?D@Q �*D�H�@���v�.h��	#;.�f�(D�t#5NW���F1-B�Y*U)%D�\j ��6Ҟ�X�)���[!j7D�P&������l�3zA (`!$)D�<J��:.j��߹<��iSd�'D�l���?���"n�T�ru/!D�8��"(r���ڂK�*Z��8��>D���GJ��o}ֱ�*X�nV��ũ;D�|ɔ�S���X�G�Y5g.�Y�k6D�����Gތ��g�����K3D��pQ��	C��y��(g�ֹ���0D�� Zt��ʜ+�P���f,@9t�X"OLՐ�ƕ�
��=�6%Y"ր��"O��z'�12���k�D[28�Y�"O<d�%'Q�o��%h�C)�� �"OX�"�gPb� ����v�h�%�'"�',��'%�'Y�'���':4����iI�`Xφa�f�'?R�'��'��'��'���'1�`�M���`=�'����B���'�b�'�b�'�B�'���'�2�'�����D-G�ꉫ�
�[������'�"�'��'~B�'���'�2�'�±��oC�YZ2�(��k�r4���'�r�'���'h�',��'�R�'�6騐j˥D�V�D�>�T�"�'�b�'Z��'E2�'�r�'���'��)����v�j%1U�O$$M�W�'�b�'n��'�'�2�'��'��8��#R=D��c�����83C�'#"�'���'Sb�'���'���'-^0ْ�K+kl�0 �%BJ
0�'�'Ir�'�2�'�B�'H��'�� �/Y�qΆl���u9 �v�'�2�'R��'`R�'���'3��'�9���Kw��SvY=?10hH��'u��'B�'n�'��';2�'{����c�*�j�ab�,�j��c�'!"�'=��'qB�'��'���'/��x�k�(k~�a��C�+<"md�'�2�'D��'�r�'�hs�����O ��5j�=""vX��cόW�Х1���Zyr�'2�)�3?�3�i&�y���	D�%�@��:�8�FG������5�?��<q�nWt%*���(�z%1����������?�7�A��M��O8�<��M?i2#a���Q�e��D��	8g�&��ϟ�'�>5��l�syQ��Cб_0��JB�$�M�Х�c���OP6=2r����|�d����56��O��du�`ԧ�OK0�)E�ib�$+���lI0�a�uΓ�y�dx�0	�Z�>�=�'�?	B�US�v����C�X86�C���<9-O`�OrQo�/�c�@�' T4x�|*���f٣�
���'�X��?	���y�Z��cC�Fڼ�xu�U:D�)R�+?���|\����c>%8��'��I�~6�D�3�,�X��آZ�&p�'v��"~� �b�Ja&L������1$a|�5�VdȀ���W���?ͧ[t�$�c
b$��&�N�"�r���?!���?Q�. ��MC�O��ss�'��*����B+�&`���h�)$�����4�'�r�'o��'<Z�E���nm����DN�x��R�,"�4z�$j��?A���䧕?a�ʒ?�xD�D��hY�Q�-X�����M��i9�D0�	�����,$/� �s�=�˴eQM;�x�	�,��ɤ-��hّ���1��x�c�<���Q3jS�,Ô�*��!���R��?i���?���?�'������
O֟.mf��% �p"pE��$)o�dP���?�_�D��6M�O�p��,L&(���2S�l�R�'J#%�7���$k���+�l��'��'q|�|��G�6�a���|�&���7 ��ϓ�?���?i��?����OE�+��X�XXx��iQ�i+dT�l��#�M���a���e��OPA!E�]��Zץ'l0�ɣT�T�I�M������ŖW0�Ɵ����Ȼ󴡙�A�=
n`%ф#7q8�����'	��'�ؗ����'�2�'e��j�Ý sLЀ&�R�v|P���'�V����4U�F<����?q���ܬ(�@Uآ ƹ{�i�@NO���I#��D�ަ���4T����O�h�tNߋ|ڈ9�jۢ.�&Q��שL�t�hW���S�Q���[�	#O���bg8e�v�0ǐ��Iߟ��	��|�)�~y"�yӪ�3G!��h@D��K��`&�!yD���O��n��a�����N̏\���J�"B�HCj���f��M���i�x�� �i��	�]��Z��OF�'>+<m���ĉ+�"L����!�����O����O����O��D�|�ץ�C�n�����B�@�L�p���ר302�'���'�6=�IQ�ޱun��J$.ZK��Qџo�/��S�S�gw�m��<�q/V�	`<���N�B�Rd��<� Ɖ�H���������4�6��-AG�4B2ʁ�[��2j��R���O\���OT˓,ޛ�ܨe����HIe�1����"˃?l��b� T�"W������Ɂ�ē�N�B+�+g��h��M'���'�<�!,��mo.d��$m�͟p@�'v�bpg	�7���� �;T��D9�'W��'r��'V�>���E��Y��>4=|ҥA��iW�����M/C)p����[ܴ���yG��d�.�ɶ,��m�HS��	�y�'+"a�B ��v���x)RwN�J$S@�	�r\���q̹1�&A�����4���O$���OT�d� �TPH2�'v�@��O^�-��o��X(}�"�'&���4�'�(�Ӥ��
#�;�ѕoHji���<��Mr�|J~z�κ`�D	����kiX�QdΙ2g~m#4/|~�Ȝe��,�Ix��'��	kN)�NH<(� �	-9d����П��	�p�i>��'��6A8�.�Dm��3!-�'=�U�U�� O��$���e�?)r^�0�I���4���+[�.���x��	*̈\�U��M��O�0�pɂ:���d��� (��qVD<�]�Q���
�8Ob���O��$�Oz�$�O��?	I�j�~%��R7*
>��lQǨTП����ڴg�0�Χ�?I��i��'���Ae�4HҊP�A�D�4:b����-��O��4�Ƒ�U�r�6�BlD �'g�4}^������˒|��J��OT��J>i/O�)�O����O"ջP�Y˔pg�̊?=�{@�O,�d�<�$�i(& V�'���'��S��q��P<V�
�H�*�$�&���ڟ��I��S���b%�1BiD�������^�A��Y!f�I0a�Fp��O�)�?��I6�$S�|J%�Qk12�ț�ݜG����OH���O����<9d�i� %b���-R�h����'�`��"��'j��'z
7m6��1��D�U��D�_}:-��`���[�[��MԻi$^�;�i��	�^�:I�p�O	�'_8��@��H�Pr�����fi%���$�O����O8��O����|�ń�,!�\u�s�f/2���0Q����%N|��'�b���' �7=�`ѭډ\����@;�҆
���ٴ�y�^�b>���ͦ�͓4~��s	[q`�;�<u�:�͓8�(@�PG�O��[O>�(O���O><1��17K�Q���~0Y���O����O~��<9v�i�-c��'��'zL��P�с��ҵ�;�2%���f}R�q�n�0�ēp�T�P+�"D�5)��@�'A��3�P�$Up���D�� ��'����rK� e1DE]O4�����'���'`��'��>��$P��F��L��P�d�ָeJ}�	��M������]ʦ)�?�;Va�!�4�L�c���Emܩi����!�v&t�VYo��W$�oZj~��ڕSʠ���5�n�z��T�t$L<q��II|��b�|2Z���՟@��������맡`)��2f�$�y֧��W������6>���'����'�6��5$�!�Y�sO�)�^�ʐB�>	���?a֚x������B�ƊfV�\�'GXNXy��?z,h�`�O6�0�DQ��?Y��*�ı<���"�ƘX�a��(�v��_m�����O����O��4��ʓ5����w��c��1V���פ�~�b� ���y�oӊ�t�O��D�Oj�n<3�FI��_�+t��p�����4�¦y�'{V�k@���?��}���g�(0�̍<�詢���po�4̓�?����?a��?�����O&������0�d #0L�"�zxU�'<��'޲6͇e���O��lZw�I B�t�AN*H�A���s%2L<���?ͧ28��9�4��D!P:�Q���!=S�ňP�Y�$7��ir	ː�?�3�;�d�<�'�?����?�$�;9^m��g��"/0�`� �?�����DJצ��pʄ՟�Iҟ �Oq��D̙Z+qc�ҟt~�0�O.-�'�z7-^�K<�O��d�w
�h��p���շ!ਘf�J�{I�I��.��4�����.Z��O$���-͸'���z4O��b�nU'-�O��$�O�$�O1�j�Ft�XS���SE%��p��h��a1Ne9%X�4`�4��'���?��Ĝ-��`�G.�;:�b B��+�?���i�h<�U�i)�I�M0�3��O4�'H�&��V�F��ʹ� �#mf�Γ���O����O����O���|Pʑ,t�|YI����@&P�!c�)��Ƨ��+�R�'oB��D�'��6=�vx�O�&{���_8ʜ5�h�矰o���S��+xNqn��<yFOǋ't��Ef�P�±�tg��<aB�P.Xfl��+����4���d^�G\�AkP"���@@4 %+ވ��O����O��c���,� W���'�B�5A)8D�7*��L�����n��Oxq�'�2�'��O� �îӭt?���I�� �����)�~�� ��7���Wԟ��b	&n�nx���3��CW��ߟ���<�	��LE��w�����ɬq+B�0�o^�	�� �`�'�<6m��\���$�O�ol�Ӽ;�Ăt�D5atE�d��s�C��<A��i��6����=1$`�Ԧ���?)v�پ+:k��81wb�Z����6�W�O/h𐅍�����4�V�D�O���O����3un��2"�MFU+��G%c:ʓ@�6l�$=��'�b���'Eh��@�	r�z	ۂ^0$T6�Q���>��i��7�Kf�)擛wEҸ* Hآpz��5`̥$�RJp�Ӿ���II���Ԡ�O �QL>�,O^}��h�Oݞ�Rd���2�f�3I�O���O"�D�O��<y��i�8����'eV��6\2���F���Y8$�"D�'d�7#�	6����O���M�e����tht�c�W7�vK��
�s?�xmZk~R,��+���S[ܧ�s�A�[
�Dd�8%�������<���?A���?i���?��Dk+D$�[%�M�),��n�����'��j��py���<��i7�'I�$�b�Q��)��	�6vp���4O�^��f�g��iۙ+h7�2?	R�X�B�f@-$fOl��8X�%F��$�2�䓃�4�����Ol�dB�:4��V�=C-"\3�/�aY\���O�˓;��f��R�'V>}�O˘Ap�� V�ėA3νzcn6?Q\���	Ʀ����Ov����G!t�2p���7i�!F�(�j�S�n�8
��|��J�On�K>YeT~A1�D�μv�$
*J��?����?���?�|
)OjUo!.A�ZOE�u5�%J�F��f���Q�������M#�"(�>���&X�2��	L�3P�!1����.��6���K_�v��x�T`�#���~� �e�h�q�psc̝`�D��=ON˓�?���?����?�����	��	E|s��F4|� %��&ؕ׼�m��\�����(�	R�s������Sd���8	pDP�V',N҄aO�4E��i"8�O�OMd�a�ir��K��8:�+�S��=2��z'󄌣��Y��~X�O���|��1}��In��! �|�&�����?���?�-O�n�W�l������#���a�D��N�0`w��k&�?�g]���	�pO<�@J�qj$�����
8LP��_U~��C=����>��O��3���i�ɧ.�x�	%�ˑ�(@��-[�s��%g�˟`��矨��˟�'ON� ���?�R�
�v�\�Z���*d�?I�iA,�g�'���'
T��i�}@ҫY<*p���U!zɸ�q����<��41����~��mK�)h�f�	ߦ�Bd��?� ���
��arᩚ�]hH�K�>kW^��;���O\�4���$�O"�D�O��dQ�L�ٵ��5ZJ^��`��&2�V�$�Ob�YR���W������Od��ʦ�3?��ǐ,+�԰���,@��ɨ�cQ��?����?��C8�fnP�&���t�ٴ	&LPu�F:b�Ղ�|�*	��F�{�f �'�T����D}"�B`�	�%F�~0r��1��$��zT��	����{Q!�����Dx�-��fk�0�ѩ�� A4Hy�L�dή��@�1� �D+\�A`\�� n�	(�;�b�E��z�@�11��QSM�)Yn�8�,S�}�H�h�?�\a0����60��M �a�0��Ӿ�Hr�D�c��sf!K�M�"�]:����g�YhN��':��@�m��rP��@_K	�k�'u��3��CN�#X�+��`0�{Z�Hk9��A��A� ��{QX�Bwpp�Ûj��j�e@�@7�Y�C�~�:��Xy�|���� �m�%ܦt@�Ykҥ��Z��!��I �uÑE� ^����TM�M�E%P<M��� �#h�av��`%�%G�2;X�2B�{|0Ѱ�*�0��A�1�&�f�9�^�����	�I�X����&R1 ����3�?�O��I��$�@�d�P�R�
� 6`|�'��æ �v
���ï^�s��>i)c�B'u�Ra3�M�b����1}��&�?!�y���J�y�� ���/?�� �/;�y�LG�.\�� ��\�2	(T���0<��	!]��hbCOҬDn��p�ɪ_��B�I�N~��`�\Jn&d�Ǖ���B�	Qߦ�p7��*Dk��HB�ɔ{CpX�ዓ6_������Ec�C�	2o�P)IC�|���hM�)��C�I'T�K���L��h�.Q/To�C�	$6p4=f�%,���RN�?DDB�/VV�l�TL
p �� P���6B�	7&���sdN&J���@�X>g�C�	� <�I	5�^�VҐ�(5튰q�C�	�	
�ke@�2;���Zp(H�NWbC�I(d���kˑت4
��+7jfB�ɪi�n��%F�O���Ù��`B䉉[����F4l�! ��OR�B�I��ހ2�e�$+YS�Հo�nC�:bѸUHv� ]�@*��S�ULVC�I�}C��S���P\����i��I\�C�	0�r���C�TJl�����dDJC�2�|�A�?D
�S��3]�C��56�l�6��pЁ���a\
C䉪`�й�0g�"�l�0�S�x��C�	�B�f�eK̎_�ڹ�PLD*bܞC�ɂ]�0]Z�l�/�������C�2Pp��o�,E������C������ލ�����E��C��5簥{f���E;��xF����^C�z B20��:p36d2l�8�lB�	(i�z�����5�	�u��T�ZB�2
KP!��,ɴzEd�l�<
^C䉇$�j���E)/�B��3@�*^jlC�	=I{ԁ��眶p*>={rJE��B�	>}��Q!fΜd`�3��b�B�	�H`��]=Co��X�/N�$<ZB�	:}��0���<#{��RPׇeOTB䉍U�F����D�f�k�nT�<B��h�\r�(/�Bm�@M�
	�B�I<b�ؒ��U (�A�e�K
��B�)� &�����*�T���ֶk+Fl
�"O��9��܇o+��seE�:3��:C"O:�K��1<��(��Ƒ<D�7"O� gi�
,�dȊ�!X�c�����"O���.J� pԯ��}�b"O��`��%.��+�/�)%B�Y�"OX��ǒ�TS��L�q���"O�t�΅��!��~Ҵ�`"O�x�ȅ$q�����KϪ!Ĵ�1�"O��K�ę[� sK]�H��AR"O��k`�E����`�Jw����G"OJ)���0O������ b��s"On��3i�7#��u+Uɗ�!�T�YW"O,�� �Ŷ��`*����W��	�"O��g�GwY������$��5"O�Q��-��|��@�b%L(^с"O�0��f���D��/
80�"OVH!�'I!3�k�!�]�"O� ��*k�H����2e�y�f"Oʼ��c�+76`���/ވD��Z�"O�H" 3pЕ`3��&O]z!ɒ"O�PRa�+��YY��(/-x1�"O�9p"��k1>�!�E�2�E"O�Ř��N�����U�E���� �"OVL�Dw�Keh� +p
��"O(��J��s<Ѝ��ǁ�)U\��'"O:|z��Z*��	v�O=<C���"OJ�2Ϋ1�N$k�;���"O� E)�n}���\���a�"O���C`ՙ$6$�
gb�4O�p�j"O
��5mC�$��8VD��#@�퓣"O�x�R��$n2��
�d��F���bp"O��E��f��!x��m҇"O�	놀јY�t�:�o]"U:�@��"OHeS��5PaöNN�-
�D"O$H�`(D7|�J�dު��9�P"ON����♐���p�n���"O����
U�<�
�I�j����"O�-B��W�h���#��h��xe"O�+�ٲC_���p�p"O.26�\#$�q2Ŋ1��1�"O$d�j�A&ډxe���C�@`%"OH42�Pvh���E��M�a"O,��"���i"��B�� �l<C#"O|t�C@�7 j��ǆE@À"O����޿swf��%��9N���"Oڐ�T���B�Ƒ:w��6 �@"OzH�Ī�<%`:�a�S�*8$"O`�o�E<N��&N�&-����"O@�QDT)|{R h�cɤ@���R�"O��2G0S�x� �|�0��B"O��kḊ1f���0�Zz�Z�S�"O���|7�Tq��(<���"O|�th�
$���Y�ZچБ7"O(Xi w�$�ℙ/RT�w"O�=�U��^kvIJ$m�J�vA0�"O�026o�3r`Y�k��c���˥"O�Q1W�Z�C�N���#�8\��<"O1�a�!v�x@D�,i�2�"OV�����T��j���6�Dٹ#"O��I��ݢ["�D{�H�%Mi�eK4"O ��T�� L6�R��Ԫ=���e"O� �,�6L���1��|�J�cp"O����Ͻ.�U�aƔU�ڱ��"O� ��1a_�N�x��U��e�Q"O��0MX�{.�S�j	�6�Y"O� Cu("@�P�A�̵=���7"O%j�J�zx���#dܠ"O��a� υz�V�8!��_���i�"Oh�u��=
l��@_#\d��"Opؠ0�4Y8,�c �({�)�T"Od=1�a�$o{^@����.[�(�"O��Ӏ�����>��z�"OV�&HR�nŒ�*�J?E����7"O��4��1\�F!
���(gx,!�"O�� U��6l��(B
��5D`}��"Oz��"O@.��y�	�=N|���"O����O�:��+ ��?3<�I	��>S�{���OW0ih�a��|��h�B�1Z��a�'`��ⱪ��
��0�L � �D(@u�y'�m��Lȵ��<�E"�Y+�x/ �-L<9�扁 P�HD�1X����#$��b��1���R7ę
>��q���&OĉPvC�pܓ*�d`���
dy����*�n��ȓ2wt 0��w���n©u
�y�O
��̤����O�v@�W9r4�'m�D��H:�'K��M�n�I;G��F��81�{������I�g�����
�i������<O�C�	,�����t�·`�i��=B�)ܨ�x�╽p8l�{c�
*
`�*�J%��<��4U�1O�Q��	�DM��g�lwΘ��"Oμ��+ʂ(���ׇJ0-�<0q5�x"�� ڤb�b?��b��{K�g��EEj%"�I!D�02��ك`��4�&��Xd�R�1�	6Y���cÓLM��A��;I�T��g�(F��ēC�*�Q���k�|��#f�2�N����p�!�$@��Fȋ����lȅ	�#�ayFA��b���:1]TQ"�[<{����9D�`�s��Mخ���[�p���F9񤑗t!���>�~�0j�
?`l���lI�Y�^�0g�T�<A��^Lg�j�o9$�*l_Ը'�j�#;�3�R,��#vI����\�D[�!��%c��YS�(��/:��@�#���2�&�uNa",Ҙr)daČ9��	qg�Gа<Q$�ڸy���%�����4~iX�Q+�2'�E��0D�\���V�9�|����~��(�A1��T=��R�{����]�\�R�I7rb���y"gќP�x��0NW�`��)�I���'ʺ@Q��2O����D'x)��jQ,Ϗ
�ئO�)�Qo�2�0�1HQ2��v��z5I���� E,D2l���C�ե}R����I�`�B�y���\��4e"��y�*a�R�y�К-a�����܅}h4��H��ēK;PiA�����D�ʥ�T�(rLHH�B�o�!�Dև#&���*^;�q0�坑X�OLh{a�f�(�d�~m�Q3�0@�p�+�;4�,��K:W��Lp$� I�\r�a��N<CቼHW�%�$��s����q\>8�C�I<ҕX'�I�Q���܇YpbC�	�<��"A��]d���ba�)�^C�I-'�>q�B�IF}����6C��;V� �:B��4��'�	�t�C�I*z��d�q+�j;*�ː�D�cr�B�ɝu�yzw�ɳ �Bi#H�Q�B�	�@�`�)�%�mzB��.w�B��["H-ʄ/ʐG��SS��(ʊB䉋@���KvÝ�i+�hX`B΃)�B��-F��	+f��-V��{s���Q\$C�)� Ȅy��F�W����J��/D�;r"O�DpAcQ�`�h��h��;{�ʒ"O�m�@bA�6��Pr埭tr��$"O�XidA
�A�J�갩�2kb`���"O}���  Y+؝��(�?P>��"O�JVh�1�a�Q��8FlY��"O���c&G�_��i���֡Y1Hl+S"O�LY�l�?VpJ$r�Ā(��"O�[�
B*2�q�	= ��\�`"O��yr��N����3�I ~D���"Od,���3��S�Kײs��*�"O6��'��=�u���S�S�@p�"OZ8 �I3!�� 9���5B�� A�"O8|j�喽n} �����-U�d��"OQ"�E�I:��HдY�X��"O�<�ӣ�;�vT�s�P�a� �q3"O���f���B����D�#]�\�"O0�h�e.6c�����j��h�"O�����<�����[�f�0�"O��YaZ�i�:�IA��$ ���"O^U�a��t��� f۹��#�"O���C"؂'��D�cS-9�\�:�"O�ѯ2<��	�uA�f�:�)BT�<I�͌�Y�����z��)��T�<�.��E�6E�E��$2��RFQS�<i$n�#F�"y��F+����t
�O�<���"�<!�3oG��hS�%�N�<�Q�غV���UB�':^N=�� �o�<�eG���`�h Ιd���C3��m�<q�
�vz	�w`�t�� �u`�h�<	G�T+|HZA��b�'C����(�n�<)bi��d\T# L�Aμh��Pl�<���K3?`T@�/[T�Y�J�i�<y��� u�D%38N\ ��Af�<!�/��)�@�ص$K'�xG �L�<���̩	���`$�"��aP�(UQ�<	���\� A�IU�G�^�	�FAg�<	���0o����YQ�n�AE�f�<��<s"�aSDV>*�0tR�n�<��"��m��l��W8k��*qjSh�<Y����Q@�h+K7"݌X��f�n�<� �0W�<�X oJ3_��E�G)�m�<�0�-��k&���e�h����_Q�<b�з����H�Q�D�3�	L�<�Q�&gC��ڃ�۹"�ۣ'�I�<A��p���������\�5�Xl�<QL�2|��L�U���H$��g�<�!$ܶ��TS����#�-h�,k�<q�"$P1���݂uW�s��f�<��i��Pb,�` �5q"Ak0
�[�<A�A��!�<�QY6)����aV�<���F�V8��PŘ�=���:!�k�<��a�[�\��f28��ff�e�<!C � �P��E'� I�����Z�<�G��9���Ca��ihUq���X�<q �ŧ<a"1�A聭
}ā����T�<�"S�eӖ��Ug�d~K� G�<I��E������tb@,���N�<	ǦE�1����Պ�7A��0)�gDE�<I�w-�1����?,X\ Q4�]B�<!o��0愴�a/G:$<y�	~�<����or����5S���'E�{�<�uB�gY`�Se�Fr���xDb|�<ad�� @���f��ai�)闪�B�<� ��۔c�5M$�X���±C@��y#"O�@�hG�.��Q�N�ha"O��s�m�+fu��fO+��02"O �i!l�E�T�J�%��A���W"O*���,I
����VJ��P2^�"O0q�e�[04�\���Z�y*d�"On
t'=c
��dD� �$�Q�"O�8ё�ڔN3:�� �
��1�#"O�X�eϚ
��)����ܙ��"Oҥp�g��.2V�1�G��Q���"O�H���N�����`�K��`!�"O��pk�5u(|�� Q�q�*�"OP�{��1�*QU���Jp�S"O:I�ƇWB���+�1��9��"O���E�	b@c�
˰$����"OZ��L�dƺ�����,H�ss"O\����u�N�s
�^ М�!"O#�,�8~X�a��L4/�9F"O��*�'Y$����F$/my"O�Q���E!V�IyWCU�<�A��"O5�C�Sx��|;���5\TPat"Oși��\�=�h�!0
T)9��f"ORl�W�J�u:��i4�@�a�@�"OP��k�J��0t��-59C"O:�Ȑ�� �������\,�"O�9�M� Qd�`Ip�Y!u��"O!S�&Qf)lJ!#ٛ|�,js"O�99@��"W��(c� �$��f"O�u�R�E�b�p���qrR��"OJz5.�S���ta�F��#�"O�m���,��d#�a��lͫ "O�Iz�eՋK�n�3��� y�E"O@������ �)gA�SJ��S�"OJ�3�l�7��Dxj6{4l��b"OJ���%ak~�����7�P��"OXi�钎` J��J�1hɀq"O��֢�l��ţ�Hӿ[��5{0"O�Ha�ڊ@hR�s��XAzq"O�,Q�&�>N���
(Ԕ�"Ov�����i:�0��f�v��8(A"O�"����@�f�B���"O���C8f8@�1E�}��A�U"O��Iw`�|��Qq��^9|H���"OV�:�
J9E�8Q��*�e��0"Ov�oe�uW��8�)W�H���"O\�8� �;.�1���?��I�"Oȡ���A��!j�dվzE>��"O ���#�>X�CDG��J!�"O> #�FA"DvTd��� `z%B�"O(ux�l=M���hrGD�B\xy�"O&�G�:�4�Kq�Q��TT�"Ov�XT��aל|kc��*��QF"O���#
�a�@@��i�7`R݂T"O�)�\�tb<��5�[�{�T	f"O�%��A�z�p�aa
'g�*<�"OR��"��=@�8�8��ݐ���9�"Oz]��	�	`�y�.R�g��j�"O��doͣ�3R-^Ss�E*�"O�|���M� �( �K�a���"O���Њ"�x��ӝA�����"O�ఄ�Z�C�4p���8p�����"Od�QFB�Eh�Tѷ�X�?�
�`�"O�-i���seR����i����"Or�є�O\*�V�Yui	�m�*H��S�? .9�e(]�I-�Y�0(B+��"O:�)�H�X�1��Τ
���Q"Oΐ�eBÄOf*� ��� �$Pg"O�7CȐ�`8;�סm�x�&"Oл��k`�EB!�F Ւ��$"O�����	rR�*i�#����"O�qqȐT�E�՝t2�*"O�$�ՙI�+t�^]�|�"OڰS�Iڐo���k�'�G�"O�9��P�3��$�)O��p"O^���3P�,�ӓ���TZ�C"Ox���G64�r��d�U�Bc���"O��$���51b.��j� ͡"OƼ0$e�!iC��S���)����3*O��C�G�9�H5+4��LP�,��'��A3�柱f�
�&���r�� ;�'=���� ;��Io�g+��8�'�0�Y���6�x�6nK^�*��
�'���
���,m1�Ɇ>,�	H�'S�<p��׼"Î�j� �;*���'��(��S��(�R0��7�0y��'m4ܪ�FR�G-�(I�(6q8]��'�bx�AC95̀!�GT)3?���	�'zn����Aa��v*.WN�	�'�`���k�6b����ԁG0$m�	�'���p�#)Kl�ܛ�D3��y���a��\��F�lK�����G��y�'�/g��$1�ɋ�6>��3�)�yr*ΡP�Z�����+6�)�E���y�ČF�9Jn�'��<��K��yR�T�^��7�E+���GO�y�oz��֕	n�����yrO�s��
T� �i�w��yr��B�`�A���0}��k&�y���j�b��s@���܅3���y2b
	��$��T�%���Z��y��B3!�ܵ��)�4ά�sƍ��y�# ��}sn/�Z���A1�ym�r�&�����i,Yk�	�y���|��9!CQ8	��}C��y��W�'VѲ��RlHy�H��y���:)5e	���ţ۾�y"��YP�bSiD�M���+�M��'���A�V4zņq*fĐ�}h�TA	�'�QcfKF	�|��U�]tg�P�	�'XUC���&�|��͇ n�F��	�'�8I�3���)�
)kUm��FUJ�'���cE@�%����� �ST؈
�'�T
�O	nj$,���(S�n���'�����i�?��H9�UI�|��'� A�wN�5���� �U�=�	�'Q�epB�Y}4����I�$2��	�'8����/�mJW�(3W+�%D�\�u�eA
�G��p��L���0D�d�2M��'���O�����0D�,� j�� dJ��1Z@}0'�4D��JA��jEX h��a����6D�p�e.�d$����+P���6�.D��x�8#���d�3��J��"D�H
 ǆ�K�Ja�G��$1� �b�%D�\AQ� �&���WP�U%D��q���������6["U;s+ D��q"lO�0y:�s���!t"Re�?D���N1$$�@���.�{Uk2D�� 8\*�j%��D��1xZ��"Oԝ��N͢b��ui!�֖9v<5��"O��k4�,1t�0aWl�BL8�I�"O�#U&رA��-S�ˉ�b2\53�"OvH`ԡ!�ܕ@'KΟxz�YE"O@�B'ܙuj������ۄ��e"O9/5�F�a �R�*��	���y��T���E# HJDp���H�yJr
Ȉ�������{`D ��y�,ZE�A���^\�Cg��3�y������`G)Z��VJİ�y!�	Y�����[tw�I�(��y�Vt-b��v���@�Ȑ:����y��y$V���K�:	4-��y"����x�HF��#A~ld��I��y��9u1����F��4"<e;��ǌ�y����z ���-+\6y��ӷ�y�.;����KQB�@2 KG��yb�%bh�EC��� %$܂����y+��ֈ�Rd�� �:�g�*�y��L�'a���QHH�rT"xW����y��% �Q-�cT> Zc�W�yM�; ��Q�S�_*jmL��+E�y��.�Z(��90�-��h��yr��,����P���Pb�啍�y2 ��eئ9�q�ǌ�&�ӑk��y"fFnǲ@@GJ�z�Q`�0�y¨U_�"�CҎQ�i����&i���y� 
�% 0,�1f��_�X!�c��yB�N�}��@�Y&ej��\��yb�ْK���� ]3W��l�V
V��y2"��3Ț���T�w�)5I�>�yr��j��s��ܡu[d%kE��y�놶O��,)j�vA�������yj�z����"@Y
�τ��y�K�\�j�x@��lz�Ѱ���y")�S�(I	�+�j����&�yR�F��= �(�Xu2={�.'�y�nʌ0'�,�t(��E:H���+W��y/C�-�:0�T%�IG�P�����y�x����E<v�@��.�4 �	�'��gEV7� ��AS�L4옘�'�j�(S��1s��c6"�A?����'tj�0��4Z��`i�@��-��'��-X���>!�^���fھ;Y	(�'L�=:`�G�/�V�Fn\3,���'	��sN�چ�"��D�B��(�'�� 3#"����F�B�jm�'̀a6)W&�бp����9����
�'!f��n�YdX3�O_#.��L	�'�l��"�'5��k�L�2\�����'G�aB
�2Q^%(�O)A�A��'[@��a��8(H�x6,�(R�+�' ��R���cf��B���'	�X�z�'��h0�ΒQ`��z�`�y�ԘZ�'�9�!�I2�;��x�Ry��'?j@���L2&�tlʐM�9h*�80�'<��y��(`LTʀ��[?�]*�'���B�I�ۄFޘ~��-P
�'hV|Q'!�j�r<HՌ� L� 
�'��0�Ӹt�Z�y�W0��E 	�'��H��J�6�48P�_����'-:h�����
5"��5l����'f��i���0}��#�dIW?�t���� X��!N Q��� ��X�,�q"O����΅(]���P�a��(�U��"Oz�:#��mg&��3���fE3`"O`��& ΑSv1��G 'xF!�"O@i0��-%3�a��%\�R�"O6 Ѳ�	(�x�1�۳k��"O|��+�3mX.�A� ��c��j�"Ox�`W8pl�x�`�1����D"Ov�b4)E�,l0��8E�J�'"O,Myw*�4v���b��"O�3ɕ1K*p�#��ʷW��T"O��Ë6����&dF�%�>��"O�|:ݎ�J+����!���D�F"O��At��U�^���\T�@��`"OU��\}9<�A��I�p��L3�"O�T��/� c61n�{�P�9�"O���}K|}�n��GsH�[�"Ot]#�� �kCӾCWhxs�"O��*� L.(����P"^7q�b|""OT��Ğ�e��T[ᡂ�6H�#"O�����,�N���U�#zY��"O��JH!	�`Iz7�ӑVt��В"O�d�g���dE�"ʜ�_�di(�"O,s���-fSj�)W@�u	�"Oh�K�d�1-����)"�v$��"O��p@�ƍm��k!�(�Шi%"O��
��
b�����)���z�"OH��'#�'&�N(���%��R�"O ��o��S�$س Ǌ����"OXHA��"t�^�@�%T�HA��"OTp)q�q����T,4n,Q��"O�1S���\a�dU��-Ĉ�y�%��bU��x��k���HE*���y��W�Je!�o]��X{�BI��yR��0�x�
�R��Td��yb����,��󆍹B�|����#�y��(O��h2�&B�8!$��<�yR!�za����	r�(p�Z��y��H�#���!d�F^5�p���y�M�L��B�T��08���y���7g�0(�p�e�1 i���y�ׄL��|+�L�i
�4��+ԡ�y�[s*P��ƚ<]�(���J>�yM	�y"`�xÎ�&*+�O�0%��-4��(c��:B;��G���RU��-@L%���@H"M���kf����t�񡷎Z9$�ش�P��.?Y�8��,[�Y�T����hh�O�&r��ȓ+dh��=K$9��B�%E��e6��&&| p@��"j� ��ȓ5��V��$'��oX�-��D"O���#�;bJ�"dO�M��e{"OT`{w�ӯb�V�I���Fo�y�"O�8 � ۗKr��3���1 ?���G"O8�[%a�/c�d�k���/$Z|��"O�u�a$�zE�uq��$d6h���"O H���*B�	I'�3o?@��"O|=�aW,H+��c'��D���"O֌�ɀ�,��<�Uڧ.�lە"O�	S�Ȅ�E.�i3��#��.D�|Q`M��I/֨�5�5C
�"/D���W��$�h9�g.�DASrJ,D���'�hYfъ6��cGB���!+D���2'�/2z�(� D��e��� 4D�� ΀5<:(�
&/G�XO%q�"O̠����i����ƯLG�,�s"OzE�bX�,��y�.��Ht�w"O�	uiԽ#;<���' h�t��"O:-�����LshEx��N%#���"O,=�3�
�J�ESUH�� A� "O2�c�o�2�2]�Q!�?�y1�"O��:V��+-Z��BG���$I�"O��1����ؔ����*zǬ�s�"O����J�]Ad�R��V�W��$��"Ox���$=g`$�'.	�f�ʔ�"O�Ł�柺b\̵)b��1'�sQ"OJH�ԇ��K\�y"�Z$�yc�"On���$���	k��詶"O �EH�aHm)��m�QcV"O(��H۳`��`i��E+q��P"O��RQ
ߵ]z�@:"��sntA5"O���w��dI�QQ�*]�q��	!�"O$�k�!�#[@L��&(p�q��"Ob�ˡd�g2<zE�[-���Bu"O��`���D�i�n�:?���S�"O������nsqN��5��eY�"O�@��%H�0���/  �$�a"O|���)�!$�puB#N�;�
Yis"O����&��LȐp��x�3"OP䘀$�7`<�{3\7I��	�"OXыF��[_�I��ѭ6�~�V"O� @c�֬E�L�Zo�5"O(�Ҷ��6E2�]#ѩ̫1W$�6"O��P���q��A���.SK���"O<d!Љ"B�aڤ�H�&bH T"O�caǱe�5�6Ǔ�WK�՚4"O�UX9� �耯6IG�@�p"O�	�[��.@�l0�|��"O~|�6�U{ڨ�F�z�ޤK�"O*�6��F(�	����.ނ�(D"Otl!Gŵ9�8a3b�*�di0�"O�)���$FV��ʝ�p�9�"O��j��� �Jȁ �N�3��c�"Ot cc�#�׫2b�0�8�"O����oگ(�,S� ̩(�B��g"O̐4�H�a"T��PO�	Y:\��""O��x�΁�/��lÓ`�Y/v`�"OP�	3AW!
�qwj�S���w"O�a��Q�E@��ʘ9	�4�"Ol�)2�`ta4I^%.��q"O\	�#���lJ((���ޠ�:ku"O�āSj�	@'�8f��,Y�xUZ�"O����(@(c�A�"M�"Or�YC.I�:�йk��e��up�"O���#�#)Er5��͔;��=C�"O̴�6�ԕ;��4��a�/w�ɢ�"O�x"�	Ӆx�L� 5c�K\��K�"O\�����n��@� ��sYr-�t"O�43�ݟmFYӃb��SI-��"O����)J,:�ʌ(L�AP%��"O@!�(I������-D� �ʱ"O�ݰS܂Xj�����Im����"OJp{���K60X�M�hQ^�B"O�PS���3$Yf����#C�Z"O���`��@��h�W���-�b"O��Ub#%Ƒ����J�I�"Oʝ��ϒ,;f��R�a�z��$�!"O���w�85�b���K4�Y �"O� \��Фӊmb�� BA0�@��d"O0�S�*���yU ��U�VC�"O��	rM����ᛐ��M��K�"O����V*�L�YP��z5�D"O��p�K+�`��r-�}�"�"O�9�k�A�*x�P�Fql�)s"O�ձF�""�8t���<>6�Qq�'��0Jt���ΐa�"��/\��� �&��5�O��hׇ���<�j����CǪQ��"O��#䊘vۦٰa�}�8�E"O��h2�\�z�4"у�0($#"O��� 	��H���qh�L��P"O����1��@��F�h�6��'"O�]���I��y�c�ʏ�z��"OR�ڒ*S�8H��Ca��-$�"O��� �S%"�>�[�BJ`���W"O��{#�x��(��E�wRU�t"O���6抄W�<b��e�`Qq"OP����j6p#�n6p�b��"O~,� �ʦը��ʁ��u��"O����\,��	�M:�LH"#"Ol���
�z�ғ�.(��#"O�(b�j��hBJ$�&X� ���c"Oʌ(�iM�.�~ur���$	��@�"O`(�Qc�	K�`��AK�#� =�%"OX�ѐ.q|L�E�.O����"O>��`̂��7$�ToR�@�"O�f&�+ pf�nQ?!~ԸY�"O�i�D�*0ɐ���
D�}n��J�"O�,0����K���!��LSd���"O� 
��K�5Y��JW-Y'T?����"Op2'VZF�A`�X!6��P"O$[ӊt��q�&�,u��P`"O�5�#GO5$�����HS,VzE[Q"O,!`&�;u��% CBL'H@>$��"O\Q�§6l��I� 
?$=R�"OD�FVX�ت��&�����"O���pO�O���Qt���{�PXz"O��ʦd_�<~�l	�kJ�nmB)z�"O�M+��I�J �%0g\,9j�t��"OX�s��,+�t"$�H48T����"O��'̘�N`��*�(*J0�hR*O��٧��w�J�Jլ�p�j�'�� 2Q-� Ī\ye�G<;�Y�ʓ7E�mHA۸o��CV"��a�ȓJ��e��$Y�.#�����ETe��s��|@B.ܸlG�q�)?d�-�ȓk,T����LP��z��|i8��?�A��ą��0�cm
2�� ��2Z}� ��-F��pMG!fw&��'�a~�*K�L1jQ;G�����Ө"�y2�z����5�AB��S	���yr,B?7r����F�z�A�O��yr�
d��u�bM�[����A�_��y��K1��IG&B�S�^ 9����y�ӥ/���D;T���!�)�y�CÅj�H2�&E����կ�yBOW0
/8���BLA��ij��Ͳ�Py�KӒ^O��r�ő.�ޱWɛd�<��
�8u�(�P(�%��$�WcY�<��DQ&aP���A�k�<����R�<�E�����@�ɪ3�ȈQrL�<!S��"B����fK�3�x�����C�'��i�š��'j�4�3&�� �B�)� ���!�2��Bq����"O0q����s���`a��O&��4"O92�N�a��Ʉ�љf����"O~D�$�(�t�A4o�a[U"O^M��	�RA�C#OH\�\k�"Or%Z��;:*,�AW�	��ě$��O��:�'B�Ҡ�ҫ>�R�������ȓt)�!�Rb@�k�P4qvo� (�.��ȓqOũ�f�?$���A�9&~|�ȓit
ɚ���.J�|���J�;9;~��e�(}���ڳq�����۷(����ȓ-18t t#T�U�ڼ@ ߳5��ȓr,��ǭָ�~� �_$��(��
m&X�#*�:���JR����=ℚ��?v�$ �	-�u�ȓTv�(L9�*���˖�zx��3�ܼ��mǩ76�٣�`��tcTu��!��j�eR2~�t(ʳ<������P��K�J�'�2r\�-�ȓ=���C��J!@��d�ұ��Q��X��p8�ɇa��t�� ^0$�����P�ά�&aB�}�.�'*եq*\�������qg^����K�@��9��0��X*�cM�3ސ5�#N�Ry>M�������c٫0)<ԉI�y�ȓy�l���?��8j������Q���k iި�z%:E���Ҥ���=�@R�cRcz�]!Kpv��ȓ6� ��'t�l�2d �T���H���shB
#�rH�;�R��FM�I�[.r���և[<�H��ȓP�FD(6AnW�b���=:�VI���$�&��4B4�9.��`�ȓv0V咗��N����N�>:��ȓF�T�B �J�M��Nީ6��I��D`��W�$��l�ɕ1Rτ���G�@@���׸�:��V$���ȓ��� ��0����͋�<����ȓOj��Z�-r�����	43ZF���{z��3s��
Hhd��d�1��݅ȓ`|L ��-�cp��i�`�9Y���!�"�G O��I4��Q.� �ȓP6 :֦�.R�r��o9��ȓ)&rH���̭f��r��N�s���ȓob�I���;����&� ��|���"�K�Mqp`��S�⌆ȓwSz��dj�3���ND;7����4�T٩CE�u1�c�Sw�,M�ȓu�\���H.ts�ؠ��3]G(��ȓ@��0����m�S	ú8)$E�ȓMw:�s�I6Q��&^4K�x��{�����`�n5(p`�Y/����'�9T�]�S��U�����m�ȓ4H��%�a�p��֡^Є�P����E��N0c.U";���ȓ:K�,U�D�H��V�ǡ.����d^a���qp�4����'Ue�4����:���d*����&�n���ȓ$���Eɺd��p�҅�i2�H�ȓ/��1�ǂʒ@Od�H�G�-�,مȓWh&�s���<y��N�Y�Ņ�Q��A7%ܛ{�40���T�C���	R���h��$�?6`}�aV!�(���0.E!��D�r��R��)<��`�5
C!�� ���B�\6�:�DD=Q�Щ�V"O�M��E�i#Xm�'��L��8
w"O.��ET "b��ۃbX��ae"O頤��b��(�aͱy����"O4�w.$�h�{�e]�*v�7�'��OX�}�j��P�ƕ�=m`A�'@T�i����pm4�/��^o�����?a��$�ȓԌ	���X�A�xݓg�Y�f��0��H[�����.��;��P�L%�-��q�8E��5��t; k[=5���ȓ+��sS�\5?'
��Tk�<k�X�ȓ<�@�B��m���cmS�a�B��ȓ`��P�ì�6H_���7��9"�I�ȓG���bc+�5p���'�D�4z��ȓr}����US�=F�ᆩ��{�X���N�eېc��T��m��d��y��mY��
�6�`��>�����xT�soX%v�<��%=d��5�ߓp2�����Y�]�|�ȓ	��A�ԩ�j�H��'`�>����%���Y�@�
m"U�����+�b0�ȓ5Vy�P#P��a�!��uV���~ڐ�3�C RdٹŃȷ\J�X��2����8	H��䮈�b,�U��j\��T̓��f\���C� 1�ȓ'7 @@\�.&�XI�O�.�A��Iì���-!�pA$�[x� ��ȓDj�;2�D�!v�k6��Sc"��ȓJ�fPi6��1�c�hО�H��ȓ	���]ju2 �TL\� ����ȓ�Ԙ1� "��S"� �.eD܄�*��ERǇ�:lv�K�fH�Ld��/��i6��36A����b͝5W�t�ȓ+�Ne��
�'$@�Q24FU��x�ȓq�||��m�>2�`qƈ�G},��I�6��!Q C��A!׊<��8�ȓ#o�ͱ��Ѵ3r��"B߼C���ȓIV�% 6 ��;��d�7
[�K爰�ȓ/6�5p1H�3T��04"��M�DA��R	Ƅs�%K���6� 
�⨇ȓ`���4��H\h0l�
�D���S�:�x�ǉ�)K��Sၧt�4%�ȓ}���"�e��r~�Sr`םbjZ���?�Q�u�ʗu$B�c�6���ȓE?:)EC�� �գخ}T�ȓyV�T$M5g�(���z|���rd�5ce/��fZ��Љ��ͅ�)�B�� ;r���n�n����"d�52d�6:���@I�`KĜ��7������A��S�"���ȓ
"!����!��9���Tm�!��f�T�����h��iA���Ć�(���q�m�@Y�M9L�P����C�'���C�Aƈ�ț M�9c	�'���P@ˋ�O�j%�aJ��Bz����'�j	�	U}ʲ��a�Y�j�4��'��Ś��غ^�-K���,i*�'�D��LN�� l37��@b	�'m��j6gûw�iؤB�-��uB�'��I��\�+��!ԅ��!g*؏�d+�'|=��0���'�b�����[=&���^�\��l$��E��ό�+�ȓO=�ha�e�wN���2�Ӂ0iZ��ȓMMf���Ȳ�@�?if���S�? �����(C�2 �bLۇB���"O���41F�1���%��}�G"O�����W�i#tĻ�$�4g�vQ�#�'0��2) V�Όz2��)$��� �8D�4�M�,�(L;���q߸�1�3D��F���{�����;ar��-D���#���^}P�
U�^"Hmd�,D�4q��ȫ^�,�W�6f!@8�7D�\����86�l�96�P�|��	Å5D����+۟$�$�{��X:!¸��2D�h�� �/]�%�꓆{X�Iq�.D��
�兵2D94+�� JyXR.D��V�ņ#1� ��_0Q焰�4)*D�d!���$w����^�o���'D�p�a�V��f���)��*jz왳�+D�p�e����()q&I?&��MyC�4D��cHE�1�p���	�B�e��A1D��pÛ-)0�8��M�>��D4D��" h4B��&�L&G�V����O���6�O�9��\����SfˆL'Ƽ��"OX�	WlS��5A��	^�i�"O"�����5
%�p��#�Tӕ"OH���@�I9�蚂�h&�P!"O�1�`��=�0�))���kW"OR���#�&Y�|�QT�5����S��6�S�iI�7�
@�7�7]b��D�	3�	Y���3W�*3������q���&D��"O�� آSDդi6\���"D�<�BD�m���Rs�8<����g&D�`j��N�,*,�Nf�r.9D�4)֊�ZD�2����@��S�3D�0���6��ȋv&ҁjS�KC��<�����(���("��S�B��egVN�-��"OFy34Z$'��1B Q�@ ��*OH���;X�H����2֝��'[���ŗ*�eB�l���Y��'����"ݝ4M��M�D�<��	�'��Q���ʗN�����Ҳ@j��;��d%�'��aPP�ܑ?�l��R዗fW���?)���~����R�Z$Q`���?�|���q�<Y���qd|�uK�%/�\�!t�l�<yd�EI�*�P>~��%�|�<�D�N���YVHR���@��I~�<�w��5���0%��_�eAT�I{�<)&Ț*ݎ�'N¬+^1I᫆B��hO�'9���h�(B�!Q��[��� $����	�D�����6߈����Ն'�C�ɨ}��\�R�P�2� xt˔N8C�I)^�Ј!+\�9\�q���7!��B�</��Y�Ā�4��=�Q	�6 �B�IF-|��U�@}����E͘:&��B�I�fX;�,X�(�����f(3>��=�
�'Hؠ��d�zit�]:B�Єȓ[W�P�U��D�pqپzR�=��f����
y����+bz��"B=+�yr�[,	������KrJ�Y�$���yr�J��!G��;�4HA�Hã�y�%ۃ>����C�\�|�A����y�\C���q���[`�)Y����yb.�x[콪��Q-*�hP��y��ה:^���jx@M�w%��y���\�hE�%#v@�4�g�ݮ�y2dT
̼�y"�X�t����w����y"�R���Y��L�	m~(��f�@��y
� �a����G��R��C�;�:@j""OD��eiҾ0��{�ۥ#�d���"O`������VИ�[���Uw���"O=0c��!y�VY1QK8�Q�"O��y�d2��]�@�2<�(V"O��paG�,Oa,��nރg�4"Oj������g-f�B��"O���>���:�Iʷ2�Hq�0"O�đ��ɊeSd%�G�\�d�J�%"O$���'��lB�	L3wży��"OX���nծZ9=�S��F�&��"Ov��\�\��$mY������#���y�Ĝ
v�lj���&�XT`���y�	T���u3�Ǐ�<x`gP��yK�w�*ic�H\�	����/���y�������7�������y��\i���Q���i���*����y�l�q�ZT!W�6����SM��?���R&8�+uE�7U���G�ǘ9�u�ȓ`�|����{�P(��O���ф�@�h)8�*��-�t�;"�FT�ȓMI��#*Q�D�6l�`G��l�ṙȓoς}�rh�)��4 �Q*	6�D��r�4�2k˓{7L�SShA���5D�`"�̦��1��>�@��]?�y�,�q����TT�๷bE�ybO�B�8t�r >ռmC��O��y�D�v�8�x���d�!�D&�y�$�6}=t�Qk�X�A$?�ybʚ�d#�e� ��+���BSF�yb�!����.O1v�"���B4�y��f��U&Vs�L�l�3s!���da��D���@�(�P�*�!�䓅i~~�R\(����t�b���"O��T��4<�<���n�:?��xr"O� 6����1P"5^q�"O��*�+�5}ځJv�R�I�x��'�1O�I��%r��ǐO�w�N)�y҅¨|F�)hVN�&� w�X��y�$��UxND+�#�P����g���y�΂I�@˶"�%F������\��y�䜬?V:P�T�;��p����y�L_5|>�[`O�1|rx�A\��y�F'A���3Aպq�<���-��=	�y��M����ف쒷 ?�7`� �y���?ä�KWǓ?�@�� ��ya��@�0��2	S�T�ԘH�f��y��8�L@j��G�pS��"�y��Q&	&t����E�.�fh��yre�R\j �U/P=x�p�l3�y��>!��ɚ�U�5̮R�.�y�^�1���q�S-\]`����Ҫ�?
�'��0C��!u��b��Z') a��'�Lq��I�j�P(@�]�'��Qc	�'[���VM&Q���f!�#�
�	�'�j�ڦH^'l�p��&e�@�i	�'��hرa��*�����D�a�]��'��yh� )��iI5o�4(�Jah�'�<d  ���X2㏬p.���'��q@�ߵ	��1@��R'��Ak�'y.���P�E�D X�NHH�a��'��=�	�hʆ�
�H5�AZ�'#�M��)��Y(���!F������'�t4�\�0h��ʖK�`����� �̫��?J<`���-X.�^H�"O.��7��5N����ģ	<"������Dփ]*az�ԁT��M�R��b���F�,�yR+F�8ߘ��a2y8�Ï%�yR�[�x��A!", y'|�����yҋ9�&�b�L�9]����×�y� C:i��)����!0=D5�����y�ۅ��i7�1���CW,P��y�*EO�~�H�%_�'.����0��'waz�C�F��t�I��h�d��b�yrA� l$�%J��^Ͼ��!��yrlOxc���Å�X�Ԡa�!�ybg�-Ji��h0�S9H�6  Q"��yҪ�0Ϧ�@N�G1�-��	J	�y"BJ/ W����� DL��y����yr���Z�s6���C���0!n�*�y���%5�R恹
e~؋�H��y�N8ܡrj�3�q�gC�y�a-Fa�R�2k,�ˀ��y�FB�t���S��:\��Y�5K�$�y����@�����1[ZlEk%*��y�G��(a$�Lq�(a5Dޔ�y��\>0#�I"��=�!�įD��y"���w��Ay�J@ 5���D�y�D7q�m�e�=+�(!`���yr L�Hꐥ���'�>9iS��y�DJTF�K�Nz�����y�6�,�F�
:<J�yZ��
��y�Ȗ�P�Lԛ���/��p3��#�y2X�#B��S�˺~�.�lH�y�K�l�U�v-�+}�
49��-�y򫘾E���aO�x�����yR���`�����m8vXkG�л�yRK�=_�	dC U���AJ �y�.>'��$��<�N� M��y��Ʀ*��	��I6���R��y��}���{��� /�$�*�n�!�y��E��ތ�%��)�tѩ��y�dӎW�05(��_�<pu��bX��y2%�>xm~�����,�:)ܹ�y�F�Q�bM�C(F�1������y2Q��tK�%�T00�/�y"*�g;���D��g�V������yh �'i�jl��Z�e�ǅڿ�y���5P.}GP�A���ʜ�yRbO���6l͙K�jA����yBI�)'�(�fIE�I��(��Ԧ�y�E���t��E��<Ub@��K��y���#��,�e��$bj,�DW�yƛ�|`���.*$͉5L���yrk�(@��y��RUXl����y�c�8ez,8�ǁ�R��X��e��y�G\� ( pB~'����k؇�y�X�r�l�H �=,���Z��ܹ�y���J$BpP���Y�L������y2�
��\�y�b�L�U;2�ß�y�ܬ8�Ƚ�W=f�1����y�%Q�� ��&��92��Jbo���y��N�2h�$0-��
�&�y�hşA�n��w�Q,�Be����yB��7~P�`��P�!+�@�+���y�J;R�{V���0S@nH��y�)�!z�0%Xc�W��zUHXh)�ȓ� ���_$%
�9 ���^%.\��S�? *ɒ3'�.6�ph��@�
��;E"OB�;�`�%%��J���1��X�`"O��C�	� J܁��n�uܒ��f"OBEI�-�!�����A)��as"O$(��ȝ�d�µ���\��Hp"O�t� �͖���R�kk�nQ�1"O�t`�L���Iۆ%
���p"O�4q�CO�V7��%$��{R"O�3�.�#`.���_�� a"O~p�$@"y��L�A�2}� h��"O�Pk��Z2H{*(�@�k�A:�"On� �A�	^�EY�N�Hn�zr"O��dE�x$�C�O^7�&(w"O$5c��H�M��K�����"O�xq���193��S.S'�،R���?LO�a���Y���Г�,WxY��iq"Ol9�AoP�{�j��w�PTRn`�"Op|��.�1 >�ä�@N^ѣ�"Oās��=Q A�U�ÎH�h��"O������/zvB��1g x�"Op�9�d�A5j�`�a�#Q�u�"Of��fs��ku�%q�0 CC"OP�`�GM:��X�͏[�v	�"O������!t�#!�A�'�t�ځ"O6���)5*I``a��h� ���"O�����T��)`Kq��=�B"OJ��tcSw�p��a�=a���"OzE�&�D�Qф�&�y#�"O|Eі��'�ਫ�!,
V�1&"O�� ˑ"eR��CGM8u(R"O�ʕ#ʰ qL!A'C;18 Z�"O|$�dm�.oa0\�lS���P�q"Oȉ�G�[j�u{0k��?��)
�"Oذ
7��,A��רIF��[�"OH=ȵD�Q�rY0�GE�CE�x"�"Oʵ���7@�\#�� �6%�0"O`�h5�� p!�@H�[���x"O���ȓ-@.�p�-�T���"O�\y�b�O58�yS"I�6���H�"O�R��z��UH��"a5� �2"O��۷l�<.Ԝ�"�ѮgL$��"Olՠd�Ô-�0\@�C��S��q"OJhWnN=Q&SR��Kt$Yj�"OP%Q��L�B!�É�SN�d�E"OJ}"#&�8������vA�!��"O4yR� �>{�*]�ԬH�ߦX`B"O��b�w�"��&L@�"��TR�"O�9��˺]�4���Ay�ra"O��rc��(�NQ�РԎ`ۺ��u"OH�����5UH����n��o:̉"OfՂ�C M4L��MU�~]X�"Ot��L�>(M�}�E�P��)'*O`� ���
���
�GA�n�Τ9�'�̫���sH�Pqd��}����'o�T�q(��B���j-	��|X
�'$|��6��
7�5{�e��ƕq"O�Dۅ��=(��P�d�Ke�y:q"O����.H�P�|���!�/d�^;�"O�A��F�1L�D��F�8��ҵ"O�0)pb�?�yH�L�,ň@��"O�y��+��b���SD��"���l4D��y,MP�D,Y6c�e~Ba''D�����'��c��3&�i0&D���B�#�"P��J٥_�R�C�6D�� ���E�5�@���$Q�)6\3 "O���E��B�)�Z7�qÔ"O:��x�b�����W�4�"O\y8į�##ti��U]�mi'"O���C)���L��Z�Oy���"O��� �Tظku ��t"OHt+�a�	t����'X�K9�)XQ"O���C��z��IJ��0H�hK"Oh=TO�=7�Ѫ�C]�W&�Б"O�ɀaO�*Y��$+b��6m:4�P"O�;���0�BY3/ĸ	���"O�8)��^<vtɖmY��� ��"O����$=��!h�Lݺ;а�p�"OT�IQ�Rڀ<1�K�\�����"O��˰k��-'hœp�Y�E �S"OfP2	��j�"�F�����"Oj5��.O$�ņ�(Bh�%"O���3mN�y�����Ɛ��kD"O���eO�a��mQ�H���ó"O�� �*�|�0[`ge<}��"O��K�d5j�k�#ZGJ@�p"Or����S�^ i���B(����"On�C�%�o���y�m5	-�u!�"O<QrD�ʧ2u ę�N�.H���A"Od�&��!c
��f�&e�ҝ��"O�JЁ�B�B�aG̬N���"O y� )��9�4����T=K�����"O0����r�h�B�I�J�j	��"O�) A�%Ĕ�a�[�a�쥠�"O>��V @�'T�����-{��3"OV<f�Ʒyd��F�P�୚�"OV��f'(BQl� Y:p�St"Oơ�w+DG�^�*��LޭY"O
ybF(�/j������0�� �"O8Qr�%F�xiaIMx^T���"Op����R�v�J,q�)9M!���"O:a���Z4��!bV�+���V"O��sѮܼZv�����?e��Ч"OJ5��(+1���!�^�W[�)BT"On���	R�(0+�Í�OJV���"O
���_3tN�Aj��ë=���"O�q�,d�����/~(����"O����܇+댤i ��x!�@�"O>m��灖w���b탁;o���%"Oz9�!B�&�\9��kW�+Sv!@�"O܁�,[�jAs­΁5��cW"O-��@Rxt�h���h���"O^�#TK&���A�1\ID��"O�\`+PD6�KG�ּ�NY�"O�q䌇~�8��r!�E�~�E"OĜ���$3�X� �h��ܚf"O������*1��Ͻ0���p"O���BK�B��v�N���0&"O ���,�/nN�h�5�&o�d��"O
Ks��mN"��5*C�T�sw"O����H�Q�8S��(eP�9��"OH)��P8�kq�$$$x�"OΜ*5A"�U�be�J
*�A�"O���a�����n>O6�Q�"O�qe��G�f=�6�.F�q�"O�V�� T>�4H�#'|�:""OD�;6�;ElaK@@�1�H��"Od`�ș>T���K�΀�P�t,��"O�|P�ӏV˰�hDM���8K�"O� ��B���Ss ����ƃ)�n��'"O"M���+h�r 
�U�Q�
= 0"On��5'Þu�pi�U�O�3�6�if"O6�9�����l5Pr���
��y�"OHIp0Y�3=H͉'�6d4i0"O|��gВ/D�����H.oq��{�"OF�� A��ai�*Y(N�
�2�"O(̫V̔ xW�����^�y�\�F"Oha�mD��*_�I�x"OJH #�T����`��2��4
"O����)vFQP���-Zr���"O���eM&W�V'f�8�ޅ��"O�u��#�0%�ck^�)L�-�c"OF�FJ�xY
�,33P���"O�58��Q�H(Q�Y�'5��G"O�|`���#l�.1cī�o@m�t"O��"�Gҧb�v:�+.G����"O�(�j�LD�Y��������"O-X`��Tk�'ލ��"O�T���,�x�a�
�e���"O:�S��OކH����n�(�"OH��Ŏ��0���M�*d��Ig"O���paܩD�*ܱ3m�G�#�"Of����(9Q��"&�L;hI<�I�"O"�c���[��m�+ә!7� ��"O
ph�!�.A���1�N!zrH��"O��IH
[԰��;lwz���"O����ӝar@)��n1iP�9�"O����kZ�e�h��P�O�Ye:�P�"O����1-����W([5��z�"O��R"=Ii֠IrC>*bF"O�	�P���R��A{�MƖK��3"O��zQZ&]nP��3��=j�-�3"O����g�f�Y�`�ۚ$�́�"O�t`�aY��F jŴl��"Oļ����u�6|���������`"O�͒����8�cbrF�$"Orm u��SyZ���.6�ȉ�"Oh���A��Q90��&�[�"O�ӧ��o���@pϔ�t��y"Or�0u�W?R�.=(�.�Y�P�i"O�����/��`�b��!l��"O��S���I "�&n��k	���"O����G�$s�P1!6�)�n<�W"O���/%8*@�*f�U�ڰ06"Ofu*R�̀w�̚��^�V����"O^l��/��6�= e��a��͋"O�lK���:��RTS�y�xm��"OZ�+rd	(H��@�F�G��Kc"O@t��nL&$�+ւ4��di�"O�й&H'ϔd��l�N,��"O@���,�1H�dp�%�\���i�w"OB@�Ǉ�!ld�R6���{Ef ��"O�Y��T�C�f�Q��L*#>iv"O�y�͇��a�%��:��Xr"O �i7 ۭ��`m��<�䐥"O�`#�c\�{dy����L���9Q"Odz��]�;;B�B�%i��Cr"O��E�N�*���ԫS R쨌3�"O�,S�g�>�|i�ʃo�f��u"O�	#2F%s©��	��8��	��"OLh��N�b\�y[@U�
���f"O�u3S��$I^F��@ ��r�y��"On�;#S"(�Z��!d����"O� x���ѝ�:T[�ݙt����"O��(��?����;|RekD"O2�#f Y�i+Ly���^IgJ�v"ODY�g�!!d:�b@��,e+�5�f"Om�iMREÅ�Rf#d��u"O��z�'΄m�҉���9� �Yg"O�U�M#*�.I�ހu�vT;S"O�Xa�5+ָ����!(�޹�r"OZ�!C꒬0��`r�,`����D"ONL��GS>%0L&�O�**�lb"O��bvn�t'v���آl+`�A6"O&H����$m�`�p��gZ!�B%5��@@����y"ĳ7H!�䌣#���cnC"{^f���`�K�!�D�
tؼ٘	S?|�Ҕq���x�!�$�"L�q���)�z�)M�@�!�$G<�F �ӊV@# yC���p!�d�CC� i�*�<������E!�$�E{V j���9�@����טS=!�:�!D�����}:Ŭ���!���[m
���/^$'��3٣c)!��<{�h�b��ϊ}��E�Ц�.,�!�+Y�b��!�`u �ɗc���!�$�8'����#�Έ{r��{� ݽ,6!����f�QG�s@����И2�!򤙦'�f5fC�9z՚�G��Wq!�D�(j����oЯ4*�!��@Hm!�͵D�
��%�/N#�tqc釒$c!�dXk�p��v��-�����@HP!�-2C���A
>k�v�:��r@!��R���s ސ/����U$!�����q	�,�C��Qc0��h!�d5��<S���*Q�@e�GC�q�!�dEj���ȳh�1�<"�J�!�$ y��	b������϶4�!��n�^�"��B3QV�q�O=Q�!�;�dA�b�۩%Nf(��M\�^�!����(dP��+k/J<ZT�N�!��ƈB�N]3e܌;� �r���$q!��;KBnA9��'�ꐪR��	M!�D@yᰀ	@B��~
���k
�[�!�ĉ�x��<!�l�f%���fj��?1!�$��m��R��?V�� /
�g�!򤑫Y��;�⍿ �V=�2ȓ#���$�X�2��%ؒEl,��Mݍ�y2�ɓ�J����[� J�@���y�HD
��ث�`��02$��Wᛣ�y"lS�S�V�)���)P��Q��X��y�ۑQs|�Ц,΁5�����"Y	�y��ĀE��\`�J	+��AX�l���y���-��D�iΗ$(��{����y�ሒ
�|<��*R9$�<*5,֯�yR̾��ʔ�1u���E���yB#ٍbr�P"eA�A��xu�,�y�o�"����KF�<�ҍbT&̞�y�bD4��뒩kM�l`5���y�E�/+h��{"�TYƸ8U���y�_�w�nM��D�?L����t&���y2����y�8��3��$5
4��'�T�j�F��7������&m����'�fz��3	8帢��T�p,��'UV� u�I��uQrΆ�R�VI��'s�`��Z�se$hx�	�`F�̓�'br��eؚ�$�QC
�p��q��� F�Y�eQ�!2l�`����:}b��"O�8���h\P�b��E�r�"O��SGYl�%����?r�Q"O<�+G�/�h9fdY,58��7"O ��ѯ� �*}��_�QD:$�"O��j��#�
�B���$JB��c"O�x��X��تv)��F�)p"O��sP6	
 h����W���1"O��s�$��'zT����1Ȳ�x"O|��ņCP�F8JE+���k"O����劤�օ�ꎷ}���"O�Ж�X�b�r���+�� �̩�"O�|RQ���V#\]A5�^G2����"O�L��cO��)�;󄸉�"O: �b�*'[�t����A;d��"O���&L��^����.켃3"O(�͈g��⧀T1>����"O|��M3E,Xz%BK)f�bk�"O�u�B��''�)#0ύ�I��LȂ*OM��a�g�@�@7���F|�a
�'�$PI#H��v���уʮCS�0��'��l(����h��!�?����'�*��RfU4v"p�2����1;�5�'��$M�n5� k��7��"�'U�M���K?,�������*B���'�<�@��B	1�%�W��`����'�X\J��+:���X6�Ÿ,b��
�'���[$NT���D%ݍm}z��'Y��1W�J5�؈���N!���a�'Y��Æ�3yC���U���y�'�\t�q"�6T)���	�"4��'��<�$p ��w�F2�Ru��'i�9&F��8��7�Qs�΁��'�4iE�0B��-B��N�k12�C�'%V�CVGY�s���'׌Zz�"�'U%ɣc���CA7;�=�'�:a����T!��C + �!c�'NRYGlQ1����M a��''� h$M��0e��C�!B�2�(
�'����(
�v`��S�&J� 
�'�mJ��E�6��A�K��e�]�	�'5��A%ȥUnj��`��g���A	�'F�Y��D5u�,}�G�o�!
�'*�6dV�q-�J�� ��6��';�M[�/��Yֆ˾x�6�C�'Lf�9���Y6.e9�k��MX4��'�p�&R�a^xa�Ή�zd��'nx(�V�n$X�����"MI�'���*�� Ʌ�"<D<��4���y��-Zu����ѾǮ��g����yr��(�P�Q�A�x
H� G��y	���"�Η) ��)����y<(�~����,t"�!� �y"4!�􅃂�{�Nt���Q��y"H׹y��� 2=#���i;�y�A^H%�Al�9��,�y�
݀���īS�014+��y"b���������[����y��N��9�Κ}�`A0�iL
�y#�F�{�,�� b2���6�yrd��}�d��R�@7m���p�*B�y���d�0��l	�.��*�*���y��N�P�ÔN >�n�W�_��yc_ {s<����+I���'�I��y
�  ���K�:���1��c�$�t"Om:`O�v�q͙��:��"Od��L�'O�P��ܞ 1�}� "O���&��1W�"pJ%U"'P�!ȣ"O���k��5�0�5�ܹ����"Ox�r4���ThA�3S�R�z6"O�
�.��R�	��;��8:#"O��cf]qj����L�����t"O��ņ:�l���� 1���X�"O��:����sF5S�_53+v��S"O"$����'}4�J��:�"O����m������5i&�r�"Ot�{bE:6�8��֢�`�Հc"O$����+3Kh�{�"ȆI��)E"O6�x1ٯX��ۇ��Jv�1��"O�@R�
���� ��1q��ȺV"O^�{�eN<n}�(jb���+"O�h*e&]Ȱ��2�ەu�}�"OF٨�)PC߆!�.��#��<a�"Oz�atC�_�i`#�K��R�B"O\�s�F&*�ɇ��R�6�3"O8��W�P:n>�R�@�;)���v"O�}���2��,��jC&|� 	"W"O‚�Lؐ�	jD��cc��5"O�z�O
�T�a�	 X*b|�"O:+�%���ɣ��"q��x�"O-�$'�J�H���e�p{$"O�QǠ��O��� b�ڰ-(ƕ*"O��x1-��n4t��T�a�`ܚ�"OT��)�Z�����<,K�h�"O$��5�
�P(�����|e���"O�@�tIС�°{U��+<8)��"O��a����`mh�W��,��"O��a��.4Ģ����7H(A"O���.�:�N����B�$-h!
g"O�i)�E�	;�C�ӉY�(� "O�va[)U���P���>zZ�"O��ig�@�@5jX�r3��
�"O���L^�$��5�	�h1`-�"O��8r��H1}����6�$�p�"O䈛!a_�C���rG��nޅ��"O8��V�5���sDcЉ3Y�Qz�"O&���ݱ�d�2"�G.TRV�S�"Ol �����5�`�:@��a?�I�0"O�#�虓d.�H�W�\)'�4:T"Ov=-)ZM�`�11��E�`d̯�y���Zx����m(���07�ٛ�y�JٯjNJ�a�"�4]��D��y��h�>��'��4N��P�%�ȩ�yү:��܋�`8IMnJ���yB��V�*x��H��:-� zD�6�yr.E&W�P���R����B#�Y��y2mZ��d�
�|nƑh#�ê�y���$u���pA�{躥��j��y�F[>`�+�;?}\m���W�t��B|ッS����0aV�q��ȓ5�b��mI̭	'�kX�ȓ9�@���;`����LN=�-��tƎ���ܞz6�x�i��h�NA���v�K7�I��(�E;pL}��l��}jС�){h)x�d�;�6Їȓ{�r�c�oYb�����ȓ�U��O3�������c��͇�]@�a�(�T��uA���8����S�? 2ѳ%�$���B���d<Q�"O��i���!R�x����>�0s"OD0�2�AX	����R� "O���A)��`��e7��R"O�g'ĜkU�p�&f�.vq��V"O�� b)�t0���Z6;_�P0�"O� )F�C1nVlc��F�lH�`��"OX�HI�)#t!��
C�U�m��"O<���(LodqC	�&Bn �"O�X�d-�$�1h���("\�iA"OTҵ@	b�|!��L@��	�"O\��˘2�|I��ʬ΢ĉ�"O@y�4Mϸ,����$��1� ���"OL9#GJC��͊sG��d%��"O�á��E�+ATd�姇�q�!�d�(d���IbO�W�|�����@�!�ĝ���\�W�COg$E㑄�=�!�䅅w�r�GB�Q�����W�N�!���,ֈ��DEԜ0@��;���"~�!��C7w4\���?JL��'�[w!�d�
��҈�5؆���e�8a!�D����ZXXY��FRrt��"O�)�lA�.�\�׌�	KP~�y�"O��r�(/H�0��� UO��#"Ob����� ��bk�.)����"O����-E��00e���W�^H��'F�A���H�E�XJ��IN!��'9�QH�##$����d�G�@�3�'�*����S� ,!4�M�<)��'����j��=�#!V?=1�\K�'515h�4���р��8^�"	�'����u�6I���*M6W��

�'Y�u	S	��-���W%ҢD@0l��'(�k��Ƨ)p4�eA&s�TM�'V�pw�h�H���AJ�V�L�Z�'%t蹶�D�����'�S(P@�'���W�:9R�p�uے�0�'��d�V-T��^8���=m��2�'���S��� 0�vBD�;3�T��'7��	ң �CfL`��e�!.��@��'0��A����\.�@Ѵh��P����'fzr���l�%��AʖJ����',��zu��X!� ��#!Y��)��'��F� kjX���ϽO�j���'M��'�*�J);A#ēB4|�C�'�j��4킥k;QR�M�C�����'� �4;p�h�"A׫FϮ��	�'2�&�CA�4�T�X+}* �	�'�����ݙY&�Ě��'R�iC	�'�x��&_�x"�ʿz�@ �	�'ӎ���:5:THש@'l���'^����'+)b�LUo�M��'�L�*c�D*e����UaYaQȡ�'���9��޽-�r4�ģ���p�'j�)Q�T�,�m�u�	�}_��ȓ|��:�e[�'�wb��򈘰7��,R��2���{(�ԇ�I0�t����(,k�!f�C!1�C�I
=�����F�L��#cH�8w��C�	�v�܈Q��[��%��\�	��C�I�B��@�m�3�l`'��%��C�I�a�2�Pug�^�tC���%�\C�	/~�ĥ!�/�.R�@��"#G�*C�	�_SX����5�<q���s�,C��	J�T=��'*Z���x�2C�)� (��ڡMo������.&Hf���"O��cd�"n�����SW2ۃ"O�m�S+�f�X��_4��lYa"OL5�T��	Z�q�AgD $ ��"O�|�$��EL��SLD�Y'"O�e���nK�!�)*���"O�u�r��@Z���gOZ$_<��ɷ"Ozؠr����$�*?���"O��� Y�a垘X��ܘ(.�Yr"Of��&�H( �#Mτ\R"O��k�!	�QU��G��aΈc3"O�)S�mgz� �^T��A"O�Y�%D�;ЖEW�жl�̬��"OJ�:���$<*�Yad��ӆ��"O�"1Ξ�A� C�߿?�V�`�ɑ8�L���E&ʧa5�0��c�;KĚ�XU
G0C���ȓ,��RM�3Q���1�CA�>�h�mZB骹[f*����S��M;0�[�+�.���K�0qg:��a�i�<�� ��%�,&[b!�1D�y?1�(ح+�h)�Rk�Ox�P;cg[�W��[�AК��� b�:�O� H�ĐPӦ���M�6�L�$f��Xp!Q�̈*i������ѧ�H#^2���H�c�rQ�?1PLۯ)6���3O��E�`�}��V�G��yʢ�мL�ƈ#�k�{�<�"��h� CY����4�ۋ$�&��"4n��Qa@i��D��'Bx٣Ȍ����R�U�xh��h�'z��"s#�;}TR�X�C�T̼�03�/35ʠ��E�
CU(��[�p<qȅ_��h�D�+HƕrҢ�ZX� m��U��cU�02��HC���/�����DԀ0>t��ǚ�)���f �z��7cq�u��"I&zfL�O�˒%œO���b̓[*���qܧ=�FC4W8~�|X"ݝ9����%􈓗끪M2(���M����jR�Ϻ|� ��������pOj�'���'��	�f`��$3��R�B���O���F��9(s��0���%��ؗ�
�Ō�,z��xJ�(����f�W8��C�	�@��E
u�[,����d0�'�m��I?j~��b���F���C�@׃���QfV�4���W�h|5�o�ؔ���S*;���"��{�L̖'��k� ��Um��Z�KZ�1�l���
;��O�nm�*\0c�	�"�������'X���@׸x �<hsB^s��yt%ۓj�����4%�y�l\��ħnF�J�,�c*�9	NQځDK2Sո(�
.�OȨ��̎+l� R��%^�X�䕽]�D�0�S�B�"l��oA�*MH����^8� ��+�q��ԫ�A	�/ELu�� �Z��mY�(�?l����$���4���%mG��TkʻG�.��A���BE�V
O�h���C�p���妘?��Dab�O��s��,1��ĉ�ː$N*y3��Wp��}�Wj뼈���6�2�!���Q�<�"Ʊ1|xŢb�!H��#!c�,_z(s'/\(L(Rd�=����F�hR$H~��Z�q]��6(�X���s�@1IO�~r�R�i��A�q(�"�<liUL]gq~	�����H��S��I(��V�Y�^��ɲ8_d��Q�>u�dG\�zQ�$�� 4U����a��O֡�_ֆ�ɒ	���l�����bƄO�f\��.}~�P���H���bəT�F�.������Ŀ@؈��
�=8P���ʜ���O��l( ��,��Q"S�Ӌ/�ƥ�
�'R�����_�:]���:����~���˵/�2��������'
f�O�X�Ɗ'[� W�� (R� �'&��m(}�zU#r"�$C�T�at��<��J��!!�]D˕�G�.��d��΀1w�%(%6�;��,pџ#Cf\����o���$�I�f0J̨qj�ET��cj!G2����E���H��Hh�֡�B�-7�h�'�|�ce �9^h��
ç&Թ�j?0��]�ʈ�6�Dt�ȓ]Q��h�'�*�&�34h@� �¹�e:�D��Yڍc��L>��T2�R�B�ձ[���G�]�<�d*Q���9م��.GTHڵ�U`�<	���ݡ�K�+%Y��sdD�c�<��M�x��0AH�3��A۶�K�<� 픷]+x�A#N�A�pKq#�y�<� .��5�P�D�~sA�^�֘q�"OZH�'��#kʈB�	�hB�{P"O ���Ԕ((���s��^O�a�e"O��a�Pŀ�B��/)� �"OFm�U�J�]e�(c$ �� xv"Ob��k�%lȖ:��'"O�Tx��@�s�8MÁ��a�±[�"OL=��N�1D ��B��s��4
�"O��yTh���7HQ/2p���"O�����й�n��-۳,���2"O�	P)�\<�ԉ��E�Z�4�"O�}!g
�u�`u�&@J�P�����"O�VR�`f�@���%J�6ᛖ"O��`�@ ��xio	ڈC"O���S#�	cM��x�H�.oTq)'"O�Rd�Xp�Q��I|� A"O8����5aU����,�k' �2"O��3 ��<P�a��:@�:��a"OJ8������M��k�L��A B"O��:7&W_����'@�ؑ��"OΘ��o�Ѳ��r��c7"O�[0	V2i�n$C#�:�j��"OxDH Eς/�N]��$Z&V沝��"O��B��_x�d����
b���p"O�M�`a��]+\�ɦ��[�ځ��"OL*H�6]l���C8 x��v"Or5���p-N	���G�^�e"O���f���%0��#!Z:|u�J%[��p���i�qOQ>��et,&�ňv�����*D�x+§�tC���$��vSh�%-&���!��`j:O�A��@�p�i�`X =��S2�'�X2w	Ϳ 3�8���.�,8@Q���\:`�1���ӦK�VU�eh�睉��%���2�>i��9��[�5}�c>�k�o�<J@� ���UKG�0D����4�9���C�5pu����Y���?0��궘>E�/�6I	6��BU2��:�P��y�dU�hJ�H�Q`��mh��3��	��	�1��'�(�ax��	�-aW���:�jéG3�p?���ϐY(\����"G��Ep�d�Qt%�"��'��C�	;a���E��Vh�(��^�q�֢>VA^{Qք�Q�&�S)��չDCHH�(�2&@��C�	�W����(B�]�x�wA�6����F��*� ����S�O-��Q/�>�Y��Mˢ4.�ؘ	�' � �HP<:� -��͞�E0� )�4��D��m�=�1'II�3�ɩT���6E�e�2Ęp��]�:B�I�U��D��L�5N�jq�cc�V��`��D?q�x�ʥR$m��-b�m��,�P�����p��ÌVFX��e�)��@��@u!���B��ܰ�i\�	�Ӏe���D{�� ,�D��v(���ON�]�&�q"O2��C��&Y�c �CA����iqў"~n5t����fETS첆�	�bLB�I�(K\��gOݺ����g�(/�D��p?�Tb^� ���ޜH�RxqG�Tq�<����. Xx�2��zL-Yd F�<�S�
�tb0�1'�oBjySNCXy��ż�=E���ׅ��q��\�!�R9j&�&�y��Ӕ"閴ᛡKP�`f(���7B;����6=�ax"������)����U�)��>�E�˩u�	��Ŏc}đɑ��z$��R��iX��!�g<�Oر�d숞/�QW�D?ʨ,���}��q&�
ʸ�Vb�_�	�;g���P�����QAA%��"�!��J�^���O=LE�\��o�*���K�<���I�h����D�"��Uzֈ��|s�uB�C��
�p���4D�� �8u"��v�`M�/ �J�;gjހR&]y����3��BP�U�p���	<��DX D�l�x,���\�l(����q����@<1�$��eC̥S��E �K9t�v9GJ�
X3�P*�}�Ȥ��S��JQ�#��=AJ`Gx2��n�����%Y���熅z���%a�m��� _���ŧP:W�C�	fZ�D�JգpX╪R�7h���x��%*�@jG���/\@`��oXK��y�X9�rH!ŵ��ҐM��yB�º7�����"5`��`��Z3&�cc
ɹ3*	����j\0�O�ў�Yg%S�	9(-���ml��L0�O:dC3@G-a����r	O2 �`�(��O���: ,��Hpc��4����DP?��t�¡L~�L�&+
���Y!�_�t-@@IEF��$�f-^��dN�c�|�ҍ[(
ͺg�y��S�4���h��Բ&/NtI�
W!L8�cc�X�CSTB��@�zJ��s��Yb��.K��{�HB�T�P�6/?D��o�>�@�[�)T�s[�0#"ě�)����T8f�P�c���&J��~�'KN]�G#G�a%��@�C�+o`)P�~����@��V]�yp&Lά�P�0���G�J�hE�c���
�!+�O��*�� ��E��5͒p��Ɛ��(O��fט/�D�7ɔx�ϟ��k�iM�X~0��d�ݸ"Oέ��)/�8�W�On�� ┵i�p0�%��=�d�Y���E��"n�	��ȫEd(]��� ��;"e�C�	�3�@eّgҹ"���k���}s��*��'x"�3?���wG�~Fz҉B#+a^�`���d����������>���D"_� $�B��2j[p+[��`ʷcU�Q $��E �Oΰ�g)B��3��V�cIlɰ��I�*s��:,�8r�1� =��ŭi�T�P2j
9*�"O���FO��s˺�+��ήV�u�[�(�&�P";�qOQ>�3A��6jY`XG�H�H�3�o/D��T'COXv�P�-�/>���M*D�����_�-x2G�[+�A*�`.D���oڼE7�	yUΘ�[�)¶�)D�<	Wj�OK�Xi�! *p��a���'D��{s���f�N�@EB�P�����)D��c�D�r�Wl������(%D��PEb��9�HA���s&�y�#%D�X˭;Y
��T�<d��ia"D��zGI4sh��M�>z� I3�-D�L�A
��iG�'i�����"+D�R e��g��ݚG	!N��;��*D���G��1sҰH���)�Ģ"D���Ɩ�k�nЃ�/@��ҁ�bl!D�<��E�'Gfp󄋕�v(�AE=D�(�'Ō,d�A���T#@J|"�%;D�DJS˕�Q:j�b'�	��)1��8D���C6D�0�"�Q ��4�8D������gtʱ���L7_��Q[�8D�T
���_Z���.��YBV4D���V*�$�v���A��g|�:�J2D����τm����)���`��2D�Dps'�(N��qrT�4u�+A�.D��;��?XQ��8��ǖ�<hA��,D��
�+ބg��55�X�a=|Z�a(D���T��ks(�wg�	b,My��;D���P%:$�i/[�Ma��&�<D���d��B���96�۳�\a�(&D�����Gn���oCvP�;D�p�0�M�.AvHAR΃�h����*D����c6���`^�t2�9��"?D��"�O.��]��������:D��Q3%��uY��1�Eّ'jJ�ض+8D�� �LBC@�bo�=U����6�4D��cm�J�����s��\2&"3D�Tڧ �nN�� �"u���[��0D����ߝ\l�a���~��p��3D�� �E���,�tx��
P��R"Ot�	�b*~�`��V0ވ��"O�5F��Q�����C%��;1"O�����
	" ��%���Y�t"O�( �_�틔���\�L��e"O���Í�'*#z�I������"O�,�DiL6]Zn���*���"O�pPE�R.y�"�p���#y�4"O��7O�.sz�q�K�+v�j��"O~���)C.\#
E2w�^�(s"O�Q���M��t�s#!zh���"Or@���ɮz�hف�^�bU~Ԫ"O�Ԓ����騦c�32�T���"OĒ�W>-%X��U"�o4Fe@"O�uQL�#zf���!�6΄\�C"O�y�B��L���2��E��I"O�L:�m�-�6H��Ǐn����"O$t�d��[]&Ł6-��=�Y��"O-#\�#Y&����2gZ�`X0퉈C�����(�'7�l�3�`K�t+����k����AB0P����P��h��߻$���l��KJEV����S��M� ��G��Ə�fa��2��O�<�ōG<'V�6�	9P%B�2��p?)�*P�bHęQ�Ax�`�E��}�r�×BY?3!��d�9�O��)�@Ԥ �>̒���|{&-z�����6��-�,��U�]�'��'�Y��ޅ`���?� l�S�"���Oϊ J.�}��H��������ޚk�b�R'b�<����c�iK�s�;���Z%t�Q!(ѳ3����p�TF��'q����(�&0�1��*����'�T(P��r�;p�M�]:�y2�ldb�Y�@�;��Ȑգ�&�p<��84D��d}�f�8`�r��$HP�  ��-ȳu��ٲ�H� ;���vH�@��!���E����)���Rd�;�0�S�%  	��asc"}��K�|i�f��E	�>|"}���+��E��A�r�Ȭg��#Gw�BC�I.|��Pt�K6Z�ڍ{�C�Y�,�ʷ��CH�P��N�9$�6袕)2�S8&��5���5b� ����ŀ�u��	'4���0 e@�yw����
�OTX�A��F%Y����;l|�L����'�l����u�z��wD:=�\�P�9�џ|���x���+�'��=�.RBc\&p�����ݝ:݊Tk'L�+
�1��?��3�G�=��K"��u��0Ʈ�<�G��	Pu�A��cY8T�8�A N2y�Z��}�1���<�
�۪2�v��s��B�<��ۛG.�Cӧ�Zp�HeC�<zᤁ��C�2v̝�%G 	Q;J�'>��@��R�t����Oմ7kveB!^�Qy�~THv*�I�Ń�J���P$ίc&~��wGKW"D��I�J��R��
zs���dA�1����Ň4��l@��UlQ��C_�oSjL8���C�](5ƀ(5��pA k��Ag�OlZgn��Px���{��9:�iՓ>���6���~ROQ�N�����%�3.���{&�>\�����)�S#;1e�N� V��#�G܆(�C䉋.VԺEI�I:�*�^V����r�.]����t��!$C��E�*���@L��'�&����	��9mY�er��F�P�T���0�l���*\%ָ�AhȺz�r)�|��y���
1������'�Z`��D(=,��#�g��aH���Of����tp�<�����J|��K�� t��l	H�Za@�!{(����p't�KB��>Z����P�U=���J���b�W$J���9=�9���-��O�P�dC����1�`��m�y�'�̀їO]iU\q�� �.)�W��~���6EU�L�)�P�Ӏ��ӫ"*��O4�)��2"A
|ȇ���Yb���'�xb#�O9
�w ��[!��ᰅ~~����N�+yh8�U�˙X���$[�3$��J�N�?}��p���]E(џ��V�:~�������wO��F�	f<t�K5��t��Q��W�����ȓv�M�q,ƣQ>�#�( �cRf��'��pHfQnâ���'(��+W�d��)we�b4~���l���#Uk;}�l$i��]�{�H��Fk.�$[�	�򙀏�L>)��U
<�r /�$
��H�{�<� ��h����L�Bu0����_R*e8�"OXb�M��:����#���>Ԡ`"O*�0Չ��J�挳�̔�M��h�e"O`Ks��i@lx�J��9|��b3"O�$���Z"VΞIrAiO�Q `�r"O �����+(e���D��i�"Omz�M'>K����B�����"O�)���g�4�j%f�8h���"O����E0%
����f��G�DD�"O<M0բT�C;���@�N29�	q�"O́4m�N�:m�)x���S�"O�X��+�"Y���lQ>�z@�"O�����|�6������ec"O ȣ!nƫX-8��AMp���"O �	W��xF����'�9bL�V"O��.
�[��0ȞAV�zR"O}��_������
5���"O^��N�D&4� ���,/ʁʳ"Of��#O��^��1�p-��N)�\�"Oژ�r�?�����͡'�x��"O�`�v�Йs�����2�<#"O uS���iL��w��5
�"O�ɰdǘ5-��4z�cB�7�H��"OJ�C�ⒿU�5���̇s�p�"O~� ���FH(�"��>R�DEx�"O����
si����C)V��Ś%"O�(ʤ K�`YJ��Gɹ���{G"O��kщ��B]�J�
�<�S"O�����ݘd"�Iݗa��� "O���Ǡ̪T]�ɇ-�<
(���"O.¦CّX\U3����,4R�"O�L�Т�&|�ō��U"OFe�S?7�P4 L�5�T�0"O\��$��eZ�,��ma@9�t"O���SB�
=6f8���A$�(��0"OfU�q�iobȪ�IG�J@�<�A"O�C&�-�� ꥩ�/@/��E"O|i{���J�l
�m������"O"�� E��x�Pś�i�f]`"O��賄V�#18{7��)ԂY�g"OVp��$�"2I���_$m�(��@"O�Ȕ��"4X��",R�Y�""O4"�.���^:Q@�"O�|q��͐6�
�rV�ī�>x��"O���Sτ�Jv�D�\ Gb�"O�  �Gl�Z 5"�����X!�yB��N��RT�^5�A�Eí�y��Ⱥ��P.d \(p#���yB���P ����@� �Հ��ݲ�y�� V��� 4r���ˁ���y�".2̂�jS�	ut�Ty�Œ�y���Q�����ˠbY�� �M�y� �)ڔ���@I0nJt���y�nԞ]v���K�\t��)�d��y�K1�~���#W�B���b8�y2�,U��$07HکN�����։�y��C�_��չ$�2N�2tA0g[/�y"A�����K�A�� �Gn�-�y���zW���WĪK.����NB9�y��fAz��2��I�(aٳIP��y"0+{^Qv WD��)8t�G��yb�0o<T	P5A�;e(�¬��y�����DI�C\�3(l�`a�G�y򁔥y;zx�FHI3�D��B]�y
� �Hէ���مa��4�>��"O�4�H�i�xZai�1j�T!�"O�Ra$Z�9�9Ag�78H��"O�e�g�e ^=�7'̹�l\�R"O��:��y����h	[w6�bb"O|�c0'�Xl
��A���0���"O����FV��=:�c�5`�>�*�"O���풦V��0�o�j���!"O�5��ԝW��)5��6̄mõ"O,�2��kl.���� e�zAU"O&��3�W�C_�*se�Qda��"OTt�S�_?
[j@(e�?(]�� "ONs�⍩JE��I�kL���#"O�!�eIʗJ�qS�W�V����G"O
���� ���)�+�eJ�"O8�C�$�Xl����P#78��"O~��s��Ds�,0�F��>+`B�"OX��服0E�D�u��Y�F"O��A��.�iX��b`1��"O��k$��:7*H��S&ʹI�"d�"O�� ��־SL�;�䌃-.5�f"O�	�©e�jE�EL���ys"O`m��(��Q�4l��(��"O�P�F#��z��R �0o�>�S5"O��Q�G�)L�ɠӠ�z�����"ON@b���q���N:+��䂥"O��Ҥ@� l��a���X�i��"O����ȊlC��+���v{T��D"O��8���M�H9��@� z���"�"O��pp��4Av��-�^G}c�"O�H� !ޅ��D�k��͉h@!�S�W���"�u��p2M�>7�!�K�@��5��]R���D���!���?3N�k��
	j�p�;R�$�!�Z�z�K&&��'�f� a`��+�!���}�L:����%y"y����>�!��ݜS�Rd2�n�8o�%B�冿q!�U&L�� ��^Hh<@; FQ!�d	I���;���IZY� �\;\!�d\Mt\� n��,\z�`AJ��mM!�:ή�4�J=�|T�fi˪4$!�ߦ� L�5�W*1^!�Ҋ�
D.!��@�~i�y��0?p�kҩ��r�!�D<'c�*�J�\�*W�!�D)I��Ѱ��Q.�yʳ���!�K�%}�qRB^�9 lH�D,�u!�ḏ�(��OP���`��mW-=�!򄓿G�N ȱ�g�ȍ:�K�1r�!� !��[���1��3ʔ%n�!��ޜ
���fRb�\���ď �!�L��>�ᚙ&��@ráF�?�!�:N�����N��	C�`��l�!�DH�]��ɚ�@F�X��1�&�!򄊦p�ԝ�e��d��I�.��3�!�#
8 u�7�[�~���b�,h!��<=��Bd�_�p������!��#U�P�e/^�[x����M��7�!��z��Xc�CF-N<p�C�%�!�F3��=[� ��F�����P�!�$�wj�m���S��������a�!��	3?z��ÏF1՚�Q7�	�7u!���Po��k��O��1��v!�d��L<�t�ݾnz�P�N	�b!��4F�$��VT8Eb׍,o7"};�$��&~F\�e��q�az
� �	K�!��vp��B�Mo�H|�"O&��Ţ��h��5;"l9�:�ِ"O�Xq eּ5����JS�H�0�x"O*���J,S���3U�ȟ[��4���'�� *�(K�P���h�)���07�!D���vl�(������ 7V��+D��� *\���%0y[LQ��h(D�j���tr�<MS&V�(�ru�8D��A��=P̈	#�C\ ��i$�"D�$����b�~t�'���V�s��+D� �k�?o�dh0P�L�� �� (D��Ve¸PuDH����/F<Ⱥ(D�0q��z-��r�qj2̘�$'D��x!�	*J�eC��I���W"D����FC>t" ���똝v�ڹ���m��l�����$x�����e9f�t�r�И�nHFy�Ƥ�ȟ�xx5�ߥ(�Z��w/�G
� �U��т4	Q��O�y1����0�4��&A����dZI<q�m�p���O"�`���D:q	�,���z�OF!J��i>u�=	Tϋ�M> �0`aB�G}�y�J ̦}9��Gd�S�O�I�cO?<Q�5�
��5���0�2a�$#� s�� Qg	�S攤��^0��'x�ԇ��]����1n��@�n,� �-�0B�ɦ��� �J(?�^��g"�R8B�	�4Ԋّ`��,(|:8���#D�4�E�xQfx:��=o��\�0�(D��y���EiJ���/�,�(�#D;D�,��^#U��-� �H�VXX�4D��g��(*햙�Z�p����<D�p�"ƴg���ؤ��7�hT1gf<D�xF�Z_bL�06ȉ�:>�;(0D����,�2�� +P��85 .D�T����:D����?SLDY�+D�X�2b\,P�h��) �s�
|���%D�����	8R���F���m@ƈ%D����gʵ��i�Ϛ:35�9�#�#D�<��
�e��٢e�ؽ`�\��U�-D�8��*��	, Xq�T <+j�J��,D�� O���"Q�R	1�NM#��/D�|z�����dU?0�Fi��	-D�d*�΄)DL��i�쭡�m*D�4$�F$!9��A���0|��ꐬ(D���h�rc� �4Iׄk�Dٺ��)D�$���֪a����Q@T�ME�u�<D���!�=3�<��c�S�(���(��;D�lҷ(]�~�[B�Q�v�Ƅ��;D�h��# �)D�ͪ1�T}x��	9D�Ē��/`�V�re
q�r�:��3D�hx
_1�Ui�^�fl�נ?D������6U	�<�Ce�"�e;U<D�P���L�)l�U`BZ==�`��,D�p;@F���I��yݼ 3֤(D�ءw�I �z�JF��
~�cQ&D��`үư��qᦊ�,ij8�F�7D��3FM=D�Vę%#H�Y��F�!D�b�"�^ @!��x�գ2D��� �^�5ڐd�4�K� ���2D��ڑ*��J�ST��<v� ���0D���%��D��@&���fC2L�YHB�	 S��v��m��yIE#�"_�XB䉝@�`3gA��|j��h��/�:B�N���I�K���B3"�7\[DB�ɻ#n����n@���A
��jB�IE��H��A)]>~e�c��)i�bB�)� |�1���/M�02�U<o�� 1!"O�i+g�@�Wy�%JA ��NZA�U"O�|KCc�D������XϠh��"OJH�B��S�ɑt^Ɖ±"O�XRi��L�i�1�Γ~K({r"O��ptA�c��PY�O�6��Q�"OH���FKA���a،1Ĥ�"O��L�,U⨑1A�WϘE{�"O�,���zc�e�o��0��"O�uY�K�f�q�MK|<�A"O���aeB y �%@w��B=�U�D"O�lRt�K!tp�+'��2,��E"O48��7^ѲЪ�\�{Aαr4"O&��f�#��A;����\+>$�"O�qIDe�2^G�e�3�	�,��%j�"OD�G�ٱ\��9p��ل;�|L�"OFu`D"ۜX��u�� ��p�@�"O@l�B������b�:%z�"OD%�$S�\�CA�'��UI�"O���t-�ko���@�>L�P��B"O�8���T�Au�T�D��T��@6"O���w�Jq׆h�*x��� "O,�"�拉m�R��c�Иrj�HI�"OD�I���OWpQA��4VH�k�"OV�H0��L�Q�nH0�`�"O�I9�"�on��@�W�H���"O�܊�aߎ3�ĤX���( � �R"O�c6I�Wۨ���Y����"O����`D(
�j�Ow���"OL�HbVkj�P�!˜�+bj݋�"O��4��hh�`"�'|�=��"Od�
��a��5�.$~TAq6"O��I��a����L�{F���"O2 �FEQ<_�,3�k�tP���"O���F虂2ܹzBꇐQ��d*�"Of����V1U��@�H��ܦm� "O��2� �-����l�'hs6���"Oa��ǅbD�t���<*Q"O@�!��<� M2%��7@���t"O�zR*�M{�|S�ύ�����"On�c���,��"����	6�y{�"OXLAdӭ~rmՈJ� $~<��"O�T�rb7U�H�S���Ek�E�"O8P�P���,k`��%�� �>Yx�"OtٺA�6w�t��öx¤��@"O��W�I�rʪ}!%g���K1"OVU�0IK�Yt��@�v�n\�"O�ʡEI�G;��3ѧ�l�@U��"O��A��4*1��iQG�iy,x:�"Oάِł�6n�� �l�/�f�B"O���D�E�+�.��Ŏ�#�,䡂"O�ՠ��ǆ<�� �K,!��9p�"ON��4�ز	��E3uD�V��qA"O″�H 9 �De[���^~$X��"OP�pc-�+�)��T�f����"Oq7g[s�L�#G�,JM��"OB�QR��DR�¢`R2�hl["OV`!��V��^]F�4��9 "ONL�(�}q��'�:<�>e  "O�[m�m�
����֎s�$I1"O�����M�*\�x��(We&���"OJU��⒏a�<:�ảw�¡�v"O~�P����r<K�ނ2(<h1"O� �Of�tb&��'�V<�5"O� �8(�՗\e�uÒ!��<�P"O�q���;��2���5��Ų"OΙ��g�znF���D<��r!"O&������~^�A��R>��"Oҭh�Μ|B8X��M6~h�Q"Or�c4#�%$��ئ���3�$,\O�E2�]7\�t���c����P"O(	Q��_-k�r]���aϚ<�"Onxi���RdP�a��.Ĭ��s"Oܽ��K� Ú�P��^�� l�"Oh)�1��f�Ii���p�� "O
<z�v�v)����!L�>L�1"O��Q��N�K�؅�g�<u���+�"O���$�ֱF����L6T�Q"O��R�5LX0�	,�~4ɀ"O���s��0��1ZD��"O& �u,
�3V��^$�$BQ"O�l1W\����Z�%��#"O1҇%��p`bIsF@T~��:6"O`�[��A22�H-3"N�X�t}8!"O4)�Wbǭ5��9p3-��[!��z�"O�du�ڠePL�1K�q�p��"O}KE#�_ )��i� ��lj�"O�u�VH��fn�$Pb��8$nNкA"O�<�OMbh��G�
�Y����"O���	��I��#�){S:���"O�x�'ƕ(13��x�Â/,�1"Ovd�'e˃[Zv(YD�ӃV����"O��@2�G
Px*	 ��Wz���"O8Q����9^YF�Y�l�-|o2��"O�ĈƄ@U�lBt邤KG�<�d*O������	2P"0x��� �d�[	�'��y  �'4�
��ً �~�)	�'��i$��x ��F)��$Y�'�A�M�{�qbB�ĕԈ5�'��)c��-M,9��-J�M�T�'b�l (�%�Pe)�B���'��<�c�>����T(��`�' ���)�40(�` ��F���}"	�'�
��Ӈ-q�)4�K�C�	�'��̫��ǹn"@z�B�u- ���'}�84�2�1�W��:*�1B:D�X��L�	z�e��:u��}y�M6D��a�f�E4.T��+�y"�M1D�4s�+�!HT��!��Gz��F�0D���$�#S��EJ4���a{D�JA�0D�����wUu��^p��"dG-D�< ",��}@�SQ�\���ٗ�+D�8�d	,Z�T�f��^� ��)D�+'¬-a�f�dB��&D���s��,?H0kG Q�c�$�rd#D���� "]�6M�	wV�B��?D��S��̘��`"��<��q��=D�`s@	=������۟����Bn:D�,���.h�u�7�+2LH!�TF<D�xI�.� �����D3;�:��/D��{o�>BU�tA!��<�.�R�,D��5��X��Q��]?,�"q�b�'D��h�COMf��s�bQ�{;@A�E'D��[E��&FȘ�xe�Q%�@�Y�"$D�� �b�%�|	c-��Di@	
��"D��zVo�?u�$2�g��9��[k;D�@#�?X��!��$[ZrԜ��O.D��s��W�҈�W蘀>��!�D2D�� ���jтB�`jgK��A��X��"OR���E�v9�t3b��j/���"O�8���Jjf| ׆�1F|p"Ol��k�*>�����3'�K��y�x�0Pڥ�DKZP" �Q�y���h6���V�s���p��S��y�*9axhl�c�άf{\��5�ت�y2Es��5��]��ya�&]��y2(��8�`���ËYg�J�W/�y� �j�>W�f��FL��y2�K�5��	!{�X�(����y2��t�X�+�k	
Eh������y2&�#c��b�(��-��9����y��ǯG��B��R|� �{���yB�Y��ܐ��I�Ę��NA��y�e�8N�-�5�9DF��3�(��y2	)f%��Ö�h�`u�7���y�g@1Y��b�%�,%��f�Yz!�$Pb.07�M�#7�,[�.�;v`!��D$,�A˕��J7���An�\>!�
1X� U��8	-KPj�~1
�'w�T��֝~���A`F�^�&�s	�'PY�1�5NڥRP��*:d�3�'5���T^<4��b'�8Q[25��'�܈� ��(r��@R��Ķ�
�'���!�6K��aO�\�}��'s�T`5���(�ANSVx����'¹�U;k����Qc˱<]����'��bE��^�@�	��8�>�q�'�$��  ���   �  J  �    �*   6  ]A  �L  XX  �c  o  �z  f�  �  ��  8�  }�  ˥  �  X�  ��  ��  �  ��  �  h�  ��  ��  ��  @�  ��  ��  � M �  [& �, �5 >> �D 1K tQ *W  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(��	M�O�
%�VϜ�8�qA"�@�!~�y�'Ƽ�G�h'��J��-��)z�'
>%'�ۂD@V�A�%�ZT��'��YE�KQ���E��.Ru��'��iS��*! z��QmE7�T���'Z���`Z8&�!t�4�>x:
�'`^��0��8�^DAŲ(��$��'|��@"`�����A�"��B�'K�I��GŨ7	�Q��Q!箸��'&���']�TQ�`G�,c�H��'���z7�5Me�X�ub� ]R$�{N<��'��)ɥ�M!u#b�{Ec�%>V���"��;{�,|��k�>0���1�Q�!��(�yr.ڄM�`����@�!�Ĕ7w5�yU��"Ip��CQmPL�!�Ү�����kd��e,B�w���[��(�� �E��o�{�4�6&������"O$��6���\�������TV�h��	�s@	)�D�8�X�a��%Jˬ��D LyB�6Pp��c�1����5�y�N��!K'�� sF; 	
/�yR�)2��Y�f�9)�ZD�Ǡ��y"��YӔ�X�P50�$ළE��y�keiظRa^(2��XV����y�Zj�b-Bp�� x6ѡ��'�y�'�~c�=�����1:��V��y�(�%-l,���h
�6@UIÏ���yr(\�cx�� M(ci����ǔ��yb藽;���2Q�K
X��<�����y���1V���f�V*:���&���ў"~Γ`�$���*�Eo^ݲ@�F.j����?�a1�Cr
���``Մ�<�j������]$erh��z�ل�fF���ӕf��a���0�.Մ�/����a٨��(G�ִ��ȓ$�rT,��� ��ڽ��M�ȓG	���J�>E�Y9!�4t�Z��ȓ~M�E�3B`�z3�^:�-���I?!g�_
J�e �-1|�S�Ƒ�<�(�5��D	�ˁ�pؼa"K|�<i@�N{�ȑ�
@��}�F�S�<���]���a®]�m.�%a�/�K�<�&N�a��d���H�B�V�h5�TD�<IW�ămt�T`�g٨k*�B ��Z�<A0+Ο/��*� )�H���YO�<Ѵ��v�*��}�8!�Q�<��h@�I�X�ZQ(P"Ӫ�� �x�<�&-��-��!� 2�ȅ8�-m�<I��4\��Dc6��Ȳ|�',�^�<1��
3�� .3'��h��BY�<�A�ϼ���tb�^����`�<�ݘ���ã�ּ |����a�<u ��0�QY�b��ub�
�&K\�<a&�>b�@�q2t�p(�7m�V�<�Q��{x,�4�:"�bz��]P�<�h��N�^�*�ط6G�1�c�R�<	��W�X�lu���1n!��QH�b�<	�oȺ8��-H��G�<���g�ND�<�S���CA�q�.��o����WjJA�<q��]�t��-���@�{z��;��<a�hA�沍д�:3�����YV�<A�"�9$��� �ס@W���G��X�<�3 �g�*����96��z�T�<	3ʌ$�麐��2Old䲓*z�<���'�~��/�#��M&!�o�<i�_0g��b'��4m@�����r�<�AөY����J�7a�
`����m�<!��̹I�a�)Ty���K"T��h� �v��:P,M�k莩�Ch7D���sd�-�(��Cü4D�D���[�u'T,�p#/�Rly�m1D�`:a"uM^��t,:E����'J;D���-�a�X�abĘ7O�����C>D���ʀ(50l<P7�@m$�j�!(D�,�g���(\�@�ݓ��u�!D�ı����*�)s⚐E�f��� D���P�o?~t��Č�W�&��@J#D��X!%��5��8Ұ���̨�!D�Ԁ�C�)c�P���#�#���34D����u�d1�D���Be���'D�� �,+6hN�V̤r�D�'vZN9P�"O��a�V阵��"N"T�`#"O��"��W��6�R�`�C̨b�"O��i&�1OL��/D_&��"O���M�^W�����*��I1�'���'���'��^>Q�	ȟ����S�2 [�LH�D̮bJ�5}�������`�	��L��ޟH��ğ��	����I�:����ǁ�JO�[�*�#F�r<���l����P��ğ0������	��I�s�l	爦j��P�p��*/?x��	џ��㟸�������͟�I蟐��k}&�{5��o��ܫb�֏thl�����	������l�IΟ�I͟8�	$Q@U(&�ĵN�"Q�Ef�7x�Tu�	� ��ӟl������	��\��2ZG$Y�PB1=@���¨S���d�Iʟ��I��P�	П�����`��Ɵ4��	O�yX ��U�Q������Q�I�����ӟ���ԟ��͟��ޟ��Ia�[��*r�����cɟI2����8�	�0��ܟ���<������4-H]S�GI�||�3�#l#��	�����$�	�4��۟���ោ���L��Y�!Z	]z;�&Nd��Iӟ`����t��� ��ğ���䟘��:�JI�6�ރ0�p��ƙ�IßH��ǟ\�I؟ �IƟH�	柰�� ����ό�F�P��b'�~Hd���ϟ���ԟ��	ޟ��	͟X��4�?��~R��z��I=*Z�ڣ�]x���0U����Ry���O8oZ�N���` NK�+;���5��D�*� �;?I �i��O�9O���ǫ�qk�@�AR&%��O����D�O⌒��z�����Da�.�O�u ĎO�X�P(�d��3�v�Z�y��'��I{�O�Z�y!�^�y��q�� 6��ew-r�0'��1�S��M�;_��rC�l��FL��~������?i�'��)擺f�`�n�<��'�&d>#f@�7dc�K��<!�'����hO���O`Y���V8�B��a�8�>O|˓��sܛ�����'q�X�����s�/��,Ѫ���D�U}�'��>O��D!dĩ���2P ���-tT�'hb!��  ��d�ן$ ��'R�3���/6ܰA���T ��!�5U�t�'���9Oz��1+Y!n��rc�S��̺�<O �nڸNl�K���4�D� NX1V�N���A9���"<O���O^��H���6m2?�O���)��j����g�� c^��ahA1�`��N>�)O�)�O����OX���OxJ�(!4�37oo"������<6�i��A��'C��'���V>牘W�`�K��g%�i�S�H1�%S�O�o��M�3�x�O��t�Oa�̪@ ��C�-���K�b�z<�����7L��S�'4��*��Ǥ?��xӴ�%���-O���w��Vm*�ݽ��`���O|���O����O��<ɴ�i�)ӂ�'E���1�&�b�QBR�r��{A�'�f7-3��������4#D��� /�>P��F·E����FL�1Y�6`[`�i��R��8#KK^>-�to�O��i��g�>�#uX�����3_��
�	W���$�O��$�O���O��$2��N��|���q���I��;^�N��I�p�	��M��g��|���=��ƒ|�m�*���dDY�(�{�
I+F��O�Unڻ�M�'�i2ش���1/��8�T��'R����&��+~���5��#�?qU��<��i~�i>Q�	̟<��7M� ��%%ݦT�еrUe�=�D�I�@�'Fd6-�]>���OB�d�|�7B��.u���64f�� h@]~��<��M���|*�<$��c@P��а
�#fF��A��CR8P������u���hЖQ��p�քZ�n�5S��aR�!E#'��L�	����	�� �)�Sjy��{�r);�"���0�H,lн�R$Q�P����O��nZ{�%��Iҟ���b0k�]�Ђ�m��%�b��4
ش	��
۴�y;��P7l�?���O�E�g�_�D�D@�񪆜4���Ԧ��'4�'���'lb�'���ԑ�F�v�d����ߢH�$���4.%����?9���䧾?!��y���e.�Y�L�%c�I$g�%l�7͕��9KH<�|��4�Mۛ'd�� @b� :ք�E䏉(���'#TI�3@韰�^��X�4��4���$E ~�%�k�����x�a��2����O����O˓v��f`X�T\r�'hBM��-v�C����@k��4��O���'���'�O^Ip���47���aŤ9p�4O���È	J�zW��r?�	�u˗������'�8�$��~�T���IdO��h�'��'���'��>��ɰ6hZ� �"P�X�:�M�9Hl�<�I��M�D�X�?9�4n���4��(ir����.4���<rvUB��O���q�t�o�5}��l�q~��^
9�(5�ӑ[�1ӥ/�&:�
dɦ��-x�]2�Q��#ش��4�����O�d�O^��ۨ[.�m��D�9�j�BC\ S�(�>�V!��Z�r�'�Ғ�d�'"�-��E�3�t%�5�޵Q%
u��h�>���iS�7�a�i>9��?�"�G�'A��y�e�߂�2|
���H�3A�&�g�����%�O`M�.O��oZdy­D�E�6�Q�כEYP�����("���'�r�'�O����M#0�P�?��9r�6Qy���"r���7���?��i��O���'�.6�ܦq۴86�jt��*5
��i�����A�4�ڼ�M۞'��� en(����������{�? �T ��L<��di�F̢]�Z��Q0O���Ov�D�O��Ol�?��f�1����GGN�a���&�KΟ��I�����4)��x�)O��oZi�	�
�L� �'�C�	�3�$NP)'����՟ �	�Y��l��<��O�L�+W�֩e!��s �M�i!jHYeh�sB�b�m�|yr�'e��'�B�&|�[��",(hK�쀴:8�'�剥�MC��Z>�?����?A.���8V� 9�� ��������h�O\���O��O��2q���Q*Ō��(���ɡ �&�+��O3>?$�oI~�O�������]2hAr��,���آ�֎������?���?A�Ş��d�æ��`4E��S�`Xr8�rL~Rr!�I��t;ߴ��'v��v��F�8�
� �_*m�ѪΓ~�l�d|Ӗe�!�oӎ����n埨�(/O(aR��]ꬼ�`��4dY�"<OH˓�?����?	���?����򉀃b#<��	Wz�xI H���l��IF8Q�	�$��C������ӥ%�3?/`��/p.��&)�/X���OzO�����U�]7�y��S3g�A�(�"���j~���3�v�X�ҩ@���j�Iiy��'�2DO:L,B����֝:1�sB�߾ZYb�'���'�剏�M��#�?���?a��P]˦ r�ST� �1g����'Mj��?���e�`���$M/rؐ�	�)I���?�����N����'��T�Vz?Q��.l� �U͗�{'���C\�u�NA����?����?)���h���D�F���ۇ!%^�"BN�1�,������V�D���I,�Mӎ�w$�� +=�d�x��lFD��'rR�'�RbOi|�67O��
ؤ�J��Y����hذhS�\�&���{(��A�+-���<��F6m�O&�$�OL�dO<gNYȲ�x��7��z�L�4V��kܴu���c���?Y���'�?B�?o6�5査`�M ���u��I��	Q�i>a�	ğ@+\���i�g��p�,@C��J03	����K��$��Hf>����7��O:�-a` �����|�#w��a�N�!��?y��?���|B-O�m��;��d�	7��@A�?pf]��k��,ބ�ɤ�M����>���?I��]�6�����on��)q��S鶸)���Mk�OL����-�(�r��t�p�p�đW��9@�٬Y�d�O2���O��$�Ol��.���8;���Q�����8~�|�����+�M�t�J���覵&��/	�ԡ��M?�����'ܓOl�$�OX�Apo�7�i�T��9 �e�F�Ąނ)bщ 9�TUY#�ܕo�d1�Ī<ͧ�?����?���_�u0�1p��m����c����?����D��ۤ���,�������?�(�l�%&D��$*M"G�>�r!�-?a�Y�����H&���ߟ�ˑǐ�v�]m�B�:�]i����)����C����b��OL�AN>9T��D3ƨ���?W2�p#�?Y���?Q��?�|r*O�%lڤW��Ӑ� M&�A0TI�&|W*��������ɭ�M����>Y��if����ӹ-� !F&R�n1Z�뀩z�ttn�����l�<1�8��lQGE��t�'R� C&o��m�ml��c�'��	����	ܟ���˟,�It��B8jÄp��+]�U���L� YR6m�/�|�d�O��D!�9O�dlz�aj���
�l(St�ơ;�0��$���M;b�i�O�	� ��Xi}�6�h�	��ɿU����E?iM2���be��[u�~�%��	Fy�O|R��9A�"qK��K��(��&8=��'6R�'T�I��M���?���?�r��kwpix�HF�W����q�����'��ʓ�?QܴS��'L>�
�蜤1���3�9��Xq�'���� 1٤h	A�������Y��+���2]�H�K�O>T(�`b�2�����O���O���0ڧ�?��N�|��ab&�؇j̄���T�?Y�i��ׁ����	��M��w��M�É���tcp�B)6�Ab�'�2�'"/�e�搟8�����E��)_"ˈ��e@7td��)$���~��O���|���?i���?a��p��DK�K1i������m�L0-O1n��{��a��蟈�	v�s���b��)b�!Z`e[�MCt��`M³���O���&�4����O��C�AZ<R��ڟw�����O�r%�6m%?	��͢94���G�I\y2�|`@�0C�A�]T�,��
N��B�'��'��OU�I��Mc���?�q�$[FL��ǬW�$�IN�<���i��O:l�'���'0�F0}4L�s�ǡ9
&L�"�իw[ 9Yg�i��� V��9�!���ߥkc/A�Z	F�q��ƈ[|dƮ|��IП���ݟ��������r�3z�Vb��F��X'���?����?���i�j���U����4��aU)2a�ܻU*̸`g��gnHpF�|r�'o��OP�8ʄ�i_���*_����\�k��%#�vs6
PHL*y��&��<���?Y��?1�m�e�9�����e{\��3����?�������������@���ؕO��@���@<0� 8���	�Oތ�')��'�ɧ��'rɁ�GO�2D`Qg�( R� �#�(�x�8 ֒���矊�2�� ;�O��Z'm�-G�f8�)�_@�+ +�O��D�Ol�D�O1�:�\��Fe� &܀�cCKӘT�<�S�;��j��'��s���,�Ox��� T�@�$�W�t�B,�`'_0;S����O�L���h��՟���L
*\����.?� ���,=��SI.9`FI�b=Oxʓ�?����?!���?����6c�z�)�u�Z(3Ń̓>��oڙk�6���ʟ���i��ʟc������N@�`i�AO4~'��`��7�?���Ş*!�5�۴�y����'X���sm4�D4�A��y��؝<����ɑ=�'��	ϟ��I6P̪ܛ���x��<��;�f��������'�^6훞`_
�$�O���	d�ִ�.T0\�P�WgN�~���`��O��$�O��O�Y��F6gp(k7d[gZd�
�>Ot�ď�aC�$���z�2�@�����1e�@|�I�a�z�q�K8g,&��	��	ߟ8�Iw�O��G�j����͝ji8��d���Dw}ӨeZR��<��i�R�|�w�
��UL��މ2�F7��0�'�7���A�ݴA��-)�4�yr�'jv9Q�JKcj^���@��%��a��Z�䓧�d�O����O��D�O��NpN��;w�̜dS5Zw���j��ʓO�f,[7���'�R����'���2�H0 @J��U\l�vm{!�>���?�M>�|�`�C	y�~���̝Q\!h�hM.%�8�4����䙢�������O��F�UP儃�.��8"DW�$;,��	7�M˄� �?Ir��f�� Hee� (D�0�!X>�?Y�i��O���'�b�'H2�1}m��Ǡ�A'R�EF��m�$�i���K\+7�Oc�%?��5�~��f���m/�aԀי!���	ڟH�I���I����V���2Ĉ�)����I\�r.\���?��n�������'�7;����I�p����~�e{Q�V�n�*�O����O��Q;(h:6�.?�$��)��A��ʚs�f8�U�
t�˲J���'�t�����'�R�'�ܰ���
��l��h�05�����'`bZ���۴r��I��?���	�&Y�%�6`]�P�w�ӕ��	���Cզ��۴iK���Iw���J�E�t���j��͢[�����8k�(�g���S�s��]�I�t� �K�!\(g��Y���	3_@����������)�SHyR�z�.tp��_"�q1�k	1��I�D�� ���f'���I}rLi�Z@*C�ȃ\�X� �0A����!���9i�46�LPڴ��dI��"H��'��S#|^��D�_F��9x��Կ5�r�}y��'��'���';2[>�!SNʦ`�4�P���Q�����M;&'K��?	���?K~Γ?ڛ�w���1�_�&�ι�U�l:D�+�m�"�o�>���|r�����Ɩ)�M��'KPM2��[��t��ꐻT� L��'$.���OF?�M>Q/Od��O��i�B�>BA��EKr�,9�a��OR���O���<���im����'�r�'�l�Z	��H�+�N��Y��D
@}-aӤ�nZ�����v鑶&q ��֋�Ys��+���I�ooX ���!�/O@��K7�~2�'+�4�� �>qX��4� 0r��'1��'���'�>��	�6;���9~J�	��0��%����M;�H��?	��Un���4�d��Ċ� Wr	�Œ*~�a��O �x�V(mڃ��oZw~�B�!?̠��?N
����S�@)H2č0x��=�I>y*On���O��$�Or�$�O�"�R�-�� ن��:�̫�g�<9@�iD8EH��' ��'[�Or�]1`�D��b葩$� ��ҳB\��#��� `ӚY&��S�?���>���a�A�(�0���'�j A�����+Od ��4�~��|�\��*@cμ��y9�!��j��x3���p�	şL�	��Sty�$}Ӑ� g��O ��Q�0!��Q�!�9.e�%�6+�Oto�p��H��I�Mc��i�7A�-����/[�Ƀ7��K��PC�Fd���䟬�SdT)��<q�'��7��_|��%����@%���<���?��?Q��?ɏ�D/�>Ea�$RM`�P��N,�b�'G��qӰ@�2�N����M%�Xr+�o��<f�P�Y\4�6EX��ē>$���z��Q��6�>?� �L�CP��7f��l*i�� �	H�������@&�x�'���'�b�'n�����j�P�I�I�
^��u�'%"Y��شS���
���?1���V'���2�0�$��Wo_���ɚ��d��U�����|Z��4��(�%$�6A|�u��F�8]1!k�hX��B$�"��D䟔u���j�OzA�!R/�4`����.3ڭ��C�O��d�O���O1�&˓ry���oV �F77J}���
$a�����'Br�tӸ��(�O��m�w�hT�V�.�jp��ʯ	Pi��M�gE��M�O�� ���<����$l%B�+A�L>p��˴�]�<�.O��d�O4���O����O�˧0����@�Y�*,�����Im0����iB����'���'i�O���m��.��M��\��N^F9<A��͇*�R�m1�M�G�x��$�U(�f8OVi��E��H�h�ãa�=6�h�>O��jU8�~ґ|�Z�p�	⟬*��˱�&d�aI��o12���U�����şT��Zy�kaӞ5y5 �O����O�\��M�i�� do��Ab�ASK)�������OR6�e≄RKVe2�L��w_���ަW��	��{׈ʷ:�oZ��D�����'"�X
u�x�yA����R����;��'�"�'����̟��FR\�P��p���й�D
ᦹ0��@yB%Ӣ��2g��i��ݑN=L��S�K�(� �I:�M;ƹi��6-�-�d7-2?a��nP|�3� x0d��}:�b�C2S�ň�.��<���?����?���?�u���v��LB�G��<x�����Цu) ���D����$�F��'HD������=��hȄe�Z��1.�>A��?)O>ͧ�?9�j�2%I�g��W�pC�O�?H�04��M;�O� ����$�~�|�X��	�A[.�1
��� zB����ן���꟬����Vy2�o�D���O�	��	��!��s����� �O��oZR�z��I��D�	�X3�JQ�3�\�-T���#%�+7�P�l�_~��L&� F���wS�(r&�U�U�v� F�(_�=ј's��B�+3�p SƔ��AH¢y+�'��n�X��%�?�Z�4��daP"�*>�j=B�MX��!  �|��'���O.�뗻i���������� �s��X���H���7���<�"�ӫe $,��
�7V���0�Q�O��n� g���	�l��h��F�k`�;�+M�1]&$KC�����Z}B�'�"�|ʟ��a���X���ҝh��b ��]�,�1(��\[���|����Ofm�L>�&�H(@v�������!Io<�i��t�bGT��T8#�M��5*����**r��'z6�&�I4���O�4��c�49�0v�
X"�ś�.�OR�dO�J�6m*?��9̨�']"B�SH���u Y�6�	jd	��.k	����O��d�O���Or��|ڑ.ܟ�L���I�)�䬊�1՛6��S��	����Ѽ�yW�͊ �0��@��D��D�6cƢS��6�C��N<�|r�dT��M��'2�q�Ը/�н��B0x��s�'�N���(�z?�N>i,O����O*�P��0%�a �� E�B%���O���O���<�¿iK$��t�'���'"��)@Ċ#X�Fl84!�ZN����\b}B�'���|匎ƚ�PP� .."qI5����X9\��Ȧ�q�b>�ѡ�O��d ޚ勄œp枱:��:"���Or���O>�6ڧ�?!�P-4n�U:e�O�
p��1s�\��?�!�i��mt�'g�(`�`���S�x��ĝ�$�ȉs�i�I�����ݟhI#O
�5�'t�����?1��dХ}!t����3�ey"�ؚmM�'��i>!�����ԟ��	8>^�;EW�q�ʠ���Ja�͖'��7��*D��$�O���;�	�OT�b �ƪ2�by�oY-p�.q��.�i}�'��|��t�R-3Nc�I�nRP��??`Qk'�i��I6�Ԉu�O:�O`ʓP�m`�뜥˾�3��˝C�!+��?���?���|�*O�l�P����I�{"�9�,U"w�n��taK�X��I0�M[���>	���?���c<:�hp'_�>���G'�G���2�T��M��O��&g����&�I��X�12��lA�I��86��t6O��O���O��d�O��?MH%�I�}X��/.~`crJ�mb.�$�O������
�nl>A���M;K>!ӾO�R���>[�z(Q6lG���?Q��|�7-���MS�O�N�>VAH��@ ���<j�L ���5d�O��#K>�-O��d�O`���OKǸ8G0��J�6F�l�vG����'����M����?��?�+�l��f2~�n�BT�N,~�tJ���p�O���O��O�0Y�V�`��{MTT;E���E�&�emջSL�wdKgy�O�J�I�-��'�̭y�-kL���OE�.������'|B�'�����O���"�M�1�	��Չ%���vLn�#B ]:�v����?Y�i@�O�1�'���+&�"��!@�G��1��nɉ�R�'�u(Ʋi �$�?وa��?�Z���D�cn½�4�R�I?Ԝ�5�|�ؕ'��'(��'#r�'+�S:�&aÀ�k�\�2d͜&	�5A�4b�4!���?�����'�?���y�j�\�i���~B���\�j�b�'ɧ�O]� �¶i��$ѪG����T��#&��U�d�Ŧn��OY�R=z�'.�'��i>��I9A�Rq�͖� _�D�2J��* d��Iߟ��	����'%�7���l����OB�D�p�H�
�F_�)����$��D|���
�O��D�O��Od!Ya���Z�AD�N�X�Q;O$�D�S� 3��|ӈ���t�����ɻbs�A1B��Vo�i���G�[�|]�	������T��o�O�" T�IdҠ ��D7aC8m��
�	�j�d��4�<I5�i<�O�0�5��'�'� 9sFV#F�$�OB�$�O��p��i���,@�����?� D\#'�J-*�d�<R�0�юDN�ky�O���'���'���;�(	��� (Gb�"b�	�k�Ʌ�M[�_��?a��?)�'��9Ob͉C��xF����cP�ĳ�B\}��'�|�O���'��XI�M���Ƶ���*E�i-�S���qХ6|U�D3�Ļ<�Ќ�!eHҔ+��"'%���r"��?9��?A��?ͧ��JƦY���WƟ 3��?.X�rA!�(.j���uc���۴��'o��]�V�v��m�;sBl�(W�ϣCL	�˘59м\���9�'���r�Q:N~B�;t��ƌP?d=rw�-y����?9��?���?����O��$XA�R:������Aӎ���'���'u(6M_,k����M�����d4 `n�I�#īZn�Y���b��D'��شQ����O��t�i��O�@�� l1+d ��d��B�唀[ZRU�4(U��~��|�Z�h�	����	������Չn�v���@K'PS<H�� �˟���xy�lq����Ê�O����O*�'J7�����o��$A��H6��'u��&ΛF�f�<�%���?�y���vDI�g��k�T��#���WC��������+OV����~r�|�ѻ1' ���V�,@�0ꑡ;���'���'���[����4���(�G5vT�c@ۃ0 ����e���?���h�f�D�Ay�i�V	���F�4��煋<wvF�*1u���l��8�fMo��<���_6�������)O���6��	yj�zeo�:��q�1O���?)��?����?����ֽoD�I0 
�/Kޢ�`ģ�;Fy�-oZ!|B��������o���Xj��������2�BY�N'��cE��m� �O^O1�Nl@��}��	#��L�䠂8'���1	Q
*���I�*�[�'��%��'aR�'4�="4,L��e 1R���gD��?���?�����DPצ���#�ߟp��ݟ��1O��z0��Ϥ���R��J��JT�	��McD�'?�'4BѸ�@R�i`�� ��� �Uk�O�+f6	S^�ƃ/��S��?�ƣ�O\0CT��JK��j��(*��2��Od���O����OĢ}z�e�H	��~��x�0M�!�.i��A���ʙ�O�'a<70�i��Yê͙v7��S�돤c~���'������E2޴4��!K�4����1V��e��O&�tr�I�`X8��B�Q�h!j�|�R������L��ߟ\�Iϟ��	�"|��҃�P
)�8)�d�[y��h�Z�x���O��D�On�����D!Ƅ[�(�!
v�:#BQ�	f�ʓT����t���'����?9�S�Xj�8�M?K#�,B׭��W�@����}�-O��J0����~|�T�8�G�׏]���h�G��[4�ןX��şx�����Zyb�d�L|�sJ�O6�"�J2>�R��=�%��	�O�)m�f��-I�	ş���Ɵ�Sdӫ�Nt2�JT��ΰ�u��>`���m�U~��WR�������O��..�j���3M�D��B��yB�'B�'b�'�r�	��	gV�cS�ѯF���i�3Ո��?a��iv�@�ΟH�n�A�I�4P��+4D[�B�)��Ĝ�l��%������SW��Qmo~Zw
��)%��mZ7']]j�i@a���T�z��I�u:�'���Οp�	��H���`z��P�%�N,�Q8���'�@��ş�'�6���*ʓ�?�,�n��n��ȥ��%W#�- W����O���O�O��Ln<,Xb,)�$��D�Y�����Ct��l�L~�O�1���K Qu�)Y�"YX�/O�j
b���?9���?a�Ş���Ϧ��@�ыt��a�5����p!S]�za���O2�D�Φ�?I�S�t��#�B���zA�)��WM=��	��l` ��Ǧ=��?�Θ�#����yrhI�$4n��$ᔱH_��EC]�ybS�x�I��p����$��ڟ��OO�]#֍Œ96�%�CJ\��]�qaz�R�* ��O*���O����Č���]�"�<xfƍ�8��`j!!�;�@���۟H$��ğ���20��mZ�<�`�1g��$����z��4�1Ȁ�<y�.K2�f��N�Oy�Ob��.1�N��7-�~�L�C�eMv�R�'���'|�I��Mkq@H?�?����?Cb�h|D&I�=�H �G����'���i�&�l� �$�����} �cd�4d`0����k�X�	�>������Kݦ�x*O��)��~b�'7� �J)m/�E5�(��qb�'���'��'x�>����0*Y��G%�<�e/G�0 H�I1�?)��S^yRClӜ���C��A��@G� e��n�@�����mZ��M��Ms�O(��2b	��J����عa�Fϗ~��{d=D���O���|2��?9���?Q�TA䈉@J��W���#ƈ�~�ę�/O�n�"pf��I��p��h���(�U�]6A�QǍ�[H���S�����O��$>��F�\ބ�_k��|�@� 5B\�gg[�dZ`�Rl�ԸQ%�O�i�O>�)OD���^�t�z��q'�|�Å�O�D�O����O�I�<	d�iZ*���'g�-q�$��7�� ��D�	���'��6�3�I���$�O����O��萨�)x��IB��/s�FX`F�W[�n7�w�,�	�x9�~Γ���;G��H����U�1c�$^�e�$M��?���?���?���OD�,�V�R�<�FfC!w=���'���'=N6�ܡL\�)�O�tlϟ��'��O�;?b R�E޲l�\p0B� �D���!y�4��ɏ�Mۜ'k"��h,����h�/rbɦ��T�\�Z4Cj?�J>�)O����Oh�d�O0�)��K�$H�`�γ#0���p��O����<�i\�@��'W��'��<�V$I���k8%Aů��xK��^��:�M��iJ�O�S�F��1��O���01l��@1�`i4L�Ay�mZ"��4���'?�']q��?�9(�"� >	�'�'���'y����O9���M���ʨh(�t�T�ԣ	uܽ ��\�ވ�.Ob�m�B�u�I��MF�5�v� V�[	�ua��3f�ƅm�MC����M;�O��K3����tZ���E��(;�eQ�2���҂�w���'O2�'q��'2�'��,X�1��@�7i�8$!u���V�c�4/p�����?����'�?�a��ygׄz��sD�5��zQ#�F���'Eɧ�t�'BDۜ���?O� :����G?#� 4�)�,�9��5O~�����?��@7���<����?y�%S&S�X8V�̙�&�����?����?������s��ΟH����#�bP"3����
��L�8eY'J|�y��I�����n�I�~��3FH ����ďg��@<ek�g��M��.r?���d��4 P�E�{�\�c��ҰI������?���?!��h����9���	�J[:_��;�
Ox���Ѧ�/�y��|���]�t,]��f�*v�ܸ@�r!E.v�\�	��	-zA��m��<Y��H~Q���?Ȁ��~��Z���:�UxqJTA�I_y�O=��'\��'%�*F�D&P
� D�)�#�-F���(�M;�P7�?���?�O~Γ[�F��RL����,vY�P]��I�@%��ߟ��ɅBj� �JY�$� �0�O�%��U�����'�,�e?�J>+O�Š�\�ps��#��`Jф��O(���O����O��<@�i9�QKq�'����G�['j��1z��;"��'4�7�>�ɧ����O��D�O�e�Gܵ!_�:��7|���� ��2e[�6�e�,�I�V?`	��~��z��*�b%H��Ƨ~��sL�h��\��?)��?!��?����OY�tPS�ӄf_JpzƆ �b1����'�B�'0p6�εq���z&�F�|R�ڕ?DZ�b�H�]�f�5�$Q]�'�2���Doߣ՛���P���(wH���=���fT��.�B�O��O���|R��?���e�L��WC �4}*`��%(�Q��?y)O̤l�	�T�Iʟ���M�%�ؼ�1�h�$\9 ��  ���j}��'�|�OI�k��SzAc�*��z�6M1�d��8Uk��Q
�F�����.���>���	~��9���|`z3c�|�.���O^�d�O���ɮ<!��iQ}�=(Y�hI���>��A&Ha3��'n7M;��)��$�O�eRUK�U*�� � =�@Ŏ�Ol��� zF7M/?�Af�
e<J�	.�� 
�(�R����bҤ�f ��y�\����Ɏ[ұ���,�t��U"Ik�Y�4^i����?����O��7=��D`�놴|�Re�[��$d�%n�����OV�O1�*�s�i��ɨb��m���8b����c�'���I���3V�';f4$�ؗ'�'���o� |��:Bk����'���'v�S���4:���?���Hg��cG��v��D"�dN0��Y،���>����?I>�u�_1N�� �Vo�

6�)���a~��ޮ���"H����O���	�{��Ƈjx�q#�!/B���B �{	��'=��''��S˟ P�1v+��q��	�b����c�ß@��4`��<���?Y��i��O��5-@|2�ϾO�2	/�<���0O����O:���S�7-&?�$,	,,�	
�Q=5����4 ����*2΄<����4�����O��O$���p��M���r�z�s�&H1�ZʓJ�B�E�?Q��?YN~Z�y�n���%�:" 2�/�-\T`��R\�Tb�4s���*�4�Z�����8y�⁺tJDmq���� X�A�a�L�뷓���ԄH��n�h��Eyb���M1�TK�l̠H�%�$�Bk���'�b�'��O �;�M3#�µ�?�@�k	�p�WkX�V%��G�,�?���i��|�-�>��i��6��̦q2-� w��1��� ]�� 8�U��lZ�<A� '��*$F���@�'E��9�ѣR�Ыt"��wM�;6亜'���'�B�'�b�'h�xy�@L�to���-2*����Op�$�OT��W�vhͧ�?٦�i)�Z��zG'˓l��9��W'R�.�е�+�ē^���bw�����$��6-y� ���w��0c4ƱH�&��WlT�il��0�ٴF��D%���<Y��?���?q�s\���� '����#ӱ�?!����I��Eq��pyr�'�#e<ْn�2<���d�?3`�jg��ٟm���?���=`Zx�*Ϳj0 �3�O�� �#�Ee�LmZ����Ĥ�'��'.�It͓ 8$(a3�$��6F���'�b�'-B���O剖�M;���1{��,9vE�M�nPAs��[����?���im�O&a�'��7�K���}U䱲W��Yx��Z� x�Vo�@�.!o��<���=���c2�?��'�D��`�(#W,8�7��8F�le�'
�蟌�	��l��ß���z����$�H��G��j�#��@�7�ݬ"���$�O|�D#�	�O2�mz�ʇ�V=z�&�x�o�
-0��r�� �?��4ɧ������R�M��'F�I���¦���R�s
��'.�ذ���p�!�|�^������p�I/^5}H$�(�
Ebqd�ϟ�������	by2
p��u���O�D�O��Ȣ���_윃��+�L��%c�O�O��'ub�'��'P�ك��F!5&�aFm��a�R�:�'efB
f�y�V!/[��?aC��'�lE�ɕ>���Yʹ����`��I�'���'!�'L�>I���:D�Х3���ɠ��$����2�M�%�X���$˦%�?�;<��Q��)�"�>m��N�(gi�Γ�?!���?	�	7�M+�O������O��JL�)k9�Q��X/�1P���	]y��'���'3�'�b����r-�ы�=VY*#�\�I9�M�^��?Y���?�M~R��M�rD��� +�h9ʡ�O�����_�X�I$�b>�ie�*� �1��cF�;��ಡ�[&Bj�p��#M�ʓnA,�"�O�5�I>	)O�� ���'�D��@�.��;6a�O��D�OL���O�)�<�S�i��@�'FXݒH�P7m��:f���T�'!b6�&��"�����8��Mk��S�(#�Й���s�\�:���6;kh�ߴ��d�6�(1���&tv����A#g-�@0�\2s��ى�iK 9t�d�OJ�$�O6�$�Of�D6��[ڢ�+��בt�9x�k^=z����I��8�ɔ�M+6���|r�v�f�|B.�9-�V��`A��t�n51琒O��D~���8?d7*?	���� �Z)�d�/&˾��E>,���/��$�`�'��'Z��'�z4�Ue�^.n,�Ō�'m�vy)��'�W��:�4nJhт���?�Ǧ��O�����^&��f��f,��O�A�'��6�Mܦ=
O<�O��X%�-@r�	qb�h�x�!H�Um��9e�i?��|�o��%�,	W��|z8d%*шKmX�R����	������b>��'�7ئ ��]x����V,�[����@0��.�<���i��O>��'x�7�ZS��10��3J8eP�4ThQm��M��G
��M#�O��6�3���[�dyP�T/[>�p�N��(< ��l���'Sb�'ab�'��'7�Ӳ �,�s���5N�V x M®��L�ٴ&�ܩ��?���䧃?� ��yG�Iרl�r�Q��|5H �3�r�'�ɧ�O�z�{b�i�dŴE���Q�v�JDs�_7#X��I>��q�'��'��i>��ɂ&�P��G�2�r,�� �s����I؟h��ПH�'96M�;b8����On��7���*���%1��{ѮY�m��⟘��O$���O��O4�91�Z,mFz<J#�%�px�К��xtD�$�f=nw̧H����D�ciW�S���f��<�)�d���������	�F�D�'�~X���U*?����
@�V���'�"7J�t�����O�l�e�Ӽ�4 �*7�h\�!�٠�|�Ѷ���<q��?��k��pٴ��D 7}�i��OP� F�����R�\55��a��|�U���ן���؟@�	ɟ�x�O��tpі���@6
9;eWNyB�|�4,�C��Op���O��?��S�T�e�
u�� �����'����O��/��)Y�X�
x�Lʀ{&L���'sc�w�b�,�T|`0���L%�8�'��Ё��
p�\�Ů�7z�m�D�'�"�'�B����Y�(��4:C�Q���oa<͈���>G(p�Ʃ��vΓX-���D�K}�'ir�'���4��y�%He��p�x�#�LF��&����E)�#A�Q>�� ���:U���·�Մs���}��8	G�ؒY!r��ӥȢ6�.�a�ҟ ����H��4p\��O@�6m:�$��:,� pF@�5;%������8s��O����O��J4�7�*?��,��᳣�>��f�[5%�@D�1���?�O9���<Y����q�"�{� �+T΁��Oz�l�>���I����	y�ă�7e�졐��>y�&��#0��D�U}��'�r�|ʟf�Ң %Mt��g�_���(�$�  -ԥ80�� z�j��|·�O���O>���S6'0�&��3]�P�=��2ܴ�� ��H�
��5;�˛%P�ƔH�NI"�?���R����n}��}Ӷ�����<���r�C 4c���j�����4h���*�4��DǶU���R�O2剅 t��`�	�@���v`ޑ P�	Ny��'p!�MȲO,�YC�g��o���y��f�D��	�O����O$�?��������3��-)�j�����?9����Şm�̄ش�yҍֿF���`A
�o^�l���+�yBd[�\U��N��9Z���>itH�� �	Z\<C!H��3T���qA�&��̒4JU1��-�Ĝ-\=���7׼Ţ���=?<$	���30�"�Ǝ"6�V	S� �<2������
�l�A�ҭ3�V�*O�*4�
�y��
�$
�uP�*r���HG�{7@O�Z�0����i1��+/.��� %�W�Qzւ߹(�jခ/ �2$
H����]Y -�(�:�ʃ#�c�&1�T�1m��=��`��:���h�j�J�Ba3�ߦU�<�0���n��/[(^���Ҫ�~~6��O��d� #BD)�u�3����dO�԰�o�ȟl$�d��ȟp�U�џ4�OQ�f��@Rd�"�&;>��i�R�'���:����������O&��-h��S�*fP@X�O4�h�'���Iޟ�
�GOp����4H��x��Iy1�V�K�؉9ӊР�M(O�����٦}����L�I�?�9�Ok�H�$�d�3�X'�����?'����''r	ʽ@Q�O��>q��o�yZ����^آ,��y��3�˦��	����	�?h�O�˓f+����Hi�vp��d��RLܜ��i�����>�ğl�CM��. y�n�r���"m��M;��?��tN���vZ�$�'i��O -Z�!U(v`��I��L�t�6lA��i*�'4��y��'0��5���C˨���TVAcSI׋�M��4� ���Z���'�R�|Zc������r�jAxSO)/��#�OvqcS�"���O�$�OH˓2
ι1ᇥ	��s��+L�|�S���u��ry��'��'���'�Z|I�͇�S���'�FX}�8�c�9Y��'M�'�\��b�G������B�]F���g��'B�r�ۦM��M�-O>��9�d�O<��CaB��I�1N`���@�a7���i�n�드?a���?y+O��#�[Z���'O`� DX3�Y�P�5��&��x ���ջi�"�|"�'�.��%r�Ot͹�\�#�VP�
�@��4�?Y���U?�6Q�O@��'��4�ҌmO�}���W-d��L�xo�O ��O�p��O)�	[:����Y�%a�FϠM;����a��Y�'�R����|���D�O��D����ק5i�&��<B�,>EJw���M���?�'�F�?!H>�����u�~Ī�
 n�,54,�+�M3d�����'���'����>a.O��cRK:|�,�, �) an��%n6힌C�.⟤���/��bp��b�:A���0���J3�i-�'i�b��\� ����O�	�H��UZ�ʝ::l�"���K��c��!e�`��Ο���矌�'� ����3�',E�U� D���M���.�h`��x�O��|Zw�RA�G�A����9���,Zp0H<�����$�O��D�O�8�j��R�M�fKZR+��.���h�eϿ_&�'\��'��']�i�	ze��>�0��AQ��u�W@o�����<y���?I����ͩI���ͧ>}0P��O:*jnp�����B��'~r�';�'�i>5��Jɬ��sʂ�A8(�3̇`���aK<����d�O��i�a�|b�1~��j����u@l�E�8$�h{`�iL�O���<�&�G�ɏKe>� !���ZG�u!46m�O�ʓ�?	�e�%����O��$�k��f��5���B�-�~P��Y�3�'Z�Y�Ș�A>�Ӻ�W��)�*Ē� O�u�)�b�Jn}B�'�L���'fb�'��O��i�5袀_ L-j�zd�ؘY&��t�s����<�v�@_��ħbt��m�#�:�yG�D41Ӵmn��p�������	����myʟ�I" �?�v	j6*
 (�!k�^}B���O>�(2
� �#�v� dW�M���?i�g�T�b)O��c����#����B)��-��������Fxr�(�)�O"���O����$dHirh�$c�D��G���y���-�I<�'�?AH>��6A�}��%߃�$�ʒ�_��'�\���	��x��sy�HC�;2��P�07�aa�$w�}��?��O��$;�$�<�;+Cv�0d�?5��	Z�`:�xm�ş`�'���'U�]��ء〢����	�i�z�c�+�"2 a0r�S��$�O��D�O@��?Q.��$�4g��H��+�&�0���`X���'h�'�ߟ � ]F�D�'i$X�/�++�\���G�BN`�`�Di�p� �Iny�=��f��Q�`���j��@�O��_?\�l���'��  M���ן����?��Ct��@聹O�Ƒ�!g�bMO�d�<�WD�{��u�J΁G4�e� ��y`�wnD ���O4���O����O��D�2�Ӻ�G�+qS�$ځ
Z�"R�i[4�ڦ���]y��O�O�~yS��'�h�jp�:��I�4?#�X8���?����?��'��?}�ˇ<~���4	 �j`ڐN����A6��b>U�Ɏ<��Q�D�����ϐ*bJ��z��iM��'?B&�_�O��OH��2w�.�K�P�@�	�C��?�6M�O�ʓ!����V?��ɟ��Iҟ`��ʌ0]U"��V��x?��j�)ë�M��3 _���'�RQ���i�HQ�{(�brM�#9��ӃE�>yp�E~��'�R�'�Y�T#�H�J h��0Ʉ�.`Jh�S�G+���O���?y/O��d�O���ϮT��q�g�5��ɪ�h�1g�,��=O ��?��?	,Oְk�G�|���8��:AǇ'2u<5�K���'_�P��I�x�	�5���q��]�������:��5��xm������՟��I_y�*��h�r맺?�1uW�AK&��+��]I�m@%(�`m��t�'"�'��A��yB�>I�Fp����V�C�N�I�_ڦ���şԖ'��(p��~���?9�'I4�1ȓ���Y�wb��|\���'V�x�	����I2V��IF��: ��S�i1�ILy�!�Ҋ�Ѧ��'�����ei�4���O���H!էu�`�.��pq�F�"\��B�1�M����?!7-��<9N>I���Ǘg��� ��!4Z  ��ȥ�M�@Ο�u�6�'b�'�4��>(O�<�Í��A��(<�X��p%Y�%��7m��-q���R�NJ�!J�}����b\�_	(4hc�i92�'��J��������O��9�(�A�OQ^�.T��w~�7��O�˓rpT�S�T�'��'�(%X&.�"����F��	�����w���di %�'R����'SZc1�K��U f�ޱBS嚦o�Z�O�0�?O2��O����O*��<�!Aּъ����%;p���ׂn&��&]���'�]���	������W�z՚� � *0$�GeU>8�8j�Ct���� �I�<�	Ay�h*f擦όܱ�ނS���i'&�"a^�6�<�������Ob���OL-��Z?Yɑ�Q=&j�R��v���q�Mj�V���O6���O��3�	iBZ?I��
F�4 S�Z�oX ���hP�%v�cڴ�?�.O����O@���%��d<}r���{�ꤱ�g��IϤ�Rh�MS���?�.O"� ��}���'��O�Yad�>�̴�fl	 ��3�	���������7'r���	ZyB֟�@�b�k���J�X�h	1µii��C9����4�?	���?y��K��i�� ��"�
�H��8�Pi6;��Qw�i��'J��x�'��I��\�}J�G�\���G"k1���'�W¦�C���M+���?���GS�`�'&��&`ר,��7$P�,by8t��ޭ	 1O���?	����'6v�гNQ;=����Ō):��Ч�x���O����
��'��۟X��x4���^Ȱ��t��4��oZ�<�'��2���I�O����O6��q��nUԱ8V,@�%�蕙�`�Ҧ����{���ӯO�ʓ�?Q/O����Fk��).�B��0�bXp� S� *Ai~���ǟ\��� �	py�A>S��u5H�#���WEL1?Of�:���>	-O\��<��?y��3�b�;�H�B�*���MRI2س7���<���?����?�����B��|���XAj@hx�*N�hB阴C�O���?�-O��$�O"�Ă^�ɴ� !+���C�LIJCѢ���?��?)(Oޑ`rhHi���'� �r`k��m8�@+Vc�IQNv�����<���?	�?x�����ɘj0C1e��!_����֡p�^7�O�ī<qD 5l	��՟����?�Pp���`�h��Ú��q������d�O����O� ��>O$�$�ON���?�r�a[�"��qzaf�I�^��dn�<ʓi�FI���i���?�'f/�I�hP�h�	�'�FU	 $�Y�7-�O0��=1Y��$=��7�ӪN��rP�!n�����"�x6m�w��nZ��I���������?Qb���~Z�8�*ߣ�갊p^�2�.\�-z�|��	�OPiIv/I�L@�q1*�o\���&�ͦ�������5,D�ĨI<���?�'���֌�0x%@�pPd�kX.T��}BH
2��'.��'��"�`tj'�A�qZ��`�ǁ7R,6��O��p'N�y쓑?�M>�1m�l@�BNv*Zt{TDT�#�U�'F�`�|2�'f2�'�剡�@	����.H�u�F�_�q�ؐ[�*�����?)�����?!�/DűR��A��uJ�F��|f�IX��<9,O����O�İ<I6bӄQM�iR�=�t�1C��hx�xV�K�'��|r�'�BG���y�G�q���PHͬ�>�91�̶H�n��?���?q.Oj���g��JX��  c,)��������d�T�D.�d�OV��޹��d!}�͒n�b�9����a>�8�gC�?�M����?y.O�]��f�w���d�Ӗn��&-�G�
m3-֍��P�M<���?Q�.��<�L>��O�>T���5Zw���̮NH�̉�4��d2re�xn�����O���Rg~���=:��ɲ�K�˪P{���M����?�2���?!K>y��$A�+~V|	p���4lR+���M�E�ÀG�^~���'���OwO&��PHԤa��#?x�m����b�xXnZ�p�.���v��Z���?���QA&( �!ܻ�1n��0��ğd��FC���'�B�O��P�L�<I@�1�o�0;��ұ�i��'z�A�c/���O��d�O9�䓕m�t-[�d�2m|�jΛ¦m���)���@N<����?QI>��O�����4b�\C��_3w�z4�'�d����'��	ܟ��IΟ�'=��kV�W��.�+���8?VR	���<fM~O��&ړ�~��@7���C!Q��j�.���M������Or�$�O����O�Y��O�a���?'X|}��m�0�� p�NVæ-�I�H��R�	�L�'M佘�4t�������n�H��a�:K�e�'���'X�\�P����'w9�S�N�J����и5�B���i*r�'��OXii��IS�5"� f��+HH[���S���'�b�'���>iR�'S��'��G��|z�	rP�K6���\��@O>�$�<)��O|��u7�R*c&�r`�U.�:4"G"��M#���?ApnJ�?����?y��R��?��K�XI(���-T&���/��]H&�oZ�t�'>����t�D�'�!��)�*"RZeZf�Poڸ\b���ܴ�?����?������4�I#pX�3�/�L�	'һe06��^pd��3�	ɟDa��QY���Y�^([��;�K��M���?�t|�xY+O�ʧ�?��'g �J�L��?�T�r��by��Ѐ�?i�O�2�'��*��4�\��j�jK�q��E�(7��7�O~ QQm�u}RZ�x�	hyB��5�C�*��a�	 a���#t��:�M��1�n���?Y��?����?�/O(��׌K+�~<RfH�4@�	3�V(T�H��'��	��ܖ'��'��MW#߲m�&��"�H��ˀ�KKz�ʘ':��`�����'����4�g>u���z|츸���'$������`�nʓ�?�.Ol���O�d͡<V���2��Zv�A!z�y����d�`m���������By��I�=*��'�?��U)+ �����:�X̉&���v�'G�	ԟ���͟0��O����:�X�M�@h�Nח0��:�6��O���<	ʝR�����l�I�?q���j�!��C�U'p�)1�
���O(�$�O�`���X�'(��K��2j�>�.��t�� b��vY��J��M���?���"vW��]!u&�h��hB�6]����&F/ 7��O�D��jp�Ĥ<y���O3�)kaF��"�]���	4�5[ܴA
��il��'�2�O�2���D^P�(����~�.���#õE�( n��]|��Id��e���?!Ɔ�'Ld# ��~��Tp�	�M��V�'��'�dm2&�>!(O~���� �1P��5DY2	t���p��t1��i�'�l���	�O�$�OT�4g$L��²OX*c4.-c'AŦ%��9
��A�'*�'�?N>Q��Su��{�ᛰz\�d0�V�F��'
F�2�O����O���<р��6W�Y@�S)5�"ű�Z�3��i�FU����柜�����?�G���J�(��ě!X�e!U�[E���|��'���'$"�'�Z}IS۟�U�s��1�XK��e%2e� �iz�	ʟh'���IJy����M�U�Af�`UЕn�O�8�g*�Ty��X%4��]�=E�����Q�"i@�.D�� �P��y��&jg�(Y�`U�&�n�j�iZ��~�bI������	H�Żte�1:@�t�0ʕJ+b� 4U�]c~ɳ1�Q62^6|[U�Q�i�Ը0��S6�05�#�άcA��9�ʂm�ҵ�^(&Ɯ�֥\�]�q�X 9߀U�
7;��سH�k�� ����o�� ���{�t(u郿Ir�g,���
���T��?���?��xd���L�g�<}�!�X�������9���S�J�-)Ռ�0s(�?u�|�ݑ�R�aBFȞR4��I31z�	r��
�P�#Gژ�v�*���?�R���w�bu�
[�T�d��񣟋�E��^��H��?i�O�O<�'/�4�u����`X1�ۧT*���Q��{�/�'}��!
īN�p�Gx"&"�S��藦M��!�I6Z"�P$`�9o�2�'�H�rKI0E2�'��'X"����L��)���(���.ЌQ a�<*8J����*VpM��	62�\�A��?�=a����Z��p؇Un������lkI�����^Pb��g�'�� E1-���fK��	�'/��h��?I��D�<�w�M��JQ��KI��|h6A^�<��ܭW��@���j�
$��(��7���'���!$�mډA�0�;��s��l��O�z�&e���?����?�fM�?!�����B

�AR�V�L�
�W,�'eT���]�uu��÷�<lO�J$H�c�:�ե���!@Vjˀo�m��_<fņ�	6,�����O����̀7�P4�	���l���=ړ��OD,��!��@�� �rF����6"O���QeՎD����UE�0`���<�B\�L�'��Uqb��>���IV�)ֺt���:d�|�lZ�fʹH+e��O~���O���kF�e�D�DA�����|�'�G��-���GO���RÈ�n�'��<��GJ/0�D��d
x��O(�ty!�U�]����$R3�=2��$##�'��X,��*�3G��l�6
,}����2O���䕺N�e��!��V��ekc�B 9a|��$�D�*� 	
ɑ4$v��(�~���˶�I�'��U>�I�������ȟ�TM�~b��ه�L�\(R�+wM�;i�\ș�`N�N�^p�F&�?�Oj1��m��j-ޑ�'�ɥ*����0OS�f�
E��i�T��0���:}>���O�AJ�!�7/xDy�Cۗp h�Q�(�%��O�=?%?e'���SN��A{"��D��L�W0D�H�2F��i;�����E�'^ 2a� ?ّ��PJ�:%��%L�d��%#O,2�*�s���?�`��K�*���?9��?�5������O�I�Ԅ��bb����J
�u"t�O��S�'���PU�,<��qXi�6;��۵9O4}��Mܜv���I��E�j�џ�����/,�K�KE��I�DD��`A1��O^��Ċ����u�V�9y����.��?|!�
<-s�P�V����څ�_��T=Dz����{��oZ�7����D�>�D�H@@�$g���I����Ο�Bwf�˟��I�|r���5t	VI��C�`}�q���؆b�А0�R�N�@i�J�V�Y��If�Ju���ǲ��+�#�<��J�dB�>y��a��t"ȰLV:��OD�Ƀ�'�`�3O��QS�ɚ.A����'Y��y!^0'���dK��o�r�)� �y�
U�.\门�56�3A�#�y?��kֲP��4�?����Έ!����L�8	��J4�L-I���a�O@���O���w&fӐ��d�5}*�s�M
:4�(�R��$H��uZ$�6rn�6M �8X���&u��-��oo>A	GD?Jvyp���(ʔ�Fl?�i��Q�	z�O�DOc��'m�*]��e�ԍ2�!�d72{��[P�_Z?z���#�)�a|"d#�+c'����SI�c��I�K=!�Y�8Ӫm�a�C��D8 ���  !��Q2²T	��>�QZ���>�!���a��(q��}�  tm54�!�$+8�� u(�lkNxk¡[<E�!�dH�0B�q��g�<Mf�Q���B�!�?���s�KN?aK�a��(0�!��5�j�K�eD�k�=s.�5@~!�� D���W�9r����c=x��"ON	�F=	t��U�22mz5"O�T0�!S�ˢq B�ͲX$K�"O�49��7o�%H��4���j�"O�u8mǌ6$ �!, ]�x�"O�l #�6	��������L��"O�"�+��
L6�s��ҕ}��D"OF,��GJ9+Aj�:5+V�wh�r�"O�E���N7���H��͖Y ECr"O"�*�a�~lIE��=u+�&"O|hц+V
]M�̂b	|Q("O�)��0n#*����M-&$T�g"O\}c��'8VDa��߇�Ȭ�S"O�t�#Z�d0)�#j�y|N��"O���i�^����h�5-�̱T"O�����Ƒz�a� AѫQ����"O�U���.AԹ��4��	�"O����.��]��̈�R�ʢ"O�!ÆM�?f��K���o�N��"O��!@�]|�i�M�~Ն�{f"O��Rq�L�H��ٗ�S"��$� "O�E��F��Ihd�J�G�,y��tp�"O�hE�T�g.���I�a�@�:�"O��j�A_�p*��%5��("Of�s�&ι
�E
��I�/��
d"OΑzD�ʯp��
l�:��("O�!� 
߮}s��R���=NIX�õ"O�M���O�|!���']��A�`"OX�	��N��]1���V��"O�d���G ͂�iV���x�"O:9ൊ�.x�d��'Җe�E�"O8���cƓv�,�6FJ?2�I��"O��
� X�H#=��eTJ ���4"O&��¦�:!%���� 
w:��C"O�#��6D&�C҇5l���"O6x�b��>��|h��\�}��"O^`aŦ�~�p�*g@/�J�[C"O�)��E���k�'[B���U��k7�(�S�O�x�u�ߞf,�1`gW�b.!��'����P�P*���I�(��9I>�bH��0=q'Oۧ���A"�
�koʐ���Iz���3�O�%;>�z���%�D0�EK9|��Ňȓ9���K�q�����
)ר5Dr��,i�>��N��#~�,�BhN�}�K4D� �W�;^�����cʫot��H+�<��N�����(�`��&������FCQ5AXR �#"O�@cm�fe;'/PptpT�P�|�/Q�p=�,��KP(x�*Q�2���P�]~h<��CۯZ�����ޥfƬ����Z�c2�݆������݉x�l�:1 ԋl��)��ɋ|�|��<q5��-��Zp(H=i83hc�<� �Qͨ��RLI]檽��čh�IY�?�}��`�8-]̑S��%��"�g�<qUi/A�H��&ɱn��48�G~��o�Ո�W��4+�(HPW��J��ߴ*w:��Ɠb f��R
N�r��'�9fA��	�`��xBD��EY�����U!J�QV����<�&��ј'�JptkЁ.��ѓG]>��"�'%jzE)�//��D�U�N�B�yҍ�O1�f%�1�2h���R4�-<� �"O�;7
�b�$��u�F64>�2T"O�P�h�! {�]���)V>ا"OP9V������E�˚cg.iR�"OD��b��!�%Ś�R�	3�I�y
� ��R���V|(���Z#9O<x��"O����/��F���$N�5c�"O��iϋ)7��1�Y����`"O����f�I?�e�S �wo\Z�"O�dAv�����8��^e4��r"O�L��S�UY�ř�%�0�B	+"O�@��ݚ(���Y$�ŧ7�t"O��9
� �tȪ��S2C���*"O`x�Bo�'¸9�sN��\,�, "O��3�#����DNV$�x���	-"���E��G�9v�����3I�0	V���]��u;�.O8x����F�R/^0L0�I�G���?E�ԭ@���@�2��a��Ѹh!�dA�Q�İsЏ��w���K��j�I=k΁��	)#2l�nO&b8�=["���"(������& �扸+f-R��2Jh�e�mP5�B�	�.c*I�A�X�FD����$U/,�=���ʚΈ��d#v���U��%+F��]b�E#�"O�)@�ɉ�/�(Q�ơL$ld,��"O�`⢁ S�d����=J�"�"Oj8�Daæ8��V���5/��%"O�96���w�0eX�C�.�&"O�,@�[5�]����FD�1"O�Ś�"���6<�%L��]���s"O؀ⳂG�Nz��.Z����"O|���!��ѵ�M*7�
�i�"O�Xz���A��(�WmP@_[�g"O�1	f�N{�`@B4���Hh�
d"O�A�&jV�܈T
6�Ҡw5H� �"O����/ȬR�G���cG�'r����;�)�'=����r�֭P�����K7|)v��'�S�܂W4������[A0�(ON�����t~%@�'g&��r��.���cF��ON��K^���f�+W�Ac��c�ؼ�ԼqSl���S(<���{Ch1�Y�Mv̍+�![�'d$Cc�߰D��](o�}��c� �iV#�������B�G�B�I�}�*tC�䊟Enz9�3�7[�X�L�1Dk�v�ҧ��brf�?��}�ٰ!]֝�3D���D/�w�Μ�J}AN�I�-4�@:�[V)�J�g̓x��x٧�[Y	i�bT9� Ȇ��y&yҗ�h�F����X��1��H(�ވ�Pd<�O�U�SdE�q�e��J�$����'��`�$[�6b��O6=�W���(O�Aۦ�
M���a"O<m� f��~G�}����?�-����FC	���X�>E�4A}.��jǆ=�^"`���y��W�|HM;�ȋh:�jQ��Z���O
iW������*˴�p�Δ3�DS:B$����jK�ᲆO�'h�#�F��{tQ;��>+xs�.)�O$�a5��wZm:�!��jh�(c��ɘr� j��ķ"��OJ
p	�+��.��`�h�;�\]��'y�KTj�8P�LŁ'�8+Pr�'%����D<8��1����0|*b�ܤN
�Kp��0�DҲjTc�<9&���.��V��e�F�9 )�#��	�J�<,a3�!a��g�'A��"�2�J�#%Μ0jyd��
�j�r i�m2,�R�`���6]� b%H �"˒
��~���
��hM��@�b�rc�����O�X���N�VQ��
�%FM�)�=jL��X�GsH)��ŏe	!�䜰˸0H3%_5 Q
�`�a��I�iy� �V��(Ќ	�ç��S�^�@̘Ǧ3n� i��d|pt�e(��q��S�iܓ ��1@��<ifD�1ςA�Ø��}��
`L4a���0�n�o���?���* ��(a’�`����"@�3E�'#�2f��؅���b�U�U���L`��F�3V����g`}j`
K���	�_>���@Z-π��	5%�BC�)� ��� @�5�@�I���G^h�S"�>��(ʣQ��:��x��DIٶj�5��쒟_��{)֣�y��	Rn��N�I���'F,���S�C�g�d��e���#m�#J�@N�`!�jPY��#W�)��;��U.r\!���a	T,(��p��m�nD!��9�D�s���=�U	ǢG VE!�$^�S��}Ha�N!2�\!J�[	�'[���Ao_r���I�9��'����QHP�jH)�I�5@ ���'x�A�ΐ�� �CyLt2�'������
�x֔i�2�B�d(s�'����1��	4�|9a2�4&��'����h_z�l �q��5!�HE��'�F��g�6j'XU+ `�EG�93�'^���I;^C����Cf�lc�'92l�e��)&�p`E��@��`�'{�xj4�I�Zn���w
�&6.V��(Oz�1BF�k���:B:�F��^5%�@�@�6�O�`����ب#�A�����rگxt���)D����	�.x�J��%�|��C&�z�L@��:��D@D ^�в�'Y�=�"C�	4z��]��nV�I�*e�d�I�`�$��߷�v��>E�dό�z��HHS �13lb�i���6fo!��D?/n�A��8m�2�Q@:�	=\���ߓ K��a��|Z�c��A������E��(J��'�^1 �j�wJ�����$�´��0��X!p��6]�l����b�F|�F/#}zb�> �|a��N�f��}rB�<e��F�������(^��(���s�<y��A�	8��¥1��(*f�<�� !VǚT���:>�Ε4�W�<V��jͦ��te6i5n٫e�RR�<1�
� KvMp2�2���r�\O�<��i�R�K���&ޔ��r	K�<�R �l�0J��2"̜HB�[I�<�b�P3q0�8�H�-�Ԡ��G�<��h�E��	M&fr��{���[�<�6�9]Ϩ�q!�X%MTC�mFX�<�4�H�3"��@�ƹ/�\��n�S�<9ҍ)Zޠa���P�EJ�L��PQ�<APC��U��H��'\�%+!�D�	:���@�¨
44`�ٳ#�!�$�L9N��A�e���{6�D�Z!�ɵ1��"�����좇���!�$�,+���Xe!B����RC�}��(�L����J~�,C$�3�(���B��p�v��u=j����qO�$�ȓ}A�lc�����
�-(�L��Wt(c�\�z������U��X܇�B�td`��ܱeD��oӜ-�b��ȓ,C���!���L�h�֏"P��ȓ:�.��+Q�]��A�eZ`�ȓv����TƉ|�YBEp�e��DF�tqG*�0�}��$S�\��)��0t�$A4K�-[�x�Hu��s%�І�O��1%eX�mK�yvcL bx�0��6V�����%/�,�(5�_����ȓY��u�l�7*~��R5����C�Bl8�Đ:���j�A 7����+�$!��ֆ����sʀfyj9�ȓ.*H	f*.
M��!��r����ȓ)[t��V����'�=;�����$҂�Z�oW���.�:\���S�? (����c�ı "&ǚn�1�"O��(I�[��(Fɮ>4�8�"O&�3� �),Xq/N�+���a"O�����Km,@̓PR�i�"O� ����<O&�#�K�'x�^l�"O� �����r,IukX����Cs"Oșy ��,\�t+!��"~�"-C�"O��&ޯ*�Rp��[�%Zy�#"O�\#��[���@�ǉ`ON�V"O 8(�f�-Ihj�0�윏>�n(�"OԻR��<'BX��
Z0hHZ�"O�0����t��<(q��&���'"O�asu(:<�B� � �OB`�"g"O%Q���X4���
�=��"Or9��[�A�Je����U�"O�%�&�1��z�O��,���a�"O�GᒱsL
P��C�8�(\x�"O~Mà)ߨ� 0[�C3@b8= "OFd�cb�?f,��ƗI�3�"O�dz0-Љ-�� WO^�zh@"Ox�Y�ρ>3X�R�#F�r��Ta"O� B֤��P���DB
�!�v��"O�E�ś� Q��V1Y��ܑ"OJa+��c�܅���0���4"O��Q�'��^@*��PL]���y�`ī[6��R����Ti@h�yB���+��ej�m��5��������yhB�a2�H0��(&���	��y���i�������0�
X����y��A�K��x	c Ϡ9r�	/Q����ȓ��� !=�^ �d�ŮV�܅�=(�#��������N߰3��Ʌ� i����¾j�l�¥GԴy�L��xl$�F�����(�� �I����#q��w�A@b죱)D!�l|��������n�J5i�	�(((�ȓM�%�c�7'6����߶���s�|r�%���Y,�O ���H%�AJc��6L 1D�� *��ȇ�YY�!�Qa�Ks�3�%d��)�ȓf&,)�����:7o�*B���'�Ȱ *	x�PmGƛ�<1��'�H`���J7n��	���1E�P
�'m�]jfFP Z��0�U:E����	�'��X��㄃J��XA�#<����	�'0�k�<t,AJ�#]�]`q0	�'�N`Z5�K0"�کQsEO�5�(�	�'��yS��A���Ӂ��$�I8�'�8�a�GY9�JLiC���u�eK�O2���OD��!�'��
g�oJ5R!��o�J=�6�B�~H6�s�mY7�!��ҍc��\��E�'Nb��ׁ|!�Ť,Tu�k �@��Q� �!�DLt�b�(I���V�ϻ#�!�d��!d))�D�y�QruH��;;!�d�#�lX	Q���N�[�fW�!�dl#p�ф�
.e�|�F�۩G�!�D�q�2���L��%��K�-E�!�D�4�0���ցP�p�qt%R�TY!�d�ev�	g��~�th�7�!�ě�U��C�'��nj �
�(XN�!��"� ���Nea��aǖ�+!�$�R�N�#���A�DI	�%(!���~�>�R&����}��Ϋe�!�� n�zB�G��C�=? 1Bw"OR�gO��rv�
6,��U"O��)e'L�~���Pr@��"OΥH  ,�dym׼Nb"�a"O���f���J���|8<��"OPp�`�	@��ś����+d��"O��`�EF+i0�&��&^),z"O��u$�d&�Ѫԯ_�.��\"R"Ofu)b萍g�`Dx4��W��"OJMhSm��r�ì�<���Y�"O��CŒ�IhP	��W(U�"O�I{TM�y%<A��֖:<P�q"O�x"��8-:����5j(fѺ�"O\�г��7*i ����V'�u"O uq��L�9g �-q=�Ѫw"O^uaR��9�6��GM+��Ҕ"O�<��1F��@�-��p�"O:�[4*+����v�M>�t+�"O���bЄ��23�� @E5"OY�����G'nLy��V�\@B��"O�3���&�['��4�Z�bw"O~�Z�lثw�r�#��)I�$�#�"O�9�#��]�@YDG��P٣�"O<��f��9C�|i�FM5�V�%"O�*��˭| 4��TfH);�`��"O�8 =e�����\�e�4ҕ"O�b���;Y�:�*F���@]����"O\��P ̓}5����Á3(=�"O�	����(�)b�� R,�yc�"O�8��.��V-88ր�1;#�E�'_(�H2	��I�wIΛAb��p�')���V��;v��yY�hҀc����'�(��J9�:tРC=P����'��1��nh,0� ў[��X�'r"����Z�ru��dOZ� �H
�'��Uk��6�5��P�U*�	
�'�̳��I�vt�]3B����	�'S�Yɰ�Wc�;u�W+<~ѹ�'C ��7n֍-��J@�!�B1��'�
�+����+�()�֦�� ���'��1+A�+o�Q��6�z��
�'2��;��)I�(�u"A(y`���dڀ0�`ӷI\��̅`af�
�!����0Yð�I8,���#E*.!��=q�D���۶4d��+�IZ&k !�$ʋ< pXsçPRʌR��7!�Ē#W�`U��E-lh���鍞9�!�[� �LE*�l�dO
!ق�ʽT�!�DY6%c��J>3En\�`H��z�!���xbr�ە%��5'�h��ǎ7AE!���/����mÀ:�r��@ؔ[-!�;վ�����}�r%�⊖T!��-<h���	�c�h��п-,!�D�84x�UR�l]zL*�d�X�!�Dսq� ��R@RN�H�`�!�� ��x5�L�c�"�ڕCTY�!���T���ЅϮ*�&�@�_�F�Q�<��
)��� ���,�Q!�9�4B�Ih=�0a$L%k=JY1���rfC�	y�T�[�����n �]h�C�I^/B :�h
�G��Ԑ�l� <}�C�	�%�\^���2Ԅ!ZБ|B�8�S�'��;7�$�DA��S�N"%�ȓE�P�J�.A�o�$��P�B,VP
���S�? ���Ҽ=��fL=�� 0�"O�"�T�p �"O�ye4I��"OX]���V �*` �Ȅ�!W���5"O��P�[�6�B�X7E'OKڀ"O���,�/��%��6Jk4"O��8�@�j�d�z���L,�X�"O.���Ӱ[��e3� C7Rhk7"OL��U>��[a��,�M�"O��P@���ly犇�9(��� "O�T�1�!{�Έ�P�Q"��t"Oe
���>Hv��f�^�
�"O6���0[Р�y��nƢ@0q"O�H)��4ULQ�aQ�Z"�"OhйF�ˋ���۠�P$�2�"O����E�k*��h�Å�z)�"O*ss��7��"^�f�� [�"Ol)!T�V4΄��+��_�mc"O6 A���[��BtC���u"OH��eZ�9��5�DȢ;"�(��	Jx��R%M�!��� T�S���1��)D�|���"%uX��Ս��W�x`C��*D� Гʋ�B��6ꍶB�^$(��(D���"dA'k��$��

'w�,��c:D� ��@��)w�=J�-��@i�gD8D��� �_"u����?`y2��ǧ6����\���"'3�hhx$'N��B�I�>���s�.M�5����'d�B�I(tF�t �V��Z�/	8�6C�	�Bȼs�GI�N<�*�\/�&C�I�-�&ͪ��n��`�@�FLo(B�?C�^X�A�]6r�h��AE�$��C�ɱ9>(�f�оa�pQ���vp�C��:Vp��$���nLKtjÃ8�Դ��k�^\@6 �2Aꘕ�`bK)"06���	[�+���H����ua�� ���Qg��/0l��R"�8W��ȓ6���[�a�/	��YW-�3%�ȓ!��T{�J��OL��@i�VC�ń�u�T��bS�;�zt���V_����	ɒɈ��P�������!~>��ȓx{\�)�$=@� \B� \3���ȓ~vX�Ish_b��Y�+,+����D)N4ӷd�UGr��l�+����ȓ��B�@O�*�hd��L|�ȓ5�8M�4,�;j唜(�ZB|<�ȓ^S�e�5�ސ'����&�/p�}�ȓt�]�'���Io戫����R(t��ȓv0){�D+�^x�q��+�x؄�;�8 �ϭr��)�"����-�ȓG�ni+&�\�<����֦A:��NhD� �!2ə�X��4��"O^��r�[&�
���-�e��Ġ�"O H�%ɜH����5.GZ��u"O>4g��VI��,�|���&"O��qc����:k��,��"O�	ؑk��~�X]�����f�1P"O��Di@��pHm�3ܨ["O���'��#+pA��+A�=FMY�"O�P!�W>+J��AU*�9O2|�x�"O�lfd׽d7.�"�(��MJ^�q�"O4 CL֕/8"!�6J�%َ`IF"O,�+��:W�h����/b�����"O,h �!L0y�h��J��L��MC�"Od��E�P�$���`��^��*�"O� �%xDJH�N,t`qAZ�g�P!��"O�Y1�jӅ^<:����&բ�8�"O^���f\�XP�� ��N6��5X�"O�})��L�jb��Xc��o��Y�"OBؐ�nً!�bE��@X������"Oy[bV�O7Fp��]�G���ڑ"Oʉ���°	utD�흏&j�S"O֩�Ǆ{��a��i�L"O��bac�;?�f���M���D"O�|�A�fW�i�eE�l�N}Ô"O�99*V\ԝ1�Q�4��tc�"Of�A�f_�s��h�v�ӻ>��h÷"O�У�!�b�l���
+
�}��"O����	Vq�a[Gk�&I�|��"O�0���6J�q����6�#2"O�b�G4sBlcB㜯Z�^A�"OxT 1(
68U8h��!M�@���K�"O�$:W��3C5��v.��s��e��"O���l�j ���*�u��hQ"O�,��nώ pH�K���!���#"O�L��$�3vה��U���*z��C"O�Т�9��PS�ݶ&�x�д"O��aun�)Υ��*H\ �YA0"O��ٶ�߫1�  b��æA��1"O T�$��C�h41�.T/,6�hT"O��Q���p�������!n��-� "O�l��lʊ%�
I	eߙ���B"O��zE��'B�i׆�6���"O 𪕠O=?�X59&�E9ym�u��"O4��b웤"�|<+T��Y�B���"O��k�ֽ
@�D�qG8���"�"Of��̋Z�Fm����k|,�"O2�N�~b���@ЊB��P�G"O�T��'�9C~icq��o�΅0�"Odq��&G�?��!�̝<|k�!Ʉ"Oj���B�4W�~,��&
 }��P8�"O��;�AJ0M���F(}M|�D"O��2̋���) �G"=�ٛ"O H�sȐ)��Y�c۴09���"O|��ыM�Xتd�%[(܁G"O�'��h�.��3�H�"���"O�jvl�DGd����t ��"OU�I�<�T(i��Q6�;W"O���w͕"�&�"�޳u�d=Q�"Or}B��MN6�Qۯ�.�U"Orh(��ݲV�Ω�`oç_�	�6"O"�:�C��|�n���8���"O&�qJ-4�t �@�;��,�"O��"�IG*��=�0��-h��4"O������@�\#�a͹L�q2@"O\��GAJZb�:5`��FL֔�7"O�Y�&��!�Lz�̏�Y�Mw"O���֪�H���eR��3"O�M��P�N��d�$ĭ6�)"O.��P�]�3�̠@�,J�uXR"O�d2"�F�^|1�AK-(��w"O�����%��P[� E�vL���"OP��c���h�2p�!�Q�.	���Q"O��;Ц׀��p$�-C����"ON,��[/T8��c�'?d츣"O,�x��E!A͖ �C	B��Z�"O>� �Y�)���8� >�t��F"OrY�ECܹY������Ҁ	��p9�"O�tR��1n�Ri@F�F�T����"O� F�ug��!��l�(]�~L�hQ"O\����bH<�	�'"D�ѓ�"Ob|���	>N|�:�CA�0�R� �"O��p5�	��,$X�cɧs���"Ot�� �$9L�]H3�߷1��
F"O��:�"�Xzm8� 3��ͨ�"Oh�"CӢ!��1���W�k�02"O��Aծ�Y�>���M�(/Vb��"O�X���о?]��q��iS�5P"OJ��"+U jD�C�
�Z>U��"OD���>l�	�pdG�d""On�:A��D� �r́:��c�"O���DN߳A:��@������o[�<1@eä`�l�5mQ%~�X�X�<1	̥=])Pa��K�ɪ�f�h�<��G��D\����Aʙ0t�`���L^�<Q�K��B"�>X(���DŠ!w�)�ȓB��]�d�mJ� I��f��ȓt��C ��=�@����"���#(8�	�a ��r�O�KKhM�ȓV�xaж�<<���7�8,�ȓ�F�2D�0�:�D�9[S���5b(��O%�lNڸ6�M�ȓH�V�ϱ(��&/�*`����8�4ȣ$L�� �+�B�r(�ȓ9��h�gL��@Bi�3OF uN������ xaƆ�{�t�!b��e�`���|�����J��	��%C�M$E��Sdt1���P�>ڴ�2a˟b�޹��&����e����Ѫ���n��w"����7Y>���O�}@���ȓQ�@�bc�O�<I��T
=��(��B��R�P�+�5U��;�~5��h4��RɆ&
"V��b��P�Ќ��-��H��U/CU*�v-��b�|��t\�����0 j81���8_jD�ȓ;�^�q��ď|Z�A`1a�m"=�ȓ
gҠ��l�}����JĺT��<�ȓiR�J2�T# 796�U�ȓOtt�C��[���*r�@�w�N(��B�N��DBWPm� �g�,eD���\� $a�اUG���c����a��g���#����p�Ei�!V7,��؄��� nlaaԯY,%�`�G&�yr,ڳJ �|�BH)t�2ˤ�y�N�(-T�SW-čL�D,����y�E�t?Z��c��C�!�E`۽�y�ԜKnTD{�"P ?���XP��$�y2&�-�6��E#��.�����. ��y���%{REj�)P�(e���!���y�Ǘ;N���g�#�>��5�M��yR�ݠe���.����6����ybaX��6M�Rꑇwb�p:V,	�y*�{Y&������ ���yrG�!]����v�����cq+� �yb#��e�����aʝ`�&�`���yR�
Q��#S�T�r,�3��*�yB@�HO�d�%�:�-��)J��y� ��_�8�!�G5	rP���y��H�Ah��X2�2��欋��y�FB+1>�qb��$&L(H�C���yҨ��e����E$!�l��N���y���=yvY���	���r�!�y��J/	���T�\�Xʕ�2���y
� ͉�^7|�8��*:E$5��"O\���i� rnH�a)ɺ3	��{%"O8����e���
' ��A��"O���TNH����k6c��T(He�t"O��ٲD)7C�t��� ���;�"OL `��'dY"��႒v���i"OH���B�x�0T���S��<H��"OnEKFMĊ ������i�hiA"OB�#�J\�����NXV+d�x�"O�MR .M�/~�r�k],d�c"O�T¥��0#�ԩ���ڕt� �"O��b#Ζ��is霨v�Ⴀ"O�qP�M�4m�P�*�V��a��"OP��Q,P�z����� E�Z=�"O�ـ,s��iw��!m�=�"O��90(o�eCn�P�i2"O�@�bj��0�m�WlR��'�!�dG��x,�eR�1�������h�!�DQ� ����Ҋi U
	!��K'�̀�f�����)G*�!��E�f�f��0a\�f�� ��h��5�!��D#J��&fHB���vG�xT!�d�,#G�x@�%,P���FG�]s!�dI ��]�p��-.e�wˠ2V!�DV2_.�d��=����X�I!�d��S�T���5�"$�P��3+!�dJ�'��d�*r ~�+&D!�d׵U� 	*��<y^�!AO��Zp!�d�M|5�t�H8Z����g��Y]!�)^J&���%I�͡�޼U�!�D�Fr|3�&B�@�(S!�Dh��1���	�ZK*�I�a\!SB!�䕟2H��ˎ�߲�*�&��v*!�dFgGD G8�x�F	 ,%!�$�tA\�s�$Y0IX�����b�!�D�*�2��"�Kh+2��#%Z ��Oj��8��)4A�4��a�Q�ώ�T٨�"O��#�C�� ��Y{��ŌS|�D�e"O���ud�z�<aɥ��jo
��q"O�d ��!-R��	r�^�c�P�"O�h[�
DuB8&"�S$�h�"O�%QqkǛ�Ÿ���?&_.D��"Oh�O�%�$}���O'7%t�C�v>���L�3�t;�=�P�0.9D���W��.1����5�B�C�6D�$��a�� 莿8��PQР7D�����v�*�B�O9(& �ct�3D�	�
�&�0A 	�j��i�L7D�T9�M�AF81�K�^���ðK"D�tH�Ct�D���kա`ˠ�Ѱ�>D�ܡ��q(L���b��pa=<O�"<��ʔ0fY�5レF0'�����i�wh<	�֌^.�\�&�%O�XT��΄���O�#~�G)�@C�bC�T* ���AI�<A���R�����%Nk����M�Z�<Ia#�:�I�c�U+P�i1�M�Y�<Q4A�%%���&��K��ݙ�$�Q�<�eI�B�Dp
�7w�Z@kǀAi��8�<W�{��1��O�fe&�"��Qc�<�W�B�aʒ�C�Kۘ	��m�v�ܟ����9ᶼ"n�d:�(�Ϣc��l��
,� ��L��TKZpt��R�<93m+
c�����	�L��Q�<�1/%F̈́�*��/_�(Pf��Qx��䧀 ��LK7ts��˧ɞj��{��'�ў�SH�' d�y5���y�
�
i��nr���ߓ��'�n��P��=��@ڠ�Kc�4���'�|�[c��1���r'e )U2Ur�'��H�ȃ�H,!�7
"I�J�x
�'�By��JP	n;��;�2BpF$!
�'��q�G.%�fx��
��k�
�{�'�R��s�Ϟb�4A���֓�JP-OF�=E��Nŕ4R�����<]�u	A
��=������r���Ƅ[�ss(�a� B@z!�$��m��獗h�,�C� ��.!�d� $�|-����=!"��+ĩD1!!� ��~,r�H�o!J񧜉0�!�d�18���(aq�`��FܠY�ўx��!x�=�֦�w"�'N�(x �Oڢ=�}��AU��������3Ĵ|�A Iҟ�G{���� �� Pt:h�r1Zǩ�L�L��3�Z�B�JS�Vٔ4(U��loڹ�ȓ2�f�j�٥}�dy�� ��u�ȓ6�,LS�OE�r��1NV���ȓIª���"W^��ze�u���ȓD�D\�g
ɐ�@��ǾQ�,��_A����'� 
1ń<>��D{��'H���"N�k���PO�&s2�D���d)OZX��0)_<�hЀ	V(�\x�"OP1&#��,��u���i�i�1"O��U���,2��@�-@\ @�V"O �z�� ,�X�vVA�~@��"O��;4
s\�����[4nIJ��_�|��Ճh R�`����R�(@ph)D���p$��Q$l=2jV�6@b�� *ړ�0<��*�!����F��jкEG�M�<1�����`X�c�@��L���I�<��jC�3yr�9(H=>���*�B�<�! �lY��F$@/tY��WF�<Y��X�NyR=�b�Q6�Y�<a%��;�T���M
�]9&Ha�<Ap��+9�d��,�;�|D1I��h͓X
�x����
[�2#a��+�Z`���4<��/�m��$��j��K����ȓ���Rק��_i)��ֿ3���ȓTvF�`��	/4������M�P��G�ȉ1G� �aʖ.X�V2��-���3�	�&���Xpd��ఇ���d�P�=e4e��J���|��
�4p�B@9hɈ@��gW�5�Q�ȓ ��Q$�Dy�Bc"��q�T�ȓT�n��UFD�AĂ��t��iꐆ�3�`��L̿s�F���!�.N8����(9�d�ž'�,��+H�I2���	�x����Q8"�]W��G�B��'ў�|"����8s|Y�=K	��Q�#�F�' ў��1^PH�I�)C1pW��nQ���ȓ
w2�yJ�'"�+#�A�:��ȓo�\i��JR�9F؛Pe��\,��ȓ��䊖J�P+bp{qŏ0��D{��O�8�n�<�bL����/�Ĭ1	�'l�9���Ɓ+Q
�3��J3���X�'�bܲg�Y�
 �֩)f�L䙎�D9�lt�
�#��k�k
�F�,�!���l�)���␺kٌ2�!�D&,m1���wQ��ã�ڪI�!���
[*��䉂-);4��E�Z�'�!��ͩ^
<����ژ&� "Q�Ŵ!�� @��aIʂT�< "�EM�$ȕ"O�� %��0Qs�tI⯋�0����"O�����UY&=*4o��`�c�"Ot�bEƎ_I6h`�����""O�)5i=5m���@�+� �C�"OL��W��X7�b�άIO��s6"O�R�m�-�����&; J�"OF�K���z�j�F���(M��"OnXk��Uh\�s���"Ac"O�\�#ʚyO��q�&��E!nx3"O�X��I�`��t�@� ��`"OXc�.� S��Щ�9N�yF"O�`˒�ݚE-:�[�DJ�3c���1�A�'0�*C�6��a@�=DD�b&�!�Dy�g"W�]�)���4�!���@��O(arxcB"W�m�!��D�NE��+rTX #r Y/N�!�d�<k�@�r�o��{�~1�R�!T�!� �jNx�6h7#�%��Ί/�!�D�w�I���oZ��#�޵!�!���$(���&WJ���-��k*!�dG;��ae��_�����,1+!�DG!|���G�>�`1 oт,�!�Ĝ3X�^]P0*S?�r<��#�!�DͶw�	RW��,|�^8Y�!���VF9UK�.&&091�G}�!��;M|d�7Ϟ {pp]���/	!�����ѷ:"�I���=�!��-���X� �1.#��K
-P!��>W�y�BdQ��l$����3'e!�$p%{�-�%�Ӥ_��З!T�<��O�,N+�$2_���傿>P!�$<R�𨢤�%JC�;���,m�!򤞬�N��VN=*D� 2��/t:!�D͢wGnA��Y�b�Q��V0!�N�?G>I�#��L���Ұ/P  �!�'M���oã �Abvo˪@�!򤔕o��%�
X� �nL��!���bŶ��A�Ā#���H�*I:O�!�d\�Hg�x��O�� -���L=Zj!��W���;��Ǚ��Dj'O�FK!��NZ]\�Q�U= �LX1㍘;J!��H4_]z��5	ʈ)��]r��BL.!��_b8��PdJF?{�-�s��;!!�$M�m����"�P i^�E�T�_�7!���"&3��)#�&D!�h�r�'%!�DR!k�<ժ�,���8%�P"O�!����r�0ӄL�+<2��E��O�!򄁚Y���谮Y=g�R43�A�!�1r�����)\��
�HӁ�!�_6a���3�O	C�6b�H4�!�
I�$�Wϗ
�fe� %�:�!��m -�4 ՙMfd��Ȇ<�!�½3������E֥gBA�=�!�D��VL��1с�<N�T��&�7�!��Uf�.9�cE�|:�����#%�!�� Q58#ŀۓX֦��A�ќ/�!��A�%�^��ga�=.(�Hi��^)�!�d	��.a�P���i⊒�U!���+�Lya��["����WJ�H7!�D�<�6�� ,-���r�h]�Y�!�6D�tC$�3���J5ő�j�!�D;9	(�k#-�	<P*����Q�S�!��׾5�<�a�_�x=BQ�v�P.�!�� ��ʆ�[�a�=BSJ�eS�"O�`���E�Z�б��5<t���"O�%[���	) �i�,�>L4^Mڇ"O�PRׂʉ���qŞ�1�b��"O��ؕ*�&;������� %2�"O�`{�S\(A$>l���
�"O�q�F�Yr�b$D�&�4�X�O���b�Չa���Bċ��v&��I(+D��ԢĻ6�pZGޓM*�Ec#�)D�hB��]A�䬫u�["z��l�w�,D�I���,�A��*"ϼ��d/D�h�)�f�y�֍J�<E��
��-D��:�^�*8Rp�$��R<���c�0D�01˔1U@^���'�	N"nu�Pg-�O��'Au!j#ꚓz<�U�56C䉹G]��q�/B�-�����_�JB�	�,ȤMS�%�)Ҭ���
�]�B�	�/J�!�e�a*�ԫb���	�B�	�f#�ez�� �x|��RBUB�I�`���Sp
H�?$x�8�ն��C�	8d��PgƟ/G�{�	�<G�zC�	�C4YA��J�t���F��e��B�	ٌdY��vb�ԓv�K�,CXB�	�Cx� *�Iϲd��� �RB䉐:� �X��3f��	����B�4f����dʈ��PD��Đ
�(B�	�m��M�����#Xd��� �-d��C�9b��8��A���ģ燀�~��B�ɭ���R�|�� �h�7a�C�ɭ8^:!�G@�_��tG��)�C��k�B�8��� cq��*�/[�C�ɊM�|j��n��,�@.И0=�B�	��V
���1GA�P���y�FB�I#RErб�B�!nKpa�R�ߌX�JB��::vdq��J���3��:%JB��?3��!����s�@��N5V��pD{J?��!��!d����ɏK �X�!=D��Qʃ�(�8�d�G�G�@�@s=D�����	�]�:)�1�K�
:H���'���*��P��4�	�z�L|)�'�H|Q5��<�^��㛂^�V�s�'#
��`I�^�=�Do�*j�&y8�'�PD�TdՑWSB�C�^ɦy�ʓ`���f��S�B	�`�.,��ȓL98,C����Җ�`��m��x����*qm�� � xR�ٝ"���ȓ1�LQt��b�ģ�'�H\���Gu�X�f)�D�B�):Lلȓ�p�Q\�G(!�%��ḧ́ȓP[��ș�)hڭJ��Y�:���_�u���ÙMhI��C�UD���J	E'X*y9�B#IST�u��"O��Q�
T#@[�R�8݆���"O�%
Ш���@	G��$����"Oԕ"e�Fwv�"�6#���c"O�u��Ċ<E�!�p���e@"O�C��K�R�< ���m`���"O�@��b	���\+���:Xܹ"O���.J"Ha8U
`Ep�xy#�"O���sO@�N�}�g .W��L"O*�#u�7RHj�*w/U=\7��P�"OН1qM��;����A4��H�"O�L��fh�YS�슾1,�xW"OH�[s;S�p �)�+1��9��'�!�� ��Z�G�0�0�z3�J�,��@"O�ce�ً=�����	�A�^3�"Oe�
�}�E��H9#O$T��"O�y�L�=��AC���\<`�"O��0
S�����w�D t�T��"O���HX�j������3�����O�)砅
Z;�TA�'�<J�@C�>D�H�Q��mS^haQ��4k��!uL<D���ӪR	k������é}+H�6�>D�p*�� &U�0��C�A1Piɱ	0D��R����B踭(�&�?�j�Y'3D�S�G��Jv]��$�"I�R5���4D� +�I+\��F�Fvv�	�k34�@�pd�&�TBW!r��r6 [m�<�����+��H����r�<)��ܷJ"y�ĉvz�(6D�C�<9��I�L�L�r��R������Z}�<I&��/C+��"F̈��~d��)r�<1Đ�8XM�b�A#d�����C�<)��>?�jp���� ]�Z\(qiDu�<1��X�`W̕��%�A(�'s�<Qd�ʲ$.����Mhz$�n�<1��6\W�ܩtu�乁��n�<Y�Ӻh��QOX�?J��#�S�<I�XK�d�B���L����Pu�<��՘=�" FC�p�a�'�Ue�<a5.6C��:
�-_pxĭ�c�<1C'��#�,ʲ/��Bh(�^��ȓ�
�)�c�r���ŉ%<�Ԇ�!n�i�:,dd�hi�r����3�Mx��G�1��m �.�7T(u��J�RU���]�)^��Ɇ�1n �E�� <t!��S�R@,�	$b�,[�����Oef�� �.;FX����ݠ5wց��Q��ȃ.P*FD����.��?Y���~j��$H�B<��!ۣK��� ��C�<I%BX������g��F�tV��w�<����餈��NO<m��3O�{�<�(Cx����Q[�N`J|#v��v�<y �(��;��&-rm���u�<��
��&�M9��AK�  |�<Qa*���H��D#�p���z�<qg������w/��M2\p���z�<��l��|���@��]L<-�.RA�<�F�D_���0A]#�� [�CBA�<q�E��;�`�4�Sr�n����e�<c��5�2�3�S�6X8l f�]�<a�톯WW�D�+ BY˛ڟ�F{���7��̚�I=�fԈ2#"9���hOQ>r�.�.1ܴ�BGȞo��WC7D������N�rC��yl�4�v 4D���0���<;.a1FF62?�X��?D�dP�X	�bCT�4I��'D���K�4C��pSΟ�;��܊��$D� DX:.,�AÓ�� ���7D��"-�8k�d�V&F�`�� ��4D��zQ�O�^!�-Æ	�;�|C@/D�b�K�cح��b�o-���I'D��ڷ�U��D=b#@��>O��:u )D�|x��"R��<a�=y_,,�*D�X)�eW�]�ȑ�F8y�pXa)D���WE5[��$G@Aq "=D���� �-o��0f`O3%m9�m-D�|1�̈�59���j��,��s,D�� B�ٶ+��~�J��$��V�$��v"O��w�F6F6���E����j�	D"O�h0��9BߎI��ghGb$a�"O^�T��Q�:	x��ϭ����"OvԉcA/F<����X*i.�s�It��)��M������ !$Xl��6D��b�2��x�5�S�,��չ��4D�d��6m�x������5J��2D���$ǖ�TР �Ȅ�ƕU�0D���f�8�@˶IA�u��"U,/D�dkUpeL��]%:�J��H"�Iqyr�'>E(�)� y�8H�D�Y�I���!D�d�I�Ab��e,ֆ=���i��=D��Q�D�!��uԐ/Hh�9`�/D����E�,$<�ՠG�0�|I��.-D�|Y���&v,�I �B�~U*t'!D��bA#�:�<��a��(��g!D��)��2mШ��m]?I�
�Wh=ړ��ؘO���e-վ?�$�@ga��9����'~� ��^+K��Ҷ�ƨ�x��'#�y�'+U-]�Ɲ�v��'M�B�a	�'����#G!hU�@���СEO|���'�](`�&��!��&>@�x��'�B�z�蒍%����	?&)��'M�A�	��y��M��7���aϓ��d&?�Cn��G��	A"۰w�<�aN^�<��Kj�X���O�rP:&�ZD�<�͘/"�~���o�A�6���B@�<a2ɞ�
14���$� )°q90�r�<�E@
Fj�9QR�R�]�8���X���IF~"%�kq��ڣ!Y�0�����)�y"J��V���ǻT���k�*�yB��7n
$['�S,s�LPd䝖�y"o+L͜TZ�B��J�
t씟�yr �%O��!x��!8��Bs��,�y�j˜=(4ه�E�� !#��)�yb�������*�}�ͫ�섛��<I��F�qh�BT�A"V�@$.J�.�!򤏬k�� R�HЙ�l���M����}��'���r�&-h��4�z0E8�!�ݘaq�eag��;X�.��&�-J!�D�Pf��'>=�ցJKC�!�TC2�b��ݷ(�Z	�iX4�!�DF�!z)b�)F�� Rf�0]�!��@/���y� �*v�0��٥j�!�D)�Hԉ#䅢@h���d��W�!�X�K��-��KY�D���1!�D�5lM��#џ-�a�7! "!�D97R�p�Kǫ^I*���aǀq�!�dAU��0S�� T<�4��A9?!���dv]�5� GM���/G�s!����0���`͚��fB;!���u��X!��kA�-Ĝ_p!�dÃ�	j4ML�[�ع`��7=^!�䏄d�|Q��32R<��b�<m!�D�8 ��(P2�|HYԁ 4s�!��Ч����`�Y?>A���j!�,����%�j4�X��Ӽ{
!���Z���c���;}�de���)P�!�<"�*$�ф'p�vՙ�n��d�!�$O
&���Q��-����@�ߖE�!�߀A����c��a���,�5!�DC'f&0�*��l+�jE�U!��-#��A�`�	!Ҿ�j��@H!�� x p���i+`$C���o]�Qڡ�'clT����ہ��7RR�2A�5
�џ��'1�B-�f��Kzm4!|�A@�"O6� a�B�"�4U����j@�5#��'�ў��8�<�6m٥bNLy:�k\�D�C�Z�<�0��D�q;qo��jآ1h�Hq�<���p:����V6N^�����p�<Ae������b��r��	��/�lh<ACȎ�Z�Zy�q$�)Y�-�����<ш��C�u^Z X��oL.�/άh�!�XB&tY�H��%?�yc�F�a�!��гh.h��H�*&:AI!��RI!���g�����S�6:Tdw�ݺb1!�Ĉ:G=(xJK`5(@[��]:!򤐵?� !��@��]��0!���5 !�H�%n69���A�c���`G��F3!��i�Y��ϋ2���k�	��O��$7�g?i�/I�i�$8c��4քYR�j��T�<�'c�*��X�� �/]�I��i�'�a��k�3_��-ҁ�[%������y����p� � ��W���4BJ�y�ƾ��#��_V����@�yB�O�B��@%M�_�H`�!̡�yR.��I�>� �Bֺ&����֧�䓠�$�Or#~ʅ�X���g�3��2#+�hx���'ق�i��V�fiP�I��L�Z~�P�������S+�q0�� ��f�_- ��ȓY�@1�"�MŔ𻃥@'�.��ȓK��P��)
�,�d#B��VIN=��c´�0D��}��a[gKP�,l*�&���S�Sܧ�`h+"�A?$,p)�G��(1D1&��Iw��q�OZڹ 0�P`�r]K���b)d [�����9U"�@(�R��i�*nB�)�*�|00��u��`�&��@\ z
�'���p2O�h�T�1w��7y@��'�l��\
��|�L�Xih�y�'4�<�B'׺h�,�3UH*N�l��$&�N����1'x���(��x��L�Y������&��E�4e�/��`�g$K�L �E@�yr�Z1'A�תq�� �T�]z�I\�����`��|�u�'AA�,��QI�c7D�d��گR4(� ���A�(�Tg4D�X���G6�Q`�ٕ�Tc�0D���J�.n l�5O�:I������,�It���S�K����3Lg��B+'i�+�ivў"~��䋣Q�D�����:�2����H��>�O�R2d˦���"1aK�Q����IH�\p2ğ�aG��5J��Y_f%�(8D�d�d#��t����L_ F��W�+D��Xp� �{`@\�&\'"���%4D�$�� Ⱦo@B}x&�[�8�3J1��ڟ�G��F�S�f���MO6����Bi��e���9O,)���$|V遰�B�!�5�Iu� z1��2 �㳃��l��"eG>D���%�**�*�I��չú��'D��{S��\�����U.m�¹۱�?D����ܑH%��r��V��	��'�O:扲\�4�iP 0�B������M{XB�I�B�2�KB�2�x���oU�2PB�	�X�Lm3��LJ�͉���5b�$���	p��|kS��%��� �O;#�68y��#D�@�/��"f�æR~lDZG`#D�� e�D��t}��$�V��\{2* D�h����1;Dfq�g�twz�x2:D�� ��s#G�u��q+S+Ư]�\dK�"Ov���H�2}.�� l�(�5��"O�8�՘{O�D�P+	�c8�q�"O�R�(#�V�s���C���'!�8-R�Y�3�G!'lF8س���\N!򤅠Z�R����Ԃ[�P�AÕ/0!�D��6�M���@0G��!$�ҥV-!���gÎ=����_*A��!�
�!�$2'Hb�B2��5E����F� �!��"�-q.˺X~m���64}!�[����h��B")��L��<�!��3w{r�KE�BԚA�sL� 	!�D |�*��k�#F�2�� kC�\!�B6d[�(��`��J�Ds!�$��_�e���'�
��u@@%7�!򤅥V� �y�%�\�
���ʳk�!�D�%|���ǉ�Lz�@�K�D�!���uf�)�F�e � �-ȧ^`!��
0t��Y��E.o��|x�kL�US!��xy��Ydț���s�(YO!�@.\Y~8�� ��!���c���o0!�D�y�!�EՐ=ݪ�w�Ç('��1O&]с��	�\��eL5�.�aq"Oʹ*-M�T�8�)�Ɇh&�۶�|�)�S�I��<r�G�9drd�E�!X��ʓ�0?т)��q���3']�-<Sw
�V�<7�[0�X�a!��=ܬ��'�n�<I��F-tJ�PC&e���@����k�<��(����O��lht$߯rJB䉁S9��7G�%J�DA坆w%�B䉌3)$�+��صE"��1a��I��Ob�=�}ҰA�(L���Cv�7+>`�t��u�<9�/��ܖi�[�*4 �0��p�<ٔ/@�dE����Gx�m�ҭ�d�<�昫G+�LYb
{�����|�<�u�N��aï �BYj'�x�<YT��E�1;��ĝ-y� �q�<��F�(�p����{���@�xy��)ʧ�DqiE�F+]ȢA2���	� ̆�l AJ���Z �q*aj��\��i�ȓs+��Km�m�<H2����q#ZM��H��T��;|l��`È6oZ���
�0�����%O߂����^�y�ȓR���I4��^1�#�	��fp�ȓ�|�	G"�"���1V��;?~���ȓr$�� ,�1`��)� 0{` %�0D{���B�t����7f�9zQ&�Ԟ�y�E�3$*�Сe?I��͓�yC�-PfV4{0��"�Za�p'��y2HH�S�e���Ю-x�a� 
Q��D2�S�O���)Dm#^I�P�m6^l��'w�9�p쇳{5�A���A�T~*�����_�$�*L�S,��

���B�w!���K��!$d����֎Q�y]!�x<�,("���4���לcj!�ьt`�b@��"r��Q�An>!��̃U�P�#� ̶0��֏�+�1��FI�-���1��,*�`�74̇�&� B��MĬA4��.�l�����h�-���m:��hw�m�ȓƚ)��ގN��p�D�?J���ȓS����3c�?Yu�x��{��I�ȓmBm��e�
<؀��Ga�00��ȓ �����͛��\���-�H	��S�? z�5nJ !Sd���i��l ��7"OZD��C���s�gًO�l���"O2-��%]�f@D+&$\<jݖ���"O*�����c�"��sԌ��"O4 �֋@g=� ���
�c��M+�"O��As̓,�Q�g`�6h�]x�'sd���ʙ'�z,Q������'���Ӆ=M.)�c���@	�'���FV59�(L�6�Y�c{�]��'t��_�0��� '���X>t��'T�C���y�؈;Vhݟ���)�'��! �˷6UT��U�^�.M"�'}��K�T�R5�\h����i��'t���R�XN�|듆�sa`i��'v��@-�7 �\KD+]���T0�'�A��e��d^}Bd%�\�q��'�h@Q4Ú�0 ����%�J�b�'��PZvk�!t�0Y;�/�z蔡�'!f�CȄ�`O^��6-�]��h�'��4���	^��H��Y x	�'�4�q�=��5�uD[�C��UK�'�@�C@0"�}�&π�䈪	�'#PS��7D������
��$B�'̸@kQ+�`\4j��ІXa�R�'��(¥gQ0NjD��OU����'N�rF�1`&�qcc
M=f�
�'����O´19dB�+�;"�#�'��[�D?J[$xyP �,(�����'��z�M�^V���Ћ�x���'��cVO #(�;�,��R��	�'�B'bʾ-�HYX�� !M�A��'�89��6L<���&��Q��'}�Pm]'"ۦ`Q�OZ�^�,�'�(��R�H�7IZ�+���	WF�	�'�h`�3�ɱw6�ڣ��<�ruQ�'�}�!m�4C�:P�,�..�8`�',��Q��tVt�1�Z-�(H��'�����ʔ"{�*AM�)\!��'�����}Y�]
�ADO�h���'hl��'�E�)��AEΚGf���'�`��H��!|~!s��ڝq����'�:�/K�G��e�Ā�$�r�#�'��	i!Jϧ0$�Qq��W%��R�'i�X۲k�%2^<H^._�@�'zQ�D�ݹ�T�جH^����'�p��b�/� �s�aW,���`�'ּ�ر�T�~L�ѣ2��C���Z�'��!ʒ9F=��ɀ24JD��	�'	ޥ�d��=�N1��A�%��j	�'(X�"ʯk�]�)�^x	�'S]b��W�$ڣ���d�h`�'Î�˱�L�z�@� ���/7ǆ(�'0^�K�g����m�&-L��B�'�Ҍrѧ�A�М#!���T%X,��'��h���հj���Q#_�7b���'JM�7F�#{�@��ȸ5�z@��'�����E#2�
 X��ؚ12�(�'c\l�u��2:1���sS��J�'a��G�B
=����m͍h7�(�	�'�P�k�hP�O� ��V�!�
�'���#cX�uo�m���A�{�my
�'�J)�ԠM6��1�����]��'�f<A��ÑG5:��@�ܓ�XB�':b((BC�A7r�!�+Ag������ ΅�ժ��l�� �Fr�$#1"O���CʄkLm0p�D?8%�"O��	�R:R������7�Z�B�"O��갮�}p,�*��!v�$�a"Opi�_�<��	A�vԌ�0q"O�Y3�
v�F5��I��'�*0��"OJ�Bc��'�∡�F����Ђ@"O��xϒ �~�8��о/�$\@�"O�1�N�v�&�PŬEjJm�t"O�����ΉzxպRiȄdr��KP"O�T:��>b����.X�Z,��"Of@q��
s��� խ>75Ҥ3�"O"���,^GF��0��>̫�"O̀���M[R�8�+�)�)F"O�!��J� �͚0M�4��C"OJ��`���#�l}�$lX T���F"O���C�5	��J�*ȣB�u�U"Oh�4M"�`,�)[=g�>4��"O���@��{I�"�&R�M�xm��"OX�$�J���i�ƐVr�� �"O�Lj�O�� ���8�� �gZx��*O
�FI�?ڽ CC�!\6x��'vޥR �;rwz���nջ��1��'��I�%O�=���o��'�n�
	�8?[� 	I����0�'���GEΫ'id ���T}A�;�'P.}y�B�{��y���.t�Ь��'�A`cO�
L�.�q ��iUh�+�'3���G�͸qْ	�L	�T��'?H5�����$d0u���w�ـ�'�0��)�pZ�q��D5uu�A+�'D�Bō�T�z�y̕�l�Nu��'�B��JC�S�q%��o�t���'��P�U��Ƚ�T���i�H�'� i���ZTtx�/�f	T5��']�Cv��Y�z�����Y�hL�
�'�:yk$��q؊u3�FT��B
�'��a�g�k��8ug��~����"O�k��	��IiS �>A��0'"O�YD,�(g:D�ͶP�8Õ"O�Y�0��+?�P��6�C!07�`�"Op�J�OA3yL��I�'d�hA"O���)�1/"�� d ;~�^q;F"O$���7���## ������0"O�:��n�B�aVdB%K�� �$"O"t#0��&��xӴC��c�,aP"ON��f�:[9V�i�Ȕy+
�p"O��q���R��eG>����q"O�Ը�Ão߀�i�ȗ\w�h"O�0�P]����`;�z�X�"O�0&-�p1��qC-����5>!�Mu��Ԡ� r����c�ڽ �!��O�rP��t��GVh#4�K�X!�$�5'�Y�u��/F<�a:�b�j_!�dC�u_l����* ~�a��ژH�!�$C9�(ѹ`�8^q�ej����O�!�$؛r�\����Q[ ;��?Z~!�$لwv�蜼4C�#��1a!�U��d@��'^X�pҗ���@B!��8����jH�g<v��ٶK�!�_+HV��eC�56&�b��r�!�O?.d�퀢/�z�f��7C�7�!�d�VW�<C���
]�t�CDL's�!�D+y(���+̎ Djf�V�m!�� �9�e'�.�ґ���K]Ǿ8C"O��!�i�Db�(Z�hCg�H��"O��C#@F�&����3{p4��"O���GG�"$M�P���+iIV���"OT��T1j��ӵ��1C��ڗ"O�HՂU��4�#6	D�K���2�"Oj|�'[�J�;�C-l�	K�"O�y��W?G> �0��"Qb䰨Q"O ���W�FG4���YY~�*"O� ���s9��#���,ʴi""O�x��@�6�J�� ��of�*�"O>���˦7���I!昲YS����"O�1�R˓�(],8����>_����"O��@�[����Ѐ�M�<`.�x�"O�YS��T9,�Ɓa���~��DJ"O���eM*[�0�r�F�P@�"O|��tcY�H�쁱ca��x���y3"OP�LM,.-�e8�o�5>����"O"�yT� 9x�mp�H�4zy�u"OvB�
+~r4-��LO�g%r1@"O"AB��k�ư:��G;^��w"Od͠CE$6�����Q�QJ�Q"O�hA�C<�L�6jǝM ����"OF0��F ,{��(�j�@�#�"O�[�D�m.�l����3"�Ԑ��"O@�c��[�$b��`�9/〭��"O �E��<���r�<�$�RG"O�����Ԛk�H}1��V�'���g"O8�B��ɹ9��T�b�� t8d�
�'�
(ac(�|�DI�h
����
�'��嚱�̲!��(i&KJ
~���
�'��D
�bG�5�.i��K�+uT��
�'�����ԁpU��C��(4c
�'��*Gk�Wь���'� 	3�}H
�'.����	Q�\ҽ֪�P��P 	�'���4~�A	�ؠK���'����"�;�����3L�\�P�'� q��D" K0�<jX��'�(hD�U%$��1ɐ��,�ny��'"�yh��_�$re�g)X� �]��'��ѱB7=�}3�C4 �P9�'��o2}i����$
��S�"OP����wl�y3 �!p��#�"O~L�&�ʎ]�p�B٬r��E"O�j����9����iJ�H��"O8�����
D͘3g;����"O4�1�#zn=#�+ײT/\$r�"O:���
˖	��$^+}\���"OF!��F�I:�EYq��,}o
�e"O���5Ō<}�PY�h�U� �"O0A#	V�=Ǵ=ь��K(M*w�|��)���BPǅ� �a�-H:@��C�I� svi���S9=�n���MJ�rž㟴�鉱z@��1T�ۑ�0II4-�7�v���>�mN�S�~�� �FW��᳢s�<!�EZ�5����r�Ę$�AX%�C؞��=��LEٸ@�QA�Y�u�}�<�5�M�5���ص��r�
�Ўy�,����2y2�EU� bp
��c�Z\�s"O����n�%�F�U���+����5��{�Pj��;��\	7�,-�,��Ū.D����!�Gj9�h@+�
�#)�<�	�$�nq@�d�(Q�H#��G<�!���A~B
�!%"\�У;R�<��E6���0>� paʁ"©�R��<�8��I~�'W�8Op�9�΋3�V8h`f[�}
�U��"O���,�3���EJ����V�&��?�G{��зɈ�!c�غF�`!e/�c�!�Y�pa�F�p2C�ؖ2��d��?��{���Oܬ��
�"^�2�h�1�"O�ui	z�`�Q@߷EU���܅�ɗRVيs�Ӷ?5�����x�B䉻Y�$�id눤O��IV	B��a`zp��A���y��[j�㟄'��Dx"n�]p�a��Ѷd�Pp[�U���x����`���nV�)#ŉ���'kў�>��&"�	lC�azQiHBij��h��tE{����,\����o�+<@��$OK�5��O���dLOBH��c�,+=X���ˆ%���0>y'd��mzː9	�Zt�@��PybL��	-��!d??ߒ���^��yrC�4�<]��D��ۉx��Y��X��d��@��}��d��UX�l���S�$R �2[�*�PB�=Xz,%�ȓb#��a����Ph`5�ǣ�8Ȱ��ȓJ���lB�~*$��`�`�Ąȓ>�Ʃx $ՊAh<��oYJ�Q��	H̓%�3q�7S�d,��/?t���;E�Y+FV*� ��Ѣ�7-8��ȓG���`'��?]���E Ej衆ȓA��qu�_�Ěd��,D]�Y�?�	ӓL�@89I��q:�]�v��l�ƓP�)�Nz|�����<Ȳ�'w����?v/�TQB�U� (#
�'!�p �#����أ��u��t"�'?x�Q�D�t��!Ȱ��k��Ɉ�'�di��'K��1�d-�S����'�U�@�?~�8��[�_�1yӓ��'N���C@�=9̦�ʐLK�);��b�'Al��dc��"x �Q3��\I�'���c��Gʤ5�c�=itq��'>�P1�$J�R�ٵ⑈]�p�ܴ��8L�)�	.nZ�Ȭ��C@ފp(������C�	ͦ�� E@(3���%���>D�Tzw�["/���IQ��x yr��?�O�OTx{✠=I���(.l&��t"O|R�#�@�p�2*�vU�1)�"O�q�U�a�Z̚rF&4K��c'"O2x�'BZ�_�D�s�� x\�k�S��Fy��I+ix ��l(0���E-_�n�0���X/��	��D�EKo;�\�s̜�#-\B�I+{���C�D�5��x*&eX�[%&B��*2i|E���J/X�bE��\
2C�	dCz�Y�GQH�P��U ē@&���5�)§S�^d ��h��\�C�Ƽf�8��{��<��#�,iS2AX��>����w�xbk�}M�V��z����u�&R�d\{��|�z�K�� c�<IQEA�iX��"���`C�h��<A�E�w��u�<.��("�!\6�<ゅ�#(�T���u~B%��rT1�F�Q�[��DB2����#�p>	���$p�9;f JE.JP���Dx���4�y¢R�d��h���ײ�(�y�gNc�"0[a�� =�2gX2�y�
��<���2m�#7��p���F��y2%	 <���!�*��`��	ǎ��y�G�&A>��N���F�x�艄ȓG�*Q���8z����Y]� ��>E����S$p�ǀ�}+8D�� ��z��J}v	ۦ�J31T�%��"O�T҇'�zE��*g��eE~]�u"O�̊�NX\�&��+[9_�X�"O��&�	lW������JK4��ᘟ�F{��I�/���+V���e���e��6<u!��1EJ�E䌾Q�\mq����i>ў\��	2x@��P'm�,���4{�B�ɂl�>��'	Z�Pd(���]�$B��>��Q�^*|]���aGB*�*C�	0w��)%�_�G�H�&F�= �B�.������k�v�a��ql�B�D!r���b��:�t X�MɯzC��D�*%ce�A�j�Eb
2d#<a�xݜYg'!�E���7N���j����t*��R���C[# �ȓ2A���Nّ.UڈI�(؃+50�ȓwd�S 蟗dD�y1'�G�Mh��Hx�����������G'��)�ȓI[t�JԠ�*S�٢d��7�m��Ip�v�dBjD�h�
h��ݟ=��ȓ��2�"X�qnP'��Dx��	k�
"�̴h#J�j�u!�KǱZ�hB��5dhb=)W�J�^gb, GőA��B��9�\P���M`�𤳆�B�X0Bb��D{J|㥘e������J�����E�<I � 9XEp�F�x��c�C�D�'��r?�K>!�M�5ehީS5���J��pD���=��A\��a /��x����[QB��'�Is����6w��y� ��Ib�͓��� �!���ִA&KI�v%s3nB�(�!�ċ�`��\��0AؘPu��	8�'(4�S�C�Gr��d��b}�h��'%8 2�rp���lǼ[10�����$��|y��,�!FNȨ��K;�!���\�z����K�_.���A�!�^�a1�] ��#6!̬��M�*9!�x�p\���[���c�9�!�u$���.H	(���;��'ў�>��׫3�D����V���8��	q�<9�ȓ!D��d��Ӧn��]� �Bx�<	�'��E_ؐ{�k��Vs�� c
7o�-��*H��Ω>��pv���&F���'N>բ��)�,�YrK�T[
�Y��Y�]qRC��(27�q�5(J�^:��q˓��&C䉻�$��h�TMH��%�ƪ)	��𤽟��=�Ɗ�u��`��$`N	�Ș����2X�`���`�E�b�C? ����=96�3�S�ӕ4R
�!U.��P6(���.Z�B䉁]n�\���#v�R���'Y"=�	ǓN.�|�dbܪDSe um�-����28�IP�ٮ���k��\T�ʈ�<���)ǲH�b���>Ȳ	��)7�!�D��|�@	9#�� ��鋒��)���x�.��i��N�x(hT��䈪�l��X�!��4_h��@C�r�$��m}4@:���0Sv �r�l߷&�@ �ȓ��y��k�V� @J��˺6-�ȓ5�&T�>����M�H�J]�ȓ|�&AH"�$O�~m�AΊ��Fu�ȓR��d��� D� ْ���g�l�ȓGbpͱ�ĕ����AW�
��D�ȓt/0�YSfT6VW�����}�<C�4lQ�@�%\^"��⑫�(ɂB��8BN2�J��ܢ<��@qp�H�`'�B�)� ����]�+_���X9��-#�"O���A<2�V�� �b� u"O���Ȇ_�Zt�����*V:�b3"O\a�2O�R2F9��f�)H�r�Q�"O8�Ywc_3�:��OE4��9�"O�|�!&֋L�T�	WD�L��]�S"OHу��θ�}8CeӐA�X�j""O@0���C�MPx��L��
1�w"O��a�^
��a�E܊ t��k"ON�r���C#�<�����`�@�"Oܨz�$�x$!4�͡M��e �"O���pB�P�@c�G���aw"O���C��W�d���c��f�P�"O�]�b�FVX� B�=-�nx;s"O�Wfң;�d)wbF�,�$	��"O�P�e.�ʘ�$��1z̍ca"Ozm�Ø+�@���U��)��"O�ՙG�����Ǆ��#"O(T��BF4G�fE�+ܱfhN�#W"OxM�瘇E� �r��դMK��[V"O�|��� <�,�U聄 2(�4O�0�c*�
W� tp҃@�fF�@`1�	�j*'�G~��\���φ/�0A�'�i
�iS9��9��R;�Q!�'뜡���M�FΜ��u�Z�[n0B�'|h���!�I��n1 � a�'��wJ<��-��!�:�z�'M��R��ݡf@ni��F�:�D��'oB���[:<�9��� {ۀ`
�'��T���Vn�8��ď��u;���'���{�
'd�꙲C�U�Uب���'Ϊ����;ҴQ�'JNR)K�'��=�6�'5-:�K�Ó8����'DB��-H ��`���>}�"�'�N�K�CY�`4���G1#�Jh#�'��BfI��!�$[�#���'5���@K�l�"K�	
Ո�'� �S���1;sPy#P��8Y
��'?\̪b ��؜�J@�D7�$ �'��ib+���9wbS�&�	I�'pN��m~��&i��lrV�	�'?|����|`e���M����:	�'�
%��J�;�pe WE�?.���'��,������`,b�eLz�t��'t�	��hb��)��*B���'��`��-V�.�B����68[>��'�0K��;R�!��Gľ2���
�'B��˔##\�( I�	Z�[|j\�	�'p>0�k��&4DT1�X�K�f��
�' P�]����l�~��q/R��y��/iJ�AG��YJ8�sq*ɶ�y���
w @�0�� �HS�ݧ�y¤
5c�$9�T�&� q��F��y"E��.B���c/vL�+D�ɶ�y�JB;^xڙ2�)Y5C$����Ǉ�y"���­���o*�(!P*���y杳���a��	f�p`	w-C=�yB.�-T���KA�&,�F����#�y"��
P֩�$�=Jf,\�e¶�y�BY�~��W��G�J4�T!�4�y� ��|�h��=E��n��z��0�J@�1/�Dem;�ym�/)"ES���A"��9uE˷��d��lG�`V�4LO��"b��IzN��B
�t�.�S�9O���������4�J�u�,�{���# ~j���A�Fi؄"¼gp t�V�'lOTP�_,*|�I ������wTB�+�A
 sZ|�`��?�O2�SfOB�R��A��� nч�ԣ=.��J�S cw�%q!���!%��"�F|H���b ��K
�`$ 48��AWER6�  b�T������)��Y���$� ��CD�r?�݊�iE�e��k��:C"�y���O^�}��Xb�!A�_5��Y���jF���' ���%�	[R\��kb��&��)F��zT���'x�d��m�<�z�F�.�(�1�	(	.��	$�[/[]�eX�CЉQ�6�(Y�Őu��̀w�� oBh�/V$�����+��h2#������k�y�tl�ʃ5JJ�0#��Y	Qƶ��a&3����֖����҃s?	�����O�$�Cw@4��Uk���X�xZ�4x� ��C�=i
xY�5K��"~n�%�i�$8 6�Ux����e�FC�	�k��m�$�٫@�`)C%o�/P�2���R%
�(|�h��Չ=���BIY�ŕ>N�z7K��61�4���2thn�Q�/W+/'��+�-�b�X��l�����"?@���еl�0\c���~'R1������hO�` $��"	�F���_I�+���)�Q$�I �`Y3E�B�ɬ.f�k$�#|��k5�C,H牾G���`��S$2�����`!
�
0�	a�f@����"Oz���.R�jP"Z�`����'}� ��-��i�#���B:�J�d���L���L��a���q:R9HC�I�l�g���Ꮝ�1c�����6W�P��v��1`(��ψ4��"?i�ʄ�N��5��@#��UI�X$(aG @6�W���~^!�DG7F�>�2�l
_ ��!dΙq1�ɉeVT�:�. r�S�O��<k�n(�
p��ͅ%��
�'AT�`riO2lЄ�r�g۵G6�8O>y��4B>�0�N�LpIЃ�j��}
uǑ�j������N�Hx�4���*Ђ%9��[�!��KJ�LA�B�!^��𑷧��|�>���T�XB�I�y����MWΜ�Ċ�#OQ.B�<uB�[R)�nX�9He*D,�V�S�kԿ$�!�䟼�D�qE�;�X�`1)Ԓax2
��h]��Ԛ|�f\�F�Jt��Er|ڴ�L�y�ǳa1�����&o~р�����ě���y�%��(3x���)Ol`��7񉏒{��Z�j@���/F4M�E"O(��OǇ�*e�����a��@ �� l�|t@���M�Lɲ���E"����Č�[Bj|���w����R�M�v��BmL�^NR	��m5ArY����F\xuٶf�Z؊L+T�m�8q�E�nlJ9���	.Y�*�C��5�X�c#jB�~�?��ź(_�[U��uDx�V�I VhAC�	j���AXv�L�#� ��<����J8U����<i�ƍH��<ė'�K��L�G�J�@�ϓ�L���E��w/��?E	�X�t����D;�2����;D��;dk�#f0�A�9a�Ҥ�����E�~Z&A�!V�C��M*�x��X�#h̨�|�	�j&ޥj��C�FmYA��m���Ğh �I����N$t9W��L���R��[�L�t��p�(Q�t��/C�U�a-�^0�!CC�1$�$PJ�� iq�m��IN�5!��1:�h�s�Tq���?Sd�
b.��p-Yc
�(eH��cUGW�"��D��S�F-K
�B�2	#�"�S��)I*S�$��'J�B��%�T��FСM��S ��f͈Q�Ok��}nxĐ�m͛j�4��P��4��]���L؟L1���78� ���+�D8�	��N��l�s�xRd�)'8��6G�R�t���#<G$��;iV>i@p�\��E{�E�64*��I�KŨE���PE����J�@�R��PKE��`Ċ]]�d!��E���Y4.ͦ�;��@��D�D� �$�=P�Ωh��W�H�H#�*�!?�Q��#���C�j���L�5p�0ʧB�fx
��F�`��ͺ��i>����F'�?6k�-i2���#l���D�B6)�3�R�z�b�!�`֮:���J��峵cN(�rݱ��� �8��$`D�N��%�AV��&-sVoN	��Y�ԩ##`!��I�m� \��^4�a�')^�#���'8��"�S�w@������h���&c�*�0�c'���|��FE�[?��9���?���au��`01�S5 �B�Ɵ�XM!�U��&�x��F�*vm����P ]��58�82o�b��S�7��X��JzL♃��$t������|����G�8ɘO����C��-RKXAP��Q�N�z�y�H�=pJ�:�$�A!
�t*�����6ʓ;�(��W���P�0US��w5$b��O���u��'i��K��O��db��J{�����������' ɉ 	�]�up��)�|�l�0�V��B�ߜ��� ��9B)�q�:1�9"���Y���`���u�Q?9q#/�;e���T��=Vp��0�'�O|0ao4� @�i&�(jDP�g�T?M�Nd��G�f�2���D��~�T��D�E�X~L�a���ƔU�&�G �T��ǭ� 4����"Oz�!g��ODl{�J1L��a2��qfP�����ײ<��J�V���g�'�H�z3
C�i�Ҥ8��r�La�1�z��D�_+\d��@�(N	;9}R��ۍ �J�*Ĭ[	q���P��p>qs�0>YȔ�)�"]�R�DR�'Kڌ"�K&�"A��.JӸ�OK0�B1�T1�J�A���Y�P�9�'��mH�kL$���ak
W���j�t��th�@ߩ��He��)7���~Jw��dUP@bQK�&FD@a�荱�yRG�f�X����1 Z��`7*�,$p�s��'H	#���u�l�rʟ�<x��M�H�T��7Т]X��q�N+�O�0I�e�Nif�ɇoE 1AJMP��p-���ƙ�^3�4�O@l`0�E1c�F�Z�!�V�lಕ���aRsV(թ�eiŜ?i�U C�H�&�"gj���1�&���ꖅb��yC"�3L_ �3�^XjQ8��'&�!�4�!;�䝥OQ>m( ��$u$H��ɥeR(ۇ�'O�-�s��VM,�OhȊ�d?�6�5#\7I���g'l�$9m�j5��/.��� _���A�o]p�sG,R�[m�I)>1�i��]�I��Ş7

H����	9ϒ�)��H��fqåE��!�����l9�O�i�`�ʏfoUx��jG��F�ݚ0r�����H�Q�̡'�� H�q��0'����F�Ӛ�8��f��dZ�3d!�X�S��59�b��W)=j��3ƢM�;�
Y�����v�ғfI:b-��?�V�0�"l�9��a�0A���
��&/�a1�y��q���[E�	9'ܠ
��
�S�x ���t�[a�qz��ې,�Ȇ<�+0<hUG�8A�U3��@��2�'t`�cd_6eg�!��Qo�{Ҁ���&�� ��@��R�9[@˗�l<���ŉ����0O�0A�&���A�������	Q��uxҋ�<!���&F7�	FY�50�	�x��.L%�=�&�N5s�RP@A�5�azRG;Q#&��P��w�hQJQ$��-���ƅ�0� ȉ_2�QoZ.��w�eD��">�@9;�x�Y��X���y{fgp̓��E#'ŲL&
��#l�� ۆ�qɟF6X�+���4��:f�*ɺ�B�$�����N Ha~��K=Y$p����M�4w<0�
��Q������W�<���(�'C����C�O����0!�-r�Z��,'À�i��3D�<B�+�]��Yd^'T	�"�N�&�|T��O��hON�W	�PʠX��'����k� j2�C�N�}�
ד)���Ӡ@~���2�IC�|A�Ԁ�n$�F�L`��|��˱�h\
���/A@���WdR>'`���!))}H�$�}G"�{*O���P�gh��ԏIX��u(Ā�?1���ם	:��R@	"���'1��� ��Z�D���n}�XE�'����ūĹL�@ń�	v`\J�Bۜ
e�t���þo���Dχ4�3����tb^��$�  ��T�V��LI>`��/D�t�1����C�7���s���݈������K4��q$�G�O~D���Ε���aI	i@j�;�'B(��j\���aˍ�f>��Yrd�/��՚�ꏋ��$)�g?i1a�m��:�M=y�fq��JN�<A��[=/i��*dm�;mʈxA�П���ƚ,E�8���,�A���[Ɯ��XXҎ� ˮ�C�G)|O��l9Bp��cA�C2�:�k0����� [{ �C�}[�T2��V�<^ )�91 `㟬G�.(��LMm�O1���%&���m�Fg�.d���'��%�Ҫ�5�M�F#E�SR̰[e��)�T5i�`\$��D5�g?���ZW>q�ƈV�@��ؘ�oYd�<��c��r�(�b"R n��`X���<!WM�*#(���,\O�1��
?#x����g�(�a���'�r���e�;w��K?n�A�fZ� �4;�B�y�K�.��ԋ��&5ʍ�ɟ��yB��=ZEje�˼�v�SO@�y«W����Dl��P-�c��y�A��R)� �{�dq��-�yB@�S[�P�&e��~=���f٫�yQ�&�����Z�;����P��yY,
l
 1F�;e0
�:��!�y�F��@RP��B� �Q#���y��[-F<�KA��V�\5�RfZ��y
� �E�٦mC�|B��47$Q�"Od�6�Ԕxu�>�"OL���̝1x�h��#HO�y+�"O�j���>�`�Qf�,C��Z�"OZ@��F��X"���;J�&s�"OVD��&X6�ڷ��܊���"O CX�3�R�lgvx�"O�����`<�E�Ǒo�ɠ5"Oza[DGGd�fA$@=F���"OF�x�"؈
U�X"�A�4E����"O�pZ�)\�~�ԩ��i��!�"O�	�F#�4N�Q�Ϡ�<��"O�H��[<��Re�P�Uq�Mp�"O^}˵-��Apd!5e� Yf, I�"O8�[�iΔA�(9����=lz��"Or�hĥ�9��� �Ň�oR.��g"O����W�[S�����n��0"O~=���
8�PȒ�3)�����"O$ˡ�±3���i^5D:V��d"Ohd)��Ζ�d ��(D<>NA�6"O80���ӤA�vi��#V9Te:V"O1��'��r1b0�Bb��V-
�7"O�Y��^66�y���	JM��"O�}�G#�=վ9��%��^Q"O��ʀ#�1s�0�������p�"O^��'#C��59f�K�A�DHa�"Od����X�XS�1�ꓰTy�0��"OZ�����]����2i�>	*�p�"O��!ҁ5�8	��;�&DɁ"O�5�u��$S>f�
D'K�+�B�P�"O�1�׈\9w��5ˇ�K�����"O�ܘ1E��7��sp��p x!"Oxt�T�^&kp,�ڧ��^��0�"O�p�G�Pu�A1F%�C6%jV"O9�#	�}�i�g��*�Y"O~E��B�1�,��S�\T ����"O�yC�KǸi5N�~�Y;f"O2���O4Fv�ɢV�MV�=2""Oڼ��D$Y_�0�J4�\��"O��{N؆Lf�E��!eߨ���"O�!y�' 4�B�lƿ4̐��`"O��B˖b�~PJ�˗�|=qQ"O࠰�M�rf� ��GVC��K�"OJ�'�Z40���-5o��"O��	v�ӡ|�|h8s�4NT�"OܨQ�o��A�^۲�ۄ98� ��"O��C�	>H�,�:�
.*<�8�A"ON�Y`��.�bE�QIN=�"O����X�B�İ����@�X���"O@�KB�'x�i���PƢZ"Ov��G��Wd�ͺIU�.��"OR�s4HE//.���ɗ�
8��3�"O�\8 � =H �ҧA�	�p"O�H�D�85j��EeN1l� �)r"O.ĒA�ЎH��%�'̈́�8`(�"O�T t��$&�F���_�M��((r"O�J6ɓ����a�#E;2�K"O���d.N	(�V��Q�F3k%��J"O���g#�faN-b/�%`�jV"ON�P�h�6B�:=;�n���2a"O�Ma )�1͘h8bP
g��rA"O��b')P#1�!Q.3\q^ܒ�"O��d��r"&�"��EnX�ـ<O�t1"��⸧��r��a�T(]b%[�g²$\�x�V"O� ��j����z���I��I _7�HH�^�0Zv�3$�xل�%
��I�W�Qr�.4� E �����
B�$2ұRA�*���"F$��	��J	�'/Z��X�> �D�$ �\���B�%�� �l���O@���bS�F�>�P�DЬKBmk�'kh�Eg˅z,]�I�5�tx�4B��Dِ�!H�6ӧ����g^��l��+��IhyФF�y2n�F��UI��н�|���	����
#d���G�=��<w� �L %�Uona4�DX���V(ъx����FY&�*�K����C��X3^c���>]����Y+h4Q�A�Qtx�Fz���+k��(2���6�b>�!�H �Lx;E���h��� 6D�,ےLј&`��W��-?\x�P3�wӖ="SA�3�$ ��'�/�~���i�L��@�֔OYX b��V�M��$s�'4��	��W����{�)X9A�N	a�O^u��^)J��!J�BH	��O*�a#Û2;S�I��	T�v^���q�'�l;�bK`|�%L�}�蜻�T%a��RF��X�d���=6:
<;g#�>C:dQ���F�aNΣ=1W� ���pq�Q�[V�O
 �1���C�����y�����'�XA �CEt���sb��Uٟ'�4�y4G�>+r5Ƞ[�"~BR̄�f_��H)	TM�$0�G�<��'Ñw6�U�!��k�%�V���I;-5��3�,��g�z |�W/*_��4i�#��2ȇ�Ɇ{�p����#�Ż`���s֠�.�
es� z��'��K����	PC0�6�h��d�[���MN���GF�T�7��/��5�����A\d���w��&?-B}���2����'y�}9`
�Dܔ�O�>y�u��.���r`�ɛsU��R b9D��q$�}�B�"/{�pd��G6��/y�zp��g6Oii�"���(�!a]%�ic0Oay��98tM��.G��]X�C�%vjʰ��'=v�y0A<
)�TY�mɀlv��)
�'W�l	'���)X�I�G-gZ�A�'j����
T���E%п+����(��L\t���[���O�$EJaS�D�?1P܄��I�~�1J�b�I�y��(	�) J�"�g�"��B�	%?D		稟�g�zL��*H	#L��~��A�*"'�8ic�<i��G$�ħ*�Ұ��,I�2� ������Y��=K��N��bQ�X��N�p<����d@�L��dn������'j�����FV?Y�.�q��R$kG�$����Wl���r�n�|��9ӢДR���G�{��u�g@�0*QIq��(|儤��+�&z��E|��$_z����A=z�XF���Ox�y��ߥ bԸq#X��x�C	W
]W�5�)�6L�<�o�V���E^J�����F!7�]�d P�IOz�� ���	�B�2����=:P�!h;m6P�Ӑ[��4�O2����I�V`�AAX8*����'�p��t��.Q�ꄂ�-�&y�L�ǎ��O�T�U��:��p��n�=��'9��L�'��<�yb�#�KCA 2��(����?G�Q��IW�A3X���aGf�ܑ&�Z�s� �Q#%I�v�TXvh�o�1)���E�ez���E�,3"�8:�"X,y�ax�g�`�j�qQFP�n���b�3>���3W�Z�n;\�P$�6�␲�H8v]�E��#�,���$�@��ֺr����':h<5���ޅ�1{���֓e>`(8e��Z��S�e�4�5%D�Q5�a��/ `�B�/ХaQ.'�t��2�e�0]Q ��*&��zJ<�2@/��K<6'���E�� �f��6��✛\z
�T!(�O.] b �b�v�����&���ub?��a�G.k���SB���c)@���ܽ28�}�S�R;�L������$'Q���c\%?�8�!iD	Y
X˧yWx��[>F���@�94s�%��xl8@�P�2x<b�˵�,-=���;����,bda���>��i�ff�B�rA�.!��t��"O�x�aǝ$Z)�&M�x�Fȉ`�>A��6>�ҥ�C�2O� R�T�
��O�:8l�4�'#�ႄI�W�����ʡ!�����j�0�|L)ehPx<9C˗!��|�rǐ~����R�'�t"0�K�-q��|Z�n͋u��sr�R�<U���Z�<� HeC'%(`��@�C��B
�@��OB	�択Y�rZH��}j0�ԔV��i'Ėf����P�<	%C!��T�3�Bq���Q��g�	�#�Б��s8�<���z�����G 4���0U	0�O5⣈ԃLfı��q!��H�B�ZC(5��'�<�r�.�&G�P��5!YRS�U�'��hFDܹ,��!�Q��7}G4�X�'����4].=�!�W� ��'��I�G*��N�d1į�v^t��'�THkd�.�VEYe���^�t�	�'!H����B[�6���o �XL[�'䢬�ǌϖEmн;��ҁj�I�J��kW��qO������&9�Q��W���I��"OU����%rP܁�Y�#:��M1��ق&0�;���d��.@�C����i�A��R+ü-G5���
hf\Ś�g[�d���r*�M�����!jOJ���M�3��$�5Eݳp"(�?9��_5$�PT3��7�	E���s���o�ȩ�&bրG���T��I�@�ғu���aTe>�q�.��?IG��@Y��A?}��I.���(g.ԗwr0 �Nax�E�q��t���|�F�7{����r��.o&��Pg��h@�'�FP��@�Z�ϸ'IԐ�cܿ(F+� �x����/O4�0!LX�sE��K�b>�c����*��4s�+U�2�b����]�fT��˒͍�u�a�	ُdz�B�N]Jm��c�c���'��$r�/F���̏�Q�ā���b�$�s
R]u��j$N�9�IRD����\8p J�S���Z�����Z��5
��Z�pPy�%I�Mp���\#A8��3��)ܣ���Z?,3F�C�iE�w��s��Lđ�d�a�I$���dh �D�6M̐�E�9Q9j�a� �3 ��y�D@��~B�"L�`����"��E�N�@а���>igB�	,sq�t����i
�A�<�wBƤm�)Ŧ	/ބ��fש$1�lb4!�%�\�Ѣ�8�x"�A61u��W/�t:��Q�V�vb�\Õc �4c�;����G�<A�߳/Y�|���Q-��� @�h���Q*xÚ��cȅ&��ŋр6(ޑ��i�x�(O�yQyG���D;l��8c��R1q��(�0"�dSQ���F데A�<	;gi,�DQ�4/R��ƫ�`�
�dB>M� %03b�k�a~�O�����@�-hԁ�Ɛ�~��3�\ӮO��pp�L��6y��������Y�sd D���d� �k}��j��Hq��i�TC=\O����2�)�<�S鑴F�f8�+k�e�0f�|����g/�$D�����F꤮,%�.31O�S�w������!�#>��ƀUƘ{�	އ`���V'\j�@Ẻ�v��'k�p5,I�u����!(��|��A�C^�B�]�E�Ѿ��[��'6����w�Ν�gl	�4r"}��'���[�{��D���+
����%�{�f��bH�	]���D�/����u!M��ܥJ(ߔ|�F��R)իi�\r�*D���f���.vT2PE�'�<��?�$�%Y�����`Y��i��N����6��5�Ǯ�v�!��v����	ԸV�Fe3Am���z0רO�T�Cu^�dF��'��p!���r��Avd�����'D�R) "s�Mi$�3�P���-�PY�ޗcF�T�鉢V���SfN9]*�d9HL� Z���p��dx�  U��a��NC� D8���ɠr;���'D��rt+MB���d)Y,��<+��0���e��0�E�ט"�,E�.�+Y���V΅�I���Z`�Ą�y�a�U�t���$ѺJ�PiC'���5,8a�+L��,OԢ}�6�!���V]	j���&�2?D
��ȓl r�*���.?�l���,;8���b���7���d1:g�ܰ2iU#'�0A	V� E��|e؅B�
U�i�ZX!'_�p�� ��c���U)�'XAՊ>�г�P�EĲ�' 
H��a4S� -��l�38��PC�'x��t�-�h�6剂n'Ьq	�'|Yc���^nT@��8Y�x���'e���6�M�
��m���N�!k	��� "��D�|"ف�-\�ld,�q"O���&���R���g����X�%"O���4��2c��0!��H��@G"OP����=���R嬨�S"O��+�!&;LȀ�Ə�)~���F"O�I�I��	,�
!��De�E��"OX`��cG 6���9㉰^l��z"O\qI]<B��j���<Q��s"OT�W��'I��� DyF�T5"O��	���5!��X$-5K k"O"�ї�Ni�Ш"�m�K8^���"O֍ 7@��Z�(�%l$R:F"O���'��= /�4�f�ؐ=��|�D"O6�`�Z<^�%pc�8H6�� "O,�9֥�	h�
R
x ����"O���E d$��p֊�-
�c�"OƴR7��:����C�M�

ݓ�"O��f�� 8�8!¨Gþ8Kd"O�`81�%ui�AIRGݻ6ʊ��"O�P��` �L�NM�'� (F^m�a"O�L�||�iuǚ1t=����"O�j��	/`�Z�f�9G� �g"O�	�f, N��$��E[�i1|XY"O��b�-M����@+�cw"O�1!��i��%�1L�Y����"Oh���C�56��1���^��yH�"Ol���v,�����9���"Oޕ�U��5�p�jM�X�q�"O=����=|�D��0��v���7O��'���	�����gM�r�a��,�B<yS��;B*��UL�|��B�Is� MR$(B�V���@e�L!H>dB�I'S�
���Qa!  ᦯�0~@B��9y�␂@�D�X���R񨉏3p�B�IR��1�o�,$�����|��B��	z��tX��^)5���f"Y�-�|B�	�$�h���6��M)cjL�`�C��-*�`h�"'YR�Ijw
��tC�I�3��A�E�cϤI�"J��s\TC�~<$"�K7%|���( 0J�@C�	$=�bQHw�N#>�\q���?hC�I��RSH��5*�;a� �nB�I&z�r��%k0x�b��u�@�>�I����|
�(���#�=&V��T�������ԃ�اȟ6p� C�%ZT#5ž?���2@NC7]�O���S�E��kc'�+N�f���	?B5\�Od��I�B4^��i[)dg���6�ٓ[���h�Ə�剄fNlA�#�]Z�)ʧQdPlr�C��AA�!+儃-H�\ϓw=�l$Zr�S�Osl�°�W=vy<�#f�C�U�F�6�Ƭj~�k�}��)�T#������9��|�� ��U�O�}�G��Ӳ�]��2�)�%��|�ȓA��s���n�h�%�#{1~Q�ȓ|���a�յP���#D�Ūs�r��'�ў"|�q�M.g�9nR>3o�8�a�R�<aU"��P���	�p��Y1S�O�<�v)�:�*%[�G���"��!`�<��o��Y�<t�� �ھ���B[�<)'�Y��R���ܔ2c�0x���_�<��.�v�%PF��y�\�Pȅe�<�CJ_,@e��AD�*,�#K^�<�g䋄g �AäʽQ*x|��P�<!Q`1 ���c
T8>�n8���ON�<���/�j�ip̺A�0��F�<��GV��(���^�thp�4�z�<�vB�O ��R�ó mڰ���t�<� V�@,��
����u~"O$a��0��!ˑo
B!Q!"OP��f�ҙ/(@{׊�v��i��"O^drG���uj���KO,���"O�s���DM�s��#��A;�"O�̙*ْO �y�(J�
���"O:Xi�Ͼj����fN�!�`H3"O$�E�K�h�(�YO:>�d�&"O����K�8B��H��J��&ĳ&"O��p.��Z((vM*o�F<H"O�(����=34X8Tm�� �q"O� �4o�05��k��� �\	��"O�5bn:`��YX��A���P�"Oh)��h��芃@��u����"O�)���N[�P9a)�!���Ӕ"O��Y�']<��m�"*E�V�r���"O���r(U�?r؁	@hW (�h�Qg"O��A`��)e��|����*��Hȇ"O�=Ka�ުB����@25�,h�e"O41�F�T�GV�y�C�
`8�"O����R.;��;�#�$��"O�U�s*T�3�H�z�.#���"O�� ���w4��F�چ<"@h��"O��I��&E*�)��?z��"Op��RH�s�(�R��.J���W"OHy����S=4(��M0A���b"O̡��)��*:����^'$�lZ'"Oh�"$�x�A� ��%.�|!�"O��I��K.�\@p�%�!dE!#"O cV��C�P4*��\?^�.4�2"O�mj�oXql$���-�B�pɊ�"Oj5��ä]=���M����*O6�j`�a͞�BLW�a�U�	�'4$XAcɖ�N��h"�c��\�8!
�'q�s�ᇅ+:V�0��qQwD4D��`���?KPػ#֋U3�%��M1D�,z�ɴ�&�c��� t�X�Ҥ9D��K󤅫:v$ek�-֊e��$D��R�6e\!��\gjdչ �7D���&/��@�q�m�-P�Bѳ4� D�t�0J��@�F=1G�I���@7!3D��i���HŨ���ē���g�<D���'K�}�j��r�&�Q� D�P�W���^��bw]N��%:D�h�3�ޞj~�x�E�ί^B6@�S#4D�|qG�L=�!��ΔU�(�Fc3D��U�۳=��S"h�$�(͹�L0D�,4aդ{z a!��<z�(�#w�3D��elS�%U���Č���$Ea�=D�i�쇅5b~,�cbR|��s�0D��� ���~
6 ���ۺ��@�k#D�L!��ٙ0´1Q� ]b����%�&D��!�D9�vԋȚ�=1���b#D�� ��i�*e�0��u�^x���6D�4�T���p�͢I*E"�LL<�yR'�jIx�2��^5s���1K�"�yb�_ L�pn�^�ԓV&[-�y�R�<3�1F��)���+����y��47%3���w$��Ƃ�	�yB"+, �'.�7������y�^�h� u�V
!6�J�%��>�y�O
dPz�շ3-�|�I���y����ɺ�IǢa$�K�����y��H���c���5 ���P��y
� ����D�''dT��SI��$�����"O�1
Ǡ֌o}����R�"O�}���+O���Pc��dc�"O���jW L�T�L�Wg�2"O�̡�J�2{Z�
�ƀ?Q��Ԋ"O�`��R�F�$�B�j�LL(6"O�$����*TB�37`r"O���RCD�.����l�t2���p"O�=�&�ιc����2 H/*]��"O)r�o�`�LM�&��
T�Z��5"O�A U$m��	5Ƅ�j�b�"OvK��� �qjNX- �$�*�"O>*�Þ�G6]e'\8 �x�T"On8��I+�x�G�Qc�N9�S"O��jC�: #���%B�|����"O*(Hd�B071ȁq��S�g��1"O�M"RƗp��@�X;^窬��"Oض�#y��aP�88ɦ�r�"O��'î��	�l��"��� �"O��ar	*m��ɂL�;0�g"O��"5��+>䐉�+))6�!�"O�A���R��J�D�G�p&����"O����b�����
�A,i�0"O����)�Hy�聦<g���"O�ʴ+L�V� ��ƗYv��
�"O4��щ��B����.l_:��"O���0.�;W�X��F�1�h��"O�9y�-��|r����0��q"O�{�J��L.�|���q$��7"O�<CW��/Og h�0�t�����"O"��� 0	���EeQ�!��t��"O��'�+�	B�팣f�ȑ"O�3�e� ��%�$�U���h�"O�� V�R4A�<9��/ �*�~ �V"O�,zᮕ�*f��狔A����S"O����ɣ�đuJ¸Z��8��"O,�H�9nT�����hU"O��8#���IB������n�@H3"OH����^�d��T(�$��Mq6"O6dkb��#�Z�Y�eB�Xfz�"O�`���>�v��c	+5Ty�"OR${!�Y7Ӹ�@
; �`M�U"ON�yA+@�zO@�aU4e��1�"O$Ƀ�	\�vR��p〙�c�-	�"O<�*���;W��t��-��uO�Q"O���V�+3]��Ȧ"�-<�,�"O����Ç2z�4��T#Q��e��"Oj�q�T�H���4���3V"OT�q'Ђ[���(@�c��	 �"O����R\��G��+-���"Ovy�a�ܘQ%4͋��X�te��"O�0�+< �V����'?{��j�"O؄�$o��9a�P'%�#v��x�6"O�9�H�u�2A�2C �8cW"O��a	Q<�H��"�_�F�Y"O �y3m[�Eʡk��Q��X�"O�urb���k#��X��<iC"Oz) �b�S ��%�F�y�Q1�"O*���B�sb�i6���,(�C�"O�T`v`�!F��I� Z5aYn���"O�eP0��Z`Y�X�6J��v"O`Y��BLFYa⨂-��F"O� ڠ��&�pA1�<��}"�"Ol!7$=�ʐ�%����<j�"O� "͛�$�*��5y��+�z�;�"Oȅ:#����)��Ne�Z,�Q"O�4B�!dx�	@�6";��b"O�Ѓ$�٠p���b��6(�qd"O.ĂU�%Cfx� b�>O��j�"O�YȔ
.]T�h˂��.h���X6"O�K��U�6DB�@��b�Fm�c"O��"���$���&̷m��=�"O�}�%��U���ƥ�&Tj�|9a"O�8� �{���R�Z�Y���!�"Or����Z�0m�S�ζB�ڴ"O��PS��^\��A��J"��H7"O�(&�
�8�N	:ei�oj��%"O�\���X�W���!&BCb��'"O�0�&
��F0�������9q"O�bsm�}h
�9�v�Ę�"O���#�z��T f�ۣX�0��"O�!s��Ԟ4w�zdD
:R�nH�b"Ot@{r�C+	T���F��@��4#"O.<�K'sdTA!��`e|�`"O�2L& ���A�#�d�$"Of�
֏]�r�I�"��H�"O�(pbh��G�
��whP)�T��D"O�����of�	�GўF̜�ۗ"O�%�"�B%�E)�e�6>�q�"OZlRC�O:^�Q#N��2a�"O+B��g�bT�#�q8��"O�%�v\�7E֕ku�!D<Zt�C"O�a ��[��]a6�M,iת��F"O� y�'Лl��,�3�U"O�l
�4=8<̙F1>�Ha"O������'=�T�Y��@�/%�i("O�Q�Iv���Y&�	�,>�-ۇ"O��*���=��|�2@�6D9�4�"O%i��B�3�����_9�	J�"O��{1lM���RDo���c"OެJ&��F�sE� (e��"O��XF
�����1���"OT����N�W�@�w�Ԧ&ќU�7"O��ʔ�-uDih��K��9�'"O %�W�ހ>*MP��D�	J��"O��؄# >'"d��67��X�"O|I�"@"r��� ��FD��1"O�|h�L�~-��' >�S�"O^�3�E�#Vt�=���� )t9�"O�1�H�
�r���W�>ya��"OPHRǠI� Y�Ɔ
`(�y"OT�P�ճ!"�ɧf�%�]!�"O����Q��rs�G�n�Nm�#"O� Q!&-'�P@�iנq�<[P"O�<�0���D�Ɣ�B�X��Ũ�"O���p#�l�s�N�[��zI��N�2��e	��Hz�l
J7M���ȓ=,�=�&��<T����`#�1s*p��ȓAl�̊��X=X�a��
��͆ȓq�@���Ɔx":�kA����<��HH���B�R�3 18v�K�z����	���T�@7-�11-K:).� �ȓ>���� @�?