MPQ    �y
    h�  h                                                                                 gKI='
���\��{8퐸IX(�H?7�-��sku%E�^|�Ȁ���"3Hg_���աN���~�;�b�b�0��'TH/����t��4�\����}�K���%�ڝ{U?��pQ��cs�	̂��2@{���,�<f6+�b��[0�ݲ�����m�ƱG�5�s7�/�������pX�r ^z%+�����ж��N*���Z��H
�o(wl�-F�"Ą�&���TQ^ϛ���~�9<�@:o��R����AK��m�cGP���ap�L2H�C�J@k��0�ڙm�-��;�&vd���L{���^�/O�G�5M\r�Ĵb�6sii�vn�r4C��?�(*�Q�lE6%_��;C&��q��H<�� jX"h��S�*q��q� ����1����X;��ˍ��'d}���4HN��K�'A��]���4��]��RDs�&7���G�b�T# �����E���x�~�hIq%vXa��%�n��0��9�z�L����2��& 8d�~v�����5���0q��� �s�y�G1�E/�R:w���dЛ ��d����!� 40�I���*�Fd��-�{o���{|����X�<-�Y���	�M_)l���,���U�V=M��n��fr����atƨ@ZϪN4]����Y���}��߹K80�h�Sl���4~P�ڼ�T��M��R�$ɌG��B\�tf�r�E(�AYk�,-P���*��t}���l���`��W*�5/~��2g+�SV}^i̱�9�%�2�U+q�ㇳfMV�Eߔ�Q���ncx���Y�d�Lâ�JƦb4ٺ�z����#Zs����;{2�M�X���Z��'z���Ὸ�%�6�O�0�z�PP~Y/_[�.�@,l��=�?8F�h�y"�����$(��"Ƣ�:/Uj|Ц.oǉ�K������X�p�0_�)2���̤���aĐ�5i�r�/Qh�"�ے�_7�G9G D�ٲ� rH�]�Qy �m�R����;���;2e�T.�vG�"#�nr�.$0Y�3$��
_aϽ'��Y<~�h�N����B~6��@��$������"���a�)tɔ����)�\E�V��	?������<�,�t���A3�JH�A�����O5���X��;M1���@�J���/VEoZ�"�ԁ7��������dL�2Νt�?�<\ˬ����(#�O��w��)`tӅ��"������Ÿ��6}(m�,	����̖$l�.\J8�A�c~��Ja��i���4�l$s�<���G٭������Tł���j�c�wV]�Z.ݫ�z�Ϳ��&e���cK���1Eh7�r���n��{�bȕ(6;6DЗ��f4���Z���S�C~�g/�$b����\��Z=l~r�M����ɧ�ԃ%�MҜ�����h��j.���Sy�c�ȡh�Ft(5ޡ���P sl�o��>�L|�1s�<�V�����w�1bl4-��2m�J�)�{�Ԥ=[�b�s��h���@tߐB�y&�e�ʑA	�::(-���+�x�QO뷎G҈�⫭T���-��.��oa*�C}�[���E
�[�"�)d	�W}F3�C�Rɚ@<�}i�kF�a���ii'L�x������m�7`P����C��ƍ�Ħ+,�**�&��`9��7U�M%�n�����%�<�V#/n3cQ��Z9W����e���ݛt�� �ATxP��gΧ{�fFJ�(�>:�Y!W��o2ƯmeBϜ\'q���P$~-o�9�Y�,��h��=o��_P��{S2(����M1�j`��}�}R��T(5�Цs�v>��� �Z	s��	ϡ9���A܏X�40�������}���C��|iߪ�����^�'��@]
S�șb��w��%��U���� �| ~Gƹ��,��CK����b]v����^PA��������j�l�aqj�>'�sIĐ�z������?�s��x�(�z��-l�����خD�V#���2���J�&#����ܢN�z�Cz��Y�fPS�D�"���rDR��B4��Za�F����kPܚ�$o�xU��P�CmR�d��P�h�w�M.͑Ƒ���e8��W�!U&�a�d�B4�z��>��Nq�f���i������2�_"t�gz��C�_f�3eP?��(��~*M���ِ�y2�-�H���2����`��E�y��/�����<P1�������I��7e � �����
/��L�-�?����jJk�(1�� ����U����QP�Q`!�t��O�vg�8e��	��l���I�:�l����L-!�ث=��Ќ�ʃ���|$���X��#��Bic +�O�/����b�g�u)v�%8ʶ⻕Nޑ�by󃋮7��$����
��D5W�o���O�|l&���آ?��y�mH�_���d����,�*�l�����ge:�8��C륙��X&]E�軜�[ =?�H�&��Đ�N2���'��&*���|���z�^n���t�Kiǭ�A��4l��װ61[��������=3��5�����f�����X��!<3�M���(6^YA��r��u�v/�W�c'���
T��LR�oj*F��1���N�{?�=��ՈH.�`�Pb�������)�ԣA>���rd3���bx"g��h6��bt�fA�疨N�5������h,�Xe*��B�F��yw��S��4B�`b4|8S=:tZ��'q�]G���;"b�	 �p����U?��cLR���@.�&��Y���uc�`� [S�HX#�\:�O��y+�]�z{ �8�����l����9a��pp�Yq�EA&���(Hs亻�{�Xs�!�$��|�ӣ���1�mkM5K�ܥ�������sQ4��'a���JR�6������1�k�ܝ��D9��H�x�q�^OG� ��Q���b�7��t6����&T
7���	�6�%4ݴ��h��A
ʥЌ���!���~�v*!,��l9��b��s^Gu�5_ ����4�6�")�~.�kE�����}��[�,{�1��c�����������y�b<�X���&�k�굵�b�c�k�������=���oM��B����(��v�x��� �q�C���wAn2y��K��p�.��� ��@�d�dZb"�0z��<|����NǙ�湷�[�8psG�r���%���2�U�Q��N%d��sBi��<��Gw�Z:F��j��L�t�^�/k��1��̔c<)7�:�ǫR�_�Z����Y&cB��U��p�V�H��FJ�ϐ�����p���t&q���:�܀L)���[gO_�I�m\������6ntaie�Ƒ�^Ӕ��*��l���_u4*;>�g�̶IH�;
 ��"�P��.vgq&_M��L��ď1�	�X���˨�"'߮p���k4��g���AC$�]��(��'ꑰ�t\D�VY7^5YBwbK�< Q�X�����;�Y��I�֜X���  =n�]0��|�����f2�OZa�-d'�#�Ͳr�5�������q��N9P��O���M��:��V����ж�T�Jl_���!!:�X0Ec\��wrF���b��{�Zw���Y���x�F5<�7z���:�vk�nќ,T�Y���1�C�!|.�G	��aU+a
{�f�[�`��6�]����L���������E�#tS��ɯ�g�~+bM�4S�q(�M-���������t��rI�a����g6�H�}�����Ө��׀g���+5
w�m{e����^d�����7���+��*�.{rV�馔*��!�n=��.鵽2jL�~�JA�b(ꤵը�Q��s�b��Ӏ^�X�x�Z"<�U� ��O6���΋M\���_�*_֡b.i�l(>���\$F�)y}*3�I��$COh"A��:
��|�ob<tK���=n5X��l0zlC2z�*姟T���ߐ���d{���A�h��ۭ��7�s��D.;r�������Q�;am{���`�H����Ti#�G{�.#��r�t�0��?ڥ
��ڽ�	Yw�2h)�v����~��@{sL���>���Ƙ<]�td^���B)3�rE�~��$^��X����~,���D��<�J�kp���Z3�AG�e8�15h�@�w&��V�a�eA���v���w����9�Q<�L5 �ΘҲ�.��$����p��*�G=%���ՙӀ��"b�&�?⍸�������m�*9	��U#��`o.����V �c4����}�D<�opo$ؗ����@r�@d��&��E��EQNܲ%���䫫̦�(����Y����y�)�1EC9��LP��>n�o�����P� ;Q�ꗕH9fdG�������~��g��-͒��\�oTZ�lrh�(�0���.
_� s7���
����h�5<j��<�S����%�<��Fo�k��"�Rq���?omY+>�{|�7w�׉�V�p#���f��/4H��2�:J�����oݗ[|���Ά�h= @��;B1K3�@�q�|%���݉#DO�+"rx\0�҇GM���W�T��}�ȳw.���a���}N���G
 ��"ƀdDEW���3��؂��@�v���1�K�����ib��xv����8(�b�iPn&��5�i�S�,7s���3��W�9VU�;�䉻2�_�� >�<کj/	�L�)Z�$I�b����X/Z�^#uAP�P΢Tf�B(�B��t�z�$N�ƊT}8a\¡��ǅ��Gv-*`6�6n级�^�COux�b[����2�KO��g�ȅ�I����}�U F8(�I.�n/�>�v� ���s�����u�}G���h4˕����+�Ia������jޒ�s5��L��a���g�;�Y
z"y�T'��!E���bU����C�� �$J~Ba7�^����K6�(�7vxo�� 
ܧώO>��:��%�{l�I�jO*k���
��5޷+�y�� ��xA��.Kx���zP�-G���I���I-�V���~���#�f$^N{+}�~F���oofKי�l���#tDm��B��Z<kɜ�~p��WUkKn��@�x��P��UR|����W膰�H.*����q�?�#��vW4�A&�Wd�/ü�c>��MqV��A|
:?`�2��0t?��g��C�R����nP�T�(�M�*ȶ�ݴ��ym�-��(�����Sh�`��Ӕ��/Lj����<R^2�>���uBI8fe�]$�"���

Z_LG�?�0"{f_j�>1(�� �t�d��w�Q��`�K���n�v¤8�薫Il�aֳ�x�ilo���6�!��=}`���x���AY�|ۻ$���ڤ�A7B�m ���Jh��_W�B�)�=8����;WN9y���p�ߓ�K��å�E��D���j͊����'�Щ�~���������	�!��zn��"��%��<G�7y�e���������&�EX�v��[;���꓆L���wI�ʲ��ӅсU��(�|�L�z�4�z� Ԇ��H�i�~���$��R}��
b�=�����vh�f�"��>�@����3ؑd����^4���Y�9�1O�v*�L�`�ŒwT��?R���j��lTm����{:k��Pۓ��`k�b�y���|�R@�oSy>m-��f�B�;}}�g;PU6o`�t��̂�wN���GI��T�n,�H&*.
yB��ԄZ��w��)S�QT����`��8n�:�NF�5剘��p,�f��d� p����)�?����L�^�ۉ�&
q�Y6�(u%3��|γ�3��\P�OCL�+��tz���8?��A�&�Ű�a��,py���@����tH.t���KӁ�����$3Z|<p���#1-��M�e���,��up���؋4N��'��i���R%��ia2�/���O���9<�
H�O�lŹ^��, �@����*��O�����T����	=1	,�-%������%�,ʀ6T������y�*|�F蚳�������?ju�F��?g �;4��[E6Y)+�9 
k`Ǌ?���9�Ԗ,���U�2���Z_��/�݂��38��a��ׅ?.�]S���|��n���ǚ��5M�����3��üv� �v����C-f���N8n6'�T���gƆ)�A��Օ>�d�b��z�ue�wߍ�V��I���A��+�p���r�E%�0��mm(��#N M	��Jm�eP�fowbISFx~���Z�v�^����Xen��32<D�]:e�R��w��)�/e�c=.����jp`�TH�J6Tu�����ト�	~&l�Ⱦ�?��_�ާ0O��<몺\賙���
6i��iw�[����y

5�*|�l�`*_�K;9Ʋ�'��H�� �6h"^���	��qa]�V���:�d��X�$g��� 'Z_0�eS!4�kՌ)=���A�Y�]��'�����O��D� 7���=E�b��� V�4q#��C�4�HI�WX��1��n;�L0c�c��Q��᪱������d�%	�ȉ���m5�h������j�)���D�¸�HC�:-���m���-��œ��gx!u�q0�����F��=[{���qA��sx��2�<c�2�������̜G�C��BG��i�\�"��H�\XB�lr�ׯI�v��?t]�(��
`�1j~��[�3���>�S�#د	��~%0�oq��ƖH��B���×t�Cur�b����̢_
��\+�x��R�6�Iꖀ#���M��5�
Ѩ�S����^_
��	��Y�+�������V��>�e���n7V��"�ږ-L�z�J���b�	�����&Os�'+��#u��M�X�_GZ��0�"�Nlv���(6ۇ����]�z%����_Q�_.D�;lc�:�u��F��Zy�䏕��$^�"�C:�K|F]'o��K�ᚘS�XEr|0�E2�Ra傺`��-o�S�9_l��Q�hT:N�ȍ�7j3ﲅDi�Ŝ6��ĵ%Q/w�m6���ʏ���4��&	T���G�r#�r�rGے0��wZC�
UZ2�ݭRY���h�+v��O�~즩@60X��?3�_�ޡ_�w��t�G����)�q�EpƮ�?�l������d,
��7���7�J�R�a^3�&��⼴��@U�1p �@=7��~ʊV�s �f�
��x0��\H����L�J�ΓPS�k��׬�̝����g=x�c�_k��{��"�R ��U���nY�,� m�H�	6����*�t
.Q��wc7
0�@t(�̪T&$�C+��d�c�����e�A��*�� ����ϐ�ҫ�P!��r0��nȐ؛��E +�G��F04n��C1���H�;lR���.f�-�Ж���ʨ~��;�����M��\��Z3�rC��k�ק�!��~��RJr�F@Eh��'j$���s��	��M�Fj�~�W�������go�^>�Z|�]��rwV�>�YKե��u4c2c�bJn���N�
6
[wH�)r0h�b�@�B�<l��ȑ�a۠p�,{J��8�x����HG��S�#�T4B�c�.�ڻa�5}	� ��
�Js"��d�oWS�73۽ ��@�nW��<�ͦ�ei��x�\���~��E�P)�u�:������z ,r� �\�V���9oUsI+䤀y��@3�۵�</�ȞG oZ�4t�?��y���+�9F}A�0P�J�ΝM;f�Z�(CfD��7���Ld�e�����\]R,��I0�-�׼Q���"*�����w�v��y�2޹��=�Ƞ"F�s"�}�y��׃(k��i��>C e��s�Y�ϗ��X����4f�����%w_�R����r��i�E�X?x�]3U�6��
�0�����Su�u�Uw!��~s8 $�+~=3���؎[jKQ֊����vS?Z�[�+w����u�K��ବl�Q'j�5���H<�?�ƕ���q��ӱr��Rx���z�rW-"�Ʉ�l��5�V�������#�Db���NV�ƌ�20��pfF��2��j�9D�kUB*��Z�W��uΏ76rkF ���1�x�IPߋ�R����,���꙰�E�.����G�݈���2=[W��&a��d=f��:h>�<�q������U�r�-O2z9otz�g���C�e���)P�U(�1*C��ݏ�2y����~����垮�`<g�ӯW�/�p��s��<�����w���Ip e�1��)m���
�נL@�5?1��v�j 2d(�t 1,2^�R(�Q�U.`W��ܭ*vú8�Ҍ�4,���x֎�x�l
3�@g!7K$=8դ��$�y�>�WZS$Q8�{��B� ����e_����%���)��88	��۴N����nZ��R}�������ZDC��e8�N6�1���v¢�����X5��Z�Js�Ű�F�آ�I������4�e��Pub!!�����&f��1Ԣ[Vcҷ>���!��	g������L�ܠ���`|��az��&�Uk=���d���ɣyB��t����c������=�G��Ode���f�_��{����S3����v�^�1��\���H�v%����T�Mv�T�H�R�j�)���i��O`{5caʫ�r���V`4�kbz�Y��m��#�
#i>�/�(�7��Y����g�6J8�t*���N�v������,�X�*�DBs,��f�w-B�S��"��]`��8���:j�>�c����=��B��&�po��Dw?�LN���L�R%�v
&`�Y�i%uپ�Ϣ�I�D\�O�2�+ű�z1�8�����bf�ŋ;a!��p�[�;+a�^��H�#X���1N^�מ$n%"|�,���s@1��#M����۾���ES�]�4��;'�����R�^$'��Je�a����;9w#�H%���g�:^r� k^���4����*���T@�0���	���%��j��D����[�[���x�Wnl�t\�*���U����G�iA�u�w�Ջ| >󞛢�6�O����k{9��������qe,�N��g��bj�f׭��M�X�����L@� ��X0�6D>��v��,�ٚy��M�O�:�'�^� vר�ktІvqCHPu�m|n�ˬ��*�Ԇ$x빜�/�P\d2��b�oz�����bS�����D#$ڜ������p��>r�H�%�c���nЇy3NV,�)s� ���w�WxFS\h�U��ܪ6�^������֭B�<_C(:�Z�R�@��ͻ�ʐ
c8�S�}�pʋH.g?J�����:�3t����&gB]���?�²���bOU��Ɖ�\#nr�3��6d��iғR�<1��a�?}*W�_l�%�_��;4ƙ����Hm�3 �x�"�;���qq�ߠ��ۡ��g���Xl�>����'�/��@3'4�F����$�A���]>��������*�D$7�pP8�Ubv� ��g�Ot������I"��X2�^�8�n��"0���?��\\]����״5d]�&�Àu(��5H
F�\��g��1mZ�����C/:����(3�����@�-�BL�!��~0{�B�zq+Fu�����{��@���J�NZ��O_<����lq�^tZ��bhK�O B������J�}Hu�W{�В}q���۪�g�]}`h�E�k�Æ�I�\�����&S��ί�.�~�����m��]�C�ɝp\�s��t���r?!��ҢW�ݨſ~�O�s�@ꭷ9�Y��>�����5��E����$��^ZY��Jޛ�cS�+�Ȑ�$�V|����l�WZ�nQO��{���L�]J7%�b�%�+�����}s�0�L��~]uX�f[Z�AU���︅�6�7~�A��5����_��.�l��L%F�yHy3�,��Ȼ$y�"7��:��3|��!o�4K�W���X�X #�0��.2p��]�܁7�r��S�Z}D�@�hvX��@<7|��ʘD�]���k���zQ�ҡm�F���-!�>��÷T�[NG���#��r�a�0�A�u�
�ֽ��kY�C�h_�����~GXc@�H� �4W��|F\��nt�Q���0%)�M�E+.��Z���N3�����,E|��s�2��JYZ.Q��A�'�7B����1���@��y�RVV���o�%�'���70����Lk��Ύ��Pɢm���:�f3"������{�� ��vch"�Y���z6��hm��A	qziY�}���.m1��=�cR ��-�������X�$D����cJپ�k���ބ\����.��X��($x�+�Q����{G�W����g�vE�^�>a��ᑡn�y]�
G���;�	���]�f����M�$�?~~'��5 �J�\��Z��Kr�����,�dY���?ҭ���h�/�j�ֺt��E8�r�%Fe�m޲P]����txoc0~>�E)|9�����V��T��+ĥb�@4~z>2�u�JI���,�K���[r�!��};h��4@�i
B'N���Б�ʠ�ҁ��n�x��=���GC>sqTo���0�.���a;�@}ġJ�
�"|�d�	�W�Id3֪�c_@m����U��́0�i�cyx���Ԉq���P�K��Uє+&�U�,�c:��2��=a9��]U.w�e��U���M2<P��/?ÀBN�ZJ/��𶓽�N����A�ΝPU�<Θf\fW�#(�������k�@���j�\�"�޽-�a�F-���l�|������`�+L����(t29H����0Ȼ�����Z}������(w�d�>��$  �7s���3�3��@W4����d��	nm&�!ْ�腪D`}�����ڻ1�'
0!���t�ȥM��
|URf��S ���~8�	�7��I�cKl���Nv./����-ʎ{����ݛ�Al�y^jEa������A�aSi����.B̠�3�x��zF�8-�+ɿ���^V�s�Cv)�{��#�B��cN1����>h�*w�fAs�U��%g�D�TB��IZ򂶜�� ��4�kA�ĺ5CHx�U�P�__R�
��s;����H��.�C'ƢJ��\�M��W*��&<�xdZj�K>}� q=
��IpAN�2U��t�LgK�0C՘E�D��Pp�(X7*���j�y�8*�^V�̫�	�_`�������/B���N�6<�ڐ�t����1I��CeQ%��Dء�|�f
�urL{�:?�kqn�j[E7(b�� L��w��-q�Q�*`�g���vx-8A�F�Om�b:��i�H>(�l����j�!��0=�i>�!�����2��$I˳U=�ABzvG \�؀v��U��Et)'(�8�5^�ӛ�N�o��ă�T߉����E��Dޛ��`�e�`8��gQ�dc�t�Y��������������H�]�ﰽ��-�e��U �����&n�`���[q&�������A�\j���/�7��N��|�jz�RE�0*��=��~b�t����0��g���id=���ي+�謥zf�Y��<��N��3z;��ޡ^���.��gb�v [������[T跾R�`j��E���x��k{0{���q�y�8`O��b����<����m��>��փ˙���L��g1�6%0�te�g̸F�N�����ϝʦ�,�`*$Q�BNϟ��dw�US�#�E�v`���8��:�+C�s�}�+��mp���;p*�2�_c?y�h�Lg��q& oY�W�u�x$ꓘļ4�\�7VOy9�+��0z�'8�I����J�f�xa\��p�N��6и��0H��,�q�ɶ�沘A$�Z�|r	�{��1�[�Mf����p��k;o��4��*'2`�JWRۥ%�d�e �����a_�9�nqH�M��b��^`7� &�H�Ѽ7� z&����VS�T�����^	�%@�w��U�e��6b��T�����o�X*2]��������b4udȕ�E �Ꞗ	�6�o���k��1ǀ�X�`]��,Ld஋�f����!t��(Ԋ��ݢ�e���Θ׻���S-u����J���G�s���eMo]��u.���{v�pe��M�A)�CcZޟ�ɠn���ʳ
ņ�����w���dM��b��z����m����?�3�������(pćvr,�%�����)�"�CNK愻����&8��wX��F.Z���K4�E�^��t�,߭�л<z�:[�Rg����I�e�Pc3�c�f�p�3�HI�J,�"��kO�Y4�SV�&b�M�K�A�}�����O��f��$\^H?�έb6_2i-�I���q�،+��*29l1�_FzV;/��ݴ�H(�� ��"T�տ?q��������aTX'0Z��=u'P �3}44B��_��AT$�]��Q��q��D_	�7/>�3'�b\� ��5�j�!��0έ�IiI]��X������n�_�0�	��M���-5Ξ��Gd�L|澗��G5�1�0UP�����ܳ�$� ���>��:������bһB7���!�)�0pj�uBF�F���B{�gq�g���)\+��� <��l�z�v�|(7/�}"�����0G������Z�R��r�!�Mkݨ�.Ū���]X�O���=g�߆�Wa����TS�#����H~�
F���B$�>X��hK�.��t��r��V��Pq��^��nD��ܨ���Y9y�C5�!1�xL࿄�^U�Z��,�m-+����x�VW�ޔ��:����n
���?�
�P�`L/�]J��b���f��"�$s��§L��9�KX��Z��b�v���v}� X6��Μ[���zf��
_GB^.��lپī�9F��y��	�z8$��"�d�:�Tl|��po3XK��Q�N~nX���0�� 2�	��8PɁrzꐉ�U�����h������7��O��+D�)�lT����Q�M2m�-s� ����h�T(�GL4�#�� r�0E���u�
K�Ž�EUY(�h��}��S�~�)�@�	�Hr�n��WM��t5{g����)DJ�E浗�u{s�ɕlꨨ9,�i�m���-J����c��\8��^���1��F@s
�t��V�������@�n�8'��L �Ή�(�F(?s��,���vO»�x�������q�0"s�3�p�-�1��"�	ma�	�������.��n��|�cm�6���'� }�$�z��}�����qa�w�l�S�����cS)���(��9�9�>����Tv����EԽ��y���|�n�.��^�ȁ�x;��j��f�!f�F����n~y�������ô�\V�Z)�=r�`0��+����P��]����h��Vj'�O�O�����F`�8�&����i�qo�ˉ>sP�|t
<Ԩ��V}�g�,3�я4��n2Y\�J$A�g`@G7[mR�ߨ�hnpE@��-B�b��|��-:n���I��<��x�k�#3�G�� N�T�0*����.�>xa�U}N�6'�
��"WE�d�� W�#	3ѷ$����@(�A�ܳ2#��\��i�xG,Q��` �s�FP���p���|�0�,���������9%��U��A��j_��q����<�c9/��:=��Z�L*���у��ɩ�����A��P�5�Γ�yf���(�_���������.4'\�H޸1��q-[���`��y���) 43����2����t��d�i�}}�!�u(�=W�_��>�� ۭds"r�ύٴ�5�{Aa4��ö�ɶ�Ze����<���hS�����	�ߓL��,�
�P�ȅR��΢�
U-�7��S( Z�~3�H�u���K�p�����v	?���W����Ay�kv�V�:l��}j����r���|]��0Փ�sr��_��x�4�z�&-؀����2��oV6��Q�61S#�`���QN�j�/kT��*f</��V��8D�]B �RZ�>�2��mS�k<�5��t�xA�OPT�Ry���i�O���8.� ���x��pD��hۼW�kO&�!d����:>x,�qg�N�rt���(�20�|t�g�KrC�벒�n�P+�,(:*9` �Epy�&��(���M�d�E`�Xs��w�/���)�1<I����УI&��e9H�_c4��zJ
�3�L�R�?g�3l"�j�x�(;� g�$�=���Q<>�`�(�ҋ�v�__8�ūj�:ݾ��D��y��l@ ���!�==���<�$�oPN��R$�e#�e�  B�*� 1�؛����h�ӯ>)b�8n�j��{DNJON�Q��vc�yɮg�����DyS��[nm��B�X��!q̢�@予���Yu��)�˻|���h����`���e��)��QWs��R`&��觋�[�	��4^>��-��|�^�Tj���.ђ���	��|W�zw䏒���7�j2�o�v�*�5�"x|��E��Ez=�������GtVfި��O��	��3)C�l�^��C�
!I���v��qԂ�Å�TGJR�j���윟�x{+���a!��4�>`jyXbpR�d�����@"q>���-<�s�;�L�g�	�6 HJt���S��N��'�X���, ��*���B)�����wc��SＳ��c`N��8�F�:`�S�N��I,ݘA�g2�u�Ip�'��z-w?��SC�L>�c��\&���YGf_uORC��?�p�r�\wqO`u+��z�E8p�`ְXEE�A��a�DpJ�&�1����YH_��/X�D�y捲�$��|��vsY1>�\M!v��C��P7�f�[4�_N'�h����R6`-�c耿��W[q�<�q9�٢H[ ��]��^�& �_c��d��%(�������TvU����	=��%���&K
��[��(�֡�����j��*�JX��G��횎�_��u?9%K�� t����6j���j5kk�����{�;-��G��,��ʮ���Ce���0��CUN����,��q��V�h�NJs����~�b ��o��MJϛ����Z�v�X�!�G����C~��c7�n�,��l�`F��ܹR�I���qdh��b��zm�(�گ'��:��R��G��p߇�r�/�%])��xXн�LN�f��#z��K8S�w���F	x���$���^��Z�i�����v<��5:�myRB��Fv�� H�c.k���فp��FHd�XJ����w�4���Ǩ�,�&]v����#�8��/L�OK��|�A\�B �i�B6Z�i��@��PK�o��r*�llI_�&@;*&<�8��H�&� �\�"Ϧ՚�<q�Ā'�E�����u�fX�����'�08��R#4o]��d=�cA���]�}�r�}^���D�/�7�+(.�$b�֢ =Y���ڬ�����ſ�I�� XhW��nLK�0�`�|��R9�yBMd�
���ޮT5����Kn��]�ں���k����9�:>�����"�7�6ʬ��!&|u0�	
�p��F+��Nļ{�V*��Xl�~��2��<4��u|��й����R�E;<�����]7���M!��S��y����v�v�]30���Yd�Ԇ܅��\��iS��s�zu�~�-y� �(�it�9Q{�S�����t� r5�����S�����i��c �z���t����Yl5v���YW�Z�^PW[� � �٦�+��� V2���G�Gsn�U������LJ/�J-�b{��������Cs�6��Z���%X)�Z&����+����6�����J#��U�_·_.ո;l<�F�F��Wy��&�5t�$��"-%�:v$�|�^o�FTK�CԚ��AXv�0�̺2f���%��P֐$o�P����B�h�M���7r����D 9�]���xQ@�bmg4��ʂ�4�ey9WTU�G秏#��{rX��0 E��>�
ƿ�n�Yc�h�g����~�w@g&Գ6�-*���2t^(��t�����
�)�f�E�]�Ԑ��D��z�,�vW��([�J�l����w¼�-�Ε�k{1!	�@6ƾo�Vk%QxL�[�������_��=	wL���΄�]���W��-�\�h�)�0���l��"�K��+q��L�����m<b�	����rl�p�.#�L�B�_c�L0�� 1��6�[��$zF6�x�x�t�e�,K�����|�k���ܞ���a�W��O�����l]�)`E�kE�<�������n�B���<�S;�ץ���Wf{K;��f.�Z�5~tGa��>_�~?>\8�Z���r�5���s��(��_8�cI)�w!�h��j��i*�q���Ȩ��F[���h�>4���QoY��>N{�|���C ]Vx�v�jL"���b4���2�b%J�������[h)�:�1h)'�@�eyB�����h�ŠA�eश�;{xHZ\�>��G9WI)GYT���4.�.��`a�I}:xQ�`
��"2�d0NgW$&3������@���+��UY�7YiN�rx␯��X+����PZ�cË%�!���G�,#�I�-����9��U�2������K:Z�l��<�6�/u�8JgZ �5��r����D�)��n6A<k�P��MΎ��fd,(t�2���Y�����i<\.$�޳U��-ۑ��F���Ƅү�Wd��Ή���2��m�n���5����}e�U2u(<$�ZWC>T�� ��us=.����B�ܶK�47`��N��2\��ٔWG��������	5�.	��'Rf
��@HS�������EUP��/tn �"~.���ؿL#K��a�Ŗv�nT��kH2%�'E�\��?�l*�j;��MyqķN��.9��$V�����ˁx��z<6 -���5 tص�V
����LU��x#�`�kN�.Ōj���`��f7v��Fõ�*#DنmB��Z��m���k7����Fx�.�P0h	R��fa��C���~��.��L�X�"�+L����9W Nl&��d�$ȼ�>s�cq�k��-���VF2pKt+3g��kC�^ܒ�@MP�(U�*��p� �`yYw�O@�(̞���`my� 8n/8[,�˜<>׿�����I�"e�l\�z��r�:
v�L��?sg��j̽(��  ��Z|
&��b�Qw�?`(:!��*�v.�Q8�O��O�Xc���X�f�lۖ���!H��=i��Wi���?x�薺$��� @�
U;B0�� ҐtضA�KGۍ�9)��78	���{vN�N�	���R����Bץ�1k�D+r�V91�m-3Ҥ<���j;�c����PD�l�˶Wr���hg��܎�#'�e�>�����Վͳ&$�i�b[�l����mcbķ|8Um����I��BW���6|)E�z����rǴ�:�jǏ�m����8�̊B�=\�9� b��b�f�j`������%3Dⲏ�M^���E3����AvU��� �~=QT�]R�e�jqo��X	՟U=K{&�ʼxЈ�;i`��b�/�?6b�>!���Q�>�8=�9��.cn��g'26�t�&&��[%N��J��>p�@8o,I;*.Bu+�F�w��`S�uv��;*`	g�8ڡ�:ۈp�)�V��u#��.w	�����p��k�s�?o	@LyG8�&��Y���u
L& ���E��V\\<�`O��P+��\zB��8+37������aҮ�p�@�,z܆o�H��J_�k��h��$%�|�"��q#P1��)M�T�,5��a���A�V4:�'h�6� R�:uU8�蛜�����_�9(e(H��X�^"� ��-��������_fT�l���|	���%��A�Ʋr0��y@w�(hx�e�|*�����9n���u�d�0� J���76ł��%��k�td�v1�iԂ7L,����]7�����^��ɠ���j�M3&����I��Gy���M|�}_@����M%aZ�먝�/�7v�`�|�aз�C�Ψ��Ĺnyi׬@DN�%Q��﹭��Ձu�d�.b���zZU�c����A�5��ڭL���p���rS�%8�l�Yf��X:MN1~�:�~�Q��n�^wNC0F��^�{8\^��\��rЭs��<��x:Q'Rk���z���Ӆc)j7��	pLg�H�QJ"� �Rs�� 0��#&X@C������JgO�DAW�N\�\��Q�6Ui��7�m)�&0!��*���l�5&_|��;%����S�H�q �i"J�#�ujqM���",��&:��U�X��]�/8�'Fa(�ђ4��Ռ����A
o']os�!�����rD�u$7e9�)��b�< �D]��=@�y����U�I�,X�v�|�n�Vd0O�h��X��0i�TSt�i�d.���%H9�!5y�U�f����?�ڕ���]V=��4�:�z��Yy��=�tұq��Ӱ1!a�^0L�!�k��F�?�	�:{fk�]KϦ߿��mg�<Ϯ�p4V�o���\"���R��x;�x���H���N�M�H��(6��æ������]�����������]m�R��a!S�"��Hn~rp�[*4x��4j�ɮ����tp�r�7�cU̎Dp�O�M�d� 꾁�5e���e�9��5Q3є���۲^K��[)Ӹ� �+Ǉ���V���QJ(�(�kn _c��G���i$Le��J���bV��܈t�X��s�{'�]����LXD<�Z�pI��L�:ոV1Z6�*�RZ��fP� f�_=M.���lO_��ᢋFԪyyD�����$�@�"�3:Q�|2J
oi�(K��2�)uX1��0�\2�@u��e��F6��,�Kp�Qӛh@��4b7태[
DUݜ�����!Q��3m"[��6�o��z�T*|T� {G�;�#��2r��q0��1�'�
Ả�I]�Y�)�h0f����~X,�@"cp�Q�Q������c�Htk.�����)���E\%�ԫٚҿ��^l�,��X�+B�#�~Jj0<M�K��l⨪ꕬ1\A�@�u:�j�Vg��V!�v !�dR<�ȧ��xL�L<5.��na���(���]n�qrtdl|����g^�")4g��d׸g[��tCm �	"&^*���.~����Y�c����,���h�̖%$2��s j��7���Tᄭ�������������U߫�8���W͸��D�|����E��T��o��v�n����g,��3;��h���}fV� �������~o��F�;�9�\::�Z-&r�*&�W,e�5�߃��Ҿ3��2WAh)��j(�3-�Ŷ��C�FVLc��0���f�o�be>)��|�6Y��m�VsՁ�Ō���H�4�c�2O�~J����SEv��[c
W��_h��R@�B�B	������Ѡ���
������x��YEG����T �����/."�aL{}��lk
��V"fdk �W�6�3�1�ts$@��<�(����i��x}���p�)�zP�PæD�����#,^��ȡQ���9�a�U_�h��e��"��G�(<*�/s73�Z[�`�K����𫥥�Awi�P&��Ήq�fh��(/5�������Y��`o�&�\�T�ޮ��rذ-�	ü�L	���Ҋ�� i%����2J���)��'	�_��}@Ism��(�*+�U1>��� QksX
�σx��đO��u�4ҍt����wSK|��rΒ^�����DT������"�o
AM���x�\Ǣ�,U����j�� �J�~)H����z2�K��䧃mv���GB��䖎�,����g�̯Yl/�tj����(tc��K�2L����5�?�٠�ƙx.�z�&-����paI�P�ZVN7�Th[��B#*�Z�űN�ό�#I���f2��f��V<�D��BzIZ���������Vk2(,�F7�x���PK��Ro��A��~3o��:.��Ƴ����s����>W�P&�l�d���Ml>n�oq38��5���~��2�lJtf�gkC����U3�P�I(p��*/q����y����yՆ&��1`(���/�>+��x<y��E���|I�a�e������q��6
QHL,��?�Sb�jl?q(��" �D���:��`Q��X`ÅR���,v�|8r�����'���*��5HlvM����,!���=$�c�r���eO�Õ$���&B����B��, �U��{1�ơڍ��)�ww8�{K�ěDN n��ك-����$�,��l[�D�"��Q$��q������W����^�>�X��K���c˱����R؎�9����b�e\�����0��4�&'����[�/Z�*K��H�e��𥲞���Hx��p|DSuzmg����ԭ2��O�{�e����e��ۥ�S���~^�=77��;A	�}qf�Ln�Ar�43_Ɗ�b��^{j��em�8oTv\�'M��9�T9��R��jLqy��F!��!{!����/����`���bf-��yi��v�Y>�{֔RA��P�wdg�z�6��tz�̉-N}�I�Q���i,6ل*���B�w���w��S�N5�V4�`�j�8��:Vg��[������w��Z �+�Ep[%~��?�2
��5L�cr��3�&�[�Y��u�e�;'_5��zZ�\wU$OJ�+���z�}8�שR.N�~��6(a9&p�c��'��ʽ�H�"Ļe�:v��CFY$Z�|C_��l��1�iM����GG�������4u�1'�6�� R�4�~-趙�M|����9cH�%)�S��^qG W�ē"6��ﾖw��iT�0����	�8�%qz��\ы�������{8��PW�`�8*C!/�A���#�u�U��u�zT��� ������6 )w����k�j�������)Խ�,@��|�)���<�R
ьy]׊D�L�z�[׌ϒ�D���uE�{�}���r�e]HM )�&�B��czvÈP����r�C�8
�YrHnT�;�{<>�%@����d�<�d��db�~z5]������]�݋0[��ʺ����p�r}��%om��t��FN���T������w�хF�%�A7Q�y�^�G{�F��.-�<���:� �R�sC���+�6tc$���w�Qp1H���J��a�-'p�
0l�$:�&S*H�\·��E��e9OA�P2EL\�^���k6P�_i>%/�(�
 �M�i�*���l�z_��; O���HY�8 '��"ő��P��q�`��]z���q��+ LXX�E�J��'������_4���0� ���AeD ]*���<���su��}�D�7 g�$j�bm�V �P�������ͭ{SI��X�h�(n��0
n��78��Hb��/�V��d���毜�;�54эā -�S�V�p�hFZ���/Mc:����&{�XB�,9܅�g8!��<0眱�f�nF����{,�4��]���!o��<j�k0�ʢFҜ���;��S������F[�CG��8	�~�����2�lI]���1��8�F��A��ը��:=S)���p<�~M�/���Uk�/�O�	�_v2t#Kfr+[��>��|���қ_�#����S�+V��L�5,��ϔ���7�^F����e�Oz�+.;���V�`g��)��ô�n��̡P!A��n\L�G�J#�Ab1���sF����s��¸���j��X_��Z�wD��u�����b6�7Fέ�G�!k�;��_�g.�b,l�_B�|��FϥWy�h!���E$��"#<:,$�|mUUo�K��m�_�X�%�0=�2\�H�� /�#]
�Z
;F&��� h����OM�7hU6p�D�"�=���A�Q��mݡ+�Q��*\�/;QT�L�G�#��%r��0vȊ�0
��]�$�Y�`,h˄�����~�]@ݿ�l�� u���!!�
�t����d�)U��E��Ƹ��:}��9~�,1�> b�K�Jŷ+\,�6��#������1���@D�f�e)�V¯j�S:���Y�ߪ�������1L����z�[�~�YyL�C���R`�L����d�f7��bGs"�<��xr������b�m�	]��œ����.�����c����S�f�b�ѩF$�=V�n���*�`��~j��[��r��g����5ϗ̾�����J�d�C���_���Ee���*
��MXn���yȲF;�%��w0f1����_��	�~j熱��8���K\U\�Z��r�?鴒܊��w���!�>9���hD�zj��H��8� rN�޺FQ���fU���{0��oO^5>1�|%��y�Vn�� 퀥N��4�F12���J�"��%ѯ[^����h��O@1�B��b_Α�n��wS�n��M� x�=��t��G/����T[�K�j��.z�Ea�\�}�6���
�"�)d��WZp�3͂�f@Y%�&*��^��w�iĘ�x�4���U��EP�b���yU��� �,��)�c�����96�Unb�+:��A+��"��<<=�/��y.ƮZ��l׈�"��:D���7A��)P��?΄
�fô5(��e���%5Ƭξ�O"\d��ީ��ͻi-�X���r���y �ej�<$��$�2�����?�'8n���}a��y(rQ��P+M>
�, |Dss������� ��,��4m�͸��k�Jl����/��R�������d��R
���ȶ 4.@����U����� +�^~$��Ya��58�K�G/��ev�.ᴂ��~����Rq��p݇@lJZLj1Oa����-�͉铡���3���5xI�,z28-irɫ���@�V 
�gů#E{}$N�����Q��f-d|���ݵn�D9�B�7Z^2R��)�>o,k-z�����xr�Pf�SR�Kϕ���F���.��b�N�������8�WsJ&��}dF_ü��i>i�qxݍ��w�)N��2��yt�m$g�*�C��c��E�P\��(��*�)v��gyυ��H��]�u�7`㲰�6�/.B����<�S���#��K�I7� e=4����h?
,-ZLg~?8T]��j���(N�� �>r{��ԳQ�%`^�����v�:w8-Cث���Nc�՞�*%gl$���Q�!��#=���̍�2��~➴Z$5�*��^� &B�� H�9����Af�d��)}�8?( ��ۮN[��ԃH�)�uiT�����k$DJ:��L/���!h�~c�rX��`M��)�
g��QQ�ˬ�}}�I�o�)m����e7��A��(�����}&��r�؎I[�rP���U�#/��-�������{�ѣ�8�:QO|_�z�Xx��Ͻ��n���T��`v�;��S�`�n������=��v�����f�N��`��:z&3z�ʏ�<^V�g�������v�9���H��WTT�Rx�]j'�U�Σ���&�{��r���e!*`���b�J7�����Ѣ��>�ޭ�����^�<�g�6�O�tQ�4�$�Nx�$�i����I�,Q��*_B��w����w4^MS�G�L�`�18��:�e���(p��gl�p��6��74p�4��_�?e|'��L���}OA&���YXQWu��8V�1�N�U~�\���O�+�3�z��8��$m��Ƀ���CaH�pU��"���%�?H�r���ͬ��=���$�o8|޻��g�1OY#MR���by�WQ�����4�@�'�_��v�RGO�����ѶO��<���ޜ9��/H,X�N	�^̌� ��=[�赾q�W�B��TG���B�	N��%,�Դw�X���ʢ9����^YN�[�*��
�����>ե��(�u�K���t E����b6{������k��l꫖�@��`,���w�x�T�a�'�������I�UA�����'ܳ?aV���6}���}-���VM���a���eUv�Ё2B��-48C����?�n/CЬ�Tb1E��I�c�Q���xd��wb� z�R�����6��+9
�cg6�x��p0Hgr���%�A��Ϣ�Ў7Nc�����f��HwD��F����|p�ܱ� ^����z9B�鋀<�w:G��RӜ|��≇�J�c�����Yp�H��J��řE|��p�&N4���
�i���sO�C��9\J���:t�6K��i��&������D�*� �l�_��;�B�Ir|Hg� B�["@�I�+�Uq����� ���Ȗ��X�q�e�'<"m��r�4 oN�ˬV��A�99]�W�W:/��0�q��DKbo7��0k>b��� n|���c�o��V�kII/�X9!����wn]Ͱ0�$D�RƝ�óM�
5����dd�3��5��Ĝy���Xj�K���c�:��*��:O�Q����s�'ҧ ���>/!�20����avF<�rkC{G��S�9���P����<X�f��%�;���JK��S>�.$C��U!�!�>
;�Z��9b6�=��W]�W�ls���Æ���##_�@3�SD�8��OD~(V���Ƨ��ږ*���d���t>Fr��G�Hy�����o�Zc�t����b�����/�k5ſ�
���+��^A������
G+I������V��ߔ�(f�^�en�������<�xL�pJ�"�b�x�R}��0qs~e��@�%��Xzj�Ze`RB��}���6�����	�ܥ�Vjh_3�l.f��l��ҽF���y����fe�$ "�&:Tp|���o��YK�����S�X�v07�Y2����ہ^�R���A�T�T%h��I�j�N7���8D�c��6H���QQ{�m�\�l$���]�
l�T�G�¥#�<Uri��01���Y�
7E~���Y��hfí����~�%@�<U������èj�lIt�a���AW)�{E�����ҵ_���i,l^�4��WJ _;��0�� ���&�b��1��@�TK�`�?V�m�q����Z�Z#��~�p��2Lr���u�$|�"]�^m���=�'�0�h�����]P,"�d��\������q�m͛0	�8;`T�����.4e��s�cٮ��"�ƎAZ��N6$Ki:�i>م��]ȷ��ܕ��$ۚBz�OP7�2c�������ܸ����zD#��E@y��e����Y�n�B#S���m��;}���Anf��2V�+v~e����Uͯ�\p�Z�retܴͬ�kOO��_0�th!��"�h_�j�j�Ҕ�;M&�y��FLX��y��o��K�do�y�>߻|`�F��]Viw��{m�	@�4J�2E6UJ�X6�S{��[YB�K��hZ�@L�LB��`�=@F�k�ח e��^�xy���׹G�����NT�����.u�Ba^h}kAk�w�
}Q"�`�d�$�W��M3�+��*��@�GA�}����Y�i��x�~[�� U��q/P�Y��ܓW�2AL,��g������9�F�U�;��F���S���$�<wp�/F��)�ZB��/*�=���t�[��A���P\�����f��(��ś1zV���Ƈ\���\��ޤ�=(��-G���/����@=�����C�s�2 ���-�Bi�U=}���2�(�_�KE�>eH� � s�"�y��z�*�g*4��ȝ9��_B�{�����T=㪋A������_�W
�M�q�/�O a����U������y �9�~B�;���]AK�$B�y�}vu���8�������m���B�le"j���ɗ�h�
�h�5��������KVxdATz�V-DX��惰؆	�V����
�G�"��#`��h�Nx��\�19f(�y��̿�D*�B�pZ9n���h��Zk(쒺�y�x-eP�dRe�;�������O�J.�4(�i*i�\#�ԗ�W��&�pgd�,߼R�>d�[q�!��^��srt�J2���t�EkgR
�C�w��x�P%(�!*%+ݱO`y
ia� �sˢo��U�`����Q8/�e���#<�A�{����DI�R�e�Ǳ������tS
k�L�w?�tGX2-j"��(	�R �����t��Q(��`�|]޾ǖv?�8��f�֒�Cְ2�e4Zl�����!Y��=�1�̨m�[�~�y�$pk\�����BA<q p"�ʪڼ�}�?�	)N�38�􌶺;�N��:O�c?��N0��5�⛏D�q��GZ��'�eDT���A��B���J�E�#���l˧�h2:�+
�D割�9@eu|:�ÒΎ��*&5ȷ�z*[��N� � ����h?&w[��D�������|z��zcjs�w�#��ǅ8��[lC� ���߈���t��=���ٱ����6f�p�������3��r�X��^1x���)b�n��v����E�ů$�To��R�܋j�A�	!��&K�{�o��>O� ��`֡b\�М��Y����">�a �J�F�_��:!fg�k!6l�3t��:̿��Ns܁�3�q�,lY�*�2eB��E��;{w�÷S�`���x`:�8+s�:L��Չ5o��@6�����pѢ���Y?��p��rL*�Q���&�lY���u;�gq)L+[0��\�'O�:�+��QzSkl8\���.D�hŭ�Ma��p�f^�鴆�f�HKⒻ�4�0�A��Yd$�Dy|y8��b��1�hPM�T�}�������h4� �'9G^{QR����i���O�Cȝ�Π9�ƱHǪ��I�N^'�^ �ⶓXEh�h�L�O�}��T�a��	�9x%�v���-��ur�}������]�V�*�w��"��Y���K�1u�<D7�� ��}�d6��<�V<Qk�M���������3�,S�rs#��f��c;��匊:G��0�V��9����:�DX����D���<p�[��M������� ��v�8O��p���C�lşO-jn
����̄F�ʐ��ղ�XdԍSb��Nz��g�ۯ���&7fھ$�3h�pK�'rs}�%�4��
��) N�+��K���Z���gw�NUFu/䄷���LZ�^�O��Lk��
�<h2:�	R��e�2G��l6�c'8�-"p}$�H��J�s���뙀�`�Z�c&I^f��l�$Ov�<O7��b\�k���5u6F��i�-���6"�>�*yj�lXe6_M�;fҊ�1H� ]��"��^��q�`~���/��g���1X���ˀ��'����b�4[
	�f�d�GtAO�]�U�rc�iOL�jD�C76"y��b# )����&+��	�1�I��X��g����n�8G0����mt|�>%���+9>0d�^r��7JH
5�tJķ~�I��&G�ȣ'���%1&:�^���߆Ў*��"(��d5!�0�9�\_�F��_:��{bS_���@�pEB��<���a�񀱐����C�1�A�	q���=����9�v9�9�����3H�b�q]�O���fGnD��}�~�u��K�S_ԟ�f��~����I�B�%uɿ"x�՝stYa�r!8���c�? P� %�UX���kn�f�ŀ�����n5��E����N�^<Ӷ�l�˸�ͷ+d����OV��(�H����fn񌴡4���xL��xJ�b�)���Ɨ)�psy
|�nb��[�X�1�Z�>-թ�@o�'g<6��R�cH쐗 �q�_��.A��l �ĲkF��GyU}�!K�$��"g�:�9|���o:Q�K��w�PXb��0R-�2R����������%�<��bD�hq|lۅ�7^���$D�A�s���Y�Q��fmS�0���'� ��TA�GS�r#٣�r�'�0�ˈ��
�����YO/�h"��d~i  @Sٝ��.��ޞO��t<+���>o),E�<����R�0b7��^,��tij���J{&k~�Y��*��3G�=�1�M@z��[/pVxt�=�8�ǟ#�ջ��Y?K�)�<L��pB�r����ѬyM��H��7�����Xy�":��� 5��\���tm���	���4k��[.���.�:c�db��&��P�G�$�V�d����[�2Ʉ�}Ԃh��p�܊�����v@� T4��H��В��fEx᠞���{n��%���(&�;)��m�8f�21�m;���C~`�W���j��\� Z��r@����r�G���J��ϲI�c�	hz{j��X��@�vHR�`�FG��0�*��f��oE��>�f�|���ԯv�Vd��������4 m�2���Jk�d��'tG"�[T����a�hB6@g�8B	W��An�T�-��z��{��U�x4�����G%	e�6�TѴ۬���.ph�a]�}&���[�
�~�"��:dWW�CK3�ت����@ϴ�\���_�ͣ[�i:�VxNc��x��:�9PF����M�0~�w:),5ڄ�0[��:9��mU�)"�adL�7�b��|�<��y/�B�$�fZl$��/�X_�0K��6��A($(P���z��fy�?(`ਜ਼L������b
UY\���ޟ%���-V/����l��<PI:�>��2[>��Z���]��б�}����B(��}�F�>��� ���s�^���V��U>�ܢ�4����âP�!:|�q��#���G��f����Jߚ;v��4
R��,s��j2*�x+�Ut��5� a�{~��6�ث��K"��vPn�����������������l�
�j'���$�ģg��ez��(��PDh�z�x�z(P�-^_�!EB�!�oV����ez.��rw#{�:��NS2�V(�̌�f#��w���1DEkB��Z� �Y���t��k#~кWK�x�a�P��>R෗Ҽc�/zҰ��.ڑi��&ֈ���WY&^"ad���,>_�;q.I���g�>�K�2w#ht>�g�	�C�jےf�-P��p(�v�*���݌W yEl���4�`^�+�d`Y�x�lxj/$���p֪<*P�����=�I���e�{������^t
��.Lݐ�?n��S��j}YL(�4a �&�h���O�kQc��`�(7޹�v��8������D5o֋�:�c!lG1���!���=U����YD��=Y�TR�$�H��f]��hB�� �O�"�3�7q!��$)��8uᑶ��WN����4�~��kT������.D��F�B����V��I�����V����W������ˢ�c��ؿ��_}X���e����^���w�&��|�N��[YU������z�ģ�i�Ԟ����Y0��^�|�=�zޛ��Rq(�^G�� <��V�L��Vΰ��"��S���s]=�����v��N]�fŲ��e����3�2��ӫ�^/ۜ1���	�\v�i�8�w�j\mT���Rn�Ej�6>�D�~���+{���(�ۆ{`�&b��w��I�*v�GP>�֥�)���U&go6G�6t�3��ZUNn}o�44�,۱,�I�*&�Bp@��2��wjIS֙Z�gݒ`�5x8FN�:��\�$ʉp��H1����<�p�����5?[o��c�Le�O���y&�h0Y�u�r[�ڮ��&�\(�gO/+�Gz�D�8�������ňIa��`pQ�X�N���j�Hr����c�U���$:�|���]#D1��MȻGܘ=$�M�5�#4&!'�N�vLGR��A\�Q������9҇Hbg�Du�^�w� �Ɠs�]�_�'H����)T}i���D�	�%�M���
����X��,<���ʄ�Q@*TS��riv�t�}��˵u�MDr!� {XN�x�61�?��k8�+�b#����G�nT�,�;��me*�
L���ƌ�ك��������9|��]׳5���*���,���;��DM����������v����0У��C7��:�n圉�,�Fg�]������m�|d�B�buLiz�4ͼOy�.�q�!U��N���pfh�r� W%�G�E_��PN�����=nM�>�w:=�FP후�B����E^��0�4�_��<�:=M[R�N��m�b�B�c����q�p8N�H�nJ�M��♻}��=.&D��m
���
�O���!�\��p�6A��iO��YO�QC�Yj*T��l�
d_�e�;F����H�ܷ x��"6b ��q9/�.A���H�<��X�R�˛�5'2c��=�4����J�Av��][63�
���'^eD�Ί7ѯ���b~x� �3��
��e�9��MI��Xo�=���n�}0;򯣈B��������t{d��������5e����˒���u��n���·�� �:@1�E��Щ�zҝON�?L�!M��0��1�W��F�L�z\{}���IUԦKD�Y�N<;�\�\Tf���w'��䚬����a�4F���4�n��1Я���N����Y]zgN��y	�F��K���඄�Sz$����~޻
�G��䥢� q��g�aZtt��r�ֈ����z)��a�P�5�*OҨ!ी�=��%��5��'р��a
9^7��Ǣ�����+�V���!VyLA�=���ȿn�2�amX��<]L���J��bɤ��t��3�st����Ƅ��K�X��Zuڧ2x�&�u��c6��Cξ��R{C��_)�|.Q�l; R�M��F�VZy�7z��P�$6u�"��:�S|7/o�#�K��F�p�Xx0m��2�.K�Z���_?�+c7t���T�h,�۠�[7ٝ��a�DAF6�h9��Qҷm6��� ������-�T|��G��w#�*hr�R0��-2(
->����Y���h�����_4~ı�@�ʳ�`���5�y�O�t���[)f�CEH���Kҫ�7��sb,�*�R���J��9t���T�┠��\1Hb�@�<�V�\Vӆ3��ⴴ�PtB�4v�d��L��k�K�֘�Ӫ��M�ë���}�P���7���S"����s\��G%��Gm��	�h�5g���.�k��c;S�������̂�1$� ��_܈�;qy�ӻ��?[���L��� ����h�m�� #�[=l�t�}��|j�|�3E����ۘ����n��	�_����;D�Ɨ��f��V��@��a�~[Gұ�;��%��\���Z�r>S�C�4��^���U��*��nh���j��q�<��c�ȯ�FB�	�/ƀ��7�=Oo�.>�1�|��Jd�V_���1�O��@4;�<2;c\JF$#��X�z[O�'�MhИ@�MB�Hh��aF���	�H>'����^k�x���uG�E*pXT��;�[.kjPa��2}����_�
s�"y.�dW�W+��3��ӂ�d-@��cw�2 �~}�iuPBx�gq��(���dP?n�(�Mg�R6,J���4��R9G�{UK7��|)������}<�6�/|R��Z��LA��s�����݂Ac��P��n�u��fԝ(�g�'�w��=���R\5W�ޚ�"�%U-��)�����T��.��i��q�q�2�����U�x+N�KF�}�YQe(C���A�>[$ =j)sĺ+�o6��0���^4>�w�����|�17�a��j��JrݪA��0i�5�$�®
�l��Mw��d���UOȊ�V�� ��~t}jPf�f	�K)?��oG�v+>��3��O�Ύ�&�#+�ݸ�Hl�Dj�P������=������y�⫴B���"x��z���-��`�\&hؼ�QV�������y�#���w��N.ڌ��30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�(ڜ4�z^��?�}qp����|��Cխ��B��
����
BH��e�]}<�>B�UO6N�̾W��n�u�H
J�o�Ɉ�!h�!-�d����G�W���\;�ũ�E��n1���^dV��	&���B7U��q�=���_b1���v�m�G`�O�{��񜾹�f��3���[���L�m��c���EҐxa]�Ehr�V��&P��~=znM�d�	9�cr�i�S&���	��I���"u��R����O@�Qr�U��6cԄm�&#��z�CI������đ�&��PN@�S/Z�vh��¢q�}�^TY)=FX�&I��P�d�z�)��`kH�)���stt�A�&���U�8R9W�7��%^;!��s�����!����`IyM��x�n��C�M�����"q/��Xȏ�V0�MG��4X1�"���'{���nf���9p)�1������0b����k��t@�2�����rD��!ۯ��j���m�3@s�4�J���,ta���N�O-_|��.�we[��-?��၍[w���G�cg�d�J���Y'(���G Y>pD�����cp������stU�=?T~	9�pR�l��X�r��a�8�_�)�;j=ʆ����]����ݘ���'��/$~6�i�{'^�$RI�Ey���VH!�Ki����[�Æ��$�^$Էa�[��0!y��~��L�����|�6$r���tBER��(�&�$C~�c�Vw�rV(�*��ػD�y9o�aӁP����VܭO������ر�+��^�jKc��i23�s|����Zj��wX��v�<��a ��2�x�L�zD;b��	~��e��r�d<���%v�C$H�Y�rw�+n�� _1`�;�-u�k���&.~G�OLY���֙2+�K�10A3�\=4�M��J~F˪��_`��@K@������3�e'�,{�bDv�z�N���@�KMe��ҔT�1���vT{,@�ռ,�y���j�q����"h讁�����;��$zK\�4� g�"�R�}#��=�/9W�x����n�{�)��r���*W�ëe���N"2c�N���=�7��&�u޿��1���7��g;N.��3��G`���ϧ���wI2L~��Is +����$6���pu��Y��G����H��%W:N�{Ÿ*���L]�u~::T��G7,�F���O��^ж�:�ڿg팳�P�D�\0�	}PO�}T�+���b���6)l������\j���]�4;��8v��c�'2�)#�n��T'�zZ�!��4h1ض��	���<Ȋ`��IF�5 ��J�$��V�U&PqW)�tz�%�p[T5u&آw��^|jM_�Kݥ�ݟ�2��I��Σ�
�?��Y8��j����e��|{�AQ*�į���M?� vT���	�H�����R�g?���Wi�KV|�5Gӑib�o��x֍�~c�u���k��l^JzE���0Ȗ�O4DZx��xm�k����w����(�|ouE�+����x��f���<
1�i�'V��@�ݹ!E�l�
Y_
�p�_ ����[�0��7N�r�pe����m,�Mg�*j!�$��rq1H���"����G�x5D,�[���-��gƝů���Ή�'��=�w> �g�ci*JCj����p��R��x"Jk�Ά�u�&��iu�����RӨoX�/K%�Nw�� ׭/F��i>�7��r���ο�:���N9˭*�]r�|M3~cqc�ħ¢�:r蟦�L֍�����㸵��݇CN���s���a�f"s�L��9�&)�����oH?OP�0as�r���3��3�_�;��<��X���Ӝ�� ���YV�H�GV飛';:�F����xb�L��15j8V�NH<;m��ړ��9u�֢W܅�.�I���A^�4���7���o�BpP~��w��o�����S�i�����p7�T�-��AH����0���!��&\��y����Z��mg�V�oi�迟�4�5"�2�*����_�ᱺV/e<;h�h �������?#(Q�4�;b�(���s��XF?}�7��܉Ͱ�<��F+�B}�����"
;�T�~��}u�"B(MsO��N|�{WA���N�
Cz_o�G�:�zm�dC2���WF�\�ܩ��4��.J1�/f�4d�X�	�����t�����6�n��S1.=�v�?�BeƂ��4E��Hl��� ��3�nj�=.7�Ĺ��k�N�Q�T]�Ѫ1�z�N�&o}_m�z=MǪ�w	��r�m�S?|��B{+��@��S{��0�f��&@�S�r~B��O�ׄ���#�ȑ̼
��8�ʿoN�j(
\Pg�6��g�Z�X�f�qC��^�=�&BFv�ikG��O`�)�bk�.}�Tۘs-l�t�N�&��n��8�ýWX	쀞ZC!Q�s����_�9źm;�y�M�NԎq�f��c�O"���'q���QB]�o�M�������S�U��'4ꇨ����)�j?h��ˍË��4ܷ�UE�'	�1,1�[y�ڟ�g��¼H4nן�7"�Ǝ����U厽5f�QJ5�
F��CӰ��R1H�ۖt��TdI�	f�s>�Ơh2]��Sy�u�y�"����`޴$-w��1,&������J�{��Jz�Х�n��B��c#��-�rz�]��2AP��;ΏU�k�&�BE{ ��@(Ta����=�k곽��9����g���� ���i#*��N��VA��%.�*��Ne��R�W��iĮޏ>;�ֺ}�"Cp�QD[)����
�~�\�Z�'݅P�g��I��C����̭����cTZK���^�dP�tug��pPAEUԪ($5� �KAN���I���A��楾x�����+?��f��[�'jkB�%��5������I)�����������$��+֩p���v�uz'�^=Z�r:����aY��߫&":�q������=�^ oXC/�^ps���G?̸tN*Y�y|��.70+f��Q���c����vT�J�ݤ�J�F��~<q���� �J��W��MVbK_��>���"�i�wQ S$�0y�� l�_��
��_u0&d$��G>��|9b�����Sl$�������M�xe�ϔ�'��f9)xc~S��K�f��s2�A}���P�OGgؠW�! W �J��Bt�͘�}�e�cV$�����.�
 ZqyE����%TeB��z�{[�PI��ٞ��qr��ʆ�F���Y'kHuo�z7��)�D��$�+Y��Թ���֖�����̪_A`{3Xɻ�/[b���UIyiplf���E��J.��S�����浲as�/^���{��|մ.��z�	�@>l�_l�;�3��)���{�Gz 8��͓b�s��U ޝ��a��Wͭ�p�Lyh�]�����.UC1��J'0No&���/;"�������Gr--���[/<	k�])�/���4�r��#�s��eg	mK*��|<#K*�lΥĳ��-�����k �	��N�����rZH�5��ԗ��	{����K�O�&ؼ�:.�{���.�h�KY5�H�[�ܽwG���>��A��Y��=[���8JI'+��� X]�;� �ގ_���n���J^��*�\�h���X#�Șdſ ��]-�u��V<�(��q5M2K5���U�I"lq6�e�}��l_�c�q�Y���]C}I�M�K?%`L*m���=�P����
/Q��X��P��RyK�%��B�����\���%{YOf��BX(�}6&�a$�I�	��K�&"%n]��5h��N�i���M�*�𒈲h�Sȋ���c���t-����zZ���Q�����G�7������&/'�X:�}�Y�f]����b�ٞ7)}�H�|�*xb������+f�K1�x��ؗ�^���
a�!e�Y�48��V0p�|�P%D�D,���+"��`R�,'�{��-����n%�+��R���_�h^8��g{��NH1EɅ�N7,�R��~Gt�d�hT�g�X8l$�;��z�*)OA�t
Pjati+����Zϼ� ���X�4/U��A�����d���y�k��<C��Lֳ�F��=g����(�X1���d+�*��l|m!%�,��J��zt67*(7�MLR�d�ab��੿c�B��X��z���-���L̝� |-P]��w����C���3ţ|ܦB��d������X9!��*`���
Bj����`6/�_n�u�M�%6ĝ��-����9�1�c{˘���������N��68BBwH�%gp�Q���[1�	�l�o �^�\'�]�]K�֐��ѵ��"�!���'��E��cBD]��"�!�/ŀ�.�m�72NŸ[qw���Ol��Q��� bD&Fxe�g�7��<Y�����{d�0���D��!��U֬ͼ��W̞�s-�uD�OJ�V4��>�b����ķ,�D̞�,y�r)��~B�Z����b
�4�p��=ש�u�Z�pA�l����W�NJ�'NZ�~�R��,3d��1�����̤���ǟ�� 
%zRg=�TG*dGX9�5ڬ�ͭNៀ�6��h��0L�?yC:�����hQ��v>�v,+��g.�/y�Y����Kڈ�ʉx&S���T�J/�����D�7���`�/�f�S?��,���#�0d�,�-�n��c`�=�DM��0Q�v.��sӛ�CJ-�5��B}�C���)[���ڈ(@�R�n�{9̬/k��u=Z5�H�Z��'�Y�A��M\�Z%���-I�W��̱ݦ�Z�n�,�VY��I��&���	B2����	3����n҂[S#:Ā���Ȯij����c�@�:�����hʕ���`̫Ȕ�P�0cZ�+��[u�"G���>�n�:ZD~�g+mf���o����"����u+4��_�.��|DqX���no�Dyt6���� =� Ia�
�%|�x!q��=�xЕ��&7��I�1���̼���28$#�d�$�Y���	����F�v>���~06?1�ނa#�U��m`u�644_�0��#>���0'qU�d�!!r�����ks��J��N�ςQN�BV���D/X�< �yJS������;! ��Jh��y�\k���3j)��vh]�ǱE��r޻��Ů؉���v���UG�2>mQe�����>��o���/�,�Ja��~�I>iN�#�x�Pt�Iod���-g�9é׋CY������=�73oef�+�*����\�Y��*���@W�D��ū�e���*�k�7J�6�HF?���#�����WV}�}Nl���kL3i�m��?��DQ������ �df�(^;L]���	Cޣʬ���x�p6*�{�^�I$�7�sj��^�C����ɦ\�1��Xh��9�~.� �$��$�x�/�E�N@��ͻW��i 3��%����"���M1Z21;��_��E���]&��:��_5��h�(߬Z`6t�n_�l�s%V�I�RmWՋtM�}'�~�hg�8�(��l�B�g9�dۑY���F%k@%4���PoX����%�r��S'���wi�[��H\;�h������� ��_?	��hl�	�a�[v�D �</bl8�5�x�v���h�1�B)K��wvYUJ��;����Z5����w�)��8F�t�PoZ�{��'�<F�7�s�����=0k)��N
�alz��^�6�mN�y��m�b��ÍR��v�Dװ=���j�.�$ϻ��y:� +Æ_e�A�v��z[�̈c*���г�Uq3�7�H3����`�C���lv�!���^|�b�.,�+�'*����Z��&pb�Wmo@y�n�u#w}Rh��z*X���<=���J���ܥ��yw��|�x���>?�Q[���1)���z)7��x�s��cY�:\?y*�Q��el#V,����+�!B,�����F�õ~���{�n�M8k�ٴ'�+i�ٰ��}#�^<���\��F��v8�M�]�b�ʲ�)r�i���qs'�/������Ȩ�(�7�~�`=.��m��Wj8���Cm&��PxQ��ߋb'�
1�XTp�EU���z�1`�ߑ�{�~I5P]߲�F59��2h������\ҋ�"�
�Iޓ��}���:F���+��HX��(wH!���p�A����
P(`�*徠F���mqSx�����e��|_2<@�(3�u�l�m,��2��q?�v>��G�7�ۜ�m�>_0��fr��5T0��u�SG�1�L��8�d�O��!�K��,�T�H�/�W���M!��Aq�Z��!�8df\���D^rI�����v��=P��s��fF���9�ߒ@�*y4�M����v���JM�vhz$����g�ukP�-Tj��5���N�bi�Cx0�ՙ�
���Y�&�\�a�o��>0��bI�Q�x�t�ڈ��1�Y�t��"4��հڬ�@�=��ҶJ����aT��N<I-,O��Z�wr��:��.�B[dg�U@�cLqKd���Af,�f��(��GM�Bp1�qB�c�ك�Lj��Eڪtb�{=�	�~V��p?�z�0���W�a����B«H�=w��b%I��3&�(#w�h�/ʔ<R/1,�ܲ؝{t��$?X}E�0��s���iӆ� 	��pS��qa$�c���8��]|"�z��~����/��o��6q�R��%sBҸM�U����B~D�c�;y��f�wU�ب*�y���ˎ��PkW�1k�ܺ���Q���hJ�؞p�|?jjxUx����2���6��5#j\K�wEݑvZZC�˄ W�&2P�&�Y�D����V�5�n"ƭ"͒����WѰv~1!�Y�m�<|���zN1�2ﶢ�8io擶2G��Yu��#�5+�񸪾M3���4�yD�#�˷���!��@���z��3𨓸�#����D���'�
N�p@n|�e9g$��tw1b�ۚ�3.{9��+������7������h�Q@�{�u��K.���K������pe��>�
9�7�x���r�vA��_�f�a0<��b�eg�
N�h3�[ר��9�F�Γb�o�՛�md����N�.v3_4`jf�ɨ�1�I��Λ��� �oC�W�w���ulҸ��|ۨ��v�e�@:{U#�H��(U�Y�u��:�͜G$��F�O���Ѓ]���g��o�J&�kse\�}�G3O4��T����G�O�S�)�� �\WIPF�Q�a R���Gb4��)СSn�8��Az�z疲��59W���i����7q�l)�%-�s8��L�f��U�n>d��!�@I ]�45Qʢ����`�j���K�N��L����iï�����YF�Ȳ�8�h�j"���rY�|(�G�G�Ĝa���F�-�P��^	;��H�>����R;�Eľ@!i��AVC�>5L���%|��%��ڴlc�v��#nk��l+@������0u��O�X�x�^��8k�R}�D �>��||q;EG���x|&ΝS�
>ۻie��M*&����EZe�
�m��HR�5J�p�ҝ�7[i���0�@�,��RM����8$~�Aq�k:�ҳ��cT���=�,�m��^}���OL��L�!��4PO���d>M���P�J��R���ԑ6����k��ɘ"3˷�k���k�,����X��%Z����F����Th������rG��ћ��:Qw[�ԭ� �r�x�:�e~𴒇;y����:�&�T�L���R(���@A*�p����KR�q�aa��j"��̔�o�9��&V:� ���6�O]o�a �n�/sA3��5���k;�g�<h���2ө.� @*��F
H�A)�0�Y;g���Q���7L����aLV��H�+mw�����69B����!��;�����j+��!�G��w�:pǕ��!z|���XQTS�PT�����%O�\_��PCA��s��A\�n���*���#�77���D�mߩ�V0���9�ş����̓y$���ٽ��q�V��;*O7h�Z���H�,�/Q��1�h��(�C^����e��}W]��)eŰz����FB��͡X�
��
�[l}"D#Bu%�Oy��N	$Wn~�G
��To�=��l��Bed���)^dWs�\�E��h(6��	q1�lh�]~d�tu	Li�(�oխ�ܾ�.I�_w1�֎vDb/j�u�#a�pe���:������d���d$Jչ���ӏ���]LV�>���<��&�FZ�D=��Ϫx�	�L.r��SLK���+ͪ�k�@���GI��eH@�x]r� 8�\{0�S#*�=̩7��ŉt��91�7�P�70Pt���9�"ZOv��S�_q��N^:��=�
&�>8�vqH�`��v`�k��/���sZBrt���&�K{r�88��W��!��^0!ތDs���,�-�'����y|M��Ꮎ?$���ץ����"Hq�P�ھ��|&=M-m�o�x���O'aW�h�+ږ$�?u(�x�����4ɒOU�HJ'6ھ,�}�yd��t�*GqX�	�n4[Oy�ė�ƻ�ԥ�b�*���^�gV�F��ӝ�R�����x �!�7�v)asK�~���/��b��H�)��a
X�t{�I�_��2�g�u�e:"qGŻ�F��O�IЄ�B8��g;������\�+�}l �O�yT��hC���W)zGꡓ�\�~���BB3�_�fu��)1��nY�V����z�����6W��c�	��Șl'�ԊP}��4�3�ψg�U����Y-݂������Pm5�������;j�ksK+D�ݭ@=�l�ݯ\GZ�X��8ÊjCZ�ϳ��|����=����G�cm��!	\�HC#���YR����_�]i[�V$�5P��x���Б��[�sc2#���]�k�@Pl,�`�Ѣ:i�0ֶhOf�x�LxY:�k����E씽_��|�ہE�y���x������
�3ifn$�na��+�E��e
']d(MM	h+Y?�q�2Ҿ��7�5��~����N,-r�M��x"�$�`q��@�1���y��F,7o�����u=3����B���u~��K��>Ϊ��*.J�]i��5kԒQچ�OkڸG����\�.14���Ӷ�DX��%{���EY̭=�-����xLQtr(��ќ��:rx����8jrQ���~�����k�:�Tt��F�L�K��Ӝ唌]o�lc�Qc���*�ْ�lT�va�!"AXe�~�;9T$�&7�Y�P
���*O�Ãa��'���3!x���P�;��\<i}����3 �ת'�{HF����;H&��RLB��QL>rC��V�EPH�m�m8�
ڡ� 9C6���$	�|6&e%��f���j�慗 �}��p�'��N����q�SV}��[N�v�Ŕ���%Aֻ����ϑK��(��5�������h�m���V)�·6d#�&b� ����:�1���B��اV�e�;kz�h.�ȇa�\�ͺ�QfqC�I�(�x��A����}��|��U���Ք"\B����Y��
�2����}�yYB��OhN�c�WO����
фoo�{X� .�Hhd��@���eWT�K\�p������$��1�C�� �d]�	�	YmծN���J.?  1<+v�Ó�b҂6��B��f��@��[,��+ލ�x�ş��J� �k�*�]m�Q����&=�����=a�3��
u	�;�r��S��-�PG�p�:��R�~���I@�ضra�ם�a���c#�Y�J�O�&P�}n��8���( P������Z��M��P5q���^��=���&�����7��������kO@��os;)t��T&4���8�G�W&g�,!��
s�Ǎ�-?�HD�ǡfM� �?|9�J{���A��jq��3��Ɔ���gM�n�[��o��&�'B!��i��ڷ��?����ٛ�}�W4j�+U��'�P,��gy@�,���9�O:4�N�م�hƜ"@��J��K���u�F���>�R�ۤ5&�"G�����s�R��vʆ������i�cg����C`���-�a,�h.��������	��J�_z��%�<YB�_#^�Y�;��z�Ӏ��pa�7]�c*���tB��:�>Y�To���iǜ�Ǌ�$� ��5�C� &H�i%s�*�4��sB�A���.������6��W���i�x��ς;�뢺�3vC~�D)�u�jU�����'��NPKO��mC��KȚ��O�T���e_^��TP9
uf�	␡A�/�����nD]YI1��R��'s�;�M���xv L�^��7��t��[r��3�%�s��� �۶	I����S�K��O
p[˜���.��1�uHD#^��a��¨���/-w�m�""����ǒͬ�H�^�ӼC}�Op��
�ԸJ*Y<�{��E$0�^��zd�@�y������%���Y�����J�V(�Y ��1���Ǎ��<rJ�6�W_4�V��_�Pd���Z��w�@o$�zÔ�Blhen�XoC_���d�^o��c!�V��9p<�Y'�l��������F0��]_1'��e97F~!B�����������ahǫ�Ѭخ+��u( *Z�P������
�e��$I�����.�b� �.E�hy�3�l(xzMPS[߶���	��d���V6���՘�g��HC��z�W��w���ς�+'���G��$�'�ܝO�x�;�xX��=�Yb�+��y�y�)�f��E�;^.�����H��ӓ惮s\���P%m{���|��.�z�.(c@LT�_:�Έ�{)�t�{�� �*�!�G���U.�������g)7�[�-Eqy6��@���?��UQP���'�� &�Y�/I���Q��⠤5G����$t��)��<���]a�/��74o]!��1�G<�	{�ʾ�R<�&���Yrγ����q�D�g��Dp	S�NV'�{��Z]�5�C���^h���{.J��Y����U	��:
���Y���h� ,5�=r���/�#���}"��V�j8q�������e�J�E�+Wv�.�l�	����#�����{�-�J�^��x��\��U�����Vړ����:3����䔷(� q(��2kܤXE�IpM66�!��0 �_s�_B<sq�;���C�M�ٜ�KM^jLل��������/�X@K�-CK���Ҋڝ��\Q�%���f���X��}�BG�o��Iӻ"�w\P�PHd%|��V*��<;���[o������&�X����c~˳�a-*�w��K���Q�u�����E����pǱt���fY�}�Z�f���:ς٬-K@�
p�*�E���$w�df��KpgxĦ��S�'�as��gJg8a�H�-��WX�^w9��p��9��@�3R��r�IaC���� %D�9<�Rn t_�T�^���g�R��?ӛJ9s�,� +��� t%�����g�]�l�n���s��x�|A�P��<t�B��!h(��#����8/��YA"ɸ�mJ�z�ْ"b���I����r)/�ϴ�!ui���(̡�F��9Y��_�Im��K,z7����6R�(�	�Mm�кr��0�v�n�+c!���f��H�ǻ��ƚ���.g�P��n^��A�˔��3����4���#��+Ԩ��!/�`i睩��0jȱX��a�����nټ�Mm,�6Rୗ{Gr�����˴{Yr���	� �(6�V�DH���g>o4�F}�1����zY���o���2��W]Ys�g;Y�t��	k("������ꑑ�˱ ]��"��!/Sd!.��7@M�)Rd�yO�:T�_���ŘND���e+�7%�<�'�Hp���>���B�DV��!>�ֺ(�{͞-�E��l]| Ve(�+�b+u���@{��랉1����L�,ު�(x|�}��p�+�t�����C����{�oZ��l̙�2q֔^ V8=r�&�^��|�@�&a���ck�h���[�s ��t@S&Y���A�8��DW+lM���!�n�s�µ��of�m������MX�ՎD���M(��h*��=q[�h�d]��AM��`d;�n�¦''FU��g����?{���>����4��U��'�.I,�kgye�z#���7k4������Ɓq�� vv�p`�dˏ��F��B��	gR��ۉ�Wܧ'S����sQhN�ۘ῵���ű������Cy`1�-����Ds��3�����p;��z�{���ɩB8(�##�浠��z��L�e��|��H͓=�B����NjT�4z�ģ6��B�T���{�����hP� �1�i���*��&��&A/2�.s��?A�[��W��i�F���sg;C��Cc�gD��f��jۑڣ)S�'��P�H����>C��B�摕tДTm��SG^��BP�ؿu�Q��u��A�0Ϫ�i��3��L���|�E�u��%�x�=���t�a����[w�U���%A���~�{�`��I��&��K|�w�ےT�a ĩ�?��|�u��}^����_K�V��44�|"�ru�����$�@^���CB8�p�f~����A�Y��
�ź�0~p����t�O��U?��q2�}&��7S)J���������C|�K10J��.W��V�j�_���)H&�wd�k$O�Ùbl������_h��dw�����h��9�Z+�^�lWլH�?������Ƃ�%'��9�Ѹ~&b�R����K-f�{SƆS�b!��t���� �OO���Ag�LZ�e;ʩ$�X��K.��� ���E4����%�,Rzr�m[��2�H|��ibD��Ֆ��i��L˪Hȑz�A��<�
�4�,+,�3��p~�i�T�����$��X�!n���b�T!�gwy��\f�ͷE:_'.�l�fa�Q7�s���F{�Q�|a��.�c9�5^@��_?EĈf#)ݍ{x�t �C�F�Z��,U�O����7��V���-˥y���e_K���U�@��3�,#���uUnͲXϟ%������)�0�7}y2X�:d�M��0Q��<>���q?��S�g�*Xy9���k\�K?rʎ�)S��=T���x뗊���7zVX`�K9k(kS���q�i��dd��m-+�nsI�`��ۅI+R�պ]Q�銺O��Y��-����nл����.n�JZ�m �7�U2����Օkqd��i5����'RㄏY�GF���8��^��L�l��.��d/��_�En�"����&�nc,&N.��n�2����L�d���n���S�fc�b��Dx����io�z�u+@0�`�F�{J|�0���%#\����5;�ZO�ѹ���"�k:蕓Z	��g�1f8�o�^k����"�'���v�4�|����|�ʇ��|�oH��tYQn��� ��HI=r9
�p|g�!v�c�Y��`�ֶ��7t��I�Î��.Ԛ7(�#fU'$_�ʷ��(����>0�W���g#w��^�u���4����"r>HԾ0i��U��W�8�!�rB���fk�GM��!�P���G��|�RX����^7�2�0��;�R��!l����;�?�)�۱h�"c�j��r��Z�*܉��Wv7�U�0�>Rhb�|Ϸ�)6��bX|���4���Oc�ê�>Nz�#!~P�jo)������9�\��	�%�������e�Ώ�����H��^U�*�'H�=���)���J��e��]*�37�ˢ6�r?����h���TxW�D{���H�`L��Lm���?+6�D�Xu�����r�.r����L��z��H�����̦]C�g����^���) j�1{�苷��e��A�	�y?5�U��Cʃ �8ӡ�B����x&WE�����c��<8 �Ok%��͒[�G�3��Z�";{ k�����x�G��x
� jϧoԒ(G��ZEٿ�d�l�)h7㴷@ Ր�0�Ľr�\���Me�8s�ŁxXB��o��C�YWFʀ %yn��c*o�;��.��7`�S����|j[R��\�0����I	A �X(?�I�hѩ�	�@�[Թ����!lIl���5��[vO4�hW5��G=E���Y�s�� ���5�H��Һ��;e����ި����`7�'|���\��s]V<GH�=�N��O�EaQ�����WL�Ҧ�A���g]���0���Ev�վ�5��	�
.JG\��V�:���+H�Ć�Tvxr[���1�Ȱ>���qPQ��ɦHxbx��J�����f�1�HІ`��c�b>���p�v*đ$,'��ƃ�b�Y�o���n��5w"���S[K*�<�t7"<bL/����Fu:��z�wGQ�|9�n����Q�Q���m�(BP)<�P�3�%��g?�RQ�L���E�#�%Ѣ��k+u�,�s�޻j�:���,k3�F8Ы�ٹ�+Q
���L}�<~���ܳF��78&q\]����Ww)�6l��3�s��T�$��_��,��-{T�#�`�H��ϗ��)��׋�C2ۼ�g.V��0���O�r1�Ќp����"
zw�V��]��N~�D�]$��F��I�6\��$Z���$����
��S�.����,�Fo@�+[�*X=Fw����|�A�x蓯	#��|�W֤� m�WѮF��5���J^2���m�Z��ۜ[mQF2�m�?$DJ>�G�e�� uG�R�a_����ѫĀiT��ou"pG�j�L�C��Yl��mm!�N���#TG��4<��/�Œ��&|M�]!ڐ�f!	g�SrN�N�Wm��9u�����b���E�W�x�a�R҉�����h�M�������y����4-YvŚ�g:��7�bNPzC���վ���"i���S�f=�vu�0/�*b.���@bt�p�=�����^a�SY������ �@ω�ӆJܭi�~��aYMN��-q�(��w��=��� ��+[��R�Z 'c�Q�d �&����U(���G�gp��8G/]cB�.����*��t��=
x~��p�C�5#D�Ka*�=ʱ
ԫͽ]=��@'Wc*+K�������y�/���ׂ�{9��$�uEq!�	{3��i��-��7\�R��6�$&����!���R��~��n��[66���XB��g���8�64\~)2c\�̐D�-�<#T���y�/��3�^P�*�@�?�ɥv���-��*����Aj�@�0v�2�b��鈙j!�w���v_��)� ���25"����6D���~ ��g�'��6_�	�:ѕ�\��oY�j7-�=U�1�Y��0�}e��x;aGx�Y�mݞ�}�+Xa���`[3t��4��Y朽��<��1�2� @���s3�Z��>
��qx�D[.L��N���@��e>-��f��1�<m����{�MR�|�ҋn��afc�F��h�!��`ؖ�vAj���xKnA�r������O.z�OU�9�%�x6�#�@�o�;�o��?��f�o��h(e�O�Ntk��6a���)��p� ^�]Hn��?N�Fa3�s�`���Q�L��IĚm�fjL =��<�ڬ@ިu�̚��������j�: ����|ju��+u�i�:f�G�T�F��O\#3������g����9�0��\�Hw}��hO��T���,"��&<S)>���+�\��Kt��$��Jy2���W�AY)��n�KC���rz�nE�r�z& ��l0�Md6�\��[ta&f�xE3�kǈ�=�Ux���F�MF�}�5�N�I��7@j�ZKo��q���[ԯ �%���Z�m
�8��jͶ��ʈ|MPhc.��!���P��؏�,P�	 |�H�Ԙ����R ^��#�Zi���V�5Y�f��ȳ�J?X֟�Xc�_/�(3�k���lp�M��6~@	0�v�OF\xK���kY����&f�#�|��El����Ƿx�9ܝ�[
�[�i����2h)�o�^E�c
k�(������b���҂KG7�)�B[���,�M���<��$�vq����WO��I���,�?��c���9OZ��
��1�ik�>w˵4J�J:ӹ�Y�֟���;k���G������	��1�>�z�>X�n%?p��L��g��O�p{w�F_r�>���K:63������I�r������~��/������\:n� �8B8L���yR�P�w�Eix�	��Ɉ��V�����a��{"�8��B��|��C[���h�����=|*�.�F�w�@ڝ�_�-���Z)���{!�- T(��/Y��SOU���)��u<��)(�Sy���N�n��MU��4��'�&��/�yY���⮼�G������J�w�<�"]/Yk/4�4�9��w"�D�		���k<��ᩘ��A���0o�Rs+��:�	�N���ۉN*Z+���џ����ږ&Le{�-����Be���3Α����ih�5���w�������˟��d�z��$�u�ڧJ�Cy+����i�W���{���(�dJ����FG�\xV����Q�d]g��f[�m��#Dc���(��Eq���2g2ؤf�	I> A6cN+0�
�m�>_�&q5�*��B�CƱ§]`K�8BL'���)M��lOUec�/m��XNX����K��� %���N\ж�%��f���X�I�}R�����I!�0��n��%
���Q���@��7���S�.��f�o�1ĭ+c̸��/-�g7��O��CQ�㉐�*<�ө��1A�~�h�B}����}��f�py���:��	�c�*����T��ڏf���KM|�xR,ڗ���5aеǳ���8�"��ĘQs�쪳�`e1�������RG ر��Q��g��k���R�3�_��@^T��gK��j���I�,S���o�t3yr����g05l@�͹��P�F�Aa�kl��t�����V	�
���s�/qO�A��-������7��J�>�E�΀6��T�����(������	k����m��,�l�1(�6S�0(�lmM;d� F~&~�|c�E������=����h@�ϼs�P9H�|�<��͔h{R3��B���ĝϹˁ����!-��`7?�^Lzj5���N~���@ng%M���6`���I�z�����M��{g�c��K����j��6� �^x�H}��g�ΰ�TƠ1����+<����4�yyG]������������&"*eŁ����߹�0�]���"��/a	�.�	�7�m4�w��ꇊFO�8��oݛBDª�e�_�7���<�g� �&ȗ
{̃��0ZDd���`��H�O��"��;����Fq��VP�o�Z3b���`k{�`4�7C���������vkc�� ���n��èp���=�����F��?_�}O���j䶷�ùt�ƁR3��3�#�ş
����hU8��ָ�O٩ &`�R�ķp�Xd�6��m������n��������0h�\y���:��%�;
Q�E>�v�H��-gJ�y����ΝKv�ʥPMS���T�[��K��."`h�*7�/�`3P���Sۚ"�HSn����dQ-�Inʉt`1:1�`�P�̯2Q�}��6^����8-7t��w��ߖ(�EG�AV��D{ú�Z^�"�H�*k�r���5�J�*����YW�H��C������^��L��U�[9�69�nB���r�f��g&�
R���Y2� �Cؼ��nn�OS?�C��������JU�i�[`�lC�@xK�?�s�����|�@�0��L�<ZF睹w��"�Y���.�
�7Z`�+g�mmf��o�����u_"J�y���4�J�J^|�M��f�o?�et0���~ Y��I�B�
 ��|:1�!���������m��7��I����=/E#ݚN`�#]��$���ց����yh��=֮n0ү��y#n]Ũ5hiuF�\4{e���>��0�s�U�D��/ !��*��R\k!��g���j�F�z��^��s+X�a=����c �;=��Ot�����C})N��hy*۱�r����a�}���'v.�UcM�>	 ��~���������TF_K彋�P���o>��#�v�Ps}o�������9�UU�߈+��ݱb��S��e^e�1{�Xt�u��*������������a�e5+*��7�[6�p?�u\�?���P(�Wr������/Lϕm���?"�Dm�0�q,�	�Q�Y�DÔL��X�%_e�?j׽��:��a� �&�^�
��ӎVj�=���<���Ǧ�����}�4ךK; 1�z�3����ex�zE�����X�W?4%+ �B�%���RVa�
�Z��;���r����2��Y�7��fx�(��Z�����$l>�}r����է\���h}�3�"��D8
�O���B��޴ �Y�F�2&%P_b�o�ot���Ǝ�VSÜ�ғ	�[Ib�\W/\�;��2� [�?%5�h [	�]�[�Z�`s���lT��5f�v���h���^�=��ӳYq���m�����5 �O�)t>������ �l�>�_='���ӧ�s�v�~sk=$@�ŻUj�a�}�zZ��	Б�).�xj��~+��T�nwKv{����W��� .�52�"?:���"+J�]�v/��[!2׈����m�O��q,Wj�ӳ�HO�����|b �R��ވ?Fн�9�z�fb5��G�*{�È$�=�b�|�o�ARn�Qw���*R*�%�@�<�gm�f7��}Jm��w>P)|�K�{}�[Q�R��7�_^D)S������n��t�?�l�QVv�#��#�ݢ�{+lj,���r�����eݸ�^J8Vl��s�+e��b>}���<�b��F���8]b�]c�N��)��R���~sCWd˶�.�i�c�m�D���)�`Y�Ւ�K��sx�N�AC������m!G�'�V�&�'1_�p�SùT�z�6�춇���ۅ~�t]��kF�˾�͜�������͋1�K
�a6�%�ؔ�B�F&M+��X��wd��.�
A�Sm��GC|���Z����1m�=��7��l���M�2��Dc��f�3�Mm�.+2�d�?[&|>)�vG��%��?��	��_LԆ4�'�ߍT��u9_%G���L�ʌ��F��k��!"E�HFT~�D�K���&CJ�i|��/�v��!Qyfx5���
�re;7�N������I���4��0��߮%[���i�^���\����Mf�T�nhՒgLж��D-pb����/�j��bY�C��z�5 ����(��}��m�G0�Mb��/ǔ&t� �Ǽ�}�uPD�J�����,v��@�z_�_�$J3�˼��rap��Nآ�-H�0�A!w��Q�v8��J��[ T1�q��c���d�ր�(�����(>��Gi�Sp͇�^�=c9!%�h����x�t~i�=���~rep�22�L�p;{Ta�Y�h�f�d�F=+K~��`�BH��v-�����0��/MVP�NF!{��$ۜ�E"�����
{i���<�������$]���mg��3����~�������(6��:Ï"VB�H���o��i~� �c�y~�������D�y��5�*XP��]�1���?���`u��)�:Ð����j����"2<�K�̥`�wjx8nw�m�vv���� s�;2�Eߗu`�D����r[�
���>�.-�3��Ω�LѩM�YY*�iX!��tÝ1	�N����T</�/��G�Yi�?�+���ڼ�3k~K4����S6d��]���>.�2@,f��03�@{��ۅ(�D������N��@
YeU���]��1~ȭ��<{U+����pߘ�7�ث��hє�������)��K�G;��fz˘��F)��&��9`��x��T��ZƂ����W�}�ꆌje��jN+ǒ�w	�����b�����T7�d�TQϜ���N7i(3$�-`��8�^��ZI�ڛ]zF #�󫘬��#u z��]¨I�9́zd:�d�m3�u�,uK$�:�
qG��XF/u�OSA�П�4�S�g'?0g���\���}Ǘ[O��T�^3��`e�Q�)��G�<F\��1b}f��O��!$����VP�8)l?�n����[z�O��Q�V��9Y���x���W��Kv������:����U/�D�'Pݽ=+\R��15L�@[����jV�K��������W�3��u$�dR�8���j��fώ#=|Ļ���8F��3j��'��~�	�d�Hԋ�"~�RW�t�Z4i���V��50��r���n����U��-c-q�?M	kw	lG�4NG���0w6O�-{x���T�kPb��`	���[�|���E�Dφ.>�x{�*;[
�ƈi�v��lܳgrE���
��:_y`�y���j�����9�7w[��\�,(�eM�3)A$��^q:f������e3�Ⴈ,2V��zyg�0����,����P����c>i�����
J�N�ӰR<ԭφ�2�k��9���;��h1�)�4�H���qPXX��Z%�Wx� +��x���p���f7��r��uѷ$�:��@w|e�s�@r�-I�5~!M��h���:%m���n
Lo�n'b��;}�\	-������'��/{5aM�"�M$�y��9��&���0�x5OyAia�缦K<R3�_�D�;Z�<��W�$�y��\� ��kpHA
T�L��;��mm���A�LF�~/�V#|8H�wsm����\"�9^B��`��W�qa��چ��?���F�8��p9қ���A��k��ֱS�b�V���UP����AQᝀ����
��F���0 j�S���#=m�lUV�2ٷ��a�/��#���f�̸�s���ʐ�V8!;F��hit6���z�Ȼ�Q��+�A�(����|�紁�T}�R��E��N���m�BFRt�tot
D���i�}�JB�*�O��N%�zW
E��7C=
L!oЧ-:Ȩ��7d�F�EvSW��\�Ԝ������&18��� �dXլ	h�?�İ�ɝ��?}7�/1w<Kv`(��Zւ������=���dң6Y�f���GS�b����v���:O�]�\.Z�o�ؿ?&�@��n=�%8��	�K�r���Sh���%�4x���D��+V�K��@��3r����x
���#F��E������8}&�S��(҄P�딙ՃZk[!��?xq�x^�R=�&K�[���ڙ��]ޒ�
kJ�$��:s�=St�Y�&�Z��8�Q�W�`��'�!���sWw��H�����Ǆ�{7M.���8��E�ڥ��,iքq�w��Z����vMɎr�ļ���'��,��#��2B?��{�ǻ�~�4eg�U��'�E�,]�y�&z���4�J��%W4��b��[��W�쥶���z,�z0��uF5�$�9_�R�+�_�d�=� ��<sg�ɠ���K�8��'���ۨ�n`Ǯ>-���ZD����D�L�����O�z�j��W�B�$d#9�v�>zP}��M����j�2���*BN�����T�5�Z~M��oӽj�I�ۯ��P}�8� %�i`��*P�a�n��AE�2.I�Pլ���mPWӀfiWb�G��;�)��&1�C9|1DD`i����ۧ9���B'F	PFXB��Cj�xȵ���ʚMT��v)�%^/A�P4��u��K`�A.>��1*<�I����.�����j�u9��N>x����*L�ɼ�k�[�����%W�8�T[{��"�I2����4�M���V ��hɖ���uc��^..��L��,W�ʙԣh�-"��b��}�����^)Y�CXېp�lr���5���Y�����0���4Ǽ�#���nƁhQ����MG�JeW��tEM���R�!#�JU��WZ�PV�_������>�wzv[$%l��/�lc�b���_>�dM���1��9�8�����l��^�)�{�.�a	u��[�'�3�9r%�~�0��n��<@8��H�ܯ��x���=>���{ %����(Q=�����e��$$�����.D'x ㆨEJ�����+�#z�-r[�C��2����r�QY���Wt�"|�H^]�z@�d�R��
�O+�K��B����Ǘ��̓&�iaX����x%-bo1��t�Ky�f�jeEЖ�.�q�|֬�'s��sW)y�({edo|�Md. �	aB@��T_Ս_��n')0�{N�� !�͜�(����UiS2�v��bCT�����<yQ�K�k��@SU���i�'��I&D��/͇�lʉ���G�ϸ�_阓��+<�H]��p/a&�4�O�,g��"!c	�k��Y?S<����64��n�߭��Q��d����	M��N��vɽZ������\�&���u�{	����L$Ǐ�#��Kp�$!��ϼ�hϳ!5T�^�^B
��Z�Q����T�Q�����J��+��.�i\7��F��AJ�H�Uo���Jg��Sչ\%���6?��QL�h3u��G��g"�_�5(��\qc��2�t�S��I�)�6�������ڵ+_Ϊq�0�3�)C��4��KQ�L�ΰ��$��y���/���X;���B�K�
�����4\�8G%�zf+0�X��M}ߟ��*�5I��c����+�m%��T���ץ+�<5������"��|���Z��c����-����Cj�?Q/���Bـ�u�~q.k(�ς#�!Z}�;ff���c���<	�6)�:*!OS��Y����f
1KZ��x��i�T��"��a]�}�"
^8|�_A�ĥA�����έ�����H�&TRt ��d�6���۹�tlmR	X_�D^�EJgH(i�7��N̓�, <��k�?t ���g]�Hl�X��;�S�/A����Ut�<Dߴ#���j�a��/~3�A]]���uJג}m6kC��+��:������\�|�^ь(z#�ɡ��Z�zwm* ,�e���GZ6���(�+KM� ��-@�K��fc�#@��p���kǶn������~HP�`��P����U�3.̥�/x5����泳�Í"!�l:`D�����jcAg���z�(��n��M�E6�h��V�r�BA���:{T�Y�I��Įф7�6A�7k�,H*��g��l�A��1V���5���G�e���E�]���o��d�"W�d���r���ˌ��]?b".p/N7.zQ�7��O�D�L���O�~���w�`? D�Q�ez�7���<���G�ȤHy��}T%DQ[��|"_�u�	��{��������QoV��Q�;Tb��Q�;X�-
h�ǔ��&�g����_��x~ܙz�t��p5p���=j����Ź���n����q/2��C>�g�|R���3���L㭊�b�U~�n���|@= ��Rp�η}m�d�CS�1���8�Va_�Iw���O��0u�hyVg]:��(�QAI>Ǘ|e��-gWIy]�
��`Kc\=�2�^SǉT��8���;?��78` |](Sv_��F�,=�d'�<-O©ni�`c��û��g�Q�;����:���-�=��TF������j,n돈���[�w�7n��X�kL���;5���#�L���Yĕ���"{ᣟ���qp�۹u�D�����nPn�T4�G�ᒮ�&��I���K2O�9�p9M�j��n���SLAҀ2����h�7/Pis^��LX@�<Z��g��ݕT�d�ɚ�k&��+�Zs�7�DP�"g޾_���Z���g��Xf���o�G��W"��v��}L4�W�ӗ%c|����_5folXXt��[�I� f>YIa1W
m�E|'(!�0�
�a6f��(7�pI8;��D��2v�ۨ�#��8$��^��%]��@�迀#m�0�72ч��#��ި��u�K�4���ɍ�>�0���U6��\U![tm��%�k.B?��R·>��<���vנ�X���Q����4���;�������̓�%�8���K)�ٌh�坱��0	[�f�7�3 ��MT��C).N��.:�s��bk����Z ������ߺ2�`��I�>=��B�� C)݋쌨����o)���O1��pKY��hRzn��V�ϑ7q�~��9]�c�FB���m�;�]���Ѩ�
i��Ū
�Z`hF��+���X3��w���r�A�)d�F�W���`X��T�m���=�e��Iţ�~2x=���:��i��֑mh(�2y��?�n>�ۤG,{ȗ=���g�_�������Tlj)u�_G!'mLMh
�R��wF!�~���cT������L��	���}!���!��4fC����r1h��wD���ۮ韁�"����d3�N�fc��	-{�WE�ZM�M�6��2��p��	�-�e�q���
�,b�*�C4܄���K��q��b�s��b�u�0�smb�_G�4�+t)zg��̼�15�������CZ��Q@<� ����J�
ռUܡa��NxlT-��W)�'w.�.��0��qC[��w�^�c�F�dwt}z��"'](�1�G	BDpm���3 c�*2��o��j2t��=(�}~9p{���~�$!a����O���=���� :���݇_�Y�$)����
/�[��_�{02;${�wE��s$��;$iI�q�ܔ"�VK�-��$�%�ɤB����6E4~D�߶���%�6-8��/dJB��ˑ�z̭��~�Bc��|�[�گ3������yb���!P'��m��v%����$�s��D�8=�j�
ɧ5�2��E�� )>j��w��6vT~ � �2�7��QD$oH�(̌�P'���͕}���(��b�Y�X��΢�%(1�$%+�������G�U�Y�����5�+/Ǫz�3h�4TƉ����sc��H�Y��@̵��6̾3,�ø�l5��)�D?7DcE�N�N�@��Ge�L3��c1&;�v{�p@�z҂;��8��޺�p�Q�dhq���W������GCKe"�I�:kN������L�9 Pxm`��W���2|���y�
g�,te#�RN˸��/��&�S����$י,�����j�]N��?3Ĳ7`�1��:�#��I{�����l �����w�wd�u�춙�w�镘�!��:��ߙQ��G��Mu��5:]��G`*�F�JJO��i�?��S�Gg��8߉�'��\Yi}g�Op1�T}�ݡ�r[�]�?)U���0&\�������!z�6����,)��n�W��}pYz�T�N~�UH�*�~��MH�s$�R��뗹�/��?���"�UϞ� M��]��_F��=5����[uNj�F�K��d݈N ��|"��78�S���,8~y�j^ �.�_|d�ZVg��G(�ӟ9�i�����	w6�H��	��7R������iV_�VpF5�T��8�a֖�~c�T���kE�l�D��X��ӳ0�p�O=[�x"��Tjk�+8� 6�z�|8��E��<���x��-����
z0ji!&҉�����E���
bh���RH���k�,���7���Y�L���[,�O�M�����$:�4q�����ǀ���o��0t,ҷ%�վ�=�NV�]���_��&��>	��ˌ��J����P<\�M#�!�kU��^�w��V���OE�����XOy%��@���ϭ��O��G�Gr��t�W��:���׭|�r�[cv�~�6��w2�K�t:�<�oT�L�����'��������X�@(S٭V~� �a�@u"|�%��9OB&���=�o�'AOgna\�f��I73��沨92;��O<$�J��,��e"� |�Pb�H�k���D(;�Y\��ߍ!s�L���ISV���HGy�m3�����9�_� ������y	�&�0�]���G��7pُi� �8����0ZS���/������yz���A��ʀ%�ɪ�Y��͡����ߎ�ݘm�j*VD�M����w�>�~�[b5���j.
V�r{;�*�h	�퇜C�h�Qa���J�(<�E��˴!¶}�,e�����Տc�B��.�M�
���G/o}^��B1؊O��N�o�W�������
�R�opg�����`d6HU��W��\���l8�ջ1د���d�v7	��d:��i[����y�'�1��v ��k�8�1�����!�ݾ[v��֞C��}�Fu�`Dl�E-�Mΐ�L�]�`����xY�&x�7�`=\�Y�?m[	��>r7C�SC�+_Ϫ����|��y�#���i@F�r'�z�3Ʉ���#�"���큿ڿ�&^��^�cMP0�o�u�;Z	�̏�pq�0}^vh�=�K�&���2!q�����2��k����M�s�'�tGw7&O�Q7�8t�WaNF��@�!���s� ���|��c@ǄB!%M�o��zƕ��z���	 �q��������8��Mi�$���k2���'����$!��Ҽ0?1�@�`��K?4��U�f�'r��,��*y[xP�0X���V��q/4�!Iـ�e���Vۘ�fl��V���F����� �Rz!��E��bJ��5�sI�Q���nx�r\�^#��H�`g,�-��'���������^O褳fE�5zBT�����B.�#�@��nz�j<�[2����Os�OB�m��0TJn���؜����
A��{١��e��^JH �j�i �*����A��.�#u��Q�Wsf�i������;9�e���C��D����1T�G�����'�v�P�ye�C
���U�B�j�hT#�����^�NGPԟ\ua����	�A��ѻ~��^4g\⺪��r(��6��O��x1�ʪy\V�H�O�)[�����%����D��@�I�y�������ǒ������=?�J�uY^����;��̰Mj'��;G"�p��"��Z�%^�jC� �p\f�Pa���WY7'_�;�o0��X���/�����nk��!6 �sqR����J�~����9�i�u��\\J�Q�W���V�j=_Q���_�u0�w�1$�E+���	lS�Sm_ޑ:d�*�������Q{9K����X:lM������<��L�x��'t�-9?~\~�Hp⊯M��)FA��|����؉�g�*�� ňJ�K���>O��w/e1��$�(��gG.�< ���E�5в����zh?P[Z�`�+��� ;��:a��m���E�H�Z�z�1����Ȍ�O�+b(��k�E7�7`K�3į	qnX�f��_�b�����y�W f]t�Ep�u.����ߡ��
�,bs��m�K�{�|�+.���&�@'"|_u;v�\�)�8�{�Ɉ �d��<#��<_�U	m��k��EحVB����y��3�[=�úE�U,t�V�'YT&�%/�V���� �G;u��B/�dw�<2�]\-l/P4*����x{��f`	VeC��l�<L����I��)�N�Ԗ_1G�4�5	�wN���K�ZX�_��%�]��3ǰ{�
¨4���/!p�cmJ��v��o��ho�+5�Ep�$����������3¾��.]��xJ�8k+��ڽ	�[�D�Ώ0�s���]�����4�J=��:!\ſ�֌\��M��iV�:O���'��]�(c�qe�2Tb���#�Ik��60��M|�z'�_�siq�bö�(C�0���lK�z�L�,}�66N�Z��~/Z�X��D�(X�Ka��Ѝ�6����\}�%dWf��AXQ.�}UK��+|I�yw���<��`�%W���>y��w�B�܊���y C������eUc��w!WM-%� ��?g�Q���s�K� ���z��oV��L�}[�>f�ǵ�uهVZ�����;*���!C�:)f�uK��x�z����O��'a�|g��8i���@�E�̍9�?�MG� �U�;�	RJ�a�֧�{���fR���_/a�^�[kg���׋S�}����,����^�t�E���Z5g�'l�����@���+�A�ЙYC�t�%��4�����Į�|]/YA��놨�b��cZ�|Q�"΍̫�J���J���~z(���A�������m�=�,~˸�~a�6@�(`-�Mh6D��)�5De]��(?��]?-_͚�h?��T�bo�C>-�����f�,�'~�W�00bOlf�>S,ts�|H䎼��A�a|�4�3��߫���@F�#�I�sJ]E��h�aɵN�5-r?M�S�w8/>�`�/�t�[j����cҖ�d�$G��,#((�JG�Pp7�S�c#%��&׵K�t(�;=r��~�KpE�ؕ�#�%��a+����-��E'=�];�z��T�i�q��@�ʚ�./�� �8��{���$E��E��n��4=ai
O�� ���c@��?U$ǭ(ɮ�6��_Օ�0�~o����)��܊6������B�������7�l~J�/c���9E��Bbخ��yl3���P�wN7��܀�˥� �)ؤJx�B�yj���1��2��O�¥J�Ej��wK� v }�jG4 ���2V<��$Dn�-�p]�t���U�5�
*�Ѷ����RYb|��ި\1�!�u~��~!��wG�ǫY�5P�iRO+�����Yn3U�4�潊��}?���UX�@����@�`3v���?�����JDI}�LaN1?�@t�&e����G�	1�K����4{� ��I�y��a�Ē��h��ꚁXj��ŭ��,K��6�>�u]��0�/�PF9�6�xw�C������*r�e��'�:�vQe���N�կ!�p8���M�h;��|E�>?˜�;N�y�3�
�`��fb����;I�굛G�� >Xm�]�ެ�&%u���#����Z�+g�:s�������u5�5:�N�G*R�F�k�O=�����g�b;)�m��ڟ\#Wq}q��O�cT2��M�k�g�T)����f[{\]?�R��i�K�� ћ�M)V�nl|�G�z��H�O5{�����!�Ƚy��܅o�g6�9������'zU�C�*��ݧ��HVc�J5�9��*�
��j�K�*������1O���[_�]���Nګ8�/j(K�8��|�(@��Ģ���ݦn���n�-�F	AY�H�U�5�R�3���i`�V�}5Z0��a�B�Ñ��n� L>c�����ka�,lq
��ϑ�#�0��O��\x��^��k:N����D��|BKE���Xp4x���ԟ�
���i��L�S�����E��?
�+ɺhR��������ң�q7!�����"k,���M�(a��$���q�ư�����ج�SP,�+��$�C�����^4�'`����j�px�>���V|8J�۽ӚtO��dF��v>k_�����!M8����f#�[��X٤+%`ff����b��/����Q9Fr͉��ᗺ:W��!bc�]�r&W@~�˹��h����:��y^�L	T�똩R��~��F���I����wqi�ta76�"Z��89Y�2&�<NǬ���k�O#E�a�`��u��3�GF���;D��<�N���oj� �޲싄H�/�   6   Ĵ���	��Z�w�J�$ʜ�cd�<��k٥���qe�H�4͔6Z"<�$�ic�6�'���Hξ���EC$7In	�M�ƿi�����B�;�4A(*L� �X����&(���:]���[W�i��qK�H�r���r���,�b�	�O]�-�M�������ɘg�)���@�W�4�Z�Eȡ ��A�w�Q$h��I��?a���E����<�E���?�}�R�K#0�H�Y��H~�#CE3��[7t��4�ɅML�$B9�$ uE�^ 9k�!\�'� �Dx�.�[�?lNM��CI�~��4I5Ɓ%O���	��`a���$,7<%r��>*���իA�i��m����<�OX�y�O�a��-�[ܾ����H���>���$�P�B���ڠq�\(#jE�]�p$;$�qӮP��$̕�O �A�"��tk����H�[�9�-xq�O�y��$�����\�rP�	F���4�����HP��
J���X����W�$�Gb��r�>pJ%A��8V�0���؊�O���1&�����k�L�c��;"�	�<Adn(�v�2O��1�J�)IZE��F�6=��5�O�I���S��(O�XBĂ~�v�!Q(��J����'�D �'~8��Ƿ��O�d�z�B��[i�w`��4-�->xU�� uy���9s��!M>	Ӥ��;s&�$�a�+�^�D�Nʽ)�� $)�'SDX<�Uk7���'0�$ ��$�5�$�� ���8�iȏy����t�)D�P��	   ���   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  ���	��pY 6�ky�o�M!6�������2��:Ĝ(Q��j��֞�j�����?���?a��|*)O��n<;T\�	_y��s0�.7�^���K6X�fx����Mˍ�Ρ>)����d��c=��8G㔣J>y;UD<��@�|Ӗ�1�xH�@����xO~
�;3)��T�DW�@� W�"(���?����?����?)����O� ��������s�ߝB�>x��X��	��M�p�\�|��ڛf�|�B��af�ɃI��<����te"+�'�r��4"׃��f���P�%Ü,Z�;�g�)�������%>�����OޓO����'��IDK�Vܪ�j�./�����Ԧ!ZQlyB�'&�S w₴�������P샇&Nv�w-�����K�)�š�&��E���{���'�]�m������M�[���+UA��>��
Q@��s���� Ȣ���R����O��$�O���ɧ<)�i?� bBŁF�L�bs�̭9�
d2���""剫�Mk��¬>y��e�Q�,>b%6K�N��+
�!X��?��N��M��O�n>h'8�	����� %0��F"6jls�k� p�戛D?Ol��?���?���?�����	H:'����abY��� H���\o�83N$�'��Ɏ٦�ݪ1�B)��� �n�j���"\�-��ڟ�$�b>e��PȦ��	����QE�/"�  3��ߒE�r�ΓU���«�O�-QL>�*O��O>X#C��9��a@�!Jܵ�L�OT�D�O8�d�<�$�ir�D���'��'�t[�����Eϑ/m�dS`}�'{R�|R���=���r��?v ����G#i�h�fnl�4c>�B�O��$���`ؘsIJwG�}ISC��q���d�O����O(�D �缓U�F>T@9�T��G���q,�?i��i�:]��'4ba�N��.��:@��0MvD�@u\��p�	ɟ��ȟ� bC���'"P�  �o�.\@l`�rğm׺�jd��	�����O6���O����O�����w�ӏ0�-Q�o��U8�V�N~���'���'$�aA�C)UB��$ ����j�>���?yL>�|�)V�*n��Ej�r��˒$�(08jشl��	�$�صH��O|�O^ʓ	���������V��QC=�<����?���?���|�/OZ�n6r�X��/|N��R#�P��}��2M*��I��MC�G�>����?���"PF�����
m�r����O�ִ�A�nN��M��OX�P'J���$���w�P��B�ّrY"�b�K�x^Nq�'EB�'�2�'���'u�*�k�+�-<�`C#��j3��R�.�O����O�1m��J���S՟ث�4��pq��"&���k��3��ڇ1��1O>1���?�'s��
�4����*�B�Җ9���CB�!IDX�G�1,�&�$Ͻ�����O���O��䆷dD<|$aV2(O"�z���2|�"�$�O$�G��V矴"-r�'�[>!u��+�8���
5a) �k�f)?Q�S�����%��'g+�E�d�+%�؜:�Q�_�q`�"P4xܪ��c����4��y��6�L�O�,�ǣ�5<̰�a͞�I.Q�"A�O��D�O*��O1��˓;����OPa"çػv��`0]+NiȠT�Сڴ��'���?!��K��L0��˖6�:��?Y�+7N�ش��D�83�@��O剞:�(1�wj�9n���k�[�1\��ICyR�'���'6"�'�Z>9���J�=s�1�J�����aJ#K�7-�>ܜ���O.��0�9O>ymz�Պ .���q��3�PH���\͟��	[�)��6 ���m��<���L
/���GC:W?�T��(��<��+�t{>�dM�����4�H��F�`c �IcO��U�q!AG�F���O>���O4�CK���L�x���'/Rb�I7�riT��Jػ4�O"�O��'w�'��'�R5��*O�ZIډ�p�C�7B�A:�O���ნ_�6Sw�S�9���O�L8�@��4Uz�H���*hE�@S��OV�d�O����O��}�;V�y����}NL�R�C]6.}�f��6ݢX���'(�7�8�i��� F3|��+!���z��d#�bu���Iҟ��	�@!o�S~r�^�!֊��S ˼�HcF4���WJ
�mY��|bZ��S֟��I�d�	���PI�[�D!�3�����'�^My��hӜ]y���Ol���O���h����2�*eZ�n4n|P2m;1R��'�r�'ɧ�O���]x4J&�3BA�(�@��R�ތX°i��I$J�s�Of�O�� �Qig?<敁�nX�D�����?A��?Y��|�.OvEo�v�z��7}PN�������p�a��s�6x�I��M{���>���?���, 丰���\�a����rN��yG���M��O�9Y2�J ������ww�Y�P�O�������nɆ�h�'�2�'C��'Yr�'��b�!lK/Fl�pAU�����q���O��$�O�qlZ�j ��ן$�ڴ���n�KlA v5�6gV[� ��O>���?�']q ��4���ߪ{���X�oN=e�ޤ[��SRJ���ۍ�~b�|�]�������	��TQ �J�?j<�튗S���孞ǟ\�Ipyb�p���zq��O��D�Oxʧ����.)Q򰼰���"q�'&���?�����S��F��L�XH�P�?�Dy�f�*:l�x˴�Ƚ,� -�O�)H��?	�/�Ă��r�AT�x���*ABm^���O6�$�O(��ɨ<9��i���F���?@]{��w-}C���)րA��ϟ؊ݴ��'2x��?� n@q*d�����1�2jW��򤏙Pr6�??����[���Ӡ��	h��Qc��_�`A�����'A�I�P�I� �	ʟ��	b�t�?@��
�![:<�T�Δ�g��6�Z�^@4�D�O���8���M�;c�޹#�W�:�V9��	�*c��2��?�K>�|R����M�'"4��ʇb�@J��Ț�&y;�'�|0� ��埄���|bW����ϟXXBl��Z"n�d		&���96�^՟���ߟ��	MyBiqӬ�j���Od��OL�`���#Y��0��19���4$�I�����O�D1��=A�Q���;$��\x��K
Y��?wTA�'������$?�W�'����I
0�ԡ�	+�C�`�,%p�*�O����O���O`�}B�S������B�C��"
ݠ-���R��B ���_1@!剈�M��w��1H�&��r��6eبb䈈��'*r�'Q�iۛf��@6��"��� ��R�J`xrE�F�{�N��b""�Ħ<���?��?���?Y�䊯s�`l�����"��	���$@ĦU`&���l�����$?�I�,��y���� Y��V*Pfby�Ձ�>����?K>�|�f�RL8� �*��y6�8(���U|���o~r�	2E$�����_c�'!� 8�����E�"��z���9,BF5�I�������P�i>��'Ң7͉�5��>�@����;q:�˔�R�����&���ɪ����Ox�G�hv�8&|
��q�1UhV��@�R�M��'t�M�>0���p�	�?��]�����X�4��*�� �@��������矔�I՟<�IY�'9����(ٛk@�䘣@�>>��x1��?��#4��,���d�'S�6M(�D�7�&lCF�;Uz�aR`�2C��Oz�d�O�)S�P�P7M%?�;2����	�!o�� �ʞ.U��2��+�?�V�8��<!��!R$~d�	���=�����LJ)�O�m�LK��'�\>�X ���.���b��κZuVD��h??�X�D��۟�$��'z�~��󋆇5b�t��-nd��W�-��x�41��i>M�&�O��O��cÁ��y�R]r1d�/a�����O\��O ��O1�f�"ś�-փ>�@�#E�,��1lQ94P��3P��b�4��''���?) ��~s��U�πE10��.@���䅦1r�7*?�7'�\����Ë��� 0KJp8�)L�]�rh��  Y��<����?9��?����?�*��ER,H���ӮB�t�̛5�˦�H���X�	؟ �B��y�l 7<�T�k�<g�<LJR�ʼmH"�'�ɧ�O�(s��i���^�}O�}a3'��9��#Q�QX���s����'��'}�I� �	�C�@Q#��Žu�VH�h�0'3���������ϟL�'�t7-֐g�z���O���K�@�Y9v/ 5>��lF�-d�⟸ЭOl�$�OʒOT0���(!�,ys�L7g*ୋc��\�۸,G�HZ�'?�;,C'�ʟ�[��V>~��cE&(K�e r�=D�<&j�=\��irC���u����П8��4Ee�/O�5o�q�Ӽ�s��t9���5�ʆ6��l�`���<I��?y��Z]
��ش���9��O?�8�!(H�K& �9@��R�Mh�Ǝ%�f 9���5o�Ɂ�O҃@�����e}���Z*�0rfjG�&Ci�6H��c�'����L͕Ex���T̋E��T�`F7�tp���^�
=�
]x@� �N �JU.Ӵ_��!Q�?.��@���J�Z�[4e�q&3)��I�&��A�)�k���2ፖ)(����N�)0� %� )13#��U=��KUi�	$�	4%�*�����4��uc��{%i!%Q?7���[@B|�>�$�O��$��؅�'$�� B�;^�eqd�Ȅ�r�l�B��O6`�!9��Pܧ7$�*�/�>4��".s�<Xm��)�%�ߴ�?����?��`��	ly2�W�j�B�G]���7�S�zB|6����(��1��ܟ�5Z
wF��"�A�\^��t�1�M���?!��
vr�T���'���O��AEA��C �a%�O�~Y�����D B��O8���O��$(�\�q֍Fj}��	ԄL0�|o�˟� �O��d�<)����#C�Y ��d��(ͭ%�*\��e�_}Rn3_h�'�R�'UBQ�x�t�[/	��]�p/��Pm���sFH�K��Չ�O���?�J>1���?!TF��ܨ&,��"݊ ��:Q�M�H>	���?����$P?b�`�'6�4���.�G�D����G�j�,l�Gy2�'�'�"�'�]��O�m�3%K-�J}���i��yz�_�����h��Sy���#/��'�?�3�7�؊�aհG�BM���N����'��'���'Re���d(3-ʔ96�Բ�|5�J��g����'�BR��i*�#��	�O@�����S� il�q�M�l1(�:�Fs�	۟T��E޶`�?I�OJh=�p�f�� 	�aN��T��4�����}n��(�Iş�����ƚU�Q@��h��4��>n3�З�i7��'��ڶ��2�S�MO��ʒ��n��XR�G�,7�NX��m�쟄������/����<�s��6�|hX1`NS��1e`K�t���
G�-�O��?e�I�v�%�dN�}~����2{����4�?����?��(
6�	|y��'	��]#�x���E�T���S�_?�OH�7�d�OF���O>�BPK͎K��{�5T��/CҦ��ɥ
E Y�O8��?YJ>�1*��a@�
�E1����,�6�<��'I(q�y��'��'�剗z�25ٰ��!���qmѤI"�`�S!���<9����?1�mh��6 ^�6�F홣B�zzL�i.��'�_���I�����.6R����3q@����o�̟��Ix���?/O����iL�9G���+�j�82W�
f��RN<A������Ol	�Fk�|�$�%�7�N4@�#2Z�d�i��O&��<��,�\≤��c����i3-�._>7�O���?9�L����)�<���`N�c�B}�E�ԝ@���4 �e��|�'�t����$����� �H�ۑD�rZ �p_��� ʚI��՟��ԟ���tyZw!*�#EM��j�V���@K<%�=��4�?Y)O�RW�)�i��3��� q��V<�u.�63؛��!:>���O@��ON�ɣ<�Of�� J�颈�;L�^a1U�/�X[4]��i �4�Ş�?�_�R����KM�)�%�2K٥���'��'��i�m6�4���D��0e#�
Vt�2�ѹA����ԇi�6�d!�d
S��'a��'r#[�<;�
�s�5s�E�s��6��O��`g��b�i>��Iӟ`�'�H�m݆45��̘S7�+f,~Ӹ��?�(O�i�O˓�?1�[`�2hK�l��)=�{sGM�C���	.O��$�O�����q?�+�6R�L$���Ft��ՄEզy!��'?���?y�����[�WL�Yͧ��(�f↑\Ŗ�wǘ)��5�'4��'�R_����B���'a�0#�U�}Fb[�g6-�Y���>!��?1*O����e���'�?���B�q�����gY�p
�`fJY"�&���OF�e��q'�T)�'
`�zXXEiH��2�&J~Ӕ�$�O*˓9�Ɛ�$U?u�I����Ӛ(�lx�*2�G�n�0c�l_(��$�O ���O���v1O�D�<�Op���ˎ�Ъc��
�	��8�ڴ��B.4W�Al�ß���ϟp�S�����h1p��Q�fU��.�+{rr�H²i2�'��i�'H�'uq������U��.0Z2���iPv�p��`���D�O����N�'*�I.w�x�R���<K�@�r��K�'缅C�4N/��ϓ�?�,O^�?a�	:ELNY���?~�&�a��]'f�HX�4�?���?���Vu���yB�'��Ā�p��i�RG������!�!w֛�^���I�Z=F�)J���?��p�j�{�lF�P!����
I�Dd覻i�B��m6����O�ʓ�?�1�x�brON�|�8�a��ӼA��,�'���'��I�p�Iӟd�'T�]@��q��2�FE.?v�5ʕ�D8 LL등��O���?����?項P3V�B6��1D�2o٠ɉ�'|�(�'�B�'��\�Y�.�&��d`�Rx\����-���qD؆�M{(O"�Ģ<q���?���vG��Γ��)���4mn<I;.('lQ���iT2�'���'5剌��=��z����pa��3
:5�Sl�RrA��iORW������8�	�<(^����(<�qf�5���I;��|oԟ\��cybK�`���'�?I��"��1�p�6�H"ݔ1�T��?��I���	柄��&:*O��ӟ���h!�M+\��IϳiH7��<ѷ�Y�y���'�2�'r��L�>��FnX�sV��H�U�v�@�ĉnZ˟��I����	x��aܧy�$���
0P�<�:�k�(nڐ_����4�?Y��?Y�'���hy�J��_ƞb�.�A61��CE�6�L�R ��OT˓��O|b�7j���I�)!1$.�c�'��|�6m�O*���O�1a���R}�Y�L��?y�� 9��`�I"3�`�!�N Φ1�'R�G$�yʟ����O��� �QWzBP#V�e�е V�$� oϟ��4����ĭ<������OkO�nBf�Z���&ukv�A��(C��I�����˟�	�����蟸�'5.t���:*RF� ��H�t� 1��lv듄�D�O��?9���?�A���t#�	(�! �d��[~^��4O����O����OB�$�<ᥪ�c~�iB�6�"����F�^��p0E@j!�if�	��Ԗ'g��'��)޺�y�В-�.�s�8	��x�'Z�>��7��O�$�Oh�$�<���ڄ	��S����v=XD��M�dJ��p-�,-}6��O���?����?Y��Sm��OV�2���pL`��&�ģȃ�ii2�'��I�-��������O�I�d#�Bw#Y���d ��N�x��'���'�����O~�S0f�-b�D�����
�Q��ig�+^Jn�K�4�?y��?1��	
�i��P�0K��0�[�M�J��x���D�O�H >O��<��T�	�n@x ��1EĜb�͔��M��K�b�f�'���'6���>9-O�V��,�E"�<}ָi��Ǯ<Z7m�?��$�O:˓��O2�?!�>:��Q�AlJ+]�� VGs�*�d�O���'�e�'��	�x�hXtРg%���~}!#�\�w���mZϟ��'\𹟧���OD���Ov�8v�|���;ׂ�U|8x��ߦ���^�X���O���?y)O������x���.P��,��RE
�V��:2i}��'���'�b�?�a�"_�z��(^�R0V˗2��%&������'������첵� j�@���/O)��T�����%���	Xy�'#��'a����!ͧLBD�
0�� �B!I1dգk}Đ%� ��n�Iϟ�I�At��	(Q����6h�*�,��q�	�|lЪO\�D�O��D�<Y���%F7�O`�!���,�DB*�0�~1��#}����'���O��D��#�B�d9}b���YШ�"��Pxj�Ȗ�־�M����?9.O�1��Cl�Οx�s�:A]�y�X�����T0��KWS�	韬�ɵo֨���k��n�3�?��&"33V���(�Φ�'����|����O}B�O���;��Q'#X�m�Ԩ�"h�5!i��o��� �I�e�V��t��Z�'U"�a��Ś�(�!{e�-}A�m��n5�D�޴�?���?Q��tޱO�aX�/_+H��ٷ�ғ'��(� g�ͦ!�D�ߟX&���2�`u�� C���Xb�bŒ�o-JTX��i"�'(�]
��OZ���O�I8�|Y8֌���D����.��6�<�$��1Υ%>	�	֟���8_@^�rBe  l�lx*�!MY����۴�?Q��3&�O���.���� ��RB��_g�,����H�l��P�8�����(�'T�'��P�H�c�Τ�*0iR�>��ბ��8&w�A�}"�'z�'�2�'\��g@�SP��FAM �.��a�<NW2U���Iޟ��Ty�N���j��+������m:2��	,���?������?��Z�,q��j��i&���|,��4�'C`VK}��'�b�'u�I�8���O|b&��=(�Բ�_�\	d�Â-@���'g�'[��'�D0P��'��]1T�ӣA�B�XI"g�
�`�4nZş��Iky��>�������t�Cq�s��y�2ϖ%^[V�r���v��ퟨ�	��l��?9�O��Y�p&J&
��[�N[5H�R��ٴ��DV�NLn2����O4��d~�W�I���3�1^YYT⒲�M����?)�F��?AN>)��t�A9sf�u�Aj?2�=�%��Ml�7C>�v�'�B�'���'�$�Oƙ{���.*+��HS�u�l�U��צ99�d�d$�P���Rа�$�r:����eݫH��dPQ�i,R�'�lO,��O��I�=�@����-:_�@bD�ՠ(kF6�6��E�?�����,Pӎ4I-<P0@�j���K)�!�۴�?���.N�����I�q/���ֈ*[������8��6ͥ<a�����&��9���DV�pE��Q�
�J$�UkO�J�B�/0)��Z�Z��@�&�L4z���>��BS2<������ζm��x#g�M:	B�w�2���9���9�k�?;@0F�ƛE;��x��)�����[��l�w��(8�1l�!8��r�n?dP	����7fv����X&Mޞ!#����p����F̿Bh����a�)
N�u��͖(T6��WA�<{�B��Cٵ }�IR�Ib��`�c+V�����8��
.P��]�zA�~6՟T��V�#?" �;5��
a4,����^.� �U
:/o�(26��;34��ň�_��m�5d�O#��AV�M)M1�Z����^�v��IП���A0�&����]�\���q���<1�Y�Q�I�4l��j�J�$����ē/Z�Q��N����T~
L�͓:1~i��S�x��O�TIʹU�R�'g��Akna8�J��7����o��l�' �����1�R@}*�^c>�$��-��FN�#S��8�b��{&�(��(N:;�!�����O !#D*��wOp��d�D
�U�� гC�,�D�O��S�SY�	�0#lPKԭ�_pD��"L�C�	Jݤ�eNW:G H����� P|#<���)��Z�V�2(*����jM��`�%�?��6���4�G�?����?��W�n�O��]���CeFl��5����/4����c�]���*/����՟ўD��J��r��J�!��X�C}?��&�<�`L� ̊��?�=���/��b��\%�$M����O?��`ß��Iz�'���3N�����6]"e����
Ru0B�	�&Dր��e^�}��h�*��lG�����?E�?Y�LIQ��d�fe����ƕ�<c.��'U@\�F������C�<�Ì��	a}"��~e�%�e�y�<q��T�$��c��M��� �$�Z�<i�@�<Dp��L
J�Ը8@b�K�<�/EcZ�+We�U�*�Ƞ��p�<y!@2GT�s��	|=������o�<Y�.�."@���C%���o�V�<�p �m8����º/qT	0чBR�<�J�<�b�{%��`�ٻvt�<!�ώ�ny1@U�R�v�[P@n�<��l��P�.�A� �T-C$�Fh�<A�uWtIS�J>	2VC��Yk�<�Ԃ�lȓG�:C��{5�R^�<��Nޞg����g�~�(%�4�]�<��Γi�y�n/��=k�bp�<�NX}�T��֍�+JOx���lw�<��ϵ#6����mѩL��� %�i�<�`����C���p�
"&PQ�<�3�B)=~��RP�#V���'�EG�<��,r��|�4��
z��b��E�<�BD�.GD�-��B�r�t��!�A�<ѷm�� �A��;TӂL��JJF�<����E"-B�N�}D��sG�@�<���*C�)z��E�6B�(Ea�y�<�!̕)����܅d*�S�I^�<I�A��^���h/��>��h���o�<� ��A!�)KE������$T� �"Or,��H��������/C�P`"O0tY�C15���V�˺��	S"O������?ox�;T�P�P!�u��"O.E���p��t@��h��i4"O�Ó���3�$�D��W��#V"ODA[�=F�<���N �K"Ox����.���-ӳ&�LXPf"O�h+᪂c�e'+�>vô� "O��
�^%� �Jv	\�t�"�"O�	���[�42�gF�Ĥ�1"O*q��M�;*�^]j��H2���a�"ORA�Hf�u�XQv�K�"O���A���I����fAP� �"OD�AA�M�`%�3�"*�����"O�e#	�n���۳�)cy��"O����E��F4��:,��"Ob�SCԤ�z���/�?2�����"O|�����?Ɉ11Td@��Y�"O���%�[��|a�D=X� ��"O~�ɇhۙ,+~��c�	5��"O$��V=��q�/K&y��� "O�؃#�W#r��	�UK��
	��"OX4q&�M>V�@M�F*�=2�.X3R"O�!vK8F:L(�IG�sx�1�"O0��0�Z44��"�	i��1
"O��� �<Py��S.J=	C`��"O0�{�Dܔv����l��7,�@�`"O�L�e-Ϯf��Z��$t��"O�(h�Y��|�R$ݽ��b�"O�YX�/� V���cD��	���0�"O��p�]-�-���ΊtG
iQ�"O���UL��M�(���A<l�5"O�d !2
��,�$*���"Oj���L
ClӢ�u�)�5"OF�H�Ŕ%��+�f��[��t� "OAk&��$��D�OS�+��q"�"Oʁn�l0�ʇ���o��A�"O\H�C��1f&
))[�c"O�Tx���w8*�ؕG�_F �"OȘ�Q�D�!H�������}S"OdC�|{,��w`�ut��a�"O� #��ƫmW�,���D��M[�"O�`:F��*������F��A��"O^ӓLI=�(`s�m��
�4R"OP���I�;�`�k��
5�\`e"OP\�Q�^�@a���i�4�<��d"O±�����9i�i3�
4�r5  "O�HW	_�z�i�Q(�?k���""O~1�
BФ5P�ÿ|�*�"O��F�1j�1 l�!s>�b'"O� ���s����jN*o��V"O(�P�L��o�a�˕ \��"Oȣ�?�\<�WIȥ$s�X"Of]��$�*A; }�ǅ�)Y�!c�"O$�*��O�,��mp�e@F:��:�"O��� �Y)�H���4�{�"OAȵf(gzh|�"�*=��G"O�x�%�'���� ��>�"�Pf"O<�҄n7`$	y����d�,#"O���F+8Z};F(B�G)lԳu"O�+hJ2u�4�u��Y�\�
"O`�iT!1�ֱ� ��+�ȱ�'1`�kPiɈ�z��!�S�m>L��/������� Z)�B��Y�`A�)�$�^��t�ɑ6
B��ddFG��d�J~�FD��_Hʨh��@�P�i*q ^�<Qb�K�BS����_5BO�@
���%�>�+2i�?-�T!�l�`���E��=�Ƽ��I�4iJ|�d�X�^5��ȓ+M�H'�șs)"����/'���֬�"�:�.�,1��Q�v
�|F|�/G�*k
�f/��Mobq��kN5�0>y�×?�* �H�KR|��@���YA`I"u+� Lk`Y� �׸L4�ɚ	�zy�-H�nƠ(bEb���"��4FxB(��&4r!X��ż!��ň�HY%wĒ�}�	h旿S�x�
���;Aވq�ȓt<x�� 
���򲭞�"u��I!͛�h� z^�x�P�K�z�襑��s�a�ƊF�v�إ[7f�ʘ��N+T���7._�sW���g�D�xU+�&�:cr�:u鑾v �CB�O�r��)G��(O�U3PCɖ_�F-��f��O,LiQ�'ˌ|agF��b,*�w�_������(t�e"���}�~��T�^_��!��	00�t�£�N�)�l���#�`#<� ���ȡ�K�<������W�o@"��+�V� �\�I�d��pHA�:;�C�ɞw�Щ�.ާLvP�J3�^�E���z��!r|�b�T�l�Z��˾7+Q>�]<B�r�/�j$���n�=|��C�IKd�T��
X>2d\���kN�4� ĳ@_�9��`��̊i}fH%z>U���	�E�vٙ��\�rբP�Q-

����½
	hqf��{�Ӵ$�ڜ�0$K��|Mb�-�b���݉�p>iemIu���!2� �r|.�BF��M�'�9�W�àT*�t�Eh�1~e�]:������ICOZ �0��'>� \ p$�&&���Ā�i����\?TJ^D�C��`�i�� �)KH�@��]�Zd:@Zΐ�)�Ҽ�3�=�9�h��ÞB���E�f��#0"O��p�j�-h���
�n rl�
X-g(�݃��H�%�:��&�6/+���$���P	\���	F��i�����%P�ca~��āi��1�r�����з�����!%�o��d�H��2%CN+^���r�IB�P02$�ݪ2�<�s��f��#>iF$:&FD�XSj�6N���ŘbJ� �!yI<���$M�&���ѩ0��������N�)����e��8���= D賖ض����O���F�.K����H~┫$h�~���0VL|
� �_�<�c�\^n��5��HH��i�/}����{�l�3��Ty���a}n9i�<���w�N�p�ҩ�
@q�� �Yf���s�xkq�����Iy��~��l	�� (��'��p�'�(�{��7��	޶`�N2,O�a��j]9
p�t�ò_�z����I?X&�Y�M�"\�����$�6����fs,�����@0l�A �ϐ!��3�j�<O,
���0DRџH���kr�� ��v伫u%�4\ �̳"(�	K��kCHޛ��IE�K�2,�R�UB�C��s�$L� =T-�&�'=�tyBm��<��M�;j���+Z�gTaz���A�Z�;8BTۗmޟF<$���ĔG����	�i8�)�
W�*�hr�9`��!�v��X��
��� �0Ahp� a� �r���	1z� �"-i[��y��@�'	�"=I����i����m��=KF(�s}�(�F<�솟u�.�s eM>w°k ��JAn�[S�G���q�9Q~��fm�|�$��%�Q�B{��oگ]_�l������C����#/�o�L>��w�
d #&^-Q�]�=��C��)'��E�p?���0�ʄ{%P�pF(�t���H`~EI#i��IwJ��;>O���)#
EȚ0E�����2����̚�;�D}��h�n���R�.�N�(�O&$㡄M�[�XSv���O3����D�$jx`ǅ:!Sd��Q�q%ў�R ��:^��p#�FشE٤5Cc�����F7���B%�?C�� Y1�*�cpoKn�����Z�zHР0�l�5����[�Vg)Z�怂��є����q�ѕ�'����5���/���:a�ȵM�H����4�yr��(B� � 4E��7L��ʗ%AGX� � ��<��.�d�ht��;-|X�wE&����:p�@ �nQ�3�`���`�d�B�ؤ�)�0����֭i �ʿ.�H��iZ�Κu�`T���8i_�Q�i)_�Q��������5
1@׻;`�h,� ��Ix�E�J���ͽM�0\�'���B���H=��`5��.�ȁ�		D_l@��KKn8���dǾ|l�y� ��\b�"A,|�l�ړ��/��4��C�!���a���kl%��d�&�E*N��ŻC�:1�!��D��f������(����2<N��SeVi��u�K[w��PЧ!�r�x睻F��t�=�f  Յ�C<����I��ypS��A���%��3W�0h�L��w�Q�O `"�J�]��I�$ �_!d=z��D�����r�R�Cx�	"$�0s푞�i��˪8�v�sR!�|Q��	�>� D���
 2_,��a,��o�ƥ�PG��n�� ��B[FR����F1
Ѳ�\M'�C�*̉7���0m��d�p
D/z�����|�;BZ��z$�����q7�)]VȓD������֖}Y*��E&	
p�H��	�nlۓ����ɧu/O2���Jἳ$̦b������W��<Z��Ex��,��*�)�6$xt�A�|��@��,a0��s+(}�<�,уS�Z�#%�	8Jr>�s�✾]t]ؗnRT�N#>CAއ0�^�ѳ���K{�LH�¥?�u���bˈ��/K�Z�T�3O��+�����)�O����E@N���SzƸc�O- vB�'%����7�8sGyE��Y_�I�Dɖ.EL\Ta�!L=�y�˺e􆬨U�͸|�(XU��Y@��YBgx��ɳd��E8�I|�>�(�+r��n��_dr��$�H�<QA��;!�
�J���>�F,j���B�<��1b��<���t `Q�RV�<1`DX7Tf�hd�(�Nճ$
N�<��� Y���S)ّ;`k�ƞJ�<�Sh'��A�"拎j��3JO�<�e� *�Z�`�~f�ѠPO�<1-�,%Vt�EG&�|��E�H�<�%��42��+Z�;�
0	�@�<Q��N3$�er%o��4��ny�<	㛲x��p8�
�!rp2�*v� �<ဢ�	�l	ϲ ��U�'-�}�<	��
7+��h�	&=����'�v�<�G �z��8}�j��@�{�<�gT+`ζ����_���:�f�y�<��Q�j~V�jci�>�2��s�<�p�B�9=q:�B��Va�\b�NWs�<ٳ���}���
��N=�D�l	r�<��
�l:�h	@�Y�K�`�&Be�<�Ѯ��':|}*E4:�0�!�Df�<�j�^e�R�B9 ��I��F^�<�v䍇U��ಈ�<�2q����~�<���B� �^�yv&�-�^8y�W~�<�a��\Q���)i���M^~�<���
��uQHȡcJ�[�z�<D^%b�r�
E�W"�,`;�@x�<�u��Hl
�cU�a�*q*�r�<)Ҧ�,j�8Bٶb��p"c�On�<�Q"�[ﴠq�V�{�8��3IFj�<�ba�#Q p����]�r�Íg�<i�JQ8h����gN�4���y�Jc�<�&�dc��]��j��8Gtt��'P�r�`�*ir� ���@ty�'	05H4��Q�� �m�	��L8�'%p��0j:h�j��;:���'70�WϙMJTe`�H�J
�'B �EK-B�.�0��3�@��	�'&H�z��J�k�.�`�F
�(�	�'���åFQ��$�e��o�Pي�'0��-�#y�f����ڂ=G�!��'>ڱ��@��9Ц��R�3�(R�'�<�{&M9�.i�wM@&4�)��'��DK�lC}>�9�t�F5/Xt!��'J�=��Jřajn��Ҧ�;+�,���' �R#
:f�J�٧B��42��'׺�C���Z(~H��&�G�����'����çS6(!�VfĒ�,tQ�'�Q���ן/�F��@�V�0��0�'z|1c�#3������=!�]p	�'  L���2:_䍊D-C;.���C�'�JX����)���I�h�P�1�'ؠ kA���wȠ��ʁ�Ѝ2�'<̑@���;8�x�ƈ�	9f�r��� *hdD˿0)+ҥ��w	���&"O���F�Lɑ7�?��T[�"ODͫeHӑH	:�0���"���"O���`�6�Lh��*�-$�b"O�lbw�ٴ��%�1*S� �p���"O��mŎiQ�X"��ۄ�T4!d"Oн���t�<F���T5"O�-xU��
^I:�s�F j���"OT=�v��0^�Y����[��9i5"O�@��i��V`@3F�iԚ�Hp"Ox���m�0��QKA\s�5�"O�ػp�܅ ����`/����X"O�(�@Ҿt��-�T5��8B�"O~�@��V r� ����uڐ	� "O�X��ɹEgN��AK5K:N���"O�0q�J�j�豒`-�;0,��'W�0�cfH�^5z�w@~��5i	�'�Li2HS#}	��)H�jZ���'��(�#��}|�5�O�~;����'Y�a� �ǚb�6�i�O"l���'�2Y3���0 Չ@�Kq�r�'���M���k_����!�'�­!�Hʮ{��*棓?�z� �'Xҙ �nD��8Lӆ�Ï=#��
�'� ®>
�i`6)��d�ͳ	�'�<qQ�a��obNE��MLFoؼR	�'\�� ���![�4r�j�J.F�	�'�F됏;��{�i9<p�ū�'�6X�U�g),P��df��y�'�E���,-Xqc��!/3l:�'�ЬH-�/:�1ҥ�H��qq�'�bm[doު{ʌ�G�Y<��
�';�9wh��(Q�\N��4�
�'P��A�2e!=aW�A��:�Q
�'80ѫ� �!i¸���C::�`���'�갺W'����	�H�3�ܸ�	�'�9+���-����v��` ��	�'op�q�v�J��&9�(i�'���%92�~AasƳ�)��'����U�	��Lx�&մehM��'1�5�hL�K�j�"�BY�S-�'���Ha���kG�/ʪG�B�'�h X� +	�H�K"�ˁ
�th�'?2�:�N�g�j(sdeݕ{��`
�'O�H2l��^��I{3�4Z���	�'���a���2W|�S�\�w�����'Hfe��I	ݰ�a� ��%�%��'�hW+ػT�ά��*@	�XX�'mdrpB�"DQ��!؎�n��'Ƅ!:R/.-�E��!����e��'\�b6`��g,� 1(�8���+�'���G$�I�Dۧ-�.76Ei�'�1���UP$��H�����	�'���g�(;�����L $CZ�S�'U�E��� �-�ሆ�;T���'پY@E� s���*R	�*���'���2Q TU0���jR�T3VA�'���b⊗��<�����Jghr�'�v% �瞟q����<��]8	�'c��V�b_L�#��,	�n9[�'��3A
��v�ۢ"�tVP@��'��������jK�����c��@#�'�^ة6#��d5�%���ñ2���'/"lp5C��v~�� �� Y_�2��� b�e�$JR�ycLO�e{�0��"O�)�rk��e�;E�J�>\|��G"O�!�Ĉ(���A�� ]N��@!"O��JA�F.RA��;@�\�D"O��3�͕%0�t�᳊=�|X2�"O|l������}�����#"O����BH-���ؗ ��d{�W����.4w&��掜5m(� X8q��C�Ip���.y"@ �1O
�hMR�"O�(�6�� 3��bŮշxӺ��"O�ٲ�ƞ`�mk��͢N�H��"OX�SS�؋|��p���M�(�ء�W�'�1O�ܒ��WY)��!�Ώ�V�� 1W"O����FT�O�iQ�)���r"O���4厈#n]z�e�t��"O,�f�gb$b��=�lt0C"O
XZ�`/ ư4��#����,�"OV��+k��Q�C�(�XKU"O�����)wT	٥�S�(���"O*�@@E��]n���O�:M+�"O�����8P��� �c�f��A"O`1
T�؀� �d`�3J�$�X"Oʠb��Ąt��% ��t`�J�"O�u��]00�@�A��R�kP�h�"O�U�ro�+�N�5*C&Ļ�"OZ���?Ԭ�`MS�Yb��S�"O��s�B�<_���A��4P ��"Or�3���~9�}�C�V�_Y:%��"O���&�"��J6�B7H����"O���FBBYGN=����	#�� �$"Oް��ѽdC<%C* &(u�5��"O�DA��G�k�$��)?aޤR5"O��c7�^P(,$\Nu�@"O�8)�"����8|BP��$L� w!��;V�V�N�0�T�X�E	:,Z!�dO�
pʀ���*�>� �ʾE!�D��k��!�Ytق���CP�v.!���>�x(P�n���X`SBǄ&!�DIO�k#�Lz���{�!�$ i�Q�	>(�����w�!�dH�L�l�ɦ�ݔT��V�Z+�!���y2�H6�Ӑ���O|� ��n����h�ofȻ5�A�n�P���!<q⧎�A_)���ˊb[`��ȓ?�ʴ ������*>(u(��ȓ+�DB��D!�X�ã��lj����A�X`��3y0,��aU�Dq�Y�����;�L�>"���,��%�>�ȓ!�1�)�Eo\AY��жe���ȓs(��ذ�ʒ:�D�B�ֱQ�)��[RС�5�R�>�������W����bБ�+ 7<*���3�48!���m�Э�d�.)-����*��s�'�x4��Y�C�$�a���7(abe�
�'���ȣ��H�|
�	�'�֬y
�'Wra�7O�#���p'D�.P 3�'�B��&7po���f��X�����'B�x�BO�K�Dq��If��C�''<1c���?Lg� dE��:��q�	�'���ۃ���?�8���{`���'#�-�g�ĠN2��[#���T��'�@ՁFD�/4��T���]<|�ZM��'�&�2�瀮r����甀pΌ �'S��r���*���*��~Z"u�	��� $���W,1Pla�BB����#"O�yW��� xs�!9�x1@�"O�9���H�@uR�ϛT����"Or���]�DӮ�;EO�<rR��C"O��
2cJ�s�nx�&ɋk���9"ON��V�U�_1 �Z��� y���"O*�K'�\'���#\!m66�;D����P*	BL��H(ԬA��,D��Ѱ	���,�0���J(n�V�)D��	��F�5�v�XW�.�X��+D��3�,pA���u�7E_*��C5D�4�D��"�4X�@%���QB3D��� �ifI�'�Ӫx~����>D�|#�*Q>$>�aj.P�c6�M*5�2D� �㜋7���$_����� 0D��R���2�h<��EJ���$���/D�����3-G�Aޤ2�+:D� :�!l�����+8 ����M:D��2VL	+@�&a:7��oVeYf%D��0·��LiA!�%K<%�@�6D�H�aG٣hi��ڶI�� Ś��5D�h:7��//R4��P`]�+VNr��2D����6l{�eb�դIQ��H� &D�`A���-�Hu��%ˠk� C��H��˕"`��Q���
�C�	�����wT%z�@�jI%:,�C䉮%��(L�=9X�A1#԰zU�C䉬�>5���'�AyCS!��C��6H�8tKR� 	���Q"m�C��b	�`�¤AG�<���3e]B䉬��r�O�-)-�&ʐ!7�C䉡*������7(��x!6o&d��C�Ɇdn�y�ĬŜp�ι�p��~��C䉔M����g$�56�����֪I�FB�	B։*�©-\���"R�De�C�ɤ.(���,�4�Z����]�xB�	+�2�xB�:W�$���~RHB�I�C7��x�K�<�
��%g^	|�B��:-^,��W���2NP�EH��1�pB�Ɉj�x��cL����B��_<�JB�I9+���0q���B�A�Ek�Yx��6D�Д$;l��PjURЂ%�va4D������HA�A��Qs�I��/D��rdÖD�0�@A�2��Ta��7D� ��
�E��0�G�":�<�G*D��a�	�=҄��R�6>����,)D��:Rhؑ~	7��2iVP�#�(D�ԃ�ŏ�^3* rj��bQ@L:D��*$�	Y��拞�CYP����9D��K��*Z���D�s�$U�p�8D�t�b��%� 4۶#^�pd�JD#8D���HZ��(bua�6D��R��+D�lS�#�t*8�Ʌ_k���`(5D��;��ڧ�j�J-�S������1D���T�B�f��p(�D_��A��+D���P��[T �!c��_5,U��(D�� �h+mh���kUY�48C3�'D��rs#���#1�F�䊱O2D�X�)ъ�.��u���W�: �!�4D��zwB�9��MXcAM�$��Q5N3D���5蕴IJ�`��ŋ�!��	�k2D��S�+�D -�q�	�S��v�:D�*w� D�j�ad/�e�Y�:D�@a��"����ǵ,b႐5D�� (�ɀlY!����������"Op���$�|�Z�s"�	����s"O��S��1?Z���4���]Ӳ!�2"O"PbP❋&y`U��Ő�Y���[�"O���S��43���D޾'��A�"Oh=YA�
h�6�*"G�T����"O"�SP T7K�Bt�[%�rt�$"O��Y�N�:g�M���јt|*�z�"OPX��sB.,�e,�d[�̂"O�h��T�� �9��N9luBa��"O��aJ�xprl�D��<1�2��"OH��L�a2�`���3���"O,����$D�z( 3�ܖ ��"O �2 [	p���hG� $� "O��"�&"�<��#�,���ha"O��;��)ì\S���2w�P�jt"O�P`�]*q	3@U�R��08�"O�P� E�XKd�*g/��;yVq��"O����H�c�( �U`�n	�Y��"O؊�!��l
x:��8(��	�Q"OLL�t ���-��ϐ	p�AJ�"OĳF�+H��x�@Γ,e�B0B�"Ox4�cٯE`D�� >�b��d"O�1`7�,*T���%��Ġ�"O����_�v!�e6�&%��"O^Dp��2.��B��TkP��"O2���L�'Y<�(��0LX��)0"O�0A$�q�qa�b��vp�pa"O�F@7bs�-[�d�Z`�2r"O \B��Q�,�!�bո/8��"OY�tW�"vX�r��@	n���"O0��6�4M��!ÕI_�NЈ��U"O�y*#��� 9��o� 'J��s"O|QW&T��ֵ[�(ܬri	�"O����߭J͒PQ�*��B�2��"O^M�7R2(w�4����v�M�s"O�y���,�`��)�iZ��"O�����_޴�3	؁PS޴"O�-P�'�#p=��+[� R��KG"O�m�
B5����;G�u!�"O��R�X�J��S���ubp�Q"O�q�IV�W�x�ZS�^�S���"O���<9�U�%��?w�z�PC"O个�n�[@��榊-_�A�"OH����;���˶(�2M,a��"O� ���`�` �Zf�a�""O����MAS�ZQy3��_R`��P"O��A>?�8�ǏA�GZm�Q"O]p�LRFيo�`d�	�u"O�|�C	�0��(�D��3/����"O���L(�a��V��H0ca"O9���$<�
����C�Z	Zi�"O4�z����+��Kqc�&S�0 3"Ov|�.^0�����-2��(�"O$�7*̧J�δ�@�1Š��3"O�Y�5i������y�0���)D��c�.��	��9���L\���! &D�l6�P ���aR�U&E������"D�xyv�((�,%���M���`�G5D�p�����1����(�5�'D�(�$��D,Y���:�����"D����P2��$���B���.!��m���?n������H�!�$Ǝ'��U$��6�����ּ�!�� �� u�A�M~ŢŘ1|?�uآ"O�}����<CL%����X8�"O2����SIH��cS�k&�3"O�4�g�ɚ8��[&#^��2xX�"O��"� )���H �-�H�$"O�!��/ �qjD�9�h�"O|�wǗ
UN���ԃ�Fq��)�"O�a2� ��{�\��B�-P��"Or��Ca &*����vJ��I7��C"O��;��ο���6�16��Q"O,��wd�b2���LX���"Op ��F: �I蕬*	��x�"Ob��0���i��=�ҋ_2G�ΐ�"O������W����&AE|Ų=b�"O&\���P�=Ybi{� ҙ/�}�B"O��Eʋ
Ș�jfn,!�L-ZV*O�R� ��nUBE��&�֥#�'��i��m
>��C�h�s衛�'n�H2�؋��	��"UA<�i
�'�Ū�C;�ahя�J<�q	�'|�hY?x$��+�A�&x"�'�D�@#�Voz����;����'YL�2�oU^�*8�'L9TL��'���B�.�`�J��Cv����'@�]���
:�f� ��xDbI�'���c���V��(k� E*jZ���'	:�'��8�J���?\GT�B�'l�a����PM�Xr��g�^,��'��H��U�.�k��W��Z�'�:9�ff�	 ����g��uG�
�'�F��ノE��lY0�^�a�t�	�'�d����Q1Xrʌ�`끨+�]��'��}Q�n�-J
�S�K�Y�����'#��B�'`E���K �V,��'�f����S#��#�M�����'�J���Y�Rw��(�fݳ��a��'s�.���ܑ�J�r�x|��'�\�Plܐ�d �R^���)
�'�X�*Ǥ�7.CF!�XР�	�'����#�'K��q(��� L�m+	�'?l=2t"���0�ed[g� ��'�>���V;(�&�KУ߲;i��*�'��A����#:���� +Q�>a	�'��ӏ՟G�\��j�8Gι�'�,8�#��h�QC����a�T�<9���D�S��c���V��j�<)�bA-4�����ό4�
�G�@gx��'Jt���쟙D�J� ��*4�r���'ǂ��%^ ?n���2�Z`x�'א��u"z�s���!/J�'�B�y`#ʧet,A.[����'�t����o�͋!�f-S�'
Хy��ƒc��h!Pj���I�
���d��u�  �-��~��Z���3g9!��\��T�J�IN�G3�P�T�ߚs/!��\E���G O>|8!�P!�a#~���X��X��	נ�!�ӑd�b�h'|"rY��*�!��ֺ+�.����>���gN�`
!�$W�_��|��I��e	J�`�(�
T�!���0r���[g�'v�(�قʎ�)!�d�2`��=㳣Wu��(xS	�2F�!�R: m~�� ���#� �~!��JM�vQj�f��D}��,X�!�� ��I��Y$h�-03͒!�Z�$"O�[�g���xa
U%3���"O�A�wI��q���x24|����'v���	��IE�=�=90�����$�S�Oj�xEnI�X��q��D������"O�L0��ߤV&xY`d��\�L�2"O&�Y֭C�iԩ��\&LP���"O��R���\��	���N}+�"O��f�H�X@2�xP Ǒ
�����"OX��B�5e
=��[؄(�"O� ��1�����`V�7� �G��7�	V̓�B����"r�!���7'� @�ȓh^���EF�4P��K�j	�D�ȓ?v�u%Kc�Ҽ�#����
�'qh�:#��1a]AHJ�*͖��
�'� �b�	s ��6d^<'>�

�'�8i҄�U i~<(�!�!l�)k�'�I�K�
�~8ɕA��֥��'3@�0q�G�s�<���M�c~�K�"O��*6�3VU��F��n���i�"O�:��S�KED!�VC�v��В"O��jR*V�|�ddʡy��CD"O�=�
�#"�y�e�{m�Ÿc"O� 3��/�����9��pE�'�@t�B-]�@�h��,�%9���OB�	�`�"5˷+��p�D�n_D�b�"O̰��J�Nߊ,T.8����y�"��^}z峕�I!�]���
P�*D���7d��W�T��#c�
{:�tA��(D���"�<K�����O\J� 6e(D���T℄~4TQ�tA��U���U"2�O��I�ܕ�����4T�`g�,TQ�B�ɓ~�H�"���5�zE+��/�jC�ɖ
͛� �(@ESQ)�%�JC�3k ��2	 )��U�� Y>�JB�	��
q����S��!�j�?&B��,R��y#@*�6��m�O� G�B䉺Af�z��v)��3��A�2��B�	&�x�R)Ph��}Y&�_	=}\��F{J?m@�l
4@x�R�"��2Fb8D�����g�!hB+jgl���4D�l�#�W���Bw@�,FW<���$D�@�pcG�>p��E�N�|.&��4�'D��P��� |�,�۱��3��%G�H�<�`a�M�X�5�^��ҧJ[����>�,`D��Uv<(t��7\}�8�ȓ1+���k\����A`�,].|�ȓ�llr�(� m`�!yr`�%cJ�ȓ}f�E��59�� ��%Ξ`���̱���C�K�:�Ʌ*�"�X�ȓi������a bո���	t����W|<�6͎5�"ApB�C�j]
x��%Q ��͝�x��X�nKG�4��[_�@���/J$����? ��ȓY��X1րZ)h�{"i�,Zz�q�ȓ�V`�d"T*�*��b��Z��ȓr�:`���к[�`�Q��|��$�ȓ^2&��Q�8 :I����<o�*|��OʹJCM\�4� ��U�ǃa�H��ȓi�̌��Â����"T��\
h$��G{����;U���b�.�d ��ǁ !�$G	Kdָ��ӌe{�ؘ��Ȯ�!�$� ` ܻ4"�J<.i�E�]�7�!�$��
����Ɇ�4F�� !��n�!�� rm�Wۗo���c��pŻ�"OP�RG�X's��5�rc��S�� T�'����DQ��r�ó��!P\���pK-D���`f��E,fy��ޏd~x$��,D����'H�@AG\�iK ��$j)D����/C�ʴ�p��ګB4l��+D� rvꗅG�X��JC�-��d!h(D�pbu	�'k�ڔ�c���=��uyr�'D��sEa��N^��g����@��@;D�l��� t�ݙ��J~8<H��9D�H�s T�3����4�um���#7D�(���@$��Dч
� *�h��ª:D��c�o�+y���0Lդ1��+fj,D�$:ՏS?'LI��/�c�ԕ��%'D���0����l%�g/;E*��0,9D���I־����d���%6D��@�e�5!�dt��%z<���2D�\p ��B�d90���)0�N� C�$D�T�5װk�0��nֻ2>(-ۓ�#D�xE�h������T�s�X��w�"D� B�4,H���H�d�j`���!D�cE�I nӨ�{֯��Z<��%D��2�`��s�8�]�` �Mt���$'�8D0�3�F����p"�i�|C�	�NP��a�F#��xc�AD#o��C�	80l���IWjFic��%"�DB�I�9|�"I����6 Y�a"D�h�Ǉ��8�Q0�� H�$q+?D��
@��������A��\(�+8D��W (� 0�$�o2�484@64�*��S�F6�C%�+gb��Èe�<�B�PA��M#8n��+�h�a�<�ƌ�z��k��6z>�i%�[�<����E�@�®�2>�N9wk�a�<����Zh��)�垅Q�\5�sHy�<�7��&b&���� ��<|б2��]i�<1���?��q��$�>�� p�iIi�<	�m�6W1�E�/�?P5��kẼM���hO�~�VT�Vb�@�M�Qa8Z46	��p|�|�����o������R4?Zd�ȓRx�Q$A��z6VL��A�,i����c:Nl-�=1��H d��L�~��ȓ�>@��F�� �1/SU_��ȓD6���3&ʽaa2�B �:6��1��N��RE�>b�\�P錶]��ąȓ;���:5FA^�勥����i�ȓk�� ����JRpIjC䝕.*���)NԱ��P����$Bs����fDP�Qפ��"�(��D����A榴�LE
eu�t"B�F���P�%���
�O'�a"�E�O�>���I��@F̗-�N��B@��dD{2�O� IPtŊ�jI,@�E��~V�]��'����ެ0'�`�T��u���*
�'���{CEF9Y����ɞ�j�2���'� =r���)9���ꎜ\H���'�
y�`	ʰvj^59��G	&���b�'L��
#k�!W1X��[���`��'�8�Ƀa��a��A$�_�yB͒���hO?�)Cj��0���	sbT +�<X��@SE�<Ia��-RU��@R+#ny����f�<�w���,��X�s�^ J[��*�b�<)FB��>Ů�(g�C�EԬX�	Hh�<Y��ì>
 �I�)MxY��Ni�<� ����Ւi[�=!��&dX���"O����D&DJ �猙�V�{V"O�s�&�8}�N8HFBC��X	�D"O.��7'ƀ
�XɋboR��|(�"ORU��K�3i��W�����1�d"O���d�C���ĥű���[�"O	y5��2"����K������"O�L{s�Wo�,s�E��I��d"O��Xfi�Y��4`p�=4,�JA\�$F{��	Z�h�X̫3
�,�w�$!�DW>)~p`E��{21���%v!��&E���"��&f\� �EN3@�!�� �FM���S+"�9�ùe}!��6Mh^\F�����H� �2:d!��N����TjO�>0L���RG!�ش���CW�2�j��!��O$kEp��cٶ<����Ԩv�!�xl`�PeGM<^�؁���'=!��	A%�D��gշ-g�FK�nORB�I)���'$�4��b��	<I�B�.����F��]��E^��]4k�&���>sUFA�p!��K�!�r��b���ch���oZ�&�!�DD4`Q�a	�"w2���-��S�!���e1d�ύͬX;�L\"K�!�$�uh� ���:Z��P$�ޮ<o!��@EhH1����j���:� Ǒ*l!�$�BT(��6e�gB(�d�%��(�'u��@{���Z�a��ާ^�PE��N�x�q�J�y��}��-N$a�΁�?i���~ҁn�J����F��"��	E�<9P!� X"�j�i���R���<�e�6j��J���m�q��%�y�<A#+@!!�)iG�x��MB�Xv�<quGT7i�̸#��T�4��-yWK�K���&��{lX<x��0�p*�:#�dyᇊ�<	�o��u�A��G��Ax��Exr��K��f�О)b`�H	'�y�`�<(�ӆ�)!e֨RB��yR�՘c�Ѫ�؝%mhr^��y�Z0#�N��F��:�k�Aɛ�y�R O�|T;�ѩ���j��&���hOq�R=�f�X�ok^5� O�:\�a2`"O���1���Mc����a�,"�(��"OL�2.ƒ-���UA��� �"OQ�U�X�?Ld�pJ_
�M�"OJA�.^�IO�*A�x�����"O����^��D3'��5��mj�"O�!��au8�`��"
�Z�"O�<B�a՗i&�����D�����S����I  �*9�_:��^7�bB�ɠZ��sc�ɷEp��o�^B�	*e� �)S�v���#�%�7u6B�I���Y1D�G�0nP�r�ˏ.B䉳GrX�bjDS6	�X��C��AKԨ�S򀢔"�?c�!�$0o��<!�E�~}�aa����&�!�ė"o�U ��
b��{pڜ5!򤉩X��l�T�4rL�-����~C!�Č��P`���5tC�|�E��q!�DX�
����alB#Hߘ�D��^!�N�&<�iR���x��0  _5jD!��$>R̀���J�f�읛fΗ	G)!�Dݝ�,����c���2s�1�!�� ��i���!,�Ԁ��JL�n�)#T"O�)x�Ի~� /�30��v"O�aZ���sa<H�r��9S��i�v"OD`0�P�Jt��GЖ\�B� �"O��@H]�b ��e
4DQ�x�"O$)Ya�2E=|Y��k`� ��"Of}0r`ܨI����͌I�p�T"O�i0l��BK�c*�⢄��=$!�D7��͓P)�t����:!���kź����?B�[Ak�)p�!�$��,	j��0��i+"`�
!�X9Z@�VEʭT��l�P�^f�!�PUf��Jv�Y�3H �����'Nў$�<IRիl�L4��b63�Ш�%~�<)$���l���57?����u�<�e���g�a���ӪB׼}B6!Ms�<a�,�7�v� ��¿���1'�r�<y%ަ�n�pq@�3Rv����F�<�F�� zؼ��7��9y��s2�g�<�%c�;AXp��K�=T��+c iy��)ʧq��8���R.�>	Ȑ��؇�z�0	)W//HQ�S��/FZ]�ȓ���@�	���A/[	z`��9���;AF�Uy���2�%,ضɇȓl�B�v+ԃP>�l�'F u����ȓ"��I��k_)u���+�$D(n�h��ȓ4�>�j!�L M�,���Rc1BM��	e�'G���)�?U�D���Q/Hy�'��0ы�2��X+�E��̲
�'ۀ�1��F����a�8���Z
�'P�����>y��2�A�	�'�0B�#������fExs	�'}���B�$r�ơҥMcx���'�N!��Ô�sZ03!%@�Wb�� ���$P�+���	�@љL.�x����O�!���":y��	�9Df���-X��!�D.l.4q�a� -�Ԁ�N[�!�$J��M(ҫ C%�� cʑ*��B�3CzaxE���ɠ�e!:�B�I�.���[�]�I	r�;)b�B�		?^���!�O�$x�@b�$C�B�%-���s��V��P�˓7,TC�	*>|�s"�X����D�ӌIV�B��-t4Xձ��0^ٞ��C�]�g�LB�IA������R���8�䍛�<B�	)d��S�o�Flp���36�B�4�9*��A�Z��A����C�I/#�s��!O�5h�F�5`ɤC�	,��P����/#��X�g�\��B�I���@��J�m�`�o�?1P`B䉺X�!�V�֑ ��H��1=pC䉽@,�tSq�̋Z֖���iT�4�C䉱]�R�X�Ɍ p����c�fdC䉟#��t��jf�r� ԭ�1hB�ɳF3��+�dE�	aR����C��4�OƢ=�}�̆8���`+���(��a�C�<@��}^`��G ��.8J�-�@�<	� 
��1�P@U=[,�8�t�S�<�'G�Y�v��r���?���X媅Z�<)p)Q� <H`��i�!Tֶ�S��b�<�N�fTBt���]	T�.�6/E]�<y"�/�l8��+�IJ���&�IW�<!P� {"���-��#Z�l0(^L�<ٔA *��U�A
��"�d�K�<� ��{���u�6��V@���P��w"O�0����Pi���>y ���"O�Q� �UBGN��TkJ vZ1�S"O��i3��
*>=�	Q�gN�E� "OR�Ab(3RYļ�v�ʪ[������!�S�	�3f��qv�q]i2%���0�!�$�#yL�geZ*T�T5��̥N�!��2�`P@ -�t�
'DˤP~!��3>�J�x1'	28����aF�m!��Q;.0x�0��r�0��� %M!�R�z�质��L `,��`�͓^@!�d�/C%|��c��PH>�����?E!�d=x�v��& �;)
�� �c�!��|(N�s$�5~z�-��aO<i�!���y�z(Y�D)2] �+ G�!���F{R<o�:b
H͚�՛�PB�	�e�Ȁ2��V �^����x�:B䉡�:!xDeS'(�F�Y�jP�W�B�I��
@�]:N�|S��7�C�	�f�����જ����2�C�ɠ*sF�؁�
�c�P�c)E,t�jC�?>݉��6X�Zċ+�wWB�	�"�@�4I�d�\\ꠠ�

��C䉌#{�䑐���R<>`Z��#�C䉓n9H�e��#�J��� 9&B�I�\I��aC����,PC�($�bC�	j���U���{�TIPa��(D8C�ɗQx��h����TYڣ�C !EC�/��yCW*�<w�>�H�_� C�	>,+4T2��њBF�8�S�\W\C�I7/���)§�0`�	�-U r��B�I
����cn�"BH^@�D�0d�<B�I�JH�a	��g� $��n�)$dZC�	�Z�fi��_
�Sf@��	�	�'E��jS�Yi<mP���>� ���'ĵI�Y���j�L:0��5X�'SV=�˘'r�t��k�29RPEa�'
ʭ�G��h�� �U�)�����'��I��L(:�6���X1�H��'\I��B�Pr�X�f��-�H���'	 ��wa�yMЍ�1��$cB}8��x���>e��e1�ĹA;��Hr�4�y��6���#cR�3�J�S��Ж�y2e_73m��j���9T�0l!�Hݳ�y��+���R%T�D������y2g�Q������ӪO��CS���yB�ϒP��ibP8[z^iifF)�hOB����=a|չ�L�	0ū�&��:�!�D�F��|1ň�F���G ?�!�D�;Ⱥ�Z (N�%4P�!QfF�]_!��_�*/�|�J��p$b�T2tj!����d8@��ɄN\!뱁W�^{!���<m��㕔b��x���g]!򄜇nC��Z	0Xp�SKB
kL!�D�W/l�s�+O R��
V ���$&�S�O/��c�O
{H]Q�C�?�h|HG"O`�����.pȔ��B�<7w]q�"O��s�� /�F��.ެ9W��	2"O��3�&�<֌	��# NB�E�6"O�)Q��F����G�\4FP���"O�y��#�&H��GO�JD&����t>���l'I6�]��O�w�8+��2D�x�AO�����̕ �P��0D�9aU�R��<C�Qgc�V�!�� ����o��P-�:��E'?��*�"O�%��H/[��cFCJ�'Ƙ$��"O�T����2||ĉc��ʩP�d�s1"O4��p!
@1"�ĉC(`7&���"Oz���-�.�p���o�,� W�\��	,<���+��L�=��1�27��B�	�IK���Lc{n(���;��B��	Q�,���N�%h`��Њ<bC�	D� �S��4�6��
?vJC�ɚ0�s��02GDD-���"�2D����K�1�Z%�7)B-�$��/=D�(� ���E�<�03H�&X`�s��(D�[&�k��e�PH�2@��T�(D�\�$!��?�4�tL�P����r�8D�����kV����W��lȐ�4D��S��Y�J}NP��I��p�R�%�1D�${��
-�C��N�K�J��$�0D���W�G�z[<�J�
��c�@4I��,D�@z��Z�ZB��!���[[0�@�?D��b�G*�M
!��@�,�R�c#T��Hׯ��(��q�e	�8YH�a"O����XVzq�dM'%���"O� ��lU)s�\E$=� {�<���:�r��5��3����GCl�<i��U x8l,����*Zڇ-�p�<�5��b������#zV��e&�k�<Q�_+2�4��C�ܘ�/�]�<�PM �^�pȉQ� Sd c&�W�<��֓�����C�3#��Jg�U�<9-G+|1����7h}*13���y�<�a8&0��0AѸ@�+��Au�<I�V +4<�wM6=�<`ǦVp�<AA�S�����]+���#�$e�<ѵ�
�g���Yu
HX~�ӣ�d�<11�D6�l�c6/J��"A��a�<I�.� !9��*�HK]DZ�G�<��m�0�z$�5
��
�]xpAK�<��݃ ��9)�T�z��88B�CI�<i��M�K�zq��J�5���	��l�<�Td�(&��<C�hQ'�T�X�+k�<#
�xt��Ъ�bXSBGBl�<F)��j�f�	�6��|�-Kh�<!q��"S�"����J#.�ʭ(���<��%Ζ/��	h�KY�^��0���}�<i���Xj*y��j*�l(���d�<!��ƍuQ��[�C2_��!8��]�<a�NR�<qp�1��	�|:Z�@�'Kp�<�F&�s
! ����r�Cc�_n�<� ˻������=h�+QDA�<ᐍOs��aG.X�HIl��B�b�<ٷ�]F�F�3"�1[����VG�<aviƐ!�Hؚ��Ӧ:?d��!�O�<�gk��e�3Ҋ�n�v��էEM�<�����=�A���(�����K�<�U�߮gMN�PR+�e
6�R"h�\�<Y�TI8�b�'ץdRxJ�,RZ�<yBi�rY����L��CO�!2�U�<i5l�i�����k�N蹸�)�J�<�s�[,b�^���/:1������D�<yc��5W1"���fQW5ԑp��[�<��� ��L��"P������֟��R��(���h�E�+��:E���@"O�-�g���N ���p�ƢDbh��"O�y���U��|L�tߚPE�)+�"O� �̉�N�T��QC� �3����"Oz�abg�6x5 ]�V+2�y"Od���̎#6�`�,�?��-��"O��q4F��@��;{8BHk2"O�@��gK��D����\+h(��"O��3�b
1!�4T��H��e���E"Ob��0���
�)�W��"-t�S�"O��!��̶X�0h
��F��s"OLPi���i�������.A��h�"O�E�1C�%?ص�𠄠,=��J�"O>��3ǉ`pl�Y%�ŏH%��3"O��0mZWVup�	ܧ%�y�w"O�!�"��\�{�G�
I��e��"O
e৉� ���q�&i?����"O�ҁ���HA��[��*uKp"O�	�!Y�I�&�� �2X�3"O\I@Em�"~��\2�j���RapU"OX)�f�Q�	�HC?�Tt��"O��i5�(m���� �ƨ�a�,D�T��G �Z��$ٰ��%y%�ah�f+D�`8PAĎz�*c1��2����
&D�ؘ��� e��a�\���Q ��.D��1�_M�4�Z�cٿ)�v)Tg:D�4Q ��1K����n)i4�� �"&D��e��KP����jJ�a��"�����O�t'
��#*�/H���"OT�±�Q����4�' ��P*O�� 5��:b����Gʲy8P��'
�Cc�R֚%2���x��L��'m�1:�" U�r��e��t�P���'(*��� 	5!6����nz���'ϔ�ے*�g=�q�
ڷm�p\�����<IH>��~bi��U�´��)��6��AN�y�M	�cj�y�k�נ�Xu�8�y2�}a�'�78�kp�WG�\�	�'�3��(�X��� /ˢh�'��䑄[�R����OF�-���2�'4����*�('�DZ��4I�'��@�C�G�BGf^�R�du��'���A���nߒcV�%J����'�x��ψ�# �m�6�ȸDш3�'����dhR	Z(�a�_0&�v=s�'SȠ/Q�ֽ��ʛ�նu��'4 A����b9:y�!ܴE1~,��'�vD"�InʌM3�Ƌ*6`!��'�Z���.��K�!���Z+7���'2���Qe�2i�N���*E~%��'���Y�ːm��I1�f��|j��'K��c��)QŎ��r���Z�̉��'�r�:���cB�F0YT`��'�z��d$��H�d�[�}r0��' �e�� R���� ^��*�'��J0�H6VC��B�ʻa�bHϓ�O�mK�g�[�Z�r�ڒ|�dI!W"O�T�����!jP`6U�qv"(R�"O���3[�A�X��٠f�P��"OD��g��7��A�D�^���"O��6ř�F;=2�$�z��t"O�{"'_�k.����>_Ddʃ"Or��Ǝ�W���4�5*`
�_��G{��	;.�e	f��EĲ��x�!���yՀ�2@�A_��m��BK�q�!�\#r�Rf��#d��Y���E�{�!�D�Z��e�-��X`���D�!�� bt�c	��DP�)��®?z� ��"O�!B4�
�busQ�:�V��5"OV�)���8��h�d'�^���"O�L�Dh��:��o�K,���"O ���* xVz�s���=G��8�"Ox|9B�Ɓ$��Ӳ�	�M�5 "O�E11��w��vG�(8�tL�W"O�Z��҆	@��,��h�b5Qr"O(`� �=L�� ��2�8���"O��V����	�!�U^��CE"OH� �I�q�ZY�#)̏h\���"O��rS냢U8�M�Fhδd|5�U*O��ˣ��z�Fs0�[�N�ء
�'��I
�~��P �H��lܩ�'��1���"4DxR��zx�M+�'dP�xU��;��L���-�xh����4�h�`��,?�v���MN�z,t$����X�O��Ͳ6�J!K�J@��ʘ7D�X:�'�D�!0HE�]f���m�*�-��'~�z���H����e�="ъ���'�40h���Rղ����9��s�'��c
�m����R)����' ,�����& �!ۣ���,>�@�'1L���I>X+f�p�b&*�ʼ+�'��`��E������ߗō	�'3J\2���w)�Q�7CT�j�z4s�'�*�� nߓ�����g�^�B
�'Mf�����*̼��&�G�j�\��	�'�j}���3FF=(w)
�_߼	�'���e��u��2��Ǌ$�8(�'����a	zX����ʬ"�HiC�'�Y�5M�#~�xtӕ��cҮ� �',������/������WY���
�����-�	��럞%���6�P0,=!�$�V�.��Ӆ1a�QSD(L�7!�D^>O�L�f鄲�����,^�!���7�h0	�a��g�2��C�r�!�D
�LF��I4��mǤ�K1� V�!�D�4C��	6R�u:��K'<e!��m��`�ƨ��n �Y�8�!�DɠE�xБ`mU.>d�8�F��4�!�D�K��U\2��`'�R1?�!�D��h����&C6H�B�JY�$�!�Y�y�Z|�q�@�, �R��5.�!�D�p*�B��4YRU ��!{ў���	/|DJ%S�j���LIہ`L9nB䉆q"�jǅ��K'$�b��)g��C�	c�|�r�O^�w�xQf�p��B�ɾF�Щ"��#sy���Th�h��B��7y�e8vN�96dP:ć/<�B䉥^d���&NR� ;F��dČ%�C�I�x\1j$�_�4���g�/h(B�	��5{tKп>��Y;�.ޚŰC�ɗbl���5��RS�S� �8��D"O��y�O�6���Q��Z�7�l�"O$q���5�:�xEoT>&���*f"OCDE�y�B\���9`�8���"O$���I�}/@��EM�BPh��d"O��J�"���
�e�46�8�ځ"O�T�'ω�bOJ�hH���|�"Ox�pQCՓ�����aׇX��yڣ"O@�É�|P($cUC��nϐX9�"O&d��&յ*��Cߐ?�Rs�"O�Ѐ��ד+�6	vLE<���3"O� �� \�%�֩TL�b�^���"O>�!e� S�xꤊ��N��"O�̑�f�4�u��@E�c����"O�@�ի^X�� ���%?�|C�"O��Cj�(Lt8+�&X�(�p"OB���mJ�`45���M�S��i�r"O�u+�%��o�&�z@	���p��"O�e�X%iy^��e�OSѦ���"O�1�K��l�%�Z�0�>(P�"OhaR�Q3�T}x��C3-Kp(A"O�-�U)O?�X��4��:oF�Iʀ"OV�[�O*�mI�Z�H� "O��J:R�0pR��D,k��7"Or1��vx�Dx���\|F�Jg"O��P��Q��i�:ʸ��"Ob���e�T� a���*���"O6)f��W���h�'@�3�j�yd"Ot"� ѴR�����$�2T�"O.0Ta�	4��@#�T�t�M��"O^X���#ќ���Ǖ�JL��"O���4�K%M���qB[�6�y�r"O�� �6�XB�#�x�);P"O��Ap�T�,b1��5��m8"OFt�r ��NQ6�+W���R���"On(B!�J�]�������5J�Z�:�"O�a��
�w���1`��B�ȹ �"Oܸp���s�I	@��1J�"O,�Z �v�(0%���F(�3"Od�t!۱
Q��Hf�M;KJHJ�"OZ�����<��h��B�d1b���"O8��$��'!�r�3UH{'��؆"O��Pҁ;'0t˴�O:<�T "O
� ��م-@mj��@�uP`"O�={2��~@��K��<0 ��"O� %ʊ�K�xM�")G'�"(��"O(�:7�=1��� tH�<Du2y+�"O8y��"���as��8q�R���"O��e�A��|ꡇ�Xm|��V"OB\�&��&�i��LV�.�!�"O�\9��g"��f+�p��H�"Od!sU�M8|�q#�	�L�YC"O��V��"0� ��EH��v�~仕"O�mxB�G�BLr�M�
��&"O��:� A��-�c�� &Y�V"O`iF�@-�vA@p�h�a�"OD �C'�2���T�"���f"O�pR-�N���\���"O���w)��&鰀^�-,^t�"OD���Ƶ[�y��c*@��W"O�Gd�E��4��LĨ�X1�"O��	Ç3g��@�P "��չ�"O\��1�] xy\����G��Y'"O�	p��N�t!��e�P�' �eD"O�\���r��bb��&%�2�$"OR	��E� J@K��Ų`�܁�"O�49�&Y�|$��A(��q�8h��"O�}0Uj�9(*]��'��j��"O\���&��|��!��1^�*��E"OR��,�s�p����(��Aa"O�0��qHX��֋f˂|��"O
��u��(mS&:r�
h�"O��i�J���\T�0$K7h��cb"O�L��(
D�1�#��%�V("O�8����(,��m�1
����] �"O� >!���VC��*�in��C�"O��S��K1���#�/qI�0�"O\���8� T�R��s�ځ�"O��B��P:QtkȖnSh%�f"OT��B�s�b���`�,+E���"O��jAQ�/;*� ��N[z�"r"O��1��G!N�
�N�1%4@q�"O�U ��% g@)ۣ���0��"O��`��4C>��Y���9ͤ���"Od�%+ |�S,
_��"O6�T	�J>q�Ъ+A]�� "O&����߾~���hN�_W&\��"O<Ybc�*Ȃt�P�#8�(i�"Oj �4�Y�@>dٰ�>X-���"O�뱄˨
��	�3��pq�"O��y��T�l>\��ɗ(A���"O�����	k29 C�iѤ�0�"O�\yD�WҜ9Ǉ_(G ��3"OX����O�kp�5�g�I�f�"OV]�T��
WZah�R��L��"O�0���Kl$�)PF�U՘1�"O 	��
�?��JīX.{���"O�X�qa�N���1�=j��hZ"O��!L�5O �QbV�v��E�&"O�#6d�$�u�e��F�Liq"OP)� ��.)�v�ă]n��0"O��R�I!cI��b�h�<)�J�3�"O���CF	:�֙k��Ic��[�"O"�C�GD�f%"��׍�8iwD�e"OJ�3�eC-r��G@�+h�y�"OL����du�`6k8C��ʗ"O�]��L�{���pH�),3|��0"Ot�v��#���8tDJ�<T���"ON��nH�zߎi������!"O���T�A�@�b�f3�n��f"O�@rq��^B,�XI9M]�`y�"O����NP>	]적��OR����*O1���ǧz�n����%O�a1
�'wB�Ra��t]0���R�E�L�	�'�*����o�
$�4,Ӂ%la(�'��I�T�ƄI�T��D힕���	�'�\!Z��S�(��)�E�J*|6�L�'#Ƚ��	C�.K�	;��	�pMk�'ktX���W�P����Qĉ�w2��J�''�� *т&t��!A!��93��k�'^��aR+����7c�"�D�x�'�T$Qp*���N	�K�(�k
�'�@����M�2r������`	�'�̑)�����Z���(~̚��	�'���W�l=���I�tKH(1	�'7�̢��G�e��:g�:86����'>ٙQl@�N�L7Ȅ��DC�'�����[{f��#��vȤ���'��\���?@��l��
�?j���	�'��cA֖ZHxr'P�r̰=��'�-[FI�4�H`�a&͸n�pqy�'Y< {��՟'�<0P���s�P���'\5C#MY3qCO�wEdD��'"T@R�ĔL�:�� D��"��B�'����4@�	����bA�	�$��
�'0@%:E(� �$s���)�}�'tZo��PX�T�A^�|� �'x�J�@%t�K�;�h�'�%.�Y���9@�_/,�ҹ���� �Aʁ
S#<<�;�� P6)�r"O��b�eN��:���ʜ�:L���"O0����S�K��¤鞰GY�F"O���k�	Ly�:w��"%9��s"O@] eU5P�4����- *&"O|��D�Y3\�*��aZ�~|>yB�"O�� � �Go�z�@\p	|��"O�;�%<S��T�7�����t"O.Y%�ўyf�;ЏΧ3�J��"Ov�"JT5��B5���:�@�"O̻�Ԥi���G ؉�V�H�"O�ţ�G	�*�>���[$"���Q7"OD�`&g8j�2ؙ�ʁAf�10w"O������
C��j���V��!�"Our�'A(S�J�FĔ�P�p��U"Oxq��G2?5�-n��d��"O�e�(]�qú��'��-S�64�7"O�����K�d��B��:8�2"O�q�N��V²@[c�چ=iPA0"O��!��׍4#*�����Z�|"O�0�%͜lR�L�b�/`An("O �@�ȺN�b�� $E�'6R}A�"Ov�1ЎYA����S큣m;\�
�"O �#1���n��L˛@�p�"O恸6'��&5���Gp�L��"OF�0p�ִq���:
�L&�(�V"O��B��HEj� 6�+�T0"O�H5c��~y.�䠛���Z�!�$�'V��QAN%Mhd�a�5C!�d��LD�ϖ�	:!��cR�A/!��l��`0!�MEЬ�"�7<%!�Đ(���� A�<����%!��U�R�(�����]Y����vy!�d�)w�i�U�!]�ڄ�b�x`!�$U�n�$�Yg�б9��y*�M�`!���~�����]�AL(���͞/!��4o��drEÉ0T(H�+'u!���0E:!ʃR��:Ȫ@#�1�!򄛞[�0l�D��D<��B�p�!�\� 8x���R�_�}�%�!��z�а�2nԓb���!�Ur!�d�[7�tc4d�ke�9u��~k!�D�p�.�va�-e��B�#g!�Ćs����͚�Vd�H�]qO@���*5ؘ���L�������k��b�ʦ���J�B|�Q�e�%��8F%D������H���0b?��ZР-D����ԀS���$�ƃ�B<�B+D�L���߽v?���2	�����5D�X0E��r�N�zT�]�S��u*6D��B�E�1 �0bV���0E�3D�T�!E;0߀x"�)߈o�a��3D���u�E�Y�<����1c����1D� ��f�	���
�Y/���#�/D��B&/�0d�4�U#�����J.D�t(���6���	N�Zf��@V'7�hO��$c�H���RE�(�{�4C�	&{ �*���'�����ћz�\�؈��>�g?���|���LWb�`���}�<�Ra�E����4+�b=�FKZ�<���h��Y>��;Fe�1.׎���qy�)h�H(U|����A�ro���ȓ
�R(���B�Cb!L���ȓ.Bn%�u�U�N�$h��!T��44��S�? �8��_���CO@�XS"O��A�3<E�M�*	� �"O���Ł�y����A'Zn�#�"O�� ���@~�t*�9LSu�'��d1�$�'Xc�!�/Y>O�<�s�Ȅ2|�!�J�F�<��	�ają�e�!�H�b�M���3Hh����c�l#!�D�&`��SRm�9��k"A�t�!�d :u;:H(m� p$Ͱu���!�D��cl�ժ��f�h�3l�&�!��ەfT�3թ�60�D�@j�c�!��X�b̌���j\$^谑W�4
!򄆝X��\ءk�)l'��9�X�
*!���A��ʊ8`$6P�(u!�d��[ �I �L֔'� �h�w�@��ɝ_��5pD��H��б�I�-D��C�I$1K�Y�c'd��l���,-�zB�ɻn���8uM7I��(p�B2:`L"=A��?1�O �Ӻ�R���B��2�Uƍ�GC^�<���݆3{:��� Z8��j֟`�?	��i��?qDG�����&���,�hC�IL�x�f)̤Y���[��D	����0?���?�4�S�H�3|�B8�%Yq�<���
"��(�\�{��L�Q�[k�<����������A�8o���w��j�<���]��ͣ�F����=�P'�d�<��C�(Ғ�QE�̚7�>�s@��b�<!���e>�c�O��ް{�/�C�<��n�(*p��Ĝ)"��\�d��B�<��J�l�Ľ��b#^;EW��@�'>v���ϽjDNT�r�c��-h
�'�<d)֊:b`���˂I�mK���<�'�OA�UA� 3���sfj6�P�
�'|�����˧z&�HY"Ȉ'<��ٴ��'&��s�nuC���� �'�w(ݛR"O���sV�R�dE�' V*@��� �'�ў"~:7� � H��/ ��$��Ɉ&�y��EJ�\)ӤƘ�}��I�ɘ8�y�@ĄK��ANY�z?l0����0?A+O�qπG���ó+	�@�"O,��6Dց��S�b:�`AɄ�z>�"`!G�,������D�	Y�"O6)�aF�R��A@��x�pAj`�iTў"~nڬ��SS��\���`�8.�4B��v,�VKB�oά1��(Cn,B䉰����lT�id��hM�o�B�ɎQ��uRҭG=�,}[䤌V&�C�	�>f�)z���m��5��L�pu���y��h�l�奞�J��١�߇N�P%"OexgG�9 �� Q�H�ja8���tx�l23�V�i5ʍ�AM�Tu� r��'�O��I0[/��s�O��Pvu���I]�9�'�,��qg�
P��8��?L�J��.O��=E�D�ȱeaL���;O���G'�y��$Ƥ\Iv�]�-P�eLU�y�"���VŰ֢��"}���s���y�"�����"��rTqb�
�y2���A��S�.���.���!]��y)F
,���2`A�7	'���*���'Da{�� v��3*�6������Pxr�iX��됫�$�@��d������ Ob�C���sn����$�!&�<��"O�� t@�
'�0Ò#��)�R�i޶B��7)�HSe΃)?TX�$��*4jx������� � ��cA�)6�)�1}0��G"O���D �@պ{��Z"IKfXiR�O@���&_@x�2�V `&@A��X��!�D�ܔs��Џ|!�Y bȁ&��;CRa}R@X�LiP]��b��8tNTZ4a���d����$��I�I�&GxPc��[Ѿ��#o��B�ɒ-
*���ā�a���ʑᕪ�al�g�����&�6v ����[�O��EK�e�<)�c"\�Ld���݌-k��v�@e}��p��I�W�Ҁ���C�YI��١7��=	��	҃A�%p�W�\�����2�'X�~2���(��A*��� d4Z��b����O��IH�O��X�s�ׄF�vY�<%�,b
�'�b�����c*v0��O�=2b|8��'��!K �D!v�
a�1�z���'�:|aT�N�W��0Q�V<$��O>��BU l���J����#>��ф�	���)W�Ѧ	�@����-F_@CEN�^4\��]>)IWaĥJY�8���lF|G|"�'�*\E���W8j�H�s��"v颢#�(�yN�2�l䡱���֨I���M���$3������k�A�t+D�Y(ܺ2�6<O�#<"��37�aIEfx������j�<d�HRԼ�J�b��{v���1)�Ax���'�UÀf0VEx]����k{
�
�'����Z+B�3��<e���c��d%<O`��@�23��ᯟ�����^8��$�h� <�fAP�a�#������h�'�џ�ᲣI7K�F�(!G�FffQB�:D��{�"D2�8���B��9D�,*��9�T)t��?��!!s�6D�� ��tk]���G�ߔ`�$2D����L�� ��Q��2}o��2w,D��S�g�S�0����@�(�r�H5D*D�4���YF��e =j�L��$%*D�x�d�Û).h�Q��s��|
�!$D���Q��[>(JRo�����/$D�Pa4�;q��pR��~��dQ�C"D� �e,u$^�ص�@����g� D�\@5&όU,�h�x�rxi��:D�p�a�2Y������<:�<�q�3D���ÛRT%�4ID1�B��2D��3�"�z��(�t�҄n�9�2D�|:�'"��H%�
[��4R�-D�8�cH�8r��hQ�,����t*D��p&�0xQ��B��G�6��Hb�d$D���)ڍ ����`癕d>j
?D��9@M�{	
CA�e�V�c��<D��Y�@�+��q!取.E("g:D� �W�		>$vT�sH�13-&=��&7D���2���q�N���/ư����/D��9R/G�xԶ�E�L:R���-/D�d[&�C�̨��C�Os� z@"*D�,PT�,ξ��S���1��p��<D��[�kϕZI��%�0���3q(D�$�1�2�8����p����g'3D��9DdEH/B�k�e<��=ф)>D�)0!��v�yBk�6u�d\R�N8D�D�Α�W��3@,\�2{F�R��+D���f�%pN4q����T�
l�b(D�,H�MG']��]�Hg��]���;D�����a�daa E�:��wB6D� �s��wA��Z��u"�!�P�3D�d�	�)�2%9Ө�r�T-`�1D�� �����Yp�00�.O�nz�ˇ�'x�ٻƀ_,]t�K%��K����*ٽ4�6)�'Ϩ5)�A�wψqVK�\bq{�'�XP� %z���u��(�&�2�'�l}�&��?�RH��%�0��'�e�$�9h��)
4O����'Y�*S`�TXD)�%	�K�,J�'L�e9��B��쵡��I@b�  
�'����n�5�$P���V%@͂e(
�'�r�"d��:�x���08�~9
�'��(��*F���QE��:���'�8�rhH�
*��d�>���'yl
�G�7�D���H��6�~��
�'|�0Z��rTN�a�,�-#h�$	�'�HI�E�%_��ZU�����Z
�'�֠2׃���ȑ�T$8�Yp
�'���Yda@�\�Z�z�z�
�'��A@�は9<��剋�'�r��'=���o��_�I���i�D��'�F�X�D���-��ݦ:6�1�'��Ȣ$��U	^`s�-�27�2�C�'�\9�B��,h�.�,Jpl�'�#@óHt[Q��qݚ�i	�'����աO0��Rl�n�F���'W�I��Թ�.M G皞`��
�'hh
e��.�D+��`J���ʓ�ؠQ�E��6 f� ���/T5֝�ȓt4���?lX`�'CJ(J��4�ȓB��Ÿ�L�(>��]�Z�`��N���cǦ�s��q��֥k�l��7��D O�)�>�Xq�(I�h���pH��SD��:�Ԍ���ԮM�}��YB:A��
6�.�(+�ɄȓM��A���#	b �D 0x��݄ȓ 6�X�G�vGFp��&ޭ$�(��C7n���ι4��4 ǈ�N��=�ȓo�pt3�n�2]�j��f��=�B=�ȓnM�
�u��r�E��|C����h�U 5𶀢v��/tn�l�ȓ�^�A��"g�
С��,Xv�u�ȓwy�IJ��&��Yۦ�\�, �|��mk���,�1�ً���$v�
݆�`�2Dl:�(U��J�JD"D"O�)ر
W3NUh���̊�s8�Y�D"O��Um�;y���A�Q�&�ČHQ"OH�������9�L_�[�d�'"OXdS�5P���H��ԡ��P�"OB��V��^y���I���C"O�t���U�<�P�a�I����(B"O�V�T@tm ��������Q�<i��T�j�|,3c���fTiU�<�g�ֆ��12ⓥ���#�Nt�<!���)@09£�H�`�S�e�s�<)w�K�uL���*M�=	4��b� k�<�Pg�+�hp��D;'L�1���J�<I�m��2AܤɅ��}"�Q!��L�<)��I�:��t�H_4<�C�LLI�<9r��H�xi�R�������r�<aC�����Ú�H�8�po�r�<a3O�e��=��%nX�Qs2��h�<�k�>Z�X|��H�~���%L}�<ɶ�T-.=
���o й��J�}�<a2�ΙK����kˁ��50�aQp�<�w+ۢ6!��c�e81��Г�#�Z�<� �m"��oH�p�TM�o3����"OJ��6�Ą1P�q7L�w�HB"O�-� ���P��Y wLW#>g��H'"O$[s�9y���Ȇ,�=�$�F"O�Q�˴$���ˏ%`��X�"O�1@�o�(M����g�m����"O�ݳ���W�RU'☿�6R5"O
IR���p�D��@���ە"O��f��� h@vEՓs��yS�"O
��
ͱE�Qɤ���S��I��>��	�d�r��?�jG�&vD��c��7|�l�fK8D��R�MH��Z���G���s�Mk�	���[�4�3扮%�`Ef�ƕ\�!��FH������GJ��r�V�C�� �D2����Ɉ�{�jY �/�Ұ?q��>�N�H�AK�myƬy'"�k�'�Z)@1�y{�bH)þ�%>=��	�m���p��9\Ě}á�3T��J � o	�����_�&IA�iO�5v����9\���5�ԟ"~�����<+o���6- �?C�Ie;��p�k���ܙY���3� �A�6�J�� ���p$8�XS�?�=�R��7j����`i@>8L�0�O\8�8�7�#9}�d�1m�E����V�P�*�N�f� �!d�N؟|+A�M�3�P�3$X6�D�c�(ʓ?c�TK�O̕5�H�K��X7�ħ��X��9|0�����@)8�������2&�M���`���<9AK+o�8��a��1F,a������&EƪbU�@�j!�|��Ӝ��C�I��PA�b��~��Q�'(�Γ.bL�(A�L�+:�I��Rn�'TL���㉋5���y�"Z#ԅ��p>���U~I	���x]V�[QcG"1������Dc$��E%��1g&q�81`M�2-tL�y'<ғ9��ÊιS�����TĎ1��"� >x-�D)�fL��y_iAhqY%o֓w��ar%k՚pA���&��W�h!Aw����y��9O`�Ɗ� H�I��A�:PuPe"Ony�5�U�[*�#Q�R��P�&�i��2B�E!|( ��i����$�P�Ax��#�f,��A�bW�z��G>�r4Y��ubXa`dN����3cd�4Ox�!���	*SG�܇��(���'���;��ABB���>J���=���J�'�ZY٥̘=;��)L2�Ӿ[:��u�K��EPթɆn C�I�+L=j�k�!8p�l�ŝN���I��աb��1���M�_T��TJ���Ov>�B�w����j�;Y���2��0,*�'�(����|��(R�˓u#���J҈!I�e�W�&=�	���-=�.�0�df�'k����*Df�L�����>�(ϓDd�X���R��(�x#��>B�"D钉�]���Õ�K�	�"��R��,�֭�u錼�0>A'D97��A�A&]>I�ac{�	�?M���#�9r^X�#C���`��3$��0n��'pz��1�֍^d��S  �X��7�ȬjE�����Qbaơ[[L-3���)P�P��L^�'l�5�02�¤&?��e��͊#J�����Μ�N��l�Kh<yDH�D�.\Rr�M�C��(1�ɰU��	�OC&"���[�h��@��cu�\#G�:p2��D������a+i��C���@��|
ϓ[J3=��i�ꎤ6Ap�UM�\th��X4�0��I��5��0��JD�p�QQ�Y��]�a"��jTN5#���rk|�$�0;� ��vbh�����/���e�2 |9j�FG�|z3+�*H�0f�Ʌ'F����$PJ�<ٰɂ�hEL%�6m��k Ps�G8�> ���0h��p�F4e{`�����`�S5f|n��;Pf��� 0���c#�GEQ�U�ȓ�|���b��BƊ�~z������~���B˃=��l��ink�JG-
-��<���&��x� ŉ6�b���r��8S�b�r���I�$:��Qr͒1�`x��Q?z^l�i1�$��$	�M��>a�F.:
���eDˢ3Ӏ�AABs�iÊ�@aٺ?7~�y�.ϯ��OW~��LJ�: 9ȣhҫ$~��H
�'֨���jS�\�
�;���@����Q
�-�<��u+�?.�d��(���V&z$ �	�u@V�8���G�NB����2͛�$�*���Y y�V6횙A�i��$X�q6�0ϓ)��u�D�+�  ��Q.)�.E��I��tE�GIBf��iX�/�5,(q1a܏U�*���)?D�T��â~��lRG۔^��M�D>ғ ���A1�g�? 2P�3ʺLQ���eԪ�0"O�xB��l�����ϖP4����"O�� '�6����@Mϰ}!�Ր�"O^h)w�\9�����,,A3G"O��i��h$`�@��E�M��"On�xA�N!~�X�����z8��&�����=���OpY:�LY��Ȳ��+>����"O,�"�EVfu���qa]�#���p�i%��B�7Q8�|�痷fĬ�q#F�t%.�Kp����p=���J�e�����:0�᪱-D�M�l D�T�剜�dYn�Ir�6ԚM@�*-�h�65�-M�?��g�, ��	#���0��C�$D���E����HAF�!b���c��|\<A!0-}rOm����!Gi��B@�C:B�"9P���0<�!��Ü=.i1Q�%mt,K7�ڲj�<��B��9D���'�l�Pr�#p�U�P�A�&><�"��PfXݔ'� Ex#�C�L�ͧ:���rD��~��@m�w�����)FP��?A.�˕�
A��)�2��0R��-
\(�O� ��c?�C����p]����V!��� �-�y��N�T�M� GT6 �D�aYA�H�*M��H�sj[P?�'��;;�XqBDe"f�e���q�f6(�U�VP�뉥[Ɩ%Z�`T���$р/{
щC��
�9��O]ݛ�%O�8t�I)P�'���kʏ`�`�V��u�Ѐ2�{�dJ�VdX)[ty2�*�J��O�&�1!L�\�R��f�Z�E@�'I���&K̎ڀU���A�Y.Bk7��o����I��2��<�eaN�Y��,b���=o�9��p�<iG��	��H��ɾr�P�/�6r~���J��!����:cS����	z>G�֥$�����L�y��� �y�͈�oK��{���S�d�EcY�y��J�,�Nly�L�FϠ��%�R�'�@���1mS�aE��b_�#z1���C>6Z!��ɰ�y2K}�@(J��8,�:It��>����J�b�>�H��	�jtƬ���0#"�Ã&�".=�B�I
)�8�q�m��V��|���F������ҡ`�5K�Ȓ!k��h�@�Q�N� ����ȓV�XhɠC,:�ऑ�&���ȓDP:�����I�ܱ��W:8���ȓG8z�¥ ]=DqX|��A�O����ȓ:4�pj�	�u4N|�Cӑ5O�4�ȓX8�����v�
<�v#��X��ȓQX�Ҕ�#�%��ۈ|1�X�ȓ;?z ��Ԋ �Y8�I�-FF@�ȓi�Y�Fnà��s'eԺe4Ȅ�a��b�����S'e̷i�2̄ȓut4I��S<,:� Vg�,g���ȓd��Ԃ���o舲��0/�"\�ȓO�:!藍�HϖY#Ǟ���a��i�mJ�W(Nհ�+�I��_�(��jl��!ŨE��D[GG{re��u�,:d��� �B��Fn_j��Єȓ�\��P"�@�����I�uHX��<����+I�&}��G���ȓ#Ff�	���++c��x�n�U��q��4��s�!̈�T�f-�]��i6�2!���<�Y0�FHz0��],F�!�сg~��M+;T%���zh�d�{B�)@Q�%VhU��M_ʽ"�I� {8H ��>r�����dy�$T�֍��޴!,�	�ȓz~<U�B��<��mRA�,���4��.	�F@�	�� ���M��h��y��F�y�d��'�<�L���c����p`�04~�[��9���ȓ]s�|X���1*k���h�5� <��S�? ��@0ۮl�q �Q�_4^���"OR�IN>���2��N�$
Ri�'"O�]d��%_ض�3�5�\Y�"Oy�w��/$ШV��H�:"OB�Q�%Sr��a(��;"O�1��� ^F�0/�z�"OFݠ���걮XdB�qP"O���⛠?��3���)"O�[c�_o���c��!7��c(D��c�fq��(�b-M/Le�탄N'D�|ppjGoz셰tcȽj���Z�"D���d�Ƭ|V��F��Q}��qv�"D�D	P`�20��Cf�P�vN�CG'D�HRt��z=��1�6)��ą0D����`��jֆu����4!a0D��Rh^=n�Kq��"�R�.D�Pk�+eJ��{ N
+�VհG�-D�H�U�T��p&̔	;�ꔠ�g)D��PQ��	�@hg�.;�) r�$D���E-70,k���B�T��D�"D�4�g��00�xE��a�r$Lm�)#D���4��-�0�2�@�5?^y�e�,D�\ �f��e����`�/IP�ѐ%-D�$9@�A�� �I/��#��!D��8fY���bA�-6��)ږ+D��r�\�e,���&��7?l9�*OF�i�$�6i�Z6T2���"O����m�(u��C.�('��4"OT!3� ;y�����;/B�1"O ��a�3'�� ��m�		���p6"OJ���'ỳ�0U
�Z�ȕ1@"O�@:V���p)U��I����P�"Oh!�授�H
Bᠤ����� "�"O��(wE
�-�H�8u�Z�6	v�8u"O0����rL"9B4.קA�6���"O T!`��R����V����a"O�`�5�pLYP������Y%"O�����B&d=��^F�<��"O��+���8sNz�K�f�=�dy�W"O�����+>nXyz�X��$�"O�@#�ԙ����lx�P��"O���6_Ŝ�*�땳u>X)�"O4�zĎ�X��i�dR�x�(�"O���1K��1@0 �M*{�>x�"O��0B��T��L����rH�@B"O��Z3�U0?ar��Dϕ4 l�"O�8j��F�j��qM�r�Rw"OHx�L��$��w��ua��"OؗU,5��+J,L�q�nM�y�&F�E� ��ÁB9<'����H��y��ޠe f�B�K^+a;�i�"���y�����7h�/`�
٨�� �yb�ɆoC$$�V�`�|���T=�yFF�}kR��2��S��̺Re���yb.��y�:����Vn���A�͢�yB�B(w;�\��
�L@`4Z=�yroKkl`�ҕœ�_�%���,�y��T�n�6M1F��/��5@q�ϥ�y�,W�f��4�C�p��+`��4�yB��[�0��% @�X��l�g M��y2eU�7zd��&.1k�j��C�B��y�j�T�IQ1#ЕX���Se��Py�lW%1y{5��b!F- 1�K�<�r�L�aCpE�gBLA�<� ��0�ȯk��9��`[�WU�{"O�� �!�ek o��J>){d"OI���	I���BD�}7Ty�"O�ܛS��)�<�1%��6 ��21"O��Q̺'�؍��I�!.ls�"O&�����}�lzG�ДH��C"O�Ŏ �0 rd��,��=
��ʂ"Ox�Ӂ��<D�$h ��N55ሙ� "O�y���.��Pd�'��}�B"O�8p�X,/�}�C�?>[�͋V"O ٘3J�E�T� A�\rh�"O\���;h����"�_*XHp<�"O %H�J$T���
ŏ�G�t�1�"O��P�J��K'#Ȏ(�v���>�ƐS��?�J��4S�!I�oۃ'f���У$D�\C�Fr�t��K0A����A�E�I1E���%�3�I��@4)�Nϱ,� HIV�B)N�P����)O�T�à�D�i��1���d.4U�9g�R����P��?F��7������	���1�@BNl�'sfE�D�N�#tD��ħ�qa!@^v楚gAMD��D�'!�H�������˲�F�Lb�8f$b@a��*Wt�H!��O?��7�v�hr҉5l��q3� )u!���M؀c�B�av�"���$�V���8T*��j�f�/'�؟ўh��EQ5>c��VꁸhCȥy��1�O�7fHA�zQ1�/-)u����0�S�E�$#�Z��¢0�O�@�cؔ~�a2!�ch$@�&�4o5�ps"#�r�IrAG�G�/VX#�ƟC���N�=)X�B�	!{��U�&m�p��̊pM&���w�ޗo�hj7HJ.1�l*�S��?�U�^���xQ�.S4"t���Q�M�<b���0˂��+��\���'��(�"���-	v`�Ŭ���O�d��|V��oMQ(P���'@�p�\�>��z ��JLBUi�l�Y�b�8��]�w����,�r\��P*�̊��2��MGz�/~<�+�	)qq���rlӶ'Y��k�Ŏ:-v�E@""Ol�@�Ǚj���AZ����'�|��aV�|�r�` T�"~���Yf��[����{?���2�y@��������D�Y��ٛU�����<�\㗫� Oax���+6�tAƆ�$��)ϲ�p?��
V����eeҢKt�YD����͂�N��_S"C��������"��k� A�"ZP��	,���wl�>j�1�>5C._.�
��)�5,�pi�E"O4��I���E��ȤU���ز�O��w�FO(�եF�L��#y�pp��DC���`�<�A�}�PK��݃�t�
s�J�Qd4�w�`�P�KP�,Wi�M�K?�����SM܁0��*���11�/�ON��ӫ��5�|���Fi��A؄��6iqhM2c�A��b��拙�0>���.p\�����}�"��!NB䧅 ��~t�IҼf`� gDa>�����N���z���4���"=D�$3#�E)$˔�g��AZ�W0&���2;���Q�K������K�OCRѸ�nQ�ԙGZzDz�'^�q�A�wg�ͺ�/�20��|jca�QZ�jO��Ѥ�<Y�a�$��:�Ȏ���q�SQ�<Ir�ٶJ|�``F!�<=V����$5�q��cH���	>^Db�Ec�h'�A+͙ri���d��h��f\�y��N&*����FDG�z����a��/�yR`����#aǃ\^�a�����'.�$�˛v�1D��&Pi��4��f�V�QmQ��y�'�g�.D�s���A�xy*R�_{EQ��T�I�H��ɽ5t�D�҈��a8-�r'ą]G�C�'9��@s�IY�-��S��ä�B�$�4v��� 	� �Z5�nXsЅB��M�"O����H�Z��(R�-mҘEj�"O:��*S+"��;@b�*=�t�q"O���R���SN��}�e"O� ����n*H���o�A�x�b�"Ol�[D	ɠ��@��8 8I�b"O�  v�X��D�,�1`��1�@"O`];���:Z����5̖�ގ8"O���D�O�;dܕ�u�'�����"O��h7���y/���;��ɲ"O2����� e�-Q
IL��l�A"O^����@�(d
���N�D$P"O���1����erf�c�	��"O���`Ⱦ*
 �Ti�VJ�G�N
���=����O����KB�j�*uYQ��J� �ٵ"O:����	��f���,�i�Z���M��t ��p>�D��q��Y�D�|�1��B��8�E�\�dع�0O,�h��W+x�0�*O���"O�]Qq�Y�0\AӓPȄ�����I)g�X�;�,�������r�H��(^�i(� Q�7���8"O t�G�^�cU�5�RN�*9��$�BBA�{���v�>Yve$�gy����������z��,�&@�y�d�3���o��$İb��#M�	I��m����	�q�� H�J=����=LL��?	��	)�4ʓbzP2��]�%����^���H6郍=Ɯ�H��5-�C��$�f����L?�&P�aN���iRɖ����q��&�J�����ͻo3��#r!�$lE��C�FE�G��a��)ɖ�{U�&_d��k�
BQo���̉�W��x�F�y?q��dIڥ�5�3N�jA���D�)�n!`�@
5�े뉲Y��&BL7z���
�j-Jwd�4k��D�`�X�{ܛV_,G�<�v�'�f��gJ��_�x�P��0X4��{R�X )��5SFK�|y�H_`�l�O%��4
N��	� $�����'���M�$TT@�b/�;MR֤��޲&�*YBH��a��<�cl�F�8j=��A��R�<��M��s����&�\�eb-a0������k��ًne�݄��1z���S���SC y�ؾl �����KJS6�	�y�,5��L�ġws�l!6	��y��Ek��ؓ�]�n�����#۠�'D�E���=*6\G��F]����X�a���[Ǥ��yHׁ.�*���ޒX��mr�P�~	�b�@�ɖ�H���f��a�#�ˋR&8��
d%.C�I"M�2���O�1�]{$�T2b�C��@��:`�iƠ�UJ�*�+j� ��U7�ՠ��.'p�e�+Z�[\����_�R���+;�v�;���  ξ��8X���M9"�D%�זR[܉��2Z�3DI\�(MɢB��oφ��&96-K�nI�L�hr�J=WF��ȓ߂\0pkC:�8|Ħ0P%�Ԅ�D�8E�w,��>�H��BǞQ���4�	V��).Q<$YF�v�8؄ȓ�!�e��=K̮U"��L9!�8�ȓ2���'�(aMf5� �2���ȓg!������&Fs`��Oc�X�ȓ..��d��\݀Q��:*a��HP��z�+R�[#����=LȆ�4Wz�Yf �!n��Yyd��?i3R4���b�alWR� �b��5bR���}��ҜT���@�0O��ԅ�I(�$����(�P}A��.�"���y3����D�Rx2ɨ�(B�)	"��ȓf���gC�=�\���Ă$Ix����%:ՊE�5#�lXW�#W~��(dP�E�֋%����Q�
7,�M�ȓ@����eV�f��m��ؿ�����UV`YA�"�=�: {�᜴���ȓw�X�81c��:˨0��VO�ެ��Zu��:P�ЍQ2������!z؇�S�? T�ABa�	g�4m� c���6"ON�Go	�s�Z��Q
X;��<!"O)���Q+��b��2Qh����"O�$r��ݬ��X�u�U�A
��Ip"Ol ��!3\jS�� ��mh"Ob��B�N>K�}���՛y��t�f"Opu '�� �a�Y�9b�a��"OH�P� �y��FJ�\r�S�"O0e��ω�C|�����L,<t�a��'5�vɒ.zN��F��f��+a!O��R�'�T�&'J�	��B8Di�'���q�N�p� ���M��'c���coܖh��;��А��,��'�QP��Χ@�D��"��G�e����
�HعX�L��U�]�xa��pҼ`�hQ��1���B
ue��w0�����ܗL&(Y7꟪+"O�����%�T������$��%s�"O0�",M�K�����F	�p����W"O�y�!l�j*$��D�*w��C1�'66���x�"��M�@���8gp��G�C*��4
@���+H���C�K_�  �&e\9���QQ˖�9e�0�+@����֭���T�j���U�I$pU�v�O9�ա6 
*_4剩>p��G�O�Bxs"��n����Ơ�@m�%�$?��0���C��=E�!	�\������4�ʽQTEЕ'�d�I�~�~E�@���ETY��S�'�H
�۾-��"�1Rx6MZ)@�"pӇ��;�@�9V�A`N���'Llq��''~���*�:l�a��W�l|z�ǉ�J��%��Q��~z'D	<v�h�&��|�<�	3@�wC��k���m�����O4b?}���|i�m����6F�;Kn`ȒG�6݄�I�H�8�y��F,x�ObD�K?񂒌�&��,H�L%:lXb�hP�(��iZш�4̆T���ƥf���IN�q՚�!U��.�d:U$��;|�pG�	�Rt����	&SD�m�ӷ�ģ~���� c��`��Ϗ@D05���#i��	8�hN�:��� T$#K��5���0u�L�ʲ�ԫw�~�X�O�:	[�<RX�\��ˆ"~�B��`�i5z�F� 8����.4D]��WGl�F"D�@�5mڇQ�4A�E7��S�S0Z�P��J[�Nl&�Z!�F�i܎B�	��iu&�;u�8��ˇ�in�B�	 K�.1W��.a���#��%dfB�I0^#�dApA�	k�� X���&9FB�ɐC�	!��ϻ+%�
�A�%O�LB�	�H TБ
��U��q$�L:7� B�ɑv�t�	��@�x�X�&���B䉥8��X���E����)s��C�	C��`χx���h3���?ӦC�-jFv%�Ǡ!��Q�e(�vC�$X���ʝ�jt^��G��*�jC��8�1y��5�V�JB�M�dC�	��.t	�V9�zYy�ȃA�C�"<P����K�X-�Gq˚B��c�*b�N�0����ݳ^�4C�1Q��-r�MK��܉*p�W�`��C�	�e@4x17I��-�`zw� LvB�5u��d�!����/�+�"C�ɘWdv!jD㏑$V�L�p,�C!�B�	%M<�t)F�mm�K��Ie�B�I� ��,xT%�>�4�[W_hp�C�I�-�b�3�� �TGP7>B�I5@� I�,�;k� �B'��<�C�	(3fXa�7�[�o��x�H\D�B�I�|�� ��Iޖ(p�q��^�2#pB��)� M����H����^3V�HB�I?L�����h?QBs0�ܮR4B�< QФ�W�9$"�؂� ٚ��ȓI�vm�G흗"8<u��h�݇ȓ}Hr��`@�(N�U����*M��S�? �Y�#!*,T�x!8g�x��"O���Nv(�%��K��Ze�"OX�D+X�Ifd�ѥ�ClL�@"O��	��}jb|nN+��8k7"O�H�<���TBϲ
AH���"O��²�C+t��c��Ƙ;!��r""O,EU���5�Ƹ�NԜJ�\��"O�y�N�)���ŧ݌|�<�5"Ob�NR+CH)�Qѡu�6-��"O1z���>n�TĄ�2�ԑ#"O�I����{�"1؁#�Gx��z�"O�!2˃�C�(��HP�/qR�e"O*�B
�`�#�YD��"OD 	E���p���v�
act"O&�H�!��x��a3i)rx8���"O&س��M�_�Њ𧆔7m,)�"O�E�s�>�"X˴,O���d"O� y�.Z,��aD-�8=_j)�R"O�"a�b!��%����f*�!�h\>xd��*ݎ�Iu��!򤄔Z�X�S H9E,�	h�B18�!򤛃IiPQ#����#�ࡱe�}!�d7
z%G�+a|�4yC�D $r!�dߏn!�l�w��!uvd`!�$4^!�$[*٤ћ�GJ)X�Lp�c'
�!�d��2`�,e	������`��X�
�'�>d)��32�L U�"BX�M	�'��`��ρ���z�N�p$Ft	�'a�P�����(D�/g�Z�h�'��Q�G�<�xe2�Z���\�	�'����o��\����c؞�
��	�'����� W�,����$vfY��'�n��%�2$tZaa�
m]�-�	�'�#�n���]���L<�
�	�'r�싡d(%�4�'�
֒���'�&��BL0�v]34�J
�\ �'A�����0[�H�*N�BĻ
�'L��)�F�7P �`r�fY�`�rɻ	�'vx�)���'|�ֱҢB��S1ꄣ	�'��E��q��Ar!�*?�Ph�	�'��iˆ�L
�cQ)��:��Y1	�'&��!�+^�`q�$��(1���9�'���j��8IR*$� �@:'D:�'�ذ@GQ�Iۈ����C$���K�'�4Mpu*ʰ~~�<{a��7�D��'x���E�y�>|8Q�P66N���'6p�5!�y-n1p%͎�.Zf�*�'����$o^�"H���C`�+j1(�'	Ze����,�������U��'g�ѓ�-�n6�x�� V{=�9��'�ʳ'�-R��X�@]�^�L�	�'h*X�m�?� H�h�{���q	�'N���b�.��\Hvb�k�9��'@�\:�L�;Y��4R�g��k�:���'�v9ps�]56��!�D�,^��� 	�'�
�xg/��`ܘ�`Ԧ[�`Q��'���M�1eNL@3/,V�"��
�'��k#(J�NWQ:�,R
��2	�'�`5ѤFޠN�\�b$A�y�Z���'>�,���� <JH��ֽ-�Q�'�2�c����ij U ��#|�H݃�'Z�3vZ�_��"PE��\�� c�'FD-��J2
|�J�V$!۪�(�'�b����Ӕ�|���O���<���� Lm���{ �Psh�w9���d"O�HR�.�*U���B��z6�]�$"O�m�"b�6"�f( �.��
���RP"O���f�6�FA�����?�$t�"O�%/�:��Jc���	c
?q�!�$£g{>��J
���`�d��!�䗞2a�Vh��JU(oM��"O@��gW%tP�z��Ȋ^ 98"OZ	�j*,�q!�n��0�~�s"O�iZ3,ӛlW�Aj�"!) L���"O����`
�px1�A�?|9Q�"OBm0G!�Wh��ʂ@>5�"O�)l��'��}!���"{AC�"O��[HJ2��XV�Z�\���3D"O�-Y6!ɴj��t��+��"O�L�R�7��U��B�A; 5z�"O� 83�� pa���O�Y2���s"O8̰e�P�"�� POёc#8��"O���ʁ9}(0�b���5>�ZQ�W"O��x����U�n)ApOM�f��D��"O�9ei��>K�L� וI�| �"Ov]�W��'*r6q ��i/��	"OD��E��Pk� A	x�j�"O6P���*:��ak���!�~�{!"O6`�䪖�3�l��	R�"��� �"O��ZG�K4q*T��}^�k"O0�)uˀC��BI�0F�i�"O��6.�ar�$1�M�6-"��"OXH�"��)$4U�ġ������"O0Ո6JV�#�H�)@`��;mj�CV"O�K�ˋ��Ή�r�H�BA��"Or�0���.i��X�9��B"O�䲐+�ON�@�dЃh�fD�"O��*$��u�n�e�P��v�R3"O�ɨEL�N q�bER;h�&�k"O���%���ZZ�h��_�9;<)�"O��;���.#�e ����K�"OTt90�#��M�2��|Rl��"Ot "#��u]�`����@d>`*b"OH� #�ŦՆ��u-��V�s0"O�����
^Eй��a����"O0RрN4iO�Uc�� OPT�"OXqZ&�޷B�ZA��43<����"OԨ
SYV�d��MN�	��{�"O8� �&Ml���%�P��y�c�#ސ�Yw�L6]����n0�yra���B"QԢ�c�Ӷ�y2�M�rl�x��A�H~*i�&��y���q�|P��K�=l��Ž�y�H��%c:���#�-Ly�03�%�0�yB�կo����'F��A U�X��y2�9��Ĺ��'^�U����5�yb���Ab��=#N�r�5�y�h�"��4K�/,L:̡Gk���yb�;x/��B���tM�%c�#�yro1U���dk�9W�XAId��yn
�O���{��2]����3J��y�㍝2ݪ4)�kE�N�@�	�1�yJ�
�rȈs+ݪof����=�yo��H$ω�3�BP�oW'�ybB�>�N��"��{n����4�y.W�'��Hb���Q���EZ��y�N��	��uф�U>�Z���K��y��|�<H����)nӦ�� T�y
� .y95�2)�œ�]�xP�+g"O
�{r�.@����-����J "On鑠��_�VDi3o^�]�(��"O�tRcMS[� ݚ�N�#�N�6"O U+��Z������W?�`��"Odı0�������W���A����"O��XqfB>(�<�1���#���"O�ɇ���	�()����z�}�2"Ot�k!��&��8��Z4jh��Z�"O`����O�,/"`$�DAL�̐�"O�ȣi-w3t%�	�aE��j�"Ol �Ǜa~ K`�܆X3�mQ"O>�#A��(Z� 2�d�%�uXU"O�A`3e�;:cWZ�d��9�"O6+K�2tP���C) �&���.+D�pK�7Ϫ���;�N ���4D�4�f���vH6=�CO��@~l(wl4D��۔�Q�<� Ȳ���d�Z���4D�l�7gI�	6��yc'��T�>�ڠd3D��AV�L%�A��@��.D�4�-D�L�bMU.s`���A���L1��-D���.�{�z���`ɌG���5n*D��{I��W1��Q�j�3b���x�)D�H��F\ #c@�$�ơ28����e'D���	&8;�툒(��Q�&E(��%D�d�#]�\�d\0�j��Z�L�9D�������H4����;(9�!;U9D�x#V�^4Z���������
+D�dѱ"���s���mu����N(D�b�$Z	-�x\� �q0¦$(D�8�� �hU@1���&|8�M&D�PSo߳(�@�����PM�F�%D�\3�˘:R@|Qʉ
+�&,��.D�  �ʕ�I� ��D�Z���+D� �a �#Ǎ�L��:�Xp�<D�c���4!�7�Z!��ՙ��%D��hV�\�B���ҁ�6=���a�%D�8�b
��<utD�0GM�p�Z��G-"D���e   ��   �  v  �  2  j*  �5  A  nL  �W  �c  �n  zz   �  2�  ��  ڝ   �  j�  ��  ��  @�  ��  0�  ��  ?�  ��  ��  L�  ��  ��  �  f )
  � � :* �0 r8 �A �H sO �U �[ �\  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6�Yg���OFD2�g,dբ�R��T)C>�
�'L$j&�3gO�d��ٮ1v���'].�0�g�l�n��6J��+ᐜ��'��0*���b��& ֏:J��F�($���UHL�]7�Ǥ�6H=�8"F�+LO⟤����o2���C���X��(D��`��̦`�8r,A�V����%�I���O�B�B%��u��]xW�
L����'c,1���C�	1��!�CHN�(�{r�'5��	w0u��z�䗷2�*؈�'#����A$)�dq�@P>�J��'Z~�aQ�×1|u�4�ƈ$e�8�'�^E8�eO��`���j1D���'�8��wg��D�jMNc$z�'V��e��:5A *
�?�� �'[6(�&g;U��9�$E
$2R��K�8E{��t���
�}8G�Jê�9"$O��y�D�F��0Y���4f�릧P��'a{¤ 
%��td@#;uԵS�����y.[�o�9	�ˤb�Υ��[��y2`��2��j�<]��C�_���Oʣ~�a��_�p�ҏЦ4-�G�<ad�����#SpYj��i}B�.�S�O�I)�.I�u0�8t��=8
�'T�h.�jg��#ƙ-f&���'=-��m@0�TJC&@+t��E���hO����o���!�4h��ڸ�䗭kʴ�UJ4D�t" " d�����ѱ0��娷�7?1�y2���	Baȝ3u�;3'��*8mh��'��$^=pb� I"�tbF	�g-�!�� f�a1)	z��R���iی�k��[����H*b�f�cV���ӎd�\3�!��+D T�G��x��`v�,g���׼�(O�>9����U�����本=�f=�#g D��S��������M�4`��H�/2�&�7�Ӻ��[�}!`�H����� ha�<���Ŭ��y��e�&n�2@9���c�<��d�:+��q"�'��j���c�'�?X��T-k>���Cc4A�EL1D��Q�U�o���`�(� �!$}�0�S�'#Z ���}I|�� �J�ȓE��mYU�2l�n���Ù5QN��<�ߓ(�ScF �_��ur���0�F���N��@�.�j������- �}͓M��"~Z���W���À�� r�S/�Ux��Gx�- t�� �A=�!��gD���6�Od�pTe@(\�Ĉ�q�;�>���'vt��8�"��y�fb37ܡ�ȓ�:T�1)Mx�:�"��*K��Ey���n���ïr��J!L�.�Y�$g�
�yRnm��wi��?�P�GN�.$�ў"~Γz��b"ޜ�±�8�����
S��'��E�R�`�ı-���m�ß(��I*���)ρ��XMR"�Dq�B䉮8
�w�U:wRŢBb�t�zC�I���s��6:�n�2Ǩ�-�XC�I�_~�
���#N�.���S?#)C�� 4N2�s�	8U�(�C��8b��dJ�]����c^��~��g M#8f!�d�W��|��Q0��(���$_!�ȾA�8�����VE����p!�D[�<�ތ��A�^0f���Y�Kb!�D�5[6� ���,3/^H�rFҳwB!�d��=� �c�S�(-{�o�m$!�d�d�b���g	�mAam��B�!�H�BCU�=�I2�ԣ#y�%"Ov� �W�T���/O�ysވ*1"OH�J�f��V��� �G���\�a�"OVqd�Ȏ��(�"!ƙSD��{�"O8���KPW���t�P-L�p��"O�bU`5gڸ) �OM<q<jI@�"O԰����8"�Q���h;��s"O`%zvC ld���#m�7z-���"Ovy�7C��Ȅ<:4�[ Bu�ܱg"OD���ƙUE,H�ऌ1d`��آ"O~!@F�gC~�c��ҾU;�#"O0鱠�Xh��-�C݌ \k�"O��k��3b;��*T��;"b��q"O�����̚S��Y�+߭G��|!�"O�J�G^�:�H)x�H �2���v"O�A24�-Tn4�p�&Jw�A�"O�Pk5k� }���H��::clec"O�u����<5�`���@(T�Ƽ�%"O�qE��n7��X�SW ���"O2P�rbH�/Ԑi��:gT�C�"O`��"k�$H�x�%�V�
v��V"O��z� ��q�8Q���%��ij�"O�Tb���?��I�e��Q\)�b"O��p��	d���D�E����"O
 �@�V}�]��"�������"OVx23e�"p,�� �&U-.�j�"O�HS���	V���`���?+���"OnUq�%����
��߫7Î��"OD09� 4����à|�:`�f"O� p�Qe�]����nf� �"O�2�ٖJ������"ON!��C 
FN�)�-P�L��"O�`��$�Z:����NU��Z���"O�bVa
28�V�ɔ��>H�@���'m��'���'I�V>�����ɘ:|��w,S,8����A��u�i�I��������	���ȟ����4��� �I3�F��'��`h�G�4�4��I՟,��ȟ���ş��	�����ğh��8y<�D��o�	�0����oO���������������Iҟh�	��D�ɊGlR����(���ǃD(c5t1������ߟ���ӟx�	ӟ��	ݟ��ɏTN���5�"<D*��[#�^:�'�R�'���'<�'���'��':�[f�ɾS�c���\q>a���'	"�'B�'��'���'�r�'�2Y��I�=IO(	��$�#x� �D�'�"�'U��'r�'Y��'Y��'�B���j��&U`��g�>�rTj5�'�2�'�R�'���'h��'�R�'ל�QS��)��)F�KK�`q��'W��'���'��'���'���'+�4xS �:-(����oZV���'��'��'���'�r�'���'� !�� �7r**�˰�
 L䆍���'r�'�'(�'<��'�R�'� �bI=9�:��33�|�{G�'�B�'jR�'���'���}�`���OV�Q�ݠf��8�mS�J�hH���Jqy��'��)�3?�T�i�l=@�	�7�:� ��
��%c� ǀ�����e�?��<y�K��@����hEN�pV��%C�r����?�!���M��O���jN?��M=4���'�ænd
1��H"��4�'��>ՈP#*����_-@�g@��M뢭^|���OGz7=�<Ց��Yn�����H�CxV�����O�$m�|ק�O���b�iK��K������b�oq�$i�%��.��$i����&[��=�'�?�����j3��ǭD�*,HA9CI��<�.O��O%l�))�b�L� &�)�6dP3F���RE#���t�J�����d���<ѬOt$��Ô62�lK�� �n#v�C���P���c�B�T�1�4��T�v�Mt"�Rfg�*p�����b˥X4����D�O?�I��L�1��2ڨ�a�A�3,H��	��M���ZU~B�g�
���/������P�%Fl�b�L�Z'2�ٟt��՟3E��֦��'Z�ɖ�?�S��{�2�u!�#|:�)  �?��'�i>U��ɟ���̟���(�z��c�ƨ�,P�bj�Ś,�'�6��N���O��4���O�ձc��2
ZިjǠQ(T������VZ}� t�کnڵ���|��'��6�P�z��Ě��G;Z@V�ar�ܴ�	�)M��?�$7�H��( ��uWG&}�fZVy�J�5�����i��.t>h0�@3�b�'���'�O��I��M7c��?�� �B�Ԩ6�UM,\Y�ϋ�?a�i��O��'�Z6mI��[ڴ>����
U�S��s6!�*a2��P��
�Mk�'�"%LdX�����
غ��;G�d������0��%�'T�F���?���?���?����O��|���{\����ڹJa�}�\�@���M��/�|��y���|2#SM��$Sc��U<}�r-�16O8}n��M�'��!۴��$F�,�B��e�ORy�Aʊ
hH`�bW�~�\� ��4���O4�$�O���H�p�m�g�F0!-bu� ���w�'�P���޴��C���?����ڏu5�U�V�J�D�d��,��Ʉ�����U��4~����٫VެZ1h�$)\�:��I�$Ğ�J����v� 6��Yy��u�H��O^�ӼSe�J�!��� 
�6��T�6�)�?���?����?�|)O�1n�=09|x���ܞ3�pX`�+ꝙ�֟��I��M�a�>9'�i�LIz��@���y����h��S��t�6l q2Xtn�<��$B��o�?�'�Dא������R�j�C����M�(O���O��D�O ���O`�'g�u�q��M&��Y6�[�9�����U'���8��ߟ'?=���MϻtIz� #��Ƒ� �A�IK��'�� 4��O/��O$�a�i�d�/��P�%-�<E�rM�`W����M�y�6�{�'����M�,O��D�O*�SA���Z`"@���<<�Ɉ���O��d�O���<��i�F4�0�'���'��̣�,�|�܁
��n92��5��OAy�'�6�.���$���0�@�0OL����޴go�	F%��`5)��r(O�4���,��џ��FEH���i�@�5{�L9�R����	䟜�	�dG���'�
� �F��
��4���\9�5���';p�d�6��'�27�'�i���%Z�9B`�။��1!���U�`�ԑ�4=��!l�����Dy�*�a�6�D����~��ͺ"(
�,�jy��c]���d��i�'|B�'`2�'�R�'W�)*B��1*4`&�?E�4QeV�LyٴT�� B���?i���'�?���7a�
��B��rY�%B�nY!]2�I��M+��i��O1����HǔTjRl�U��2`�pr�I[5
V6�UXy򦓲MƬE���d��'[VH����m��񛲠
=FY*� 
�.o�����"_�AG�s�"\h%bE�'3��4B�!B�a�F�D��O��d�O>��6+x� oW	{�Jl���4$���dp�l�Qk���ŭ?�'?q�=� l,�	[.	�v�3��=��C�6O��D�O&���O ��O�?i#��ȍ@\x�b�Pq��ic�������l��4M���ͧ�?�v�i�'�$3&c�8\�L��v�<#{z�h|r�'��O�V����i��.������T�.+ra�\{?����1��0�I�\��'��)�s��!��̹"<���V,$�\����$����#3��'�V>�£���0`c4���blDt�'�/?�Y����韐0H<�O����t�N��2�C ��lp���[_(18��i����|*r)���$���Z9m̄H[e�ÏY���T�5�\�4G���"��["T=���V�M8�U�iL��?���m���F}b�'D�؀h�X�h�{ �K��~�`E�'�d7MN�`h�7-9?$P,v����~y���-:�B)*%B�{�M�c��y�Z�$��ş �	����˟��Og�Qj&��J�{��	9:HI��p��1c�OT���Oؒ�P���Ħ睾M<2�a�)��
E
���3'�,h�ܴN���"��)T���6Mz�|)�B�C��t�%��'b��䠔b��:�N�[��N�	QyʟDI���?�z�q1�ӺI��h��'y�6����0�d�OV���L`�%2�C�.Q�1����%Tx�(C�OJ���OƓOZ��� <a�U�@�"3�48r����2��+2���nڔ��Re�	˟���-#w���S�E/vHH猉ǟD�	ğ �	ɟ$D���'8ĺ���J�|�@͈�Oc���A�'�6MZ�r��D�O�Xl{�Ӽ����:|�
���U�t $�%'N�<����?i�u/�w7�%?y@��Rs����:X�093�O�1Jm�)P�^!V�M>�*O���O$���O�$�O��S�3�!PnV�
����<�&�i�B��g�'���'����#�(�9M^��0
ί�d�X�#�x}��'0��|����߹V��l�GH�,��i`d(I8c�@�+A�i8�ɡ$ό�
�O
�Of˓1P�Ȋv��P�$
d�2Sa������?����?���|J/O��n�WT����4��dP7�̷o� dd�! �I���M��"A�>����?Ѡ�i��E��<H}t��cT�A��uQ�ɖ�L��F���;�@�yT�t����F��rc ���6�߬p(l��4O2���<"粨H�A��5Qנ�z�V��O���ݦ�0�<B��i��'R&���J\b�%��� ���d"E"���O��4������{Ӫ�(�iC���~�Xr$��[�L��@B?*ߤ��@�ITy2�'�R�'�鄲̌�R �5�����ȃ&y��'%�	6�M�����?��?i,�8�SC+ƺ&zd	Yt�^7{������W}�Gj�x�o�M�)*����V��t�1ʺ`;�ir��ɳ0H�Y���Q�9j��X�|��<���H�[w/�O,'.�p$�9�P�F�$�:����؟H�	���	ߟb>U�'�7mғ9"<�8m�,>`Ձ��sU&|�3��O���_ڦ��?�UW�L�ɬC����gKɖ{8���)O�Ք�����MFV��M�'s��9%O���S������|�Ρ�樉?8�^�: �'G�ļ<q���?����?����?�(�zd��ʨ0�-����9��o��9�s!��,�	���$?%��$�Mϻl�(��]�x��(���9�Ւ��'��7�4���D��RLj�l�	+�I��aA,O�a@���9X���I�[J`Т�'�n�'�d���T�'^$0Q Ɣ:
ɒEF�b�vt١�'���'��_��R�4oJx͒.O�ͩ]�E��R:g��d�a�եW/�⟤[,O��}Ӷl'�`b!�=-�$Y���`m<]0�f!?�hQ��"͊b��s�'�(�Dͳ�?YE��/�,�+G/P��\�ah�/�?���?����?I��I�O&�i$�1^��9��ہwy�9��Ot�o��D	zu����X�4���y��Z�`|��JG�U�,Y�h���y�'i��r�6�iӢuӒ�]�������H4��FR�w�X��#,{���"�F����4����O����O���A�)���勝k���Y��ҧ#
Z�]D�fKU9_���'�R�i[�
�FI�r�#�8�z��ۯ*�<e�'2�i�z�O���O��D���@]`b����H��A��E����S�@���� ������n�O���@�o����5�Q p|�x���?9���?���|�,O�m�`��	]�$�	6N*!/��(�d�I��M�Bb�>��?��d�l� O�m�`�q��ٷ00�����7�M��O����j]&�(�����.7L��U���}��T�#����O$���O8���O:�3��|4�a�@jU5-sh���'E�.�}��ןx�	��M��Ð�|��HF���|���!<h����u��@��7��'5B��D����v���:�
G,Z�$����BiVk��ym�Z���$�ķ<�'�?����?��Α;)���ɉ&h/�a 勩�?a����Dڦ�0��ӟ����� �O$��J�"�_�1��L�4-`�O4l�'�B�'#ɧ�T�'y@A7�U#yX ����4�|���t�vj5�i{�	�?��U�O@�OV�8#/Ԟ*�ub�!]	+(�`���O ���O����O1��˓>�@Ƣ8g�:6L��r�]:��z�0�C�'���}� �䙯O�$��b���bA��.���Ï�L���d�O����o{���I�%��#��<� \8rL�J2�{���P)���s>O�ʓ��=a��tc��Sq�= s��h��
��G�2x.�'���	�զ�h�~�R���<$�!d��xtB��	���'�b>Up�*Tܦ�ϓ�������`��pZ�d\XJ�)��V1`�鬟�'�8�'�R�'^d)�f�O�7�(���E�&�J�a��'���'Z�#ڴ���
��?��g��D���^��X
s'Z5}�H�@��+�>���?IK>�Ej�9q������)�ҹ[pe�K~!^�nm�Լi�1�&���'�"��]�r�p�L?$��iĵXu��'���'���ȟ�5F�/7>�I]�b����	���)۴`�~�s��?aջiN�O���"5�ͱ�b�8DϢ<�6GS&�$�O��$K�]��J���'Z9��hD�?�����L��lIūpJ���\�m�'K�i>��	埼�	ڟ �	 d�&(�G�k�A�/I�D2X��'��7L3{H�ʓ�?qO~B��3�.}Xf,֫E�XKࣞ�u58�[���IꟌ�I<�'�?��'qU�qa���vJ�p���$cNp��E��;?�0��'Ŝ�y%ʈ�t�Ǟ|2Z�4�¤��j�Ia�	l����Eʟ���՟�I˟��ByrE|�j�2��O�`Å��]Cܩ:��ѻk^���#��OTXl�{��7
�Iß4���M��"�2�fM��ЃV�zEѵ��sn��ٴ��$׾j��`�'۸O��j�0H���+dDЪ�;"����y2�'g"�'���'�B�iC�zd�f+�]���"�F�0���O��d�Φe��(|>��	��M�L>)��Y��Q���8�(*������?)��|�U�_�M;�O��qش|@�t�QH@�;�)2�M29Ʀ��7�O��O|��|���?���~07�S�^pQ{�]�/��S��?�/O n�9a�������IW�T�C�J٘�� "Op��= @į���LY}�'��|ʟ`��� �ZBBI�b�_�!����V+V+��1eF~����|:����'�����]ƉhƮ�.��j��W��0�Iϟ|���b>q�'�
7-�0v�x��Ϛ$!�6���g�j�ZG��O������y�?��^�T�	�-;<��%��Y��#L>966q��ڟ�7��妕�'jf1i4͟V�'j7��h7�$z8���T���͓���O���Ot���OX���|2�%_�`����q�����(��g���Z61��'�2����'��6=�>d�񋉏+�RQ�`#1J���`���Ʀ1�ٴP։��O4dp[E�io�R�Ќ��7m˪$h�h��b��d��!Ӏ����\�O���|:��.�ҭJU��$ ~|��$A%w�\PR��?���?�/OX�m�=��4�'A�2v0��2���3�d�4cX"u��O�|�']2�'��'!�i�B�L03C\� ք�%����O��@Ȯ|q�6m:�]���O��J�)l9��K��w��,x���OR���O��D�Oޢ}���-���C�X�n���J'w����@K����'~7�$�i�e	a/��i��-z&�>f2ݩf�c�����۴t*��qش�����\���y1޽)�eP+A�y�O[�S,�0��=�d�<�'�?���?���?)�)M��� /T��#�I,VLQ,OLn��vB`��I��I}��1��X�~��B�@�o�Ik� 
��d�O��D�[�)�S�0���-�!�&��R�z���Z���?ժ����^���Z������ߌY%& ³�^U{�1e'ņtB����Op���O��4�ʓ!I��gٹ!��ʇ�|B�PYD'Y�		a��$��l���m���$�+O��D�l�J�~��7K��]h�`��pE�SO������?���<�����Y~��O'���	��(�	Ң��  �_��y��'�r�'��'���I�<@��E&))ISr,geO9[����O:��M�M@�Ak>��	�M{K>��ǟ�b- �%��2t�a
1���~z�'v�'p�v�)̠"��7q���	<<J��'�P_R���hl�@A,�?Rt�$�@�I~y�O;��'���<(�,�i�~�����B�'��I�M��Z��?I��?i)��3�_�_�P+�L_�[������@�O��l?�M�7�x�O-��ˑ�$�B�w!8��Q��@..�	H��OL�!��O��)��?�B� �ě	o�@��	.@JMPD�ʰ�<��O�D�O���<Aıi�:DcO@�l�5�+��sr�"ƣٷ���'�:6m/�����yӐm�������e��W� �H�j�֦p�4[��9�4�y��'S���ueT�?���O*=��g�N��@(�ē9�|��8O�ʓ�?)��?Y��?�����I�MPjq+M&2�:�s�͉K�HpmZ�
,l���柜�I]�柤����ے ��w{̰bMҺf�x!�vb���?y��%ԉ��O.X�H'�i{�T�K�Fe�`ꁇx�t+&�=~��T�!�4p��`�O6��|*�$���9@ư�0H�����?��?Q(O.Xo�Hm�}�Iß���	S$��G�� P�ŁL���?a�Q�0��ڟp�M<ɴ��v^\xA/8�V��!dAE~^p�vD��F���O�rP�ɂh�	P&N�3`(V0让��'�c���'��'j����H�U�ԭ"reɶOa�]@Zt���̦m(E	��X��%�M���w��l`��v�<�r�nH'XE����'{��'���T!H蛆6O���ܐY��|�π ��8���|\���@L5}��s+>�$�<�|�<y��E�dT�G� 6����N~"�i���"��O��D�O��?�sP��:��9�d`$]�R'�.����O ��R�)�S%������P(I���0DX�0�<��vƛ��	I/O�����L6�~�|2V�\�U
��0�� �h],�r�k'�Op�oZ�C�tL���jJ�TQ`�
���=j�Ȏ-R	j�I�Mk��E�>y��?!��Y�N%��C�m	&L��c	J�MB�J��MS�O"(95�׺��$��t�w���""hÛ�z�@�đ�B^���'���'z��'�2�'���1�ҷZ�t����`N�a1��O*�d�O4@nZ(����	�4��3���G�:օ�2ƌ{��K>����?�'vs�$۴���̦n��P/̺PB�[��^���yC���?�4�Ļ<ͧ�?Y��?��ƕF�t�����]x:��e��?����ڦ�������|�OjX�
Ń�~������}FN�q�On��'&��'8ɧ�)�a%�	t�*~v(��p�ǰVn��T� ����'���Ӆ<�OVE�ɍc	��Yu�O0��\�4��(��ݟ��I��)�Sfy��8��%b�49�f��|R^T��m��U�6��]~}�'ڼ�%�/I�0Хm�ZQ��@��'Pb�N�c����LI���,
q��U�ԍ]0р������i(t2OL˓�?���?����?�����Fݶ[���r�*Mˣ���~T�l�&D�2ԗ'����D�'�D7=�2���ܖ,��$J ���p����'�����ڴ<����Oy�]�w�i��Ē
B�<���Хm�Z%#N����3�0M���;"�O<��|R�2ֺUف�ːH&8�#Ђ�;<'8H���?���?�*Obm5��m�	՟�I�V��ز�C;o����"�����?Y0R�أ�4Vܛ�b'��	l_ !��J�
臢T�F����<H�eL�x��c>%���'��=�	'RH����� D1�iR@��5��1�IߟL�	����b�O��`Y�dx��"B�F"8��O���}�h����O$�d�����?ͻH��q��C�.e��ӥ�9z6E��?Q��?�r���M��Of)�q����4��/�.I��^>- c�3�'�i>!��ΟH��П�		�,kс� \|��g�	# �0H�'T7æhO���O��D!���O��3�"Ĥ��$�' 9��r�y}��'�"�|��Tk(�|"��#E��t�!I��װi ��5�4A��O �O��xP(�jw�!#-�P�/�}�b�A���?a���?���|�/Ov(oZ�.�����n8&��a�Õ\��DЄ�3(�0�I��M���j�>���?y��o4j<p�c\%I���@�I�T�����M��'+��!�j��'��D������o���P膘ǎTّ��b,��O��O�D�O��!�Ӻ;��T��m�	r���i�.�#!@���ş��Ɋ�M���G�|��`�&�|"���&|R6jN#^}�s�C)��'2�'��/N�Rɛ�7O��S� T����Q�v��u�I�
�XP� /�e?�L>�/O<���O*�d�O\��7M˔^��8Ȱj#&��� �O�į<)��i.퓆P����F��,	��	�H�����0*ڃ����e}2�'x|ʟ�� #B^��lW5����@�'"�1�Din�b��|zׄ���$��'�I
2%�����=�l����� ��ƟH����b>�'Ԟ7m�Jx��c��N WD�f����9���O��dȦy�?q�S��`�4^�P)CX�ttۥ��12�ձǵim�6��O��6m ?Ac�N��`�	2��A5F�Z!����=~򵬄��y�^�D���� ������I��@�O�L	���Eu� �!��P�Qp��s��=q�N�O��$�O,�����Pצ��)p�T��f�K;i"����җA���I۟�'�b>ѐQ��̦5�bR�!G���k�1H�J�F�| Γr��y�����0&�`����'�&`�W��"�R$p�J���D���'2�'��^�8iش�<��?1�%�\8BlP�<����� @ ��K�Rd�>9���?�H>��Z!K�8��fY8,��`q�G~±X�{�,�Mӎ�Ԍ�?��x������rD��A�O�i�h�����?9��?����h��Nݚu
=(�D�f���M�x���$[ͦ	Z7,�L�ɫ�M���we���1�6���V�H�'��'��7�U\��6�'?Qv��Y)d���>9� m�N��P���2� ��Fg.y�K>9-O�)�O���OJ�$�O��L�)|���[�I�:>>��{AK�<���i~H����'���'��O���V��Ƣ�0�N�b�JT;���?1ٴQɧb����Vʎ7	tl���^�;T�8&뒎f��� ���G~BL�1�D������'�� <�x�F��u�n�!�J�D�l`�	����	ȟ�i>�'v06�K 7 ����GҐ��w�D*d�z�cׁ�"A���$�����?!2_�t�	� �	�TY�]�t�o�щE��iT� �f�Φq�'j� ��?u�}���%�򍃆�&7�H{`�ҦX�"=ϓ�?���?Q��?Q����O����`OOq暉8e�K+Jz��H�X������M��|���Qћ�|�a�3Yk>��5	.L�z<`4΃�^�'2����N�~=�ƕ�xX�I6� *��@��;b�x�1� #�Fi�&JP?�?q��7�$�<ͧ�?����?��	�k��Å`�;*���:����?9���$馅+�������	֟�O�X��G�@��6��:T���C�O���'5b�'{O���O��24M�1�QB�G5*��\2��)a�(�hC�t��ݕ'���Z?�I>��\M���)��/&vΨ!@�ɵ�?9��?���?�|�+O��mZ�Q�88��X/x`H�&	=E�U��C���I��M��B!�>���v:9q�ʺ-�d�B���W�uk�Λ��[�;/����8pFa��Y7���<ѡ+��[ah	��(;X��yhҠ�<�-Ob���O:���O �d�O��'y�h3d��1#Pc���]�d#e�i5�T�w�'r�'����oz���N�J`;gȘ�#�.���ɟ���6��Ş���ݴ�y�Ƙ�Pȶ��DוZ�r��G�@�y�lۻO[rI�������Op��H����
q������Q��$���D�O����O
�z�����O��ڟl�b�%EH�P�rlݸ#|n!���w��f��	ݟ��I8�ē+v܍��)ڏ!p~�{B�E>T[�a�'A��3�O�:Kޛ��#��\.�~b�'�����H 84�>���o��<�8���'���'���'��>睦[�*�jD��57��5�u�� �`Y�I��M�"b�0�?I��o��6�4�ȜB' �q�*Y��J�fH ���O���z��HlZ7;s��n�q~�FB$���?�R����M�v�Έ8⇝�5᠙|rR��ԟ��Iߟ��I����S�E(_�(X�RdyjӰ��W��<a���'�?aB.@�RX�C��D �C���Iǟm ��S�SL^Dju�\�e 81HJ���y��jϐVcB�S1�tDC�O��O>9,O(K"c,c��`��]�&�!f'�O��$�OR�d�O�i�<���i[Z���'�����.�,U,N�H��\a+T;C�'��7-%�ɸ���_��-C�4Vp���Ҷ'���@ƭI��S�ƙ7��	�мi��I1��؊�O�q�X�΋�*�$���l���ʣ@�	\��Ov���O����OZ��5�,�*iY�/�##mH� �4����	ן����M�ԥ�|��eZ�֔|b��/v0��T�(X DF�&M� ՘xB�'�O�$i�7�i��	)Fܾ�1GL�F �d�������{A�ʆv�"���<����?���?��%
)/��ksȁ5(b��� ��?y����d����"ßx�	ןD�O`ָZ� $h)t�j�ф9�t�h�Oؘ�'�p6@ڦH<�O��(p��{R� {@b0h�"9B�K�/+Pa�$H���4�h���d�J�O(1�F�� :}���1,� ���q��O���Oh�D�O1�
�a��ւ�W���	o�bR�m�42�2�x��'�2�uӪ���OZmnZnB�����`���
DoG�&����ش�4�۴���_ n�R��'���(E���AIj-��GK�uٰ��Ky��'T�'��'7�W>���$v;
���><fx+�%�	�M�!�?���?�K~���M���w���q�>7�Zx�De���b��n�"l���Ş��8��4�yb;MBԴ�"�>�6a!�%�yrDM(�h�����'��i>��I63QVܲďߐ{��(x�H�)x�	��|�IП��'�X7m�	Lw����O���Ӌl�r�ߋ'_��(R�Z�5;2�H�O���O�$�L�A�mg����&]zM��G:?)5+	�3ƶd��Ȩ8ļ����?W��*Ue�A$@��}@�tZ����?����?Y��������,��ޏ'bX ��Н:L}�0�����4/�8����?q´ii�O��Q/3Z�b�5"Z��P+W.O��O��$�Ojd��'~����ҟ%��-\����%���R(	Y�u��# �:`��O���|z���?Y��?i��J�� ��8
X��D�ݢ�-O��mZ�T'8�	���IG�I���c�
,!jv:UC5�Ҋ��d�O��;����g^,ˠ���hXt�*���,��`���uӜ�n�"�����$���'cބ��O4
4\]p�o[�#��a4�'���'������\�`
ߴ����r̢)�����Ty0Cič[���!��NR����S}b�'���'�6�P �5O+�4z�����$�i�mʲ��������4MQ>a�]�=2��R�L�(��Q�*�/+����	���I��I[�'U�� S����V�3�O����Γ�?��)��6�G������A%�d�@߷�BUI]���!E�T�I�<�i>	�ҏ�����'Z:���LRK=���2R$A�0��dŗ?�&������4�j��O��D�,&��U��iۇmj>��m��^j����O�˓F��a�C�r�'"]>��#c;�4����3^��E��m=?A�R�D��ޟ�%��''�D��wᄙ$7.��a.��)�@�{��8f��aQ�4��4�����'?�'8����@�r)La��՛[Ԋ-:��' ��'t����O_剛�M�5�0!h(+ᘸZwN�:���5^���?ٷ�i,�O|��'Lbi�G������z]4У��f���'�l���i��I�%��L�4��^97������̱e�d�zT��e��<���?1���?����?�-�� *��ݠDn��ˎ$HJ��N���k�����I�(%?��	8�M�;[��1P��Ai��!�[�>j���i*�6M�s�)�ӭ\�ְo�<� ��"�ZK�1� a��a1!=O��D2�?�1J0�ľ<ͧ�?��ʑ,4&��b�I�R��%R�l��?����?�����dǦ��@�dyR�'C���b�ҔSh�� OFS�і�Ă{}b�'�b�|�ᘗLFBa@2l�-
��s��Ф��$؂s�u����L�1��q���I�<���FF��$�8JLS��A X�D�Op���O �� �'�?q��|0f�� &?Q�� )��T��?Q��ie����OPo�k�Ӽ�� ��"m��`ϝ�W^�$�#�U�<)��?!�W�(��4��䔗��LK�Ov*X9w��	+P������S�*Tw�|�Q���ş���ʟ���џ��G�'U�v�:�EX�b�d����Xxy��{���97;O����OP���D�gW��G��r�&u�Kܗ�.-�'�2�'�ɧ�O�B4��A) Һ@@�I^�A����l�%]F�F��H��(_:U��d:�Ľ<a0�U�~��ERQ�F���c�_��?���?����?ͧ��D�mR�j����)�kk���<k�
(B��d�@Z޴��'ծ��?Q���?�7'�F�.��G�F�7p^4�W�V�}�n�!�4��^i��9����@`p�
q�f��Am�(O����T?O��D�O����Ov���OP�?�{a��!@)Y� 
HQ����$�	�\��4��Χ�?1ıi��'�R��v/��~�X-8�!Q L�.=�%j5��O�4�r(JAg�F�T��a��䘏\�X�'d�Vl`�S��)BO��$�1����4�>���On�$U9�*QP���8�Ҥ���[.L�f���O�ʓE����<e�R�'b�]>ih��S�=b�L���ǰh���)TN/?��R��������K<�O���a�A A�*�W�^+�P��s+�f��ҿ��4�>���}%h�OT��	 V���b[k�h-{��O��d�O�$�O1���(/�v����NI�#*�1"�Ƿ9gz�9�'�2�|�:⟘دO�����sNB����ʡ;���H�0G?��dTئ)�R�æ9�'��p�ㄐ\*O"�T̙1GP��1�Ο�h�&��3O�˓�?����?q��?�����	44�� �����A��&� 7&�o�!bx�I���IH�'��w6As��L�}ڥ��-O�E�}�a�'�R�|���/H�ț&?O.�Y����sX�X`%J[b&\�1OJ8H�%΅�~"�|rW����L�M�X�ahϮ4�HP���͟�������	Vy�t�6���<��^���%�4*�`�P��f�*l�����>�ѵi7M�U�ɬ�Լyc��m\���R���)d�u��10*�,S��|�pj�O*ؑ�1�D�s���5P�2]B3f+EƸ���?��?Q��h����J����'E��T1<���I�&���d�����Fǟ��I%�M���w���+���}�P#P�_L��l�'�6��Ҧ��ߴs�~�ٴ���|�@-���z�0p����.��
�JZv�7)#�$�<ͧ�?)���?���?a#M]�5�4t�!��ԋ�	�_�ؕ'h7-��gN����O���'���O��hrf^�S��L㗮Mc8���gDH}b�'�b�4��)��uj���E�X�h��xj�m�>#�e
F�+[��	,8-FD�D�'�@'�\�'qT����?��D�է�������'x��',�����T���ٴQ��͑�.�f�Rp�[���B���S����!������e}�,qӌl��M��&�]n�-�D ��Z`J�$v4aPٴ��$U([j�����O��F�o�J�Su��j�<���O��y��'��'���'���i�1mB �HԝKc��*43P���O��W��y0�Df>��	��M�y�Ȟ(B�� ���L�%�4�޽V��'y�7�N��6&�Xo\~j�-`(m�@�תv�y�s�� UM�Y�R��jW�|�W����Iɟd���Ǹ}��|�s��+H?l-8�H�͟��ILyҥo��U�׃�Od�d�O �'&5:�x3�ͯ6~�0����m����'(��=Ǜ��f��&��')�8 ��H�}6�}�C�c�xɑ���p��a�V~�O6��	�-��'�N4	4��@�~�g��x�'�:6-�/��8��aǩB5�TVaF>:��4�u�Ot��G���?�S]���	$IB�����)�L�J��f� A�	�M����M��O�x�������Q�p�3f�6�t}XT��+t}��I�y�Е'���'�2�'��'b���F�i��̣"@�D͊<Vx��4�`�i���?�����'�?�e��y'���NY��b&�/�XP�AԋS���'ɧ�O�sӽic�DA�`��șL!��9��Nb���܌H������VL�O���|
������6f�AȆ���'�6zTʵB��?���?a/O�emڹMX��'#�N�NVb��'�]�p�(S�IG�O@-�'��'�tOJ0'�.x��t!�V�,(�k6��4�BԤeErp���0擡d@��ɟ�P��ӓ_�r���)\]�1	�ܟH�	�������D���'3��#ԁ�;R�f�y�e%/8Ft��'C\7� =���D�O�o�R�ӼsA<,�c�e�#3������<���?qc�iPb�QC�i��I�R����O�H���7Ǭm��=x�h	�&�T�}y�O �'��'h��d�j�qWo�%3�=�ĭőn��ɨ�M;�#���?���?�O~���Y�Ԩ�5*BH�b�B�M���Z�|���M*L>%?!�r� � ��b̑�-��Ԩ�@j��1MV�.�ɀ V�)��'X<&� �'Z�* ��)N/n|d)A�&8b0��'r�'����S����4a��i�p����	��a�B�7Q�&���(P���S}��'B��`Ӵ �wc�$�. �$�!ʮ�����7M'?���.'���) ���Y���?JwĔ�F 3�Q1"av���	����IП��	����5��2T��z��ѡ�>�Cф�!���O� n���꟨�ܴ��ڔ!���U�9��T�V
M-R,1�I>���?ͧ��iIߴ��D�6r�p��5�Z�\�*e��*��b�ϖ,�~B�|r[����P�	����.�"Q�Ui�K�:Yh�`��p�IPy�"g�Xe�<���)�H�R�1��8���y��ѓo��I)����O��$]�)"d��;X� ��@<��QJ��
�C�8}Ǭ�>4n0��D���`��|����$�(ƍN�0�$�s�F%(��'�"�'S��d_�� �4m,p�bW�p �a#זL��5�4�V��?y��9*���ĆM}"�'Ǽ�H"��I��3D�)�jQ*s�'
:7-Ҝ`�P7�2?IЉ�$H���&��L@�� zq�ޅ<�����y�X�$���|�	�����ן��O^>���(S1h��Qa�yB��tӎYy1��O��D�O��?�@�����M�iTqG�XZ�l�0���?��s���O�Eó�i|��5ОL�pb�f5��B�<VT�ɔ''�i@�m/��O���|���n0,�@$�'{��s5�e ����?Q��?�.O��m�'Y���	��4�	-V# qq3.�<b�% �+��-<��?1qT��b�4T{�@0�dG)}�Z�w�1M�|��6B+E���6c.��C��V�b>�c �'���	�j�����0���9�DH�6�*��	ݟ���՟��	O�O��\�u�:�)@-	�Jts�C� r�d��XP�"�Op�$���5�?ͻ,8qKd�C,��%��^���ϓ�?�^��f�6tƛ�����@M*aZ�􈛢K�����`��n!�Ԫ��
Qw�-&�Ж����'S�'��'�Jp)�����@�O��8M��tX��sߴ�X�q���?����'�yr&�&jo�B!q��d�rFP�Y{�i��iSʒO�O}j���fh=���$�@y ��Sx�A�O��𤂔�?q� -���<I`�֞\��ePn�28�� ��#� �?����?���?�'���񦅐�K�@p�E�@��a�$=�`p[A��ğ���4��'r��?�� ��I�G�q����]� Q@څ:^��źiJ��iG�0���ODq�6��֐_�ܐI&NT.	�9r�k[���O����O��d�Oj��6�Syx�{�*
	0��uf#��Ctdd������I��M�4K�|"��0|���|bˍ�De�T��녏mVb@+��,��Ol���O�	T�oD66�#?��F_�n��!C��x`�Ռ���ĺ�&��P%�P�'UR�'<��'�h���G�:�ڀza�
�w^���g�'$�[���4w�fL ���?Q����i��J�<��������u`m��I��d�O����k�)j&d�&��H A*�X�
��/ٚgB~�1"ی�MC�_����6���Jy��K�Q�T���+��`��$�O0���O���<���i�i �.�kN��sY�R� d��������'{�7�3������O�YѴ�ٯ.�8�ӆez�x�N�O��$�t.~7�,?���&���OC�� M.���u�����$�H���Ny��'�B�'bR�'g�[>=z��B�[��X�fOǩw<R5�@�M��Mk��P�?	���?!L~�d��wfU��·/��p
�II�M:C�'���|����رo�6:O��5�դ�p���ɲEr���6OZM:b	�n�§ *,�6CX?����1nE+rHA�@G6w��b�JcD`�BT2G��D��CR�':�@p�L0B��ҧ(B�B����E2�-��&��v��Q�^1#_�Y��_�H�T���U�`�	"~�0Q2e��S\���,�k��B�H+O�H�5@j�����## �W�ڜz��*�[�tl��;K)p�iε|`H��d��=m��ԃՆN��kGV�XZ�3�K�0"�~�����='pf��s��5(�=�b�\�Y;J�a���ݨ�j���i�l���O����*|,>IB�>	��m�$'��<Xm����$�4�����r�rnOn�iV�[�j��D�%5ap0��i�R�'���'�����\>u��۟,�S���-��J�~�����	�'ڐII<1���?�I�?Z�(��<�O�Թ"��O�-��a���!�.؛۴�?�������?Q-O����<���p�ɦd!oX�:�
�¤mZ���ɶK���,�)���F�xv�%d���_��6��+����O�ʓ��*O��RZ4�G�pƚ	��KҲ[쒔�Ծi'�1��!������P�$V�k��(h2d��P���P!T@��o�ğ|�	ߟxs.����D�<����~/; ��,��㞯5�̨u�ؕ�MkO>��D�1���?��?��V�NA�n�x�� �h��o��L��������<�������E�͚*z�	��=��H��q}���4p��'^��'�"V��r�P*<gl�B�)[36pMHFfD��٫O�ʓ�?J>���?)��i}��e�O�	�
�ᧉ��o}�L�����O����O~��Zl��7�b���m'R��D�s�,p�$`H�i�����'�������q�B�[?it�U?cڬI��g�.K!*�s�e�W}b�'�'
剃\�L˭���U�? %��ʅ�dth!�3}�|���i��|�'rM.qOJ���ǭ7T���Q���D��i.B�':�I�8��K��|�D�O"�	��	��i0N�*���#���=S���&���Iӟ�B��\���'����%�P�Aƌ�$g��c��^�0XnZjy�
Y95H�7m�OZ���O��	Py}Zcd�JFN]��Irf��m3Zixܴ�?���)�bM���ȸOF��z�*�@�*5��F� lL��Qܴ*���!�i�r�'x��O����ѣ"a���ע��r�^�+��gۜmo�Jn��?����'�Jh�`�=T�i��C.]֙�GGz�H��Oz����xE�'U�	�|��HO\�C���FD���RWr,�>�b�B̓�?9���?y5n	�	p�8�f�K()J��o�'ě&�'��Q �I�>�(O�d7��ƨx�P�Ԛ`����Tᢍ��T�t0�
e�IɟH�I🠖'�<�1���7��@W�+�HQ���H�Sr�	Пt��֟H%�p��֟X���L:��%�K�[ՊLegC�0�'���Iٟd��yy�d��b�Ӥe5�|�RQ��a`6M�<������?��ZQ�x�'�8�����O�:�ڣFɷ:�4%��O����O���<�D��/x����o�04~jL��eB0gF=����M��䓵?��6r�� �M/r�V뗨�&U�� 3�p�����O˓5��^?1�	���?q�>�jƃb��=��S�2���+K<q��?���J�'��I�_\`���υ_-<R��ރ"<�&R�t!$�Q��M��S?]�I�?e��O���ȫ[��S�d�$^�=+��ib�I⟘�	��ħ�������ː�(�� �2L���x�Bf�V�K�`WܦM��������?M�K<ͧ%_>h��T�{Vp���y��"_��M���?�����S��'��NI�PߪT�������$��KEP6��O�$�O8�WC�i>q��n?��5ws⭓F��/Ȅ�	P�]���	|򉰀�9O���O���m�~4ӑ�R�'~�Ȁ�i�0�����4�?ib��m������'�ɧu7�ԧ��ig��H�X�
ᄅ���?�,O<���O���<�ˌ6�(��-`�J!�"�	��A!4�x��'zr�|�U��ݖ2	�;��J; �	(�.�7��O.�Oh�d�<��*�2-h�O�ĂeJZ-CIx�� )0�
iش�?q����'���'𬬙W�߻�MC����F�{b�%\�Dn@{}"�'�B�'�ɐ,EDL�K|�"/	fm�ӎ\ }�2�� -�G��F�'z�'��ɆrʆY��M�	�'k�ZFi��-������`����'���ş�+��SJ��'��5F�����g�xB��cŔ��ē�?y��@D�����B�S��A|�T�QB#L�v������[��D�O�DA��O����O����R�Ӻ�`ʀ�RHP��LԺKo(���.���I�H"2hɺL�$b�b?��Q��x�d�2@]�^�ܹ�ab�np�ס�Ӧ��ןl���?�`J<�'kuB�2��<PQ��R�+{Z��ƾim�U���'zr�'�B�O���}�䋑�V7��8*���pf�N�6m�Ov���O�Y�ɣ<�O�'���y@� >��r.�J� 5�u��4����~2���~R���I��̇+C��QT�E7�M;� ��(O��Ok�O�-`v��+�4�fi/{�f�0�r}2Kny�3$�S~��'�2�'2�	�{��$`��ȱ{|��y`o�-t��(� N��ē�?������d�B�� ���G�՚,�l�C4.ݷ8} �$,�$�O�ʓ�?q�%�8���(g8@Q	0▉.8�]��.D>�M��?9���'f�L��f�q�4%�Dr&��7/b���C'W�4o@��'T��'�R�ԺC��ħP��YY��K�_M�uС)�	D�1X4�i���';��,�I�`�TX��h�i�4$'��
6j� }�C6E�3����'��I��LZR���'����5�$H�v\ʨ�V+׸0�|C������?9���ش�#a�f�S��b�l�j�b�71|�	�,��MK-Oh�C�G�ئ�����	�?)	�O��A.h�
"M�4,"HbG�߈I��6�'@���D�<��� ^�t���`�"�{� A����M��M�3|O�v�'X��'T���>�*Oj�c��v,��)�6Hw��@�ܦ�!��g���ry2���O��9�n�''u`�hA�Ŭ�Z%��F�٦��	Ο��IO�h"�O`��?I�'�y��a�Oq4|�T" #Zn��ڴ�?1*Ol$Ȥ4O��ɟ<����|�0�L޺��v[�D>"<a �C��Mc�:��e��X��'"T���i�	�Q�̦e���i$ӎ"���$��>A��O�<���?a���?�+���D~�C���GI�="ti˓l�<	��gq}�]���	jy��'Z��'G]�2�9O,t	�o	��G&-X\)̓�?A���?����?A)O��Z�I��|" X�S�� �\���,�HT��\���}y��'tB�'�JQ`�'��|
��ѻ\�0�!�&/qI~Y	6�>���?����$��"E��O9��ъc9�Ͱ���7}i�|�(V�eR7�O�ʓ�?����?�q�H�<9,��fBQ1}Ɣ`IbG�/����$�M��?1*O�Dڰ�E~���'���O����� ��lΔ!x&d�x����>y���?���e�Y���9O�ӾM��� ���!EN@8d��,^Ю6m�<�D���?~���'���'�t��>�{�? �jj�#Ppqb�.w.�@�i���'���"�'���?i���▾F�ce��{�2=A�H��M�˅�$��v�'GR�'����>y*O�7-�f��a��$D�g`��H�ş3�M!�<!���?����O�򁙽$O��B�
��#�ɋ0�A4
6-�OD���Oъ3��A}�Z����w?A�1�B,3@S�3#�|aAJ�����	HyES��yʟF��Ox�ć"#	{ (ǧ,�Ru�(��	{��l���bEFX����<�����Ok��oƦVQ�f���`R�]_�.�l�ҟ�9�{���Iş���ԟ,��yy�޵Yv�C��
�ͫ�	*0H�#
�>9/O��D�<1���?�����z-߫wRʵ���Լt[������<I/O��D�O���<I�Ɨ�_��2}\"�#�(ňP���9@�D�&_� �	Ey2�'e�'Sr٘�'�@h�H΃~�r�I�£-ظ`BP̫>���?1���ā(�P�O��Hw��H�U���6�ɋ���h��6��O�˓�?���?�F"��<���~B�s~��Ej��oh�������M���?�(O��I�y���'���O,�q�O�Q����1�X)b�3g`�>)��?���>�L��?���?)�Og��[WKΦqZ,�Հ��@@��4��$L���nϟ����D�������<�@��u-�)�S�Re�M�p�i��'n`���'n��<ы��
*N6����n��i2�I�U�ֻ�M��jA>m���'���'��$��>�,O qr��(%0�p�Z�?���P���uCq�h�H�	Ty2���O��
��][�']�F8�ۀ�Bܦ=�I؟��	'g&����O�ʓ�?��'�NP��덀<BPh%��(5��xش�?(O�3d6O�S˟��I��@12�.�ϛ�k ���͔ʦ��Y^���O\��?�)O^���.\��!�q�J)��0�$9�Q[�h��ez���IΟ�I埄��Oy��+S����D�m0�:gnAHeja:�F�>�)O�d�<����?)��e�r����L��Y�劌|:�I~��'���'��Y�d�qCЃ���<<�8d�W���Q8��)��M�/O>���<���?���B�@�~x�%p6CF1a
�QhЧj޾ ⑾i�"�'x��'=�	�q��}3��l��ٌ6>�Y  � 8m0�1�
��^���l��\�'���'�aG��y2�>9����9�\�`e_V7R-��oΦ��I̟�'�t��Ơ�~���?I�'zn����NͺS�.�!��H9E'|�ʓT���I�,�	�]�����'z���1n�`V�A���e�0�։%Y��S�HS�5�M����?i��b1S���d�t�A�N,��ȓOF���7�Ob��'Y���O4���O2�>�1d��D��Q�#�3T�F�P�oӞ�J�h������������?MK�O��W�� H����J ����< �iV�	ʞ'RP�������M".����p�G�ʙ^�Q��i��'����JO�듑��O���*A�.�ȃ�#pX��U	�+mf7�3�d��h��?%�Iɟ4���IvX�[�(ض�C� �\I����M��E�,}��R� �'�bT�$�i�y0Tbʅ'B�d��"D�Z�s5a�>o�\~"�' ��'~Q���++�h�p� 'Q]�e�o�=m�P�J<����?)J>���?�$ҟi-�����c��AUb�rY�,�����O���O��$gX5h�5�!�� �,�陖�Z��H��U�p����$�t��쟼r�fq���n�d�d�z�bϣ1�N�yd������O`��O�$T�9�����/�z��d�Ȏ(�3G�1d6��O.�O���O���'�O��'��`�u�W�^���#�Q%u��;�4�?�����D�KV��&>Q�	�?!⥅�uS��rˊ%6n�^=�ē�?�^�N�s��������L�P��5�ϯ�x������M+)O�����J������B�D��\Y�'�T���  Z�䰳7*��/G�S޴�?	���m�����OμQ�+�QŊ%��n���|�ܴXa~�y�i7��'��OWFc�@�Ƃ�y(�H�(t��Y��Γ��M����?1M>Q��4�'$^PsZ�k!�2y�
��4��7q6m�O���O���6�C��?	�'V�ٕ B$Lz�
U�P�6P���4��6=)�5��d�'I��'sv�RE�	"\�v��g�ѿ$�*��	p� �Dk�<5&���ܟ<&��X�!�`yADO�vF�@�.�=	���p�@}J����O��$�O�˓5��U��I_L���@���H��&�r��Of��>�D�Od�d�	5D�`Wm�J��\�r �pKƶ~;1O~���O�D�<����-m�󩟅b�"iI�,.��󋙛?��	ß��I[yB�'��'׌(���'ƈQ��� y�fԱG���HB-��>����?I���d'��y'>�*�f�X�8�9׬��
�����/�M�����?�� +�������I721��A�T#�M\OH6m�Oh�d�<�2H�~��O�2�O2�H��R���!�.Ä7����J#�d�Ol�$�L�$4���?=�`�9�4�L@R!$���cӮʓF�\���i�:�'�?i�'��(��`G&Rq@�A��<5 f7��O���ذ,�8�$$� �S��T:`�5��ЉJ*�v7��?�o��p�����S�ē�?��%ö �X �qAN�0�PT��
(-����I�R;�O �'���Ob����53W�]�A!֟"�� DA]��Q������ɫO,H0�}��'�� ��p1��/8��SY�@y�S�i+�'��#��5���Od�d�O^̸��I�[7d�褯��A !�eeP�5��w��(L<ͧ�(O�b����0V�el0L���x2�'��ݟL������'p��� �K^�3C͗�X��� B �_��O��$,��~�"D�r�1�`-�E���C�J�M������O*���OL�`�|U��<�VȣMT��vԂ�J�-,X.�x�Z��It�'��	ߟ�ж�J�R`ܡ��	6J�T�jbH�����O����O:�lI�4�q��D���]]ԅ�ЭK�-�H��ӄK6fB�6�#ړ��$�O<�O�@8R֠��j]��5�֤'8"���4�?����d��"�$'>I���?��g�Ra���J�2�Ywi�>�c�X�'����,�ISr � !�e��^�\7��O�dG, �H��O �d�O��ɦ<��!��W�?Gs
�@�hV�TTn�ß��'M����/�j��E��v� ���˚�M��U����'��'��dl�>I(��P#��\
h6`1���0�p$ۦ��	C�'�' r+���� .�2��y�T̙�9?�6m�O����OZ����<	/�������{G��I�:!�2��a���dR�Of�%>��I�t�I}R�Wi�6cƠ��+�wX���ڴ�?�`]��d�U�4�'*�'����aB� o���"�+b5d,*B�*��?(;�Iǟ���ȟД'��D���б�Z�Q��c�Ze�BD��>���?)���?ьB�$}��E@8B�Y�m��a#n6m:��O��d�O��$�O��,�?EI��#2٢��+���(&I�H���O��$6���O�ʓ6\Ynڷ(��!�IB��B�B�/��
��6��X�&L#���(��0��*+O��JE�/� "O�ܩ��Nf��Ag�G�8S���g�O0t"3�L;(;���r��?$eΐ��O"8���cr"�&C�L#�d
�v�x�1���Q�|��#�?�����E)�2}p&H�� �� ��V�����m��8頪%3�p� N��ыAڡCCЁ)猙\"H���@X��C�K�h�h�[�W�Hu�򋗺t$����'J�'�2�A*��4�n�9�	�`��[6.I.��H�-�u�L�	��D�_��@�'ۘϿ�ѤP4n�JYcч,S
��
w�L�ԕ��m��!�;F�P�G�((�!b]4X݈�z�����;��R�Kё@��r+ ��(���IШ�?�������T�|R�����q��ꕸIc�D�蝸�y�fJ,M����s�΍��p �ے�Oj�Dzʟf ���z�hS ]�zi��0u�Oz�d�0�T���Ot��OV�D]����?1dA�k����EX�p	ti�-o����TRv�`U��MR6骰ԟў� ��b0��/�6�B�CW��?�����{���P2bJ�$V��3���k��7|ɤ�Ȗ�������_��a�����D{rS�8��.F�WϞpZ&��Uw�a�e�7D��  �+v_B��𩀊C�v����W��HO��oyB&��H/6mկ|��ū���s�$PCf�M�H�D�d�O&�D�O��@��O<�d~>eJU�O^�DؕE<, �RD�� I~��N]�|�.ߠ��d�/E#��b�׽%5�T�2�+&��|Bi˴�?��.�	3j�1)Ү�Á�ǌt�\����?�*O���?�)��b�(�v�"t��eb@)נ|�<�D�+Ts��('�I�ʉ��(�<9�X�ܖ',E�U��>�����I��3��I�@̑+АP��@��#�tx�,�O���O$�AAlJ�@�>Ѹ�����gd�O�Ӱ7?�DjN�D��C����6���<�qM�* Q��[L]&t��zO|:A�Ʒa�`�Zm�4+;�H$*�d�'�$M:���?ɋ�D�E�6XB!Ϫ[ X��fi���?Y���;r�}�T(*�@1	c��BI<yD̄;CD�3�����h�+�<�CMİ���'�BY>�є
͟`������	��4�|5�%&l��4�4��%�~�K���Lp��%�O,�'���<�a+���#n�og��!%Ь�D�)ߤR�б��>E��_*Փ��N(n�.�84�O�
��ir��R=�?�������#|�	�JM*��D�ѷ D �3�ɬ�4�̟dG{r���Y]���V��0*�m�#�M��L ݴt�f��5n���Ѱ��RmO/\.�Q����ɤa�s"�Rݟ��Iş����u��'�"A*�}�oœl����7��p|����_�V���Xr4U	��hO�dQ�GP�V�r$��܀�ҵn�ϟ���K�h@�
Ѱ!���I�*_X��6d�@�~8IV�z���	�#C��$+|O6l��LǄ+.����W6�>�#"O��A�͟UY����BF���	Cc���Ps���ܦ9�%��Y|pT���K�B��}Z�L��������ɹaB01��ܟ��'k�dU�%F��eR~Ȱ	C3�}����5kenxi #Q<�〉
ϓB���#a���r�`�G �i�� .@a���0*��9� .��������$n/�sǄ�� ,8פT֟H��{y��'G�O�3� X�q�+L�l�&��;Q���"O��+0��g��U!���A�0O$\o��P�''�Y�1�z�����O��'J1�������Hn�A��k0�c�eߟ�?���?y�'O-�����Ņ~c��S��Θ�t�z��	/�2q�D�Ϯ�(O^L��I��U����%�Qܧ%��Y�k�'��a�"S,"�Dy��?���?i���I�%E��)Tƞ ,$�Ҕ�Vc ��D:�)��<YA�׵]�ʌ9���3�
�k�cN<���3@�����K w��Q�K�d̓�?�y�J��g�)�����о1- ���'޼��pX/D�����. $h�{�'�v]������d)�h|� �3�'�>�ʷDT�5�Hw��!n&�!��'>���4�j<^ii�f^�g��1�
�'����U�Z<��넇�+2hf��	�'ΆiPF�2LӸԺ�oٻ#,f@�'�\ ��&�A�pa���3Pe��'ŀ4��K�LB��d$�Y�d4��';>��WF[:�����G[���
�'�)БbO�{;yhCG�A'���'���"C�^�`	�3F�>,�MI	�'��рU�Q(U��S�P4.}����'�� �j��P`KB>�~���!;D�p0#�ǣ�$p��y�$=�S;D�4 u�ɲ>1�H�rB��V�ģ>D���i�M�����&�T2F��e!D� �ub!"���cۯ=,p���3D���+�w�$T�X)�� �2D�dn�&��2��זR�y���/D�(p�hƺT$X��-�:Vp�u$#D�0ɤ���~�1���J8y<A�C�+D�$0�L	2�����ꓱj4��W�)D�$�S퉎xh�����+�*�)L;D�h��ʙ�:����Z�-�
���,/D��CI�rDP�ȗ�c�:<Ѕ�,D�\��"Ȩ�:A.���8��+D�j�o�3)VT����Q
#��8wj(D����ݱI��	�@	K�[��h�`	,D�X��6݈"�G��^����W�(D����T ~�� )�3r�`��%D��"P�!/�a*�B�E�IPN1D�da�C�|H��h��A�JJ�Xr`0D�@H����2�� (U��I�|ّů/�Ol��E�Ɵ<�D	�H����E��@]q�-D�4��Fǉ���	"�N9A�0��bJ,�5����"�'2�Lͣ�%�H븩��S�9���Q�T��#�ò��F�c�<-�I�;J(���S��:����#[�l��0G��H�v���%&v�ز.�c<n���{`^�<pF��!�a{)]*�ȸ��Ӄ^�������>�d���7�W U�� HEO
��})sHV1!��۩%�X X�؈oF\�3Ŝ�$
ў��j�' �>�q�hΦpv�����F�uؤdq��#D���i�9�����ßxN�(7b����d�d!�g?��j��-b�)��)۸=�����Cd�<� �L�Z����AZΤ��A�ǟ���5�O�����56Z�R����Aq��'(.QZH�d �*�`���P5%��X�B�)D������3��b��U@�4�Tj(�	�"�Z#<��T$���V���:��G q+.ūu"O�� *%.��0�(�%#�p-�"B ��OT�}��q��i?(��1�eH�'�L�ȓW�t}9��֓*���Q��.U�4��ɕw |��d�.~���Et����JՑI�a|Ro/�$/Q�r���R"_q���@��Z!!�� *ċ�ަ#sh�c��5y�� �"O�MYѯ�z�1��m���U� "O��	�?W:�L�4a#"OnA��ÖS�z��Q xt�dB`"Of�A��+MعC��V"tr�9�"O�D��BN|;�qh� �"O,YSa�W
KF(Y�dB��k���e"OV��	�
��egE5(> �Ӥ"O�<�#�0
S�\���UL��!"Oj�V�
�#u�ѱFf��b>���"OZU �A'\,h�#S�!;�1��"OL��p�ٛO|��@�F�-?�-3A"Ox�@�R/�<�ˀ<+ ��"O�I���2�hQ!��D����"O]�3�	$mT�(�s�ԄZT���P"O���䥔�}�D���B���b�"O�I����$~@����6	�U����� ����X��+F�^�8��Dr��Dh�"OJxP'hP/hnp�$	�v����E��_1��|�'��p f��-� �#�i۔���'�\����?3����E�8/��!p��Թ5����D>{0,�2�,�]��Q����z��zBh���E����i��K�t���H�8;����\��� c%>AR0�#!�	u���=���>��O�O��S�`��S`<�t�al�I�'�:��I�خU�cc!Z�܍��R���'�V�G�,O��I��:I�`��(��H�d"OԤ�&��o�*x8R�M��XMM�i��q�6�'v(��D���$���ȡi�=0��'�x�h�E~��ͦ%1��Ku��$�������yB)�U��M�Q��s1��04��'Hn8Z@�s>!�ba� � H�]y��{�C�	?5�
�/�/d���P���el��Cу;��02qQ>���!��>���4�Q�d0贅ȓk6X Tb�Ds�0���M���#�F-6�����͓v`ߠİIq@E[h���5dB<�OH��"C�0[G����ח4��`�"OL�:�`_cl��2D��!>I����ʏ��t#ç ����E$h��ӭUi\ؙ��W\@a�%�?$��W�U�%��0E4.�"��GZ���ҟўd(�D�*�\��H��ab��8�OnA�p+�~j*|� �2�0'd�2�F��M���Va~��-�0���.�8���@ U��O�(�cYZ�A`��<��@��P��Y%c�>u�3��D�tC�	#T�"�x�-J�t�r�(����^��0@� B�gY���!Ny��9O
@k�(�2&�D�h����9�"O� j�䏞0�&�¦Ϛ1<p�(�����ʤX�xQ��Z�G��3�Y��lصHU!`�H�Apˋ1vK�ԇ�	�ތ�Y���5��	��'\�~��ĸQ��s�"��㝒:�B���'����ټ"����؃UO~��y��ȣO~��@�/&
�h�#@��=Y�\>��� 3]��j��Z�|� �#e/:�O�D��%� �(�d�v�U��$�7�-�����f�C*��x��bòB�̣|Γ"u.�����d�zѺCF�+�-G|R�ޅPT �dB��O�ީ�"
�e �@)�a®EK�ㅺ."��[ �`T�� �B�����DR:�p�pg��n8�`Ӂ���)78��� �6֧��i@�m96���P��h�q��.@Q�j���4k��xg��!F�'�r��ˎ�T��=�v��)cvzs�%G�I"ͳ.���0ڴA�<�)��-u���z����sF���4�0���l�&�<	k1�Lo�h8���'Rh9��

K`H���J�e�L����X����r4O,D�'Gjm����#����g-�R��<��l;;;|�¢F���"�K�y�'���`co�����ʐ��a���*��#`m@G��}k��_�C
�����BV��r�'|�Q�ψOR��sh�#dM�ᓷ퇁tEѥ=O�9@��9[~J$HG4�1�1ODMC
Q�7�@��w�H&a�t DL�t �z��
Et����;I���AAM��wo�1�Tl��H��L**BԽ�S�禽�4�� �	v��<5�7��!�8cW�'��)gX�^2%�%!�mԂA����s;����-C���I�NU��ٵ%$�)�S��V�#�Ѭ- ���B׸$��#>it�Ǌ�$4����v_T�O4��Ӂ���M�X�Ȁn
	���bC�\ܓ�X�G��O�<��M�de���4�][1ָ"s>O��JR�Z3�4�k�r�q��T>E����yc�t�W�.A5.�AS�V�O�)�3�'�8��B��?>�V����<�̍`���*l����fU�{��÷U�֝���禙�:�	
�O�l"~�R�ᗤ&��K��'?$4C�oN:ʳ
@.n��c c�Z]`��6N�����m�hu�uo�A��� ���a��?�I�ҝ���)�Hjg�ķ,%�#<����t�ޤ9ы�=xҀ��Ƙ��S�'Ti3V��l�01�����~�xF��#E����\��8��w>#>�5DZ�Q�FU���?t~0@�Ɉ�ä��gD%�<�A��#D�)�)�L>�a�l�gD�|�B�)0i��gPYr��Vi��T���+NZ�8S�� �J��M�yzn��Ũs��V�!��?1(����;7m�@5!P���O�`p�"	x�|�k�W����2�-Cp��jr�U�7��5JF1�ؓO�4HB#qz��0 f7^�y��~�=ݬ�H�]0�H�{�p�Dx�h_��X˕
�� ������?�'{t8�d��-�=ѳ�ů�j=�4�2�-ӗg�6��QhF�'"��F}�dϦ	���K�Kp5���N�mX�hX?*1�ѹ�G�Y�~�����L���޺C#
SN B�A��s)VIH,Lt"0�㠉0�O���q)Z��q ��~t��R�)�?\�"<�'��	=6T|̻7~���S52��@�7G�p���	/r�:���?~7@�O�;�����[^�q��'"P܁c�>�s� y�v�i�,����#��$�b�H9:0���u B�z5�G�Peў��C��j'i�P<^���/��<p�J# &`Kk�TƶA��.�O�0 f*�T1�hCad�m�<r��I�0P�eZ�S�,�|��7!Ό1��I��:�����
<����Y�p��">$E�����â����� �C��x� )�O��y�3��BŇ�>�~9��
��7a�9�E��K�����$�y��T5{Ij�:�,�wp�ܱvnF'��?!��D;��b#Ș�$���ND��������31�p�N�Q�8�n����	�OZ��NP�g��a�K8���$�����A�2l��=胶0�2�:b�ܦD��8��i8e���V!��c��lHP"��N�Q"�M8�l�f��+�Y��ҵ0�v�p��>}�\�+�p�r�Q�X���U�8(aSUA߷s�\�[sǒ8=@0І�V(<�#j�F��BBY�T#����D�x"fQ�dl��.,�EI5J:扜n��6��\�r&z��8�O;F�μ����Pd�B�J8�Ot�dJy�h�g��9�������?2�
��6�&˓��u�Ol���-�'ϸO����.ͰO�x%��%�y.��c�����wrj�d��%�Ր���� �Թs`RrH�<�����Єvd��{���p<�Q'�n&"�1�ꜿ0O6�� ,S䟰��"[}��L& "���Y��*񪇵v#f��`� �O�@%�ÝR/zCቛP!H�C
_�"1����*!���:1䀰5(3?q�'�䁲I>��{]E���>�
=���W�	"�B䉌:E|�*�B�����b���!l���W�<4��I?+���q�k�Xp�\#4Ƅ�
x C�	 uT�I8G+Ӵ/� У#�M��B�ɞ�ѻt�6j����s���B�	;`��:%��'x(=�/�%2�B�I
A����#Jg��(z���	$�B�	�¦8���
�|�,�,z�C�I�I$�)Y4�@I��Y&�C�I�
\Q�w�L�M�M��d�1��B�I�RA~�H�� �����k��B��~&�§L�?�1JGĥO�C�	�XX���l��O^��cT�sF�C��0 hL��Q��,[�@E�L��C�I�L�n	;td���a�	��1�) �'��R��U�7��x��=O�X��'��[�E��n���ɖN�})�m��'+�x���z��'LP.����'¶U3��Ր=�N�����?y�HX�'�|$��N�!� ���Gx}��3�'��s��ܓA7܈�iǴ�E��'#tLcRU�Mǰ��#�S�z�̠��� ����0u9��M
J�X�7"Oڭ�ǉ�����
HD�5"OjdqF���)�l�3'�J�:� 0"O�̲���i9�k��~jXPA"O��+��!M���g^�@�"O�d�Ӏ�[��\�b�� ��$��"O��	�+V�|�"��U�th�t"O�5�N ,8�����&"O����^6:���� �ԡE�tE["O��vf��=��0'��SR~��p"O���T��uȡ5e��kU����"O�-dQوl�D��JT@��"O����V�C��:,+���q�"O��{��:g�`�R�j��c��;�!�dɦ>�$9G.�%����FS��!�dn�X�k�B�x.��#�7v�!�䃒i�Z��ҥ�,�Cb���!���VJ	��S K�((&cU�yP!�d	�˔������J���0l�yB!�DX?��$N��):B���cm���ȓj���lٙq?��sl�l�J��ȓ=�N|�GL�g�Z]!�Ɖ(*�
���R�V��j�.x�ep���<)�v��ȓZU��7��J�Re�"�ݻD^���A2��!K��&Z�Eh�-4���ȓ�Taa��#fF����؂]�� ���<���yb|�ca�Ž:	^��ȓp'X�{���J<|{�nعs�d���8k�h�"Ǎ��=��cֵ%�ȓ4Fތ�G��(&AL���y�b�ȓH��܀��+LQЩ�$��){k
����xRu'�>mcJa�*�[����mӺ`16�,7��'K��Zw���>�P��i�4|����&Ήćȓ;����D U�q���x���(��D��_��="g)�9�5���L�g��Ɇȓ0����߫20f�2!% p��ȓ
^�AW	S�4���2��]��e��^"Q���5����a�9C�~t��DQZ���T�T�h(��%�8G	D��I-l��5M�&i�\�a�T�:IvфȓPMޡ�4��{�f�y�A\�C�L ��p޸̫!@Î^�x�Ԍ^BULن�>��@�%�8� c��ϒ5C0D���4�`��q�Ţ�P�*D�p+R��<ph2P 0���kB ��&D��2��������A.w<T�F�%D���j�C���9d�ޗ�B�{�#D��ʢ)�x��e�%%�X�3��!D�<[D,�%j����mZ�<�&����>D����aا"�����DQ_Fq��-)D��i0��T�����[ 9��L��k(D�@�&VN`�f͍gk�Hy M%D�苳&D�]:n=�f���+v��R�6D��!�	؁nu,b4H*+Qv��4D��Q晕l�@�:���a:��%D��x�S>kN;b
�$i��R�!D�`{��A�NA��)�& V��I��,D�pzF�-`�Y��/pӔ��$%)D��Z�,�&�f\�e�lU�\��'�1O0yXv/Q�c�ʶ�8^?mЄOcp�B�9��$б��3�\4�W-0D��f���:�i6�-g���t�.D�LGK��ʆt�w@��&�Т�?D�� �e���+�m˒��wV���"O����?�,)e��>I
0��@"O��`��Ϸ(�Jyk��G�(��iXA"O}�"�R���ƕj�|$�"O�`[7H�'I��o�L���"OДa��*-Uą�gN�=n���"O�Q D�*"K>T���P��x���"O��Ӫ�2����ڟ7�PA�E"On�)��c]�y�� 
��� s�"O~q�E�hր��q�$7t��"O"�"w�6�Ѥ�_:�%"O�]�Ũ��yQ�%J�3���"O�y�&f� A�"�# =5�����"O��Q�o�"7+į3܀i���y���'' x�,Q]�� ؜J�����LP0�6�mN4G�$=�,U���Rr/�(t�R�����<�@�B7D���G7 n��eM=gB�iB�a)D��ȵ�_ jҜd�tf�j��8k�2D���#
��̀��E�r�f/<D�l�b�Z���(��L	3EJș��9D����ힹa��L2cˇ'4�D뤍7D�d�`��7vɚ�ˊ��4i���3D� �Ql�	�U���0��#�E&D�4�Á	*��`��ŀZǸ�@6�"D����)��y�7M�L�r ӑ% D��;�B��
$�m�%(�>���'?D�x �� o ����JB:z}ڠ��:D���1�ȹ%���iG[�h�Ьa��"D��34�іTj����-\�%:��+C�!D���3!�0����X`~���� D��c�C'\L�#��3ж�Y��1D�@s�
%"���qT�D�I���#�B2D�t�3�W�(l�#c�����Hi0D�t�֭�6	F�U��&�!@겕�T�*D��2��@�{�N���j�(}����*D�LQg�v���zT�C�4Y��PѢ=D����n��Aw
b}A�n_/d�!���Z�ƀ�g!��+��@Q����I!�$P@lp��W-�L)S����6�!�D˛����ƃ��p��iA�F�s+!�d ?7\������{�pTR�/ȣB!�D�0S� bO�=������!�$ .�q��]8"���K�!�@�m��i�jφ-4 �C�K�e��}◟L�0�ͯ]@� ��!A�4yd�1D�T���[h�(0�e�,&��q('4D��{ H�<k��)!з�}*�B1D�|��
�
vfU	S�Чw�n��2�,D����IF/D�~�JF�5H��	�,D�4A�b�O�`	@a�'	���'?}2�'Mn��P�K�c��l$�У#ߚB����D�S"����/�qf]����!��ĥxي�����GQ|�qpB`�!�dW�(#6�M�4hڱq�%Z	w�!�d����[u��e���$��!�W�X�����8Ni.�J�dD$;�!�D��E�rx��`I�	N(e�¢��`�!�$Pd���AS�Ш1?
��뙫]�!��*nF���Ъo/p�3��2{z!�䓲t��	��MjMPhR �A5 =!�D�5]����U	b|$��#:!��;��M[��Ϊ(�\a��E9!��:���Q"�U4&1�CʍP!�� �8F�UFH��z��ӯz��5Z�"O�rPt"�Q1�`� "O�0��]6A��b��;B��=7"O�� j֭\�H�3�M��N4˔"Or���o? ؔ�BڑQ��
�"O���� � P��j�a�"f��hR`�d7�S�S	:$@�CaC�nXH��	��x�~B�ɟ(�i���F�|u�$HO�30B�I�=�&��r
�w�0�(Ϡ[M�C�I�1T�@�!԰r4 EN:.�C�ɢ�����iB-(c�E�M%�B� (=8fG
>u��5!�Dٿ��C�ɸ:W1{� �8K�Ak���9�0B�ɎBǐUwj!��kם=�B�d���y�l�+R�z��A��)�C��n��)�7N���UF��p�C�MǺYs*h!AU��r-�C�"#�����T"4Ah����ZB�� b$���ڀ�n1�d���^�����:��I"^ ����z 6��� #]��B�	�*����`OQ 0��,�b���@�C�I�k��������X����%(�2C�	=(��(��6�8��'���B�ɪst����=pp��ţ{>�B�	�v؉����tM�Dca�&=�B�	6X?�d*]:@|P�6	�.��C䉠.����I[��5�0�N���C�	;$�+�ݐ�0�-п3t��'�0�3wb�&=3�UA�O��<�Z���'�B=��`�[$N�p��[�>��{�'�v��@�2};`4)QO��$�@���'�D X!��'l��e�'ČP<DI�'`n(x���y�����[�5�8���'aTs��>�0c���E�'I��#��&�XS"� w�,���'��1	���;f��!¢[ k��9��'-�	x�Փ\@���aA�%]je	�'T�s!�<{�!H���jPJ�';P)A$C��TT`�Q��3#����'�x��呺#^2h�.����|�	�'���R����A��}C�7��!��'��0�%ݴo��$���0wMv���'���Qg�C7fOƴ�Bd�>t�Ft�'�|�hǇ
�1���j����C�ٚ�'�(�S��O�DY{�8��=0�'7�d�ͅv$�� ��-�:�'J��R&!Nq���Q�V�����'��z�M��i�>\2R��JU�D�'q�9I&L�/M���ڑ C�JF]��'��a#ڍa�ʡD
�S&���'.H ���ܷ)6� �;Sp4���'
D숖 Z�5,Ҙ��ʝB|
 ��'�����b�R,�']�D�'������j�:��c��S�x�'�KQo�@xd�!%�J ����'�pݻ�
�O���y�(̐*ͪ-"�'i��QC�B|P '��%���i
�'^�����
FY,�@r��9$&b�r�'�m+�D�!	�!�	R�ٓ�'�������~��♝2"D)�',���HY�G�X �M�
i�f͋�'�^-�'�>���BcĐn���'J��9AH�;��0���_W���'�ЕZ@ᓚ(����*/e����� � ��%�%u������t[. ��"O@$�G�X6V�VLW�Y"4I�ԓ7"O��C�oW�O��<��ڂy(��0"O)1�(�����G��B���"O��#��6�<	�5�]�m�4���"O�I��AĚ,���b�*��:o> e"O�j#��l���c	, za��"O��a1K�.Li���۝pf4(J"O��Qv����&�/=}���"OJ��s`�Q��J0$Ӆk�}!7"O�	u�_�R��ɒ��b�p�"O�M���]$�J��%AC;)@���"O������� B�B_+fm�7"O��3��R�}��W��^"��b�"O��C�
uNY��-��N�
<�p"OP�*���5S��@���n�у"OZ����X>qR����~�n�p�"O�(S���"��1aT���!q"OP�y�LƤAMa��=5�E�3"OV�B�	%W��ղs�.M��e�"Ol�� �R�~�	���L@cR"O����Q�v#�P8��y@�*t"O����l�%8x�V�O�deεq�"O��KC�W/����a	}Q�რ"OH��1g�V���#D��Q�yҕ"OFm"�SR>�0�-+GM�cq"OX��ԡ�,���s%�єyC��G"O�;SaD�xt	)A��('=> �U"O�Qu�ڽH}(-J�N �X��M��"O�(���Wbܐ���D�\^1b"O�-���1orXq�lA�+�F�K�"O)�# �:V�*0�t��#G�eˣ"OvYhf��,W{��RD�	�+ބ-��"O�H:�i�4�Na���,{2�!��"O:�9� ьF�m��+��'���"O(²�֋ܺ��*�!r��3"OBɘe��
\R�C�)�
�T	�"O�A�R	5�����M�N���"O��	# B�yO�9i�M�5|y8(5"O�p�@�M2V�6�yE��pN�(�"O"��bZ�[@� /����k"O̙xՀO4c� ���c�^�u"O�e*�&G�U<�˕AS�Nl��c"O��1!��"i���SG^=[�1:�"O �1�<
�`� �P�y��Xq"O�Q�p���X��KA�\q�"O��Q#��h��T�M* �h=��"O^�c�	 �]��@��V4��@�"OXQ�,���Е:7��
X̐��"ODК��҂o�\A���T���"O��ʠĆ�,0tu�W�p9��� "O&��tP?w	�(�G��RÄXQ1"O�YS�픾xe*� elJ.˲�a�"O�iV�؀g���#ػ ��*"Oh��К���R�n�;hX>1""OXݚ�e΅;\|� /��jjLŪ$"OV����
�d��m3�nǝɒ��Q"O�0��ڤsJ�B�[O�꼂�"O��Y҄@fTɳ�oS�g��"O�5���׵Ilxu(H�{�\���"O<tY�K�L�TE�ԦK� �1�"O�@��K�V&v��U#E�E�f�X�"O���Q�r�Pc���B��I�"O �p�ǠB^�����H��"O� �h sA���H��G�w��� "Ol�ұ��51@PEA��T�[���8�"O�%iq�!4c�������S�B��"O���woȠI��U��G�!P_D��T"O^)jq��#����E��N�fQbd"O��*$��	��1e֠4��Q""O֜f�ĵ�t鲦Ƀ0P��V"O� *2�&��˲�֤R����"Ol���ңAU�\B��2� xJ"O�1K�&��� �(��	^�H8r"Oj䑰D�WV6eʔ�Qsm���"OZ�`Ɖ��-�L�֚5O���"OΙ�5
љR��� �0\�H�r"Op���� b����ρ�w�D��b"O,H D$�0o��,*EIU)m�}�7"O�\� �G��9S�PK��;�"O&�S�dN'�=�U�J��2�"O<�;R�W�o��9� �� Z���w"O:a+���M�1�D�Q�U"���D"OD��T:	ߔ��7�èVs��"Oxu t�׍ �
F�ݭ3���1�"O�	s�b� b�BC��6���"O\P��j9q�p5��'.>N��W"O�* 䞚F�:E���*)Zt�Hc"O�Q$�)T�,-�=R�8Q"O�ИvBб'��E�̅�*4 �!�"O���Ձ��R�M" !� �C"O��&NO�l��N²$0��"O�hzBi��l���z$�A�b�2K�"O��3��$<�hV��#�p24"O��CQ��>r!n�ڑ��S` "O�p�w �����H��~py��"O��a���6�-�����X��T�"O��1A����`H!�W�A�y:�"O�\��$� ���2�쇂<+��5"O>�1p��0V'@�aj��m#Du"Op5��$ZI���c���<��"O���S��z^Ƚ�w%�&%H�j�"Onѫ�-�I��%��0k�ޕ;f"OXD�əvA��z*O��tJ"OQ6��>v�~81J�**S�eQ"OfT�(� 6Hp�"h��h��"O�q���S�*լ��t�C<��<9@"O�htdT�vz,�A�$$��Jg"O��۰Ӡ<�.!�G;s.a"O%z�4^��K٭4a� �"O���7�J=��h+H%^&�1"O�DB�#͛����iA=:���"O*l��$�4:n�X��˲���*�"Oz`��)�y���BԀ�V�~��"O�	
ߟoI
�Q�.�;���"O����d�!Apj�8P͗eG�I�"O�Ӌ[$^9xpLfA���"O��
1A��� �iM�$�<�Y"Ox1�f��,!�]�ahH� �v�C�"O|QBաבt�q@��	�E��m�"Oz�IV��3EF4P����%���y�c�>)%����Id�����	��y��z�p!���O�sb�9ۡ��y�ֽP�*�Ba�i�>%*���-�y���(�ԥA�Ֆgo���`Î6�y�bP�D~=���	�"�Yw��yrc��F�D��@nL"�ʧ���yҮ!V.���(ڒV�f�ڑ ԰�y
� �EH�K HX< qJ�1�W"OT�z4�Q'��I��1y�"O���L�XƔ��u(��.�D�r"O�m�I�2I�.��2�V�򐥪�"O�(;��T�%j���pf�y�~�X�"O����D���A��&?���#6"O�ВE?}pyy���w�ZI��"ObKD#^��4����C
e���1f"O�Y� �C�V�X=I6
W�*up�Z�"O�TRR�\04�b5�3�C7�pp`"O������bmC�ɔ
��(�"Oh�l��[� ͱ��H-�0�S"On����<~�'�*h�y�"O����͐�y���TG��#���U"O> �/OF�<�� ���ZRmX�"O�Svn�WU�s�_�e�Ҡ"O�\�wΓ@����`i!b�[�"O�u�d��.S^	�%�,���Su"Ob�R�FF����Λ06��AV"Oz�C㨇$rظ$h�/S44�T��"O�@���ܝ.G�L�d�vB�9�"O�<@���Ċ�зc �.S��g"OD���݀53��(��ʚ���b"O �����&#��u�BBXs-�YV"O�y!eV�H2�iT�K������.LOm{���8�� �`(HT`l×"O<�HS`ϛ�q�ձi=��"O�ْ��A�}���` �#�"�"O2��"'X� m��;�fd�"O����GU1Cy� L%tzu��"OX1�0`V?�X-@A�� ]lD���"O2Eзm�,~��X����Fp����"O��TI pl	h0��=^�8��|��i>��'���$w�(U�ш��w���p�'¡3t�[�Ea̩9$d�^�4�
�'\�@2�lC�f6��t��PJ���	�'h���µKҘ�QGI�=1�-�'�:�k���+E�}@���4_���9�'��D���û,l �+�'PUc�'�l�h�L&��]�t$[�+�,���Y�j�L��1�V�F��Q�t����'�a~K˅a�"��cE"�ې�޽�y���p���p���;u��r� ��yr!��[s�I����~�zd�GΗ�y�Vv>\�k�ɵM1�II�kC$�y"�w�A����Hƈ ����y��S~���b5�| JJF����O`���$��JDI�BB&k)���u�t�!�F�P��]�d�WQL1+䁍�q�!�d<Ў��͵/��d8V �*
�!����R�viI�1#�4=�d/!p{!�$_�t\��$o��>�Ԉ�UO2{�}��!��N��5���ܪz�QH�?�	x��\J��xU�=����|���j!��П\F�� ߷U.�	)TQ�Q�y��f�3-!���54ˢ1z�F
�D|�}�A@�!���;C���W�R�}�H@1H͑z�!�+e�9��^�j�AC���!��U7j���b�'eŊ ��/������?E�DG��TP�(�ʎ,���t�V)�y��4�~� Q��B���m��y2J�I~Q�B�H _�K6>�y��R)o�z�`��Vh��l>�yba�l�6���
�����I^�y
� �\	��6o㜹X��*"�(l��"O�����ؽ��a�O�Z�REh1W��G{��)e����?�a�j!zM�{��G:Q����JF�ƨ)�R�$fJ�M���x��L+��P��U�Z�&h�q';D�롄�*j\9
�(��!L�����:D�D�2�%4��q�tO4H���j9D���� #'�ri^�3#�A��g*D������;)�J�s�}z���(��m���ӷqq:�� Lo�a2�hB0����2��k��[3>�̺�`քsX{��6�OL�wܺ%;ED�1+���C��V�\70���!���B�a7:nD�QhٴUB0��ȓgjn�{Sj�$Z!d�*T��+�0F��S0-"�ap���H�0!`%�I�p-C�ɭD\���#D�<DV�p��kڒO��=�}�RK`���V�
!T�Q�D��d��)����m��r��$сl�g�>���E��8S��Ă�Vx�֧&IL��� �:p��{V~i���ܥ0��ņ�'d#�m�5�j�GL��U�4��ȓ�b��e�49a�"qj
�[�T�ȓy'��l�Q�QRNF�eGZ��'ў�|Z�+��x�dѰ枚#nH�[���۟��� �\T
��I�~�d�a��� T:xh�'�R�'p�Oq��Q�]�#��BU�N�D��@�$"O��i2��Y�Е۷����tI�"OpHɒd_�)�� ��;ߜ�)�"O$u��ü�+K�5Mj%d�TQ�<�4� !gq�ZT�X/P]��Y�bAJ�	}���Od����L��`�-�'*ۊl(�'�r� ��V�����Ȑ�YW" I>9�'�Z�AY[�Xp�����8n��ȓe�@4��;|�a�&@���v+H(ABB����A��"[i��ȓg�3�*šGK�(�,[�=?���ȓ3�@��H�v㲄�fN$.��ȓ>.b�CRF�*p#|8��)�A%�ȓ1��Bf�����Tb�&�:Y���K~�N+l&Q	�-A�c�p<X�I��y��]a\��FÒ�r
)�(Ð�ynBz�=B������x��	޿�y��G$EI��`۳�E����y�mO,QUΠ@J���a9Ɔ9�y�'(!l|��FJ�{v�5[EE3�yAK�r0@��՜�E��N�y�ς)���#-��`��ȩ�yBiǶKU:U9�%C%a~�D��y2%I
O��
�fQ�-��Qj!��y�[sZX��$/.+�@!Fl���y�g��Pa�,�u�"(j�D��$-�y���7��� #�3&X�U걃P��yB���Hm`���G��(�8�`�y�X�<�5�����
�����A�<���>X�� GSDN`�-C]�<��+߽���
2g�*ߞ<�Ao�\�<���͟	��rAŔ�?���Z�<�����#�ȉ[�@��;V�i�W�I|�<Y0�U�)�dPr��Lq`y���N�<A D�19�h����^# i�4i')_V�<��`�?Q���j���CH�x�<�/s�z�34�}38��A��q�<�&
-=�Yy�Ss�(٨S��X�<	q��3�@e��W ��p j�T��0=� �4�ь���d��hI�v�i�"O�7�,oE.p:@�SC94��"Or���Ƞ��0�L�5V�8t�A�$1�S��<
𺶢�+o��m�.�PP!��y�l��	GSLx1�Q/ԭ:!�$�
jZ�SEg�,e9�urr�t,!�� �)F$����hѺ��c��K+�O���ă�c� �&p�(�O�&j!�$�s�	FƄ�Pj�H�ęs�!��|"��Qc�&:����cT"!򄄆%����&�+t�08�#B#'K!�D6v��PdU!9K�m�ThX�'�!����9�m�?MA�����j��y"቙,@`��4Aܢ�f(�m��"��C䉍S�*�{��-+�u�� 
I9$B��2<�0�g�B(��4heL�&WcB�	�W�j,��@�o���[wkH/Y��l��	�B|���3��	֚x��Lʏ,�C�I�HBZ8�ȡ_n��!ꆠk�B䉴:Y���(�ƕ������۞�y�M�-��ɛ!C�;`v�l�WO�y���oD�mb���h�n��֬���y�@��cN�"^%ޘ`��Z��yB�ϵQHl�'e
�@�~Q�g�,�y�.PT�`�ӟ1�(q����yr�e����&]�����6�y�*�?�pï|H�[��؈�yĉ8�4�zR�A4)��B���y'Z�(�E(�j6e��� >�y��N�}٦����2�Dsg���y�園;�D��dbS&�޵h��A��y��͐�}z�+�=!��H�l�yb+N�G4F�k����F�8q���R��y���aL��Y���`���]�yDEqN�k#
>5��xD�L����=�O��Ƣ��bTQ&m�K[��f"O�)�1-L�O��)��T <��p1"O|���	�(R�0�D �(:�e��.�S���T�~|z���]��0�%M�
(e!��.K��ي�mإYӘ�����!J!��4BؾdH�-~� ��E
En�!�������H�W��c&I��9yB�|b�'<��1����@�H���v吜I����c���	��c8���6-\�CM*��s�?D��j� ��p�����ǡc�X-jp0D������$;�� 0DFS�r�N���.D���7M D��KR���R��XwC.D����-�#u�,aAc��]�h�Z�/D���DK����
�6�:�s�/<O�"<Y� G>��5JG�F���C GP�<�QL�mڔ�5;Zd���s�<) ��δP�l�w�:`��!R[h<�wZ����F+u~��r!�5�ym��/�����>`݈��2O���yR��S��)a�O�"X{<1�0�O��y�
Ɖ(9<I+`�Q�����L��y�eņh��QbהBȚ�{���5�y�=�v� $苢1ni�&��y�M!{�F����J�.�|�����y�m]�_Xv�v�I4*�L����y��ΉP����%��
�� ��  2�yr�X!d$��`*²PXT���I�%�y��=�l T��H�A�
H��yr�\����uhAWB}Zriؒ�y
� ���Wa������J�+�x�s"O�QR�ճm�$�"�(�d�2	Y�"O�:��)©�u�	�L��=��"O�-�w�.��,⧍.>�$��B"Ov�r�R1�z94�ǫ��q0"O6�`��ٝX(f؀@�T���@�"O�7���8���r'�^Q愹�"O6�k!!� /J*����(�~ѻ�"O��١��.!��6n܋bM��#"O�0�%�(21Z�$��,m�1"OP���c�8x�  vM���P�c"O4�+@��	`��Z�*W��b�SW"On�x&��&u�Р�#c#�ĺ�"O�'L�U�ԙ`��*?4 ˅�'�1On0�'˃&�j����5�p�"O��#PA�-�T��*ۻ>��Dq�"O ͱe�"G�����`h hB�|��'Պ�#C�)�As폒+B���'����U썄�
C@�*%[6�{�'�l9�I�X��\S�
^���'e�%e$+QF��q@-&��x��O"�Qt"O�4�F�SvE(oh��"O�	v
_ Fp�S5��O�� Q"Oʈ�څ-T����D�k\H��"O�;���%'�.�Y��Z�B[�A�"OZi8#���|!!���(ܞ��"OBA��ț�L���<w�X�;�"O(��AQ�[/,���e�k��u2Q����B�S�Ol�Y�uF��J`H�
A>x��J �$.�Sܧa����rF߈Y���W�U�h�VT�?���~j5���_�*x5Q�Uf�I�/Dt��H� ����(��H�(=n��2�6D�����Y�H�F�&cBq#/D��T)
8(.uBw�ø#}&�ye�.D���1^�`�{S'�R��$��a�<ɌB��L�c��X�y�"ė!\�$�OB����O�a0��6|,}��;s6Pҷ�|��)�S-�԰8�J+ZP�$��˽o���$9�@y㈗K(�kW�+9�`��,D����(��l�F<@�dV�0)Ҭ(D����@J�kh��*7 H%d�Mhs%,ړ�0|Zc����4��čY���!L�Z�'"����4��H\4�J$��(o�˓�?����i\h�pkT�
;"H3lީ[/L���O.�$#�OИU�S=ZC� ��`X!)�n$aՑ|��'=az�c�9~>i��C�I�>]��څ�yB�@�8|h5Kh��9d�aaQkг�y��f�Ș(��%5Y�u��#��<Q��ݩS��Bγ*�N��b�/}y!�D�q�篆�"p =Q�� �dx���>"�t�AD�# �$��ሏK����?q�ju�4��uQ,5�T��x�P��ȓVʖ�H�gQ�~���D�E�<L��<���Ð��(���+�$ڎ�ȓ#���A䃺:p�x�7�ީa����s�xap��M&7�<=����_n�)�� ��݀!0�%h�hC-9�6��/O�=E��Ě�a%�h��ʏ1DB �F,_�Z���'��~B�z�J�;eI�
A)���Ă`�<1���0{ �81���ucʜ��g�<yjP�y`Dha�JH7"�&L�e�<1��UlL�AI��2 1�s�]^�<y�\���jE�D�tЕj"l	C�<1�,�(M=#�o�^�F��T�|�<� f\C�fM�60�`�H�f�<pKqO�q�F�d*)	�ꎎW��i��)�OZC�	�(��m��C��<O�|��"2�B�i��x�k��#�Zu�7%V�T�8�	�'&B%#DH&�&l���GS�mJ�2�)��"¦=�&�̉�,D&ٚ�힛�yrB�L"<I�#!V�N�zj�fƼ�y�!B4(6��Y���7�hy��g����x�o	�B�9G�ƫxP8y3��R(G�!��+h��x!G�)E�ph�FN�
�!�DԆ �r�p@g�n��@ �{�'"OFu�vʌ+`�0Qڶ��~	��U�|�)�!w~�|h�j�5M��M�];1�C䉘~�TTXe��ma���B㙌���0��	%�i���M�>�)�I/|�C��A2��vE�7�.�z Bt�C�ɢ{0��GR
-9��j9L9�B�I����T��-����&�6��B䉋#�H����^t7��o/��D'�S�O$z�)�֯)���AA�O����Ig�O����\�c3�Kr���
�'ɴ܋/�.��Q�N�s[��
�'�f��'�.(�`7"ҍl˔��	�'zT\r��<^���P����kB���'Q�`B��7H��i���'Pc�i��'BN9kŁ�P@z��τI��4��'����,��p�j��������OX�17�4P
�˟��A"O,��O	,��0�dL�̝3G"O��&��5A���� #O=�f)	Q"O�(X�";FtB Zq�\�����"O@	@�Zc� �B�e�&���"O�U�`�&rk�D���	1?2Ԑ�"O"�37�_�r
��;c�[6'� MK�"O���ꖄF/�I8��P�i�Xe�"O:aH$Ă3t���I�㍍)�"� 1"O��ig�[��h��u��*}�0���"O���b,J�[^,�0��F_��u�"Oj���A�SwҘXV�P�U܆Q9�"OV!sF��`���8F��ܽ*��|��'t�-Y�A� l��n|��+
�'�^��1X!I&�H�G�5v��	�'��ڑʓ?� t��ԯ3����'���"��-X��z'�EZ�'�V��r`��t����q���T:]8�'H���0eָx,�q���K�r|���'ީ��A�r
xp�p��?y-O���D�
-~���ǎu��u�C�B�>�!��ڞl4̣CGW"t{S ?�!�X!���!��H�W6hN�<z"O� `��V�R֊쳤�[B��P��"Ot �,l����Z��m{"O�]X�^n��		��G1�5y�"O��0��@8U�� u�D.;��R6"O�H����$�rP�$�/J��m#v"Orp��O{�L�Ղ�8l��p!"O<��6

#
.�S���T�t`�"Ozdj�I��	��Ѹ�3E�n�@c"O�-)fi��r0҂�K3#��V"OB9H�"� b�Ġap�Y�z&��2"O�|1q�<&����"Ȧ 0�q"Ot��Ī��+��h��]�0T��"O D!�@D�H�����֋- �!�"O�3�A�m7���3����"O� ��s4���)�d1�"n2Ҽ�W"O����9 eĸF�wȼ"�"O:̨e�B�8�0��"�k$"OJ�+��,>MpY"֠*(.}�4"O���ݑ{�
i�O�;|��W*O� $'�$b�R���!�v��)C�'��TE��1(_��a�E�~����'u�xQd�����^�"���'�R���$�2ph���*�'d={T��|,���'L�D+\�h�'^nP��> ���Kj3���'��AU-M�2f@0�ʂ�8��(��'_2Q�N��X|�����<c��(SK>y�u>D�1��L�tCԡ*V#]��X��_��+��7	k�A"q+H%}Фp�ȓ/�I6ᚹ|���y#�� 茝�ȓ|l#!@�_�h�D���EK���ppxM0@�Y-s?�ӄ�\v4��N����&�z��[�����g��T��乲	-D�����vQ�M�˃tg)y &D�����E��KC.�.>��)"D�dc�o]0�����F�\��IIvj>D���7�� L�d�*�@�XŬ�vg;D���юX�XIT	�Ba@��*��7D���̇t�l 6A�3���H��5��0<���0�ʔड��z1[�f�<A4/ȆF�"�j�ș�1)�X(�b�<�S̴nr`40����zʽ��e�`�<!L��mKб��n �tRg��c�<�/��Oe��x�e`�ʀH�<�ëP�V!��@��}�b|�O�C�<��͟'�r� �mT�R��}�	ʟ|�?�}�D�HY)Ӧ� >n��7%^�<�&�jzz����|�d�Q	�A�<a$_�	 `���^�U=x��J�z�<�B��	9��mڵF�� EDEQ#��w�<�,Kd����0nK.���P�HSw�<��H��~,��b�޵2��}� �q�<1!��E� �+"��5q!N9�C#�C�<�7&C�gZ2e�T �32�	�a~�<�bh�-��٨�7B%���f�U�<g�}[���W�S����:׀�\�<�td�y�\хA̚)�,t��V�<�&�%
��"�) l�J(��k�<Y�� ��8ȃ�Pt7DI�e\c�<���$J`��b`Ⓣ]�*p;���a�<if�N���E��� �$�q�[]�<�ÍI$"ɔ����^�<n����Y�<!䍈5E� ��a�O�5@��`�M�<bH���<��&�07/4ŋG*�J�<Ae��	���*�a������Co�A�<�̓0:�����)Fl����<yȍ�F��"�� S� ���nV�����.=�|��)&=�4b6!>���ȓv{B��G!�7Wx�h�Ī�=|fY�ȓ�~�)��J�H��PZ��n����k�:%ʤ�S�[i� Z�I��re��w�L}*a/�f~ā���	5̰��@��	��
F���-��9�֐��}�D\J!cҼ(��Ɗ37{f���,�"a�qm��d����"�jSDD��tJ4X�#枔<��la3+��e.̅�l��Q�a�*V�z�����i��@���l�(����S��͐r#������S�? ��`%��$H�$�T�L�NB�#�"OTt�`�ںb���A�ϺyBz	)p"O�<��o�,���h�%��2�"O�h)�o�20�ipE# f��`"ODUSE�ְ_&��RE�6k�B�1"O(��fA��c�ZIǏ4!6X"E"O��궤� ��}�Q�@�f���""O��c��,_��&%�e��19�"O�e�w�K�Hy���jC2+���"O��yM˪"z�E8�b��H���P"OZq��]F��W!�#�0 @�"O�C�#�̔xs ̱l�Y��"O(a���Q�0{��*6 ŘJ���S�"O�����=���E�N�8p��"O��i�����r�#�!�C �9�"O��{��;�$ �a�[�U<\�R1�'�ɺ:[l���K�#G�!)D�>9�"B�	�K�x�r� |��j1�:��C��rO�	�Q%,�f����Gh��C�	;�8�'J�l�B�5���"\lC�I�ib,��UK����@GjK6\"C�I)k�e�k	�0���r�!	?��B�� X������[�4	���2����x��(d�/6� ��nR�T�R�)1D���$��3,b��T�2�r�Z��-D��� � n�n-Ho�'bX�5�,D��f荃o�`*U�9��Y`�+D�����"��\��R*!m��1 /D���0'��t^<(�l�K�:� g�7D�(J��R�L��k� !�"(�5D�dC����5��ڢd.2��0D��y�
�nKli:7ɍ�v�@ٱPH/D�`�D%Sq�d�h��%��-���?D��Z��� M@�*7�δQƢ��)<D�`#��Ny4и�������L9D��a��$*��*��ɇND��L9D�,#R�7Y��ت `H�9�]���6D�<Y�@��2�bq{�3����c!D���q �N�z!��E��Ĺ�� D�$�(�v`j0{BJ�+c�L���J!D��&�W�C���X��ȧ�(��*O� �BQ�kd�pG�M&�P"O��2����2�������$FR�+c"O����d�#����b%	-J�OĘX#�?I��ے���U0��O��=E�ġS�c�$���>y�0$@B7~�!��C8!���G�8,�0q����B.!��O��=�E�߄Z��b��D�n!��\���Sgm�	�2�Q�#�!�D��PO(!UH	�^i��R!}�!�$�l����� �R��7. ,ء�9i�[�!\�l_dXv#�9Z�˓�hOQ>���"�I�x��D�(�NԚg<D��<}M�<J���%$r:�2��W:+�!��Y�R}0����Y�NO�o!��4��0���J�D�E.S6?Q!���SBe`Ԍ����4� 1;!��S�}M�H�pl�P��U;�%�6 !�DN�J���8�f$l�`%��I!�$	O�Bp�S8m��š���P!��@1X��+��}Q.���ZG�!���O�t�(I�� 1�a�	]�!�^�[6\�P�Q .��kԏw�<�T�zI�e�[�.��AD�LC�)� >���K\�t-�7�K�.3w"O�@��'E�е�Df(\�nE"O(I���0|\��✷4��Hi�"O�Y;7��o.U�d_��婧"O�u1Ƨ�4aȌ��'��2iN|�1"Oڈ���uu~("$�I�Z"O�t��@�wa��Kd��+|�X��"O���g0L
�+��ͨ3=��ѓ"O����H�00D�v��rN�@
`"O~�`���~1�C�F���f��f�<A�b��Ʈp��@p䐱��T^�<�'��:�8cr��|RJ��VW�<1�+���|}(�����fૅ��Z�<qb�Lz��):�e�.��-�C�_^�<�P l*(=@䥔�Rj��#�X�<��Q'\jع� �~@����Kz�<�� �F�╓���n��1���
x�<1FdoɚF'^6b��)q�p�<AP��ր� ���~v��Ga�<ɑ�L�E��M�1�� {�z}"�i�^�<���w�y�����)��[�<q�*_"}�$P& ���kt�S�<�2#ҒB�x�x��S"~P	qjDj�<����$︼x�n� |A`���iP�<��iN�PkJ�p�fE�V��x��dF�<1��.i��0` W?+�Αq���W�<�#�U�x	!V$��BVje����i�<��E	q4e	Ħ@�2���@�b�<��*�>GO����iō,ÎX�@�D�<�$�o����G܈	����e�Cx��Fx2��C���eFU	�~dQ����yR�
F�-P̫72=�e G��y�����z�ǋ�6�Ök��y�l��A)����F�	O���f�A��y�[}�-p��{c�p�Q�^��y���	��O��q��8�G`M��y��?� �&+D�st�պW�����<Ɏ���&'�̃���R���	�-E�~e!�䊿/:������pU���
�!��@|�#.Ā0x��v�!�䐦(Ep	�.�!nL8�
7V!��P�/?���%H�bI��k��ؑV�!�$޳#�%����i��@2h��U�!򄔿9j��SNh��b�'	
k��{�Z�`biQH]&kJ��:q�U�/�!�$		;Rl��/�z4s&�2 �!��O�J�>�Ð�Ȩ��8ǊS�F�!��mxP	���Y�&���I�0@!��_�y=d�
�ML�Z�����I(!�$�*��%2�O9{��h��k�"?L!��6L����O�?cd�
׊`>!�dP2L����A�HW�ʂ�#;�!���?�`̰���/�	H ��!�W��d�T�O1������!����JMI��	%nz�1�Jٶ�!�ޏ,l�LJ���o�����J�!���{��A30�'\�v��0*\��!�Lt�U�$�8���c6IB5}��}⑟���O�;J��u�ؽ%��x�&�9D���E��G��v������$D��iG�$=�Bbe�δI|x)��!D�ܑ�I֥�zy��/؍mF�b@,>D������=�|���V�K^��*D���G�F��d�3����,�*ч)D�� ��3BT�Y̠p !7�|��"OV�8�fǖ]0�l�@!l���D"O�$��G��TQsTlT
7�\q�"O\)�hXIФY��YbM��"O�TÂ>��4�����\��x�"O��pD�@Bf��O�
)=�z"O0M*2DY�nv�@�ԁD5Jl��"OF�g��,��$&��w!:�)�"O������#m�`Z�#1�v q!"O���ú(*�떃�.v���z�"O��i�@�}�쉱�c����ˀ"O.}	2-M3P%h�{�C��Hk�h�"O�=!0�P�0�d�)�m� !�P�@"O�����U�TXڝ�C�F�h��i�s"O��4L=Vg����BT@�"O���Y�� ��F�/0�0�C"O��Qb�ÿY��fǒ9���q"Ox�Z���M3���:!%|-�"O�m��˃>��92ٚU�l$�e"O�̡�䏬y�@�Û%56
�y�"O�dP @����'��!�"Ol�D.]�J���O�$����"O�p���(� ��Q�RH����"O2l�$�J4:����$��g�\�s"O�-3�"��aV��6a�u�XC�"O�ũ@o����'�ר���"O������.!�8��͕�m�<�"O���skG�7��xဪZ�{X~]�B"Oe�oV�#a�M�`�$Ch�u"O�2�A� �BI�Dϒ:]�ЅQ�"O�Ĩզ�A�qS�l�������"O�X�Ɍ�B������8��|(B"O���q�� ~����<>�`�"O��B���<$�4�+?�]�"O<�IVg� p��VM�
,���"O^X�Ө��),9���[�$��a8�"O.�K�+V,&�#�	'�(� "O���O�p$�1��!yp��A5"ODA ���~�p� iL���"O�ɈS뛐JnP!��^I�V1IR"Oly�v��&���SȂ�!jDat"Ofh�v��;�`��A��J�&���"O��ʰ
�fh�\ɐ��5%x��s�"O�c`����$�j�	h�P"O�	�3�ЇI_����\��b"O$�K�e�o���@0{��Ę�"O� R�m3Ӯɣ���i|��:b"O�D:�Y�hR4�Hcgۃ�HP�"O� ��K�>�\`�֣ɿ-|��C"O����V7B�P1ҰM����"O,1���.#�`{e�\T$Ȫ�"OE��g��H9L�y���a�$�V"O���4H^���7%@6!E.��"O!��+��bA�sD/l���"Od�b��!l�����(�! �QC�"OJ�f��45H|#g�=b����"O��`��	��U`v�8;���ɷ"On�[�3Z�KeBJ8��őW"O֡��J�>(B���q��3$��l�"O̑%�Ў!BL��cO���3�"Op)J��"�͠^Ҏ��͙�y"O�R��B�;�����[�Z�ņȓdז,*�kJ�w ���.ڂq#"O�9��5"-"�6�۳ \��q"O� ��чE%U[�d8b�E#PN2�+"O�)!��l���1�⍰$0X9Z2"O>,Cv��>�����f�ǚH�2"O-��$^���	�Č�<�^���"O�)Bp�ɡ"��܂5I��]�=2�"O�pR�J)gf��Ve��{���"O�pm�A�R�X4'Ig`��y�"O�"�D��nM�Uyc�U�]C��"OT��4�UC0�`W��#l���"O>q�bQ
W�F�xT
��+�ہ"O�T�r�X"3�MZ@�K�@��q�"O �b�oЯK�X�Ff��tf�l9�"O��؃I55p�#�!|l2eh�"OB%C/�!*�l�pI��0z��D"O��*��=��\[�MAS��"O���@hۖ9c���`��S@�+0"O��c�)�3��I����	BN$��"O0x�b�[�<������1i��E"Or�Y����f�~A	�i?.gF�;2"OB5;P��8���9�h��4�VXє"O
(�eE��*�b���f0�Cc"O��86aڷ�H�D�o�$I�"O0�{%'�MWĥ��'��x	t"Ox=��M�+ ��A�Ȟ9�|}��"O��[C٩�zqx��Ƈu/��ە*O�MC^tH�%�O�8D�v��'x �Qd�	c��y�!�X=/�ș
�'�&����Y
Tz}`AI�^���	�'Z~�*��Ϩ V�Aȧ��,V�H���'	�Ũը�<#�h4�E]h���'q�q�"��"S����ANPJ�'+�T��[�v����@�=m��8�'��$��_�xΖ�á�E0�
(�'� ѡ���un�Y��U8dU��'�BR1#õq�Xqq�Nv�P�'�D���;3�2������N���'p¡��H�4���x�oQ��;�'�bU�qa��u����愺Ffxa�'�j����޷V=\��'�����)a��x���O����'��6K�[0u@e�@|f�y�'1���.X7�r$�T��!ap �' xt�6O��nB�{�|uz�'���uMV�@5���V�'�R�K�'Vm@Ț)RZFB���T�A�'���mG��U��	�����'�.LP��:#�� ��"Gz%��'����r�
&7�EBO��h�⠋�'�Dt���@�2]XAل�RaǺŠ�'�Tb��ȩM����e��V�I[�'��i��3催��c�Fƛ�"ORܹ�+L�jɁuə8��-�"O
�H�� �zy�R�� |�`�"O�)�O�N��D�W���b}�-�Q"O�蓢e��\��7���"O��7�E�F ��	V��$iq��"O>��fԽ~ `�Viy���"O��(q+� UN.�� ,�5r��1"O�`Z�&�?(h����S�)�$i�"O<�3d�x���`��Z�^�B3"O��Y��O%C��&a�?�,���"O��P�읫�u˄�L�Q�\�4"ON�8&�C>K$��2g��)�US"O h���,'`r<S�OȌo�
���"O� \y`G�\ZD"Ƞ��=L4���"O�I�U�I�Zb4 �a�	AU�1"OĴCeˏF�NQ���ƝJ:��""O@հ�
̍Tp�;��ɢN����"O�I�͕� ������Y�B�R"O����� I���	��#c��͒�"O"%RD�9B�͢�Mȓ5����"O���E���Ё�2��n��q�"O�P�#���G�^:�K
Ŝ�a�"O�ժ�A���>��H�Vt0�*Oj`	���,S�Ř.i� ��'�^�#�jX�m�(�a��kt��'�� �5C�D����)4�����'�IA��� �~A#��C!+;`<��'�ҭ�t�2jϔ4�+W	��l��'�Z�2��S
t�ȩ��V�����'� ��V˒8���	�?�F0��'⎈��D[� ,1.jaR�P�'@V��cM�:�ޅp�ՑbƄp�''�0��9�Jd��\"b`�p��'"0��`A�Q 5s�?E�`��'8T���X�,/�{�͈�D:��c�'��sB:QA��%�߰F��R	�'���gBE(9��mcUhK7:S����'�¼;�n]�՘�mζ+X�u�'�K�	�V{��E��"�d���'��r��6�Ld8d�Ĳ��	
�'�8����S�:<Ђ�JR$�F�
�'>��F�1�i��bt�,��	�'��lq�ޤ1È��&	S�h^�	�'q.��`:}<i��f�?gP��	�'��BTFdr���N��\f:�x�'�������)��
�ҡF����'̈� 4��5|B�kłք4|�0[�'����>�,��DI+�!��'Z��р��<2��č�#�Ф#�'�"��P�2V�N�铦Z�fj�}z�' �d�P�D{-�j�'Q�`D���'Ҏ��Ʃ�-�j������$���'ʴ%��	2�1b)T�J�,��'
�Te�)+�2��q�҇/:i�	�'�![���."����.*��MP	�'��I���U�K�?oG8���DC�<!uO��,I�x8Æ�7=����33T�|P�L��G@(�wIZ*s�$Z�-9D��9v
�:���C�X�
�b�8D�� '�ةU�pZpNҶ?	vۆ�)D��{%��3\�v�S�GeD`#�5D�� ���32]((��L��A�a�n&D�\���]�q/p�eL�;tC�1�0�#D��s��>6�麰�ۼ?ږx;Rm&D��b��8NT�[���@��I�n"D�,�d� 14��֫օz�p����>D��+�N�P)����-X()�m;D�����ŗP��$�V�3�F���A:D��A�C�Ϟ�%�]�2`ӥ�;D����%�|t����g����5D�4�&�@�n�J!��ڮK0��E/D�4�F��\I�6��=�8����-D��bC�'\�x�e	�,��"5�*D���dnǛr��  mG�l���CE�)�:Y�azB�W;/͢9 ����',�s�j��y2�S*(���J���xߚQc�B��yBmY^xa�E��j��� R����y
� ��R�4O����r�
-�y�P"O�����4��m@aϓ,�6u���'�`h��?h�	gϑ(u�����.H���X&�
@��5FhR����*D-���U銁�e�2O�8,�H� �+D���`)�D���K�Bҳ]�ɶ.�<�	�FZ��D%�V�� �oS�M1j���nt���n�]�Th�c_�@�ȓ*dL 1ŉ�sk�9
��D(
V���ȓ|a�T	��G�% �T����%u��ȓG����	LttQ���-�iEr��DM��a���*��3tϚ1`�B�It��(�(�;$F��j�E	�|@C䉇Vꪨ�@�D<iv���ǰ{8C�	}��!���:fA�a�eX�wZC�ɖX ,��U�� \� ��V�X�@G}�T���'����/�<aHEk��RȦD���������:�	����!�F����,�d㑳m1@�=Qçk���r#��..Zx�ਂ�J &�E{�����^�v<��ݚ:]:T��)��?�g�)�^ ^��w�[�v�a���%8�0�'�,�p�_!}yj�pK�8"w^tR*Od��d�?�l�6�٣R��=�!�;5��}b����'DE�{�R]�vB�5R ����/D��*Ŏ�C�8z��X�8�Ab�9D��XU$�;-ht��+ʊs�hh�5D��z��քg�h]�C���QN���d.D�|�&�� ��*4ET�jL�qj5H,D��@�,��&~"E��A�Z۶QJ��.D�8��,]�U�[� �HX�,��1U��<E�dǕ`�Ap�״ŵ�
/!�y�f�6p�txȴ�F< ]�T������0>Y�gB�*�!�A��x~t���GJ�<��)��u���L��P� Q�Q���.�S�O/hq���
D��(�L����9��k�OH��f�5�R,�c�;,�	�"O��"Z�7��80��͊j%�=r��.�S�S�L�ฑG�E6?-v���@J���$)�I�M����soJ&T<'���BC�I!��!F�) D8��Ʌ�vb��E{��D%��9�z�Ѕ+Q�^�Ɉ�@��yR�7T�.Q*R#ܝ��Ȫ�O��y,��2�A`ЎPLiW+��y��)s6A*���P�6�������hOq�<��T�� �>��ri�p�(�xc"OH
KQ0��͙�ʘ07�����IH����Տ{�j����	��8�$�gax2�iI�PЇiB�*��eb���B�I�%L8!cP��_��@"Ǧ\�DT���hO�� i��0-�� ��L͍C��y��0���<q�+�2�x����- |\��LZ�<)u�]e�D��%?L!��A�n�R�!�DԀ@9���@�v�kW�θ��z"��Gu���&�Z�X�!��b�!��C!��� ��T�tsn<p�H�o��ȓ�nQ1��օq����s镈c��r��Dn���9O���Ed�c]���G\�T�h���5\O6�p�K���I�g�2��]��2O���O/AM�A L,�Z0"��B5u�$p����?��� 0�8D@�֢~��ș�KPl�<yG	m��H�A��P��d��-Is�<�t�$ov8��v�v7Z��Mf̓�hO1�Q��b^6+(^,ʳ&p�~��"O�-�EĒ+���W(M�f�rtAOh� Ԑ���֣J�B��4�.��A��"O�X�6̂9E־))�Cr������'��O�6Mä� \p������z�掗z�!�D�|��@��8%~��#�2��x|�_����İv�K�Y5-x��!(3D�ث����8R�E'`�fhS��$?���?&��Q2�O�n:�IpWV�=<�b�5D�|[�,S�C�0�W�*cHt��l3D�Hq�ON�:mfPÐ�E�*���>D� ���[�R/�b�B3=+�y���8D� Y�dĐ^	p�9�@�qt�-H�$6D��`�������+ᜁ��3D�H� 
�"vصc�
RK}L!�`�<���T>�0e�>�f"[*[�� �V���LU�<��G�!�i4J�E\0m3���9��OT5B��T>1s�N�Jk�c"�J�c��x�d;D��(6L�B�#o��*r�ذY򤽸�y�O�b>�ԧyWCf��`p@K��OZ��
�I��y�j�C
X[eΏ�AD8�y� �#�y��IN������-AD�HG#�y��HQ2�)c��q����@��yB用��|q���+j��p���yB윱d�`)�r�xh�����y����y����W<R|j2��?�y�	;�
Q��&�<u�9��@G2�y��Ӆ�>�`��.r�r$X��K�y�i��&����8{+��~Ņȓ bL��c� (��q+1�����8��!ftE'�Z8-0��*=I)�t��a�^����$T���p�N���n�ȓ@�j
 �	Q�}3 
��0�ȓ)ܠ9!�(A()F�h�	O�>;����Mo�p�tMN.b~U���RR��u�ȓ`���&��=+o���'!x��GB�j6j���*X���#A25��C�I���H��/��ɳF�^�u�q�'�1O?�I�`G�
��|�`B��f"�B�	�=�9�e��%��EA�/ǋ0ʐ6m2��+�H��	H��\��O�.��6���dB��?-U���r�-K�d-!p�@�'TV"<����?=��Ѫ^R��@cZ�����.D��HB�6,��H0�����-��+D��3bKӪ]�YЧ إ
.�=I,g�$���<Q.�q�AG2d��!�#o�~ڬ��$>?�b��Nj�8��_/*s����ɜզ����)�53�}��-E8�,HC/�oi8����B~�F�o��semL74c̕��Х�y�Ϩ;0�${�!X'It��@)I,�ybO9O���"���U�'"ش�yG	~�*C��kx�k#�V���d�O�6M� �yR�~��y��ĭPɶ��`��[BE1u�\�=�B㉨a���Jŭ&�&8��
� y$�*O���uw��B�?�n�ڭZե@4dm`�$,�y�!�$�Ab���#�09UX�2��;A+2�'D���$ �������>����3 M�z-D|�Kr�4[hv��`Y&e�u�@��y2�.G��a*�j����ݙn7��m�~�'6Q?7-
�[((T��P>�|IĖ��!�DF� � Ps�J�^�8��$P���8��HO~�8�f���DZJ�&V���'�z�8왵�L�HP�qJ��q5>�ȓ�����Ս"�(���\�C�& Gy򞟄D�D	2f2���t�_��j��c���yR��y��dj7	��{k�� V��ē�hO��� H�a��C-Qಓ�Q#����"O����ΝX��Y�U��F�
T�v"O�P�%=:q��iu!3!��s�"O��@4�ӽ��]�$טyE��$"O4����<%H��2�M�".��A�"OF}�g��0��=icU�|,xD�T"OX�g�A@1�d°B)�=Q�"O|ȡ��)<�4��$�7���"OV��6hC�\K\�!�bF�)j����"O��V)��-(�u���\R�ڒ"O*йGA�04�� H�iM��*�"O!!��ϼ�5�D�
(VZ�ad"O�ԡ"�Kt.����N�n���"O.,�'kA���]i��/�(��"O�%r�aP�L���oN��̈@��(D���DCw����$`۟|�����(D��)�Ì!'�L��ߵL�ʽ�c�$D��b��D�)J񸄬O�Дi7�?D��B$�&7�$���+�� ���<D�0iU��Y\� ��
��<u�<D�D36�������ãw���";D��;&�i�&�Q卄K���@f'D��bcdHd����Q��J놀�!$D�; ��i$��Z�׷����@,5D�$� �A_��IKʔ�h��U$>D��� ��C���I�F[0�3�:D�l��cE	A����`Lf�,�8�	;D���6O	�Ĕ�BI�|�8R�:D����*μ+h��������ȫ��%D�<!1R9"���ѣ��E{�k$D���ݨG�<K��Ξq���r��,D�pc3��32���c��� �Q�P�%D�(�Ѫ��+X�$󐨍M�v�	0D�,iFIK���J_�1e0D�l�$��,�0� ��.a�H���/D�0y�Ö���e�lT�l�p�m�PA L��YRH���%	%X��+"�q�.LP�DH��<8@C�E�ĆȓL��4��Śj" �vĄ1ݔm��?B���-F3>'\)��"�<"/���ȓ9*�B�� �"M�TO�z��Ն�8vT(iQA�4����e��w � �ȓ"<,��G%�$)!�$ �F1���d �t���11�a�d��ȓgȠԳ��.GO� ��\�}��q��W�t�V��_Lqb��'jz��ȓ;�tyfjB�U|��3ץV��A��|��=��+l�Q��c��OY����HeQ۵��	x^l!�d�nj1�ȓU(P�B�9n@��h��O�|��!��P����*��W�`�R@�>oА,��\X�����
u�Djv)
�z��H�ȓJ~=��*ŭ$#j����ȱ)���W&�Y4�Ɖe�� `�`�%- R��ȓ2�����Y"pH�y���\8ښ�ȓTT�H��
	q����>_q<�ȓ<���0ʃ%HX@�k«:d؄ńȓu_����4��DKDν%����G������l��Ц�4NX�ȓ�f9y�*;9ɂ�2��4l����ȓ>�D���Ծ["�z�(M+|��L����}˳ �
�&���ޤ.X���w��<PE⌽:_v٩��qN*%��e��钋Υа=ٵ�f1�����V��`4"P��zp�F"��J��X "r @r�݄����̉?r�B�)� |���#�?{�YÀ��8�HDb��	Jj�zg�Ǒ}�."|bVn�.IN�H��I4�dUd�u�<QԄ�n��C�9Zׄ�a���7GK�X�� <�P��'��>�		����I
'x��-�l`C䉯"�D�գר7E�,B��,.�f�X7b��DN�7h��R;H��qs6�J�Q���+̦'��{N
��\"K��J�8ѩ��_�T'�Q+��.��T"O���3mB��1#�4u����'-�q��C�e߀"|�GP�v X͑ǯ�h�
�{���j�<)f��*1�|�Vd�&>E#읧`pH�BSk@mC~t�'��>�	�OF6�z�aθq�P���6i�|C�I�CH���I#8�тW��3A����9
�(��i��zB���~�Fl#"
��Kz.ݛɒ�SEa|b�ލJ����H�Dw����B���33��LN�	�'d�8����Rs�D�e��[��D�df�(3�,�'&�RH�̂/lA��(S�R(��m�.=��D���a�V�ʏDhчȓJH(���F�E8�]x�n�+�6D��o>|��( d��E�%#^�-6�ȓ=�yaU��)v>�!p�[����ȓ!��At�
�!����E/��9��v"�Q5b�)/	�QTj�o��|��	��@$.�l�92(��hl�Q��i~�0�"��s�С���+�|$�ȓ=����(־'$v-T)Im~��ȓ5��52`l�x����ԍ�L��ȓK�bTX1�Ƴ9��݀���l�h��u�j���LG0_�]L��L���7��Q3$�%}�����H&Vq���ȓ:b4�QQ	�����ڠ	�6�hM�ȓ>"h�y"/�����>̈d�c�F]���h��$@�3�f�sd���W�P�s�ɦ6!�$֠�
e#���^�`�#��a��V�� oC����	?4��9����_��1R�eĈ����9C��� )Of�	�"	&r� 0�ǟ0�"�"O� �v��7X�d�B�ȗ�ewDCE����F�����Ϗ^Zn,���V�~d���¡\f!�$	A�p���Y
�@���=_�<@d -�I��H���D~6�A7� S���hD��4}�C�ɂJ'H��	�	���sA	Zd��7�D�?�.q�pJ��c�&r�Z�yW/U詇�v�T��'x���g�,H�(��ã9����	�'�.��s��f�:�Jt �F��q��'���E�T��Do^�>��ѩ�'�΅���>�zIR��7T �A��%M,���'�0��"�XO�S�'oQ���ȏ�  �����4��8��	$Dz��@��D�	2�9���ڕ�G	5=�(�I>�g�T�?��>�O5(ƈ=�`�CRm��z����q_�@�Eω4Z]��v�>�}*� �C����p�
�Z`��R8��t(:e���ā�p=.��d��Y�<	xU΄5`�O�i"pꑞc�S%u����' ��1p�`Z4j�,2�
I��dϖ.ꨇ�	:3w�P�SL�0�ژ�+!����3�F�:��"��ih9��D��{ѤO>��U�ؘP��qS�"ǎ�&���)7�cfL�6͜	>�x���,E	B� �@E�N��3�*w�CQV����]�x�J��u��<,���G�Ģj�����M_$˓���SKʖ0c��JË�~�ץػ��ˆٛ]9�)�1G�?2Ɛ 	A:oݔ��C�?�;5hԌD�q��[�Q78��O���`4�b��a���q�	!:\��'�iZ��Fl�ЊGl���y��':�}j���/ظ�ƣF;Ɣ�h�l�'��M���h>lp���X��FD��	�ş�������O������0��"�I��J�0���'F��V(Lk�'o���򦖴u�x�G[��`�ی+edE[ Kr���@����ݨ���ƎIznT�ǎ�;@h�[a���i�w�2�8��"��]�t�8�8��B�'���a��F�p��da��K�����A8Yg��YD�W(O�~�.�s�K�,q� k�Gf�<�<y���g�>S���Q���"G� �}&�π ��r]x�� 1�Z#i��d��"O~��֊J�6�h ��dػ��	n�����&�8t!��F�ZQ?���Bo��8��T��)I��[@�!�q` �Ʌ�ȴFa4,"��Q�"� 'P]܆TS�fB Li(%۟ўܩ�)P�Q�%
l,��rn6�O:h�0aD�w��x��ŢZxS���K6���`�( 	D�QaŶt����DN;�����8�>��a��$��t�D������$�t9�e�ѣ@G��bӵ3����f�Ƌa2쑡�!T��y�dD�H��P���f�,I��؍uK@���d�p=Bq ��A� |��@��s������-���zc֖H��!�B:D��yqE"�QY���O�@���K�Sr �Q�۔a�H1�������Sb�'v����'U7(�������'���*O���sj�'븧�ĉڂ%���H�g�(��pMZ��|HJ��Ï/(гFB]2Ю�� �'�l�V雬�(��# +ۂ%�M<���S�cd��)�<M��B�v�P�C�O��(#"[�����+@819��NND��B�)����'E�)1/
ͳ�O,g'�)��zZ��JC�Q�/���ZF��?+���?5��U%P�SE�1v��Q���C *{�UE}r�U<Q>�4#�ɟȨ`��YXP���!w(P���i1F�[�S��0	�u��r��?Qx���P	/��8U�M�G����*9��D�(qgr H�����~�HF�!�N�Ԩ�����aH�ֲiK�A̦�>��c�N;��Q�'�V�y�NW������:��T�J��I�o r*$Q�f�	?(z��*ܺCp�݋IS�iͧV�(xA&�:���'�W��Ԅ�ɲ92N9� %�]�^eY6NK�d�&0�ࡑ_���5lT�`��a��B��UP�_�����,0:pEp�) �2N ux��*��>��W2���D2�ӛ5��-����|�p�	���$%��a�hY�b���7�ǟr�)Qb�韜=G{bמ���D���Ls���~��U'q��� &X�T?�� ��B |��Z��0wKR�0E�U&Qi�i��k �r�"=��	6/F��իɧd��R�=A�rO� ��F�x����6aE�V�x1�S���ߟ��)�@G�7-@�:B����X�W�'t��9���o�`13�'��n��!B�D�����L�3RqOf�}�I���K@���h"Ltɢ�4�<C�ɆL�z��Fl�/,���C�<EC��3j�^�ȓ̖O��%�B���O�-�����4���I�]��i
F�V�"b�6 !�$�s���Z��`��\s��2�F#q���*Opűh�i�g�I�j���xT̘63/ޘ��˲dvPC�	5R�d�aǛ�]td,�����`��O4������94��Q
�I�����长Z�u��>�*A�㉧U�z��`U7�,Ċ$1O,������4�̇n��YAR"O�@��m0�z�h$Ď>�*�Sv�>���Ȋqn}�glӝkT�#~bw	]:F6jt:5"��P�Ԩ\H�<�'-?(e,��a�<k��������}�l��"f�y��I�By�}&�l����@�PCê7s��q� ���+Җ�<h�6����b,��(6]I1��%l/x�ذh؞@y��ZvA�Yz��ߋ2-��kd�%O�a��z'ޜ`�TZ6��T�}W�U:!�0Y�qK��5�Od�r�?O�1�rȂ�Ll�	��|�p5P�>93����x�R� �8`V M ���,�Tp|��HJ44s+�v�@<r%�GW<���؋h+��;�A�8������1=���vB\?��
k���X�i(��c@�FGy<����ǐ'bX��&/U�X�u q�'Xf��A���ã�8�rWdуW��d P9>�!+ҨsN(�ϐK}��Ȉ[�L�K�*���i!6ɻ�PGu��I�ƥ�j�0��dޭcHx�W�>YPjƧ	�~� S"s�չa�9�� v�:�>�K��>	D�����W�ߘu�ax�$��I��p��.�@�����L`�tˏ�+2������}Hb �%Yx�|:�@DA$L����
�4B����w#
Y0 (��x�hnĄ��ԝ2�vx"�L� ��0��&L+k�Z�c.g�Z��́laֈ���U_yZ���Vk���W%
9
v���뙽��=��G�Y���� �kӖHc�E35)e��G�x���Rӽi�t96&� ��\��O��͊D��%>7-S3hP#sL��uY�a"r����O��7b��.hİ��Z�T��V#�,��'��!D���n���g��!��<��bE/��l�Q]'S_���A'CM.Bd����铻�`��@�SW A�@M�#��=��Jb$L�"O�u�1�/L#��Ha��/X�X1��'Q8���b
�`���ɻn=Ҡ1&�P4(y|ܑ��2�����G�wp=��Z;�M� ��Pu�K,�BZA���V"Or���T(��aQ@��y� ,���I��M��k���h��q��80]4(#�U�h-�E�s"O�0�gޅk�Z�8��]x`��"z�U�����Ol��gH�
EV���M�3k�`�"OaZ��Ϳ-� ����-AQP)s"OV�+�NS�1��$j6��,@0����"O^�u&$4����ĥ­(Z�iU"O��Q�)�5��:��ýDp=��"O�仧��>r�\���e�=��"O�x�l��iT�9bN^?Y�� *"O�y�Q���M�	����'M2@E�1r<�h	$����'ܬ��-�0#%��*Х.I���	�'_�d1ǭ_� "p�g�ς�&H
�'#�`�N�&R:�Ȇ�.:���	�'�����JX�D��I/��%�L���'� 8���6Zyڠ��$3n���'Q�%�ޑ$��0���`�' b���,öo��HЪ�~)���'��:�酞	���!�AAp#,�1�'�p=�D�0_>1� S��n�x�',X�9��M�d%B)���η���(�'�V�;q���n���!շTX�;�'�����^�/7�*3e{x� 9�'e Ъ"�
M��m(� ��k&}*
�'Vj��を,	p�|�a PfG���	�'��Xxp�,}D�ԠӄE�^Df0�'����K�d�C�U2Uòл�'&z��P��XJ�R)H�h% �'��
5��T����#� L�rT��'
VĚ��@�v ��CոB��ܨ�'�Ρ�d�S1E,U��EP�8.*|��'��0�u�ՇJ��-���><\�
�'k�u����h(� "%z=dB
�'�*$R��	�-��M`M6M��] �'�lU���ՋG��8àE0�Ҩs�'�1�	�3Q�����운2��(+
�'C&@��܂o��䨆���!hf%S
�'������b�f�c�G�$��	�'�q�C�-5�pb�B݁�h��'Cܫ�*�+4���'9 �<�a
�',����lRLi�Q��'x���A�'�0�1��k$���%�x��ܱ�'�EP% �.&�ġ!�1�b�k�'�Va��%KK��uK�
ʅy�"��',0pIL�0�D� ���%p�
�'˨} ��$X����ت>M�̓�'.�9�&P2i���a�HA�>f��'t�����$<�x�tmX�*o�9�
�'ሜ���O�E�8���Y$plt
�'�|����	 Э
������i
�'��C���b|����{O�H�	�'Z�S�ə�����~���q�'�n�H�/�S���Ibd�6dcLJ�'�zؚv�°
�H��Q��Y�T)Q�'�2Ub�*�0h�`���!��a��'��\�e%��B����%3�	�yR�C�U�l�4b���誑�Z,�y�M2G�X�Bl�!	t������y"Ņ=�V=+���5#�`9@���y��MH)\����R~�y���yBLT�DLѷę9 �`q���ˠ�y�P��bͫE���M��}Ƞ��y
� �(�Ӯ� X��ǆ�_�>��"O\@2q�V ]��i�(@3x�١�O  ��M�#F����)'���k��"ȉE�>}a|N�*��}�ÃTϦ!C��>]�ȥ���V/@V���"O�{ �K�*�,����.�"�1a��ߤ3 �!���0W#|JR�ݮd�Q��҈嬭㖎@z�<�PcP�`��[f��c��3M���a 4�'`�>�	 e��z�iF�I�(����Y1I��B�I��8���\�(ሐo����S!���HE�S���Dx���Cg�$Zjv<ꃮ���{���;�AP�ؙz�����$�1�п��dQQ"O&yq �	�-��T��ŕ7f(���DžA��}�"�ёc^z#|�T�H�|�r�@�(ƶ����v�<��
���ҭ��h̹S��ʭh:t� (� �'��>��Zw,��:��d�:a��C�	�8��m�s�Q='���b�fݦG��Z�8��K�KK�i���d�PꮸR1��U�ʁm��Q�a|hT�n��u#D(u~��5�J=m�(����L�I�Y0�';�,z��۝L���!rf߿O�>]3���S529�$j��;ҧTh���κ:����y�؇���)Ado�R����BI�
���a�f-�͒2��"&C��Z��ȓ�1IGC��>i���'�B*8Bб��?��54
� W�~���T+*[B��ȓV�X��7ą�
�b��oO _�2��c�RA�C��N2��u�Y�E�L��ȓbf�3`a*S�T3o���"O�T(֔E5�@�@�-�jS"OL���NP�?�����J�#�P���"OD���C�� �� �u�3{�� Z"O��X��ރ`��l�O�4-���S�"O^\&�Իe��$Z�!��$���W"O�X�-tRY:ԀP�M���[ "O��d��dF�1(��ߧY>:y��"O��b�N��`¬�'D2\#�"O�=�4��c������ֻQ0j�A'"O��Ŋ��8���� O >+�8��"O��YP鐂C�^3 �R4�q""O*���M�o��Mn��7"O���+DQ9 ��Mч_�� �"OD0�rN��?�5����L���!�"O`�+�
��(Pl7�֕L��q�"O��1�#�N���.�2�ڠ[�"O���g��?c�hF.N�0�YZS"O���G�U6=Z�Vm�ȓ�"O��ɖ�[9�0�2��9�4��"OH�2��+8��bkL2D.-i0"O�<K҈Q�4il�TiD	�9��
O�-yT������⊼G�vx���YW�ɩO�5J�������O3"���ﶪ5�`%9D ����&v٠-Ʉ���`�5�.3Ф��'H%��*�|�gH� ���}&�L�բ�>&ܑ��Fϑ'e�aRͬ<yg�֚>@���i)}��$��y:1(P/�a�*`�\B��!@ӂ�&D���$(��H���'N	$�҆�*v��]�J�8h���P�~��'H�2�di��]��'�ɳe�ߘ`2|YS���3��"�s����e	�g�:@�F��v@�%���"R��A6�c�L��a�	�"�L��J�"|R c�W��X6f��eHte�q�d�'�T9;4�؛ٜ)%>��ΪoJ��0��f��ճd�T��o�˗I�k�g�!��ȱ^<X�z�S�n��hN�M�'�j�Q�T�TŨ1�Oq���S���.J�@��V����c�U�D���¤KA5�p?��5��9��BK�:��Y��؟(2�?qx-{@N����&�3b�DX�c'Wr��.��|�sa�"aR�k��ͪ��X/���AL� |� bR��x����� � nZ�BK~�bѯ���S�O"�q�d�� �ȉ�@�!�.��Ó+�5 �̄��S�? R1c��O2�0L��ɣ>�	R��2��ɓElpC6�3�I)Y������
}ֶqy E!�f�'��e��J@J�S�)X��P�-��]z2��`�{�D��w�Ȉf�.Lȵ�'J\9�&o�p����ǤV[(X��e��������g"� #T�Ϋ|�\Y�b�.R0�����n�:%�3���ۆ����X�$��s�M�	d2qO���lX+�S�D!� ��p��jB"O�ԩ"H�e��M�Y���Y�"O��j��_溈B5�<�4QP�"Ov�餪�4����'���$��"O=I�Î)	�����=tr�S"O��C` ��~���w"�?ξ�E"O2�a���r]*���BJ%`��|Ё"O�XX��1��R�B��q�U"O|a(�HN1|�!!M��j8ٵ"O2��RO��n/��"�Rw��y83W���"�KqO�v��q(#7O�!UH�{�j`YF"�<��qæ"OBU�*��Q�`�Ѕ+ǲ/��]yПx�KWgZ:U�� )hXT$�P��П�� �LR#9+�� _*!|��i4�'c��c�3kB�X1�i�mB���+J�^Ě@�&��0��e�6�>������~�e-=�l��B��E_��*�kԼ�OB�Ⳉ�E"hiJ��d�M�'l5`�lþ5؁�3HL��?i� VC�"�K�=lO��B�c��\���`P)��m�Z�c�O�B���L�2x�O��K�2D�ꝙSzb7m�!-�^��b�</&x�wt!�ͥ��p��um��{�B=��O��L1�܇z���Ta���I9��ϧ%S�y "�2bA�� ͍��م�ɰoq�|'�ħ�x�!*� 6c�1%�]�uV|� 	.�� �O>��D�3����!���xJ.�0�i�c]D�af�:�sO���0��b>��#(��Vs�R�#Q��a"��OY�(1���y��`��O!������*X����e2ь�j��ҧ�I�j����4a<�M3Wo��vf\�j�NO2U���"�|�<��A��
�+@�
�c�2�x��7)� Be��s&<,�|R%�a�K<]���R��:P	�h1�]��܁%�< YfBR�� MH3������%�!%wN��=����'̱Y�z�8XfFI	5V�C�' �U�)~�&��%

p��D��'��
�;�8��a�yu2�N>�&!��xw6�V�1�}�N�cdʖ�x�Ip���J��ȓY�z���
�j���TC�
 4̸�W(b�ʓI| �`��xR��h��x����%D�pxӎŷ�Pxr��(�d���M�w$�|�I�/U,�R��(8�Hb�w���C��� hҡ��#�>nw`�Cf6O�yBǌu���eϙ4�y��<��C@�/v�P<�`�J�y�.�!���7ëjB��@�i�4��IҐ��A"ҁo�ȹ��P���;#LB�G(�0&G��k\�B�I4DvP�W$�!*�&A���t@�m#4ᆧ~@Γy���!��<�3�d}w�r�K߿\T��e��z���D�?8�V�S�
�R�a �I�g����T;3���I� �`����&` s�L�]�(3��Z2
J�x�L�2uRb�c �͔o�80�b�i� �O�1���v"�{(@�	�'K>�0�E/`I�eQ���aI���,#'$5S��$,�D��U
7�� �@k��Wrv�:��Z��y2�U�R�|��dC!?u�$S��A�~�VmI� L
H2�	2D� ���S�l��d#}�?�rԳ������%Pr̍*8xV����'���Ie���,XCFva�'�*7��� J�7fR|HcF�$dXM�£;����Ub�m��$�H���$3����(����1k S<n�@�ϗ����)���������u�)�
sA>q��K��K2�\��雟����%Xi�@���N�ay�A0,�����5Fyx��\N�8���\�� I���P�Gc��>B���Ip!Ս5��=���֦27x%�K�.FB�C8o�!��T^n�S�Ԫb�(p��L�P��i`�ņ6�^�jV��<��݄SWp�S/�h~Z����ˌ^�:\k$���QZ֝����=	��]V7��iU�k�4 n+'�������7;@�¹iΑ8uĐ>zYZM��O�Ԋ	#x���&>7�� �l�A��m�����D!<��O�$�Д! N�Ɋ��;Q�6�{���X��-)�a)@�\n!j�DH���<� ��b�Z�%H����!N'y�<���?/����$�|�d<�'!�d�[��
�v��w��*��L[#�T]ӴE���My��]�0����!�M�2��I�E�m[s���>a{�f�#KЎ��2l��[�FAST`X���=�uʔ�F�� �F~�L���0!�(�3pL�� 0)ɥ"Ot)��)i'8��ae�4I�h�E����zDfDg�Os�2��^N)K��m|9��'F|5��oA�>�a◈K�~ �g�׳[����{���'g��C���R��S�P��as�'A�qz���?˂%�џ���'n�\J�gZ�"0�x�a�(
�.�P�'�`�zCk�,=��{�=���'q�D�\�Z"��Ap�������'��� �D�����@�����'��"F�͞�c���6!,uY�'A�,���T�W��\rr��	"X���'��!Ɨ��x�aFב&�p�:�'�d=�`.�*= �Z�j�er�'�EXŦ����{ K��I$��*
�'r�ԍ��I4�a�N]�=����"O��p��51��m;
��H�ԝ�"O�E8�L#z|�
' ��(�q�"O�p{��֜Z7�MqщQ�h]�@�"OȰ��Q�@��z�G�*!HR,p�"O��q��S�%-������PƄ��E"O� he�+6]А�0G��$�� �"O�=��HR�f�`�&P�#��p!"Od�$d֜%���3���;M�~��r"O���$�]�$�i��� .B���"O��*�n�-S�-�'�X�\�n$9�"O��xq��U�p��c�<��)�"O�ٸB�WZ$�V`�|h��""O��d�P*k�DMc�U 1�:@H�"O��!lF�^)�,@Nq��@�"OB�K&��9B깉��ܟm��hi�"O$H�",}�$�C!c�f��*�"Of��l��p�ՠ!� p��9�d�<�c��`�rʞ�&�����Z�<�%,���K��>��x8�i�[�<�#Cw��D���Y�i�D�R��T�<�e@r����c��-C��QWoP�<�V�K&��%�Ţ_���qC��O�<qe)I���]��G*��لD�B�<��-�s�4���j�������<AG���Gp�0��+I;_U�|���n�' �L"G [�VN1{�ei5����'欱r��ͅA�%	��.Qr�
�'Uڍ8���0q	@��n�X���Y�'���`sˊ��
]�0$ݍV�Nx�
�'t��jU�g��b1�Ի]��z�'8� j�n[`<��`�B��,�
�'��Tj$�J.t*ԣ��SG$�i�
�'��1`%�^2!ll�`�L+���2
�'���s����zp��˝�v �
�'V�A�"e�6)+�J[�l�
���'S\��5�ֆ}zL��)�!m��H�'%6	�DUT\�P�Z�Rz���'��Fy��.pP��<�d���+�`p�P�$]�T�ÁM��M��,F$�M�O�?ip�a5��1���{��DB3�ކ7�������$�0�0|����U90)�f�Y�""t)����<Q�#�>9 ��d�ʧ���Q�AH�5\x���d+<Y��ũY���_�%�Z�S>}��X%Ԫ�k�(s�2� U���,�F���~�=J��ʧ��O�TQ��<��BSwH���� �%��I�MX�%)�S�O용�E�=�J
��+<t�M�׎�>yG�0vn\��O>9�牡l����@7z��<�E�~��N�`�p�wo����3� (�"Fõ�%:�a�+Qp8<��ҬBa6X��"#Լ��Oq:ʧ(�`i�'�ԇy�!p�ǃ������/�6{Hy�W�Q�'z��ղ��O��:LF�0Ԏb;R�Ç^�&φM��D�C�:�)�#ſ|��1a�l�T�s��s��(bAZ����Z9U��H�X;"���?O��[�O���	�ra���e�S�JA#�A�	kL!��#(�N�Zү�4����@�1(!�$�94���hPʑ� ��Q��o�%!�䋥zW��2���u����[��Py"KC�nE�C�b0=�`�)�yk�1N�BTۄDX�H��AP*Q��yr臱n�4D��?�Z� !O�y�&��j-�(xtӷ?:��B�Õ?�y����K�\�����!F�Z����X8�ybn\91��̡W`B�;﮴y���y�Z�)�=`OP�0�%�#��5�yB�;	���c�.���s�O�1�y��O5-uL�I�b�j��3O_��y�`�+���[�C�,G�t���.� �yB*N�9l����6FR�x;E(�yrE�r(���%C�R�)�t���y�M�;jጹ�c.Bh�����y�$�/�:`j�� ,{i|�Y#ɫ�yᚂ��{5�AR(��KD�y���T�8��Ʌ�@r�����y�ܓo�dlÃ�M�E��q*�h���y�`ϸ4�PK1�X)P�1Y�j�&�y҄��
\f�b�
^=R)�lqu�H0�y����Eh���	C�teA��6�yb�2b���Yb��A��Z�O��yR�B%����T�+<0J��ќ�y2"_'�`�h�T)&{�����Z>�y��T��Y����5�`آq,U��y�枏O(��"R��'��5��i��y"�@�wvi�3�@�{=��1� �y���<���q�������n��y"�C�c��2��W�rڎ)4"�'�yr�̵hB�tc2��n��= $���y��� �l)c@��^�֍˓�̓�y���,�҉I�&��Uz���&��y2!Q�r��}�Kճ��%!���yBI��h�0�LZ�
��Ĳ�yB�l\��w�U� AУ���yr�N1H:�}8�ˌ�L<]2�G��y�kƦ����׊���=��f$D���)O0N����&�'>�eK�-6D����K�2� ��1�����3D��:sJ�-s`E��\� y�L�,D�8�C�6*��;a�Y� ��X*r�-D�L��t��M���ˀ Ѡ�9D�v�]5�\��b[�CF��&6D��`DO�o�"�1V��v�&t(4D�X;�(]Z���K�=1^xn0D����F�y�q0͘�1�1�-D�\;���:`��욼i����� +D�@k%o�e0���j�J���(D��K�Η5<�~`X�ⓧ=���z��:D�H;�M� {F�
p����j`e=D�<���(%^eA�AΖ���*�<D��æD�+/_���9�l�#l:D���"@D=X�C0	B�D��S�,D�djSW�1NBWAϟ<�����)D�h��'��G�"l�g!=O+(��F)D��CA�L��p(��7��1yB�9D�D0W�ɠg�D�r�ݷ~
��ِ�6D�� (��t��!V~f�ђ���8)��"O`XC`��(�x�y3���8n��S"O�����'�	r�I�1�"O�\J��I�_ۂ��am��.� ��"O찐T��?-zT���	N��5QG"O6Xro &��8��������"Oܹ�T)3�X�j#�9����"OF�A�뜭�8�$i�;�"O@IK���(IR��Q�v�V"OlոL	�T4���< �T���"O��P��O�,	��	�*0Dt.��U"O���S�l[��0��Ccδk�"O�Z `ÐB�({���+\��A"O�H���P�I��Ϟ�"B�ȡf"OBq�U g����A��Ch,�u"O]�Ѩ�XI�����-k.���W"Ork4�� 9J��wk��H)0�R�"Ov���L@$0.�%ᱤD*��S�"O0Y��%�t�g�g&P�`�"O�]��e��X�Rڶ_�q�3"O��z�o�� �󖁈 C���@s"O�\�r�΢����z���g"O���R��h��kԉws^��"OB�S�K.	���/�`Ib=��"Or�b&@��g�R]�O��=��"O&0�W�A�q�����g�8  "�:�"O�dfL���i���M)Q��K�"O4	 ��c��*�Ԯ���3�"O�hP�@
g�F�sb"V)^@�JC"O�a��)��<(J� 5!�Tx�"O�u�H�
ZbX��	�d*�:!"OtQ��� ڪ|"�M�Ch2L��"O�����iq*  ��Z%/K4%J"O���D[�l$:x�Fƞ�8b����"OHe�g�\����P��zI�"OZ$AQ"ЎN��Ax�#D:�(��"Ob|��'X�%�V0  G�p�'"O ( �FF�)Ƣ��` ]!��Ab�"O���RbM�!�Ia���Yq��� "Ov�V	�/9*�a���POdh��"O��coםZ�$����O��6"O��8���]�3w��/W,!s�"OL@2Z�=d|�В�?m�)��"Ot�T��&}�.����%�5{v"O$���- ���KA"K���"OL��$J�3��Y�d��.ג	"Oxai�[0��GCL�@�DI��"O�q35I����bs�O&A�D,�v"Or����C#*>�Q ��Ӂ( ��"O ���d�!B��-�����HQk�"O��ET�j��Ӏ�>0$%Z�"O���U-Z2�i["����ٲ"O��� �|S��DM43�J�
u"O�}��.\2"c�7D�lY20"O�颵'�3-���Uh�9E���i"O�$$^�R4>q��'�3�`s�"O� �m�
y��T�7���x��h�r"O�]�C��
&�p��X�h����"O�A�C61��2Ρ~{R5�0"O�D	����h���� 7c"��D"O�qJĮ֮Dp��Zt�J�mP���!"O�i0��3(����+�'�x8h�"O*�0�ǡ<`�H!� �xB ��"O\E�V�8��a�!��Cj�M��"O� (%�e��C��	�C�;8��S"O����F��~y3!��U��M�D"OB�(c�ά.�bP��O_�X�i""O��s"	�8r�#��L�iXa"OH�I��(%Mf4bU�/bZH��"OЭb4�
�Z��\є�M�n��S"O*�q���
#��{�B##܈!b"O�4 (T%FŢ!�1M�$�����"O�h�C�ىZ�h�p,�*xŐ ��"Ov�� �$�'�I
F�4@C�"O��r��?Iih��c�2.:�	2"OdY3쑔%N�(!�I�X%�ͪ�"O�M;UKLj-�Q�;:��`1�"O�̓@��&�.��$Z35��x��"O��2���@}H iN��x�T"Ohi���Bo<}��hS.VmQ"OB����Grt���pY�"O���#oQɴ�I�b4��]ru"OԀ8�fݮ���ʣ$�
Ύ��"O(|Hi^�{�8KUH����a"O8x�F-`h�c�̦x�P���y�Ā,�x����ɬ	d��؄����y��̟`�ei��
< Z�̵�yb(�9!z`Q��"��s/��y�J/s��I�P$R<�̹;�%�y���@Xx`�:e
$E�U�ƛ�yI�&<�1 �lN�Yu��@��?�y�e�7	���q�C8%��Uhs@0�y�.�lA����45�x2sk��yBD�4�n�X�/֣��#�����y�h��qC.��+�-
ӄ��y��"\��1;f��5�%CG���y���+| =aǀ��QY %��HԎ�y��9^��8!
N�=f��+����y⩀���̱��2�PbdmL2�yR)�
)������6;�&ɸ�+���y��@ ����W����"`��ybɚ�)0Te����5|FL�@�	���yb�	'�zi���v�^�:����yb�P51�̈�- m��p�͈;�y�ș4� ��'N:�U1J���y����i ��U��,0,�ɔ֩�ybɛ�F�@Ż�aE�*�����
�y��)��Lp��W>(,:�����yr'7��z�.ݻ��Ab����y�lW�R��=��'>i=fyr�$+�y2*�^@T�bA�w��!-_�@��mG�di�X6vE;�CQ�+�虇ȓGa����և]�j\��Ɉ/=7j���y��#� �����gY]�v��ȓ�x����ܬy�B�1���j3�i��M��i�gͪ.Qd8Jc �3�d���h�=ۥ��U�DZ�\� �d�{�<�!`C�8��$(�MZW2N`�w�%D��"� \j��T*�g� �"v�%D��	LW7G2�Q��Lj`��j#D��b�N�A8���C
F�Y��d��"D�D)�m�tD�a�E���<+�+"D��:c�Js�@��ʎ��h���h#D�XZŪ@|�d,k�hH�LbF4BEK$T����'��td��	�T���u"O�2�!dI�4@a�Z 7�Π�p"O���T��� i׀G�1� �H�"O�<8�-�=�hĲv� ibN���"O� 9�� Y�y�R�]�d��ɘf"O֍a�'L�zDD�t��I�8 k�"O��GG�7S ����e��F���"O���#�N2VHifD
M� �"O�L���ыmc�Y{���ZF� k�"O���℉�cϒУ�ʚ]�<Y;�"O�����BS�ca+Y�?-Z hq"O�`i�
�"(��1#e�Q/"�5(F"O���^27x������)z �"O\   ��   �  /  �  �  �)  !5  k@  �K  �T  [  �e  ul  �r  y  G  ��  ۋ  G�  ��  ��  N�  ��  �  ;�  ��  ��  	�  ]�  
�  ��  ��  &�  ��  ��  � 9 � � 6 �"  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�9�x8�� |e�o2+̒Ѡ���vaz���O��8�[&&$)�ޭiJ�:ǎ~���	Cx����ԊE ԁ�)�p8�k�>�����$ʌ{B��/���2e-P�n��%g��y�B�v��`���<��tρ�yR���,�wI6d���1o��y�FD? Xp��T�ԥ�1n��(O���D� "� Q����
7�<@��A�<zQ!�	5t����W���<&�-b�@�;�B�ɞ�H̻�kB�9d���_�Jؼ��$�O�c�4�C�
(�<��쓧aɈ���8D���K�&6t^��Un>{Mn�yRd1�d<�S���\��@��e}P�2.�=�v���6����I2cS,��&��:z����y� �+X�$"s���m��	iܓ)���F��#^�.J�e�u�nԄ�k���E4s�D�6fٓ����'2ўD+�"�٨Z��\q"��*o68H��y2��'"��
�(|B�FJ���'��{�Չ8༫��V������
��?�ԊaӌyZ���k-�\�dG�MJ5��"O2T"��Σ.�B�C5�6x4`��D�'Pў��"��12�Hҷ#�ui|x�t�$D�0���� �BMK�EVNfHqȡ��F{��iC��FhZe,Vu�]BD-I,!�Ą�4y�FR�\?����S�?�qO0�=%?��@�e6p�i��7e����4�|��!8�0sf�O�,}K$~*C�49i\��ה1��Ɋ�n
�<^�x"�I�]'$��iغ]��=H��ʟ {B�	3YPI�"��F�di�&	�Z�C�	FYrUh�ڵ|(0q
H-�C�IpE���ӭ�0p�N��`���HB�66d�{q#Bh�|c�J��d9B�	jNm�#bN
�����"9�C�	�r#��0�����5� �>@�C�I�b֬�bM�:ƌx�rm_ >b�C�	:P�4b�^�3�|��ӨɊ(��B�	�*}(�JJ��N���(b��B�	uA�b����X؀⅘ � B�I�l"��P�V@z
4���5DüB�&j��kT"D�iP��1��%�B��.�ҍ��J��i��-
`��=�B�I�Fv˷�[/>�A)�%�5D��C�ɜY�&�8u
�%w�HeB�K��5;�C�I&
����T<Hi9+^�y�FC�	<p��4O35�@1�h]�ZC�ɒoP6<q��Т=�f�a�]#^ЄC�ɢ ^���.��37(�(��|yVC�	�Oˆ�)�,�+��kTU�8I"C䉕*�����d^p�s�nS7;�C�	�?�(AD�ȿ;T�@TL��C�ɤ8�P�A@�#kU��B�Q;�C�		gN��Z��Hx��L�ƏA�,�C�I0U�d����'��5#ȟ�:PC�I�>ъ�!��M5%iL����P *�:C�	QNu95��	��m�D�ɪ|�XB�ɐ|�,x�@X�{�u26cC�B�NB�	�}H��J�Wr�TAD� �"�XB䉩ߠu*Tf�;O8����H��CB�Ɋa���󢌂�qtb��O��C��^it�r��u�(�OM� C�6h}����,��P{���C��B�& ���23o�����%�FH�C�)� �qR��ToJ#W�����"O~��GV[rD�$f��xA�Pz�"O�a҂d�)Y�	�gK�Y"a��"O���'^~��R��I���!"O����O�z�{�d�/V9�"�'��I͟@�I����՟��Iɟ��	2S6�T��A��$lR�΅�<*���	�d�	��<��۟<�I��H�	�����3���CU>�`�(�#��I��� �I͟T�I�X��ПP���`�I�Ȥ��,��9����5O\�'��e������ן$��矔���L�I�t�ɸ/�4P��n�h ��/�������O��d�O���OD���O*���O��$�O����ۘGo�s���:�r���O���O����O
���O��d�O���OXu4��Pg�1��
�R>��3 ��O���O����O����O��$�O����O�p0"��	��]�C�Nr��Z�m�Ol�d�O��$�O��d�O����O��$�Op�S���7�"��kO�[�P�ª�O���O ���O���O����OD���O��f�ʯ��񋏫"=�����O����O����O����O��D�O����O���!+X�-ڂ�X�cU�݅�	5�����O���O����O����O:��O���[�Pe�e_�"�x�{���������O����O����Od���OT���O�.�ddX�� ��6�:��1bV#w ����O����Ol���O����OD�m�ܟ��ɣ:7lxȷJ��8�X�`�- v��+O��D�<�|�'3�6M�<& �d3&
�q9� ����L����܃ڴ�����'"B�_�,��)���]�bY�� )ǘ0�"�'�t�
d�i:���|j�O �x�R�0ŋ;��H���L��:,�<�����"�'`V�4,��xm|�`��D�h.�y2d�iC�t؈y��Ϧ�]$^ �y0� *HЃ'C�2-��E�	͟T�����g��7�g��
	"U�6L���@�k��K�iy�Γ
J�H�z����'�dC�D��d.��yǣT�w��ѝ'K�IO�I�M�w�{���t� �H�����o�i�AI��*�>���?1�'{���y��Y��M�f�%��l���\��?�&kډM)2��|�6K�O0�[�`4�eB��a�
�Kt�Vq�BP.O�˓�?E��'�Dyˢj��\ъDHVOG�MJI1�'�B6-����	 �Mc��O�l�"���1e��R��&vrx��':R�'X��Ƕ�����Pͧ_���DO\r�@E\�&��J�
XӾ�%�������'H��']"�'ވHh�E�{�Ƒ�e����� �\�
�4ubX�����?�����?i���
t��Tȇ�
' �`L���\�i
�Iޟ �	]�)�o���H��T�*������t5��C��UҦ�*O����m]��~|�^��K�Mѫ5��ل�� �\U��N�����ןl�����my�n�N! 5�O����E_a3��!IN��r!�O��m�b�vd����I�����$͹�P��V�P�^l�@�恉]��$n�}~��.<)�vܧ��� a](�zR������@��<����?���?���?����9:��-�S!�>R^�3b'�u�2�'�}�l81��?-��4��p�v��̆+_�aHs�7@pIKO>I��?�'-�H}�4����0�JWUF��X�iN�n����ƦJ�?eD?�Ī<�'�?����?��lI�B�(q�ō�A3�)�G�>�?�����$�զa`��쟌�I�ؗOи�Xa	�%F�
�Zp�L6d�%y�O�T�'�'�ɧ�I�^)��C�ҎG��&�#t�f���"G,<D@7�9?�'����w�Pe�T�"c�-}"�􆐥ehv��I�`���X�)�xyo|Ӻ@�񏟚Zv,y���a�ԥ�]������O��m{�fo�I����lG�	JeNZ}b8���hݟ����u,�ql�p~2���P�����$ݔD�(��܀G�4麃`׸ ��<����?����?����?A,�ʉ:�B�JDF�J�'?�V�8���	B���t�	蟌'?}�I�M�;4d�Y'�oE��t'G�Iټɓ�O�b>���cS���3@&N4S'<L�3�i�a��@SUb�O*=;K>a-O����Op�a��O�q��j��D�x�E����O~�D�O���<�s�i�ƄAb�'�2�'���{�*@4���C�l�h�`��SP}��'tR�|raZ�z'P�郋�k܍�H���$2<H���-�1�.h��(�,����}��)��N���Hh�,��0����O^���O��&�'�?�wB��_a�m�b\9������.�?�7�i-��"��'��f�����7<��h5B�4��*�c�(�������I���rG����'��!�����?���a�\����`��S��U�"�'��i>���֟���ޟ��I��1��âBy:A� �ǣ�,d�'͎7�<W<���O��0�9O)��Ĉ� v��k1��4w���ْ��F}��'�b�|����sJ�"�3��y�cė 9�$m��Ē���/[r�M��� GB�O�˓#�����X�sn�XAG�>{�^�����?���?i��|�.O<�nZ�/���I�1gn��b��$]��1[=�h���M�J�>���?���"ŤgFH�D���o;r|� s#^�M[�O�=PDB	1�B��d��� ���`(z�l�:4c݃_�bcu0O����O��d�O��d�O�?�і�B>>���k�vXx�e$�ݟ$�I�0xݴk��`�'�?Q�i
�'nlb���T�l�k$,�8h��A�`�|"�'��ON�|�iS���EJ0�U�;�$�BDlL�9�p���LF'`��7�ĳ<ͧ�?	��?�FL�h��yelN�A � �/N�?�����D��Ǫ����	��O�R�2vK��W8 ���aȗY�U��OLA�'�2�'�ɧ�I�9d"bu+�mM�|��
���
���3'"B;J��6�'?ͧ�.�IB�ɥ u �T�޹��0j�����ğ �I�l�)��kym`�,A���	�����r Y��8i��G��I�ʓ.i�v�dX^}"�'��30@��v��8�߷X)r ���'rF�,(G����(PA�#&Mq�>�0aY�-{�
cFY'8�� �0<O�˓�?����?��?���)W>G�XkE�V�My�XB������nZ
x�����՟���n�s��2�����Va�f�cC+ݢ��ԘD$�?���S�'J�$̘ش�y�j����T����LC�����\�y�hˮ/3hm��䓛�4�&�Ā��6t[���F�̘S�ӎX�\�d�O*���Oj˓2���&UZB�'#�܀Ch8�(WJ��Ѕ<uz�O���'���'��'G"�i���T5��FF�t�b�On��r��8"8�8%�!�I�.�?i%��O��ZS�5��6���ޜ�ӆ�O��d�O��d�O��}Z�jB<"$đ;td��=x�J���` ��O-"��+�M��w����48�n�Pq�Q�o#�LЛ'_2�'b� :��&��P`T�ۍ?��=|�nis-�GA\�Q��rpȓO^ʓ�?Q���?����?��J��1	�Nϑ�BD�V���|�:�-O�8n�,V�'�"���)�&8ʖn/J��=�m��[�V��'2�'ɧ�O	���΄&�ԅ�`�N6�d�E�["P�L@R�Oh|I�K
7�?Ѥn5��<iw��=��bF�@��Q�����?���?����?ͧ����=�g&��W��77�z%eN�� �D�o�0�ش��'���?���?��U�(M`��mE���aB��{(�̫�4���	�g��}`�Oq�O���,j��9)r�ϗ(�t��eߓ�y��'�2�'Cb�'����B2%��E9���\C $�V� �V�$�d�ON���Ҧ�z�q>E��,�M3J>�rO�$K�&t�'��	=��DC��A]��?A*O�1/q���*��MRƟ�Q�:�8C �qNA+�ϛ�$g���������O����O���eN*m�G$��0�y#c&ِ[�f���O�ʓG�6!�'�2�'��\>�y0*�Ed��(4��:��@rD�:?1UY�@����@&��'$x�9c�����cG�6�|qJ�'�Y�T�۴��4�v1B�'~�'�K�<�����8~L����\��?���?a��?�|/O9n5]�X+ĆC�{��ٱ�[�rXP*#�HuyB�x�L�豮O��$E�I�"���\�dP!�Q<0���$�O�m�i��z��:u���@�O�b�0$���F� LYriS�[3D�k�'���x����8�	���	X��ˈ1숩(Gˈ�/'�Yr����6�Z��l���O
��6�9O.]lzޑ�#�Q�Ov��2u��:����m����Ih�)擟u�fmZ�<�!
�r�8Pr��7��LɐØ�<9�	�L�t�������4����O	%�Ȫ�D:d�F�Ծ�����OP�$�O:˓�F陳Q:��'M�
_g� ����:Gc��P���,�O61�''��'k�'��5jТ_�<rNh�i�vF�J�O朠�I�5{�6�&��k����O5�SD�h�{���*���7E�Ob���O�$�OF�}Z��LFN�9�KT�v�RX*ၒ�,	Nݨ��b��V E�K&��'�6-8�i�	{Q� �s��m������f�
��e�0���H���`� nv~2-ǳY�����G�ո��o�}#�	�P<V0R`�|�Y�b>c��*�AQ� ������Ոn�eh5&,?�ŵiC��j��'��'���
 ���.� �رgT7�d�Z�Ne}�u�4��Ş����"mN%ȰH��I�t�D0�M�$P�,�%�ӌ$�d)�Ħ<�`�	�y�z����VӾr��ǭ�?���?����?ͧ���J�m����ǟxr���=��@A�A� ���w��Z�4��'8���?),O�H���cjɢ�A� =qƝȁ�ɝx�"7�6?w��2�L�I��䧶��B	�1蘨xЍ�����QCÍ�<���?����?���?��T�Z���Lj!̎"ܚMp"ۍ_ ��'���q�~Ek૤<�b�i��'eH�;SS:�i��Q6|ݢ! u�|��'��O��hr�i��	� F���q"�l�����[OȐ!�
#��5�D�<y��eE'z.a�2!��Ths ���O��nZ���i��şH�IF�d@�&]�Z]��,��:\h�0C���$JJ}2�'��|ʟ� ��Ć���9�Ҥul���YL.IC��oӨ`���thc?�L>�1�
AH�C�䈑8�~$�⇖��?���?A���?�|z*O�Dn�C��*FgI�j�Hph4�k��� �\��ɣ�M���>��U��@*���Z\4��S��ZX�P���?Yw)^�Mc�O��P^:�ɔ��� �}P��ЛI$
�F,h���v3O˓�?Y��?q���?������0q"�"��5q�r�R�ʅFK@nZ�
Ƕ՗'YB�i����]!J @��7L7BňP��F+x��I��h'�b>A���٦�ϓX%S��KpV�4�Bk�@�T�����O�"L>,O���OB�J���^l�s婜2�>9)5��O��d�O��D�<)��iS�����'���'�\IR�9,<a��';U�����dYw}R�'�B�|�� vFҁ;��<e6�+���=��$#y^E%'e��b>���O �4�֐����Gg`tA��D[,��O�d�O�d=�缃צl��tD��?�>@�2�^�?��i� Y��'\�o�<���-{�
@Z��1 ޝ:Ӈ&���	ğ8�iyo/)��o�v~B�L0L����#��U P���l�� ���,pH>�/O�d�O����O����O�7�ڂN�Q�VM	 c4���O�<Yd�iB���'=��'��O9�ȉ  y��I�
D*[3��ɂ@R>h���?����Ş��(��P
=JR�3��	݄�@��	*�M�'S�H�& ��4H�d/���<)��=��Й�*�-W�:-��m�?�?I���?���?ͧ��X����P�����] �Ճ���u5p�"���� Zݴ��'v��?��ӼV� tt�9LE#��e�='�0]��4������Qa�O/�O���G�/7�Ukg
u&R���L�$�yb�'���'�r�'��	S8!$>�J���4p�Z	k˖_i8��O���Ʌ
m>m�	��M[O>�� �clQI���+r&�г7������?���|�P�Q�M��O�n�,I$)�E(3=�l��⑸�T|H���O�1�I>i*Od���OB�D�O(�ˣ�9���[�J�Hd9�@�O���<��i��Y��'{R�'"�ә!���i�֝�s�Ք}��U��������R�)rV�P�Z�b�y�F��PT<�K�f��� �� �LiP@[*O�I��?M ��+�����^�\���:|@&�d�O����O���I�<�Ǿi�P�
�F���Bl�E�\)��
��|�2�'V�7M=�	�����O� "VaR�F�	�OXts�!U�O"�$��`�*7�5?�T�Y�Oè�Sqy���^݀���ԑn�pq�R��y�]�d������������ �OU�8���ŠHQRay����2�gӪMi�O&�d�O����$R���ݛG�z�{���7',�Qcn�!+����ܟl'�b>ai�+�̦)�x>�M��)(;��r��Q�G��h͓l��B�C�O�qL>Q)O���O�������l��H�J�-��i�#�Ov��O��d�<�ǱihdLB��'���'3��PW��	�ư�4�?M+�$����^}R�'��|e�$N��SbQH�\8�����Ģ>���Iv�~�l`$?Qs��O����j���s�Q�if��+�Ȁ%"��D�OB���OP��.����N�|�H�X�!f�z�qfEK�?�ſi눵I�\���ٴ���yW3:�����k_�%�L��G���y��'B�'9��R�i��I!S��m���O��|f��Md��`�Ig�����w�Gy�Oh��'!��'����f+���EjE�ؘ:p���X�剸�M�����OL�����^-�~�!��n��� aD��Д�'�R�'+ɧ�O��q�%II�V85`�^�:�IQG@�rɛ6����%����!�D�<�H؁eE�CD�D�I������f6m�O$�$�O�4��˓w��7����,HR�L(��U5F��+���y�j�z�x9�O����Of�$Z�4B�< ���l�>1�e�`��$!w�fӼ����ƣ��>M�]�x� ��S�$1#� h���c0��͟���˟���ߟT��o��B'0�;ä��C��� �\Q�����?�-��&n�7a��I��M�J>��.��k@�\B�	5�ʠ`GlW����?a��|"oى�MS�O$��oN�? �����6#zT�4&|v����'��'g�	�|����	o���Ж!
�B�<$�B|ī���?��������̝Ɵ��I�|�O��ɨǇ� &��q��bI�p�\e��O ��'���'tɧ�ɘ!6�`dʈ�i��Kg��(ߎi�c�ߐt�p�˦���S=!�2M�C�ɪH����� ����CZD`I�I�����ɟ��)�Ny�nz�F@Q�!^�~��S��AR�d�g��$�O��la�3�����5GT(:�Bth��K{�M1CFGvyҭ��;�������-ąI����FyBn0f���"`�Yh�/�yB^���	���I���	ȟ��OK������L��3�t�� s�����"�O����O��?�Q���3@�e�zЁ��a@X�MQ*�?Q���Ş-�R)X۴�y�8���˙?zJ�<RQDE+�y��*!����I!�'��Iß���*9��@ Ѩ�T��Pv���!}V���̟\�	Ɵl�'u�6�X�!�8���O��dZ�,��J�e.�X�"̄=]���2�O"�d�O\�O$���0qRJǢu ���,O;~�	�E�����*|@i%?��t�'v@M�I|�aU,�,XP���Am�<=t��Iܟ�����	Z�Op�ͭ��
�n������St�Ҭf�����O*��Cߦ)�?ͻ5]2�bq̖4?J=XDl՛�>l��?����?�â�0�M��O[�惴��� ��)'�H�l)$�3:��
��"���<���?���?���?A�l̫�$4s�F�3|���D�4��˦�
������I˟%?�	��h��Oq�R�:��M��O
���O �O1��}zS� h�s� �)=�n�Ȗ�X�$���Y`�����(I4JL��A��ty���m^�Z5��#B((kT���0>�b�ix�h��'yLd���E	J������H2sl����'_~64�I���d�OX���O��KF΄t�Ʊ�b�$��I�Þ
4��7-+?q@'U$���j����:¦Q�ժ5���M�iJ=�A�p�P�	۟�����|�Iݟ���0��d�R=���V�T��댜�?i���?�B�i����SQ����4��[ڦ��ׅW�r���+߾0��Mm�	0�i>�YV�A¦�u��W<!REY��è2��g	�"V4�ca�'!8�'���'��O��Kd���˨�B��9Gʨy5���M��n�-�?���?q+���� 
�������1"邃���S�O����O��O���DW~лF����zfCA��lIt�#_�d4lژ��4�:���'��'�<�ꂉƭJU��Q�ꉁN;��a�'�B�'���O��ilZ�9n  $f�:�l0@!��x	��ɡ�����I&�M��r �>���d��hX�-��qHn1�a�ߧz(\K)O��Qիjӂ��꘠tJd�Iߧ��DP�lM8�rTo�w�,��VB��ģ<����?����?!��?9/����	ծ/ �}9r�ĸd���)4D�ͦ!�U& �������
r��y��*X��P��G�3U�I5O��d���'�ɧ�O:~-1��i�$�}H�L �ǖ�C�-"TR7Ee�D�rH�
�'��'��	�����^R$x�dػm;fHBu�8mN�`�	����	�ė'��7-Ǝ;2^���O(�� -�1
�Ĕ20H��ℭh��2�O���OX�O���<"p�Є��wr��F���b�
C5I�d�ZM)擶vԜ�0J��.I6�QY��Y�''����ѭF�(?��M�ev��c���2�3���ϼ���f���x����#_`�s��S4֘�T�D,�m;�
��{�*Z6B�����˂.V8�A���Z51�fa�P�ș`��Q
�^�������L�Wi�&�ȡAu�_?%�6��шÏL�.1�j�tM	a��*lTAP�ǄJ�Z-L��4
D(�Xت��D�z��hb$hM?�x�!"G�e��+�4|�:�1 B�$T��R�E}��JC�ڍ�M��'�Z�h�_�Ȕ'��|Zc�Y�FP_��ic� ��-H�O ��n;���Op�$�O��KzD�
�� !R%�	y��u�&�ք}��Qy��'*�'���'������wX�x���YQT`G	0H2R�p�	̟L��Hy�7D�p�S.��l��� �d�I�⊫u)|6M�<����?�=j&[�'���w�[*��I�͢5㢽өO2��Or�Ľ<IQ��C
��������m��}���k����f�0�M;����?1�M0�T��{��0�U�&j�p��B�Ǜ�M��?�*O�!�a�G�T�'?��O�8l1"�H�:8���Q#�pXZ�Q�I-��O��d��JL��h��z�xɡ'�'	o�-i�)�1x���mTy�GP�NT�7-�O��f����q}Zc,�py��ӾY8���$ГW�H��۴�?��WJES����Ƣ`d�5莦s���"���	D�*�# 7��O �db��)�`}RP�� ��V��P���&��A�:��pcY+�MkC�%��'��:�$V�
�މ� �Hr6��&�\��l������<���1��Ĩ<I���~"P!$���' 3�8� �����'�T��|B�'���'���P�$�2���$㌲Jc<͉�kӐ�	(����'���ğd'���&�5�BꅦIP�R$+�y���g88�zH>���?	����DL0���PB�0=
"�����m>x�B�	N}BY����J�	���I�v�������DV�A�,�<�.!��c�Z�ӟ��Iɟ��'�bE��r>@&mПZ�>�[d�	�L ��dӮ˓�?�I>���?)0�� �~2����S�42��V˖����O��d�O��@����R?]�I�A�!Y��D�N�,{�\��@h�ߴ�?�O>���?�'�DB��X�+���w�����hif0l�ڟ��	`y2�*\���'�?ᚧb���$�l:��"�&�B\�e�'E2�'�-����?����^�ԑ� ��J00�ǯ�>a��Yi�]J��?	���?Y�'��� ��s#�R�({��	G��CG�i|RZ����K'�S��'G���5	̛]��e#t�R��6�_�S�@��O��D�O�)�<�OF���+Jo�-Jߐ��#�y��,l��Ex���Q~!V����-���
@O t�$�o�����ԟ�A�G�dyʟF�'�Sg0����!댝)^0H���"V˱������� @s��1җo1nd��v�L�D����˓I���N� �5L��K�T0�%B�}���t�x�͔;��'�r^�D�	� I������?a\k�f�15D����oy��'V����O��I�z���z���m�ܙTi�$i�7I�"����(��ӟ(�'=��@�x>���Lm���7�A7�`m�0��>����?�L>�(O��O����	M@��mG�`/�=����l}"�'j�'��	�]��M�N|be� �س�*Ʊ��(R�l� B}$c�i���'��I˟ؗO��Z>�cU�ӳF�4(���X�p��Ǭ�M�����O���ɹ|����?����qcR�jd���ͥA�"��H�b��۟@�'�m���f��ūF�6/r���9zbX�Q�i��Ɏy��`��43���۟L����Y�����5�I$v�m��!�^ۛ&�'���'�bi�~�-O��禅�fE9y�q#"��a�B}9�Hn��)���O����O���^�S�tE�)��j�DDJ�,ec8��YN�Ex����'��5���$������2�h`Ӵdi�|�D�O��d֋o�f!�'�������9��ň_�#�~���.�K]8oԟ��'�*|Y�����O��D�O�� UG�Y��%���)�� �B�M�	�z��u�O<ʓ�?q.O>����{�,q=�)3F@�]!��a[� �aq��'V��'�1�vUBņЭ��$�㞈Vؠ�5���T����D�O˓�?����?�%bXV�֔����3��k�es�i͓�?Q��?i��?�.OmёD�|���v�T1+D��6L�YrcZԦ��'��^�����\�I��(�i��0�GX~hx� �C���@�>9���?�����S�2y�O��Gع[:̬cd���lW�kP��<t�,6m�O���?���?����<�N�T+�IN>���J��H�gӶ��O^˓$��W?�������#9ʆ��D�H9 �l�aAH9c�6h�O����O��K���<�$�?ݻb/�(��I8�hQ�j�Z�HF�l��˓X��Q��i���'��O�Z�Ӻ�U�7\���.���9�d�Ϧu���PЍy�X��5",�9`w�D�7'�D�'BKF|7�»�P�lڟ��Iߟ��4��D�<�@���K昗�l�d4�)P�$p�m3�4/����?�)O(�?��	4s&dd��A4_�8y�3W:J��ش�?����?IT�ɕ
�Ity��'����[a|RQ��.`m��h��A��f�'(�	Y0��)���?�O�NzBlY�lR�9�b�> ��4�?�"��9[��IkyB�'��	�֘1�>��aH�M��Ai`�,gOr�������D�O����Oj�'H�S��H{ڀ�X�يrx\�񄏎���<�����$�OT�$�O�G�M4 -��R*Zg��9�K��l��$�O(�D�O��d�|Γ!~@���>��ey�2i��J��kX��&�iG�	���'F��'�2�'�yZc���� Ozi�Љ�5)��UH�O��$�O<���<qS�O!�ǟ�ׅ=܌
Uʞq{���d��.�M�����Ot���O
�g2O����@x���k�N5��Y!/$�)3�~Ӏ���O��E�.8��\?��Iɟ��ӂg�Xp p-��O jH��΃-�U��O&�d�Ov�d���D�O����O,�S�F4��2��X�@�!����}��7��<��L.���'>��'�D��>�;m�n�hp��7X�I�c�29 �n��|�ɀA���	���9O^�>EZ�L�l�����@X�U@��MK��ʁ5��'���'���ͦ>�,OP����v��s&@Z8��hj��ڦBt�o�L'�����.X�8�m@8j`��#��֘) 9�Ƶi%��'�rDƥg"������Ob�	�9DizE��L5�Rq�H!:��b��b�'�	ß�����%-�{��Y�P�&W� �Lݟ�M��84��T�ܕ'W�^���i�� ��� D���-L�,����>���D�<y���?����?�����66�#+Ԏ9P"��$(�0��s�a}�Y���	[y��'0��'�r%�r��K�DTۑ��F���	�E�y��'+�']R�'��	�vu�%z�O��,�aJ���)�z)XmZ޴���OR��?a���?��OW�<)��_�{�P�D�--4���]�?��f�'��'��W�(�R�=����Ok̄�z��JǬ۸\��л��C�{�F�'����I����cp�ԦOԬ�#A�"g̈�n	�B�)�U�iA��'T��"eT|�H|
���:#ɓ���c��C�=Ӝ(�$�]c��'z��'�E�!�'��'��IJ�!d�y�Ӫ�,���b����&T��X�gV6�MS�Y?����?�x�O���f�)��s��Т� ��i���'�d�Y��'��'/q�HI@C��/.f�h�dXJ�y+t�iUN �%�o�\���O������>aCI�[�T�s���9L@��\�|���?M�|r���O�s�	-Xhh�4�Z�jTaL�}�I˟��I��(l�}B�'��dF"fP�y�E:p�R��"l�.x���|�� �.�����OL��1u^}P` �R,�U�!�"���m�꟠I�����?I�����+�jJ�'1�m��A�)C?����A}bKO�yX�X�I柨�I`y�Ɓ�Պ��ԫA'K_Vpy����a����(��ݟ�$�`��ݟ4pdB|0|8���=8ѳt�ʱnV���	cy�'�b�'��	�����O^:eK�h�^s�51 �54��1��O����O��O����O��x���O��+�fA�u�.jԪ-����=v����?i���?,O^MbT��uⓂ,�$�Ħ�)8R(ak����# y޴�?�M>	��?9F
(�?IN���b��e��тFmT�@<�T)�/s�����O�˓@N�\�e����'��d�\:
�\ihg ��	�����C	Oz���O^ �g�O
�O�S���R�����`I�-��6��<Ag��������O���PD~
� n��QI�~�t����W
@��i2��'� Ii��'�ɧ�Od��(�B�	7G6���S?Fhi�ڴ#�>�׶i���'��O�b��(����h����e�]4L�Q���Ĭ�M3�)ȧ�?YH>��T�'ܢ�+(^Hz�Ĉ>S�
A�Um��E/�&�'N"�'�|Y4�%���O��D���J��J� �2H��7XW�y1#�'�	��@'�8��䟀��?+讴j����NȞ�PP�U�}0�ڴ�?Q�B�e	�'���'�ɧ5��S�`�CR΋.��dⱧ�!�� �e\:�d�<����?1���&\���m�&�ެ�U@ůkH��%�q��˟�IG�˟��<"��ě*��-���J�K�Hc���'f��':�OiN �"|>集�,��1�僉2hu��2��>����?!K>���?	�B�<a�D�L��l��/LElyv�C%K)����\����\�'L��(�iS!)>-�3�$W��(�i��xDn\l�w�'��I쟔�����`6x����PO�$����<rԜ�=9���OjU�D�6�8�(4�D�G!XȈ�"O�1Q�$۸s�(�	�!���q�O��sW�V<iX��Sc�Q�1E�?}��C��-V���g��q�i@�h���(�O$P�e�D ��kE/�j�����$PR`t0oM�\�
��YP��犓)$+T�2OVi����%`��Y�����u%"�jG��L��KD��R7�@�d���?���?��u��ΆD(8��k���@V��"3�AE�CP0ٳ/W�d��,X1�&擝���|ɲx�'�0k��t���$���/Mڸ�E	@�|��q����''�L8gt��a�[��4����]�@ ��\ӟ��'0�@���|Z����y��a��E&'B�H
���y!򄁓�\��"Ɉ�h���QQ�P1	s�I��HO�Sgy�*�2C��H D��[JD�3IT;:�:��d��P�'���'B��]П����|j��NL��9SP��'X�JX���+�a���[(6����'�H��eӫ0���ZCΜ vI�O 5
5�=r@�<���D��G,��ba�C,?tD�� .��:��=P��'��Q�]�$���F�lE(�˕�"Nk�}�ȓ<����"�
�0aя	�<,��<�&P���'<�M� M�>q�^�bъ�9��aŊ�4|H%���?f��?������o3UܝÎ���t�i�.a��a��2`��*5pPI
Ǔ/Kn�!�H�v�:@ɂD6�M��
R����Ao�������Q8����c�Oz��<��b�)vW������
/�FظRD�r̓��=��*c���BSe��fH�(s
�k<y%�i���Oӿsa$��"f[��]ɜ'�ў"~�d)�)�E�1E��i�h����]�<Q���!YG:������xl���GNY�<qd�)K\���Ld��@��~�<�#k�jg4���%=;%���1��y�<�O�\�L�"�H7A�����s�<9�A�2��(a�2 ��Rx�<!V�޼�nl[Q�oő�P�E�!��ܙa��`S��I�k��ٚ_S�!�d&+؆�JT��:��(
��
u�!�DC6$� ��4�-GE��� Ρd�!�DY	m6�+g�%\%�}[��̸w�!��/o�U��[/L����P�r�!�C�t�=��ˊ�[,�
S0O�!�D��`����A�R;P�؄!�q�!��,7�¹��NR5h@nh*��/q!�P�|��$�@����y���2c!�ҧu�>p;w�T�Fy��`��kL!�$��0�A���];c,�%qc-��!�$!"G0���6+�9cU׭]�!�!l+^bD�=�H��dᆸ1�!򄌨q��m@�.��hip��A�!��]��y�ώ�F����e���qH!�dM��X��W	S�P��@�>o>!�$�H,B()C�d8�EH�?i�!�D̻!.� zF�'h��"��;g!��A)n���
[�)t(����5!�$�,Ͼ!��mR�nt��zP��2#!�$J`�j,�Q��:��:�i3!��3aYF���✢%D:��pIݺ!�d��I'��i7j�W�M*�N)]!!�� �iB�8l��6	�0�,��s"OYh�'��2����j��HTٚ�"O<��Bt�����ɒ!P2� ��"Oje��e�*/Q�i�Ɖ@�6�x�"O��iD�LVl�͒c(�R�!�"O��S�B߁.�̨�w@�>:	�d9�"O<,��ǴC�ҁ0f��6|���"O4�����rh�x&%ǫye��1�"O"c�e���	¡�_V|)�'>�AB��!��X0�B>l��x�'GDՃ��W��DA3�J k����' ����fU?4P�+��J�e��Q�'�@Hq��%<�n!3�a�OX����'!hI��!,�Du�d��>��|��'Ĝ]iħաB��@��NǠ-l6A��'�U�`�ڲ8��y�C�����ٱ�'��x��[��F��BeN3uP%z�'�:p �MF�}�8L��f�}�����'� y�veWZ+��8`�,#
�'���ꃦ��e����]�2�'���ƫE9	ݔ�(ԕZ����'�\BզV� Y�qkS�ߣ~�zDZ
�'Id�s4��J&/�#yM�X�'T�Tr�ի"�BőFآz� �R�'���Ӄ��!�4�[v��1y� �'7��
S�K�pI��+��@0y�:�0
�'�d��U	��7��\B���q.Pݐ	�'�d�RF
�_�C�ٻez� ��'6h�hw�F�o�@���
�aG���	�'��]�"aR	5�:�ɴ�K#n-H��	�'P:��i���01K��q�n	�'y�]�%_��8�ۄ�Y T�@���'A�}�N�:	�j�CÊA���
�'~b0�G�7�ޘY��9/6A	�'W�EӵJ�,I8[�+�1��%��'�,�)��/bkxZe�ǥ��P�'�^�B��yZ~Ш�iR{кŪ�'>Iz��KZ�.����v���'�E�V"1�,�3�'|�Fɛ�'mh�h���&�(ab4�_�b����'����R �8�@p+�o�$R�TE��'-N��D>�����4	�'_��a�*Np�P���W�B���'t��
c�W�X��$�6g�1��4��'�B09�/�t��)��Y �R��'"J�K��՜^&[�HZ1#0vŰ�'ޒh�b܂#tx���3 ��P�'ʸ}Q���+N���1��9<���'�pB5퉤����ٝ	꾄��'Ǌ�ybf�^_,m*�F����')BlQ4BE�!�*�@WkΧ�f�[�'�Qk�^9XU���6�ְyR���'��@ZuhY�
"�,�S��$o)�P�'Ru��+��� ��-a���!�'�f�1�nRg�!H6)�
XjH��,-$!b1�V.HK��Ҍi��B�	�A�`YB3�I�I���a\55lB�-}|9�l�+DXE���$Y6C�I�0Aɉ��A�{�4����P��B�I�DL����כ����-��`��d���v	��~����;U i�O��0}8���Bq�<�7 W���A ��F�P(xn�;�p�ũ:��Dѫ0|�?�'8)ٲ�ۛ{^��T�DMS�'�m�4cL�U4��F�*>�� *d#���ƅZA�_a脭�W�9\O� �<y�,@*�M"��{k~t���'�R��$ePU��Y���/Ӟ=h�gՁ$���hG�I�&@!��P�y��?-0�<Ӗ�
�wt��@C��$�5 o�C��~L �����'Z��?5���-KqvX��.QV0�GN;D��[�a�*[<
d���Zo�*a��
�U�f����P�Z��6�@lqP �|
�x��G�6�2�A�E��!.>�p׎4��╢��y��\7
�^�:Q�p.Ϳ? �����0#@<��Ig�����'�J�J�/f����Z�pޑ	ÓXT@y3��H%$U��Y��(2�`$��OU3]g�Ts�@'8�t� M�zTB�07��b�%9).��s
�:e+��
�R]��5JVA⎀=!��t�)�=}�[K�<Xb���O�V'�C�	S��X8T��s�8	U�A0��p2a����
�3��O�B#:�e�kv� !�!!O������y�|���+��!ӓ���F��(�
��$)cw/�!y��9�d
�b,P0�EF�6w�����6j^dлu��a��Ĩ�ax"�΍g��*��U�F��co.�bJW/b�BH�1��!1�!��O(<iS��C�n\Qk
-w� m�'ŁC~�,�4f�`�G�#G�
Y�s�ȭ�?�}B��.A&�t@�Q�d�;�bS[�<Yq/�E{��ɗ�Kjِ��ܱUw�,S�o
|X��/J�I~�P��/B�<ͻo<�֫�/�����j3.�����F�<�g��Np�8G,4�E����9N������3Db�D�N�oX��c��=�hO���B�a����IԊ)s8���'����������/�+&�*�B)�&N���ɗ�D,U^��yb��h���D�8�Hń�I6f��r����i�K�o�c��k�[�/��da�aNH��Q�r�,��`G�?Mq0Kĳ/�2x���]�p*p)Q�/"D�̈�� V���*%��0��@�LѬh(�baaK�B�p��틄�p�.I�]$��pc'�/u�s��@��B�	:A��CƎч����<m�����)D��}���Ly}�K�A�g��&����#h�$2�t�Pq��0,�*���	9
�h��PM�6�Z5��X���
��G�bEx��f����ы���@��D(P��-v�0Jt�hݥ��' ��O�xP��..���� �ۃf�U��k�ႀ��RP=*Dd��h���YH��)�}�(�XT�E�������D�`��� pZU�P)m������$4��h����=j�E��dM�{L�L@�`��a�,9اJkVd����TMfi,O,��ߝ��E���AR���u�����"����j��v�ʄQ�	�u��d���҃j�6�i5�DE���'�:�S8%p|Rs�Y&k,<��a��6S����&S̄4pS�S��6��D�'L0��]�	r���g	a�>E�g�\�nᆸ[W#$���AN ߟ��j��U�RA1F��_d��c�L�!�X��-ǐ]�"	�3n�"j:>P�IY;��Tt}�F��6�����KA��lSBA�7J�(h�'v�Z�MڛJV�2R��9ċ�iG�eZ����i�
c%�{�_������a\:H(�4�T3@ ��ȕGZ�Ƥ���r�F�k(�i>��/�h�qq� 9rԡ� +��y�.C�I���)��Qx5�%
��Э1�p��Dϻby�Op��'���� �7��'�r ��"&�p�Gߖg8�X1
�b��q�O϶'��Y3��@ G[�
sm�=Bn�7�ӷ|7���ck�l�C��{D8|�s+�.6��?6ņ9�l�C$��|����)�s�	�U�����!� �l�q�2^➔�`/^5N�5�aϘ+M�Q�e VOv�T��	p�ʡ��I<C�R�Ћ�5����
A��1 !�A=Q����1uf�杠ti���.X��@ �C�L �B�I:+������'�L��K�#y�mq�B+ߙm�~��Y�E�ؘ��!����<.0�#ף�)�@��R;���W;�4$�2臅p�>�х�iF��Rֆ��s�Rd�Aw]�5�blX%�8�:s!U&��r��-OXT�c�K7+B�Zt�ǤL�pܹ2�x��B�	x�wm�
��p�bM���'Q���po�;/e,Y�$��UZ��kMHX(<�5'��W1f���n�5&�j��f��B)ykF9l�Yaf��j��n���{��H�zN�sqf�3L�v���̎xH<!� ]!An�PQiR�h2�q�	�7V�O2 ���Z��壦 dQdu�4�>�q/[0$@6dYQ��:P  "'QwX�lʶ�Ra��%L^�.��d	rʇaޞ$z���]����C�2!��}��Y�자ر�ߘzd ÓqR��\�r�@��H�C�ƹ&�@���0aR�qQ(^�b�6��W�,��.V@P�P�*NP����I%n4�`�	U��8�!�گ^>��Pl�H�|�%���\���蓪JE6)���Rx���w���B� H@�M2��[B	����'蒄�JͷO���
��� _�ҷ &Y�(�}%��)O>�l)L
&�|�I+O.Y���ȂeT� z$h�*MS��#G�'Բ!x `�
Ӵ�!C�5�� ���C'X59:B����N
8bhY2�i���d�{����a�\���O��㉕-I�R%�V�5(l ��F�u�l!��P?yXؐ�#E2��Y��p��,~`P�@��AHԚu�I*�N ��I#�| v⃑\��H0�@�� �4�$�! �>�g�$c�h������|�'���RE&l�v0�Ńց! �-�"O����bR�m�,ts�H=v~6�+���\�&4؂�R��a�oß�p<!�f�'.Dr��Z�(�4�!�\[؞X�����D�iGn�:\ ��ġ����s�f�'V.��� $�(�Y|����I֡;���q�-D�̠0!��e��r()��Ď��B��'�<�bg�a��H�Q�K<m��C�	����� ҅(�,���
mپC��uY(@BwG\�O�¼2P�X {��C��.L�����N�`���k �7ffB�Iy� ��R�@�/L��iŀ�Ki�C�ɡڮh*w�ּ�r�8�@�F�>C�	�c�|5�5�4�P�����;R_<C䉒�(��V�21xV�i�
_��C�I�UCh�`FL�#[P�1�Ȁ4'�C�ɚ~x!cTCRY��!a�:��C䉓1����I�*u�t̃�I0��C�	�?�T��ɐ0�|�T킁lfC�I�M�l4Y�+��0��'�
�NC��D�@���f&�f��6BC�*�<C䉄Qq�t��D3j�=���"BC�Ɇ|84M�CA��[���N0B䉂Z��Q�#�[�@�nAp�n��|�nC�I�G`�Ͳ�`؞
�������U�6C䉾o��(0�E>����B�k��C䉱;�~Q�J[�}�N1Sbo�q��C���F�ǣM�T�����0HI�C�I�EvTomR2���:$`�(b�C�I!�B�B7I&7��˛�t��C��0��z���'qJ��H �	5��B��pN��	�`�-6�x���Y�S�B�5*�䴠vG��{�XUS��Ӭd�B�	!���B6jL%�-
�,W�f	B�	�R0��{#��;gf�1��԰c�C�0e&�Q��*y$y4�M)�C�Ʉ[L��e��z�<8�V߷��B�ɤY��t`5��,�2�Q�\:،B�ɔ�<"A����bw#ٗ4-B�I�b� Roأc$8,�w�֣)�C�ɾ:f\�cW�ĤyG���'T��C�	�{,�U�T&C�Lٴ%���Me�C�	�.�F�8b�:q�jr!��2lI�B�	a=�ܑcF��	�JM{�EH|TC䉉7��r���M�D��GA�6C�	�]fઔ'�-J<Ĩ�C�\B�Ƀ*P T��5�����EJ1IHB�I9IV��R�F�,MOօ�2�	�3�DB�I�O�4�s#�,/����Ʈ��3�PC��3hi�q�ɗ�\N�}� A��B�	�~�9��.ЃH��4�M� 1�B�I0o�0"EȩB���7o 3vB�ɗ0�d\�T.��f��Д;�B䉑A�h{����8c�-͊;XB�I)6LRn��W����R��g�dB�I6����AC� N���A�oX�`��C�	&Q��q�'�RU�	�CӚEz�C��Ĉy�
�&^�9� �-�B��2h9�<�� @�
Uf��MʞYzB�ɘE�)����!L�p��'hTB�	�)�l��2�QH`�ăÃ	K?"B�)� ���q��:gHUQ��Ǣ��a"O���%�ضY��У�<i�Nq�"O��ї�^ RȰ����M�z�d�*�"ObD�ȊYmn�!��`�p�"O�Eh��E L]2p�<^���Iu"O��R&p����lКg�� ��"O9���h��e��Ƕc���P�"O�U⢩�yb����Ɖ7� "O.��EIa��y���oZ��E"O� B!�A�p���(q�#G����"O�Taˊ��k����0;�"O���S�UB�Jm�FϷ8z�x#"O�x��F�K6^`�P�K�B�P 0"O�<��n��a iF�_�k��}�"O���2B�Y�8$�t��!V�4��"O� ` G�B��Q��"�p%�"O����M˔y��E#��O;�V=JC"O�dH�a�!��I�w+C�Fv����"OL�P�U1}m2��kQ�q�1�"O�m%
\�,&m2e��0m;�"O5[&X�rg�}3鐶o\P���"OX9S�� >�8�&� �%FF��"O>����:$�l���׆R���E"OjC�EېLS��Z�F�`��i�&"O1 �7P�5�޷'�m81"O�A{�+42��T �����`"O���GM� g�h"eG�B��,Ib"Oj5ug�:�Šw$��d�\%1�"ODI��耲-�i�!c ??�tx�c"O|y��F�%XNyJ��� ��"Oj�ᔃV{2N�kE�"�<��"O�`k��
��E�B�<{�F�c�"OL9p7�?H�,���I�[�.)	�"OP�H���ltY"�Ő![�,1""O�(�7K� �����'��{�"O`�4�܉M���¢LIU4uR"O��+fm�V���A�K�o&��"O݉��X�6�sb$C�L��`��"O�����݈k
 �B7�ڎI�x�t"O�t��K�o�;�ț0��Q"O�u�/��T X���#��A�"OFh� ^�[�2-�S�{��`��"O�I�d͙������&�"Oz`:v�U!1�px��c��İ�"O� k��v,i3SE��3�浣�"Ozc��@l��K�d�/z����"Oԝ1��6��Ms5�V�{r�cD"O��BA%Lp�.��"��Y 3"O��R��V)<M����S�	,�"O�I�TiK b� �p
P��s"O\A8E%@; �H�)���!r�$k"O E�rDŻw
1��!W��t"O~]�Ql�"�����L�l����"O&��p�_=T.��@+�,l��9�3"O*¡eE�eudD�0�h�2"O�!����4�ʭ��pV���"OV��tE.��S7[	+H��""OxA�²<��1jQ
�-	(a�Q"O ���햗r�j�)��P�*��"O~x�r�-O.��F�H�Z�~��"O�A�S��
Jzfy�a-;_�lHr"O��j�:+Ya��W/ ci��"O$�ГF��:Z�k���O\�Dx�"Ova@c�'Y��ah��PFU��"O� �U��S?P#`h#qҠL*�"O������i�v	�$.-L���"O|�` ��Vy:� G5&�RD�'Q�صM��/���1M 9��J�*(D� SD�B�F�*w�\'d�$��g%D�ĳ&��o (5�B'=R �-�f8D�,
�I�!!h-���<С��3D�����O�v|>�K$��Jvtu�R�+D�$H���d�d�SÅї$�j���<i���ӆ:3��i��5����K߅kt�B�	����	�
���{���BfB�/A��`y�Ȕ<#��8��S�i*B�	9O���g^�g�,�e��0QB��pK�)��N$��`�Ϙ*f��C�I
J�H���l��!�X�����e��C䉙�N|�QK,��aT�8FtC�I�* �	E�Ɓ�A�c/RG�B�	�_�vM��n�:�A�ʽF,�B�I�;A1A`�>w7���"L�:��C�I1@������:D^��J$@��h�B�	.?�zY
Wd�r��L�� �,��C䉱|���p�S�z\!��.-�C�Iq�&�8�d˘_fhp²��4��B�I������,r8r%"��}�B�4I���C��`D�t�3ԑP�C�Ɏ%�|��"K�?..lLR�k����B�i!b�Ӣ�M�L�\(�Rˈ2U"�B��`a\Yj�钂&��$��fJ��B�	� sf�ɤj�&��H��I7��B�ɋ(_���O�0�-�CF�hn�B�	�*	J�Z��D佀�#�vB�3UR���دf�h+"�Q�hB䉋Y����b]�9�hx��͉{�TB�Ik��) �A}^D�p�ϝ1�B�	o@�D%)��#��K���C�	&�.%��*��Rc'5|�C䉬2�l�iB��
b��MS� �H.�C�I�Z�#B#�r�J�9��C䉆�d���\�!g�Ѝ�C�I
��x��'Ȯ�h��M�opDC�	�X�ɀ�}T�If��B�hC�*���0�c�	U�*�*V�L�
C��"`�Y�Q��>ʼ`b�!��._�B�	*;�}�Qj��F���Y�DH ^ɚC䉺b�H��uM'~ɐ�i�)F8�DC�.]���)�#ڥv-:Y���7??C�	7` b��!@���`u� �+��C�I6k��<��.׆F�&<���{�C� y>
���Ar�JE�̞98��=q�'c$8��FꞲ*���qW'
�o%@%�ȓ;b��pM�%��#�բa��@��PpR���!��M`1,F��!��UHv`��I�2\��+Tb��0#�E��P�)��F�2x�>E��b�:Ї���!��4`�$��+?x�I��
��tXtǒ,7R��1�n��8�ȓ
�:ݘ�)��Dk�͑�9T����ȓ#Ϧ��EL��";(�q �V+�����Gul�3� 'I����(<���ȓ;'���Ӏ��<�$�Q�W<`O�	�ȓsZ��1��y�,� ̑H�V̅ȓ(�*uXT��2��U�!���6��Ԅȓ_3�	!+�c��A��AH��X1��eU$��� �'����	X1C�T���S�? �-9ԅ�*|�*<A�ӛ&�ȕp"On��F�ۧG$�{#g@�)�F�)�"O��Q�G���l]�x� t�V"OD`��JK���B��	�N��f"O��y����?�H1�%ȇ4?4��v"O�����
@��d"��Y<�5q"O`�P$	%i7XP�[��2�"O�;[r�9�o�%Q�d�i�D�?�y�F�}���"	�FӞq�l��y��M�N\�rIS��Fk� ��'���-ȓi��-����;?-��'i���da�(~پ���E�
B�u�<!��N`Dܺt"��e��0��[�<�Ř�Mj�]+6�<��%v�W�<ф�8�NQ��V����T�<aQB���c���]��j�Qh�<��:���oY$oL�AB��\�<6�	�~S"eY��Fb׬MQ���~�<٣�]�cQ�!�q��{Bi� f]x�<�p�@�U�Y�!؇+���`���o�<y��\�3#���C�8�v�2��V�<�e �&O�511�le#VaO�<�5.MY�R홲��2`t�@M\K�<�&m���`�� 0q+�QL `�<!uDM�5.���� m��*�.�X�<y�d�wS4��0�ƒ8܄H�!C�X�<	T��Ymh�8�A\�d���ԏ_�<a�J���,8�EJ�	�́u�t�<	%`4")��괯��H�yejn�<9eA iؼk�`B�3�:�ˌh�<�Qg@�Y���	�~�� ��dHh�<q�AP�X`���(�mA���l�_�<�2�A	>ۚ���	ه*\Qa�"�X�<ACO\�6�����ʅ �ؼ�Q��R�<IT�ݨr=8��%�_�ɘ%i�
KM�<#��� ��:�%��*6��F�<Q�U^kj087��g�F�I'�>D���8�Z�kV�� ���l(D�({�
R�¹RA��? t�*D�(:�GE�{a��EC�g��D*D�I��7g�j��^,z>����)D����.ܘ� q��$:>T����)D�t�g�L,~.���O[�Y�*� �d,D�<3!VZD?v0AQ�<D���c�w�0ك �>T�`B%0D���p��5g��"��4"І"D���Uo�Eh4K�,[�Ҙ�!h"D�dP�L�4r:��IUFʷ=��hs�c;D����MD�?1�y����%�p��%),D�4*T��<' ��FCZD��u�&D��g'�Ui@ܸl��-�<�hR�&D�(X�B4{��` b@h��*W�%D��GI��w�А�RD�a:c?T��/�������sr�"O.	����"�@���'!2a`"O"@�����Is��&��e"O
����*pZ��͓�e��(F"O�d�`��Q�d����DȆ��4"O�$8c,�2k�je���&k�`�A"O��vl�0+ݢ-�Ś�ʼ�W"Ob�p-��v�:$���ה{��Q'"O�au�G#N3p�U���7�|dK"O�(2��]; b�䳐��	j��6"O�q���90z��(ƍɺm�F��"O� P���d�!�n�!J��9� "ODb���ݳG獲ak̜{�"O6���f;(*(��ǉ1�1Xf"O�I��W*H��Ȁ3Y��1�"O؉�G�ȧ0*4@$L4yW���3"OD�صdF$�L�3󃃙?��"O�cU�_/P:\[���E4�89�"Ox�����p�D(�w���YL�
�"O�t�S�0�h=� '[��F"O��hn&=Xd !��IK��;�"O�D�B=]��$Ic��Gv!�"O�͛f�S�K�r%����N���"O��O"�A��Բ5��]��"O�D{7Ɖ���)91�ҳh0�0�"Op��G�m��l�H�(�����"O�ъ��ԙY����pgB�s���)�"Oh,˃�� �Q�����܆Lc"O�$S�ꃬ*Ʊ�į��(6�q��"OVb����;�̛Ԏ�>a+��f"O�P�L�"
��y�k>+x���"O�J�fV�)� @s���7%}�#�"Ol +�8��@�wȋ ����"O>�p ���2D<`�c��8�:�"O�0 ��í'e�e�Ɯ���a"O�������,�,�f�\�N�R%��*O:��H�$("\��bL RL�!j�'44P��#U�q����璻EQd��'����3�X)=D�"���<��
�'�n�A�Xm줘���%���	�'��Q�
�f�lI��� ��-r	�'7%9�G�*w�$�˱#�1j��] 	�'�4d��̗-�L����L`E���'+���`��51�����ZbLH	�'�F���$܂<���@��!R���'��]�JW�H[�\Jf�ޡҌ���'�z���/��3�	�ϗ�<L��'i�-)�Ϭ"�����]���)	
�'���S���_h�7g�?�����'��miC,�RB�	KKujR���'vP:�!O��E��N��g�I��'ZF���
V��"P'@Y�x�Ҙ��'����0��<��p�Ct��Ը�'�,��FjZ�g�zp�Q	v�����'w�m! e�=;b�@2Dq��MR�'�	��$ap��O�
W|ވ�
�'���($kO<�Ĺ�p��#S�.��
�'2D[4Ɲ�*�i��	�w�X���'b:t�Qo�q���Ǥ?n�BP)�'Wz(�RI�o��=ۧ�B�s` �'���"4 �(�*U��	F�d;�r�'�ڰ��L��PE�1c�z���'L�� ׃.)Q(�`��Q��(j�'��,(Ԧ�aG����E���C�'r�X�&�;l%WK[�r*����'\<`a��0���`�iE54�*�C�'�PY	���Ea0L�C�0[��i��'E���aDź43��� ��c�Ly�'�A�@�P�]TZ��'n[�i��Ui�'+�uI!�B�@�y�.į_#Z�C�'��q�m$��7N&(�
�'tt@��iɺ�^'x����'�H�O�0b�&���� vG�Yc�'�V�[jҝ/{.4�f�gc2��'�ق'��-[�n�k脘n�*���� r���
cnR�@��^�&�<JG"O����X9����Oqܩ�""O \:B��1!��*7�+��us"O�+*W&8���S7�O�J�H]Ӆ"O�A MJ$��p�e'�R��"O ��r�X�}���+:LHi�"On���-Y�"�y���â�bb"O6,��
&4��`�ЬL�<�r�"O�@��*+,��J�
�6��"Ox�s%]�ڈ2�%� �"��q"O�L�����*�H�(0�X�/�B���"O����f̔n�>�(�Q�<�|�["O��cgnYQ� ���+E��HX�"O�D+PnËy&\m��mO
�&�JF"O*p�ԣ��jk�,DV�ԓe"O� `GЩ����pM�6o����"OF���*Z�p8�(RBք��y��"O�H�0�74���ʟ!�� E"O�4��f �x!�,�3��$�"O@(���1@x�P�b��v�	�"O��;W�˺j�A���x����"O���rث��D�ъU���"O���5��_M���KU�uۮeY�"O.�8t@��=��@�\ժ�"O���"@
;o^|1Vɜ�J]����"O��� K�3�xPK��_<��U�T"O�y`��Lt�E��T�Ѷ��"O�DYg�C�m[��c5��\��%"O؍� BP5����K���YkP"O��ѢCo��q� �$�Z���"O�D0P!_�l*ZY٢�վl�y��"OJ�S�f˨;�D3d�,�.��g"O>�A��l
��5�(J�T,ã"O��p���a| �GB�����"OZ����,�LU��jֿi�2�;�"O���fP�[�TwK�v?20{�"O؄�6�2<o���oU5(��a"O�,�F�3.8Š%O
w@�!��"OX�8u�&&�
�Y�.O�.0�:�"O��r1ކf1������u���X�"O��[���F(�h��Ŗ`�t��7"O��5m�-C]H��� L}��!b"O��֤-Ql@���Ln�uw"O��������Y0�EܖNj��&�|�)�ӯ:5��ōB�k��D�d�̭I�BB�	�~v�5��H�3$�v�%L�jI6B�I��Hh3��ӏl�z�2 ����C�-RZ�c�@�n|��J���C�I;W�P1�E�ϥW�b�[KԤNƨC�	'V��pA%��>j�P���b�l�Or�=�}Jf��?Fp�� L�����KDA�<qa� �(�_�!h�]ZC�DX�<yq攋}BS��٪ir�{��	@�<�u/Z�b̹0��g	b$�P�T�<��սD�E�&�&u����`8T���g{y�I*D��>G8�"�,D���1�ֿ�,a�E]�`-0A��5D��qaNW�7�.P�BbF2m��(S�4D��+�*[&iDV���+��� �.D�$c�M�5��%��"�8�¸�tF.D�dS��� x0)&��e֜p�h*D��V+�=$ ���_�^��c��'D���'��0�<qA���:B깲`�%D�\Y���C��-x��#aXq�	}���O� ��a޶	�0J=H8�Q"O���Ti��B�4�f) �0��I�A"ONA�e�-y�Y��ӞG�f���"O~�悒2.�]�f+]!��Ev�<�0k�Q�h�+s�z	K�m�<񧀆,2/�Q��mM�]Ul�Z�c�R�<�G"^J|�F&N�2=��ǒRx��'fTq�I*S̬�;���*s�x�,O�=E�D�ެ���`)
9;���F*��y���$	 ���KV|�E�	)�yroT J�D���^�I�)c�H���y`H�fs�(�ET�GXvmBd�B��y2�G��x@��(G��t���yB�<Ҏ	A僒>US��:���=�yb�˛n��y��Dw �I1��I�hO����оL-�Iز�U	5�9�o��q!��К0�x��A7�&q�7�B6>i!�dA7z�|�笖$��1��O�	�!�R3EL�8gצLaĈ��H� Q�!���+$K����!LY��ْ4E�4�!�d�&X ��5��>�ʽ��� ����A�'��R�N��xx(�0��)z.P8b`"Obؒ�_�E����	�B��z�"O�Y̊�#u��)Ԉ4r�M�6"O����D1c˖mTBJ�i�4�"Ol�)�	.H*�qG��xN4�1#"O@�psd��4���ꀏ?�Ʃ�"O%�@��-3��8jS�E:$�&����2�S���B�L�)���}�>�J#���=!�d�����+�dW'pvN�Sa^w!�DP B8��Q���Z,i���=I!�d@�h��Ip$�KOzR�+~ !�$Z�e.\�0�PZY�Q�7*!�DH�{���G�x \��X�'!�A&����#v^ଐq�� !���_����Q5mtD����	=�'Ua|�b�?e�@�WI���\�2��-�y�j	�)�nl��'�H�jf�گ�y���~ ����b6ų  X�y�hܵ �0KB����ۇ��y��L��R�Z�.�I^^�9'͛��yҥ<E�Ȉ�ĉ<Vvd����<��'�ў�O��̺p��[����D�׫Z�dU��'D��炄�[�� ̶Y��S�'�T���B�{�<��Q�۬W1`���'ĸ�1��A>}��i�	�
=�Vx��'�|}{����@)����-JT�x�'��E"�0�& ��/�-D�H�'�"d���TQ<�����-���0�'p�RI_<f+��6ʼ��ay�'B(�٠$	)Y���Y�Ǖ)Kh�y2�W�gE��ђ�IQ��+��y�%�j4B�j��]�SrP+�+��y�%�\��X���TQ~Z8�v�%�y�lS@����d��s�ҡ�����y�[�%qޱÕ�Ԑ5�`"f��y��U��2	��{zla�r◻��=�$3�S��݇0����Y#Y���WC�o�<Y�2z�,����
�< �u�<��υ
����T���a�'��t�<�6k���|j�'��Q��5�ƏPl�<)��p���OP6٢%� i�@�<y��
.�H�ǁ�9h���Λ��8D{��	�x�ҝA%kP�`/Z���Ɇ�V��C�)� ��񤫖�+M����F�A� ��"Otu���Y�&�48��)��b"O`L���і%�����"�!as"O ��7#ܩc�lĺ�C[�i2���"O~Q��
���f�6��i��=	a"Odx(7o"CH�����e��ѣ�"O�����2
����7��:��Q)�"O2� ���$���9�#��C_�#F"OȤ�t���Z>,U�h�R���#�"O���Qㆠ3:��G�)	n�4"O��a�ܕU��-Iq �!/ ����"O�����h=�� �8� �T"O`�� ��:n�p�f�[�#T��*q"O������9��|�c�H3Q�u��"O8�pV�H��|f�C;�E�"Of칑�ٚ��)���r.p�Z4"Oв��T����͈-4M�*�"O\��2:2�^�[6�*#Zi;W"Op��@R5Ȕ#����:�x�"O�i����m�x}u��i	���T��G{��	�J ��QH��N ���2!��#^��ۥ�פ4����S-B�">!��U=ˮ\�"oHyͺ��ҭ¸p+!���8�~9yd�_�M��Ku�M!�D���R���ְW2pSg��!�L;
�֔p��B���<I!�dʃ.���I�%�
d	�o̽xGў���ӷu�0�0���RFy
�ɞ#{�DC䉥v���I�i�j�2��%eX��&C��H��m���Fb��s�*�M��C�	,G�r� ⪜�}���qlU�>U�C䉊DRpT2��X Lt��Q�V�MkNC�	&z���7M�Qt�dP' �
WlC�I�!���6,Q�>j�@8b� 8$B�ɷ�.����ð�*���O6�6�OT���] H�AĨ��4��< c�*j!�DVqq��I�XW�rT#��{!�dƌt���@�B; �q'�4B!�dH�D>����	Z5�)3�B�(p�!�DUJ���bvJ2x���]�n}!��F%�iXs�m�Xh��(�"Zu!�D�lij�q$�g���{����*�!�_��v�#�r�+"@�!�$�14���Z7�[=(���*��lj!򄃌=(L=T���B��A./]Z!��	1�I�ЪXo�����&R!�D�Z�	����W�"3!�M� E�Æ�:$������c�!�D�j��J�46|�̗�$q�O���$3B���%&C#%�`z�-�<0c!�d����	W��E��^�P<��@�8��h�����z�$�X��фȓo�0	Z�ʇ�7%�  �j��:Y���MZ��$��޹Ӂ�͐I�^���<�����N
�$��6(Y�rH���O��2F(Z:�N8��U�v�j8 �'����_<4)�H+8e(�'qLP�%��$�5�n�%@Ȟ�
�'� "��pTî�$2��z�'ܚ;ɕ�2w������-��P�'���	 ���y� ˛)�H��'��M�W��PCp�2MB�7ʤ4��'P����NK��l�Հ�+{gDQb�'�K�\$��a�(��#�(	�E �{�<� X�[TB=8�`9��ހg�&��"OZ��ƣ��y9AR�\�F40�"O�����)V��-�4�ݨZ��M��"O.��I4Cpݙcd�P�� ��"O�����^�&��rt��4V�T� q"O�M�$j�_u�=H�RD�����'�!���K�\Q�#B�=
�y��(�F�!��^���FP3~�t��1G[�x!�[�4M�� �Q5p�*��LV+�!�(Mr�,s��H�(d�b�
�J�!�]2]����#@S3� ܐ�h��6!��5Y3�@�eA��"rFLI��_�a!��6%��x e�K�pa&�k���i&!���A�����,5�T)ɲ)͓�!��k�D:p�I� �$L�gi�v�!�C�I.��r[u�t)�@��u&!�d��q$�j�j�R��@%�ʟi!�Q'���Ĩ 	$�ز'*��d!�dȮ�a;�E&��<3��X�E�!�9L���3!��T�Z�
��E!�$_+��U���J<��A�V�A	n�!�30�a�	�L�:��v�
On!�J�^�􄠥`S,�Ճ��ւ�!��;I~)(���%uh��wgN>�!򤕫^�0Es���L9.���E�:�ў��I�)pF ���%m�Px���!^��C�������	"�>���%C���O���
T#l�P0��8l,��F�ad!��(3e+���Zn䱅�Q�TN!��V9�(x�5�Ї?�M�CWD!�d�)Sn���Âr�遐M�,4!��/���'h� �܈6k=A�s�	N>ł�hG�O�A��U S ��3D��ӇJ��@�=�Ǚ`� *�"�O
�=E�$�Q|��j7� R��Ã)͸e�!��D�@3�-ÀFKxdʆK��!�ߕg���g��)O$#ꀚ-�!�d�'S\�!R��5v6�4(�1?r!��èRV���F #��wHĊWD��F��|ztÝ
d]*�jSAC:M�!0�+D��q`�J��D=tH_�g4n��3�%D�|�I��KJ��������S�9D���#�]���AaG�,��� �8D�L+ E  "�y@7B] c�ظ#� D�<��Ô
a���	C�����>D�P0��êo��l2U�V��8KC;<O*"<�V���?��5�# .4fT(�Vu�<9��>Hk"����ϩN\$P�c�o�<�FB�xy�*�#[��4��Vi�<��R	DA��!4/)O���Kej�^�<�D��B4HD�
D���$�Tp�<I�`U�d}t��m� ��1��Mh�<і�K�k�,u�£��^�u�' �f�<���-Ks�	�^$[J]څ*�d�<�r�1�t#��W�@I2���^�<�`b9}�`C.L]&<�H$`P[�<�`3Ӑ�Q��T�M{*�	҅�^�<���ÓE����	$��1
X�<���/7��	ad�mE�<q��Y�<9�m![\��b��(��)��@�<#M�M�x��D/�/5�@�H�{�<��۠a��[d��<U�e��R�<9rl�m�ε�!Ѕ�x���K�<�b��P{<�E�B��P�&�r�<� �L�틶}H�"����:l�#"O�]�+�&ݫ�EG�׎��"OFhs-4������R�P��R�"O�@�ÀA�xޙ�S���d����4"O шT&־�:`xr��~lv�(�"OL1
�cG?c`5ia��":�R���"OH�ׯJ&6�\|�T�L�@�0�W"O�����f�@�
3jؔ~����"O.U�`%��z���#*G�/�؍�&"O����Xa�J�Ǝ�E蹢TV��D{�ɔQ��$���L�3�HB�=�B䉥yd5+B�J4c}��d��:�<B�	7��zB��Ij��yDi��XK
B�Tm��а!E�P��S��:sC�ɞf;�
�T�k$� ���~�B�IW&p���60c>x(�C�&�B��:�v���X�z:d��-��84��D-�9�`!�>Պ0��;��U���;D�`��F�Y�0����5:V ���8D�4J%"����]��JR8!"�ba6D�L���y����3Fb��c5D�,��(�	~�.��C(�8��q�=D�af]*S� �s�E]Iw��;D�PH��z�������$������O�=E�D��e�8� �n�/(��]˃m��~!��Q�myd�&��%l�X�ӫ!+�!�DLgIt���KXXj�h�D�D>!�"Z�8`d�!s`"�H���'�!򤃭 ��q����G�L۔�Y�O�!�d�5M���� 2�86���N8�B�	�y���Yq˗Y�8-�sk�"^ƒO��=�}FI$w&��򦀠e[��(��U�<A Ό�!<�pw�M"^"��ReR�<��%�[Y�Ts@��($��u�K�<A��&L`9
"M�����ME�<QsZ!M0�耏�)�2�)��y�<i�(]�x�A���'�h!$�y�<�C)ҀAh2%:Ҥ��Mh��u�<�Ye����'_�\�J�E��)@�!�Ă��A�!NG�1����Oߠ p!�	�`��Gը:�P�yaB8Hx!��T ���`e��3�x��B]q!�DZ@�fDᄠ�1�`b�bh!�$Y�s6�T+ƀR�C��YuYGP!���?�ЈR�Q,^]��*3`!��T$��рK"k��}��Ǖ�eK!�Ę��@�sM�.��"%�4�!���/'D@�k�D)B���Q�}3!�-���Ps�Whp`��[!��-'�8=p���=z�hP&$1!�E�M��T�Ɵ�F0���"��6	�!�d�=Ů}�%g� .Z�5Aٔut�	N���B!��:�̐�V;D�H��
!D��ȱ�?X�D�U���s�tKB&3D��z����}q�ɪTe�+\'`��L/D�,�0 �&j��`S�A�rGnt�� 2D�� H�B�ęq l�NP!��<D�X�ӊWw�����
9o�v��%+-D�@��o�[Ԣ��w��L:���'D��!6�8�� �a��ޅX�@B��k�ޠxf��<7�zqk@���PMdB��?���e��(~)Q��M&��B�	�p/X�� 7�NspeI?C�	�fn��4���]o 9�1��U3�B�)� ��X�ʚ�@$���(��ި�B"O(E�dc���:-��{8�u��|��'�p\�v��B��"7��i	�'\�0�L�\�@L�%�"Q�����'G^�:1��DM(Q{���FnΥ;�'B�[���o$YҶ�=�x��'�
���:��%;�#�0d޾!k�'٢�xCɕS�"��v��9`.���	�'�����Nc����v��;.���x�'|��+g��yg��A\@a��'�)�AO9z�
�:���J}x��
�'dم`��jY)�J�E�L�s
�'�R`�c�B�(&�]��&q�	�'� Y��T�.ܹ������'=z� �-:BHi9F�ݧL��]��'����/��F�BE�B.K:�l��'nx��$��x��$Z�	�(I�J���'�@ه��<"����0nV�n^4���'
f	�5�R?=Q� AE�Q2�'6�i��o!}�|*����+
�'��� aL8/�vL�n|�6��
�'۶(�#��u���g�'���'��{�M	�}�n��K(:x���'�`�bዉo�̌�&	��i�.���'�|��( ���Z��{�D���"O�(�_(xfO:	�T��K�0[}!��<�"th#����i�4��!�$�'���劄6�����/DGH!�D͋l)�Z�K�3CΉ0e>!�ĝ;0�2 �q�k(,�I�-�,lU!�D|$����CZ�P��a-D�E!�$	�\ �Aa���Ѓǎ4&A!��>[��l�1��%�&��p�.0=!�+d?L4	�/��z���?~E!����bt�UlV�.��q�Ƃ���Pyr�3L6���7���Ls��pm@5�yBK��*n68r��:H�`��tnP���O�"~��T�x�Դ����O�x�!FW�<I���4|�|@3N@4��T���k�<��C�w�uZR�H L�Rt�s`o�<��n�_���� "Z�Ȱ��k�<��I@7'�
	*���WT`pS.Ne�<��eޓa�����>Xi��[d�K�<�&��+�{�)�0�R,9�ƂH��0=р"�-w���kĠ8����J�<��e]�`'xI�����Z�C�B]�<�BC Z�Dp����c�� �`��W�<it셷o_(<['I��&(�x�I�P�<C"��Y�����I=3���J�P�<ye���cR2�)r�f��	Tc�Z!�ď�,jh���B �L���"��rW��DƔ?�Ra�A�"y0-��G�_#|B�I/c6�0�oW:	��Z�"؆XvHB�ɬ9}�P)f�� ��8�E��i�TB�1O���.	��P��jE.Ecw"O��:��J<�Q$�3�6� �"OI�Ǉ�@5�1���O8`Y0qZT"O��q��1
��ț�j.	�L���*LO�i�SK�`�%JԼ(�>��7"O
��FCҐBT$`�����)!3"O�}�MI( �����g����"O�8#���T"��@��zk�"O��w�
*BL	"פp�t$�a"ORTj2"7��:���)���p�"O� �U���CD��#��d��9c�'w���V6vpI�ӣVy�T35D��!��0Kzu1"n�4a&�d)7�1D��f	(>��L���m�A�R���y��Êj��[5��X6�25��y�
�Evc���*Wd�q�.� �y�ɑ� ƙ�����  ��'��>�y�i�S$7˒"J,"�Ss`@�!�Ă.#���f璥Y�z �@�K�Y�!��4j���c ���|`����$��!�F�pE�AxQh����b%*G!�0.�!��*1챀"!�!�!�d�+n�T�W.Q8Zc��CC*�!��D�^l��G<1��EF�0]�!��H��ҥ�)bJ(t9��H�!�=+_�IHE���$�0r�m��!򄟸6֜so��Wk�})��-(!�DK�:L� ֫�#
�I1�K!"!�$?h2�: I�`�s�蘼�!�_�c�aaD`�'\~�2'@�*�!�%!�ִ�7���u���S(.!�$�#HΦ�1rK<�n-�@HO)!�$�;IX��`f�����qU��Lm!�¥	��u"����-�� �V�vS!��O0\�.�a`�:gs(i�#
ʟT]!��'LT��%�B�CT��ZpJV�{!򤗲^ ���t)�l;|�H5/�m�!��O�C�v8(4��f���9cJ9H�!�$��2����&ߵ*�f�i�LT�
�!�/Y>tG�+��!��.;�!��\061j$�ҔV�$\YG�Y�}�!���w�,�K �Q
i�P�3t�� t{!���&��Q���@�	~t�¡�)r!�їB]n�!B�;m�(���LLC!�D��n��Qr#��H�b�a̮�!�䟽T!z�s��9����!��N���$�:]�P��EC�Fzơy�G��y2"�4 ��x:bD�>ꀡДƓ��y��y<ȕ� � ܺ�h�7�y���J�س����3�^��yb��vu���tCR��`c���yBF�9k�} �kL�	Q��y��_�c��7Ɠ�gx�E�gIޅ�y�BU<uH�R��A!w�8�xoO��y�/��F�.��eɆs�E�Z��y�M�%8��+��� q��t#�)���y"�C.[2`<`0�DiƖ-RT��y�� H�8�P!�Iw��,h���y�N�Μ��$KѲp��&�y��0Y�d���,)����ޜ�yRe΄t"��f-���4R�y� a��9��҆�����yb�ݶ0��%C��÷9���k��ݩ�y"aL�X���D��0)L,#ֈՌ�yR����9�U(ۓ&�z �_��y��1L &���f��2L)�l���yRȂ
pd�����J-���K����O`#~�`�D(��\�-�VA�q*����0���t��:kD��V�B� 4�ȓ
 �ԋĆ�:Y�XԯC0m���C���i0���0\���B�"n8�I���
�p�FL�a+�ܫwO܈3���ȓ��Uy$�*GE�Pʢ� <$ �ȓR��$J��aN�@ڴ�4$$��S�? ��Yg�ғK�U��j+.��y�"Obb���* �ݫ��&|��"O����g���ȹs�E�����"OdQg�ԷY9�S1��k�����"ON3D��h^Q8��XѲ�"OƤ��b^vu���Ԩ�?>(��q4"O�Yv�֙��1�^�R<�hR"O~�S�O>G���Ғ�]9Ү��"O$��I �.�W��`�&��F"O�a0���YoA��C"��"O�8H�3%��A�-� +ti{�"O� uI�6/ �	���>-	�L B"Ob�ȧ�]xZB��U�.�S�"O���B���~�ƪ�+NF�{�"OL�d�0l"�D� ��5q���["O���	�Zu��!��8��b"O,Q�H!U�:əQ%��9�tt�"OHH�y���g�\~*��g"O�E)�-�� ǂۂ`_�7xp5`�"O�р*ֹA�.�xdO�=� ��d"O|$�se���%s��#K����4"O�t�PBA�t��rge$w� %G�Io���&JPK��I톛0Z��j��6D���S����0l"�,��l3D���d��rȬTs�&p�ȹ�'�1D��W��O���ϙ6��K��-D��%�N�sp�&�/
x�T�/D��ٲ��]$�-�F睞Lv�C��'��O��S�]vb`�Ɉ�s���X�D�^6���0?�!+7�. �*�@m���$�l�<��ʉ�9?�9�D�!-�\�C�E[R�<)%n�i9����)Ƞz;�D��O�<�b���� D�&+���IlMJ�<�* 	~~�@�Kؔ$�n����D�<�S��L�JI:�O	5�����C�<	rɝ�'j^(�0�����V,�T�<����#Ҹ�ҁ▰ Ű�£��i�<���;b�ň�� �5`�Am�<	��ֶ5�bl1���>RDڥ���S_�<�7�4<,L�:O�j��A�<��e޲t�0��g�՟lQ�(B�Q�<�Gn�-�*��K�U�Ft(���K�<Y��'~��}SQ-Y	I��@���l�<� �<���� M|��X�
d�<YE��L��c��Z֍�#�c�<�d,����&#Q�?�`�A��H�<��ɇ�,���N��.��`A� B�<��g�L��ك��/{tZ1�b�Xg�<�r�X�LO����`�)I�~�B`�<)3o��0S&'R�h���4FM֟<F{��	��M�>]��儚+�`�k�⁻lnB�	29o�)�f�
/��X�e^�f�B�ɘd��P`"��$�n��(�ec�C��R��p�Y�3"0t�"P:��C�	�0���#G��6A�Y��IκB�hC��/��y'jJ�P/8�(̸C�TC�I0r�����fܗ@� 9���S�l�$:��jc�
/|Z�ۇ��ظë!D�tR`�ۤy�Y��͑)E� �T�?D�9�e��'4�TS�0v;v����:D��
R'��H4r�
0�h�zs"8D��Fx04�t����.�`C�	Ihu��nǚu-�MBr�םb��C�ɄQ���`��8��\��(ʢkZ�C�)� ��q'*K������df�v���"O�]���{.�����)l��|p	�'b�e�����P"j�3����MZ���'�	#u/�yezD�B�<���'�j��N=|Luk��	� ���'�R!�ěBbdxCƍ"��!�'�hC0oJ,NXv���.#9P �
�'�ލ0�*D`xNh�b@A8�`�'��ڱ/�;=� ;�)�d���'h���oLC�쀐)%6���'<1灼;vfp��b�� �����'U�Q���8�9�@�$>���'uҭAЭH�F���2ä��?�rp��R�'�B����4IL�4�3���(���-O�q3F�R+�xe�_n9`�"O���h]6*���Z&&�BI��"O2 ��GǙL�����*�x6"O�4y5EB\0lk�`0c���"O0ScgP�H�%A�^
)U"O���f�^�����9"d"��"Oh����ԓB�� �Њ{�v���"O�0����v�^r�� �*(!���7v�$	3)f8|!81��5-	!򤃿'8�d�ΐP0�ɖ�R�i�!�11���8d�ޭv0f@�Ō���!��Eg�R���f��c?���qe�R_!��A�-�*�+��T�!�E�S@;!�ϵ����)Y����QbD��I1!��sņ�(P(+,
%��#T;B!�5}�F�q(�w��(�PV�!��I�:�;S�[�~al��b5b�!�$��<X���D�k`z=�w@�'t!��D;N3��y0i@fV�rE�R�t�!�d�G9z��@`^���Wǟ(�!��\8��)���\�ЕŚv�!�\#g���R6�
l�d����:�!�	��(�ʂ/4PȤe�PǀBw!�D���^�	o������!򄜍M�2]�#����L�0�%_�!�^�0
�m�Ã��q��a�U��6p!��b����0(@�M�>�{7��}���9OZ�9��o��Ԣ���4L���"O�1�|�xf�e9j�@"O�\*�i���xp��cū$�xS�"O�� F�>7b��CǸS����"O\�xv-�fi,H�ȇ�,��qؔ"O�@#���:�L;A������"O:Ԁr�B�6�@@'��0B��t�"O*IYvf	�`��)FA�jP
 "O�h ���\���с��6 ���0�"O� x� l8UA���c��-j�"O4XDl�A{�Q`&Ke�:�"Od�L� Z���#��s�ۦ"O (c��	[ۢ5`�M�LF��b�"OTuSpo��h��E;dK[�<��"OԨj'g�*
qN����6�$\[a"O~x؇�	�R��y�@�v"O�!6&ܥ���u�\3����"O���T�I��M9����"O��C�6/n�ģ�,�#t��ae"OvP��? ��h(���>!+6���"O�kr�+���(�B�'@G ��"Or�[�a$�tcT���>��3�"O�@T'�FcRMr��ד[�: �"O� �4�!���eK���!�*��8�"O$LYqk+7T�w+Y�8L���"O=���!<0&m�'F��"O���1�E������ŷJ(PD��"O�	���p���A�
�S��q�"O $YE�L
��04�R��ެa`"O���Ռ��L��x��ܚw�4�"O5�B�=0
�!E玷m��;�"O���$��	��@�B��s"O\,��,K�'�5�I�0J��ݙ"O`d�Q�Њ#������/N�n��`"O���c�30�0��Gb���"O
�@Fd�u��Z.D�)E��7"OP���:d�$[�4Ԝ�`d"O����5X"�\ڵ���.Ѱ�2g"On�2į!%�9�����hx7"O��,�$+��Ȕ&�zS�"O���k�Ր�rD�NA���"O~���o�JD� c% �q�"O��2��/��Tk��\+�r)r"Ob���#UG\�/��x�"O��Go�$J�@Wh����"O!�V�V�u:6Hq���7����NK�<��ˁ�����ƙ'�4�apa�H�<i��J oPlڃ��>�0�eC�K�<)�Cn��}�!B���<�Z�-OH�<i�E�
�@U*t�QY�i@�N��y"�@��^�Z��k�,�c���yB ןq���U��z��}pC����yR�o�����fM�@����G$��yr
K7!�8��`OB�6�&Ĺr���y"�^�9C�i��C_�-�<�"�DP�y���.+^���B� �섛 �8�y`�G'"��&�#W����t��}�ȓ'YyrR��3<��{�"č'}>܄�}�����c˰re�� �@�#A���G��ۀڋA�	�兗,W�h�ȓL�r�(2�'�,��.�.+M����.˔h+f�%c�Ƞ�q.�?�>}�ȓ��0��`�Qb�а@ F?+��4��Ғy�c〓]�P��� ������ȓ� ;�LDc�Mp�J9FȮ��ȓF��Q��<+|r����4Q��P��75�D �̓�2W�S� �	U�<��\�y�	
E�d�97�B������\���EW�-���
��N�fą�Oc����)P����3ʤ>6b	�ȓ5����5Z 
D���/&����\�s��Ug�H�m��/��Ąȓ���Q7��� ��t/ΔZ�Ԅ�{��Q/N3�"�x��
>1��J��x[� &"Z1�iʏ~z:h�ȓo�j���- �5`ׄ�	}�ȓ'�Xr�Dj��;r�ٔ,��A��i%\�t����bqΈ7|����f�3��*{�f�!Q$2�����w�S��;J$a*wL�~��D��`��A�١'� ���\?�ڼ�ȓ��g�*>V}��	.����q�p�w���'
�a��q:D�D�D�ɩ�����1�9@E#D���#(�"/�4�9cV�}F1�p$&D��Pg�Ǎv����S�S75=ڌ��(D�<���_)}|p�p�\=(�a�9D�� |��E$�\~m��@73��HD"O�=�46�ơA�/ըi�~��"OHE��I��R�n��¤S7]��W"O��X n6Hk���:R�BYc3"O��$a����A� �W� `Z"O�����S���AcB �3�"O�$"�ˍ�� ɍ�j��t#t"Ovd��g�5E����
 V��PY"O����B[�*�0Y��D�K� (�"O��+M�w3�taE���
!Ó"Oz Ȑ@۫|� 1�����=ِ"OLhPTE��\�
=�� �:#�|@A"O���-Y	^�� ��\��`b%"O�5 ��Q�(���3fE�����"O���D/y���fA�A��Ma�"O�)�%K�(�p��B�"Op���*]�_ih��eb�3��8)�"O^;��ÒA�\XsK�*+��8��"O��pr�C@�}� �-،�Q"Oi�_�j�T�CY(	ʞ�@�"O.mk��C�-{���	O�ڴ!�"O�y���1Dk���(��V���q"O:�3��T��4��'Gq<3�"Op@ɠj4!Ӑ��GHY	|>�<��"O�i��j��������#Tݮ�"g*O���`ʂ���c������T)�'� �K���?pԜ+�E 8i����'\@'���E ����GE;h�P��'���D�̍X�b-�AF���(�'XPbWe��Nj���ₙm��h�'���!�E�,BC�10��/c���Y�'A�jr�K$uڤ���ÝWl� �'.��(�m
�1��rg�Xb�B��'�.ґk0N�	[Ġ��a�\��'Wp�y��6x�"��B��&6P�
�'&z��$��8eg���I�,����'R�`�Ί!�����K��|����'_(S��[� ����J�]�z@y�'�xa24�"|6X��[�[��H�'X��s�HG�!�t�Br'�IL���'��Ey�f�k���!�M��(S	�'L�]�4���Vz���D����'����?Wg�*"��;UR��'+\�я�_"@�Ɂf��7͒�i�'Z�܂"gX�$*=B�'�5^]�J	�'?�yX���J/�ܑתӘP�|�Z�'Ğ}�e�U�\9�P	7^A܄p2�'�d"��37L):��_2D�:T��'������MW0�	@�ȗ2T`Y�'	�``��V��
m��%�TTXY��'=U[����`D��Ms�r!���V�I�������6�Ȯ<�!��;S��H�"�J$I��@��� �!��Ǿ9v���h�ot�bt�Ѩ>�!�d;3�3!�M�7�h�%D�>(�!�d�#e"���B�A'g�H�`�Aw�!����I��=C�l�`V�U�6a!�+@���� �\܀�0h��8a!�J�-Aba6Ȋ}�T&Ñc�!��PA赑B�W%���EHR	:t!�$��yYh�[��O�k��qa�[�V!�$� �*@�C�J�9V�
(l!�Dބ��1�mLYE4-���Y�N!�DP5S� �")�}�d��6!�� �I�"Y5]@����)̱��"O�tS��L>@�����7z��0c"O8p����/|��d�h�=�~�b�"O�h�v�\�dv�U�'�1��F"O�ء7�Ӯ=R��3��d�6"O����0 2%�C#@�'c6���"O(	)V��8���Q��/@����w"O��EOV�S2Zݨ��C:F�P٩0"OrEK"U�#�!�rm�0�@���"OԐӥhL�.>pr��,S̸I�"O������i���V���f�P1S"Op��C��+U����4m&T���"Ojѣ7Dζ�`���KO�9D�y"O����ß%0��r�d?s3@qt"O��)��k���2�=a�\K3"O���!A5!���	ƞ�#q"O�XY���[���S�mW�:�:p"O�=��BpJ8P���& @�"O6��ra˃�H�ǟBk`"OX�p5���>�T����C����"O��	�/��nBI��)66� w"O d��˔8t� �b�F�8����p"O@D"���7p��ūA��>a�6"Od��3h[�iA`h�Ӻ�4y�W"O���S�>V\��`R�fX P"Oh\�F��U���v�"~=~��w"O���P�յ5�:���>`%,)�"O�`��.��|�f�3�ܽ�R�3p"Od̛t� �b]�U�6<.m[`"OH��%Ϟj��#�I�]*X��r"O25P�&@����jEH 2"O4�Y�%�>�,h�"[c�DC�"OP�L�H��r� ��Y��"Oz����2#`p��֦Fe��J�"O~`pF98��Ї��j@��"O� @IA�m���e���Y{JX��"Od(�5L+��YU�O�'_&Г$"O �x&���|�k3c�:A��YD"OXͨ�Ϸ���)aT�%0#"OԥAc�G�E�r����}�:���p>yO<��c�7>|r��r�27\�`����t�<��!��^�z-��ҭ+HA�"�s��+P��<���9pHk�  �Ҡm=���Ng�<�Ҏ�&d��B��0�`1�bNW�<Ɇo�EB�ҡ�IW\Q�<iu@ �oʮh�qʙx/�(:S$�N�<�tM�	�H%���242����B�<I�KR�=����d�P�X��<�JA�<9p�.�%c���Ȕb�ŝ�U2�C�	����j��BR_��ۧonvB�	"9�AjE+\�  {����'�B�	�E6�C����F��mܲ%�6C�	'5[��ˀ�߂'�l�p5~�w��!|O���,�S�
%.M�**�0PE�'ݰ�l0�t1�q��Dz�����,B��-12����#PA���㴅8V����D4ړ1i���ӥ�Mzn�"W��lÊ܆ȓ"y~�9��^0Bi�?Dl|��u^T�B-��y����#+�9l	Lm��t8, �1��$8�9z���7`�Ԇ�}���e�O� xٱ��5,��%��%�@�j�h]�OPy��Aa���ȓ'��y�hY�x;@9 �iH⼄�S<���a�G�`:掞*����S�? |i��*'�z���M�$�04ٴ�i���.�)��}⤯�	4�:�A�I��r��h�8D� ��7��]Z"�^��F7D��
@�/유���џA��YQ£3D��*�"U

ZH�L��#��1?D�H�G$5�Є(� �2iǌ��g)D�\p���'MZ�@�L�m�r��:D��(G�ٙ:lXp���#0�h@�.D�p醉����A�m���\9��*D����U�=gČ�櫓0/����5D�󪂂n��9���B*D (��3�O��D�:��CS�k�H�e#��j@tȄ�RU
ݚ���2a���1�K\�z�Ȅ�6���0
ft���w�Du��Q��Ih?�(^�6�{�H�WβX�����'��I3�H��Ic���#��?<� �O#�zB�	�:jPM1r"�P�����b D�48�?iӓ\����Q�C�D�<����p
\��	B�'��]���/&��mʷ��<�Ǹ�yr'X�C�`I@�)o�’�I�yB��e���"��&7��<�DOI�y�H�>L��� ��:${������?�y��2\�Da��/��@�z��5�y2����]A���7�6��5����y�K�>l'Q�U�����t�E��yb��8c
����1�4($�؄�y�ĉ@��@���I��Hã�	���'#ў����{�Ç%��  �ư-T�p��"Ox��s(�2a���Ri\;Dq~���i�D������ēp���舣~����/�2|���ē[��D�T���A"�Q�R�
�ѳ�$#|O��� �,\�`6D����p��O���@[~
,y@��=⩛��6D���$��7�Ƹ�����{[�,1e"'D�@�����/f0���x��А��%D����P/H}�s��}���Ԥ"�`���OD�XP��\2:�	
�bU�-��a��'��ECP!�"N>hHk�k�8T&&����D+<O��(�#7?�ة������E��O���1�MyȨ��lԶ$ɤ�����]�<����."xu��F�5����ЩZ�<��a80����@]).�"1y�i�U�<�W���m:���'~I����T�<��E+^C,�b�%N�{	^��-j�<Q����@��Z��ވd���l)E�!��E���a�%�[� �)c�]�2+a~2Z������j����ɛ�FO� �&>D��b��?(�2�¶�Z�V5��b�g<�	�<I�}J~�gu|M�",q���&��t�<�`'�$όMQ��`,�`("LR�����y�^���ƻ4%l����P;���	L�-0GĄ�Nޞ`�ِ~���ȓ4�Ɖ� ��<I��[0�
�j����ȓ3��`�+ߙ|T"hq㬅%2B:<��BZ�1��iK�|�d� ��|��	l�	�-�@@p,��K�\]��-"�C�I)�ȱ�/0^G�HP�=���<����*牝'T9p�F�#7�b����C�ɭW=fiq���8�X;c�8;�2"?9��S-||�!�5�'B��H�Y�pC�Iߦ����j�(�����Nh�Q7
�<����	Q����$صU��U �a�4M���9ғ!�fEK6�T;�$|�O��s����ȓ��=�VD���Qk���6���I��O� �$�E��/��p�.ݱ6�ś��'��M~b!Fw44�
c�5|R�l{�e	��IVX��0"�8w y��/�<��y$ړ�ȟT��d ۓ�X���!�1d���a�C�<����Dj��r��/D̈ek�XX�\�'��	�n���Pe�Z���q�����B�	�O�d`��/\r��h�wd�0l�*��D7�T?8 �t�t�K`��$������/D�p��EQ��XI���A"��Y��$�O�c����Y��S��؋x0R�t��I��*D��ztC��nu���l�5�!�'�,D���R)��P��p�B��K�NY�t 8|O�b��C� ��w9��@��	�%�IS� D�p�Q
�4t��k3mǤ!�"Y�R�;��Ʀ9��%=�)�S4������8{]P��FєW�^B�I�^*�i� �:��M�7���u4������O>�w�  �&%��;2l2�Ň�5Y�"m��z�����D�D������d6LO���@��}a� B7l�2_�$���'Xў"~B�-�=Q��|zP�`�d�K��'�y�
eB|��!Qz�{D%	�䓯hOq�|9#Y�X�4�tP��" �a~�T�����e��!vV���4D�h	QK��$e�u��=Q$)%3}xR�ǟ�(���c+|	P�U"o�]��,0D�d3AIŦW���G�rN�ف�!D��rmT�rWp� U�L�=������ D�p�6��hD.���/́Y����f:D����Y�}"�X�k�(�"ȣg�%D�\
�
��.�F���/FGеh& %D� �0d��r7E�z�t�%D���%E
�y�0)@�遾/L`eP2 D� p�Ƒ�ZT�\AQd�&�I&�?D���"����L1{�k�f?D���'ߠ���D����%��y�!�D���8����"U��rET�!��̹)�`]��l�;���C�a�!�ē�t���Uj��G���*��ZS!�$�-�����/Y5��4��P3<!�D^̩q�J�#xD��Ϲ$6!��S��E��-�5e��@_=S/!򄚍E��i �N<<�
�jՏ�G!��A�}�(j�T�~n�Y�$��!��-�
ʵ�N�p�<M�Uȗ3!�|m�l��/N� �y�a 1!�j�h��	4;԰("�K�!��4��8�J�'9�Z �cnӣL�!��76"с�
��^�$�p���Y�!�Ē:a	
�S!!s�X���L�\�!���?/9�+� �%pn���+4u!�%ab~��&�T6:d*]AԎ®#�!��:M��S�
�S$��q3FD�!�d�=b��X2d�$�Tc��A�u!�	�@j��:$F�1���Ȇ�ɗ?�!�$ bJQ����:�� [`�^��!�d�B�&��P� ���P4f�-+|!���vڀU2��L9t���e�${!򄌅D���i��֏\	��qt��==�!��!E�^U�eC�`X#m5!�$�*Q�ԥH�oI(�%
G*�3r~!�$\̮��p� 1�D�"w�єy!��=%�N�2`�X�6���J�v1O(��V�� y.�+2���\���$:%qJQ��dɆ-�^�S&�^	~l!򤆃{6�Y؂ƤX ^��� D�]�!�� 8äN۟ i�Vo�'��8��"OZ$HiA8�"���)�y�T\a"O$�*D�D2vq:%����@6j�c�"O6�����%z� v�O�`)����"OL��a�4"z��b�	/p���"O�(Y�"
���`&��D�l�"OȠ�fK�g�E��n�^�^��"OK�{eR!��eX&Xt����5�y�*�N_R<9�oϏ_2^!ɰF �yR�N�~��abS΄�O}����%���y2L�4.�#�NY�;�Zp�h�&�y�c_�^�@JAnT=-�);����y� |`-`R-]�$O�A"�׊�yBB%"jX��C
-���33�8�y�M�)+s�Y�q�,B��e�2l��y⇀ n�*m�m�GM:@��ϝ�y��IF��#7j�:Ef�+�a��y��ۋ�b���Z�!(�eH�B���y2F'pv�}W%�,�%�`	��y2���T�lUl��},z�!��!�D���rt��^eP S�ٔ!�Uq{ؘa�gS�Ig�� ���M!�	0#/2]�n�5Z�^%��a�4!�'C^��2C��e�hŲ��O
!�D�|8�p���˨>�hP��1^@!��<@���8Ș!�N�Ũ�k!��){�D�����+�����Ş<�!�9P0�=qp' ��Z��Y�H9!��		-�\�"�۱����c��6",!򄀳�6#�"� B���L�/!�$�S��r�Gk�LP�!R�U!�$�$=���SĜ���%q���[!�ݒ5�D���6����o��!��6�ZXy0f�c3��8&�V@�!�$�O�6a�g͑�E'�a��#X�!��i��æ̖ ��l��a�!�Ԡ%�P�zpa �>����UƄ.+!�d\���#��6ov͊E�&!�d+dWb��g⑼*X�೰���!���O���	i3�u�b.A!�D^�i)�!"�]3:�3F�'`!�AB�=vR\n��"�D5*�!��D#lے��]�|%��7Β�']!�$��<SB$�BR94�i('*�6Z(!�ب`�
`�V�V|��w*��?!�a��y�`DR��A�#L!�DA/��!	rK,O�t�2��.�!���I;B�q��f��H��V0�!�D7m�N�C�Җa$���4�!��EJ������xS1A�$a!򄚕~�"���N�i�~a��
?n!��9\�l�qq�!}.ČK�hZ%(Y!� �G�D����[�����7!�d�&`���<@I /�q_!�Ҁ��m��Ɏ�K�F��#a�3|�!�D�'d�n1���Xt������R'!��"@���`�k����OڟB7!�D�H%���m#w @�S!5^!�$:,���(E�S)aH��"f�ĨJ!���P������y$�8����F�!�d2l��X�`	�B^ �� .�!�\v��#E�1��QSd荴+�!�dW
k��,��5�tl*�"q�!�D�3kT4�g�W��\��	�gp!�� \��DN��Hvv��r�^�%)���"OJ�{gA<q�q�[���9�"OR��`kԚL��ݐbQ[�@d��"O���%f���݁�Q _d�Q��"O�PYr��-u0�2a.m�qT"O�X�3K���}36"M�\R� i�"O�����F�� ����
Nh1 7�O�<:�F�4�0>��
��z� �*�/ 2;2	���C|����阼.�y��(Ƹbc��0�ĺaGB20�C䉐?��!ÓE[�K
(X��͗ �O H��M����H�v�w��	Ǽ�J�b�<AC��!7"Or�c�I�0/0N‚<b�@�W8r�P �bc��<Yᣆ�6����'�]Ę_����w*K�g�s
�'�*����[�H��"d
Us� -�O{}�	��JO#D�D)7�'�d��W�P�}���')6���Ǔ_V`AW%&���8����M뇎�*'�ͪ�D0490ks�<�V�DOY�"�hZ�w�i���Y� �b�oU,b��Ĩ)�'1Dt�'ܻ|���wf�2q��,"u �P�Xs8��7i�8F�ȓ�"PuB-��'����d��g�I,+p�� ��	xB�|��C�	�:�Q�܋4�)Ѷ�Muκ9ag�2Yލ(�`_n�ܰ��I�9���+�)��B��%KB�H�q������ZQZl��'Q�Q��'�Hxs%!�5������2m�PD�	�'\������,mwJ��@"��"OO���9~aJ$��Z�������v�v�+1���?ӢQ�g&�>(!�ɠC�,�`�KH��P���N���tI���$S�8�p��~&���f�Պk�@E(��Jx�8��l24��"M��p���a�Ԗ�	�D SӠ��pgK¤��7G�~  �	xcX� �G�V��D�:�ŐQmÅ�y��]�7��@�E�$F�j�mW2�y�O�1���[��ت��1Ѹ'sf�#��y儑D�T��	s���4�B�k<��BA8�yr��d]��]g�� �T)��C !v�A���%)�8��4�་�)�72�quBK(5��:��A`�<y �x_FMӅ$�(	��5 5�7�y���7XO��� ��Q2�u{ �[}S^}GxBa)(F\�	�A<H�H�XwG��p=yPϒ-W6½�#��@���	@Wb�K%A�6|���3e� %+�� !4�>U m��?���Q�H<+]D�i%㖹wJ���=�Qk\�&�R����W@�A�bJ��Ʃ{B�E[t���b��,��H�a}"T* D�c�k��6��M��\!N�P�m���Hy3iچ�5򱤎b��	S��7��O���]�uv�C�nM�0�i�P��	ўB�Ir��$�0	M2s�v�p*��jx4`��ϰ
��<;W���
���f��,�I�2r�xc�����աZw��*�I;4��9���;�O�h�f�$PDD�Ȧ���D��RQI_�a�Ԋh����D. ����څر��  �R �1LM�e�ĕG}"��W�=R�+D���(
vN�8|܍���S ?�L������4��*��7��xªU\4���-��rU�I)��ێ�~lLl����ro˫+�nd9u
	,��`�����1h��`��Δ�8�H�ل�4�y��ڄ_�օA�NS�nǐ=�D�P[��u�u�@�<���2O�M�M?m�-8��(���� ��"�䊂�u�a�.V�4;ZLmƵ1f�1�D̫4t	��A%U�plk��FEԠbC!�`x���"�<s��qq�o8Kz�  �@�����=0�)ԈT�����UE�d���n��)tx{�V6���dM4�d0��K@,<ђ.�2��I�}��@82e��h��ٶb���d�Rg��;��p��,�*���n��<q%퇐5�vXp�	�+|�Y��h�R�h$	3lFD����ؔ*�v��|�J>�G�V!ug�%�BUt�yل)[B(<1w+�
PqR2A�"<�䪐`����T%  ��C�
"��ٚU��m��k�8"�NE��ժ"z�x����愈{�[�R���a�&ի{��y�#e		�1�#"ś�L����E�%JEr���'H�'�u�?�0F@^�
�B�D��[0x��ջ%	�,a���Vi���yr��(��i���v!v���`�% 5�"*��Qm����;]��x��L<��&�%t$D���W�4��A���Oh<�� rM�Cf�@�N����>�����W�8g.I!�m8P���퉗&�h��V�*Q,}�b�N�Z�N��dJ\�����V1S\�زa��u�Ub��_6Dkt$�r$~C�I%.21�' 4��tH��&=�㟸�ф�1J;^lBd�@jN�>�C�.�D�G,�)Pn*5aӋ;D��Q�����V
�4U�x�&F����p�X5Q<��R�>E���L�b�J<��"1pi� �"	��y�P"�YS�Qz<N�Վ\��I�8�h�b䫜�6ax���u_�!��ϘGP֐�MC �p?�@`� @z̭ �$ا6z1���E�X�P��G�cL�C�	�{s��g�r9���V�P�@���>�g�A�{9���C,��\��Qu��!	#����ő�.k�C�1[�f�	ڂ�x�E���I�5TZ���Ć
;-�����	�s^�#\��Q�D���9!���J�.����%SC��ˣ�D
E�4��H��cf��w�\�.J��'hTs�Fֿ�̈́�	�S
�,���şQ=��������>1��N�K�V�1�C���(���u�A�!��Y�:����c ���^l�a��� Hp)�F<$xX=�Q�.Y��U�4���c�ȏ)	t�^��yV���ָO�����dV�:T#�n.N�f���'��H��߼L�e��Q'x1�|�-O09{䁂�B����6�Ԉ�j��'�nU����f@�D��jօiP���(��ڥ�_��P�R �\�C� � փ^۪-c�N5�p&'� �ք�enA	;����#9�fw��`0��:^�b>�	��i+ȍ�wÞ/��!:��=D�\B�'�7 ����!)l�˷����y`�]�c�Q	@�>E��I_*m�p���aK���ꗐ�yb�8IJ��"J�j¨N$��I�@�p	�D�I�ax	��+;t�#�LP�%(��p��4Ͱ?���R�R~�y 憧	����q>p�Z�nW�Pxr�G^D���X�u�ԍR��Oqek7��O�����߽* ����ӠD,��9�'R��c��F�(��7 ��aM� ��'�P��B� @��i9�Ċ_ZX��'[֩����i���Hg
�N�=��'6T� o�8��+��FV���'u����@�H5@-���DK�l�
�'00a�����o�ԁk�.��v�	�'�Ę��'�b���`֥d��Q��'H$��3萎4�2	�g�d�$�:	�')H��M_Z�A�C)��������AI�>�@�<:wp$�Q��|�<1'F��mz$�9s��sd�W��t�<��EN:�@=R����R~P���EM�<���V�8Z0�1���~��U	��P�<1�^#oe(Pr4 �+R�1��!�{�<I�j٨]�^ձҩ�F6Ld)�N�z�<�"$Acn�1+���X�D�9R�[t�<3N�9|��ab�O��`iQBXy�<a��F/���� ���Q�@p�<��!ԣ��;u�@��Z,z��l�<�q�JI2`RD"ӓD����k�<�杧G���6A��d1�ree�<�FbҵL>�S	����;��a�<�3��%�|����G8+�zmS Oz�<�2��+ t�3v�W������p�<�1�_K�� h �>~��r�y�<���ڿb�ޥȱF�M�.� dB�N�<GG�fA�	�s�M YP ��l�<�r"��~�ps֪�(����c�Do�<9�G�G��I!�M�����R�}�<��RB�.�c���&7�>���ALy�<9��ƬEV�s`���3�Nh0��I�<�#�ȵ,��6
_�m�AϏG�<1 "����Š���h��|�<� v��ƃ�#Fܘ��͓9�$�A"O⁣Q�@�) l��1�.��e"O��A��`s�)�ad��p�"O�T���\�ٙ�KK���S0"Ox�ʲ�Fp�-�E�ȱ��\P�"Ov�WI��9%@	���R`���"OyrCӥh�^<I��,l�T�a"Odj�o�2ف��f��D  "OB��e�cuZ�1ƀ� ej`�1"O���fꀚRe�Q�� D3;��v"O��
b
��6�^I�C>��E*"O���s+̲%�A�A�Ɋw� љ�"OX�/�.� �)_���	���z�!�D�Z(lȕO5f�4��F/�@�!���v&��Z�铑xV�ݡ1lܤw!�ߚ<~��F%L�=�4ˆ'<C!�d�Y�$=���<+�����)Yk!��5q�h����Ѷ/�B5Ȅ"L�!��h���.=W���% �
[�!�@s8��J#����	� !�d�$4���H���]��R	4x!��JVW��9�i&Y���aaL F�!�$̞P��]�Gi�@M0&*�=�!�	�5��8�d�ɐb�`�q��D�Y�!�d(v'\�:@/B�$���R�J�!��6j��4ӱ
�+o�*����03^!��Z���I=J���+X�:C!�D��04A���/�����@4\!���/%$Ē�mQ-{�ŁW�{m!�)3 i��*/gr�1 ⟊6,!��:L��T��=o�ذ�q��,y!�� o5�=X�IR6 ���2 �Z e!���=u��x����'��t��g�FX!�䞑U-�y�҇�f3��qѐTA!��\)�������(2�|(�'K�yS!�$Q4|��d�T�Y1�|j�\�~H!�dЕgC��	�G.p���4!����ܪ`j�R�0a�+O=/!򄏃�<1 �*G�d$T@���3I�!���S�E�� A0V�'U�^�!�DN.j0�Ycg�e�t����U�!�D��
$R�&�7<>���ݪO�!��F9J:���»Z���A�gT�4�!��"�f!��*'�ҨI�� 4V�!�R*�(s�Q�'��e#䈳0s!�ć�n2dd�7.M�[R�#b�_S!�$�L��'(I
hZ��B!OI!�Dx�bcϧ|�F��E�Ι _!��F�5EjU���r�"�ҧ��"do!�d!H��OW={8�����7nT!�Ė;0��u �&	&^0T��1n��t@!�ʵ2t|��B�>6t�T��� �!��*"�fB�<c��J�͹Q�!�ě�r�N�s�>�E#�`�6�!�<���ۓ�=Pg�К�A�:{!�@�k�& ��90�X���"Z!��K�
]�Ʀ
mr����P��!�d	�8X�J�:(o��c�@�-(�!�dY�o���DA8���Q���!�V:�$c��C:GXA{�%T�3�!�d�\�P1���X9�p�dJ�U�!��q�
0��X )n��u��/e|!�$F�f,*��,�y�.P�5
	�T!�$��l"�1*�B�$U�����;�!�� b��U��$g � +EbL����@"ON�;���PA�|Zbπ�ռ@��"O�1ڇ-��cZ\
���2����"O��9p.��R�B���h@��P�X�"O�Z#�!i'�] 5FΒj�
�!r"OZ��G��lY`�98�x$Q�"OB����7D �B�^�"�;�"OR����A�!߶tS ���$���3"O1�g/H�1��B���^��C�"OЭ)�ȇ5!n��q�6�����"O�Т,�2Ղ��IN���d�O� x���0>�UOM*p}�UA	6U��eZV��U��Z$��3xѨ��I�R�|���)�J����œ!�B�I�;et"P��������$@&�O���M3&F(��3�G��H��H�'�9E5��a�b�P=��"O(�5�
Y�RMC�KZZ芥��N [9�h�ծU�<��.J걟�'"D`ұcZ���J&h��zHV��'#4���EV�3R
D,��1%��bN������0Ut����Qa{B�_�(�c N�=5�	�����p<	�N�:0�d���(4 .��ߴy�����W�xz��a6�X�ȓ<��5!�����E+g��:��ȧO-��NU�s$���WG\:E'�"}�aFL�aE 9ƍ
F�Bt�J~�<Yw];m��!� �?_��u���p�΅��H� "	�8�n��}&�0#r;ug�K�O�r���ï?����H�@tȳ$A�h!�Q6b��.w���OE�:GX�FP\؞����͆Q��9G���4H��)OB!rgH��J���i%ir�ѬA=�8K��ܮ5�b�K���ya�p���8êU0 /����6��	�aRL	a�n�.��S%��=��e�@+\!�/)<C�I�b�T(N�q~8!rKٍn�$DfA�C��-d3�����L<�r���Ԍ��/Ƭe220QAGh<��=F����̊d{FaL�{I��KT�#j9� NlS5n!x�V%�X���'z�  �.3t̓C@���I�2uf|�t(\6�0H�ȓr��{��G0p0qp�³ʾ��=�#YcSj�S�e=�'z�*ᚥ� ��3G�+JV4��Ht��R�� ��1aB9l�фg�$&��O <x��Y�Z�b 2G��T2��.V���:q�(D����r�@�2�$ =@�I��6%��t�A�/��\�CT�%����C�U�m��۽R(� b��zR�7�p,+.�e�� ��2 Q�D3.�XK�@,c�Ṟ!
O�Е-%\�iОkkX,_1:%�=q@a]����P�ˈTo�)��:�Ӕ!(�<8d�r�j���\%)�B�ɪ1s,�����cfJ�Y��[8{��2cgR�@/։h��U�&��7M_�����l.u16�ъ}� ����xZ!��iϔ��(M3c�M�e��O�	+n��<�@Fۇk]�U���'�\``D��P}0�M��$q��8	��>7@�qX�>a����$mPD�'�/@d�M��3�b�U X�r�����T�)� 3R-�p��("
b>ћ���^��걌�?�Դ�"�:D�d��hQ-E��$8b,�W[J kq-�� �$@f3~��r�>E�t�]p�Ȉ(���$�b��a��6�y�Ĥr"d� �+��-فJ��	CR4Uc��_�?[ax�Mr�`���*JJ<�QT�	x�vl����,�.���K�&�Rxb,��#v��k���3#� �HztB'�D�=`R�0�N��*V��D�I����~Z�����~�Y���2D��Ke�E_�<1Â
�XF h�/��9���X��n�<�4ď���쩱`I��2�$I�g�<�3��ZiH�A�.oBD�hW&=D��v$^�̽�uM1#�BQj�A.D���c넶e�0�A�i#V�B��E�,D�̰��ٹ\�P����WYL��r�'D��`��Ÿ5G�Uyw�[A�`*A�$D��  ��b7�<]�6���H�6Ȱ4"ON jm�MY�3�,	4A��	�"O��Ā�H�z���y.���"O*����2�
��� �H�J�s@"O�EK&E� +����!6&-C�"O�E�)C��H���5\Α���'��M��D�S��1A֢H(=���N�0�N���v<���W+���G�2'72�F~�	!D�pH)@�ɏ�CL �ZF�����O !�$ҳd:��kg��<��x�j��ܻ:���7mF���)�'�� z�N@�AZR��懪tf�u��b"�:A�ɻV@Tir��H�ht�O���R��7M�:��Ó����D�:4��z����2�����I�?bfx2c��l<�7�7X��aQ�A8X�"��aO�DN�F�>��"&V�:o�E����B��y��?/`1��8���{x�(�do�m@�l��"O�,��P��tmqQ��,?@���OV� �Dl��D�<�O�:��#����@��9`����]�P��"'�O��8����(�����\2+�6��C�0�t��ү�>q���6�Y�%O���U�ێ�0,A���(WW�b����Z ��`�ʃU^��3�P�q(�
V�`��f�TF�r� 4��I��x��V�z|0"�����I���O��~�cm����͚u}��!�X{��I�z�xc#Do�,^#PR	�'�V��a�Q�[p!��f���z)OL!w��^��5zs�%�d����'V�Õ��<����R�O�a���A�oh,8���e�:�G�܁+�������i��#�	s�R�Q�\4��
L'ujN5��a2�1� �{%H�!��b>=r5���S%�̡�%L�v��0�Si1D���%$7WݾxA�NT���6����ʖŊsl��>E��D٨`<QG�E�p� EX��ߖ�yb�_�2�����Ip�9×k����1�J��;vFax�����8%I�����Ib����?I��G3?�H�b�/=/��+��p,�6�
�Px�AD;/k8ehGF�3�~c��R��O���᝙��O<����Ď�7F��:��!|��x�	�'�l}�f�K�a����;q麄i
�'G�-��n�[�f����(_��9�'ɪs�j�9u����a�Ĳ{�0���'dH�������0���Od, ��'����
/�챨sk�<h�	�'_0`A�d�1��P֏�(%�j���'8mC!LP�Ԡp6D�:ʶ�h�'�)����_�4�+���>{�d���'��e�T���@�p���$�8��'�`�)0n����Z��H�(���'�ܬQ�^����aS�@��I�	�'p(�)Cƚ�!d�22��<&�b�[	�'`�t�P��={����A�;�h��'��#�0j���!C�����'1�pw �[��Q "o@�Nv���'���@�K96e� ��P;r4	��'o�,S�G,��!�ш��ҬS�'�8����!��괊����2�'������-O0���H�qbd��'k�c,y�¼QÍ��s�H��'l����IO� �BXB��Py���8�'ubݙEk�')��*����T��
�'��؉�GѪw�yj'�֛i�yb
�'�RE��Y�0�=��1?���'GB�[��	�X
��
2L��4#fM{�'H1"�l�n5d3R��0�����'L-��Έ%KO��:�ݭ?�.`�'{��r"HH�Py�`(���r�	�'*���H�)��"Q��"s�zts��� 4�g@��N$��$��R1`Y�"OjT�ɓ�R��1w@�e(p���"O0H3��0H���ԠS�Hq�"OXH���YA�}X�I:r�8��Q"O\����!B����DO���QY�"O�`ڦ��|rpȢ��00�~D���d�7�`x���%j%t��0��+1O�ͩ�̌�z�	8pI,�`��"O:1�CL S����s�S���F"O���զ"L�8��@� 	��@ "O�-�u.�SS� "E�	C�j��7"Ox@�Ԋ�>g|�u� %K��f�j�"O܄1���'9�4�9�m�q�y�B"O\mR���-y61�c솣ng��A�"O��rA��m���rk�?\>j�"O4�ρ(hI2�5@FX�Q"O��QA%&B�"�q��&�|1	2"O %�P�Ň;v����Ǜ�T�Q�O<С�.�)�'DH\Q���  �uP�d�b@�u�4��%<��;}�INZ���)�2t{�fQ;Az�i)G!�%�p� 0� wy��\����S�
�䨛���8B"}�2NB�.O��(O���E��	 �8�ç/L*��a+�!j�����%.*,}�'�UӰ��&>.uYq�;�'/M(�C��~��L��/��S�����Tӛ��I�IF$T�m��Xa����0|j׃Tl��|�f��<;�,�Sr	�ɖ썇kǜɻ�����ӊ�\@�P�>^�չE/�#O
R������ �a��]}���6��CWA[`�R4 㮼�d�M(|�>py�!Q4w,A�'w܀ʧ�O��1Z�.�DGt�eD��8�f7u�)r��J"#;�Ͳ"�x�s#�;�
�k��(gӴ���ʄ�7Ϛ4+S��8&!Ȍz&m۟Y�NLp�	32��)�~�v��p�)^���X�,T����N�.Δ�e*��@A���Pp>�D��I���PI�5h��|c��P�nAv̓�	Ϙ�fX�vI��V�����	u]
�h��
�X/4��D���q�j�l��>X���&v��:$�1�f���"pl=���)�����>qVkE�>S���˓pJ�US'̷e�^@X���t���@��fʆ�y��j�'�hX��m����DR!�:���ŠM�5��{H��˳�=AL�-�1f�_�����zg�T)0�DE�A֕OQ�ȓF�����|l�<�3#;� �ȓ�(�e����D�(7�D�g���ȓ��-��F^�;~���O[,C�24��N��uO%h� y�w鏱8���ȓ��0����-l�Ĝ�w�A�~)�%��px|�t�[�L�Qς X퐔��t�J�P���lOJd����%6l�ȓ*�a�T�Ԝ
0娃��"(T�u�ȓS3.�Zś".�\�xAh'XT���ȓJf��0ЎN/*G��zBgA���ȓl�zr/Q�%����� JV�nq�ȓqZ���D#� E�Fn�,E�  �ȓ���1����X`E�M�Z��ȓ���&H��9�@!�M�.$wz݆�ɮq���S���A�c�ʴp�-�ȓɂ�!�"&I^��D̰y�zɄȓR���S�U-"�8���Ù�1G��fQ�d����gG ��� �sG�Q��^��y����w�x�#�"aAj��ȓ����dւ�  �1Ɯ�K5�Y�ȓdB��fb .]1+�@^!R�TH��(���[P�
�X��,V�&:�`��ȓq��I�
_��#��G�^���me&�X�.��S:���P��P��a��7h��K� ���.Tb�ރ!�Ňȓb�H�)�	�I��t��j
⑇�}i�r �6��(`��"��ȓhX !Y��$!Xt� B�}�$���S�? �EK��ќA�8��s�6���"Oz��6Μi7nI�`딬xϬ�s�"O�I�A�/!Z�@��j̔l�HM�"OT*�!ܚ٤�ǚ3ѐ��"O��Z�Z�o.5��сV`@dpS"O���vIF��u��:E|nA�3"On����E�\�`�I5���D՚���"O�X����'���䈊lZ�PB�"O�	RQ

�7��J���Wd ,@"O�DbkH�st pCFlg`��X`"O���vϗ�5�H�!k�i�0�"O��"�DU�H�\q�����,�"O�pJ�@�ut�1��D�#�ޤ�"Oz�� *U�X��q�敛z�~��"O�u�kE<��)���I}��Z�"Od%"��"
4�"ΩN����"O��x�Ʉ j7R��aش5�X�j�"O@\	R�ғ!�6��Q U, �,Ղ"O��ؗe��+��Y�4��"O�����D��1�5��|@3�"O�I��I��hU�1KF�+lf�h`"Oҹ�鄁7d��1'F�]p�"O��#Q���m�`����=�$ݳ�"O�m���<M+t0��-�hq��a�"Ob��"�V���#�ZϲA�"O�J������x���h8�ȓ\r��ϹAJ��aC԰~V�%�ȓ�|��� �(+wXÆ�+�:@��x:�yŉ:`�h�rrlV>h� �ȓ�P��I���"7`�\���kL�1���1=�@���Փw���h�n�@�� �g�2vlB�"O�T�e��6|�vI��Y���ɤ"O�}9�+�'�}�BG�&�T帢"O��� -�	V�\P1'�A�-Su"OZxz��X���C�&�<Z�I��"O���e�2{"e� Fܒ,k�-I"Op�6'H����9D�ùr�H,0�"O
 kc��'%E���m՝[���H�"O�9B��1���4KL�Pc��Z7"O��(�K�:P�f�!�)S,$�R0��"O��U�o�@�{��؀/�z�Q"O����H�P�HH@�бD��8�Q"Ot����$q��0zu�$G�q)�"O�a5AM-\�@}�d�1~���"O�@n�v[�2��ٔ*��y��"On%�����A�$Q���O�����"OH4�g�	�8�4���X�,{��S�"O.�a`@U07��a�g�Ǎn\��"O~y	0�B�?FDR��#$��=j�"O��*�f�2CD��UNT:��]�!"O�Q&�M'D�|$#�� w ��p"Ox��,!�XEi!�d_R��"O2tt;ӎ�q�k�nYne�1"O
|��eJ"Z�l[F�K�_;�A�V"O��7���<��c�j
D3��1�"O�5F��BD�s��*F4<+�"O ��� �&W�` ����+n#��p"O4U��Ć<���"��)wЩy�"O������:������'sD�"O.���} 5ʄM��SHZ��"O��a����#��
�O1��1�"O6�1 Z�`���D��v�XI��"O�u��c�k� 9Qd�J2�Bq�S"O� DL�`�H��n��ՁP�����"O@��Ek_�9Kh��U.ʦIx4��"O�(��G��@Z���� !e"O��7��;�֐0�!�)e���"O��K,L6c�`5��� D�"O�(Q���y����]'9��"O
a��.�N9�����X��\�B"O���D`L�A�� ��mX5N�rQIV"O&E���҇O�q@�ݶ2}��Q"O`�� h8_MȬڤÒ/�n�a�"O�	�Ԩ_�sF�i�GCL�n���H#"O4�B$�5<�1Q�L�6�r��"OZ�٢���!V���!Gb�UjG"OH����64���a1 \R�8�"O"�1�b�Y`����e��"O��7e&c
N�k�'�C�>4S"O�!�-��i>�}��G�")Er��c"OuH�H�A� �16�S V?@���"O���3��t+��I��\���"Oj��ѝx���s�#�,Rj���'.�B��sB]*�#�.�|�K�'����CF��lo%C#�3{���'���c�g��%�@#J�k^y�	�'��)A� �L�����	�'��1'8��h &	Du:;	�'+���b��X;��7;��d��'��9A�i��.�A��?A�m��'� ���
�=2B,1!�@�0�c�'�U��NF0f�`e���+$���'S�=Q���&e�jc�˴y��p{�'|�|#����J��2cݳmD�� �'�&$��Cн}	&qS���dv�U@�'�L���I�^v-��Q־Ѹ�'ي��6Ĳ�ѱ����$�0�'�f@�}-z}�!�ޝ#�6�"	�'��D2gN�$ת���æD����'ZDP�.ZXG��1E��q�'R�h�S�b���S�d����j
�'��g.��g=�LC��ԥJ��	�'��� S$�=zЂ�C�مH�R�	�'��0����-2��r/�?�:�8	�'
��cE �6��X�
\�8q����'M�q�d����J�$65�i�	�'�vH `+׺;-
���4���"�'�������"T:�c���b�J���'ۦla���4<`���T6Ĥ`	�'����m���`�@��bk����'M��J�H�-�@끅����'�U�u�M�PG���nYְ��Ib�<��L��*���e�D�w��w�<i�L,���rh�	��52T'\I�<�dC�x���N)3��9����[�<����0 Q�ʁ�)�4C$�Z\�<A'X�U��(��4�vp�7m	Z�<�0H"c]���B�QZbе�Q�<�ԉPS� TP#A�*tT���J�<I�狺�jA��Ά�+��l9�]M�<�O��$�[&[�^i)ӌI�<����2�4��6C�q�D<)��\�<IףE2k��*�,Շ��i�AAX�<i�L�/��I4�C�8�h���QM�<Q�ɟ�\iC���v$�&��}�<)��\"�d0J>z)����u�<�U��"�t����� �4�	�)�r�<� x��2 Q�s߄�;5!]�hL�l��"O�$�W!!R�б:�`�^�T-�4"O�15ǜ4!�0ා��1'���"OL�0�ŝ�j��p�t��8W%�""O�˰BÈK n�i�P�H�@�"Ola��'�	��:Æ�P��Q��"O�\�0�K�`F��`1�̍z��Q�"O���4�I�8Ȕ�ƈ7`�V"O(�;��/Sm����FQnKء9`"O�`���^[q$F�[9�U"O��B�/^ R���iZO��b"O��G��_ޜ!�R�Qu�*O�$�e�:&.� s%U�nq�a��"OrA!�N�VZ�z��6g��kW"O��Z� ߈O��T�n�&�Q&"O��R`a��`}ޱ3&DP�z�"O>�hG��]��I���6Q�	"�"Oj\���l��,�E-�	s�8��"O��₇ :�ݺ���/m�J=�D"O����+f�����\�N���"O4�J"�R�B���6FI�q��a�Q"O���CY*P��ׅEn��"O�A�aO�3A�^}���Ͽ4u����"O�}"R�L�>4�[RNӲB�)8r"O��g
S�`զ�m�+K�S�"O4d��F�Mf5��̍l�j �'"O� ����;0-|a�񋌍w��-�$"Oh�4�
"p�9�)�'E���Y�"O��ɳf«%¬D�`I�&#�29��"O��x�N��*�����<3����G"O�p)G��(u��V��Qv"O�كEY�P�@Ę1k �E�:	�b"O��  �Xh�Q��J=s�ĕ�5"O`�`ǃM4~�����Y�tX�"ON��E�?�4�k�F�a��q{C"O�m��   �P   S	  �  `  �  y&  4/  v5  �;  B  TH  �N  �T  /[  ta  �g  �m  ;t  |z  T�   `� u�	����Zv)C�'ll\�0Dz+⟈m�Oh��5G��DB� �8��GPz�إ�7&=Ĩ��(C����AL �$�e��I�{),Ȯ;\����'{��@��'�tp�g/;�ԩ�aIg=ZaRFT>*��m@�I�5iR^�i�7�Ͱ����LsA�럒�D��.P]!4Dљt�rh�bO<[V��X�̈́�JZQ�	>�I�
0
!���ٴ5x���?���?I�'�2ubAC���V�Z3m�j����?)�%�>K�R��,O����"o*�)�O�牵s�v4HP.F%P��l���ԔZ��$�OJX�'���'[�M͗���z�t�jBzLF�H�*.h�89�r$9D��K�V�N����,�� L�O���g0�A����Į��u�㙖/E�ٗ'�<�ӣ(tI�D�	�
�ry*��'�2�'���'���' X>���'%���	$��h�
�g��{i�@�I��M1�i\^6M���	��M{°i~P6��A��5s��(�O��ɩ����zp9����9�ȟ<̻�	Γb���*�P�b��%�ƚ
c�\;��ڏǤ)uiv��lڊ�M������c�-Q��T���mx$��2Of�⡃����?��-A(/b�=`T�:@%���#k�q�(�r��OZv���d���nڥ!x4j�n�0��+�+�|Dۦ-@�*O"uK�+^�M�v�i��7���*�c7/ȝt�6H��#ާD����~#�\ &�3݂�� ^�}k,�7bH�db�$lZ�M�$�i^�51HY1��x�;O�4�%*��[j�Pye`O�\ѥl�>-��D����Ȫ������3H˲��	W�:L|a�%
B\Xa���%;@aB���'�|�藝���%�XM�0"g��(htd����$�y�B��hb�@Z�!�� � -�y�@�?G���8�瘁E$� ��y"�@�Q�ƑSU�L�	���3e�y�+L/t�0�!�W=s�F0�'����yҭĤ[��p��ĥh��9�EQ�hO҉����\CZM(�������A�4�B��6f�Lбb��9���&N�:b��C�I�A0}��/C�!
�帧, @�C�I�(G8}땨�>Q�1@+�(`�:B��"Ze�0�=o=l�F��"WB�	�NP����
<��ȡ?���?!��"~BQHN��ʔ[Dj�X/�li��-�yҡ��`��T:��HJ�̝��D�y@�	�����j:>��0 �)�yRe�C�$\�Q�2߶U�M���y���+�`�'D7W��t`���y2O�k�}RSA]Y|�9��lǉ�򤒺
��|R� �5VY1�M�WYr	�e]<�y����}��MF�:W`y_��y�+2u�bj'�r蛢���y2i[�h�t���ʎ�d9����ybؕ_ Ȩ�QI��\���Њ���<�a!X�X���'���
k��,A��K�4�|���!K�o��'�b�Z��'�0�X�0@�Z5&�<���'jp�EHW?@���8����:�̹F��#��MF~�HI?� H�g���?�ܼz��4�ɳqq�
snt�L�7f�/
X�D�A�P���|���m���C�ウzhݹ#�/��=HDC}y��'��OQ>�ZŦ^�~�|Ѹ7�ʿ,$��g�'�O�i��A{0ժ֧ (+R��A� 4%��d"�d�4���C�9O杣>cV];aϖ4�� ��^�c��C��%�����ꂍ,���3̗*9�C䉞g&�[,��up|j�!��y��C�I67Q�B4]���!+U��LB�ɵd"���%|<0P���9�nC�	u�4P05�7S�8�����E����ܺ,��"~Ұ�<vI��F��#8\����y�&�'�f`���#|���-�y�fC"��!2���%B�yEK»�y��/���:ŁR�|֔� ࢙�y��E�gqF	rE��w#\��Ƃ���xbe�6&�����! 21�T ���d�ze��'a|��VN��9P��B�rV�!��߰kdx��'�&�q�V�W;���'+uQ�F⒫�xrGV�U�|���6	`�(b�%"n��HA���2d�y��)��]u��#���y�,[�M*��8 ��1��r3��n웖�|R�B��y���$K%���+�w���X|I�?O�� 3�ٰ:���O� ¤�tMěc3��#$k\�0Z�&�'q�
b���n��'̒���+5 o�M�hS�|�
Ó_x���	��	П䚂��B��!θ	�SDPMy��'��OQ>9{gB��6����'��&Q�m���$�O���	*I��)XD�&B���u�=3r�$�<�AK��?����?i+��a�� �O�Ms�퍭d(b��z��<s�e�O���1�R<��B*W\�b+L�dg��O�S
��K�H�K�h��I�H�6a5QtLx��#��8n�Z`��_�E��=�O�v�
�J=(������%m�D��Oũ�'x���<	�㜉/7j Jgkʍi���J"�`�<1��	E�R�-�$ ʈ�+]�'ۖ�}�bӼM<Ctk�* n�kĠ��D�O��$ g5>59���O��d�O���l�a�e�)G8 �;ԪQ�M- qiՁ��	��M�1R��z�O��l��/��v48�Z��Gˎa��1Kh��bC���`|b>c���PN�|'��b5EZf,i!���OMm��h��L@��x�|�'ra�+o���d�+m����U
��;^�{�����p��:ڊ� �(��Fb�,�M������������b��9 l�j1
�	�Ŗs���jcT��$��/HEc�%D47}���F[�"�!�H	fl*����/`L���$��!�$@7CE�X�2IǶbJ��5c�1�!�d?:��u)��d/u��Y�1�!�DZ*S�Z���
4N���r���*��}�GL1�~����x*���1�l�r6G/�y��٧j��)1� �w����6e��y�!I kH�f�Tl��LBW����y�m��z��D�i���uaĔ�yR	2,]�ѓ���2C6���ޔ�y҂�HO�����G2@X� �$���hO�H[��ӱ�Z���$^3K�KG��9Kq�C�I!j�`����<��! P�C�	-Ga"�0�ވD�b���p5�C�ɨN�Cd`�.#jk�eXbZ�C�	!�n%	��X-t�� �-�0Q��C䉕)��ذ���5,�U���
� ��Q�t"�"~���Ŗ��bRO��Q�m���y2� �6=I0�
2�mZV,5�ygԝE�,a�֏z<x��Q�y�AC�VN*��k�̨���T��yrbU�]F$y�rmƸ_:5hd�Y��y �<�"�͡.�Ͳc���DUIx�|��g�t1����c�湰�œ,�y�F�C��� qȑ�hs&�iRΑ�y�*>F �Sk �(��I3�yr��@�u��̝bTн�m��yBbC�O��M(���0W��)��G���>�c/�^?�l
6Q������<$r�Ec��o�<	go�75�p��	�l�MAҌ�h�<I�4��Cυ�y��Pd/�f�<I����q�P3o@�Q"}(V�Qn�<�e�\[4����oڄ}�l�l�<ٓe"�dupц� 5~$M)��p�'=����i�2cdc$I8�^�3�#�)�!��+>Wr ��ȁ�Y����'�Q$+�!�R�_�<���O������b·s+!�Ĉ+�NQ�1j�<?v ���AB�R
!��<n$�fEܷd��"b�3r�!����rH��4�K2T�u:v ��r���O?! KG(h��5��cR5e< 	���P�<Ir�C
0ӈy���΅2�֙"�O�<)�*Ǣ	�l�3�H��@d�g�BL�<��B<g�b��be�;g�5 U�SC�<��I�݃��CZ��е��i�<��&З�B�p�G2{��<JM�dy��p>�1���|X���E�	�ܪ�B��y
� V��������3B# gY��i0"O(���U�.��Mar�<7bdȣ"O�ݹ#M�	�����H ^���"OX��e=1����u�/?F:t�'�����'���R7a�?���*_�q��'F�ٚp卹& h�3�T)���'�L}��i�-v�s�i��c��"
�'ւx!�� {�T	���>#��D
�'���x#�R���Z�ߊ1�(	�'+v��v�Ɩ[ԡaӤ_"�����D5b�Q?i¢a�:F����F'L�]�0�8� D��b��M�� �c�]�K�,=	h2D���1R������ꂪ,D�̓�l�5E���E���g��m���(D�t��`V=C��:�M^)irFlj��+D��藪V�P)@�g�\�Yn&`Q��O���b�)�ZL�a{�̃�)�dI��%�3 �>$��'\�!�P�[
�U����t��%8
�'�(D��o�;cEŃ�G�Ԡ3
�'Y�q��� �#���g�<Y	�'w����C� ��6"�*�Y��'X�P5F�2���Sa$��� x�*O6)I`�'戱��@��Te��m��}W@�
�'X�L�wk�w脅��eX!,��Z
�'a�� �&l=�pчI&�
�'�@4��,O�$�"�����i	�'�1�O��;�9��Da/�����U�#z�z�E�o:��A��-L��Y��O]D�s�*Y7D��(g��)M�9��o�tL6 �V���h��k���ȓ=>x�*�˓�p�j�92�,��(�ȓ^\`��6�)�d���愃u4	�ȓc'�u� ��Fy���(�<x�5F{"6���"��.�*���.Vu����"O<t��f@c=�t�Gc&�d�Bs"O<�if���.#�d"bl��denL�"Oz��A>��P�ԫ��{��\i�"O�m�TĎ�����P#�d]QV"OVɑ"��T�l����D� 	���'�f���� �@Q5ק"$j% ��L��ȓ,���[��>�7!M�Y��ȓ��T�a#��xdH"狛�z��ȓ%�x*"���Lx�`��;@h��L-8,k���!Ec��B	Y[b����s{��P �;�0B�*ȩI��'��8�8�b��틊P�a����1ĠH�ȓo��2g�A\��q���"Zi蘆�_U&�Z�_`���C�ڢtB ��ȓ:�D�	�ad�\�0��T�@����A\:�����z�\a0J�5:J�-��I�E�L�	�c��CU�E,$�lDr���-]ڀC�J`V��nJ/oBL����#7RC��
V�����U�e'4���#z�^C�ɴ<_�q�6��`g�U��JF�%�(C䉔~��Q����'[��P![��B�I�]+�Oq�~0ȤA38��=q$�x�Oh��cO<]���Z�(��(�� �
�'� ܉�μk��S%��� >A�	�';�Y�wٮ�p����g���y�	�(�8���BR>y9J�	6���y�ĖhhR���"j�������y�fC�\W�����U�9�z�PA���?1�*�a����r@��q��X��%1	(h�C>D��rĥP�W�B��'P�\����M;D�� fH;1��X��4��%�u��X�"O�e)�@� ���p��P�� ��T"O�@r`N�s F@�vc�!�J�h"ObI ����kz@���a��;�`�T��2 8�O��3�j@�`�����D�z&�"O&���G��Qт^�4ܔ��"O�����L�n����9��!e"O���E	�/~Ֆ������&��G"O(���#��a� ]#D�	��'A���'��d�VHˋ\Ɩ��7BK�[���'`P3%#ZG�d�Wd?*�"b�'>�5*�%G=O5 �d�%|�y	�'��mP��^0����!,�tw<`b
�'g�����P{���7�:p-�)�	�'�
�1��~�(�G%½��mӉ���}
Q?u���
$�d���\��`�! �$D� �uˀ�W��`�\=n�^�i&�$D��pe^�b/>,!TJ�fKX��b�!D�Ī��@�U�����o�cĊ��$�=D��Z����\ٚ���=K���d�=D�, t狵<�t�6�W<b��&N�O@�0d�)�/2��@��A�'U@��u#J8V���'��4��'ж1Mu"���X�J�'$��e�A�v^�t���P4&��'�&ip�8	��f��5$��X	�'N��۶��
������;*�9�'b@�`�	�e�<�aE˖�<`{)Oh�	7�'�j;�@��/kU�Ȥ�t���'\|+fͥc�:�e�6Ɔ���''��ۑ�S	4!����Ϝ�H�`M��9d�!��+0�B�H'��"4��ȓ��Q+���U��@��Y��Մ��� Y6�I�$ i�t�?f����Kz^dB��#=N<�"�dS\��j��͚,`B�I�
�"0�k�]Cd����.B�I�����,�f�[F�
e\C䉌7lE�7e1%�TՑ�	�3�C�I�%��c���h����-C��P�=�f�X�O���)������C�/�ձ�'S�4�*#pN��/ӳs�Z�	�'b����IW�5�}�!�-n-�p��'I@�yŢ��T$`����O�r�	�'��,��+Nzx�45T�qB	�'�N�B���.|��� �
� �p��KҀGx��	M�7R(!�!Ł&/$��C�3r͔B䉿t���"��+^��'X�$z:B�I�;�ht����o��C���}��C�I��)t��+4�q����%��C䉃A�V�Q�˭w(��"*�:r0�C�	�+$�i`F��S7����C�_f,˓I�� ��I�O�Tak�,�B��b-�9�C�	�w��h{�!� �2��N�8RB��=k1��RC��]��آ@ML�QcLB�I�=�1�����-VB�ɪ/�Xl�� ����dT��$����5yz���/���ڧN����0`!�&4W���@C5;��i!�W/Y2!�$�7��X`� ���B��q�.>!�$]~:D���'�?��	Z�� '!�d_�w��$ �E�M�2�*�
Pn!��/#����-Ŕ,�tiȱ.˷\ў�[$7�_�v�jwi!1X�1�V�Q�����+�NĻ�:0������E
����(��(�d�/#ޘk��%6�,��S�? ���į��#m�L
uk�((���*O��xA�\|<m+�"9	�����'V��g%[]ny)È�p��(��4�ȬEx���Ҕ+Vb�j�FP�2 �,�4C�I�������T�ڹx���3htB�	�"TJ�"�!u���_�3�jB䉏h��IH#$��5��a�h�/_h�C�I�N�4)�ՅR'	:n]k�*�
`eC��.hZH@�ʫ�PqI��@��ʓWP����	'm;�P����-U�JY�jޱ��C�IqH�
\�N�t���� 0H~C䉩9�2���$R�O���9#J�s�C�I�l��B�oT��v-"܊b�'�nI��	�V���b���~)�n<����]��XBWi��' U��f�H��ԅȓ5���-�C4��!���h��u�ȓ4�Hx���S�cp(a%��&��Շȓ]�h	�hɱ��t��/ ��ap��] F#䀑��Z:/�����s��iɦ#�y�r�*d�C6_zZ�F{�%�������ӊ$0��yp��;q���"O��V.b�D�F��;CeZI�u"OtH{%ƃ�B=y��ͯW:\�3T"Oȼ�S �:
#�hja��$�8�T"O�᫡�bht GL4k��mµ"O`��f��-,��K�?p�(�bQ�'Yd 	���D2�<����8I<��o���x4�ȓn�F�G��{0^R@N�5s"n���`e�pS�Þ? %�QR,�-k��!��!�$ɳ�SmP�m�2R�$�<ćȓD)��+�〄��$�D(�Ɠd�:W�\���a��C;-�̨;����	8���u����'�&���d�%�	7+�HA��c�TLZ[�şP���T��(���(�G�j0���aܛd �5cDm��N2{f��ؒL�����;	��9�E�Bݎ�Z�'�(جAc��^S(<��BE�$���D��)!F�:5�]!EJ�#<�H���	F�'m��I �D�2&���s��;y6��'�a~�(��\���2�*�@7Ȁ)�`���>�q_��T��.t�V͂P�0pE ]sԨ�<U�]0�?���?�)���As$�O�ir\A�F��n�1@�u�g�B�8+��i����O�����S�t�)R�e�6��NN�L ��p�dZ;Y�d	d�:���Dc,d�s�>�'Q^�(�g6�`0$�S	m���̓}r����ʟ\��'����_<d��/�|rUS�!E*�!򤁚TFV]����&hN�9jd�۹=�ўD����ȫo�U �)����@�� �L��O��d��P�����O��$�O�����N���{X�h��eY�K|���@������D�]0��d暷8+:ˀ�3J��䕝F᰼s���7�Zܸ�EZ=}��i ���;Q�0����EkXhU���?ݻ�a��,�h�oO�KL&M�8tp��z֜��'��q����?)���p��AW	�1�kP�5l��A#+D��c&ײ8h�xB��1~��n�O��Dz�OJ�U��cЅ�$�B���%Ճ]���T(^)_�
M#UgD��8�Iԟ���6�u�'^3�ܥ�'�D� ��낭�-&<ɃBCA�:l�S�8��t��I  sÚ�:��(�F��&D0�P� ��+�ذ=fJٟ� h�#݊a{�	54m�LП�E{��Io6�p���{����L��MvPB��
u�Zu���_��i�THÑ&ʓS�V�'U�3�����$h>�A�ӫU����T"� K���O(����O����O��8���+/�!��d"Ҝ�i>�R"�̌<��Å�\�0ZD(�%L9�r���O�*XА͒=���V�g��x�g4p��	!ٌ@>�Ē���O��D(��
p��p�Հ0�d��vFΝk���0?�`FPD����A�	UD�R#�Ax��C-O�	�uE�vW� ���!S��q�Z�tQցIҟ���� �O@VY ��'�r�S�6>
!r	�K>԰�Ʈ 2���
��@���N�6�է��'�SK��ъ�#�R�H�	�8BN��I+ٺ�K�ˈ�4�r5*�O?�sv��3g��'�fպ1[�jy�$Kp��O.��=?%?m秀 r�FK�.F�ш�� l�)q"O�a;�Z�{���1�I��b��I��ȟܙ�I�l�^9 �ҍQ�,�Y0��O�D�OF�s���L!��d�O��d�O ���O&Hr2����\��+��:��bk�<����Q�
� ��P��8;���#V�O`���"B�u�tC%+Cx�+��=}p�A!�'wk2<� D۶F�� y���g�%?�#���@�!�ޫf��`Xu�J~�#���?Q���hO4��r���@ʇG����B�#�B�	2F�X!���<��ęG`]*)���d^p�����'h�?
Z�4@q����e`�9�܅stI�8bu������I����S̟��	�|��Ӡ#�X|I��1x6��:6�LWH%c��]�����t�'�&l���<e�<�qV+
�hV���0OB]�"�Y%�׋W�`��$�0�҉���F�J#
b,(�K�G�"F�B�t�'r�@����^Z�����^�� T��'-b0��Kf:��8c��n�~��(Ofo�ٟ�'��,SP��~�����J�R1N����5��� �Ҫ{����ޟ���(/9r�����m�ty�d��47؈
���p��g�L��|�u%KY�v�	��^-�Ta���D$�פD;K�]Q�o���<�)�n�s��A�)�'Z8q��ğ�|j��^�-���sU	��Y��kyr�'�Dl�#bb��s2�όORbl��0��	 2%J4jU��ʀ��d�T;SG���?)���?���L��AŗS�n�ڗ�)Zf	ZS�5O��=a��Wi�5��Ig艺�j�e��S�Z�%���~��MY�z s���"������x~򆧟���0}*���\�m5�z���s��X	Ș���??��>���[��i��]~�<��E� �(\����>	��O��}Γ:PŚ5$Hj�&�7I_�p��sV%�S���x�$V� ��5�SG T�Z'��#1��v��x�R��U/u�����D��*Ć8��Hv��>8r��)�i��P��I���,'�'(�7͐�-X�D�4cwϔ��&��E�I�8y"�'�"�$�*�� �c��-9�ً����O�������S��'��X�O,"fW�*Y��[���r�ȑ!br�#Y�y����?�ED�<)��ī�{,ر��;��0�k�?qQ���d�qo&?��y�f���~B/�V���6��܃H�?ɑE/�O�a��G�/`2h�6�"/30�V"Or��S��5#GPM����`#N���i}r�|r�'p��N=O�R�r���x��*�O��BPn��$�����1O�ip|��.�*?;��I�|��E�M<���)��u4�a�b�$C(1��S�!�Lb(�0"�&(�E3#��]�!򄊄df����S12��� Oż/�!�d\)K�N���DA&�( ��Ň!�D*'�,�Q*�:�F��!�6
!�d�43` X�P��W0�3f��!�(R��u���(BT&��u�X�=�!�=L�b��0yL���* �N�!��t6�[�m0oB�1`��5!�S;	HB�"���,
�CR�G!�I�rfp�Ui]�b��{@���!�䆘��m��T���h���72��O���^�27HY��^*}?ƑI�NC�e|ҵ�3��z�LT�Q�϶�Q��%Y�t���HF0���a���a��~�����^f��k��|�)'�R�rZ�P��+ƙ7�>I��D�G_ ����J̙iך��h�?��={��N�)��w"�,��Lr��꤃�R�n�:U�ߞ)�T���Ij�)+�r`��l5ze��釛X�i�ȓ]i@��"ؓq,�(/��) � D�8s��VB�|�;tlW�ˆ!��#D�� �t$��c�<�j`!��6D���O6N�&+BO�+|���!s�4D�P�
�;��!�!��=3�d��ԅ/D�xJ2�W��D��Y�8�� lŃ�y�m^�s�
�o�y_����¼�yRNG�l���D�E]gK�y�	�g�ll��B��8��\��y��F�N�StJ 	t�F�۷�y�)f����쑯}�xĘ6���y
� >�k��ˍf{�1Y.�$z1A"Oa��eP*)�>�`�MJ�g��`�"O$a��13�68���� O
츁"Oh���版�2���_*��U"O8h�Ԯ�(�x8��ԍd�1"Ot��E�P{I$\"�����"O���C��f$����!�R��"O�|�v�(�ABC��	�$*"O���2�̕|}�yPb�)7�0ՙ�"Oh|c����7HdJ֏�8V�D�0C"Ov}��C2S��X{�/Ծ+�$)"O��j���zb���s�1D4@�Xa"O0��垸�t`����#'d��u"OH�D$-����'�e#�7�,D��#S��Y�|� ���,c�H,Y��+D��1�+o
�pI$#_/##�xѕd<D�|J���&bɈAb�o\�5��D��;D�0F�&Kr5���Z�(֔I��7D��Is�S3m��Ih��Z��y��n)D�4I׌^�B�`b�$E]68��q�(D�8�ݗZv�����N* �j#D�d!1*�*^Fh��m�17�y�B>D��K�%�6���Q6�;V+����:D��#�-�7����p�[%}8�0A�%D���C�/���4��'d-x��!D�\�um�[u@ ru"V+(e�l��H?D����?f���4`_0&E.Փ�1D�P�b��i����(�1e�FPG 0D�����!z#��@#	�?�~�a�-#D� \��O�5ز�;��G< :C��E��E�+x��U!$�t�C�	�V�l�E�4Sގ)ۧAB�P��B�I�v\�a���$f�i�e�
=_�fC䉇C�XjBK�)�^ՊW�M�2C�Ɍ �jaf&p�Nu���؂bR�B䉻!O����t�v�RH�?~��C�I�qt< ���R�:�HÌ=A6�C�I�������
QT�
��#�VC�ɝ�褺��|��IT�H_�<C�	W�l�O��!�J`��ƌ�TC�I��6mJ�@88lSS� p�:C�	._�h�� �/M��y �k]�C�	;S��JW>2���J�JAFB䉬p��<�N,��s����B�9f��l.�9%�}pd�D�b�B�	�(d�����H+b�\Ԓ��׈c<�B��?K����!�A�`�J�h��:c�|B䉯S��{A��=O2L���"cM
B�	.���"���.w~ P��(L5�B�	(+��t����8p���`B��C䉌k8z��t$��l��ɚ�J�6B B�	�cM ���ʁ73�yB��N9�C�I��r��M%+q<�P�)B���C�#����ã[�$0P���,��B���
p��*M�6�M�♊�rB�	*.��XZ�2��<cB�s�PB�I�*�8 I�gE����i����XC�I�W*�����E��I��mO��lB�ɐf[��ö���/�
;��B�8NB�	&FXyтD�/�1�QS�S�xB�I�;<r&k�������lC$ �C�I�p/� �Ĭ�7P��)h���\=�B�IfH�H�u��q3�KW3*!�DҹW�I)C˫�<6�U�!�� SQ��&k�y�$_�H���!"O�r4�,S��a��"m5$� �"OnM��"�5�{�(&*��9c"O��y$�Ɛ��A`%�^�2�(E"O��"�S�7�.| �o:�"q"O���,R0i`�!�d�7��<��"O@U	J�3���j���!�z�2`"O���I�!d��X�C������"OmЁ�Ɏ�\ Ȁ�-��M��"OD)��b<
�h��AF�.�xC�"O�93��ts�jqe9\�~���"O�=I`)��b�<2�c١��H�"O�9��N�H�t9�C�s�,@"O�LY4b'q8��-�"T;@  �"O
�@�K�*�\4�U&;C>���"O
 QU�=	�q�4�w[�.)�"O�\:VLQ�t�ĀP�Vw�I�"OxqVb�R�)��^�H�� ��"O�d�q��:[|����
�x��"O^d��FV5�j�$��h��:�"Ox��Ҫ�*Cy�i���)5jޠ�"O��E�`W���RE�`2���"O*�'�Y`�,��6E],�p;�"Ov �2�>e:>���%�~v���"O�H􁘟~i1ˠÃ����"O�U��f��d�\SG)��@��(��"O0�xW��o�FH��%��0��Y`"O��[b�Z2�|�y�O+��b"O�K榈�u*�!6O��g"O~��C�K*ƔH��D?�Z��R"O���Fכ0[bq���d�Tx1"O�!q�O-'bp����L��$"Oh ��NS.G�|�� gRC�sa"O� Q#�ӃYcZ1�e���|9�S"O�8q&�J$��,��C�Z�*Ń�"OP�#���  e�@j#i
/7���H�"O�9�'��F]��6�	a�f,)v"O`1sU��'X�~ApB��&jzj4�F"Oh ��oƻ)J�zw��8E�cD"ONd�g�S�y�8}J�Ò+r��8s�"O0ň�B��\���%x4r �%"O ���hG�L�D� ��+%n�� "O�a��ȇ�(|xr�\h�9*u"OP�b�#Ϻi���©�
j�1*ORԡ�.�|������y�����'p�$Y�/[�"1NM3J�rR|�P�'+��z���@<�"bK�`NZ�'����疙QbiT@���'o|Z4� �;�=��x��j�"O@k�#ƹuhܜ�Ca��~3"O������T�`g�78�&�k"O��;� �($HѶ��E��E�@"O�9Te�Na�e�F쇸 �h5c�"O���6�B	���ZW�J�0*�)�"Ol������T�f��N4Dm"O,�!���?b�Ehef��1�1j�"O�-�g�
4d��Q�B�$n�(�"O�y� 	�%V��(���0.�Y�"O.}���0V�-�T��#bX�"Oh�A���87��lQ���(r�0�"O:\x��	)��rR˄�|
�@4"O<�KWH�M��(s�6\gvh�"OȰ��L��0)���"Pd��c"O�����BH���3�
N_�� -D�� f�Zv�u�ڝ����K��0��"OZa��͌��<�:7o��|��I�"O��8�$Bj1�l�EP�b�d���"O>u��oɋxb�@��ҔZ��dB�"O��wI�
0�� +���=j�"O���gT?p �PQs�.*�p�"Oղ��HAt�V�F�[�$x�&"O�qa��g%��P��šp禌��"O�L�tEٮBl�\�׋Z�R��+ "Ox�����4wTdX3J����(�"O��kg+���H%��ꎲNT�{b"O��:7팴,�� �eK�!Q��I�"Odh �Ds��M+��Hb"O|��kJ�7���ܦS�`x��"O |f�.9��pVcT�i��;�"O��@�kL:0���'c@�g"O"U q#�,%x �r�P�w�`�ґ"O꡻w�ӆG��q�(Қd��M{"OČ�!�{�d��6c����?;�!�ĉ�Lf`X�J�p���a��!�q̆%p�I��?���"� [#t�!�Ă�`��e�ҟ�.l��@-mx!�dWUp٪������@?!�$�$k�d���EJ����
�u'!�D��da�M�&R$P����M!�DN�N�i���@C� ��!���!���fG6}�D�K4�Ȋ��~Ih�'��{���P�l2��Qc|�!�'��qhӁ:}ȉ!1�7;	��'�$�ʤʞ�h��x��M!Dʦ�*�'M\����v)���%E�%�	�'��:���Q����H$4;�$��'����U
6a�\&1��ɩ�'��)#�:q��)fQ�,�x��'�n}�@Y#��ʦ���P,a��'^�y[R,�����-@T��'ԚĀG	�����@� �yS�'PF;��@�嚰�Anنv��H
�'�TH�����:l��S��]"[��و	�':�4	'�[�:�j`+&m_1b9��P	�'��5�؈itY�vJ�%Cà}Y�"OF�ct"�uFZQ�V��3s��@�"O��t�N,E��rS�E+[�Y�"O�P��	w�i�0�Q����H�"O`E�2�^%K� ��zH�"O��@0�-�ТSe�#�^�#7"O�a�E�)F~�0�7�G����ʗ"O��P1k�
'j6lY��ǜ0�� ��"O����ҼZ�t�"��>F&n���"O��jՌM���Q ��l�l�"O^ps$o�3)�JBh߸O��-1�"Ox@i�NH�Q4]�r�	-d����"O@�8��+,�hQ�!�ZlP�  "O�=��	P&hr*T� B�']�Tu��"O��Ce��*at��r�׊�V�Q�"Oj=�Ќ��a�����	��^�r�"O���G^�
G1���_B��Zv��?<�-:b�H��:�9b�F�;H>��� cVH�7@� ���)ֆ�o�<9uAލ\�T$���=���F��i�<qPN�:?� ,Q��fV	��Ug�<��n�ssJ)��i9��(ϕ{�<R�^��HlZA`�9c@=� �b�<�͞�|s����RU�m���b�<�a.�&ʔ0p�I�C��k���S�<� ށ��*�=K�N@`�C���M
b"O,�t�S�s��|2��A�,�k�"O�(dł_��x;G'MTf��"OJ���6^��ؘE���9}�Q�"O��al�)4�����kFl��D"O X��O([���A�rڂ@�s"O0y�*��w)�M����xȸ!��"Ot0ر�F�"���
��U����"O6�h��^�Y-z#�ED���0�"O�5�f���?{x:U�O-��u"O�鳫C��4���6W,δx5"OZ�sm	E{�KA	ɅT*��" "Oȵ��K�W�(�	2(ZU�"O�4²Ƒ�."�C�	Z7鴴[V"O��k���V�$�G-%�z�s"O�	��D@C����q�Υ[��0g"O�$K�K/"pS����T�C"OZ5#��ܲ$�:mҷ�F�"��=:D"O(Ȣ3�Ȗ;tԈ��N߱}� �Ӵ"O����B4a������͚A���	�"O�@y�mT�b,����Oz$Z�"O��RA�	� Q���M	�Zh���f"OVY(`G
S:<���%ǱjV���3"O����F�Ĕx$fK�_����F"O���$�>pZ
E��T��t��"Oft��CΞ-,]�1��:!C*���"O`Lq���;G2�2�iH1�D��"O�a�p���^5�{�c�YbN�y�"O� *���B墍;X:H�"O)Iu�M�Ԧ b2N��q"O� j"/Ev�1p��9=�`$�g"O��bf�F�"0{���	k��Y"O����)6sȱtNWG��`j7"O�\�dD8+�4��ˋ�#*,T��"OP��F�K�.M�!	@,6���W"Ox�tB�xS�I�g��?bnH��3"OlXڶ�ѐgŪt�%�̌��mS�"O��2�,��}����JZ)�t"O�@� �x/�1��Q�&��#�B�	�V	�g�A[����h׉/�B䉳L@:�g	�Uq2�S#E;6B�	���)���"�p�[�ᕌ$B�ɰO�Z5�����<��2��p0b�-D�xh�Krϒ�Cv��E��M,D�8�:r�LEfF�l��:�7D����fF�~�أŊ�4&|�K4�3D�D����UӒM{UjAt����&D�;�W���I�O:Xͱ��&D�0+b���� �f�Tی��J%D��ɃE��)!�q���G�[n��*#D����8&�� ���mD%pD%D��C��-(aĸ�QaǄP�@��j>D�� /�#W��}��H�N�<]���<D��+g`�!�L�J��/Q�	��6D���V�@?5 ���+B>r�uP�N D��Y6�>05� ��!���Uo8D�xJ�L��mDj�td��%OdH�D<D�삁��>�j��ړz��(�/9D�LA�v.�z���<+���:��'D�����Λkid��q�у5�0u���7D��œ"jD)�)�91��X�(D�Ȱ�oS o�
�ˀOZ$3�Y
`#(D���f#HG�e��I�+�֩��7D�h0�N�B�q[0�	�6Ð�au�8D�� �Qd��c�C)��^�	�"O",����PJS.L>V�b�"O��b�/�n���:8���c "O�p9b2��ȇ.��T_4}�6"O�%�C��`�����:T�)�U"O,a�RA?)��`��#ٜ��"O��BN��t�>�1�%�0���"O�\��&|<ā���6y&�"O�2`S��4c@.S xr�X"O�ՈQ���0EDA�`��"O
,AA�����;�#�I�D��"O��+�8P��<�A�<e��m��"O0E��΍A�%���?KK����"O�й�*]�1�$�+ d��Ht�[�"O�U�KǽG��\(��^��9p�"O�i��ўElݳ��_�<��\��"O�jg��3P�\0ti�1��"O|����	3$T:@�AR�b!"O[!�l�f���
l��M�"O*4� +O��ʕʊ�
.>��"O6u�=6B���޹c��`"O��	��G�g�,���$� ��R"O���d�?��hB�f>�ͩ1"Od0��E6,Nx�tb�b)h��"ORm�R��#2`���@98!�H"ON�'N��0f��H ]�Ǩ"D��xG��@��P �m_�u7�q��'���*4*Q��ÉPf��Ta�'����)׮&��a�c���c�l���Bv�Ը�F�~��eE^�����j6Ƞ
A�I�=�� '��ʙ��S��A��ȚA�`�Ѐ��"G}d%�ȓ~���R��=n�%�
3�Ą��h��6��`z����)���̈́ȓ"�`Y�f��3�!T"A'��ĄȓQ<U�@�	�>�Pm�2��-TXF�ȓ#��G%�tt٩!�3#x��ȓ=��m0�KF� W�y�C�RdPp���t�#��ʙ?�ָz�A5��Ņ����D�M�hBD�
P��]���M�8�����G��fa�Wm݄�c��*�ˆ(x��$��@�2�!�ȓRC����L�
��A�&S�]�ȓ)���ގ$�VS�	^� ���
!�����qw�I*�Ý�M����ȓ^Y��z�Β�lx9�c�<elĆ�N��y$�ԃRg<E�e_�>u�i�ȓQ����@_�[���D�FbC>�ȓF	� �H�n!P��H ��]��T@u�P��#oD	�`,�z���ȓ6��m��ͦ~��d!�E��W�⩄ȓW9�XPf.���U��ʃ0���ȓ9��<���t
�F@��]��nP�Q�S�X��$X�SF����ȓ�ș��ԯyj���H�
1i��N�"͓��Xjl�p�$��;&��Q�ȓ3� p�;�Nc�hWX���v���e�7)�0���/M�݆ȓp�̴!��N9p���P�R}��6I�iB�B^�9��Ÿ5��
6�����	<,�PA��7z�d�����T@$Y��}���#�;f�Hȵ-�%]b��!>^`a�gĒ)��`��K�#�z���h�b$� l�j ��镺,t^���S�? � �� s��i��g[�_�E)0"O��2�o�+��Xp�ِAz��"O�܁��?<�X���W�c]����"O���dA	W��a���S�j���"O\�@g��-d_�-�de�G5|���"O��З�\o�U*�ŏ�S�ܴz�"O�x�S�	�$	.q����/$"�
5"Oܼ� 	WCj`
 K0 �w"O04��	K�N�0��˚f4+"O���&�H�w��
�Q@�"O4�r�8%+|�4�G�Xfᓑ"Op`���� �T����="bc"Ot2A [
��$YsT)B�q�"O���T��(m�
G�=S؜9�"O���Ą�B���S�#mjj "O�@ �M\�c�����Vl�A�0"O�a�Bf�AK<]B"�:7\4L8w"O�(ĖE<��Sҫ��8�.���"O�Ͳ�,�"��4�v��;���"O���q�
�r#i�Uk�s�T铦"O�1�h�J^���
\�\>pe�D"O�4��L_/���MN�t�u"O ��"�	^����X�M�(��"O�-�&�������n>ـT��"OVeJ�%��n�Xd��lU�H"$ pA"O|�{5�G�M��Ac���fE�a"O�=���$�2��D��AD@�"O���ț $��Q'@��^ ���"O�����*���2dݖ"L
��"O&��%��*h���ćWFbm�4"O��� O/>�y%�ɟ$��*�"O�Q8���3B�������J��b"O֧�i@0t[�'@,ҰI�"O�qX�*Xrv���W�+'9|]�a"Op}90a5C֚�rŃӬ!v��#"O�}�"�ώ�(8Z�B��1r�X�V"Ot�#��&��8�O�a{�U� "O �[1O+]LX�ȉ�/{!��"O�\���D����O�(,z\@y�"O�X�c� �^A��Cyb�C"O(@�i�D�����#�-kܼ��"O������W�x��ɛqeyf"O>���G�<aMf�42���"OV1Y��؀T��� D�A�$a�"O���Ŧ�v,�8�ce���A"O
�sg����a��IS�0(��"O���#��?S���)2s��KS"O��k��S�IUs�hʨU�d-��"Oy饍U;y����U�ӕp��|��"O&1�fe@�8?LY�%!,cSv]:�"Od Jt�Y�O0�k��Ǩ=jޕ��"OJ�!G,Z�SX�
2ȗ�1��"Ob`���y���"��*��:�"O*����������هD���"O괻q�L�Q�M!�Ѥu�L�"O\��W�6�༡�eZ6���8"O��3�͐�Yo^�c �,ծ��%"O�M�D��w��9�4�,+�9ؕ"Oj��ac��MA`Hu#HY���"O���2��;��ل�a�y��"O�y��>F�zE��'�%CFz��"�Ě1}`mW��p�p1��/����'�Z|C"¸6TV����.�(��',zmx�	��Si|m�󄚏x28tR�'�+G�i�y�w%3��Y�8D�� �\��h�3��eFḚhӢ�i!"O�q�B�O�7��� ��1���0"O�uqq�Js���T��Eł�R"O�A����rOZl8GJ�)�jp�"O�yѶgP�S4���
ɝI�|(R1"O��Q�L -��q+%kQ<;/��7"OF!3�!�:��2j�:�C�"O u�pj\�Ct�k�J�8]�4�"O��� �D.E;F=i"L/;>�X��"OZ�"��J]�2��e��"OV�*A+^�_p:��ǩD!$�m)�"O��a��� /�Qza�ߕ
�8�̓rРh�p�K�Wt遵��Nz�͆�U�$�hT�� Ia.�I ��ɆȓetX)P�Ғwը��WF�Z����ȓyqԠzu� �<^���C� >Z��ȓr��T��'��+�*Mq�̕A$��ȓ*o�����r&|�`MD�8~�0��dy0���@�S݂9CF'�A���ȓ�
ak�kߤ�ȱ��H��Gu �ȓ7䈽jT�ف9Ł��-7��t�ȓ`�.d���^�rz��Jt�][�l���� ��#ت�5�*tִ���(���"�#)������Ȟ����:}��6O�)t0��A,N�u�Յ�Z�*SwY�&��Əǲtj �ȓ7�ԡQ'	�B�pP1$�&z����w�z��IբP�be g(�mtlC�ɂ]�.Q��N�>K�����7 ��B��,e=�u�R�]�:�й� �"TRvC�ɩ&�P��B�rEj��B	1�pC�I�Bi ���T���V�8C�w�bpt��e�BU�8IG�C�I�5� ;E�ь:��mRDO��DmC�I3:���x��͒�va��,�/n�0B�ɋa��y'��&� �i3�
�9c�C�IN�tUk��>����qǺ��B�	���� Τ��Y�tm)�<B�I�eX�Aj�@�)�k�-#�0B�I8>��T���=��J�m^� �jC�Xlj+	�6��Q,G�DC�@��1�OY9@ђ��j�r�C�I�`�P�DgQ�O���pG"�1��B�I�&��`��aL�Q���B��;&�B�IJ;с�@}~�)�(���B�I(]9���č���DG�]��B�x<v4x����jҊ��Ƣܵc�LC䉗X�R�"O?�L1X�왚�.C�	 H�q��&� �hSL�:^C� `�&a�% ¼K�P��A�FB�+�pzfC�g��$���T!0B䉯lM���G*�g�VDJ:��C�ɒ3����F-X�k��#�iS��G"Of�S��_]G`@�{&8�
"OZ C�"�$[�����LT#[��"O������3S�02�i��5-�e"O�y��l!9b�$�W��<$=��"O�x���Ģ)1h�a�N�~�B"O(mȷ��L0 @��F�0c��tK#"O�1���48h��3�K� �i�A"OPL�%��L쩐J���H��"O �+Q����z��9�(p5"Ox�a�]��U�w�ŷm�ŋ�"O�DIu-V�&Mj�`�%%���)"O� @���D�T�X�sM��h�j	(T"O`��f���8�M �h�&L��"Oց0��S�kƭ�񋚺'�b0Z6"O�����
a  �M��$��"O� cI����i�ҎD,q�F��"OL ��e>C�D�{S ��%�%"O�4 �,¹~w��@v�͜tL͘S"Ob�)�Z�(B&8ŝ�:0 "O���KT��Qk���+�� �"O�E���h����O!T��M�0"O�]{'%C�w�R�T+g�lMS�"O��H&A��8Iؒ�U�b���E"OthB�D�+2��@��&R�a��F"Ox� T�k~ܣ��m�R�B�"O�x3$�<'�h�Zsŋh^��"O���%��)<����'*g�y��"O`���R�c<��˷�XZ��m;"O��c6�@?J���4kKz�{ "O�� U�]�5�<��a�;Ht�s�"O����>-qx� Ǎ]��8�v"O�r�o�;wIN��f���6"O���D�D3 �܂#�T>7�l�ٷ"Oq����7�� �֬�(2�J���"OrX�I5�`ڔ!	��X�"O���2AV�};�=qc'��
H<�zu"O��0'�ح��l��Y�DL���"O.	92dۡ���x�$��{�]p�"OXmp��˚=�V�sBM�gJ�ذ"OV0�c)�?o؍�U�qd>�*"O�Z#��+��H���U5%F �v"O���j�4��͚rl�UL `�r"O�1�$h�J�N00�i�0BXT�(V"O@d�4hT<r��`	Th�*@�Q�"O�X�qa�,޺�D�"��R�"O��Q�d�u����0�N�p7"O  �&��x����3��
X�M)�"O`��&�۰|
և��Pe <Ra"O��;G�ь,�[Ռ�5��Q�"OdUc��^�.�:F��>ݚ$�c"OH6��b�����,�X���"O �{c(H����!N��$��x�u"O������vP�qq4�Sk���#�"O��@!���6V(q20�Z%P��9"O�BwC�Zafٙ�p�X�"OJ�J  i+�8a�q� :U �*�"O����j�y� �qOTn�]"O@h®�4�!-�f���/�9S�!�d�i�[�0�L��NHw�!��92�3PBL�
E`U[��F#9�!�_ Ft�wB�3{�|h@��`|BO|�g��"� ����-��+�"O���%�i�tP�wo
�z�0��"O:���i��@��8n��L���!"O�$ըR�7+����Ύ�1�!���X3F��%�!>����)a!�Ȓq�vH���Қ}��-�Wb�.�!�ğ2P���w�N�x̺�e�!���_��$3�+��S�)3S��2!�� 7Z�Q��M'W�v�`�_�2"!�V:2/~�A�&ƛ6�ti��O!�?dxb��H2/�hq���I��!�dN�X�F��V���\�P�O�Z�!�����37ܺ����!-r!�ӢA��iq�H*�6�8&F�]!�� �i����/^���êFhS�ȓ"O�1��8&�}��n<s��0�"O]K���Z~|ipm
5MN~�9"O��'΂�^3�qط��)[dY��"O��`WL͌'�� ���t(�(3�"O�� ,M�|���cɇ��6"O����?Q� ���.s��S�"OBs���p�e�Vkr�DX�f"O^��w��#*�8q�B�P̠�Sb"ON�����,���Bt��#��-�y"+[,H���ȱ$[�G���`/K�yҩ<O׺lZ󋉫h��u#����y��S�_��xjtM8� ����F/�yb'�4z������#(�,5���P��yR,	j
�%a�"%$A\��� ��yb���oi�Z�ˆ�G�Zݠ��yꇱ@bZY2�#�3]t� �Z�yB뛴(Y>i���:2E6���.��y*�b&��F�TKlI�n���y"�ċJ[&A�d@A�x���	�	ܟ�yr�,7�v�
#gƟo�lRvFF��y�mכO�x0�3'I�1cB!�E�F#�y�j������M"r���<�y�i�.|+#A�V�m䊅`�,��yB%��>�4p�,՝c�Uɂ��3�y"/�	Gh����4�#�K���y"�%��|)�vJ���+^#�yB��Y~B(;�".=7�4���3�y2�ߐD`���H�9�*�-��y"�ÿf��E�+h>��"#!� �yB�P6i̺Ӄh�<W�p� ���yb!Sh�5�fF�0K܀�s�@���yrNU�d0�erb�=q�E�A␅�y���Y�PÔ�X!:��y��j��y�G(4{n��Do�#���A�M
��yBa��8<�*%A�������yb�HYn��섃bq����
��y"���K���&Y*�Y��lȅ�y��ڋ;�*��EK�O>���C��y$����{G��I 6������yR���~!!A@
?��8����yr"�'VX�h��2` X�G���y�!�#E ��ޫ9	q�фN�yBE�0ER� E-�,���i-�y�_9b�����7�B�(a��$�y�=����\�l�f=���2�y""[7ip0c��a� �ё�F�yrO��'4�-�ͅ3Q�8Xr��T��yr��	��&E��R[*3��@>�y��ߵ8�ڜ�S��3Q��x�A�8�y"�]�
#��f%�-y��m���y�Õ��"S�� �Ta�鍕�y��ҌVC����'�<�8��e��yf�LH�X*'bO@/�9J�-\��y2
�e�.��@���k�zrBƏ�y����.����֯0`����yBAVQ@<��[�Z���֥��y�	g1�Dr�� gY���(�8�y��:]��lX'�M�b���{���3�yRe�eޮTrDU'�b	������yr��_cȐK�E 
YP��ץ��y�/\4������~΢������yb�D�j:��7�Ίm6԰`F���yf#f ��ږL_��䫤�D�y
� �1 �l�p�'ʧ#4$q�"O���cӃ�6�����)�4��"Opp�Uς�O�FDS�яO�(�"O�D��.v$�UK�� (0�"Tyb"OJ�`�W�$��н�v�"Oa����3]�1rV��$�V��"O�(s�ǋ9hH��	8x,�<�"O�(��V�L�v���2b�E)�"Oj=@�H@�D>�x�� �J��xb"O�\��I��-/j���*ӕCJ�Ru"O`PiUZj�	 ��-<�l�0"O��a��K���c"��Z���f"O`�3���#1��C�͍�x�"T"O�Ac��+�4L��N���UR�"OD�3jWqy
]0 RS�Fqm&D��e�U�a�(���j�~q��8D�4��ۛS��x,M�,p�q�))D�+��ȘhR�����8s�2Mҳ�)D�h��eW:9�^hz1�N;�*I�F-D���R��W�h����%Mܰ��#�*D���祆����RWd�_d�!��#D��J�n��&0�t��/%�v�AI/D�<��� W!~�6(̓I�����,D� h���f���R��"Z��,3І)D��yf�\.*t������	�*drs#*D���E�#�*eht�Q20$(c'D���&D@İ(q&δ��05*O�a+wK�.2ذ�0�/	:�x�@"O��c��ĊbE^tp$lF�9�t04"O�0�Ağ�6�6Y�ӿ\��d"O��s�o�/2�<���#��B��4�!���s[�X���ݐkW\4pi�3�!�$��[r~EbG۳MQ�9*W.��%m!�dōp�@��y=�p�P��	!�$�����'�
6����>_!���q��F �$��B4�!򄖽X�$,��W�<�����*�y�!�$M0����Ŧ/��(JQ(Y��!��
�f��OӐ0vJA�A"G�H!��G�;����$�"Xb��bW�6!�Z3z��*��!1��1"Z�zD!�Dك��R����E> l �����!�$ )�@���nwl=�)\��!�$�T�उwɗ#>.��Eϔya!�$�5|Q�0�$s,JےZ�=c!�Ğ8�Z$�V�۸#P|��֘R!�d̿8ϐH�B'ŝyz�H�q2!�$ۢr��c�,����M��!�Q�DĤ�j�-�l�j���J�@�!�_&%�-����g�0)r��<9!�$ߑI�ik�H}��Yj�I�!� W���sEĆ�B������("!��> ݻ�B֫O����'K6JF!�ą�H�D��J3a��1Ȳ�K;p6!�DX��������e��Ǔ� !��-���ڒG�ֱAf�Z9i!򤊃�t�0��LD��|sC�&M�!��)7���ej�i�B��p�O�Py��w�T��# 17zD�P��Y��y���^Ol]��nF�#2�TҔ��y��@�fF�0@���lv��S�D[��y��F�,��x��G��K���P�B��'�>maTR�V�(B���3��B�	�`��Ŋ6� �SN65bP.�,
�4C�)�  ����.:�Z�& g�"���"O�98b�LXD\�Ԣ��B�@��"O���sÁ1-�Tx��L<ai���"O$�Ig�G2�����'p,b�"Or���"a
$r`@�p(�;�"O�B����p�K��&4C$���"OL8H�]%1��	���7)$4l)�"O�h�6j�(����(��&��V"O^����=��4�bgK�"O��6O�7U�1Xc$I%f��$ �"O<X�+��Ŝ�	SJѫ1�b|�"Oܽ�e��/4�H �9N���q"Od4
s �g�Tz�HO�	jl��"OlH�P��QZ��I��U2�����"O�C�y�J���K�ka��)�"OnRC'�0���z6 ��uN d;�"O@Ek�ʏV��=ځ΀#�%%�ybi
�)�F(����^� A���y�V	[�Dx&IA�X�0�Kaܑ�y«�	��	yc͹O�1�P��yrmM���1He-�p���2'��y�m&R�|�h��ATʍ�k�y�
T�e�P����Q������yr
� �X<�lF$�����F?�y2��g���!O�vV|�ɢ���y�8Y��X`��Zm�hP����y��6.^����@;L\�����y"�N�[D8������J�n!�"����y҄A�Z >��bDo��r���y�b���b���)^�:X��#�)ح�yb�Mv��aW;+��Eq���y!�1�H���a��V��C$��y�.��i;����O
%��tRCV��yB�\�2{v�vh��lV�+C���y2#�@�=��΀bAD(D�"�y���!*�xP�s��8`�fa�s�
��y���	���[�ݴ]B-y�ŝ��ydE<#�8!NWjD��u��'�yri�	Y��S%+�0d��)i�D5�yb���(`	��d���S ��y��K�BPȌ��F��f�(�!��ޤ�y�W�1f��KF�F����"«�y�O�f�������dy8��H��y�
ؿ RH�×n�Z�n<*�ˊ"�y�E�+��h"��{�61�#+���y"IɇW���z��z��ܳ6b-�y�
��mav�A"n�>�8&�	�yG�#���X���^����E����y�&	5<M kr��Tr�]p���y�#ڽ]���eo��yׇ�\�<��oL���U����7[&D�e��]�<q���X5�E:�"�y�>P��f�d�<A�e	7b���E F	*�(�C��\�<I%�H�
t:H��F��+���� �Q�<��kڞ3��u C�5�ŒTLJ�<�gS�JSB�Х0��
�B�<���Ճ7����m�>;�2��P.�{�<Q�"@3QX!�����)՞�q�C�p�<�֦Տ�ؔ���	�zB1�5Sk�<��d׊e�6\�bM�oc���Uf�<i��L-����t$�n�\EyVF�_�<�wa;|{���P.J��Q��UX�<Q���ݪt��/�K ��s1+J�<QOQ"}���S#U\��D'I�<� J�
!��)���sGC�$M�ذ3T"OR����)PI�ai��D#C�F���"O��1m�7t�01;f�Qը� �"O� r�d��0�c�CJ��r���"O���A��-��jvd�H����"OF����&Y[�u�e�O�s�*��r"O��{���Y~Et�N����"Obq��ĔnZ�[�ϑ00:E��"O�����C�~�P<���H �$��"O^ؚ1ϝ3U,����{ bHf"O�⑆�	����c��B�ؚD6!��Y�on Ad�\9�����#�6�!� �/Ծ����<;J����[OL!�䝍(!���	C�t�"�H�\G�!��y��\�T&̮0f�pʐr�!�d�($ZAH YS��(	��e}!�ĉ�"~�xPL��&�ɰ�ӟ	�!�&7�6�!2���D�z�tNR�$�!��ԨH��E:�N�7{d��,��!�D�g�ĵn�%a�����	�!�! �V- ��(��}��͕�!�D��u��Ѐ5��b��m8���!�ė1Z�b% CY0���@���:s!���B�b�2��z�:T��v�!�� vz(r��mv���DKp!�VY���X� �9)�)A4�H�K`!�$��|�`��EJ���$�!�I,%L!�D�Hξ '�T�D�V���C%!�$�|#ЄSg�̾ay�q���'5!�� <9%���`.9>\��G�Ѡ"!��(q/2�)򎅘vP���s� 
!�ǈ:*����D�4��)����!��Sߺ�YU��D�P��wE��P�!�$�����Kcc���,SV�ar!�$	�}��lXD$Ɵ|�6(d�
2X!��צ$.�YSp`�9S�ک[aϑ�}T!�䙺iWd����E�� S1E٬S!�S&J���&	�MrP ��e��"O�a��L1=���GF��(;�`��*O�9��MQ�
Oj�r&AMw�h8�'B�9P୘�P���� ?Eb���'���r��̧m��d�)I�7��0�'���I��
�tkpT�1�4-�Ό:�'��а#&N��ٛ�N��8�'�0��ԮN�MWP(r��О����'פ�H�\�<��r� ].-�
�'�D�XwC K���!�᜴��X
�'jZ4�1� ��aQN���>��	�'B��r�mP4c6�aeBù(e�'*�P�U����ǞI���9�'�x��e��'MҾ����<ȅi
�'a����ϛ�` ����)/\��'�F�����'�`xC��Z ,���'��X Ś�6��p���C'Rq*�'��L�w��,`��.5��̚�'m��Г�#^�� �.�R��	�'����+Ē]3�#�c8�X�0�'˨���Å�R@�B�:��p��q�<1E
$�8�(ЩU�z�![���q�<q��
n0���aY#`ܪQV�<���G=+j�1�) gj2��rj�T�<�V��?��A��Sg�y�]N�<iA��>"������N�p�)G�<q6�1Q`��`�J��҄H�W�<� p��t"�'R����C|x��d"O&D��HW�}��!��ms*��T"O��ط���J��R�o4vgXc�"O"-&e���M�@�6�lZW"O�%�A@���k1�� /�=�D�I��؃i��*�6�	�:e$��M�U�>݀��(C�qOl�$�ho2)�#I�|h� s�N�'6����O�����w'��r��k�D�����&z6E�hȻ*���p4FB�U"�}Ҥ@����=p�Ǝ#o�[V�X�E�����3���{a���O8��7\�Fde�k��?����������w�ڟ"~��k�<#펟>z8�醈rX���$�٦e�	���ӰO*�[�g�ds:$a�&��4�W
U��M{���?y)��T
d�O��DoӒ 3G$�4�,�`�l�2.I�R%�!@)O;@-���ݱ �z�J�ҟ˧��^c]�A�?Nn�}caǔ8��޴"Q������"]M4HsacɚH�\�y�D�G�<�|�1U`�0�'eT,#��4 � 5�8)o�g����O���?AE��&~�	t�S25�F 1��  �\��㟔����܁A�B�X��p�,%V"��&�b̓)�6�'2�7M�!l|��qɛ���<�N�fS�|Q����MS˓`��A��O&[J�� �1r'^`�u�R�3�n]���_�
�ґ�%�H�`���[~�'���IƇD�lu�*����}����`���V�8�3K4�ٶlE��i�J�[�� }Zȵ��K�2Huc��J�9�fh��O�I���'S�|��'Zb^���4M�(m*D��"�!C�a������L�Mɇj�3��`Y��]�t*rY�i��'O������'5�S+m��l�nߺt3$�C���`Ęa��L�'����	��<�	�4�ԟ����O��	��ݲ��� ��|a���%�١j���rfCM�"��`F_�L�ۍ���,�\A&Ć>^�*,��*��r�x�M:��}pF��*��,Qc�%���9`�	�2P��a�T�'�D�P�Z��D�^'WY2��A@���M����D��˓����|�ɭA�Vlj�O�Q��\����}�<�!%Ǎ?!�){���$I�8e�ck�%P�x�v�$�O̰mځ[��`޴�?a���?�]f&��
��A��Xy�)� 嬡z� �D�O�d��pIB)�dퟻ[t�=[�#�xT�Xs�O'���!���XL�� �H� }��k���+�p!�N����wB%r�T�: �<c����9
�F�2�՞zY�����I�2�d�OB�$>9l��)��-	�뉫�
��q)J�QR2����������\�,�Z\ ���-�D��1�"Ọ=�|�°iy�,r�L����$ez�GŻ!WV��>�=��O��$�|6�� �?)��M3�SfGr� ��w�| B�P+ntV��&��_ Д�Ĥͪ$���ן˧�b]cLf Z���92�,tB�����F݊۴oc�D��}��y��ڠf~A�M�Kd���|��[�"���2
`�B�� π�m$Q�����O��i�R�sӠI�P#U�#+��ag�"r�|�S%�O���<�O>���Ԉ�
S��a���;+�
^A����Q��B�4�?q��i��Sͺ��ꏇ29
-IR.SX����$H��`'��퉍wBf p   ��   �  <  |  s  �)  5  H@  K  �V  �a  Dm  =v  �}  `�  ��  �  5�  y�  ��  �  H�  ��  ��  P�  ��  '�  ��  �  Z�  ��  ��  ��  R�  � � � A �% - �3 $: g@ uD  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�Y�G{���˾R5$�Qb+�jBƅ�7��Oi!���l8��Ӄ]*W>�\����]O!�ė��ތ F�8#"J��7Lb!���P~��#���(%l�(.ԜoI!�d�0c>��=`�r$,�
�!��LP!���6HٮsX~��!ݺ�!�Ĕ�m��G꟯i�̥sQ �W�!򤃛]Q���D�o��Z`A03�!��R�6j�l��B�^ ū@��;Ol!�P9��$`b��e&Ī���c@!򄊡jX�QTυ#i��A(PhˢF"!�D/2��`pB�]�6�`�6��9!�dEE����BݙB~�tK�`I�W�!�DV�=�i�H�!(^n8�䏔$g�!�$��mMX���9OT���n��O�!���-
l��WoР>J���NE�ni!��K�4�VYP�ɑ����+L�xT!�$�4<{��J��! �PhX6*ʨI�!�Ff^��PR*C�lʹ����F!�ͪ&�����'�4j�\���(�8\!��/�:��������bN	i!�$�<PⱫ��53���{J!��@�S�vL���?ʀ4sW��*t!�DT��`Iȧf yƬ`�c�]�#�!�D�p�,l G�.x��ᲆ�T<@Q!�@7_�����=�"|p0��-N!�"F^�cbI��i��,�g�:'�!�0�@1g�żm]�,�Ҭ�
3�!�d����(�qKrأR+�<q�!�ںO`�i�눏`�p�5mܒ<�!�d?B�>�1f��~�>�#���0b)!�$C6h���@焐K�и��)4!�� 4IAI�R@`�g� @K�C'"O�ِ��3|�V9Y%hS?<v��"O�y���<9�t��'��X=�"O�a��Q�/k ����$�Lu��"O08DF��D��6.M02㼠���5D��")U+e$l�ȶcX�6���Hu*8D�T�N�,N�n��4h>~��ǈ+D��@� Aƒ���eT�VD4��%D���q'�
1��Z&�Q�9h� 6D� ��a��1k��T% ���J)D��(�f�4��US L��1�z]���4D�p�3ϐ�ѡ��R/BI���&2D��I��.��s���p�� -Y����@�Ta��ցE��1 �oÓ�y��SZh&/\�SIRݲ2��y���(@��Sʀ�9̸3�j#�yB�ZM�z��?~�t�>�y�NÙ[8,�kWG!hQ�\�C��+�y��/����C�úkl�Y�-�yҎE G���롃�f�P}��eɱ�yBbӣ6OI��G�s�@�a�NI�y���(�=�"#�1lu�l�7' �y���8l<v1C�G͌eI^yD犠�yHг w�Ժ�=S]��������y�c�'�8*QE�K߾ț ���y�]*�������9,�ٸ o�#�y��M�j��D�2|¤{�G��y"#̽���h�A�a�Z��1Ů�y�)�s�0	���\Z�����yr�	z�H���+1��	Pj�3�y��XZXt�-�%`��ʤ`%�yR�IJ�P�����XWI /�y2���U?E���Ԍ|�j�!���y�c'�V��p�P��Bh7�J�y�:v% �𥑮r?l�i��y���T[�)Qg��}�`P1���%�yR���.���8�C["#�v��AOV��yBn�b=�A�X<� ����M�y�eD�_"J���t2a�5�̂�y�*��X`Ht���:�xED���y���1�J�Bc�"��,zu"OH5�5����\�B�ʄA��=��"O| [A�Ȯg��c/,�,��"OBy�hP3&>(��AI*�H�s"O��Ru���d�B�@(�&���"O�j�"�	�S �W�0�P"O������n[�}���>K�Ь�G"O���#��q�)ڒ@#Gt���"O��S��CT'��kR�Q�11��)@"O60�«�j_���hٶ4#�"O|P�d�I�j@@�2���4�,"O�@S��W���@�����TwB�(C"O��C�C׫Ix�Qi2���H�X�6"O�ɱ�dZ�{��ͫ�/��	l����"OY�!/\  ZR��BHW)+pD�ٗ"O�q�@C�lx�#cgިk���P�"O�lK�&T<T�����o�t�2�� "O|iA�,���٧��#&�YzU"O\ȲX*��9[V�C��|@r"O�-�Q�j ��	���`V�lA"Ox�ۡ,�:m�d��qJ�i��h"OD8bC ��\��c'/0f���)V"O� �/<]���z���F:z!�E"O^���'�����+�"ԋ$(�S"O� �x{U�jHXAY�̓v�x2�"Oࡓ�O�B"؈ �Z�6�1�"O�Y$�ِ$���RS���>-vd��"O�����?Kr�HA���X�=��"O4A$!8<���M��L�`��'z��'��'7��'��'��'tj�1���<w���G�B���'\��'cr�'?��'a��'"�'R.@q��y�|$�QՁx�ځ g�'��'~��'��'�2�'���'6�0�M��
���U��1�� p�'�r�'n��'R�'2�'���'�Dq���+K>��`�3������ş�������џp��ݟ�����4qlڌ^Q�<��W P�t�ǂ������ԟ(�	���Iʟd����\�I������Ԫ�^�h�c�I���3��P�	�����ޟ<�I�,�I̟����h�7ɘ�!���4&��W�����JΟ$�	ڟ������	��	�$��̟{�f\�`��<h�c�� �x|��iP�������$��ƟX��ٟ��	џT�����I�Ε�!�����P��
V����D��ޟ����@�	���Iʟ��I��|�&��D�d�r���>�D�$������ ���0����d�Iß��I��$��6&��,H��[�e�6!W/_���ş��	џ��	�t��ȟ,���,۲�%M	����[�ТZ��Y�������h������	����7�M;��?Y�R��"��8a �i`��0k�	۟8�����
殮!KE����1@�x�Lj��@i�V�6��4��$�O�T�'�A�N���k��1Bj�O4�DZ~�,7�"?��O���i#��fZ�P��|�a,�!W4�}�'+ϝ��'52[� F��$�p=�j�C��L �S'�܉utj7�c�1O��?�#����/��AH �ʒ�
b��h3�k���?��yX�b>%�#E����%*�1�%��:s2� r�� ����y"�OR� ��4���d�2��1q���P	��TÄ�4c�D�<aL>�ҵi�� C�y��
�iܸ	�c#M
���@�#]�O*�'�b�'�d�>Q��^nX�3��E>�`%�B l~��'�@�g�B�ژO�B�	�Z���W�j�v�0��?Ѹl�թ�J<�	Xy������N�tµ$м²u*��2-'�L�E`e8?I1�ia�O��zϠ�٣`��_��A�N��"t��O����O�ԘD�lӔ��������ݺ ����diF�B�d;F_zf"�O���|z��?����?���(�����{��\�$FϏn.�	�+O�o-;|x�	ޟ��	�ޟ��� �/l��1	QAUF�P��̑�����O���3���MT����!����h���B�Y�"qmx���A:��tL���'�x�'�Z�9��@�Y�1���JWl�S6�'���'��t[���ش"0-k�f�����>(L���A�6PP��U�f��VD}��'-B�'��롮ֆ2�Y�r��8d6����4ț&�����(!y�Q>%�蒷�&mp���e$Ν"��:�:ON���O|��O����O`�?�3Aʻe��Y��=̼Ȫ��@y"�'%�6M������O� nZH�+(���c�/- ���oK#��%� �I���S�E(�}nZ~�
,7��[��O�N�ֹ����=%`,�#���|褚|2R��ɟ��	ǟ4��
K:u�P��C���wC�t2�N��X�I_yr�m�J����O����O<�'�~��gbڻn��p��:���'�&��?�����S�T!́yB���D�P(��|9�S)!¤�G�M�V��擖;k��?���a&~�R$NX�lG>8�DcʘB=����O����O���i�<��i��d�Vɘ�l:���C����є	O-k���'*6�1����$�O���	0���R�>q7�(zr��OP����1Pt7M&?IA��9���>�3�j4V�7�(d�4�JG;��my��'��'���'f�V>�q⦉j�Х�r��([���UnD�M3 �W��?1���?�K~:����wi��qC�OK���"�lK��'T��|��4�U2ۛ�:O�8�� �N-�X�6�̌.��:�9O}a����?���/�Ĭ<�'�?Yv���*�PFF��) ��R+�?i���?������F�-��N̟�I��l�$&�]�,YR��
�^ӴժCdHW�Tv�	͟X�	d�n���qF#��H"Z�`���sx����-ʆ�M�}R�M�����+�palQ#M4R��p�L��>h�I���I͟���L�Od���>X����W�ASԼ�����|`�l��5�t*�O:�$NǦ9�?ͻe�0�q� �\�Y�G ]�G����?���?!ìʸ�M��O�@�c�6����Tt
h���,��$i1��.3��'��I��P�IğX��ܟ$�	1\�8-�1j�$6d%��)���'F�6�-_	����O���.���O>���o])�li����&��ON}��'|��|��$L�J�~�1���YO����%��_��!���i���| ~i2��OڒO8�H�*Lp�m���zɣA!ܣ
�B���?����?���|�.O�����X�&�$_3���K� U�A�-W��$��I�?!�_��I����8V|$��I�$�ܡIW!�n��Ť���5�'cl�ծ�?��}2�{�? 00��$o
�Y��G'S��)�:O����OB���O
���O0�?��̏]��T"\�^p�A������I؟Ȋܴ0�}Χ�?�ӹi��'L���''�68B�h��+>8^�B�|��'X�O̶(�2�i(�i���g1+\Q���Ǆ݁ޖAd���h��'B�	�����ڟ���� ��e"�� \ �+�Bʼu�,�	韨�'Ɏ7��S�@��?�/��!���%#�ڰ�u	V�hLZp22���y�OZ�D)�)���^)'�[�ݘ[ͶA�c��*:���J�@ԙ�/O�(�?yg�6��7}y����Hi,�Z��T�,����O��$�O4��ɧ<�&�i��2G$ĕ|kh���-�C�>�oB�s@��'�7�2�������O�YA$k_\N�`�*}i�d��O��Į��7�-?�;r\f�)�'��_�����4`r�o$7���Rgp�ܗ'���'J��'���'	��R�~e�]D>�dK����*	�+u�� �I��%?��$�M�;�����d�}��D1:�(����?	N>�|J���+�M�';Z� �3LMC�A<l:Q;�'��y:��t?H>�(O�)�O"�����G�6��-�M�bH�Q�O��D�Ov��<��i�:�ˆ�'
B�'<�q�eE��͂F��lu������|}b�'|��[K*�$퀈Y�v�jfT���d��p��1�ɨM�1�b����H���%\`a���^������z��O@�d�OB�$�'�?��L�6�����%~T9�!Z�?�r�i9l��R��{�4���yg�]���Ź�K�5FC�l��eȌ�y��'���'Y�M!e�i6���1�|Mr�O7f�U��6
Б� �<J��
L�Iqy�OV��'�"�' Bm
 a�F	��,A
(�٫� =��ɼ�M�a��?����?yN~ΓG��)�qAރ����"��P�e��Z�|��̟�&�b>)8&��;�Ȑ�U�5���CP=A+��nZ��$8��z�'��'��	23�f�`�B]���Z�Ɏ�!d�Y�	ޟ��I��i>Ŕ'����=t��
�/R�9�u �
:����GW�q�2�{�
�x�O4���O@�D[�_0��C�`,[��؛57.D�uFe���bo�ܨ�����>}�ݭ��!��\�`�챳/��p�Ih�	ӟ��	��X��|�'65�}0�@� !���M�غ�J���?1��7�f�<�b+On�l�Z�;��aKW�
�4����烖)�lq$����Ɵ��oZ~��N�wl�r�ٖ"���xw�71/ڸX�G�p?�O>�+O����O��d�O܁��e�%1讠#!��+`W��T��O ���<��i����B�'�'b��P�t<{'�*^�
DJ3���[�Iӟ��Is�)B$�'cլ��U'ɦQ/JI�PgK2E"yꒉW�Gu�xZ/O�iɦ�?I�I4�
.SƜ��,�.e$$����8t_����O�d�O���I�<QC�ie��� \�:t�,�zs��� ���';b$n���l��O�d�
j���f�^9^��ز��_Hv���O<����lӜ�;`
G.����d���Jb���
 4���'��I����	ʟL��ϟ��	Z�t��,tsF�I .��\���26*�=H=�7mCu����O^� ��/�M�;L�;�B�1�ƭb�%	�H�R���?	K>�|jw�
)�M{�'r��T��?"(��;�)�'䊠x��s?9M>Y)OL���O�m�婍�<Xb��A�Ԙ�+��O��d�Oj���<ac�i�
�c�'���'��]K�b�.%����S-�[�p�J��D�N}��'�ҝ|bjM# �RQ���.�2���J������9 ]$Y�	s�pc>@��ON�$�1���ャJ���7Ȅ��b���O~�D�O��5ڧ�?IՃ�.J �`ƨыfA���3��?c�id�up�\����4���yG���NA�Tju������!�y�'�B�'ꂔ�Ƶi��I1p��H� �OP:��Я�J@����ŁXF��i7��h��Ky�O&Z�M����?��2������5uĹ�㍑�B	.()O�dmڼf���	ɟ��IZ�ɟ�D -T��3�g��qWS���d�O��*��i�{���Q�nJf� qp	\Y�����x���p8�*'̾�H%���'�(賷#E6��J� ]K$�B <�"�'���'��O%�1�Mbm@�?��̆x�8�@�.VMn|�qgʜ�<7�iJ�O��'���'\�Ӄ'K4գFظ���:C`��6�0�i��I�qJh�ПR���n'�,ٱ�&c��H
�f�/k���O���Oh���O ��:�O��qC��	;-�U[�G�!x���	ڟ��	��M;�L5��dGݦ�'����d�JP8!�������se�JO�	���i>ywa�ܦ��'>�=��hX�.@��9g EV��j',Q/S����������Ot�$�O~��=)v�ʵIŇ�Z�Ȇ�@����O�����!����' �S>i)�`�<'G�����1A@���;?�2W����Ο�'��'[��!�j��0��D���D<�E�5! �H�
-�"+��4����5T>�Ot誐���U�0��#A�0�`ub,�O��d�O��d�O1�z� ��fo,8��L��%��t!��d�zЊ��'Ol�v�t�O������J�G�5`�@�HN����$�O����Cz��Ӻ���V���H�<� ���YT��xÀc�zPI9O�˓�?���?9���?����ɍ-"nά1�R!x�aI�7-�hn�T��@������Z������;V��\Kj�Z`c�o6F�I��	��?�����S�'�ܴ�y2D-Bf�T���H$�b�a�_��yrM%iʈT�����d�O���[<M��p��LȞn�B��o�=+�2�D�O���Op�4p���D�b��'�RM'fd+&c�
X�m:�B+Y��Oj��'�"�'�'!�K�lr<�"��G�Z��c�Oz<�D��b���#��^��?q��O���
�������%��I�@�O���O.�D�Op�}���e��Y��ec��isVMK3}��4;�3s�f#��m���'�r7�-�i޽�
�?Ed�����D�y�-r�x��֟�I� �:�nZQ~R��j\y��T��!��&z��Yr��$��J>!*O����O����O8���O��ؠhG.5��3��Ol���� �<�i�ljC�'�b�'��O���>q`�z��?J��8��{&���?����S�'8Ո@� ��>J��Qg��nٸ݀�EF�`�m�)O�e3t�P��?���/���<���N�|TX|���^4d�>��F��?y��?9���?�'���-��͟� �*Y>H��T��Ok ���bvs��de;��O���'��U��C��J8|L�<�p�҈r
e��cӏ$֞�nZV~��ӃM�T��S.G�O�����u��"X�"�E�f��D��?����?����?����O���&/ʪ9����CJ1>Q&�*�'��'�6���ad�˓s���|rh�C����ψ�YLH-���D(��'����b����f��ZW��)JNBm�A��I���ͣt}4����O�OP��|����?q��R�x�*p�ż-�>��3ϝ�
V��8���?�(O^�mڳXPr��Ɵ���D�$�W6s�\�sh�'����,G
��DX}��'Br�|ʟ�y2F׸]�0��p�`��x�D��0c��{�d��|���X'�$���{��hŀҨ��$�d����Iǟt�	ӟb>y�'��7- QA�1��G���lP	���5F�!$�O����զ��?�AU�$�	�l��I�$OPL� ���G�B:.@��՟c��L����'TrD�$T�?���|��6L
'qf����JDL�v��"7O�ʓ�?����?���?!���IJ�z�ܜ��d���䱐־)aЄl�+��`�	����IV��������K��N�������^�J���?i���S�'x��z޴�y���+^�$��gU�0~��1T逶�y��	NuT���䓸�4� �DU+xDhd�R*�&R]��TaП 9����O.���O��"��v�(.�b�'���d�Ę�g�͌8?x�	ce��g��O���'tb�'=�'ː�8DB�p���Q�����O��(!�DbX����k0�IƘ�?��K�O�[��� �{��M0n��c'I�Oj�$�O����OT�}J�a��|��3
F��ϑ;1n�aJ��Û�m��b��'� 7m#�iޡ�Ŏ�z}pp��!&����e���wy�n��&��6��������;� ��7�n����e�#G,��p�|�U��������	ڟ����lZ���tT�Q�	:6�T��E�wy�
b������O��$�O<����$A�k�
S 6��"7��: (�'��'�ɧ�OĐ��eD�.-�65!#��^4uȲ�U^����_�p�t$�V6��l��Wy2��t�^�g"@�h����/ U�r�'�'��O��ɶ�M�/���?)�-G�H�ȴ�P2%��c�d)�?9Աi��O4y�'��Z�pЕ�\7J��	�E���eb�Ǻx�B]nx~���5p����r��O�ɗ�E�F��4%�Wѐ���l��y��'B�'���'�b��"d[>dh��ޣ/��Ĉ�H�������O���LǦ��� :ZǸim�'(}�A��(qf�#�/_�Dd\�q5�|��'�O�:H���i!�i��A+Ǆ >���1'� �LPp�@�0V�vP��:�'���Οl��ӟ��I�G(�� $Ċze*�߰}"&Q��̟��'��7ق`���O����|��ל[�%�C#�=)�*����_~��>����?�M>�O���AD�4_��=�����L�Ȥ
������i=�i>r&�Ot�Ot �!
� Q�"��R%\"i�`��3��OX���O����O1��� l�6�Ή!���T�*l.4�!۹Bl��'O��b�<⟜��O>�$	-qC�a����+Hvqy�M�$R˓J�-�ߴ��d�+>���'e�@�	�<��0�]�D[(I�sH8 ^p$̓��d�O����O����Ov��|*"!��1��<l ބ� ]�?>��fڢ3B��'r����'d6=�(���&�*H���}h3���O�b>!
��ަq�7��$�Ы��&�L@��I�P�ϓ���Bn�O�T�J>9*O����O�Ȳ&$ڦI\���%��jY6Dzs#�O���O��<�u�i�z��R�'R��'���X��H$<�~P�Y����D`}��'��|�� HM󡪞8�"i	�=��U=\6B�V��;~+`��{+|��]S�F%;�ሳo�&�"s��!=Z���O���O��$:�'�?	��N/~ϒ��BL�S���gi��?!6�i�ց�%Z����4���y��
�"����ZE��R@��y2�'1r�'�J���i�����D	PП� Ԙ�j�x��/V�M���ge$��<��?)���?���?��k\�!)ބ0��8~�.DYT+����1��
⟀�	ҟ��ґ��h���x�m^���!�e�����ß��Io�)��]��L��nV�L��m�P�گ:�L	�����'���2�h S?�L>i,O�";�Y��O=K�r��EZ���Ox�$�O��4�2ʓ!��$��-���R<`7��&O�n�#.ͯ �b@eӢ�lH�O�D�O����+ �����aiՠ�ǂ&��R��c�H�:�P�j(�'��[R��U��L����l�$!C���<Q���?���?1��?��t+v�T,���;=��al]�R�B�'L� dӬ�C�<�B�i�'��@r��g�~��5$^7��z��|2�'��O��\׺i��I� М�Q�>&�3���4�V����%A��4�Ĳ<)��?��?����.W�0}IEC�T�.��$.��?������p6A���I�h�O������z64�*/�R�e��OVd�'�r�'�ɧ�鞑)�Щ ����M��@�Աs�����X밈�����=��)�W�`L|i𓈆�-�X�-ul��	П������)�iy��}Ӻ����ɭi�����)B�T��a�*��~�ʓV���DCU}�'��<��F
�%
�����=F�إ��'d�bJ�*�������iI(oq�ȵ9�
! ��p"��,�`�1O�ʓ�?���?���?���)�?d���gċ3\�m�����U��Mo�T����I���u���i����ck��	��Ǧ���>�[7螭�?����S�'�<�ݴ�y��J� �P���Y�[|X��*5�yRU/!y�����a��'x�i>}���(��}{db]��hIܟB�`��	����̟P�'�F7��
Z `���Oj��:���$����m���{ �$�p}�'�2�|O��^%&�a���#^����ߤ���n+4��
i� b>]h�O���3P��m��
�F��t��C���$�O����O��S�OrLB$d���Њ$G����ɤ��~�*��(�O��D[Ħy�?�;��2����Z���	2��HzP���?����?QŘ�M��O�L3�О��KAk�qjD�S�w�L�i��X$�OJ��|2���?���?A�%��X`r��{W�躱� A���(O��m�#M����ğ�	}�Sğ��d�M���4j�/ю �"�n����O��b>IZ�(L*R:r��'� &Й�F��	N��#��[yrN�($,��%�'-�$?��,��̑8�~�j	&D���	˟p�I��i>ŕ'��6m�6cY.�D�W^.Lۀ��i-M�p]�� ����?�0]�l�Iʟ`��-}0åmP)g@&L�ᝍ^y����(Z��'7z�2�G^jO~���
�`AKV�*r�0���":6!��?����?���?����O�`���Ҷ�rzg�P8!�)S\�h�	��M�4l�|z�f:�Ɵ|�Śj<��gcc:�xDA�.՘'�B]�� �͔���'=Pt�Ƨ�,eZց���҉W�̹3U/��Sw���I	-T�'v�I՟����<�ɆY�X��B�	d�$m{��,	�0��֟��'�6��)J�����O��D�|Z�씪{�Bt�CLؔ%I�a5�f~"�>a���?�O>�O�\��0�I� �
=b��1U�ct���F��a�iI�i>��O4�Oj��e�O�T@��ǅ���i�1��OP�$�OT�d�O1��ʓGK�Fk�; I��ɐ�|�n4j@��&_b8���'��f�`�L��O���C)m�a���j����#^���9e0��ڴ��d{�(9��'.�t��ʁ�T��*X{�d���+5Ox��?A���?���?Y���IT�kl��P���"`������M�0�mڶt�$�	؟��Ij��؟�������"PSb"�/Ѭ2��)0���?1���S�'j��@�ڴ�y��h@�i�F,D�=���B���y��o�@D�������O���`=��r��Up���/X6V�����O����O8˓z���_�8���'����)L2.�;3�D�*]a	ǅ��v��O���'�2�'Y�'\B|�Ǎ'c@����l
)^y�`��O�������L����A�?�ĭ�Oҩ�%(B:G� �br��0���y�b�O��D�OL���OT�}�;c1L��'	�$Af��Ɗ!��Q�W�bP�;���'�d6�$�i�]y3��hy�T�da_X��D��Fz���Iş|�����l�N~�֬9�����s<�2ekE" 9
ճׄS�g���rM>�/O^�$�O.��O0��O�p"�fсV�&ਦ ܤ6P�I4��<IA�i� ��'�'�Ob�	g�ȉ�����h�@�OBQk���?A����ŞiX8y�V�"VL �l΃cV�Hg���M�O�Y#�݅�~B�|�^���V��>�6��R�K�8 cB�L�Iϟ��	ן�Ay�iw�ȑ0��O$W�.�Ըؕ�{3�Ab#R��?a"�i��O��'v��'���	m�.!Q����@p�H[�6L��i��	#mx�	0�OBq����J.v$ �p0ج��.�.�D�O����O0���O��D'�"b+�BuNˊ|N��4Kɫ�-�I蟀�	�M{#�>��Ć��Q%�$PW��(�����ހ.�"娦�P@������i>��6\���'ԭp
� Bd���F81�ָ�wK�fa�t�`M6�~��|�R��˟�	Ο��T,�v/��Y�T�"��8J@l����ITyB�dӬ��O����O˧�@�AeF"`�BM�u���'�<��?���S�$
\Mx�08Ǝ�a��G.S6J�����Ŵi�(��R��*��KX�ɬn򈠙 ��:<�
(3rGȭ0(����̟�������)��ay�(~�d\�PD�'t��Yn�>W�AO��D��d�OZ�mZ~�k��ҟ|�6m]7tN��Pe;oW�`��d�gy�=v�����pC�GZ�P�$�	ty"E�<�`���A	B�`�9�!�)�yr]���ȟ �I��0�	��<�Om�����H�S_~!I�jh{����r�{�:	b��OZ��O̒�X�$�Ԧ�݅t�B)�c�%1�Ą��T{�����ʟH&�b>A�	�̦=�?��8�҇�	9/r���*��dV��̓(}(�(��O��@N>1+O���O4H(D�M�k��q$���;��0"�OZ���O>�$�<�бi�r=��Y��I&J8d2�jc�V�)E�S�t�?�@Z�d�	k��<��9�%ܻL�\IHF���'���'�
a��枔(����T��՟��'���Ctm\6C�-*P�D� R���'�R�'yB�'��>�I^o"�����B��}ѐ�=(���I��MS�M�>������?ͻxs��#��l���"��b�lϓ�?���?�U�Ǭ�Ms�O&���L�8����"QzQ��I3J�*x�k
�T�2�O ��|"���?I��?	��GX��QOʤq�<���	��8(O��n��z�'7���D�'z�6ʻIb��ѕ#��X��q�tF�>���?�N>�|:b�S�(�>��M��y� h��G|��i��4^��Ɏ ~��Ӕ�Ob�O�˓pf���^��Z��TEc�)��?���?���|�/Oܥm�<"����ɯ!Ƶ��iy���Vn�*v*��	��M���>����?�;AX0��U&w�I�C!��Z��£��M��OP`ks���d��D�w���R7�ˡ�	���!z�	i�'�2�'���'��'=��˰�PaG�L�q�H�S�Z���O��d����C@�Uy�Ga�j�Op����P��t����B1�:�&���O��4����(j����^<	a�A�S�T}pr��T^�X�@�N�'�ԇ����4����O�$1I�u��_*:�|U�U )�T���O�˓K��&B�$�"�'rZ>�Ø
>��u:E	�X�� �&�.?DZ���IR�S�t�J1�A%��R�\<ï߃,��l��M�YNhE�Y��<6tB	Tu�	4 ��`{�(ǻ"��G9��\�I柠���)�y��e�R����>	����U�K3�Xc� ��iHL���O~�m�S�Qi�I̟���ԴL�J��zkH����f�p���O�h�#y�6�j���"���"�O:ܱsFħ4}D�R�	X.�؊�'e�	��4��͟�	͟L��Y�4/V�!�ũSh8:����4��i�:7m��+t�D�O^��?�i�O|�oz�)Q�I<8L&��b�K7�N���F���@�II�)�:[4<n��<!1�VV���JA�]�\p���<q�dr��' .<$�Ж���Łxb:I�,T?	7���t/�>3�axr�wӒ��d��O��$�O�5�bgh8$��C���&Nn��O���'k��'��'��xa�Ϊa�\�C� н����O|�P�BZ'FG�7�C`�0N���O��s5�G�p�ԍ�QæG��e"O.=��gF;j_��ZU��Z0(�9A�Oo��(��I�(bڴ���yǊ:fԜ:%�OvA���<�yb�'���'�8����iq�i�)Ƞ���?��IȨ4F��Ñj>؀�.�s��';�Iv�'��T�.�%�\��T�ƅ	~~B�bӢ��G!�O��$�O��?��̓%ٔ�	AJ ���%]���$�OX�$%��郊,{�9�Uꌿa�~�3��.y���cv�@��'t�J���]?1K>Y.O��l�7) �����y�fXB��'Z\6m� &���I��йj/A���A-U!�����ݦY�?�CW���I,���I\��XT!>��jEAZ�R�R� R"ҦQ�'GJ�J�*��?}�D����w�hp��D$���c�/Ǭm�RLJ�'��"�C<n0u��ؔO�����K�"�'�"{ӄ��w�?M0޴��+����j�6��·�2eP84�J>���?ͧ8��e+�4���ʷ%�tIipD��9���D�z�AՔ�~|�Z�t�?�'fS	?r��)��I"t���Iw�'�,7���O$����O>��|�q`EQz�hp�ߐN�d���x~��>���?AL>�O��Ɂ�ڛfn� �f�U��8�؉6�{!�V�$�i>A���'7J�%���h�c�\�����~v��@�3�<bڴ�`�kcѩ*<����,ٿ(�����E�8�?���@ʛV��Sr}r�'&h��5瞹8��� Rkđz�f��O���A'(�7>?�s�T�pq`��py�9Z�`�c,�
~��vH��y�U�,��I�n�����I�`ٓ%��<���شt���)��?�����O�6=��}��킟>�hq�
	�.�1Å�O���6��I�; 7-k�� ��b�b�/Z�|j0LB�0��X�?O��������~�|�U�����@a3̚2���+e���_:����ޟ�����4��eyri�,�!A�O&���O�]�¢P*_�x��֦{� ��f�:�I#����O���.�]�.o���6Cdd���çI��I$l��(� �ۦ!M~������ɛ��|�ï�U�Ӂ蔕 -h��Iퟘ�	��@�IQ�Oj�L2|&�����Y��F�T�2�gӀ<���O��DZ��?�;/\Bq�L-��=�-!SӐ�̓�?����?ٔ� �M��Oq�DH�4��T㒷Gͨ<�T̡�(�A��ƌ|�'��Iߟ,����p�	ݟ��	4F�ݘªнi*.�
��K#1Z�'��7m͠_���Ov��?�i�OT��j�� ̎��&O%)"�49���E}r�'���|��D�X<o�P��6m?��I�F��
7� �ӷiOd�4��T8ᇹ��%���'�j��`�E�.)ʌkpNN1|��=+c�'���'������\�X��4\w��I��6UF0��M�V*����$+��{�!ڛ���Kv}2�'��w��l���Cb^i�F�Cà��&��	g0�&�����۩/����J�������9@a����ПI�ଈ�Ev�����D�IٟD�I��"�� AuB]�̊�3�8���mQ&�?���?�r�i��<O�bGxӺ�O�Ek�M&�a��@)e�
*�e9���O
�4�<]��bӞ�Ӻ���0�t�PGeZ� #����"� t 00�pT4�Oʓ�?����?Y�����R ˽a{�l�W�����%J���?i/O@oZ�hz������	N��:[�1b`!��laa���y��'���?y���S��.)$@՘�Y"�	�EN�/���CR!�f�
aU����(�G�ɦR��Q�md<x�G�:r��,��ҟ�Iܟ�)��Wy*qӸ8�s�3���!W0g�� �R�z� �$�Ov	oZZ����
�O��D��	��I��  ~�sэ�5d����O,4vGhӰ�;hҨ�3��?Q�'ܔt.T��;�
I�5�z��R��y�Q���	����I՟�	���OZ٪bg��Lب �LJ&g$u!�#pӬ�s���O��$�O ����DE���E����H_�]y8t��V�2?BM��Ο�&�b>���F��4q�ؠ����s W-<�ϓ�Ĭ�Ai�OdՙH>�)O$���O>��G�:ਤP�^8j��hC��OF���Op�$�<� �i�z9���'�"�'L ɒu��w�D� ��B�=��a�Ք|B�'����?1���e9N��b36vW�� g���	.߅hb�$(�n�`�ӁieBn��427��w�@uKR�� D���"g�������I̟�F��w0J��QA��r}hS�׈�1��'.�6�E�l����O|�n�K�I�����!Ϟ��C�	���y*����x����O����O�u3!�rӔ�Ӻ��BC�J�L֜6�lp�" Q���\��O���?1���?i���?Q�.֩�q%�\k��R�(Z�1!
}b+Om� %Sș��۟��In��ٟ��d�� 4�:R�5�΄:����O��!��	��"���`��Y�r�&���ɑE��|Y�&n���'��(+&��C?qN>�+O�(�j�'���<��cKJ�a|B"h��u�a��O^-��iǷZ����/D�l�2C��OVpo�_���	ן��	�$kg�)>��p�!O�=���&���1��lS~���j����ӯ$�O�w��e�$�q0a�J;(���y��'z)Qb �8��L�P�H:� 6��O���O��m�B���ZC���|R�ǸU����'%�$P��r��C_g�'�����f_ћ���]�U�p!
e�� �>�{7� (hBT�O�㟸	p�|B_���?��Ə�	N��GڻI����c)Q~�'At7K*~�x�d�O>��|���I�yN !{d(�0,ѩG	�~"��>����?�O>�O��g�#7����O]�@�İ��X�q�D�B��i�h��|r4ʵ��'�DY"위�ʜX���3��xrU�:��9�4<k, �v�6(P��v�D�#�4���R"�?!�dԛ6���u}�'i�P#I�HiM��,�.<� �(��'7�H��{K�֗��HR'RFW�)�<)��ޞN��҄-5)�ѕbK�<�,O�D�O����O��$�O��'d�E�c+F&p���3�N��TR��i����D�'t�'5�Owb w��t��Зh^���(u!�?3n��$%�)�S�`1��n��<�Qɍ+?8u�C 5�(lX�<��CU'/��􉠨�N�l�9r�Q�ū��N��ҸA4JT�5�f�� aI�%�a�f�W*&|�D��_� �T�R@_ڢÁ�F	T��3�DBG1	D�]�2t�D�����̉l����0G��a�FE�<�"�B`t8i�OA�ccY�=���E�y��-Q0�!TĈ����:B�|9� C��hɄ4@��o3v$��Θ4Qd�8sת��8\x(P&�J�I����G�4y�B�(�	s�ֵ��GO�U�H�q�E\�!P��^,�G+x���s�ːN����C�Ѳ
&L�WA�\d���'xB��g'���CO�0I��[��U�Ti 6��O��O����O���O��'t<ۦ��k>��H#ᑆx~��I�4�?������O�N`�O+��'���n34B�,p���nG�	` ��:�O��$�OX9�7�(�IG���1Z�| Ӱ+Ɇy���9�k즑�'AN��$�l����O~�$��Ԑէ5�l�.[��Rũ�&X`�2���M���?y)���?K>���� 4j�M�}9�<*E,��N�*��iE���PCg�:�$�OH�������'��	�h�L�UJ�*_�M�5�ظ��Z�4C���[������O�	�%Z��Mq�ǔ�,B��2@��7��O���OJ-��v}�W����^?�M�B�(�j��*~P(�`�k���$��W�
��'�?���?Ie��, U͍%�q�1d��a͛��'���!�>1.O:�$4���`xǉ����4�Q�� 3�IWQ�x
G��L������� �'�@�¤�,<e�𪉣c�|�F-��L&����Ob�O<���O�-�T�כ`VPb�UY� 8Ej�Xn���<���?�����.z��!ͧK�J�	��Ǳ��p�kN�v-h�lhyb�'P�'?r�'�j���OTT�g��#W̵K�F]�VS��#�R�x�Iڟ|�IQyb�W-v��ꧠ?�g�FL�ҳ��`>\�
����.
�l�ɟ&�$��ɟ��w,�Jܓ��$p� �ᐩ���ؔ32X`lZן��IryB��E����?!��:�l?�@䱃+7;B�zs�6w��'w��'މ�����?�XSO��`��}*&8!�n hvjz��˓4�f�C�i��'��O�n��;�"X7Y@���=R0t�c��Iȟ����G�׸O���`,�7[�<�Zd"�o��h��4��`�S�i��'X��O�lO��W�rX\��ޤ5*4��ʆ��nem�˟x��͟�$���<���W$i��8yG
�s�:yb���i_2�'�RJ�A\�O��O��Ƀts̚��
!�|x"�Mׯ/s�6�OޓO�������O��	�A
I�b�2G���!�҉#��6��O�����<I�W?}�?�P�/A��Y�Jښ
.���Q(��V�'��B�O�D�O���<��b\�K�&�U*�h���[q������#�x��'_|�R��]����1����4� a���RY�7��OJ�O��Ļ<i�g���Odx�:v���E?؈��&�
޴�?�����'0"^���ih�ri!����w�I)w��x-F=cpT������ICy�R�)���,9�X}�B˃�!�� j�[9(6m�On�Op��|z����ӡ"����������	C�0�6��O�ʓ�?������i�O>���k�\�W:�`A�[���|�S`�M�'4�W�`C%f8�Ӻ�0%�#��@C�"�9A�ԣ�P}��'�`��'�2�'V��Oq�i���뀣X`>� Y�/�% 7Hj�|�$�<���G��ħT���!��'}[�1#��\�knD!m� yF��	����	�,�S^yʟ���T��(ujr9jB/ۨB�Ea�N�D}b$���O1� �D��S��a�g#����3O�<@ڊ�mZ���I��(J`[���|R��~�M�E�v!��ݛAr>����*�M�����C��3?���~�M�9%���(��.)��� ��M������-O\��Op�O�)�Ϛdy�)����(8%���f�Ɉ.��c�D�IGy��'5x��B�H>d҅�%g�kl�5�	/5�	ڟ���h���?�'Ū�*��?=�R܀�f®4�	ٴ,Z���'�b�'�_�� DiS&��d�ֿ.f���3�-�l9�/�>���Oh�+�$�<ͧ�?���H�4ʬ��u�^I���OJ�L��I���	��`�'+���AE)�i��^�v�B�дo�~�P�CC�Z\tn�ޟ&������'7�'Z\�	S�	ZI�\�P���b)��oZ��x�'	�KT�.��͟`�I�?��,#I�T$B
P��p0��	:g�O��ĳ<��J�_��uwꘌ_U1�t-[�5 �	�E���M�)O������1�����d�x�'��b���%���P$/O�!�l��4���O���x�H�s�p��M#ٔ ۀ�'nR��@ǽi��H{Ӑ���O������d'���wCv�����y>|�����91(ȑ�޴�?���?1O>�����"�yIC�6��X��
�
���n�����ܟ 
Є�Zyʟ��'֒X��P�>��9b�/뮴��6�	��O�B�'Pr-DL�.�r5$��b�)
q냁�~7��OV��F�a}"_�(�ISy2��5v��j�r���۱&Ϝ��e`���M���J���?y���?)��?9/O����J74	�T��\�wj�"`陘~�}�'���D�'�B�'��@֔�8�@CBטt��"G
��Gĸ`��O����O���OJ�9P9b�5���0�� +[�@s,�G�d��iN��ӟt�'Or�'N�FG�y��%k�=AbHI>�˴��]��6m�O:���O��$�<a%�πP��S��Hc�Z3D���@�-ؙ�@�ΰ�ֳi��R� ������Ɏkj�I�T�I=D�N���m,
iS�F��0ܴ�?	���Ǭy&2��O���'����&X�q��QY��[Cnʓ � ��?����?��m�<�M>��O��i�qp�
�N��h���4���إbt�l퟼��ӟ�������PD���-R��w'[yx���#�i���'|����'}�'�q��0ڲ%S b��)�EZ,"s(}�6�i��|�u�"���O��D��0��'D�ɘ-b��a���9&�r���?�i��4k>dΓ��d�O��?��IV�t�K�ҟ. �٢�	d����ٴ�?���?���A�B8��_yr�'��Ğ9a�@|�A�ȜA@v��4)7:��|"*��yʟt���O��dXd�? 8`׎�>z�t�rf�Ԉ�^<��i����^6�����OJ��?���f5pBR�;��S�� *�H��'7@�@�'��⟤��ğ��';x|��m�~3�X���I��ٰ�(K�8'����$�Ohʓ�?���?	 ��X����޽<�pY��55$H��?���?Y���?	-O"��PM�|:"��LY�&�#,�,9��Yʦy�'�RX�|��ɟ��	1RG��	6��a!bh
6&�$�S�U�o65�O���O����<��'݄���d!2k�5<$1[�& 
u&��A���M�����d�O����O� �5O��'�4�cE�	y�ua&U�X���4�?y���$�2i"��OT��'y����"}/����	�af��H�	Uf�"듯?9��?��Lq~RV����%WZL2�� $(��H�Æ�IR~�lKy�N����7-�OH���O��p}Zw)�$�
lc<,���l]Ȧ!�I̟\�Ut����ry��W.�.�8�#D�s�Xp �h��iTG|6��O��֛6�O�z���D�$S��RG�]	�b!2���
<rl�9K�*����+�������B��ar�~��K9�MK��?I�""n��0_��'%��O�M��X2oڈ� ��.1p�ǽi[�]��;��|��'�?���?��i�c��e�3H�L^\	t �uܛf�'�d����>/O��d�<�����c0Jl�G�[�T�3w�[v}bcY�y��'�R�'�^>�	�F���jwcG�R} �D��{�$Q)�/X���<������O���O� �A_�b.�M��ۍ9�%��
05��O��d�O��d�O�˓hL��5<��1ˇ���`=X4HT"��S;qS�i��	��Ж'��'�rb���i�#$��� ���""�=r��=����'}��'^�P�0�'A���i�Ok�^ �d%˒���\��$�g7@{�V�'J��՟�	՟,�A�'?�'�B�;��٪��ݐf�[�-�1�޴�?����$Z�{ (�$>��I�?�;�/s9�Iq��!7��S�����?���k<���������I%Q��t�d;�P��ďǓ�M�,OF)��
R�uX��2�d��h�'�噓c�"u��C��Zΰ��4�?i�Y[��Γ��޸O������)X��DD]�O��ժ�4zB��3�i���'���O�`Oh��Տa3�0�1���G�L�c���5�dmZ,q�u�?	����'T�!H1������%�:���}�0�D�Oz��E��'���I�L��i�uc�#
9b&�jG��*f"ao�|�Ɉ6�.�)���?���z����o�3%�vyЧ)7	n��c�i"�2c�L��D�i��y�'Ӷw��)@�����9"�!�>�%�Q�<A-O��$�O.��\�k��U�s�t�E�%�\�	��L����>�����?��C����שP�X�8�HD�����w|��D�<����?A����$	�@o:\�'OPhȹs
]�Q���A(��2`)�'���'��'���'�$��'6�DB� O�5W& �󪄨�T�9�ϲ>���?�����*{��$>%���^�HJ)��_P��0�#�M�����?	��=�:!͓��ɬ�h���X!j�pY�c�A3ha���'���- �d��I|����2F�<.�j�����c� ����C�=@�'�b�'�V5R��'��'z�I�+Y5�	Q�D�/-m ��!�,$�6[��9�,ͺ�McCR?��I�?M��O�`"��Ѓ)V�x�3	�k�BQI�i�"�'E`�!U�'
�'yq�R��<[���ɑ��cf�A�2�i��0ћ&�'�R�'���I:�	1lƙȲ��Z~�y�a�V��lCش8�� ��䓓�O�2&�+ߺ���$&�X��ф�|�67��O����O
�k�/�O���|"���~���Dp �c$��a˄��Ջ��
��	;��'�?y���?��Ȝ�Kq ���䌞dޠ)I&C�f�'������>92T?���ȟ��OԵ���E� gj�Yq��+RL��xR�|��'��'-�'�-YW!1j�"��R�K�W����Zp(Qw�'��'���'�'���O�@�cǻ>�ČJdgAO��=�iW���O:�$�O���?�uf�#�?��=s��4ah` ��}q�F�'�2�'q�'�"Z�p��l��$ٗ�Ӕ\DA�-I��I�V���	����y�,ò((�����싵]��8���'^��B��˦��IZ�I؟�D}�ɣV��H��O��@w^%H�M���?y)O����k�S��ӧV�PИ�AV�!r��q &K�.�~xIH<���?)F�NS�']��M�ꈹF�J�(�x8�҃��<���Q�찄�Y$�M���?����J�S���8'�X�S�:~�� vA*CB7��O���CW��Hh��'�q���2����nP.�����g�A��i���[4aj�����O������A�'��I7d�y��eS�q'���]�3��jݴ^��Gx����O���v�\��`��NG B�`|@�-�æ��	П��	�l�Eb�O�ʓ�?�'L{�ꏌ(�0´��#+$"�4�?�)O����=O�S�P���{��{�l|z�K��I��,+c���M���;�|-�Y��'�T���i����$C�$c�8iR�ε<��Q� f�^���
	T��<���?�����DËU%Bm��&� p� Io����xA"f}�X����Ry��'��'�x�e��!iH�#S*�
~ �Ң),�y��'�r�'��'k剽����π  e)u�$)�Z��PgP �L��i��	ߟ�'�2�'}2A���y��>�=#��U�E��˛�u�7M�Ov��O����<Qd��&�����X-1}r�#�́�qv�\�uǌ�Rh�6��O���?I���?I��<�+O��:P��H1��!���e�v�9�٦	�I�4�'�"�$�~2��?��'Z2B��w�E]-.��*vGA�����O��d�OP�D=O����O��D�?��V�O�N�	���N��FJ~���V~�4�F�i���'B�O,N�Ӻ��N�=�� 
sC�7Y��!��-�IП���ep���I��If�'}�M��Ĩwނ��j�z|
��I`g����K�]>�����U�~ 
�C�Z!�4+���)Q���6���>!�<�r(Șɠ��q�Q�'=@8�SL� ?��\iЏ�
�Fuڒ��45�lYR�j��.�*�@R���1Z�F�&e>�K�)	*��|p �SB��e��:�zA ���+�њeE�2MnS+��H�x��S�ciÄ!]<b�������|���O���OJ��;�?A�����"_�<0`$ֈ�@[3�V7�M�f^�4 "����@�`�#��0�[���3�)±n������5�c�D�b�b��e��+�NY(R�_:�JJ%鉫x1X]R��{�Yj&J��cP$����O�D?ړ��'n�р�Ë�7��13tLA�"h�p�'	ta���9
\Jpġļà��y2N�>�(O����M�V}��'�\ �Ƣ?kr����\<Y4�Y��'<"� /	X��'���$Q�H�acP�-(�U�(�Tp�۲�BD�F��R�,��I�X��{×�c����'��`����?X\%m׭qƐa�L���	����'�p�!Cޭ**T1��U�k.	a�y��'-ΙS!K޷b���`@Ô]��|
�'�06�ǉbQΙ0�&�'�Ήʠ����Ŀ<� I@�RL����L�O���'��Kd���a����F�7B�Q`��'��(Q*�"e�by �l�O�Sz��j^�(�l�J�bK;;�=�îY����Az��
�eЪْI
�_T�O�$=�g��6r|R���$9�eHL��ऀ�O���5ڧ�?��m-sV>��/ϼOC���U�<�W��k�V�2��ϵK4 ��
QI��8����Z���(���t:�M�$�(nZß,�I՟`��E�M��	�h�	ҟ��0{@>�S埌Q$rPIۀ��'� b.�9����,��t�cJ�#�d�v'W�q��U���"?��+����>�O཈c�D��� �+ܨ�z��O\�	T��)��O���O����*�
�d�R ��G�hHbb�)��!|O�#���su�A��G�����u���{�4�?AH>�OM�I�[R#���H�
uXVѺMN*�qc���>���ȟ���ٟ�Sß��I�|��@ͱR���R��6(��Z�KN�/�Ԋ������>4l�+lV�s�7+���׍K�(/���$M*��>	�$�
�l$�J$KH�����[�"
����ϟ��I���'%����==^(�"�D�9���Y�n)\�!��-8��t���t��M��͚�1O\�l�۟��?�O�x�dH� O@ ��a&��0�'�(Tr��"��	���"s�	��'�VPĪC�'v���cRh4Li��'>����ה�-뒠	%*�ҩ�
�'P�HDt�d}��F�ObJ��	�'�TY��H�m7>�����#]ֆ��	�'�0�SN�2v	�cM-W�|�[	�'�P�����S��T����R�~M��'�-�VC
�^�Č�G>��+�'��Ƨɰp�"�Ɣ?gZt�
�'��l���I'@.�lK���KP(J
�'7I�E�.�>�@���C�\X��'����<�Ty��/�`�1�'�j���(H�Ҋѳ6'Z�+���;�'הaЂ����Y���� ���'qF���̌"@}�9������͊�'��ŐQG#im�`�$b��ꜝ��'6�����������I��)�'`������6Gf|L(wdL=Q�T��'�����ƨ&�r�/�V��yC�'�65`�%/�J�	3B5� j�'o����
B�]��s¬�wyFdc�'�,L�w�Т&��%ÒǚtrDt��'{.q)�B�����ܞd�4���� ��RD8���ٳ�R�B�<��"OX(I@��(����˟ :��8�"OL5�h�%����׻0��!�E"O֨A��8��Z��J$��"O%��D�r8r�@K�6�Dx�"O���{���6j:Fe�a�%M��yRf ���9)�B
-��LCe����y�_'VR�9yf�M�+�H���G �y��];<�]�%�n�Kq�ײ�yr�e�H�'Ć�oC5�`L�&�yb^::�t��iǈXb�"��'�y""ӘY���$�B�dZ�
�a�y�GU࠼�c��rî�
�y�ߠ(����˫?���`��B�y� [�>��b���;�b-dF�1�y"l��+e<pXT��==:�	u�2�Py�E��8"|�X2	�%��Cu��s�<���T)����h��66�3�E�G�<y�ɏ����7h��I�8I['��l�<a#�ʨҷjz�4m�G�
j�<i�NĎc�� nI�����rTd�<A�^9��g��_�����BV�<�2�����2D�i��08�.j�<	f�1kбp��݇`~\i�&�P�<��
tp�r��P���Bd�<a��H�wy���fC"��k@z�<��C�\��i�"���JA�]�<� @� J���J4�U�f�����/�[�<�g�U�_:ְ���ү��%藯�Y�<�)Y(H���F����+�$AY�<��� "*	�e�vK�<;��)q��V�<9*��xpe�RK�*�<m(p+�R�<Q	��yԁk��-��z��N�<�&OM29�a*�iצ{�b�Z�DQB�<ف�[�#X"C�  �1rQ��f�<1�G�HJ�T���<�0�Rf	a�<����b9��i S�r5��&Q_�<�3mˤ+�T�Ƅ��o�t;�Pw�<����ybR��g�*��'�Wh�<�T.R��Ĩ��]H�*�	�e�<)Ǯ��%�0�� GQY-���y"X.Wz�Ap�ÛG٤q���yr�� _���L�k�:=��G�y��E�?Ȥ�"o�'^�6(��(��yB&�3�Ĉ�t�C��l��c��y���!O�*|�*���T���$� �y�� 8{��uH"�
h���p���y"O'<�N���`�4u����y�W��B�a�&���L	d�_(��'���K�$*�'��$�A冷9tB`�E�.	XM�ȓW�RupW��	\a���Ub
�Rc�u9�,Ts��+M{��IU�����e7�a˃�ɧW�l��	<a~���'z��Mв.�t��dJ�8�����T��?��I(E@����-�,���D|�WM� ��'���"� �<�@���C�E��rtk���/���B�-��(�$ r�FY�"O��×B+ d�S�=65�$H�
,H�]j2[�Y�R+Y�d����F#0D�S����w��87$Q�F���F	��P`�H�'�z��]�kEFi�`L.*&i�SR^R��Rl��i$��m�$Yu���'#�ls�'jS4��'�b��/�[ǆl
�$V���Ó8	�x�lBDa�9#� �3���Zᚖ\Y�Yjf��6�ځ*�FI��.�4��yUU�1B��$�U�N��ТΎx^��L����I�]q�b�$!�\x�FŹ2����S?)j`.�Q�����]����cR�c%Ժ#�!��C�X\@�ģ¡!-\ ��]۸ŉ�	�- ���n�5,�j�3�C�\TP�AD�ã%%]��Og�@�^�8�C�@��������xb�P��� ��(��؅2���fғ&��q)�^�f�|kebh��*D�����Z)�`5�Q#���U�� S��7�@�{���g�ax��rߖ�� ĻFv�<�ӦH1�&�x��I��J�$��&`��[�e�oy�*�<Ó	�t��Lm������Cl�'Z44 ��`GX9!2m��<r�J��O�O���Zh�J�$�(A�kн�y"aKMT���4G�`��<�S�]�_���Bi.�� �'=~���x�^�����!�2tIW�Z۰��Anƈ1�a2�Olâ�A�?ʚQ����4tz`mR7�a�h9�KIJ�tT��F�j�0:���G�j9`�	��2�u��ι2�
�>q���#�X%+H�]�)ץ����v.��~�<%���P�c^�qf�T!g����#BH`E"#^��p��+s���'x(q @ӵZ<���w�ӨP�X�J�O�O�r�c�
\��|mmk���
�'6b�V̇Q��zP@��4��$:f+��-E|�q�OL}�,�Q�ӣB
��)O���PM�i�����h��R�@�ʴ
O�@�ү�-	LT��o�L��0�KQ�}jҖ�T;x&��0aZ s=���Qh ��G���1B�I�����	?��3F�Y�?i����0�IC4����]���EzҌZ�+����L=5%�-�&�D1dIjg�<�I,��*�J_�suԕz� �Hܧ
mh�3�}�����P� �%��%� ����sd�
���%~x�(PFP0l��;CnM� ��D1�g?�@�4}di��֝��%Zӎ�^�<9&�Z*c��]�D%�J�l��]�<1b����=��f���<�R��|K�����T��J�QX�4�� c�
���M�R��,	��
2�
�qb��y�Y�\D��T\�.q�a��k�9ÈO|0��3�'h�i���CR�A��GJd,�ȓ2|���6휕4�5��	D�\�ȓm5��f�lV��	�u4y�ȓ6.$d�#K"	xL�#~:����o�i�I?<n��Cq��=[�H0�ȓ8q*s7���A.
����@vC��ȓ&�:,�s˗2Q����P�͎C�#��i(&fz���bg��"A�jC䉉AB9�6DG�-$^��U��-�J���%2�La	�҈ ����(D$ވ!��܇�	�|+�\��?OV�3i���e���!L�$$�'"OZ0
K�$W�Y����O}�����I�~3JJ��5N�3&V���Ⱥ���4@��B�I/E��2M
 )R�J�Э5����Ě�%۴�"~�ɸ/
^(��	�h��"M/RbB�	�Tu �	�M�	iL�a,�3	��j�^h���'�̽���϶$��ٶmo^�"�'T� G�����)Ua�)�����'-r�smM�dm6�u�!��1�
�'H������m�hX+e���: �ĩ�'��|;C���	~�|��@�9[�1@	�'�����"����-���?~P]3	�'� O�-���IFj]"!��'h����?E�H��0NLR��i�
�'*�9p��
�QF���J�L��	�'����["J�UgPt���1ZC��<�ڑ�Ԍ�YO|�˝E�B�I�� �A��.�,��0ilC�I?���`��P��%�sK >u$B�ɨ(3�z�E	h�昪6BIFFB�I�+�¨����?zM����dW~BB�Ɏ"'F�q��9h<ڀ-�g�BB�	�D���������. �C��~�XB��B� ��mR�;d��B�kc|B䉩t�*���)�=��b�#�ZB䉼��0��I�[�����NNq��B�I�eÈĺ@i^r^Z}��-�_�C�ɛ"#p�	"�Z�%�Fej�Fŀm��C�I�Ys�Y"�J{���s!�@t|B�)� (�����3�"��B�6!�
�K�"O���`�e���[��O�� Q"O�|��'��nҎ%H7�Xg�2�"O�Q�-w��3�/ן,f���"O��M�Pl�e*);D�@ 9"O�y�Poف6�&���AG�:�@!�"O�y�V�T+F�v��p��]���w"O.L��&I��5p0�����"ObxRC�\�J��)X�Þ-p�0��"O��J3�9�*4c��h��"O�e:��F2v8�a�<Y^�Qq"Otu�֠l&y���oF�"Of��AG!ތ�(��̸O�$���"O���W/�K�f@�/��(��qq�"O؍Ru�dx��P�F�#�p��'L��"@D��	�ȟd��t��'��Ǎ�wک� �ӷ[�t\��'Z0�*栃�0j�x�ɐU{~t��'F)��癡,Z T�b-ɓ�L]��'E�*ZU��@e#Q��I
�'Y���6��o�شBM�EX
�'nd��CӡSjTI�GJv$e��'K����Կ4�mtI�zV���'d�yґ��E-��8D�	t�
���'"��]�+�� #d��8���j�'Xn9��CM:eZC�^�6�����'�81��+G5XD�A�'-����'��;��|��))%ϖ�'��9�'�`up��J'����1iU�"�0�'�x�:��
*qHޤ�⍺"�PE+
�'NT=�3eݮ�ڨ��A#%-�
�':Lupa��(\�>yy`E�#NJ�8�
�'+bq��3l�ܒ7Ȇz�2D"
�'WppS��*v�
TK�%�u`
�'lƱqǡ�lO��٣� ���	�'T���͂�e�,S"��~����'+���"�ŠP�uH�&&uA��	�'��z�q#bݠ��Ԙp3~���"OHɥ� f�&���Ē����ʏN�<�ucٕMN�l�e&��o�8͸�̉K�<����U@�m¢�Ӡ�~�� �FL�<���1��(����%.������Q�<IG�T.f��ի%;!��HB�~�<q A2_���RA��AG�����Ev�<i�,F�R�\ic�H�b! ��u�<q��Y��H���B�'��H�"s�<i��(x���,-�JQH�Lp�<)N��H��7߲"��1s��s�<��(��F��| 6�8�]�(�U�<ѧ,j28���/H�J 0aI�Q�<!�-����z�ō�;̺�S�&�M�<��(��v8�a
�H�")LЫ�̞F�<���E������6�d���d�}�<���.�U���b�6}��
Nx�<����V���F�� T�u�<q�jۛD+�e�%�u�)��ϢT=hB䉭-s��$�O�b8%��$0C�	�qv�Xv�D�{����j~�B�	)~�{fk�& 	��	�g��B�N��$�]?y�d)(ԁE�c��U��DeB�+��ϊ�*�֧��2��t��P{�0q2�5��p3f�; w�t�ȓY����E�1�P��G&����ȓ(������tbѢ��hu��S�? J�0�$��kY�d�i�)�6�P"O��6"8�t�2�ߩQ=j !"O�$���HX1P3A�.n�U"O%Q�V.l�����@�a+~]�b"OP����ȍ"ֈ3���]%T��"O����gn��A`L߅O� �6"O2,��	�*~���?)f8�v"O�9��xj\���E;	diz�"O�Y�$��8��,X@K��Y�JY!g"O�%�Ō�-���v�]2RK��y�"O��Xw��7?#�����0�y*"O:pr)�����S�H�y�A2b"O`YP��KQH����n�q�f"O��Y3%�O5�!pc(�o̘|j�"O\	9#ҙ_�bm��F�P��&"O޹"��[�G!�]��g�,����"O@�����_!rx�@��P����"Ohd��#�e�P�F*^9E�`���"O�l��I�Cu�GJϖi�V�B"O��be�q�zd�B�D���x�'"O4�@�,b��&i
-~��a&"O��1�-CWxb��z.%h"O��R ��U_`	"�Q�/_0H� "O���D�8%��:ck�sG��qb"OT-ň'5R��ak�+��a��"O`u9��%R��tj�2]<=�"O��b�MG�u2q��^�"m{S"O��HC&]����'�ǭ
�!��"O���`�V
T���4&�7D����"O�[��ĿE~�{ &A�4��H��"O [��$�r�j"�
 ��2"OL|���*x�LPA�M��*��XP"O$�K#"И�h(�&��]+h�"O2��c�ַ*le�u�l��"O�Uh#�ρQ�t�˴c���"O$�s$����@�I�8�R"O���#�1f�*I#���ٱ"O�5�`/](&P:�
"`CF"O^�P���?'-Ґ��hۨe��X�"ON���Ɇ�� U�
�p��@w"O��V�R�T%��Be�ɅF����F"O���ύ�q���#w�՘,
F=P�"O�����P%J�X�ѣ�{�rL#�"O6Pz�ꄰP�zd�N�g�0E"O�و%�A�9�9�H�C�T�@�"O�9@�Ό|�*�W�݇�6Aiu"O������P��!(A��	�ڝK�"O8�diW#0(\X
f�߁0�Ѻ�"Ot|�0C[������$���T"One��b���B�I�%b�qX'"O �J�c�at	�I�!�D �7"Od��᧟�9ѦR��j��Mh1!�dN�V���3�;`�� �3���-!�C!�^łGJ�(tx�9ssA�!!��T�!Z�@&XZ0	�aBA�i!�$K�x4d��Ł���
uZb�G�w�!�]�"&%��Λ����R 
�F�!��"����E�"T�z�KqMMv!��C /�ĠP��$ߢ�Y����W�!�ą�t22\Z�M�*{�t$��� /�!�$��!�� ���O�&�>��!$�!�ĉ�(1�����O�J������8;u!�DU�Sx��5�Z�N���ڣ�D3zu!�$.��qH��L�^�����%h�'��|
� Pm`q�S�5�z�+�HI����"O~8����$��9��h��l���E"O���@D$Ҭ2��҇^����"O��"S�T4��)��H.?p���"O�����ݲ�g�1v��i��d_Q�L��i�$`i�Fb�jA!�S*���S͔ Kr\r�!]�],!�T�cz*����G<�a!y7!�Ube�d��ůEz�ɀ�]��!�ēA.� �^��3�9E!�d��j��s�Ʒ'H0|�c-�+/�!�$
_�R�����]d-����2Ex!��^@ሠ34�&>T�艥�)iX!򄑩	$�
�*PM�c�N!�D��&�;�#ڍ2�UP� �3;!�$K�$i�6ɯ?䨨ȣa�!���	�\��*�!E����	i�!�Q eWF��F�R��X���!�$�=~h�)�*¦K��	�Y$Q�!򤝻0
�4K��\�?����&d 9/�!�DS1� a0Wş'��4,�1�!�ڼel�h�Պ٪k58z��]-b!��(�T�+$�SO%ڄȁKB�?Q!�}OXEၥ�j$y�
["J�!��L�y/z�g@�3΀�$R�ZA!�βL&�L����o����4:!�8S�}S0XJ�Xl�7 K7dL!�d�#$��暘ksd)x$�Z��!�ta��H&v���h�<n4���'����0-@>���۲ ���$a�'���P�n�#_���Se�}���'q�L+��S�>D�Ód��^>��a�'�HE��*Gu@�a�K�Pa�tz
�'F(<q�-Z���*W�P9Hn&I�	�'��LhuJ� �6p
�I�
@"v8�'l8�IRNH�(R��6�S8I��U)
�'�v�� ˭>Z�l�V��A޴�{�'�f�w+10RtS���
D�c�'���p�@n�I���s�Y"�'߮M��b_-b)��:����M�F�Q
�'�PA#�Z$��dI'%U$F�"-
�'!��"���� �̏�E�ġ��'�|-����P�Q%Q!��l��'��!
@�N�3ҡJ���'�� �E�"�#����Lp��'vd�b��?;Tℑ�/	
G�T��'7P�e͑7d)�q�V�MR���'|6�����$ ��3}4�a��'���Z�
Ja�LF�y�4�
�'�q�����]��� ��jx`	�'y��1��hWfI����&[�z�'�*�"F�'@,����LG�&�<�@�'�}��FKF�A����U�
�'7�x�ĝ�q�h��a
'<L9��+<O�e���S�4��T�@ 9�t�A"Od��F� /��l
��:�b�B"OI9��P�k:�Ɔ�+/;�t��"O\��6H��n�;1�]�}2�	b"O����-O/k8&�Bs�C n~���"O�h���/}�P�ԫT�L1���'9��ps���R¬���F/~Qp���D�s�<�!�:'�~��6玟?.$�C�q�<!�iUv|y�2/��Ey��q��k�<�R��%��L��$UD@�
及k�<� ~�1ǋ>XA�8"�%�!�ހ# "O���(��,�DF�!r��q*C"O�
��2T�E�S+������"Or0YS�Y�s� qDA$8�� "O��gMK�l/�b�b���rl��"O��AB�Z�PT���lI�-��| "Ol�8%��{��2G�i� ��"O�ڢ�ץ@������#cv��q�"OFt��k{�Z�!!� {tΠ2�"OBE���S\U*�A�o����"O������9���ᄉ�%li,#B"O�qģ� � 8B��K�7T��!�"O�x��q��@���!�R���"O̜S�f��Vq��˟��u	�"O�(�(��7����-��I��"O|�����[�|�%�߄��`6"O�U/��q! `Sqb�%��S0"O"0b�d�!m��� �9^��h��"O��JV!*��U`2��".�����"On��vfJ�M��9y�fB�i��1"�"O�,3.%
��e�% �t�h�"On����|1J�d8g�v�9�"O��03�S���lQ�H�E�5�v"O��(+��rO�`�\N�^��"O�L:!싮{�r!)�٦�+&D�2dG�uB�ɵ�\���Y��h'D�l�A≽E�ꈁ�ޖCd�P��&D������2T'$}�0i���ĩ2�-?D�����/�Fq����4W��1ȅ�2D�(:���:Wo�����E�kŭ5D��XW&�lF.(q�B��j}f�-D���uBY44n�L3E��/;��@�H,D� *`/�!}=�5�ٛ'��=��*D��������A;w1f���#'D������)�8Lz�iϩ(�F��$D�0�&�0H��刢 �*���"D��2� }^bXz���h��ബ"D���TL�f��:$�Ǿ*��"4A D�����#�9x��ڟfg()k��"D���v凄W��I����[^D<p�#<D����.�G��T�7ED�Fw�p��%D��kē��>i��`B�
d����o D�\�f��'�Z��q/�f�Ny�b�9D�Dzq��?BiD����&:�BR�5D�hA�#���	�)�'�ƍ�Ud5D���/Ґ<Ւh@b�9u��	 �$4D�0QPC�v�8�*f�F�C��mz�M0D�Xb���NC�H��!L���8D�:D�����C;��d��E�+n��J'L+D�PI�a\<lܨ�B� v_p����'D��s�ȅb*b�ps&2'�J���#D�L	b��7&���Z
'D,��6J>D�@��l��s�a�#<����<D�`�I�s$��`�c�(Kc�<�'D���`	��mPX�����(�Z�a֌*D�8���ȕ9�H#�F��:V�<D����^�RQ�C K7�̡�=D�$��`��b�mIcd�5۞Ѫ�#/D�+��,n��k�GE>�b�	1D�,`Q�2A��:u��)(K|]c-D���eG'b�0땏QrB)��C/D� t�.^�H�2���J�6�+D��[��T-��II��~��9)�%+D��R�H�	�vm����d����(D�� :1���L�����J-]���j�"O���4gJ�g����F)f�H0��"O�䀄%�	N�"����%!��b�"O 9�P��J6�Ԡ�9� h�"O�͐���?Q4���i���:��"O�\��⓹r,@	<IAP �0"O.��FhڨV^u�@��w�L%��"O�t;䊖%���[���1c�����"O���/��P�H���I#��hw"O��`���L��_�f!��C"O$�lG#6%@̚�ƒ�Ru0}S�"OX�c���t���!��Qmd�r"O@Ź$��j�b@zĕt3T{2"ONp���*��8��%^up]��"OX$rSϚ&U ���� �u�ɪ"O��h�HÆ	�ݨ��]�Cd�%��"O2��J �6��X� �حj9J��"O�b#
_t�d�+J�n(jU"O%:%H �v^���/A�~gFQ!P"O�x�g�5����ͲPR� #"O�$��%�A=ՓSb�!M-.�bc"O������+���v!��#(�lx3"O���EX�<(T���F6uPM+�"O=ꒀإXr�`1SI]��{�"O�IR���4�����ʬ	����`"Oʘ{d�E�����U�H ��"OҔp!��" ����֟,7|j�"OV%@�B�5	�H(�Rl�7�@�"Oز��zZ����jF�E
l�b"O�p3���zM�1!��6|�Y&"O�h��T�Gez8�7e�g��5"O�iC�
>ʀ�C��$�DM�"O(LJV#�-I�:u��G�x�aw"O���8��X��Fr�����"Op4򇎛�6��Aˏ����"O,�y��S8V=���!D��P���"O�Q��A�3~�T}���1Gt�x(�"O U�UME��� �Q4��
�"O����׃up� �c�]��l���"O�쩕(H�i�z��E�ة�Q"O�P� T��#�D�ح��"O���R�9p7�a�TX�w�H��"O&m�gO�n��8��̡k���"Oб�&h��] �Ӣ�� ��D��"O����U!'��:��l�K�"O]��a�}�޽��@�"�(�S'"O}5�q@@�*`*ԅ�T�"O(�)B'��I�(� )�
�a�"O׏��Xu��C�-Ţ�I�"O�L �kJ_x=i6���Z
P�q�"OTLx�)S�(p3�,�ZT�"O��z�hJ9��H�*ǍL��0�"O����\�>�(�)[�t�P�"O�I��7u���8�Ɂ�i��%!�"O�͒cĈr�
]�w'E8g��Q�a"OL���C�sk�����	�����"O\���"V�T�UhY%�����"O2�F��BY��aW\��0+�"O�x;��_��p����itn�@w"O�p@D`��s�fpi6O1up� PG"O��r��O����ɉ�fU`�y0"O�)���'WN���$��O��D"O��:Uĉ�7��{3IǕG:n���"O�Y�a���@���?(���"O� L9�!L�-J X�g���Ta"O��ycN�FN�a󐄔�VJڍ�"O�l�o�mp|�0&��+\�@�"O�8�7Ƙ�L��*�b�.����"O`@wH�� �x�rp�Ɯ��"O�l��Oϯg]hKQ���e"OfM�#΍�AdX�0!g� ZG��4"O��0���Tm`yJD��"~M��"O\���.Qژ��$�(��ݙ�"O�M�2gM�.A&� %����U{ "Oj)��e�6v�|Cv�Ĩ֞�B"O$ds��+W-�P��@��f͙C"OhX�
ȟ_{r`p�@���2�!"O2���� L��ܨ�e�/a�V��"O��+D�sP�ٺw��i_��"OԜ�j��Uz
F��}ґ��#?!��ձ,{�qa%O�&���j�/¿�!��/&���:b�h)8�8#���!򄗎8D��*�Lׇ�9@T�F:C�!�dY��J$!�B�,j�]�K�ws!�DC,���s@cZ�+���� m'yc!�Ý6���׆��ы�(_!��bŚx���/���k\�0/!򄐖|ڜ͑��ޅP%�T��j�$m�!�A���9�2Ʉ4")��I0�!���D^ d�(>zdhX�刀�{!���I|*9�I�,bc�eb�NX~e!�$��� X���ґO!�+C�^!��C:lª`s�"=5�ѩI�?Y!��8PM*"�o$FYH�ʉ

�!�d�@tzu+"��#y!z���iȋi7!�䂣�Fȳ����=�E��8!�$îg���A��[�z�!�@j�&R%!򄎗MFd���Kצ�
��f�y#!�$k���a7*  ���խ"!�؄{���Z��U��ڵ�n!�����izEiۂ� x "ο*�!�$lh=�d���(��1��T!�	{B�cBK�G�>9�5��u�!�d;_�t"�J����,�		m�!�B��t�Ӄ\�'؆�вg��!�$@;J���Sf������4�!��zV��U�H)U�<�x d�%f�!��ߥ� �BcYg�dE*b��3K�!�$�-6*9�����E�^mJ���8�!�	�o/�����Z%Ɣ�be �"�!�̘�^��w�;2�p���o��l�!�d;��8rqL�4�j�a���0I!��L�h�y�)@��L�Տ(:Y!�dr��0��1+�:!X#��?!�:����w�̰�J ���Ĭn"!�[tݮdB&Nэ-@�pC�G�5!�ӶtT�!a�k�=�-�#Q�!�d��3>v��U�̸i�깃��� �!�D\�SP�
4�ʆX��p��a4�!��9I�@�׵9ΦqQo<�!�$����O&Ǆ�xnթR�!�D���N8��MR.%΀J� ��W"O���`��XxL1D�3�i��"O�I�te���D�B��$\����"Of1�f�"lNH�06��.�����"O�qR5ԢM�q#�O6�:��4�'	�ہOT=R����7	�;!�D#VyzP��%��LA+%(Y]�!�� ���b�UѴ1�ffȴV� �{w"O��J$�I:g?}S�/v%��""O`Z��̊W�~�Pt���PM`�"O�q{bo��"��Q�W�	:La�"O&���Ŋ3.t�с��hT���6"O�u*B��MrV ɠl(UI"Oz ��l a�ڔ.:�X[F"O|쑤�� |j��
�c��)�p�"O�ٳr��$�*�1���:^Pb"O�-���Z֚	�Ń��|ؑ�"O4t�L	{P��`���)�v1�"O��ÆO ��p��B�
�$��lp�"Oz�j��
\�P��DKՂRxD���"O"�ag�{��9��I�vu�hx"Of� �Y��(�*BH�"��0�"O��@��Y'D��=�����	"O���7�k�/�3jV� "O������V���Y�¿G����"OJ�8q�IG,iZ��Ɏ*N����"O��+Ҧ&^[|�8T�ҥ+�V��"O\���.si̤�4� !��<xV"OH5b�!��A�r�JP8�S"O(��,T=���K�"��"O�$Ka�9sp`�)���)S�@-a�"O�ةC+YQ����ON�V	JH%"OTx� NX_��@�r�t)"O����´{�-*r�	�Eb��q�"O@��e�<,4U�X(%!`G3G�!����e`�-aAC��`�!��^:l��R�6@���"�O�!�$��by
=@�����kM�c�!��K�����%�Z��3!�
!���?%k4H�� �˚�'yx&]��3�x��$�ʄ0T�{B� �t����R ��Ɉ�c���p"�m�d���J�
DH���n��͓�H"4��:O�%Q"T�H�*m��c�)�N5�ȓ*�tD�"F({� �� �
���ȓc�bH����R.詗��C�F@��ly���Ѯ�).�ppɂb�c����`�2hu���T�4PYP��'li��a%��e�R���h[V!� ^�H���2i���`�.; �[�D=St��ȓ#�,�V�]�x�t�$���RB�	�2��E�&GR|Q(��V툏?�B�ɪ+��Pf�{ب(��0��C��5B  �C#;�`��EV�4�:B�I�����S �dpD�TN�^C䉿1����mT�Xt`��s��
C�I�A#X���V�I�:h�jM�]��B�I�yz���WAзIj�H��g���B�I�&�}�M	���VJ��*LhB䉻!قƠ��m�r�r�~B�I�4�4�(��7�6���]h�C�(o㢩y�F X4P��3�+-U�C�I+Q�);�D�4 �ny���-��C�� �|y�D�� Y+G��7Cy&B䉳|´��׮]�w���ȓ{*LB�	�&D����nO�?>v�HuE��Hp�B�	�Zkb̂ S�F�*�I�4�����,?!��҅SPe1�n�o���@c�]�<�TB�5� 	��ι�x�⪌V�<	�h9x��E��2)B>0Ic&�M�<�GG�-�������/$O24�+�M�<� �2���nް`r�� ����"OF�2�_�D�ʳIW.N�f\	�"O���&#�%�Ve�$���;��IF"OH� pBO\0\�[�,S�$��D��F�O�rq)�.�/v�Jdc�H"�'�1H�W�)��(�`�W�
��!�'-���� �*&4TTk��̸ �ݨ�'�$��,ٽ\�T���	ue>�R
�'��y04č%�L��7�ž~,P(�	�'h��D�*F�R�`f� ���k
�'�z0�'��2i>(�E��H ��'�!��O7\�"���@'`	�'� ��DF�6'���Pc[y�P��'%\�'�@'RuP�v��h��'(�[wD�c����8T�Z!�@$D�k����*�aB�N�F�Z�"D�L�V�/f�"-SvE�_`��q,"�OR�b�J%���K� ��Z寙(Q��C�l��E7"L����%Rg )�ȓ\����aE8d�
�r3�
��m��$����Z�\N��� �T�GO����֭��f��@�R҆{Q���!Ir�s	4C������X�^݇ȓzy(Iy I�F��M�W��@&ft��	ӟXϓ*���&ѻp_��4�֮c��� �:��R*¯]ܪ�L�$nLXX��X��9�d-(3H��$� }<4�ȓQWEzkP�4t�]#�T�7*�I��G:fI�F��]�6Y���Ϳ#��d�ȓY[f�����./��{�Π~N��ȓؐ1��5q;&�8��%��3�� �!�M�:[�D7RV��ȓ=��s2��33�*����q-�ԅȓN�b��o|aQj o��t�$�\�<��Ӎ�� x1�g.���M�<�厓.���Y(W����fM�<��ǉf�P �rD�0:�x!�F�T�<є
�1I0�rXQ�İ�o�v�!�ę�p�f�éUfVk���+5�!�$D�$W��k���(X��c��o�!�L�9�<M(��Si�L��D3u�!�D��X�Z���坔e=\QH�'
0V�!��	��0���UV+���5G�!k�!��R>����%FƦu���Ȑ�1!�$��kV�d�	���iG�N� !�DX�:���(gKX>t�����A��OH��ڼĢ�RS�G�||ĥ!�"O<�����N�V�{GL�-7q~U �"O`���|�I���<j �:�"OzD�џi��P@%.R�<aT"O^�0�L@����!	�:�)Cw"O��
5�@' Lv�9�ə4��1�"O�%9,O�>S�Xs!(�>^�V-B"O��!���T�
�c�e��#zѡ"O2IY�VL�*���$<�,,R"O�	���^�$��ϊ%lJ�8�"O�P�7��9h��5+��F6m��C"Ov�����k��@�f[��<��$"Oޥ�LN�i><ey���� B�mk�"O��ɤDZ	5�0Fd��4
(�
"O���i�������W�μ&e6���Z�D���	&,�L8�sjH6hz�p�ȓF؜���	C�F�c`L2	ul�����k#LV�[2,�+n�
���S�? &0��M$&)>�3팇%�TLa�"On���A��n"(�#��|�P0"O�����Pj6q�!�#aĜ�Ч"O���pdË\;v �v�\�>��@�a"O��S�"]�Sh,�Y3/�@�f݀"O|����;��S�_�Zզ\��"OJ��*-���#%��X"O����S�R��S˘-eT�Q"O�X����89d��V� �b"O�	��!ߨ	B�ma���a�e���&LO�	��H�b�>$0Fנf�#�"O8�1��[�MU�6�φ@��CQ"O$��ʏ�?.D�&��H�DS�"OB�`.���`���"�<�*O�9tK��?��A &j���'�,���&4G �*�a��X�'���3��ەkZE Δ�Z xz�'IheQ���%f$Щ�&Kb�d�'6�IH�-�O}R�C7BG�I{�D�
�'�f�Q㊁�d�d�I�!k{ll�	�'��XAd�W�J����dy2��	�'�p)�1�1r�\�����3�l��
�'�n��B\�v�L�$��c���k	�'rLA
0��*s����d�d�E!I>��k j$gM��M���Y��r����������h�%kN
_����H74�t@�O��8W���@F%{�zрu�Ir���Z=5�����%�V�K3�2D����� ژi2��˿�6P�R�.D�T*a̘��D���.h����U�-D�$9��F� c�г�� P����l+D���Ŧ$;��-��\�u��ra�*D�XI�ˑV�|y'�Q{��;� ;D�X�C��ਭ��W��5%'�$<�Ox���K�1+���a#'L� 8�"Op�a@��:\����q�5	�v��r"O�x[U��h7А�EH��¡�V"O�Q�b�]2��S���K�2�"OP\�$�Īg�պ'�S�x��P��"O^��gd0V3�5k�oχP��x�"Ol=1��[bp���مM~R� d"O�$�Ь��(M1 #Ýy���"Oh���L�; ص��c��PX���3"O
�("��	q>�j���l6�鲣"O�sTcC�~G�q�����_6�]�V�'xў"~�K�5b�$]��G/}pHM�҃���y���b�)y�n�u#n���>�y2�_:xx�Д 	�!�du�  ��ybe��nБ���߶/�D�g�ò�yR�M�+����'R!��)�&�D��y�$J�=����Ҭ� I���yҠ���X
�B��B��ð���yB.��L6�����:��4�Wh��y_*~S
����T�e��@�X-�y��ѥ	����6���^VD�h&�ȓ��O��D�O�c>�+��C�Uw0H;�j	�
�D��)D�t�ذ�Bp��ɇ?n��E��i'D�,0�N�#�&][���p9��*D�9�.ݺW��܊D�P���,R#*D��f�U	pSh��͹`�nd��:D��ѡ�Q�@M�%�?:��l��`<D��+�+Y�-ຘ1�!��V�%��Ո���k��=fK^��Q�;~-��8f"O�y	�j��Sߤ1�͖>/�N���"O� 6�����@���2�ýs�M:�"O�D eW����b��C��@��*LO @���5>Ҿ��P��W$�s"O�P�o�j�H��� �q`"O��ak�|�>Is�&��@n@���I��D��C�'v�4�*�DÐj؀��ƺ4�v���,E�My�*ĉHy<A0g^�U�d��Fخ�s3M����)�^D�Ņ�!vt\[ΉB��U)#�W�Y��p����E�)2^*��7 =;h؆ȓ#���l��N�Dc���teZ��ȓfoD��F�q�3�Dџ�l%�tF{����K
��ؓt-�^] 5"����yc��t�P�𠕾j��D� Ǹ�yr�	bzec�E�t6e�B��y��H��2�j�E˦O�t�s,@��y�(̀=�@tI�h�(E|�{����y��ԥm`N�@,��A�|iȢ�3�y���$�q�U*�33
��Q�Hֆ�ybeS).R��P�Ç/L<��g��y�Q�	pDK��ֱ!����b���y�ؾK}`���k_�D�`��$M��y�Ñ�q��萅�7a�fpK���y�k>@<\�� VS���K��y��"r'�1:W%OHF�������ybD#�V�h�ֱ>� ċ��н�y"���@���a��f��nW�X��'�䄣��춹�")�.m��h�'�C�.Ǣ6J�U�*�&g�D�!�'.�|����

2���>Vq�	b��$;��=���%;���y4"N<���X�"O��ɂ-۞	��
GN
k� �"O4	��œDf���;a��Pz@"O����`�{ኍ!�(�0o�N���"O0�`O_Xь�
��Y1Qоi"�"O�EytF��[h�-H��
>,^P:$"O�x�[�P�Ia�ؠ��:�"O2�I�]��]�4f�ָb"O4�XA���l�ZA�ߛ�n �2"O�X�Am�J�p`˓~�<S���~�O�rh�Fa�,$}�,;�LV�e*��	�'y�)��H�A�Z�P���
�Ό{�'}���"�H�%�t�Z�x�
�'���������ag����
�'0h��TJ�r�p8vdϜ{vtA	�'�8R����� ��",���'�Yg�O.hr�; ��e��' �D��L�hL�w�E�@̈Ő�'���
cbҟ7�v̂g@�K3rd[�'E
�JGV�!�������&x�~M��'P0YPP-;�1��;w�v�Cϓ�OT��$�"e��e��o	�̛�"OP%QQ�0J˪hB�ހn�Z}[�"OhM�B�M#��o�<X�R"O5���*`o�I��i'~��c"O����g��A�6}�◿/���`�"O�P�Ԋ\=oS�xg�Ɂ��� d"ON��)�Qk2+\�C@d#�"O�uP�a����tE�uqg"ON��AǃP)���k�`Xbm��"O�lkҠԵ��� GսvDb)�T"O�Ր�[�%�a�`f\:M~U��"Ov�a ��3 �A��F����B"O�����T�#yA���9�L�p�"O� ���g吅��\b�cޞ:��Y��G{���9T�k`�'�.��U�b!�1�������M���q,T�K�!�$�|�r)��	�dPm{�@G5!�K�#�Z�P��O�W��3KĊ�ȓtLRԚ`K�h���C��vV��ȓ+�
��d
нZ�nLp���&W�J�ȓ.��E�U��"�H�QSO(X�Ň�	�<	6�ݚ|���D��%΁�p͎}�<A�;Xc�(iD�L"�<Y�#�x�<�hJ�[2�H�R"<�HQ�2fx�L�I�<9a@�+$(J�cC#_�j!P bGx�<%��c2|p�㜊�l�)�Ŕo�<Y ��6�DT���?j�N���BZT�<q��-$mp�2i�E�Ѳ�U\���̓+8�As`LR//׀yѬӏEʮ��D�Mw�'U��ڄFͣ&�t�ȓ����դ��0����X�v9d|E��S�c&|9��A5GI��g�M�S*�B�ɑ�̴��'K?�>�X-Q�:}�B��z=�0)�Y�m.H��KDnNrB�ɉq{tDx�o͵'���` }�B䉲�<0@GF�G#����O3^%2�Oʢ=�}�b��6�ժ@��zd.��kHF�<��LP'n���RBB�� �d��~���Γ=Z���3�P�^�Tӣ���pY�i�ȓ1�ђ���:ʂ�����"8��ȓ
�x讬4~���+��i|\���"Oj��N�!�j�ҁ�V*mh���"O YqԣG���X9@�������"Ob��,%S1�\#è�~L~�0 "O����
��1? �9V��R;P�j "O�|J5� {��Rn��H2��8�"O.�)�-ƾ/�)k�M�
$�!ж"O��yW$<\�p�%lR�c!4�$"O���ZEc��j��94��ZS"O�tB�#,d\���@��$�i��"O�\{�E�)3�E�A����*\X�"O����-c̘)��
�u�4P#r"O�X��p;�U*w)�/ �����"O��eD�TUl[�B�c/.���"O��I0'� Q�
��v�^ Z���"O��:���E���Q��Nr��Kf��-�	L̓}��h�6 ��[�d0�u��xE�ȓ*��\��"��S2���KT��@��Ɠq+8p�U��KG�8�cMc+>��
�'�h��g+�P��|:5O
�2j���'e�xp��M�� *�-c�R�'4f{w!�-e����G<1�1�	�'�t��bBg���I",E:-|Ѝ9���'\4�B��MS��9���#4D��'6�81EK(:¸�w���Q����'�����B�%��#'�OJX��'R�!zB�Ќf�<{�͕�3�:�	�'Eva����7a������F�1����''h� �S),R�9��%ƺ���'W4p���נ!���4-֡K	�'�97�J.�6؁p�IY����'��ӷ��q�.LrWņ�	b�3	��'�`R慼5��MP�ڥ+�H�҈b�	B~B�4C�XŒd���A���IX��yB�3�� ��4>�Q% ��y��AO�b�c��[�&�f�3���-�yLJΘ�����lbJ���y
� ����������b!8��m�U"Oj�!1�b��tJ�ËI{�(�T"O�!��Z%�^�
pi�2�.$@�|��'���< 4I����~\�h!'�2!�d�Z� <��(�;eV4�@����c�!�Õ�t�i���`�D�B0�>C�!�d0N�d@��c�cM($	6H\�F{!��V�;nQ[�!�65�4ȥ	-c�r2O�A�':ȲR��9b�h-kf"O$�����9���A�Mĩ/�8���"O�4A%��k���Fky�q"Ǒ+W�דLof�0�f3	` �5"O�L�&�B�e_ȉ ��?`�����"O�m��BV.��EB�D�L���q"O�-9� M��$�I�1/���`"O���A:M=$Y�&�L(v���"O(�S����Q�>�8�F��.�T�3�"O���Ğ�V��Eb�B�.T��b"O���$�^&D�m01�C�-�l(�"OrIk�\3^����F�6T��}:q"Ov�Z�J�7-"�M�&���Y��	F>�8�Fy���"�L**��]:Q�&D�� /¹R@J���ρ%e�Y��D$���O���>�r�n�	r�$����6埶�yrE�1>u%�Xw��ȉ"�J��y�JI(_�2��e+Q4�@�Ao���y��,}YhͰ��X�Z��4���y�kEF���X��ם���3o�4�yG�6Jwč���y��������hO���$�-f�b�q&�ڎ~�V�{'�	3�ў���65�6D���
�+�-�PF	�%zC䉣G3�D�r�24�`a��F�Q�(C�	o-l����1m�2�B�׳"LB�	�w� �HZ�_�B�*�aՐ] C�I�O�8���T�!�:�g�(4�B�ɭ��,�(�\�*��5�OUp�=�
Ó���,t2��M�J�� iU CMyr�'�(���|�հ㬚5g�8����yb��5�<
gDM�7����O7�yb��vh�����X�� ����y�DȄAѪ�V$6N�R��G���y��׃ �X�uM�'x���6�̥�y����VyX��t�͂�MF�yb�w�UF�4"B֜�T��;{�=Y�ZP�9rS.&�aS�-W80���
B4-����ôA��I^"y��ȓ�dI9�d��@ܦY�pdC��3$��ہC�S���)�#�C�IP4ܔɃo����!2�_�<o�C�	1�z�PԀT�%@���	3(8e��L](�Rj�*�,��2
��cz�ȓU��W�f�*���E 
����Sq̠ �'T�V�h��]`�Ȇȓ������\�@X9�m��bp�ȓW��0�ă�J��� ȉn�T���:�Nћ�OM	PẂ�n�,hxG"��6Va��a�!*�r��3�^�)�vB�	�������)�$��@�w��C�	G�����HX��T�6n�/�BB�	���d)�O�xH�KIiB�	-gkt�#藤Iy.�����?�B�	�C�P�mJ�=�q��.^�#�B�Ia�	�J��9��1��]�czNB�	�l��qcĝ8���1�[34NB�)� .�`FN� �ҕ���
�����"O�=k��*���*����8`��'�1Od0a�m�+:�$��w��>^�8��2"Oh��Dƚ,�R�s��+x�|@W"O|L{�^"|О]��՞[>I�"O�ևV�]��	�% ₌�G��[�O>�����H�6���P��!?�����'���Ab��x�T�K�:L��e�
ϓ�O��ӥ
4>vI��˕�:�&�
��|r�'!N�P��)Pa0�*8]�2�S�'V��C@.W����c�XH��9�'H��n���|±E��9����w"O�TN�5M�����37��D6"O���Ά�bm� 2&�lp����p��y�d��,ZLl̲��sSx�Y�����hO�c���Où�5��-��T��I棧<9��$;打LNdc�͖2|Ȭ)#�<B�/����H�3-�R��󨜝;.B� �x�hr��&6�����Z�c,C�I 1�� J�&V)%Q�!i���	e7C�I�[�H����[$	/�ȓ��+�B�+���´לn�IBP&�(�B�J��Aר\�4��M���5`B�	9>Q�����#	��"�Ŏ�z�B�b@�q��H)z�ђ" 
4B�I�z6^hA����Y�2��'Q{8B�I.��D�0]��{O�,P$���$?��Ip�â�;(�2 !d_E�<�t�G)BHr4(��m��� L:T�f����I!aP;Y:�,��@9D��(��X�g@���LM�|��R�6D�8	R�o�
��	�	D0���5D�t9��D,v��X���|8��d3D�0�E/�L1�1hvA�5`�j��1D���v�\:�(s�LR�:X174D���0M��'��["br[D5�Ç1D��F���0�6�C��7d*4%A�*D��)�i»���2��D���b�*D�ā��L�jpxXd�D	ۼ��1�&D��P�X�e��(����t�vE�l8D��Yv�\��Ҥñ#�4����"D��K��4u=�4C�*��-�'!D�ȢU+Y w.U#+A2l�^�X l�O��=E��lЩX��0 %��>�Z��t(�&�OZ��dU96�������b��F��8�!���9��ċ	+��'/��!�d�==BY2�֎E�ZQ�$��!�Ғ80H}�V�Cn���3� CE�'�ў�y҄@	va:�
�S�r&ZxZk���y�M�V%)#��	u��� %�F��O�#~�#��aXf%�EI�@=�a��@Bb�<���.c�����x$�]B��Rs�<q�-Z*v��<�b�\)���R���m�<�RN�/`�@�B��ɤL�����e�<���J?�0��e&�ؼ�$\j�<y�ٞV��!ǅ�W�bub��[fy�'�V��CFQ7& �S�̵�v����C�(#��[��M�(���,,�!��V.�(;�T+(�5X��.i!�\29#�"�$�H<FDr�(��g�!�D;"�$���	OS�� �@.pI!�D�3oW����� .���SUJE�,6!�Ā<��a-�4N1h��¦�~!�dE^-�6aI14��&O�A!�� x['Q�P��u�`����a�6"Ozuh%��1:VQh���� F�)�r"Ot,�aJ�	xy:9P��;� B�"Or�#W�KF��ȐMϔk4�2"Oz|�fҖJ�z�	;_�@J$"O�}��X0hP�)�O]5'Id�Q"OJ���:V���`��\�o)~<Pe"O4!�1_m����?�����"O���珁-��TA&h����A"OV���܍W�j��7l�9YH$�"O@|brf�]ò|C+�lA*�Z�"O�3��
qo>��i[`�X�"Oz=Q�N�I#<�1����0�lp�"O���2c����@WHI���m�f�'�1ObA(E�٤ye�s�,G�q�XP�R�8E{���ό`9�Ċ[�䍁��"h�!���6�"C�;� �v�Z�}!�DP�|5��yPO�*�F��D�� |!��A�6���!Y��5��ER�.k!�d��&6��e�
4��37DO	!���l0�ĦR,peƥ�cb��'[B�C�'TQ
C��Y�U+E%�$֨H��	Vy��ɼCu��S�N�xNjT㱁�7�C�Ih=jh�'ޖf��5��U��C�	�M�1j��LBSV\�3g�O�xC�I�HUZ�YAU�D76�±'��	�B�5dl8��F�.f�1S�B�$ٜB�ɤ����C��,i���©^��O�=�}�u�_O�JM��B\��) 0��z�<����	A"���k��KS�s�<Q0�]#\Y�-	\J�l���Kq�<�u�	�HdKw�@+O������p�<��`Z�A����c�� -Q"�k�<�&3��Y�R�J	.J���aTSx��Dx"��9F�����6Q�P�ʊ���hOq���y��ڀ
���Sg�R���5K"O٘��ک �Ls�M��b�N葀"ObAj��W$pj�9�Ӄ`�i�V"O���CAM�BCXlҀR
$�̨j�"Ol����G�Qjl ����`�Ȓ"O�]�7�ϗ/�-;�D�d*謠s"Od�� �	�b�$`D$7b����!LO���&�W+���K��9~� "O���%���U�Hcd�Dz�"O�Б6H%I ����%]���P"Oļ�a��:r����өf=�ԛ�'����R�=]]lUeI֓���'���r���gu&�$�؂��@�'�P�kEM�r���V���l���Q�T��'���O5f��,ÑPRQ�˄m����O ����+���K�H1f�"�h�"O�׉�w������"T�"O�u��'��MP�����2L�b��w"O��g��sS���r�×�\�Q�"O�P#�Ģm)�H��oX8ڴ��"O��Z��8�p��T	X�Hx�f"O\���,K Z�r�Lɸ.���c����hD��-�M��ih"B�Y�l��5@�	�y��N�W�:�9��=_�I�D���y��[�zN�[F)�X,��!(��y�G�1B(�\�֡��S�8$�d�O��y�lY��T(�	�`�����&��y�FF3'CR�s��*Zl&��Fʉ1�?I�'?�E2#X'?g�ɫ��j �p���� -��i<9%f<�b��\;�"OF�����8�Τ�'�Z�j�)e"O��zU�C$Jh�"JL"Rt��"Ov9��N-
�<P�����g/z�su"O�u�fnЯ'3�m�F�G�\=nP�2"OD8q�ހ`;�U���Y/Y���W"O����Ǐ��4i �<U��"OZ��6mC�-]%�Ӏ�J� ���"O~��A�-�v��N}z=i�"O��ڃ��Fj8�K�0 �a��"O�E�aK fhx��A/�L�*LY�"O|M��ɩq�H�`'�}�<�"O0�R�ґW���@bm]�C($��A"O�4��'��v�|�,��%�eP�"OlY@�h@/~]�y���I�f����"O<�s��	*U���  ���w�^�`�"O�dAm�;���
Qb�$3n�Y��"O��y���>�:6�S,��݇ȓCל�����G�����C#~���}G�`�6A�=;�hْ�i1yN��Y�h�vDP,rـ�z7�U)���ȓGW 1&g��� k@TD�����L�bgT-��$P7��N�ȓl�LT��ʹkT�p�Ղ M`��ʓu����L�P�x��B$N�D8bB�I=(eȘ��gI%:4�X3j��ȀC�T͸XA'�?	�H����M�Z�C�I�zQ�}��͞r�D�W.H,��B�$N7��5��J��K�H��.��B�I�t��<��M6&��S�J	l~B䉸p���j�!��
U�� a߻J�C�I�&�@��LF��֐#  �7�0C�	5"C���� �/�Ҍ� c�FC�ɱix( ���1O;��؂���"��B�I�r����F�
]&Z�c��V�{RXC䉿f��	� d��i}�mC�_�N��B�ɠL�"�y!  �E�s��	��B�;Q��t�Ѡ:.�%xg�̩�C��s� �$�Ыh�r�KBK�-��B�	�x���kP'¬�b%pq�a��B��g�uQ�͚��P�@�.�lB��8.a<�Cp$�=M�К�	V�`<:B�I1bd�-P�VYfq��`�7+�C�ɭ!�z��n�#9lz�2a�Ň<�C�	�Wv�D�힛EzP��E�s��B�I�@�i�U(M$q</sa�*T�����Їp��isƕ�H���"Ol�ٕ��Q7\t���I�Kn�X#�"Ox���ܟ}9��o�?��y��"O��-�"f�Z��T�4��(��"OB�0ī�)����1��xJ|�T"O*�0���o���cm�#"�8)F"OL�K�N�.�uf�k�n�c"Ox�(!��8̊<��Q�{n�܊�"O|`[FK��Gܬ��G��/$|d�U"O�m@���2O8\���/�4]ځ"O�4ٶ���s��<S����H{
"O�	�v��j|�q�E�NETi�0"O(b(L:g�
e�P R(7.\�qu"O���҇V(:�a�䮔r�Y6"O\��w��W��Q&DM���a�"OD�#-�+�h���f�:�"O�lH�h����J#�K�l�`�"O8���E*G4�18�j�3&5�;"O� P�	�����=��-F$��i�"O���MTgpd��(A�'��4�4"Oܩ��Hǻ
��Y
�HX��i"O �a���6�F�����..x�K�"O�y��O���
����rN�Q"ObA`�=��"K����)"OR#g��{|�pu@�&E�<dc#"Od]@��?:|��/ߠw���Hb"O0}��9�\!kD�I�b\��"OJ�9����� �	Ϡ]��T�"O�\��f\5z:h�Di_�Y�-�p"O�P/VFE���E��l2y�"O���nP�>� d�Ōh��G"Oh��5ǀ2x���J߳,�R���"Oꍙ4�����M���L?�!�"OXyZ%g\;��BQP����"O��y1Cݣ3"6��E��B�R"O^$A%a�D�@&τmf(�"O�4;�c��g�S4MQ�4�"O4��c�>-�u���#�thja"O��,u��j2hǎ%*��E@�yR�Ķ�>�p�E&��<h����y� �,�^�-� ��ʤ�y��Ƹ>2y�l)Nvf�Ҏ��y�<?ݢ�3��?A����nG�y�˖�]@����Ǭ!͢�cj��y�)��:��}i��}�(�gĝ�yB�U+I��p��0b�hD��&�6�y�c��P�j�&)�Pա�F��y�·�0IF�"t/��,��E��y���,�а�@
�8��M^�y�*	q�0�r#��)Z�n!� خ�y2BʔO�"�:�H��Kй�����yr�֪\b�beoȊm�Iх�8�yRʲm�[Ř�UsX	���
��yr_�5K�z4A�(z�> ��D!�y��p�R�z끿-�CK3�y�*�>��9"#�}x��qǉ��y�EF>,8�xU�V+e�9�Ԣ ��y��I�*�2̸��φ��ᄫA	�ybc�V�y��H�I&NTU�H��y�F�hJ�%
pbHq:��4&T��y�)���h�B=A���pS���y� M{X���팊<�� [��3�yrE��`��G� ���@�����y�8��D� o	I�����o��y�c̲Bm(8���=5'<���Ó�ybś�b���I�!-�&AA���yb�ˀ /F��a��+����+	��y"�>7*h�P�U[<|p�E�	�y��	f�D�A�iZ��zyA���yB�[�Z����QK�6^�������y�.] Nc�h"f��~U��ZU��y����!R��{�+�f��d���yB-�/E
U	M%)NْD�)�y�H�p�PcV���`gN>�yB�-rȵ#�ˊ}��(�u�L��y���8�Z�!.|z�r�%��y"&�=M����g�	�lʎ���Jߴ�y�+��+�K�D�:�,,q5@ϡ�y�(�9�Bq���X� �
,��+��y�͐,8���!����PDX��y��Z�\s)�F�̼bgF�4�yc�xA���+BXʨQ����y
� �%���D�pS1K#��@���4"O�� �"�!HӜ9`g�I6G�� �"Oz�%���q�1��D`��+W"O�|��)O	:Y>�)��ۉGIvQ��"O�u�R+�_x~��0�V<EF���"O��ZbF
F�T����S��.H!�"O<�;S�$U���nŝE��h�"O�i@Q�R�W�ⵀ�À�Z���"O�:�n&�*H��B�0�~X"OL� @���m��ڲl����A"O�}�aͳ4e�1����	A��"O�q3�D�fZ�hsf �$d�n���"ObUc�5;��-@��`�L�"�"O���4�FE��[�&�;�"OD)C���T���0�"��.��ų�"O�͈Q�ݏ R�[�X�{P�"O�y����M�c��M�a�j�"O>!�$KV��H��g��_���u"O�����GI���m�"%����"Ob�!�
%4��j^4Z5k�"O�\:���y�(�b�JdB�"O�$���,[g�d�TǊ�pԎ�!�"O�d!��?H���r#��{���1"Od����I�Vn1�u石1��#"O$���=O���P�o7��B�"O ���Z�3���iEU��%"O
��P ɢkq���'��q<:�e"O@z��[�Z:F� ��<�Fu1#"O�R�bۮjL,5��%T��E"O��ZBC �m,�XB^By� !B"O0�����Y���!�3(B\3�"O>p�Sj�e�u��H�)�uR"O$�
fG�'�r0�Ҩ��4�0yX�"O�j�KF]�Q����	0}à"O�̢UI�)L}��'�
�&"��"O��Jq�M6��p��%S�����"O����C��-~� ��˃p�ܵX�"O~�)���ir5G�/P�FR�"O���Iȟ{�`9�%2_{�=��"OF��"K�`Yud�t�,�p"O��)����z>�!� -v|�9p�"O.��t�͒%`
k�Ę4�b���"O=ѥ���(׊DrF�:2� Ԃ�"O ْ���8X��7��m{�-��"O,���7\���ʲ]�1"O E��N�!W�)B#��'"O���5p.�Ȓge �w;T��"OH�6G��MZ�2�Ğ�X�D�CG�x·iO�b?y��>$��|J��nY�yZr�6D����eH�B��۠�D,BBtc6�Ix���81��11Z�)�l�	ﾡ+�#3D�t���Q�]wL k��ۀn�J�:g�+D���V2!�����*Q�NAAt<D��q���'�  �#H�(��L;D��eD�3[��P���mcޭ�tG?D�(���N�S�����'���hUN>D����'3,GmCq�Q��	��<?�
�e���o�7r+�
���=ޠ���@y��C4N}��R:!&j�$ G��y��=��ڵJ�-�bT4@��y2�W�m��s��N�~NM��kR��y2�E�TB��X%�J<�.ؙ���9�yT�S� ���X�~�p������y���/lʼ��kQ ���B�IR��y
� ���`��au����0\Lr"O��AL8��Xv�Q.q#��p"OJҷ�6��E�T%� �"O~ي�#��P�V��c�/["&["O�HR��uڬ;IսY���q"OH ��N�l��xT�>��a"O:��vm�(`�a�dY.G�Dh�B"O�	s3�Ƿ~�F!q�j �("Ov�� ��W˄�{%J�	�T)��ቻSQ��S�D��a��| �GܲG3�X�ȓ4��Y��D��a�x��,:!���n]�T��ꆠ4�D���I&F��8�ȓ�����KՓZ�f��0G�%K�pM�ȓ�Fl:G�,E����!���Iu(����i�	�a�4����N-&�ּ�r�O$HPC�I�]S\ej��͚N�a���3S�L��*^����-�,t�h�Q���& p����L�'���/��9���h&�S�����	�'�����Aی�肄U3|��҃T��26�>E��'Y���0���yx�FJ�@Z~)�'��`�yR���a&���r0@O*'
�pEzR��,�ȟ���1��4�N<�e�"��Sc"O���g�hju���\2s�FmȰ�Ot��>���i��I�@ B8tڰL�@�7&4az���Ñ���Zu'z^�� �P��'
���^�qYY���#��ܹ�̖�n���ȓK��89�$ʛ*HaY�#�-����ȓ)�𤌁3��%�w�7D�hŅ�	v�'��$��P�uA :����f	b!*
�'\!�/�h�pv̟"�(
�'̮ #�P�Zn� :�"�:�'�L嘴��2$��a�����˗��L���<a�홿>�����b_�5���mB��HO�ʓ�y�)��	1�䚧���/���呔�!��
Z�m� �ȫHN��ѣ�c��VV�D��M[��s��9P�!ܚB��d�T��1�lU�"O&��l���r���C�T����IxX�4��n��[��Ĉ�j
/��9��/+D�`�eL#)J(QAe��<UZ���O��=E�$!�=I�.�j&m�y�j�B�L�.NC!��B	:�|s0BM�����+ʥp.!�D�a�$ɳ3��(3d8���(&�Du�d�OR����|�7�
 @Lf#"��'?�@�G؟`����EyC	b? �m V)D�O� ���I!�
=Z�{lt3�f��;a~⁹>�A-	���i�GՖt���B&	F̓��=Is��&13�d"DcْFL�A��F�'s�?��������SSg� �e��d+D��p�$�{q�pEɭ��(��)D��A�bK�N���X�F�-~h��j�2D��#e'ֻ5� �w���g���i3D������^	�]��tAɧ*O�U�D�5Q��`���̑�P�d"�Ş��8#�L�ta
�I��^)N�l��$��)C�DX�K�Q��Oƣ]�$��>��(;<O޽�G�7?\9���#4��&�'ў"}:ش<��Q�v��5e�&�� Ls\dц�[Uj�F�&��,��\�}D��/(�Ex��	&l~a2��C{�<�V��4�����C��Wg�j���F�PP���"�'Qўb?�)p�ɷG��i��n�Ή�D�:�T#���i�s:�	aehF%�~e� 
�!�D� �8�9Rm�']~��w�9�!��9mj�AF�����c0nQF�!�� 6X���(a�2�PA�� Y�x��C"O.鐐*\($?�)���ɕE�yI"O��yE�yɧ!�d�V�@��x��'�����L��:-��q�iJj����?��'�B]�f�N�8�k�I_�=�NU��'B֭��A3��Jǧ.�T�ٌ� ��?�nZ�L=�oO 	lIa��J�_��B��=���k+75 A�a��"?���5ڧ\[v|*���^��q��P%U@����j�j-�V�0�$T�P���`3�Ș�'sў�}Jd"I(W�z@qA E
l�� NJ�<�a�V�U<���$L?5h$Q1$�j�<��y'&k%�S�d6��!|����'R�	!T����5 ��[`�q���h�nC�	�sd*бW*�&q�t�A �%+}~c��̓��'F�'�h��B	�&
I�(��ɞ1Or��Y��HOj�a��޲a�}�EϧS2�,0"O�R��P��ȐE!Y)r!8t[��I^���	 (�<�D߬n����_!��&����כ.:F���L�_�C�ɧ*2���'D�^�Ѓ ΐ-A��C��!6�v���ǧ��т��,?��#=�
Ǔz	��
H�4Yۚ-Y����LчȓPޙ2��1�q �mF�J���o�{(<��枧Fj�,�V��7 ��s���O�<���R� /��#�U+��
��O�<1'&C��*�C�%0�>���Cu�<��A�*!��#ȶb*���h�<��D�a������3.����f�<Q�o�U���0�fe�g��`�<���4�j��� U�$�z���nM���x��e�p�ytQ낰�s��+�p>iH�8␡Z$i_�P��$�0! XK�<��IE���dc�B"9�CW�J�<�gHr���!�G�q��I�2�Jb�<�&��<BG��� ���b�nXy��B�0X���5�+Sm�Y0�*�Ho�B�I*�n���/�.7�fl#����t�B�ɪu��@r#�Tc�x��f�..٤B��9]�
�� ���D�L����B�	�(�ɱ
�H�p�x�L=-�B�ɪZvj�Cޥ�J!#c�7!��B�	3@x6��C
��(]��.M�~28C�	#b���b��=G��� �K-8&C��"M �ĥG�D;��J:G>B䉄T&Hբ�'.4�u�L_�C䉈S��B��g9��x�+�P��C䉲!�h*���0N-�pPu���-��C��)wt�A�o{����a��s�~C�	�;p�@� ���'��x�&C䉝E�0X+v�A�f"v�L�4UC�I����έv�j|{5�[�˨B�xr��pr���2L@�#�;�B䉆z�Z=S7��6A�> zAʋ��RC�	�S��͛�
b���6f��Q�C�ɓU��i΍E�!�wL�"Cr�B��J�͑7@��wK���E��'!
�	�nW�xjp�(g���<���'��t���:���f%¼�r�p�'?t�P��QV)J�(��T�sX���'�za���K�rwPݚ`,�=l�����'�hL���=AZ(8��٭kc���'�(��V�L�]XX���r=X���'�� �@�/C&���A��x[�h���� j0h������LY��ǳ	֬���"O��i�� �n��眒d���˷"O%:��Z�Sh�¶H�� �0v"Oz�"�O�����s��U���*#�'����"�)A�b�i!K�
{��Ư����y����*6��'~)�@�A:�nM�`遾-9���'9���s�	W[�LɆ+^�ar�'�(a���B�}5>ԪӇ�Qg�0��'�`����%]�P�T!R�E2 ��'@BQ�  V�IB�dгL]�3� ���'��ݓt��P
��*�7)U��'�J���\.~0J�
�gۍ�̬�	�']�DE홥�1��E� cN	��'�p�;���#�h�C������'�r�S"�Ez��ՇM�x;��	�'�(ܲ�љ9����cԺz����	�'f�]�;D�]��j�%��Ձ�'ג�ؓ.O�%���*F�23r��'�D��j�-Y�EXcd�t!8�
�'ch03D�^�=d,�Re�زº�	�'�ހ�'F�1 iU	���fl��'vM����:u�|�Q��"�����'��-�@c
�{n����H�r�F4��',�ѐ��*^qd!#�ĆsS����'����C�T&&�Nh2��Ȩ��
�'���k�X�'��;BCZ�[`�(�	�'����f�$e���`�V����:�'��}�%��I�A��0ۆ4��'3��S�iW�m�j	� g�z���'L�h�m^ 4�8;���v�z���'0A�Ыʲ|�Ʃ�ц�'nH����'��\���Ӌn|��{�Xj(��'KP�Cb��M�̩���ل&���R�'9���r�^�o�h;�eÌ+�D��'�0�u ��(�L�կъ
<��'�NH�"J��_2�[�

��'S����d� L��/��w����
�'�ثfɘS�L�A) &j�콡
�'�lH�&nIL��D�3bL�d��`a�'�r<�f矼�����-��u��'{���eQq2�X3�ʂ�i����']����Q�z�����m�L��'��Lh3�\B6�#GaQ>y����'�t C���Nb�;&+,=���'H&̹s�A$˄��#� ��\0�'��'��2,�v0�vXJ�@c�'����1�ޜ4��@&�S�y�	��'U�]�e�Ɍ��X��[�{ߤ��'����ӊT�z�4�Av�_OҘ�;�'��c �*dc��r��L�_�$D�e"O�X�f��C��଒+I(��x�"O0����9��ae$VM� "O �����[�悫r �@r"O戰DC2v�`�Ӱǚ�HN@� "O�,S�(�)P���kH�,2�"O����؟~�\�g��5����"O���n޿w���"��
��X$:d"O$y��/�-O�������Tp��"O $�`b�%j�V=����,{
}B"O��ЈV@����#��]�<x�!"O�И�H�8�
������0!��"O�yaI�1��I�o�l��d�""O�	,���wT1��e�b��1v#!�d\_��0��.�Z��K'kJ!�� 0����,|�P�1���b��8[%P��R�z�a{��Ⱥq��[#� $v:3��p>��$�l*�N���3��*�&ARbg�!fB䉔arp��" �:�V����"�� �+����ŀ,!�}2��z�S�a�`YģQ�[%x�OD@�B䉳�����¸���	7��z��4c!.]O*��a�O�q�t�GL�����ͻW�`�W��QH$��c�5���ȓv�Z��g-Cg�Ԅ�3��04Z�P'j�.�<x@���8� �c˺c��4�����3�L�`7�˘vX8�V� \Oڅ�r��O�uc@bCL�^��'L��T� ���"�K0,��zȀq5�
�0>Y#I�^�8B5�ju�(Hd�@ܓ;\0��C�L�b|��Q+B%�`�3���x= 擦ٚh�R��7�r�#j�
B�I�D�&�`��U�Nq�ԇ�b��}p�H����e��Hw0TP6��G�"b>i0�N|��V!� �Rx�����?_r��u&D�˃��� :LHŐĂ�3;�!I�Y3�t�C�ՍJ& 	��!���1s���?E�P�] 
�=6X��C�@:����I(�����Gm��2�)h��c�}U��Rg�I�$������;$|����-wÒ�i�o;O�僡��Ɓ��
͡]/��x��$�_*��(u�ؽ$xͨ��\�m�� �"]�Vޘ���ѱ�Ԡ�f�3G�x��� �$9�/����	<��\��D���%bW�L8b����aȈ&+@��ꑍ#t�+Ɗ�<��|�r������8`��.كdT�� ��i�����$c�!�$ζJ���ғøl�c�+v��h�4(	+9��mږ�n\P��l�-ig�":,�]��LFEy������%#�b��Q�ԉU��1�0=a�)Q���t�Y�\��ɂt^�А�#hL��5�K(�$@�'*]3�nV�$Y�HE��mℝ��H�vA�X��.�1��'X&�:W"��T@[���:F"��OĆt8��Z�cNNP��a_��}���D�k�D�e���`�MV�N"EcG�W�`�d��(�
P�|m�t �6pf�96N˦
�,�]7[�*ش���]w��êOwÏ2 @bTy��3{�ɘ��QG<�VC�3F�v �Sǆz=$;�c@4A��K�퇓?z��ǳijf$���W����~:8kS�A7��䍸�R�$��^�0�j�b�72�џ|[ŃR�`Dt9�Jɋ~�´+�.�4G�N�p�+	�
����&O�撁#�ITOyB��>�H�[�'8�)G�s��9@��M���.OʥsǤ�3cW8e���j��b�]9w@
�؜��/m��tX��0i*`��&�=XB�	%T��@+'��b��g��!Hz�J�5p'�ə�:|iIq  �i��l�j������~݂��3+�S�f}��I�h����'6,R,�o�&@�IQ$>��8�!B %Ø]��h�M���L�(U���l���vk�+=�>�?�A�
���C�cڮ�����R LH\��d��~IJ@��Ǩ}�8��#$���xb/�6i����A��X���w�<��_bnv�r�_�i�����Z�4	�E &f6�S2/x�x�I�F�u
�GѦ0��B�I�b�rب`�ݜQ�n��C� �J��	���!�+�>K4�X`�-���I6
�	��ђ���7%�"	[TBT�0�`����	��Œ�J��f�!d�O�
&�I�!S�[�����-�G���0�ڕ<0��$Ԝ
��e+V<IÛ4g��x���Q
(Xh�diވ2Eg�#z����,�o[�UXu���<j!�WO�Q��mV(���s�`N(xGE��$^F�t�Y�	��\'��"��������T�}ST9Z��;)i!��;^W8�5	��}E��eZ�hࡳ�RT��ى'�^?Q���O� bP.i��\*	�S
���"O�$��F[�\�����H�DX4�(��'l�튕ϐ�:��D��SNX��pdŕ�#��V`'&���ю=|O$yJ҉������%U�b!R��T�Sq_j5(��T|�9�'�V���/�R�ڥ��/�c�Ht���d��,�v�����j��~B��3;j,�Ǭ��k�L���`�<�%��m�L���K*Osb<�ŏ��a[����
�ʲ��'����O.�Rҡ�i�H9@��`�~@k�"O\ !��f�Q�ء~���E��,�s
0A��-��ɒ>?�az�>Cލ�0H� &�b���I�YI����L�.�6Q��
:U��E�ϗ�y��i�����J��'�Ɂ���y�ɜ~�"��"���UQ<���c�y��~��$�e)
�D����&
?�y�M�*-���A��߼�25��I��y2��(6�d�`Z$�psN�,�y
� �< ���<��JA�/6�ep!"O`k��JЩ���("�q`d"OhDj��Lʪ���3����"Ojm���~�-w���CAfi"O(	��Y���'�ޮm�j�9��DW6W7���(��%�ġ�pH�I���+P�ه��(��1;KђO��CYнpt��?1�%��8����`F_7����v,��L�>tGB#�~b�`�O�q��	nx��#_,]o2<Y�J��?�BB�I�D���S�۪p��jv���r��ʓn��Ac�اS�ӧ(�p�����FD*�� �V�m�8mc�"O�8�ɑ(N�5�W�TC��&O���(; � hu�,����(쨉��ߴ\��\S�#�^n��)������;6*�,)�!�NM9A�Z<´��ɴ5&�� �M�3n��c�`���?��� 5kԐq�/��H >�t@3����R�� �H�g�!�d 6[x�d-ЌO`}*�`�)W��	�B5N�U���{��S�O�J[<ԭ�Q��d���J�''�đ%痞vuA�u$ipl$ Rb.}"�?!���x���{��A3W� EK�J��\�L�3���xA�U��_&u�V����K��ج"c�l��ԛ0K��Hs���Ԑx�����/O Źv�ʀҘ'��@�D��\�Бë�yJ<��
�'�����cǊUAּ�S(7z����'8e�Q��;z�Hu�2��$�|�{�'{��+$H�*1u4��1�R��!=m�Ѐ��'5���l��U��*�/���ă�'4���'�ӻ����*�0Sz<��G*F76����'ɜ}������0�͚+:�(�����+58$�� O��ħ*B<���ѭP��u��'O2{��ȓq��h�g���$В.g���'Bd��3 ʸxF�]�OQ>�h���h$�L�w��i�r�!��+D���%'�(�����fso^�$���I� �ʌH&	�F�3�	�膅�`�0��[׎��X���$A➍ؐ��7���
�)Y0iv���� ��i��F$���U` %7N��C��-@dX�G�j�����Ӯ�F�ӆvS��b�G�6�h�6D��ZD�C�I�T�8+a��K+(u A�Ϣt��Y"��t��=��ӧ(����c��ppzM gӤV>�p"O�ÕN�6�����~@�P�j�p�$��`�(����5����4�j��S��>b�t����*f�!�č�6�����$��> A�1j��\&<e�W	O�-JP��D��%��D��k��l��=2�T�%�x�ׯ ��<ajP�{��X���Ҙu�����_A�<��S B�xpS���]r�Ix�<�%ș�K�0�!"��J�/{�<�D���X2��H�F�vf��KSp�<!2�D��hl �j^5X$d�Ir�<�-.x�DP��O� �,*���i�<�3�^�ufn�����q�l$p'��<���Z�N!�@L]�a�	!�Jx�<�7��H�����\� lRe	�`�<a��V�\5l�K���sH2 ��*^�<�DT�B�-)`C�!4��zw�G�<���l>@%brl|h]b��JB�<	!�-Q��[?�I����t�<�P�حd7(9[�'GkT�Z��J�<)��܋���1��b3����UK�<�EL��
��:gc�=&&�Q�[^�<A�L�?xxIݵu�\��FF�<��f�Awd���KB05�d5�D��B�<��h�)$����T�2���`KE�<����i�< q�����D�}�<1���,B��S��ʍ_��ͪ VU�<� �t�Ԧ-�ܘUlU)k��1�"O�q�C�ˇY܈QEHT�'� tZ"OTЬ�.Kڥҳ)	��Af�CW�<��+R~��Ȑ	�9����4a�o�<Q��ʖ(kx�bg�@W�A@B��d�<Iĩ�:' �� �)>fJ�arF�K�<��N+{ex��g�1�D�[E�NA�<	RGp��b·Df�+�M�C�<�#F�.-I�G�49)�&{�<q����F03uĚ(_j<@Y�L@}�<��Jصq����gS�S�t��6��\�<q���H�MF�#਄�3Gs�<q����L)���r$0�9'k�j�<��k	9Ĝ�R[Ph���b�`�<�b����җ�	䔐#	�^�<aG��,o`�ʳ�S�
���aCS[�<a� U5Js,D�b��@\�0"&�O�<	Q΍;yp9���12P�qV��E�<���@�S�4x�����ig�y��\}�<ys��$t4p0�H��<)��cT�<a� wP{�哫两�7���<�ga�#s��I�dǛ!h -	���x�<aR��1`).��3�@�s2`Yp���2s��A�{U����'�~hҤ�ȓD�t��չJ|,���4>���ȓ6_0E A��p#,�vN��+�ЅȓO��$g_�V� ��P�F�J�a�ȓbތ��a�<c�ʭ@T�J1渆�$Yz谐�۫<
��#�AɊU�H�����$��(�L$8��s�,��Xs<�u�L�?�}�T���N���z%����3^���(Կ
�4��ȓo0u��e13�����#!��ȓ7 �� B���p�A�'�0{V�؅ȓ7�Z�vĜ%:�p�ኆj�~��ȓe 6\�0ˋ �j<�ժ߇<(<�ȓ!����R$�)&C�d0@BY�u#��@�q��ж,;���!�֓1?�8�ȓ|�b��A����R�fݑ/�����)��h��N�FV ���ȓNV�{�'жL`x�&�� #�L(����31�Q��la��<D�LA��_�.lȂ\(y���ٖ�լm����Y�px�AHU!`� ���Z���9�ȓf��@�,	��)��͋{�8t��<,]:� 	44הQ11��m��M�F�8��K��fX!W��^���ȓ5�H����X��cJ3�ȓ^�f�i�Ǣd=�@o���,(�ȓu�~��'�O����HƾmT���La��	EF�<Ms���1�M�5�x �ȓ\"J4*�$�JĢFP�HH1��[Bq;d��x��Zb�ϳ�T�ȓ_؄�u@7sn�<)�M�*oz���I�,�yRA��᠔"!<�Ly��8��9Ѥn��H�An���ȓ,>%���C?U,���"J�f>1�ȓQ˰�B@Ī�*��ŏ�C�a�ȓE�0� w$O�:��iY�%]9�-�ȓG���$	�6-0Ե��iR�] ��ȓn�<nܰp�4���m�a��!�'B��x�� &@��%���5"T�A�'�^e�qǘn�A�N�~��5�	�'3�����8�|�"P�D�zV�<c	��� uZRdNT�P��`͈�����r"O�����#��)BÌ�����&"O�� ��Z� ��a�,��b"O��ȖK��@N�e@�a�B6��"O�K#��j���SE 4lՁ�"O~�R��ޣWw��J1��R���#�"O�����&� Tr,Y;JZ:��'"O��j�b�L�\>N��;#�'R*����t����,���Xa��/%Ƽ�`��J	��C䉗��X��+�6�x�KT%�d;�c��[���f>�i��2"�P�dބH~\q��F,%_�C�I'k8P� ��l�>Iq�N��8�ij�f��p˓)�T���L�$0�OC5{Q�	I>�x�����x���Ps���w�[��<q�O�?���@�^�~�}�p�'�0�;��]�Dfz�HE�X1$��<R
ϓEct�(�EY2"��(B�'�2���h�A���"ό��'%�L��'j\h���b�΄�M>�k�d�ָ����%���}�լr���@� �ĉ�3"O2e"ׄ
Jc(�ZE���:|�u�R%tA�\���TR�!��
^���0z����3�Е��͔)?��Ņ�	9o�H��3�O�l���}�0|*@�"U���q%�'Y�9�'H¥0~(r���1U ���Ш��,2�c�p���!#�7c�O|���d�A�l�I�0c�=jTG�O؄T
F�5��lڱ�^�%�}h蕁q�j	a�N&��?!��Ż�8zW���J"2) %�+AP�� ͣv�A��ӃR.���ź�*�A����4A����HҮ쳖�̵)FH�&��`�<�t��}�t���nK�0��JD�K@��'��	���F�	M�@�T@��y�\�ph��lN�$�,O����D����ȉ"4�3c�'�jex�"���L���d�x#�bF"!� �G.v�0i6 �w}2��U3l�����s�'z(Q��	�77P��GO��%;B�ȉ{f�-|Ԁ3)�H*���H�|�4�GO�p�y�(�B���;�4}��2����I:q�$��J�SƐ[vHO'�l�sgJ���zy��卻f���a�*fݡ��)X�bT9cNY!�����ЃcO�B7���e�2y��zO�أA��/�MBf��A�NH��^�HJl���Q�Ai�	4JՃQP�9�TP�Z3 �!R����_��Q��8m�ܽ�DE8�z�`�"<��JᾝK���WZ���"�sy�p�d�:����gE���Y� �%B|t�`(OF��S���*�
���F��������  �2%��6��uY�(��1z_Ѐ��#� $��0���@�t��C�:�R�ȯI�Z@aeJ^�f[�ij7��o(<�wj��T{0��D�[���!�7g�|�8T{�ӸIH�m��i��|'?]Ҁ�q~�_�n���g^�C�$��ubG��?QF@߆hV�P�O��3D?L<ux&�Ċ!�L�a.ڪ<I�͓a$��0<��� X+��j��Sjh2d��o�'j� �D�di*|�a�Q�y��1P� !�����`*�d�d�,�"hƆ#�!�X���X�E��PJ�Xh1Ɯ@�	?�RY¡v~�1yff�?:�@���R�'���"o�{:��e`��%;(t��K���3 �Q?Z́�^-&[\,�	�>��!��B`��Z�c�S�Ae���'�2��2�� m�����U�&���'�6��R�S\o2	Ӱ��Y�ĨĎ �Y2�uf2��X�e	H�$��I�s���! �<�6�FA�4��dÄ�����K(��/{�r�x���D�b|�a)�vX�AѠ'$�����-Ivl��r��&��,8�.:�ɽ;@����i�0���j*�Ӿ�v�����$�kf��O��C�	%5��ڕ/X.bѠѨE��@JfE�#�[��B��Z��~��s!$���
�`T�QxN8��*#D� �SfR#N&q���,Tj "�O"%�a$��[r�`�!���<��p�z)#nд��3�8|OEñ	>��zA�֫MT�p�%19��k�1?�$�
	�'	r9�'$N)x����Iu�8�Y�����?��2ɞV��1�~��bS%|��a
sO�7�����+�q�<a���1�Ȕ�&��>g��cE2F�8��K��n��c^�"~�I0U��j�F��L�����؛h�B�I*��$��(ߘ,�h����/�1[2�����'��<�B-G	J�F=�b��Y ��kS�v��i�͋�$D�1��]p
H@n��~*��[d"O�eW�L�0Zj8� ��X(J "O� $5�I�t��5�J*�i{g"Ol�k������R,T�|,��#�"O̠ZPF�FN8�a�k
h�a��"O�*�K�*S����t�U"O��/�'d��<�W�P� 
�h"O"���,�.�ޑBN��&t*�"O�l�Pb"n>�$N@^�0�x�"O����N� :z��R�Q�B��"O�HK�͓pE,�1p�I�H�ĈB��Τp`@�ZÓP������F����#A\�
ڱ��R��+V��\�kƅ�;WT����
`��X`�K�*�	�![I�i�7b��B�:PDbf�oR*���H�Ӝr�X��꘎EKz����]B�C�ɀ;� ��W�ut4��l�]L�˓^����J��^~pӧ(�T����])b�a��Ð^�����"O�$�EBE&<�ccS�u �@����B���'{����K'����L
5��c�:LQɓ[�Z��@@Z�h�#Hm��ճ�����@�s�j������<�C�$�/)�`ȺsD�>~>�?���M�:���q�.�IA���p�IY<���c��E�)!���4
���k=�����Y$"z�ɯC�D0Sہd��S�O� Qb%@W1���Z���"7$:�1�'R�I�p�LE+1B��4U��%>}B"�+*n�����{�Hݭ^Na�rlر|^�}2���x��,\�Z�	��q�Xݰ��k�)��Ŝa���i��~�� �d³Ir8� � �p<q B��$c������zL#"b!/'�U9Ջ D�x�v�ʹW<T���W 0��ݩ�C!D��a.�/?�����IG>�9�f?D���'��*Z,��ՋF���%ڃ�9�{��Q��'-��[ �I����D�ͱA*�|@�',��s`f���u{��P�:�6!*e��Wc|)���'}�y���<%���s��\��y�����i���o�8��'}IL!Z�'[�q,�8�C��tkء�ȓ���"��[�A��`c����';��'�n^`�OQ>i{wG��~[Ɣ�4*�w@&���9D�Ui�Qd���CQ�de@4��
���	"|�ް O�U�35U���ڐ%��(ڲ F�	ކ��$�"6�C�<b��! A@�bH@ʱl�=˾�3�����P�K�W� �:��	D�D΃�+�FUS0JHJⓥ �l��" Y��y�t��K�B�n���!�#dV���*�ؼʓ��y�Ҥ��?Dҧ(���9���'P*��Tz{�xP"O�47L��!��}��i� 6Uf��6,	S��S�j�����8���1j����e%� �(��#�ӳ9�!�ğ1h���b�(�2v�r��M)OD��a�,t� ���
���W�ĳ;ψ ��E�}��xR����8�<�'.E�:�b�)#��"i�x�<�����Y���QMn��4d�w�<yR��%w�e�)��y��%�k�p�<I1IY^ax�:�h�9/ּ`b�TW�<�S Ԃ%�ف:.j�Qs�RF�<Q�� �&}�l�RJR�T;>���`�}�<	�N#r�R��%��0S�x�#�y�<!c�V[|�D
w�C&jj�}I�D�y�<��F�x6D�K3eբz09�+�r�< g	����@Q�x �#m�<����+B�ܡ&Ù$ȴ#�g�o�<Q�:���(%�Q�/�f�b��e�<頪ˆ�ѐ޽A�1���Pe�<1Q�A3w�2��R	[2xW8��R��d�<�3.͝�m�uo�/8��}2�%SH�<a�	�"��l���_�Ӥ��s,�@�<�BN��4�>����ٹ,�
��^[�<�  �v�<f@�+DmQ���1 "O�Dف��<�rI�D�T�x��a@U"O�����d��h�����zt`�"O�]2��eJ^�0C��]!,�	�"O��À��G�����+"xtH "O00�ъݨ�~EF�=	4�LS�"O~��DѿЬ9i������"O��+�AS2�����F��'"O����ѤY3(`Yc��3z��Y�`"O�IUG=,4���#&�U�#�"OHX���d@=�$�1�P�W"O�T���Ks��hb� s����'L*����Q�e`5��E�hjp�BAB�RKr��׎��/<��)
�'��I�5�U�'�b������2m���'~:`���~`d1W�A�;�n 3�'О��V�R">��rs��, B���'�>|����){R��Y"JX�f%�' x�a�;/�`���K\�M;q��'�@���7_i��t�شE����'U�-qjr���q���S� ��� ^����CMk�H���nY�9����;��d�^�qÒ���=&�)�T}���/<������$�0 ֤F�x����J�{�B���<E�d�шa���
��_E�0ģ�U�r����O*@��˓T ���	�RR��B��6F~��8�.~Q!r$�>���!&�c>�%?M�%Ø�B���6�K,6>������]3�I6Y\`��1%ިT\a� E7[^�&�[�5'l�Ȱ,@:��@�A߈�1q�e ɧ�O����MI��J� �%@����O�Fꘘ���H��A�[@F�,ȶ�4E��h�=O���7|`��$�8z�Db�J�&�f1�ȓ�T�c�c�!`u�&H���̄�(��6aY:w㙈�.��ȓRd��.jv��2�̀G_���ȓ�<pZ�GJ��C#��4�9��VR����-�B�AV�6<z���6L�="�F�1MK�ـ�'в&P|�ȓR��t�cA�<܀I�0�JM-f��|p$�2W-Q�͡�� QT��ȓ_��Ď� �,1�E	��9�@�ȓuN �UJ��{�rA���Ŀs���ȓ=����VŦ�5�������B���fN�!M"f���I�J�X�ȓ4'����b�0*�;��*a!�ȓ6�JH ��}Vd���&�.P�ҡ��Uվ@2�`��a�XmKF��?9.<��ȓ���R��Ap�͘e I"� ŅȓT�#Wߡ%�`�8u)_�8��ȓp���H-'�b��,�-I���ȓ.@��G���:��SŃxW*��ȓX]k7�9�"��������3��"!�&h���k2n����P��}:hXHF�2ĉ�T6���ȓMT��go�+\lႵ��\��ȓ�	R�@@�\_�I�`�;sAd��ȓ6K�j��B?  ՂT�ݠd,
i�ȓ����ڡl��M[2�Cnb���ȓ+�h	�����3��]���ݴdغ��ȓME`�p���'������>[�	�ȓ"' @��],j���ڂd��A�����I�:�s�gE�*t���B�շ}+����m�\h�@�[Є�jq��U�pŅȓx�H�1IݡIE��3� B�g�"���'�D����B�[v]顦A�<�ЩW�jH �a��@A1F�@z�<A&�R1>x�QeI�*��  �FN�<� �񁖫��e�*C��A)b||P�"ON1 ���T��
���$��"O��"�C�38J� S�+M>L�4��"O��Z�
V�| �M��tD!�"O�8�R��Ty-T�i����"Oٙ2��']~I�K�82@���Q"O|��Bf|��
�(x)���"O��c�L"
�����ȓ*k �
�"OXhX�%��>:��B�E�p$"O|�b�O�bL( �`�=N`�"OB`��Ϗ
$3��ڲ-��k����"OZ4�5�
7��9*gF�:`���"O�Ȁ��E�0�B�#��,x~!b"OX����
H�ns5d_�V�X��"O���QJ�0��q0�@ "O�Ba���R�qcC� Ll�Ay�"O��[��b�D50��� `v (�&"OX�3�@�(�H�S#ܾ���@"O�Y��ܖ���[��ƽ:��� "O|�����L@$��0gj��T"O(�B��u��5FlI��u"O�qQ�䀆t*�H�J�~0\%��"O"li��É21�gݏ1���q"O�)S�&�+OP�e�G�ϛ@���"O`���"C3����2%��2V"O,��`�<o\,qe�<v4Js2"O���fҢJA@�9Ů�4q�d�K�"O�I�efa��Q�~:�iQfeΐd�!��7bu�2g˔a�B��Ę�9�!�d��l�D��� �DP����]!�E��l=��ھ/��AY� 3�!�$-��2Ϗ.�����Q"0�!�$I�(~(ת�602�"���>X�!�DQ69�j%�B�M*�fa���j!��,qL~�i�k�m�L kA�0f,!�G�S+�5���V0٬L!"ꂭW�!򤛩,M�=�f
�t�p]���!�
B��IX�˄�T�-����!�D�e<�a��� �P��߼1�!����(K�CAX蔩2�F��=�!���,��]D�d蒷�_�}�!�ď!c���D!��V�9#�v!�Ы|��y�b�3l��8�d���Cp!��	�Uir���nG�s��qzw+$QW!�Q���:t�O�w�XPq$ҁ!�!�dJ D��Y�����@#]�!�DUt TX��kZ3#2��!R
X9�!�ſ}آ�bd�ϰ@��}��ɡ)^!�$�%)s� {Ä��{{2*�h�6S!��Ԋ��` ��ޯjr���  Q!��L)
1�A=k楫��!A!�_>8Z|�	�!QH�I���a`!�K�./��� A�&�V��/�!�Ջ��Q�R�t���0b[�&u!�έn�8X�P/�4�(�H� �Pk!�$ۖJx�+.�d<����N!��b���3�x41����Sb!�d�G/�U(�lY;t&��#�O+cL!򄅕�İ�b�����_:>!�dT<u�mx�I�;:xTj�.2!�d
5d��+p�\~��X")�)�!��6k��`��fS<�uː�[�v~!�d��d�I���|(�AHH!���L�6���_��qt��<!�� �|��Z4V�� ��5b;l�Xc"O��p�#nBx�6�3k	��b�"Ov�[d��'������S�@	���c"O"��#,Z3+��CM���u �"O�u�Q�U55Ɖ�R���_���r�"O� £cU�(\!�c�	�9$l��"OM�ۆ'�@��`G�J�b���"O��������~�D`T"O
$���Z07�~܃��K�a}*��"O~�I$Ś7�p ��d=�p��"O�0�.�� �����W|x�6"O��ؠo�:��؈���^Q�]�"O@Y�'�y�v�ɐ$� R(��"O� * E��B#P2��ϛ"����t"O����'P� 4�gl�0�����"Ox�C@̈́,tu�q������ "O����-�)}����d�0r��	s"O����� [E��%O:wm���1"O�P�2A�I¨Di��ԋc\�:�"O�X��(<�\XrG��$Aʔ:"O��8�b����AD� '���"O�H�.(kjd�{���n�y+�"ObCNB�P��!�`҄�v"O4-2��(��4IY��J�"O�%���4���@OO�K�^��s"O���3�A�y�L��o��՘�"O
��'�p����_�w��!�"O}���:"���	�Q[r�Y�"O��ʚ3{�1�����B%	 "Or��U-�� �x*voZ�%�J�W"O���i�"�T��K).�|�v"O�$�îZ�����"a�IЌ���"O�E���)=�����Pђ�16"O�Q+@p�� �c�ˬ=о��"O��Sa��)Ϣ�e���=�ȵ�"Oz���I�EƲ����NE4� �"O������>@p^�����0A`%{s"OTY����i&
ݡu�)
)p�(�"O�h�`F^)��a	�^�l�""O��q&l�5K�X�8HB�I���Q6"O��R�^�4"�A�t���"OD�5̕�X�(�*��R1=p
i@�"O���o�7_��1��嚺PuAV"O<��q�Ga�}���Vr���"O��#Ӯ������L�9�)�t"O�ȳ%)�7+��1�fI�:���"O�`u��5L<0ѡ�
.���`�"O *��K" X�A��%"�,+$"OJ����#�h����2/P�(Z0"O���WA�
6�l#FHϸ1�ɗ"O��/K�#�h�1@���5SR"O�S�G�v���13�[83
  ��"O�2Q�U<+�a�8	��j�"O�eۂ[��F���N��9����"O�z-^�h���F�E�`��r"O����IuKx���G��-��;E"OV�gڷ^�zQSW��G����"O<���-�,-8q"E�Ȉx>i�2"O�q�C-�8=��m
�gJ�e����"OZ���$N�ll���'��1�*OȹbP�� DV<��B�3���9�'�����ҪMB�3"�&H xIB
�',�	D��*
?Q��C
�'Q�GO'�4`$,G8oY���� ���Ѡ~#z�q�����yxB"O����.x�9SӉƨ�RdzF"O�q�5n�<��É�%^}�$i�"O���]+?<�eF���G"O`P���KǄ���k��d��"OP�0��\J=�3吜nnY��"Oi�F�1u�r���c�&e��P�"OnͲ� �g�� y͔,H��a�"O줉r�N�X��f)��j��xK3"O�xP"�&}%�!�"�3���b"O�!���ߞLO|X�/��s�FU�S"O�-��A�
x5��O�}<d���"O�T�'+g%����*xڌ4nt�<��K�A��Sf�.�B�)�j�V�<�F�8�D��1aO �ڣK�T�<��d��ݓk*�hks$IM�<���q���]�2�P�b"��}�<9aJ)U�(s�W�0�:k��p�<���N�Dy`pi
PCH�Z0�Q�<�.[?2���Y���=�F����N�<Ic
A�S��`Q�ȯ0�xt��J�<����8H{J���³w����o�<rۧV��*2��D�2%C��Fn�<a6	��a�%+g�F��g�h�<Q�
��Kڬ��7�0_� �}�<I7 �SV�l���
�,\�m�s�|�<��J�`CbYhE��� ��;p)�{�<��	r��-�����u(��:3bc�<ѵ��|�t��V�Xm" �	c�<�6�G�FF�9��/a��(����H�<�'R�橘�@[�{��ic�{�<YSJ˔D}0�����7?PX!'�s�<	��"?����V&A3�g NI�<`AY9E_�	��Nşt�hH9F�<�ׅW�~��̳6�Փ|1�)�KAB�<I���&6�4i�F!E�e�j�z�<!3H�	! �`�fR�I��q�-L�<��$���(����j�0��w)NA�<ɱ�W���(9�.�m:z��ʆt�<A@��)���6lT:���0 l�o�<�`��:g�D�\�RYbу�(�d�<	U/�4 0  �P   G	  !  �  5  �&  [/  �5  �;  ;B  ~H  �N  U  ][  �a  �g  )n  lt  �z  h�   `� u�	����Zv)C�'ll\�0�Ez+⟈m��>���ɪ�l�D��'O�����o] �P4�ѠO����N��H'�tP�l��BY4��D��<L�;`f�K�'G�d��'TD
��a}��`��U�	Re��/LZ�ҷ��*=�p�!j%e��KǷ��a�"��Z��D�E�F"0� �ՑrǦl*��)U���,j��ɣV�:�3Q��#-z����4m���1��?���?��a� h�a��73��Y���4"�&���?i!�i��P���I3`�P�	ß��ɟVznX��ܔ +�)
7�Z��4�����OR���B�����/j3���?���=��a�5������T�!��ʲ��#�jO�+x�4��,���	s�'���Õ�Y�͟ ��k\:3b��`�j"��:T�'���'2�'��Y�d$?�j��k�d s�	��yz@yÁ�Rןh��4Td��%�|��'��7��Ѧ���4j���'�f0\M� ��B �#;.�B�'�f9"jU
�yY�a�`�J=Z}��h�	J���Q�����rT�˘�Mt�iȐ7�����-#N0�PZ(VU�"n�-d,e`'�32O��$^�и��A�a��$[-,T���5n�(,l��M��iE�\*�D�&� �pe��I��Y�W��!|��`2�͍W�6������4R�b0ْC�+R�M�j��:�� �ܷ$�>�	&��U\�0 �i�� �}K��B�@� �еi847-æɠ Oe�FÃ�������[2��*g�҉0-f�%�Kɒ��ٴr�Q:eO��S:�����2w��Y�����',��zP�%>*��iri]�W
0�9G�'��O���>���N���>m@#®��!�0G�L�+�!���]�XL�TmЦx��zW�ǂ"O��g�
-���ЀJ�K��Y�"O<-�AH�E����Pg��2p2�"O2(+'R~t(��Œ�!�Pl�"O8���C[y(����k�8!br�	�qW��~���
�,�F��GH�-p�I��
e�<q�K�&3���cE�>4�T�(_a�<���E`h���E��(�Hr�<A�G1v�V��B�b��HSl�<aug?bf���ȏ@P"���Vk�<y�*��olZ�9'ṇ�N�� a��$1I*�S�Ov�T{%o�Q&���/q��=#�"O���p��1)\M���:M��q�$"O�����0�J��D���q�F"O<Hc��H�0���P�R�t;�"O���g*H�VDÕi�f���!"O��ƬWt���g[i���Z��*��(�O|��o��.���aDۦ[�z���"O��&� �l��A��&�Ԃg"O�TY��K3spЄ��Ϊ��|�T"O�I��]v�X�ϐ)w����"O�9��j��o�8��V
�p� �'b���Mvӈ�d��YI�#B
$�2UÒ/Z� ���Qy��'���'WB<� ��/��ɇ��! �\���3����'  =�K�Ɋ6Qxax"%;}ԜpB��1tVv�� �'�����@�O�"��DKY�u�*�	Ó���ɱ�M�]����4x�3A�$@e(�QiOےE�/OJ�!�)�'��P���!3(5�-?;e�������?!VVT7�8�iC$%�D@:@����&�:4BO�:�b>����$j� ]����Ļ+��"��IJ�<��k��c� 3Bв&�l0�F_�<	'jE�|���!�/&! ����\�<� X9Q�r��k��F�N����@_�<qү̎Qt�Ub��4p��t��]�<Yg���1�c�`R7*��-��!F៴㔎/�S�O�]
`OcR��, �*&��S"O,tQ�Y���w�L�a��)"O����ɚ�C��YV��;.��!"O��p�-D� H���ǂ��.�Y�"O�h�G��c�6yF��<+����&O%�_�m�E�_ ��l�S%��\��>O�����As���^�_�.y�D<s��1�tOr<�GB_;1k�EІ�+�%�<A!�_:1m�AP���-���cAb	�5�0Չ!�'x����}�䍱T)�!oָ5Ό�y~!�$H�j�N���C���}�`!#f�X�ɰ�MKN>y��ەb��ӟpC��G% ༕k�Ă�0��ݸATҟ�I[�,���ɟ��'(�T���F��d	�� ّG���� D��PC�H(X�#���N9p%@�)���lH�q�V&̻/�P�Ո]4j�Q��g˿H	)C� �M��+0ғ_����I���'�|��H�^�Y������K>����QA�� ���N�4!��ɍ�?1B�T��yY�h�/",N�	��Y����'�Е)��'�"�'��7�!�I�0�"��)ɲ41�U�g5�T�I�@X_$҈Ct/U� ����"&1~�'��	��1.*m��9B�BP/�p��I�ETV�X�B�z�Z�Х ��-��Ŭ�:�� (A�N�KȜ���&FƬ��d���!a��O���>ڧ�y�-&��ѡ"�?�vH�g4�y��{^m���5��-���Q���O�F���V6vs�k7D�_�d�A�5�?i��?i����X�	H��?)���?	��yw�ɆyV�j�Q;T9]��"C� ��L����a*eJV �8
@�4r����|���J32�C2�ۋ*�M`S�2 �l�'�"d�m�b��0�:�{����i���'xȥFP8	�d�S���u�`������G��b�'�ў��
ۋHr�)�I����L�h�V�<��?���Їi�v(<mR_Vy¬ ��|R����ę�6s�$���ֲB����	�"*��#��P(J���O��d�O����O���c>�ZR$�� ����N31�j� a��;�Jdy�l�5$�rpmR* E�  /-��Aԋ�2]�FH���K�>�!׬O�s�X���Y�3^����i�BeDzbJC�c�T,hUCˬb4S�ME>?�E����?����>�~�d�₪)�d��C��u.��ȓ8��\[G�7�PY�����%���ڴ�?�2�ݓ���Y�W���7�
K�x� ���y�HP:|4�d!��B.e�g)�%�ybA�������ˤ4P��7��*�y��) �����19�k�"�-�ybb�v���[�1�v8iFޝ�y�B,��!��. ɡu"�!�hO�xR��S� ��$���'.�L�[�� 0C��0(��d�V�Ҩf�����B�I�+WlΧX+%��CX
�JT�V�<��bT�u@E��W�W��b��[U�<�#�P/s0LJ�� ��bG�
v�<9��(Y*Px&D�(i'�i��L���peJ=�S�OثD�M��a�Yj)<��Ŧ�v�<��펎;��+�W�7H8���g�<Q�(�%@�) K�!9:��ӰFn�<Qtkޙ��)�l��\��r�mj�<�Tg��J���.?�&t
#E�c�<�ꊥD�8 *ƥ�k� ���+�`y�G�(�p>���ΦSd���#�3GM��Kf�<�@C3A�h  -L�&���V�<�'ギQ2�=;���%���I�I�<���%^��t�d��K��IuB�A�<���؜g��)����*e��+F|x��bĹ�0T�Z�4h�Ałf�@R6�=D����?*7�eZ��AoM�d#Ŏ?D���ぎ7�� s��@��`�Pm>D�x��S�>�d��eޒ?Mn�H7D��#�셢Xp���T��˖�x#k6D�\�ʞ�;jV*ԊM$t������6�$��|E�o
	M��<P�@�-X��H�$A��y�A�/N��T�s��0[�ҕ)ٸ�y�@����L�P�A�@6P�*Ea�y�]cH�{Ĥ1H_|���[��y�6��D�ç��B�f�:�,W��y�_�E�@)��!˪'����B ���?���Km�����p��	7h�@�kM�IL�ȹ�?D�d�.��p!���>Ԏ�!��?D�T��EUP�P�V8n�8�i=D�����9�=!f��CPP���;D�ܫ2"�GNnE�e$�+V�z���<D���`R�W�v���J7\:T�j'�<!"�Ud8���A��V_H�R¬�6}�>�RB8D�� 1�G&I��(5
\-����"O�H������D0��N;~��u8"O�]0i !ܺ\A�K41p �#�"O8QK,s��q�@ ]Rpѷ�'���*�'�4���ʜP�J����F��!��'����A�'��p��-@��,�'L�a[W�ɰv��-��L�(,�
�'p�����RG�%(wh��L��ĸ	�'�D��Nd�p�RG(��x���'�R�@$�U(��5 ���h��D9{FQ?�� �>� ����m�84��F3T�LٲAZT��rV�e*�]3"O�3 ��%5�&���Ɲ
��|K1"O.�r�&<\�`���/��a�ʀK�"O��ⴊ��PY夊�6��91"O�m�gaѕ8�}Y��_�M�>�Yv�'��ҏ��;���S���VuT����#cȅ�'Rӥ�S�9�<̙�:)Z@��F�
-1�b�Y���@K>.�$��F�����e�qy8�0P��#|�����y��ԋ�L�PC�	�J ��ȓk�x1�B_� ����%n� �=�'��m��2y¦劗�~�Xs��L|�ȓk�F8�!ډ��p�W6COX��"�^A�Fܮ3���w��3D�̄ȓ
l¥�E
����e�"��K�vh��m���E� S�@�U�1��1��ɬNx8�G:P� �ʇ3f��0��%0L��B�	��x��P����*��G7HC䉇J����5�8v:e�4��8] $C�I��PֆH�&rތ	g��n�C�I�C=L�dcX�\�l
�.B�ɹ9Jtx0���]Q<�C��{;��=��Qm�O��ۖM��2O��� T'%@�+���� TJ'�єh00�ɒ׼y�!�$\�.�*������Y1��W�w�!��YHPH�OB�"���[7���!�Y;K�P԰��_�I+��$fR�zs!�dW�Q��x9`i��*u �%��7\r�U(�O?�*gmM�E� ��B�(5�����x�<a�(��;���ϟ$�4Ad�CK�<�c/�"�ɧH�+Qօ(��X{�<I��ыV�z�ys� f�>���u�<I�@�	�k�S>��ѐ�RG�<A�i���)�J�6@�҅Xg�Dy"H��p>a��@�@|�����Ը`j�����B�<�� &x�V��R���f�ja3�UB�<!�e�1	G�թ@�/PKB� ��A�<y��Iv�x%`ȧJ��p��t�<��JZ�m��,���Ԣ9r1*ƏZwx���1`����'�	s �Iӊ|��)sR�?D���	�c�F�P��˾RĞ��� D�l��D)v�hX�I�$������>D�d1£Ãv�n�����S ~�D>D��a�	����Z��� z��v�:D�4�"a�7w��u���-^��� �7ړ!2P�G�4��=���x�E��JfV�Cw��;�y"���G��X�W���ID%�f�R��y�F��z�ա�dE�4�Ձ���yB��
%�Hb�/�X��`���y�]�'^�52��PX̤qw� �y�!�#�������0V╺6�2�?�u��C�����hծI�,��h�H0lp[2�0D�lC�K�r�4���I�e�y���0D�� �<��IR
}r�@増�z�~	w"O๢��+�t��vK�9��i�"O�y��#�Mh<Lq�ʉ�m�` �0"O�����# �i��wph r\�p{W !�O8��An	N.
-��(�W]�8��"O�T���u�`���W��\�D"O��� 'D�aj9��m
7"O^��ra����eh�Y��d{$"O�v�/�����ą���˥�'Eld0�'�H�S�N�*��e���V���x�'��`���L,nd�1�f����k�'�� FE��T��2�.��yrF))������G�Q����DҬ�y�� v����GH�CJܼ�S��y (dTD]��f[�f� �22�P3�hO*�s��S#l��򡚍��Ѐ�^��C��.	1�(1C-٧\R��2)��O��C�I��C�\6���q��7i C䉾w�p��Ǘ���`��}lBB�:/6ѻn�	�~|8��=W�&B�I	�����H֓[ގ��@X�Hz��D�Cp�"~*�E��e`CE `^�l�M��yBB�b��a�0΀�Z3��34�_��y�+�l�pu��#�L$"�1#َ�yB��;@��Z.�>���8bݦ�Py��6~m0�I�`�#A�X�:��N�<���\��0�J�ƨ��Yr��HTy��֨�p>��E�pX��Ũy�4�
ǯ�R�<1"'��hR����J�!=��B���Q�<	��Yw�"�Sb��4��a�kQN�<A�ʚ�)|�=��L��hPP��~�<��k�1~�U�2��;|Ϫ%�B,Fux��"�ù���D��+����eÛ�f�4`��6D�� �W�2���Ӄ0ZDx�1D������^�",��lI6s�慺tE/D����-׌Ed��R�e�v��!"D�	�U�	��d���?+,Dr�5D�L���̍va���iøE`�P[�K1ړ:��E�t��:u��e��E�%�v�Xe�
�y2��,=�f`�3��k�|��bF�"�y"��bQ�젱�L�f�*4Q��R�yRKmɖY��<bg܅f��y�'^�N05�$/��)fɋ��yB,@0r��ҷ6V�@�H��?�� �T������q! v����0��=�m�,)D��c��~�8�@�&Q�#j�1�'�(D�d#񢄭vp1 ���"E�P��%�'D��B�o�I}x5�d�@8�1���'D�,�ť	Ԧ��Pe�#la�%CTD%D�\84�����D�]5�T����<�@��~8�x�s�՞"<eQsF�b��\Ӵ�!D�|�#��.3ژ�"
E/���W�5D�D@QOxe��1�%  �E�7�y⣂�;".���N�4��8�$��yr�^�xi,4*p�\�C�&4GS���>�è�Q?��D-�>i�F��X�N|�6k�a�<)��I�fq�͐~��騅�NV�<��#�/K�Z��v`�������X�<�5n�c��� ��w���a�JR�<���t�!bI^
����t�@M�<A��*L����Aۚi�	P�,ZB�'�.�����)<:��A�_*d��
�@իX�!��@+L��a?.���@��J)�Xɂ"Of@Qo4NH1��Z'ttq�1"O� �Ŋ�cMr���n�o�4���"O}ц�ޜm�� ���TM��"O��)�n+<�|�(�n�=5��Yh��'(L9���::W&������8J�H��Ċ]��ȓ�H	#"#�%OL�\����QE��ȓ�8���B��)5�Ms���<x� ��h
�h�� �Z�d�0���>v"�ȓ<ƹ��I:;��Ie���/��8��͆� �ٕin�aBԍ�1|�|�'�XD�J�~�JWG'p ��B�9o�dA�ȓ!N�8��Qe�� 8ӣL�92��bqx�z�.�;�\m9% ̔�v�ȓ<�f$� !�W 	���3����9D\�B�݁g;Hi�����Q��I�mLN�	*����"�:� �r����s�C�I�lX �N��P�2az��<7<C�I�~�e�0ꊝp�0��5Z:(C䉍;��`����F1�q��9��B�	!юm�QK�%��r��K�
C�=E\*�{�[x�u1i^�+�B�=��h�O؆-Y�,���ױ~�"�(	�'>����m^9J�TY� �&t�&�i�'��!Ȋ�;�r�x�"D?>:
� �'�h|��B�a
���μj�D���'E�l���Դ��3��-2^=�'�݂Wă|8ڝ)���4"���8�Gx��	޹(��۱8�ā�ႃ<��C��p��+J'J����.«I�~C�	�F��{�eIk�<���jA�t�.B䉣c]<�ȣ 
ua���A/o[B�	�1H�:#�C�LVƠ	򯄩T?�C�	�`֔)�oC��LA�_��ZP�=�O�<�bA�����O瓅vg�`�1��B@�0F�ȭ`����e"��ON�d�A^1 5��RG�Q� 	�`o���r�ƀsD�с.��%Zu�D+j�#>��ȗ�G�ȅ��+tǼ!QF��-�ug`�Nh!Ap��/��EGD�O��Ez�'�?)�ΘOϦ`UZ�N�4��'�1p�0�)Od���-� �j݃�֩:MѦ?,�}⢮<�㑕=�jjg@\#Wrt���fCByA�.`�R�'\P>��@HW͟��	�de�d�Ў��ufهȖ��I�dy�IQ��cG�1CJԥ:�����ן�b>�!�'�9�(��� C�Q0�"@z�����_�v�ɑ��kx �����؊�$�ϝb�!��텚2��a�W%E+�y�."�?�������$��p��f�
8d�)��5;��P�4D����@�U�)���95.ړG��?@�"Y�a�~�����*�N��G֟(�Iߟ�a3�P�t�!�I͟<�	ݟ�S֟��Be�s�N4A��!m�ƍ�Ч_�8�u	l
z�����n�=]j!�O��O.���Z׎�ؗK�X}v�����t��!fkߗGն܋$��".������1�x®S	��Ţ�'˪S���A��3��d��U���'�ў(ϓmҖp8f'�z����R�'9�8�ȓR#&�`C�h$�m��J�%��Sןh��4� �d�<�E��}*r�4$�!Y��P��KˈR <Y
��i�2�'0B[�b>��O"W2���تo���sU�p�hC�,	)������<�CC�gT���B��xQ���>b�ؚ��ؕ2;�%P'O���<���ܟ�Hӆ��V�P��˜3C�u�F���D{B�	'VZ\���P��ĺ1�R�y?�C��A�yynQ(yz�����.OA��:^�V�'��ɢ^�������C���y�+ʡRę�VQ'|1���L�Iោ@"+M/6 �qJ�FG��{��|J�DH�q Ԑ
��>�����F�'9Nؠ�ȉ�e���"5��S3*R��@���ױz�#>-lT8�	Ɵ��|���!0H�f!�2 ��q�q��xy�'�B��G�<BX�"�V�����)e��DpLd�t'��m�����J1ê<����?i�����|���?1"D�"% *MB5�Ʌ�tB#/ӡ�?�E߹`�B�0�M����T򧈟�����16��Cp�>.���(�=O>����'X`�p��"�|�z7؁2Ͳ0:䝊`� �^���gYV��O��S�q~
� 
Ii'��vt�&��!k�x��"O p��'/c"\�w-���퉏�ȟ��ᤫ�({�
����MS��?Y���?�o��j�D���?)��?��'�?!���v'D-�%N٩u���P�Rb���Dԏj�JM��C�"�j͟d�8�,��[  QIf�0Z֮ 2JޫW��e�E%c��e�0�.�'�M�J;�D",y  �sQ�@��c�J�	�8�����O��=��'k�}B`@�#���
��ԑs����'����RX���KT�}�$���F���S�4�'Il���#T�b��A�Q �ȶ��@LB�'K�'J�)������"D�=�â\�ᱬA�leJ}A��;I:��ϓD
��j��P�E�@-��o� �̤0��M�E��\k7������8�F����	�I0����E�rZ�z�nK���Ie�'���p�H�>��]����IpT ��:D��+���:N���ȲiN�vMX@8pi�<E�irRS�,��g����i�O8� 8qD�ق:�:a���"<Y��D�3(���OJ���� B����(G�*���<+����ǀ�>@�S�*����">���YS~>���!O�J#����F�?�R)Ɯz͐� �჎G�s�d(�P) ��I�Ms���$H��f���J*�6h��@0���O���� f���"P	���j�MF,)0�}R��<Yv�S�4`}+����+���&�Wy��'��ꓘ�Ϙ'�N���':� !�cE�UB �Ó�hO����3r*�U±,_�m���r�DB���'江n��'��%-���׊�:�D(����!�'�@�L���<aV�]9r�q��ʑv�le�%�ݫ� ��O|��O:Ł6�>�����S.�j��$P�T1V���D��F%:�Oj����h��䀁]�N<y�%� o,Hg���y���u�> �>)��]i�s���ȬZq�� 8F���&��%�?�eg�N���K��?�2Ĉ�9Xc�����ʝ]�T��_���	8\b �'��'�.1@M�<۴e\|��,�BE[Ĩ�F��vy�����ɋ�ȟ�t���ʘF�p�;QK�:��H��l?a6v�T>�-W��?݄����A >�x\�A�_�za��Km�����G�~x�$�O��C0Oxb>����Ob��(`��EE��0Z�D�O��x�'+�,��O�s��"���B�KղL�u�ed�.s\����O^s������G/�`@�i>C�r��ozRI�-��Q��!��!��R��l�'��	F�)Γ�?QuĒ�=d<�:s�(�����(�;|��I۟��'�ў�	:�S�/^�L�p��(���dy��'��0�C4o��[���?[�=�ȓh�0��c|V|<�C�v*��<N��c�C6c6X�FO�Q'~4��R7|1�t�8e�$�9�������ȓa:�,��'�D��k^�S6*	�ȓ	8��`$bӀ}�<aw�}�pC�	-zx ���Z�E7� ���X�O1�C�I>B��A�@b�h}B(yShj�RC�Y'�@�JCVy ��`UU�C�	�3,Z!��&ڬsE*|`p��'dlbC��7p��a�G�ۀ�]/66C䉽2�PuKa� >�!�ӯ^cW��ЛQl�<xbڅ�&B�*s��&�ў�c�'_-G��4P���G�4�� L�@թJ�$L�����CG�=a�)k�R�Q��̩so�	Z���<4�RV�G�4�%9�ߣ,��a�`ꄧt��*c[���M*���͖����B^�(Ҋ���DŉK>�w9Yu`�eM�{����E��v�<�&�M*w�"T��#k���$^�C�I�x<��C�K� Y�#+ʎ=ҘC�I�kd ��c��`�����oI�3�~C䉚B2���YcF\�xc�pQC�	�oװ�8Cl�1v@-�%h�Q��C�I�<�Hi�IǗq�h�P�"��I�C�ِL����$�:)�a� X|.B�I �d��ۿL�@�X��*�B�%J�&�Cu��f ���L۲e, B�	"97�s�]N� 0r���C�	�&�Ρ��k#Z3���r�ۊ'�zC������s=@$Z �)3`�C�)� �X�a/��@L��J[r��y�"O���2�R�(��������Ez,�r"OH)*q%4HX��V cb]��"OlŲ�)�8��@B��;ybz �f"OD�H4,R�H��+! ŗ%��m20"O���!�	?/�Ȱ��:
�F�T"O��k���d����g��A"O.�J#̔'�pP�ǥ/��r"OF��s,��;}nP1�&C�2���@�"O"�@`�D��[2f9�� �"Of�`��Çk�"��֨)�R��"O��T�K+!� ���<0��H+5"O�Ay���s�xY��@�e�
��@"O<C��S�o~:L��M�!��m��"O��j�Ə;~��(�aO�0H��1�"O�����Il��R�nȃp��0��"O��H���5�4Ⱥ��8?�+	Gi�<��ҏ4]P\[q�½�FB؇�!�$
�cx\C�	{�k�~s ���"On��O\q��`Q:����
�'� �2��3-���j�1B���'vŹpƐc���w�C70`�"
�'@
�����J�~�b�	 -):�E��'%&| �aI?vF�	R�HD�	X�
�'�Ȍ�G`��^�����Ĉ8n�4���'PXᐉ�-���� 'id�:�'zF�����#It��@�ޜZJ�]��'3\�ݤY)�E��&ܵK���'D Y�$�2ZH��! �$<�@5*�'r�	����,E��4�� 76��x�'��d�֫8p�֨��� +0��i�	�'(V��@�""���f�"�.!��'f}���	T�(��n݃�^X�	�'�x18���G�jE������p��'G�c&��p�:�Pi��"�%k�'�fd�`��Da�öE��	x�'J�\ �k������A\7n���[
�'J0Y��*&�<R�슫Z��	�	�'��%Q�n�)��${�n��Mx8�*	�'�f���
M�8,��I(L�
�'"f|��N�]՞l �k�o��lc
�'1��"��9G�����d��a�\��'�����P�|x��P�� W	�[�'�Ԛ�� }��=J K�� ���'ʎ�2ǭ�=������,<p�)�'$�X)Q��6��8;��V�X���'�Uj�&�[�(��c!79���

�'YL��$�>Jx|!#��*�5�	�'R��[D��C��<#�cN�$D���
�'�a��ٳ7Gv*��G"w�Z�'�)��';P��3������	�	�'ٮ����=�Z!b���
5���
�'�(UN�n�^H���>X
�Z�'ed��$A�$�&��2�ѶI�!i�'_�Q۵fǗH�*a�R��	Q��@�';��)�@θA�``��$>D@`��'�N��q�F�n�z-s��:c�h{�'I(�Z5���Id.�+�O�6h)�z�'�:{�lg^�2P�a3r��'l��s�ؚ7T��B@
Ͼ*��l�	�'=�}�A��p���喉��:�'��zv��V	J`�ƌĀ\��'q�5Q�l��Z�@&��Wh��';da0��8�T����T������ �26���fș�䓀I0�Q�u"O
���=:��p`Մ6,Z1YV"O~$+�B;.:55��&��z�"O��� �	�����U%I�M�%"O� �
�5��t׭�K|���"OE���
 �srN-�
ȹ�"O&�����m�j��@N��v��4�1"O��j԰�@%:ס/�"E�1�I�<)�A#6\�5A�ҶO���yU*}�<a)�08渀�K��P2*�aq�`�<!��@3&��A���P���3�^�<�Pn�t����3� 8�q�\�<��8�Q�n�I��x�%!T��Bc@ҟ��DI��
$,� 03J8D�Q�j��7f��a�ۇO�\�)Pk*D���mF��f+�/o�XԻ@&,D�����M	T�Z�O|dQCE.D�08E�����T��2xLF�L*D��Sw�GG�@A@��6T�ԯ<D���@�]-\�!G�X�+s��9�%9D� iQ&�a	�gV�%���S�f+D�`2�N�	NiF�T(�扸��&D�Dj�%�#\]�{��P&0���B��$D��Cq�8W��ӵ	ЕOi�lSF� D��a��*j��V-�`ec)D�������1�~��fM�R���4�,D�,�6�*-1�X1LM�__z�S�%D�<�׮R�&� ̓l[� :G�(D���D��E�X�{fl
';~6Ȉ�3D�� ���#�;&�j@r��4D���E�_��;��8,8,�ZQ	 D�����6a$��aW�A2���b�D?D�ZѠX�'p�qjR� =L�IpQ�<D���A-�:�Y�0�+|@��!ac9D��nN�A7���U%ُ�f�Ӊ)D�x
�͎�!3��3�Nn�!�w%D�4�ӊ
`P�|Y�j5D���3�r�k7̓�M4h��C�.D�zA�Q':�d5��fR�
B!q +.D��ZC��1a��D�#T]23"D���,ޣ
��R䊀mA���w�%D�8����X����w&Ho��$��l%D��� ���+3&C��t�1D��4�D^�4]s�AݱT�f�`�",D��j��3[�����""S�-@U�*D��`�m�&����O2`I�]"e�4D�(a�
��5�1*�/@�f����D�$D��(�"��(��B#j4~��W�!D�4�$�Ɇ=������(R�@rwM*D��QQ�@?��1uG�!�%Ӆo-D���`�\�'��-���K�L���d�)D��C7h��&-f������t�A��(D�\�U���S���	��C7Dn)�'D��:�C͘~(n�ڡ�L�68����(D��Bd��>�9Q��H�>>œ�+D�8���H>G��[����8њ�)D���f�܎IT�1�
R�H'D�ؘg�GF0�S2�
41����&D���D�y�jP�U�p�扉��0D���Hu��[eL��S���S2D���׆��-TS��0;^��J�+1D��yL�P��%+$D݀��u3��1D��r NAI�fx��.�whxIb �;D�X bb�!
����Q��W�2Cu@:D�� ���Ե�d��9t2��t"O 9���'J����O�BQX��"O�:�Ƅ�1�Z��Ɂ�zH~hR�"Oވ��ԅQ�����";B�r�"O�����\��U(�F�-)�ᨠ"O���b��n��s������д"OL�bmC*y��܃$X��v8�e"Ovi돎"�yҴ�4R��Ljv"OX���ݸT�|) ���,y8@a�"O�P���&9�t		0�_"1���"O�k��eo���⏌�5|�,��"O�x�NȔ[y��� �eh|%�Q"O�t#NA=%���G�~�^�q�"O�$������(�m�%����D"Ob�[��s���
2�d �C"O,�6*�3-�i�v�'m�ƭu"O�X{0�V<}ስ/�Z�r���"O���۞8�b]���%�(�"ODz��L 0b(�U۠%��s"O�1�`�$�}Cp��}�"�(�"O&��a$��q����F�U|���YF"O:ɺ�I=b}Mɕ�/��	j&"OH�����H�IL�p�X�P�"Oܤ	b��1T~܁�2oU2h�i�T"O�3���3�`�p&)�6�2!a�"O�)ңp���&Ǐ�xX�9�"OJ�K���46�-XtK��j��X�!"O��P�[!A0��dk,���"O�!�3C7E�B�C
H/�ֽ8�"O)v��PԦ������K5"O,!Z#뎯gizL0�I�L
Xɰ�"ON�
��>쁻	_�t��W"O8�cH"Q����&S�wTUiw"O�}��*U�8����ӫ �3�zYs�"O�r"oM� Gd$թ\d<n0��"O�0h�M%7�N��F�'f�4�yG"O���%!A�=d
�Qc��'G���S�"O���l[�D�Z�A��Y��"O<D� I�3�$��@��[����S"Opyq��:S��5*�/]*xpD�T"O4�s�K�3��\)7�(f�	@"O��F�[�w� ��BJ>,ZN��"OD���΍[>8�����8b���"O� S��e[r�Ca
J���aQ"O!ia�ש{�Ό�Aҋ���"O`쪳,�^�He��ΐ|wx({�"OE���6�+e��cN8��"O�嚁a�����&�./4�4J�"O �ВlIr�m[p�ǟ3$q��"O(18�
�=��U�dƞ� �"O�Q�c��Va�p��C�_���P"O�X7Ɂ�U��1f/�����"O\��B�S� $е�?Uߐ�T"O$A�$�5t+�xY���=���BP"O��Y�'F� �&�U� ��ոd"O���9ټmE��D�Yْ"O����m�\y� 3�PI[�x������3���t�T�N������	��'4ꝰ#�)�P%��'D>
E����'\��񣪃w�x�DS�l�J`��'��t��D�,?R-p ,C?Y�^,a�'�,dB���2>�!���N�z��'K�qz�&�@�0��"	-B7*u��'��Y���ӒmN#�ez��'�����ŝ;:�6d���L��vL���� �˴,Y�d���7K�K�2�23"O�jdK̲Y��-�����W�dy@�"O��9��;� �4fԲm�R���"O���dAM+@��U���q�L-��"Or��/B6j>X8GX���	{�"O�8�R��Y͘e��Vb�L�V"O:L���
^:nAzЪىLV�"O�RS�Q�H{�������"Ox�CNޕa���b�R���"O2��viٛ;E��y0 ݛ.a8��A"O�=��a�k���b$�,Pr��d"O0=2!c�(}��I�˖:9Ѝ*�"O�y�bC�=��8�"J�m��D�"O���ՃˊI-bL�S��N� H�"O��R��@|�8�#f��V}3�"O
�� �ŝ3%�h�T+�G�L@k�"Ot(�� :X�H#�ܹj�H|8�"O�M��"w���T��%D�̂�BA:�Tl�+��4 �#D�<)���r)ؙD,�;"�� �RD;D�l��eQ:<����H91l�蚣D9D�����^	bb��3��^��Sf!D�c��G>�����f޷QҪĠT#"D��s�ķ@��l�S��$�n�G�!D�\��mB$#�`q�A��m�Di
�  D���F�t�Y窀�Z�<Qs�m/D��`6�d������#_t�%P�/D����o?��f=I��сD�7D����
�V+"h��"�C�ֵ�t;D��{�&�/TD�DI���tв�Zeb&D�p�`痘{�,�9s�ˊ�z��'#D����O�wC(%��	7Kl�M���/D�����%M͖�C�)V 6b�@�g�,D����E
t��G��J�-R�'%D��v�Sfڸڤ������D!D���d��v��c��6V��p��@<D����&���q���}��S#(:D�h�DO@64
*�Ȕ�t���k�&D��bE�$ t���f�n�00D���$ ��8�� �b�X$�N=D�̹kS-1���;�'I6pA�L�`D;D�d���A��� ������N�!�L�8�
,SA�bLVL���Y
M�!򤚂o��@Ʉ.Q��L8�	�z:!�$�(*hh1�=�P�
�&!�Dݎ7�J��'(���T@ ��-el!��B;9J�d��%\�g]�����1!��W�YV�r��ȻK��R��Ө1h!�\�n��a�J�����$K 4!�d��o4�U1���Z���Je��V%!��͜g�2��E�A�tI�0R#�!�dH��� .F�*��)�ȇ �!���=��a �G�|�ʖm�y�!�TH�[��
�8�:��S	8!�	0b�HB��A���C�s#!�r�洺�Ē�0�④U�֚|!�]"l�~0ꓩN=KvLq
�nUQK!�D;�n��@�E��Qpr���I�!����B��wE͕o9�pȟ !�Ƣ%W�z����2 8j$��8!��@4.L�5��3⁳㭌!�ė�=f\ئ	ښmxn� g헥`w!�d�ڮ[�,U�}�� �A,t!�dA38<έ��㜄k>BX��!�g	!�� �(8Ō�� �5C]�m����"O�Q�mH=jsha 1Qv�d�`"O�YT$)�܁$�B(2fr��"O" ��CN��(b� q}�0""O����eE�7.΁����Yo���w"O���@���=9��Аj���6"O��cŌ�>���A kޫ��|�6"O�x��苵a�мc��� �8�"O~h�+�/g/�����ݙ:��1�'"OND�6d�_ �2��ۚ&�N��w"O�� g���&x������.:�3"O���qLA�xs8}HB��"�� �*O��0 םY�<u��
+���'�n3R@\3N�dYӻ4 �z�'%R�$�����Q#@�R�e��'��B׀�$|��-�H ,�c	�'<,yR󮄹q9�`�P�Òt��К�'"�Ss��r�a�&��eA���'W�Mb�����5Q�OP�����'��Rc��������Q.N�:�'l�=�` M8;�|��K�56�$�2�'������|�PcD�r��'��:ƪZ����Í'�vL*�'��s��ܱt�@���b�?g���	�'(��l)!�4u�皝.E"(B	�'����mY9xtP���0)�����'k����)6T�GmߊW���S�'�-�ׁ\�<J���7��]���Z�'ߨt{7�*U���c���3V��$a�'�JP�o� ZeJ��GP����'�����8D��!-LI�|��'u�xcQ	�,��l�v
�|�z���'����Җ tTI e��m�+�'+� k9Y}Z�A�O?̌0��')��@�[�u劉�đP�Z�'��� 4+�"XS�jN�<4T�@	�'��!�W�ɫ/	0��<0ZXC�'؅c��U
Ui��(�� �<�5�	�'��8��M@��y�'J	f,�J
�'���J�"�`5.	2
S��'�85�$J#;��q�[��(��'G�}�AF�3S�
��#ޥ8���[�'٨y��
=u�8y����/"2����'���S	9���#]Mɔ�C�'�p��E��boR��c��1Z�h	
�'�Q;�*A
eBL��dJ�Th@�i�'�*(x��=kI�N�Im�L��'��"v�m
�u��u JM(�'J�ڧ���8v@�td@/="�9��'M��!'�\&%4���#'5�c�'_��^�=vu�vҍ0�4%#�']�g�I�J褡�N^�/(.��
�'KT\��N��V9Ό�a�-�@�
�'J�LA�MH�L�j�hC�%JI
�'�����������CF 0rp��'�5��cذF������6`��c	�'��R���n��d�T���jl2	�'�iq5��?��P%��;c=���'�D����qZ�#��=-N!��'�¬#5 F�T?v8!5���4�����'t,3WlS�P%
��O�,�Z�P
�'��5��2��s`�4^|��'��0�ƅ'��x��W�O�I�'= �W
w���Bǋ��N`* ���� pM��c:	
r���-��n��B"Oz��F��4<zr��'���!����"O
�ф̊6sD���G�MӸ���"O<a��$1�h�rw��|WA`"O$���7��!'�!@VȰ"O�۳�V�'/F���f��j�����"O��娏v@ ڄ�Y�F� ��"O��Cb �2�Qz���<P�XX�"Ob�35�ƅG�������'"O�5�����Ru�, t�X�qy���S"Oj�s��?d�i�E��t�
�"O�ػi�Xܠ;`DF�^d�Y!5"ON��L�>s6�K0+�;Nl	�"O����L�%���b��#�0�"O�L���At��%(��K�����"Or�YU�W>&]
�2'&K�1��0�"OB������a{@���!W�jD�"O��wl��'�d`q�-_</�Nq�"O49sč�9r��h#oW�+����"O��Dgҟ0�L0��@�*2w|�	"O�Q�c��5 �)�	��z���8�"O����h��K%6��pjU�Z�1"O5@4_
���1�	[(:���	F"O\�Q/I� i�$!�$���"O�(b�%ū
�*�cDo�s���q5"O~�CD�# m�D���.,d)ʓ"Oȭ22&O�EirsFOW;85"O�li�$Y,g��qPc�#d�p�"O, �ǈ3; �j��B�u|�8�"O�@ka/P�Ie��S��p�X�G"Of4�4gVb���"�ޑ9��"O01�g�,�cB���"O� ��J�9aF+5��0C"Oέ���V�2����N8&he"OVT�c O$!���@8u|1�G"O<����Uؘ�(���A�\��#"O蜨�c��:��|)%��*����"O����D�:�p��ʀ>-p�$"OV�S��_�a�ޑ��J��F�<�z�"O|�d��Z�JdrG�� N�����"O*�𥅒�g�h�CרNU�RMh1"O܉2�@Zw�Àȇ1<)H���"On$"���7;|���L��!�w"O�0"ql$zx�#Cl��	�r��"O�4��l�s]S��5�>��"O�E��J�u�)���W�E����"OL��B RH'dI$�5o�ơ(c"O��H����x�T���H�	Cw6U��"O��I��-`2�߰U7.�I�"Op"d�W!;F�Ab2���d*�q2�"O��R!U/[��w͐�g^X�"Ot���l�h�*"��	(�"O�U���ZM�Z���ha��"O�u)���gt|�`��+f��R�"O@aՃp�H�ߎ����1"O���B�Ƕy{X���G��( �cw"O���Q)7A��˶hN&#h��"O�h�M�8��S�� ,�ܱ�"O�q#���)h����
M>;'0�"O��w'��-6,�0�	�4)�JEx"O��kb^�l�4
��
�dBr��*�!��U�0��d
�Y0U��'��v	֠I��qB�ޒq��Y�
�'�	�N��*�0!�%�4\��9
�'鲹�s W�(LD��TGτF�L��S�? p0�%.��k6�ܳ�'V/�ּZ$"O�Z!+��\��y�'ٔ+ҖD��"O�����>>�I5fۢFà} a"O��q� >Jl���e�
�����"O������B���2"V��y��	6��V�k�f$zb��n::C�	�)�H��aC�3�l��E� .ZC�I?�HDpϚ�Q��c���V��B�<0M���oU�6��K�͚I]pC�������X��e�F!6T_,B�I��`e���g�LC7C�7vLBC�I<E&Q
����xD�P�"a��g��C��� �f��<F�L5{DoD�jgB䉍8����tk,B�C�F��C�ɉe<� �F_�}I�Ր��PiJ$C�ɍX4��9g���yΘ����(>�.B䉏kD�ř�lD�`�87�c�C�I�}��\�F�ξ%(���FÇ5V�C�	��fx3Dl �>������%C�C�	��6x ���G)��.�z�hC�I�}[����ؑh��x{��XB	�B�ɨn����/��\t�ф��ҴC�	>xJ^Ac6�K����l�,	1x,�����sMU�)y��0j	+*������1� !݌$(lx�K�JX����nɮ9)�Q�8��(�M%W[���#k�	��k��0�֙��
�$�$��6Ժ�UF]*Nn��tEK�x��ȓ\4�����]�@��F�Q݅�$j��֧��khn�s���ZtL���4e���J�e!0��*]!t����ȓ�� �Ф��P)����aV�
�*��t�"x���R:��iS�d�=�����?� ��&q��� �c��фȓ9�4D+W���u2�=�uE��[3���ȓ\lY����d�T	Z0� �4P��s�W%�%��ѱ���W��%�� ��B0	�z���)ej�e�����-H�ZC��^AZ����	�c�.0�ȓF���k��?��Pi7E��`cD$�ȓu&*YXBAQ�բY�I�",y��;�.9�W��0)k�B��K����>����FJ�s�B�p0���,��Z�DaX���D<>����N�|p����6�F���"п=��٢L��<4�ԇȓk�!J�	��@��P�I��L�ȓ�F�t��7J�9(�B��䨇�c�>)���֢9�Dų1�
B0��ȓQ��9�`)H�s�Fu�"^��.l���P�yf��#X�:KoF�8��h���XX������5��]�؅ȓ ��,���IQиq�J���8��ȓ0R���g�5���ѩӢ$�6���~����E��/ΞHHd�AZ���ȓ�耦�
�����*:@��Pž��h@ S8,�)�nM�hMN-�ȓ&�������iԂ��D�!�(���i��ؓ�gղ]t�(�@��>S&ȇ�\�J��o��`���S��p-|���L㔘x�[.��J��Z�+h6��ȓKی�i`(�;yDN�"�B�?��لȓ�2�Zo�j���;#�	�N�\��]��8���7yR�BIK�P��L��1���T�+`|8�t��2>6�ԇ�S�? �s���4Tb5��V�r�!�"O��r�Rk]Zs��T��x��"O�(p*�*~t���Ih�"O����[},5�%%��2��;s"O̛��.�lL��c®�:c�"OX�a� ��=���r&b�n�N#�"O�iW�G��R���E�Nm�X�F"O����V�\�F���
�
5
���"O�b�@��%�d�Z��8Q"O>,�$�ׯx
.��A#`ج�"O2qI��*	�TD�d�ʷHp(��"OtT���C�G;*a��V�-c��[t"Oܨa5!�.^4j��u�B,-��R"O�y���S�
Xh��J�k:� ��"O^<B4��/m{lX�D��^:p�"O�eq����L�7�	�8�Y��"O�m���_%p�z�
p,6���"O8-�F���ۆ��E�܏]���W"O�������� #s)\$gQ�e"OЉ�t�ä��So�S}�q��"O���E�.��<Z�HLgL���"O$��#)�&~Ҙ;&(�`��h 2"OJy:�a�|� �9�Gϰ*崄�4"O�xW �FbԠ[�fG*;�di&"O$�⥉ē��\HW�����ˤ"O`�����#B�.AhS��25��u�4"O� ��ض-j����R�E�"OQ�wdM�[z1٦k����R"O2��tfz6�iT�
e�>ݹ�"OzmiLA�$��� t��%K�eZ�"O���@ݷ,��ŏ�)*Шx��"O��HG�Fe��s�o9�����"O�y ��	o=��H�B�6��"O|4�Q��-��'�� q�r"O���
ޅ vT|a"��㰴�&"O6a�E"PM88�dկ]����"O���r&µ�]�q��!6��aS"O05���k6*w��v�n�;�"O��yV��N�⧬W`�.�A�"Oʤ�@�L�&ox�`b��] (��&"O��rD�Ӱ, ����]�0�"O8�␌�B��u�@(@�uc�"O�1#��:Q\��hB@/%ŰQ��"O�r"(ֿC��pS�H
.��å"O�e+���$s&�%�R�Q�7�x��"O��a��"#�:݋#�֙�@�+g"O0e:sE	T!8���,�<14Z�"Ol�'L �J%�i�
�[F��7"OJ,2�:u����)�Q�dYb"O��掏&0��A��Q���"O�5bBi�hvܒ�N�@���a"OJpZ�d�,I��䭐%�Ե��"O�� #Ü�P^�Q��H�_���"OX�;�-��]����'^g�� "OmzAG�%w �5���QM����"O�s#EH�vu�)�r�>8A�]��"ON����@l)X��45����"Od��Ǎ n� 4!���4�I"O�r�φ�~�ZA�ŭĦ\pv@��"O����Z
)Ǧ$� �8]��Y���'(��D��١+�e:Ŏ�- ���D*-D��SW�@4zZ(�B'�,�t�p��,D���q[4\0-��*9������ D��QIԮ$/�\;t.[�U@�%���2D�� ,�:��ÁRn�9�˕�L�H8{�"O�Ur��	�u嚠I�
ƻ���X�"O.-0�D�D�:5c�DL���0�"O
=�`����0)K�Ã �P ۥ"O�R�#S%��T��1"�6Z�"O* ��]�Ȟ��Y�x�V"OT$���G�Jl[���J�$ə�"Oy�0R�QI\�cb� �PL.D!��4�t!)��S)%b����G�@�!��$sP���1�ݷo��}i�,�/$!�dY�w\L�KJ�$�|q5��	�!�$V�^���dP2�>1�JX�'E!�D�Z�y����bE�Bi[!���%�z�iQ�MR�K�(U#�!�dջT:ƍ��ʦW��U
�Z2:$!�Ĝ�<oV��B��iK���G!�ď+_M�H��
C�$~���e�	�!�䋈F�("T��Xh��ЄJ�
�!�D�)6�x����?l�l:��Ӕm�!�d�> 0i���E�P��5gR W_!�d�9e�JX�C	F�!Jh-a��A�!��#4p��!@"\- ��P+��=�!�$F-o�=���Q�xҎ��G ^!��3K�lY�bE=i[j�p��eN!�Ԡc:�: �_.w�lh#6gP�h�!��Y�mpPe� O�/�=�w��k�!�D��՚c��:XD�� �Ԍq`!��S3nH�dJE���iIV)��$�'*�!���4#V�0�JΆs<ZH���;�!�$F$`d4� w)ZbC>P,|�
�'�d����n��C��̯L;�x �'�!�an�|�x�tRi�|i�'���Tm�^rLa�@�H�zm:
�'�t��	Q�B�xXP�I:�v���'���#�'�9K��j����+�6%��'h����号a���k����2Lh�'
��"�ŝ�v5ȷ���S	�'��&�0ٲW�$�np���yr`�\�ZH;P�͟%�@��ʟ��yb�Z06��e���� �����yB�Z|�0"	�4Z�R�J��y��B@�d<�b��M�Z���y���S��T�D䀎�
$�1��%�y�AD�[��YQ�߶jFDA�yrBŮz�Rh�%nU�^_�ó�Q�yb��w�R��Ԫ�Yy�lRì�y���(��\[�(��>�ĳs	,�y"� �P��1ś2;Q�= cBז�y"G�5�*��A��9����F��y��V���P�gˍ2�P�B�F��yb�F.Y�x��E₣#�K�$�y�*)��; Ր ��,B�f��y"$@���P��^�A,��v�R��y(�&5�� �Bȸ0<��%ۺ�y��s� ���o�p��őƄҩ�y�-mD��qsl�<d}����+�7�y�l��3Ffh�4�ܑ&7�������y�^2�BP�5%+�8akg���y2��1�r��ā�K����˖�yr�اZ
�p�F <K��1���y�K%���0j�H�Q!�ϵ�yRD�����)jW*G��%��y��E�q��Is+�=���`f�Q��yB�Ӡ,-��)�!Y�e��1WI��y
�  ,0��ܹ~���t�8u�9��"OU���)_�`@ۭL����u"O�)H��A�(d`���f�l�;$"O��3uG�R)��٦!� �	P"O�����F|@{򏔕Q�>��"Oa��� <��M�4q�(D+��i�<q6B��FakG�)0]�a�<�I�O�6Yp��A�N�y��u�<�Ӌ���+Dנ��n$/�B�?I���@R��X.��b��5�B䉪a�h����!�VE�)edC�tְA��n� "��+�+C�.C�I5M%^�iצ �s�~��᠂<�C�	� a�Y����W�&����Ld4�B�ɺ&�9 �Tdb�L�u/���zB��"ؐ=Hql�L����ކ��B䉥��Y1L���$#�m�{��B䉨8.D�q������۲
�3ZL�C�ɣRqt|���2�������&B�ɰq�� U퐓P���bhX4Q!�ڎu$� ��	�}��h���!�d�U� W���t�����!�Ğ�AK��+��(P�'%6*�!�� �v�[�E�R�(A����!�G��ʐ�+G��U2g�[��!�d�)����o0E~`)(bc�>N�!��϶'��}����;m�Qr!���!��]�G�Jek�)S��[Ҋ�	 �!���0S��Rt�t�*uF]Nv��'~s�gC���k$�F6E%��(�'I�8��hċ �^�Q�GZ�B2�h+�'0���.�n�Ȫ��Ƕ3��h�	�'����٬n������[�@=P	�'(����%#z
��WQ�	�'�>�j��Qڀ{EI����Q�'߀��1ɑ�lHT�t�G�(�V�0�'� �T�P2y@us��.�&���'� ������	����/�>�J�'����K�\������5��!��'�بJ�OX��Ic�V�6����'�Z #���� �� y@n��.H���'q����V�)����w��Z���'=�=x��Y����z�阻)����
�'��0�aU��d1p�I��#zT�r�'m�t��T>\R`�����q�'���Dɚic@ ����	q&P�'�%�I�8�9��@��5�	�'���[��H1���j�MP܍��'�d�BN��^���ա�y�J��'�2@�@�	
^|���ʬrn4ua	�'�^@�w�]2"����:�A�	�'R.3S�Q�,Uuj	69բ���'z�eP�ބQ `��/ҳ-B�ݒ�'(v�1�G��`NJ�2E��&F�X:�'[��KG��0&ry��D�+7��A�'��!�3,2�ڨ��`	(y>�d��'�4�!�2���h#�W��4�p�'�NQ���0SF�#s�F;��ͪ�'���"H�h�Q�� '�����'��0-�\���	NMQz1j�'��dr��U�.\ 	�S&E
HP�Z�'(�YQ-�?e�	P �S�F5Ш��'�8M�Ǝ�|=<��JI�(��p��'�>��ᫍ�r�.]�vMB�p��J
��� �ĉ!(S+0���rTm�\���@R"OS�&�@gf���
�FJ�@�"OP�s$k>?�H��ugz�����"O�M#!�	>r�H�2A�N�X�*p"OFu�U�]�j)����K�>��٪�"Oh�"�(�$ {!*�h� �Ѵ"O�2��׼|H]YJ�@B<b�"Oʴ��EX!O�F=A� +x˨�8�"O���a锲{K`����=�H�Jr"OXL��΍y�ڤL�+d���83"OD�󷇈9^K�A ��&AT��"O��#hÑa耸cTj�>���"On�ӁA�O>�*0�ʅN&r'"OΑj�M�ET	�N��,k�}�"O$T�n �s����lѮP�(�w"O̹��8Dƨ]�#nѹSڌIx�"O.0k5`�h@�ӭ�x�l�$"O���VJO�=F�B�-�*&t�J�"Ov��7�ę1���!�?V��-j"O��!���6�����ys���"O���#H¦X�!`_�y�d%Y�"O�	S�ÉN8B�f+[�,��!�!"O��S�#�Vi4��#�ʫm��	�"OP�(Ԭ l�� ��H�p����$"O�{0{��|�r��e��X:�"O�d1�	�[�]"��T%y�����"O�P@���1醥"���`3p}��"O�����801��0��g�Pd9&"OnP����Ԑ��PW�:PIE"O��BMU�������x�'�ސ�R�hl���ǟ�+��Q��'4�}�G.y�F�
5X�(L [�'U�E�AL��V0y��A4�ʄ�'�>��S@�;Wl�R�EN4���p�'KN�QI�D�����DF?�d�#�'v<�X�d�<1�]�č@��R�(�'��Y�@J�.��s���tz6y��'怭@�O�=K�1r�h����'�pأ'W�Z���	�����,�'y�+��?�N�9&�C� �޽k�'f� !���7*�h���@~Bֵ�
�':�����;A���z6��a�䨲�'�2�xc��>
|���n�T�|��
�'����iʭzh���E&@�	�'�t-�G�I�I��%����,r�'��bq��/O�8��a٥p��Q	�''|!�R�Ǔf�vH@��L�y!"t��'C젉eK
�x�x�GG�w�&���'_J�Q�*� رH	�eb�J�'�ȡ���ɿ"�v\��c�91�N%c
�'~���&
"PH���! ��.��'��9C¥4w?v��PD�%*O���'dx����'����V��<O} 9�
�'wN��E�^�.���Xv�_�?UҸ�
�'W� ���	q���@6���1�t`��'�H�ђ�ם<���H�/���b�'�6����\�>Rd��F!4'�2չ�'���#��ǻQ�8%p7�y�'�ڡ�cTT&��g��$`J��	�'N)�PgW�=jD�:�`��R�x�p�'��{�A�>����q�W����'����=�htr�K_�U��C�'�h=��
De�M!�����y�'5���q���z�3s ������y
� "q��'ǣH���r�>OW�i'"O|<Å�߉�P���E�7c���Р"On�#� YM�P3�د9��`3"OrD�'�!{\Đtl�1x�Լ�1"O�I�Dg�]�B��bF��M1*O`�c���q��$Ȣȇ�*vLQ�'�8�x����ԙ�c��l���)	�'�
��S%���
�Jj%\��'ub�ۤ�N�,T�g�9t~,��'�`|k0� �q.lu��!MkkX !�'��Ygh2.8P��'
_[|iA�'�*���3}Q��ꁣ��%^���'kH��@0}�����$�L�'Ƥ�S�S�v�b����gJj�*�'nj����6�rL���d���k�'*A���C�yW~���ͅ�U��$!�'��%�fCJ�%E�pkA��N��!��'Z()Eˀu�*����^�J�C�'��ZDnQ%Qz8ba�A�I0$	��'DBl���ΪH7�-8�&�E��P�'�@m	F^���� #�/o�޵!
�'Ȱp@��3�,��֩e|$1x	�'�VIxqa�2D|�1�gNX���	�'f�9c7���Ż��
a��`r�'�tuRs��*D��ub�I&T�> �'���!� *kh��i�	��Gجuc�'�Br	��´�x3��qfщ	�'�vXcr��8L]d��5���$���'C.��҆B�T*n�+%j��<��'}"�"R$ҥ"�0���N�,��A�'�ayv�"@&�@�'@��x9��'C����A.*�.D9��P���X��'����(�)Q`T��KٍP\*`p�'؜�9R�а7���T6P�h���'�٪�L7e�������,=�����'��P#���H).�u�_�4�ua�'2� aA� !:���*���-��'L"��ׁ�-�4 @�i���D�y���*| ��#�}��:��2�y"Mϧ�P$[$cX-iZ��V�ط�y�H��1G�J�{�j�a��]�yR�	q@l�-�v"T2�k��y�H#PU�mq��Z�us(P��)���y�H�+b��*d`Ưs
ؽ��$Ћ�y2�΁��u���ä7��ԓFo�>�y2�W�N@0Zu,�73 ������y��Vo�@bl��+мDSu�ŭ�y��!]��T�2&��7���#�K��y�E�%<�k�9/���EQ��yR��fg���r/؇S���k�.Վ�y��� t���3R$�M�ꝫ&CH��yi_�6�~�D��/�ƍ�֍�yB�U�]�-#�c�#-MH5��'�y��
j^d\�wÀ��t@�1��yrkS�z��T�q�Z(e ��	��y�"J�M!2�!0cǂ
H�ʁ˚��y�.+F�jaH��-��Maŉ+�y�	�_� ���"T��������y"�ݓ��S�.Q��4 �M�y��4+.A��(�]׆%��?�yҤI�7�Ԡ"��^�Gzi��ׅ�ybc�`�|�y�%�7�@�5�@��y҃�: < S��N�/��xU䑠�y��G�"�`m��(�* k���y
� ���Հ�#������=0�2"O�5։�{�J%�CCW�]7���"O�I��9]{�<�sa��+��pf"O�B&m;z
��F|n,J"O�ES���k1�a�� �(t��Z���՟�[�EА8ߛ��I��Y3b���EW[NK�F~	qO��$�+4E*��b�ЫDI�����5n�L:�Oj��r'�W.r� ;��J7>�%���d�����I� %\��ף[I�DR����#1V0�� ������vnG���Gz�ݑ�?q��_Z�O4�FM�5/xl+��X�ʈ�P��1g�H�D'��i�Ͽ;0e9,��#�I����qS��e8�8i�4G���i��;6bXC�ɻ�0���p�'�~���O��ī<�O��'>�4c"��Ox����N2����CH�\��a�E�j�@���:JT�����Ͽk��M������2�>���צ�P��цo޸(a���6�Bٳ���6s����\c�8��!CX~n6���1%ut���44d��I��Müi���s��D� �yT`ve�F;�(��O�D%�Oz�a��҂V�x���H�������O
�m��MCH~r3�]��u�o�He(UX�!�u�8J�I˰6�Pʓ��E2`�iYay�g�%H�n;`�[�} `�uB�j�����[� �^E��ϛXĴ��G��lYz���$+s��s�i]�"kD,"f����{1gE#�8�2�F��Rt���Y?��ǩ����'Y��)�
�N�l�#�/�x$�I˕��O�����OZ�O���Y�D�	Q}r#_�7����v��7t��q�>�y�c��\\���5�
e�l��棉� ;xr\f�l}�i>q�_yb+_<�����cj.}*3��$��P�"N`�R�'a"�'B�X��'E�'�tԠq�iऍ;R�7V��{%��hW y�dg�,I������Wf����$�����ۅ9B��I�hԫT�q3��= 6��"S�2��B�,CD`HFzc��?)ߴY<�Q��M����UZ��ʸ�.�W���'��I�8�?�OB��a��,
��|���[�f�4���2�����`0�A�Ь_�Ki�H!���0�(����MCB�i��Ba�H )��O}U��n��?j��pm�?K�iS&~rqO��䚫�Y���Qz��91�V+q�~I�O}yy��	y�}
�kG�k�H�Њ�$N	�t�$���9����5��5^PD��3N�KӚ�i��Y�l�0��0�*1.�uFz����?���0���')�S�W���J[Ha��Y>N&�<p�oL��?������,L��_�&�FD3��׾SU(��R�'h7�ԦAo��6PT�q�%b�(a��|�����':%Pc�OF��|z��?����MK烝�=G�3o�
Z�Q�ܷt/~�PCà!��)�g�� }�tdb�/�"��e��r��%F�Ԉ�O�U�
I�@�{�pt��-7�� L_:)z�� )�����\c��ę�_��3���?~R�B�48R���ܟ r�4�?ы��i��9����[��1ipDU�-��!��'J��'�ў���R�K ��XE!���S��+Q�	�M�Ӵi��'��ĺ��F`��-�� �1B�~��L�I}؞+
   ����0d"̍�I���p�{1��(�O,��O����˺+���?)Eb��X�"��31���Qr?٢�4�Of�q�и1ȠH��ݝ?L�� �O@	��n
�#ڼ?�1�'Õt~�������	���$���	�t��ґb����H(��,s�vB�I�b�(�0$�,؄�@�΀kV(щ��?	�'a�`�s�xӜS����C��i�`(؜SV�䉴��Op���O��dI>3��D�O�d:^���O���,�"���p�\�ydd��'z8!�.O؈��Eb�p��S��:5�,�u�'�ܔ����?ab�A�{"}�� �^��SU�g�<�rl�%=�ac&��*�h�]|�<!�PN	2e���Y��-���<I��$�)QֽoZ�$��W�T,[DFhY���36^})v�u�C��'���'w�M8�'L1O�S4)����N�	-�l����T�j���<�DLTm�O�ڌ��b��_1��C�?O�l����$Ʃo�R�S�fpT����ƻ7�LD��P�rB�	��p��^�u��#JԓO�H���Xb�I:?��9���"*+��Mܤ6BB�b�jw	�*k�ؙ��o�>B�)� ��k���1Xk��J19���;W"O�Q�#�P)MG
%��NV
B���	C"Ob� ��UW���sd�&\��kG"O�� TH�2l��	�IfVa�R"OBEa�剩b���#Ѹ�~�	@"O�d@��D'ԠK�-�&]r�x'"O��'
�*���y��Rl2�s%"O|�Em�!
�L�@�YK�<pr�"O�\SR���{vN��S6y2�"O6L l�@QT�;CG��-�1"O�����Z#Xꐚ@g��3P�"O�%L5$6h)�b�D%a �ٳ"OZ�auf�ƙѤ'���z"Ofu#S���i:
����'?x�3P"O�:TL�/e�X��e	 5�9�1"O�Q`��	2V6�����*/(n�`�"O���(Z�!"df.s(��4"O�U(D3`���(���(�U1t"OB-� �E ���Y�F Zp��"O�x0�ڛC��1B�@��Θr�"OxD!��+v�&m�:'�ԁ�"O�m�$�@.#�%p�,���y�"O��%$��s^��d��P��d�"O4�����sV���2(����"OƩS�+E�/F�"��w�JpA�"O��j�ݾn���`W2�B�j�"Ox���]f�{�!p>e�d"O��@&G�&t�0��]��C"O�kA ��x�&Zs�T<V2���"O�4�E�@����RcS-1��R"O�f$Z�+f�����,<um�#"O��h3MLhަ�9�!H2CktU��"O4�'E�T���K@�܌%k49�"O6�2p�����
g�.U���;"Oh@�h44Ђ�o�,bc%"O�rW��C�0�[�.�4g�x {5"Oy�s��!`>�P�]9�i�!"ONR�-~GX�q�L�� 3�"O:8#�HA���'�<b�>�d"O�} 'M���R���*�>;�>�d"O� �lܷ_���B�HKO�iD"O(��d�J�lD��G�T�\б�"OB�{�O^�I��c��k��(;1"OT����� p�D�&D��0��I�"O2H�w!�l_|P��"H�0j@�"O8@H�Ő|��r2aH�2�꽱�"O0�����~�DS�D+Da�:A"O��@bm�;$vT˗�ޤo!�*R"O��!H��
���H��Đa"O�1�V<��`�w脺�!�Fyr��1H�c��|7���{�X �⌍��;5nX�<�DCPh*t�!tBw�Ra�Љ�T�	s�BA�ϓZ�Ab�)�?w����U��25�zP��	�{R�a"�(���L�e���4�k3��#��x�Ѻ	r��bu����������O6���_�'! ���!�	U�"4X�L�~K��!Q�����~ �U��f�<qb|��'D�0�m2�)ʧ��%���L+���:G��h�H��ȓ-�<C�(�Tr��J'Z�~e�H$��
�[���<���t�d�����K�
x<���$$����@a��:k|Zw���k-nHbO�	4�R�F���u�;�p`@�"O��pM�@�
Lc1$L���tq�"OyK�j��D?0��b�(�| c"O� ��XqKעUVtm9AL�P�p�"O&ř`J�%vZ�2C�H�j���"p"O�){s���x$�:@�����8�"O�]�IL�2V������
�F �"O��� B��u�ʝ�㧂�
Rr1�"O��;��L�Y8��Ɖ 	nu�4"O��� �����6� H���"O�mC�-�>)~��p3�@�Ҁ�R"OʁA$D�Z�<}���[�H�8��0"O`� ��-�9H��N�u�DT�� 
.<��ɀ8�� zVj�1rF�E G�[3m������{�O�,���A�"�(�/�(7:J�2u"O�eڀo�<-��-�.R�^ ����$Y-B�⟒��%�g�C�ބ�n�<_(Ӄ"O�"��c���]2G��n�k�Jʣ|�')�����[�d��b�^m��' ���0JמJ�]ڴ���M��U����d���"H�B!e۩[��i8��Veq!�$M�I4�R-�1P���FY�!��?8&� ��.�4�Ԁ��f݋�!�SG�������W�XP�CLٟ^�!�$Ӳ8��Ŋ6��y^��gj\�%!�$��y�I��a���)��1!�D�+(�jՂ5垈zF8�i`遧#!�L�0�l���wH��u�!�L���"~��9i'�}�!򄆓̜��3S��Y����z�!�d@�6��\��`"������!�<����5s���)�!�$L==��PG�B	}��;AO�!* !�d^��dy6c˩�����F�!�dЮFl-�����*��!�>�!򤐀~�U�ТƐNj(�ЁI�@|!�d�+c(^��4$Glr�5p2ϱWu!���, 
�I�Aˎ	�P�z᎜%	a!��Q�?�Fxv-7}�ZuI��ʶ"T!�ę�WZ�Y !L�#5����@@�O�!�ĉ�E����n?z�^�)�� �!��7XHI��,��m}hȣ�ǆ`!��\�n2j�XGl	� d:6ս7�!�˱U46�h���- N���%6�!�$\�h��|p��4m�����1&i!�d�p%�5�̀qߪ��ƀ�*y!�D;�b�ɥ�ӏ"/�`Q�l�~!�Ă�La��J���O$X�Z�՘#�!��:cȝ[0$��&���G7I��y�$��"��Sr�<q7�N�F��@�Ȃ:�4q���v�<���܈2\���ЦC�|f�"��u�I�tv�bs狷�蟊���'�q�L
���	��8K%"Of�K���#�Xp{��̠9&�q�hW�`��O\�P!0�3}��r� �4i�/Kg�)2�i���xҎ��qS��8yxX){���A(q�A)5�^��+G����tK� ki|4�&�e�y�K�"oal�&�<���	h\����J�3���k�{�<Y3@ /an�ۗD�;�Hʳkv��?�h�3k�����s�EV�b ��.,[F0�E"O<��QΙ���cs�H�Z��uʒ=�OЕ�'�5�3}¡V�L��M_�m��� �6��xB�.E�@�# �O����FmI ���$��;
b���I�|�(\k� }�����W�,"��ti7��%\��D�'d�JP��9h��R/ SU,�
�'���s��U��m�0��3Z�H:����){~L47�?�J*dOL��y�ΟW쀜G�Q�t��X�I���y
� phY�[YD9�&L<iJ�� ���(P�p������Tڢ�����>K�!� �_j�<�7	�#��(���B�G�\��!<�=`����?�	��G�DI�$�-��)�Pe*D�ě���qy��+&����*V�	�6Mn�=s�̀2�BĬ;�0�3���k|�ӈ�$lqK��̖$j6��!\�:�-��Mj�4�F�7��Yf�U�K�H��L? �D�zW���%ƛv��2��',��>}1`!�Z�vF?���!�<_�n��T�!Ky>�b�ʘ�s�ӧu���3���SB��	5M�ۅ˟ c�zp��0����p<�t��k����N\�xFDI3�C��~1�R!�k�tk�oT���`�Ʃ�T0�Ft*��'�p��$�§F�x)�ϜK�ؘRB J(<	掏�j�*�RlğD��xs
Ԭ��@�J-9���L�A�N���?et��D�R"L���!B�1�����G��|�ff�6ѫ�C��
!nm��n��X���g�G;`QT(��>�I)��	���&:ofX���ϙ0Fz��'��FM��#�k�-m�0ӎ{�Զvטhq4�X*r�}*�.���I��<��JJ\E�q�ʂ3��#�
�� ��r�MZ׬-:5+	-q"џH���/Vn���JQ�g0�w@��o|>��e�F*h(Dx����ҝt��(�� �18"���
��e �'<�v,�d�
�J�,����!��?y��N�V���n�%q�0iƈ�W�剪M�D� 32\�a�њ~�#�Y�8ט�66���ߒA�����ĨV�ƍ�	�?|@�h�ą]����d��x�£��R"4����%r6��#��<	#!J3
HX!�l�,]r�y�ƫНp��5��\�t��nԚM@0�ra�V�X�'�!�	�q<�Dg͈u�ax��*-��Dȳn4V���΅&fI�Iԧh�� ���GXPl]k�m��n[�|���l~E���d�Ie\u��	�Jx��"���}V����T���Y�VݒP�M�8�!��+Nb���'���,��t���;��@�����HH�YJ�2��;LQ��q���6c�f1��:�?�:sf�Lp�g3n�l� 2��[?1qc����'Lk��1��`gf!�&��ڼA��ZH��Ab�B4n�Y�&L�s���[e|�z���$#Ɓ�!a�>)�Gܳe��4W�X�QʟXy�@�(ly�	�P=�����(Ol�@���'�|�C�H�-hWR��W>:��A�� �+-�p)M �z�ף*k �&D��0<1E� 0H\�S��(��)3��C�݀� ��'&��i�����/<�%��._��l`���k�<���P�f푰��9/3n��s�Mp?�3c�����h�*�kD��YZ=�sGDj���Yd"O�ڣ`�w?<Q����!6��|�q"O����ɸX�H��T�M��A�"Oji�bI0�BmZ�	�V���B"OVT���U!P��i�(��$�d��"Od)�H�j�����I2�xt� "O6���dK�k�L���-����U�7"Ov40��9m��eClIt�l�Õ"O�X� �̆}�P��@E�Y�hQ �"O^4��%��XURЂ&F��D 8�"O���B��?pX�H�C#Ӱ;�a��"O� ���-(�Ƹ$3B�RA��"O�A�A�)3YR��C���L�"On�	�mD,Db"eg��*����b"O�`��,�� ��z!nJ�U+t��W"O@a�e�E����[#/E�H[V"O�p fNܒb�q*��O2*X�"O@`���G�vY����;>�`�h�"O*t�r�)u���s�Ĝ|��|S�"O��g �7	ty���LxP�xw"O�Dj�L��2/��7bY���d�D"O��éޮWG��C'��2`�~L�"O�h��J$X�Xeڑ-�(�B|�g"O� 㐊R�\EBtK�)E�4u7"O��$�(n�h�3,��S����1"OrP�B,)CN`@�7�L�)A"O�a�2 �fiJ2N��tȂ�"O���G�d���'��B�n7D�P�)
'DSHA�"�"kj$K�E8D��z�ѵ �*Q�����*4�5D���A��Q��5��ψp�Q�3D�� �ܱ�)сJ����e��T�b"OT�3U��/T�~��1�Ϧ|G��E"O�q�P�.߸I��Y%}��}��"OT�8@-8^|H9�i[q, �3"O���dj�))�0�q"@�gx�q�"O�z�L�&n��M�q�K2��4�v"O�D��%�J�I���S�]	�c@"Ob5����5g���&���5K"Ov�`P� �_M<4��A�T��``"OR���Y=m���BR�; ���@d"O"��,�4i����튮$y���#"O�THG��l�dS���(+Z��"O�zP�]�o��Fm�qF���"OfY2	��1^��,�/+Fj�"O����U�/��,KSZ�"Ol�)L�5(�M�ĀP6g���P"ONX� !f�bH�v�ť"��I@"O����'בU�ީ��m��~Ո]�"Op�1 �#18����C�;�� �"O"�(Q�(;*��1�&v���"O�������:%$��_�٫"O��5HJ�B���r�GբA"O�t�T�$��x��2�2��"O����A;[p�;fR���TÂ"O���ѧ޴b�G��T��"O�GI�]4P�%�ȚP.�"OƱ�! y�Ȉ%��ln�p8�"Oh�1�� t�ra !��)ZWl��c"OZ���n�Q�
���)�;k72p��"O�1��	߅���7#G�K���yr��z��]qK�: ��\���
�y�IGj5U��;'Ԏ�ٗl��yR���!�b���l6,�����y"�,3\|T#�X�G*)@!�S��y(�(jxy1%�x��0:Ʀ��y)��f�ap����<R��z��yb  ��̝#��A6<˖���e��yR$��oZR���agNڊtr�ͅ�IC}rd�B�~DQՊ���٠q�I��y�JUb�	Q�i��l�D��HH�y����\�Ҕ�3OL�8����4���y Ԡamf��OR�4���CT���y�b��e����Ɓ�	D�>�	�'̬T��#��k��|hFɋ�	�'��LY�%�:X���� �J�'$�3�18z�����Ӭ��	��'���e� �X�'O�E���'���{�CM.��yӠ�ݎ��L��'6p���E@�R>���k�<76�lJ
�'ϮZ4BN���5��\45l�As
�'y����<	��c"F��6i0�Y	�'�T-�b�����ҡZcd���'c��HV-#�޸�#dQ$�Z�"O��r��B���1��Q:AL@�"O>E���ɢ>��D"6h��W)`�g"O�,	�%D�J:�f߆1'�M��"O(jQ*��?c�4�F�g�d��"O�S0����xY�ӆ��.�x`��"O`���<��� ( �H� �"O
�Ge��&�\Kæ�u}��""OU����.)���[�A;��y�R"O�$��i�g��"vH��Hq�"O�m���&4�NKM��<�g"O���-sf )�#f�,��A�"O� �ö
��YR�l���Qܜ��"O�Ma��ηr��5Xgǉy�*%)R"O�<˳�\��T�� ��=�n!�g"O��w(ci,ɋ7bQ?�|���"O��)P��P�P�O�3Q�����"OJ 8dfV �b�S@������"O�ay�Aӫs;�y��6:�DH�"OTUP�FF'n�6�sF�Vլɻ"O��5"Н��$0��<�X��"O| �Uƙc� ��+�X���Q"O\�02MV�6)� :�`޶O��}��"O�����хP�4�CCnFW3(Y�"O"ɛ��U.ܮ��G��oB�@C"O�]�e�V�n5&}���%4�@k6"O�|�'�'��`hE��fZ 	*G"O�L+�ӢO�x��Î(!�(�"Oq�f�̊iu~M0�H��;�����"O�mcr�?S!���AǕ;��Q"O���"O�7�&� '���\�P�"OT����؄,�����e��2��%"O�M�"�X�'QJTړoX=H��	�"O����#nFJ��UEGф�;W"O\��A���1�e�<��PY�"O�hB����L>RQ�̞�M���t"OP�a�NثZ��|�G��tv��"O0X	"�W.�tL���N
-tb�"O8:) ���yyS�G�V]���E"O ��T�Q. w��r��$?�A�E"O�U:���� ,U�7#Z|W"O���,]�U���1'mT�"O`M� �_˒��1G;]Ա	f"OԤ`Q �6�l=��=V{�Ę"O"��rJ�	B�����R	fo�}�"O:	i�o��u�LLj��H0m�B���"O���R�u� ��t � �d��"O���#��^�pM�	�M�4Ғ�|B�'�bB�r�H	�6���y4��+�'�|t�5k��~���t
�_�<�A,�rL��R@ѩ,K^ ��N�<a˜S>�)� � #T~�+C�G�<�ϔ��Z�C��8}�ƽ �g}�<�eJ	�VP�gG�4���a�_P�<1DJ�"����<.�|)c�BN�<9sE�{�4D���L�IXШ��AGI�<�!�*I�*�C�[�d�Y�)HM�<�bU$o���2��g}Pui6dt�<a0��/�@��+D�d|z9�G�Z�<���B�[9	�fD�t�MXD���+�(X87���g��ɝ
0�dh�ȓ/7nF��w��m1�J�h���e�'�D��E̩Gc����ۮ^z���'KV����+k�4�6!ΎE��'���`�/�4BT�hJ�-O�%V<�i	�'u�+���42�.Cq�Q6m� ���'X�r
�:D������]:~�
�'�T�F�v\�k��O�O6���'�yz�ě)C�՚�M����� �'���昢We)G��)�Fz�'��M9��V�)k�3��7��}��':nqd�����Xsܨu�j}��'92�7-ͩd~ ���e�p��'��z����ڙ��+ζY�����'D���A��}�va���VN�	�'�����/#$VbB@�E��P���� ��@6m�&�2]�BDԟ2rZ,ڥ"O�i	B��uS�81� ²;U2��"Oh���>Z%�5�o�9
@d�{#"O0�A.G40LP�N��U=� E"Obh:D���T��a��_�:���"Oz��fIL4kr]˔7Bٚ�i"O�Q����!h&��#�O�`��a��"Op= �G�1z�89�IQN2�#�"O���[�-�蹛v	0�R��"OB�2¨�	T��&���Y"�"O.�*b����?�ܘZ��!4��P�Ν	P@)91J�Gb�5�b3<O�7�:��##Uvz�""2��`XBh^ed^B�	~L8��O�?����D�� C��=��S3�&���,��g[x�/�'L�\B�	�3^)(Rk�Hx�%��Ba*O6q���ՓW)l({�c��?�d���"O,80���=q�9�!��V��@p�"O6}j!��\U�q�C�Q�!����"O�	֌ưz�ZQC@�6��u�A"O��(�&
$&�J,j�AT*I�
͉�"O����p���j�^�^� �"O���qH������˂�`*4�G^������/_�1q��6@ExD Y8�C�	�HB@[����89{�,�y�dC�#zB`a�Q��}�+�Qm_�B䉞)�J�A��o���"�C�)"�B��R8�pC�=:IbMpᎍ�&����%�$O_����	6{���
&���cd!��p�6�P��X�X���p�J3X�!򤑟Z�peЦ`�T��T �7L!���Ns�T���%S��j��ؐ/�!��@
���y�
M?Ch�W�AU�!�d�hJ�M��a�����,��!��+F�LaIaL� �%j�!���Z��` �'��U�g��#�!�D�����1�Õ4}��M(���K!�	O�x T��aC�Di�۶-!��
��l�X�B"$d�mT!i-!򤆄�0œ%J�-�ȉ��)]�c!��)I��y$,�?{��mRU	C'i!�S�4��
b�S
�2�G�Q!�$R2�T����R"A�Ap�M�rY!�S�>�$a�/��y� ��R"K!��J=}�t4��D�J�Qx�E5rI!򤖜I����O_E t���$I/!�D�8`�Щ;�!�-�(�'m�Oy!�D�gY���b�C���=0�N�>5W!��^`��J  �m{���$�ŏ�!���8*���:v��nv S���~t!�ą3x�a{�l�l��A�A7i!���L�`�&"U�0=��'���P�!��ſi�E�
�T�8-�r�W?�!�[��j�O٪Zr�1윭*!���*\	ラH
/e�eR�h��5#!�U�J:��r���,hma%�#b!򄛱 DyJ�J^����DڪC!�d�3.N���D����S��B>%!�d}>|4�cq�����g�08!�DI�c�ŰT��+*�%bE��7,!�1Jj�D��nC�R�J��O1#!���f� �ie� �����^>e!��б$*ʡ���D�d�i���!�ݭ�<�aoɠ,G��g��{�!�� P���S�&e�l
�I�2&W�y�"O|���V n}�Qk�h�=)TA!F"O،i�F�;3�����g��w2��"OR������$h�H� $^�)�1�"O�U���P|�%Z�\�D���"O����M�{h��pPa��L=�"O����(#�@I�5A9��Aa�"O�|��iܬ 
J5�@@D"�*8H�"O��`�A o�����@�.F0�S�"O�#U"R;:]ۇ����E ""O=r����l4�PNڶ~R�ѓ"O� ��B�`�h)iDK�O�D�#"Oj8��F�,2�U�Eg�o�U��"O�U����(~����fR$m�(5b"Or!3��l��!���?vNP�"O°"&�נS�l�H�
�)8VU�V"O��#��t@���WK�W<�R�"O����Lf�=���U�4��s"O���g�&^[2�9F��a�}��"O�1 ��X�k�`KB���4�N8s�"O&Ixg�8�0p�Q/�.>r�[D"O��I���vp��2NA�3ؐQ�"O 	C���2�`I���@g��a�B"O�M:'E�i���ؕ�� ��"O�0!� mΌ($ �о�`�"O�k�"�9j�j�u	� K�P���"O���=eQ���&���h���"Od�C����ys�͗`�N��f"O����*�BO��9�3"O��K%�p\��K��\���"O�M�&愊? < QK[�#��i�"O�HR��pfv��J�<9s$Ha�"O0�3�ʐ��4̠�(D$]��"O8���o�:+u���#��BP�C�"O<�ɧ�
0��䐲e�� ��p�"OhT�c*:!о��#^% �쓃"O�@��\1)I�ȪvbZj�y�F"O�I GdN#MJ�8+g��}R���"O4u��ce���#G��|ȷ"OT��	B7x�����n�6̨݅4�!�d֩*_����/L�80� �.�!�d��"�.�)�!�"-�┲�1!򄅶T��%�C�ƄҚ���(&!�$�>5j�D��K�F�8�q��C��!��~���z�غ3��1'��"L!�$��]���7I[6W��p���RD!�X�"lz�qD���������8!�$ҋQخ�˴cB�B48�P��YZ!��߆O�&��c�M2}�5yկE;Z�!�dF�F�`�w�ҤrdD�1�E8tJ!�D��I؄�����;ZX�Pv���qG!�Ę�z��rE��;W�1��I��|-!��F�����ΗM:�0���S�!� �GؖmYcN� |=��� ƀ�!��d�&�i@���Q&�4{�瓕d�!�$ۄ^���Da!�.�n���"Op�ʖ�ݭ~��+f�A-P��<�w"O����N-�9J�d�g�93w"O��"�菙 �(P��"�ݘ"O�� 4�H���P��C�eex��"O�%bAO��	 � �n42\�E"O���'k�� q�^�>��`�"O�mc����� ��ȸ'w��"Op@�Ũ�/jր�1'�A ��Ě@"O� [W�*>u�"Ύ���*"O9�5��N|P}�u*E�
h����"OR���]�ol%�7�L.UCv"O�JuG�@����CHJ�#���"O98�!�$�^� H��g�}sG"O*tZ�m�&��[GɃ����a"O�)!�hR1?��8FC΀Aր�j�"O���Ŝ.'ZI�-W�J�J��"O
���A
�H�v �Ԇ��g&5�#"O�\��^�)׊�q�z��4Z"O���@Z�➠��CŤ0�6u��"O�` �@�%%;^�[��M�>D��sv"O�aP��)#;�i�a��(%0h#Q"O��Q@G�s��24eC;`7<-Jw"O�{�iV�/����X�W2�`�"O�X�E�ՍC��)���U"a'"Oص�@�E�B�v�A�ϛ�Q���"O��(��Q�t�3�G&.\�"O~jq;3,I��LR�'2��e"O.谳Oɢ*�T2��Sj��r�"O�u��"	uR��ʢ1���XA"O�`S�ͤ��Z��˨,�L�d"O�1���u�@�%M�+.3�r"Oơ�U(�77xc,Q�x�'"O��(���j�QL�X���"O�d(�`��^B.��a�3`ȴ�d"Oph�#ș	�58��7���V"O"���@�p*䰒���ڔ�%"O�Ԙ1��	o�
䩟�K�@<�3"O4�� R&f���B��L�ֱC�"O��@��@:�&���!�`�ib"O��9Q�̲f�x{�)D^�X9��"O ���B�1=8m��a�j߆�#7"O���$ۥ@#�;�Đk78��"O��!��b�16/϶k)`)xC"O �C���@� ����n1#"O���p	81:�[@�d��9��"ORM	A.@���P�V�1�n �"O(A��5 *���Ĉ)B�J���"O��x��
�v���8W���H�ZA"O��C�i�h�M�H0$"�"O:u�@��%�4qD.;��C�"Ov$b2,	���$2�*.�Ba�e"O��c"תyr�8���'�V��&"O��1� }z��&%]�"O�Ha�_��D�:bo��MK���&"OҼ24�\�O��\�!���m���"A"O��R%(Tw�e�S��w���"O�@��@�9^��T�����ő�"O�k��Ś>c��&]�k���J�"O��e�e��	�+W�C�2�SS"O���TO�xcZI��)B�����"O�5��'�/n��J�9>��=W"O���f�Fp#�T9����l}p���"O��å
R�s�¥�B]�2��$"OV]���@4�(��g��L��ْ�"Ol�C�(:Z:黳o>|����"O:-��
�n��}Г�
C��%9�"O�x�%N�
x��̚� Q).z��p"O�Ir
�dt20*w��6}Ѡ!"O�����3�h�з��1Z��"O@I ��vAfLs�T!�y�"O��[�茱��B��9[�ԡ�"OԀ ���l��(��_Ixxh�"O� �,'�^�=��MC'�:h�a"O���B�=!%T�P%�3s͔	"O4r�$qk����D�8�,8P�"O< ��8��X�'a��m��\z2"O�H�d��[�<I �@W�n�\�i "O$	�6&�"�\���o�h��Q"O��PR! "|�ɻ�-���"O��2
G�R�LT;�+Ȩl��E��"O��h��K�N�n��K�m�.a�"O���TK,]
�ʊN�>m��"O.� �"B2�e";� M{g"O�2%�+�e��Z�b��Q"O�ܺ%��0�ތ)%DҊnCLR�"Op����&ȼ��ă5l�4���	i�O\*�K��6��d�Q��0��MH�')��j�c�3��as�	��PL�9��'��p���� �֙��V* �����j�+R)�r��m�$-��JzY�ȓ5�Y��l�8&� V��n섇�d�\S�H�z_Ν��j�qu�u��c�4��! ��NT��Wf�"ar0'�����;E���qeOD/$L�4`W�
9D�vC�	e�Џ��\x ׶y0N���r����Xݜ(��0@���}7F��$ePd�'���Sj�l(�
r˸H�`�J8o�FC�I37z�1��^I���AΣ]�8C�I>P�Nк"���}�vc�o�C�I�jA�E�bN�f��D#U�˓�?Y	�����3��P�����.9�(Y�ȓl���3�.�@���mK�8N���,O���ĄV�Vp��n� zM6�E{�O"Qѯ�:]���qOё>�|��
�'�%����$/)�x�����	�)�	�'e�a�@GX0+�H��o��Yp$�
�'_�p�� �YPzDB� ʤz�=�
�'�;FL\�Z��p(�>y�
m)
�'��p�!����h4Hp
F`�&Ű	�'��Rsτ��T�8�)Z��и�'���ۤ�٭G����"-X,a�,��'m6�;�o�$gV�{�j�.t,����'�VuH7��e���b@��m��)�'����疗{0��ɾaj�x�
�'O�x��N^��4Z�(-�X�	�'��<���Ⱥ1͞X�i�B�9�'Uh`�&Yp�E��������'e�A���O@@����?ql�)�'�V�h7yST�g� �^a��'��̚�"2�U�f�E�'�����'�	���2��)���4-��Q�'����>S楩��S*4��'���xa�ƝR�ș	�ރ(T��a�'����� �XȐd�������'�ʤ2e퐣z�t��g�##N0 ��"O�U��D^n)�S��PM�\r�"O�8Â��;p��E�Fjk�"O�����^>�ZX	�E�h8����'%��'֕i�h�*�����G��ʌ��)����/LH���/L.e����)���y��R�0� �eΝ-L�H�F��'�y�L�ph�R�M&#�0Iم�M �y���'c�����6Ns�-��BJ�y"��u�pZ�F��C��0�B��y�+"���C0c�>Co��9$H���?���hOQ>I"�o�qنo�[��h�7�!��0|� V=��>F�0�����&R�L���D.�S��0X}��݄)��r����!��7�h͚���1�$��1�!�;�-��)�}����f����!�dق$b�*�˚?�����T$+�!�Ik��%��"Yv���X >��|��(���Ag%�,��[���/j��-�$��R�O4�`�N�&k�� �L��PZ�jN>������f`NȢ7@O0X���i��!�d��k
jyA�a�<!�Ԑ����7Y�!�؎D���u��j�z ꓈UW!�ě�G��e��I��-+��(�[/A�!�D�('�j�r�@S�5b}�!�ټb����5�g?�uz�K��=����G�^���hO�o�\]�cεf�F�B�+շ����/v����/Մz1ah��ԍ��e��h��3�U��Y98#�L��4 ���m+�!C"��:�x���^n(����(A����"LAa'ִ���P~򋙴c���C����
�� ������&��O���ac�&5�6(:�+�!~��R�|B�)�S��l*�FаȈ!��7}��B�I��٘�� +TɚX�""K,��C�	 $�n���rR�xI5e�)U3�H�
�'���񔄂�4��p��FQ��(x
�'�0Ч�^�6,�XP�o������'Z�����޷"��$36j��"�
�B�'��9PE�
Ō,ƍ�'"b ��'�dEI7��U����	�W��x�'W ړf��,�Ҡ"U�3:��Tx
�'�h*C ��/������0�LU
�'�-�Teϲ)�}s�`�8?�LA	�'����,�0.��Q���[� ��L;���+�p�h� �+�8 5���HE�6"O��ҧ�<S"@
A�;aH:���"O��p�� ��yd��C���`"O5�6��yh4��!�.b]+"O�|���M1c�	A �=K4U{�"Oz��׀ʛT�<��E10���"O>Ei,�/M4Naaf_)0"��j��'M�	Vy��Ӿxs�
��H��Q�0ˍ6�!�$ך�.!d���]�:L���� q!򄊯�$�*4N޳y��͢'茭$�'�ў�>�b�$H�3(��zh6D�����U�M$LP�N��d�@G4D���.Z��\ɉ���D�(#-'D�<S�.^?
�hq4� 4� i#|O�b�Xc�N+I^@�Q��M~��ɐ�3D���T@U�ʵA�ܻ#"����0D���U*��kp��0"�O��H+.D�T��)�+ÀM1DaM�ZD�Ф8D��A2'D~��*C��]W*��$`:D��j�Oӆ�<aඏ	*sb<�0,%D�@'��I��|��c՛Ng
@�#D������ ��;Db�"V����"&D��RU�\ւ���T�e<�R(.D�p� F0%6nU{��љK>��b��O�=E�cB?�4�''��6��([F�!�;%`,�!���'
j��Ǘ�r�!�$}HH��������t��a!�d.&����8�����Ы�!��Y�C<ؑ&�p��T��&G�i@�O:���#uG�=X@��<q�x�����3
��՚��� !��Aqx��Q���d+�S�π �ItlI�.�0h9��80*��Y"O����I�h*�A�"��%r)���7"O�M���1)xּ�f /z�0P"�"O�Ed��U�b���
+w��e�"O���fDn���3��M�B�{$"O@}��,�9	��Q0�G ^��|s�ONA��nT�	_fJ0$���	�0m4D�0��He`08�D�X�I(�)	6c2D���!�K��<J1jU5�P��/D�`pի��Q�(�aԸn�Ȣ�-D�̘�(X$U�Q3�%/&���I*D��ђ��;'�VU�E�8#4�ۃM"D�`��k���p %�k<���'i!�O��䃁D��*�p0�j�◵HB��5pr�M;eN
�G2�|��C� '2B�	7f�����b��*�>^S�C�ɦP��ӨܶsV�iU�O�w��C䉾4R�X��Ү ��iT�6Y�B�ɥa*K�[b�U�#DЬB^JeyV"O�42��� ��0Zcʄ#����"O��H"L\�"	��B�$��q�"O��9�
��m���QD���; d�!�"O�$�7��S���b�ذ��"Oݛ�!�b/��2v!��x�Z"O��S�*ܙ?R4��^����P"O�a��CT7��EM$�8i�V"O�4 �śq�F��W.�$V��h"O����^8`&�A���)－�W"O@�+�˄���٣�ʍ�8��'��9P���8(�f}�I2Xj����'�)3�_�Wؐ9�S�@cRq�')v�B0���IQ����!�(UʴJ�'�!ڱ��>jܐ��Y�!74�0
�'�n�f�B<x[��1�X�
�'�"�+�ȅ*A�� ��Ĵ@�X`�' N��@nS�Z���A$ŬJ�5!�'P(�1�C�a��d8�$P�P�T���'֪�� 1e�ՀU��-Ml�`�
�'�Qq̀eI��ۑ׻O�n�
�'s5Hՠ��@�M�PG��|:H�X�'��!���܀M<
	Y@K8t�����'����B�ec,�!�@�Yf�4��'����n��u�d�h��$#���'̮�u/Z�]��݉�fډ+n��{�'z1``��]Y�y���-�����'␽A�^-D�$�рI�L�襁�'?&X��GM�\KTt�ԁ�{����
�'��� A
4���#�V�l� `
�'��y*d�ƽ��S�n�yts	�'@���N����h�%��o�L���'�0Yx� �gs��qp
��7����'�H���dO$�.�2Aǈ�2D�J�'pv�S�F� 1����>���'���1��n�^z�O��7�T��'��y��\�VH*�1`.½x����'t�	�nS�G��U�$�r����'�&��G/8�mb�.R^Z`[�'�jgi� Q6*0#�
A��UB�'<$����նe��� D1)Ɯ �'������I� �"M�4-d��'jV�a�!�H��p����1*(�
�'����`���|}�s��2\8@j
�'H��5-F:%E���3Ōz�L��	�'Wn���j�x�5����zY�Q���� ��7�C�_�� ��,+�TMk"O,)j�.�$0jZm�VnBm�� �t"O�u�c��17`BA��i�eP6�'�1Ocd��	*�(�,D6O���"On��5��u�n�S�E��U[�"O~���-\;\���6%��ym�E§�|��)� ����uj '�<!s��o[|B��'0f�H�'�M�g�:9�AgβXZ8B�	S�j́ �ƞn���B���**B�	?9�(̘Cꇨ+��� 2��4b��C�`�l�A��� G=��]�Q4�C�I'�n� ��.N���yg�[�D�XB�%E��Х��I���J� Z�V,T�O��=�}�1'�ltH�1�=OJ��D�C�<1�᝙%V�ţ�ȁ�q�*e���G�<I��K�]Y��s0bƅ)�01��O�n�<9��G(EW&�����A~�qK��_�<)�Ꙟ\7 ��gET�N�(�«�t�<1� �{�|��!�#o)Pd�%%s�<Q�BH�%
�3�,�h����fyb�)ʧ+����eK٠zH�hY�Jˠ+ap|�ȓB�(����� ���~� m�ȓG�p��F�:> [�n�2U��(�ȓ����&`ťlm�@: e@�6�M�ȓ���1�I� {�ZK&������(�rΟ9w�^���hQ��܆�\�~ԠUJQ�^Gz�Վ�.'"P��{���{�b��iC4��'���@U��Y(�ԃ�Ӽz��,�S�ǊA���ȓ=�$)�ȿ��T㴀O��h܄ȓD��蔋�JV��2�@O���x��e+X���n��k��)"�%HD��g������%e�|@hƂU�#z����}<���N8�A�
� ���	��t�<)!���Zl��jS��j=2�o	j�<Y����&�ع8���/��H�b�f�<����~��d{V���?�~��0��}�<)�V22�5��o 62�x��M�R�<)ǓY���,�_"���K�<iͅ�X���L����e�fFğE{����2|������D6e�X�0��BB�	!h����I%n��
��ͅ%8B�	."<���H��Jl�a���k|�C�ɾ|r����%�� �T��&D��K\�C�	�T
�00��g�PL�� �w�B�	�:�l�
�.ķ�K���;�����,�x�R����ԞL�t[׍�'t+���y����X�x�� �3�H�@0����t��*(D��	�&^�> 8���
&�|8V<D��IM�E`Phڃ��ɥ�9D����IV�D���$�׀�v��& *D���S�֠
B)y&EX9%�&$��'D��
W�ˢ'ɚ5�W�U5U`�6'#D���\
�Jݡ�H�,e1�䰧�=D���� ��<��	Q�4��I�GG(D�8�w�[�$"HT�bA�-�V�Ȥ�%D�$��O��� K��W3l����6D����*��2sq��Рmi23�&D��F��-��<���� ��-87�$D�PH��¹�F����FX����#$D�\X��V�>�ɰ�3�M���-D�8�l�)7Ā�XG�
�;v��BD'(D�Xa���
�T�Ul�q�`�I�&D�x���fJ:��e�C�0,x�:Pf#D�� ��u��+t5� ���%���8�"O�U�C�U 4�|�A4��:yDT�w"OD��̌�SU�{᧞)/c��b��'(1OJdA3E��z>j�# �!pJ̤JP�|��'\�����@���
���"���'��M��h�(p���&�+�����'�<l� *C5e� ��.�2T�����'��x�A�NȾ�ʄd��di�
�'ޕb��=Lc����� $wR�	
�'880��W�� �9?/H�$"O��B��G<H�����BŕBUXT�p��!��џ��'�R��qE���}��Ȝ.r����'=��[�/[+R��y���xJZ)X�'`�1� �V�$	����l�R9�'#�Rb��2��Aу�F��'7�}�G�L1����#bCN�fY�'�� 25)�(5o�]rS�F�wX���';ĵ�'�C~(���I��n��)�(O��OV�?��'{�8�v�X$�ޅp��� 1�ֈK	��O�}���P:�`8�ZZX��`"O���sǗ:kr�])bb�0dy��"O
�@��Վ=��졡O��]G�|��"O��А. �7،�醏�\,L��"O���#�H�8'�Z5���wL�@E"O4Qؗ�J�j�
����n�H4���'�ў"|r�'���S�g�W��1����>IF����O�}�E`�
%;�$��	Z�l}�(*c"O(���_BŌ
�iЉr P�"O\8�dR�F��Xq`	�(9.<q"O�������5��-%KC|�"O� ;3E
�5�@��ˣh�����|��)�S�'��D8 �X�}�	� �P ���I'�T5 I�%�����eG-�\���	^̓n8��!���W"�!7��=m��l�ȓH�	�3�Z9�9�C��\��݅ȓ	�6	sh��*�LP*�V�0��d��q���S�|Bd:���9:��ȓ=:���G�ɍD�>$�t�J�0R�F���8�j�&a�e.�����Q�g��㟈�Ig�'���_3 �R��P)D�|X�B��&f������I`���'�p����w�lT�S�-<�D��'b9Q�� �g�j���K.t�	�'�tap�=$x�򭈒q@*��'�B����N�H��!�M	�@0�Z
�'�x�Q�L (����F���x����
�'l"�TgI�f]���eo�8^���C�b�'�:��@�O�譱�IφWqdp)O�O��}�A�����L�4����'[)�"Յȓ	�X����~�\�x��-`�"�� �q׆����(p7$'Tf�ȓ(�6��e����ĳ"���ۓ@ D�t"Ĥ�������D�R��d�� D��:\�12���Y>��g�?L\!�dȓ`�2E*d�c%�|��	ay"�'��O��?��{�
Y���7�:$X(��(\~9�B�i�� 7!�<U/Pa��3����B�N�N:�����N�H\�e�ȓi�N�#�
@�s�N>~Q0��ȓt"��Q���)������O��2���`N�c�#�T�{�@�9�v���y����IH�)>��#�JlJ�'���>\JB�S��|�`�BuI�/H�C�Ʌ$�)����T��Jv��{��y��v�z�"T�g4�"��V�Y]�y��S�? "�#��9j��(�a���]:06�'����D*��;�Z�Q�L�!oDp�e2D��a3��!S$�p7S(.|؉��0D��s��4�D��b�7/�F8�-D��p�j��D��BCJ�)�
@#��'��hO�	�a6����Dgs��J���4r��5�|��I�v���h�81hܼHj1D�t�t�ן�и��a 2f�Yw�/D�,03���c~�yZ2"K�z��P(��)��0<%��9ykN��ҍ-���@{�<��@P'�`�TKO�Bm�!��Py��'�O�#<�D[.A
��'��J=pLx��R�<Y�8X�p)W�ïm��#M�<�$�݈@���M��m���� Cn�<i%F��\���+_+>9[f�V^���hO�Wf�dP�J+l0 �Q�A�6۰M�ȓd(q�0�٥$�-�u�B�P��!�ȓ b@Q�#8ߖp2�
�HJf���ٟ��?E�D`�9y}`hs��j%��1R&K�|�Ig��x#Q�*-��˦�p��h��7D�,�fK�Z5��!��	ʆ��І9D��K�
�	�ԋ�����y��4D�(�2�B�?/�����NF׆0i�'3D��9Gh�����KZE,�Y7I6D�����.�x$����W�2k.D��8@�9xY���T)�`��Mh���O���S��}� ӊ\\*�K�:mr�B�T�<!�։;Tlp��7��R�R�<��D�A�V�����;G<e�a%Vf�<)Oۉ,�T1��1F�\"�_�<�� ?����"[*a�����q�<!��P�q�|uP$C�(Y�`�w��x�?!���Oݑ��kNC�ӒP=r��t"Oh���Z$%��@#�P�bV!F$!�Y�4�Ƚ�pܔ$��r�C�Q!�D�2@r@����N%쮥2��G!��"�4���Z�
M��L�pb!�W�=g<8���S�#��1KY;LN!�TsWk	�<<���۞/K�}r�'��� J.ҹ��G����a����&��)�'��H  @�i�� ��iS/l���p�'�VՁS��!LW|��7�EZl4��
�'���*!S�ց�D�?��%��'X>�kw��4G�b8:��̤DAf���'����@$�l%���$G4�ѻ�'麔���"
�Ͳ3�A}Zl�I�'����@a	��C��',0������d-�O����!o��)&
�\i�"Od=�UnL�E~��r��FU���"O���׃	 �M�ӆB�m����"O*�3f�Y+�zИ�ԗ2�pA	u"OD;ec:��u�
A�CXd�A"O(��%oѭ���Q "U^j�!�$˥,�*hi�'n�9��ҪOD!�D0܀A���S���Bf✝g4!�$��p���`b�@�y��`p�aA�|!�$I��h<#�$��8��D#A?4�!�D۽u/�U��H��]:�L&�2u�!�dʍ-Lqe�U�pw��2uϐ���'+a|b&�%��1� G����cf���y��P����큠.� ���O5�y"��4�h��b�����0.�yr��a�$�J .�{� ������y�Y4����G۷?��U`r�ȴ�y
� Rs`�:��ڀ��?{�T� t"O�Y ��-�(�QǧV�T�fW�X%���ቮj� t���@��M27�XDrB�	0*2��#CFB�pf�-CgD;lt�C�-���Ċe�z�r��C�I�%��c��\Q:f�k��B�,ל���b�#g]ty�T�U�"��B��%7Pd)��Y -�l�6BB�B�4 _���7fM�9V���T�m4~��!��=���y�l	m���J�
,�Ĺ֧��y�M�&p|0��!�N��`�6bT��y���o�F�铠I�%�X��sB���yb#H�%a0��!�Z����s�i��y��N-*�#LWZ�3F�.&�vE��'�.�C���.^�m�Sa�% ����'�e��H��e!Ҽx�M\�S0����?y�'�ҍ0��!
jd��Ɵ�I%����'⌅�v�X�I��,�u�RA�<*�'�.�Z	T�K]'<�d��z�<i���}ݮ@�*�0)d����Ys�<��$E)3���ITÚ+�\lF�c�<I��h?d��7	�q���&O`��C���Iw�J���Cc��zi
cc0�t�)�O��	8B���G�I�~�PS�й}��B�I t�b�`O�t�`��d���tB��;'�!)��M�U{B	G)֘C�	�-
� ���#���yB!�1��B䉢 ��uAQ�ĳG�hC4L��}��C�;m*<����0d�$������C�	�EI0D��Q�M>�C���:�C�I�M�x�=�$����p��B�Ƀx�������$ש�:p��C�Ʉ0����ѪM�`�� �&��r��C�	�v�Zȡ$a��1���7!�3Q�pB�I��=���&of11��� LҤB䉨%U��� �k��r��fZ�B䉣p�t���o�8yt)yu��O�\C�I�9p��Т���Acg��C�	�`Q�!���\.Uc�D�Z��B��.78P{a$p�ܪw�ФO�C�I�_���YB�' ��kƀ�TR�B�	UO���0�CY�.ț���H.�C�	4f�
����͂N*t�����_BC�I3~��Hcu
Cd6�9���64 @C䉑|Eȣ�˻X{�� �Λ@|B�		��@�"߲k��P�
L�vH�B�	p�����N(G��\��B�	�` .��DM��T�c��7hVB�ɛN�Y��U�(gJ�)C� �B�Ʉv��\1F�?g�tk��m��C�	�ej1�#��1;�Q�5�^�[q�C�+�>�s���
�Ԍ�$�'YcfC�I��X8�uA��܄�q�C (8C�� � ��$QT�m��D�z��B�I�ʀГP��JM�� 6iO;|2B䉡v����'�X�J�Q�̓�B�ɦ���ҡo�0(�iU
��B�	@�p��d�D	 �Q�4�bl�B���:��"�_�,l�q���8^��B��%��t��A�9y1�-*5m��i�^B�I�f����!���'��4B�I�M���SbP�B0��SVl� B^C䉺Av���XH�^H�C���B�	:S�Z�ŮA�,�7��=�|B�)� �L�7!��z��{�#/j���"ODX�o�7N@�H�#NE}���O��r �J]4��� R��BЁ�];!�\�&���S"�H/tZ��q� ��z1!��$1����
U<@X�jj�55.!�^#t d"3�)��o�~!�d��Q��ň�Ε��^!� k]�?�!�$���:�����L��8���y�!򤉛�4��!ٱ0��R���qsa~�-
�?aU�ݏu��0�$�f~����=�y"�L�r�C��!8I��s�K��yB�T�S����G��/�R\&�y�D� J��Y�6�G�)�x�i��F&�y�/A%P���#�B��h[s��'�y2Iͳ&��\(��־-��/
&�y���*�ڭ�X<��x�@h̐�0<y"�
ҟP$�|��#��w�E����=[�t P##V�<��^�|E����N 	�8i˷��N�<�nR6:�j�؆�	�9��(��C�<u+�?�|8��a�1D�p@H�}�<��HTkZ���E����\}�<	��n޽)�n)b����Vz�<��Y1^z�0P!�[&9��[1��x�<��K(f��x!��8+�ec���_�<y��V!��� ��	���rRl�]�<�V�U|~� /@�:,�j�A�A�<����'��y���e�1:�a�z�<A�G�2c������4BC0h@!�AR�<i�
����Ө�B�<���Di�<YÍD�
in-�	J�<Q��ƪf�<tbC&�d5�U G����M�}�<�P��O_b�C↜�Q���Q[S�<�� �"78d(�ڙP��H"`��R�<�A��2�\�'�À"2�ŀG�Q�<0����u�2����
�����N�<���/MAVQ@���@e��a/I�<�D6hd�I��{�2U�o�N�<yag��(Kz ��nY+䙴��A�<u�Ӡk,~��� 0k89C��z�<1.�d3�	:D
P�il�����p�<Tf ]�Q�rk�X��x�<Q�%C�*����3*�/���) Mu�<�@��T�s��W�tp�2�Yh�<q�B ��x�s�fЯ:ʎ,��o�o�<�2�]-@��u���@�H�~��k�e�<!D���ʅĂ/�� ;q�R�aD p�ȓ�X�)2�x�B���G���D��?��	j�ǔ���R���qN �ȓ� �:����\H� ��>��ȓ,�����&k���%�̭[P��� ��l�Va�qA�<;�	ȟD8,�ȓgb�h�$)�<[�S�F�T!��n0���`!	�e��5;���
Rj�Y��"dHԻB�!��`ju'L�++���6"~�9u�n�ʢ��y����D�9�wL�mxV��"�z�%��_��Y��%~����C�[ %�80��{��y�gR�,.���Ȓ4F�b���kЕ�⌘x,����(����y� ��5ij\i����-:�=�ȓ|���[t��̼\��������,>�8suC´x��4�C�R4Hrp���:ġ'GCWl�bbh�$	�8��T�4��"E�1�`N+r�����S�? *���O��Tm �&�0���
�"Of�[� %A�T�X���W~�]�"O^xPw���U��e!ƃM;;�d��"O�s�(�pXuB�oў9܄=�"O���I	D|i�u�d� X��"O����/ujȣm��T���04"O�x�%^-N(�4S��<� �p"O�,JP.Y�1��h���\$j�(&"O�0��薍i��IS)�&M�Ըg"O0���BEHk���A�k�<e"O|� ���.U�ؒ&)E(HD}x!"O2QX�5]��|P ]�3�V]��"O.A�	�
|;!fK
Œ��g"OV����Hk��wE�/Q��"O���k˃Bɨ��q�Xcp��"O:H�dI��艺N[#<R���"O,�@Ѯ�L/��MTJB^	�"O��8�IE V>�K��U�Z@���1"O���qJnB"e�P+P,H��"O�!�y���)�� �}��$Xp�!D�x"3���7I�]J�چB��D�%2D�D�&@	;h�p��ʙ ����E0D�������a��G6xC��S@�-D� �.
p8"0E�@ߌ��m*D��FB�50��|A�	sؒq9�`=D�·�ų[�`�gkQ�?�^a�B >D��Qb
�9#g
ѧ�.�-B�=D��5 �!͖�p�*K�E .� �:D��A�G�<� �v�ތJ�d4`��:D�B�h�(��u)�7Njd�Re�9D��gC�� �|�XFK���R��sB,D��)d-�	(��3O�;5E��T/5D�P"��ɺ�	�A�-V�ģs�.D�[���N��L#jۦ �
P��7D�kq	\>(�B'JY50����K2D�|{��ν�&��/�]�I¥�.D�<��"�D�R|s��,EB�Ƈ*D� �p\�*�z�GW6PI
���%D� �@�T.y�E�'��7պ��#D��S����O��C@����N�q�H"D�l��F��>��E��42RD+�?D��y��%f	B���؄3,8�!<D��5�e 혔�S�*_�P��/D�|���K0.2X�Q�o��@�V�*D�$Y�n�2��� �<TRG)#D��A�HV$�Z��v
hx���!J!D����,��]9�-�����!,D�`�@mJ;d�b䉗��	D��E���)D��:��\���x#�9���i�%D��k�Ã8L��W�&]����@O"D��!DF����2FO������;D��"G�J<���q4�))O��c7D�`����� Kɂ�K���(�E�5D���P��i��� ���-a��`kw'2D�<2�#��b$�R�-�v��	,D� *��7�����i�V��g�(D��xDd�6�f�
1Iݲu�T�P��$D�L�d��N�q{���a�~-9Aa!D��RхA7A�Mq�Æ9�h�B�=D���!�Ĝ`�b��Ʉ�8�R�=D�a4����25 ԱN�\��l%D�f�\�b� ��TW'b!��>D�˳b�'g9��W�Q�rx�bN?D���N�3��<��@�F�4�'(>D�� *�K�>*(��k���E�6�&"O��c3�҆aKR�{�\	(��`"O�dq�oʴ\�
���1uu���!"Oޜ�0���
x>�;��tb�m��"O���qgA� K��o�\4��"O�=��-�lJܢf��&Z�)H�"O,}Ƈ �X �ɐ�02�"O�]��dS�A���*E��-y��ԋ�"OZ�B�A�9 |2��e�VK�
�PV"O��{�&�)tw��$C� �@��`"O��P����Px0D˥�!����g"OL��W�H�!�@(�AL�s�tq�"O�!��K�`L�@ݹ_�h� "O�L���~m��x�l�dcN��P"O��щ�o���@�	�M��H��"O��B���.BŚ���J��
h�a"O؄�$��2*�.i(�	Lj\��ц"O~�{cȃ3z�,"w��'G�`#�"OT
�O��e��3��y/��bR"Ot؈�Q��E: �[�Q1pQ+�"On���/�
8KX�@�4@ؽɤ"O��@T�*D��(d�\�B0�`(�"O~�D8]�l��ԩ�R	�u�"O��ZqnT4t�Fi�ǩ�j��d
%"O��p�%I��^̚'��#v�8 T"O&� ��vw�0�� T� �`�"OyP0��T``@ɯ,�v 0�"O�qS�"�^�4��s.D�m��P"Oy���k�<���L)�0��f"Ob�"���C�z���MV�k�Ɖ1�"O	*�]~u`ɣ%M�;ͦ���"O�\2�)d�P��[��Bu!�"O0�S���#Y����j��Vb쳶"O�	07�^�R0Hp�7��. (Vr�"On �VnH.���;�OT�3#�-9�"O.h �A &�mїn�|��""ON���a�:i<;f�RP B�"O��SV�$2��D�Ŧ�#����"O�8�K�DP��Qr��d�5"O�9�"�Y l6��@��R|�kR"O����T�Q���3bO1"=K6"O��k�IJ'�x��':�(��"O��AҤRǤ��`�.I�2��"O��ҕ�Q,�:�,���"Ol�
@ᐼ�Wh�v�B�"O���W�GY���鋥p|Ը�"Old��� �@�b�Y���#R؈���"O@}9��P�B,�K&���X�9��"O��y ��6�(m�@���|�ࡳ�"OB��A�(,��d��[��Šb"O��h@(*vbpuY��:pv��9g"O��yя߷Qv��J�5D�X1"O�=xuo�
i� ��-qjq�"OT	��cx0��=9�Ġ�7"OtU��IQg6@낁��m}�Ӆ"O2i"4)݋��J͸����.D���sᑳO��,kQ�Ƒn�b`��)+D�|��f�d��r ���`p|	�qi&D�X2���q0��*e��.x��i(D�L0�k�&ZeA'%}�$�2D��Ig�$s{
���\ ch�	x�0D��1r���=%.h��V���+F�/D�X��+7v�TcB�ҝ)䍳��,D�k��� u$)��ϔv�A���-D�� �ѡ�і�x��2G�)`�tDy�"O\첵��N�x8������r�"O�I��bAZ8�P��'(t1��"O.y�%,��7���
���,��i!u"O�2�G�6t�ɪ-���k�"Oҽ�Bۈ7��M5C=Q��q�Q"O�҃/N!Ocv���X
/��s"O�5!5C�M�<X�a(�v�ے"O0-j��M���*�C�Rpa��"O���a�)�j Jϗ�Q
�r"OV-b%�V�E�$m�1�X��"O�5B���H���a�l��y����"O�``��ϬtTlJL�7� ��"O>h��E��7�A�:����2"Oƴ����-*��RB!}�%)�"OT�PErě��R#z@lh�"O�e��
5�>���eM�:O��x#"O�D�%���5��5� A���b�"O�r`*�����:u��p��"O`Q6lF�Y�f�I%�I�/�I("O�t
a�#;�6�<��r�a���yraN-���Tf]��lJ����y"�ٳ9�"��#/����R� ���y���G��Ƥ @dm*�����yRJ�3�,�x�"Xy�}	��yB+��u\$ȶ�����5�й�y����^=�LP�-E�����B���yr�7#�b|3PNV�N� �*���y"�i��hJ��9P��"'��y���0��HC�-٠K�Lܚ��H��y(��;xBuRp�>p������H��y��4�����J��*�y��
�ydQ�&����KD=�.��h���y"
B�"�Y�1	U�1m"�)�j��y5��7K���ٺ�%��y2&ɔ~��-�U�N W�ē�eL��ybm�������q�4�H��yb��9��)9��
��J$����yB�̻G?>FE�Ld�b��ɢ�y"�ˍx��ˢ��E����jN#�yB�O�݄X�/8U���4`��y��\�Z�	�fN�?���ȧ-��y�+�X�NШs�R(2x(DS0!��yB(6�,uxī��,l�B�e��y"�ǭjZ�|��a�8Q��������y�a!PL��	�I<�9c&L&�y"��[���q�[!,��JW.)�y��/����㌈;R��I4a��y$�5c���Y7bٹF�A�'��yrh�5�f�����;!h�*�g�y"�ǘM�J8��œ4/�)4`��yr��&I���ibDɷ&�4��Ƚ�yb ބ{1re�̎$�.�B�-��y4�L]¥O�(FP+ �3�y�aQ�Hl�\#�k�5��r�!��yrmW"#'pEb�H׸31L��#�y�-�30�4�jf%P�u/�=H��)�y�mܝ~�Z���
l��h��W��0?�-O�I�v"W�	�`)"���[�H<ST�`��������D,6&.�`2��~lB��`�pyWfER��D��i�
�Jb�\��ɣhY�aB�	�X��8;D�Ph">Y��i�>?栁�#��IJ�����T)!��H,��� ��L�����KO<��7�S�π � ��f��2� �*%�lZpO��v�V�G�
h�bZ�:j�}Z�GnyB�)�',���a�c��=�!�2��|Ɇ�II~B»$���3�F�n�|b���yR(�~�Ĵ��InU�P��+���y��=<��EAǡ�+m�؀ C?�y�^�z�$����a)��1�	�,�?ً��S�Y�ژ@�m�\%$Wp�����f/)ck�$RX�@���C�504`&�O�㞼D~���%-4ЅA�lɒ?�0�W��D��䓎��|%a��I� |z��[B<��*OJ�.T��!A��V=����j����D �S�Of���7�9~�8))�h�$����'U8ٲD��(Uށ�f�:~}X�������9�)�'K�*8���[qD�lV7H86��'+�x�U�S�=�f�z%��2B<Tq/O(��䉵b��@��%�$Y�*l#B�C�1O��=�O�rj]�Ns�t1�[',v)0a��y�˥v�2�zF��9NbL�+�8�0<9��d��D�@�3�c?�i6`��2V!���6S�d� F��46'��`�<�r�)�'k�~�pP��	��ܪ�ā3qL
�s	�'LJ�c�`��AC��bd�^>|�P���'E�\���8Um&8k3���+ X �'�^xa��N�TK��R�6��%��'΍���Քv���µ�K�j*� �'_���F-3||�c�F�(<��'������-&��Q(ǁU%;�>����'�!ۆ�9'X%�6
�:C
���'F������R	���6%<N�l�	�'�@���KQ��{̔�9�x��';n����?Q��UN>�z1��'ʦ,�&�>fO �a�gI�j���K�'�E��dU�[�5x0A��b�U	�'���1�&9A��Ф�9V�[Z�'�|Q��T�U�'���^�6y2	�'�g�Zd�v|���ݬF<@a�	�'*�!��*
��8t�Ա8+n��
�'$���[0`����*3<��p
�'�:=ʤ�)n�d��Q"wL�aK<9�]��Z�lݢq�<��5��4�� �ȓP |�8�B�-<8�%c�8]�T��'0a~��%�n���<qef��g��>��>Q���y�Z�z��bKчk{�0[��O�����O$$
דm^A�S�Z�p��D+����h�tD��I?H�6���'B18�Έ4�~X��'�Yפ��h��I���-��Ī�'��rg�b��E��癮'W��a�'����l�2t���0e��b8h+'o D�L�#Ҡ �L�B��S�xV.���+�O��O���I�-{��P�v�҅P�,8F�x��'L|8y�D�XӘ���iƀ[>����~��U�,�DS�i˜`p^�!�B�;�y�F� �bM@��*U$�� H���O�v� ���;@�]�������V~�'F2�� UdD�1E�>} Bdc���ybm�XD�����vľ0R����0<	���'�~5��J��sR��qMܬ5e�82	Ǔ�HO�t����'��A1�Q�?gb`I��	y.�>��d��'��ai���%����b#J@��y��L� "'�=�{�H9,�.�R��$}B�xb��	�E�q�J�/1�L�w�|8dm�n���m�3j{`eW��#c�~��r�VR
B��19`���רZ���X�S�;{����b��� lA��H6"��P�7�Q�k�|�c+<4���`NE�v����c��A�����3<Ov��}R琟BJ������O�̼Br�Ϳ�y�.ɒ1'~A�_4�8*"��èO,	qB&ҧh�j��s�!;x�p�Z�9Ҽ��q�$$lO��0f�E�\ �BP�2~H�>����	�)qZ��E�ғ��q�m�\!�$Z��8� �mX*�����M�qX!�DČ������O�:I~P:"
�J!��8j��y�|��)�A�P�Ie���fx06�
�6��
[�S��:�"O����~��傪k����#���{B�'(��%��Sgd��&�
����	��?ar�iFt�*����%{'�-D�R�'��:�"	���1�T�� 	Ǔ�HO���p��!��e��ϭK%T��"O�yꡎ���eӐ��O\�rW�>IT�)�S�~���w�,"��y�圊*d���d/ғu�>	���ˠ ��ۦ �B���ȓQRi�����1L���t��[�J!�'_�F�)��)t�Uj�7 ����f��N�JB�Ir�6�s�&A��\$��Gn��"<Q	�*XM�a� �ȁ]<~�5�ȓ5� x���d�\`WIN8��i��-�,��g��m2�KE%#�F�E}�;Ox�|d�.`��2�@�h������@�<I�fZ�H��y���v6c�@~�<�E�/UG��S�|�0�D�P�<��p�T@'n	q�HL3���N�<��@�u������X+  DH�<!g��	�2D�@MP�Ǥ�j�C�<!�'%|4�GƏ8��UJ��H�<��iA���j���'�0B�JDF�<I�Ɣ�_�ź���KW��3�Vw��hO�O����I�j�!��Ӓ*���0�'� ��5��&�d}Cf�!��u�-OO���@?վ�j� �^Ap���$�!��;� ���_bPa0�"L�t����>y�(2E��A᝝xxjpp�eqX��O�1�$e�w�2�0gW�a���"O�Q{ӌE�LR|�&ؒ
 ���"O�����O�yP%�]:��L�e"O~\��1�]���/氰jcR�8��	;�ѱ"��<�D��͚/@B䉤�����쌟n-����"�6=����M��h��P�l�#g:�9D N`�j�����V�'�󉉈b��Tr��Ҡ���M�|�!�d�<��uɄ�29�p��Sl�8ǆU�ӫZZ�S��?��b�.��T˅�^�ln(! ���l�<A�C�`Ā�(�w�R	��c}E�,��D,�S�d[*��cg��Ia�(X��>�#�� P3@<�.��׬A7*��;D��:#�R�LF����c�*>6�p(�D;D��R+آK�)�'�!߮<ST�8D��#���v;J�Ν�!�	p�	,D�<RN����2�H\b-����n=D��V�[�pZ�
%"�0z �Y�&.D��V�N�e�\���3m4a�.D���f�Ճ9��� ƿb�I �"*D��:���,���!D�	��ȋ��:D���M��c�ni�5.�#Zy�l�r�,D��y�kQ'|y����#!��;�*,D���ϭ}z��k�^��#$C(D��ƣ�|2�
#�P'?8�-���;D�� j����ճ)��%BE��41�A�"OH��A@\D�j0��<J�Τ�"O-#��ڞdVT�ˤ�ŕ��5��"O�]:F�\Bs���ԋ:sشh{�"O����*N5<���	��,�kD"O�(��]�i P\���Ԑ�2�"O��b4	���x���
I�6�"O@�D�E^�n��
C��"�+�"O�I�D��[y`���ǖ���1a�"O�`�WyQ�x� J��Qb�"OX���)7R�I#���/z��P"O��X�gC�	��E{1 ƈ ���ZW"OQ{@NʠWN�s�P�"{�LY�"O�����S�-T��p5-�ӈ5��"O����#�e끪:5�Xe�3"O����N�(~��&��[��(R�"Oz�bA7���ť["6��1r�"O�)�,Ӌsn̻&d���b�"Ovi*7%��{;�tI�o
�����r"O�% PF�(4Y��iۤh;��"O�D���B�:iI��(ڻ7�9��"O,��$�D��1I��
���t��"Od8J����2��2���!KZ4I�"O�Q V��4q�
���I	:XLQ�"O�\��b��p�
Lv+p���"O4���бN���d�U*�4�A�"O���%Os\$(䈍,d
h��0O\,��'�E���:V`׃=�����	M�I�jV�fi�qEɁ*�<B�	�`����P e�A���!&B�	<d��(H��߃�A�P �9Ee>C�Ɋ%�̥���4E��	���ޥ��B�g��嘶B
��ux!^��B�	�JO���!��iR��E�_pC��::w�<:�F[(A�Ċ�{,C�	�-�`5����Aft�F"
,;��C�	�;T8Z%��<P�*u@�
�bC�	גg��sv��`�V�?z$X�"OpPBt���q��5r2@��I2 �@�"O��b5o�$|��Q�@Ϫw�:P��"O�0�ፅ���aYЉ�p�"�q�"O"��*��{�@=�-�<@��4�D"O�lYT�E�e��EەW�h(�a�"O�M�c�0?�RH��� :ĭH""OFig#�R��@O�M��:�"Ob9#8B��`�/S�t��UJ�"O���ʟ�zp,%������y"�=
�X��1�I$=<�P(�'
Z@k�b�9f��s�8\e��'�*�Mt
�K��+0|��'�����ή{���5��j�j�'�x�1�мYs�8�'�K_�-��'�p�3r���B��N�A�mP�'�n�8V��.j:|��R�O-�]�'b���e�S8���h� ��K����	�'$��g��:�ph	���VѨ	�'� y�ϊ |^�X����2ZzB�'��Pq��%��B���@4T:�'��؀�\�s�\D�"���xۄ��'�`�ȶ!SRU`����$X� ��'(0��`�-,����4JˊQǂ���'���9B@
j~L#
�qR\x�
�'e�Q��%���&Ui������
�'�F,���K	p�р���t�HC	�'!0h�t���2\E�W��;c�H	���� �D�� ݞD"<8��J�dzB"O��`	J20�XI(A"�q[8���"OҌR�ȝ��A� ��0ۦ"Ont�3cX/^�Δڑ�E�a��X�"O�l ��9��-�&��-_tmJ�����#�ʚB�'���8�h
_J<�Jw�?9JR��ȓ����V�9�L�c ,��͓8dѰ�耥m3ҧ�����O�3:IX��hMR��yP1"OR)����vn�Y��������W���6���	X�B�.S_��)�
B�l��P�V&��$�7�O�4 !K��G�4p�tn�c�I!�GVm����4��N�C��^<��C�Ɨ&N]��U$R*��=a�a�|��X�QE	�ҘO
|�����D��f��YG
�
�'@H 8�KPad��%[2/�%���2�
���Ɨ�P�1�*O?��2/�N����,B��4���bg�<9��'y;r D&Ȓlv�$��by2�И%G�顳,Q@�ax"�v����/��0�8������>ѕ#�$��91���w�NpC'E���`1����8���a�'H���p��'C�D�3�#Gz�����+�4 ��)P�&�b>Ia)C.��|2��~W���$c!D���0]"0���V�P�T�1z�$�e�C��f���>E����,_=@�J�R2z,
��@,�y�H�%mK(�y�C�Oz��������ɰ"�����_MX��(p�PV����` 0�(R`%4D�h�B
�
P����}��-�0M3D�#�H#b�闢/# ���,D� *5�(e��"!�DR��j�l+D���p��$5���5#_9명�ei+D���g��1bb�p�뛭d0��v�7D�8�H\(k{`Ƞ!�V���F9D�L"�d�88�@������-�rO3D�<�R ��U��1�U�5��j�A3D�,���\->�E���hd��r�-"D��R(����B�-}{��A#D������K.���D%V��\���-D��!�C1hܨ:p.!M'�|JK*D���j�7:������̐m�Fh��@<D��PPGIl�2l1!M(]����:D���� c@��A��
��bޞ;��"&$ިvzӧ��BΘrZ~�Jp�J�S\���f���yrˍ�VZ6(�0�^K*�D������y�%���䅙��Km�y��*IMR!Sn�J1���R�R��=�4I�/�&m��IT�K�<�#�͎�N��IzA�Lupx�C��3$�h0�*7��큥��,!��v*)��4B�^���#d
��#�	�$:Ժt[����b�M�7!򤁴"*Up�J�*2Ꜥڤe�(T��"Sr�̙r�n�j?1���O0p�DOY(rZN`i� ?b@���-D����PYנ8y�ʎ�0B2�R3��OѨՍK����h���+��<�k �5�\�S񍛖v��J�$]��`A����BF��a+��h�Z�Ԧ"4�B�[mM�=_T4���Ao�$�=����'�B��2�,X�T>�v����P0�K$(T`,��~JS)}��S/T/���Q���<��G��<�J�jߓVv�a1�{ݞ�zRJSe7�4J1���&���-�&���1�	WP��4�&Q��Måύ!>!��B&��/d5j���cFB�<A�C��9�<K�H��7�q�#H���9�CN�A���R�!��>��6C��=�2��S����є)��0��/�$<����dN2X��|���R�����GR�@��K-p0�H`�Xފ�6F�=U��'��>�	><��Q�feE�b�$#qJ�
h�>��qq-߄{tXA��IO�i}���g�;k����0+��y�]���C�_����D�4ҚY��&��{+>���ELo��Q#�-�6Yiر�OT�ӳi�Ҹ[!�=?���B�շ�M�
�6g�&] ^�\0�0�b�<I� �<�N�x�׃'�����8����#-z	�ILhv�E �<ϛVDŭK6���3�D�e�2A��
K~�q�'���pdVR��oZ6��T"�.2C|�R�eL���Y��ύ�a�x�-O>`���F�j�1�1O� HT�t�$T��a�!h��6#Yr��$��H$���	F���O'$u�QhI6?!Fr0m�7y(M��bJ=��H��"���<�i��'��m^�8�r�͝{f]��i)f�~�ٵ.}2?��ٸc�"Z���S���J�������aҷ{k(8�@�(�!�[���z"I=A[ I�*QR�bܡ#���{�%A'�A0M<񧨋��'Y���y�o���@��uW���}b��1X���oء<`E2��Y�A� 1t"��^��c�()4BY����ē&�h9����d�rX�#��2�t`FxBf��NH6�b0�	B���0�ٴ86	
G�ˎh]DC�	^�B-q�&(c��᫕�P1�hT���"~�ɡ]P�s���X���k��R�`�XC�I�:?�<���P���CB�uK>C�I^;�TāW?v����g��lVB䉡p]n�{P聪i��U�Q��0��C�I�=$|��ѩ"���B�K�U-�C䉀{L8�y`B?rFD����>Z��#;g�����s�B)ӆJ����4�B�-'�)�S�p1�(4�/A�.�!�˳D��C�ɱr#��Ⲏ�6��!aRe��#$�'�$q��! �c>c��QdJ)Wܦ���Ł<H����6�Ob�31��]ZeZUMU�.8ءY�OH� v|Qx��&հ?q I cT�y����F�n�(�H�j�'I	��%JL?Z�JL�\Ĩ	��A�`,��P�H+%�Ơ�U�'^ZM����g���
��F��&�'��)#DEW�#:Ƹ��>i�,!Hh�Aɟ�m�E&��,���S�EF�-+�A��"O�إ �(�RT+�]��h@L?aP!�̘��'Ddʧ=Wf�#ꄿ��ݑ�V`c��׍QQ�h�S�	�
��$B=AM^�:�%�I��"ej�H	�tE�'PVE��ΐ��԰��!IR�m*5�Q�J�Fy�%�<�nUI�Y�ڵx�bĄ�O�ٻAm��b$�5�}�H���=�H�i�)��Q*�e���=�<�
6n�u�.L8Qł{8�Hs	�	��u �H%Z��؆� h5��nK>�� %�����4A�W�*0����On`��;����f��/���C�5�䪡"O�}��N��������J�� �5h���IH?��$��]��m�%ٟV\��ǧup��
�w���G�@zq)�F�d3&a�	@R���_��&!řk��0�W�$����ќcV�Y����0ij]"��̃}��Y��N�Y#
��j.���6"�b�V�E~b͛S�&Dc��O��{�0`���K�V�=����G�Xx�M�n��,R�E�"�J��DW.*����т��OJH��aGX9Rp�Bˈ,L���DX?��K�YC��0�jE�#(���S(��-
D>�ʶ����k�E��y2	�6P`�""�I(��!bb1�M�&�L ZD����<=JT@rf�Ro����J��O�H�íT5*V=h����"JL���UPxI�� ��;�ڽ	G%��	�=�e��+��p�rP4����2[�n<�P� �"�Z6�(�3$!i���1����'�� ã�MӺ��|�3�Jݠ� ��$#8��[�3�\��S
A�WB�|j"H�6�<��er%�e� =7����Xц�v�VXQ اO�)�,�.&��4�G&Y#S��]	b�Z�s�G,T&e� M��e�<W�Е{bǘ��y� ִ^}rͳ��ߡH�ȃ��yfY�u��?oR��4) >p�A���V5\wj��v%��ɘOC����/I1{@�A�!ʮEf�ѫ�#@^L�r��b���	�?�B�YPO]��0��*�"Aʱ�㍔����kC?c�\ґ�=���fW5(��<�VeY)Id��@(N�ٸ'0BA`��Q�0��I�~"��/hV���pM4c&`�镥ѥc�"pK[�	��ls��p>�2�ɗOZ��!�iC�%�]�zfy!�K�/���'�8خ;&]8e1'T�A��{����?�1-�P\ &��''��i�dj�4j�D��ȓK���C S�~; � �²
��o��uet��o��E�h8�������	�|9"�>��@U�8����,ef�Xf*6|O2��r&���$�{�8��ՠH�U��ya��/�Z,�(�\y��Y.��}&�8Ӧ�O1t�,�:�&�`�f"4��R���1�*�h�,"�0�@���j4��l�0�a}�B�Z�2Q4�]�S�B�i���"��<Y�'P�L�A�͢>�w�m�ލ��ޥ�e���DN�<��eR�N���B�$r-1g	B̓&z9#a牂������U� U�0�Hی�҉��"OR�U�50��j�(�p�2ā1jU YtqO����Y���5DO<�q�CMڡ�����1D��  �Q�:��,)A΍"��iZ@"OvxÐ�&K���DK�9%J��"OHd#$��"y�x��vй�"Of�k�E��+�h�ЪٳE���"ODq���Ch��F�@�8���"O����gT^	j'��j��"O2P��>�Ȉˑ,Q�1�&�"O�qb�oX/_0`e��썑b�vR�"O~h�O�?`g����-�`�"O������q���I�V y��m�$"O
,���4^|f��g��g��t�"O�Ѳ�d}�x�VE�;pT�"O��kf.E�N3�l�D,ԉo$�u��"Oȵb�K�(�*U�ݍQ��Bc"OAC!�NI���JأhW�f"O��CWa�`��Q���	TC�`�U"Oą���$�j9��) ,Un �c "O����M�y��Y���a^�=('"O&�� *L<"M�*�Gގ{�hM�*O� �a���.�KDL����$��'&���I&c:R1��N��!4٢�'�P��D@�%E��ls��ЙX�x��'�="��ݠ7b@���ͺi��`�'�p!��a��a�x��˝1-��'��|��eQ5_d�q� O l^.��
�'�Љ�U�SQ�J�`�	gv\��'��L�G�9�Bh�E-غB�����'�b��q��v�n�
�E�68�d��'�P<[�)�-g:�çn[,
���	�'G��0C�ϤQ_��#r&Y<yN����'7@�Ra�

`$����rSΠ��'U��U�oF�!��G�����'����e��6� ���af�Wv�<I�(ރTb�M�c��:��	'��T�<!�TA-�*�a�?BX�=B��H�<����3�t*q�^OR�H��@�<)d��^*AJ�Aվ2H�@��e�<q�n��}Â��!ǹ�b�@�N�t�<I����*���c��?tp�����}�<��L�/�|L���;BoXy���{�<i�.�?u<���kN�<������q�<AA�*s�i�tN^�V�>���$�Z�<!�C�F~z��C;6��R�[l�<	����s���b�ˏ�0�B��C�<�0A�'wNl0P1��^��\��Kd�<A�
C�d}R����TQS��}�<���3���k#^�i��xSKt�<�QǄ<@�
ɦ��d�1�TN�<���I��@t�L�t b�T��v�<�%ξ9bb�����S�f���_{�<���]�A$�d&΍nh|�@F
�t�<yw��LK�&�2D@��6������b�X5�(]�2x��R�"�F�ȓ!1�Q����1�
�6�>yN�܅ȓA�4�ᖃ?d�K�#�O���ȓd����\ke i�����`��� 8�ȶe��=��9��;y�P�ȓH��9���*R��%y���5}���ȓY��L���K8`޵����2%�q��X��X3�V��@��o�5P|,��!EI���<Vu0�g'7�l��ȓ~^*��G��3�NH����dS
�ȓO��=*v]�g�L9��T�=��r�j��eꀸ^I��p"��r�Й��S�?  �˲��5�4x�ыE�WZt �"O���"�ܼ�pפ�9/$<�#"O�`p��PQ�\@�"E�#c���"OBm�2e�ut X�V���a��,h�"OB�S�F.:���Q�D����|�"O�}�􊅝6 a0���y?.̩B"O^��E�^:�8�!H�P�r�"Oh�0��9�0xZ1ᑙ�����"O���,�3	&�@���x�c���.N��4�� R�L�x����L?B�*hj$�6E�����iB�Px�Nޏs��8���2&vZ�7������"CLҧ��2x u���[|�Җ�iZ�h�"O�h�)NE�����M�,E�icU�l�vbV�5�Y���U���(�%h89��5��]2vF5�O�M�3o��Tp��ąq,�Q�K�e�����Rd�HB��ZL��'L J��Lc��M�z�=�qa�sp�9s�dҢ��O]�|q�]?��Ec�.Ș!�d�J�'f]8�e�!"p��"���3�$���bYX4B�g[+$>�++O?3���>��ip��X�8t�g��n�<�ס�%G��P@��,T@�L����~y���0N�H1I���a�ax⭅�:>��#�I�KZ��x��Z���>i� Z�<�N���\u��1���!O_�8I"Nw�q��'��e��%N*+j.�r_�I,hͳ��䒥i_n}��*
I:�b>q���?[�V9��"G�Z�$|0��3D�զM�z4�5c��6Lqڙ#�r�����t�:|��>E���X7#L��mH-����F�S2�y"#�iXa�GT%�@�Х���ɨH��؁�oX���qF���|rӦWj"Y��1D�@k�ò`k�xҤ�F��I[W�2D�4�V�]�z	�5ڰ�޳q����#D7D�@����
╙�G�=�h��uC;D�$�����R�T�QQ+ܹh�t��<D���n��6��Lڶ[�w�,J�:D��QC�ϚN�41��׸!9:��1'9D�Li���;6������:c��*�A D��(���)y"�X"� Y�L����>D�xs��Z�C�,�p�a�#C�n�I=D�l��"�A8Ιhw
�\,��
$D�x��4Z� YkNF�Y�
.D�(��X�2� MY�^�&k���d(,D����
+��赍S�Y���1D��s#ٺ=E(h��]7���V�(D�8#�]0}��L� �Wl�����Rk��
H��~ӧ����ˌ����H�y��᠂��y���N�<�z��u b&V��y"��)Nt�8 �ҡ g�y�	D$)��=Z�*Ѯ`��q�ˇ��=f��`�d`��ĥ+��� �H/oƀ����	���Iӭ,$����#��l�Ǖ7U"���)��tqpI���0?�5����x�����O�2�(J�CБ]�!�d�g������J�,abS�[&%�,� v阨LŶ4��A�f?����O��q����-B�J��s�̡�"O�|�Va���l�񳅇�
v��?�`)ҍE��й2�\&g2��$��]]��j�a�)>G(AJa��yk�{R$ҥ�xh�w���XZ4%R#�%.� cC���G�ܑB��"4p
Y���d1��(�#�/,��G��%��AYgf!�	3*�� �G�7=*N@B��i��"*
 #T�
?�(��ի���2@����"|O�#��3M2č���)��y���0!J �T�M��8���'orP�T-��jv�7�K5Wd���G1
.R�Qv�T�!�DF�Zi��@S�^��7垏W��f�>$��u`P�~S��8u
ǚ^m��O�ؗOh�qQ�ޜ{�r���*U�@ߓ��1%��Gm�yYr�� ��Ik�	ȫwQ��D��O���aRn6e���'��>�I�V��P�T��$m��s�,�°�lZ� 5S�����:1�v�jR�
�*�`���0���2F*�('������"o������c����K�j�V=�2�L�2�R��FͿ+Y��O��{Z�l �+T~����Z*�M� 橁�#��wl����]*.�U"O\��W"G!A�h��Z�0*� cv�''z"���.㼑2B�0b-H��"G��`���'b�����!�Ɖ�+fԨ��2|m�8آL�`ܛ��@7E��[�B�4�-�ճ
�hk$�=*f7M�: T�*����#e���:\�t���,�O���@��A�8J���0tp#d8=����VJ�+����!ƵUJҜ�s�N?m��{)�L��Ay��8>e�b!R���h�4�t��'�_�+� �Iw�M�YA(Lz�0O�Xz�;1�6QH$F@D?��0`"OJ�x�/Q]WB�����O���*��'�-��eՊyx5�����ē��RH|z�fҸNn`zf�|��4�ť�t��T���_[v]k��i�dl�Q�Y�Z����Rf������&�	>�����L<1tm��miz���)\a�0�0b�u�'Bܚ6H�v��>����+��x#C�G6�؉�#�;D�PCFc�>a�ZPI&K�?5�hM��(�d6B���%�)����T$.T���"��&-�^E��A7D�D�����1�<���ϑ� }c�6D�t;���,?aB%�b%ʔc�*5D�h�ӈ�
m�"��V,L��j0�<D�py%M۾>B=1AW�^��V�4D�D��mW(Y<�=���`�j��u2D�����y����F��q�nA�0}(z����=��Ǎ[��x�JԮU���r'�j�<�!��3p�6�E
�*??��
�$���q �c>c�X0U����@Hqs4�9��,�O�P5 �{�q ���V�2�#�
[�q�G�����?a4.Ѵ$��A�Ù9p0�1r�]x�'���� L�ܑK|
4���$]�%�̗l.R	��O�<�D�I9pX���d�j����-Q?��D�$��e+4�F�����'����6A�Lu�EH���bäB��
h�����L�G�`iBA��e����.Oq�%%�W��Q�J?��w�K4�]��(3l<9kV�)�O�A[B��(�HX�!I�]\�`�!I?:�Z�������DSMv�\�"�ÇS�gG4h-Q���'ϖ.^.Tx��p��f�~5�f���$9�L���C��7?�Y+uH�7a�5I��
2zkv��)A�L�i�Q�՗�h���P
�4Y�!�	-}~�z�"O8ݠ5�8#�J�)�.�;`E�{4�3?�D] rʞ �(0��b'֦9�;���"43��S!��p?�c�[���Q1�?i[:�s�D��pi�RG͝�B��*j�R�(�'���1ʃ�q�R"?Y���F44� ����� �H���΁".�H1P���y"��Z>4�hcB�2��9C�J�R�>`��c6$��1c����F��'�p���TbM��@�6@X���'�"�x�g�z�µ�����)fe�ڴ�x�/�8�p>iљEg������4��8�/M���aW�Ō="B��V3O��Ag��|s܂�W�Uw�qC"O�]�шC�!��Ѳ�bllL˥�DK05>�͂s,Z�ǈ�qJ���

����P}K�Y�d"Ox��ՎF9,V2<��*�&N�lŠ1��]�|��B�>��(��l׫�<��'z5���%]c&�q�E����Y	�'��l��)Y���� �ƭj\@J0���hvh���͌�h���f��ɧ�O5|
`�C(B� ��'�@�~�	"���!S ��G����{��l�E
ȶ�����㙌W2�nM���3�x��O�|s�4�p��FL���rd���_\Zb$&���h���b�#M&8�|���X�nB*6�Lғ��6�>���ش�.%"��<���jބQ{a�r�����i��2�]�E �!���Ǿ&��D@E�J�t�l8R%�t�!��F�O�0e��G�|Y�lأ�W�G����'.w�鸆oq���R蒌��)[v��Wʕ���PJ$ʅB���$��uC�T �Ot���ePpL�@�&f*�h��F�y[إOP p�,�3}"k�ג�S��C5$|V���ϗ��xR�˾U}�c�BQ�[�@��P���A4��uǁ:r(݆�I`��X��E2[_��`�,O�k����ŲYY�Xм���'2����e���0a�OB��.��	��� L���,R�8�8�˛`�:���b�0�&�$��1kDD.�:Y�L�b��<=�ڨ��Na!Deۄ9�zHI�D89���4�Qr�\�|�'��@q�U	��+� v��Y��'IDex�Á��2�X�2̒�'߶|�0�� �24��dG [��z�'J6ʒ*K�i�����iΩQKԡ��'Q\|z��
]xjh+v ��S��=0�'P,�R�%�?w�t8��Ԣ����'����		�AŊ�de��<�q��'�r)���sw
U��a��ȇ��'Ć�3&���qD�5 M߀H��'�"� �!t2�*Gʔ+zah�'��`�#�G�H��j�ʬ/�,��'VXiK���=�X�nm^��'8���k�c8B��j��M�Z��'�@2�+�B���1t�^;)�E�'#J�
�H?'�,��0K<,.h��'�^��ƪZ�	� �*�/�XlUh�'�ZM� Ádqdb��!|���'|6����� k�Ⱥ���':���'��i��AlE%�aR��'D�l���-6�p�Də�J�կ:D����-�.��j�M���6D�TS3��Ϣ�� ꍌ)��e��8D���@�R6{;�����<8���J�)8D���ʝ'(8l����5�iK�h%D�$��L�t9��:�jڐ2y�����/D�(f�U,K�Tɋ�$�"�8k��!D� `��� ���GOԡd��8�a?D��3C��#>#����EYv��F?�y�A�X�� ɂ�Ҽ=��j���y� L	I�Y�S▋��8�3�
��y�C%lhL�YA)A��M�rH��yR��;y�){e�ͮ5XRu�n�*�yb'Z1P)��"sŔ�)�h�
����Ohe��f�<����ѥH�9O��E"O�PP�Еz+�q�S#B14J�"O�P�
ʪr�:����89-0� G"O"��*݂�H9*fb��h"� 9�"O|��T�X�&ؒ�o��%0"O��r�o܍e�uCP�H�$��4"O��cD�,!�p9���)zX��"O.Q:7d��j�eNYQJ�\ۆ"O�4ja���Y�4pCʡrQ��J�<�2� D��c���2ZB��(E`E�<�4 +)�^�q�2'�2 �D��}�<����5������^{�ux �D^�<�`+Y0G���C��L���f�c�<��%�\�,��rir�xp6��b�<a�%]	p�їN�"V�ؼ�R�g�<�Sd�2y�d��5��� �VCa�j�<����ڊ��c�� m嶸J�Ś@�<ibbƤM�L��̎�<�^8:��X�8�"S�@���M�'��7^f�ː"ԈF�A�'�F4�?�u��1(@�`��Y|�l@��#}�A��eKvf�1o�������� 6df���&/?E�.L�n�Z�˃0KԠ��6M��p Q��)u/�8�'��O`���ځh��#2���0�^�\��Њ]�<5*���>Y�j��0|�p)@?_i����9�)AgZ�� ���&J�O|��ْtW���~BN?E(ֆA�SЬ�*�eŨq���۵MblP3=OT�W�:�)�S�{֊�b�
�F$`P �><D�B�I�y�(J�Fٌ7�Le����0��B�	'I��b��M*^����0��(a��B�ɕv�"ȹ %�+P�<�U�d/�B�0o��D�Q#�.@4�Ġ�LrB�)� �d��ĴS��(�� 7/�I""O����
d�p�R�o�"�m�f"O�|��@.��|SE��"�����"O��E� (��:��oDR�:"O�h9���[�pd�ʙ��x��"O�� _�a�������)^.(x�"O^��Bͦ	R|s�b��*[(8K�"O�q+��Ϛ>��G�ΎUL>�!"O�	��D'R$�C�OkS>uȳ"O0���$s]JF�$x�!ӳ"O�{�b�8��-_?�a�R"Oeq�L�LVh�6��`�"O�t04��r��,��E�p���3�"O�l��`-�~����$sE��`"O�|�N�{�4���N58�5"Oa� ��;.���iCE�쭰�"O��a�i�@��]�eJ�T�� �"O��S�X�,����4k�:���X"O<aCdFO$
^ƱG���,0E�""OبqS�V p��P�Ń&D��!hf"O��W$ܩX�,P��0&5�"OZ�zg��:���5��`*�"O~�za�~�̸J��$S���"O��:7���5)��B��-!�$ǚ�h9�a\�^Ub0{�@��K�!�$A6=�smP8>Q���#@�:&�!��X�jtX���{<��f/�81�!�7Nt��f�-�u�o��!���i�]�5g "�[�Ȃ�n�!��G�p�fN2W���S�&�!�آgfڐё�4���\!�ĉ�nK��ţ �D�a`  D"!�� �^]\�m��JHġ�3IM�<!����L��''\�:B�A��
�?�!��L	g]B��SC��d-2�
>�!�
!�Z�§
,j�@�` ק8�!�)�pQ��I�3
y��dI�3p!���yg� �цV9{W�؊T��)e!�D	*2�楪��DML�	w�N�b�!�Մ澽��D��>��Q�n��g@!�D��<!��F�&9�#'(� #!򤅕�2��o���"(�?!�dڬ+=�\"B�'�D�s�V8!�W�v0L�q��݆:А5�Uk!��3GdF0�u���!p�C?X!�DȊOK���f�ؠ/�t@딾8B!��
D0��t� ��]��J�&)�!�d^:c�P���)��~�l��')Z�Y!��ˍf�@M8AE�/)����IA�#
!�O=b�&9�X;b�6�y��1\�!�$� 2a��ȥc3ڨa���G�!�DE��V����A�_A^�"��D��!��!��9�#C�K_�H+2���s�!�$Y}�0�4GD40R�I�Fې2�!�D�68�x�3�ŉ�o_Ve�G��l�!�#]�Ӆ��-/^����^=;�!�D���h`���i�X@F̛�Zߡ���.k+tJ$%��L�VI���yR$�U�$R"�+[Z{"Yb�'�����,R
>6�i��C�3U�V���'�f
'�!CpT�4�J,Br����'����T M0F����Ά�4xft0�'u6��۰9�x�&ؔ��e��'�H(�U��&�����JM"�t���� Ly��JV?Ő�8��K��4�1"Oڼ��J��j�~�#,�R��a�"O�8C�N�G Vh�� VC~ @�"O����!5NF�|���N1ffQkV"OB��Ο���� 1���"O�lA�vCPг� �c��6D��ia�&0v��I�(�8���5D��"&�I4l�� ��EIl'fș��8D���"Lf��X�2C�6.{�`y5�)D�l�VI�x�\(:�G%A��@s��(D�Y �˒ �x��.a��i{a@*D����L�-7��)R�7I�U�@,D������-�Zp�QϿ{��z�b<D������D
2��^JJE.D� ��`ՀUK��p���v�v�hDL,D�ܒf0�0�?	a4L���4D���E�ؕ'�Y��FX1 ,x�e�0D�Hz�Ie�&�k�DD9��,!D�t�Ы���T4���y��1�a D�(z@`�S���V.P�r��kF�<D���%_*P���������� �>D�܋Ԇ3+���	�
�H��Rv(/D�,��l��C{JT��M���"/D���-ŞH:V� @���I҆-,D���0�D�I�t��$�(Wy0��(D��	a,Q=u��50P�d�&/�*v�!�$�&-)���E�\e����Mۏi�!��� N "9je��>"�	�"�%%�!�d�4Rɴr�C�9nذ�[ ��,n�!� �"�0	�"���ۗ@O�a/!��̊i��q����3��\�So.�!�L�h��I���
�T��ar6�@�/!�O) ���,Y�]�Ƽ��.�$�!�$E�8^ɡ��9St�e���}�!�D�u��M�Am_|V���A�z�!��f5� DJ^?<]�z�'��Ux!��G�l�~p��O�pL p�DL�pr!�D�?s�:L;�I�i�w	c�!�dP�(EV�JF���^��т�@��!�d�X�0�(��A��fd�7��@|!��8/J���X5�dq��$�VB!��
	<�[tcM�Hu�{		(!�䟾F1x�ҠUh���D6,!�ڦ='� ����
������W'!�$�[�6�1�a-. x�hV퐾7A!� X���I�,ݦv��1�➙)6!�䂳$���"V06��=׏�"!�$OY�L���>d�|�1nҘt!���n�"8�'͘Y�@i�#��P`!�$M�=��2ajM+�j�X�	��|[!�D9al0�R�^N�]��&ư�!�$�4G�{�d�&[�|��d$�;{B!�)A��y2 I KȈ���LL4e@!�ė0(\���k��P�05x�œE�!��A�̠9��i��q�Z�F�!��ѓ=��H�!�Q�d��FiU�)�!��,HȔ;f��[r�-�U�ѽg�!�DT�@�&��eN�Wд�&��.!��W9{Y8��cUp�y�O��r�!�c�ԈhM&:��t���!�D�� ��*$'2��01D�ɟ�!�Df ��r��^@�"��`���e�!�d��#�3V
J2��-J�J+!�$ ҍ�Hw��!��Q�{!�� \���M�.� `�Ңr�&� "O��CA�F6�hy��!@ M肤�"OPq��.
��1��N]`�"O��j&N�L��t BnΥQ��zF"OU�r��Z�B�)1MH4bo� S�"O�xi�ȝN�uU�ϱsi���"O���h0F�+�ʗ	1[����"O��`7�ǃ��8H�iJ�}Fp�ђ"Ov{d�P)R�n1��.֋q@�$j�"O�(�G�B�+�rIr����~)���"O��d��'VLJ.@ٹ�"O�PۧDü/pNX�QP�[�"OrD�F�{M:m2gH�/BBlq�"O� b��#$����P��1<'��r5"O�`�"��eB��� �X*T�"O�Ы�j�&P�Q�`I�@Y(r"O\��5���p�er��53F��"O@-�߳G�5���7��#"O���Կ2��@ �O�0� ��u"O���僙�&��<���ʸ�I�"O�����$vd��pU���F��"O����<vbث����Ͱ�"O��%@Ыn��|��J�ˤl�"O��M��EX�eڐNb��)��"OX��gMġ\҉R��$��<�v"O*��bn0<:�C�����-�G"O*��` ��,ԐPM['mZ�]A�"O��r��rу��I��	�"OPX5iӃp� �S ���
prw"O��C�$�A=�1���!,k�"O"(r�'ĸ5a�x@�c�� �r-@G"Oh݃��U8��2Y�9=,��"O��[@M�	J��)�&ݏ>�x "OX���IU�3l��4T?F���"OȀ�3�F��B1���Ѣ���A"OD�K��V��)P�,E�~�	"On P2j4U�-��
�UE�!�yReZ�
DM�I��CN��y�M!�Q�G�7u�U�F��y"��5G��k�
K�F�p�h7�[<�y��b=
���7E��Xf`���y���(G����a$�<<�a�Pj�#�y2/�,�N�k������͉�y2�H�uV6��a�F������dL��yD�6e
�lxP��gf���uM��y�	����E�����Y/�y"����f�@v�	�Y�\�cO���y���xڠ���<�r*�yr!�SLx�KU����~���+��y���O�e�*�:5�a��J�y�e4�$��-��0��9 ��@�y�jJ�Kl�P����=�H�$����y�ǓJ�ݪ�dX78z����\�y"8}t ��d��8/q^uz3�Y��y� �sc*�Z��)�\�ђ)�%�yR@��1:�t:��%*E�& ��y�Q�S 0 �l��;A\Y�9�y��M/xq�OG�8x|�pE��y�"�<6E�boQ5v,1�X��y�G�K�p��̍='I��0U��y��;r��1��U�Q�d�Q��y�<9��1%F�TC��Sb���y�(�l�<sg�!�����C��yRaϚq�!�4��>$��W ~�Dȇ�S�?+�ş   �   �  <  |  s  �)  5  <@  K  �V  �a  ,m  'v  z}  `�  ��  �  4�  v�  ��  ��  B�  ��  �  L�  ��  "�  ��  �  R�  ��  ��  ��  K�  � �  H �% - �3 %: g@ uD  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�Y�G{���˾R5$�Qb+�jBƅ�7��Oi!���l8��Ӄ]*W>�\����]O!�ė��ތ F�8#"J��7Lb!���P~��#���(%l�(.ԜoI!�d�0c>��=`�r$,�
�!��LP!���6HٮsX~��!ݺ�!�Ĕ�m��G꟯i�̥sQ �W�!򤃛]Q���D�o��Z`A03�!��R�6j�l��B�^ ū@��;Ol!�P9��$`b��e&Ī���c@!򄊡jX�QTυ#i��A(PhˢF"!�D/2��`pB�]�6�`�6��9!�dEE����BݙB~�tK�`I�W�!�DV�=�i�H�!(^n8�䏔$g�!�$��mMX���9OT���n��O�!���-
l��WoР>J���NE�ni!��K�4�VYP�ɑ����+L�xT!�$�4<{��J��! �PhX6*ʨI�!�Ff^��PR*C�lʹ����F!�ͪ&�����'�4j�\���(�8\!��/�:��������bN	i!�$�<PⱫ��53���{J!��@�S�vL���?ʀ4sW��*t!�DT��`Iȧf yƬ`�c�]�#�!�D�p�,l G�.x��ᲆ�T<@Q!�@7_�����=�"|p0��-N!�"F^�cbI��i��,�g�:'�!�0�@1g�żm]�,�Ҭ�
3�!�d����(�qKrأR+�<q�!�ںO`�i�눏`�p�5mܒ<�!�d?B�>�1f��~�>�#���0b)!�$C6h���@焐K�и��)4!�� 4IAI�R@`�g� @K�C'"O�ِ��3|�V9Y%hS?<v��"O�y���<9�t��'��X=�"O�a��Q�/k ����$�Lu��"O08DF��D��6.M02㼠���5D��")U+e$l�ȶcX�6���Hu*8D�T�N�,N�n��4h>~��ǈ+D��@� Aƒ���eT�VD4��%D���q'�
1��Z&�Q�9h� 6D� ��a��1k��T% ���J)D��(�f�4��US L��1�z]���4D�p�3ϐ�ѡ��R/BI���&2D��I��.��s���p�� -Y����@�Ta��ցE��1 �oÓ�y��SZh&/\�SIRݲ2��y���(@��Sʀ�9̸3�j#�yB�ZM�z��?~�t�>�y�NÙ[8,�kWG!hQ�\�C��+�y��/����C�úkl�Y�-�yҎE G���롃�f�P}��eɱ�yBbӣ6OI��G�s�@�a�NI�y���(�=�"#�1lu�l�7' �y���8l<v1C�G͌eI^yD犠�yHг w�Ժ�=S]��������y�c�'�8*QE�K߾ț ���y�]*�������9,�ٸ o�#�y��M�j��D�2|¤{�G��y"#̽���h�A�a�Z��1Ů�y�)�s�0	���\Z�����yr�	z�H���+1��	Pj�3�y��XZXt�-�%`��ʤ`%�yR�IJ�P�����XWI /�y2���U?E���Ԍ|�j�!���y�c'�V��p�P��Bh7�J�y�:v% �𥑮r?l�i��y���T[�)Qg��}�`P1���%�yR���.���8�C["#�v��AOV��yBn�b=�A�X<� ����M�y�eD�_"J���t2a�5�̂�y�*��X`Ht���:�xED���y���1�J�Bc�"��,zu"OH5�5����\�B�ʄA��=��"O| [A�Ȯg��c/,�,��"OBy�hP3&>(��AI*�H�s"O��Ru���d�B�@(�&���"O�j�"�	�S �W�0�P"O������n[�}���>K�Ь�G"O���#��q�)ڒ@#Gt���"O��S��CT'��kR�Q�11��)@"O60�«�j_���hٶ4#�"O|P�d�I�j@@�2���4�,"O�@S��W���@�����TwB�(C"O��C�C׫Ix�Qi2���H�X�6"O�ɱ�dZ�{��ͫ�/��	l����"OY�!/\  ZR��BHW)+pD�ٗ"O�q�@C�lx�#cgިk���P�"O�lK�&T<T�����o�t�2�� "O|iA�,���٧��#&�YzU"O\ȲX*��9[V�C��|@r"O�-�Q�j ��	���`V�lA"Ox�ۡ,�:m�d��qJ�i��h"OD8bC ��\��c'/0f���)V"O� �/<]���z���F:z!�E"O^���'�����+�"ԋ$(�S"O� �x{U�jHXAY�̓v�x2�"Oࡓ�O�B"؈ �Z�6�1�"O�Y$�ِ$���RS���>-vd��"O�����?Kr�HA���X�=��"O4A$!8<���M��L�`��'z��'��'7��'��'��'tj�1���<w���G�B���'\��'cr�'?��'a��'"�'R.@q��y�|$�QՁx�ځ g�'��'~��'��'�2�'���'6�0�M��
���U��1�� p�'�r�'n��'R�'2�'���'�Dq���+K>��`�3������ş�������џp��ݟ�����4qlڌ^Q�<��W P�t�ǂ������ԟ(�	���Iʟd����\�I������Ԫ�^�h�c�I���3��P�	�����ޟ<�I�,�I̟����h�7ɘ�!���4&��W�����JΟ$�	ڟ������	��	�$��̟{�f\�`��<h�c�� �x|��iP�������$��ƟX��ٟ��	џT�����I�Ε�!�����P��
V����D��ޟ����@�	���Iʟ��I��|�&��D�d�r���>�D�$������ ���0����d�Iß��I��$��6&��,H��[�e�6!W/_���ş��	џ��	�t��ȟ,���,۲�%M	����[�ТZ��Y�������h������	����7�M;��?Y�R��"��8a �i`��0k�	۟8�����d�hG�N:`pLC¤׵����&K����_3�v�4���O>�&��O+
ͫV�� Wɐ�����O �$ڛl�07-+?a�O���5�$�<iZ�]z�)�=U)5/�)��'T"_�lE�DƷ�h �a��8P��u 6m�0�1O��?5�����@���b�h5��k �;gᕅ�?1��y"R�b>iѦ�S��Γ6!���֌��u&֝�$c�"~b���yrB�O$,��4����-Rg���J^�fL����]�)D�$�<AO>�i�Z�j�y����ة��V�U����b	��]�O���'���'��T>�05Ù���fѐ\��b#1?���bj ���FF̧bk��F�?I���gb2e"��F6�E�� ��<��S��y�,T��Sv�n^0P@�H��yB�|�!qӝ�@Rݴ�������y����\;]��Eh�D�,�y��'���'N��1��ic�	�|�#�O��)4n�!
6�%���w�=å�X��]y�O�r�'%��'3�i�3J^�<�W�Ւx��dC�B]�R��	!�M��V��?����?�M~��}�n���G��rS�4`�ǻ�Nu�$[�������$�b>yr�O��0f�X���
R`�3x���mZ|~�*Ȋ]����������;�
�j�#1�0��$�.;qf���O����O��4�|�
C��Ǖ8��-jN��	����!�3fc��t�*� 8�O��D�O��$��I_��ఫШ1뤔�'b�1\�Ĩ(%x�V�!�,�3s2ʧ��KT�S�U� �h- �c��0��<Q��?A���?1���?���o^�Jn�9�F�U�_c�hh@��8a���'���l��8)6�<a��iR�'�aI�� 3�@�x�ט~u\��P�|��'�O���h��i?�ɠDҨ�L�6]���"uIР��~]"��+~�O|��|����?	�N�
��S�l����"�C�Hb�����?�,O@�l�e�j�'R�Y>9���%�X��b�H��6�cw� ?y�U� ��۟�%��'6����'��ec�t1�O�p��k��Uq��,�޴��4��i��'g�'5�a(�F���|�cv��]�v�rv�'T��'o����OS�	�M��L,���b6�O�s�T���(1z�����?!��i�Oة�'t�d��8��H}�Z��V���'��Ġ��i;�	�f�:�����&�P�Ju&U�Ev4��b��fu�D�<i���?���?����?�*�2��GLؘh_̱�!�*q,�C� ��I;u��� ��Ɵl&?牟�M�;L�I�l���BǄ0u4��Ο`��z�)�(p40�m��<93Hڟ-����HE$P����<�"A�8"�^�DT��䓢�4����"X
�h�(�dZ]K0��/�O���O~���<���i��)��' "�'��|rp��:D֐yR��[��9ѥ�Du}r�'���|�\c�]�� 
���1ሂ��$U)vy{�`�^c>����O��d��G`���
�y�:��d��!���$�O���O��D!�'�?��!�~DŒ�O(:����?i�i*Z���'�c�X��]�h�=��J�ce$ٲpĚ5�x�����	�� ��Gצ!�'�,�&��eʀ)SF�iAL��lJ� C����$�O���Or�$�O��	�b��婒h̎$��PE��B��)�f*��R�r�'�R��d�'�`��gfG?IAn�#��[�~�Q�O�>	���?	M>�|B����L�jq�q�Ũqb C�_�CҌ��4��$]kM+�'1�'��	�$@hq[��ᐝ�g����D�	�$��ݟ��i>9�'G�7m�{����2F����� իmP�re�������?yZ�@���|��4ik�4��@S�(��(��#B���tB�����)�'�20��m��?�}��{�? ���2I\�*9l`���:rP"6O����O���O��D�O"�?u�� �-$1��@U*`e�!w�W֟��I�l�ߴ;q���*OPunf�	�2��	�@D2iM�[ �	%���	ʟ�/ƘmZB~Zw��Q[d��\��ϼSUXy��nٰD��L�g�	py��'�R�'���K�jz��׫A�9�@�@�pr�'��I�M��	��?1���?!(��� ��ׁl�|���_'-9�������O��$:�)rf���t#�&Y��N�X	�g�챂��_?|j�eX+O��C��?I�A$���(+t>2���(�Й��O.N���d�O����O���i�<93�i��E�b���Z���J��	�t4��N*��	2�M��J�>y��j�ё%��|���gR�R���?�3����M+�O���v��)S���B�8���2���8��U���ςrH��<Q���?����?a��?�)��pԬA�:Vn�b(ܚa��9�b�ͦUі�
myb�'s�O�R&m��n �k�l��ǂB�����47����O��O1�|�j&,u�6�ɨ;�*)� ��2n�RE[pH���c�,��۰n��d*���<ͧ�?�v �-��P���^O1R�I4��?	���?!����N���E��������,J'����p�ZԫƟqh���b�Mc��h[����l��]�'_� y�e�0lD8cG㍓���`����W�(��|���O���OD��3�֥BlR�i���/0�%���O
���O����O$�}"�MDd��5L|�Y�-=��I��G����/<���'�61�i޵C��ìZf��+t؛4,!�w��æ���ٟ4��mU�9�'fҨ�t ��?����5L��(�)����pJ� [��'��i>��I��<����4��"f�`);���5��v���)���'K�6�Ӕ~t��D�O���/���O��k�+�	�j�r��a.qKG��x}R�'�R�|��T���K?�4+�4P�`�`@�l�ݘ�i
�˓����n���&���'� 1��`QRq�䊶��
]lc�'_��'�r��dQ��;ݴ;4�Y�:�&� i�B��k��&Z٨��:��v���d}��'���'mژj"iF�Yd���e�^8� �*ڃ:��6�����ǆ6��t�	��Hɚ��5#;��jP����5O��D�Oh�d�O&���Ot�?E�-�;C��j5��ؾA���՟��I�P�4�n�ͧ�?���i�'h\��C.�!�%��$��\�uI!���?���|�#M���M�OҸ ��g�И��D�7FrF��al
 	x�Q�'��'���`���	.Q�*��H�D�ԣ� �UR���ϟ�'47�[t��?�)�z���)�0�VT v��%� �R����O����O6�O��;GM,��a
F�-H�q+&�V`�d�st�B�>LvD�"�ey�O��,�	�"��'�ҁ�`Ӝ�88�a���O Ɓ��' "�'��O��ɷ�M���O�T��s��X�(ڕb�,�0X-O��o�o��^��	��0`�ȷ{iJ4j�� *U<}9�oßl�ɹ�$�l�C~��^������W���\����a$x�a�i�)��$�<���?���?���?�+�5��ّP��5;���9��y!�	W��a��"��������8��ŵ�y�.4&�}H�7)�H3��6J��'Bɧ�OO|��űi�d�<"���*�c`���!	�zi�䎭b?��q�' �'��I��@���*T%��#����ƌ (N���ܟl�Iן��'C�7mVG����O���,��"OfaWc+�p��e=�	�����O��d3�d��s�>a��M�\�N��]��ɐ8D;F�P��|�f켟��I)#f8d�~2�t��@ʇ@�&�I̟\��ȟ���G�O'��O�*����	,�r�#��6U�Al�1�E�Of�$�ߦm�?ͻ�5B���)̳�nuɶXA�4Oz�D�OV����*6�$?Q�[2*WX�	-��zQ#��2ڜ�js+­e}`�xI>a+O��ON���O���O�=������P%���˓�R%QT�<ɔ�iӸD���'�b�'��O�"�?4�ai�h��zb( �f�2 J(듆?����S�'|F1�%��JCkT6d�N1r ��MC�O�JĈD��~��|R��	�n��zh"7A�Aj ��Dܟ�	���	ߟ�Suyblv�(I�v��O<8�v�Y�]i̝
��\�Y�3C�OV�n�y��a��Iោ�	Ɵ�j��@�" Y2
KH@�D�O E�J�mZ`~Bh�>���'��ֿC����L�+p�	Z�I(��<!��?���?����?щ��
ܟM�f��Կ�E�N� L3� �럌�I��iݴ��ͧ�?��i@�'Z%���*��T�'�Ŕa#�ͰՑ|"�'c�O�@�/�MK�O<�J���6a�*�	���-3|~0� ��2s�h3�'��'s���h�	ߟX�I���j�ƴI���PӯO6.% ��I��'��6M^.j�"��Ov�D�|��a��_l��V���V�6���ECR~2�>����?�M>�O����a��>��MQ(7�� C�N)�\	�#A #s��i>McU�'��y'�����X�!ؕXC�*.��d��K�ğ���ş����b>y�'V7�r�RT;Պ�<n$u)�#X�?���
G��<���i��O>u�'<bK�."�T���'N�M�d�P�:v�'���13�i�i�=ʦ���?e��^�� ���ʃ��u��MC�b���zC5O6ʓ�?)���?���?�����]�@������'�Щ���W2>e�m��Ti���'������'Ԗ7=�������K��A@��N(�Z�A��O���8��iT�z�7�j��s��A?"��K�SM|J ��-z� �#L:Dt�$0��<���?1Cb$�8��H(B��8H"K��?���?����d�Ԧ�kf��4��ڟز5M�.X����FP�{)�u�m��zy��Ο��Id�n�VY��D�m̺��W�ѡn��4��u9"��9TȀ�|j2)�O܀��_�N9���s��,ї��3(W�A3���?���?A��h�r�$�e� x�-�66܅yU��,���Φ��r������I��M���w R�cBFJ<
:<��ϿS@-8�'��'B��	�E�Ɲ�����P�iF�D�j��r���a6��$ �1{���O�ʓ�?9��?Q��?I�l��D8(�*9����҂�%V4�2/O��n�3\��=�	��(�	\���D�q���P%�Z#O�4O�aCu-H����O��D;���M�|l���7�y���Z	O� ���Ҁz+�M8,O8�S��X��?�7�9���<i�$�����l�9��y�b�>�?y���?���?�'���yQ�@_ʟ�P��͆A�������Q��l���{��	ܴ��'��?�-O>��Q�Z�X|��9t*H�y3<�ȗ�!'�7�=?���Y�
�h����'���c�KF*i+��:���H��Y�<i���?A���?Q���?�����(�\���%s�B� ��^�P�2�'��(b��+:�����!&�HY�hռ<�|ѳu-߷p�8d�2h�V���d�i>-��i���'S�Z�#[ x�2��c�{��-
 �E72�	���䓙�4�x��O��dμ,
.Q悈9�$������b�$�O ʓ~����\��r�'�\>Ȇ,��@�fyY$b$kH���??��X���	��%��' >mQ�E�<��,�!Wu8�[ "�$�D�k�4��4����'"�'o�� �M(��<�2,Ƌ;��E�F�'�r�'����O�剗�M���*1��D�3R���`��>u4�+O��l�]�3�I��ĸ�.Ϝ=�mۃ�se�cU���ɒK��m�d~Rg�5A��4��[�	�.�L0�/E�X����n+��<A��?���?����?�,�h�I���> ��
��3f�V(��@Ӧ�@������	ȟ�$?����M�;B�v�Q��=(�H����*gG#��?�J>�|�A�+�M��'�����)���;�N6R�R�'_�9���y?�O>q,O�	�O�e0���j��^���S!�O|���O��D�<y��iX��'�B�'��Ї%X�>;>��VD]�Q�����D�]}��'�r�|"�v���z�i�y�3#�Y����Ә2�(�C�Գ[�4��, ���^���$#,Dɐ!.��AGKN �d�O����O��&ڧ�?�EEݼ[�p�	���?E � ��ô�?94�i�\X{"�'ج6�0�i޵!�ʈ&h� �
�d�4r�xR`y�h��Zy"�X�TU�f��HsA�Њ& ����6�v�F��4��T	v5&�$�'���':��'k��'����_c�,�D�-�B�r�\�H��4*��i�,O���,���O���6!X�p�d����.{Z�tjդ�_}"�'�r�|��ԥ�4 Pr'+ѥuB呅14+P���'?��6l���P%�'���&���'z3F)6~,\��!�'/ ����'�r�'R����]��	۴5�hq[�N
Zd���9��h���G8�$���K��V��`}��'���@;��+ n�;Sΐ��Pc�/�R�ZV���'��J�E��?��r��4�w"@�DE,uo6��� _$A"��'L�'>��'"�'Z���xV�����S��#3U 	����O���O8�nK�6����|�P�~�b�n�"a����"��)��'�"������'ԛ&����Pd�2�c�<��a�̥(��Z�����|W�<�	ߟ��I۟�zd �Cj�R��X2Mh����4��iy"�c�vm���OB�d�O$ʧ/�`�Ӥx��Ya`E�;-v���'����?����S�4f�\������W���1f���vbF��� '��擟�����6�D� !��Y��-ήF�������l���O��d�Ot��<�4�i㼔��#Z;�
5Q�f��'&����9;剂�M+�"f�>y��P��:Aɖ j~�B��8$�|
*O �y�b���� 	Q�F��$�(O���2l��b�j��6�U���#2O�ʓ�?Q��?A��?)�����J�HZn0S�
�������Tn��~@�	���	U�s�p�����s�ې;��@����;yg������5�?����TOO�YK�v4O(�9��� ����9c�x���=O��/���?��>���<���?���F�?�X���&h�5���1�?y��?�����CȦ���LƟd�IƟ�8GF�1w��I!���,[��N��Q	�	ǟ`��E�=r��m�\3�bC�-��6X��	[PE�M~�3'�ODE���K�X}��������!�B�?��'�'���S�x:��>/�|	�#�q\đ��� #ش�bp���?�W�i��O�.C7�i�A&	�����c@O/.m�$�O�D�Onaʑ#k���qyzp��?� �����-��SLߵI��T	��$�d�<)��?���?!��?�0@�;80(���Y�EB�i�ɟ���Qʦ�1Є�˟���ޟ����Ży �X���@���a-_��I���L�)擉\I��ˠ#&�*�b�L� 4�Ȱ�Lꦥ�'�J8�dB?�L>9)O�i�A��8�pS^���D�Ь�?q���?!��?ͧ�����N���`�7Z�>�Z�&��1se�`�'�S��X��4��'>�ꓣ?����?�A�X�9�H�+)C��E�ఖ���M3�OB��cF��(�t��Ԁ�0;�$��^p���m\��OR�D�O��d�OH��4�S1C�-���N�J'��dK�@R� �	ӟ�����M��|B��N����|2l�#Nu�T�SHŅ���sa�-��'�b���tB�<*ƛV�����:D>������fq�!�g�œb&6�K��O��O�˓�?���?a��~g<�AC�ȲU�z"@�Zw�$���?/Om�Q8��������o���ȗ:��ōA&3�`��������C}��'Hr�|ʟ�H��Ř.�z���i�j�9�d��H*��h�(_�LI�i>1���'��&���(ð!�E�3�*
�����T�d��ɟ�	��b>a�'�\����6�RJ5��jU��J��A�Q�'�b�h��8(�O
��3O2��I�V9��Pw��h�&2��?I�Å��M��O�mSO�O�t�&�,T�\�ё��tMH�H�'��	⟼�I���I����IV��'�
L� �鐣ɴC��Q1NB�,N�6-�0*v���O��d.�9OAlz޽�׈Պ^� �-S:46�9���러�I@�)�847p!l��<y7�%�h9����y.AQ�<1���"[����1�䓢�4�����*3����ɝ�.���	X���O���O�˓p����̓���'W�w�$�p�A�hx��I���O�<�'�r�'��'�){�(B�pԊ0D�ˉ@�.��O��I�)��7�!�nP���O`a ��!J�5�FQ�Jx�w��O���O(�d�<E�t�'ᦘ����6��l(��5;o�ar��'f~7MB�D2˓DQ���4�0Š����1�$�!����~YV�QC=O��D�O�ZB�7�5?�U�_z�@?,ڑ,#j�Q��A�f:�X��K �$�<ͧ�?����?����?�����\�Nyc��_������������E�c��vy"�'m�O��i��Um��PP!�!D�0ohj꓊?������Q/o� ��6���}�:p���/�M#�	�!��I�w�Xt�g�'��'�`�'��t���]/j�* ³ ���P8r�'[r�'7����dP��شV�<���lo���VJ�>���`ac�Y0�����Y����d[i}��'���'�f��w%M�Y�(D�A�5ղ�`��&_�6��Pˢ��#Yi��?�	��p��^B�ur��Q%gOp�(0<O����O���O���Of�?1�s*�zo�Y�2�82���{���,�IןX�ڴ-.v1�'�?���i��'b���ڴTCV � e*3� 	�y"�'P�	v,��lb~2&�'AҺ9a��S�8�``�T+�`iP���ҟ40��|�]��������I���0Pcլɢ ��#]� u�u����۟(�Ity��dӎHȢ*�O��D�O,�'qxL}:��;����R�:(�8��'���?����S�d���O��(A��KWo�mr��?����t�7N֛擟�ӦK���-�ԮR3"S�ϒ��b��EQ�'���'����OV�I��M���$/z|�����tA�֍�l% �y#I�<Q4�i��O��'�Rb��h5�����5=V:-�E�V��剠$�llZJ~B�̓.d�H���\L�I�"8�����4���"�T"
����jy��'�B�'�R�'�B\>�H@�e�&X�̺-c*e�⛒�M��ŋ��?A���?�K~R��X���w��f�uT:�r�(k���'&b�|��dc�t�?O�J��)l�ȁ�ՅP��PP6Ol�L^�~��|_�$�	�������N�~<x���j�.���k@ٟl��՟ ��\y��uӌ�jPB�O��$�Of�;e��+ ����Ǜ�gcxJq�&������O��D;��Q�n��|S��!0lz��$�/Ft�	?B0ؼ#�Ŋ�_��c>�+��'��5�I;Vv�Aj �e��t`�I�<��������������Q��y����z���a���0��h���*A#"�y�2�Q��O�������?ͻH���Ŧ�9^�8)9�BR6K%^e͓�?����?��OF��MC�OȨ��M��������U��D�U��.�xb�'E��؟���(���ɯI�����m-T��Y���0�^zy�`}�6�`�<a����'�?��iR�$=�t B�*y�(Q&�9(��������`�)���H)ϐ$"{n(**�@#����@���Y�'? 5@bˋC?�L>�-O�hIq�R�N@u�$��`���M�O��D�Ox���O�)�<i@�i��i�&�'^F��GFE�*��D�q�I�w�Fl؟' P6-5�	����O��D�O��y���_��j�	��e��"��Z��7�9?���V"-���!������do�"ھd�AI�4�ޡq�fa�(�	��IΟ�������"�!mNT�`��vW���@a��?���?�v�i���O��hӸ�O"���2����EDY/5u�y��.#�D�O��4��qEoeӨ��|D� D��c�C+$˾q��Mע.V�A�b.�.�~�|�R���(��Οs�䈖W�y�%��%8زٱ� X��0�Ilyr�h�J�bb�Oh�D�O��'U|v=!��ʒ^�X�t�C�2*Z�'�4꓂?Q���S�DɎc���'�U�.��H# ����0��A)p�X]j�\�據�ҩYa�	/R���f��\Jb!p��>^������	ǟ��)�SQy҈r�Ƭy�/�8&�y�!UYxPsg�*G���d�O�n�B�����Ɵ䙇̔�;F���p+F8�T��S,Xny��?�������
���M�Hyr�T�t�=���O e��J�I���y�X���I�T�I����֟$�O����U,
Z�p��/C"�jU�nӊ�pP�O����OB���D	���CK��`���u$��K�cP�2����ԟ�&�b>s§�ئY��Z$��3��9�%U>(͓D�,��si�O�PZM>�+O��O�����;}�0<�q��^�8D�O��d�OX�$�<��i��0��'Z��'-�݋@"x�}S ^1:^T([���J}B�'b�Oʱ���Y�P�)*���G��Й�$R4	��i9�i)�Ak�h<�����ॡ�;'��#7��X��`�b�ڟ��I�0��ڟ�E���'n�4��ѝ0^�Z���7�%�'Kx7C�ʖ�d�O�mP�ӼC O� �*x������q�͇�<���?���j�n��4���F�t`Bm��'p2��a�,��~�<0ۣ)Q���Ó'?���<�'�?����?Q���?����/ZY�
�	nfJtd����D䦩����p�	Ο�'?y�	�c�ܭ���#@c����.�ʀ(�O��d�Op�O1� ��éOJp�i;�Ȕ>��]RԨ�A�i�Z�t���K�Ƶ��'���'�d\AN�.z��!%�sbvXC6�'�b�'����Z��H�4w��$C��oM���t ��]JL�t�Z�� ���&���A}"�'o��'Ά�G��h����8N��!��yN����rV��6ai�)*�	��Z����Ֆ ,T���~}L)CP9O^���O����O"���OT�?�"2��1!���P/C�'����L����۟t��4>�lϧ�?YP�i�'��9�˫��i(@(��sWj�pV�|B�'��O�M�¸i��	'e�����^ƀ	��)<hp�:(þq���`�	~y�O���'�2���)�ҍ&�̗�t]Jd텅x��'��ɹ�M��o���?���?�.��d��HeY慛��Nd`�r��l�OT��=�)�A��y��!6�8�h#� �L�&nݗJQ )O�8�?1D�-��E�L�T5C�HBm�  [�5(��d�O����O2��<��iL�аu#W�'�	���b4�H�Ci��[5�	��M����>��i����gB(�cOE0:�
Q����?�ӂ�(�M��O��3Bې�I?�Y���L�d0f&R?^
��yD}�8�'���',��'L��'5��_�صrB��F���C�B׺a�E{ܴ
��Y��?9����<��y��G%b�I��ׇ=|���U,ӈ#�R�'ɧ�O�j]���i��bQ,�B������t�r��3/��-<*h���*��Ob�S�jC.in\P�7(��a�&�r����0<��iS���'[��'79�'�#AW�	1��l�25�� V}"�'��|�z'iɃ,�18����2L.��$Y�:�B��	�MS4��d��R?���m��3��:��m�Rh�]�\��w�ma��;e����썅\̸L��8_�f-���!�M��w�pA( ͞9L*�r,@ 	��9!�'P��'����&J�V����	��%���F^�
��h8�B@�s2]��|\�8Dr&�g�!��J+6���nA��dU٦�;��������ڟx�*�/:]�� �G�+8�5���&��	ٟ\�	e�)�ӈZq����
�`�j�R�HP��5�����.O�0`E�K�~�|�U�ĳ��ݏ}.ĸ"�$��,�h)��%�O~�m��p�R��	!8��Y�LkE�x�R�לVǄ�ɂ�M�2f�>����?1��:ʭQ�Z�<o��P���>j~<ە���M+�O��)�l��V+&�I��<�qOL9��C�&C��0�;O�����d�D��7�D>?�%E��6�d�OV��]ަI!�5z��i��'�Q�s%��mOb%zᇎ
����|��'��Ou\��Ʋi��	�`�d��OϸP�l�ڒ�I+�A�r�A�Z���<���<1�B�
�Uu����O�t9DphG�J��OJ�m�a�Tŕ'4�Q>�ñ��9`�Jq�2�)k�	�N1?��U���ޟ�'�������N�<F�^�F�Y�I���PL�8&lUC��:��4�.����ꢓO^�2CJ�����$�+;)<���O<=n�%D��+�׎b�l@ڕBA�v�R��$�����	��M��i�>9����;Ԁ�6��`�>������?1��^�MS�O5 ����U����i;/Z.-�kɾ\��Ӈ+k���'��{�C��c R��f�w���Q��)|�6^�4�����Or��'�S7�Mϻ@Бa'"�% ���ZPbN;������?J>�|J����M뛧� H�@��L�BCV����W�w(�(&>O��*6D(�~ҝ|�[�p����0��.
�r�҅�`��/?�S�#���������	qyb�z�v<��'�<Q��:��$�shW1H�4Ja�6<<=����>���?YM>	u'̗�p����@�� ��Y~"l
;� <�p�i�ғ��EX�'�g$"v�1zN�7uЉ`@�n6��'w��'���Sݟ�P����w��e ���]�"LV̟��޴��0���?���i#�O������[�(�:_�V%����d�O��$�O6�Bd�x�~�T	��Qi�?��JĢ_�,�ĥM�] YyS��B�	Cy��'��'J��'M�Bʱ}��vhͷ<qΈ�b�]�j剭�M�aM��?��?qL~��e�yʲ(ٺH<���b�ܼ�rV�D����$�b>u��$�j���h �E��D��zP�o����dF "����'0�'r�I�m��p��bC!Z�@<J�n�8�9��ɟ��	�L�i>Q�'��6�Ъy����8
/r�Q�Z�7�P�/ �B�B��ݦi�?�eW���I蟌��b�f%H��S�D��� ���*v��ئ��'�NT:t��?����t�w�4�=WFR��p�V�t"ސ8�'B��'���'%��'h�2�97�J��*|[1n��i+6� ��O���OԸl�9���ן0��4��l�X�{łG!#4��X�L�b��=�N>Y���?�'e[�dk�4�����٣�Fݧ?�"E�jЖ�@'�"m���������O6���O��>��83+�2�����~\�d�O�ʓl6��@b�'^>����FC�Z}`2%]��n�`�u�8������O��)��?]����&���+�zV�����SJ�Z4ī��O��ᗧ��E���J�|b!I�Ga>�9��Y��b0[1d�F��')��'m��^��,�h�!!Ꮔ4�&��"�PT�@D��;W��$�Oȸm�j���`�O�G�k��S�daL���	�q����O��R�ai��w��U��?�'�ƙ�RŞ'a��q�`\�L�P8�'Q�IX�I�|�����M�t�[�h؆�S�w�Ms�u֮7�
��x���O���=���O(�oz޵������E�Qa ��LP��"[��l��D�)��&|â�mZ�<��P$mXi�w�W"�\����<����u�t��������O��d�$�i"%�ў_����Q;%��d�Ox�d�O~�U����ݮ���'R���!0�&�R2W�|�GC�)]�'\�M�>	��?�J>��	8N�6�S��W0�&TJ��t~�ٹ`���g"��!�O����	�!Z��F�qA�x��a�.V7�J��	�
��'Wr�'P��s�}�r�{�e`Qa4f��A�f�ԟ�8޴\�"H"��?1 �i!�'}�w��b˟�|}>���.ۘS�e��'��'���%��&���]�S�y��*!&~����ׁk2�,[0�לz*ԩ��|bX���Iߟ����h��ϟ0��O�\�4��&qT��
&�y��dӔ�����O��D�Ov����$·c.��0J�.�lׁ�1�T�C�Q������%�b>��%���D6�a���{�ɉ�="�nڢ��dN�l��1�'z�'v�IjC�]*�kϳ@�U"�	̣Y�����ݦ�8!�OϟD�U&R%���e��XJ��$�j��A�4��'���?����?��,� ;^<���&��8���P;xD�؛ٴ���n�!���`������J5���bL�f5�a���ޚ<��?�O����E'@����!�8�,� 	�<�> �fC������ަ�%�Ȣ� �B��}HgJ��$�� �Gl�ޟ��i>��a`ۦ��u����@ A&�A��IN���B��,��|�R���?�џr��ih�����4�x�'��6
~����Oj��|�֡E�(��}��J����;S��}~2ǵ>9���?�J>�OR-Cp��(c@<�L=}
Z���!�"nR��p�i���|��J��('��)T��u�T3���/��xRT
O��nڢl�d{է��a-�M t�#0}8mI�&��l���MS���>���
�T�d�۰=�n��Ɗ_�ح����?ٴǒ"�M��O<��4�M���d_�<��&��"�2a4�P��e�	rk�Idy��'��'�R�'�V>�J�]0?	����vE�1"pg���M+�A5�?����?M~��r��w��� ��U���kD�E���'@�O1��H��ff�T��5g�V$XC�>�Vl��N`���	�%v0<��
� }8�E�)^���)���
����&�Q�@ �D�'b��(y�%vPR�䐇<A2	�+���������=/8�)�#Z1O�t�B)�1''�1#`Y���y<�(F��'3�(p���/,��	�f��,.�n�5�9�X�`D�Dq.50�jT�PGґ�C�
����h�5IT��&W�yM�IP�����T�KT�%{C_�>�xX�Bo�+C1�d�� Z�M%�����:s�@5��c-%5ʬh�+��L�����Vf�e#����o��y7�#@����b�ݔ�,6�O��D�z���!w��o^��ͽ��<n���P&�������Pg����O ܸ��)y��9�F����ıi���'��	��l|X������OH�� "R��4�]6�L�)�eT�a�T0$�����`J"'�K����h��g���pD]�1G�Lk��3�M�(O��i&��æ	��Ɵ��I�?k�OkL�)O ��t��0�f$�S��J���'�B-��ub�|2�� 6�0��H�Jʠ� �ߍH�LEa�i&�1�%y�P���O@���&)�'���-tV�,"i�cZu{��V�r�J%Zشr��������O�"/�	6�@��_h(���X�J�7��O��$�O�PA�[x}W���	?Y,	91�N���F�s����#d�q$�ȳ�J�<��'�?���?AB�NX�F<��h�(�����$F����'8%�	�>�(O�d7��ƺ|�p��7$�Jȑ$��,/`�	�[���Ծ8�O\���OX��<qd@#W�l MFAt��J�12�\�l�'�R�|��'�r�J�Ph���T�RJ�@��G�@�%�G�'
��ӟ��Iɟ,�'�6�
T p>�Q�L� �Qs�*\��H[��qӖ˓�?IO>I��?	BPt}"�

ɴH!E�Z�@څ������D�O��d�O��a��Tk�S?9��

'8�hp��w�V0�@�ڹ|̖�Z۴�?O>���?�����'-R�*��IsF�PP#_�y��=rߴ�?������ſS����O!�'?�4���Q�X5�D�S:�]ʠ�2BOv�d�Oly���:�IPr6��>�0��6�Q�<ڶ�#����'-����j�@�d�O2�����ק5���#A*��b�`��&�i�F��Ms��?�®<��'q���c"b�7Q9� d�	f�Ř��i���	&Lj�r���O����TD%���(t��m i�&��E8��y������M�)��?�W�Q&�ӡ���W�A�����';��'�����4�4�\�������ƩZ� ��MM%9��,���rӈ�d+��e��Od������Gf+�xx�����. ��ye�q����ޚY6�~���m��2�! ����}�"ɱ@㍧EK�����x�n���$�Of��O�8#4ș�E��w����
56�U�5�Ϝ=^�'k"�'x�'j�i�U��԰3�
{�^ x�>l��{�F�$3�D�O"��?Q�D����t�(�V �T��)vb�X
 H���Ms��?1���'��Ix�7M޹P�����'�a�YY2�
J?��ܟ4�IޟT�'�DpҢ�/�iT�_}��j��S" @0��7p�Z�l�p&�����t�'�'=°��e�ԣ��P�`E�.�Pl��D�'*"`Ȉa��Sߟ����?�X�G�%8E�K�M���`�R']�.O@��<��V��u7���	(sL�e��������d�O�p�u��O����O��,�ӺK��o����KG+=O�T���ݦ��	Sy�I���O�OA̜	A.�F��颴��-���:شvz�8��?����?9�'��?�	�LC1`^L��A�-Hp�4�w�ϛ���J�w��b>��� `Ή�rG�&'��s���F�1��4�?���?�w��#׉��$�''���,.f2t֝6�rxb�l��~���'B�'�\�g~B�'��$�!I��[�,S�qvm+AlE�<��F�'#4c$R�������L��I��~u"��#�z�إ�A��ēL���<	�����O �S��iZ�AZ�j�(>��=�2�	?T�ʓ�?����'���O�(���7"��;�Ęm�*b�i�I��O��d�O���<Y�!R���ӊ,��:�iٔJ��Y��G	W��IٟT��u�	Yy�O�B�ݱ0�d�	M�0P|d� HN0[���?���?�*O�� WOⓌ"5j�Sc��N͚�a�=.�����4�?YM>+O�i�O��O�Z@�$g�&�� !���2>�Z�4�?�.OV�De,"�'�?�����N0�b��j�Z�1���=l�̐%���I_yҀˬ�O��9f������D����;hG��\�LSuDԵ�M�tT?���?�P�O��ʢ�U18ǌ��.ŵfJ-�M�*Ot�d�O@$>�&?7m�i� �'ة��<bR�R�k+�6b�� X�6��O����O&�	V\�i>MoڣT�F���#Y��X1���h���'���'1ɧ���h���цE�$`�L˺W3����
^.�M��?!��D���-O�Z���An�����t�z�C�>�f�Gx��(���O>���OE@%�ڞi�(ٱ��(�1:�
Ц]�	ߖ���O�ʓ�?q)O�����h�fN5I�B�z�ύ�Iv��+�i�B��y��'D2�'$��'�剔kG�U���mxx�Q�)Q�	�5��Y����<a����OH���O�͑�,$k�EC�/�<Y��#g��,e�	���	ޟ8�	y�d��k޾�S�p�@�SPmʵXGHP�Gϗ�|8�6��<1�����O����O(T(�>O���5F�q����@ʻ#���� � զ���П|�	Ο�'��H���~r����h��!ʍ0�(p�"��	��K��M�����O`��O�ԣ2O��D�O�(I_����
>�r( �)ǖ��7-�ON�D�<���Ԥ[Y����d�	�?=�Ł>|C��]7g�M���8����O��D�O�)�6O��O��S�B`�A:%��}>4 cf��47-�<ar�P�a����'j2�'d��c�>�;*Ϧ;b�Q&4�\�]�@�4,n���8���Y��	F�	]ܧ%�L�M�:= ��SOL���4}�zD���i���'"�O.����d�4-P�x��iC4\�ܰ���:�l��l���Yy��'e���k��3�@ ��tsU�N@���o�<��Пp�#����<����~b�=5�x�h&F5YB�-c1.��M�O>�g��<�O���'*Z� b�h5�U aT�8HwQM�aQ��i��������d�Oʓ�?�� @܁RFB��S�� ��#���*P�'�ᣞ'j����L��۟��'f"���
� �BI�f�2��X(�]
qG������O�ʓ�?���?	�#����}����"m����C�4�N���?���?A��?�(O:���(P�|b���+NP��a�9j @�IUƦ��'�2P���I�0���6���CL�))�g������
L3m��@�O���O��$�<�u�S7&��S֟,)G呲f��2�'�S�2�"�c߱�M[�����O��D�O"��4On�'2 ra�I"q}��Rg!�(SG�,)޴�?����D�д�O�2�'��E�Yﮁ����4� ��W'���?����?Ajc~�]���'H&��������=+�!ݚ5��Xlby��(�6��O ���O�	�Z}Zw�&b<��B�)̦e�l���B֊�M;���?�f
�<I����3��=�R`D�Ȼ`�r�Є凥@�H6 o�(m��@��ퟠ�;���<I�"BM0�
�dƻ:��H��Vw���h�����<���t�'�4�`�M0�� {`/3;�����sӒ�$�O��D	�|�0}�'���ʟ,�c��'AI<'�N!
Fj]�r�o�۟ �'��K�����O��$�O��Kv`��[����pc%��P������	lL[�O8˓�?.O:��Ƥy�E%��z�hY�����z�A�A\����Ee����Ο(������y���"0���BҢ(�|�sf��4VC�0
��>9,OD��<1���?�i��e ���RP���S!+�J��a���<���?a���?�����1�ͧLYP%�=3�L����<�>�l�hy��'���d�Iϟ��Ʊ~F��"L�h���C�'r@"�s��@æ��Iß��I��'��e�!��~j���7*ɜ)X����ۼY�A�W�릡��Oyr�'|��'>>��O��I�3���1'�-h���*Ǩ�"@7M�O��$�<)�͜��O���O��in�0=ѸA#t&�9t�.l�E�0���O���ٝ
����:���?���k�-7hp��9(�ݚ��l�~�=� ���i���'�?����I=P�68C��
*�94��yY5�i���'��r�'��'�q�$I���I�R X��"I6b�v�Bb�iN� �aӊ���O����-$�$�ɅM<P�����XP�d�#R�7��"ڴw��9������Ox2
ݝY�<XRhV�L��r��ئ���ǟ��ɮ+L� K<���?��'7��ЁP�/�f#�K�UT-�ڴ��g��|�S�$�'���'y� �Ǣ�DiٳCO ?j�� G|��Dӷz���>�����S7�,��lڷ!Α��L���v}be�y�V����Пx%?��ӭC;v.J��6�$3f�ԉ9�8���}b�'��'�r�':Zt�.ц ��!����Y������?��]�|�	ҟT��wy�(T�`��S�d��f��X���ø�,��P���	�t&���I��z-r��S��H�>��X� *�m�px�����Oj�$�O��Cj�A������O�={ڨx�$_D@ఊ��1?I�7M�O��O��d�Or��T?O�'�ШB����#�����'ܮl�ڴ�?Y���Q	bi�,'>e�I�?�B6Ӆ\b�|!���cΔ�����ē�?!��j�< �������K��dbe�
�]ZBiP���Mk+O&Ż �Y򦝡��0�d��l(�'r:�+�eѨu׎��R�nC��x�4�?���	,�?�I>��t��8�j��r.ԋr��iF�
��M��-}X�F�'h��'[�$`+���8Dt�2��ф41�5ka��3I,%`�4zg�Dϓ����O b�\�"�:庲�S�+o\	��dR���7-�Oʓj(���/O��?	�'r�����0[���蝫7�U��(��OF��'���n��hPS�+[$IQ@��:`�"7M�O�1�eeRd}"/�~���?�K�X V@Ǝ��	�jQ��X�1�d4���Ov�D�O���O�%��X�xU��F��1�Qg�4�>��?A��?yH>I���~�J�?V�F�ps�C��u�t�M0%	W~��'C�R���I1�"9��Z|ڨ0�m�o�p��ӆA��P�n�ٟ��I֟p$���	Vyr���M[��4Rt�q���z� A8� �|}b�'\��'�剢'ґ�H|
BB#d� pA�2!��C�!B�s�'>�'���Iof�<I#O�~��KO�z��7-�O���<�a��7Gm�O�2�Ovܔ��цg�![%��=�,Q���9�d�O��Ƅr����K�(٦�\�K. ���R�V8��m�SyR��WZ�6��O����O��ITZ}Zw���:�&˂E�2��!k�u��@ڴ�?Q�R�h�͓KB�s���}��C<j�F����S)�6���
Ӧ�aV\��M���?�����[�l�'#�����x�Zͳ�!.)��l�G�e����O��?y�I1p��y+B�H7j`h9��	i�r�!ܴ�?����?q���B��Iwy��'��՝*�.8�d�X�tt|i��ǣ>t�6�'���(x���)����?��*�Fm�Q�� ,��Sv�S���c�i0���7~2����$�OBʓ�?�10��xiFFQpӼey�b��;�Ɖl���Ky���'U�'�2R��#E��t�:p'ˊ8Pi8B흩�	S�O�˓�?�.O��d�O���A�d��|C$�8bU4�Z�m *8�8OF�d�O�d�O�D�<�գ[�>�� 
$*sb��s����c˫M�.�pS�im�	ܟ �'lb�'q"��*�y��ěs&8�PTm6	��Y����,��7��O����O�d�<�"�K�p����֘)B?����[�S0�����.��7��O^��?A���?�se��<�-Or�P�D\�xI�X0e�H�C�d���9�	ş�'I�Q"h�~z���?	�'<�>,��c�CX�Cpx��[���Iߟ��I-���	ȟ��	՟���A��b@h�uc�(@EJ"
ynZ^y�n��Rm6M�O��D�O��C}Zw������N��(i�R�h�Pܴ�?������?��?I���(ܭr�z!�^
tI�p�@�?ٔ���0g��
A����cH O1D��0�0D���r)?79�!@��)\��,Q���/�j��Sb�@d̢�,�^�)R�+5#�����'@ښ�!��%�:�V B�9��Z��#�@|
@@;b
�x#H�o��i����0|a��"G�-�Lp����-�0�J�B1v9Z@ �	�U����I.%ư0�2DT2_��e�D&�ܟ��ϟd�I��u'�'��5��K�EU���q{��	1͘M+R���83���1��S^�X0jմ<�AG~R�A��]�p+ڀI�`�˖FЍN���� ��=?��-�G�[�[IG�ę9� #=I7�޵1-j�z"ӵR���3(T*�b���⟘G{R���BA�����]�)\	(!�M���6�&"W���z�1OI�'��! G ��O@�$���.�蕞x%^%����%}
���O~�JP��OX��m>Mh�Ϛ�3���s�Y��~��?��� v�A�w���p �p<)��+1^`0�(�sy��L�]}��z�M�	����
�H.�x�Q��?I����	��t�JY�I�x�BQ���k�1Ot����6�V�ؒBݪ'R��J�Ka�!�D�I�s`P�g@&h��+	;f����|�@�'ӈ�� ί>����iH�f�����!�b@��%#�]P�b�6�j�$�O��r�B�%a"ʥ�~���|�-�D!.�LI���D>����>'�Kv*I( ���|���ɖ0:,δH�Ο*��tI&YP�<V �	ܟF�T�'}������zQtq��&� L`P@�	�'�Z`W�1iD��rV���	�ґ��;ҍ٧z��Y�G��f� 8���A.�M���?����Xe�3�?���?a�Ӽ;4�]!sAq� (T/H�r����Tm�%+�MF�p��/�1y4˲cҋbS��:��ϯ>����'�t�BvB�g�ɣ|�R虵 �3Iy��y�o��E�D��|~� ߌ�?�}�Iϟ �ɐ����fG�!M�L@$�8."M%� ��I�}/�uԂE�@�hٰ�fq3 �~���'ɧ�i�<�f
� GH�'�Z�޴�&L�"�J��Q�[��?����?���|
���?	�O���eg�0M�r g��%t�1���cv�7�'Q���䣐�0 �b�%<,�Pf�	rJJ1���'HH1	�_+Z�\EY��؊ D��5����?����?���D�O��X҃o�Gj�IP�c�f�)4g%D�LkF +�"�Y`/W�JJ	�!.�5�M;���������a�q�� �>�{���\!��?y-b�!g�:p��k6'A�!�$�@lHC���!0��I��S�T�!�$����� ㊰i�H��U	!�8-��@qN�-`j�:�M]�^�!��2H�fH��m ���&L4?!��Y�:�3��.U�,z�"��mT!��և��D�U;
qP"t��M�!�d�a"�r 2=�4ѫD1�!�D3Z�ȇ�N����7D��%�!���&$C��9&�P�tNP�CD
NG!��RO���p*��Ts�pW�A�`4!��9f갥�a!�)w�N 	�!ʏ+(!�䎂Xh��hp��P�/3y!�D�SK^��uƞ*&�2s��	,x!��a�L�t�P�l��ゟ��!��é6���4S�4���ǝ�$�!�Ę�[�8�R�A�L�\�� �A��!򤎷`n*T�& �Yk2!R�aԁ|�!�F+|M�d��:w^ P����%�!�$�;�d[b#N#2L*��*9l�!��D�uBr�q�	�#ScD�L�!򄅠M����G�U�N��	��M�!�ZnFT� &�hQ��!R�!�� �M2�K�Pk��i�o�c�^��C"O�t���ޢ�f0�g[�V���I�"O��: MZ�
�q�C�Bu�IB�"OR�6����Z�R�F$,V��d"O�d!��*ME
�J�7eENX�""O�+�ڧ'�]�%	�):l���"O�����0$���(7�̿�t�"O�ّ��ܰ�Y�" �P��چ"O.��4���ѭ�'A�  ��v�<a�CV?U��ZS+�Z��6�g�<�d[$p�tA�
��G$���	c�<��C���@}����3��93$Mu�<)3f�S���"� 	$r���%[r�<b���(�
A�ƀ�b3b!�tnk�<Q���:,�M��慔;Ŏ�Y��i�<�Ɋ.��kq��|&c��Wz�<��	-s��s�ÊR���q�s�<y���}�vf�1#�^�jbH�c�<��d1B�x��$ޫVQ���'�i�<i%�ۑ �걨d�N'���c�MZK�<A1��2W��h�U)L<]�����K�Q�<A�ܑW%��f��F	0�FS��yR��+=M�A�W�_8�|�ħ��y�HY�v�H���اb�j5yt�ٍ�y��)"��yw-NR�NL�ҥ�y�ƞ'1	�I�9*���+�y�KʅH��̑�%'B�"��O��yM�{�Ptkt!ЩHN@�5@+�y�e\��Mڵ�F��3�'P�y
T; �p�� �ǳrW�q��2�y"H� 330u�D�S;d����E��y�A2FҺ	rK�%WRЌ�e���y"��#j��l��IKo�`bi���y�I�4a����Ɯ��-�&EӢ�y�6,� ��f�`d	ֆ_��y"R�q�@f���尕(�	�y�-�%��1J���s�`��ȓh�xe�N�g�j�ضk];rЅ���$��N��ղ#f͑x����R-�F�B%�䙓t��<�� ��h�E�1
�b���:��5�ȓU4L��bƝJg*��@Ɋ-�P���0���i���F�����M�9F�Їȓ{ ����I�j֐����V�`��nD,)#hF51((�2��ʁ"^Q��h�p<�c`ʲp���14jT�kZ���c��Qg�҃)�r}1�׼5��ȓ����Ҍ`|�D)�e0���ȓ\lX�s�m�Y�P�д���t��?a�㓬��?M��i�N���q,�2�Z�
�#D���So�J�n��S!ٻ@�$=)"��8�ư�ܴVr:;�O��g�'K�ܙ��$�t50䮛�Aɢ ��`Y ��V#fD��E��=�$��PD�6����I�KW�����'tJ�q���S���A;3}�=�M�<0��
�z�x�WUF � uB�Cv0�"禮|�BA�'�e!�%�6])D� #.Pj�<��J
̠ !��_�y��JSI\�h�"�(V�����m���B�t	p���'0����Owk�0X@�;���^ۨi��MΨ�xrg� <tQ�Tf"P\@��s��9�V `��	�.��A�	,Y���d`}�	J�p�z���|�$��g@uc 㐔g_N�9�B'�0<9�1|O4�t��t���(�E�)N��P�RgMGRhEC���4Ӓ � g�>��+0?��9O��'Q�[r��BO�MT��C���z5�<u��	E�_t���+A��r�������h֚9'0;Q���j�h�WA:(,��3�B��xb��9X��8�ذm�����	�T�����º���2��T�c��;P��xgٲiC(�ԧ�[Wř�'<9qIR�_a����U<YQɁw�? �<:�-�f�adf�;5�6��Ց)���Fe�/"�V��`!���6.�n115�:��$=��`��MԬ*�>�	B.��(�ax��b�T��W 9�Er������P@f�ԥ1jrk �hz"�x�ey���<9Ó.�t��F��}�x�t�Y�|���'�z���R9�MHщ��a�	�R��8O��T����p��s����G��#�"O��7�M�O�|�1B�ǳD�m2�G֛�Z����G;c��<J6��6��O�=H2��V}R��m\�ٹ��Q0;F�)���?�$���G�e����jA
��MA�>��I"CTi�����0XuY��_�d�DdG~r�)Ҹ"Pc�xx�u�	�Q���&�Y*7�ꍲ��bn��U�뛴`��\���T'p�aY1�uN��
���%|�a�U�В�.�0!DE�3�G���Dފmք~5bD�`�W�a4d��"Da�o���M�{Y2�)vЄ&�C�	�`̀�)�$�r#���E�/*~l��ؾr�2"3�i����Gɗ]��:Z}���+OBA�d��~:8�1U�6vs>�2
O��	��@�5��#%U>�B���(���T���<PV�z��Ó3�����Y�{ڦ$��v���I�;Z�,��6��9�:�AXFoP/���`*R<�'g!�43c��|z�1:0&؎eL8	w'-�	3���K�Ĝ�SL��c���xܧH[Ε:ġ�(>�,5A�	V�t���ȓi��);V)�M�����Q�>Fd��2���#¡�d,>��D4�g?qQeB�Dq�4H2��O٢	)��N�<)��0���k�W[�U�Q��<�e��0ax�I���<9�A)=c�߿�rXQaK�gX�䲦ʆ<�:i�a���Ip��Kq*@�-Q��y��ހ��%y@g]9EP��aR&�"O���J$�'���;��H��� �PhC�v�p��
����K8p�YrFn̶V%��ȓaF�Xc��U0 �$<���/O���ȓ'�L����;C"���
ѵ�(Q��!�Np#r�D�\Aޜ�6MV�=��ȓ~8�pa4�ʺ+�&X�E�ŉlhL��H��y�Z�(�D�Ӡ�P�Z��E�~����?e `����b��]�ȓ/��1�´M���b�%�
D���|�M���'��ݐQ�V[
�ʤlW%�fu����y`�8�y�%�,H���lÉE�(�6�م�y�
ϤI%^���h_�7a̪�"��(O�P�A
Φ͈�$dX��Ɠ[�98t%Q�J���"O��$fߟ'mp���nY�N컇nX(Dj��9R���O��
b+�(rN����'Q2'�>x��"O(H{tiN<1���%`��@lZdR��᭏,�0>Ѡf�%�,)�em�= �`��$�G�<� �f��x3� �5�ّ��@�<���̟N��8�%�zi�Ap)�B�<����:;Knh��A�4G|�P�$�B�<��a��3��H2e*J� �#4b�@�<�@� ~8���2l��UR`�o	W�<���
%�d�t�� ���NT�<Y���;9&�|+Ď% i� ����M�<�`I�j)�I2qH�*�Z�Q) H�<�t(��!Ą�,b��L��G�<�I[�n��Pr� u5^��VC�~�<��!� �j��t��I/����b�<	���).�8��$Yp�Bԛ���[�<�v.N)cT�u#X]�FT;���S�<q��%�p�*O4.U�IӁ��f�<�����FM�% �~�� C5([^�<���Y����d5:� ���S�<yҩ�3��q��ذ,�`bg�Z�<�ƃ&|��&IvF�`�O�V�<aƭ��.�&XXt��S�H}J��X�<y�-�9c4��!"��=TV.�8#J�<���]�d$Yq�OO�g��M���DC�<u�0%�֡���zR��I����<� N���I,��z�E��b �2�"O��4eHs��`��%C�	y�"OT���(��ɱ�/׈ā9k�"O� ˀ'x� ��͕*�˵"OhȈ&�͑ \��P��9"OXMz�NX5
���Y�� )�b�x�"O}�&�/C-�I@k�%�|y�4"OvZ���lH�́S�C@���+�"O6�x �E&Xl�0�4H�<��]k�"O&ESF���Ib��g	�qFh�{!"On�1�F�$�\�Ȑ�ú:=���v"OԤCH
�Jv�T#%�9q"O�T	��(��	��'O�i��iqf"OB�ԽL�N�:���"�"B"Ol�%,��Nd���jA%}��"O��]2��1�A:���#�σ�y"-�3�*�I�ɕ1/�(Đd���y�ġ��JW/�qB�M�cA?�y���"Fx-kF�X� ,�g�4�y"bZ�T��#e���C`l�J��ǒ�y��ϴC�nwA�6S����G�
�yrO��8.2�C.KL���v���y�,N6,t�y�2i5o����'��'�y���-�0Z,��g	�˓��y�k�a�Q�&�N�w&�UV��]�ȓe7,��SQE�;��'s��?�*�Q�/�& +&�Z`K�H���ȓL�x�q��Ăx�!�2N�<]�ȓ�����B�H�ł4�ٮ��L��D�I���XA:�r�2^8a��-�Z����6jj�Z�) ,x��\�ȓ/�u�b��CI��l��[7��2t�eJw��f�~I[� �1�n]��Z�4]؆�ʓl/�Bv$_�#ŀ4�ȓ���"P4�آ��̗E���ȓTz$�1�"�"v(�Z��:=&ĄȓI�����ڧe�}:T�T$��I��V- A�˔;hI����F��\Q�M�ȓL����Zu�\R�!Ĵ)�d��ȓ.����1f�'0�j�h�&_��2`�ȓ^b��0���,��jѬK����/ �(���H�
�b���)Ѭt�Їȓr��	D匳i�h�h��\�V�X��HT�0��
m�Af \|�E��'�(����[9(MX�h�$0�
�ȓ  ��¢��6�|���Z�T��Ɇ�=0�Xe0T�z�*��ŔwHNԆ�,��3)V���	�$�Z
%d��� �p������nivp�,�%¤��	�t�0�jN��9�tC۠��H��A�	1"�,�@L3@I�e�d�ȓ:��[РH8v� �֯��	����k񎭻á kb��!@�D�Td1�ȓL�R͘D��1
�i�`��W����M�~(�	��BD�
EoV�)*���2�&,�l\V���n��4��dq��� Ied8�7�G�-2X)��i�D�r�bX�F]���`ߜE���Bc�E������>%�C��3��`��!�6љ��2R��8 �X�p�؍��=�$,BEȆ�[1�4�'*^�9�ʥ�ȓ%+&<��Ş3Ԑ�H1'�*n8<̇ȓ4	@A�UA�%^*tA`�n�* b�|��n�.�I013��3�!$-�\��S�? ��Z��_-�Ұ��ΐ#R��ݣ�"Od�{�CT�/d��2���'r�8��"O~)i���>-mE���%W�!�""O��k��L��!ȧ'�`=��pq"O�`�%�G��"̲T��%{��!�"O�0�pM0�2Y� mz�p�%"Of%@a�A�r+�ÑnrF1#�"OԍW��-|�� (��&n|ꩣ�"Ov|R�V�?�5�ś6Fn��q�"Of (w�٤m��C��<iF�W"Oj��`�q�ѡ"�T �@"Of�+SoF j��T!���<%[�"O��
��0z	�k��+32	��"O���4M��d�	�4u��t"O��
7M̿��He�'�@�"O,ň dU��XU��q��%��"O�����*{It��)����B7"O��We҉!�||[�H\	f��p�"O��p�#ߛ:���I曇�Rex�"O�d� UǊ=�&��p�Q`"O� ҧ�n�$TZ�W,,�]��"OL}��琉!���`*F8ڢ$3�"O�́��أo�E�p	X�N*��Ct"O��P�,�|��'D�>�`!"Ol!j��T�I%(��M�X��P�"O�`�ǆ*���B�T�u�kF"Oƽ�R��\i�QX��Ai�}�P"O�a�Ꮭ�bF�kh��aM��s�"OvDaG���2��Я�++����
`�<9���/��|#�/N1M� I �F�<7%'R�Z"E2[�h�Gc
F�<�§LA ���e�`~(B�@�<��-M�@DT0R��F,mH	
�f�x�<��E�1B0�e��Ą�v ���Z�<��`�46�,��U��1����7�N@�<i�*G=iNv=���U-H� ���f�<��%Y;=��!u���~ ##f^�<Y�jԒ.�@(�R��]��u[���\�<�G�ƃIy��� �� ORm�Ҥ�X�<92a\�%����r㞞�M��B���yR�P:���gF�.����HH��y�I��]�ՋY6"�$�Q���y����nT!�B����8� �fG��y"lY�eJ��c�����eHA��y�]���m�z�D�s�� �y2��68WJ�gOӀt�t������y�'�e`��� �W�d�FAY� Ӟ�y��
4mǲH� �۠����y"@Ň_���Tkβ�LiZ�C!�ybB�-�E��b�n��,�=�y��	�F�ZP���	�il��z����y�C�ii�Dx�OZv|�����y��ݍ}�|ZR���Q�D�yb��	)��`R
J[Q�-SC���y-�*<V�+�-�OՖ���L��y�b�4]{$,Y;s��,�ĪQ(�y"
 *����0dz�\�%I���y��,��(��j�(@,����ܛ�yM�3����F̾C(�f���y��T�c<Pr6k��eJշ�y""��u@L Ȅ��#���҃l���y2�R�.#F�Y���,6p9#����yRe�2<P��-��:84X8nT��y�oc���0�ݱ*5&R`�	���p>�  ��Ơ�(����Fݵ�m�"O����ݶ>!`��c�K
~
<��T"O�ahP�_I�� +�
�Z%��"OBE�t'��U�ء�OM�
�<H3�"O��B�ٌw�,в���	10h��i)���Z�9q>��@�}c�ူBV! �!��nW"�Ԯ��4U���䡊��!��R�Y��mz�Z@T�]���a!�D�)ô�@�f�18I,d�с�+p!��+�إ��a9�Pp��7DT!�D;P�0�A�_�^t�`��5:!�$��~���ZU�܄��A�یY!���*�
��E	�9�tt�%��o|!��Śc>�I�4��h��S2�=a_!�dO%�daE�)����c�7[!����Xe��&C�vt�a�\�1�!�dW�<UD\����EYʸБLW�]o!��:>m0�a�*�aM�1EL �f!�H�G.�+Ѝ,X~�QFŒ�:_!�$�2�m!� �".��QJ7!�!��'J�h�c0����XB��RA�!��oTę����&Vhͪ�Ə4e�!�d��0!�w �^��˷��!� �������L�V�%hϽk�!�O�xA�ݛU�^t~رs7��*�!�d�R��q��S=my�c�(�5E!��Âkb���g9N
�� �g}!��E8��	�ib ���u�!�d�TH!����)Abĝ+"�Ă�!�d_�5Y(�Y���DxT�x�݀,w!��S�@#��x��܉f�iP�-92�!�$��_����@eN�%���S�!򤚈�8M�W�=5Yr�#�0�!�䕧z��-���I {10}�#B��!�d	*`�*�ڱ�ȑ��*��ۧ^m!�$��2v%2�V,�l�QP�C8V�!�O>I�t|I.\�h¶NƼ�!�d���]:��D��6.F�:0m�[�<aנ�3^ؑ��m��^sX8iB�O�<����,���������I�T��I�<ߡ5<�����4S�����E�<�t�Ǽ#8D3��U�d��8�L�}�<)�L��:��1/�z�|��WI�x�<��S7	6�K1-FV����v�<�#�6Ux�"���9���Yg��B�	2(�Y 0l��EL����* �g�LB�I��[r)�^��zV%�w%B��)I�x�kA"�s��W�<0B䉇8հ|0w��9y���s�ȬB8�B�� u��qЯ�(z/� �'� {�B�I�{���ʔc���Q�A|9�C�I9fҀdBV���b(���
RB�v\�d��L�-1�!��/�)$]&B�I3R*�j�n�-(����sD�,V"<iϓ:�P�+�N������^�C��i��g�㤉V�Qt�P��gZ� 2>��ȓpU@@o�9�(���ړl?6܇ȓma���	�M��IZ;Ygt��C���	UӾ�b�0�A��kXX�ȓZr�)��kN�oRp���e�/ �*e��	k�'���a���:|��]���k�d��"Ol�����H��0�ʵi��Xxr"Odݚ�a�g�)r5dR<P�d�"O4 )��X{v���E�|с2"O� �M֋�?0@�9��Ц=�|�jC"Oh-ٶ�B�aFa�ᅼP�����"OH�ɕB��y/���f!�szP\�"O
���N�S3N�9AϯA!1"Oxa�f�y�ܔIt ��O�=��"O�{��� H��A��:%vej"O�Q�r���
���9Gϑ.r����"O�1S�	�+��;��XK���J�"O�p��G�]z,)���l�R���"O���Z >�ب�D C;M;=��"OBQ�S�߃~e� <*���"Ot�*�%I0:V<)�QČ(l��t"O<�; ]*E�AQCc�b�d� �"O�����^�~|b�@����`�4"Ob����7��m�'�v��Y �"O.yE��S�8��w��K��9C'"O�@"��ַ�ң"�-Y��4 �"OF8��-G�x�0M�p���1�ʍ`�"ON�Y2�ӿ:7�LzFb�n�6L{�"OR%����&v�xDcLQ#tJ���"O0<J��8Z��=Y���@h����"O�ɋ���.~����*��#nڬ�"O�M:�Q&yt��"'��Q 8 �"O�kSk�z�Z2-VcZ��#"O��2.H5.t��E�8I���q"OD�D%�e�D�aR���b<K4"Ot�"�� Vh9k$䅡v�ٚQ"O��c�T"M�4hu�����l3"ODj��S�*�X1�⓾5���V"O8��D�B�h���`}�.���"O8h�F�Ʃ5��AM��5@({'"Ol��G/�0N�T���N�E �40w"O��Q��w.��酨
�٨�"O�q��mR;J�8����4o�Ls"O D��QE��i�kP�[�m��"O��#�!����)I�O0X�ش"O�6#^���ޚ<NEҤÍ�3!�ĕ�@^��)G#�,,�	����'���aD'B�����	?aZH��'/*�@�l�l3�h��ٱ2g<t��'*�a3�,P$?"T�Ud�?10����'� �K�`Pþ<�QK�t���J�'�Ta30g��^3:���a���i�'������8�-��L:1%@�I	�'�|�c���0~��S�&S.Y0���'*��M��y.��auG�0�A��'�\�ł{ӒĚ5L�=}�c�'�*�I��B�5H&�z�� 4O}��
�'����*�?h&Y�s�Z�@*X�!
�' ։zQ��{�\�zC�ɇ0-���	�'�ᒻ�!��Ĥ(�p,k���yRàf�(|�3��N�SO���y2&�2��5&D�?�K�.���yҢS5v�j�K`n:Rra6 A��y��2��آ#�F��u'̎�yၣ5B{wM�1Q�B�n�6�y"#�s)��r#�D)���TƋ��yrFM�	��M����eɊ�y��"��� �`����yւ	�y�o��a�ð�L8�Τ{D�Q��y���Iup�+�	��6��9�F 	��y�K��	r�y�`(�(r 9�f���y�g��Mm���)תl�"���.�y,Xm!d؀NR$r/������y
� J�8I��Z�xE������k�"O
m"FL$[�L�B�ΉO|�\�!"O�:PDP%��� Ͽ�
���"O�$�%B�A@UC$"y��4"Oգ��E�x�z�{���=Vb,8("Oxt�i��D��Q�k�:|Qv�*�"O��G�e
��Zk��!Jn�Rp"O@��'�\�vyr9����04���"O���QM�$4�Y�&U�1��"O ����Y%BB���� �.$�P�"O���"���
�]" ��y�Zݳ�"O�]+��*��`��W�i����s"O*�k��ۋB�X���甛W�� �"O����Çz^
���E�u�^��"O2� �A�ȒH���8��!��"O<��⋘�a!n,��m�)�l�C"O��ĭB�:��$��b��4i�"O�U�T[]�-�o�-�m��"O���R!K<[x��sg.Q	�<
�"O�$XR�3tvx� 7+�8F�"�0'"O��NgU�����1&�܍h�"O*T{ ✀F-@�d�64@�1�"Ov�k��X��0���8Kf���"O�bjEsBm�%K���p�U"O��V��^�6��%���O�<LZ"O�u C�˞oa��/�,-ovсw"O*)0d"!2~z�#��"Qe�@��"Ob�2��L��D
>Y���E"O^D�Wk_�Z`P�;R%WRVf�H�"O��3c�P㖁��D(|1���"O��0��@�V���bX	:��C&"OVI����u�����!�Aװ�d"O���b�?8��E���Tʹ<��"O�hJ5��5. e�7 E�U���d"O�Dr�K+���-P3i���ӱ"O>	�uĞ(5a�K��s�z%��"O��1\&9�,p9���=o���e"O�4��$.]��U��DP�{���+�"O
q��l��P�ԀK��$OV�M�<i�'צ=t� YF`�X����L�<Ab��30t���-\�+��kp��m�<����J�N� �h�3j�؈��Fh�<)�-�<E-BH����Ch�ɻ��a�<��)�#��u�IZ�3� K#�E�<1D�A�,���4�p��\����<�1�Ӻ9��C�N��h�^��R�x�<Q���r̶Ɋc��vB����Lu�<1�I�u��"ʔ�� �Ik�<�2M�m>�l����,�XgO�<�p'�F�� P�3��Ñ,�K�<�'L�JZ��p�NS�!}B��1GIl�<Y��Y�L}>��a��",�j��!+V�<��_�>&�0�
�%S��kF�[~�<�2���*r�b���mh����I f�<w`�(o��9Rp��'� %��Lv�<I�cȶC��
�&M ���b�ğZ�<��h�92Nu�ፉ6<9�s��V�<q�ǈ�^�!'#D*?����3 �S�<y�b.s\f��`�ӻ#���Hd��L�<Y&H�E��s��9����FJ�<�3d�
%��I.�_���$ I�<��nW���a��T�EB�ı� G�<����0��	��@(c�Kn�}�<��M��Ar�Y�2mM�
|b0:��q�<� �<�1�E�20(p'�@�G[¬��"O����b^n��s��=K��3�"O���aK Q�v�J�b�i%f]�U"O��0���5 �F���Sw�pX�"O@+��Ќ?�$�0���ke��v"O���qm\�C�����/�[a��C�"O�d��Kηf<�bvn�;u<kt"O ����#ea�m	���b��8�S"OȄ��MZ,&X [a�U��A�"O ��� M�s`���	�?�ڍ��"O����
ё;��
�+׋�Z�bC"O��C����B��[�5��ڥ"O���񆘺a$��'�ǘ4�`%�"OЭR�M;�
�ң ��I���"OF@���J3�$�I���(s"O��c��RG ~��R胢� �v"O�X���<u����7��ʜ�� "O���Gە����GVS�H�+%"OB�x׏�5i���D�Q�@��E�$"OL,9�m0$5�a��]rG�)D��S��B1M���F�D)��.%D��H0bX$`i��c�T
��E->D����d��~���F:p��P)�7D����#�/��9��$ܣ��8#�8D���C��k|��	Y�,�X,1 8D���d&U9:�н�Ə��YD$pe�2D��@�(��/����(W�3x6X(&�=D�$k"�@�����)Ѽ�j�K�B<D��k��"fO�<�r�B�Vq�y��E:D�(�ŀ�6,����R��,R���2D�X�F* 9c���E�^�R�h1D� ��ʽ!X�%_�V_�=��)-D�К�h�:%ΚP�ٯ��Rb,D��s�!I�a:<ͳS�X	R� ��'D�X��BXX&�HC�W����� D� *�d�.�NY1�� �����-0D� А�7]��@	�n�I��m-D�H1��Τ{5�e��l��A�x}�q�,D�XJr �?b~Fx�� �-��-؀/8D�x/=+��#u�سv�
`5l�)|�!�ۛm���\�Y���:�^�2�!�$��}^,*l
)�Q�dX��!�"�D���+$�*�LV�W�!��%+,h-��N�+|"���� �!�d�%l=̱�F���d�!��&�!�$�-6���#���#H�h�F�e!�$B2K>@G�Y�d<Y���?�!���qx�TH�+ģ������I7݄��&�ї��Ⰵ�Ҡ�(]���b!��ZS�R,x�8���D�x4T���v��qs��5}P������ȓ�N1{
܂E�xyILu���ȓE��[�� "5�� 无���6%J�f-X�%�h| !,\���y�̱��J�Ml����&E3�x��W��=i��S�5NTh�"P�g�4�ȓ
jq�wFBku�E� %�*h�ȓ$�8�*$͞�wtΡ�R+�'��X��r�a*t�ʈry\ݨ%�T3����B�(sE[�[u\Y�.N���ȓr%��3OĄ>�ٸf�Ũ-�|�ȓ"z��a�5/Q�r&�*yT�@����<�#e��N�PN���(�EI ~�<�AX�?�MP��ͷ�`�Z�@Lx�<�  	��^�dr�x�/يL́�@"O4�C�!G�����@�
��"O)!�JtB:�y.2ޒ�D"O��"�
6XXd,`@.��$� �z"O��"�<h�dQ�퉶���w"O���8l�bI6�\!R�"Ĳw"O�"�mX!]ָYp�V:� �Hd"O�a� Ȼ3�ldnڻ�8�+r�9D���4-iBTZ4�S*̕��8D�Ӷ��q�H[pB1�� �5D��C$�·(����D�DԌ|J��?D���ˈh�4s5A5L�N�{��"D�Hi���vmN�2�G*"D�!�K�%w��z�"M:)Z����3D��K3+WU;h��A �UB��p$3D��cR��3(�LY��M�',���C%`0D��qo�/b0���.����j8D��Ќ��]�*���)ǫ4Z}�3c8D��7��5k^0�����(mJ�{s�5D�Li� �+`~^:E��K~�PT�4D�����/: �"e��H���y2�	�1@9  �:A��aW����y�	R6hW�!����i�hq�����y�H�jP�P�.��d�25"#ݴ�yҩA� ��a[�)�Z �$�%5�y��B:w�ƙ�`l �]� � 4F��y2`�W��M�Hζ'�.�	S���y�'��-���*6�%jZ�C�gT��y������!U�X$�NŹ�O��y�Q'i���q������y+ �y�C+`+��z�B9ιk@�J-�y�!h�f���Im��O��y���!�u�6�_�)�
���y"��v���'��/Ң�Rڻ�y�O�J,��ID�|��8�K�.�yBm�5�H���������9�ybO3,ܞ��"�V�ݲ������yB�֎G��s4�7}cNa���4�y��8-�\�1�N�q�j�sN7�y�΁/Uܴ�P�G��U�`z���y/֊2 ��DA
K+≻n�!�y���i���M�m�]@k���y�`C6-��ܯr_8<I���yү
({�lH�E2p[8�����yRE��o�V�R�g=v�D�d"ڝ�y�ś�v`��v!�*�t}DZ��yd�-y/����33����
��y«�;J̮,�t��+�޽ �A� �y��&�,rg��m��`ccCɸ�yr��,>�ƨáN�Y��[�L���y���,
OB|AGC�P��a`�
���y�)�=1NM�e�Ñ3�H�B��_��yr�Z}����f��&����A@���Pyb�X �Vd�w�r[��G�<��hV�L=��R
 �V�H!g�J�<i��K�� � 
�uZ���I��O֮:T$�� �K0,*��݇�9v����C�&e���7��,,X�����#�ڼD\� X��lB�ԇ�S%�A�K�3"�-{�D��J����I[~ҭ܋{R�'��2^��P[s���yb�~#0�̸j@Y�'���y�#B6����E��4�qAB
ѿ�y�@
/��k���pA;�I�!�y
� D�p$�=+D�ʀD_�O:M҆"Ob�Xdf�;"���'Ɣ_R|�"Oj�Цh���p�A�Z����D"O���SE�z�:aF��(
��d�IZ�O{l�X�
��N� ؚv]�v���'��@��o�.5�B5��N�Z`�<��'4����*EX0�v��Yf(Ⱥ�'2�ċC\ߚ��TC��S����'��p*Dvl�<�Ƒ�9�����'`���JI�dB�.F]i�H�'���2/D.��9P�F3�h�p�'���s�.��L��"E턽E��(	�'\�$�ɕ��ܲSI��<��)��'�� X�-��y�Q��ٝ<��u�
�'�l��*ښn��D;��?-����'EX�`ٻ+wvɻ��ѭ,= ���'Lҥ�#�/Fo����G'*����° -z��EBU6. J��d�c�!�D��	�i�@ӠY��eJ���7�!�däP�쬚��Df��Aےd�'�!�סJ.(t �ԏ���YT�\5�!��ɫQ"�u▉<n���䀔x!��U�f��l���6}�liפ�r!�&4����*�8T��{��bp�}��'{�\�$���.��^;������2i�!�ğ�\:<�hn��3��bS�X�J�!���3T����$�~0:|:��\�!�Č$)[�mJÛ�t����
Pl!���_jB�nÂ.r`�Bd���|6!��Fy���HTm��pL*�PF.��8!�ď:3�����D	��iR ��?�!��(��ᘰ�?/͌0c�.r�!�Ą�P,��U���A�
�!�d	pi���u���0�����@,�!�dӔ<�h��&�	�zt
���!�DY�>�yCT�";�*�۷jJ �!�	q�`�qƣQf��R��Y7!���9O�:���d}}n���(��!��[���ȀnZ
e�s0*�2!�(L�t�/��>L�q����!q�!���p�M�P�ǽDe:�"K�Y�!�
R^D�T+P�H]�� P�!�$��I?��Y�L�,),P�Fږ9�!��W�Ҥ�'�)t�<`����HG!򤂛H��9Ӄ��xbdD[��;B!��Пp��8wl���ɦ���9O�*WIC�6d����k��a`"O:X�� ��C��� c�?⸙��"O��T��8��g��d�F�/�y"���	�`4�a:�N�ԋ�/�yR�T`��h'��!7h �
��y2ϓ�Βxb�P�^`��m��y���	��ģ��=\J��1�A���y"DS���=����CHDC�	��y�F��C"�ZAf�??S�-� /�
�yo2`_��¥AI�v�� oҟ�y"�վ=�:�x2���>v�ZcnM6�y�k��@�ly`�# :����2A���y�ܝ1���P*N�/��S��*�y�L�
�(����'ҮeJ"� D�$���̦oJ� "Ç�Dm���uC<D�Ȅ)M�X�j�E���}�Ȓ�4D����A��e
�C!e��qBy��/D����`F?`�H ���!���$l!D�� X�CR��C�pX�1O���lhR"OfQ �N��80�MS�;��,�F"O(x�!�!X�ᙑ�^�<�V�9b"O�H���Z(~���,�]4�P"OL��VL�SԚ�:Dk�xްP�"O*��#V5_���au逤/j�2�"OrP��"�'��@��5v�j�"OZer�ëB�d�9�lĘE��(��"O��	C�M*N�Fd�kT�
��"O©�E�J��9��L�r7�D8LO�e9S.��^L��"o2rJ�%��"O�svi���j��v���:4T:�"O��	D�����Ù�G0Ҹ�"O�� �D�E�|�bA�jث�"O~��r%�:j#l�4��?>!Ne�Q"O�ث��_*N�bl�����"OPy�� ���*v��i%
iY@"O�[ �*��c�>+��I�"O�ux��ɐ*�8��f��A�6Iq�"O���)B8���r���Тq"O���E��`��9�pG�"��	�"O I�q/��O&�11����\bD�t"O2@k�Jվ4���Z'�<{M���"OZI�p'_�ywLy���L�:Q�HS��|r�'-�9�%���k�,`�EAߖ��Q[�'dZ�'��<>#�i �((�.=Q�'�JÒg��0����- �h;U($�|��'�ND����"G��^�H��'i(�)�8y�}�&g]+ ��hr�'Mv�r#OF�l�qG��Di$��'��t��I�
�90���C&����'�D
t���лc���7��]:�'@�U��,���1�I�)4�t��'���Jbl��<熡�d�4_Y�ExK>1�8X��coÏS��	�"�A�|u�ȓYk8e�0�����ȋ�C�5�ȓ4� �q�斬\��
�D�P��ȓF�|���-ÞV���2QOS�
���%��3�eԜ���@�+] ��ȓ(��eB/-�L�"@Ƞ �f݅ȓu"���K�>20rP��q�|���V)�4��-��$����-|� ��ȓ=]:��iT=R�*A���&d�V��ȓ+)�)��٤?�$���a *�����c�@�Z���2|h͂%卞J��1�	����bu��뗵H�H'.Ѩ �t�k�'.D���VŖ��'�= p�IA�&D���'��8ޢt�&��!)810m%D�̉��ĬqF��'n��z�%D��3��P:���S�F�
 �)��("D���
�	_�� ��$0ش(��>D���1$�<%N��B�8Yt8
�n<D��6�@�#��|8��j
dD�W�;D�����L<5����4'����4D��sb��|�� q�b�tc��6��?)���O֢�!� ����� ��PB�'��		�!��Q'�y�p�@�x!Y�'��ⵡJ�":��b�˰P@��P�'�X��J!����I�T,1�'�	0!$��\�ve��EG�>|v�p�'->Q����ep4�����BfT���'��yJ��o�j��oF�6�����d5�B��xCc��~�ĉ��N8�(��ȓh�� f��8i��QIW�B6E$���S�? z��adۛo��@�#�&��y"O�xGE�6:��Є��\���9LO&�����USBd��ճS����1"O�R���%�����=\���"O�䑁/��'����-	��Z�A�����o�')�H��D�۵qI�l�D��0E��ńȓ4��!PC��
	��#����X�m��er��'Z�}��p�p/S�B,��lz�x�#W�M)�b'��$P*�܇�O`���eL�30�CƩ�!CF�Ї�ybU0���$:���#bI l�}��@�4��T2�`Sc��C�ҭ$�F{��*�Р�pu_+^q��*��yr��>O�qPa�ٞRy\�`U�X
�yə	�:���
]�AV����E��y2��Zx
��p�(p=�(Q���y���F�ё�;MT���b	��y�$Э!=�������3�2�*j��y�lH�fH�R���=��5���y҉�.�0(jQF�2�vݪ@����y�Ɂ��D�3�^7.*�� ���y��PaEX4�� %�6l�b�܉�yB�� :r�S2�2�8!C�H��ybFX���B�c��flD�-�y2��8Du*a�F�ij���w��y�D_ND$8��I�S�j�kֈ@��y"�׵[�Eq���I~�-��̤�yl�%<�̄kB,�B��0(����'���t(N�����i�:#O���ȓ'�����Kfp04�@H̝A�0�E{��OcJ��$�6��0���F����	�'dB�3�O�/@�h�$��<����'�8��F�5Y�������~��a�'׶]S�@݇�nYa�ٯ�,���'3�@�3���lw(��F* 0Z��'Hi�޴G�U���$`>�8�'��ABBl��g4���r��g�� p
�'��pӮ�"m%�ib��d�J$��'�t�%OŊ�T!b�G.K�H���'\ ѩ�a�{�x-��Kβ=��ي�D3�[����˝>��2�(5�h���'�����N�L�=�t���p��ȓ�lUs�d��U��`����+i��ȓh,�����L!�X�`)��.��ȓBΝjg��D�l��e )�x��@��Bv�نs�U�D�D� �2m��<m����γ]�<����z &U��o�P�k�`������i_v �H��6�L���� v�S��ٙa+�0��1[а0�FS�]�c�oH�5��ԅȓV�
ؒ��ҥ1��9��ە-���	`�'���R#(�^zzuB�߹�x]B
�'�]�H���ZٙÑ�A�u�	�'�L�i�n@!T�&ea����Ի	�'3N];PE�P���QLB����	�'��
� (3�<Q豪V5{��l+	�'�x�H3لI^�A�ԇxNN���'Ѣ1�g+��{�мc�wH^<�	�'6���aT
H�a�(�{�&1I
�'8 %B��R�L82���q���	�'�|�+񢕂C�ay��_9V�y�	�'��A�*Y2g���C��O)S	�'(B��D� kdP��-�+�pR	�'~D�"�C��W1� P
0Ǯ�B	��� 4̓�G� ��!I���#%\�PE{��+'͢%�wH�� �"��t��z�!�T:N�"���#a늕1gʍ�3�!�Dطm��9p3éQn�	�v���\!�S{^@�fK\+0�i�c�\;9
!��Y�H�C�d��htC�6!���k�̀)t��4�h�c�D!��&qpvtjQ��N��#3��
9.�r2O���p�T�a���R����,u	`"O���7�גK�	�I���W"O�h���$Q��Qe�,�v�	�'�R5O�"�$C.��}�wƑA�0�s�"O=cC/�&i����OE�n���"OH��e^}�z|[�m�!�\9�5"O���2h�1Μ��%��Hƨ�Qc�'���|�X �Y�Z �;���{2!��
S����#�/>|х�V�!�d}2�$�2LM�  � �G倦y}џpD����2E� A� +Y�Lr#���yR@�4r�T�sf�8%�0�!DcV��y*PHmz��2(I+MPU3遡�ybgո_\<\2�
�f��1��O��yrˡrјr-S�	�Fi�Jʹ���hOq��y��	�/ḁ���F�j1n8{�"O 2��	"��P�fτ�F���'��8WE.�I���|�(�CkR�k�!�$��3� �↸^|l�F�Oe�!���2BΑʰ�V�j���	�^!�$��T4�W�Y�����hX�R!��(;R(�!Fz�.�Y���=!�d�&~����Ryм�z&]�!�
�z�0yhfȎ-�Q�9�!�L>J��a� ��NР�G��+,�!��X����Ŭ�.I:��4�!��8�4ݱ2E��OՌ S�$+x!�ݫfx��nOI�Δ�q)�	cr!򄆖T��Hʷυw0��rThFW!�DJJ%�$��Ïh&�R���TX!�L��I�`*$�p�"��Pyb�D�y���g+�,?x�]@�aD��y�ӷ'X`F��ڔ�`Ϥ�y⍖b��р�mQx�B�����y"�5�V��,�`��0�-
>��'�O�c�2��I�5�L ���f"�(77D�ʒ��hr��8$�H1�S�44��p�HG'z�R���W���Ԁ�p�<�0�/5aRC
O�D<����l�<�%�OH�����J[m�HY�I�N�<����1
ʘ`Y�Ɂ#��!���H�<���յw�z�i�R&8԰Xq#AI����<y�j<fH���ԐE��ŜY�<)U �t"�!���(N���HLX�<y��^4����@dHS���_�<1DD�^� 43�
�}ـ1K�ȟZ�<����C�2	6�0a�0[��+D�,���$J��R��[�4�Z�.D���Da�j>�3�M�7?�N�K� D��Z�H��8@���eԆ-<B"<D�TR��y��%�3)�$��Q�c9|O�b��&ȿ5��)Jb�ſ�x�+5��V�'U�ɥ�� ��j�cЀ�+�����DC�I���:7��"\a����!*\>C��2i��@�� RL��5�P�\��C�	z#��ҳ�_�[:Y��J���C�)� �r��G�Tu�VH{G��"O�p�v	G�v6,I�����q�θ�C"O�\��M+�: �
�~��sb�|��'��G{�\�Ҍ��f*�$i���6F�!��^9u�|�a�39�T� EM!��ݭ)��X�,O��<!#w䛈H^!�䂚p� ��e�]�x��UxF��!�$�Uf�d����'�ra #h��2O)��O�$�}hR(ӿ/H��!B"O�)�G�
|&�H
��
-�,�"O��v,��6hȔ�LG���k�"OB�R,�.�.a���8��}�s"On���G�"	u�5����3B@��t"O"�v��@�,US�f�q.�TKB"O�U�nݲ`q�q���� �"O~h�ħpfZ���. )��"O��$�W�j�Fui�Mǂ�f}��"O~@��
2Ak��Y3��"��Y�u"O�<�� &�2���̢y�H�"O"�h#�4�01�Aݛfmn���"Oj�C2#�8l�f�c�
T�g����IX>�cd���`�LX��A	���$D�`P�@&Nhji�iH�q,��rV!�D�O���>)�q�J3��ɵ�K51��? !�ĜP��X�o�Z�P���	Z$s�!�$��E1Z�
��'Ѳ�3�h�:5�!�(Cn��bB�� �L�%h̕9�!��ʖ&A�G�I�%� aȲ�Y��!��6d=�˔�>dG�ЉG��72ў��ቕYZ\b���p�`�����	"��=!
�',��Y�N�,(f/��p���}m
��!ϊ`���Dn��K����ȓ� U�w$�Ty��+�[�R��]��;2zX�K]���O!s���ȓE��A��X{�≺V�9O�Ňȓk߫�4{n�j!@��z��x�a�IC�s0Ă�A��0�o��S�Z����<Q�
g�����C�Phk@�;ݬm����<���)����b'U�DF���dC�I/ؒT�%�.&L`5��/A!bC�ɑ�؀��G�9+u2��/whB�ɋ�Ҡ@�z�\��f�P�7FB䉚t���w���V2��c�'v~B�4���cA�My� �C��|K��=��K]u3$T�6��&��|U�ȓk�V����(W.uA!(�(+$y�ȓ���Y'�;خq����OM셄ȓ�\�Q�-��p����$]�䕅ȓ<޴��N2L0����!1�<���*S��C�m�y�D!Yn��
�'�p�Zf���2�LD��Ė"mܚ	�'�	�1%8h���R�Z�hD���'pVl�FA�:r�d�q��J]��c�'�t}8s�½]���Iڀ0%��'��-G�\	��
<׎�'uN�2F��2M�a`r��"/�Db��:�'O�*�@��x��`�ͅ(0@8ͅ�?`�/�*p�2)+P�6���1Xv�����6I�L9*!�-QJ9�ȓ��̂�F���s��a>}��"O�x��G%舕����aL(��T"O  ���
�P�a��� eT��"O"0B�� ��m�o��Z�"O��p@�M�l�$@���M�Q{U"O� ��Q)��gL��pG�lE�`"O�<�"*F!1�]s�lH0QE�Y02�'�1O�li׮�<a�����˃�o*��ʰ"Oh9�eD�,F%ޑ��͘�(�=1"O�)��&��W^�a{��S*�s�"O��3� ��$E��ɒkΝN$����	G�Ob ��6H���TV0 �6�;
�'Nh��i�DTPɰ⨊3"��Y�	ϓ�O�4IF�C�"��i3��ר=�^-���|�'#``	�3Q�@|��.����'3$H��Ș�D�Ҥj� ��!�'��<�q��_(L�2�]Ya��'B�;���"13�D����%�N� 	�'��S1�K �^�� �="'�9x��!�$*j��n�!8��\|xt�#D{�ID�'=1Od|��i�2�~�I�oW8-J\EpT�FB��#�`��]2�B�!ƌ??$!�d���� ��j���D%�y!�dB�or��Q	�vL0[u��3!�dn�����&<o��a��ܵF!�$�E��y)�Y~mP��D��l�!��թg<��D��'^ UICn��N�!�$>O4�A�sOє�Ľ*�mT�8͡� 1E���$-���m	����y�����Hy�_u����`\�y�o�-$J�����ɵ�\��y2�5k"��4b��|#�U��F�.��>��O�aPm��&�����
�~�lY�"O��z��=[��=����h��b"OlLI�݅v���q#։OkN��"O�x����2@HT�5bU����"Od!͋�I>�Y"F�6���P�"O�E���rh�p��#T�2 Z�"OX(�炣==E��@B�yt��Ye"ODt:WO�y=�� �!	�@Xԉi@"O��Q7)����aΐ�d)�"O6t�t#φH6�p�՛6��X1�"O�p�ς�K�޽��D�a� l�3"Oj��1�I�iWZ�r!AI=`˺DaD"OI+�D,$��o�b�^=2�"Of욧o�)-��"�S,'�����"O`�Å�M%;
�}�wd�" �d�`"O\��f��pD�K��J�F���'�ў"~2�`_0yڜ��d*r(́� ���'�azrf��%�8��B�Ĕ~+���u�O��yRo��tx��3��o40��ӇO�y�'�8~��D-ŵd�.�j��j�	�'�X�Ȗ&JOE�aр�D82%jM>!���?��7v$��7���9�a�)oXI�ȓXY�Ԑ��x,j�Y�
R��F��_搅S'�Rz���pI��)�C䉆)���A�aܹCw-��$�B䉖s[��0�Z:O#�5(��	n0`C�I�U�
�3�Ԁ;�8�b�l�0��B�I�}��A��ȕ�JS4��odh��'e���H�D��z��P��N@�)OR����=���h�˗e���6bA�}��� q�	�@!qA@��]~nhI��6D����j�'G pHQJ�$7Zx�k/D��h�CI�O>��x4�H(��j�-D���뒌Yy��#�C3X5Н��J+D�d��k�(�R$� : �T����(D��9�Z3T�P�c!J�3�8I�"D�`�Ђ�Z�|�F�^�F��s�� D�� ,ѩddÄF3lQ*ao�y���d"O	�)Z6�9�v-SV��1�"O١�GjՒ�.8'����"O�<�3J	�$q�dB�G��p5J�"O��3%�Y�?���b�6�A�"O,���� >g���`��*y�Xkw"Oj���K��.�<�㄀�/U�`bb"OH��EN�f�L͙C�/-���"O�}��m�IK�+{��:����yr��.3!����X�x�}Q�+7�y��@�UԐ![b��� ��������y҂>Ċ<I��xi��K�%D��y".Ϯx�mcT�k���C$�р�yҀ׳O�<A��#p���o<��=��y �k�ɡ֢N(��-1�����?�S�Oa2�C�^�<��Q�G`ʃ�f�
�'X�葂K�
Xl�RתQ%�@
�'�@ $?�j�Ag!��v�ހH	�'�Fd�1�
p�9�6�o�J`
�'n��0Nۣk8�xx���s��܇ʓp�����I���"�؅���CC�'�ў�G{��3FE�@)WÇ�.A`�%��|�ў��'p�|���\�u�,�Y�íaA��3��6D����䛙9�0dS�KB�qfb���4D��r��˜���!f��v�p	�E2D�`H/ɤV����j!Jv��!$D��I&�ŨR�\�6�n~���n"D��C���H��	"���4#�Tq��/"��8�Sܧ��Iª��x�S��%U*^X��]�92�ʊ�"��S�@�}DX�ȓ�Z�9��2)I$0�`��L}�l�ȓ�N���ަ"�M	��֣9HƬ�ȓ��eǀ�@`	�"��9I�z��ȓ4���!#��H��� 'd�UP�-��u�'B��éߨvۊ�6��ZؒO�=�}J��6ux�y6����<�d��Z�<�P�.�&dȩ*�����Rn�<�r�϶A�X��գ<!0�ı��Ej�<YDo� ��14�V:�X�!ŀ~�<y��<;�5��15ܴ�zrMz�<��jI>�&Ah�Uhv�ʡ�MA�<�A�ՙ(�MKB�ͻ�#�w��0=���E3Z����
�@�A���p�<i�(�+I�!��F�	:�ĬQ�<�4��� m^8o~�ȑ�w�<�`HĹ|f|,��F��U��a$��I�<�r�0P�OD;�H�B�G�W�J�ȓ@�^��B=�V\�bE�gY�`��F�Y� �]U���`1��-8�P	/O.��?��'�rV΂?;F Pd�-L�Շ��m�'x̀هK�.+"*�j���TM��'i�!��b�~@�*��x�����'�>�I`��Ft�!'�Z! �b5��'���w�1#�~qŢU�wِ���'�=��	�8Q[Ĩ�$G>j���)�'W*�Z3��5OR��0�A�<<U�	�'�l8#Re
9�B� ��v�����D�O�"|�O�	�n11Bj	6�
@�q�<�u��7��m�Dڳ���� ��p�<Q�͖jт��*Y\rTbIj�<�҅ۃr�����@�*i"�m"�BNe�<�`��G�.=���B�.�Ѵ��a�<���C���4��6x��)�%蟨���Ywv��" !P�n!c�'�-�X%��S�? t�IȂ�2Z��V��<��q"O�u0��t8q���;XR��#"O�!���b�~1y��[����b"O<�3�oP]�<���+�̑$"O���R��u2Y1㊅@���C"O��U	F�~0�(p/�/�����"O��JX����3*�!f<��A"@��y�E�<e�D�?�-k�f�C��(M������ڷx>��)�ds�C�I�G�`�M��@S&9����7��C��]��Gh���d��R�� P�C䉀O"�9X��A�1:�3ER4ɜC�I=:�<i�Z�<H���A�6|.�B��O�p�5�Ƨ<mh��U?�B�	>h@��j�,�cP���@З�B�ɏEP�!��T�O�0c�g͇G��B�ɳi���A&���Q%T���	=[�dB�	�g�P�a��?�&��Q�4k�\B�	�:��䲖��Y�|���lA^B���0�@0Q�	��5��b��C�9_�4�@��Z�|���E����C�	�K��Ś�LN�1�p��	��C�	lL�R��N�+gDwF�1I�C�&hUx�;$O�[���gd���\C��G��f�Q�X�#7f�(V�<C�I>q*
�Rv��xQ4`K��S=	8C�ɂ&C�y�C�e��v�8'��B�I�h��x{
�n&�%
Q��B�ɷZ܌8�O�������^(C�I�P�<Aj0f�+%0e�+��B�I)U���X�c��0 ��Q�fU�C�ɱc[*q�WM)p�Xyr�̒M/dC�ɥ)x`i���$	Q��	G1�PC䉨)XT$�G�E�07<ە�P�C�I�k,`��N\�{ ��Rą�P��C�ɰ)�f)8�"��y]���%�^$0�C�ɚ6`j����$Tw�Q臣Жr�C�1&�8]�S파r4�[��P�sB�	g�Nq` "��+��#	���B�	8o.l}C*FZH���4�-�DB�#x:Ԩ���]	Z.nT���I��C�I�}��r��=��(C/@<$�B䉷K�\9SM,�d�X3�.l�C�	9O���:�h���dؠ��t0lC�ɼ2�b��gh��k��{b�B�a�jC�	>1EY����|r1�g�8�4C�I�R�H�����\90t'�u�C�I�S��ZTe�?2Hl�p'ȥp�B�	�'Z0���*ܔ�(w�G�Y�B䉧2h�4�@�O-^t0�4�"R��B�� 9r"�����Q�ت�hޠo��B䉲9/���ҍ�),��="DAݵh-|B�ɉS�� �]K�2�s&�۶A�~B�I� Ş|ˆ#�1=��r����+&B�ɵ@&�4(@�O�
��ܘW�xc\����D8���\�\���&6���3:!���=H�̺�T%l]T��lXu��ǔ�2�X�j�A�A�a���X�k�荒5$�3@�G��M�ȓ{hiۑ�P�mE�(h'̌5q> ��ȓw}��y��,�]�/~<����:E��N��w2�����o�H��ȓ!/L�[�̓E1�)C��!�݄���d
�O?:@r(sGn'Y��d��S�? Z �6 R����1Gˉ�0���I"O^�����gȊU�%�ۤ �Ա"OR���}4B5@�D����B"O�]�H؏a��䅼Z}��"O.iʤ'F"_���� (�3w<|{�"O�@8d!W�N��ɑ<\l81"O0m��� B�(MōZ�q����"O|�"s� r�(������"OR1(�"�+z|�e�F�z�:�+6"O`fkʟM���c`$�:d]��"O�����O0�����	H"Ox�*�
б5Uq��>pQ�1"OX�i�
W
��j#g�54"O���ǧz!��!Щeݐ�"O���LՕsQ�Q��(��PQ"OF��
V3q}�9	㢈&|���"O��ʅ�?�M(ӡI3s�&Tp�"O2|��N	�� ȵj3HJ��B"Oj�S`�!rVE{�LZ8+�9(�"O��@��Q�v��sU�Y�^),��T"O��c�"׭y�����!5��d"O��q�	
d��I�%W1�E�"O^TtǞj�0$�B�şsŐ� "OHM2�K��'v�$dг�N4b"O�S�L�� ��I{E� a�"Op�᳄P���H@+.���"O�A��hR�Aw�ݙ(G�!�A �"O
�ek�9X��-KeFI�-q�ԑ�"ONK���L�4$��#ҡ
�r!s�"O)��+A��L�b�QraHd"Ob\��I]	*�4MR� �vU��%"Oq2�-Z�0�؋Ձ��=N���R"O�ED��8hA[3.�1'"O�)! ��+}(��Fo���xX�"Of��S@K�$"np��J< �`E��"O0�7�$YׂyCMѫ#���s�"O8@�7}���s��S�����"O�̋�@��:���ť�A�"O=�F��h<@8Qc �`̲�Z�"O|�2��K<8ed
P��)oP��b�"O^�sqB�f�t���}Np�s�"O���Cַl����!��+����0"O�D@��=�`��R�
� �D`�C"O\�J/�,�
U{�.�2��,hq"O�,k�hU���#���:�
T "O��3�R��r��ìQl���"O���1�I1m�䤈�oɰ)Y��"OH�9N�LK��0vF�LZ�0"O��5(xP�P�5��Gh
m��"O�����Y{�|7�ҳS�j9�"O���O�s��Y�,T�U�L�G"O�Q#〉v&��aC�T�|�<E�"O�����s��� �I4�Q�T"O4���bɜ.�����ΚON@9	w"O��g���H�!�p�?c2`� �"Ov��nPyL���N�:`�B$"O�Eh�yY��I3�&1���2"O�L�$ɑ +�X@�X�N�HV"O�I�#��F���q+ֹ����"O� �Jʾn��`�R��4i�4W�V�<��� {Rj=A&�D�,��S�I�<�$@�hIF�6ȍ�xfA��G�|�<A�.2 `+� �Lz���-@�<a��8F����I�22B�:%��}�<� ����H�
�bA� %�4ŤlC2"O���Cђ?v�]�E h\ زS"O.�����l��Ł�d�Q0$�)"O��8��}�,��Bޝt���P"O��#4nˏz=�Q�k62��%��"O\Dؗ�Z��1y �V��<Ó"Ox��JS� 0!��T@l��"O��!6�
s�ޤK#�?%H���&"OZA�'�\�}��� Q��YU"O ��Pd�J5>�R�/SA$MBr"O8���8x�|
�-C:Q-�(
%"O�%b*��G葪&�[�q@d �"O4���!Ay|%"�KEo^B9�"O ��ǧ��Bn���/kR��aA"O�	�2囇^�$�8-�=E�6y�P"OR��u�6�ֹ�g�G�J�^X��"OZ��𮏠P��,�9�����"O.�[qT�)f��: ��b�ny�"O�8۰��9�.]���Sg��ԛ6"Oބ:�C��c�l�H&�@�6�)�"O`�*R)$lV�B
��R��0 "OVA�m�,^>H���I��Q�2	*D"O�T��l�'α��-Y�:A�r"OJ��W$)@Q\�鱌�-�a"�"O
��r�8dt���G!�j�z��"O����a��;���{�%��+t�ur�"O2K�m���E��D�2f<|ae"Oh<���@%RU�T�vP�5"O|<8�,�4Q���r �Hjj��"O��i©8qU:��p�C09i^��"O�)v��A�D��D#]7y���"Or̺3���1,쬓�,fX����"ON��2!�5�"fǇ\P���"O廦g�3X�B��՛
7�*1"O@z��P�QM@�A@��F8d�!�DʏR4T�&,��B��I1G��!�DΖy�9�A;R̸�I5�!����	�B��/�P���ͳ�!�� �:��4��X6��@`ۮ!�!����P�2�U����t�]�n�!��$n�E�a(B� �U���!�{������*� �U�!�!�ٯ{|���-�Nl��[�eO��!�E�X,�8�m�GV4������!�T�!f��:cIt�F��?
!�C+	�8Ma2��1B2�#a�p!�ə7u4�3�h�'ya|1�R��69T!����,�c����hc�tF�'|�V�)�:]jdY���.�8�vo�C�,C�$B�H�BԣL5�Xg,+�<㟨��I�(��$zw U¤�CSB8:C�I�*Z�Y��$�̙  T�4C�	�R�pa@��ՙ20����	�;YV C�Iy���*����>,�w(�4C�.5({�iݪ.�����NB䉶��l��Ji�f���lEG�DB�	�+~���`�M�C��&�����>�4%Z"52�}С�@$�ʓ�U{�� �'��`�1@�g�|袠J�Z�Q�'θx���6�E#��:�1��'A��C��s5z5B���?��3�'�
���E�B��s�\�9��ջ�'�~E��'N�4�<��!Đd)|Ez�'ʸٳ&�Y�z�B�	�*5^�x�r��� �=�ʍ/.$H�ҡ�>K��U�"O,A�"[�(�6����#V�ށ1�"O!�W��-�%ɟw��"O~4�I�#��Y9��B�MC$@�"OD��Dع��̋ ��%[&�ӣ"O�,;!���I�R���Oٍ&�Y��"O����������q��j�q[6"O��r��D�+����ѭ�A�*���"O���㎊�<'r�)q�![����	.~�Q��VA@�ȁ� �i0�pi�EA,?��9��i5��P��I?g6liF��݇�jcHtr��	���[�ꑮx�����mj�[�G�ͮqc`�N)3^<��K9 1:�bV
m�9s���%J�� ��I{�$g]��X#' ^Ӽꆎ�8, ZC�	�SOXXƤ+���6�2^�b��D<�V��e���K�@#�\�`k˒a+@ ��Iu�'d�e+L�-	�Ŗ��1Z
�'K�512C*<� Q�DK:E�>��P��$�>E��'��! jJ�[{�q�0��5�,���'���y��ڇ\��X����6� ��dڡ�HO���r���b��w�K#�̡3����B�Ҷ��(Q�1p�[�a�ц��	���'��?��e?�z� �3~X� �	*LO����ͬ@vH���]�1;a�;��`��"<��y"� Ô� 	�g�̕b�i���yR�Q��=c$��I\�9玀!�y�kC>C���q��ˑGs2�+Y��0<َ�d*&�U#�$p��8��e!��	�9;��\WI���W�%h!�D'*t|���:2J05�&�R7{g!��,O̊�P¯�-YB��B�G�Y`��c�'�̉��>��\C���	{��i����<�'�1��x&FC�&e�-+7�K	�PS�"O@�R�p,�h��c
N�!��i����<�۴��?7-^:��Eh׋Z�]���re�&88!�D��p�j�"@	�咴�@e�&0�Q�T��	,���{��Z8%����p�	 �C�	w��h��M,b8��3��z���$�S�OK(���B(I�� 1�Ԝ[ Ԝ�"O�`:uB���^$1��ӣf���"O�`SOڄ+��ʄL�~gY��O��	D��<�L<ͧ@F��2M�l���C�ئ���	i?Q�"�5RK.!:�å8�RT#N�P�d�hOq�,�ǧ�z&��\�\�����'�`�)�N��B�:T�xC�Ol���<Iߓ0����3?��᪀c�r�F}���E���A�e[��t	���${�C�ɴ�^� ��W/\�;3�Ɔ*��B䉅���J9j�B�S�@8o�B�%~ �Qg�T#$����b�OSBB�IRdTq���&-�YJDcD�K��C�I��i8�NM>sI�ģĬL�(z�c�HF{���ǅBN�!7 m�H�p�gI�yRѻT�
��m�(e��A����'!h���Ib���xp�O9)�q��ŕp���$&�S�O��V� xU1�l�T4Z�� ���y����l	�p�\H��9����~b����O,#=��F��{R��C*�Ds���-U}8�$J�4i2�+i�ġ���M�$�D���1��:�S�'oA�H#a�;�ģp.�/�ƸGy�
v>m��k�S�ʬ�E�)�@��?D�hsC��}�ڹ����8���d;D��K��U+Q��+�C�)��3�:D�� ~Xi�;R���z֡R=g���"OH�j�eK-�T��^�R�����"O�)a�H�m����� <�4R��xR�'�9�b�ͺ0�����
.=)�(���?��O�,�R/[�S��I��k�
��'@ܱ9�!��3y*p����+1^\@��$-��?�n3C@�p��!��P�B;3�DC�	'{wXi0Q�Ԑ]K*��5I
'V#?Y��(ڧ+w��IA@ȟ{���f@C�,���L����w G6���:�n�'[�`��'aў�}:s&�8fHe5(��p��M���XK�<ai��Y�t�㋜�P���21�WH�<��ő���u`VnʉJ�Z�!ԫVH��$�'��	.�9���=��e����=+,B��
N�����/ݒ���Jb��c�ϓ��'��'�J]!,^+_K�����04�L�Ǔ�HO<8(��!9����+Y�uf@��"O�x؁$Vf�~i��	�.X,�}��Io�����E������#w� )�׀G+y�!�$�
�)�-��1���A'�!�R��|!ˀ`�ot��C"�/@�!���MM��oμZFHM8E�L=l����I�\��(�N����s�&øB�	�n�аk�F�{~�3��C?F�v6�:�d��ݖ|i��p" �F���m!D���*\�,���$S��<Ѧ�*D� ɇ�ʔn��P�T��T���&*D����)��-�A����d��F&D�xh��)�����(�"4�׭.D�l#`�]�1����fQD��#d�!D��Qt�I�9�r��V��I�f��M�Dh<1a�ӻV(��/ȸ-^*�x#�p8�H�OT���.�7[�$�:����<<�"D�t*fB�$wh�!P�+\�zk�$D�Pɷ�{� ��j4��)��!D�Ăq!�4H7�|B�̓g�8�f*-D� �jͧjI�h���^G[z���I(D�T�r�O�W&���dK+YD�1�Q�#D����K.B�	[�kC<PLV��2+#D��[E�ށuN`�Vi�n.�i5D���$/��䐸��ߘp�^��w'4D��{���37���q��L�VY� �0D����a׬W����A�?��#��/D�,K�F��U�L�@r엽D0Hu�#8D��)��]M�����?�x![1K5D��!l4!���*#J�	u4!���.D�D��$�)#��m�L��,-+qO2D�XpV��6G�2���&W>�vm/D���p.����0@�F!j�h��d,D�T��Ǜ*� �C�y���*D��@���zfv�8�,@�3�H��*D���� �?s�X�����-Q�q��#D�4�B]�	��x�V ���5D��z)�/X��$��%�F�x��6D���gEz�#�ɖ6��I`J*D����0i�lX;Q�8>8s�I(D�P�@g�-����"���7�P���:D�<�@��1(S���t�3:��:��8D� �B��e�����:W���a�+D�+�b�:X���e��f����Ѧ(D� K�ÃU��Y��"��%����	�'��<STd�3ʜP��E0*Dp��'�!̗�6���f�%xD	�'���e�	H�J����ݖ�4���� 
q�0�[�q����iQ8�dR�"O�XC�F�3�4m��J�"��"O�����T�tB��`ߦn���"O�q��`Y�R5j<��i�:���h��':��ĩ\�Q�f� bl% VT$[p�:[���u�I�Rx�%q	�'Tf��5�� � 0A0oU�Uz�dH�'4�Qb@�oZ��G@3|���c�'�\-
��'��l�_|ذ���'Q:��6��S'ĩ�f���-���	�'r�A�R�Ak��B��U�
���'S 4�0cX�'�&1�L��E��'V��է�����V,�\�'0�q�S�D�l���@�Ў]��'{���6d jL� �_H,�l��'~0�� �<�\Q���Z�2��A�'F �)Ѐ�<ꖔz��R07_ĳ�'�R�Qgc�%E�ġ A��%�.� �'�*�� �!q���լ6�:�`�'�ށPM�;�|��������
�'��kek�XT����r���!
�'��]=-6�$y��I�y*���'�X��k &o�1G��5%@1��'��9�d�= ���P�Ϩ\�B�r�'���Ġ޿-�����l۸B1�Y�
�'+� *�N�}˨�z&�L�;�FmJ
�'~�)��,�%x �yq 
�*�nt��'uh�H��u�v�iP���Āqz�'P�I��h���w (c%��q�'��l��U�X����M�"�|P�
�'D�T����;��)�e݌�-X�'�dA��h�쑰��[:fHY�'�����Z�P�\� !�(UH�'������V6��z�#Qr44A�'HHt�Mۜ� !��l��C
�'�=���V��i�J^?[���'m4 ��� C0�����Fp����'��@�B�<4�^h�c�7
h�x��'; ��ǈ�5^��5�s!6 ��a��'�P�;�'�^���V9|[*���'��$0fJ��/>J,��mz�(9B�'���MO�x���V��/�f���'OȽ �&Inf�� �M2��*�'w��'M�#��Q�' �;��A��'�ʵ����<z���i͝4:���'�l���(ܵ|:��)6&�<7:���'w��P�G�pa�i�%�
��U�'g )�d��as���0g�xa��'<<p�[E���ؕjX\p$i��'b ,�	��ٔ�Hz���'=�IS3��<������#A�����'�F��!�хC����*�A*�T��'��� ��)"��Pࣦ��1ˠ�[
�'��E�b���Rt����<7e,	`�'��AR�DM�a�����A�u� H
�'�.��c���ҍ	�(H�]�� �	�'H2��M��Z������4��
�'(������_*m��B�K�4�
�'��A���ޙn" �\91R)�W�)D��{��Fg�*aD�85�TY�P�)D��!�`ί2�]i�c�5�"�9d'D�,�K%o"����.�JBj11'0D���#`�$.�84m�Y�$Z��5D�Tf�	�,���Ώ8��p�F	?D���dɀl?����/��B�8D�� |]�)�D��2ė�b���v"O��J�d@�r���2O$}=���"O�]Bfd�`�
 �&C�')���B"O���A�H�Rf� l+$,���'���H[
���?i��$����B��00']�B��Dz���F~�����GQ��b����g�S��,Q��S�M��]��GԻE
�8��X8xB��>f7�h%��z��B�jW9n�TH��\�U�2h�/O�Y{A)��pX�&>�'�t�z���!vz�Qq
_9?,|+�����M�R���JAhR�h/���S�՛[�Ơ�GaĲ�2��v�X)�0>y֎R ?�� r@0=ހ٠�ˉS}r�و��FLƥ\L�8�O3� ��̎4f:<�Z�4�v����5>�P=�
�$Z^ʥr�"O���"�/zO&�I���4����ъ^.6��I��t<3m�;;g���ҟ���26��˳6�Bq�үS%=��+��r��{��'��!*�m�>x�@�B��5��	g+*���Gh(Y�)�a��q�R���h�{�N�r��4��>��5}���]^���Ǌ����ؘ�ڿ����'�J�2�P� &0���IP�N=��@���>j֐�q�N@�]�܁�&n*z�6�l�s7�'��ijp�;G$n���)c6�M;�'�6�[$V%��z��X5��aΧG&d� �ب`0�E+��Y'{���d%Lt��`b�،P��\��ݟL'��#&x�Z�Ѣ��!��{��K�5r}���ަy�W�|��@9  �,M���E%B&|-�W�H��Ɓtf8uq%m�r�����c��}���a�|8�fͶ_���8 �ؽK\"�*�� �T�����$%C.}���̵Y��h��Y�I^*��ת�<ѱ���EX%�׌47t�! E�'r|���$}L1��C�[l���7P?�y�6��0@V�0���F�-#�ߖh��ɮ��
�-�0�џ�{-�R�������Y����5OP �k2]d�0��^-x^�7�ڋ�n�Cfk�W�4圻b�J�`֯�F��S��PC��z��0�Z��kvXP�
x�VB�}�xYZ0捲`;�m8�n�%i,B�gI֦n��]bP�spɚ�Tr�M��Ok�o������&�4KM	J@�}"+M�HF�5�Fi�!yF�t)��T���k��7�(��d�7�V����X�Cs���QS����j�F��	��V��1�k^�]7�y�F��2]���w#"�p
�gc��|U�}�$L�4��ɰ�GA��t�ڗ�W�N��/\����ʱ�W���$��rL��'O�l��KA>D�P�4�ʐ~<��2O�c��4Ii�$�G�/�`��K�<N�H��?u�b�)f)��@���:H�� ޴V�^�r�
O���/�3?fȤX�EEc���;�!���~-���	rQJ�HvͼV�S�躼���:?�4E��1�H��$Ǝ8޸��1��A���s'�Ll\*�(�%i4}i�g��v�x�!$%Ǧ�q�F@R${r���֟@Pax� �	T���`d�9W�,d�9��O�Ȁ�
:J^��ӥ�gJ���2���hRJ=}��3�n$%S堚��x�c�Mb����:ƺ�3qk���D���|�av]�^/>��p��5�2;�N�]�'M-p! �^+�b`�R$M(s��t�ȓ0N����O(*:|(��A�R��[#�\�Dm����BC���5�	}����'�b��#ϐ�?�$XU	�&qD����'�f��s�m�r���Y%l�����l:	�&iƞ*���`raVxk\$���+�,����O�G�h�2n�`�p��D�?�ъQ+ԺW�q�����	@��pq���@�&I�ӣG�+L��!�?$����- ޒ�6�=M@(�� 1�IK��)(t�ߵX{r;�ӱT���34/O~<0�é��VC䉠mY�9I��?*t{� �=���6ř�G�\ٛ�@��~�\��ϑ^�$b�΀-�ƈY��-D��[Ƨ�|l5���)	��O�<�G�בj���pៈ��<��C���M�f�E=HMH�a�ϐ{��Г�DD�E���@_�
X2���N�>��CkW
~B ��Oܝ�# NК$DB�>+V��Qቪ3@����-�%Y�����V��c�h �1G\��y�k�'�`V_H�ɖ`L�~P�-Z�K&�j�ˀeTn��S��?A'Ȉu3��!c�%V�Q��x�<y��|�~���׮o�N���w~2a._�&���'�P�� T��y!�$�N���d�~QRE�;��S�j�Qy,m�Ї�5z�VC�ɱW'�}�Z�z��$f��B�ɌT1x+��[:�f	R̛�Z�B�	����Y�E�Bd���[�JVB�I�en !��?%/���j���B�II�����' ~��S�O�<��C�)� ��)w�Q�>��mV��("Oڀ� �ӨW��&�6@�"O�Y�e��@����ao�*V���"O>h;c�	I�}*�%�(bQ����"Ox���^=yb��Ό�[��@��B�,b
H(Ó_�N���FE�-���)!'�+�����_�F�z��Q�6�:����Y��R���E��`� �����Y������#5�6hE2��y�h����gⓠh��FR� L��!��77&B�.@Y�q�!��h�a�K �+2�ʓW T�1��,|�ҧ(��-h$!��Gwlܨ �B�+�H:@"O�hqU�����Wh[��xЁV�䐹=���� �-���X����C�h�;iE��1C��l������IA%�0�n�p���_\,}#D���S虇�It�(�`fѦ6�����K�E�̢?�`cB��T�C�#�i�u��W+�͞����35^!򤗌 �6�1pg�7�B(���<e9�I�[��=Z�ڕi��S�Oz��󆤏G�jҢ!73G�y��'�`+�@��%x4��ٿ\G��:�*&}"i��|����%���{2ኜ;�~	�M<Bl�����=�x"��94��,R9^ZDhJ���#KRū��0���k(.`�K!b�>��Bo׽�p<�!o�@>�b�h�W'^�!QD�r��	;g�����9D��1cmE�*&\xfC	��U���4D��0�C�_��,A�Ǩng�S�3D�@U.�ʰ�h���;uX��.;��xw�'���Vf��,ގ����	;E�I�'�����]54X��@�%34�[��C�+N�U@��'��e+�ϥ
Vnq E�E�M�>�j���\�>�$D��!���ħ�}v�9%���� gc8���\34Yj�K�2J���f���S�f,�'� �+P�xF�OQ>�cϔ19�x!�ֆ�L^v	r�H$D�hm'J7�P��ى!U�Em�����3Vʢ�K�3�ɘv�B��1(�9.�CQe۸$u@��D�u�Z��KUlV$��)G6���D�;�Zq���sT\Ѓb�.R�����ޥ�.4GR�ϋH�PK䣋z�S# �a���:k_HP{q
Ѷ/�C䉀i��P�UcՉ0`la����FH�˓T#Π�%mG#jӧ(��Y��	r@�� �膐)w"O �8�gL�/��hK�O�(qߎ]h0H�H�$�S����0��� (ښc��6U��l�r�٨px!��� *�^!���J�,;~�B/�q.���FU*���d��P���Um놴�G��<R�x�k�eV���<A�O:t�F����)g�0�Qu�GU�<�T)I�M0���RJ!;ڤH�⧆R�<i�	�YP!�#ef0�7�LS�<1G�<\B���RKP~84	�NPN�<��Q6�x�qd�r��� !F�<�1��R�dQ�1�H�=h4ᘱ�B�<�VO�w�V�@�B@=SÐ���a�<IE+��m�	���F�9��s��P�<�2h��	/���#;w(�3)Sp�<���]<!
�B�0U���+��s�<��O_�7'J}���.[�B]�K`�<A∅q�t���nҢA�Ċ��e�<����7iz�r4��4(�
��i�<�i��uI�p�e�m���j�<a��&b�� Kg.HVF\RA��N�<��#�q!���D�2f^�y�/E�<c`	);SNLxg&E�Mb:}�1i�|�<iU�S9"ijL�eǇE�Ĉh�O�<�Qd��(A! #B-`F���˜`�<��#����k��Q�a���v�<���-���͙bN^���IHn�<� �9�FøE�$��E�S�(<�""Oڭ�N��Pe��b��pR����"O�=a���X`)R���h�p�"O*Y�P�,�n���gI�i���;a"OZ��d@�7�H�{�%U�`��P"O�����٥NQ)�%S�9Z���"O<T�Ю3Z�t�Zq�ηA8K&�y�f �'�2'D�	��Rq䑋�yRj<v��Ud (
�����y&��I��y��8/�!��G��y���D9nx�`�(f�Uau���ygS����+4����q���y�	�}>��{�cK� ,�0���X��y�$�)�1��k���A����yBj<	Ș�8 �N�zo#�yr䇇Zބ��I��~��X��Տ�y�M�E���x��-]D����ė��y��y�F��#����H�	��Y��yb-ʘ�\��֙kA��	�3�y��`G� cĈ�8cF�C6)_�y�H���)��_�g��U9CD*�yBC�
`�2}��Qi�8KgE �y�D��"�����O�D�~��D��y�C�J.iP4�O9���0U��)�y���!����hͧI6����A���yBk�cSj|q�jK�7�} b��y��l��9%F7a��D��y���pT���E�t�c���y��'\�s��2ւA0��Ң�y�kƬn,�<ĪUf�tU�D��y�ĄFƮ�%�@�m�� �F�yc�	K���ׯN�V��l�&!ԡ�yR�LY��l��6W�z���mF��y� ZU��IU��M"� �e��ybOD�#z�<8�H�=?�V�xċ��yҏ���<
��ȗ\��(PC���yRK��\��Ћ�ƳW�ܰâ�U��y�`��*�X�!wf�X�3b����yZ�z�Z��$P<���+�e��\g��I�*M R�l�Ң.�[<���.W���F<\��a: 
g�8�ȓr�t�Av��y��+:�ه�~'hY�VIDu��AA��;/\��ȓL�.�;%J ?�q��|��]�ȓR�vtK���^��b� MW2��ȓ�AEDY�Ft)!U*͝#/�Մȓ,ƒ�r�H�Z�p��R 
�̆�3��;%��$ƀ���ĥ+iD���$n��;BB.�v��BJ�=�1���:+��uh�0��Ʈ>����ȓ&T	sF-���g�J(2�u��
{4<h�C����fQ�!��фȓo��PH7a��KHV�@��/)��!�ȓD��x!�Ďo~�x+W���4wZ����W=M~�5"OD�v�ۊ*o����W����G"O<�[� � ��ulϊ<���7"O�����5?/�+�99�1C!"O�t1�ů�=����$��q��"OX!W/ݙ;~��"��pZ"O�,X���v������-�TA�a"O�1�잪8�����
渹B"ODP�	O�*L�8��L�=�ұ�"Oժ�٬dӒ��j��.����c"O� Z!�R��n>5���UE�(�c�"O
<��ōP����􇙿0U��qf"O,�#��ԫ
B���I�6E%�w"OE��J%�vI���Аp<p�t"O�)�7Ć2�Qa2��/,��X;�"O6��q%�]���C�^�+����t"OPbr�J
t��8âT���� �"OH\�']-�0�!\7M�9!��'?x��͓uO�I�Y"({V�
)L�W�F:A�B�ɪ,�8a�Q�r< ���3hYlb���aE�j\f����S�j'^]�eeM����j̛n�rB�I&I+�� ��j����*���u�:�(H�.O�Ӗ
"�3}�M��K�H�����0^���sڠ��xRIĴ�R���ڸK�`P�䇂�>]LT�h��KF���d�'�,�㖎�5i�,�AL�?i�L�	�4l����M�9c�X��'�%iT)I="��BL�x��3	�'���*�A�a�S�#ܒu�B�(H>A��\�s�Z�HpoʭÈ�L�	H6	�T(*5�O82i.`X�"O0�b'J0,���5!�M�Z,hP��-pδ�r,��[���t�)��j� �nE����M޾ 	�Y��I�����O^�`���+?�A�o��J�����U�ȹ�R�7�Ҁ�di��B2J��$�Ϯ4�ą�.O�
q�L���O��#����z�p�I_�0�`$	:3r�g�2mD|q�$�Q ؕ"F۲g��Q[��D���?�1*�*,@:��dĐ_��H�a���|��R��ND��ȅr1�j�+/H.������t�W�[�N��55Ҹu,��z�s'�n�<ᦋ�>,0
�`��?�T�T��$o�D����шq`���a�@%H�.@�?(:� ��]?�@�,OZ��"�C�(�4�.+f�Iq�'`
��FK�m�L�Z��^�#�taV�z{ɐ���Ԙ�"��WF}�$ �؜�d�UP�'�F8;�]�c�vPs"�6�Vq��{Bb��W��LREbY8S��4C�S��Eө��sm�<6���w"цlV�5��4М�����7!���
��*֬D?"�ܐ���/�>X1��P�a�J�3b)mݍ0�&J)	VDPz�س�����VF�F}l����
�
vT��O�8&_�]����F� +l��2��NO������٩n\�R��+F�h�_�p��@U�5jT%��W��`���%xG�렣
�d
lҰ� �f��IdN(Jt���+8@Pf��5��8��! ��spCm�"	A+O���o�f����E�F:�H�
��W+���Eo�7��	*.@N���#��?aԤZ���
/F��dUJ��b�"B*�Z��$"D�n�0s|d�J�o(<�6��4�8��(߈<㦌k��eq�KA�6����mI0h�\�%?9����p~��{�rXhE�܋��%.���?�B��}�<P:ȁ�FЬ�c�7U�T9�cI�'0�0�č:;�D35�բ�0<i�޷\�J �blW @ZX�*U�'�x�{A䋲Xa�	+S΄:4-Z 6/\U���$]�� ���c_�J�O��y3u�ZxRw��.T �3R�0K�I\?5�L	�΋/t�a�����|
���<��|�tc�:��uVœN�<ӈڭ4���G�.@6A�![�4���sJz�~�䓵c��$?�R��u~�@���-*��̛CU�hc���x��@	I�(`��.>8�& M�Z����Č��aA���l�`���_y8�10�y@�G�f����6�H�y��xB��1K��zj�3$��M/l�Ԉ�ǼP�H��V��.7� ��v$�)_!�0^~�S��Ԟm��=�3��w±O�Ă����1F�P�O��Qy��d`{K"_;B��E�
�ތ3�"OARO ��㷩�<Z��SG�L!��qQ2��9{�0���h��W�q8lq7 ��G���yGd�a�!�$�^�� @W9k�9��C�#���
`��f���:>8��ɤ4[�b��W
>��c爠O	����:p��4@ѧ2Q�d[r�ɛ����$I��7�B$�fn���x�K��&�4�z��ׯY��Z�G��O ���g'GRA:��	o�g�H"'��wq�`u�� C�.l���Jq��A��Єˁ��x�C��PhH�q��)�)�矘�#ŇU:8]X�#]�����l;D�<��+q�n��ADH��423O6?����	0��a�@;�5P� 6 *d�F�Vx����_���� �GC�lh�ł8T��H�KBV�!�?_�j�@�	�?B62��;!�� >h����
y�(⮀�#�8�P�"O�Y�d��ҵ���L�l����1"O���p�.Sw�c�Jō Bj\+e"O��J�O����`7�H>l�\���"O8�`ՠ�l�ΙAI98�y"O�T��#Ǔ=��4#AIC������"O�%�Dd�3B*j���@(&�:���"O⡨�Dąo�}: �ϛݾ�{5"O��C0�E�HW����A�P�B���ƨa����	Ó^�<PELƽl���Hr`�.S����^�4 '�ӱY��9�a�V	Lu�@,ܸr�4����x�����@�F8he"Ѐe�J�D���d�U+���I�S�L	z�P��Q�:�@�fĭq�\B�,��a�cD�={�< (���.*!��ॣ ���e��ҧ(��YV
2x>�y
�2�U0�"O(�˶�ڧkT�#����8�d���-}�d�t{8��U�;��$\� �*� �@��7��C���⋜�%����B�e�D	9qiؤz�+T�Y�-s:8��ɾG�Z1�  4A%a�S�̢?y�@>4��$D5��ʹa � 3�U�f-����+X!�E;�T��.Z4bʌ����+,]剻jטyx���t��S�Oxh�1H�q�̩
�C�	;����'K����	e�:�2�N6:䀖d)}rj �bh�Q���{�d�c�~P)ǉ�p�ґ�P����x�$'a��9e��B��<S��&=̬1q��N�RG��G.l$�t&d�o�^�E��=�p<)��p��c�D�B�0jQ��X�֠IqRi���$D�0S	�n~L3ţ[$M_2Ms�,D�D ��$ j�B���
=�TH�A-D��J'K�3J�}��Ҩ;ܤtI�*=�oP��B��'���^�ʽܴ#����O�1 ���#��J��S��0��)������?�thO�&NZex�F I,��1+�i�'�,Y��� �$>U��V/z�MX�cA��� �Q
2D�|A��"��%��M�?
3j��TB�<��̊4 �<옵�2}��I˸d���sA^_�*�C��&Z�!�	,E�Y����Uݠ1e���p�b��O�U�JI���qOf����L[XIK"�I�_T� �f�'dl��hюlA�=ئ!��*���ełZTݘf$ZC؟\ c ^:j�D)�v �>8��Yx�&�y�Yreh[���]�4�^�\�,���R��Ic�"O�M�w*ѯ`T����t�N�;7_�X�"�8
����>E�DC�gۢ���I#k�)��Q��y'��av�8�O����`j�`ֿnr��' ���&�|��ϸ'�~�S�X�(�(���I�nj��	�'�z�3���PR���OW�ڪY#1��%o*x5�'��d�7	��g�����C�T$y	Ǔt�R���:��9�00����#�Y�Q�؅s�2B�I$W��E�u�)��Xe�)L�ZB��L|�%�3h�h���U�7�&B��͸ i�@.p3�@�۔P��Շ�n@�E���U�\N�0�KK�m��h�ȓ��d�b�V�
AHڗ��,)\�ԅȓBxdP���G�������z��ȓ� ���O�"���#0�[�J'<d�ȓII��r�À��q��/Rw�̄�dڌa���^t�2%�2;b���ȓ*`8�¢I̧um����<��(�ȓy�D�b �s��䒡iB�Z2q��+�zѩ&�!of� �V?air���[��L�$EC.p�� �!�>h
�$��Qhr5��E�(�d�c�#�\\�,�ȓ��V�E�������Ea���[]�e��J4/+�$�tj�U|:\��S�? �%�ӂ3(1�ىSGP�M��A"O,����]$2>=;�>\��+""O�1�뇴3(�P Sf��6<����"O���b��0:=����ft�{0"OH8��7ؚ�Y��g��@i�"O�d�m0���5��<��XC"O��mU	6Bq�Cd߲�"O�J����y�f�2�IW?`�\��&"O\�h#��$$�T�$J�*��D�"OD���nà���j�
PX�1�"Op=q��S��DU+�)��H#���"Ols��[�Q��l�Ub�V/�4�W�'u��R���(I��SU�Z Sߔ�s��Y�.~\d����53�`���'V��B���&̍�`��0No�Xd"Ox2�G�;7b���g�0H�Ti��"OD����	#��yxƄ]��,ɫ�"O�$�1��9�+Q��o��	�"Ò��&��eNX�T/�!`��J"O�0�QaD&~����^�#�0"O�mK%m�zd.R�4�����	=�HO��$�jJ�)]@��J��3��	�P�L�
m*1r�S�'���#7(��	�>RR&�Y�@�v�5z��`^��+5E]y��II�uMVI���ǴNc�`1R�٬Nn� S�Dդ^~H�'�8��� ��� QiX�6���+DD�1o�D	�윏��	�"�v�q��?�i�&i�-0qȒ@��|8�FL�1T4Tb�O� ��ƃ	6cx��
�'LM�"�U� ���3�Q�y�5�'�@ �P1��ȻN>������g��\ 
�1p�=�&o�I}�B�Pь��=E�$�ٔI��[᧓W�����%V;�y��Qz�����k +En5��'��:��S��6D�@Q�MB��p��l�9���'D���b`?M�$[E��7���3�$D��z�Η�Ń�ć����5F.D��C���$K:��6Ʉ*Q�,㑃-D�,��B
u��C� D�E<Ը!�+D��{�Wz.���m��9�s)D� ��]Y�N@{��[<��ܢЌ:D��8t��;����v�X�hk|�@	4D���V��)��1$�X�
G.�c��3D���2 &4N��4�,�$�&&D�4�ܮPHv�;i��v2���, D�@ㅚ�!����b�/� 5��<D��)�O/ ���G�}+J>D�@���'ܰ(�t$� g��3!/D� �"�Cy��:����j1iG�8D����+�d����)F�_�n(�B8D����{"�sD*C�Wn���B6D��	� S5S�*QZuk�x�zMh�4D�@q����S,�{�A�DR��0�H7D���f1�`1yӦ��wnt�9�*D��p'�4dҢ�IF��C#V��4�"D�ل��=L�֤��D;OW$1�1B;D�xzCb�6?�[�CiP�H��]�v�+D��h&�1��,a6�A$��2�*D��J֬�.q*���B�(7�`;�k<D�����{D%CvmT�,	�pc�'D��+�oCC1�mb��M0@���r�/D��A�ϖiEyӧ��	�hi���"D�dZ�`��zs(�j����N�;ь?D�\�C�4;E�1{n�IlިIRa>D��c�/E8�T����@�1�$R�� D��x�%O��y�Q J8�j@�d�<D��˥&�P�Y{@G�%��q"	?D�x���$<�L��7j�
���"D�ԲSDʡKR8�C�' =]1�@9�D?D�� �,�cIR'@ܸ'�_�;h0]�"O pD�87L)b&��)h�`��"O(@�f��Q�.9��� �cHfA��"O��t��h��xsm]�F��"OP�ڴ��+����,B��P#"O��hR���J)�İ#)!CR"On}�A��	\B`|(CH��T �$B�"Ol�cCa�c�6�.�R�"O�m+5`Ҙr2v�S��)t��2B"O<�+�L�"ר�*S-�� 邭��"O(��@@�.Ka0a!�,��E�nx�`"O�Id�A�!���d��,ժE�D"OV�ť�)4AN`���]��@t�""O�QukA�+�.��0���{�$]A2"O��%&�\��y� $�lI�"O� @�D �
0�շF�n��"O̚�Ojb�pѠ�9&t�h�v"Op����84��ҷ�*B[�9�"O�͠#�%~��)z�OK�Kq�{�"O���dW�^t��0�G�ϊ��b"O�h�@%-i�n����BQ���S"O��1�ܔF1�a�&�Ƣ43��!E"O�\�gC
NRh�
 �7#^�"O�t�G�7g�$b��<�"O-��]|	v Qf9<
\z7"Oze�aE-Z�DD�.R���%QK�<��f�1N^��8alѷl�2�PN�O�<AEO�+ʠTˠ`�FLn2Ӂd�<��j�,��iQ�ķO��Hy���\�<�4 U�JMQ���כ�]Z!�D�<#;T��I�H�l��J�T !�Ɋ=s�`P¢�#:$�yb���~!�d��G:H� Q	��G|�%XCaM$i�!���m�DbpU N$]���P�����A6o.J$�ǉ$�"�⬈�y����4�Х��	Q�E{e�)�yr(ĉx_�d�T��-O���o�y�a�4�!3 ��!�HZ�m�$�yB!�O��hA�.u�����X:�yB��7D���I�S�y�,��6��+�y���c��Y$�wt�!
�Py�ˋ>]hѸv�Y��X\`��Rp�<��ᅀ.��X���'|X�HVi�<�B��1H?�Qi$D�X���[tIJq�<�b��-~l՚���9z�Y��̑b�<Bn�J�C-�?�T��!�G�<a�j��رW�U�f����a�E�<�N�-X����b�Ab0��1-C�<Q�낂r�
A�a�^�(�J���c�<��V�%��q`%ǞsD�P0I�c�<��L�[]HsQ�"A�4���Le�<q�^�k���ɵ[7Z\ѫT��k�<a�P,/���2ȚwZ�-2��p�<�̢2 ��С�\ z�|9ƨ�h�<��@ߞi��km��=|�BG��d�<�d"��S�<[#b
��2��%d�a�<��'Q����Pj��ug����e[�<�E�<E���@�OO�>�m�T�<Y�-�'���z���u�R�[��YZ�<��T�����!n��\�X�R�V�<Q�I�7%�>@����'�|9�QR�<�ʒ�9�H�C��B$bh;Cv�<�&,��z���#��yZ���*�o�<���]1x��A!�Z�m�@c�[i�<� H��î�?f*.b���C�I�"O�q�T��5@ZVa v-D�+;�=R@"O`���W"?>�Q���݇L*��R"O����$x� !�ϖI"(�g"O�@sp)C !x�1!�7:v�|P�"O��#��DF�|Y�J�9AA>��'"O@x�G�W,�X��U(	�M+&T�R"O�:�/�K�6�Y�)�,���y�"O��dʹz0��H��o�� 0%"Ox��Q[x�|z1���h�z���"Ol�XO']��#�j�2���"O���Vg7t`����ڎN�
HA�"Ol݃�f<H���ZD�ɖ3����"O�|K�!,���61?�԰Y�"O��ã��y�h��&ުb�����"Op�r�Č12Eh��_�4�X{�"O~�B�k�w��p"�
��U��"O��͕1e���G��|�n��"O^�R�)�2a�0���1[D��"O!��kÞU��l	ƥ�|��v"O¤�SD؄/�:��7d�d�cG"O��Q�@O�q��!%y`�B�"OD�qr�٢]���H FXj	½��"O,�u���V@�S�M� ����"O��[�@A ]r�@�'�T�E"O �#�$0������,�PA��"O^�˒⃅"ul����]GF|yC"O��S�/ٙ]S���D�hV4!S�"OtD�6���jF�+zh"O�!䦙�yil���*��<���[Q"O�W�� =�(�F���`��5O�\�<q�J�Ȝ��
��7`H�"U�<�RoQ�^?�E��?x-�C�F�<iș�*햅�� ѕX�:�	%OP^�<Q����wy�k_�HCL���\p�<х�?aΕ�َ8���a�![n�<�ؕf��ya�E�|���$i�j�<�G� Exp����$3���_�<�"T1"_
	i�ȅ-2��n�Z�<�p/�v�#���9� ��J_n�<iV�^>=\H��K${ܚ0VO@l�<aը GvbY�V�ψ[b����R�<��D�F��`�_/��r��N�<�⌗l�R�����;��)�!B�<6a��4�< 'E��.�uk B�<!� �2Ԝ����6I�Q��"]@�<���:a�\HV��V�~�0���p�<g�Jhd�C�F�s��l��#Ul�<ɅH�)�R@���nխg�Yr�"O�V���0���MS�P�8(�"O��hc	�	fBB`'k�#p��j�"OB��'@�
{'����7����"Oi��D� _fda"`��#�\5ڤ"Ov�zf��H��	/�tt2�"OFT"�n�>?�8�2σ%w�p��v"OeA/�4����P��/�.�8%"OH��.U
�4htC��W�rmX"O�M�b^!Y�4�QC�	��a"Oh,@�f*y��M�S�ʩH��h"OX�������H�!��9��١"OH�3�ڧ�(�!k>3TDD��"O�!aG�X2,U<�0�I;IT�\
4"O�e�.A�!G"|;6�Т=~a�"O�t���:@c4��ף�m#N���"O� ڰ��Ȫ�,��֠8"�e��"OF�6�4W Z��d
C���"O���되=��Iʱb#x<��"OT��mEsI����k^!й@�"OJ�� h���� ��#=f	:�"Oly���O����1��7��p"O4�Ra�̩	�@��G��`�Y`�"O��R5d��>z�$�֮�6��d�G"O��AI�0`���s䋡S�B	��"ǑK%�@�A�ܜ����@�P�i "O��S�-H�n܀UO��6�����"O������LI�9���E}xx| 7"O���6D��DEd�΁�^���"O��%̉z�� ���^�\ &"O�-P@f�9.5ryȵ1QT$���"OT�P���,ܪ�`��a�rU"O�D�&�#�J�(����q�8�"O�� M��]��͢��G��~d:D"O�Q��TY(�Uӵ��_�"�Bc"O6,K+ې$��<���̭:���xw"Oj�h�

�Q׌X
��
;�����"O`=��S!��D�3���r&"O�9��*֭~��o� @c�`�q"O�a�UL�0�o�\q< :�"O�hsq(D�9;Xh�U��uYH��"O"���O\<-����D�Ԧ7=�]�r"O������#;�貁`�'hD�1K�"O���H\Lߎ����\"];!�"O��x��B�^���Q5���J.؍��"O����/D�IC��&$^�V"OL�	%	S	H�r	7���T�f-{�"OSWJ�~p9K׍	�d�֬JQ"O�  G���{�8�9�+A��` �"O5��LĞ�
0a�Kʝ^�p��3"O��͖�8��agJ��N��0"Of�!WG�Z�>}�hײ����"Od ).!W#�S!B��k�LmP0"Oj��ǊJ�K����@��O��Q�"O�����T5YN�`� #��y3�"O��dO�'䙐7��eH2]آ"Ov#��2{z��R�ͷ 88i��"O�L�`   ��   �  O  �  �  `*  �5  >A  �L  �X  �c  $o  �w  p~  &�  Ǝ  �  W�  ��  ܧ  /�  ��  �  k�  ��  y�  ��  &�  h�  ��  ��  }�  ]�  � � � � �!  * �1 "9 d? �E QI  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(��I|�O���#�H�R!��њ]��p��'_��uʆ�vӲ�R�c�*m�'�*L��܉�` ��ڭ\�����$֮w4I�1O�,��g�W�b-h4��Ӽ9�HMB�tX���;%�2���IЦ�Fx��2R^zmC`� �p��#�ȵ�yRO����!�L�q�tR� K��$"% �"|���6U3��B0)зez��%�~�<)0��.)�#U��4��뵥�T�<��۞@J9������
�ĥ�F�<���R�}��%�	2a ��`j�<�d��W��aP��ۆ&Z<�j�g���'o(�TA0g�]j�ȺS�����'���G U*=�~@�g��J��p`�'X���	B�z��X3'�R�m�4u�	�':��D�K���@ W/�S<������ �\q�C1������h=�A�#"O8��N� Gv����^�g �<#��>���tl@aM�/Dc��2X���ȓp_�B�"'���BQ �萄��N5[�œ�J�lU���V ��-D}�����Q��*�	��ȴ�� �C�I�qv�d��+̅Z�����슃'�B䉌�����"� TU��gɭ 6#>��C?�'w�6��![�.v���a(3�i��j�X��`	O̙K�aX���YΓ�hO?!F��*e�@y�FP�@�XɫA0D��:4��(N���q�S�/�����,D��z�K��U�TǄ�'TI�9�+$��g0��9�� �:�����o ����9P�M���4t\�\����ayR�O֒O�0���xb�Ӷ���V�{�"OQ4�B�|;z��&T���S�pG{��	�d�\@A �K���)��/�!��>P� L"��"GBi��&K/}�ttFz��9O�I��rL,y`��hX�xp��'��+K�Q�����T��������1��]m��<)�]~��ʆ�&O`�3�X'>��1��	k}�K>!B�;q@ηn��l����yRaA�90�����Zcz����Y���OL�~:��N�8aޜ�A($}�q��a�c�<��R;/xВ��E-�:ѡf�c�<Y�Y0�����j��u�C��i�<��#=uL-R��	�+($Q�E�]�<񳋟�%D��O�g��,P�I[�<��g�&�:�r&l��G�.a��&A@�<6��_N^�R��:���� �y�<�w�ґH�yz �3�`��� �j�<i7�}�2٣QO�p����2��q�<�5�̏�xq��T,�s�F�<�#��![����UN�t˞�b!W�<��k���≨��Q &Р��|�<�ƤS��ڑ�UF�JIj3�Mq�<���ߣ��� �M�1vN�Y©v�<�q#����g�)��!��v�<ag��R�F�� �>���Вd�V�<�����Ttހ	�[\��,3aL�i�<�a�C�2��-�I��T��x���F�<q3 �jT�㶦ւa�j0I�~�<a��WB�<�S�	?sC����j�o�<�"��P�:���=bJ��&��n�<�/�"��ړş6K2zD��c m�<�6�P�*���^�B�ވ��ŋ}�<I���1�0��#�3c�R͒��LS�<�$o�^ľQ�ԀR;1�:�Ns�<�d�)0��f�g�����/DG�<i���B���UB_�&���SFG�<i���b��C�Hܭc�����<�k��FWL�#�M�%j(X�FE�<�ä���8�d��&J ��DoV�<s�T�\���9�2M���Q�<��/	�P�RfD�<��l�F��e�<���G�#�H�1�K(v�d�4By�<qB�"J14Y��͏%�B���t�<�PHZ�:0v�a�U�E��!Y��p�<A&	�W�� ���~tb|��o�j�<Y@��.k�:��m�9pt
Q�5%f�<Q�4F�(�3�����k�'�F�<����r��t��v�J�{F�{�<!ݚa��	���.����d.�z�<� v�B_�0�q�� �f�2���"O�}p�4�V%Y7b��i�!("O(h�`�lB���5�B�	��""OJ5�f炖l��1��Åw ��Ҵ"O�IȒ��&$.i�Vo>)#�ı�'M2�'�B�']b�'V��'P��':L�Ye	�#?�T�*�j����ͻF�'���'���'N��'���'���'��q��(�.mZ���x��1r��'�R�'���'SR�'.��'���'�:�`I޽f��PmK;�8h�t�'�b�'�"�'?��'b�'���'���# ��4a�R�QB�Ɣ�f�'}��'���'q��'�r�'���'s.�[ukF<7aq����`%6���'���'2�'��'w��'/B�'��p�D܊o6~Z3�E$#d����'���'b�'-B�'��'�"�'�8}�#ެN:�J�MI�?	����'Q�'��'��'b��'7��'B���
I�s�t���ع5sx����'�B�'"�';��'/R�'�b�' ��J]�<�K��ӧc%tQq��'��'0�'�"�'*��'/�'�b,!a� YH�,ܲ4��>�?����?���?)��?����?���?���� #�d���B ;�
1�A��?���?i���?1��?y��?A���?�r+�
�\��,O=4���+� W�?Q��?���?����?9��k��V�'���Y�i�"qR�)�	�~��5ET�3����?�)O1��I��M#�O�(���h⦇Vvb�S�"��'��6�.�i>�	ݟ�P��f�~�d��Vp~�S�M�ڟ�	�a�zym�[~�<�:��S\�IDL��i��.�� Ƴ"��<�����/ڧ��sU�8!�0�밯��J][S�i���y������]
)����t��r5���Z22��������i�4Ҳ6-y����]�[�Rsd�(��v��̓5Fr�Rp�����'�N���W>hӚ����� SΤ�R�'��	g�,�M�K�N̓n��.-k�̺ �QI~��{�Mw��t�������	�<ѮO�x���[�"�Y�#�V,1,dhǒ���I=F� ���/�S�GҎOݟ��	¸� �J�/V8�SmxyT�<�)��<)�C�*����c��O���3�+�<��i-��1�O�Yl�G��|2�ꙷhHQ���N^���Q&��<���?Y��Sܞ ��4���`>���'煏�\�}�"�L�m[l0Bt���b]"�Of��|"��?y��?a�t
�2T/�D]�)�Ĝ;]���p-O�5lZ/u�����4��b�����$d�*PR�*"i�͹�*X9����ڦ�*����S�'U*��P�h%��N�B������x[���<)��*1���6���򤆱Z��rF5�����	FL�$�O����O^�4�0�Sg��*�7�
#�Fɑ���v~��-W<-Ab�v�����O��l��M+B�i�F���� ��h�An͸7��!�#�H?����L�F#,l�����$9!��ɭ+ ��$��YoN`8t5O����O��D�OP�d�Ot�?a����h�3�K&3���v/���@��d�ٴFk��.O2�m�t�Ie���H#��Ք����Ncs��YN<ᴽi=�7=�TP�u�4�3ʒ���	=2��x���N4E0pe���DR?��d�'����4�:���On���{�ƥ(�	QZ̈���兦y�@���O^��2�4R�7�'���'&��5d)̱d���WF�qY1C�)\d�$����M���i(O�3@(\X�-��&�����,&8!Ԋ��pn����l(?�':���dې��a�l��ӡ�.�r�P�&#�j����?���?��S�'��Q����ANW��p0�kb��ӣB9y�v���˟T��4��'J�2�b�Zܼ}Q���<;P��+�O�~��7���EqpN����'ܾ�Su���?駟��k�(QKnD�&&�}��Q��>O��?���?����?�����	A�Q�F8c2�P?Vu�b���$ �oھj��������B�������Ӳ	I�@���$�d4{�:m����a�4�&�b>%�t��Ʀ�Γ^)��	g���㉌./�(�l�Q a��O���J>1)O���O`����,	�ʜ�׉H�W���X���O�D�O���<&�i������'t��'���@Ř	
��)S�`�#R���'��_Y}�'M��|�j�jz�/hP�YRGQC.��#�OJ�.�ƌ	*�8��O�Ę�	:z��+\#Y�1p읊/��(���_��'�"�'}���	�V�%0�U*�ʅS-$d�U�؟��ش��]���?�c�i3�O��8"b�%�3S�%�F��W�+1��d�¦�ٴS�V�DQ`�&���Jפ��Vj�E�
9��1�F5	E��D.G4BP.�$������'�2�'���'��;QG)S�����+p0�R'^����4M6�Y����?I����<1chٯ>Y��p�CE�M�6h��<�����X�I7��S�']Ԃ��o	�<�(*A%��w=j@q���h����'�z���G�П,���|�W��ا)�2f\�H�G�5b@�*� _����I͟��I��zy��r�r䊓O�OB�⩌�H!�U�����a�O�TnZy��4���ß��	
�M�S-��W��)+��K0���Y4y�%3�4����J��\3����Op� ��QHV�(�8ĉ�'8R����9O`���O���O���O��?ɘ��ي�@���@��}d�5Ӣ#U̟���ٟ@Zݴj掠�)O�og�=�����ߊ��@(�"rm��eO/���5���|�d
���MC�O��!Fm��{4Ht�IR��#��52������v� ���<y.O�	�Oz���O~���gW@c��q
���t��O`�d�<q��i�"4�'G"�'�������1��.���yd�^���8K�I� �	���S����n�ja�rF ��:���E.V�P ��C\�L�:�O�	8�?�u��O��Ӓf��HЌ�����,}i�{�ͅ���������b>=�'��6݁xFr���,5Zɢ�s�`B�#��btD�O��D���]�?�^�����~蘉ȇ��>u�^%��`�
o����
�M�B�߲�M[�OR�V�:�*H?�0dFԽ^i2i�qӈBt��{�ؗ'"��'2�'br�'��S{�j���
��$:��bo��[���0�4
@�+���?	����Ou@7=��E��=WE�<:�G�&�4�� m�O���Nc�)��&'���l�<QÅ-x�|�AG�H!|���d��<��nʷ~�dG/����4�^���%����˼>���YG�����O��D�O��ac�6	\�L���'^��
K��j�,�qQ&�JQ� C��O���'E��'Y"OHIǎ��`e�X�@L��P�咟�����h!~p���/�i$��Oɟ�Y4��9�HTbA�ֻ���ȟ0����T�	џpE�D�'n�0@ʂ�b���E�%uL �P�'M6��C�����O�hn�R�Ӽk o��z�r3ρ2V'
�##�h?���M#U�i��{$�iC�ɩU�A�A�O~&h0b'� �$��e��g���A�G�F�	Wy�O,��'r��'4k׭s�l�9cc�9j�ve�F��%��	��M����?Q��?�I~�Fe�p@$õj�$����1X��$W�T�Iޟ��H<�|��V� o(E�&�8=֪-:���4�̜H�fS@~B�1-|���	� ��'}�?;Jh����/C.A
B�~���ԟp�I�d�i>Օ'�"6-�	u����3	���P�y05!�W�j���Ŧ	�?IP���	֟�j�4 <��g�n�B���k��/ �������M;�O��Ф�����$�w��=���C�j�����nǴ�rQy�'	��'��'��'��ء�.~|
ђ�b�.;�X+c��O��$�O�0nZ�E2N8�'�F7-.��H�?�d��F��(7V�o��N��&��#ڴa5��OL�}��i^�I�X��C�e�b�Yy#�K�x��Y�T�?fTb��U�Iy�O�2�'��gU[lr�H�կ|9I7 9ri�'�I�MKdOǭ�?)���?(�z���G�M�f`�3�Öj��Ý��x�OmZ��M#�xʟ��¤�\��uBB+�~���+5�Z/�>L��.W'.��i>���'H�a%��R`Q�]^X8Cb"Z9h�4��Z�p�I����Iԟb>�'�t6Mȿa��`j�"�\#�	�,Q�+���?���
����D�u}�t�J�[v�P�`�0�j�ı0��!Ū���1�ڴ7����4��$ѕ:��:����S�[8��Do��{J]H"kN�h/D��zyb�'I�'���'
T>UHWk�m��2a�ΦV����C�̗�M�vHT�?����?�H~��Xj��w�b8� ̌U�
����`Sj=�#af�։mZ���Ş��|2�t�;���m@qQM������P���hC�j��,TF��Ly�O��c��m_�qG���h���4�F�[ ��'��'�剉�M�4���?I��?�S�0"3\��q�ŤA{����	I!��'���?���Ez�'�I@��ەM�������>o�� �O"�1�!�F�KA�Ʉ�?1A��OLD:�ǌ�>f(��c!-$�^����O����O`���O~�}*��uV���Ūՙ��H�Ɉ%^)�t8�����M�	��	��M���wr��R��1���8A!_�f��R�'��'�7MC"j�6M7?���K9at����,�"a�C k-j��n�
PЩ�J>�.O�	�O����Ov���OB���+P��pˑ܀WFy�Dj�<A��i�pI� Z���IX�Ο �pHR5,Bp�C����e�h���B�����O��\�)�S�	=�e����<j�� �߄�T��V��j���$��O�ՒO>�,O�����ٮ\:�x��
2���K�
�O���O����O�)�<���i,n `��'dؗ�*Sx���GL�ܸ�YvF��?1B�i��O�L�'M��'a�@.|�B$�����0�H�&w�:8T�i���"q��u���O�q���+2�4����VV�X�����d�O��D�O����O��d5�ӵ0A�LI�c��K>�d���ےF�nQ��՟��	��M�-����$�M%��1�@�JsP�Cw ɡ75�)�Z�ēm�F�h����hϛ����1�KE�n��s�ڎm��D(�f'i�2��@�'٠�$�З��4�'�b�'�|�e��g��R�	��5>@1�'�"^�y�4,Q��:��?��������$"��H�L�v��FѹqD�����O�6��b�|���&.	�I8�#�6d(!�A�EL�8m��n�<�)��dD]؟S��|�璾C"p�2�
6*@ 1e �(M��'�R�'>���Q��8޴	��$���'��$A��W�9������?y�.ϛ��dvy�i�\��J.By��U�S��S��e�J�m�z8l�}~b
:Bm�z�� 0���"S��"�.��K�X�:�>OP��?����?����?�����	Ї,���� ��p���b��$̔=m��=x�,�	��x�	b�s�({������-v�5�a�A1�!h����?a��5���Ok�����i���G�/���4c�B2�X$@�D>�,i3ؒ�G6�O��|2�X���"��O�[,I�Ei�<a�� P���?i��?�/O� mZ&1�	���I�G���PC�=�B�!�%Z�Z��U�?q Z�hH�4j!b�x���5A���HWf].�pB�AB���$̺�=��%��@���)�������M�̚T�C��_�F�c�Z(5����O��D�O���*�'�?�IӀ91�m���#��0�*3�?��i�VUsD�'���p�r��]�b�\��IH�(�R�gڢ-X���	�M� �'����S�[b�柟�BTo�$/W���&%��t'���
"�֕m��$��'4�'���'l��'�`�:$��a��MC�N˅NMvy�0]��ݴ5HqJ��?����O<�6�'a���&��JƲ�BE �<y���?�N>%?��P��:sAL9��OO2���r��'yu��2�ĞQybOȻv����I{�'��	 }.��ʦ�N
/Ҽ���+.E�T�'�'��O����M��*�?y�gN�7y@Ձ��2`�|�� �?��iY�O���'`�7�������4D���:�	��W\��A/�K�Ę�#X8�M�O$qX�������w���3�\*i,`�yVi��&@���'b�'���'�RQ�b>Z��B w��SCM�0���:dE� �	��`�ٴE<V��O��6M:��*&�*!����\�.m �t}����xr�'e�O���i��	%UH�!ae�0�Xq����߆���Q���P�IXy�O���'z"�*N2��0�H��a��Ȳ��U�T���'��I�M۵�Z'���Oʧ[��E1�/
�kMdX"MgQ^��'ȴ��?�4G�ɧ�)�z 8-x㨝,q��J� Tcfdq H��\�jǕ��ӕ"��v�	�D^�q1�Z{��!�?Np��Iџ�������)�Sgy""{��X����&:,��_�{V)@�����vқ��d^q}�'�� ��"�M-��'��J9�'$�6��1T��7m.?9Fئax��-���V-'����S&yP9PǭӅ�y�X�4�	����I�\�Iȟ��O{6<jW@�N�;R�Dq�@Xci�zի�#�O����O�������ͦ�ݺC��(�&Ѩy�AT�7,��ៜ&�b>9j�.�զy͓bL@�ToT�Nb��.\�H��̓@��ux$��O�u�L>I,O�	�O��#����1�2Щ|xV����OP�D�OZ�$�<ǳi6y���'�B�'���葭
�}�d��aU1'!��;t��GQ}��'i��|r�ޖWT԰��W�"�ʕ��4��D���XqA�ïlj1�8\Y��ij��Dٞo3,H����pXT��;����Ob���OP�$>ڧ�?q#d�($�|c�g�'	�¡&B0�?�@�iTt���'9�j�4���h�� ���m( ���J��9�M��ii�7�@*Ү6!?i�9��I�D̂��E#�6�*`1��T+d�Y���<ͧ�?����?���?�F�)&�]��߶ol��
���ʦ{��L���	П�$?��I�M�"�@��/������3D2�`�O��$�O\�%�b>u���(K�A�b뇻.������:[&�B�5?���}�>�d	�����E*	qDt`ta�;>��4�Eʗ7]v�$�O,���O&�4�l�]�6��./��Y�D�$R���(mBb���i)=l�p�6����OD�lھ�MC�i�\)0�P5�Z�㧌*G��=�3.��Z�敟��7#�W������x��tE�
�t 2�� l��
�4OV���On�$�O����O��?�#��<���9�i��>r`���������ڟ<j�4^Ũy@/O��la�	#`�b=R!�)F�|0teԸH�N<����?�'_�,�rߴ���0}����'J*A�a+w��x�jAx�.��?��8��<ͧ�?i���?�D�K�_lF�oڣ!~|�CuQ6�?����D�������dy��'��ӥL6�P��5T$�}˃��!()��d�����\�	@�)�W�� WZPXQ�Y.R�(�	���z�r�C0�����ġGǟ4KW�|2C]N����5� #Y�I`s#����'�"�'���\����4`�ҥZ�#��Fw^Pb�]��5����?a������z}��'!��F�F*Ϧ=XK��%<V�q�'@���Ŀi���Y�l���Od�_�|��C�5Ґ%DM�#;�<̓��d�O����O��d�Of�ĩ|:��ev�TWiNV$�Ҥ{��-T5
�����%?u�I?�M�;F�舚�L*?.���#[�tБ`���?�J>�|z���&�M��'����+�=u�, ��Jױ_n���'��R��Bß4�U�|�[��S��|#�O�ZZE��,8�n�j l���8�Iܟ��	ayB�|�"4pd�O�d�OH�*���n ɺ5�Y�r�v���%�	)����O�d9��ͅY+����	H`���©X��2C����@�S�b>����'���	�'pzlj0&A-:���v���;�D�������ߟ��	T�OM=x_z���4[��ɹ�H�4}*�m���u��O��GܦU�?ͻF,�Z��
]
p�q���)-����?�ڴ��vc�p枟Ш��đG�4�7� �p�5FڷJ�n}1ǅ��H@��Z�)�$�<�'�?���?i���?y �L&C�D����F��t$U+��$����``O���I��'?���*9UrMy�L�x�NK1@�%�`�*+O��d�O��O�O�VB�Y�G�@����ØzJ\cs��6�y��_��)��(��[m�gy��3�t�B���; d��"�Z�*�r�'���'�O��I�?A����,�Vl�;D�6Ha·c7�8+-����ܴ��'�˓�?1�4AЛ�ŧh��{�l�*��`��fޭ"q:U ��i�I�y��cQ�O�q���.�>��ш��_]=��c��,��O��D�O*���O��;�S�vNtx��ʔ�tp���D ʡ�i�'2��yӾ5���?���4��5;t�ɦLޓu�f�Bsd�x{�1��|R�'y��O7�(Y�i��ɛ��\�b%�$�H��EgT1O�x���/\�D~�Sy�O�R�'W����c��!��?F�J�A	;R�'2�7�M�%臱�?����?�,�$3p��{�BJA1"05�4��@b�O��D�OT�O�142��Tֿ7�p�H��A:H�C#&ȿ~-8�z�-?ͧw�P�����Y�*91�-�mĮX�v��8>|�����?����?1�S�'���Q:�&f�ƌ�P��M(ر�e��!Vnh��؟<aܴ��'P6�A����V�[Aˋ2bN�Ԋf����6-����ƝƦ�'TY���?���F1�!����5�ƌ ,�����0O@ʓ�?q���?����?����	�Ȱ���!V�aU��:v�Po�?�����˟���Q�s������{FFך%�����ƅ?5���S ޡwg����O�O1�ZY1'�eӮ�	�
V(\���Ʒ!¡0ĉ�
����ul C��'��'��'���'nD��rK0{'�M��B��@ZS�'��'�2Y��@�4($�����?I�����#����i1 ���R�$J��k�>����?H>1�
�E��B��#Q����jK~B�F�5ٶ��7�U��Oδ���
>����[��H��(�Z���C��E�B�'���'�S��ST�ќC? X����>F6q� ���̸�4# h1�+O�unZN�ӼÅǟ"$�)��q����A��<!���?Q��i6����in�I�t�5�P�O�|lDoէ+�8$ �E��|�4̊f�Fy�O���'["�'�2'ʆYBTP�!D��h����)��^�	�MC������$�O��?)R��J��ʎ
(�|��@����Ц�a���Şg�H���� E���(���!���  ��t�rM.O��K��A��?�5e1�D�<Q�b�'NX�Kդ!Ф	h])J�d�O��D�O�4���$��v ��%N�.��t���ʌv�2ŋpGñol�l�6� ��O�ln�=�?��4x�}�G-�Ƥ����<�@���J�M+�OL�B#���Q�)����Dq�E�M�t�T8�Q߀�Z��3O��D�O����O���O
�?�B*��b��,	u��+��!�$IE���	П���4P���'�?�b�i��'�Ơ�A�.��<punݐb:�)�5(,��X���޴�z4Bˌ�M�'rh��p[Ƀ,/gj!�4��蜵�%	������|BY������,�	��P��lQi䞈۶^nV�I�!������py��m��J�h�O��$�O �'8h}��Z�S� ���N-`.���'����?����S���	I��]d��%��%o'y���A�x�|�8�O�)���?�q�$��c�3���*���BӺ_�n�D�O��d�Ot��<F�i΢�Ղȁv+��� 	�����Ð1_/��'�6-?�������O|űC`�ަUc�@���E@ ��O���E"�6??��@��c���)$�/J%t}tq�
��)�:�{3G��y�W�H�	۟��	ٟ��I㟼�O.T�� L��;� ���ղ�!�:2����;��'"����'6=�52���J����a�#~7�B6��O��D0���	vA�7mv����n�z�0�� ���5���f�t���W�#��Ic��Oy�OgRʁ�W�Db5bI3}|Q��E�@���'8"�'B�	=�M�É�>�?	��?�!��A���J����b��b"����'S���?I����+p.X��Β4��q��k�Ф�'jH�#ΰ!�0�ɏ�T%���g�'��h�l�6"��{ ����;R�'���'���'��>��	��-��(����āS��|�����M�iL��?���;��4�&�3GT�H=�%����]��b�3O����O�Uo�n�*0oZH~B�Z�{�F��S�8I���7���;�z9!&B�u�Za��|V�������֟���ܟ웅"ϪT�`9��H��6���rqH�pyB�h�DkD.�O����O����B�/��8�bH߂,�� ���?8h�':R�'��O1���M�?�B�&�Ӯ���rK� n�D@�#��D9��: ��GH�{yB�
�WC��9�Bĝ6�A$\(uR�'2�'��Oe�I�M�q�:�?!qF��Z���� )u|�����?aдi��O&h�'J�'!�㞧
��#�%�I_�d�	@���x�i��I' m����O�q�x��H�Q�=sBK�d��a�GfĘ���OZ���O8���O��$*�3c�|h	W�	�L��Y*���&Ae�=�	֟0����?�&#z>e���M�N>��$�{�pI�7���0/��AX3jL�'AZ6��Ʀ�S~�qn�z~��I� �(�"m
-~�lbUK,ά�BV��#�?q��(��<�'�?����?�F)ɒ-+ #r0VtvMٲ�*�?)����$���C�A�Yy�'Y�ӣ	C�`U��5�N���DN� |�	/�M{�i\O��F���dF��K�]�!ŏ1o�Jei�f���$�4a6?ͧ����,��K�*�Y��[:MA�'�8�
�����?���?��Ş����eI*�+X~�e�_hh���=Π��g	ky��y���XҮO�oډ�zqI�	.o�H!A�"ez��4*K��cK%6�֒�DYB�],e��~�pk !-���UJK�Y
�0�Œ�<*Od���O����O����OR˧_-pX��M�,���U�6���׷i����'��'��O�2�a��W,I���Ǿ���B�M�mOx�m��M���x��I�R	��1O�	 �Þr�p���o�S�`�1�3O6�2
�.�?��)6�$�<�'�?�$�E,u����t��x�`�a����?)��?�������ћ��]��|�I�IU#�j�t�dhP
R�(:�`VR��r�O���OB�&�ĺ�G�.m���r�'���9S�>?���E&!|Hq�i̧#v���)�?�FE�YnL��N P�� ��Ï��?	���?����?�����O��z��#�f�Eƙ�*�|��C�O.�mڛ��4��ϟݴ���yG*J�/��xr���+�l�f@��yB�'��fӨMˀex��|4�a��h���}A�L9qH �%�
X��zc������4�����O6���OD���9�\9HCiVsY❻��5,&
˓|)�V�ޞT�B�'�R���'�r	#q@Z�.�>�ҬӌUIpٙ�˵>)���?	��x��d����XȺv錢���̎P�]�́#�����3 J�Od�L>(O������>�n%�tDO�o��L����OZ�d�O����O�i�<y�i��rp�'@�-��1(���{��yw8�1�'8�7m3��	�����������M�4o�}����B`�HȈ93���
VR��4��D��r*�c��c�.��$�����$i��'ƫ8���"�&F��d�O����O*�$�O���$�S�$���Ss��:-kP@sc��:;�L��	����	'�M�"k��|���zM���|"/�)BXՈg��tæ%�1IW�S��O�Hoڌ�M�'D�L�cٴ���^0�ZT
b!�!� ����]\�R���?��( �d�<ͧ�?���?�ÌR�vT���/� �0����?����ঝC ��$��ԟ<�OG��jS!6�Ȍ�­�(3l�O��'��6�⦩�L<�O?���e��"�
(C�F�T�鰵�\u`�sb��7��4��Ģ�e�ԒObA�S�%3�T���"X������K�O��$�O���O1� ˓} �V$A*Z��qq%� ���;�@Ni�=�%�'sb.}����O�,o�,Yb0IV�#mNjM���� #�d���4$ț��\�f?�V��0A�
Q�mF���~r�IP9���!R,åz���A���<�+O����O*���O��$�Of˧��R0���]Ere�ǔq9J"�i����'���'�O��Ob��׃;��P�C���TC�Mw�� ���D�O�'�b>U�
ϦE�|y�1@s�ؙuR����74 ��͓5w8����O"pKK>�/O�)�O���tϘI��3�AˮX��lB�)�O����O��Ġ<ie�i�Zʐ�'��'D .�>c�8闤�2C�"x����A}�'�Ҕ|�㉵�\����|e�U:�.ۿ��d^3}� -�GP�z1�)���p��,F`
h����s�(4S���G�Ot���OV���O �}R����a)S�!#?�T��֑z�٩����fC�j���'&.7�%�i��맏��ti	�L��Q|z ������4#��-t�f��F�r�h�o������ܑ�p�ߐ��ԠA�0u]2�p�HѰ����4�4���O����Oz����B��rf�o��I��  3�ʓ<c���Q�B�'-r��T�'���r���5%�p�`}i��<���Mc'�|J~*����Goj�Q�̐�/��eJ�
B&�j�&O~�;�*d�I-+�'��	$�!B(T�%P�y���%?A8Y�	柼��џ��i>��'��d��Ns�덥m�ِ�F��F�����N���yr-r��⟖ay2�'��&�m���qb��#j1�8�'�OqXUhdl��
y�6-,?IU!��<{��	8�S�ߝH�����2`S�C�TY�es�,��ޟ���џ��I֟���Fރr)�D�U�z�~�2FLP��?���?�ջiC!S��pܴ��j*�� ��O�zG,�.���醒x��'^�ON��־i���5����	)��
�ύ;?>��'$P� ��i��|y�O�2�'�"�O#a�����M��2�`@Q�	�)b�'��I4�M;���0�?���?�,��0�
�<$B�*Q�1���O0�d�O��O��'�rm��͈�<�LA���_�l���q�)W�f-~$���>?ͧw�P������,��գD$FI���;;i�hq��?���?Q�Ş���JЦU�5K��b���`��vϠ!i��I�02v���ߟ���4��'<���?��˩�x�y"��(Hc���v�HH��ȟd������'!�a�e\�?��:�"�c/q8�PZ�)>5���G1O:��?���?���?)���򉀼l�`5�.��X�6Q�T,F&vf��n>m��-�	����A�S柸p����%�%1�H�`�;:F���E�?Q���S�'	i$
�4�y
� JT����\V}ԭ_>lW�4"�3O��AgE���?�vE(��<�'�?���QԒ �F�+[����iS�?I���?�����d��ғ�U�x����g�M%ǖMRE��/oX,$8���s�p�I��M���'܉'E��P�).3��QI$��<Њ���OP��T�(L酠!��8�?����OL=��I�*y�h�a�N�0WLdY�N�O*��O��D�O£}
��!��IP�ڱ_�̵doR=��LC��"�6�Wv���'l6m(�iށ��SQ�舋��<��#��w���4���i0t�i���=�ʩt�O&0�"�I�Q��`��I��Ѹ��Ty��KyB�'��'��'��ӳ
��PSH[�;��M�S�HI���2�M;P��?����?1L~��N�ڭ�S�ۺ�9'���L ��TY�\�޴�"�x���*�lm �J��Q1�A���>1�̘P��J��	3ds���'(�&��'sz%�.ݗ.�2X�pǛ[;����'�R�'Ib���]�p�4W$؁��SQu�C�^�٢�v�Ǭl�͓5Û���uyR�'��jj��F2�0r��Ȃ|���#�B�f5�6+?&B�M >��'���0AO���8��I�4�{t�c�$�	̟ �I����ݟ��R5(O *�\#hJ�\��hZa���?���?�7�i��;�Z�l�ܴ��b��A�Jրr�Tx��]�'ЈbF�|��'%��O_4��i�I0K~ � �NL
pVI�D+L�($�_ �"��D��Oy�Od��'"�� 'V2H#q���$u����3g��'N�ɀ�M����?i���?)*���a�<��H�Bf�,1JFY[���D)�OFPoڿ�M3'�xʟ�X�5�*6x���T;R@�ip����Qb�X�GN�i>�Y�'���&��� Iêqad��r��1;��4�'AV蟨�Iɟ�	�b>�'��6�X�����.]6 =,�0E\&(����`)�O����䦭�?�TX�|�4Q}�8J�ȝ_J����Z�_�Č��im7-_�^ 7�'?I�H�PZ�	8�$!B<tC�!a��2���	A��yrT�H���L�	ޟL�I�p�O+�l�u!I-,)ꍡ5D�6�l�g�n)��e�O��$�OD����D�Ԧ�]?C�	�BC�Q�r�`Af*$s�u9�4QW�I4��q��7Ms����U�f���W���� w�@P�f�#"ɏM�	my�O,�GI8�x��D�(?<a�Ff?��'���'��	8�M+6n���d�OBm91�V/j4ܩx�&.�|�� B5�I����惡Y�4l��'9v��ק�'|�a�W�x����O�#���c�j�����?�O�uؠ�Ö`h8���!u=�"T��OB���O����O��}���E����_A��!&��acl�������.-pR �s��OP��R���?�;w;����QN�@\Y�Y|ʌΓ*o��/u��m�k@En�O~���  ����'7�ZAv � �8�0���5S��|rZ��џ,��������0�T�C�W��VO_0sP���Q"�\y2rӢ���-�O��$�OJ����S�0'�M��c��-�:e�c-�.���'{7�֦5I<�|��eΐ2��=a�f߯g�D�N]�_��9)��G~"-��\��m�	���'���$U��� �b �5�\	ز��|��L�IП��Пp�i>�'6�TY\"���' ��ȩ���:7���«��R����L٦��?�#W���	����ܴ}z��[&�_0n���I�%O`T�%�?�M+�O�<aT���B����@*B������"w�y��o�,`u�5/L8r��qҗÝ|�n�a��W�BǪT�v�,k-��agm�8HVՋ�*G.^��h��˖<c�4%�5�ɲKd!�5K�8#� �G�D����%Yx�	ɣHR��u�6�֧llJ]�@	��2�Ř1�S��6�j�%Ҋ�hL�"JW��d�Y��ѭxD���Ŀά��"�K ![ٸ��Z]n�ڃ���&��T��d��m�m �f�#$2ˣ�N.=c~9xf�Nu>a���*
��$��a68�(K�1d��@b����)�	֟��^���'\�S͟���xƴ�r��Әe;0`ߜS@�p�󄊨J.�'>m�	Ɵ��ɖXj�(6��Щ��>�l��6!�{y������<I����cy69��ȴZ���K�g&x�@��c]�`դ��@����?a��?���?gJ�'w2<D $���x��3�fS�vy����?(O���=���O��d��m�³��5�8�C�B�@��� R�C������������џ`�m�H����_`��.�	+��H�q�'|��'̓0N��(�4_V��`����-h�c�-RW6��'}��'|�Q�TȲ&����O��u'(�Lg\�uh��:�b�ꦁ��]����D��=���[�2`����F��,
C�˦%�	D�'b���Wå~���?���~-D�A��;]y���U �:~�EB7�x"�'t�J���O���5F�x� )u��3dEe9�7�<�)ԡPa���'C��'���F�>��(���摆F,^�sg/;hV m��8�ɧ8�&��	�[���ָOwT}�(
�b�U���ͽN�PL�ٴ��A9A�i�2�'���O�.����M�_"�!��R�! ��EQU]J@nZ9wZ"<��T�'7��g��:he���S;2�.� �K{���d�O��dH=7E�d�'��X�DҸV�m��*�[8%��5�*z�D��F����wh�t�Op��'�Zc�V��*۳6X!��<��A޴�?���J+ =�Ieyb�'#ɧ5�h�>�`hXa�TBR�Jv������'w�l�O����OP���<��� �Y�d��?
�69��bϘm��	B���*���Ty��'w�'���'��iV���f�*m�᭞2=$�a�0x��F9�y��'\��'k�	x�z8��O�f�zE%�9`)B]چ�1F���ش����OʓO����OҨZg뵟�k��ۣE�@�cόIc��h%��>���?����򤃈 {��O��ۨ6�\-�Ƣ��0V �P�G.�6��O�O^���OA����O5��]�L��X�d�֘�B��;v�`S��gӨ�D�O
ʓ3]�uI`\?�I���S�bDɘ�bl��J�O�R�&� J<����?���U;��'2����:��2L�p��X ��%j+�VR�$"��Z��MC���?����j P��X7f�d%9�`�8.:!�7a�i 7�O��3�"�<�}��$��d�4̲5jG�H�ڸ����ߦE���0�Ms���?����B0[���'H�Ђˑ�2��)w�o�����<(���O0�������W��|J2�[!y���b�F�W��iub�'_2��
q]:���D�O��ɼkܰ�{��A	od��N1_c�|R�KV��ן��Iޟt��"%��� /�3H����j���MK��7zFa:0Y�|�'�BR�x�i�-��%Z&Y&����E�м�F-�>�dK��䓭?����?�-O�$1�m]oT�,�AN�0���W�����%���	ӟ $����u'A��oB�|ʷϝ#5�d](�L���M����O���Of˓���b1�԰a�S������~� c�Z�h�����$�l���$�'A Y.m~�(Q�M����j4E����	ɟ���@�'=Z�`��?�I?��qSvg�3�t3����K��m��@$�D�����'��%��%��S`5�a��iY�oZݟp�	`y"��c�����D�k�]�8�u�V�I��2 ���mƉ'�I��t�I~�s�֝�)�@ݒ�mQ6:pk��ĭsJ��?B
�?��?����(O�.ӥp�Ib�� 3n\�p�?!��'M�I4w? "<%>Q�����r�0K ���`�~b��O�D�O������S���^���$�@lU�P;�ۍ_� �^���Dx��	��H6�eXF�<�DYG��eIڽo����럜Iw		{yʟL�'-��� � `�Z���XpV*x� �1Pᱟ:�䲟@h��X6!��P���۪0i�E!��xӦ��3$ِ˓���o��$İ�&� ?,�P����E�xR�ƍҘ'��T���I�%��X��Q>3�F(��d��wXhxG��ey�'���D�O��I�l�J��4h��$���;>O7M��
m�I��	ǟ�'�Z��sJp>K�>���X�5�ܬ�'mȓqs��֟��I|��Vy�O���#!�n�7��<�H��LD}���?���?/O6QʕC�i�S�[	t�i�5���{�A�?�F��4�?������ON�'�?�J?!(�+�Y�v`j����L �\��j��d�<	�M��-���$�O���(Z�!WC��� ���m� t���x�'�B� �H���y��(��$M@�\pk�A8Sz�K�i���%$F��ڴA�ʟ<�S���Jt�1H��!���C��N��VY��b������O|�I~n�=M�P�ǏH<j,����0zH�6M�,d���$�Ol���OT�I�<�O�$P�ǜ�f0�ӁCV��L# d�5ɂa�9�1O?A1珖&+��2�A�\
�������Ms���D��h/j�S�4�>!פT�L���d��t��Uz��ɩ�1O��{)V�Sʟ������*!�i D��%��X�����H�+�Ms��d
"`� �x�O�R�|�fe���b!*�1,(�
ĥ� |9��V�a�����?�*Op���\\}.
�Ճ��\j	�e��.������e��?����@)`�c�$`/p��E&��6z�A�4-�	���'W��'+�?�i�|� ��?u��0� ʔ%htu�@l��]�'1�Z�X������	��u�|�V��.ꀀp��Q�#�R�*2����M�s�n���?Y*O���%�Q�4��5I��;t�Yc���z�CPʟ��M�����d�O>�D�O*�:';O�����@p3�6\��`!d�7 �H�"�j�l�D�O�ʓXe,���W?-���$�Ӡ?jn��tHH	M/~�+��4�ڑ�OH�d�O��%M0�<a�͈�������Oq0�i'?�|�ـ����M�.Oz8��Ʀ����t�I�?a٨O���H�*�R��o�p�`�5���'B򪞘�y��'��	wܧY��8�$C+i�R�5D�?M	P4nګ��Hs�4�?���?��'���Zyb�.x�$�0sc�-�ڥ�Э/��6�8z\�1��8�����d��o���"�ʳ`�䡂d��M���?q��h��5_�ܖ'x�O�A�!�N�`�n�����w�4��\� �'Ŕ���O���O����Ot���-!�Щ�Ɗ�+�H��Q�릑��."�޸*�O���?�-O���Ɛ��f�H�5�VU#����#f>�R T� ��x�����I˟���Py�M[/}R�y{��_16��YS/�C�J�اj�>�-O��$�<���?���q}@40qFg^��!�_"SG��Y "�<1���?�됡�?9����$�@�ƍ�'k�99���RڰM�w�U( �"$lsy��'��I��	�L�mp�8sB�)�F\�%��R`��h���0�M3��?Y��?.O���ςi���'�� N,3�KH�2"��Ȱo�6a��أ�i'bW��I����	�k���Iq�dJ�8��ըT��r׀ !���0q��F�'�B^��T�O&����O��d����z�m�_m qkf˵~��EO�i}�'Y��'��58�'��	�>G��':���굀Y� 0Z�
u̟2e�inXy� �)cB�7��O����O��I�r}ZwF�1�G�i�j�n�i d�hߴ�?)��>@͓�?y.On�>u8
�	S��!��ڢ>(�@��|�`Q������ǟ8�I�?Y��O,�L�@�v)�Dq*$jH�KUp�0��i ���O,���O?r���Q��N�|�,	��N@��l7-�O���:�FA�ej����O���f��+WF�A�Δ�b� L07�#����^o�?��	ԟ$�''IV�XƁJ854<�'�Ήn\�Ln�ʟ��N�8��$�<������Ok��).�j��J\57��CM�:���<&|������I֟���˟��'v���	5,p�0��,D*�#��	zt�O���OʒO���O��un����@��	���!U���<	���?������ Eb<�'bX^�a���@����8m��\�'��'?�'��'���%�'�x�)���Z�Jl���#32��6�>����?9���DH�l&>5A�F�Mt����(��K�����
�MK�����?A��_��͓��:Rj���Wu��؂u�P�oy�6��O`�ĺ<!�]6�OS��OBj�c3G����LA4K�Z�!��(�D�O��d)%p�$8��?�w�=,f
��cJ/�f!�׉fӬʓ6.�|��i�h꧳?���c��I�bY�㵀͕|����� &�B6�O�$�'\����8��=�Se=��K7E/Kx)"��$�.6L,Y�*�lџ�I�`�S;�ē�?��̙a���� )�O�r�!�&���lݎn|����O.�Q�O=Y�(�#! (�I�!���	�I� �I�i6d��}��'H�Ė�I`Jl�q��F��=����(�|Rb��y"Y� �� �i�5���[�xS\�@�é_`�`*�yӼ�d�43idm�>Q�����+�&�(C�D�s���qIF�n�g}��I�yZ���Iܟ��	hy�ۦ<Z`����^�.;��f	/Q��@�#j6��O��d6���O��d]2}��E閼7�|�Ӈg�BL���s
=���O��d�Ol˓]?�5y�:�zA�EN�~Y�[���"z1"��x��'T�'���'ՔQW�'m�HjĪ�5jT<5`�ЬI.��&�>���?q���к,�L&>�jE�
Fc�0C*я9�8P���S��M[�����?Q�?�ؼ�����IH��)	���q�Ұ��lާHF6-�O����<�d%K$8��O���O��顁	�6m��9�/;m�	�!I0��O���δJ��5�d�?�{�jD�J[����/�:j�>|3 "s�Z�|~U���i2맯?��'e�	8F:Y�Wϗ��L�i�$�/4 7��O��L*=�D&��0�S�u���4mA{e�h��6�ʤw�(�oZȟ@��⟐����'��i�0 \0p�a��I�J>�3UIk�Y3�1O:�O�?I�I�pj$����C��c�5YT�)rڴ�?���y��<9M�On�d����
�� `��r�	X���t�h�Z�O\�!1�Q�矼��韼&a�{P��C熣fE:�IK.�M[�'�ذ�x��'r�|Zc�xԻP�S.\\&�I�4�x�OP,qV5O���?�����Jڸ� ��ߢ-[pz��ʨ~q�10��TڱO��$!���O�����aX�2�!0}�\��R�� *T2�դ�O�˓�?)���?�.O(9{Q%��|b�/�c���02�E!,]0�jBi}"�'L��|2�'M2�&�y>\2��Po@(����!��%3L��?���?�)O���� �]� ]�5���y�TP���A�E���4�hO��dV:fv��+}�o�D�a��HN"6ġ)܊[�'`�X�x�\e|D������k��Q�8 �ά1�Z=��E�e*�O���!A���'�T?AC��b6�c�#�>d6�y�3�f��˓
WD%��i�l�'�?i�'���Kdp�d��p=�4���KO2��?�l$�?AH>�~���ޚd^1�$EB��T�Qł��y:	B����ߟL��?��	͟�O�֤B��E��p��D_�_�	��{ӂ тmJ�11O>��Iil��c&�:}4��I��-��ز�4�?����?a�?���z���']rC�+np���ݽf%��s��7y�c�0�bd=�	˟h����T�1iB�Yz��d$�,�ʜ��,\����4*b�'��Iȟ�$�Л�e��$��qj�a�:C����-58� ��\��Ο,�Iqyb+��J�ܜ�V�z�Tp�D̠P�񠤤�>/O�$�<���?�~E�83D郪S�Nxr�wG��{Ć7������I����'v���w�m>m{� 	b0������:`h�.l�ʓ�?i(O�$�O����� ,�Ĩ���Z�hW�0�7LH?e��l؟���ԟT��SyB�+���'�?	�n�6
�B�!�T$2]�l &\�V�'/�I��	ݟ��0�y��O� ��Tҵ��;B������M����?1(O�`��D���'�b�O�"  # �-(M1��OA���ŧ>!��?�\J(<�����?����^	�2���J�8n-��hiӘ˓0g^��F�i�B�'���O#n�Ӻ� hT�VGK�4	��AH(X�\0� �i�r�'�� ڞ'�]���}��E �0�3�J�(�bp���Ϧ�"a@��M���?����_�Ĕ'*(� ���cy�@	]6���baj�6HK�;O.���<�����'�`Qq♡#}�̋5�%Z�%��/g�����O��D9dv
��'}��֟X�(U� 0!��j^�t�G�rDn�ӟ��'ڈ*�����Or��?ib�$W(���)�F�� ��iuӔ��
�= ��'��I͟L�'�Zc=���K�; Pv���`ųqj�8�Oph��=O����O���O��d�<Y�B���\��U�u��d�C �-xFP���'W�]���	ϟX�I>r,��t#ؕ7�@������}�D��۟� ���Y*�NH��)�	!r�@��SJ#f���b'� oh!���#�%�#)K�C݊M���]0^IqO^d���X�'Y�H���NV�Xzf�H�����R�������To�hZWd�
�$`*!��3�r%V���Q>!���(FR(�p�Y[�����c�8���k��z�� ������ل_�9	���#t��)��7R�Œ���h�<�@E�/���G�irh��������p���#|�%�2�S�*�3��˟\�I&
��~�S��O�x��9��� ����֪4}��w���O ���,I�F~�,C�l� �q�I��I�J�O��d"�I9�	�p����S��+_��2���M�1O��(<O �	"�I����BF�&c�sR�'�"=á�-z�f_�\Z�j�%�0�����F�>�y��Dş<�I����iޅ�� y��f�çW#�A��ٓ#�{�Q��c�*��@b>�OF�k�)ޞm�2�����1J�T����� �C}r)��:0��}&��HrDJ�Mq��ٔ�ʘGgeC�Hß��'��0���|����H�b��c��h;~mz%� S0!�$� ��L{!l�7�4�����	��HO�Scyb�G�I3:0����)#6P�c�T��I+�	-zH�'���'1:�]֟ �I�|j�+Z���0�Z(S�*
�*^���@+���᱋�(r̢��	��J�x7fٳXЄy0�L�)Аa��@ց���t�Te�	ϓC֙�&G����� ��@�ֹ�e�JП��IA�'�O�����$7H`qc��1 :̜[C"OT3�0[z��jB++��(��T}2Q�h,���M���?�� ���-�D	��ːLHD�̭�?I��X*��?i�O�l�Ғ'	�5��'E��X��^� O$\�d�@��8�8�S���0s�Z�ē��h��,Qq�|ՙ0���l�XI��3Dy(���Oz��O$-`Ũ�}e�X���ɓhyj(XRƲ<����������M���9G���W\v��3Odn��C�9�ʟ�C���fBʜ(��	a�����1�Qh�l���34�%K� �"O�,{CM�:�4AB�Q�A�Й�"O|��FI_�^�X)K�J-9
�DA�"O)�'O�bX<	��K*$� P"Oz�s�F�.|�Mk��%���"O\����R+ؕR���L�|-�0"O��E�O��<�(F��$#a&�S�"O
1�VA�D����U�5"�"Ox�R�/2)�NqCS"��e5�@�C"O���,�t&2��ӊE�9�PH2t"O:)�$E�Egz���J�B�$���"Ov9T���h[��xc)�!���"Op% ��$Y� a)���m�r�"O`� �F�8� ��g,�%F�����"O��*���z�H1�)҄��%�"O�$�I�2�A���� ]~�D��"OP0���?��X
���i�-��"O�P��dŴw��9��_14���"O`M�G�X};��m� L��"OΜ�3�ċBn�(gI�G�^XJt"O�y�뎳K��SW�hx��"O�H��$T� ˂p4���`Y#"O^��0�I�'ttS��O�R6~ld"OTpҔ.�{�!
l؟%�Đ��"O^�s�,�i$���\�����"O���%H3��p'�ёj��p9�"OH�r�'d0p�&HB7i�R�X�"O�-Be��
tS&����R"O� �x�
�6
Q�}�1�\�Y�`��s"O$x*��!l��]Rd�l�`���"Oƙ+���(�|����1�P���"O�#%$�`d&�@�OJ�l�ptk�"O�m �["D4�ű���)R¾��"O�`#ҖA��ũ%�o�h��"O���!�Z�f����@���C"O�jB�H�!�HiS�h(��ˀ"OA�&�۱8��1ۺ�R�rE"O\\��/-�������^1pF"ON������&� x�`Q[���Aw"O�eB�Kx�6I�w_�T|�p"Oh��N�&�����K=�I��"O���0+N*����`k� β�Bf"OD���KVt�4H�'�ĆH�a�"OH�YH���]yԬ_	Zƹ#�"O�آŔ2;L;u\�2����Q"O��jL	�.qTmb�������"O�]��|5�1�wM��|Ɗ�)�"OP��&䖯T�@�[�n�$9��s�"O�u!E���K�F�>�� ��"O�a�!�]7�a���,�0�"O�a2�hا8WF}s��)j�X!��DL/�� G�tmM	�$:%�/W<�a��ʎ�yR�]8�|zJϘM��48���i���A�d;�g?	�ܛd��;��ϥ2�ZZEF�M�<A��/k�$��ᛜk��9`�(���vj@��0?�s�A`�U�S&�?��"��3|O�Y�c-�iy��$�:���5e>�����y2�۫lDy��4M�I�	��'� a��a3��9Q���8��Y$��	7`Y��#{����9)
}!�Ɂ&O�Hs2�ٚ��'��>�ɕNJ��`��
"��:&��f֮C�ɧ;^\�y��9�l��oD��牜S2L�����%�d�^��t����P�J�ȓ\�� H�c����Bӗa�,�ȓLx��*���1���1��������z���`y����Y�6��q�ȓP1��A�MX�h,J��r{DA`�<�Q��U$���p�*�qPt�Tg�<��c
� +�C!�L'4	��0jN�<1BK�hl��2��K�I+B�QD�<!ザzR�B�
�E1���5NA�<qD&��.��̳s�_�6X���"O�eRP�E$v��`�	ހ`b��""On�Q�+�G�F(�0 f,��"O�2���7o�%#UA׎k���X��>	ƪ����=R��@L�#g̗"ȑJb�H��� �bI�����~X�%�	�+шx!d�/D�*�n�z�,0!�P�|��#+,������I��=�[�dT�A�R3\�`�
�'�)Q#V�Wi�陑K�1v��u��'��
S��S<nz�mH%ɖ�R�,��K�B��C�IRI^�z�!A"%&��ۇ�</Vh�'B\�7�'n���2Ʌ�a�����V��yr���Ey��ʃ�7iX�,�Pb�y��԰qN,�$�]F��B�'�&�y�KTFD��)�ãPN���O?�y2L�r厌H�&�N��\S/Q2�y��� >���H��@Ƭ����y�˛�jgV�)���.�,����y���U�����D,+S�]��BT�y���7�����ܤ*b��y2hO���C���X���eV����� z���%!f��Y�2�K�Dц0�"O�ea
_�_.��R�U�"�"�Ѱ"O��{7@J�mF0��ҥR�zBM��"Of�*�lT�s�8��E@�4�6@ a"O��(	�!_�s��$@�L<+�"O�-0�+�$���j���>#(���"O<u1%�4U(�aC`>8k��s#�'xୃrV���q�\�L��v��J��H�&7D��%n�7-n`%����è�Hg6�^i��p'B,�D�^eq�G��9�Nd��a��A��i�ȓ^�����*XlH� +(zD�!gM<i0�"~Γo&�����	�([��T\��~�z��	� ��J��_�)͓hpb��>�O��*#E;�)`�i�#uG�q���'&9Ps�
����^�L�F��JZ)/���"O�	��~�]�%(��\v�� �$��]�:�0#�
��h���;��;0�,]��G�%��P"O�lr�M�9߲M9t.X����'���ߴi��A��@˧/Y�O��kt�D�L[)��R,B[�Ј��'�i㕇��7�(��͓�>e�y���Y,NT踱�͔�9\<�W.�j��Ą�,��IѤm��V�b��dG��OQ*#=����:w�I���N ��a���h|�I�x&�c�iͻv"�+d+�!�dZcꙩ�ӮUR����Z�4Ǜf�Rw}�A�1�RZ<P]i��ȔFF<�E�\cK.���e^�n�Z8@�Ԕ�����'Dl��A�P3��i�fT�B��`A��]$4��oQ�r�V�i���������'������LL(�%�5)\P�	�*ڨ�x�K&~L�:W��
N@Y36@B�@0���3��Ph���u� ����TW���WA�f��i�3Mء$��4b��C�o�����v�ћ"�@#R ��c@!x|��A)�㐃�4�y�İ<��@�r�`�h��=�M�"6��b�&�V��x����!�>�|�1C�8(�d��\�t@c�J|�t��ȓKи=�ALπL6���ࣈ�W��Y� ��]D�-���I*O���;N�e���	�ggb��ʕ�8���\�~�(���X=F�8{�>G���`�%�!"~l��Ql�;�0�oZ�Z춅:@�'��Hå#�a�^U S�F;H����z��@p�h��T����-E�!
�a�.^�0����2D�(���7�-�Xxa����=UJ"<��Z)eY �~ڷ䎩��r�S!�e���Z8��ȇ�)�I�T��	�eW�o��-[������I�A� !�qO?�ɄN��S�a�/�Ai���G6��H����>�r`тI�4k�����(fQ��	6�����p>vh�X��g�³C������ ��4�>�*<mږ�V�9L|�̟�Ė�M��I��Ɨp�ذ���C�Zv�~ң�=>6L�4l��~4k'��1vnfl���CF����W�6�za�n�֟��3�ɐ%�������K���8�e�$?qQ����"����X�'�AY�r�Q��OXY8���5{��L�h4>��CdU�ؑg��Dk�	K'�b��gc����_���,��+S�An��	=8~��Bbn��2p�e��q��O2EZd��?�P�@n�`�GO�RC���Mz���(&��|�fֳW�f�:�-�2d�>y�1b�q�f<y�d�SX�'�v8�4��Pp�ʠG�hX�	�
g�f�iG�'�ڐGMЩi�he8Ma1��bg	��F6�̓��`Q�}̓3QtA�6�ij�i�)rhd2We�;j� )́�p�^����d�'�&��P�2A�
��
n,A0�$v�d�N�#Dt&�c^V���BP��s��6J����&B��Q���'@�O��S/�-y��jw�ؐnfҍS1X���3�E�F�u1�f��Vrͫ�&?�`*�uC,�U���:�ܢ��L�BUUG�::ti�բ�*h`ː#$|O�����-r��/\��8q˸l�������Byb��1�21��jKܨ���%�*E���R��?[�m1"�P���?)�-�
\�ȡ̤u�X�K�kذ������<�@L[����T����n4�Ԥ�1dH�H�x�� V. V*p��H�W�h!�� ,��E�i��cm^Lp���{ �58���J��I#����7�ڠ���T�Fhg�i���ZTxZ�؅��8b-T�B(M����?a7��s�L�PB�=�\щ��RV����r&�����]�R���Q�L, �Eo؜/�0j� O��ԊC�@/4���vh�f�(��'�&�d�;���)�� E/�=�I>)�����e
� �� ��ƚ|?9䈯�2�oW�}&Y�%n2���)f�p(<�7+ � j���놺��܊� ߵl_8�" ���/w��W�՝x��\��]�|�q����!i��|�m=h܈���G�xsp0���p<a��ic�c��Ɇ+T:X$0b�Ă7'���%?a�̙5e�N]	4%�uYp��F�d�'��h�h�,�((�k��+�Y�O<���O_1OuST��2��=r2�DkC�ʫHS� �aH�6ufB䉢:��d �Lܾ3�G˄�o~㞌�aJ�W�S�!���"Zؖ��C/�� �C�ɼT��mZ���-%�v�J1�ܖ% B��* �L4��h�5���)H.bY�C�I%�U;�C�06�BЀ���`��C䉐BF�=5� pR q`"�B�ɭwn.�9��C�� �&��3:�C�Xrha&�P�@ָ�q�E��1�^C䉎7UF$٠��Nmܽ�TE:m"C�	�᪐�vO�G1�q���ڻ}�XC�I-,�D����P=x����F�c`.C�	"� dY���QxD%�E;�*C�	0H�,BTf�XN J ���C�	�
 ��`�,�L���N��22B�ɡt�c��� .J���-�&��B�&gtZ#cܾj�\ug._% ��B�	d��E� )�|-8v�����C䉓.�6a��ĒNS>�Ғ�]�`�C�ɥY|1��]�t��8�V�A;XNB�I&=24;��)S&�@��΀�D��B�#8 �cT�V�=���kp�@#D4\C��2@�r`�' �}Á�u��B�I&XS�41"��t̊&�"UTC�IdǒX��̖���r'�(C�- �Zt��Zx�I�(�o�0C�I�1`"̓�*1s���!0Y�Y�BC�	�e��xc��5{�б�C�0C�ɣq F�`rJ�\��A����X�B�ɬ�&t[vM�i�d�)�*r�JB�I	x|���0&X�[$�_>:B�1M�^T���;b<	�BG�DP*B�	l"z����{T�!Y����C�ɡ1�H�ÌV[��Q��K=-�C�ɐQ���1'��7�\����Rr�C�	�u��H'J5f�X�S�s��B�!������1޵	��]�w�C�Ɇd�L-���I�T��-��*.I�C䉷mFi{���Cа���G��r¤C�		�0죓G��;�����Ƅ8LzC�	'gj!���I�,�ՉֲN�VC�ɧL$U��f��;�d�BW��O��C��^�(�ٶ^q,�a���KT�C�/O�L��6�R�lD����N[�<��C�	�����dI؃p?J�)�
 ��B�>���;`�'P��Z�,��L�B�I��8�Ɂ������F�p=�B�	���B��ؐQ��-��$���2C�	'v�1	��Ej<��B�n� K�.C�	�mͨ ��<P��ũBJ ��B�ɥ^R.Y�+O�>���"�#�_^4C�I
.t�T�/U6�]j`�O�X��B�	w�v4獄�a�@�#a"-a��B�0:F�a�D�L
H�Tq84B�I��B�A�Q�Ū|q۵�6O��B�ɞ2�TX9e��J������fB�ɿn��Y���^����%왠9?�B��0'�E���86���X��Բ+�C䉐SK.���ѴY����Bo@*\zC�	#a���Y���펰#0i��F�pC�)� �㣌��|����ͩ

���"O*�V!UjG���r�?O�B�"d"OD��7��)C\��`蛃l�*살"O�X{%]�ȱ iT0R��p"O�H�"-�n&��Ӂ�'a��"�"O�� ��i9(}���N�y�Z"O:�����F�YCo͍4h�4�V"Om��n
��6���&9DiB�"OΠ��k��U�r8�@�9B/!(�"O�h�f��0�,��x9 *e"Oh�ʴ8	^T���� Q�&m�&"O�`cED�j�*�m�<���A�iH<!EG�G��0��1P>�����<ya�]E0�E33
C�I��,R��Hy�<�����C,�u�h|4H�(�jQZ�<��a��JNpk��c��Au΋V�<�V��W���7�_c� aѐ��S�<1*�{����zF]�� T�<���,]�B���K<czx!PO�Q�<�2�ؖ \2؀s��*���(NX�<�e�8}Y�~�pb��S�<�5˒�w����$��9Q�E
+H�<����� �Fɐ�d�d��`I'cC�<7cW�/�qڒ.UyZ���}�<9��PRC�"L�X+����!z�<YF�I�u�r�e�n�2 �� �s�<�1l�Z�i�k��f�T� F
�u�<A�%�,wꆀ���ތ�fՀ7fHt�<�d��9@	*$
�p�,��"H�K�<yp$A�1*�ys%���@F�<v�t�MT�W�oi&ؐ�/�\�<i%j_L�X,`���(_Gx��$��U�<ٰm\�j�F���ʈv4x���J�<c�&N���a�ɉb!��Q��H�<��΀3>�N8���RUR5T|�<qC-A7-8r�r``C̒5N�,��B��{bn�S��B�.=<�YBi�$~�B��9$j1(�%L�k�`�4y�B�	�	�D!j�e 
�4��"N�y�~B�I	k��Rу�+*!����P�2C䉗%h��pc�^	d t�̍�:QC�	\	Sd�����Nn��s�H0D�$�Q
�1~�K2 �.��ū�#-D�Љ���?@�����O,\���?D��Qt��x�L;�gT��`Ix��!D��ʓ��-�t�+A"��]���A��!D�`3,�<���ªE#G2�}I�?D���A�	��0���Aֈؕ�<D��KD���h�횈n9���5J D���Հ{U``׉��O�����L0D�,���F�Z�n�I���0>�$�*D��֧��ivep���0Y�P3�a'D� q�/��!RQ.W=O�l��&D�8���-L��1�R��x�#D�t�B��3[�HԱaE pOZ�;�%!D�PW��%�n��g,Ű.A��h4D���fR�!�de�����2D��K�G�m&؊��ͿS��%1D�P g���p��bֆV|���9D����Iìal�$��6�̥*T#7D��Gƚ�	��1V"I�Ρza�'D�p�+ǈ1 �R!�6+�b�h�h*D� 1!��W�R}:���+.b$be)D�dq	^�c֔X*���"0��Y�o%D�� ܸ�я^�̅�&,�n`,
"OB5゠�'H,��-{T�<�0"OX��6a��*���&/Ծz�f�Ȑ"O,��&9�YAH�3C��p*�"O�����d��pF�0X�{�"O�D���w��i�Kǿ[.z�!�"OR�a���V<h����.p�|���"O,R���Y��T�D�]2$�$@T"OD|��(x{(-��Z�R�L9���`�Рv���
�����3o+���B�.D��ǒoD֘r�ֿ=b^�AG�,D���#Y4RBB���!&RD�CN)D��"���hQ�PcQ��^��@e�&D�\⣊��x�@d*��\�
!,:q'#D��ؖl��D�����:��}��)!D�h0��[+q��u��$>��=��"D��!��6��i ���v��8��5D��86�׸H,H��e�
%�i�14D��i��
�7yqI#�I�zAZIt"2D�p��/o����q�F!/�pY0B(/D�Lx#᎛2�&�8u��&5f�µ� D��@�.�Lb��iwa��_�1��>D�\A�@�7Cv�Je�P(9�!�h?D����!���t9�� J�Ryö�8D�|j��R4L�tP��N�T�,j (4D��A���v�y��a@4q,II�D0D�조s$`�_0vQ�9D���g�/q��@��*qJDH�g+D�b���-Wfmr��ؾH^8p��'D��z�̓�Z�b-�dY�1$�i��"D�h��8v�D�VM܌>��5�s�"D���C[?$���ɛ,$f�0��L5D�l�)�F|��"i�-_����B1D��@	!WQ䀊���4^���[sn:D�̚�+2	&4p҇�=]}�UBa�=D�d��ø�=���E�<�9�,=D��n�\f���C69V ����(D�0��jį:�B�ې�J)��с&<D��0���iE@4ʊ$/�3am:D��jW�"c����'�|��	;�e�s�<���{!�x���6'`��S`�Z�<1��/��#�.ش*'&�����l�<�uIEO��t*�ă-
b���K�^�<)��@zZ=x����y�(`2��[�<�AQ%$H���-�QqHɶ'R�<�¦���4i�`"��|��@!j�d�<it�ӣ��q`1�������d�<)���u򔄸���f�h�
 G�b~��'0�u����q\��a!ʟ�D1ΐ�'�X�
��Cf<q���X�C0(��'2�ԹNP�M~��zq�Ŷ7���Hӓ��'��M� @?�[Y��G -S��'�} �gI��$�(�n$	6}[�'�<��&�#A�J���2�4r�'����c8\�R�0��=l����'tݫ&Ȃ�+E�\J�ϐ��,�	�'x�Eð�7{���F�΢==|8��'߈�:�m۶OTLr6�?�ht��'�:(c�O�j�P�cψ6`ġ��'��<C���9p'H��N�6(�X��'��Aӂ�&(p���X1Qܴ��'Dr� �C:\�L���"d�	J	�'��!R'!�@O��O'�D��'*����� ��q�hO�2����� 2zB�P*LX�KVu'ʽ�"O�DcMó�����P�"x��"O����[67���.֦~����"O�yq r���dg
�e	��)�'�`a�4aC'XVu)6O-}�x��'�x�ؒ�P8]4ţ�#{'�l��'v��RFϑc�R��q�I'kl|ٲ�']�pRp�[�&���!1`Pm@�'N� y1�����w(����X�<%n �"@R5 Ղ1K�yQ׏Q�<!���&HԃU�� Cir=�c�WL�<駅řN,� 5�S�^�H�EJ�<�U�Z$z��	��Yz�j2��Ї����@�9'�,�10��-ɮ$��vӖ�a�Î�@(yIg&W,L�.��;�p�@b��]��U�q/��f����g(lL�d�ӵmU�����yF���ȓV� �*BFP6@	b`���3(f�$����q7���2��zf��8ZQ<��{�>8Q���'���*@Jҵgi
5�ȓcA�JmI�	fVE"-R�	��Їȓ]�N�r�-Y��|��SM�.H¢Y�ȓN_����C�"�������2�5��X��R7l��(\K���A�Ȇ�}�(�� ҤK̠(`�D.Q=����^���g����KT�)&�	��wC@�гG��Q,*���L/z�\��w�r���1P;(Q�&dE��>�ȓ��æ��$-#4�Ә4�"e�ȓq��%�7�TZ�8�ޘ3G1��S~�B`�Uњ���E+@�p�ȓk;�YJtO?x� 0�B$GW`����o������,t%��b*�lF���ȓ"�Lr`J�f������GY*�ЇȓI(�c�<!|&����Y)}�BY�ȓF|�<sG�ڞU"�%�G�J+�n؇ȓ��)��HҜu�<u��b\15Z �ȓ&b����]3�9y�C�+,��ȓT%�j@t��$k f|t��>P����"�Xw�A�9Tцȓk X�FJH�O��a�vL��, �ȓRl�)������I��D�;
���+B&�S����/h���2�Ab~��*G�m�o6�D��N��̄ȓE�ḇ�Z�� �T��Y���v��U�ε<�F��Ɣ7⊍��;�<#�oZ�8��ħN�Zd���ȓT�*�;�O���D��	��(�4��m?2T�QbC�t���j�EA�F�i�ȓV�`� �C�`��Z��V�@��ȓi1� �KX+d2!�͆O��E�ȓ0����e��t���&SOm�M��)�PP0I��r����f,NZb݇�VW0 *�$
��F%����"9�l���O�*���)U�q�<UX�u�"O�y���1�\���+�\zP"O�Z�KV\�H��
:�t��"O.��,ؒ6 ЁW�f�f��"Or�[�#A~Z�8q�D�K���E"OZA�0�ڡy�>��c'+�2  "O�D�*�'_��Y�$'Pf�
�X�"O���C�H?7�
�S�K�p�R=ie"OH�IAHJ�'VXIE�C(f� s$"OZQ�r!ːI��������g��l$"O� �����7o��4fсZkB���"O�YS%^�e�����A�|�P {7"O��3��9�:�� +AL@I8$"O��K+	dh)�g%5MA���"O�3����J����n;��6"O0�S'�S2ND2|2%N�	2�d�"OZ�!�Qj(�PD�,t�h �"O�)���4�����aK!`[l=s "O"�	���jx��%\ FER@��"O���2��,m��X9�%�"h����"O|̃���*�vEJ��J	�"O�9����q�&f���L�!"O.�a��Z�����Tŕ-Y���#"O"I����I<I�V ����!"O���,ԂJ� @[ScN�i{Z%ȁ"O�-��B�o 4a���ԗu>�0�"O�����lM\���G�Ne�dW"O�����9'j�!�F9PXv�ʗ"O~�B�Nۜ-��Չ�=W��"O�\['�FȄ����P�kQ����"O(�0�D�q���te�(���yv"Oxm�Gϒu�T�eD�`�V9�R"O�t��U��%�^�,��r�g 	�y�M[�@��l�iă��@��y��Y7İ[R��7A� �	���y��1N�� 0��<'.�)��̳�yB��QR����c�.!V]�����y�g��h�z� �G��H��g>�y��$O��Yavb�9?0J�x2OQ��y��Ѓ0?Ȑ���*>G�qq�y��LZz�)k!ϔ52�B%����y�mW�����b�+�����		�y���c?���M6%��Ű���yBI�{��<�QǏ�?zy���y�UGz�����a'� 1�!�y­�8eq��q��Ѷ�W;�y�"[W�Y��jN�xjì*�y�Af����R�r�b���1�y�eXE�D1qN�Pb��K� ���y�#��9�Z<B�	�G�4���6�yҢF�_�eIу�R�h����y��	s�z��`�B
R�LH:��9�y���#ul4�ehK"[�!�'�E��yRBU�u��Q��X�_x���
��y�<�(��e�7\���[�EZ��yB��\ʱ�o+Wf���A�y"�ĖU��\��c�(Q��#&�^��y��2u+$��#"9�B�Ő��yr�)C�!��$���!��yBK[�'$Qr�hԖy�ε��ԧ�y�àG^)���U2y�P�xd�@��y�BS�b���*� ݛl��(�L�yb�C����$�5i�Rq��j��y�L.��Њ�f�eR�@� ��y�a�nN� "h@�?��D���yB�5�n-��E��.R ��V>�y"�S:sZ�������RU�<� �D�y�ZRbF%�IޮG��qQ �J��y���f�`�Ĉ��k�QB����y�
Ǥ7�m�t�G�:��g��:�y'�J����TJ��5h����y��ʶ2�X���jF��>�i����y��N�B��+�~,��٣OG$�y���H2Ptx'�Y5s��-���W��y
� 68b�G TBf�H1�bo�U�"O2��1�Ε\Z����Q��0�"O���l�,`�,��V�L�	V$��"Ofq;�"�&b��(鷅�8���Ѵ"OD��fIN5@�)�M!��<�"Oduz�<�����"ׅ��0	�"O@�@��G
���� �X�@�����"O���g��:�J�Jp@U6����"O�q�IV�p�:�Y�n��JN���q"OX��IA^W�`���R��I4"O4����ʃLK��S�!�r�iW"O�{�B�h��t�8�	��"O�cB�	�}�٢�c_%e��ำ"O�I��l��t�H�B]�$���"O����/P�R�0 s0B_����"O~�sH��x�8�jg�Wp`ȡ�"O�a*2΋%�����_k�ĉ�"O���a�E�jτ���Y��=��"O�}���
ixQxQ��W.���"O���a߻=ߒ�IsKB�I�|�r"OJX@��<�P����E��m"O���qI�:s'.�I[�D��"O�m��B��#U�Qȁ�. ���"O��H�%G�W[Ā�'D�c�dA�"OjE"ŞR39J$�ڡB����D"O�U@��֊0(HK5��	U
I8V"O^MH���$f�t���W�Vnh�x$"O�a��E�ȪР�@��Y3�"O�=J��A3_:ZA	`͐n��0��"O>py�M�9L�U��k����4"Ov�aB�O��R}��D1Z�+�"O��Дkި:�e@�����$m��"O,dc�NLS�|�c)Y;�@��D"OH��AGW�2�R�G��F�(�"O�A�'��&�@d'�6^���"O4���ؑo��`&[�R̈"Oȵ�U�O�@,:�c􄏆NF��i�"O��#��eM�����%�D�"!"O %�lNudB@˕�,J~���a"O�I�)̂e��8�bC,Y�0x"�"OP0�k�7-d�-)��I�l!��[���u�\E�l�Jtj
_!�D8\Jj��d�>:�&�3��W�Y@!�$Q�*:U�'��e�TD�򁀈,!�$���%D����a��Py���
A���N��	� B8�y�'ۨߒȂ��9V��Q�B�y�s�J튤eB0p�Љ�ς��y�k�A����Ǯ5,v*4Y�cF��y$@(k�t�E�G.:�=Z�O���yRh�	~�PZ2EV�0�*��I����=y�y�㋲-rT� �`V����y2��r���K� ��^)؄a�Y��y�&>�݃� 3^����$͞��y!:  I�3���AC���ToC��yr�ڦ$
6x@'B�569ڡRD���y�-�7pڨ4����+��Hk���y�ߴ"�p��_sz(Q����hO4��$A�`y�q0IC,����r%�#V�!��a����V�ɒj��ty�DA�*�'�ў�>�����mz~$����i�6���� <O��$6�I(m��*�e����RFV*�
B䉘n,�`+B8Kᰔ��-���C�	K&e�'�V��X)g�>l'�B�)� 0���z�手��� W@,����O����W�B�D�J@�]�B�x("e�3?!�dU> !�Cd���M֒%Z�B��&(!���Y�����(����¢A�`
�y�ɑsG�m�ŀV_~V�h�B$O�C�Ib�l�EKX�P�B�B����C䉷 ] ต�N�Y��$�_�yĬB�I���1D	N�FoJ����2�hB�ɺ
��A�g�h�6�2Tj\9bB�I�+h��h0�O��Ve�S��<
��B�-  �,놭�p�(	��,GC�I0?��Y�!d����L���V)L�B�	K��X҄O�v����N�1/�`C�� _0�q���(d�8��&U��`C�I�v�|\�Wk� {l� ��͹39BC�ɛ*�]� &A�-�, ��V��B�	~�����J�)`���a�h�/D��B��y�h��c�Ԭ �� bqd\�o~B��+Pǈ���"�:C�x�j�o�zB�ɟp��xa���R>	F�	�t;!�J�1|��h���&m�9��L3�!�d�K�R�K��Y�RX��0@E��!�$�/W�6i`wg[�|�P�7�U�D�!�
[䡺"n\><������	1�!�_./B�`��>�-@�(��5�!�d�/k`t�+�@Մ!c� �A��h���N��@�)F�H$�`(�K�+e:��+�g5D��ٵ�`��I +��C�X(�4D��0��\#{�>�ò,E�(���<�$�Ox���#B-�F�Q�����Ju�џ<D�䣅��DA��/wV%y�CЊ���;�Ovj�"�3j%j C!�Z�8��;%"O�X���G�>�A4�1^�N`�G"O���؅#�pY�F-��2���Ku"O�q��d�;��1�i��'d@\2T"Oج(nR"inޘ���ƟFPFP�p�|��'iў�ON��퓶n�4��¦G�i��`��ODQ�hڡV:� ��&.;��-J��Ik�OI
\�AD!�z,kB�.Ĝ�Y
�'����a FӀ��KW�^Ϭ��'M����L�3m�,[�.��D���
�'��ą�'�2�z�"U�Aq���	�'̖�)HI�!���W�3
Z�2�B�)�$k��Z���A|g�I��C���=)�y�X�PLRb�O�D�ɛ��hOt��Iׅ
dhp���B�8 Iq�̓,�!��Q5d�D11�~b��(AW �!򤏸A������>$=����\?/p!��AW�h�!���-A�rt05	�M�!��8q�l��fϘ'E��,�������	���?E�$I��c_v�P2?5Xts�C�<��O<#~r��̓B�։���L�j�x�R��~�<���]=���T�%��ȣ���v�<)A��U��1BZ0�� A�Xp�<iK����01�eN4@AX�ğh�<�$N��� a��ϔ�@{|�R���hh<I�o~xљF���u����'�ўX�'�~��Ө�3!�V
�R�L�(x���>�4����]=On���jЯp/�"OT�u�-
�"�R`��:p5r�"O���^!���;`n�?�����"O�k�ŵ{����$����hq"O&�ƥ� U��y��-, FН�7"O.�����0)�V�Зl�?)���J�"O� ��Y��5/�l�q��؍)$����"ON�����y�;�g�`n�*�"O��q!Ԡ`��@��
�0�̘�"O����g�s��q&ٻ ��0kG"O��:Щ���P���D����*D�X���^.n�x�!n��Gu��� L-<O�#<	�i�%]��(�&ɜ.,�k�N�L�<yb�	<5+!��*3�&iIDKOJ�<���
~m����
ӧ~���1#��F�<��-�/lP��O�"^QX\!�DJ�<��M�)�zt9��
s�ف��ZL�<W@|�$0������w�K�<�uF:�.�r�c\���4*�Fx�З'�>-���1���S��H���P�P���l=��X�hɭt��P�W�r�B�	2@��t
�h;��9���*��=�	çE�~p�&��% 2�h ��+3b�ȓwtX	��L�`�t�t� g��p��zk��r�F��O%he0���r���ʓE0�lj���x$� g��9���Dt��Ґa[[��`���8�((*I:D��E�a/�L��m�0_�$D��5D��X�- Q�J���:P20�*�f2D�dٕ�L&��BT2'_��IU�1D��A�̽&�)j�(�(����+.D���CN�)���!�0�Čpc`!D������ܨ��r�X�9G����� D�`�h�tE,| &`���tH�Q$<D��q&��3iﶭ���H�d���ҧ;D�����W$6�A�	#\�h�Bf;�$!�S�'x$����Hǆ0�i�FG���ȓY/x 蔣��h���`JI�.0�Ն�.Ap��l��9:�	t!FJntمȓ(- |B/V(R��!�� 3%@a��j�t�2���?{n%Rh`���Iq����l��M&<HTI�Dӱ��q�qC&D��&$ߙh��)03��4/B�}E�.�	e����3}���P�����3����B䉻J!����`W�f�`��a!OfVB��K���ҦH�.;��"ʕ	v�>B�T�fH"]v%� `�����B�I/#"} �&�����R�j�B�5H)��ǹ vaɴGQ��B�	1O/�iQ�ƃT��O[�~����0?����4�h���#HQА�%�R�<q�L�M�%�TK��RQ��/�x�<��l�~;t̙s�O�^�C�t�<y��̭fxH����u�=ʢ�E�<a�м2�6E�4{�UJb�Y�<I$eD;R��e��!>?���ύX�<�$�C�ڥ�a���W��!� .՟��IQ���QTkI�`�x����/NXT��-D�X
�PB�����R�1�D(�8D� ��L#oG� �f�U�6 ��5D��w]�̀�!��^6<{R�7D�d��Hꊱ�����75��s�0D���B��)F����B	Q6
���F-D�@�$F��^rU��<���D6D�졣.��D�Lm:Q��S\� �BH3D�8@2ŝe�tdJE�wd��!B/1D��!���1%H���(v�(-a�%5D��+5���8})r�G�Nˬ��5a5D�hpD��7n�2E녟u �D���1D�(�a=��8�OB�g�|x`,D�� ����\(+���#g���B��"O愸�.q�jy1��[S��d"O�=(aȌ$�Pl���B�[O�|q"OJD�"��2��b ���7���"OBAJt���[���IF�:��,�v"O��*U' &�R �I����d"O080AQ�c�͸I �J��5��"O( �SIɛko܉z�Dq�6=C�"O���/r?:Y����.�p���"O Q*dI�"}8g$L[�<��"OLh�'҅�,YՀ<H�Va#�"Oj�J��'|����B�n�4�"O��" Ȳm���+D�6��{�"O}��l�P:�Ap�� ���"O�I�M�%Ѯ �Qd�n��H�"O����7������~�t(�"Ol-1$L�z��#C�{�4�g"O�!¦V�B�\�[��őn�zL��"O��ɃK�������S�>e� "O�!����)b�;�g���\�"O����H͙����3gI+x���C�"O����ʕj� ����z��e��"OH��V�� �r�Qu�1�D0[�"OD���'ְ+�h|��bV n�T���"O(��)���J4raKF�դ)p"O�T��6I���3A�+u���Q�"O�`��eG:]�����d�,`"O���!Ѷ~yJ<�ꕼiH�-R�"O�����\���%+�6-b��t"O�;�@V�Y���VnV�{v�X0"OF0�ږ�&�:�Ĕ2I�d�"Op� ��(}�����g=��St"OvA���
x��ߚCL�C@"O6}е+��i=��Y�X<B1T h"O~��@	]3�b��d�)t�>�b�"Op s�j����R�З.q���"O��)#�
j����D�2�zp"O,�`�NB&:Й�CCp�|�6"O~}9ei�r���s&I�(
2��"O�p��$�¤�+��# ���T�'[�Ę�(o�5b#'G�#5Җ�x�ބ��'7���V�%j�r�ZT-�$lj`]��'��k��Ip5h��F*_|BM���D9�6��b�K%Be�a�Ns��	8Q"Od��L��d��#�����U�"OPP��=m:�����Jf�q�"O8�aQc9����w`P$BPu�&"Of�5��S8 Y�+O,!@�"O �c��3���`H �rp1S"O�\C��A�8��(�)��/ ��K��Ia>e�s����a�'F��g>��)��7D�س# 6a�J�y�g�0b�|=���?D�ę�j�m������R'_�����?D�����E.T�����d϶)2����1D��4�)0�H���B,;��y�pO+D�|�G���-�����J�0�i"�=D��j3��7��%�SG�K��Ƃ<��O�����G7tQi��hV`X��_�
^C�ɑ/���FL</ ��`��c�8C�	,D�,�`��Үj����―B=PB�	t��,+�J�2�j�2��H�*B�I/7t���ϝ>@�����[�CغB�I.?�V�)OV!
ܯ\
�C�I/[$81�Q��W�*9�p�#HB�)� ֭Z��@�q锘�V.�sL�ԙ�"O`�#��;��ajNۀH�^��"O��gi�(:��q��jF�^���P�"O��QvbE�l�D��=��Y�"O`!�e�5-d!C�?Z�D���"O�!�'��� EcR�A�@�tX��|��'[��ʣ��y��
�]�̀)�'0��d��L�F��ʘ,�¸8�'�pU#�X-@�tt�U-��m��'�R���FӪm6��:dg�*N}x�'(��rd^3��A��Bϓ{���"�'t$8�녾�N��򊏔x���3�'�F�0��|l�����_v]J>i�����&�������;|@����ڽ�!�z�̸b�	�6K"y26ŝ��!�$E�!0�j�j`��DN�x�!��H�mǂ����c�,��c�(~/!�DIl��9I@-�� ��ţ2h�2!�Բ������]ΤHyj�2���dB#`�`�Q�Y
�
��@���'�ў�>���A1�\�bJ�%B���&9D��Kd�A�t
,D���6)C>@��e5D�����r]p�0G���<�n�Y�C(D��H��!��;�B�=cX��b�9D�X#Ǩ 8f�1T(���2���4D��;�I�*aC,�&g�A�� �<D���U
в}��("0�\�)$�kp�:D�(��'�j�$)eb��Y �|�ao5D��U��+)� t�en�d�)5D�<�Q�<%Ȩ�"s!J���%D���Y,{p|�� �Q�h���a1D���c.�W��cu���F��|�Bl<D��խ�c��y"�{�b����:D�X��A.~�a n�z��%��"D��0Nˍ43�%y�NU���Pe�!D� ���F�-�2cT$����*D��k�!L�*3���ߏy�~�چC*D��aCb D�h��V'��T�A6�2D��Õ�����¡�"l	Rh�0D��ӵ�Y�f�0pG( �ܜ�e*,�On�ɂGh�h 4�(9�y�⠍"P�=�
�#������S�$�0���P<L8�Ն�\����&M��9���7d�8���_k�L��+Әau�y
��^0U6���/� ��S���;��l" �?��*�P��D�J3Q
̄����J��ȓoI"Iia�I�<Y� 1�	D���'	a~���9X�H�A��ߚ��լ��?ٌ�8�	м�A�(o��y��
n�|l�&�FE�<كD�8>�t��IU�b�4J�*�D�<�s��[7���`ᏜFt2/�|�<q�B޲X�BxrSi�Z��	�^�<y�ƙ���E1�]r������p�<a�Mǡ]&��R(�S���:UF�o�<�enH4�!	$D��ʌj���jy�W�D&�"|��غHR�	3!�AB���G���>y�O,tI�
mò�j���,\/�c�"OMPh/W���y��R�L/��A"O�H����֤@���W�>���"O���p�ʕ1��]�<Ĕ��"O�!�u�G9Bi+�oLc�>��A"O���3�B(�`T���HI��
V�|��)�B�Jѡ���Rp�	`$��B�$0|OD�Z��������0��8��}��S�?  ��6F��x�'_�~��"O�ю7(��pK�kb�
u"O��d�X�^�j �	D7X*13c"O��M"hX�	7*�r�ށ�b�Ix>J�-5���{C�!��3 E�O�=E���
�3c���t�Ԑ��2`̍�r�	i����i��"��\ x�����I�,5$.8��q �Zt �Q4��C'S��ȓ,ت��K/�h���Ȅ</:n����J���ˡ,�.|� @/S͚؄�n��m`�V�$�5�,d�fe��	d̓��ln���f5E+�!�x��	�<�?E��	�G� ���_s���Cτ�e��|"�'���4�\�cLb���#�[+����E7�y��E�d;VIz�˰q�4�t����yr�ZQӦ,S��S�s�6��㪌��yBjM9z(`	��� �v�B�Y����y�/�p*^�� �v��8�ugR�yR.Ƅ\c-D�w�����8�?����S��LyRs'�/��ܢ���ꘔ'��u�)ʧP��ӎ�,z%�0�%eG���ȓIt�����K�E]��q�E̞7����ȓ	���F� ��̇�5N�U(B"O�m��lX9{�؝HW
Pi�Ȗ"O�� ��0#4�m!%�&1=*ؚ�"O��p�Q,c�<�A��V'|86�
�"O��� �l�;�A�`y��!rW���'<�	o�3?��N�I�R4���95������۹�ybLU�1��T��.^�)���j#�y�O݋h���8#IE��D�3aF���yB [?*; `@ԨƸ(�9g���C�I�y����$��d�>(j���$>�C�I�T�%�Ԋ�+E���)�*V��C䉔v��XZ�l��P�y*ѫ��]�:�=�ÓCL�}��?`�СCh���!�ȓ]�hP �C��CBL��Ǌ��J��Q�
�+��0S�v�:w,��&��ȓ(���D*_9fB�!!�!M�4%���t~bʛ�ܔs�@�d�H��O��y�E���6QCkmxⅣ��y�Vg<���!e�����Fڏ�y�́�n�����9]��x+B�L"�y������ms�� P4�M���C��yr�Ħf(�"C��tꆴ� �X0�yb�>^=B-H4�D%Y�\���e��y�� ���V�W���u�Ķc݈4�.O �=E���"'�ju�Tb�=W�0�u�R�y�(\�VM���aH�&{~��3kͧ��'"���Ï��WK:xV�D���k-2D��)D�"�j0�䢃�x"	�`�2D��p�-��uH���5lA�_��y�
2D�d ,a��	�C
��Ie�(�G�.����`U�ʯ~_$�+V�Pg)��ӄ"Of� U��*&���bث��e(�"O�\Q�Q�b��jt+L(�6�P�|R�'��Oq��k��ұ8�5 �`j��t�r"O�4j�lE�y_\4#JH�aDt�p"O���U"´P!@�J0�V.H��	�"OJ�.��}�(�ᆀ	U��l�"O���'N i���DN�dՓd"O�]H0B�?KV%Aw`ݞ>�����"O��	�� �(�����aU.v��yc"O�Y���0QB�t���lؘKT"O[c��%�vP9e���-\T�("O� �<s�����t�U�F"?O~!��"O�a�t�U8@�z=AW�� <���"Ovu:�+˛85��x��	Ծ�13"Oݹ���jZnx�v�ӷ;�`���"OX)dƕF����D�[��)[�V�8��C�S�O���X!HM�[���X$�R�[�N8�
�'�x�JZ�5;0�!Tj�C�Z��
�'�RmRQ�[�L�r=���5����
�'#fd��Q�k���ɞ	*� ų�'SP�A�mM:kn�vꉽ.6�k�'tx��Q�-y� 5�hIP�}�<��BÌ����M�'T�A4��u�<��nE�$ne��CN��01�p�<I6�B+
N2�;�H_<T` ]�W�Xc�<�ĭ]�����"�[�_1��@Co`�<�1FR\�T��Q5\�ݡ��_�<Y�h�:lX��	hy�1s�%�`�<�6ɐ52G�%b��V���)�`[R�<IQ���J������^�^d�<9cB�{I�tc��D*4�Լ
��-T�����
��~�!�G��|d
,�p?D�\r���?�T��H���ٚE	=D�h��$H�E�h}� ��
ms.���D9D���	��F|Q���L>^D�b�6D��1�>S���Rf#�7	��E)D�\I��=P��������s+#D���e$�,4.>H����9^dص8��"D��Z��5HŠeI%��a� � D�8�7�ۓX
�r��ۓnXa��=D��8 M���}��ܐ{����u�:D�$�`L7)O�yC��\��^���-7D�c�/�w㘬c�f�Z���<ړ�0<	
��lɉŕ�fB�| 7�m�<y�c�LDD��P�-BV���!u�<1�U�R��E�ԓ8��d�CH�{�<Q$�?�u�c!�gA61��]�<9�� |��8�ŧA&�j(#�MJW�<�a�ܡB�4��ƙ��l�&_W�<�C�z�Zq��[�E ZUp�m�QyRY�8%��g�ę7GE+Ѧ�3�� �"#ըVF!�&V�@e	�e`���q�B��m'!򄅏i�~�3�	�]���֧܅f	!�ĮA����00O>t�&�ˏ	!��׼v����������:��չR�!��A�w�(��;d�p��ɒj&!��Ɓ�H8�Pn����,	@�O�Q!�\�p'��g�d �Ѳ���N��I{�IC
\��	i<�䦇6Q��Z P,�ְ�'%FZ�<�2̛2;���N_�RvȔ�t�T�<�bt@DM�P��G|�����j�<Y ���L��ȫu���d�d�2��Rj�<1s�� ��`th�=��ҧ.�[�<��Pcz����I6)~��i%�Mrh<1����YRL-dA.@(����?�	�'�~�v捒]����e�W��\4��'Uԡ8E��6~ID����Z�Di�'�$c@B�4!̔#�)Ӝx�l��'H�y���Nu^�Y�	l	�%y�'z>!���>PC@
�J	<f=�����<�*�����{(��k⨍�KR<lS��'1!��ͻc�fp��ְ�h��5#B�nJO��c�/�Zaj1��)��<��5�V"O8��Be\�)���
 �߄j ����"O�� ��K'c�����/9�x�"O� �aQ�HܥyN���FT�L�h�"OT�+7KN�"LP� M
�V���"O�����F�L�!����d���"O�b�(��)�\��[F��x�<��&͘Z=b	�g��GL����Z�<�U�(Gք�p �6
�p�IQ�<f��/(�\��i��P�!��X�<QcJ[7	��pٖωTRy�`�T�<!���%��:3aW�IGHd�V�Kv�<q��å(�:M��ЇC�L@����w�<��@�F��@pB�J�m�W�W�<	gd�-"�6e��7[J�aଞT�<� 뚭�<%	�!�6/`P٦��g�<I"T�t@��c҆N �%�p��d�<A� ܗUb �S@���J�`����U�<Ad�@(����6,�4�t\H�EP�<Dc@."�"�.T�0*�AxHUO�<���[5%���v1�#�kH�<	ѥ��^�,��e&�X@H�@�<kXT�IHO�<g��e	�\�<q�H�>b���r4�G 2W�)�dM�D�<��|Sµ1B��%`���� �LC�<�3��K�Q�#J8E�f��A�<)���4?1(�1���5Ն��'��t�<A��Z:D�y�@+2 />�1j�s�<!��M�)B��:��ޱ240��p�<Qk�=+�,�nʰ9��YpN�b�<�Sf&#��(�ߩް�����]�<�$�V�"߄�1�n�m(hq·�^�<q#��#:b-is*�8��jLc�<���W+�Z��Й�|���WG�<�N6C����b�;s�ji��@�<y�Fʅv+��zH>+�9h��@�<q��>M��*]�M�J�CGk�z�<!t���,�<p00N�SZ���҇Yt�<ّ�]��� 3���U�yKQ�Lq�<!�@�*Պ�G�8���E
�F�<��L�< ZI�9J�7!�w�<�@D/Q�P����M����ˆ|�<�w�-,��9ju��3���VK�x�<�@��"�*�9��#i>�]��N�r�<i!N�'I��i8�� �,;&���_S�<�fNK������OJ���w�ON�<e,J	&�pM�#��$a�)����P�<gDT%:�k��*Z����'�A�<��	�'�.m��#�$���`bJz�<QPcKִ��R.�d��ؒwR�<Ic@�k��x�̜�ePv��K�W�<��H�#:���&�X��Ej&�[V�<!n����3�#����N�P�<�c`ŋ3�8�@�R&6�P��#�F�<�TiL�(e�)��ʜ$Y�x���mTi�<�ӭ��YF�N��1`�Yy#b�<� ��*��Y9&���L�A�c�[�<��+�$$�n�z�MQ�;�Z�Hei�_�<AE�F�lL�dY�Jw X#L�t��y(Le@3�
>�-�7-pZ����J�6����񮁒�d�x���ȓ
g81ir��0Or��B(s1�Ԅȓ9lD�s�G�
{�	�B����0�Dx�#P��F�an��zH�ȓ }�	���+eq&�2gJ�k(���ȓ(*�h)C	·L��*��VT���F�Τ��i�:E�}b��ѬrΤ4��S�? �,����Ae�p�f�d��4"ORD�ǩܗV(Z�%$m�E "O�,1�(W,k*�XqaDI�`@a�"OpL "�32��u3�E4;�3'"O@$a�����	�1�HJ�2}C�"O6)pD��ʁ��/U�y���K&"O�Q�1W~���2��.�����"OL��@k%8dTS���e
�Uä"OĴ��� ��		A6{�"��'4@q����0�(y��H�u�#�'�s��0�Ay�Ŋ3?�&p"�'ע�i C]$bI*`)P	V�:.D�	�'�J�䫈�k\�P �A>8BnM3�'����
���y�D�#.(�H�'*4I�-[�h>0zgᙑ�����'����W`�{�=ӶH�\����'S� ���B}�|[�
�XtJ��
�'2z�GoQVY��Q� �5Q�^�b�'\�Q#�n:Cq����&H�5!8��'`�xѦlP#ڹ�@ӧ'n�%�'�>��M��If�qk1(O%w�h�'3F���F�D��k�CJ,���
�'�bm�� A�X̊EQq�В{c�P�'��5ã?I�D���
woZQB�'�{�l-� �V�Cި�	�'�`5)u゠ ����u�P�jZ���	�'��<��	�"h�1z
�f�6�K�'����.l9�p�vƖ�^،�[�'ŤQ���G�.t9�.+z�D��'���P�j��m(�[:!�N�q�'RZ�i�56@�uA3�[�/���
�'�����#G��\A��K�����
�'����B	@�Ln\�� �(�
�'b���6 e�}��IS�g��	�'>�����,���*�OL�1)�'�����G�̀��,��F]��	�'�2�3S�G�����W�'���A�'��yS4l*UNt(�i/��LX
�'q y�0oT�3�
9��R��0S�4D�`��/׏MmJMs�FL�Y;�rd&6D����BQz�0��uI^5N�%�"n8D��i�f� �6x�0)^?i�����4D�|�E��%��v�A��,�#�!�D��j�<��$�f����F%!�ď X�(u����
@�d ֩e$!��-H�[4b&n�F��.˾�!�$�[-P��Gɗ$���C�
�!�DV�U�@�$��Hi�+c�!�䝇�8�#eg�a�*Lے�r�!�D�c�Ha��R�8Ts���!�$|
U��n�\Κd��iܪJ�!�,�p"S/�]�`\��S�v3!�䗡k��ܸ�&72WM:%�ɫ�!�C(T���`K
_��!wj%�!�ě�z�8Q�䈑12�^Q�"#ՠ�!�$9���'�]mLųS���0�!�Ċ=�DH����5b9��� �L�!�$�U��bP|��DP1灠X�!��� [�|��Ʉb���s�
:~!򤈖?�̔�ql��
�X�i��#{!��1{r0���J�!�#�+7r!�!&�
	`b��{�<(!l�M7!�X~st4�$l�2B�d麡`E {!!�d/�`l��K?=����3��&`�!�� ����T%�u���h}��#"O�l�r���S&m;Q���5	�T��"O��8�c��-(:���"v ���"O6���0>H���*�\eb "O��)db���ppO�7;�"O&Q�wkHU���I�e��P"OИ��mȅT�
�q�� ��q�"O$\U�(ft88w`JI���CT"O��$c��|M:���.�&�j̀�"Od��dS�K���k&��:z<Y�"O.K�4A&ƀ����A��-6"Otm�QeȦlT\�d�}��i��"Ol|��KO�}"�* ��0*����"O�͒�
�
��+��ƙl��R�"O�Ր�G��r���B2�ːD�Iڶ"Oڝy H�����a����"O A�C�	X����ݨ;���"OƔ���m%�99S��@� e�r"OL�R�'ߖ7����C�21�*`�&"OD,3�χ)�����4+��a"O�~4HU��_!+� x�l��!��qJ|@�^�w��p�C��	�!�����Bt����ǎ��!:�"O~|���Ӵ��� �o�$K�>i��"O�E�V� =�ʭ;T�ٖM�$���"O�݈'Bʉ�٨�/ӫv L��'"O��X�└|�q�ș�����"O�i���?�V�#�f	<��� �"O�ذ�8fa֕�2嘨�|a0�"OX%���"+�4���^�l`�{�"Ov ��Ӛ�X-��Gʎ���`3"O<`���V�x-�AM���d8�R"O  4��g@� ���*��Ec "OzH�&���B<�H)"��"K��H��"O2d`C���v��1h�Q�o�Ҵj"O�a���+S�f=�2#�D@���"OR�#$:t^Tq;3"&@�Q"O>���B�G�F�ɐ�ǘce���"O��5�E�u�$\��xG�A e"O $�N&��RT��@��K�"O�9p�c�7|n�p �ȠW���"O&-:$a
�@/�:�h4�V�:"OL	�']a���8䈎-��
7"Of5
PnҴ)W�8	@gץp�� ��"O���P�-����EA�ph)��"O,Qe�a@1��R�fN1��"O���F��%
^�h���|�4��"O�3���.v��q9��Wm�pp�"OhL�d��������%�b	�"Ot ȃ�Yx@��7��4����"Ou�`�E.aKdaH��$@|5(�"O<@Q��]�!�"hB�|>��"OV���wX�q`��p:F��"O����m�8
whe���qDzт6"O9��f�~6�k3��h6N��Q"O`q�**u�H���֎]GM�!"O���b���|l��'ƍn���"O0���
�=6�����;ĞDA#"O֩p�	�>��:���-��I�0"O�I;5���y=da�K�7G��(��"Ol��7?H�<����"l��ٵ"O�h���&!C�,��T����D"OL$�%P�d4X���fr\|`p"O�`FF�+d�t�p%!V
��r"O� f�����bI��7c�88�%*"O<d � �  w*�@u,���c�"Or����!2l�P�J+P��i�"On��6.�4��}�fJؗ
�Ȍq�"O�����X�v%�D!�^�c�hp�Q"O���W�k���t���=b谅"O>�Y� m��aʃ�(��"O�$�� �+,�(DhCN)��hQC"O��K$��*2(]r%mۮn�y��"OIf*ǒ-���re����xQ"O�h"�b����a˔�*�d䨱"O�	�ue�l\D��g�MZQ"On���$mv`���ԝ ��]1�"O�}@��84�
��N�N��"O�d�ЯT���(b��%���P�"O��x$
�}�,Ӈ��>V�X���"O:����T-⴨�����;t"O�y0-A&� (�s��0R�K�"O� 3��U����wf��PSw"OX����>Q�s%�,*��PZ�"O>TAR�6�v�Z3�F�
�����"O��Q�C�kѸ�D�<r��U�D"O𹣗��������P���"O�آ�͊�,�<�kK?Iy��Qw"O=J%��b�����Rsd�8u"O�	�"ď�Ԋ]��
S�]4�*"O܀3��D���B5I*����"O��e�x�>��#BC,��p��"OZY��#��D��ٓGU�j0I�"Oȕ ��,�ȲUGS� �ju�"OrB &��#�P���I�t�B�)�"O<��ڟ$UԱ#�+Z�l�*�H�"O��6�p��I����	��i�"O�DH��ػ/�$2��n���;3"O���P�j��0c"�3�P4��"O�9 R����,@D��!^��z"O����o� x�H�K �9H@�"Ov�i��6n  r3`Z !X|�$"O�P5j�y���hVMՅB�n���"Oܨ��-�!�`9X�Ů���"!"O��@Ⴡ5 �@�V �{����"O���F��y9��[�n�"�n�(�"O��B38wN���m�G�0��"O�l�̎�Ƕ]�4�:<!ӳ"O �h���]���:v�4'��T"O�<�J��E-h=K5W�,)�"O�1Ҡl�r|�q㥫ȉ#��|ca"Oj<yђ}��!k�yՐ"OX�
��ȗWk:��&���~T,���"O�t�P�I�P�R�ݨm�va�"O�KQDЗ���y�"��v�,���"O����%?9(B4�V"�c�"OT���
��h����1"��Y��"O�胗�E�m/����	�;��i�"O^�r�J:A ���h�>!�pbB"OpU�t�N�:�d�"�I��|Ļ�"O���3�߆1h<��'� 8�2,�"O*Z��"!�D쏗|t����"O�����f>]��jȬ{�QP"O � /�zQz�"#�ĩ"�@-�"O~�zS!�.8�w�X MCr8W"O���G;Z뒘`ׇ�P0P=��"OT�J�I�+��}�b��1~ȁyP"O�s���&9�����)��t���"O� ���� �¤e�鍺i�d�*�"O���֜U��\��F�V�����"O�5�t��j���y���`� "O*9���O�|�j� �|q�C"OT�y󭍄[�R�iB��^
L9 "O�p��d��,e4Ei:/b���"O\����!��9��.{U�Ъ�"O^5����YL~�� A�QS*hy�"O�#4Ϙ1bzJ�� ���X8�q�"O�a2��#��eI��ס0+.���"O�h�g'��
i����Y�p�<,#q"O�Y��b����;�@��m�ze"O���)S��G��)$S�P�E"O��
d ),^��bOզ6��!"OܴY���$d��3$�J���"O��Cڈ�l�ע�C�Ic�"O�!�l�(Ϫ�id���Y���Z�"OHd�Ҁ�A
��;!�]@���"OJ�D�ƨg�s�Jۍo�6<;�"O�\#����s:Zl�
ϾU�`�3�"O2b�&�.��$��'�LyI�"O��;�G�:R�{��J�s�l��"O��(Ǐ	y��QsT$�� ;@��"OL��i�h�^Q��[�|!��"O"��'�0+������P$��P��"O��kcǓ4��#Ĥ�u{��[�"OX	��@�8'�\�!��S��$"O@�j�(}�(؉`��Zc�Lô"ODxˢ�6$������H".���"O�F��X��O΅�4Q��"O�x"r�A0��R	�>���h�"O�mz�	�:��Ԡ#ذ ��EA��0��a���H��U5I���ɬS�8La��9D�T"&ɛ�gڒ}iC�Bl%i��x���sӌ�qD�\�|K�5�t��3��	2�'R�O:��W�]#WHp�c�N!��ɩ"O���g����#�O�k�20��D �Şm"�����vd0���ëIǨ@��"���w��Y& �`,�p�H��'���q���S�`a(X�DJۊۨ)Q �R,�DC�ɔR��T��ϥb�`���\�QghɅȓ1��#�`�'<Y�H��@^& )�ȓ;X��IRB͹^�8�T�!RŇ�Q�H�aDg�"��]"�V%H��%�dD{����k��fh$?7���"�ٟ�y�h��`��C�$�/Ak�L�q�ۣ��	A?i�{���.	[�0�f٤Xhb��ŤN��B��|��i֜2�1xTG2c\�ɊbP�ad!�D�6@�d�ǯ��Z��u��#U�O��=%>! �
>hhT7�T0a�"�pu%D�,8�-��$�8]�2��%���8U�$���>I�y��TEN*���`���BDr��W����y�V�Q��, ��=���9S�I���'azb�F�j�e��34،ͻ�b���O����FڧJМAb���!��PЍ�<����DP�-�8@�D�]�q����	z��	A "��E���%̬)� K�Ji�C�`�:���j�Kfr�K�o�+���O�=�}� �kv��C�&x>l×�DU�<ɳ�k��]a�j��Ք��$�N�<���̐k�\diS*��#�6��Cb_G�<���	;�8<�B^��±�����<��e��@���j�B��ZA�Xb�L�<94�]H< ���#V����C�`�<� �����D�[��:D-��!����F�'9�*�5�+�6�2ݓ4�[���B�	�a]�y��ʴb�ĕ�'YwC�I�Z���!AA��ʕ`C��B�Ɍ���!�h��?PN�:%,T�WB���LU��ޜs�6�v�\� (�C��w��Jd%[�2��P�1�C�I20h�uc�ϛ�hy*�'����C�	6�����.M�$Zhp�֎��GT�C�I9m�(�9v"U�{�^@q�C�T��C�ɂO�Es�8���#EJ���C�I>qs� ��I$A�5�t`�?Mo�B�	?7��p'��p� i!��[��#=YǓm�d5�$��&t�*9��SII���ȓP����a�9���R/%f `�?�	��&�%��3�� ��W�i�,	�Ɠ^�x��	_�n���c��HS��ⵈ���'9�g�'`p���FgN���6��:?�>Q��ט'��K��M������Q=���O����N#�JUA���w����2�Џ(�!�CL�V5��4*�t����!���b���np�pϐ�c��	]��|!�eH'��Ι>K�؍YG�5���	�30<��N~a4�S�&ܵ(B#=��O`\uJs�á>_j)���P�+&���Rl`W!͙$�p9�+ fp�lZ_(<a2 ��b�j8(�G
�4왕�UQ����?����>[V��c�ʂ��%Z��FL�'��y�/ή�T�xT ; ��`Ȍ��y��':>�"F�6�<�W�Y�n������,d�D�@����(U�޿n�z�͓�0=�L<Ʉ�W>�F5�tǀlJ��3��Y��hd�x�͜4C�}S�jS(b���ʴ�ݛ�?9�'ұO?z�F�ʆ����\�y��iR�
H�'��':����H�
-���+C`X1:��@C����lZ^�tb��bMtd"s�a�̕) ���P��I�*F]%$�K�J��p��0<�L<g�±`|x\r7�Ȉx�6��$ZX~��'��ѡ�ꀔ]��P,C�Ry�x�
�~y$�Z��tPň�q�"�y@bD(rA����|<X��Vp`j5Q�&�#1��d��ɈZT�'��
q)(Nĩ����ĵ��Eè��IR����{���7A��w")��s)W��(O��=�Op�M��n^�:;���{
�'�����%M�Y�'��C��M�	�'�����nI,��/ �@Bl���'��zv�Εfʌ	p۸6�09���1�S��Þ0&,�UH�&m���,�)�yb�$oFT��δ��j�D6Ƣ=E���o�X���y'���ÆY,�^���H��$BƐC��Ӡ�N(eFP����hqaR �f(�h׌c?VQa�fX�p>�O<A��I5u��X���(�t)�C�<���(�~t�CAK���d�J�'H"=�OR�x��O
$4�-S��4f�H���V<"�P���tΌi# ?(��͆ȓl �)�Sn3lh(�I�kۺ���>	ߴ�hO�22�A�s�/|DR�Z'�^�L��C�	/0��)�]	�>)0a�J ���IC����V�K6,׃&S9#�HC5 7�]a "Oi��`�t	�W�)@�LŚ�"O�P�tUN	�e/ܚ,�TL{A�'��'}��R1�����V�l
H-�I��y�DE�֜���+a�@�x2��y
� �:��Βq��m�q��K��"O�<���ٲ:P> ����NH�S"ObY�N��)�j[���mږ"O�;�"��vLX����n�^��"O���kԱR�m�P.	�|��%�"OR����O��51��-!�9��"O&D��C�"�����b��*?ąr��Io�O�$L�/�	JWVx�K��t����'`�Q���S�ԐP���-iNd(e^��'"���3}2m�8@c\Đ&�7g�����#��y��W,(����`�
�d�����II��(O���Ą� pA�EYx������!�ArV<|�$�F
i�L�0h���^���/�2��K�'.z�ɲ`�b�4��ȓp����@�"�$h!t,[>4�݄ȓw�\�S�O����m_�ȉ�>��>�>Q�g�&б�`��8��ȓR��T�֦¿m�~l���
&���=9����D�+s���z�O���C�	��p=Y�}�	$<C��p��C*V��AU�?�	�'S��@DbS.~�6���.��l_�H2O��"�]i�S�'2�
-��(�
@�<qp牊e���ȓ7~��٣O��Z@� o��j��>A�ÁV}R�I�:����1_�ĳ'N?H�C�I�qb�h�0,Ѿ!bܥR�M]��"�'�\-�@A���y��.�� �V���'�2%䊃.pSa�� 1�'3�Y�An�>"�}KE*��tݢ
�'UL����-B�t&�"	F��K�'!��+���3L��$���-Ԩ��'H��B!���f�ش�� �<u��'�R(�$�.�Hx�ė�{N`��'[�D����v\0��lŬt�dP��'�v0�Ac�uZ�;�NT�j��0��'�`h�pbvL��*��6E.��'-(���'��un�
�lU�('
L��'�<aْL����|*A�ZL�n��
�'N6Ԙ�F�5�9
P�a��@
�'<ؔX��0?��q���4=�$T�	�'΄š�L�X!��{�M��Dt���'�ayS�ǨG�JA��DD L@�'�Ĭaq���G׬��w��#L���R
�'	h����]����ǰ�Z�	�'m�h�Ŝ�h8��c��6�`��'�Br���:���aV��$b�,� �',`�au釞
n�Zv��e����'�%W�D�H��q+��γFCD%��'^����ъ2 >�8�*p���k�'�����ş�j�L!�'P�r,��'z�#��H�MB��B�&�����'t��(�gJgL\8���-BZ��'?x,a���J|�EhGi�x����
�' ��9��B��0�V��#�y��'��h2i�-�2��gkI��`��',`����3#����(�). ��'��{sAӦM�~�j7�W6}�����',���2�!�.�1}�*��'�4$��Ռ(|��ɬ]�p y�'�d2a��	OD���U<Y���x	�'Ǯ����+ Ø��@N�S�R�p
�'��]�P-�2�>i��C���ǘ/�yRHu8<����� ��DQBi���y"'Hb�B���c�0@ "�.�y�o��$��N>d��0kG-��'��=H����q�(h��S�)�z�;�y
� P�T!�R�*y�FAN�+�H<�*O��i"#@�B����C;b��t��'-�*�#̇K+��`AK�"���'�4�@��F�d��0h@�ӑ�R�B�'P�I1��#e�䣒#��|�����'�ֽ9׫Et���²�\j�T��'li���ϗS(��c�ą�Yf
�+�'<�tB�D�-U��|�H�j� ܩ
�'����Y;!{�%�Cd��e �'D�IR�Q�$�S�ͽ6<��	�'}�mp�������#Ԥ"|���'Bb�s�,�7IA���e
�#�8 �'�8��֡Z�]�C���'�^
�'����¢�c:F�3��F;�)�'���&�7i������4< }�
�'�v��V��%�h��A�YC
�'�z�@�o�,;S  bT��*a�4<*	�'ĶY�6� !� 0P���-����'yJaX�R���Wh�)$ܰ�K�'J8daǌ^�H�X�X �U��6�c
�'��¶N�P�B�0���
���a
�'O��r��V%id:a���x�%D��I��)�\�x`�;V��U�4D��S'��L¼#��M�҉a�b4D���mU�a��h���0�dp�c�>D� s��U!�6T��� !��CR�<D�x$Ǚ%@B�s��&WÄ��r.D��e�;<�j�k�W���1l/D��Q���"�0s���o�����+D��;�M�m���8[<*xY"+D��k����ms\�!@����(g&D��c	4�ze��K�SǨ�I��%D�x2�oٵm8��c2b�#`?���P� D��h�����-�gGװ����:D�h��F>(�)(e� J��qb�n,D�0��"V/2�V�C`�"�Љ��"&D���֪'��U07�ɫ eTMM�<Iâ{N�(�E^&CKD@���H�<�R���^8 ���� �qmUQ�<y�1P�&�
E��5'5.Ȋb��N�<��g~f�pZ��U7N���R��b�<A ����n�'aW��&$�b�F��L�5l�˰\�'�r{R�[�\5��9�/��`5�	��'!D�0�E�(&غ]��@-7h��ʎy� �5m���V�L�O���(�Ǜ!\L��ܬ8YxS�"OpD� mH5	,�X'&Q��2�bFՊ@��Q���J�|�g����>�0�t�ϴEf����Bס�$.��ER j�=#!�P�ïؼ=Ub���i�& ���Rb-�O.�8��C�~|��.I��I��'�t`�Ae�-O��a�:ON�"c��U��	�1. xb"OZ��
�6��%��MPb 4�0�|��g*�j��Ę=�?Q;#@
�x��4���R�k,D��9�#��ML}�d]�(�@�53:Ё���<!� ����m�&�J�b���RB�G<8�B�I����k$�H�9{X�@e�؝3'ب����C�����N���&��(}�xb��#D�h�l)<O�pJ��E� C�@�Li��Q�i�D�~���f�L���ac@%D�ܐ��'Y���${����&�Iz ���GD�h�Q?�vΈ�K��ʓ�߄{�t9�VE#D�D��fC�0�qs���)� �z�H�{o2��H>q� �gyBW	8^n|�Ef�o�V�z D6�y"��	�T<`l��T��$CH2�yR�I�aB� �Ԏ�
c����˱�yB���|���R��t�X��y
� �a��/e�4A��)t�BX�U"O^jB����<�:�l^4=7f��"O��9t��QnЙr�<8U�2"Or�{b$.ELt��798���"OX-).	&^y���ΫU�c`"OLa �m�`[*I��':�$]�"OV��i¾p�t�Q�*r�nYb�"OB�e
�f�| t����J�"O�%t�?��T#��X�J�S&"O�t��c�A��%h��ƛP!���e"O@�AD�bTt䳧B܀�u"O^�S��W�b-dDsBQ?�\�9��>��f����S@)�82���aM��ˆBΞ)��"O*����3|��b��ưg�V�8��Nnb˓���rc\K�g�$�|E8G�QH�B2��gѴ=���#%�pY���P3�`�e���T����ǫ�m��19E�N\�a}���C����Ɗ�>nq6��dܭ��O
�fǚ)_����В����'l�zh�����,9�Хl5!�dP�~H�Lޏ.�V�C�4C�	�{8�;�N���!��S)�6aQeԟDXA#��.|C�I�.����!�!��eI��/`.��@"ͮ�~(,N^MQ����{2aؠq�=y5�O��0 Sc����?�g�X�w.غ��6Aa�`dfG*Zs��ˆ`��A+D��Gdr���{��i�>C��J���G���᧪����$ήV�c���+Ԃv�q����������1A��
?.�ܣd��&�س$�P���c>c���?R%�%�1�M+!���a��<�� ��6���Sk�l��	6<h�Aԟ��w����'n��Y'T��4p��`5lX@y�ד[n�0m{�N�)�5E�d�vJAd� #A�!-���Rv�(*����T��k��(9X�H�8��Ԡ{d�C���⌠���d�A�0�{RA�"l�ix��۸p�:]ðH�B!��ᙅr۶�4	�lp�'��R�d6§1H���SҲ]���!0@/J�����;�6���Oa��ѲČL���I"���Po�AA�MB({P~���'�` �I�F�0��ǥ�{F{�Y"�� ;��0[�H��m�>�ēf����V�[^�����]C`�����_��f��6p�ey��Y�>����fkKi
��B#�'�j}��'66}�'�ę���6�݄�XTa##3}��D�;����'L��x���X�F�o�0]���/~;F���G�YŀEpH��>�p��D��}1^H��ӨM~h�1B/҆R0�r�m��(��D�ם&�,qeCA��M�o�&S����D\� `��pbl� Q��h�c(Z�џ�QÃ�2~PR���$ə hp�����&]:u�s+�J�2��$�j=b�&?��	�$�	�{s\�)@-^|�
fύK\��P�P�1��?2*ӧ�ԊX9<:Y�c�o�:1�AaI4�����1��U��&/�xb�n!�q��A�8&ʄ95B��'�$����uk�`Y��D������!�l��$�ΞK���BKur��W�#�b�C�	8
���2�ڇz�LI�!��w�\�� 
�8��'�Z����i�Zh!g���x�&a�=CO�rÓ+\؈�@���h��8�&��gq4� M�"�ʼ�ȓX ;d�x��m�Ө�p#$��On˖�љ����O�Z�HTh٭C(6�5��/R(��'~ 5p �N�LI*�p�/đR���	�'u��� �%�p�!A���#�
1	�'�^`Se�˵a9�m�'�ۊ,7�@��S�,�d�V�B��q��=�V��ȓP�С{�aF� Ī�Տ�2H%�(�ȓ欪�.TQ�	kC�D�)O��Dy�$��	�F��H�6���sS�c�2�O��yr��O\BlƧ��D|1T�P�[�4Xє�ė`}ɧ���DY�P�M���&_n��[��(-�!�d�?lD~��6l��rTƎ"�R�W8h�ؽ� ʐk؞�!a�Ć@o\Q�"аu�ٱ��5lO�	:v��0>\,��c�i��Pj��K_�УtC�gZܫ)O,y�S�����=�GL�K�H2A͒�:R@ؒ�/Sܓ)"fQ�7?d��I�O�Њ�Oۓy�Е�䄌:(�b���V^�i�r�L�<	GB�y�`Ly�i�,l�;�*�t.��I��d�Wr���=K3���,�XUЙw ,�97�H�"�0��R&�h������� .QQ"�Ʋ���S�$�5���$�R�%pt�@OY;"JnPS�J�.YyR�Ǳ��������^�qC�(@�P��f��D��Z<�
��� `6mŎN}�{6�G:d�~9:¡̋l���Ot���p��^.DB0�a��'݀󒯙�o2�x��X/��-��{bW�[��v�ؖ}���#>�vu��o ��?�e/��" ����s/P�Kb�ͽ\�����F �	��ɯ@���F��>!��+$AS�����'�;"�:�?AAII.B����'R���/~f��p7��W����ߑp��C� -��h����x����7bV��h��p�p���H͜C#8jƕ�-��P�iz����cy�]�]Z<)�M@	W>4�BM5Ȱ=!ac�$�X��i��<�HE�Ht�[��Ĭi�*u蔴~�L��'$��S#^�Ҧ�ɭP�L�?����!I�رP(Z�0'�3���Pyr�¡i7Ƙ8'�Ȏ2A|�����6q&��̋vȔ�H��)z���V�1? �b!p���%R����f�'�O��5����q��.�-����Y���fi�9A1����N$>5t�	�`��i�(�#$��;G���4��pa�%�%ق���JӰs�<���ܦMx�x�O��z� Ţ$/ 6^�̰�c��n����ѯL�H���
:�2��/��	�(<z�'ʊ��į�.��ԉU(+����䘨N�.P `�0��d@�g�"��,�)0�굠 ���9�4���� �h�B��	Ĵ�cJB�C�FR��6;���g#ٻp�{P�1�~�W<��h�c^CyB�^�f,c� �~�h6�M�iq�A�F�b�6�q��ɛQ�wը���c��3�Ѱ3�Z���L��<�Fd�'e6�ڥ�uv���� M8}�P *&��*]�Uq7g�����n��Ԙ�O�S��I���_�p?��'��OdN0	��"��b�-��3p�غ��� A�
lk�u��!#'�-[J:TI �<@E �'����an�����p�g�'V�8R�����|����8(Pv�H�"�qC�i�V��=G��/�^�+�.�=Ѭ���ɜv�>equ,/�,Y��_�r\��ɫb�T�@���-��Sr�	.�8����O�}��=� d�.)/�0�2$�p���E+X��Px��׵w0��zwT�w&,+���h�Xpd�V
;Z��6�ǻ[����S�V��'^H�9�Ѥ�E� C �%}�<���	*_J�1�®ܮL���{�.�u_jd�$G�(�����ؾQ�v�r�U��G���;q��x���'��-�I�1oH��ȓM#��9A'̟u���P�3.����'}��k�3 Ȱ(��	�'ĬM�ְ�����Lx����*N~�mA"l�0��\�@¸����)3�K	�'��:�"�7�����N>"C���X�WB^��3��`�r�P6�Y�a.f�C��ծN>fC�ɱ( ���t�C_�nj�l� �ɦb.�d��ӸK
�$`�ķF���0�,�1$������y	`n݊e (HTƚ�!�
(%6������_�B$R�F�D2!�d���B�m��B���pe.�#!�$A6�杸t����)y��X?{!��D][�E��J�J���'�!��t+䖄`�+Ƒb��[����!��Ҭ>l��"`�3|��)x��ڠH�!��$w��i���)���A�ȝ:V!�dK9W�` #2OMڴ�@�A�EZ!����X�I@+�V���A$����!������SoGI�z��Q��u��'f�� cK�_+*�ɀ�S!�4���'���;AX)
�^�р�ۻ!΀���'&N�bq(�<1�ԅ�mS	r%����'PL��b%�9\�,4��jRs�4�9�'��
VK��|x��u�U/hz�a��'��1��$(���
n>0 q�'"9��-Ԟg%�0�B���
wi�i�<�eЮ5̆�c�&��}]N\�E"h�<��b�. G�Jlʔbй���g�<rH�]9�D���B(/Ќ����\�<��bA7�Dl�-�'IS�y'��_�<�e�<ܒ5U8�,9w��r�<ѓ+� �5P	�?�B#�o�<�@�I�P�J�*&��ɑ+�k�<y�fN>Ĭ$��a]Ȑ�f�d�<�� >y`��Dm�.�P%!"�`�<� ���pm�J���iJ�OK�U�V"O��3#n�25��	O�E:Z�0�"O~9�Ц^�:ۘ]���9���v"O(iY�.%4���钌_bl�g"O(��W�A''\� wG�7iV�!"OJ��#���1��<R�FֆHdP��"O��@�Y�|�ޥ��lB/(�^iP�"O� q�o��<b:�R��9YB���"O�H� Ri��hC1LJ�G�t��"O!��#M�dih��d��"O�X�R"O�Q�i�S���K�	X�2�.az�"O�D*p��g.4�g�2�D5�!"OB=�¡ѧ]�zLr��)q��`K�"O��j��c�H�@�%ؑ-�"O`s��b�(d;a��̴Ua�"O�0�vl՛	� $RdL�=KE�m��"O ���d�8��%?�@�"OʔjE�PD0���і7����T"OL���#�${�DH�Ph�:}���@0"OLlu�O}�4��w	�Of(��"O�Q�Ĕ�"�kƏ�;��`�"O�4�P��Xj�q�J�xۣ"O����OG��0"�L��~T�Xғ"OFhQE��Y�8��fi_�1~t;�"O������[�"@��häU'"\i"O��YAH0E��9� �8U�l�"�"O��c��V{�EJC-ԇ(&���"OTՑB �$u���3L0X�S�"O��Ud�/t�XI�kCW&&m#�"O\��܏ˈ��iX.J�AI6"O��֣�1jPH�Tm���"�2&"O�ؓ
�R�%�W�����t"ODm��m̕<�e��oT#r�P��"OЀd#�#zt��R��<����'шa�'��\��tqDh�Um��'�pQ���Q;e8�@H8FîA�' ���e�.>&6�����?�� ��';�(Y��˘G���r�H�FV�	2	�'�0HUL@f��%��W
���	�'=�= �g[dnX)�I�C�#�'A�r���^t�%@�T;�lP�'C��83�
 ��i:�G*I�h��'9��a���n�0�A��L�@��'����1N��U88���BM#:����'\�La��-��<��DY_PL�	�'yt�ҵ �<MH`��L�n��i�דZ00b�?����"WǤE+EBS�dS�m����3,�!�$��[`��*$Kҋ @�����s�1O��ȧ���q�j�����I����B$M.uO��"T Htr!�$wJ�HyR��	_��9���jLMI��ȕ&4�IY�:���OJ��f�TX�@���%K����O($ㆦ��.8pWb�@p� ���H3m`�U`��t!���� I����2x�}��E�!~9�y2)3}�M�'A�|;��@ [�t@��olmH#f�C�N���ȓ[�)��5X���9���	�\$�������B$����[�O����D¬5�>y��/�px@��'b�ph�έYt$Aok~�"�&� ��Ȋ-O��a�9�3}�k�^D�@*�m �l�rXvK��x�K��-�]��N�y����*�{���2aZ7�$E�G�'�ޭC�R=f�H)�R�2@�ϓf�P�_Q�8H��'�*�뎱�x�p��G@ɉ�'��yQ��v#�tk0�P�8R�q��y"�P:W�e�v.P�O�(��'�)5�q��i�g���'�p�z@�'����әs5.]�uN���.�O,U���Y�� ,����_'0�Ԝ�(ԧk�&�JG"O
�bF�׬'}��K�%C7ߤM�`"O1��	�W� #�D�zV�E�$"O�\�rm/����$�$Lx�"O�])��<=���`���z?��0�"O��"�nj��v�������Sf�<���.S���NJ�P�S'��I�<��Q�N$����\1m������K�<��P�ZCZ�{��vU�I�g�Ql�<��ώk��)�՛QK&��`�<A-͊
�� �Ο/V��ٴɌI�<A�	�y������
�@tH���J�<�w�Q3F\V}�1ٍF8���A�B�<9�Y"Y�x=z�kEY}�9���~�<���U#:��q�v�Xq6h|f�v�<�s�q�x����ڈA�J�8�Eo����l�(Q���0|Ғa	��BɅ3��D  �j�<9��^�4��=�1�L��$����,aI�@+OL�T�O5D�1�1OPd�bɐ)��s𬃩u�����'�Tp��^=�� �1.	��J@���/Q2��s���1斄����9Ny�T���~�^u���I�ͬ�?��R�7��F�y�%ɱS?�UH��a�r�֬ܯI��)�o2D��3D�T���*TI�vz��	�<PK�'_$��᳌ɤO�#"�dy
FF�*��YwgF�<9�C����A4�.`� !���*T2���@�Or㥈�;LH��qO�)��.�JUQ�I��L��pIf�'��5��� �,g�4 ��V�]u�Lhh�=U0��J E�b��u'N�7�qOVb?yX��[ޔ�R���
#��2T�>��o|X���3 �k���~*��Ow���"kOP-��!����P/�	�KB�g�1��,8��2d{�lI&��=�8��'ʔ����Y<�v���
q�O�� �à�Xxl . ���礝U�>��IP[}h��IZ�⩚@e�,e��e���N��n�j}���3ǔh�O�\U���EͲa�O�y�N
U
�i��֗0 <���(?�O�m ��y�驅��7��Ssi���
�s�������4� �3Ӊ����a�O��]��/:H*T�T�4���Vd�h��I,��'l��q�n��.�h�q0)E��b���'��9�"���F��inF{,^P�6�r�)��/�
��$N	��'+ �J$��9���?5�S�?!�����$B���+H?�z�yC�7A�|B*A;�?�!�=1����J�����IZ%l�&>���4L�8��g�PpL)� �s�6@�69�6�(G�*}EP�@6j��rΨ�'�'�<�x���d��+���8l> u{��_0M���r�*�ݷ��%q�xӸy& ��<1Ǡ+�\�bG�$D
��]�'"��#�k�vVd$>ٙ1	��-����f$�1)2ޭ�7��ݟ���-�>hM�1�RC�+}���E�(D> ���dj��j@0��F� 2���(	�1�dB[����?	��ڛ2�Ǐ6fT�J�A� ���YA�V-��<dVC���-r�ys�$��q��k��+Δ��J��1�J�6k_�-)��ζlk�O�c�wcT��?7�ΑS҂*���	�a^�;�\�K�L�
BB�6���2!3��Պ���"'�c�ܒT�4���&Z+T�nx`0��5�>�Q��0OX��%cC�3n�c�H�6��	c�~�B.�ԣ�"O4u6&�/��qW�����2c�>��B9]!D��?% W �"��Ȑ���P��1ӆ@=D��U��[��9 �R�v�J��G�<D� �u#ν<<�뤆�6yW|U�:D�H��@D�#i@E���6D�ܪ��ۨO���
�-�Qs�5D�nm�6��|k��ȓ|jt�p�/D���P���#�����M�,�x��-�ܨ�p� �'4y2͒̒<��jwF nr��ȓ�r���î:���It� =`��ñ���E2�K>E��'X�9�d�"j.�YSd�;{��}��'����u�ĸ�t��Ճ#@,�I�_�B�CQ�Ǎ_?����Fa���G@�<ɨ������l؞�YM�0<����kӀ�1�E��{Dx�1K��BDZDH�"O� ��"�{��y�����<���d��UR%�Wg��Z9�"}Z#�΄N��J�iVY����(A�<�R��o����'�em&�rLP>.O����ώ)Lx�I1C�Q>�BlM#C-X�	�\��� "�F��ȓ P��)�2%��=ذ�	�p .�k ����3��a{R.V�u,�<`���0�s�X"�p=�_
���sH\��Mk�I���^%�J�8n��9��u�<�Q%��.:ܵ9R�|@F�
��s�!�B-��N�)_F|ى���	b�Z(�򊅞k���J3)��$!��EUj	
�c��t�2���n�6l@����:��l�>�|�'�5
hpx�
?u�ui�'xd����"v��i���j�B`��g-HR=Zǩ��0>��F�f�$��-͢0k���N`؞�ITƍ�c�����Ua���jXt��d�5H�,Y,���3�����[�WG��*��H(�}�'�Z���X:#�\l@׉LE�O�ey���|�@�̖�I0p�	�'CV�+�l�PɁ�ǭk!Z�zI<���WY�J��Ǔz�D��@�H�uG� ��6GL0,��I�*��V)�'�;-�N��"�֞sDLA�Ot٘�f �a�P�`vMRxU���	�;mhH�
�d�1���D�:)�ly#nFE�D"O!�5/�-V���sC2*���d�O�x���5�E�H�b>��D㑂^�j=8����c�b�'�]�@�A0�"Oh��W�muP[�&����Q �k��Q�b��D��D?��$��S�MиهL�J��"H��0\<��dL�_N!Ca�jFl��#,*���0��(T�FdF/>�ܸ�Q�!}r�ӵ~�����&]����"e�tE}r��"�I�e@J�'}!"���2Wd�"aK��T�'D�Da0�
�)�~\��II�&��
��^ (Η�)<0��0V�� �R� 0q��S��gTlP��I�0�,5Pt���cI1h�##O%{�#��8L���`6�3�ēi�`�#6#��q�9+���2D�O�	V5����Aڸ�NE��U��2K�4�jؠG
�I�Ɓ��ߗ{�q1��js������U��u�O?Ź'@R�#� ��d�N%�t|�a�Pk�<15�E�¥itC��V �+�J�my�&Q%$NM��/DjX�����֘3d��JY�����h5�O����U;lLd%@��W��i�,�R�^��c܂��x���Aa�13��Ϗ]k��+��¦��O��Ce�L>d�?�ӄ@�YB
�K'��@?�q&�*D� Q�Kr:�ДK�$e��K�̫�X��i�-YqO�>��lλAd�Lx �ϑ|�l5b��2D�X�V ��K[�}�Ӂ�>X����3D� ��#!�\2l�$,�B�Zf�:D���v�^�N@P�پ1tp��@7D���KZ7-8YaCԎ-�~|A� D�Dj���K�Qc��U��A�1�3D��X`MK	F�(� �)$\�i��1D��0���Oy�Xا-U2�f�as�,D�@IIʩ>b0	A ��B=�	+D�z$�^��	Ҫw�Ƒp�<D�!���&B���T��
p�e�4D�ѷa'N��Ԑ�Q�[炠��C2D���1c�w�����&�-b�iYF�2D�\1���i��4�r#�X�S�0D�@���N�R�n�4̉)@_� @�1D��{�o��"4<(����<������:D�d��[�S�8ze���Ylڭ@"�'D� ������ݪ'�ĥD��}�'�6D�H�2��(�81����#8�Yc�3D�IQǉ&X��)�lA��dm��#0D�`Z�M�f�ư�I=�D�Zv�/D�`QfM�k���1g�ڑ�J�s�.'D��c�l�8I�v(\�P�m)D���d����1�C\�.�ڀz2":D�� "��P��aF0(7���]v�B�"O�a��J�R^��K�C�F�c�"O�Q�
�?L�Ԉ��^�/M�a"O�2�,��\:�5������x�"O���'�Á��b`L	b�L���"O40�`J�*���a��� ����"O�Rf� :cM|�#�#�-I�@9A"O�]2׃_H� Hq��B���%�d�9E���� �T�n�u���1O�
gC*N�0��J�/�  ��"O��y�O��H|ekr#�u�Hq@V"O^��		o�Q9�b��� e�R"O��TFP��rT�}�"<q�"OAH��+���'/�]9J(H�"O�u���\Љb��T5dY�E"OȝX�֨>ҼE�c�V�1��4�&"O��u�Ͳ�J�;�萑E{"iq"O�;v
��tf����c�s�"O�S!?��W��+PV�D"�"ON�ɑNÙ(����>c�"d�"O�qJ�T*zY6- ���,a�z�(��'.�*׹i�h�a�	��&n@Q `A�	?�>�Ӌ{2��z��O�OĒ���n�S���Ӏ�t�%ǁ���3q�
�}���F�,.I2Wǁ 
.����3o�����Фst�'���I3,�`��!I;Q&F���ҜD\v5ˢ*V:��$\�Kru����l5��+�$�$�Q�j�2<��Q^�̚`fI*A���
ç.>"�r�܈
^��q�� ��=��mO���'W*���K��Q9U]�����]]LeY�Y���Sť��t�r
��u�dMc�OԨ��`���7Á/*�P;�a�j~�Oƃ_U2ĩf�Oj~m���L�7S��c�#H��f��(O�H�&�� �X��!��b>W�O��:K�e.`� #A+H�� G�'�V(Y&�B�	3�ڐd�>E��C��2����Ƅh�M7Ş��M@ƞ8Ԝ�M1	��{v�� 2$����D x6�u�Vi�R�\=M���I�!�gRR�̓����Oaz�]�{z@����^�p��$�	�'8�E�2$�#ۺa���d���	�'V$m؄i�A�衡�R�D�\���'&�E	V�悝����@!�P�'s@�C�Ή�s5"E!��	 k����'���)�끁lc~L�2��(j��i!�'4d9��K�e�iu��_h�	�'s���AL<�Z!��-�7J\���'��k��A�7*�M�ÁY �J�2	�'O�p���4F\$i!�E߰^�ε��'�����9>!��D��V���'O0�����!t$���]z �A�'�.e� .%1���'q
~E��'bl�`� �=�B\k��Z�!�{�'-\8x6M��(,���I1���)�'�LL��
�;���O��N���'՞9�	տ��̑��J9=m0��
����,	�%��K��_�44
NZ�yr�V����mƫB�RP�,A��yb.�+�0��4C
�8���	R���y�(J	m���S�\#'�6%1�*ϛ�y��9$�"���]�&Y�YQ���y.S+z�xq��#r�H2j���y�R-$LLxڅ`��f���$I$�y2�&Y�
-��R�\���Q��y�0m�v�`/cI�G`�)t�xy�ȓ:�l�)V��1V���딭ؤz��t�ȓa䰓�fF�k�����J����ȓP�*ܰ�Hϖ$�5dN�/Ҩ4�ȓb�Ē&#�EÜ��2FL�]]@���l���@��3Vh�[e�Z�>��?�@8е�oѲL��.S�e��S�? �@h�BT�pz5@�aN�KpH��"O�ic�iF�{KF��Q #s��C�"O�4�"���U-��rR쀃�"O�D��,��)u���.��c"O��P��O�UɺLq�GO's��'"O|�0�Q�M��u �e�]�h�� "Oʝ��4�n8U$ǣ[�ɫ "O�`�@U��n�2�bP���P�"Oڀ�Q��/��U��2<����Q"O�|jQG�!1~*��A[��V��"O��R�J�/ ���#!�Ry��"O�P1# ֍�3�1�(�`"Oе+Qx��Ҧ�V����"O4q�bT:
(1��� /�n\i&"O �J�bY�a�<S� I�J�4�"Oh��b^�A�(ha �{�=#�"O k�o˒SD�#�dO�T��@v"O�#��=@�m�De�"0PH:&*OȰZ�BD���Q�R���	�'��	�\�w�!�n��b%�@r
�'��p��O��m��`񩀆\%n��
�'���K$��$.�*��l� \����
�'��ũ��Ըp���`�܆A%l��'�\�`���&I�p��?*����'a��2G�طiQ�l��+�,p0X�3�'S����㖡t1��̎ur����'�fAi�����,ġg%
y��'����6L�p�ҥ�M5�R�'�ȝ��j0�2A�eE��
��'��<��f��+�B]�da�'yHX"�'
P2d�Y��C�,Y{)R�A�'=�����D�>�A��Pz� �
�'�ͺ�*ܟOg֭��;D�N̲	�'׌�X M���@ZQ�@*?�J0c	�'��
Ηa�h1�󡖊0���J
�'x���� E(�@�&@�� â1a�'�D��n1 ��a��� \-J�'�"�Ò�_��>	��/l�<�
�'�ʰ����jz�yƬ7"��'����L]-�j� ��©��<h�'�q2�)ا|�E
4F�g> 1c�'C�I��c؀��i�[�q�
l��'h��7�Q;HQ�a�˜Y�Rx��'�@�q���c9�b��]�"Ƹk�'�aY#�ġ/xd�"A̭+;0 ��' 6�Чg�8K4�t���)r@ɪ�'���#��̷��݃G�@�J�'d֝�a�V�"S���f ԾY���a	�'�:�f�.�0I�ŏ�P���	�'O���࢚8Ǆu ����wq��'8ԉPV<\�r�#Z�D�L��'],`�Ɖ�d�me͝�9D^���'�", �ԷYUT5qg�Z�/:�1`�'6��gׅII����뒑Bf�
�'��uI98Np��s���!Ep��
�'�H�1�1Z�����̘�c|F�
�'S��&ed������/^��R�'�H�B��:�ԨSm�%&�����'��� #�M�5���HR�Ƕy��'�^�#���!%Z�x��.�JH�J
�'[H�(G#בh�:��W"y�H0�',y;�C�%~��uh"�hT	p�'���!��C)z��J��+]�0��'�69�f���=��I�ǝPꐘ��S�? 2铤�'ʢ�ȵ��� �<�I%"O(h@ �ՠ �Τ�A��J���0"Ō
$�X�I�!&B~Gj�"O����Ή9�t��"J�T�A��"O�8Ʌ�I�<���!ćE,�Cw"O6�	p�^�x�ִ���L71�l§"OR��Gf�
k�̬��hT7d�
�C"O�pQ��\��l{���2O��̣�"O�cU��,�S����.Xx�"O�|��jD� �r���`)k�tyi"O�@����5f�y�S/���a�"O`I��l�(NS�E�
(2T�@"O|�! ��i�eQu!X�	ܨk�"O�^r�Pѣ\6b2�H��!�D�Z>m��Oơ�2����$!�d��F�ig��#c�5��"�K�!�!��\z$��>g҈9�q�é1�!�dޖnH�@AK7W#�p���^�!�
��̩�	΋nZE2�	*w�!�Dң,�P)i�eX��-���J']�!��;>��I
u
��{��#F��E�!�;4G�PQ�C�\`
�$�72�!�S6\|\�x�#"� ad-4V�!��ߐ2mFAbgĊ �v��FMM03T!�䂿X���8p��,k\�pa͉!E!�dЗX;��q� �;L��E
�&#!�dHB��Hyw�� �i���;a!�:oKT�`�@�G�a0�ȉ�cI!���h.���D��M+����a�D2!�dG�r{2�蔩ޓ*��0�֟|*!��-$~���펇&��q��͗.!�D�1S�8y`�
��L�r�_�]f!�Dx����/�T��1Ü� !�da�P��v��2�z"L8b�!�dZ�N��U���V�%+S�T6Y�!��Ƞ���hY�g�eCP̔�(�!��̋s,��z��K�M�@��F��PyҮȊO��1�c,�+4m괂��y����PĜ��V��-n��ԡ��yb X",��a�u����a�%L��yR�*C,�{AI�)p@���;�y2D���1Ӣ�՞4�Ʊ��(�#�y�� :¸�ԭ�ΐ�C,L6�y��);�񫡢�{~�0����yrHC�5 �r3�A�`��1���y˔����uMX��٠�y"�hpl�ː��a!؂F�>�y�I] *l�AC,Ə\ V 
��P��y���"��(r��׵Y�⨙��� �y��¢)��Po�Y�0B�̝3�y�ۮBs�kA��y\n�dDL�yb.@�Z����vfV�q��]��a �y���9e�T�I�d�v����6MЦ�y2%-d~ꨂ��L1Pd���۫�yb@
�T��`+dC�xߔi��e���y�
!Ԛ��uk�&s�TM[c�*�y�Om�P�(� ۬!�V�yA���y��W�c�j���%�E�.���oM(�y"dģ+dr��aÁ�̄c�I��y�eA�/��<�Vc�'�hY�]��y2b��!��T���	�xh�������y��&c�NE8�@ �r��U{�B˳�y�O֫D8�A�íkc>�Ɂ�D��yR�Ro']�&�D�rV�31��y
� $0v�@�T���SA.]C/Й��"O-c�6i�Jջĭ[(5�H��"OR����ϘQ�r�ѫ�6�D�F"O���4�K�k`����S1S����"O�`[f�C�?�@�	�,$����"OH�p�����(��a��J&"O��(���(B���t'@�EW�I�"O$��.@r���� �B���5"O���u��x�m�3D�[�"O�$"�a� jC����o�-\$X�"OĀ�tIT�Cv������`���"O�I��>4Jb�` ��m�|���"O��G@�r[|���	���y�"O8���Y�P���2 �_�*���"OT���D�QB�9�O,Os�"O�ȗ�V)Y�](�D�Y�Mj�"O�|�����Rp�)rS��WMır�"O� AVF 8�V��l?Z���"O�P2�ǌ'�6����'%�Q�"O�ɺ$�� 9�l@���D	��y�"On�!�O��^n<��f��=M��V"O�x��΄�Gǖ�!@�d��=Q"OؠYC�4F�v�#�dN?���0F"O��`�'U�N���ㆡ�@eb�"O2�Z������a��Ce�j�J2"O���+��j�By���,`�bp{�"O�C��e3��aw�%X�V	JR�6D��*4��z���IS�0�X�F4D�̰U.�*HNt���ܖ'��$�1D�li�l�)�$L���V�E>8�UA;D������]#>Lё+�,t��`�e-D��*bO�� ]�R�P�?H� c�(D��3�N߮���Q�2	�!6�!D��"��Q}��q3�p��|`P�<D��S���u4�Qa�"Gx����#9D�\�҅S�[���,*6n��T$8D��[�Э
d�z��Æp!h6�5D��0�N   �