MPQ    4�    h�  h                                                                                 �C=W������՘��w^�eO��p _6���P�9���� �EP �n��q&Z�=����^��o�
?B�[�j 9��1$�CSd�0&�����G�I�#pa����f�?"�F/Q9%���w+���	X����� ���_m�d�8���w���=Z��1`ǻ�=�z�U���h塶d��JL�Ņ�F�s��~@h0:m�4i�	���x�r�N�5 Z ˌk}���3�ٜOG�ܜk�0�XlqJ����=P�t���׸���R���o`f��Ot��%�`��w�XaVx%{J��#$2�[M�j���>��D��Hd;)��ꈎ���3ΥS|h���A�Z�Е$G���)*���VT�8KH'yT-�7�a���͟&u��".=��ݩ��~�a3�ڕ#	��}6�O)@\*����+� މ9~��<��R�g/^��}�����f�V�����]Xɯ�N�wݺ��ss
1ε[y��h.��5m�bk���|^�;��X��+#N�I�L�;�b��ǒr����#?�&%�S�_l~K��h�	�L�*5��
�Ls�O��j�����i�����L*n��mE*�X�v�Tuo��f�X�*�4û�a�����J�%qy��z�`�L������D�s%��
˯�c��ǅ���'cv�z�K�����e��M��χ�T!����0Q��,����y���qᐙ��XEf�z�"m�kQ�P��{d��`!�- ��.���*}�@���;�]��1 RY�؎�9�=yvq[:�)�*r��6cj�ҋ�U�s��Q�}�I��#k�S>���U��)ܨ���o���
a���ep���_ƹ��+�5H�M�*\6f� ��3�&KkX����ధd����K���)p4!���Cw�GB��F�!�<��(VWZ�U9_���-��H�v7T�0�tF��n��������>����
�H*C�j��pt̸l0� �(#�(!\�����Z���i)�?�M��m�w��/�T7���m�� ?3S꣞m�����Ї�Mbچ�D��(����-M�B-}JO�0��_��t�ٰ���pRs�DLW����@�ȱ�O��6�-�Z\|�����K燌�E�m��Fa_���PDQ��p��*t�u/���w#U�h��dd���9`ݱ�hί�7G#�7aZI=�;�K'F�S߯$��ef<T<����\�-���#���7��e�")�Ɛp�up�g����ϡq-��@Ѐ�<����c�	�r�Áh�y�2>0vn2Zޥag�F�쪦�1b��"T�,]�[�0ϗ�<���km�Z�W[b�V���Y�M ��k�&ʣ�XID���LI`��{Naߙ�Yp/�{5��N��b
s5�9���כ+쏻��q绤�A�z�0o�4)�Xr�EB繥�:�e�v�D�%��CvL�{�4$�}$��'��<�[��19T��1�DS@�/&2����}�5�R�ngM�|I�5��$�!XݼWGOa4��6J�j˿�k����N��i���1�S��õ�8��{]s�0�3;��H2	���+S����n���e �&���?�!�Y9���90H)c[�}Ri��F�i��A!깆&���_�����+�1����oJ����[4R�Uk"�/�n�i�)y��n��fU(_ح���e����K�y����Uۡ��6o��=³���H�/T`˾��=��e�*,xk��t�vN�^���׹�5ې�N��X�j&�ٙ�[�7�~��2�o�J��d���5F	ϸ-lx����,G%~B��Kgօ�G��)��+��j�=��_Po�&Lv��R7�w>��gM���s���Bg[�q��~�����s�7�j<ᕸ�&I��S�=}J(T�r��ɮ���]�$�{lm���t�q��({K�$��=�h��q=iG[��o ^�v��nIIzM\�\�o����,m���C��|$�ݥ_�U����WJ�t�2�5�}�SO��ަ��i. �����k��-I�vA��sc)�b6=��� `!�hǿC1>w`�>Y)ˎ�;9=hփ�Wj1�N��-����(D"�J�^l�^�A+:%Oc$&n�j��تl�"%�CDҢ!fƆ��;l2QۈL�Y���Y�R�2�3O*r�1.cp���Q@q0�/`G΍�� �w�����#6�&���-�;r�;�s�&��̬��F���������������<���ܕo)#�'��y	;�/��}�Q�^|Te��m�i�^_���6r�.�:��j{�'mr�k�u������Ȅh��?�[�וY�v���	��.O�z#X��YepG(��՚�O��t3�.�} �c>�=y�&�E�7W�s��h�0暃F�����*��%b�M�R�`.�\�F��������U��d����Q�R��N���	/5�׷42�lw�L�m�qN۷q%*B��)�B/����{���m�_��5�Ë�%�b�8j�4�S�[֕�iM�y>T^�Ǉ�n���*��Yy��=&���G|���~$��0�,[D��ɴ���e�|�XZ��C���E�"cH+���'��X��~_�wF{�q�Y>\�Q�=Xs2��Fh���~+1Y��T'��k�i����r�Ax�;rg���� =	zS��f<2.M�n_�&;c��so�\��l��x��S�AS�.^1��)&��K���6�4�"�	�m�s�+_�8�A��`�B�TP���?˨9��m��@�aM�
��F�u �-2��#K��­PW��MJ��"��+A�6	 ؔ�1j# *�_A��cd�d����7�F�0��S�(��^�u�>��o-���T�ـ�3���]���%-#s5������s����jA��t��-lA������Zъ@��LTW�zg�-��t�0��# h���.�0M������gg
w�;`-�ϊХ�����K.� "2]��p��l�6�۬���������-�F�σ�b� ���Eg/ ��窅I����\��E�J���lٗ%���(`�?���8J�tp�}Շ{�.vӖKv5+j�Hy��D��)�nKL��d_�UZ���P�~�q
:��Oi�f.?儿��[�kR4��t�5���c����uD����Sj���!IUOsad��4Jb�<% �ա��Ӌ8�/i��a�=c�[�DV���;v}AdF߅�×��uys�����(%w �uը޹Mh0�+f�B�4�~��-m-�K����ڵ���8�h���2 c
�A�<9�4)[�s�.�����c8}����8o$�Q�Q��ɕ�`#r4OV����U)%�f������FV���h�#�,�[�&��M�>���̣��;���IM��3�K��ɖ´#g��0�+��GB0�)E�>��u�8&S�'����҂���6�����4�.X���$__�Y��3>4���gͨxhO���3����!����f\Ƿ�Ļ��}W4��O�g���|��� ��� u1`�o]����w8���.Ҵ%;F����Ӽe��v8m7��R�|��w믖S�FP��z�����j[rN鿡��?�Co����6?Ol�.�C1�ׇb�5_��G�0O�н���L��4���.�'(����SE�
>X�j�T��XáEZ�s�,������
��n!J'qFyמ�`%��+ֱ�7D8��^^���2�M>��aR'�?zj@���p�et���΃���7A�0LJ�,�ɛ���y��"q\뼓��f`)"�LQ�p���6��Yk�H�A�'���{x.�3�]�����f!RA#����=�f�[�N�emg������|�s�6�Q�sI4�$kw�7>L���)�)\�Uk�taݶo�p�;p�,�_�P����5C	��c�C*ƒ�f�|��3�'�kCt��j��૾��D��K��)*i�!��CR�%�i���Q�an��I�W߇9zm�̨%�H��{7��������B<2��N>�����#
�C)��YD�g���{,#���w����֞5b�4�������wk{�/B�>���
� �	%�m`�����)��A���ԇţpg�0���}�om�+o���w���w���B��0���?�G��J���O=��6d���d|0���\l�� �E��!����_��^�B��C�l�P3���
Ue��h�)d|C����(O"�㍦���S�Z���6�;'�&D�jT����T�F�Ч9n�hw�m�7�����ƫ��u�૓��
B!-/�@��<P���˴���ׁ���7v��
2��Xab\�G�h��2��=<�,��Y���������im�����b��X��,fM��k�,��t�q�g��?�Pba�WSY��{z�N�l
��9��r���R�vj�qeN8��U��o����0E�X�w�:�b�v��%S��CQS8{}ݧ�������9[�bW9o_�1���S2�&m~��.od�]ׯ��Lg�Iϟ�ܟ��X�`G�YH�l6��]��#���PNY�b�,S4���x�1�v;�l��3�c0��	 �+.����|ֺW;���)�l=�?�DK!��-�"�0#�Pt�}���AA��:��t�E&/���څ�����+R���Q�u�ji��۹����pl�2T/I���PXْ����a?Q_3�D������$��Z���Uv#����!oY��n���c�ܭ�]˙��x��e2�xftR�9�g�]�����Z;��kRP�Ψ/j�����}7)���{�e�idBt�����pM-;����fG�S��p�~֠}O��:$�l65ۥ]=�[Pj��L�����]����ꑊM}�����T�B��q}&��ǟ��R�<����ϧт����}E�
�j�rz�%���]b�~{Gyܳ���#�(v��$X_��#S�q/c�i�"���&�^��KH}IuZ�T �YEE�G�g.0�-����@��U�����J�7�2LA5J�OS*�ԋO���� ������k�A�I�\ASc_�6xH�z_!��3��^8w�~YD���,�h��W��Ե�%�-�<�$�W"��^���:��+3�c_����إp[�}��C���!���Jvh;G��]���"F�T��jO���1I�V�c@L��/�&�������k����6��o�1(M�{;�t1��ٰɀ���yi	�5D��$�c����U�5���o�R!'���	V?���2|���|eS�N�d`����I9<�1k��}?wiu��o'�Ñ��҃��݇������_��ie�z�5{�T��G�l/��VW�jԻt�j��oߞ_Q=��@;!WOª#:�浡��9�س�~�`��M8�`)�0\r�B˄������Q���?x���bR/Ъ�����f��r�ֹ�k"Lf�D�L�ط�g���$~�/p�ς]Ţ�*��mI"*����R5%YWY8eKY4)�y�I���my�aJ��Dn���*�@�Yt^�����\E����[$&;���"��,`�p�e�׍�Z�Q����Ea�/c#>��4\4���9�g@�D{���YY�sQ),+s]
F�+)�1�ϯZׇN
�i�����xʤ�g�F�ņ�P=���EŽ2�vKn,w��e�;>��s�B�ղC������D}SR�
16��)�yJK�Yq�Sڱ�	��B�΄_Hx�A-PԽ�*P��|?N �g�� aE��,k
;ͥF��V���a8kK(����H�0�}�F+��	�!��#����F�B��_WY��7J'K�D��N�(hD�4��uP̄��X�;\����N�����v�;�#��,������T��ab�C8٨�z�}^T�$7���>S�#�W$1.T�.�E~�u  C2��i��MA�8�~�g��Ϻ�l���.��þb~�;�]uG�p?�l3C~�g�+���+�8d�����
��b|���}�/[�G�e�~��`�\]�N�%Tǧ��%:��#c�?Qs�`�gΏ�[}P����E���^�5��Ht�qDx��)������Э���~��:%�hi��c��m��[�1�J4Mut�B���'�:֢u?�7芰j��<.lU���s<}@�o~��S ��	ş��n}i���apr��6l�V��x֜�A_@h������Msy��VEh��%w;��Cp�Mc�r��FBL$�~�А-���K���g���cR����c�
yA$9J�[�8c.�\���3ت�/��o�)�Q���D��`���O�*��T(%��6�-ʁ��V�U�@�#�G�[Ü����6������;��� ����3���J$�O̤�_#���G��p)`b�L��8�T'�L҅m���½���!d�Wf�.sTaݟ�p�43y�S�Y�F�s���,����<���7�Z��]��A���lg��7��?є\C�ҍ�T-]�RZ����w�i8��@ef�ӗ��7/om��΀||���j�Q�a-�?3���FZ�.xr�u�ޙ�?L��x��Q?~lt2��x��0r5��A�B�OR9���l�� 2�w+[�FJ��_�ES�X�~)T+vP�\DD��{V�G`����3SJ��Sy�}�����´ı���D�I�9�c�8"�����')Iz%UC���e��-�u�o�����Z 0G� ,J��V=�yÓ?q�el��rfYe�"�3�QΰP�1v��9�c���{�\�凶��� KD]���ЂR�������=ow�[�ē����lH�^Iq`lsXw�Q I�'kR��>�������)��0ǰ��n@�a��	��Ap���_<�v�a/�5>u ׾Ȩ*��f�<k�ݷ3sH=k~� �l����ܟ��Kb��)E�b!�$�C-b��L�|���c��7�W�K�9�q��#��H�tq7����Y������m;��>���톏��+Cd���]T�b��֪O#t*����v��/y��t�u|����w�=�/:P�:U�cs� �`j�m�a,������!"��]�$��S�RF}O���&hό�����
����f/��Ǹ�@Ц�v�w�s\O]�t��>��F�|�,�7�o���QET���D_s��Ɨ���3��+Wa�G��U h�sId\oӯ�6�C���^m	��İ��k�Z c�1�'��4�%����T�pJЂ����,k�lZ��\�7j�����q�ƴ�ufV���ΰ�E-��@���<��$��0������^Fm�轏v�\2�#�a]�M�����#(�XD�,S�C����Q�[��^m��li�br.����M$�kyR.�K�2z�(c`��i�a6'YfRH{�J�NB�*
��w9��\�Q�y�1��q.@���0tqo�͎�E[��oh�:T�v���%�4�C,z�{Y��B����:�`Uq[E
�9��+1v)�S�%&�����#�ͥ,�Kg���I�)9�p3X���G�q��V(�pm�~0�>IN��� �ݕSo�.��q����J�3��C�B	�c�+	�������02�X]���?]!��)���80�J��o}�
��<�
����/$&J�,�U���+�$���a@�e�!�6�M���鋍4᭘ $Z�֋��#���\I�_� )��������qW��XN\U�o����o��t�)���~�&�%���t�,�A�e�#@xa�t��E�"T�����`|�F'��	�j\]���7]�2器�рy�d�� ��%.�.��-�_��+}G�H��+m�ֻ5?���
�Ga����=�PPe�&L,�|����d2�T��q�]����B��,qI�4�Z6��m��<
d¸n��;��}@�)
��r5F� ��]�=�{"���6���(q��$� ��jqJ�7i=
k���E^���A)Ip�6�!����b�\�`ϐ����~����U�}�@��JGۆM�55�X�S��T�ퟭ: �je�A�	kH�*I�C
A}�c�6�6���6��!�d|����wք"Y_���1@[h�i�W�쵄�
-������"a2^�����u+�`�c��aŠ�ؠ����K�C��v!�r��c;"�@QQ.ʏ���Oyȗ�NaO���1d���њ�@'�/�%T�5�b�l�Ʃ5���6�~��g)��;�~����{�w��4�P� ��xm=�����z��\�oߡ�'r7�	q���y��:^Ԝ
e����_��kҬݲd������ݬ\>�,u��:��Ub�7��#�F��la��:G���zY3n�O�G�<��K2�'�t)!��tio�٠A=�g��;�&WlJw�ޠ5�������������M��3`$�\����?����[�����T��Z��R�_���%�m�-_���L�|��'<Ʒ��rx�U�[F/�j���;E�~m�6��H����%�k�8`�74��-�����y4��}!�nZG*C�)Yo�F�󪪯c:��q $����JQ���_�H[�e2�"ZZ�H��h_E܉1c�p�o�����pC��{k��Yt�Q�:
s�:�Fޠ���1�3�
�9�	ɩi��\�h]�x�-Gg��!��=��2ߠC�2���nG�K�	�;�:s����M����,�	�S��1Qe�)icK[8J�Lf�L'	���)Y_��A)���8�Pp|&?A۝'��`�,,
���F��T�#�<mKcn����Q�C�c����+�o	6M��)#ֱ�������z�Z�PD`7(�fԁ�j�(Cϵo�Tu�yv��������OxLi���S[�fq!#����ǠB���k��9�ix'�"1��#���X?p�_3M�v��(W�Q�����l �金`M܊��
@�g�������e��\	Ù���v&�]��p��l�od�"j׹ZN���S��xL�E��b�����/�:�� �����N\�b� �f��	(%���K?��5���ΪZ�}˸Ǜ�}H���5a^HotDu%i���r�%X�K!��v��~3�h:��yi����uֿ:�ߡLK4�3����}�(���FAu:{�C��j�_4�Wt�U�s�u���f�Ӻ �S�d�+��h�i*a���P8V)[q��AZZ�;Q�\�Ty��h�W��"/wv����!�M^�1��N�B4~�-c��Kb�D�P��6��^@�Zq7c��
A&�9�C[�-.'ݥ�)�X.SR��d&o�O-Q�P�vC`�q�O̵����%�Һǈώ��=V���ߖ#���[�2ǽ�>'����Y7^;Z+
;B�C�;3_�1-�E����	;2��GG���){ ���I8�Tc'*���ʛ��dO�7����?.��-����G+3��Ε��n,��`ݺ<���W�����"u��: q��J����g@���TF𞊔ׅ��c���l])Ǔ��Gw�p�ʤ��[�.�����r��r�mm�����|o���%r��|b���s��.N�P�r�^��73?��#�3��l_�l�U��6����5R�ѭ=NAO���> R�/+��򙓫݃��7Y�E�+�X���T�)��cҡ�q��� 񻏼��nW�J]h�y�|�¤�}^w����D!M�f�s1������%'t2Zz��u��ej��P,L�w�0BT�,��U���y�J�qR ��Z�!f��-"> �Q�{��f���{�~�q7{�7���廂�]�3$�B[$R�̄��=ꧪ[�P��������T��4s؛Q��I*��k-��>�B��&��)͋���),�a]��fpb8�_wM1����59��ԭ*<`=fފ�r��3N�>k�J͠O�L���K��)`�e!
�WCN����:�م柒�@W�ؘ9��-̞T�H�W7��EX�Ք��4��ܤ>Ӟ7���m�C��2�A���]�a�1b�#/������1��/�5�����w! �/�}�U�ݤ��o Кf��m�\��I·�ڷ��Tř�j�k�S�� }���!���p���H��t���M~�յ��{y͂�s�W�O��g�����|&���~��8I�E�2�|�_�(������Dԝ9�A���UVU���h���d��z�j���^'y��l��ȳ_��5+Z��,^�'W�%����;�Tv�r�]M����P�Y��l�7ŷx�S�d���u��8���ˀ�-T�2@��c<ѫ��׉�4X��&��í7vo2+vGaXD��z�b4��slW,����Q���j��\Lm|MĨ�b-�_��2PM��;kT�8����9��d{]߃Ə�a04#Y��{�;�N}��
D�+9���׬~`�쭪q8z.���oB��)�E-���yY:�]va%I�}C��{�;��Y����L컑�[ Ү9��1�ˤS���&㸋�d����crig~�IԎܕ]>Xn3G ����+��ؿ��f�&N8)��Yz�%OS�7n��خ�l�^�"53B�"i�		��+�s%�P����F��!��"�?S!�:.���0٢��}#��7I�����ꢀ&e#��И��^2+Ȉ���MC�`��������Ω�(��MW������Ws�_�/� [���8�}c*L�m���U����۵�o�������������O���;ehP.x\f�tUq�����3�*�P���!�D�<j��ș���7����c�_ћf�d�B���Ÿ�i��-= ���oG6^ٚ�-����x�ݣ"�!���=Qy<P`��L�[��7�=��'���z�Lv���H�B8��q5D��T���[z<�՚�I��G�f���};D�ew�r�l*�.o]X�9{���Qj�B`�(lq�$���qeKQi�����^X���[MIk���m"����}Z�����8H-\4�v�IU����� �J��h��5@��S�iۋ����:�\ �M��� fk=I
��A��c�.�6�a��z!���TMw��*Yz���s�hgRW�x��-�#�ڑ�"֥^��W0]4+ˮIc���;�o؛�=�3�Cu��!�x@@�;��@�e-�*:��J�ݗC=O[?Z1��L�k@��/EՍВ�F4�!�6�=0�6[a�'�q�W4;#���Dy�������%��"�k�	�YzH7?�1)���rW���*o:'-�
	��֜��{����3e�*9�Z՘p,-�gçS��'�f۸��y�CuUH;��[y�y���p� �(Μ���p�5����z�PY�JxhG9-�.a᠚ t����O���=J��6SHW�e̪�'.��=�/��5���F�Mnͤ`�\(+{���ũ�c�G;���O*��WIRemk��"�@)��˹���L\4��㣷"L|8�X�/&G�����`��m?΋ƚ�<Mf%���8[��4�I������y��&�X|nS��*�_jYjd��N���Ҡ���fm$L�Ϗ8S���e�e|���Z���HEWmc�Ö������YV������{&�Y�]�Qi�s�8FZx_�z1շ�e!<�ħ�iL�����x�ֹgV��żE�=�V���� 2_*�nb�.w��;�HJs ���������d��SȬ1l�)�x�K67q�&m��&		���M�_�WAD��Գl{PK&�?|�ɝ�����#�rK
�F�;����G��K�^<�!�A�>�R�36�+rk	Q_U�;#��)���4�x+��U����7�H������](z	��u�G`������|��
$T�������A��#$	��b����
K$���=?0ٞ�r�3@<ΚO��f��	1�W��������k
 �iD�߱�Mw��"$gx"�l�8� �L����t����X]�lp�x�l�J��A��2)��.�XӾz禀۫b�n��M�/����MU��x\S`d�ۍ��R�%pA�ɔ?���֡o���Z}F����)�G�5�9�Hj�qD�򘳟U��/���ƴ�Q��~n,�:[݂i���Pn�����g|S4C���}��c?��p��u5-��JjH�u�r�*U�1ks�[��F�U�Y ��h�Ax�i�ei4{�af;Ƀ�SjVdډJ�AU�*ߖ��wy��;����(w�(�y�MY�l�<�}B�c~'�4-��K=4�����r��Y�A��@sc;`�AAV9�R[�"'.b}���L�)�^�oA��Q)���:�`�!�OaE��-{%�8����D�OV�:6�_#���[9�x����H�̴�\;��V���3:�Fh��}h�7]�<ÍGs��)��
�B�78�"'e�G�����+H��N���)�.��Bݕdx��3�Y��CB�i�_���N��	�r��u���{p�uU�Nt���`g�����v̔R�$������]�[e��-KwI�*�_�Rv���Pg�M���xm����;|�M���ɗ��5�6����r�g���E?\���5�ه��lj������8-�5�Y�8��Oj������JV�m(ث��f�rr}E�l�X�(T���ҡ�ć"��٭�j�⎩{J�yț�q�;�8(��,D�E���=��`�"�����'�[Kz�ދ�'��e傾�+��@Jd>g0=	$, T����y�!qͺo�5��f���"��~QĐA��T���K≙h���'�>�,	��V��]�~���RE�.=e�U[���������jw'�[s�X�Q6I�>�k�R>�����k)�l��f�%�7a.�V���p=��_����@54�c�t�R*���f��}� "3)��k�'�;S���ñ�UZ�Kح�){�!��C�YG3�Ҳ����,��mOWF�w9�����Hp�,7@����v�⎯S���V>���|����JC�ߥ��<�X����9�#�s�Ȝ��l�i�(�pJ����o��9Lw|"]/��;p�.�Y�� �Rְ�m1w�����:C��r�S�D�����F�5�{/}�������� ��C��OK�\����ZƶB������[dOgy"����n|���6U�s�E�w��w_)�	�<k���ڝ������4�U6xzh臞d�f�%� �y���T�ˣ��� �Z�C'�'��'��ߛ�+���T�%'�8��H���\7 �i��{��x�u\����x?˻�h-���@���<ag��O\O�ޑāT'����/vZz�2��aS
��X �e*����,IOܨ�[]�����S:2mw޳Y�b腩�f�M1�k/�ң�m������������baKRGY\�k{�LdN���
�C9�������2qS ��3U����o}Q1��,�E��%��:�v.U�%�wC�'�{�}@�x���{[���=[���9���1l��S�[&����Õ�����g9��I ���k�XI�G;��=������4ux�$\NS��������XS嚤�I���g��}�3���=	�	���+����g@�(|D�
��}�c?�!��:���h0�`q��}�+\�2��KO�A�&���K�k�_�o+��"Y~�[���t�G���/gᣁ��a����Y�>�R��_Du���/��2�'����b�UGh����ojѫ���S����*m�)l�e��xWFtc4���H�N������0v�Yj��3��G�7���D8Ѷs�dx��ࡅ�ϤB�-�B����=G��v����ׅ�̜����VP�=�!P[�L���@H��
ڑ��U�'���NB�}qA��/��K��)%< g��$j�����qS}6�-�r��Ү6�']��	{�\γ�Q��.�(g�$i��T�q���i39k�ZL^����IfA������P�����%�����hY��2gU�͇��7�J�?7��Z5���S��&��<�լ6 {P����k��7I%�As�c�F26)"P�l�K!�ࡿ��gwL֖Y�K��'�)hB�YWV�x��v-����5J�"י�^������+�hc����ؖ<�Ԏ��C0M�!Ҟ����;���Ǚ������E�.��K�O�1�����a@��/L�*�k��@֧|�����65Wv�F&��x;^�˝�
İ�o�-�_��5���z�
$#Q��l~%�&o���\?o���'��	�U^�o����J=�e$�B�U0���.�"����,�ۓl��X�u���l�����+%U�Cv��b�,�uP9�h8z��<�Ei�G�=���I,�-/t���*��O��=�8�1�W"���T������Ex���
�әM	�M`�\���˵ʎ�����e��k����zR �ρ�t����ףg��#L�Y�ݩq�]��e��u:/����<0�{�.m�)���w�%*�58V��4:1��Ga���5y*J�3;zn���*ycYe����������{�$�Ǡ����s[�~�Ge�s��lZЫޖ�H�E�p�c�6���f�R������X?{�Y�H�Q���s�V�FT3}��1�W���އ��i*"^�^p�x[��g��U�W��=�5�V��2��n}ZY�i;ϼ)s[��Ճg���`�俠pS��i1��+)��KV�"!hڂhc	�����a�_y�A_�N�.��P&�?��̝8`�����͊
l�F
�I��f�6�K�n"�����9������+-�	l�%��#�����ٲ���PyO%7{�	�d��(�D���Zu!5B��2ÏL=��������I�[�=V#_:X��1٘�zԔe�Z���Xm��r0�a��Ջ���)¹h�W5�����0��U� �5U���Mȉ� $�g�O�'SZ�;ۛ��K��Og��6]F��p�ElD(1ۘ9;�M,��{�ә����8�bMs���,/lIS����-�J\�}qضZ��X��%�)�,�?bZY���Y��Ć}�iD��M[ӂX�5�dHe��D+�(�Z�)�Je�AhX�,�~���:�"�i�����(���s��d4����K5�������u0����j�[��`�U	{ws͇� �;��0 �Q#���$��iO�a��؃�wlV�y����AP���cݗ�;�y�a���F���w�K��LMT�#B}�%~BF�-Y!K�̓�ʽ�P���T���0�c�:�A\Ek9�J[jGQ.�=O�_.$�շ@yo���QD���`��^OB,"�%`�%��W�>:����V�n��#kX9[t����Y��ؙ����;�q�9p�3#���E� ����R���^�G.��)��I��;R8�֐'����>�0��}���򈻐.�O��Qn���3*Q@�*"Ĩdp�����������؎Ȣ�ް-�����Ag���h��&����j"��f��(]_���u�w�����$����x��(�>�Lm��H���5|%�����ɲ,)����^&��7�r�S����4?]�X��~�٢�{l���诼��s[�5�u٭3�BOc2���g�e�O���(��_�㭫�E$͢X�z�T<��Í ߽ۡęxӖ�E���J���y��M�ޒ��)�'��D�9���a�鯄�X���i'*�zVS��B�Ge`)�
ջ{����>08��,[�⛇� y�qH�Ó�f
5�"t��Q�0��B���E�l��J�-���l�gy���Q�]�����'R ���'��=�h�[�0�Q���=�������s��DQQ�mI �bk��;>8/��\9K)�m�����c#aI�	�\�p��_�Ob�2�55/y/��J�*��vf�Chr�3kQk/%���vW��Zܰ�}K��)��D! �C���nF#�M7��)ϟH>WR:9�=�̔�HK��7{�*�{����� ll>	p���X�Q�Cݟ�w+�S����0{#�V�������U+�k�F�����:w�D$/k9��H��l �*�nm̱���D�����-�UOŏ��!|�Z�} F��U�&����Ʀ�7J	���l����+ׂGͳ��~On
�ݱ��7�|�������E%�"�r��_�������
�)�/�G������3�U�^�h�A�dm�2���k��p��˺�~�?*!ZP�=�"H�'��VSA��i�Tl�g��T�T��B!���7{6{�����u�vv�_�����-��@�ǹ<���
"�����GU�y�wv��J2a{�aN�J���2�ص���r,ĺ��f6ٗ���7mr�Qz)�b�aw�,�ZM��k
����^�K�m�< ���<=�af��Y��?{|}�N�5�
z;9���b�n�bq~qnI�$�d����o��E�_k�E�0L��K:���vIi�%?��C���{
�i���v8��qj�[v�9ۛx1�p�S�9&Ys����=կ�g�I;�2܋�XX$�bGvz���tZ�i㿏G�oB�Nn����)�x�S /�䍌�bS����T3�F�X�(	�M|+�����K��������?�Sk!qO���0�>]<�}Y��-�Η��"�` L&�/���+�:P]+>�A����V%��G��e�ܰl�&=��[�<U����M'�_���0������s"��A�	YU�i���oťG�Zg��u5��8���yd1�e�	�xRF	t�3)�S�4�i�T�F�,��e8��)j-�V��7n�ٹT�Ѡed����|e���p-s���}��G��s�\���n�G�ء�ۑ6�=���PVN�L=<����֙�:�v'����@bBn��q�l�E��ǋ���<{и�Jʧ���ט}1�*rf�?�Q�(]N�%{��i��X�x�(b�$Ĥ�F�q���i����5B�^Αt���IaΠ�#FD�Ed���m����ܣ�vݬ�U�%��Q�4Jx�����56�FS�c��0)�p�� vs��R�ky��I@s�A�4�cp~�6dU��%�!��~�
T�w/gY����:sh��W���U|-�` ϐ"�"�}?^�R&&��+��cKT&�q�jؑ������C뻃!��6�[;�Q�G�`�<�@���y�O��1�L�B8�@�c"/��S� Z}Zԧ�U����6Ps���FtU�;�]��z�W��T$���e�L���s�"�����c����Ѽ�o�O{'��	�G���H,[����"e��P��&�p���]����U�n����nu�ň��;�/�����^>R��c��P�ھU� z*��@z�G�m��|�{���et�����ߊ$�=�ay�,��W}�V���!Zu�%��q7D�LM�/`��\���p�#V)�=t�ë�֖��R�������k��^DQ��{�LR8ȸ�/���Iof��n/ܟ��I�g��PSm5l��|�yò��%�iZ8Q�|4�8	�T��Iy�׳�x�nɂ�*�Y`�x���H|V���$�j�s�����V�ۿe���CC"Z��?�i-EM��c��;� U���S�K�T�={��Y�SKQ&�sy�nF�,���1��h!�:ňiE��)Sx6��g̗���<�=�4D߱~D2�]�n�;�m�8;�P�s��=�^o��*0��,S>��1�i)��6K씏];W��5	�ԧ:��_4�-AzI^ԩ��Pڃ?�"��,�� r�(�/
'8F%`@��m1���K�<�W-J�4�d��*�+��	�Y���#g��2GѲ�P��Ko a�76���ܩ��|�(�/ 3u�B���ޏ�7����n���N���H#������Ș�����
�|O�s��ٔ������M�G���(W�J�@�M��i��a�( �!6�U`�M�U��E2g.�����_�V�R����*��'Z]�mp�2�l���SQ�h'�$n�t�M����b藬���$/� B�Qs��H��\I�*ؑGyǓB�%�@���[?�<K�L݇���z}<�e��ӽ�52�H`��D�����e5��;��_|~�H�:��}i���k�����|49/�|9i��qu��X�u+ǒTXej�k妨�U��s� 6�[�4�&@ � u>Q��^ij}�a\�4���>V�8�BwIAKh]�L��� Ry��1���o��w'�cկ�]MO&W��B8#>~]��-�aK�G*�����K��O��k?Kc�5�Aw�(9�u[E��.�����,�����ko��Q_C&�0��`j�1O}S���?%{dpǙ�����V6�,�#F��[��8�T���
��j��;����m��J3�h!ޏ#»��������G� )̚��8��8mǯ'۽���$����H�*�Cm_.�8D݋]����E3eh7�� ��_B7�q�m��񨡘�k0���F��&���'�� �gQ�#L�A|�H�x�$�@�]������'w�F���/�Mx��g�6�#PSm> 7���|�Re�V������+U��]�
�{4rU������?����d�4ٽKl`��芯�׮�r5#�Q�.I�O��o{�ހ��c���n����~E�M�X��T�p�HU�����쫻 7��$�J.˺y�9�'�Ϯ(�B=�D��!���V�$T���z�'��z�d�]�e����ᨁ���H��03�7,�\)�B�9y/0qÏ���3�fE�J"&�Q���� ���L�����	���i]�t��S��R���B�N=[�[\й��5.�ؒn�����sD�/Ql��I�� k�4�>s����")��\�xZ��adF���"p�\_(ٽ�т5*e�*�}*m�	f/51��<3�ckj���q�T����g�KNQ)�& !{V_C�������kʫ͟��W�>�9��H&��7���� �\��	�\'��>$�X�rOj�CP�t����N��BH#`Y��0"�b��|�q���z��z�����w2�+/&���W)�OU) a"KLw�mg������ ���!���
2[��K>X�}����$��1��yj8�Re��Ri��f?=�,5���������O������R��|��������%AE���m�_�y�����%����ż��&��3S�UleBh�ddȺ�ӛ���[��J+��Y@�zT�Z�̉�1'h<��#[�19T�Z4��ڶ��Aw!��\G7֥���i�2��uRl�:���1C�-%U�@�<|V������J��T=v���2�-�aI���kշ�&��Ĥ�,?F%�A1ŗ=bP��U�mm`���b^]ɞG,�M�Vk�)��7���ri��ln�����a��YR@{WμN.�+
�9}v]׽���q����쿀���o�.���{E�b/��m�:@2vd�%�R�C�U{Eb�ݮV��q5m��[1�P9���1bs)Sb��&� ��56����th�g��lIV����gX��[G���s������9\*��N����yS�[S[���?�]��3 �3szs�E	z15+uU��˺^G7��;�3g6?I�=!+<l�v��0j<�w��}��)�(ŝ���ߧ&���A�����+yu��XМ�Q������V��Q���>���w$(���#�H��_����.�(|��1�ݒ��D��U}����To ����+��쟭����^�me9��xMf�tS���D��Lf��6j۲�*��Wj�{1���E7�\��O�����dn���We9�K-�7�xCoGG^њ0��'V��#ߣ�LM��<1="��PQ��L���hx�1���"���{
B	�Dq�������FQ���%�<��,��K������zS},)�v�r!Rp�l�q]��{��ճ��,�(]��$ƴ�ʒ2q��i)���^	�:Rh�I\{��~�՟ <�g��jŐe�i޳��G�jU� ���J3�#����5��rSqN�@xJ�, q�M����k4�UI[�Ai}QcK��6��*��v!��7�e!�w§�Y�K��Ψh���W�\յ�
-�9���:"M�R^Ι���+\XUc��:�،dd�D�C�J�!Kc�;�ga=bc�����;u��TȽO�,�1�iPĽ�2@�g/�bQ��fx�.�2�z�n��6k��嘥�O�;��L��c��Y���� h����� ���D�∶�\�~ѷ�<oKb'^b�	�Yf�e�6���]�eZ�}�KFp���Ҙ4�����M�I��*��u& N��-焊��*�y&	�XOh�+�뾐�=z�i�;�=GJ�|�7�N��t;�������=Jҵ'�UW�w���{��<���(��L�-�K%M?hH`y*\9�p�+�m�>����@Æ�F}ZR6I���x�Q=(�Aj�,L��ȓ�ݷӒu䘱�/7�z�,�����m��ދWPB���%`�8L��4�_=��f΁�$y �����n{�*��|Y[��_4ǯ�3e$��ڠN�,�����Ee�US��7ZF��.��E��qcj|6�[c@��z���j���{W�2Y�~Q���sT�oF�EC0"�1�p��v;���i`. �T�x�2g�iō�*=�S��}�2�'+n�<���S;�Ys��չt�����u��S�J�1�U[)g K���u:ڸK�	��n����_�IA� ��$<�P��m?-h�n�砃��iq
�sF@"��s���@KO�b�/,��DՄ+��	��4:#Bq��m��I��F����j7�j �t���K(�:�[�1uWp������K�;�����?5��҈�#��v�3CИ����'[U��)���0����Kd���z��5�W�Q����<��.� �-���MH�x����g�2����I�qCr�w���� �b�q]|G!p�?l�`������V*�����O@�1Sb��ב�u�/"�P�6��c��\���lT����%A���
R�??}�+���6}���@������5�)�H[l�D�i��q��%+�7/ʫ���~�:,oiz�5a{�&]����4�m(�WG-�;��AI�u&�o���jyZ���uU�ms��+��c�&�� ��L��݋���i�.a�X܃}�V��=AF�ߧ�*�H%�yz����J��wbpo�J(�MJ��M�QB�Z~x4�-O̓K���<����]�J���n�clP�A�	�9��[ �5.���I��or&�Qz��䫸�`E�TO�"ح[%f%v*e��$�u��V5~��MC#!�6[��F�����Λ���8X;FZD�NY/}�3������V�B��ꆏM��G���)�?���8H�~'�>�tإ��@���}��>�.�A1��>�{v�3���`?ШZ4����J(E��Õ��槫~P��&i�������xg�D�3!\[�����S���{^5]��j��e wZΆʐ�5��n����^��m�_݀�c^|�"��G��v������8?�<��r�Ȩ���?��p��l�#<�e·���5����)24O#4�*��ޛ�6�ޓ�I�J�#~�EZ��X��xT�6��t����n&����Z�TJ���y����{��iE�]��D�rV����_��%��u='��_z̜'�xYeV�B��g��%�V0.��,p��;WyJg�q>��Ɲ~f�_'"�r
Q��=������K��n1#U4����ݹ^�'��]�����+Rvcy�]��=֩ [7�������s���l/8+s��~Q���Iъk��^>����4�)���wra�a)��RbAp��d_c��h��5%qׅA*({@fJG^u3��$k���������f�K	ӿ)��C!�2�Ct=����҃���M(����WwKl9fo̊21H�N7���9���e�d���{�>?����E��C��]��T��I�-���#|8����gAW��!��|�����Lw��r/�t
��Ҥ�]� <:���m�i���ԇK��ڣ��<�#Ņ�����}yvt}V�|�%������4.N�m������A���g^1�}NT��&�O$��S/"�m��||��~!��$ZE[J��h�_:�/�m���@ɟ�%�}�r���n��U�*h�Qd#�j�V����W�ŪM�4�|����Z��҉�
'à���y�"Tb%����(�ʖ,�I���715��?��M��úd�g~�l��-���@�] <r6��O�/i����A�/��v\�2� FaD��iPطN���L-,��L!�x�/�$��mhQ�0*%by��b��M}�"k���rA��}����H���jma�l�Y�Yl{2?qNi.n
�+9x�s�X}�شbq��2yg�w�Mo.��͕H�E��n�6��:��sv��%5*�Cs�{���I@3�lRp�'�q[�0�9��1ݕS=��&ϭ�ЊF�����O$gj��Iq�v܁S#X��G����i��޿EL.���N��_��z<.�US��@����X/�Ď=�3.����J	�4�+P��<r���ܤ���%���_?�!F'����0EZ���u}�ʹ�#و�\���ݧ&ѻ�ռ>����H+�Y���;��L�\��O�xX[�P�όk]�ֲ��*���C[�_Uo
����"�b�ia������pU����lo{��ІJ������˻jS��e�B�xH��tt�a���x����<�Sۍ/M�0*�jc�ę�<7$�F�OZ�[d��t�2��U4z-�jJ�s�G���pB�B���db��<�c�=�o�PLpbL󜧻#D��4t�lT������MFB�'q�$��n�����S<q۵��lh�3[B>F}'`H��r�3e���]D,B{i`�=�w�Z�(X�
$zY���^qћ�i�o��^^D���IWHT���f��3���V!=!�@ @%���PU�5���J�gІԈ�5,�JSL�)�{��� l��jXk�JIv�*A���c&NW6��=��!�
Ϳ��w}@4Y��5영�h��W�1����-�2�F3N"��^)i��+7&$c�F�ŧ��؇(Tԟ\�Ca��!#�i,O�;i�!x�2ʖ��6���6uOGfV1�ڜ�8A@n��/�#�<�s�䧍h��)�^6�&���*��;����簫~��>w3�g�����{C��^��>��$�Ѳ�%o�i'=�	������&��e����F��մ�S�$���u�$|�eZ�u�R��׳n��Q<�\��є.���Z��am�ˊ�z`��6�|G�.���\����t��5���� Ǡ=�RC�"�W3b���y�W���ʤ�'����7�M�ۙ``�\�������Y�p�3-��aÖ�tR�'��*��.G��]g�)��LHR:�n�{����t��K/��6�����n4m+Q��2"�(¹%��k8G�4K���x���&t�y�R��Q�n?�*J�YV�F������׽�N{�$��)��$ K�O�8e�3��]�Z&.�I	�EC;cEO�����#p1�}4
R�{�
Y���Qcs/pF˂�1�����.���b�i{d����x�egB �(��=�|�g��2Kqn�]�c �;`بs>��T�?��
��ES���1�a)��5K�rn���S�B	�����^�_��iA�ԟ�P�h?h�N�	&��@1���
�-	F[&�����U�K�_���2�*�g���Q+^�j	��G�|#�������x�A�|ϝ7���,M�w��(�e���u����
�]>�����ͺ;��^�#����~ĔvrKʞ᩷يs���MΆ ӊ}4*���UWF��Y��1<;�W�w eYh�ˎXM�����g��G�XY�����������a}]A�p�l�lU-����o��������*���lbbA���m�/}�����~ݰ\?���G���	� %ܿ��?sa���1Ժ}2c��u��3r5hd�HV��D<h��x+��5$��B嫽D~Z��:ǳXiu5T��d���0�Ө�4/�p�2u��O$���Y�u!�h
 j4i�޲�Uz�s^�ѫ�WB�� ʾ�+�*�U)gi���aRMЃX�SVP�x$7AA� ��Jy06�'Y�%�pw�zo��y�ME2���B�b{~���-�V�K���w���!�x�ERb�!��c'� A���9�jI[�u�.N>��0+S���Q��o-�eQ���&�` !�O�M����d%q6�O�q0�VP�z"��#���[%ɽ��b��L�� 	W;6¡M�3<3�T<T���_��f"����G__Q)���.�8#	�'Q6����������'��0I.kf݁��VR�3�����}Z�UF�'4_��*�ީ�a?�Y���a�m��Z�Ժ�g�/�;bwZ#�>�c.�����]0���uw�u��K5t���Fӹω� �mt�;��֌|6������LA�!&���öwar��n��-*?n����f��ߢlV���@�G�$�+5Y*�$;�OtK����޶B��Y�c�$�a�^�E��+X��vTM�@þ�6�0 ���Z��($��L~Jd?y�W���$�r�x>Dv��[)���]�����p�';A�z�qζ�œeр�F��,sN~��0)<,l嶛��xye�q����'~f�$"E�Q��t�S���v6���ڐ�~Q������x�]���	�R1٠�x"�=Qz�[p�����0�%���s��1Q���I�� kt*�>�r�-�)�0�����Цca�,R���lp��_�Â��d5 �;���(*�fe��&3���k๦ͧ����������K�t7)縯!q/�COɀ�n��E�ߟY�JW2x�97*��zH���7,�e�L���VP�����3D>Z���h� �mC��Z�H/�DK����#־�4E)�XE�2���\+7����pw�k�/�B��AD�E�� r�½�m�!������8�^VhWEj� ���� ��s}��c�޷�7ª���و�s�H�-�;`Ƣ�<��ȱ��O����|��9�YZa�_�qE�%1�c>�_���(��[�Ɲ�N��M�~��U��jh�/�d~M�����s�@J9�>ܞ�9Z!JQ��_'%�߇"��=yT�rФ.���W8A�ߜ�7��o��~A�h�huH�]��K�˧#�-[D`@��=<��;3׉JFG�@ij�
=1vF�-22��a?b��U;�	h���g,5����헳n����zmcb�Z�bԴ��}r'M���k��ݣ�����p�$�߃m1�a�
iYH��{��N��d
KR�9s���s�$���q����%[�R��oin{�0�rE�&
瑰�:�˳v�e$%�!�CN�{�ƞ��I��g��삟�[���9,Y�1XؓS��&
{o�k�U����*W�g%��I�����X�#�G'����������~@�[%N����oS�	m�S�gǵ�.�S����U3� ���7	pXk++P�w`'���
���A��W	?��n!a2��l�Y0 ���}*�W����\��K&���7���˪F+�]V��Ǜ�G��X.3$�-�-��&F�z��"��ţi�>%�_�xqa���=���䰺�����U�.���^�o��Fm� ;���˖TXA�eo�xCvt��-�4���p������hğ�kZmj����3�7Q>�
�B�"�dd����ϐo�-D5�nG�������]&���ѣi��B�5=X}dPG1�LN}��/��O׊�� ��#���B?��q��Vz�Ǽd��a<��j�����nh��!q}"��,G@r�5���]��B{DL�x.I��(Sۊ$�hݓ@�oq��i}�Ʀ�^����IR5h�4���vKD�fG|/	�B&T���}�U����bU�J�
��5���S'�5��h)�A+� g���cL�k��I�A_n�c�6�U�ش!�X>��w8�0Y���U�h��WBy�&M�-�Kϡk�"��^D$����+�c���B��؂`���XC�U!>w����;Dy�����1$��1�̗
��O��1l1ĳ�3@Iϩ/8�ȍדjnh���!^��g�6���厄1��;J\��K�㰦�*��[z�ת��u�������C�X�����ѭܪo�'�7�	��[�����6�e�p��A�7�� nE)���6��k��E�u\���Y҄@����ѯV/�N�T���^��z��z�1m�G �O�����'�:tg�,?�;�	=Q{̵?�W��ת@���r�r��������C�Muo#`gf\�j*ˡ�\�t����9��<r����Rl&Ӂ��@F׏�H�D��Lé]�I
�I�/L��)�/���z�&��-�m�����c��%��X8B�>4��3쬁A�y@����Snz˦*�]wYQ#H�9֯y�בiH$�&���_cC��z9e�1�T�Z����d�$E���c B|���>�����F�e::{͏fY5�Q�1Cs
#F@�Yf�1�x��,B��k�,i��B�Jox�Ig}dN�ß�=��r���J2{n��ބn;;��sG���,��H��+��SoT�1�+)���K}FJ���}	���K�_e��A�.��YP�Wr?�R���Rv� {�9�T
X��Fv�ޚ^J�K��í(���%"���^+�	��8~5�#��k�㸲�� �<r�07ġ���0(e�=���u�+{�����~��^8X;�5b��T�#K?�i�'��j�����ˠ<��eZ�x��z$������x���FW���q���LՁ�҇� @���V�M~����k�g?���F���+�m��û����3}]�Z�p�l��ۄX4��I����dধ��b�������/�����ə7#\�3_�"�<�D��%w��� �?Σ��}&��L}�Kϛ�lB�ne�5��HQ�}D��)�F�I��e�-v쫘��~��f:by:ip�n(ο��͡���4�JŰ�e��-�w��u3~eB�j�[����U��as9�'�lW\�� ��f��7��i���a�a�3G�V�64+�A<���]	����TyK`�d7� wؤcՀ�aM@���	�Bi2�~���-E7K�ՠ����弁+�@�p�|-�c��jA�MQ9u`�[��.�~��rzխ��"�o��pQ���q`�p�O.�ޭ�j;%l�Ǫ��덆VknO�D"#׃�[`X��%$��{�{��;�1z�J%
�3��!�S6����ڏ�G�_)Uּ�v8�Y-'���������Yna�tBd.0����B?�1N�3n���<�Px����S�^��������x4~ޜM�U$��Ϸ�gb]ATc��y����	o���X�]�"g��Յw=�������d��Ӕ̭Ը�mR��iw|��[���A����F��=���ur&�����?ɮD�����*l��W�HH�_T65􋊭dOϓ\�����>��������UE���X���T����y���K�ޙd�����\J�M�y�d8�p��������D�ۣ�6}��,�%s��k1C'�
#zBfY��Q}eL��rE(�gMk�N0$r�,����s�y�5�q4?��|эf�	"�k�Q��Gﮱϧ1A � ����Y���Sz��]p�]��;�d90R�n��o�=�j�[�o��=�c��ZVи����su�HQ���I(ckO�A>$�Q�ȯy)����-���R�a�O%�HO�p�[%_�Ե���5�w�;��*�Țf���T�/3p��k��BE������pK6s)�c!�KC*uZ#�ҹ�6���ԹW��.9R�̀�wH�4k7gԶ����X
>u�B���z��^Cl���g�?�<�SN�#�!;O�(��B�Ie�s㪲	I��HOwC�/W0>��}��� �� ��m8�j�� ���ϧr՘�{����3��}�C��{������٣vR�ä�������܂�OU��N�O����,-�qL|���4���"E�!��^��_����	�vK6���(���pU=9h�i?d��#�̪�� �@��	����+�+�~Z�H��0'y���BR��XFeTX���=�@���tѕ�l:7���9ƃ��u���P�����-���@�s7<(��x��eC���	_���v���2�Va:���{���8���,��}���)��$K�Zn9m^���Mb�؞�E�Ms�kv�H�裞���l[��(�a��UY�<I{��Nߦ
��9nkU�΄��NxWq�-��-W�o�E��˥rE��쁲:q��v���%+9�C)
�{����s'�b���ݛ?[b 9Gإ1�:�S�@|&Eh��������~�g�LI�p[�w��X��gGb�<�D�Y~uʿ�В[��N�G���K��t9Sk��Pxi�N�m�D3�)��		��+�u��n�/hh��vZ�D 3?zb�!|]��40���(�Q}�.�a��0��L;�&�ղ�P��+*�ō)s�BᲜ�,�˰�H�S�
�!�%�(R��`���9�_��=�X�h�_ OnO*��EYUN�ͽ�o17��F&��;��b��q^mP�Se
�=x>��t*q�?�M��2��2�+�Cy"���Fj�"��~\7��u���o�=��d�E+��$�����-����i%,GX~*�HRO�x�0�Z�-�Dj�}�=�!PB,L�}���;:�jZ�b��n�J�,{B�8�q�\@����w�ĩ*�<gL�kǧ��x%�}.���rrRW���d�]:�{X����^��(Ng$0�A��8dqui��O��]�^�F#� IMB��7��1�����A}����+��I�U�����,[Jd͕�
�F5"G�S�q������B b?s��N�ke/I�ǰA�cܝ 6Pb��s�!�Ƌ�vI�w�ёY�E�H�h�}W}7G��ҷ-�������"~L�^_�$��+�!rc7���݋��}��UC�C׶�!Y=�"B;2��~�����,�J�es$O�9�1!�.ʦ@$3w/s�B�rZ if�C����lt6�#��	����;�F5���W��(%��_�Qg�����q�j���'�->�Ѩ�o\M�'�R�	.Pߜ�^��\aq�qe+x;�<���j�����!�k�	����{��P�u������<M�����ʞ���Ѭ뼶��A��z��6�,��G[oy�h���B�t����q�/�v�=��m��`W����w�m�m��ݺ�8p�M#�`�^\Jq'�\�����ء)f*������RE�����bq%�J��_�FL>!��$l����z��c���/HQ��5�n�6m!�܋�%�Þ<�%1|�8=b4����^ҁ\�y�Mߛz�Bn�#m*��YLv�p�=�4�5���e$�~�߁Z��Ə�Ee�O����Zw��)GE9bc�TǛN��Y���/��B9{��FY1��Q ws���F{QC��1�,χum�&�Vi�0���O{x�k�g��N�^��=�p��8�2�DIn iY	n;�s�<Պxp�̒T��S*	�1گ)yu�KX�I�ډ�0	��'����_ ��A�e�ԕ+�Pm��?��	�?����`����
��F�(���C9_hK ����K�� �Z�U��+�'	�����e#�P��t��a�7�i�$7"��#���m��(@2�Zu(�5��7'�߇�l�X&;iͰ�u�cj�#�|��w�|vF�,i��~��3�ـ	|�U�v���(���2��ZsW�ch,=��g��Md� ��A="M�����g�v��R_���@���?Ö���&q]M�p�&�l&��?���ԣ$�x���%ܦ��5bTjꑧ�/3>�=><ɴ�=\5����:����%�h����?)��8���g~}(Tp�фөx�5�98HLvD�b���ˑѵΉ��߫s�R~�}:�^ikG�r෿WH�	�04%�%��0ڟ�V��9u���%j��u��)Up�Js�-�G� �T� ��M��˼�i�"aH����V�u��Q�A7�߸B0�y�ryfK䁈ۊ�w�K�}SM;z��^m&B$"�~ɉ�-��ZK_�=��46�W~v�;R�׼|c�`�A��9�u�[���.�ކ�f�Y0z��Io�׿Q�w4�z�`���Oi`�,=�%g<l�um��V��s#��{[��)��M�п\��	�;wM[��N� ^3\����d�'���澭�^G�GՌ)8�ݼ$Cm8��'�.��E�z��u�����/tC.K��wϱ�ju3Q]�1[w�K�7��6(Y�2!�W΁E5��ﲚ�����g�S�����4�K���,_]fw��ֽ2wk$���]6��x�o�qym�>!��|����Bb��9V��w�������2r�股�	�?$���P�'�)��lL������ך"�5�!���O*�0�[�%���͍Or�ڴ?�ԩpE+��X{��T���4���f�I�ߒ����e���J���y����V�Ϛ�ͱ���Dl����K���I�f��'��Tz�zȶ���eǿ��Md���G|��~0�0,"�D�.��y��Hq����W��f16"{�Q�0��	�&��k?�;���EN�4�������]��|����R�$����7=G{[ȏ��x��D�Sˎ�I�-s0��Q�N�I���k*�[>_���c�1)�RJǈSF#aВ ����p_��_}�9t�5U�ז�T*Y�f�-y��3KϊkV��{�~-��w �K:s)�_!g��CA~�j�T���`�	W�1f9m���h=H���7�&����
zЙ�u�M�>��K�^��ֺ_C<o��~9�:[.����#L��j���N`&�l���êMy6�ɫ�w���/>>��;7J �A�8�umӶ������\�w��gK�����?��h�*��}'b���;��Ҩ�e9�پ9�>���Ҷ����N ���O5���(���|��Q�,��նrE,=S�Y<�_Ks���흖W���^�xUؿ�h��@d4`PӇoA���6�T�Żk�f=�ZW��	�}'ԍ������s��T�D��Z�{V������\n7B���p�ƞŖu>�T��un��w-���@�.�<�%���޳��`��6�����v�]�2h8�a5N��z�!�)��0�,+�Ȩ�\֗)�����mY�+A"bJ�:��8�M�W�kQD�#��R�Hz�8ں@��=a�jY>��{�Q�N�n
�89iR �)K��	
xq�����&���o�<�f��E�jU�Gs|:,��vЭ�%�p.C1�{1������]ib�8��[�b9bwE1N�.S��&�uW�H=�e˯���g��4I��I��[^Xk� G��%���ey�Z�VC%��N����ed���#SG�ѵ�}�Ii�ğ�63_r��i�	f�Q+���S��]���o����?56�!��0�b�0�sjc��}`�����m#����&"���-����R+e���>{�= ��K����c��<?�x��c������4�_f��ױ�s���گOI�<�0��U�Q�͸�o��T�&��V	���<��L����e�Ux9&�t�'��)���=���Nծ�Tj4�Ι��75������XbwdZ�8�äF�F -z���d[#G�s���֓va��Qu�8�۸�
=���P=�L��Tg]������N�I���g�sBu��q�(��p�2lɩE�p<�oY�F�~��5Io}Œ�er�ܮ��f]��'{�����\��(I�$�����=q"hgiƎ�|4�^�����mIHo�����ց:�+rt}��%#��lݳ��UԽC�$5J���%�{5���S��30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�)ڜ4{^��C���p�?��|Q=F��|#�@��#(U+�R�,
�ޙ�o�ش`�Lv=Qb8��z�W��+l~���9}�H4<:3ߣpF�|�8�h]��qʵ�t)�H�����sJ��=j��P��
����+�߁˾`�����#��z���5OCP
��z��)�ߎ���m.�1�"ap�G��;d:z�H��]ң�{~L�]B��F�ɧԧ���ܦ�ب�~��C&��aVP��	B�R��_�g^��g_���.!L%����k,�������tw�2�HU�gtuJl����Ǉ�
��A��0��tIp�{֬:���'=�8J�/5��A�+3���x�����H������ᰳaw���:�՜(�]��t���q��m��,����u��6�(�=M���D��B�����c�3��8!"�Z�^�w��,-�� �9.Q[]Ii���ߢ�8T#=&��^�]MPԎ$uaƮ��MAΪz��*����s4�⺹��r$�6��OG�x1�_�y�|���O��[���l%�����	���@I�� ��׳��������7��"�J�)u��^�̿;AV���Ij6~�*"�?�"V��Zw^��1C�oep\�ُP����Y7���;4*0�i��UR����n�D�!E�s`��˘Jpx�E��[�i'Ņ���J�`?W���V�9�_Q���_�4u��w�_$�t#���lBڍS�*_�@�d����Ѡ�9K�r��g�lM���W��~����x��'t�9n�~\��H_���"��;AQ��|�ԫ]k؉&��*̷ �w��K�~�탘��e1� $�w�탖;.�ö ���E�
���ˮ�zh�k[Z���ZP��T��)���<����TH���zࠤ��1��~+b(���Z��/�7=�3S�	��X�����b����!y�&Wf]#Epc�.���K��%��;Xs��%�K�V{�
|��j.����u�@'Q+_uJ�\�J)��{�x7 ���<�Ì<��U	���z�4��VM�b�y���[��ú�|U,�:�e�'YC:&��/�߰��o�G;ļ��q�d��<2y�]\��/��4*<�����µ�	V����{�<Lr$����ZԭNpՖ_�Y�4	�	�N����:�ZXQO㞢�]S�36�{�Y�4���/0��c\{��E��ouho�j5����$ ��J���y��u�3�l�����p�J��z+��׽	�D\�0�����j��g���kJ����\��t�֛���<r�8:�4�������(cA�q�2TqT��Ik��60¨��6�z��_��q������C�����K�))L��V�6�Y�����!/Z�X��o�('vKa�fЍL/���\}m5%dC�f��XQW}$3���]I����@F�˯%W �>��w�k��YX���9�y�y��������5c�^!F�-%g���g|oQ�/%�s�@� -6�.i��o�Z���}}[H�fz�ǵJه�������*�*�Su�!���:��f�qzK��x��������?a�K*��B�8��!E�E6_�9%�M)�� ���;k+R�^����{N���R���_/P�^�*�g�G��D�����H,�,�m"t�4F��)g���l��������z-A���YRt����æ�S���]/�#A�"Ć��@�"�2���Qzp΍;��J
��y2����(t��AT��S��#/mʬ�,~��~��6@��(`$Mh����f�Ʒ��ʆc�xh�A������V�:ƕ�ω��P�ނ�1�缿����3�h8�Ϩ���φ���cz�!:�`�h{����j~�܉�W���Fn4c�M(�6m�ї���	��:��{�0���#�d���e6�2\H�1gyQǐᦇ1�߄��UL�m��E��&�a]4%o��(\�����"�ԁA-���H�,�p]�
�"��o/�c..�p7��]����c�O53��:��� ��DOB�e�|7��E<�P�-�~�Db��G�QJD���ǵ��4�6�D�H���>�:8��V=~y�Clob&���-���L��G�;������c���O������pgw�=����>�o�Y�<uK��.1��芐\����R@J�3-�F��KP��&R��]��v��" �y�R#��d0L�����>����%˟�[[� 6�� l0fy��:�k���W�Q��>g���qg��+g���y�3����KM�����Sg"�T4̚����a��7��`�
�TS���ص���pdǫ�-�J�n��`�3����@Q>(��CVr��{�-jf�򲐥�l��rOMd͈�B����vl�̕!�k�(~�e5CvNõH'�WYdV�U�w�CM��m���ۦ(A��:nO����2�!&��P�2s62�z����
1�n{��S�U$��9u��H����i���9EP@tIQX�@̿=ʕ���i��Ƚ[��y0bZfn����"���~��W��ZM�,gT�fG1�oo���?�"Wʼ�>rN4k���7´|m/#��y�o1�t��j��Ɇ ��IZf
�9|�O�!��&Z����g�zI67��I�.�����~��{-#*�$Q��֎�v�lL�_���0_H{�'��#;M���QpuS�@4(��i�#>���0-I�U�����l#!����&�k�V������W�iϫ�o΋���@�X>�"��v�v��(;*j䬞�,����m�܃�j)[�h&:�.�7r�4�������v��uUЪ�>+֟�꣱�L��T܃�-x�D����)�>�#]@cP]r�om�5�V�9.���f�A��ݾ�� �ieOZv�J�����za*V�V��t���*�ӎ��e��*�;�7s�m6@?�?�M]��Z�]'&Wp�f�����L\Snm�A?��D�扑~�ж̟̉o�1 iL����R���< ����!�%9��sy�^�T�`ƚj�fi�il�-���l��v��tYׇ�� �Y��`��1MxO��E��)I��ͤo!YX \�%��e����wWQZ�lR;�_�Ϳ�ߒ�ҟ��؞d�b�3>�(�a^Z	
V�7�l���_[��{�����������y����8�*��٧|B����t�YGc,F��~%���Vo!���h��{�0SPB��`�[�(\��Di.�X� ���?z�h���	%��[�M���f-��f�l#5j>\v�h�h򤍋�;�X
tY�)k�䋦�_e�5m�����R|���U`]����$:v'��5� z�s���=Q/��;�۱a}��'���V����IA��������ޝv��/�yN4�͔�.����#l:nf��U
��p]v<7[΅��eƧ���@�qY��à[�H�,���`�)����L�u���J5.��;�b�Z���+*�(sp�����b��oin�mEw�S���-�*�W����P<&(,�S'�
Rݥ=��wo�|}��Ɉ��ɁQD��u���U)�]�3�i���7�?B��Q�0��b#
}��.�+9.�,AR����~�n�w��8����r+��ݰ��}�<�i�E�F�-�8�]!]4xE���)������s��h��Ȧ���E�qz�縐`�2����� ���7CvG��y\�H�����䓎w1l�/pXI����5z�K��C:F���~���]h��F����zﰹ�U��p=����
�BZ���x�'#�F3�	+�BBX�PwQ-ޠ��yAs�/�!�g��ʻ�mZ[1��#e��5�0��2�r��}*�ZP���cm�2���?���>V>�GY/2�dw��ۺ_��� ��"TY�8uf�ZGN��Ll��(���!o���5	.T��x�g��*��������#	N!��:fe���mh@r�J����}�c�Vj��/��}~Mߛ"sS�����i��mŀ'{kMs�C�7����Pjy��-�+Ԛ����M�b/.CAn�Ղ����c�O=����>�:W�0s�b��A�ft֪���A�ݢ�����o�6@I�l��{�J Nt�B�)a�SN�{-��Q�Nfw;~8�üs�7��[� ڞ�c���dDM���/�q(�ymGV�pZ�����c�]�������t+ҁ=�=�~_U�phxX�y�_X"an-��u��=`�$kϱ'�od�н��>��=��/�xܛ��{}f�$h\�EOF8Q�lw��i��u����Y��z��$ꀉ�1���Ƈ��U~������X>46zf��\B�h˾]U�zr	~�8cc��N߯��>��y�y�)���vP��C�&�܃�<�:ͭ�q�o��v��Ŭ<j�k��t�2IqiR����X�je�wn^�v� �M;e �2����"��D����_J������k�����M-0�Y���|�YwB�E��.16K/X�����/�<��G���Y^�ʞ,R+�l�Vz38=�4!A�`ܞˀ�r�����:@��n��lV3Y|O��d7�5�DLV�F�N�du@�zMe�*��*�`1�Ꚍ{M�kd���Nz�%O��GJ�~7ah>���$����DU�v�K�%��6���}��]쓻9mTxz�o��<����0W���5�Y��e�N8�$B����EO����dkٛ!�ܜ7�ND}T3т�`S3%B	��I��*�� ���� }ꬄ�uUH�����#�ͮ��:���h�@���".�u�i4:���GMU�F\�O e��f���g�Ӊ�r��t�N\F��}���O��_TJM��h��j[�)���),a\�(������m�͎�+�����d�)�{tn�O��jrLz0�P{@9��i���ʛ��� $2�|��6R��n�l�����JU<�i-H�
t�IR3��5K���!(��jc�dK�:�5���kO����۷1d8KGFj˧:�;��|�M�B��Ž�`������p�T	�ڷH�)�o� RDv>��8i��GV��5�|��E������yc�t�lpjkD��l��k[7�0^��O�>�x6��TTkh
���O��|E�eE0i���px�湝W�
�I�i�R���׳��EC�h
�E}�!��3��Ԃ�����F>�7$d
��I�4,�s�M=G ��$�[qGJ���gY�L�\���,�x�ѧ����̝�ۆʆ)K�M�,�"�:Z�«)|���EO/J�v�x��ҝ!
Fim���Ux���EbU/
�^�Z$��%R���xHMҥ�!7c T�%3��HlV,��M��E��.$�R�q�ɯ����kTϺ�>�,��5�f�߾����[Z�)�{�<���U�>Uq0�X�J���CEԙ�����k��*C߷�|=��?Á4�3����X���%b����7����\���F��rOJѣz:Y�Hc�o�� �rؙ�B��~�7F�C]��bW:�,o��ML����Z����Q�HL��xLI��8k�yp�Ta��|"�%����9�[C&^�t�u���L�OeF`a(���7,3�٩���Z;��<p�1�^�ӱ� Hj���sH����8v;o�1�Y�`��:L��)�V��H��m�2��rP9J�Ԣ��>�C&!�eq�r|��)1,��*(浪p%\���W���۴`)S�)���a������n�A�T����k�v ��2l��i{�?����h�m�N	VR	���;�͇��ގ�'�0�o��߅Ť��~V��};2�3h��u�����4]Q�`n�p�e(����/a�m�}_Us�1^氂����h�B��|�`Շ
��X��u}*�`B}�qO��lNvWvI�#՝
���o�d��"��K'd��1��W{f�\钶�pO�븧1��t��d�&�	T\��0�յ�쾫�S��1��vL(�7XP�}3�i��mS��'8��"�D����s�,9���b�7�&�k]TܣF;��D�&�otb�-=�(�d�	�r�ST����ת��˷H���Z���ٻ@�m?r�X�d�c�[E�#2Ţ̱����$��5��?G;�UjP|�*�A�\ZW7��[�	q�!5^B��=��&�䓇~��h__�~�Ck��~����sbNDt�w�&���a�8@�WW��Ā�P-!��s�3�4	b�/Vi���	M�(�Ƙ뀱(�����>�q�����һ�%5M5M�P���W�׿'i���pŸڞ��?}���1��6�4��U�1'>,+Xy'�#�|�Oa����4ca|��� ��j䥢��2���fU�^y�F!�ӥl�R����˴��)���~��sS�p��Q�7���j��UR�w��b�;�̱Ε&�f��E�o��k�cZEß�V "i1�p�2����Z�bgjf9�!o��'�@."	�!�0�S4���ө� |����o>��tWt�Y_� ��I3$�
�|yn�!�� ���s���,q�7���I
���V>��/c�m�>#\��$�q�@���^��ױ5�b0���J&#m��su��4�,����>��70�\U�6��.6�!m���L�k���湣��S�]�C�}38�r�X�T���a��h�0��L;��U�^���^��Zf��*)3hr�`�prY��䠦T����v-��UB��>Ⱦ�������⃓,�j���&�y`.>��%#O�P��o�2��p9����މ��"��p���a/e����2��ܼ���P*�*1��O��t,Ӏe�e��[*D��7%�;62h'?�����E�"W�Z�*y��QL�tm�?!e�DLf�0V�Ш�z�+�ڣ�L8�i�Dx��>�齀c�����+���-�^K?Z�Ohj�����������S��>���:+��n pt�R_���x�5kEL�;r�����7� ��%�X�Q@"���Zc"�;�����.4{�\৞V��e�'(�z.Z�Q)�)�Kl�ю��޴-����ధ�p�����í�8�:M���B^�)�?׏Y9�F�ɬ%/ֻO�oi������>S7�Ҳ�[H��\6�,��� ���?���hGi�	�[IU�?������l��5���v3�h�
_�}�8��YP�o�A�Q�5�ޢ���'������K̓���('�?�R��s�I�=C޿��I3�a����]�򪈧=���cخ����M��v:�g�kg�� v. �2�a�L:��R�!���<lCv�j�[�%b�'m�~]�Ў3�qKt���H.zS������N�������M��V�b4Pn�&+�*:�Ibڈ����bS��o#�n�Zrwߓ�	*bwG���.<X����[ℼ��/��w=-|����:5k��GQv�#"����*)r�~�"���ޕ{n?4KFQ�(;����#1�r���C+k�,�9�1��p*��%�OO8Fs��8+�����
}~�.<��tw��F:�h8�N�]&p�M�F)m���M�s��<J� ʍ�עtI�c����`8~�]�k��դͿRC� �+q���&�(��<1��pJe����z-��������\!~�]�*�Fa�G�l�E��#�tZ��p��
�ԓ$�<����F�@�+��NX3�w�i�m��A3M��
[���n֤�m��0���U��h7�"�2�e~�#���п���vmGhd28��?���>H�G��M��@���;_눮��E�z7uTM�uXKDG�-�L�:�q���
��!���⧍�T����jN*�%B:�H[������!�t>f�k�yr���M\���B��!vZ��`o�K��Щ����������M%F5���4/��+�_-�
M�Ђ��I��b� �C3v�մ��R���列lX�l&<0�P�b���3��t�4}�B�Z.xݔV��I�|��	5��@;xe�ޥ�J��G��ka�c�N��-'KlH��w-�N���YΩt�[?0�ڐ�c���d�����!�W(��GȓLp3�}�cc8��G������t��=��~ѻ�p�]�k�:�Ga�|��'?3���=�?݇٩1a���J�c����c;/�>���Bn{�p�$�EA�/��Q���ih%�ۦ��H��f$�kT�#<ڶ���u�Z~c�ߵX��6����آB�s������	%~���c��!�:&���\؃��y����))Pf�p�>L�u�I�l�\��#��y(��c#jV����2��D���6�j�o2w �Fv����5 R��2��w�cnD� ��@��I��]K,jׄ����$� 4Y�D��6ی��m1(x����3���5)G�PXY�ݍ���A+ΦE��Tp3jQ4��|��@�r�R�'�v���@ks6�=3�k��9��sD>P]B~�Nf��@I�uet��\��1]��>4�{������A�b����9}��J~h��O��*{���ج�^�K$���2���E,���9��xl&��6����:�L���ㆋ� ebװN�顯���~��k�=:�VVSG㜩�TN��3ÖE`������@i�4�RyP�fY������7��Q?50U�9���1d�@`��>�|2�'�('#{@��sĖL���=4�pա�z9�a�*��F��>�9^A�����������~/�v�E��S��F�.�u��2R+:�l�21O�m�=v?�[1>��*��/V��_B�q<�����RH_c����Ԍ~K�bv�ޘ����	���bE���W��*��YӴ��M�b�o�)n��w)�l�:J*���|`<�%6�v�p���]� �wN�B| ��ɋ�kM�Q!Ԟ^�o�])c[$�e����掠?�ȺQfT?�3>"#+0��_�+|{�,�G�ނ�y�ሩ�uˠ�08��g+�i����}�<%pGF�18m$�]��^�)��0��2&sS���ļ�>�M�s���Tβ�*��`iC���������^��C��l����}E��7ln�6P41o}�p����d�z�&���y\���~�*,]^'F�E��X����%���A�D
٥O�5����sF6�+_$X�evwt>�A��Q����1��j�z�-�AmI��Wt�|�*��{2����T-�!���C}@m؜{2��?kX�>9:!G������p�_\�lDͫ+�T�*uI��G��RL�������{��!2�)�X�lT��*�[G~�6Y�yT.��	����!a��f����l�ru��^�4� �ۮY����`��@��߾���s~�yKU��1*���hMv�G���բ%��6���E-�&����z�Sbc�C�"�E�?�6�Һ�����}A_0�Ob�uǤct���.�6�+��݅4�Z<δ�$���@�檉o��JC���Ŭa��N��-X
�{�w�K��6E�Zd�[7ځ��c�b[d���r���-�(NrGy�(p�Yn�cI���x�����et��=��,~���p��\UK!�a��x'��ts�=#Y��ڻ�R�R|�,���#�@a/]{�^��{��$랜E2�8�v�fi���L[��몲��$m�Q��|�	
ە��~�:��&�[�*6�ʢßD�B����sl�0~�cf"��L5���T�T5�y�<�:NdP�r���z��;N�����p�J���xj$�?�`�2L���f�p}Sj���w��v����	� ���2�Q��|mD�3��z���Nq+=ń�_�\�]�)Y:�?h�9��5�1Cv���d4�?�pG,�Y!'��Ohd+����� 3{�4İ��c@	��)��%>x<@<�����3���%�N�8��D���ɱNa�@��ee���mN 1����(T{e��.�?��7ߨ���*���w�h���'���B`�9�.K�z��(�ۜ��V���6�k9p�x�fG��h
���_�*����d�� �e��N;!ͯ��y����r���MG�y�d����@�NG��34�V`��H}b��L�I�;��m0 $���&���u>Ͷ	^}�Y�T͑��:'���tp�C��ㅪ�u[rl:��GКF?�%Oc�Я``��g&�O���,\��w}��|O��GT�>��
���=�)�:�L3�\xr�r�F��1������`��)|��n�;��0{z#W��a�O��k������x��i	[���0��������U?�G�C����Ll��	w25.�y�P�v��jf�"K�~�����?p�gH>��)}�t��8��j��{Ϟ_�|�y�ʈ��Hȯ�C.���m��H	�nH. ��2L�Rg/o�j��i�]�V�<�5@�������і���Vc=���O1Ck��lWx^q�%�K0!e�O��3x����HEk`��pAM�ꕻ|�'�E�B��>��x(=�:?{
�L�i��H���6��E��
���oK�����jx��&��Iq~7��D����l�a,8poM �eC�K$��qJ�F������B��r�,BHwъ�X�@�4��;��_q�`������>y����6J�����qԽ�����Ykū���J��y��9�	�X$JӁ&�X�S�%��0��s���෈���nr����!:��1�hk���r�]z�C�~����^���':5'F��jL/�6�~g���}��l�e��B��R��ρ?�1a]�8"�S����9��E&���s���O�]xa̅��[��3,Nr��1;jE<����4��Ո� �Ɏ���HQ|o�\cg;F�}e`��;3L)����V3��H���m����lhW9nJ��p�كg�q��ږ�����%���U�H�pI�𢐪9�Yg��S*��f� )�:�e���&�tAa׀�K.��͊VP��@�I�cw|�3��m�xV�lc�!`��q�0��D�ˢ���	�����cVHk
;V1Phy���"�؍MQѥ��'(���D��8<}q��U�ϰ&0����BV�ϡ��D
T��|}�C*B�kO%��N5�W��G��
\�o�ckJ����d�H?�U�0W|s\]۩%��'1HD��0*"dh�	x1��Ԇ���5��O�*^1���vpH��|u������嫾�T�FE��v]�wuД����U�y2�Jz]��j���=)&�WY̯=̩���	�	�r��Sx��図i�����-o��ʿ[��@��r���׈)ʄ���#Vu��UF@��mQ�H���ci�8��P�x��1QZ{�����q�N3^�Tc=�C&[������c;ޢ!�kZ|j��/s�t�a:&���d�8�?W��71�!
�;sg���X׏���P����M>�4���ۀUm��u�y<�q���j�仨��M�|ouW$<�	']��[f�BE]?�J��$ō�(>�4u)U��g'�ˉ,*��y�p���^:�X\�5��4���o��g�����������\�!FE�T�IA�R�>��oB�M�A�"�sw/��Dq�[��܉��d۸r(`�&/-(��j ��4�\z������z�0o�g�B��#Iߢ��?*z`�j��_���-D�.��j�B^>�)gBT�rU�j�y����z/����`������ IipYA*`�t�~�<AU4�.Y���d1��'4W�|�ig��W��;�kL�6�OCI�DT(�����۷E3#b'VYPV�}�R;Cz	��ŕ��tT���9��^?�PD@uѥ��[�qA>&�A�Y�]��Hl��*�{0�����X
�n_-�B�ќ��;�����}�m@��y�O��)�=h�\U�z!�r����:�d����vG��U���>b�l���9�rfʃ-[�D����c���@�>^�O#){BP�Xo9�Θ��z9��ދ�@���� �T�Y�Q����l^��/�l~��r ��	U�'%S�9�.�~Mh�Y�ߊ�wH-�-�<��J<����Z(A�� �13�|ɡ.p����e�W-$u$N�T��.�` ���E�:��U<\lz�	�[���޷�������z����Hoxzq��ߣf�{C�+S���R�P�ǈԗ̤�=�XC�F���b n��%��y�f���E�\.EVɏ�{���l��\�s�|h{V@|�H.1�Z��@��e_f̖�mF)�{?�# 2����Ҍ� �U�da�]��u���t4�+�yb{$����k(�U�����'j.&�d/��˰}�E�L�.G�x�м��U+D<C��]���/RJ�4��]K��s��	' �ꁘ<]6��_S�_f���������g	�s�N�H��'	Z�8���ol����ě�{Zqs�ç� ��t"������=h���5IW��X��ϙ���0����d�n�B-���JP�+<V=�ڔ�5�~�AZ��vW�Fx�ݳJ�[���\��<�ǆJ��q�9�����*�s�6�(�wqԥI2E���݉I�ڽ6�T?���m_nqS����C�j����K�|�Ly���$�ʆ���5/K+\X캷�Yu�K��������4q`\.l�%5Hf�{SXbj�}�����I���#��|��%(6��/X2���C��)�R=����Sd�K>����c�92��-V���48ؽ3Q4�q�$Z���\���9ᱠ� ��}�jf���f���X^w�⫶{�*�ƞ�r�M���f;�-K���xp����,���a.`��8����U���}�
��>ދ�13�l �ReT9�u��g���,4���0�R��0_@$^��g9���H�Lae�,q�x���
tщ=�� �gN�l�չG%O����A�J*@t��p��E ����ΒaL/���A΁*��s&R��Nk�\������+��s������'(+L��r.U�s&��M�m[%],/�w�OqB61��(qu�M��J��`\��D~cM$O�%_.�t��&OwU��-�S�n�L`z
��C�UqkQzpO�����-&����_�(���ԡʐ�����[��/��QLik�Z/�5w���c�Y �x��6��.��k�^�Q����eÅ���n�:�[w����&�t���4�2+���̲��FiKn7	�S(�]��X՟�>�ȓ=�i�L$��a�@���ڃ���t��6�֥i�yQ�!lZ�~�� -�"s�W�B_�sZ���g�Ef��to+���{��"��z4'���s,�|)�)�;cno�Aft��&�c�� B�<I�h�
I�|��.!�
���=g��6u�7�x�I�� >e�(Ӛ��#�F$���J8��42��>�ǒ0���c#�Q5����uЛ4d���%��>��0�� U�6¸m�!7�t�VF�k
n;�p���a�g*b��K���Xz�B����&�l#�;fe�h8%h��ׁf�ܿ�)2hbIα�mr#v)䪱��
D�v�� U7�>�>��u!���{��郝����͋oY�C1�>���#�GfPa�o�X���9Hs�hS�}0�z���<7�eEK�ZC���%p��;m*�ډ�t��2���?e>�g*�^7/b6||?>2����:�+�W[��"}����GL�mտ?���Dߛ�:������h��m��LB�������JR���hu�/T�^7`�@-j K�hB��i����݋�e���K��ÐF z���I x�,EV��C�`��]�� f�%����o��?UZm\�;�FG�{�[���ǟf����Z��
�(���Z����s�lG���}�7W����Dty��Y��ͻq8�	��n�B(���I�kY���FJ��%�t�Y:�o]�ց$��Ʒ��S�����0[�_&\ ��%}��/ dO�?N�hQ@�	a�K[�
��	�e��B�l=k�5&��v�zlh�K'��#	���Y�� c���4�5)?��R�^��5�x����'�&+��,Vsݜ��^�=��N�-��a�LԠc���N!�RmS������v�;g�#8vD�׵�p�?�.ʍn�km:I�Ië�]�1&v��[
E	����HwoИ�4q����\ �H�h�]�{�eNg�[A'ޱ��w<���b�w ��C�*D��M��Fz�b �o%J0n9c�w��q��a�*l�����<��ۏ��ƋO�yaIw��|�]��D;�Dx�Q ���㫄��S)�J���v����ޟ�Q?~��Q_ú�L�#;<C�� +��	,}�I�;��úEE�n#��e�8PBQ�9�+���V�3}��t<���S�F>8��+]pٔ��-�)7�1�W�?s,29���W&�׬�֭��ߣ=7`O'�g�<�\�ɤW�C�!��5~Z֡�߰S2��&u1('�p��Z�]�z��8��Wx� �{~n{�]��=Fk�˧�G���R�>B��z�
2����@Ȕc��F�+��eX�3�w�{"�wHAN�R�/@�%��#.5��Pm�?���A����l12a�����������m�<�24?��>�pG�FȠ{"��f�_5�B=�\�D�cTֲu��G
! LV���{�V�T��!+E��qG<TǬ���������2��Rf_9!Z�f�O�)j�r΃���#������ϓk���9�<��XN���8��@�}�co/M/����՛R��F5�1-�\e�Z���0bΦC}���>�����3?��h�����0���b��x�}�t��RG�(�d3�������Lg?w6@�3{�hʷJ\t���vaٳzNaU�-���R��wwa� �sT[I	
���cq�d�s��Z�k(G�&G��tpv�Ǖ�c�œ����cftg��=���~��,p$Z�����Ę�a��(�1a�M�=��� �����H��-�����/6L��W��{���$$6�E�W�����irF�%^�IA���r$�V��m�ڶ���?!�~moY�����q�6�����-�BW���z��̶��~��c��l��|ү��؍Gky+��˳ҚP0���rdܿ�h���Q�S�؃@����j���ɰ�s2���6	�i[j���w*$v�}�	`c ��2����^lRD�f�ğ�S~n���F��F��e�=6�	Y3a��ꌽ�r1r������k���?G��)Y䊞h��+�w��CG�3�U"4]qu�O˼�)���.W�z@u�����J3�Ѹ����NDD�D�X�N0��@S,�e�1��1'�ŚHNT{>t�'s��5�����ރm��:D�hz(>��.�����2`K����4�|���8���M9)|�x��4������gd�D�������ue,V�N�A`�`�p�� ��o��G���D����ɜs7N ��3�`�a���JyID���6 ��,���5uC��"M������(:���y���u�^=6uT`):��MG	��F� �O�Y��H�|��g�^�Hex����\_-}0��OY�@T�!L��x��b�)���e��\<�K�ں�Z���ݶ_�c9��)ufn��&��zlU�7)�����S��͊;��
s��:J��g���g(���+D�U��i����V����B��5�y���жd�j��K�1S����0"z�����7���@�8��j��|�wq	|����t,ā7�圄��R����ֆ	��'H���+�mR�$&ģ+i��Vh�5و�;ʯ�n��ʵ
��YcvvY��k u�l�q�'��f�0m�O��{xˣ�z�k�4F�	-���p|�]E�3��WvxaPc����
cCi*3Ҳ�W���WE���
����QQ�o�ؠ5$��"�7`� �������N,q� My�#�f�$C�0q*
��>��@C�
��,{�R������,�W3��bk�9����>����5�uJU1��9�:�V&��Jh#k�Έ���h� ���r�ā�a����XXue%�F��	󘭁z��'E��-�rl���`w�:��e`�|@.r��v�~uO�`T��:�����L(&J뗿���r��Oև��ˌI<����}aV�"�̔�V�9��&{5�F���A}Obm&aŐ�t
3e��q<�;��C<-j���&CӮa� �r�N@H�R � 3;�������J�fL$���'VLx)H���m�s���09+��)���@TCjSٟ.�	����#횴�D�*��o�5�t�E;��j ��#I�k
x��|�PF!������9�ŷ17cqI�0��O�|�ؚ�BQ#��O$<�O��ou���j�Z.�.0*��R�[#�b����u�P-4�8M�ty�>�"0��U�I�J!�b���~ky�c��e��z��v�Iζ���˹�X)PT�m�	�!�;���x;���w��Wғ�P�9�n{d)��h��q�9�rR��乾���v�x"U�]�>a;��kٱ�%�����MU��t�>���>]�j#��Ph��o��J�!߀97 ��7�t,� �	.ߜ��:eZ_i������~��g8*��lX��8��9p�e��f*==7>�6k'�?;����򨣏W�u|qUѣ��qL'��m���?zTvD�@9��'�aM��ڜw�LQ��}��ޗ�_���Ѧl���z~��^D��+��j@�7h0��E�P�*�h�{������- �Թ�������x:K�E����Ɋͯ.��a '
@%
�9��S5�b�UZ�o�;j����к�'G�uR|��u|��M�(vbZT(���l�����l�F9���������5��\�8b����_xBW���X[OYr#3F�]%���課o�d�suH��OS���4[���\�N��;�8�� ��c?}�Yh`�d	PH[j���S�0�Cl��75u�v�҄h�J��C����fY�Ѹ�/1��
��5x�����'��$�p��W��*R�o��'k��+y5ssZ��~=|�fyh��oa`X5��8V�ay�k�����`Ȯ
���Ʒdv����$��I�.��#�zGf:8��z�ĵ�v��[y�^� ���w�Ч�q�QA�+��H�{n�������	l����������^b������N*�o��흕!�bL�o4�n(��wq�v���S*����cV�<1I۾C]���ۥhy`w��|h-��� ���xQOm���� )��2l=U�T�r�.Р?�2�Q�U�{Z�#J�����+Ē�,,H6���*�)�{�F���W8_u,�(~�+]�^�c.}��<mTPU�F3\�8�Y�]_�Wʦ�)�	���s��2#вʆ1׻�q֜t�r.�`�Y���B��B{��©C��W�D�+ų�����~pt1���pRS����z&+����E~=*�]SF�F�6F�%s��N��m�ы���
!�^�}N	�{;F~T�+JA�X됇w�� �A=n~���wԩe�
�u5xme
U�����ĩ �[?20Q���K��i��ۋ�m X�21�?��>��aG��i�O ��a�6_�
�����s�T$�du�G٪LLcڙ
������!z��J�T���-��~����4�5���n�!���f���8rxr�����kd�h=���am�����t��ZA�����q����M���d��Ⱥ(CD�-�d̚)$��}yb]\C�DsՍY�K�����F���0^�eb=�A��Mst�1�vB�s�=������ȴ����j@��Y���bJ��Ƽ��a�8�N0x)-�R���nw��P����΢�,[X˄��
�c@��d//e5�6��o (���G���p%�E�	c��W���D�9��t��=�0�~ʩ8p3Zy������aY�����!��Ed=kt�^�_��2s���܋�ʈ~�/���ܦg�{�01$3t-EzW�ܽ�b��i������d�(��C$�3��\ƶQM��f~�;��n��c��6妩�穤BF���IJ}�e�.~8t8cKX?����^w؜b9yn˂�[P���%}��.�<�E��܇�ؒ����Jjlf�_��2��)��n��Hljм�w9}kv��P�8F ˰2DA�����D�Ɩ��v�bvj�����	!�8�:Ѥ�S�>Y����U��̂11a9Z�g����懘�Gg�YiJH���I+�N�2?�3�K�4!�櫹9�+Li� �X���@��}��P63��+�m�����D�W�}�N_}�@b��e�	`ҵe'1�����1�{��lvv1�:�X��3�r�
�	W=h)��o�.�e<����jK�>�^�#{_�Vz�~��9��4x%)>�tق�R�S'F��n��o7e�@�N��ٯ�/�ޠ���Vw��6^��.��"aiN���3|��`^����¨���I3r��/� l���K۬/ճu`��Q*������ټ':o~噼 �^E�͌�u��V:�"G�>F���O������Po�gn�}����߈�\�f}�HO(E�T5G&�;T����)�a�W�\K�{�G��Ue;�y���4�)�@~nL�>�5��z[A��d�P�����<֨�+ĉ�
8���[�j��&U�(��u����.�Q|$5vc������Sj��K^{o�@^��_�ί�e��}���86	jX��S|��*Đ]S�lǷ!u�[v�	/h�HvB��z�]R�Ĳ��id�V7�5�gi�~l�����Nj�c��k��\k��l��>��;m��0i`�O�AQxڦO�Lk�7𸉓�2��|�E;(��*1xp򁝂��
2t�i��V�A��^5�ENX;
����< �K>Z�����ґRW7�:�b@��x�,���Mh�����$�3q�yp�F���W�{�9��,�Ud��c羈��jP��3�P���ܫ>���D��JDm�`��������k���۷O����]���j���5�XL$%N�s�x1h�ІD�Ƚ������
�r;�~���:EUn�ZA��+�rD�.q~dk �/�!�:}�;�'%�Lw�����	��r��+q�d����e(x�	�a�`*"4�~�я�9�&J���e��0�Oѧ�a<����3t�p�`;��<�{C�|n���� 4%��8H��"�Y�;[;�������Lq\���V{��H�Xm�KRڴ�a9����7�����x����v���8f��S�p�"����k���Lh�SIFc��5�qH���E�n��A���7~r�bk���4���?������{ixmSm�V�=?�iZ/ɹF�R����˲/�"i.V�';���h��ćT̰ �%QLߣ\F�(�nu��s��}KD��*��n�}�G 5B�/����v
�,��g�}��B��Om"N}DHWb�&؏�
��o(~��i��;p�d������WgC\U��\���W~1�o��x�Jd��	����,�!�$����r�1ύXv��b#b}��z�U�d�%�Xݣ���о�]����B���Θ/��]@(C��0��&0DUNA)=�I���H	S��r�OS��J���Ǫc8��4k��1������@�Cr�:
���I�G�N#��̝KK�9����ī��%�P�!�--Z���G�qD�l^.��=`�&����Q�T���-�k�'�UsN�8t�QR&	���8,��W�?��!R��s��+������O����M�'�2u����PC��IqI �ڲO��M!x�N�ml)�V+J'U�e�ܣ%ڊ�?�İ�l���pj�4�ޙUF�'*��,r�By�_���;�p�}ȕ4OOz�8��Ư���;������
J(�F���ӑ�FR2-�۷�ܕ�0�j�ms��	`���5e�V�x,� ��`��-g�5첚^�K��]�\����z�w<ٯKAB��@#�Af���Yz�����I��s��v�+cOB�?g�q�GT���zr�L����=��3m���p���� Y�i���*������A�
�.���-��	��W+7"i�����f;�`Һ~S�C���D�x��=��ǭW�,'��@P�g(�J�=C�8 ���"��T�.��0 ^��.P��-u���}A�媉�[�������r1��*�t��{�D�x�!f�1�Uj��M�[e�-L5�%�;K��(��N��I�+Ո9q�ѥ�ԒB�t�o>�q��7cu��?^e����ф�Z"V���@�";-���ڬ�B^���C�yNp��mԸU48Y�G��V0l��M@�sf�& ���
�+�ݥ)�J��1�����0��!�:�y<�J�(�W�dVc�'_	�����-��wҜ�$}]iÇ�
l�8=���_�ŭde�^�m�����j9��L��l Z�]���:�ݹi��0Ǥ',
F9��2~�� �ɊgZx��Y�ܛ�4�B�ж��A����s� }(�C3�ǘ:ʢe�7�$|	�;_6.��
 ;��E��ԲF-1���z !8[�D�v[�W'���8S�G"0�z�
H�ez�K4ߪ��b�?+x�Ԛ���1N���?��4�XJ�`���Tb�5���e�yj|�f0
E(�.l]�Լ��*�v�|s����{�{��|O��.X�a�@�1�_-B����)�ͬ{��q y������	U���ΩP��Z���@y��5�o��r��U��]r�'�t&��~/\�+�Ě��sj1G�W�����&u<��]j�/�#s4��ρ���z?�	ULʱS�<A�Ꮎ��ƶ�d �����L	��NI�=��@�Z/��V7\���؆{aSZ���j��w=��|[�'Bh'�5p�8��Q������p�������Q���S�?FJw��+Cf����u���"��@@�`2����ZC��J��կ�+�\}��������#O���;��$�H ��O�(�q��f2�C��1�I#� 6�n�U c�2Q�_u�Oq:�u��~)C^v�K`�LL7������js)/��X�}Z����K�/�E �[/b\5�%��f���X	�`}7�u�/�IF��J�ē�ia%������/�L��/Y�nHU�1��z���Ĳ�8cqH��|e-�t������Q[+"x�؍R�֥���l�'- �y��}��f����my�?�>Cb�]�p*y� ��&��^fb�K���xWz���c�z��a�T�z��8�����s��]��-��Ib������X�R̝ܱ�+��Ɂ�3XÍ��YRa�_��^9Pzg�}�菎���ol)c,X}�����tx�)�i�ig���le�{�nҹ���iAf�~]tJ�+���{�7�A7�ιE	/�Y:A���`������� � �	���E΁���ച���Ł(Ң���Y�L���v�m�w�,6<x�6�U6�l(��M C=��ͫ�R��A����@��+IZJ��9�?�oh�_	oZ[;����D�Af�l�+5Ƅavoz�hw?�g����-Y��F�@'��;l�5�j\�� ��e���������q�'���|��s}�
g�<=-<��8���)aqP&�3f鲹��Lbab�����ۢ����v�O~�U�P�)K�.j����:�֬�K�Ħ��v�=[��ֈQ�|�薉�8��q5>���{�H�X	���������Q��Ц*����Ab^�C���+*�k|LE��e�b�Koŝ�n�*+wB�f�s�D*7��uA<�N6�/�u�f
��bwgc�|Y-����䯍Q����\�Hl)\R=Į�E ��?Ow?�iQ��ǖ�˱#�o���?U+�Z���'JJ�ӎ� y�{����W���'�ta)"��gH���{��u�Nna���q�����%&d�۳D�2AF��>޼�o�n��S>���d���Z���Ѱilӻ�cl@F:�j����)��35�;��ϟ����{Z������U"ɼ�вߕ�Z^*gfH<f�);o�v�@O"i�b��C�4����	0R|Wn�Q�Ao���to�����k X�VI��
�	|�iW!=�i���{�֌,7
�Ij�䎶�y�u�ͻ�#�[
$#0^֠�O��|=��:��m�0qFt�yq#�ߨtn�uec�4z���Y�>^�n0?9yU(���v!ͯ�����k "��Fݿ�)�Ͻn���:�ҜSX�ϊ4���Ȑ��B�O;����r�~'�W�r�U��)m�hxiı��'r��'� �Q� �v��U��#>(�k�L�E>�xR���ǯʚ�EȌٿ�>$2w#��UP�o�o?B�h�89^W�>�e���J�Rye��`��b��8����9*��2�So��h��܀e��*�O�7�jN6���?���~��on�Wq�I��B�^�LnӼm�_?��~D�ER��!a�(�^O6��L�G�_!ޞz����3%��(P��^�.��r*;j6M�>�������6��\M�Y�f Я����T?x!5"E��.�Ʉ�6#��� n<�%1'钱3��I~�Z�m�;���Q\H��CL��ۚ��'l��D�(]:�Z�꿉�Bl�h1M�����&�$�$�r��#��8	��k�B�����Y�CxF �F%�U��-yos@���ź�M�SbRN�s�[��2\�͚{���C :��?��h���	w��[qj�����!-lS5G5�ve"�h-�\�����J�Y�|���8~���M5��/��^ db�K�����̅�6�j']�Բ%Pss����=���$����a'��y���輙���<��ʵ�Q5��GUv�c���3i�_$�.`����:_�QÁ^]Ĝ�vNvn[ �5��g���,���-q�)��2֤H��7�Q��{\�1��G���\�����^b�� ��
�*��F���,b�A�o{�+nOBwx���i^*¢��
X�<�G�%K���,����w�?�|O�:ɚ�RZ� Q���q����)ҕ�sv�;B��f[?���Q5l��O#�r����+��,��ޑ2�����DB8I_�8�nX�O�n+d!n��*}�.F<߁��F�?8��l]�F�ʭ=	)�Ǧ���UsB:�����e�0�����y��`����-�r��-�]CH��싌��z߆O��e�h1~pBp�T�3�z�s��U\�DO~D��]:j1F��4��,عz=	��I)�Ъ
H٣��(�����FE� +�2XrOw#����uAd�������yYn�]�m�&q�\a���ł�N27Y�T��0��2�m��2��?��]>�j�G���6 s�(~�_K���`�ڦ�Tk��u�YG��L�Y{�ѽ��jL�! ��]"Tu���u��U�Ũڵ��UGur:!08�f7�3�(mr�����_�O"b�h�ѓ������m�heNZ��w���f���<M�q��v��qo���;���-�Q��0�W��P�b$�$C�m������֢�a�æ���̹0EP�b�aǓ-�th�ݧV�����]C���ڴ�e%�H�@�/�>I�J��D�T
a��BN7Ob-�
"��9w�r�U���	��[������acGxrd���1��tL(+�G(c<pl���c��S�{�� �t}�=ga�~1��pz�|��4���a@\oʇ
1�c�Z=�;�=}9%��� �
��o�O�~/L�H�-�){O`�$z��E����Ia�iȰ˨;���닁�Lf�$��SɃ���Xz��ՙ�~��q�����)6L�x�.tWBmλ�P��Li�~�	Ec�ސ��y�R�$�ベyA]�ˉ|IP�jq��d���w�̜M�C�	��rg�+Njs���F�2[&�N�?��j7?�w�L[v��:��f �N2\;�t:�Dc�L�1pX���<����������k��L8�Y	h��� M1�_��vW��(��NaG�Y�`����8+.��Y��3�M�4�c�rY����W����*�@ˮ`��~3����T9_�G�D����^N�R?@�"Ue���Ҽ��1�!����{TЭ�Q�ҡ���7�yޙ�,���h���6�>���bK�wy�H�~nV�n��0%����iKFʍ�ONm���s�nj_g1E�᭳b��\���}b4O���T85;��h��*�)0�y���\.���kj��~�|%��Q�Pk�x)熼n��E��z����2��佶E��v\�N}���V���*a�������U��>����8�7��4=�5�@4�;~�Hj�!K!BZ�c�͢����	�N$�_@|89�jyG�ϩ�n|?/��b�s����oo�����^V�	�HH9/M��<�R2-�ĕJJiQ��V�j�5��t-�����<����f;chgn��(�krj�l�B	A�0��0�ˎOx�x�fvO�KkK|��b2���D|��VE^��	��xS�O���D
ի�i��3Ҥ|��!n�Eq�
�4h��4C�H�1��}j����7�M��4&�7��,c�M�77.�I$��vq���	�4�z榺��,m�9�ln�+�	���x���k�=��!>D�J�'siJ��ӫc��6Ά<n�kВƘ9_��N��dOw��i�l,�X
�%�O�;ɨ����KR���9B�Sr�z���x:�3d���.r�i]��~��_���-��:�IO���0L�f�I�������V��C��f���l�Jگa�I�"�߲��M:9Ja|&�����3(EO���a7uo�&yV3W�벣#�;U��<����]���� W���SeH|������;��V���$�<J�L4f��R�V��H�e�m.��W��9�ʈ�Hx�r���-��aF(��8��{,T�3�p����;�p��~�o�#S�r���O��V�POV�q�A�����Ʌ��!4p�k/���y��޵mVv�V_g��,�A��,�y%����0.�nݤ%ňV���;a\ah�S�׿*��XQ\^}���T(���7˴�>�}n8�� ���Q~�Պ�VBA}����
�YL����}9F
BljKOP�~N�|�W;�ؒ��
�po�y�Cc���AdьI����W
w\X������3�1�������d�&�	V���<��$�3���~5�e1�MKv;i�� �,l��1�s\�vf�Q�����3
��&�@fq�@���M]���u�|�Sg�&��&1�'=W�����	VؕrR	'S���N��u	�Y��tP?�F��@��rBb5דڄj �#!{̀l��|Y�3 �Įc���HP��ޙP�ZF�x�*��q��^�l�=c��&n㇭�Y�wx��m�}k�� �}�s�V�t��&jI ��8OpW�NƀbHf!��7sR[Y��"}�~�焽!QM�K���À�i��̑d��qL8�����MDC��eOI��G�'�`
���^���e?�J��k��lZ4�1~U��L'͊,uAyv�(��9�^��� ��42���{���R=��T��u��mL�F7U�t?�Ru��ZwVܘ�-��)s��.�,�̿&���9��Y�ۣb�`"B-ʾJ�ul�n!��'���?��@�z�۞ٲ#�BI��#T&+��g�z+� ��N��-_�n.��B	�h�4�zT%֑�5oB�/|f�_>�ֶ5�����y�H �i��3*+P����PA�b.D��0��l��W�TZi�iЮ"�;�K\���[C4�D��P�������|z7�'!��P��T��Ce[��%/����T�r���^
�WPou\AZ�F�hA�����db
&���D��
n�1 ���Lx�>���d-c�*�[�U/��%���O$�Q�I�p��������ũ��Y���4��%�u��^Ȭ>���ѧp���b��]�"~榫}�Y�ɝ^�b�Cs�p7�p��� �8��Y2h	���a0o�����;�6�*�I�[�\Ըj����J`L�Ϭ, m���i����J0.�W��V�A_��������?w�x5$����
�vl�!$�N��_9s�dh79��J&�Lye9&����JLl����vہݼ3Ɠm'�9� f~�{������7a��Ɨ����˧�ddg�e�� `���F�8���=%�eL��$?1+�^g.�_ C�E���k�XVz���[�����X��o�� ������H�2z�l��miǌ��z+�BH�}�&��ǒC���$��XP9��w9bJ�pԯ��y���f���E+�.ϙ.��0
���{��k�s��Fw{`G0|R�A.��$�y@�t_��|��a�)��W{I.� |T��W
Ҍ�)�U䆄�Q���A�Q�!�B"y�s��v��5[oU9���E'���&��/�h�Ǎr�ֽ�G����ڲ����,<�\�]WS�/\5)4�=H�� �=P	1�(�4�@<�����:��i���	�Ӗz�)���j	�=�N�Sl۱�ZS>���.��k��NE�{$LW���j�[����������,�h*#)5Ӯ��]���7������..�L���B��Jڌ�+����݂���ˌ����I�Pu_F|VJ"|Q�n]y\�1k�:G����Q������KX���(�_Dqށ�2����If�B6�%_X����<�_8,uq]*F��CA[D�ϗEK��LO��Q6��]�6M/��iXv�{�#��K�<��H1����B\�l%?2�f�zX�.}zi�%��IIx������F�B%2���y]}�3���iK�ˎ�4�p��G���N����c��y�-�- B;�>��"�Q�lM���p��b�Y�����j�,�a�}Y�f!�'�0C$�b ���ԫ@�+*���|�ʹ�.�fńwKuz`xz�5�/�i�]?va��F��B8�� ����ލ�Έ5��]1�6rURo�ɱ��{�����Z���0�R�#_�N_^|��gC�t�W	��/?�,{K��F�gt[�/���+gX�lh�ʹ�n��n�A����t-�K�k���D����7/��2Aؿ�����:��egf.*XxΨЮ��B����o�9��(�n�<R:���Ջ�m�,�,��}�Y�6{K (�15Mc�Ӻ(�����5cG����!?���ƐR����OPa�Q�����7�V��&�3	�r�j����~��������!U.`_͜���j>��$���+n��oM�2�6����q������ul{����ꃿ[��0w6����V�H�Mig���|��1�<�0�Dw� G ����]U�ݸ ��KC���"R��be����˧^�]���"	_R/�fd.g7�������;�O���g�;B�D�\e
�7�Ç<E�x�HKRȿ����X:D�ĥ��V�p<��Оc����l{0Vx:8�ޯb!�1눪7�X5�����U���2QϞc����o�x�᪥p"dS=�������4zK����JR���H���:�R[��3�Av���i������f�	ɰ�w� N|�R+}%���d�Cގ,�ِ���/�D�;��ç�ef0��y��:�^F�c�=Q�[�>��=p�s���gr1#y�ִ��HK���:�SºeT�o%����V���7�N`[=��E�Sr��pR��#ZdBu-�Cyn��`Y���+��.TQ��O�^G"��s-E
��*��F�m)�i}R�l����&����pp\k�R`9�@5>d��jY��С}��ݢ�uP��W����^�Znjg�Ϛ���\:&�:~�ͺ2����k,��zn�f�Sg�퀭�f�Ó��r26i����
�@/�Es&��:ɝ��-֤M��Xy�t�ZnV����"�2Q���2��Z��g�fB�oʛt��q"r(J����4F1@�r.�|#���$ogw�tX�s��� �?jI�U�
Hn�|b�4!�������_�֕}�73�I����^}mH�v*N#���$�%֩����:;��vN0�|��"yk#��]�un��4�X�D�u>�X00��fU�^<�W_�!�Њ��kI����O����F��ΆT�כX�ۮ�=ҵ��vh��{=;e�b�G�'��� �f�>�5)v�h�h	�	�r"a��� ���vVj�U���>1�Ɵ;d���bC����|[qs���<��>-by#��P8�$o�a3��u9�5�0����s��{��e*Y!�Y�T�����ϋ*��ˉ<����s�	@�e]�#*!�7i����:���Luy Ч|�0�殤G����v�J��~-�r,�.���8�:�=�8�ď��v� �[�q=��ұ�Q�a��jwq�m�Œ<H�H�v�.4��D�޺E=�/t�,W8b'c	�y��*�Q�u짝/��b&��oN`�n�>"w5@�\3O*a��5|<��ۘaa��c��u�w0�}|B�*���E�vQ���J��� )�����.tx�H ]?G�	QH�e�U�#d���N�+^�,7����Ã�$�W����y8y��ق��+�/��ߋ�}1.><��y��Fb�8�*]��e�@/�)��!� �5s�&��|��`q���Û������`����?��%~�@i�C�e�^C��b�XG�1�X�p]G��FY�z ��(6�IX�~ׇ�]-WFc}�"2����Gx׋���
{p���[����F��+���X�%w�����#�A�􂓘��.���*��X�m����ɠ�Fŵ�2ʜΑv
�������m��2U�?��>ۊKG~��)���{��_���&ͫM��T>16u�Gs��Lߕ��$x��Q!�:�zZ�T� ����)�B#śY�O�(za!C6�f�[;�R�lr���@���B�j����4�G�"���]8@٩�	���i��ЕM�H�NՄ3��^�O-";��Ka��� bw��CF~,�'��%�ק4��/FQ�_2P08�^bW�e�FAt{��Ptk��$��'��<�3����@NF��Q6�Je]L�'�a"lNʍ�-zz���w@-�hL��|6�[r,R�#�cڙ�d	2QO��4��(0��G�xbp?��W�c+�|��S�3t0�=zwN~��%pM�	���7-��a36��"���=�>��/���E��ؘ�<�ʢJ�/��
�@�0{¾�$M��E��v�L<��i�������ಿ�$��~ɶ-V��
��<�~�����~��˅6��7���B�����5O�?O>~R�3c�ա�����Śnضyt�#���P��W?1܈-�������ج+<�J��j��9�32�zW�ĥRe�j�l�wS(�v(�r� ��U2^�8�'rNDv���`��|���g��j�޾Ѿ�`�r�Y���y;��!�1���}Y���]1�43G�%�YU�qRU+�Ū�{�3]Z4�ۤ���k˅%����h`d�@���HG�3~���G􍅚�DQ���{PN9Oh@|��e�K�O!�1�#��;]{o���A�
�=��Lf�h�Ϛ�5���CZ��hK����_0}�D�8�X*}9қ�x�q��`����9�m���/M��~�e��N��N�)�6�x�7�� �pl�Τ�F���w�N���3� `�a�ju���H�I��*�Oͮ FԀ�e�a���u�{ֶ+X���Ԥ�3�7:	����O�D�'6�u=r>:�G2nF�U�OE8h�ѝw%ϖg�i1PQ��*�\+��   �  R  �  �  O*  �5  ?A  �L  X  zc  �n  �y  ��  ̊  D�  ̜  �  Z�  ��  ��  ;�  ��  ,�  ��  g�  ��   �  f�  ��  ��  (�  j 	 � 2 � "' d. �5 �= E L FR �X pZ  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�xR�)�S�y���u䐷Y�m��ìS�4C�I
Nԕ�d��Ų��G ܜ{����p�qb쐪a��1r�a���ēc}��[�.��m1����cC
QV\��"O\��G(=t�,ya���:�0e�' �p��Ü-�Q�� �t5��&!D�<�F�8NԲ4�g�Q/.�|ZVK �v���R�P�V�Q3m�$����Se��ȓ*�.a)�%�54�����͌i?��S�? ��: &&<�tHp'�H�G���"OXui�JU5m���p�G_[�xHS"O�(p!�#Se��N���(0�"OP�HE쁨3�r�htn�@�>-sE"O�YP[�8c�i0OY_���)q"O�LRAH�%/$&�J��Lh�r]�"Ox��S���C�l�XD)PUݤI�"O֌��T��X��1�CC��0Q�"O�|����)	 ���@OH�-"��!"O��;V,�=g���JA�B�3����"Oh��3Y�,*�Qxc�-Z�t��"O4`� �3+��EA��}�I��"Ox0��V�f� �
��L�P���C"O�h2��Ӂn��<�#%	l��a�"O1Y�#�3��� D��|2�Ȑ�O��=E�$�(�̥����%VHjD� �y�-.Zxђ�A����7��ItX�8s��A�1�"��7��r�A<D�ܩ7*��!�y� �|�Xh
.&D�D�Z�D0F�VH��`�8D�X��i�"~�䠅l\,@�
(��`6D����k)Tp"`��h܋^�@m�Te5D�����rVd	�bM*b�1�s9D��hSB�x9��c��?3��`3֊8D�	Wo1Y�L����G2 ��D� 5D��2Q�1Q�#��'kVq Ã1D��Q6�^��p2dD�#1c�1D���� A�ds�k�$5� �!�<��2����-$q��Kc�X:�Re�ȓ%y�|�t��:x� �;tP`�ȓ~���ƨͳ>�p��K.IXZ��'�ў"|�A�&�<��3\BBש�D�<��'W-�*��5Nۨ%�J�q`����=i1�� q�jT	����
�t�1�B|�<�&H�1Z��`#'L�
6X�jG�@�<q���X{�pW�H!%�>q���~�<)���kv]�Tg  ,���-J|�<�7�ׅsPXӷ`��H ���an�<a�͉�%��0s�Dv�$��%�L�<�ኍ��rU�-��pu���d�{�<�֥͹�
�G��.�j��f�Jw�<Q�-�#h-������E�$���Oh�<90�Q,9�(���# �ZL@��Y�<��MV�0�\�8�HԪ��u��T�<�4ܱoF�cR�Ӳ����G�E�<aCP'o`�ĩ�-�����n�%�y"EJ%㰱HB����LU�ͬ�yb+��"�e�r@H����"�GU�y��l�"����	�`�#���yB���H�+�fN�M�$xbV��yR-P7D+�l寅�bh.ABG�	�y"b^7!3�����#�tP�a'�(�yO�)��Lc��)o�(pqρ��y���.�`qD� %�m@a����y"b[�7"���k�4D�e������y��Hb"Vɑ�c[,3�>(#�(	��y��ki𚂤#f��6���yb��<��9u�^pp�� &�X��y��Z�F�p�I� �f����.�yb+ܥ%.�<�W�MY���
5A��y%Ϟ#y0��Y�KT@��"=�yR!�,M��a��4�	�B�y���M�\0 ��h�����&
�y��ˇh�@��HW�_�"�s���y
� ��giѩU/̼��/Qf���"O���2o�&K��9C���Ĺs"O*��熗.T�Qk6��*��!"0"O�AP��L�:������`�z�K�"O&9�UH�,$��kCK�s�`��'���'���'m��'�b�'��'������G����X��)2U�'���'�'��'��'�"�'���
T�B!٪a��F՝LS�ʅ�'ZB�'Rb�'O��'���'YB�'TXm ���/�b!`�ޯs�>8r�' r�'Z��'�R�'�r�'���'.2I�d.�9���Zt���O��E�V�'�"�',��'���'��'���'�l,�C�#PL��_%~�
��'���'�"�'���'r�'�b�'�x��%��K�TP����&��=k��'}B�'��'���'���'�2�'s��ʦgҹy&�q��M-�H<j@�'e��'�R�'��'0��'�R�'b��7M�pXf��ԣ]�{���.�?���?���?ͧ�?q���?����?�#��d�]�3�G���P�db���?����?A���?����?1���?����?�q�Z����c�C8�9C]��?Y���?���?���?!��?i���?)tI�"�U;���ju|i
�$�?y��?y��?���?���?Y��?	@�\���;Ge�g6$sS�(�?9��?����?���?��87���'R���3�r�RtÓ�LcJ����
ʓ�?!)O1��I��M�ČFm���K0M�;>r�%	&4���'�6�6�i>�	ß����&�$i����;b�d�៼��� �(	oZI~26�\���E�)�2�H����<%���0�aL:D�1O��D�<a���P�qO晀��f���ʔ��/0�j�o�o1�b���g��yHZ�`���e�+C��-[�j/F���'�D�>�|�'�!�MÜ'	���WkK�e�rPb���i�9��'��G�$���i>!��1T$Fd��%9���2�Dſ'y��	vyb�|��qӎ(j��Y�Y d��[n���CB��j��D��O����O��IG}B�(Kf  �t���}g^h�����d�O�H�1�B�vO1��L��vOj�� =I���K��W�0�ߕb�ʓ���O?�I��b�[Ƥ�;��E@b"O	��扲�M���t~�GfӖ�擴n$� $.MxΥ��%��J+��ݟ��	��@�,^���'��ɒ�?�� ��	V�&8��	��k�"��ъ�A�'��i>����@�I柘��%)ݴ�p�I�s�����D"����'TV7�C�&�ʓ�?��4�� \��Uj�0_���I�	ؒ4����FC~�*'�b>�#�Y�e���!7�=��a���rtd}9h�̟��Q��B�GVֺ[V�x��<IF�oc�Y��^1�e�ǟ�?����?���?ͧ���ӦQ��O�d9T�]�x>�#!*I8y�l2�֟l��4��'�2�v��tӺ�DJ�H2����
�&z���D�e����d}�p�ɘs��DHr�_�9�dp�[w2R�O����q�˶[^�X ��/ ��sօ�h�	ß|���\����4�J��L�'��2B��_a8��=�?i��?IԲi$�q��P�t�ݴ���䔻%��;q�� Nہ6�r]�Нx�'��O8(���iQ��n(�y��T"f,چ��X���&�ܓ���`�Ry�O��'Y��+LQ� ����,��:w
�*b�"�'��%�M۠�[&�?9���?1-�*!�@�!np���a��B�s񚟌b�O����O&�O�SI�jŁ�9{l,i�"L�>6i�ĩV��,\oچ��4�����'J�'i�5�a���>]�e�<�u��'1��'k2���ON�	��M���j�,aa��"�x���Z��.Ox�nZi����	͟D���R�^�Z�(dO&���VI䟸��>54l�[~Zw�Z� #ԟL˓-X4$�6`؊W7��j��^���̓���O����O<�$�O�d�|Jt��t���􈓠&�:S�\��G��s���'&����'�.6=�Ypf�S�'�8B�	C#3���)��O��d�c�)�ӍQ�]oZ�<ْ��<Y�n}�A	�!'�(�R���<�խݷ�N�d�����4�.���b$*iJ$�%�`i�@�ɵ��$�O����O��t֛���O���'��NϚ1�f��i�:D�-�f"�l��Oz!�'���'��'�f2�\tx�8$��|v�a��O8��sȖB݀ؓ��7�)��?����OHI��Oʯ@[X��ň�>T�(����O���O>��O.�}�F3��r
�_>N�Hӡ���	�7�vZ�m��'t6�,�i��0���cw � t�n�hw�t�`��̟�I;x��	lp~Zw�n�x�O��!2&�gв����x�8Ђ�A�O�	Zy��' ��' ���yG��&~��i�u��:$�P�p��=x�剭�M���?����?iL~���� xh��]��)[�Je�xaC�Y�l��ҟ�N<�|�%"�E5n�i�,��4�PI1C�A�`~��U�Z~R� �&����5��'�剪U�q��]��=s�J+����I��	�(�i>��'�D7M�o�R��-P��*���}�� �aV;O�8�����?a�Z����ğP��4}��`
�AL6��ez����k6\J�	�/�Mk�O�ur���j������ �)�)�.���ʶW/w@,�=O����O&�D�O����O��?�jB-P*JDy�"?����B%���ԟ��4fn`�x-O�AmZ_�	&b4H3D�Tb���ٴ��7�hJ<���?ͧs���[ش���PP�3�\5<�P�t��(�\� ���?�C)5���<�'�?I��?�U�I�|)
��˥���wmԷ�?�������%�ת ���Ɵ�OE`�
3 M�e�t�	񪕳=`���O���'nb7�D̟�%��|�@J#$I���� �BJ�~t��
�&51�!_���4�� 0��y%0�O��+R�QX0�'�)J��#D�O�d�O��d�O1���$��6�kP,uc�n���
�던��Y�FU� 8޴��'���]���ז
�%���C(d@ͩq�х�z�$}�Ph( k�B��fP��a�����.O����lL�Yȝ��m^�7.Lx��?O���?����?����?Q����	D:2Ց�Oڦ=�r���ⅶq�"�nZ�pb�Y�'&���$�'��7=�v�:'�W��������+D)ij�O~�:���\�- 6�v�ЫZVYRGj2�ـ��p���%B� �0�'��'��I埌�I8C���%��"j���@�/Ԃ%;��I�����ʟ��'��7�Me�\���O��D�SHq�!#X����Ǚ�eՌ�T��OunZ8�?�O<ɕ&���4f%Jw^0y �w~2L
J�\d��O,��d�B Ig�� 4gŇmB�h֮�%B�'k�'�r���P�"/
�<2�|I�.!*zB��R(���8�ٴ;�R���?y�i��O�n�2s4P Zi��G��p�)�hZ�A�����McE��M�O���i̦�bG��*����e
�#���@�b�OK.�O���?���?��?1�6h�9�LU)fIz3��Ć/�D*O�l��#C4p�IП��	q��П8�����o�B��R=+�b��3c\%��d�O�6-\�)��� ����S��x	B� @�@"C5���Q�љ8a�ɁD�jPIS�'~'�X�'N�
�R�7NHs�`NBȼ0��'v��'7r���U��ٴK]�)�U���i�DJ�N�6`��%Ɉ_|��@�F�V�$�Sy��'}��v�4Ƃ�	T�J�LV�c�ia�KP:�7(?!�Œ/GŊ��#���������B��B�Q�����u�(�	�D��֟l��͟$�Z��� c̨{�IE���,�T�F/�?9���?)��iL�R�Њ�4��&�� �\r,��T&O���06M	�ē\��6�x���Z6-6?yrJ").F1Hu��/I5䘚����d�4�"�O���L>1*O��O���Ojt�g�Q-)-�0�4�'*,V̺��Of�D�<��ivNd��'e��'!��������;IG�(I0��#E(�:���낄�MK!�xʟ�����p��c���-VW�KE�^><k�aH���a��i>����'�t�'��H��K���!�c�qYD`�� G˟L�	ܟ��	ݟb>u�'J7����B@r� ש�h=q&.D�w#x�ۣ��<!a�i$�O~=�'��7�f]�x��	��ZBm�0e�����+�T���'f��𤆎�?)�6T��"c��1�ݰB��>����&ku�@�'���'��'
�'��ӾY��m�S����2�L�3�F)�ߴY�*d����?�����<q��yׂ���L�Bډ?�e�s�YB��'y�O1���S�Cl� �	�d���D
�w�$�Yp�@PJ���8h��'�$�0�����'>\�{�擑��Y�g
17��Ñ�'LB�'^"Q����4>�.��*O*��� x7�そ4^X �&�C�[,���O����OH$&�cǎ_(Jɤ�@�K�=��1%*?ɁB��+����a�Q�' ���D�?� M^'$B��A#>�����؇�?����?)��?9��	�O$�b���x��0Z�!�_��4����O:o1�6T��ޟ$�ݴ���y.�,.����r�A��9�&i���y��'���'C�ՙd�iH�i�Q�f(Z�?����6��t��>�~�s&I*U�'��	՟��	��Iҟt��%/^ƕ�Ed؍^`�ă	9���'�6��7&���O��&���O0p!���j���P�NƶV��EjDcPU}��'�"�|��$�Նc�)��)�l�LX��Q$UDvL�+�#��ɂG�TU�A�'��x&�@�'��\*�Y�jf�(ib읐LMF�R�'c��'�b����W���43��@��bd�ػ��<i`�2�"^$b��A1��"s�V�ě^}b�'��w.y�u�Y�o~Fċ�/�M:�����#A.��<O��D�6(B*X��O6�I�?y�]'�H�@-�&B
��B�VI�^�����I⟌�I�D�	E�'@�F���5� ��,�"��"��?��C�������T�'�x6m0��'�h�c�M�>Z��6��
`x&�4�۴*a��i�$��4��D�'�n�U��@�$=���9���'�W�?QTn;���<���?Q��?�$F�<*�qa/��AKY�WK���ٟ0�'��7m���O^���|��΄</����؅ ݾ�J� �X~���>Iװi��6-�K�)����7@�ŀ3�F!£�_�.yK6`��tV����- ���`q�|�I��Y!���#@;|�}P�F�=*���'r�'@���R��2�41h4��.U�;��;Dd�g0�m��
��?��M�F�dQy�i������++T��v��G�ysf�m�d�n�8<��mm�f~�=+@����}�� ��w��$q��9���U ���9O�ʓ�?i��?q���?���I[�p3"L�Յ�8�`=q��8Z��EoZ�tи��Iퟨ��w�s��S����d;-�&� �*T�&UhV�Q�m@���wӾ$�b>YZথ�kQ���,�� ������%��ϓ.˶x����O�]�I>�(O��O !(S�	�,X`��bZh�bd�O����O����<Ѳ�i�d���\�����?�pd���]�z��%Q������?�'Q��ڴL��d!�Q^H�a���R�9�H[��Ix��]���>Pc>���'
P��	�W_N5��f��tcJ�ⵌ7P�4��I���	�h�	^�Oa"E�4����Gk̕���C�_�^�b�hh�ᏺ<I6�i��O�nh���'��t�m)#��=^(�D�񦅘ݴAZ�v$E���֛� ��C�z���-խ~�Xi'cO�W;���m�?7�<�&�����4�'`��'�"�'�ҽ�"�b}�"�E�~>LU0�]���41b�����?	�����<��.$=���![�n�+0lF�<��Iߟ��I���|b���GƑ�w�~8�&���3���&\;l������V~�oͮv�B��-��'��ɚ9�:u���H��0,��Fe�4���韔�Iӟ��i>u�'|�6-�{���d��S�
���QAb�ሕB}��Bݦ�?a�W����ɟ�	�G~���D3g�C�$;g�\+�$����'��$��CQ*L~��;/f�	���ӽ+8�J6H�� I͓�?Q���?���?Q����Oq9YR�QT/٠@�B�`թ �'�2�'I`7�J���Oh5nZQ�/x�Vp#�(ڽAB
Hc'(M�F؊O<�ײi�67=����֫t�"�^�歐vȅ�
�	��8���M0�J��>g��O���|Z��?)����Py��6�2əFaԕ6=&�:��?�*O��m�9=1� ��֟`��[�4"��'i�G],2�h3�Ţ����x}2�'��d0�?U׮����ɺG�O,��áʥq����V�{~Ҕ�����Ο�IÒ|��A$%�\�u͜%:@
I:A@�y"�'���'����U�� ڴg2Y�@R�%FTsEƱ2/ݕ�?��k�V��X}2�'B20��Ѻ1�y�,�#.S�#$�'��f������]�1�
����$̕	Tpڷ��g�JA
4�Cj�ĥ<!��?����?)���?�(� ��C�,�@BUi �B�%Ҧ�CW�EZy��'��O��q��N�
���7�фw�Mk��ѐ3c���l�H$�b>�s�F����͓bap�Q�JV,�@��B�9l����$���+�O@��L>�*O ��O4�1@,�]U�u��+x�*.�O����Ob�d�<)s�i�>A�W�'��'�&�� �B��\�
�%ۤ�u����a}�b�.��	v�-h��ͩs�D�}v���A�o��=�Z�@7k�<,���O~
+�O�̹�j�̸��L>l���W�UC�����?y��?���h��NB�E���B�=il�Y#�Do�>�D�̦����M�����'�M[J>��SdG��1�qo�I��`�'���<A��?��H�p�4����`3k����ArLJ�)p���A�Oƪ�Q�Jü�����O��$�Oh���OR�$��k��u�J�2ZV-�������ʓ2���,��,R�'�b��t�']�P��EMB6V ѣOÚtj6�Rf��>���?��x��D�ҹ
�� �ŪW����'g��"F�P)���b��C�U�O˓p� ���H�8d�Z$�X.0�dYK��?i���?)��|�-O$ymZ�d֮��I�&d�6a��I醍���5ڤ�I4�M��d�>��?	ƴi���k�nU�+)���D�/�N���`��6���;��h��$����j�3���'Z�D�aj>G��k1:O����O\��O ��<�|�`�(^T"p��# �*]*��:�?���?ѣ�im�q[�O��a��O��WL��_�Ձҥ�{\5y�k^@�Iɟ8�i>Y����%�'� �*ֆ��;�(�R�IP4[#�8�f*izlU�I,E��'y�i>��Iӟ���*MR�LXs��=�f���#��Jp=�	��'��6m�>~���O��d�|R�ƝJLl�Th2��f�~~B��>���?�L>�O7<UХ	�X�hE�BBΒYCd��V��]9�D����6%l�i>�8b�'є�$�@K�WRhش.I4Y�8��b����	������b>9�'�7M��J�h�W"��*�ݒ��ݫ1l<;�$�<��i��O���'��o�T9�un�"��9�򡔺h;��'xrI0C�iF�i�Q�5/T�?�rU����⎟[�PY#A$�dm^a:�#f���'�2�'b�'�b�'��S�aTʀ�T��$�.��q���㦡z���ӟ��	���'?�����M�;���I�h�k��ж
�
+�M`���?�N>�|�r���M;�'�z-E�ٮd�Tј��^�YĴ�+�'���K&�̟�՘|_�0�	���Ka "%�zHf�_�H4Y�P����8��៼��Py��`Ӯ���o�O��D�O�YY@'��&���M �f����>�	���$�Of� �D�Bz|�A��U ��� ��O���#�@����Ƞ#<�H'?����'6�l�	,4�<�0�	9�  ��A� ����	͟��	ğ��	j�O�b.�7F������G�T<�!�$\���gӨ���O ��Φ��?ͻ]�씊Ū޴3�`�ɋ )��Γh��v �O47�ό1��7-6?���� ,����Oi�? �h"%��3X����f�da3&�D�<����?���?����?��-K�*�p�0gI�T�T���L"������0�nԟ���ן�'?���n
��{�nCpC��F��9����Oj�oZ��?QI<�|r�"!5��Q���_5���[fb�&1���Rp����$��4�� ��w@�O���Z&�ȳDt90SA�J��4����O��O����O��<	B�i��eq%�'����%n�:�@��H/�ਚ�'r�7�#�I���D�O��I��m�sA�h8��KN�Vfb�FQ��V����57����'������,X��(	$gĜ�@ެY�D�O`��O����O��d1�S i�؀h�˩m�Tpq$[�}j(��ɟ��I	�MK�E�|"�0�F�|bh��� A!Th(�ؼ��
|��O��$n�����s�i,�	�q�jt�ǍD �I1��ê 4�#r
[~�rN�F��Ey��'��'bjҙ*����Ó�`}�OǾS���'��	0�M[�j ��?���?�/��<�'[tt�P U?R�Z�I����,O���y�B�%��'t�:@	�3bA�ͫ���<7��[G�b���;$�y~�O�\����s��'�x�0s!�'P���/Ef�:(*�'	��'�����O��>�M�BAX�IxLL�uo��(K���-D.L1���?A��i"�Of��'h� ��\�)���J�@G�ы�%�:S�2�|ӮD�4md�J�� �RAE���O$�HvlC�P�T-���V�L��T��'��	������ �I�0�It��MD�U�ڰ�.����!�oۗz����͐v��Iҟ<'?5�ɷ�M�;�֤1Č�Be��
$@ȔQ �����?9L>�|z��G�M�'�$�%�6?�l���M�K����'@� �s�V������|B^���I���K�Y��@r fO�i���oI���	�(��Wyb��Јs�ǩ<�!,�)Rl�y��A4,�1��8��O�>)��?QL>q��Y�PD�j᠐�8��Ё��E~���7�`i�c͕�F�O�du�	�ڢ|��Ա�
 �h8)s��j���'�B�'���� ����y���1<� 9Kd���l!�4ce�".O&�o�W�Ӽ�jH8>:��0��$I�|1�-��<��i8�6-Ҧ��+O��E�'B�<�"��?1)�E��h���'e:�+�`�.Z�'a�i>��	��$��˟��IE�H�g`ȕ]�
Y���%3k���'f�7m�:u�&˓�?�J~���4�xǣ��a6�ljTʊ�2�bU�7[���ٴV�r�x��$,�Ku��U��5&8��B��5���{�aS��� V֔�#�'*L'���'����� ?�4<@���3���P�'*r�'�����DS� �ܴ=y����g�B8{�C�m��Y������a��1����N}��}Ӣ��I��k'�./� c5h �`R�3��J.t�Eo�X~��H�+����S�;��O�g$�X����5���Q��y�4��y��'���'���'����Vz�b�����0V�,i�ŧZ�k�d��OX�����eaVI�my�cy�N�OB�����!D0�<�vm$gc>	# $�x�ɒ�M�5��2����M�OF�K�^�<�
!�ĬrW�\x +��}9��p��ؒO�˓�?I���?!��Jr��L)K
��#�W�o���ȶK�O��ģ<���i~�1��'b�'��S�A�ְ#祐�i�����K�|������MK'�'剧�)ӭƠd�E'O2j�"P�
�a�6ݪa�ځ9SRq�d��<�'m��ē	��#�0̀���2 �Dm�0�؂)'�����?����?�S�'������z���+5�\(���j�[G�ơ����ҟ��޴��'k�듃?�&���r,�8i���G�4�?1��+���Aڴ����(8�M�?Ֆ'@��i#�Uẽ[�F\Zh��'��	�,��ܟ�������IZ��N��Q` m ab��� �d�N��6�@�5!D�d�O���=�	�O�ilz�=��E�N(� �^�C�������IB�)��5,2Po��<YbK��DB s���G��i����<�A�	0"�	I�IPyR�'r��=\�@d�$�������'t��'��I��M�G�C��?���?�0�?�tej�KLn���ň��'Ar��?i������ijuO	�O�@�� �{��'�$�����Wi�v�-�I�~B�'�X�Jg��P<�`C� ^}�\���'`�'��'��>��I|���k�2�p@KG��r�I�I��M�p�\�?��a�6�4��i�
�hnūcR=�e��>O �n�=�?��4]�
l�ش��$=�i����n�`#�di�h��(�-'}T��?�D�<����?���?����?�v`K�4�25�p��6�y�cѳ����Ʀa:Q��ʟ�	ٟp$?�	� �^��b���l�q�_�R<A�Op�d�OƒO1���dG;6V� lJ���(�K����3#�<���/
=>�������ߋ9�
�ET'7��L����u�����O,���O�4�J˓/��ãM��"��zԚCT���i�T�8�yҀf�p�X�Or���OJ�o$��+ �N�o]3��8/m� ��b�ᦅ�'���C���?��}���%I��𩙀��y�ea.�͓�?����?1���?	����On�a׏2��k`%D76>�HڢQ���	��MS���|���T��v�|2��}�*�X�&'������"COx|oz����Xdc�,� �2�� �m�S)B�v�N8�6������&�?9��-���<y��?y���?�7��`5���T���>I6��A�P��?����$Ʀ��gD�wyb�'3�S!	Dp�p#�S�P"���y�L�`�ɖ�M+6�'���)1p����D��v�17a�-h&ӆțE��`K!�<�'h �d���)ؖ�q�� � EVf�>k��mq���?����?��S�'��d妽q"�I>/�4CףÐK��AP��f���	�L��4��'H.�)͛Flɥr��h�@��]f�a��*�"����m�@s'Hb�R�^nx���$�0/O�+`�_�G���z�0"�a 3O�˓�?���?��?����I�3X�(��6{�V�`�o���	n�9��ٗ'"�	���ݠ5�,g�T�Aʲ �$�Ɉjb�R۴U⛖L0��Iau��ڴ�yr�;D�@�5T+�N��Vč��y]�D���,kD�'��i>%�	'_Z����/�m�<踃-޿}���������	ɟD�'�>6�8jN�D�O~���x��[�)@�3��w-L3G:�裪O*�$�O��'���s�Γy��e�$ŔD���P�'?�6�B�>��k`AYJ̧5����X
�?Q��$�a
sgL�:���	M�?����?����?!��	�O�(��i�6<�z�3Ć'�^�� �O"YnZ�o�ڜ�'φ6M2�iީ��	^�3(襻c�*�a!��|�t�IҟЩ�4uJ&=��4���N�|���i�'K��q� �	f�ص����X��k>���<ͧ�?����?9���?y����F@q�W�U�ɱ�)�����m�AhN��|�I���'?u��-lZ�<�%�&k���3�
N�s���.O���`���$���,�c�P�
� !�4FOH⮠�S��o��� ��PAC�J%�RT`��Ty"lJ&`�~A#$ڪ~�F%q����r�'��'s�O��I��MU���?Y��U��`��
�2(|"��c\��?�$�iR�O
,�'���'�6-D�J�(+'D�gRM���� H������o���.���E���>���
�N�Qj��K��x�i]+���	��H�	���	ܟ`�	[�'�)�+,;�`AqӸI$�(O������J$�`>�����M�H>��Aͬ`�m1��	'<��kr�I����?i��|����M��O��,V�:A �V*(=�nN6~��;Et$���'��'���'Q0<²n˦q���c�L^�dӀ��'��Z��cܴ,��e9.O���|ʢ��)�^�C6oDZ͒ �<����DԦ�X������|���6���yf 	�M!l#W��(@�
8�h
J�t��5����?��?�q�<��L_�U�����4(Ĳd�]�l���Ov���O���I�<1$�iq��D�$5�@㖑L2P�D�&@ ��'�|7#�4�p��'!bIZ�?6����H�Q`y���m�R�'�	 �i��i�A	S��o*-O*q1�͠9��D���[�wl�t�;O���?���?	��?�����	�R���s��=�>���B)5Ǣmm�k��1�I�l��x�s�0b����!�ֈr����0�`�za�E��id�O�OS�����iq�$5-�LѢ�V�֩�Ui<� �D}��\�l�OB��|��E��1#�Nؽ�yk&+E��n���?I���?�(OJ�nZ�3��e�	ƟD�ɃE��l�� N!hB% 3��$�?��V���	؟($��Q�'@�/�b`!�Şp<�#b�)?�BHS�x�D�͖��'Q�����?�`-.bY�Б/���D�)����?���?y���?��	�O2|�QF��DHq+DP�<
���O�l��uEl��'�,6- �i���)O)GB�Q��24��lf��	͟�(�4\�Hh1ڴ���D7�P�'HyD4IG���8q��e.a`1��g$��<ͧ�?q���?���?	�j�8xL��k����dy������ЦmP�����I���&?�߶���HҦFx�e�ˁ#�$��O����O
�O1�������oT����H��m�c��z� �G�<��i�`a"��������d�$_zL���Ȗm��[@���r�T�$�O��d�O��4���U���g�2Og���J������(2���aX�G���q�d㟐2�O����O��d�{%��ZW��d���p�Q1Sv�xa{�"�FŸL�����xK~��R�T���+�Z ��(T3����?���?���?����Oa�H�v@&Ҡa�͆J4�|Q�'��'�B6V�x"�ʓ$Y���|rĞ�ek�=Q@	"������E�';���
�z������e��#���'

8�r�D�7��1X�k��Xy2�|�[��	ğ����pAs"�=S|����1hc�,C�̄ޟ�	Sy��h�J���O��$�O�˧`h���X.f���F쐱J�zu�'����?	���S�4�;v���HP�$��Ы���Ѣ�F�:V]�RU��|�ҡG�I}���ao����T��Ĕ� ���I�d�	ş@�)�Ny��vӠU��l�!}y��h�'\(F��b%h��ʓA��V��g}�rӜYy��]�u�6�rAH·޸Z���՟�mڣ|!��oZA~�M4}~��S�'�I�:�,<��/`R,K �2P�ry2�'�b�'�r�'�^>�;q��
�B$zW�.PA�q�����M�(��?����?�O~ΓoǛ�w3$�H�gP�.�ؑ�F(A�jZ�\7�':R�|��T�3iߛF?O� ��� #�$�5�˙,�|0jd=O
0B�� �~r�|"P���	���HP�R�����_��P�cş@��埀�IOy*}�F\�F��O|���O��$J�X� Aj%�/$Y�h�R�>�����$�O��d ��^�{�0 :w� <������E�Ri�	R]�R�V���M~�娟��	�Z��qZ�iU�b���2��������ퟘ���<��T�Or�A�G�����ƒ�c����5^�t�0���O��Y����?ͻ_�Diī�W�����m�D��?���?!ł@�Ms�O�N�j��S�q�,�A�� �����A�5�*q$��'��'&B�'#2�'���rI��za�g��d�(d1�R�8��4sp>$���?����䧕?iT��44�]��l�7�Ȁ�t�������X�Id�)�+gӞ���lUco���4GD�Y/
���hӺ��'!*t{�@o?QM>Q(O����n
��b��Ї�=~.��t��O����OB�d�O�<�0�i�谳��'���:��ԨY8 XpS��>/*�I��'(X7M'�ɬ����O��D�O�4!�k�u�̱:s֕�TP��F��4��S5w��01�O��O|W+D�t���[���8L�<��w��y2�'��'���'�2��"vL~�)6b�Q|Tizg��:}���?�d�iPC�O4r�d�6�O��Q�֦Wo""zJ� /�b��O��$�O�i5,v6�-?�;HP�d9פ�騰�!�W9<�6@{&���?���#�ĩ<����?����?��(Hj��@q���v�5[Ce��?9���DƦi�'៘�Iϟ��O�$�+`�R*~Й�񢔚X��(�Oʅ�'J2�iN,�O��-C��
���$\$��&2 ��2k��+��mK@'?ͧ#U$�ā��1�$� "ھR���XS��"}�������?���?��S�'���Gߦ��5iV�m<����Ņ�uJ���H��d����4��'��듐?iũ��C���pL�M��Z����?!�1�(,�ش������?�'ͦ�GW#)Dĩ�F�[<Z�y"W����ߟd�I̟`��˟��O�����N�!�l3�T<>�{
r�<3��O���O6������]#Ev�U���$)�SL�Rе�	��p�I<�|�b���M�'I�X��*Gh���S# �zY�'�r��j�� �0�|�Z��ß�"��J
<�J����I�I
JG��ퟰ��ޟ`�Igy҅f�����O6���O�lȱ�I�W�N�!�Ñ5Ub�1#/�������ON��1�D�)ea��S�`~&��P��"ro�I��� eL��J~j"���l�ɔ,��}��J��"r�d9�Ş��H��П�Iџ���S�OTj��f��IRm13DJ�q�B�-���h�
d u��O��d���5�?�;
���sHG�/��@PᇃD��d͓�?Y� ��/��&���P�A�lq���Ј
LȔ@͞'Q�$�t�]�5J��$�,���T�'���'�2�'��l����g��b)�j��#Z��H�4��P�/O��$#�	�O"�����b����-άn�c!OAk}��'�R8��)��
`z�4�ڲo�� tl ���ҡ��-F��	 rE}���'��Y'�t�'��x��ϵa@�H�k9@�FDr6�'X��'�����T��z�4&�={��Y(��SW��^���Ԩ�T��͓>,�V��\I}2�'H�+e�jD��A��f5�5,�@�����,4rV7m5?1�"�S��)>�S��!��g�MHY�!&L�	%t�`BEn���IşX�I۟|�Iܟ��%��6�zy�'J+{!�t�ԝ�?A���?ֶi=f��3[��۴��B6i��W�'72h��ខ��5*đx�c�V����	�P�{��CBi"��ņ��d���P�რ��E*L��M������O����O��d�(}
��0&�*���a�ˊ�FX����O�ʓ3j����>B��'WU>i
R+��v�x���	N�MzH���*?��S�p��4]@xʟ�Hk��D�:��7d;?��V�?�.A�A���we�<�'�~�����@��sG������q���!���?����?��S�'��$�U;�O�F�V�#�����Ek�D�2���'�6M;�I���l�I�w�� �}�'�0�P=�����tl�TZ�	n~R���8���t�� T�f�9�d �` 5�F'WP:�	Xy��'�r�',��'U�Z>	��@�p��#�K�w��Q"��,�MC�&X��?����?QL~���'K��w�K�3��`�'��|j�ڳD9�?1���Şrys�4�ybA�I�^�,��`�	#c���'K���@㟴0��|�P����ϟXC���?�j�8e�߂o6t08��S��l��ş���Jy�FfӼx�/�<���4��W�B�~)r���?p):�1�-����$�O>����;�t��4�!6b!�!�4YF��C���ŉ�!#����|Z�i�O��y��{���E��4���g�V62w�����?	���?a��h����I'�܅�d�BO����+���$[ۦm;�	џ��I5�M���w0�� �g�10�={Yy�BE@�s�h��4���Ox�LIڠ�t�(�~º�*`��T �p���f�Ӱ����U�,��H�H>�)O�	�O��D�O��$�O&4�SɌ-\Z��D	�|���Ƨ�<�мi����#�'4B�'+��y2O͘ $F��D�u��I@.�@h���?1�v����OY�4K� �P3/0S��@`���k���9 AS�2��I+R��s�'j�A&���'�vdbs�[!�b�J��L'o�V��'��'�����$R�lR�4'?����P j���?wVNl�6DI�Tj��x��OC�����R}R�'���'�j�j�U	L����͓hE�Q�W��*%�Ƙ����!���4�I��j �5�k��<��']�*�╫!<O,�D�O����O&��<�|�ge�8��%r�I�O
��A'S�?Y���?Ie�i���ØO)��s�\�O�y�N*yyxm{c(E�Z�v��@'�W�	���mz>�p�ɦI�'ڼ`j��ЅJ �"�/D�#�8���oF�3�
A��,b��'��i>��I���ɡ_�MP���\��Ċ�3��x�Iϟ��'��6M��T�r�$�Op���|B��1휜 V�L�V�@�9��Y~�>9��?)I>�O^�r�g۴w�l�A!k�1W�"��6U�����i<���|�bG���&���T�C��P�Г! +Ĝҕ�H�p����`���b>�'��7���x;0�5ɉ�fOjA	����	���O���D֦I�?�U�4��(v�T4�C�Y�TtD��B�{����ßd���ئ��u���Tv��<�T�.6x|�rD\�]�zX�G���<�*Ot���OX�D�O����O��'2ᮐH����!cL���I?e(ݨҺi�jM�v�'8r�'b��y�a��..�dJC͋�Go�5�Z�5r�D�O��O1��x�/i�B托)�b�p
�	�$�"f�9L�I��0�@��'h��&���'���'�6��$�\�l	�D0q �,B]� �'l"�'I2R�tQ�4[�~�h���?y��5:׉�vm���dPY�9�R	�>���?�L>��^=?�D��-Ӡka �B��n~"D۰A�&]�g��W�O�"A�	
WA�&ar,"G)X�c�`4�g"�?"��'���'j2�S۟@3�
X�vT�;pl�v�)#�D��$�42�҉����?Y�i��O�ڎ ߪx�O؜�>٨������OD���O� �umiӖ�Ӻ{�/N��Z�MJ��
x����"x���"#K6�O$���O��x0	 #E�����c���֒��!�4_��}����?i���O�L5[�cH-r���P�*��>���?�L>�|��ұa�4��@��7�u��dO�&6�	�B���S�����(�O����u��
C��+ҫĄҩ��	��M[���*�?9��
m���)�8���s�bP)�?a��id�O��'B��'&'�
(�)��D�'nVꭐ�c�s��Ͳ��i��	�-y̕�E�O��$?���4ڐ��
J~A~e�H�3,���O����EO��P!@S�[3u@�=�F��(�I���3ݴ/��l�O��6�?�ȧO��BI����N�	X��O�D�O�iő�7�;?��b�:���
E͔Q�
'{̸AKѼ�?�l0�$�<�r�ޕLgʠ��?���sJP��O 9oڭ1'0���؟`��h�d�H�`~*�nO�/���FV%����\}��'���|ʟ
����rMf��%g�`p���,~^�[�Bc�dؕ��4�^b?�I>a�'] x�b��ۡ��Ձ�� �?���?���?�|�*OzYn�	@Pةo�@����Z�ǮP��&�ܟ��I1�MCI>ͧ$�	���UoZ�OL�eۑ�
'3�l%Xs��֟��I0���l�h~Zw�5���O�l�'���@�a��4ʑk¨Wv��'�	�	��0�	ʟ��	T�$D�y�6���aV� ��� E�[-6�6��(w4ʓ�?�I~��$ԛ�w��d��+�;v]l��+ѕt�)d�'9�|����?��9O�A��*��}����cRrM�d��<OD���Y7GЭ�T�ɻ��í	2|�J%C0�ޝ@)���j��&�Fhj��Y�iwD���0u�T����
��ȱ1�1�0F�  R���5Q�/W<X���q�Sf?�FM�?,Y�� ��%�%ò'zy"N�i��0,J%��)Sƍ�BB�t8�I
mՊ��lD�$Q��@�o=u5�����V	-�l`�c�j�N��%²=^�EqY��@x��
�@KIjR��!ߚ� 7f�1�0�U("
IJ�i�K�,W�:��GL�A�:Q�%��P����6�]�E�,���;> ��KǨ_��M���?q���{1r� AGTZ��!��BC�f�'�'1�	���<�	��~{�#[
KH�)S����^6�O�$�<�qƃ�<�O"��O�~���P��Zaҵ� t 0�hS�.�D�<�Ix���IB3{ֲ�q�A
"ז�����yP�v_��T�+�M+U?��I�?�y�O��BJǚ'&��	%_�Ia�i�副�0#<�~:��S� ��-��?�� ��m)�% 4�M[��?i����0�x��'��XѓLW�cD�HXb<���:�~��}���)�'�?ѧM -jd�bđlH<A�&)�
U_���'S��'���Y!�+��Od�D��4r�nE�G4R�Cn�x!
�
��4�I3h:`b���I��d�ɺ�UQs�X�:<�x��T*6���4�?�� �'z�Ob��:������ �ށ�P�~/Yye^�����+���$�Iȟ��'dȒ��S�}�|U!��� -��Ӥ
��i�>OJ�D�O ��<!-ON��e�׺d��܋Ib֑kC(�,1O����O���<�)D�D�I�N�����T�6��&+��쟴����ly2`C����-;m�d�A��T��[-�82 ����|��ǟ��'
Ș�D#�IN[�? ����oǄf�d�Q���p/�6Cd�`��=�D�<�SHB�l'��  `Z� ࠃ!Ȉ#<���l����I\y�G r��������xR��^-��8c�
�"un�B��YJ�	Uy�$��O�S��ީZ6Dܡ�ND���Ԓ{6Z7��<�F
��"��&��~
��jT��`@Mȸ5<�-хC�8~��j�'tӢC�	;!:B�P�&Ϲ�X9P�'ց|47-��9�`�m����	Ɵd�����?�ʒ�5��Q��Ԡ$�<�T�m�a��'vl���� P��`�E�Уyk��C��n����O
�d�,Q�$��'������mby��iF����d'P{��ml�E_�'����͟��i�a�r�F9�Ж�]�=:������X���q^��q�O
˓�?�J>��F ���q��%B�)�cѰ�B}�'4z1���'��I֟(�����'����
CF ���f
<Vz��XW�;$f����O�O����O�!i�晌���F���.	����*S��ON�$�O����<�bFS�V����6�n4��d��RE2��`�M�*O���<���O��d[{� �E|��83�glb�A��O̮PV�T�'��'XBW��ch���	�O�8#��I��|�G� W)�0�h���Q�	Py��'�R�'�.Y�T>�@��H*%�M�@���H��T�b�oğ��IHy���[�"맒?Y����#��9��4K�a��~�D9��B9Ɖ'�b3O���R�$�?�s�H��:H�C�mSd s���<>^q�i_"�'��O���ˇ	�z��ySaiF5Uv��#��妅�	���;��I}���ON��d��p����������q���M+���?a���S���' e04�M���#MU�t�����oӦ�8���OH�O��?)���BS
X��D�$G�@�%W�/���:�4�?����?����3D��dyB�'D���=B~̙�b�<����`�ǵD6�O���Ӫ1��ON���O
�)�
%da܅��Oo�l(�ceΦQ���%в�O˓�?�L>��kl&Y��ᇶM��H�>o2x��'� ����|�'�2�'���YNM�bVH�
�.�nuB�����.�ē�?9�����O��Ӻ��	U+t�b@j�<�j��ϋ��	Gyr�'eB�'�I�X���
�O���Ƞ��c�\���O6.�n|Q�O����O��O���|��	ZiX�A�x�s�=J�m*F�xB�'��BH�\���'�����pdX�����"4[�l��0�	cy#;��AE4Y���X4)�4��ȟ�L���n����Fy���9"r����$��klFĈv�>�$\�qe��qq�'|�	����Iz�s��]>lV6@��˕�ְ��Ń nq�6�<��!A�s��E�~���z����@1���q^��w�.K���s�'k���?���(Y�O���Mk��'1&Ѱ'�����S�[ئ}�!럔�	ޟ,���?����ɐ'
I(b��D6S������h�oژ,��e3�E.�)�'%�@Pr���8*S�%q�'"�d����i<��'5�E�2ss�)�H�,3���8�x�'!�)�H��s����'n�+�n9�i�Ol���O0���I4XaĽr�B�U�P�&FT��9���mX��K<�'�?	I>��-V����Xd.HY&�SL\8�'@@p�'H��ݟ$�	��$�'��q{uAܚ�B=���s��X�Q%E.W��Ot���O��Ov����5*�:k�`	��_$bҡkb����?�/Od���O����<Ag�Q�R�	���$j�-�5i^B�`���,��۟H��[�[y�
c������ЁWb��(dMs���V_���	�����wyrǂ�m��8ā5I����@�	A`���2�Z����	�D�'���'�n�[��'R�v/"M@%�:杀cׄ1���o�����|y�K"y �t���klS:kNL��Q":lu1W擽	Ӊ'u�əy����	F�D
fˉ�;�uв�|�P|�P��J}��'�����'�B�'�b�O�i��J�l��7 ��x�,6vm��(#�fӐ�$�O�U sLүk�1O�� x�ΗE�􀀷- �B1�N!m�%W���	�|�'���[��'g2�
�c��K1l�q�FY,M���w�ift���Y2͘����p�%N�$_R��C����oN������$�	�k��ɕ���:}�F�2�|̃�eK�/J��"d�"f��c��y��ʝ��'�?����?�Rf�2М��4'�+\M��2�*	�`*�6�'���xĩ>I.On�d�<A�����3
�ԙt Yo�`j�PN}�,:�y�'�r�'���'a�3cfԘk���1���a�2K�m�%c���$�<������O��d�O�i��x,��A�K�JM�f�$:-�<���?q���&Ra�DΧ$����I�1�ȀС�k��ش���O���?���?�DJ��<�C����5;v*#����hR*y^���'�"�'�2_���F-����i�O�"���8Z��b#��T�!� �E�Iuy��'�'���K�'@�i��b��@��Y���5e2��3bf�H�d�O6�=1Nt��R?A���<��-<�Cr)Ĺ0t��"�D�ҽ��O����O`�����'��',�ɉ�w�^X�#M�'��x Mџ.,��^���U�@��M���?����j]��=� `��Ql�Q�nM1���:#���R��i42�'�:���Ojʓ��O����ÓA�v )���z��42J�|��il��'�B�OM����C{d���LFL�\�B�E�n	F�l�\r��ӟ��'1�4�A�i��
%y�P)e4?��	o��x�	ß�ɦbU���Ī<	��~���j�L���(���������M����E��?��I������j����3ƘM�����*z���۴�y�I�'#��zy2�'\����ؔYd�Yi�B�g���Ѭ��KZ��{���?����?!����9O�l+Ѧ����A�# IcJ삢��8l���'@�I؟��'AB�'`���2�J5s%��?3����"!֌y���2�'���ʟd������'2p���%l>1�D�Z!R,Ҷ� !o M�j�x��?�+Oz��O���@�O���5x$���o�Bh����(A~�nZ����	l��oy2/��D�2�'�?�v����s�U�H���(�ٙ6����'��	џ���ןd����[?I��D�FK���㌟#TeDe�T��⦅�Iߟ��'b�a�L+���O��F�x{I��Q
t��P[�L� s���%������C�j�$&���h�������s#�F�lm}y��ӁaF6��V���'7�t$?q�d��..XdQG��UN5hC� զ��I˟�8�@�$��}��F^�T\��%��0�p�[1E�Ԧ��F�J�M����?Y�������^�p�,�!땼	� �!�"]`��l�M:�	r��E�'�?YYy;&�I��Z�u�#�c$L	nZϟd����PY󪄗��'5��Oj%)$d޽6a6�
�e��-�X����đ��(�O����OP������h��7׾a9K�c4lZ��P�q�ډ��'5b�|Zc.�,QA�׿:��[�(+J� �ӬOYۀ<O\��?����?y-O��i�*[6lo��2W��z��$2`�� R�Bh�>!����?)�{�\���C�DB0�xk�)�����<i,O��D�OT���<��"m��iZy@8$�\`���B�	�'�2�|"�'�R̎(:B�$'Aĉ�mR5Xl�[��	G����?����?q-O�!#�VM�q��%o�CV�w��/Jfn �ٴ�?yH>	��?I��<�M��fDǇ� �����;j[9�Ԍc����O\�`G�Ts�����'��dE�pXe�'�ީVjzS�"
�Y��O��D�O$��=O��OX���!_b�X��X�9�X����C5t�6ͫ<Q�� ����~Z���Ց��#��YL�
�����~�j�EmӲ�D�ON�y O�O��O��>1;�L�)=�d1ckϫD�|a�!kӞP�7��֦a�	��l���?�Ɋ}�LT,6�;rꞘ)W�A鴀�!T{46M�PZ�*�� �Sߟ�XDM<n��2*ԶE��i"A�Mk���?���M���v�x��'��O�Q�ኄ	��D* �Z.B�҅9W�iH�'*>�yP�,�I�O8�$�O�t(� �1��1Y�C�����զU�	5(0|�8J<����?�I>�1h�н*���%:R��閛"�L��'�$`z��'������IޟЖ'�fIxb"�'hy��3�P�ծԈ�kF'ބO����O��O����O��ڵo��o��-[��1FZ��8%
c����<����?�����$�e��l�'z�@)4�`!pͺƧ,��X�'���	~y��'i�p�k�&Z��8��H@�2	&Ϳ>1���?I�����5"F�%>�Z��I-�pr�	t(Uf���M+����<���	%6�9H ��(j�QT�{Ԃ6M�On���<	u!_ƉO����5V���`g�@*a���v�I a����'p��ܟ��?��\��:gbF� ��$>L�2��'
��%%���'{��'(�d_��]+Ǽm)��
"�U�.��Mj�6��O��ExJ~"�	Y	�v�*�*��EQ��lӔi�0�	�I韸���?A�M<a��I�>�bf�J2Ԕ���ͶX��l���'	���pH��F�V%��/i����i���'!���OH��O��ɗ3�J��bi�)1�}��j�w4�b�$z�7�	ßx�IǟT*�N˱cT�$�KTJh�FmG-�M��Ry�q���xb�'�b�|Zc����@�)�d�C��L�d>�-��OX���d�O��ķ<Q�p#�8At��i�6}�U���:�Δ "����O��$�O�O������Z78��$�%N.~?(Ă�Dpӎ���������~yr��(��S�u
�hx]p�1f�s���P���џ�'���Q�-��!b\�N`�\AS㓴G*���'���'�RU��z�.�!�ħ3�Μ�tG�H�=��W�r#,���i��|R�'�Q��0tnՒ=���P��6 $� d�P��OH�ɐz����'P�toՅS�NO�Ȫ̋��_33�tO��D�O����~*��R:��D�,��M:�#[�E�'��tr�<E�O��O�&�	\&�i���<"P[\)(1��m�ğ�� �#<������'�.Q�`N,�@���O��?��j�+7��"�ϟPt���I'��ݪ�C�Ib�5����OB�Im��ׄU�J��a��M-C6��% ��vQ`�
d(�
̄d��⅖@>��V�P�V�ځ��J#W6f��",� �DX���m��]����)	�ۗ�A�o��18f�ܠW��i�SB��g-r���y͜�����51����D�{�F��<�H�bB%.׍q(yqS���?��?����.�Od��u>�!�B�h/��!��TB~����ߴ-:6�� ��	J��*�"ʐ[*��d
�=% 3c�#i��P3s�3������6*-���D��I�0+#H�
Lܸ2�'�I�V&PMQ6��$��&/�^��P��O��d$���'��,HS�Y(M<~ �V&~Pa�' ��MU3��B�Ȏ�N$��2�yR'�>�)O�@q�NB}��'�차��* �icP13��b��'�� �V B�'��	H19y҈k�\��\Hc(b�\�xR9��8��	`A��ڤ�'�4	U$��DB�1�%L� H����A��-�E�V
rS~��� A)�p<ɇ�����	Oy"�>-�LHұ�бb���b� ��'�{��Z5$�PpQ��&�BhA-� �xBCe�&-�N�td�f�6#�;�=OF�?��A�"T�4�Ig�dcFo�'N�<_x�@�c@2#� 9��@8`��'+�����͋��Q BQ��T>)�O�;R�W7
�}�� �/I�2!ZN������=h�0�C5��J.�dG�$I���hҦJU��Ĕ�é�;��I+--R���O@�}��b�MzdF?јY`VdWx�i�ȓ[V^��H�rv�KÆ���(��	�HO��և��G��يb�ڇr�9��^}��'���ճ6���C�'�R�'��w��|� ��8U�*�ce/\آ$Q��ů,��9�K�Ob���	�1��'�@�V��� �������˘�M���Aqi�Op�AS	�����y�����Y��X��ܬ_^�	_r�j�Op��������I�_\mQ�L8�H!�(�/dC�ɮj�ڑP@�Ukt���f�4-�z�{)���'��d۲>|��r��k�&ƀ.ʄ�Y�<D ���O��D�Ox���?1�����P�{�����c¨�@aJ1<�j%�T�8;XѢ"�� :s�yR"%x�ȉH���1
 ��%�2��˄I� 3��8�dg��y�)��"
��U�]=��dɆ�
�ry)���?y���%��#~-�̓B��▼Jt�f=D�5%��y�����k�X���>����$�<��Ē����'��DV�6TL!��}n�c���1!wB�'���'�'�r1�ʥqw�	4](O� �"a�)pu��j>Q�7�'��Dh� �1NA`1a�/&�1w♄]��CE����qU��D@џ�z3��OP�d�<Ѱ��9Fi�'��/_K�p���<���?������BM�5C`a�-I��ժ�oдbO!��22�TE�)cn�< ��<A�f�\�'� ð$a����O˧[8��p�akPmO�K�(	tDB4O��=B���?9Do���?��y*��ɲnezU��#��Ȱ�+�{V �' �-�����G60:��p�L�$��-⅂Ɂ'��'M��	P�S�'-�8�&<2)��҆�je�ȓ1��Y���{����c�����	��HO��*#b�3n�� qTm�V���Ab�˦��IΟh�ɨ0q�#I�ɟ�������iޑ�N�tG�,��C#��;7�ɐ;�"4`��@�Lf���¢@SD��|&����͔G�&�[�q{�Ja�	�=�P�K�"��L�� ��'V@�>�O�|���+L�ر���h������֦}��П�PM���Sҟ��I��	ݟ�x"�ߟ3}XL�f�&��;GD�Lh<���}��i�C�ПxF�d��A~bh9ғ<�	sy��ɞb|9T q�-�k��u?ΥH��Q�A�2�'���'f~��������|e�D&u_�՘$
��}����&XT�����V0����B7�h9;FN��pf�x� �b<��Ƃm���8F^��r)�Ǔ�9x�(�IN��,S2�׶9r�Q,5�z��H�c�!�dK�<u���f��P=�9�SN�Uh1OJ��>I�AY�0���'���$(Z��cS˅+�,<hF�׽%���'�nd�!�'I��'[BU�oK�=��OP�ąX [����Pk�����'�ڬ���u`bi���J�g-�q��nH3\jP7M߷Z�d}��IBv8�`�A �OX�df}"��W@x<��DMx�XM�M�y2�'H���S�mDy�$)�X�ppҋ�ja�hO1���ll��m3�G���	 fo�.d
���4���ձ8qHqoZ�x��A���ݤB���*<�tmч�S=w_�}Ӓϔ$���'��i��'�1O�3?	F���t[�tf�ɟu��ɒ��E�$Ԉ	���?�h�Ìp.��gg΂8QQP��*}�OΜ�?i�y����3R�2i����^H�x�?�y�
ހ<�r��tHήJ�&��e�ܠ�0<ab�)� ���֠ɄK�"�����z�f�����	֟��I�kV�0
Ģ�џl�	⟔�i��b!�W���:���k��5G(�@�H�Z���	~t��)Q��ڜl�b(�<1��XH��+<O QaN�/{��9g�֪r'����!�	�p'����|�P1\^��%�/I�	�P�B��y��]���q��8T-Pʀ.��]@���8�s ���e$���$ �dH�� V晙{ڄ�A��O����O��������?a�O5�Pp�K�[�lܛFG2�0И !^�dD��'�����D 
�(���=ŖLTaG$f
���'
c	�2��񃰆���ܡ6B^:�?���?����$�O����R��*ePԢq�6M�lj��;D�����O�����)M1���v6�ɥ��ļ<9U�^�Jd���'!"��>�(�@���?`2�@�d��N��'PT\���'A:��E9"���a�Or�Iv�K5J��\��&%`Z�u���'���1b��d��']哅��9Dɠ=(��!$���ǓJ�%�I����ן,�׎tv�Ѓ /YVoZ8��_cy��'I�O>1p��Z1�����)�v���=�̋�4V���g�J�m�z]�lU�@mϓ����󙟰qc�2�D藄
��D��7D��rA		QV��:��ɑ&�@�(�6D��`G"��H@�)8��E�|�ZX#4�2D��"
�����D�_�hXc$�2D�̱fBD?z��4�A͈�\`�8��+D���A�K����N]M(�l<D��J%�M5 �(�80�ʿ�y�d"/D����V��d�6'�
8�y�Rc-D��8��M+���hCJ��1�Xe+D�LC�N���d��D�>>���� <D������!�:�,سK1tՑ�7D�p�B=u����tjȕhj:�!��3D���@B��� �3��*s�8�҄	3D�P���k�l;%J�r��u�e<D���QoΆ6��	� �3j��YX�*(D������$���ΈV"l��A&D��E�� �z`��HèE8� D����0�<1���6T�ᱶ�=D�4����4h&>���c:*��PA�<D��!#oT)0~v]!����o$ۗ	<D���(�>]��K="��hp��:D��c#�8e%�$9��Ƿ+���f�7D�T�wN.( Xe
ı/a���0D���H�!3zQ��h�71�-�&�.D�8C2a�-=KL��eǀ� ����֢9D�����Y=71Θ���:zk�"D�,B6��^�љ8H ���*D�����ǉ
t����K$��ى��<D���P/���vn� I?��c�K6D�H�cNق]-HH��J�jR�9"''D���6���MTp���b
V()�s2D��p�X2԰)���k�́&C#D���+W�`�rIh�兴(a���	#D���V/Z�B�Pp�?Z�(tg.D�X��ñ�X��F�j, �)D�����M�R`X}R4-B�_"I�N(D�`z!K<� A�-Kr�&����0D��C��ɇ)�`�s����q�P�R�<D���ԡF�0�8(r�Ѳ~8�+�k<D�8'�-$O�ـ��R!w�X�*&D�$(uo?WS��D��'U��;7�"D� �V��(�~��À+��=:7)=D�0�æ�R\�ɫ�@ ���FC<D���oA�P�� �SO]���'D��	�G�;5�X)G)O�68�AH$D� �%��@[����DZ,��b�=D�� 0�ZU)�5Dɳ�.N8(���"OTE����d�6�{��қ&T�b"O��Z$�Q'��IS�B�t^�)@s"O�ݸ@�вp�,��(�*C並"O�}q�&�tPAf�Z�"Ƞ�QS"OʍZ���l��銤�ġ@��|rt"O�5A�7h%>`��U�g�l�#�*O4Y3�޾71�i���	-66��	�'��ݣ��Ц`'R���jS�E�
�'�Vy��(a�^ �c�X;
�'(1��C�&��܋��p���'�P��DA�|Y�=�S��!,���'7N�+D*�.T�rq9�D��u|,���'W�m�&�U��r 1�͛bɎY:	���ɂsb.LH���t���f�K�<��kK	 Ѷnǅy9D����J�<!�@�g4^�
6���[�Г*VR�<�W%s�c�P�h×�QO�<��FK�	�	��F����M�<���7Q�2���OU�<��� SDQF�'ME���5�h�y l1�$�S��<$���"O��D��<&� }�2�āE�,`� ,D�,�#�	�e�)��,  ���� �<#�:x!CN�D!��J,z]��e݅-�Hd��GݓsQ��ö*�>L��":lO�b�L݌-�<u�1�+X>�ʕ�'�p�X+V&��6@A6a�Lx(@쒛>\(�G��0�y�Ӱ��Ƅ�29T<ѷ�@�(O4A��Ҳ�#}��)����I"f טR}`���
�f�<��!�{����@x�Orp�7��2+7ɧ��Ҏ<r��������0Y��2dMڷ�ybF�\YLp�#7��sk:�~�J�$H����'.
ѸSHU1N� HǔF�j��[
1�Ѭ���M��l3;���%��r�q'ʒ�<���* ��Q�U{��Y�A�R�'L@�F�(�>i��+�1M^�/%���z��:D��&� s��=Ҳ#�i�
mH��zir(r��!��S��?I�V;u������K�p{"�m�<Y"I=�����9j��!Ml}R�F�z���Q�L^�`�gR�f�	�v�K,-�ɀd�~>0��'R$҉𙟌K�,�5K�e� g��lL:)�d�%D�L��M�c}�824)O�V�,�I"KĶ~Д�qV'�!G�����@f�\�Ƣ�#>��0����(5azR�`r�ܐ�I��y�j�	��Q��aK���0���y�N����ЂBG"n���`+���'����+�=�$0����M6?�U�@S��)��Z:�!�䙇� �����g���H��R�Dp�Yxp
��n��	�h��"|�'?t(a4Ï/hR�c&�t4�@R�'r\�Q%#C=_�DU`����j�ƕ
��Q:"��%KU�0>1�\�֮�C�5T {'#}���awɛ.���ӑ��x!p&
2�F!�Ί'���K#i<D��aBD�G���9�o��F����d�<扞B���䧝"L�"~Z���=���$ Ϛ��p5�x�<	���k��<��m���=���ݳT������Q~�+ȹ����/qR*p�Å�7DjL��=d�C�	�#h ��u��"$���ܬ	BA{�Z�ljRA#�O���[�l�5[¯ >��8��'ي�� ��z<��'f� ��7g���F�%&�j
�'�kQ��
�ڍI���͆��y2��Ŗ%�D!����D�; +ȨHX��j�nM�[����"O�y��ї+��%�!�S�"�1�W"O�\ZT�1��(2V�e��z�"O��Y��34��12C���yq"O	j��=$�2�	�	�d1�"O�p3����137�T�K�J 3"O� ����ӌy�����6t��h"OF�ǌ�wD�`Q���>
�ѵ"O^��a�44��33@J9$@��6"O�<`Ӏ]�����Z�n����"OFY�A�5� �؂�5j��L�a����yÉ}���'���k7�N�{�gY[ߐYדs)��[J<a��(�f�a��� M+�Ƀ��@?I�#�p��jر|�ay",��R� �q֊�9<є8�i���'���2�D�g���'$��f~����7'���uF .�����Y(<�⌱n��aO/%���MP��N�<AI�u ޖ9sk�����`R?�p���
�Ol�"	^V��"O�T�6�^&nH8 )q��,7���7�_5�zD���V��0�^�xU#���M��W�\��[���v�U)V�����N�,�jS��>�����4US��#Ք	-���%��ȟ�"D$(Y���$��t���1�G�WF��O�T1O���C�4��X$�����?��f�,����,��>;j��!![ ���'=�O���"�?�fu��M�#��� �j��"P��P�����s{�瓽 ;*P�"�'�x3�O4q���D� )����@ҒNm 1���'�R����DyBA�P0�0@[�|�� !b�( R�Ǚ'l0U��%�0L�cV�U���3FC��	�g~"g�e�T8��I���R)�� ��g�¤P�#�<���I�+B�FQ���萳
��A����1	� չ�A�T��FP=Tz0��B�{�$1��EU|�`�T9�FM6E�U��� �fy2e�$��ux���gض �I^��LSB�|�  �y�>pC�R,�j-PTC��R��I���W��֘kvy�dI�M˖3Tx�4�G�%�<A�&�O����
��O��JU�,qV�5(ѫ�zN.�KJ�Dt���FjX�\ &,��X����������ֆƲ;�D|�'���&9"�lˎ%��AĶY�hm��'�v�*�o�/�>̐Ac��Z*O��P.E;5���ԏh
ѓ��xR�_���#ϳ@�ʤk���#1]��7U�p�IR�h�1�;]�I�d�z)��!h��[S��ё������
Yy�'�����ʸ#�̱���Wa䐰q�[�ݮ�9��
l\�pB;g8���fXTa��.��I�r9��O�cE�l;��M,L`�����5�
l�2,�b�O�)��Hj�B��h��d+�b?�W@Z�7�ĸ�|�SHJ�w*Ĺ�A�;����҆ԅ-a�!�A��5��	�K�A��7��ir��>rpL#��åz~$�h$OL)1��ar$�$m�\��C�rĕǢ��M ��ە����=�,8r�z2�>Ld�e�d��Z�d�m�h@�!�/ߚG#���H� ��$�s��R�����QH�J�4:�P�k5��	E�#E	�D,$���	�N����cG¢��1R���Y�a�P"ʹ~��-ٷ�Ujn�)�Q�ؓ�`ׂ?ԩ�O���@�Ξ9V���8J	�!�'B��DJ;f���Y,1����­�\v�b�U��`��nO�ٔO���wG��K�<�cK&��}ҕ���h��J�>������\�&D���@�%\�$�� <y��ɇb����:�����ȉD
�GhVW[��d�z�"Ђ�����ǆ��� :�{�@�
������J~䀈 ����T(=�T�'T$0�0�A��%3�H���GDU̓k���hQ#}G2}§@��w�ŻB	� 4�s,�<�a{BHϷG� s����Y�L����E�}�s{Z���w�<ڄ�	!SN�L�D��9�:�{��nވi�`C�_B���d	D�g~f=A�LНI���Pm����
ܛ`�Z��IFkT*`F�2u��0�ԉk3G.�wIh�H�ػ &��r.�1���ϓ}��x�W�~!��c]�p�:4�O��@REך a�tj��:O"����$U�a��zu�[&JZ��hte���$Q�׺d��M���6�:�$E�!B���DK(l��H���;W�x�ʧ�Aަ6�-�i���'uz�"��	p��ɕ\	�U��L�'���`'��wL�U	�X?Eځ��dؕ��+�H�֔a�Zn�&��ǅċKY�� ���)�:D�'�.d{2��i��9i:E��g��J�d�p獦R�HB�̄%fؠG|RKY�,���K0	Ș��Ox�+0����$�2���V���>�a��7n-2�A�>�&����D� 4����R��ΐ T�!y����O�$s�1$�ˏ�D.^�4�x"���5�T��'���EZ��E�g"j�X'E8�ʰ��ə�ڔk�	D����b`Q�+88B䉞�v ��BU�>�qB�&jrB�ɓB���qW�Y�o)R�ɻ%nB䉏?|J�P���F+L�K"剋Kl�C��:~(��W=�����&y��C����Ɓs֜@A�X�B���:D�L+��C�e��5��e�&1݈���M-D��IC&\�>0�E��2!:�╁*D�� hYkV�]-F�L

s�y�A"O�LR!�M�ȑK�
ٕl����d"O��IcHM2qG�ة$DY4z@�{�"O�8�7�֊,��L�tcP;�xܠ�"O��h1��2>��tc��t�L�"OD�z��F�H,AV)�~�< "O��C$CV�̅��i�ʡ��"O��H &Kl��Ig�N�w�L�)"O>ihަHPB��0�C�y� 	+�"O�=y#����+��g{�=	%"O�ai����
|���Q�8m61	A"O:iSə|^@E e'>zP$u�"Oj	�n�!-�|D�ϞzQ�EKf"O�e��L�H���#'dR�Ej|=�"ODqx�a�S���#Z1;Gx�� "O��)��� ��M��D� 3TCP"OP��b�ݗe���1���"rl�c"O�䓡g�

�Ɲ؇�Q�al��"O�HA3�8A)ZQ��Xh$T���"O�9����2��ԓ��3��9�"O�x����/	���l�n��9�e"O^�)b�B1�|9�AlD�p��	H�"O
�7�W7�HA�kN��� ��"O�az2.U�n����1@��9ȥ"O<P
m�W�����$�$�#T"O�i���{4$��(�.{жIs�"O,�f�_�Z�X�PG\<�~ �"On�q'&�-`jQC&�%���!�"O������H�G�xf��y�"O�!A��2��J��5���q"O��[D�ΜvL��*�B�@�d�p"O�@�c��#�"�K���!I�� @�"OJ�!�-
�z��຀eېe�N���"O��H�e��|���E�\����ZB"O{��	` T�g�	 �~��"O�yq"��$@��%�;�`8E"OhIPA��ZN�MJa�Ԗq}p	rT"O�e[!G�,|����A�N6m|E"F"Ob`�C'�YxTr���aaXh2 "O�M`�i�2^�|J��+S�A��"O�)���S�?�\�	�fP(O���"O��ɐ�F*7��3�KWIA�s!"O�A�  Rɼ�z��ɪ)F޹�s"O�H*�̑	,���GO�&g�|CS"O�虄��z�i�#�wj�詖"O�B��1w��]/qwj0�$V��y�h��t81�En]%h��H��yB$�`I����ŧ8���q,ܕ�y"
R�n��`"�g\�%F�8�7� �y�a�V��A�O�L�r�
w@^��y���1@�#�n��Cr�k�&��yb��'9W�| �ۗkyA����y��&,����r��	.tF�21.��y2�Ƭr6@u�㎁/9��)�C���y��!@��H1�i̅<ښ�z����y��ի/�t���-״
�`9`��7�yB��"4�}arN�s/�0Yb�Y�yR�?;��̄�7�rtc ��yBd�8���e�-���X¥I��y���-`X�C��U�u��p+�*�%�y�e��t@r2���m��p��"�y���(S�mڕ*�/�vqÅ��(�y�┐-����p&K 8m�U�֨�y��ށqK�K�Ӑ���҃,�#�y
� e+���5(o:xJ�K3�|�0"O]!�9Q^<��`:_HY9"O�4V��o���r ��{��,�"O�=y��	�i��R��(k��-R�"O�,A�H�Ktl����?���id"O�#���4$�ҭG(��x�"O�qKB�Z�� 3�M�~�><��"OH��f��9g�X�`�Ą�"OF��C"�x�d��A��kcp��P"O U�fB�8@ܹ��F�Ab�A	"O��bm���A)�ϩY[ (��"O4��dƂL���0b�W�oN���g"O�*��Z1��j5Z(5�"O<eʕ'�n����f�mq��W"Op��"^�`��#\oa��"O���ˍ7/8��1e�xr��hV"O05XDkP�+A��.V��HY� "O`l G�Z�O�ր�gk1�4uc0"O��A�X�`�:�7a��j�pZ�"O����:&;:��`Z�4&�'��OȈ�v�J!n	��Ѵ E�>t��"OU�G/T�R\zd�'�5{_B��vEH<9vj\�E����U�*����!�\�<���'?�35c�z	�����a�<) (]��;@m�Y���0D���W�Z�.��)��)B,~B$}y�*D�p�G,Ĵ���M �*��(D�XHŃ�4 ��P�$*$���K�(D���7�I<�\���8Ns��(r�:D��%/������e��/r^�8��.6D�T"��7��A���_�o&vU��5D�𚳀�)=��awEI�z�;&�1D��@�`���A8�d�8O�� P�-D����ꔻH�P*G�Q�=g��1$�.D����W�"x:�
SHO�F^��Ō/D�<�")]'��`2`ډ7�)���.D�4��0��]h��يΪd�`(D��j@�n�!aǛ�x��d�,#}��'E4���㜌s�(��6��.$tƌ�'���u�����hp��/!܂�
�'ň�!ʛ�2db�ôJR%g٪\r��&�&����S��]�M��P�ꅾ#���B��i[� zA,�� 8�y�ˉ�I�A��Q }Q���_	�y"��
D�&���l	v�	���4�y� Q)�����bP�!��q�F�&�yb���&pt���m� �F��'�yRIɃG�+KY/E����6Z�B�Ɇn��%8�eN8�!#��&��B�Ƀ�2���!�&p��)?\B�I$n�&-�d�-\�<����\��B�ɑN).���)�Z���F�(,~�C�	�	b�L�A�Ԑ&P�	!���7\hC�3Hx��\6+~$�6Y�5 B�	<s@�:a�S�Ȳ���
T���C�=�@�!ɗ�Q�=�)��#e�C�	�RZ(I`L��e�B��D�͓U��B�	4LA� ��s�(H�a!�;|��B�	�q�4(
4
� kc�0�S�+|��C�I����� �	g���)6^�!�DΣ~�l�
s@�?>�����i��!�D߉l�<(��f�;�&Ei����&K!�$�>lc�`���,|x�i0�ר{V!�d�%�e��Ƈ��>�R��2[!�� �}��Ю�Ƹ����Z��"O2-��NU&02ub&�O7X�4�B"OF]!pʜ�[���3��'t����"O�8�&$ rQ��hg$�H�2"O�XQ�H���HmρG�-1��'!�OQ(� A�6 i�LP#��3�"Oh3��if�U�""�>bf�r"O�,r�*��8�����Z3ZTj ""Oм@r�P^[�Ԫ`�YlՐ�$�#<E��2'��R-	�,F>e�UL0󖍆�q|s'�R�:M
8��CdD��'S����I�Xu�Ex֥@1SI���f�H4l����$@��y�i!�U�
ΉzA�����<N�L�
�'82옔iW� 	� ���ǅ@}L�"
Ǔ�HO�+���<j�MᠧM� �m��"O�4�tDI0,����a��8��;�"O�iၕ�u^Zu`E��<�^d�0"O��A�H����$M!eu�P�w"ODLH5�ѽ.9@ͳtC_�fh�ࣵ"O�%k�jNFu86�R�
�����"O�E����C��(Y�+A1��IbF"O$��Ԣ��P1X� UA���v"Ol�;�䏇mxl�A@x�"��"O�ՋE�X�X�8�em�;|Z`�"O���'��#u1��0�,�;@�z,)�"O&P𗭍a���h���*��ZU*ON����9����Ǚ0@{�
�'p���?f��y�L�2��'V0���ݳ7 �<��m�I4=��'�h\��1�4U���� +�|��'�:�;�k^�nLs�J�=y�&�Z�'�Ry� d�I��K�o��mr0��'�XR��֮��-�`�=Y@4��'Qj����9Q�ll�l������'�",��#�V8�o�%�$r"O0�H�M��+{���F���
$�$��"O�%p �PB/��`�/�+l��"O�3sM�4lD��$�+zN�%B�"O�b"kW��jQ�
'Ol %A"O�E ���O�H�����h�z�"OT����<8lL8Ǆ͋���#U"O: ȥ��|��� �#Ws�����"O��g@�7F�E27����x!"O���6D���6�"g��Z~, ��"O^4�a�J�@�8I����<t{N�("Ol锯ҒAY�@��U�D0	!"O&�3��� 8��v��%9�,�+�"O�A��gֳ0X.Ĉ�i�m�1"f"O�EZ��Il��1�!�_�Si�Hk�"O8M���MNhx��U�3Tiq#"O8]P�"�
/)4�xPɖ�E	�"O����� :�@�a�P6��kf"O$��3/K�}�6�(�Âs���"O��BV�՝nO��ۧ��Bس�"O� �g#@�|k����h�H�Б"O܄��@H) RÅ�:~�L8�"O>�w�vj|�0*1`�L�V"OU�g+�V��H@�ANzp@0"O�9$�%/+D��쏼67����"OH̓3CM�m����#%/b�""OJ%�k�2DLhx�#��	�0c�"O(����/=|�ЁlJ�Ah��s�"O�4;ǡ\#�X�B�ӥMY\e�@"OX8���n������LR-�S"O� X� uHP*���
���c��0"O�q�2�
f�$�aG��,�#�"O�$+���0��V`3A�\�#"O���!iT4
PHs��C�v�St"O�:�B��Tn�1�AQ�"Ol�#�E�~ȸl`G�ʤ;Fl "O�Գ��Y
kD�	("M��XC�p"O��Q��ϩ��My���F0 䛢"O
$hC �&XpjG��b��E��"OVzwA9?x�K*��i��l��"O����(D`w$��� �f�As"O~��e&�RQ���
�B���"O��q$�y�X��;��0��"Olq��_/$̀Lx�FK��\Up"O�5a	�U&��R�H�9)�,�Q"OdY�q��=R,��^r#�(k�"O�`��ض'�͋���$N�IP�"O��`��9]������	;K�D�A"O@�@F"���(���8-4 4"O���Я�!?Ӯ��"K�k��9'"O���mȀS5��b�o�,�lEA$"O�p�`֘D��KvOM!v�=R"O��0�ȏ�d��X��ԇ=`~���"OȄ���$�VH��'��`��C�"O�Q�D�,f��Ճ3�=R`"�a�"O�M��'_�7;1���}Z�!��"O�|2��f�vp�7O�OK6��s"O�)If��&`�
�	�P8D@��C"O���J�<X	FN
1�U�"ON`�pՎu�B��	����"On����+�v�K��ҕS��#$"O<=����9j�:;�R�"OؕQ�B�!"�b���Z
��J�"Oԁ�ph;R���y ���FW�t3A"O�xT��F |�I�6#E����"O����(C2^xaBcgK��T�v"O敹t�A!,���G��/k, �@"O�	)�k�3@v��(w�U�u��-�`"Ot㢨]�F���hծ�X�+Q"O��:�d� �@�����8�"O �2B�4#��caOMj���B"O�����Q�$A��jN2yJ��@"O�([�*��Q��ߍ./D�)�"O�X��.Ϋ+,mAW��&.�	5"OШ���T4Ƅ:��Be�M'"O�� H��j�BK�'���"O��V�f�Eb��#>����"O&0�#@�	!�a�1Ɇ!�m��"O�	j� '�t��ɉ�x���"O��6FN�j�2(���_�=��q�"O&(r���6��T�;¶�Ȳ"O6��L�!jײ-��ƃ<��|"C"O�Tb�nD�4Jj�$e=Xb���"O��A5��93��g�ςCf1"Oڐ[�%V 3G*�Y�eǯn�^m�!"O�P�%�@3S��ѡQ��>V�D$�"O�,�&����0!̸/�䓳"O"Qq�g��l����o�<<�Z"O����'�.!�N`+���(X4`�@�"OƁI�L�8:�h�&*J�KJ�B�"OBI #��8y�(�s��*j8�tW"O�� �
浡�h�JTL�	�"O6L�W؂y-ȡ��9��Ș�"O�|ipd� OZ�͛"���B|�e!"O� �q�� /��@�ݪEKH�1�"O�Y��Yg�vmVOA�t1)� "O�}:���y�p���M�
$,B)�r"O����f=	SR4�bJ+|P�z6"O�t:���(9x8p��aӮb\��@"O��:B�ǂL�q�f&Z�"h���f"O�i3�P$��BU�,vz��"O|Xcd��_�3&��[<x��"Of�`#�m�t�C�D��"On��
A�<*N��v�1$��p"OJ�(#��=t&�s��ҝB$���"O$a`)�D�p.J�!sr���"O�H���]5�:�an��dlb�#"O������S"�E˂Ï�|P����"Ob�YP�R�Bs��Q�3nN=в"O��!6ψ�z�*@��
8~S��"O�����	6QB�d��ɍ�@:Jt	�'[n͊�,�+PU�y��^*'��8��'�EJ'��y�����"$
p��'S�!�Ve�<���g�/�����'Kl��A�(�rܙC�<cr�8�')�ĺ��N\%�eH�-&���')�0�7�\ug
��Hȥy|<���'�
��7�Ѓ����'�ܟnM؜Y�'ɺ) ��͚Y����M��z��/D�,���7�d�qa��"q��-D��!�$�.�4���L���u�5�=D���/(�����E$�E�;D�T8fN�*sʤӡa·-̬� �=D��q�%ؠD��Y�J*�l5��:D�̰�`�/�����k��a�Xu{�8D�h0Qo+8��T�èJ�z�x�i��3D���m_�/�����;bR��0�B3D����ć)j���r&;vD�1D��Sa��Wql��G�����q��<D�苠��� `�G26f|hБ�5D�:ơ�&^�E�u�i\��o3D��4��3e����G"X6���.D����/�63�|��DDZ.�T-D��Æ�Q�a�0p�CE�|p�r��)D�(r����m��M!p�p�,D�DiS�:V��ipk� 3!��?D��*����v�Ѕy�m�6~��=���"D��Hd��~�a��1-���c!�;D�p1����=�>�b!Od��R��7D�0����$��$D?;}��"D+D���B0���5M� �0�v�=D���l�)VeN<)�9{�E��0D�@�!�
X��	#�"!��M��i9D�\��mL_� ��� r,����6D�l��.�&t}롉ӿ�%���5D�H2A'oŞ0X�敊8���W�9D���oD&n��j¯��a��!��6D���Q���UY �;��O�<��h���4D�����_�:��4�M8+����U�>D�\k��ɔa}�aq��!y�K��9D���H��V�� [�eׂ[H���E7D�d U�	G��a87b����)`�� D�lHa�5T�|u$�32\���-1D��j��a��UX�g�/"�B�;tc.D��H�F�=$�:�y�͑�l�:$�8D��Y�Q�U��B���L�2mY7D�����K�b@���E�˩p�TM@�� D�pH�ϾX0�|�����OGDL���� ��w�2�h�i& N�~m� "O��aկ+&1dl�([&/��-Pr"Od�@�̼t�X-*��L/jn\5��"O愨�
K�-��	(�,��b�8c"O!xs��g/��3Pm�?"5fIZ�"O6ݨ�"\<�(�q�f^���Y"O&A��CE98�̽KP`�� "O�)"��.-DࠖO��9,��`"O�h��̷Q�\��Q�	3�y"O��r6��.��q�@L,mZ�"Oj<����Y��%�Fʾ�9��"O6T�Ŏ�=.�	r� �2S�����"O��B����Y��@����B�"O,x0Ýi��J�h[���]j�"O�m��@E&	~�����#~�\�8w"O:0�Ϝp��r��f��<��"O�1 o]�W&1�҆��B�����"O��Gj�4�A�ř��2���"O�1!��%��Ұ�,��e��"OD�A$�:Z��u�ˁp�4�C�"O�CE�Y�Ɍ��]�C���c�"O*p�&�Z��>�GD)�d+���3�S�)�)Tt��iV�N7�m�'h
� !�îmH�a�c�y�>�r�(O�!�dQ&B�XB$��9��l�eѢ�!�D�L��$�L�N�Ҍ����:!�D�7s��!�)�$(�i��O�C��'}ў�>9���-�z�X��U;F4�t,&D��v$V��Z��TDΣ*��.<O�"<��ɣ.��E���ļ��sF��Z�<�6�ϳu�`� BiN�p� 6�W�<au$�	 ڞ��f�P�jE��S�<�) �L������<�����Q�<�����6ZVPj���1i�V�� Ps�<�F,�'A�4�`�)��bN
t�<6-��GO��bI���#p��{�<�k.6��l�0^d����b�<�e�:6�V�ag,�=�̕IL�H�<QG[+��	�v��1���sQ+�E�<q��r��8���bV@l�FC]E�<��&B�ju�.V;O4����A�<!0C�.Uؖq��cG1��qv�zx��Ex��B�]�T�@FkZ,T�L��#�&�y2�J�_���5�	�M�ٙ`���y���!o��(!CѠj�x$q��>�yr�'HN![�A�:\~�
 HO6�y�Ȼ����	*>8�cP!��y"T:̑BV�֨;,��NC�y�ȫ<[��h$�F �x	
���=Y+O��I&��h��E��'�B���Ԗ6��B�#���ԧ�!+T= �v�@B�ɢ�`�N�6z���4,P��B�IR5�-�A?{�"P�5G�jx�B�	�=�8�Q����	��ݺV��PݠB䉹Pl�С
M�L�޼(�D�q��D>�S�O����5��s�����۟;��a��'�\[pÖ�~2"胁����z�%�	k���%�v0��9	i��垑j�jB�		���Ch��Jl�0��B��C�1l!��2�S/w%��!��_0C�	=sV�i�����R�.�3`�LC��1X!�I;�B�$;���·'Ǖu�HC�I��M��K�0iu��#
6p��D'e��Q(2.�`A��iE�����S�? ��#��֭n�b�z F�#+��!ZD"O�����Os��922JK�	l�	�V"OT��I�:��R�M YH��"Of�q��V 9��	�Q@x��U"Oޘ[��M6WH�����?v���"O���uǽ|�p8FZ�B1�%{'�'��$�=l<�%$��vH�sqbJ%Y�ў�����M����3��yq�ĳW2DC�I0�pk�d�%6�E2��V�B�	�-������L�$oh�2��L�p��B�u�~p�"!�7�T���Xc�bB䉮Okd�a��Ǐ�z��wo�r�d�O��"~��OQ+(LҩР\>�>�b�G+��>I�O�9�V_<.���0�[���E���	l�Ov��"��L/A�`�L��	�'7�l�C�ޜ<�Xȋ@G�"?��`�	�'�^-PW"��,��7K� 8��z	�'<�5+��]I��A�h�1"��ȳ�'����
�t2L���&ЦH00�'�P��Bc��1��1	 *�c	ĥbM>9�����t���R��N�|���t&�y��$��?�����^�b+R������^�bB=��"O�Ij֋�j���R��{ʩ��"O��X��V�J��A�;
 �"O�e[#�L.��!;0��*�6]�"O�I�'ǻa|(���(�g���i"O�-�tI4G�-���&�6l�s���O0�}��N)�LR��6��߮{n�G{��Og>�EM��'�Xg���P�'u(t��jڸ	���ψ[)���'{F�c�Z@T����X�S�0`
�'<^�`�*�H�A�[�J_���']�����SD�@a+�V�d]�
�'�B��*%� ��7X%N��[���'�?Q��-��5���G��	p��S#V�<q@͠8rb�e͘ 7,kІBG�<1O9�nE��*�����.^�<Y�$� Z9�|+!�H�'[�EÂ��Y�<yA��:�t�rȘ�Xm�h�Ԁ�{��0=!g�A(/�\a����(),p���s�<��� 2�8��&G�]�h`�q�<�D>@�X� J	_f:���$Qu�<�P��:TR���7��+&	vd{0�Z�<��V�E2,8ۇ�$\Z��6��T�<��k?(�|+�o�W2��7�@T�<��i�=Ĵ�@�=��@A��Q��0=#K[o�����j�V�%�T˖U�<Ɇœ�d�����!F�mf�-�D#ZT�<n	�]�+��}�~ ���t�<�p���c�^�
Q�<��4�BX�<I��{�P��'���hu�U�<1�͘�=*�uA�ϱ)+�]h�A�G�<�l�k��d����19��a� (�G��0=i����Ԇ�`c�AOL��S!�\�<���kޒ8��/��v�s���Ux�P�'��ej�+F5�ă <GN=*
�'B�(�B0��ɹ�f\�0hhș	�'A�h���4N=����2���'��i󧟟m����ƨ^Y�h{�'v�!��'�� V
��,9J>�-O��$��(R� g�ŷ��0��H�=!��,Ιk���= ��%��k�џpD�t(4���h�(Z�r���*���y"H9a����/��V�|���/<�y
� "���P��MIԋ�u���""OP�V��/9��3,��g\�S�'U���"ڜ�6*	|pQᅔ�2h⟌F{J?= !AW�,�~,�0*�8YY�c�0D���L�$$�qW&����Wg*D��P�n�*��(�u�1�⑫TB(T�PY�JY���B�l�Z�
�"O<�£�)1?B��Ah����z�"Ox�����V �� *Tq E�"OD�d��(e���O��/�^�r@U�8��	F�V,�1��7���@A⛬m��C�Il6�Up�ͤ+T@{b�.8��B�%�u��/�T�Z����*��C�	�5�*��NY�� IMvC�ɵ^�:P���Q S�����W�C��uƚQ�Aɘ�h�b�[����%��B�� 2�����0um��r�5�D-���͚��aq@�I��� k0D�T�&�M�	(��G�Y/��aA�<a����'��@�'��L�H���'ȶo>�A@4D���@lǴm0���ρ�a� �ԅ-D��*w�UUT޼{A��3i𜙩u�)D�hA�o����CQM��,:� 
3.#4��c�F��zQ|�8�nM�&�	�O���'h2T��g�Yxz�c/\:Q�l1�o��pW,��uu�|���	9�V� ���4�	R�����,*���@��ٺ�'�-!0��s�4D��AĐ� ��!���C215n�R0j1D��ڑ.��YS��򅕁^VV��e/D�0�U��a�tm$ ӃI���1��.D�x"Ui�O�ؔ�7\�d�v��<�)O �O��K~���"��=��*�$�j����?Q�'�b1
0��q��E�-�3�x�C���hO?x��_=��@j�I2z�aSmHly��'C8@��(�7G:|�$�	4ȵ��'KF�����-X ��� .�Ь�	�'񂨡@,�4Y츍�pL6s�@���'f�y��]1�hrH�/�谸Ѧ%�O��	;Yl�����& � �P�_<�d�O��0=��D�	%"�DHP*�b
�!"��Gx����f�ɟ{9�ӓM��֤��{��p��ex���	�fI0�T���gN
B׈B>`����r<���'���G�T�>��p�qlRF�<�r&̼9xj�P����PP���B�<Iv,Z7#k}���!�X���[���G{�OD�O`�3�aZ� ��*e��L9��`���O~�D�OP���7lp����F>p�V����D�zm�{"󄜽5�✠�)��-�` h��?P��2O-�3h)?f1���N0���H��'�!�$�RF�����+�ؽ��셽QG!��Y�n�A'A#6�0h.׷M/!�>7�B�[u�]&��٠�ّ;��{��_!_�d����
(�؅y�cНu!��G,T5�<�!*@1'LF�Yp��V��y��	�B� $��
�&h��T>{�C��7FƮr�&?le��!g��{���I~<�C��87ڱ��&��3kTbŊ�x�<G�XI̬
���S?�ԙq�Hp�<�gbW���cԠ�)B��a����q�<QT-�,w��i��ߍ)ծ�c�)�H�<��O�
Mi*���D�?`��ab�A�<�$�P#P@S�i-���� �A��lD{��)�65!vp�G�Ȼ0^���-?�C�I�,��X��X�J�p<I��+
�C�)� �$�"�L�z�d�5B�)z�}��"O0b!eA�(' �r4���Hg6`��"O�<���Üw�
��Dc�`��C�"O�����zOj�9%���au�p�AOH\SpED���tJ����;z05�`��O���=O>����ƤL��:0KZ�*��DX"O�)a�D�Y��2��Ӯf�D�1�"O�S�L6~���"%G[ti.\@�"O*��a`I�:����ȟ�OZN�y��'-ў�Sj�'�3TnΞQ`x(�Bh���
�'�����r�&:����"���	���y��(Y����p̛�44��kD��?����'v�$t撿F��!���
.ƴP�'m�0�[~��,Y&� 伥��'���q$Q�s�P=8!�Z�e���'��8�0#�&-����0��P�"h����|��'81OXy���8y��r���ة�"O�]곪��w��s�oœul�h'"OޡC�f�1d����Ht�a2"O�y`�-�Zf a��1U�dc�"OђϜ�3�.�B#49� ٵ"O���ͬj���]�
�h�v"O���i+@wx��% Ik�"O��;��+s�֕� ����i�"O����3F	R�$Ճ�T�"O�p�o˝b�0Ű��*��x�"O�]@2o����|���A?�4l{"O�$9%((;"X��Bi��[���w"OR���H1�T��Ú?ϒ)�
�'?��s��-W)x��@l�a�<eq��?�������i���:f��Ö�Ƀy+J�OB�=�}����!hR�k�"��a|�@�c�F�<y���0�v�y�H�
?B���+�X�<A5D�x�n���_S:L���S�<��l��h� �!K��䈪"��O�<)5$�!n�ѳD�Yox��TL�<٣��b��sOTVN�y��_Qy��)�'R���SٯfndD��R����ȓ!��3��Z��H3e,��!��`�ȓ(��j�aW:�"��ӷm���?Q���~�vϗ?^:���*f�>9{��V�<!����N�$\��IH�.%L(���O�<!��u���:��7���R�Q�<���n�^�[7�]-&�¤�2DCyb�'l-Y���i���D�P�4���R�'�JR"C�3] d�1��R�,�$����hO?)Y�1�ؕz�@
;4U)�z�<�d��tȐ+W-ZL` �a�<�T�:ÚyW
]�q�@GO�Y�<���J+~�yX $Ӌ]�ru��'�m�<Ԡ/y\�!�Nǣh(Di�	�g�<�$+�!d�*��6ϑ	U|f�ؖeHg�<!t�NO^ �	�h�
�N|9�'�N�<9h�,3�^���.�>�y�4/QJ�<��oN� t�Գ5����
�O�<!���.��QZ���0A03��TB�<17,Å$�E��R�]��y
&�[e�<i���9?���Qf�/L~Hr�B�a�<�SD[$�.=�	��F;�l �/Rd�<y嫞�\�����ڨ����F!�$Բ]��ݱ��Hk��e:GL̛Dџ�G�t��'�������Jc����X��y�J��4�b�/�$x>D�!,B��y��X@e�G)M@�p��FF�'�y
� ֝(�֍����b��>v� p�"O�x#����y��ע{��x@"O��[W��49����"�& ��i��"O|����I8e
J8S�O+x�������O��}�'!�5SG��#+V��S��1��`��'ӌH07��^)��8J_�H���'R�Ĳ�
ثh�T�ƅ��=\�q��'�f�iwj�<z��SE�G �բ�'ٖ��"�A;�����ǝ�*�����<��yr�Y:#�㑊,F��}�OӀ�y2M�h<���oX�9zy�&l�%�hO���.o�n���oGYN!5��6U!�d�"�Z� ,� X�;�*�'k!�ċ ?:���m�:��E a��3hR!�$W0z��GP}���q��R�y2!�^�)�聂SY5[-��!��O�v0!���~ع�흷$�q�/J*�!�$� P���hB�ڔ���1$O_{�ў���	�e�r\����L�X�`f�9{��B�I BI��rNV��ac��[�L�B䉗lܕ��<6=�����B�I�3��Uԏ_M�0k��-4���13f �pC�+n��:c-��|<x�ȓ|���LX"c{F,�&��p#&͆ȓf�֘2&#���t22�ϳa��؇ȓ:T�QuI:�츤I\
\q�x��%��̐���
���Î#���ȓZ�8���V�'צ���X_���Y�Z�#�&D���\�&��Da�d�ȓ7�* r�/�*r���b� �`E��1Ð<qM�@Np��T�g�ͅ�!}�-+V��K!d�*�֌�ȓ"�6����  2u#��v�P���v�dp�3LI�I�X�ꑫڞ*�PA��wJ�����!V9��0��R�����ȓ%�������TY�G&K�
R-"ړ�0<�&&ֺ,/�͹w(]�
��xpg�C�<A0M�p�N�kP� ;�t�%�UB�<aW�[�R�"��2��:�D�B��}�<��JؖT�.(�ţ��D!0�gd�<�e����&�|{��-_`�<!�)U�[(��y𪇈1�n�ۗ,�e�<s�}44*pDZN������[�<�FM�	�(I�F��-W(��d�P�<q��Q�t.�Q�g�+krL���_r�<�ˉ�Vh�!D�, ���l�l���0=!� ��8@"ѵdSj�К� f�<�aN�l���B
Y�2ׯ�k�<)��^$b���ˁfnrБ�j�<��jΪ���������cD`�<I�"��8!����Q֊�@�<��H0]S�ݓ�.Mgd,X��B�<I7Dٞ::�<�t,��0�9���FU�<I���0fz�82��Ձ�6��H�O�<	go�j���RCͼH .uZ£�r�<Y�A<(-�\�Gȷ&q�mz���h�<)�1+��$h���2]�XM�n�I�<1H�
���B��K�K�<Q���(��lC#���.}�d�q.�L�<�uE !�X�ґи�H;�͓ry���o�'_8J���e7�-H�h��Y��)�'�����Lpk�H���%��c�'��i�g"K)耩ю�$d@Q�'������*`"5���[v�K��� �4@Ä7.�$Ցtm�&A`"O�Q���{vd* ⚒Lβ$��'�T0C*�$�`/R�^�U�v<%��)�'��q0b���  d��fg�a�j��'�jÙ�U��m�6NЅ(M���	�'�������#3 ���؄KL ��!"OR�S����(\�za��A�v`���1LOr�ʂH[���3�NΑyL���"O���C��Mk:�е��$o���"OΥ�B/��T`����АOSD$���I~�8� ���n�Nh��+�h ��o=D���p��_� 
��*�, �s�%D����0p�F�s!�*:Q � Vh6D�ȫ&.Ô{�����R���v 9D����B�Z
􈩠��DT� �G7D��*�� U�|j��R"�yp#7ړ�0|Jկ�/�Tm��^�}���
�ǃf�<!��-/�
�Y��G<#�\`aV�m�<I#�!Dv
!I��H���:�B�o�<���ѿJ�Z4��&5,d6�7�Aj�<A�/�x^���á�(C�cc
�c�<�Ӄ�<�!1�"ʚ�kǅ�y�<�!k��@�p�埛=�J�c���w�<��FĀ1�~d��ހ(:��@�r���Γ!��mb�ꕏY��D�"�3�ج�ȓ=U�(��O H����M-nXQ�ȓ~H�-���+``2)�'#d(��ȓM��x��� �h,�f�
�}��4�ȓ]��G�|�`|#Ō]�+P �ȓ_	.l1r�Ҵx�S� �Y� �������gJ�I<��"�՘A� (�ȓa���XP��Cw)J*AJq��?��Y%]!�:u�!{[ (��_ ��bf �?.��59׉%�)�ȓO���1m��f���Xv�E>B�lI��o \�Qԇ�@ Y��n�N�	��B��0�&�"5�Va�b�>J��H���pȉ��0���[g���`e��g(��8��;���!�Z�$�C�I$���҄o��`+�ř���&MfC�ɺ	bA����f�6�ش�I�7*C�ɉ]vv�8���
c߾-;��]�n.�B��Z#��� CD�*G�Q�]�.W�C��xJl�t�e�r<�L�3�"O�`	�C�B�f��[�8�ز"O��z%ظ��ݻ��	|b�qc"Or\�$�z�)�BO[�dy���v"O��k%�O]p�̑��Ƚ	�I�"O�8i�	F =�P&�5	�r��"O����j&j��m��+O��H���"O@m�&����ݠ�+�=g�p2�"O��3F`8	�LBŉ�2b� ��"OJ$;�����rFB̾n�ܨs�"O̵�Ҍ: ����a�,#}�pw"O��H�a�@��IFbM)�"O�,�cS$%��E�u��<;�1�5"O���We�/�r-�����'CF0�6"O���6�:��J�v�i[v"O�e*G��6DS�H�K�����"OT�X��7��%�'Y�z"O�m ��(i~��S��sX���"ORqI�*�F�Z�95��'%��6"Oԍ�E�Lc�����`t�e��"Or�@Q�"l(�#��g ����� �E1R��!�����<�јS"O�0����FjM���?f�4m)"O�����:Bni��aE��$��k�<b�.2"깱ա_6K32h��p�<�A�	�su�<Y� X� �DD�Љ�o�<YΙ���8˖JŦ ����e��l�<ye��Y�*V��"~Tf���ml�<Y!ĂZvјŅU�N����bA�h�<�)O>zWr S3̓�\H*� �oYh�<1�-�>�
�sŎ�67@�h�mOK�<)�"�Y�b��X5e��@(�O�q�<�3��E��`��FE"i����`+D�PӰ�� 0���B�Gʊ��F�)D��zAE��/Ă)R���x�
T=D�p�&��7����p�6;N<Hp&�<D���M�N���3GIY�F=����';D�h�A�rN�\#�&��t���+D�0���K8lخM��?4G2�0��(D�t e�
�F�)$����Fّ@e&D�����.'e�`����+����/D���l�
��8s�o��R� 9�"M:D�\(���c�TH��.�(wy�T#�b,D�P���U
�� ŀ@ ��(D�����]�J?b��gF���:�RgG#D�P�`�S(nTP�)t2V9�R(4D��Ӏ�G�B.4cϟ����ũ2D�܀4��=IV*i�C �7s�5���.D��3Ę�a��ad/[7"�=˧F7D���M�r��3%��QY�&2D�<k��@t$�f��0���S),D�D����4: ����O]�^�@�	/D�l�V��w�&Yj'�
{2$̀��9D��Y��,Z��m�󠇱V �R��2D���c­t�������%��0D�p%P�:��)f	�fD���f/D���cA5$�j�)�Ƕz&�5zb�2D�Hz��D����AX9:킕��"D�����ϲt�$\��J�.y��1��#;D�(FQ�6d�3�Æ<�'#�Z�<i�&�PP��Ɯ5:�Ե2V-�[x�pGx2⃂ �VԘbOcc0iJ��yrjkT�d�D�E��h�&�+�y"��$���X&b�Q̪�ʅ4�y�CN�3.|Ĩ�)(Kd�<�"%�yN�/U6�P��H�/�� Z#�.�y���bsءۤ���%���P�̊�y��6	^+U,  �����9��x� |W����W�-�X{�	Ɓb!�E�>�F�A*]4I|��B�D�U}!�d��dT:4��r<v(�
sy!�$^�u�l���^���I�x!�d^�*����2�A��EQ�H�&"!��I�~.U�H�cd�l����2�!��2]�d<*�bY.nR0�X��T�!���`_P}J�D��B����E�%�!��<VG� ��ֶ��L�'�V�;*!���	&�$3q�[�%0��"�bޘ!�$Q�%�j�t&�<>.���O֖1!�ă�i �H��g�'%R�7�N��!���8%����� .�:p)��E�I�!�$�X^@�1�C<s��p�(ٞ^�!��])��<K��z���aAݟ�!�D�&��1�NG��priT��!�ˑ`
�<3Ro
����Y��ـ7s!�� 1&C G��x �)��8��F"O�I��!�2F*LP��|��A"O��aj<��R�
M���(Z"Oƭ�r�"�*�h��M�^i��"O�,�2��c�h�\�^͌���"O􁺶c�PJ����T�xq� "O"X�6�Cָ�Pc��Ҡ�!"Op��1CVe�2BV"@_��y�"O�p��X0��#ab	=IS�K�"O�ab-������M<��k"OF���8{�9��Ϫ(�Ш�"O���N�4 d���pB��%�p�#"OdH��`2���#k@�a�R�˅�'�!���%9�4I���`���1��ٳhg!�D�'2��	b+�!x�PH�"A2\!�d^@��RB�L�5�,���!أ[^!�dC�x�vD��_�u����UDL/!���<�l�v�Oa�^�a@� e!�d�e�B����?���!�I�D*!�dץ3
�H�ŉ0Z\qj�ř�9!�dS@���a�xl|�J�Ø$@�!�$+&�B\�M?�`��q(�;A�!�d;�>)�O�v��$b�ݲ �!򤏾���
x#`��o^�u�*�B�'��Hy�A�]����R��=滋{�'���U�X�aΟ3M���'�(H��B���+��P�_N0��'H���m�%4E��P�T(*l��'��}���ɴwV��@GҸQD~�j�',̙Z��ǵ)��m	Ă͡^��)��'��a�#(O�\�#�8^�N,{
�'7��뉗M�hY�A	:G�&��'�ڍa�(0Z�A�2O�)/R53�'c&eq%k=xd^|���J+�A�'�<q�� /"s�%�(�O�%��'T�PQ"�N4$I�X[�f��Ĩx�',�IE�
~ȲuH��[�V)�'��2%)�Q�d���9��Q�'������*"x��O�y�*O���!/�T ����ɤ\�X0�'z*1���6�6YCGf��JP�pB
�'1�E����F'��y��֟KJ���	�'Z�����h�	��4Gp�,�	�'������� |�$��E�� D��Y�'���Q�����j�LX&Z�t�'�&�HT�X�2t,�WKߋ|U���[A���G��I��T�Պx�89�ȓ-�J�G�p�@Yf)@P�Y�ȓcQ@������H�@[\�i��Dm�� ���mqW��<>��(��
#�gb�a� �61�C�	��p����
���֌Z	D<B�6|��)Rf  S����&*�b�JC�ɕu�M�����S�*��tjU�u 8C�ɳz0N0���$Q��Z7�0+�C��=;z���L��"ӥ]�f}�C�	7j/��11��`K^��⧝�&�B���%j�B���c#�	��C�	!C�`U�d,X%D�e
n���C�	9������7ɸYd �3
C䉢)�N�P ���{�Ɉ�� �U�0B��&U��E3�G�JL�t.�A2!�D	�tx&I�`�\�vW�
�!�D+IW
���G�C������C�H�!�� ����
ѩ9�F<�2G44���"O 1�7���4\�
�%�����"O|-h�EۥC��L��㐧+��0��"O�
��О<ڼz�L2���"O�l���l���Y�L�e�����*Ol1 %ŪR'L#s�A,SzF��'��8�"��
 �Q!I*B��A��'"(q���S�Z >$A҂�8*x�J�'��H��N�8�J���+({f���'��mK�N >d�����ğL ��'⊉����� ���A����'dVpK��@�
�Ԓw�;��Q��'kF\C���5C�8(
��-� �'b6�ڰꑲj��Eb���y=���'�X���>d�Hj�g�5x%�܋�'�
,�Fʎ�z=��dôi�p�B�'�,[��]�TnBl�dIWx���'5���T�p���!פ�B���'x���ۇM$j ;�õR<�b�'�^lB��=w��cmыO��T�
�'n������ g���*LSD
�'�(0Zd�I��¡���ZO>��9�'*���Ȩ$�����_�H�%X�';Z(c�E),�F])�FA�2b|�i�'�|����0c=д���D=}���y
�'F�� ��
���K�w�p	��'jVTYq�$P�zc��@����'5�0RR�
Yb�I�r,�=H�#�'��TS�c;
Z��B` �#����'�(���X� v���.����'-p�Q�Q��dQ��[�&�����'}���I1�	� �͉%}5��'Ϭ$�3GC�P(�b��_!�b%8�'K�%�0a&�@)2-�C�D���'!�L���Zo@a`E9^f�:�'Dx5E��"
&��MEG@�-b
�'N���jR"�*�i�5>=(��ȓ�6}c��	=�V�jPE�X����R3�� ��Pށ�&��af|��|�:i����*S��w�_�[��Ԇȓ/,��ߨLB6Db��Ѵ= (

�'H��t�x�� ��ؔ2�8D�xZ5��`�:v�\y2�����6D��A╇h�RљV��>3�$��4D��x&E�i�ء��)ȳBd�0�/D��8p�(`��Eaqg��1�hy��y®�Vqh��4�$^�Τ�����y���F��d����G�|�(��/�y��X�Y�$�5����2��7�y��̓[��-jʅ�8)�� �,��y�C�T��ZDg)7��{5ȅ>�y�f��2DC�iK2���j�J��y2��:�Yӥ�:��H�dT5�yr�=����QN�	cj����0�yR��>���H�HJ"��O�m�<A��_#w6�c��c"T 9�Rs�<��`d�l �dE �G�v�P��n�<�3��`���._�Yn�``�Ln�<�r*J�_��y�枇}F�pC�Jp�<q�_���P/� n�(
���P�<��d\�@F|���f�o����^P�<ɒ'�>�2�*�=�2�lw�<���?������X"乓"�H�<��jۨA�U!Â:*dᩓh�D�<� �-��cV��y �lq�0	�"O2��H�:F����'�ڰ'r`��"Oօ�*�N����r���3<T�"O�`�P���x��Q
h���"OԸC6c��͐�ek�;[ҝ �"Op�9�������\|¼�%CF�<!�N�mJr#f�Y�,��x���LE�<��/��#Z��;D�K(����e�<1b"p�R��$5eJ�bC�CIa�<���C4R�ЃZ�r�M#p,�f�<�q#�0>���6��"iʲ��e�b�<1���5:B�9�
K9��c�#@`�<Q�&Pi��5�'͆0�M
#TZ�<�#��%v�6L0���[H��d~�<�N^�8���Yf�u.$�ąMy�<���8O�:3@EE�EȎ�ȡKy�<�c	*hdΘ9���j�By�p��j�< JZ/JU��rD��/���j�b�h�<���� ,6l�⧤L�_�*X:H�K�<95&�|�\а�E�B����S(F�<A+�+K�
9 �M��"�ʠ���D�<�++�̪�	'FSrݹg�A�<f�^@e+� [8v�v`Q@[G�<A�/�sk�<����v6�����}�<�Lb��9E�B�f��}Y�EC�<1	���3c�4{��*�,�s�<�
ƱLO��a��qF��r Cp�<�$�E�:G����6��ڠg�R�<����'F�y�\4X���XF�P�<ɐ�A1*��HBd#�4{V��L�<a���,�h���K����L�<	�h˜a�)��I�>�"���N�<���B�I�0Z4g����w(�p!��ؼ�"p�1`�HB�CvJ��f!����NQ� � �nG�svgµ;Z!�$��` �1z��N4H���f�7�!��߼Nqt�xG�"jͤ� �CM�S�!򄈎��ق肔<�8�yP�Qs�!�$��r�r�%E�7���0�E�\�!��1�H����&�D9�AH�9�!�H�K�h\;aoس�d�{F��!t!�d)8d9s�C�Cv0-�d2\!��Q��9��yu��qw*�5>!�$=j@&`��� "B���U�åA�!�$Jw�9�e��P�� �G��!�$Ȕ?kJ��4ƂS�,��$MIA�!�D]!-n5����c����[�?q!򄇿l_
��*�.l"M�P���!�D�]l8A�Cd�sŮV�L"!��נ_��5z��'�����\�x!�DL�"��q��e�2�q��Ȅ+�!�ƕB��0u��C��|Xf�ֺ�!��GP�J}xCk�b�ި����>�!�d�(�p���hXX~~,�r�uy!���()�!a�Ou��0��'{!򤃦>�<ٚ$���R^������l!��Im'N��8P���qˎ(`d!�$_�|r�и�GʻnK�-�4�V�+&!�D_�,0x5��`�PX1 	N,F!�R�^�0�E�G�4�6R*!!�		q����� �G4�|�R��<!�٩^�0�8�LQ�1������
7�!�d�3 H��97%������h!8!�$Ѧ^p��c⟖#B d����)@.!�� �pY�`R�q�,9q4C@6;�P��"O&�@�L�#�84�)�l��"OظJ�ȎYF�k4�A	=A:�"O���d�Z�I�I2�@M� �,+G"O�P��:sgd���h4~���`�"OrrAc�4Ş\Z@H	�p�@�"O�h�A��<}b���%�7�U"E"O���H)��ȠǤuٸ8{"O�hA7��U_� ��đ*�����y��>�2�kB%����r�HΜ�y��9yH�d���(b��o��y�@A? "ҙ�4h��"�q���yF�&f3���6`޾oM�)J�&�yB �ڨ`S�K�b�޵Rì��y�J̙4�4��[4V��Ie]-�y��-V#�!�rgGD����I�yR�W�|VƄ 1���K��-z�Ə#�y.�*�Dq�!b\�G `'��.�y����,d�X�m�)��:�J��yR�G8k  Kw�޶7� ��߈o�!����U�Cc��h�`��j�!�Dђ0��Ec��֟cl�9�.�"e�!�J�D��9�"��*k4k�l+�!���"=���L�"�I?O!�$��|�\�Q���u��)�
�P�!�����!�p���2p��IP��+�!��1A3��j��FT���4#�]]!�dG�֭��C�F%G$LM!�dΩ���J�e��^�4,㲣ݔ&0!�䇈HP��� L�h��ktb�$X�!�d�.p�\�
��b��`��"�!�D����7�1��9��@Z�>n!��A�����B�W�f��S*
/>!�dű^�X`z4$��k�T5ZQ��t�!�\�!~����@MYG���g�5!�d�	�&��4`Y=_-*�S�ژ%!�d�n����4����
�� "R!��V)&:VĐ�C�b�0`X�&b!�ܢ�ڸ0��@����@��W�a�!�d�|Pb�r��]�@�~�r����PybOF�
	p�K�O�Bn��ꣅ�,�yB��J��;��
h�Z����J��yBiXI� %��ʖ�D4���I[��yR�^s2����A��4].�y2m� '�P�q�@U�S�J����5�y��W"B5jy�q��]7 ��ا�yb	ՄxN � ;Z��`��N ��yb$Ϛt�j�˧�	�.���h�
�y���<3�-v��>6�p2�é�yRZ�B�"h��O��&u�E��.�8�yr(��l���уKŤ%*�h37f�4�yr��C� m*����h`$L�$�y�ȝD�,Q�U�J�����f	�y"a�-E����:ChÃ �yB��$�ƏQ�3��8t�
8�yb��5U&�ix5		//䌄s"����yR��0q� n�� ��ƙ�yr!�\��]���'Z��寏��y�b���xA�'�ݚTyh����B�y2�_ ��= v�?��a�m��y�
Y�U����K�9ް{"���ym�M6��K�c))�R-��&+�y�L	m]�\p�V9t<Y��O���y��4Πm#f
�=w��1%�U��y
� �����P�9h~�rA�셁F"Od(ꁍ\�m,THz��ѓ4��*%"O�1C�L_:�tU��-�-"�p�"O81â�B5X�xU'�jl�r"O�X���ܩ�jA�ƥ�'�A
%"O"�u�OS�"��0y��{�!��	;<@��N�(.���l�8��y��!,���"�� ��Pd�ֽ$>�B�	pd#�Jl�	 ��R�!�����S��(S�.{q�C0h+'���=:(�R���${�jM�f�*F�ф�Y�Rp1wk�4a�<Py#���DD�ȓ6�����N�N���ؕl�d���'_R�kfE#6pz�8a�D&!R��4�hO�SG�H���X�D�[ct<�t�J�W�ȓ(�4la����Q.���!5��Gx"�)�3�S�?��S5���EHCd^D�<��Jm�`t"�(C��&'Ʃ#Q��G��'�N��J�+K�N�C��؁=�65��'8�8S4ğ�~� -��ɾ3�Xܩ
�'id��pi�(4�H�w�	�%LdB
�'�h`�Ԩ���4��fU�g��I�	�'�`,xd��.pg��#��J3�\���'Td��h�?6����F���'t�i�V# &U���8g-�!ƌ�I�'�)e-�5~��=ʖdM<Q��'���N�Ā�a
1{c����'�Eq��� #+�0�P*ñq�th��D*?a��)@3Y�P'��HN��2n��K
!�Tk!\ey�&�(eF��vj�
g�!��5GR�p`�D(�Z��QL�?X�!�D�V}�BAs�tL1��_.s�!�'$�q[)V�	}�$���"�!��
l�f R�"рt����Tʀr!�$�#D/����+
;[� ��$
�Ee!�ņi�=��M	Ep �k&Zj!�?.hM�r�F�kRz z�ѮXc!�NHTaHq`xP���JD��2O�x�%�oh5�ޡ.N��""O�|YD�6��u@��zV�(#"Oz��Dj�u`a���	0�n��3"Ox���S�:���`4�D@�X1C$�O���$

c��d� n㶱��o@-�!򤎖,�<�0'쐆s�����G_"�ўt��Ӵw�Tp���d#4i�nY��C�;�E��8G��`���֘C䉽+)�QhAn��3;H$�O�#(f$C��L�z���m�<�D,� ��M��ʓ�0?y��L l,���Ui]�QtX���NeX��Oz%�'N	������|���"O $2�-[�:�,��Q;�,HB�^>u 4J�l�@D�s��7Z}�aL%T��r1�H�u�"�!3�;&�2,��<O�㞐��I�~W.y3%ŗcC>�s��۰�R���1�$�0�8�PA��)8 �UJ�
��f
Ob�{W�ѷ�t��T�֢0��M���n~"�'01��8YqO	X�X��܈:�:����':���z��=��H���p��Rdr"<����?U�#! ��鲲E�$��1�F'�L$��d��*-�.���)�uKx���c�>Y8�Gxb�'��l���&/�DJ�(@0I�����'y�"=E��+�HT��D.�� (�P$�R��y�`3Z��if��Kz�\�^�nM���@�f�<�~������T[��#{� �o�r���֧� �m�ԭW�V
Ir*�CM�i�"O��X���<5���h3^t�P�'�9�'�R,��/J$>���+šE�z��}2�'`Vͳ%��?.��\��#2ǘ��&�S�T
U:%������=g��	IR���y��+/�$�K
��luLt"U�I���<����OHK0j�gf��B�[e��`4�'�d�.�����U�r�l��9�0?���Ŕ�T<kV;{Ü���l�'C�����'iiNX���)q�Q�Q��&L��z�L��&9O�<;Ԍ�H�P�Dyb;O�#~�Q�&H���J���KWi�	�#�y�c�;n���c��,ԨI��拚�?�*O<�Iɦ=�O��I[y�
MP��-|s<]�0�K{l�|r�x��z5�ħN�)�Fe+�A���HOX��$Ѣ_�zxhcg�R<t\�3T<'9���$0��IFd`���&\�1d�5*@!��S��a�C�
�
܀����_=�	S}2�'�L���m�:��nS�}D��	�'��X�5�L7<�*E�D���y�e1	��Q=?����K`j�5K3x
!��[�Ee��9>���!땶4��'���H����˖"p�&N�R�����m7!��Ң5�x���AήG�v��A_!�Ă�l�\�Sc� !���D�X�t!�D�ed̜�'��X�:DؔfJ��!�ϫc�R$$\�zn�`9�
�c�Q�8G�tg�?9E,��O� �	���M��y2�ڥ�0\1��.
f\Q����yB.T#Ar7$6Ec�b�>�-�
�'v�F$�#}O*�I���62��1��'o�!U�G#q�[���`����'�@�Z��.���Ԅ�<f��1�"O��!g
)R��� �ڳP4A��'�Q�lh '��?�|8W�Ҋl�4!�	"D� ���ã;� I@VН|)2�"-�D�S���OT��1�Ư ~:!���70����'�6�T`��������z>5[�'n��@!�%J�5�5��=���Uh<Ym#`���S�ӛN��4zjB䉙b�R-�<L���Q�'7����?�I�"�aS���b���a���5q 2B�I%~X!�Q&�>`�'��d�pB�9��,��-�(ٴ��GS�=��B�03�f�A(�QmN}��.��B�ɓϖy��� &�N]�5FO'.�B�ɀ&�
��!�<\�09c���H�B�I qA�E��I��}&!Q��!x�B�ɱ��)����8D�k�GB��B�	�Rh�IQ�K��\�x�R��GC�t��p�����Dh��ǙS�B��̂O;2XIG"OTu�����  $�KUKE<+z
u��������(x�a�>��ku��$"�B�	?zW^srÛ~���[r�V �4B�ɢ��ٱw�׾qK��S�)�NB�I|<1U���Z��8��D7���m#kݝBm�U���!\���'�ў"}���Q1�~� q-�Z����S$�i��Ԕ'�Z����Y�~���i���03ДD��'�ʕF
O��5D�0pެ(	�'��t���tC.�9%f�>R�^�q	�'�C�!צ��JS��?�
����5<OXh
��ԍ%�lH��:ZwEj�"O�aRT�W����s
E?U��ˆ��$\O� X���a��E��}�Q�/z*�)�O�`8�ϭ1#�P��m��5��#~�<�իU�.Vlkp���.��S�I@�<9�&M1yĺ�s&��8]ݠ}A���d�<Q�AȦ~,�\�5J�O���6	��<y+O��d�<�|�'������F�7�9#��O�n��Y�	�'�&]��5.]�Kŀ�^@�Pc�Of��$�nL�+���lC.h�'�W�x!�L�	,�R2�̓=T�@p%�R�b�!��>&��q0�L/0� �bY��!�$�!$*�嚷��I�E�g��3�!���.�Z	�"��O�H��!�<l�!�$bиŨ��ʍ$�~��g�4!�$����
�A9�����q�!��G9b,l��%eӈO܀JEAɃa�!�Č�=i�у���^ �=�UA�	�!�'l���r$�	9w� �6��
u�!�42��X���/\�L!d��!�dU�v��8QH�F�Xu�b��,�!�d�'x-��"D�oۘ(�M���!�$�5r&̐�ܥ=o6	��k��/!�d_�h��BP�G�L�����1!���kԐĉ��хt۾��$J�*>2!�$��HG��b�n�	҈�Q��.j�!�Ą�u����%�.	�� ���F
P!��ڐ5�p��N^�a���XfLĂ/9!��8qf��!1C2Q��\�F*!��șQ(�l1�ꡣ @!��\�s�xف�W'�h����$!�$ˀq���BS'f<qc GH�2!��+}�l���6Z�Z�� ��>�!�%��M����(<�2��6ɋ��!�$D6D�%E喞qe��+G(��F�!��7H�z��?r�1��g��X�!�D�`3V;"�£�P`#F�m!��Ď`Fđ���B�h@Pӏ��p\!�تxy"�X1D;Q�Д����(7q!��e���&�6=�I!�t�!�dʲ�`t�D��7�X��-ʨ{!�DL�d�LT��H <n�Ȱ{0N�?	!�%t�&0Cu���
D�!��έ0�R]��C��O�*�[��H�@�!�D�~�<)2&牳��X8$M3�!�d/&�XMK�˔�.+Ɂ0I<[�ȓh|�ZE�-t8��(�@��R) ��?�b�AcA�pY�GD�23p��<�P��05<n���ɇ;����Vv�Q�$D�QÂ�|�2���@�1-uP̅�;nI2� �8\���i�$�6`�ȓ@�M���X�d�^Y�%GU7�x(�ȓK ڸ����F���E���N�����w��aTK����5��n��*m�ȓ2<+U���nG���gmΐmX`�ȓ5�p�#�!&�h�	QB�)K���ȓ#�.Y�NݖC���@�!C�H�������$�)���@�7���M�\�8��J'29܄fN\�N*�e��G�ԩ�f�"�z��G�8���;}nL�0E������$<U�ȓP�,l0�&�5d���r��w$N�ȓd�J�1`�N�tb�p%-8�L��ȓg�Z�g�1�� @)�OO者ȓ!�͚�O�4��'S�5�f��ȓw�(TCW�"�4Pb��`�� ��t�^�A��0�8��K�9����S�? ���e��AX1 �)�2��P�"Ox̪&) 9�`4�e'��!�$ AV"O��b/'4�D��"%���G"O��	H&+3p��V��s�Jze"OZ)�I6(�j]�� ҥ
y��I�"O"�� ^:~^@��H��#mB)""Ol��Ԃ�.0�Q�EN�7Y6x�"O�y���	�{�t��w��=|�lX��"O4�-�&��P`�B�6��d��"OB�yw������@�:0_|L`q"O
=�O^?6?|�IF�C24ܱzc"O���t��0�0(��8RE�)W"O�@�dCSf�^�@7)�Q?�$A�"Ot́������)�� 0=
(*&"O�i�kJ�i���y�Q�1$��
�"O�8�G/�\{�ܨy�3�"OH�7�ȇ4���.Ө	�l�g"OV8 �A��X%�D
fn">�@� A"O\)B�ܡ$w�ATjҼ��S "O�YBC�v.�q��,����$�5"O\,��X�i������;Y�3d"O��hìݐo�9ô&St"Oc�B-d�T�CU` �w=�,xD"O,���Գ2,�qK3n\�t�n���"Ol�є�x8S�ݝ�� "2"O(���͘�m�h��BK�<��ݒ%"O���C(yS�����Ik����"O�� ��ّdT�A1��ۻQI�,�U"Ohܲ�L��+`��Q�\6xkBD3P"O ��_��И��H5GI�59"Ov��UA�~�b<K�f �q�R$��"Oh�X�F�)�ᥦ��&��B"O�mY��ژ&j�)䄹A�@�"O<+@��3Z����r\�`(�"O��`ㅐ�%�>�Q���$`T�1"O��c�
ͬ [���I��8j&"O�E�Ø�=/��S5(����9&"O�A�2Ŋ&{���u�P=hw�A"O�|�`H�L����PS<-��"O��(h��V��ɹg�S
Z,\�0"O:���-�66Xf���ȍ~�H3"O�a�rI8`zT@�`%��|�jQ"O�9+�Ǝ9�pC6mS?f�����C�d䐋{��9O~�C�O@L� "�-TL�z(��'&��R��>�����,ldi۔e���mFҟD�i��C��I��I�~*��6W�Zʀ���ңA�z���0	�m?�'˄��i���'��)b��ۜ*)��	�f��E(��'U�V&X��=a���xp*��6�vO
�P�U�/o��Ҍ����ļ����(q����ȗ�N��q*�m�<��Q'��F��ˇ��)��c�P���O���D�џ�A'>�Gg���&�g}�t"�0{/����(��0��K}��4g�J��;tF\p���=�M����Gf䩺'�.|O؁�����1�D�2��8��do`�NT~yB��)i��!t���?�qV�]u�FM�&�ý$-J�;o;D���J/­+TG�:M�PѺ1�V�B��Y�r �>y�J����)reO*操��ܱQ4���*��3	��!�,<LlXb�J�iQ�FF�f�����$"l��t[�0�T%��p��3H����De�F�P�0�k��џ<�"��`��CM�8�D`�'�d%+s��?�9��
��t�	�3������_�p�f��
��L�1���IJ]�r�>���Z;1�Dz�Kd�Y�G�?����P�-6��|*Դ����<<rႆY� !���k�R` šL�L�8e�~�����jćRΈ� @� Wڵ�7�~3 (�ēt�.L�6�<L��q����.�J��	�P��A\~��mY7��	n���`��'o��m��_�p9���Ə�8Fy��S�? ��1�-	��8�S�l�X��8��ɚaچ ��Β�7�ꑸ�R�̹	���AJv��%^�>��|(��K?~�5
�O�p22)����)�m2���d�O�]qGe��IK�|�A�q�(�K�qVrT���*Q�-WHm� ��(���O��y�-��W�6Ě�1!�nԛ�����s�L�-
3�4K2��n��	�Xw�X!�0��+�nG���$����`X�Z1J�3%��%,�zr��F�F	��tJ,;'JS�^$�����#��,{�H��w�<��D�	��X�Ggx��D,X�8��Oʒrv�$ �fNqO�B�I��&*bɪ���,{T����OB�%��7q�fy�Ƹ0��9F��GB�@��w<a���!��!��ьK���W@ɰqV	n 5�$�1i Ӧ7�� 1��@l�!���y��R#�S�AJҜ%���e6������{�
��R�|��HXn2:���>R���u.ǀy����Lyb�H�?���M~2��銷��Xe�K��L�F"�`���C��|s����umO#u(h�v�]�Q>8 ��#�Ď�f�vd`2*O��!�/'���3cZ0 6�Ė ����(5{L��㩉��ճ�D�R��St��.>�!�d�I�2���iO��RӬ�!���_2�2 ���5=���@x�!��I�l�������38�b�) n�x�ȓ55`���':S�arI�A��ȓX["L�2��	���A�cr�ȓ_<�T��	:�U�vD�)=�H����^Ԙ� ��-���R�	+{�$���R���Z���'nfx��E�%l#�<�ȓ'D��SBM(NybUkBJ��X�b-��J+��F�����\kŇ]�ND���dA�lT��9u��x��A	 ~���u�)�ŀP�,#�$+&@��K� �ȓ=�
9�re����� 
bQ�ȓKӛԂ�ZO��J�V�.�P�'��x�֠֟N4����@
�	2���t`��,)Vԙ1ի�!{s(�#\��IS"O~��7*���];�HQ)m~n]�Z��C7M�G���%��|*7j߽O"�Q(S&����A	gX�@ �&6M�'7́��&��<��'�.5)��c�>q`oϟ^m\�����}�E�}���@b�`�!��"���� ���[��Ť��)��\�,���S��e�J2Ȓ�X�%�`(��@��G����i��u_HǬUC�&�`$l��~R� �g��bv�g�-�A��E窈 �>�1b��Li�cH68>�p���%�����I�%���beL�C�P��QE��m	�b�b�$��t��S>t�f�O�E/��'9�`���4%-$
�2V�F�� ���,�1��O��b� P/`�f�H�� ��@�l�~=rD��7�<E۴��|�"��N�p��)8z��Y�O|�>��I�2�jex�n��bH�Q�F���<)S�VE쨨j�h�"X��i1��kq*��ƶB
�b�^M�0� ԪŹ"pt$�'��1'�%:pqS�Qe�T�1�ț�s�FT����5���
��u��9�b|��%�|��ƀ�k1�>B�p��9n�a�'j��X<>�C�D�o%����Z(H�k�ҍ=�^��&�XB<JL���|2�X�@91��[�ՔsɊ��FL�S��#P�	�F�$"����$1�=SC� (�Χg�1��e��G}P�z�
�x�@�<q�J��y�B��$B7�U��Չ&|����+H�bc^4yH�0�`�.8]h��t�B�6�>݈P�^�}��$Y"n�= J���	Hm�<i��X�sc�(;p$��,�s6 ���wf�2C�Ka�:`��O����-@X�,ӧ��NAб���)�Oҽ��I�^�
�
v�W�n�,�i���#6��}®�g:`y�&,Ҝ˘��dR1#G2DsS�L��t	AN �ў��lH���8!���$4TR�{�f��|�QI��I1��S�DT&�N8�2�H}�<�����%!A�g#s�G���l�hޓܚ�)�⑲Ctڑ��D�V�OZL���&�Չ��Ӻ
�R(� "O��!F�P��A�阝$�z�X���aa)�Qlޤ}���	"��00�3�4��#�K-|2	�T@���	*!�~������?펍i��G&C֮XBf�̽�t��S��u�th"t�'A��H��%��Q���5 ]Ë��_�Vxl��n7-�
Lz!�~J�i4b	�'NE:4��	ҍZS�<)ԯ�Z�J��)�a��hc��k?!v*�K8[E��yZ��'�"Lڰ�� ����j$t�@9�N�_j���"O* "���u��P�]0O��J#� CѪ��Y�x��t���1�O��3F��Cy�H�]/�u*��`ح8�"����?ٳMȘ[T�}!� S~YgiRHm `��E]�1Ԕ�u�,M��性X�#?9�	�bw�ui�E��7f�Y�D�Sw�'^���w�a֐��oCp�b�^$�`�J� dY�ᡓ�/�����/��Q2a���K�d��� :*�������$�.�TxSޒ�~B�_�[Wf%7�CX�S��l|)E��nJbD�3e���C�	��*भT�V�jVN�uB�u�Uo���⢊�>�z�C��m�Ӎ9�n�k�]�X���_�H4�Bs`;O.�9;�6�OdM�0
��(�Τ)mEy$Ҹ��NågW�"��~�f]�s6�@HW�'5X(�"��{�<�K�����X��D��]*���$���~�.�
aZ��YGD�w`�
�C�+3y�ȸ2�ɟqB��ɁjШ!ڑ �A�F�Y����ʓlF�#���.5�H�I5E>|Bh��<*�OC�X�`�' ��AN�|\��c
�'Cb@RR�*-h <����,kYܜ3$T����ޟ%��uY3�0�'��q�'�L��1��� �vl@�k�i��'�D�(�d�!g��}�P�S�,[����CJ"�O�ԛ�O���0<Q�)ۘN���P�G�|jVa�Se�Y�<�c�R(Ny�0N@N3� A`�Z�<92��O�x���bH�0�V��V�<14H�	Wѐg�.�JLD�L�<� �#ތ�xao�	+�͂'�S�<�����&��A*�(P�����!�p�<)�Oͨj$���[�b���g��s�<`�G�R�v������<����v��t�<��)��)��a�+D�޴�Y�<!�@�T�#�L�"A1^e`!�T�<��E1B�%p����x��
y�<��!X�h'�4�a�S��24����u�<a�h��a��I��l�&�HPa���Z�<��>sG����ǉ���9a�
VQ�<�G#�.5|jt�P$�0&D��� �S�<)��Ԃ1��ɻ#"�J0n�ks��N�<�!@�:�hE���O����OED�<�S`�	aL��GI�_R
f�@�<9�o�%Pv��1s�N�9���fʇh�<�� �>D(H(�&ӠOc�ɳ%~�<��b�=H����j�d\�E�y�<��E�-G����5'c�x���r�<i6��[��Pp�/��Q��L��+�k�<� *�9=-�=�u����b�L�<ї&��	�x�rqH�)������d�<!�Q�N���-�L��#p)�c�<ib�F
'����J��w�Z){cLf�<���9T���Cǀ�Oqb����o�<�寉�F@���Z�,�i��_h�<9��.;+�]�����%�u��j�<qǊ��R�@�"7��KAl�<�'G��cw>(�C�ٷh�x��b��R�<� ��_?�B��,n�[@`b�I�<��"P�9��q��Ff]��!!�X�<Y��\?:�v����R�TyQ�˔P�<�M)}���bN��w��8̐g�<����&���A\/�h �&�]�<�� ��)��s%b VzJ\�a�IM�<�b�SC��St�N�Un=�cIIC�<�jRO\�5��C&{@�h�B�Xu�<y��[+#p���uNڝP��9�Il�<����6<�7�E,~�`1�Qgj�<نKLR~�j�
�L��=�uN�o�<IƂG�V���1��&��h�Uɐb�<�WŃ�B` Y�E��Zz^���n�X�<!Ǧ�� @s�Y+X��r�FT�<� l��QnC���1��Sذ��q"O�Y�w���F������³z�.�r "O`|�R'80�jE�g�:Xޞi� "Ox��d�P*PH2��D�(���h�"O�A���E7��j�c�>��X2�"O \��i��v0:&��CD%x�"OxD��)C"Yk:I��M�$*��6"O� "�I�RP<ȩ�Ɠ�()V-�S"O��Х�ψj)�pJe�ű.d]@"O~�)β^����$,��I5"O���Ł� �<�0��%c{�rG"OX��'�c͜Q(�ÊcW��"O���p,O�f{��4�|�D"O�Ԃ�/��U�uz�M��U݌�z�"O�)q�
�_V�= c�(s�����"Or�a�E�4K�|[��-|��1�"OT����EB��a��kU��k�"O>h�A�[�Yh��%�ʨ"O��"��]:�8\;VD��F�x��0"On������@C�C�!�iu"OE�5�	f�@P�`B-8X�"O�e�D�\�j	Pe��2�D(9�"Or��f"�mଉ�Bꃲ��Q"O�9��ߊEɳ�
3{l	)�"OPa���@.����H�u��]Rr"O�\��AP0|,�Z�ݬ��@A"O���W	��h&�2��Y�Pz��3$"O���$Ng�`RAD��LpFD��"O�E�cȑ�AN�%A�!I"X�"O���яŐ)U�Q���:�c�"Od������UK��١8,�0�"O0�KV���wH\cg�H�?����"O���!�Q�H�B�^�2�X���"O%�aָB�8ٖ�Ҙ�"Ov�HU�š{�ыZ=6I����'��Lap?ED�=�T�2�D	�'��bb.�o�P��ǂ$g����'Ld r�Bؕz����?(���'�� �_;'V�|����--�`�;	�'����g�ɺQ6M��i�� ���'5��B�͟S����)�*Â���'�{��[�f��$�T�D�wvq�
�'g,@�Հ�v��{�׌i��< �'�L�K�3)d�S�]�3�$�'_"��b���{ѲBM�:4� =��'3�)��Z!��C��$�n5S�'&����O>6rp��Ŗ Ҝ��r"\?<����=E��'9��8U�5`d���mX�H=2�
�'��IÇ7��5�4�2Hm�p��D2tl��k��0>�3���}���I��4+q�R��B؞��6��\-L`C0�'�^	v��8
�Z��
�Q���)�'�p�9���cB8`��'�+W=t-��}�J�Y�vĂ�g�Z�O����Uk�c	>x����Q�>�'jbl��DS� $:̛3 ��=/�j�f�5C ) `�>���>�ҠH�KE,��FTz$�h��u���g�Q�)�	�)$bU8�Ȟ,+X�4�G`C�D�7�-	����勛��=yrBPrir�:��)_'1�jH�G���TbI���䗨\-pb�R���qo[N���1�`զd�a���E�<���*�rX�+� ��iR� 8Y�r�n�A}RO�.��2�J�'*���.d�Ԁu�"|1�"L>5$�B�I	"�pDEM��ƼH�IQ�aր �+�7^�`+p/�>i���\>�)�&;�	/]5�#��ٜU�m���`S��?'̘'fqR)M�9:X�Y��Oè8�fOR�&tzL����Z]�l��l�,qB'G�0>�s�_D��]��dDP�Dٺ�˜p}�Z5'&��Jt*V�X�偡o&
��j���3� X8K��C��=1�]c�b�p�"O�H��K�E��rQj];��")��h� �p�ɑ.��]�����"��'\,@��H<�v�ԥ3��	ؠMY'JP�9�^\����wg[W����%�[�"�*0�@ <G��R�
\d�{�[� !�#�^	�p<�ꝸY������2��Pp�Z�'�ԕ˥n��.���xP#��z�)�
]�E�b��cW�B����2S�C˪=kn�n<IwF��Mo.��&�J����V?i#�7hx
�o�t���+cߤ2Dy�A'擿Ax���2G8T�у?/�B�	2<քw�M?�8�뷯Ěd�a�G��Ĥ�aߥv���LD��ýM���K�O��!���-F��q�w�Q�<��'"]X�M����o��`YRrhX�gH�ъ�`?�V+�E�B= � OtA���,_��`��Hߕ� d	��I����O�X��d1�����5kZ�(.0�Ij�Y�*2�5��&J<	t�ǧP�D�gO�!h;�=:���x}�eJ�y�Q�A\��ۑ)�([��3V�)O�Z}�������(o�!��=<eH=�D_9� x!Q�ى&��ę&����G!	#�L�S��OG�I<O��9�'R���G��6"�B��7hJ�SS(Q"~�MX%j���O�E���3'(��2��ڣaą#�BA[���
����2˪d@�9/j���a�T�`�)W�
FH<)e�֕i!� `�(���&!�A�<!��R75Ƃ�)k��u{�m33�]|�<ɓ�����P(�'7-�@� �H|�<�1֮Kmt�
��hNĈ4ǐz�<��΃�\���+c�Zb�U���@s�<�́8#�~�(��VuܤS�Ij�<��-	w�0Y[��=��ȇ��S�<�'bKPU>-K���=8���L�<1�Q�2Z�/� ���qg�H�<����]��șB6��*SI�<�NF�&��1�1�&/x*Xz��G�<�҈26)�%��X�?���C�}�<�$I�V�`��O%U&�� I z�<���=WaVIK�!�er>�Xq��{�<��"^�W*2�+Ў�,$�#�}��B��܁wqOԁ;uk�[N���X�<�d ��"O8�5�-48x��N�E:�a��]��(�@�8M�$��|�C��*�gG		(��m��Vh�<p���l����J��];bF���I�%JՃ���g�W&����5A��2o����q�\�5�D�Y�(����I�j�qq�rZ���'��13�ƂZ(Y�vd��Y�*9����
?��)����'`�
�y创�O<3���l:݇�F
N%x.r/���ʄ $l��'��+�ė�XW,�O�>eppꀗ%z *cԥ(��Ġ`�<D�|Kt
<����k���t��!a\w�ė�>�ZS��y�3��\p�R+�:X9�����ԳD����D�6���d�<��Ph�BM�e�`bw�YH:���pJ�QX���/V��K�	�M��%E~R̂�_p�� �Z��(�s�̑�xX�]R�!�/.�C�Ɏc<T��E%<0p�ݙ*��>������a'��(��S�Odb��P����m˖Mͽ(��X��'�:����B%�칒T���ӍyBK�������n��0�M�(1h(E����o TC�	� �n%rQ(�k�!AF�@'/�
C�	Af��Uo��(<�2A/C䉰8�,`����N.�s��2x0B�ɖ.�u�փ�6~��IHA�

sI�C��)<@P�A�{LЭ5Mɼ&�B�ɠp��l��"oz:o�G��B�I�56Y��썫>�J�c�C4+�L�'|Ɲ�#�DG�S��G8BP��5�����D�;/��ȓB8؅#]�x�ᄄ+�2�H>�a�)�:�|�<ADI5g�������;Z����3�[I���Pωt�? `!)��A�2���Y�\. p���1�֓A�P��I-)Zya��W���zB�/��?y�E�Z�zP��)�Ɏ#\0P�ޑ2��|"��}!�dټqq�@�A�wz�r�␟5剕IO���A|�I�V()a��I�����th*fz,8Y� K�V!�� ��K0߹]iz! �W�>��9�'���r�K��"�R��O~Z�끢#����u��鑯D����V��,'����� �ḣ��=[i�����Z�x�����=��̣�'��ѻ� ��{�h�E~R� |�u�a~xe+'�΅��O���WY&����'͢Ţ`��f-ș�T��<+_�A�S�ǭ�@*�Y؟�(�`9{���F�es��+�J�<��a���ﰟ$/��$۴�@����+ùI~y��a�+������Z/�y�j�D�Ε��j's��L㐁޽8����'U�,���eڅ	���%?��U%���*�ƝKp$�$N��(9P�W�6b���Dˇ)��e�c%�-�Nx�6J��.%R���=\�T��'x�d����X+*�E~�h��Z58(P�ł�1�ƌ���7��On��  �����'(��k�|:�����\,Ťd06�V3*�X���HX؟`���y2֝J�HԆms�,3G`�<QW�]�R��Q�켟��c�;P��ʠ���Μ'���cs!R�x�6��l�?�y��]��� �R'v~-�0(�'w��I J��E���!��c>Q��L�ayb�V%�}�Bk��iaּz񡞝�PxB�u�v�{ ���y�q�fLD �Aw(W�DM�� Hp�Ŵqa��J��i��9�:���1���HF'Q����6h��m�ȓi��T R�K�w%�LyW�~|B1�ȓx�����)5���.�.'���ȓg?4\�&Jc!p-�d\�чȓq�MB���#d0�����k���� OX�+�LI� M����J�>�*h�ȓ9��pQT��0Z�h��'�$���Ve��s�&ҟ8Tl�����b��ȓeL�0�l���%lСGmY��h"�{u$O3� �����"TQ�ȓ�xŪ6m!����ȟg�@��)gr��hb]Lݺd	P���ȓ~������Lo��aA�,J�x��D �"��'b:��F��,��ȓt�\8[�)��s�H����#,Td��k7��{���7I�Eb�^ذ�ȓ4���A�N�7{|d2��P�M�ԭ�ȓ�Us�� CT2�C�*!�ȓJ�m����ހyQb@W�,���J���Aܠz����o��5��e��`S]=��i�+���"�ȓEPl@��!��gT20�V�̎��ȓA��R�f� R�("뒅*��ȓa~�"&�c�2a�`bK�5�ȓEɄEy��֜u�e9�o��L���+Ǩ�@���a�"Y#i�-3CVi��=O,��� ���H���X>�ȓ~�:@X`bְ1�|����S������� NϏK�lлՋ�+�~��c����W͆�A;�ً,�0�І�\:����R�'�t9�Ώ�|��0�<a.N6{���0E+6Y��V`̓zf�@�a���m���eD�x��ȓ|l�:�-É{.�S��U�
�:@�ȓop]�"oN�dD{���)\�P؇ȓ�JИ��O�{fDJ��ܤpsP	��?w�U��OUF�9����ȓ}~P�k�l��G3rHYSjI&�����E���2��!��uX�ԇȓQ�
�B7	V�m� �%V�VEL���+�T��%�):R�Y��-r�]�� ]��2m��@���1���H��ɇ�S�? 2��CѰD���@%� v��U��"O��7�
g<�U��G�ƕ�7"OB�`���fYvɺv+ ?����"O\I��j��|X���8@5"OL)�*Ȇkᦕ��$�U��E��"O\@��(w}���K�~���'9�zO<)p«�ȟ�l��֣`׈�rLY�F�����O��Y���+`˛&IY���)�O��r����<u2E��`O��Di�G�)?���4S�ɨ�M�s������<�Ot0�U��=O`J�c��K��h�ώ1X���=���ن%�]>@ ��/�rȨB��aT���T#�<�1�J�Si�U��M~��閟A�M1�A�	-�̑1���H�$��S�`���������>Ɉ�H���&���GY">Ȋ��>QgG�r>��r+.8�5/��(O�e�ܙ-��	�uP� 
$��y>�+f-��|M8���ē,I�<�An�<�F�O�6 �� Gy~��)J#G�r���q�H\���`r(�X��$���{ɬ<
�ǨO��*&�ԈT��t��FϢ*�.�3�"OPT�V@�e9R�0��U�)�6"O	��b+3�D4��#t��la"O�µ��x~aP�`�� �"O��g��	J`�ۣ��C��I�"OرH�c��ip-�	=�uB�"Oج��&ž�
�l� ˖�b"OD�j�����@�Y|����"Oi�R�t?t�A����>�2"O�}23j��Q�d�oެ!�b�"O�YR3�G��*�#F��"G	FD��"O�m�a
ݢd3X��5V��!��"Ox�{f�)$NJ�m�s��=B��7D� ��  g��*d�ä,s�e�T�4D�d٧�ȱ	��Q�ÆCNN���<D�,P!���4��Yy0�T�y��S� D�,;�K�<�)kp� Dt��v D����T,f��A���&1�B�c+*D�L��?!�ip5���X�(%((D�T�G��96�I)��݂]ېY b�)D�D�.�*���i��ߺwv�룠"D����[�p��]����)1v:Y��D"D�@x4*�45v 0�b���L�j|�GM,D�$�T��
l	~dxs�(t+f�C�6D��p�Ĝ
â��c�;Mrah�G'D��x�-�`� <A�� ��cխ"D�(C0��!yL��@"�?t� � �=D�DA��x)�v�Y� �)*�	�^�!�Ve	F-[��i���H�K��[8!�D�I\�Z�ϧ#ɐ�yB ��-<!�!D���d�ΣeŔd��o�H*!�D�7X�*���n������!�P�D�����0D�,�X΄2=!��N$>4	`�.
�~c8��a���n�!��-2�\8ץ׫8�t,�C)m!�D��;��ZsD�'�f�P��ؼk!��Zp��pȭ%�Ĉ�Sj�J�!�$�<�d�`	�]����ֈG��!��3p�a2��Ӡ/�j�x6�%I�!�T�� s�UM�\u3�&�	�!��/T,�AiR;�����D��Py2�X_,�"Cm��8�:`Q�B���yr��B�,��(��7����eC�y�ܠ|�is+-����')�y�)q ذPa��=)h5	�-�y���N�dA��̴$�f����y�mΦB^24��� �wT�`�g��y"�]�H�:5)��&��괬��y�LԈy�5�� �>��|a����y
�   �E���
������*.D���"O�1���6��)�^7��!%"O��s�F�9Vl�2$��n*:=��"O��SAL�H���� L
&S�"O\e%�\?8yB���Y(R(�q�"O��n 0 FU�OςO��0e"O"I��f<к�.Zo!� �"OJ���,�T�Q��ٌX����"O
�!Č[=bT�9R�T"\�&P�"O�\b�G;.���6h
	33f�[�"O�%b��]<tD�A�dG�:#w
��"Od��f�4ola ���Vb�mؓ"O�� '���j�s*�:1[�	y7"O�taֺX�X�3��]OY�'"Oz��������5HT/F��H%"O$Xkp�U�(I�h���4��"O�-R"D�%�����ʶq�ܺD"O�HA`k'&;��7'�"0���`�"O�A��C�X���Տr��ͺ�"O��� �̾p�ޔ�d�)ul4]�"O5)�C�$]t9��)y���"O8�P�k�#��{��ӿf�`B�"O�8
T�ߺ9մI0HU?z6��"O�Q`3��d�J�R�ϵzq�i�"Ob\	�H�G:�5��d�F���ȱ"O橢$�D6F���k��i!�/M)3M!�ė�[�=1,��s�ԡ��� p>!�$�"���d%����G!�!�DK7.����Xc¡�2�N3K!�D� �:` ta�p\�Aa5�8�!�d:bq��9!�8;��%I�Mƙ|�!�� �B��L(g���aN�1�!�$3^�%�4�%������2�!�o���a��tP*�(	$�!�d�X'��P���}����SIm!���p�k�&y��8"�Ց=O!�M�%P���0`v�U��S�rI!�A�Y��a���%Ü���x0!��	~�6$;6�U�)���{�m�B!�$SC�88��3�
l���֚/!�U�1I�M���.e�r����D�!�;�ި�@h�3�CƤ�6c�!�*	B:MZb�Z���Q��b�89!��$|{�)%!��y@q@q䑵)'!��t�(]a���.@D��T��Ws!��A8���"��.-�u! !g!�$�up�(j"�#'�X�0��T]!��U����%C۵u�Ѐ�P�U!�D�+gs�Q�¤X
]�
��4�O�,�!�FQ����@�P��qyD�۔�!��N+�Z�P��M|f�r7!��P�B!�1��~�T�V�8!�D�������&U"�A�+�^�!���Rm��zg ���x�*�7V}!� <����h��HmT�h�*R�F�!�dV$�� )�,�D$aS��F�!�S�_��}2� �'/�0���	o!�$P�(���ѕ�M�5�a�M� _!���JC4"B;Ow�	�֥[w!�D�d�\(uDд!^8��"Q08!�dV4f��T��F�@��*�O�!��˻S}\��@I�&��1jW��;!򄜢S�9�B��'&���j#���{!���?8�$���#ƶI� ���K�	L!�� �1rQ� 0pi9 IK>a� eӀ"O��z@E?G���X,��}S�"O�����M�m����a��%��͂�"O �h#�T#ƶ��%�Y˖̓"O��0v�ۦe�B��u�Z`�p"O6�g��c\(��Ym��C"O��tk  Eڵ�L�)_*�2"Or��ץ	'T��Q�Z�}�@ T"A�!�Z,E�|��hUaŰ�B�ᛴ\!���$^{�+��P��o��9U!��#�d�`$-^O���1`@��1A!�d��Aʕ9��ǟpܰ��싼+(��*R��I�L׷:�,YC���yb��D�|��#���3�`�q$�@;�yBG�4!t��)���B�s�R?�yB���8̠p��35���X��y%ݺ$@3�`'2�@9[���yR�"O�Ց�"��}�����
�y�F�� ���#��E4}�,m��I�.�yBH�kW�E ��?#���dN�y/�&�J��Ɲ!#ʰ�ġM<�y2��_��|!�"�P�+���1�y⪌�2O5�c�\�f`lY�dܮ�yrk���"��M����Bϔ�y��ڕ���'bCaC�D�8t!��5.�TI@�ʒ�T֌�q��15p!�� �Ƣm��n˳fI� z2�?<!��`�ޙbg葨21D��qJ�q)!�$ޒ��L@�j�(��[@��I�!�D�m�#��D��r �ݹ�!��F�N���M|��E����X�!�D�h�(�����x�� ���*v+!��	�f�{p����� 
O�Yl!򄑏9��k���+ �r�@R	;:e!�E�!a������6�2��	�a!�[F6IV0mh�ER??�!�$P�U�hg�������e՞T�!�ƫr�h�T�rC� `KE�!�D�Y����WH.x1N�`r���!��/UEY�J�"+7Zl�`�V�_!�D^�R��E����Q~�p����-�!���1B�s���"yl���eY�2�!�DP�u�&|���Z�xj�1
��>L�!�$����m���B�ab��WZ'HQ!��8BX��х��V�5�]-k@!�$J� 1FUj� )*;,�#�� �!�R�-A�\r�ڭR9d�) i�(�!�Č  %\���	��W�ֽB1nU�L�!����r��9�M�>����w�U�!�O2}��p�Wi����Q;�D
z!�ĉ&"�ASPiRv�����կ<\!�dC�X� ��Qa46��ӓd��kD!�dEN���W+K9"��]*�$�+i'!�&r�]a�I�~hEZG!\<j	!� D��D��>�	���� eY!�dQ�5/�њ���"l�x�cW4bZ!�$X"��s��S�t���(=!��
�cr��0��O�O@�E�>-!�/]�t r��B�"0 ��џ*!�D3k|�1�ª�&1)��+�� �!�Dɷ����,=
Q�Q�G�!�$ߴa���Z��/
V���
��\�!�$ͣ<d<���U+u&h����\�RB!�<�̥��!T�=rt��(5!�� ��t��W>�����8M��I"O�\��S�$��D���
�g����4"ODqh[Y�]�M��Wm�����x�<)%��J�xYd9NZ���$�q�<aF�� "YelN�dr�����k�<1Սފ;��]�#�#4:���@D�r�<�HF"0���z��]�8Ma�i�<�q��V�p�k��k��ģV(�b�<�%B�PÖ�C�^1��V�<)W �4?zS *�<9�5k�O�<I��^��cvc �.LT�
  �P�<�թM����L�R�z=z�!�H�<�5M�(6�D�to�T���E��j�<�t-J�=:���R�B�!��m�<vgߞ���hU�h3j�ks�DA�<94'�����
}6-XH�s�<�m?'ި �S�Յq ���i[m�<��

I0�oO,:1ޑ�g�~�<����4=�d����Ϧ2���$��x�<��!    ��   �  G  �  �  v*  �5  �A  M  �X  �c  ^o  �z  !�  R�  ��  ��  b�  ��   �  H�  ��  ��  F�  ��  %�  ~�  ��  ��  ��   �  c �  � � �! * p4 �: �B �L kS �Y �_ �e  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&��Q���I�8bE!�۽}�6����>:�!��P�K�`U�1� !�,Q�~�ўx��)� h����M�+����&�R�z����p"OH��e��%�>q��/�*S�����A(4� A�'��ޙ����3J�Z�H!�OR�O,j��I���a�)� �|-�"O�Y�C��"Њ�ÇC�@�"OHh��ϟ�P�Yɧ![�T�T1BO��D/ex�5�qL����eoĶ+!�ʻvBPa!@��P��NF0�!�d��?T�5@�Ή���\�D�Ӄ8!�Ğ?ZJx�mN�`+8<9�	�,K�!��\�'d��Ǎȼ&���r�I=�!�dR	�n��*�-Of�����L�y!���H����%�� !,�D{S�QMY!�$
-t����&H gl,�rao۩N�!�D_� <�9*��j��0��ÃO�'�a|���10�Q���§'R�A �Ԩ��?!�'�J�r�/E�3�v�(b�Ȏ,�����D�~�O t���B�nm�Q� �UY<��'_(���.V�d�<���?0a��O�O>\F��O4�a�7V�`�v�S=6˂��"O���3k��d\$��ѤM�wY|DR�i�����Z�H-pu&֌3�2�8�B�%JUa{��C�jj �X�`˩2�`�����G#!�Ĉ��,d3a� �+�2xЯ;7!�d
�)i�4�q�	)����'��B�!�@+.Q�!o��Q��9��n�0tf�IB�����2 �I5/��x�Wi�U�F�:�"O��f	�)��)cQiMV�Nur"Op��#�Y���,��H,)�|��1"O�x�7�V�a�&���HB���"O�m���E�d� ��#DHj�"O�e�Q��m�\Բ�G�_�Q�A"O�5���G.m�
\ ��?c.m�"OQ�胱Y���	`H�/�V �P"O(M�Z�*BX���/��tc�"O�J�D(�lA0�%A!���"O $�2I
7b��ˁ$�
�R �$"O�`G��$��b�O�^5��"OΔ��%Ŗ6����GB�-�	�'ӂ�p2ɜ�#�*`�ąz�p�*�'�!�%oEgH�����9KZ���'TԊQk�$H{�A��ăs2DaK	�'yR	K&�Ҧ�!g'^�q\��*	�'�.��w+��	��5�'Ă�b>�K�'�b���(ŐD�m�E�^�T�H��'��u b�I)�~` �KZ�,���'�V��"i��+��CO� `�'�`)!!F9c'li�'�DYb@��'4��c �K?Qy!���K�̖p�<�ԄS�N;n�hE
u�Z�!@�]b�<Y6*� TT)�vb��@2�PV�<Q�j/\��6N�v�6�{$��U�<٠!"�H��2bH]f� 5�PS�<yA�d�)Ӣ�ק^��ٓ�χj�<٠����v�ɕ+��l4r����b�<���S����5 �;{�Ҕ{4�	U�<Y�l/��st��Nr(�p�G�<�R-ص;Π���G�캤��F�<���K�Hi�)�\+�z�jDY�<16L٣��\"���, &p�qL�m�<�"n3v��)��k�r���"LN�<�#aKM�H�'kɏ9]
��g@�U�<�#�U�Wi���(���� [�<�� 
���)�9�ȠA��Y�<� ��jrF�,JOX�)�4=Tf��"O�=;���>�1��ZAn�z�"OШ��Qt�A�r�_�'\TI��"O��ɇ!��R��T�$]��c���yba�)v�Nɡ�C��.����6����?Y���?����?A����O����O��B���>�ɒ��S�
[��B�C�OV��O���O���O��d�O���OJaC��ƹGBD p�f ���U�OF���O����O ���O���O����Oh80��3dZ�A����O��(�d��O����O��D�OF���O��d�O����O����SZ@�>t�y����O�$�Ol�$�O����O��d�O���O�f��g����n��T'�l���Or�d�O��d�O����O0�$�O ���O� b�ٗ���W�$#U���OJ��O��$�O���Ov��O��D�O��O�Z�6-�A���&8�f��O����O����O"��O���O2���O��
T`�$;�&�t�
򺵲%��O����O\���O��$�O����O����Ota��c��5.\h��.��R9q*�O>���O��d�O��$�O���OX�$�O�e�¦�?����,�8�pl�Ѥ�O����O����O����O����Od���O��A�
��@)"\�#��$'V�T�7�O����O��D�O��D�O�d�O��D�O�L�H�1���X��Y�t z�B�O���OH���O:��O���Ǧ�������F���icFパ	��]�ả���O$�S�g~��cӘ�w���j�IW�4t��#D��%P�����Mˎ��yB�'>0E�t!U8K�� �Ï�,Z��k��'2�9����8�'9����~"ҡ�9l�0�0I���,��$R}��?�)O��}j��SZ����v�U�<v�"�H��2�ƥ�٘'�	nz��)ܭ���KW�E�_�T�K�(������<�O1��xӆ�ɀy{ڴh���O�4Љ�	��>��I�<��'��,F{�O2.^?Q+�\)&�ɟz�&+a��"�y�R�x&�`�4=]R��<��ܹ�2����:��������'�b듵?����y2[����
f����/�J3:�S �=?��ȕ˦`Zs�'���DZ3�?��+P;�`Q�$xb��r����<��S��yb!ʐ� 8#E�
&OC�\B���y��i��q���`��4����ԣV�q]pltϊ@��I�PL]7�y��'�r�'����i����|J��O�Ɓ#aU�*E8x{�G�m���Xx�Ily�O��'�"�'���N�2��ЈJ����I��	�M�@"�?�?a���?yH~r���"Iy�͛�D�L� � Q�s�L
�Y����4@
�x������rm���]��9j���q��D�S-�#D��P���W��O6�hH<�_�`�Ѣ�-�ʉ�6(@�>a�`Z��쟜����$�I��Sfyrff�j-��6O�P�q��D�x���ȹ�)��6O umN�GS�	8�M���i^*6����Y���JȂl�&��  �M��'�X!Y�.ۑ^X����_��'�u����vM1f'��0���&	������;O��D�O����O���O��?%r� Ůu6^�)�L��ԉ�'�v���Iޟ���4-'d��'~�6�,��Ջ5/nu;bC@�Bs��Ps����N�$���ٴf���O
J�)#�iQ�ɪ?\��c��9~�B�#�"c2�`�!�S38n.|�sy�O�'�r#T�J� ���&ɻ[��D3�ӊA��'&�I��M���<��?Q)��x:WJ@�9S���WЮxBF��P�����O��oZ'�MK��xʟ��A�ԚvA��PnͿB4z���*�N��P���)��i>E�r�'��%�h��f�'�6�@��-#�۱�T۟`�iYn���)�ayBgg�$�f�ɽ�xUp�#�Z,}�I �PG��?�M���>�i]^Ѓi@�����Å�+��aԣe�4	lZ22t�mZ]~�I@��8�S^��I)�F�Y� �Z(��C6*F�i"��<����?Y��?���?�+�P[�n��#�QSa��H������-�v� ?i����O��7=��  ��;�ҥ��bA����������z�4q艧�O�S��i#�d4] �!ۡi�?�dh;@�L�y��d�7��8��$ȒO���|����)j��ѾNf��#�
�$\���?a���?i(O�Pog�I��|�ɅR����3$:��Ҳ�B�@�T�?y�X����4FK��++�
� ���	ڼ4ʃ�7s�ɚ3
�hrh?o5�P$?iH��',�T�I=$���]�6�@ԃv�II����ߟ��	��X�	{�O�rb�'p@d�
����pC�� f+��m��� �Oz�$E���?�;������Ւ���t�#�@�����%|�(�l��H�m�E~2���F�����Hx�1)Q�Ej��
�-<XX��|�Z� �	���I����p���{_��+��ю�Ҙ��!]myBmy��	Z�F�Od�D�O�b��
�__�$�#d�	�v�QT��=��H�'��'O1��9���T;T�� �āS6�ླྀ�*\�=��7-�@y"��V���������5&�ٚ�'?Y�Ή���I3t�R���O��D�O��4���nl�ƨ֬y8"�>e�����H�Ң=1�k�x�Bjz� 㟨�O$Uo��?�4:b`�Ac�ΑwH!P&A�{��X[���M+�O��2eM�s�4����� ��s�M*g�R�`�HJAO�d��;O����O��d�O���O>�?���Ɗ�}�t�0DN<@�x�%��L��ϟhs�4F�r9̧�?с�i��'�d��ӊfmp0�-�*^�.r�'�:6�ʟ�i��c�J6�<?�'�J�ɸL�0��á#D�7��=Q4@�O�HI>Y,OP���O����O�ep�5��2��ֱh/�h��O���<)B�iP�Tsa�'���'n�SG߮��W+�'X
rY3���9�\�H���=�M���'����	� d�>l�D˔�i��a:��Sf����U�1�޹9�l�<ͧX���d�2��bURp9��~��2�c��F%����?A���?�S�'��d�Ʀ�+��P�7�Uy"��{Vv` �@�.Q
���՟���4��'m��
Y����$I�(ub��Q�h��MZ�cU3y����r�t����x��[��0������+OvqVg[J�(B ,Y�'zi0O���?I��?q���?����׊mL�Y����lÐ�b�@��-&�m��PT����D��m�S�P����#���/'~��C�ǭ�԰�WeR�����O�O�I�@�I2#�`7�h�,�w㈭#���xЧ�č2��l��:��Y�$W�J�z�	Iy��'~R�̗8\0qPAň*��Y!ek�3��'W��'��iu7m]<T8���O8���5��=�IF�t8n1��E�Jaz⟈x�O�1n��?J<�G��'Ŭ�6��#2� ��EY~m^��I�DZ�"O~B6��OZ����T�K� �5X`d�r��\��=?J��O���O��*ڧ�?�EP�` s`Ӣ!"B�Idi]��?��i<� St�'���o�4��6ot�˗L˾!B��x�hʹ
����M��'l��@�7������`�gJ�	�[��n�"˅���䊚�xh`&�ȕ'�r�'W�'n��'Ҋ��� �q�>�C%�;bgt<�#Y�<��4nfj��?)���O�E!��Ӗ\ܠ�7�[�,�s�.�>᥶ic���"��Iͥ�X����$��lBD�CE��A�1@?{���-��gM�Oĩ�H>/O����.�v����Y0r��䋴��O����O����O��<���i�)S��'�(�D�jzl%���2VA�ɸ��'I�7�/������Ħ���M�τ����ra�Sb�m�ǯT�4�rĐ�4����*����'f� ����Nʝ~�DbV�xM `օ��i��D�O���O,���O���1��2?(��  �+<�{�'U|p�9��Ο�����M+h�|��U#���|b�(:2�"�"G@����D[^v֓O����O���z�&���A"Jm��m�uG�0�\���̡t�R!�&�'c�e&�,�'�B�'���'`N�r$�
5I����#�DW�n����'!�X�,��40x�=��?����i
RvU�B}rq��h˳�����dS�-P�4X����ɑ�{���x�i�<u��q��F˭5g�K���+w��擴,���r�tBE��[',mLhǊl����I����ן��)�SFyl������	�m�$wn�d�1D�7+�ʓ@�f��B}"ml��]���,�V��U`|��q���i�ڴM&����4��ăQ� ��'W`�ʓ�b�k��Q+s�]��k+��̓���O����O���O��Ĥ|�⅐�-�x
0D��?�Q"Q�ہ>���F�B�	ʟh%?�����M�;��
P�W�zؠD��]�`=1���?���x��4�D�3I��6O Y�2�G�|�,�2M�s�"��b3O|�	ç
��~��|bU�d�����b��=Z
�ږ��1L8����䟜����p�	Oy��f�v�t5O|�D�O�Pi���'J�aR�ě�;��h/�I#�������ܴj�'�4�5Ā�/Τ��yݠ�O:��ŕ�|Z8�a�	б�?�am�O\[�,]'��:��h(��Ќ�O��D�O����O"�}Z��|�5�@D�hւ\8�,�4I�������&A�������?ͻ"�n�l�~a(V*�G�H��蛆�zӜ�n�K촩n�i~��T�-�v���B���������k�/&J :e�|�[���H�	��d�	�4�0�	����C�Y�l�{�#�Cye�"��w3O�d�O����p0R�oY�
Ja�o��'k�6�@榭KJ<�|ZCD��}�6�8'D7+t��#@(��E:� j��BE~2�P��v��Ɇ
��'��xK�Ѥ�nQ��!�'M!
���H�	�|�i>	�'�27��(�&n����
 t��Uk�M����Φ��?1CS����4Aڛ6.s� e�V/C�d�8܉k@2C�q#�GL�s��6Mt���	.n0���O� ��"��g�8T��bZv�L)�S��A��e��?����?���?Y����O1P�c��lz�z�d�'�'��'��7-��R���O�(nZd�ɘt�qq+�>ʴ*���.�j�QO<id�i2�6=�@��Reeӎ�2�$���<L(���Y�@:�c�f@(EP��A�����D�O��D�O��D�2Ɛ1j㇟\�J�@ퟁci����Ox˓hH�FP�c���',�_>���H_�<,�4�v/��d9d=�F�-?�]����4e���j/�?��S+�=_J�jC���+I�x�b�V�>�0L����6������L�P�3�|�͖ ij��Y�Y?2��mQ�&[���'�R�'���4[���ߴ5h@
��.ZȜ��B��TƆ\�C�M���ċ¦��?�BP�D�޴KFN�:�U�v�x0��.��o���s�i�D6���j9r7"?'b�y�t������� ̔f�T�ۨ���$�"[��jA0OF��?����?����?����iڟ}rPaX$E�&	4>�㵀�T���l(XǦ�'0�����'2�6=�
4����x�-�3I�9}Y��+�@��n�1��S�nX(PnZ�<�4ѠC`��цS
jS�����<��i �Ȏ�䓓��Ot��V.�N	0c���5c#bG=�����O����O��TL�F���'�B�[�8�`����p�q`'I�C�O��'�h6B̟�&�
���
�0�	��C[Z�9tL7?��χ1���uh&��7�����?�'*W?F�����I-��C���?a��?���?ю���O$L�&��5f�\R�C�-�(�rf�O�o��:Ӛi�':6M1�iޑ���w�h���MW�I��X:Qf� r�4^��&)r�|0��%o���J�(Adb�|\C�IX�mI(�Z4	E�NW��X�������D�O��D�O`�D�O����G��q��k�b F�2�#ۊ,@<˓��6�/���'����'V\��bM��R����I��H�;��>���i��6͚i�i>���?!��D%_�E1� ��>�tP#�76uT�Q���Fy2�#����ɗ~P�'��!}�0��P��nX��ۄ�͓u=����ޟP�I��i>}�'�7�L2A��Qb�� 	�䔨N;0��%�ߑI�D�Ӧ��?�T�`3۴^E���oӴ AĬ�hn��i��ʍY�B��#�6�)?15@$"A������'���g�Y~��� &K)t�L�gk��<���?����?����?����ۼk�dmp���U���@c�	]B�'��C`Ө�� �<�g�i=�'�x[d���
�ݒt
C�v�6`�!�d�O07=� �(â~�`�Ud)� H(=k"���`Ɔ-�r���M
���������D�O6���O���D�<-PF+v 9	�MY%;�����6�<!��i�P���'1��'���"C�p�Z��4a]��֤ד~�o��ɳ�M[ �i��O�',RVp �-�S�
���K�	!�p�¢DE�n�:E�Hy�O���I�Sc�'q�͂��C�����������'���'���O����MK�� 1�>��'�:�ҽP�G�Lxv
���?���iN�O�X�'�6�U$nM1D�/�.�(b��;=\Tn�!�M��H��M��O A���.��b�<�r�G�rH�	��$2M�<	/O��D�O���O���OB�'q��a��,��(yE-�^��@a��i�,����'��'��d�nz��!���5���J�3'����M��iK�O1��A�tӜ�Di��T�%!*2�u��Zy��	�H-b<2b�'n�I%�$�'Sb�'Bn2�D�t;\��N�h��#��'e�'R2Y�,��4|�����?��9)����ĩ8"@8�G�8}�5ۋ�c�>����?	ӗx�!��w�h��2��2/d��!�Q���$
1!dN��~ӂE%?��5�O0�d�A
�ݙ�kI
jE���S�X���O���O^�$9�'�?�r(U��^�	��Ta���� �?���i�d�!�'%q�>��)q����U(l �\��
7$�	ɟp�Ƀ�M�&	���Mۛ'a�)
)1�����a�KW���8�[/>��K>	-O���O>���O���O �j�_�H(�!�"��D��+�N�<�g�i~6���'�B�'���y����&��'��f�芐f�o�4��?���5
���O�ui�K��r��_ LQ IĻT��F+�<� ႂF!��	@��by"�T55@6�q�˾[LR�j��עO�r�'���'*�OR�I��M�f��'�?�H�C�ҠI�HK�3d��L?�?)Կi��O��'���'�R6�[��x� k��L�����I�{��𫕄c�$�&�f�+&F�?m&?i�0b��!P�Hb��p@G\�Y�	ܟ$�	��t�I����	L�'aBr5�6=��Y�ʀ5N�FD2���?��F��%�����'t�7�0�$�:E������)@��8�kv�'���ʟ��g��l�X~�k��n�豓W�^�-�v�@���]��"�^z?1M>�.ON�d�O����O:�R!������&�960��Iܟ�'�D6D]Q�ʓ�?i/�
T�*��}j
dhaV�}2�ĸ��,��O����O$��#��PࢂO�S���!bR��*2��07��r޴�i>���O��O��S/S
a�HdO�L�P���OF���O`�$�O1��lΛ&hU]�l��!aTv8�:"BݢB���u�'�Co�B�̠�ODAo���Δ�wEG6���H)H�$h`��M��I�)�M3�OF�;��
�jA��<��`����`�̛G|�87���<�(O���O:���Od���O�˧,TBt�e^y,�;��R�Pz�=���it��'���'Q��y�n��NݞSo
���4c�U�ťW�mZ��M+�x���B�;G��3Of����ʣK�  Y"mP����?O�<6oG��?ّ!���<�'�?!'�\g���ft��A{�"M;�?)���?���d�����R���@�	��0� ����C`
�j�ph5��c����	��8�I��ēe�>u�&�άK:tAZ��޷KwE�'�t��\�1ط�is����I�'�2J)r�"�̓&?��҃����'���'v���D� ��:+�����VG�}�G�t�ٴ�x���?��i�O�.F�@�޴p��=`>��q�K�70����OX��ۦ�צ-�'Gب�5�[Y� �7f�0��Г��x��-
�1�D�<I���?���?����?��c��CJ�́�c�+L��
e-^���_ܦ��T韌���`'?�ɼ��9�Ŗ)� U�T�ݜ!��۩O����O�$�b>=x�$�YY�H[�aJ�]�*����"j��n���'<.]��'��'����(yu�'�U
0A�����Ɵ��	����i>�'��6��KI��D]^�Π!�C�)A2�A�F& /`����٦��?Y�V��I����ڴfD�R����A��Ũf��+!+��h�(K��M#�O����BB������w�^�@-͟Y�p%��4I)�hx�'�b�'FB�'���'��6=J�`��e��#U�H�y��ЂD��O��d�Oڼo��m�'ђ7--�H�Đ���Սh-�� ؑ[ T$�`�	���"��}o�C~�� 5bȪ	�g!�i~>d!Ҁ�J0f�3W��Q?�I>�.Ol�D�ON���O,�d�M!{�x�HѬ�.k�p�����O����<��iE�E;�'���'2�cgZ1Q�$���f�5$�r;�$����M�S�iDRO��m��lrC��y`BA52���ж�
�w@Py�O&��I�'�b|b@A�O8ij�ǀ O=�����'�'X��OK�I��M��ɕ;s�,Z����CUH!�w�b4Ľ����?)��i��OU�'�`6-��)�c	 v�rѡ�Ɛ6l?�Qoڠ�M��陬�MK�O%Ss��j�Ƹ<!��ԵG�B�K�&�b�h1����<Y,O���O����O~�D�O��'zS� ��U8RR++Ѩt�P%���M���?����?�O~���	��w��ԈA!�G�� �c?(ԨM��)�OZ6�\�)��� mN7�~�h�7�4
��͓�k�����Ӣ�x�\��[:[���l�I{y"�'t�J�z��g獤'��؈B�ȶ_��'c��'4���M[t̛�?����?YU�����;��ʏ87\�S���'P����vDk���$��zt����9zd��f+���I�G�H����!"7��'?��t�'.���ɐcN$�sĔD5&�	�e��HǎE��ڟ �	П��IX�OAr���8�H��p�@'�T�X��`�b���<ɤ�i4�O�.	�(�6�pm̶W8V}�u�6iI�d�̦��޴T��(�<.<������p�\�l��D%���=���0-�z���䛛@D.5%���'L��'���'L��'p��U$9�<�b�i������Ty"Mo��aqC��O����O����<z�R�r3`�5�,t�-D�9n���';�6�Ǧ��I<�|B�Ŭ6�B}�Q���O�vr4�Բ^��٠�T��DѤ�Lͪ��P=b�OF˓G@j��D�ݟyqʨ	D#J�M�F����?����?���|z,Oz�m*��5�IDȠ��Si�j|�	��>q���I*�M��rJ�>��i��7m���CQ���,�̝���ּsdvv�Kh0Z�lq~BDX�/�V���;s��O�'(� �܅q�*XB$|�/��y��'�2�'�b�'���i�V8��)4i
��aŜ?lO���O������	��)?1��i��'gl���]�P�Y�MΜOJ�$���6��O�6=�Y�W�r��0�T	㱇�[jf(
4�jp2TiG!
z���"�䓈�4��d�OX��KJy���#h�?x`�$H���90[��$�O�˓u���.\;<���'j\>e`gI��f�P#͜f� ����*?�AV���ܴ,��� �?�[���/��І �+2S�=F	J�5'<�In�m�����G��� �|"�ڄQ4T����
	)A>�Ҷ�W�!���'BB�'����W�p��4_쨚4 ����cpCA�����vO�*�?q�9�F��M}�e~�4qA&��5S+T.g�*�å慠.�6��香x�$_��i�'�N͑B�G�?�åR��d��
��N�3&q���j�ؖ'yr�'8��'�"�'��S�N�$Y��_BdE0�L�/�,��4yc��S��?���䧪?�2��y׉��.6�,����/Bi Q�r��>s�6�צ�(K<�|�uh��M#�'7<0�j�5$R�!2S���-?��Z�'��9K������|�T����ßX�K�/F�çI�1��M��ڟ�I� ��Zy�JjӢ%��d�O����O6�����"TD���Ej��� #��#����	�4�'��y+d�L`�QI6ϋ�R8���O�$c���+����;����?)��O�[�NM�S@�P� �<v�!s�h�O����Ol��Oޢ}����٫��RG���C��zX�AH�����C��R�'+�7m?�i�eQw�`�ưҤ��9��������46���.d�@�'�dӴ�t!�7���\�C��ʲ!��0�wg��	B�tq�����䓋��O�d�O����O�N�l{X��Q(0�r��rE����P��+Y2�'���)-Pz��Ц�/U���iG'�%Ni�'�v7��ۦ��L<�|b�jLk�b�I�1x����2򰱃� C!��d�w�hأ�� �Z�Od�	�	�#�f�(�*�:_�����?���?��|z)OĐoڬ]��a�I�g�	�Vo)��Xy#��HӘy�	��M���$�>���?��i%�H	@��:���Y�[/A&lL��"�6k�f����q�;W��=�i��(�p�*!�R�0&�"l�;B:O��d�Of���Ot���O*�?���m&@]��c��x��k�d����Ɵ|�ݴ~f`�ϧ�?�лiX�'��!��X�,� ��&�%cNm#�>���O��4��	��uӼ�O��� �p`��\���x��M��!�6=��ȇ�~"�|bT��	ğ��	۟X8�G�����C|��9���ʟH��gy�&}�F13�˺<����iK�F5y�+���|�nT�%���#��d�O��$S�)
懇�~�8�0�(�S$���،a~�8;�߀�Ms�^��i���4��� Nf�`b�G�{{��Pg�N):G����O,��O���)�<��i4~�s�E*z�⎇<*�[��R�WYr�'�d6�%��8����O��M���|�i���P�N-�7��O0<nZ�^�޸n�s~��QF'� ����č"cxr��(ԣx6H�Ѧ��(#|�d�<)��?���?���?q/���;ь�5@̂�3��^>G2�d82��񹑭�Py��'z��\lz�)"ժ^�[��(�և	6 Cq����?�ݴ�ɧ�'@�J��4�y�)��4&8�)�
!L�x�P/Z7�y� B�����	��'����H�I [>��PaܯZ�D$�'@�40d��	ȟ �	🴗'�6�k#����Od�D�4Bf��ǅ_� ���"%� 	���a(O���}���&�� rHީ+���{��G�0�2�!8?q�f�`��0!ajø��'m�����8�?AD'�(%2�Т䞵)����BY6�?Q��?���?A����O�]�'ߡH�������v8B���O�%o�d͒y�'�26�:�i�;@!�=T1���7(Ҡ������s�XJ�4.���e�h]�PihӶ�B-ht�g���"�#m��D\X�a_Na�J5�S����$�O��d�O��$�O��DܯJb 
�g������=�J˓v�vbW(_�"�'"���'������Tou���V�6Z�2�%ad�I�M+ði�6O1��Q���Y$s�J�J�^�p��k�1:j�D�·<����.0������䓲�D>��,�d.W����j��H�gA���O���O��4�Hʓ����- (�*Tq�Ep�eʯO|<��䬅�y2�}Ӵ��	�O�|n�;�MC5�i�Ve��)�MX�U��/=�t8(�%҉�����A��"T���j�D�S��a&��O/ʑ Iֆ"�H����i�8�	ڟl�	۟`��П���A���WF�hQ�E,w&a��-��?Y���?I��iФ�ZbS��X�4��Z��!C�f7pq�xi�`	,H���x"r�� l��?ѹ�ڦ�Γ�?����d�5ˣ`B�Kr���s��KO�x����O,�N>�.O����ON�d�O�`��'�f��a���Hw��iǪ�O��Ļ<��i�ޠ��'���'T��� ���67�I�@8�l�6b�I��M#��'C�����O$��A�]8V>H���ʲp.|�0��ߜ�&t�u�G���?=���'Dt8$��#A�6_Vp�0��
��H@Ē㟜��ϟ���˟b>�'�\6�Y�C,*�S`@X95d��%Q�b�����<yp�i��Od�'��6��k(Q�@��"q�6�Q�x>}m1�M#`֭�M��'�"�8 �!���)��ɻ|��lR�G��I�(h)Q��
)���	fy��'2�'�"�'|bQ>�ka��K�$���,=V����f�F��Mcug��<���?yO~Γ^ћ�w�Va���H�� 0fh(�,�bu�4�m����S�'[�^�h�4�y���4p��B��*	 `�%���y2�-(����I#^��'��i>	���7�d�V�E�6����e��VL����h�	՟�'�7�T��$�Oh�d����+�C��@K�90�R��C/O��dc���%���PB�)�=�h�,}i��b<?Aĥ�0jT�h�IDp�'}U���E0�?1 ^�A���9$�N�4�|��̐��?���?���?َ���OP����m�Z����ˈ	�p0C!)�OV�lZ2Thv�S��&�4�@Ei� ��5r�%�3[{�Q�79ORAlZ�M��i����ղi.�Ig���R�OB�EKo�t�w����L�q��q�Qy�O��'r�'��A�L񐸲a��/ORu����c��i�mڻ�t������IP�s���3lۨ(��9s��6_�,�Ê\��������ݴDp���O�����,�K�R<B��X��
�bN|F��eY��SD#8bB�Vw�ILy��Q7+:6A���3I����ښEQb�'mb�'��Od�	��M��E�"�?! �C��F, 2�\5Q�A��<!��i��O��'D�7M�Ʀ��4'�XcO�#��Px�4����aeT�B@�N~��ҷ7P����OKw��-S��!����#�h	[�Ð/�yR�'�B�'d"�'���)�3��Bk��R��a9��P-��$�O^�d�Ŧ����E~y�
zӤ�O�\"e��P�f�jan�"�X��@Ne�ɼ�McZ��ɜ>�F7�8?�sɇ�J�$�r��	�~ESf��2DSR���O�`�J>)(O��D�O<���O� f� J�T��QIV�:�b˔��O��$�<�Ըi>�:��'<��'��S^?�53A��M2 �Z�EI�$�C��	��Mkһi�HO�S�Ƽ�:D�	?9���y�
]�}�$9�ŋwh<���k�My�Oqڽ�I�m|�'��ٙ����H��I�ML�mܺX��'��'�����O���%�M;$�!���Ƌ0o�.E#C��#��(O��o�X�i���1�M�DJ�� @�|��S!vi�T�#����6Dh�u3v�o�n�#B�}y����T�)O�DYsi4!2��K�d�is�@��?O���?����?9��?9���)��?�����9- �ʃ�G[�^m�1
O��������@�s�̸���#pJ\�/�	Z���=2�b4Q�@�2R�����O0O1����z���)� ���%H�z����"14Ҽ��;O�q)�\��?�C$�$�<	���?�,�}��QT��<����#��?���?������̦��`L^Dy��'CDD��`I�´$ؓ�� j�kC���N}�i�Dd�	Y�ɲR-��
��+O��� ��=��T���#��&a{��L~��l�O��Q�5~6D@t��D�����GϢ0x���?��?Y���h���D@�}xh��CI�%�8��@S�9�$�ަ�y$��Gy��i�4��}�
�A��"�.�qMY�5����:OD�mڝ�MK��i,¹�W�i<���W�����O�<�K2�˝I>���P�Y�\ �uxT"�h�	dy2�'S2�'���'��+Y)*ah�`�g�_�&PA����=��ɔ�M�B�A2�?���?�K~���m��s!�B��8��cF8{8>��6^��!�4{:��x�����	T��4pE_� ��%) �Xa	a��J&�	b�e(D�'�D%�`�'����r�ޟb%���G��:Q��B�'�"�'!����4Z�<��4�0X)����$;���s���0N��t!���1���B}2|�҈�	��覂�Fm4�� 	�F��P��}oN~�"C�&���S��O:g%��	�j����'`��|��,\��y��'��'���'����!�8�A�%N����TfK˓�?���iKL9�ȟ<in�]�8U�ΜaA�B�@o~��dF�cc �CM<Y$�i��7�����2w&}�:�����S�ό�)��cPb��d@bB/U��ȓ��' f�'���'�r�'nb�'4��s���D���TN)X�a�7�'�2X���ݴ������?a����	�_��9��n�4P���) ?~��I��$\���*ڴp̉���^
�j q���/�����&̼.������L���z H�<�'=:�D���r�f��&�XІ�6��ir@����?���?A�S�'��dY즥A���@ D� ��-��8e�QeS>)�'S�6�!�I��������FF)^f���B�O���ѭ���M3�i�:�Д�i��I(_cd諷�O��)�'�l�� ���ݐD&.��m6�a�'����� �	��I�T��]��� -���s�)�"�z��f.Ԗ6�	U�:�d�O���?�9O��lz��r��r�k��@&�>`Y"X5�M[ �'���Og�s0�i�󤞬	�FmR�&�#e��`�����&k�%���R�O���?�-�4m"�h�}z�k�kB�g������?���?�*O>	oڌ7f����ן@��0U�8����U�-h�Y,�N �?��Q�$�޴W��x��02X 1���Y��f�����)l��6F���
$?A��'�
(�� b3�<c�!HPm�R��;�0�����������p�O�"+-`���L�HԪ�Q����i�X0c���<���iN�O��֫��r�H�xtM��J&������M;2g��MS�OxA!�f�'�ꁨ ]5֨J��`p�(�1/��Or˓�?���?y��?��hF��15�T-}B� ��탣-e�1X/O�1lڒQD}�I�����|���|z�DI�~�hTK�(��%����$W�q���S�''�^H��n���*����j�XEo²K�@I�,O�P����?�%�;���<��EچU]PJQ���ł��HW,�?����?A��?�'�����Y��՟PXG�53LB���*WXq0!��şDC۴��'���yW�ƫ�O�7�ԼKEi��Ϲ�U³
gI�#Db���(|$�U/㟲=�I~
�;��k�$��;�
�S��E3(�|���?����?����?���Og�� ����R\cv�B�aP�	�Q�'	��'��6�=5��'���|r�Y<�x���=X�
%�v�W'`��O�n�!�M�'�����4��d�]xꠠq�O2m)����$̚A!͊�?��g8�d�<���?a��?yB��,@p|+�GK�}b)�3*��?	����J��ɪ�b�П������OˌSaJ#	�0Y ���6lR��O|Y�'27m�Ѧ�BK<�OD�z �W<k���t�lԊWA4ɞ��b��7C�i>UsB�'�� $���%�G�"d���`J��9��N�����؟��	֟b>�'��7�Hi b��?hCؤy��-`�}[�a�<Ys�i��Oʤ�'I�7��4�e�«w᲌_3 � hPć���9��4a���ڴ��$��F90��"��ʓj��������m�&&�Z ���d�O6���O^�d�O�ĭ|��O�V��j6JWgD���r��>z�����R���'P����'W�7=��R���9	u$���C�9�╻��J�}(ߴH#���O��x�'�i�󄖖R=��u!�5��:���'&?��0i�]p�Qhn�O���?�X�1�G���(	����L��b����?���?	(O�o�+t��Y����h�	!2�Z�n�
�u�a�[��^��?pR��H�4<���&��˺=t��3���8�PPl��a���
Q΍* ��3=��Q$?�"`�'��}��B�,��Ԡ�NX����0Yl��	���������\�Omr��L��R�i[�!����!\4�"e��ݡ"�O4�$�Ҧ��?�;@,h1!s��U"�H7eJk&D��?Q��uR��`�%�斟���O#4�醝�A* dɋB�<��� ���Oʓ�?��?a���?��P�2�۱F�+�6Aq���($z�/O��o��VF1������	W�S���i��hRv���F�Q�Iن�"���Ԧ%9���S�'? .� tչ�M5YM��1ĘW4InO�Ak@�c�]���O.�IK>�(O|	@E],~��q�F��sNpda�OP���O�d�O�	�<Ie�iG�'��\����a:��� �gh=#�'� 6M,��(��$��Q��4l`���%Po ���-J���"�EPi1� ���i���A�u���O�q���Λ�M��<zׅ����	¤�%>����OZ���O����O~��=��0S�Huj ��A�z��B̔aF��	���I��M����V~҃qӚ�Ol�s��[�y@ G���-떤�z�I.�M�����t�,F�f���P�IM!X��x`��F0L;>�Q�ކa�����'�l '�������'�'4�.l���v���@�BtiG��-R�'>剞�Mk�E�e~"�'P�g$��h�2o_ 	����(f2�c��� �Müi3�O�S��=2`}h�m�{���1Ɯ�2%��tFl��O�	+�?��M/��@�J�~�H�M� OĆ8`�$Y�����O��$�O���ɣ<Aq�i�<��R6��1%n��|�6Ty�"H���\ɦu�?Y�R�m�)�`�0��E]�Iwc�Y)�}�ڴI��*H�.��P�p�_6EU���~*@�ʳk��x�Ck�3w'Ɖ��f��<�.O����Od�$�O��D�O�ʧEO~a�!A��ZXd�@�ܣ�X(�i*��:�'��'���y��p��Ε�Q����.7��,��� <C�qo���M���x��E� N��v<O�Ż��C�sH"�y��֯'�����=O2�����?
.���<�'�?�A��\P���A�RB$9�K���?����?���D�Ǧ]��c���	��dJ���RؤI�c偏;�
�Cm�g�~o�	 �M�g�i5�O\A�alC�~!�Ya0�&X�@1������E^@�41`�m �ӝ@�Rm���#�iьh*����ܜ> -QeŞ���I���۟,G���'\�a�����g�,|s��7L%đ#W�'Ґ6�K�Wo����M���w�	�RCڦw�P��O�K��Ai�'���i�V7M� �b7/?��Jȥ\������01@q	�.�EM, Ag��;c*��K>a/O���O��d�O
���Oʍ��`�p^� ;��Q+g%�<	$�i�����'�r�'��O�oE�F�R��e;oLd��F�'�J����dӄ�$�b>�#dhRu#.	Pv�ۓ;����dHV=o�� R���Py����Y�M�ɈZ�'�剃ܚt+QW�nY���8��Y�	�p����i>	�'��7m]�z��d������L�����Q�8�D�Ϧ��?�S�,��4t��Aq�����^�PĤN�X}�]*COP�Je�6�/?yw�=u�b�i������a��,j$���ˎ�`��d�<�
�qV�ԡ5nեG�P���-��/O���m���=
԰i�'������7l4P)eG5%&����)*��Φq��|����M;�O6My#(�8sʄh�q(J�N,�v!]#!����4�O�˓��'��P��-M'�]�& U)^�9���9��my��'R�Ӡ5�lbௐ�ND�!#0	]&o���$��I��M �i�O�ӂS�
��S�ܩ�#J��(=8E�	Yd�"��hy�O<~x��f��'Ŏ(�ڈ^j�Hw�	c��!��'�6-�&N.eS�lM(�N0��JKd�2q��d�O�����Y�?Y�\���ɚI��= #�� ;j�!3$�#�.-�I��M���K��M�O�1GGS���d\���i�6���x��0��q���'a�{r�OB�X�D��W���q��0DL6푪,j�ʓ�?ى��y���W��2�-/x"�P���Zu��mZ��M[�x��0|�v5O��T���%$Bi��\�|�l��6OR(�F"W��?���/��<�+O$��&��({(����*�$�a�'X�7�^�>�d�O<�$<�V�sR�	�P4�)��GZ�	�J�p[�O����O�-'�, ���>wǦ� v�B6��Ё�F3?�Al~���P�i��������'
B�C���4�sbN���J��l��P�:���i�'k>�G��3630�I�i՛�蝱<�剫�Mێ�w����Gƭ������'f���I�'0��i�6mH&qUf7�&?i'e^�lr��I��$�.� � ԿEՆ�36�� C�qH>!.O�?�$���23��bž)JBXj�O~�l���s�<a���Ox��ARC�s�f]�!�R�Zp��`��>1$�i,7m�|�)�S6n�@��DJ&E� �t,�#꓉D���'o��-��V�|R]�pZ��D/n�n��6�d�JP�1�OLn�Aly��:Ғ��#�b��B��q�,�I/�MC�2�>�&�i��7��ݦ)xC�\�g��1w@����<Xb��E@�Im�t~�`ݮ5�L�S�x
�O׉?rl~�!��ۛV�j�YAI�y��'� �I�c"2�I�B@�TA�(���'���'�6-�;=���MH>!�PTX;�ɟ�@����Ӊ'�����FŔb_�ƛ����L&lo8ḵɜ�\�|�3DC�C�Lڦ�O��O ���'�N�{C
M�<p��!LZaچ@I���^æ52�ʍiy��'���:��KE�г�@�3J?�U;�C<?y�[�T(�44w�Fn5�4���� H��&B�S[���S�#��)�g윸(i���d!O�8�����#��O��H>�*P��Xu�&Ώ�c:��/e<���i����  k�QH���;e���Q$����'Y"6�2�ɕ���O8и�����Rd,�ڽ1��O�Dm��b�Z�l��<�OQ�l S�?��'3�r$N/1 �tQ�=h4~��'F�	џ���˟p�Iǟx�IJ�4"M�-�$Y�!�ɹ�$� �L�,N6�F�6�˓�?)���!m��CgZl���G�6 ��಍�tC��mZ��?QK<�'���'4��zܴ�y��
�M���y����D��"���y��̣7@��*b��'�	�����*Jw^�	�O�$IK2�@?gz��	ȟ���⟌�'^6M�L��$�O|���TRq)��4<]}k���
`\�*�O}m(�?�N<�#(]�xo>�0+�	0���*��<��)�H���<q�z��)O��)\��?I���O­"!l�1�p�h�n8�.1��f�O��D�O���O��}*��'�J�X3�E�3;���D`Ͳd�((!�"���c����'A�7�(�i��s��������FV�9�,P;7+��� Bx�:mZ��m��<a�oC� ��U�Ѫ�5gubъ���Sp����@	����d�O2���O��$�OH���|䎁��dLJ
��cޫ$��ʓ&'�f����	���c�Ӟ:�Hph����)�ص��oS�hh
��+O��d�O��O���Ob�C�Jʡq��NDܵ��J�d��G�� ���9`�(	S�AУOQ� ��!�N\ ru_*o,MԤL�n3��	���~\����t���ߜ
�P�h�aĐ`�f+Dm\�Bk=H3��,n��he��H��E�t��]��Tr��UP�����RUbeɔ�,�ḎSVjq���'8h �*B�d��T@	���q^>Iz"�\3=ʝ�b&ɲ|,F	��d��)�����"޼
J�j��E6��;��QE:}
�!ƬHD�����Q$?�)��(��
��f�F�R���< �!@��&b���%.Z<o���G|h�C��Ms�a��s�FEѓ�P�/���z���� �&^�x�	[��ޟ|��-^Z���Tp���H���&%�,ӄ0�'�b�'�2T��H&����OVp˱L!1G��*7R���O��m�IR���h�	�!�Ib�D�qL1Iq'_�?�v���Y1h����'�W� Ȕ����I�O��쟆�AEǗ��ȖJª8sj(s��R��ğ����&0��?��O��)�U���R�t#ŏ��l�$�ٴ��A�W��ho�<��۟��S����Ǝ@�1h�%y�� ���aь�Ʊi>��'��Ճa�� @�4[f�Z���fg	!�B7��0J�JToZ���I����S;���<��ə�'\����_hӰd���Z�U9�����O��?m�IC~l�d�,[�&���(~�A�ش�?���?Vʝ"L��ly2�'��$B*���iZ�v���#Ty��OX����>���Ol��Oys�Q��dY,����-bca�9�I ��ʬO,��?M>��O�n����uYh���F�����'�*� p�|r�'���'7��-�|�k�*�� �0E�I-��ܱ��	��$�<������?��Q8l�C��	;<	XhS��P㔹+d X����?����?�+O�����M�|:�(����E��2Ǥ�+�.���q�'�W�t�	ޟp��9VL��QBU���@�&���AK�-�'7��'�R]��C��>��)�OUSCV����NK�iذL	 ��e�IJ�	ǟ`���dcre�=�tG�O��UxgM�&t��S�צ��	����'�
����~z���?��')gr�؅�آGLu��e��bx����xb�'�Rm�$�b�|؟��քl��I�uJI�;����i��h��޴�?����?��3��i��X��J�K#~ ���F'>�U���uӚ�D�O��;��	b�'0�da&,J
�z���T�=��Xn�<Ɇ�3�4�?1���y�� e���4�ȸClr�X��Z��z��&
X� 7�(&��d�OF˓���<��9���CL�<��̀�(�d�zLR�idr�'��IB�O�	�O�����c� V����!�
�7Y��6��Oʓv�3UU?���L�I��
 A�->IB1 �f�.<��z2-���M��'��葲�x�OL�|Zwg�$x�#G <�3GƦ�R�OT�#�m�O`�O$���<!��\F����V4����o�J��C5�ǿ���O�$=�I០��.޶!�¥�rRft�w�ŸrF}�a��=R�b�$�Ivy��'SXX8�ݟp�(!�\3�$	1��)jf��r�i?b�'�O����OH��$$�#˛���;5�̘ �CB�09VM��Z��ē�?Y)O���R�6�˧�?1�f�&RXLx�&g��G�Qr�� �a+�V�D�O��d?6���ʱ�x2D8\����aUF�;���e�t�D�<a�O�&�/���d�O����6�&o���$������ ��qkU�x��'@b�6 .P��y���LR ~0���g c�D��!S����[S*,����l�Ih��byZwG�4[!	D�h��1x�!y�Va�4�?a��_ώ����u�S�')|�)3��n	1o̴tҰm�`��x�4�?��y�'o�����㏪_��D��aT�󲄱�
��
\�6��<	n��OZ���g~�(w�}I6�w�l��6Hr�6-�O��d�O�5Yi�<�O��%�:`0VJ�;N�~��$
�<~LL���\�B%���~����~R'X�g�����K#�HH5玚�M���fK�|�+O��O��O=� ���'��6F)rP@B�@�R� &�xO_;��d�OF���O �]��U�	��"ٜ���'6s ��p#%[��'m��'��'l�i��aá���Aa�/�ʴ�i�z�Ĺ<���?�����  -�'t{�a��J@	4*�� )�>P���'��'��'�i>�I?l�1��Ņ�+1(�E��a��E�>��?����D��v$�H$>9�%��eU��@k�XL��*�6�M�������4����%����Q�hRp�
�m!��[��M���D�O�@Pd��|����?)��&έQP*����j���Z�"N�����'��py���z<���'`ب��N��[�|5���i��	�D��<�ܴ]���<��9����
f�F:���X5��� 6���'��g��7�r�~"���.���h�<Ը��2%�Z�&��4�M{�!ZAX���';2=O��f+�4�k�]~�!ŉ5X��Bi�`�֪?���'_�'�TZ>}�O6��9c恼#!�h8��a���
#|�h�d�O �$�}@b�S��>a�-Db���څ���ef�����i&1O�d��A�[���|��ǟ��a���]�|�
e��;wL��Ӓ���M��'��}:Оx�O�B�|Zw3|e�R퐾Av���J�4oU��OR$� ��O�˓�?!���?1/O�Ƞp��X�Ɉ��#%<t	�t���x0$���I�����py��'���2g�E��^d�\�ř�W7��d�'��	ڟ|����p�'���s�-`>U�w�7=W:H@�ˍ<a֊�a�)r�~˓�?).O|���O��$fg�d�o����� ���î1|[��o�ԟ$�IڟT�I_y�̉��ꧺ?��GO�MQvqoL$_����
͒F2���'2�I��0�����J��v����c?��X<}�>�;� �;5��bK���ӟ��'���B�~
��?���j������aR�=�gd�`�0h�S�������6?\��Iq�IXZ�I�)Z$h���� iL�zqRߦ1�'�~x@c&tӂ���O&���<�֧ug�T*m�<9����1&B�1��"�MC��?�4K�<��?���ԸO��A��K��-0���˚#� ��ݴH	��r��iX2�'���O�ꓵ�MX,�X���JG�RV�
�l�6�nڷD�>���X�'b�D����%$Lx�RY%JE��k.t�ynZϟ �	韌� �����<���~��;�ux�� �����n���Mk��?�����L�S���'"�'e�4R�,�4裶H�0K�v �FldӐ���R���'��I����'�Zc� @e����X +-��[�O舫�4OT���Or�D�O�d�<��	ʦ(�2�"rf�T��a�@��V�hJ�\���'��[���I˟4�I\7�Q	 �
�<�['A	�(B���r���'62�'F�R��Jw.�����A`$P��Lz�ʼ�B@�MS*O ���<Y���?��J���$&z)��с�Ԕ�s�Z�!�t� �S����ٟH�IQy2�g�q"����D`ӌ��җ���b� JN�K�4�?a*O�D�OF�d����x?YF�Y;O_����P@�Zh0���e��ڟ�'}0U�Q½~r��?)��n��SC��=�������rY�@�	��d��Y@l�IFy2�'_�IڀV��LC����
�9�|���Z��S���6�MC��?I���X��,)gd�r��H5t3r���6N�<6��O4��<^�D�O����O�F��m�/n����Uf[�Ci���شi
�:�i?R�'�2�O�����DZ�R\:y�5%J����h^��llZ
}L�Xy�'���ĕ�+eE��(X<|��)�l�V�.�oZ�$�	��!Oֻ��$�<Q��~�"��ڐ��/A
w��
4#��M����D
��?A������I�"ظ6Z)<�ڀǁ4]��,*ش�?IdF�>��`y��'o�����*� ԑ�Ay��u2#g}y��L��1��?����?Y��?�+O�� c��_��-`��YZvh;�j\*=1V��'|�����'}��'��A66%$����K=t)pZ�jW�D74ᰛ'k��'���'�V�Xytѷ����$�Nxz��Ǧ�,�se���M�,O��ľ<����?���2�8�O��(3�&l% I��	��Q���ܴ�?���?9���D�=�t��O�Zc�T���Z�(��@a�k�پ��4�?Q+O����Oj���%$"�|nZii��b2N[�vi�Z��C)y7��O���<��kǴ@{�؟��	�?��3��A�<���f������%�����O����O�"�;O���?��O���: X!r<�Z�h�3H����4��dΏkRrLn���	៬�S0����~Ij�BP4��)�����
����?I�]i�q̓�?q+O0�>A��뜥m�,�	�A��#z�����LC�mLŦ���ʟ<�	�?m��OFʓ@�1���N�!-�z�S�S*ر�i9���OJ˓��O�
6v������p!KX��7-�O,��OT0Ks}�Y�,�I\?!���]N��X��\����K�ʦ�$�S�u��'�?������� �AN̽��Z.ǚ�YPj>�M����|T�S���'V"U���i�m��%s�L�K�%�3 ���A#�j�D�d�rW�<)���?a����](x��["NU%c�y�W��6TzQAn}}�]�p�	ny��'���'9�0iև��~	�� �%cr���Cۻ�yb�'�B�'!R�'��I�F�vP˞O�d��'�,m?�P˷�]��۴���O���?���?!� ��<��� �)4��7S�(x*&nT��4Ѵi���'�b�'#�PJ>���V���;-nk3G��$��U� *t�Tn����'���'���	�y"�'H�dQ�S"�|S`$�<ʎ�c�L$/����'�W�|:Uٓ��)�OZ����n��d��s���⁗4+�p��Ma}��'�R�'r���'u��':�֟az�l�3o�l�1�ϭC�����i��	�"l��ݴ�?1���?A�'l��i��YB'�6�&�F���@Ejc�����O�;&:OXm�Oo�IU�l����p�X�*���p�߳@ݛ��Y�R�h7��OL��O ���m}�R���WiA�g����`Z�f�vЊ��Ǣ�M{hz~b[������\ϖ�٧�׊�v�`�A6I�N����i���'"dǷ6�2ꓙ�d�O<�	?|%"�Q�`�
\u����pIi׿i$�P���P�|��'�?�����B>�:H�*��Z���Q�����M��%���Qb[�8�'+�U�<�i��9���"�>���d�-���D̸>ɣ��<A���?����?�����$i-��ѡݟY�2wʋ2;�����"�a��֟��	n�֟���j~����(��v�
s�LQ&�;U����'Pb�'��O-0ZƂt>5�e��0�����h�rH���/���Oz�O���On��`�OjQ��^;~R�}9��X�$��`%XR}��'�R�'��I(JX\xI|��._��٨�	9,���$�UG�V�'��'�B�'4���}�.��n`�E2�lÑp�V �󮚛�Mc��?1*O&x:H�w���,���n��9�,�6~���`�@:��N<����?Yg,�<�N>�O^��s�J��.�y��Y .'Ę�4��� �3�v}m ��	�O<�iW~2'E��tٲE�y7��{1� ��MC��?q �_�<�H>9��TO��t��m�4;:���D-�M+ӭ[Eu��'f�'}�$�.��O8x���H���׵;�]7�7�ޙJ��d4��(��̟H,/T�����:[��`4.�,CB�o��t��ោ��n� ��'@"�OnP���p�xp�`�@6Y#e�9w�J�OV���O��dY.'�\�S���:3���PA�+ F�ho�ʟ�I����ē�?a�����C���vM\R"��~��\�".g}E�0�y�W����ş��I_y¥�*�j�VÊn}�$pG�E8Nx����6��˟�%�T��˟�q��t�f��Fʖ6�Б�p�](K-�b���	����	zyBh�4wI*�ӈ0w��I6�����S�\7D�O���&�D�O��dɎ%�d��Α�J=�#�P�O�mi7��3D���'���'Q2\���l��ħPϼ ��=.=2�)�J�K��T���i�Ҕ|��'��×� �B�>��ʫ8����E�_H��B���	㟤�'��5��5������+��f	O�;�ej"'�"Kܨu�'y�'�J�g�O����VrQ36N�z�,q����)��6m�<y���{�FI�~������ta��M�J��x�$��
?�h��Am�2���O��PF�O0�OF�>��vK_
�)Qu�%����Ӌl�"t�@���I���I�?�HN<�'@�zE�����QFe�Ӄ��kE.0A!U� �	[�Ş�?a�oX�����%�%PV&�9���qb���'��'�~�Ȱ ,�4�l�'���i��׍0�r��'�B�Y$�Aڴ��'w������OL��O�*2�����[�2h×.�	v'��l�џ<��S����|r���_OgA��L�^��TKſ	#��Y��Isy��'
B�'�"�'fJ���,�zQ"u����?���vNA���	͟���<'���a?A3.ȆX�6�����6L�.a2��Xڦ�"�$?A���?������=zX�ͧ^�2�����J�� +;pܘ��'�R�'R����1��S�?ծq�b(/j��x���I�>��?���?���?�k	5��鲟ؒs�
^��9� �#f�� ���L��5���ON˓{~��$�4�aN߂ Ā�A�6᦬�mjӈ���OJ� ��p����'��dO�
J���e�C�R�Ԝ��ưA$�Oj���O�IB��I
�B�BL����P�c`�ѦE�'�~�R����꧓?���Y%�	,��%�ŉ�;~>L���>e�6��O:���V%���}���#_g
 ���EG�uM\Цq���Ο��I`y��O)2�'��I/F�~����46$J�%.@�O6��)�ޟ����NN�#b-ȇX��i见ݦ�M[��?٘'6����x�Oz�'�:գ3%*H���R.e�
iQ�#�	.��c�����H���\u
8����QO�q������A�ش�?��1��F���'^�'��B�9T�#�.L080YD"�ݞ#g�	ڟl�I�Ĕ'�<�)W�RPgq�Ҹ&�0Q2ILr�*O��D�OZ�O��d�O�-#��
�l�S*U�� ��.W�1O�D�Oj��<�R(���)A2Έ5p6�E��@h� ��	��IA�I���ܴ�2�D�ӨÃ�z��!�s�ZQ�']2�'"�Z�4Z�"Y��ħQ��ۇ*�$]�>@a LB:$;�8���i���|2�'��ˉ��'q� [BN�
��@E�C* �;�4�?�����$�:rP %>��I�?A[���nk�8����;Kg�iۀ�����?���tN�QGx��� ��)��z�~ YG��Œ5W���	�s�l������	�� �SRyZwQ��vm�v��cQ$�-?���ڴ�?Q(O�S�)��}�J� �j�F]z'�mL�vJQ:<X7��O��$�O.���k����؃�!��������әw�����CX9��?I�^�|��ʇv��c/�,d��=Kq�i��'w���#g�c�d�Ip?��ŀ�_�yX#��1�� �(�T؞��ß���IDn�B�G�I���Q+�fDJi��4�?�s�M��'��'�ɧ5�Z�EHUɋ9`���"�ٷy�R�*��$�<���?����򄚑Gڪ����.H��h�3M!~Q���_��x�Io���|�	�?���fB��F����A`�>��4�*hc��ӧ���+~��T����'Q]yE��-d�⭊'�3�=�ȓ8G A�Ī�0qB�W0>@��"e#�I� �@���ΓL(������b����"���li� (_��5P�Y��"͓'(��6$P�R�J\i�J��'O� �2k�<�P��T�"��-R�/��L�pV��&�J� 2D)W��A�a6pw� �a.
.�x���OY�cQ����@��&��@)Q�@�c������5$���>m��"�&�[j��,����Ob��ֆK��n! �\�m�]#�۴���]>�1���?_(蛖�J�h�cQ�>}2�� ��Q���^��ڝ���˝O�.�B`��DI�>c��a[��o�������|���'�(5j��?Q����O��
��N�WZ�1�ѾX���S�"O�IAָ�c⌕6}Ђ���h��poaxr�%ғ2��{�ÎOJE�
�#g�I3Q�\����T�Q*_0t�}��ğ�I��]�j7����L�"8sB��b��M�u!��z����O|8�E��w�1��'9,P�ȩ�����@wif-�L,s#��O�a�������p���{���+'BbS�B�
�������D^� /�Oў�Z2��v岉S�����ݻwo8D����A�d��t��*��e��K"?1�)
.Op8Z2<
�ȵb�")�)�@ �,I�v7��OX���O��dܺ+��?��O����wo�/fY6,aՇ�1zf���nD�N��}�cǀd0�`��'�4��� O��f�:&i� �#銨`.��ShR8Q�$�R�'g(����E�u�����MP ��Hɨ�?����hO�⟜8@�M($��‽)r*8Y1�,D�����!c�: 0AbL�8�p���+���d�<�� ϕ�	�����T1jCn%����4v���s�G�T�IŊ�	����'B,��h��+E�J��`��"�M��m�A�6��iL2*L!�OUN8���7#��01�dY�#���k���q��ؐ���lti��&O��:�'Q�^�l"���@m�i� s�:��/$�IA�����8s�D��Q�ȧ^|`0j��#� �ݴDĆ��&�3yF�$��3BM��͓��D��5�'��\>q���L� �֭���\p��Fŕq�l��Lğ8�	��`��
*����ū(�?�OG哆pJ��
#�6��	Sd�H�K0��'<�5ZU�-� ��h1k�>�JPj�.b�jdC���#ydx[Wj5}�&M��?a���h�n���*K�*�1�g]���3�A�D�!�dQ�Ss�beg��P󢀫��@U�ax�/ғ`�ld8�D+x
��҂��y��Y9�V����џ\��O6L�2��	�������]/[�iW#D���u+�!���q�C��fe��i��W�srl8o�g��#:F���E?M��� C��Ƚ��ד O�<rG�׌ [�}��I0�I≴VO������4CYXʥ�٬a�2�1ݴ+�副T���4����:�	W�|@E�
�}Z��'",�C�	Cg�H�%u¦`�c՚B�T�C����O
�O8��4���3 �鳪G?O�4*���<"8���?����?���6�$�O�����0L�v�/o�j@�d%�� zQ�ge�]�~�FY�ZT�hN�RV8��Cȓ��`�fƅ��>�+T��%�����c�,���µ]�bIQdM�5
\�@���'�B�6��O��d!��1i�p�Y@BԋKb���a�6Cq��#�ēJ��u͓��x��y:ׁV:I]J��HB�)�/O&��_}b[�8B"���M���?y��^����(q���1�����1�?I��N�Jhy��?�O�|x����'/^C*��w�&(�g�΅&v^���9,B�P
1@|�;S�4�\�p9OF�U�'0�X�����O'�H �GTM(2I�c`w�<��Ɵ��?E�d��+
B<�`F�G����6��C(<I��ik)�.P�1�*T �EB�2Z�Y��'�ў"~�)�D�(������BM��(W�<qWI�7qe��MΧ�X��/_W�<)2�T��,�8�
�E2����GL_�<��L�q:��ҕ!�z�Qwc�Q�<� ��ARCD�$�h���ބI~�!0�"O ��7��+
}�҇�Jy΍0�"ONHC�GV�e���;�Ϲ2��xj�"O6���d�0m��eB7w�n��@"O�(H�$�F$h����պ�"O���p��[�&�i�DѬV���"O���B�ZR�bq��Y?r=@�"O����L�BT�+t�Ȱo�D���"O��[d�ПE�)�S,	�O�.�(A"O\:��Nk�!�a��I�H��0"O�����D:�!��¯k~��p"O�4 a�33Z�W�7ndu�"O~��4���< ��+�`��mx�"OV����5bN�]iAd�z~pi��"O<8Y	c���C�� ����"O���7���J�zCI�7�"%�"OԲA�ǓEP�bAB�	hȺ8g"O#$�P�q@p-�TaL|9;�"O�A8���qh2�O.Az�qw"O���q�^�#mh z%� aԠJ�"O����J,41�K�lW�v���'"OD�8q��7�h,Ɉn��sp"O�՛��F�Y�x)�e�եt��;7"O��r�L�0�T����t[`D d"Od����N?i��A�U5-' ���"O
�x�c����"�%\6$�@�t"O�9$��L�fU���ɖ:���a�"O�M�'�'�M{ƀ���H��U"O�݈5,ߜ++go��m�ȅ��"OҸ�L�T�����-8~$�sQ"O(�3gP/�"�P�o�3,iT$��"O��1`Aut�ܩ��1BH5�F"O�P8�僕z^.qA��*(���"O�X�c�`�,U(c Q���c"O�)�q���0=��`���^��-9�"O�Q���u֩�4!Mwc �"O򧠆�	fp��"�^�~Tz�"OL[��,R�L�1��kjL��"Of4���W�P��=Q�Q����"O�k0C!�r��
�W��1�"OVX����^|B9��M��b��!A	�'P<[uT$�X&Hק �qj�):D�(ᶏ� �N��r��j(�rB3D����+U1<�j�@�Чae@ sĩ=D�,����9�TEP�kY��J�:D���Ď�3W��0[����T�T 6D�4��W9"0�Jrퟍz����	3D�����A�!l��r�]��4ԨF�2ړN7h]#P�6<�n��5�>n�	�w��%?�fC�ɵn��(A�B0�f�^�5$,��G�L7h�R�{���F8}堸���I|U�/\��C�	?p����N�pƔ�.�a���	n�X�"lOh�t ڋ$�V�c%�܇�D����'�T͐D�WӦ�yAF	�	#��1IȜz��R�5D���DIۇR�&\��J���1O.�FzR듊(���1�k�#~n�4����y�/�1|(qR��K76d��C߷�y"�P�[������G�Iւ��ā�(�y�J<)Z���$�	R���ªL��y��	����M�w�-�w��5�yr�\��$�ˇL��ZS�lI  �y�CҽJ���s΁.IO��'$ޕ�yb��#��%Y�JS��Ri���y�/��a��aZ�ؘ4����5�y
� �-��KÆP!��f$"��l"O6��e i���dɃb���6"O���U�ANdZ'��V� �3"OTIC0�H8` ,p3�٦0��y�"O��Y0 C[{��' �5��=��"O,)yCȘ�X_��#6�4%��)��"OR�◭ۺ�a �B�"N���"O�(�t��8���($�QlҀ"O�Y��^�*���!� �R�"O�Ur�(��B��T���L�f�'�R�����4i��3ǀ�%=�L����P�!��^���a�PK�n�"��'�pt����3Op\��Bϝ u�i��Z	^�!�*Az����ص>^0!9�!�V��O$�ZB*4O^(��nΣk4x�;&�)��@pO���R��Z~K�J8���#��z\�qOjM:T�̭=]R0:�C� .Y��צGm���S%a}"�S���'O`b��7D�y�<�P�Y4Z2.�HG�;D����-�j��9+si���>̙��y��1�&��6�V9+ۓ|�D�D�Q80�bP��ą��*���N�{�d�۴Q���N۱0S2UZ�/Bl�.q�ȓm�40�"N���W���V���<Qע��R���VM1+��>Y!D�B�/�� 1���$`EI)�.?D�к0d�V�#
yF��Q�k�; @Fh�����YS>�_�%B�bՍ��<a4N��}U䌆ȓ
 u��Z2G�`0�Q�H��Y��Q5�3T�a{���g1���G � �̴9��ބ�0=a Cmn�<��o�)@|�V��"��eS����Q��k���y���-�)�1�\�yef�SgI�Ә'mv,��gH�W���r�.9ҧc*,��ϙ�+��]�ĆW/���ȓm`� &�Ҧq�:��%$�7�Rh� dz8MZW_��!B2�g~�M�np.<�SL�
+4
h�/�:�y"B�y�d���!VR�nl� j�#\�0���H��Yr�`�'lOzLI��/BQ����K)\\�r�'�H������t��Uck������ 1u� *�3t�a)�"O�5#	�9U�pX
R�o`\���S� gp|�V��X;��D���9�8H���IqR���c��y2��d��Q�D��F����)��+��	FK�O�|�J�d�D��O~�1������S�۩Y��3R"O�%��$�2U"}� n�)�X�
G�	3�%��� �퉴.6�B@��x�"��SO�%l�B�1;r������ �0�7����C䉷1
!B��NH �냀B�J��C�ɏw#tq�`�~��x�0(��
�HC�	�p54��t$T�7\�����'C�C�	6~��%��JS���X	����'�ЈIPc�:�(�)�
�0}A�'�Rxre��/>r@��*�=z��R�'�f���G��ؠ!ᄥ
1�%��'�R�xB�6z�)���1P�0<j'/�L�����P
]��y2Ĥ,#��ɣ������Į^��&ᅦ�\�ȓvF��lM�FSn͊V�@��Ή�+~��c��2a�ƌx��
��?)��8����1E�=�c�ˏ2<z�"&�'�ݲ#�'}r�ْ�(�BGa֍b&�����3I��)�4h(͸��?:H��9�����%�d�='��`2(���8Mۀ�O�z4��q�fP,fBY�ɶ	���G��a����0�U8u�֔a�'��KT��"�/N�L��kLۦ��h���V���a���O�E�D!��rx����z&�qa�"\O���U)���̍��4*N��Cw�:Ų�Ð�U|\6�Щ4�,PJ�#O5����c@%��<�w)�d��u��H��O|a���΅��܈�M�LChPgb��- /��д��D�q.f	�U
ӓ��Hq�i�	�$��N?I�'�T��LT�fr��QD��A߮]*��O��#�ŉ�HM����}�Ԕ?UAql��<��0`�p�$[�v7-â1�A��,gQ�D���4F�˞w�>�[g�˟_�|���"L����C�5������]����]�L��OL�p�]	4����[�|iZ��	CʔB���7SlHw�+��.[�  �{m����`�o��(@�^ɲӎ	����"B�s�����S�? Ρˡ���A#v�1��S)e��;$��X�
)Y�j�Z�'J(���1������un���p�W�f9Ĕ�Fɜn��Y��K;KW~$kK]�*�x�J��V$��2](������"�#9� tt�0b��J��M�'�X��)U� �}�"�[`q�%C��6\�9"�J�	59*��w���W�bu�caj�Ő%E[;naA�㔺\��x�ݪoŎ�Y�@L���)�c��ƭ�R�ȹ�ą��x� 24�Oލ�*%�	�2�.�B�L���� �JX�F)�tQ�5�D@ށJ��E���tU�T��>nT�sEI69/���OdQ�r�S�
1O>�b�лDhp���	��@����G	�G���3(����p�g��vM�"H�5�8Ӏ� ]y2ܙF4�vH+�i�5Մ�m���r��L�����.Ғ� ��3ǌ��'>��3�6r�nU�����ji�شY���D*�=h:)R��Z�gJ�R� @�p�$=˔)�w)<}B�D7��(Q��B�'��P�P��$�1،0i� K�M .����N-B"Q������ �B+O���@# �Q1j�S�-����Ƹ���%`� �R�k?~D�+�^�g7<P ��5=���Oԟr@�4yr�3��S�E� �Q�cu�)�CM<Z�8�R$*�9T�ȉ|A�Ƨ�O?7m�4/-�-9�,��`��y6+Ô6��I���+O��I�)ȌL����;:(@<�G���p������T�|���O�)hB�I��J'��W�,OV4;�F�o�P�z��^=~5��N�h�,P�&���'TƬ�#J
�z���`�)נx�ܴU9ĉ@�Rqu|��ł�(-)v,��@���iU��9��'�hQ��?��Жjײ^�5�,O��!b֫(f���P�Z��2�=b�f��f��!=� ĩa��բE(ܜ7�L0��Py�O?����"��W�+f!ȍ+�:��-=��x{a)�"���ڵ
��0<4m#_���1v�H�
��-x�g4S��C����>����m�9+��mæ`�,B������x�43�`�K����r�'�Mau�E����i׿s�Ub�g�(7\6��C�O.E��$K6���p�m�-}z�dǟ{�u"wg�J?!�+��M�4�]/�.ݳ�b��}�vPƧRG�!��"]� �Bc��`X (�X���%�:9�a"�)�'}��Ѭ��J���0#y�A��~I$�[ū�wqX��%k�8�
M$����c�2<�ay��(���@����tT]�e�E��xB�, n8H�O��h��M�KӞO21���'$��p&Ζ5V�pȇ�K�ةH�j D�����\(5T^ģ����1qUA+D�h)����~yi�aa	KIh��(D��b�#++�8;THX�����D#D�4r�Q&E[
�s��V<dk�Mb1$4D� �q-�!�쁰�:'6n-��)3D��x��M�k����)ݘSL��%�/D���cX��6�f�=u�,�c�a;D�x
wh�,���D�Q!�b�i7D��R�LF8^܆t�gdđ_+�q��)6D����Φ��ف!���/�U��J5D��IS�:^G�Lka����N-B1,8D�$��͊7T�Q)�%�� 񺥮1D��je���?
��c�H#|6mKT�+D� ��-�8
(���a!��q�eH%,?D�81ԃ�ʸɅ�,8��9$n/D���D�ґyb2Q;�b�wV��b&k+D�|BHӇ=�lJ5�F"d����37D���n��K]ތ���<0�����3D��ڀM�-%�� Hת��~G��u�0D��( *�a���[��#��k�c0D�� ��ڃ^+R��L�[y��y� ;D�,R��x/VP1���}N���#4D�ɣ/�>�����c�j A�(/D��i�F�)R��4+�E�->�N���-D���.L�\�x�fX54�J��)D�XR,"%FPyf�/ p`��)D����Ŝ�$dˁ��FF��-'D����k�JJ�e�FA�USv��1D#D�S���`A��P��!eur���,D����q�ЕO]�B�S3�*D����ܐx�8�S!�Z+���*�'D�x��g�n�y��)ׇ(ޘ2n7D�ܡ֌L�zN ���_���j9D�$�f���Dz���r�؊~����5D�� J��B�\ @ �K	�K>���7"O@`��E�Bp�Hz���T*"�[w"O>��$dK /�����dD�/�H"O6x��.	*z��QH��H��Ia�"Ob���]C��6I=/�F�k$D��PЁ�1S�0�*�^&,�-���$D���S�3^^��b��']�4LB��>D�d����:���x4�C�*�p�z7�:D�<{���=	�+�}�8{9D��	'GA�,<��'� j�9D�PjN��G�Z�j�+�8~¦R�9D��dV���� �!�x���6D�أ���-&E�R���4M�(*r�4D����C٨/ ��`1�"�bp��1D�<�2��"2����E�?�(�1C:D��#
�<9�x�S��i�JX�e�+D�t���@��, �Q�Le��z�*D���Ug � 3j�`t!ҥ��d�-6D��
�@��:��=2��Ψ�����g'D�8���Z�Nq3���1|�N�0�(D������(L(�t�iʲ: L�
�e(D�x"ga�9F��a7%��J�.qA�"*D�T"ޥ@��9�3��a���&D���D��g��T�:�!f�$D��(T�Y��� �%�_��,@Ä/D�d�i�(P�z!)sI��� ��h3D�X�T@�*���D�Y(Wm����<D�4�u���Y$B�
&�|���h7D�T�!h�/�,ەi\B[�AUO"D��#�'�+/�6�kao�#��ewd:D�D:�E�!�rآG�új��0`�#D��@n��J���ÿz��	��#D����-�+|� D���0Cx�21A!D��b��7CdpAK��JT}97�+D��Y���7@�ɣ�+�lH2	x�e)D�\��A=pyT���T:?�1��(D��ga�P��f�Q67+��H�#D�$�P���b���hr/�;		�hb�"D����Ň1I�����:�
=�"D�"��FC`�u(Cj_,U}�(© D��
WkNW���3ś,"Y8D#b�?D�P8%��&�=z����B����<D�T����*�0�z���7]�0�-D�Xk�"ۻq�Rmy��R>����� %D�,� �j{�Ѷ�2ZGR�%D�D���,
A��F��9��B'B�hO?�$�A�2�Yd��cEt�d ��!���$�\
�PS�G�u��C"Obe��,� �5���%��`"O���V#�(v	,��#�M#�ViQ"O�`Qg��/V�,�ǃ����"Oj�[�nߙ3� �b�A�����Id�O="c7��>��	���&+*�3��OF�s0D\0w�L%2W
}N���"O��9F���u�̉Rꀠ!�hI�b"Ol����<\%p`��
�&�!��"O�a;!���v-��V���0J"OV1Y�σl�Bȓ��
�6/P؊C"O&�0v,Õs��TbK�0-��""O��pr��8r#�Ʀ[*�	�"O�Mٶ�$��ce/	�?Yf)
r"O�p���%1��㔨J��`��"O�U�ð+m�I#W�Z�jq`�:1"O�U '���pz�&0l<��V"O� ��2��B��hR���et���"O���=L��0� �46�ҙ�@"OD�i��6���]�+v:UiB"O�q�lS1MJ�����,W|�Y�"Oxa�dY�pd������86e�7"OX-��Hڹ+`,��/�� �"O�(�tSq��\s!���)��"O:����M�,H�@e����3"Oh��c�f��ӊ�_y\�2"O���tm�p2T��ë�"W�(�g"O� ����?g{�ț�� �T�"O�K��(���q�Z�Hɪ��S"O� q�HMh_�����m��XӦ"OdY�lT=//�4#w�I�g�0�1�"O���P-�/tŉ��]���ae"O�0'*G�>��P�?w��	+T"O\K4�+	6�@�ϐ�>��y�"OT<*a��=8xHz���/u�r`��"O���\)5�����!����"O�i���5$�l��/��LPg�'��'�y�@����p���{�l\�
�':��V��ndh�"�	�#7v%�
�'��c ��1DwjL��-!X,L�	�'p�Y����p�|1"� ��n7��9�'��d3ΐ�5�hă���7���+�'����R7|z��c��.y�s�'i�1sv��;�P���.�)�';4���GT�1�.�R�A�E�$d��'�(���0oX���B�<D&�\�	�'��atM�����Ã6ö�1	�'VJ�����\f��b�#?/=֙��'��|����)�j������7Հ8x�'t1��J7.����Y�*�>�)�'�&E#P�ƙL����Mה/ֲ �'/��ucr��ꑈR�&��(s
�',�3DH�0^lکсL�,T��
듡�I�}wBL)�dJ�)o(t����xB剟%uU�t��ó&کa}!�$�a���IQ����j}jĢ�
�!�d�3b�`p�B��&-�ܐ����n�!��/8��:#B ��$E�!+�!�9D��HQ��@}�Ȗi�g�!���J��ځA�+`8i��NV!���*3�\���3|D\m�֯V`!�D��k�>���L�Y`�1q��^�9\!�D���s�kNOA��F�^8y�!��<b*��	@C 4����)]!!�d!G�,l�!n]���H�k��]!��A��B֭5~����IT�P�!򄎟J@C�Z�z�H3�K(zKQ��E�$@22�� )$��/��@�dˌ�yR��1.��mW�|���ٹ�y��K�/C^�YR̅/V�B��ꃒ�y�hT�����LB�O@��R�:�y2ǌ�tX�c@R�: y)A#��y"�Z�{\8x��X�7z9"@�K �O<�=�O�.����%>�`�¥&v��i�'ܸ�9�ŋU�2Uab%f���'�8��R-�����XI- �)�'�l�9`*��r��(p	�u�\e[�'y�]��DW/��ˇd ;n@��'l�\����h�.�q�AW+��TY�'+|tA'�7h�"�����pZ�'�@�R�P.����������� 2,H�o��n�{���-����"O~!3ՅVNF�0���)&*l��B"O����E�hnPm���F&5��"O��b	DL���hKH�#Xq("O�ݘ$ J�z0B�䄌C��C"O�y�b&�	Ԕ��0� �f�X!S�"O���4�>�H�b%�R90�E�"OM��B3�t`�O��
��h�6"O��H��8�x8
�+F�H/�\��"Oܔ�T�I,��0h�i�4�0��"OH,��
�'3��b����1�"OpM�����8�"O�+��|��"O(���Ae�<-(�װb�\�A�"O�i��*dA ���Y��(�`"On�z����BIT?�4����~"�)�'�,�-�DC�%����sf���W��	ʤhc�\ Qf�z%���B
X0��hW�p�h�1��̫�l�ȓ%�(�JSE���)DHӥJq^���F�܄٦˰v�4y�BG� �D�ȓ>0��$K�1�x�4�N� �ȓo��h�9��+L�E=D�h��!I����RC��I�i�� D���$�xX�$9e���x�[`,=D��j�"_�| ��) ���6��d���:D�,�bIB2��!��oH^��p�+D������C��A�m\.zFB Q��5D���"�Ƴ B�;a/��e�J�C�
4D���@�Z���2�'�.0�l0D�
�	P�'.4H`F
L\���`3D�8[f��9$�ػ� 
�%;�9	t�4D���vG԰~a����	P�yt�?D�(L�DW�Y+�e�I!<@QF�;D�<����[��RU�֣9�b%?D��!ꁁ[3>E{T+ѷ_����':D�����?OYh�M��Ac`	�@�#D��X��	�.<b`�t�	��,a� �!D� �6��A��kΜ?a�*��9D��QqNA)%*�!�F��`�4dQ-6D��	�jX9 l��8CD��X��"8D��jB-�[�8q;֫*Y�꽳�m"D�h@2o���|�x����*����� D�0��N>�,=X`i��
3���D:D����K�a���G&K�M'�񋠬6D���LځIHV��`ɒ]Z� 5G?D���Ή�F���:(<Ai5%?D��9�"�lF\�p���4���J>D�x�d�#7��#�0*����c1D����)�d��� �e���0D�����˓�40�7 �;��z�//D�T��$Ҿ	�ABе&�| Db9D�d�G
ff)1%J�ΐ�9D���DiJȪ�(D0 ����4D��Z���++ܠ����Î����.D�<�CΞ�v z!���j���K!D� #�>M{��+���� jH���n;D��c��]�xIH�[����,��Q�,D�D��..Jd�P�2PX3po?D��+� bv|%�PiC ���E�7D��@��%H�XD� 8{\��Jsm4D���s��#U�B��/˝c(R�XF5D�8�tO?`֐��(^nZD��.D������sh�i(J�1-����c:D��#G�L:��ac�
	f�
��9D�� D������ON~��ɍNs�(
P"Or5��I4p���βB�n�E"O>���$�/G���΀\f�,��"O~3f��6B�(�a�L)b�*O����M� �� ���,�Q�'��T���9ij ��e�2J���B�hPN�}���kC�$+�DC�	&[D�qu��K�\��1l�+KzB��X��=%>���s�lʮ�ZB�I�+�~��u?(X�q�"݆<��B�I�[{��󃈙y,��T$ۙ61�B�7<N�ұȃ��=�&˃n
�B�ɲ546�J̸ׂ"��A��׌9�DB�	�8Q�=�Q"W:C}b�p��B
K�2B�I�&X��L
R9y$$�	TBC��7~DHi�`���6�S'V/_6C�I;D���R��̩M+��R��S8/��B�	1@;������-lZ�8U
�>btB�	�� ���;}AP9�&K�W�nB�	~;$`�M�v(\�AP˼n�FB�	�0�A$B�&S�D �FΖ2
��C��,$%�%�QNZc��P�D�Qq�B�	C�� '�wc���d���B�	��8����B�NY�B`6D�Pk���q���Q֭Ŋ��(yf�2D���%`��\��8�f��9ܪT9C%<D�B�B�5(�x�lG|z
=D�\)AC!$|�E��Ԇ7�m���/D����H#u�����O��p�왵D/D�Л�BC34��ɫs�ڿ|�d��2D�� ��O�/ł���&�(�4͹��0D�<���Y;_��̻b�U�9� /D� �A!���M^6*�
�a�,D��[��U��I	��<?����7�)D�����
&ZcR}A��Z.�D��L-D�9��K�0��cf�/Ԅ%�@,D�d)�C����$�A�P�l%Q�=D���N�J#�[�j_�ux%q`+9D��V�R;B�:Փ��b&�ɚ6D�$�T@\�9����p��a�d5h$�&D��W���-=�ePӅ
-���!�8D���˜�]���w�͚4��� �)D��X2$�!����
g���n(D�d��O�z���ׅ�1P}2t;#&D���Ġ��3�j�@��@�����#6D�`Jb▏~�&�R0��3m`�}�@5D�H�P���L�x�
R>�i�co-D���'%G.!��A�󫆊���ڄ�,D�Шף3Q	��FD;W	�����(D�(�Ï?#��\�F㖽7��qF9D���@��~p�̨�
�2P���`7D�,Ge�j0�`��m6�-I��4D�����!�Ub�A�n��qp@2D����bJ�Xq��NL	 bR�P7�-D�l8AJ@3�� ��ɒ}�XUB"i)D�b$�/5�<)y�E�*I�Txנ(D�$!��K>@1�tG�s�P�*R`&D�P�U�A xZh���9P�<�&�(D�T�p΃w�ؼ��)�&|xҘ6�;D��3�HU�s �y�DN<O����f�4D��9CM�K�ɠ!��<�:B�(1D���Ā�~x<Ї�ܿF�$@��h+D����%L=z?��A@�[U<5�wn-D���eӁ&�1�7�_�!��h!�� �В�h�&��A�O�!uLѓQ"Oڌ�� ��8ɶ�^QeLq6"Oxq� $6Ia�N�W��|
�"O�5��K{���pm�M�>��G"O�,(G�èLeN�RQ��+y���"O���倎�G@L�:�	�2 �1"O-Bg�*��0�D��$P����"O��eCQ5��Y��"!��髀"Ol�9���
�ܸ 7�Ⱦ3����"O|��@�Ij�h$E�I�q`!"O����6~��#坦5g�]��"O@�S4�A�[���z�#*P>@c"O�\b��1��yrB�$A_N�1F"O�%;�!&��9&@Zz�V"O�� 7��6��#HY}I�ҥ"O�Q�bk�@�������=2�)�"O�œ�B73t�	/�7*R J�"O q�L��]b����$�*P��5"O�����?	Bh��$�7!޵j�"OX�n&EN�4"`$&&�r"Ob�����(p��Es��#%�`r%"O�x��&Ӭp�^�;U$��l#"OU����/��,��iV$�@)�w"OLt�&���1	�s� >t�ٳ�"OJjsH)/��!PFQ7iv���"Oj4	3e���)x��s�
1A"O�\,�G��bt��,p�$��"O�� �&"��4J
��J܊�"O`�����QMx���D$!|��X1"O\%z�%ɬjL4}JVa�< `@��"O|�[��;Rv��7"EaШ�S"Op�[#K�?X�$�Qbצj:nɁ"O>��4�J�Z��"��"G��]��"OFq�r��=@���cb_�^���9�"O�5��F��")���KՋx��w"O�|p��J�o�t�Q����4�e"O����	7�Cu�W�c*�x��"OF�ÓB�_��!��3y����"O:�!C�K "?T��d�������yB!٩a�bd���� S�I��ώ��y�)�;�|5�Y7�%X���yb�I<>K�u��k{\XQ��y*�
XV�����qM�a��H��y��C6�����n���9��м�y�Y����@�ӋiB$u��V��y��W��(�B�>[�U;7j���yJ�t�h��/�b�.(S��R��y��ܚJB -�CX�Z���k���yj/m�ء��N��{�@B2͓��yr	��E%j�i!��PB"�"�y��Q?Eh2x2�h-R=�Ə��y��=>��+T
�� ���
��y�#�gD5I`(!����j��yr�2f
tP�Jb�PD�ܧ�y������F�D�	.��q�I�8�y2+�!F�c���Q?�A���#�yb �u�V��(	F�J1��Ί��yb��G� I�V��9>��@v ��ya��U\����49�� &@��yr��-z�:�e`�1�I��X$�yiF�
�L�K��|l@S@^<�y¯X}���5`�r;8�˵C<�y�H%v\	��Jȼ?��"��_��y2o��K�("�N�2���q����y
� i3J͜o�n�䥆s����"O�lC�c÷/ ,���G>���F"O�U+��	��tb���$��"O�-� �A�d\���\k� �P"O�]��m˱9�iSȏ�h�:�"O����ڿC�Z��b�Ր9�R|Ѕ"O�X�H�}1�}ss喫.IP!#1"Oxhz&��M���eg]�'.���"O��#@�}Ԉ�f��Y��`@q"O��0�X G���7�W�	�؉
t"O��ψ<H��@L69,�u�T �O�=E�d�\�e����!WBRTk'`�*Ui!��`d�X�2j޾X%¡�a.ۢ�!�s�E
b�En��2���6!�Ğ=%���� "��]�b!)"!�� ��$F�m����`!�$U�b�r��+F&c�f��e��>i!���!d��0-!^���A��q�!��@:�I#�O6$�H�	��'�!�
$ĸ��pe�*��AX��=$�!��^�����&�U��ͻ2�	�=�!����8�;��C4p�C"O�xy��'� ``BU͊1��M��'�Ԁj�mH.󴘱 �Y�f@�	�'�r�6��*e���6kE�L:�'��qz0I�(IE�PV��~��ِ*OR�=E��F�=ot-�g��b��4�&@L:�?�����4��AV(Q�dy^�2���(��؅Ɠ>��@���<Hg��0��zP5)�O~��8�O$�)��/@��z

2�Ա��"O��.�5u�tPS*�
{xY�u"O�T1�a�yf|�QN.PUrЛT"O@˶!A�n+z`�tĄ%.����[�DD{��,5��!�̚�QO��S�/иd��Oȣ=��H�ö&�*�`RA�07Zi��"O��B�*#o����b�s`d�s��'�!�D��O9ށ��'I8��X�E҈vI!��b����Dc��)��p s�_$y�!�$���d�8 @ԃ�:�!�D�* �0�7HZ�|h
�$B�!E��'P���i��X���"
9��LarcP�i�!򤝭/a�IrVf�6�ށk �W!�$z����OP�E�^��$�P�k4!�D��&:AصHf�K�6#!�W��4�+W@�PH	��d۝�!�$Q47c����oޮ*����`��5T�!�� <�i�kӓ3y�0���( !��0q�L�t�:��,�r���=���â#��t�V	ӗX����5a�?z%,C䉴#
�򅋗/j� 9�QB�\RC�	<$��6�	���}R�� �=�B��(p�B� ƣU(jPV�xTbٻ(�C�$QD��a�
-�$PZ�Ř
' :C�	N� }���٬I�����6��=�Ǔ]�& ;���,��u���:>Y��,KPaR�b��0]�zE��0s�8�ȓ.��a�0�%��i���)O�R]�'7a~R(�a9�Y�K ��s��y��M�R��%�Y'Kg���%��y	�8&�؁�1��@�O��yBa�CA*<!b�3z� X��* �yBm�*T!(��f�B�F�( �ք]���xr�h���kf-��An�ܩ�KS%+�!�D�'eD��rB�+fJ4�q�.�B�'Ha~
� \`i!([57����Ձ~v
"OBۖ!�:��!ҍJ�g^(p�a"O���n�?L�5*V�I�N���4"O�+�g��2�B}K��_��C�"O-
��=4�P9j�'I zS�b��'*��R�̳&�ʚ#s��'��o:�O���d�%6�vU�C�Y�=��хb:
��f���Yu��4�ΈJ�L@7 ���G=D�dV�L�T��􇊏*�T���>D�xC�.����G��&�(��?D�(�ŁZ��v�@��&�(	D�!D��if#¾S��4qw���/��P��C%D�8�JT�1k�9@�\�6�x�3a�O(�O���>�3}��4(w^�A���n�,����yBD�=��t���f�(���ҩ�yR�Cc����ʛ�bM(�Q(�1�yR��w&u��K�0�v9k6��9�y�04&�!�Fs��u�M1�yk�hr��Y��9��$�婁��y�(��?�ZQ�	�'7�d�c���?A����c�@`�je�,s�D��Pm��&�$��	 $�d8�5Șm���T"��	\C�	 ejPp�Ҭi���2G�B�ɏS�45��)$v���B�9!�.C��K� R0O5j�:����$]&�C�IxW���W@��O�0�b!�	�[��C�ɞ6��XC�$�4 ���W��&�\C�ɽ}#t�j#Ԋ.�ȕ94 ���$�<�3_ ���`�~�^�C���gB���t�2��#.XE��˶o�Fd���h�D��B�?uh`dYS'I>�%�ȓVO�(+GK�	$- �i�N҃�օG��e-2�����#@��!��@��C��83���x�(��B�8�j&IG�IɄC�	�a�$	�v�)*��k��߁F����e��<�4A�mDDp�AM��[D@���5�$��MB!6����Rp���ƓsP���~���W��F��'�:���P�hZ��ڥ�,����'xa��5M��X��L�&Ur��@�F>���hOq�4�p	��V���ЀD �|����w"O������/�� �C�CZ���Ӧ"O��F�F5��ѫ���!!#x�`"O֙����2!w�C�(
�!A�'���O� ܖ�a��{A�T�E�-]62�' a~��ۆ<��#�X5YL�j0�N��䓏hOq�Z�K�jJc<��`��L��,���D8�S�)�9\1��Ĉ�N���F�\��r�'Y�De��)p� �3���U�x�c"O�·�O�rw�b���j9>�"O��C�EI&�@1�Y:F.�mJC�	���?A�$��k��Ȋ�B��i��K�<�yr��=��1ڀ��P�)����Pybg�c2e�W =^�H"��n�'�a��Id�A:Q�ʤa���,~W���'q( �'_!d��1��`I�>���Z "O�	�F��/c��r��ϑU��h�"OX���L�0m6�CvƝ�>����1�	|�O��DQ�B'J\4�S�	�I�V��	�'=�,��-7�xak�dʈ3��H�	�'C2�2�(Y1��̙7�P-1�l4r
�'�^a6�Y�]�G#��/Ht��	�'�J(A�_��1K'��1p88J�"O��H#'*�uS.�1v*T�@"O� ��2�V�2�dѸF�x�̱*U"Op�s/Z�b���:){����"O���E����fD�
"x�͂�"O��N��A�yf�<�r=�6"O��[�&O�K[4��0Z,<���Q�'d�kg)]�<j�1��ڀn@�;�d7D��R���偠�Y�q�8��r�*D�諃n��k�DBd��&( )*��4D��J�A�	'"Ne;U(T�+��%��4D�􀅠I#g���:5�רlo�Y¶2D�XY�מs�N�"�ɔ;.�iZ��*D��3"-��,�cU�sh29�Ҡ'D�l�db�k���H0?�M�#,3D�,�QlKm�j|�2�P�T�m�rJ1D�|r0G�I��˦)��t��X�Fa$D�|��������K-�x�IAk"D�lɂFH�M����K��<��m!D�$�c�\��H���n8:�d�1 !D�t���	�VA��&����H?D�lk!��B�Q�Չ��"����9D�� ��+������>����1D�X2�J]#�FӇ��4;6<��j1D���@�ߓ)�<��@Vvk6p�d�$D�p��)�UV ��,T?�`JG`8D�Hb�	�	G���W9D<���(D�l閮��C"�){5��I><4J�<D�Xr���Tnx=���Q�/UV��D�;D�d1���'wa���`4��0�8D�X���	&;����@4 ��Ր8D��b�]sd}҆�B6@�*Y@�2D����+S���SA����)��	.D��� 8p�>�����NG��"�+D����c�5\R��B�]>j��  �d+D��Z�¿5�F̺�[+|)�p�p .D���$۰	�zX�Y]oĠ���*D��	q\�'2�M�4���2e�<sp�=D���t��m� �F�_�8S^��5O D���GE��b�A�asw,t��+?D�hA��s�<��Pg@9N����*D�007�֫7�x�)���(}ҥh"%)D���ۥ/b)0ʀH��̢��%D��i�.A���q����\PFE$D���9`�J<�����3�-90$D�Pr���b��ґ�e�za�c�=D�Xz��ު?���{"% ol��0D�y#F�!�����ؑ`S����+D�[�mja�HU�a�0�P�re�B�	�+Fq;�"Õ�,�"d�?&�jB�ɹ?���G�7E=�2�и9�"B��?���#b��H�KT�B�	�|Q8!�4��F�N ��%/f�B�I4X�tU��NKdV���̻f>�B�I�E]�RG�p�Q�%�-DU�B�	jO���%&��n���kxB��m�5�r �uBր��K�6P��C�6F���m\�eR��`��$��"O6�@ҢΛH"�Z�g�Q���f"O��Х�ٯ-~|(
B��
K\�B�$/LO�������,ɑ�'�}v����"OLUp�ײR$��ŖPX~�F"O$�`�D4)�.��u���0I�5P�"O���H�Od}�b#��7;:��"O��W��m!ԅz!c��d�~�1�"O��R��\�D� ��*d|�d�D�'��� ����G>5~q�a�Fs\ŁW"O���!Rj�y��I�"*Z�И0"Oj��6,�2r��HI�)W���"O�	 ���l���[���_����"O����&�����;���c�0XC"OJ}`UJÆ܀���V�JD4�"O��;��� z��`��\'9�`"O�����,���B��]Ҳ��P"O��PEgPx����f�$��ѓ"O>���HҼlh�@�x��h�u"O���#M�6��Y�x�x�+T"O�`�@ޮ~���������"O6e����i~`CqD�D��hR"O`	��eD�L,2$�����H�D2"O*����֤��N6�}#�"Oj)��F������^~�m�r"O���b�4� ���F��BW"Obhdi�-��p;v��w6�P��"O0AZ��8S,�C��;c�2!�j��]���^�-nd0R��BV!��%FS�Q�cA�l���v��G!��$�|�S 
�a-�p;�쓨XJ!��şi_b�E��?'�	��mWO�!��?7�X
��ۭA�$��-�	R�!��E��U@ԂՌl���̆,i�!��%�x��FOZ�	Φغ��� !�Z�=>U3�h��`�HӅ@*!��
)$�D�7ij���p��g��}�(*�MD&LnX��g�I:!HxH�<D�xQ�,�0$��R�ŧa�x�k�l3ړ�0<�ƨ܅����Q	F����͚r�<9H+p�b]��d�:w9`���k�<���&�!��8X�u0���<�&���0}��g��>����b�<Q�E\&�(�FE�cm��3.X]�<�W� �:Bd��� �$}���*Ԍ�}�<�U�M/G��ɉ���r%T�j7'�A�<Y�Ł�{�m����T�\s�Zr�<�c������q�O�W>�a�D�S�<Y�(J>Vj�0��#|�`��L�<���H-Pk@�+E��=�h5�QXO�<�M_�>��D�%[
��I�<��ŝ�pլœQ�$B��fH�<��iV�LAE�W,�	K����h�]�<yv#^5�!е�"%�f�¯�W�<awOHY�D`e�Jy$ہ��Q�<Iv��"��A�-W�:���A�Q�<�%'��~�2�f��z�`a��@TJ�<��
G&h�Hy�6�ك9 FLz/�B�<���҃]���7�?��!z��A�<	��A� hX�R��9bB��)rO�e�<q���`�aa ��b ��u�c�<Qu���L�нP��ҕ(k���eLJ�<iRMB�Bi�� dW7E�d��I�<�w$�r�rG��,��b�&F�<�3C�~��J@�C?#�y��O�����'���Y*@�#�CԞ��D���y?�{���-dT8�J�"��e2R�4!�d##Z��#�5�H2È$!�d��(_2�Ƀ��>��*%�Ѥ;b!�d��Q���r�(�rو��ÔoT!�ۯ?�䵪0R%&�~��2"Oz�uiU#1�di����$Z���u�'K�2O*���B܂M�nqV�7���3��'��)� �%H�+��d����7��ɚU"O0�3EL j��X����2����r"O����v6%��S�1��"O���!�ۈ0�|�0��A +�\�"�"Oz)@�L��A�)C�FH�yt�1D"O�e�0�2cI8Ѹ!,��v1�G�'��i�eN�;tQj���A4hxV�/�O��W����@�=��T�w���Y����"�P����!?��÷�/�"m�ȓ.�LB *O?���u��UF�t�ȓG':y�a��h��D�����.��$ �-xS��B��)r��
�ՇȓF�x�c���o�ڀ��Ň�vhX�ȓ�
�c1���O�d�v�V4~`d��`�'�E
%�#+Ţ�P׶1@ �'h�2�AX�D�.��&L��y�B�)�'��`CU`����%����p�'=����ӟ+G4��	�r�UC�'��q���t��0��oR+l�ҝ��'��q���
Y.N��Ԭ�UC��b�'�xl9���z���"	��؁��'�����Z�"nv�Ps#���}���xb�ݚl�b���H9�2Y!U�H��yb��$���s�eמD����C��	�y�C�U�2��C�"5�v�3r��$�y�S71���s���em1��!���y"F�֌<;p�N�(	�rA���y�&Ыo�h���¦	�<x ؊��'^ў�O<䥺�͋9���&�>�L���'䶩��?]_�dy�OL� M����'>m2jT��NQ�&�'D�M9�'"� Sr-�O^jPu.�),��	�'i���Y\l�۱	Y�����'��!�C�'�Xy�O����'$�I���M<,0Di"!��2�|q��'O��ICR6$@8M!2��+�������'Vax�(wW�5("&�	Y.ٓ҆_�y���;!FP��l�+T�@��e��y����up4x���5JJi�R�[	�yҁ��p3F�L��fs"���y2� �8$!e		ɖ�kr ��yRI۲@� ��c�v���A���x2�՟E>�m�ye6���C��F��?��
���a�F=v��x�b$˝s�:ԅȓ3�R��a��=V��;�G�.C(�ȓf�($�+�l���'�C8��ȓ;�!!2�T�)A�p񎏙(2t���a��J�*Θg�M�钞R�TA�ȓ,�|�f@\�r�l�3ណ7]�xE���2*���A�M�.�:�2��P�"4�x�'�B�'��D�C�S?W��HׯB7<)�E��'�h�F�x��(r���e�l���'�T=P��݂*
P�n��X�Hj
�'��p�l��9�2Q� 芮~Rn��	�'��x &+�k�p�7w�&)	�'�p��VOV�S���E�%�03�'��y�1F�	�8��S�I	�Ll����$�5�5�c	�A�Z��^ǔ-�FT�l��ݟ���*�t��/ہ?���fꋦ/@,C�I�-�<��������1�o}�B��X(]�Ѥ��Zp �+FH.C�I�y�~��wOʡk�Θhŀ�6<"�B�I4Jm�DD�h�<��b�qA�C�P��`:�)��eYI7�A	~����:��t�� ���a���Q�J4P��Μ=E����|��'az"�EXa��:u��_�xQ#���=�D:O�Y�k�ch�2�*��ϐ��ƛ|R�'�az��H�:���O�T�eS��^��yC��-��
H�G}"M�*��y���8U�ɛ�iѶO���[��?��'������k.Z�4GAǪ<������O����p��\,4Ö�5�+R"C�	�?���j�f4�P�k�|�O��$�O����==�0�*0�к`ծ%	1O=.��O���M�Q� ��S�ygԭ�HE=wS!�D^=l���8[",��-�3Rh!�N-|@"&�(f�$U�p+�dE!����*[Ы\�mt1Su+�t��{�'��I G(�z�"
ߺhFiV�B�0B�	|�r�xE#�skތ� "y�.B�	2T���#�I�wD����[z�"�d#��C�Ġ��5A��Y*���B[R�[W� D��0s�(�� 4��/*.����=D����Q�Ud����M�6��}���:D��(�#ۄb�d�C�N��Au:�O��>3�hd�W�V ��C�E���x�ȓw�ӵ��U¬@��B��S1���ȓ\O�C`!�"��
��E� ��؆�6<�Cr
�`�0B�G�mT^�����}3�_�v䞁��Z��1��z�`�'�9h"��1���+K�L���v~BOL*r�����u��H�AͰ�y2�&'�֭���N�l��F�I��䓪?y�����c�F-��*�;d�t������yҩϴ;_(Z�[�b8B%��%�6�y2��Y��Qf��%p\�g&���y��ӸO!T�ጅS�I�\��y��B�UR�2�a#�D=��߬�hO���	�"
�L���3)�QFځ�!�d�=H�DdI-�&7x�I��_��!�0,���L�)�bܨ���XX!�D_8�y�����%����J!�$��\D2,�sh@;7�~�b��@��!����z9��z���Hă�"�!��iv�8*�=<�j�	C�Z��}���K�Ƕ-ˮY�2�4��Ũp$/D�X3B�%�F� ���W���Ħ1D�X��*��p��6T`G�/D�<�u	_�h�W�Vsf��a/(D�8X�h�c�~�Ɂ#U*=`�M$D�Dٲ.C�A��Z�钢|�P�ґ� D���&�;V.\��Ǔ5J�.�!
1|O.b����$�@�����T�,@r��-D�<��d�	Kp0H�l����H /<O�D#��2�x�Q��R�`�t�pK	�� C�ɎX��<���z4%����=yJB�/2�(���n��<ճ2�W��8B�I,*���2d�Ɗ=��8��.עP�8B�6Ir�k�o>�qI��ԑ/n0�=���?灋77Wz|[0��n��F+4�T�Ș;Cб���J.}�M`T��ɟ��'6��4����U���50TsA��7��ȓu�e@�A�!����C�܏\t����Iߊ�
��A���� G�S"6�م�
I��*�.� kp+�����H �@*eDN��}ic�S�5M�`��g�V�Ƞ��r�x�8lԇ�*}��NԈ��
/(0�(� �'
NfP���� | �#��*dD�5+˞�w�d�P�"OJ`b�FD���|���A�\)·"O��J�ѿh��Q�U�;�&���"O.�B���'G�@���� =�ʩ�"O�{W+X㒜��J�O��a�D"O��G�<��R1�M�l� �r�"O�q���Hc�%��@-�c�'�!�D]�1岉8�c�(� 1G��!�DUpyN �c͘�m��E��f�6�!�d�.R<�� �n�L��1:@i!�P� "v�qU��+�ȉ�ƪK�Sf!�Bb���A"�̡_�-0��Й>�!��=u�[�-�K͜,���)w!�DБ:g�!�g���y����@��s?!�$�B"���%�_�|�����	tD!򄋦 d���g%�1.���r �׃�!�-�5�p�O�N\�ҫW"R!��A�.I�I�>*p�|��I��!��6,d�bg�(\����ȃ:O!��ܽK�ژx1ぅ!W���4���b�!�\*n1���_�&��̘ �V- !�V<\�،ك�M�0�Le�wa�=~�!��' .���&F)f��qh+�A�!�$�?dbt�A�ε1��U;�HV�jr!�M?U�<Zs���W1(�`�V%@�!�[u�����#�-$.��4h�7d�!��^��Q9eρ�jb���K!�$�7�^p��eߣ7���hH#&!�ƫ�2��D�K��F��q��V!��ޮ7���jтS����GA�_!��%?j9�tOB��P!�F �%�!�䋜HR�ᙳ�ի��U�wMI�F�!� 1	�a���7v��)�ꑔ`!�䏁a��]��  "a�eB��)s!�d�\�x�D-NeK��9�ʈ[�'-���5/!��uт�T�'��L�
�'�<������j��Q���!?�8*
�'�L�8laD�8+X7/��
�'�b�"!mH�~�!�ӣHaډ��'�4@󀦙)^W�����A�740h�'��� �� uCt���� )'����'FB��խD���A%D�Q��a�'c�$ಪ_�?o XCO�!T�����'�������9�v8�W�P��D��'�V q7[~��uDhV��rAa	�'۔���2j0x���V�w�8*	�'{���/�}p�1j�jU8vg����'��2�e�/C��� ��=�:�'� h���Z?v-d�cI��<wc	�'s��5������IШU�2����'�툧-E�h޶�CgIR-3�`�	�'�j@҂�ǫ4֖d�֏C#2dq�'���0� �+F�B�9�"J�.�L���'A^���/��w��	�0%B<4�j]0	�'�,��r���vI�X��H�A�>�Z�'6�$pu 4c�����ʓ�2k�(��']�
��ϐ\������[^�D]H�'FV�H��-Fc�Y	s�Y�;�l���_��xBvLT�����%D�1��K-hD�B)�g̦�`qb@�:�N���#MRl�"�+@s)��qoe�ȓ�FYpe� :9
��#�ͻJ�	�ȓd{H|�$bE*��C���3ˊ8�ȓW�l=r�EMd1X1��.4�����S�? �-��7�U(�M*W�|��"O&]� h�*o%Z���W�T�&@�`"O4�����}NL�ң/ 91��	�"O��d"�$��-�O�f��S�"Oȵ��� JIy�@:{�.q��"O�Ըl��I
f���d�O�>a�@"O���f;�:Y�'�Z-� ��"O�UB�n�ހ���Ïk�4��"Ox���j�����)�8L�<��5"O��סs	�����P
Dp�"O������p����(!�He� "Ox��CR5~�r�GĲj}`�
s"O`h�Wd�Yh�BC�6MtTyc"Ob��"��)F��	A�ֳj�|�"O�	� K$���CG�
���a?D�(C�Gҗ v��h 僑t0^�ؗ�/D�,��rX�V�)%��X���.D�0p6/�>EL�5�F�Zh&pn,D�8��K�jh�T�� >!)��(D�d�C�	�!���CD�Z��|��*1D���J"���spȃA�X5{k.D���w�I�lPgMA�ErPq	�+D�@rP�4+$��СjRw�<	Y&D��C�J2� ��·^)��a$D��D�5��|[����X�=Z�h D�T��~��\�ҩ���"J D��CF� &`������ͅ+r��B�>D�DA�,��P�f��ƈU s��h�1G;D�x�Ї�eV��fǔ�{A����h6D���VeB�.d�p��oѶ6a�P��4D��3#����� �N	OВ+3D�@�aĒ/}��;��o$�Ya�k0D��w̝.@����)���YzD2D�H����
I��&��0 �pc�3D�T��*S��T�hRBQ�v�"��1D��:R�
�e��P5M#�y[��5D�4�w� �5��q!�Y�z3�ժ6�/D�xqq$��}:}���UBR��xCK)D��P4�%�x�D��T4��
(D��؁��b�y!pLўYUV���+D����IKd����1B�PX�p�)D����=v-�c�/S
l�.��C�'D�H`g�)�`�p0F ��Q���8D��Q%�S/s��X���7p~��Vf6D�Xa��	N!fD�o	1`x!�2D��T�M�:�f�F�>NI�0�>D������!��fL@R�8�R�"=D����
?H>!�t˜�;W(-�!��y�`�H�k	�V��)b��¦]�!��,Ch-b���=2���N�	Z!�$'i5���>��p ɢp=!���)e6d�5H�T %��͏p!�dGzJh)G���kըy��ٕ3t!�Ă+"���r�v�k�+��]W!�D0� 51��c�N��ūY�U�!�D��ga��pH��}�,�w�Y!J+!�����4��/;�dQ`e�KZ!!�d�C �r�����q;%�Y�:�!���?F��D��$-�,����.:�!�]�X��X�b"�u��ih���l�!򤗋E��}B�fA�6�&���͋�=g!�d�T�Jl�f��-p��AU!�9Y�l��A�-I�2�#B�[� !�DR	Y'���C���p�3�h`�!�� ���D�5=����H� [����"On�RVJɆ1U���Q�0ipV"Oީ��#�41f����G%9 H"O�=�u�WIL��
pk�:�!÷"O�(���ѭ)Nʇ�<"��e"O&��[�&�R�c`ɉ/I*��"OtM����b�R��B�\���"O�T)r�0}���R�ȽD��Y��"OP"7&�%[���\���Ze"O�+��O�G��RbD�\,B"O�,`w���Bs.�A��M�#7ji)"OI��,(W�Ζh 2� "O����h��Y�\�+��Ѹn^��r"O8l�#�J��-�$�I�;�e��"O��y�)��4�����EU��t�1V"O���P$X+|�RU�: �����"O��Y�e'6:h`�O��ih<�W"O8��	܉]�����4�qU"O�C���!��!si�s���)�"O�u����].�j�NP�l�R�+�"OTɳQ�B 2���J�� /,��� "Oz���@  ��S&�̰n��`e"Or�0VB�k8�)i[)$�$R�"O�����vՎArFm�H Pل"O�ek����SV�r��Y�A.��d"O A��o <uAV-�QC�; ^ݫu"O6AgɣS��]S�"@�st@��"O����#+���5��L��l��"O�����I�~��!ͽm���[�"OX�:�B�0���
D1K{�<I"Oz�I��)�@pؖ�Gg��×"O\m�Gɋ�d}�M@�iش_��a�"O�e
֡�D��Aݒ�i0"O*�����\DN���@���``�"O��
 *I(@UAF-Q37�٪c"O��	�Κ� ��A�K,q�c�"OZ2%�j$�8p�ҍyʀ
a"O�`�#ʛ: �k�C�"K�u:�"O:1��g�@��l���w"O&���i82����Y	r|
�k�"OR-a+Ik������P��-s�"Od�9S�����#%!M�Ф$p"O���t�W)Sgt��Ņ�VE�v"O��z�)�~�ĉP%�R�`�Q�"O�P�# �Kf6�;�K\"�����"O����,I(��Q���@t���"O����'1d}�枓3�*ͯ�yȒ;aL�Xg��"�#����y��]����4!���,��RLQ=�yB�\/>UZ�(��Z3% A�ں�y�]�Ya5n	��z\��%�y���!nx�(e��)n
z��SIʒ�y�C�T(6���ũc����B� T"�E+BFbi�&,�=5ԐB�I�_pE)���m�V����z�B�1y��Ѓ	XcV9�U@�QN�B�ɞ(r,3	H5;(�����A�#pB�y��	R'K[�Y���02#�'p`B�I~�~����Nl�p�Mڱt�C�I�D#�D�3n�35�H�;@QC��:ڌ{C����T�W,Öe�B�kZ\%3�,7LQ�x�OA=�zC�:�N샔�L(���x�D�.	C�I�پy�󩈢@�fT���
'��B�)� ���Be��t&��"�<:v���"O���`�%>���� C��0�V�$"O��R,�hab`��s�����"O�u�,7J}bB#/�PZ�"O����lC0H^�p��S��$�c"O��Z�]�v(�Tr6n	� .鉣"O:��,X�1
��ˆ�Q:q�Xa"O��g���a��mQ.���"OhA���8���A�f�<?����"O~��w#�Kĉ��Yf�H�;�"O����Ɨ�V����`U)J-q�2"O�D(�%[�1�BԪ�	Tf=Zv"OT��e�/XR��������"Oh�Baۑ ���aQS8V�P�"O4�;�Bd���1HF���:�"OB�K�G�y�ɦL1=����`"O0�V�̟Ps���3�Y�x�4�J�"O�,��@۶P)ؼc�C��x"O��9�ɒ������ƈ�W.\E��"O��%/$3�@��Z�BL���!��7c_�0��E|H�� �6;�!�Q�~������K8,��/A4�!򄄭
v���/͢h RUʴmR�&�!�䞡n��-b����4B�+ޡW�!�d�<��c*V<f�@tkcm��n�!�$P;$
r	PΔ���s4l�	s!�DӺAQ�yH!�^�l��9aR���M!�dY�C\�ƈ
&l�ڠ �-�-J!��6_�@�iC?��I$l�*O!�4��AjћI��D��	<?!�âZp���$�ë$^L�g��+d�!�DO�:3J�q��I�jX�kL!�D�X(��hb��_�(�;���'$D!�D�J�`���鈔m�PC$Lэ>!��I6h�xd!L!?�m� �!j!���l\Vg�>*)�E�B
�>!����֍�Q���J7��n�!�ĆX;(��Bq�h ("�ՙr3!�B�6ذ����Ż/��I���/!�Hm�4�#ũY�g.�e��T�vC!�$O�R|@���:�]�B��Y�!�D�>?��,[R��0J��I�%fr!򤒺2��p�V,bd�ڗIH+`9!�[(Hرs$��`��$B.�"z!��"��={��^�B���!d�I�!�ܟL���aT��"�n�) ��30o!�dǎ]0��F׬7��a�ˑ.�!�D��-�p�8)p��p��ˍy�!�D��G�����55V��r�NO�(�!��15{��*GK�%2�� �M�N�!�%z�A۱��j�j��cC�{�!��@�
��'O�CT�X7bR�{;!��W������ړl�f��/�K*!�$��tƠ]����}Ş��mI�1�!�ĆoU��;1�@�B�����8�!�=m��8�;,����e�ə�!��^��1Z�+�UQL�"�'0�!�dP:mU����,J��\x��)w>!��	�H,@b,D&"6�5�!�ŖR��e��K�Y� �w�+	�!�D�nz`�0c���fQ�t��q�!�DʱTɶh��G�I���a��>?�!�$Z�CG�HCF�F� -��!�,�!�OW94�z�%ׄ o6|�B6X�!�� Z	��[�A*�D�&�6I�G"OE �k�m�"t�&TnC���"O.5#'�^.�X���* <2F"O� Z�����:�-�ruxR"Oj�mֲt�N�!��$1_zy��"O�]�ҡR.1��K$	BLLH"O�`�U/eƐ����I�1Y&,x4"O���c͊<Vz�e�[�^p�h��"O�8ڂ@L���	�,�2F9�"OJ�r#�XY������kblC�"O���I4J�X��0��C��XR�"O���ۨ?BUK6�8j~`9t"O� `�Ό}�pȉ�dK
ov�pa"O(0PvdK[!����L&*/��A"Ov����މ35��!�a �% j��"O�ɭ�^�,;pM�e	�S$�s�<aU�T9;8��*�!� _xh��� h�<Ɇ��
B\Рdc�������d�<1S& 
g�*�)2�7v��p��/�k�<���%|�l��t��5m��6�\�<�	,H��s��ʻEF�u�__�<��n�d�2@�;_�͐B�X�<��[x�(�ԎU�I�q���H�<�g��=M�P��JP���T�D�<a�*:HÐ��j�<� 4�O�j�<A��5Z�D}�"�{����Q)Tq�<	�%B�A,���dJ֍"�#!��F�<y	J�
�^��WM2�ԙ[2@�<٦ϋ���9QYq��U"q�Ch�!��[�T�k���<h�v�pIi�'v$p%�*$����#�L�&��'��x�O	�)L6�CQBюC��Mj�'*�E9j��3q����  9=�!k	�'��8Ј�3GPn}���_:���'V
��䉜s[�m���۫&��t�
�''��ف�Ϯ:K���l�da�'���a�2;������>��q�'�
���݈	3R��7����*Y*�'M��x�j��U�)p�����4��'���r$���,�c���
j4�@��') ���L�_X�p�$gʐK#�e*�'f6 ���GI��r�Õo����'�"�:%�(x�}�B��<k�āS
�'7�<ӳ'�;GDR�����M�Zm�	�'�z����D@hXs�	M?�<�Q�'�F�ȳ�Ł^��Ȕ#�k�A��'�p̫g�AJX���S_r�QA�'�M�B�	pe,@���W��J���'�nH�/+4�@q�����)��'��K�l�Ԅ�sJv����+U����	<3�uq#�671��5��+'��C�I�C��9B���YG����a�+&�D{�����h�e"�E��q��dJ-]�N��Fe9D�H�7JfQ�X�)M�4"m�T%6D�D��S没q�N� `
1��2D�� Ӌ5����z��2�a<D�҃�#�$�Is/9oh���%D�0���T*cjh�S	��N9@wa�<��M��K�'CW��={S��)-��̇��w~��^�~)z��c��d�pZ�$��y��;T=�xA�lȌe0�A�'��')�z��F#sOn�jÑT�6l�b�P&�Pxҷi����4�S�$�RD�D�O��y��'ў�S���'�`I�
�4\��Q�I�҈�8OPHEz
� �rq��%��!��ԯyIZ,���;?	�]_Mɳ��.1V	Z7d�?V�`��Ƀ��'A@��R�
|
ջ��
�i)�'�@uy�L�E�ش0�(F2��I>�q-f���O�L��t�S�Z����¡�~��,K Ob,�@�$�̙�So;C��RT��7����#RGVR�N���h�
� C�!�ߑ*�L	C-S�(�t�@D�0�P��ȓ�T�S�	Y)���� g����'�)�� A%�Bm�2�J&E�;��}p�/D���O�5$�K�@B�!��1Ԅ�����I4B��a�O����4kE�l�B�I2NW��&�M�@�viH"(�!d�B�I73�8j�f�+P.���D9W3dC�Z�k1���,����Ɗ1R�B�	$y!\���*�1��_>5�C�ɩ}+��6B��(K��v�4C�I�r��ęeE��z)̸ۇM�2�B�	..R c�cY�S�ke�[�6'B�ɧ�"h��Fʬ$�T�Rc�D%B�I~�*���4g�� IɺV��C��1� ��oկJ���y�%L911$B䉫5FMc#w�8��6\�B��~�m�w.˽Z�t谀�݆������p<��(I3���)�FB���["
�Y���'�h�* #�<2�)p��@�'���7斌k/�"Pǚ)Wd�#�'v����N�-zM��o�#\LX�'�lXP&�Ie��aw��YO�!��''v,�v��R�q&�M &b�
�'V,�����^�B�{��.�p��	�'\B��g�W3D��I�&����'�A� �Q�(9�i�H��mA�'=T�9'	��L���C��
�p��	�'�S��*CTz�&��1����'6��Wi�4K.hH��h�8��Q��'4
�;��}UX�	&6�H����C�zPvikT�@\F9�3e%Gd�V�)���1�z�4��ڱJ���1�.�*�O0kC,�.3г�a�)3 ��(A�'8�N-$�	83J	>W�+��V� �ȓ.��%�(ڼz��Mb4���Iv�'��x���1 �XBĢ�-y״����&D�����+I���0.�t�tT2� &}��)��%Ӱ�a�[Pdb�L{�U����s�Hണפ5��l�p�D�������5D��:����6Y���A�NFn ��4D��ɇ��!��h!J��^�(��0D��9�d�U�(��E�d�͙ �-D��� �Գ\��g�,+��c3?��Q��ħk�)��LQe.����M�1�Ňȓΰ�s��6���APD��B��@�<I�
��b��SQ�R�B��ܓ��<)ܴ1��XGY�S�RQ'K^�B�.����>a���	_ކH�� �j�� ����B�#?�M<!J|R񄙞
^l�h�IMK����y����-mGX5ƦZ!L�h`�v�Tцȓ`����6���!ɉ�%�*�FzB�'p1KA��9�Pa�`JB�+�Բ�O�=E��ꄯm��;��@�%��! ����M�'i���v�Bt��h���w�@��'�(p��&W�Pk �@'�
�k� J��hO�ܨ�Zy�乹�K	T$��B"O����ܠeWH|���Vڌ:�"O� 2U+���0A��R㕰X%:%�P�D{����?�Fm8�:,;8�a��8V���)��]��#oF U&G%M..̑W@>��#��U�'7�T�D=v����S?	n�t�O���dУ#�Q!d�$��sfb�s��yB��>���P��1����q�sā	y B�	%��9����"�2�ȧH�,��C�W�^}kƬi74���ޔBYC䉛k���QC	�h��p۰B��J�C�	'	�3�,	�{��I5N�7m^�Fy��s>�k5�	�E��y�$P�~�Qo��d� C�I�Z���v+�`�����+\t�b� G{��df�.+�4sQ+ƃ�hl����=	q����I> ���z���iI�l0 �%)΄b��@�'/�d��B.W��BDL4������?qI>QgD�<,=��Z�f^�y����2��x� H�O�p�$ϾjY>m�!�����O�˓ɸO����ĭ�O�B�x�,�ŐA����x�fGqY�=����`,��T-����')�	!�$�#l����m�7
:8�B՞BN!�G �h�`�<h\lD���0�1O�l�)��?T�Xl
�N.�$2��&�C�ɱl��y*���73����G��*s�C�[�&�q��"n�(�ֆP� SxC䉣R`,UƉG�Uh%�A�{ph��6�O��Bl�M3��I%2�#�~�����>�4�j��b!�=(�F��Gx³i�a�ā��Q���36J�4	i詁fJ���yR�Ƥ#j�0��K�
BFqi�M0�y*��	�\Ŕ'n�UYQa8�y�V#��A;�e�>T�`�[Q�.��UX�� ꌵ$+�u����$D �f>D��q��ΞE{�X�g�6=��� �+0?1C�	H�'�X1#B!ؒX���ydB��TG���}��|�~�0U�`y�a
�xFM�$��y��h#��t���O������E�̍��$�7{��ˈR�xR�UR�,��B��o�̸�VBђp�H�$�鉇{HF ��Z�?��T*"hXDc�x�'��>�ɴQ�N�&'������+�xC��,U�dN98��w��2ml#<�ϓ)[����@�� roW��(��%�����#ϳ`9�!P��pc��'��}"dI3F�`�v��P(�@�7o8�yBĊ:4j� ��HQ B.��)�̌$��'�a{��#U����Fg߮8��ʕ∪�y���#`PS �5��\YI���y��	gE|�ŉ�	1-�DyG����y���6=����3#,!�Ԕ�V�٣�y2�JI�D:�"P!J�r�6�yBN�p�4jG���q�ï�y�E�YZ=+���%_wP�#��\��yrCƠ�r��ʔ<z~h*�5�y�X7)�蠺���x��8�
&�y��߄N؉�T+����l�d,1�y��ޔ�����ʏ�	��$`�����y2��5�4���1��mÈ��yr];R���J'�!?��8bI��y2�R�[��`���d��@Q���yR�ؘ^Fj`/�
^"6P�0`ʭ�y�&�P�s� H1g�F���n���y��	6t��b� g�� G(K!�y���"��Y���`�iٖ!�y���!^ÀM `�4ҩ���T�y�B��H�����	53+���a$�y
� V�"�kI�h�P  ��1��h�"O��
s��f("����Z:���Q"O����j�~i	���<zs1"O�D1t��-j}�%��BV�V>���"Od	�aE�4��p��a�*F�Z"O��`��N'��T����R��"O�\���ܗ��'�6:�m��Qp�<�t*ѯB�!1�/�Iy@@l�<i��A4ቒ
�S���Pt�]B�<�Q/��l�Jݡ`-oDVD(��Pt�<�e�Z-f6H
Ň�L.aۣ
�l�<�!��'��`��M�H���{�l	e�<�2@I�S�H�{'��bDxxKc+�c�<�c� ��ܹtj�5Y����I�b�<٥���w�r!('"��6��xIbL�^�<�P�T�_�B;�D�+��i�I]�<�6�A��	"�
�PYlh�th�t�<)vKZ�l�59S��r�x�[ %�x�<��e])o��HV�_
�vG
t�<A�
��S�X�3���CF�<)7�;Y�Ee�K2BJ$d���_m�<��J=I�vm��$4 ` 
g�<�!��u�(t	��5c8��Ki�<��6P���!Ʀ1Z@�	��n�6U^�q�C-��]{5�#|P�<ђG��Zh�� �[�pH�ˊp�<����/n4l��,O$h"�#ŀo�<YG���|	��<�\Y�#�j�<󊉑��(w�R��P`���j�<���O"\��J�~� ��`�<y� M[�x�9G�m^.�PS[�<)�a�<RdWR�m�h%A�b](x!���w��\k�CE<%���`���9!�Dz���#pk�7�F�!F���<9!�DT�T�Y�F��v�F�í^!�B�PD��/Y�o4x�uJ�`�!���+L	҃��P���	AD�!�D(��l(rO��v�Hr��Ƀ�!�d ι��l�(�I�Q�t�!�d�I/`\Cٌ�� �"�!��3$���eF���%�"6Q�!��Y�=N���NG�*�֘�Z+O!�du^���F��7v�)���B>!���#1�DX��R�p\���c̘x�!��%3,p�V��a.���!W$-�!�ŮZR6�8�Bɧ:*:�;���h�!�D��+rب,4� ��a�|B��u"Oj8�W� >�TѲ�!Ctu�7"O�)��A̩XN����G�'G(|�I�"OҼ���3Z&��gU���:�"Oz���R�� �Ӽ���"O��0G��$L������s�z�
�"O��)�b�3S.�#��F7��`�"O\y5�D�2Et� �z�D@�7"O�92ah�/s� ���Q���q��"Or\a*[	��U`����:TQ�"O�IА��xI[�Բ{�0:&"O�چ��LLڀ���"@�:��"O	x�C��H�8�J�U�ıb�"Of]�TD�0�������xxLDj#"O�(0���b�b��!hR��"O�8��D1��тe�/0���6"O�5#�E�5�Ƒ�e���*r�"O�"��B~0*�3hC����'�NX�c��cUX�� b�"��	��� @@Y��Ҩ���{v��_�H�x�"O�<0�I�I�2��Ц�}� �8�"O�1z!�ý0�=���8}�ZT��"O�u��G�	(y�'���B�"O���EY�$[:i3fD�!���"O��E�,c����Ԙ2섙r�"O���8�4�B"�|�*!:e"Op1R�C�h��"& X�I��(;�"O"���Mڕ4��IX���p��"�"O� ��G� 6�N�zFnu�Jd��"O���#��)A�	ꕊw��zU"Oxk`͊0%7V�8�I�wi��s"O�A����2	ʤ�`H
tl�8��"O��J�B�y�`�(fE��J�QZ�"O�,pƏ�?T�a�@��*v�>Q{�"O̴��㒴v<T�"W.�A���"O!��@�`��պpdY�:���"O\t�v.�C�h8����#;N�c�"On��ը��P���mٲ)�[�"O*��iR�lr؝��,X�b�i�@"O��iƄ�8L�FU����?l�1�"O2��4ɒ�`�hq�Ձ� ű3"On�3��T�5;< �F��$�n�6"OpAZc�X�h� �v��$��g"O�=�#��,t*J��VL46�N��0"O6��C�7y6E���B99y���"Ot� I,�D�$�Մ�Z��@"O��"�AJ�"��Yn��)J�S"O=��aЉ5�`)�-FPݺ�"O*�V��o�ѓ�)7��a�"O�XR�C(W�V�B�h��8L%I"O0��f�:i�g�;M����"O~�0��cX*0I�:¢��Q�O,�r��2�?6�N�s=���O X�� ݘ� �H�^���i�Dp ຕOͻ�?��� Z��`�Gl�;(��Ղ�$f�e�/���Y���d]�U�u Nض0ƈ^�&X����P�I�����J�5�H�:�KGV�2��h ��jb��֥��%uh)sH΋�a|�,4f�:Щ�2HZ��C<�����#� ���'>�{�hLp�(L��x�I�5��d���X_��q����W�VB�,���YĩQ�+�m �o� p���ĝF�%ڒΛ ��!b'�����'�O���0Ro�<<��HJu嚺|,kߓUR����aA0u��6R�~�yON=N:��#l��O�4%�7�Z���N�ܣ|�'h���SA!4�6��n��v�<�a���Z&9��p�QH�O���Ruc�3U�CV "y�����IH�V=�3���1�0>YVԔ6p�9Q
�=9���ˍ�g�Pe9�M�����*����N/5�� 5��n�	/�4��1&N!�$J�9����	
S4tI4�ֱz��g@�"o䀐`C�E�b���
�8��ħt���[�!��W�b蠄"uBԅ�I%�;���0�5�PK�:TYE�4�D �k�X�U���|�+/�g}��J��=Qm׳Ϫآ�$V�(O`=������*Kf��jݵx���'1L�k技����qa�O�Ik2��=�>I!ٝ�^Ir�&U����e�B�'��8�LNE��>�@�*��{`�Ҽ1�h�	�"O8d�p)ӡp�nzT/N1^��xH&���>2G-��F���8�>T�d��w�X�mסH�HA(YW��X��'���yA�[�
}C�ʎ.@���޴<m(tR�[#j�L��%X��	�X�U�=��ȅ8>a2 ҕ��,mۮ]��V8�d�)��T08ZA�;��M�⣕�1�$��a��t��D�qEA�6�0=A�CFt! !L�w�� ���R�'ZT<�nBA~)�'��8�%��@�0�Y �ŵq$pe�e&���J���A�<A���5Av��2�2#��$����*$�"AC��(vV5#��'/F�R�6Dq���}��1a|5�o�>�F�C!�);\C�ɘ!1h}�&�A���c�i�v���	BcV�Fff�y��:s�
�q��|
��D��c�P�nAd�����F�ּ�qM:�O�s�nG7o�c� �'�
+�P���
ßRk�tIG.Ο��IԌ~�$���'�L�f�Ԝ=u©���"�D���D�U��<K�*8�҃��}�B�0JL0F�V�B<)(���A� �E��M�ȓly��Cg��Y��0�"��4���!>sRy��a��q)Rj�o~��'�t�'B�l�����/e<E�O���/g8M�@��(�T �A6<�`xC!�ZX��%�R�K�c�r��W,�7F�1��� (Ϭ�Vmg���,|��<H�CC�)#�M�!�>���k�ȝf80��OH���:�p|`cń�+� �I�M�C�L�bv��BlU���P�Ж'[h�0��O�L��<Y��;UQ�TZ"��?0ՀL��C!eD�cee�$2.�3#�H�I:��	?WR�\JCR���OBL�"ėIo�۴�E��}�4�'].��.R81e���'@l�@1g@,~	��&��2N ��sOJq��i�,=	f���Y��'��F�	p̓?92��tF�'F�l��4#�dҴȦO��B��G	%ļA��gg�4�1�)�<Y�$�hA�Y5(��Ԩ�璲��-I��:����'���TX:5��O�Y��m��C���g��&����6~ٌ�8���Jw��Ǔ^�E�'��D���$g0x2%�e!5z���ZwH�:��c�`B9+�<��"n���rH.l��D�BϦ� 	rF���ht��K�@&�TZA�Ѡa�|�&�j��`y�bϦ�:�[�P�EBJ�]���GCWB%Qu)^�p<c�<tY�դyG܄�2��
���j�:;25����Y�����a��(����C�R I"��u��@)Ŭ̜�\:�W�BA��\�f�zDӢA܎_��R�A�"J��*�ԌC�7C����lkP,��Q�S�D�8\j3�I8]�N�5d\�v���f��'n�	a`D�XD�q�lb�*B&@�H�D\G�'Ɛ�Mި1��M�SC� ��m�3���P��2j]�89L{��59Ô�3E�)3��I�S���m�Ì��Wo�Y��O+A?�U��$߾{i��HS&<��2��'y�Ճ���W���x���A�8A�UkX?=(�7��ʡ���%M�~%�w'�7m�Ɓ�ah��O��QΓ{r\����;�>IBꁤe��0�C2�O�5pb��J	�Q�SD��`1��3�gI�m�d 	�/�,}M:!2fC]>2v�$�&
�v���4O���G)�S8@BX$�p@�]�]�G+ޢn�ޣ<�j9CEH �� �Z�I�k�b���՜\�h���C�dV�`�D�pDH���5O<�x��$APaO?���5/T��L��
a��Ô�R�yisb��;�RQ��O�'X?H�F�D�Ǩ^:����fV�se�H��IB:�0:Ef��H`rk�����>��!�v�py�嘘P�6����9�`aW�ǑdQ��Q�钫/�Q�;<Y�A�!�ٕdoZm��ʫ���"���Ra^�$����K�u�j���T�Z�0���
�SN�u���9V$���mA�*��Qu(�5Tp^��C%¯]�t���AT��I���O�n���A��R�ƨG<m�d�r��RWkH�0E!�e'��"�l�z�*˧(X$m��F���z4��!���͚�e2�G�b#|�'�L�h�%�5P{R�+"�G�À0��
Z�Ī;$�!�cc�bE���9��h�>|�*@
`�*���"O,]��G?^G~�M�J�L����
^p��%$�%
�$ʴ�O��)'�b� ;B�F���uz�j�9Y"Q��#Uh��
����K���.ؠ)kT����V�����& Ux��(�
ԷN�qx�4�Pv�7�d�r��
U�H�Y8uN5�P(�E�FA0G���v@ĥQkTŇȓNmDU"2�ڜN��d���;{4T����% ��ѹT�L�2��wEl��?�$W�E�� ْHv�1�R�k�<�@�S��-����B��t�F"L%'>�D�}���h���l"�D��HO 5X�+ֿw���r#L'��ap&�')H�۠�!�p%a'%���-�aǒX"%���ғtV�ԛ��'o����W��U��3ي((�����.9bԑV@�8xnQ!I|2eE��[����A.Z��8�6D[G�<	�T�jT5�c@7������B}?)����iU�'}����!~�8�
ï�6P�R�p7@ԩu�!��'N�Au�ŋH���0�M'��'�ċ �YX���#L4�P�C�8Y8���I7D�,���Л��X(�C�T8ā5a(D��p�ˊ��݀��B�QUHI��(D� !4�_�,��@3�;>y�1+4�+D���H7�1��o��S ��(p�(D�(r��� �0�2��>.�24�v
$D�p� k����|�B�0!c2�Qq�7D�\� ˛!T>�#�N�H#PAX�?D�\BV�ZQ@�
p�C�A\��� h;D�t�0�ٿDQ�ֆ%0�zt
��-D�<���\;A�j���<	����k*D�p��W75bܢ6�`��G)D�b7EY���O��|�:6�O�<� 2���f�O'� "�ӆ8$ �"OzH2����D���OU�] 1b"O�T��e��>�t���Hا�,��"O����+p�x��2���p)"O<q��E?�j5�Ek�k�޵S�"OŻň��ىF
ōz��Aː"O(=X%拦0|�k�%2�(�8�"O$���N�d����Aj���ҹ:""O���'�%.����`D�vl�<�F"OR�c!Ö��hWj�,lC�h�"O����lA�������\�8p2"O�- ���<D
[QҁR�n�q"Oj<�Kӓ=���ag	��(<H1"O&+Yv�)E7�pQ�"O�QT�Z� �68R�J�Gr4Ћ�"Oа*�� �ePl�d�)2f\�3"O�,ZS�����+�'52��Kv"O:\+'nǰq�ٛ��ՐM;���P"O�i Vg�p7�)�c�)K�	�"O�1��*N%U/���ɷH��e;�"O�dc�(B�%�*����Etوy��"OMr�/��h��	G�2��+"O"��Ӄ�"��`�'6�Ч"O�b����$d;u��5/����"O�� �DU�i�~�W׫J𱹧"O�y�n�L.,�"�AƨK��$�p"O�q���C<6���%��?v�s@"OR$����bhp���Pd�j0"O UKQ�%�VIQ�kO���2"O��JQ�U�
n� 22�������"O*��4��,x@�)�-�b�J�5"O�5P�
�-��8a������2�"Oz���+K�0��B�z�yG"OJ��1kٿ/�XL�Qj� A�ɘV"O@�y��׷|k��qWB��u`�"OB�z���}d����*��T٦$��"OrЖʚ�c�*IB���D�"��c"O@$�䍺-3V�ʱ(E,'֔!�"O�52G�1(˔阠h�<?+����"O���d�L�_m�)!P@� 9��	v"O(i�*R*'4h��f�,!�xZ "O�X!�U�i�ءpV$ݫ~a4j�"OLu� �F�A" ���T�0PJ���"O� @�͘���8�@�"�4a!"O������z=d��dR-9��Ȑ�"O��ʴCҧFΆ�EW-@ �"O�Đ�N>J��S�e\�^�$	�"O����8!%J��iP)>޹�d"O�u�Q�q:�-�H��*r�'"Op�Re@��|�����t��T��"O��˔�2:����4[�� ��"O�l5�]�q�z� 1��2���S"O.�����	HD�!0R`�3s+�p��"O�$⑈>�Z�P� �#)�ɠS"O�� �Ɔ&������<o�R"O�DJ�ٱ?#@�R�G����"OB�[�X92 t(UV:M�����"O��(T%2��d�3Bɔ|A$"O��"F��B�ֹ�qH@9).:!�"O�<Сk��p]<�3�
�
���"Op`v�@��p,k���*;�D��"O ��ԍ>(��)h�(�"B0D�"O,���j0M���Ш�%D�ʰ"O��σ2 uID��E/~ŀ�"O� p-�a�5F8:p&@�`��6"O@�؄CV]�� "��&eX��R"OJ�5�O%]̚L2�U-_n���"O��A3C�ti��]%L��"O�\���D�
���GG%���P�"O���F+ξ~�����x�  r"Oح�`�+��BUR�����"O8�)+���aK��Pk�"O�`6�^%��T�0�^084"O�5{ԡK�Xw�%�ꒋY!D���"O��׎Lh�����[�,)�蛡"O���f�J M�>Yҷ��v88k�"OЄ�AA�پu�O�h�vի�"O�]!�OM�.���3�NX�0�T�"O^����L7�l��&�H=�>�[%"O�a�<)���Ж�!{�(h�"O�)H���3�fY �0]�Z�� "OޡJ�mR�E�bE��gQ]����"O���F���F��(����D4
�"O��I1IN�UT�H+􋍧%��q�C"O�m��jXp��S�*�)��H�"O.,�� �.M��ka)]�zs	��"O�D$g�/WZ�'�&\b�t8f"O�^'w���+�FT��	w"Or����[�V����bQ?'�jx�u"O4��'��!'nD�yRf�<�Z�c!"O��ad�ыd�,\��%G
��u��"Ovi��H��J	��W%9��H��"O��r�ӌu��)�A̤FdxK6"O$�{����}���%oƻ-X ��'"O��ڥ�

f�n�㕮�&8��#�"O�e�r��ؔY*'�]�r%z�$"O� ;�"	7�P���Y��Pf"O��b�.��d��bK&j����"O�X#��Q����u�Ȃ�~�Q"O�p���S >!B䀕:p���"O��v�� ���D�D�7~�D�O�Q�g��?�H� +�|��O�����].���$��1>� 
�$t�A���?F-X:�py�� ۖK. ��'�cшa�C(7���X�����p����[N�u����O�蔠�>&�ҍ��P��l�H��V&Z$�<� �>Q���'`q�U�'Ox� �� s����#�(dl�L �DE��) gh>}"�~����:����rt�(x0Q�Jx:�%��_7,��	3D���
:Ƹ�Q��ɹN�N�!��O�t��s������V4�S�*}�����#P=�5bɢ-��Tx��Y���=���ˇU����g��	���*j#�2��$k��x �j�#H�ʽ��>��5�gy2'ҟ����K!u���1��U���'���.:�a	8ҧ�%:� W��`��F��'WPF�)Ѯ��vh�)��VL� �@�[Z���&D
MƢ3*i�0e����[�	��x8y����y�Z20R\|+�{Y~��	��y�"�#�I���٦he@�b�ݼ�?12�%k�u�vԭ#���㐂����Ih��1���	�"�.˞��w��f�������9A4$�wM�O�aa���a(��&jFq(�s��[�D���N>y��>�D/\�2�T �Iѐ9��!ƖZ�'`h��dou�cR��Z�)�!P�H�X��@�Y�v���p�'��t�_X����)ҕ�v��Rdۈ_�T��$�0'�P�Diʍ�(���hb���:%���Q�I��$Q�"O�X��I_�Phղ�B��>����5_��!pE,*+�I;9�|u���w}q���ΧnK�U�ck)N�l�	���ͻ\�b����Z�)t�`!T��>�Ms����~D|����.���f��c��}�w��)B��_r~� ��n�'P[���	:S�T]���\�q�l}X�B�Y#L%1�A;�|Ъ�O��2�	"�I�o �(�ĦO9�$e��I9 �T,FyB�#j���Ϲ�y"f�8�@�f���8C���0w�tP����-!G0ԅ�S�? Buа��"$C�*��]C:\*�'ԇLn"�dP�=�Q�I%pVE�p�V�&Aq�]�c�Xab�Q�O��yҥ�K�
����ٕ	�+)P�v�tyWҠgn��e�wp5
��|:�f׹b]2b�����	��9J�ϗ�_yy7,�O|�i��\
69���ʹ?B�д��=J7�!Y�	��$��NѲ���CY��0=�2LKiԡ����c��<�T��K�'�ZD!�	D�2��Y���FYE�f��b�\l����J�$L�`�L%7w.�z1m"D���e�Ǌ%����AhK�_'�A*���O|�`��	�����RhF��fG'���?�b�� ��9p7DJ�P�|`K�f�	�R�t@�f�O�pd��"�:xY�ue��7�`X"p̙�p��ɰ��YR,�y�/'͌a+�>O��̚}8qO��r��>	��#ɏ\, �34��/e�|�'�\P�7�\ʞ�X��A� |��~�b���-�������G��E���7��*�'5�l(B�lx��0��3��H���i���ڥ�Z���US���驖(߮\����2��@鰡\_�'Ra0`봢׀s
b-���T$Iv@8�Ǔ_�	�lεV�(����>e�B�4������.bu�mAu�*�:`X�4^�B����Ϻ)�F��5����7�-�I_F���ᇃX|y��_=k�:�'5���G�|�@i���i�&hб@�]���/�Hd	x���ng�(���/ݸ��6�X�E�&���'�2�K���)�I�哬d��s�R:G�X,9��_7X4�J��X<>�<�+$K#��Y��-g��ãoS�E��l����L��(�8Wa�<K 	)�O�x�6/Z�t�h�挶�J�`�FM��@��.V`�X+��
Ra�ty��@]�f�x����B�0�O��Z'1W�l�QvɌ�z�6x��Ju8�Г5FX'6 �����*E֜�Y�L�.'W"!�!٬A"1�CiA�L���"��S�@��b$��=�����O��(Ҭ֢
����4�N'�y�#*���
�Q�@k��Y)��I
�h����Q���bd��9F7^� ��g*�)��خESv��!�ֆH�,-��)V�	TQ�`G���h�I�H�r��A��	qz��1�6�L$=�Z2x�̴*C)o�B�	��R��M[V��Pi0IqaM�+7!�XRr&_5f�ĝ��8�r���!���@��b�$�7�8�B���>Ip!�'
�|�v,\Z����ӈ��u5
��C�%m��7�ܿwv)K4�ǣ6�t �tMX�7���;�g1A�t4ΓNҊJ2*�/)!�Iá1g�t����"�O.bR��*��}�Ј��vAly1$@{U���j&�<��DFj��'%@�<�(.��O�e(��:sv�����>�z�
Ód؍�CD��v��8,O��QR�@�)� �Y�`������cH�&`�I�	�h)�Ώ+3�g�(H~���΍�-	�\���o^
	�Op��M9ݸ���ˡ#V��He�նN�&����$B6,�C"�$�HE�mS�h��}LIc�����K��&X�lT���O��t�\�\���UaZ0��铄~���
��9/QԪ ���:� �K�+��R��<"�cB�����2���I��l@� �g����(�B,��S������86������	���T�Fܧ# R|9vE�}�p�P��4�]*" %��*#|�'9���hG'��X1���d�4`{�'��,
���J� �O�>m2�n�Y:Ɖ'/B$z
u�&9D�d��ѹoF�#��
�a�3)2}2�$  �����d��*EȵQ��}5��*x$�	�r$3�O���+I'X�@��E��$QV���l�@�ʍ$�J%�x�+�+Z�r��l�	2q� �`�/��O���%��#K�x�0��$.�13��[�eV8(�y�C��y�b\w�X$!G18�|��Ï�~R #5����Ep�퓡0}��Y�CU�Wj� c��+g8*C�	8o��ĩ��S�}��B�A�01��'�,8y%�ed�5�ቔ3�]�A#t�D�b�3����ÁnT<�X6�J�N]���`B�0��eN]�5����'���*�>
:yyt�	�B:�	����'V�.�q��+�S�����t1��!�*����B�I7"�*`w��U��ۣ?�ʓ|N��v�&�)ʧLAї��	z��.�1>�H�ȓRq2��ʐ�@�$(�&�ܤ_��}��\�N�B��K>%-��
�ǆ����ȓ7�l�E�N���r��'@/]�ȓ \��@7�8�X���,S d�ȓ,���"��P����w�	�H1������W/^�<�h�p'�#�̔��z����G��W���p�X�Z)����-�vx��'U) ��kܱT�!�ȓGd@�;���c�ʈ�dAǱCϐ��ȓ�6����ɨ|̔�[ר^�&8���S�? ����_�_ި����Lp0})�"O�[W�גP��s,�}}�8Xg*O%��*7<]vl 
 .���{�'���3��6�r�����%B��`�'��x⣮(d "��f�ġӲ|��'Kz�Xw��<Gւ|�щ �:]�	�'�@XЁ��M��I�h�Z��
�'h��:�UsVܹ�c̅~b��
�'���;sCȧR�=:�a��k��=�	�'��3��Z�0�戢���l�L���'�
�)� g�f]H�Bɖ)�p�')t`k�h4L>���`�''�tx��'�l}�	<I��;���"���#�'4"m��,w~RpȢ����:���'�TJ��ʎ@.`-2QW/s��X��'����!�J<~� qA,�wk�yA�'�a@�:c�ݑcG 6���;
�'W��j3 ��)���;49�	�'�t��������)�0U����'���h��-��-P1��0��=;�'N<U�b ��t��4��-|�@��&.D��!���$_m��%f*HȨ�
.D��s G�gc���$C�8wN�ar�3D��Y�E �TtHl�šRqH`r%!/D���GB��ҩ*q������(D���ai��3�lN�� n$D��S�B�<"v�xU �Z4�ӫ7D�XsY�1*B�
��ˤK���'>D���r���"��`�S��54�0��?D�d�ԬJ�w椡��T�G���B/6D���&N,����4�FВ��5D�|`�ߣw�蕙$�m�:��d�2�ɞj�$���B$��gh�N�c�Pd��BN�A�%��3tv�Ek)>D�`҂���Q��
�$)�m9�#!D��si�;D�������
}{R%�v�?D��Q,�V�̩�J�a�i2�	<D�t"��B ^�^�&N�KD��=D���N�l �M�U�D�N�,�{�:D��A�J�B^��TG�iˢ%5D�4�����v`T%R(T�PHg�>D�*"��%	�R�4KS%	��|:2*;D�Dstf�kX�u䅴,f�}�֥�<�V��(HE3��"�	B??S�)�ȓ<O8��/��^I��z�>t�E��o�`��m�F���Ⱞ�2���K<贌�"9�\�JD͗L{�-�ȓi[�,1v(�{ m;�aYvrza�ȓ��e��B�/j���LA�q��Ex�N�?:�� ��O�@] �[m4�)�G�q�0C�;O���V��z5�-���0|:taQ�u�f1�'�ʠT9�M�VIa~ro\A�p��6�:�T?7��2�p^P��I�[��婁$EXϖ��=I�#�S�01�f�^�5���3O̺&��˓{�г����E9&֤�Y��D Ǯ���dO?=rm
i�OQ?�q�FΰH�@�Ph��Or� �`�Gh��h��ӥZͪ�0	E?S��}�oD:w��\�Ō*}��t�2����� ��w
�;����X�!M�>Oȝ{�F�F�rh͓ӆ���X���B�<ER��� ʓ}���ȓa��p��I�<�~P��/#<�x��zc@�k�@6v6�$�f��Q��4�ȓ��@�$5ָI)3�ԏP�^��ȓ4@���RM��,�ڌ���@�V$舅���qF�
0-*\#��A�>���ȓI�q�$�$P���w�}�:؆ȓ?آ�r�.O�Y׼��L�C���S�? Tq"Cnذ0���Ɔ{�aXQ"OhЛ!��$4��֥�@�̛7"O.E��jȿlͶ�r"e�	<�~�""O
ŢT�^�j��`w�&r(�0��"O���וf�8z��>�du�d"O��s�S�d�Дh����w�v$P"O$��!��	���F��"�"O��iW6\ѐ�R�)fi("O2�+��W)V���*!mɠ[�x�Jt"Ol�	7 �anU�d򤸹"O2���!���(tA�*́_�T��q"O��˔L�7[�P�6�[�d�J@C"Or�	�Aq��2i�3�Z B6"OL{q'�B1�I�m{F��w"O
P�6��5g���PD��oJLѧ"OU+���;��i�g���zA|�"Oj�{��^������̬S^��"O���W�� ;���5�	<ZN� �"O��Э1jKD}B�)�$ao���2"O(���
<;����h�QO����"O>��/��(����ҋjX���"O���oH=h�±��H^l��ԩF"O*�K��.�z��1��"O0i�EMƈjcHi�SE	�6��ܩ�"O0��#NE�@����z�%�g"O��1G��L�t ڱC�#r�y��"Oٛ�@չ&�FMiQ Z�X�a"O:�Ѫ�!:D�����M��ڇ"OA�A�2b,�\�GM�5$�
�"O�J�g��`�,���5�"��&"Op�Y �߂"��h(��
�V� �g"O2�����i�2�f���@�#�yo�;�-cO��.4��UI]�y��T:%����Ƚ.��P�����y�e(6b^�s�[U�Hd��,�y�MC�r�ah&LP$}�(u��H�ym�1:���ic��D���@$N-�y���4Ĩp� J��@�50���	�y��k�ڼ곤՞mZ��$���y�M䂖4���*PO';����ȓ4v�T(F畴 �J����+�p���M��ŢDF��- �]Ҳ/�#>�h<�ȓ=:�m���V4��H�j
�'��ȓq>!i%�@�<8u҉r�̆ȓ)����3*������z�ĸ���� ���(��б4W=�d��V`(�-������� p<��ȓEwNA��a�Z��i�&#��:؄ȓvM ��A�B�A�(�%����@��ȓ%�-y��B�|�%c�����0K����N8%�,;5B1tt���wʠc�@�+�0�j ��8�0��ȓ\e6��&lߧ|ΰ���L8X���
"�Q�Sm��f`LU�$�@7."����S��(� � b�WYװ(ab"O�5�tNF�_l��Qw,�P�l��2"O���4&(NFp��K�+�8���"O��	�[�r�J͏�n��"O�9;0FLJ��-k�̍&:��AS"O�@�C)4h�qr�f�X��!��"O ��`W �々�;g�b��"O
%�0�Э}������N.|A*�!W"O�T��.\	؞P�BD�	a��z�"Oh�"#b4>�:���"Y�B�,��F"O� Z��f� �Hs���5�LX��"O�t Ӆ�eh�U�g��-�lH��"OpJ7�_�WR1�´qNT���&'D�x��O�^M����5Z�r��b)D����SY-֐�t4%��x�@*T�8yٱAE��"@D��P>b�:�"O��!*1OP��d
�\% �"O�"`EE���5#�4��"O]@���!���N�8�0��E"ORͳc'^M+R���O��i�"O&��ӂ/�h-+t/A��X��"O���Bi�%:GE��dI�c"O�v.�0�T:��W���9"OP�R�f���i�d	|�m��L�t�<�,O�'�l�p+�@��1�F�p�<	�d�@=ڌI4N� F�tq�k�<�)�{�e�Eȇ"�Va��g�<I���L&P���/���Q�C�g�<	�Ø@�p� �G�WY<� $�}�<)�<P��;#�<p����w�<�Ad�$�V�*�
�. �,
�mw�<I5dA$f�|4���|���� �Lj�<���Y��(G�V���Y�4b^g�<��7T���9�f�� �0p/c�<1�h�Xy����:e�PDg�<�v��t�D`�d� �D��$ƪ�w�<�HI�1�	s�aIMhڔ���r�<�i@�T��.�=�bAK�I�c�<Y�`S�R�F,��kGv�ɂ��J�<9 A�7M^8�to�v�����DZE�<Y� ��i��r�M��A2��B�<C�x H:��%Q]�JY�<Qs`�!R�:��86�@1�W"�z�<Y`�[-r�������?�*��N]x�<A���%���eH�-cTZ)Sр�q�<)шV'&
9�a`�g�Lzf�n�<�
��~��� o:H
����h�<aU�մL���+�f��)�fdCULd�<�1E�"�S�"��P��KX�<���U�P�ij0��_c��9��~�<I.� � ��*9���Nz�<94Ô7U���r#@ǜ"B �g�Fy�<�� =a=D��pD�{f���r�<#�W5U:��T�ҖZ���c�<q�U�>�8�A
��G~�lB��{�<��M	T0�+#����D,*���y�<a���U�Uã��6f����I�<���*�aahS "P�Al�B�<� �1EV����ào�rQCs�X@�<qf�sz�CGX�ZF��A�X�<)�� �����Y� %�5�S�<���'�tTG�{0�(�h�I�<9�-*Yy\@9`�M�T)x���yrO�nY���F�a0�9 �G���yb'�g؈tI�ǘ�`��������y�fT�z��9RPՍK{�q���y�'��wgP!Ã���Kg�$iG��/�y"D�+;�,����@FL�2�5�y2!�<�@i�fR�=h���ъڽ�y��P�%̄M�c֎.L�8�料�yr��<Q�H��@�C~��i�a���y�ᚐ}�L���cZ�y�N!��y��H���!��@�H���h���y���*�0%صL�?��� P�N�y
� R9
so�*�괺b�V�VZ�Y�`"O$�#�*��	�$�x�JX7A>ꩳE"O�I�@�B [)��׆�;�9�"OƤ(fOH�+��4��2+̱��"O��!v�«ZI��DdD�3@zq"O������z����� 2��9�"O��sdеHZ��C��[�?�����"O̍�2镰9�Hۿ$,�#R"O`- �>H�rI�dL�>L1�5"O��HP���`4����ݘwni:T"O�(�R�]
5�\rWɎ~c�ث�"O��Ѓ�: d6����l^ ��P"O�kq��
>�R@��lΘ7��ܺ0"O�����?'L�c�D \��� �"O�|���9;���c3jC�)s.��"O�	b�� �< ���Uu���W"O��êӠH��TOԮgi\��"OR|����,��+� ƣP���2�"O0T��O"{XlPd�Y<R� �ѳ"O$�d��&���s�(��K�����"On�Ht�3W� U1�(�	^}�d�7"O��U��'���:3H�m�ؙU"OL�!rX�S�A"p!(H�t+!"O.�C���*0;��M�-3 "O^-Y�C@� U"�n�82x�K�"O���Q!�dM��P�=s�"O �:��ܻ=�T���لj�41�e"OR�K���q���@$U2l���"O�	� R���	B��m�!��d�*��5͎�)��Bg��<]z!�䙯z�n���`|x�(��''q!�d�'������ҕBb�a���&3!�ڇ8�$����RL���pƓ�L!򤓶G�Jd�%c]:��ht��%}�!�W8{��E��Ŕo���Y�É�a�!��!Mq����EX/}��IqR$_�l�!��%\�XLWˈ/	��-�G��
v!�D�	��4PB�ȝ �t��(�	2}!�$��YoB=�reB;����'AI
!�	�g�v�ۄ�H5�Ly�g�T�!��:(��k�L��k�6���kG!~�!�DEZ6\ܸ� �: �P�6ˋ�A!�/b� u���56�\�HD����!��Z2xb� =0\�pKT��!��4l�,J�m��f9��wo� L'!��ʕMh Yւ�P�ȑ�m%!�2+���EB^q�3��/f!��\ӍȐ�ܡIQ j�!��U-_�L؁��!����z�!�d��Ld�j�OM����Qf���':�	ph��A��-�Q˞�W�PIQ�'�,�؁�${!r�Q!#?a�j����<�@w�[�(AYH���$Rvi��&��(s�T)�xP褉�*e�Q��i���*��?,�x0觢�g����,�&�>��~$mXCeC�y2�ɐL��K�	�a'ܩd,\.�y�垫3"�q	�h׳U�b����-�yNJ-�0xc���% �JQ�U��y�&:Heh��י��-�GZ��y��z�������� ��S��yR�P;3 @  ��   �  T  �  �  J*  �5  +A  �L  X  +c  �n  �y  u�  �  /�  �  &�  ��  ѯ  �  Y�  ��  I�  �  ��  ��  *�  y�  ��  ��  @�  � ]	 � < � ( �. ~6 T> F gL �R �X �Y  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A��bf�I�ð<�䄝+���Ņ��.'P:t��m�<駅N�C��{d!]O�4(�cS�<9Ҥ��Q&��pɒpP f�R�<�'�
30̖�b�LdZ��M�3�DC�	$a���ށx��`i N�{�+�3D�4�GŢ@�f<IN�e$���J'D��W��!��K�l�)}F4�w.$D�k�O#V:�b+7[�0T���?D��I'I� -�]aD,T
Z���+�*>D�$S��H��azVE�%E��)5�8D��/�= :����>�h���C,D���'܂HW�H�R���Nd|���)D��P��Q�)lj��3&ʾp�zt	�j'D���A��p��R5���C�\��q	'�"�S��P�0��JY� ��T|]D���z��|i�.S6N�ha�I?����?ɀ�'�"9C���e�� `�懐^�H�'��↫�o����f�Ev��b�&D� ��� �z��gE6i�*0���8<Ov"<1�J�2 #�3�Mс!���c7Ln�<IJٗ����`�:Иx���m��hO�OY�d%�]��h�P�ڭ/��X
�'L>��KY;��d�j�>^\Q
��� xёק�:}	��ҧ��m�ĥ3�"Ot��I��8����嗟X�L�g"O�k!E+j����7��8	9<p��"O>d�4�M���˕A&����"ONe���R�K������`&V�G"O���h�7O,��qU�ڛOi �E"O�xr�3� y1a�U�p�x�"Onf��(�d�a0�O����"O��XP�̷>�|5cԉ�z�I�"OB���M�j� ����'x�H$J�"O�b�)V��1�eN	6m�:V"O�����x̔5ˏ5j c"O2!�q�ǂq�,�C�ȾU��Y�"OZ�PƤʐ9Az�qDו"5ra�&"O�=�ŉr�X��9y(ʘa��O��=E��n+;���V�-�ڠ�A&V,�yr�	n���:!�(��(0nG���	cX����Um��	��I�
o84 ��%D����c��� ��D�gS��y2ǞK\�1�:�<Œ����y�!�'<)N�zǂֈ������y��(2��ygk�l���!����yj
�y��˟�ZɎhc���)�y��/��p�P
Ń�*5��E���y2��%�VTQ��(f�0H���yR�[�2�. �CB>$'<�3gN��y��ӕ
�(;�
�#1rhɆ,
��y2���+-J �P�&�5sF*���D1�O\��T �_��QEJ�,�*u�#*O|���%��G����g�,p����''(��國<,$�o
�aŌ ��O�=E��k�<D���1��Q�>��@Ӧ����y�چ<TB(�#�Ԑ0�"���`��'{�{R[$R���N��t!�} ��E��y"h�I��(;�W�d�*�
�(M�y� �82�cFD4�r0�2�� %�!�$�![bm
2�P
-I�=k�?Pb!��cu$����<:�y�4��[=!�q��@a�3 ��T�R�D=!�$Y�vY8����@�$���J`�8&�!�[	-@���
�8��R�2c�!�S�K�-(u�� 2���Ⱨ��!�$�Y�^5!cB�Y�jYc1F)4�!�Dȿ0�J�`��W5x܌�aD��	�!��$����q�+;rd���� \�!��b7T�"w�(sL6r�@{�!�D�!)�t;��y7$a`�	_�k!�$;�69��mH(c*�x׍�X!�0P����%�3������^�RN!��Ԝ=�B���:�(	D
�C4!�D�󾁛�� ����gHS�m-!�)`�8���8nW.��4	I!�R1F(x����#?�ؘR�˴7l!�$�(��<p4$K8-����ȩyd!�$A�� l�� <���ݥ�!�d���9G�W�b�j���ƃW�!���^��$3�	�whf4k�-<Y!�ʓ/@@�y����gp��1MA;8�!�$D��@��.f<��0����!�d��%�����j��;2�ٳj�V�!��}ŀ�+�S=.p"vi�$�!�D�6�0�f_��`sIC		�!�DN�vx��"c,۔�6h�o!��_�h��!5�=w7�؊�4�!�� ȤP�*J�/��$ء��/>M�b"O ���Z:!��]�ǈW�mz�jD"O�8���	�`'�j�Z�Q"O�5riK�X���(BK��HG"O^����@����CA0A������'��'q�'��'��'��w�T:q*ި?%�9SHB=
D�A��'���'��'7��'3b�'N��'�ԑ#���UFz�b��s�@1R�'���'�R�'l�'p��'���'���Ȍk6f��f�7��5�C�'>��'p��'���' ��'���'0��TBP'E��4Z ϖ��Ĵ��'Zb�'��'��'�B�'�b�'T`��2n�<,6м�s� j�rx҅�'���'���'��'�'�"�'�Ta� �7,�N[�l�T�R�'4�'���'r�':��'���':H ���؊T{���K`���q�'�b�'�R�'�2�'3��'^b�'�P v��"h6�R0�@�=Pеh�'=b�'$r�'9��'���'XB�'0`<�3
޷I`��$���' 	�'���'"�'7��'vB�'-��'�r�cRJ�j�\57 4���'�R�'8B�'f��'�R�'��'��͑V���/�^Q����:2�����'���'��'
��'���'�r�'�u�w�B1�~m� ʳc�ؼ��'���'u��'���'jj�>��O�8!A5�4�3r�>EOhi�g��Sy��'��)�3?A��i~�\�tΘ��W-L�`���K���$�ۦ��?��<��]y��!�؇+�	����@������?�w����M�O^�
�"M?�h�՝o�z�مL���ʥ�9��̟�'v�>��u�@�Y�t`�� 3�y�4bB��M�"�X���O�07=�G��r��s2)W�3��Y`�O>��k��ק�O�~Ĵi:��8=��0�gJ5[�>�Q�cF�}��{�P���%>d�=�'�?)���8�p;�"S&NN��e@�<i(O:�O�Lmڱh�0c�0���!��x�о.\B�	\�4�?��X�0��ߟ�ϓ��䒟+_�y�%^U��YUؔl�I��P[��L�)�b>QS��'�X�	7�Ќ�ءX[,!�ߎH�ft�'��Ο"~ΓMH�8t`->�>E:��7����`O��K�?��d�Ц�?�'���ˌ'.s)J��I�+y ���?���?)c��M�O`瓞����T.$��Ԓ�,A������YN�O���|����?���?��K�X�����z�3'E�?"V�4-Ofam�!o{��';��陖6ւ%� �����@�]�w��P�'��7M�צ��H<�|����^�U+��l�
��t�R8�b\C�S�?�f��L76�[���5�u�d4�Ky���9u��z��<'3��;Ӫal��'�r�'��O��I�M���0�?qp".o���{��i��!�'\�<��i��O�]�'�h7�Ѧ%�ɣ!Re`i�)��7!�"a��d�C�:6y��A��(L� :�"��u��'c�D��4��2b���H�Y��كk�+#d��Iߟ4�Iן<�Iϟt�	c�'���X�&Z�da+/�{������?��u����5Q<���MO>I�aנC'����j�.X�*�� �'��� ��=����(�n� *�����#i�-�&��PrlL�r�'/<�'�X�����'hR�'U�Qf����P���d�����'�rZ�<Z�4g��-���?1���>,<���'͚����@�PPG�I�����O��d)��?A�ŁHW;`k�	��J�T	��B�4^r��H�Ǐ�S/O�i*�~2�|�̕2)����R"V�S��M����'/��'����Q�$2ߴ:0��Ac�$N��$I�b*%�*�?A����v��d}R�'+j�b��W�y��R̈́1x��)S��'xJP� ������݃v��'��D䜑 A��a��+:��<)���?���?���?�*���؅@��ڭأ"	aΜTsR�Tܦ)s
[��`��џ�'?I�ɺ�MϻC�t(��㘔&�P��0;1d%;��?�I>�|B��O!�M��'������1���"�NJM6
䡝',��cj�j?�K>)-O��D�O�]�'��<lJ��'�?�FY!��O��$�O��d�<1��i��s�'"�'��P��&�7"<~�JQ�U�Gل=�c��s}��'\r�|"A��]I���+X�<(���1��$W)���(H'f{�������c{&�$L�U�1qS�G�!�0H��@22oZ��O��d�O��D*ڧ�?yb��<+9�����<~����bD�?��i`Rq��_����4���y7�Sfv�����i���r�ƅ�yb�']��'�f���i��iݡs��E�?y1Un�*��5�4��r���a��ގR��'��I��	8�	���=01���F��1���sQ��JX�m�'�V6M3vfN���Ob�$7���O0�3fٺ ���kĩA�>Nv9#��z}��'�2�9���F���%n5>\M��C42����-V����h<��'���'�4�'�Hbh �`�Qzd
��LI��'�"�'�����d\���۴@� Y�wD�R��W)w�����"��=�I������j}"�'���c��� ǐ�t�ñ��	��t�4b�	,'�6M8?��!�r>��%���� �=b@'�RWlU��EΝ
��� �1O���O��D�O����O:�?��akV�W�A:e�ϐ� e�������	�0�ڴ0?蘨/OH�nZA��0>`VƖbC�A��̦$+f\	K<����?ͧ�b���4���2e�GI�'��iHS�?IV��@���?B=�D�<�'�?!��?��]&k��pj"�P�s�~8�W`��?�����DWӦ!@	����	����O3m9�K�0.y�1�!��3vh��O�Q�'j6m�㟬'��,���95IO�2���ʊkkj��R�ϜA�~5[�.O���4�E���9=D�O,�wǋ`���9�@�R A!�O��D�O����O1��ʓ&Û��ɝ`7 �p�j��zv�)ڒ"�g��, 6�'��L�Z����O:mmZ�L���3��M�����7HȚe���M�"ݲ�M#�O��I�������<a���C{�#�G4+(�� %��<,O����O�D�O����Obʧ2fLR���
@���j�!L&�Ȣ�i���8�'��'�O��e���B���qqe�+Z�"!��Ǖ�,�D�O��O1������b�f�KG�$��Z�zek�K%X�扢-��m�U�O��O>��?I���>��C?����׺'Xv����?����?I+OX�m��u*r��ڟ��ɢQ�d����H�)��� �Z)�?��S� �ش0<ҝx"�/:@��L��`I���d
5<@y2��4�� L)������:l+��ՈG/���t��;z� ���Ol���Oh�d'�'�?�t`NTժ��筍?mr��P�A��?)׹i�E�'Q��H�4���y�@�=� �6-��Mq��W1LvHE�E�����O�7���L�6m ?a��P1Iu\��^kb�X���X(tӂ)�.l9� �O>�*O��d�Od��O����O������V��q
E�^%�邷ʿ<aE�'w�4���?������?a�ΕG"��$��UJ=Ҕl�$L��	ҟ,m�$��S�S�JM"i4��D:�I�!�J�gĨ
eL��F|j�+�z��5*�O��JN>�-O�ѫ��W�Hea4�pX����H�O(�$�OR�d�O�I�<yG�'�F4b�G	$�$h�;�z�!�ӑ5��-b������d�`y�'��FaӺ�ZT�Y�$�`�v�ҟ&=2A����#�07-$?�)K�$���(����cǋ(SӼ�pW���~�4�$�|����Ɵ<����������4�4"`�T9w��'D�H�����?)���?QƸi�V�Y�LI�4��;�&Hi��&S�=҆W�d�JT�c�x�/k���oz>��� NƦ��'t�%�bm��3ԬKwf�5�+ԇ�5h��T�	�tf�'��i>}��ן��ɿ.Pz����R46�4��nC!ɤq�Işܗ'6�կ�,��O����|ڦ'�G(z�!�L�J|����r~��>���i��6�PJ�)R4�L���{�/���=S�g��D~�+�oļ<��5��T�ɟ�k2�|2�ȳu�	!��95�vA�]+�`!��˟@�	�H�)�oyR�aӦR�Ӌr�t� E��F7�
PiU$[Z8�d�OJpm�A��HR��:�M[����h��`��P&�h5�6�U{��i�~i8�i���4e>F�q��O��I�'�t�3*[���P+i�ћ�'��	��������͟���H�t+�>60`0�EF� v�2ũ�Պ�b7��*���$�O��d7�9O��nz���sIƅs �9&�ٓ�.�rq�G������Ş59�Y�ߴ�y�e�yL�1���+ң[D��̓'k��('��O<=�M>9/O�	�Oĥ���Y� m䅓��*J�� kb��O����O��d�<Y��i ,��T�$�����)�(�(g�(YF�[�����?)�R����؟xN<����<�>bp��,S�hBFI]~���=�~9��R���O�z%���'y"靬F�� ��fj$4��T�$�b�'�2�'������)L�)�th�G��� ^�@���ޟH��4U�,�p��?�i��O�3g���2���G"�YJG����$�O����Oj���{Ӹ�Ӻ�E� �"q&V�#k�� (�d~��q��^ ��O�ʓ�?��?����?��,��CGn��� V.�^c>�2+O4o=j����I؟��	u��؟Hx�ł�A\�T	ƯÜk��r@`������O���5����P9H��PAG2lp�{5��	*����.��#Ē�����O$��I>�(Op]��L�<�u�ր�>>�q��%�O����O����O�i�<�!�i�|}���'U� �.ۜt+�d[$�'X't1q�'U�7M%�I���$�O����O �aP��SR,j� a_dCt���ii�D�O@컃�����\������ñL[4Gd��8@gɕ1f.Q�6�s�@�Iޟ���՟l���l���.��D���; D RȽ�N
<�?a��?1��i�칈GS��r�4��j���[�a��ɿ?�F$�&�x2,h�~���2�3Q�s�:�k�r���SB�Ub�Iօ	����db��K$��P������O���O��$)
�fy� 9v�����,v/���OT˓����Hj���'7�V>�`V{����A��m(��)tb"?�]�8!�4f����>�?aZmG�i�����Zo�������v��A�*.���|�c�O>L[H>)�%Q�fNʠ���V�&�9�@Ѧ�?	���?)���?�|z+OYlZs8R42c\�*2`��	�Y��"��|�	��MˌB!�<)�49�B�pv�)<��F[.#����i�l6,�7�!?)f�+2��:�� ���o�/����29~m<ORʓ�?!��?Q��?������/)����gH�Vn�����X&ML��mZ/e�� ��џ$�Ie�s�Ĺ����6*Ul�pq�K1A0*���}����}Ӷ%�b>�g"M��U�c�Be��Ǵ�n`�׏�K3>X̓H��L���OY�L>�(O��O��P����%[Jț��̌
�Qf �O����O���<	$�i�&(c`T��I?*��db aX�iH���2����?�#R��j�4��&9��ѥa���;QEM���`@�*>i�Ɋ���jK�;Ts�b>�z`�'|�8�	+�z�S"�(2�t1�� �֙��ퟐ�I֟x�	N�O!2+O�~�DrW�T$Kd1�$�Ɲm��Im�JAv	�<9p�i��O��:0'�({�m�4_ʬ�2�@�?�����ڴ6*�Fk�n�Ƒ��Q�`҄Sx���Y� J�RlDAA�"��
5�#�D�<ͧ�?����?����?��Å.]����i��G�����ǧ��dV����J�� �Iԟ�'?�	v;�L�q&ɪE���hPʊ�S��O����O,�&��Sݟ��ӌ;*dTR�nߥW��C	��@�B�Z3�=e��|����O��L>�-O�}@��P/Y��SUgW�
��U	5��O��d�O��D�O�<ٕ�i��C�'f���'��FFU�"���U���E�'��6M"�I���D�O����O��tb��xࢀ�M36���A�R�D	.7M:?���
-~|�]��ߡ�Q��'G�}�vi�(!|ZD�Cgi�T�Iҟ���8��П��j4j
�C�q
�KAoj8�����?Q��?�$�i��ы�O B�v�0�Oj��Ѯ�Jc7b G+�+��&�d�O��4�� �f�0�Ӻ;�.�SlXB�/Z��F"^�nh��(n�O���?q���?q��DȺi����BA�ao��9:|�����?q)Oj�mڱn��m�'?�W>�[�덯؄��(	���I[�h$?)�V���I�<�H<�O�����b�ay7d��jB��� H�~[:�;�Șj�i>Q���'X�	%�Tpn�$th���S	ΆE�e��Iܟ�����b>�'S�7�H�(�:p����
��Q1C��k
��V(�<	��ij�O�Q�'i��DUH\�T&R6ɴM��$F|@b�'$��x�i��i�尤�T(O��Dґ]h=�2%K*y
�Z�;O,��?����?y��?	����)��v�(q�@�:fA�!)2g"x�~�o(�x�������_�s�<1����d^r��!f�Gr+(��`S��?�'���O�,L`��i���B��py�,�����uj:(�d�z�ޭ���Z�D�O�˓�?��.�d�D�����f��&b������?���?Y/O�1n�N{�)��������Cr�@D�I��Y�S��V�f��?Q'Z�<H�4P�b�x�*S&&� 1j�c��y]L�p����D�,N��`#�9�Ɠ������T���1k�1Z�Y1I�NL�T�;����O>���OB��%�������^Mr�+�.N9� �ah��?"�i�MЅ�'2�xӂ�Or�4�h�P�Iħ��ՠ�oF�"2O��d�Ob��Bc74?��9"Ɯ��'��$J_ni�X
W�Q��F�[�$���<1���?q��?)���?AV����͓P�B!Ed M`������J��3�L�런����\$?��	wbLɁ)8k��5�&��+�� �O ���OXX%�b>�C��mR�m�B�O������`�F��e9?�e�1e���D�2����ʉsqٳG�B�U�y	���*A���$�Od�d�O�4�V˓r��6IS2�� �(YrB��<�[�'ۑ�y�@c�X�袨O�$�O}mZ.MOJe �f�>���K��m?ƍH�]ݦ��'����
�?��}���Y�n! �mQKR]!�	�,3���͓�?����?��?(O1��1�@�S�!P_␐%���'��`�tq��3��ć���%����� �
����@0Q���D����?���|��N�M��O\	g�J�4Y�]�F#.�>�3Ї�nn��p�l4�O���|"��?��{����ɛR+�ŭآ��ؐ���?,O�o�d_�t�	�����M�d �d޺�Ǭ���� �BQ����d}��'f|ʟL�Qt� ���Q�<n� ����h�L�J�gV �^��|����O�(3K>ف��j��#r��tȾ�x��۫�?���?����?�|�/O�@nZ�g���2��<R�P෢�%�,e�Go����I+�M�����>���"Xr�(W�-G��q��A@7He+���?��.��M��O��-M����@��P֜h��M�$v�ʸ��Q� ��<!���?��?9���?Y-��,�m��@�xzG�z��A��g�7m��i�ʓ�?�J~��Wԛ�w���E�*��Lq'�� Tp4��P�'��|��TeY �F2Ox`��G\�8��u ��D�[��z�2O��[A�ه�?�5�7�Ĺ<���?A��P�s��R%dD3-*6�T����?	���?������\�ݒ�Fy�'$�Y
�"֮er��1F(4�(��DUA}��'�b�|�䘒I�`R�iH_k�X��'��<�e�ƼwyX��p��d�������'��M8'��y��	d8�Q�'hb�'���'��>��I(RD���<7����=U"�����M��'��?���
��6�4��-J�M��$
�]�`śc�00p�=O�o*�?q�4���r�4��$��~�$< ���� z�p�P�[H�k1�7)��'�.�d�<����?���?����?�HB">�j�����aLx��H�#��N����ן��ݟ�$?�	\�JX���J(rB���eό�M=a��OoZ��?�L<�|�����X7ސ"o�A4yf	q^�v��'��	9L\�)��7�ʓOT�`�!�-�:���4	�~������?y���?1��|�,O
mo�({�ןh1�V6(v<�G���D�5�֟�ش��'���?1�'g�6J9`8���AD��ɱ��ҕ!arqIƴi�ɖJm��
��O�hp%?��݃Y$��Z�Λ�4W6˖�}~���I��$�I˟��	o��d\��gF"|�, #���|j���?������͓�C��"�M3I>��cA�=���ӷ��;^�8S�a�M<�'��>O�tL�_�����`�#��g �=���,4fXz�:s?�`��'�(�'��'���'���'�Fh�'��(g�	!��W.�	�e�'I�W����4��S��?q�����=���J6�+NzFq�JN�������O�6�m�|���I5�f(RU@�A�N�@kB%)X*T�5C�-n:����*F�H�3�|��B��$��[�+̽Ȗ�VF���'j��'7��Q���4T#�ш�	�<�6\��&rb�A�Q�?��E�f�D�R}��'{B�kw� b� jש<5���'O6m��P�7M(?ab �p�	5��g2l�$d��J���CPK��y_���I��l�	���I�H�O�T�2��	+7:��#�-^'{�%�IlӦ�����O����O�������������J��N���$ϝ `E8���㟠%�b>1�����Γ+���3���!Maz����������\lj4F�O�8pJ>q,O����O�ܹՆ�?:�����%SZ`!���O��D�O����<I��izQ��'��'�|Xä��yⰰ��N���1�DV_}��'���|�)ՔB�m��)μ*0f�sE��!���S�TU)0e���F׬���P����'��\�Q��"}4���Q�H��(i��'��'2�'��>}�ɋd�P�
�N�dz��뎐&L�����M#��
���d����?ͻ�4]�`��Hn���l�Z�8�ϓ ��b��(o�8�nK~BGY�7��m�S���� G�Ѓ`�����JECR]��|�Z��ӟ��������������)~l9aw�U�O-�LXf�HVy��t�B)����O����O�������5i�`D��65���s��70���'\�7�Uɟ|'�b>��'�-UR )s��O��}��'F�
.V4S�e�`y�%��,����]��'�;LJX�KgV�S'��s@fB;�@L������	�$�i>%�'��6-�؍�OBG�Ąt�vP�"#G4H���3O6ulZL���I�M[��'ƛ���i �'�"�`lY`���C�i���5zd�p��OH�$?���5R["m�uބ|���T�h�(�֟��	����	��	B�'b�Z�c�b�Vl>���g;�.ON����)r� p>5�	�M#J>1A�V\���(� C<r����A&�'�z6͎ڟ��ތ07-7?!�Xv܈�L�K1����h0+�^��U��O���N>�-O����O��$�Oe��B!v��q�pL-@�,} ��O���<�v�i��{�T���	g����Iɲq�V�@�8t������Xt}r�kӴ4�	v�)� ?�m��-Ӂ�\�����	b�!���R�&�+O�^�?��'�_�j<8�JG� <VY��cԔ%�P���O@��O ��i�<��i��!⡄1_^��ԋI%ڞ�d㋾"��' �6�;�	-����O&L�ց��RbXD�Uh٤hZ*���e�O���Ҽ{�h7-,?��ebF@��O�剚3/�|�����o����fΌ
�@�Fy2�'b��'K��'�P>�B�+��(�B4��&�sݲ@cW�=�M�"G��?!���?�M~�2⛞w>�p��+T�e��t�q�[)m�����'���|��TmVx��7Oґc�iU�-ό8� d��H��eڠ8OPի��#�~��|�T����W
�=�,��r���t�/���������I[y�Gf�\�9�ȭ<������a J04脹��Pnrv�؉���>���?�I>yK��/����;'�9s��^~b�Aw��$2c�iAN��|Y�'����.8^ZAAQd�5o�:y8B��#���'h��'�����aF�Lu��X����^:[GmFޟt�4[�u�)O�	o�U�Ӽ�I�6 ���FI=S�\�Q�$��<��i����y��܊��{���R�(��d�i[���(~�Q(��M76��b	�+�䓷�d�Ox���O^���OF��
 
l��n=z���[�L�A��˓��ƌZ/`r�'����T�'�ԙ��a��j:�ً6L�(6�E��>����?�I>�|Bb-�"���Ed��Q�f}Ƭ���T�8Vo@0��d�F2�k���r�O6�&�y���Җ?ƌ0�	1Q�� ���?Y��?���|�+OP�o��Y�D<�ɖ<��Y�J`V�A�4�դG9"��Mۋ�ɷ>����?���i)�xs�
�(-�|2���NGx}2ύ -�����U�D"�������0�D���T��J���8��1OL��OD���O����O��?�I� Ѝb
(��-Ն�x� ߟ��IӟT��49���+O�]nZW�I_U�� A��2�V��a��(W��M<	"�i����O��%Z�i���_o�� &A�W&P�:YB8��(P #���$���?��-�$�<I��?A��?qQ��O[�D�-��N�䙺��A��?!����$���Ձ��������@�O�y�WKZ|E��yC�ޖH�m �O��'A�7��L'��e� �u�;����Z�.�V9J���\*���*Q���4�n����AY��OR 4�%f�8$�%P�M�=4��O��Oz�D�O1�0˓7 ���}�r���T(�x�25i\�j�,a�W�'��Dv�4���O�]n�=]�(Pa��0<3��PA]t]����Mˢ_�M��O
���A�*s��<IWM��F�µBI�'���T�<y,O���O��D�O,�d�Ov�'y�����ױH����hE'����iE\�3&Y��I~�'}���w�DX˄�E"s��hІ��O0S�odӰ�lZ���S�'u�4�9޴�y���Xfn�`Ɛ^P��`+�yR��p��	
��'r�i>��I���W�*h12i�88,hu*���O �D�Oz�D�<�ֳi�v}���'���'�.(�L��ڍ*D(�c��Z��$�c}��'3�;�Đ�`�u�%��[˴ݑ���4j1����ѻQ��i�b>��!�'��	h(h!���F�6��%@�.X<:�L8�����ɟ���_�OR��N R�䙣A�W�f����EhY-;Hw�8t�,�<���?ͻlzt�ԍõW�d��cY�&����?y��T>�������f�����A ��$�ãsq����mA�M�2�rը�%k��8&������'���'���'$�59��H�E�Z�@��E6�9�WS�D+��6)��	͟��g�͟T@`oݟ���iG�2	�q��O(���O&6��\�)�iS����΀�)�h��H�!z�����/L��I�#�|�'��$�t�'R��2�-��z�b� 􂐕l�h�e�'�R�'����_�4a޴0V>����u�БҤ��i�dx0��0��QH�uC�f��KS}��'��c�$9���.Z0�7��2�j|�Ҁθ_��7�"?���AC�|�i%���߅怞q�<�X�뗺��Mb�e���	ڟ0�����ݟX����i�n�qE���H=�����?����?��i���[�O��@o�r�O0�������N�P�\|��g#�D�O\�4�*��T!mӦ�Ӻ��J�S�
 ���3[�����KO�_�P*�'��'[���t��ʟ��	��6�s�L�gl�J%�ۓ��@�	���'	�6��|����OD���|�b�
L���Z$�ĝ�I#���<��y��	��M�q�'艧���O��4P"��4oX�p�f�&�9����%i��a�Ŋ*#�I-�2SM�OBTQK>a�mų.:yං��;����3�?���?1��?�|
)O�UnZ�9��m����i6l#e!G%7�4�� �������M�L>��i��I˟���,K�ߒ]�Nd��o������6r.��oG~Zw�,4C2ٟ"ʓўa����:-N���!-��	Lyb�'B�'}��';2W>��L�[TQh���?B�����C���M�L���?���?�M~�KT��wq⵺� -o��̫��0c:2��O�6�TQ�)��ߺN�T7y�`A�톼6����₯s�bUK��q��k��;)�(u�Idy�O��ܳN."���}n����%��1n��'V��'H�	��M��>�?Q���?�� I���`�/G��t�E���'6���?����?��<�%F�WTI��`Xx���'�����O�4��<#p��䍏��#��'a��h���$���3'�8,v����'`��'K��'Y�>���4_^~�f��#	�E��O]:&�}����?��d�dyrvӄ��)*����!$��|��QQ\)6��I�h�	��Ms3�@*�M��O�,Q.���NQ	?o��k!"�/`ެ=!�lE+�O���|���?����?)�!�����ٟD�d��FS14��*O�	o3(�(��IԟP�	a�ԟ�*C��W_,ZS��a�� ��e؅��d�Ox�D ��	�!b��qk�f��Z�T��t�ponH�+�P��wt�q��OZ@�H>)Oh�(�ʁ�_t��)�A��A�Q�D��O��D�O����O�<i�iz���'�]�FdǯCi��A�@?� E�U�'�j6-�I�����O&�4�����&g)�D_.21�)�**m|p7�+?i��Ϫ~�J�����'�����Ĳ/�~M�䋓�OC�D����<���?����?���?����%U�N5J�x-�V>�p"s�4~^r�'���cӶ��?�l������%����V��q��:��Ԓ���q������i>�a�'릙�u�Ñ��<�V��"�"����7��i��'��&�ȕ'�b�'XR�'Q�	� a��p5hūK�$�v�'UBS���ڴm�e���?����	^&Ѵ%#��Ükh)��BR:��I���D�O �;��?I���hMT쐳@� ?R���CxC�h9�@+9�)�������,H6�|rD����R畩G���G��)Eh��'ZB�'
���]��شcJr��G�
?Є�q�#�n6����H��?���H6����N}��k����o�eX��[�Jڪ��a��tl[dpoZx~�C<,����m�I�q?a�U
��4�b20��9R���IGy"�'�"�'Q��'��\>풑�G�"�@��Ô�wiReؗ�G?�M+r�@�?���?�M~���V���w#��*r�T�p2�	�7n�I-dI0�'��|��$D�J���3O� ƨ�s�4���e�(���R�>O��9P��~2�|2X�H��˟��w���zvL ���G�c��)�g��ǟ(��蟴��Xy¨w����#�O����ODD	Aܟn���A�������l$�ɰ��D�O|��+�D���D�;2��"��S���vx�``�צSI~*р����I�!��y�MҳAiТ��D�x�Vy��ڟ�������O���[a�AC�b�ȒO� ��)��G����(<��'��7�0�i�q�a'U'ZҰ�	�Ǟ���XH��|�t�	ϟ��I
��n�d~Zw�d@�ݟPȢr�-Y�����XD�p�V',���<���?!���?���?)H�Z6�X1o
�{(F���#����P0�՟��I$?��I#�&�"F�3OoD��+I (p�C�O��$�O�Oq��t�T.Y�m¤q
d`ڞ~��{T,� ~�N�<A��ңg�T��p�ryM�b�peKS%.{�P%BT�G�gr�'qr�'��O��I8�M�ᡑ3�?���C=j
�y��:l�b��	�?IC�i;�O�)�'���'}�o��2����.
�W�CoR"	�����i��ɼI�$ȓ�ޟN����.ѱ|�6��iR<=��`Ac-�D�O����O��$�O��d7�S]�Ҥ�eG�T��� ��7��t�	�@�	��M����|�|���|���t�(B"̳|iv|�D_�4Z�'����$�A<��&���t� H��ŲX�VȘ S�J������@���|�^�4�����	���)�GNRB8�QE��h�J� �Zʟ���qy��m�"�У�O����Oh�'(1&����0L۱�ɨW5p��',���?��4*ɧ�	�9
3L�36�2J� X�Q�X�:�V�s2ȟ%��!ۤ���S�>LBIYD�	��<��7@G57a:�I�ō����I㟼�	؟d�)�Qyb�j�)�r�"	�����5-2
X�`:iF�˓ڛF��u}2�'�L�E�a� �E;
{�!v�'B��F9Λ����ݣa������ݪJ��Ir�I�b���"�'���<���?���?����?i/�V��b�	�+��� �Oʘ7(�1�����p���O����OT�����;S����rF�6iQȕ�4��$"�8�	�L�N<�|��$G��M�'��-�d刃C�h��f�_�F�dy�'U�P9��F�Hk��|�Z��S�̊CMP1ms���$W9l�DX*r�� ������	cybLr�C���O���OV��We�� r�}ò	V��؀N$�I:��d�O��d6��I6���f��z����ף��|���� U��#H~� Ʒ�4����F��5���?�aY���:J�Jm�IΟ��	џ���Q�O]�2�h8�'�@�⠚Э�
8�B��>m���O����ŦE�?�;�\[��Õ���a3#��y=̓�?��22��O��ƞ�����޹�t�ڹ}Cԕ�¥ŭ�fܒT����'�Ԗ��T�'�R�'lr�'U��Sv��C<�����S�t�����T��aܴs|��+-O���'���OjHP@YN��1 � �3�@Z�.G}2�'�� 2��I4�ڰ��C�U#%��	U�k0�Up���?��ɪ�`����'p4u$���'A�b�L�!;�n}��$my!A�[9�?q��?���?ͧ���FȟX"DN�OB�����1X�0E ��g\ �Q4O�$o�@��i��	��8�I*�M�5�X�\f�̋��@�*���@�Ɛ.��U��4��d��7CH�����O��d�h��ꇆ�3ð�01��yB�'+B�'���'G��	�>�A�2,,�qjy�x�$�O��$
���r�Hu>�	3�M�J>a�ÐFh�[g`�Z��X��O>v:�'�*7m��	C�	��6�&?q������*�_+�P4��z�|t�q��OƬ�O>�)O��$�O��D�O�ӵ$K}�܉���s!(t�d��O4���<�R�i$�S��'qr�'��p�bvaC^Nh�j��C�z���R��I�M�P�'͉����qX��� �N�C�@��l�N�ʆ�T�6lH�t(�<ͧUr����!������uز=��1��F��FD����?���?A�Ş���N��@�5PPd<K �/X|�x�*�w&I�����4��'�8ʓ�M#�`'-}Ƚ���Y�	�K',	·i���C�i��	>�^LjB�O��'�n���b��ʽ�q��(S𑋛'/��|�I����(��Y�4`�3)���� �azt���²%E7�Ž4���O��$!�9O�elz�]�c%Z����w�V�{�d���͟d��Z�)�Sy��oZ�<I���7��I��B�p]Mkth �<isΖ$S(z�d�4�����O���E�^J���,^�br�G���u����O���OF˓����������J�!��l؅�(k=�I�A�c�~��ɟ��	��ēa>��J�Ƀqٴ�3vnC"tz%�'�07�I-mA� ���T����!�'�@����V�I��,4�P����'F2�'��'��>��Ɏb3�R$BQ�#�n��åO9]j����=�M�d����?9��G˛��4��}���K�-I�r
��h �)B3>O�Pl��M�p�i�4\25�i@�Ʉ+� C��O���c�Hkw��%.
�q�PCG}�Jy�O
"�'��'�2$'W��uDE'>� i����'e�I �MsgX�?!���?qJ~ΓdQ��K5h�>hz1�H�A.:t��U�t��П,zI<�|bBƝp�? 쬫���'�X8�$R�DV�Ś���:]����lӬܛE�'�l�$�ȗ'�NE�!.��w�:e�� �%$:��`�'��'XR��t[�x�޴PSRu����,��#��I��"�J��q���g�V�d�D}r�'���'�@x�_/�0� �I�
��r��/;��v������݄6��<�����"��^�A�v��SmS�\��1xv=O����Oz�D�OJ�D�<�|*���(|�p\�Ä��mL��� ��0�?���?�D�i�p��5�4fB�֙|2��"ov Q�C]Xf��9���a��O���o��	ҡzL*7m1?T �rb`D+$����p풯. 7�h��|BR���Ο��Ȁ�+ȞQ��lʃ�V@ihb@�ʟT�Iay¥`����$�O��O8ʧ7�~-�g�T��<
�b�,�2@�'�듌?y����S�����T���֥[�x�Ӫ��BL�iY@-�=3ě�(�<�'o���	@�I4i ^��㗙o������ Y+����ܟ,�I��h�)�{yrIs�@M��#���ૄ~>f� >=:�LH�F���Q}��'�h��������2�W-S�q:"�'��ѐ%Λ���֝���������*�j����Ϯ@��|�E!˕*3�Ķ<���?Y���?	��?)+�&|PtE�?'���H��B��qQ���զ9r�a�ڟ\����P$?Y���M�;G(̭�%���1b�re�RM�9p���?	K>�|z*��M��'c����3L�����D �V�Z�'8`T�+Ο( ��|2[���I˟t�d�
}�DX�i��/G�-`������I����Ly"Bv�"���Od�d�O����N��=;މqӤ�,��"cd.�ɭ��D�O���?�D/Ljx5��dP�VR��H�o/�I�by��:��@�z�(�%?�*��'�(����������|�`$�݆k�y����h�I��\��K�OB�OM��%��g^BLӖӧq���sӼ<q�L�O��Nܦ-�?�;+F`�[��!	b]���J13@�̓�?���?�sf��M��O�A1���']����O�\i���q�U��	��$���<	���.K���[J���E ^BX���O�o��z�'E��	?3�M@T��R� ʀX���'Eb�'ɧ�O���`�5;�J ЂH	��	�n��O��uk�^���F"��0�r��h�I~yr)_�F�ֽ����<~X:�@�(���0>�P�i��`�4�'wB���C)(�n,�gH]0[
���'�$6m0������O����O����/ºnA�W蒽.RƔ ��F�J7�'?	S�7h$���Z���cU(E�5*�5¦�E�&v	�G	�<Q�j[H* ���e$X*c垍(��.O����Ǧ]��5���i#�'{���6-��T�
hDɀ�5t�!��|B�'U�O>	��i��i�јV	�Z�ް���X74zE��ͭ}��������'��	y�����R�i̿.���W�Z'-0�Gx�!k�JT
"˥<����IX02Z<�ƞ1t��� 9�������O���%��?��c��4T��q[#@�1��ͺ;�H1 `�ڦ�)O�II�>�"Dؓ {��  �EHL�d�$��V�E#7k\��Z��h��oΙSB �� ��?��-!0O����,X悏�fu�`L!�|4[��)��"�Q���r$�1�?�wH�D6{���J�4�Ԁ��o��$��#�*gg�1�B$׽,�a�L�s:|��� PZ�+�L�!��[t&�<K?`Q��"ڧ���y�C�OY �!��ƒ�юK/4�$��S��8���
����s�0qP�+��2�.�����7��<����*�|0J�m+�	�S� �%� ���'�B�|^�ЈLټiɖUYt �&x�U�Ы@�axc���	��	UyR�9I �S9F���hS�f�ZT��f�%3'���?�������S�Inب!��hQB"�13G�h��^�$���@�I}y�Ȏ $`D�6�a�hɰWa�$�u&ʌie4�r[��7m�O��O@�L�t��>��g\O�0li������,��Q��ʟЖ'��)���(�i�O��iX�v���AN���K -E�nu�N<�/Of�j��~�qg��*�� �CD�(cc�!���_ɦ��'"$}�`qӎ��O"�O��� d;s�3�
�)C�ĎPlZ@y��Z�O��,�K1&έza�A�A'��n�0�úi�*���Bl����O����>�1�Ԅ"��0!��%YNn����Ʈ4��� R��O>����Δ�A�Z�l�X\`��`E�y�ܴ�?����yr#0k��'V��'�����p����D ��֪^C�:c�h� g?��֟��	��P�/$�d��CE6kq��	L(�M��'�ج�P�x�'a�|Zcu2E��Ă��<:cq߼��O��V�$�O��D�O�ʓjN0AW'?"�D�:sk9k��ɑfOv�'���' �'��$;�ȑ rA >69�Ee�&�xe��1��ʟ���ğ��'����k>�p� !�:x"��W���p��=�D�O|�O��^�^��'�����b�1:�~8���k���8�O��d�O����<q��3��O�<I��)N{pܸi�n���Kf�m�0��&��2O̤��+�D4�r3O�*��ʣ�i���'o�4P��M|�����K�${Ƙ���́+�-�3�/
5�'V�|
� Lua�C��0��P�%�h�d�i��ɜX�x�j�4�?I��?��';�i��Qv�3�`my��X(&��7�v�l�D�O P91��O��O>�g}�e��"�x��"L e��%�p	��Mӵ"Q^_���'�r�'z�D��>A.O�q�i� ~��c�a��.z@ȁ��+����\'�����'��vd�4v���!��A#�8�3�i���'_2�I�G�`���D�O:���X-~�2��e�H�腱R�@b����g�y�I����I��E/K�ɓҦ�+� )ۂ�Ձ�M��<,��@U��'���|Zco�}���Éjz��-R%n�聭O0�4��O�˓�?����?	/O>e�`H��ʣ%JĹ�\�1����'�Iٟ0�'B�'d��އ%7>��@"&�<\��7K�TV���?Y��?Y(O�i"uiI�|��k��>:$�b�ڂ8jƝ������'W�|��'V�$̈́z�����m�8�rS��F����͗���ן��Iɟ�'.�9�CF�~�m�4����-_��c
^%Wz�T7�i��|2�'�Y'c�qOb��
6�� ȅ�˪L\���i���'�剋`��ٯ�x��O��I>��x�_Kq�0���	v֌'�$�Iɟ�;s*�П8&���D\:!�#Š$���>H�J�n�Hy�+u�7m�ON�$�O����~}ZcK���D�x�����(��ha�4�?��d���Y�2��ֆ+��E����F�/>8�֧cZ�6m�O����Oz�IT}�W��Xl 5l&tI���k�y:$mB�M�`d���'�����,���kԃ'?����G�,3�Htl�۟��I�h�S#3���|����~rf�Lˠp�&GW�S} ��[/�M������?�*OF���Ob����"���0^��(Se
 �:xm[s�if� ��eBJO��O��O�,�!�b<T ��cҍ$����Հ�m�I��'���Idy��'ِ�B���'H�gڢY�0y!���4Y��ڟ���d���?��'E���*B#�4���ɳC�E�޴Bl��'�R�'��Z���].����1)���2��=S>�M�qg����d�On�"�D�<�'�?y!�I��ȕ��K�k�����ފJ�����	��P�'d-���1�i�"\�lA�c�G�xo¤�Q, �m����$������'U�'�L�Lʵvm&�j��")�	nƟ��'f�X�s'�S⟔�I�?�?*�0���F��8:�q��N�^��Ov���OF��e��9h.1O���n^F�0�I�6���I�KB�&���?i ���?��?�����/O��;����.@�9ݾ� EOU�E*�V�'2b̙![T��y������&Y*�1VL�0kl�8�ɀ�M�H%^ś��'="�'O�D�8�4�4�ĭ\4!.l􃰣[� 9$����Ǧ+3���$��dyb���'�B*��j���{g	B���|Dһ0��6-�O.�$�Op���\�i>�	U?vL�/1<��Ğav~��#g�����Gy���l��<����?���iJ��ω8U�D��$�V�-]�1��i���Ouz�O�I�O�O�Ńu��k�x��E� iD@�o�d}r����P�\�������CyR��O��,�e@ +H��A�ף�-c����c-�$�OD���O��?��B��,@�ʉ˱��)�\�"��?iM>	��?a-ODE�`�V�|�o�{�$ze5GzD��à\Y}��'��|�U�T��B�`���1^�8U�U*M,�*ܣ�J�ē�?-O����=xh�ʧ�~b*��4���2BH�(��q:�E��M�R�'��Iҧ4N\�AI<)��1l@A�4�ϖg�^|���٦]�	~y��'�H@�`V>��Iʟ\�s�y��#����K�@G�d��L�%@%�d�O���*d���J �T?m�̀�Pn��AK��hL�'�>1�
`��X���?	���?��'��J���TA� I�@�2u`��i��'�� �����O��z�<Uٌ �f�ՖG0��ڴ_f<�X��i�2�'���O�T듭��ӛ&�$�[�ԃ=Ҿ��E��~ mZ�HP��	ן̗'����X?jX!	���vǢ5KQ$�	Y�p�l��t�	���za.�����<����~�פq�����2_uޔ���]��M�L>���<�O�2�'�"i�[��%���³�h,��D\�7��O�x��C}BU����|yR��5��Ϊ#�Sa&/��G�J���$EU�$�O6�D�O����O@˓EN�`	�M)"��+��۱�����C�c�Iky"�'*�	���П`�I<��\�����K�@��l��Gy"�'\r�'�	�(��әO��d��D�v�ӡT�E9�`E�M�*O��D�<���?9��G���*�q��T�ML�"����x���PQ�����h�IGy�+��R꧊?��f�/m�@�����e�|ha�ߟj����'�	˟P��ϟpcw  ?��1�Ù:'� �gU��|����r�����O���0|��\?�������Sg��5K��΢|�հ#!Y�.n���O���Ox������MyڟV�iV��>:��bՈE)6�����i��I-BxHu��4�?!���?���6�i�e��-[�6��Yy%`�_`�� HkӴ�d�O
�=O��<	���F�U"D�@��D�SJ�qQ�K��M;1A�({k���'��'��� �>�+O,�ʵ�S�f��ň�BT����ɦySbm���ty��)�Ol%� ���D�w<�q�F��eC��iUr�'�rg�$l�6�����O��IY� q��K����b4j�J7�+�dM���?y��П��	�D�T�q�
���s2aȔtʖ0��4�?!Q 0M�	qyR�'�I��X�'��I�˿dȻ%c�e�$�u�f��?����?���?�)O�!��`i&��"vc�W�6�!�Lߞa�'���`�'��'�BD�\����@S�|�.��B G���+�'��'.��'��P�,�с����:;�޴�҃L.M,)ӒF���O��d;�$�O���~E�D��$�x���pJ�%��Y9(��'�r�'{RQ�|�iə�ħa ��s&%D6t���ar,��@�h��i���|��'�I��Mb�>I�̞2E���F��e~��h������ܟ�'n,�I�!9��w��ɜ�b<���'�8(�l��dd�"��&��������0ob��$��'V�F��j�>{��� �8��n�hy�J�82�7�l��:O��<?I�d�*&�= ��
�� �aB���I��6�R���OB�y��M������0����ش=�\��i�2�'���O#b�h�Q��*Q{���:*gJ� ���M� ��<QO>Q��4�'�Dcp���B]�NN<� �רg����O��I<;����>Y��~�">���I�b��&]��s���McL>4�S�<�O�2�'�����Apn�i��TY��q�d\�ш6-n��
�*Q��?�M>�1jKR�8INPh���8*�z��',�R��'2�	˟|�Iğ̔'I���B ��h@���))��rv�1_�b�X�Ir�	ʟ\��3*�p�!Sf�-�0L�e(F�xT�Ia����'���'X�W���Pb�������bB
�8|j"�#��$�Oz��1��Ox��E/,��d��Fц�٦�R�/
U�D�_��m�'�R�'�2^�t�`@C��'az;WlX�x[|$�d�**,P"�i��|"�'��iV?�b�>ArO\�\`%a�CGy��c�֦��	�d�'��E���9��O��I^3z �	0weُ5)�(@ËwQ�%���IƟ�;3�g�$'�,�'#N"8EȻ;�*	`�>dV�ldy�)Ж�7��H�d�'��T??y����p6.c��H�)�T j�̓ĦU��ş�[F�ʟp&��}�s`Z+w�UI$E�,c�`q�čR̦�����M����?���RW�xR�'�j����lcFQ�'ǎj��Ģ!�'&2j$�'p�'{���$F�F]!�	?qp�i�P49P�l�����	����b��ē�?I���~�c�lD�B,��\c ��]��MKN>	��i�O|��'��,��M���ܓmo(\
��9�&6��O>٠��E�i>yEyb��h��M�aL��9} �83�3�ē�?A)O@���Or�$�<1`G 6X��PʷnL�Έ�2��ϳ+g�dâ�xB�'ў\��z��X�-B�vP�E	�#*<��m���h�'���'��Q�`A������bV51��@S P�D�إؓ�M�����O�=i,O����m����5����\�˵�S�7��i�'��'��	ӟ���g�p����9a�#g{
%����`.��K���Ms���䓴?y/O���Ƒx��@�,����=M!�4�'Ϻ�M[��?�/O�1 Q��V�ß�S�,���˧�]#,U+Bߪ!�N;I<���p=��,@�j)�r��.{��� Ʀ�'�A�c&t�:a�O���O�D�*��]#dF�8>^6�Pb  F��yl�����}@�"<����^�NM1����8f��!��`��M� ��yԛ��'�B�' ���:�$�O�tJ#̀R�2wdѲX�P�a�Ȧ�0�)��O�Bb�7h��)Q� \ψ�2!� �
6-�O���O0՘��O ����䲟���f�D�s$�W9jUF� �d�'�Oj�'>e��Ɵ��	�I" ��n�-PDp��"b�zV�k�4�?���E]�'���'ɧ5�C"U�m`���+�d�If鏾��O
�d�O$�ĭ<	�+i����+eD�[2ed*�Rq�$�Ot�O�����
sΞ# 2ld�8y�dPiw�#�I����	�P�'�Da`��c>��`]�v���4�&4z �oa�>���?QK>����?9��A}"F]�x�.�� J]�A����#����O��D�O�d�ح����i�QjDlө%������P�C�.�o��� &�X���|Js 1�	�IQ�m҅�P��Lj@G1j����"�8a�|9��j �^n� �g?��S�0�F�b�F�gu(-���|�<�v>Ȍק�%+������Fo#jxa�M�tq�`��.ؽ#FtP�#��"���ׅ�:�����C{:���!H0)�@LW��,R��.U�ɣB��6����J_:eҸR��;$ ����I|Eer�MB�*����V�ِZJv�W�X#�)���\��z�J��=FS"��g�r��}���[�8���O��d�O~��;p����D��)*h���ܻ��hpċ	�3-}�㤂O&�m2�l���OI�'�@|�U��<�`��EЅp�8ŃA�ȏ}P��#��9�Y�t�:1؊����tm�'�y���6|<L���$��8)$n�2,┟�iRH�O��/ړ������%]{tm��)�t���k��i���N�Q����(8�v��'\�"=�Oh�)� ��ǥ�/F z��Fʄ
wn�$cB��0#>����O�d�O����Ϻ����?�O�\a�J��T���f��.���ʾ2��X�#�ߚ]�����'�v�2T��Up*��Y"NpY�땽w*�q�33"uX%��'-�q `��KW�D��HxC�!ѵ�Π�?)��hO �@*�%ʈc� u����E�(H�q,.D��"d��s&�(�"�R����0�I�����<QpÕ�}���䟼�A���1Q���sng�鸗�ȟ��	�E����ʟ ͧ>R� �g�6GL=�Tꀋ�M���%h�B��]�v��a b8�\��-�#G��ڤ��56��=m2�$ADʺ*� �c㘰(�����)�"�'��	>B�����]�xۀ(X��b�t��Ɍq��{7�'h�`� �%T�4B�	3�M�" �Z�x����2-���d��<i-Oޥ�!m�Ӧy�	��\�O)�� �'P,P{Q�(D<K�!�2p�X���'�B��*i����i�=���|Z/�j��͕�R ��#�ښ9���곘>����S
]���=����Ɠ�L��ѐb	�QÂ�
�>!�!������p��T��>]F(;"lרDXU�*M`$��<9���<��N~�J�@?/�h`B�H�T�3�����ޙ1�G�+� U����9k���'�2�'H�����>Z���'���'��dE
[^�'1g^�i&�\5<#�$�g�I����T=Z�����|2�X%Wq"��?ME�P��AҘ3,F�"##�f���`q�58��L>� �W8JoX0ȡ�]�n��"4���?1�O�hKE���t�	�'�pd8P��'��pAS�=NWdB�)b6�,a�H�n&��'GH	z�B�n#�����J�j���7l�X��� d]X�7L �����O����O�٬;�?����$�Ҍ�bH�C!��t��M��d^%c�vXs.�4q�}B
�(3�h�j@
�.�"���,�k�
�pL
�>�����ϣH����	1(���q0�8먝��*x$��3��OJ��;�$�OD�D:�	#OD� ���X}�����W�>RvC�/LX�)5'�mN���I �Rc�0�O˓EH�C�iJ��'��]Z& �+!s~y�a������D�'��A����'���0�|R�]#o\,kG?�0��۽�p<IC*D��s�tmQe�� sU�� !"�r�v���I ��%�� 8^F�CC�R*��Hh�fS|�!��,�\�
Vp��Q���y�!�d	Ӧ=S�M��zZ�f�J�Rt���s�1OȈ� 	�������O��A�&�'�mS%'́F���-�ui�����'b����-)䠞^���Ƈ 9%�Z�$,�ڪYc!NK!a�|�%����I�xWt�q�0�\1s��RE"�?�x��A�O��x�1`�Y-.u��-!}rC���?w�i ��'�O6�)ȳ?�%�3B�8v�{��w\��'��'��y�N�������)-�Șbo���0<as�	�c7f��� �O@@��H�0qЌ!9�4�?����?1�D�/ZV����?���?ab���!"��%Cj�%Aj5�9��?�Ƀ]Y���T[���	�U05ŠR"
�qO�8�'�}��e�.��#s��-��i��$�-���L>��'�/�T�6᜕r� ���f�<�e'��_�(81��)L`�U�,�x~��&�S�OM�m�0(:/����!L(^��I���,��}��'�R�'�r}��	។���[�X�#��s B�8��7:��`���$R�<��'3� �
E<_��Xʷ�N�T~�7�E�t��/��|7<X�'��!�1HÀBU~��B㙹?�<y2'P�?��;7�'i��'b�Ot@�vϟq��8㞓(��D1b�'�ў���`	!q{t��w�D�G��uXE'y��M���i�剴x�A�4�?	���(Ӂ
T�\�H�2����3�����?	baJ��?�������Y��?aJ>	���rY�J�
q72ݓ!�ZG8�x�$�1���%qr�� oK��)���,T�����-)ҕ|J�3҈�6��*{�xi ���y�̙K��p[���&�p�z���xb�s��\��恣L���(�/ ��X�d5��nZٟ��i��ihd�L�t'b�2�5��M���qÌ���OR]��d�O�c��g~�D��6�,C��¬_||ZQ�\��	n�v"<�"�m� a��9At>�PAo�L�d
r�b����::��2%4Z����꒴�!�\%ntD�H3�	)�@�i�(j�ax҅8ғsS�x�N�%���]�}�� '�i�r�'e�
�94�y� �'G�'���� 2٫�B8J��HQ�ڼn�v=��^`�	�Z����0 3�3���DL(��woy��q���e��a$�<�F�u�q��'C�q�Lv���C�!T>��w�'���':�B�������O�`�� A+���`��r���E ����xr��#t|4���6Z=,ay��ڒ���N�����<�q��;+0,�O�&V`05�r�<1�֙s�Lu26hݚM�:tR��D�<&LD�N����a�-J抔A�<���x7"(��x����q"O��j���O���`'�]5Z}֘[�"O��$ᎎ,�&�jtW�wq�l�"O�ѥ,���h5b�!T�%bbY��"O�1r�n:Gn�$� �N�E\<�Z�"O�aK��9j�X��B��,E�&�Q�"Ob	FnT�M�a�7�/t�4!�"O*�����A�$��n�1|��J�"O�0j��F<]QZ���M>�p��"O@�y%��4.$�)U)t�*�"O�qBf
E�^4WfM�p��u"O��+���O����接Q�HY �"O��Kw-@nBu����0W��x��"O�4r	��qԁ3���\���a�"OTЁ�5���J���nE�"O~56��.g�mb�O5��e�"OV-S���~L�� ��_�1` "O�|��'��M�Rx�6.6DKИ��"O¥*��~e�(�^7v��"O�M��@�F��x��߶cʬC�"OJt $f�������l��I�"O��bB��;�z ���C�L�r�1"O~�?]J�D*�>F�X��v"O����Ä}��h[��5��=�$"O���hU1k:�=cf.W�Xļ���"OHX�v'��Uz���F]Ѿ�("O��J���a[��A��x�"O�5����8��D��A½1�xyq"OD��0�} j!�-q+��{u"O(�#��9��4SA/M�N°;�"O.թĤڧ0	��1b	�Zd�xp"Oܔ1�k��c9�����J�.�Ш�"Op��u��O$���h�!�:T��"O���P��R-��h �˼o�y�a"O� it�B�Dz�l���E�A%)Pb"OdA���
)y�J2`Aѱ"O�4�毙7F�>�x��J�	�|"O�Yg��U:(��b'�7Y�6���"O���1�W�CV[�	�ʁ�`"O,� ������E�s�����S"O�Q
i����!K��;��AP3"O�P2���;�� �_�m[.P�Q"Op<d��Q�b+��JK�:D"O ��1	Ât|A�F�>H�}�C"O4��L� ^��]�g�)��F"O�����]�9�tX+'ˌfd���"O��rG�ԛt��Ak��H�]�<1�"O�9�$�+��H�g)��'Gh1�"O�(�d�͏{���?G�xIAA"O�5Q�mϤA�Nl�Dn�0 �ā�"O����y���i��O� $r�"O�I �	�{.��i�J�6�2��"Oܠk'C���
��0�Q�"O�0�� �/1�*�/� u��"O½��� ;�H�(ߚ|����d"O�-#g	�=�Px�� .O�`�"O� Ĭ�qIJ�r)�u��0`~��"OD��g�~V��E�]�M�
��"OP����(�Z%U8V�]�"O��;�l�"f����70���&"O�@�s�V�K������Y�C�"O���V�X�\�jCI� �&PC1"Of,yb˧ ��;#���H���r�"O���ߟ|�n1�Q���$δx��O����@�~L�{��B4~&��g�Ãw���5픒�p>�gNֶWB���ش^yƼ� ^�dHZ�D��3�^(��	�ri�f�[�p嫳�ڦWH��Dy��	�bI����"\�P�Ju��]vi;� �3g�jB��Z�έYT�:k�=I�E�2yF�<���ݘA�L��N>E����J=���ĿUvR��`��z����-�\2��Q�0�h���+�9L�\��`���1��ٰ=�գ˘R��y"o�؅Q7X8�!��I?P�p�0�Vͦ��7J�`xƤ4�J�^�lM )2D��"'�&G���p�[<OR= נ,�tڄb�'��H�&�ʄ��j
>)HD�(�T���'	h�zm��J�Mp��g�����$O��g��Z�` K���:O�|a�L>	���'y��ZEF�(�6�{�J?]֌�"�}�G�#(��#b9I��]�0���5u���a� �`C�Y[�/�'k��$�h� [�;lO(�1q��n�D���\��yBU��;SW���CD��|0��4(��>��.��8�m�8j��#@�a�Y�D�\�]��B�<;"MR��ܕ^F��)�+�fȳ'j�%_�\[�m�=�Ve�>�l�y�՟ �QH��	��ѪVF�d���@��'�xti������9��)B�R��� �^� &�����Ę��&�#0�D9M�H%��!�T�4��<�6)i��!�ŝ5���d��.$q�Ȁ�G��W0h�@��YH�j�v"Ot�3D��'��*5h�6a��ˠM�,����X�&�cfH�R>�aQ��"['�XY���L��8��"O��@LG�Cp��#o�=O6�%�r�Q��dTx�Yuz��`KL��p<�!�Ծ��0��(�Z1D4�EJ��p@�*��b	T.Y$�\袡�]:4(��
�G��:"ϥn����^-#DH��،{Pb����O�G91Or�� �N�C1��rƌ� * �̺����	�{F�1T�Y2+⤡:��y2��
d��#���8��5mV�n�Z� 6��3{r���S-]�v��� x"��7(Sr�:PgN�<_N��S(9D��m�B�ذY2.��J1ID#=[b�h�l��	s��&AM�TD���ރrm����ʋ !�!+�H��/gaz��D�Հ5$Gڵww�i�H��q�T�S�
���S��"	�І�H	mť3a����<�D�<���8�dp1��AQV]8>�ӭY�����ʬU������F� B䉎u�Q��9zEsH��Ja
�*ԏ ?Ԑ͓�A Tꐮ!�g~r�|\QjX:�\���e��y������s"%���@�	�C�+%`���	c�"��������I
>�Vб���8l p)R�� 2wQH����,�p(P��7�H��b��z-�LY\U&q`���9�&x��
O�i�D�w�,��'`����Qa�x�Gв{���˧ʐbm����懅v|q��A9�I(F������RxQ"O3P��0��l��
/C4u��$@C�̡
�ۖ =��2LC�Iͱ���'8��A�Y�*�(H��Q8Ri|��'��ZbK�P���b�O�Z+�hA�O�e6���of�u��J��V���� ;+�8���@ py>��[w6�x�`�C���toD/���2��*�Vё��R�j#p@q��EҨ5!Tc%���Ƙ�tiİ�3��`��X�փ5}RoF�i@�س ��|�1�&�8�M�;d��x�Vӟ�H��ȓ���Zf�}�X��"OJ]0�E�1T0Ƞ�:O����ĥA�ZuG�,
_Ȩm9�F������T?��#he�bT�J7&,j噒�X�2a#1�"D������U�@
L�N�t�$m���$CK��д�`T���@�$Z�}"��'��ɪ	�
�L��D`���f�&���DEpP�R7N�CNVLz$�ħE5I���!3�4�W��&o�D��l|�i���~�&:�ba�Y8	��'*	#SHS�&�%�<!W@C�f$#3`�'I��z�H�;�RP���(W��Md̞�78�h�t#�-�!�� B���J�x�J�R���oR�5�*T_L��s��~���)�-^�/-x��'P�x�w�l\hbH�����ڄ���4b���'&k���J��	�0}���f���J�:gğM��-���y�@�P�������=��s���S$�ؑ(Y�u1 ��C�"�&�t3$��u�D\�cѲ��"�8��my�d�`�@�u�Z�jG��T"�ӒOMJn�%��Ոvl����|�؈����jR�p�� K�@�Rn�my��Ճr�,ʓ(�X�h�.e�,�h�
���:*��9�bC_�U���������=�O|��o�)C�ȑ�g��9�ra�҈�|?C�C�6-$�8Ɋk�9��D�P���'�y'��
�b:�*eS�N���4d"�'��TȢ�ZyBESVҘ3v��/q�J	R`-7W�A��!�+GG,�E��p}� Jo��89d͇2%(������$њZ�2��([/-���DͲrP�'�� 9����%e�%XW�L�p"D�!M-�	�<��	#U
+x pH���6Y^41�Ǎ��`�Ҥ���DK�l��MC�'`<�) 얙a}b�y�KH!\����ӺBBn��/�#6�5��}B�A���
e`(o�
i��>]X�9E�B�6���Z�&� ��i���#�I�k�:)p#i� ���*RB)�ɡ�� b���.I�'����Ѭ�0p�4wi��Q�:�(�쒦X�X��@�fX�t�Ul�1�"2K�,a.�q�l���G+F�ƊU"�a^��d�I�Y��	�M�B���ʣ>sh�
��H�*���a���1���W��q��Ȇ�9���%��ᦧ�-��'�D�~���{�#�ɡW1�őf���-�O�f�x�A,Y��Xs7��"!Z�ekb�9O*L�QM��%�F�)��ʈ�� ��Ҥ[UtZVcT����FxR�qu��C4O���OI�?3B��"�0�ͪ��=4�(VO@,U�U���]Ϥ�.�&=Ex�Ŵ��I�MΠX��DZ`�&<RGP�`u��/��q��R�W~xԆ�ɘH��q+`���0:�j�,D�8`���ݖ6�x��$�$��Ͷvhx�� �T�JB5�V{�qO���0A�7f�
��F2>Ǝ�6S��{@">[I�9�nȬe,.M���=ʓ/�����T*7����LI2#�`��ff��H�pG�_�^A����i�& z����"�d�c��H�8)�Bc�7Xꨅ�	�fa�ӆ2�z�b�ש)�H��	#	�(����Ӗ}*<�&���,����
��<y`!\:1�X���5Lx�}ضG8��庣m�-A�"\Y��Ϥ�����0&�=-�l���F�&��{�t����@NRŒ&G�ShFXB�>�!E�*w&Ѝ�0��.0|���aPJ��]\�0�0L:������ȶ�ʜ��!B0����͗_Ķ��Q��n�qF{��!,w6��mG�~����9Q��vo�Xv5��'Cb�IC�v�jH��Q��
�3,F�tD��c���ՙ��/*|���Al:����.�O�q`v��<HL�j�ꂄx�<�S�LP("��Js�'��P��F!�]�#�-y+ڼ����
\Ql���U�r2C�g�'�:8[�#�� �^�ⴢKn��ϾC���	fI�-���b�D�
v#�V�0���8UlF��s���}A,H�?Q���"ʘ��h˾E��к��<)����[	��Y�"���">ѧlr��c�SHbmJ#Ć�>�mS�\!:��/Ɔt��{R��`�l�c���{���dd����E|D��1�qO�U�9�5Pa�C��).��ń�Ɋ$�°�7���1�i�Ed�hn�r�R���	b��Eit��t�D�F��G�9UV�`�i' X���Q�%�<��M��C�4ф�Ti�+���+��a��
ܠi�ȓ;_���b�9>H�x�i��F�3�'������Dh��b������'�!@J�*)�8]f�Т�p�'Q침4d�v@��Ao�p4��'EB�H0/�?h.l�4�V�%渰�'Bڭ[en�:�(i�d�ʸ k��	�'�� �ҎM?Z|\  !���b��2�'��\Ƥ��IJ:���E�.K'�$k	�'�8�Jv��G�$��A�;E��;�'����#�ū&�8}�2敽:�K
�'����C�55x-qՄ�)��|{	�'�D9 �bɨX �X�v���'��u�̀Xs��Stk�O�	0�'����6��k9T��A�����'ݠx��O	�h�CH�%�B\�	�'�"�	��̄$��Sƥ�>K�P��'{.<I���k6|���A$B����'��� Eܠ���"ŧ�c�H��'L�4�e������.[�#�Z��� ��Xd�Foc��!�H r=s�"O�G#*�Ta�@M(� �"O�*w�S�gsL,��'
�+��隶"O�\�&m۰lN5KC�X��,K"O�+�� ���Dg��>�$ ��"Ohx8ᗔ�XT0�$��o2�<��"O���d�B �R�s=Tyr�"Ols+ں}�`y�Q�Э
P�3�"O��h��!�`y��	8��3R"O����U�,��� H�fbw"O���^���C�ӟg�F]31"O��@�1L�hC�_�xċT"OL%�⦑�u>0Q�
�}t.�ڶ"O��d`O7A�d j�݄C���"O4�
�N�X~AEZ"*\,��"O~m�`�M:�M��AA"fD�B"O��avC�7%�$�C��ZD���"O,p���.����L�<5.�8d"OHq#tn	�M*�֫�y\L"O*E�s�=yP �� �)}k��""O*�#U,ǻ3��RR�M�]U�<�"O�Qy'���"62M���{��s"O�����m`t��GI2 J9�R"O0y���^A6��	�F�2"OF��7M�%0^&�1�IܳI���:�"O�xKg�V�������<�"O"�!3(�=�(E#vjP	r�L�#"O�z�$�0F�XpC�? �DĈ�"OF, V��R�h�BR�+���[�"O�ɧ�،JǦm`f�S?RQtq�A"Op5sR.��w�v-ʡ�E!`�Z�+�"Oި���� �
�*���@o���1"O�Y��:k�UC@�ș6��|�"O�ȋ%�V;T|���ҏ��}��"O
16K	�n�$�	��F��|q��"O��1�h�5:M�q���D�pS"O<���,�\�'�S*Uvh�(�"O��6J��N�����DB�o��Q1"O�U�dӽ�\u���;V8�j�"OZ��� 6@��td�")�@P"O��+v�T�)��4@�(�+e���4"O��!���Q�U�Nq��ġB"O�� ��]d�����N�"OT� /ذFuLU�#�(��M�"O�p�χ�4���#'�)��"O,�a���_>:��`��q$
�@�"O<<3EdC���A"&kC:��{$"O*A�3&��~aBܺ�l��u&�8Bu"O��(@��E���[W�_&P}���"OP5!�Sw8by2W�өq�t��"ObQ!�D��4x��k���4oX�4�"O9�f�ߑk�H���ѝ%n$$k!"Oܺ�k��
���5�	�Ab�>�y�,ʨ-�L����&Z� ڥ�U��y"��. �n�
pf؁�\��ĤD��y�J� �Fu{g"_�Z�У���y2�5�t×Ɇ�f��@C��F�<	0�?r�B�y��D,p�a�cZH�<��4Q�Z���dC�����$
�D�<1���B |Q�L�bŘ�����<1�lV_J �5�_0&����B}�<Qr�:a�x�ڵ`�?'�����f|�<���	1N�X��3"�P��@��DTR�<A�M�=X�l�ڐn�����PO�<� 652�#�KS�!c��-_BB��q"O�����7^�©��E�+).$yq"O�;6��"	v�j��Z+y�P9T"O���+"(K�	B�%V��Y�"O��S�6y*>���n�q�§"OHezp�%hu�����X��"Odŀ�D�	��A�ϭ"�b �"O4���$���+`ȑ��	fX��r%P!A2���P�ə#j,C%�%�Q���37�I�J@�uQ<	��45����R�<\j�FH�Y��h���p|��}�ʐKA�]�7�XS 
��m��	�ȓ� @��aW]NLPT�	1FJم�����U_B֞M���+xh��NĦ���O�8*!�0f�J�Pꬕ�ȓ&h���RbB()�)B��K��
Q��QtuSqMY7	;�J����j��ȓ��鸖Ɖ�T�n��h	�I�z����4�3��L���KqiT-���
�&,Ct�&p$Ջdɒ�eHZ��ȓ6`�)���1S�ԑK���zM���ȓx ��q��@�����Y�X��2u$с᧕=����g�Q�i�ȓY��I:��ޝJ&\ +яOj�(�ȓ7�tuIRJسr��A	ЏĬ~C&UF}�S�,�X9�"�B�(d���^�G��B�	�a��U���͉TUJ�#�'}��B�fw�,��mU�/P�aJ]�NX�C�ɶDop�B��ɝu�S�B�)n����0?a%LS�Jz�=6)Φf���3�$�W�<��$v���d��?I��;� P�<����Ih��%���Rd��*N�<A%�G�>tz��'���akUP�<v�iaUgLog���,ׇw���F�����`��u�f�1�&��ȓ�ޅ�T�	'dp�aA<V=�����P�XCg�?R�(��>=^I�ȓKn�1�J�D�޼�CZ�Hz�`�ȓB~dQ�Zhi�Nݦ� �(A Xa�<q�k�p��H�*/�գ�K� !�DӲ8>*IcթDN)��^�!�+%x&�QŌ�,�a�D��?O%!��W[�ȳ��ۦD]^Њ�)"!�DI�(WT��%jڗ�H�� oم!�d˘z%$���͟5��3@0!�� ��*%�.ck4��d	�;�!�$�7Hb�
�/�9hX�4ӆ�
u[!��H��P#"�;h\��MZ��!��5$j��PB��Q�|�u�ǭ�!���'������2L�D�V�T�6�!�A��i�!KhC��O�C@!��r}���'<(=���H�!�$
s�zL�1��+��MK)"R!򄇾6��� �j��I���
!�$��j���� *Y�
H�!�f�D!��ٶ��-���]� s�Eo�!�Dϴd���o�&x,����@�!��޽������O6C� �D��!�D��^!*ID���\I����+[!�Đ.= h�V.$}0�k��اDI�|����́4��2�eX-v=*�!/v�!�A�)9ja3�%��b*|Ui�j�"Omўl@��ӱD~<iS����)�1T�Ӿ_�B䉚n�R�5�K	���Q�[9�8 �i�R̓������� vZRO+H�``�( �xLPV"Ov%)�O�/jqi��(z.���D:lO �±���2���.&@S1"O�-ˣ��&=Kf�[$F_�9��	��"O�U�rL�^Z1IU+�婓"O�р5I�r d���L�Tj}( "OFL�E�4hR`[sB��_�@Y)5"O�HQ��&c -��]�Vщ�"O�x #A>H?���G�7��Q��"Oĕ3���i�Jg1Q��Y�F"O���@M7L�4�T&� �a�e"OP`�1)@+6��Xrϑ$p&���"O�h��Gץ�4�8ucX�m�@"OU���^�Kx*d�#š#��`�G"ON�٣���zr(�x�H��Y�:�B"O����LA��p�h�+}�\�A"O,��RCrpG'_5�{"OL(�#I)Ք0��A���,��"Oh|���;W� Z����tԪ��"OL�@B`V�j�������Ԣ�T"O�	�Y/D�����F��fP��"OĤ{�rd�k!�J�_
���"O`9(�������_v4087"O��v&�{al���.Rsj�8�"OPt)	��h��d��
G�;h�`��"O�ɉ'*�%�,����rI֕�&"O|���4��[1M6�s"Oz����m.B�) 7 ���"O,������t�*䱀ʵu�<�[#"O��� +#]��U1��=]��2D"O�6�(�h���,� �D�!�"Oe����%���+Ca�7�$ W"O�\i�� #�8�� �#Y�f�"O$!�S/�%�b��Ԓ"����"O���J-��dZ��Պ �,�@�"O�a����q�	�� �y�l�!�"O��¡ +����7B_�uVr�� "O��P�t |L���.5@�U"O �DGN�� �3dg�Z2Ĝa"O�S�A_-j�
�c�,
� �G"O+nS�ИĩT�F5x���C 	!�3v��T��n�+	�:ңJ�0�!�$Ýl=���a�Z�
Q�ƹJ�[�'l����X1,*�$�R
`�^S�'6��V@�Hu<�����]@�:�'&���GT�*Uȝ�@7]Nl��'�@���)L��)��[�)��	�'�XUZrf�3a��s�-�$��h	�'�B�����3�p�R������'3�=��M�#$i�M����p����'���P͐�v�\j�H/y���'LV50!�N�Eq��[�Aro�H��'����0�
!��!��f�贃�'_H|��*#�S���5�pA�
�'�4ȱwʌ�/�LD�s�ǈ'~"�		�'�Z�J�@Q�5� 5�#�P1����'7 ��@fB2x38�/��i2�'��k�9_�Ҵ��쒿	&���'�j  ���	̽ʐ��
>��'_��i�i˂s1�PQ�f��@���'�������^�Rƭ�t�B���'!�(�Ӓ>l����Lol�e;�'�N����G�@3xa��B�������'��j�k�>r*�h��ċ��;��� ��钆O��b!A����A;�"O>Y�-Ȑ,ps�؞vM�"O��1�\�T�v��T���2��P��"O���u�%NU�Q���+*$Ta�"O&�IegI�*��%�B�a�b"ON�z��KW@$!�r�ZH����"Or�� )� ^]A�oR��9�#"O���(>)��![���fP���"OTys��ꍫ���1��*�"O�x3+�9g��J���8r��t"OP�9":� S���H�X�X`"O1R0�S�:&��!�Ûv�MPq"Op"��
�>�`x����G$1�c"O����J�?Dx,�R���7�d�	�"Orx`2d>T�DH���Y�0Ѭl��"OH4��ǤdnD�h��_%$��U�"O�(��J��*�^�#w+92@���"O8<p�H�671؎O�䑠 )D��r�s<��YT�#qk��B�c2D�P	��Px�<�Ԡ$ol�0�3D�4�����!;�*׷Z�Bd��(3D�0�K�%5��ْ��U�K�"D��L<D�8 ���K+"�z4�S%r�"���;D��1��H!!�B����ay@&9D�<h�&
�dm1s)�Dԡ�%D�����+>�9�BKP�~��h��!D� ��+���#Aͅr`�TZ�=D��(���:m�iǂ� �\#��<D��r�G����Ւ�mհpЉ�Pd%D�p�N�В�#E�4z�����c$D��(�'ō+��XB��EVri5�#D� 
T$�"o�H����&lq��,D�$�Ά8%����g��d��P�*D�XJ�ߘB��WAX�gj��@��#D�<q��
�G�P2B.l0��$D��&��{����!6hX�[��#D�8��GJ�,�ZT�p�I/'�N��� D�D ��(�N�:��M�.@0��<D���ŀ�$iDz��5�ɷ;�L�ā:D�px��Ӿ5�����H�uY�	p��2D�\C��� '��Ir"eJ�c��M��&D�ā����T�YV�I%���S��"D����+��Q� 
�[�����c=D�\�1���:�P�WG&��Ч<D��Y�4~8x� �ԈMz����:D�pZ@�H�b�E#d+��[X�[1�7D�t0aCݻ7�f���#L:3 � 5D�X�0��7��贀H1/F� �1D������Jc���©?Rs><��1D����$�l��d�� Pl$D��S�Cv_��j�.���te7D���ĩ�$���\�Z��� :D��ddC�2�Jth����,�%�e&6D���`aУF�f�Z�HM�8��s7D�@;c�ܪQ��Z¥G-���Fo2D����FŎaP��A�凓.[�@�p�%D���lH)��3�
�N�d�`�>D��2�#>S2��zD`�v�3��=D��� �5�F�Y�]�+����/!D�k`k��{��)ʇG^%[y0p��!D���#�Y���̈'>^��ؤH2D�Р�W;��H�͝�x���V&D�T:�����Woۯq�aqQ�"D�	f�B�;QT�$�"2��]2�-D�� ��;r��T*):KԲ|G2���"O�=�
u����D�2cK�"O����1��9�b�2<؝ʒ"O�-�� A:zH9k�g.X��#�"O��B��I�Ggۈ}�$�"OjK�%8q��	4"|ŒG"OF�;4��z}���U�yG�|:"O>��U#��	p%"S���E?b�i�"Oؑ�`�_ ���2O�8��'"ON8��LƢ�~�)�C�<D�(2Q"O�L��X��@��^1`9��"O�J��L�.�ɦ�ӐT1F��b"O��c4T�*s�=zϴ��"OА1q�U%I�X��F�lǈ��$"OH ��O8u�v�A�	R�ybf��d"Ox�zNX'o��x�eH�<BW���"Ol���	M3O�8$� �	|p܊w"O�$����	Q���rɕ�w$��"Ot���"K�\�ȕHU��N	��"O�-�&�([��9�g�j����"O���3�L	��lPv��B��#�"O�@ U��L�8 ��!Ўd�s"Ol@��S���3d��� Ԡ�"O����BG�M�~����>�^mz"O(��0�S�VR���"�?j$�Kd"O~�vk� "���"Ej1�g"O�l��ˈ>�@$С�0`�2u�p"O@�Br�ӄ
b�B��#{ð�[`"O��"C�P�
��`�T�I�� *�"O� jF�#Ez��W�����"Oȥ�䋋A����&O�|��e"Ohlr�������Qd�f�Th�"O,����S��<�4#����x�"Ob�� ��d�h�@�</��p"O,��s&��n��]��-f��X;B"O�tb ǎ�Q�b�@�%��6��%�A"O�Xk��1g�
ݸrE��b�´"O�
a)�1%(%�25�x@�@"O�Ee��o��iHd�"���"OXa:r�ҩV��d�Ҁ�ct\	ys"O�С�>uR�i��n��mz��"O�V]O(ԔÀ�C5y$l�&D�S�<!�聥lШ��Ò15��(��D�<y�l�l�(Ȱd��428��hOZ�<)�J��1�\l÷�����{�a�L�<I���!��x�0�)�Li[#E�A�<�5��J�.�� 퀱+ڵ�4�{�<9�(+�����kO�w����� �x�<���F�Ƹ�d��=U���5��r�<��N4��N>����jn�<1����H}��-�;;��<pҡ�k�<AS�N!bB4Id��C�ٗ�]B�<�3I�����XqFJ��,�*#.�h�<�VCZ�Cj��CD�aF��r��y�<Yow��X��[�	��,��l�v�<᧩
�}yLu['�	.	6����|�<����h��e��~���#��P�<�������+ŕ@�&���d�<Q妆s0�Z�d�m2����^�<Q���|�Ĩ�L��������Y�<AfǰbK �0�ꞌ4Ȁ���|�<iD*Ġ�����B3Ed���t�<��`B�dF��(�͉�QN"�Ue�h�<�
�o��1s��(dHt!����d�<� ���)ǡ*��r�)��zC ��r"O�	〤�3\�>xX�I)S�4�Z�"O2��1��"q+��7�� ��A��"O �۰$GȦ�X��ԘYn�,!�"OZzG�Ѩ'� �j���;��]��"Ob���A���\g��mhr�P"Obrj��\��2���qU�tk"O�Ҥ֯��x(�̓�r:�Y��"O(U�ǅK��"X&g��>z�9v"O�hbSH��v�Ȁ*q'­m����'�!�D�s6�Q�4�dr�L�����' 0Q��g�2���!#Lm�Z(R�'�6q`�@-,(pb��3PE���'�}����K��%@EDݮԀ��
�'���;0O?A����w���A\Dtp�"O���6 ���@�k��#yD�$k#"Oܓ����O��X�g�Y��h;��9LO��@U G�|�b�z�%̪q�d��"OT�C6rp<f�'*xY�"O���&��w��ʧC�
 ��D"O��+�@�7S�������/�J� !"O��b��A��|��(�:�L��"Oұ�p���N��Y�FgF�n�6Ez�"O2�����/f҅��暓�f��"OV=�u�2/vN�Z�կ+��}��"O��83A�/�R�*`$?�U�F"O�6�؞*�$��-=t,S�M;D�`�d'�w��S��(9�}x"%4D�  ���lx1R�X�蘲��1D���v��W|rm*E�8Tv" 	�!0��\����O��̀&+TX|�#��,D�����S��HY�fBF�?�rAS&�*D����%�/[������$`�b9�(D���1����Z���!�gk*�#�f$D�h�բ��<�T��.|���#�!D��ۢ���)A���AG��)@s�!D��è��q�l%+����(�@��ɰ<)L>y���O^��ŧ�8`:,T{�b���@&"O 	Ig�֣O��b�A� �b���"O�h:��d��[�@ \���9�"O~X�� ���8�Oޜs�#B"O�����<<�TM r��L���V�'��	8G2�ˡ�҉h����avaC�Ʉ)�
k�g(m�͡B"�;O���d���W�<		& 0N�X9��<6v���9��b7��f�f����ǲF4X�%D��Aڇ;���ǩD�@��&G0D��@�$�.�h����F�#ZJ��Ĭ,D�̨V���PV��bECİ���()D�	!m^�Y+�ㅇH x"+D���@.ԃ@�⨈ ��zu6eh�#�	��$@��>X:�3�_��I@P�#D�P�f�ߢ�֍r��N�V�܁ڳI#D��IuM�#k����6��l�C@7D��sPiT�gZ� ��W#7mH�k!�'D��A��w�(��s��|N|��#D�3�/Yq)�us����ȷ% D�\��	�������{>�|��I�<���S�#�����ω0m5TX�'Ɉ�I R��0?	��L�i��=h2��/�� CISD�<)�o���L��<�ǩ�y�<)��ىErV�a�a=c&�{��Mn�<�+�/V�8+w��5�~A��&�ux�����<9��S|��8�Q�\�(���)z�<� ��a-P%���S��ݰ$��e���'�ў"~�6�OM"�9z�J3�Iµ��䓩0>!d�ğL����cӐRJ� ��D�K�<���M�v2l�ʍ7fܬ�11,�A�<Y���9ޤD��,A�z?�x��@�E�<�u�I�mp�&LѶ i*ZD�<��1,TCs�L�'c��o�Jx�T�?��(���B�#�EA�> >���?��'�^ IW��#l੷C��8��O>�m�A�c��j�.ܪe�>4>�i���P%B��R�ktlȅ�C ���@5�RP�~њ� � �|�ȓ|��!�ӭOc���f��s�A��z<�Q��4nC�%Iw�	jJ��]̓E<��fF�_��eC�
_�4��IW<pȆ�#Δ,r�0 Ȍ�j�uyR�'oQ���W�U��m"�:27����'��@Cσw��@��)X� !��'�@,ӄ�		�|�W�%_�:ph�'ϰ��g�X�D�&�N?fX*�S�'�@@�i͢g'T�3&LM�bo�q����ʌ^�N���y[�����1t��F�����N�g��A�#Sgf}	��:D����L����hB�Ž'�B!�)9D���w��Zhp�r�(��_eR��9D�0p�`I�)��y���'�@�Hp�7<On"<!b�ܼX�\p�)��X��yJc�o�<)�ƃS��ÆÈ�orV$R��j�<Yf���9b|��#Kܕ#��F~�<�gl�C��r��$;�Wv�<�@F׮*��@�F���:d,�F�Wi�<�� d$hd��P�ȳèg�<�u.�"�pbk
�00�Aq�mPWx�<DxbA\ qt��W���LL��H/�yBf^�K�6py��9��������y��B&6,��!�/ް,��¹�yRIǇ]h2t��
J8"�H��3���y"c�f0�4
�%}���,ޞ�y�-R�Tst倣Q�:���y�^g664��H�h� �*��_���<����S�0���c��SUpӲ�W5�!�dեNA0-�%'�I+~,ig�Ǖh�!��V�(���b_���(�ӎ<���)�M\���^1��U:bM]�<;<���'1f0HeBG
!�<��$ 
#L���'���RQ��,ɨ`Hc��!m�4�h�'���S�G�%딱��
�-�`��D�<���
Q1�U�u��+������y��
Y:$Ѻq

����D��yR �2-
��W��&���n����0>��NA|~�#�d��ƕRO �5�!���?���ꕈ�۰������s�!��t��"�L�(��qp��K�Pm!�$�k̴�J�H�I�8t����$?R�)�'f��赨��{�ap,G=Q�QJ��x�Ξ�r�`u��#T=�l����Ʈ�y��9wh�IP��ہoZT������yr�σ0��b'`K�j'�� V��y"MG�:� (���%\����	���y"�� A������iJ�"��'�y��	`V��E�P *������hO����I���ʳ�R> ��({4bAS`!����ف�	�	��ܢc�
�9P!�đ�C۾�R�W�}��h�/ ;R!�� �q@�$((A(��!�� p�"O�UY��G�>�����D�s�@a�"Oډé�^:���.�t��@"O�1�&+l��)ѫ�9W�ȉ��d(�S�I���K�O�2!H'E6!!���x)���M�<,ˑ#<]�џ��?��O�&�I7BB�0
 
�$�<����'R��ń7d՞�y2%J�I�i��'���iLф �DEBB�>U;<DH�'��p�$i�9�.ыA��*L5���'�b��e�S�X�����y�@��L>AK>y���5J�LĴ"N�� g�ȗ�� ��Wf�<	�Y)�>�z7a˷K�*�c�Vx���'��塑LFVl�7��*\�2���'d�ʐ�K�p��w��"b� �'y���P&M�8򥡗���J��	�'^i�sٙ;k������D��	�'����`ΘZ���������	ϓ���yBA�G�5)�I�{)\Xx�d���?�I>	.O?E8DG�>D;��³�C:(6��ō~x���';ƍ!6EŰN�F��vdȡK�)p��7�@��Z%l��H0vLՐS�`��"O�i��Ο�_�N��U��BO��>�!��B�Ƭ˔�=�6l�D��>�!���Kɸ�a�X!%��JVC�/c9!�[�=ݒ(K���]����@b�b�ly��'7�	s�O�J���f�WD9�#��,� �S�'��U�e�ݪ:��\;�g�3_� � J>����?1��䙟p��r�Yqƀ�U��H!/�<A��?)H>E��J�y�(�j�1R 5��ˏ��y��հY��	� HHxtx�B�f]��y��*]֒���n�¹�B�@���>��O^�k�`yH,a6
N�Q]�S�|��'*��'��OF�S�p~h�1/�z�2��5���B��!Wl���s��2Z�{�.��<�ޢ=�
Óo�<B��X�"ip�ذb�dj�'}�I^�)ʧ[7�]!RDN?POh E�?nw"e�ȓy�����eZ�N�T�em�	�Շ�M �ԁ��б?�����utXd�ȓ|$����!��i��I��E{��'����8&����� � ��ܠ�'Z޽I�q��݈S߱�N��"�'2ݺTGQ0#�I�jܖ?_4d�O>�����OO�dom�6���'�#�~a��'�$T�J�5��b�`�^
�!�'k5h��]�E[�`2��
�d�`�'I�����M�& ��R�­��-�
�'A��q�NN%��Pլ��6�u�
�'�J�N��&��� �S�:@
���d��
��e����	��Mc�iK]!���2Z`�,�ED"F�!0�AX!�ߧ}����ԏЈfK\�f�ܴ%�!�Ė�G�i��d0eY���㗳\�!�d�'1����$�
 CT���kM�$�!�$DK��X� C�SP&��Q�[��!�$A��d�����{>�X� 聂0��'0�OD��,�
��XpI�
{,��r/K* �B�I;7��0��ۦ<�8`�f�N��C�I#;�BQi�'S��q  ϯE��C�I�,��X`���43���R��Y����)?�  �o`:�@�F�a�81��3�0=��T�r�(���/C�E��12� a�<����Nq ���i�2��T(RDy2Q��%��M̧w6N	S�S'~ �U�H�0h��S�? �E�7	HA�-	��N�uI>}�%"ON����p���*婓O6�9� "O�a�l�i�}"���Y��*��'�� �	��g5ΠJ�`Ϲ�@�#�=����0�ብt�����Ѡ7��$�A��$3��C��&Zт޹d����㚌0�ZC䉩o�.�z�fP�U��h�`�9~BC�I�*��Q�*� �z(�`n	A�^C�?+�Q���`�>d[�ጫ��B��DԾ�����9q��5����N�B�I�}|%�f� }t�{�H��:B�	����e��uZ���a��,N8B�'""�t01"Ŝ�����M<R`�C��#k���!�Q��u��e�!�[�kn����$��?��<�R��){�!�D�h��Q�&ȢwDx[�F�A�!�dҙCSD ;��ٹq�i�%��4��}R�'��Dp�R٩�ʇDU���%� ~���7(|ʰ�Ġҿz���c�+��s�C�	's��<�$K�q�|#Į:�PC�I&6'*�K�	2'�ȳ����%2PC�	,,�̑���|6��A�A�W
^C�I�O��A��
��#��-ê_�o��C䉳L`��i#�H	r����IûeCd��$����yD�`��e[?C�V=�vi5D�&H�$�XX�O�C�:�Ç)4D��ŁG.y5�ʆ�\�P�*��5�0D�  ��?F]���G��L}Ԍ�Vl�OC�I��.����CrUr��J���B�I�^�Ѳ��I�<�R�,L�c8�C�I(�6d�@m��+$tY�go��v��=Y�'8Qx�YEI\!iC�lR4eHdP
�ȓB�
,y2�D5(����DS�H��8���CɘSRj�iB��;`L)��_N�����PD!������4���wE�h�����FY
q�O��R1�ȓR�H���2
���SM��l��ȓ��+.�&��PHƊGgsZI��\�0�.�� � ��E�=a��ȓ:�n��c��H�)�pBʻc���ȓ ����ȉ�娷H�7R�Dمȓ���kCl�Za�cb�w�(��ȓ2\ã��� ��|�́�8���ȓ �r��NP5{�����z���ȓ}�B�V�ރZ��)z�\�3*:Ʉ�7r֌���KG���k�3<�4`�ȓ ��ؔ�XR��T���/-H��3�E@���5ת�kT�P-&:��ȓ��A�U/.*On����H�-�P�%�܇�	�Zl�� �`ЭD��		GM S��B�	�	7�т��u����7���Q��C�*2}�%Q����"u����=g&dC�	:z�$��AB<H\"}c�k�
>��C��!]�<E�#��j�Ds��:5�C䉓E��۲�̰d�� z���x���,�	�rH�N�^x�x�����(Ld���O����]h4A0*F�I>�{���+Z�!�d�OX�%Z�fQ��6��Q��{�!�$�<G��e�>N���J��H�O�!�r�|�(��=\�5:P
�3��Oƣ=������@> �@,�6�E�_Xɡ��	s�,k�,E�.'��Aa&F'[_�M`3J;|Otb�ؠ�EF)��0ؑ�Kc}��#D�����G�S�y�!��+���� D�� (��Aⅵ7% e:���!gL8�"OȈ��ρ!6l���S�lk�y��"O�q0CL�S������56��lS�"O�h#p�A6}x�):U`�
���S"O�9�1߀aLڕ�n	�B�W*�{"�d��kWZ0"���*&Fȁ�䈔I;!򄎯�"P�ܬV+�����!��߁n����1��ї"8v�!�D͉|�l�$&O����0��$\�!�q���th͈(ᦌ�vc�1A�O>����RK�!�C���v��!����yr��8M�nx
��̩Ey���p���yBEd�(�2���-�e��-�ymP���0�G��<hY�v,�%�yO$-sn!Y�c�69�^}&��yRaQC������2�������y�a؛s��3tJ tCU�FJ�y"�Vt�Dp9FE�#p�j�f�ڇ�y������<)EJxp��TD��y�B.{�����Ԩt���"�:�y�)&1]"@��Z�qD���y����B��ƃt� �*�oP��y91��e�!-y�$i�/���=1�yª� ,�	$��r�������/�y��644��{ԉ֗@6>���"K��yB̆�_3qX��P j@6ՙMG#�y�'ڕiK�!3�a��Z���������y")P�tr$e�EJ-U���'J�yҧ��B��[�K@)N���)��yb�<[�� ��$E�]�z �����yR
<K��H���)S�L,1���y2�F�/�l\Bto]�G��DϚ"�y�ҿ>��\2&iA�Ia����!��<ю�DP5��u��x��� 2K!�D�^^M�u.ѫFv�؅�/!�ĉ�>>扈�@0!]N��6!�$ڹ.�T�b񯀀^P>֣͊��!�K�k(���ʩk�
I3�L�;�!�Dُ/XTP���B�����÷yp!���5d���Ѝܷ-ބxQHK!��?t:��f���k�rc�瀒p$!�䕵E�.��$�\����%�I��!�DL�*���v��w{���D��H!��Α2zx:�nՇWVP�33�!�dƼ8r�����x�6M)7��	l�!�D�[Q��3@�Q YJ�`BX�s�!�d94���,�t!�8Q���E�ў�F{�<O��p.��R&)���d>�P�"Ot-�u� 9(�q�;��$"Ov�9� St����F�ǈ�l� �"O\��"瘽N�"� ��ʟE7�#'"O����IݓN����+?�T�$"OZ@ e��6
ޘ�a�͜#+�� "O$��$�:7�d⑨��@=�P�CX�DD{ʟ��w��ӥ)C�z���qRK֟�F�ȓDE4`��9?y쥹iH��Z%�I"����?�9�%K�k!�܅��0L�����QX0I�r�v�r���	x�'h|�J.�@H�a5�4���'�p@�o	Dr���JG�B����'��A�-үDL�9�i�3D�0
ߓ��'�δ�ՎW���� �A�)�����'Hp�H9r�>��")�-�P�!�'���vjۂu�z�����&�Pa���� ���O	
��EzB靆6-z�1A"O���� T�O@Q��b\$D�*U"OP��7�++�����f$V�(�"O�U���A*j���g�Nf��G*O��;�Yz�r�*� )|��j�'s��.
�X�,H$>����'+䨻��&YҔ(V�ݗ*P���
�'� ���Q�Pm�(����Q�<�r�Ɲ1���&�$UfȰ�c�L�<Y�F�����cW�X:��� ��I�<���Z�#CjٴT<�2rcm�<q�	�@6zLq횰 �����A�oy��)�'0�X;�f��8�����-Xr�݆ȓp�ݳ�I�!;�����M%�~���޸�1tn����E�!�6p�ȓ6)x6��7����JW  ��=���eYW+ڨP �� Q4�Ņȓ���vBԽ7�}�bv����"O�� �.Dд��;/g��"O�% uL*J愴�7�P�zh��"O�x�Ŏڨ;���:4KJ�gr��Q"Ou;Vk�ajh�����`uB\��"Op��Ql�0g]|�;�k���"O��ՂAb}Yh���_d8Ds�"O@3V���]L�`�p 3#]܀"O��8�@�%"��Zrn�S��X�"O2��e�Q�~M�E3 -�UKԉ�"O��1)<F���l2_J�	�"O�Ah#��8��h�W��8��\b�"OL�;��\�(Kס�I�z ��"O^!h��۹I1�!����>�T �w"O�q#DEJ�ꑒ��ůV�@D�W"OPAQF��?��q���s�yۅ"Ou����$hd�ذVDL0X��( "O���f��b�%s�f�1"O��ATH9�X�(�� v����"O�8a���<{�d�hg�$0@��"O�]	c�N'.�P�,�F����"O���"ǳWb�XG��`�pz4"O�Vo��:p~a�5J�/!|�dE"O���,Y�mO����qp�"O|��4$@2y,XrF-U@u�a31"O��a$�!e	�6�
��)A�"O�P�(�wJ�h��B�|܈yx�"O��Q�I�$b�+�NI&D8Rp��"O��0b��%���#a�Q�t-J�x"O*tp�i���ul�;v�a"O|���vubR�Y��j�J4"O"YHt�K,D���I�g7��L�'"O�i��I���4cC�$��h�5"O �I��eH��ѥƒ$�����"O�DSE�!�41ҕ6�H "O��R���N*)��D��
 �x! "O|d��BJ5�|ݼOS��D`%D�<B�8���"��	/.��Y�yRD\.K7B��n�;��\��Dק�y�"֖'W�T��G),Q(Z�'X��y����a�O*+p�Q�!\��y�ĳ\B�j�,P�*
�x�L�7�y�D%�=�I>(C<��#��y�P�
�z7fA	"yb�(#���y�䑊O��|Yf�גOT�MC�yr�-�
H�u*��B�V쌌�y����d���Zd�Ń=h6�"�J]��y
� �h9�.�EcΘ�Q��7 B,��"O�d�₁�6���w�<),����"O���^�K����N��R�"OZ5�!T���ToѓU
�i��"O`�X�I߼=��!e�Ԗg����T"OFh���84�f.kr�1*T"On�r"+�Pbf�Co���"OH���E>h���IՌ�meb�
�"O���-Ԟ]�,��jL"6cb%��"OJ��udˉ*EL�*C ;�PxA"O`�T�O�j�̵'�Թڒ��"O�E8��!xUD��f��d�"O�ܩ�l�M���ɱ&�R�1"O��E��*9{�T�R��3P�^yQv"OF�����/`��kS�B�ְ�z�"O�]SU�	�1�����8Ӻ�b"O���Tf� s+"��e>�F���"O��y���7y��Pi�&�_N��)�"OyC-�l$����R?
7��ȷ"O��jG�ұQ�1B��N�yz|#"O����Ɏ�I�Z�c�(��D DjF"O�i�c��,i��i�I;	��Q�F"O.Q��
��_�`	G�Y�N�vS�"O(jJ��`Pl�0`=��ie"Ol���.I�qp-��+ݗCF��ar"O��@�A_��]j�,�OFp,�f"O,h���#la���@�C<O�舑"Ox�S�*o!~�[�%��L��q�g��5LO��E(�C��Y8УΔ:�J)(Q"Oh�K@�<7�Ei�b	'� I6"O�Mf��z1�0hP�E�ep�"O6���^#`�I�%l&��b"O<�����0��l�g�U.t(�"O�8JR�LC����W�Zc!��T�%\�J� [
�ԙ��f�3J�'�ў�>�T��9Z�
@�M�Al�j`�#D�����4]�����Ik�h�"D���bX'g\]C&	�)����k=D��0b��RXh���.Bސ5*0;D�8�Ѭ���HzA��h|�N%D�X(A 	�JAg!�&5XaI�G6D���d�R/� 4h�OV�o>���1D���@�'MY6A�j���iÌ0D����oԢ�k#]�C:QR�B:D��1���ٛQ��[�0�)�>D��[��ƌ?���Q4�W�Y���k6D�J���% ZAq���2u�]
��&D����΃N2�
�3����K0D�LIц�(-�4���MѶRBd3D��j���^R��X��&܌��P�%D�t�Ȃ�NQ��:���NXd�W%D���v&���|A�#��#Щ�`!D���R�ЭJ��E� +�8r�KY9�!��nDBt*@�P�HT��o5�!�$	�O�~<��*�;�Rȑ��)�!��#q��K9m��Ts��î~�!���Fn�Ku��{�uzܕX�!��Y�j��;dC�y�)R ���!�D.Nv�6���
�����	!�Dáy��2��/3(4�y0*E"b!�$< �@�b�T?+s�h �"t�!�҇z`t�gkK�D��T��e�2�!�DI'��d�� ;I�����J<4!�d&?��!���F�^1`�*Y?'�O�=��� Rx���[�zNh� D�y�z��V"O $�u�,n1k��F�O�V,��"O�\�qQ7C�(ed�#q�X@	E"O��A��_�rb,�cO�lm�"O��B���}��V��6uK�	b�"O��KQJ��<���t��=.@��"O�$����7l�)��� ��b"O8<���\��ܳ��OE_���'"O�r�Ҥ[�Fis�n(��1��"O�$1�HX
�pR.ߩ�$��"O@ː(].z?�*1�C	�\Q��"O>�A�i���H���.f��T�"O(�	��;	���4I�p�S"O� ��2Le찂ơծ?�L�#�"O| Ѳ��H��,R�/K;m���"O,I����R=�ᩄ��fɨ�aG"O.)��혎#׾�����82"O^��B��а2�A+�d�A"OZQ�C^j�\�k�A�'}�.�R�"OF�Yj�}�������$2"OT�y����J���j^�`�`��'"OVd�*]�2 4�HqIS��y���~az�rU��6���#"��yR�6�,1`S�/k�A %!ߺ�y��Z��E)�� �>�9J��[��y�B�sN�0B��<sj��F�F�y�	�)D�`a�a�7�  Hs��y��I"_,Y����,��X�`N��y���j,����p|n|�"���y�m�|�"��@�V�}��PR��yCѬ9Y�hqPjP�'��e�I2�y"� �<Tظ�.�9'2xxZV��y⃞�e���it �|��:��ԭ�yRa_� ͼ�Jk�:��I`ïҖ�y"�% ZD��92�8��QAO<�yR� C���)�����`��n��y��g�ᠵ�����Gm]5�y2J�ki X�'�[uH�&�ې�y��ɏ���!]*i�!rv"���yB���1:UӒ@A+@X��ըY*�y��V�	j
Y����B��:�y�F��xgBvmC�l���CI��y¡�52y1DՙbH���yB�� Vu��`�� 㮆�y�; �`�Z��B���o�+�y� R��ҽ�T�6u�u�&�yr�G u.x��a�A���*�A���y��ޛpg��aI�;��p�(T��y2+�&G}"ܰ��Si�Pđ�H��y�!<�����@+vahE�ʕ�y�,>.0���	�b���r�ҩ�y�B������*���#-�vY��s���J2g�#
6��%�����ȓp�<�`�A�p !z�N�'w�؈��Έ([3���{+��q�'E"W��ȓ�4�� 54�
��	<�D�ȓ%�T���V^�2�	1f��Dju�ȓ�=�"�k�؀�2��
~wإ����PS��J��5IR��#$Z��ȓV�6<�΀�[تĨC�Ҥ��-/Jx�h�('/,����ȔR7r��6�����'�&4����'i����O�"��'fǡ'p@�"��튴�ȓx����d�(:/f�kgcOc�`9��S�? �@j� �21������I
A�yR�"O�DBF+��u�\�!e��:��C"Oz X����,�5n�#0>��"OV�A�L���Y�w#+[-�iz�"O�`ID�H5��"��,5J%�"On(�� 
9�� �q��v NM�1"O^������>�C^�ka�#�"O�<��@U�X� F�8M���"O~HɅ"B�<P�cl��:��e&"Or$c���<���GlU�^��I�"O�ͺ
]+4e�7�� \�<�"O<�����<�^�4�:���"O���!h^&zX�0�g�	r�1�*OH냯v$Y�`�:~
��	�'2��ۧ�ۗ+b����Y&�]B	�'���! �6�H=C@�;}'}
�';j��q�V)GΞE�Dj'ƥ��'*b�
W�I�rqb���3a;>T��'h�<r�'�~@�6C�.���
�'k��)Wǔ?X:p�Ջͮ%��Q�'j��cP�+m��Ȥ!�d�3�'����K�Qg��t.ڂ�9�'�̤�䊇�D��ND�?�S	�'��Ę�&nR���	v�z�	�'�����敐Ij�P��^Ă�h�'$t0�b`��[RH�Y�����'��	Ѣ�U; "|�����.N�.l��'�xa�B�<Bd�c�>P�z�'��L��m�(e�t��>8�ҙx�'0>�yV�	�.p�Q"+ �4@(
�'�-{��̠L����.�A�2Ui�'B���f
M?L�ZY��e_�@c,���'��C� 	��w%����'��T!�	Ơk�֐1T�D�,7�)��'c�q�����ܑ���N
��Ԁ�'snȳ�#�5�<��&\ ��'��IAg͒i^��Ѥ`��|T��'됹AS�O�T�64�#M�{?F�3�'�xbB����0qJA�{<(e�'CN���i����HI�.!)z�K�'9��+T���t�yD�[�'ڠ�
�'}8�e���Gp���E�5v��0��'������)��<y����V��'�d�R�	�e�Z\� 
�H���')R��o�/ah���á�*�6P��'�`[b�\WH�`��e�5z<�H�'��sC��?��x3A�x���'a����H���Ps�9q�( y�'�^�Y� E�.��u����j��5��'�(iJӄ�-[}�d��䍶m��!�'&� ��i¤@Fʈ�f�Z�7�
4��'�r�9�Zg
p�v�_~�x٘�'��"d�0SbL���B�����'���sg�^.Cs�uYǜ5�t���'�B�b��Q9<Y���u�ʔ��'v>p�a���%2��	S��w��Q)�'�`R���J����q��n�n9	�'v��aV�N2��� 2>� �

�'��+�N�R�!����4��
�'��ܰ&��c�pС�L�� �I	�'E$a�e�6r\�\ ��U��@��'�~���&�,�����?P�}��'[����H�<4�:�RҡVeV�'���k�	�x�D8KK%i�\`	��� �����>���mT4}͢5x""On၇�C�s~9�m�X)�3"O*=Å�K�c��9
q�\�=<����"O�AAX�/�^Ё���
!!N���"OZ�2��](y�d+ѧU�.&� u"O�𐔀Ψg�~�������g"O@���~|�!Ņ��s�v� s"O x# � 3X��Q�䗸'�����"O�e���u`��'�6�[S"O��Y��d.�����4p�Д"O�����c:&���|X�[�yR�8 ���F0_�(����yR�B-r2p:T)W'-b�`����y�َ/!�`٠i�$\&b7�y�HdtA��U2D`��� ���y숈Bt�����)��i�"�K:�yr�lᖠC�F#L�*��X�)_D�i
�'�
`����1i��A2R��58�"
�'Ղ�c��a�4`�Z�}T2�H�'�J� Vj�>s�,��F�L���'�F9QiƆr|1"AB��H�X`��'�F��G�-Q���{��Һ
�|8��'��;�H��*�(�c(L�z�'"@}��G̾�����[W=4�+	�'�~�pV�~��)��Σ�\���'@��jF�ha�#�Ȝckz���'�4CǢF�kX��Mf	����'F%KC�(y������d���'��9�(�?X��s�#��f����'���b$&�Z�,�����M��xR�'7*���S*e���+At���
�'��qۀ�5!��5�V�9��Q�'c��YO"G�T)З�*bz�t@�'/Ʊ�4iJ�Q8��ᙡK����'�p1�g)�B�nZ*X�N`0�'��0�CO�+���&�A���s�'pJ�1f�^�z�(Ј�bW��A�'�N��4ϔ�rf.��#�+n�i�'�Lш��h��m� m� Ug�s�'�ve ���E��ّ���J��LH�'p\�S@: ��X��?=�dm�
�'b�A�4I�'��(q�
ϯ-(�Q�
�'�=(@�zSڼKP���2x��Q�'i*�iqe�*v��kGIF�*CZ���'��8+g+ǂչ��Կk%��0	�'��%c�(8ud)�`h�9���'���v�A�,�V��i�ՠ�'؉q�$� ��RHсP�6���'Ԭ�a�-T���׈��@�'��!AO&s0�H鄏�FL�R
�'����7f�R�3! �p�n��	�'&0�����nb�����t�T`��'���{Ul�LP�������B�<ɒ��gG)(!���"P����Q|�<���ڣx�"�\��g	Q�<A��L-` �DK�\>G�8��o e�<��OG
c
�u�f̶=�бz�d�]�<9b�W�7).�	C���*\�<���$9�l�S�N�ݢq�!B�M�<٧���U4�k�퓶`a�,�J�K�<��'T����@`�.N�!dh�C�<��o��V[���[0k����g�Re�<�o_��%�G��/A�r�0�Wu�<)G@��B?�E��늷q�rH�j%D�� ��bp�&�4e�����`5�Ȉ�"Od,`��Y\>��EN�k��)�"Or\�뜠NB��B��ۆ2�|pe"OּQS��/($D`�dGĜt	�"OvD��Ñ��Ѭ	��A�u"Oµ�En�V|X8�h�hy!"OִKF��; ̠`���p 8��&"O�L �k�[ȴ)
�0�Tm��"OV�z��]�{4�LK�'8r�I�"OZԒ�a��3!�X��A� �
�[�"Or�{)W�C`fu���|�F�Q%"O���`G�W��p�%�&�0U�W"O�T"���94��i�0{�2��"O�IfV�oTXss��`|���"O̙�F� Rv`��Ao�3e�F�"O)WE�/_������O��u�"O2�ӳ ��,��ɠ�֝-�!�DA<���B���`�iRmŸ$�!��Z)[���J$`5I�.�a,'p�!���c(��� +��&�V��Ҫ̺c�!�d� �ni�bE��9�>(sB�s�!��ϱ}{��1֣�f�d�k��#5!�d)�d�s�(U0"��4b���%!��ר	�b
@%C7�i���T�"!�ʇ~�8�c#	��=�՛�� !�d\�e��3�9P�1@�+�,�!��4`bf��5T�@j%!��L)u䕌z,
��I!�d�'NK:�z�
��T��`�E[�I\!�d#}Z,�(��{�ĉR&��r�!�D�(w�AQ��͵,�F����<�!�$�\���-L	����G���!��U:p���T$)&U2}ag��a~!��9	����5Bd*��V��$=!��^"gA���
WpD�(m�!���=7̸ E��y�ȹk)u�!�D^(�����kB�bs��9��ҞU�!�d�L*8����"�Ae���@�!�d�r���p1�@&hd��-�!��!<��u;���N%�Phqv!��F�*��W�))����q!�;J�&�VJ�p<�&�K7K!�D/���x��W�T0�q%��y�!��Y@8C��Ԍ�x���K0=�!���Ԏ��aT>��m�p�τ{!��T��3w�H�6�2�8��G�k�!���5CG�T���9p�tUc�,��&�!�$�76!�*�9nm,Y����_|!��\t�X�z�%���,p;s̗��!��6`��rKmf����ULh!�� ���scD9��"X!�L�{��d�0�A�\]���f �&e>!�dƃZR��hF���(?�ia�$O5nD!�ć^q�X��jN$"����j�!�D�&�����/�%��9o!���{�y�1�vd88��X7�!�DX �P+t'ܦZv:����!���g7��3�Ϛ�
g�X��� (!�Y�^����cA���KH��O���d��֩��*&.y�B�F-!���^�XekM�$]/rD�&H4$ !���fl�H"�Ͳ�ra���I!�Dϑn ��%bW�z���m�$,!򤞑?���%�E�n�ᵬ��>1OH�=�|� P����КU޵Xg���!$�0xG�' �<�b�Bsh�>\e�:��N�vX� Gx�'$Ă��9?��p�׈|��X��'��X�a!K�6Z�tz�k̟v�h�'N��!� 0��a�o0h>L��c��=�#�(�*{�>MC���43��&!򄂐!���C��j�b�S!��h�!�d�1߈��aES�h1T��A�Py«R$>��-AF!�
��1��]��y�,^-��*����P>�yc1�y�(��{Ji���P����&C�'�y ��4��mܺ:�4�P�뛭�y�$ �y �O��h� q��FM��y2.�?X��,�3kN4cRV)��ĉ �yRk��A1N���M��W�� A����yB�TfM��� U(KqT;Wf����=?iӓD�th��� #��!ʡe�2a��gAq���bTL���m���=�ȓs�Р'����{ĥ8(e"��>�k���
5�-q�F�4��ȓ=�4����E�����A��?�R���@Ǻ�0�͂T4��t@@�L,L��u�(ѐ1�M�>!���T�_3e{$��Xr�8 .K'h���鏧g:i�ȓW����B3��|l-%P����P�\(�-Q�Nh�*�K�uV�	�'�ў�|���%VE�ꓟ>��7a~�<����{5�����QE���vNBp�<1ĿZ�Si
�}�D��cX�'{ў�'uj0�1�N�Gʄ��
�m�R��ȓ;pȸgY�bt0U�6���ʤ�ȓ=((��
B'o �br�t(T�'�a~Ӽd䂴�'�=\��t��'�yRh6/<�S�΅[ݠ@�0	3�y��P����� ކXa �z�H��hO���	��,�SFI���1�$�؀t>!�$��q;��s�F';�AR���*d&���)����c�A��MS�oEXT��PB$D�P�`�E)T4�TR.�=dw.�q��<�
�0-�h0'DK;Ml��bY�K�2qDx��*��p��ȱ���<z��ѵ6�B�ɖ Q$]�B-6���`gm�V����=질��D@�.�*P�d� �JL�i�w� m�!�@���X�EcH�{Hq��&���t~r�'�ax�(A7�M��LϷ
���d���~b�)�'"b1{ �%t'�t2�mN)7��I���?��$ jz���v-���`H*7*p~B�pӀ�`���'�;%(�#��u옅��� 
�0?�UU��{#��6�~l���0�`RW3D�\�H�{r�P�'Y6^��DpU`;��g~b�9	���k�f�.y%�8h5�h"��COZ}x�b0��=�A�<=*���v�O(�=E�4�E���2c`*ڥ���
�yr	�4��5f�� ��83�@V�9��<��ԟ �<a��%����j"1<�c�IZ�<!&���	��I�$�u��G�� �'�O��1,�;+͎�J��A0CR`�S�'��&�Ty�lφ::��!aLwL ��F6D���2�d��A�r-��i�b����>K>���OӠ��!G�j��3i�����`�'꺩ᓖ����ߓQ�>Q�O<��O�(H&�Fμ�4�U�N軣"O�e��*Ė�Z$�i��d^Y?٘'՞�=�}
�oǤf��WH5w�PʇPV�'��	ꟸ�π <��m��M	"�0v�J���
�4OVO��DD�-�2�y��["+�n��H�DD�D{J?��=P��^�1�dɯR��)LQ(<��4`�h�dКG���R`DB"�.����?Ѳ�צ'�ά���3Lk�A1Tw�'��w�OY�Չ�ǉ'�Xt�%N>�@D��'>���)�8F
|���-h���'��<
��ǉk�%��
�/y
�*�'Pў"~z�G�, ����=��8I'�F�'�?]p�Ҋu��B3,P9\r�cH�>�	�+^T�����^����W��XЄ�|�ΰЅ���7����υj�~Q��А�	��q��yѕ���E�����	�F�J*8lR(�0GH�[��܅ȓd���_�1 � �e�.C�@��O���(g��p�sMԯl�P�k	
!�D\ ��q��4t��Q �\!��g&�\��o$�`k� �2,!�$�9b�H����Q��a�XD!�dF�h����V+̶]|��7Iǔ�'Kў�>U�@^=:��۰k28mX�B%#D�;AƜ�h�Dص��I�YR��<�Im���s��/c��UJ���K`�8���,4��4�
�@���DnY�s�v�aFe����x2O�sڔ��Ds��`��%M��y����Ex���]�8b"���yB�kBt�{�.�d�����E����hOq� ����?R���H�*�/�d�"O�E	d�!~hb�@�
�5�&����IaX�,�`�" *�@��Mx�h�Hu�:D�И!��Lݮɉ�̡ �\��6!+D�d�U��.!�"Q�K%_��xa++D�裁�Z�w�Li����yR�$*D�`v_�+�P���ǅ^�zYc�%D�艳�)(�b�s$n�'j^�3��"D��I��D��r`"B��>}zU�!D��b`�j�@��i��B
��($�OV�T��xt+	����t��D�hd�ȓ6b���̧�����6,�v�E|��S2I~����
,>�PJ�B��B��=W�Έ@6�Z�b�)�$�n�B�	�I�����Z�?��|�"	�T*C��a+|;	ɼ����UMo��B�I�N ���R����ɪa쌗<5�b�dFr�O`qB�`�1gX5�6FϙNT��"O��G�Ƙ(���FO� �(!�2O�=E��J1Rt�����L.+��}�CH���y�GM�A�l��M�0�U�W-�!�y��M���Gn�W�p�����0=э��"|�<�Kr �U���U(ؒ�y��t�� m �_s�`��Y��<Q���D;=@��¤���e��	˞%e!�ła��3Cj(����Bg���K<����� �\ڬ��M�%p�fF�<x!��fpV���pY��p����!�ė�e@D�s$�(1pR��3!��t�azBY�l�'�R�hbNX<dgJ�ӑǹ	�F��O6qB�R�2Y�Ćg�xu
W�I}�O���LC:�X)�(�9�H%��'�;�,fB +$b�/�!�'d*}P���Q��!�B�-�r2�'@�)�X����sOʭ� �'8<u@��$;+��c��q���'��a��F�0K�ņ9cN�4���� @����^�c3�dadE� 	�	"O�L���@�� �[���:m��j�"O�"�鈽M"�J e�&��m��"O !C���S��� ��@C���"O���a�Ľr�����DR&Ow�z�"O�eA�	����ޫl ��p�"OԸ�ƠK�L���R�U��Y�T"O`H�SG 5��� Jϗ/�.y�"OHa���z�d�b�"̐A�8��"OL��
��!���P˄��"Ot �GgG�wt��1% �Y�R�	�"O����ԳPtf09��������"ON���#;Y
B嘂gÍs�İH"O�4�B��D89��FA�!��t@�"O4pt�B�^L�4(F�6�`ڦ"O�����Ҍ� Z!hT����"Op�A�jA92� �� n�1[�&��s"O�5��I�r���g
ASb@QA�"O��I*!DXů_�PIJt��"Onh
!��)�q�1o'���X"O�s��� w"�	7��"*��0�"O�@��a�
Gs�� DA*~&��"O2t�'!�M3"�[2�Q����"OX�`�ܩ����ŦA�����"O�Ԣ��0P��}RD�I).�P��7"O8,��g��32l��f$��`y"O����H&yg��ɱ%ˠwc�L�f"O.H��޶j:�a�D�YrfXۂ"O8
N+aY�\�A#��-Z�AQ"O�U���d;̸a�R/A�9�R"OZe�b�X��xXQ��M
�]1E"O����	�|a�s�Ӱ�ԉ� "O@� a��2(��acU���T��H��"O����(<�Y�%��9��x`�"O�����ޙSF��!�"Of`2�"��B�\8[OJ�Z��I�E"O�y�7/�2]�
ya����ye�`�"O�m��)��@���Ie�oR�I�3"O @R����`����d�Vܹ�"O�u#F��rS��d�i���"O`<���m�.yӒ@D�F�l���"O��ōX�b�NisnF���P��"O A�޷Oz�\*�'ے;N���"O���LD(��\Q�Y�.n�)T"O�%�vCr�+ʍ����p"O��`a��� K�OƬl�F�zV"O!B�)U�4��hڬX�zYr!"O`	(����_�rY*ƌ2Y��"O��Ä�Q�	����W�e��\x"O��q逜|�z�X�$�J�U*�"O�=*W����`b��!5h��"O΍����}��9���ƶX�j��"O�*`Q�Z�=���^y���"O�U�G��1R��%��n�]l�+%"O6!���%)S4�P��\|d9G"O�� G�҉?fb�`K����4��"O�"��l&���]�\�&�	�"O���[��.d�o0{B�R�"O���� *i
AB%L@��*%�"Oz٫�D��v
��,�1&�n���"O
��2鎢 ��h1��i�6�S"OXp�Q�Jr����cH��J�fT��"OP]*��ד7�.02T�À&�l�*1"O�n��#�~����P�$��`C�)�  $+ENI�2j\�B�W�Q}@}ˤ"O�!��_�+�p� e��ra"O�<�rh50�������%}	�	k "O���E	�
�ֵ;&c��x��A�[�.[�O��}�?�&�
!3֍6���!��W�<�]���\�u�Ϭ ª�aw��צ�C �I��}��G]k�e�!H��ԂB�&��=!t�Q�_W��v椁�W�;�2=���Z	VQ`��ȓ%�iP��Q+�Yv�[-Y���>�&+W*vDN�:r D%)v�rU�^�:e`�G�u�<���" �-��*+�ܩµ��D Z�8�{�'�g}�N_��V(M�����h�M1�yR��=�h�kuf@4Q ��ͱ�Mk�'�,v����$֎'o����=
��Li�⟒<
�{"��W/��eX>Tb�DǸQ^�A�	h��C�* �� �LƱRf�*T+ �V	�C�IC�bFț24z��q�_
i�C�ɢm��x�F�Y�^l8@�
�C�?b�|��'I��2.�� Ǧ�*s B�:d�\)d�F�j\	"���B�I6h�BJ,JT���4�?i�6C��!�xAå}�:AcAi�@C�I$Q��ڒ@�.�,���#­Wo�B�	�d���PCV�b>��b��2r�B�I !��Ɂ@Y-6�0$���=x�B��
z��p��K6@԰��I��B�	���s�LR�{��<��A�>W��B�	�V��U�r(º2O��e�Q�~e�B�Ɏ@�dX����FLaa��kL�B�<�yҤ �44lUDAM9C�4���Z h���'͂�����(ّ� (����'�p�Z��& �����MV�V��A��* �:�~�����;F�$�dǶC�R<X�I9��B�I	6����G��=����t�Q�!Ũ�P�?~qzاO�YE��O��c��CR��x�G�9Apda�"O�����*�mjt��kw^��ѳi�~�R�eU�I��Մ�ɘY=�0cbj�un=a�'V(`p����,$���j��N��?��$V-�,
"��*k���j6�SI�<�`�c\
D	VD��a,�]�M����*֕����)�Z� pIU�iw��{Ф���,ڂcݺ(\�����2D��Z�,L����İ2p�(k N��0&���Ιp��	��u�B�N���?)ՍE�ȴ-8���dԋ6I�ą�I7O�20!�b�'p��Ӑ=�~$sa��
J��T�f]���V�`$X����I���ZF�3e����S�O���t�)�I'qmijv�V3��	�O�2�cSȒ�'��$ @	��Őq�7T�p3@���yRn`��qw��͘1w���a��?��̙�q���� ��9Oĕ��c�E�t��RQl�C6�^6oh���F!!�O*,�vI��V��'���(�sÀ_�5G����}lD]��/R}~@�+�܌Fy��F�*9h���K]jLb�aC ���Oj��c�Z��a�f�0��j��Ʈ+m�$�Wh�!r9�ħ�4>�� ��+$��i`eRKsv:��[n����P�ӫQm��R3�Q���,�)�$;����4 ��M�x)ZV�`_ɫs#�'�y�

#הd�c�"S�t[B��?�~���9�$ 25�iA�)����S�G��-�v���x��ޮ��AC�ǒl/�X"�/�O�����G�eL�:�����$HW�^�4y��q�g�q��Q8��΀p�䭅��e��H����>V�s����<Ӻb��{�JO��!��S-y�⍘B��vnP���1|P��4�0$�d�ԯ��	�!��ċ�N�!�dA�qe `�4N���S���8��1w&A@�e����?��[1h�sb,X� �L��9Ow�]B�2c[�*i���\�y�A�<�4{�/�9kꎝ�#��<r����ͳe���f�X�8�2y��'m�1���4v����'BN)�U�7���+CJƈ2-"�
ד!�ܬ�A"l�H1"�ɩ(�2d����J?��IЏ>����>��N�{.����i4O�(���5̀%[td[�Eo�)�b���2� t)��'nL�y&�|Z�e�F������A�xMn��#J�[����G.(B�)� ��p!�n��C1a �Ƀk�qO�U�]w*�j�b�r)ɧ5v��,9ވ!��A��Qf(�Κ�yB��"H;hhZ$BL}�DSs���MK4��L�@�y�/�C�S�OZ��P"΀y����gÂ(
a8�'d:�RD�3Vt����k��p�'���r�e͓~���EC�=[���'1�h���;��`Pt4x`��
�' ���A2Ԍ���]+g̬1�'�DT��>"��rc��))�b�x�'��a�u �.���i")�� �B��'ѐ�c�̕�d�R�$��!�'ˆh�q���.XIH10�<a�'D��jP
sI�q�������'�NAjQ��W	�`� ۧc���
�'+�p��IO�;��d���È}�����o]? �T�E�Tė/cR�	�ȅ�7���w���y"B� ��pzV�Q�{(�,��N!�=Bl�'��#�Q>���8��j��ܻ�mT7G��$���$�A�(Q��z���_W�؂�.�2��2u�
�v���U��m8���ES�}����(̱I^�"�c/,O��ALa�0���4Ǻ|ҷ��*F���#�]�r}��� C�O�|��l?<uX')�9��� �K� I0<%�رA
�!gG�|@�-Ǧ�(�
������O��@S!+}uD��Qbį\���	�'Lf��r��4	:]Q��T���4�@d�.��U�`�R�\e �,�2��O�> H.O�D��H+4FT�=�`
O�D���c��Z �G�SJ�MY`�r��x��ج �n�	�$ڗs½��ɨ[�����ji�
c�LZ~!���DF�TvTK���!a���K�T�f�p�����!�*ׅ�ZU#5���tt��d�.�4�� �r�pl�hH�+��I��*���g�[P�ҁ�D�C��'��N�^i�=x���[TL	r�܄ZXC�	8:��Kr��7x�� `�Y!^d԰�@c>!n`�g���d���&,��b�	�'��$�����R $�vhչAo����'��4�wk�����WB:S�h�:S��K��d�`h�z)b�s�L�*0B̠�I
l�P�h�/��!����J�G���D��|LZ-�W��]J�G�E7O�x�I�]5F�icgY@3���5�a��:%
�� B�6z�M��ۈu!���'����/���Z�Q��#~NX��Opܧb�|#* (��D��U�c� Նȓ{I�h�#-�/�b1�eDJ6zZM�'�K�<�RE��O�#ZD��Qӧ�v̧��s_��v��8��%����BhH5�.����OQ|�|0f�ۛ��١!��R�ё�F1eᴩ�p�9LO��sa�%CTصX4�ݶ/�Hѐ�'�]A���rӮpHR��;�X+� U�@�����?���c�b�<A� |n��P�	C� p�G�Q�I��50�,O &�1�o�M�O۲�r,�5�R�����	7�
�	�'�Z1{��X�R3�����J�I� �EOm��]�l�Qg�'�� ��C4�x��'h���Xl��I���$j�	��ztӇ�ھ��q:�X���S$�J .����+��L@�ؘ�p%���0����:cA�H)�Q2+>i�w#�=2��G̠ �ԡ��-��ӺCF� ��hh�g�b�`���GYR�ؐ&�9v�p�ٵ�?D��Ad�O$0x���RhZ�Y|*���g��I���x�s��>�qO>�G�}�y�Ԁ��[��P��Δ7m	.	yЬ8�O�m�t P��q�m�T�P)����	S�������dR�B:"D�
�4�����/hF=i6�/9EB��	p��I�YH}�����arjG!H�X�O
25,��vN'v����S�(>T��FI^������K�&s4�&���~�ǋ_Z�4��`�K�4hߔ�h����^�Αsb�����C��c9��K�Ğ7�Yx�g�!F�, �'&��P� ?�,��O�$$���N}FE�zˊ,���ɦe՚P@ͦ��?�B�ł|#�@�҄� �@�5�V�p&�1�b�&*H���-;������O�y���:E]��n�B�բ*���b�0�t�p ��U���	�[ ��3N��:�ÆF�t�PH�� ��d=�� ��'q�dБg<2�0mz����E+O� �i��}tb�'8�pч&�H(��'>�a��VY�����M�Y�Jh� L6D����!|�&}�v���W&��0*�)�~i�'m \��AĆUG�Ogt���DF}
� �1n�*1�  �����R�'1���A�5P:Q.���0�P��ϑ}4�H3��CQ?9�)�y��1d:�G�>@�C��'W���J�<w�`��I{�4�J�`_]y�hچj�`!�ƇG��: ��/�s���7�n}�b"������U.gWD���fȡ��]̪�Q�>�b�ǸV��c>A���Ū�,�9FO��/��I�C7D��R�� Q�>�[bL�(P�Q���8D�HȀe�BB��BDe
�e��yY��7D��	@N[�SM��+`�H�fx�iy�)!D�h A@������6������<D�(�4Ί�\������_d`��W�=D�� ңЏ73Ry��\(
z�F�-D���G�PRf�=I���+�0�5D� P���R`��B	�z� 0�4�?D� XG"��;ֶH��H�/�4��a;D��aႅ�3Ăm��m˖6&�/<D��H�hC�t��L�,�`h@}��� D�L��ƫr�ts�B���VaB�>D�0ɶ�ެhDf�aP��������?D�L�Ō?�6Y1A�%��98b�<D�D�A�͜-{@���\�K��1h��8D�@�@�˗/~��W���~�H���3D���rY�K"�5�X�^/|��:D����l�$�|կ�"��%qr;D�t�V��e��rckV �${ի9D�dj�/����`"ֲLI8 �,+D������:��M	T���8����)D��R�À�J+�q9P�Z�$���*Ӯ%D�D؆���<�1�/r�+�O,D�`jQE�}�$�1J�":wt��F D��!C%�p �M���M܊����4D����/��\ʺ��� D����$D��K6�ӻ	���&E��@XE�%D����gQ�:�Ľ��U8.�h�ks'D�d3�^2�V��6蕞;6ٓt�+D�����*L;i��џbA�x�&D�(:j��rL�yt@N>~3���g+D�t0ց<�]���8~O��0-,D��T��<{��q���g@��0D��qE�;�Kҝ�HdYv�(!��;I6F�"��.I%F�z�
�]�!�2�ṗ .����4-0!�D�D'��`�`Y[�%!���K!򤚮r����#���5@lՒ&m�-)!���[��!a�
Ǳ,LrѰuc]�!�DE;�nL�cFN�H˪ೖ�H��!򤝡��� "�
.X��D�$�!�$��8�z��6\-p��QElV�!��?څ�G�*�`��Y�/�!���0�e�N�_,���	%�!򄙑Z�0Qp2�X4Q9��`�a��!�g��	��}/P��v�C?6k!�ą�,�&��ER(Jl9r���'
b!�]�N�B6jѨD~��ܛ�!�d��E�r 85	ˈ$�Xx�g�-P�!�DJ�fa��gчG�@0�f���!��S3DP� U�È����$��g3!��ΫcWJ����>�̀F��3�!�Dʳ������|)|<�R㞙�!�� !(E�%>�*�b?S�!��1��@p��#'�d��]�1�!�$:��0f�^�2��M8fnR�&!�B�_�0h�!�M4(�6���V�U!�Ę�bo�D�V�u��@�۫9[!�� ��ʢ�:0����~I��"O���C	6�Ȱu틱f�B0�q"O��*c��?~��Mճf��U"O��Q�Ѹ>t������B��	�"OTac�F,*�������7�m�"OVL�遪I�,��Ğ�0ʔɋ�"O��4(�@�����B� Q,�p"O��Wn��pd�A�bA�6Z۠"O�E�E��(��!C ��Y�Z�@"O�\�0�P�*�|D�$$E�^R��"ONɉ�h����D��x.�`�"O��kǈ`��!���PK�m03"Oр'�[���a�遮4���"OŃ�1b�� ��/��yht"O�1@2�E����ɀG�(x<��"Ol�Z�ႏSCP�0��ܛk���G"O�4BT�]3N��A���OH��"O���@�[�?��́�j̵	7`�
�"O�lH�^*u]h|jA�_�5�X�3"OR����U�J�L5��׍i����"OH��&RF�!0囼"�]�"O�4Y��
�0`�d��m�(d��"OP cGK�|Ւ!���[ݺk�"O�|Qp]3:;���7.���x�"O�8�o��Q-~��#�!���!"O:T��/K�a�b(��C�v� mb2"O ���L�h�����'�<��0"O@���J�7C�����Śf+�%@$"O,d�菢KBB 0� ��©�"O�d�¨Ɗc�іDL$=�pB�"O�5��#M���^�z�"Ov��,[sN�b� 1�8�"O؝�f
�-Ī`��AՖY���q�"O�Yx���,?�La�%oW� ���#R�'�v��\Q?)��̳2��NG�	���!H�<����=2jm1�J��0�څ^��^����sm!���ܨ��FJ�a,:%@!��g�d"�"O\u�d���m��k��Q��T��lՖYGx��<}g9�g}�#2��)��[;8�j�̅�y��� ymju�h��db5۰���M`oM�\���,|O�� �'߽"�8��䌕�7��82��'���B0F�B�r�ɡ~Z���)� �����\�d4BC�	0e^����76ͺ0���+	�x	C��ν��D�4T��b,���O���aN4@���R�U��	X�+�U�!��чM�)%ʶ~�|�S*�_rU��P!mX�d�/Oxݭ;M�=�֥*�I@��ui�D�JP��q���x����:z}J�O���y��^��n9��jM&A8��)���#�M���/\N��dH'|Oh��R��=Re�5t� �`	"1� ��R��q@ǫ^���DP� ��9��h��b D���y���(����)�z�<ɴ�� J�ʵ� �Pp�����I�f<��
�۟�%Q�I�N�����`��'�"e�?�0ڵ�X�k��f�*�z����'5�5H�ˍ%��!�A�ԁ6c�ԉT.�%J��v� �P���3J��$��	���	=Ut�4�Ԩak~8��C,k���>�q��&K�B�2��x3\銖+�=WDb0��H�9�M_JF<�HԸFB���R�lH�P����P�L��D�O��� a8��r�^%_�8av�	,P��}"�ڂ1�R1#��+2����M�j�<dn�k��D�RO�7bzP�l�&B�`�F�	�.���fF�?��x���]�A�M����c ��DJ��Ŋق3(�~�@̋fl �I�L'��d��h:�\���K���|���i�Y�K�m�����"�T!�G�����dB�!��>�p"�Tvh�kIJ$ � r`.��v���s��`	��AV�`��Kسo�B��8'�`QC�Ì/3�L����J�8���`l�ĢL�U��	�[��PC+�#��O�(j�	byHe��J�C�)�'r�R�$K8Pz�m�nRAJ�'[��h`@�k�(d��Jr�I�%�E��O� 6� ��xU�h0׼2��q��'�~}JQ��O�N�f�I:d5��*�kU��,��T\�(�Q.֋Y����E�'��[���i� 
5���H� ��DM� +OJ��A96���y�B'N�|�{ƷEX�/�G�Ҹ���pdp���İK��L؉
��F~�K�><#�M���	¯���bteP��L#�D
7�!���$�z`[P��s��y�*@?��	�B���c��6z�s������q��Xb�B�I�iq�u��c�H�����n`�C䉟+x�r�T������쐀IJ`C�I���͋P���~��� N�:bC��2\l�Ȥ�U
O�h4XÅ�p�C�Ɉ V��� �QZRjԠ �!�
��#sb'i
�:RꒋuQ!��h�HU����<gPx��I���!�[�q�(����7[֜��H��%�!�DR9Z��PI�2/1���槑�^�<�D�[�j��|+���f����čA�<A0&P����9^�\��� ��<�TJ�I���[0e�X| �x�<	�ĕ���br'C0��m�]�<��I7dðMz�����\jŋ�Y�<��	�$�d�d��e^�-�@��_̓e\�%�`�%O6h�b�U
�tQ�ߊJ�v��!�'c2 @�Z+�12��X%P%|�g#OV��O��1N������lP3 M�IT�I�pol�W�Ɵf��OW,�H��P�XAq�*.L䔳�'�8�ڇ�rѲ�ʐE�T�ШO:l��	�P]�<:O�"}Jp�Q��rg��
��aЉS~�<���%;mpm��C>��l�����{t	�f�ܷ��g���
�Oʘm�֭x�L�L(��	�'8!���P1g=S��\?�H�&ǟ��	9S�'�z �|�ݰtb�
a6>���Đ�+ Л�Ƥ��W&2��ǉ�$Fc�������I����4�� 7*�!�mM10]t��'����ᏻkm���O�>Q�Ň2.ʅ�4�φH)|qq�g+D�8Ƭ�Pv<\�e�J��\yaVd�S���9^�ʢHJ�3���-���裂;�LTJsh��%���$�/��u����(v�0�#fD=V�6N�	��B�ɴ&&N|(&�L1X�0���C2Sg�����1Pd��z�{��U�y�4b���Fl3�$�
�y�I��_9n�D�K�K�*��#A���y�%�,6�\����7����v�%�y�I�{�t�Cיm�m �B�y�D�!z�2t���]�(�jc���y2K��z{��'I��%{�]��I�>�y"N�a�P!��/I�䰺'd��yBl�E�<L�"LZ�}����ԛ�Px�� ",J�dnп���(�.;�����z<afl@;�=�r [���'�Qh��!7MIY��&�\ǎ��
'��
�jM��*�3�4D�lKV�ίe�\���ƚp	XhY��<�Rm�:l�=H�E)}��I Dl�+2K_����X�K�!�dS*pv��G!���"ӈ�>��O�u�cMĤ� ��qOd��v�	2ӐM��`��[�RA���'-n����Ӥ3���Z�"�"U���_?Z	&}j3�ly�#�l!�ቁ_�|��`�:P��J.�$��?�!�ہC�X��h�>9�ЎVqn�W(� 6�P�!��a�ACEgF���?��\f}bB򌌴gմ�v��qyR�	27ކe���XY?���-@O���֌:�i�i�n�フ8�|��n�<:�!�"@��̘e�$ݔ�C���3��!�)��F�*[���L~���(X��&^�`P�\.xX
�h��5?ɲ�����$Y�PP&�
0�zd�GO�,'Y���D'�a<���Ob-�&�'<{������D�5"tS}��4��;8uџ���юK�*��Op)� �]�NHZ�n��@�!5��1c-ߦ;쎼��� "<"�Y�F��&�>n�ʓg� 0AB����IEGpK��ɠԉOG�D�6'�6�v�B��o3�݋	�'�ʀS@��o�~@����5\P�����p��9���R��N�<���r]�d���M	2���dc��1mPq÷9�O�m�M2��p��^�� ```ս�60Ӱ��7�~2@@ ��	(���F�'��r�72�����Ak���huld����8�� 7R����g~�
1�O'qv՚�Z9^Z��D�AC��B���).*4CѤ�#��QX\x��)}bK����|��m]SX��a��Y>V��P��b�V�<����q�0ɀg茿h�����*V�<��4;x��'��50Y�����HS�<�,ρ�e��iK�*�Tm��cWv�<i� �.�@����ν1}�pQ�%
D�<����g���J"�^�,k��@G[�<�q��IN�D�4�9z���� �t�<qsK�a
 =�b��7_@ĐұGT�<InWe����&�Ĭ<��C �W�<�5S�tDf���D��r�i�M�<��cZ�o`
 ��C	�ki2%覫D�<"�ֆ�PZ�CشZ�X<x2c�L�<��ō6Y��k�v~�9�F̘K�<i��6��(X���\�9��LC�<I�M�NB�h��"G��(8���k�<!��[;O�>�Я+R�s'��N�<������iz���j�dx��"_H�<)��S,^�v�ZQ�$7j�`�@��K�<�6F-Eʆa��O�:ًQ�}�<Q�l��a�R��dK�.�L 8�
�<����3��آ��D�L(@�
|�<	���5``Z�/ y0�K��^B�<�(Os�Fm#�� QVT�����<fh�2%nJ`����-y2�ժ�q�<Y�G½)5��cF��Z���J�DZZ�<�g���D�PL�i)%���*��V�<A#�`�؜�"g^�A� X�!dY�<��I�P�^�b�j�=b�LҰ�[W�<ѲJ�r�uS��P9�̴��kZR�<ّ�؇mN2\+�Z�\�1;S��H�<9�l�#� B���b�4����LD�<�r���^�E�d
��L���Sn�<Yu��n�:�q��C� `tN�l�<���Rq@�{A��/;Әջフf�<A�
�'z-�0�Zy�Vd�O� !�d���X�/�j�c֧(]
!�1gT�
�LH,D�taP'�!�E#ޅ]�j���#_�Fl��c"O�Y�&ɮ�����O M\(��"OjY�)�jS�@xҋ�L�q:"O�(��V�"�؁��m*��jg�O�t�����1O�>�H �>k�X�С�q&D� �
t������ē��mJH�X�r\X�OD�+
���&�f�$�f#%§���șZ+���fӜE�����Õ\k���?��K-��tC+�;G Ś���"a;����D�0T�⟒��qk�
/-'\��⥊�+:@!��5O���b�,_��'��}Z���-+H\�Mݼ!$n�Ht+�7;�آ��5p���|�r��i@/s�U���+}2����G��7��:�Uy�N����}n:�Ĉ���Y�`��E�d�����ٵ�<�9q 4.@T��شX"�>�H �^�y���z�D�:s�=�V��֟����/gJV�[!���n��l�����@��� ��6�ȪX����ۋ����[�l�)�8�R0�`&f�F떃�*(\9�c
E�	�2dj�L4?y
ç*j,��_�-&9�&���rܠR���=��*Pᰙ��S���/��8�l��lLdPU�"����Wؚ̨4��D+z�}�z`��A��tm2���I�z펨Γ���C�C9�6ҧh�J� ���b�=XR�L���	:Rj�	࢈�.JՋ5%����%�'���_	�R] D��)QeHd�4�Y~����	5?�VI�3�0|:�L@�G��9�tL���R�f_G�<!�K�|��٘T� �R�0���A�B�<i����{�B2��p�dE�F�|�<�3/	3,������=. �J�-�x�<Ah��@	��J6xPM� v�<�&�F2���cg/7Հ���&	l�<y!�m���X(9+�� G�h�<Abg �ᚷ���ʀk���g�<)���<6�P��Kʬ��%�`�<�AK�:I)4�	$ņd�#�]�<Y��#D%�Zd��q�,����@�<��+��S}�%8F�C+A�脡C� X�<х�H�QeL0!C+U�ʘ���̞S�<�M�)z����K&è���Q�<������D�s�P%6��� �	h�<���)y�@�bSM��,NXhQ|�<A1�~�L��	[s"��#Ęs�<Y�)> ^d,�d��[*�D�VJD�<���a�
la�_�v&~Q���B�<���ڝ^�p��.�w��+���A�<ip�×4��M�`O�0jB�r#D�<�wD�NF��pHԓC��@�$�B�<��
�,'E��vK�U˨���g�<�E��#0��X��)�9a�p�C0!�a�<��ܰ���+sB3�,,�0nPZ�<���	1��ݐ���R�<�cC,�S�<�(�(+ �3�OՅBl{�M�<(Y�-�fd�1
:_�\+F��s�<�4�A�mP8 ��7c� L���D�<���9��]�3��+��lpG�C�<�r+��T���_�"T����i�<9�O��s��$��4{#���rj�<�����D.e���,1	�Sgd�<�����T���ÄM�R8n�*��Z�<1��M )�X��E�+�p`)LY�<���۱.c����bɅ���.S�<!sD��
(��ǥ�
�ܙ",V�<���ʲ�0}�'�;��A�#)j�<)��!Z�$h�R;8�P��CJ�<a� �@�8Yf��4[�:Ńɞz�<���0�`� �ַo�e���u�<!Q�^p��!QeB@�i\�u�lt�<i�O������ح+��b!��m�<�`�54�J���-i�����dA_�<�d�fyp��Vݸ��,�Y�<���s�������3������BQ�<Y���"�r�0�gX���i��Jt�<����6�pq��PJ���c��K�<��*S.'m�̛��#���M�<���Ь5|&���#�&"�z$Bï�E�<�3��	�dtZ�M�&E���i�-
�<AM�g?^��U<+���i#�}�<giH�7�$@�cB;0�]����N�<1!�N#7����9Xd�%@�<��'��[�^H;5NǊQ���+�~�<���>! ������'�R|��(
~�<�w�� u
ވ�m�"bR�
!�O�<��kY�s�Z�l=9�Թ#wFp�</�!��)�A(��Mg8�
�� G�<yS�Z�eت�H3cP�C���*�
�[�<qrg5M�\@0W 8��(��o�o�<�RI�*!^]�")ӧk:����Q�<� ��9�^��A#�IԌ2�켨v"O"���� e<��C�^�L��QA"O+k�?C�-�GgZq����*	H�<�0ȝ��bM��ܜJ�PH���i�<���8z�zH���� �<�i�GPO�<y��#�tűBm��]V|�Y5�L�<r`VO��h[ǧ>�$Ɂ�K�<��*̓͸�[fM�xK�-Ie�H�<��ò��}�֋���� vCM�<Q"��F�h�ɇ*�n�`�(�h�b�<�p,���JR+��=(6q�c��V�<�A�A�5``L!�@_�I�aВ%Sg�<5M%7��tJ"g�}�l0ëe�<�����4�&��'/�	c~��$]�<ї���Jg�]z���='2��fHp�<1r͇2'H���ŅJ��,��i�<��E��dh�b�Ql0���\�<ёC' ����1Ǐ�3�j��'�m�<�sfϮl�t5rdf��MZW��i�<���!h4�m�C��-�(US��Ic�<Y0ǅ�Rx*a��":-��$��)�y�<7���!��	���*α�whGr�<v�%&HM�wE�_��	ӅSo�<�)mzds¢�5e⢉�"�m�<	�%Q�<�BD�Z|\A�GH�g�<��.��D�.`86�M�A�\=0��`�<��C =l�p�͜@�Z�:��A\�<�BI�K�n�A����VeR#F]�<1'Y�/���P�_;)�rbtV�<�E튦[s
�'D �M��Q��w�<!��-Κ�H�E�5\6��%�k�<A6��	O�$� ��Z�2�>�h �f�<9�J&.��!��]I�\�h�'�Y�<a&��?e� ae�M��y�b�W�<I�m���^�b�\5z��e�e�J�<q��Y%�N��%�T�{���"��C�<񴮔R�Ȭ��L��	xxDq!O�x�<���O�[��8��S�G� �wo\�<9�c�C.L���&��R��H�gLW�<��S	Ҟ��SD���٪���Q�<��ś�G!�8�WE�l��7�XK�<9�d��/咴y0�&=8�1JS�F~�<	�喭j-R��f�
+�4�+x�<�5��|�F���#��U�n��CO�O�<��
C�. 
!��xH^D*�"Zu�<��I�j+��a�D� ��a��͝s�<Y%��?��[�B�)����ƄY�<��m��O�X��/G��,�Z�<F���c��w������GY�<�#��I� �&)�cн��YO�<q,�����`���W"�@�FJ�<A����|��E��<p�=�)UD�<�w�GY��a�
�-,�8x�#,C�<i�k��C�� �R-n��X��}�<��ύ�]�a1"�� �2���^�<�NE�J)v��$ŗo�>x@��CW�<I7��p.�,�#���-�dLHd.�Q�<Y�`@�d��L(��Ոz�VM�A��M�<�����H�8�򋇅W���:d�J~�<y��Ҭk��4�r�D�L�|���h�v�<YS�O��ls�J<q[� E��q�<�T���o�~tZ�̞9U��K��l�<�D�#5&����R� ���o�j�<i��ڈY��et$��@�p�C�[�<� @�CF�6�q�#	X�R��t[�"O@4�ekNW�|3ƈ��V�I"O��Sa�_����1G�;g v��"O��[wᛕ@�J�����aBXC�"O`����O�a�@̐F\�;2,$"O�uQVC�'r2��eb��;���u"O�����)�l`D�G�1B"OԑQ��!m
����ع?'�`Ya"Or|��� v�����8 Z�cE"O�q"�h�6u���4tt���"O�}�D�$��L��S��P�a�"O���N�?^�>�	ӂ,^�ɛ0"O���7 �u1�`�X�\Q"O�e���O�O�~K� 
1��#"O� 9��	�7�P
�A�!̨T�0"O`���ES
\Q��k����x��"O(��*U�tՙ*J�^�P"G"Oh�3 D
[Ҝ�SG#̾V%ޘ�"O��@Ƅό#���쉛ut5:"Oޕ��F	*;�0D٥A�g�B�b"OT��B�e8N�#bǷA�|�+ "O숀X/,�%0ԋ!j�pa "O ���-�.0yJ�qˆ�ad��b"O���!K�%vC�ԈK��B,��p"OUh�A�+f)N 8ƕ8���"O\���ج	
I�тP�6�$ ��"O��(C�W�i�L9�%1�Z	$"O��B�E�����S���"OPpR-�u�欂%iǭ2;& �d"O�̫��A�Z�i� �U#.���"OE��m	=g�^Q�@e�&Q�*���*O��RR)�6�a�f��F�ޘ��'W�h�PBT��L��\4*�`�'C��7��{@���#lM��*<)�'FJ�#�n�jx��!� �.S�'�ԬP�(T�=� �"'YU�	��'HZ9 � �+̨�!�	O!,j6ŀ�'�����U
�x��L9)v�h��'����B���W]�|�� ����'��D���$.���JFʌ
Q�]��'H�k�(�"5F�m�5�Av�����'�����3�q���2��@��'�h��#
T�J�K��pP����.e�<A�'Y�CmD����()�$-��x�<���ǬDI(�5��-;��@8F.�s�<1���d������* ���sQ��x�<��a�8v�*@C�$W^$	a��r�<4�Êc	���@j��)â�k�<��R�hIj���	�>$`���eEg�<�r���Z����$-���eA�f�<�oQ�<)z��1
{�ڑa�n�W�<!5H�y2HHY�ǌ�&�ܘ `a�Q�<)@�'}��X�X<p&�^i�<�` �x�͘�pkV x݌�yRg �R������Հ �j�s�y�`v�ޜ:�G�'�����y"Í0.iV��#lN��ᦇ��y�b�*77\$�a�3�t@�%L��yb$��h˰�r�e���#�Y�yrcN����QJ�	G�^�iu��ya��l���{��
lfLQ�F��y2�� v~P+�͊.j%ȴ;�f���y"�
�.�12UMH
d�Y�l��yE�P��2�'V��
����y
� 4��F��J}�F+�d�&A �"O�q�DM�m�i���@0^�F<�"O @+1&˰�oN^�E��"Ob`k�Pk\�����53��T��"O(�zU���H�9F�ڐ�����"Oz$���5d@3-I��n0r�"Ot�!F   �P   x	  1  �  I  y'  /  S5  �;  �A  6H  xN  �T  [  Ua  �g  �m  t  `z  C�   `� u�	����Zv)C�'ll\�0"Ez+⟈m�˸�ɼm��D�	G��ط/W�F\���g��݃DjȐ}� �ɵ��*Ɛ�)�ޠ>] %�;]'P�*��.a�)��� kB�kFJ�=^49#�d�`XT9��^5�L���=XX6F6@� %����(4-Ꟍ����,�k��4UCFl��nN�k��EK���E$�OH-����)\X��k��������Iٟ�I㟀�2l�T�De�1O܉|Lp��̟��T�Iw��?� L�8�?A��?)RA\d� �Z7��Y�]c����?�������O��� �������'�����Pu��F�=�]Rq�:���y��)�O��ɔze�ݳɔ>;��HY�A� 3j��yR��>>���`L<����'Y@��2���E���S0�˟�����	����I���M��2���`2��6��H�6F��}
��'s�6��۟�lZ�M+�9D��}�J�l��M���A$6��O�v�h�ħ^�e.t��O����:fy�lA#J�:v�H1g���ܺ%jK��4��-���hӜ�l��Mk���2�!�9cs�`�A.@��1%G<p���C�Z�?e#�V����<Tw�@qq�.�?���F�XB�ks�T��1 '�)�O>�:6�	v��p���Q n2�@6����h��M�'SE����h�3���*ӫv��Ԕ'kў"|�C*��!(��W�q�48��+�,�?ٌ�d?���sM���r8)��,a�D�[u*F�!��K� �q�@�&p���KB�p"!�2;�pm�!�'f��i���9!�ʆK|��zQN�X��ݲbJMc!��B�qr�a���P�|@��H�RI!��Ѕ4��2�?9h�S蒲ў�˃�2�!�l}��*��5�<T	����`���ȓ@L�q�Ne�4�/[Pd4�ȓQ2U�v"]%&���C&/�8�ȓHv0�#��؂`�t�����"WU�]��5F&�+��`T�B�|�X��ȓ6�┉�a�!K}~ ��ʧj�b���&�"<E�T��]�J@��	�Թ�eΑ�H�!�˸f^����N��l����b�!�P*	Ŏ@+���-&��՘aM�-m�!��_"-y����-n���Q��M 8�!��×Yk>�jsa9Q����Vi�d�!��b4�"��&�ԙiE��um�I�,e����QeL�i��!�v����bR!�d@e��� ���+��tS�[� 8!�䎂 �nt{R)�<��c�"!��+���z��]�~<�R狯i!�D!;�J��&A��x�i���#�y�M]
�~7+?��K""��٢�OTp��b�#��'r�'�r%��P����ҚY&i�/4<C�
e�y�l�	�r��0�-��9qx���	e���� � �89+�'

Mb�K��Ǖ>݆u�����O*0�1�'���sӢ�ď'}��ULV�7(���FA��c�˓�MCS��OhV%"�.\4��d�n| �t�D'u@�Y�@Mm��OH�=�'�RH͐G���As��GkX1��)���?i(O@0%J�Oj�ı<q��<��'�B�5L���r蹠�ъ1"Q�O�1���������@[��@�'Q��)`���,(�����0`��+qO>уƎ�Pz�hAh�$b����1?����	o�p̧*�n�Q�Fǯ�����Q���%�<�	S��0���9#7(jq�Z�^�~ba+�t�>�B�V�ɶ�a�iڞ}֮yB���Ҧ��Ivy��2p�T��$ ���*%"�W'�1����}��H���A��;@:@eP���]�����<+x@C��9^� ��GT�/<����èA�X@�F�L =i���q󩈼�Ʌ}&����lA�X�u ���XlZ���$�j���'f��'jܩ0����-���c��+s�Z=���'	�_���	c�g��C�%THa��k�6���fX�_�I�Mc��ilɧ���OR剎b�D<��G�>{�R=��l��Q j�kҊg����aP֑3FeP0AH4��w� �hb��:��J���A	v�y@ʚQ��K2,H/c�C�	C	zts��I㶸�&�+BP,�#q��O�H��ɿk�:�Ɣ��`l��̟ӲC�	�r��4 �n�qS���^�O��lZ]�I�d��I~R����|�,�'M��(�������<�'{��'��A�&2N��CᆯPQ{��ܺ|~� I�3��EU��j �k<�S+�(j��
CsȨ��;F��
ٟ	sڅS�͐K���!Ǥ�-��O(�i�'�қ�<B���>D;��ƒc�DIq�2�d�O���D�cά
���� ��q!�F!1����Or���-���lec0�{�i�T�'��� 4%*y��4��'��)�O�Q�a�?��4�U N�	4h#���O�$��hw<-P��"fK/��iz�	BH�'G��dBtG[�5����A^� >\��O$�r�I��Hn�8�e���v�"����5�
o�P�惊.U��R����v�^��y�I��|G���'����j%$�drQB�l����5"O挚��T4����-�4��� �h�ة�&�A�VV\8� �{��)b��}ӆ��<q����r��?�����dX�uXV�M�
&���'��a���A���R�|H8#ŀ�O ��xEC4�H�ɚ� I!��_:y����-ߋz�4�a�]	5�^���]�,��'��I�%�� �bS:N�� 0�瑒i��8?9Pʏ㟨�Iǟp�?A�'��B�� 9(v��x@Ȫ�y�%[�3� ����mJ8b/���Y�����'��ɀ�J4�#�� {�閡
�|��蟸�I���ty��$� 9ͤ0�" @L!�C�D
B�d�aA~��'��.��l��)��6`��P�!.�r�:�F�mX�i�#��9���Q�2(t����>��O診�nxq�bMFV;�9PE�s�L�k��?����'d>" c�>�@8���@=Z��h=D����ܖpM�U��͐^���0��;��尿�	qy��^
�z���5��g��g�m|��� �'��	ߟ���ܟ�q�$K��L(�`R�l�P�ָo�-��A�4�x	'k&P�������Q�>�
���$E��qKE���|�d���ꏮf�F�D-��E{�ɲ$�+�<����	�|�'F6��@	C�~��u��*/���N>q���0=�D��7^��g��i����f��h��t��_1u��&9t�*�J�CǬe�	ay�=)73�)�|���_	%W��Ag��D�d�(��1�?Q��'`p0���uF�HJ��Z=8�|!��	��e��1�V�Tt[2!�T���9|�����<��¶��+'`��PE.���Ƥj�LP
hN~R��?���h�Z�䆢9��(��OI$�����Q�p�@B�I;aPXbȁ#"��7��W' �?���Ss��ppTiH�'qL�'��vx��'�	�]����ܟ|�	ٟ��'~��H���GS���o��f�
��C�}�,q�c�/t�:�S�n±c�1��O�ܛSL�0N8������Vax
 JB�?"�:�I�%� Y e��>��I/)S��X��Ȑgɚ]��i��mʴ6mzy����?����r�2�B*1�T��eg�	�. ��⑌|�!�dӣ!�e���	���@k	b��I��HO��'����?gL�PG�d9���d,��ʓ�n��	���qB�M#l,�`2�o�1]$B䉚-in��c$�5��y�$�#j�B�		<o*P�$�P7��|� %�+1�B�D4Ѕ��ڎ�^��EL�=�vC��'�"�QR��eb0���
gXx��T���XBl~���$x�l]+r�� �!�1|��$&S6!�f8�u�C%�!�d����%Z1��!SΓh�!�D���	��%_5/���4v�!���>h�'n��GU������y�!�DDJ�(�xA�^*Ix�2.��f$ўl��m-�'[@��$�W��a�t�l�r��_iJ�c*�=5o�y��C�,���ȓ��!=v�,%!��XR&���[��iDGX�s�|t25�Є{�����-L���f�ѳL��@*�D�*�ȓm�=Å^/xgXl�$���9c���	�#�"<E���3��D��X8bc"�����-����P�_����5��J��ȓA�2��ܫWw \=wETE��
�̼�P(EE�P�%툺7�X؆ȓfV�![�ub,UYE80�!��uSv����`b]"D�[@�� ,����Z�oWR�RN�z��=�� ��;!�� X䲳Ib5NK&��4$�YC"O�9@G���#��Bc˟1�v�HT"O�����M�+���Iq  6[ x"O�Ȧ��e^�J5@U�
Eb����'��)�'t�P2O�>1�I��΀<{�'3�u�ׅ�N��i����zQ�	�'� !Α�a\ɱ�fD�~k.���'{�E�DȠ���BҞnO��2�'�5 �.W�0Xey���l�(`��'�<�;�����E*��.S�41�����0
Q?a�@	μUx�m��x%&��SC!D�T�B��8wlDp�̄�|���&<D����S�Vw����o@� 8)a<D��с�7
�H���n��� ;D�8����2S���eDQ��և9�yr#H�&/°��b@������N��?���D�����D���/<	2]�k�>IRN*�-D���a�X4��@	���<��A�(+D��x��2W���)
V�I�`'D�8��2~�Xh�>[�a1$�?D�|��`\�����O>h�d!*D��pV�^S����G˃�p�Y$§<	Ĉ`8�����VA� �7O����r&D�@P3�/8����a\�=t�h�)D��)؉t�<eYʇ��l�sR�<D�P�M�)��KŇƖV�~j�(D��J�F	������8(�t@cb�#�O�����O�͒�DH�&N�LzԬҀ1E�"O@r�O�;�<��k'��)"Op�4C�2h{�Kv�O�S����"O�H�s'F	mڔ��Q�	?<�����"OV�ү�\�|���	78�.�r"O���t㞊=5.9@�вP-�|Ab�I�Y�̢~"C�\c|Ii�D�|������x�<��Eʮudb	3G+F�A�lAG/[i�<��N_;gNƌ�wA�#R�^��FEo�<!4/״�&AJ��S�X&�5i���F�<i����W��0�V��M���X�i�<!�d�x�I�ΰ`I)��/��$�!b(�S�Ov��2�L2>�j(��[��r	J�"O�qTO�C^��
f�X�\ވݣ"O�l���Wt4����Gϰ'�4m#"O����%+��ki��T��V"O�	6G�%(%/��T�d)GR�!�Dڥpk���sf�8a�XA�e�<D��	&r���d�n����U.-ұ�ANV,f!��@��]˵��x&�U`�Џv�!�5F���Dj�#�4g˖=<!��Йg㐁�FkO8+&
���]�C"!��/>t�h�!��		FUɄ&�}�&[��~֍s"��aT.
�\�/�&`y	�'�R�HqL
& cr����4P"�A	�'��)��'��(�I�r���@	�'��G�|�D��0�NT�6`"�'"L�Q[�%{�K�Er�}H�'S\A+ck_
�^!�AI�3D�Eˏ�� �(/Q?i2kݗ/肨J K��Kj�K;D�9֣k@2�3��ݼ�u���%D�@aG���!d��""�h�"��c�"D�@v.ߏ[�ppã�T$V
����;D�ȰF�Ms�4q:��R>4�$�s�`4D�萂�W	��7 �Mu(�O��;f�)�^޺Lada�a� �*�B74��E��'�vx	G�It�-��&�3�H	
��� x��j��2�\�����a4����"O����UW�9Y�#�6:>�@�F"O�uaQ�(ܚ��d�6�dH)�"OjP����KJ�r�FEb�ABX���2$*�OƬs���fث��ѣ{*�!��"O��C4��(o��*d��}:̍:q"O�{vD��N|�1��c-S���"O��ò�۹;�ѳ����4	��"O�� 4�ٯS������Y�zU�E�'���@�'0��Q��}R�![7��?s��(
�'�T�)V�^	_T��a!`�'@3J)��P|���"��3ò4 df\�
��܇ȓ����d�+���f�X7���k�n�k�xd����_��(��Fe2/�<a����.[�ǈ9F{g:���Ԕ�&�Z�����VixH ZB"O
tpbI�I����KV,1�)iR"O:U��%ΐ8T��Պ�[���j�"O���%�E�drJ�V�T/7���"O�	�u��6��\����-O6�E�5"O��agY�qD B	'3�0- ��'�h ���`�&�WG)u��i�@!Y=D��ȓfZ����:X��g�T�cH�E�ȓU��A�N�*T�F G3N�&��ȓ+��y
U&Z�IB��0�ذ�������� ��2���2@���J�f9��M��9	ш�R�x��b�I�zrHp�'�� 
�o<L�{�� �*?���3LfШ=����8�ȗt�p��0G�3�-�ȓ[2.�i�+@���7� }c0e��)$} ���+�m�n1���ȓ]�pH �l2\��$�,T	(���	�+���I:K�a�aH=l�,�a� $�^B�"/��Œw���� ���T!G^B��%Q{�����(��S,G�kdC�d�BV$�:���'�	qHC�	�x5h��C�*Rj$�`�k_�t�C�&Oݜ	��I�E .��U��#Ӽ�=	Q&�H�O�pJr�6ԍ�%�>����'���U���c���f���v����'< |Y�S=~���@h7�ȝ��'&��%�B���؀�C$���'�F�"MI]X��g)U�i���!�'k$y�C	T�o
�c"�p�<���Gk��Gx��	N�2� �)zl�S��<6��C�I�� ��h	"����A��B�I�P���C�<Ԑ��KO�t]$B�I/'���i�[�z�ı�� �C�ə.�NdK�D2l���I��i4�C�-$
��Q�@��� ӍS>v�˓8��X��IU����F�> 4|���|�hC�I�̶�i�F�^Y&Й%(�;=c6C�	�Z &�2�	!ODR�� ��2M�C�6ˠX��̋7I�@���E��$��B�ɨ1���OX����Ņ�(
���d
�u��B�F��|q`��f�xъ��Y, �!�VL �#����q�%%;�!��L�<@
��ޕ1�D��eY	>�!�䔚<�h"�I�V ��ŏ�4�!�Q�4��e�M[.m*����e��!�ƌaFYx���Nĕ�e�*`�ў�Qƌ'�'6B��j5n����\r�R~����5�t-�f�G	���g�܋�P���A��@��[W	�����<o�$��S�? ,�1ElU#7+�p��
��$]�%"OB���[+�М��R�ƺA�w"O�y��G�t����ġnĘ����'�����E`��Z�e�$����C15,��}YƩ�'I�38��Se�`���Ӓ l":+�\�5��t�(ؓ#D�k�-S��XS��_Y�4�sD?D��1����`�"9HLrT� />D���B	Y.{V ����!6��¾<�-�{8�d*Ti�$?2ٔ
Y!nq�8*�!D���(V7kcD�'�#�ʜ��-9D��X����O��Ӈ�3�0	!/7D���ԭ�A�6�����7��44*:D�X�1e�0K�ʙ�@�V���4�O��cG�Ob���_��� r�F]44Dq�"OX�sF�] O2�ػ��ȏC�J)A�"O
��j�>"I�D�Uϐ	i�����"O>�	�lk�U��ԂHMj��T"O"� �B �{��]���^U잝(�"O`����uc��r��q�<�z"�I39��~���պ�Ft�g�Ha��P���K�<isO�Aq y8pΈ��ܬ����|�<�V�ˠ{4ͻ��|�N�r��u�<�A��AK4��C�T�T��r(�{�<A%cV:88����)\�p	@nUb�<�'ϑ�'��\�δ}�2m�*�?i+�c�����0��ӋY�����ȕUbD���,D��Y����BY����2�L�b�*D��� e�iE���tCX�4��Y���=D�����.?C�����փ]�6�hR�/D�D(#,_:*JR�JU�'�
蓱�.4���`.�v5��P�Ğ!C��4�eaN՟(�O(�Y(OZ�[�#��T���Y��˶|�p�!�,.E�*ia�̪<A��?��#?���A��c�j��ܠM=X�:1�Oݞ�2� HU�IÖJV������X98����6�ّ�/Ƽ9yb����zn����ɄwC|�I�)o��(	Q��OR�$.���Ġ`����'rTa��J��*��0?�U��:Hb�:�e�5qy"����`x�[(OH
�_8��"��c(b���Y�����	`yrQ>��I��af �n��49e��0�0Wԟpj�	dX�,;��99���Xe�N��h�
�3"�L6A�|�1D)Ee2���3Olزw/�S����O&+Rĭ�1E!�'JQ8�f�H$|z�"�0̓c��D�I퟈�䧉�DA.�D��1gʹĥ��o�$[�!�B@���FפQ`|[V�� 	�ў�Q��I��޵x��g���{W���=���<I�aѪ�?���?����ԟVИ3��^���C>u���a�N	M�K�n&��YRF�Q2���g��~��Q���=�^�db	�/��h����m0�0Ro�wH�<ˁ��_����`n�3�+��o���s��/w���\�d���O��=)�'��:,E.^�1�!b�X9�Q
�' j^�Q� �`U
���W��?�V�i>��	vy2˔$&����Q�
��(K6e�Fmt�'"�'p�_�b>��G���~�IT��ŖZ�.̙�t�S7�͘w�,���J�:f�*8��D+
 ��LL�-^�xL>vvx�Z3Έ'Z���ƙC�z��t:�� �h)�	�
�qiA��r���`��4CJq�I[�'n�8aũ¤`[r��%!œ "��;�,D�,�&A��K���Ҧ.�b'j���(�<y��i��Z�Ⱥ�A[��O����ߚ%��
T@�n���qtP��	��t�Ʌh,ЀT`�Y�����ּa��i�'0�ʝ�񅙬[,Y��FJ�e�=D|cQ$[b��͇�95�X�*�&7��Ɩ�.�h�p��	:�����?��O�Բ��'b�I\�*9���C,V��"ÏU�U��o�����ф*@�Ycf]��&�Iq�2�O�}�'���1b�`#",�aK������,_+�O.��O�pJF�C1H��5쐤D���¤"O&eQ�+���u�G�LN�B��P"O 9@�jݯS�hi�3#H�o��sq"O� �5Ñ��vX�@@�G�v���"Ox0�*)s/�%k�����`�'"O��Ф�>+x9��Y
ho�ād ���O�}�8��*��@�L��������)��L�ȓ]�����^�a�ș,r򆍆�}~���5�F ��|0A�O���O*�L:u��pMfL��/�n�1�ȓǒ��- [���;�O�>�Bq�ȓ"B�iUC������,zJ���	")�Z��$A�:��]1��]&-� t�b  �!�$S!`F:Œ� �Uy|��Gi[*N!�D���t1q�Q�Lp����C�!�DV]R���n�V]���`L$t�!�DFe�x��7NnIk3'I��!��aĜ�s@cN+'3�L
%�7�!���3�S�Ν3C.^�g,̯!�$�'���rw��L1�J�}!�DJ�k�����
W(8��Y��0!����
�Q@�ML�U�T��_!�Ƨ;F�I��K�^����MI�a���\�	t�)ʧ'�~�8�D��>F��R���L@�'2�~��a��� a�W% k��*��'Ȃ��J<���d	P+r�%ڒƨ~	��I�"�3��l?�"L�T>�	J��Y1��AX��IC!#_6DR0˒�W[~�B4}R��>���"�ħA�~� �74x��ā"���9�(}r���E��'(� E�G�)*Ν�6!IJ񾩓�#I���	��`X�'٪�'�.�s@�G�#Y��bB`µErx�ɺ���'�>�����c��@�L�d�`�[ aY�D�
�d�	[�Fd�0���Oިl��F-�`(�!(�>1R���(7b�˓y����Or�E�dDޝb7*I�CT�O�ZH��OыAM8�	���ҧ�9O8�c1��+p��9�M�营_-�Ԓ0&�v�J�Z��'��D�$�	�FT���M8KﮐZB�ӎ�?y�E��@
g�4?��yBd�'�~��X"d���j�C��
�Tá�S��?iV)�Ob�@Jά&[&M3Q��&g+n��"O�zbI�S�����<B�p���i��IWy��'�B�|���5��� U�M�&�4���K��ե�M��?+O&�D�<�|nZ�c�y���װ���ߙF��C�I�7Z (�En�!���
����C�w�^L��`�5k0��
!Ð�6�bC�	�^R���(Q�P	�$�6n��C�	�z���w�3}>l����^B�I3j@�XqeP! �~���ӆo��C�� t=�S� �$�@}�@��qBB�	v>n|R� 0�9��dªC�	�.%��In�-���wJ9w�B�I*:�̙kQ ��|�n��֧�E��B�ɨ@�v|)�mX/<����Ց3��B��'N(a��[�_6���"f�%.��C䉝n�Z�r$���!��Y�&�ϑ_[t��)���/8ږ��U�SRL8Q#��ؚ(���bc��W=dSKM!\,YG�@G<�AC3/��d"�@ǗPPj�B]�{e���M@;(}�̘��|?�5Y�GN�+J*tˠL��_�X��@�N�^�c&@���W� d��������ړ�ϥl����I>��A�eqN	�3�Y/2��ȉ#@�W�<AE�*L��2�Γ0Y�g��O�<QB��_��<��L؎^�´��/QK�<)��r)L�!��N*4�[v�QF�<y��=d�R}!�� ;k0q;��Y�<����,ReC��?SH��XV�<Ѳ��-�҉[��>���#��Q�<D�eP����O5.o���AF�K�<�gn�7=�Xx�/F�Q�8@$�E�<��ͣ��u�
W�fk^���^D�<���x��Hb�C;�^�c����<q���{�����#I#��ӌ�a�<�D
>
6����&��D��b�<� 
�k�..�Y#5�͡'�q "O.�+q,93�HAADK��"�A�'"O6� +*
V)���V�Y؎
"OB�M� d`q8� �6d��"O�!!c�@vzd�F*żY�6�j�"O�ȡ�de]|M�p�ݢ�{&"O�4iS&ܱ5Ҋqȣ�ƴ,��]9�"Of��g�<?UBͲ@mW>�|��S"O*U��]��#�����4e�"O�a[�ۻw�P�ĉ�LQ6L*"O��2�Q�v� ��^zF�h�"Oډ����b�*��&�K5nRT)*p"OJ�В��^�дq&FE�ua����"OJ���-���(���γ:{h�["OH|�A��"Z9p��H�atư"�"Ol8Y2*�5Jqn��МWyv�k"OR�#���2=֌�I��}YR�j�"O��Q���{j8� �G=\:�-��"OP̡5M��V0�	*FΖu���� "O�}���؏+̀� �͠%��<)�"Or`��Q�<��8$c��|�� ɥ"O^�۵e\�T+N�Xc4K���X�"Of��D�#_V����Y�H\�"O�	��͛�w��-�p���}Ҹ���"O ��f-G�4/aH5��&&.8a� "O>�q��;]d�%I��$��H�e"O��ReGU�A����nA�;�\��"O������%.�U��t���"O��Qg�bs������)c�`�"O�����U?@6k�"3x}�"Oڵ�`ˎ&VV;q*�5YfDC"O��w�a����*-> ��d"O�m9�H�YM�%����V�Z�2�"O0u��� VE�$-�o�V(�Py��
����1������e�<i��ȀYb�S�j]) o^%j��VK�<1$g]�\�C�hG"i�]�4�[H�<��*U�Y�duЦ�@(k��i�3I�<�w�H�m*e��c�j�D��$��D�<ɑ c�浉��/Cm� �IUB�<A�m���l`3 �*o�h�+FI�{�<�wHV"6aV�Jv�^~�D�ćC�<A�	Y��T�DBѦh�h�)DB�<cH�*>��'Q�" U�ҩ_~�<��n^�s#D�1AI'V����r`�}�<��"�yY:��W�_##>�CP��A�<��ۢ���#�O"R'����z�<�$�J/F���k�Qz�J���}�<I��B�XRVyɁ,(mR��r�b�<���C�Mh��w%-~\Q{!�VE�<�Vo�!;��y2��G����	[�<�C�L�R���+�+TQĜ���)�Z�<�G�T0�)���C"]�y���T�<	�`�G�0RЎ�<��X��l�<�"�E� ��)�Hη���N~�<`e�+F �� #
�`�&�w�<����1�r�{�ET�$�H �\p�<iƏ�>i|�0�LY���xG��n�<��H�dC0M�6 �o�RM(�^e�<�1�Ə/��u��A���#TH�y�<�FA4Y<@+�͐�YSشk%��l�<Y�Ҭ\Q�xx���	�Ca_@�<���O5�i�f�Z�%s����q�<yeA�9���⥫L(If)�n�<� ����1���h]�p�~�Y�"O��$+U�Goj���!�\���"O�\���:h� ��1�2y#E"O�\`�ń>\���Ꮢ26���"O�����0a�����φ�#�q�"O�t��Ֆ+���K"$��?f`�"Odᡓ�C<ZBpVlҨ$��"OV���	 CI�d`�ꕲHhM11"O�Q3�dG��U�A���&����"O�L��nށ`�8����f�
��!"OT�kb�D�/T��&���%"Op���e�#G�� f����&"O�p�G��#e�hȅF��\\��"O�Ġ� E����02CԨ4�Z��u"O�PI"�J����X��6���ȡ"O@�t�Oe��K���<:�"O"�R��-j�����C��.�4�"O<,0W��W�����G��4�f"O�i�6EE6�`)��5}��]q�"O���̇��ݡ���w�vu"�"O�������m���>��@*3"Ox8�&_)J�����M��å"O̐�fjJ:�T���R�g�!s"O��x&Nf2JJ��ӫV�M��"O��ڷ�U�p��XR��	[O���"O��j��:�42��U2�A�"O>���ʈ�=�pȈ3r�w"O|�Z� �+�0غU��3�@�P"O�ۧ���0��iZ�P��"O�t��O�72��	��9j 1R"O�p�d�����(3D\"O�@�""O��:e����T`� 5C�L"6"O������$����- cX���"O���b�Nސ)A�ǟ��>l��"O�r�`�@ !��!Ո�0�"Ov ��Ί/6޸@��ОX��"Od�b�l�%��Ѣtl�0��d�"O$șUI	�+ ��K��S�Q"O�<iQa�5F���ы��v2��"Oc��Ρ5ߊq��@&O)����"Ol�Al*~���a)�q!Z��q"O�|�/�
{M��`t� 	�
 "O��FǏ�R8��e�<l6�HH0"O��1Ms�L����	QB4B�"Ox���/@=v���k6MľVX~Ԃ�"O�z���]&"�L�mW���"O:j����
fd���ҁN2lt�"Obl��N
�-��W\2M��匔I�<Q��J�[��cQjԮb� %y�mMa�<Ar����i`���%�����[�<9�"ϩH�lQ��F�3lI��W}�<Y�Ra�,%�0��:N%�mp�$`�<�aƅ�P�2�j�՜.��ջUJ�Z�<!q��]e��1lHkF���a�<!g ��bj8���C� AZ-;6L�Z�<��,�$���{gD�:�^l�FhZ�<!���W�iKb��6H��K§�R�<��6,U*�蒏=�`�����P�<��]����YQ̜s�H�<aC*_����N�Fi,��rf�K�<a3�Sz��=���,x�# H�}�<�7�p*N�p��Z�S
�x�"�S�<I�怣%)���U�01��3 XL�<٤� Tm$�8C��7[_Ձ�r�<� $�xa�צQ��]��H�|o����"O�40��-hV܉���pY�b�"O�$��<����@TV�%aC"O4�p��8(�l���C�(8�`;�"O���v�4`�����n�N���"O������|��V�BY��%{"O�D� PS\��w�ƥW�|s"OT8�L�=��+�AX;��9(C"O(Y@��ÑF�`I&Ւ���9�"OB|`Q	g��ss�J�&�9�"O|�[�AՀ8:Mɕ@�`�(�"O�����	{c�G`Z�'��h�f"O�`��I=4'2�r�o���T��"O�kP��4:��'OU'�����"O���Mf)����a �����3�y2�	�TL$X��@0k��tn��y��O+}�� x�JE��M�1�T�yR,ǱOb������
��QH��y@Ҁl�X�OV�t���1&���y���e�:���I�6�tx8�mB �y�^΢�u�Z
1���Pd��y�CIJɔuAPc-���q�IS��y�T�s�	E��$+L�C��y⌓�0�QR���H��c���ybi�>V�0�f,ۯ(?z*c���yr(O�i��SD#ɒi+Ȉ#m�5�y�V�~�)���ɔc�,�I3���y2&�"�r@��-޵]�R��רR��y��@0[��8�!`{����L��y""۶N-���%E�{^ٚe�R��y��β:^0���լ�p���\��y�d�=	+r���ΖRl�t�E���y��/^���3I9!����/<�yR������Sq��"L�CBD��yB��n��Ń�9(�A "/ì�yD�.&�P�[F��6�0������y�N�^�㋐(|�����y�nV�%��h�4<��5˥`�5�yRk�.y�$8EÝ�2�&12�CW�y��F��H�9�A"0}d=����:�y�e�.u�4j�#j�aT	��yٟ҃�|��q���~�z�CO�y��	{r�`�O9��`j]��y��һmމ���R�1f2� �n�"�y���F �pIBS�[`6�y�O��)B�!9UD
�LX��x&k�(�y"�
qv8
� �-/���Հ��y��=8��<cB�� Ѣ�9�i���yr��Z0=R�%�RT3����y넊b�V�j6)T�_:��(�o	1�y�@7��tB�1X-|�`�dX��y­J�0s%�B�S;\��7����yr��;�ݸv�Ӑ]ծ��փ<�y��y(tX�%Z,ո�@����y���s���+d˘�Le�������y.O'ĩ�s���<���@#�1�y�a6��Р��	 9��ip��'O^4�eO�/�0��V��%��xN>)�aƭf�Zơ��U��Z�ϐJ�<)0�L+h.��{pJ�P�`TsE��k�<�c�>q�=�"`Dt�~��t@�h�<���{�f�����p�h�a�<)�G4Qo*I�/�$'�B�)�!S�<��V1?�(Dk�ZG*,��d�<)p�Z�M���yQ��Un���Tc�<� D�8�C��VA�G��,�t"O�q$�� G&p��
�k<�u#t"O�	�OP78��ƦK-V�8�"ONU����/)����'R�j��В�"OlTT��*ڢ� �"]���;�"O� Z�K6�#�g�Y����"O*���	�F�����h2�"O@���ěG�l� ��h�vX��"OHLz�H^6N� �ZQ�ʯ<�"8{�"O舘�!�=n��SG�N$B�y�"O�÷�J	zܲ��6�R*u�ͣ0"O.��� Q�g� 贂��X`��"O����`N�M|bY��FV�Y@FPy�"O���ʄy~�����ƵI1"O�ш��+� ���46�=�"Oڰ8�A�c�f�a�����m"Ov��v$�ko64�EF�#��\��"OR؀0��g�i3c�@�W T:c"Ot���Mծ#{TA�Վ���@�:�"OJHQGGّv{n� mY�"q"O�M�r�;4�iGL�
C�8�a"O��W�Q)b��L*r�B�f� X� "O��q�>)m Y��D�z��*r"O�KfL�gr�cDo?�J���"Of]�$��%���ÏW�6���"O��Cw��w�Z�A��]��1��"OJ����V�� �fO�fr���"O�a���\�X���I�e@��"OZ�*��Ԉ>�����ƶp�bhK�"OV����'���A�-^>G�fy�C"O��J�`ʝS� ��S��$5�&�C�"Oi@�ڂU�T�
�7m��آU"O�D�GB%:ͨ��X73�Z�2P"O�2��#����LΖ-LB��`"O�]�v��c[��	�&�"L #"O贳'�A0K�x��i�*��"OX��oB�"4���_+��=�T"O@	J�N	?*�~�g$Ϗex�8t"O>�9Sb����쒥hE)P�k�"O\-��
�"�b��6�WC�F��0"O\hy'g�8ؒ���]�Y�H��"O���,Tg�lfhܲ�x�a�"Od�a�]-��5��-Q�^���G"O��:f�:DȒ�j��*A�c�"O¶�8J:���a ��<ʐ"ODE� Ɍ�6rf��f�]�:I��R�"O|�a�F<qn$0�@�.�nP�"OL�21CTY{�'�5���J"O�h���\��違�ʠh�hEb"O��&`�1V4����!A.ug����"OxIqc��))�Չ�,<e �0"O�	B�G�SYz,��OǶVK���"O����Lإ���X��	1-�`!��"O��/B��J4L��?�D��p"O�)����y��$B!&�P�h�"O�)��-6CR �9q��"O
ԣUJ�-Xj��Ҋ�K]��Z"O���W���(���	2���f�T�P�"OP=��AE�2p'j�$4��*b"O���W삋[Q���T/�&:뼁8d"OnP`F`�/NX� � �;tҤ�[�"OX�觢��i���¦�0>��"O�y0��3x<c�� i$�x�"O~Ԑ��'���z*	�_�s"O�   p�B�+�J��@�X����"O���6=)�E��fߘ[����"O���� ]�z�.4�$ߡ7~�Ѻ"O�����&�U��*Z5�Q��"O|�� �D������(�c~H��"O�p�iΫ' �ew���7!�A"On�"6�[,q�D�g �u�Q6"O��B3k��xe�I�i�w�vI�"O���@��ѸS��3y�ĸ1"O����nZ�~e�iK��������'�D��닉��p�V�5Rx�9�'����%�Š� h2�lY�BA�	�'���2Ñ��p����;��$H�'Nd���{g 1�ucR�Ob���'�ri����J���(�E��'�R��5�\��+t	ݴ@��X�'<j�rw�IL��2�L/t�9!�'�`� �1fFi���T�s��4[�'�2�(�#b ��s��K�7;� �	�'j�i뗈�7Y���цP*�`��	�'-��b c\�f�4I��]�)����'�&�cw��" ���A�[�)�'[�ي�ҫ#,�"���M����'誤� �E�8���p�g�C^lؑ�'�@]A�ZB@��&O�G��Us
�'� y����X�N��1,Y{F`)��'�  *��u�����k8$L�'�R�:`đ��&�����fMhL��'�&��Ae�*s<��Xt&R��.��'�<� ��&Q>�2��֡�S�'�D�k�*��4!�8}�� �'2x�1R�*z
��ߑ$J���'#�p�3|��]��&�k��|�'�T$
�b��1t�D(0�>���'ʤ�\�O� 0o��[t���'�n:qH�?Zg�ccb�d,���'�5Oͽmr�I��T&*&��'��S�����`Q2�^�C  }�
�'��P�!cE2%���E�-
S���'tԴȶ�Rk�2P�E	 ' �'��0��΄���y05 L P{"���' �����4��i�g	J�D0�'5�u��׮�h�4�Q�t�T݉�'I����F���!��\::N���'��Yĉ&e(⼋C��i�����'X�!*�GI$�հ#d]�b����'֘���$�F)�\�D��	\�!y�'���0v 5v)�%;B���`r�'R���&^�����ed�&�~\��'}��!W@ʱy*�r�
^&L^̩�'� 23�����$d�K���'�j�K���G�/{°A���yB��2a
 �q�{�j(��y��X�(��L�a]tv�9��I�<�y��Z�LG���Hՠq�4�c��-�y&�t�V鰆-�m���C���y��34bF@����<G��0aD2�y�C�{G�h0�ֿ.>�ͺ#�@$�y�h��+
聅�Sb����k�&�y�(���2��U�4�ÅB�yB�S�2��X��:�����<�y�Eō�H�F��~yr�E��y2�ֹV�.���ɁZ�sE��-�y�P6I��xr�Ĩ=~4��%�*�y
� �eᆤ��d�e`��g���CU"O`XR�D<��a��!�xL��"OlP!�P�6q��PoÚ8,� H�"OzP��([��H�%�H;�"O$m#K^!s�<�9���u"f�1S"Ojʁb�:?
�ٲ$�N+%"�̲2"O(�&��MQ%��^,����3D��
`FIs8���̘[Q��2D��#�m���)aE�*Ǽ�(Vh;D��zu��'k.��q!'Yq�L@��9D��CO("|��*NY҈�!��2D��{�g���F|���A,'�YQ2�?D��:Տ�sPT9�`�E!:����`?D���۵��=�L�LYx���O<D���'W�eZzud *�<pq-<D���B�֟y�<�5jEYt��!<D�x���9��	'�o(8���;D�ȫ��F"+�Q�Ԥb^M�f�+D��8bG��� ׈�0R��`�<D��H��	�,��UyV��X��QD�%D��kÄSby� I�"��s�ވ��g$D�����?��dZ&ӵc����5D��2�ț�Z&|��ѻ`L4�Ҏ9D���dB�/
��P9����K,v��&D���āŭ ?�X���a�b���>D��;b��oF�S�7�@�(2D���Q�ƗI)ܸq��Q�D�xE�7�;D��1� �**a�X��E�,>V��'8D��83���Qq��@���gj�	�2D�1�m)�������C��>D��P��ىB{XY�UO�$]cbuR��<D��$'s�%�ƤI�0i6� X���ǷZ�\"r�$�
q;�@.�y ��>�V��A� ����B;�y��(jS��'͒�r����Py� T�0��P:a'�$)@���N�<���T.y��&
� d#�h�C�a�<)&g6Gf��)E>jK]�w�D�<��o�04�D	��n�b�Rs�E�<Yg쓧p@kO
�8ݪ]���XK�<��N�[��0�(]�k-�����F�<	E(C-(��h׋�>8�<���]�<�6�ݍb�L�Z�(����@&R�<����@Z����/�T����OG�<!��2]������T�`��C�<�у[�<���e=��d��\�<�ƅ]�jd
�T�pd�((e
a�<i���n����#@�C\``uJ�{�<yR4*K�@g\8�:�t�<��iC�p�D��k����S�aWZ�<yTj��v
�y��
�_df(S$'U�<)����HVa&}���8GIx�<ɇ� 8a_��:/ΉO��pH��v�<��{��@�BH�+h�(���O�<����Ol���bI
K&�鲨6T�\ �b�	"a�W��K��t��@#D�,P��Vr=���$��E@��Ѥ*Oq3Ul��)�tq��l3����*O�T9�`G�]��8rR�O�>��=��'ը�މ*�"%Aw�ѐ�� ��'/f�3�A' t�&jõo� ł�{��ҧo���{3Ǖ,b�8���&��%��Za&+{�p��h��%�Նȓ`��ĸNպ�:��s�ĥ�jM����P; _>�%/�v���j&D�� ����={�M���>1�X�"O��9WK4j^���G	��l�T"Ol�(7�V�.	�qM�A�Α��"OjHӔ,H�)Y��@��'hI\�p"O�`S�L�X�v���c�C�!0�"Ov�{�7
X`P�cl5.�(�@"Oq�$�=�h���N�YGBe�q"OpQs�L����M�S�*,���"O�x
S�-x��bg
�T(����"O+�J�k>YQ��֙,)�-z�"OY3UD�.`~�� �ר��R"O쨘�-]4F< �HF�]��frq"O�{Ё�4t*8�kѨ	��H��C"Ol��+16�a�Af�2*��a"O]�����l	SƑ��^��0"O��j���qAR26J�s�$8�y�-�F�Z�:_�$Ca"���q�'����U{Q�ݺ C+s�8���'��9j�煶3� pJe�Bm�.0��'y@�b6��"E��lؓ�ް�����'���!� G�$QR��
��-�'����$��?U�AQ�G/yٶչ�'�H���ïau�ղaCۜ��c�'�JY�T�݄Y$�bǡe4�C�'
�@����6. ��EK3qp5X�')��]2iD!��B�>1�aC�'t���
ǝ^�
Ы�I��}�
�'���Y�o�9FB���oG+}n$�2�'i޴ৎ߬0�P�+�bG?��|�	�'b��4)�R��}� �9�\�*�'ߪ "��C�F_j����%E�ҽ�
�'��r�F6.��k�	�h���	�'@����j��%!�!$`��R�����'�r����,:� TsC�@:n���'����C��?#�����U9/��1�'Yd`4W�U�j�k�%8�X���'���1���+��Q��
+Ϊ�s�'ʰ�sҌÿw7��ԏN�"�ͨ�'�������z �/��i�j�(	�'�r����|� ���Fd;6���'�$eEޘG#`x�(��Z�-p�'h�%@��V��������P��Pz�'��&��=zR�h�~�5a���y"AU����(��C�e�u�7�y�JVDY�]���4���T��yB��$�T3#���V�L���ybÀ�Yo��!'L/y�@�(�L��y�c�/m*Ɣ[�" �Hl���'P��y�-@�Jo�!���$H00%��NM��yr��>p�� sբ�A1d}Q���y�%�5<a�H�6�¸7��h2dM
��yB]�=��$�E3S��h���y�k�v ��g�·*��q��H#�yb�P*sd؃C�dSCQ��y�M��[��=yc�ɺ���1��ܨ�y���VhXE3�(�[`���@ˡ�y�k_n^ �b�b�-K�X�	F����yd�PzАFۋ;O`e���H�y�۞�C�� ي3���d�C�	��l��c��(k���W��bE�B�I�y�"X2P�O1SX��2U�V�k��C�	�A��'��m�n��F�RaK
C�I�$��@��F-�8�A9 1�B�#G�(m:�V3a�|Y�H y2�B�)� v��!tl��1�MɿyTx�j�"O``@vJ��{*�A�W��6^��h"O��k�/٠Vk�y��J՗*w�D8!"O��h�Ӡ�ADp(,Z""OB�bOS�����&!c�"O��KY̊��)y� �"O|H�GKG��r��H+g���t"O�Q���,A�츥�ٙ'L��Q"O�
��X2�Hi���>���"O}�SK��5[�iR��2Tq�"OF�Z���E/�aW���U�D�4"O)@FعTz� �F��U"O��i0��@��(�D�o��P��"O����/�0\�2�"iN�Nz�mH"O"!+dEF�&�*�yѱ`�mj0"O,U�hæEi�f�?l���I"Oм��'�x*w���b��#"O��[ĊR����Ȝ�dX�"O,���;=[ԍ�K+0��%1�"OX�2�PԤh�q���	HzT��"O�u��hL�'$�HS�A�_)�\8�"Of)#�L�rո��,>%bqqT"Ob�{fl���k��v ��a�"O��R!�4j��L�J.d�Ib�"O�c��`Dޙ�W�Y�hXđ�"O����_�*z��.��	>
� "ODu��	��$�p&+��H^��"OB�"MC�bӶ-	��`-qrg"O��Hen@4a�"��6���t5���"OTt�IQ�9���!c)�Us�"Oj\���ѠAV"�s�گy��"OT�e*F�Z �ܡ�.	^�򸁐"O6]j��.iar	W �2ܶ́0"OHP�ϴB���U!�.x�"Olщ��;TZИ2�s``e�"O΍���ƴ{�YB�HG�t��a�"O���:l�a;
�
J�Ĕ�'"O�M�� =+��<а�_z��z#"Of�H���d2Z$��$�4�2%{F"O�h�qf�_�4c���c{x��v"OJ*J  �ڐ���ټ�D�yr"O� �T��X4I(3 D��L(iC"O��5�/{JP�������D"Or[�ĥXCP2o̲b��X�"O��P�;j�\H�̜_� !�"O���Q��/��a��TDRQ�"OP��g�ZI>	��a�88P�a�%"O��K�)+����݉w<�f"O:�"�
�rV�@�DƱ.
���"O�I��E�{^�*�]�]��h�F"O�y���ZL���9SA;p��P�f"O�e7
�<���
u6`�"O̥X�̔@�h�2�:c�e���'dў���3D�y��nK�?���;�%D�$j��>.�j1z��ްXǚ�!�)"D�$Ⲡ� A�tӅ��V�J��F�?T��sf�w�Bh��͂/s�A8$"O��dѥ|g�P��	GVE��"O��_�`x�3]�zYRRB�3^�!�dI'��!+AMXv=j���A�4e�!�d '?H,-������B�H.!�$U�9�q�g���\р��i�!�T���C3��#u�%cV�8�!�ۀ_��p��$r�y�4d�'�!�� ���фS�QŦ	�%[�N
fuH�"OdQ{�!�0Kc�S����"Op!�2��"I��)dc���-�1"O����G�^�[gC
<�M;"OzؖK��:�z�1�2ztX!�"O����������įtn�@iv"O`�s���-},�MâhE���!"O�0R"��&�fA3U�$w-����"O�! N�F!#Q�֦6��D��.D��i��܂@�a&�Ҽ\1�fB7D�����̃��=�A�`��ৌ/D�\��@pi��	k�`b�';D�`�B&��Q�"eΖXƌ����9D���g��x��=J���6
�|H��M%D�|����%Y��՛��@�bx!A&D���B���;�9����̘)Qm#D�L��f )̰�pumğu�z9rt�5D�,X'd�E$:|0&��y����'D�\�3dVZ���B�&Q�M��1%1D�:[1@
����T����0D����i�N8�
�&�,�� $D�Ze �~|�����k�2U�&D��B�ɇ1O=`!1�W�c�R�#D�p#�I	+΀���V�e�X@`�,D�((�ɟ�X-6��i����ʕE=D�H`�k�d}:x�6iScZ��pq�'D�4�/�) ����6kO�$nL�2�7D�l@���`1Z��S' $:+v���7D����(�.�`�"��8�^�@0D���EJ��P H�8���/\J����g)D���w�)]�"�F#X��s��9D�������T��Q85��	!x��Vi+D��h�4c5�p�o_�pLY#�c*D��dB]��P��	E�t�{L(D�,RP  n���Z(�b< ��;D�3Dm��\�
4��
~o8S�:D�P�M!�6䡣��'��@��7D�X�1ĩ��%�`�h]
�1SJ)D� �q�Z�S��d+��de�*&m:D�4�&�7o��J����� 0�k9D�Ӆ$�)0�j��_�AXn`ye6D����Q6{u�8�ń�#NJ�5D�|X���I��-��N��q I��(D���B�%7�،�B��^}Z5 �L(D����@O�Qj,�U�D!}׊s��!D��a�DE&[A�-I&�C�C1���Vh>D��y�k�*oI*� �N��m����!D����o�2%>4#d�dr#<D��C�\�l��t ���V��IsP.D�\tM�*��mp �����y�R�>D�PiԂ��AL�z��Q(a"i��O!D�HC"�A(F_t�R�,B9��A�%:D�,;���={�S� A��@P�"D�0q�i�4
�Z7�O�4M��0&�?D�lye�҄V#"��g�ϼ	ώ8{�C"D��wƛ�y�Y@7�L�Y-�	�3�2D��p2�3b��T��g�T�n��0D����&�J(rB�;Wu6�a`3D���`��ak�	9vC��0u2���B1D� ��`!_3��R4�]0	�� f�/D�Y��������)\�|x�8D����	�"c`( ��E��f���7D��J���:�X���@ǟ>J�x��/D��"��jAp���ٗF}X���C.D�� ���D�o�ȁ���"�X �"O&)�#D�	�p�q��щm�����"OLę�Gݾe骩�Qo�0�r�#"O�DѫSM���P�E�d�D�Q�"O~ɠa�� ޘ�s�--iu�,��"ODh��F;V0� y5-@�&�����"O
�1E�J�I��ԐD�V'��yqp"O�!�Q-_��9(+ضS.R �`"O�z��x�R0�
h)��"O���E�%.���#ш�%L���h"O���qW�`�Z$f��z�6��"O�,�.X�
@�H�F��[��A�"Oֱ�C����z�/�&k��L��"O�\�ޛ}�|��&/��3�^��"OL��� Nx
���6|�B���"O�x0�a
,�:tJ�σX�~���"O�=0���;����@D�0ذ�ɑ"Oҵ�pB \�lI� ��n�(�"Ox��FmGX�P�(��1�b�
�"OD�U��'aR,�R�B������"O`5����&���#�l�W��"O*Y��Ԇ��X(pO(D黠"O�]A2�3|k^p����4j��A"O����޹.����!�|�"O`L�(�QI�h��.VT�Z\*g"O`��AQ(��U��n�3~����"O2l��k�;`J��lK�`��"O���aL�x;d��j	�1����"Ox��#h�(� <�� �ru����"O(�`ň����=��$�-\"��"O<�bpa�
j�n��7�� Z1B�'.�L��ƞ�-� �#a.�?+ ��C�'��,�mD+$0F��A�.7����'�<U�0�Be���0��������'?�t�t"Σ
.^M���\4*!)�'u��@�@L�.�v�"�L	Nb�p�'�Z 2���^f$����?�T��'�*d�ᒹU�P$�?/�v4�'���	cn[���QjA�,�h��'I��!��H�:T�&�ɰ�h���'qf�҂(�[�,{ƫ�(}i����'�4d�D
S8��T)^�6�0�'-����LJ�&0��"Vq9�'����e��R-�Y��ҽ)�4�#�'�L�`�	��ܱ�3D�J� �H�'U�j�������m؜rV��
�'O|8��+�Gd���
�'r�}���]���rG�WY����
�'r>����#~�T��������
�'�$�[rjU�v�L���g	b
�!
�'�쵨7B���Z��Lr�,E�	�'����3���K��e���	�'�Vm����2/���G�VL	
�'�ȍJs��?w@>1��+R7�M�	�'�\�	��?_rŐTd[%�2�:	�'��e�w��/�H$MV!_�v�`	�'��L�D�OC��C�ڎV��%��'�=!���\�2!Xr� E��(�
�' �|���;�B��t��3�|���'>~���&�6h,�$���:���8�'!��KF�P
�8d�G�v�K�'����Ġ4Q����@k�0�����'D�l���S6V*��`JD�^�V���'��!	1�B�z�e�SȾ���� 2|ȷL�/2`P��� ��ы"OlqX7�ܕ�V�ȗ�]�� U�"O��`JD�K�Dg	'k�����"O��t �攘U��/
�(P�"O�q��%�/p�԰�֓R�9��"OB��B�W,q|\���áOq.� "ŌseHכ|��f�
o�|C"O�%�iǶ9�!��%T�)8� B�"Oj��uI�]1��"��5 <r-(v"O����jֲ	9j�� �R "2F�ғ"O�(�k��`H����@2@���w"O$D����q"�0�D�>.�2q�"O4��"+G�9	�� ��0`�"O<+���<����h�*�s "O��N�]Gx �k�N�ֈQ *O��6�âZ �2.	�"���'�x�IK1O0���΢`�'�t��cçI���!�Z) ���'�BA#E�C�P�h��ʄ�P)c�'��'�
>H��ۣ�J�M��M��'<�BRIW�\h�s��$7�s�'�8�x��`N��ڣ"�@�ԕ��'UN�ⲀDq���,ĺ1M�@��'��"˛T���
�Y(�`�'�
d�ՌNd$E/YN*��e�n�<��6e�V*`E�)�6YI�DVg�<9��`Ậ ��M?V,���s@Xa�<i���2��LC�ɱ�$����_�<��,iR���b�l�P`J��Ww�<y��wMV,�5,L!�Mb��V{�<�E��qJ�@�d���x�@/�\�<��>;�x(���B:����+�\�<i$��e <2W F�*	�u��HZ�<��4�򹲴k[�c�������R�<�cMH�r�%������S�<I��@\X���.O��S`�Sd�<iAm�+�$)�`�"��C�B�^�<���*C�⍪�!��F�@�ZEG�s�<ɷj�,DK��d�a�e�<	����I�pBU��P�L���_�<��+�3g�D����Oj���yq �Z�<1 O��KH�À��SXZ���c	[�<y��֠(��r)�+=���
V �|�<����t��8�s�S���J��S�<����8��fM��P������J�<���>|�����3e��"D�I�<��MH�仳�:S+̍i��^D�<�&	�.�FU˰N��e9��P��}�<ap'�m���R�����c�A�B�<��A�z�6!kRHE$��I;3�@F�<`�!k_�8�J�(��}3�N|�<9�ߑZI���%��|�P Kը�x�<A�ؑ�N9�#*�WBf��h�z�<y�*@�M{@\{�� ,a�\����~�<9��B�+�O��$���b�<�"&�޺���ATv^�a
]�<��ωm}~)ɐ%\+�pDib�Jo�<	uNT�(����O�ZZ��ԫ l�<!.T!�ra�Ck]�a�,��OKf�<�c�E.z*��c`^�I�p��c�<a�C6El�<�7�̴��RU�	z�<�j�)U0^����׻Q���u�t�<� �K��r�0rh�9��H��)q�<�U�4����ԉ��dM� �'	R�<� ���#��]�2�a�e �<l�K"OP�hЅ�6�B3�<#ȹ��"O`�
JX���!LԌ;�"O�]��
�/����$���GX�D��"OT������A��3g/�3�ɲ�"Oub���	� eႃ٧Ɯٱ1"O~ �DdĜz�|R�aX_��Kr"O��Џd"���@k	0R�(H1"O��YŃ=�3e�JQ��Ed�<���
�2a#�[ٶ��� �Y�<i�6k#n]����-�dh��T�<Q��%�* �f��dI>�KF�J�<���:r�3�o�e��Q�<�5�D+$㈠@���v��W�<��Cn��Ks��|z�VQ�<9FW!��s2��+F�!��c�<9e�TD��I ��!bQ!�JE�<�f(J��D����H4F`�\
EOPC�<�	ʘM��a�'�4v!��U�~�<AwmUae��ht�@'D�n���*�R�<�&-�>��0�f&$z��"�M�<�B���s��#G_�r�9���H�<�!jH:�THW���q%��AG�[�<�tdZX�����$��^�<�S�$L�<	�EUs�p9���6P�V���@�<qk�=q�-���0���J�R�<9�Þ�pK%XW��"��]3ģR�<���Ʀ
�,��W!N�\I���X�<1�L_20�	8�m�*V%�b��T�<qQ�P�0ѼH�Bg��K5�=�v�N�<�ଋ�rUh��5ت0���@h�N�<�#O��h�m�25΄�!Je�<�c�+;D�e�Y�X����&�_�<�@C74 �h��h^�\l�aL�u�<�6 �!Y���P��T��8��J�<�B E�1��[7��).,��fE�<��n��d��S"�(�x�h3�Rg�<9X����נލe"BE���ùS��C��H~�YрQ�
\��
b-߿l<�B�I�8'��e�O((�l��#4�ZB䉤hR�]J�`Vv.b̸1��]0FB�	;`�vo�0_�N��� ����C�I�|Uඇ�]6�4����<�C�WA��e O,��a_?"rB��_vFěE��#�Kr�E��C�I"F[�XS���0t�� ��%|��C�	�g<�v��+}jj`�ܕo�C�	$|���q��2(��V)	<HB��w�@��+��A����&���:B䉏�j��֡Y�\��m���T&u�B�	�G
	J"�L܀�K0��I<\B�I�=Pny��`U<h�`��!MJ B�I-n"�����]�!HP�)�kĦAv4B�	�D3���ҫ�-:.x��?9>VB�!��h�&[3R�2�J�,�12B�	)�N4�Ej�?����NB�	(�*���l���M*DC0C�	v��L�	��{n -���9@fB�	9P�m�&�ʞK�.42"�W�ya[�-���{���$G8u!"l^��y�)DK�j<�h��,��|i�ǌ&�y�e {8�p�ɛ�!�<��O �y2�J.xyZ���r���-�y��&B��58�/�~���)Ϫ�y
� �C�ȏ�Q�li �$��(LD�Zb"O�9�!F9' X7E9&���"OD��Š:�,(�ᬃ*-9��a�"O:`�!<2�� ���D�("4� $"O�X�'��.|+��/�@L��Gz�'��`y�Tm�X�'c{n����ߥ ���$M�E�ڽ06&Ԡ|�R�'(�镖R��[�Oӭ	�V�@�� ���'%�F\���_6Vt:� 
B$��Fz��ފTGn\��I�oX��
�I��)�e�B�(�9C��^�n~�)g�ØB,p��dNnb�'m4�x6M��"�������*�d�b�$+d���[��"~�I~Y
}{$@��D�0G��8&����¦YQߴ�M�ɛ�O}��� "�� ������Y?��ٛ��'��i>�8�&H�,�I���A��W�(���#Ù`�J�s��HiB�0R޴@p��A�H*D���Wܧ��^c�!���h�6��E"u��3�4m�f�"�K�Y��1 7��Ǧ�[w�_�ZA�U���\c�ld+w#�f�R�Ƶ �P��4m�n��	ӟ|�.O�D�sӶ��@�^�q�p8i"cI�j�B"�O���+���'?�Ѡ�ǒ
�}��
68ز���D��m�ٴ��O��N�_�^Y�5mRg��ݨ�+]:jf���'�*x �bёt���'6"�'0:֝z��oC�t�F��D����L8����<B�o��&p(8�-�#��`��O�DԪ����-J$���̞`D�U դ�7]��1�ɩJw&�X&�Rd(��20S?�o�W"�%���	K�Ci�i��f��? ���C��?�ƞ�?���Ei<�gyR�'���0���Ɖug�-�f�^���h��I.,�v�S�䅖k�Q�c!��M���:E�i�6�:�4�����<�퀬/�v�Q���� � �E]�����?���?Q�"���A,�J�d�K��K2�\
X!�r�W�,�p����P&ky��6�ݳ!���(ڗ��O��� ��)�\q�� � 2���`F^�꬀s�.R�>`~�#�I׎;:mx�i�'����D�OD�*ǪW�6�l� �+�<{���3*_�>Yl��t�'���T>=��D11
��E ]�>��-�G�#}��)�S�>���RT�Z�$��-�A<
�
���M���i_�ɗ9����4�?	I|ʃ��#U�*��g�R�S����e&K�< ��Q�'�b�'w"��жi�~�S�j�?$�$�:t샍��ti�O
��u�Eh2qR�a���HO*D��N��`�e;愊���)k��G�K�����I `~��@1kV�~z�8���#kL��qd��O����l�Ҧ��sl�3(fHP�H�#�ER� ���?qJ>	�S��?9-�>t�d���RLƲ4�'�UU8� 3ݴ�?��4M�(��L�P���x5�ʱIn ��#�z%V�앧�䋟�W"��'q���\zf�m�`���N1v����Y��<3'0�aN�	[q�Pؒ�
͸O.�d���b)	�r6$�����I��i��L a��b,�T$3O�In��,�s���	Y1u�
�R@&S�)�v�XѤ�>%+&�'��-�P��0��	�����O`�{C@��vYq�？ �	ܟ��ICy��'s��$���0=��H�B��P�`���I"�M;��i��'at�'GQ&�XmX7�`�Xš_�1A�qT�|��'����� ��"O`09��4�RXx��_K~B���"Of��T�&m��i{�(��tk�=��"O@�����?�Ƥi��4Uc��D"O<�PAe��^2���gWZ��7"O��ʁ�d�*9C`�)6�%Q""Od-!�����t�Q/L!p��!7"Ot�{V�7fm��M
�T��w"O� ��Ik�:4�FuI4��=V�b"O�D�w��%��)Y�A
r��"O�@3`�_/6(��
s_(dN)2r"O��� �x���ES�P���"O��I�ZO����j�O�4��%"O�5�«
�`������Wb�dH�"O1���z=� ����2'�܋0"O�1����4� py��	8�@�*�"O�tȃ�Z�a�V��Mf�@8*t"O�]1Q�D5Lf���P{�icR"O<�zr���>���"@܋d`��ۧ"OX����[�2Uxv.�'D��0�"O��+-��8�FL��
B(y��HW"O�P��(H4�p���3L���t"OD`ɡ��+]E>�� ��6ED��u"O���	�.�A�ă�m4�8�"O�r%%�X���s��>��f"O>��d�� �����	H�x�"O��3F�!8cb���?�B""O�4��20��t�V��B�raXT"O�KS�C%K�,x#[+R!0��"O�X �m/5�r]�Ԣ��=l�A"Oֵ[�Ü�K[X\��A�2C�0��"Obو�A�8D�Y��ҷ72ZxZ@"Of�k��?zy$ �t�F-�Đ�"O� �a�][+ Y]�)K�Ϗ2�y�	P=V����_{�ْ��[�y"�OC4)���e�VY�GB��yRF�m'|]�d^�d�������yb�*/�hs�]�Z��d(w#�4�y ٛwT|��(�=X4�CN� B�I��l�" d���d�'��$N�8C�2e\����C%,F�;�LC:��C��%|��؄卸L2�[w��u��C�&M�1��-�F��E E-�\C��8�^Q��D�8rG-����uC䉀:�Q��
ބj�2-�G¨WC�I.�����@�^L4�@E���B�SUQ��!�8��a��S�`B䉯{T�\�d�>s�v�rO$t�8B��/a��a���-t�C ��gU�C�	�Jꪩ!��O�u��)CA -=�B䉑I��6΅���uX4KK�.C���4Qj! >oyЩH��D�@� C�I33Cd�   ��   �  ?  �  �  �)  5  E@  _K  �V  ,b  tm  �x  ��  ��  ُ  ��  ��  M�  ��  ݯ   �  ��  2�  ��  ��  -�  ��   �  w�  ��  ��  N�  � �	 + o �! �' </ 28 �> E OK �Q R  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+!��6*\�c�<4�d5h��'�B�'���'	�'/�'�B�'���U�W9��m��Ʊz�0�b��'���'�2�'��'�b�'�r�'���k��.Kªa��͎ 5���Ha�' ��'���'�R�'���'���'����
F	�>]�&ΏfEP$�b�'�b�'��'�B�'�B�'O��'�$��zm@|XpjC�6�D�'��'���'v��'�'��'�"1�)ֽⲵpa����j5�'���'���'t"�'��'��'�%؇�Δ*��� A�B4%
0��'�R�'��'o"�'�"�'/"�'�f}�b���Xs���]��X��'iR�'���'���'��'W"�'g�=��'��"��	�Jw���'���'j"���d�'5r�'}��'��u�1� (iL�\r6e �t|:\���'�'H��'J��'ZR�'vr�':h(uC�=��)��G-P�����'��'u��'}��'���'u�'�;+�'HhufUmzn��`�'���'|��'���'��'p��'�J���R�h�����*|h�p�'���'��'���'h2�h�x��O��"�q�R��t�T�)����G$�|y�'��)�3?	��i�&��#�Zyf��B�º�1x�I���Ŧ	�?��<���i�X�p�ޚn.�R�FO�D>����?!pm�,�Mk�O�S��K?�Af͇2m����K��CS��ą6������'��>M����I�,=Y�fɝ��Ud �M{&%�e���O�26=��H�N�:Hm�y��[^|<	���O���n��է�Oj.��ѱi��R:28Zݢb�"bw��:R(�3��$t�$*�#��=ͧ�?��&ޙC��Y�S\)��<1,Or�O�Em���b�����C�R��f
���"$��Q��o���ޟ��I�<9�O�A1���X�`,�wf�;��"����	<���U�;���B�����z L�4�*H��M�+\�����my2U��)��<��%�	|��0�K��)��i��	�<	b�iV�|�ORtmP�S��,P}b���J�.����g���	�x��5��HmZG~"1��)�ӳ@��˔kJ>L�b}�Ul��Y۰�|b\���8�I��,�I��H������eЕgB �P�[Dy�Ooӎ�2��<���䧊?1 I�D+!�e���E�Ȉ!�N�<�����,��L�)�N,�*����d(,�Ƭ��R�;Ej���-O�4X���)�~�|�_��!��������_�f�.8�!��ܟ��	�������{y���Ox(1��'�����ˇ�?}l|K�O�A�aR�'�~6�.�I-����OB�$�O���c,��£,į;��#C�&JL7M$?1��J��I*��߭iN�F����uq0����f��$�Ol�d�O����O��$<��Qv���h�`K���C&�@!���	�����/�M�իK���d��&��2kY�1\*�����
�촑P)@�柴�i>�c�`�٦��u�n�,���������FJ�{l�-����q�	{yb�'�2�'�R�{{��*mˋjm�JuO�2hk��'��	)�M[p�˽�?q���?�/��|a�⇽l�.t�9r�	F�W���"���O���&��?I��Ik�6mS�lG�H��i�Hɑ��(Kf@3%�N��|"�L�O���J>�� �5|�5z��V=u���a����?���?I��?�|�.O�l�7)�ys�Y�Bq�ayGHʾ;)H�cf�ޟP��
�M��B�>���,��SW�J�J�� #��U�Q���?��\��M;�Oؕ1"�(��K?��^'�QRD���y�%�|�'f��'��'�b�'��S�KŨ��
�bE�b��Yf�I�޴�������?����䧵?) ��y7�B9b^f���<B58-2�#G�9���'�ɧ�OG��d�i��āt��0SG�;C�%k	;�yR�3~VM������4���ĝ�p+�I�l��7i*)[���@���D�OB�$�Oh˓\��,4�r�'��哏�B%����8&+N\��ȩa\�O��'���'#�'s�%`��0�މ�H3R����O����!Z/x���Q%�I/�?%L�O����U��e ؎AJ&�j�O���O��Oj�}���u�b���S�#-8�C�G%.�l9�v���Mz�,�	ҟP�4���yG��*%~�@w-��8�����i��yR�'W��'��;�i��ɶ7A0H4�OΪ��K�`��|`2�n�B�&�HA�	By�O���'3��'?�(_3}�(1�'�4�D�c�T�J��Ɉ�M��$ў�?I���?�K~�Ch�kSA�Db�I��%[�*���ɗV� ���t%�b>I����LE�p�,�9;���5�`�����#?�U�^��(����䓟�J%7��Ѫ�ͻe�rU���D>&���O��D�Ol�4�f˓T����	�S" 0`��k3,�eTJ�����yRzӒ�h��Oh��O���,9�)�i��:��he��F�x}zӠ{��[p%zs����>��=� l@P��A]f�x����*�@�@4>O���OR���OR�$�O��?U9�.��o�Z�kʗ�'� �e�՟�����Hڴ/<h�*O>1nZN�ɇ_��<���6b����)2�z]$���ɟ�1%���mZK~��ס1ސ�dK���Z����!�$h���i?L>q(O�	�O����O�+ש��-mƨ+�Ʈ9�v���c�O���<A#�i_,����'?��'9��u�<i*g�܌@��-O+ˌ�&*�I���d�)Z��=:��	:С��gS֭	�,5��V�Y4�Ms�O�I��~�|"�_�W�m��(V
Q+S��S��'�'{���T�D�ݴ6�Ũ�af���w�ѿ;\h������$��i�?�wY�l��ԅ	�h�.8~Y����ob����ٟ�2%�ݦM�u7�V.�����Hy���/uz�H��ݹ	���7�6�ybW��������џ��	��ؗO�lHk�+�C��9��IЂK��yYS�o�Q�r��O>�$�OT���D���睗I�B �`�M�%�Q$�EM�x�	���%�b>E�WΦϓV��H7 �Eo.Q���o����t����f��X&�|�'�2�'p�ѱ��H�vP�X	�!^>� 7�'�R�'��W�Pcش"���P��?���N��!���ʂ]�VP���(�,����°>����?qL>�`k 4v� ��l
�Yf	�a~b�E�����Β���O����	��ֳE
���Q�O�|�\�Зg�	6�"�'|r�'Pb���#��c�lX9f["v� �"�dA��k�4�|e[��?�7�i��O����)E@3c�
��� {��D�O$�$�O�#n}���A�E�Pf��h�C�L&��!���:_��9s��\�����4����O��d�O��D�T�����o����W�-o�:ʓ=����	5*���'�2���'ܸ�*RkX�my�uSu�8"��ų3��>�������O|r�8 �UE"@�pg@�U92�An+H4Z1��V���t'�����H�{y-��B�~E��cw��@�����'��'�O��ɘ�MS��G�?Y�ʚ�l�x<��¤P_����?Y�i�O���'��'j�f�ahY@��Ǉo=|�$.��h�D�մit�	��2��q�O�$?��](q�����Y
�M��#���ݟ�������	ݟ0�IE��}��Q� �̤�����b#=0t���?��tg���.�剘�MSO>yq#W�$h�!�P�تuj�{qiG����?y��|b�B���M��O\ܸ?D^�u��&���m�Q#	�eٜ�[�'��'O�i>���՟���<r�J k�NT5pt�0b���v�������4�'�N7��9D$��D�O ��|R6�ً\ˀLs�MH�dI��#�-�g~g�>!��?�M>�OE�B�oϷ:Ȅ�� �S�AOHi"qd�<t���K�N����4����v�b�O�\뀄N `wX�ʧ�� �.}�«�O���O����O1���	���h��;�T��ܿ/�l�$)�+z蠳3]��sش��'���?yg�R�Hސ���,e�e��h��?��H���۴��� 䘠0��G�"�`8�oĔJ͜�L�/�y�X�0������I������(�O��9s�_4}6<hY�(k"��Ovӌ�˴��O����OP�����K���ݿ��h1ȕp���E�(�Z}�	�8$�b>�!�	���̓	�FI9enF�x�й9t���\�d�ΓR������O.��M>)/O��O��S�PX�����ud�r���O���O��$�<���i�Mq��'���'Ͱ�B  p���낯ˌ(��� `��Z}�'G�O�S��G�D��D
U
Za�������-$����B[p�/%��B�".��M_�c��jxy@�	�ܟ������˟�E��'5L���۪��	P� L�S(ܐ��':(7�ޖ����O� lO�Ӽ�4hچ��}ࠊB7 �J����<���?��O�(�ݴ��dȷ2�h��O�Z��`��lk���լVc?���`�|�\����ޟ��������⟼7Q"4U(e�E�̼�I�Bny� }��5���Ot�D�O��?Wr}�I���%&��Q�2�Ӂ-���?I����S�'}�*J� ��}qLIB1$�~ȑ3$h���M��O�PFN� �~��|�X�[���	wG���j� �a�V��h������Iߟ�@ybn�J cK�O"�Q�)
�z�Ҕ1�!G�O�ni3�J�OD�lX��.(�I���	���/q�@͓g�8�`5���U��DnO~�,R2`�`����'��k��U��
43���lw���L�<q��?����?!��?y��dO�(b0\����M�J��L�T��'VR�}��Y��:� ���æ&�l0���B��e0R!�y���u�^F�	��i>��E�ͦ��ug��:0��M��	�=��5��M-����'��&���'���'F��'/��pA����d��J2,EHHF�'6�]�Xp�4NO
H���?1����)�.
0P���l��Eb����	����O"�D%��?aJ�B��r`�Snʋ8l�mSb���dqT��U,�-=������{�|��|%<P�bN�]�Y�f��'i�r�'b�'���R��c�4(}��8�/E�$d�ȊM�st����ǎ�?A�Qћ���t}�'�V�:UV�R���Y�BƔ:�̬���'A��V#L�������gx���~� x8�@�Vqr)"�	űPh)�9O�ʓ�?����?���?9����)H9m��ʲf@�!��%����>�$�nZ�\� �����P�S�h+���#CAG�QX���%��u�ҭpu�6�?���Ş2����4�y���A��1pFHQ�<p�G�א�ybigk����%~��'o�i>��I"W��sFO׃n��BeA s�y�	�`���� �'�7�} �d�O$���T�Z��Q�
H��+�4�Li�O����O�O꡺5�"p���_X������n+x�g4��n/�g�����֭8oB��vCn�A��ҟ����T��蟐E���'q�-K���5}�H�Q�V�@.<X*��'�6-U�]0����O�o�B�Ӽ;2f�9j�f]؂b>;�)���<�����䀨N�6M/?�c��Y2��ɕ96�N4�B,X���Uk
N�'��1)I>A,OH���O��d�O2���O`5�h�֩��� �b�C&ļ<��i���T[����{��a�x�d̔�6I�0CXi�P�D��n�Ş<�$��o׀g��ra��f����Y�{�|}:,O�)+dG.�?���9���<�ͽ/#-3���>H�1� L��?���?a��?�'������x�����eA�)A�Np"bH˯Mn�d�T�4��'�듏?���?���_��+s���9���ZA틉h4^���4��D�5&�������O]wG@�-���Q�A�(�6������y��'��'C��'���M6?4�q �R�>�9�x	��D�O���XȦ}��
a>!��/�McN>q���+�Z���y"=Y���:�䓴?Y��|��e���M�O^m���Z�n+���dm�9*��	q�1��'�'��i>�I��Ic�
��p
�+.��t1T�F<�P�	֟ؖ'~�6Gr���D�O��ĥ|�R�6^�"oH4�$�PT�f~��>Q������Ud<��i���� �!B�Xe��#�
�Q@!�<�'/(N������F�4���Z��ȍ��%[>������?���?9�Ş���[�=y��3c�&�RBI�z�ٳ�Ǵt0�(��̟$��4��'v$듩?����v���9��6?�l �'ר�9��i��ɿh�����OGPH�'�t�F5.Rz��g��8��'i�	ߟ��I��t�I؟ �I{���1x��UŘ'�<���_�H���$��YP��'�2����'��7=���3UG�2*�z��#)ʵe�v��O���7��i�$}j7mi�PFB�s���shP4�!�k��9�J��=���'�d�<���?1��4��y����+:lJ�.���?���?�����y�GEVȟ@��䟘9�I��7?�H�M��X�ؑ��U[��M`���H��z�	#D2—�3猏_�����%:?!���u��#үJŞs���K��?��F�"��t���B�i\H��4Η��?���?I��?	��9�.QU��tIcB�(~BuX/^?��`s�\����<AW�i�O�N����� �#1�4'��`.�d�O��$�ON���%h���E&����)S_~E�F�M9&"HI��0�O.��|Z��?��?i�,	�U��
G<dV����R�Yl�	p(O6ql��Y� ��	��Ir�Sd��V5mQ,ep!J��[;&P�f����$�O���"��)�4��<aa�y��v��Z���a�G���˓H����f�OX�JM>�.O��a�Z�N'0���B�A��4+!��O����O�$�O�)�<�b�iь�D�'`L@ѡ
̔^-
Tj7�^�w��IC�'��6�%��)��d�O~���OJ<:�C�?rU���0�H�U5�����X(^~7-9?�C
Ғ��G����uTm�!3.Г��5��(ו8���O����OB���O��7���e�o�w&܁JU�E�����Ɵ��	��MC�o_1��$����'��ےm �R���Z\`�3�f�~�I͟��i>%zA���)�'���K"wj�(�qn�bDr�G�R/X�F-�����4�
���O����%^O� C�&���o%~����O�hޛV �9'F�ܟ�O���cu��`���	��i�h=��O���'�B�'?ɧ�	M�u�h s�A\d�����H�\���(&����d6??ͧ1��T�	G܍
����IW.�'�)ɞ������	����)�ny��x�L����]�m�mJD!���8QtJ�5`N�˓vE���DQ}"�'��HhR��JB�,��MZ�}۲)���'�2�h��v��pkׅR�/Hq�L9@QM��)����	۱T��y@g1O�ʓ�?����?9��?����I�'-0��bH� ��0�"���=��Qo�ŕ'V��I���]

�$`A3�̜sm ���f�}�$�	Ο�%�b>�f��ƦQϓUXJ��w�υD�
�!�!ZP@�e�z�\$ΰ��&�����'C^��@g$K�J,�`C�'�6����'NR�'B_�tH۴۸dx���?	��|H�
u#��~�V��v�
�?�Xm�� �>	���?�N>�DѾ4�Js�}�@�$�z~��\6����'Ƞ��O���I�;B��V��`  3���0��0C"�'A��'g��s�e`�kY+O���:І�ج�֬Iş��43J�S��?1Ӿi��O���dI�/Ǭ+ L��Œ�QM��O����O�A��e�R��h������ T�z���7�P�1Sf��8@�J�d5�$�<ͧ�?���?����?Ag$��J<���"�H�0�V3��$��т�GF���Iğl&?�j	��p�d0CKV�r��������O ���OܒO1�H�i�Ê'��<�e5|� UQ��#�$6�)?	T�\�L�R�IX��gy"�_�qf�2шݒ�t(7J�,]���'��'��O*剤�MC��.�?1a	�
j�DW@VF\����%��<9��i��O0��'��'$�%�y�g�D�[%*]�eIH=y��{ói~�	%!��=ٰ�O Ĺ'?i�ݦc@ܽ�V�ҵ%������n����������I�X�Iq��P&:Y�櫘��n�Q��< �Ĺ���?	��8ϛ������D�'R
7M.��҄�hM�#b��J	�)�,�= �O��$�O�)�,V#�7�2?�4��JY*(�UM&@o"��l�)Jv�� ��O�d
L>	,O�	�O��D�O�i�B�jn )�b�@�����O�� 9����d�O.�'i䠍�'�G�{��[so��\��'�N듌?�����S��P.%��0Y��ހ �ΠI���:vC
�SR��9N��%��O�i�?�3��L:c�(U��� � �j���2����O�d�O����<�1�i�r`Q��Ɣ|�8��˝�4�v|JG�ɀ��I��M�b˽>!�� �%I;;�`��ڽ�yS���?�����M[�O�D9�.����O"pP��ҬߪW8L���㳉Z�<�.O2���O����O"��Od�'�"͙�H�!�����9i0yC�i3j�:��'u��'9�Z�lzށ@%�9o�zͱ`��GJb]�Q' ����I\�)�Q�:ynZ�<��MK�\�ZaZ��Y�x}��BÌ��<ٕ�&���$O��䓟��O�D���� �њ+4J �r�	�I��D�Ol���O�ʓ�戙�b�'��L� h�����Ԑ�Xڅ� .o��O��';���8E�F]*��X�kN���U̇H���"��ۂ�%3��$?����'6����Y1:��gZ��j1�S����	Ο�	���IG�O^2�ۀ|꼣(�,���1��+���g�X�q���O������m�?ͻ4���	Cqa�uV�3'>�ϓ�?��?iG��&�M��O�N]�9%0�)� qv"e0����pء"�ʙ�~���ZM>9/OT���O����O��d�O+L�?W����N�=��yqJ�<�·i���Д�'b�'��y�.Ĳ!RhE�&葋��8y%+�;N�@��?9���S�'jr�!�P�1�ؽR���>�@JBi�9�M�R���J��D,���<�4���������V��1��O��?)���?���?ͧ��Y��Jw����df�4��l)�̅�48D��4�����I۴��'���?a��?�2D�>mHH �$��h�2�XBL���ٴ��˔K�+�'��ORצJ�H�´8c/��RA�x@m��yb�'���'�B�'����ǟ9�� ��߸��	f���U�~��O��$Gæ�OOyH|�f�O����H�t\�xyu
&P��2�)��O��4�y���f�v�#xx#�K�N���ffV$1�:�s��-6���	v�[y�OS��'_ҋ�='1�X�oF�?�z��A�5\��'����MC0�Փ����O*�'6���x��R�^!HQ�!�$=UB(�'�@��?a����S��mΉ�9x@˝�HŊ���B���$�蝴��֐��#w���8������Yq���`� &�H��D�Oz�d�O.��)�<!��iz��r�5&�.T�6iW��#��.4��9�M���i�>���(=�ȷ蚂]^�	�F�bI$����?�(��M��O�-ʧ ָO�l��`լ̒��؉B�A��'��	���������I�d�	R��D�w��اC˗R~���BZ	J�6m3�r�d�OJ��(�9O�Loz�yK@  a,Q���(*�,��	��	w�)��!`m�hn�<A�왱o�\��R
�ck�!�S.��<�
П(����_�Ty�O��o�ZD�x��Nk��$���^���'R�'X�	�M��5�?���?)t�Q�<*���d
of��2�k���'Yx듌?����=��y�`�Z$:��u���!X��'u��ҋ�H�FC&�	U�~��'؀���S�����`]�x?<U���'	��'��'��>i���o~\��bB#8 ����GnX����M�%��?i��2:�F�4���Z��քTO��ʰ/�j���3O����O���V�+tB6�8?yc�P56it�)�}V�X���ǔ�c#,P;��O>!+O��O��d�Ol���O�����O���o��i;���<�Բix����'Ab�'���y��]N*-�) ��(��!@c���?���$���N��s�
�鎘[��Y�K� $��<y��	gg.}��'��&�h�'(x��%t �9��;(��y�'\��'�2��tT���ٴ-ּ���Z}������Pd~�k���%���ΓcK����R}��'��I-m�8�ӂV���Bb��o"!�������'5�����?�����t�w���j�G%y���%	�A*ظ�'z"�'���'���'��R  ��6���$x�bG�O����O\qm,��П xݴ��u!��3DF��1��9CR�%�NtO>���?ͧ���4��d]�3�� ������5q|X�A��S �8�E߬�~Ғ|�_������(y���z/��0ևM=xo<��%G�ԟ���Jyr�~�V�(c��OP��O�˧Q�ř4j?��d� Es|��'al��?����S��Ș�Tp�l��N5N�z�H����qJe��8��x@^��� f�B@k�I5����3��b�1SǄU�ag`��˟�I��D�)�uybd�vqv �0BZ�1��H
BFɺ�m�C��D�Oh�l�c��%)��ڟ�C��/�Ԁr��<AuK�ߟ��I�xR�oZ~�K�,5�����A���y�f����K��T[�j� jc�D�<)���?	��?���?a+�>���ϼ|��@I�ȚW���=�"�ןP�	��L&?U�ɝ�MϻBc�L�2A���)�bf�%���(��?9H>�|��N��M3�'IP ��J�!Y�:�:�U�S�`��'�X������9��|�Z��Sߟ�ht�s��Jq�
X�,��ɍ͟��	���	Uy�uӀ�x�C�O��D�O���"e­/���f	�`M��V&+�����d�O&��=��k�|X:v苇B-��bU`�<a�I�ZT�QJJy:�c>��'0�����|z�M�`�`��)�����8��̟���[�O}��wm� q��
Ri9�/�:B�#b�V�!R��O���æ��?ͻG�@腯+��l�6
%��H��?����?���,�M#�O�N/���I �}�N�S�᙭O_��%��
6��ؑM>�-Of�$�Ox���O���O���u�D$TM�F戡BI�sկ�<�°iB��'n��'�Oj��ΙL�2�z��7-�&	;ҍ]�o����?����S�'W�t�2��]�/X�e��@U� pt�4�M�U��2�&3|�#�D�<��cՓ78���bEE�\[����O��?9���?��?ͧ��ZĦ�`Y͟���,� *���m\�JE�"�Čɟ �4��'x��?9��?y"�$�\�ã��_����٠�J�Z�4��$Υi��?��}Z��wGT�q�)R�q1��'��Nޡ͓�?���?���?����O�fU�ė�.q���d���Z���	��M����|z��E����|��
�=�ŀ�A�� �T����ճ[��'5������P*pC�֝��Bh�4q� 1;�d�bF�)��W�:uG�'Ff�$�p�����'��'$�4@�j�,EF]"�)��K�t	��'��Q�`��4h�����?�����	�-� �ZGd�Dӂ�����,]i�	�����O���2��?��b�{��i�>z!W��*���b�<c����!$?ͧ(y���B���W�V�yE葪QZ��g�	� M�\���?���?1�S�'����q��L�3 H�1�7�W}� ��I�1�I��x�4��'F\��?���Ȝ~����֩�rޖ��˄2�?���Xup�*ܴ��d�%Kq�q�����Sd%�R���� K!a2��{y��'B�'�B�'�BR>	�l�d}	j�!�,t©�a�^�M�pC���?���?qJ~���j2��wX�y�a�'PG\�*ExN�|)��'�|���@�[/��9O~AY#�\
���фՖjВ�t5O `� މ�?�9���<�'�?���:� $��Vm�E���R��?I��?���DC�Y��	��d����t��oC�>�x��+ϰ0 �	Sh�g��`�I�(�?AM;q$ERS���@X�1X%An~���}^z�L�%k�OR~	��$""fH=S����ac�p����A�!G��'2�'4�Sٟ��v���0U��Ɯ;���6�_ȟ�[ٴA:��+O�\oy�Ӽ�D�=XB��B�I����,�<q���?i�H�ݴ����v�34��P�A��E�9Q��'�X�����䓅��O<��O<���O��$��
�b%��Nu�׮T�UѨ�{F����'v�R�'����d�'ٌ)�CB8h�)���<lh�8����D�O��D-��锗|�����Df�"��+ò:p�� t���&��sB�Oĝ
H>i*O��` eV0na����#�u�ب����O��$�O��d�O�	�<%�i�E@��'r��#��I�D��h�ߒS�J���'ؚ6M!��)����O���O�j'""F��gR1X�T{��ӟ;Q�7�7?Y�՞I����Z�S��I�F��@UlU�ta��'���@i���	C8�m#���.��F�ʃ"��	������M{d�D�c�T�O�Q8F��"m�j�($�ے K��d�:���O��4��,Q$njӼ�Ӻ�De[.��xX��Ѯ3�� ΍�{Ò����`-��O���OD�E!L*|,~ѡ ��ah�����d����Oğ�������O=�-���݉,$�0P��	�(d�\k�O���'���'�ɧ�	�9M�4¶&�_�8���ϪZ����nϕ]]�����<�'6Ux��כ��b�9Y�S�0v�Ю^�\ ���%(���{6�bd�v(�h��@F�"Q.����'E��j�⟐��Ob�䙙���T�Y�������^�d�O`�Rg�.�|��E�?��'� ���ON� �~A`@d��D��@�'��IQ����v��(��S>f]�L��ؽ�M3�탓�?����?	��Ăn��nd�7)�	�"�_��Y26��П@��\�)��,��o��<� ��b_'!VDJ�Mõ�^��W8O�u0���~b�|�S���'Bb�kq-�d)l8��TcWF4j�B[��I��B�'N��)�6ic�@f*�@��@��O���'�b�'B�'˼�ȡ�����w���
��O�=H�Xva�6m�`��5��D�O�좒$�a���.�2\��M�d"O��!%bX	h�`*�[:i��YA��O*�m�	$|u��؟�(�4���y.	Ė�Y'�ȉ�X$! ��yB�'���'������i��I;	P2�ӟP!7�J(8n�mL!j�З��'`�	x�'0y��[���J�M.�
�OJ	oZ��4���̟���|�'m
���ޤI��@[)Hpb%+�P�L�IןH&�b>QX�ǥu(: Yc��4)M�2@���,�oZ ��ĕ2�Lh`�'A�' �I�QT����� ��;���UrX�Iʟ�	����i>є'�Z6M�%	��ȇ�j��g��)i�>�dn��]������-�?��_�|���������VfS�z��IېK�vt%��Ŧ��'A.�ڡ"��?������w�詢��ӚQ��r��G�=∋�'YB�'�'�B�'��l�դ�&0[�,(�I6�U9�O�O^��O�im�7���˟�P�4��_Qt��`�Ϲ"d��OBsa6(�M>���?�'l+���۴��������5]�l��۶:�������9�����䓺���O����O��D<u�@y"���b�MeU�Nm����O�˓}���i�:[r�'�Z>ISȔ2$n�c�@W�.����u/.?A�R� ���� '��'P>��2G�
,d�99��	�a�z��T�y�ƈ�A�����4���#�k�̒O�e�¬�0>00%��� 8[Z�#��O���O�$�O1�8ʓA�f���u�~P�P%�?mΔ�!
�tv��P��'T�ky�T�S�O,�D�zP4��PCX�j�p�U�@z:���O�Qq�o�R�ӺKR��3��Ué<&�U��v؁Q�ʑ�Qh��<�(O���O����OZ���O
˧9�8�qNE2r>���߹\���ѺiֶY��'�B�'u��ybLv��.�c����eC�?@�[�F�e����O2�O1� �Ab��8+�\X@!�6jn\q�oJ�,<*牀N�1���'�$�<�')"<O~�s���3π@x��(b̩3$�'Y��'�"T�(�ܴ/�"�����?q�`�E�u��p@���Pe_`:@N>��X�I���	G�1y��Җ�ܯ_6��W��@z�_��\�F�A!�M���t��B?���|��n>X����4d�\4t�;���?����?���h��ŧx�GH«F��1���G1$�H���⦉"�h�����	�M{O>��Ӽ{�m��ޢq���$0gj�Qk��<����?��"6	��4��d̙:9@�:�OOYb-Z6eR Ej%*�VfQ`f�|Z�������I�����ɟ���+Ǆ�jqGS�_h tR6aWry�l�b�H �O���OB�����)��
R��X� �b��1���'��'jɧ�OK��&�� ��:$��!^�Q	H�D��	�<���B0I���I@�	ey�Ƴ�DL�T�R	D�ĠB�ۦ7p��'g��'��O�剶�M�B��?�sd�%E[�Yj����d�R�x5c��?���i/ɧ�th�>I���?��c1f܈�����-��(0nڪ2[f �4����D��͠�'3������nZ6e%�u"0���`F��'@K$]��$�O�$�O��$�O���!�Ӆu��Y�HΠ�P��	�b���F�O����O�,mZ X[��ݟ���4��;��E`�$��Ir���Tk*�K>q���?ͧr�D���4���&A�( nL�o���1�O�GՄL"C��~b�|�Q��Iן��	Ο��R�Ȩ/�8Bk�l:��q�����	ky�t�v`�p��O^���O��'#8>��PC]'T��[���At����?��_�����P$��'	,����L�`Ә�4����u
�L^�B���J.O��V��~�|b�Dd�QcAH�K������Q�b�'���'���^��j۴!,��"��j�����Y-M��������?��&���dF{}2�'~�!�J@l12��g�~��5s��'�ҎM�	����p�tq�j��vzy�eb3���8�ąj�1O$˓�?���?	��?1����IJ1N�\��� �_��]]��
�i& �q�'��'S�qmzޕ�v`Аs>��C+_��d)2��X����X�)擟7���o�<"܂6��h�֊��'f.�ʡNO�<aS�j���	N��uy�O�����,2 *5j�>n��@z���"IB�'���'I���M��k_��?Q���?�S&�8��ybDN�6 y�P,��䓥?C\���	�$%�dSe�&N��$�Z�Vʥ�L$?9�I5 ha��4_��OB���?��p��\ĉ�D��!H;���?����?��h��5~���A+Q� �3�d�2��]ڦ9���ş,�	��McO>���p�:Dp4!��۰k.K��C�<���?	�5��E�4�����K�~ �$ݣEИ!QS��/aALT�r���������OF�D�O��d�O��$�(i����5�h�	��	+�r˓1!�F��UK��'�"��$�'�L�e�Q�+����rE�Tc�`���>����?	K>�|Bg��j�? "��׭�
ǈ�Qʑ�j�ε�֮}ӂ��'�TT�W��u?aO>�/On�C�ΐ��E���&�X��� �O����O����O�	�<AĴim��R0�'g�����)'G�!e���:�:�i��'0^6�(�4����'��'e���1Y��3)Ts�:��cR>K��0�C�i����I�,} ��OJ�l'?5��9"�&���ӏh�P��FՔ&��Iٟ\�I������4��_�'w�Ka���!�!��2ľR/O:�Ʀ��7�p>��	��MK>�J�Z&��nG�Jm;� ���?9��|:g&5�M�O��$B�˕���ֵ ��
�F�F����O��yJ>�*O��D�O��d�OFU�r�ٗ8�p�����t�8��a*�O����<y��iQ<x1��'��'�Ӫ�*xӅ���)�*� � �2.�I��<��O��d�O��O��(a�p��`��"ii�A
����O�܍vW�D���o���4�D ��'��'1��IB��
�T9��?i���c�'V�'u����O7��M��K�
\�%9 +[�B�t�U䞤p6F�����?�w�i��'�Ȣ>	�h��{"&PtR���@W:�B]����?��$�%�MK�O��	ֆ_����S����4G0��ذ#�&W��3�
b�T�'���'���'q2�'��өf���ʑ� ��`�&����4#/�T*O\��4�i�O�4mz��$/Tl�r��]�v�P �៰��o�)�"���n��<��/���t���J�� v��<���үD�$��������Ov����Alj�p%	$80��9E�U7a�����O<�$�O��3�f�C����'nR�[�'��K���6�����.��O���'G��'��';z%��+�=I��`q���%l\�q�O��� �W�An�7M�\�*\��D�O�)��ꓵ?�@|��a�g�$����O����O��d�O:�}Z����x��+u�`��D��⡙�6����T��'�7m �iީ��KS�O�48����4�8(j@Ep����㟸��;S��m�A~�&�&�@��("�s(M�r�� �gL�, �2}�H>�/O2�$�Ox��O2�d�O�ຠˏ�045��I�6g����"�<Iv�i��<cu�'3"�'���y���� ?|���DE"Cd���?����S�'k��au �o[�M����<?R�]�l�1�M�rY�����
�[rvM���΁�Si�v�e�Փ0}h8�$(�H<)QG��t�`�X��!t�i<Q�Byg�Y �-�|kҜh�A[1Ԭ8`�eY�mBc�)bS��!��"�h�x`7�	M���&Wΰ�ɣ"ƉM:������(ArڑH��Y�F����:W������B���1��F�P3�����wD��G�m��4�v�$k�8	�w��v�D P� D�Xͤ����,h$ ��C�>S!�T6#��fJ�$�4E9���4�����L�WھHR��:���'T�9�<��GVq4b�0�aZC$�6��<�����?���!�ڀc��Y��R�
��@脬����M��<��_������ ��m~��
?*��쟬i�AżTbla��,�5�,��C2�M������?����U�{R�� �
�c�X�3�������MK���?��O$@+���~����?!�'Q��!eD�p�Q� ,��CX��	Ğx��'���*`;b�|"؟LY���B8�M�V�Àv�P=�u�i��	�<n`n���h�I៤�ӿ����ܵ ��� ���c�n�< :d�9!�ie�'�
ۍ��!�ӕ%0���H�x�±:t&�h�l��#?�6��O���O �i�Q}bV�x��V�zY�Y:4��2bj���-׾�M�� #��'v��dI=~�|x��f�J�TlyV	�xuL�m�؟��ʟ@�P�����D�<����~rU*q��D�U�+�Jez7��0�M�O>ك��e��O\��'��Jܓ6.�A5(Ox�����:S��7��Of��}}Z���	}�i�Ak���<s�rp2��Z�N�|��a�>S�LL��?a���?)�O.��U�̅�A
G�W�&���j�� \������O|�OR���Oz� �9$4�	���h��s�+C�;pL�O����O��d#?��$W<��4u�(қ*zh	[�ͱ^��}�q�i%�x&�P��\*k�>aE�W1}�`]З�I����i}�'"��'����Ox���O�򫘴a<
!��G�%V+*�s��*7��O��O����O�0�P�%�	 N��(�&�ҟA"��H�4�:6��O��(?aP������O���l���j�k�THx�,��mcz51�o�	ğ��I�5�0��?�O֖��J�)�l�?!¸qݴ��d)	 �6��Ob�$�Ot�	�P}Zc��d9�ʋ�olz��K�15D��4�?����	�b�i� 2�z�H�d�&%�Z`�#$��'�H���'p��'��m�>�+O�$sG��XU���#���F��Ȧ=��Wj����O���F�fy�"�dW\���"'���#��6��O����O�$�d$K]�?�D��l�3e4Ҍ���j0p���Gm����&�D�Z��'l�'D�	:���DF�I#��CV��9�6�O$iYX�?�9�d�:;��9��#����,�*�$����~yb�'%��'��ӞA�=9�O��}K��\�_��KÔx"�'���|2Z��ݰL��i�k�n(-[ES�bk(6��O6��?Q���?�̟^�#6�b>=Ѐh̔+bQ�1hP�.-��ծ�>I���?qI>A)O�i�OJ�a�f��%2tː�����'��'f�V�|���A<�ħ� R՘@)�	y�`R�]#-sP�iS_�l��gy�O�r�~�逜z��4���̞	�������]��ҟ��'&�i��..�I�O�����q�I���hIr��;3ތs��x�P�����x$?�i�I� ,��O���H`B�L�\�S5�rӂ��a�вiG(�'�?!�'|.�Iڑ2���08`z����6ͯ<����?�֕�4��ܴ`�Q���-X,�qcݻp�>um�k��i��֟��I�(��Fyʟ�QJ���ELNY+"�D%�U��U}�%���O>ig�R�@"A���1>������E��Mk��?y�O��� *O��w����>~v�� �+4] p��>U�DDxR�"���d��Rl��(FH� ���@" �:Ȧ�o����CE�@y�L�~
�b�Ǿt@�(ɗ�9}2Ś�ps�Oz� ����	���	q���L�<ʚ`�� �^�u�%ʓy�V���x�'�"�|[��]3��Q�@���CF	���7��O:�O����<�
�\��O~��Y�)Y���Qփ���H��4�?9���'P��;H`ӪĲR/�#?�F�{�
�)�ظ��xr�'P��՟x�fo�S���'@�Ś3�ț��	b6e^���Moӄ�|��Py�����ēr^4숔ŔK����d&`�n�՟З'b�/�ޟ��	�?טm	�h"Po,ڠ���f��O��ĥ<�7��~��uw��(>yu�vk��aY�MyW�E>����Ob ��OZ��O���*�ӺSBLC�c�R1Y��/=�� 
�m�	jy¯Q/�O�Oj��p Yi���Q����7��!#�4.� +�i 2�'�"�O-�O�iNC��J�@���PAY�M�L7�OZ��OʒO�s�h��6k36�
�Yai�E��,�׉�Ɵ��Iڟ��ɒc�Z�{K<����&�X���̑��HⓍ�abĠm��<&�8A���$�O>��OZ�p���dA+2���mx�(S즕���r	�Q�K<��\�'�b��� ��$�矹)� �ÇrO|���<���?�����D��zݴ�i��(�*�B��Cp�D��M�]}�Q���ILy��'Y��'�j=� �ТF�V�Pp�#T�X��4�R�y�_�h�����Iy�.]�Kk.�S�g�6�#�Jݖs֐!(�E6-�R6��<�����O^���O�!�r3Ohm�Lٌ�M�f� � MP!O�ۦ-���P��򟬗'̹x3�~��3��=1���b	#� ��Lۦ��	PyR�'db�'MD�8�'���Ƙ�1̞8���@�C;N���m�П���Vy���o��맩?����c�,�Ҍ�oʩY�H=��C.w������I՟���p�X�'�ޟ�dY��WT���`T*W����iJ�I�g�P���4�?	���?I�'O��i�E@�F��LyiUm �l�E;�l�����OP���?O���<���TjDb<6!�\�� Ѝ�`_�V�ߓ/46m�O�$�O��ZF}BP��A$�-�*z�(��m�d�I���MC���<I�����6�ן�pE҈[����nw�I�ӭ��M���?)�]��E_���'�2�O���� 82��6O�&g=�Yd�i>W�
%q��'�?���?�b��8%���!��� 
P(� ;��'�ްXRM�>A*O��ĸ<I��K)��p|0�'kH/YҦ�g�c}��I?�yb�'Z�'�2�'W�I,a��Z�E�rX`s
Տb� ���"T�/��	Yy"�'L�Iٟ��̟�1)�.wH�|h��J�O�0j���4���?����?!�����y��ͧV{�bCU�$�A"bC�!K���m�ry"�'��������j4�t�0;���${B6U�"
;0;l��#�:�M���?���?Q/OZ�x���X�$��5�/
d�J���(ɼaC�dZ�M�����$�O���OJ�S�1O��D���teE>7�θ��gc2�D'g���d�O�˓zL���R?a��؟��ӑ�\0�G�.5�L��b�Ѡ :~Y��Ot�$�O�����|Γ���CR�  �r$�(5�@�:7�N	�M�.OD|������	������?5:�O�n�~Ͼ9Y��ŭ+h����l*���'�B�մ�y"Q���	UܧK��;֊��qt$�i��3#�(l�L�X)J�4�?���?��'9���My2������ä�D#�Рs�OX5wh�6mH�����O�˓��OQ"H�i��i����CҲ�
� ��D1t6M�O�d�O�u��(YN}�P����v?	�iđ춑	 !8��a�H���vy����yʟ����O��Dđ�@�!r��3�C�D�Rx��lZ蟸ʇ@
���<y������Ok,	X 0%H����P��2��]�W/���'���`�'���'�B�'��Z���#ɕ�Uk����4F�{#̕:�^YC�}��'��'���'ښ ɖ�F��������xF�Qr�ျm��X��	˟(��by�R����q���(s�ϐT3�U "ݘO��$&���O��D��OY�Z�#ӊ��n
7��49�.��]�'��'��^�L�s�R&�ħ`Ǆ܀�,�$^WP��A�:%��! �i1Қ|R�'0B˦Z?r�>a���6y&�����%���IFbͦ�I��P�'�p��*�I�O����La�CY�8�b�H��I&�X���ȓ��c��%����/��u������m C��);�uoZwyRH�Dz7mYw���'����7?� L!�ւ��	"l�{'�3E���s�i�"�',��'��'�q��0X�`?
���yvd? 81d�i���7��.�$�O���V��>a�  �1Pz�᐀��N�"lb���:������y��|"�i�O�@�FD)}H.l�5��'��a��ߦ���ş��	�M|���K<����?��'��	'�(a�-*���?����4��U��[U����'�r�'r�u1%/ˌQ5Qj�l�5I��5{�m�����?llh�%���	���$�֘�zĄZ��ŉO�ʐ��I6 ��EO������O����O>�IґU� j���FT�q�|y�]�-V�O�D)�D�O��J;r�K§��{:�,!�-	�YP�!���O@��O˓H��lhP1��5x�ӫD�\�Р��\d��HP_�,��V�'Z�	ӟD���8UÀ	2�Ş7�-3���&����O`���O4�-%⤘Ė�N��[
�VA� r4��iC+G�b��6M#ړ����O��'��h�V��;�x0"`�(E�,cߴ�?����?�5u�����?�(O��I4f%�a�F��v�����M \'�d�I~y����O�.�8	����I%�ݸD��{6Q����Ȇ��Mk'\?}�I�?i��O�ub�	��R��,���4Ƴ��'���p��D៉'�����I'�`�c&��@|��ݴS��<����?Q(ON���<q(O���)��-jĐG,�	jH�צe}r�Y��O1���$��3�0� �@J' ظ�@�,�k��%n��L��������ē�?���~����*Cfѩ`�����&@���'����yr�'���'�n�H�ߞ<�@Ƌ�,��HGbӰ�dR(W|'�h����P%��X�\����A�.DiF�
�dR� �	�<����?�����	T�fؚ�@���
V�K;Dz����mYm��?�N>���?�dQ|�q�&&S7��A� mހ9v��<���?��� �6�ͧ?��j�'7�8a�o�5ǌ�'���	x�֟������'�ؕ�R�H�J4����n�;\�pM�'�'/�[�X	���%�ħv��P@Т��4΁2$ƞ0�,]�r�ii��|�'h�L٫��'��e�4)�BfN����w����4�?A����dE$(��t&>����?%���e���c+K�~��0��B����?i��h��Fx���҃� oG�" ��.#�v�*rZ�|��e�t��Iٟ��������ݟ��'>�8��A�oϖ\�uH݋G~@nZǟl�'��Í��t�]�#L�	�@��LE�`p��[�M��@3��&�'b�'���2��O����6В�9���@@:JT\؟���m�la�U����3)�<g� ۴�?a��?�eH�]c�O��d���aY�@s2T��hγm�؁�+lO`���O��²v�z��i�|�Ah�F�$$�(mZΟ��'�ς���?�������"~=��+s� �*V�UhĄMW}����'���'G�I۟��UK�+Qz���� )c
��S��^�f��I蟼���� �Ik����$��T��� f��> �m���Y�Z���oZ�k;���?���?�+O�XjG�|�2�կ�Z��d�#�"��W@�f}��'q"�|��'pb��$�3#�H#�	�98�=���\X��Iޟ\�IߟĖ'T��1�� �i�FHP���N�:�� �kN��,nZџ�%�\�	џ�!Q�:����#����Y��)ò�U�NI�6m�O���<١�x���(���?!X��N�v*�8ҩC1@(`��f۽��D�O��d�O���5OL�ĸ<��O�.���@�8�|�pc�Ъ[�n�[ڴ���*��nZ��������������Ԡ��#7�ҐG2��U�7�i�b�'MPh�'��]�d�}:��!:*֕y"f.3��y�ϙǦ��e�M����?y���UV���'�H6)\�7��F@˺BI�Bcw�^���1O ��<�����'�½� �
)����K@�fmtӠ�D�O���D�L�\��')�џ��~��(��7l�Ti�Va�<n�ן��'�j�"�����O����O�(�3E��2�k!�I#�<���ަm�I,wF�ҩO8��?9-O:��ƪm��%=\e3q�A�Xq�V��#0�~���'Z�[�G�(�J��J?�ء����D�����/��Pǭ>D�D��A�Z����6DpޅI6�2��h��@H;5(~A#�'��l	#�K�
%�xQ���0�`�����\�C(M������h5r�A@*� 	��1sg� "��1!��2�z�1�^.I\�;!��<I��Q�*�1b]l2%CӲNr}3��Y�
m��D�#+����c+y�p�p��,V4��S����{���£�7_�l���C�(2�����8�	� Z�B¸4q����Ȫo���+�
Q::-�i�+,��x0�,W��|�f��r�Q��XTLA0�h��P4a�0�o��)����S���5{��0�*�j�L�2PV�"fʪ�?����O:Y{��X;L<��v�e��j�'��B�Y�"8�u�4�V�d�q�혰�0>!3�x�BZ �@�yedF�\���KӦ���y�h�zGf든?+�L{���O����O:lqv��^p�W푘?eZ `���PC���.�i����`�۟�'���?y�F�}�t�YF����`Aw���G=ځ����RBX�s�,DC������ 
�CG�PT4�@��|I��Pѩ��uH���O��S��Q�s�H}S����?�T5p��,8C�ɳ�l�a!��!R�x�,{�Q��J���?��Ԫܯz<P|��&X5���Rv�����"uF��3�������	�u��'����#L�ر5(Z�W��[0NY �~�!�0u��<:�)�A������^M��O;W�R�F��d�R)��ƚ��LI�㉕�P���������À�ϸ�I�d��d�O\�=A)OvI*��P�?��g@�i�Xi�"O��[��ɧ	N��6E�1{.�@�(�E���ɷ<��O�+h�Ś�uڄa��L ���q��T�+@��'F��'����'�b2�PP�gfG�;?`y-A#S��Eu��
x����(�Є{&2<O��!
��8�;���&�A� l�Nx]S�ַn�^�`��3<OvQS�'��U?lk�h�7/
z	,6'b ��=���d�!��qw&"|�L1a
��`!�D�.oD��`.V߲�iV*��88�t}\�Pb������Od�'����P�}�\t��-�A�$v�*���O@��'P���l߶5b�i��Y��'m>@@ҷ���DNdb���`��uDy��Q�YQ���ԁh9x!���'vp��D���<mX3��Z�QDyҁ�?	���OK�u#0\������IV�ت�'0�R���<�"2��4.{�qE�R1�0>!��x�AߘW%��0/F�ؙt�9�y�����`7��O��$�|JHW�?���?�2�U�X�H	j�o��NใW�E�#���������	��X���b�8Z��̱�ؒ [jq���a����"m0�$j���0$��ؕ�U��� ��'1O?��Q��| A���L[�ī �!��E�FV�sUL��&�Ό�G�F�\�� S���?PE"G8m8 �	�����BQԟ4��&!��@0�ڟ$�Iß(��3�u7��y�� �X�ǂ�h���3���~B$_&��>���8D�l�MծcH��OUU?��Ix��{`�PԊ�\X%�`�Zߤ�ɡT���8|O8����^���1�]E�8���"OLmy�K̉`S��WB�NmH"i�����х���͑&�Ռ�Dpdh�?d���Y��ܟ��Iן��I�m~����؟�̧G���	ޟ��6�̀S��"���,uڜ �=�O>h0P��c�)�47/�-hP�C�G<�+	<�O��'�'����=4��T�ۜ{��P$��3�y���:��A7�-����ӏ�,�yR ��GF(�y�M�Z���U�y�k=��)��R۴�?������!qHJ9U���M��#�X�~٨���O����O���Fh�O^c��'F�BE��3i=�����Ƚq�L8GyR+�(��d�"���o�l�G�?{8b,x �	�"l�$/ڧ5�,��ɅP�ht��Z%��ȓ4VqIAk�h� ]�Љ܁T��l��	:�ēyH��3�^�Ha��c������s��1��iG��'��S�h/���̟L���(�L���ߨI(�5B����'��X� J�柈�<��OV	��	�cy�88���j�ICdU��V"<E��V�9� �ۮH��=SE�k��ِ��?ٌy���'άXą�;t�#6�,ҪTX�'�p��!�۽	/+�؞w�R��U�*�`L���w�<�s�G�55�=��\$"vM���?�4$��\+&D����?���?	���|�4���iΥP3D�J +Yjjb��O�9�b�'�~EҒ.ҹ���Y	ڈUL��
�'����X���S�.rt"���&���P��{������2t�� ���0$�E�Æ1D�p �ݏG3*IBӉK)[�Pv����HO>�Ӫ���M;��Qr-�Ȁ-088��m�>�?����?Q�u�����?	�Ob������?f�4l�&�	��B��q�W�B8�|j�g�<�q"�<OVhi0�g��D`��r8��Z��Oj��U�=���,����`0^�T�O���OX��'T�V�I�ˍm
�)��" {B��ȓ@������/�̅���Ѿ�x�C#�Ihyrn'l�D7��O���|�T�ˣhu�Ű#!��uc��M�3�R=���?�N�$��혧�˔b��8H@��<h��@��-Y�W�Q���	'�'Zv��$	y����.:>v�GyR��8�?Ɍ�� ���c�ʶ:���pԣ!OG�( �"O�\�Sǘ4�x��K:k1Nca�'�,O&�p1�))�8P$�` 3#"O$8`�
e	�d��K��@�`�"OL%zr�4Ǝ�g+Z��a""O5S ^����3�J�&w�v�q�"O�X�%�c5����@�IƼ"�"Odm�B!;��0	dc�2���"O���c��i���K����LPw"O�$���Z��~�1��Q�Zl�1kF"O20	�@�"}f P��٬qY�M˲*O�T��MΖBE�h����(Tx��'���c0A!�~�˶I�3�:z�'�j=X�-�hk�ݰ��O���0�'B�;@��?"Xpy�b� p���
�'��\��)M�*~�u�U��@�'"�MI �G<3$���TB��.9��'�F,xe+=Q.�8)�@�Hd�	B	�'�ة� �	7G��Ԉ��)@�Tx�'� pZ��ӎ)��<�7 �0n�ɳ�'�h�P��X�q�.��� Yf�p��'��=����]|���jإ{CpK�'����"�6D��P�W/��nѼ�	�'9����$W5��J�CO���'���@�F2?�d�YqFN�3�����'E�����*\��1��i�*3 UX�'�z XY/F:�ks�Оv+���'�Ψk����i�y ,G�o�д�
�'s$� m@�^��T���]�f=b�3�'�6���&ǂ4����(�dK̑�'}�
PJ\��1�XX�-��'~��35L�"����Tb�%NΨQ�'��Eɑ��L��	h�EE��*�'�	�Պ�>!�bt���8G,�=(�'�<�֋վ,"��"���6I�' :p���-[۠x��Ԡ� ��'zX\i�'TFCT����i�	�'�B�	�DӮ{� ��� E{���k�'s�%:Sϗ
M��9�i�;d)�1�'a|�1e]�:r�K���j��݊
�'F��p2OzzS�Lٹct����'���FG/@�<b�D�?[S�u��'����4�*\���b%J��K�µ2�'�\	�%	ڿf;䐂䧘�+ �p,O����
�]��ܒ�d��[B.� }�P�b`.�O@�"��xr��1tZ�%�.�w��K��-D��fbS��$�`�@_���@�,��<��bRg�O9�@�`���ք8+ԅ.�ԭC
�'�ԁi�/b��a��fM( qQO��2p`����O�q��9s&H��<��s"Op���C�!7`(�G��'��\���O���C�,<
�{R-4,Cn9@L�=8$x;�&��p>�`�A�L�u�	�4p9P�c��>L��M�?X-�C�	�I@4Z�']�0qW ۉ}�"�<�W+�MHF��dۥ_2��`�ѝ)��Qs���"�y��0r� �D�Q"۫�J�;4H�)��'H$F1O?����g��p7+߭o�\`1Q��c!��U59zJ�*'��5�2�)��P"U�~���Ó@����I ot��(���������\4s)���]6w!�$���8���V�z���Q�ى>>.�>�ci���H���X�nؕR��܊T�,^�:�y��I�3���4nٗ�(�V��ǇM�iI:ŀ��\�O�681�O�mR)'�)ڧ}�t�����;:�,�s H�XL�D�K��M�L��##�`���OvrA`�|N��3&�9T�i�C�>agM&��=� �5˔�,���E�ȅ�"�i��O�E� �.vM>D���dLR�7��
^���� �+��"U�&X��|U��pɺ1�u���`�b�f� �>�4�G}�K_L�>�B�K�Y^��e�:1�e��b*ʓ}"� �J�]V"|J�g�"-�	�(�	w4�PeIV}�L��O�>�0���Ϊ1x��0��@w�*�q`��3�.ҧ��«�=\�x�
�_P4���N���y"B5eb��@i��G�P��uO�����	N#�zbl�����/b����f,�%v����+D�(�ղN�p��oK���a� (D���0��7����o�-E�6�:�&&D�X����k1n$hfh9+�@pÈ$D�A�
�>=�����!�yg�j�5D��H#�щXq�Á̵j�TM�Bg2D�PC! k�$��&,T-3��<D��BD׬>6���`$�LL�A<D�|�6��2{�҈^�.�kԮ,D�$�$�1Rh@�D�pa
�� �(D��O�'e�M��րN��ԧ'D��(��)�f��G�W��"�,'D�XCD]�"�L- �F
	�l�� D$D�x���+N�4A��/�z���b$D��h�e�l��L8��N�qo`�!�� D�D�W��=�vHے�pk��W#D���Pb�	]ޝ+�NQ�_h��`C-D�LKfT)[(A��!M<Wr�2�&-D�Ę� X0F��M�n��S��G%D���$.�L�2E�𠜍*"�bE�"D�x�)Y�nt2���2|� �c;D�<�"%X( ��՗��C�ɠ+��H��[&~ZP͂�鋑J�C䉨J���0o0�Poާ
��C�ɻAX!�s�C�yo��ӳ��o`�C�	+6����Gl�\t�`e�7��B�I�c��=�D�ׯ l��A�,�B�ɶR�!����X���p�탺U�B�I�b�* ��� �j.p�0���N�zB�#T�x�o�#���tH�Q�B�	:i Dpف�A�Wۊ�!��@P"BB�	7G��r��r�Z-:�F�=-��C䉱	E�HER�VLp(Rv�C��!!T��$摼E٫��O�C��?2=8yw%��4������+��C䉓i#@`8���yZ�c<o�B�I�l�J�r�hʠ1�Z-�f�6=��C�	0A��9ʶ'"j�:�!QO�C� r~]AC�Q;E����k�8�C�ɴ?�$`��N�P���&N�v�fC�I?��A�ʚj�T�!�O>��C�	j�������Ud�ũ2�����G�ɉWmv:��|r�dɅ�S�w%��kJ�4�Px��
R��$�E�g�9�J�d����ED�N��	�1��1c�*�,\ъA��\��č78_�<��ME)����C`r���l�P!W�E���V"O<$q�J�ho���ꎖ`��ԁ��>����)�j��G,�@��E�G)e���i�i�м�5���S���~��!A铁E����A)�wlR��RO��.�'�Ȅ2��X���]uJ"�1-#p�3�P;G�mّ.C�Px��5� �YZ��!M���b3g�y��,4J�O�����b�#|� �Y�f�Д�ė�� ϐ(\�}����j�� y<�F@dN��3j��l��,�5F��M�"~n�2"����m�+>� ��2�[=2�C��1~���d��>6t� ����S]�ђ6��5X�>��DL�I?��i���`�Lt�f�>A�a}"՚B܈J6�?� �5����|,J!P���c�hA�h%4�ī��G?}��p��}=��I�d3�F[b�"p���^�t�?�hbC�0��(��+0�����+D��bN�>q	H�b�
°Y�#~�Bۡ"�>^�K�"~n���l�Pk�	4�T���:��C䉢$j�= �N�����H��J��6ʴ��V!��&������2��(V,?D��sIZR�a}�늄zl2�cЏO�G��8%MLbL9egR�D.�Ą�#�V!"* <_�DY��F!n��GzB��!c1R�_��E�^�9���.k��8���E@�X�ȓ\ \(��6
��a��P�E�(�l�;%����@�Hlp�S��M;.&;� ��H·]�pA`�F�<i��W7Qh��*`F�$-!���0�\yB��)=4�K�'`��B��*�]��d3w��
�'Z��  ��%r2�H��.l�xI
�'8"�5�Úa�A���b��Y�	�'Fi� `��N~��w��Q��Z�'Z�{�mG۸A�G+�0O�>�Z�'�J��1��>;鼭Ɇ��5�:���';R��
��%����[І���'��5�7��;X� �+��I+(�V���'���i� .]tT3���,$�t�'��@�h��w�*iB���ը5��'f04 �>;�VDz�n	�T��'S�5#�c�7K	�`*�ƾARȴ!�'o�˧�5|��wBĉ)c� ��'f.��u��k=��7�JS����'NDM9цD�6�B���ℳ}��9CדTf��xa�>A ͂�z{v1hb�6"��@��S�<��D�-Sغ�kr��/?�|D�U&Lܓm62�j�'������ʭJ���Y&e� �F���"OP���"�(�oF_�d  �<:�qO"�I��Y�Dゃ�BV-����oi�ó	+D����'���"C ֶr��8@\`	-�O~���޳�p���Ӂ@hL͒��'��Yz�,?��ضɘ�[�F͕P��,Q#�N�<!�EA7*��c'�M��18g@H�<I6���_��5h�m�ds����V@�<yeh�0t�P:P)@1����W&�}�<1�'!APֵa0)�Ph�r�`�@�<�G��x)Y�Ң�r	��*�+S�<��ش@PՁT�B�V��3��K�<I�˒7bj���3:�.�;נ
l�<�G�K�!�½ӳ�/-W0<0��g�<yS�� boX�".�(QI����#Z�<�����ghM�B�*{'o<T������Đ���"^�,��;D�tW!��?"a�/�n�h��w,D�8!���Y�TbA���jtK@',D� �UL�nW��PK�B"�T��.)D�l�`�ׁ�8�W��M�vd���)D��bP'�1B��0�3�G>F���e�9D�,r�n����ٓ�R��F���-D�pe�6�@�B�r�y�d�*D�4��D�j!���Ύn��#J*D��g��>\M{�&TV� 6D�ة%/�
-z���K;U���CRD2D���ۡU̪�AT�˴k��I��.D����E�5+'5X��ȩQ��5�7�(D���Vjֹ0�1�B�ƪv� u��"D�|y�T����z�¾Y ��4�5D�H�G	��A�2�O��&��L2s &D�\y֍�s��%���#s� �@b� D��H�j��Y@f��S��RE�s�?D�� &M�Հ]�AP�Ո-����r�"O��c�e��E��(��	=I�҉X"O
�1q�V�%fH���7I<�t"O(]��H�!^䑒�%s�J��c"Oz��ǐ�<�5�֤S��R�"O�����F+I�L����_�{�xpe"O��Y��3v�1��$E�B���"O�1���P�~=���t7B��"O�cb,ԌB�f�0snȕi��1Z�"O@M�Yw�Ii��y�I��Pa�<�cǁ�z
�����%0����s�<�CK�3z�"z�Ύ� Ԥ�Gg�X�<icEǯ6�@Ga�'�0�0�JV�<�$�Q�(�"�q0�C�P�(��Ł�T�<y7IJ2ѐ���I!�����K�<!��	��|�!k� ꞡ!E\�<�um��!,[�Z�**�� �[�<�G)۠v~���Э>T\���d �b�<�5NȊd �A�O��z�B�"FE�<��l�����5!(�C�.v�<ɣE"���j�S8�C��Ko�<6��_y����e�2��D1�/�g�<9�#F.6Q�'��0e�"�ؠ��d�<A$��	����E,T͢�"�fJx�<�3H3{	��b��ϫg��qVƉX�<q#����䅹M�+\�NDk��PL�<��C{��ts�u����\�<�����ms��s�LMw���YS� V�<)��ًv����"I��p���G]�<� N!-Ų��!�PҘ��p��[�<9��T+Fvd(vc�l�^8�!q�<��T x>>�郯��2��0���i�<AH��D_��u+
I��	�v�Ti�<��ܢ&U |�ՠ��|n4�R� b�<ن��6[�d�Q��Iw�r-�c �s�<�w蚏o�\�X�V!��0�7j�m�<Y�i�O��)�у�R�R���g�<I�Ɲ�G�p�a�	+���!D�g�<�rm��`��y�/Ȃ+�@���kx�D�'I �!+�}|��ƙ��4��'��ݩ�T;j�tCB��*;p�I�'�X��@&}��P����41Ķ]��'� D���&y��z�/��_�pH��'@��bv�E�����HV���'���/� ������X�,�Ш �'Y�с�_%4h��� k�/�H��'�
�P���Pt$�p��M�F<�-��'B�$�`�\�Bݫ�ď�0!����'r�b��b �%���;#] A	�'�v(8m�;>�zT���%�t`�'��lskܧ6T޽T����'��F�,?�8]��̈
J��{�'����e;�F�82 D�{܂р�'*Z��� g�$y�q�u�Pd��'�ɑs�����b�ūv��'������Ø_�t,�c�G����'J-�P��i�����0@��r"O��K�e>/���p���<l���Q"OT�0��%oa�w�4k�h�"O ���BL"�l�� f ��sc"O�Q��D�h03�A�c���"O@� R�9=��=����60\���?c��@�H�:W��9]�.��ԖOQ!�Ć�He�P ��O��m�"eO$N�Q�@[��� �0B�P&���ץ�P%"O&��I�)��q($�B�9��y�O�Dz��)N�R�T��V�[25^4�P_�D[!�DF*���s�H�"�PQ�eQ�@1�|r��OD,����͉{�T�Pd�yb��36v
a�6�o�a��	��yңT+nҥ�P.��&���y�b�-T+t����N���X��ϝ�yBH%o\0�QƏ_�f9��
�y��W� �܉ZU�^:t�`�pFdT�yRdT��	A$D�W �Y�ш�y���� �	�U0ag��&�y�ܑE�*�HvbG�F�9�F%J��y��9GӼ��LG�N����3�R%�y��L"##�Dq��B����y�b�s��lSC-��s$E)�y����@���[qQ,x:��	�l$
C�	 �:�%�V7$<��c�8_��C�ɋu��(��-�)]� �u�D�\c�C��&[>��S��� �D�C#s�pC�I�qG�a�Ciʤ���?�DC䉸=p���gn�36���h�o�7=�C�ɤl����CW7
r���Ɂ��B�	<9[��"���TD�L�d�8D�B�75�l�q`L�\�� �"V��C��G�xK�O��d�<AVW��OƢ=�}
��Ŋh� ��ԆY
*+Z�*�FS�<�ƀK �N��Be��:���a�|�<�2B&�i)��F��:�/z�<I�&�kپ����N{8��g&�t�<A�f�\J�I[��V~�5Àu�<�U)F�+�~Hz��\����ggXl�<�����e���C�ͻ���s�<�$�;	���`A�ag��a�l�<���9��$�4��9L�\�9V��k�<)�b��Rծ�S������[�
f�<��v���s�cv������a�<i�ϛ��h����� `
�j��v�<)c���z˴l�5�,�1���p�<	�KHk"�BAf�Q&8�C[G�<��m;c���YUK�}��p����A�<Y��!Eu���#
�0�����C�<�7#����,�]�N]*w�YR�<	 l�2($�ڇÝ�k���b%WK�<)��5�bDk	M?a@�� d�G�<Q�)ձP
��s��L�H*��`O@�<	��I�u}<��׃B�Ҥ�P��y�<�k��p�4�;��bin)��u�<	2�÷>�h����i �8A%t�<�iJ�h$%���rMn� aa�X�<Q���Q�B!g�ةs2u�0�FU�<�Ҋ��8�h$p�����*$l�T�<�L$Pv=r�M�q�g�<Y�]�0Ҋ|��K��^��D��f�<q��7�D�,Y���@ۧ�_�<�Y�P���0���`�B+5��Q�<��L��*�eY�޲���΅r�<��Nۋg�x���N��P�%A�q�<�A�B<fmjw�ҏ?��§MEq�<)�B$k5S6EUxі��ǂ�o�<��b�0��x����L�Z�Zt��P�<�����u���޿W�l0g��T�<�#A�e���2��;|�A�6e�k�<�f٠��(���S9٠@�*_Q�<� �cC�Sh,<J�O���g"O���ˉ��(���C�ح��"O L!�R�C��!r�3.����"O*����Tc@3GLM�H��zd"O�j �V�Q�d��j�E��H��"O���5�X�`��Y�iI��$�1"O.�Q��@�l(m��'X�E��$��"OD%��G�,%�hl�% �pж�A�"O4J�O�\�(�'��.���B�"O���/j�p�9�-Ԯrt�P0�"O�%�@11&cٮ;c���"OJAS4���^(��e��I��  "O�H��j�,l������4 ��*�"OZ$ZQ�:j(�S��W����{2O������D�٥ė��A*���T�!�
�A�pɣs��X�F�25�)�!���e����/�>��E(>�!���-l����PqTGѿ2�1O@�=�|� �׌CS��Ҕ��+MW��G�i�<q��4y����e��MN��� ��d�<I�P9Kwd:��Ѧo�	�y��)=J��Ӈ�)3fE��A#�y� �	ɖ%SE��0c ���'A+�y���b���Rh��,��b����y�+�G��HQ)	:,�n1#�/���~r�'��q�Q�.�Q�r$E/�*��''Z�#��E�!�� Ҍ��IĹ�'�:��֬ӷ0V�xvN�m��z�'i�
ro�2u Xf�Qc��	�	�'���w@��&���	_G4��'�d��Q� "N@4*֊�)R(0�[�'�:}(�Ϝ)/fȃ��S�B�����'�L��M�;��D��O�0oI���'��J���h�2�8��v	�d�'^��i��ytB�򥂽C	�=#
�'= �څ�T����A%�F��A�'���e"\�T�F�B��=��'��,P���02�^)�`��ib��h�'I~�r$"�y�V]�W
e�����'g>a���	;w��+'�:g�d\�'o��QG޹j	�TX��BI<v���'kht�q��EL�ع��Т����'a9e,��/[�Ї�߼[�e��'KfL`7��eE:T��	�(qLj�'�.�:��;�.0@���B���'3�b@֠>հ�N"8I��
�';<cw`ҫ��������;쮼��'^2Q[�F S��Q0H����'�Qcs�(��ʧ��O�e��'0�2�>�%"X�o휥P`ěn�<���#Q��5a���5*�<)�rF�<�S�@�]�T��#�"N�L�`��H�<�"��#2m�`�Y�Z{��g��]�<5��G���JĦ��L�'�E�<��m5Ξ���鍏m(�Ij�h�j�<	3-]8.@��2���O�X���d�<a��'7�){	����0b�a�<yT�R�~v�0�� ťR�x���Sa�<��!�2,��@�QPbV͑䢚\�<QoU�;p��3@�Ù)�"�!��O_�<��B��\���P�M��#?����`�<�)N" �m�7���v���U�<��l�xxt�%�͒RTV�2��L�<ه*��h�[��Íg
zyЀ7T�� ��A�g�=g���"��_�]a�a��"O�Ix��a�3�lV PG@��`"O����$a��|�F�P�rE��$"O���cE7��e�r�C�P��	�"Ohț��܈^�P%��N4(d���"Ob`k�5�,�UcQ59P*��5"O�,��D�'+@4H�ЀOaR�1`"O��0�b�!w�^�sbJ+8�I�0"O��J鞎�&I���`%DQ�"O�	�?�}�e�A�%�!��"O�c�*�7 G�8�e���:q�"O�h��L#���՟.�(A��"O���3*'v��p���d�J�J�"Op,0��%�r��� ލdC����"OdEȵ� Rb1i�i�/b���"O��ia_'�`��j�%J��P"O4Iu��C��=�2hզBE�CU"O�yi �1,��i3��ME(��"OJ� �K�>��FDN0v`��E"Oȴ���[�d���#��8 �d`�"O>q��
���£o�9���"O����bة:"���H�!$�Dl��"O����E�H�;�EB�=��DV"O^��l�l��tZSKƱ�tؠ�"O���!�,BE!��P�%pp��S"Ob(f�L+�8e/ݕN>�"O�=�֦�@�8;��
x�<��"O���Gm�+�8 ����k�LI[�"O�ɺdfΌ+��i�E5ELh�*&"O�\kc�3wˮ`�Ĕ "/sT"O�Y+�#-�hP��ʘ4�@��"Oֹ�D @'�: x����V,K�"O�lhFE�Ty�W2�q� "O�Д&��т�c�>E����"O	t۝<`�t91#D�/�F��"Of�@R%��Jy�tOՊ����"O(i`�Ϩz�LD	ao�n��%Y�"O����Q�,�:�+���	\H�F"O��H�HW/XzJAR�"�y2�"O��;�	^`Q�Pbc��$A ��p�"OZ����Y��\��q�B�j��U)�"O���?y:$5����<��e�Q"O�I�A� �3l�<q���<��"Oz\
�V�BZd�:�H�"1�D�5"O��f��#39T�r��I4EM���"OV݁��\�֬� ɓk���W"O��!����4��O)L�`8�"O����QO�5s�&�cے�c"ON���GV�)���Z8@����"O�@[Va�<dP3��]����ç"O���w���:�^�#Q�.����"O����݀\%XT�T�x��2"OZ��$$_�G��%���A�<Ь�"O�}�C�<n�\�`
��^mڧ"O�`N�6�nh��Pk�BD�Y�<��ø.0 耦	�G V�{2�p�<Iq��Pt�� E;$�3,Uk�<a(I�rZ���![�0�
�L�g�<a�K�i	`�%NP�T"̽ʰ��f�<)���)2<M�bo�8'�q2fe�i�<�6�NkJ����Us"���)�d�<�q)^�3�V��3$� ��x�E�]�<%���.��d�ak,h�a($ȁW�<A����^�����T�Y�<� R��AO�c�B<"i�-L\0�"O���(�@\V��(ѡQ��"O�)P͖�F�|�#���k0I"O���"@<"B�x�C��g�-�"Oz��s��^DĈ��Q�'�:ͳ�"O��ՋL�"W|���*�d)S�"O��P���R�q���3Y�@�j�"O��WkȪ�� С\�^�1"O�UK�ّ/�LAòd*ذ�P"OP�bg����d�a�L�Z&N��u"OPcnD&,�1�	�f����"O����BN�<����0��.��"O��+"땭&KҔ��$�
���Ae"O��cS�%k4��q'͍�/�Ν�r"Oh\�tD,�N]3Ҍ�4:�!Ӓ"O�ݫ���& �	����Ȁ��f"O��IE$1�4P���!�H�r"O�m���(K0����%a��A@1"O��i�j9[��xK��߇(����"O�`(�"A�4\����=�N��"O.��`�V,T�˃J�
M�e"O`��s��Fq@�IF)�<{�c"O��CE��r�<��.).h�I�"OR�r�^�)Iꀪ�_���"O�����?}o����B_`���"O�y�B4m����e��R��"O�I�5!1G
���'=F4�c"O�@*�-����P��7D(����"O��@)6G���!"!f�"O���%L�`y���E��{yۀ"O���*M�Jʤ�Д�̢ZoJ�0"O(�H�&�4ʺਔ�$R<��"O2MsP�X=.G H�1�n��"O���ۃi���w-L^�J�"O��j;Z䱠��X>~T�0:�"O���j�52��{v�O9SJ�p� "O��#c�<wf$��j�v?phK�"O��t�Dk���� �:}��"O�sŉ�:,(,���E�a��$��"ON�(��I%�ȕ�1���y"O�	���ˏC @��D"Z���!"O@���=D�`�&�?.�2��C"Ob��BI@�KӼ��]��n���"O�+7%[�8"��pǅ&Y���{Q"O���$�4,�:,I�b��Pm6��"Oح�q���5�f����֭Gb"t�r"Oh3���ކ����JR�� "O`�X��Nj�Z��g��*Y< ���"O�-����#�Y���N�e�H�w"O�@k5��a�,�R1Z$hq"Ob �4���^]�%�����4b���"OH|�5	��J|.�@v��O�H"O���O���2͍*UF�i�"O�)�'�)�v���QdHl�"O�؈ǃ�=�su�:Ojh�"Ob���ӣ|Vȱ��Ʊm^8�Y�"O��ѠC�mM�xaܸS[DS"O>a��%@�((��m�1z@�m��"O0H6ˎ(��\�e�ͳ$ܠ�"OҜc��ƫ4x��Arj��A���S"O��J��͚$n������	pT0�"O����mJ+0F|sA�"0ހ��"O���	� 3T�pV%�,��U"O$|t�ҭ���� �!t�B�"O� *�Ig�*c���"�C�arn�*�"O^��r�Ξ�X:S�\6>*Q8�"O�w�A�Rm`���x�aA"�s>)�픒;�@RclDG��t��OD�=E�t
��:0��(�`��&��C$O� !�dCB�1��E��h$
A.x)2�|b�'�ܬK�Iߝ#�^��F�ۨX.ҹ�	�'�l��L�.]��
�KA�j���'�H8[�˧��T�����>�l8��'��1�U���Nz.����nUxy@�'��3���ΩIѫj�p��'V� ���ӽ2���
������yb��Jռe��4���Q�_3��>��O�|����Ѓ��B��i�"OJP��o^&*9�܋�@�v;TJ"O�<2į�Z�p��Eh�2!�t8$"OH�P�,;\�p�I�7��(qf"O��W��X��&�Ϙ �,�)�"Ot�2󇌚`�Fyc�S�8p�Y�"O:4a�oD@Պ��3���\�����"O�����=3U����=��E���	N�HH�Ή>�\ĳ�
J���k�%D��@�I�>W���2,
�%Q��!D�@�5�@&E��K#�;rK|���";D�`�3�
�<���iЯ
�I���<�
���D�6�':�ѵT2�Q�ȓ��hR�n�&j�.E��̋ v���?��?!2�+�(�4-��cTE�2�n8�ȓhX�Ѳr o&T�h�"Z�p猘�ȓd��=�SK%&R���Vb� qNF���pz�3M�d8Иh&�	&�ȓQ(�}�B'=!|ɴ��7����ȓ|B��Pp㋔9�հ�)�a���Ijf��'FJ���GK�!<|�	�ȓ �Y���%�x%j׎$4��ԕ'�a~���9|���ɐ'AmLjI�s��y�m��"��$@U��_��Y�'8�y��ŁV0p(�ԣA�S��i�!k���y�.���<�a�D��G�vT���y����o�zY��%?�
 A!�%D��9VG�>	��T�L?O�B�,"�O���*q!QW=H$��E�ҁ4R���IF���������O�?����u�e��<D� KsO(T㚍��AV�;^5�=D��Jt�K%t}(0,U�s{L�s� D�,QR�P�Q��-�$�:�k�*D����"Q �\�Bb�Y��xV�2D��ؔm׃c>�D�G��2Z�ؼ����O0�=E��k�d�L���Syv@��F�x�!��A5+,�pVn2rd�P���	�!�$�1l�4�S�R�~H��t�˄l�!�'F�]��fQ��y2c����}r��,CHo�H#���S� (C�A�O<�=E�d�	����V�C;n/v-iD�]�$!�-d�]c�kH^�F4�eG��L�!�,U�=�5��rxA���� !P!�$����
�N3P�pijEm]oJ!�䐉lJ9[Q�/~�d�+!�2!�$ĭu�d��D�+}Fl���R1!�$� ���q�U8.ƢYW��>&�'����8��$[�,���B|�{�K2j���?���)P�5ǖ({` ,�b��4�	�I8ў��ᓙ)`�E��FL��uy�(ې9r(C�	�N��`�;=Ǿ�`EJ�
%BC�)� �,�a��PU�!�× ��!�"O�-pS�ԷB�RE��ɰp��e�d"O�hh�ȋ�x��E�\�t8�"Oܥ�A�P�t�챋�Iƍj_����W�O��Q��ș>f�h�@).�&�����D��V�e�O
(��뵥m5!��Ρ"��A�w
P}B|I�ě4|!�(T=��Q�HQ M��jGC�:!�����eD���rd�Q!�DSez�z��Ϡd�����3L�{2���m(z��6��<S�X9��Å����0>1��
/-V�\�F�+�t����B�<����1>��Q�*2J8Hw�
g�'�ax2&��=��C$F{d���Ϣ�y�"K4;�X�G��:�ʄ���F��y�m+�0ˇhG*41��95��7��>��O��@�R(���P�$��5���cW�	Y��Bw
̫`'���樕�0�9+*�IW����K�R�òMP�c9jD�q�K�N�C䉞�ĩy�*.���3��I�4e���0?i+ĥe�L @ː@ܰ�U�@�<!�O���yhۏ?1X���!�x�<�Ì#8Վ��D��`J���"�t�<J{�Y�a��x\�r�u�'�ax2H�"4T��0��Ƽ5��Rh����'{ў�OGt9Y%��$<�x�k�v��Us�'�q1��ڈr΅�@�t>\Ly�'���{fA�WK�E��%�9Ǻ%��'hء��)C�>�K����̽��']d�맅�3)��H�cZ�H�'�|���揓��q�@Q!xE��'-dM�X*>@�2��Q�IU>��/O�O�|c>�e�+<����"T�%���p�=D��`�@�2�!Q�S+4(H�8��:D�X�ׅ_ v���뒙y�ީ�e�8D����K�w��0A�b��y)�-I�;D���q�B���ا-Qޱ��+D����L�;X�,�qs�9 �+D����A!�H�2d��qy�]S��*D�@r�O^�W�Q���� =����,&�$2�O����܌�!di��F�>�S�"O�UrE�\6�i�#K]>����3"O�Pi��߂l+
}���J)� !��"O8U2�JM2}�f�9�	��F��}hS"OaS�n�X���X�i��(���R�����S�O�,�[��4t�0�!�D�}&���'�p|�B匲5Lv��S���3�}�ȓLՀ�k�%�*��ta�]��d���4�d:�b؟'�$p/�at(p��M��Ze�(o��g(�����e�<�`Z�4zX���W62
\���D`�<��Ҹc��qb쉵{��DS���_y��)ʧpʢ�@\;l�0Ԇ����ą�0m���uaB�@C�Q��.V�\Ѕ��ev�_%x1��Vi�#,1RU�ȓi$��Pπ>,[��ޡ5�х�2r��`F?K�
Y�ΞI8��ȓ��A10��"z�:�#A��(U%��H����T�}�"mU��c�	�'���'�ɧ(�p����]�g��.޾}�"�"O-�B�A$r.␻���0|��3��|��)��Z�(`�g�
�d�\�jC���Ԣ=çc_�0�e�F	�f��7oP2{��ȓL�H���>�h���¥C�8X��S�? rؓ�JO�na<�;�k�&z���'3�dՠYp�u�q��$t|��rץT�N�!���3L"��9Eo�N4�H�[-R!�<a�|�#�ںxG6ܪ��J�.!ў����zu��2e R�G:@�� ��Y^�ʓ���hO���6)�P`�)�5y�)$kB
[!��ե��ݠ��`ɦ�8��*<&!򤕫J���$1@���$���H�!�Ě�f���`�7N���Z��P5t�!�X�ef\�@@EſiG�P*���$O�!�T���n�5�å�ێ#�!�o�]����k2����L�F�!�$���l
�H&�g�Ɉs�!�
0
pRhy�-��(����M�!��I iEj���ϪgbՈ�F1O�!��A�1�(Hw��=f�:9 �	�!�T�R�H�V�T�Q�	_�-���x�b����dڙr��s�A;d�V��!� gx!���	.3r�gd�.�*�`��̶_Y!�D4s�@])��J��
d��A�zf!�[�"��䛢լ�c��OYZ!�$�<?��8qp)	4�d�1`G0KY!��ٸ.G��醗��Hp-V�H!�$�:1�I�� Y�56$H����595!��i1��R�@̉*�xQ!SN�?�!��S	0bH!��oZ���M�#� T�!��"#K�%�P�۞qQ���^�!��&,W^�"�%G&�6�y��͞0G!�ā/<1V�
V�˭;�ޥ��$_�y�'�1O��h�f�="�FDA.�!D�tڂ"ODu���Ӂh��0�2NO�6�͘�"O<�2SM�<\��CN2F2���"O�$�R��̩06��B���"O��0��N"�3�IU�O�N`��"O�Ԫ��U:d�KXQ�x��k�z�<���Uww`��� cE&Y w,�P�<)3h-e܂ �u,��x1X=�D��H�<�hG2�\ᘑ($IV贚��m�<QP
i(J}�̠t���9FƆO�<9CK��;޶��6
Ýv�4k m�Q�<	�ɟ}�9rs�o�h�
P�L�<r`�i �!�$�-F�0���`�<	Ţ�4O�H�{��$h@�ҫ�S�<�wD�f9lp�EWmoD��e�<qS�Q��|�Ud.{Q��q DL�<!�ʏ9[�"1�ר�-x[�2Sk�a��0=��LxU\��&��h��&b�<a�J
@��PV��.a.�
���E�<�/�,8�fɡ�%V�d�`�bc�\�<頢SI��E#$@�$9l�]���|�<���A�'�ƴ�Ea/�Hl��Xx�<�Dğ17T`ŉ�͗$�0���s����`��= �M@u�����^� A���#q6`a0�̜>�e(�ɵ;$2��ȓz
�(��@Q��\)�R�@@�@a�ȓ ����˛$X[HY�3�[�X{�؄ȓ8��h�E�B\:��  
vN:8��2=��s�ֽ	6쌘E	0s̥��9��(Х���^ء��^!� ���5fL-s���GgJɉd ϝW��E�ȓn�"��?�
��/ԯP2�5��?�8�n$}��BMв����ȓ�Z�8`����Zc@'{k�]��S�(=�6�ڼq}�l��$4��u��S�? �ˇ�ЩG����f�3�jl��"Od<���
	����AI�;_���"O����C��b� 4��'I���X�"O�{T�]	� D�V!E�l�h���"Oniq�	xah��EgK)`L$�s"O��[s-@�k�DI�уD5}��8��"OJ�@5.��&i��±��*/I[%"ORMk`닩q)(�A�C��F"O~y7) �(���qv��qIlл$"O:T�@�O�Foh	#��(&/�I��"O�$�4b��I���"@Q=&��"OP"�HeQ�,RE�[*�Փ�"O�Ta��++ �ł���:m��F"O\t�VMHa`Xa��D
�`)B�"O>���!H�Z�`T��"P�u��4	�"Ol=�����-��Mc�BD7Q�pPp�"Oq+��[3hB�P%��6�т�"O0�#EѸ+ *����5Щ#�"O@��NX�B�&T���8bZ �"O��:�%��0�z`��K�:y� �"ORh	c"��1����jb8���"O��@Ͷ.�BSO5Z�(��"O<$3䫁8w�n5ɓ��,lU����"O�l�`O��C�@�y�� 0�#�"O8Ta�풯)e\��N�! �A�W"O�C�.ϳ'it4��ZN�X��"O�:7c��E`\R�,�)���!"Or(�A>Y��`+&&v��r!"OB�(��9?>���� O�`(lh�"O8 �/'	�m�� N�n*�("O�|����0�{r��.�2L�2"O�ؐ��(R2Ѐ&$Y�SȒ@!@"O�)#�F5s�Y�(Υ�p���"O\Hs�@8=n��h�������"O�+����L�q�Ϫ.��� #"O��+@��-U�M;�/̸ �~m�"O2!pEB�}{�1�P���0�Fm!T"O^��5ܓ����k�jpB�"O��!�'
.�4ř��YXr"OR̓`�F�4�@�S�!��"O�Y���d6��)A����T"O�ܒ�� 1M*���"�|�W"O��燏�"��qፘ�V,�,��"O����)L��\;��3o��#�"O���󃘟PnQ�a�+vhyR"O�E���!Fldhr��^��\8s"O���U�i�� #��ph�`"OM0B��~y���B��#�"O ���̚,�"��DA)j�6��"OF8�� �&.�EJ�E� ��hJ�"O"q(���( ��Ȁ�$=ga�i���A�O�`�d,]�
�*`�an�/�����'�y�"��Ut����(/��P�'�L�B��-;�\�h�σ�u2����'DdAg�P�y��}�wI�7i�y��'���c�R��'`H-��H�'� �y����q��H�7E�T�'ҔH���E5��`��T8~����'����HԻC�$�`�@ԺYL���'ؼ1��M�HMJ���	On����'@d��C�����K�85Zqi�'�Z$`u�Q�8�H��Ĭ'��(�'Y ���%�em0��sG�����'�}�go�.�������8x��� |u�â�L����0%@(%"�a"O�eJ�\�r)(D��M~	����"O����l��,��ԩ�%�=�� ��"Om���R��1I���^��e�"O�1��b���n�V!����x�"O�!bS�<b�dAZ�ꤕ#�"O��j�W�H̡t�F��Y��"O*���N�3U�miR��h$�s�"O� :�/A�8ʮ͒��L"2��mxV"O���ѡ���0��SlX �� ��"O*�ru�a�P�P��"�����"O �ڥ�UD�A)֙6��K1"O�xb�/��M!s�-�V����3"OHX{� �, hejd,�9ZZf`x�"O2���4O1��ۂ�����]�"O�E�`��(C08����x��"O��pQ!(~n:��$�O�!}�a"O��z��������.V��F��"O�=p�S�V� ��?����"O�5���֊|�
�F�L��rp��"O"��AȂ|� �+�#��?7<��D"O9B�E1"���&1��5�"O�1)!BԅsbM+����*x|Z"O��JB�լ�xY��C9^v��RR"Oz �p�r�:�BW._Q���"O�i�@I,'H,�co՚lG��s�"O4�귏�,����Ї�,6�AF"O��Q�
5����쇗FV�"O"���n���;�-�:����On�(�ZI�ڥy��Q��][&n7D�d	����SS�+�`���uy��2D�������K��aa) �0X����+D������g�H:1���m��+D�l�/�	-Lvɱ�*K�@��X�1D)D��ƊI @��	r�E+�ڠ@��+D���-�s
��@e�!��|jr�/�O��	�G����G�hl@��L=[�6˓�?�	����M[�lPs$C
r���`G�Є��A���񩕆[Z����=�؀UH�ـ��":�Y�ȓs��t�W�ߏ4Ό@�	7O���#��``F�e��T�a�ߨ��Մȓ?�2�Z��[].�(��!}����CHf��Q��`fJi���ʙK2���ȓ.�lX dʹo�`@�  �u�ͅȓ7Δa�K��{�$���>a��0��.׊���o�i�\�!�T�j^�Ԅȓ:@���t̓b,��ۺ}zb���l8�Ya�ɝ0=���VÉ3;d��se�p��E;fU���c@�A�ȓR�҅z�
]��Gŏ>,�@�ȓo�"���K�,��a�v�<X��>tA�_�vh�Tip�XM�ą�LC��q�JʻAl�}Z�͞0��=�ȓ-6��)��0e�0� �"T. Ąȓ- �%R�V*�b�e�[  `��+���	Aݲ6���M�'K*$�G{���,�9l��<	]6�
��W#���y�AN1_X��֔%"�tZ&�/�y��ݯ}�n[E �)JtH� &�4�y�l©"&,�UkS�j��P`�ϊ�y���+<Ӽ���cMbY0��7�č�y�%�K�ҜS�"^$lG�y�욬K��L!R�Y�%ā8|ʘ��S�? ��R'aV�M�<�s���!)��"O�Ա��4C2��:gL��p��"O�A�S@ŭ\��6�.��"O��
��E��|�Ů��(�N؛�"O
(I����y^��贬]>z �lA"O�����oEl�[E郯6b-�4"OP����	Q=ҁh0x�z ��"O��b`'�L�Ɲ钅��F���"O^\�2e�>kXD�p��v���"Odyx�Y�3Ɓr��#3Z�]�3"Oܵ�7.\T2��E)�4HT�a95"O�푣�R�p�d³(@�S<!��"Oj��*A
[FP�����V9&0�b�'R�'����h[F5�S���zh
� ����f�!�D�J3����Q���aPZ= ��l��0i�O	sR%��+Q�F}�� D����"��e�آ�H�1���,D�����k��I�eŏ#��@�g�5D��� �j;J5YUGM��\�ڲ�5D�� �U5U�
D�uB&� !�3|OL��y"�+=X(��$�5F�*��p��6�y"�0}O��P��YdnJ���%���0>�/M*T�ź��A@�N���bNc�<A!�|,TP�rˋ#y�|�R��\�<�� �~g�j2Hװ.4��@�Z�<��(T�i�������/p#�A���z�<9�b�ivp��BKʥk�L���Hz�����ȟl�).�ʁGןx����đ�I��9�ȓ���b� w��qCh�fة�ȓ$	<�Hf�R&x�b,i%�%:�<��
�غgɠ�x ��H�¼��s���b[;,���s�I�+��U��#�����B��cf��O�����c��x+�!�-3#�d�C�-4��4��L��8�E�Gdn�@"��R����5pE藚�Rd��T:ӊ���/$@�r��#�Q0��V1֥��Xߞ8��h-yc�0@�ܼC�u��:��h$'��2�(��$J�1�*���
hyQq����vEB��8W�͇�z	1V��c����D��7��̇ȓ�H8@����P0�c�36���ȓS�P��H3{��b`
8Yc|��Ol���az5t���8cR��*
t̻ �-/2��b��3qw½���z!`*�%q3���&�72�r��Rx�k�K:/�<�tm�=���ȓy
�f, (�6���3 *9��j`��J�>�-�牔,5�����l���o@c���m՞Ql��U����(�=2x2�BP�P�"J����`�2nן-}8	�񯊋1̆هȓD���(�ʏ�	�Y��oXX:ԇ�9�������4A)3��ۍ=�杇�^�>(��L>D�:�!�#��m⽇�`g��� �w�ց����
�x]�'T�	C����&��@+�b�����#5c��'�fB� ԅ�BW�I��	4m�EB�I�Y<�}ss���<̘����N!8r�C�I/o��������p���H���C�I-�0T
FnR�
vd���Э��B�I�[�(G�0� 脫�/�(�Ɠw"��(2�W�>"����X+�f�)
�'!�y F, �z�s���~=x,
��� �u�emn�ؙ��j�.��[�"O�ABqO��;��aw���<∰��"O&�(V/ʀy��p��!�$"�3#"Ol��wJݠY�i:�w�P�'"O�YXs�'-�EM:��i�OF�GkM7 Y�(;�H�^d۴�;D���`�� f�=@D��]'�	�:D�t� ��s��yҠ�ҺxT<D� ��"�8 H4�3��;6_�`��m:D�p�`ă+Z�Q9��16����*D��x�"p뚥�#(��^ތ��4�O�I�qy��1�,ΤF�`j3֣/�\B��6:	r�q�(E:oȼ�D�H!�?1��	�9e���w��x&�����9�'9a|��O"M��k�Ń�Ρ��ȟ&�y��ݦ15����@�eJ���yR��v��a� ��<Fg>�yB����gB��H�풤�G	�y�	����<��V&P���Yw喂�ybꄻz��A�M��L:����CI��y��07R�
%EX�T3�q��S?�?�����2�jW�G�LĀ�Z4�^�Bj|܄�ed$���A }�]�R��,v���ȓz�\XX��ª(͢��P�'	�H�ȓ&�D��'Mݠ��2�$&1����s�йХO��{���9�(�D`V\'�DE{����98�A�U�6Y��Bc�V0�y�M�>[H��b���4D6H����y���+z`r�8f�Ͻ��j�d��y���J
ҙ�� ��}��"E׫�yҁ��TI�}c��v��ҧ��y�Q8&a����#tc0I+��ˏ�y��.ϲᐰeN.b"�>�y2,X�{�l��jk��Gb���<���KUM;a�s��*$���U!�c��`�j�^����m��/�!�ɲt���(GǱ@�X-�v
�H�!�U
hw��%+�Np`��֥+�!�Aۢ�p������BD�� x���=>�|�+��HO��{��'��B�	�q���w U�ga�Qs�&fXC�	'6�#���	�"�zq���&ѶB�ɥ �2@�D $F�(�v��B�I+�����R�@a�!ڋS�C�ɋ:��y���%&��y�EE��+��C�I$1���L٢���Ba+�*o(nC�ɥ`	�����%/<�zD�\�F{��O&8E��`��}��&6xAK
�'3\���K ������T~kV����?�#�B*rb�ZĄ#L؞�P����y�!Q%x�Yb��E�o����V�F��y�f
�!��I�2+��qGrẆ�jI�ȓZ�䈕ߧyC�@���H
g����x-~DZ O���2�z�U.^�����e�����5 �\�f�	27����b�B�x����V�J<�C$B%$���'�a~���?Ot�����EłQ��#H?�yb�!]%��pë�'oX�jP'N��y��آ<n�H���;tA��o��y�d�� ����ل����ˊ?�y���qn��N8 r���胲��'zaz�!��a"nQ{�Ę�n	���� 5�hO���)��B�q�rgW��1�d��yQ!�d��d�ea��Ñ�1���>-!�� �s�$Wj��s$.@&d�]pq"Oڈ�AEɟX���2x攍��"O������Z
�(1*4Y�܀;�"Ob])��M�N�������Q�>���"O��(�@�1@M0}�$"֟,�>5y�"O� �S��0��xg�V5s��#PP����	5�f��e�^N�jJ��� o#�ψ�,!���C�m�"䘑�NR5�4��"OT,� mV�2͂|[�n�/BD q"O͛
�?*[Zt��6/� pG"O��x"�?=`a:$� N�j��'#1OD�R�;)e��SL_=x02��"Oа*!G*YJt]�k�|�Р��'<!��	�C�R�YSDX�-��,8��g��'�ў�>�3�	�} ��pfA�',w�����9D��eY�o���d)�Vݖ���#7D��:��J `��V���+�y��-3D�, ���!_���ǁV�\)a -<O�"<��JX$0���W.�(+&NT�<�f#ה.��d��p���@M�<aR��CS4��e� �T��q*�$
�$E{��i��8�����D |((���M�WUtC�:J��q�6ʝ�CNQ��k�lC�ɗIt(��#��/���S�`���B�I38�>9#v��� J��)z>RC�	z2�|�GA�27����-�#֐C�	�_��T�D\M��"�(n<9B�'�1�f�ūcd�Ē7���N���'g⵪e: ����ĝ3�nx�'�d��%G��)X)Qd�N?-ռ�3�'������3d$	�����8\�P�'�|�� n�� ���Z7A��P8:�'5��f)�iB�18I�$23�BL>����IRU����UƂ��&��+�Sl!�d�*{ j����dwT Z!��Ƣ<p9���61ojZ� "9�!�ѐI����ʱo���n�'g!�D_�`F�x�ƴT��BѽPb!�$��Ϥ����OJ^�Kv�A:{!���Kl4�#'J�kB����ɖ�w�	U��(�Lȑ�n���p��iz|�$�6"O�U��B�Z�����g��<cj�T�	\>����^1
(��ጮ�(���:D�*VÓ0^�t|�#�̹-���X�"$D�l#2�:Npt+`�+g�L�W�!D���gc�<;�%�`L�<�L ��,,D��X���K��� ��m1b�ѓ�(D�p�6�Bc���@�״^?�+��:�D4�O�0��h	� �0��|�^Ep�'��I}�4�4���B;�� �m�����v"0D�8�ԩ�8O���E�-?��J�-D�p��������,�=Wn� q�,D�l��H�-��,�'g��jՆa��7D� "Sk'1`X	A!F�5o��#�7�IF���<��J'Q�d��|X�C�*�XC�I3��իu�2
�(��Wӛ)�jC��*V�.�ȇ*	��1Q5N�?EpC䉵���BU�h5JC!I�`C�Iw+�mK�# �$����NB�>�2C䉾=����,�Z���|C䉍T�����Q�>�&x�g��> #�B�	5	a2�b��V�YWL�B�@B�	J��pu�@7X��a�f�4UG��� ��Y��'|����E�I㠍Bu+(D�� PY8��\���3A��=	�"O��k���VFT���b�!��"O�!�h;$�����)F4B"O|�⣏*v|*�����+TH�"O�ј`�یl=8@R�F,}h0Q*�"O��!'H��8x"�fB�-���*�y�ݣ,��\��
W=0Cp,��%��y�h
<j���"],���E����'����ÌF��~5so�A�\E��'�
��c+��a�>�RI��'�!�R�N֠T!�U>7��p	�'z��Ǣ]�U�jPF_�0U(i3'"Od�s�f��Q*a�DT9Z4XK�"O�CNT�*�����Dٯc�Z���"Ob�i��C#zԂ!��a�����"O�}�#�6Vx��qB8m�4)�3"O�8jf�O�[bTX�C��s��P8"O�,� �[>0�r���N�
�pX+"�`>5����+Y��j���Xt�3a�.D�<Y�j��r��P��Ǘ{�j�p"�(D�l��MF;�������d�y�;D�D#��W1*0� C<l�2��3=D�DkD���X��3)'qH�Dxu�<D�Ȋ�HE�B���^�AQ�M0�*:D��(�(��B� F\	�ZYH�;D��X@��q���x�HV+6.Y"e�8D��0B�O_<���k�^��I�	5D������:F~��T��"���KB� D�|�_�Yse� +ː�j�ǜ�P�*B�ɉ _lm8�@!M�x��b/ƟX�B䉦
��5�m�</�\�ۀ��Id�C�	�-��*ƥ�s3*�R�F\2upC䉂-�l��&�5jBȏ 8��B�I9O-L�S@NZ��1��S�|H�B��6?�(BQ�O�Asc�,&Y�B�	R� l!!c�$_�ΌRgOP�#s�B�	0\f����D���ÇmY��tC�.]�R�Xr�G�V�l�k�*�6C�	$h~�� ��4-ߺɫ�EO�?��C䉓&&���O�Y[vkG84C�	�	P`hj��Y�\p݊6EG�.��B�I'g�~!˂�F�F��R��4V�B�	���騇�R,	:հ'��3}{B�I�D)�IؠB�E�F�sS�B�	?���a��G}�)4�˂�B䉎J���2��=8���f�I3+w�B�I�/@�Y����"���k��	or>B�	?,�[h�<����ѨB�I)�h`�1��,}��:�+��>��C�ɽN�f|���A%MaZ��G�Y2c0�C�ɀ6���A�s.���GX�"��B�	o������0s��a�7Y��B�I�"X�0JQ�c�P��dֲg�ZB�	�΁�#�W4I�v�q'`ӐY�`B�	7s�S� I)GDb8�g�Q#,�\B��\�B��d�@�TZ�ea�qdC�	�J��	���'p7��.�$��B�	�[Ҙ9�,U
 ��u�ެRJ؄ȓ?0v�fi	*{�6�1��J^�=�ȓt)�iK(@�X�p��K��H��R|Ĵʵ�-�֩BC��[X�ĆȓuQ��/P�A���Ѝ
��� �a3D��`A��< �P�	WF�P��ey&*,D���� A��d��[���K�D*D�� ��A��K<���=a� �u"Oh|��^8V��A1����"O�P�cI]	%̼����T+f��Գ�"O^�����+bH�0��ҕuO.%�T"OV�dh
��B!�^
>F�j�"O\X:Vb�1CO0U�A,� 5V�zT"O�p:df	�}�V�q�a�T�Qp�"ORH�q�C�>0�iS���2"OlQ7����~�aOܗX4� �"O:r-�*8E�c��]+��k�<�W/o3j�����	\9�Tj�m�g�<�@�׮i���
�m�WAN�K�ϜN�<���S�92x����%^4�˓bR�<Y�J	�p-����!8�uL�d�<!bg߷̘�2VN�t�c�u�<�"�H9G��5� �>,x�o�n�<Q�ct�څ�GC�1WĈ8Gʏh�<�ro��\(�p���J+v�3v��M�<a��/��5i�J�e��%p�#�@�<	7T�.`b����r��4�z�<a���'��	���X����_�<���ڼQ&���G��w1\ԓ��B�<)3d�ks����.��-��K�Z�<y-B�1Q����L�*s.T��CAS�<	g�I/�L��S/�� pA��H�<��'�5h#,A-L,����"�k�<�D��"x��Ea B߬��+"�R�<�#�aߴ��g��;i,�K�ƇL�<	��X.�*P¬P2X��
L�<�I�"D_<��6�Tw�Ȱi��]K�<�6Iú5��)B���7nEa2�G�<�L�"�,Y�O2�AjD�<ٲ���YҰi�L/��U#$EHh�<)��;�Z��bg�$��Es��b�<�7�;�A����5��ɖ	\�<��Y5M��d���HYJY�<�t�&�ꍃ��?~�(��R��]�<1��'�0ͫ�H�8t p��[�<�`�+$�WE^�8cԑE`V�<�C�Ә�bԱ7��Xل���ABN�<�耥4���S%��\�%�"�^�<��F���xI��]��$)#d+T�@xRlM')�m��e�vFz�A$3D�ظ+�r���#1jD)Z5��q�k/D�T���3x����c�/\ ��C3D��z �A�ܬZ����&�$� rI/D��+�ύ��Q3���J�����+D�0Ps!F�}�᫵�
�M�\�w�%D������R�Q��I.C!ԩP�%D�����T/�����M�/D^8X��!D�4��qf���5�DQp�%��.4D�lSS�@A6��W-�w�ލa2�1D�l�դ�R<!'E"���ñ�+D���c�� S�ir�N�n7z��N-D�4a�g@�m���J OH���K�X�<��ϟ <+VcH�rFN[tb[T�<��螏,q>�Y�E,C1@1P�-
V�<�V��t�=ÁO�K,dPEd�v�<y��
!9� qL�@�����,u�<9�V�J]������=#\H��u�<.�&�����H����Q7,Og�<Q�$���j�2�C�_p`�H�,�a�<�f�8}ո��������ձ�y��/�"��VJQ�t���aq��&�y
� p����{���x�)��i��"O���ħK�� p�cCv�PAqS"O�xe̶�����	�%�ڜkp"O���@3TcŰ��<,���D"O���4�R�-�n��I�!�_� �!�Dʳ�0�Bϙ2�q��J�l4!�$I:1?z��IY�-,�y[q�@r!����d��$�^%����&!�D��CG`p��_@�D�%�D�J!�+b*��	ޑU	�[^���	�'����`ͅUIl<��BM))<^4�'�N�;'cC�"[�q���@�	굘�'�:)��ǃS��;��-j`4��'�d5ؑ��پ��W�[�|�"e[�'rF�d��FR��`��r�����'[��g׀J�&��$��p4����'�UB��$'?Te���+r�� ��'��T�P�'�41H��ؓc���#�'$�j��]�P:����TjZU�
�'����4�E����R�.KHn��
�'� ����m���ȴD��Ւ
�'��q+FCC/\��($A��C���k�':�HY�)Ѳ8s�5�s�D
jw��
�'��i����Dl���H�0n�Y�
�'��:UE���81@��J Y�ܜ�	�'�XảǢ���%�y@��	�'t����5^�9SrCw?��h	�'t��R*��x�؅����2�	�'=FA"tl	�j�plb$��/�t�a�'ߞyJ�	ҩ&x�2����z��5b
�'+�@@�KӕQ��Lx#νknE+
�'��PX��u>z��F!Phh�	�'d: ��OA��5+R/5xV���'�h��q�K*g�Q�23���'1$��c��WD b��L�t�D�1�'��Y�s �.�xY����!�1��'p.����}9J�z�_��pݡ�'��iS���7$P=qw��ĺ�"O
�U��S�.��3�Ra4(��"O��q�nÌpI���!�"O��1a]�@x����H׵i	0��"O�e�Ԑ�AǑ�[N2=�4"O2�1�*D�#x|�3g���'@���"O�p�h�� ?`Yc5�? X�"O���3 �A�\QR���'L�I""O,y�u�*���;&�M��1�Nd�<�?S@P���Q�P�R���x�<�񫄖l`8��; ?���!��N��uqef�>�V����ѦRZ%�ȓ9P�)h�El�
AkA%_2<��v� Q:�ϜZ� �g��x�.]����"ڎS�xp��	$D*�L��;����F�|���DSh�<��Ezr����-[�R9��+��X ��k#���1O	�Z��R�~� ��XZ�}��/f���jt�v;U���OR�=�Z����pe���\�zɊ`(Vk�<q�i��)9��J���0����E�j�<Q�m�5	h��G�%@�Y*�QBX�FybgVt~��2q%YXyv2�k�4�y2�\�[J.�aPETI�=aT C�����hO���,8���
����	D6Y��8��'��O޽H6��[�8�C�%�ft�$"ORԻ�L(=��M@f�˭A����"O� v`��/�5G�6L��� }�����i����.�i�p\T�AǇ��c���>���<Y�'��'ٛ�� {W�ɑT���-E�y�֯߫�yb�S��4��R�k�����H��p<���ĝU�jU!2���=)ūE
XBa~�&�|?��&��#T�<�z��M�<�t�^4���b��.�*0
��a�<��J��6!��2$g�t�!M�^�<	�b��(�)@��G+5���^�pjV�z����O�3���Q6�l��kƠ/� �"O�����ߜ0�\� ��~�
%8!�Ol���=Ѡ��	6\V4���A�~�.�ұ
F8�0�$IGU}�Ɂ$,��ْ&��Dm9���M��'�8ͱp�6t\�R�nL�1����'�I�e�%.��W@ķ2�ʹS�4�hO?7mչs��p�+W�49���Dњ���-��?��J>A�4G �1b�J�,x�,kgK^&|�|Ʉ���[S叵:u�Qa�A7h����<����i�> f��uH�3'3x��a��$ab�O����$C�4�&q�c[{��u��1LO�8S!g���̣lgN<���ɼ�h����Տ��P}�ce���A������������)�'Ƙy4 \6F�xP3@	ը,�.���	�<�{��E6}�:-r����h!�*Bƭ�y�蔅h��Q�\�S�]���K����wX��2���o�ܵΎ �%7D�$AãT�v��U��(R�a�6D��(1�2(�@��u�BZ��� D���"�
1�"�ʙ�P�@�1�)D��R��&��:�֏<cհ�I'D��6Ɉ:9$dr�H_E��=�D�8D�8��H��_�D́�nФ'�X�a׮5D�@'&�w��p�Eܔ
�jy Ԅ?D���Pl�$O��-I���.�"��=D�X�ōȌo�XI�m�N�xz�N&$�D"b�ׅr�t�w'O�4I#���y� (O�H�˦d�+@�V���Ł��y�|�tx*͓:�|��2%�&�y��%'���
`��<7�Z�c�U�y��עb3]KF�8zqR�۷��yBK�J�e����gX2e�c��y���.5����I�tt��'H>�y"F='o�U+�*�>�4Xjg�[ �y���1�8���14��ܲ�e@�yb���~����k�3&�=�P�L�y�B׶2�6��b\(-�F����y��Χ
�:�J�j]$��u�� �y2��0 ,|�:GY� �%���y",P�Rt89W��T�@][r�@��y�E���]�ĤV�PN�aԢ��yRD��#���(��L�|�r�3o��y�MS�f}�mZ�}��吮�yr`¢KI�Ah@GR��S��%�yR�ۛn��j$�_�S��y�պ|����#YXa�乁���y�5~�����J������y"Eʼ ��iP@��B�t�9��%�y�[8e�P5C��Y�n�
� Z��yb*O�CG��{s�M�vI��"ֆ�y��l�XQ�p�V:�e(d�Ҕ�y���J��ȷ��x�2h��hU��yRÛ T0~�q�a*u""�B��yB��=D� ��!ޭq�h�q ��yB������h�ꡩ� ��y
� ���S�M���r�R(մ�pB"O�C��Y{@�ؠ�O8|��DY�"ON)���U�!$����c�l)��"Oᑶ���VM��ru��,f�`��Q"O"HCF��a���q����0(��Q�"OD�we�7a�R��k�"Y��S�"O�`A���|�v�h1
A�#�"O^I���VY���G�V��#�"O�� �r�p����i"O
m �ꗇc���Qa�Ӿ]�������9LO��*w��B�$�F�Nf�1�"OP�����/y]����= >�U�C"O��K�HAuV�؃��X% 8n ���'o���b��2(;v�v)�><PHʦ�=D�0ɂ�I�>����'ƃv�m0<O\#<��$��O��A�aQa�����	Qt�<Iu�'2>�![��M�"84���@�k��0=!P6�\Px����?Yb1ZT�g�<�c��u��934`�4d"Q�C�ʟ����7$R}��hU)X�`ʠ#W�.]����_n��Fb����`�i�,ip"Ox*�Ȝ4#�G�V5d��;��'Q�,@���+��=�V�y%����?D����"Џ9+��&��p��\봩#D��+���*ZH�	֕^:��s�#D��
r`�'`�U)Y��j��e�?D�L[�쁖{�u��&�.$p��-=D����
�e�4AtJ׿2MJ�K��9D�L�� W�nv�m�ԋ��Y�H�B�mxӨ�1�)��ЖG՝k�Z�5�W9�lMڲ.;D���#���*I�pO�r�,��c��<Q6�'�8@ȷ,Y 1򋗾a����'�dK�(1�%3F�M%"���M��l�`�Dz�X6M�J�'���O�4q�AT+%2�{�J�OF�C�"O��P-����E�(Ic:�q*t"O��!2�J�)>�s�~/����'~�ɓh��i�%ّs����k6IV�P��,�|���צ<��X ��̓3|��$2�d�6V�\�s�K�JG"Q�"�!!�!�dˌ[�ntP�ͭR֍�oT�MJ��Ay��)b�M�0ɴ�bS�Ǽq`z�S��O�<���	&	�.��E�$	���K �QH�<�%otx��$��c/Z�8字G���d��H�*�晒d��J�H�EI����
�?y�Z���PB��2#�Rũ��=�'a1O����� ��A?����@	�@��=D�Tv�=� 3�Ý� �Rm��O^ꓮ����N%� i(Q�*@хc��&��5C)O��=�e풧>��@R�'Q0-����$(�צ����'�Q����ǂ�<�̩4�6O�����*�O7�;?�c�CC��(օ�+3*�����P<��ɝ�hglp��F2��yU��N�'F�b���ћ�T��8�T�B֙^08Tq��3�y����|�z JL!�Ⰸ�k�6�@�͓�򤨟�g~���X�EA�l�V8�p&A��ج1��+D���b�9(�H��r��*u{ʘ�CT0��'��Y���u��.O�(k��� X�9!�?D���0e *s�	�Gޤ��)�1*>D�$���^
9�X$�pl�*Ԩ�"cN?ʓ�hO�I?�%��A^6._��Qc 'DB�I�x�
! ��>�$-�th�-�S����OJY�3Hժ7
�k��E?�dJ�"OB�z�`�)64����0��	u"O�q��ԡCҰ� ��ӯ���!E"O� ��B|6�Q��ȋ<5��<�U"O�}:dw*�X��ŕ�f��Q��"O�������M����撑V��5�5"O��a��Μ~`D[T%�5L�� ��"O���Fŕf�ıG��q{8��"OJij�MʄAʘ�#U��	\�6"O�a���{p��6�J)B"O�ڱ���f��E���_����"O�a�ccR!��-�!E
x	�u"OĹ�	�$0��$��5��I"O���ɫUa�E�Ԏ�51J`= "O�ѡ���s��x.Z ? !��"O����զIxp3ã_�3.|���"O4��@��W|q�Q2�j�"O
A#RF-l�������"O����&��`s�֐�5B�"OL!��B��1�	���.$Dk�"OF5`������_+U�Dd9V"O�cs�#��`���=���"O��H��۞Sj`�h7�E �z�J�"O~t�ǅ�4�Ɣ 3G��B��h"�"OP
�N�=sC�� �#o�ċV"O�	q��/�x��W��,[d5hd"O��p����Q�����OV�#"O��ku��{E�����̀H$��X"O��Zv�P�F�ɂ&ȅ,B*�L�"O�!�)TTn�1v�]?����"Ov@#��1G���'G]&UG�Hz�"O��c�K�e�I[��ߵ \F"O��A�@�RfF��*B*�$"O�� �Ɂ b���aQ9����;O4Z���F��H��.���XC�*&�t���e���ҡ��*��5��'�\�:�O 9+��1O2>��K�'<��vc�9~Pt$��
3t�A�	�'���q*Ԧc��y@�K�^��(i	�'}�V�ށ��%��[�#z�U��'��X��h�;H��CI&����'�/:�@WIʑKG�a̞��y���-1��Si�@!o���y��W�)�i������H:�	��yǆdd�����.�
�P��Z�y���6�ܨ�
	�
7��p�<�ӭ��_NN�փ�8��8��UQ�<i��ߥc@
̹7��:v�+E��L�<���#M�-�'Y�q��s&�JH�<���0¦PIT/��Fa�E�@�<E"E�p���ȵ@�$d�ې�Z�<�4����{e+Ǯ]���z'�U�<��DЭ#� �@�*`΢����k�<Y��6(�j�PŤI:i�(8���f�<�f��퀴J�=�X!�E���yR��-M����̌�+e4J$���yB�T4հ%S('�тs�ʤ�y�GǊ3�*DS�֝NlN���E��ybN�@�a��M	2�I
�T��yR�C/����7�H?Q���ۡ+K,�yr ʈ��P�P���Lr�d§D��yr���H��4�d=0fV��y�ōI��eYDm5z�
���B��y"�
�}�,e�!�J5z���p����y�CS�Ӳ�R%*�܀�ٶ�yb�GP��y�)�/U�4�V$��y"/�1�dɆӛ�|�����y�H+z��9�W�?D������y
� D�E�њn��9�/ڳW�,�s"O��p-)~�N��g2t�"U��"O�M�#��d
�!KP��=l�YH�"On)��FǬ��Kͣm�2�v�D�M|�����@�9n`�S�C�C�� �T�Z�2!�Ƶi_Ȩ�w�E �jMɕ�6�`H����z�ɪ7�Q>˓/�>@Cǉ
)1#�Y�FB'aZ��\����KM�,�ه�E)p�Ʌ�
�J_�����2�O 
�N&u�~1��Ϟ!�ԕc��'�БǏ�z��9�C@l��0a�K���@�j�&��Gr~u(B�ńs͚�q`�(�ذ�<	!�]*���It�7�M��*���'m�� �*«Fj"��ȓy�.�� �*s|԰$��$,:���'n�|
4�'Z~�𙟰���W�+�Ʊ�W+��5,�)�.D�X�Pb�RӖ��k��|^ t�1��	"�`K�-X�c��|����D��,��V�2�A&D,�0=a� �)G��0Cb��?a�ST�82�L�t8����M�<17�U�N��h��j��pU��gWE̓�~}�3�ևpVe���&
��z��N�J/�%���'|��C�I�hR���	[��9��A�qȍI!&ԑ}F����O>����3?m�;F�y I֕=���b�Bm�<I6�6wʤP+gLY�EM�=���#d!�qK׬
�ẁi��?\O��qRO+N�Q��ˇ�>���'@�tˢ�	�	�I= @V�s1��"gJ���g�ǘ��Nv��3e��*YviC
�Wδ��>	��ղn� �q�����(�h��U�>o�n������Tx��	�"O��2�ER�1��2�_I��Mcp \� W<�Z�Ï
��)��<�3�4(�q$���P���D�<�����=���%NG�.9@m��E�<�C��.[�`���C4\Ojl��c�"6&p�&�<P�@��R�'��Rt*D�Q02x�!Ĉ��̭Ґ+Ƥu �`�ح�y��L�W:�T�C�w6,�B�Ĉ�(OL�x��U8�"}z� ����ȗ%�2QƐ@��V�<�S@5��H!��)	:6u���G�����(qO?7-ʂW��1���m�,T0eEI��!����!���N�,�tѢ��g�!�� 8�X�O9rd�u�f%�!�DT�
^��g�B�Ĕ�%U5a!򤑆>u�� ��V<�h��&�x !��ĮfB��� {�ڈ04�D�4w!��E�t�n\��@W�����FA�H�!�$�{�F��F�	y�Z����/O�!�ěS���Ӱ`|������A�!��/XVM$T��+J�E�a�ȓE�L8`&�v�P����D�Z4�ȓxM���Y�z��ؒ��%.r��ȓvM8<�GI�X���A$ L������L�T!"�� ��Op4��-B�`�V�] L��N�ON�ȓ|84]��N߶n���B%�L��Q��{ü 0�	.WY��BC��2DH-�ȓ6�����w�d F#���֡�w�<iIΪ\M.�rvlƤm�j`AF"d�<yA���5=�{e��CL
���$ n�<AT�P;�8��d�R�Eְ���Yk�<�����RR$��`F-p,��a i�<iբЖc�B���#N\��G��i�<Ʌ�W5���S!n�y�m�j�<)�P�
��I�f��u��ӳ�e�<!rh�:| �91i��eڬ���\�<yBD�X)8�1oD�� �GX�<�CHU�~@2�'��h�dM����a�<A Vl�l-��t
��ɼ5Jt��C��c`C"+fT��Eɕ2�T]��S�? 4�AGm�&f?6�3�=_��
�"OB�'�O{�fM�7b�K�2�"O�L´�)-����RM>:�"O���R��@�`�F�V���"O P�F)�2fm|�B)�.X��X7"O��3�'Q ��	����J� �:w"OFK�(� P2��@� ~y�-pc"O>�㛓�H�1MS�\���`�O<�#��D�;�f2;{|�x�Ꟶ_U	�'�^k2N<D֚D؃K�L�L����I8k�MK2A/�S+`��K��>T�@��Njb�C�I�d=J�@�����D��qI(����e�R	dj�ӧH�@Y� ͚5���`'d�:hօ+�"OZ!�J	b�����QO�mӣ�5}"�K*n�����+���ƪ����9\R��7'a�F��P$�D.9Mp����PJ�8�5&L�H��?��I\�s��|�$�*c䢹��NV�N(��
~�'�Zs�-�<r� |&?MC���s|ȁ2���
cU�Ӝ<F�C�8S"��N�"~n��*+ lvf��x��!�s"7-o��2�b�[��H�ӧH���0C�ՇA&j��CJ��N���?OXyT�F�>�\8�`��p<A�9�(q��ZR�T�#�N5��������7��'i<@moݸl՚�i&��73o<���B_Bn	S%�Хf��p#��'���6&͉TflbuDE5\H<3�����x�'�f�	�u%0����N�����k�ģ�z�(�K�)	��'Ԣ'��Eb�H�w�.` W�IT(tNA�2 �YT���d�'~B�j�&)P �%e��NDO.�H����P�b��q@R�l��M�i"r�6&�b7�)�'}���*􍉨/�@0��*ʸc�bQ�G(��@ڔ���N�j������%��Oj=�M�N+ݺ���<P�^��r�OJ}J��V����B�R���'[up`�w
�	1UX�*����0�𤘃!�6b�N��Ҋ�4+oT�:So�
��?��kʲhhD����0�
���+��8;��Fm�A# @x4��0�˱c|`���4�*�G�����qص���8��(��Ox� 8�J�[��s�� �ڨpq��v���4H� >wfEb��̈���!��<O���gצ#�Դ@!��^�O�[�J��|�
�rB�� ��U�Ɂ�ƍ��&^�F����"�4�b̧��T��G�38�`&l�Kt- p�O;Xj�`C�a�����׃֑�0�P8�7/�
^a	Fb'&#D"�bC8}@���aa�e(N@2R��aj��ō��(CaBR��B �ɶF�	Ì�)x��Y��͑���`c����x/AU�`tau�_8/�xD�pO�b�Xx�HG�Q:쉋�l	���`�I��
(��Qq6�c�թ�� �0�q�T�'%�1�UB+|ON�R2"ۢY/���f�@05Z6tK��0��E�r��G�x9僷�.	�!o�*B�Px��23V.\+�S�����c}��ѷR�vaR4F�-�Ҋ̦��'ZR��tg��k�Nłf���m6�h ���O��
3��	!!bn������C<8dl�m�%fE��(��0Уs�6�)x��" �$6N=B%��<vk�i����(�$Px#�Wp�S���*}��2 LC%3�$G�uc�A�GX���](��{��":YЧJZ��?��(�@��� u��423\���JW�k��,�h݋U��D++O�12�h#v(V��R-L3䝒��w���C��B�݀f�Y<a��t���'Ԕ�C���p�դ�(fL�m�%�]57)��Av�.>(\��'ꤥqQ�O2	�|�0��< �"�:���p�4�p��^~ҏÙ\d�r��BV�Nd��O���'4��Apច7��z%`X��t���Yh3D%a �Qrb!�
���G�ƸpPHB�"&"��� H@�|'n��j�`�1�fY�������$��ǟ5\6��yd�M �XX�o3zy�Q�UB<�(�'����KF~b<s�@�.c��� tM /�����'���#�W�D|qf��
F��#�n�����C�
*��q�'e���%�[���"�P/|���]!�qN[B�tݓ�kU&X���d�T�xh�3�A�B^V�AN��:�}��)L�H�iJ�t�`j�8T�l���$�:m�Fz2lJ!0z(+PΞ�M�A{E�>�0<�ca p�e��'��!Y�呚}�Є�$��.���Q�BR��u���J��E�
�@�����baIB�M��Ii�A��j%}�� F�����d���{�`ݶ���?�BA�z������:I;a�"D��cH�EҤ1ʵ�ř-���AR�L�����c��&�"}�vj߄D��,����REΔ��Ts�<!��ޫRI�l�5BǀGDb!1�)Ta�FFf)!��'ֺXBR��"�l�6�Oc*�0��'�.����H�*����._����'�l��D'i�Ŋ+V;CC����'��궨�u�A�M@4;����� \�IeH�6+�Ax��D�5ev�p2"O������2q~y1sCC�7lH�Q"O�p�4�MDjgB��CC6��"O�ؑ�ڶxU��SEa<R��D"O0�a���J����	u�H0�VoL�<�f@���D�Z�*�  �(�Ga�<١�ؓN1�ɗ�O&c� q�U�z�<�wSq��x��jܯMy��aҫ t�<QD�++�!��ʗ�u�x���	N�<���š\^��"g�M0*`��J�<���F2Tt�����#*8���6��A�<��D�W}�����&-�ȐG�H~�<qpn)n܋��U
4&X� �{�<�q�J+$��%E݀~t5P��O�<���0Ez�ӱ�Q8>��$����n�<��o:k"�D�KF,�m�)�e�<	�dܧ�X�{���,g�v��Ǣ b�<a��ЪYQ (�a�XS���k���a�<94��A|�`%�6�pX���@�<���ɰՀ5��B�?'�Ir�O�e�<	`��x��(ى�*���% i�<Y�睹6xRLJP"��C��}!��Rk�<y�j@2֌�����轛�
c�<A�H�\�<�{eE�9ihX��$��f�<a�`ȫ-9��°S�AQ/L]�<�c$��FlB\3h��Q �����X�<	QgB�s�~�KiX y�D�K$��Z�<Q�G��v=� �Fk�t�a��x�<)2�� ]� ��
�v���Jßa�<��J��%a���<l:�9�*�+{!�]0s1��襬X����Q�dB9
t!�dON�8��@� 9p��ງ���-C!��T�����74yʱ:5�K!8!��� ��˔�I9'I `��/4!!򄘾]��Z��v���	B$P!���(a
�1��)[�l��`. !�X=6_�a�Cݺh�r�8�.ųE,!�Q�Q����F�*g�pB�MĮB!!�Dya��؀@^R��LT�q�!��ӑ����	@Z�Y�+�9rF!�DҒ1����r�])ODZa���I�ZS!�DE��H,p1���\ �ȥ�d!�ӀU�fP����9�⍣u��7	�!�$� fJtӑG�i�"�s2'֘(�!��G�@E��%�
�|IYe_#n�!�E1I�~@��Ϭ&�N�k�ҹC�!�d�"l���E�b4��� T�!�Ě'uXԝ�j���z�X�"[2eC!�ds�YɃ)D4��ɛ"��8S�!�Dʎ&�:	��F�E��H��Oҁ?�!�D��~���r�۱!}"8"���v�!��ױi�|m�J�;m*e��V�3�!��$0��bakA��ƈ�k�g!���,V�|�4��:ђ܈cL�*!��.���,� �\|����)�!�Ć�bp�f�V�&j��]:v�!�$H�+���,Q95F��cR�c�!�DŜq��Q�S��~B
�����c�!�Đ�q?��H��>!@%
�BL1�!�$�� �Bd�e�=F\@g�F�ym!�ث{�r5k���P,\��eMYE!���B�(5�e8 ��#W�/2!�ݣ{��PР9��m(�b!!��8l`4�#�"�HXpR�S�D!�� L�������42���g�\K�"Or��%��	��$���.�\iS"O��)Xњ�p�Oek�H�"O�T끅@)gp��d$ �lf(�x�"O�e��/B.d�ɵ�Hr�d�"O.l��l^� B@Z�}&��"O`�0$����:�R�#]�5a�"O��b��4z�e:1c��o��DD8��*��I̾T�&��1��R3��)VE@�!�d��7�$2���E,V��!
8(Z�QsAb�I8)^Q>���9�+��:QD�h7�#K���ȓ= A�3j��/מ�b�C��!��������=���R�9�O�� ҄��kM�C6��?��p��'�9�Q@���V0�"v����FoX��4dш&D�ȓ>��E�����e�eG �3���<�5���5��9у�=�',j8�
ͣr	89�w(�	UT%��pA�ݪRe�Tr�!�&�L�xha�_/)P�'�<퀊��[5�N4>�ڑA�-J-%�^�#)D� ��U�E���y�F�FLY�Ή;J�8��U��|"�e1d�ICE���f���C�2�0=�r#��I����q���?�"cނ�x����F�Ui�D�K�<A�(%H�b8�sfɍD��8�7a�N̓E�����R�7��A�t�0��2��L!c$�����8&�8B��4~Rq0�/�Ik�A�
��0d��!Ԇ@��D���O���3?��V(m
�c��)cx�q�H�<����i����3#�B@j*p��h��[Պ� s�,\O�����6P��C�����'Uf�x�'�mM�I჎�^�ƌ�D�0W�����/G�O#$Q�ȓ/����J�NfP�ءʴ�>	V(D1'������+�(����5� N���F�QD���"O��z0)�CEмK���H�n���a�(��P�䍺��)��<1��W.Av��ȅO)m�Rcni�<Y쎆��Hȡ�^[�H d��<y���ŀ%�!\OzY����B-�-�鋦��Z��'^0	H@��E��L�WK,{��zե�}4`H�$���yB&�:~��$�r?<a"c"݆�(O�eX�� 8 |"}:3�،-�8w!��!��$H��XL�<1Uj��� 1R�$�M�6i�ɦIBU��$GqO?7M��Xi���u/ɱ>�V�Y3��l!�d#<mB@��@�>+HMJ��!�D@��.�{!D�-���ռ�!�H�a��l��I�&�
b포4�!�D�9֔�����"X���RF���E4!�
�x�n�[EB�1�~1P�̃� !�Dg�9�ǝw�dђW��K�!�$�7|l�#�d��!� t�c�J!M�!��[IȰZs�	o�r([$
Z�b�!�d�DX��`�1L
�)�U	»�!�dU�R���Q�2�yį٧2	!�$ـ~j:`�9����k޾A�!�ϦK���R���ts�!����!�C�-��yv@H;]~̀�WL�o2!��U4̐Y�v,��`d�y9d��\3!�װz&bL�P*͈]�p�a �Q�O�!�d�z�l��� ��ŉR��,o�!�d��^��8�JƵi��8Q�[�!�/dw8!;�*#$$��T�K8m!�DCQ��1R�
\�d�M3���(L!��ę;S�7�ֵh���/�B	!�$�:P�M!}�h@�W/�!�I�z��`;ҤT������;_!�U]jИ��R-�d�0�gʪ|g!�I�7���0�I:4��x�e:C�!�Ě"�P�է�&6Q>|�pM�6c}!�� ��9s��;\X�PA�;-ȅ��"O@t`#B�@w���IU~�z��"O AgBµ0��a�ǥ��� �"OZ�xbB��	Ԗ���g�k��@!v"O*<!DEp��t9� �h�V"OQ�#�F*c�x2E�z�z]"O� �ǩТ,U����dΆ�u2�"O�A9�$ʜR��%�!!�c����"O,ā���N20��`�����f"O
���p胀�	9���B�"O,�j0���k�����n�#a�r��v"O���'
-��d��T�3���KO����`5�+�"�VΆ�������U)�@6���gQ4���L�*P�Y�)�E�PxL����O��j��[�W�-`Q葫<��i�ȓR
X�p�Դ~��`+_�<Q�'����#��\��O�>!��b!�*ype�j��T`w�<D��R���JФ�F"�E���8�M�k��D/q�@1��l�o�3��h#�B�-C4R�+B <�����U�
�ʣ�H�=}��!���![h1e�X�:`����?����cѝt��B��/P4D~�lP���̘P�a�����lG"}4��K 6PC�	�{��u����%C��ŰB8L	|�~� 1R$���ӧH���6�I)
*w�aP�"OTV�{�&)��@�Όx��=X(�2<�9��*���&>c�l��Ȉn�f�1c@1_��\9F(�O
	���x���RI
7~��`2h,Ԭ���)����?�4��&R��@�m�Mstkp�'^�X��E1��m˵��hM�p��D,͞1�D"O޵
#/E�e����1(ͯ8�nݲ���<ѓ#К^pqO>) n��4xp��/U�s��+`#?D�8�_(m����:jj,�w�9?
��	qJ�AC#�r���A��}�O�"A�s�̳���&Z�.-D�@�'A6!O�T���PeB�&����P�S�#� K�Ɋ�P,d{�oX�����f��#��*e�5zK��aT���dcR�!Y��� (�M���B�@��q�`��$i�&�2�_�z8 #d(>�Oh�Jf�L�"cU�BA˝d�'�p��
�k�2-��ٗ=�@�R9�~,�2�U[R��FŜ�Y��5��"O�8��̕INb4QQ�Ê{+�p���A��@�$�G��b�ľk h1t`���(��d��b��Yi�_�]=�������yBaАY�|�;c�^=�~��s@O^1��k�>0���3j�8:���O�x���$��E��X�t�ȃn�����{�{�h2�෡��@�@��
<#��2f�VS\U(0�G����b��a���(�\4��d�1@V���΀�6\�@EE���O��8��]6f��h�A��,zM����35��/5���ZV'_�tF1 u��d��B�O�)gq����	=�B Xm��+���?.��/�L̃��;!�=���~�V !D��*��#=,�ٟw���Ha+A0@9bmF6aSd���'D��Aլ9J09�@�LS���'�R��$R�@�ɗ;J�����%"��B2)˂6�����$���H�J�v�ҖGu��{R��.hu�@wm�!�f�0��ⲗ|"�ʐ�ų��$�mR`t�cɔ�)����֑� �'%ς���b���w^\lx�f �	���$P�O�2
��S�ˤ-��ԎMd���	���(���Џ�>Q¤ ���D��B�	�a}"���j����`�թ[�
ɓ�lB�q` @�v�
)�V�ڕ(�
�"D'��$i�������wo.ɒ� ʄ6�0!��
��I��'���j��C���Ή*d� �2k{��u�BÂ�g��=%�|�2��>`��!-|� �5�DtAU�=t0
Px�b�39�� *b�'���#��X\I���Ջ!JJP1�ki�by�� �S�䗽�����!$>�Rd)ғ<Ô�!VD�&-R�@���'}DA��I�#�<}��G��<�c�Z�d@��[.��t�:���1;Ѹ����ּF�h%°�mx�����Q�%ľ\�6d\R�Nj"�4}R-H��:����c2K����?ٸ6 9��@�aQ�n��@�j>D���Q-�/kl�EH�J�?�n	k�&�>i�#W��HL>E��<��H����\e(5�'�yb�F7kK��B7"YjV����5&Qzv(,,O� �Qj#l\�A�(�v!��h�c�"O>z�D�-��iJPa�$!׈H`"O���ԧ�� <>�#@�S���X��"O�q�C�֦D���jb�[�;�ց0�"O�\���՝*�-*fM\M.�(�E"O�< v��OXR%��Z{.YQ�"O�#�
�bX5�C!�%-Q�"O�< �@'O6l�"@%y�T��"Ob,��#6;R�H$�͉X̐$"O��:��Hx�n|+V�[:S��d��"O��(0%�#=��"�H�k�"O(C@O�3B� �VK��R�Z�j�"O�٨�D�-2���x�,äv�j��f"O��g�?�Q1��4/��0"O��B��$���;�����L��6"O$u�7��@\T��ႈ|�De+�"OXm	 aT9��JU!e�D�D"O���ӊ�H$z�j�	>��dp5"O��z��R�F��
�L��fl�"O�*��̺wP��Q_�s��r"O��j1Èغ$3Ǣ0~���b"OF)��@���Txc��42��)h"O���*U-�y[S�� ��"OT�(���u�8�ڦ�O'my�U��"O������#+}*��F���y|��"O�=0�`�,�*�*5 �he̸A�"Op���!ޖ9�@�*�-T#Oe�B"O0ٻ�O��l�(���]7��A�$"O�I(%�۔g"�x;��1��,��"Oh�b�_�l�A*��It
���"O|h�+��jǴl�d�
ZTlHyP"O�aQ���WȰ����eW:�ʱ"On�K���V�L�D��@i6 *2"O��Y%�E>0�nQiD�V���v"Oh����"�^�l)R�R�5"O\%��ǑU���㣉M�c��up�"O(�ˀ�ȤpKء��
�u���"OL�� ޿	~�hAh�{�z-b%"OD�0��P�&i;���::#n]C:O�up��S5$W�����S�Z�{��	���4�4M �Rc�q���R�ZC�ə���qG重#<��s�A$L�DC�f\��3㞜=۴�3ƞ�C�	D4p��'b�qQm��UזB䉟7޽3F�Oi���㦜�xnB�I�2��1P�g
5�z��V�g�$B�I� v��+�k180|(�d�!VL0C�I�V0��R�SЕkj��5@C�	�]�25��
�����,v�
C�	�(� i��Nph]�D�
�U/�C�I�_H�PkҿJ���(�ĉ W�C�ɖ.+�8�"e�2]G�0����*�C�b��`H7G�2=�L*�
2h:�B�Ɏ;\j�p�S* �@�DmH@�C�	f<x���Y;t@@|0��Ƥ3���D�Y}b�̾(�%�u�{i�U�`�R�ē8�Ш���8�)��=~,�aRe�G�7��A��i?e���s=��ѵ/*�)ҧ`G�@ ��6 ٮ��$�G�̽lZ���9���Ӝ
p��%�^#M�i��jC�	]ɡ'Yn��0|��mO�1�V�R��	!.S�0pci���'�\�$��>1�l�o�p��:E�����F��hO�O�8�&K\95f�����x�[�'���rl_�L%�0b�C q�ڍ��'�����K\�Ui�I"U��T�� �'�����Ɂy��q �ɟ�Q�%2��� ��B	K ��!`6�R��R1"O`�C��	���T�5.{X���"O���!V;s��
� Z�����"O� ���ñ^�8���BX���"Oe*����ݠtM˱}9^H�p"O}�D��lFٱua�;��ػ�'P�i��\d��xb� �Ȕ�'D�tC���-n2T�FF*m��}(	�'v��k�Ƒ� 2��D��:�}Q�'4� ɷ�H
P�IiC�Ւ+'���
�'#H���kR�>���We�?8ɸ<a�'W��P�Ϭbe|T��`�78���`�'Ph��jӟ��E���1��	�'�� +��֒6�Be�1�F "��H��'Ҡ8X!��Ow�|1�˗�
܌z
�'n�9��Up
*��+���4���'������ ��ؐ�W
m80H�'�@�4+��w�[	�� 	�'?�%qaH�"�ĲƤ�/�(��'Y:��HS�F���U$ 9l�$)	�'����	�8r�Ht�eAČ^�R�s�' ���u�,L�|;5������'��쉋�X95Ɯ,��9�'���څK�:�� ���W�Ys�'�NyjF�8 	���p�Z	��hc�'���	6�@](!��-�D��'ά8A�
OT�vիsO�t�����'�����j��[B�yBĕjkD|��'^t�g�������Gʠ[�N���'J��iEbֶI���˷�I0Qh��I�'��,Y���O;>LZ''��y�X
�'�68�c �*���	�FN�D�F|q�'Z�0���j�����k�.8�Jl�'�h�@Qz�H�ZǇ�1��Q�'���*�$���I
w�\;/��4�'+XPgJ
eI��+?")]b�'s����@�L*��n�f��'��0���f��=�!�7b�Ճ	�':�}
"��4lۘ��f�C���mR	�'���[F(�'z��X���M����'���Z�'L%�إ�L�lT�'�|�PJA$V0�1��I�T�l��'8����,��8�4D�Q�U X$D�
�'��TЃE.�8�[A�\Nw
��
�'�0��!���ddZ��Vf�	�'�ڄ"$�,����'D�C�4��'��d���2x���斡6���x
�'TTj��"V� �S�S ]�	�'>��S�߂5���0�bĹ{M��:	�'��們2S_Z	X�Β�py6�		�'Ơ�
2oZ�\੓̚�3���'�6�3),,��8󢍔%||�'Lp�S��Q�T�S�����y��'&$�t��2ȅB��]-�����'��)��X�;d�ㅯǠ}��Y�'fl�DΌ1ga\�zt�_ b�P�	�'�����KD�Z�Th��hZ�]82hB�'�d���G�B�Cd�ʿ@$�p�
�'�t���Ã�v�lD�3mĲAT�3	�'Ӵ���K	^���b�N�1�'H�Pe�
R���iE"��<I��'z.�3@.�=c�x�t` �
rq��'@��b3�K|�j5j�H�d�V���'☌��h@3V	��F��F0����� �܀ѯK�~���q�F>@tm	�"O���E_�x���v��;T�"O�	AE�/1j�=pp�?G5*2"OLzF��%#Tx2"jP�/�\؄"O mrU�K�;����Y�%�T{�"O^=��უ���B�X��Ţ$"Oz�Ң �7RZ2�y�a�D�`A"OX�Q�3(n�C����+�fM3�"O6}� �18����U.ìo��Tc�"OL�J̓�78��
�GY,sh��(�"O�����V~��	���Z� �""O-� �� �t�
���E�G�!�$Y:>�B!���M:dqe�b��V�!�D�C6^Ȋ.�9DH�� ����!��%~�A��aڟ*�a+"Ύ�8#!�DS&]XKBecr\��(�x�a����P�p��Q�O*>�l�5N�@�<QoZ�7)�е�U�D��e��b�<���x���B��^�Q�=둮O_�<�2�.J~	��O�rc�W�<ɷ��Gt����׆Dkv5��RO�<�Pe�*Q����Nɧ_��{�d�<�2I�5(���)���4���rBPc�<)իI�1ȅb ~��y!A�!!�#2h���M��*Ѐh��Ar!�d]�zV�i���b˼ajC��>
�!���$�����-�1�:̛���l�!�D#�=�s�4RQ1É�m�!�N�-��x�G
O���Â:�!�D��u� "hHz�ԘEݸ�!򄖗+��aC�̭#2СQ�[�7�!�$��Ny�n��C*��K�?y�!��xf!�C�,�H�K�O/8!��QKX1��ЧIgtQ{�I^6"!�$$3��p�$o�5Z���'�32!���H��-9�f�G[ �ǅ�+!�DM		"��U�@9Lb)�c��dH!��W+}2؂a�D.~D찻�㘹'�!��UO�dM���K7	*�5R��{�!�� ^(�*UJ%'<˱��4m!��Gkb-��eK*AA.�A�I,V!�$�'^�T�@�
�@:���S']8!�d��m��b�L�L7�%"��S(:!���< @�(֛T!�${cG�H5!�$G	��%vbT�nؕ@䁝�i-!�䙐P���ҶX�d�6FW8`!�$P�}����
�$@�b!��%!�)���+&+= �i�oM�e�!�H�DU�!b�.��|ﰵ��m�;,�!�d�d�j��?_ޖ�6L@�!�D?"3n�H����3ՖE�gj��p�!�;q�.�@�P�U�p�I�5v�!�WJ����Vc�:D[��!�!��lV|�3a�=?��f�79�!�6Wy�B�I�BԻr��<�!���&��!#��.t�mQ�`���!��%�*��7u��Ba�Y�7�!���^�Ӱ��aj`T�1�R�[�!���m�����6�`mrG��JN!�D@�P6�iy�j	7J����3+L!�DG�+ɼx8p��6t;~i�g��mE!�Tx"���M
G;��Hwi�%iU!�D�:�����֫.�ZUP�h��&n!�D�O�`[�n�
�A�f�B�c!�� ,��j�)����a".tV��"O����N�{���x��_�}f�}�"OΤS�,̰6�LPBA�L�$��"O�����T�8N�)҅ @�wB���R"O�e˃��~���ڇ��?��	2"OhУu�&M׌H�醰rȎ��5"O�Ր�ˀ�Z� U�� ����d"OD�J7�ڨ
�\:�F�i"OR-cP��s71jG$*� �HQ"O�L�!bN�Y��aGj��v��<B%"O��K�BГ3!~Mk�
�:B�p�Z�"O*��Tc��q'�@p���0��P�"O"p��CA��ZٳS�\�b��)�"O���+b\�T�ňB�_X��ɖ"O���b���*0ʈ*��Q&?��"Oz�!s��>I���p��	)E3�x�"O����Ĺ>:������>�-�U"O��"n�}� ��b*ǃj�
�"Ot\�W�ŝ��!�o�9a��G"Oҍ EHFt�ZT:��PIa"Oa���={�drElĂ7�:��"Oba��8j�Ό�!L�2jB���F"O"	Ju�d��,�#͊ANШi�"O����,R&N+�Y#U�NY6]˵"O�t1�+��aU��2T�D�b5���"OƍC�.�/O��X!g@$X-l�(d"O8�&m\�1�Q�U�.B��K�"Ol�ծپ?x����1L�Z8Ñ"O<d�p�O%؎ݫc�ȓ�T ے"O*�C'D�@%0R����!�	�"OPIJ#j�(*�ZsWA;?�6�*w"O��˷a嘬	Q�^[v���3"Oʉ�a�e��,�0J��|p����"O�ȅ�1 :�e�s��4yp�m�e"O
���E��U���HA 
��I "O�(؂ě"x� ���F	ޤ��"OZ�H�HR�Vxd �=��<�"O��࣋�m�6���OU.(�HY��"O�H� 	ղiLū��� 8pt	�"O�H����v�T�kF�0GkxS�"O�%�dB�5k�"�
�
�,=�1i�"O��*���o�I�c	¶tP�i�&"O� Jw��a���G�<Bx�"O��Q���Mx�L�$Gñ� Ӱ"O�%�PA�
2��@֥��5��9+g"OV�""��#㔐X���.9{��"�"O���	�y����0-
�'\�`t"O���dŊ0��i�4i��M��Q"OX��2F����T��"��<�"O1����k�q��,Y����q "O>J�P4"�\��˖�J���#"OLA�^�NĄ��@6�؈Q"O��� Tzl5�d��6�V�Z`"OLH7l�3n76�U�
ҕ�ybI̢@����B�A�TFީ�y�*J��1�Ƙ�R�)�/C��y��^�
V|���~V�e!�/��yr�J	F̎=a҅�y
�D��E_��yb��HK��ԁ�<s�x�jԃ�-�y��s�,�pEbV�k���!�g��yW�M!�]Q����4�3����yrDM��� �b��FN��yȟ9l�V�#(َt���3悗�y�oA)`df�U�_�k�P��r�ق�y
� �pbG�F�<� 3�̓wZ0��"Oܥb��4T�R�Y�F){G�|�R"OѢ��ҷe�ꀢ&ˁG�)T"Ov4�F�ˀ~ژ����G��)�"O���	   ��   �  l  �    �*  26  �A  M  �X  Od  �o  I{  9�  ��  +�  b�  ��  �  L�  ��  н  F�  ��  H�  ��  �  p�  ��  3�  v�  ��  
 �
 � � �  �) �/ "8 Q? �F M IS �Y Z  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" OTp�t%D��1k⭋�L���ctFR�<����� cE�+���+��N�<��+�7ƨS�g�s1V�85LL�<��C؇N�=Y���n R��@�<��(K> �H���"?�B����A�<Q�+٩$�2�*�%{F���**D�� P	"��)Ku�Z�5�&���+D�H��*�5s���i5.��en���(D����gR9&��J��F%�@ᆌ#D���3,�&���bf��*1b1駌.D��#�aիd�Y�(eot�zѧ>D��y��@~pH$�@���	3d2D��%%ǐGi*E�$�Vd4�;0�#�IB�����MN2D���8�HPd�<�;��"�d��M�0��l��,� GD���R���ƓiV�e�@N�(Z�b5�k�7i8)��	7r��#<�G�ω(�����<D���o�<���~�(\��`�4��y��Hj��x���ODZ�a�T9mVd��#�	c���'����$�O1ք{S+��(g恈�'�<��$m֟,z������8�[�'p*��)�E��lIb�I^0 �
�'[����ʊ#t��{�$] I&a
�'UDKfK�|���NP�FV>��	�'T%���ߔ*QD!��h>�A��'������6��^.�4�'��=��ZX�>U�`�lJ� �1�I�"|�']F�����?q�� B���8\�C�'��P�	�u��i+ M���� �'Z����ȑi��	�w-J�
��8�Y���|Re��y
�iB�L ~�B�[ `��yB�I�m��#�F���T���͸'������|� xQG�>g$eB�+�y�,g�$��U2`B&�A�%R��y���(#c���-F�,Hm�Tĝ�0?)O�Mi��O��xA3g.@!��3�"O� 
��u�^ڨ)�Č�"G:�4�q��`�O�m�%�9����Ù�J�m��'�*��/X�90��I��FmH)��'�4�Zr������l2l%zx��'�xa	�j�_��
_��x��'��1��ۃ�j��� ^#�"��˓1O@�DZ�-�j�(u�ƷVjf%���_%o�!��E��tK�Gc��A�+��џPP����C�v� ����x �%!&A^[!�DH�h���q�u��C"Vj�It���җX�nrݛ�K�}���"O� % H �:�LÕ}�"��Q"O*��s��s�~<;b*\�a��Pcd"O�\���A)=��4`�bZBI�`�"O���4���Y������J��Z`��"O���DB-+�|�f[b����6"O&�+ ���t�ܘ�/V?6{]��"O���V�L[��As���P�0#�"O"�R�C�`���� 7��UA�"O�DT�h%�9	�kBzTD��"ORv���L����	�ƋT�!򤌖���p#�6�QI����_!�D�-D�5	�cRxml�a1L�.,X!�DX�M��r�fԀ<d^��2��#!�ӵ=Ō(`#�;HO=�g�D�!�d��y���C`Hy��I\<C�!���-w26GD�EE8̣d�»<%!�� b�y@�I_�$�(S<!�D�:��8�ri� �Q�f���!�D	{A���j�X�iUQR!�D��������J���$!� ��0��3d0�#d�1Z�!�d�)h����wP%.J0�D �-,�!�dF	T��Yv�H���P��O&bp!�d[�r��3Uƀ'M��(�b�Ap!�J=��k��S�x!v�iY!�� �hm�qV`]�.C:��/w!�D3Q�����tM�]�S�Z�K!�=HP���h5w%�1h�"�}A!�$�Y:��9�Vtxb�*)�!�D�	*4��֎].9�[� �!�$Ocڄ[��D7����Av!��U䞌��K-3����"�- !�$T�,� 8��������+#��2�!�D��2q���Q�t>-ش�V .�!򄖥G^d�)GF�\A줂�
�.�!�$����"���_^� I^��!��O9�����o)pd-	�:�'$bL�'��� �I�kH.W�p�'zX�'P)Q��Y�S�1*;�}��'�(����a�XI	SC�v�Ҡ��'!�anE�`�U��B�A[2���'_������4);�����*���C�'A�A�@�P�.�����w�ܥ��'E2ͱ�%6��L[�T�3Ҥ��'i<]�c❡��%�K��	�'�ЌK�$�3�hh6E�{_`���'B��Q�Ë�L���n�5#�6���'ܵ����H��H��c�[hȻ�']�����ȃ
���Aԩ�4��'�J��"�"E��Hs�/ ��4��'��d��C��������  ���8�'���*�)�p�b]�E��!qh���'�|�Qw�X,X�� Lϧ{�(Q
��� ��[�H�>H�lu�c6L:R,�"OH���,��(��-°b~��5"O�PA�.��_�4�fc�����"O�A�⟅�ܵ����� $q3"On�3QG���L�7��<O��`���'F��'�R�'�2�'�"�'���'6��S�%�9XV�3à��3��<Bq�'<2�'�2�'���'8��'���'2��2��BU`H��N�A ����'b��'�R�'�r�'c��'*��'����U^wb�(�`E�r�^�pr�'�B�'B�'p��'aB�'���'�@�&"�0�� ���Hg(�U�']"�'�"�'���'���'m��'S~��v��K�qac� �"}ɩ��'��'��'�r�'��'wr�' �l(� w��`'ȟ-����q�'��'K��'�'�b�'���'�n��d�J/����	-PD-(�'/��'bB�'u��'���'*�'O�T�I���|#�F�| �  �'�"�'QB�'��'��'S��'���$��V�ԉ�5�U�h2�����'���'�2�'�b�'�'�B�'�p�i �=�(��&t���'?�'Zb�'���'�r�'��'1p�	��6����A��(�境�'���'oB�'_��'�"�'"�'�Fx��0Z�`�'u:�"䔇{G�'u��'G�'Tb�'�86M�O�dR-D��UC0��xIbi�r��~��Ж'��]�b>�MΛ��P���iUA�J���#SnłA��� �Oj\my��|Γ�?i$뜁HTH��O_��jg�Q��?!��O$f=:�4��q>uH����Ӷ)A�|���v!��!�!&�zc�$��ay�퓈2|-"s!Ч~!����Ɗ36n41ٴm�� �<��t�o��$�4ssWp��2�a���D�OJ��m}��� ��3��65O�Q���K:"zX�z�ś�hkDiR�3O��	+�?��f4��|��� 1hf*��������������"�D��m!S,扯iJ��d�D�z%HpU�H?1�J��?!2W���I��L̓��d��J>l�C�![��0b�k�z�����L�!�[n��b>M�1�'��h�I��h��W�4�P�����D'�@�'�I֟"~Γd��}A�l0��)����x��(͓3���K���N릙�?ͧ'tZ���	3_��B`�B�=e ͓�?����?���M��O"擙�b5��G.�$��7�	q)V-&**�O���|���?����?�Ψx�s*��h&&I�k�&���b.O��mZ<Qe�4������t�s�@�"i"U�����.?I�0��!S���Ĉɦ�(۴`P���O[T�rưi��ԛ�V����q����x�3�'�jQ9@H�=5]�0;���Ɛ'���*O���I	+v�T@��I+-èl��o�Or���O���O�i�<1��i�Ƶ���'�"� �> ��LR5.҄O�d���'��6m1�I���d榥�ݴI���Q�g���Ɂ��8\q�23��;p
|��i��䏂\f�P�N�#|��;��'q�_���6o�`X�EW�2~	�'0�'���'A2�'���#�����9�Ӫb� ]rB�O����Oj�o�J@�ڟ�ڴ���h��a�]��`��رs�H�@��|��'̛�Ot����i��	�شHP$W�9����C7yb`a�%F"MrO�@�	cy�O�R�'���Y7j��X�@�Y#�г�e�0"�'�剜�M�p�P5����O�ʧg�N�+!�2�[th���m��������H��=
�����|2��?��ð⟠7��) ��\�S��H�R@�� Ѓ���n~R�`��xX�M��+�<���{v|�T.��v�NTˆ��zL�����?���?�Ş��@Ϧ�i�hNH�
d/�bydl�*T��
�H�̟`�	:�Mk��>93�i�
�R��1�J���=*��re�`Ӥ�A|0�6M9?��Z{�n��/���PX�R�bޫ1TR<q��@�yRU�T�I�D�	ޟ��	ޟ@�O
��F��ǂ�@#�p<>��C�i�2 QG��On��O��l����睗	� ��c�/����$�{�x��ȟ�$�b>Ya�$��ϓ,(0�yF�σ!"`����	:6j��ΓfX<�2��O��kK>�*O�	�O(q�,����4�t�S�[�N*%�7�O����O�̛v/ '+�B�'<�$	%u�
�p�̔++ìI�5dOG�O���'�7��1��~y�A�%���p�����֬�	��D���]�K#1��Q���0��Q�m���S�hK� z�p�	��\���D�O:��O��D3ڧ�?��"J�70BA*W`ռ|��@唣�?�b�i�����'bFgӂ��]���X1�^����fB�>>���ʟxlZڟ$��!�����'l�������?A�B��	���)���n��(!��J5�'��i>���ܟ��	쟘�ɚxq��� n�#%�iAwj� |)ZI�'�6M��w���O`��1�)�Ot2Q��y  ��,��b�D%BB�c}JxӲ�m�)��Şq�Q��GO��̵��`���
x����\xܴ�'����'����iő|�W��qt�۔A���1와P�z���Eȟ�����<��e��4��Gy�|Ӭ�ʲ����@�x]|E�$&���`��OD�l�����d�<����M�Q��arv(яs�p���ʟu�֠�G�;�M{�O�E듶:��	2�S��� r(p@�ȍ2�Y�ǂ¯A]~a36O����O ���OZ���O��?6�ǐf��|A�#>��$ɆƎ����ӟ\3۴T��ͧ�?1��i��'1�:g���0|��!ľ"��2��'��I&�M�3���4b�<U�����ɜ:u�9d��1X�@���	�&M�-K��'��'�$���4�'+R�'�X˶�^��h�
'e)%�HI��'gR\�<#ڴp��a+���?���	
�x�.��D� �J3D�/w6�	����O�6�O��S�Ԉ��'���Ƅ_�kbd���dޠ\��Ap���&Mk��:�O�I�%�?Iuf,��$%����	Ȉ;^6�Z��̵-���D�O��D�O���ɠ<�f�i��H�A`�;/I�@7̕"B���d����'v~7!��3���ئ��c�¨>8���5@ܛo��Ԡ�L�M;ŷi��Bv�i���(>������O��'d$��r'_#K�5+�R�7<�̓���O��d�O����O����|��$�=Vd8c�FG5E������n�F���g���'X�����'��6=缾iQNה@[b�kЉp �dJ1��ۦ�ڴ�O�"��C�i��d� ߦTK�nU[��Aqc��_	��J�����&yP�Xx����O�N�?��I(Q���p� B-p9Jġ��@y��A�℅�����`L�5E�m�	�?�@\w$�!A�OX��'�R=pƠPr 	A�
�r���'�I۟�0�CQ�4�ݴ+�&�u����'�"�*&�$P�-�B�A������ء.W��c�.5�1�����9�J�$׸{�R`J��=4�AB��8>����OL�$�Of�2�'�?)��ϻʤ�׏��T�bY �$���?�`�i��Q��'��%a�>��)�ј�a��7=*D��� ��	��M�׶i�7-��6�.?� �8��G1|6�I"w���h@����jZ%��O>�-O�I�O8���O����O���J�b,�(��ư�1��g�<IշiF��D�',��'��O-B��C��@�q%�����X%K��?)����Şi��m;�AW1�~lH䮒p$CƝG`%�'�hI2�͟�J4�|rQ�D��F��BC�=��dl����4`MƟd�	ǟ�	��ry��s�`�âF�O��*�G[#�H� {���W��O�5l�S��$�I۟��	ݟ��Rm�:\�!�W�<��)���WPh�m�G~R�P=n�XG�$�wVtQ��n͠H~�� ���g�n�z�'�2�'���'JR�'b�҅O�R������B�2x�#�O�$�O`�lZ.:f���P�޴����$�� @.<��ěӢ��
~�p�x2�e�>,lz>�Bŉ�զ�'.-K� �(�Z�!w)R�u�x4b��9	��Ir��'�i>��ğ��I���D� �[B�����M��J��`�	��'(�7�v`\���O\�D�|�	�O�y�I��C>!�4L@A~bO�>��iD6m�S�)ҵ���o�@��.0BQ項�I2_KB�)ū�'�j����W����S�|����t/l�9#�.�|9����5U�B�'q��'F��dZ��۴U�FQ[�]�(A4ay��VoL��c_��?��M؛V�dDr}2�'�F�J�)�� g��	§Ǳ4+��S�'��ӇL����t�#*��8~�Ԝ~�w���J}��ě
!���4��<�,O��d�O���OR�d�O˧$�⦭A-�r���/��9Ӹi��T��'��'C�O�R�g��Ҡc�p�J?�-���A�8�*�d�OВO1���Ռg��找=P�k�'҉R/�p�T�l�ɰf)"� ��'
N1$�̔��T�']���Ӡ�����h�$�	��հ�'22�'q�]�pXߴ-I�0����?a�Z���Q!���4ls�qV\����>Q���?1K>�F��0�.4�G�T
U����P~2�J�:�7����O 8�	�y��)�
\`!r0���D��V'��y���'���'_���8�BJ�.'j��hM7��S�j����ش&ߐ����?�A�iM�O�N�1�1 ȥpMNu��B�y��$�Ц��ܴQܛ6��,[!�F����6ğ��t���p	������M[rP:��Ò|B]����	�t�I͟<J�6`@�e�B�$R�i��Wqyr~��p#A,�O��$�O������ s�0@ph%���p4LW�X��H�'+b�'�ɧ�O� ��1M�:�cV�O��mr�i+�	(1:�{��O6�O�˓8)�1b�`ץ(4T�k��� �p�`��?!��?���|�-O�toZ5N�Z��ɩ}.����m��x��%�����N��I7�M�B�>I���?i�3�D�zE�N� ����L
.Z�Mp�c�6�M�O�h�6!ͱ�(����5{�t��U�O�q7��{cN��	��d�O����O��D�ON�D%����p�q.S!L�Х�<�,���ǟ<����M�ff��|���~��֘|b�OEa���S��5N���@йt�'x����	�C�����Fћd�^� թ��!T��ᄜd��$8��<�'�?i��?	f�2v��%��ϑ�O��ٸ��4�?����$GΦ	�v(������`�OX� ć��h���4�P��<���O�q�'>7S����	4��O�<|�G�!9��á G�s{Z@��C�h�*!��;��4�fݢ�{��O��Ł��.�XT�V�C�t��E��OZ�$�O��d�O1��˓W��Fa߹%�1/�ʄ��C�!���X� �+%���'�v6�4�����Y��=��e5�*�s��պ
��@�`ѓ�M���iN9�7�i��	�,*�{W�O��g�? �"��T�[o��B�� �u�6ON��?���?)��?����)Q�MB�Tc)�+}02y"�eI<INN�o� /�"��'[�����'��7=�t��DI�'#2�)ī�'q��H�CG�)#�4�?�(O1��-��i��?z��Y&�X�n�REP���7H(扑eD�1��'2(%�8�����'W����Ď�v&&`���x�y��'h�'rS���4P�2� ��?���2��<P��^(q�	�C[�)�#��n�>Q��i��6��O��l�����f �U�����n��(�'��EG�֜<�э�D�Vݟ�ѕ�'��@��a�$x�
�%f�����'5��'�b�':�x�e�O��K����O���F	�0�N���O�O�Amڈ_�*��'��7=���O�nZ�0����
C�iu�s��Ōm��Φ�۴o��f���U�&;O���^0I�dȘ��:��`�i]�X�"VE
;(*f9QH/��<ͧ�?���?���?�q�Ǡ?�zt��Z,h�:�Zt�����꟤��+�O���O�)�V˧a$xb&\zQ���A�'$�I3�V�@�I٦��y~J~Rӄ	61ӀIЁ{��X���D'\ ��@_~beG�-�H���&>�'��	�4�`�ƞ�M���� ,�5q����	Ο<�I�,�i>��'��6m�|V��n$��FG����:%�]G��D֦��?ّT��	�@��?��(��)�w}Z�1���2�>�"v�����'D�������?I�}Z��]��I4��6=d5��-U).�tP��?y���?����?Q����OU�� O���Zq��e��Kᆄ0w�'�"�'t�7-��<��i�O��n�]�s2|��M�r��4ru��&��I$�4��Ɵ��=�"\o�p~B���DF����<T���I�M�0d�|�RET��Cu�|U��S����	ݟ� ���
���j�!��%�U�WOɟP�Ijy��w��%�d��OV�D�O�ʧi�-��AGa����/ک>���'7�꓎?�����S���a.��F�-z}�����#���˄v�>�"�O��N�?�E�/�đ�WG�sF��>��P!� �2�H�$�O ���O���i�<Ŷi����q����&J!7��X������Q�'nR�|Ә�p��O
�m=vx�y�	I
��t��&�0o@P�ٴ=��/.ݛ����q0ɍ��ė~�tnR:8���X��L�@���SN��<�+O �d�O�d�O��$�O��'W8M�@��g/@��1dE8r���inM��'9b�'�O8�hl��ٷ��)A%��:Vg��0/�*+/�uoZ1�M[�����)^2 � 7�s��ZE�:h�h�ȃF�&�m�4dc���6��=n�C�f�	Ay�O��Z�0}� K�e�")Fe!�n	�3b�'��'��	�M;�Gؔ�?!���?a���- ��+�F� ڢ�[Cb�<��'�j�`�V@qӊl'��@��;����
�&Ԭɑ�&(?iAD�h����!IO|�'e����M��?�&jF�ErT���Ӓ���T!��?)���?9���?����O���T �a3���e +k��+���O�ElZ)���I�d�ٴ���y�Ob�PZU�K�"���*��y2�'b�'+J�#u�it�		(���Og�Ik�E�� �+q'�� ��p���t��Uy�OqB�'��'���&(,��C��=�����P�}�6�M�1�ƍ�?Q��?�O~Z�8������sa%��4d�ذK&_������0'�b>����ɔt~H�ڱ��'���Y�('~��1KG�2?a��[�F���������DB�J���O��Uk�jQ�|4����O|���OP�4�0�A��+T�?��gD0�<�c�'Z���a�"�?I��id�O`��'�B�'0r��> Ra�E�u���3�(B�NHI�i<�I�g��V�OMq����W<�tP�q�{Հ pl�S=Ov���O����O"��O��?��F�ƬYE��
�lؔI2�Pb��Ο������4FO��ͧ�?q �i}�'p�rɏ�{�����ܚ(#z,HE'!�D������|z��C��M��O� �#��}�#�I�B����Q$N8�����7R��O���|b���?��OƚM�Ѫ
T�*0� �$v�����?q/O��lZ%̤�������Q�T�ռ>$V��`�//~Z�KԌ����d�^}��h�ʰn�ʟ�ҋ���!d ,�� �#t2�]�sÍ�A�AJ ��Y��O�)��f7����\p� )dϊ�_m���ω<Z�,����?���?��S�'���ͦ� �e��q��C����ܙ���r�q�	���Cش��'H2�`盦�ԫJ�Zs��4fP*��5s�N7mɦ1�Ŋ�˦U�'HhX����?��V�_]������VӚ�z�;O�˓�?��?���?Y���	T8q��E;���j��)�F4e�n�)i�P�I؟���i�؟4���{��<2�6@�p%uF��1�`B�'��Fu�8�%�b>���h�æ͓i#��X'�J�D�B�M�+h�\ϓw��5�D��O�عJ>�,O��O�`U�j���$ȍ/Cg2LX
�O,�D�O@��<��i
h$�'6B�'���i*ϓO1����BV�6y�Y����p}ho�"dmڊ��j���0�%?PۀU(�Ӟ%���'��� �Ҩ&��������꟤�Q�'?��(tK�B�̑D��&�����'/r�'"�'w�>��	�~9c��Ñ+,��b+Ʃpgz�I:�M[���?)��x3��4���%@_1����D�y63�;Ot���OP���\��6M6?I���Ê�3� �� �Ip� 1�RkW0J��B�8��<ͧ�?A��?���?9E�ˑF0 ���A#\f�iӢ��#��$N֦���i[֟����x%?��	2�4 ���� ��Ѓ����٩O�D�O�O1��u�х� 7Gx�2$gˋp,U��B	}�t6�>?�T�3$��IO��Gy�#�q��Kڸ{N��EF� 
h��'���'s�O�剘�M[aI��?1�.G�����"��X��ᱦ�Zn#�M��Rc�>��i��6m�����E�*-6��y���W�V�pb�"^��o�|~��¦il:d��Hܧ����n�-�|�A�_�4�R�hu�@�<����?����?y���?i����%}:��c�Q�`��C���'Y���'*�ds�.�6;�����9%���&��]�2�BT.B�_�p��.�ēj���!t��iK]�7-4?��C�Ȯ|*��إ:��sS��+\�����O�]�K>9)O���OF���O �CC�z䠑C�oP(8�^��b�O��D�<	��i���(�T�<��J�d�ߎ�b]�.�$$ yK�NQ���t}��'���|ʟ����Ż��Q#a
��������!��4��i>��C�'cDI%����g%x,�hi�(]�J+E�,��(�Iџ`��ӟb>�'��6����
�apN�GԼ���AJ���A
���Of�d��i�?�vZ�Ԉ�4j�2�)�@_f�	�$ś�Q\:0�!�i!6�Q���7M)?)��Hg��I9����7쨐4ş m�R���yBQ���	۟��I՟4����̔O�ٹE��?v,,� ���g�c���)��=B�'$���T�'��6=���C��.)�B�H��d�"������4�?q-O1��i�Э{�4�	N;浂�gS�� R�ŏh@�	*(�z�hV�'\Z�$�����d�'aP�%�T+ֲXA@�C3�y�t�'h�'�W��4DԮ$`��?��c��͊f�K$v�$���gƣ��9:���>�E�i��7m�O"�l6���T�^ a��㣤zqk�&?9�Z�w;�E�Ӣ`�'g8�����?����B#�uL�)`�|�*����?���?)��?�����O�\{P��4.���i֭��$�t'�O�a�$��)�O������?ͻLD-���B�&�**��9�KM�fnq������`�7m/?���*;���iҲ@_P�`u�.Ȟ ps%�!,D��L>a+O���O����O<�D�OX�*�ԟV��{��5r�ک��<9�iG����'k�'��Oj� ơs[8�Q�E�8� U@t"כ�B�:-��Mp�P�DVH�OS�Ag�� �А���/`"Y�s�T5���O4D�P��?�O#���<��̦Nô��P�G2an�q���� �?����?����?�'���ʦ-��I@П���"�H�(P�m�ip�!���]����4��'"��?��4�?��3m��Ӑ�E@�t% 7��9,$�{ܴ��$�]�.� �'ȸO��س|����V� S\�atMV��y�'�"�'��'>��	J%^���9_�T����ɾ3�es&�'�2�'��$L�����'6v7-:�dɝ0�x(5���K ���n���O����O��A-472?Ir�
r��2�c�Nsh �C�K�@�	�0G�O���L>�(O���OF�d�OJ9����+�(	Ml��-yb��OP�$�<Aװiߎ�Y�Z����s�4��(m����MY-wU�x`Q�����v}R�'�b�|ʟ�h���w,�qq6��(dh2���i�"b��i>y���'�fu'���G(.tj�t�o�7'�2H��\؟��	ğ8���b>E�'p7m�G�J	X4 ذ;�@��v��6X��p���O��Dۦ��?Y�W���I4K��݋�j˴(���0���'c!�E����$�Cڦ1�'�b��Js�'D����RIF�1>!���D���͓���O��d�O2��Oh�d�|��"�3C��a"�
�8�HU���m����L���'�R����'.�6=�8���.@�҈��lK�3��}�gD�Oz�$,��)��u�&7�~�T�e�0�z�h�/��lYM�6Is�T��Gv��D2�ĥ<�'�?A�탏6���ff*q��?����?����DC�=rE+�� �	, �mͬxf 87�&#1Qy7�B��v��ɴ�MS�i��O�� ͘�R����v,V�/K������S��X?<<�ʓ$�S�?4����,�f��0m�|���[2N���������	����	ʟ�%?%+Dџ$�	�x*vIX�NvX�=�b�A�>��I��Mc&���?��.����'m�I���]�\ߎ:����d��9j�+N�;5牉�M��i��n�W�v��j�
�:3�d��'�2��$KM�F:<a5&=Q��'�4����'32�'���'4��{���	кq� M\� ��e�2Q����4ix �-O��d;�I�OZp`3�ʃ1P�H�!�%@(U��RC}RabӸTn��Tj��	��LCP�䎟�b���A�f��m�A^��3
2�UpG�'���'�@�'���� E��^�N§<m
�E�$�' ��'�����W�r�4H^�p�g�m26"��C��ȵwj`z��9қ��D�p}��'o��'�ҹ��\�PȎ��&[=i�Beɴ�SJ����P� �0t����i��Q
��Z����vL�|�j!p7O����Or���O����O:�?�8pg� ÖDi��W�ps ȴ�ʟ�Iן�;�4T�̧�?Aǿi��'�4th�������C͛�+R�|x�|�'��O��D���i��!MZ� h�S�͋?�&-�$J�4i�BX1b���?�SO2��<ͧ�?����?�CB?
"K�눜5��ۭ�?��������j���ğd��ٟ�O��ep���'j��}�����Od��'k��',ɧ��&)r*p��lX2�����ϒ_�a G�>�8%�є��2/y���U��-�X�K���J��32ʞ�U�������������)�cy�	k�Z�s��
�|�%�E����Ǧ��zܶ���O>�np���I��`�fFX�yT��ˣ$�y���rƟ��I�)�nP~c��~��$�}�䊈�SQ�Am�}[�/�<1(O���Op��O���O�'����f�}@4�X���7�,1�i�� ���'���'	�O��	��?����APJ��ĩ����/�j�oZ#�M3��x��tƖ��F0O�x�b��1V�����4U��� ;O#d�ˉ�?�S%8��<�'�?�e�؝0*p+A�^�j�"��Q��?���?i���ăݟ�E�<���F@�qcl��fhp�c4P�0�T���T}�xӒLn��ēVy��"�ۼw 0�V�A����'�@��*C�L]k��ןk��'֜���N;c+}��F�4'?����'X2�'[r�'��>Q������Gʋ�|�!3�z`�X�I:�M{�܏�?��� ���4�<J�ܷ;?��J�4l�%C�6O�to	�M���	D �ߴ���K�?m�)s�'q�(r� ��~@؆c^7l2ȸC+�$�<�'�?I��?y��?Q@��l�H=1�Oo���'�������;#������I�<%?���S)j�[` �qH6d�f��=K:�(�-O��z���d9?%?U+#*���h�Hӣ��(�R���mY�z�D�{`�0?Qc	�2(���!����Z�s��C��8O E�\H�@0���?���?	��|�-O�]lZ:b]"H�ɼ�na ��ތ�(��E�8���I��M��� �>�ֻi8�6��O���ɞ|Zd�� �T�kM�n�R6M=?IP���'�J�	<��ߩ*aMV�S�r`��eۙG�R�h{����ß���䟜����T��KI�Y��ӄM�0cҰ@��.�?����?a׵i��۝O�2"y�ГO^	ېه"�z[��س�˩g�N�O���O�Ɋ_>7� ?q%�F
zGH�b�B7Vs޴��`�8X�P%�g䴟�&�엧���'���'�F���KCX �yE��┴!��'��T�0cش Tf@C��?����N�BԎ,�Z4�xh��ϡP_�I����Oh��)��?�r�kƔp��4CC��Cv��=Ir��4C�r?T7�3?ͧ8S���J��?����УQ6&Q)�Ө/�6��	ܟ8�����)�vy�gӘ�a���Y�ȑs�ԬRu�-���;M����O(�n�v��V��	Οԃ��h�Xˣ�H�	T�X��Aݟ8��+���mZz~�@��3���}�q׏Q�f�3C�>��@��l��<9-O��$�OR���O����O��'z
��sJ�z�(1���ߐ1�6Mc��i��e�s�'2��' �O3��~�󎏱V���O0pyUxЭ^>.�8�d�O�O1����E�s����G�L�FG؟>�,,[h��#&�	�hZ���s�O6�O���|��P��y��_���Q�N�r�������?���?�/O�]m�!D*p������	� p�@�Ą�� ��EG(�q�?��Y����ܟ &������2�8h#E�b9� � .(?�F̏(�ڈPߴ��O[ ����?i�#�W�(Y8פR�.	�7���?����?���?�����O��`�X*���Ai���#�OԽo�6xc*A�������4���y	��s����$��E�Q	G��?�y��'�B�'mM���iW�I!Dz��b�ߟd�����'U2H���U_њ�A�k6��<ͧ�?���?���?a��6J
�@	J������Č����&d]؟��	�<%?����Tmi⭙6n��:gO�/S�*�O4�l�M�u�x��D$��rq�殛_P��{��W_���*�!�9���W�`��M��ypޓO��e^���Æ��L	�E�D�q{�����?Q���?Q��|�/O	n�y�V �ɨ|HF�cuo�4B��@��F<%�&��ɑ�M��⏵>����?1��I��q(ǩ�$�����ݝAР�;��F�M�OA$�>����d�w(^�A2��b���[夋�])�,��'�r�'"�'b��'�����sB'�r��,�6�$�TA�O8���OZ�lZ�a�(�S� �ܴ��oK��0�����Te�'$�HH�N>���?�'?�Q	۴����
"T�s�'�r/��(!�����5"��p����r�oy�O���'��,Ț �^iH�G�`A��c�~���'��I��M��l��?I���?�)�ڍ{h˒3"8*��[�do�Y嗟���O���O��O�S�?��`J����2�x��&�
�wϔ��cm?0(�m(3�1?ͧuaZ�$���U�D0�E\B���Yc��s��p���?	���?!�Ş��P����'� Z!�%�	NA���04ꐦq1@ �	�0�ܴ��'5�=�V�H��]��j��#�����;9��6-��I
�ƦI�'����K��?U��\\!�`��,�h��b <��J0;O��?���?i���?9���@$#�\I�(�;�XU#1"�?n�T\o�h� ��I����A�� y������i���5J�Hׄ�h�#?9�b�i�D�O�O�K¿iL�� �19G��˼���@/UҐ#�1O \`�L؝�?��-��<�'�?�aO�j�Nđ�տI�qP��W�?����?����d��͹��_vy��'�䣢��=[Z$j��Аr����Dj}��v�v�lZ蟌�'�v�2`����,�Z��޸�O>}�2��8	 ��!��ϝ�?q!c�O��ґ�օ�����(�3@��Ă��OX���O&�D�O�}b��:*���B��;�Ҭ���ӑzO�L(��8�f�u\B�'�v6/�i�%zRȇ�?�峆�:\?PX�6N����I����I����o�c~W�t���'�V�:`�߭�T`���,�f�|�[���� �I�\�������5S]FqE�ׂz�����+�yy�}������O����O�����D�%�{l�"ZQ�)ZD����V��'��e��6��D�K�OX�p�@/P�Dj�H�o= �'&h'X	�&'?i��,_�B��N����ε_Yv0��&g�-I�J����O��D�OL�4��n�fÔ�r���62��`��("���D���Rjm��pЫO���O��RT8�3��e;ƈɢ�J�|kP�:%m�:�*9R�!De���>U��6[����E�dd仃�'K�v����I����d�IO�'h�H�s�4W�d	���Dh|���?����K�����'�7�&�dU�WlV=��	M)^� 9��^9�^�O����O�)ϣ��7M.?IU�� gL-0�a�%�Z,&�	s&Z�
p��������4���d�OD�D�/!&�`aJ�n��  �D�OAF�$�O˓_����"�'�R>1c��W0����I�'ʰa��+?��\���	۟t%���jX	t��#b���[���5I�&�8�����A�E��P~�O3J��!��'�����J�?��)b�& 4��Z��'�r�'	����O-�	5�MT%s�b�I�e�:R~݉c��]�ru!��?	4�iy�OpH�'���Тy�R�� E�v+���0J�'�DQ�i��ɤ�Tq�e�O��'�)�&�67i����A�l�����Ov���O����OJ�d�|�7���k�")�dH�Z�|x�Aͽl5�Ҳ�?���?��'��-���4�@*N�N\D ���Ѽ@݀U9F����۴�?y,O������D �T�r7�t��
��ѳr������ҝls�H�Re�(+�iۑ_[���d�Py�O��bZ��\��DL�
��ъ�<
b�'hB�'��	��M��E&�?i��?#�"&�y
���<M�=K1�̂��'����?	���CH���#/��nd~�c@��!5�'�ȼR'N�M���$ş0�g�'f"��a�ەf�؊�M 
D�����'L��'��'L�>���[&���g��0�=[�=4l.��	��M�� ���?���M��6�4�\m[��N���o_�	c )�:O��mڱ�M���i���"V�i���>D��X��O_��H�L�
����T"eF�d`�F�L��My�OU��'y"�'}�D� -���`֔>Ϭ9�E),b�	��M�T�@��?!���?AH~*��`�Y�� "
_ ��&퇗Q�^���P����4=Лv
6���^-Gk��fkG�c�	F R+D$�Ae�I��8��'��$�0�'h����"��_�]��m�>a���2�'`R�'�B���W��*�46�B\Q�x���S��ƺ/��a�%�N�<ˬ0�������D�cy�'ɛ��'���;�
E���qf� �ֈ� ��O<����$ZCc*&��4�	����V�$^�)$+�%�4��3O<���O���OB��O��?�- %i�&  " 	��!*�-��L�	ß��4H*��'�?�U�i>�'|*�ã��pi�ïԨa��	���2��5h��|*-���M;�O�T"`��4'^�0�A��5[��T*Q��I3��Df�O���|���?9�b<�0E�X�g0	�c�My��s�)��?�)Oj�l��tll�'#��O.wBP�k�~�@S	����(Pv�M��y��'Jʓ�?�4�?Y�O�T�O�����%>5�N�W�Xi0���8SƬj��5������i��f���O\qr"��V8\�y+J7�țc��O>���O\�d�O�)�|�(O ioZ6z����1��T��@B�#gԅ��[ʟT�I�ML>ͧB��	䦽��ί~O�Ɇ͈-H��h2ߛ�M���_�n��4�y��'��e1DD��?E��O8e�AK��0�1E�nh��E1O�ʓ�?I��?����?���ή;=jl*'��#Rٰ	�$�?b���oZ��Fy�	��H��\�S���k���C�)��_�j��&�P-Y�:��7 H+�?����S�'!�D�ڴ�yb��*�$�\��:M�p*ۭ�y�N�$	����I��'��i>��(@��Ȓ�R%J���+5l�HJn��I��|�I�4�'�(6m�8@�|���O[n�a�(ʔi�-)�X;B� %t��?)�U������x'�tq�F�a�A�L�*��y��h7?���{��(�ݴ��O�>A��?iì��Wu�� ���h�R�jL�?A���?q���?Q����O�(�
�-[�6劰ƦZ��VO�O^�oڄt������4���yG���]�:H�@G[�R�	��Ǐ�y��c�haoǟ��A+��-�'R���G�?��ue�[԰�1���b�X*�iV�'g�i>��	��0�	����(��� ���$Ϟ[Nŕ',�6킜x����OD�� ���O`1r��ãF�$ ���MZ��S'Ag}��'��|������� ����+K-��y�QfԊqD��U%��;�I���h�
Ժk��'��	��}�P0�є7r 6 ړh;�;uj�O������8�rAl,X����O��	Yº�$���K%��T��d�1`�����+�
���?1(O��$ Af����MC�4ӿ�,LR��8�#Ś�����@hT��4�y��'�D��g��?1q�O��I��f��Q�C-O��V�]T�Y�2O:�$�OV���OX�d�O��?]�ş"-$�A�.�)���C�Dş���ߟ��4j���̧�?Y��i��'&�1�V���WFލ��@A���9!�|��'-�O�R�qƽi��		h�I��M-D��*��G�x���0�e� +D��n�ay�O�2�'����^�4}A���)*I���EG�e���'����MkD

��?A���?�*�Zuy�`�-*�l�k�#�3X'��c1��<b�O���On�O�ӋH�A �����Eƫ\'l���< hͲa�)?�'p(��Ó��c�pB0g(z(!Uk]������?����?��S�'��]ӦE�i��W�)�׎B�'�jl���G�E�$%�	L�ڴ��'�ꓶ?�C��F�;���O�p�EG �?��>\8�ش��d��д)��,�Vh��j���7��ub�	��O�]6 ݮ�f���X"��9��i�z?�*��= �ԕ�
��S�^�Ag�L�D�ڨ�U�޷K�*蹑f֮hZ$(*��Uiԙ{�kēZ)
W��d��\�9�I�[~�����]ڳ�]�J�Αj�āef��POӠ7��5h�|d8�� ��l�2�Z�V��1*�Ē��jWdFc��$����m��x��M�|Q^dѦ.J�b}x)��̈́=��$*�fCw���J��q*�<8C�H�&���3�0U��`�W�M����
.;67M�O����O�	f��L�"]�� �[~�H�Z��i/�a���S㟐g�ޜ(�J8�S'" ��xg)���M���?Y�Yl�a�c�x��'2��O~e�s�V&��ٓ��xG�M��^n�1O����O��Ή'��i	�b�ib���d�;]��)mZ��L��h����?�������l�ml���!
)!���C�#�I}�J��'L��'c2U��n�-��$z&�V�t9B̒�F"��)�J<����?QM>�-O��V T�.dQQ��[���g-]rM1O��D�O0�Ģ<�C�յ �N��n@ɘ��YkB���R�	�l�I[�Iky� �����jx���Cg���9�.j��	۟��IğT�'��Y4�n�����3|~�� `��*�Vm���'���'r��}B H	lg�XC�̎����Ĥ_��M���?�*O�TA��v�؟��Sl��b6iId�)� #�).ij,�4��d�<�E�z��O�iR,�'�Z�ެ�q� �{/�R�4�򄕴#��oZ-��I�O��Ɂ}~� ؒn�lH�b�O�E셀�	�'�MS*OZP�A�)��}�v�[BɈ�G�,L���d87��QJ�m� �	؟��� �ē�?���B���R�X�L��&��'~���cD�O>u�I !9�=�T��7V�t�E%ـ,�z|��4�?���?Y$ �~�O�䦟;b=@�r��6K� ��0ţ(�I�s�>c���	� �I�=*̸��D�&�8Q ri
�j�#�4�?��$]'nC�'/"�'�ɧ5�� Q�xY�BB� ;�Q�XQ�n�@����<	���?�����DA�=�4ȡ1/��:W�w+ qۨ=� KZ\����P��|�@y�"�b��!ԭ�#XT�Q­���¹R�y��'�"�'��	� �<x�O�5#�K1�}"�_2��4����O��Ox���O|$#�M������$8H!���˞� ���>A���?���� 3Ѥp�Oz���OZl���DT�i���{�h��1Ū6m�OҒO��D�O\���2�I'C$~��R�0 ˼���N1}@7��OF�D�<iD`�!f<����I�?������es�.��#�z<pD��ē�?q��h�
y��՟H4!�MX�R��j�B�3k��ї�i�I�D,��B�4�?	��?��'?k�i�Պe��� ۆ�C�$��� Hg�n�$�O�����FܧP�*E�D��"��u���8��@mZ�Z��4�ش�?����?)��B�	myB*B'@%xc�� 4�� r�R�d6&|1������Hq"���E.�W垛4�\)8��i��'����o�����O��ɦ>F�T��
����[fB�o^�6-�$U��	=�]�J|:���?��#m쨑С3t �m3.S���x���i���=mn����$�O�ʓ�?��'�\��!����w��3�||�',(t	��'8a�':R�'�S�(�uX�`m���-E*N��5�2�C�y���OX��?�L>a���?�&�P�}�z�j��͐����Rc���)�O>��?A���DR�frđ�'$ XA�MW�>���� ���9oZAy�'��'��'������On!�u���m���aD$H`�Q���������Wy�a�;Ԋꧭ?�u�V�gn�Lq7��'Lu�/��C���'��'���'������$Αb@��Ť �1��]�	���'�"R����H����O��d���M��A9:ĸ@H��;w�C�ECD�	ן��I�y,9�?��OEF�{5,�e40;� Y�`��!��4���ɂoZ̟��I����S������ڄC����SG��_�Ɲ�гi�b�'��f�'��K�O��>�z�eΨ�&��eK�U�,8��q�Z]k�Ħ�����I�?}��O��6s� ��0�#w0�c�d��Lܚ��i�B0f�'�d1��O��?���_v���j�aq���6SH��j۴�?I���?I�̀�,n�����'Z�DZ>Pg(�lO{`8A�ܔmW���'�'����<���?���Pg�"F�%fT`�F�*���a��iPR�M�
�O��O�O����֒C}�7�/[�qe�3���?qK>�����O,$Pӂ��0�{1��ꁢB�,jʓ�?�����'���O�4X�)ɹ��2��.��LX��iT��y��'x��џ�{�A�J�$ϕ�k�� @���;@ޘ�r��֦��Iџ�?!���d�$�נpGJ}���; Mxѣ��U���?�.O���Fu�˧�?aNܘK|�0�t �'��17-�9tЛf�$�O��a�&�0� ��D�`��
�.`lU��m}�h��<	��?��Q�/�`���O>���d,8�H'tB8���+����W�x�'5�	�X��"<��9���)C��a��=��M�M�x��'�!l�"�'g��?)��u��g+DY&ŭu;�=Ӓ�0�M[��?A��E-�L��<�~A
�9Ox h&�Ļa�a�,NɦepϪ�MC���?������x�O9́�b$ުD���V��;)��ؑƪd�:EA�O���<)J~�'⽪1�C��K�/S 4"B�gӎ��O�d�lE
�S�$�>�CjW�3�`0A�����n�#��.G[1Or$R�G\Q�ş�I���ʒ�Ѳ3���RA�W�:5��J˅�MS�H�	�֚x�O��|ZwX��*�k�\C���9	7�<{�O$��Od��?)��?�)O,��Fc"p,���C�-P0��۵ �4V,&���	쟠$���'�Tx"#h�T�IB���:F��) �!��W��I֟@�	^yb斦���W�0�8M��H�F!�T�ӵz,���?������D�7��t')��E8\
 ���"Ğc�,��'`�'grQ�AeD���'DJr9jcf2Xq�Da��[;Ph�a�i-2[�D��My¯]��ғ~"�d��`�4� ��V�%C0qAe����	��Ж'�i`��,�I�O���ƜT2C� \�0)�� V�Jndht�xb_���QdҟT&?9�'Q�V�)c���Vw����m���`�T�n��t�4�ij꧃?���=`�I.��ԑ�[�
+��S�O)_�7ͽ<`���?��������4��ٻ$NA
]��a�c0�(amZ4_i��S�4�?���?���)����^=�0H�pLW�o�D{��	|*�7���s0���O<˓���<���jd�b���S���@���0���in��'�뒱YV���D�O��	.B^��!�����f��$8{�6�+��Gy5�?Q��ٟ\�ɗ6����T5QB�����,Edhcش�?I������ty��'
������
*�2����Y�N8" �^$�	*��ϓ�?)��?A���?!(O"�����+"�v8d���'��8 �]?sξ��'�I�0�'b�'���$ �i����	�0�b �$ē�'���'��'��_��E3���$�yw�����J��������M�+O���<����?���u$��'��U�g"<8�5�Ee� 4��4�?I��?�����3�J��O�Zc�.5��X>RΈz�M�d��h �4�?Q/O�d�OZ��$_C�D1}B/�&kVU;���
�z��EA��M���?Y)O2TQg�S�4�'���O[����lŹ'���#�&���
v��>����?i�z�a����?a�6f��W���9v/[)bx�Y4�q�����;�i ��'���O_��Ӻ�IV(V咡��M��[u����	򟨹�h���I�ܸ��a�'L:2���	x���:��A9>Z�yl�a�|9�4�?9��?��S$��Cyb��~�D�fk��d &㏊=��7M���d�Of���O��JT�^�.�
�|	�����?�7��OP��O �1��P|}Z���	e?	W�k&�����{P�|d���&�K��m���?���?1��Хj!�}��-�	O�=ȃH�tӛF�'a�d3��>/O �d�<���5#R/�(-j�W
`�qI�Gr}"H˺�y"�'���'���'��I�&h�]���p^�K��<�Xcߛ���<����$�O����O���*T�1��dA��;�N8t��:#���OR���Of�$�O�ʓ{>�Yh�>��jrO�az��1oP�}���iE�IП��'D2�'@bNM��y��l�^!�fA���'��Q(7��O��D�O$�ģ<�NȠ,���ş���a(��L�Ht~4a��L��M3����OH���O�K�=O��'����/	i,ΈA���._���4�?)�����4{���Ok��'����*.����ǃTf(PZB�Q�C\�듞?9���?����<������?��ciۘ<��Y���ߔu�T�Rf�y�.˓c�����i���'�r�O�T�Ӻ��`��[E�"0�� �X�Zu���	��០���v���'y��cq��K�Sf:�#��r��q�FG�uD���[�v�~6��O��D�O��	 O}"]�p2C��CNpAC&)S�T+M�aJ��M� �<���?�Tlɠ��OX����s,��3Qo�y�cR8\N6��O����O�Ȁ�I}W����m?���^�*ђ��(a|����Ȧ��	ey��&�yʟ����O���^C� "�.���!±o�0�<�oןd��O������<������Ok� L�� ݜ`�r��3�ڟ&G��F_���u@c�<������T��Sy� ){�j$҃�!'=�RU拥5N��w��>�)O^���<���?q�xi�E �,�v���i��D,Q�L��F��<)��?!S;�?I���QW�ͧqr|���Vmƴ� �d�
���o�My��'P��͟����0Zs*}����X�Mۺ�a����q��厴����rH����O�˓Ur%�����`<!m>$賆+Q7z)i�,��0�6��O��Ob���OxuRw��O��'20+eg�+e 0x���A{
ŀ۴�?	����@-H�&>�	�?q+U��1a�*H�U�J�Ks�%�ē�?� �v�̓�������zZ4� �F�Z7b��,��M�+O��RK�Ԧ�������A�'���\�Na�,�t.[���L�ݴ�?!��,x�Fx��	[ #����#C��Rz��4!UY��6g�9�b6M�O���OF�I�L����ĀYL>�p����3��Q�7O�?�MK��޶�?�O>�����'G0�
5��6�-��m��T�j�����O��ۡ�ZY%���I���_d��PgA�)�V�2������io�R� ���)r���?�&<f8+�!��$L<}��#зʡ���i����0/"zb����L�i�M.�z�;�ٔ.3@���n@�� �7��������OX���O�˓`�f0�FY�K�&�d�ѓR���� Om�'���'��'���'�h+R-��-� ���+�'jt`9[`�����Z���I�'?�5I����� H'3��qԩZf��%�1�ē�?�-O8�d�O��$ոc;�S�G��	DGtTXM��Gr���?i���?�+Oȝ��k�S7s'���1�W4R�
y� GQr޴�?N>���?�����?L�|��%�,:DRرR���<0"�r�����O(�r4}�%����'���$��+�a�1ǜ�v1�X���-Mp�O`���O��T2O�O��SY�m�� b�a!���"U��6��<��C�+���~"���z՞�����A�>�j���/8E����}Ӛ���O2��'��O��O��>��,7`�L�i��ӿvo�	�2%}�P��lL馭��۟H��?m2�}�,ǀ- H���M$��dS��xZ�7�L� ���d1�$$�Sןx ��o����5!أ85r|Qu �
�M����?Y�'�Ą�v�x��'>2�Oj�J���(��m[Dc
��cC�i��'�с׆*��O���OP=��L�T��� ��J^(hs�릁�ɔ}O�}�H<�'�(O��1�H���$�I�&�- �\8q[�4�!̈Ɵ �'��'
�T��I"�^�a¨�eF�$�P�ʳ<�53H<	��hO�$ӕ(yP!(0P#s=@����´��4�"��O.˓�?y���?�,O�MXɖ�|_2P�"BE�:>Z��r`η&N$듑?�����Op�����O ��NS���ʣh����P�Rb}��'��'�剒]���bL|����K`n�rs(�"'�-)��!J�v�'NBT��'�z�R̟�	4H�J��҉	_,#��U�b6��Oz�ī<qЄS�(��O>b�O�J�j�TH~��2��42M���f�e��˓��DC�X��3?�禹JGm
6EX���Z�5{�-���pӪ�S�Z���iI
�'�?q�����^��D�z�6����).�6m�<!4�ׂ����L<���l�h�V��]"�]�f�֦����ͳ�M;���?	��:��x"�'���Af�ʃx��@�Qb��3�^T�A eӴb%�3�i>c�4�I����#���s�&��t���j�a�ði7"�'�넥ld�y��'t��X�:ݜHaG���R�.W5�t�DxRI*�I�O
���O�t#dͫ	�.��������s�.�Ц���W\���O��O�B�'F�m#R��Y2f��z�F�3=�$� %������(��ğ��I8G�L�����Xn����-�0��W�Tş8�	hy��'�'���O�9"���"��Xtg�yC`��i[��O���O ���<1�ݎ-���87�@*TɌ�MW�+�"K9	ڛfV����Eyr�'���'��(��'a�Yx�AH |�Ij��I�y��mx�6���O��D�O��V�1�T?a�i��[��\UY����F�")8C'v���Ĩ<����?��6�|u̓��iCZEH�O{b J�"�80P@��4�?�����Dӱ]���O���'J� ��2�����ѿV�h�q0O�A$ꓴ?��?��<i+���?�#@)پm�r%��_��P
����˓n��b��i��'���OԲ�Ӻ�7��^��W�#���JA������0R�
p�4;�����.��S��1
�Jݴj��q�խ3V�7�9i��o��`��՟��?���<�dͅ�9�p�B�Yu��8�"�3xțf�[��y�|�)�OhXДˁs�
���ح(�����F���I��	�Ir4ӮO
˓�?��'�P�n !ľ]�D���j���q�4�?	,Oʔ�`9O�'s��xಆ]\�䐀1�T�7��ј@d������\�͇8fHB0���ʸ$b���?{�0��I�.���/ޠ�H���i��A��A��5"pꤋҠÆ$S^L�Q�#f��C$H�>!b<�rdǣi�q�#(Z�JP�Ȝ;���ҁ�)R���fT5.�N�)gTS0�;����uV>�C�Ɂ�D^�p��;=&9�'�W"P�����_�;1�Q���|m@�ivl��P�h!�R�f"���O�Ժ�.�O
��d>�5K��Lͮi���0V"�lɗ� ��Xy@Y	C�\t�\e���O�|k�,�b��d�q#�0[6��Tbp�S1\��>x+�ǈZ��i6�ۧ'cE�?��d�ꟴ�	]yL�Ƹ��_0�*,��C�ј'��{�ʖ��,Ii�"�,�f�i�m��x"%iӄ���ā�`�``gW)D���2O.�>�*�TV���IM�$���Rr��'$�ј%像b��AAR3
�B�'B�D�@Ѫz��"�+*T�T>U�O���VJۧf�ya����w�EQO�h���N04�#�� ���F����!1���`�# ��M"�����	�F ���OT�}��,�	���=��
T�F&Q@x���-v^�:�! ,+�@* E��HJ̅�	>�HO�$�g�׹ 6v���7/i�3��Hr}��':�T-%p0��'3��'��wpT�CG%�&�n��nʞ��u�I6P1���2�OP�3��!q1��'Ƥ�$d9\���2�D�bF@���@2l'4 �FI�O��+��������?�-��o��Ym�m�ƥ˨����O�󓭵u���$�	�c�q��'Z�?S�yz��N1t^"B�s�f�*��KY�bI8�MS��eM���'��D�0BTxI�:n��\��٭�|�`�e� ����O���OFT���?���g��\L=Z��
�:��	�f��iBR�6��+B�������[!�y2'�6U�(ظ�O�p��������L���d���W��y�,��4��l�@C! m)7GHN�V,s���?a��D%�I�s�2�b����)
�	s��g��B�	�8H4# �@�O�"mZ'/$�c����O�˓.���Q�ir�'��\�B90�����ߞ]܈`�S�'9��?��'��"ҡ�l���ߖy�JЃ��e����fą$�X�`2	@Y��LJ�']P�Z�Ŭ)r���0˘�"/:8 �*e���!Z�/�I
�)Uu�!
���L9~;r�'A�7-�O��rg;W z\0�)Ω��]��h�<����?	N>E�A��cdt�0#nR�wq�\cĎX���<�S�'	�f���=��fR�q�r�׷+6m�OEnZ�e�"˅�O���OT�ɖ�W"�d�� �ܼ8S�6H�N��,Z�+"\���O�-�'
��v�~}��fٙ6�� ��|�.�"�bŨ��/χ[Դ 8F�ݶ��
>�v�`snˢ}k�]Vn�^�O�(ybC �|ZV��@;*Jjd�M����k�O��$>�'�?a��~T�)Ѱf�/,�(\�C�\��xr��%XL��aS�!�f���$��0<9��	�qf�b�ٞ4�r0s�2;G�8��O��$�O
A�s��'D3x�$�OX���O��w�0���@ߦ_0r�iT�B�k��(y֮,f(�����.�.|1��'�B��Wʆ!<��|�!�M;=\�E���&Z����@-�O|8B0�T����nSl���(!�Mg�\�>f�x���$ܹd|�O+����4ha�E��
?�d5�s�:o!�ā4�,�%��)D�|��Lk���O�aEzʟ�2�fJs�À%�bx�2H��
�LY��
A/J��P���?I��?ac�����OR�S�3� i��$�2Dd���
��!kLA�g�>�t�4"F!>7��� '�}�l���14$�B�� <7i@Qj�1R��C��	"U��a��O6��D��� �;�	%:�b�r2d�jd!��{Z�y#���_}��  #]'1O`\�>I#�P�֛��'52MU�
�z� 7$[.5|>�C@���'��8Qs�'Zr>��a��'v�'�J�C����>d�r�ؑ�"��Ǔ1'���?�0k��`qČļ����D�|8�, pD�O0�Ode�v�S�Cv x�`m��;�"O�����F=B3���t)�)��$��O$m� ,Z��Q�M0�:�����c�Ph�@��M���?Q*���ñ��OƐ���Z-6ޑ�e!
�'�j`��Ol���-jyF �A�A�5����W>a�����Y��*�V#eo�W��< �(���J?4�L�1�L���ħ ���rt$�)�6y��Ȍю��OXi��'"�-s���*���D��fZ�P)B�9ǩ�I>�v&�d�P�b=O"���O1��d�<��KϚ>`�K���&x�-�@��T��1�O�A'��m��"2���� S�S�%�u���R *۴�?Y��?1&��9�&�����?I��?ͻ!NTj3G�)P�^��bH�K��8��y�E���<�uD^<��R���($��x�McܓW�,��I�mK�BPH�"$A�@��Q6��<� �ş�>�Ov ����!�-��i��Q�'"D���b�К7�!ˏs��R�>?���)§F�������?g�i��ڙeSpT�H�q�~��O6���O�d˺����?��O�^4�E[�Z�L8X#��D�9�����xb�Vr�? P�z�£L�\4p3"G40J��9��ZnZH�聃�(g��hD"$��d,�O4��;���WOH�-5�T*"OZU ��:g��trG)��(������FM؞d�C�R,	���	ܹaMP��':D��! /S�m.~]�O�,b�$���#$D��b�L@6\�`I�i�^�
)�("D����'�3@P�1�U'u��er��?D���p΃r��SA�fK�0` A#D��9G��g5\U�"mp��3C?D�@��Oۄ�(����/hIZ,c �;D��ʒ�����ЉrcހkH`�9��9D� �aKK"�h�`�d��#Z�Hwk<D���q���+[D�p_�$̙P<D�c&� 5>IH��ѯ��!0�,D��a��M� �!���0^��9 �*D�Xr��U�L�����B�s��$D��cbO��x���Iө!긩 Vf%D� R�����C�1d�MaC	"D�4���X�`���t��i[Z��a4D�<����k��IS6�F�����%/D�|���Ut�hT��N��F.t��2D���7��
E�H�#Ĩ�����1D���(@*���0j^/Bn�8R�9D��a&$D�dn�g^Z��	�2�6D��b�+�0�1 rH d�$;�5D����n�>O���pb5r�0�	�C?D�D�	�) ����gMȇC�:lq��>D��ѲGڡKS�A;rg���u�U=D�����&YB��5�"<[��4�<D��3a��w��-���ݑiʪA�=D�t+��F�j��.*dz(�dE^Q�<��
 4��t����-Z��2&LG�<)d"�A�|X1�˱�V� ��<���8_8�U@AK��\w���~�<A��S�f�0���(��c�|�<�#現w
�����3�|�<y@�WG�d|9�F�_:i�!Gu�<)e��$r��ջ�� ~��	CQh�<�.��f����)��@�<��d	f�<ٗh��n� ;S��k�5��jM]�<q�Nٲ���S`K�
���0F�V�<�t"j��)hr�A
p永G��O�<9c��M�H��#�/>u��DVM�<14T*xժ1�'�_a��ZFO�<!�NFO�\|���>�`	PA��o�<��ۓB�R�@/�c�܍˶nD�<�D��I��,A�,��<tcs�}�<9 ��6��H�R����{�<���b��z$�T )�(X����s�<q���"�(\��
�?�t2e�q�<9���v|ڀ��I Tg�͓ҥ�j�<�ҍL>4�4I��Z�	Ճ`C�K�<a�ǜ�uX��(oQ�������H�<ipo�2X�I�&�F�<DK�%�E�<����,���e57٢cg�<Q��hg�����>v�<=���De�<�)��]S�����0�Xa�<	�&R))FH Q�I2p�|��f^�<�g��(���F�T�f��1�H�ڟ �R@�?i�X+�<��5Sa,��D��zVC�t�P�c=�ɠ�g
8��i2+H���bX�Z��E ����yr�P4"��,Z3��&%�yX�HB���'i5�ͣlL�E�4ϟ=Wa� � �W%���" *ƃ�y
� x���N�s<�8�����<��ֽ���xG�C�d2�g?��2z߮�%Ҵf�j1�eo�^���٧H�n�|m��@�%똰���8�\����'d�2�{(8��	7����U���0l�Л&�:Gϸ�=��]kkt�ϓ&�v�	$��1j8��
$��xS���z�E ���� �,�3-E����-b�ʐ34 ߟ[��MI�>����G����ζi��?�.'1�dm�AdK�:���[�K�џ��5�)a���ͫ��ې� ���MF(�
	s,߾~�-��ӻo]d��'��iX���c��a�ꁮW�ո�E�T7D1S�d�<A��Gq@�據K(n�`�
وt�T<�@�̘S��1X%l�?A>����yܓ��=!Ai�b"�PpV�-xD<;�[��/|Ly��;Rf}#"
??9�(�~ҰB;��e�u�C.!���p`La<�0B�=�b����3��h�Q�6d$|���%�=?���2�'�<�f�v�����0i��\
-��I�vN��H!�d#�@e���\�aM��K".�U/�f��^|��6�Y12��z�Ĝ�6Ɍ ���� H� A�CΌ��= h���u��/m�<k�i�Z�$�A�'�=e�l��'�ͣ	��U��*��]h��Iy�s��݄|ߌ�J�����ŧZ9��p����ևZ��i(R�fP0p�f��{�!�dɵ.#����(̛TQ4�!ե�"g�]�6J�½KM�<�z�)��b��#}�Ji�pc̎BT��)��ÈG�!�Ǔ�܈���[>g��
��ĈtLz�\��;wF $�F�a��Y";��LGyB@�X">�����X|�Xqf�0�p=�a,%�V��2�!9�`��G:0U	����O��q5�_�:�`0r�C�0���D^�`ċ��_6"4���K)�1O$!�E�Z)m���V�X�da%J0Y<���60���O��3+^4�Q��l�.��"O4����=e���i���4t`q�sO.���2D^�&[�M1E�>�4���	:�	�~󎔄&=��K��� |�l��FI�Bn!��4l-�r�⃤#�����Y/x� h�V"^"".hx� 
,a����6(��$0%�2�	����a�(����]/\������-J�٬S&��R�G�h�Ґ8�j�\ ���J�1��=�"�#,�}���b؞�"�".�@`�GΚq��{��3�ɘu��; ��*6�2ᐕ61��� �G8<� _w% �K�?*E>9����4o��p��'͸���ֽ��!�Bτ2�^1�T��<M�~���FO��M*��M����&�	�)b��N�9(u���T8:T;��Z8Q�!�d
�%b���c���ޘw-�$����*G8l��9$���1W���Cj�{-r��bc�S�l.<Rf���:.Ψ{'T*�b���Ioĝ˓*�D9V�bw�A�L-�3Ƈ�2���`���y�f�*���x�|�)�![/�=�7ǪH�nH�� ���bc�J̓w�4��cЈk`����4
�
A��^�h���3���i�a*
�Ik�9J��aJFV{�<�EO1X���H�1TVbTR��S�eT�4��P�O4Aa-V16.��M_��'q�.�ϻ2�0��4� R`V��Eݡ=�r���4
4k�,X+���HAeE?~�īQ�bÒ��#��T�V��sH@1<)2$I*��'�\Qa$
�9bC<0�d��ʽB5)�O��S�*vl���e�L��A*�-�/�`b���);�&8�`D��۳�O��;� �2wO� I��<��3f��m+�f�6H>��G�#@K���|���]�ZЈ|�������6.�ryr�J�G�a|ϊ�3@@���f&����mͶKq��K4�$T�bb�Z:^������1S>��.�r�!��#VCP��eψ�z
�B�I6i�
�p�������!�9ve��GA؍��_��0j�kF4m?��>�Yc7
b`uȮU��/I8t�p':lO0��!�.9��E)�*�>>pX��~{NP���:2��r����l��}b�0���Ӱ��3_�����/Ѭ`���@!��5\)
�i'>���O�A(�T?��+Ĺ{T�!�I�/3k\�Dk�<E��%�0>�g*�n~� ����"&ꔵ�p�ٰ?&b���O�{Zn,`�FI�O���)§�y�
ˣ�z�����1*�H�h�Ɗ��yª����㗥�f��`��	2b,ڹ��>��0k2i^-Y�!!�O���EyrE��o8��k�P$�V�� � 5�hO@"<A�
�k��}�&-ĀI��K�#�8�4����L$)RB�����D�2��$	N�����Q�	CWe^�,w2�Ⱔ�O��PE �<ɜ'54 CK#,B�T��(�ݼ�$��
�fi��?HETx�r!KX�<Qpc�@� ��`=1�,-ܮ,͓�~������um��[��� xם�E�O��������y�kլ8h
�+f�C��0C�~Y����t��!��\�0;�21N�0��ɨg���u���1ڄ��sDTQ�� d��bl�8U�>x�G"N�E� աg�	�ztLɪ���b�\�R�\�r��';�I��	�5t�����2#xl�9��4
 �SG�m�s�W���O������h��C� E�)�AP�-˝�0��l� ��5�D&4��$
�ez�4J�h� �Th��w�����b�<���(-0��9_�������$�>;�M�;'i�	�#�I�nLI��k��r�� ���Ō�d<>9�E�	C� (�%�Q������%�:�@f�E�=v��"U,ϐ[9���$Nr����!E��j��@w��f����AV�F�f�jQ	v�S>+�����F%%n�i���~Bd��2j��'�~�r�0�T�#�NM�A�D�2��B\4����V�:�A����?!�A˯N`�%ˋ�����U"[�.D<��������>a��y0"?T� i�����	4>����X��	�0�Oo�C���;�� )�����	0.��F�X��)��닎lX��w�;s@�;`l+_��Ȉ�'�M�D씪$�*���	 ��lj1M̤�yB&P�B�(�AćӔr���*>�KФA� ѡ��}���A��4�hVB@*F��`���.�OR0xA˗>����,YV�nȈOR�.x���w.X	Pz�"c埮q$��/I>o��!'A,6^���|A��9��>1Gk����!3r*�:�X�14S@�'�02Cc��xP 0t&�>z;X�3�'�\�w��%t���s֪� X$蓬^�=Ǫ}���>��$@�`��E~���o~0�Z����Z����z{������5/J��c��> �8��_��)���;+�,1s��$2B��r�,�3C�����*�3��A��a�Pc��5�T��c�J���N��ӧ��0q���'C���w'�i��(�`"O�H���!|3g�� 6�lM@Ĕ�(�bƊ�A�ؘ��'�P�%��zd��br��>����	����R�*��@��UJ�;Q���b�F	(v��#	$���R�ԃ ��\r4�F
a�a��I7�m�J<
f���O��}��j1��� ϫX���2�'��8�%o�{�(��Q�HbXt�'�*��%B��H���+��Bv���'��\��K!Q��uA3�S�1�'����招�78vЩ�.�<�@Y�'���"��1)�`HO�spR<�'�` ��@ȭ,�:��v�������'a��˴�1#�x`�H�4.���'�����k�-r��Ъu�W���$��'�����7��]cԎD �����'k���Q8w���0n��a��\��'�Y��*�	����ǕYɀݠ�'~` �C�A�aB:�SԂWޖ�X�'?D-�h��#��l ��:�H�[�'�b����~�@�z+ӟA���)�'�0�I&)7x���kT�cd�l9�' �I��f��%B��Ja#ɐ1�5�
�'�,�1EBO>>Qq��((q*t�
�'��%A`�J�jV��w��N:D�	�'l�13agX�A�li*��.@��'���)F��o�>�bw��K�Q8�'9��1��P�px�)B6�30W6���'�.���b^�w�<�e��#"�mc�'��\(��v�h{��L���K�'%��k�c:V%�ِt��?����'Mm�π�_�p����A�:4z�'�n�HP �h�T��6l �(�V�
�'��HS�.S�@��񈑩�&�p�'�HpZ��U�7��@�d�]]R|��'�@�xᦅ�B:1)G:V�ܵk�'��%�6��(<)
�J�RT����'��U��F��u�<+�GQ9IH�1��'rVI��$�~�IPT�������'�hrR ��p���HY�(��)
�'�^@�F`�~ufL�Cđ���)	�'1�$�<h����	��Z�'�z�1���C���R`� >D��x���3c!۵@Z!p�j(z0���V(��P��(A��H%#־���s��t����0H`���ͅV���S�? ��oQ�s�pAoA*P�Q"O�q��T�/, �����k���z�"OJl�p�G3l���Ǎߞy�!�0"O��4lO�y�^�ag��+0����"O:IԈԛr���9��@1%d�尢"O�I�A*�X��=sT��Di�$��"O:4��Y�C+6�k$�9Nf-:G"O�ĺ �է3 l�A��#j�M�"O��It��kZ9h��ȁgݼT#�"O�Y0s=4�#'� }��P c"O�
Ѧ�>��|�&��^�.@3 "OF}Y�� I�/��{�$�yBK�2bVhȀ&�$#�A3����y��V
4*N�A�	��2ReB���y�!M6I��}S��X����E��y�#Џ���z"�ۨ|���P̑��y�d�%Lf���#�nNXD��&D�y2��Z"|9�mLaX#Æ��y�bY�dR$�����, �C��yҀ�=@>�m�bA�n^�3�I�!�ybO��mXa��A�,^�քz����yrI�bόd�GOA�R�VU�p�9�yE}��ȳIP�PN	�ԋʷ�y�)P�MՆ�r��)JĶd@w(� �y�[��U	�mD6��c���y���8^��G5A=��م�W�y�9l@$�Iцܱ&�*���	�yª�1n�,� �A,'Z`9�	�y2n�&ƩC,��
�x8�S�S��y�e�&_P�}y%�)����R���y�֧��}*4͞�z�Z���o%�yr�F�<��hvo��[�,�P0���yR�ʾR�;�-'f3�T��EF�y" )����ύJ,Lt#6aИ�y�BOG�(� G�� G��0!s@J��y���<�$ �C �24�Y"�ǒ�y�o�*�� �f��.�B����yȒ�o-Z�ZE*�*-�ڱ�%N���yB`�WlȄҤ�U$/F죤���yB��=Zμ$9�I��.�&�#���y��
�`�9w �1Yp�p��@��yB�J�x���E�>W�= !���y\([��<c�@Č\��H��l΍�ybn��`�\����WSl!)U��yj��EDb���Id�Ii�/���xRK�vb��=N-�׋Y�A!��4W���p ߲v����N !�$Nfܰ]J`��2�T�!��Иo�nX�Ŀq'~`��G�O�!�d�./�,@�4����r�p�$�!���#\�ݸ�e��f�8���0�!�$�14Vt��Fk��PA��N-(�!�U)u�lТ.ԇt�"�Q`$�k���>��Je�N�9rM�Nur0#c%a�<���ߤ4�]R���k�# �Sx�<��O�?���4��/L�8��R-NK�<�E� Ud�H! �1����F�<4G.)�̡��!nl|`��K�<1F��V
����Rot��㨔I�<�K�c�hQɢ ёI�ƕ�%�G�<��L�\�]Ca�J��Y���Y�<ad�V�YE4�+�J�����4�XV�<Y�'�9n�d���Y# p��@L�O�<�3�#����[�u��t�z���S�?  �"ÊX	�P�a �-(̦�Ӷ"O�1��œ� �� ؗ(A",��DcV"O�mQv��jnQ�4�Y�F�D��"O����ٱW��H�hn� �h�"O��ӕ6���'B$�tc�"O�M3��6@creP2e�~����"O�i��@D,�|��r�p�"O����J�|�e�Sw�� Q�"O��h�� ��̫#'
�����"O�H���P!f����(%┴�d"O�@Id�@7-HljL 2i�zq��'f���t�H��f��C�|�r�9E�,D���	ӈ*Μ![�KW�G�X�dC=D��q�I[�riP��HH�}�F(�P�>D�<h1郮�np�զ�~+:S�<D�x��
B8��|��O9* ��F�.}"�'Ɖ��D�`�p�J(O�0�
�'�(T��� J���IT�>���'�:US��R8�(m��A�X��;�'���*�mZ�m��Iy�"ޛ!�D��'�Y��)`�MJ;$��a΁Z�<�@��#`H�
�'� L�Jԡ�)�T�<��,�0S���Yt�O�$%H�<96JݺY���C��`H\z�<���,�Ba���(��ڀi�w�<�g͕�(�` �%�8jF��ǙO�<������s�Ή$��@�G��b�<Q�C�h߄���	�zeJ�d��yRe�SU��gC�	q�0��\+�y"��_1��r�4��0-�����'kvmq�G<'-3��8*1+�'X���5�A���2�'����'I��q�f��0ɒm	;��ܱ
�'�[ ��C�
 [�䒚6q����'D I�PA���R��1��1����'B6]�BB�]b�I:F� ,� � ��HO���Ӡ��ç*��J�չC"O���'�P!n�8IQ�E� �4ط"O���-ۻg�Be�'IC�L����4"O�<�wk�9�B$;��+ 'ɚ�y��ХE���'12Zb5�ף���y�c�4�B+�-74�)2�)�yR#H�Q髥^���DS���=�yb�O�Kn�]��=u�i��$� �yb��l�*��B9�^�ȓ��?�y2�Z���˃ʏ"&���`৑.�y��380	jW�/"Ͷ�����y�F�g_$PAM1X>�
t`��x�uӘT٤��I \�bK�q"O4���j�8��uQw��q݆9�C�'6��$�	J; 4`���Mܸ�� �Vt�C�	-��8��b
��Q�م7&�b�D{����$gN����W=�DAB���yr���,�d߂U�t�`��O����A%/X��펝���c�b]i�!�P6�M�T0Z�`�gЌAV!�d
�P�jU�R��C.���W&X�O6!�$�� J(���+�c�䃻Z$!��*�\��"Ę?�������3j!�$��P^n=�[�=����#);u!�d� I���c"��TȤ̂w���u!���E��lF��J��	
:�!�$��9gB᪤�L#�z�RI6j�!�Dī���c���ā�)ĚM�!�� Ќrm�#5Gv�hv�%}�P��"O��P�m�Ľ��� I`��"Op\"� /��Yp �DFT��&"O�ab
Ù���Z�
!>���"O���`Z(4��m��-@3M:�"O@I�Ь��혽зL�c�C6"O���i��mQd�H�����"O:�ZK�%<���/����"O�=kF��,SK*�Y���c�Х��"O6���%�}lk�fA�y
�����'t�'䔄�p晽E%q�� ��y� �'ݨ��7.��"���P"�s�R��
�'�\�T�a�ظ���j� ��	�'�H��ĝcĉ��e�j`�,Q
�'`�q�*'y��9ģ\a��A�
�'Fx�iѭ_�z�d�x�Dj���	�'p��R�D_�H�1F!il^dC�'�F��yL�M�&䏰� �
�'���I@"̧NX4E��#(U��ix�'��%�M�G��yr�"��N E�
�'��ٳ����jo��a�E!,��	�'���9���>$z���eǁ:O�(y�'8�I�"kC3S:ܬp���0,�j�'�n�����#�vT���W+)�����'kέA��O���](%ڎ�b	�'k�(��S�_�rjt ��P�v�	�'2<���䝣;c�\��΀L���a�'5Z�3�O�%G 85��
-�U�'�L��b����v5xa�Ɍ"�X�
�'������ѼX(�+�Ζy� 0
�'9J�ʒOWt���i�+�:qq�'�И���Ћ&.	5�^!�@L�5�y�	����g���,-2���'�y�A�(B�qm������c���y�����|��-�x_�ͫ�����yB�O&5E
)PB��!3���E��yr�
kKbE� �4l���X�ybc\dI�Cm֬)���B[��y¡I�cŢ�[���JnL D.�y��{0�˒�L�VX`k�;�y�
*<ε��1 �dL�r�� �y�Y�n 0�F�${�JPx�e	*�yb�N!pbl8C$�!���6!ə�yюU(����-,�����ͥ�y��370Xd���O�H�
Z��y�h�C5p0�f�<s8�,`�/��y��/P�ԙ�C� kI�hR�� �y��A���Fl<~|�#v�+�y�kQ�w8�h	3�#�v�
F؅�y��G=3���$�A��E��yb��*v\�Ӑc�'
rx%�V��y��êU�샂��!y(�y$O��y���'tv�8�nX9��Sd�̄�y@�./��Xq�d��=��f���y���Nx�JVY�����G:�yR���Cv��@Y	��BPh�*�y��A��аFa-e��#0�
��y�ݶ&�^岁��%(�p4H���y��8/ĥ1)��~��E���y�gMv�6�#V��SZ��S� �y�g�5S����gnT5@L�b����y샇gҺ���͚2��\в�\-�y�
�]MLec�C�$*�(����yrM�;:��� џ'��L�����y
� �9�+�N�t[CB@����"O��{ִ[T,���˚o�rd�7"O�����ݦm��E�7��(�1"O�����+#�@�0$	�5t�E
V"O���#��?#sP,�D$	?|xV"O���7��\O��H�BL 1�a�"O؀�CkA�[��!�(@��i�c"O�YH�%Rv�r�0aօe���"O�1�Q�
�2���	q��ZB"OZ}��6X<b�mr�^1R�"O&IRa��#y��Y`�ȣ)��A�5"O�Y0&�W " ��(� ��9ä�["O\`{s�S�:��m��9���Y�"O��Zt���0O��3��
�Hz�!�"Of�۳�Ǌ�Lx ��t��"OP1Z�h0qP�z���>%�	Z"Of�{���8�^��-�*m��<�`"O�p��W?�툆��|�	I"O6�Ț,k����μ\��ٺ�"O��,Q�M.'�9*��a��"O��SH�)e4 �©��a�bZ�"Op���Z�s\��uh���m�6"O��k�6zC�q�#�\�6e܃�"Ol���E �O����7�5`�\��"Oα�m��_)А1G���.kd��"O����@&rP��g	�}q""OnT�'�Ѹ1�A�m���0!��"O�8� '��<��G5DD�z�"O���6���$-�FN�6�$��"O����ȗ�Ǫ�ф�0~y@C"O:Q�'[6@�s��ǟg�@Q�"OTAG� hIR)!Td�Z\��"O�p�u@��f|�F���P�t0�"O�DC�nˊ�#a�Q9�ĉ�2"O�,8UO҆,�Xh�&��(�2�ۃ"O��B��G!@Ld���D�;��A"O.�@��� Wt�1���%�$��"O@Y�`�B�r��2wBR�Cr��"O�e�Í�l�rD����w���"O�1i�lR�[�ؠP�T%�Z�r"OM�TȔ��Z��TDQT�4|��"O��U�ٯ|��I������:"O��r'fԎV!�����5�,݈�"O���F�8TSxU	�a�*N1�19�"O�� *C�t���b��4���"Ol��E�֧-aӂ@s4}��"O�|�p�]
�� �OM:��"O����2*.1� ޼;�h$� "O��3��.T�p�RȺf�\��"O }š��9.���1(���("O��b�J.GaM�߳<Z�S"O����j�$7��lA��?|&8=0�"O`���Ğ4v���C�Ʌz���"OV�@��S��U�����b���"O�H�be$g�j��nZ�S#0a��"O贙�읚t�Z�㤍˒��RP"O,���KϳI@>���˖�,�H�Ҷ"O ��(� c���
��
�C�vt"O�%�C΍T�|�dGa�E0"OT`3�ɾX�F�s�E�-����""O��0��B�,왳��%}����"O� !ׂ[�p7=r�  �`~~${�"OL�ve��AK� ��O��(o�H1"O����"&���w��lD8H��"O� �T�2�;3?�����2<z��b"O���DH,(*��բ�4]=����"O4�;�'��y��ًP�O4V9~�[g"O(��@"C=�� pg�gH�ݢ�"On��'�U�O*hhq�I<f<�Q� "ODi�u��0Nъ�n��X9�4Z!"Op9���+x��p#$�`(��"O�+tD�p� ��B�p	�	B�"O*�f�!s�*v�U�X����"O>�#���,Pt8��&��4�T;D"O\��FF(O<� PhS5S�F-�6"O���AL�N��q����	��a "Ox�wa�!-zb��倃���0"Oj%� ��ۚ82�˟B8C�"O�(��ǉN��i�S3�>ux�"O�E;�蒓zz�R�B��+��UU"O��zT�^?]��8�g��N͊��"O]�wi�U���QE�R� ����"Op  ���^���yc��#I��)�"Ov��$�6ըD�/Z�
0��"OtH���N3��[��}y�"Ona���ԉ(X���� �r�a�$"O�D�`�G,�� {!�ѝ?��l��"O�pH�fK{�P@���y�b9`"OR�렂ѭ+�ĥdAN2Ps���"O��dmQ����S�!���$"O2|�r�z�����F�(/w�q2"O�i3���]2�`��
�3M����"O��RA�82[�e�"�QyI��Z&"O2��שиr����Gm3<`�"O�Y8B�۔H�h9#�ϾN*X,+�"O�x;w�&�A� !�)�V"O( 0Dƛ�B1���D=)�R&"Op9z��צ���T������"O�%��d�1'��2	%�O�<1O��f�V ���$���8W�Q@�<Q�D�H��賧@�yD�+���S�<�A!�39�n����-��am�O�<y�΅/�@��a��F�8��P�<�k�+�ejӦ �}]�X8u��f�<�T�$?��Z�fT�?.5��K�g�<��΅-μ"��.��p��C�_�<����b���(юܘ]��=F�[�<j��~g֤+�(�f���ǰxC�I/S�L$x ���o>ɘʜ:%�B��:`r�Y��!d{���Z8.�pB�	#m"�9�揁1w�D�%G�quXB�_�.���A�;	�l�j#��}2nB���^T12�L�g|��h�F]�-�NB�-�Б1�#3GlV�V|$��'��U�&!�.U`!A�G�K� T��'�q�dːZ������L�I=�u9�'���Ê�G+��5%S0F�L��'��Ѐ5��V%����Q�f*�q�'��-�iD�# `�ڡn$OLp��'̴�:e��=R�j!v�ůB�$K�'U�)�ٕ��x0C:=���X�'��]����-��T�שԤ))�Ń�'���y C�E���AS���S�'�.س�J]�r��Q��b1��'8V�Kb�@[8L�n�$Q��X�'�R�R��=`O��3��ΗK�@��'z�A�$A�cnZtH�CP�J�0j�'�8�#���V�z���B�:d`	��� \yHaHG<H됭#��ݎ.i6q�q"OИZ#��"1����Co�_�J��"O~���8<��e�R�-1�g"O� �Pe�.W�,t�-ɘ4�r���"O��8 *�-\�r=��k�z�:E �"OЅ�3C�8
:tT@ ��)|g�`�"O�� ���j܈�L�]`XXF"O� "�nf�p��WI޻0�P�0"Opiq��Y <1J!`
T(�p�"O���'$ěA�l�u��6u�-��"O�Lc�/_�L��4��臻���S"O��c��~w�Y!Ѩ�.���e"O� ���{#�bc��!f�⬐�"O�M¶%�/dZ
q@Ca��w�����"O�|��L2u�����'n�\8K&"O������o�Z����Y'#���*�"O�l�E�BU�+�Q?�XE��"O�m���P�q@�*T'}3F���"O.��f��2_Ƥ��F;t�*��5"O�=8��ҳ$�Ɂ�&%!�:�!"O�	5���e�))P��z�VmAd"O��b���N�]�ׁ�J}a���N�ذ�(�U$6�+ΐz꺡��&D�\�'kX&[�����F���Q5J%D�H�X] �ɗ�P�N�:m`m#D��0)-����e���,I�FM&D��1e��P6 Mq5iD59�� �pi'D��[�k��Y�x��#%�3T�b«&D��aפ��R=��T.��X<�@�k%D���p��.Z��h�(n��&��<����Ӑ;�~�rp��J&h��CÇ.B�I,��@��G�U�@�:�\2�C�ɯ�V��
�#�`H��?���$ �S�O+ʌ�⩄�X~���럎g�@��"Oh%���&m�ikg%ٙ��P�"OfLXG*��\W`q���[���i��|"�'������OT�u{���H{v���O�⟢|��!�gy��H2A��Rg�B��Wo�<��@�L/b	jf�X.v��A(&�p�<�w���L�0���d��t٠���l�<�^�1ق$XpO��(��5Aj�<Q�X�\rh�j��;�8Y��.Xb�<1��sO���"�I Z)PQ�@^�<!e�0���"e2hC:,1c��]�<q�ړ/���J�Xc����M[�<1s��+����� �la�0��CA�<�fM���� �4=�)��Dz�<�E��>�}Àʓ�;��UB�O��M���O��M��"�/cly�A�)(�p���'_\IPB�z|�2�W>\$���'����L;f��iaG��OĴ���'�؈�Pɓ�RN�}�u��'A���	�'���ra�����T����y	�'�l�c�	ɧz}l��ģP�{Z¡�	�'��!3��T%1��0���#(�<�P)OܒO�����}�]�Kr��83�S�Q=d�9��'	�O<�}��@J���p�Q��}9��S���C����Ŏ̞<^(Q�kQ�.��p�ȓ���)W��
��X�NG�u�܅�:zHyc��9a�YF��2�l}��Q���p1AĢM���(m̙D{2�'������W�y�T��O'A��J
�'��	��R%l'0�sFN} ���
�'Sp`i���0V6m�âV�s��	���4O� �IgbHS���C���T�l�@"O�0���O]�	p���D�!"O�t���W�2>xp�"$C/b��1�u"O��5��t�@]��&<�*X�""Op���e�s�=�0V���0@7"O�D��N�����^>=�Pd"O4���l�|"� ��I��y�`�D9LO@�0!�٣*�.�j���x�t�+�"O�Y(��J� �T(�A��l�!"O�]����*3l�QƑ;B�c"O|`�g I(n2���ě\�������Od�4�O��y���^�b�h&�n��+O(�=E����p��)�
*`rL�EH���>a�O��3�T�\��A���RG:aZ��� �S���<�h�2�M�+�Lk�bE�y2!�����BJ��j��(zv!�Dˮ���'B�q}����:7u!�$ý}���ă�*`Թ���-^ў<���U�`r'%�1���ó:��B䉹A����S�(���$*�/��⟼�IU�}y�OP�R�� � o������jRu����:�$@R���"\i��!'����"OL��rL� R0�T�J=-Bذ�"O��H!�N8@2����eRPT"O0��	�#\�~�BMq)��LƼ��?q�^6�hSd�ͺ#g�C��}]F�8��x���7P �"`ң�E���T�hOD����!GL�Xu�`�� �����"OD ��P�=������'��=�$"OhU��B
�`�u8���K,�k�"O���V�,\�����qz��"O�t Eܭu�6�	w-���^	{a�'��'!bgP:}^�rF�gf�X��ܱ,!�D��?h��0ug	?^zn�#��V�0�}R��H U�aNh�kؤI�\�E�>D��S#U�I'D�(��	/ꄝ��?D�`2�kŔJӀQ�P�AI�(D���v���`�j �	�\����1D����:څ1g�X����0D��z���%* �t�1Qhv�"m�O�C��4o�9`�FE�EB�,i���, �lC�(0��`�D��h�R�h�O����Z/8�,�����!��A�P���J�!���(���01��M��𲂏��9�!�{�R!�Qh^:n�8h�����4�!���'Ef���.ܡ1R�p%�T�џ�D��ᚈ~=+����g9���+\��y��H�*K"UBQhܰI@�A �.�yBJʅ`���$�A�?L�
�-N3�y򆇣F�d�94#�rp�:W���y"�00*��棈�y.r9W�+�y�V���K��ޅ#�=�Ǟ��y"oQ�(���I��n��%]��y�%�KqT\��>�Ց� ��OR#~҇��9(8���cV�m�b9�&��Xh<ARNOlT�Y�OXPMʠ�A���0>Yv`E�8�NE����>����'��U�<yp��6ReDSsa�1|O&`���Ml�<E���n9X��%+�F\"�H�S�<��G��]���6�C�r4M1�"O���4(��R�Ԃp��FY�����+�$E�G�!fv��f'O�+P�ೠO�]C6�F�A.<�3w��N�n@���<D�����"㾸y1k[Dt@ч�O��=E�D� (蒈د�0]s^�2�� ��"O(-I�E�3�؈��I$>�*@�q"Ov}�q�ʪ]��agG)-d�"Oܴ�Gl�scl���Ԝ,���hy��'NJ�A�>!J��gF"-�PU�-O���dN��h��f\'Gߤ!�$K���{��(�X {����(��U-D�_Ƣl8$"O�9��| �=T��&Æa�<�TmES�`����X���Z�m�S�<9t�޿U`JiiVAS'�viZ��Q�<��IUL�H���%�X�|��0�O�<�2�d�I�ѦкX�F�a��E�Ih��`k!��^���Y�U;"綕�D�_���'�������x����'B�V^p�1���>&�C�	6B�QʂN�L�>��"��$*�C�I�T4L�	�g�53�����X�q��C�	�yP�8�E�M�X���V|C䉼��T[6��.8\����s�C��72~�SJ� "|�@���-E�TC��0�X�2��k��0"M9U2C�	�O�ά��B����#��(�B��)u
��[0-�~�%h���Ph�B��3p'���� Ń)����i�s��B�7]w��K2*N�P�h���K94���=����������b�a�'A�^�ыc"O��{@�Q${�(i8�F���T��"O�ȗ��z��0���C f� Љ�"O����DПt0Z���d�{r�pW"O@	�!	 :M
��QmT4{�*5"OB�ؔ���r����f��G@-��"Ov-(��v<^0Q�ľ(��Ʌ�|2�)�S�7)��"�͐w�x��ת�6p�>C䉫�"��F#�2H#bТ���_C�ɱ=s�@0¤X+=-0|b&KH���B䉅`
"�ҵ�	6Zy|�4%�
�B��=l3-�Q��(0>A�ScO�p�C��5Q��R4�M%A7��y�FڔC�2r�<��(�4R�|{E$K�TT�C�=��$����.%Xƴ��� -قC��4YO���EjI:��Jg ֚�zC�I2Y�)�gI؊2���P�S�M�hC�	/om��휘o���ː�3�C�4C��x���B�{C&��c+�G��B�a�z��3����훧��b!C䉠+l��@�l�bb��fD@ Z�B�	EJк��܆cj8u��+�D5���0?)�J[�_dQ����_٠a�EeK�<����"l��3�i�7��m�	7D��r�)�)U�J �4�ƫnC��C�5�$�OQi�Nd�Z��;���C�"O)�r�& >��BC��P��"O ](��G"hٖ��g�J�UX6qsT"O.��u�8:�|���/R9I���"OB9����9Ie�c���A��Xa&"O��g+
NH�h��/˄m{��*��',�LH5*��g� �.�J.����%D�P1�L�pC�ҁ�0cc>���9D���%k� ����{BV���K8D�А���젫�`W��&��"D����O���!*�a��l�@!�U@5D��Nϛ}[<��b@ޙf�n����2D��@��K�H�Zh�P��?<6���0��������� .�:�0`h��C�p��C"OX�:��ˁ;��Y�RJ�!e��"O� jŢ���*�� i	:\�u��"O���Ǆ�e�HLj H�6����"O��7��� �#��<)R�-�"Olp�W�4:���h�( "Oέ�S�־C����@�ҝCS��q�OJ����M]� �޾}�d!��'�ў"~Ҥ�ψ�ˆ'Β͠��c�)�y��D�h
�*T�U����H9�yB�U��A�4LQ�	J�
��y�N]�H��A���̼sg��CAb߹�y�%S�=y�Xaa���g�E�  ����<A��dR~�xB$((�\8b�����	S����<=p��I�DeDܩB	,A�0�B"O��%J�]^�9![&2���"O��m�*2�H<q�-N�=��M�"O���Ǝ�SƜ1�s�ڥv�^�H0"O���*��tJ�:�,]�e��D�P"Ob�"`O	)6����0hvpM��"O�Y��WA)�0��R>f_.�t��G����6���n�0t��h����+�y2�O�v�*�L�. Ґ@ٱ�ƙ�y�N��BH��0�x)2����y�&�%1v��ŉ�ƔI	���yR���4�2Us`�V�h��K°�y���&!X�����Ą�� �GX��y����]�vhpe�*d I���y��W�@50�rV# )��Sgk���y����}�:���HU"q�8��&O�'�yBB��`��I�oG��v.�%�y��:�h���ET��I9�iR��y���9�d�AN�M�&`@�'�>�y��?Xd�j�O S�p�ri���y2@-n�x<�q�ЯI�F-҈K��hO<��)R:��P�MR�Eu�mk�"����'zH��gCXgJ�l0��Ξ�H$��'�D\J��ϐvR�2�`æ~����'�,�0u��]ᆦO�{�N���'Z�@��L�qʨH�,R�?#���'�EI.�	���SV�j��`�<�a�>e��
G�F-m�4)��BM@�'tB�ӛt� Pۑa��Gn\���˗6
8C�ɚ��m:�@f�Z1�T�׌:C�	�o0�M�q쓝0���!��8*R�B�	�=X� V拥M�]����i��B䉽>���3��Ǯ��8K�c�;r�^C�IN�d�AF[(���TF]�#�LC�$`�LZ�j�9���Q��tQ*C�	0r��] �$�!baR��G/���C�ɺB�tݩ�0n�(#�T�C䉹V��!S��%�����H��=�|C�ɘ;1�s��<@�xQUdǃ�tC�I�w���ЮL�A:h(z'�J]�B�IO0h�y�cœRP2�)��$V�B䉎@�D���օ;Ub\pň)��B�I�-����3R�6D!FkG�I�C�	�k����c[`��J�Ţ t�C�I�4�a$	�)�F���� 0nC�I�B0�%rrc�+�X�b"J�0��B�	,#!����\"[B(`Fȕ/p�
B�	>e��h��m�!C2аԅ�$-�J�$.��V�1����W$Ay�N��S�2D���G�B�|�t�@�
'H�s�6D�$Ó�G���eG*��xEL0D�PڔfP||�I���s��p�/D�� L���O�W�޸x��[�M��;�"O����oZ*V�*����J�~�v��"O�j�kA9x���욂[Q�J�"ON�Q���Y�(�h_)9�h��"O���wo�B3(e3�*�t��M�d�N�؂dB�"392� �gF�U���-;D�`[WcN��x����vӎ�j!g:D��`�N��
a<�kn#
VY��7�O8�ɔd"J�R�]�f�Q �Q�6�C�I9f��x��ɀS���@�91���$��Jq�'w�8�HP��<%`�ȓl�>՛+O%y�������q�<�?��$�t��k��i�B1��KUel�ȓDe�MO Ӹu�e�5kF@��ȓ^�Y�B�≢g�Y�v��U����<I���b�!�G�S%vj�����P�<ц��Pk�H%�N�S�����MK�<)�'��z1�3K	Gd��tF�<�#��ncJ �`C�
�d��KE|��m�|�R�P�Tdaa��6�qY0�?D� �H��H���#��Y7����	<D�ԙ 5��`�P�ې,�6d���<D�$��ѶD(A%8��:�#-D����H?}�u�"B�Lqj4��F>D�X���X���P9�����<D�pI�D��
�T�q�"�E�)�$�;D�`5*�)A�Ty���X�2"�-X"�9D�	��
g����� 1���Ŧ-D������"�r�Fԑ�n�xD�-D���1L��{��q���ҷBȄ�� D�<27Ƽ��Q�%oܘ�N��V�,D�H�ԍ�X�ZM�ǕfC`-))D��c��
4�H��	��*!�Qd<D��A��V�@�R5���ȻT�!�d�-D��sr�&K�Z=��F;\�(9Ȣ�*D���3�a�}Z͂	mF����)D�tjrMO0Dr<�ӠcB28Ԉ�#fn)D���OJ�NmЁ��"A�(C�p8э#D��c�m �� ��@<����&�O����*Tؔ�<k�J����B�3?V��B�W�x�rf��'e�B�	��
�˥��q����UCs�B䉝e����3�7S��Yt��,m~B�Iu��t��'ڂH�i�kx�B�I�^D0aA>��Pe���e�~B�1}u2�m�x2��`%�L!8RB�	'33�(�5�رt効x��]�'��B�I5}x�6L;^�"ʚ�MݠB�	�>^���n�"~���%^#%T�B�I�c�LAi+4�vx�3��G�fB�	�zyb�`P%�s.^��0c� BdB�I&EF����4i~T�1�%�)��C䉉'�t�R�?/:�bq(љ{-
B�ɵ��0(Rh�"B$K�?	��B�8�1Z��A6M���
�4��B�-'���q$j8�Y��k�98zB��;l�ȰSUꂄL�)!�X��VB�	<a�u*�-�-X����b{��"O�H#,��x:�VF�1(�h�a"Oy�!��~�<� ���v�s�"O���ԓ?��e�4�'*�qC4"O҄�LS�ѓ�L 5Az���"O�0Z��+}l�)�ǈ���L��"O�8��A���09��esB��"O� �1�EDZyL<St�I s���"O�iIS�D!:�h���U	~�e0�'��ɒ^�M��I�r����噞'ʐC�9'~�AǢ˫b���P�j��6�JC�ɈK�조�a�&_:���e�Du��C�	�m;x$زfű�% 7$�DB�"O�iC�m�:�,�	0Oup��u"O�`�4�N�����gM:Kz�{�"O(9�e�4:�d�WG �uA�Hr"O�]`��J7/^tꔫO"��4�*O�����Gl�P�A��C�P%��'�f�z� B�<�nQ����#4XX�	�'f u���	a|�t�#GG-Q���z
�'��!�ui��lH�����)Q�D�`�'a�!�P�e?�q��'���=�
�'p~cE�ǆjb�B҂��EіY�
�'l�m������<�k��=�&Ū
�'�T�
@�'%�����	�*�X
�'PNe !/X?`���ѣ������'L(��$ʹK<i�'�ϳ�pё�'|T���>� ��b#T��c�'���q��A�A��YPb�c�����y2�	r1�$ #��iQ��ѕ;�b=Z��D�������$!�J	�x��\-6T��rAJ�G�Z��ȓ�DU��ł:h�2e��de�ȓeepU[R��i$�����N']%е��g]:]"7W)Z���Q����{���ȓ� �	��<w�B��sh�,���G{��O���$��7��qyeB�9�bQ)�'���3��L��@� �&5���'�HT��G�Qh<���(��z�'�ܭ�B���	s
.(��}J�'��l�#/��iP8H ���~a��'�h��� � AN� �R�_=����
�'�d���>Q�����2���i
�'��Q����Q?x���Ƕy�ԈJ
�'|<�A�T�_b*�"�h9�p0)
�'c<�K&�İ/�eI�E�.�H�
�'|V �!"�]�8��"R 
M���	�'/T��wJ MW��UT+*e��'�$<���m3�����6L_�M�'�(��6@S�H;�I@b��<T=�,O"�=E�T�KH��p��-���zpϓ��yJ���*`I�,'�A%���y��E���q�Q�R25B'�\��y��U���Y6]đ���̨�y"E��b�Pa��E:5�8 �B��y2	��`�T��d�	� F��v�N-�y"���U��!�d@�p���!AC� ���hOq��Đ�N�Ct=X ��k��$��"O��!���&/jeBg��M�D���"OZx;V�<1�I�'��6�-��"Oԅ;��~����'�#��M��"O�<�qE��,cyKt��d�޽�"O6��7�I3)U��ă>:R@@�"O��s"�z$��Pf#��N���bR�|��B�S�O5$�H�_��Abj��g�]	�'�4�2#�;��XѠ\�Z��d��'���#���,l`��EA�L��	�'�j���ܵ5*�wKL
F�f�h�'T���+��R	{g�*bVԊ
�'A��0�Ex#������H\x�'ў��O�$���z�$		n����'��c.��N�k�8>�,�p�"O� �Y7�~����&�!/wj�S5"Ozead�Jh9:�Ϛ�K���"O���A�E�	� x��A 6�T�v"O>0!e)M<����u/æF���!"O�m�W�Z�h]l�)0E�UJ�"Ov�Z7,	�twl���C�U�����"O+R�F�l�p�u�W�`�j�@�"O2�B@��c� �`a��>�:� �"Oh6,��	fL����ߍa�d���'��\�H�8����'3��xHr@G�!�DO�"=�١�c�it���Q��+���7?G�9��bۈ���;�y�*��5Ѧ���nFf���)���d5�S�O-T@b�XD�BM��h��o�AH�'@�ـf�ҥj�zeʤ`ٱz#���
�'3�����*�\Acםy�l�
�'62�c�Ǚ��=�eÌ�@�:e	�'����B�(A $	�[�e��e�	�'Z���wn�99��-0DQ$T=&���'V(���C�clZ��Rf�cu�I�K>���)T�C��e����$C����h��Co!�Đ�T�b�aaԕ~�h��Hfe!��"1!���ek&j�>�Rvh�"g��$�k$t��V`���T�2�ͪKb�B�I�F�^eӡYd�=s��ʟ:Z�B�IOf(�+�"S�P�"M�	E+.C�I�J<nx��F��:+i��P*��hOQ>�Hĥ
&/L�F�(Qb�rg�#D���$O^�j9�tB�Y�� �Y��"D��8u�F�(�h-�����g*O���a)5��`�,��m"4"O��*`�ѵvOXa��W7V��� "O|e ��
,CFҨ(4$�4m�,M��"O���Wḏ<8 ̹�C:c����3�|"�'��Orb��r�H�l������ �� "0D��*��a�^���B�yCR��׊.D�`���́moP8�)� u�UP��1D�,��AX"OB���Cn�> 
&(�%0D�4����96���T�"'[�@�gh8D�䨡I:thaPh�5G�v0H��5D�� �Β	��m�R�o��c�7��<�t>�+˜/Fx��1ņ�|��D��V1Nع!C��qu�4��bОDݮ��ȓ<X@K��R8k`�Cデ�:�&����,!{>�0����TA�H��L��B�I�]�����d�r*��:c�B�t��B�)'i�)���QB܈�`�+PYvB���j�jp�M�<N����ԯk��Ї�3�F%�O�K����@�9#0BB��?'_Թ���q�0�p!�4x�B�	�.od) F�W���[�jl|�B�I62M� �
�,��ip��
�B�	r�����R?PJ$!ە�Ǻd��B䉇0&�d�ƌ�6Ԩ�&�C!��B�	%r>��@�|I)��E�I��B�I
AX��q ��	�LY
u�^C�	Z�$�	�OA�U4u	�[�}O�C�	�A
���jY�p_ڠ��=C�B��$ow�`�P��0x�|@&�SwnB�	����䏄it8)���*�^B�ɖi���@�n�D���n�B�	k�Ҵ�V�R��څ
�:�VB�I �L��T�xH���,Ѓ9qBB��-x1N�@!)Ʒw�(�+�;%l�B�)� ��An�EB(����R%.��6"Op�D郢T�(|��<H�~�0B"O�]���-����� 4e�\��"O�0��gُl��0�`,�o�ޤQ"O>T�vm[��Y� ��4&,]�O>͚�/Ϊ'�ؔ�T)>�4@��E+D�<�(��z��%S�+N�$Y$��A*D��"-�l�А"� �wi�b�(D��j���N3�dC�M�{����3D�L!e��w7��� ��^�0Yb&�-D�8�S+�f!Z�Y���
M�@ٱ��-D��ÄOZ�Z�b�� -ח�$�A��-�OP��4a�4�t���{j0��T�λ=Q�C�	 	�L��S�V�(5y��@��C䉠^�P��C��b��L#!7�C䉲<	��:��/�� �KFgh�C��&^b��Е�
N�<krjW(<�.B䉒Q%�(A��#}���)�`֘N��B�I�yd�T��%A�}�a`�I�-�����0?q���!B�sNZ�=l��É�C�<�e�U�SR9I0GF�	)���6�B�<a�Y/7�>qcC���0���'�8T������x�ɒ��.IQ�Y�g D���V�L��*��Hĸ2��C��?D�6o�mt|)���;8�i{�@q�<IV�.HF���P u!�˅p���hO�*�h�^O��Z�������[�D�'�ɧ��>��c��r;a�(��8���CFo]h�<�a�#6l�����-z=0��dBM�<�Eh��}&X�;% �(b�JܺBBO�<)��
#m��C�I;��QSp�[I�<ɇ�O=C-Rx1��Ð�j(���G�<�t닔	�n�T�)^ZC���A�'a����B	��V�U�6=3�ٞ�yBnY�^�0-h��H�%�Z��K��y��D�3T�0�	�|ּ#uZ=�yRϨp*f���I>���r�o���y�,c�J��lE5�*m�T��&�yB��	P��a�2"�9�y�A�ڍ�y�(J�cmv�{���`�f��d��yR���7V(ĲR+G\P�2��i9�'#�ڔ���N5�U�E��7b��`(�'>�H��R�")���5HJ7rlQ�'6ȜX��%X�Di(Vd@�@�,�@	�'�hQ��*��R��$8��U
D��P�	�'�T��aȚ=�Bț�F��6��X	�'n��R-M+B��<�F.%Av�hK>����*Q'��8A��+e�l�����Ak!�d.�Sab�4̜��̋*g9!��2#���-�p��u�%F�Ԛ�'�H�D�d��1!�H�wI$�z�'��	3��� ��Q3�D$uo���' ɉS �Pn�D�!�0|x� ��'X^�b5F��.��`�{�Z0�'�҄ǹ�N}� #K�~���'��p��VK\
Q��H�r@�'�� !lײm�T#oR�2�����'��x��hN]o��ip�F� 4�q	�'+�Q4�oO$(U�S.{�4*	�'?�`h��bl[ծM�t����'�p�� N� *�$Kd��5i�\��'��4�p�Z,z��H%�ěW�j���'��]1���0}2��D-A#DPH	"�'�MC�/�39��"d�ĝ5!<k��� X%@��v��Q�"5l�j�"ONX�w�\9'����e?V
�,�"O��Bv�*L�<���S�]�NH@�"OB�k�AC�8툕��;?�d��"O�4P�Жo���q#ܙlϺq��"O�����J�	�Z "�L�)>���"Onq�bH�.?�MY��X�V( �"O<�s#�����b�	U�ţ�"OP�4�B�T�j#R��:����a!��#3�48j��$? �(�INd!�5�%�A+8�]�/E�uJ!�$��&�p��'���������%L!��L�4%���4���2y�f�V� �!�$��]��uӤb�H��Xu���T�!�dW�<�J��֠M'|���nX�!�䄮�d�D��wh�Y��G�1�!�dS�|� ���t���b�l�A~!�\F�J����qz�<�e�J6TL!�D�	���6�O,�� ���#9!�DD�P*D��5������bF�"/�!�DS5E���9p�ϙX�nx���	%~!�دem>��RG��j$�w�S�s{!��"��P��IGM��'�!�d\�4�a��R1X��	d�S?}�!��ѡZJZ�rBG^�:�d�Ȃ^!��߲�X��B~�� (�)��F!��KQ��M{!e'Z�V}��>c!�$S�V�P&Ğ�u���X��'/�!��Q/:�����@0�c�*�!��Q����@�7{iYa�!��$S�Ze�S��e����a|�!�D^�f�4��C��$Is(�X#�1�!���?�Z�(����K�"����ѥ`�!�D |;ƙ���ψb���O��C�!��@;Av0 xBI ;)N�a��=gO!�$J�6��� G�1�v��k�A!�$B�;F�����2�bI�EjR#!򤊖3�.������	�锝!�D@2/�DA�(E=U���:ЈO��!�D2l�F��
�.��q ��ͪ�!�$4(��G[�Vy�YJ�f(�!򤁎/�.4 @P*nr<`h�E��1�!�D��v����O���Hq�/(!�اc4�i�tG޷,]t+pO]!��
�s�T%��d-'&��˅�O�N�!�$QdPA�������盆2�!�dئ!	~�:¤��^�9WG;g�!�$�w�:q�r&J�r�����E8�!�D�1D��A�l�����J��J�!�dYz�(�� �?i�"H�VI�`�!�$�}%(�YU)�Z��_>�)[�'��,`�F/�h��,��6ݜ�9�'A@X���&�6@3���5�j��')"��ro��N�m1�h�3)���`
�'c�B���+aO�I�HL'�����'�T���M�]eK3�Gp�: ��'�=�kі�^�����l����'�	���ē?X�LI�ۘ_3�5�'ɠ= D���]r�"upD��'��Y[�(θW p�ӂI(Ȍ���'�B5c6O�3Y<�u��J˛b"��	�')��2��,]�`��H"�؀	�'U�}h��>{�L"`BN2>�<�[	�'����K�z:���WϘ�N�(	��� �	:�R6�t�p�?��"O杠!h�7��4�.��T�p��6"O�u�3%Q��X�l�R�*\�P"O� ��)O��Ͳe̖B�ʼ�B"Oua�K�dL�� 6P� -�W"O8HR3"�_Mv`�&�	?�m1a"O��HF&�H�B��7F� "O ��3&��+����Gb֏��,�"O⼰7H�����#N��R�BF"O�Y�-Z�07Z(r%�Վu檕�s"O�i�W�8C01K��^Ŭ�S�"O��EC�o`8�u��I�����"O��2�I5Sd�A�SD�)jfA�"O��.Qsh�R����E]�Q�"O�%j�C�7M�H-J0 �/<"x
"O�"2ǆ�r�ӡ��B'�I:"OB%�f��/gKD�6C��=���C�"OZY;�-:'d$�C��	��<�@"O2}*�V=_zh�ڔ��zn��i�"ONU�"R,գ����1�8���Y�<��Q:4c0T�af�&s/�4B�C�R�<��G�����Q��l��ű3g�G�<���Ζd�:|(��#x���y3�DH�<a��԰)��%QrƧg F��pi�G�<���H�s� ���dX�m� ��	^�< MK�l���"�
gG�y�(�X�<1bED'p�@��#8e�]��*O�Yy4G�?A�\�%O�C�z���"O��(�+�X2^��BU X�Ab�"O�Q	vKL�/,�}��&S�,�����"O� Ґ�@}��#q���-�y��.#a��#�_,I���H��yr���<�Ұ+����Nx9��o��y2��+ɬ��.P�Cf��*�J��y�b<�|A���5ݶY��δ�y��p��i��-�5xӅ��y��زQ_h�b��:���'�/�y��^�OWZ��סF'~�����J �y��Z5M��#�9|��IT��yRO�,4�j�i�)V�rN�����D��y2k_�$�1zv.#q��h ��yrM�*q ���$"�>p�L8����y��:�\��F�Pl�*`�c��y⇌�E�x�!2f�!rQ	V�y�
P��MX�dpfQ�k5�y2�T�?�l��g�!F[�F��yr���
�� U"�#:R���)[��yrH�,@��Q�C+G�$8���4&�C�	&7�C����|D81���ÞB�I�,ʈat#�/ے\�c��q*�B䉢$�%��⚞h�\� 0�J�T�C�	�b�N	����gy����=��B�	�
��Mj	lcP,�&���0�ȓxj���!�{���x��ߊ�|��ȓ-�hH�JJ*W4v[G��i^����	��� �f��"��C�� T�ȓX��H�����4�sf�l��ȓv�0���
����Jb�<9��[�f8r�_#�y���HWy��ȓ�6����5�n��lRc}<��m��erG!�~m�X$�U+,�f����l��(˷J�,P8��%2݅ȓ$j ��T�H?L��M��%���W8+�ޕ"�V`(�eȈߨ��S�? ��	Uj��PX��\0�s�"O�!0B2?DЁ���@��9�"OH�s�ZnnIbg�՛bN��a!"O�,��(�6h��� �;dI""Ob]�ʊ2'��(�,X e�:Q��"OB�ܭcV��Y�˥tfh�i�"O�m�t��)dB1``�ەP�Dq�"O�8!� Z�6)�4�B�Y�XJ��`"O�Q��	�a��D�r?��B�"O� ��G�5x�9��X1+<lp*"O� ��W�Z��rs�	�~*y�w"O�����3p2�u�r��kh�"O�,C�'G�WP��[Q�[�M0��"O�Zv��L,|D�5D���Y��"O�\�F�o�F�Kf��
�\�s"O~�µ$���9��ǯ}~�e"O �!�H-
:���A�;�%A4"O$�y!G�ef��g_2$�ȑ�"O>�"��py���4��1�"OlL"6�Ҹ ���*��B*bxQK�"O>EC�OC+p��)Q�Z���"O@�J����d�q.	8^�:�3�"O�P[P�N�)��t;�c�<{���z�"O��rK��8̙�W�
5{�x\0&"OnM�� c�&��$Q2h�(�a�"O6*��Z��²%܃BG�R"O ��Rk�W���EO���Kv"OF��U
W�����IUHɑ�"O�e�`��� �&!�cF&(t���"O�)��ꂰ;�x��[�e��:"O��p5-C�m�Б�@�85�5"OLRC���2<K�-��j����"O��#��W�������Sv"O�MHT"�@Fԭ
e��D�veIu"O��1H]4SO`�Cŏ�ٶ}c"O�P��b��Ч�X����"O6�Y�Ðx�@ØZ�M��"Op���y��)x��@�H�[ "O�i�㘎>tt�0q!���)��"Od�a1O	;
WL����%�m(�"Or�0�� /Zh���� =y�@{�"O����'N�L|4��p��;:����"OFH�v#��(�����إp%�L{R"O\�:��z�FM�3o�?�x�"O�j�AS*���qN^0�Vy�B"O�P�cq��1ƬA���"O~ua�F�!��0b�"TfQ>��"O@+3o��?�(,�'g��tB�0�4"O8xc!ڽ�ZIE+ƉV2 ���"Oz CGH�*��%Z�Ĳ@�XSR"O�9
d/P5� 		�CV&�����"OF��bH)0�pX�̞"�� ۂ"O2q��ڕ��=��.7�*LBf"O*�Ӌ��AY$��G��p/�l��"O@��®��
�@(�aꆿ}����"O`e9`�@>��J��() ���y"jγtb�80���0���@��?���d/ғMT��E���zc�@y�E�$-��ȓp2�}B��0�"V(k#9��g1D�0����#XEQ�τ
}��Kbm<D��Y�소=Z��i%#�1�$P�./?Q	�k����e]'c. !6�\�Ar">Y��!�O���L0Ja�|K�E�J�����
E!�ć<m��t��_,+�B��f��+ў��3� v]*��&s��L1,��%���򖟄����Q)�H�����[�M�3�R$}�� l�����>隧���l�P�°.
Y�ܔ���HPh<���̧`^�Eb�����
�
,�Mkߴ���;��?�O>��aDF/��³˰M�(�
O(7mSn0]�P�+%����	�/q!�DR�e��,B��6�$�"2=W1Oc�dF��6��t�&� �S��$�EA���y��P�ZR��(1�ŋt�N�@2�T�Of��X>'xܼ���6��AgF͎*%!�B�C�\� ��>=XDZg��+!�BO΍�����m!�� =�����'Y1OR�����'gA0�׽H��(2�"O�@�S��!JN� �@��J�B�"O�9Xt��"9t��W�D�"��e�"O~�!@���zת8=P,�
 "O�%1e�ۺ�Jh�D�[ 6��!p"O8!7G�V�T��R0B<��0�'ў"~�c�8{��@�`ƨ%�2\PD����xrν<��A��0 \�� �Oh��B�ɿK��B��Q� F8LqElY�;c&�=Y�O��	ئ��OnZ`	�{Z� ���qs�Uh�'��T��ꜘ9Q,Myu�B�	���4�c�DxÈ�l��\ڲ'
�%��a�N}�R�G� �4L���j�؅ȓL�P�!a˜�k������IV�9�ȓ��Uj5��S򄣱��<'L�'�~҆R�E
�I�K�y�VQYcHK��'az�cJ89�\�'!�%0���W��y"Aՙt �P1ӭF�d�r'�W0�y�Ԅo��LñC���jW��y"�W�	$X#�� h�!&L��yb�Lu.�u��6��݁�`M	�y 4�A�b-�-�R%{�,�1�yR��m��5x�":���jT���yb�-��q��o�+�"(��5�yB
ƹ7��jW �ȠRC��y�k�k�t ��M�w���#�X��yR
��!���iJnlB��
��OH"��F
vT�S ǴH�Y7(Rr�<���]t~��B̕t�R��V}r�)ҧ&-�u8�c�G�4��Y	8;0<��IEy���-�&���*��ꐣ��HO��p>��lT�!8ށY2�� @���D��<0�O���u�dq������4�;��H�)�B䉥i��$3f��[�2$�r���o��6��������|����4j� 	vGϟ'RT e �s�D���h���x�ϑAPHģ�J,���<�E-j�C.74a�6Eޅ%!�h���z�'�`Q"�^:�!�!�.�	�'in�b�K
�r�6���L�, Ҩ�	�'�d�؃��<?ZD
b���i��'J 4H�"��B�����+��ř�'V��ɄH��M�R�I�0�֫�m����d7�d���8����;H	�I!=<h!���T��瓡j( qB��M3SN�OԵٍ�d�L�$��1`�uc2����|��,���ybϝ�NnJ���@.��;VI���M���)��		ꍍRm.4�0�6�x��ǭ D��#��oJ�t(tJ 0��cUC�O�M��	�+�&����҅�1�%*A�
�^��x����!`�{�f�H_�L#��ր-�(��ȓ:��1J�ͥtv�u�S'~��,��ē�?��'����ա�f?��°&̊I��p���O&��� Z���B)T��� �^?ʀ��2����<ٍ��O�,|H����t�н�![�r���'���ecĎf�f< ��`)�F}B�S
�дQ�h�Z�XvoG�C�n��M���Ĉ�:,c� @�ZDB�ɂ���q�U�Z4��H��n�H��t��h��|��׳\v��hW2x����r"OFU�P�Ǔ(���`e�u�g"O>��7�!;�R�Ӡ��<�H8�"O���]��P�C��T%�<��s"Op`I�͒A�z�{ �Y4ڤ���'M�'����i��\��c���l��'0<(k�i�*Xd�(4�����)ۍ}R�'|(��'�B uX,�TEW���9��[�4��	�Z% %A`��.3;��Ì�+7�`��X���N:4�����{J��V+�4��<��8,R!M��)S�|!�H�2+����?���~��,Y�Űs�hZ@�7_S�<a�mJ �nt�⧛�/�J+#/��<y���w����q��a�ԁ�4;0C�?�fy ��=]� ��e	/Nd���>�#�Y�	�p��\b�	1�f�<� 8^�|��F���ED�W�<Q���7]
��.
�Ԁ�kܓ�y���!�Dԣkr�`5	�C�:����wD!���m��@{�I�%� �D,�Q�!��4Ej.�͗����R)ؔg�2�F��������c@mX�P��$�S�!9D���KZ%]�x3���' �2)�G�:}�>A/O$#<1�C�!nƖlqg�ɧs"<̘��|�<RD�>g�l��B�"I�$��Ү�:!���)�矜�A� ;�4�Q�K�5x��$Ej;�c�D�'����&)��P�B��	d
���|�B�=�O�a"�3���B�M���Y4����<�O?�m�l�Iݓ(bl+�ΐ�fISS�!�D�h�P`1W�%z����� !��O��DzJ?K���34�,L�N\$<U
�# `2�O��!U�qk#Nˇ(tLbJ�g3���F����ĥ�~`��E���'b"@�ȓj�~)��O?oG,4{��9U���ȓgx�|��"��2z���D
ѱ}�PM'����_*��9�Ԯ?�ԝ�b��'h�,B�I*i:�Y��Nֹ(��ib�יX�B�ɾn0�	�1M�CA<캡�ʌB��C�>h}�1	�LF��`�@�!6B�	� ��R ��Wc&D��c�J4�B��۶dЎ͇DB��T�	$>&B�I!O.,���]���]��ᔳ'RB�I5I�#��L�`E[RĐ6e��C��=�,a!LA�` �xЇ��C䉍��d��(��҄U�z�C�ɶv$B� ��V�`&<+A�Q&dpNB�I -<�@�	�$�.Y[��Q#�TB��:u����5��t Nh�*B�	*o�(:ի�)c��0���4"~�B��>,b�2�b�6���煞5�"C�I�d�\!�6
���iU�>B�I�K��1��_�R�����O��C��"u���ɦ�݊3%Pb���B�Ɇ|xl�a�+}�ܡ&ީ	��B�I�q��z�.�7��\��
 ��B�	/�J��oS�M�Ż�n�._ƒB�	�~�8���4tzޜ��C�;�B�ɢ�n��A��"U�P(��B>b�B�)� B)�-_�!���o$�z�"OV̫����2ZPĢ���f�T�j�"O�8��K�&t��h!�b��8"O�]+a?}4|*��l�h�"Oj��5,F�Br.�Y���7\�"O*9y"
�"m���f�6��P�A"O�u��M�4v_6�H���+{N��"OP�Y�`��<�-��i��π��y���1��T��D�Y�عc����y�݀i2�r�B�М�C�D��y�QVj�����Ch���� �y��E$#�j�Ғ-�1	W6�a/�,�yRFF�-Oʀj�@�)�؜)��y�ē }r�Ƀ��&8�&�ɪ�y�혍q��H9�KǢ ����B�B'�y�@/O.��+��_%q�>���6�yR�J�P�d�	`!����I�����yr'˪=mv���	X��-2u��$�yrA�_�N(0��ٶ}8T��yr �=f��Д�Ѡ�0������y��A�&�Uk��	^}"Y���ɯ�y ��,B1��bʸ�Za�)�y��C9@Ʊ�4I�*<�p�Ž�y�`A�F�*L�b�N���s��?�y V�P){�c5Ex�IíL��y2 M,b�Lk��MC��2B"K��yR"Z	�mx�I��0�B)�A@��y�/6v�V�A�Y@o��������y�F�%IHL7)3v��� �˽�y�kJ�K��u�ͣ.���'.�yR �*&p(�!ǚ�zy��a�۾�y¡�;&���Ȍx#`���+�0=)���?���`Ԗ	zN�!�T�c���Ra%7530�k�+V�<���FuZ��O73��M+7��Q�<�1�%S�
��F͏�l`���\{�<�c�T��ص�sM]/3���q�J�<�"E�-3v�U��	'C�0yq�E�<ᤢ�v����O�' �Е�5�@�<�3*˻5�bML��v4 ���<� -��`�����"+�Iy���R�<�eÉ8Ebx	�P8��C�G�<�#�I*?n�H�ia�>8S�nX~�<��	ѼWXp�K��_"�,��7E�y�<��Ot���IK�-H2��B�<)@�)\V0����<9ȼu:�.W�<�h(nf^�"�;dtTԑDn^Y�<�ڏX��ȵ
��?`�Q(Z�<��Ή(�@�Q�M�1G/6Աb$TT�<�SS�&�$x��動
bz%�b(�W�<y�B&4/�ÖH�&�� &�2D�XBd"�*;
�QF�R�<S��X2�%D�D�$꒦8�>(�auX��U�=D����$�6*�R� ^��1�S�8D�<rVF�'(�"����+v�mz� D���C�+>��jA"��8���;�H*D�h��l��'�d5�$=��uqW@)D���g@�h�2I�u��}( �2D���b�IN�i�l¡y+�ŉG0D��k�"R:^�䔂gD�%s(2=��1D��a�هf ȭC��H�9�r� D���2�?�T�#!�S�h�A���>D��2��ڬ���1�
ڼI���xCm<D�\�#�,t1̓�lվf~����!D��b׋8���E��w�|1W:D�� X�)��3_ �S󉐟HMh�"O�3���"7�Z	A�ġ@5�""O��� �̇!�j�Qc`F�k�X��W"O̥��Tf�u6V�c�� �p"O�T"�bZ<ĉ���v` 1�F"O��aB�G�EYt�2E�$8VdD�"OT�J��
�)v������K��E0��'��U(�0O�-A�M#sX��l��E�"TK�"OdBf Ҙ�z�P��U:�Z��E�	�x5=0�S9	!�e�˖m4	`m�E��C�"k��嘽�*���Qw;p6�!�� ��{���iԞl �G/~z����=�J�	�'jf%���5�1
 -�aj�O��)u I8��=%���u�P���/mYV�	��hX����@�S���C�;O�x
愗"S��hY/Y�y��6(]�%�m�V�*�@f���HO�9酢[��h��E%�&�PQ5��1s� �BD"O��4�E (Z(�r�$h�õ�'�\
���ӤY�X B`��]A.��k�9�dH�ȓ|c�m�7.`6�ቓ�g�9��i��93<����*�2���ȓV��a�� ��D��$�f�
7|��TA�Р�֞\��g
w	�D�����Pa��V� ɤ��,�<���0�6���d�L�#e\*-�Y��W��b�Ζ�\��J&2�T$�ȓT[,t��b� ^����)��� ��~"ZHE��\�|x�Й7�,l�ȓ>O�d�f��$aJ�bd��@�l���f��f��%b^�rVIźl��܇ȓ?Ix9a�H-'@*S�8N�Y���zI��=P�H0�Q�G���\`��r�G\;�@��׏p��ن�c� �؂�=����yHB���B��	rfϟ|��Ȼ4�ˊ��U�����B�TJ<�� ��	�ȓ=u*|X��"*[Z�"�a��OJ�ȓ�XQ�Ɗ)�U褠Z�Kl���7RD)w�B���Ur�G-ON�fHY�Oe��S���1�K��0>��̾q~�2�'� V
�����j��\	1)��-J� ۿ��?��(��8�j�8��H���P�C^����c�FIyr �Rv%��oN�#@���dK��y7���[�æ�ޮ�x��m�yR�Дi��l�Gh�*�VEcC��� m���͕{���B�.T65�8�sjЕh��|���+��)�ʼ{ �ިA&�����G��m���Q��?z6�j�iS�0P L��](6珙j�D�g�
� ���/Yav�ɶA�6zS�830�́��c�Ѳ!
�	)��j4��L���r�N;�	�Wh�AKe�H��
�,9#%�\7#]"t��hѴ5&�̓��R��,#vƁ3�Qs�L>l�~Y��'�}�� G����@`FU����jQ�*hL �N�Obi5��j� U���Ǆ���ذ%�
��-����-<o�"�9�߀zP�����e�<q �[%�~�ƨ
9/؆�/�#���)"���d����m��)��
��%�j�i�˸-��4�X���Q�*ͼP��Eہ�˶�(��"�O�0�НA�<{ݴ|N�L!���&"۔�i��F~K�`��H'���1⍉u�b ��$U��Y���^Dp��2�͢gB���u%��O�O�4�6�H�=����DˈHQ�K�n/�؛è��v<8x�g�Hr�4 @3j	�x��C�Ã�|�LpW���=	�bN��vD�S瀃t�ĘpQ�R)��Aa��9t����a1����rL�s���u�ȄH!���Q-k��� nН�Ӏ�L�&DA��>tN!��5_
�)��B?ULQ{v�ӃY(��3#�d�*��s��O<5���?5Z��)I}Zw�T���� 8	t(u���T�Y�,S���D�>Pz�(���#�y��	�al��dI�J����D@��n���ƍI�Lؑ���<��`i� ����=���q
�el�(Ö��(?�qO�}�4U��7z�I�4��Y��7��>\1�X��YS�:��"%�!�d�)F�r|��JѮ,���R���ZD�|� �뾬2�Gw�ӗ��.Ū,����ؚG�f3���L�!�	;�J�鏤e��ȗ`����	`#�#��@�O|5Q��ǐB>���� ��B��/#F¶�ըߪA��'����>�2#M�*�X8g'� B�
1�rh� ��O� pq0�'=���N�v��0��/T��8��^t��%G�5�?y�lS/8�Bֆ�%kP��aF�H�<w��}�����دPdp;��}�'���W��P�O�%IN&$
,@ e��+6��u��'�!�E�?Bm8eˍ� ���	�'p���}ֺI��j��rsr��
�'�����R.�X9C�d�Ge��K
�'�2��t��,(�
������:�Ts*O��#���Ƹ�(�^��VÉ��Y"t*�,;m�X	"OH�8���8,#��d�5��څ^�!�sfݴ
;����
�0��� ��x�ACQ�c��}B͏�b��p)���*��tò&��g. ��lf�dV�+��p��ɏkxέ��Aߤ1�K�x˨�Y��<���ˆ��d�r*F|���2���[��^9��j��X!@Q!�dN>_�6�1#M˙V�"%�2� C���Շ?c�q�jܥGV�D`(��5� (��U�4��­}%P;�$L(�y�S4O���g�.y�dy�,�(>M�T�P�|B���M���`���hO���5�J�۵o�.���s7�'�6���/ݒ{�H���5U4���0y�~5��#�*:V�A�%M�� HEL�^-ҩq�c�"[D��aE�,�1�n�1�����L�s/F��+�*h��
C#(\�wk]��q��D�\��y˓w04y(�J#3�9"�%\�xI~x`G������#_!W�=�ׄ�G�O>:���	Ǔr�j<IRH�i��ta� �1z,9�OXQ��$"hX��6���RaaU$R��A�a��d��\��]/�.>~��h������i�m V�	�R��ҨL��|���Q$a�a|򇓯,�2!�wA�� 
��m�15�i��D�T?^I�f��2{ڬk�n�JQPLhՓ>�f=���7a.}�6D�8#�0}���АFe�"<�(̚jg�p����wMxA�2��!��i;�:TeH��8�$!it��
�R�'sUh����O<��A J�Ș$&°A"�����h �D���On4$���B�i��|��-A�n[�H:ay�q�Wk۬#4��k2&���D�
54!�`'.6��S�K�|�H�8pC��s�"Ê�0"��������A�Ƥ�J����A�+���b�h�d@�<�B��S;��K5���DT(9k�GČdD8�R�^�b_�PiЅS�uyL�p6�A +��) ֕>�����Y��'>2��Ή���1p��#"%��8&�!�c �&΋��	��#'��V A�1k�Dj��iR�qFߎu���Ⰾ�d���?�na[e�]z�3�	%}Y
<p&oH�n܅��F��	=�6����٦B�3��Xr��K��8(�,>��I�<p��/1����G,R!�(l�wW.<���<d�9�
�oc� jB-ԮZ��t�c�M�Q���v�H!$�H��em�׺k3DT+C���)r()}Zc):D �.�7���jt�� ��uI
� ��yQ�"C`���P5�w�ތQb%�("z�=�4�
T�`p��"Y��*J>y�M� \������ $�o>�)��R
x��Pd��
A0�!���"ZJ�ۉF���$c֢(%|�V+�*�~ţ�@&V#1O|ͳ� ���p<���C�j�C�0Z�d,(6�Iyb'L�T�ji�'#��"��v!p(Ad��|�ٹ$N�u�B�	�d�� �A
H-V�He�(��B�I�21y�0f'�Hi����z�2C�	�6�<Xq��	��Zv��2u$�B��$0St��e��Vip����݈HւB��=��\�$%z��֝c�B��� ��F�"��i���-ԸC䉤t��0��o�ܸ¢��6�B��:lɂ�)0� ����f�s�bB��78z`}��C�A����zLB�;T�3ƥ�P怔��BN�v.�C��5˦�aE� v�F���$ʕB�B�	���Xx��\�I�j8&�\)žC�8R�]���#X|T��R�I�C�1Zz�CDM� ,����S=3�C�ɲu���t�U��T0��QP�C䉃,Dt� B��f�������2)��B�ɥ1^9�Q�@�:k�-yvdť	o�B�/|V*GU�o����>h��C�)� 2�ʦ��d�ā�˿xBp"OZu�&&ײW/�Q�	CBT$�A"O`,�r���}��C��CoT��D"O�,z��[#1� �2fP�T&���3"O>41P�Y�@����%�ę0eK�"O���D	����kFꉃN���"O�YM�7x� H��@�5 ʱ8�"O� YRD����`��'W(\���"Of��6#M�B�ԁ� f���S"OP�
�lO/u^9ң&�u��aX�"O�9��[�!�L��A�8��鹣"O*KF���f��dR*
����T"O�
�
ÿ&k�MhD�O���࢒"O���S��vԪ�*�cGeن���"O,4�3�J/=r�R����C�@��r"O��� �V)Z�(I۱"O�M�̭�"O�Pӵi�x�Bh2^�Wʚ��"O� a�&�%{�n1x%.�{����D"O"xZ!��L�V�P/<����1"O��r��[�� �n��,R "O@u��6C�Q9� �M�Zy"O�pz��_T`y�e.T_��(� "O$��E�R&�d9���4nT���"O@�#r�9}*��� V�nE6\&"O.��WE�:<��Xð�G�yf���"O~� t��(6Tx<pD�
yFd�"O������
;x���*K9t���"Oִ!T >���U�wM�Y"O������Lx�:��!a��Y�"OQtgY�w��o�;>��Pg"O�Y2���o$�� ��ǔ�P@"O�\hw�Ӑz��@��N��i�Ll
�"O����i�'u�8l�d�F*trd"OA�0 � I��9i�ʐ0.�=��"O4Y9U�C(Cn�j���"O�\����)�������Al=B"O2�J-4;%���KN��3"O���'�	vz�afI�p��je"Oݫ�+���mP�	�ѾeA�"O>��CKH�V���U���t�ūa"O�  ��(><��p fܻi����"OL\���.�� �c�3�.M��"O�M�����8�r��ǀE���� "Oh}:$"�I� �" O�C��L�"OT0Y$�*m����#�F�Z�J�t"O&���l��b0(X�Y_m��٧ˋI�<��Ţj7��ą��!w�QZC�r�<��?\��i�T��p�L�Phm�<�@�0� �k%LD^�轰R"i�<���:@� ]���<����O�<�"M�-�L��L���!���P�<y��\N�5�R�@������RQ�<A/�O-"�I7ҟ9Jj��.�H�<Yl��X�R�C&βP��شER�<V��[ 81�1F�|ސ��(�I�<AՏ����� `ϡG4e�"�JE�<�*�ݠ "A��))�$�F�MF�<q�-�m�dHk�̎��8�v�H�<�F�B��Vm8`��cU���f�D�<)W#@'IK�@�&w��(��͏}�<���P:;��qZ�!]�F� ��Ҁ��<��荾?��|h��a��=��u�<��!�)�h�[��Ό]T�t#�	p�<Al�<x���g�� =��r�OZ�<�  ���!��"|��kuGηD�|86"O0LҲ'�1`�<̻2e��x2�d"O(���d�T�Qⱦݴ8��:"O��Y��2;��ᆇ"]<��PP"Ot�`�o	�Fh�9�%�0{'�!"�"O������.]� �3�J:ڝ��"O Q�cT&	�&���T:�HR"Ob���A�n4�U#�!?#>:1�U"O}y%�ޟ�䄉w��85�ç"O4y�n 0�t�K�&N735����"O����tV��F��W"��Q"O�%����'b�����&"X�j�"O&�Ұ�^�Z�@D�6�\6HJ R""OP��V��%d��B��/.���"O�����<D?P\2'HO����e�<A��H�I6��f�Q�U҃�a�<q�F�4�*�J�k�B�D!��[�<9Po5x��a̢S$�Q��Y�<	aK�|ݖ(�P
��t� a[�<Y�O LW�822�q��CQ�	T�<���2%G~���)ڠY��U����y�<a�S'�8UAЁZ���P�w�<9�M��$�h����e�R)�ҩGs�<1`Z+g��M��
nT��Aq�<�v%Z
�.�Bd�M	&��Tk��_l�<	�i�`ͫì̒:�٢'��m�<1�EI�/&��
��IGF $be��\�<�Z����+��}�d�av*@Z�<��!@{G�|�S�� 5���QP�<Q�,(u]�M��h/�����J�<A��:AI�#V��D��F�A�<�R��*rC�x�E�h/���dIu�<i��0��"B��W�s�<��C�k�,ȃ�I�'����A�<9І͍n.@��[-�� Ha�<��I�g���&�N?(4���K]�<�����9B�Đ� q�T�̟f�<a��޼=-2�10'E2v20�B�GTT�<�qˆ�b���D�4D((:F.�P�<�WT�m��=�7&E5Qq���@�I�<I��ǧ	j��"���N��3B�n�<�%,�tqk��Í~�(��̄i?��ۛ|l��e�Ƚf$N���M�3F��� �@7|q�
�5n�a|��ÑU��a;�f��Q�I�"a�����=G�<�s5�.���@;P�܍V^�l��Js'�xV�Ո]8��MB<�!h��T�u刉��K�/����#~ޙ�%��`�	��>T�@!$�?D���k$U�~�rs�?i��+��X
l��m����6K��æO��Ci���F+$T�t�Z3�LjS<�~��r�F$J���fې����'l��P@Z"nz�m�4=��	�B�=����%� ��X���ݰ.����H�KR
�i�ɴ=���⎛��'��u���[
�X�V�	H}�ဨk
���@�����
䭝<��v�[�~n]1�S/�6t�kF/��$�&�:��B*�5K�n���I�
�ִ��̋"�H�b��A�.���p�L�Ʋ<1�'�l���I��ؠ�aL�$�F�ZRK@�(���Xc0�]��ȤG�(-q%"e�>���'Nb�� ��~�@��)�#�(e�G�W<
o���a��~�R� ".�5}Az�� x�h��i��,q��;�Z���U9v"GloV�	��s�xY����x�^6�?�`���-Q;!��H�4k	NԊ<����	?��#�ϥM�H���=�t��#m�z�)� ��7��=���sU�/8���?�EgB�]X!��/�O�g��'[x&D�5%g8y��Ə8Gٜ�C����R<�%&��ii�#4��8'�|��EE�-��E8@G�x�TI\)*�T �*^���ɇH�ȉ��� @�)���8AF�l�$��()�T ��"�h10�%/iZ �C�ާaE�M��">TX1b�A�!h@���#T�9�|$�C�&^��+�?�ck�� ;\P1B%#m�i��X�w�T+Fۢ�P��9b�`�G��i0�}�����mWL�pҩ5���;��̈l��4��e�=.�J+O�N̓n]T#<i$⁃Wj9!�"V�av�BW�B~��l2�'֨s�:�C�� ƠZ��F���sƎ��Љ5"O
<b�H���̠&��:`���9���Q�3͂%d"��H��X��m�-Qh�+h����G"O
P"�IT4M@�P�s��Z�ۣ,�$f�Pm�dD�e�9�g?yQ$%�������%�|��C�z�<y5'J�:�4)D��ts�"����#�S�Fȉ���'Xx�P0 �.U^Tڃ�T��i���B��pΛ��?�WmLl�`��˔<t �n�^�<�`
�5%�=A7��}*�]��*�R�'�6$�@J�u�O><I��o�\_�Ȋa΀�Cb֕�
�'�b�т�
M���+A&U'��0
�'i���.� $D$����L!	�'w�%��LW�
N�+��	t���'���a4�P�h&�!R'L��cF�R�'��p�ՉB�|��3wH\:Fe�8��'�Ҁ@ӏ�9��*aȔ8-�m�	�'1*��W.��f���P&�"g��{	�'^)���:1�İ���8^�����'��Q#D��<0����"Jsd,[�'9�Ȧ$H��#"�ӔFe�Ѻ�'3�P�P��]�n-s�HT�4���
�'* ���*r2i�Aˡ+6!3
�'�H��H��Qwz�a���%Td$*	�'Yt��7Dۦ?mFy��h؜E����'>�$�gı#(�h�ԧ�}r�a
�'����M��V��	k4h��:����'H�!8��)������o�iK�y�C�n�m��I�u��t��O�C��@c���"9���ͮw���a�,�'/`8�S��7TϚ1Sˑ4�0C�	�f�L�`Ɓ&͈l�����Q�"?���چ0	:�@fD;�		�k�,��ET� ���8�!�D�w1@�����Wg$Q�v�'Y:�	�2:�j��C��S�O��Pa�ŢG��\Zè�)�)��'���Kth�/y ���Mގ���钝>tc�������}�� Ҝh� N76�Db��?�e�G�M�5�Z?O2�cBa[�SSxH�GL[&[����R.	��yu��)P�4g,E]��xaplΨ*�P!������8b�P�c���,�1�'�)�yR�� ~�쒖n%	|p�`��-��$�5w�0u�#�E2��)�'J�.1�
F)0¤X��I(T@����bB���0w�y�h�=q���0N�h�P�)}�^U�I|�>ᶦ�t_d�B�/�h��1hDO؟�ȡm̭0F�4�l�kKv�;u�	�P\�h@��ϲ����.�2���h��$��f����O�x��>G]���O~�!D�>�bH�%n�$�h�G�<�����<"a(�#���q[�Q|y��v�Lh ם|��	��l�<J���#�t]�G���k�!��y����������� �L;-1O��� �̻�p<�OWL3��aC.A(e�(���X�<UB54�"��f%;Ť��S�^�<�s��Y]���P�
"E#���3�l�<	a�'p6Ș��^#w�ޙ�N�Q�<�+�,gm�T��燷� ���[T�<�ǍEH�!��&P�[����QN�<�O��ϖ|��)�/{�����CL�<�I�МB��V�?*����(	`�<	g)��1�Ɓ����<���J���K�<q�/�0R9.u{��46Pb�"�A�<������������q�fz�<���ȣ l�Z��.O@\�`��}�<0,9�:�km�$\$X�%��B�<�k��}��!AX%bcN9��
�F�<���L'6ɠ�ud]!K%$���y�<���V��A���:P�q�b"�u�<� (|C㤜:/M�`oƖXC&]
�"O����̂��DI�.��L�e"O�ܡ��"1r��$�l�ڨhb"O� ���6@�uKM�*�l�S@"O����@�4�ȕ�A����]:s"OZY�'YA�%��E�:.�@D��"On�z��όD�Haj��8�V��"O`E�J�%U�Ω��Ε��uIS"O�R�d+�!yP`�θ��"O (�Q-&���3WF��s����"O\�#"	Z7I7�4�`�G���p�"O��������!�n�@�P I�"Oa���sM`�	�m ���T"Odt�3� ,DEM����4r�Z帒"O�UPUHX�Lvl�tR7~��0"Oh�	��TV���E�ڀ^�J�0"O�`��m�n0IT�W)84�R"ORD�G	
� 5�C6�A #���"O !x�-��!ˤ$
�C ����"O�ȃR� �8�\(Qk�=i�\[Q"Op�.7k����)\: �����"O�pA��܏0�fT��I�&b8��"O�l@C�La��*�n�,��ae"O���oO�!1�y1U�
����`"O��Q1�Q�-��AVl�k�]p5"O�0Y���a���4�\�"뾨��"O��(�'H�Mx��!�+;]3����"O\�a3鍔+���,�H��4��"O�@��$L(�`�Ȱꆜp�X���"O(@An˳9u!�)b{��F"O��7%U�<��B)|x,d"OZ ��[�l(����͍}T�iB"O���LȳVBHkU凓n)|��"OT���&BlΩ��$�d+��2"O���AR�/�` p펼�̀�"O��+p��Tf��'�� M�E"O<�!/V�M�� �$4�F)��"O@����SY�A!�Α�6���R"O:l�@#Z={�D��2-K/n�P(*O�m� *ϋ-�H��6�\5t�LdHӓu+�Q�N�9Q),��B�(��PN�C����&N.m6��ȓ`�4�H�&#W,݃��_�m�ȓtn�C��̚"�U��%�57�~8��<b�)*�Y��A��%�0LB��䪐9q�^�K��;@��+>��ф�m�51PE0q�����$.�ԇ��*��#<�P.&&�2;~<#�j� c��@Gf�}�Q>��O���+�	_-L�6���ܯLƦ���{r��cRV̇��,j`�aeI>�b�#aL� F&��'}��RW�ؚA�N8�'`�O)B��>sb}y���Tt���j�4�?�#�G�@UǊ )���)�>:�L���3T|Ѐ��?8qN����m|4Ke�G�8+��ק蟶�����6u��)�0O��Pn�d�Pe���h[�j���S�O�p��+GF%X7h�"��#�t��&Hk≒0Fa��oŉGI��C����=�d5rT��6L�T��'��5��#jǴeF�ܴ%����	��NP����~���N�ΑxҠ�NW���(O�>%xsE [p��w��*qv�<HQ�K7VTh�%Ǐ|6~�g�l��ym:�'}BF �$۹(fz��dG�x��D�7DD�:A���b�� Ot ���	T��,�S]پ�C��ЕX����Ǉ,}��م��=>Y�E�ϞK}~���)�^`�w���,3���G��u)~	B��zv���"�ڻ~�.4S� 5�>�$s�-Z�B����|��t��-�3�"%+Ͱ�j��Q�r�B�'B��i�Y6��wJ�"��N(�t�u�ػq�&$�=E�4憡 �3C�˚0�4��#Jbl��1�Ie��~��(����_)+vi{!Ҭ�y��ߦۚ%�ՆC�$6��k�c��y
� ڑ�c#�^���D��q�RP)�"O����n��񑌀%-�l%RQ"O���E�+PJ�E�F�8ي�@�"O,�����/ެĻ�/\�]μP�"OL�0��_)}���4.ӜK�U;T"Oͩ�U��R��R.Z�Y���e"O��s���U$������ͱ`"OJU�P'���� �ԟ��P"O�H��S�1�9�g��"���R�"O@	ے-șU!^�xs�C�z��x�"Op�oT�5�<K��\-"x�Hj"O��k"hJ�%*0ɀ@�Zdp#�"O�0Û�b��5o�/
,(,1"O���'�B�̱0nZ�=/pE�"O����U`��ٳ�^���c�<ٰ�ϦUg�) �Ƃ�s�33k[E�<�.S(R��q2��2F�"�2cA�g�<��J�L���±%�J�A�'a�<Iu�=g��5���1, ����[�<�!m�]�tP	��
�1h|Q��d�A�<�b�
.Zi@��!���l���`Sh A�<�&�4d	L9C��2$�6�E'�}�<�Qk/i�1ER�j@5��!�p�<��C�gڊ� �NON �4�AU�<�t�Zbq����g/[r����M�<q�C����U)%�V;(Z��Kʆs�<1DlL�E[�`���8A�4\�d_s�<Y�*�]��M҃eR4ϼ9#G"Pm�<!��(���j��ڮl2ĔӶC�t�<��<.��$k��M�,��OAq�<S,�v�|��F�7t�\D��!�G�<��kԉ{S����é&p6�P��E�<��a�9��gH	����	�f�<ɓK"k�Q��0aZ�y�֊e�<�C`3(�0��� .6�.1��B�g�<���W� �@��L(#h��:��c�<I"N��N0�E�APB�&I�<ل�_ :̬�2���MF�q��a�k�<9A���4�r�Ԙv1R�M�j�<YJ�F*JD�}ߒ1�
��yr���xA���OLK�CD��y��E,��p�
�+1V��2c�y�m�3�%	>nx��
U|6��_�����(�5rE4�6��]ʘ؆�;3L��B�с����$"H�Y�~T�ȓG$Hݠ�E�� ��H�dǇ=R�=��~Q�H��#2�$�"��8�LІ���HH_�i�<T�@�ݚo`H�ȓ~y��C��0(;H� �"J� �ȓ\��%K���AX�l�D+�/��ȓ}L�(�KU]l�:���A����ȓgy#���ON�u�4N�Hz܅ȓ��a���'{�䅘�B�7R��p��V���j#�A,*B����A�--�̆�qZ"�PV/T�6�ܱ(��M��H�ȓ+윅"S	}T�x0���n��ȓ-~��q�o]�4mRa�G!A�@���ȓ����̋�n�Z4���>-J$�ȓB!B2���@�>q�2m;�Єȓ�@ɺD�0o¹1+��fظ��l~nPsw�҄Z�<�E� �W���g� 5�`���rM�D����ȓH �dÑ0ahtz��D!�����UL@�p�ꄮE�9���fB�e��S�? .Ȩ��D?}s̜���4��(�"O���q�J-Cv��$��5A^$� "O��@d�QfD���)D�r"O��{U��/!�r�3ċo1脲7"O����nϦ1�r	�(9~`[�"O��l�8��qH4BZ�	**�p"OD�)C�Ě�>��&ܹmt�v"O�!Q0��U�Xa��U�	ˌL�B"O����EX�t�PE�6��,��"O������T*p�F /ǌA+R"O�Й��ӀT`l����J4\YV"O\�r2lUL�q�#��d���	�"OFE HE]�ht�s≴6�z,�"O����׃l�|��b����� �"O�1�OS�2��4��X���"On���>`�r`b���~E����"ONU�TA��F��qI�`�<cA��@D"O��D*��l+�DJ�o�%m�n�b�"O��"	�S�K�2�칀�"O"�hG��. �p<bf�5ox��2!"O2�BD�G�&�V��b,[m��Y6"OXXA:`�KG�@:-����*O~5��OŹC�r���;g�����'}������0�W���_�1��'6�(UKC3TY�ɷ��U0͑�'6��#��?|��GP���;�'%DM��4a��0yWG�CGd��'m�RA�ʕ��!�� ��e��q��'#���4B�O���󰭘�^�8`A
�'�����f\+2����аB�*G�YQ�<� f�*,y蕨�g���Jt�<��"�(-4��U	��;[�-\�<)���|LZ��M���Ēn�<��@�0��bg�e�ؓ%Kg�<Ie-�
T�$�q�Dٯ5O�dF�[�<��b�T2w����X2g��U�<a�/��a���RX��@P&�S�<Y�j�31'a�3�޼fS�`H�j�<	tm�L��� �&	���@�b�f�<Ѱ��(X� �yU뉪A)p���\h�<�Q�ÈK&d"��F*/Y�-�E�Ap�<IE7ibA��n�ҼaCEl�<�Rd�s���v��"�P4x�(Uf�<Y'���V�Kh�
L��%J�d�<��I����j�B׽`nR��rf�K�<A�6�\���
�:��pYr%�@�<Y�g^:D�$2�]�;j�p���~�<I'R0!��I1��M�N�ӓF�s�<�	Bu��S�O��r�]��FI�<ɲ!�n2X0��|u C�oXH�<��Ț�2��ٳ��'Ub̴ʁ��F�<ɷ�J�+-��y@��"&d�q:���E�<	t�
Zr��5�U�(���D�<���>���'�:�)3�ID�<i��H�|���+`�/0�R���|�<����R��X ���p-��22ME|�<IpD�M�TYz5!�z�P��#��{�<�4�`�8���_7H�I�D�Bw�<!�)>�݈��G�T��#��Dp�<y�/(��t��!�pȱ�+�a�<Y'@�4<�!hR�E�TX�)B�Ob�<����;j}�(*�T�(�2��D�<������h�h��C;	���X�@�A�<	�A�6�v��T� �Dp��O�z�<� J��&X�,��|��e��C��D#"O��XP�K>7*j)�e����8�"O��b�䂺.	*4 �
�|��A�"Ob0��
����)sC��F�튲"O�%(�E�t�6aW�R��rs"O~)�Ш ���{��	"�2 "O<�����a`D� IѻodQ��"O���b���$�P�U1��e�C"O���G��z��3�I r���"O�X`� ����UJ3'��ѵ"O����R�5RaӇ�=x
�ً�"O͙�.Ť� ��fD�=�I�"O`����!,�^��3�C���"O�]�u��?5ԙr�e�I��q��"O؅�`�=fu� ���KR�x�"O�E�҄
�vOd�I��Q/3L���"O����&�7Z�0%$ן~&�u"OzY��F�?f���Lә!��3�"O�4��Ԏ)�lx�����0�7"O�a���T==��$	`H�v���#"ORd�D#2
��|�F��jp�T@A"O�a�֌�y�r���/HX4؈�"O*=qe�\SF�}���W�1V �q�"ONt�?<�6��bd]fn��0�"OfH��Ŝ�;\,(�!�("�&��%"O� �LW�%��ئ��D���c�"O訉�g	��ݰ�l�+H`� "O�X�l�4��`D-�.	پ�{ "O�T15ϖ�8>2���ڒF�69�P"OF5�Fm�'_8>��3cV$���"O4� ���EJ��K�;�c�"O��ر�Z,Hv��F��= ��X�f"O<����֒B�va�K9l��M["O�rp"�7��a��4"����"O4(���
o���D7j���"�"O�a�L��XT�#�نP���"O�qb�\�O=��K 8���"O�x3��u�V���@�f${W"O�I`-�1!|��(�.O�X��\j"O
U���9|����J����"O�Qw�)���
<GI(�V"O�����"��Py��Z�b9��"OX��s�ʿdF^��B�	�av�d"O��S��X�������-'�~�sF"O�u㕀�|x��3����!:�"O��r���7F�]�d/�'��`q"O�X���^�Y�*9��QM��{�"O�� ��BwK��Z5h�	J���"O� ڢ�o�T�Ȍ2�!�"O����n^��8$f�4��e{B"O<���'�H<xHy��ρѰQ{F"O��ZL�+u`H�Gk����"O�����ð��\�@�"�&d�"O&9AS�]�1}2`{��I�-�L��"OP��tf@ .��ktH�&i���"O~��4ֲ`؂e.��р"O�Z�䋰E�8�Y�_,����#"O�i�g��D p!y������1�"O0��޺2�=�����"O��X%`\D�pbHNv
h8�"O�U�U��p=���D �2k�LRC"O���A��O��M�tfP<sn��"O��^�H*�-��C�O� �I�"O�e��̞�6~x����R	����"O� J�®K�o�J����"a����"O��X�@Ӥ���AEvn���#"OF�`"o��_����c�9%��Iq�"O�Ii7��I�T�7�0I"m�"O.�B���8=x� ���;IJ �""Oqs�	   �P   
  �  u     �(  �0  97  |=  �C  J  ]P  �V  �\  @c  �i  �o  v  I|  �   `� u�	����Zv)C�'ll\�0�Ez+�⟈m��e���+gR��D�Ԭ0h�� p"�e`�o�ݑ_	n�R� -�H��ՁU�Jp\�@��!Z�矀�Y����TT�C�C9|>ԉ4�ϲEd|��J�a�����#�/����	
t!`Iӥ���@$�4���Zx��4fܠq�N����5D0����P�S�����'6F���I�!C��x�b�y�B`���O��d�O����OZ��Ea�[\��r@�ɔ>��Q��Oj��˗x� DmZ\y"�'-6�3`�>���\� (;��ylȂ�'�Zā��?9�V�<�'f�aR��?�'r&ҦG������33s�`AנC�a��B?O�H�,�t��U(��� n�X�A^��ϓ��'��}(�#y�ɘmdn�!���+���B$ŀ�-���d�O>�d�O.��OZ�D�O��'�y'Il(�B4��(yR��BR��?�C�i��DlӢ�l�ܱ֟۴ol��nl�t�n�П:�Mˡtw\
0F��UL�ܠw��HOn<�����} !
`�4U��(�@k ��!�	�E@�S�o���mZ�M�S�i��T�rݥwGM�
�<��
S�:�Rݢqi�}���w���MKE�;��LєL��C���J� GF��c���A޴w����e�bP!D*���£�,k ���i�+J��9S�ކ)=:�n���M���ii4=p�ǉ���Ma*��Mk�E*k����	5	�H���M0UN���@��P�<�� hk�L�m���M��u��|p�' Cߤ�ru��^�&��_(r�KԒ*�0	���M3��Xy���a�2i@���3����d�
���än��4Δ��Vƒ.{��;%�9(��=����?1������0�ޱ:fc֮���MDU�4K���ԃ��$@r	�'��XڦD\ M�p�B�?̝s�'�n�c�A�*9� x���9�Ό��'txMS��[��ġ�-�$,�8`�' JqIB�Ԗ�p�)�>�7"O\��"�ǉx��e�D�N�n�j��퉉h�H�~R��Ї�@l�F�?iV�l3A��t�<���"��qa`�%$�Z�
 �r�<�VI[�=h��5�M35�����Sr�<����P ���@R���SRD�<�S)�c�d�$��NQ,�"i�<�r��d�|*�D�5r�ցM�<�A 8�S�O��ˢn���\��C�FN
�"OH9CR	�)���P���JFl�i&"O�X��R
]��qd��3P4�"O����^�<�A#��# "O,��(�/I|�10f� 9�^$�""OD!R� ĉC˨��C��s�H��w]��X�-4�O�ȱ�G*(�� e����"Oq�Ro�Mx��� �2l���C'"O�9�2.�����)_�L媵"O>�
W$�"jو Yfm�?\����"O��;VD��PJ���JƐyFP�I��'���X�*fӄ�fd&�R���[R�=�m�3
�	ly"�'F�'��1bb�{���0��v�V7-`�>� &�c�d��0����E�'%E&H1
v�*�8j��i���&�s��:4�
IM�X���@��KO(��'��6-�O28��Kѯm4�b�)Wm2�&lyr�i�2����g%�A�!ɢ��P��d%x�ւ���(�'1�I^���dG�O0��+�t�T8u��3l)J�X��'9�	A�l����'���'��W;XLӢ��'C�8�"�AT�8��	#u����f��Ӕz�����:Ԗm`D���I��Tcn����$�)§AՎ��O}Hz��bG��I.���'������?�N~2��ԏ�
.0���a��5E=Ĝ:Ć_���?i�yN�\��ʌ�X\jԎҙ<���F��(�'6B�[��Ǫ`�fR!��'��"�4�?I-O�<�/���#>� -ʺ\h����F-�<`�m�-�x�۴�?y 	�=�p�!,�Q� 2TD_�4�vT�u���	���P�*y->�PLH5db���ç�c>��,?q�������D<E�������MGS�$���O�b>��O����;[tћ�,�b�� IP/ˣ^(��d�O ��?ъ�L���@�0��x􋀶(�zlS��<���i$�7'�4�
�ɠ<�DV�O�Ѣ!ɻ1��� х��&���͓�0>q$��>q?r����N���1� cU�E�܄��RP�(�U�	I�H�A�M�B��c2�CR<�G�K�-�Ӈ-5P	��n�%f��I��?1Dkٳ!B�(P�p�,��(M{�<��(ӱ=�ܝ�2KSNzAw��y��MJ>0o x��O-�E�C��TqI�V�fv��������O��D�O��h%Nc|a��iT�K��		U�#� ����ݚE*AQ��9;�@#�^����;���ܗ:KB�3�	؄F���P��� ��{ �^	��O%�&�'�����٣�F�CtV��#��= Ә)H�#�$�O���D�$<��� /� i����	>����O��)׋�Gk(��^*Wx�P��'��IznD�ش��'���Oxa*���"T�(IZ0�@cǸ4`�%�OJ��P04�֔Pun�&��[ǡ	�h����~"Q�̫)�"=(րߖG�� ��C>?�b�Ϥ��p�%�՗ ��~���?�B�IJ�TK~)�5
P4=��]�v� ?i�kT��,��X�Or�[%�*��Rݪ'|Q��6Z!�D�<Wm�����&v��T��.zџH����	�O�H`��ʋ
Bmf�Za߀Lg�6�OD���O�5xRl���*���O���O��]�Zx��g��L��A�aW7+�4����N6mX�G�m��ұ�.�SH�I�,�Lգw�{-�h8���#j�@|�C-� M�ڬ!�F	R����5�)�SR��j^:8Q�GQ<$:r|[��UaL��:?��(W��	4�?�pGǘ���n��I�d��ybi�����A�cR*
�lu
�����q���T�'��ɊI���z#�Q�}U��#�H]3=���҃����	����Iky���+�z�>A�"g���J��5�΅(�k�4��Ҕ^�q��k1�M4("Q�P.0Rd×#��x��_4$���0����+v<@��|��B��5ʓ'�\��5�A�@��& �Yd��w#M������`�?Q��	?$WxExU�]p�SHܳZ�!�d	���ȧ�Y�U �,���;Z��'�7��O��KoN��6X?���  �8��0Y�1tMĴu#����ȟ�y�Pܟx���|����Q�L} wo�.GM:���H��JQ!�B`j�2����@���D��u�1�d���ġ�L��߶4#�\8=i���*܉hDTK��&�q�������'�&��d�D���,S�M�)�vbO>����0=I����YAG!�¬���u�����o2�4���^$�3dNʉp��	Ey�h�*#6M�O:��|�R
��?�$��F\`�7h2���K��?��	U|��E��H�\����g�����V?��O�ⱪ���U�b�E+��y��k�O4I�[!�2�{%��'Fe 0{��4�S%Hr]����jQ�1�aZ7u�T�:ע4��Ɵ�E���'�(l�-D1���T	S9k���D"O
أ7�N,	�H<�'L�� ��&�	�h��H���F4oo�܀v}5D���jlӾ��O�Ĝ�LfIPSG�O~���O��d��ArD�"�h�8�!ȧW�.)rRN>~\)Q�O���V9�1�1O��#\)"jMR �A�2� �)� W����$�O��i�+3�1�1O|`�d�f�V�jV�ν/���5-e�vЗ'p�}1�����'��'K|q	T�,(`���9����w"O�)��MK[�xP�Q�(e�IW�����dKD}���l��ݡ �Mq�"�f�0 gi�<��*^t8�� g�+Ւ�*fʄ���rGO9D�t�A��@2��4"�1TWt��,D�*$c� t�4)�c�?i01��++D���q��J�X�)�K�Sf>D���P0
����(Ȍw��wA<�O�:��OT�rbf��q.�B�۠jy���"Oj$�5��5Ҹ`��MD�gl��7"O�I�%��&���̞N���!e"O��rfǂ)u�X�!^��lĉ "O� �v�A
��Ӵ/�~� 9`�"O�$S����f:Ι`5�����I���)Y6*�~�R���M�pB�2Lz�]�d%j�<i���
F�����-�-A��U���f�<ѓ���P�V���*T�19M�F�<�P�ݪju���ԅ�O&�X'/�A�<��"�-c;&`�`#D#l0�aӉ�C�<��(�+!$�) ˰H:�(�ß�J�-�S�O[6��"��*`�D �WiA�Y�Ό��"ON��o �@v
	9�g	f�Y�"O2A{.�!9:�����'kQ���"O���BU�m�P	��$7<tEA"O%�ӈ����9��9�"`�S"O�,Ҥ��^3���ɬ(uf��3V�0��� �O�Y�%)\W���:�A�>�$h�"O� ���䄢Q�te�pj�	^����"O����Cn��������� "O��JDH�w/��2��תo���`"O����S nR�1��������'~�`�'b<���Q�>�����-(��LB�'��P��	@ղ�R�$��p)��j�' 6e��則K��@�G`R�}��%Q�'�b�B�'xT���U���b�'��I�����D����'� (�
�'z���b@k�8�Qt�^�)9_�'�
����&� M�F$H�N$�􉒟6�!���/�P=k�]� a��Q�ǘ�K�!��˵stI�fB�_C���ġK�!��E�qOr�[#���G�5����Y`!�d�xk\�w� /�-j�W�Z!�Q�V�$13�o:]�� �4��s���͌�O?���(-��R6mo0��Ph�<7�U�rp~ܻ�KT�e��C��z�<����Xj���oI�A�q4�k�<��Gʯ7lp(�t�,W�fl��KOe�<1�ꔻ1q�i��ɩ,�*$+R�	y�<y�)��Vؔp˄@-~�J�P��NNy2�̵�p>a �ƒ
V8Y1)_'(�8�ԏS�<�A�	+��4Ab�Ҩ:``��VX�<S&�t�R�!�]'/*9����R�<�XT��F	-�����D�<9wꏫ�<�HƀU�lt�р�Bx��P&o��|3 %�8�D�P�b4*� D�\{P�)t
���d+ŴF�<�)�O3D�H�BI >���qCH�>x�g�#D��v�ަ}Q�4��䘶o�`h�&D�Dj�F��� �ģW%� `�&&D��H������CT�S���(�
#ړs�,E��B��,�`��%n�BV	2"F �y��ݬR����nFm
���d�<�y�)C� �):]�d�����ybaP�)�5Sb�ĲRZl"�H��yB�G� Hl����%6�l|�MH�y�FT��$�i�5y��9A�ă��?��/�m���� 3��K(ި`���<`��ؔ�6D�����8��6Ǚ�����&D���"/L�^�R� ���Vg�� %D��T	�1f�i���� S�pA;ń"D����L�X$�v��2JR�)B�:D�DC ��a�[r˕'hq�@�<�ÀR8�0�i�&AXr-2�@A�>�0� 5f8D���Pm׮9~l�{��_�x�h���"D�Hpt��"g**�Z���F�IH��3D���W&�O�8@1N��E[�o0D����+-?��]k�l}��o0�OL�;��O�H�%C%�@@��G�oC`i&"O�hsEH�
��Q�Ê�-H��D�S"O�.��� ����|L��c"O��GZ�)(V�ؕdD�Axh��"O��Q��!2�x��*x��Hɗ"O���G�A�3z(H�6k�,!�D̀#�I#[��~5(G]�v��g� %Q�DA�Ip�<ɧ-KITȝж.�\���A�<��N�-$޸�9P�
�jR� G�A�<I���+9����*H+tG��"i�|�<م�I�eb��3�g܁S1����S�<��H>on,$�� C(�h8K��I�)=�S�O��K#���G}`�yu�¹u��"O:�SLEO���sn�Q�^� "O� ���&S/b�I��_7S����"Oj�a��1@� |��H�/��-
�"Od��[�!R,�Bh���S"OT1I���Y�pI��-ҡ1�<}ْU�`8Ң9�OTVA^V��c����D��@�CV�<�R�ÑmS���e�L.$��ç��V�<֌�)#�j	�ʍ  '��GN�<�mC�\��s���?	�����p�<�GI6GF]co.iV�B��Ijx�4�f���d��_�&���F5�l��Q�1D��C�\���ls�i�2̂و&�-D� �5��.RD��)ę$�b�ˑ�7D���0�1 �Ē� [*\%[W�"D��b2FF�0����_�0<� 9� D����;������kH�Ē�j>����E���׸�v�h�#Mw΂\j�� �y_,ƙ2aS���{#�Q0�y�nթ_���e��+n�e��NM"�y"!M�1�S1�G�f65�"��1�y"�M�"�0��K��$��зIԗ�yRȌ:'�`�0���6mRy���!�?���t�����\�쏕�Z�0C�+�@ѥ�9D�ؒ����bd��@E�]�6+V���6D��KW,Q��LM��7h`y1�(D�h�5I*u���x���D��t�g)D��G�Z.�b�:B"��o�����,D� �2�S�=�l�m�?܂<��b�<I�k�I8�\��Y ڪ���8,�|$[�i=D�̪�c�$Q�Y���9_&(��Ջ'D��qd��3a�(<Xr?�u�1$"D��F��^���#h����$�>D��*���V�4����Ը?���k��=�OvP�6�OlЅg���Q%�º��<Y�"O���#��P�6�a�A��ĥ��"O��ԡC5.F�)℧��[�F)3�"O��BVj�S�X�ᢦ�#�X� R"O�$H���SEh��F����A�"O�ѦHO�vpq�� A�����	A�J�~�B�&.�Фp�3�)�A�v�<ѐ�	I
�U���M�_���j�h�<1�	H{>L�� 8�(�1�^d�<��l
�+B�	���s�Fq!Si�{�<ɔ��$	Z$��g�²5�и��y�<�&���L�
��DbǵE�僇���1�F?�S�O��	2c�N$wb� �ݔj꒕A'"O���nI@�p�	�J���Zq"O`�P��D</vL"��®+��X�C"O��D�mi�q{s���S�D�˦"O^�آDߥ?P���Al�p)�[T"O���� �DxhX:6�/l�H�U�Z�'�OZ���% ��x�\;@q���"O@�!���(#�6�0u�wg��G"O��8�E��w�
ʵe�D�}��"Odp���&�2��#_��xtY"O �ՂT�W� `�B�(l�TI��'`���'��K6nɀ��Z�U�r�		�'�$D��ə,ì�( �^J�����'�n�(wfߟAt$��IJ�F/na�'���!�#w�1P"E��Dsli�'J�a�V;#��=�aj٨<���q�'o4$��}��A�.4
|����rvQ?�(�*Wtji+�j�S��Tk�7D�(�4�ܟR(=H$�����dP�"(D���u�K�3���5<��z�(D�� ����߄yհ�XàH;a��4�P"O$���g��p�v�:$�?v��EI%"Ob�c�H�Z�Z�D�֏+<pD���'s�,P����_r��۲k�X`���	�?�r��ȓhF�����W�&���o�F�����O�0�CB��i$p��2� �U���ʓ=df(z`H�U� �Ac@��A�B�IeHBɒT(�<D��$ϋS�NC�	�US�]JSo�*��u#V���`��"�Tͅ�ɴRj1��� Eҥ���֗bRC�I	"�؛�̒0,�Yhr��\_�C�ɒ!i8���T�m��5�"/��>d�C�I1 f��w�1W��q����t-�C�I@i�Xc')S `�ّ5�T=g�b����v��-9�����S��l��	L�r�!�$L}�-�p(��5c�5�&��E�!��R�b�,J�q�haC3%�2p!���w�Z���(��%	�,��Ĝ�Pa!�$n:������, 	J�H��V���h��`*�g�7K�� ����Ȩ]F{��Eۨ���X���8l��j��0 �"O�hXe��&�|I��ĵ
��إ"O6��"��'�v�#F�׶I�|��"OH��a�N�ற�	ҭ!����"Or��r�30����V�+����"O�@��D�T���<T��	��'b��J���S'KS� )P��)R0!�@��І�D������	0cTZ�!"ָqO�E�ȓFA�e�bZ^+��  c"��8mzmr��#Q8��9#�cJr��
�,�"�l
�|����pI�!%Lv��ƓP��P�lO(*|^$!cNjk�ڌ ���I�L�ɚl�I����������#�,-2�y�"��0l���'���'�R�H�IXnEIҌ��Z:t����w�����'JO�iDŗ�|؊D�g%��#>y�oG��D�x�~<�ڴt�(�3���]-��
W�"�`���	�pӠlGyBmʶ�?�����O�*����N:i�r�Gw���{.Ot��DU�2�"I�pW��1/ĳu�}���<)U%�<��q��Rqа�3�d�{y�ڬeWR�'��Iw�T�'���\\���s۾��!�WR�m��D� �nUj�:Z�����ky�Z�F���U@՚}�`#_�;��FlY��yRH�:9Y.5���S�N����i�r5['�F#�O��X�u��XxcΊ�*{ج�'���Q���?9�O�OV�ɜ"FA{��� �ș�"GGSHB�Io�d����'��L�6��
i삣=���S� F��q�nґf4�A倍��9�	[y��$��'mr�'^�?y���T�^�}��X#+52]"���/?���nکL������x$,�OO�O|]A��c�J��-E%��$X�ێ`�>6-[�J��2!؏��z���2rC-}�^7:��
eo��F�`b$�	b�$ ]���'�ўxϓ���B�B5�(��W��"A�ȓsְ�'
V�\8��v+H"h)R��	/�HO��O��a��*�}�f��7�#}B�0�so�
�?Q��?�����I�)V^�Y�ҳj62�3E��wBu��"�y�����'e}�ln���O�t"w��&/�:�̂�<:L���'M�Q$D������؀@%h�8�����Q�T0q��O4]�ĥȼqS�yX�M:�b)��(�O�=����LL�`��р<^$��k�$F-!��K�:�p�2��*��u���!$�	�M�����]&�,�O��2�LP� #�uO�� �.�#ެ�b�'RHY��'���'���;���e0lx`�	�b�4�~�)Cϓ^�� ��q �ɛ�\1 FBh(�#�"�z�����bx�u��-�n�lA;��ÈOV�Q�'����\�B���#Ǝ��J�I��IF���0�ǨC2 I��k��g����"0�O�'��"�8v.�Ʌ���#RLP9,O*ms��Wަ�j�m��t�Oɬ��O����\iz L΅��I�b^�1���_�>�<���U�B�r�I$˄�ؘO�B���N�w���DA_.
|�	h�'�B)$	]#r��۳���~��U�%�' �p��'+C0�T`�d�1�|�	~�0�D�OV�S�����S�? ��[�C40x4`���;���"O�P:AAO$$�`�����;/���k5�	�ȟ*�T��2L��@LǱ,vx!8���0��$�O�����[�h.�	�O��D�O|�	�O�䓂�B�z��J%K��TU��#&����	9c��e�r��,v��g�'�$�Idc 5r4JD��t]�X�E˟�sQ"�=p,�2������I ��S��,]�1�3m�+��?[�(�Iܟ0G{�<O�t($����+gKˉ]�8�"O�P�� v�`��T:NR
5��'�#=ͧ�?�y"�qHa3�Z LL����"��?�p��I�����J�V����V�x�D�W,1D�0icF�-Ȁ��Q��;�hE�g	=D��Z�A��S��t��^}��@�&D�4K�AI�SݜՑ@�K@���9D��(��-@��!u�D�e1HY�6�c�T�ɳV�����|"��͘r�\�1����)��C�N����ߟ��I��2A- �Z~�y���	~v����|���ǆAߜA�2)�*^��r��q�'�bE�3
*�m�C'�a"��5�H�3��ߺ/�
�j���4DX\#>�������pߴl��OoX��#��&`�x��ش-OB�$=�O��J�L
6D�f�/��Ҥ�'� ˓�����X�:�BP�Ggh�0�'<¥}��$$�S{��'�����a��mgx��E�nԔ j�OĢ<���&U�`LY�]���})�cd���}s�'���z,��Եo,�PbDC*G-���t��\��'$��yK���<��CA?G��Ј%-� =���!.@�U�}y�Od�O�R��>	W���b�p˰�A�F�L���ǉ�..�l�O����h����Qj�H�cW�H�@�c��)>�~�`�>W�>��Up��P�D�@�\�Ԍb4�����&�D �?�NW��

@&�?�"��ީs�Sg풾r����E럀z7�#}�c6}l�5��I�M����ܝ) )I:�R�"V��iy���$��	�ȟ� �'�
 Np�q���Ɔ%���!��i?�c�Z�T>牮�`�	ҟih�<���b�C�j�H�ڰMަ ��I�؝�'�tG��bJ7FxH��T�R=���MG��?1�������(?��ybI��~2�[*�a�͇�y{�mj���?yq�2�O�-YA�!2�;����Y�t�d"O@`b+�6���v#�I|ڔ21�iM��vyr�'GR�|B�5�c�>ۖD0��L**a4c3� 2�M���?i-O��$�<�|n�1Ln���Y�al����Dgt�B�	-+R@��������c�
[IC�ɂ5\��aC�"~�^�RT`�Y�B�I�U��X���!'�h�#U�J:H�~B䉚fX<�I��@)1*@3"�\�*צC�	)o\((Q�I�K��g=a:nC�!־(
"�ɬ,=��R��=�B����r��c(Փ ���_�C��9-#��Z�ضF��+�B1>B䉫
(H��:b��|���:��C䉂C!X�6�*6���0d�=n� C�I*�zEJ�/Q�06zd��T�6j�C�	-0���3JF�C��e�e�ߒe����K���<Yg��צՏK�m[RJ��.�&�s��\;>.H��.ðD(�SD�	�݂" ƌz�
|�� P;O0t��#	�0v�<I(Ϊpz���ŕ�5��}á�X�8�Oّ%����"!�+f(���m��k�)$yzՆ�!w�Ƽ	�ɕ��h�I>�eFE"j�b�qv-�4>ƭ���^��X�>��b��#����iF���!_t�<�A��~`d�ԄG�2��3nNf�<9����(�#\C� �z)�E�ȓn���C!��	j��y��^�x�6�ȓM���8A
�8}{�i��dJ��z0��w��h@�w,��`���}����ȓ.�"Ur0�[�9%�up��+&���7N9�1��!��UP����y����ȓ��uPA����td܆r�:����~����S�q���IW�B�j�,�ȓ�̵9��S�%@��)C@�o��L��o=f�b]Y�\y%���Jƞ��S�? 䕨6��>e�A��[�O8�L#�"O(�S�,l�0�bb�3V&`[4"O�M�2w���7,�9� 8�"Ox�h�i�H(�t@��_,��� e"Ot4{�Q� _v�`קʁP�� h�"OhQu�Aj�v��U&�H ��&"O����m̟[
��FQ�hX�-�"O�p����B���KU���T#R"Or�`�H�_�A��*UWD�=�6"O��gQ8�А ˁ�@�m�'"O��Bî.A�QX�'��DA$"O���c�L���X�������"OhP��LJK���qI�&zp.`)f"O� +�e�3�6��t���MD0� �"Oƭ��@ͪ���w6ȍچ"O��`��̬?�K�	- *�"O�5�b.��c|��J��*$\u`6"O�Y�-Z���*T'*ڌȴ�I_�<�+ؕO=4{w��|d��	��R�<yA#Ȩ����Z�v��-�M�<q&%�2'<&�Av�A��ޥ�ʂ�<9�$�-`˒}�"A�g���E$y�<�ĒLV�R�d��/1��!��r�<ɲ˄9g<Q�T�Яi�ea�fEt�<)%iO��:�R%�*_�R	V�He�<�d�E�$R�� ��:b�`�1M`�<��K/����۽^D��r�d�<�%���L��*f�7xK�h�+I�<!�@W8|Q�
�o�,W��PүK�<Q�@Kv�RSl�6�49�E�D�<��M�:9%n�b����i�4 �Lf�<�w@+t��8qr�H�# fh��UM�<94C�hK,�ҥB>��Lt�<Pٖr�h��e��	Z�jGK�<���^�AJN���S"70���E�<	�)�E+^��t!F&f����SAW@�<S��	T�aB�k f���HIf�<�Uˏ��άq�O�$�B A$�]�<)��}At�kd�ۇ�Ɛ�)�N�<	4OB>zD�1�H�KUS��VJ�<Y�i�:[�23"`�4e2=��ZD�<�cҿ� ��Q�R�,���b�U�<��/��m�@3��� p��؄nEU�<��*��k"h�p � (�X���IQ�<1#K�_��e)G._�\����ÈJ�<�Dk��%_@�Е��~%XA�R��C�<�5ET�q� �3"�5`�h�G�<9�,�	xb9�ģK�r!���H�<���*":�q�SN�+v�X @AEH�<��KtL�m�Em�3
G����O[H�<D�S>[Z�Q�M
��Ke-Bz�<I7��
Δl4BC�T
��6hUK�<�p�9��(X3�آz��Q�@@B�<1S�S'B�	�c�9{p
��c��t�<!��\�R;�C1���~�
�nYk�<�!��Gw@-��H�N(,M�S�^r�<є)̻+6�@sÊ߂"��9J�a�n�<����%e��Ȳ2�G \������Dd�<)v�/ԛ0���i�4	$|�ȓx<*@�u�Z�
(�s�7�8����A�GC�u��9q���k�f���o�`!����f�.� RE�; 4�ȓ
�j1���ӟ?ǔ��%��'&5��_���*�[�h,^4��0���S�? �8�#���8 @��A@"O�4��0e��T��Nr���"O"A�A~�l��2��
W��4�T"O֝�6�ڒ���ǖA���yb �(�J,��傸1erl���#�y�L�3~M�I{�^�_���b0�yB�\u��B��9B�X�A���y��]�R��а2���9�d��:�y�$�4.\PR3lϦ�Ěd�U�y2�7 �j����%l��3�,Q��yr��!���N F�A9��D��yh���(�*�-ɇM�$�u�\��y�k	� e�V�W	�I8V"��y�'�+�Da��]�R�>�zT�M�y��//KD>Pm�a4g�_~Ć�X�\H�UQt�؂�ޖ}�M��/��T��ǊTׄ�[p��>0�ȓ>���a��׳��C��$�T���e��x�#,<C6�a�I��hq��8�t2bˏ()���ȅ!_�IFN9�ȓ4���F�Խ�*C�a�^t��ȓA2<ŘgI �*�����g��B�^�ȓ �ʙ��������W�������$&�2�"� c�DD�Sӑ,DT�ȓ	���F�	^�Db��Δ����X��P�Če�Լ�ˌX���ȓ5�>ՠ��L �d0�%aEX�,)��H%��q�Aˢ�IF>b4┅�&Ā�sī�=�6�¤"L<C_�|�ȓ+���y�� Sf�J��A���؆ȓ!���q@��	�q�7	#6,�цȓ: ́���K��p� ֟~�
���-�jQa�A@�m�Jׯ�qRT���,�`�`�i��D٣�2�I��r��2���!\)ᠪցT䰅ȓN��Z�v��mK J(�>]��#�`!;�A�yˎ�2��#,�$���pܩC�ڊv�X驇I�&�����x5���%V����O��Y�",��F�.����
��U��O�e�xQ��1�rСa�J�K��/n�25D�lrf]?uK�AȦ�\�kJ�i%D���D�w�� �ٕs/�à$D�p�����r�.a��)=_�L���,D�D(�μW=�!N�4
��* D�8���6��T�(z�
y��a3D�@9��M+ � �� j��:h�L��5D��[r䗸�B풐k�#��܃�9D�$	�߀J� �˲���m&��� �1D�xB�J�O�&1��.e�^�N;D������LN�4�t�_R�6<�to#D��pS�.;�Z3A�݁ �3�%D����Y Jp��������ٖ�/D�X���نf(��#�b��WQک3S/!D��C-�#�,�,�� 4�y�t�?D�$��EB'��O��L$�a!!>D�����
~:5
�K�+b$��>D�(�eH�S�@�RfW&dNUJ<D����i�d��0HW�k#����;D�L�F��n��D��&Ipq��$9D�H*�`]�Z�*5�!�P�y�"<��+D�\��$Ъe����,Ϟx�H;�C*D�D�D�ԕ%�Q��̇'+�	P4�&D��i�2k�\��d�@*.��&D�� Zi(dk�`�J#s�L�4$�u�b"O����-P�R[��E�(��]��"OJ���-�<k?�d�4b�/Z�J�w"O� ��˽om�a2"�g�^X��"Ol��+��~�4D��A�(;yNٱ "Oؔ���k$��9u'x�C�"O�X:�D�&2K���(3w�Y"OD��5A%q��[ve �>I�9� "O"�Yt9h'���P��XDQ�d"O� p�Q1H�-(�fف3���"O$��c�O�=N!�% 0d!�0"O<UB�d�!/D`�dV�<�`U!�"O��)�&�R;� ���z�p92s"O�EKG"3R�q U�P�m<��"O���1@�t��yX�NcsU��"O� (ճ�:�e����9�ŝ�}�!�(r8�D�J���)����!�ě:i905�0��z����+S�[�!��ЛDEa��+@Xaǃ;]�!򤓮p��*v0�pHt�!��;-Ĭ�s A�5�������F�!�d�6�"PACq���+�BF��!�d�87/F�ԁۚ9���h���D�!���7Q��r&��襙��\d1!�D�`��+b�S�z�h$f��u%!��0Z����XOtvx�#f�@!�� d$�	�K�	�.�9f�BS�!�đ'A_֡�QE�1Ѐ�r�)�!�DC�8�C�@="�ԅ��)ҙ-�!򤖱 �-���L9���@���U�!�D��+y��[6��(A��q�α�!�Dڻ`<4�Rb@ ]�p�p���!�!򤆃)�~I)a�C2}���M]�6�!򄉎Q|�Z��QcX��C�mW�_�!���q�L��1i\�O�vPI,BD�!�D�HW�U*q%��Q�p��� !�&j���, �(��B��@�Yr!��_�m���yg �r<I�g Y=3X!�$#M*Dp�!Mɒ
rn)�o'I!�D�A��<Q�a� ��X�0O�.r!�D�/fD0(R
������+<.!�d.oP���Ab,u{$|pQ8g�!���3�:��aM�i]����s�!�Y&t#�t�G��r�c�c�f�!�DE.8��M9� X���ث��/:�!�DӞ"3�}˴���+����q��?�!�E.��Q��ǖyh����3Z�!�d^�����Nv�d܂a��71�!��&Z��w��lJJ�"�Z$�!���Z״l����%,�U��̸y�!���3c4��%jS�Y��#D��+�!�ĕGH�鹐��$i�&�s��93�!��^tw\�3�G&s4��/ù0�!�d	x|���Օb�B��B�!�$�	ZP�5�J�:�/P�u{!�D��Kal���A�)�e˚i�!��*�ƹJ�e� :*(��	�f�qOI� I#P�T 7�]��. �S�|2n�$�;��\}�)��Ƅ�yR�/tp1��.�"eҰ�p����yB��<=�a��
�"��
��\'�yR�LD �1�O�6Ta$,��\��y2�	3f��I��fp	�����y��;5�~��/��
�ڡ@�W��yr�.hȉQQ��R�n]��nAs�<� �hE�I�B��Xè�M�h�v"O��z'���rq�)���x��"O�P+�2 ⰸ�hЋ)�\��"O( ��ǟ�WI��U��`2B�I�"O�M�妋�T�Ri��m;�M�"OR|{e���9�b,���x��"O
2� ӂE�<0��6:z�8��"OJ-sp,���so�'!����"O��j����xR,<Hc|鉰"O���%�1�V����J ZHxM8�"O�Ԫgl��Ό��a;���`"OL�A�ۘ8� y񠜌��4�S"O����"�N�ĉ���*?��ٴ"O��:��x����h��$pӆ"O�T{!N�^�2�*V9���"O�Z���=a�ēa�Ϋgנ��P"O� �צѢs�x�C��dg�h�"O4]�2���/,���0� 1c����"O~�x0 ��y�$X�|�i�"O
 mʳdHLT��$�x�;"O>\B��K��<�d�֨d#�ԋB"O���GI�%o������_+p3�"O�I�&�u\�ِQ(:��3d"OV� X�a�'$H��Fw�<Q��{�x�I���P�;7h�O�<�I�F	�г睑T�j��0�B�<��N�p�L�c�ḫJ�U��Nf�<���߸S���Z�m�!(����u�}�<a��,2/�x91���t�~�umy�<����<G.x)k��OKz�M�H�y�<QS�I�Z�$1u)�{�� "�D�t�<�e�0?�Y1EL��!��,N�<	(#"U�5�h��h�R6�H�<)�聎7Pҝ&ċ�Y\�1���D�<�#nU#KU&]�cK�5�T�SI�{�<q��ӓ5����N�! �@�Nm�<�F��
p���B�V�&�R�<A�͇�qv���N_#?�����m�<���^)q;v��톉p�Ґp"��T�<ѷ��8�"t�0d�^�����*
h�<�
\`8T2Fh�5-h����n�<�G�!x�<M"a�D5r&%`�MXg�<) �Bww�Xx��X�`Ne9�Yd�<�A$/���ZBK�G�HQ��`�<��l�/dDP��)a���Cq�<Y�сID�`k��H�L`.�"�JM�<IW��b؜��Uc���3���A�<y�l�v0<lA�-`�؀�-b�<!�01��ਖ�(]f�����R�<I@DΞA���x�)Ƞ3���Z�G�Y�<Q6�j7����MƸ'���2�
W�<���/�\�"�̹ ���oHG�<Q�(�!l\��R�G��|�cv��E�<��K���Mj��ۄe ����C�<�E!(Jd�+A�E	�z���d�D�<ĂA<Τ��� *��D�r�v�<���7ÞY����g�Y�2�W�<Y�l!�T�Sn�iP��E�l�<��	T�9�T�+?(��IV��d�<)dI3c��Q�r%��@�V��@�J�<�q㟣YlRȻ�l��^�$4���Q|�<q7kаr�t�
�$_h����z�<��	�a�j�À�O��d��x�<�e̤W�
�(��U.�:$i�i�P�<� ���e��5��\��Ũ�"OF([�d��z'fȐ$�|�u�un?D�\�"�L�
i��z���3�x��c"D�02�G-6��|	���{�����.D�(*�`�N$Q��i�DL
��� D���	6]'D��`ՏH��x�b D�D�"`�~�r��W,C�����G/D��YF�S}& ��'"T�N x�7D�L䋉?m`赀᎓�R��=(6D����P�	E��m�V� D��6e�w����W��-5���5/)D�P8u�P�~D4��k�m��3��"D��`֌K$/���'�Ү/�`uB/D�dЗ�΂¢-f�����q�.D��X��[��tU�BPJ~`��-D�(3�kۀ_����U/#��E"+D�x�͔m:��E�P�4�z����7D�D��ȑ55�d�t㒣g|Dp���!D�����*b��Pd�7^�ań.D��ʵDU(��0��D�+�@B�-D����J1U�@q�e��k�`-��&D���D��� (|�ミ�?>)�p�#D��h�ᑓ.�D=��F�Iz-"D�<�e�^�)*ZP��L�j�X-2ӈ!D��(Ɣ�+@�l�Ҧ �dB(I�� D�D0D�I�)B���%�X�5R��F,T�<PK�=B9����0�"O&�+6!W?`�eB`��
)�4��"O�8{��4D2K�D�,��"O�9�"�I�#ަyi�5R-N)��"O�CFj�8,�P��w���$"O�)xBGK�h�\��eU>�]Q"O^	y��;��I�@d#\�!`"O�8�b�/# ����
1A}d�aD"Of91��ĺ?j<�C狚NS���"O���ק+I�r�X7�V�*E��X�"O�`�C��	w�xu�H���̨b�"OR ��:��%�I7+�T��f"OJ]�VCӴ}��I�Rm�/%��p"Oi���_f���jB�2��t	�"Or�A��C��M#e�Y�~�n�B"O�����T�J�iF�u���"O6�j�o���� �(�"O��8)E�z6$X�b̖?l%97"O
�8� ͯI��bL ,X�W"O��j�[�y�T�e��O���sd"O���1�e8fD/9H|a:�Gй�y�O��_� �˥��,5(H���;�yr��2T��рS�]�$�� J���y�G�4Rp�'FR�-��j0��%�yR�:
.$PS�Ҳzي����T��yr��!v��
�)��;��`��O	�y�ꏑDݲ|c�"�=.�xQ�aF�yr��l:wF�%��부��y��E�O�X��(��"ՠ�H�)ۏ�yrI�.zp�!o^/=$�ۑ A��y�&��!2�ᙰr�V�dL��y2k�.��y�фZ�4�X=�FAP��yҩ�P��1`�+P�2��5`Vℬ�y��9���@��1��i�Gϼ�y�\Q:V@k�o���J'�y��2#�b�5�T�q�l��y�I�!vְ�����[=h�yҧF�y�ꘄ[5d��S���Z�!�դ��y
� ҍ+���6Q�	̦x�JR"O�<3Ũ�� �#	�}�T��"OJŻ�L�L�9�1���v�:pI0*O2�J@��{��%:�F@6gC�1�
�'�~ܣ�/]�
����&N@j&(S�'�֤�áԖ�Jt�f����'1�H3�K
��E�Addjy�'V� ��^�L���jW�����'%Hp"��(>�A�C\'��
�'CҍZ�'
�e1/T��2�[�'.hÕ��<�� cE���l���' ���4A-W� Ke��'����'�j<�DiY�k.2��'IV�!̈́	s�'"H��!o�W8��#˃1��-��'	�<�6��}��� 5b Y+p0�
�'*,ۧMԎI���A���D��z
�'e������1"��y��e�(B�v��'�,��� ��f��3*�1v��T��'r*�j\�pa��ڃ�_�_ż��
�'�4�C� �%s���FQ�f=�
�'��8 lвH������@2�Hl!�'�bz#��v11@�[���l�	�'���Q��Z��NP�Sb�H,#	�'c����kX&k�2��S%]��XE�	�'׼��P�F�Qd�#+�(k�
�'qt)R��:'r
QP�����
�'�M�T��|F,�C��ݒv���'�n�aK��_�B�S�C�"�jE��'��M�c)��E� �B3#0[w���'_v�г�Q�9ͲȪ���T# =��'�>-Sq	��e����W%VHnl)�'��$��*�$[�r�FV<F�.��''��뒫�g���	�j�"�'.tCUG�"�XXK���;`�p(��'_`�)�iڣX�~t ��)��e��'����	C�'��i�T�� ��5;�'�`�c��ƯV)�i��@8>_lq�	�'��+s$!�� +��ѥ#�怸�'�n�+�3:��� 6UM�I��'8����x�\����G�qq�'S�����6s�T�V�DƱ�
�'6���&��0�����f�R���'�´���P�ڨ @�0�İ�'y�ɰ�jˬ]L�@�L�gD�1
�'�Lٻ(�4LY�� �ȅ�7��L��'V���k����=1��Tp0`�'�lD� �[D�da��J� <؈P�'=F�x�N3^#B��F�J��Z�'���Q��
@9�@�Ŧ�%<G�P�'YJ\�J��g��Q��Y�2; \��'� 433��2�1��3�z���'�
!3�b�2h3<iסA�/9�<��'U|@҇���&��3�N�3#H��S
�'��̉b\L9���r�`T��'�4@�ݒL9��3���`h����'�hY32C��N!U���ށj� X1�'���˴L4��Gm�N�9�'bF����M?A�h(���u�!S�'�$�qe��#�h!y�D
�Ws5��'"L����"F�fq�e��RC�%�
�'ԐM(�j	�N��,��ؓaJBi�{R�� �4��hJ)u�u{�`�=��="Nik�mZ,���(fi8 �ȓ�̡�HM�I�0@�.��9B�̄��Z�8v���ܕ�Sl�#>^���S�? z=R2E�!"��i ÃL�tq�'"OB��Dƒ,��aQ�i;D�FIP"O�MiT�G�\�2H�,o�,Y�"OĈ��M	�?�P��t��t���!"O�=!ы'YU�Tt#<��J7"OЌ� `W:O�\���F)Vx�s7"O��c�@ؐ
���j:��W"Ov�A��9�LX�a�/���R"O��	��J ��J 7�R�"O�S��D�2y�̓�&M�8�B#"O�X�A�+�0m�ǄR�)lr�u"O0�I��4g��9�4�W	=c􀐆"O*���˭3I�����U���5"O�P(\�w��X"��>@lu�D"Ox�2jC����sǋXk����"O"�p��[�o��l���,l̹�"O�	���.I����X4i��-��"O\p�w/�tŔ#�M�^��D"OfQHQ.2%�I��!
B�P�R�"O~�J��׮!�l=BS�P!6-V�2"O�Ű��1VL�c�O�Z|ۄ"O�!@�V|�ƭk4GVa PB�"OJ����=2�mҗ@ RfαA6"O�P�t�HO@�$cB�/Iq|�4"O��`q�D4\�U#�O�4Ml*4	�"O0IC%���.���2���+
i�,�"O���W!EL��S�Ě&v`���"O���o��f����eF�g��Z�'�X=�QER���P���$V����'c~qZ����d�Q��Yj�I3�'ܴTC��؁�`�b��?V�Ys�'` /�2V2��b�g�0h}�'{��{E��� p���S+�F� �'A
#	�� �&�V�4���Z�'J��ũY֠�lya܌��'�f kqሗx��
Ն@	h@��')��@L��+�-�/�	�b�z�'�\���.M�le �!$?#F���'�B�Ӣ�'BL<j�삃}pp��
�'"Xf+G
ļ�xBL�>|�pU2	�'C6�qG�]�%ON�Iː
� q�'��p�䛶�hd:�KL�u��H��'q>�h�BS��:GK�}d
]R�'�p�a`E53�x�P��0aX�`�'��	�6*F�4��Y�g@W1	���'i�D���:n�x��F�!ѐ��ʓ��$-�9u�]��L6c^f!��IB�cD
��0}<�B�%C9�(��)��c¦�#-��:h�}h�\'�\E{���A޴[�%�TA�4t��C�N��y�M�aX؆(�>�h��%bS��y��Ϣ2�����/������!�y�1�#�Fͻc���a�ħ�y�� (p7��@s�GS�U2A�[9�y��,t(h����=TI��	��yBG� {g
�8%`�;[���	����yB��j�<!:�.iY�)!W!��yr�ԏ)��x3n�UG"}����y	^�)퀠R�١ AHɋ�G��y�)M |���!�� �6���,��y���4��<V�Ý��r@�ɵ�y�"�22�l
S�E\ ��
�=�y₾?uR����W9G��3 ��y��K%5D`�"\*��8ѐ�(�y
� ��#��Уm帍j���%�)�"OFi�FD��Ӆ�p:)��"OT]x�C={�J�c��Q�Q��d)�"O$���m�=3��|c�ջ+�"�pr"O<xe'��69{0"�lth�Z�"O�p[r�~�ڤxw�:p�I "O��� �9��Q��P$%&�4�"O��3a(C�z+~�����: ��Ԁ�"OySFǯ%_��+P��%��uhc"O��b�	�,����(]���`3"On�� J�W��y SO:W� �b"OP���O�����f9�:�K�"Oڭ���6������*��8'"O�Tn��L��3Dh�@��"OT|
5E��$&�-���3aJ؂�"O��r����j�N�Ӏ"]�LP��*�"O���6��L8�`��<(1��SQ"O�M���K�q=tLGA	U��pP"O�eN��@��98�R�P2�җ"O&;s'�6��1�� w���Q"O����S��T¬�K��&<�p��rtƭJ�jU.H�(˔/H�Ub��ȓ>���c�6ǺS�.ʶ*"��,�0l�EOƿ�|)+
�X��y��7BN��k�S�P� o��)�*��ȓ6��Ax�
��]���b��8�h�ȓ
|e�0ʌ��bu����3E�\�ȓ=�9�d���X�n]r��30�<����I
�j[6+��*���2LD�q��kŸ5��WIZ�񢏘"Nzt��2k(��c��	��x�rA�$�b�ȓ~����Qo�++x�ra�[35������d��CD9�����0q�V���h���L�'A�������I%4!��h�J	D�O� x����+VΕ�ȓY�ִaF�(Lr�5*O�"!�T�ȓ�)���F�t�1b��=~���ȓ��0!ը$Cܑj�m 3E��%��TNx����+Va���
Nv�E�ȓ;{����J�RV����ǈh�x}���LA*��T
AZqS.�,s�H�ȓ=a�a���m~�����9���WR�)3B+,z�9��o�#8�¼�ȓIn\���"kCH�UB�T���ȓs��,��}��`��Tف!4D����%w�x0X�OC�&> ܓ�2D��D�3���f
�g_��)=D�p���߱@��e�'�Ӑk6�B��6D��b��:m=��1e�B�ݳtO D�H3�]�����`�~��"�>D����O=��s $щp�h9s�8D�J�����X��L3#�\j�3D�\���_�v2��pt�B�Z�+�2D��a�B>[6�&FMj� l!<D�dAq�?5:�6��=w���2z�<y�lU t���t�^gȲ��'�`�<��o�@���Mґ	
$�cwH�^�<!�e�D&����S�$M
1:���]�<� ~�%��C� 	Fd�p,�q�<�(��2=�`刑��(�j�<��M#?iXp�GL�4j������i�<Ѡ΋�+����!�h8؁h�M�b�<�sʗ�8º��p���.`����a�<��e������˻	Ԭհ�N�Y�<� ��Q�r_X��cM�{F�ͺ!"O�9RJ�$"�а�'F>e��"O��A��2JB6y�4k�6�8�@�"OT�C=7|n��1�,�X�j�"O���$�-�d2bh��y��u��"O}�'�˯9� �����,h"O��[&/ҁ=c�I ���D���"O�5��A�>�E���۩	�(p��"Oȁ1"�$!XV�H@+F�0�ӥ"O������a�֬ΐ>�$�Bt"OȰ0���N��dS�&
\\h$�"OʴK�eR/?� R���M�@�"Oڜ�Bd�
m9^Ȫ3e�<E���xu"O���N�Y�b�ٟj�Dȸ�"O�]i�M8{6�*W�M�i��"O�����<�Y#����D�C"O8ea�!;S40%PV�\1_����1"O��5��+k�m��a����i`"O���%���rH2s`O���]3�"O��)�\!#8�j�\G� ��&"O�9o/��!͝_��l�4"O�R��V�8�%�W�G-Hh���6"O^�)Ԥ?6J��a���I��B"O�)q��A�r(]�"��|4�=yP"ODUu�FN 9��D�A4�Z�"OZX��G��̘� ʱQ��[�"OJA@�UO�R�ЉhJl�Q�"O4��7�\�H
��8L��"Ob�����e���.�6L4��"O�hr�L�z�ʜ�_� ��V"O����	UB�����C�y�(9q"O�%����[o<-ꃠ��H*��C"OAj֫��y
�y��N�(��A�"O��'M�q�-Z�,��b���
F"O�I&���0<B��q�VLA�"O~��1؄L.��h`FPĠ�"O"��e*�-�Q�O�X:��3"O��s� N� V �r���r�"O\l��"$P�%���ڽYp��"O@2vgNuI�T2�/˕uB"�!�"O��;$���f�`Q$�F>�X�0"O��)�E�|�0�Ya�Ռn�i�"O88�O��,�y��`J8,���E"O�g�ކmpI9Y�a���� "Ob(�W�C�vJ U�j�Tu2�"OH��o6usy�aL�\�pyh�"OX<+V�"B꬘`���^v �r"O�	��d@@�^Y���$nl�$qF"O`��1�Z�d�ԩ�������"OpAsGm62�� @���_u$=�"O���B���` (��Bo�3G"O`IF�ֶK��i#�ǒ p�ȴ�s"O��Y�n�	f��*Fe���HQ��"O���T��V�4$
�2�:�ȓ|�R��dΙ%�|)� ���V��ȓPQ��@P�A4&d�Uȃ� <V����4����Y�5��+�j)5@2�ȓ<�N��$d�*���I���BX�ȓ.�`�a��׻h�\	��x�
�ȓU��y����>=�5� c�"���oX����q[�	qek�f�<�ȓSf̡Эɋ;��HpbC�'1BY��C��Lk� �18d��3��7�B�����I�aJH�e�f�J�(a���M{�<� n�C�ܧc�~�δi�~#�"O�|�vm��������|2��"OB8Z �
n� @��b�.8�]�!"O(u��1X����C�<��"O�Au���o0��mӓd(��f"O,�0���.�h��lU𠠻@"O$q��k�X��h��@�sC"AZp"O*|A�)���p@pV�8��p"O2�	@���k�X��K+;>\�V"O�����j_ ���M��.��ݑ7"O�����{fi��o��^���"O>�{4)Nr��-2�>O��"O\ɨc��V�l�A�6i�I�"O�	�ƠC*}��]�\1�fg��y���$3Ӷ�`�1S�����|���LZ��*iP�c&��V
�j�@�ȓ+ł��mG�s;ֽB��ȏ
2��ȓXX��.�&�z�ե��:U�ȓ�P�X�+�R�`��6f"�PL��jZZ$J�(_
1֬e���J�!�ȓ6�B-�Sn��a~:�7͑<~$���-:\�!U�Ɲ["BpZǭ��kT���X�Hf��gb	"�����i�ȓ{f6�	���3&�d�Ȇny�m��e�~�)�F��>0$��EK�+-��E�ȓV���#�(�X�(�IpA�,eb��"�RD��L��:���j�D�6,F|�ȓ>�]�A���$�NPv@G�Y��ȇ��,��+;6�Q�ThW� ����E�^m(�Ȓ��`P�-@�����pٜ��4�N��H� �]7"]�������Z5�RUP���	0���ȓ�iJ�HH.gv��-�(�d���(ř׉��#���!�H�XB�ȓ(��d�'JŪ �B�K��*ir!�ȓ*�����6�����˔���^/����	�<j;���CG|�ȓ&<F���Os����T�
ܒ�=D��1晏AΜ�䤃>V��嚁b=D�tY�I� ��ZcD�^v`�$�;D����KD�t�`�x�Pq#�;D�xx�lǉ2��5�Z�8,�c
��0�!�	�q%���Ŕ`پ}a��S
f�!�D�cr�+�$�n��(����.!��@u��	v��9��$(Wi�X*!��I&W�h1���H�%���fe��H=!��5�"��a�
�5���2'G!��;>����@�7����k^�j�!�d� 肠��[�.�R��?g�!�$62l,H%��e�����S	z�!��3��9B*��4.��e
�!���3� 	�`%��T��K�'a�!�dA�oy @�X.Qذ�%j��u�!�d��qb��(RlI�5��<�! Ҵ~ !�d�W�T=�".��.�bas��'E�!�D�xe���U�k��c�[�gr!�$��~8`��.�0;4�a��;]!��[k�y�&�K<@:�ʆE�� >!򤂹xY�$Qw��s׺��s�[�Q)!��:��Y�4�΃ ڊ�ِ�	1�!�'f���\�,�� Ǯ�7U�!�E��4u[C	�2j�颭�k�!�dId�!K��'
!�H���9C�!�$A��yq-�F���$��9�!�� ��䒷uz��1���.6T�P�"O�<�""�%E+@����W�j`S�"O�(ۡOTOB<Y@�������"OI �UH\ڡq$H��F�b��A"OtYCǯI�Ș�N�"%�����"O���B�#L�T�1�m
�Qvz�p	�'�<xqu�N>{؈z��	�\V�ű�'2�D9e�ܚ$\޸��lĊR�����'�\t9҇ߞt`"��gd<��Hi�'��
���<c��rD�3ǖ��'�����G0��s,[2(��'�l3��� k$��qJ���(	�'��)R`دt��az4'�X�(�'� �u+�9�&A"�A��R��u��'پ�z����E]����C�Lu�<��'�t��e��(KT ���Epf ��'!,�k���e�-r��ӡ܀��
�'V����"_�� ���K��u�&)D��{SKD��H���1Y-���@G&D�@�@#�%Ĭ�1��ԯF��ȓ�#D����5X������јj�z)��G&D��w�栁3�Kf$�%x��$D�<�����/z�D���\qx���j8D�t��!�6�y�Q�GLȴ��4C7D���eg����ZB膳3X����. D�`��@R�"� ��5Ѕ� D���F�ǹ.
D%��a�@�~)w:D�ܚ���o�|ya�G�+6��H�6D�|Ѵ��>�R� o�i�|u�! D�� �aS[g�Y:�k��w�B�Ps
#D��2�h�b��1���Y��h0h6D��Zl�-��ܲ��j���V�2D��C��.��y���K�f�A ե>D��CTD�">�`�[�ᝆN�&LS�.D�� �o���y@��?i��=�U�*D�H�G�ِJ���h��$m�����#D�Y0�KkO"i���#6�U��)6D����?G�a{� ��X���:eE5D�� N�$ܠɃ�4Z�<��6� D��`e���\�~$��X�Lw:��I?D�:��^�"]�ȃV��*Of� bkH�A�¡V�{N�� "O��[B�Vi��"�ϋ�N��!B�"O��	FI��6�̩�ƍ�T�> ��"O�|�N��0���Pf�Qj�B���"O8ejQ��2����@;0�Je��"O�4X��X�������8"O�ջ6�;��	��(�5�ި#�"Oܴ鵫��x9K�'U��=��"ORe	 J�Sj&���	M�>�E"O:8���ЎOC���ηH�Y*F"O
@�F��&��ġ�%� W�~y�"O�ұ�Ţ~N D3V&�R�PA�g"OX� ڍB�P�����o0f�b""OLT1`%��/�t} %.�;ui�g"O:�B�m�*}d�1�����
�1"OT�(�ĉ�"��5 �Vp��(
b"OhT��:p��l��y���cV"O,1AmF$Y��1��
Q�"O�i�Z���sC"C1m��	�A"O�yIe��+T�"S5�\�`���"O�(���c�>H�QN7P���S�"O�T��	T+V�x�lC(?J6 �"Oj��w̕4]]�5��.�,]�2"O� �@[���IQ�=��j��w�j��s"O�-�0`�&�����j
:"�ݚ�"O��$j��-�J겏�~�D�� "O�u�F��g"5y�ΐHʤH1"O�EӐ��6���c̀���d�"O,����c�N) �B��H� m�"O:{d.��JhZ��U���c��s"O�����m�~-��-ɭ��@��"O�LfN�R��MI�,��a�B�sv"Oj�ch��e�~��ѫ��N��TXq"O�]ZbY�mqI��ʩk�"O�@�w(�|�vD��m�NZ�"O�\A�U�^�V٩Ǧ�=��x�"OzݚKB_ ����S�Cy�=�""O҄r�L�4Q�8��.�5Uu`��c"Oz��CdW�|�ɐV-';p���"O)�f	�&rs0p��j[+d^���t"OdIsdF4c��HS�iH��B]��"O���d�P�^f�@H �� ��"O8��1��!e�(!YT�
�H1�"O���'�W%	�d4�qk3\�ܽ��"O:���H�d�n�g+�$��
3"O�@sUb�	5����2h�M�$]S "O� �e&P\r$1䁎$}tx��U"O�-@���c��@!d���J��U"O*�� k`�*P����E0C"O�U
�.�#*�l̻��)$)k5"O恨��ݣ.n��R��r�uY�"ODE��d�
R`T��"e��^���9"O�8�0M@+�b}�W����H��"O0���F��`v���c�
�|��U"O~C�W;.���V�ևozt�r�"O
�穜�C�eac��z���c"O���@��
3�h�ȵJ�;bj�#"OUz���8�������M]��"O��#�R�h�q��)�I�}p"O�y�T�L$p����c����"O^)!��\�(�r�S���ls"O�(��M^/���A�L8\����@"O��2��X5�*�RE�7.{��D"Op|	ШL��<���9Gd�(�`"O\��`��8	¸��J��@T�]�"O��c����Dż`�'�7+8�P	�'�*��wn6�����n B���9�'��A��r�49yD-."I:�0�',`�Û�fmr�RT߬h00�'L���fƔ('t����B�����'bB�_U�q�o7����'���h^�i�T*c@��gd}��'���叇�7Dd� ���$Z����'�bxǯ ��BEP0�/c�^���'�X��߁f�|qh"BR�]� ���', ��ժ:R)���A��d��)+	�'�J��B+��ҰZ�(	�'�e!$h��;@��A���X�"E:�'B���7�Z����!!�bzxxx�'?�A_�@wN��p�ڡ[�8�2�'�|���k�^�@a'l��V���
�'�L�1f(��U��8����5���
�'�L��`Y?I�X����}�p�'V�t
v���m�e�V�D����'�j�BEE�<�e@՚>���[�'m�,�U�ڵl{���� �8E��9��'n6�:q��U���IdI+A�Z\B
���  �Ї���Z���A��!y,��G"O���E�.��s�H��_��"O,�j��h��h�!�H�!$ё0"O �#EK�AJ`m�0A��"O���ː>���#eKT�B���)��Iٟ��w��"u�F��G�T�.̓�N�}��4��ޱ{MqO����S�u�T�ӹ?8�iB�c��h�\a�O���#쏙E6�I"d07`��Dz� 
8T�t�E��9-�½{Ǌ��L�\B�ȃx�P���L.q�.l�c�Ӿz�B�����>�r�'>�7��O��'F~ҀjDMJ;�@���R�)3��c�'��O�h�?�@Q�� �gc���r�O<�O�n���M��4{F>���$TP�G!I�{Ԉ��C�X� �i�U��ē=��40��[�6ܩiUg�'h�d��3E�gdtUhDЇgu������(��}���ߝ�rCD0��
<< E�e`|��@q�`Z�
֖����	;r�4"��� @`����8���D9�MS��i��eH�1��iZ¡����?�Ƽi���s�8��O�#�I(�$@�l_Fm[��O2�Ġ<��\O���Ę�D���X��T�T�FzR�i��7�)�������3LV`���ڧ�2�х�e>B=�(Olu⣤��剺A�fI;1�Ƣw��!��"b'l��'.f�C�̐�x��C��:�2�+����x0ϗ�1��$�!�A�*&r *�j�6�إk���$!>�a@�z���Ptw�i���>����q�@%�́~%,�,Q�|�R�*u�I��M��	z}2��.h���#�E�j�7��F�˓�?����?���'2��X�@�-\��a� �<<1֥!�ϦI��4���|��'��t��XPM�f�ځ#���Z���"<E����OX��D
e�(�+3�i��jǖL���b&�4�(�P �T�oߤи���]��!�t.G�>�x�7�B4u��Y:�&5���� C�IZ��J�/�nf�À�7�	�w��f�L�2���Pn"��΍4�����D��ē�?!������5A����7$�|H�lлF���>q&�L�e�
�s���<�C�"�j?���i�b7m�<�p,�=r�v�'̉O�4!��ꄲO�9�!�W'T���8�{��'�� ��M�aP��8X&�l���GY��\��X�L90:|]�P��8#=�4�&yB�u�X�)�fH��� �i��`�f��p�ܙ2Q�+����Af�W�te �ª���?��@)���'=�S����0��б,�0m�lR��Z�?��Oh�� � �ׯ-9�٫�"D�W�b�Ui9�O�pn���M��4��+c��"�|� ��ƌX�pFB	� Ї�?Q*O�IW���,O0��׏�=*U�����nA�`��ïV��Qǂ�U�o��Mcs-�dܧ���]j�ա�,���CȗZz(7�7D��\#�fH�
0 ���d>h��4\���k��4o�������l��!#f"��������?A��i&{R��a��M�p쒂k��x[qE�0M�0@goM^?-�M�+O���Đ�u��HR��S�h���4d���o��M�L>i�j>���cK87�D�j��'x����O����=� "�    �m{EHY�B�F��OA��R
r�Z������^����H�9��$�����[?˓�?��O>�&_�3�� 8DH�:2X2k�O��=E�t��F�n�X�兌9�d �䔏z�� o�!�MkI>�+���O�6��  �  �D�)�D��'RY	�@J�W�>�Y�&M�%yb1��'d�W�=b��*�>�p�)��4D�,���L�Kh��(s	�%J:�� 2D��#'*˲P�
���ψ�D`ԙk$M0D�pҵ�H�F�d�7��gsNu�C�+D��EkT�2�(:�-�(�$�-D�<�G%��1�{Ў�0dP��閎+D�0)C$�]ݴ1H��@�?��df�"D��	�),ra,=
�j�qܨ�n#D�Hا�O�t�hQ��%_(��i��� D� �斚"duzM�8��0{��-D�0����q�4�pe�)|�f��I!�Z?*$\����N�0�%��?#!���y�F��eL�x 0xJ3Ƒ��Py�c�{V4��3�ӻ�Ą��Z��y�@K����@�-X�e�(�6�ybD�as8�0� Ӧ)�l�X5�P��y2�G*:���b�])�PȚ�o
�y�E�)�T)Q�V",�H�����y�mA�`tr�JA6#3f�3����y�G��]xQ�Wò��K��y�i�'.p�)�`زR\��Ӣh�=�y
� �)Ag� 56��V��4#\Q"O��D$J/	|������W$�""O�%��8)<�DB��X�{�"O��a*�e�DD���Y�!�d"Ot3�$U!k\A�`�#�6U�"O�-����?&I��O��s�-C�"O2$��"�����c��DN\��W"O���b��|_����_� t�ȓgb�؂B��-OX�۶����<���0� >6z�A���&of8�ȓ(�j����ٞ�iJ�L􆰅ȓF.�81�A7&NL�y���#�^0�ȓFW\�3
� )�'įt�"8�ȓ(�[�f«s�Is�Ì?|6����FYh��_,�r{WKБ?�ȓF��`�Fe Sd2��ҫӥ��1�ȓ7LL�%�j@:V�]fu�!�ȓ)�4j��ɕP��!f�S�oE��Fo�(;�JD8�]IëG:RBe�ȓm�"�����5�ƕ��MQ�r����ȓ98��"L�+qV���.���^=��q�\i���N����V"�؅ȓp�-3���E�Ryu`�\�D�ȓ{��r��5-�a� �l��݇ȓV	�-#�V�WJ:��Ca�x/���"ޖ�����R�z�+4e
�x'px�ȓkZ����&Q/��'CQ�x�`!��iBuaS��U�&y;��"o%TԆ�=΄�(Z�3$+���5I�`��Gd��ؒ%��e���1r�j���fW�3�k�);��� y�������.H��IA��ʇ :�ȓN$r��# )P�^��w�Q}Nĝ�ȓs��Œ�B�*����L'vu�ȓe�t#����$	��gB�s�Z��ȓ�=j�CX F�}�w��e(`܄ȓ!�$��&�D�X?̩@�X5��E��27&��Mq��I�BP2uB8�ȓE�rL�W�S�r�B�J�6�"u�ȓv�$��D�
�Nz�N�<����h�%�\�h1u ��Z�L��ȓb����փXG��P-F�����>�X2�ʔ�����䔍� ��y��UZv-,l�ܴ u�� n�C�	?v`X��"
J�"@��G�sg�O� sT�̥��F;�d�Q�P���OP'lE�"O�4{6�'��Js�G�%����2egt%%����<!��8m�>��GI�?����T�<�@�L?�AJ@������ِ�p��c�%V���dݟLK�ᗅ}h�� Ώ�$�az�KB?>�h@���R?��K� m����M�<��a��n�<�K�Ex8�,|��d�7j����<�W�5l�����D+�'j�|� ��!o�����J(X�0T�ȓ*9���1��%ej��5�S����b�,&��'�:�я𙟘AUf�S0��BaY' d�1�)D��J�
͍B�, �+��c�b	�V�+���8��	�r��|�*��+G�0g��3����i��0=� %��x�t ��J3hS%��0
a��'ՒXAD>D�,�$�@_`<D�Qb(g�����?�I(f����I�#I�Q?}@���6\��1�G��Dt$xqf:D��b ���FS
��U�N�D�;�aث��bL>1��8�gy�/�1W�@�ғ�R�J���)����y"!	�����R�ިL~�I�$�-�M�`=XXH��ןx������E�4 �ʞ+r�!�� BpZ�a�7i�� 7f@��ֈY�"O,T:%���rmtLpP�[�$?�AJ�"O���0`O�D���Ä�,,�(4Y�"O�� ���tX��3��tĶ�k�"O�ty�
ǬW��pSa�r���T"Ov0�w�O/�bAQ$���x����"Od<p�X<���� ?fRH�t"O���[N�f��Q�U� N����"O���Zcu���Q�Z:?RP�Q"O"Ē&��MX�yf��jLx#P"O@�{7H��{�.T�0�GP&�-�"O�4*R-�z���g��
Dp	3"O&<��G.I���5Fo<���"O��Ql݌o�V\�AŖ�@��"O��,X��^��*� $̄�"O��"�9w; |QwjB�= �Qq"O����$ص6�v�q��F�mpt"O<����%bb��iG��	qF"O> Q�	JBѴ����C1\
�!rt"O�-(RLG�_ЦEa�CMQ�j�C�"O�!�f��	A���h&z�X 7"O�\�A���k���Hvr���k�<���%M�	�kI�Y��I�Wy�<	�M�3~�0c�=����v�<)�*�5q+Z!��B���@\H�<a�� :��s%�	n�P�[��RE�<9�W�m�B�z#�� %�t$Ii�<	V@��*�G�vo��K���d�<��e�1k��+�ǂ[�`�9�x?A��ؙ>�'�����Ӳ�5���'|���O�P%�i1����n�1�����w�l�AED,c���`s茝
��gdB�8J>4j��*6��̉P�ϱzC, ����O\�BS�,��>Q�Z�y�ؘ�ڸCp���G�
k��W��MY� �4B��	WH�4�O؎%8e`�/h�D�(���\�NM����Q ��V�T
`����IT�0<y�CE�<D S�T3Q� �ŅڝE.����4ZS��ԥ�.�Z��[ e��@�shA�5��x��aK�R$}�`��f4�aR���x�"�H>�f����@�f���?�����i���h0+Oi��DX@�J1�����p��O����ޠn48�j�i���E�ɭ��=�f�_��G�h^���5f"Yb �a1�
P �
���Yi�5���Y&��@@*sT�����,O8���σ�&w
1`"���Y3�$��=a�A2QGA�<
2n ��#lڴp'#�s�1�u�\�d�!�F�	q>�U�ag��^{��56O��
��b���q��4E�ջV�S��8����m��OJ�O1F)���I�~���j�x�4Hr�z9|�i�'ȵD2��7��A<i�C��c��@� ��4,���V�
�N$���K�3P¸�[� b��l۰���(3UlK�|zVe܋%�
L��D0��������a����SŜ
q]p�Gfi���ED��6,�����:rfd9�����YFF���/s_r�?�=K�l���14��u ԁ1H���?1����Yv� �M�bj<c?A�C��'�T��%3[R9��OZua���_�R8�u`��<At���8L"�P:*:�GʘFъ�ۃ��!p"��h��dV��[DW�!��e�� !��Q�Э�E.��tw����0]��A�;^���y''�A؞����C-0�����K�FI�f"�OU�gꂑ7���X�.ĈCg�����Ȩ�`׼/�!���z��Ğ?T&`9�K52�������?K��j��$ҧ�0�`RC=P@���R蔙itvфȓ	��q����#BA��@lڞ1'a����u�)���q��G#Tq����/MvKq  D�4 $%M5:�r� �#�y�4س㣟����$���'m���slI�4�&x��O.j ���@��!�_�2���`
U A)� �� �@˗1D�D��o��. B�pP�]3X
$��o/�A��l��+-%F#|�Rʗ�2��AS󈇷����A/S�<qB��عٴ�\�9~�qÓJ 'v�%��i��H���O?�$VV�őf�K�����l!��G�-�ΐQ�NJ�)�0w�:	���̫tX�| e���0=� p(#oT!نyx��>d�Εz��'��]z��<����臰e�f�ks�J�3�~�	�.Hc�<�ÂO7T����((zP% ���Z�'mڹ��b�6W���E�dj�
P��C#F�"��#G��-�yb��_"X��.^�&k��¦h��M����i2���K>E�ܴl�zh&Տq��p ]�<���ȓv��jB�$~vBE0�S�ZL�@�'���5� S؞@P � �z��򤝗K�A�e4D��ٰ��9�6 �o["f蚕��5D��1[e��C�G3?�@m��0D�X�-J'�>,+Vl�6�*%Z�*2D�$�� @��W��Fa1iԇ6ړZKj8� @Ю���CC��<rw��3g�ۜb�: �"O���"	ئ2� �sv ]=B�|A��	,��yc��:e�듟h���K�B���v G�����^*�!��3�uٱ��4�,5Bѥo�v�A?,>����F[$EN�9��J�f$�s��	:��\"�D�4�х�	�/�(iE���F~<1��l˭{���G��'u(���B�iz�Ԇ�T1@%� @[o:�Y�f�Hl��=Is�Q�<ވ����TlÉ�T���)�L�ٱ�.e�&�� N��yB��!u��q!Cͽ�DPP"Ɣ%2-2ǌܔ=��Ca�OfXa��Y�|q�F�7�zq!eF,uM����3D�@Y$�8M�h�7gſMA����l�D72i�#D$|N̻�d��<���	!�F �'��V�L�2�X_������2H��bv�c!�e!���s6p5I0H�i�D���F�V���h.��f���@�G�H`f��R�B<pׄ1�r�B=sߐ��f	�Sv<�$F6��;]��a�j�z�s���i�b�>��n�+�������P�e���1� ��H���UOR����X&je$��o�<�ċ&�gy�G�Q'��D�Byz�z ���yb� L�`����j��S�z���2��4����a�0Ÿ�HN�,�`y�KQ

4���(m�v���B˿pz��[i�X �	�}�䬱S�3��'���	���C`n	�t��� �L
7$^x�Y��)Hnx��	�&0(�S4�{�6�)�@��fPF�x�.��M��xҠ����Jݖz�2#~R�)I�(M�\��dM 1<v��Dx�'(>9��Eȝ.��}.u��AK�Ά(P
�|��F3|�εIcΞ5&�n�'�.�G�,O�)��\T#B�W	Ѣ.���Q�3O��y���w�9�J�"~�Bf�ekֽ�PȀ)/�B�g
ʦ�!�̍;��I2�49Ó�)a�M�6b�,}l>�R�><�V-�<Z��b�8�vmE<[��	�~��qy��5���[ �«9G����U�"0L_�y�PIj�Ň	"�):�h�1E�YI`J�d(<A�kP=Q�uaS�E:@.<�#1b�|�'�U�C�]7��^��@	�80�F�iRÊ*rF��f"Oz�� � ��hؗ��*B]�1�uZ� �C�EqO�>��$ƛ ����X{v��d3D�,��
'bT:���Xl�R�Y�3D���ë�S�61Y�g�+@�8�0D�� R�w\f���ۗ�D\{V�,D�4a O�31r����-b�^9�g9D�h�ӅK,o�R��^�Zx�B`8D�Dr4,�%60�_�3-7�*D�l:W�;;4��i��\�u������5D���$�Uv���.I>
��)1D�T"���*7��h�I�vؑ��.D������$#B
�p���;��¥� D��Y݃Kzn�@IјF��}#v-*D�P�f��4��A�w�O�l��1���6D�RX�SN`��`��2�#2D�dq�a���AR�I�2��H��0D�PЅ�E�:8pC�$=�i�( D��֧Z�1MdPɐ�5\�|P��d?D������ʽQ�ĕ_�FH;
;D���I^!w���b��QV�9 �;D�H�'�Ð6��q+Y�z� �"7D�$�犼l~iq�V�nr(��"'D�� �j��çLZ:�DjUm�\�d"OH���M�@DIEV��$��"O��"b�l�X#�h
�gk`�Ґ"Olh+F���;����C�Ms�@1�"O��(�
�[�ex�/K�ph���"OdI����	Yg���qH�c��዁"O�M�e�O;`�Vm���19�8S�"O�\ڃ�G� ��Q�f*�w/��i"O��TM�:=��"�	L�2j�cW"O^�҅���J3��đQ��P�1"Oj0c7�[l�X�0�Ȝ?{"�Ъp"Odq�ԧs�8x�&K�\	�H�u"O\S�/P�7m4LACE�*��]b"O�8���5k�(�
ㄝ!@���"O�y��N�W��$��T�uB���"O�����S�����nJ37
,M�'"O��`t+��uܴ#vmn�vh��"O���g# �x�4tѷG�%N�V�S�"O�Bǀ|G����GQ/XrVݸ�"O���	�F�����C�'tB=��"O �s	R/0p1�Vi��ykK�1:�>�z��A��n����w�)���+���e��]��R&^� ��8,��\�΂H�)ڧ��Md&ӫK6����38�po�Ag0�ҡ�|��i٥U��5s�D�$_�@���,$��YR��s≫YI<�����<�íW3�����fy�Z�%�4��ˍ��xםK�>��Qx�F�rW���NWjy�L�4�Y�+\�ݨ��7m�?+�1f.	m��y�G����c砕�FAN�rק���DW�͸N��J�*�6�>Y�r�q$ވC��)t� l[览��^w�t��tdĦ@�pٓ䃞Z�<�Cdj��IFDhT(׽I?���O��"}��O��x�)ݐ	��8��U�P?��T�G��	��/[/\����H���O*H��e\%�P�1�١I[H�2���l_�!X�Auy��0�ɇ<g�$�S	$��P��?�,�X��	��1�`�d>��a��ʦ��"!��0|�eE'H��Ր�M�S�ʩ*◢\W�u���ͦ��a��U�@�Zç��5++�#!��7�D�j%�b ��O�9�`�y�J�F��a���iGv����;Ъ�A�ޔ/RX;tD�+K�8�k���D�I�r�O�>�ӵ[p�e��7U�Ȩ�ψ�&rJY�G�X<|[��y�a2�4��<��-�ƁړEW~���@�N)��8�M\(=Xvq���'�����K*
2��j�[�HB���'�Ԥ����.��\�RnW�A����	�'ĔY� !�@�΀HR"�:2��S�'S�J2�ܴG� �,��"�|��'Yl$������m���Z�4V���'�r0�WDӬAxD�KB[�L��'���g��&��)��$�!�.�C�'�6a懙�(t( ьB�'@ܻ�'�"8`3�6��3�n�b���h�'��ؠ�k^*v�K'�,[L\���'�d��gW	Ԓ�8��Z�Op�� �'C������P�zЙť\�EP4A��'u�m��$�#NRjp"�N�A+�D�'�����\�i����ģ=�
 "�'z�K�X	��}��#�m(��h�'[XP��l�'m^���s���aX����'*��Go�Q�3�܇Z�|���'
��	c�!u�ԭh��E���'Q�P��Ё&(ֈ�a�Mcb���'��:6o�"$F5�#�Tw��DX	�'ix`A���Ё�3@�vܢ|��'<���o�2J��Tr#�،\<$��'�t�hQ-F�$#H$�b�[:���'�x찃G��X�8�'a��
��':f��E��1�$1&e�>�rt��'��|���Ιu��ɫ5I��#����'�p���Hn\8��٥,;\x��� ��o�B�؄ 7�l>�-V"O�QQ����h��e����I=�|�"O�틀L��q�P��1��1#D}��"Ov|�EG�>�di��
p' ��"O�,q��PV��,��hE�$��"O���I%{E* &! p	���f"O>-��jV�u�́Pf�˯�Di�"OJ�p#�m*��¦%p򞉚�"O�y�S��P�x�K��1�ʉ��"O.�B�� {�AC�F:�ءRc"O!aa�2�6U��lYe�R%bu"O�p%�9�p�Kí�5��|H�"O4�h��κU]d�;�l���b�#"O�MY��K�&��u�^���ܺ1"O2	gg�,Ю]J�K�c� Ur�"O��$��< ��A���t��	�'W^�ӰJ��q��5�&��q#���'�,�3�Ё_6^��拎�8e&ٹ	�'ް��M��vb,ͰE�E;)`ب!�'�ЕZ7��M�th��(
.m �'��I�2�ͭ�y�C52x�`�	�'�~��0?3�8��&��\�Aj�'=vt+��*O�L���ߌf*֤i�'*�t a,ظa�
Pp�oZM�Y!�'��!��K�h�~P�4���>�89�'�E�g
�VY�	c���#|eD���'�v��foE#"�D�����
9:D#�'�R� E̗�y�9IѠ��f٨
�'�,��s���c��У��|�[�'�F�k1�I1f�B���"յ��${	�'���(Bۃt���j�A��e�,���'�E�dm֖���Ç�enB�`�'�`���$�	_�iu���y���4:u�)	p���o����ʂ�y�D�D�� c���{����d���y�F/Q~ e;����k���/H�yB�E i���	��I\�^E[Dɖ�y�/�}T�t*���k���Z��y`�*&$�]�d�˧�R� r�͝�yr*	�)��hC-&a<�9�����y�ŋ�nvH���/����j�"Ƃ�y��E�I ��f�*~0�3�Y2�ybKT`S�᷍S�C$�m9��7�y�	G�pp� ��2sSt��dW*�y�,���x2��e�Π�WiĀ�y2��{H�#��0�6�����'h��sk��%��!���KΨe��'�\� ᎑=2}LARc�I�Eę��'��ӱ��+yx8T"͜E�^��	�'?�E)0�05�̸��\�:����'K��8k�Y�P�_�����'�� 3F �4E��"�[W@���'_
!i!�>f���>�����'��� �Y�&��`�nP�8���S�'��'H�q���~��,8	�'�>I���a�a �ۘ}(�l��'�����L�46!�!�	��@M����'�,�!`�'^��m�&זk{�`��'�d�0c�*����6��c��s�''� �@J�**&Y�$�M<a��Mi�'��0P*��W�(�	#��#����'��}bD䥬�-vY��NV�<����K�@�"�D 
�Z�x�(�|�<10��"m�h8R��X
?���#Z|�<� H}!��"_@�� ����� "O`|���
Dm!!\��<��
�'���`���;#b=P�mʴ	<��'�������1Trf\�"(3	˖�Q
�'7"�#�j���xYd�.rXP�y�'���[��*O���^�{$���'��|3��C$_��a�ėfdT��'Ɔ,0��EP���`G4Ű���'��I�6oMg>���+�>�e!�'k��P�V�I�zt��K�
���
�'`����)Bp�)Z��xH6"O�(���f�80`�(Y�~
�"OB�hF��A����X>H�Рw"O���N$����$n�:j�X�f"Oj��$d5NiN���-M4aox�(�"O�V��~Ta��, �d��&"O����)�p��4�*v}�9"O��D��U���	$MK�_c~�+�"Od<��l��ܲ�I϶t#,�"O*��B�BU������R	�8�"O蔂��Q��h�SE��9��r@"OnM��ۖx/*XK�d��~W�0�"Oġ;7g��'�pD�tM��X I5"Ot裄'*��K��ϯ;L�S"O��1����̋���K�(`��"On��pD�H�������!?�����"O�a�"�S�D��O�A�D"O�h���(Z�}���h��s"O&%�#� yP&���Ƿ,����v"OB	q��h��`:'����0�"O@�ʀ�_
_�� �AKȩ,t�a%"O@�B%eӽdԐ<�DI��Et
��B"O�9��<�Ȥ��&�:wτi/!��N�A�<�i�CT!RN�Y��-_�!��B&[,A�t��N["���[�s�!�D�;	 �rc��Dƙ!�A�!��ԋ[����i�=f�.uX4�V�7!��<zrc��J,"A�>�!򄒭s�����k�DhE&��	t!�I�ODj�*�9fތ`{�c7W[!�Ĝ:z5���q	��+��D��lޖtE!�DZ�E��,k��خ��$�A,E �Py�L�+����'�
�Gfv���@��yr�ޚ����/W�9Q��ӕ�y���L�N��D�f��F���y�/ݱ5�j ��b��,,m3e�^�y�+�k�����*
Ai��O'�yr�$��9)� �������)���yB���v:~�r@u�I��.��y2猢5Lz��(�;U��B��\�y�л,h����G�}Ir4��K��yb�El7ȅ�����kvb�s�n��yR��g���W�H?A�%�U� �y�F\�<���nҕ	��)�,���yB��.x;�4��nT�8����sS4�y���7WN�J�F@/2	�4h�)s�!�>d�t,�Q��k�� ���.?!�d�.Z��=��h;43P�IU�
=!��A�$L	���8CD���6'��	8!���pu�}��(��gB��S���N�!�$O�.�p�x���U��!�/_��!�$(J^\,C��0ۼ|���0qO!��5Ƥ�A#K%]�t�:ը�-!�d�.}ڵG��+%����%�9A!�� �4�3�B@��]�򃁝X�-J'"O�-S��=_Ж�A�̈́�k���o0D�p�G���P�wY�m�<��Wi;D�XIQGO�U���jg`�L
va�V-D��r�ᜌL0� A!��:3�d骑m,D�pb�b�T`�رQJK3u29�,D�H��	S�(�4���!��U�hɐq�*D�PcqI��(d���|�T��Q4D��z�ɐ/;	$�Yt��#qDx�X6F0D���&���1HsC
94*p2��/D��C���M@��zr���: � �+D�����iڔ��v)Њz4�q�&O,D�4H��P�2��rGDJ�x��)D����MK>6��	�g�;r�ڑ���2D��0mS�|�3����nܔ���/D�@��H�NU���.9�q��g;D���C��zP�V�Ԟ@�*l�;D�L��̂\UdىbaN. �5(Q#<D�4x�j�)���b�:z�ِ�l;D�$��؈H �d+�`�lՂ��cC:D�|#Ƃ[f���̛�B�U-;D�<(��G=bz�Q��'r�B�*�:D�����6 ���0�/�s��Ѱc,D�t#W���](\��dV�,��[�$>D�����S0:�,}�� �;��ԛ�0D���e,�9 Z&�XwEB�)�t�V�.D�#Gt>��P�]�l�a�/D��Xb���gu� �寜;"�(��."D�0�'��8g>��u@5P���I��>D���)N��#�)#����3�'D�p)@MQ%�RĨ��"j�$qTF#D�P�qEҴGj*��k��o��ś�J D����gI�v�:��5��+����A4D�x���--�:Qkf3a��@��1D�ȸS��*VÌu���»<s~����;D�\q���S��P��tv")0��8D�4��J7>u���	�be
ţ�8D�x���w�u@�mJ�9���7D�D�g�W!xUh����|��9�Ĝi�<��*(����L+	a&Ă���\�<Y�'�:έ`�ͤZ��tZ�#�X�<��L:��ň���$�Y���S�<����0(h�H�E�1��bU�<�K��.����OS�Fh��R�<���,E�XQ��ǈ�p���pI�f�<9�H	C��e��0�BJ�Id�<y�H÷v��	iƋ��I k�]�<��և&�Q`q�Q�*�:�hD��t�<Q��až���k��x`aڱ�Dl�<i�gZ�s�逡���m�4�!���h�<17�Q   �P   �	  �    �  �&  q.  �4  �:  NA  �G  �M  ,T  nZ  �`  �f  <m  �s  �y  ��   `� u�	����Zv)C�'ll\�0Kz+⟈mڄc� 特m`�DB�6%p� �f�q�䐻"�m�|Mi+��.�c`e�	��IuJ܅b�"I�;0�4���'Y8��J��}��1c��)U����	��l%ʡ�bC� b�Ԛ�@�����B&� 9� ���X`�-��H���9���=vr�,��$�3b��4�WEXB�b5���1���G��z�*�4yir���?A��?A�⌽�g�X���`�r)X�������?��й0��F[�(�I)es2���O���؊\����6&���� T(�����O�ʓ����O���'	���O����tI���R�~��AY�8�O�牐�>�+�&�)������۴0�(��y��,���I<Y�D���ⓤ9>i�1ӑe��D������I���������q��?�P�wB���Q� �$/��5R��'~�6O��m��4כ��'=�6�	�y�޴`����'��3�
��K���{#��<���*�� �G�?}� �Ϊ'�0�W���LF�IX0�����@��m-m}[��i��6��1����u�?���lY�Ik^��5�<"�J�A��;:Ȕ7mP�K�V�i@DN�Y6��PA�,�D�tk>E�mn��MG�i���Y���` �="�5�j����B �ŷ!��7���ec�4v� ˃G�)�j��!ǔ(���@�֏�V�K� AO��Y�*M
g@x��pB��\��	�´i#^7͎Цu��\�Q�qR�,� zR����G(3~M"��ڵ��p���_|�,�I=^5��u	�"s��31��
d<|���U��sA6y��N�i����9=�6][U����2��'���'	���O����K s�I��'xD@�P �-nY�T��N��]�R�:Q"O�mA"�\�VƁ!�Ə�7��eB�"O����96��3R��-��%��"O���#ȁ1�И�F)��D��S"O��Jq΁�.?�	�R�7/��,	A"Of���Aif��Aj���j!;F��fU��~Z���<�n-�4i��	��y�5��c�<!v�@�U��y���G�]t�Ѣ�v�<�f�3Y4��*ʢK�H�!ʞt�<I�͝�3Ft(��͠q|�02�I|�<g"A�������ic�c�t�<	�mS�f�(�n�>�h�AR�����3�S�O��lٱG�;C"�,�B�:.�ʧ"O���a�ލ+�D*4��:�F��q"O(�#�>�:��R�� ���6"O0|�D�K�%���*�M&��"O�峕�O?CMh4�LZO_��z"O�ep'��8j�XaP4+�.2T��X�<�r�.�O(�LN �0�"A�C�(��"O&	���Rvސ�AaJ�M��%�V"Op8��K�3s��
0��[�Lpu"O����MD�ufp��Å0����4"OB�a�m�d�x��з��G��<y��X�!��������J�x�2O
$��3#A�O�ʓ�?����t��$0�npʂM+s��!C ���2㟿e�X��B�6�t�)��I�F�J:c�M=���� :B�rL�%�z�:e"��C,!s�,�z/�� T�ɏ@�F���O�4oZϟ@K2�žM`�V;dI�Y�3GSy"�'��	S�OO�Ɣ;� �S0	�K.Y; #��1!�$e�����.\����G*s� `P�f�Ox�D
ߦMr���ß���sy���y�2O�T 􎐁CJ���Ba�>�XQ��R�ϳ>qO>�ف� �3ܑ�&�^�K��i)��;?1*Ƨn���"|R�O�F����N�9�H@�ľ����q�j�D�O�c>��N'bhR�Z�o�J<�r$4���O^�����j�
tV�na
3���a�џ�Q���L�WMJ,{Şb��c���$2K(S�O���	k�,@@Y�~ni�%�Ҩ";<B�)M�Х+0��\�>��"��:-�B�I,}c��zu"��c��|`V�P��C�I�=��d�h^�+J�]��I!�C�	��lE�$�"V���#���
��C�	����0�˟.I�Z�ASKT(��KeJ}�Ć�d����P��*O&6�8׍v�p7�?����	<kD��"�[;����W�c��C��=
kN=xw�=T$*�j2�Y;s%\��Ӣ�O�̇�I	|%P�8�@
02��M�r'];��Ǳ*5��h��'eI��a�h�vr�'�`6-1�D�=o�`�$?�a#A�B���z���o¤�Q���OV��?���?���>׆$�'�%^��s!��� ����ۖ4���艟rb��*s�4�G8�l9��O�^b50��1eڽ�Tgۢ �8��0��	f��1.����Ox���'�򚟘�� �Ca(�!��7	rte��A%�d�Oz����T���A֫M1�89��+]2�O�O��(�Ȏ}��S�B�_������'��	$O��2ڴ�?�����iI4��Dд2O4�
���(_�0RR?���D�O\��c��Sb�z����(�T>E�Ow�(�`�f��s�k��+�\�X�OaRT�Lw�-r�Î֨��tô�F�v�t����2 L����O��lک�H���)�7<��ѳah�"X�r#���XB�ɖ$1��X"h��("Mh��[=?�N�?1��ӆ!�B%'��q�Hd��E~��8lZ���'��D�a�X�$�O��$�<	�����	���RV*Y�������8.:���\5T�N�(���)BS�	8�䜁�*4:AF�2i%~��0j���	 |�� i]�!�1��ORP1-�4_N�a���U���C�'k�6��O 0�*�O c>��?9�%Q�+� �	� X&xC�j����d0�S�O)X�V��>o �b�d]?���I.O��m��M�I>�O��	=vp	��K�d:Jx ���}�z�*L��M����?9���|2�O�B�pE��f�% ��Hb�ٽM��]����Vm�ق��N�џ�\c	J3�$Ul����J��!�X��0�F�jm��s���iږ����%5s��Gy"'�u�+��
F�d�I���0����?�b�i��R�@�	Qy��?��TI���V9`��Y��*��6�OJ��"��7<�	1��	�(/���'�6��OUm�ҟ��|�	�LF�H�v����d�B<��Xj�J׏� I�ȓ�T]��n���GC�^���䊵� ��9��=;�F�"p�ȓt��gC+7��� �[�Qoj��ȓ~�^%��(�,(��S5PB���o��P*S)��Hf�
!�XR�F{�'D�̨��9��^ }Ŝ��A*��wR���"O�ܛ���O²`��7m4��c"Oȡ�r2-lI#�oÎ+���R "O>$���B��0q��Z�`�� :"O�T�0`�Q?�=�Fni�X��"O�Ճ�i3L����-�>��d���'a��8���7$� �#CҬJ�R�8&`F�n&���Exybe+I4%���u����o>~,�B�͇~onA����P�4��8�BL+e)�1 �UY`��� ��ȓ$^p@{�;w;΅`������ȓK�^�A�S(M)0p�ە9�n9�'^�X;�)%I�de��8�$�7g_�-��A6�Y�3H�	8T�zj�
 �Ą�`�	(���:+L�" �!�D��ȓb�ڶ@�p�-Ąe4:���c�R@#rG�.��сD�ԥd�Ņ�	5��	4��Ȁ�@�Rs�� �U?�B�	8"<R��3\_�1�6�Wt��B�I	P|��VI�C�8����U�TB�B�I&�<��%o���G���a�nB��0JJ�$8�"	(�[�O�2x �B�3%"�s�����ѵ&]ZȞ�=��}�O�:ܸ��j�&�Xs��=>&�B�'r���B��J_4E3���0�&;�'�
�����p���pKԺ ����'� ���ΰs{�e��l�;i~��'14�X�+��g��C@�-��c
�'��)y�$�m�(�C�R㖝��X�||Fx���I/\��,�Aj��5�u�U�8�C�I�\�Xb��ω(�^5Ps�S�J[�C�	Pl�I�튦a�Hkmѯ}�&B�	4>�`�1v`چ/��D�P�mPdC�IjwvM۴�ʈ�&Q����&C�j�*��5N57g�{"LY n6˓R+"a�����(c�*K�*�"��C�)� ��ZĮ	�&4S�n�*4���@"O�9Z���24ҵ@$��*+�P�0"O"0kA�&?74�Kc��.t��"OP�� a5^�[��H�]Ӗ����',hP�'j�d�s��%^L��u+��4��'�hr4EY<E� Eo�bO��3�'�H��I�l#�'�^A~���'�FpE��7�|��D!#?���'8�U�ax��U�cF?��T��'����C��am��2��Q�v>����d��Q?�h�����(���L��aZ�!.D���d!��U{��sd�L�fy��K�9D��y�����t�4��"6��1cS%6D���e@�#"�U*�HM�6�~���6D��B��!�heHV"�a�
YR��'D�a�L�_�& �flG;-1�D�P��Oz-��)�'!L(��_<F��)6`�',ҖDZ�'���DրE$�"�D��:�a�'��|�P���_��,He([�<�2�[=|%�DR�e*��k��TW�<���d�]��f��ea�T�<�T�Y"8�
U�e׶O�\5x���Ry��+�p>1 -C���ʆ�ʵ��)f]N�<��+���D�χj��i�2�DH�<��اs��12EoT!,q�3��G�<)�e�,t�j�m��aB���&X�<�5�A	/���:��8AU6��⪉Wx�H`E��8��_�6�Z#\?��;A�4D��	q��$��)'��FƆ��e3D��c%�8K�Ƚ�g��,�z�"1D���v��U����C
';Uh4�� 0D���D���1�l���Ʈt�*p�Ec D����.	-gNb��P�)��SEG*ړVK�@D�$/�F��4w
�}���G���y���;>��a#�W	n�s����yr� �Fd)�R�/Pت�j6 I0�y��P�v� 
���O��e����yB�Д6��p n4L��1["�P�y�� b��q4-E�/�xҪ���?��F�h�����Ո�π20 �o�@���"�g%D�`�ƥ�� ��r�mK�F��o$D���*Q�PR���$��MJ@�J3�"D�(
��##t0�kG*�B��>D�����Do6��7�@�?jr(�A<D� ��+ʸ	��7��d���<���C8��A��ݍC(� Z'�� aB�\"�(8D�$X �M\C��Q�̡U��SrG"D� ��K4�R\�sb��{ي0A%�!D��z���n����
l�p�>D��C�!��erz}���_�B���R��:�O$-� �O� RF%���>��0.�9;v
(�#"O������A���P��a�s�"OP��d�_8J��d"�E k��K�"O����!O�/Lxsu��t���`�"O|D��%R
)pDE�$�
lO��	`"O�A�� H�m���F֌6�ځ21�	�o��~��F�I�(M@�2_�LҒ��B�<Q������0���^��� ���v�<�p��>e@ܨ�B�� :�*]�ȓ|0�y+D��~���4H��n���>	�Z$�+{�t�X���
|$�ȓ.`>�gb� � �R*Ɖ3�9�Ʌ٘#<E��N�1��lPj��r�$q�S�	�!�$\,E�ʱ�d&�����!T�
�!�� ��)��!<Bp⇭��-�>�y�"O.���cǚ2>e��͉�cw@��"O�hQ�G?+!���E�*`�S6"OVm+���6Ծ�3��"�yQ��  '�O�)��Mê2~<��E���M�"O�͑WG�d���u�I�a��9��"O����V�M8M�D�4/�@��"O�]13(�)$���AE	H,2���"O6�@a�"y�biI�N��Щ��'�.T�'~�<��U���{�e�-u�\�y�'f�mz5咽O�~D�fH�0��T��'3�m�S䖰W+��*�.!�&�s�'�t!�@%�z�ąkENCJ�
�';~� bɇ(+���ڙ����
�'Ǣ���gslr�˴'N�ڪ�+��DW�Q?�#�,ȋEg&�2�:yq k(D�|T��q���b����{	*D�$�F�(I�y*G ��:~�(b�+D�LZ���#�"t��E �)Lp)��H*D���dI�l�lE��\(W��8*�"+D� �ٝ{���4�A6�Y���Of F�)�'f^��q¢]>n�j��s�RU�����'c�mK��[���#�M�TD�x�'����'U�Y|E�@zkt8��'��3��Qp��07�P(h4u��'�.4�R��J��C+X%xdB���'�L,yk x�8-�d
e�l+O�C�'�h�����13�}��Aèl�#
�'⁓D�G�H.�� $nzǮ<�	�'�su�1Y����y���	�'@���T�O!P��52�]�v�\Hx�'�j�%���%��!�R�&eff})�������Aք�=���s��{���ȓc��A����3��`{Q��!���ȓ&c�Yk0 ��~B0��Wc��,@�ȓ[?��b	*Mو��c��SU@���cm���IB%��{`c�\T&q�ȓp��ㄭԃ^�@u{�"K?=��mD{B������8tI[�P�jy���^��"�rE"O�Xs7�[6&�i���'ͺxK"O�L��`��NÚ���P�j�"Oa�tm¾$��Ac��A{G���"O<��-�F�D̊�&ۜ��ɛf"O4P@#�$�UI��V���e���'�Dݻ���@CX���m_�� sA"/�B�ȓN0��+��J��8� M���Մ�$��r� F6T(t��,9
q��fۘ���ԈCm��HO�x�@�ȓsLLр�kW�$�Ƹ� W$?�n��ȓ�h��OY�U(�=Y�/�[��ї'�\S�I��	V�?f1ir�� ʡ��	#(�S�V)H=�1�d�^��܅ȓx�x(BC�CY Vjb��a�A��m���#��>E��4qvO٦El�Ɇ�I�:,��H@�Bu�-�s@]�k�����h:��*Yx�!CS!28}R�M �C�I Y;��H��͹K5��!E 9
�C��0l���g�.�n�PsF,	�vC䉞rD<1�j�2T�Ҵ!�&6B�ɡ	e�m�VIR=�:ܲp�K�C䉪y���於��P�ǐ�_)�H���0�z$���;
����rb�D�ȓ~�"h�"¿?�8( 'řg���ȓd���� !#y�4m�� L+�@���S�? ��R���M����FBWY����"O*\���A�p)��^��L�q"O,<�W-P�w_
m����t�2�$�'*������S5k����FR8����%(s�8�ȓxo@���_�3�H���i��B��Q�ȓY��:P�T	Et�[Wk�� ��ȓ<	�IS���<�����r�P��ȓ?�� �e��]��,�g M�!2N���9`iy�͜	�6�i�C�76h,�'�ڹ �g��E`c�!&��y�g����5�ȓ>��=����/5�TŘ���m�2��ȓr09� ����X�Ɗ�3�\ȅ�%�\5��D�-'�:!�l��ȓ]=�@P���xJF�[�N�?2���I�M��ɹ_ܦ9PV�j~�5�vHɖBwB��* ,SN�k~��e��/C#B䉦a�by�Ff�C�Iس��')��C�ɤ;�u���N=���s�� �C�	�z=ҙA�˗<Z|j��F,�6chC�ɩM����D%�16V)���9A���=a���S�O�`Ʉ)34���6�( ��'�H㗩ֳf@<�h4�
|�L�
�'n�5���T�'��l�@�^$yT�p�'TT�a̙6A�[Ã�;k+�� �'^rQ��h�lHZ ��a����	�'����HT����R��L�K�x���#v�Dx��	$5'4̹!��
*�`p�C�U8B�	r��A�
X&��]�+,,\
B��M���ޑj��=�Ph@>P��B�	
}�2	��{g����C
63ĪB�Ɂs�vL�g��,2��v�y�B�I�8��|B���2E�T�̒xc>��=1H���b�J?9H�x�w��06�CqN%%Z6<a��	Uy��'���'DN�ӣj�����o�9Ai�Qb󟮝K2H ?p���d(D!Z�t����!D=Ե��^-r��I׭\7cd��r�C�� �&mE�H�]&�����-T�2����I�f���O�b>I�����.^0D��΍�>5�xKSξ<��wu�aҏ�
aE�LCc�}�j���	����ѩe�H=���jP�5���W	9���!|�^E��ҟ���d����Z��'�j�R��C4���G!Q6����'E<j���P��R7�DO���T>��|b�N�md:]8�L� svJ��2���<Q� �D��d��߸�Z��I�>q\��A��h!1�X2 M�d;!R�'��)�	:?A!ˈ�!�z�D��:	Z�����H�<��FL�JI$�*Q�	 �e�P�B�'��"7K^�!��+PB_9���䥎��?)���?�3hÔ#?�r��?)���?�����d�%�����B��rp�_K��������Ò41�)�4�<Fx����Y/����< B����d����':z��8N��i͟��DK�%(d�����I�`��)5?Q!X������?ٜOp�Ԩ���,w��u�5	[:@=�U��'�f����2A�i�NO):^Ȝ��0A���Sٟh�'a��@�鈶2�2����A%*-@1&�9
�L�(��'�b�'s��h�������'q��Pa��;\��rM�^]���B��%)P4�ǅ��X�F�'�h� ����=y#��q\z�@�y��V쟁�� cs�*,O��+�'oy��/� � E����]��@�P�'����3ڧO=
���	�;��ZD&͚K��	�'��X����x²uZ� �!HD�I,O��)�Ir�:�~䥟�p7H�	j���s'��L_>��@"O��`�$&��Ex��T�bkz�Iu"O�SPo��8�<0��F�=}6nYX�"OTX�dI�:g����8º���"Ov�҂L����+�dĪ�۳$"O�hr��/~T���.f��t���D�+q���O6z�:�ٯ[&]���V�E�\9b�''$H)����a`ˍ�6�b\�	�'�P$p c5\�J����6qd=`	��� ��5Ђb��Qx��PY�EV"OЬ�ѭ�$}��5�2�.{�6�!4"O����)j�0u�!@A�28\P�@�΢�O��}�A�f��D�I�Jȶ�C���ZF��>��kB `�|5+@W�Z؂8��	��5�&���A<Х�gf΢44t��(��5�wL��MC���#�(u��ńȓR-��b�'@ a�;��>)�h��ȓXX�����V7q��EM�W��<�I2Q@���d
�E�R��/'T2P�lZ!��9v�䃵L� N������%�!���~���K�w�ʤ+_�!�$97vbPKa�� �8�	�m�!�K��q�����%2A��џ,hf���M��?�O�� *�[�@�$��ӏY�]��K��^�H�Q���?���\�B�˦	Ir�d���ITY�6=�2���L�O�Ș#W�ޗ3������7a]v�I�+� c�"L�1aU����!��127���4�b�LK%x��##��O�#|���Վq���CS�ӔAI��c�\�<�� ��M�EM�JZZx���.OZ��=XB8�9'CE
��D�#V���Οؖ'�O���.�P�0���rT�Y"�Q�Pׄ��:�|%��C�-Y�,yx#��[Rn��?�4�ēA�8b>A���Ԏ.�hdq�6z�y��(?��O��q#�>��y2DJ�@��{4E�41��Z��ֻ�65[㓟p�I���.}Rk/���ck�8hUƆ�n��t�!-^�C�ti�I��a�'��>�	KG0�C"�$dߔ$�ƀ̋aHx�dD>}�"}�`	��I�����pE�-3сv\��s��A'Ę���I2�N�*R���F���cb���6�N��놫�?Q�(@��v�$ɷr��V���.��B}ތ����)�$����)��$��c��sQ�?����?A^HQp�2Ad�x0��{��I�/�ҧ�9OhT���*�&�5H^�ʶ��`�T�⮃�to"T�'*�mJ�O��x��)�r��cR*D�;1��AIɸy��@C?��MN~ʟ�dSq��$@+V�9!ꈁ}�i��8N�2�_؟x�uD�<u2�)���A�R>��2D�.D��)ai��q]��h�
(��lm��4$��٪���O��4E���x��E V��k��^�Jh�&T��$�tG{��	{���g�H(�C�0P�d���"O�%�P#�\�d��SD����
E"O�#��JV�-�d�3{f-a�"O��k�#�/���"ʆ~eP���"On9�W�M����!/�5\v�4"O4A*I-+n��b���"O���៫(�h�3-:c���(�"O�L�d�9Ȁ�5+K�6"O\Б���<k�0���+ި���0s"O4�	�Y.Yt��kC��#R�0�"O^�JtM��`@ ��d͎�	�"OXh�i�>P98��ad�/\T��"O���Z�I������,{��D�dZe)«^���=�FN��<X�v!V�,��}�gꍋ	"y�QL�sͺ%"�֬k���8�C���<��*V	&��쀑=J�ٙ�K�O�J����۶_�&\
�� E���1�0I�|1���îF<�Y��J�P˷l�(�$���t�6h ��j�>i�dqQ�%�=[O�m�tc�7x��B�	X�lL{�	�<��@�K�G�hB䉍:G�H #�Fֈ���l�2�C�ɼV�
�%����9�L�Xp�C�	/M�0�AB�F�݈U:�+$-�B�;R�L���-����"��+vB�	� 	���h�1B�����x��C��qc�� �B�m'P�J��^,;ΚC�ɫTl�IQ#b�.f_��#���bC�����yPe�~ �0+g(X$�ZC�Iu���h�P7(����ɿt�B�	.7Ťd�!�ǖ������E�I?�B�I�x�Ɲ��"#A���ڱe�8{!B�)� xys�w@�����
��#"O\�z��?i��	vLQ�|�~���"O���'ď$���K�7A�:��`"O���`J%z��S��;]|�x"Ob��Q�K�y��H���7�<��""O���`bB/Q2�)BW��7�H�2"O�P�*�T|���ӮH��Ss"Oh��q�W��p�u��bD 2�"O�y�ai�4��"	�7C�}Z"O ���˒+-�ry*RF�#8��%"O8M��y��\ �ZEs"O����;O̘a�K�$5�U�"O�vH �����	��q�� S	!�F�"�Tepօ�!�&�yQ!�q�!�D�6@^)a2�ܻh�"�)��NL�!�d�F��ѱ�I�)�N�P W h�!��/�la� [�XЬE���0q�!��
t���&�lDR�b�2�!�$V�(G�pC疿u-�}�5O�}�!�d�h�ˤh� L�x8�߄�!�d�!UfV��C�^�&���)����!���*l¤��2|���h[�8�!�V�S��(7!ގES�@��gOi!�ݽr��)$�XC��ArM̞Z�!�d7D%P&�E� ���P��ս-�!�d�Jl���K�C�,��3Gو�!�<q�,أ�~�<P�fV9Uk!�D\#Z��hfA� +����μ^g!�߾J	X�AчH|�� @*[��!�$[�z���E��dj��xц�t�!�ΪU�\��&!��ze�4�ckB?�!��	T"��p�䕑:�v�jBj���!�d��d5��hM�'�q8�+^*�!�	�}�d�0���N����7��}�!�d�@2@���ڷ���D��&�!��\��H��
�J�f��	�%�!��=~F<<q�ʕjmde�I�6�!��&2���h��7&V/'q���"O�!-%�Дӵđ�c>Q�
�'��ժU�է_�� �fU7����'T�8Pe��`2�tI �)b�p��'����G�3J��Y���R��<��'�4���#�	GT!@�(��X��'���H� \9Q��ǡ��mR���'���`�Q �B�ҡ,�h2(tc�'��<�$�X3Fm�l �È0�R5��'���(F��r�NN�QV�@�	�'G�At̏/o�0���-xC��H�'(���`啪*U��PR��*#��A	�'$dɱN�"T�4PP��H-j- ���'����/7��<j�ɂ�`H*x�'v�����Ύd$����)c���'��]H�BP�@>���й`8樒
�'Y�HX���C����)X�h��'�L�����T�A��}:�I��'�)Z�	_���Q[�ɍ�|��|+�'^d��'�1_FE��Oc,d��
�'��1��Ї�x�S挐'!�
�'�$�CBDR G�PE�0h�
�d$z�'�ƥ���]���E�;m�~ػ	�'X�ܓ�k�:i'���`���;N�1��';�J5'D;k���p��.��h��'�^��Rh�3#��ʑ��,��
�'o��'ˣd��P�Q^4<�s	��� ���K�Gft|2�K���"O���a�����bg¢ ؈�"Or`9W"�5�z����>��r'"OB ��Ԑh3̨*2���T�)"O�I9f$��
��qri�+��`"O�!�(S3
�r�����T�8�Ys"O<���g��X�0�`�*�*OXH��`�\��:�g6@��P
�'Vr�fk�/=e��ҕ�?�z
�'��Xq2$V�zش2rD�=�<̺�'.p����9}���4L��.��9!�'�=@fI��yAoܘ&�ތs�'����B%��0�=4�|<��'��D��� 2�u�� (�fE��'�XU��b	����Y��B�ꈡ��'B@d�G��;JF���ĉ�j���'��Y�Fl@-��QP � ~��<��'��<�u���4@�)ҥg�h�h�'�,�sB�U0��$��g;�A�'�ju��B��BPY3ˀJ�.���'�����H;?	H5��BH�>7(h��'��u+�J�K�=F[(:��y�'0�$�LZ�`ܚ,X�X;
�'r6��L�L ��)!�S0[.�q�ʓy�xą��,���B�!������3��I�<�X���f��&i�ȓ] d@��������j�*C�ćȓ	*^�b��F�;
 ����ц�� ��I�T�%�d��MÚ����LU��հ0@�|�0��5j����N��H� �4܀l���'^�6y�ȓh����,į;^V�����\��fe�����I���G�	�3Q]�ȓ0(f��q�9,���:�냭D�"	���}c	A�E*����lH�l� ���pXe����~U�Iz`#��>�ȓH�F�`ҿ���I��׭q��ԅ����j��ѝn� S�.N#�Z�ȓM* �ЫVÜ�&Ό������gm�4���`ü%F�݄f���ȓC��ʀi�"ڠ��	Z=	�e��tڤ1��c�N��)sΚ>&��	�ȓ^m��h�0t�����>~����|�h������Y���̷GNP���:8�h�\�p�6���5r��ȓwĠx��kN�S�9�B�'x�"Q��D�Q�#�*ihuu�[�JH�ȓn���yB�VF���DL�v0��ȓ@��L��:/*���� ��E�� H%�b��4r�H�Q�1#q��ȓN�X�s�>�0a)&�FLj]��Z-�xi�\�Q�v�*Ba_�L����ȓy����>X^�j�疳>� ��*��r)�.�Yt��M�x��v��(��dݏ9:=@�=h/�a����`�uꉘo�0ĠF���q�ȓ.6Vv�7]6p��t&�A'�܄�K�B}�"L*%��SEHN�E^�Ʉ�M�\m@��2�h�&��S8΄��}m�!���"��L��G�7̴��#
���!+}��m;g�^2��ȓ?Y =÷ ��#�
\�ၙT�Z!��y�dيG��/]����_�R5x �ȓdF�ծ��r͘#kQ[�j���S�? �P�,��JEN����(\Ș0f"O2�:c�IYB(�e�q��٫Q"O�A�f�?	�B�Y�bNd�"�;P"O.X+�d�(�vDrrˈ?+��U��"O�z���<~͂ܨ� �>����"O��B��B��\�4NZ�~�V�qd"Oݚcn�X��5	b�>޾�2f"O��L�"/Ў�r�j�2����"O��``F48��BQ�W�^,�6"O ��&�ր+ D%�"���x��mP"O�y��F?q�\Հ	]�()"O��&�^ 8��m#'ϑ�Z��"O��k3+؅n�*u�EG.2��1�"O�(�k���O��1�zR�"O ����΋h�<K��m�Aq�"Oz)���)T��I+��=p<l��"O�9 ˀ+���b`i�%��"O�=IG��H�������W.Yr�"O
iQ��ÈyD�suA�RQZ�e"Of��Q-��a�(�Z�/�?k��$��"O���
�;��a�`Q�=�����"Ob�d,� b�tq�J�G|xU��"Obq���юd�$Dqīyu���"O�	�'Bۡ*�4ܻ/
 r�̊�"O��R�߷$�����o��qzن"OT��"^'HlH���Ƭm��ca"OV$� �"H`���"�_�f:�"u"O�9�6�.B�Z �eKGd-�"Oh�2����T����<;E�Xq"O�+��զ\�Υ��H�o�L��"O<�AVGq0�5���W�|b5��"OH<���#�X+dgYx8P��"O6 ��J��n�&`��[?��#�"O���o_��Q���{/�)��"O�4z ��Z���ҧ�����AC�"O�� S�=� 䂲�D2�j��"O�1�"��O6�(�bϟr�N$�7"Om���0����_� p`�S"O� p�O
Fr���U(�1Z`�x�'"O�����"R��xg� ]"���"O�p�@N�X�*-�pe�~o�Ty�"O��Q`��^rr�i!D�0fz��7"O�U�1���l%��آ��eZH<��"ONdB��ҜnojU@�W7F�L��"O��ؤ�G咐� �zͩȎ�y�Ɔ�S\ �##N@;��`h�A �y�� B"Ver�ڶfۄAJ@"��yB �%F�h��PŖe��X�K��y���E�Pԙ���,� j��
��y�H�q �ؗ.X� 0q3#���yBNθ7��H�%��`��x�U��y��� N����͙4by|���%F(�yr�(K`�}�6ȃZj��H���yBh�0�M���5T�V�P�L�6�y�M
�dnБsC�M��U۱���y�>_�D��t�@��P�ƫݙ�y�g��>}8�!ɞ5<5|�21+V���'~��Ȁ������!h�,�K>)�!
�}:d-��B>��rmd�<� ��>M�I*A��K=_�,��'�~		F�Ր7tQ�c�
;\x� ��'���l�+N�<PZ���%g��'l���$�T�IP#�gѶ��
�'\YT&�$c�T���Pv��`
�'9�Q�/��r��4 �ȣ=�<�
��� &Dq�hףdz�2�!��+ژH@�"On	&�M�-h�u!�4��,�"Ovɣ2M�1��;�g��m���B"Or��B�ڣP~��ކv�P��"O��"
�>�`�O	�vfҨ�"O � q_�3'�4��-�r��9Qw"Od�D�PF�d���앻
wLi�""O��m�m'�$�0# ^��x�"O�U��4E84�c cɐ- ��8�"O�1�1��C���Z!�ݜ@�\�q"O��ǬśX�V����9u���v"O���P�T�] \����6�:��"OP�q"+�-lf���g6��4��"O��Xd�3[�Ȝqvb�p�q�"Oм�oR�X��I���*|hx�"O~A�*�@��D�.�."��""O�u�mί����UǍ	"��c"O���2�D�K��yӰ��].D�g"OԨa6ȁ�K8����c�B�4"O*в+\�C%xqs�dǸ�""O>T�Ҍ	)ܼ���]�N_j���"O
�#���n$�9���1��X0"O����V�Wh6D�@�T�#"O�����E�`l��C�� �/!�	V�Q���7��1#�!��XC!��0+�̰��`!��b����!��_&q�Fف���uk:I�g�Z;4G!�$͕=�$��ĄnV"\QԦ�$e�!򄝺3�FDy�m�"HK*,i �V�!�$� -��V�^�eWJI[$��#�!�DZ�fƎ��-� T� 4�W�޼/!��4l�MK�E�$�b!���I�@�!�d��eh�q�5~>(��E���!�^�)����D�2V>�P��M�%�!��a�����D�x���7�!���a��,L�!ihI�n�c!��ÏE�Pt`�HвL�h��j�#v)!��d��@5L�^[���`Wc�!�$ˉW8��p����nEt5���Y`�!�D�~�ԱQ,ڰp�m@7����!���	_� v�+wOH�q��Ѧ&�!�O>�Z8k���B�)zaKF�$�!��(ꅬ�(<P-)��Ȑ�' �%��>�𼛓`V�p��h��'�\1�@U�<^U���ѳY�l@��'i��R�?8�UA M�q��'ɠ�UǘYq��HVAͭ[t���'�p�xe.S�d��x����Rj�x	�'.V�H�(�(0�i�¯C�]��'K"�A��0Y��!�bD2u��%��'�� �V��!Jޒ��4�CAV��#�'l�C�O�"��T�a��-��4�
�'���1Td^T
��c�Q� ���	�'j� �w*Н c�N���%n�}�<���jdL���J��i�͋R�<�A ̀=��!#��[�`R1���m�<9p%Ԁ���������H�e�Zu�<9B�!����6��wi��&čO�<9�/�{#Pa �Q$�wJ�<�g�E1M�`���$U�ЉF�IG�<v-3��А �P��%:Q�VC�<�(��fuR9�wF�9zD�Q���M]�<����F@0�a�@�2Y �I�C��X�<�� ��v��"#�)-%̨�LF�<� @�Pq��7D� p7��Fv�1�"O���'h
^<{0� i�t��"O8�"�"	(k?�Y ���6$�!�"O���ϐ9~�� �ַ2�^��"O����Q4 �8��Ņϸ���0"O�x0G�̹}���%��Q� ��U"O���lQ&8�F��@���t��"O$$��IK�7�,���@�NY�"O�Y�V�[6~�Se�^����k�"O �Uh(������@,F�<-�u"OU3$j��W���Ĥ�=s1P"O2}ZƆѥfGָ��O#bh��A"O@Hz�+P�p��-[�͆5W�aju"O~��f�����	G"�f�@�b"O��[�#�!L،8��2r�`a`�"O�����Jt����HŁ��4"OΈ���Wv��[�
 &��Җ"OD�sJ��%���T���dX\K"Oj��%Z�9�V�Ď^B=("O��؇���(�;�MT�kG�h"O�� ޘ+V�����C�D� x	�"O �x��9U��`Ze	3�8X�"O$s3O"Р5�4k2'�H�"Ot�:୊�O�����i����(�"OL(�2۝]������W��()�"O�͓E`��?�fL�7cܑi���j�"O�����>���85�m�"O�H�
1{�N0y#�P�*��5"Ob�S��>hO���C�p<Q�"O���PÙ0f�m
�J
9�4r�"O��k�C�%&�����/�t�ñ"O�,cv-݆�H��'EMV��AIw"O�#�)�6�&��s)�==�;�"Ol�#n�&"�z�k�h0O�Z�*�"O���6��5�L0I2�I�.�XHV"O�	��B��Q�(��3-��|�u#�"Od�z)�t�5y5#�9�`���"O�p��*�,4#1�
1z�� Z�"Ort��V�&�*��/��t�"O20��׎57�x;t�¯ij�e��"O��Ĥ��mƲ��4�	g����"Ore���+%y@8#@��;\���"O�H�-@�F���oҠj���G"O����$[R���ΜR}����"O:D%��{XD �3�S�Vξ\J"O�P��O<1M��#��2G(�(i�"O�M��� H�V�z�eG7	^�X�"O0�S�'�y+���W�
nL�b"O.̋W(�7o �#�*�,EQ~���"O� �)�n�}��#� i�X�#�"O�arGM'�����,�h���)�"O����*�8�����8f�P"OP��T ��j����a(��2���2�"O�(���]��谛��E�8�t�c"OB5�P�Z"!�^i��'�]�x���"O���5��k��,�v	�g�.4��"O8 �KBM�(��"�S%I���5"O.����M�n1"	ۑ ��$Y0"O��@sM;��<���L:$��"O�Ԙ���]�@��Cd,��"O��ˢ��
%;D���G ���:�"O����Y-'����g�-j�DM�"O��y��[:�.u��޴j�"O|9�[�f�*�srJT�"�[�"O� �`c��A& }��������C"O\��3g�3e�\([��X7Vh��j&"O�K��Rx%45��acT hv"O6e��̛(
� ÈU��"O��j�Ë�\z�`'H�m��Y�e"O51�I�4N�%�l9M��1�""ODT2�#����Ӡ=j�(4�S*O9��ʇ+�T[�FpM2�'HI;���J�t�1eŔ4���'�0\�6B:6��T�!fa�B��?DjZ]+�'�*��=	fJ�$y�`B䉾3���B�,�2anE��S�|��B�ɰ2p��W�
�M���QCаT��B��5>pj�⡯���d0G�"��B�ɺo�|2�G �@'6X�B�	�Ni���'V�.������A2ԚB��62�>� �R��P��#F.pPB�I�)I�\2�-�0�4����=J�\C�	/E<m�-�]]J�P��?k�B�I���}23��P��y���ʒ&pC�ɑD�VaM�Ll�������P� B�	�_�p1��F8�x�apmQ�z�BC�I�C��@��
�0h,nAGL�&C�I	CNMX�@�\|�p戕j�C�	�[��	IEBޯ6� ,@
W _:�B�	0k�
�gl�#!O�MT
�~��B�ɧmd��cH�?f��i��װ}֜C�	�<(8��앎c��쩓���RB�:h:+�='QV$��ՋQ{��P�'k,�c�H"`	F���O�4�̼y�'��	4$�:��H������ޒ�y�`͡[���Q�	{hp�X�B��y��A=v����ٹteĨ�uI��yB��M|�05�]Ѧ������y�M�Rw��� ��%��[�GP��ȓ-@���B(�l�8�0��g�rh��V��Թ �p�)��ȉ]ӌ��ȓd�D���\:�B�3fo�)�ȓl�v�HcIW�WvQ	U [�qr��P}dU�'��4X�zy2�I*����'�,�k��
lt%��_v�����!�h���PU���ŇU�VM��,P,Ms�W&�&������i��.���gg�duI�Ro�t� ��ȓt�KǢ�4"J:(�0��e���ȓ]]v���h��t��@�t�n���D�4L���0��Y�2��D��W�r(1��?��9�j�\Q�Ą� �@�[T(��)̰�B͝�b�fY��nB�����-U�@��OC5$H���Bې$�c(Ӗd�����
3K`m��'�"TP��^l���Z�-	l3�m��v'�#�n �VM��N�1K�,�ȓw�i3��ME�.�2�K
u?J�ȓl�.���@R�C�d�8�K�K�
Q�ȓ??H�)2��t�*��bD���,��ȓq�@B&D9��p(�L��6<Շȓ-? �{V� ^�Ni��'//�F%�����`��S�ipv�!�ì��%��ih`<Z�N�6`�r�G�V4|l����X���������FC;&��5�=�#�w���%��5X�$���f�	�-�,	����FȰ&��5qC�I�}d$T���H�.Z\|��76�$C�I'X�֔�l5#(�E�!Y�C�)� �ZQ�<��a�v��%*p!�"O8T"B��q�� :�.A�~!Vp�"O^���ɖ[>�+��R�;9(LrQ"O��S�̓�T1��t,
_+xd��"Ot���	� ܢ�%;.6��"O�0x`��"��A!a��M��52E"Oƽ"�ߴ#���a��)�����"O.Ԫ��ݵK�p9Vb�z�]�W"OfqX&ʣP�bL����WbA��"O�D�w*�%P:���O�Z,Q�"O@��� )O�mH��pF�S�"O�M�AdX��I3�P�H_���6"O0D1Ɠ�}J���g�>hOV���"O����14�XY�2�T�*6|���"O`��ꁻ{D��X Y�:#��H�"O&�I�uԬD12h�<�)A1"O��B\?,����W�I2"OEر"�12�j!��>#��V"Oq�L˹@Z�뵯��:L<A�"O:Ta�G��39j|�c B���ʈd*!�D�q|�+�$���J�.�+�!�?N~a��V��%�����!�d��5y��1AI�(M2ɓ�|~!�d�4��䧓�$��AzW�*�!�d����aXtc�x�hp��CP1!�$L�&�����^29^9ӧ�լ>1!���	-��H㮔y.���wh�%!���
d�(D0�/S)� Y��8R�!�Ѷ>�}z1��
Y�( V�)r�!�,�.�je'J�f�¼��DVV�!�DO&^h��s�O�jP�h31m^6xZ!��1L@��N�I<�x���C�x!�Ď'za�#�N�#CXP��!J!m!��/�J=�Gb��N���#��Ο]l!���|,����;�D�82jɐ@l!�d,�ݩ[!"� d�U7H�|���'wB��*�ޕ��A�8ʥ�'C(0�!��c���#��4��(��'�~X��zL���L#.rpy�'-xxr�2e��A(�o'\�F|�
�'�P@�#�̂q�JDi�)	d"O 1�ˑ�v�J��\��
��"O���nO���a2���s	�q�"O�����_֒eA�� g$*�Xb"Oܠ�
X�c������E~���`"O a1�ڋ0F8q�e]�>d©b"O�-��
�,9���%EU;G^�)G"O �cS�*P��e��M�%�T�"O��S��f;I[c��hm���"O�<�"�Z��U��FA�pÆ�r�"O�l˷+26:Yw+O�\\f5p�"O|u��^�gN\�9�꓉wʵ�%"O:�CD��#������$Ev���e"Ot�Caڀ2>�usq�1);����"O�)E@��JC����p��8�"O08J È��pPU���R�5T"O�M:IG�b?2�:a�]�f����"O�1s���W,��U�
-�H��3"O.LP��%XC�\y�IY� �M�"O6@�g%�Y�jܨ�����D��"OdyZDe� |����/�xI:,P�"O�$�����
���Α#���X�"Oz��@��î���2V�2 �&"O�	�#� Z6"ǋ��I~|�ѓ"O� N��>'�=`Ԭ�Yz��z�"O��b�mF I����TA>~u�@95"O�`�WCW���xtIĊ���"Ol+w�ˤA4}�Gԟ]�~���"O�ꖩ~i��#Bgkq8�0�"O�Y9���H�V���P�@`
P�U"O����J�_ � X�Ꞙ2T���c"O�8�(�NZج��,̽��pu"O���,)z�.�@��X9:� A��"O�ܨQ`њ+0x)�r�[�D��exA"Ot��`N�T69���2*�"Obp"�oH @�AiCmC�h���[�"Op�h��'YW.�k�k���Q"Oz\1cM��f�V��1@�?���7"O�����|�`4��!�8�"O���D僧#��mi�/B+ֺHҒ"O��9�(�q��M�/�6I+~M!�"Op�(B$٣����Aώ��z��"Ol q6��9<tMb%o�!r&��"O��1i��$X�I�YYh��"O�p	T�\�t���&ʴ\eV���"O�OGZ=�h	��4THP��"O�7 G�b��IKw�X#<hM� "O$A����#,@�xa璯^8<p(�"O0�4��9|d|E
�"M��35"O^��Q��x)Ԧ�	����"Oܱ�!�G����rfͨm�T��!"O�I9�'�2��R%�#.���p"O���6kL�R���p*he��"O�<KaD�S3��ꄠ��m���:�"O��C#�A�ne��ؖ�$�{�"O�T�!�7r�>��/۷j���"O���S�Z�&KBE�B`P�!"OJ���G�^lX��ڹ��a��"Oz�Ca�׷�DA��q�@�g"O��UDS=�ju�F�o�"�d"OԴ�W퇤6�N|Hҍ./����"Oz����Z;[F� �q�����"OΡ"f��$� �96���&|5"O�$�eA+Q�J��B��ٲ�"OҜ��EE�m@��mJ���)HB"OP��"!�5:��M�Uk��%���"On�&�%���s��3/`lEh�"Oh�
�Ry!��JY�zD�Y S"O��I!g��B�0�	G$���� "OT��o��$���iP��[#0���"O�ɋ��?+nNTʄ�
�	1f"O��0�0/X��z�E�{�Dkf"O3E�ۅ �4ӧ�Y�%�x���"O��0����R ����.�v"O�1�fӐ|���U��L8XJ�"Oz�	�U0i�e[�İ_ї"O�!؅���lM�pA�� 2}�B"Ol�Y�M4M��Pf�1]L!#Q"O.|��K*n��`[�6"�\��"OB]PO��R�n5#��,w���"O�(	��X��p���F��5�$���"O �:��V�l�9:wkJ.h�.�8c"Otu�q�Q60{Z��#�7vrH�""OL[eO�x�2������]h8m�u"Olh1�&]$��t��L�q\b���"On-� ���� �A�K�5f�I�"O̐*�-��dp:Q��?\�@��'?�DG7Dv]bUM�R���C���%R!�� ��f�B�^��rm�?TE��"2"O��Ԁ�	U��ƍ�*o9�I��"O��!c�F��dx�+Z�����"O� ���8� �t��j�R\�t"O���i8T4�aÏ�l֚��"O%8�&h�H�
T@4��4p�"Ov(@�kG� ��Mkq�>V����V"O���V�T�XD�B��˟a����"O�pKrJ��k���(D����y���;��"��T�B�L�� ��y�6Z�Eqs��=֮�B#f\'�y�-W��]����DlQR�U��y��X�j1>�[V��4.�Qq`:�y�C��Đ,R�#��{������y�P�Ix�(�"�R���B�yN5��ʓ�M�|ָ(	Sj�y��Q:R���u���s��A�b�L��y"ғ`��x���V�W�4d�&	Ƙ�yr �� �6�:i�"O�$��ˌ�ybn�Nv�� � �K���ZuC�?�yB��*`��=�vi� G��ɨq��yRi�6F%��
�ǅ�B��L����yR�ۀ)XL*�L�A��1Y�iѩ�y2 ��(���	T1Ì�q�N��yb�+��- �Iw��8��һ�y�C�[��ɳE�Hk/\,�v��y�l?nNĺw(*^�9�RD�-�y��)Ť\�'MGD�`���^4�y�bV�Vv\h�����D���k_1�yR.��[��,�B	D�\r�T��yrf�7`G�q��`;
x&HH��I��yB��$���i3���*��������yr+���ˆ*+^�s7�P��y� �[䡓t̗���m���B��y�膮�0���J�C<v�Ӑ�_��y��?>~��GA.5;>�@��y��T*�N�(�fЧ43,iY`���y��r�Uh�!�DL)e<�y�AI!s!\ jrE�|�L[Q��/�y���\Q̘`O��AH�� ̖�y��6O�h��⭅�Mp@-�"JR��yJ�(x%�ys�J6V/H��(ҕ�yҠ�=]��)�@*�;}ݨ���E֯�y��[�$+����x��h�϶�y��>�������6#p�q�W�T��yR�ƫ+c����^�{��#��G��y����z'4�� bK�U���qL�y"`�N��RA�J\h@�Q=�y�����(���^����_�y���_�L�w��"��"��y≔�3���Q��M8��	��y2�ќ>������5j�m��#�y�#��;D����W�=X��)�9�y�MS�1���,�/�a�n���y�J[�l�f�砏?)'�MY�`���y��G�� �$ا(rV�ӥ�׊�yb���&m�$ZA�\� �Iه���y��X�ع� U6!�c���y�L�� �˂�,�u�N��y���#�\����eGlX����:�y2A��Nꓨ�d:Z�Z��@��y2�[�}��%��*�0]����eڹ�y���<-��2fnZ�Ud>Ei�����y����p�ک+&�N�xTXQ �-'�y
� ���%��	B��
#.�q{1�7"O��#a 
F��bb�'6z�x[G"O��2�Ϣ%�`��a�h~H��"O�0s��M�b@+� %"}�<�"O�X@!.U>Du���f��b�b�"O.8q�E�h&@�$ωzY6�%"O�L#���\v\��� L�T��"O�I���Ѹ=�x�*��[e@Q�a"O X秇 hd�$�&���0`�}Â"O�H��D�5"~�IB������"O�ڢ,�ms聱2�L�u���3"O��s`n�N(V�j���-j\�w"O}X��moj��D�O�Kp�"O�@r���
'mĔ+P��v=H�� "O�Uxr����٥�D}D��*r"O�d���ŻB�NM(j�h�"OƘ� d�>c�bx[�T$���'"O��(U�
<WYHDx�M�  �8W"O�3J���8`�i�y.Pp"O��Icd�k��	Pf��(T�|飥"O~��핃K�p=�Q
�&,�B�t"OV �V�Þ}J��IP�N���U"O*���\ Y���#e��y��J�"O2�9���#Va�}�I1s��"O~�(1M�*U:0�5�$�
�E"O�2���"s�R�:�j��܉(�"O��A$](Fx�T��c�k�����"O���t�@
j��
dɇ1b�Yh�"O\!`��R/J���)�.�"m����"O��T��p��1m
 ����2"O��I��B�ᶽ�lC��Ecf"O�xC-Os�fêD�4�Qˆ"OR)Q�gM��HQ:��\z~Ř�"O<���+`<^�	2�G�A� �"O�yeH����٩D��v��j "O)hdB[2�J=P$����6�JV"O�A��[-*f�@��9.� Ʌ"OZ�D�;t��\[���$�B���"O�(YuaЦ;�p�ȏ�g�zMڤ"O@���շ]]:m�R烂Q����"O��sF�g��0KF]-�ͺw"O�,����T1'�	��"O�qJRaPoc`4��΄��D��"OL�8u��]���C�	�}��\P�"O4�#b�5Y�lp�Ē�Z�t��3"O*9� c[)>0�ãM	|���"O�Mq �:e��WMK,z_� ��"O�8���	�=2&�I\�
T"�"O�9���J�7�P��AkD-P3���"OƐ�e��'O�4Q�H�?G1 �g"Ol�g��!`T�1�C\�@�'"Ox��C�*.��s'R�1�8(�"O�{Ќ٦LpB�[� ʬ��T�u"O�A�QM��hP"�-X����"O�=3`/X�m�^X����"�A�"O ������aEG�1��E�"O�0�v��d?.̉sg
�=x�X�"O�[��
�"e�&�s�(�"O�iyG'0\J�]���A"Ox��C�&nS�K6�#up���"O�����j���s���b|�x�"O���D��-[�Hh�˚�pH���"O4乢H��O{0�T��F:��"Oz`�b�	6aYP��Ӯ8�Ep�"O� �����n�x��+^�x�`"O�}���ws�m�F��+g`XM�P"O��(w�������S!*R}J�"O֌z6��'3>��k�/�7F�$a7"O�M)EI�\�j`�vDF�Iނ���"OBL���t���x�<�f$� "O*�i689[�(�!q����p"O�Y�%o\쌲5���;��1{ "O
#��K����K�i�ܕ��"O�ڄ��3�q��f�?D#�90#"O�y��'i�$@a�c[�o�5��"O.M�Я 	Jj���p"�
�*D�w"Ov���ӛ'��$�� VQ���2"O�Z��[�R�l�Q�7s�i�R"O*�Y/��̝S�8��qD"O�]20O&9�DM�uc�-R��k�"O���B�E$�H����/?�1�b"O�Q��RIBH;"�B�5�ճ�"O���+��2a� ���Գ9��ܑ�"O<�;�����s�\��F��"O��)AHǕ1r`�8�M�'Px mB�"O��J#E�][թ�-�'m���%"O��ҁع >�����kN")��"O~���j�>\�㫄�<Ne�7"OLHZ�Cy��@��GkC.��Q"O����G)4t�a��B-`�"O4�@�Qau&�@g�^���ʢ"O�d�FnȲ!G`S��B���a�"O��"�g�hHF���B�.(p�"O2X���)S��pq��Ԇ|��D��"Ol�3q�k�d�.N#U��h��"Od@���3{z<�sa�I,<�Vl�%"O:���M�x����W+Ιi�p�yS"Op�;V�P=*�<T6K�#BK���"O��a#��:e�,b���+����q"O�E�� �Gz��ҵP+���U"OP5�+ֲw��3!ݣX��m�"O�aIA���f���(�E^�:tP"O�Ts��Q�"Dv�u�&+~��a"Od�i�bɺ��ҷ���Π:"O�8*aJ�:}ڈ��n74<���0"O�a�bɌ9o/M���kW�=2U"O`1 ��!A���S��$� ��"O�a5�̒9�*p��'P�m3�!�C"O���̛�vM)��_�x+���"OH���,2C.�{G;����b"OHd� Ȳ&������Z�у�"O��k@G"��i��� ����"O���$���� ��GI�\�rmZ�"O�!
��A�d���q��[�"O�Mst�;s�TP��D��,���"O��S%C^/24���^�z1��"O�dbU�P-���j0G��af"O���!�[?T��2�(C�T�x��"Oz����6_��"AF�N���C�"O�Hi�O�A�c��
PM�d�a"O�Yp�
����(��[L?��a�"O�d��ᔙ��5"�m��_�-��"O���c%5��Y6��*e(�	"OJ(@&��(����1�Ŵk����"OH(+�k��ʐ�	���}��qH�"O��s�a��J�)2K��@2��p'"O� f/	�9����J�	:.rm	2"O�� 7�C
oKHЈ�A����"O� ��2���"*�ȉtM�!g�@��w"O�dȂl��f��ӟ^���Ae"O�mX���.��Uk�e\�Ht�P�"Ozթ�i��"�$� 
�Ҥ`�"O���(��k�r�b�早[؜=Y�*O4��4�I-+j*�S�RD��*�'�E����E�EjӃ�+�<��'�*Ƭ����B�KrސT��'��ҕ�^,.����OҲdU��'~�]�s瞉9D���ٶTB=��'�n��팬l�����f�&�>���'f=��s�,�p�戄=!j���'�����W-0�e�"g�^ɎQ�'�rs��!�V���׌W(�1
�'jrm{��S'�*��Y�N�Y�'�52�L��X�p���*Y��}��'6�}3�mJ�V/�Y�U�O@���'��-@)��5�V����J�&���'��U�q��!�|=�CfMpT�+�'��Q�E�D4���MY�X�D��
�'N)��G��j�����S�~�Y
�'y�]:4(��N��)�6���Qφ�
�'�dʲ�Z9*�]J��9��	�'���E	�X�~��!��-+NH�'��wf�U���rCD�V�`]��'1`A�B"��n�<�{&�UeJ���'kTղ0i+�މ�����[�p�x�'7��3���u <X"g��!I��
�'����+��Ed�,��l�:��YJ�'�Zt��N*DP�[7�A�	nn��	�'�&ă�%�g��m�`��0ș�'�����@�a�f���~Ѥ��'����d�4�z�q��N�s��b�'����u�0	�|�@� h��`�'{ DZF	�N{x�7iF	����	�'���W�L�r&ӆ�5cDe��'z��1�l��qʰ��DH..����'��-�&o2C*�U����*��Hi�'Fh�m�
x�\hd�Ϫ���0�"O�X��&b�\ �ȑ=:�v�s"O���F+"���1jT�$V�:"O�ic�JQ�k�Z��q��;��L�"O6,�����<�f ��g͌K��`��'3yi�
�_L� 33 �,`��'�*�3��3w��y V'S�k���'V�;4�ۃIF{�*ưcD<�B�'�n���ٔ#0R�"PJ�'M�$�:�'`�8#!�Ո.�d��̯-z@��'��<2ЮA.���bD��*���h�'2�H��,+*@�{e���ԉ�' ���>nD���ɵAF�
�'c��+��K5��
%<���
�'/����K�ޑC�����1�'�pܻ�_�!Č�)AD�`v��
�'-��� ��7I�rDK�J���'����҂F%�0̚!=yʡK�'7���&n��Y0����Ϲ%tjD��'�ȤZ�`	�iY����p70 �'㞐@��,B���ޔv�D�#�'�D��f�=15��X��3S���'�(�1� =4���G%D:|@��'�*� S�D:B��)i\�.�`�'�h� �+dED��s��4S~���'�RI��CI�.�V��Ɖ����x��� ��0�M&�� �
�'��"O�<��EW�qq�qqc�G� ��Y9C"O�k�*H�I��+A�6�Ae"O	�r�ě*�,���3	� H�s"O��s H#��2���{�½H����,AS�LN��iũzl>��%�M"�dJ�GA#g�qO0����SL�A����8�F�s2�=~ȅB�O<�+�������bpO�.7�������̴9�]ڢ�x.��$h��g��p���P1&˼�)�(�+q\i���.-�H�r@J��b�`<�"a�<)����t����MS���)Ǻg,p��%}HcǤ!Ȱ�ʱ�'L�O£}���$ΆP�eE�pHƝHP�T����Ğ٦�(�4�Me���)8�q�LT;%����$#�w?�*W:g��f�'C�)�L<��/�"m7�]S�
C�iV��2��G.,�4�Sݴ]���	�i��f��e�Ţ��O�����b��w"����Ȟ�i�n lZ�z��,��'X�[¾ �2��;6xȜ`�d�,�>��%L�kl��j*�h`坘F8��:�ቯ �MC��?i����O,>7��?+x�2�ᖈ
Ұ�$�W#
����㟴$��G~R�U��ʨr���_: ��L��(O¨l����j�4�P�$�48�
q��]B��]�pr4�:�M#�|���x�g_	N��f�J_�d��NE�����4`�RĨb�Դ4��I.�OxQ�A��=x�X%R͌�\E4���"ۍ/t�}����|�%�],�ݐ��Y���*b�n6ܕ��4��j�<`�LE��(�!-:�`�DQ��g*�O��Oe�r�$W�p"�*ؐX�nA�2�")sjS����hO?�ĉ�wܒ��Eӓ"g�U�Á�(S�����4K��Ɣ|�O���W�x��	�sܬ@3'f�w�Q &H�L
���Fʊtx�T���lr.6��^�����/�3��5��'C�<�R�p�	�l�:$H�(]�o�"?i���
{ހ�ׁ]/ ��xE��𐪥 -��{AB�1Q#RO�h�伱/Q'#EXt9(O�����'_����5���ɵ���{0LH�H?�7-�Onʓ�?�(Oxb?u+ ��r���އxN$�ӥ:D�TK�4t��@�!N���zRa����ٴ9�6T���׻�M����ħA�5Z�j�MDD cGS;����=��X�����(ܲb�P�A1�O�ڱ�vKz>Ţ3a�4�0�;Q@ߦR���k4ғy¤E���R�b�M)�ɟ1Qr($��,V�;3>$6�5,��a
"��Uè��R����5�+4U�H�.��t�	ܟljٴ�?����yBj��:����N�e���f(_ҟ�?�|�K<�F����ఁހZ�pm�4��g8�	ݴ=C�6�i
xu
wĔ�I2��R���P�@j�'�R�ۢ�v���<�'�zL<���uz�u
V�M�Sg~�ڴ��;��)�!_�pZ�y'�3yd�x 2�Z�'���8����F�9= ���s�^�$6͑�f����I�A��b4fE� 3S��"��åU*����hi�E�3�d˂,@1u9���7�i'x����Z���<%?q��M�&�;E"yXW�L�i�
�-s�<�GU->$�MR��^�)��ӓ.�y?1I>�p�i�T#}*[w���� �ց`�a+D��>�~5���(��9lO��9`�  �   ;   Ĵ���	��ZP�viė:&���3��H��R�
O�ظ2�x�I[#�x3۴|f�v�J=|L��gJ�'��l� j'�6-�轢ٴ.q�$0��\�I�F�p�� I@��4��X����f$?�!�r#<) �d��&�R�~��� p�<
'��`�^�xQ��A�Μ��'?����6}6-L}�D��$�A����36�̣ln*�c�CN^y�C�ODcs�ʎ��9O4�y 
�/��cEI�6\��L���X����b�8��D�`�葰1����'H$�n��$iq��%F��P���q�'�dS�	�lu�'�����K �R�	�7
�j�h�'B,FxBDH�'I���vjƓ4�T����ܥ/I���O5Ku"<)pI�>C䆚�J�PMV�M���/�H��OT�R������'s<!��m:����)�*rY�8i۴;WH"<	s5�Fa�*�Ɏ(75Z� +|�;qh�Z�>��#<1� ?� �B����P�¦.x2�Kc��Yy2��~�'���?I��ؗ	h���'��MY|[Sj�?t"<�e8�2����н)����B�R�]v���s�C1O<� ��$����~B���p�� 7|��ukƐ���lT"#<�m5�k(:�R�^6V��-AfՈs��x��o��X�K���i��mGDq�����|y�@�3z���*��$�B�<a��"T��P�<�2k�3Uo�O�2��>R��#%
�f�>I�s\�l���I�-C��Qe�:2z���P�:Y�I�"7D���'K
   �a�N>�,OrE�h��y�ޅ"#ŗD���8c��O
���O��O�<A�iX|����'p��12���P(� z�p<p#�'�~6!�ɫ����Ol�D�O����C?[��}���#�D]���_�7�!?u�y�n��7���)y�J�1_`@2��j4�e�qK`�0�	�<�IܟH�	� �ґ��)i�1y�i٫b�� �/ֶ�?��?!$�i�ЈӞO!��r��O8!%FMy�jDbWHLD�ސr�J!�D�O^�4�b`��k{�|�N����-hm]@�Vz�<P	1)��I@��Ty�O���'o�k�$)Wbԁ��	"{A2M�G�A6T���'�8�MK&�۔�?���?-��P�B�@�
��@����8�ٳǟ�p	�O�$1�)҆,
	���i���[~�R��m�Ρ ���A_���*O�	���?�7"���H����    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   �	  �  '  �  
'  �.  B5  �;  �A  H  aN  �T  �Z  >a  �g  �m  t  Iz  �   `� u�	����Zv)C�'ll\�0Dz+⟈mDԤ�57���DB�������$)�9�R��<5G D�Eg�  !Xm�@�߶>���VƐ=-�I��~)�U2�'Wꊠ���(I��A��{�>��`��H�t)�#GJ��x�R�<2�¶^5���Q���������,���0c�Ш�aA�H���EbN�R]e�pJ�8Q���5 ���"J�9pX�q�4gn�<����?!���?a�K����_#>�xؐw)M;9
�����?�1�i�*7��<���hܘ�'�?��v���aD��[2�%��_c��X����?S��Ɉ*48!�	�fl�l�p��A7�̠$�.r�F� A(�,q(@����<� d��1q������℅�F�g}4O�㟬���R*-��'��8�Q�B�s%���Pl@hܼ����?9��?���?i��?�)�,�ݾ �j�[4?S0���%C�=m� �d��a �4(���i�����nZ��M���i��fg֌
f	�E��+ZŌ#=!v��s�O������9Ahd "%.��#0�,���[Q���EG�u��� �i��7��ԦY�Ӯ�RdK:*��X@f�z�Px�E�I�lQ\{r�t����P�[�.�s����h���I�Dk�7���޴�z욁�X�E΄��r�ZRːH�𢅮)���5C�����GyӸ�lڶ ��9s��%{Ӳ���D�<(tM�gힲE>�Lˣ.�:yע	=��i+pcϰ{�I�ߴ��/o�L�X�g���Y���� cvO���`�ϒ�d��CĪO3d�܈�iZ�dz��N�`xv�a���AR���'�O��aNIa�+r��R�
���g[��� �f
����شj����O�4�;Ć ���@+"��l$����ވF��i� D��'!�D�h��p1�`�V�#�25�!�O�W� U@�G�0�H�֯��!�$I%Yn\�PJ%M$v�&�O ,m!��JנxXҁZ�,��cl�:=!�$�0@V
�bağ^���yeL24ў r��/�NothP��'u�(y���%���"�X ��-���#�Z $~�ȓY\��CHĨ}�x1� �M�r����=�u�8l�]cco�b,��ȓo�$�D�;��\��?l��d��@���:�遌|w�!g��72��	b�#<E���שrm$<��%�"l�Lp��ږQ�!�$ۢh�n�iUÍG��\��NLA�!���#�QN+���5�F#�!�V�=��M"`�A�\ 8�,��!�d�3H"�B(�_�P�	�`R'�!�dBn&�C�Kg�PR�	C�)`�ɑ2˺��ĉ�s�(ib����0R�y�B	��js!��(&��x�Ņ4���x�悚 !�D� V�����=B�&�CE�	!�$ݘW����I�j��8C��܇/!��.q7��i0痍i���A�����yB��>d��6��O��N��B�y����j�c5��$�O�H���OL���OF�p0��O�˓�y��Z�uÑG͙t����A��0<�BnU��h�	6mz�		��M+���N���В�W���D)}�2�'x6��O���IB�L��xd6R$1X�%�<�4;��O�d�ɉ-��̣#�OhQj��ܓOcZ�QSD�2yx8�qd��*��|J��'�L�	<:�dRQ�I 1x�������!�����O�˓�Γ�y��7���6��(e�M������$�`g�
�{��	S/m�>�2��ڝA��q�q$�K�	%� =ʗ��S.P����%BU6 ���
 6`��K�� ��ٟ�%?a�|����O�����Ul�-� ��k�����	�q����ʣj1��ň^EF�?)���A(|��@пD�hEz@��>X�H�� ���3ʓW�����/�(*f�$�<0���/� �)y�bܲӈ� <��z�\j�̢~m�Y#sL�3�����yZ؋q��cr�$Ӓ�ŌBv����&0���Gݝ.�	��^:E�H�Ɠh,`�#q�&Xk�Qņ�.;-n��G���<��q���]Z�L�p�T>]EZ��D��z<��#p��)��wL$i�ā�}�ֽ���'p�@�"˲Lۀ�	b�"����B����� �ز�R����e˹v⁇ȓ���+0�ʉGR䢑\ ;�,�%�Y�4���� ����N�;Bt�
&�O�l�L��w�@��?�,O���O�����,�\���e�.�.�P��!D��� Y��&����(1���ټA'f<�}5�l�ab ����J��Fd\1pq��!XO(�"��N�/�3�BN ��On1�`�'��u�"}?8����m��2!*�D�O��(h�)���'u��1�D(z�����O�yH�f�aI�!��xq�T�'p��O.���4�?I����9H�b������Ԉ�7n�d`JF	��.g��'���r���t��ɣ�@Ը2���T>U�O�|,�@*�5�m��K@H�O�JWO�(�\�h�֖\w��}J4�U��!��F�R��h�F�e~�鍢�?���h� ���0��88�kR�N�>C�<-�iʷ ��g���,*Pq�����h��d�Ԧ�St��&���4�g#j����<�wS*P��'"�'��I�H&\ӣ��	MӼ Z�a�z�>�d���b=���P~���d
�K�d�O���O��s���0�@1I4@�
$c(,��_$7Vx+�L��1��܊rL�~�UFI���F��,$��p2��$�?�´i��Dp��Y���	�N��8����;*a�����.ٔ'�ў�Gx�)�>R'���U^��`J���$cӞ���Ozqn��(��ꟸ�O��%#�)�-9�6�kF�ܰ6#4�b�ሄ*�6�O*�d�Oʓ��Id>���_���1yÊ��&���'�;���"�Ͱu�Co�@�FrJe�5��+�.8iꁣ�"`#lR-�=r��ˇ����_�+W� ����(O�E�D�E�$�1U�~ĉ�B!j�b�'�6M�O�ʓ�?i,O��'[N�]#iL��Pe9�,G$R�%�l����}R@& 9����ނC��������M�����?YC���y�5F�F��׍ _���� B��y�kҙ���$��5mzy9׈ ��y	�T�P�Aci�!�4��Ù)�yb��~���2�
�;�L�����yR�\�k��ѴǏ��(Qk�I"�yr��(Et��� �={�(0����hO������&!�,PmV�\���Kp ]�8�C�I�
���cAL�v�j��v�گ&�C�I)ee��K��0@`~-Z�� o��B�ɣ>��рh#���7-E�B䉆CVZy�'덡m�,�`�ҵ:�B��;,v20��\9~U�aQ/us���ܬ�"~� �G��t�ڳ���:ǔ��d��yj��
��c�� 2 �c�� �y�b��c/���A� �}�i�A@ۥ�y2G	�&�����jM�
Q�U3��B�yr�ТiF����YkP��#D��0�yR�I�^���XP�_�c&*4������
�|R̀*��B	1Ea��flW��y�%Q���Q���&��0��bF�yb�_��b2���Q�.��e��ybKq�,x�5>�`ti��V��y��Η,D`Cf�$n�n-�%f����>1҉Nm?Q�%�\u��e�)]�ڡ: O�_�<��(�,"�6*�I��X�6ِ&(�C�<��R�#E*a� !�䀐�<y$)�CO�� �K�� �2�+�ov�<)A��;,4�U�Ӝ+B8<c ��r�<�1ǉ� 4E ��A�"�0�Vr�'6�1����>jT���Pe����J�P!����a��F{��rn���!����!*��X:4Xzx�,Λ"�!��t����K��>���t*^�!�$�o#��6��=܊,c��D~�!�ą/.�X�ѥ⏬-�Na0CF��&2dZ��O?�J�"x_$�jĤ�)Wԥ  ��T�<)�m�E��ҖL�Kl���k�M�<	4�VH�8�2��jT�1H�H�G�<���&6Y^Lk�� ly���� �]�<	7�S�|���pEWc�h� �\�<�F͗�%dH��B	}�̸�Uy2l���p>	��p�9����&�^����6!�� ��B�HƲh�:=�-��N$�9""O`1@cH��'K��D�E	�B��1"O�y{gǁ�3�܀��+����(�"O<�c��ҡ<Tu!@M�='��"�'� ��';ƘpP���f�{V�T�}�
�'vt�ڐ��:c�v(���S��)�'a$���G6� �vK�-I?+�%D�z@�Z>�ȍ#%n��O����g1D�T�EC#��I��E؇eq��"6f$D��;�ۻDx8c�	\�����.�D�AG��gZ��T����s�M��ݝ�y���?L&�m��[�'��)I��y�	��V��-���K��B�"�ybMŶQ�YĄ���}؆$��yRV)��ǈJ"y�Y�����y���GG���`��0�~��TeǑ�?��W�����Kr/�0d�"���a�h��o���y�"Z�I%���dC�
 R�)q% ��yb�
�t̠�)��u/��p!���y���
3J2h	�)��v��o�4�y�-Ղg�e2���^���헣�yR����l�O��[K��"�����D؃*��|B��%�:��d�CH,�[ƥ�y�HE1��J�2D���v�ʷ�yb�Xb���qdű7��M��&3�y2�/t�0-�q��4�tm�����yҧ�n�0��B�[� ��H�������>	sdWu?���0`�i��;vtҀOB}�<Iw�F�F�81ƍ�?P��h��z�<�TO�G�ޡ�2�Ć6��E��s�<�cD  ���h��
�T����j�<�r��5����LǔVT�Al�<��h�>P���@�i�n�1��L�'��š���L2R�D�Q㘜A�0�[�o'!�)Nנ��u�W�`Z,"�cҥr!�Ow�d�F�*&xǌ�9$!�$T=Sz�+�8-�����(_:!�D#�������8���zTA��R/!�J"2����� ޲�ˑ�Ͻ�R��'�O?i �PSK��3�h��q���@�H�g�<�nW:DL�	��:3�R�x I�b�<	�ǩe'��G!�8>f~+0�Z�<�VI̸n�������5K����ΌR�<�5 Ҕ!��3AW�8�bl�vʟP�<!T�Sd;p��%FhqRĪ�Qy2N�(�p>�!� �c�:��e%R�>v>�a2ɎQ�<Q'���P��'��s~�ę���L�<���� �§	kn$����L�<��*�Hݰ�� w��R�%$D�X��ł>+D��*��%-|�uB,�O�E��O�9��-Z�Vİ�ȖM��Y=�y�"O�]&�Է|��Hp@4�!c"OV�����A��ʕ�k��؀�"OB�ʢ�<M�A�O01�hPs"O
,�P�X�.�NUCb�z4���D"O�mqe#Y]�d� ��@�iE�DB��	����~27@X0e�ؠ��A�O�\���g�C�<�ǃD�2$IWS/�<Q�"l�g�<A��ןo|92򍐑K��8���}�<���ϦQ=��Q�
$����+�a�<���9̢�iˆ+V!2e$�`�<��oR!Q���'�Ļ>��Y�fEß���j&�S�OI4��Rep�,ЧO�Bc�M�4"OX`�,B�B��<+& (�)u"O� �XG��$��x3n@:a�.q:�"O��`2���ex�J=G|��"Op�rW�L>S�����;4�Р�4"O�hr�n�Q�΍(q*�� x��V�d��M;�Obu 2�ͳ
h~Y��IB��c�"O.pr�Io�z�#���%����Q"O����&	)Wb���&H�H�q�"O� �X�0�썒��[��Y�"O�UM���+͊(��T���Nx��e��"�n
���ZR/ĿW����3H!D�)�%-b%bC���dp��`�#D����⑓��C0�IU��wA>D�q�O�yz��CE�WmB� �?D��{r�6bL��$� �3�F�M=D����Ϛ ]�.,� .�
o��E=ړ
�D����`>�T! 9?Z(Бp���yG+V�I;'#��9�M�l��yBÚ5�|4�E��(]�`��DT��yR �*JB����[3"��Nޒ�y�"g��裌��H g����y�R�d2� jE%�^`r�ܑ�?��l�]������&��"bi��Bu�ޭ?۠�:��'D�l!m;/K<-�bG'[�L���'(D���HO��
ࣧ������*D�p�#��'h���D�BF�1@6�3D���-�d��ɳ.T8*��]��`0D��X�G�$E�(8c�7/r>d���<Y�Sb8���ч9I���ф9 ~���)D�(���-��Qr�9�Z���(D�(�.E.8�2��mQ�xeN��4D�$�2.W�I�,9����H)3o4D�4��j���`H���5Ԅq�g3�Oz�p��O��rԤ56�����JQ�N`x�A"Od�0�����M���_{��ɀ"Od	yV/�NH�a�M���W"O����>1���"`���""O����(!f�Y,1�Q�w
̎�y��Ξq18e(B�����d�&�hO�CD���:�h$�E�{�V���W /��B�	�\>xܪvdN�l&K̅b�V��1"O�����b�*0�0`ȶ&�8Di"O��Q��_���$�P��t"O(P�7EΤ"$9(���L�9�"O��	��0g�$8��5h@�d�'�0������Vk��P���
�2��� h<��x�]�ޅ&�1��C@���ȓ^f�P8e�bD��R�Go	.���QH�)k��L�'<�è$f|��ȓSX��� �X4X�B�x��ZC"��gt��4��4�l�q$dԜ	)J��'�.I�e��@@��68��X��W&���ȓt�Jp`G�:zG�YCc�@�oʝ�ȓP%������+'9����-�P�
E�ȓ=��,�!*F5��4�U�G8m�=��X.�8q�^�%�Z�2�"N	c�<	����}��	8
X��OR>�bJ�5��C� ,0��5l۬ļu�� ?w�*C�	�+XZ����:(�H�'�1Xt�B�	#Plj�j��G�Q0H�B`�ж|�B䉩�D�:�G_�&}ZQ��a�a�hB�cU�E1F��2P:��BV�=�)�j�OD�[Ƃ�4� ��tB��;�@I��'ۂqj2�ӬL�h�B�1�v�(�'�Hl"1�%I�@{���}�J�x��� �Ð�V�f�賓�*Yܪໂ"O� ���6j�F�� F�@L�t"ODL2w���z��p!N�C��%i��'x�R���ӡ��\C�ȇ6~�$L�I�+C�|��<E�	:�I�Aߢ�L�4�^̆ȓYҘy��!�#��؃�R�dԅȓVi��ע�$m�|K���;�&I�ȓ��zC�G�
A&�q��O�q�*��ȓK���΃6���KL,��'�$��W��*r�b���Qe��\��ȓ������S������ۥ�꜄�dC�y	���+��l
3��%򪑄�O\Ea�i`OV�26���i�ȓ�Ф���R�<��Z�+��p���	�m~��ɶR���H;7�Y��@�7M:C�	 v^�� %P"���b���<C�	*+��m�F�פ�����B�\�|B�		�;�T	.p�Ѐw
xdB剷=ex��w���%W��2��V�@�!�$[��=���XT�2`��_�ўаt/)�5�~�xR�e�px[5$W?v�L�ȓ]�PP��{lB�!�M\�uT1��9?Sq�j�E�Fg�
>ε���Nl!�����	�$��&���ȓ�2��%B&��m(�չ\5N-��!�4R#)��C��ř���3=8|T���Jm�"<E��CL8�S3�ZMc&f�rh2"O� Iwb�bT�A���s�!Sb"O���⏿E�u�r��7���E"O�s��4 _��)֋��E�4�t"O�Y�B�%������D�OPp�F�ޠU�����/<�z@!�f���'{��n�,��'z��z���B������� 8#� ѻ,O`���OL�䐠G����;=�2��	'@������!B�D`���L��I�]W��">���F?�TI��+U$ �j2�j�U*ld�eb�rj�%T1r�S��à�(���jD�$�Oc>��pj� �s������V,�<!�hp[�e8;�[�8�H���0��D�j�@%�#�"4��#%兪T�剟8	&\��ԟ0�'c��П4�I�!�<�Մ�4���: �g����ɷu"0\9 �~q `ī`�"�	!��u�O��� DCO=9�(��D�Ν�`�'d*�@L�!|���P�(L,؈ )�eB���x�}�`=&�(����%*p����<Y�����	M~J~*�O�sTAM8 �dQ���jޠ�E"O&E��Ǆ�T5"0Q�*�i��]!����ȟ�`�d�}،�ʹ-�lK��OL���OF��C��(<��d�OL�d�O`�)�O&{`B�k`�C�Ş������Q�1Oem9fiZ|j@F\�*;���O�b���G�Kf��R�D��VQ�5`�[$G萰� ��H].c��&Yt�'x�x�)6,i~��G�.��]zGLZ)-"|e��D��dX�Rz2�'�ў�� sщ��T��)�+c�)�� %���fM�'A;�A��]�S>��I��HO���O�ʓV�8"�8OȲh�� �媀����7y�ڀs���?����?Q���?9�����F�����')��DU�	�N�-���8Aa��*�haGC�
6��&#�H�'D8i�酞A��]!�l�1g=tE ga�A�Qiۇ0����E�@x��q���O��Ñ�'S h�wd�����F�	fE�yzD�'vў�E|�����[�:FJ'oH�o<R�ȓKyL��dJԒV�����Q�T2Bx�'��6M�O2�\�9��N��i���4�\JЊ����_&��B�_-�?a@���?q��?1Q�2ۦ0��U�gH8��|�Cn^�w$T����G�x��1G�[H�')bH���Rf����Y�C��8�*tH�	YoS�M8 �	�7�4���ORc>��F��d��ط�̝US�(�b&�<�[��!a�ϔ}yx����l&q��I��d�-c�F�C��1xI��	�H9[��O�4ِ�9���?�	�K��v=R-��YvJ�$�C��&��c�p�uy#�;�PC�I?I�8��p��l`�E$	�S��B�)� (������huRb
�z0��B"OȌB���B��юV�0���
�"O���m��T�A-�)�LtR �Q�O^�}��W��p�b
n�13��+�䑆ȓHg�%�F�X�-6N���7�
@�ȓc�n�A!�N�1D�Yۡ��N�F��ȓ`y��P�LyI6i`ceٱeT��ȓ!��kPck�X���/)Ϫ��ȓo.R���:p��+%l�6.p���&>����$ۊe��	I��3ΰmƦ��C��G�=��*��L�x0��1|�fC�	<�q���ɻ4��ك�6YbC��'e�L�ȀGH&3Ȫ�(���u�VC�I�7�ȳ�A�A�0��g����	Z�P�'N28�N�
f�@�n@�r��U��i�'n�d��'w��'��h�u���~?�iK ���a��7-��uw�E:G��pW-_�8�����m��O����fekA��-�p��)I0��*���E����0���(6��  ���On�d-擔6��[Hsj�󷥍�PI��0?�p�-���R	��
.ȵ�V�U@x�H)O��J  ��m�-��N�?a����^���I�����|�'������� ������JMm��	U�'�ў����ʄn��z��X�?�l�!�
:�Ɍ>�Oxb?�1��6��	{c�@4xЊ7M;?��OԂǒ>��y�M�x�0T�T�ؔY��$�$��Lk��8�O���@�,}�� 񩄒N583-�I���g�ER�B(K���'��>牎^D@��6��?Rɒ�[$DT,����U�+}�h+}�������i�h�@
�m��\1^�a�F:Dh�aK$��ɍr�Т� c֤j��q���J҇�]�?Q!��S��@��r3�_��,���L�%���p	TⓂ��:$��`��?5�"���CV��r`����XSv����~�$	���|�fL�Z���?��n?'�)S��JV�͑�a�7M�d�'��H��O��B��i�8�z���պX�r�yrc�_�mV[?t�MS~ʟ��T������8팯[c�1�ԡ�>k2ie؟�أ���]�������,P��5D�4��>`����Ĉ)���e�4ғ��'�"�'�Paɳg�~�ap��X)/�	��Ʊ>�K>1��T?��\M/�4Ys��/ZHX�
�M�y"b"F(�(Q��|{��Yw����y��Q��Ь1b�������V�yR��0
����!���Zgm^��y����X�v�֕��`6�U��y��?dZxU�0JM��Ys0���y�O�!ҹ�w�>J��5�FN��y�Bߙ�J�[fF0,�,bvl��y2�� �FAqf��?W&^�yBM9�y��fL ��g�RI��P�fA��y�n�r`���XEN���!�U��yB!��$�����-g����f؝�y�-�:��0�&��2	�6iy�����'n�}¦l�-q:����m�!r���"b֎��7a����̀>њ��͎�X��@�
��%�4��Q,�?�48��b*�8��Qˍ$,�jH�0ʁ�!0N12L�!?���b�L>`���h"�7gp����
'*���fiɓ϶���6$^lq�1�'T�j�O��&Ď��*p�c£
�ؘa�IBx�X� Ϥn��Y`�ƥC�Ĉ�'.D����a��L����FR�ZLK��*D��8�ˌgY��2A��(�l���&D�0HrKM,>� �����Ufh�A:D���-�=NZ���Al8}"�6D��A6���zV��x��A5D�X�a�'7#��;Gb 6���HT�1D�T��,˕1�VP�H�U�r��u�-D��{���Q"��J��c.Bգwb*D�`XDA�)i@�r�CU�HWڰЫ&D�8�#-�,qF,���2 c��d�#D�P���ѮVxz��Q.(d�v��+#D�� �d���K�?�r��O�9���"O�1*�c��z�����i���e"O�0q�/��Haܵ�W"z,Y�"O���ōT|�����v,�1{#"OV�K��.ঔ�vA�;����"O`HЊP�\���h@o�!o�&��"O��i�˲8�EKȗ'���g"OT����>Q�M���M8p�d�y'"O �P1��� *���.,-:x1C"O����D�n�x @��Q"O�(��$�1}-N0DŒ�N�aQ"OL�`b�Q�q���S:Z-���U"O�(��\"��� GŮ/ (�"Ox(P��I�2�QO�&2�T� "OЌ�E,R+ e�M�;�*�"O��з=l�3�^�v�Y1�"O:� ���0��V�]-O�0�h�"O,�)�j]�s>a��	33�"O��Ħ�ck"M�'X�c͎h�s"O>�S0-N|>����׆�b�"Ov�h5��0s�����0�J��A"O��9�b"+UJa�����a"O~����&��!���A����"O���3!}Luk�	̀��]C�"OHa�@Í�%]�պ��\�m7T��"O�Y�if~�u�'�V��"O.AS
��O+(� f╖��ڑ"O�E�*讁(C�W$+O�"O���P�ӧh����HQ�(�c"O4͘�JW>�<�k��/�x�"O�Q���k�8hKed�lG���U"O��B���NV �A�BJ�J��ܑ�"Op��`c�$����ʠS���*a"O`s�V�p�T���W?{����S"O`���# ���h"�t���"O2��U�R���0c�� D����4"O�ѱ��8&^`�"��>m"�ݨ�"Oz��cOC�*�$ɣR�V�IT+w"O�=�@CY8@��O
�)���a"O�l ���[�(Ĺa㛃V�z�#"On}�A�C�R��$A�4�T"OX�VF��)6��86bׁ_p�yC"O����%�GY{��X�eD`M�5"OzH1�ㅅ��A�" P�q�-Q"Op(s��2;j4��W,��G��K�"O]rRo� ^j��&��CӾy�"O�Pq�b�&E��@
!'}
"Opa����{��8�&k��^4� 8�"O�y2Vㄺ���E�?��J�"O�ev�_�d[49:���dĳ0"OV���D	)C���eش&�x��"O"�3� T�/V�C�ot ��"Od@c�I'C�	LY`��"O�D�$@B��y�e�D�ȫ�"OO�դH� ն��gA��y�Hʐ%������C���Lkf$��y2F̛X5�)1g۲|��ı�$�y�!�*n�0�Q�b�+�|�a.�+�y$��H�~YA��n\��sH��y��/}Π�Hs��b=�t"$ۚ�yrl�.�dD�QIюU5lK�+A��yR�7
�h�b���L�,��'%��y�Ws�~��&L����7����ybH�W�N�2��_B������y
� ��P2 �Yk�%���ƈt�~���"Oލ���'Y�Bq�2�¡Q#���"ON��	ڵ7��Q��Fdaː"O|�3l˰A��PS�ζ:i�)"OVѪ5��%,iR%q�nT�tc���u"O���Z!(�� p�+�%��)�"ON�R�e��jg�X�
��V�`l{�"Oxq�J�g�@���5��Eڐ"O�$��>���ףĭ$�b�H7"O��* MF�G�u�5h�o����C"O���#�P~ ,�(4�ͮ�HT�"O�T����-��,�t��O��mE"OZ����ւU1D嫒cU�t�$�s"O^����1$��y��A~�U�"O���g�A���{��
�{F��"O�������H3a��"CV000"O�U2�^�>�B�Ceꑑ\2�x#"O����P?lq:5��O6��"O,�����(�J�RL�5Z/�X��"O�hR󀑴C\~,�jߪk���@"O�չ�f� Bh`��)��7�LԘf"OvK��&-v�:���9�B�8�"O��'��OU\��ՏFK�483�"OpL"��)+$T�z��:@��z%"O:���$B1eAZ��6*�p�<�[�"O�T�t��|t`4I1�Ƚqˮۂ"O�\Z�\9CA�YHUO,Wa
%3�"O����ރXb �@.�(#�(�"O����GZ�v�X�C�Q-Ӛ )a"O��O1�>Pr���W��)"O&ؚ�ƋZ������3|�p���"Ol�A�k՜W��G�)*��â"O�a���rWT@T�&�v%�v"Ov,���a��D�o4!A"O�Ɂ����Qj�
wރ>C�-��"O8�)g��*\%�
@]:���"O���"NF�gj88��Z�k�ȩ�"O��BC���a��8@��* ���f"O����n�n��'��Z����"O��!��h�T1�G��W�д �"O�l���B�Y�<-zD;��	C�"Ovy�B�X6&	�5��#�P���"Ot�#��U��� x�̯F�-�v"O�`���G�.!0@��8'~�k�"O��n'��tcl�)s��q!c"O�h������R��ǻBB*��3"O�D��Eՙ;L�X{egՉ)4x��"O���'��Z�2�[�^�=��Cb"O�$qC->A�5�C�(F��p�"O�����2*H��$�K6u�t�K�"O�M��EQ�q�5�2ۜl(�*O��'邉=C����b�W\+
�'Dv�r�E���gI�!xF��'�vu�q�ջ�.�" !�����'�F=j�M�-W�Q���ދh��j�'�����=u=�q�ʼft���'��% EQ�ڍ��mޛV��Y�'�����@�_�fe	��P3TZ�-��'˖C�
�O,���V��B��C
�'uR�ӂ��'&��aN'�r����01펩Z���h�Ϝ[
�'!^�ze*�.
\�BqnZ�\n�@
�'��t� t��|����&o�Y	�'HD��V��?fLm9S��F���� @�`�])^2�e�d�c�"O�ȑ%�3�L��PТy�F��"O�<�t�L�a�pdM�|-:H�"Oz$�bO���C���<��B"O��p&�=��RTEʓy�T�q"Of<�b↑4�"���M]���	S�"O(-1��3$Xm���q˂��"O�d�-���3�ǴJT>Hh�"O������3*��b�l�wD:�`�"O���4Hú0��I!�K7�[�"O܌#0�Ӓ�(P�@j݊=�p4:�"O� �b��`>T�J-8@���"O��9e��5�Af/N�W*0q��"Ol!�CM�d�1�/	�D��s"O�1���V�AmF,���()�x���"OnU��)���i�(��M�"��"OH�C)�-Q�N�'R�<I�"O�%�W�� 0H��r�&�\�"ODIٔK�m0��Ci�<Y�v��"O��V���	�vD�3�ˢ9���p"O�t ���+}�R�S�~�,��a"O8�Q�˥@�2a٦�FH�\���"O�8
��$*{2s!�^1d�h�H�"O��y$��
3��*���/{`]p"O�+�
SUt��m�T"O�!v)V�T��y�3�[0-_* �f"Od��7���P6>0��Ù�;��)A�"O��Q�X�(ȅ��	YΜ�:�"O8x�bW [����@-��,�C"O�m�u`�+t�@�MN�fL"ZR"Od�wM�-ilts���X7J�"O�p����n��ِ5mT��H�A"O\�j�BU5��yUꎗ8�h�"O��Xu`�7 �|R��4m�ѩ"O�@{V�U�"��"Ā���Ѷ"O�!6mַ��Q��%�<��"OP(��_g8�(��b:�d�C"OBm���R=w%���1BE*z2:TS�"Op�aC&P�>�"�hG���x�+�"O���0��2"(��2W���.pPI�Q"O��R�� W��q�S���h_d��"O�p"w
,{�6	��ϯ,Zp�:d"OT4*���Z�ֱ0�%�}Qp=��"Od�(�+�M_ �q$F�>���c"O8ݩ� �%q(W-I���q����yr̦V�U�Lď.���k�G�h�<��P��j=R�.�C4�x��.�i�<y�	Ȓ�\9ȥG��AP�Hq�<	u��*rK��p�`ƪӒxy�-�o�<��R����'�V�h(��ۂ��n�<y1`�g@-�B�<�L ���h�<ё���3U�@��J+���t�f�<	�H(p����X�<� �1&��y�<�'�2
L `�ڢTa)���a�<��JX�����ݜ*I�"�_�<�J�li��pbAN��QdI_�<�#.sZ�a�⠘���XQ�Q[ܓy�Ԭ�ЬE8�����'�,�%��i�삌i�P1%��6x0��:$'/D�@�b�:2j�ܑ�ئZ�Z}Q�!D��`�o�Tx�a�G����*O�l�F�O�{�YPB�� �x}��"O.�q `�0ā�,@���2"O����G��С% مq��`""O���t+�v������| �*���y
� 0�@fH� Le1�Ŝt�B��t"Op��%�d�"���%֭tߠ:"O��X�ǔ��h����#!�I��"O��pB�� E�ڔcD������E"OX=��M��/ڶ���*�	J�q2"O0-(u���R"��8
��2���Q�"O8���M�g�.��ЃZ��) s"O�p�'���?���b�CP7la�I�!"O�}C���+,I��HJ�xE<}��"O����c��|;�Ua�����"O*@��oX�L��\�.�&l�ԍ9"O�y� iƘpQ\�"� 2T��=+�"O�yzF!�	G�t$�W�� ����"O�iچ��|�\�Y�BJ�r��Ȱ"O ٗ �%m#�8�@C/5l�L�X�<1��R*u�豃޸^>N���c�\�<2LR�G4���
�9�4M�t��`�<צ�!?�\i�"� �<�qS�
G�<iǠ�_6�5,���2���c� B�	�%X�eҷ��;_� bu�E?B�d�p ���4.�b�X<'0PB�ɸT�
@:r�˦q�L���,.gA�C�	�o%HX��}�p(@�tŘr�'*l�0glI:Y�1Rc��OުT�'G��#UL°ilf ��JNL!X�'�<�K��aϖ)�5�ȸG��9[	�'G0���&zdd��M;L4�a�'VF��Deڴvqx���H,B�T4��'�"�)uG�� ���cW0>!8�'�-c�/�k.e룁�"����'\���Ǉ�5c7�@�F֞XR�*�'��8z��X[tU�h�1:���'�@�G�?9(�W�ܜ7�!	�'>���V���r�6qj���1���8�'�X�aR般Q�Z��рNP萫�'�\��E;ޖr'�9ox�0��'{<y�e&��T Y�HW�d�ʼ 	�'�N�cc�m����sǎ�nV�Y�'���a`��J�����Yz���'rT]��&X<����	�O$��	�'�z���L�}},��-_ L�Q��'���%��z��a����B)�|��'��K�E�l�`5�`%)�B���'G^xU`;�l3&^2w���q�'E�D�"�$CH���,m��'^.-h$cW�^�~)��d�4A�0��'Z��D�4�� }r���
�'A�8��h��J��f��o�Ȩb
�'��r�N^�)�`X�AB{�(��'B�Y��'�-u�8	��쇷p�^���'��t(�hI�65
�������
�'֪�r^� j��S�l�����'(��;��D���]x��1^��}y�'��t�d,��A��AcF�\�����'ͦ}��
Ì���!c�=Pzyc�'O8��ߛaU~��E犢is��'�|1SM+-K���䣊�DA���ȓv��z���1yǰ��`�B<h�lЇ�� dkTY3p�`L1N�Af����a;Q�БTH1�u�͊s�D��s�9�6I��Ĳr@�-C�6���W�����À-;�j)*�X&'�T ��E�re�p, 5'a��I�#j@���^+l�3`Q��-a�.��{��͆�S�? �D����SH��Г�T'A�|��"ODt�m����h����\���b"O�QQ�aוe�ư�˞&~��s�"O�h�1�No�p,X�#�
#�tX�"O.���h@^L5xc�.=���*`"O�IBFb�4DL�yv���tY�5"O�ly��/��Ԩ��4��"O���W.9b�2��L�=�D��b"O i��b�#' �1.@�e��-�"Oހ�@��J|z�K'l�gN����"OZ!q�.V4;�<�"cbTa�F���"O��ѱ@�8$��,�GE�X��m�g"O m�6jI<I��1۰aF!EW�bP"O���dc�v�� ��02��1"O����6 �������$*�2"O��ց�M�ʁ	�̓(#w�p�"O4a��GU!e[��c텦D�|0�"Oܽ�b]�yC61�`e�
a���W"O�!�M�y�(�if�D�J4��"O҄�3b	��D4@b��Q )c"O�C4욃f�4���I�J��"O��2��ɹ{�ZM���*jR�# "O��#s�^�tRRX;DK%bj4I"OB��1BU��Pacr��IM�@e"Oj9�*ީ'za���q��Xr"O�<)Æ �,��	��]6E_�p��"O^X�'�P4+�YABL|���"O
X�t�%3�-qUA�Eʴ�P0"O�Ը�m^76�L��'V���8�"O�$Ƒ�2�z��� �K>��3"OP�;(XXH4[�E�
pj��"O.�s5��	��)���T��1#�"O�I�H�U="9���/ߴ�s�"Od�#Bd/�:]��0<���b"O��0G!��LE�|�ŇϥP0h�kt"Ol�� �ȍ��(��d�!	7X��U"O�US��_V켹V�MR����"O8Q+l��:xX��"�$��v"O���7ꂚ��1�D�P�J}�8p�"O@�W�S�<����%6�4��"Ot�H�	 V�d�H ��9bf"O �B��⺵�眃�J��3"O�P0��t�U�U%�2!�֘��"O��)ňr,$+��7P�H�7"O>9c�dw�~-qAj?Q"ୢ�"Oh�r��؆h�tE+�(I�pau"Oez��7N�#T�Y��`�3"O,�i4��1.JQA�M+I�b�� "O"����Y��@K��	�e�na�3"O�xJ�2R�ah5�
!k
�E�g"O�t�AdKj�t��왕t(X��"O �2	B�~*�)I"E��]b��pU"O�C�F]&9�j욲ˋ�d=���"O�0�AC-pcr�� ��{|=�%"O�8��)M<0s�i�@�r��1�"O�)Jp��1f�*7g�.Y�D���"O���%K�{D��@�E#��j"O:ؠE�)R,�p�O��Y6�(�"OlQ�`��{?�l�Ä�y%�t�"O$=��^7��!󇢊�M@���"O� (Q�&wH2�1&��2L�@�"Ot�����~Ā�v�"B|}�"O��Z���Z���X�`X����"Oj0:M�	If1��cU$,_hI�f"O� xl�@�f$�E��Q�TB��""O�͋B�]ۘ�X@��f�YH6"O�-�����怙�S(�&}��"O��9p��3`�@X`��2;V�"Odm�4��(BY��^=+mH�!�"OJ���D�h_� h�N)T9T�u"O0X��'�%V���4-]�<34��"OTA��X�E��@�F,1TŐ�"Oܘj�)A2{�D�hV�T�2P�ȓblܱ��!V��P�%`ڿF��|������щ6���y�eć.���ȓ2H����.r�$Tw��n���!Ӑ���Ѐoa���vh=8�`�ȓD�H�!�)m��8a��A,	\���ȓ7��BR4�tY�SI�*Q↩�ȓ{l�;�հ�ĵ! M�R��(�ȓ�T�����;��Ȃ5C� �ȓvǖ���f	qx�q��|9��}����$�/q�*컷mҚ(6h}�ȓo(d(�KĢ#��[ ���@�ȓh�����*r�2�AC<�ȓZV|�[DE@>L*�jd�@�j��m�ȓCx~���d�*re��H�� {T	��04�Rp'�����S�/����+����U�N6]|��dO�0ʐi���"��U�V�s����TeL�T��-�ȓ(j��h�M�n�&�üi�*х�7v9p��S��1���K�$�ȓ]�2�tp؂H�i�c�`�ȓU�V�cCJ�1m.����Ԓ/K�e�ȓq�Q�!��~#�M��A�Bh��V�( #`bN'G����1�Ss���ȓڂHRĬA�T�HP��Ї��i��Z�$���(�+��Y����4l|���5<T�D��`�A��!ɚ���1�R�3#.��کP�A]-�Ɲ�ȓb=��$���ȳA��'��m�ȓPQ���gA+TR0xs�Y+E)��Lx,�FTq�(� _t�ԅ�K��֌��d��s��
L/8���P�8��(� ���"CTB��ȓ_�`���/*w|��񃀟1i�d��,�. Pv郅E�H���K��*g����;�Tt��'%%�`��B_�-�Z��ȓb���Y�A�0-���A6#����d��i�F:(Z,J�,� p*����Yr*`Q�&�y�V*�m�m�������giԧ_� ���x��5�ȓw#��s��m�`�R�� )�Ň�n<$�'��5H���C����ẍ́ȓ1X)�P`Q�y[\Kfƃ�v�*u��@2,iz%O	, �6���f�8�d�ȓK|���¥�~����A��`���{X���-��d~���!�T�0�ȓ*� �SkU,�0�"�A1Dh�ȓ�֕3f�Ɠq��Yp��96���l�N))�g��03��h\+`���XΤw�3vX�@@�̞=�p͇�q�έ!(5	�Jq���`[.�ȓW#�� 5�3��XPwB��,uL��jy�Xe�X �ə!�ׇ2���=���K� �Q��j�:�b @�I�\�	�g��A����?9J(x[�K`�C�I�F^ȸy�A2pQ�Z�I����C�ɐx�7�H���}��,9i��C�)� n�@1'ZG1<	�1Ĉ2v����"O�zG��gj�Sc�]AFL�G"O
��K�FIl�ۂaS�*<��G"O��@��	6��lx �-����"O�I���:|�� �E��J$���3"O4���ɕ 2D�PnHP66��"Ov�
 �1C����mp'V��"O��� 6N{��r�e�BL�!���+~�٢�d�nc�T���T�!�d����s�-�(-]+J˚$���ȓ<Fj��q��:#�P�j�犑{�*@�ȓcl�{��oT}
v�]�v=�����!��Np&e�$�@�2�d���!�p���~t�t������a���ڥ�wf3.Uj�	1j�:>w���gF�Z�	�(j�z�*�K��J[a"O�7�^��@L��`�o�̅ "O��B�*!�Ip�����s"O�U
4��^(��7Ξ�E*]!"O�Er(���a�'k�)d'�<K�"Oċ����V��j }d`�d"O��	��
g�P��D�ñ?=*�q�"OL�zS���G���(�=;���"O�q�F�]6�u�#R�B/�%�S"O`��֮�k�yCU��Ы"O�{�ʘ/Q��7��<_�٘"O�E����4�L�G�	�kSV���"O� � X����#��8:�t#�"O�����*{,�P�ac�?p̕�"OJp����$�d"`�1
�$�&"O2�#��$]����vR�}�h�`�"O8ȓ�d�#�UaQ������	7"O
I��B�I%Jy�`�C�A}x���"Oz�e�?ÞM���L�e��"OB�O�	�5cHXԖ(�"O��	\�t@{�j�
L�ʉ��@� �y�#ֱDŲ�;',�*@����y��7�X�� �f[ ��f�՗�y&�*�T9*S($/?d�a�́�yr����N{��-)��A �,�y�I�'u���S!�H�6�B��y|�@�\(�J�KF�nK|�a��5D��!�lL�f��(��mD�qz��ZHB�	�7�2H��%C||`�ch�5}2�C�Ɏx!�͙�gV�g&L`��&"��C��;qu��� ��F6dq�k˛��C�	_��b��~'�@3�Ŋ�RlC�Ip�b�*�C%s�p�!�J `C�i�� V�@?���W!��U�m��'rz�S툼n�()7ŏ4���'4x�1�g�<�8<�'�A!u�,A�'l��`�F�?� !�J�|�����'x#�!uA��K�o�Lb	{�'�B���1S�L��ECT'�m�'�\x��Q$״̳�
��Wu*-��'�z����%:h�B�ՖR��|��'9����C�c�Z� �d�;%�Ex�'����Diو@���4e�n �
�'l��b�-D�oݶ����оeB<��	�'�jw&�;h>���
Y l�X�'a�M3�Iscԅ�&�Ĺ�
�'l��悍?���`��t��);	�'�b���ŢU��K�
;t����'>̭���7v(�B�F�x8���� D�C�՞>؎\"�B��$���['"O��"D�6L��� ��*Mʠ��$"O���P�����b��_�ڡ�A"O������0Z�	K�E��I� "O��,���1�??Fz�#"O�@��nF�T��T�@l�㬽��"O���R�M�B-hƭO�����"O~- '�#A�~l�"M��?&���"O�� +��3��@��[��Ÿ�'�t�PCn�1'��;�I�2V���'ܔ)�͗�)�F-S���<YF�h�'��bA�4XKvA_:Xv����'�.�LO6Y�$�Vc�8J�8��'��X�mɉ�}�����LQC&C�I8�d�+�� �TEy��ǜo?�B�əY.E���D�3+B�$d��6��B�Ʉ_d3�Ĕ�D�R�U*l4�B�I=$��0�&HI��9
�	�>�dC�	A����B�8^?�ո �$o�DC�	�M����dl\\jP�0�f��y�h�,� �A��Q�"-G�4�y� �
؈$i�D�
O�����7�y���+�D�h���^/�M�s���y��߁xQ�鱇*P6[8����)H��y� � PyD��!\*<���D�yR�¤n���S`"�=�� ��
O�yBHR)H[°r�Ț�5i��A3��,�yr�4D�l�#B**2Xɓe
��yLF\tA�1���zjxГN��y2�S�*�x�*6(�8lDIᢄ���y�͑��
��ƫչLu�d�� ��yR�қ/o�M�ե�;@hIs� 
�yb�^�Lz���!�L:D������y��sQ��4IN�`��ҡ����yB�=
�D�8�gS(eb0�t��3�y��ʡ���C���$%ҹb����yBT�S��]��'�3�phB���yr�'�r��eUI��@#��-�y��ԣ]�N<���:.~ET�ھ�yRj�"[l��チۃ@�:H��HD��y&�=v�^���,2A��ra��y��U;(|u���M-�Ȍpc�Ґ�yBD޶*L�$@3f)�f������y2cB�2\0��!�S�P�J���y��,Q���Cʸ�$a:3�J��y�*F6�|M3Vʍ=[MJ�K���y�-�wc�a�j��r$�2�u��jb6��E�$��eG4�.mE{��'e�<�EA��b��"�.D������'��������<|��Ɠ�K� 3
�'͠T�g J$#���8���F��ِ�'v��K��uH���@�˭;�^|(�'r~0�!�Is�\�0ē1�䔚�'ƴu F��0SCE˗JŻ;����'�L���d�&e_� ����/߂a�'4��"�柼<U"u+���j����'b�!��ȏ ����#:�L��'v�DA_�C*�� ��^�7��
�'(nsVB_�3PNtc2H^� !��'��)*��۔+`F�c!hz1lX�	�'�@=R���lD	Q��E����'n��4�Z�y�R�c��R�Iu�Tr�'~����4�����˼,�\���'�ʴ��kF$x���2#b�9vIZ��� ����2(~�}3�E�%F}�Q"Op͒4fV|
��z%�O-Nu��"O@��T��[jDMѥoSO��(`C"O�b��0I��m�����b#"O�T��'I�����=�Rq�V"OΑ��F;O F�lǘ:���w"O��؃IĤ}J\@�X6ry���"OBqc��A�#C�끊L�,��9"�"Ob5y��w�j9����O�d	XT"OzBB�̜����3�Ƞn�ԵH�"Of����n�AƩ��k��E��"O�!�a��)�B!BFW�n�.T0�"O��h�,Z7v����V�*��yE"O.D��Ϝ1V�b����9y�j9XW"O��Z�@qS|��R2A� ���"O��J��t#�#��ԅ.�j�@'"O�F��L������3�f��d"O���b-�X2h�"j�$|�X�J�"O.����yY�݀�		U�r�R�"O\4��P�V���P3*I*F���@�"O( 2'����j�O΄Jä�Ȳ"O.�I��Ӷzܜct���K�0Y[E"O���ܲD#l��B����`�q"O6=��I8RxC�+ʹ�`	2"O�����͜̡ 'k(d�|t� "O8�;� XE
�a���\(���"O�h�!�O#Uy�pbŗ}�(�e"O$D�kQ/sT"�"
+� �R�"O�U�e���Fo�����!�"O���P�7�`��E�}��@y�"O���ukA� �>zP�ƦTR"O���?PJޝ1��NM�y��"O�tB�� 
a��d�U�I(�R�"O`�{S���12��3aX� �8"Oh��F*l�.��D#a��a"O�hk�&IY�D��/�/Y���"O��i�-
�c��@� _�t�r"O
�$%@�J�d���P�(�ޤ�$"O�Hr�S�Ah�X�c�:����"OL@�B��Gr1�r�D$�<1��"O���S��^����GO]$`����!"O�%�pe1��0�X�u����'��,1�рO$��+��E�:zT���'��=���˯q�4e�th@,
pdh�'�>q����`E�����$�9�'�L@�Аt\ĉ��͜	E�d��'�^�D���r�|#0�֒v*��'� �X�oX�9���<YL���'�e@�#�5� z��S�3�*x�'�t!�E�-?��x�`��%S�Ё�'�Z�
�jW���H��"ـX0�'��P�)8����F��d���'"D�GiT���Z�+HJ���'��U�h��'�fx9%�����'�\��H��0����̘�2k>���'�$\R���.�f�+���.?X(�	�'�Z,"`��?Ш���D�M�($��'h�e"!CU����r�[�K�Uk�'�T%�i�-1��K�K�P�Z0y
�'b:�@�-��"Ud�W�Id�y	�'�2 `�'�x; �ޟLA�'�,�g������7���z�/6D��b��P#�,X�D�:i*��2D��I3h]�upt2�BK$i#���+D�� <�2���!%P`�%�@;q[�m��"OV|�в2ǢYB�B%l��"O�$�#ШJ�v��BX�i��Y1b"O�h"�
��'��y5�I���!�c"Od\���0�L��D"�C� �J�"O V�#tR�`�b�C��x"�gLj�<a`Ş�\�b�	�1]�1
"ʝf�<ө�	&��d@�g��h�V�kł�L�<9��_9/ (Q��׼*$D���D~�<ّ�U�lϤ5����5u�jt�6Oo�<9gJO==��8y�-������R�<�7�
�#@���� Z�<�a �%. @�fnՉ(�ȝ	�N[M�<ဢ��@)Ze�e�Ӌ{Zl,��Qq�<�,S��IZ�`�/q�A�J�i�<	�� �&P�R��ۄ	�F� ���]�<ц�*Y� i�6<��T�G�[�<I�ݾ'�ݒ׈��%�r�`�T�<A'��yF`鴪��lŶ �g�[�<�g�'Q΍��A����"�Z�<a�	���ji:�lL�B"����BR�<��,�kZd�FNH�5�[GI�<q�h�
f}K'�7.����ƊB�<�]�C�� 0�kݱh9f]څ'YF�<)�x?<,k"�P�5��Q�!�}�<�2�H�'��)��Z1x�����_�<�cEċTBQ�lR-fu5�@�_\�<y���?f�N��ɚ�;
�!��T�<�gH	�4�^8;���"=+�X)V��R�<�P@G5;c�I�E
�%~���Qb��h�<���N� �� �Ŋ!h�,1�o�<a���?����%�G�a'�Hp Sm�<�ÅFG�,�#��D�CnTՊ�,�f�<y���B����eL@�JH����G�<�E sx<��5A�	4����D�O�<!�/,-$���
�#H<=��lGW�<	P�O%8�9Ο�#��R"M�Q�<���0ftq32,�?>�I#�JN�<��b�uׄ(pV��@��U��j�H�<1e/�_gp�E�hi�#�E�<��#�������^��ഈ�}�<a1��Q����{+d����M{�<I6�ȤW�\�x��O5���c�s�<�s
��v��1���2*Ѱ��I�<��b��K��:���+	a���"
[E�<��j�+:�Ma�.βW~줚�g�<��KܤE?<y0V�L�_��T
GIZ�<�&F���5-^=��8�L�A�<)o
�q���eOe)"P�N�k�C�	Hc(��"�#2q�p�ңr��C�I�Hz!SF���@�u�7�P�GۢC�	����5�� d�)��B�4E�iS���M�ָ3!�0��B�ɘq>��M$Q��;��[�u�lB�ɪ@�����aHQ�U1aO�k�.B��%FyP�F��`�v�Sv�L�>��C�I:lKpU� $]3+J���-׳-u�C�I	V!�1�*��l�(��3��n��C�	�Mdq���2{����b���B�I�]18��7`^9�d��Ə}��C�ɀ#�,��J�vo� ��L��7h�C�Ɏ4^�@�WJ̝X�fL�c_!nC�I=��0�q�E9iTi��۠@A�B�I�`[F%����o'��*p�B�)� ,Qs��$[�X[0E�(h�Yi"O��rˊ1�{^͸Q���¼�ȓYZ��/�� ǲ�0vNA?�J��ȓi��H��'g�& ��ٻ�D�ȓA����яĘt �U�Uc�:Z$����:T�а��޾?Ղ+���6W��TZ���C!PS4iR�^�����ȓVad Ⳮ�	%���5�˾Cc���ȓz�F��`��
\�oǠงȓ!���0k׷b������݁eB��ȓ�d@է�VĜ���λN�Pq�ȓ)5�s��*j�Tېƚ:jD�t��C�IA�0zf��rU�L�rZ�|�ȓXy��!�;B2j��S%�?Tie��&RTQ�fKn��Qg�7O_}��%�>�C(Z(�XuL�
v{ZX�ȓK�|� ��1n�0�iC�LV��ȓz�;���pϖ��D�a�ȓ?��y�s�"q>"�yv�KZ,9��@т=!�@�������q็ȓZ?�!�uǀJ��X��&^p3�ȓ5�}�� a�Ń�Ij0��MR6��%ČSlH�� j��i��|Y@,Eft-�aQ6�>}�ȓmɤ���c�'��=�q<�<�ȓ�9[�(�+� 2�	1
d����83慈E��7B�m�d�22�����5ΰ� ��A�P#
O7� ���$��<Z�Wk�b�@0�Y�6k�܄�F�P�
~:�I##�(Yq���ȓm����f��m�Ht��ƌ�@�2������g�ַ!p���ǥP�:�(-��BRj��$\�7��9�MY�LK,��v�d�SwmH�s0Ґ�v��aR$��N�"�a'm��7-Z`�A��?DzB�ɤTy��I���->��y�lA�/n�B�I�nK���G��:U�La���]<C�	�{N���K�?#(<)�萧w9�B�ɑ9 X���Ǝ0��a���Bj�B�	�d�F�@�o�l��%`b��B�I�a:r�c�k�+��-(P,�f8�B䉼=�����x#���fԶW��B�	7L`�M���W+T�xᨳ+�j��B�ɹ`��$�U�ۓH�)6!G+f�ZB䉽g2lY���"�"Q��㊈3�HB�I#L�hP�#��2�ElH:T�NB�$mERI��-	j2�����Ĺ<�LB�ɗ�~��`(Z���0N�6��`�'�L��G
��t���u��tX�'ހP��H�[����@��h�lm�'���wÉQ�i��?_���[�'-Ly����n�|0��@��5
	�'e�5�R0P�T��"�25�2��'�l
�_<#���n91��l��'���&�
<F��V+=�8,{�' �|*t���S��-s��� fƴ���'�N��6��l�a�&m�3t�jl�
�'}<)T��;a��{�Z�Z�pI��'�,��m���V���e�j�'`�x�  �$��a���
[�.��'�Vu���I�b�H�BQ�_	Z*a��'<���t�Z�A��2!
����'�(�cثp�"xPcS��Ԑ��'�v4#C+禙ز�AK�A��� Bm��@�=��ةV�P�Z�����"O&�"���a�|<�@ͷA����"ONA��NH>�y$c�p3F��f"O��'��!�B�����wD�z#"O� �@U,
>�33�O���0"O��j���H�ް�a`F(y���"O�����@�p�*	���>��т"O��ۇH58t��@3w����"O�+%�п4o���2O�0�\�Z�"ON�zwG��w����-�.H�쨋�"O6	���
k��5���Z$QB��"ON�#��	2K׌ ���L��|���"Ou���B'{ƪ �M<3��R"Oz�K��
l��a�G�K�"O�����]�^�)��#'��q"O��q�͛�Px#PG��Y]"�G"O,�Q�N�'je���.1��g"O��8�p:��ڲLt�チϸs!���@E��e�?-JB�f'o�!�$��k�!8ݩd��Z�\�!�D�-XO,5r���Y0�y�@�l�!򤞹k25���Х`ݐm9��"B�!��4+�8h�&^�*�0f���!�J(H����Ą�G��M!F9U�!�dW�i��,�7mB�Z➽��-�9�!�D��h���E�N�8Φ���ݙ#�!�$��"��9���'V�ʴ�޹v�!�d�%>�r�P5cB�J8���u!���~�8�6¬r���� �� e!�d�q#��� �B�W3rh�7�>M!�Ϗ��P�!�'6mf`U tK!��F�j���uC�����	5S,!�(,V2q��_
>���_!򤌸)��ݪ���]^�p���a�!�䎚:����\P\�vlb�!��/Dh$�mߗCx��Ta�4�!�K4��-xp�L�0(�|qQ��)e�!�ӆ��PD�߽�{W��	H�!�D�3'L�́��ɝ
K��De�!��ոMXdmi  � 0���@�L �j�!���zݔ��#�ʻB�xX5,��7_!�$_ |Ʈ]��J�;�N� ɍ�!�Dt������z��!'m�3�!�䂆G� �������#�%�9X�!�$w���Qnͤ�6���%�&�!��dp�1��!�&x��F8,�!�$�c�.��V݀v���&��V5!�W�e�.1H`h�	���Є̃I !�$ޗKR�`�J��w�N�K'!�l!򤜷5��ꤋ� �j%���C�D"!��@K�@p��VL�A���I�,!�$Ҫ�f��
�g?j�h�7�!��C˼����B�m����\�E�!��� pV��x3k��"U��^.$�!�Ĝ�V�)5o�\E:�C�Ѻ�!�$Q)��5{A#y2��
�S5!�$=] �	��-K!�	���!�Or����	�I��%B�`#|�!�ă�k*:L�"J�`�x��`�c�!�$V�r͢���)^"�Bm��Y��!�Dʔ���x4I�SR�\���ēy�!�d��9�q��Ą�t2�-���U�P�!�D�,6��Ұ흽6u�2Ύ�h�!�ET�T+@�� �*�LN u!�� �(��F� r�`�\��-��"O��!�@��$���Yؚa86"O>8�b�6D0� /���@p"O��9�(�m��8���M�!����"O�m���ӻs,�5�5�y��3�	���+%��<u�)�&�$���)pDj� @�7qO ��9Jb4�և�X�.���4u` �O�t���1Yf�K4�	wY�����ĦpR�Y4B�8��Hɡ��@*$��_:�9q��/uf���)�M��-���I2%����O�nZ�(�O�P��+J 5N|hPBj����E�a	�O����V�{}��hj@���d��ۤ��p>�w�i��6�f�8૱	� 9��ѫWb�4N�$�a�
�M�fV�p��	qy�O��4�x����D��d�#�9t�7L=�¬/{=,<���)z��ڂ#ܨ��O��;-�`�����9��� ۓw]P�lZ�FM�5h��=A��ncC\��I�<"k�t�|��sj��S�׮r>Yk�J�d>�o:}h����ٴ�?����il� AwJ�%����-�.���'tBT�t��	<rL�Wb��DSD�3=�#=9�4Hq�֟|�U?���I��I�eA��N:H�Q�������'{04�lZJX��@��ƂLy����-սs�����b�&����$P��A����/��H�'L1#<�Æԯ-�8�e���t�Rt�!�ܷL�Q���I(e��E*5N=)����O!�fO�d��'B>�q�3�a�&��kâq"��OJY�0��O4dlڰ'N��<�����d-+�T0�� ���HQTBѴQ�Q�P���6@��m���xiv��,uq�M�t�i�7 �����X�����$�����Q��G3��1���ox���	��P�ȱ�ٷ)ab���oMƨۗݙ+�`X�h�2n�
Š'�� J瑟@����+T�V�Ru�5+�"���a��2����LX��c�'�+��h�ūN�)'`�h��Iڦ���E�E%��5��j�jy��oӪO����O�O���h�(��k��h��آ={"	��OF��d�9^^�X��/�1T�\X���y9���	��M���?�C�i�BL�q%l�z�d�<��89_f8�a�]|��MҖ�oRT�l�ɷ Gy�1�ђI�tBG�ܯC�x��A4��a�צ`��B�AF?���i��	�C��A��]*~z܅�c��7O��;XjV���̇]��DR��?%��@��cJ�OrHi`�'-��nӐ���~B1�ֆj��h�eJ�O̬TZCN:���4�"=)1$-,%n�r��93f\�v+	z8�d�شM��i��2,ߨ[F�u/��(\���'aLĚ�jy�N�D�<�O �']�aJ&LQ>��,R H���L�.Р�ru���es|PJrCϹD`KY3�q����w����t�I!0�MV�;� ���4z�6���(9�hI:`aW=cOl��6�	:'���|��5�Bp��J�澔ˁ킒��`mZ	�����O }��r��i�ZU�eIܛv�0-���ĀME@�'�b�'��P�z��N�XLX�H����~�Q�ߴJ(���|2�OD�N"<�ik�OR;;�A��!��9�$�&����	K� ��   ?   Ĵ���	��Z�:ti�-���3��H��R�
O�ظ2�x�I[#��y�4g�Բ �I�n-s�E�_�]	p7m�䦕��4E�� ��q�	x8�Ļ��My�֠�B��H(�Qy��7U�#<Q�
~ӨP(&m�r��xp@DB4F��r5X�T�$�����1?�E���/��7�f}2*,�1��l�?)��0��0L־�iP��uy�`�OvԚ6F� ��9O��@qJ��0~
�rt�
[bZ���(��L�@���'�,��$�ȄyQ#��!Ӹ'=�TΓ�|�YՌQ�����fn��hJ�$�<�ቭ!�'���#1���{�L:�I�h$�'�Ex��|�'�!�f�N	^PH�$$��}��-��&#<���>��I˟R��X�H>C���w�Y�D���O(��{��]�Jr؉[�B��K1�=S�,�MSV�1���"<���	��pˀ�8���(��[�HI�>q�	)?n��B�9Bw��2b^�H�����<�fȕ'5��Fx"��N��|� �%�L��t��'	��F'|�1 �?�@�"<	(�O�e(����.��L8��Ev�����$Z��O�D�O<q�	�W�؜1�O�"
�j$�wL]?y�3(o&�O����*�1	�D���N`!GK5F���l~.��>(��4w��	�/^5� �O�h�q�סe�8��F.[e�0�X����M b�\c�0�'�ǁG�'�b�S�������$�C�2��ۨO�����d[3�OL���LR&����f��0��:F"OL�y��  �~�s��A�X�"Oz���P
��)�#�;(_�P�"O2��*Z��z�1!�.Q�H@"O����Ic����B	5�jS�>D���/����+-d=�@=<O^"<����.(y��-�9��Q�G�u�<�eA�<�p��範�1ZX{A	�z�<��a֋���3��(�d�J�b�<���ȃ ��q�bC�*(����o�g�<�5�fe6I�3�P"#�Qe�a�<)��ɶ,D\
�g��bA$_R�<1b ^<�~xqP�؃o\x�2'D�d�<����,�p�J�	_4���A`�<i��Vp��8�5%7NN��U�^�<�p�%i��wIBYɒ�QT �]�<qա�T�)rU��?�t���h�A�<Y`�Y�.��|�@YH:�%1�JX�<�b���h�f�;A��D	��8�EH�<�I� +2�yC�''Zbu�J     �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   �	  �  -  �  '  %/  i5  �;  B  IH  �N  �T  '[  ma  �g  �m  3t  uz  �   `� u�	����Zv)C�'ll\�0"Kz+⟈mZ�p|�57���DB���H1�ѯ&q�5��7�$�b�ی>��+�FRH XY�f��%e$���;F�FiB�'>Հ,y�'mx�a snQ�)�8=s���(-��(:0Lݧ||<Z���I<���@�'�A����4���蟺�d	�
`
�c땘,�z���0�	Z�DΐzRf��	��<��@*��ߴ+��9���?1��?a�n�>Pc�(�[\>�j��¢;����?�
�;���q*O��ğ*K�����O\�ě�a�n�AU��8C�"��%S��v�D�O��'�b,	!���C�?ٚ'9�t-K1Nz�Q�m0\�����ؗ/��2OP�Z'i��P�2���UI֥��Q��̓��'�P�2�#L�	?� �[$��)��}���/� ��O\��O���O���O�˧�y��ېj@�@SS��/m:�A�c��?���i�R6MSȟ�n�˟X�ڴpr��md�lo�Lce'������3�U1�X���J۾�HO���k6�'x S�����0�&/���v��o��@ؖ˞�x`���ڴfۛ�{��I���CwM�
P0����W�k��f`H ̂ �fyK�4c$z���� '�YP���,S�h7�5��aP�d��4l���M�V�N�0�rw�<8��1��!z]�}`pA��G^~��u�i��6��צZ���A:���v%�	Xh���M-�4�@�D����G�#`���pKJ�H����ώ�M#&�i�>6-^�q%��φD����fo��XJУӂYO\(�g�A&H"qo�����1ʉ/m���d�c5�m9U�ٟ��?�C�. �R��$�¾eu�`a'ǁ*Su���$�
����n�8�m�?���� W$�2�8�	0|�8xC#Z|���K'�5�ؽ��t2:9��(٫A�#f
�T�ȓ&�� 눓��#!�ӣMB$B剄�t��+�Xy�p@ѯ
sVB�	���'��Cf��yүY�3:B�	 
�,"
(�J0q
2"h�=Y�g]T�O�d��q�KiP����\�"2�R�'��jT"J"{Ȯ!rP�X2�X���'��:�� �ĥ�WH���
i��']�0+qo� Ub�@�7�������'ق����[z�+B	Z�wA.l�
�'5<%���hS�I���8l'4��#R��Gx��)W&��4@�T�9�%H�K�{�C��05��e%�� �\�%Iרz48B�I�c(@�ȋ~��Pi�㔣p� B��o�^��f���b�+��b��C��,9ej�j��+_%"BR�1p�C�3Z�ֈ9��0m��:�H3M��˓/=J̇��-O�����)e-ь�)"C�%��I0�F�%��̙cm��C�Il��ӷ��2���	v� *o,*B��������Q���h�fѴZB�%"�ޘ�R.#�bro͏�����9H8�n�۟\�	�)p�E���9�nek$�V�T��I������V��`�I��Lj���ƟP�'��N�zΠ� '�
1Ϝ�2�F7�ax2!Z�ː��X�CQp���~�pgN�P��rF	V3{ f����;8s<��O:�o���ء�+��s�$\�Sp��U`Sy2�i�R��)�=,�J�h������L19&JE����'MP�Q�m5��a���D�O���B R5$��"�&V�J�ã�'��I�L��u��ӟ�'��'K�$F�L*���]3�*M1Q�z0�	+.�A���;�l��9���p���M��)�@��.�)§m�ȵ��.�
J���U��j�I�'�����?K~j���h^�Q>6%(%	�9@�bI�K����?�	ӓ*�\Ĺ�Hϵ6�N�Q U-��D�9ڧHՎ��wȾ�p�C��>f�	����?��g�'P��F!�����B���<Y�'�(+�&k�|�ǃ�^KؔC�'&��@��Y�D����DK��MLM��'�T2@��9�V�kW�����@�'�,d21-�3< I��#~�r�'H\��H__t�R7қG��ܛ4�Ĳ�yB�'aH%Bg/��q�6����T/���A���x˚�Cw ����!o�`�2q���Mp�m��'p(���(c��Ш��~�q� �?�@�'��AB�'�(Dô�D<��0��'@�s&�1
W�49�A�7˔�N>�U�i	�'1���<�I�;q�6�c.�d��y��@R���\������	6$ $j�ݳ^� �)�-��f�,�� �I(�산 4^l��)W'.*���*0�"�flr��o�����?w`�*��-�FYJ�f�'M��, �����O:�u�'V2��XY�@%�JH"qO?��M���%���O���D�ilĺp�
>e�����۳�xR��O�u"���Y�.D�G�<ɼ�A�'��I6fך0�ڴ�?�����2��R,)�7�����(��kρ1��'#�Dh�:�p�%B�k��T>��O��̓�*K�.Q3T�ߍZ�����O��3�.��ڴy��A�@���}�El��aqЕz�b	NPx���M~�.Œ�?	��h�@�Ĝ�i����r��!��"J,B�	6b1,��4�ȡ	_����!r��?I���1D��`�@V�bc�z�j�-ZC�$l�ڟ��'Y6��pa�����Ox��<Ycl �����e��|y�"݌�F��"	�;�"QX5��&D q�*�>�I�o�	�$L@@h������9���E*H�2�a@sc,�6p�)��>�u���q�O�L�v��p��
�T�(L�bR�'{66��O�����O~b>˓�?�EG�*D�40fe�:d"�ec����8ړ�O̸)"o� p��x��3���{В�$oZ͟��I��M��������)��#�T@ce6ţs
7\�X=�4�	Ŧ���� �Ioyb^>�ϧ�^���%B�?i��c�,(]�0��A(�5������R�쁪V�����O���t�iY7��"B��<��D�W���D�RN��#���;R'l�6N��Ipޣ<��ݍY�
��b�("y�h;��O�UL9�I��	�4�?I,O��D�<A̟$�AU�͗��Rr��;qM�K!�|R�'� 2��̍1�4!���&{Z�����'��6M�O�b>���>){0�	/�(X�g���5'@��cb]�P�C�	�u��%f׎Xp���e���C�I-���ac�Yr�8����B�Y�&l�p��j��:0E�[R�B�I8
�Xy��U�;�z��'.�"�nB��;g�<T�ʹ�~a�f
�<�,�=I!U�O:Ԍ�P.��z�O��n���''�9��ҚE��@�EP�X���
�'��ty���	OS���f���M�
�'T�e@���G��!K�����4�
�'~D,J(/L�V+#a/\TX
�'v�H@`��`PE��?R�^�{�{��Dx��)�.���c'C�b�YҰ�ƓSTjC��%N�VH�3Μ�-�*�#�MD��.C�I�x|��`�U���E��>]�B�I�$n��ӷ�ˈe����`� >$B䉜3p�l�'+�%.�ΰj�@�� B�Ɏ,<�'�jh�őp�P&F>�o�T\��I&<�~��"�ŷ���%+�F�hB�*D}Иd���} �!�'jȖi�,B��v�ي��Y�X>~qK��E(�0C�ɲ��X��N�&n@ kH<,,C��
U�N�p��c�,������$�d
�$�6���`�K�(���*R�Ūe!򄇉v@ة�	M�o��I�V�M�{�!�����ʴ�[�ER�P�%[�ZB!�)pL}z5AQ�.�k�e�%!��RT/˗'����%_1E,!�� ;��K��C��Պ�$8�ў�P�/1�'i�PR3�����B��Vd����N��h#�c��M�le�q��\A��h�42�ԯ?�����jР�ȓu�Z�?PvN����479��@��x��8h!j��&`<QOẍ́�t���D��`����'*H�	 ^վ#<E���N��9�S@W�t�bEkuᕯ**!��+V�p�o�6�P�
ӡ��M	!��ؚ/j,�8 ��Z��XQ�V��Py�&�S�\@ё'��X�JiFؾ�ybI��S>)X�O�6I&��y�ə�]�����+�\UP݋������o��|"葬�"U��ŷ�eҤ����y
� ����,�nM��ʟ�v~h �"Oܝ�눢��£��t_:
�"O� ���4h,jO�DZ4|S"O�Cg�4�V�����cS�p2��'����'��AR��
�~Yj�a�L����'�4kr��q�Z�;�l�6Z�5@	�'���1I�'H�`�6m�T���B�'X$�$l�b�Y�#�Jr��#�'NF�ph~m��5+X]~�X
�'�`��엣G�}�ŅM=���ʉ��؉~gQ?=Hb,�d�J��"�A&d�,|xB)#D�ԣ+Y�rBi��!=3���@��!D�� u�V��@��2�da�W;D���W�6x۾���O�a��0+5D�xA5�ǄU���Bb���t��2D�܃�n�gl���ȑ�vU�0D��O���a�)����B�Ɓt��ѳ ��V��	�'=r�1�n�Вqy[v��#�F�<T�� H"�sw�H�mg�$�qO�A�<� �ep�T� 	Ѵ"�ZQ����{�<I5eН=�*���K�3���AK�z�<ٶ��
d�xh"e����"��OyR�W+�p>���WC�����^�l��z
d�<�!m�;Z~舡�Q�\,�"�^�<�v�0vo���f&[V΄�,O�<ɵ�;'�	)�
ƊV��h2S	�N�<��
�吠c� ��>d�B�Bx��Q筺����^�b��Ȓ�)^� ��!D�tr����O*4H	���m�Iæ� D�D�fl|_�Yk��� ��XR� =D��Q��4Pn���I��r�`ມ�/D��Ӫ֡@f���8�Z(���?D�L C�j��-�`gD=m0��k;��>mG��Y
�T��q[5Mj�zGHߖ�y��H4p�N�~<��c���y�@�O�n}2�B�,q��M�W�G�y��$"� �5"ޚ{U�1�B�(�yRĝ�6x��;U�G�x�>�@S	D��y�m\�}�B���_w���i�%ΐ�?! ��c��������Ŭi:6�� �Z�+�U��;D�\ÃF\G��<HD�9�؜�5�:D��B��^�r����KW*m@n�H"�7D�Ęu-Я����
Z/+�`A�g�4D���Ԯ o���i7�W�'�B��)4D�x���ۍnp��.
��"e�v�<9ƍE8���u��+
� 9k1�
*f�H��dg,D��6-�'Dv�4C΃�)"��C�.D�lZ�J 0�Q��_6F�L�PD-D���d�+N>d��蒱V�ȸ�N+D��@VgW�}]��9tH�\�l��F-)�O�3��OX	ad�8`�>�k�d��?����"O�j��.��!��c�/<r��"O��Q��4Bk��J�f�B�"O:����Σn��,�'I� �<%�r"O�,"�i��s"b!a@A�Rh�"O#p��A�r��r�2.^�xT�8<��~�$+T;J. ���)�~3܀���e�<��.қC�� ˳&����/�b�<����3���:��+G���[�$Rc�<�Ђ�2r,���4��le�W�<	T���&��6�W ]Ö��|�<Rl���P@�ϋ�@�P����@��*�S�Oʪl��oٜ$� ɜ�X[�4��"O�x��!�����)uX�SW����"O� ,I�d���Hsjȉt��8�"O�����ȇo�8�Qa��#6�ɑ"Oxh�e΅�a���	􊕙`��5"O8�X�"L-�����e��=��X����(�O"A��ÃN�0y�T�S�~l}��"O����U�;\A%�F<m��4Q�"O�9�`A�z���ǩG�D��"O�$Ȕ��K�RHh��z~D��"O�Y�ԫHW�|xU��΀�a��'1~��'�i��6^w�H8&�ֶ)��i!�'	�p#�E22V>�8�k'�����'��QG��O����ⅉ-��h)�' �<�nI�	a:YR`A6!X�j�'�N�1��r��ԯ����
�'�lL�t�B�k�^��ceF�"�҉��X�d�Q?�
rO�(�Q���α'����D$D��PB�&hL�zG�A9�>�2P� D�l�a���%��ISID@�B��?D� Jգ�9L�-i��)Ya�b8D���M��]���In��3��4D�L��%�>��z0O����O@��)�x^���^��X��荃�^U"�'�l��O�IYڐ{T�+Qެ�
�'Be��$��l�xȁ���?:�ܵ8	�'������N�BM<�X
�/���	�'����bN����h��H	<�}��'�y���ՂW�$ŘdD�6`|,H/O�$i��'���窎�"��k'��%,�}X�'?lt�B�'[G>�KbjT'�`��'c��)DNO�{N6AB���	�-��'�A	�˂�8�l��E���}!T�p�'�ܬ�W΃'�I����p ���������HE��
5�@�K�1h��ȓ��})��ѫ �B�h��L-q�����h��iծ"�X����E��y�ȓkߪ���#aB�Y�.^K�t��_�Y��D/[��H5��3;�E��DA���`H��Y��#-(�&�D{�쎯Ш��0B��M���X{���	�ňa"O��Ru��"�n�����,�>t�1"O��(��6=�(��Î���h�g"O\�w-ӱ-��{�b�"u���{�"O�͸u�2NhjUX��T�5��%�A"O�Y�%� V&"5K��߄$���'�'��������>��J��Z(,x(�S�f�4���ȓ=A���p�ʩN��T#�D	�i�ȓL쎁�2#�3.<�����YG���ȓ7�͋���ҨQ�NZ?588܅ȓ	i8�hg�S�&r�8A3��/b�D�ȓ��U��*X�#�X��#��S�`�'�p�
�>���+�뉂/������X5zd}��J>d�tϜ�S��H��R�U��4}h��`���0����Gʘv��T��rnd����U �p�q��0옅ȓn�����&��k:���eI#ȭ����r�6�ɲ(��Ɉ!��|�f ��R\���מX�̼��@�)=`�;��L�G@!���
��ٲê7�hPdeX�B7!�$�fJd���$8�:�i�c/f�!�_��E��j&;�aF�L�!�DK(I����̅�+>�BЁS�:ў+�%>�'W
��#B�B4 2�h#�ʆ?r�̈́ȓyun�* N^�)���rw"�ԄȓZmb���")��h�6!������S�? ��o�-6�%Z�͔+�X��"O$���F.©�FK�7&ۊmY$"O �aS��G�႖�{Ǝ�t�'��p���S�q��)t�O�a̜�y��Z��z���P����
 8(�y���ͩ���ȓ#ҒR!Ҟ1��i�@�nS�t��q) 5�ል�*��D���E��H�ȓ+�D4���'�8��Rk�-d�v���g�����3�T1HR���V��'1`�
�8�r����@e�bICS��"k��Q�ȓ��Aq6E�q`pQ��[.����i/�Y� �<l���R�י
|�ȓ;-2���'�k����Hx������j������4a[N�a��QAx�h�&��XqW*�G��m+b�ԡP����Ў=D�Ԉ7˄!09x�Ȥe�*|J�31�:D�$����	���C �A}*X1�e9D�$���/;|�Qү�k��d���2D�<*�{��a�9M� ;��5D��AnǴ����Gf�3a�2�4��yD��+����7��E��)I�y�k��P����tcʚ)ZlA*�.$�y�h
8�� �A/|ک�&E��yDY<l؂�kς!��t�&N��yҫ�}2��j�f-/2<�c�=�yѐj�(8a�S�Թ�J�?Qb������R!�Z�)�����"4�|r:D�أ��W3I���26	ɓ�|���4D���!Zd���,��>d>@ �3D� � J(�4�P�*�8o  �6L;D�ph!mu�6@� ��th<���/Mp���)L��C��yR�����O� �Ϩ����O��`��ԮF����ʊ5+l@ັ��<����?�cujFm\�;�qKG�n�y��O�2�I'F��mI�IBL*��@���}Ԁ�1Z/�ik�ꀐ��$����j"8z��0X|�!���R�&Gy�R��?����On �1����o1h�8��\pz �,O���d��d��") y4Tmr1Q�2q�}��<1�B�.Ǣ��D��5�D�[��\y/� #��'j�I{���'k�BͲK�U< ��	� PV�-��.(�XP��J��K��x�j�}���!^�
`��D�Cd�X����<a�)N9"�4 G�Ƽ	52Ё�E9h���c"8�JH�!�<W0օ��(��dF�I���$�O��S�V~�gO)"�� ��p��y0�`�>�y"R'5
� ���kji`����hO��F���э�tz�+�+ִ���ܱ_��'�R�+�����'���'5��O^��Y�H*-h�L 0W���$�Яs=\��G�}�J�&��j�Z���
+���D�4+G���`*�׺u��E	������A-;�ΥH M�@X��#�?%�Ɨ�ysh�6��I�i �qP�av�8�R��'������?����r��:���-d�$H�7KH���FL2D��	�鋊H���+Iغ�#�O@UGz�O�Q�|�ՈY�k���wa�u�\$WD��mY�;3	J�踤����H���?1�IΟLΧE6�\`S �8&��,��"�:���ĦG�k�PR1,�+D�I��4H�"?9��O�"�2���:��\j��`!a6)�h�N=j�A>���� 	f�ʽEx��_��?�%%Eq�P�0ð1*Z��� �?���:�hx��k�v@���>E�ȓCOHA��+N����c��U��'�7��O�ʓd�Չ��h��1�����&��(u#��� �i��	�?IńO�?����?Æ,`#$��@➆=����|����?`ܝ�d��Py�SPE�~�'gŹ�3$�L8�#�iK":y�钮�Ow�d��k����pQD��O���(��1]��㲨�/��D�c*ɪ!�˓�0?a�	�~{:��5D����elSx�<�*O��1ŋ
J���t��7B
^����4J���,����� !V.��9��`��P1�Ix%�-D���%V�E�d0H�ڕ�ne��$)D��9�JB�J�4Mrb հuI��<D�� >�xf�:���1%o��rl�M�"ORYR�»B}���-& ���"O�萱(�*Bt��#��r�����Q��O<�}����Bs,C��3ӡ�6�(ąȓp=���.��8�a�1
Ե}�Y�� ��!�ł�:XRL�īƭ;��0�ȓJo2(2�������$�#g����ȓ^���5��;_UB$`A�V���s����GQl���D�r���Ƀ3>p����&L����ō�:`����Ɣ26!�$�����c� +l� �c��?%!�Ď�*�M�D@[3����C뚈R!��?5)~P觌�K��%J3
�n!�D��'B��J&�p18 r�[џ�����M�I>"��=�|�[7`�{�p����X[~b�'�"�'R���aؕM���!I�����j#�����J5�=4�<؀�sz>�X��I�fƚ1��0i��x HK:.��M�ڀ�a��ŋ�Ѝ
��˃A�x��2�I-���d�O���Oh�S5���;�T�۾	a�A�r�P�D�Oh˓���	>?q���L��"� ���,3 ��c��|l���d�u싮Qo�E�f�[7�ʴb"�꟨�4�?Y���?�.O&�d�OX�5L�Չ�iMt�r(��)�(@���'+Q��F{� G
W����e�5d�V����D'��'���K<�g-�O:�'	���qE��i=��2�OW���d�'�z�	"�ӧ�9O�@����$I
Y�'p����t Pb��Op�,�&��OV,$?�H�E�<U�܈��ꅣ:v���5M���Ɋ�~��s�L��M�M�V�K�a(�`ABM�rn&�'t�';:q�J���>�B�`��!�8df_�mt�,�?Q�@�x���U��?9pK�$wҁB�M�bxr�q4gV��r�"}b�3}R*����ə�Mcs��#\�b|)t�Y��`���ĝcyR��9���ȟ�PA�v���f��* �����z?a5(I�T>�I4�����֟���'B�|��i`�:eo؍� �\{�u�޼�'���D�T
�B�B��GL	{O�1�p"��?9�L�����!?��y2��~��?J�(�a"D\��䙈Gヹ�?��m �O���f�J�pt �Ie)ʿ�Tcw"O� G��9_�Y;�A�31�x��xRP�0$��Sٟ,��9S>h��o��n�I���#��X�O��O8�=�OR�Aqo��CΨ��Ȁ�P�؍}�)�	��~l[ЄW�z.�z�_+!��ش���*�3����7�+\u!�Dc��� IX��h$��*�=!���yAb�1k��� Bgk�!�D9;\���(ʇU���goi�!��0�����B�ks��`&X�!��3n��p�P�R7Xtp� �i
!�$Q�'Ʋe
��K�9�:pz�
ʔ�!��/l)X5#�O�:m�=Є�ūE�!�$K
A2�V2I~�x{�"M$Vs!�dO�������@S
����O`!��Ao,U )Œ&A�pQr�
 %d�O,Q�$�J����	"]��y�E�KR�P� ,F�h1�1�!/���7DU6�W�Ly�a��C�t���"�M�DY24p$;��4(4)x=椨ԤA��o�D�NhUÀ�o���BD�O�& ^y��o�X!$������s���AG�u���Q��F�	 .���C/ �D��&��'Y�#<Yϓ 0�d3S �"O. �"��!�ȓJ�d�A�ʃqk�}��J� %�Q��Y�Q�rI�dn����B�\��@��<���a�N��S�.�����M#���ȓ �&�0k֦���C3���0�����_@Y���	�2܊$�	>j����	��sXn�
���d1��b���6�[�r��b��;�de�ȓ+��31�����6�t]$p��rX5S��|�$B#��*ʢ,�ȓ	leX*��f"u��S�"����@�2i]�=ҵ�4�ʹRFp��S�? R�)�D�."~��RfƘ�N@�D"O�0p���wK<3GG\Q�b� 6"Op �#Q�=��L8U�D�{��|��"Oܬ��V�4����Cx%`"Op���*zX>��B�%<ʼA�f"OQP���@��<;#���z���hD"OV]�C��$3���ϖ'�<ɪ�"O8x	%�Ւ9��T�%��P�v"O@���Ub��En�2X
��"O���a)V�C\����j�>CR]��"O������9���)�<\*�"O���wE��U���R�G�' ���"OhU��.J7?�F��򋝟uR"O���(�}�H���F�Np)JB"O��)gf�0L�yp���%�Z��@"OdY�t���+�)x��\	"O�m��D��l`|�k#h�.�Va T"O�@Ѝ�{e�0R"hؑI2�̀�"O�$���C�V�)�MP�2�R*6"O�ݲ.[��t��
>7�
�s�"O~��mX�r���WO��D��"O��QV�{� u��JعWmz�5"Op��^2s�J��J�RUjl�"O�!��� �"��sc˄Y����"Ov��%�C��||z�D޼;B 1X!"O��0X����# O<�A6"O��%�:x�!��eΐ\1�"O���R�B3�� fA0�E��"O�h����>���B�
��*����"O��#M�9,ԕ��)G'}� ��"O�лэU�gj���A	���"S"O2��ݧh�V #� �2o��Q"O�)�TK�]�$�O�-/�>�Xc"O���O08���z - �Iߠ)�"O!��0Y����Nk�B�r�"O�M*��Ӫ�jPY�#¤��E"O�t�mշ �r�8��+"����P"O�L��F�{%�=lc*��Q"O�%�.@z�����1{v]RT"O��!��0�b�ģ�,Z��"O�S���RԠA�FÃ�S4��8�"O������36
���"�<mмI�"O�	kUă.Q��TCS�Í��"O� "�F->�����/.g�~�iF"O�D���Q�a*v���ӛav��"O�ä���y�,
��?U��"O��.\�,���-@T kRkɅ�y����U�ܨ����h����y�DŁ HK��+jJ\Ј]��y�d�2��	xԇ�&�\0" �2�y�χ�k�`@��"R�'rN�@�9�y2GƫJ��ĉI����O���yrb�I�f���ӊ�v�	%C��ygE�td&\[BB��}�����y��}��E��*� � �bE���y�5Ѻ��ī|6���Q�yR��-��b�mtԞ��Ѭ��yb�A�\���D��r}�+� C�y�e�5�J)ЖAęc��yK��N+�y�� <XЅ�«U�DQʷ%��y�#��;\�ьȋGdm�G,���y2�W"<ـ��@�7L�p`�Z��y� R�"�I�'
=6��)�#��yb�$o��8�����3�Z�hf�4�y
� ���a�E!��#BE�2N˘�2"Or}��(V��^��ġ�'(��x0�"O��x�o�2��
�J��>�c�"O�ɡ�	��\Q�*� 	Ϛ��"O���N̈́`t^��lѰK�`�	""O��@V��hچ��b�F

 �v"O�̀��ݍ'�	��
m����"O֜hG�ЙT1P�1�B�?��Ȃ "Ov�cэF#A�j��t�K;\�Np�#"O�yqt��0F�2��_�K�����"O~4��+�i��u�0����H��"O�ȷ�T]I���q��l�]XG"O�(�#��|q>\{������"O��(Gg�cTt-a%N޴N�^ْ�"O̐:$O�P%��m�Uh&�b"O�`�T`�s���U�X){b8Y�"O(��E�W+(��L� PThQE"O��qB�I�>}j�˶�j;j���"O��A�(�w�Z�X��	R2��`�"Ov<����!X��=KGL��p0&`b"O��r*E#d/�����G,P�Yj�"OK#m�����C�?�^�"O>�$�H?аt���&�1
�"O�H&���t!(�b��S0%-;S"O����&��Q�ɣ#4���"OLApщ�����6��� �P"O�+��=JWF�1�e�	>Feڧ"O�4�4���?KP���?$郖"On�YUm���l�$b��d+6�s"O��3��Uv!y��H5�5(�"O�=4K�h�����!R�W����"O����#�3j��b��0j	;e"O Z4���D51��ƕ^cfm�"OZ2sn�pFD�:�O�CEJp�"O��{�n
�\��܊�gܭ]).��"O,�3�+�q��Arc��	u��A "O�4	 A)����!jņX����!"OjS$h�6A��K$i�6l�"}��"O m�nB:=�8h�P�h��$r�"OȘ�Ƨ��sy��P�փ>�L<s�"O�>;���bn(=�b�A�"O��`�CK�oH8�(c��k����*O����`ؿL��r E�T�[�'ֲYѐ���2l˂g�PڒQ�'�FQJ�)��䀡a���3/X��
�'fZqh��h�"�!�
(b�<�I
�'nd�Z�f�"�����ϰMK>͚	�'V�p��\(�t�ǌ³?VD�A�'�E!�֓X:
�@7�W7��`[
�'Ω��.U�u��Y��z��
�'���Q��/=�@���^�b�t���'W$� �dI�;�l8R!�0O���3�'w��eG!T�e�򍊗PFν�
�'f���f� AD��ѫ�H�F��'������\�%���H&ԁ�
�'�R0�L"FwV� ���r����'Ȗ�A�܂8�����lа���'ȶ�y"/�wġ2eˎ/4Z��'��[ATU�"�i%F�0��}
�'ܔi[a	E3+�"K��(�z��'� �j7`]�,�N �đ��z�;
�'���b���&��@0�� �$���'�8E E��l���J5D�	{���p�'��tf�K�3MF����lf}���� ����	���@q���3�(l2�"O(QIըW$r��8�D�	f��
`"O��A�іxI��� �<�\h��"O00Q�70A�}+�$N/(`Y�"O+d@�e�V!,��\q ��.�y2+@=b��!���""�
�b��yɜ8;��0��!������Z��yB`�뎤��E�K
�R(�0�y�l��Mo8Q["�D����a��yB@�#�D@��7x̠�搕�y�h6��$Z"�^�y���A�ņ3�yR@�(-p���Q�n�xqi'X�y�ؾ+��h�����3(N)�y�ܝBpf�j '�H�u����y��+Y�J�@��6"��b�Ά�y"ƌ�!&����9to�������yr`�D�ȓ4� �g#&�{A�G��y�I�_`݁�GAg,,<BBj�$�y� �#gY��I���X�"@wa�y釻J8T���%#��P���y2�ћf�.�*scM#<id@���y�� k�
��$\ANlz.��yb,O�.���D��UP2(�OC��y��
�p����� A3Q�����Ͷ�yB��n�T���!��5h�8b�]��y�$v}�s�� ����a��;�yr�^?*��55g^?����0�[��y��R�t?���d� �RXd �y�d߭K�T�g)9_��J6����y��6>#��b�G"u)��;����y¯\&G��	��)��$�U�Ǩ�>�y�D�5)��cҧ��r5ƌ�� �yC��dN�a��S�oN	���y"l7'&a� B��hh:�.��yr�N�@>�r��
&@�s$�F��y���9��,;�"H� ƨ�+� �y��@�OI�4�������u����y��:7�n�V�	┽�A�(�y���
��L���L��d	��y��Y@�qQi_�J�>`����y�F	:��c/�%U������8�y��ǆY%$����µO����%�y©��66x�k�D��������y��M:*/H�q� �F�����f	��yR�~*A���9�R`:��3�y�
W��H8�LΏ!p\v����yBF���h���z3T=�%�[�y"�Dh��𢠉q�0�T'��y�G�[�1H�V�d�"XCi+�y]5_�渑�	�f&L9ٔ#t!�$�q�x�WD��e��eqq�ڊBq!��j$��A��7ux8Ԉ�
��6f!�d/v�������,rR=R� F�'f!��G�$M���፹t�����ԜML!�_�w��z��Y ��94�z9!�'G7�Ո�*�F?hѤ.I8/!�6T��B�02'�]2�F2& qO�P'0T�������6J�8��|"�ֈQv9{'�A),�mh��yr���Ko*�y�� r�B����W��y��M�O���l�":o��U$B��yB$��>Qԑ:�E�&*T2x�Ȕ��y�h]�orhQ����R�\���!��y�
U�	�"L�B��T�*\��yb��- ��8خ
�fI��/��y
� ���6�I�)���c��ϙ}0RDJr"O�)�	�;��!��D^p��"Ol��瓣<� ua̵�J �"O�XQ�g@�hl
����y�L%��"O���b%�9qw$L��+�>� "O�����؇q���{��:8��"O����W�M��I�bG,d��K�"O�U[a�*6an����D8DP"�"O~��E*؄+>0��[Ve��!�"O���jV?x�՛���+
� ��"Oƙ3���E�>H�Ħ�<ǐ�!s"O����F
N�ԳC���1��s�"O�e8�jG�.|1�w+��n��$�4"O�Ջ5��=��ɞH�@d@Q"Oh8R�/ż`���7��.Z2��q"O��[E#L�@
ژ��_2��h��"O�h_b�8{���i9�"Ozܨň�)C��5�Ġ_�m	�hs�"O�D��/]�a��Qs�I%R�0}��"O���@��$�RF���@["O*	�,s4�����èi�½��"OL�"���,�p��0E[���+�"O��q�AP"����Q��,E�"OFˣjT��}c��Q�97e��"O�e�`��m�v�BT�̡(+$�kP"O꩘T��,y�PȔ8��5�"O� ��`��F�YC�׷q�t� "O�|�-�8���H��E� �:Mx�"Or<"Q(R�^�RmA��̄s8 ��"O�����ɑ�예 ��O��"O�d���7[�t[d	�:HA�1P""OrM�J�)V���$h����(˴"O̬g'�D � ���[s*��E"O��
e.lDj���ݒ[b� Br"Od����PԀ�����, E@�w"O���'� �u��胀
*����"O@�$D	-]"�B��A��.�"OTx9v,�:O�L���+G��"O��B��6Fl�P#�O��,���"Ox�ю�P�XՉ� �!P�yc�"O"�
����%-ӖH��T����	�y��N���Y6
X@�
=��̉�PyRHT� -<�3Sn�O��!p��e�<R��*a�=RC�ڙ?�Ʃ�b�J�<�w���.�T�����.�>�&&�D�<�$��T���qjP���Sg�I�<�k	J�����?�Ҭ��o�<i����LДcɾ�[�'�n�<�$���,�$	;�Y�'�S�<�flL�T\���� M�n��-To�<�E��d���×#ZԐB���l�<�r�%pPF��g-O��~����Us�<�S K&{�>��$ѓ;��ۢ�M�<������"�I����#�e�E�<�cN<
Kʽ�e��/B��D`�B�<����h�n�Ze-G� hT���y�<�kM�@�&�J3	�-�֦Np�<9��7w�n������ZW�ɑχc�<����,0�a0���hRpԲ�Kh�<�� O
��Pum ",���S���b�<I�%�"SX%���=a�����h�<��ԗ� 1�kŵ� �N�E�!��%95��j�(X�N]�����$�!���8%��A�dÕaun��t���!�� ��A��*8����J�U�"O�,H����r!L�ل{�s�"O0D3r��:�"�ó�E'���zc"O@�"��B�T�8e�'�ł���'"Oh �3*P�=Sl �bj��X�����"O����N�.�ts&�
<�H!"O�݂U���F��M2�(u0�T��"O:]���B	\��.ѨB�0�D"OƩ�1g�(ֈ��n��}��!z�"On�S�`_�q8��r '\�'����"O��S�s�"m��/�8�>8��"O��¢�H�}~��s��^R}��"Ox�p��M<&p�ؠ��ٕoB��Zd"OԹ�$iNJ�"Ҫ���E[�"O�J�J۔P0n��ǬY�T����$"O��x"
 � ĸҥIA�.�a1w"O�E�G�*u��XpH�7����"OX�H3h�nвI�O� �"f"O��h�K� E0�L�ٴTP�"O08��Z0��	r�@4Y�ܔ��"Ox�s/�B�.�!j�|�J� �"O�aP�Z$Hf	Aȋ�v�Kt"O|� ����M�`=�q�֝ ʆ��"ORq���ɭ0�F�ѓE�e$�TPv"O5B��!���fD8p�� �"ON0� O�N���.ǽ&4T� �"O��5@��~�X�
�D.�#�"Ol�P���6,3և�(,���C�"O`,����9G�sG�h����"O��`F��s�
���e�-���"O. Y� X;�����R,#�"O����3w���X��F�Y�xK"O��0"��[QN0;f�^
U��]�"O�)$��~x���D�ޚS$�T��'p��+7��W(�Q�H+6�^���'!(\"�a�V���㍴.$nU��'����D�
+R�� �g����y2�'��$j NT�����QA]m���[�'O�X
�KR�4b�9ڰS�69��@�'L��L[<"F�K���=f.��!�'Y�`:C�K�\��H�@W!Q�� �'�|����1�N�����FԈ1a�'Z��r�F�9��10g�U=58
�i�'���y�oO=)�.q���\�*���x�'�m���s��LP���*RBI�
�'�~C��4tJ}0�ܾ$��Y
�'�8�r�L�3$�T����>�D��'�np�[Yf:�"#��H\�R�'���b���:tĉ���B�8�>y�	�'m�2mR"s�(���bZ 2Ƙ��'�D!0+\�ځ����+��P�'��� i�?$�|����Y�� �	�'�\(
�O[���CʳW���z�':��u�#X`��3�� �	�'}��`g�00�����)�\l��'����e�O�7X(��/��&�<�K�'@#�$ѦZ$D�&�����p�<�PE�$h�|�@�ȚzZ&�5��H�<�ul@�_�Ƙ����*6l�R��G�<AAM<E�q�D&�$J�3�CW�<q�b[z.!B�uqd�˅h�<�iH����sA�;��h��˃l�<�A_�U窜Q�CFhJn�P�/�B�<�d�?q��=�&�P*&�^U�RhQ^�<� �,���'E%<P�FK�2�=1�"O1@��R�c���s��@ψ��&"Oj��e)T�QV*�2iȷN1�!�"Ot���h�^���
I�"#.��ST"Oh���O\!yD�! �"}��m�V"OLi��
�bF��!�:[��D��"O��(q�X'h�hl��l�2o�&��"O�Dh�ꕢ�0l8��"�.�p�"O@�:G�ڌ^gtq{G��aϺ�s"O���TƑgX<�J��V�_3n��g"O\�"v�A0k�f�����.���"O"�A�りTE���+	z´�2"ON�!�H\;l���B� ր���3w"O�1�bF��e�<�yQ瀣9����"O�p:`Έ%�pS�]���*�"OvA�F��L�r@��(��	8�"O4Y�ʖ�O�xѓ`0;���1"O�� ԍA��D�d<J�Nx�"Oz(�E��Z�P����J�r"O��墈�
��B��06��ڡ"O�(�մ�H�yF����,�"O����1��L� n��r}�8��"O�qx��[%���Y��(JA�=D��¡o�7�I�+B�Eh�<�#�0D�HZ懊.���Ǖ
=$��l=D�(y%�E�x��lU�F��U��?D�� @*��W��y!�$_�t�cN;D��z��6��h�����H�a�:D���!�0PQ�`O�Q�:��Ć4D�СP� �|]��)�k�B��%3D���E��@O��{��G�"��X��2D� k8tز1$đH��@�1D������)M���m',kڌ0��3D�|q�n�?!�蠢ҴD��2�'0D�T1&"K�'��\{��%\����1D���A�_*u�a�.O��m	��#D�@�E�~Bz�X�O�=��xѣ4D�X�����H1.f,�5n\�=蚌���Z����;V�f�R��=:�
D�ȓAX�|{�T�a]t��`(��4F���ȓm��9ɕ}0mj���F$B��ȓtAn|�e��v���SQ�U�¸�ȓ@��XQČD73�xHk��7I�Xl�ȓX4r�;�e	e���@1f.���v�,(W�ю&Y�x&o�05��ȓ��8zbH f�lD����(3�I�ȓl��h�MH!ft����*VF��ȓ\d��#D�y��ӓ+Z%�:(�ȓ}�t�D����}�a#�5/�A��3���9��9�: o)�4$�汄ȓv��؆jʖ"�����a���ȓay�Y�
_�{G�A@6�	)kf��ȓV "aԉW$��'�6�v��ȓb7�P�吹�� 蓪��]R�Ȅ�NV�� +E=���i�C�'q��q��d�e�K�]`��ې�ˠD��ć�_GLգ��
\��|��S�/���z֪e�`(�lhx�f/Ɨ&*��ȓW�^	j��2Z$��g�J�V81��P �A��aȏ;�� ���$��ȓs�la#��714�q�!
��d�=qԍ�v���a`1m>��S�I�v��,M
|6ܝ�rC��;��C䉡@�h�Srb� .U��W�N�s��C䉠{^��`���~>qH��MtU�C�)� D�A���&j<����H2E��"O�Y(�l�!�B4#U:m:�	s"OFHu'�X�zM pk�<0��@�"O�\��E�.tY*Yq��<[��Pc"O0e�l��|i�!�Ĉ�0=*�h�"O�"����셄�g��H��=^�!�d�r��ے���;�&U��&�s�!��Z>|
e�`.H�5�J�0�凩!�œ.0��쉺]�be�b$�fY!�d˾R�2��ӎ8?�V����>,o!�$
�)��T���U��-���	$ZU!��\
yi�M DQȥ���\�!��@�C�����MY�,!e�
��!��0�����l�F��#���{�!�ϪI$(d� mD�x�`q��K� �!�ĉ*�}B��>W\Y����0,�!�D��Hwň��%BZ\�d�i�!�?#@p��G��(Ḷ�#Z!�d_K��9d�E
^�lI��E8-�!���% �����L�fE)˽
�!�$� ���
w/o���[�x�!��05�2Ap�E1+�̂�Ոw!�DW�.��t���S�6ǲ���>a!�$��Ԩ�IueX(��U�
շd�!�$�z*��V��
�k�?GY�� �'���v
V�w|l1�&Csc��{�'A^<�4��x,1s���_EB@��'���ӭ��y ����: ����
�'4p��%$�5J� �UoN�t�8]k
�'��9��� ����+B��N 2�'��!!�Ð�慨�᎐y�``��'���L�60���C����'w�PC�M�,���eiU����'����G�^'1z@���N��*�'0F�QvEE�Op�9vF��-W�(��'�0T�6�G�"��E�ΦTr^��'!$�A�O��r�#àFƂ�y�'c:X*Q�%<���ɒ�˷@
�<��'���rO�{�V���kC4;��	�'�����ŋ�6��r�K�[�z��	�'�K�(+�Zyq��	�x�,�gQ�<aԀ�7	��$[��yG�PO�<1����	�� �;4z4���Mv�<�O.i���re*O�?N<�`�n�<)��G:
D5&=��9�Pl�<	W�̌_�d$����5�^�q�g�<qu't���!�	�O� l�f�	=�!�ZP]>�sA!Q(~20�c��!�$>x.�;�I�|h�=�s��cA!���3n��ʠ�MM 9iDT�j	!�$I/T���t'�a=XK ��!�D��1Q��R�mF�P� 9aQǜ}�!�$ٽx��������r�+��b�!���2d�D�&R��� �Z�!�$��@�e����w�a3�MT�d�!�31C��3�h�,�I��,�!�Ďy���pQ��;���t�Ѩ�!�Ą?B�h +b*T�X��D��!�Ě�j�<�����#�|��\	�!�	>X�(0j�	�*��q�`�=#c!�D� д1;������C.l7!�D=I�Rђ�׫I�[�CP�MT!��Ϩ/v�P�F�5if�y�f;!�D�/����R7��Q�NG�Z�!�� �1!W�0��j��߮`�~L�f"O��'IX4}��M(Ǧ���̡"O���r�Zy�h�҅��`�$(;�"O���&#5/�\���e6$E�#"O�`�t/��F��s�ɐO�~�H0"O��{��ٶN%@vd��К "O�T��	ɔw�X�"�B@��l��"Ov��0)�((~q��!So4AJ"OvP��)O�ಯ��8�X"O蠪�HS �����m�6t�����"O��6�Ӧ0�dm�VL�fvD"4"OVP�t�ƷN5�	���΍aO�x��"O�E�'g@
f�P�D	!	4b���"O���ƃ��n���B���7a` "O�X�mM`���iG�y
���"O00���/����b���/�1i#"O�ࠧaHPH*Pʆ#7����$"OT����<2����\3F�00"O��NK�7a��1H[���͹�"O�Q	�(P�WT D��[7>|��"OH�P�e\�n�*l��a^6h�pY�c"OP�`���VQ�<P�'{*�s�"ORI��(����R�e��Ȅ �"O�-xa���]!6�`�E�d�zl��"O�V̙"<D��$�w�4䲥"O��9%O�7���`J�"'�X�@"O��b��E+�nH	gh�ZaXf"O�֭�*,��#���`���0�"OJ(	R"�iL��SE˪6vq�$"O:�yf���H�)!���#DEbs"O�p"cWX_�$:�C��ޘ�"OJ�c� ԧc�����- �4-["Or8%��E\r-��	U����w"O^<�bX�^���
��E��"O�Й0�(�Kԍ$�v9�&��yr���j�r1�׀I�"`	&���y���6w9�6�@wN��	0�ybgל?#�xaCjV+l�D	���y�F�i(���	8g	DD���<�y�ɳ}�RI���u�������y��
	�Pl�w�B\&BɊ�	ܬ�yª
UR��E�S�
���$��y��̓(t�=��ā4�d�D�ޱ�y� �E`:�jT�('܌��O��y�Z�4��IB�l��H2C�N��y+݄]��� Ym�ک���Q���!�S�O
���o����K 'Մ͚�'��l��lM�0������h��m��'����ߵ��P�"C@�~�<i��ïS
t�x��E����~�<�烅$;����ŗ�U��2wo�E�<A1,#q�RE�e�؁t�شJ�MN~�<�5�G�en@;q+�>	9X!�m}�<�C��(i�qWo�7u�u�R	Vz�<q�o�1L:����˵H���A�t�<YQ�۳e7��D	_1{yF �@ m�<��!�"#6Q�G׈(��M�ao�i�<�l�t�.ɠo߆d�(`�d�Nz�<���
��&��Kn�跉�}�<��/TOnQ"T�q��BBR#�!�$�@K�ak�˓�]�ȱ�@̰T�!��2_9^ ;a�F<h[LЉ���'>�"��L�+ɲ1��囱a��p)�'E��y2�D�.2�(���Q%3�P���� 4��H��}��{R!>��l�V"O�-�P�D�[u��C1b*���{�"O�1�M�v� т�g�+;�� �V"O$	 ��aڂ����=Ђ B�"O�Ģ�
".�8m+����)�b\��"O@�Ԧ���E�+ݭzD�@�"O�ݡ5K�<E�P����2:qa7"O�`�u+�(����u	X�f�Ա�"O�A�ՄU@��(]���S�"O���S�D�F�9b�'��Z�*E"O��)���&~��bB�� �T�#2"O̴�j��241Jq恷<�0И"O�)�@@�>��@����@�\)c�"O�� �O�{�p���c�z��j4"O���&�4LmӆB�*8j�i��"Or����݃"�P����gĨ@!"O^����o�0�e�Yv�����"O�e`��-fWb%1G/�7_��"T"Ot��%*��qS�9�#�Id� R�"OR��H�8�8�a���M�f���"O�	��)#��\���|�|"d"O���B�,a�x��؁,��u�"Oa:wL�Ȑ����Ĵ�.�y���d�T�oH��#�y��\~D����*b�:ĭ#�y��E�z5v@��MW���WkA �y�	Φ�؉yQo��}�$�foS=�y�]�&E���� �@s$����y���u���"��}��I�)���y玄H0�Zv�Y-�|�3�yrc�'j781xEI׺b���H N�y��X�9+4�欝.a<
d��٣�y�����l1!�T�] B٩��[��y���kB�x�1��!`,��L���yR�c  �cT苠����y�G�25��s�I� ���4�H��y�(��<���{�Gճ���0b����y�_�}_ح�q�� ��L�К�y,�6|�Xz��R�x �����J��y�۲J;��[��]�^�Q�i��y�o�O��D�S�C7u;L�0�y��U�������;qBx��Ś*�y2+N��u��n��I�Ԁ�PybG ���Ɛ+'���5&�\�<���
O��
� ��7Z�lH�JU�<q2o�?9�`�" "5�d�Q��N�<)�&	�)랔���ܹ:�a�`Ht�<飡�/4����6jI%��n�<1�C~|���1tn�Q)Td�<�!�T nE��!ѻP��t��T�<Q�F�t�8������d�5�f�<)7�B��&FazR ���v�<��E�A�����=F�4h���x�<�u�d0�g���-^'^�C�I����f@;$D�M��b�>C�I�qy����H%�m���Oz��C�I���@�G?�����xC�ɶt��di��[�c�P�Z2oã �ZC�ɐ{�QÊӚ5b����B�@[rC�I���h����t��3�A+U^,C�	(-V�[P�6��͡�d��VVC�I�l\:���E=5�����1.G2C�I?V���Ɓ~D>�0�E�X�C�	�j۬|x#aN�M\2!��o	,� C�)� ��s�a=Dh��H3W�(�"O�T"Ĉ$�21j�<H;V�r�"O���c/�<�l��"i�48��"OPQ W+�%xSHY�⊋<A��� "OnȐ�(O2FL���cڋC����u"O hC��OGZ�=B���p��)"O��I�L3h���P��Y�[�{E"Ox�;p�ѣ
��4&,��&N�b"O�(c@��*2:Q)��ƿ|�qɇ"Ot��/[ }_~"�)�3=��qZ"O��K��)�([�Mq����"O�D���$38�`�'6�j��S"O���5�Q'H�h��5�]�5h>-K"O�Hc��>nZ��ʳ�X�g"�3"OLP��)WII��,[�,[{"O~L���_�,u�A��]B��s"O�%�fFD�J��h��a�'K��@A"O�1���jzhM�����T��"O��G�Mo|�ya�*C�J��i�"OB�{�LX���:4�����[�"O ����L/$tE���t���(�"O�@r�D�.��І͌�;k�I�""O���W
��!~)[�[<RS���"O���K#W�, ��	�a5�pj"O-����>T���t)�$\"����"O8����˩V,* Ѝ�yA$� �"O���i@-{��D��+	�8D�Pzv"O��Ɗ�c������]3t@xK"O,Zrn�\���$� z?H�Z�"O�ۣ�ː"���$�G53�2 B%"O�}�v�D/h�+��ߠ3.;!"O�R��MlP�f�!>�m�e"O8� q��)���8p��(Q�؈q�"O�����.3GP0���`����"O�a!�	:5ܰ�PᑻZ�t"OB�)t�vbƜ�B@Ѥ���j2"O�� "�1�H�e��Z{�i�"OԀ2���m���y���"O�Z�NA�2�$�x��Ͼ=&d �"Oh9Bc��m.؈�'Gu@|!p3"O�(�Iw�Hi���a*p(��A6D�kC�Ժd6�#�Ή	^��Ł�'D�4�Gk�'����B�<���2D��q��׌uv� �'ϔ.�M�3D���2 �[��������
1D�C�%�,ZP{�E�z!�`Q�,D�ԪP�O�2��3AL�!�X9��+D���˗�W�`!���H�B��@�+D�$	�/ơa�аRug�'�t�Q(D����>/�� ��`xh�l0D� �G@Lg�� r^�x��1Ao1D�����Y���Z�!lr��p�/D���R#J�?*|dHv
� C2� �B/D�D��E�7�P �e�4j��u:�+/D���S�K5W�4�ZR�� ���6�(D�Q���f_n�e/~F%��h&D����ޣmz�5 ��� �Ҙq1I:D���i[�)y��$E_�K��X
!<D��8 �L>�~�3V Hf�|��#'D���æ��:v�[�!ƄswD�6%T�:�#ܔO�E9Ң���� �"Oʤ��%��&jXpR'P*�8IKc"O<=��/Z�B8�H���S�&uB ӧ"O�8��%k��)&$D�xX4Q0"O� � څ"�\�����ᆺٞ0s�"O���b��(��w�0f�e��"OtIBf�RVH�P&��OO��"O6!9�ObIF@[���B⦁�y�Ⱥ��Xid��>H��0�A�]��y���T�����
�n�6|�� ��yr��!3W��j��Z�]����yb鋮uX��j�BZ�g6!�P��+�y�K�Yu�5QU�A�s���0 
��y��I�.|���E�D4c��A�E2�y2��41x����̸\�z�S�'�y�怭0�~��g���AHN�1����y"��7i��ITlڅ:�`��3$���yr,�n�l{�&�4ڪa����y�Ā
(��9ya�P�0�9�u�'�y�ۗ:��;F�V�3 (P�+E:�y�Y���RnY�*fl����y�V?')
A���@�D\Q��I���yR -b�X��K;�JUX K�y�+�MO��jr���$�/��y��;g��8���J�MP��F*�yҧ�RۄAY�G-H����+�/�yB���:=���q��8�Ń��y�耀>�1�'LǠpe��hX�y�$@|�sFh��ѓA��yg�`���ZKJ]O�����y�i�4D*:u��)�"M�v�j���7�y�E�)<�TmbNܵ.ɾ4���5�yr 5Π�q�nJ�#��Q�Py"a3�N�i�#�mn� ��J�<GI�* 5�y��F�p�����C�<1�U�����'�H�aʕw�<�e���}M�����A$Pʑ��Cq�<Q��ץ^�L5�'a�<���l�<Ѵ�G�K���Z��N�s�2�cgc�<I�G�p�d���.=N�#��t�<)t�	?PL ���(�<`�D�Es�<Y�E@�x�^	�UKҌ�`�B��E�<�S�J	B��Cg�
6��	����B�<1��P���"d+nt2a�]|�<��I���؈�Oۦ:���A�|�<�� W\���#Ǌסg����E��v�<aÁT�0z�� P
q�81Ӥq�<1�dF
|p��p*Ŕq�n,Y�a�w�<Q�)��(t�WeO�jw�)�g�\�<�t,�
p|҉���D�4Z�U��Z�<��C
�tl���ě9	`���QW�<9�&%Qm��Xn�x���S�<)�)�6j&�*���zP����N�<	��R� H��ӫpA�uXeęS�<���4a�ebE%	���ˆ�Q�<�#��*) �k�g^&=����.�F�<u� �Qp���c� S�:���C@�<���ru�yY�Ƒ�@�K�&u�C�	 6�k�L����i�C�O�C䉔q���!�Fͭa7�,�OދHC�I�uV���˲hd��
H<>�,C�
|�A��Tpb��Eż�@C���!�G�>q f�(�p�jB�	�R�`dBC�	�O�nX��.�v˜C�<�n)*S.3-���	@��^?PB�I3=uR���E��hn:����S��C䉨$��Y�4@X�� z�"G2B�|�.%�C�C&l���Z��N���C�)� �䢓EQ?���26gM�HH�� "O���dƆ|_�y�Te
;_1n|!q"O�WK/q��Ǝp�l QJr�<)��:t�c��L�.�D$�DD�<�Ս�;	�~,R�Ɲ	k��K�g�[�<q�Oٲ3�$HI�!BD;����<7$�)*��-��Y�+�<�2�KA�<!��Z$*�k�>l�b�9P,R@�<�MA�~n;s�f|B�C�IWx�<!�G)+a������1AѶU�K�t�<����z�Le� .)qU^�2��Cu�<�a˓ 
j���`m����_{�<�c�27�P�����0s���BI�q�<�Q���J[,��aŝ�uΖ�[��l�<�6�L��,m0w��X�VYyF�~�<9$KAO jPhPoЦ��Dq�P�<9ݼ1��c�� Y<�ts�#C�<9�hӹF�����&HN�)&��u�<�3k�R#���ߟv��M{#B@g�<��O�eB����]&aYT�RU��f�<���(}F�r��C&	�8`���z�<IS��08&tb�e�EM��ɧCN`�<q�m��Yk��z��@}��8JU�_�<�+��6r��"�T�����]�<q���#�'��3�<�T�HW�<Qf�R�@}X���nF�@൐�`MU�<��I�;G�� �J3a��P��H�f�<	��=1]LԠpׯU�,p罞!�䕫P��hC(ٜ%��ɰ��)�!�D�W=��R�@_�QT��XU�)�!�dG��¦������Q�	�!�_�|P\�BD�C���@�)ʲ)�!��^8�i!@ f΁"¥	c!�$
�� �A�ŏlX�Yp��,#!���0=`���&͝;S.m�Dd��I!�� k���kP�"�r����>.�!�$V
ž��dn0>\���!�)V�!�D�,)�hHT�Ϧd@��jbY R�!�t�~H�c+��2v�jf��}�!��A�T��)U�B�*��9H�����!��Y"Kt�ר�+u����ϙ�yn��$��<s���=DpZӆ-]:�y2��^8�u��W?%���q�]��y�
-��r���"v*$h��ɛ�y2Ň�|�RL $����� Y��yBm��8p襑sl��h�����I�y�g[<���Sk�>deh��B��y2OH�X�: �U��%[���(�y�Ʌ��t�۲)�*Z��0;�#Ʊ�y��O1I �IơFM1� ��߯�yB��<����$�Da����y�T=��y{�Ǘ�D�BF��y"�5 ����� 	t��83�I��yb�� �N�.��	����"�ڳ�y��+����c�$q>~z��X9�y#N�]zQB*jC$��'
7�y'O.
�#�
�c�=��	7�y�2�t����X��wg���y"���	,@uR���N�HL�qE]!�y"��~v�� f�R�oh(	�h�$�y�o�u��H'
2� �	�'�0�y�@�o���K��0yb��(B%ަ�y��X4J��d픤({�!1�K�y" K�dy��seҞU�n-ÓO!�y
� lQ��݊�ʨ�v�֠@��m�"O������'�P%�%DD�o!����"O�Ź�8MG�$��"V;<@�"Of�r�䒫�l�e��G;0ɑ"O~Pj�%iwP��@��(� ��I��P]����i����AsV�Ұ.�<`y1�[>������O�h[����S�huiŤG@`˳� >���JJ"���0g-JFײ!:sD��HOdk&�X�L>$�'9Y��9H����T:��G��G���*W�3X�4A�%AޤK��̓ti�O��$������F�oN�i�Z����b���4+0A���!�i>�$���'���xV�Q�0�zN��I8�@�Û&/fӠ6�	�U�|��-Y�t�d ��FS�P`ݴ'���"3R�ܖ'���O�'�'���z21iC�\>EB�ʁ�ɑGC�ć�&VM�3�X6,�J�i���Ͽ{��Ko���$�L�;����l�ʦ�E� C�����x������w~A�t@�4{�1�k�L�dK�(ɢ̈*%� 1 �	s��L	��?A��in6��O�#~n�-
G�eQ�������#��| ��ß��'ayb����ȴ��[?�	�%E�HO�7���'�(�O.�rhQ�F2��*E�ʘ]�HQr'A�<�Co�7(k�v�'̈�{C���@�*S��@K� �D �(0	P����X�F�2k̊��ψ�O ti�i������;,ޖt��N_�� 0P�+KLV��q�D�!���ڦ���g�ɽg������7a~���T>s��k�(+
!H�aݛfI�t�,O��ķ>1g��v���To���%��A�h�<!�  2DÔ�^�~�Ǡ�,#�� ��a���oZ_�	�����<A�����0Q)��?��BcωG#���E�_���<I�GpDX�� �h�)J<1�|��CÛ#�  `pN�C�H: ꋝ[R�"?�%&��Aʖ�#D �d�Xxap��;M�m�c��3r�~�A�,I<gd��ѦF�Fx�!�?�۴Px0�#�����Y�T�X8�jPlD��͟\�	[�IF�S1�~��P�I�A����$G���IE؟Ԓ,A�.T��[Æ�*,a��r�A��?�Ҵi���'B7-B��mZ�t���[b�Q
i�t�5���q��a��B�B��?y���
�L���:c>�Tb�)�#%�擩X:����,R7H<��EOr!�#=hX�{�
�FR2/JV��s����u�'��-�U��.-Ԁ�b�se��	!l]p�d�O���	E�����T��V%S�	�d�7�H�eά�D6�i>�Fzr�8��Q�ʕ_ �8W����p>y��i��7�wӆH�ьW�O��6�F�D�����Oi�7����	Qyʟ�O%Q�&��M���4d>�5aTk4 ��caH9j�����P
q���x����W蔻Mv6y@�E�o� ��k���M3�O�=�tH�c��OC��{S���@��̻��e�����X�Uƌ@��H	�f��x��˦;���ON��_y�����V��?�8�I��+Md8����~"�'�azR�O`{�䎖%Wj'<):Ф�M�Q�4*�4(���|��O���ʿYP�t��Z3vJ�(�LT� ��4'��퉏e~p   �   9   Ĵ���	��Z�:tID:,���3��H��R�
O�ظ2�x�I[#��C�4e��B��.�=H�n�,��x�$�#f?V6͂���H�4;p�1��\�I�$U
E9�`[*P��2A
��l�tD�UE/�7�T#<)�&i�Z%��MX�J���$[���DX���'e �jm�,6?i��K) ��6Mp}"��t�Lc��&q�N�3�jAg� ��
ry�.�OB�6d����9On��$J�)Q����Qa�dL"D�#
(6 ̋v�H���D�==�������'���D$�q��Ȫ�`����H(��%����3##�'(����Ð�> ub$��T�M��'��Exr`X^�'��E.��!���Y�P����(N.#<���>ѧ*�4e@>a����Ty�F.r��)�O�ڊ{@�Y�V-;��ΠZ�<K��F�Ms3�-}n�"<��/�G�ld"sf�|e�Z0�E9Z�p�>�Vn)�n�4�t�xEY�(۵#H��U%��0�� �'(��Fxbn��nfR�� 7{x��K��Y�0վ�a�:$"2#<���Ox�$��q�E���6[�ٱ���OB�8I<Yf�;t5���Q�I^��p��ZS?Q8�\�OR�I0K��p�"�Q�Љ�ޢ4�.���h~r��97�]��4*��ɏ1qࡉ��OT�qakHn��SӨ��
,MɁ���H��܄N�Q�����>%f߷&.T���	 ���3ǄI}R��j�'ѪGxr�H�s�NS;2F�� �%�y�n�J�  �O���Q��U"�GUy�Ne�
�OȔi�)��8�L�)�A�2�"�����Y��M�@����nD
V������)��3� ��w�?.��E�d���V�>ŉ&͚0�?A��:���<�'�?���?9 '�!1r`hlA:���`�O6�?i���ċ�	����۟ ��̟P�O� ��F���ӈ���t}��OJ��']p7����O<�O76��U��v�>e"i�%cLY�c�aA��4��(�� �̒O����>A�#��19�B)(3��OX���O����O1��ʓY��O�=�0��E�F�;!&��em)C���*�_�H��4��'-&��M� �z!��C�	����yZ����a��od��Y�a�|Ӿ�|#�틆I����O�Zc���p��@x�`�:By
�h�'~�Iß����	����IV���3e�4�I�#���@�syB6-ջZ!    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �   C   Ĵ���	��Z�Zviʗ&���3��H�I�
O�ظ2�x�I[#�<��4d�v�V��$�s�ի-h�K�GЃi^7-ƦR�4WU��!��U��) ��|�t�G�,�B�Bc"�3���uH4�,��"<�hӐ ��g�
8��b2�Yo�p��X�`���gxN�Ѣ�*?�W L0
7m
P}R,l��)s�R�9��\�S#Y%B���k\6��aqB�X�i�JC�x�+��,�k�
�tj���@-Y�x�eӋ��F�� �'��5�����'r�[%C�^:�nڠ"S��PM�p�Z�Y�ǁO�(�O�����$����u+��
��$ӬqU��-�Pp��"<���>�]B-�S%ۻ[/�,���К�M��I�)�����Z��20���3j{AM�3�8�� K4}��e�'���=�LB[|��L�-,��A' �⦵��I����!m��o7����R�ԅ1�Q�1b�0y$�	7&p���m�j����ؿW��@�GJL�T��˓��"<)� �	�f�z���@<i 4���	��i��ɮ52���E�'��Г'&թ]
9r�ږ!����yRi�'�J�$�T�7;%f�;�j��T]�aX�����2S�ɄZ��'�f�ɱ0�\P�+x��f��O6���~~B5xt�l��4��	S4�x2�O�T0B��@<L֘aI�ߧp�ڑ��Y�T������c�X��Q� `�'ApE� \E/�|� ��[�X��O�)���䃼�OHt�c`A�M�����E	'Ӕ�S�'�@ �����d�5�?�!\���ɬ��ˣ��&�F%�P�l�L�������/Q�
�B�{yԠ��ĳ?��'�de����;;ب8@�J4�|��'�I� �I�������0��w�4��e����倗>�Bh��J-
6��B����O��$)���O�]mz�IBɆF�
�{��̧L���Ċ�����z�)�S)G����b�$��ԜTDi�G�x��@���h��IE�В��$+�ĩ<����?!��1-����� E9D�	�7���?��?A����$���2U�C۟��	�hh2��^��p��0c�*a�n�D��3P�	ޟ��	p�)� (���̔�4Bx����$�5�g�����ƤXw�QbV�W� Xs���O �(wNҊr_�AQ�٤�r�t��O����O���O��}���<�F�@�kͫn'�J��3p�y�����֠Q    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �   F   Ĵ���	��Z �t��8-���3��H��R�
O�ظ2�x�I[#��q�4�?iU/�+SM�	�pMW�0�h<@P�\���j�6Xoک�yb�$6��[EBhR e���B!N�v�9R��Gu�p�i�vu�o�/�z)���&pF��'�DA�.I�$�*O0|B�99#61X��9��ϥ�̘2���5f̴ �PBP<Z@_�L͓Ooք��Jʻ�ē%ha0P8y�l�3��y�D|�4�%^�態wH�<)�k�����&�����nu���_��YX!�+)
�˲%S�?4`g�5��L�OH��O>	�/�o��z�&Qg@�:�V�<J!i �"<q4m�fWd�G�Nz�<�#�����̻��I�y��əR����5e�9J��,Ӑ-�ۄ�'k0Fx�a�Y�)��	0&Q	t�3(_�,lnڭ:��X���I6kH)2�����FG	��Ȥ���/�I2� K����P�L�L�XɆKǺ2��5`%��<�e�$�R�4KԄ��_��lb�l��P�������D���a�	%}��G�9wH|�,I^�ܬ������'%�PGx2�Dd≋wD�{�Ȗ|.5�q��	�EI��D�xrn��� CIJ�G�n����N=��(��o�O��'De�aߌ�M����9��Ҕ~+�ŉ�}��Fi�F�Ƀ���.�剄��I�1��L>���'�xb��<=�`/ݤ3*�������N��O��1�����
@o��d�x���R/!�$��#� �  ��O����<�O��c �ۜ^Fe�0��b��Pa�zӮ��g.�S�1O>�	�n,�E�Ր
thaäj�!pt��Pٴ�?���y�FGh)�O����PR��T��ŃKզ�Y�&I!lO�$�OB�dv<��s�CW�X�"z��O$H���o���`I\�ē�?������f	<#9�gcH�F���AQe�o}��U"��'v��'t^�LRC�){��U�Vn8�eA�Z�(�J<Y��?�N>Q���?�ebD�&�z����B6���
r�z��<���?����?)�O�ܠ0�Oތ��FƋKL�PQ.J*#��ݴ�?i���?�M>a��?At�J�C]B�l��Z'b�ru'[�f@R��/��|ꓥ?���?/On@B��J�D�'+bU��Oތ�8��.L�HD[RdӢ���O0�H��7�I��������`J     �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �   A   Ĵ���	��Z�ZvIJ(���3��H�I�
O�ظ2�x�I[#���ݴjk��&ֺ+�j��'$[=Y�"�a��<EV7�����4=�$>��E�	�!��l��d,)���Q^�(p��J2q��"<Y7nh��(��+S�@}�U�A��P� �3+��@8l^hy��ćayL���D(��D;W�,��H���R͡�@7`���0����D���/R�-&��r�ʛ�*W�����E�Op���G�V�~ ��|2!��'�pd�K>A��� �� ������0�OaZ\�Qe��M{�D�'��ò"�i�'��d%��o�ܺ��
C�\������yҸn��hd�� Vl���� D��2�"S��]���$
<�O�Ey�O����K�$L*{�	>0�T[��>���,�u;`�`��R��V�r���/�c�d�l\��d��O�MH�f�@[���nҼ6�$�ע�<�O�������$j���J�~&��ѫ��\��!*��p3��Ċ�f�.%�؄���q��8C_RY���T��O���E׶����Q����4k�%����<3�<�c�O�L�0�|��Q�  �L��Q�OV�ۉ���
�����ѥkdtMi��2�� y0H�ZPr�WUy�d%F1fA��4���W�\ɩ��Of�ٓ� /G�dأ�L`eh�qS���/��1Y��O���Ư�=A�'�8�y��"���1�/��U��O�9���_��O� V����D��,۩E��+�"O�q���  �  �"O<�iea�F�8x���-?��k�"O 90�
�(O\x@��D�Hks"O�虷�K�?�|�/E�b�0D��"Oz�:�a�$���{���T��t�Q"OjxP�Ł�a@�c�1y_��0�"O���C�Ι0���p�ၑ==	�"Ox\��AT�tQ́@7�7i6���"O�)�RKD�SK=Q�	
��p�"Oި��k�2"G�p�vZ:u�f]�"O�m�F�ܙn�@[���,��Qd"O�0,]��Em�)���Ӣ.D�D�r(C�D}��ɘ8QG�e"B��o1n�{�)��]������00*B�I�/�Rq�X!_��mawɞ0k�C�	8����W�������G	S\~C�ɻ9���Q�aG�Q�%�6G�$�<B�ɒb<�� à5�Vye�8B�	�Js�M'�ef��`-�' HB��wD�p%��6 c\���C�	�4ìLja�M5z���/ �L�C�3i �� *݄8��q�Q��0��C�	��q!Dȟ�
v��H��r�rB�	M�h�Ǎr⒬���)T�B�	�^�:�J���Qt4�#�R�|B�I�^7��teY�]�b\�Nsj�C��kP�@@,R yh8C��:]_zC�=)L���I�0AyX4��*ޫ�NC�)� ���@�ܑ��â#6�2�`�"Oj8�d��R페@6��dXB�"O�M�`E0�l@�J�d� "O���4
�:ʌ��AN�'�Q�"O�����7k6��ʇ��x��q"O��3� �GS�U)�oCYy�TrU"O��b�-2]�	�0�7re�s"Op�j"$��<�F�R��13T|��"O�<�Q���4V�P���P���"O0H��Ih@�rb�>oN����"OL��.�= ��t
�730�}�"Oj�[���{wx���0D
L�2"OzqC��/:�(਱�7` ��"O�XG��-�<5 FB�%gc��ks"O�4%"�?
�$��!�ULX��"O�Œp"��xPRC��1o9����"O���u	ҙE��a��
�9.\�f"O��(�[�NKV1�Ώ�62�[�"O�Lb�a� _;R�{W/�g�HĪ�"O>l��Y"el@�$�&aʮ(�S"O"d9N��0�*���㟴���Q"O4$s�;N��ɻgCރQr��A"O�1� |$Lu�g��;3``S"O��!r�3HVl�J$]���i�"O�񀐍X�kz��n�!�,��"O��N�3�Ġc�]�ov�s�"O>�!��B#㦉����-/B�e#S"O(Bnۛr/�c�a�1.��"O�S��רk��	�2.���0"O��2Vc�!f,�ŪH�&|�)[�"O�q��۠%
ƀR�A��L2���"O��cj>-��3� ףN��k�"On����0�-��i�4)�"O����� M�L�M�2H����"O^ ��΀�����	
!&^J!�"OH,1Ѯ���F@`�EP�)�Z#"Oܤ�U�\�O(��Ņ�&hj�kD"O�Y�M���t{���!:hx��"O�� �␎K\ �f�Z*&�N�S"O��J�,�?�4q��A����8"Ohqc�S�^���`W?d�$"O�x�����O� ١���]���"O�HeB])�6題|M2�)E"O��
U���<3�`:
�+/(4�D"O�|�weǼ9r)����A|r���"O�U�fo��
���c+�o����"O2���mUy&��R� :q���3�"O�pp�#r���E�9,戣�"O��	4͏�1/$�Q�HסW��A7"OH�x2G�RF�zH��kn٪�"OJ\�7*��&�6<���!#�t��""O�$3�OF�{Q8������t�H�is"Od���k�
vX��6/D�v��Tk""O�x�P�?kҶ��d$�7�tYt"O P歃�t�X"�?+�R��"O��[RM��"Y��$�ɉ*�p"O���x�۔)�w`�]5"O$�KqOP&<
�B��	DXq;�"OJ��U�rpNp�I��<�m8�"O� ���A��� �1ba���[�y�䂁)�.�8�&��Y(�� ���$�y���CT�rD'��
}�qG3�yR�
I�s�
�|���¥H�y��	:"/�,�$C���@ƢG�y
� ��C��ĸ,���0(E1
`41 "Ox�C��:%j<m2���;$�
W"O�XC	���9p
DZ�h�t"O���Nz��]2B)�q
��s"O�3�j�SԾt��g�D��9;G"O���!0ڨ�{�EƂGڒu��"O�%���Q*[���n*݂�#5"Of�p�?�4�A���>�P��f"O�a�` �BJ<Ժ��2�K�*�yrc�]��@�!�CLO5�N5�yn�NKF���)W2i�jW��?�yB)�3���a5��3"���Q��L��y2��6Ks��agH��T� �)�y��%S4 ��BhpՈ
�yB&K��`�V�G~�Eߨ�y���Ju���/ܧS^��Y�.�y"�����������g	֊�ybۖ(cda����:s������y��, vy٣gŴ�BD��cS��y2@�D���m�Z�+w$���yr&�(<�HؕF]?R� )7-��y�o����i���B�6@�*&I��(O6����_�^��F�S
��s�jG3G!��REIv S,�>5͐�P6ʕ�9!�č?E�|�WjW��vD�b/�� *铨�>!f�_*��-�čD/K�8��U��C���!�����A�l ؜��)K'-��eK��:D�4�qṀ;A���`�
�s�<]���3�Vb�D���l�(q	 E�${�,����y��˫B8��5��<"��r!��y���>8��W�7ޚɃC��=�y��4��`P��߅'p%Ȃ�� �y�, 
SÌ! �I2�� ��yb%�����*���(2k٫�y��Tl1�A��}� ���G_7�y��΋*-��Y�HEGX��Ј�yl��k��X!�!��:�^�!@Ԑ�y≓7X2`��7�`��JI�yr���}�Q����e�:	��<�yH;z�< ђK���|�ae΃�y�j�����"HL�����1B�=E���X�RD�����L��X���z*ȇ�[�8[W�E��V��g��\ 0�ȓ[!6JB[�iq�ԣP-ˣk�:̈́ȓ/���gZ�V�p��a�H}6B�	=}�͙���p[��a�bB]B���>�H>9P#�' 乹!�3*^h�r��f�<ф�ٹ3��=��M���|��O�L�<��/Ϡ:�rp�peY�
�� �H�<Y��B�pM�uPHL�Z��M�`��\�<��2�e�!j1:0��&�>Ii!�Ğ<	�.�P$O�6,0��C��0Z!�$��8Q��A�'��M��vH!�RQ� �P�ƛ`�����FWU!�Da��oӷaq��&.��*J�Q"E"O&�Z�	X�_X80��N�*6�,�"O�͉������M �h�T����"O�U�T�S8v"�H��C�S��33"OD�����;|n(�!�'V�(�u�$"O�T¤�ŜH�H��a����!�"OdC���kǠ٪S��
��s"O�b%G��|t���i�l�B"O(�`(`-�QѕaP�:#�1""Or��p��*��u��Y�u&���"O� �YE*�2�X�*F�Hl�*��"O(�
��ªS4`B劇��1J "O�Q�'���ޘ���ʫ[���2�"O*���	&7��E2�q�� D�4��)ͧ0Aj�zgG���͋�1D���U㐶�
}��R"O�es�@.D�8���E�G>b-�%ύ=ahA+B0D���e�Դ`�h��P�0{I�{�	0D�h���[ ��ZƆr�fQ��#D�d����FB<�1���w�2e��C'�􈟸%�2�<�� ��,wi�Q8'"O�!K�\O�u�AB�T���"O88���=a i�b]�zQ��G"O����_���0@ŒjJrTk�"O���0K�����$��+���'"O(}k�L%3���h��ք2�"O
����̔Ȁ�Ѷf"K���8G"O6��g��U]� �F��HjV1i"O��g@w�(���GT����x�"O�Tb�hV;.�����+f�Z�q�"O*��7K� ���N��C$"OB��P�@:k,Ը��Ԝoh����"O�\6&#T��TP�x�ܠAe"O�%caE8XY��4n6e�2��D"O����aFA@|�7#:� � �"O:`�C�
@�R�ʢ�
5Ӡ�:��'$qOZ���n]�]�U���64�0��"O�P��L>M6�8b�P����C""O�49w)���Y�p"����!"O
i�dH��z Z�Z� �6� ���"OШ���:�@����B�C����"Ob́��QgZ]Ҵ��� ��"O�xCMڧ`�@x(��B:W}(ɊS"Orp�<v1ΌK��P�ko�U��"O�0�h��G�̳��(ø��"Oj��$��e��)��̺e��A�w"O���SL��#�m�d�\=���8�"O~Q�%���d�%�Sd�0��W"O9���=+D1�r�Y=7o���b"O��ࣄ�5	�0��	~��aU"Oֽ3 ���z��#<����"O�đ��ξL���j ǖ�S��8�"O�سU�lܠmHw 
���b�"O�0��i�I�n�7ŀ}���I�"OԴ�5�5�`0�aD�S"��2"O�,; :IP���+Qr�*O�����7'h!#�W�l:���'����ȷ_��Ih�MI&b�b�Q�'�Rl�t��,N�PA���D�nՋ�'��h�I��8���0�N�?����'���%��@�d�W��H�Ȭa
�'�X�:��߄����C�4>��x	�'l>�P#�V�6�q�S):�Д��'���s���M��a�@�~]~H��'�����e\Z 2��'*A�h��';,h�#��;�6�zЊމJU�� �'���ۦ���lȉ'�F2H_�4��'`m����{�M���Z8:��Q�'��lZբ�U+HcD�(:����'���D���M��!˳㉯�����'�ڽ��b��&LZ�k	�b��'�>�i4E\�Zid�P�Ǖ����
�'M���ł 2%��� _.,��'[���r	�3ߴtA얬\�t���� �5�HW37G�y� ��<AF"On�	$K*.n�S`n���<���"O��+��ƺ����#@���"O�tS4@҄R����֢Ąe����"O�xĎL�wb���2GշM���`"O���a-�#"��-HC��J�b�R�"O�%;�&֜!��Tsw	ʃO��3"OL�b�^�5�ٲ�(Q��T�(1"OR ��Wh�) M׏@�
d*A"OxM	�HK��Yu���F�(�"OJ��
(i�̬�G�U&`7
b�"ON�9���
@4*�%����"O���%���"�(X�Y�k"OF�aA�V�n�jx�G�+,����"Oޠ�W��3$�� ��;@�
1 "OJ�VÂ=Ft��Rb��cj�:D"Ox��7�^�"�q#M1�t�f"O��CdX�O
j�A�{ (3u"OP@�S��*�|���oJ�VQ�!S"Of<���F��f�a�]�/;�( "Oz����V�[Wz�ϝ�:����"O�P"�ͷ~��	K�`�!Yb��"OnDR"o��$�m
���8���"O^I��Ь}⁮;�X""O�Y��J&n��ٵ�ɭaj��"O��)dj�1/(F�8q؂�,"�"Oi�t�O$�<u�կ]�T��Q�f"O0 (����U�(�� E	R����g"O���֪a��!j�i��	{T%��"O�F��)���A��Ra^���"O�8����-o���B"
D�^U"OT�TM�,&�(�LU�љw"OP�pu+�4R�T�S�A'C- R"O��� ��7c|qk&�R�b/��"O@XY�,�!g��1\�9��I'�yROL�F51�ÞZ��i�#�ݛ�yR��+eT@9"�`��4 �m��y�AW�M�f�`��:<Pá޷�y�#��<kX�)�D�.)�>���]7�y��X�+i���@�'&�`B��J��y��ɨI@�-����dv�� W�yrE_ ,!�Aa�HO���x[�e��y���Qd`4P����ea��y�9�� �g�6���b���yҢԸ_���,ٴ4*��LK��yB��_��x���TqB��O���yR���X�A�dҵA� g���yR��%)|r�1���n "i�����y�a �v*�PdD3Z,������y�lٕ;���j���"�
=�wB�3�y2ÙN���+E�0�\&��	�yb���K��H��FT	*!^-Pf���y�*ӻ2��p�/ε@�Ɂr'_�y2#�^��@{��@�pQp���y¬�6�(g��x-`Ur����y"�I2����DtA�Da� X��y"�K�
��͸g��j8a����y���mJD���'d��E�cd�<�y��
�~��q#T�U� ��ӯ[��y�B��_�ހ!S�$;�0��#`\��ymBQe,$���U 4��a �����y���X(�\�����(�,mB'o���yR�,a��]s���v�['��:�yBj�(V/�%0У�K�t�y
� *	)F��(d��p�A��J�@D{r"O4��j�8YC������c!��"O"��� �%�Ȫ��Z��q"O|5���h� ��#c&�a�"O��0��� `?J� "�ѷx�s%"O����_�@h��0W��N��\
V"O�<���Dtj�`Ɓ��Ai�"O�܁q'�.:p�a����~�ցk%"O����ܲ)01L�'y�p�Q"O�p�RKV`��9CP�Çn^|�R�"OF0�7#zmZ�,M���a�"O�Պ3��"�6�q��O�I�1z�"Or0xe�W9.�����xÈ��"OI���?I��4Ӵ	E3O����1"O�=҅
�2�"v�V�OuR`s$"O:1�n�T6ʘ���c,܈�"Ot��a�O�>�Vaj��WbO^�� "Oʌ� a���,��%W�����y��G'O���G�)o�}�!�D�y献Ae9IW�Ϸx��@rE��y�,ֿ+pT�p���p>��1�S7�y'�#/��rDjR�?j�������yR�ޒa�؅�H�!�L�����yRBM�Yh��{囂�z�B*�5�yR��(7����Q�g�~ J ��y"-�C|ؑK6m�P�ے&ت�yB���Kh��iH|�t�P���y��U�Ҙ�e�oG|4R����y2�D�K�T�r`��c̘�&)N��yBG��?�"M!'�כ[1X��e(��yR�_�f������M|6I#����y"솽H�	Q��J�7L6�Sa�\;�y"·8	uhذ0��\L��˻�y��فsL�1��G�O�ԁH��ũ�yr����;�ܝE|������yrϟ�wI���"�!(?P9��
=�y�+G	W^qѢ�P>�x��L^��y���9�,�[���+Y��l�R�'�yR�*E��y �h���h��]��y���>t��	��%�D�kO�y�Bۃ%2�a�-�6x�f�a���y�fA�YSȕ���r>�|Б�ݽ�yRO�FL����P�=>�A����y2�](Y���jA-�>@�i�G��ybJ�&���Q�֫=�F�'��y��D9%���x'���.�dAF�)�y�+�9e&��(�.��e����yr�6����hT9O�`W�е�y�
�>=�60����)%0Ijv	Q$�y"� Gת	Z�c�(v�I��g���y�F�)���@j"J,�{*Q��yҨ՗S)�=���6h�.�y�@��A���Aa1�����y��+f����.��4T��g_��Py���"E��SG��
��Ɏq�<�6f�%(��"Ň�0V��U��V�<9�[
#?�a�� �-$8֑ pHy�<�1Ϛ�1�-Vv'p��E�8D�L�U,��r6|iqa�ҁX�Z<��j*D�B%�C'-����"�	u�	�4'$D�X!���<	 p*���2Y��D��>D���G-��Q��U<ڸ� �:D�X�#�E�|��su�s�LP��9D�kwA!#�9"�ʰ7S�@��9D�� �xs��N�48b��p]`<:t��"O:��e��0��P�S�FJ�"O��Y���3]���E�3Z��j"Of y���&�t�A�?NC�@s��'��$K*&>a��`s���&�)r�!���(5!IX�����Ы@��O:�=���T��,I>	�1p��	��,j4"OD���@5$��<��ƀa�v4��"O���b̛����xbeܻ(3��c`"O�@q�Y�;�J�`Dװ�d �"O��)U%@9�ԊAC�9I��	�"OR �f� 5����:C�AA�"O��RӏG�z0(`�I<:0�	�@Q�h����i����/O�&�
\9�mC"9�C�ɧ\
�Mic	M� 0q�v̀Q�C�ɬxZ<�c�f���z����B�	!D�MYP`_>#&-����'I%��O���!LO��Y��}�<L���x�� 9�"O�tq�M3�.�:F͖�"����"O�� ����L�4H
0g7J��|2�'�I���:X	���5�^D^�Y�'o,x���:!��UJEj�����'���ۀ@9(5�
�BF���y�O�M���p��%��F����'�az�U����`ݟr4�-Y���yR���-R��7i�<B�`˟�y/�<Y��J�%
+a���aN-�y�L$}]�X $u��Rh��yB�	?C���G5O	�<��&�Py2�^(�����$zH �6�_t�<y�_�XUn	ib�����p�.�r�� �ɹdt���`�JpA�i��"J� ��jF��{DOY�G�����k�,ȆȓD��@�@�!�<��G�T�5`��ȓW�aÄ\�h�l��gkM�l��=��^Yʕ0��5�$A
1��^?��ȓP�@�f���wHdb5�%>���Dm�HW�˛UeL�"Å %5�� ��W4.�c��W�<�.$	�&��U�$i�ȓA�u��������AK�+ ��'��D{��Tcd��	��\1�.�t����y�J��`��6Pp�հ�y��R�e1HHc���-�,lY`-�y��K�#}�!d��<<�a4m��y"��+ ���!p����=ғb�	�y��B�g �Bq��'c$���X$�y�U	H�,i��Fºc!T�jC��<A�����P���Lد$!�8���3LoV�OL�=�}2�-ʬ~D�R�� Kl�$�I��<��E�\_`%�'l,���D�<�W�ZJ�����#CyT�zd|�<Y��O'c� R�lãf�\\��Ba�<	�͚Y�Pӣ"*e�tC���G��4�<�D"��Xʬ�S�R�$����	A��T���OP�Tz���"K�-��!�%��q����5�b�� DD1��i7MR�E]:\�R"O�����_�!N(@f�PQ�t�R�"OH�QB�6zϔE�#i[�d�"O�а!�yM�p��փo��8��"O�+�6'Hā��"O{��C"O��a��5Zr�M����ٸ)��"O.�(TeW?���'�4��1��Io>���2$�f�V%K=kZ�ukSG7D����G�$.��sɈ!sU�e��:D�� �]��	�e��b�@ǻs���:�"OF�ʧ�ٿf�x��V�	
f�"ݠ%"O�Qi�H�@���)!���2�L��џ|��'[�h E�=G~��*� �BT��'�&PcD*�wB�I����w0��ڎ��7�X��j�_�6�I�!R�5~@P�A"O��	�`�4%?t1"�n	r�L1�p"O�U��D]�e���&C # �����"O�%;�`O??&ı�g��`M�I�B"O^���ʇ��KS�\%��id"O���Ai�z�8s�d��\�"O��@�
)U��
*@���t��U�O!ʵZ�`QR�n���!�� �.O���7f�^*�C����T�1 �f�!��B]+��Krt�ݪE�!�d �t���@ /��!���I� �!�d6��8�]�3�@#�K�XG!�D�M/�u9d�V�O��!��Y#�!��-v�$u$'I��E�5	O%n��'�ўb?�X�b�M�>L��"ִxV��g\����I3I� ;�9o,#V�pfC�+&WȠ0��PL R�r&�8
�C�ɉ^!h�P�M ADؠ�BP�C��B�ɬ%n�9���>2X�q�N	"RB�I�1�Z̢��H�mlTC�
�&\ B�	�_$P u��>`H rDG��bB�ɂV��q�2�F"6���"�)��C�ɰ �j@�	�	7��YHr�9$�`B�	!S��6����&A�p�@�m�2�=��'@����l�zL9�E�B;`���FR�����@-F�tٱ4�V<�܆�wv��WJ�4�����̺Z��0�ȓW��TJ�		�JSd��R�R���ȓgE�x�dX a��-��P8$��=�ȓ~���aea�������1^��ȓQ'$�kҨ0(rd�ThZ����ȓ����1������Ŧ��ȇ�B+�1ah s�b�H�`ӭPJb��?��,��q��B!N�@x�ç/Q���ȓX���I�2���X�&Zeȇ�;9��R�C�@�Tp��g�b��|�"�)D�J�)^,q)����`B䉗nY�8i�+ɋ7�
a�C�{�|C��/kG*�� h�B���:nZ@C�	=*���4iy ��	PHӍk �O���D<�z�9�+\�-A��q�(�ў���	�z��ar�ǄS~���smJ�\�8C�	h\ Ku(W�L�H�����.�C䉘N����[�[y,�HrK��r�C䉲W�ٕ���u1@d1�(� x�B�I�`�CV�V�6X� �7D�D�zB�ɇ��-+��?bM� �Xq@`5j���'��`o�<�4�rŤ���ۈB�)�df�Me@��c�'"������'��'+��'9
�0:`�D=���!>!��V�g`0#���-�,��F�9-]!�$�*@�nUa�fX#͌�x�&�%!�D�7������1`���d <!�d4e�4�R+ʕP�1�6���)!�d�
ir�����˙&BdMS���)K�'bў�>��N�z�`4�2"�x):��A�Ic�O�"H��K�	70����CF���'rN��a*FS���؆dX�'��U�g�A&Z�x��7c�<������ �X�so�sd�)%@$i8�X��'����0����#ԉv��x�u�X�]�!򤋞y��A6J�)�P!`�C�1em!��Y���#c�_�TH��o�<�5O�����=,�Z��v�xq�"O���@V�J/��1+�>�TB!"O,�!�
π|�.� Ӓd�X���"O��ʤ뜬UT���cE�N�`I���'�1O��qBӯ(�՚XY&����ៀ�'�ɧ��N�"�
��H���w
��/��-<D��١� ?�����f�	�G�44����C^�"o� �'�R� 3��b�<�#]�����_Y��RP��Z�<9��1J.�q��"��C!z�#a�*D�|����7 9���b��40���1eg)��䓹?�ʟ������P���@&�f1���S�XG{��i�U�Ddc�T�j�D�b����*D!�D�4��JcG�..i� ��34!��D�� aAʖ�(V�K�CB�9�!�DQ� F�$�c
�5
6��S�@6O�!��V�]�����Ʋ7�I1��#!��P`a��+N
tVոC@U��O(�=ͧ�y2����%�T��v�`C�>�y�F7X�Y"E�K�$��!�n��yR�@�~.���WGK3;�X�+�l��y�jte�)PBfV(=b�8���y򩆻X�|5c���D��A�����y�/��.Y,YX��֍;��Qe��y�*V�w 4(y��I:,�`�����䓫hOq��i�ݰX��e��4M���J�"O*i��;��u8oH���T�"Od巤Q�@� vhbY1���y�*Y�� J�P�A�ZX��gX�yB����.P��$��9�d����y"�_T��qjB�9D�0�cT��1�y��Y�`
Z0�/�Xi�Ç���?a���S�q|��� q�ȴ�Ӫ �ގ&�Ԇ�+�ruӢ�_�"���D5
�C䉺)#ެ)���k��Y���fǔB�IV5P��A�Q���l�O��.�lB䉎u�2YH�H��QO��ye �r@B䉣xك�i�"������(qu(B䉃0�z�� �,n�	��\�p^�C�	*�#"'M#���\Y���$�O�����/^Ǽ����Ӹ	7� �L��'�a|R��	ejH !Ő�n�L	�Wl�=�y��S(��ժ�!�h�i����y
�lƎ<�bC��K�bQ�v��,�y�!A�CJ��%�X
lc�eI
�y���c�X���/B�܁�ؙ�yR�	(g�[g�.@��:�/\��y�-R.K�,h����<KF���y�*�Og�����-J�q�&l�y�D�(;��ȃ��Tp�!��H��y�˞%�bH(�`��`B�І��yRn�2Ud�s'�'�Xd���G�y�f��F=5�
߯/D��6Jլ�y§ 3	$v�!�G�)�,щᇇ�y�*�w:]0gG	� ��Õk���䓓0>1sJLL�v�[ �H�5Z�|JG�WC�<y��B�6PJcn�[���1�o�t�<��d�a@j]�C
H:usNHie��n�<���K{[ެАM��=x�t����g�<�@.�$�|kB�[P/�`ąN�<� n�Y��)#W��B0�Έ52��j�"O����FO��8b��D��h!U����	��:�BGm�@̘9��C��B�.-D��mL��0�b�'Z�bB䉪(pHt�C+��,��b�/q�B�I�JlhUXg#H4x�h��L�=!ĢB�	���%�C%]��e3�/	��B�IV�,H��aܖ8c$lK�ύ<BB�	zd0Д�Վwd��'�=��O ��č	^L9ka��=T�ft���	U�!���n�2,�@�ߵ;��H���u'!��ܡe���u(I� ��Qo!�3:4m"fm�̨�n�)�!�	-4��=a��s��ô$n!�� 	�<rB�@�:�\q�3+�!�D���ӀfT�j5�P�PI��[�!�dӪ ۴�"7�E�! �=�u��	�!��C�lq��A�
e*��� +�!��Ty-�A�M_f�b�c+�5"�!�䆞>h$��ʛ=��b���S�!�/ڎ�r)�&4{h�[���3��O���$
�Np0�a�@�"�E�D�!���J�P�K�zjT�JS<
!�$�Y�U� Ύ�+WĻɍ1H!�0��}`U�Y'tFRp'��-�!�$o�1�'�ەB�r��匮f
I��R�jT����3'�<t��S�eǮ4��0ղ��Ei�.P�d�0l�� t2I�ȓ�b-����	"��f*F�O.XՇȓ
n�}��C�n�D�QL�ȓ>��4�K�b'��3D$!5���V�.�� ^:O�x�Uc�:����8[n����0{DN���0mb�Ԇ�:��h� W�.�,+rH�ȓ�Rl�L�H^���E��������IC4!
�,q�Θ�	��ȓl�z`��%�S�m�Fn�#�nهȓ)����jtN|=�aUV�4u�ȓS��q��!��JP��@)ev��ȓ��h��K�����j˧=��цȓbr�e�f�C�g0 �F�P#]k�U��m)X���;QpR�xª�E�q�ȓD�M�V,�C���4m�'�bx�ȓ(�.��͐�Sd�u�I�F�*-�ȓR{�t�sa�V�����"�h��iԒ`[����h�!Jǁ�G�����G=B���,�y_������Qz����>i��LFS|���+��_��m��,��A���C�/�QG)��@����t�������`iH>'!�9��ʞ��툤�/D�H�6��*�<EH0�����UA'�-D�P1�HJ(Y$Q���D����CQD,D��B�� �`�X$��KD�w�iJ��*D�,J�#H.���J��Td�Q�s)D��"Ro��A�6kxȪ1R`&�O�����UѲ@�C�me�yhp/Z�Z�d4ړ��OD-jb��L�H��+�,%�*��"O `���&�N���B!Y�m	�"OД`�(�<z�zh�ǡ�zS�"O�1�$Ŋ&�1� V�8t"OʝJ��CJ��Ю&<�B�Z�"O�۰aw�ꔘ��	���-I"O@�
!n�4ͺ���ܘ�:M�#�'��'
ў�Oļ�)ŀ����M�S
�b��� �#sH�1�H]�w�#�9�B"OT0f��J����ܡe�""O���7	�� �  ��)��q"O��׃@55�QǮ��Y��Y8�"O|-C���";Ă�����R���'���ߡ��9����,J/N5���7]�|��)�d�T���8�	_�1�ޓ�y"㑼^.@pB��L���� #����'9ў�Oufm���\�͋��UU��
�'TJU0��ޒ{����.��U#X��
�'{:�� BC�!��KS
?v2�
�'ܤ����g��� 4X�/{�� 
�'k4\���1�x�dAǶ[���Í�'0ax���d2��x��I�Z�#H��yB,�P�P�ޜEX���a*Ѫ���hOq����w��i!p�YÖm[�"O��2Ĕ*���0q!���8
�"O|}���*{G��Q�{�xY�2"O@�	�@�<\`*0H��k���H�"O�	Ѓ*
���RAG�[��md�'�ў"~�1EƼ}��є$�#9�z�yG�	���=يy��.<C�D�k
�C���2tό2�y�X�*�ȥMT�)�6��>�y��Ģe�>Չ�& !��,x�����y��9L�J�� �Y1����y�(�����F�X=JB�A5�y��*[�!��y$�����?����S�v{ٻ�f�)Wa$�A@[�j@2�ȓH�������<��	��M�.�=��W�l��Bb�7�V��I�*x촄� �2\��枎8_b�����L����ȓ#��49���?�`��\Y�^ԇ�.1�0� �T+�2%�0`�T���	��)�a��͜P�A�X��8�?��.\�y��K�0�q�ë�o"  �ȓrR��c�� 9�HP%�`e���rz��1#DVzt�!ůs��Y�ȓ���jS`�i �`$)���F��+�\�#bK�(R@h��F)�X�ȓt�H��9&Ʃc4G��cptȆ�|y�Ԛ�L�8'h�SӅK%%`
y$���'��>��4:�N)Z�����c�O<��B�ɌY&ب���� �.��-F�B���x�r�`�+���:�lZ2hfB�	�,	�l;� _!=��`3e��U�C��:Ԯ���M�Pv�D�fA��ftC��<2�b=S�7����a �~\C��^a�����܂��[B�a{ C�I�od���"�!xt����H�HB䉵<��mIsg%+X�v�m(� D{J?���	��S�:\�U.MX,���H D��QFL�6Up�i7�xX�=�5�1D��ca�U6E!��aپ��A1D�@���y(���0%( ��q5�0D�P�Si�>Q2�j֋UlxQ��d�<�H>�
�'L��h��P�[Ȁ��Օkv�A��x�N�Q�o�Ojv!ڠ*�_N�?���~:d։%l�`��+T�"�ӥ��d�<�s$L�L�h�'�&aT� i�^�<)��M�#����gG�Ei`X�D�N�<)�nG'f�(� Cl��[%\r�'�@�<YR%���C��:���A5F�ПhE{��IY1K!��X��"em4����H��8B�I�N���AE��u�8��%�G}6^�HE{J?� ñk�<S6h`�GFd�1�"O�С�lL?U���b!�&W3�@�D"O6!�w�є^�4�Bd�W l�I�"O��5�K�%�T�$�ڷD��b�"O�����R�a���_2G�^5��$�OF����-�=*5��*J�`ҡi�=r�b0O�EY��х9��ě2ٜ9�`��"O��jj�	2f�;bwD�B�"O�,q��
?�8mP K/Xh��1"O`�Zf�D��ur��4FI0��C"OzH��'m�P���P�YLxh�"O�$볈J�~�v\7h�.,�͑f�|�Im~�e
�`��T�c �8�xU�p����xB��V�zh�B�SV��훳 N�7I!�d(J����!Z�c�t%.d����"O8��@S�p0�Q��H�Q���"O�x3qH�55=\�S�m�4�|]��"Ou�$ͯ��eyb�d�l�1"O&�4�		1�~}�NN��\6�'w�'!�)�L~'��0��ɥ�@�
&�	� F��y"�ߧIIZ���0f� aˆ�y�����Q�S)(萣�;�y�+ЍG�*-q�l�R�XM���M��yb��:T
5�$�C�0������y�)֔P���e'G�,�Ѷ�W�y�V;�h��7D+`�|����D,�O�Y��fQ5<ײ,s&%ОO�V$�0"O�0�_�g��\��M<h��`�"O.��D�,�l��"J@���$��|2��5h6az�CPԆ��Aa�]�9����y�E��`q`�Yi�)�D��Q$��y���9I^��r��3�Hz� X<�y�*�>-���E��9�>���Ɲ��y�E~}�Cě�3�.C F��yN��.^b��}D^Pq����y"�\&(mQ��1w<uI/��?����D�<a����5e�Ԩ��-�PSE��!�T({��b�̻~��ј�,��!򄛑F�9t-�##MT����!��K��er�(��a�б�rO[�e�!��-)XP�0��E)�ʍ�r.�<C!��
	Z=�� ޠA5��hӔ^���M��4���̰>A�����"�,�P/#D���G �Y�c������ #D�8��`�&>-����e̮>�p��$D�,a��(���y��ԣ$�D��&%D�@{�F@2Bh}	�n�3�M�QE=D�h��J�?p8������ "�%H'�?4� �2oI:o���h��'H~٪���H�'ya|��ߊ&wf��Ӂ�$q���Co��y�g��R��H� @��i���*��3�y���sfz� ���a����(C �y�%6g����Oٖ[ ԼRbJܦ�ybM���B�jG���V+�I�Q��yR�߮+�,�"L�G��:��Ż�yRkOi��0���̀Ft��i��+�y�̓�%+ڬ
����f�iY7H��yRnKd� �3F��¡�f.���y��h�.]��u3p=�jψ�y"��E�%s�L�n'�!+�
�yr	�8��܃!�	:��p&��y�j��-n�����V�8z�x�	�y�_L*��҈�5�@�Z���1��$%�O��d�-8�Ĭ8&�6"U��9�"O� dDzI|�|h��\	5���b�"O(QI��!&�e�FG�7f�<rb"O��C.�%3z� �GJ{�=�""O��+����_�ZV�]$U̸�p��S>���A�; 8�a�G9�d�G�5�O��uP8��`¯>�j@�SiH.W��D+�������9L��U��"�6�a�8D��r��0����w��U�t�"��4D��6��.��Y�c�B���$ D��:�ڲPM�؊`c	
,ތ�uh8D��aө�#9Y�4l��]��)�Aj�<���#}*�(�(\�w숵0w�^h�<��U��} �ϝ>2F���f�IX���OҐ�`�E�b<��'$'9fm����dЬ'?�u���H��>��'V�^>�IJ��\�'%W)x��&ޠV�@`�J2D� y@,ʄ(�PbdJ�ޤ}�A�+D�X{욇37�t���_H�\PGf>D�����W� ��ز���;cƸW�8D�L"S͆-[: "�J�Z����7B�OT�=E�dC��'�$�U)�kj(�Lg�!��"gҜH���̆&Wb�
H�*�!��:Zn�I��O$%�\���� �!�DV:wJn9ڰ0 ��$b@�~�!�D	�'Z��a�ă%Ŏر���pzўL���+q�6h	���A��+�H,ZO�B�	�\Ppəu��7p��e�:R����$�S�O��`��N�<JƸ�!E�M�7�C��Wl�x��l�@�j4	��{���ȓc��1��Ȁ�!�Zy��*�;>��ȓXġ#���l*%J��j�����^~�s�@��y��m��-N6L���ȓ`���cI8\0��p�Ҷ%L*��ȓ2��`͝ 0u��:F�I�&Z4E{2�'�$z$H�1J"@�jE7)t$�����y�C�gH��OE�|X
R����D3�Ov��
ܡq��K�/V�e86"Ot1���ЎW-0�0W�WI�lB�"O�хJ�/.��6G�&b6`���IE>)��3@T\RA�ֳs�l����3D�0K�%ʍW�8W�S�q{�$	�
�<���Ӣ�^�#����5���h.B��D0?���؏x��\�%�7d�v08�kRAy��'�����2dI�&�١+#:1 	�'����)���͠v�L�o��!��'3VhxC*�m+��;eoʋZ����
�'1r���n��eQe\�=%V��
�'j��Y�T�;�p�PR!��O�%����hO?�p�.��V�rVJ�
�}�a�Hx�<I�̌A���Ǌ ��`ht&i�<���.m&�a��+��/�%ȷ��d�<1�(�
5"2�P���QCRd�2�K�<��ήr~h�"�T�]���#KI�<95��b;��C"��Z���І��]�<��B5c�N�хi.�\�e�@y�)�'M989���K�p�j�R&EXC4�ɇȓhfh�gg����ӈ>����_x�<9��ͷ+�V8�CL`�~ YŎ�u�<Ѱ*o��Qr+'|�<�`��BX�<�%�()d�&.81Zd��H�J�<Y��5]�D1KF2v�()B�L�<�	�*�5�a�	��9d[J�<!���
�	+�.��L�0��HyB�'��c��x�0)�@=�(���� |a*BO݆�\��ր541�"O�8�gL�	�����.����"O�c�� -�V�QɄ�.����R�'T�	n�)�=qBΆ�?ST �񄁟��*�	�l�<�P�\��`�A�8��H3�g�<�Q-O�d�>����ـ 0h����b�	I��`P	�x|M�n��!�tp	$D���4E �b;�=愁�;&�K��"D�8+& %r(X�_�B��SaE6D��
��X�d��v+�gG��P�A�<��2��m�Ba?8jh@ C�KL�|ՇȓS�j��g퓃f'*��؏n��݅�i�`�6",(��˧hY��r)&�0�'��>��*V	�!��B^�^�е0�k �e*2B�I 6�Y�� �̮i�d����yBȌ�d�B�&�dT�@Y����y"��ow��mG�X$��;�G���>a�O� Di�=zԠ,c�ȅ�^:��[ "Opܰ7-�7�����b�h�%ZG�|r�'�az"� �Ӡ$���(4І`_+�䓑?��D1?A�f�D�16bPcy e�wM^�<���Z+�� ��?i���@�`�<�eo6u }B�"�����@�OV�<��/�vb��Yr"Q<b�HŰ" Sx���'�dK�P�8 ӆ��$ڨ]1���hO?�	�.���P�S�W�h4�}�bdU\�'�ax��ޜ\��x�M!-�t(��ǜ�䓉��3�SJP���Oʠ�JW G
1)�b�<!o��4{���M�M�^�q�[g�<�A䜬1�)�ɓGݠ%H2( J�<1�/F�
�p���ʔz�(У�͆D��x�<�S���@	��"]�uk�˟p��[�S�4�'��	A$��$�T�K����CY�1�LB�Ʌq�8�����~���e���L�B䉅%��@y�k G��Z��<\�C�ɪfÆ]QT�&<?��s/ӫahC�Q�v�;�e.V����!�mVC�I�qcl��@���C��1�N�'(cLC��7��`�H�8}�W�̲C�ɏq�xИ��ԁR� Ŋ�x���2�S�O<����ތf���ZW蚶gq�d"OV=�U�V ����Z�nWU��"OD��:��yq�KE�8�H��"OB�(�cB
FJH�3%��o��T�S�'��Ez�٢F��ly�:�jY	a�L<��'H~ɩ��I L�h��dĒ�^�-(�'����	��7=YYtcί |dK+O����S�L�@�����P��OC��P �h*D� -��OUd�YUN)3.�ܹEm#D��%�]�m p���*@�.m��.D�0+vN�)���ˇ�4h��P��84��	�>Xr�ҐG
�Z.�t�Y�<�"��:X16H�ON�_������K�u���O�\"ыD�YI���C��b]	�'��"�N�K�R|�Th���8X��d(ړ�y�NY'_�"]����q�h�8�h0�y"J�+e���:� J~dp���ֲ�yB"۶"��HA� �p� �"����>�)Ozd��G��e�-�ʖ��C�=D���!J]
tT�T`��att�" �ON��!�)�'	�R�`q���t�T
E���Ѐ�'k"Y��o�$���)�l����$%��.���k�X	J&"p[��Z�O|�<�炂�56�����ڜZK��Y�B
u�<� ���	�&l�2YB�U\�2�"O���cD�2)i6����&gJԨ"O6|�F�x���P�M-N�6C�"O2����
���⠁�bp�X�6"O�DȤg���Ȋ���;G`��7�|��)�ӄ'�PU�ˍmd��˷�H>�(B��,yθ�ɖ C�L���ʀG�/R�B��7�Z,�� ]!�켺�H0��C�I�	�Rp��NT�|�h	c�:]r�C�I%\��y�"~�8�@�dv��B�ɡ_ hA4��`�J��QHS��B�ɶIT��/�o�>5� B v�<B�	�Hd��l��mx8�IF@´B�,k4���� (=�T��,Q�0C�	�AB���T┦#$4,2�nY8#�0C�I�_�}��"Z$7"�ZtN�e�C�I.8;�k�)L�)�K �n��C�ɅLX���7�[�G�|y��ž|�!�䙴z���2o��߶��vD_�m!�M�;��(Q�/:���_ �!�Dֻ�R���
[ͼ%R����!��ȓY	20��@>0^"���,�#F�!�ײ�x�B�8cpvh�lTG�!�D � �"f�~*��j�!�d@�`��BT�З#FP�2)�(�!���MP�����LKx�`��!�!�NJ�0����$�n�i#���`!�X�<9�h$�˶��R�˚��!�ĕ��45RI�Gޢ`q�
�&�!�$�X�8ڒo`+��*
9B�!�H�o��
�eC3(��HY��!��������+^*�!2���-s!�Dډu�Q1���4%K�N��!��u丼�$�ؐo�h��C�xm!򤈪N�j쫇��2~>�j�@�8�!�ό~~%��ס-f�e�P%�=@�!�d�(S/���T�XIv։�q	p�!�PA���5�,V^�-�d(�.Z�!��G��P�t�L�JK�5H�5<�!���d�w�}W�TA�aX
u�!��,���
�#F/g@�Q:6�_G!�$W��"��A-��s���;G�!�*���(7熃,r�<QnR:�!�WY�����N�8h|\գ7�>YG!��	Ħ��@�[���+���Y!�$��!
`4RS!��[B�����X�!��u,��jǽM���"f팅#�!�d	^6�<�a�@�`�;s�(+�!��
+Μ�"�_-8V����	�(�!�$C7*XZ�e��-	p	�эݡk|!�$��@��j
�,;0-Jti!�M�x���փ$|���=|!�dB�4�t�@)�He��&Z�6�!��֭\hT�%���Y�-Q�nʩ5�!�$ϳ]
�Z�з�.���U�!�D�;ef�����$8d J05+!�D�+��}1� �'II��CB�o�!�D��<٪ �E� 2\H��n�iD!�d@3��I�^j�]"���Z@!�`3�H#0�؎�̢�FK
yhB�I�&e��
�.�H��K�ƅt�~B��C�f�G,q�à
DX[�B�,8{*P�R$��M0�e�r+xB�	�z�$�A�K�F�}��e['EVB�)� N���H�:��h������"O��)�-���6�Hg��	n��T�P"O�9A�HN
�u3��ݬD¤	b""OTA�@��-hb:���K�X����B"O��qG��:�R�h��b��	�R"O0�`C�؛*��1�8V�,�W"O<\� d����B$��zF��a�"O�]�f��S�l�9�A-Hu95"O��褢�.�(���F�Li�"OBura']4���=��M��"O�f,X�6�Blr��P�G�|-��"O lYW��4� ��|Ժ�ѧ"O4����o62�Sd���M t"O�5����5�@�)qi���~|�D"OL}A�n�EHƅ2E�F.*��u�"O8$�Ƥ�-���ɶg5C� ��"O$�82'�.L x@iB ��Q�"O���g���BUʂ(ƅ_����"O��RKe�`乲�Lgj��z�"ON�����2X��+�	E<Upp�"O�q��`��}�tW�qq�ѹ"O&I{����_��-��G͠jEb�	�"O����I!~�1w�V
�"P"O����,�5�Fn�]E"O��q��>i�*�X�o:]:n�K�"O���2�ڤ+�}y�i�*R�*�"O�� P��e�(�JG4�@=��"O�S��̰ Fh*R'^<E���E"O�}�ǯ�}�fb&a� ���2"O$�9�kR�0�Z��Q�_M�X�@U"O�4��/7GT=����`}(�c�"O�(��o�A��M%KӶ�y�"O��'�� ���Gɱ%s���"O½ࢊB�/�`F^�I�.�!�"O:���AڢP 9:�NC/6���@c"O�0�ͅ�-��(	�-�U%��1�"O���5.�H1�����QD"O ��EK?=�&Uj#�G|���Sa"O�� $8E̪����4�9�"O8�)u㊕y��ࣰ�I��.�D"O8]@�݌Oa�ͪ���A�>�K�"O*����L�?��1&K�q���`�"OR�@�Ӳ+�0)`s]�!�"O*؃֚S�U���?I�$�s%"O���7 D)9"�|زe��|�&ك"O��bC$T.XQ ��&d���}�6"O��b�e�2wn~lxg"5z�t�h�"OIs��A(%��Q5�N3o��c"OX�AS���r�lXC�NX&H6"OF0D��-�����O����T"O@���a�lo&(�����x��&"O6h�H;���tm�R����"O�Ɇ(ӳ>���DmUf�~���"O��FC݆L�ݘՉ�K:(��"O*�3��H�*j�Z�Iӿq�D��"O�4�5�ʖ\.*I)p�ٰ��L�"OL�їG�F;�Z���\8��"Oԁ����$�<��HF!t�1W"O�1�"R eR8���۠I4���"OB)��ʨ[�0��Nߞn���qP"Oα#��
|���3�-ܢa�XrP"O¼��kP,�-��ٖ!h�BR"Odts!�R���,Ʌ�� ��i""Ot���>j�^���U��)��"O� ��hǄG�`	⣣��Q\�{@"OT��K:����@�ĳ/C��"5"O:��i��"ul�ː��+p B�"O0���K���1Unȭ4i��"O�K&&��+���آ8 -��Xs"O(����A
9{Z�B�@�r yI�"Oh�[�Z[Bp!a(�?C-4!�"OzI�!��8��+3.˱:�H�S`"O"-	��.�* ��N�n�2�"O��E��?��T�SȀ�,�`"O��qCg�-���`�F�VL�"O0ui`�T��d�J���+�☰"O|�	E��"H�:P��'
?k��9��"O0��! �,bx���f�>�9�P"O��:sOQ���$V"s�D�"O�)*�$_�2 $yQC.����"O�	�v)؆r6��C�R�u�X��"O^��S�β%p�:Go
)$w�s!"OF����:@��1�R��]ї"O*7�8(l���En֋oΝ &�#D�4��gΨH��� �T%>< �Y��#D�8a&F�7d�D�4+��'���5�4D���#*�#qo���H�3@��x�3D�̹�)7<�`,�h64�|aiw�1D���I� %���ĤslAS��/D�\��(̄I��I#�n�wN����-D�4	���c'�#aFB�f�$���,D��Qr�M)�F�7f߸$;�X��+D��GJ�"%ZDx�E$��rA�Љ�e(D���SF�D".ɰ�D�l܊5��� D��O>,�ƝXC��:�x���*D��pCLS�hz%��I�mV<ͣE�<D������	��b�/�4}��<D��37ɂ�HT�� T:��%���8D����׍Y\�m��hΚ8��9P%h8D��s�(��A��p��Acg6D�d��
�����5&��5
:D���w�͙��I�a	��t�U�E�;D��@ԫ->���7'�qb�IZ�%'D��CǏھ!�(i��ɢ/�}:/&D�\��ꕝI_(�*�j��#@VB䉏D���rFK�$��90ϔ�+�B�	�J���� `�	'P�4j��H�C�I%K~��F��:d��G�Y3�B�	'X���m*A��j�|C�I�#q$UZb�W�}&�1	�&��<ZC�	�ob2Px�خv�5���E`�C�I�E.p�yV��&_h��Y��B��4C�I�@�j��\�FN���_�r3C�I�ަ��7�Zl�t�Ŝ1F��B�	�\X6|`��N$Z�dز ��K�B�.h�4:��Z�{�zl�E�[���B�V졻�O 4�HT�b��N��B䉔�@0����7M�:t�w�V�MڄB䉬��f!�Be�?y)L�Aq*O�͚O�!�qisD|���"O��Pa�Q�����U.ظj�A��"O� �� �/EҰ�%C߄J�!�!"OJ��(ٕSR�5ءaF��h�"OVY�b�ϡ}�n���@�$��(�"O�%�Ң��\��p�!7Q�<��r"Ot�h�ܥA�H���;q �8�D"Ohĩ$"�3��!�C����'�qO��/C&"�X�rI��1��A("O�  �(���m����2���`��'�L��'�b�٥(�A�����C5�=Y�'�9�5O.���H�9�|*��d'�S�Dʓ�]\&d����A��h���y�#S��9�TZp�� �T�/q�<���O�(�-Oe������n�H���I ����!�[3Q9�Ţ0�׌�b��Y�hc
�1�2�4��=[��2@�)+y����Ñ��'}}�'|��#H$T]��S����z���H�'�&-�\��؋&q�Ɓ��OTY��O(�	j�Ӻ;�O��36+�3I�h�b戅�3_l�[�'��U�s���hy�!x2œ!F������'�ґ|"P����ʑ!G0|�D
U�SaRh�cVh�<���E3'�$){��&~��x�b�Za�<� �&�,����׼cK\Ը��Z[�<��Ƃj7�T2���yl� �,�Y�<i�E¥BP��Q��8I����eY�<)"�ҰV�2u���\</�B���S�<aL�%����9i��;ui�P�<�f�dl�Q�v�̭8�:a�$!�$�	O�$aA���T����)��k�!�DK`I� o]�h�V�2!�!��˲=�R��Gtԅ�s�\�j/D8��hO?M��9N�$�H�BѧMڢ��U�#D�p	�Ƕj�� �φk��$�!b7D�D
�gH-�y$���G2����*D��e$Եv0V���@C�sh�ʷI)D��Ĥ[�3��(�fj�L�d$�s%%D�p�  ��sž���6M�b�r��5D�H�s�*�`*��b  �))4D��ҐD؟+|���ߞ=�
 Ò�p�E{�����pB� E�:�Ą%-!�D}���c�ϥ9��y��IݪW!��(h��d�3�&��&��N!�d�6jB>�$�&j���0���n�!���g
�51���,�rf��X�!� ���ۦ�L(x(ٛ �ΏC�!�Ԕ|�i�筇h�����,^�	s��0<�I_ʺ1Pd%	�@
��$k�<�% �/\ph�3G�H�U�0R�e
릑���/�T�d�J��N�Ť=cBiF#C�ZP��6�q��VP��G&էg�D�'��~�#w��IF��^~�p��Y��d5�S�O,�A�BG n�&��B�L�a��Ep�'��+�ߓ<6�|	����T5����>Y��	��t|p��PdY>Ti�V*�	F�!�&�>,��gڟ�Kѣ:��p�ݴ���1���O�@A#��a� !��Ȋ2�nM�'F$ы���1�����gH-0A�xS�'�д��	
��uA�`ԛ'�LJN>����~��tR	�0,U(H����ȕ�y;<\�� �K�j����RKD��R��<a�O�ܣϓp��@gٖ���9��$Yݴ��=t��ifjݝ_"�-H�	�yr�Gx"�'���X���1���ׂ!H��4���d>��UeC-Iش8O^3	�(�0Pa6}b�'SP�zg��G���ж�M�C�f�9��?	��:1�ѡp��5ͺ�Q�g��k�!�_�z���j�$�@`�4p6�N�+�ٟ�'��;�Oq�
$z�H�]��dCr$P�M��=A�"O����♎>��<k&�0,��,;"��3LO��x�
�+I}H�Sdl�(%l�q��"OL�l@�Q�dЧ�U�`ܩ�g]���I�G��ʁ���fL(�Jː*��C�)� vh���ùl�����Yk��	tX��Y��[7D(�(&m-YV8��.��1�O�� -a��� qo�; V)0! $�\�f�E�^��p��Q�H�Kc&�z��D�?�e$څ|^x�K#��2�4ъ��L�<�#�U;]l��@E�,Z�D4Z��dΓ�M�O>E���d���B��H�&�2���J��'�H��?�͟��J8jYP�dj2
M��֞~���'��&�'���3k�u�q
�͉���a��>�e*�>�N|n�?'v�,Sp�)!�U�ƍ��l����ēMj�H���؀"N@@(�nLE���Ml��u�=q��T?��r��.�
|�&g�g7�A�:�c6�I��P�p�圜`��xT����84�x��)�S�9�ؙb���-�`���	��b@>O���۴�ا�O���t��0e�`�+�23+�y�O����5**PK����Z8�D~�Gx2-�'�?��w���d�ЀII�58�Bʇ:��ȓ�6�8����+�@D���T�����p��>	��3�f�r��AM�Q9D$����
���ȓj�Z�q3�
�;fE�p��_	�@��O���G�*�(Hb�/Z��O��@u�u!(�21��/����Pe3D�L�� ʗs��yu	��P"��#0D����P��8p`j��a��� /D�dY���Zc��` �]&t���XAM+��6�SܧVJq13��};�B��5A\Xԇ�A�&	��d
��J�ふ�(�Gzr��d�O-��i"���x��2�@83�4��'2F1÷Q�h�x��B�G��4ճ
�':*��'��,}z�;�A]�t�މ�	�'��U�T-S�$�z��T�6Mq��'�p��K;3�Vp�қ@�^5��'����%�ʢb*�<�D�)@�f�8�'ˮ��D��i�z923 �iD�Q�O���$߉j�X���l��&�.�Ԡ,�y$��asCnJ57��Yc!��~R�)�'n:T�b�J"�� S�ɫb�BL��ID�k����D�Eh	�eXe�$(\(�ȓF���c�<A7X��`�Y�"�����hO���`I�/ԨxS��������T��DR���'�(��`�پJ��5#�;6 8��'� �C�Tٜ}:E�92.`x�'�*��1ڬW߆0����[�s�'��,	�)��p�왻������0>�N>!WG!�H�3��	W�F�zg��<�'�Ă�-��؆C�8��S�Oq}g?��(�9$P�-4��R�S/0�����"OP����L�o�D�������'��<�	�O�8{��H�cG���Fįw���/LO"�`�ׄJ�[����&�@px�� ��>1��-�b��$'��3��C�&T�J����8b�H���$(=��ښm�TXb"O���QMX)?�`�6nC�U�ݐ���d�ڃ��D�$@q�%Ŏ8`�Ҍ�S�<�6`�F�8A�_�$H�-�t��<Q���6{�Ѣ��
2R~xx6NO'��c��D{����P"a<8���?�$������y¯�+a�� V���r�|�"&���y��/qGF��'X:w���!gk�%�y҂�q~���T�E^F8;�N[�yr  ���3�IF�T��X٦ ���y�!H��#*�Gk�A��V�yr+45P��"@L�.D201)5g��y�̖�r��a����>%"T(J�7�y
� ���#�uZT�ħߡQ�����"Ox]9�D��b�C�ĝ-F���""O�Ȉ�,���1���N4Xa6"O���dl?��(d�9�1H!"Ot�S�Q�:��eH1�P�U���"O��y!(A�4����0�-\�r��"O�����k��P��B��zG"O^�S KF�Uw��KDIQ�?� Y"O���G0�[Ղ^��ڰp1"O:��ЯJ�j�`�Ȅ� :��՛�"O2e*@�B�\ܰK<�fl�S"O�]��!W�/�0��-ʭ0��<�"OACU�^m�Hs$���1���"O���U
Ĳ+H$A!�ю� "O�e�"���DIpӬ��VÎ��u"O�]��'�:F�nX)�+P�nI�"O$r���j��݊�)|����"O����:��H�$�)cy� '"O�b��E/4%̽�6I5p
�"O���Dbϧtd\*���5@���"OB�K���?A4ؐtȮh*�At"O�$��˩Gz&�j���v� "O.%ఊ��l�\���j!�i'"O
�§�˘24v,�hF�r�us�"OD`�
�z�`�f�C�~�xV"O���'f�.�0hӲ�&O����"O��6���e� R�-=��B0�J�<��
H:`�h�@�pN���G�MC�<��@N�?C�$�I� 3Zt�v�XZ�<�#D�>?~��*�o�1��bX̓`��s��;M
���=w�t�<)U�S "B���^�xTx�Z
Q�<����G���-�#
U���T��O�<Qテ&ݺ�`��5����f�@�<a����Ҍ��Ѵvʍ���@�<� ��&�{Ӈ� <�āp�<���Y�B5���׳*V�e�3-�v�<�v���p攕P�Ƃ�wvL�ѩ�K�<13 �/m"&P��NZn�! fN�<id���Ԥ�>p6�Q�VR�<A��9 �:��\�2�����K�R�<�t�Z� �����y�6u�4�QM�<�C��T��K��K���{S%�f�<�d��P�R���Ki081[P�Vg�<��E(\��}�D��tJ<3���D�<����$$ �X�B��r �A�<��N$(��SpC�P�� �`�Yj�<�
ߣ(Y�@��@�
�y�g@e�<A���VTllá���r�J�a�+�a�<�剓>;W����Ȟq�l@��"D��3����$�3��pVp���!'D��3`ڕN��r��Ȉ	�Ppq �%D��W"Ҭ	�n<����TB�r��%D�Hy�o��#ΚQbpmF��v��M/D��"�%K!Q�TZCÙl�^ҁ�0D���Ug�m��� A+{B"�.D���Ɠ	2m���9o~	�I/D��F�V�H	���� 	Ap;F�-D�$��+D�g1|�q����&�[��*D��������Ul�#m7ܬ!��*D�[TQ/X����.߳2��J��(D����혋u�8ys4�V��`�A2D�0$b��+]�a��h�H��ԛC�0D����(=7�yc���7IJL��0D��`��w#�1�u��.P��D�,D�� ����C�%8tY����L^�iv"O��C��Q���� ��_�`�( "O�)٤�&S:�q�`�4	���"OR䠳�!�Ψ*D�*���H°iv0#�'��	rC_�cd�rǋ�\�Lu�(���2a7?�s,[�xAXݑ�GК~Dp�+��Vz�<�!!Ö9:�<��	v �+��X�
��9�c,��A&�M5.��TrA�;u�=�"O�TQ��]H3��b�!�I�"81�䈗V�qO��#��Y���DNݫ}��"�$�)ۨah�M2D��ۆ�M8l�fbt�+l^�X�>lȨ��6�O���*� __�D3SiR�m���'��H�da�A~��G�<z�Z��O�tP�'�Q���x��-��!��l��	��a+�+f��Z�x�FV�cU�O�On��b,I.A0v�v�T�# �9#
˓]�n�S�.���|"�  !(�b�P��R��'!�$]-���@n��1�a�F��%���VhZ�[6qO�����"GƷp�`<J��m�PE�V"O�(�b��Ey��FI;d�%"�,�	��-)��L<�Q�H5>��k֮�$�f4(7��vH<9"-?ԨhI��M,Uba��E�9ɖ܃0�*�O>��d�_U�`	���R$���Q�'�D�*�K�M�I �j��aD<1U!�$�!XhDC�	�2�\u`a̞��l��
�&��O�`��J?�)�(R\�6��[�M����P+B�	6Zժ�L��A򋝷V�B�I�^�F�ߺh���5↔r��C�I����b�S��";}�C�7s!L咒(d���N�(�C�IKe0�KV��0c8t8׃�G��C�	8��{@A�� ��@���C�5kh�Iq�
6�8Y�	,A�JC�bX�{'D��q��ATIG�#-.C��ol:8P&l�j����BB�I�n����ٱ��	��ЂS.bB�7�P\[�J�1y��ce �׊C�	�H�]0�Q�9!H1�Ԃ�Yo`C�	�.�o�;FR\mKB��e)RC�	<�h�aԈ̕e�\�8dmA�(C�	�7�\̺r��t>���� ��B�I�9a���ҥѤ|�{b�"'�B�IC�b1�FG�-OX�������4�⣓�5��?M{a�`y�,�7��5�|]��"D�Db�(����Fه"x��`_��ؠ0�|rO?�g}2g+4J�D��?K񌽠'�,�y�]�)��񨧭YA��L�fD�ڽ���yܐm ��N��0=ɳM.^��e�Ee�"~}�|�0�Fpy�-��T�����|ZwV^5�wO�`��ͮ5�4�i���+ ����'�҃0�P�'��t(�"E�k��+�/��h�!���01V ��%����X��T�8'�b�qq�]�<&�=A<��v��S�	��/F�9/a|Х|3�Q!'^�_Z�)�E�]{
	ӧ�Z�t��Ј �T&UP��2~_��a��JXT��e�~�B�x"E9z�r�3gۿeI2�6��э,��ں��<I3ޱ�'�^�&��i���	�@�	?q�&iʠ$S�R2TԠ`-F�s7�$@*�K����<)��3c�D�%/ "D2���	�0��%&n�5[�*1B�d�Z����3a�l��/�!&N&�ɵi5��%s�?����u�ˢS8V�(�*��u|R��Y��(2�7u
��T,��t�D�Zӫ�u�RLXs� /L��1��E�6���׈�4r��,͐r�L�3ًs�@\`s� /q���2��G���4bU��#x����D�~��@N�|�BE����JJ,���jg��qPR���v�m��D�;��0��"H\r'Ϛ&KL.����	�g����ٓ�I�a�ҹ�N�*V���8$FX%�c��9&�:n��zg9�L����?E�D�Q�e{HQ���_�,�#�$\2�y#6g��:ޕ�%o�?F�|�UcX�cw\M��A^� �sԛxr�'��lذ%�"k�n��&�J�Z J@2 �]�1���:k�<��'��L�e� h�j��<+�n�1��Af ��VH��Ni�b�	Yol�(4��o���)�$ΐ��,3L�"ׁg��,�PC[�_���2��)ql0&H	�7�����*,1B�B�A�g��,l6� |��FQ
>ԙ�'�Qf�P�=]�6y��]x��@R�^�^�:m����؀ �	Sd>�6	�B%B�h�|t�B ��1D���h2-^0doZ�[蓦ɾ5z}
&�
�o�\��0� �?qX#V;M
R�4.
	p1�� ��!�r��fl�Ojf�j�'��nEr���n_>GAP�I���)ts���D�y�ըH+0/2�
�n� ���.?DF^��'1.h
�m	2*�W,�/.�LM���Q��0�B����铄5$|"�k�W.*Xh�#�!_d�5	W��	���Ae�1*)���]�s ���o���k� �6��j���%���'�Zh���]��)�'�)�^�n�;,�=nG��AS�V3{]���G�-��	�d��k�(a��pE����i�&}��含mV��OI/|�d�4F2a�� B�0}r	��f�Ʊ[�D�}����o��1�8�P��vܬE0wBΩ��yK1�	�5(4�����rڤM�~J�G[�X�`0
��S�G;�Z4�̌@p���%� G�.�P�C� D����Ox����<���&��ƍ�9�z	�Ѩ��[�������+ݹB�:&`[*t嘨��g�-U�ԍC� ��f	��"���-��J��'�X��w�@-V}�%��5ΆP�'`%(p
ʌ/%��Y�>Ap�T�XZD1LI�P�H���L��\1��y�G���(��2k�I�b���5���E�S��~	���Qي��c��1���A��ӱ��bL-a�¥f9f�R�9~��>`�gّtVdk7H?7*�x*��/ʓS��80g'X�|Zt{���o	n�r�@#@�}��,��G�"��L��.�
0
t�WoO�z�D�𙟜��F_�xE3Ŝ�ed��"�)h�=Y�n��PWƑP.O?��Ӓ=�1{�!K�?Ḅ�gMZ:)a�#_��8�s��}�d�5��U0@��a�C��6 ��)�J�>���X�\� �l!�	�]�(���9T��z��0az�pV�H5X�|�`g�-��(3�'W�Y�b��3b���a϶~/5�U�Z$6�����V�zt`����8�� ��׭dl�ȰgG�|��&��p�N��T���x�@A$Vu�<YW�-F��IP�I���@
u�j��R0e�,AQ)xO�pl�����y���Z�:��+�(�DA�����y".�Sa,���
�UG�������j䜰	e&+R��`h���a�Ƀ��T��E��f.����&�?h�bxc�6A��~�2K��pA���q�"R��X6�,�B+�u�<r�UZ
a{�<20&Yڔ-�+h���ܩ��O♡ai��n�B@����x�ZIZa��������
�$�g:H)�"O�=��(�"��s��nz� Z�<��bL�2�Y��`�mCr1����G=ꌺ`�B$*L,���C7JrB��*@*z�(�a&��UJ��@=0�b ��A�.O����Y��xgOٽ:�,؛a��� �:�Z��%D���$M
��s��?��0� a�qՔm�@�=����,`�vKƶjWh!��Ľq:���C�4���@lڗH̙���ne�<uK&eJjB��/$�2��& \�̌L��M��-Lc�h��K�G����@���4x���_5���A!�z��C�I%^ <d�͌7
�Ip g�%+�R]�%��&k�ΒOP�}�j<�c�lΩ�8`A�DN:oq@����Li�f�U.,*�q��;G�*�ȓ"�(@�@)-�̵H�FF2|jnu�ȓ � qU�
M��w�W� ����ȓ���Z`�zAZ,���1>�\��O�T qO,�}��l���*cx^��]�TI>�ȓx�%9��8�J�#�O�<+��n�%�
`�B�i8�P��D�a���-��A	��25b6\O�ac���}�F���'��b���1$�������Y8���'A��9��_�x�噲��َ�!�{"LɀhM�8J�MA�O� �`��;Uz�2 *�� �'�����Jҷ)]�F�ζ!����e8�*i�J�����<P��̆KT%^,B� ���i�<��NI�kw,�8򌒠c?~�  j�X�'S�&�"��(��(�&�ްDA0� `V���A�RM�Z �E��y���in�9`�W?R~��0��N��yU�?�.J��L-��K����'����Ņ<�b�E���!���(�/�F�Z-�pjS6�y2� K�n}�a�Ō0Qh�{Gǉ�rL��OV7���b�Q>�|�����b����;Q��хȓ~�����kd�P��1'�Z�mZ�bҚ�K�!�L8��b%�\�i� i�BJߎ�S ,|O"�ԭ������=ZsV��`�ζJ�	��}k!�d�5^1��Ǉ�q�M� *K"o!�� �8"��U+�RQ��r�n�3"O��� �5�TXJ%�M.0�8bC"O&�A3e�S^J	*�͕�-���S"O��FG�|�3%0�*�ѥ"O6� �j�!�`�wn��@�@"O0�z�o�;�] ��� i����"OJ�X�lO�/J8T��� ��L�T"O�dK`(^K�t}��Ͼ4��,��"O�Q��S�Fs��9��5�V�а"OT	�����ĈF��0�d�"O:U��_Nj-���y�4���"O&���N�M��V䍐C��-j�"O��JW�Gk2�9FYAR6��S"O*D��5p��	�@Kj(��"O��z�ƀ>"B�����"*TC1"O*x�
*D4�i��3"�|<��"O�a7���x�ɑ*Dd�:�*!"O�-(�k�&(���Y��w��l��"O�l�f��&(C℀7G�&�\)� "O|\h�#�b��� ,�|+&"O ��2,�7!S���
��8|�1"O���`�1-^޸J��d����"O��� ߁N��E���>��Ԓ�"Ob��c��CN^YH坫Y@�i�"O��@"�c��l�Cˏ�G��\��"O�Lv*K<){��Y���8�����"OL]�]�n5
��掹1����"O�ܢ�4�b�H���!G�����"O��H����>�NE���7BK�؀�"Oh�Q�.���d�aOF)S�m(�"O^)bU�N WVX�2��	onµ{�"O$9�7�O�J�}f�8]f	i�"O�ap�cL�5��H7gԓH�B�H�"O�%#�H�>L��Q�2)P��|�{"O*�9�+�~�ڐ+R�Nº��R"O�pF)f�ȸ�/�@�|��"O��3�R1+#1S�v�K�"O�U1pBD�FW�d���N�bx�|s�"OK���=�ѠD�ie���"O��h��O���H�U@^@����"O�dH�`ћr��lbA�N=v�\�Q�"O:�r.W�����H�;�J��"O�D���i�@�cMW�>���Q#"Oƨh� ��~:­��L�>�4��"O�Vdݫ)%��j�?V|�S�"OR�q���G��H��
zf"Ovq3"��	�,�+bi��ڂ"O������7>|�*&���`�"O�9�5�`a�	9\�:��iW� !�ě�B�f��eG��.���v���#-!���)��@�C$Y�ڕ���7!��H�����>d"YC�o͚C1!�$��6]H���JW#F���ڝc\!�@�GU>x�qo��k]>p(��!�ą+,|<�b��:Ui��+�N5)�!�䄔��ɡ`�V=,��-ΚE�!���4w�xCV���b�LqslƎ&�!���}5�����t����Gh�!�$ܷ\�Б�tȄHF�D����`!���Mt k�A�H7���u�!�D�n��ʓ)�<@֕c�c�: �!�� �2	��)F�i�*��0���!򤍴�Yy�N^�^�H�[��Ȩy�!�$V3*0��b��D&�E2�(�6nS!�� ��!��-�.� ��ڂ\K�"O�(��	�V��2	��d�s"On�� ��|����3��6~����"O\d��i�N�hr�$d����"OԹ�>�� s�D�0S��"Ov,(ԧS+eu��j"�W	�0���"O��#S��Y��$�#A+5��#�"O��	Fa��X�ZY�'"O���r�"O�x@�Ì�;�T8��8Eyv)�a"OT���Ɔ:-)�n��;f�4�"O��ycj�9	���.�����"O4�+�C�y%چF�X�.�:F"O�p�r��|碥��o�7�$���"O�H0P�Z<�#X�4��䁡"O�Ly�Díw�n�����6��M�"O ���Y�S:�l�˾���"On�1���� QJČ)(�^�p!"O�H(��2" tԘԬ��+��\�"O6<Q��¸�u�2��%�>�"O}[�a@2z��P��	�/K�*��"O�m����g�X�4�
"{��IZ�"O胣�ѦO��5`�ۖ>�<Y�"OX��pR�e����	��LUc"O�9�#�X�%j��G�3�N��r"O
q	E�G�A���# P & �"O����➖@B�q	���
	���"Ov�3��F9�~,�A&�
�i��"O�`:�[�,c��S�/L�u�T��"O�L)�E����Ϙ��{4"O��G.�)^����qM�:\��"O�5�vFF��0��NR$��"O�IPӌلPUً�ʄ"!���"OJ��6%��M�|��B�_���Z3"OT8��Mdܰ��s�ǲ-s2�R�"O��˛/@��ї�_�
KDd
�"O(|4��0�G�U4;�X�g�<1g�"S�H2˂7�l�pl\�<��ŝE��3��KM�T�
���f�<1���dk��g>1kr\�u�FH�<��
De�t��";�b����p�<ADf�5QVLK��`� ��͟r�<1����z	jE�PH�$��Ēw�<Ib�Q���X�&%��+�F�h�e�<��G3q�h�pD:$�^L��-x�<�7��!_�$�U+I*[����⇂u�<��l�ր���ռl�d�f��l�L�h�ō9�'| ���<�TiAN�',!^��Z�a�U�%��1�	\f�v}Ұ+�^�OtuF��O�q��o4;pp)`����jr"O��z��Q/*��ڴ�K�%�V�&�ɨ&���Т��L���K�'�0���>Ro���V�D̴.OJ��f�9N`�O�ۙk���L�c�:	��\*2����FH��X��QЫ��dP��d
��Hg�ղy�c�\;y�$�"%�}�Ƈ�:r��e�"��&�+r�Z�my��Cg�x�}X�-9x��e�C"��`Ä-9�O9x�G�&m�20�f��p@B��*X� r@$�Āԗt� QI�$�O���JB�DI	BiaWJsEF�O!�O�𱳩� |���ǇZ?Z�Z��R���#�SD�$I�O���hM8��P@��9zNu�5f� {MA��h�7(���'��&Xo�=�$�DX�4�F�^3:���C��Rj��
n��)��-�g1�hI�AƐyШ��^29��IV���W~8���k���¥�X�D�<!�BB�j�j!I/]k���ȗ��IqƇ�2�@��v+G��t)�N�btVCp��)k�`h�����Yq�1 �T���F�
�k��Ұ u�˹k�HR�.ٕz�����'H�9�r��7�V��j�&(�ja�!R�Rd��#b:vH���t6=��Tf�23���Ľ?��R�Y~�U�UP�}P����,*s@^���'�� ��FB�R�Za�Wq8R���O��:v��($�]�U��?64ɱ��јoӠ���Q]Ǭ�S3�-3����� ��9�NU%:�"�3����$,~%��*L��L}�S��0*�z���9�����$>�6�s�BA���N*6{P�+"+�'�VD�`��(�I��酊'�(q���zǼ��ثD��ث��E�6���w��?h���
�H=;�^tP�I�zŲ��FX�D�����)4���R���c�Z]t��;0�o	�x�퉹x����lC��9jDHEdH1py�m����9-i��s�F�WL�<S�޶t�Â6O��x�*��X,P��WM8�۰-�{Հ4�?	P/Z$ ,�P��i���̘c�	��E�
�f�L�1r�"���~B @7Xa| ��k�U�hᠯ�V� �3!�2A���������0p%J �9��S�O=�x��	�uZ�BS&ػc�Ų��ƃ~tlPJǰij�cW�\�ZU���� 	��h`@�$�d�����d,�	6f4Yu�F}�	28�!�i5�|X�'���X���6>6�p��"d�r�	��p>ch]�'�0�I�m�iR�h2�S�?:,t��Y"Ym�Q��}���n�U�M	���[$e��1xx�H�뇻{��k��I�D�9�%�5~p��~Z�)@�Q0��-.s7����gګ�1�E҉}ڼ�槈��䓄9�ƕ9`��v������7p>A��,]�:01J�y���'��fL�A��@�D��gΜM��'�کC4O�&B�Uc�L2�Keg��JC";��˗�Vp�:2|z�!�W�0P�}�@) ��"��y�f	Y�hL=e��[sM,`��I6|O5����.�|!a'm�A���c��> ��lXՠR�&�R�\���M����GB#��O�2�a�&7z��p�D�X��q��$�$�&�1bf5y��b?�0�ժe�9�Ӫj�:�e��z�L �0 �lj�G}���iY���� �),�p�*��y�f��
)\	���2A��M� �S��?q���֩���"�N}�aO�Z�$��F<J��v��0<9���&��&GڄLtL�*�DR}�GƱ;�,p�#�i�'M�=iaA��7��Q�Ϸ!,ԃun�*���(c@�y�����/�3����gEi=I)v�д{��0�3+
l�'}\����g�E��H�<����'%#� �H[%r�0�C�^��P������mڇm��I��@�1��t�o�0D���������
]��F�d@D� ݶi�6�A�-�H]+�Mг�y�L�a��� /�h]��)��w�
���'<�����W�]�N�PO?��>�F獏'�4Ec��;+{��2 %�]��LY#��49 I�#I����{@,�*���Z �Ѕ8��(��ڽ�*ń�	2�6�i��:0��"�b{d"?��i�"Y.ؑ�_<< �S#�ٺ#u
��?�v�]��\����P�<�b��N�*ĺ�k���BiOy���6R��#�#
&R0���|�OӴ+g��0Y-�ɲr!+@�xc�<�S�^)Q(�k� �>�2��ݨ=Y���<db�u�Q>�X�.� 	o�.�@�EQ4�p�ȓVݔ%��e�=4��@��#Ŷ�0h��ٳhW��#ꋅi<a{��;CL\Ѵ�W9<��a"֤�9�p=�u��9t��)�.п�MCu
�����(^�l�lK��p�<��
*^0i�C�74*\Kb�Pl�WŚLD+S*�z�}�����r�L��W�e���"Rf�<�c��q�r��3Kψ0�F�`� A ?4�x	goN�	`��~�ւ2�-Z���
+�F�7�y"5{ �u!Ӹe߼���O=�y��Ԟ=�T�pf@�f���)� �0�y�	Ԕl�`8p�;_Q�墁��y)S�,��іo?R��`���;~�6���?�I��~"o��|nmK�愂���BW�y"��H4�t/�7@�9�ɉ��M[#�Ad��Y�)m����F�%8�!��q��=��	Oy������!~��ی����S�	Y �{G��O�!�-z-� �m4<,V�N�9�qO�gQCld�{����QN�����
mk��V�&!�d���`*$a�f�(�[0�:zS2��Qa�'@�u�|�'7�rt��-�\�K�Ϙ��C
�'N�LY����{t<��=n(�(��VQ�5��ǁ2�0>Q����,��A�%G_	e���W��Q����'����I�S4ON|���@�\hqa�/ѯl�J��"O*|g�>�"���A�6s�d�w�$�8F�l���!�9����:�	��,x�®^φA�G#!D��+EL@���P�:0~��#��8Q�
L�J>}b�x����Y�)����a�ԝR>�y&�ÓV�!�� �Y"�F)a�t(�w�;i��iE&� u�$��|"��"u���F'�H��A˒��=�d*Xu�.��t��g 
��9��!�4I����ȓ�(}���s"r۳KN/T����8b`��o5hY*����]9�݇ȓv
U� ˠ/'�����s\���Ny�غ�Gܪz���;e�<RU^��t�BDQ���""~��`C�' cN���x3�\IB�
�u�n|���c�|���9�j� �❍v)\��H���ȓ,��]�p��7�l�� �F	�ȓ|��h�ML:=D��Å�j� �� ���r��z�J�@P�
W����D���� �	q"���վY�bD��S{Jx��,�Q�h�G���ȓ5P���j�*mzI�	�"mqn�ȓ2�1q��߶?�P\S��"z�dI�ȓL���Q�R�waɲ��X�EGh��ȓ�4���ѓz :�b�bT�^��_�t4�b%ATb�E���,4*�X���F���R �x��ce�,���Y�'���xT�ΚS��5�A�(�
�'��J�V3_G
��
ݦ2�� 	�'���蔣�jd��� -��+�'����qf��T�B" �/ ��	�'��X�B�3}g�9*������
�'�d}����i�<�Ï�;e`�Q
�'zq�r�Yj��8aF��zʌ	�'��Q�A �E>fa��EN�D��'�����L�\����ň>��9��'�<�y7Jʹ
ă�҆ �a	�']�`�פܛo.��УK*��3	�'|p��9�n �S,��w<�0�'�A���&[��3dS�����'o�AhG����\jqkW�p_d���'�8�)�扎p���PNޫsh49"�'�p���le�� �a�l�@Z�'?���+c`8ya!�0}�lLَy��O�z�rp��ϋ�<�A�fR���'Z��Q�|,�i !�7r��Y�'��ᢢJ.j�<��R	p����'zh��e�G��\=*R�����'�D���#p�+��J�4ƐH�'�dEz���Ta�Tb���g	F��'*�s҉[�a����v��'t�*);�'��Z׬��m�b���ɲ_�$<i�'�����;u@��"1e�Q�4���'H��BP�{�$+��V
Ji�MH�'�D	 'P� ��!�劆��x��'��"=E�@C�4f�0��>�
t!���gg6�Bs�Ocy¥�6#�����-KE|�ʣ�އ13L�X���{�xݺDT���q
�
�����O�8�ZF�?Q2��K〉\�����'I���1��M.���]U>�YR��	3�ݹ&�K�%ņ90���%��� ÝkC�|��)�q��b:`�8�d�m�����^�~m�%(�#�CJ��h�����������,k��Y!֬ɉ,
�T`��>�R�X�=�����/,r�9���4NҪa��'��	�h��Q�6,�)���5����g�I!B���t�:qp��+~W�*��<�)�'h��mA�6v�6Q�$mR�z�J��ȓW��@��3"�d\��������ȓ��0lɂp�V���ٍ �5�ȓN>�ٛ�
R�
,+�hJ�(5GzR�'�tӥ��?� �E	[�yg��'v ��`J�	�.����Hz��xp�'� 4a�f�4��`(�A�'r�ٹ�'�lKd���#6����HПǪ�	��� r��l�`"�Ѓ�{$�h�"Op<���=J6�0��"k
��R�"OL�4�Ű �l��'�#h
�uRP"O��b�ր �hb��خf����"O��btJŊFX$��C��f���H�"OVec� ߒP��P[��)E��D4"O���D	JMA��K�
�R��8"O�	���GT4:u��F}ϊ���"O8��@#�&�VI����&dv"O��
��'�貴�D�+�P���"Oh\9�jCb��5��G#<::���"OZ �c�]�0Q��fi� " -	u"O�	A'f�$-{E�ԑX�A"O$� Fē:�A��Q�`��Չ"OL�c�A�T̀� ��.;��۔"O�u���� ��4�0C{X}��"OS�&*^�P��"Ɓ.Xx�"O浑B`�2_�,�+���Ie4���"O�R��k%�ͱ��P';O�p��"O |�jIx���A>=��W"O:��t��8YÜ<i�l�+U>P���"Ox`�ע��ę�+P�x89�"OV
Q#�x�������"O �D��i���ҷ+�1`~���"OlmS��1}�� ��.p�dV"Ox�����"$����(��6i�d�#"O���&��;@�ذ��GIPf ���"O����@�6I���#���dW�@["O�@�Fd��K^�!��D�3cT||zG"O�x�u ��pz�!�<���R"Oƕ҇bU�~s��"� �O�N�y�"O"������i�/�d�	p"O�h��B|�H��%�HQJ�A"O@u˶j�>�N���7�b8a�"O.�B�&�yV�b#Êh5���"Ox͒���z���*tC�-���S"O `{!���^dꑄ�=>��"O�����#���$cEp.Ƭ�7"OM�È�2p��ⓣ�r�
"O��3��ri�+w�M��D1	�"O�e���P\�V���O�C�蜒b"O=���ڑ�����@]�� �"OF�b�4��������HՑ2"O�!P&"t�$spE>P�|4s�"O�x��iI7[]r�٣������U�!D�t� &?K�{`b\�R$��u�2D���0g�\����Y�k%���2"2D�����4�(d��'V
o�Ыa..D���f��3�-i��8������)D����C�)��mYↅ�.1bQ 'D���&��^ncf��:~if�0��0D�PQj��=�Ed_#f�D�I �.D�\�@E��WGd�w ��oO���+D��R�/N;/[>I��YQ0+D���a���7�ѝ��rPL�Z�<9І�j�����/ra���}�<�ckS=�K���d���fN���C�ə D��:��;MaPE�aI�8��C�	�^s�Sm�(J:Ł�-E�M�C�ɬ&�� ��U3E�R@#�	�D$�C���֐�pmW 2Ft3%��$��B�	%Nm�šd������F�T!�B䉃}��@��Ή|��cP��]L"C�I=3jd�򷫆t�����k�6x1(C�)� ��	�*!�j n+zy�@"Oj��s!� p�5��ְ�T%�Q"O�81파E6b)q�9(�4�kQ"O�-��.ΆZ&LT�}��U�g"O��� '�wj�²����8F"Oք�6�.�*��؜��(C"OԐq�6�yF)zZEС"O��x���!L��J��Z���p"O���p��=&f Adb�w���f"OL���A?:0ha;�c��i{�)�Q"O ��oX�]��<�C��:9�Hy�P"O�|���	O�8�c߾n���yw"O�遥��C�.T�g�Ό>�xf"O`�H�B
39x���H��t��"OX���-�68��B];H^�"O�x�pgC!n�V 	�CʰTiI"O�] GㄚJ����U��i��"O�$��\�c������)���4"O�Qy�!�'I� U���Y]�t`2"O+Í�;C��Dg6����"O
���M�9�,ܐ𭀻�|Hx "O���cD8)¤*���\�T��"O��±j�%b1<�{�j��Mf2��"O�	��i�2gbtY�L�Fk3"O��a�ތ{	�������H�8��b"O��x3+�Rw�L��Z�s~�YX&"O(�seMٖ �B�BaB� %��a��"OR=����,1�K��ŘVX- �"O8T�ՎK%Ny�5��䄨p9<=Z�"O
��ꅰAD4�z��S�+
pa"On(�S�:L����!	8��� 7"O�@�
ɽ7���x���Yf�k"O��藠
6�T��6Ep �"O4�󳮜�JIĸ�w,�+]-&!1�"O�\���\4J_�W�^�#]ó"OB����>/WN�9�,��&x2#A1D�|Js�Îo\`�˗�8a�TX��-D�t��	����d��`��1Z�+D��'N�RA�YАg��T� ˵)*D����T�2��礃�l�����(D��)V�3}�l$��hC x��`E(D����A��r�3�\�#� p��(D�����Q�i�>�k���:�zq)5n%D���1��n���
d�9$���-D�JW������-�H��(���-D����b��y�6᳖��h�hP1�O?D�$)1��2	�zLZcE�!�|Š5(?D����P�e,|��!R�d�zq��=D�t����*q̰c�
�%]��y��<D�|���45����������:D��7A��II�����[$����9D�8;���68u����3:�k5g)D�Y ��t�ְ�¬�<fQ��0�:D�|ɡ��.�t�$M��/���#D��xujɈN4ܫ��[�d��4�R� D�T;e���,c��)���cP�>D��Z�-T� �T�#3XP0�!D�8ٱ�W	�Չr`V�uzu1��1D�xB�F����U�CZ`�Q��3D��r��ڗ>;ne�fL՘GU�YZp�6D��C'O_N� �̔���M0u�0D��;��E*n��Z®ђ���@<D��Y�)���H,P�Q���w.8D����%AB��⨎<ƀ�b�;D�� �̳<����/<0V�\�"OV�$�#�p��͟�NFJ�{"O����{!^�[nY,eǖ�Ce"O��ᢍ0t_���Ae���#u"O��f��
ٞؒ��Uhc^C�"O�]�i�/`��"�HX�,q�m�P"O($�iH�E��y@���>7P��""O�!B#H�W7֍k�aUH�8Qa"O����K4>�
y:��\>���g"O�0q�	{�d�"����+xx�"O�!����jk>y�㘌}�:��"OȘR��tL�"�a��~�쳥"O�Y���[dd�j�a�!=��H�"O�8�6� �S��z���!"��q�"O\q��*�8<[�C�Tv�!!"O�	2�
;��A��c����"O r��.6r���,�>���Z""Oq37�@"zw�}@�j�p�b�S�"O���� �9�.��(��޽��"O�8�2�UWu�`��L�(7٬�j�"O�Y���E�0���O6�^� �"O>��3�M"}�N$��m����"O,)D���xAd���ǂ��"Op���E��W�L�ci��U�p��"ObD�aL�L�z���U F�y�"O�q�K^=pO<���ܲ.��W"O,)Ss�P<_�,Da�7+BM��"O�����4/�:;�տ<�0��A"O�ܺf$OT�S��Y��|�"OX�3*X!�V��EV9,���"Oz|��K�b�� D��X�A��"Ojt��3׶��AB��w"Oz���	T��pA��r� �"OHX� �ʭ6hJp�r���@��:Q"O�]�1�d��u"jv�y�"O��)!�^�q�t�����A"O�(�"D!z��i��C�6��Sa"O��ӇF�#qp��C�̿@�Z�iq"Oΐ@�DT-V���s���4)��̐�"O�M�c�R�?q�(4"��0�(	��"O��R�aĨ&,�X�A��<<����C"O��P��I�m<�[B틏7���T"O�Ԁ�F	�xW:3���[�䨦"O� b�h�1]�|H�l��)t��$"O� 2�'x8�Br����'o�j�<�nKTj1�A'۸'dD@�W�A�<9���:m�e�B��t?�,2Rf�A�<�W�Ʃ-��YIQ
�Z&�av�}�<�!�IgM����ĎC��KVgv�<QuLC<��,p�49�-�r��z�<Q� �"d�B �R`��#*T�<�`�J�rb�D�"�M���j`��_�<y�fQ��DE��F�<$�fLҤ$�^�<)�F�>���1'��Y[xE*��V�<���ڤ����Y�NY�����N�<1��N�m�4A`FO�)3���I'�q�<a�ID35 ��VKJ"����D�b�<�	Ծu<d�b`�K�l-���^�<�C矚]�TQѥMΉpv*��e,�~�<�a��,}�,����̉!��2�)�{�<�cR%/��a�"�ڼQ�0P� .Tx�<�6EU��~<��f���ybH�I�<��D�$H�H�r�®~th�G�]�<qA�Z�&-!헬 �̱� J[�<� x��K1M�!J��9Gnm�"O�Tۤf��!�̸@�<��b��>D����9Mf������x��C�d*D���u�   ��   �    b  |  �)  B3  �9  =@  �F  �L  S  FY  �_  �e  l  jr  �x  -  �  ȋ  �  ]�  ��  �  %�  f�  ��  9�  ��  ��  ��  u�  ��  *�  n�  ��  B�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�VO&}��a4/zY;�#m�����#D�D1���'�01Vo^w:,�U�!D��1G�;(�x���n�$X�6@?D�P�$�Õ�ha�v�C�y �a=D�t�+�p��xj�N9N|�C�<D�:�K�<M�N<ca��*�Ĥ8��9D���������%� .�7Ẕ��<D�L�p-��h�u W$�[Ri<D�������e��E��V).�&9D�T*� -5��dKq�߾{|��聥*D�\�t��J�9��D,~|qR�&D����O�RtN�I0�6S�L�jUC&D���f�a�R 	!�j�T���$D�d8�FD�p��a���t�L�b��&D�|��揺-����e�˳I$Z��A�7D� �Q��,YX\�;5M߾[~X}��5D�p2'����(��R�,�^)#��2D��"�V��V��7-V,�^�QEF#D�(!�c@�x��V#�FP�-&D�\:�英B>��aι�m��#D� ���9SO�ؠE�l��В�'D��x��̎j=*���?�J�A&D��Z%��.}> Jr`�89wQ��N>D��TBԖoƾp�1���HIF	!D��-�$[� ��T���p`��1D�d����S�����K�,t���h%�/D���Cn<5TP��޽2�x����-D��[#.1S���g]�?�d�Q��,D�,��'i�踰�E391`�֢/D�@�OH=�)��ƀ�M��4�,D��8V"J�Rxv&� +�4U��*O6�E��#Y���d�Ѯ8�*�HS"O�H��E�<X�b��hF�U"O�cQ�0��s�;-�q	�"O�P���,�.�8qe��N�% �"O��HE*UR�����]U�T#�"O���HIi:�֧�\���"O��[����d�@��2�"��"O�kҎ��.����o�-|�Q!�'�B��P��B_�TQ j��G�II�'<VEZ&��9/<Փw�׳*`��I�'ސ�������Щ� /���
�')�9�#�W�cp
��
тTx�'.ıRV�A�Ws��id�D�o%8���'�΀UBDE7�³j�����'�@	�W&ŬI���K���-!س
�'qPȻ�+Ӽ	��E��
.�R�
�'(�D飦�"�`5 W:�U�	��� �<(Ĥ�
N��Y��KUR��ۣ"OvtSqJݲ>,8�&��w�2|i�"O��S��^�@�
�5/ɬk���2"O�X	A� ]1앪1���
1�(��"Ỏ�F�>�`y��-��He�'@�'2�'R�'���'��'N�
 �A"t��I��޵R�0�{��'���'B�'���'���'��'��������)�/��{jP{Q�'�'���'�b�'�r�'��'�Qid&Ǹ Ub4�^�l'邑�'y��'�"�'���'Cb�'-2�'w�td(ګ6���I'Kx��G�'�R�'���'���'~��'A��'��%�B/�K�lX�5�!?�.8*��'�R�'�2�'���'�R�'�B�'�V�A���mО);�,ӎz��Ybt�'��'���'�'���'���'��Q��L1�tT�����.̋W�'�"�'��'2�'���'���'�N�Y�D�%�.A9 ��k\T���'���'	��'�B�''B�'ab�'���4��%%%�!	vMIx�J|��'���'�2�'���'3�'�B�'���X5 Y��N�3ӭ�`3x�҆�'<B�'�b�'���'���'9"�'2�p��f�_��Y{��JZ,����'rB�'���'r�'���'P2�'|�Ju�ݤi!����늏"µ ��'x��'�r�'X��'�b�j�����OtUP�GN)J|�!r�Q9���`&$Ey��'��)�3?Y��i`� �*�Ɣ`�@�,kx�С������O��<�'��A��`:�#M�Ι��l,[��'G�����ia�	�|RC�O��'J��}�f�<ܴh��FԤk����<����$,ڧ �ԝ��@^iۺ9�F��!\r����iH@��y�i�O�.�rP(�{fb��Xz�X���O������O�	U}����b��F7O|*ĩ�3"�L��D�Ew
�H�9O"扔�?Yt� ��|:��k)����� t��(c'w٢��p�X�'d�'�v7-ږL?1Oq� cH�GԸ��`�2r�|���0�	wy2�'*b>O��\"&!�2,[p?��S� W)�+ ?a��Q���NY̧Q���N�?A��W}~P�&Lܼ3��Jb#����ĺ<A�S��y��!�9c6O�3qm2��b(�y2!r�Ft�4��h��D��|2�IU80=x�h��\�* �	���<���?��-)ݴ���i>�0��U��u�3��O�E�5������K�=���<�'�?a��?���?Q��ۧJ(<�pwc�"s�h�ivD�;��٦�RM��|�I柈'?u���0Q 4��@A(�)t"�:*~D�'�7��ᦵϓ�H�����eZ�8S��@��jx����6Q�d��X�����ç&���I�Gĉ'.HʓPL�y���Ig>�ˇ��n4�{��?)���?Q��|2-O�mo�0T����ɽr]��6������部��;b��������?�+O��m��M��Ee栙�J� OӠ�Q$��B�n��+�M��'@��km=\b��I%�ӽDfk��-2T�PTm�-h�����l��j��d�O|���O���O��!�S�A��0�Pȏ�w�@��C�*0Τ��I���	��M��F��|Z���?qH>���~�6T{�Hξ'�\l`�R{��'�R������Ni�v��싧�R�(wL\K�E��;�ޑp ���(<���'K$&�0����'���'�	SE�7Z�(Y�F�*l�Ea�'tB_���4h�������?A����]�75\\�bh�n��T�FM��e��	P~��'��f�:�T>U��g 8y`ezB�� 6[�ѣ�]�&5��(��'�P��|���OH�L>!��N4
`���U�@�9�!eL(�?����?����?�|2-O��o��HH4m�qϚ��`�8�^:���PaFyb�'��OZ��?q#��xy�B 0�T�c
"�?���i" �ڀ�i]�	�L�P{q�O��/b@' RnPb���K�ϓ��$�O���O���O����|����5c���V���m�(�����ϛ&*��V���'3�����'��w�l1��g��H��I3I	� ���'���:��)V!ch�6�e�����	�7`޴JeE��N,x��{�M�US��DQ�Iny�Ob��j�� 1իS�Q�����0W��'�B�'���/�MS����?Y���?�폦z䒘���M<:=����mߨ��'A�IݟT�	���L�b`�
)p[�IC
C�]�'�|3��\,���[����ٟ�[��'��y2Ԍ���$��s�T|��'���'��'��>��	3fA$X���B&�ң/��h�ɣ�M� ������O���k�a��Չ;�m��g�s>�	ޟ�ɤ�M�+آ�M��O �i�B�RG(U���jA#	<r�����.2�P�O���|z���?���?I�U�X�a�V�h鶸�Q�Y7D�\�j)O��n/\ɸ-��˟���u�˟�ңˋ1�HP�E��iW�I�"�KyB�v��Do����S�'�^}��c�Pp�3��/� <�靤);��'Z �z�ES��L4�|�U�xc e��Il�9b��M��|��%n�����i�6��O6�4�.�ep�6��/-�BX��2%V� 4�v`O�$f�'��OV�?��47��O�|�̜`gBC��^�y��!�sW�i0�$�OH|��b���������� ���4b�.v>:ak%"ScZd0�$2O4���O`�D�O��D�Oh�?a����P)���%N�1	�����Ɵ�	�hڴ�j��'�?����;&9 â	"���S��3{������x2�'v�O>�I��i+�����w�R/r��C�YQ�z��B�_}�R�K{�IUy�O��'tK?J�镊¥`����u���'��I��M�Q���d�O��'V���ua�`t�:�I�?i��u�'[�ğ��I���S�4I��Ӱ�k�'�%�6HKr�"g�ԩ������O� �?u)1�$ˊ}���3V���;�%�f ���'mB�'y��OH���Móh!tTL�F)�J���#!H�|�NZ/O��%�	fy��p��#pUc�:��U �80�V-iv�����Z۴�ة��4����9����'��S/Ns�PC߉Ch \ �@��6��}yb�'��'�b�' �S>j�C�"�\,��*.���xY,<�nZ�^$��꟤��b�'�?�;PX)�ɏ��5#�
��7�i>67�g��֧�OTlP��i����o
���KKd'�Q#��\���A�����!�B�O���|���yȤ���F�N�⭹��S&4�v�����?y��?�*O�eo�S�Ԍ�	֟��I!#,e���@��
�2p�P�s#��?q�O(��f�J$��1�A�!vÔ=K�T(��08d9?Q�B)=�~��t��E�'0�j�$��?��ٴ�FĈ�=mpR��M��?����?q���?i��i�ONbf�� !���z$P Lp,rR`�O<@m�>[����Ο���F�Ӽ���Q��lU��m@�Mحz���<�r�iҺ7mæ�	s���e�'�`Ye�B�?a*"�ʿ#h*5#��:<vuځ�A�T#�'�i>�	���	۟<�ɷz��A�@�?V�ش�5!|�N��'��7-�'@��$�O���>�i�OX]b� r_���e��B?�9��<A���?YƜx����5w!�͡�nH"%FA+��ۼ"��ɒR+���]�QEջ��9�ԓO˓8�8�@�W rE�RVog,�����?���?���|�)O��nڧE�\���2� �d  �P[#�Ӝ�$��	��8�?�O���d��pl�%I�Р��И|�l4�f�E�Bl$9UJϦi�'
�$R�?Q�}���P�H�s�ҖJRz1q#�_SwP���?����?Y��?����Of�p����YNVHq��J2e)�Zٟ��Iџڴ`��D3+O��� �DѶ�D*W�ߣ:�QQ�HH%he'�8�����!H���mZ[~�h[�����李p�f`�Ug^�>���Z��̟�'�|�X���՟����D�D�G�=,��c"T/4B�43v����l�	by2�r�A���O�$�O��'j�z�xw�]-y���MY)�T��'i��M�g�i��O��H�eꎎO�bAx��!,�}�t�=�ʴ�4�-?ͧt$���P���*xU#�-

�V�H�KR�؍k��?y��?A�S�'��Fަ�p�[�}��Ѣ�7]@�D��9���<��p����O�űG�55�J���D4`�B�ODQoi��m�s~������Sc��H34���ǐ�Y�Tѩf�ȦG��D�<Y��?���?����?�˟�hE�V��.����̫x=���AbӨ��#��<���䧎?1�Ӽ�A�-"���֌I,A�=�tO	��?!�eω����'��$��o�F<O�;� �%+]���3�6X�~��b0O�\2ЅY��?���'��<ͧ�?�`.��Q	�5�� ���(H%��?�?�cυ��?����?a��LZ�.I . ���O��i��|��ޑx��9YW��DY����D8?���Mk`�x��@7����B�R�nX������y��'�*u�V'D�=�8݊�O��I��?�]
��_�M���&gV��)i� �'m��'���ǟ�H��5l�v1蠏J%h]�< u@�̟<[�4n�U�,OH�9�i�Ia���Vq���yZİA冡��lZ%�M��i�@���i��O�s'�+�j�LĒi��E%�	�Ԗ8z�T�2�|�V��S��`��ݟ4�	ϟ(3��K7GIFqA]�Z������}y���*���O��$�O�����dD[��	K�#G �����Y�dp��?y�4cSɧ�'q\}����i*P�0�J��N'0 B���1��'�N�BT�ş�!#�|Y�@3�]�t�Q�D'C.PZd�F��I�� �I��Dybil�:	XVc�O$Ͱqi�
e-T�0ʔw�\�`�O�$4�	f~"�'Ǜ�)f���U��ou@���C�"o�P%Ǝ�H�7-5?Y�`;<Et�i;���iʐ)I�.�j��w)F_�h��z�`��� ��ퟌ�IڟH���b�#�P�#�̅���
�3�?A��?1�i�رi�O)R�'%�'c�A��̆9�PHRX�rU6Oj�2��ֿ�\��\ǖ�n�w~�7KKv���R1U^t(j��I6J�f�C���ꟴS��|�W���$�	ҟ(��WrS���!+D�.�� t����p�I@y��z��z���O���Or�',e�AHЍav�0�!M/H��'X剞�M��iE�D ���_����n�͎I�gA��)��/7������ˁr�i>��՟4�0�|�i�i�,QH݃xK��W"]6w���'�2�'e��tU�Bߴ
>�M0o�I匁3#�J��Dkt���?���?���V�����0#�7x��%�5e`�x�	1�M��ʞ��M;�O����<��J?� �%@Ü�?�|��+	��X��6O���?��?����?�����I�,�$d;��a�F`���NRx�o��)z���ɟ��	I�ɟ��i�����)T��ҁg�V�����(�	��Şk�i��4�yr	]�e�:9q$��C�b	��\%�y⮓GrLD�ɑ��'v�i>-�I�3R 	jgꝧN� 2�S�^�b���p�	�P�'�|7݅/g>�$�O��3O�d<�!E����w�N��?��O���d���&�,2��J�]��`��9j��dj(?�"�S;I��c�i�g�'A´���'�?	�T/,���Ƿa�&]J%V�?����?	��?��I�O����X�h`򂎎��\@�e�Oftm��I\ܕ'�b�4�|%;3�.f��E���2�::"�Oj��x��mZ�'��ul�O~rL�L		���q�ViX�B@���yG�Hnm"D�|W��͟ �	۟��I�l�@�4,U2L�3#O�w��0� �WyҠe�b�����O��$�O4�������>�<�� N&A�ؕ�4��*\�ʓ�?a�h����O1�F^�~�*�84'?%�5�s�N)"��1�OL�� �?IB6�d�<s�PI@�pp�Z�y�������?����?q���?ͧ���ň��؟dZ��qn�Y7.�*�¸s��柌��[����զ�a޴I�����'LN=��h_�
�ҕp�B�=1�y�u�iL��.
-�@S�Oq���N�:�F�sE��t=�V���<m�D�O��D�O��D�O�'���~K
9�(�\��X�%}���I��	 �M�G�|Z��?AL>!)�t���,��X�U 8F��'�z7�����o;�lo~(R�3.v��f�LfO�|rRg��~B�6��)h���`��'t��͟�]NR��?A�Rp��mU������˥,]���%�H���?��B�@z�����ɔ����<]�Z�ZѬ�g�l��O�1�b�	ǟt����d��ğ�Jٴ\1&$	(���$˩d���'M� @�h�&�{u��t�]")��(ԓ�(��EW����B�'zU�gi�e�ێdɎR�#�1�?q��?���?i4GŧDǌ5X��?��2����j�)"����&�@S!R�T���O���3���զ���	^���I�!��[�O=���"���Bk�˟�Jߴ
�� ߴ�y�'��9��Ǡ:M ��O ����ܼ?Θ����i�"O���%!W%=,�A+x���B"O����a�#Czhk�����%xR���l�t!��h�MQw*]�1��q�@c�)W#*�+7��c��Ÿ��� ���d���h03@AT�2l��#�m�x��q�@	4 l���0�N�)����8�s�BS�.T�\�0o�l��Zt�C�2�㕮X�"�p�[�6r�C�-%�5�v��)�2��%-�#lC�T��CK�'B�ҍˢdY�",v�`dB�0��	�4�߽:f�����Q|^d��I�-^�m#g^�6&U �fG�PF�P�0j�qIB��ee����u�%e��N��ץ����ގ�J��	��&P�'�Fn��) l[�Nz�\j�ΉJ��ɀ�}��I2D�8��^�qO\����چ5٦�{5D��B5ʍ�R��[��U�)�S�,-D���p��*�D]S3B.
p��iFA+D��$��\M�9ѐ&Ւz��hQ�*D�DĬ�1IǞp஖�9�yQ�-3D�X�������X�!n�3%�8Z�
-D��Q��D�	w�H�K��� "%?D���V�H+DA�`��M�l��.>D��*� _/i�E��&H�5o�(��<D����k9[�i�c�ӹ55&<���?D�����&d�:�*�HR��-!r�!D����,B�HHY�M?9�έ[BJ:T���D��P��h���^02���PU"O"��@I�|f,���܊330@"O���'!,~�Z�dG�[2$p1"O %c�bY�[��$����/>�:!�b"O�ѱd�0i���uR�c��t`@"O���
S5�2d��m���c�"Of�)�,�/|x��`ކQ���p"O���s���d�xdE^.w����"O~Y�c$C�EPj���@E�>`(pB�"O��#F��>��}�7 ^S^���u"O���ۃ}�	hQ�߉g��I�'���q��EV^,��L
3�
��'YƘ��	�f�J�C���3��99�'���ao�5K��j5��1��};
�'� $��c�m� ʁHȗx��\�	�'bB�8��=�����4:G��	��� ��h��HN.��#�<Zd��5"O�x��%��2�Y���4_WT��w"Oh0�!U�H>��gGD�ei��H`"O|�A�lS1'�"�
�H-ޑ�"O���*�vq��Q���:�x�f"O��(��8J�q�$��@(�x@�"OTԋ��Y$O�\T?~�x4`c"Oȋ���F�a��k߶y��3�"O�٨7As����
�F�*Ò"O�E�¢�:P��;JI+*�n�Ђ"OX\Xo� c*lT	C� v T�X"O��DN�E"RX�@mZ=.���2"Ob<a�υ� z�1Į�8�:�'"O:M�@,�J�ӂ���̠��"O�Xi�F��B�l!6�E�1���e"OZ5�2� v�8�B#2z����"O�[�
�Ky.���C�5*�,R�"O���!a��Z�u��	6B"ObEzClʩf�T8RLJ�$]�5"O8�z�F� j���re-͉4�ƥ0"O���k�M؂x�5�K�Z��!�"O�dA�MEL[�M�"���zz���"O�x7�߭ �ƱY�i��9`��`"ORx*p�BLl��
��k���b4"O�mbw�5�>d[���9�N�Y&"O�$���^�l#K��8�i�Q"O����G�e�Iа���u�Z �"O4x���[��ؠ��L��,a´"OΙ��Id�P���;O)`=�"O�=�f��R����	O�V�
��"O�]j�G֊<�X��-"����"O"����0|(@ F\"䠀%"OI�ѥ�8\p9!vcܦJ6��s�"O�)�K�%J�RL�B�,nX��"O��â����'O�Jx8f"D���`�3��H�G*̫q�(���>D�����G"[S�q�`$ʾ,E@q2B;D��c� n�
�C#��31���P�D8D���#M���܋�B�U����N!D��a�)f�����L5Z�e��!D�|��.B%<��S�ꈬx�0���=D��Se��#"�mCq�2�V�68D��2�(A	O{�|����;c����C)D�1���`X�ܙ�b��Hж�z!�4D�L�LF����3eE<i�ޝ��.D��!�A>F5��I�-W�{��)C+D��97��=	�N�(ᓛQ�D�҈6D��P��M�o�lBfH]�A��
�5D�haT�M�?�6��3`��7p ���3D��X	�"�f̣���:Y�څ;�n3D�h`ۼYqd��2(Ŭv�Z���TJ�<A���.
-��Y�H1$5Vy��l�O�<�'�q�^�AU�ޭDÀ��ML�<�MA�

t��&9�1���H�<��ꇧÈ� �*K%���#�
i�<Q��M3��*v��4{z1�Q�]f�<Q�m�t�� 5�����P� �^Y�<�wJ�2hX�"�Tk�d%�T-^V�<����J4�A�7��3aD�ٺ$�y�<9���`�ly1���� �
��u�<C��qt�SuU> d�X�PLk�<���9M���[�|�P�Q��_q�<��	�rÌ1��6z���Q��EU�<IǦێ^�&�X6!�-���p��O�<� T�JB'X�+^��dQ�,I�@r�"O.MA�L�E�0h�� IH8Ĵi"O> ;�k�<7s �S�E
�C$- �"O�ёG�>{��a�v�Ȋ�*ܛ0"O��ڰ�8w��qa��[6CےA�w"O�]p�"[�_Yl�2�bH
^��"O��1�ϨGR$��@�E�)�����"O���"�txF�Q+ݍx���"O�ԛ��^_�jƇ��J00r@"O` !�:obzyr� е+D)��"O��#�-A+dA���nF
W�-��"O���W���qF����mh| �"O��x%OQ,;��m�AI�P�j�"OLI���}P1B��\�2E��)"O�e#����vp ���� V)�es"O�$��%�%v���Iط}z�X�"O\�i1g��&l�����^�@ȁ"Ox�B���b��Q[�w�b5:�*O��(�@&�j`J�rKx��'z9�G
�*���yg(�;�9��'��mIc˚ |�\�f���5�؊�'���P��L.��G�<����ȓh>��J�фG� ,�7-<�<�ȓC�Z�@���'?� �q־T��ȓ}U8AW�4�J}�2�S7$�2d�ȓx	���_��D�����H��؅ȓ\wvQ���ϰ�6(��'<[�N,�ȓI� S�����9@d���ɇ�^�,�3/�;B�,�Ӥh 
sHR�ȓL�� H���4f`X07ꑃlA^��ȓvn���� �gȄ�f�ת���D$����L�_�`)�B�t��%�ȓ9O�����ߠi�����Z�K�Ĭ��~�nժ�Ő�DY2��ğ1w��ȓv��Ps�!�ɺ�/	!�|��E��j%�΋{�j�``��G@Q�?�@3,O�pr���U(C~�ҽ�On�+�B�'
��'�	�R�%1�d��B�tB��+Ho���h���ܨ�G<3����$�$���<��BOf
ze���q!�X�<i6dW�L�̐�MO,K���i��TL�I)j��?�}����^�<]c���bDnA�҉�F�<AQ��3Q2$aH"��$.��g�[�A�|�q���2W ��v���x�"_7C����Ɠ 2� [��ͬaP���ώ�b�Tma$��e����ܪ-���sA�F�e�4�EN3Ű<��ν�J&�(:��2t+�M@HL:m��-D��{c��5_��pc�v�����7�x,�4A�{����C�z����Ls��Z4)Ö�y"�-��d9�K+f��X"l4��' 	�9OVQ��̘*h<l�x�ҀzBO�0�F䓦/����BC�$~���4G��h��C���0�Aǎs������9h-8U�剾}'
��=�ͪ>F����K�*n� Ӕ�j�<)�'�����&�;p����Q�I� j0�}��D�]����Z�p�2��fdɍ�yR��l亡I�#c���P����'��U03�3O��s�̈́^�5(��H���rO�q�O��`�2�~�����a�2�pu��~��8HFM�`�ej��\�b������>PqO>��qK��А%
��8;%���y��"c����S��Д�й�yү�v&!�s��97IB���C1�y�,Ҡ}�P���ɩ6K���OL��y
� <���V������4��KC"OB�bاjiX�pA��cP�� �"O �2%B�5r��1���AG�g"O�eiv@�6�ptr��ܼ55l%��"O�!��/�$l�� ړ$Zu�"O,�Br��9gL7��-hv[�"O� `͙�I��5gX�nHJ�!�"OZ�i�   �l �eO�%���"O���DGۂn:2���$H�V	��"O���o���D�n�"O�,a�[=p՜�����"H��"OR�� �Ɏ�J�(v��cҤ��u"O��� ���H�i�����"Ot��V�s!�MbvkU��Xб"OV|� ��!O��e��D�/_Ў<y6"O*%���Tff��W$;�J9$"Ol)ҕ@C)WM(1QS"	�+��{""O���T��$$ \��?�<��q"O|�36/�w�T���*s��R4"O�
�DV����1��ܘ!��)�"O* @A��-N�&���@�4AiR�3�"O.�
/����oB�b7�4Ya"OD1� ,�&OXi+�O��d̰و%"O�5���#+�r�;�Q�t�<�3�"O6H�及,Y#Bݲf����+#"O6�[�%�7Z
$#��
=;�i��"O��x�`�8@֐�1�M�/����"O�uj�/�SGl��e��>fp"O�]R��"fCꙑ�dݫz�:��4"OIHB�ޝ7v~���T{211�"OJ�{#��=����Ꮽ/�H��"O��8f��p0ѣOC�*���Y"ObtH�-V��y��ْ>�:��A"O0l�Î
 ǌ�:TÂ\��X�"O�����
��
_)tX�Cϛ��yr�3�%�6㟎W�8TSoV��y��O(c|�[a)S<xk`����6�yb�
-?��!5��s��u*a-G��y2f� bQ��G�L�p?��p��!�yb�	�@��i�P5p.�H��,��y��R<}(����7n�(��+���y�.N�=<e�wC�z�n!��ق�y��5�0i�@�qז4��!�y��V5jf$!5�S�\.�PgW+�y"`\�o@X	!�Y���!���]��yJ�>��MhT�Չ0��u*��<�y��\!����4.��)�� ��ϛ�y"@I�W��q�bַ�^������y��Ж	�f����R ӄ�L��yr�K%���@B�l�T��G<�yr��<< |���b ��.H��O�y����푅K%f8���eլ�yO��n��(b��>uU��c2�M&�ybeD ;h���� 8mJ��$&��y����V;�lC#KZ!d.��3���y������!	�0,-��Ϟ�yBH͌=bT�)�F"���v��(�y�Lنi�uB���/W�m!����y���X���#$G*f��`V�y��3=�}h���(�jZ��4�y$�*�v��B�I5�VL���@��yR��"a�x������)���1-���y2M�
N� `�o�+*r����J��yGQ�G<Z�J��Z8��0���y
� ����O!o��ia*̜0��]�"OJ��A⒞Yx��B	ʿf�<�"OT,�卐.6��=���Qhd�3�"O�J7O� _�\z��ƭSMV-9 "O��b 1 �z��'c�r�J�"O�X�ǫ�|��MRv�],	�\,i0"O�	�׉%�Vx�7���">lġ"O�a�dF1CP<� !��"~���"O"��F�"�.d��۵f���0"OHd�w� |G����Ȝ�^��,*"OB�A�C_��\-١�Fo�^l��"O4���046bU�7�C�%چ��Q"O(Y�q�H �д`#GL�r�F�V"ON ჈H�h�6H]�.�Z��"O�D��d��>ˤ�ё;�&�q�"ON̨3"�5BP�av썥�\��"O
�Ђ��s�i�Z0y��h�4"O�0�ШyQf��#t���"O*}2��K�i��()�
�^Ҕ��"O$�ʄ
h�����ϲ4Il[�"O� �C�>,]bt
�#Z0ٰ"O��k��$5����k��a6���"Oة�����c�Ԕ�𫕺&=ʵ�""OT,�Q��0���n6�щ�"O\��4�ȼHQ~)�@bҜc6()�"O�����D�*�BG>;
�+r"Oj`���v�x1i�ҰB$(�;`"O�1p����j8"5��87�e�"O~���Ži@������:/��a"OV{DO	W�b�F�8or�`�"ON�c˓N��ūs�F�
x��"O�Q3R��3n��č�x���"O��u �&n�����E�و1��"O
�#�L�D�R9�o�3���h�"O��C��I!Yl\���Ң!��\(�"O<w��o+Hy��R�
�^t
b"O8�Q0��+6칀\.�1�*O��*��X|�-�@F�;N�{�'p�eXd�Ҏs�!���1�� J
�'J������|���Ө<�V�	�'r�x�cG�X�� #���0�h���'jtA��P!�"	�Um�"��e��':���ញ$X����lU2���;	�',|��7�M�5b$8���'��-A���V�U�� �6kJ����'�eNN9YV�AEB���,��'�ֹ���|!���b-޲�i�'vص3%�hǤ���6h{�l��'m����숩 p��QŌ�3dF��	�'��� c�J�i����>`�f��
�''�R3AC�� i�@�+� ���'5� h�GHP��E�N�v�l��
�'��A�&eά"4�Q�9�D��
�'�V �$�
�V����/�&aP
�'E���K�t&�X�ҍ�>!v���'f���N�A�B9��'M�2�[�':�u�v��/r~������?HX���'v���		�A��4��[ NeJ1��'���p�܆Հ�)�i�G�0!j�'{\�I�O�<bߪ�ۇf�1G�!��'�8d��J��4>��W�8�R�'��<qG� jˀ�PE�L>Q5j\�
�'@�	�t !g� ���D�#af9�	�'�.e�S�Yhֺ���(��Q��H
��� (܀w���H�ք+8�`U�"O��3H��8HI���g��+r"O��p�SgC�EQ���}~����"Ot9� �݊!9@��ra��\$��a"O"�c�J1���P��3@tlJ�"O�	����0dj����20�Ձ"O��IR�Z<xB��o����c"O4�#D�0V(��㊤M�h���"OҨӂ�U]�F��b��b�~�(�"OdT��!�b�R���[��\@�"O��4Cbp�3'��2?{���ȓ���2�)ȩB�FX93(��-Hz���t����F�0m
��8e�@�n�6���h9����i����u�uS-r��ȓ2�8���Aĉ%r�h��8d��.@�ه��Z�ҁrQES�K�Ḋȓݰ�*�	N�O��0��0_�`��ȓ��u�w��'l9����* ���$�ȓE�=�@��>^��b�ɰ��`��OD}`�I�O��Q��%?�|�ȓj�-Ζ)�vɠ&
34�H��3��Ti���6=��b�`ės}�̅�Nk�����I���		Ɛv���I� 1)���+q��r�A���Ą�L�n��F�!+,��� P�Ȇ�q�Ȉ��CŀXƐ�g6+�̘�ȓDF��:�4g�U�1H�0,6�ɆȓK�4#��:VI��wCҮ7r���f$�]j��-�n�R$�R�d��͇ȓT\m��8~d��BT�H�0�ȓZ-�	�Bj�/C�X'+Ř`���ȓ��}�P�!Nr�J���6�v��ȓUl�����4^Ȣ���K܆�ɇȓ�m�ᮇ�<�6h�%�+Ha�|���6��j��Dٞ��7��d�4$��5:� aPV?@�a�C�
$O:�ȆȓD� %p�&X�6NZ�0C�;Q�Zp��4�fܫoܲd=��l�
m��U#�'�hd�!bN9Q1��<���',lD�p�U9p���qR��zȉ�'t�q���V�����P�{�z�9�'>�#%�R�5�xā��={�����'ي�bTD�c�=���r�\q�'�R�����-)�P�)�唝t,
���'����F�]80�6�s
��e><Q`�'Z�!��_(`i
���eA5]x���'�N���U�(G�P�B��[���

�'n��u�^8&8��eT�h���'� $�q�����o8f�X�'��X��Q8x�~[�.h�PQ��'"`Y�N��v;K��U�غ�B�j�<iq(0x�R��&�z7@���_l�<�g�����tꏀdօ�D�WP�<ipa�?z�z�*�댹�8XB�V�<Y�씘4ĭ"���5a�8
� ZU�<�'�H/Y����ώ.%�b���O�<A�D2�����OձQ��M��B�<�q̄�FMbq�w�\�����FG�<���(\��@�J���9U�ߖ%!�$ūf��@M�%g��B�c݇>�!�$���Uc��M5~6��R�e�3t�!�C�Mz�$���ͽ(�\�+���!�D�m2l�;ԆM;Ant��©�?!�X<<�d����֏kc�8ȕ�^+�!�� ��VFL!�؄i��L�}Yv��"O�\Cr
���ɂ�DYH�����"O�@�$������&C>#�0<��'�x�3t�_�5?�II��T�]Z ���'�A9�^7���Ջ��j`q�'ΘYS� _�(y�#���x�6@�'6�bt��9X�2(�L�i���
�'f�m��h�>��BC_�3j��;�'�l�;p�<Rj�Dx���C<���'g~@�T���s�$�:��<��89	�'������|z��V
a`�%8�'yPh��L,tmNɻB�L1�J���'� �h6�4���2)C�3�8!��'F�a9�ҟE�x�VJG��iI�',J�$傴L+q��J�,D8���'*N�n	��!�\!��C��0��'�i�J�-��}�^�O�0j�'�% W�V0W˦���
ǐM�p��'����%e:��d��Lpr���'����-/�@	���R�KU����'�� ��FS��i�R�D�q��'&c�!�)U&��g�/@̙֔�'�
%kԏ֦/a�Y��6���2�'��Aԧ$g}@�8�ߤ;F���'.X�� ȝKkf�3�C��$��'��(�蔤!���C� �#F@}k	�'�J��+I I��\µJ�7;�����'�Ω�0B-0t�����<�HU)�'���;㋕�¨��M\̩[§���yreߎc�P�k��L�<
�ؼ�ya/x�|9 �nޖ<�D�0��ǯ�yr�4�V͘�)�$?H`��y�]8$`.�8�fΠ_U��[��>�y�%�qh����0FHeivɞ�y2B+���խ�7���� _��y2aL�U"p�c���+Ln�ڣ��y2��D��(�[�*��M����y�k�G; 4�a(��(k<��C
,�y�%��~X��0��j����QJ�yR�@�`���3vc�j�:��I���yB�ؔ>[� �A牝Z>�������y�(P��@��CR�X�D@����y����J���s$� �X�ẻ��y��Vq�$��B�6u����dë�yr]�����OJ�W���/���y�	��r?p<e��%(���M��y��yK�@:g�Y���}�a%�-�yR�-$y �$����q�&
��y"��i�rh��j��A2y+���5�ymF9d��*Dr�vYs�#O�y�h��[��� �V'l�D�ٴ�ӑ�yc�oT�yXE��%j�,��D����y��@�_4Hp�L�c/0K�j�	�y�� �%`�jA[t>T�����y��� �F�bs�P7B����bgʗ�y�*�[)* �Kʆ�3gj�/�!�d݄Rh~��0w$�Y��Z�!�Ă >�cb�W6kl�X�P�Y�!�D�/�\	�R��-`�y:deC�P�!�$�*}�$��%� uu$��I5P�!�$S1jd>� w�Y��P�"�ڧ�!�d�"a� ӣ��7�2B���!��N!�#$ �t}��St���q�!��[?�>}��e��(zD����:cT!�� �c��A�k�dUp�I��A��A"OT�Kҗc+&�Õ�=-լ���"ODLـ`��0܄��g�H%nFlB"O.���ܓGH�0��pZ���"O�� �t�5sS��H����"OL�ٰ*F� ��Es����)�t�"OV��M
�a`6�)¬C�l��I""O0��a�m���J��?ݶ��""O�Z���Ű7����4�NZ{!�D׾#�=)��e>� ӊ�Dg!�ĝ	_f�����D��E��^�J�!�dT1<�-z�.@A'�ȶf�!�D��1�Z��Z� pK���3�!��`,����!,|ZfO?5�!�D�7���.tX���v&�)I�"O�ث��K�.�q!s�H�( �;�"Oū�h	8�5K�!P���q"Op,��̚�{
���Ə&x�Bqy%"O�h2B�5�E`B"���bi�"O¬�s��(�������{�"O*�s�P5D�����:m��4�q"O`!;�ʑ�h{��s�� 9�"O
���H!}I �wc�$F+!��
~��<f:����W�g�!���8D����#REYԂ�8�!�d�*!��|�J�Yg>2�S	dU!�D_�"�@�b�I4Y2Ĕ�"�L0!�D̗ �	���ۃ^�,�ۗ�҇i!�D��IzaF+K�e;��^�N!�d�iR��SdE�lhnqoA�pV!��4A�fH)E�4?^4���9_C!�DQ3x�:`�iE��˒��+a�!�Ā�zz��ü3[.��PV�ԊZn!��خ!���J�<5lD����>h!�$F$�21Q��$G���ڳlÏd!�$ �9K� � P2A���R6
�!�D�,T�T(���í���C�-	�N�!�ݹi.T�W�y�NP��l��.�!��B�x,(�KL)�hE�S�X4Q!��7f1�E����q'<�@�^*6R!�81$Z5�Ṗ0~�b Y#>L!�d<_x�˖,�9m�U��6F�!�$��)g�E�Q��<hj�A�� �!�$F2<���dH,��d��7-!!�D�_�m�P'Ӱp���aa��!�$JW�Q�s'�����%R�!򄉿~��`��F�2"�R ��!�ݒ42�T�@W����c��LM!�V�:$(`*]9&z@����:L!��G
>7(1r0�Ѩ����H7:<!�Ƽ��� 1�H8�bV��""!�䓁b(���'g��G���H��"!�G'
�<h��̇�ް����M�j�!��#j>� �B/ۃ}FYٖ�_�j�!��ɴ;X�G��<Ci��h%�^�6�!�3n(�b��ΨUJp IWG��Py"␽T��t*ŋ�$=*�&ߋ�y��H��L�ڤ�Ϥ^�(��T �yb˓+k�Ւw��'�n��N��y���u:���w��`Hb�R��y� @3�
\�CL�3Yv�〉̦�yRC�'D��A;����ـ`�L��y���#VZQ�is�p��W!�$�T1�T��oT`r���e��!�� Ȉ��㇈Q0Ҽ@�K�*
D�t��"O�X��*�&�d|����8)��kw"OJ��ϑk A�˘�=�9�"O^�u��3�RH��i�(9Mb�r"O|�y"1q����/W�?��"T"O�����}�n���58 61j�"OV5�I��k�*M`���.�kc"O���`��F�b%��.�:hp��
@"O�M�'	-"��+f��7CzF��7"O~�"��96�G�oj�%��"OH%��n�fM���(NP@�S"O�i��֓~�u�U�^�Oh�|� "Oz()da��-��X��Ң5`\��"O
��E �f���ц����"Ov�#��PPd��SJ��zS�"O�����X���1z�ƈ�zIB"O���$Ⱦ{v���v�Z�L�2"O>�Q���5�6�'��e��"O � �һb�t@�1�V\��"O������r�j����HR*��"O��i3HX�_����b��jE�isU"O�<��R�ʚA�`�!)�䙆"O�H������Z�����I�"O4	�P�� qč*#�I��ɢ�y҈��<H���$Tgn�!�M6�yN;DCҠ�R�W�A���)1I4�y�
�e$�	���7��L� Hͤ�y�d˫~2�i6��,)�`� )��y���Y�:%�2��P�`�PG��y��ٜfP3�ܹIp�㖌U>�y�_�*�"���B��"N߰\�`P��Y_�(r��Ƚ^_h�MO�"1�ȓe��[���Q}^D3����Q��ȓs�bܑ#MKed<��V�$`���[��`�v풓S�н"+Êc~@4�ȓ?���w�O>5R b�
.��ȓdf0� ��#���W	+���4�������g��"�"�\ �ȓ]�����!�?V���˃k�.��������k�	;�%Q�AS�Sb܄ȓZ\�ɸ��[�l$�MH�B!:�R��ȓCSإZ�!�~xݳ�B6T���ȓ_�1'��009IR_�2��Ʌȓc�����O����w:-��x��p�H5p���V���`	�Q@��e E�V`#|Qa�K��ȓLIF�#R�[
m�0�@����݇�@�PK�������
uG��q�"��ȓk?�Y��-ź�>)�s�F�[PZ���m��4��
�5k�,�a�L�[���C�"�y�W�R�y��N�d��<��BN�%�'m L�f$*4��%e��ل�k�4\CWa�7�A��%O$.M4y��RW�XxS煵c�I�!gK!H�T�ȓM)�\�CL�N}�4��Xr`��	�"�7.J	.<H�GY�U�8���&�}+����bQ�IC� ہ\�H���jO�seܲ�XE�vi�8�^1�ȓ1j�Z���x7h����1������� �@�H	*#�	�2
D(j����p�� !�*HKn(s�J=W2�<�ȓ=��H���H�dph95��?J+
y��d� 4�S�7߈Aɗ�;�z��ȓ%�T
����lP��V�j�����S�?  :!�E�<x���*�3��Y"�"Ot��"�������c�'
] �2�"O�@�O�8<xUC��;T��F"O�)x�N
`�a���8͑�"O�ѓ3�>I*��[��5��< !"O�ݫ����eބ\kE��/,HA[�"O���OV�s; 5�FI���\�"Od�QA
�e��gF(9r$"O���Jۮ/�(Pr�'_�mB ��"O|MpDE�l��f�!N�#"O�i���W�kr�Y����>��I[%"Or%Z�,2cx��W�Dzeᘍ�y�@�:l3�d�U�F� �"��T�]��y"��"� EHĉ�8v[U��䝳�y�ʈ*��J�I?l�2��bQ����hO���<�ňٯ����I�2W��q
�@�<	"%�:#Z�ԲD�ê,W
`*c�<	!ܦ?�6 ˶�L*PL0LCԈK�<�a�-�6��6��Sþ�`��p�<	nR�<��9�E��v&�P֤_o�<A�� ;�JA:��.-���Gk�<yf�!����-dN֬)��e�<�4�x� �B�U�~��E�Id�<��Ā�g#R	4 ��h��y!lZJ�<ɶR�7{HT1�J�o88���D�<�&E�b�\<y��PH��D���<�䄝�d��=��ɋ�v�� �#O}�<Y�D��d(�YU��1���p�KFA�<�2gΜ(X�@���-)�!r��F�<��R�0��@�#�'W
yX��VB�<!`
;^�x�� V��Ś��e�<���0i��gʃi��Ē�*�l�<�e��WtݑCL�d:Fb�e�<)fj�,A.5��mF�W��t��b�<a�ɥ[811��=�"<+���^�<�5� &�\kQ@H�A(Nqp�D�<q^zH�bv#̵U���ó�F�2B��"K��1�f�9rc�$Tč�VOTC�?����/Z������%���Yh<y�ՐnP�up"�^�gDu����\�<�G%HC�l���N�a�F�@���^�<I� ��1=��q�鏇_'Np����Z�<��Ӊ{�fC���w��y�f�\�<i@�@"b8����ʆP-nU�cE[�<)���w�@a��*�7�N̉�.�T�<�".�9�pU���{��Q�͎U�<qv�^�@�h]As�.�l�h�L�<��"%&C�eL�V��h1�I$D��1w쐏`t�-��A];)�8�Ej%D��"W��Vmr(� D�&*�̑�o#D���`�ϴMF���$U?zθG�?D�4�1�8e(��[@AD{�8���;D�Hz5(H�)=���B��*v(3�,/D������	9Rs��O�{TH�Ņ!D�,�E�BH���/Μ=T�*"D�(`2 ����)Fi�q����M*D��!�m��6�j�G
�
C ]xV(�O.�C��zC"�l���K��	EQ~e�ȓ]���JR��?>R ��Im �ȓ0�)9�jϡ%�2	� ՅFܔ�������ö1��yҔ
X>S�����s��D���ŧV�,�KE��^��}��-��DaōN}*�KЬ�i���ȓrU��3�M�p+��#�I�tm䀆�S�? ��
�!$�n�
���1C`0Qw"O�(����9�>ѫP���[a��(v"Or���.}��tZ!J<ZHr���"O�S�J������$�?#\�H�"O�����p3�4`��v'n��c"O�Up$LF4��<h �_�;3����"On��c���	�`�A���i+�d�'>b��;\� �!��{�a�D�O�h�p��ȓ2�2�����,�n`���=a����{k����!��Dm�%��Y�Av݇ȓ.��Q�v.��Js��Bƒ���ȓfe�,�`ΘB_ XZdd��ˢ���1��m����3 �0r�66�� �ȓ=��!�D�<� ЂAU�T;$���П�'��D��'d����+��q,a+��=�$���'F���n�+�*1qF�e3�I��'�c�Y�$61�D�LX ����']���T�_��*�E���y2�]F��ȓ��A�@AD`���yR��
3�f��1���$�lt��jS��y�CK/_�@�ʃW'0������G)�yB���R�Խ��-P%&��e�2ꈼ�y��)G��|(&៫%=��3�Q��y�!ħ#�BL:G��I�Ԥ�Ƙ7�y�˛�h��C.I<<9��
�
�y"�,m�fYId$�l�X�C�ݓ�y��O�f���)%j��Q��J�y�C&g2�y`��<75� I����y«�D��pS��!L̍��+��yÓ=Ҧ�CB� .� �ή�y��7P����ՆpR t�GG��y"��	�]�������OP2�y�!�h1��ţ��p���ǋ�5�yN��[� CG��sz5	��y���6�V����@('��91�]�y�$$�j�;1+r�ub5��<�y�b
��5z�&Jm99��\��y©æZ�J�[�Z�d�\y1��ُ�y⧓�N��9��e��I���qD()�y�'ҹz�V�z#k�42V��9%Ɛ�yb�7�؍���5\\XQĢL��y�.��/*@hJ�l�9M�
��yR`��5t��I�3=�t���U�y�O�d��z�I�ľ};f�\2�y���7EI�����M�P*�yb`܆]`�BjW�Ύě"�J��y"�� 7���a� �5���9�y2/���q�T��<Y/.-VDɜ�yb�׫�J�̭Se�R婕#�y�E�<y&2	� 'U�L�X����yB���_��Ys�G��Qc���y2b]�g�T�K���9�)顯٥�yr����AQC��CXVa�A���y"a���XܓD�?��2��yb��S�8���ܷ'�rT����y�*ِa���qh��"��4�vk@)�y�LN7����DW�(6�*�y�چzt[7��:9�Y!&`� �y�,_(z���9��
.�p�P����y�M\�u��{Ƣ�)�����y"ņ���Ԓ�iŐkO�=���L��yBi��|�h�%%^�e������]�y2��wH9K�c_ /��1j���y2��|`�pR�71P��� ����y
� ��;���X���&K΋@��p�"O��)QO�t	�yz�iG>|�LqR"Ob���ɞ(o�ұ��(�$�j "OF��f���t$��Ǔ�F�:�I2"O2�K�f�WR����R�&���!�"O��:Aā�!v�3d�	E�.Ԩ#�'I��'��
���7f�B�1�I��`H�'nH��@^�t��5T
�53��a��'�v��5:H���ş(l4�!�'�8Az��Ț)^�5�2m��T-��s�'�ʝ0%*�}�6����/@O0���'\���c�q�S�M��4�L��'�^�Ɖ�-6= T	��1������?Y
�D�|Ys�Z�W@��q�n^�H���A,�pC#�J?*d�hG�O���ȓl��Bv�4�>�����~@����ް�RQ�P6l��'J�??���ȓ|L��x�&��<�9� �ɀv�x��ȓ:�(`2��ʦ	�.a9�e�>��ȓq�p���)��V��h��޾NIH��ȓĒ0 ��T�B� a�5ϲn���!��}iqiŰm�J�KP�E.��Q��,�p��gV�
�D��2O��;�4��-�:���C���������^��ȓad�X���_�v�kP�`x*��ȓJ$6u���\�$�nHo\���L��'H��q�.#A 2���|�N ��'{�<b��8��y�Wg�80�B�	?+�$�h�#�� ��a
±��C�I�}��I�d�R/bW�������DC�I�0:\35�!rx���
ܾ,i@C��.�q�AaH4�,"ai�1�^B�ɯs`�	(�I�s� ���Nػ~.rB�	�j��@���͐��t�󇙵q�|B�I+MX CG���,Hr!�p�U>B�I-��r+��P/�x4	�:��B�	-+8��𢎐D����>)P�B�I��!��%|r�
��B�f�RC�6`��hS`	�$U�� ӪG=�C�Y�h����
�u�bD;p�ۃa�&B�=yf�@rrƞ�gBjLc����JC�0l�a�&9?NdJUI�/) �C�	�A��X��FI�
r��xR��M�C����س�(E_3l���ܱr��C䉂 �X��7/P��� A��C�I4Q���fe�y�&���C�Z�C�	�Y1RA�7c�+pMX�w�ܗA�@C䉰F��EY`@��4Y��nЩ[��C�I�3֧?̶=p�
OxX�C�	�.�h;E�z���H�ΰ��C�	-yj�(GΓa�\s�96ؠC�I0&� X��  ��K���w��B�I�d��BF�ȸV�0�M5(	�B䉵!��i��K؃ ��Ti�h�c֦B��1[��d���&Ln<[t�Z��B���zi����p��e�'%�d3VB�I��NQ�cW�-g�-q%ġ+��B�I9kŒe!
1*¥YQ��N]�C�	�0�Vq�"�Z���\ ��3=v�C�I�B�,�*!��$��K�W�B�I�&(�4[��G"��଀8n�ȒO��=�}���2��ǌH�f��0��HV�<!��M�O5�<P��)�4�ub�O�<���1;x^P��f$�<�!`��K�<� X���a�4e���vG�,gČ�"OJ9����w��<��GM�\6V�i�"O>����R���i��ۮ|I1�g"O�%���$�:��6�̋;4���_��G{����Z����iF �����f�!�$ܦ@�v=Bum1>ɮ4hݽ<!��� Hz= ��V�TP�!��*�!�N6z�}�iG�^���u�O/)!�d]"O�I�Ѩ�s� ��/ԋ!���SX� �F/
���U�!��Y� hip'�����H ��'�ў�>�3�E�"$
���-Xd���5�?D�\'MS� ��'K�G���G�2D��S!/t�1" �n���E�;D�TR��?U"�y��^�#M$�I�N4D�����P�V�X�o�I��kq�$D� ����4G<i��J�
XSZ����,D�l8�AY�d=pay���5i������*D�H���ܒP倩�"i	��P��N=D� a!�/2d<�Y�ܼl���J�6D�D����%@���+�hL���(D�t"� H�L��&ưW�Z��w%D�(ð�:w��y��O}>!�#"D�X�H,v�"�2o��5e��6�-D���ħD./߮�B6�Q�&�ٷH,D���1"ޑn|�+ Đk��[�+-|O$�D2?�b�"8�|7$�Kεч
O�<a��=h��*�MռZ&^�!�$�M�<a�F��x{�h"c�:E!�g�D�<�E(?��i��H m���a4bY�<)��,Ly���
}
�d��T�<٣'�b�P�r�BYKF�"��_Q�<q��I��J�jZ�7Ϣ�"�I�O�')�Od�)��\�\�@|S��E�0����ȓr�j��/��G���jU�&x� �ȓb
�����[i���Bv'N�Q5,��<?>� �4p	�Թ�'�t�5��u��=@��ڦk2x% R�V�8)����`2�A���EvX�cU���\��v\t���HfN���M"AZ�'���Id��DUg����]�w�U=��a�5D���E��cYB�Q�+�M]�Iq+2D����)y85b��ԔW�֤��5D�H��EB�W78URD�l�b����4D�@;�,ԝfblQ˱� c,@�rA8D��*��V<��K#�ޘO�n�0 �<����
fT���ա�R�ҙ�Cغ[�<�=)Óa!8E�i�/� {�#��D��w��A`)b�"c��R����ȓ2�Xly��#�r��������y�BT�1I^�G�,��1�ֽː��ȓ{U@�W�EZ$u��F�h��!A�����R�;��4M.�F{���<��3XG�tq`��0{���3�^�<كG�i	Tݒ��U�:@m(�CW�<�G/����a��,ew�H&l�O�<A��įo��Z�����ț�A�<A�xK�@��C:�P�3��r�<q#BY�1�C7�ۄl3��"Gl�<������t<��O�>\�q�l쟠G{��ɞ	~�h����B\���E�F���C䉟I{^%���T�*����oD�k����0?�p`��itT��m
.fQ��h�<`"\+~�p�) o§LYJ�g�<� PM#��5�؀!�O���8G"O|��*	i����%%B��Xg"O�9�ת�C�pը�*�+><br"O�˓�ǅ4�F 3��yq��{'"O�|(��
0z�<D���Ӕ']l���"Or
�+���z��ǋ��W�<�""O����	�\jD%_�@D�p"OHrt.\2_J|�ˑ�py��4"O�Hyq�Z�*<���#��L~�#g"O& ���	Z� Ѩ$h -�R"O�<[���P�FP����H��1��"O�yQtbA�C��`���=[�Z2"Oe!îӊy20����̱<PBRS"O��+�ur\�ZCMK�a�U[�"O2���Ef�٢�J�`qQt"O�X��
-=d�%zw*�)&�xQ1�"O<ا&B�VP�Ǣޕ#�:�{p"O� �b-�<�$�r����:%"OdE��BV3Kh�h��a	������"OĀK4(U��@��&E�W��x��"O�y�Q��/kUD�	��G�#�4��"Ov�eFj�<���ގK�$| b"O�E�b�X�i�:r�i�{P��"O�9���R,WVl b�B]4^a��Ie"O\,rGQ�(�f�xᄖ8]�a"O�f�1J� ���Bi�F铷#�<��nnD0&NО,�DЧJ���|Ş<ó������a�-��ԅ�'}t!@�)�����gP){H}��V)��S��5P�+u�6 �`�ȓ�؉�g��zT`S""T)F�(��p�B���H�6
��*�bG)M]ƹ�ȓPSd
e�1^|��NĥVN �����!g��.�D�9D����8p�ȓw����M�"z�h`�P�]�!���NI�lSqA�8��If�в4!�D�����[�I6AVV��E�ӳ�!��1Z�*e��g���1�9�!��qÜ�ۢ!/�\����Y!�d�A�L�R@/Q�.%��	�m�!��V��:�"��w�lв��;�!���r�����ϴ�,�c��Z,�!�d!⺰;�L ���T	�M�!�DN*؜H�e�6>�@ȚVl��]I!�$G.$(@)v��79�Jy�#�BPQ�2�)�dk�B���#��W9O���C"B]!�y2����ɐ�Ј���Xt��{Ј��SH�UT��cf�愇ȓN�������M�X�d��0��D��P�H�Q2�	�u)���g�����8h>�aCM �p��ӡ[�$4��u.A����tw��(���7��?ɉ��~�ч�Kq,��$��4Ct�jՁ�D�< ��=:@i��+�0b���g�<� �]��2l"��_��P��u�g�<y�b܄K �P'�?O�1���b�<��"G�7]:i��:r|��J��QT�<	ã�9��T§B��Rx�����V�<I$/� v5�X�^�1��y��NQV�����n~�  Ӝ!V��'`��,�q͛��y����Tb@$���Đh��� ����y�bŨN���LȨ[�n0I��M�yb��VN ����҈E:�y�m���������"m�t�٥�y
� bȻ5!O��hԋ�g��E��|�F"ON�K��K�2�yr�Ha=08�e�F�����J~"��FҢp@�M�>�L� 
���yʛ ��1�°I��b��y��m�@-��.M6Hlԡ7Ő�y���t�ƀR�%�%=\�ؑ�W��yb�%�-R��Ҕ4Ѿ!�ai�=�y�AY;vI��S�cW���1���y¦�7	���#c�(<@`�/�y�͇^���
"���_��p�gL��yr(y�F��0h(�� @�б�y�����0�+Q����n��yRJ��yf�`�����H�� )6"ƺ�y��kۆ�Rq�į>(�pJE"��y�!�*K�l��./��tp�ŧ�y2DL s���Q(�<��݃����y��D�Wm�QI��`��M0@�N��yRM��;�(�3%_�S<�����I?�y©�.$��B��M>�:A�1�y"m@�n^D��K?3����k��yr�R M���Af@	�U��X�Cͅ��y2.ӊuΈ0D�I�EF&	肤α�y"��/I�t���U�1��ZK�+�yr��$�Dm�)"�� Ӧ�؊?!�D%�e�� ��5z�P$ 
w�!��:WC��95a����b����!���EPh��Ӫ?�l �BH_+b�!�$_��4�Ⲋ�1��|�'ȣ)v!�d�)%��ջ�(�z��"��#Ov!���
��R�Ԇv� ��C�X�^S!�$C"h�x��ԦD�2�(�2��� !��J�q�th�F$�c�<�4
M�L!�Dҟ~AZm�L��
"V0��ȟ5b !�d��h�e����)Q�hH�ö7�!�ĕU˄䒤�ΦJ'|����In!��]�Io�X J�V�j�F1g!��U-D���
�9A&�+EPȹ�"O���C�Z a0��A��#|;�.���"�O�5���Шj�z���DW�Z�J�s"OL�r�Ӌ5�Ή�2Õ#}���@a"O蹲兙�ok:�R%dH,IX՛�"OV\�i��8[x���m˫26��J�"O|r�h^.PM���K��e��E1�"O�T���!�|����͢#ll �`"O�X�!�� ���K'�@�4�X�i�"OJ��L� _�6�����3j9��)""O6��Ũ�.m�R\x�kG�*�0"O�d�G�����C"%N�cr"O´*2j��IQ��Ӗ*g*�J�"O�S뛈.% *Sp`s�"O�)궉�m�l�T��+YN��{�"O�#��P�H�H%
7H^5��Y0"O>i�F@�b�����@�*r=`p"O���q�X�Ty��R̶6�8���"OZ�hƤ����Ƀ+��yZy�w"O
����["�C�ަ.u"��"O���e%`�I#�F�q�#d"O������v��QVF! Y��[W"O<D��R���B%��<Gj4��"O�
g�v���qoG�4aH���"O�M�u�G_W�\��+I�Z�d\��"O��4o�;R�e�jJ��(�"OB43�b^&�X�
�fF�j�±b�"O�Y(ՊW�j�Hb���R�~�2a"O� ��c�ď�(��W�LĀ�"O�lk$�^T4`B]���l`�"O0��ހL:B �V�e~�k�"O�x
���^F���5�ާ>� 9Ar"OX���R�B��"U�@�X#hiH "O���q�_�5u���gcWs� x�"O��x"��X�9p�":R���""OF�9g�'�@kUŢE�\rgO�m
�U�q����N[�� �	9�!�$8��(c%1x!���i��u�!�D�c�L9C�Lb~�XXqIA)2!�D�U���gE�.Ey�,`r��-C!�Ę�v沘�l��?b��i6j�$.�!�$�$�fxR$�V+-�<��0��/U�!�D�5T���*���	���L����
=,�^����.Z�H�9��E�lE~C��2 	(����7�PP�PJ�7�hC�I��R�Y&-TWhѱ�O �O8C�IN��93�ߎe�6db]g'"C�IΠ|����a&,��Hk�B��81��}"`�K�b��l�g
"
A C�I�sIPhʠl����v�4B�Ƀ\��DБ�F*�Rl�'(D	Q�B�9g��=��T#VU:��%�C䉟s����� 6+P��^Q���	�'�Da�t
Ÿ8~�t�%M��Gv�`
�'&0����+(P4��Q&T�P�'��Q�Dj�-%���J��ũ#f�T��'���@�bQ*l��-֓RA
���'��A�TNJ14 ����@V��-
�'ӆ�餦L�wL��Q��*Lk�U�	�'��u�W�S�:�Kq���IuT �'��(��tf�BKΞ<5f�(�'LȅHDE�.L������7]��B�'�����E�h�p2�1$"�	�'È塑���� �v�$\+�'3�C&(ď ͠�8��B�!$X��'a^43����u�����W ���p�'n���!���M��oT?��'k8�2�� ���X�+� �ɩ�'��|�ѫ�%�dH���	<aJ�y�'3��p������!v�@�D"���'���u��>A�}R�#�%�h�<i�_8���Aƌ�1nҒX�FLN^�<�b�JJpz��TI�91�)�X�<�%*�mR~�XW�B�x3r�(��NT�<1&���
<�v"$eĚ���n\M�<Y �T�<1��ag�["9�8b���E�<���� ���:jX���JI�<)ABnt&zp�� �%�o�<!�G��1"�L{��LS�N�tʐj�<a��5\�$h'D���Л�%c�<�u9�z��R��= ���y���[�<A���$'b����P�x>B`9�Yl�<����<c R@S��-B���@��I]�<����n��<���Z�=!����S@�<�p�σ ���1��+����\{�<�$f[�b��,A�#λ;�*��v$Ax~re���0>Y�K��`�����4�^,�P�Z�<�S���.x���ڂ�h� K
V�<a^ɠ� �-*�p`8�gUR�&=�ȓb0��ReKߊ5H��A �$��ȓX�d&b�%n���1��A��$��Vs��;CJ�}���e!6r��S�? DT����D�v�� Qv	($�|�'�֥Ǎ[<��;hR.���9�'��0dg��r�
�Bч�9d�x��'�r�&�ݒNr��b�L5E�q�'��ۡ �8x�F=!0�n�j	�'�v�C�\GW�H�ܳ��
�'�$�;����%�J�+��,��E�	�'�l�W ��	�ō
՘}�	�'�>A�ɏ$8��m�  )�|��'4 -���^�?�V9[�G�3��<��'��h��X'�`[1�_�G�N ��'��ih �Ą-����@ �@�����'�^m@Xh	G��)Sd1Ӄ��y��&>n��SgDF���eFP��y2�*e��&O��Be�X�����y�C�$2xa�"P(;���w"0�y��i�<e��<7�9��+��y¤O<b��$�3�؎?hcg�֦�yr�� �.1��Gl��h)��y YH{�D �-�J�t��yR��o�,=3Qj��4EV�j ��yrb��
�($(��Y�&���y� ���yb���xID3��E	Rm��y� 8] �Y����2�4���́!�y�i��X����)���
��yBA�z�T�*(8����F�Z:�y�Î�,�h��߭-n~�`�*	��y��>gv�2�������6�y�,jA����!H�hѭ�y2`A:!�jꆦJ9r pS�J�yb"�s�8�E�U9����RLH��yg�	�	KW	J88r���y�E�Dv�P#�}�.�x�bK��y�j�&4�fi�U��3y��r�m���y�Y��QRĎth<q
s���y"�؊ -�pk�,C�oe��QŮ+�y҇C8_|,paǭ�np�����y�M&D�0��DkB���R"�ybG�x�X���^�e�D(���y�*Y7*
���� {��B!���y2&חK�HL�֯h-l|�kQ��yB�04�Uɋ�c�@h�'ſ�y�g�7r���E+?Y����邬�y2��%]�-�Ɖ��x�D�S��y�	�=	�v�^�jp�
�S��yH���U�	&�<L�f���yB&�d���c�gB%y���y�̎O�b�����mJM�V+[��yr���M�*(h��H�8{ ����K4�y�L	#�����>-4�r���yrn��o~���N��y����f��yBȃ�H5 � �PrԨź���yr�ٹ!2Ȱ��_�e�B�v���y2�	<�6�C�@
�
��)+V�ė�y��(_�r��6d�����s`�N8�y��]A)x�*2ɐ��ǅ�y� ��+Ȃ���΂vl�d��'�y��G�3�uB��2_�����(�y#���aң��-;�t1��+�yr$�Z^}�G��P��\)P��y�mB�4���ؑ{N�P�C��y"GզW�X5�3�ìb�dLpN���y�H��@>��v��]d6�7�W�yB!��|V�u0%�\�9����y
� 6urH�p��8cg*ߘ�H�A"O����LѓM��a��3O��I�"Oh�kQNص/؈p4%�]>F�A@"O<qS'�ԭ%���:U�͂!=l� "O��)"��N�	��u�H�""Ox�YM�2U����W��2�a`"O��ȟtt (
S� ;�:yZ�"O���v��Y��1����u�L��7"O��Z�$|ԙ�o��~#�]+w"Oy*�(�2�L���c��~,��"O6�����.�ؑ���	���1�"Od�ِ�/w��)cb�J77�~��"O��(�A�(+�� BŮ��6tr�"O\u�u�Y)^�R� 3.ɮ~ָ
"ON���!B�b����wLX�=�M2D��� �A���B�V 4Z He##D�Pi��t2����g 6�R�/#D�l�5��8zR���AI-D^��"#D���5�3D���YwaF�`�B|`�&D�h�Dֽd�"	S���rB�� E�'D������&T�8�#��7p֬�6�!D�|Y�%�8��X�c�vqtY�1�$D��+�$�H�^`GX!L������?D�@R�gO�Ͱ�BJ6?��eQ��>D���ckk�Fׇ�pn�@CO��yR��v%�e�R��@��4J�o�yrIQ�j5��(�ȋ��8������y򅛨c$M�u��z�x� ���y��<y��F�V���f&%�y�Ϥ�I�(���!�!��y"����`ǧ �"��߀-?!�DV�MX|H�%A�9Ft��d,�=:/!�DO,
1�Y!�F�OG��23��"!�ǁ"��ኴP��KBbA!�D�'b{L}��X#`��ݢ�˙�Xa����b���J������Blߵ�y�������̴X��U�Ⱦ�y��L���,��%@37�3�I��y�%K8.ɑ��&-�P��埞�y2�(}q�C)�Q��X��y��T�6�D���eܙ"�(��FN��y�m�F �m��a^���%�Љ�y���Lڑ9�
��4.N$1����y��P? ������\�E�wN�y��.���[��ǲ���q��3�y�c�[P�E�Q��y���4���y�Xo.p��%F?�ࡹ�E 
�yҏW�}���Pd��l��%*�M@�y��D�=8�� �ߐ_?�PC�٣�y��ѐ}@���o�7n�"]3����y¨]�uj��Ύ�=mnihݵ�y��E�J���I��Y�:آ(��A��yRL�Q�Ӎ��>a� ����y2EԺ�,T�V�� {D #�_5�y�MI�A��R�kWL鱣���yB� (�Ĉ�닂3��}h�&�yoD	8$qB� L,��aa�� �y�bʂ:H$�+�c����ph��y"�>;����Pꅦb.�	G,�5�y"�Ix����6�M�q�F�N��yR$Y*����1�S�F
y:��/�y��9���qō&l�(=�%���y�aTt�+R��f�JXFcQ>�y�n\:_���2/�\wH-9tNÀ�y
� B�A����,��A���L�v4@pv"O0�8%4-$~̂��<<���"O����M�-߰�Y�7S:��"O���V�6CF��i�m�4�I�"O�����[5LƐ�Wcʔ@)I��"O��� �H!|��Tb���a��"Opq[5H�2c_��q����SΙQ"O�哧(��Q�|���@\�=PF\0v"Oj}I�
T�v��٣!fJ2-�AB"O��A�ה�n�C��U��`�"OPq�ʙ�L�)sd�(&{ U��"Od��0�,mJ��[�b�:���#�"O�uh��7F��S�/W<�r�X�"O �)����;���w�>�Tyic"O���E^? ��Y�.�g|z3�"OV%@A�T.!�����1~cN8��"O�)P����<�WO/V&��E"O`! �bP�2�iFC4ZC�{�"Ob�ÖfY�/�$p�@���>�`��"Or5x�K��t�=��K�BU��sT"O>���iK9�.yYa�������"O5�fK�\���T�T?>�V��%"O <��,Z!@�Dx���V=4��}��"O"A�Q�AzJE�� N�R�Ę��"Ox1��]�;�|�������4�� "O��I��g��x��ݰ_��=�"O����;]�AH�#ތ|5�"O�i����%\�̩C c� �
"O�H5I��
d$Ԉ�h�E�"O*�aa�^�����ao�?�l�"O��* S�X�p$��x�"O���a�J�$�.%�jL0�`)�0"O�!؂@1Z�`(�D��r���� "O�q����!��)�'�^���"O��3�P�H�r���HK����"O��
tʀ)Hh�b����4�d�z#"O���`?,�A�"��n;�9q�"O��Kf�9��Y�&�Hd��"O4@*3��@f�(8rf�9$<1�"Oʨ��"�A�fhɖO-:&(��"O�����/K]�qc���6�1��"O-2dܵd|�5�îF���A"O�Y�"����qbb�H��- #"O 4؂hL�s�µ{$���qt|�"O<���cOa'4��10T�ia�"O��у��|���g��t;9�"O�H��_ %�ph(�eL�&/����"O`PQ�]�+t,�H@�L11ɼ$C�"O�@��30��*a�EL��z0"O���e����hȉ�d�-����"O�`�K+ H ǄR+08����"O�u"���W��p���?5�MBb"O��z��8Id@��p�_�h����"O�dC�N�%k܎p�S&͡*d<���"On�˞�a2���o߬((�)�"Ox#s% }�� 	��N+e4�hr�"O(;��
#.R�Q
<N�`��"O*�"`��G~l�!�����P�"O��b��+�𸻴j_4�ؼ�"O@@�����L�+���84M��v"O�m�#ц[ʑ����&����T"O���Pa��`{�M�����('"O<<CR�Oto���bB�'����"O���I�F~�A�&� :'[����"O� >�C®w��h ��/,Cƌ# "O�k�f@�k9����F c$4!��"O(�I�C�I-b,S�O=$�H�"O�rD�a��U��q��i2"O^������L�9��'��� @"OZ�����mr���T�x��I�"O!�eL++��<���f�abr"O@!A��I�+���"^,�:QR"Ol�sEN8z(�ș�.��C"O��@�Z  ���z��8J�R�"O:}�5��59�`�ő�P5Q�"Oԉ9����Y,��D�*jp�	"O��X���=�(Myu�R�Z�6�yB"O`: �@���\D-�Q�*<�"O�T,�,Rp��߈K�v,h�"O��ӭ�0L��jʨF���V"O\A�RZ����,�&��lҔ"O��*H�:`��!G�~�J�bu"O�E�W�F�W���7�y�"O8=�"lݨ` ǭZ�^��8��"O�}�bfJ�y׺�HmG�h�t�؆"O�$Ja\�P̜�)qO�>����"O��[b��t~�Q�ɓ3k�����"Oȡ�nӃt��YU	ƪA}��*�"O��ǒ4�u�P�Ґ5�b�""O t�Vŀ4J������U} �Ҁ"O�a;�`U1T��q�BT(|��4"OnQ��N��Z��'�D�E]()�g"O��AW?!��/����	�'JZA��D��U�g�X�kL����'0� ��AIf���Jg�]��'��$���_6^t"0�b�O1gt��'���2AǕT�a�g̯2����'�>XZcZ�Z �J�	��i��'�ڑZ0֝q��4���F 00�D��'��x:U�~ՠ`G�QE�Y	�' ���cǾt}Ҡ�W�8����'x���_�A���r�H�d�j
�'��; `�?>����a�HWvL 
�'/�h�F�Y�5!n$kae�Dx�)�'jt���$�%e��Aa�Z98K2 z�'����+�DٷK�1m�1@�'"Z�ږ��$r���G��=,҄b�'���)�dtÃ�b�ذ���:D���C��5�U D�هM�h�7D���F�2Ű�� 7���H �3D��q&d�3m���b���IȐ��0D����d�$�@�#7e��(c\9٦�-D�L3�җ;�#�ɋ�>%�*D��b,>��I[g.�{d�`rpc5D�Py�˙s�fU��哢)k����@7D���2J��J���MB��i�m4D��C4��J �]ذ�(O�ܐ34�4D� �"�!T^��� ܠe%0D���pcH	2��m�$+�5׋.D�D�FK�2H�P����$]��F*D��ڦa�����׏3�xu��%D���p!N�^�L�A2-�p�d'(D��80�ܐs�tP3�@S�S`�4�%D������
��Qz aV�roj,�FD.D�P�sʈ,[ru#�/U�w�x�Q!,D�j��
�I�8ȩ��:d�/D�;�-P��p�ʄO![�1:�l1D��f�O
>��ICѦҨZ^t�9 i0D�� T��gOI5��
���J���"O68@WY�;G�-���I9�va�"O2��$(�x�V�ҦhD�JP�=0C"O�<`�ټE�Z�*���O��`yU"O�j-Yrx$��dL�E��ݻ1"O��!��y-3U%KA�N���"OLM�fɏ �x5���e. �r"O���:!�Y�F w&P8#"OP�Y��X�S�]�O�!c�P�"OV�k�b�x8ғ�ٙM�es�"O�\ӑ�\f��9��L�'I���u"O�qp�0@� ��%M�V	H�	e"Ox���u�\���Ƒ#��"O��3���'��IVňM&:#�"O�\���A�{� ��B�"i �"O��	��B#?*n��P
X7 R�c"O�t3!M�.�����e^���"O
՚w�� FD�e�ܖ�:5ҧ"O�@ӑN��4b
XBRKC'��(�R"OB��a��lhD4bᚄN�v���"Olz�`˷s�z�[E�]|��2�"O<5���?���	�9]�ӥ"O"|�dl�!+}��za�C�!�����"O��K�eҥ)d���Lc�"Y�u"O m���ޑ �6�{ׅZ+r�0��"O�`8#�  ��9��L�&Ҷ�"O~��J�6�"T�#�P���Y�"O�YG��
^�����E�lU "OT���gղ6{r0��b���¸��"O�]�S�+
Xd��KC$x����"Of�HU��:^����G�M[rq�"O� ��u��@��L�	���D"Oxe�#k�2},4@Ѝ��f+��J@"OP���jН2�����B+
�`"O�0b��Iz�؊�;�e��"O^(��$æ!�g�Q/]���g"O�<XUf�0Y`D�p� R�4)�r"O��qE�#��Lٲ����R"O�9y��N6>E����(@+u���
�"O�]�Ԃ�TU�$:�}��(�t�3D�����M���Y'i8�xY�`2D�8Xd�2��]��Y)?�~�3�4D���'n��i:pI�K="�b��$D���jA�!L�	%�R.O"��2i$D�tˀ�Q�*-�R������ D��HA���%ې��%U('!v�{4�>D�`��hM�lS���z'dmr'H"D�X����~5t�q'�
�*a{�'6D���0͔h�T(@f��n���'D�|�qf�13�\�#��'� i��9D�4�Boӥ,<�t�O<�P���7D����7WVvmQ���,S�X!Qp 5D���-K@`�&�'LZ0���g2D��rl��-o\���@J�3-���.D�L��ٽM~`PÆMI?��H�
-D��y��AP�B�Ѵ��x��(�3� D�$V�* �L˷�E�W���d+D�,�q�@��5��,z���*OZٚ�ꗬI�$i�F��=���Y�"O��A�i	��2�*Ҥb@���"Oj��Pd΋c���,&���'f�\��oY�p�♑��G�*`)c	�'���h�2ZV�h����6lh�j	�'�bUb�ֺ�2���LJ�|ʬd���� @(*A��
���I��ބ[ٖmC"O��)��ʥ}�0����C�Ԉ��"O�)�VG�4IJy���vҾ<�S"O� @�)e�J���#[�E`��K!"O�XʧBP�.y����I^�rs|!!�"O��( �p��5�4OS'©�"O������*~H��'X�쀀�S"O�������S�F	����(}f%��"OZ8��ª���jg�G5=�|���"O1"TG�n���yF+��^�PA��"Ov�1����
Ba� 7\�Z�"O�\��Wn�<��E
�z<��E"O����H�Vs���Y�1�hf"O~p�e�]+_w�h��唟|)�E��"O�dBU;�-;'��>?ò���"O~�W���6��L�@�R�5"O$x;�m�;}N��kX�pR���"O�i��ۥm%�؃���-GKJU�q"O�i�r�ߒ1V$\ g�{,�Q�	�'��')Ԣh� ���X��ح�	�'�8��Ꟊg�dс2�V�_
F)q	�'3.5�H�7[�������U�<��'�ƹSpR�M�n����2S1`!��'$U"w��?@��A޼M3Ե��'��i�#&_-Z@��Ȑ,E��0	�'}�D�AD���d�P�X�tez��'
t�*��57`��`�]�e8�')�L
Ѩ�*_�`�7)��
����'~�Ac��*B������7�����'��l*�g�7E� `�7@ /:D��'�@̉�Ǎ�Q.�Ap-��v����'w���FD��\r�`10�ۄi��I�'�^`3��Vצh��/Z{B�2�'F���O`R��g�U�����'*�sa ���lX*��"dx��'0���F	�s���	�_� R�B�'ɖip���b���@�B�
���'���A�ԱMpbmJ�&�	@"5��' �Aq& D=�F��ѳ7�J5�	�'�� 閏]�]Y��"�Q.�&�{�'�0�/���2�@=R���A�'-*���X��L�y¢��
�'�Fmi�X.q }3v�U�j�dP�
�'ξ r J�<�ځY�7t��*
�'�X(A1 ш)&�C��:��4�'��l9�m �"%>-)�mЏe2��'\8�Xq�#%9�Bc�<s�'ꎘ�'݄/D�9!��X�P�0�'�B�c2 ��W��@�N�B��h�',�A���2 ����#PKX�x�'o��J� {:I
"mV"E�B�	�'�d�c� Ea�(����5���1
�'�
�O�ii ��b葤,"�x�
�'���%�Z�L��c�!��	�'����;lnyHb��(yL}��'`rX����ʸ����.�Ԛ�'Y�8j�0A����']޲�j�'����Ǽ0���'O�d�
�'ټU[��\�G�$E�?���3
�'�N�x�MO	A
�`r���IRZ�Q
�'��lX�I?T�n���1����'��鋴���Fl�\)�c��n� �'xFm*�b֨^���C�H�4Td��'^x��@�+
!�DR�h�x�
��� (�6�C7~�4j��N�`�q4"Opd���h�|(*bcZ�t��#6"Of����c�|! "̑�.���"OU�6���8f��@�\=�\��"O���RGISn2|{嫋�&��T9�"OhL[�*��%��A��i�7k|��Q"O�UJ��o��鑪��7�V�C"O�M�VFF?g���3H��%+V��F"O�9֥�8(�����	�%��Q"ORT���<k<"PAa0��h�C"O>`q�g�K�����@��G�<e"O�iDf�&+���1�NȶL���X�"O6m��c�����d�:
�� #g"O�9�`kD	,ۂ�(����QUt��"O�b�P)(��a�1-F�VD(9I�"O&|qpd�6*r�(��757�!��"O,;6$�5_��6��"&긛G"O�UѴDΘ,�"�9g,��5
�Xч"O�<�4��>/���&����L0�"O��a�ꕷХK�@�<-�����"OT �e�.޼�#���'p�}�"Oα!�j��/�a��EI4V^���"Oi9�Iڞ� EQC�S)&}D�'���I�H�嘧��>�0G��G�bP��y`�|��h*D��`Z-�P�z��[:$̲��5ˤ>���
��-y��'A��,�!<�6��%k�,�F5"� �<�*�HܑD*��H7J��b��dPP#Ҡ5M"���"�Oh<�U�*N�:��(�"8=bt����]�'���#KȲW�m*5�1��F�T-A孂�q���ҧ`��bu�B�I%:b�X@#�!�5���P�:�X�C���P8��Z�mQY��,�g?��̤z)JH:ǁ�Hb��u� \�<��BQ9FWl��
���\�7��ݟ�{$%ւ/����} h��D�1�4k�fL=_����t�N�y�F�=^������
�H\5� �[�H"�| �C��$r΅��D

�Ś�'�v���S�N?xE�C#Mܲt�L<���F�,�}і)�\�BL��)���O�ơ�uK�x�V!��A�?�U��' :`�e�(�H�Pǭ��"�l�j``�'[-"��A�Ռv�v}�����O���'����&T�{���"f �@jԌS�'��Ď۝qu I����V�6IgΪw��!'�R�mq�M�
�wp褆��2id�Z� ���!��a[Xz�?�s�]��HX� �mov]�a,[�;�c��w�
U�%�<iSl5J��x(<Q��^}J\;��-.�՘ �yb�Џg��l��C�w�B��#���P���P5�q3�� U���pc���y"���.1 �8��НqL��i7nՑf��<�£tb�1�d	r�N)N~
��[�$0z�Ĭ���ZL�^��c�54Qa�FJ!c��y2�.��E��i@�AZ5x8�
�mK�%�"DoX��q	g��r��x�j��9i"\����
I�}��A���O���|w$��g�{.�r
�"::�m9��N@.��b�&�t��c\V(<���@��[�h�;_n����{?�%�By����7a��ɫb�\��K�韓^n��;�E��F~�P����!�Np&H��s&�U��#l�G��y�b�:h��#@Ś	5��h	��~��`
4h�e��18��d��pe�H4m�,��	1I}�����������ؗt�0��A�:�R���\-��I��g��g9��ǓN�0��u�	3 P�i5��Ul��E}r�]�{��\�V��} u��K� �(�/R�~��a�4��?	/h�4�`� C�	�H��Y�Ǌ�mҔ�{��L�H����?T�L�fl�(Kh�iz��Y��[%�I��OAb�Ҫ�i��5�<� i
�'$T����Ȳ��1�0-"~����;jy�0��H]2׶	�G�ˍ��S�g�e'�,��(�^ћ3g��Ih�0�O��	��O!$p��� �*"IdI�EC�qz�x���ʪ	���5CY>��'�)G��� �R5�Ѥj�X�b���9��u)V+j�*EK��*����eG�U�n�KQoD%s(���e�a�<��M7���[ �ǧ�ȃR�Py��!�^B@�
 1CxMy��M��(���6'�>w�z]�WBO��("O� R���#$Jh�
�(�~�� f�ŁK��Ɋ{���IAL2�3�I.s\��c�)C5)V��� X3[�~C�ɹ.�d49���#Lu�q����#�H��	ƓBJ9��Z>���L80p�`�$D��.�Z��ȓh���pr*�	}��)��6l�%�ȓ@z���hSos2��&a�f\��&"�|���_+o?@ ���
����ȓ2Rz'���T�L��
�� u(��ȓ/h�YV�c�Dp���SNh�ȓC�<�i�J�N�� e�
;]0�ȓQR��� YqR����U
�n���`��-c$��j���ځI�$�ȓ<�)��GInހM:p-E�Q�ޅ��M<�0��J W��	jdbYH�L���KqD<y�+	�'V���5��v{楇ȓr!4��dB-���GC@�����8��&ɤ91�!�e`B�&E�I�ȓh>��PN�9�ht���z!B5�ȓ.'<�cJ�2��5!7k�9��!��O$������]��<���O�A�,Y��	%R�Vǉ�g^��3bJ�	�a�ȓ^N�UJg��[�d����('jT�ȓ � =��bE [#:X �o�?>��d�ȓe,~D0���&~�@��f@�K����:-� �,�g�}�P$'> ��Ge��BROSF�\�p�S<3\\��}�s�5E���S��'�E��j̬���1Rz��s`X����AA쌉!���>�ȤcJ��)ޅ�ȓJ�����N
�2B:����%��ȓ{nlM�b�� %���*���8`9t�ȓ9۴u�E��$�����9,����"�'���!琴q���2~޸M�ȓTl���VJ�"G����'nI|�f5��|�P��a��w��ԋ�,]Bn����?�L��	��
gL�^�P�
�� D�|H�i^� Və�}�@��w�?D�����[����xEO@�y*�!�vO'D�x0��W9$�t�!F)��Z��!#�/%D�l(GjXR��0Xi�-��-j�a#D���2���D3VM�n��I�&d4D�����R�0L攡��*3�i�*2D�La�mJ��{eg��xָ�9��.D��jդE�������'=���.-D�dȥ��VD��u.��R���N>D���G�3<��xp��E-?䖸i��?D��c�aݷ]��R,��(��5��*O�(#���:TӶ��@ ��_�P3E"OȠ��Ҥv���r��I&��h�"OV�K1�56J���E�� �"Od��s���Q���ԋH�u�-��"O�<�-\!Prz|X�
Ƙym���"Or�H�B���L���D�4��0��"O���`�)������3�<�2s"O���F�5�*���8L� �0"O��Ѝ�l� �e��$ ���"�"O��Ӥ�]�.-*�+
|m��i�"O�1�s��q�t�آI��^m��`�"O���Z .π��P�Ո%�$A["O ��6
IjwN +�S�`�dA"O�^
���% �c�	�&!�y⣝�a-:��a+���,<ju�B��y���-@t���+R�b@J4�D�y���v�\�����0I� $��
��I�" ��*,O� �@�dN�-<n�E1sƇ��~�`6�'<�Ų2�R9W����M�XuY�O�>#h�I\<���%z�p衧O�M���[Z�'i(�v	�%^r��sA�v�� X*�Q�c��R���$�}s�B�I^l0sF�0A�" �>^W�7��g͠)(vH�[hM����}��M��,K	��u��'Z�~\cA�Rx�<��X�$�l��IW�>�
��Z�҈��M�~m�3M��rG����HOJ� �;��˰̓d���pS�'_�Ւb�4C��H��I����0��jX��)ɯp���I@�NL���Z��t����L�c���C'% �uQ
�jc�P�q���Cq�a���=�hM`�c�Zl$��wC˭��L�ȓ5� ����+�����CٶQ���RqK�{��b0�>	4�q+UJ�-�h����:��%/�4-�ZɗL\# �!�dA�M�<:VEĿ`G�Q�b�P}��t`�aPH�C�D�,�VxCU7�Ԣ=��[zYkcɂ�0ĉ��^��ǁ�=��<�6K��r��Q�r/�l�� "��F�xp��4.��M���a.6)9�
��k�@y��[�53n"<A��,�H@2���!W���JK7��6�`@�&���
O%!�Ĉ>q1�eA5�NB�k"j�����3GC[Q��`���#������(��s �� D�r��F��?����c��t�<��ꂑɨ�CP�ġ���S��.]�&���9�\4r�L��0���'�hO$�y�$�+`�N�i��-b����V�'�lˤ��7^��B�[:/j��0��
R<�ST������[
��}+)s
(h��L��kѳ�(O1�P��(w 8��ѻ D�˟�c�:6,
"P�0x�MG"O���3H�7�^dI��37��I��	�>�,DJ��D� �:,C�Y�>Q?�$�0|T B�.4Ρ�Ȝ�|!���B���F��$1T�G�X�R��rhD����#dL=St_?#=���x�4�3�4�`��gqX���	ϯ`^
��7�T#Q\X	�d�z�:�Aц�(QF�("��U����`^jT�h�N
'�>H�7k'��(���fܠC��)��
4P��1�)D��J�t!� }��)���) �ti��ID�]��ΡNH �K��)�'M0,C�<d�BC�M�:����.��(��	WJt�"�n�3b��t%��*�Nճb�ay2h��T��?2�J�"S��w�!��6<hZ+�<rTLzr��'?�M�ȓ(�8!8�B*W����4��!Q���ȓw�"$��	�����N1艄ȓ)�\� ���/"���y�EO<UF������T`O_�pmAQga�z��ȓ��h3GI|�u9e��>F
��ȓAtJ��3����q�"-�>�ri��hĐ)��ۙ6h�qqC91#D��ȓT}� �����"��?�����8g���?�Q�u��-ȅ�_s� �q2I�Ԫ�'u���A�"��'R�*�F�`奐�������6H�fX������j���J˺"U�]�#�X��E-��'���ȓ ��ћ5l΀$�B!�œ�B(�ȓkS h(�%:LHIF/ϋ%�$�����*S,E̕���	O����|�̬2��B��(�z��E?OLr��XUTq�BHG�w��%�I��f�Ʉ�%8j���i�FH����qG\Ň�IO��2�+�lնuT�W��*���zEtla�i�*;�ꙛ����o׮���!�ʝqS%@�BFf}s��v���Q�Z��'�F-򖝚@�V;h�̇ȓ5�f�i�"L�i#C3d��ȓnR�x��ܠ��!�60U�L���J2����	Jqr���eصHN�H��u��}Kcc�#0�Q�V��
/� ��S�? L�� /��Дpp
Ax��Q�"O��i�nΘE
D���85�52"O��@q�N;�@����G��'"O
$��J�"�d�T�}1"O�0r0��4��)څ*ښ�ر0�"O��C��+����vN�p/�%i�"O�\+�W�	�֬��ښ~�@AB"OMR&�ǁj�P�zB�۱oh�z"On1��%2z�p�{�cܩZ#j�p�"O"apu"ז@�6�+���3 ���"OdX�4�%&\b�(� �s�
�Y�'�y�$�9 &t����.%t�`��'f�}Af+V�z��7�ȅ�t�1�'�{� g��\��	�(&���'��d�A��P4�bd`!�,K�'8�աrc@�^��4�^*�hPx�'��< o��Nv�@���
� "�e��'?d�s׌��:`ī"J�F���'@����א Wx�6�ɬr����'h��l�2 B��D�]�dVĝ��'A�$�@'�<-�T`� �ޡ^�ua	�'�x �%��"|DꐅɜJ!.)J�'�j�['�]
#o�q1�A�ek	�' l�!���E��|��n�A�����'�L�i����p�(�굣��0���x�'@dᅞ:CED	��H�y
��	�'Cx]`��YF�;g�M�4�C��V<�)��E{�S�O�Z���'�� ; �2���!@"ObEQ$;)wةP�'��.	t�R�@��΅�=}2xYӓ&UKG-*��	4f��N�\��I$�0�Be`��E�BD�a(�^��8���t��!�6n$4��臅@� `F���.�;2�As%N1�i��1��� O̜8��I��lAr�f��>0>�`�>b�!�H*�D�`��9ghX�n��0φ��@NE��ڸ�F�y��ʧ	L�dI$x#t%?`ȉ�U7D��ٓ�E>Y^�p"'I0�r���A�O^軕%��"y�(���G�[�x��ЄB�̒�.K���� �+��<��ϖ.J���RB�ڨe�i4� ϒq"�2)b墠g�
l���G~T��N��|��zCÂzh'�<���+ :�VhN	P���
�/�cܧz��ؓ�B�v{��!��0��#6�HID_�:��ғÔ	o�c�AM���CG�)>?N��v/�aܧ��OL��QvD �B�^V�9��~LT"BL�:�F$���,m�e����!����� \6B���k��=���񤌀Et��$��la���Dmџl��Ȓ\J`�m�-N�A�@P�����뉔a�XD�7,[)pAB}i��>��j2��*�J��\�S�4Âè<!��w�X���lʌ&���a�)Q��%�}���0[,e�T�R����HFg�<�@�C�1p�D�Ve�*x�P`p��"pq�'��o^t��g�I�+*�$?��'�)}���)r\��{c�1ra*��t����?�⁒P�&QR D��D�����oޡW}�X�� S�OJ$3��I	��12�G�4�p<�g"�v�� ����h-�9+�x�''�XQ�K�H�b}�&�4�l���L*��E��ȮXk�,C����4�Ro?�,��Y�E�Z�����y�1�bO��(j�B� ��T��l��|�ȣ��S*V�@��e�=	���Y{6FX�Ē�y�i�"��[B�¯cbfQ����X]S�+;"�>�26�WH%�,�I?Q������IY,Lmڶʂ�MV8 W�B�6��䐵Vv�X�ưW�\S@�׻xD��'j�0|/p0/a�H4K:)��#u8O��[Ѫh���7O�\�ȗ�	����ض�P;�~=AQ�	y⼀�JL�Vm�x���?�V񃔍Ǩ&�Hb�'�H����@�be8X��S#h���'�S���k3��z�ԄR-Zٛ�@ް0��>uL�=5��m@G現`:V�	�l#D�|t�ŔB��り��Y�6X2�D�VP��9-��I��	� (&�O]Vŋ��xR��-\Ozl2��o*(-�� ���p?	���D�biCD�4��`R��}Z���lδ`I�$
cA�%�rU��eQkx�� |��ց�X�@1���������60d�tj�S(���휆6:�h� ��}�bGE^�VL(0dh��yRB�L
����샘f�ԡ#'�����g�5�2GV����l�n�Q>u�qk��a��̰�K�D���Zs�.D�t�`�ƃ2�t�7Jɰu�t;�O5j�`8�H�6�^�g̓=��0��16���-_NHx��RM�u�PF��B����Qi��F��"�ݗg�1"��'QP���ׯgޚ@C��qn0��'��H�w���Z�!c�� �rM��'�ĳfC��8#����Bi:�]2�'BL�ͪ���RgI�m	Vp��'L������,D�H�`�Tp��dJ�<�Y`4\0�iӺn�V�Ff�M�<DV��hmx�e�9���ᓁ�J�<�0쓃m庄�t��:m`��z���}�<a i�?Z�� ���>/�)Z�b�<Q�k�"9�y"�Y54h{ׄ�]�<��ɃF�P����6�dR��G�<A��޵s~�|z�nG��u�p$��<I��-����� ���a��~�<�`1פ�aV�0���Z}�<q�c�(�^�c��ܼ*�(0��@W�<�Ƭڷ��)2Ǚ?�>�+��Y�<�Fϕ�Od��"S�@�Q�[b �U�<��n^ �6T��%Úg��![���t�<�tiU1I9�Hc�` �YT6}[��Ty�<A��@��L� )�f8	��@y�<���95�Y��l��I۾�_�<�!��RI��b�6�"�A��A�<����P���Co�h��t�Sa�{�<�G�+`�n��J��:p��ąv�<פӎ.��@f�^��`�w%�u�<�6�˰5
���ғseT��Ev�<Q�K�D�<�,
Yv�=4�Yp�<�Uo����Q$Ǥm�ko�<��'I�y�0��l���jW�^f�<Q�N�h�����B/�Z DOW^�<�#\�x�R�� +khũ�Om�<�e�A'xDBB���&��eqM�<�ɗ�\Le1 뙢]��)g�\�<�k)1ZG�xcx4�T�TY�<����6N���c
*��	��A�P�<a�!��QS� ��e)Bˑ�M�<�3D�l��2w�K�G���փO�<Y�$�	9�nI؃�_�d:A	�K�<9�L� g��@BHW<��ҕ��L�<��nK<W$�Q
	�X`�
��a�<1�ۢaj�[6�8g���2u�
]�<�
����6Y�#�&^B�<aǡM��&��l�0B���K2̀v�<i��B�[))p%`�]��{d��q�<A�+�3
�hi�qaܰ�.5µ#l�<yL��&����A �,i�H5m�i�<���(�}�M��7fACV��L�<�uF�7f�������iI:�
')FM�<�BD�h���#0+�+N�`��GR�<�U��)$� �	�S��D�W�p�<QR��6~|����mZ�;]@�H�Fo�<ѣ园^�r�2EM�pӈ���^h�<R�T�LX�d(��W~6U�H]�<ّ,�.>�xhaL�Ɉ�a�X�<��N��Nx�􋀻lwL�+�aWc�<��dEQ]�s
�(�1��p�<yw�ą}�n��ġ'9��dK�q�<� �=Ѐ�èk��=����`D9�b"O�䋤-�k+Jp��\)�xzf"O����ƶ6������ʼB��C"O���&	�.!.����oӤ	a�"O��pJ]�9���A֭��0���5"OB����il��!4�(�p�h�"O��քI�Il@�dK�_� ,�"O� "�e��J�'.�F�� "O$�&�)= ƀ��b�.3�P��Q"O��Va҇/���r�<�n���"O<�h1���~�
,H )[��Y��"O�Q�v͐�5����B�5�4�(#"OB���{�l��Aʡz�<Hv"O��	����Ĩu���:�$lS�"O�!y�&��o�HaH#6@�0�"�"OR0��0����Vr��R"Ov�QW�%<E�Ad�xB�hG"Oi�{�H�A���6�Vؐq"O�9�'�L�%�@yPm�<f��u{t"OD��*� 3�F�x6M��\Xd)��"O�{&�^*[�d㠌�HF�D"ON�s��\7%Sh|�V���nl�0r"O\e	�؃6���j�G�$F{����"O(�"Ø w���rS� c�\X�1"O@�y�֫+���/�_䔂�"O ���/@�Q�	S �C(}D�"O(�'�=H���#d�5nWz ��"O��K�a߻Z����]=��	�"OLQ('2��3Ck��Def�r0"Ol ��[�.�bJ]�jf �'"O�t� ���a��ɛY�t��T"OP��G�98��,znM?k�ڱ�"OuH�h��sMұj��3"O~q	��Hu`�6���zDJ4"Ozၔ���u$�@pqiD�i@���"Oj�i�'p8D=���B?���d"O�A"YC �* Ǆ�<��$��"O��27��^�i ��\����"O���?!��L�$�K@�4Ҧ"O�H���/5}���wm3e1��C�"Ox�Q��
C=��C�L�n����U"OV����>y9���PACqy<�#"O`��"�D3���O��S��h�"OT��5��)�]HA��K�<�"O�d�E��j���4'^���R"O�d��B�:CA���o�/Xbe/x!��K�>�X�v�
tr�"T#:1�!�_�/�a����?Aȱ0QBG�0�!�$^�fk|�9�昣]�`�c!a!!��l�2�@�]�(�H��Aʠ�!�O1������Z���r��-F�!���<�W��6��s2N�>�!�1S��-���@7%�R����Z0sx!�D�*ޮl�� Q!x�0�P��k!�DY)E8�-��������<|!��߾uZQ1�LK��9���!�D�F�� BF�M�p�ڦ�Y�"�!��J#"Y��\�J��AOS
|�!���R%⌂��t�l�z�/�� !��>.��ۤ��1yL�S��; !�S�h@�쌉^{�9��.��,R!��}"l���M�Z\�A��My�!�$N�؈�c��+k�
�L��+�!�DSJ��Z2���Z��@+M�8!�� ��[ +L;8��۷�	b�� ��"Oҙ)�l34Ȣ��b��&P�g"O��P�%�L24ы�W ��"OD���/
�+�r�y�MˈET詓"ODE��mG�=�.�n_�7�"O��9���O���H&�D���t��"O^x�a0w��l�&(\<���h"O����ZtT������7T�\P`"O�Ա��CX|��H�;;�X�*"O�|A�D�Nl{� eFܺB"O0)�T�$X"��{�/��1��)�"O�,� 	�8򔫴�Wg96�|��)�Ӵk/L@�Έ%ݚ���Ś!i�B�Y�z�Z'�S���4��珍<�RB䉥J�`�hg�>R2�����y$B䉡>lܴ�u�_-�<���O�	�NB� 
�r0��!MV��1Lƌ�B�I�D�P��;���@fI�f"O 1��G��E`� B= @ի2"OH|b�C	r�liU5߸�ȶ"O\ �Ƥ(LL��C��0Ό�b"O����^J����ՆZ���)D"Of���^#Y�lLR N��9j�4��"O��X���=6,�i�Q�ٙ)�T-H�"O(Qс�ڨ�Fmp�8pl��V�	��� �"AT�n�N�#�.f
����������	�N�;$҉��..)H:�XA�x���\S�O���5��V�[(�9�o�,89x�V��J�If��|�>�u��?���E ͶV��2��Zᦅ��7�S�O�F�0���
&��y��،uD5��)���x�!h6E��'ʜ]��Q4�ϑ�y"�d�$���jIc"MϤ~�}��,��s��_6	bdKǠ�q�8��OGP���߻~��	�FG<Y�
�ȓEs5c���!?,���gLL�%��%�ȓ�(���_*Kb���f_a�~��ʓ2m��f��@kX�i1�.e��C�=hMJX���A�88�c�|C�I)u5GZ2�c��r� C�	�j� b��J�u^��v�(,��B���d`�EH��4	�C�<0� B�I�ikB�`�æ~1�ak�6N�B䉢*��Cs�p]ا�ژ��B䉋�V8�,�n-*��ֆV*B�ɮ~BtX`f�Ĺ8��:���W"B�@����t/M����&�W;~N�C�ɺ�[�K�+B�Ⱥ0)�Eq�C䉛HZhɳ"J�	�=�H!w�RB䉘[𹱷cŮ9�t�#B���ZC�ɝ������9~�(��/?PkB�ɔjl��
�f��	���Õ��'nJ�C��$":	��(R��A���C䉯V�e �� ��#5�4?B��)5x�I��K%bݴ�3��J�B�Ir/�@(AG�Abr*:O��B�	#(�m�P�U��!�t*ː<|�B�I�l�� qR\�)��mk��v~B�I�m*��u�U�o!^��r��=�BB�I�jU�ds��I�-�~W�v*�	�'��E�Ū��i'R)۵��Zh�
�'.(s�Ӑg��I
�o
��|�1
�'R���.Y��Rh������	�'�2l1��(ڥA���԰Q
�'���H�ˇ/>瘈 %FE;t���@
��� �H���re<	٣hMe �Q��"O�$��$ �yBm�HӃQ�tTq&"O�H9&c�#$$q{���j��7"O
(��L[,���c��� [Hh��F"O�<���%T5� �@L3E0t!�"O6�)S�E�==^�����%!?F�:�"O�8d(^/;��u/��}	���""OX)؅�sĞ��v.�?dKz�x�"O�XU(�b`P3.��J��5"O$<�Q F��]Ґ�������"O�,�5�ߔ�&���*RQ�*���"O��C����	�mq4�Ì}\����"O*�PE	��q �Y"4���&r�#d"OR5a���Y��D;�(OJj"OdH�Q��P�d��!.�髆"O�%X�ԟ@����a�(Z����"O���GcI<$P�+g	�n���"O.��5��jѪ<󐈐>�z�s�"O��#F�;��Q�Q290��I�"O҅��̓G���ʁ���F�z��d"OzD*�hU7'�2P ���<���9�"O���$甥muʐ�V��f�����"O���@aԉ��;�'2s��{�"O�(�$o��cV@3�JW�� �"O�86j_�)��iw����@��"O @���ӽQ9�%)1�Ñ-�x}R7"O����\�B�V����R.J���#"O��B�H	d4�+�Á=W��@90"O"��b'W�)�=����*�c�"O�@! ��
8  �eBI�Kt� ��"O�`Zc�L1�n�p�
��8$�E"OⰨc*[�i A�0J\��i�!"OZ��@B�(3DA;2�}"<��"O��Yq�%h	C�A��Hܢ=��"O�����Oj3v 2�@��K�6;�"O������g���B��<X�6�i"O��`�	�?��
֧ol�MXB"Oܜc�휧0�P(�cGM�syi�c"Ot;�ᚵWU`D�f�>�f���"OL�cF��p���_�-Ӳ5�c"O^���"]� �	�� �,�s�"O��`�$��wi\"��6J��@%"O�1{�EA�55%EV'F��"O�	s�+�/U%zU�"�H#W��Ѱ"Ox�X��H"���"�C�4)�"O�@��ɒ����3ŉ�?���#�"O.iAa��[w%Y6h�2w���*"O�Y��
�z�|z�AS*T&H��"O(h@��8>�CV!�?8��!Z�"Od�z���C]�t8�	P�0�r��F"O��C����2��T	\8}"�!s"O��*�Zmޝ��Ʈ��PR"O�SQ+�^��=��>���J�"O��1��! �1�Ƨ>�6�
�"OX\�J������Ƽk~B-	�"O(�*a�OȖ%@�cĴEi&��f"O�\�� �-ɦ�`p��;Ng�C�"O,�V�N(}inQ�u�U/-K@�X�"O�CM]/Z�J��o[8.�$2"OvI�Q%��U?�l�W/JF ��"OnyHP�R�x�kƺ ?(�˷"O2��G+Y�T�\C7��;,�]�"O$R��*x��{JZ
't0��"O����G��Pr�p���cH�I�"O� v ��F����a4�[=m����"On��1��6:�����"-�y&"OĈ�R09�tP&�=0��Y�"O�	)q�F�D�6�@�f�X��"O����(R�h��$�>1�y8�"O��i ���x:nM�ctUkA"O��a�g��b��d�$c]����&"OL����W��$�TBO�[c���"O!�R�N�&QBR!�<���d"O�#�
2]����� U�t
��H4"Ov`��F��I�t�s5 ؼܙhW"Oj�TO��<�bd�� �4�(0Z"Oޡ{�NT5馤���_2C��#�"O̽9FƱrQ �s�73,��y�"O��OJ�� ����аaC���Q"O�8{A e���еaݪe'�8�"Oh`(�BZ�qGU%��>�]r�"O(p�Gě�f=@��P�a�"O�)0�F�p��%blO.@jrģ`"O.E1���8�X��Eןe%"O"%�mӇ8.�:���F�0I"O��q�F�%n(�����r�H�٧"O��&OP5=Iθ	Fc]� �q�Q"OT=�CFl�9��a� -���`�"O8�s�CV���5?H���"Ox�IƟ2i�,�c�A�5.�Yjt"O	�ĭM�h	X���K�=y�"OfQ�a�,*���ɧW���Ӡ"O蕸�傳<�h���=.�5��"O�%����5 �N�=�BeB@"Oz�9aո;]�d W��'��TC�"O i0t���R�lBS&͝R��p��"O6)���_6Z`v��SjQ����ç"Od�y�m[�u�uz�
N�^�N�� "OH�K�G������"��IW`� �"O�4�Hܫ	�0�V�9I�@X"O((	W�)X0�L�� B�� "OB�@�Y'e�5�5"J3D'�}�D"O4قR逭h�Ȕ�&��f�b���"OB��gb����uP%�����!"Ort�'�
�.M�9�Aʃ.��JS"OH|A�o�Q!��K����~m�7"O�-����6P��`W�U��j�"Oz
!J��ؐ��.�J��"O�i�p��|jH�)U�X&6q��"O\�b#�
nq�w��;YCrH��"OV�@j:Gj�h5!��>���"O$�ʶ��V�$;$�h\��"ON�xU��:sT��g ю6_@��S"O�1�V��8�xI���O��(b"OzPZ��H�u� 	k �|���T"Oj��*M*���s�jڼ=#~��"O�x7��nt���&Mm�X�"OTp�Ej>oR8��'�k[v���"O@�� �G�����iQ3�:� "O���F�J/i����/,9��؈a"O9���+5�L��}�ZUkQ"O ��nTM��:1�;^_����"OZ!9G�M����b3�/N�"�9�"O�9��,H2+�Z�R�L�uMX�;"O�u@E�֝aSb<�r땬C>B|�a"OhQ
�g��u��,@C&e%ʠ"O���DaH��2Ɵ� �l��"O�@�� �[	��"�d�uѼ�U"O� �� �ސX��P��:�Z��2"ON� �L��X A�\!�"OXh��I�z��\z7��>B���JV"O����)4;�R�n�34����"O��I��P<jZ�Y"nY[²���"O�!�C�	l��=3c�J�#Ȝh��"O���D<f��*�kVf�@�""O`ɹ�'�;a����"Et���"O�l��%C%V^n����8Uy�$*�"O���:m�N�p�ʉ4Ds Qc"Od�x�L֩Z�2�Ǝ��5s@�l"O(-�n@�o\@3ȕiF�@�"Oh�3��^�	�Ua�m�U$$��"Ol� jD�� ��j�g�`��"Ox�8�G
�\�N��l�9vu�lb�"OJ��.��d
`�#����S�rp��"O��tGX���Ѩ�*!	v"O�-�l��N�b���Fy�q�"O6�ѱ!T17lD@A�Q�a�̩b"O"��J�-6�.��ĭt3\r"O��aI\��qGT �!8"OȘjMW�D,�0���=t�Պ�"OR�i�+a��X�@���>�~��A"O�!S�d����Q�g�����g"O~��áҧo	�E�T���L�y"O&ъq֏�¤H3f�(\�@���"ONX��R�T��恘H����"O�\b��0�� ��\���	�"Or1�Ud�9<��1i���G�<��"O����,%RP�BᇔRؒ���"O�(QEBrvR�K��D�*L�"On����Ў;3M�%�:�╉r"O"�s�' ��DŅ�
��x�"O���r���v>�{��G>]��)��"O q����(��9zT#� ���j�"O�k��ΏA}�X�C�'l���07"Oȸ�   ��   �  ;  ~  x  �)  5  Z@  �K  �V  :b  �m  x  �~  g�  8�  {�  ś  �  T�  ��  �  \�  ��  ��  [�  ��  ��  ��  E�  ��  ��  ��   t � � � �' �/ �6 2= uC �I  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C��I����á���[��.�{c2��"ORH�^�Ua���C�xb���!"O���㫇�(�<��[1oT�KS"O.�s�
�jB��([8(T�� "O�DRG�X- �R����P9S)|�"Oz���OJ:B�ppP�mղ��t"O��� �1d����E{d��y�"O��@A �.�d]ʓi�9SJP3�"O��ceV�xt1Q)L��nI�"O�	Y�/J�,D���nV3���)6"OXsO�*ZUp��'m#}Z���"O�]�'��>�<��s�4\���F"O��x�f�F{�lqA�ǵ��x�"O:���ǧe����fO��I�Z�"O���EH�)IݪM����2'D�Ű�"OPl�#�O�/9�M�-�&t80"O���dC��H$5˂��<$�s�"O8��*Hza@�-�%r�P�A�"OrAsl,>|��s�b�z��tZ�"Ovh F�7O����) �Rq"O�43�ϼ9��9D���YQD"ON�r�a�7%V��f$y��t�e"O*c$A(򨹷e�H�9�q"O(��gj@�$�� r�BLz��9�0"O��D�ΥAy��ʁ� 6���1"O>8��`��m�E�@�.�8��B"Oi�O1�ة����i� ��"O`�H"��$��a���:u��$�"On��DP*<�����nA�N��"O �K��{a����-�x��A�"O0�x��ԀoR���7��M]��s�"O��j�d�~���4�	y�$dB�"O� �����#j��5CX@�, �"O��b1���_2��p������4�Q"O.��A��(��L1ӯ��"�#"OL��CV j��aΌ.Ƙ��w"O��+BO
5=�h�@�퍛D]<k""O֡`Gh�7u�����c��`��0u"O��Wo�0��D	�"����}�"O�D��f��+v���W�d�6�b`"OP� Qmɀ]�R���a���ł�"O.��f�P޸��!�+�p�0s"OlYP�%��!;䠝�/x��ZV"O��;��B��9F΋TT�]��"O`48Ќ��S
-�sW�~Z���0"O>��o�R�bG!ܠFS"O��U��(N�xQQW`Z�z3��I�"O|tZ��� S���-�����~�!�$� ~�I!��:4H�j�49!�d_;b��@���9?)�\���/>T!���!g���CqɿlP�CV�]3!��y%Y�.�4a�)�I�>H�!�d��#�6�P`��2�D	+�H�[�!��Mt����9辰�(R`9!�Ā�v%8=*��f:b�U��G7!�$�u��ਕ@�l.t��6$,!�� �����$J��*���,!�d���`hM�� ��6��1�!�ڏf��U	�������(̍�!�*�R�Y3?���x��\�|�!�F�S@��H6E@1~���@�$�!�A5�,:�-�ds�\z�gN0_�!���#I$�T
v��"_�t٢G^-�!������EL��h��D�G/!���(@��H��/ ���bA@ V-!�D\>_�T�1$d�=*u�
@��~!��(�V4�e�(3���qAM=+!򄓃E �=Hv��00��)�s�B�x!򤐌gnѡ�.�(�x��MC�K�!�đ�X��u� �N�9�@HR�̐�U�!򤘔k��Q$��}�ũ��H�7�!�$�(�����P�.��:��Y�!��\!<��M:5*B�&wR��
ŮVz!�$�k����+S&r��b%�@�b!�dͤ8��� U��Q[����ITa!�D�')���Kغ-I$�;�" �g!����O ��r�G�Ej)���ɋ K!�V�$������7<*��S0�{<!�$�;6(�p'�3(&:iЉ�/+!�$	K�XJ��֝O#�����= !�d��+.�غ�R��$d��L!�D_/�ԲT��6(��H��B͆[!�$��X���0�BɊg�$�׭K�!�����T�GL��>4J����4�!�N�v� �S�ˌq��5�]ȹ!�"O���#Oo3V��i���Dh�"O�Ap�eݦv
��'�aq�"O��k�Ad�FAb���`e��#"O�A'�� r�@�(A)�&�`�"O���pm�l��e��3��#"O��M��p�$�A�S�j��5��"O��J�"2~�J�f@�*4�9@"Opij��;[�z}�%�X�����"O��Q���%/;�t�Uk� �� "O8���ǖ+GК4Z���|.\���"O���f�$p	�)�Q잊)ʹbs"O� ���2��|�n��J۔ez�Q�"O�ׯ��k�$4�̗��A�b"OF��f��[r:l�BJ�1^�ā�s"O�P9c��
>���HAgL1���"O�jU-�/���PF4^����'���'_��'�B�'�"�'�'������~����F�PCt�j3�'7��'/�'"�'�"�'~��'9��	�Z�ds��U#ݑVnrP�Q�'���']��'���'E2�'d��'�2��-��,0��Ӕ`�� $X����'���'�'�"�'&��'.r�'����P�H����dB�z(��'
��']��'���'��'���'����_�0��aQ.�+)n@u�'�b�'���'�b�'�2�'d��'͈q�H�
j���Ӭ��x� <���'�R�'�B�'�b�'���'�B�'�j�`�+N&[�Q�ס��#��؇�'��'2�'�R�'���'�"�'����2�ӊ-�J����("
�蚢�'�B�'���'���'_��' �'��8�D�(H�P/_�>�0���?����?q���?!���?����?Q���?�riļJ�����\L�H���?���?��?I���?y���?��?��L��z:�y�f�LSN�����?Q��?���?a���?��?����?!�	�Ld�������H8dpz�=�?1��?Q��?����?I�9���'Bb�-4NR�� =l��c�$� 
 D˓�?y.O1��ɾ�M�������きA�C���p�ʦ,��i�'@�7�"�i>�IƟ8�p�ȅ;���
V9t�����	�,2R�mZW~�0����N�)�"�J�G�٧z�P�{�"�R�1OR��<!��	��R��P���.Q��	h������hoZ�V36b�D���yGc�.:yz�x���|��h�
�ut��'��d�>�|�pƄ�Mk�'6����h2�iP��g�(C�'L�����`�i>��I���(F��:B�(	А��7�V�	Ay2�|�%}�T��T���4Ah j��YȽ1a���"��⟤3�O��d�O��	Q}�J�2o8��Q!��"s���4h���$�O.��)خp�1�.��p�\��Em��W�P�oãHҐ.�"˓��d�O?�

h�֠��QJ�|x���b�����M�e�[~�gӄ��� -��D\�|p�$@OD��������	ǟ�����'�	A�?]�2LJf��B�o\�2!F`C�c(1��'"�i>������ߟl�	.$�^�����e�pɸ@&$f���'p�7MI�&˓�?YI~��^�`�jF�9|�)r�J��S��Xۃ\����˟�&�b>-KD,�5C|�
Ej�; b,��5(B� 2z�mZV~��W�� �������DX!c�eB!S�'�d��j�i���d�O����O.�4��˓���F�N��&��9�L��T�0(���F�&o"�k������O��$�O��$�J�B����F��CKŋ{\��"�.��P�旟x���D7���������#����iˠ!�W#4�bA�0Oj�$�Oz��O����O��?��+�d)�E�����-Q�%���Qy��'S�6-������O,�n�V���� g�����c�c��oK,u$����ӟ�S�u�nZZ~���-:8�lAu�2�f�sB��;D�q�"�W?M>a)OF�D�O��D�OA��H-b���b�{_�R�G�O��$�<)�i����$�'-r�'U���
8�P$�WzJ�{E��/���w��	џP��Q�)q�ԮZQ�8`�뜞 ��{�+W�W �*��̈́��u���Oڟ�� �|�ƈ�m� ��ĩۡw�X	�$U��'��'q���\��P۴�V�����-	G��kR�a�v�����?��C!��$HI}��'����A��3�>=yf�
$$ ��'�"B
)_.�������E+OK��~"��
Ij��[Y$<��Gϑ!PL�Ĳ<����?����?��?�,���p��_ߎ�"�K��g	f`(��PŦ0'��П\�	Οh'?�	=�M�;r�t9[�`��U}J`ag��#T�� ������On �iP��`c���.Q9Al��%n�?l6�d �`�=��^�ԒO˓�?���Hq��B��R�R���50KP�`��?����?�+Ot�m�GTJ��	ߟ�	�{��sb��+���3IZ�PWRp�?�PZ���J�c��x���$x��)hGoB�tR��'�]S�ǎ�c��������џ��p�'�pT�@"�(C�vx�D�]hxf��'d"�'db�'��>M�I�5����l� r�,��3�:��		�M��Ǉ���D�ۦ��?ͻo�`'��!qP�!g�S�I1 ���?��?F�7�M��O��Ս���T3�.e��'�
�
ti�#�1Z$�'��i>]��͟x�	ݟ��	�ְ ��Qya6�Zt�U
$�4a�'%�7��:�T���ON�d/���O�#�-(���o��ju�
U"Qq}��'+�|���k�v����s��A{�+�$΄4 ��Ӽi���8=Ұ��O��O^ʓB��u��R�&���s�+_�A0���?���?)��|�)O,nZ�"�	7F�r�h 	�|�v=��
ʽ��	��MÉ���>y���?����
���X�(�R�+Ӑ0�*Q�f�B��M3�O�8�E�%�(�t�� Z`J�� Y�zqA����P27OZ���O����O����O��?����G${u�����N�8R>�@�ň�\������ڴi&ͧ�?qa�ie�'`�̀��Rp`�n���A�Z�	Ο��i>Q�V��Ԧ��'a�t�u�W�Xhd<:f�\c��*F��Emx�������4�V���O���;Q�6@�_�ഴ�q�*W����O\˓s��� �	f0��'Vr[>���N��`j�# ����͘�B'?�P�L�	�'��w��0�%-��M<l�٥J_�%��Xqw)�o��=��4��i>)���Ot�OΩ�� H1��K�o��SŌ�8���OD���O��d�O1�*ʓ_F��.�gw攸�7|ώ1�@!*�y6�'�R`x��;�O�����>@��8I�d(���/�0���O8��Ll�0�ӺK������<1���6	쌝SP�_2}g��)���<�(O����O*��O��d�O�˧/q��X��М_bL�m�d��@צ�Y�M�����T��ѹ�y�⏑zB��@�"���$�N-{K"�'�ɧ�O͆%�7�i��C�)RRA@�ˏ��0Y3E�V�~��>�ꌉ�Vn�O���|R�XI$-Ӂf�[�&��}��Tz%#�����I�4��qyR�lӪɫ�/�O���O�1�W��l���S�H>nQT\Z��9�I�����O��t#O��/?@���+�'t���0?ɳCQ m:DaZ!�����'j8N�$�8�?yU(��z\��Jâ�ud�Ya�ǳ�?1���?����?��9�N��C@c��Y��&R� mL=�r��Ot�lZ�g(�T�'�P6M6�i�m�!O%v����`�I1&���I�r����Sy����PțV��cb�͞58�tOT7w*�AWN�T��=�'nL�zlLQ&�8�'���'hr�'���'#Xʧ�P��<xV�F.ӸXV���ݴ�t���?9��䧱?)�
�2�ґ�`�H92�������I某�	^�)��-v�r��},vcU�:F٘H;�E;�D��'�bR����8�|b\�x A�#T�Ix� �+����Ԍ��d��ԟ��I���gy�Fo��U�T��O
E�qjր_1��0���>�x0�5O�l�~�\�	� �I�1,��qr��
[#���"	B�Q� H�Q�q������`+�'ܿ�%�;mC�q;�� f2ڄ��j��<����?	��?����?Q���N��5-��JG��&9��x��4q���')b+{�8�4>�R�d\ަ�&�`뤦F�KƲM�`쀕CaX� e�v���,�i>]���WѦ��u���w�<3�k׊D������]���h7�'�v�%��'cr�'*B�'���`<��p˂��Ix���'H�[�D��4>�fiP��?�����I+s/1����&�؀{��;��	�����O^��0��?�
��o�2%��J&r�" B��+]T��g,!s�Y����S�XGR)N�'&��C�ϟ; ���OA�0�d�I韐�����)�{y�il�p�ɔ��f��Tia�V"D�>��4!H����O�4n�G�]��	�x�EN�R_�a�«��f��	�q�؟$�����n�c~���}���Sy�)�C�Y�E.ѤGA����*���D�<����?���?A��?(��p�rE�G�\�z����]��-i�
ܦ)��-S˟(�	�P%?!�i��N��_�$�P��01l�q���C":���D�O|�O1��5�P�h���I��t�-����n�,,-��(S�l���5.)��d&�D�<�'�?�Pf�� ��u+�C��}�V9(b�'.��'%^��9޴9�^9��?Q�IJ��C�L\�z���0��iy����B��>A���?�H>1&��]����lU#������K~�#ؾ0�d��(ǭ��O �p�I�$���B�z�$��'Ƹ�tU�ET�,��'>��'�ڟL�Q���E��ZPَ)�n�B��柜9ݴlQ�$���?�r�in�O�$Xk�L�F˗?n&"9�҂V"��$�O<ʓ3����4���#4-|�	��ZkVpy0$�4N���f�3��i��K,��<���?���?y���?���̃�8�oO�
�X��	����d�����6��OX��ON��^�D��m��겊]�k!�T��������',����XK��OC��(��>�"i��K�5�8ʓ�T���I�OR�J>�,O��$�N+鞀���W���E����O���O��O:�$�<ɖ�i��Q��'<����&,��T0q��8������'�X6�;�4�������`�'=`� �ڏz�h��`��2D~������{��&9O���Ώ�nȒ�'�d˓����U.B��bQ�dH
�b��y����?����?���?1���O5�I$BS��P��N�����'���'�x7��1����O(-om�	�@�p�"�����6�A�b�l�x%���������� n~�%�&\v�3+�^ZI ��D�S�E�A�?�H>�(O,�d�O(��OB�"� C$	d� D�H(	���{���O���<AԽi���qU�4��t�4�#��ś�� '��~�8|��O�(�'�2�'�ɧ�ɞ�WĬ�)�"�>��	�X��	�A�X�|6m;?�'V"f��G�=p�D���E�4�`����-Em�5�I���՟��)�SEy�Ja�e�U��1*����8>�I1s�zԠ���OH�m���q|��՟Z`\ :"��b��:5^�s�Rɟ��,&��LlR~Zw`"�c�O?^���� �л�i��xV�Y��J5Ͳ� �:O��?q���?���?	���	�Gr�}���`j�R�+T ��9m�;Hc�X�	̟��Ij�s��)���s�䕑����Eؖ$&��"A��=�?����S�'�Ա*ڴ�y"�/E�E�B+�4-�~\�d�G1�yBd�,�@A������4�j�
(�'�=֙bD��5Z�$�D�O����O��=���F�B�'�^y�J4�$�%A��J�9e��O���'|"��	w�"���Ԕ;��0��S.����)A ��e��\=0Y&?��5�'80}�I=��!��I�w�L�й#��0�I����ğx�	m�O�b�g�8���0�3&0����'DD7�@�#a�˓Pt�V�4�\�T&1Z�u�E�3�~�r7Ob�$�<Q6��M�O�i�������T�]��2u{�/950�6.O~N�O��?���?���?���v� �Ҁ�_�4ܸ��I*p��!-Ón�5`�P��I�8��m��|�H�^d�D�E'RYj������$�O���=��@�C1R���D�=�ڀ
e!\v��['��O*�ɸ�q���'�TL&�|�'up����b}~P+�ł�;	b���'���'v����D^���ٴ%,��g=ʃ��\^�%�ᨓ%f��ϓZܛ��Dv}�'�b�'�X���88g�#��R�Jl�8r�	ՏT�v������V�Q>��]�j�܁�w�F�sѶ��$>M}��I؟l������៌��O��S��3�V\Tl�ݣ�J9���?���̛�H����'6�$��/Z�z��e��O��)	Xt|�O ��O�)
�7%?�;w���h��Ʃ�l��Q�<a=�=RUE��?��?�$�<����?I��?9�ϑ�M@F�dӴ<k�Q^�?Q���dOҦY���Z�(��ܟ��OV�)p4�O�U硄�^���Cg7?�_� ��͟�%��'HK~��"ߎ/���Y��]N�\��$�>����ٴ��4����'��'n|g�M��r�1'Ί7��`�a�'m�'0����Oo��M�%��g]���t���i��p��	�)�~�c���?�@�i��O�A�'�CE�P<��:C�U<����F�@�9~B�'h@�i��I�e��lqe�	N�dY� 1o� 9w����&_&ak�d�<���?���?���?�-���p(��M�|ԉGҰc���x3ZƦ!��ϟ@��ӟ<&?E�	!�MϻF8���S��0}��E�;,�^i��?qH>�|2�I���M�'&����ŉ^Pd	�)��wyN�ʙ']���D ןDx��|BT��Sݟ�p��R/��M۷#�
��GLɟ��	ߟ0��NyR&q���-�O|��O�|8U�ӰE��٠�4N�NT!j*�	�����O���=��ه&:&����]#,�u���_1T��ɻFBi����:L~b蹟8�ɇ	ŀl�P�
2|!��>'{0�a���$�O����O@�}��Y+b �va]+��<�%K��������i���p�[��y�4���y�`�r��Ę��%i�yA䔚�y��'r�'alkB�i���pjD,1��O�ʥ�b$e�$��o�L���z��Ey�O.��'1��'�2�Q$T=x,2�ʈ:GBd�tj^�,N�I=�M��ǜ �?a��?9M~�K�X�o�tc��qq@ �m���Q����۟�$�b>�`���e��y��}�t�v*�2e�r�m�K~��Z�tĖU�����D#J����J��0��$+M�v��D�O����O��4��ʓ���(b>��}�.D�e�ɿR@��e��^��bb�@⟴��Op���O����4y	(��R6 ���(�d��*�c2�|���,�,���^$�N~��;HA(Q��
Ш6���K�n�&�ϓ�?���?��?9����O�����)bQ\lZdR��b=z`�'z��'=x7���i�O,�l�O��*2H�|H�Ȉ'50�A��E�w�м&���I՟�S=mQ�o�~��7��8`�C��m��4��(��"��`�V�|bX�������蟀ѶMK18�p�ҁȍ\��@s �Nʟ���Dy�Hd�j2���O,���O��'����&`ޓi��`	ǥ�kk��'0��?a�ʟ ]�#�[�H�0��b�.=��"�%�dk/�O��|Ҳ�O$<J>���\ڶ�+��1hd�S��@=�?a���?i���?�|�+O6�m��z�zZ�	�E�l)�#�2 �)au�G����ɥ�Ms���>Q�<x��zA��pP`�aڷM�e�0˓L�h,��4���b��I���۔��N���$R \�,a��/r>��Γ���Of�$�OD�d�O��$�|�Շ�'�^@df�l
��z����sQ�f'Ӫh���'�қ���'(X6=���f��'i�1R�'O4
Ӵ��Q)�OX�$1��a�V6M~�$�T
�a�9��͑hqD��`�q��FHЦZ�d5�D�<Q��?1��AFL�D�O�
�+�FN��?y��?������Nۦ��&�@ş��ӟX�����!	���cAif�q���$Tv}r�' �|���70<q�Qi�`���E������3�ԘI��Ľ,a ����q��)a���~r����*i��!�, ;T���O:���O&�D%ڧ�?��혪Ev� AN$_�ެ����?���i�ʤ���'Z�{Ӧ��� ;��iR���#&�ȃ�a=�(��������LZU��̦��'���X�e��?Ũ� ���O4_*�+5(�>�`I�� ��<ͧ�?i��?)��?a�/J�>k8B�CȤ��t�����FĦ�!�[ϟ��Iܟ�%?��	�=��%���2zZ���ȗ+n�<��O����O��O1��(ԋ�*8o������$Ty�*��i0 �҃��@��)տ��~�IybU�<�#�)K
_� ��`�A;"�'��'/�O��I��M��c���?�G#بk�`��F+��=��B�J��?�P�i��O��';��'���TL��v�>y����̉Xd`��i���3'R`ys�Obq����Ԥ{�vٻq",I�hx�@�3��D�O���O���ON�!��� ̜��a��?��S�ʟ�V��	˟��	�M{R�
���Ϧy$��H@�U+q0@4]{'������J�I蟄�i>5�G�ަ=�'"@o�y�cw+\��hRs�҅m"�l��s���O���|*��?�"u0��+��?�*���σ��������?q)O�nZ�O����ʟ���D�ԧ�F<�|A�D��
�P1�+ʰ��$�i}��'���|ʟ����'ګ%�:�v�Z?$�hŠF%�}8�WH� h��i>%0��'��]'�83a˕,΍�����X�x1�M��� �����Ib>��'��7�˫0�H���,LBO�M����!5<h��<�p�i'�O�M�'^r��$5J(��,߄kT�B�� 'r�'ߚm�2�i2�i�A��m�?)��V��[񍚾J�)c�@= �J��b`���'�B�'���'ib�'��	D�@��	&Ah�"�� ��-"�yk�O(���OV��.��[Ѧ�]�,���RA�ܻn
�rf�s�:E�I���'�b>m��Gئ�ϓ#���OE���ԁC��t�̓,��d9�-���%���'z�'_�M���>{*~eZdiV����c�'�2�'�b_��ݴU8(����?���r~�X ��E�
&�ۗ �.��Ԩ	x��=��	����V�	�1�J�86�T98��ek��܄R�H�sp��QcP�4���|rA��O����&�qS%(&�j��%kV9����?��?a���h��$/`}V}�r�̱"�n�駨��P�:����Q���lybw���杤T2-��_�,I&gω9�V�� �Iҟ��1�E����'H���3C�{B�n�w��`� �7�E�$������O��D�O2���O���9-$tʇ��6�H����_O�0�s*��"�7<���'r����'��p��@�yB((P�@04�)2��>��?H>�|´I<�L��V�b$���&l�l�@��Յ�򄛰~�)�SĒO�o�<���M��c�bB��i4=0���?���?���|Z/O��������?9��4Z�p�`%K�] �9ŏ�<�?���i��Op=�'�r�'���;�|hCG�A�rd�p�B�u]�9��i��I9t�)��ޟ����.�����O1=����Gͤ����O���O���O���&�S�J��P�W�\��e�	5�]��ݟ����M����|��{���|򠙴r�l��$S[z�u�c�G6\�'�b���J)6���4h&�\:j��Q�V5T~d@q͟�=�B嫖�'�jQ'�����D�'��'S�)Vl�*A@���B��u��=pD�'�2V�|
�N��1��ٟ��	s�T�F)�Z�"�]L(��ANR��{}B�'%�O���`K��y�oA�h+G�H��<��,�Ҩ�Ц\cy�O���	�r��'�r(:0˕�W
6:%R�Sn�2�'��'*�Ok�I��M��)P:#����,ѧ�`���P<|Ѧ�+*O��o�G�
��	�8�4ǐ/�M��R".�8K �ӟ���1�%lZH~r��&G\2��}r@��/"����Ī^��9!�<q)Ox��O��$�Oz�d�O˧qj�uˑ-��XQ4��+��o^R�e�i��ԘT�'�"�'��O��Ak��.�_��	��&nJ��#�F��*G���O>�O1�����ce�@�I�C_X�ZF$ �It�����h�	�e؈4�'�|�&���'�2�'����V~Ⲭ1��S 5ȝ��'�R�'�BP�p�ܴ2�ܝ����?!�AC�-ȔY�.�΀ ���>Vx������>����?H>�����p{cAR%�`��#LR~�Ƃ�*�HR�����O<�\�I�ª�܆�!5)��aՏ'���'b�'���S��+�`��	�]�2��p�M��k�4Cք��(Ol}�Ӽk�K�*zN�٘�D�yt�eS�"��<����?���5'�p�4��Dz�
�(�'h�H����o���Ӳ�ļ A@�4�D�<�'�?����?����?A�nV�`�rp�D �:~9�PK�޽��dʦ�q⢚⟜�I�|�:�A*��ER�LD7!n�z���40������y�)��/�ؠ+�N
9�T��b���'��I��B�j�Op����O��(O>9+O����I6�e[��	,ի���?���?I��?�'��$�¦��"*T�l�í	&���։z�0 .u��C�4��'7���?!/O6X)֊�.M½[C��-�F��q�F S��6M%?e��T��	K���'���G�������^�Z�X�<y��?Q���?����?	��T�
2K"��w	�(P	u	�돱D��	�Tq�4c1(!Χ�?�B�iQ�'�ܩI�� z��	gE�D�ʭz�|b�'��OD��ÿi��I>wD�� �a{�b������(tδpQ�dZ6�~�|b]��ןd��� ��W T2�tó,�J�hUQPL��$�Igy���O�$���'�B�'Q�SQ@Xh��Xv�у�P%0���I��I���	E�)��dsh{h/7�|�V�IY�`�r"J�"�M;aQ��sQ��'_�'��`���>�5;���(A�+c�'�"�'b�OO�I��M�� 4x�!�^#8�Ȩ���2d
E����?م�i\�O�p�'R�1*[0�
V���81���)9��'��k�ia�IL����OD�'�Ґ3���Hf	k���(��<!,O���O,���O���O�˧F�8`C�
�(����C�pƈ����i?� ag�';��'���ybBx��N[w�d�3�W�5.B������*��D�On�O1��Mjd�p���		�`�7�@��4�o��7�T�1x�0���'�6�$�8�����'�J���%���9��@gr)���'��'2�W� S�4$r���?��XNy	$�E�2�����+� ��	�>	��?�N>��D�;V(� �q�<K�p���Pp~��6y�nu��O#ӘO�le��!SsH�	e�4��T�>5��J7%W8F���'�b�'e2�S��l)3Cȑ2�Bܐ�D$��=)��՟XHڴSG�����?��i�O�N���H��_tj~������d�O|���O&c�)f��� ����?�kG&�������TB樃�ɛn�Izy��'#��'�r�'�B�L!a�(�aan̕6���qc��5�副�MC׀ݛ�?I��?iO~�3�N��b���'���
�Z����8$�b>��4O�n�-Ǜ���j�%�
_+h�oz��]�>���륟%���'-P!��n�����s���R&�5�'���'Gr��TZ�|�޴?LЀr�^����Ԥ`��Fk�6~�Γ
����D�c}b�'�B�'��q�aܕ<�FDAEg�53R�s��#��摟Li`�N4rQ>m�&b���Q  	a`�Ԉ$J-���I�����ݟ�����`��Y��ň�3�eB8��n%
�1��?��C̛&�ϛ&��-�M{L>�.
A�>�yPG� *(���e����?���|ҷᑏ�M#�O����ʩ(Ÿ�m�*<�Д����E����'��'D����8�	۟��ɭ�"\p�M#%=�E�GiH�}����I̟<�'��7mK/h��O:�d�|�bi�)��S��6:��`�jP~��>a��?!I>�Od`���Of��M�G��-�Sa@:�|(ᕳi'`��|��é��%���-N�Er{fl^�pd�V-�ȟ��I�������b>�'\�6B�e!�]K��8G�Di2��[9�|���OD�č�u�?I�Y�P��0�x�[�
L8ONaH�><��������,�����'�V��@�'���Ѳ�B�r@�0�V蟪g�����$�O��$�O,��O>�ħ|2à˘r�@(���3� $k�e�+ �V�O��"�'���'ʲ6=�RX�%@��)���冥s�\��*�O�D>��IR�'�~6y�@a�*Tf���e�#�`��u�pa�TB�@�	Sy�OCb'�	�|%�E� cV�:�1VO2�'c�'`��&�M��aZ�?9���?�I�<<e�,���C�ccT�B����'�`��?�����gZ\ ƅ)v@ �5�GUM���'P����'8�������TП����'RT�0ҋ�nr���cB04����c�'�b�'l��'�>A�I# �	��"	Ö�z���b`�	��M۲ψ��?��%��4���8�ΟiM���ad��.�)qq5O����ON�I4"(�7-%?)奎�gKV���nF�*U�	'9�08��E��0RDx;H>�/O�)�Ov�D�OP�D�O�5����7 ���ǅ�)�=E� � ͛F�aU�'�"��T�'X�E�.N�%�-�5�C�'�E��I�>����?IO>�|js� c���4�3@9>���c�`��uBܴh��	�p\�w�O4�O��/m|!��J�Tu�����
mÞ�����?���?Q��|j.O��m� Z�t�I�q�Z5��K
�M+�(�N�/~,�扑�M��h�>���?)�AN�͓r��=�T�ŭ�� DPX��oR��M+�O �`�������w��M����W�\�[�m�y�B%۞'�B�'��'�B�'���9{@�;�么��_��<<	���O���OR�m�Z���Pٴ��_�����-��S���Z�I�o���M>Y���?�'4@�y��4����,l6�����M�u��ΐ	Z�uJG��?�D�1���<�'�?����?���	�6x��B��&~\�ff�=�?����Ҧi���Ɵ����`�OG�J��S�NcZizǑ(�"Xk�OH��'�r�'�ɧ��I�U���9�ˈ��ѫE����$��j̾�����}:���u�	���(b�$S����F�� ����ȟ$�	�)��hyb�gӎEJQ䀷9;���ŏ�/i����d�׷=D�T������o}��'�N�cn��h���,��w��1�r�'��BEW�����[�ƪhq������v&���lQ!F��a��3O���?���?����?����i)�X`��Ғ����"k[�	!� n�8�@��ӟX�I@�s�p�����'Ȇ�D+��B����]��A����?I���S�'�Ĉ޴�y
� �A�"��13 x��.�2+�Ȉ�>O���E��?q��!��<q���?���E?,q�%��GI�� �A��܍�?���?�����DצI��ş$�Iş��?:&��BG�?Ma�H�O��C��	֟d�IR�$F��ak7(\�+p��T��oP���"�SS#��|2�O���^��t��a�la��xᒒݪ ���?���?a���h�|�$׺a��w�Z�^`��=W�j�D��q��@͟�����MC��w��e�O�bA�i:פ��P��)��'��'O�� -Yv�6��8)f/�a�i�-�İ�)ݓ(y
Uh�	N(6�T�O˓�?����?���?���ӎ(��a�K�����"�L�)O��lZ2#����Οx��f�SΟ@@�"-�~���HJ ~����7��5����O�d6��i�8`:0{gM�1f}*���RdN�S�(�rA���S�ȴ���'%���'4��C�|z6�ӡBN*��a��9^��M78bI��5)Rl�&K�]Ih! s��$0�"�e��⟔H�OR���O.��\�A������@���@��	U�e�Zx6-?9AaJx�M�S��)�gS�lL	s ع(��x���i����	>^q�	�cJ�SLx�rr�N�(�P��IП@�	<�MaOXj��mt��OP=�p��1k��)	��ȥ\��6I5���O��4����")i�~�Ӻr�IM�����D6Dnr���Y/�����
N�O����'�$���P�<H"ɹ/Ȓw�����ڦ13W��۟,�	����O�2�2qSW�HU8!I
����O ��'��'�ɧ�)Гz&l��a��ll��A]�Q�=y%!Ψ������<�'2�l�$ۂ���q@&b�$� X�#�I<(ئɅ��1!�F$E�U�t�C&�8{�@1��*�%R��'gkj���ع�O(���_��la���\���UdD!�J�$�O�Y�p%�D�Ӻ���*��Ud�<a�E$R�N��dO	<D}����<-O&���O���Ov���O��'>�̙�Λ,N8�0���
�B��#�i�j�:��'���'*�O�"�t��nX�"qٚ�˭"L�E�')z��� �)擬`���mZ�<A�ă�.��kR*�36�Ig��.��+r��O<�M>9*OB�$�O�\CN��~E���6�+9^�gE�OF�d�O<�$�<��i�.��'<b�'��Å���2�RQꢋ�9�0A��$g}��'$"�|�J�,p]�h4�A�,��D��fۅ��DB�8Y�аկٶ(1��Ԑ��(R���&��]e�2d<vI3��)Fl��O����O��$;�'�?����:ܘ1�IR�9�b�Z������+\2
p��Mk��w�2XR�(J8��A��m�)i��E9��m7m�O����'(Mn6�9?�6a�4J����*J��2�!�4!S�,t�cK$��L>	,O��O�d�O ���OI�aJR�o�vha�C7@e�󀫹<c�i�Jm#�'���'=�O��.E`� �Qѫ��#8L�� ��.Z꓎?����Ş=B����υW=�D*�"�j���i�FS�y����'�%�̍����|"\�LyUAJ��*!��	Q)W,�+Sޟ<�	��<�Iӟ��ayrMpӊ��	�O.y�u��	[UF[f�3�Qc��O:�lH�-'�I�X�I�(�L�(F��xkO�)`� ��L7(w�lD~l�3E)��|�'��#2�
"-�ڴ���գ]�������<���?����?q��?���O���S��.��Փ��*b��'��)~ӆ��A�?	ݴ��*4��ೃ�9��!�FFJ7!�D�J>���?�'W�r�޴���
'&<|�p�"I ��٢Z�&�"��c�7�?��8�$�<�'�?����?�7�
���h�AY)5�x�e@��?������RܦŠ@aEǟ��ٟ,�Ozt{�'e�8�����NM���O�`�'���'Xɧ��J�s�h�%�PU�t-"P��>&ӮT�ƠC:[u@������t��
�n�-P����ה7�����f?�-��П���џ��)�@y�q�8����G2���<V�IX��
�cY
˓����D|}B�'lܪ�j�#�
d�e��� d�t���'��A�L��f����u�<]���<Q#D�Қ��c�E_��kB#V�<�)O�d�O���Oh���Oʧq�8�c�>n��D1�h�0@���ղi��җ�'���'���yb�h��ٜNC@y���;(PqQD�w���D�O��O1�̜�eg���I"&�\�CDF�4~tL�v'�":0z�59d A��O��O�ʓ�?I��3ډ�҃�~��ea�4Rܺ���?���?/O�DlڊGq�$������	��2l�%y��(���[rFY�����i}2�'t��|�ʈ�;�N<��	Ȩt�  U�M���$�q��A(��m�T�'?���OP�DX���D\%_�Xэ¿"� ���O@��O���0ڧ�?ir늞N�|5*�&��tsp�95�	��?q��'J�b��?Q4�i��O��2
Jp� �O�7�$��� ;���O~��O���«z���8�츑H�?�s.T�-���"�Ú==k��Cu�n��|y��'���'���'�BIF�j��V���bV�I��!U34��I��M3����?����?O~��\�`K"��?l��%ј�t�S_����՟$�b>e���3� Z0��	
<%1�|��+^	{D�a��$p��a�'�J�"�-l?�J>�.O�1���!g|6��-G7iT�񵣲<����?���|+OV�oZ:d�tl�	�E���Hѭq����H�7���I��M[H>ͧ)����<���Dqrc�
Z)�šҭB�����HqL��l�r~҇�#E����VB�OP�E�T����>դJ����y��'k��'�"�'����=b�$i�Uh�xT���_�X@b��?���i.t��O�2O`��OҼЀd��U��I�0��7h��x�b-���O �4�B�:�i���Ӻ���'nK��,ͷ/��i�$,��S u���d�@�O˓�?!���?i�=��0�ĥ�}��!k�-8׼����?�-OP�o�"'�}�'�BW>E�r�Q�cIbO�6��(�8�	?���O���1��?-��� �rAv�  &Ƃ,�>}`l[:�C��W!h�����NAן����|R�~�Di#��2�J���m��':��'U��t^�tHشtִ�� ��3��e�Q�U�`����5ʋ��?y��Eq�6�|B�'3���?��aB�F,��(�-�����O��?��Q Cݴ����%˄-j�O;��a`�(T�H�f0$eNn�IGy�'1R�'Qb�'MbS>�j��N�{�f��N�u��@�����M!Ȃ,�?1��?�M~r�T���w(8��S�T�f�V�΃&�QW�'�|���oC����8O�D�*Q�V&�ȂK�1P�%+63O%8cŐ��~�|rX����Ɵ����ο3�퀔O�+;��Y��������ݟ���vy�ni�Nݨ�	�<q����ᱰb�E�ʡ�^�R ص�I>������(��m��Q�8��e�&.��pM3q(��L\��5�G�?�D�ZI~J(�OP���CXz��# �^)ڨ�E�1�8Z��?���?y)O>�3P�����ۃ}�,+���y����,�M�ƅ���?9�;��v�|��y�l�\hH�s� � *�e@��y��'�"�'_D���i��i��%�?��5��02�<���`^0�h�PE�K�@j�'���ڟt��џ����x�	�;�bݢȞ�97ұ@���;-��ė'��6�������Ov�D<���O�B�'(�x��,F�Sxl�{U&�`}2�'Q"�|��$✿xu���e��Bhz�J���IuBM�,A���d5'�΀���s��O��#�>���g٨����C!GV�����?)��?)��|(O� nZ�_��	��e�s�A�A��c!ˣV��5���M��R�>����?I�?F0H	��,t�D�k�EW�E�� ��E��M��O�2�L͑�����G4�dX�d���REeЕ�"Y��bI�[X�qyq/!C`n��X�Ե��'� :����$>��<ؔ�W�'-�L�.M�	�4;��
âȐ��]l����7NM1e� �+I���A����!0�G%e��tA)�'dD���h	M��2�(N���ᙂ�ǎ��A�B�u��8�"�X"}<����i�"��u���%������R�nْQ	X�aܨ�1��_,a��uk�(�6p%k�>m�B�fх ����s(؉h��o̟<��ٟ�qQ� ���D�<���~�c�eߨ�:�iȱ�Z,wj���'[phV�|r�'b�'n�	`4�R	q2䛅� A�dI��w���$�V��4�'�	ԟ�%��XyN�l6*�	3�
��ө�g��r�M�O>���?i����M����l���B���C��!$��
�@ꓐ�d�Or�Or�D�O�L�Gd��<�ڢ!??"d�i$��9H4�Ī<��?�����D�l���'K�Hp"��.ԕ�V(�9�� l�Sy��'B�'V��'o~���O����
��IP��N)gTr$A�Y���	ߟ��IByRcԭ	�t꧆?�kȒ]O�M����?H|J�c0B����'��'���'Z�tr�چ�^�#MQ�G�Y %!����']�X�x�EHC���I�OJ����J(���,���"v#!y*H�����s�	��I�>=��?��O?R�Vh�cz"(yР'�+is� �-��Sմi�B�'���Ob���cV�þf�}�a�)���(�B�ڦq�I��(#s����O�RL��I%r�ЀRPm�T d�ٴA41aq�i���'�2�O��듮�DԄFI�xC2�V�}�81��@� f���l��Z���?Q����'d�9#��^p@�'΋#�0U��d����O���D�`b���'��I����}^��b�Q�.=��a��*����>��������?���?A�"�%W��+��L	��n@�i\���'�"�i��>�.O��d�<������5�9P���� ����{}r�ǆ(~�'�2�'_Q�t�u@����@�_�Đ�#A#b���O<����?�M>�)O뮗"�N@��h�E�:E!��w9���'|�IџH�IП��'�Mkb@g>�#U'@$tx��y%���0�����>���?M>�+O���O�`��4:��][��T�J���9�gG���'���]m��S��̂v/A��^e�-A��䉨Á�M#���'�!syO�i*���~�N4��Ns��Y#�i	�\���	�s�6�Oj�'$�\c��]�s.WnX�Tz� �s��D�N<������!F���A�pD�@@0D�ʸrUC�p��듂?a��+�?A��?	��+O�n¹`00*��T�PB��:�ť>̛�'��	� ��"<%>9�"�
K��X�͚���r�x��4����O��$�O��D��S�4�&� 
��RG�eX�<�T�ǩf<�p�U��8�	>�S�Oo�0:�nר
0�;B��3{�(�CfӰ�D�OZ���N�b�S�t�>� ؎��2#$.R}�@x���3^��`�����'.�D݌QVR�QQB�2<P�Cà�a���'::0PQ�d+���⟈���_�^K�u���ۿis�aꄇA �� ,5�<I����O�B�-O���ю�!'�B���$�K� ��?9���'��O���K�&|K��b$T !D��ֹiㆴ"�O|���OB�$�<��ؽ���D7�8THA4}�ډH�A�*��I����r�	ay�Oz2�>D.��Dn=q�l��bX�O����O���<a�!�85�OF.�f@�̬Y��LA??ͨ�p�Ogӌ��9�d�<�'�?O|:��O�M�4�&@6Aw�� ��e�N���O�ʓLb�:��d�'��\cV��V����*��t��>]&�-�H<�-O�D�O����`�$�.=��8��!o����i��u�
i@�4=��ޟ������3(�Pl3�=ad��Q��Ll�U������bK|
N~nZ*e�j�����nv��I���6m ,:��m�ϟx���,�����|ZV�Mg+]�MR�RՈ��jD�gI���'���'�ɧ�9O��ߊS�Dѱf,�m�"q{�iM0b�Im��@��䟌�B����|��~R�N��!b�O�h��țB��M����Qi�s���쟠��NN��k2��:tB!�5��o�(�ڴ�?�((P����4�'��'����7BJV<���Qɔ�$^�Y��'�d�O�ʓ�?����?�+O��`Aą�-���2B�"����4�$E��'�p�	��'�]�֝�.C�[c�-����b�8�7��O8��?A��?�(O��!��\�|�4*�����"k�5�h��C,HҦi�'�rZ�l�I�����0:<L��4JY8-��B�b�lxp��ưD����ٴ�?����?������ݛj7�5�Oy�l�W���X�m�r������*�
6�O���?����?��Z�<a(��6�<}&���F.��]T4���ը�M����?�)Ot�8� C~�4�'���O����EKOQ�,�$�z�r!Q�Ǯ>1���?)�,���O���^�Ƥ���S�2�ܱ!�+{��QmmyR���(^7��Ox���O
�	k}Zwm���/� +N�22�)H}؜!ڴ�?)�>���?�-O^�>]�eG�LI��#�hF)U7���lh�xhp�����Y�	ϟ,�	�?��Onʓ&Ңx&��Q	\�z�"#6��ڑ�iK�R�'I�V�0��T`�1qF��9�Nl�უHIz�	�i���'ve\:3YZ듹��O���&@�*�
�)M"/;X%i��&/�(7M�O:��Ȅ�S�$�'�'�*���M�"W0�$I����/@�%zA�rӰ�޲(�X�'<�I䟌�'=Zc ���q�ϐ<0}E�E R��dK�Oh\`8O ˓�?����'G��BVO�U��SG�]3����L F��xy�'#�����I̟HP$���H���
�<.����+q.��˟D��֟���П��'¬uxv$|>�S�cQlh�h��9:+����,v�bʓ�?�)O`���O����92��""* Y�ҥ̕n�Mx1&�2���o��p�	� �IPyR�_�rk ꧤ?�d�!�i��m�!� ���6�'!�I����ȟ�4Jo���M�R��Q���Т�ͅ3���0�Ϧu������',�Q�~2��?9��c^Ջ!	� �$�8��A��Q(�\�����Iw��Iџ��'���A�x�dEZp�� s��0`�
�H��_��j�dF��M����?Q���bX���?��5ᆌ��-��p�?_��6��O��$ړ��gy��i���Z����R5&������{��f�G>p-p6�O����O����N}�_���䅗�B�R3gez|RE���c'�x!�4���Γ��$�Oj�?��	9�Q���&��E�7�Ǘ_(�l�ܴ�?q��?�T�O�q���Qy��'���Q�t�2�p��7 ��(��C!���'��' �D�����Ox��O���׏�5f,ɓ��Q�Xr�̉�I㦁��	G����K<)���?)K>�1��H���=e�Zp�R�+�l��'eZ��'���ҟ��I۟��'��m��I�q"-��Fʝ���DK!q��O����O"�O����Oz����	Z�z�s��@w�X$�
�E91OR�$�O����<�W�](lQ�p;��	|���
���.]��p��T���	ȟ�&���Iȟ�YQc�̟�s�	�B�ڑS� �*L 
K���1��$�O"�D�O��V���������@X����n(�d[�D $6-�O��O��O��2O��'�������6r�{�����P۴�?Q���$�ڀp'>�I�?����IxD��bH�~��:�eO���?���<�a������C��,l"��D��|D��`Z�M(OB�2bG��!!����$⟆��'��}c$R�%(��@ٰlm�i�4�?A��gϓ����OJDh��#Ua_<y��D��p��y	ݴg� ��iVr�'Z��OB�O���æ4��P'-J�4�w��5\d n� R�Iu��~���?E�ш.{ ݑ�h;�\9�"E�xx���'3�'���`/��ݟ`�3e��; ��?Z�Pmڂ�S�9�=o�x�  ��zN|j���?���r���C�c[!i��|��c��"4�����i�"��ONpb���W�i�� p�7G�]�&�����38-�đ'[�,�%�l����H�I��ĕ'�!ƂN>Z�� �H�X x�-��b��O����O��O����O|��2)M}���A�])*$�S�T%/����<���?���ğ� ��XΧo�"�z��
%�fh��C7��'�H��C�I՟L��Bk�8�ɤYt��0`%�,3�v�X�)�1�Oj��O2�D�<Y����m�O8��	�ya��܀$<�E8�i�@�-���OB���3����'}�EI� ����@�V�R�@����Mc��?�*Oz�����P��<�S� G�L#����CJ�D��tJ�$;I<����?)0/���'��iS�����"�7B�M�!�˦'���P�,+gI���MSC[?u���?I��Oj! U��8Q����I�u�  ��_���'�"����J݃%_� �pGӦH�n�'�	�MK�n�F�V�'�"�'y�T�"�4�p,	ro�UZ>`b��|�����u}��'��O1����ˁ���`%�=sXR-0�=6�t!o�P���` �i꟤�	t���'���ҷI~v˲B�T��-{�[��ЀDx��#��O����O$����>(*��S�[��:5!ŦU��2O�zP��O�Q�OKr�'�����Y��	_ԼI��-�'Gؖ�'�<'�T��۟(�	П(�	=s�FYAMqU
1�$� 	01,81�cџ�	���˟P%����K?5��i�V�iT��J��ыQ)���"-?���?Y.O��D�0���`WB�����;��thɁx7��O^��O��O\�$�<7��Ϧ�����Z�|q��%��<�0P{�&�>���?y�����ձ$5jI%>��p�B-=���`��4딼hG����M�����?���dJ�8��Qe�L�fMlM�� ����'��\��@�*_&�ħ�?���0�hX9�)��p�y�b�˽id�(y�xR�'�R�V�O�S>Z ���Z�t�+��|묒O`��Sl6LO���  B:|�R!:�2�! "O`)�@�����n�8�����`�	z� ��@�k�\`H��F^��a�:��Qgl�,��(
uc�B��(Ai��4��)X�r}@P�@�(�	)0F���A`U���&���l��W�Q1+	L�"����G�4�^�Y�G�)�J5d2�Jb F��W25��	�G&�O����OP�dպ���?b�
:�h�eNA�Dx�>��pjB(��4�0�wE~���ugQ��s�'Q*�q;��;[� ��ޥ7P|䓷bP�5����Iڶ����"�j�0�ct�ɰJX<�X����*�1R�l\_ؾ�	+}�R���O�=�+Oh$�R�@�J��L!͓~w���"O�m�pNŰXq��@�	�q�}��ki����<��a�vۛ�M׭5���mʶ�!� �3_���'H��'l�����'�2�p�W��O��]!%X�Y� E��h0k���#G�k7@��V�><ON�����{X�5�$�_2��tOPk
,y*��c7<����#<O"u*��'¤��"��@�Ԁ]z��E��0	}ў�E��C�Y��1��]�,��4��y2I�j2��
[�B�G�2�y�,�>	.OP�2�YH}�'}� 9P���O	QpC�
[�O�މ�����	�tyFn�o�飣��aw�H{�S��c�9�� W�o8��u���(OP�����)�Ĉ��&[[m����3ą�?6���@ME"�r�ٲ�	,����Oz�?��tOM8ئU��eD�x�1d�}����I�t�6 ��1#>P9�QH���dN�ɦ]�9�� ����͒U��� Z�T� �O�d�|2a�
��?���?��Z�`���h˽X|��wꑽ0z~h3˛������>�Ox1�2��! y�8�l�'�h��'Z�M�������j�O #- �)��Sn��#�� %+�$dڀ�J۰3涕���������Kg~�jCL�&�\ѷ�ܡq�H �ȓJ�N%��P3'4Ι�!e�#�aDx��;�S�	U��$[��]�z�^��'#M���'pP2W/>R�'��'�\�'�?)!�<2; i�U��tr�p��hD�<)�]�a�\���~�� #�A�wB�=��@�`S4��Ň�)K~��
ƧP8؝0d�:/�^l�g�'?��kq�.u��[���'e�����'!��R'�'"b�o��Y����Ky�đ�|�0�+�-ǋv����%�HrN��R�ڹ@b	�4���H�\ nZ��MKJ>�,�rʓ{�����is�Yh������*��B��a��'�"�'���ϛp��'��J�>r�&<��v�T��	�7l�T"'R.x��	&�'��th��m�v���/�4:`�p��Oɛ{��ig(W�
�nѢ#�C-j�џ��7��O��%J8*P#"��1�q���DIn�şȔ'T���?A`�J5��e�v�n���z�A-D� �W '{V���KAV��1�I��y�4,�6�K�	-e��	6�H�^���x���-]�C�k�t���ơy���HB�G8[p��� ~yA��UG���!3=��'"O�����)��*�� �a�u"O��	���`��d[�� i9T���"O^d�WB�$�t�d�1L�2�y2�F� ���+�8O�8��y�!Og"��@4A�����GG��y�d�.V�=[C��;k���{�ŀ�y�J�/I�@7o��N��bp��5�yb��ZD�J��Q���Gɋ�yBk���e���]?@@�����y")W�*"�z��_1V������yb����z��@̈́�o����%��yR%��(��(�c��!y"��R��y���|E���ԛa����e���y�-��1x9qG��䠽��N8�y���)hT*Ö�s��Y����y�ʈ�ik�9Є-J>�8���8�yR���YO�`P�;:��{�%/�y����f��+8,z���s���y��ٓB�����W�$3�K�+��yB��n֕[Q��; ���1S�U�y���u`	yG
�=:4��̌w�<yW��	*�b������X:�'	p�<!�P)W\�@L�9k��m�d��n�<I$)��+	�y�߳? �XbVDd�<i��n��Y��-4��0G��Z�<i��� P��M�'�Ĵ>�z`(�i�V�<鴁ͨ|��Q:rj3
�� H�˗k�<i�� *<��p�T#;>&y#a[j�<��O68<��]u�d4�E@�<�B
]	k��`��,�3D�Uy '�~�<q1
�"*�� ��/$Y���o�<�d&�6:9z�f�]�q����r�O�<i�a�h��9��%Xb��(�.Xb�<G�;0�d%@��Π,z�q�Z�<���Q�}6܋$]�eP����fb�<�&��L�RB)�\� ��F�x�<���ZR嘽�T���uT��"��SL�<�p)�({V��	�$ �)�t��H�<���U�# R��'�8�\@MB�<��cL���$J��o���0��d�<�@���,��e�S�0�@���i�<1��M֨��  T:��*u�c�<A� ױi��H�#�K� �B�JIH�<�E`ѩR���U O7U�X͋A�p�<!r�Be�AP����̳�h�d�<iTFϨ5������-N�,��fD_�<q ���h��x��M%� )R��_�<i���?�=�r���{��H"N�r�<��e�"	�p��R��#Nr,д�n�<Ap�N�vXPܲbK�5H�Z�[2��m�<�� �X��Es��
'8����h�<Q����W��H���ц��df�<��I�vO�U!�-q6��Sa�^ܓ<nՅ�	_J�ha%�)�Z��g��H�B቏+��!�R�8-��ˤdH�"�R]
DoPH<�Mď^n�C ��fm�qR�Vp8����C�0�(��aUiB�x�� �Ȇȓ[6t�21��`���I�2b�ئO.-B�)3�)�ӑ6��Y���M�a"�C�J�15� B�IfGdhZ򉍰d����$�,v���TX����"�FW���@��s����3d }���*g�O1�>��� �
.]�0�Ս�Х�T��v�B�36������R��5�����OR��1��E��a���>� \�I۔B�$��c!͋y~4�!#�'��	q5�����$��w1�	Б�ߜ	zt��fL���?1�ǜg�!�u�߾D�^p��Oz�' z�{�� ����IH~�H"+�<;1OQ?cb�ڒ �r�<!����$	�c`չ� \ڒ��<�D�0~�V��t҅����v��,��G�+̦��Ӏ�4b��B�	�"H@XD�D�n�\�U�ȆZ~���']$� �
�M5�����O��d�y��YѴp�ԂЅ��?��KQ }���`5���Ղ��Di�Fc��:ԡ�,���I%N��?�~��GՖ�3u���!a���x�'f�9��,��c��q&?��b�@�'��ۄ
ZoH ��%���0��㉛s�N\�B�J�8ȸ���M�e5J6�éK�hY+��}5��S��V)wg�S<$����'^p��Q�V�m�2@ə�a�*3cSh	�|K��>j�E�RC S|�"��ǐ�M�C�ђH[z�A�.?��S�AQ6����={,�n�{����P��-r��Us&�@�H�|Rŉ(CUb!�gΏ�|�>"�ʌ U��N�N����X�0���S%$��u{7�H�sa�#K��Ë�~bbΕC�p���J�� o��(Ov�fj޵I`$�F�[0^���	$���TaI�:�M�ko�p�vA��tU���+ȔH1Va���פYIQiYx�'¦��)F?%d���dB�7ڑ�#lZ�Jb�QF��L�6EZt��~B�I��Mnڽdz	��Ze����lF3z��d+��ߨ�S�m��9	�~BM˓@�S��C!(/n��K̼
T�=�D����Gר�ӥ�їb���'��9��N�[��a�$u�F�(;O�a}�+@"6$HFh0^Eb�@pG�39D8��h�<R �	$7Tq9�G�(�F�"g�b�BtO�s�D9��`���$�&�������
���ãF�Ƒ��2��3VX���[%���U��>iQ�K�y�M1Q�P�h��ȳW؝6%8t����4S�����E �jU�;�R��ԠD�v1l�i�шx�����!�J�j�Ƹ<���@ɊFҰ�(X�L�cƬA�cS��(:g+_���aSe�Z�D��I!N�d��DʑtB����>\>�PAF>�Q���B	TL�n�;p��}�;-(.=�4��(����%�.t� h��	�2�4hCu��
yV�A׍�ii<�0��ĆR�8ORx�c�}�pX%��vh�P�&%��]�X��T⥟�c���Y6�5>6�[�n �v0n��E��%���Z�kÙh��� B���1��M�xaֽw�6m��`�F��!@/ ͸s�޴��x��F�-7���	ro"`���r�>р�_�;� 9���3x���C�Ɇ{�'<~ �#-H�Pø�� �� �h��0�x�_�/hl��u�V���Ô9@�����F�G���yʟ�H#ɗ	3 �N�7u�y��C9��*sGG�s��ͻzҐT{��4/�\C�D�qQ
�I,O��p�3��D+�.�dU !�I�h�N%X�Ğ4},����	
�(��)zX]��+R3l��PHe�	E���1l]�W�D�@¥�E��IR��PYC�dx�'^�q�n7��G�%����yO �eW�÷�='o�pQ���~*��pתH�z�fT ����aNf`�p"O$9���D�G�:|�.��t�b$�M�3Nx ��1o�J�&V¦#}�5O5�̈�qB ���!0���9�"O��acZ ��ҳ䁭w#`L(����������}��x3
֤B���d�UrY)�AZ�+)�Cw&�3M�|�͹$���bD���N�$�<��
�r�F| B�9�d�� D;`P��h�i��@��%ړVY�#��ITyJ��պ*0f1�C�JJ�<��\O�9����k����nC�<�	��H�Jd�֌\��L0�[�<9��
$�������� $�!�	o�<��۶Nj[��� ;�r�q!�kܓa1��DxJ~�V��f�&X�#gȼov��k�lYk�<)&��bj�1IP�W�[*D�⁊��O@Q��Y�(j�̎"Ut%KFGR�A($ D��`�흿�<��!#�1O� t�E꿟xd	?�	9j��#|���*JxJq�և^����b	�`����֬q�'�0�"*I�g�4ݨ�&\1)���'A�'�G70�a{R�V�,%��1�İq9�EB�'��b��Du�|7$|u���D,�U�H�i�K *-!��-9��kҎ�>p:��#�ʀ yz">�e 1��E6��]�R������jxR��6C�[�B��2;eV��a;I��|�c�2�\�	�
��i��t��+�4?mF<D��aQ,��B�Y2�h�BA�x�2y��I!�@�O� �nQ@��ap��;��m����M˃�3�0}X��)�f�3�r�-r�S�.VJ)Лmԡ�=ɔ��M}2�L>J�xy�(�|2���0<Y2m�"�R���g�i\�#sÑ!���k
�(�%ڐ��k�ֹ�!�K�B�P���O�|37�LeU�5r�&�,O
�8Tv]
T�]�pB�@��g_�~R���ȓC��11�m�c�x�T�C�2�"DxL<A�Y������B�6�2d� Qd����U#��ۓ-�=���$Yt�C���qpe��ېw����R�<Ɉy�?0�ܰF|bHMV"�YR&��j�2��a���0<Q��6	<t�<�� , b �V�<(�����O ��-��"`�����65|�`k�\3:`�J� '\OJdkƍ��d��|"le��)�?P�`Q���.6!�D��ƹ�w.�9�8("�]�O�hx�DE>�P�ȚXC���T�K�|� !�"D�h���Py�.\{�O�3l�1H��+D��:g	Nb�6�CҬ�D����CL(D�L����3o0��s �B9�@�LF�!�dړSu���i\|���G��Y!�(lÞ���"��&�����(�!�D��Vz��\<�ΰ��/Y�!�DM�� W��d(8����Ab��~��\
1fV-jP�[�m�)˖D��YĬ��4���(X��0����ȓf�Դ�EJYX��Cl�]�6���#r��"J)k�t�#�Ä�21�%��{��	mZvР(��; gȝ�	�'f6�S���x�� s+ŕq�H�@�'̒��MÜXe*P��K/2޸i�'-�Ep"���Z�����f)��lc�'_tk�VF:�S,�2�E��'Tl$Ъ�#�lZ��*,�{	�'����ƀ�'�(,�"��0�2�'~�:�JB=ba^��qΜ>.�d�!�'Q��Ö'\ Rl����̵�x"OP��g�A�|��0�o��m�"OJmz(�.`�N���43��<c�"O򔳒 �#��l[A��>ag0U��"O2��@�5��A�E]�^M҄+�"O� ���i㞡p��5��+5"O¹jTk��ľ���3e��w"Ot�����9ș�E��|X��q�<���E+$M2 ]R$�|�C�n�<a�cV�3hp9��5{�dbl�T�<I�ٙij|Ĩ���&���u��P�<9�M�I�0�ig��7�V,���N�<��e̥8�ta�/׬`#��R�oYH�<�gN�,�
1#WO�K��c���@�<y6��j�b��#/�(l�1�2a|�<�㧇3p��h�@�?ݼݘ%DRN�<��NU�V캝��d̋@�aDa�<A���(CK����(Q�!T�qh�]�<�U��>�����Z�[,l٧hV�<Q��7[`ٰ��Ʊ
�ty���X�<�4���]��㦘*"U>�!T�CP�<6��Zti��.�&Af\���J�<a�+;%vщ�灟GL�Ym�k�<AF�ڊ�R���y����f�<WHT�6�����
F���H#*J�<i��7�= a�@oM~�����^�<�UnA2Re�1�Dj�)�h9��LVa�<����|�Z��#��]��@�v�<�`�2�.�)���'W��,�tp�<qfMF�'���"�I�!"޹��'�k�<�U��6G�&�!�Y��<:M�k�<� ���b���o�� KC�8Z`�r"O�Т�O �`�ɋ��Z$
*���"O�Sr��0-Cl��⛂��9��"OL ȵ`�4��*#+%x�l@�c"O�m�w��=R�+ȈM��p�"O,�@FT8��\��C�V!Ne��"OU��^�fo�@ +)��X�"O��;T�^��d�ٸ-
�z�"Ob����� �w���dP�"OҐ��`��fre�@��Z�"}CP"O���f,�y��OT-x���q"OT5�`<=�F�k������"OP���k�: e+6�F6)��-��"OhK�ڀT>��7,�=qv"Ox(2������F�ți�	a3"O*0e.֚\�.l��
YyAƽ�"OR��Jư^���BUiU&$�Kb"Of��DDŋY� i�ĈN�;T8�t"Ox�:��0CW���g̅<�����"O:�����&��pq'�, �"��$"O�킠�O�M�Ԩ�p�4�v���*O:���>?���d N]
�S�'��	s n*,j��=L�Q��0D�8;�䅰6��e˕�<Ck�=�1-D��9s�QT�~�Y�'��a�ҁ?D�x�$V�����J�>:��
��=D��ɀg��^"irp�0x1҅9D�HZU,�Q�bXz��)E�����$D�X(��֬A߰�pҢ��������?D�h�0 �8����n�,����;D�hj�&�b�v��V�葂�"8D����́T� Q�Ƌ� Ԕ4�t# D�,�E߯������vB�k0D�t3�i��Y�0)�B��N�h���,D�|����
T�*,��j�)PTN�{#�(D�Rg�	�4<)$�әY����*D�$�6Iٶ$��	a� ��!�-D����-�+^@�'%��u���@3�*D�|�$�]	���`�_�2a,,D��s_�A���Ǫ�U��P�"0D�<2!����,+��C�)ܞ,8��3D��3��9b2>�fMC79L^|���/D�İ�K[m�B֤�3-7�H�.D�`���X:!|��B�^�O�CFG,D�D���K�׊��3.�@����.+D�lH�M��œ��\�0ھ$)r
*D�`�0B�:|�Ι��E�m�P��b(D�apgM* �!�7�Dajd��&D���%OԛE�h�3I�����m:D�L�UUlD�"��V[�.�r$�:D� y��]�4�gIV�';��b
+D�L�u�ڲ��n ��e��i'D������.Av-���#s�Ybt#%D�df�ߑJ���&=O��6$$D���wB�E4�h�q�-�d�bWh,D��ۀ�N����9  l�80(D��V��R�H�2��KV�H(AH D�4S���,;�~%t>�4z�')D�̠�i��j�q��k
=/�9B��1D�t�SiЎg��8p�F= 
���B1D����)�5`���xW���X�윓�:D�����8sp���'@��I1�Ix�E8D�X�֧U�[M@|�&��<�`3c7D��u�/~��h�%�	k��
6D�� ^]QL��_G�-P ���&Y�#"O
�H �Ԃ2Jx�+B/�7Y0 "1"Of�8 "�"P��=�S���'OF���"O�����<bV*�R��{B���"O�	�2'�oNn����{7�,Q"O���2K�W�P4	�d4%��"O��k�w�؄�"�Y�!*O�L��'�j��J!+�+D���J�'8f�C��C:-:���p+!<� }��'����weVO�,8�d��2���'r�#&�Q$m"�0�.��0v�����!<O$�5��4򎝺�JͧP�8�`7"Oz媂JN�=`@�Kb�)}?�5i�"Ob�
Q��x\�A�B ;Y>��@"O��H��XU���=H@*)b�"O��Y�g��
f9�k̐=$�:�"O�]x��Ǫ\�6X�C�ʷh�X�c�"O���a��:��V����@"Ox�p��E�S����HG�m�ԑ��"O2�����P�v��2J��U��"O�yh��JZ9�s6^2{���S'"O��!�a,!3��Pt� �"O6�(���!F	���<f�0/�ybA��`�P��<9ֺ�a"���yҦ �s���1IW�2����ޕ�yB�ʺ/LR�H"dܴx���Ub��y�M���k\�l�"�!+U��y��	!+3��Ӹ_1f��'�Ή�y2)�
�NH�3�Z�I�����%���yr���F���V��	���Z �yL�+�t���΍�r��i�e�%�y���[��Q-ԐQ�B��y� 
s;leC���  ՙ�y�OA����'�3lQɞ��yr�֜0xE��{%�p���y�Ԟ,�ڥ�Ȱ?�����C
�y"�"<,�͇9�� ��ٌ�x��'\RUmީR�r�҂�S�,�Ѹ
�'���8f��Ā���+4�h��'��d���z�H2@$�>2�H:�'����4�׎+�p8G��)N���'� 9cV����l{�W�����'".����$�fs#�ԫ] �#
�'ep-�&�G2�.R`(^�N�t��'b�B��Q������w
��
�'j���CǊشm��Ĝn��H
�'�,9ч��TdUx��"_
��'IH�!@��$��y��Q!F8>�#	�'+`pR�m�28�x����	I����'�<ػ��?9�TOύ(i{�'�E!���R��8˲f�F+"�`�'�`!��7XA���T��!C�)1�'��c�/If92��.[�JC䉰p�dlI��^��� @C8�*C��]��R��uM���˅!^��B�Ʌ!�v������S�^\K1��3�C����H�fܩj�f�٥J̯�%"OB��e�)_� ���/F��s�t8����I�>�b%Aa	
uzr���',D�X`�n�"qۂ	����5m�B�sc�)D��z���C8:E �@�N�8��Q'D��r@���s��e�F��L����8D�����
����]\��o8D��@ROQ�,���1`�I-nȉD7D�� bM�p��l���R�$1 �I��"O��g��r�P���MB��M0$"ODM"@A�I�\B�� 3A��J�"O�4������`����u|$a�"O
��g��#frlt�5�5AԲ��"O�b&�=9�\[���|��\�u"O����.�l�u.�>0�(�w"O�@b��� z^[�	�L�"�"O�U��-V��0z,�
�̻��'Y�OY
qB\#���ru�U
f�j�ࣞ|��'�ʀ@"��$�^�D��K�T�)�'Д4B�,�nr����Ie���'��|X���0£�޾){���'
��sW�-5e�I��M1���
�'c��A7�-�&�ΖU��
�'"RmQ� [�!�Z����2Ox��"�'��D�+�7Jx��4�,E� eP�'��4��O��)�*t����B��E��'f�����]	��#6��P��'��u"g+[�)�~�:N�((͎�{�')5��$��A׀=I�薷

Ze�
�'� <���3^\P$� �C
�� S�'��0Q��������8���{	�'�T�H�������߽F�:�Y	�' $9@�lE.��L;�$ɘ>1�5��' �k� �x�J��s
�%C�j�1
�'��$�fݩ!�(�s�03X��
�'���R$�/w^=z�/R�uz�԰���y����BM��7e�q���?�y�]4r�L�C�!nH�ձ�m���yҥ��j�bO�+7�,����Y�y"��9��Th��ǃ?� ��-Y �y��HFeRܢ�^75��XS�Ʒ�y��'a-8�Å%�]1�=�%ᝋ�y��A�9���,M�2庅��yB��"P�q��)>�f`�TOL��y�71ze��T hNl�s�ڣ�y���&�䪋�b9�-�s����y�(S�,%x���H/Z��c����y$B�G��h׌P&?ʌ�H8�yb'�'�����A4�乩���y�L��%��� (C�Vf��K�7�y�C��~�R董��UE� ��C;�y2i�5�:��0-ϱ83�q�ф��y�9Q�8l����-R>i��9�y��������!F"+�@�@0g��y� �:)����7f	{�T�D폘�y�Ժ<�5��F�*�Ag'�y��E4{�d�@�C�2~��rf�]��y�J5�P��۝*��=�%���y�ٹ[� P�LЙ/����
�y«C����!玥�\�1#���yr�W�e:������X:8��cˏ�yR�".s^���R$J�@��̽�y⚗i��lRFe F����Ҟ�y���#t�l�X�`�@�JU�G˛�y"�c|Z�9�
p���	���y�̔�ޘS�D���>1!v�O��y���$��r�OD�����HP:�yRAr��)W�Y%C,��!�!�yRL
�*��p�d-�Y�Y�M�y��	M��KS �'�f��s�ʼ�y��/6���$G�
��ʓ@�-�y2cؑ*;|E2�̕)�Hs�!ˋ�y
� (�8� �%Z" J6�خbdb)�"O�S0!P����U���&��7"O�%:&�:v-����<�X�@t"OL�u� .��I� `M����"O�d�V�W#E�BU���<v_1{�!�D�,.��1H!i\��Ɖ&!�D'X�p�04�\�KT͡A_5Tc!�d�0O`�
���D@^���鈔n3!��y@U	��ǵp)$�
GK�)�!��(�4�QP��R�8�`�6w!�$�y{
D��0{W�AL�A
"O� �$,��(�l8�qבdZ5��"OJuk�!-�ޡ�3��0M��r"O�<���X�G�X��#��h�ѫ�"O"��%c�6E"�M��b]6G�Bu� "O(`+A*a�ޕس�͂S�"5+�"O�\(�	"�XK0�A0��<K�"O����F�4Qi$%��G�5�j�cg"O~L�P.�6V�M9�-� (����"O*�Pr+�si"��Dl^��-[�"O� �vE�(��qX�JT�@e�"O�܈V�F�}�Vꁪ�68�1�B"O��z*�d�X)�%ɐ,/��1"Of���K�plV)J��Ӂn��X�Q"OjICvJH{:9	q�Ґt�F"O�P�T,Z�n�ܱ���2*�e��"O6�{�LK�.��p1ւN~����"OJ�!n��rzp��0�8�x�"O�y�D�]}���J,����r"O>�s�)� J�T�+�D�RuX�2@"O�I��AR�r���B�"�Eq ��"OЅ�F�U/JG*�9BF�cnFĚ�"OHU��̸P��Ze.��eE�d"OP¢�'b�Z� �/��?)��"O��䒵 ���e�	�x.� :"O�����y3N�y$A�~@1"O���QGC�uB���`Z/ �"c"O��r��Ѡ�fU�>-��W"O�y��
��(��e�r*��x"Oj��4�T��N�$:tQ "O@�C+еk�&qz�gRp�q("OtU��
�t5�2ǟPԡZ#"O~�����?��01��0�� �"O�i�-�g,�8��%X�W���"O\5��fܛ	9��8w$ )�;4"O�mٰ㒍Ժ�B���E��ٓ"OXi!ekS2�B$��
4�`�{	�'���Jddъ�J4:uY>cq6e��'���Rs����p��k%$ب�'�!�@�Ҳ��60k��
�'��*���hkX���(�(9�
�'#ؑ�0�B�����-�3*�E�	�'!`�$#ZH��1i@�˱"H~�y	�'� 1�I��;�H�T���`�s�'�V�:�"ւ{>����B�۠L+�'��9zr�
v(�����.����'ǔ%ڇn^F�H40��"r��'����-+-�n�&o���-��'��U�ʇ�h3�ÍO�%`0�'��ɲl�*D1�u3��	A*,��'�p���+�9JMd�sjR6PhL��'��LZ2 W�)#иC.Ήee��c�'���@���Tz�P�/J`~�pA�'|�ś`H3p�z�H1F7X����� Ҵ���ް��4�M�~ ��"O"��o�l�`M�r�[�튤�"Oz��@��2(��WD�<l@H���"O��gE�2���ڐ��f/�I)�"O��h��&�D��	?j9 �  "OL4X����S�d�C�OS��nl1p"O�1�dʋ?�5�F�c_�� W"OЂE��#�$A�mA=&�
8S�"O֝�bۨRx������kլU��"O���W�1��z@��M�v�(�"O�٫��]�=P@yR�N�o�B�S�"O�\�R��G��0�B�'��L!�"OmZaI��G8%qb�!���R5"O(T��@ɸ
�\}p��FSvR�W"O&���AŔ'2�-"3:<�:�"O�%Z��8��s�D�/�0U"O8�w�AFM���1�O	�Xs�"OJ J�#
�|Y�
rD�D
�p""OT� %�P�l�� ,D?�H�ʖ"O��S	*v#�l:udr�u��"OTx�Ç�O�
� ��7m�:I�1"O���R`A�D4��SriE�|����"O��I�ט���!f���u��"ODșN����h4%ʻ$ƦA�"O&|	F��%.�pRfc�'H�Y�"O�Y����3- P+a�[�h���"O�	YD�s��aܬO��	�"Oʵ3�LEz�d������lĘ@"O�Q�vF^0:v���@��;��@�"O�ġ��	;{=���/�1��P{�"Oڹ�AŢM�nM�P.[_x�;#"OZkC�E��h���~�=cB"OV,�j�
Dn����Ϸw�����"O�A�!E'Lx���Sk�&U���"O��Q�D�z���CЩ9�����"O��ڤk�}(P,�P�
�H��Mxa"O̙�E�ł�5�����A"O���ӗ;֬`l^|�6���"O\�f�,n�$qlۇj͂@Xp"O�`��BY�V�ԡh'� +, �xc"O�c�@]5R�&<Y5�\$5�"O��-e��2©��CIԼ!����yR�4Q�����$;PA�ʊ	�y�"S-h`�����{����)	�y� ��,�3�
�s��=ؗ�y".Q�U>Xi�(��r\̜!�DY��yb�A�}�ȭ�F�Y�W�>�ZW����y�m^3��ї�ү;��d̨�yB�E�VpR�(˝�F��u�S��y��VV�K�&�D�"l��➲�yRÃGJ�C`�*-���B� �yL�,��E������@�k3�"�yRH��3����N�Ez�Q�l�<�y���7�����#W+u)�����,�ya��z�K��U'HZ]+�(�y/R5w�e{ua��b��u�g���yҬE���Cp���A'o��y�\$��t��>i᠇L*�ybbM0dm���jLh׍F��y�
~�r(���;�� q�#�7�yR��z�.@i�����%86ꍔ�y�lK� \P��!�Zv�R�	�*�3�yb��JA�\��hӶo��%�&�U�yB�#R�Ci�ܸ��%Ϡ�y
� ��@�AZ�!��wC�2�@��6"Ol�:�הo���_%r����"O�q�#ǐX�t�81�ψK�^�xq"O4����,kw
�����F�b��"Ob�1 ��8��#�!�3���U"O�,�to�	>Y�Mx�IE�o��ͻs"O�$K�J�����"���ln0�Ks"O�ԋ�jP6�Ts�g�"E�f]�W"O��`�۷ �:I����c�^�B�"O*�ń��=Y(D�"�6g�Ld�"O^!��!��)b���z(3"O�;g'�j��"7�:~�@�4"O���*�!c��x�j�[�<h�"O�@�ˊ�glԒ��	���"OF�c��p�  ��HR�ny��3"O���.��!^҅���By0�J�"O��Ā� �l4
���M��(�"O:�rծ��sl�QҴ��|ļP"O:-��b̜C�<�U�E"OX��d�\�z����A�TΨ��$"O����q�|!� A���"O|qh3���F��$���G�u�=:W"O�t�$��/�Jp��hQ�h�`�5"O�ԚK�?L�-q�͝9&�� �"Oh��D�Y	�L1�����~�� "Or�i0�K�Vа�K�E3z�!��"O��8T������0ǅW��x��"OrAۃ�7)�D��KW�]ި1�w"OT���(�%�jH�wKc�nh1"OZ���.��b�1�,j��89�"O���I8;R���Ec��*����5"OR����68^��QB����I�"O�y��ĹDz��!"Y�Jq�I�"On� �'�@6v��S`��X>,��"O2���J�3�*��� �`W��"O"�r��>��Y�.&|W�M�"O5�
6T���/�&U�Y��"O���#���zDKЈR���e"O��Q�.U�C���i�H�v����"O�h��	�u�l�w���;�Ă�"OH,Ȓ��L�2�٧���&|�	�"O|bv��)�,���e�� �T"O@�9#E�x�x,������@�"O���deO�m`色��=� Tcb"Oڴ���9a�R�[Ў�L �	""O�ѻ�	
��4��M	:#���"O�e!$��rB���l5{��B"O��g	��G��k��۪DM���GW�������X)r��X`�%跏	�0B�B�:>V��;�.�m�,qꦡ91U�B��Qϫ�Ͱ$�d��o� 6j9
�'�hP�"��R�JI`u��8++���'�$XA��PhV�s���$�)��'� ��I�	P��J���P�''V��2�l"�1#�j��C�0�����d>��S�Ja�`1֏^�j�f&џ,�%�ȓp����-�W��M��͔�U��=�ȓ:��ؖj��4H�H��O28��WW*mA��<��8��]I(���5�[V�M�/2�ay�` ;��P�ȓm�̹cl_4r&��H�F{�����+-���[�"`D��]*�n��ȓK7<�e�F)`�n��F/��E�'�a~�m��z�l���Q�c�hp*AA���y
� 2X*���[���ڀ͕k���G"O�<��O��`n�p�k�9 0�""On	�IĹz�H�X�i¾&��!�R"Op������K���iG�O��^���"O��  ��!tp�r"C��8�.��"O�1�0�уC�,��3�
�/���b"O�� FH�^��#	2�[f"O
2��$&3P\8�c�;&�EV"O��w	2fB�<�6�%(l��W"Ou��*E-��9F�ٙAzy�"OZ6#Q2k� UB�m�
x���# �1D����H#<{fغC-��L,�|���2D�X� �E"?��e�X�zK��e��OLB��5{c2�10�Äsar)B�G�D�ȓ ��M�Q�ù:�� $:�!���� т��+!1��r��7 �ԅ�L���b��5��͈�솰�ȓV�\���[�G�Pd-ӸѲE��^x��FÝra�����D3]��<%��F{���C��s��My���j$��@���hOx��D�o��d!b�oU �j��N]&!�@�Y���T�	�_`�B ��B�O��=���%���>#NH�毜���yR�N56�����;,�8BrG[�y"�.�@\ ���r�~��v���y@ul�2�.��@��&�F��y�C�&"#X��g&ÙM���dS�?��r�'
ԸDl�D�����j_8T5�E�'���qc-U�F��˧n��`�$�Y���$�'��h� E!��ģ�	��qԠ��ȓAݺmX�Z�YBh���T��4H�ȓE/F0KS#ڡW�+q��M��Ąȓ<��m�����F뮴"5i%U����p��fbA�/d��"Ѐu�ԇ�5E8��2e��+��i^9\� �����`j�%a�� �oU�J:8�'��'��O��.�x�ꑀ��	�����G�F�� {	�hR�4~�j3��.�� �ȓ	��,˔'�
�B	��#d���ȓ�Dy�g�_�4'���6?��!�ȓ_��%@Ŗs%����uڰ��' a~���F�đ�e�J6Y��͢#i[�y��=/�`��W4'ވSD�	���$ �O�	��N�c��h{C�G ����y2����9G鞱o�hq�@�*�y"-K���yѫ.9�L�`g����y2�޼+����mG�,�0��IĀ�yrȖ�9Pxi�t
3�lq��y2�J���X4�"�>�j7�ĭ�y�A�H�4xb��'��ad�X��'�ў�O~�@��,�P���q��;?=��Z��xRK��g�le�S�ɳq��
�I��y�M�'
�%�q� & �6����0�yR�
��bgڞu����c[��y�*ֵk2�S���7V�����Ҝ�y"eOl�4�KG F���*��y�h,��j5��0SԞ\�!X�y2�C�Iuf�q�J�@\�`솎�yb��"�)A	$0�I��$���y��[�g��0�oS�*�
������yBaw[Z���g�
�����&$�y�f��O.,m�5�˛F�`]0R����y�N?P&X����[*>�|!"I��y�Q�`���Gf�7.z�#���䓪hO�b�� ���p� >�>i���Eo-J��@"Onib�ߓq �X{��[{Z1��"O0�`'KN:��5�ѽʬ9y"O:Р��(��ZA�;fƨ��"Of�� �V�A��� �P�Ayd"Oԁ'	��g�F�C��4����"O���E�G�c��M#�4��M8�"O��T�ΙL��آp�G9Y0�1q�"O�p`�Y#Ldbb�إk�p4zF"O~M�Q�|������):p�t"O�����:u8QG�	�-�^!��"O�S`��T���ӌ��D{Lx�"O|!і�Ž1�lQpc�\�;�r0�q"O��svM�rnt}�w�Ph�&�! �'�1O|� ���$s�d�K���>{T��"O
�Q��ܡ5sH��,U�:��m"O@�G$�� XS@��P�N�q"OL�� ��x��p�F���	jP}(�"Oؠ��
�5~��5XDL�8Y�#'"O���W�L8%��y��%�4:�* �"OP����&�x;�6~X��2"O�9(�%�)A�RD��t�8s"Oj����Y��� �F�/<v��"O�������S�K�i��`��"O�� CN@���&m�TF�ԱF"O�ؓE���:Lz�XP�ġA�d ��(LOR�T`��%���VVv�B���)�Ia�'9!6|���v��zr��0��%��G{����N�+�jpfX�b�Q�S1�yb
<jX�J@
'�,�怔�y�`M X�Ps�@NP�mj�ϓ��ybY*y2fI!�F��.`��N�"�y"�`{��
`1�u��	�\p��
��҉5KK��
dҖ,ijh���a�lnx3g�sw�0�Qe"Ņȓ�<���j�m�T�{u�@	�t��:�=���0{�u��@�o�����҇AH�Y�}*� ւ>�f�Å-D�P+�	ߦ[ ��N�$>y�3.+D�pq6(�"+�"�p���H��a��.D�p�G�>F�T��ׯ\��5�*D���t'�(l-���WE",�P�)D�<W憷{N�=��JN0Q��	�)D���1��xb�1��0��� (D��C����oн��f�4F<!
f�1D�HhCY�L��;���[p8�60D�2�Lۃuh��;�a�/�Hð`"D���mW�o�r%�`N�e�&��`$"D�<�e��+`-�"F��1����,D�Pp���t1������*����p�+D�Lk�l��~  ��8f0��#t+D�ؠg�� _��]�6
Z��p��3D�0 �mٍ<�"�&Q�Hm i7D�L	�̞Y��@�� ܶ��7D��Ȁ�]�͒��"("J�! b5D�0҄��3;�P�ʢ��.4/�Mr�b.D����=�x7�@�嫗�-D�VQ�n����!��)��x�Ǐ��y�*��.����[� L Y����2�y���L��ըb,N�
 ����E��y��&6���c��~�����ӳ�yBh
�31Ġ�Ƨ��-p öK���yrb�2H���»w��,ږ���y�N %���ƃH"4���uș��y
� ���d�E�n���q�b�D��y�"OBqX�K� &����5j�j�"O����G�o
�ix��Z ���"O*���Haێ�h��D�G"O�A	�@D6|z@	���ǲ
���"Ox�P���l��@H��Q)iR "Ox�1���JT�� �"O0H���%=���G⇌G�<U��"O�"g�M;Lp�y��īz��j�"O�����l|n頓 ��uА�:�"O�����n����
$a� x#�"O��@�ߍp�z�Z�-�ɰy�"O���B��/F8�:&���c"OL}�p��o�B�H`��z�d�3 "O>̰��� *���}$��z�"O��S�K,.�84�J��I(`9S"OPe�夓�;~���Vi��(V�K�"O8�4�ǆ��p��G��:>m�e"O�T	+ ����v�ɽ6��I��"O�9���0[����� ��z�����"Oڅ��W6$�.�#��/l<�[C"O� Ґ�ˤy��#���(#�x	�"O�t+��V�mw�h#O&z�T�`s"Ohbv��%�䡑��O':� D"O0����B�.%��2J�+J�H@�"O�@36�׍c)���)�$r�,x�"O����M<m¦( �-��lU���"O��E�Z��H��Űk@P8��"O.��(p�t!y�D7�,�:&"O�9�����qh8	UᏖ��Y�'"Oa���=x"J{6B/i
 ˧"O(�k2�:Q��=	D��pS�"O����D�Vr�!�"aF6]CF�*2"O�� `���T�uˠO,�*"O�,�z��H�@&�heB�"O('KE9��hI�V�NmP"OdL	�f �[������Ţ���"O����.<&�f��iOp�v"O��AǨIC%6�1g\98H�2"OX����г)�0�Dc 1+�v�1"O$��`ė&x��0*^P��#�"O����N�'?����O�
�)x"Ol��t� _8r! @�_8;�dJf"O�-۴ �T��\��ԣ
� � ��'�1O�d�H�����TE�و�"O�	#u	Ź)����B�Ʊ����"O���b���D�2�EN�'����"O�D�1�F6e���Xgm�<O}��ZA"Ou1e�"7�����ǀK���p�"O����F�Z�b�b��u�P�K`"O�y۶)�:Q~�q��%��0E"OV�c �ţaq��c�
f���q"OF`ʵbW�M�H�Ī�>p=`�*"O��G��$k��������#"O"�%� �ZH�� A���
&"O���&˂~�����탶"O}b�'5�@P%�A�k�ҐP"O�i�"�_,<*���@��rQ���'O1OZK�B+G�؋�+U�bD	�"O>��$���0��YBr��6\��0""O��	��B|Jl�����D?|�87"O�@;�b���x��n�6Yp�4"OP�*� ��l�:A
 �@�77vha�"O����gLD���':-X�z�"O� ���+�<C|ސ�S��t��"OJ�@"Q�*����� f�[e�d$�S�IG�	a�Axp�U7~٨T�9u�!�dס�ٹ�NR�H���CBG^�|�!���u�� �/�9^h�=�6&��M�!�dX�z�����S;g�e�"C66�!򤃬�|}h�dӮWJ�`R`[34�!�$��	c�����[�$F�� �t!�DVr a��J�!sL�h>[)ў���I�pȴ$�Pf�`i�X�PlP�B�ɛ2�@=��
$J-68���%2��C�I�5�)� �`�(@AF�ܠ-ڐC�IXB>�DK2� ��4l܃�>B�ɍ�ru��4,<�f�+�B�	�H�3T����&)��#Q�q~�C�5�&�{ŉ�6(H����@S�Q��C�ɟP�L0����s��� ��>r �C䉤aH�z��Y�H���+x?�C�	�_7���b�����#'�0�~C��:T:�!5I�w�88P�>�DC�I,B'x��X�@s�r�ͅ	]�C�I�[$8r��0q���b��������<?�w���+2l�C�����1Hi�'�axrOF<kn< �aE���X����y"˙4%iL}�q
�[�b ��L�$�y�JS={�r�@5��WhU	ԇ
-�yI��j�-��� :͖�p����yR�T�L��"�oõff@1ڵb���y%��|�`��e
�J���"�(F��y�΃�~��b#�$1 �kc��y���|��l)�C�z�D�#o�7�yE�1f�$�/A�z�(�f���y�.��gbns�&�Y[��Z*�y���A7��:ŅE���s�N���yr�ݜbt���'�'\�kt���y2T�K���5���x5�ֆB�y�n��v���4�
��L@�n�<�y���GLj�*Qk��Dz!Ȥ�ۛ�Pyr@�&�A $�����aYY�<i��)-uF���My�
L�P�ZP�<�A.	�9K��pS/���.����h�<Q
6Z�]s5�ۚ,�9 ��f�<Ү�Q�<�`���o��g�^�<�ΟUd�A袩_rb�1$��W�<��<�6%��*���h����J�<)�h�78|�����
x9F�b�~�<y�.	[~�;��	�:e1��wx�Gx��5 h���	̟+۶0����y�	�)B�����9*zv!���#�y�/ �@� ��d�ű�ڤ�����y�F	c�ڝ�E��D0#D���y2D�ܠ�Zw�ֱJN�)��NM7�y�-��h3B�&+���F#�ybl��T�y{P݀S֔�c��ۇ�y" I4�x�!��"F�B]�$Ɛ���:�O��r�����(�$-ʡ_+B�{�"O&����5GE�aB@�/s{�z�"O̴�e�	�i�jH�F��/i�PA"Op�� �֬� O�q^0,������pF�d�
4]�V��ԨDq*��ò�P6�y2AD�MP� "�9 ��a������=ъy�`�ev���"��؍HF���y�O�8,!S C��,�<��3�A��y���		��葈Mu�̡A����y
� ��)��MO�!�Ċ�2L�p�7O���Cɘ;T�<K��Q�y�0�!0D��32�*gbxh $\�r{p̲�C�<)OL�=��l@�C�iz��P'��g���
�"O�x{_d�й�4��%����v"OLq
�+�/z�T���D�(aq^�E"OFi��)�y[���dʐ:ю���"O�h�@���00��F�vf ��"OQ0�'k��)�aPkH�R�"O���/k��`�w ؍ۦKa�'�'�azB�ճ9PbY�����:X�r'͞��'Vў�S�<�􈒵An�40�O�jHy� \W�<���Nz:n�`KC	zV�x�Z�<��O�/��S��Ƃ2�#&��Y�<�D��G!H�+�mϰu�j� ���T�I� ��Z�s�"<`��F	Lx6e3D�@��`�����Ҙ@�D���OOF�S�g��Ĺi�E��#�K|*Y*t�A�\ў��	�@�\� �'����X*A�^3E�N�O���D#,�pqb�ӻGV�ՊW�T6�!�K�-���`��W�.�ͰÌTz�!�D��hD����#�&�����G�|��'��u��~l+u�4��x6���׍��yR�T
5��,2� ��ZOpiJg$�#�y�� Jّ���T�F�����.�y2��(,�N<�bhѸQ��9�#��y�H;�T��E%��Gx(��I��y�Sm��jwL��?/�LH�Ю�y��T��T�Xs
>s��CN}�<�aX	Q/~�˒�N�`SNd��`\r�<�'��.r���Xuꑕc�V��5Ėǟ܇��*���ҭ�gz��"�֔'�<��ɆW��Y��OW"v*RH�A�*h�C�)��Y���_A��l��B��bGN��%��;S�œW��Z�B�	���LR�R+����)� 
�0C�	�yU(p��c͖bK�ɣ�f�H}���(�-LOV1��W+i�x!��R�x^����'^ў"~���,��P##���)�'���yR 
�3��;�É?U�ڵ+W����y�� u�E��&ךS�v�Q%���yBH� `Y1V�I-Qm0mZ� �y�OKt""�A��veTX�ď�B�	�H>�x���u��Z#C��"�=1/O~#<�1����Mr���:f�ҡn�D�@y2�,&
R�Lh PM�X�`=D��`7��@ʜ�ɣ��Xx$�PG=D��9h�)'d�L;�	9/����-&D���%N�K�����A�Y��2�/D���)�AP�u�@�R�i�6k/D��Ӭ�0De�w��ab�=�c�'���1?�L��@� (PgP);���+Kr1�?).O"~ڗ�i�=K�aU�BW�#��W	b�!�D�x��Bc͎<{/"D�QIA0/�!�D�3Q�bAjbBZL�`����+�!��D*�ve��	�L�<y�f�4�!�=Ny���Gŏ�z ��↙��!��n0����]#r�D��D��4�!�D7X8�`&N�:����D��{r�$ˉ>����1��"
qC�P����)�'|&�͚��N�W���A��#}`v�z,O���D�uq�� W�6*������U�s�!�dʥu<B!a�%��,��y0�M&>R!�J�W �,��.��U��=A�}b��� ژh�牻mĐKЎ�i�^��	O��ү�T�|ͪ 	ϣ
��i�f%D��)�FH�\2T��%^A �$D���� O����2$h sTc#D���F��p������w�6�)`�5D�$�E@�%�,	���P�)��8�h5|Oc���	�"7|���Q�/����c�6�O��&\C`�cQ�M)B ��YjW�a@x�d!�����y��4<�V@kU�P$�δ��F��'R�?�J�!Jb��X��*�! n�%CL1D�D��SqW��s�	�R4�q�H-D�X:�Ks�Fi�p/##O$����0D�8ٖ#��IpJH:�F��!�<=�G.4D��`L�$}���Z��	��`,D�\�R�Ö>\^�!6iȫh.��&�$�	ܟ0��I)�u��JÇ��8ri��u8�B�%\�8Ջ�R�K��i��_�t�4�d�O̓O�}��C���im�%7G�Y�HV�J�����e����*<9XQ4���3��e��%���q`±gvĽk��A6\���ȓ �z�Z�MY"�l���#�l�ȓoF)��Љ6��$��F�w��E��(@�WhU.,(��
�v!*�Ȍ��=O(TK��(��y9�K��*��� P�&��E��'O��)�ϕ�0��1 3R˼��
�'�l��V�o���S��fI��"OpX�â��t�n�r0�*GmRA8`"O 1�%)��w�m1e`Q%Z�@"Oe��K�4rHy2���64%����'\���ec�pY���X��ت����џ�E�T�?���Ӗ�
�9piy�?�������@7��N��qӣ�d�ʀh�m!D���D
h�P�(ЉΝ.(�|� �$D���FI�q�>�KWe�L�dT[�!$|O���.?qG��?��q�T6\�n-��ǚD�<�!�
Z|�#vC��DZ��d�T�����|*����ٗ3�,�X%����F{��'�|K��2����-��D�DJ�'۞����ݛI�0ؕ���
q�$��'�дZ&�EX~�X�G'��!	�'��Dp�	W�bQ�(,ߧ۴X���=���kR
��2�R�P�cA�*��B�ɬE)��`ыǆ4R��EE@u�4B�I�\vA�0��:J\��"!ݡAx�C�	�M��=['��L'�;R \�-B|B�	�^Ix�`ΓJTZP��+�lB�	�^qP���N :@���X��rB�ɴM��}�F��)��ТehA3nB�	9@K���B+ƾvڜ�hn�<�.B䉮4�<�S��˻Bx�Ӈ�J��d&�L�B�� ��=b4�O���G?D�����Ri<�+���81x�k�J:D��Yg���E'V1B�� h4�����7D�,��D�,���ӏ&p��⶧5D�p���l�F`��@N�l@��:@)'D� jue��qn�<��K<����I%D�` �٨/?�J���?;6�؂f?�IS���qb�� Ģ�����k�<0`W�=D�X趉Y�.p
�kТU�o��-I��!D�,� ���j�jp��5j�Ω��(+D����ϛ{�p��D�"/�5�%�*D����ȟ,>n�Q*�Bj6����&D�H����<���K3n�p�Ivk)D��!��v�8X�P�J>xqfl���'��H���3� ���3��NSpQ��d�������"OJ��@��,W� -s�IY$(x�C"O���C�k����(O?Qe � W"Oz��)YB�H�&��PR���"O4�@g-��ad��:�);&"Ox�`#�S�XJe+��C<Y7\��Q"Oh0�-ȵBFP2w/ؒp!��'�|�'F2�ᄁ���ܼ �m�	����'��4P�e�v��1��o؁ymR���'8����%�f 0'�tٞ,�'��hP�+�Dx�e��X}u
�'�A�"��^��i�E-�?aq�	�'g���P��Pd/&G���/Od��0����$-����G&��`��8����[��O���$�(V4|��g�Ƚ!���҅t�!�$�S���+\rT�Js����!��KP��5!�ʭD"	K!��׫zR!�f'�U�I{�`�E7!�Ask]� ���z9ʓ`Ҝ.!��
-�pأD�N�y��D�f/K<��y��I\, �oǜkt\������C�I��"�K��1�� dh�j`vC�I�f���U�N>��rAS7?�PC�	�Z��AJ$�:`��x�bIϦq�.C�I?wѠ�H�O*��RA��*B�.C䉌8�qv�M�g�@��I��<W����h��)�'�"U;-���G�\f���wM�O��=�O1O��#���M�� S�;Ru�"O�}X�I9b�IpAM��5�ܐ:�"O"�Z:�A)��V�rP~��w"O����C�	�y��
�;V� "O�,��k�
�:�i��#Zt���"O�T��O/ 2#�Ϸ1V�ݺ"OL�dBɨx7�i9�n��mB���'�n��pȗ	i-!#�f��������xR���P�@��შ8����t�R�y����tH�֌+�J�c���/�y��)Wd`YefR�(���"��B>�y"�F�9�I��#Y$O�8G�E�y������ή[g����A�&�y�l�F������K���u�����0>9r�H��d�� �&9��L�q%�I�<���*�̡��F&�۲���F�<i�@S�H�6Ղ�F)Ed Â�B]�<٥�")rMXW�:�l�J�/
O�<y���z�٢��ޠ%$p�Z&��B�<a'��18d��/�B ���� �u�<	���e�&� �:&�hQҔ�s�<,��O�@)�ē Ī��%d�s�<�tmȈX��P�� &38<���s�<���	
 �,��7igʰs�N�F�<���o��"cB� �ba����A�<)c�T>uU��t�ϻ��1�
_U�<YO�W���IS�8�����%�M�<!`a`�f��`D� Os��:��DJ�<y�LS7[��YY�\ �b��G'�]�<Y�)��	��)�t�m?~i��r�<�2�R�"Z0��%�<Ġelk�<Y��|,\E"����� �g�<���2in��"�bY=x�ʼ�BEJ�<�à�<��8���[:W� T����\�<1��N?
��1x� Ơ�X<�CU�<if����9��F(� � �K�<��,��Z���hbMp~0��n�<� �,�#�#]�J|ia� ���@�"O�M3b�_�bӖHr�eP7(m���"O��;��]�u� ��Ï ���"Ot逄��*(7��K������"O�� �D�$,
�Ó�ފM��)�U�'R�	L�)�=�s���`O��� 
��R,JM �J r�<�ǈ3Vt�ѓ ��\+�ͫe�j�<���P� ���w�B����Yn�<�̕_�5���ǌL@�2�GT�<A���]�r�� ��<�@�2��P�<���D�lX��O�[`�ʶ��P�<!fǃ�F�4!��H�D����I�<)��l����dET�:,��	�O�i�<9͊�.����"[� UpW
�^�<��M�I����$�#�|12��E�<�t���=T����kH�V}�4��AA�<�����f�^����%1�8�����v�<���W�OL�lR�e��|��P��AWk���ϓ�>�r�hW1[`z��Z�ZG���a�,�J���O�:Qz�I�9E%�ȓA*��{�\9"T�u�Tǌ�\��9�ȓ �
I��c�q��RSd�
���A~�ԩ�'I�-���7kAL �ȓe~i���)Rd����[V�@\��ÀLçoE�S�P��G9ๆ�О�;2d��U=H�!Ljl~@�ȓn���!��N'K�L:椝�K�ꨅȓH.�y���@w<�1cQ4��8��Z����R�O%n�tمƚ+�����:�df�Q#|<�-Ad�J3O�v]�ȓQ$�36�Ҧ"T���2E�)[��5��RW�ȡ���d�l�8�_�dsm���{JZ�4L���7�l�ȡ��~V~�9�J��C/&������{:�t��#�Q�jQ?W`)�0�]}�Έ���D����NS��CS�E�[����N~�uCf"	!䜁�2�2D\���BMْ��W�cwnԪ_��ȓ3U����Hˌ~�8�V�A�|@4�� �>�ѢO�
ZЊ��N��g�J��,W
<1W˛N�=w`D�� ��˞Q���ڃR]��*���L欵��J�Ȣ C�#Pe��2�-V� ����ȓN-I&�E�J�&�R5��8���M�&�ʷ.��y�3�N��}�ȓA ���ә-p���H,6��c!ʱ��g�7'$��F�fR���h5 ��B/B�1xq�F'�,��b��|��%�:9���3��� i�hY�ȓ%��3�Ǜ6�H<(Smؖ{�*,�ȓz�Ƞ��.Ɍ48x!f�َ|�ԇȓ]1�U��U����	�<L��j��<����9H8���R?;.��ȓi^��#�O�<8að͂�`e($��Dg:������j�Q<@:�8���*MРV7A�L�K-J�84��w`� �f��x����T��p���ȓI����׼+����s��Th���*��I�q#U�LTǬ+��ȓB�fM�4-^�pVf��leQ��6}�1��'He< � �՞`��h�ȓfp�ؤC���0���`X�1�ȓp0��"
��v�DB�DT�Q��n�|QV�M�P�Q�Oߕ{D���S�? �x����6�d��$��[$�X��"O\Ғ�T(@����ᤗ�H���"O��IF��}�����:|Ԍq�"Oy��*�Ul�$�B�}Ќ!K�"O����ˋ����['��MVƔ;�"O� p딃)�N`�B��_,҅��"O.��#,��P	,B�"!��x=!�d����ǉ'\����#ω�B�!��.+2�i���ޙz�h�2&G�25!����T�`���! ��+J!�D��;�l�P �'PL ��	57�!�$K �|YꝹ>���BOʕl�!���[I"=)�	�(X.��Gd]��!� bh�ʑ�6Q�r���C�!�!����1P��=�؅�c�Y��!�D�J��A��"W�(�`�Mn�!�ٮ���R;��� ց�w�!�$Ͳid"u(�1{�b�����;�!�$N:H��/E:k�x�# Y��!��گK�ɑ�LЛ��<�eܗ&�!��p1��He* ���ksL �$!�䟛b�VhZ���z������)8!��Q5ex��F*W�"ߴT���Py�l�}���Ӛi��[R��9�y��9�>\{�`� 
ͼK�G��y��W�r��Q���"�`���
�y�+^a�ݠ�,��+٫�y2
�(s*��t]�G�T��ώ��y����p�I��P�E�����6�yR�L�{�a��`A�B�zYk�����y��Y�IVH8%�'J�TQ(��1�y"�M4R�6����n����K)�y�ȑ )-����#>����܁�y�LJ4>,�ѫ1��:�JY�#/*�yr��&I�^$�R��!};j�(fn���y�ʅ8ec��p��I~R~��`A��y�.@�>,��Ke�כ+Ê�X�K�yʑ����f
��J�\x�Ɉ��yr $��0���٣{`�� ݠ�y���1\#xh�
���2�9���y���6Y�~���L����[�y�A��`����50�x�` ��y"�;
Z��PB :)t 9Pd���y�fMxL�yb�R�2><�g�Y��yR��8y�|5�
���P(u�Z���'0�!��=V�����6�1��'���ɧ��9b�He+��*@+f( 
�'p6({6΂���I ����x	�'���&j�M�T�GǑyr<���',���&$f��@���*h�а��'�b�Q�C��X-��"�
`N��'��%x�AO� Q,���e�1��Pi�'΢�+F"�9|�z��A�P`er�' ��Ē=P2رq�*+)�E��'h~���+��QÖX�-��V&a9
�'��ŘS�]-XJ��
���C��	�'�b-#ӈT���I�I}V��'J���*�T^���J$D
���ȓJ�0�c��xΨ16�A�&@��;5�x!�f��[����G%kye�����ڼe�U:�d-����
�'��{W��7OB�0gƛ��X�
�'���a
��zH�N�v����
�'����fC�~�'@v������� @��#/�4l� 3�K:yb�"O��r�B[�b�$�8�&�+
1���a"O�(�T
��<�@����w*l��"Ov��!�j~4���Aז;s��"O���dg�$D��-)b᝺9�&�ʅ"O��Sg�����:2La����yB�ԌB�
lb�&>r?���'>�y",��O �x���,Rr�A��yb�&2N��B,��Wznd����yR��{o�U�5
�=��I�Q��ybOðzAx$C֣��(�b�@P�Ǉ�yҤ&H^�5�Q�Qb�ɲ���+�y� <-h@��QC�X��I�+�y�ȇ6Rn|�㮓�9)Н+A�N'�y� -3o:PsskX�7)�xj @��y��ļ?��1�5��7�$��'�%�y�H�}�V,�r��0�ug� ��y2�P�@���԰Tq��폺�y�Z?C�4割`�^B���Ҧ�y��P�&��7��jK��jE*��y��Ťu����u%Y \2D ��(�yb,��/��p�@/��P���5���yr.B�ǔ!���O>IA`L�K��y�G��I~]�֫�:K�$�(��y"B�{x¬����} ��4@��yRϗ%�Ba��O rN]a��ً�y�g
rOn����Е0��4+Do���y���P�m0р�.�4��@hA��y��4{x�(�	+��R`e�
�Py��K�T�`�E� �8��A�<ل���w0�MK�Ɓ�?�qӣCt�<�(z"ٸD[ PJ�(7ńs�<�1�\92,���I�o�Fq�6N�m�<��������W�ѵ'c��J�!�f�<y&S3A{:��E�8rrX��3je�<1Μ�(��)"q�P
WP��7�a�<A�4���Bc�d�4�Ue�q�<�4�I.�N����R�/ih�B�ɦ��	{�#B�m��'+�B�I%�Ԉ(�	��>LUq��^7&T�B�	�k�`=����"���w�_�1��B�Inv�i�G �:,�p�Y�Q.fo�B�	��X���?�L�yu)L@<\C��q�~��0L,G�8=�ԉ_k(C�I�d�� 8��"	B�x(c��&3�B�I�WR��D�Z(V%����ȑ"t�B䉷r��ŸD,I��p\�Ak$�C䉵tY�P�tÄtX,]�c*.`��C�ɦ:�.�ɠ�/��J�� &ҼC�I�9z`���E5uM<Ep�-�+8��C�I���Y2>$0�TE�AC�I=�4���W�Y�jȱ����C�	�Gv��c�B�;�NܓQH��'�&B�I4?�ZaFAq"2�qC�29�<B�	V� )�G�܁ClsFܪmB�I �p�B��c9,̨���I^�B䉎u�����)�p�C�J�t�bC�I��8�B6g�?���QD�����C��:�.�:�,�b�2�P�,�|+�B�	�n�\��0��B��<�'�/$�B�I�;��qP�&t&�A�Ab��c�B�-_�:�i&EU�O�fE( �C�;JB䉆>��-�Q��:�l�W/B
-*B�* �:���7��å�\�TC�)� ��0v)��ȵbV�.��́u"O�YSG��=|Ep@+J-\�f�[Of�nZ�q}&�*`�W�*j)�"�B��#{z��rD��P�.D�ǋS�:�"��$�E�'wLy�ҍҲa��qp�ϤF*��'�T�hWF�$&���rT.b�Ekܢ�ē�hO���-�l�#a1~��Qn �;y�4�"O0+���%o�>������B�ܽ('��7lO�yPǕWiT�eL)'��pr�O�$�֙O�u�P��\�>��4l�J�<���;�����g��:1�'lF�<�H�
���H�H�dY�<A���L�<Yf,DR�|42c�רxN����LO�<� A�p0���#=<Vi35��J�<1�dT�01f��c���|��#a�<	1EM|��$,^/�	��`_�<���9��Ͳǂb!;�j ��yR�Ӛh����*S�B蔬R` ؜A�
B�IR	fI�fm\�<��%�׮J���Ir�����1Sd]�;l�0šڷR���"O ���C�q!�
�a�Z��QX�����'A�`*�%��|�upE�
L#ne���)�'���n��y��lQy����BhF�8b!���"A��M�cB�gf���&�a0	��?��m$z��W�M*[�赳UKu��8�ȓ=�z�H��F0�R�jG���=b��ȓ^o$ ����!q XD`�#��-��	qyB�r����&%��}z�(p�M2�yC;n��0a�,����E
�yb�>��'l�?�z�o�.�Y(�z7�4a'i0D�� 7��)��S���*G���r��V�����D��X�ƅA⭚� �v� � d�!��X��li{��M<~��)+A��"�!�Դ{����mK�A�p%3�[3N�!�ɺc����&bˌ'������>�!�D�/WV�B�*\�T�p3�!�� !gl��7J�����cΘ'1k!�D̑V@F$x�%m�CU!�$AE�J��ʏo�ޑ2aL��!��U�*U5X7ÝV��m���[8N��;�O\x��̎�`cՌCIQ4EF"O�A2G�@L���(,ٲ9��K�"O�d�w,[6{U�J΄I��T��O�6-?�S��>Atl ?|���g�P��R�ߙi�!��c��`�g��(8@1�3�ŗ1�!�ż?���ʚ 4���熛=�!�d�8�J8����{�h��KB3v�1Oң=�|���5)�x3)њq�����w�<�%ŏwDJ��S�R��s��j�'�yB)^�4H�˰��'����
L��0>�J>�����R,iZSa�H���w�<��G�5Ye\�p�kщ
��A �M�t?�1�)����,�	iׄc� �T�t@��'����z��A����6�C����]�.��hO>��$�̑#��u;Ԉ�~� H�t+2ғ�hO�S�fN��D.�-7-A#�A�c��r�'H�6��x����� C�&@@{k�6m0��O �)�C��� ���4��eQS h��'m�������qp��@cn��<+����hO?�������e]`�\�d�ٖ�!򄃗p�p�pQ솲OP��c(,$!�$Ԧ9�8�� �xH��N)z!�$ճ_pir�ߜ�{l�C�!�d9��@�F��_$��hP	J�!�� ��05ɃbΊ�!eo�U�@X�"O�-��]�+B�M�cm�,�j��q�'�1O"� E���U�E�ȑO�f����'S��X2���4)j��D�$>�2�Z�L?D� �h����5YQ�[:Y]���0D��d��2?֒h8'�V�Dg2��f)�0o�B�����Ǌ+"\T�q��5rt�ĥ�<���<-��9����Nci �.E.^B���^����#P�8�XRE-,�0B�ɠ��m(�O��"4��){�C�I�� e��+)	���6���j�z�$=�P�&]	rt�Y�f��J� �z�N$D�D���ku�Q �I.�=��&$�8�Ԡ�5��x0䌚�Xۥ��yR��2vF��%����u�5l��<����"/�[�n��?#�� ��Ցp�� a�������Y� ��u'��v�NQ0T-���y�O �6�k@醽B{L�Tb(�y��K�'��q����5�RhI4��y�_���k��>A�9�t�V���IhX�L�t���1M��I�m�-����O��=�O���>��� ���Ӳ��'^%tpӇs��D�'���s$Dj����[u�0%��'(�O�?�gM��yY�M"��#f�~�{�
{�'�?�nZ��T���)y��X���ނj�
�'�a}���C��06�І)|`�`�y�^)_��5�5�B,$6�j�Eǝ�?��'9����l��>:�t��K�7N�]x�{��Iv�KG$��֊ŧ%�꽐���#6�4�ȓt����C�tPn���#$] ��?i���~� �|!�͉�,����q�<!�HذTf�0r�%�D��Dj#�b�<�g�,/�ڔ���49�f�8fL@Y�<9��hO����IʆJ���q�<���ESR�����ךO���k��p�<Q�O�����=k�α�Um�<9�Up��h1�n6~yc6oP�<I�FՌ*E��TC[c��i;t'^y�<�u�''��ԓ���(m&�z�<i�K<w.q�����v4�8�g��~�<Q�R&�|�sq�V5D���F��<����@��d郈ϯ����K~�<i ��4f�|�$�W�W�6Ȣ��E|�<ᗈ�qhf��f� `0U���OL�<!J�.fP�qBk�b~�3 #L�<	4 �s�2���8#V�S�EF�<U�����Be��	��h�Q��C�<���.W�9x�ϊ�G]�4���TW�<�s��:X*���ӱm0H0+�Q�<I5�5T���$�?�Y�%f�K����>�T�ʹ���� ��p�PĚfCD�<᱌�3|����J`ڼ�Ct��U�<�"�Ȱ-��,I�)߄[�`+u(f�<��V"4��{W��9V��a��Oi�<�1e�Aʌ�a\�?c|-1���e�<�R&�:dX���1��/u��9Rө�b�<�pĈV�� Su*E��~�Cv��c�<a"lS�L8^�
�H"
*���b�<�⪓�hj� ش�%n� ��KS^�<	�育`�ҭ"QD<���X���\�<�ib'p��Ė�-�px�oZ�<��'�"G|��S����nm��P�<q�P�3�8<�s�HpYEJPT�<G΀m8hD �Xh�T�� S�<� �y�Ń w�DR&cٞ 2x�
'"O�a�d�+*���j��f�bc�"O�|[� kn�!V�&��e��"O��8eC@�~�&A�!�_�Ҍ�D"OV��ެw�0 ��N���0r4�/D�����
7�(��-L�0�p8��-D�,W�ƾs��@��/|�� D�,D��;��	x�ՙ��[/��p��m)D����&ȿ?�LTI��*:�V���%D��@6�ģ�����,]�x{�d"D���hƟu?T)'ʓ%e�ћ�� D���G�pA)2DҘ���G!D�Du�T.>@�� `�ح\��-rč3D�����		r �s��/�`�ye�2D�d�7H@	�NX�o0u���'�2D��#��+ jL��ԤX�l`�'/D�b4�R���Z�=d����?D�T""�8R��5�ԃ�:�~ q�<D�p�pˋ���X�6��|h>�B%&D��;6B�q8P$�-T�(H�f�$D���4��1MY
���BW>���A�=D��h����Y��i�����i��lꄮ<D�\��qpFh[̆	�t��҂5D�@y���~�ޑzp,=�T�[03D�B�F���^*5�S��M�T'0D������&l+��F[.1�_#>��\<J�Ḥ�l�5[m4��+��<�eC��>lhU��s8LSWUX�<����0d&9B��E�\ |���"@`�<�o��D�,�@��ܠ-��ې�_^�<�Ӧ�#��Tc�"yc�H����@�<�ĥ��,RA�P;rL=[$��}�<6I�7�$}�"-�;���F���<)v�E�qXЂ�M�3'��z��Ho�<y�Z.bF�a��f^b&��%��k�<�%�V�X�X�hf� G}���a�<!�Õ��H]{���z��%Qqj�E�<��AD� ��5�����7D����i|�<����'�h���'-ƪD���Ew�<Y �_�\�T%k��'7������<Y���W<�<�S�P�Yo��r��x�<WA;��=@OĈt�0zf�Iv�<QG�(^
D�pgN�r��Ebu,K�<�I2��l��OT�Q�,�Em�<��n� 8= � �L�0}�v��m�{�<QAA�tB���)],m�L����z�<�Eh�u �њ��ЩO�`�Q���t�<�'���3m<��W@ĩpz��d�q�<�b�B4r5����D�.P:A���d�<�5
߶V��C�*��,a!�Ie�<!��:b[�d(�Q�@dqІ�h�<!t��2�� 1��T�z�d���mf�<���.Q}bx0�JO�o�r�z�+�`�<��$����t�d�N::k���֫LX�<!$��1+�`	��.�\�(KW��o�<aE'H�<0�Zd �k��0�vc�h�<�&�R�km�ͻ2�8��Qf�<)���$����Iư��%���o�<,�6�l҉�4��Ȃc��o�<a`ᕉ3=l�H��S�&Ω���^^�<y���|X�:�jSG|4�9�a�^�<�U�7�Qㆯ��a�v,��TU�<IrN�(58T�'3w�ttQS�U�<!s��<*�aR�C�/͠�('dj�<qE��j������K�:��#n�<� (�����"I1҅�T���s?H�g"Od��� \�[*sq'M<|�3�"O� ���	��,����T���"O��G�]�r���D�/<�rl�g"O�@������8��F�u�l���"O\x�3���]���T$l��D�&"O�K�Nޝ'E��p	��a�����"O*U�i�h����t�=6ZЃ�"O��j�ރ4d������j�#p"O~a��� �R0�t@�(�Xp�d"O��ʀk	�ș��B�E8pB�"OE�R��O�nl�G��!;2E!E"O(!�3�6]I�HO�v*��V"OF�����r߬�jaH��sZ��B"O4|i�Ԛ2�����.� X�c"O� r"�	rGD4Y��3o�v�[%"O���jJi�������5�EI�"O �R�ܪy�`�8�L���ʒ"O��J��J|��M�4-ՊR��"�"O8pP��1["	P3��Q��H#�"O��AO<8=~��f�} v�u"O,�F$:K,pF
�[�Q��"Obiڡ��3@[J 
T&�V��H�$�>I��!�L��?]��b��H����rm;z�J1Z�F"D��(vKY�J�)"���+�XA��@��I/V2���M\A�3�	�]{�$�Q�o?������.^8���W��p��2C�?lZl�P�&Pa���s�N q7��ۖ����0?ipj�a�sD�Z�c�,�9p �h�'J���L�`��M�4LY�0�S��N5��O�?�DL�QCQ�g�C䉦C���E�9b�<�v�̇���ɫU��V+�0iQ�h���f�O��┊R\�j�{Ї2����'`����GP�-/0�G��"��m�c��.}���b�sB�ya�(ش���ɫ'o�5�!,��V��9�ƛ�������:b 1h��4�+��]#�� �(B��?LF��
�14*m֫�=hTz��
6o�HEzbJ���)���߶/�rU�c%��6V�i�����SRoٱ���҂ܡs�!�$��8t�ÈR�n��R4�Ҝx����Lwu:a-�G�r|�s/V+*�>�ؿ����PV[���χ�� �>�Q+�Wb#|Z�k��DQ��2(�1��!E.ō��{��#��Q�YU�J�X�+�ES�<iWoB1��i��E��� mҧ���<C�\l�AI>�'[l�aa�&ﲜ8��Í�f�y�!��U0����i
'm�H��P�ǚr��z5�8�O.�j�\�B&>����4��i!�P����.yD�J�ED�	��dh'&��	�"�җ$�!uXJ�8WC���a.Q�M|�QkQ�E��$Q�F	�#�$�#��yb���%�n����� z.$p2L% ��2oG�	�ux@Á#�1�Q8 �� �5�	
.~t���jB�ԑC�!�hOTi�b�輩J���%U(����Χ�}�����4.H���{�hzA.ۄIs��s��)��8����Q)��-H��
���
6˗�bRO�1s~�� No�4��Ԙ�!Y�h��L�T�eZ ��)����'3�>���ͤ ��ʰ>�	�0B����-�/E�
��\y&��]�8���v6MjQ�Q.~l�x[��
}�̤�7�0��i�75z�|yD�<h�
ݡs�'��ç�Fu2I�'MO�UB�Y�v$P�M:fW�{�� Be��j-xh�`e��b�bY�ga�S�K��ɺ�2CH���� W�D8���H�h���Fy�+H(1DF���HˡT�H,���~Z��ߛI����bVҥi��ĊD���d��.{-�xŝE�k�Q�|e>D{	�W�\��7�U�Q^*}�B�w�4�A���~�P�KE�Ӆ2�$�T?ճ��߫(�*��g!H�M��BVl]41"�pK�#P�	��2f��I;0BI����e�2F����w�γyG�RV:�?q��N�~�� �'��� &�T�0�9V��:Eƞ�λs2rt/�2�v@�AA�����W=xo�	�n��# \���t�H5j�M��;���L�DPz$i��ѢR�p��S��P�I)?�`G )Qo�88G��Jz�L �kq�'����*Th���s���O��"�G��*)�](��P-nt�1�!AyJ��B�'���A�GX�c��A��� ��&D-��sTI�D��!؀�K*T��S���)
n �P�d�e�Ό�x����h۔
CN�P�
#W��B≋�p!C�(@�_,����\��T����t�<b�%(���2`��~=s�(@��?��	�/�^睦e� T�P�������k� ��;RҰU��QE�? �i�Qf/�:����W�]�0�""�7gI��	ӹ|-x�O�}����=��A A�)�%{�'���x�(��u����Ԁ-�qP%͚s����%��5�A3
0LOf9:!
M"������-_u�)r"O"�٢M�5R���F˻z�u#�"O4���AK9�a$ʹlz|#"OF�`�\SĂ�� Ymj)�"O����dI�@m�c��&tY�X"O�(s�ƄD����7g0�)�"O�$�P�+o.R�
�! ���"O�	S6�Q8}kt�QZ� �ɳ��DT#x4��L4�'F���N �f!�I
�?Y�<���3�8dᑈ)>R0ҴDB0_� ��G A��J�D��Y�x�k1�0��b�2o:f�8��<D�D�-Ȧ83��+��l4�d�mD�Aوt�C�;2��`�ۓP:V��$�Z�>x�H@�A�9_<���뉞;�]@ю��-(J�lZ�]~"���G��(��u��$!�(B�I�Dw�e�b��$�����,/�n�PRq�D;:�C��U�O�Zq���;��شK��1f0��'`�A���!P(�X�B;<{�&ܧFh0*PŢ<�9�gy�ԴZ���@�"�1j9vd`�@��yB+Q-��(��<��=cA���	��z��[�d<���S~�
9���"بON� � �:_b�p	2��?%2hT�'^�ԡCȃ	��||,��"*�y{��sG��Їg�/����	&���B#	��RDT%q� IA
�<I��C%#>5PƇW�I
D���	�2ʧ{q����J�Bp���7s����lȬU0�AI_r���h�2�L��l�q���%��^�b s�I�(��D�;~���8F�
�*t�(�$��ȓ�ڈ����
��a����;ߌ|II�);�L�@�kZ������E�I�t�4��N����adX�%� C�I��>�Bä[6M-�:7�o=�ɠe�J�� ����Kx���pa ��`qc���	�H)+�L.,Or��f$_p�B.O��	�"A�]����s@��2��v"OVI���K5<+N0�Cd4v���"şx�Hl�f��%
_j�O�hG��� �ip�A|� b�'�P�◯=7��l�7�]
/v�I����.��\������x"���	Gk'
R ��k�ϋ��B㉄J� T;��#�*}�#��̐��41�5��I�z�i��O������߄PT����O�f�XH�dZ�a.>�"�;g�
'���R�+D��#�a�+d%LI�܆^�V�P�G%D�dC7"�<��8�D3|x��C��7D������<�����')��I��&D��q׏F�B���#��.l�T�&D�(��kZ "�֑�#�V�H�D)D����_,�6B+b�y�VF$D�� ��C3f��7��Df|�37O.D�ӳ�G�-��a��-��_�Py�Wc,D��s�k]�P��� ��<_`�b�-D�U�"V��`�R"Jt*�+D���rO-؎\�"M�7�b5Z��)D�T�#j�6S6H6�[�6��8�B%D��Ʈ(-���A��25�+�c?D�@9�%F�q��FS��qs<D�xwCo @���z�|f;D�\�S�b���r2�0�ڂ�9D��A� !w"%s�R�����C�5D��	�l�4r �F�N����P#/D�LCS�+�P��Nϥ\@�1AH*D�Lr�C'�8��2gL�_<��؀�<D��3�Z�i��k �6)�,=n~�<ab��/2���: �j���y��{�<�t��AENM�ՊH ��� �Z�<q��&�XI���<`��E�eYV�<� ̀(�9L-Ι �:2➥��"O.!)cNđP��D��8Zل�a�"O�$趮4_e�AbU��0ăp"O�X�2�@)3�F��BF�!�F��"O�-��b�D�+���� �"O�UɆ����0�#����X�YZ1"OX8"tLŘ<mz0A�(�	��	��"O�@��KU�3���zծ��k��Ԑ"O*����ȈJ܉��앤d�:�3s"O��{C�i��rM%sی�  "O$��[��U��
���X�"O�1k`��iЎ��AK��c�.�q�"ODL�")Q�)4"�c S�_ ,��"O�yS�M�*jlJ��D7:��""O.x�d���<���m3$��1"O.�Xo[1}��a�B���,����t"O���
��6�`��c�lv ��"Or$q�����6�V9Y#i�&�y�#�
e:�����@�����y�!����a"$9y5�%cB�yB��.5�(l��́W_���Tm���y��%PgΌ;�&ʢD��kԌլ�y� H�W���S.U6d��y�o�y��¹z$�98n͆^k���Ě<�yb���c�ٺ�G�B:�,�B
��y��I��(E�Y�8��8�r����ybl�&q9��ȴ(%����A��y���P$�0�0`��x9Т���y�T-�r)c�%�3���a����y�FF6/�T�[f���r�DQ�1�H'�y�$�0J�EP��[�j� ���ל�yB�� (�����!�k8�C���&�y�9Aj��4L�Q8���܂�y���)w-�L�dEN�$H5T�Ơ�y�[ ,���;t��m�3��pB䉂��`��Vu�q��`:7bC�6&d�բYC,�隠$��F�C�IiO�E���ZC
ֵ�W�ي-�C�	�s0�� �O4"���
�D�B�1.x�csa�Km�d@C� t�bC�5ż���ѻh݊$p�H��i�hC�(.�sP��;fj~�Ǣ�" C� ���(��n�#v�T�-D�B�ɑt���2�b�4� �z�	+<�B�I�B0�PdFܑn{R���G�@#�B�I�ZZ��+ge���j����@t�C�	�-8M��p^``3�d�8a�HC�I�ڵ����J$jt@eL���^C�I*	�(�g`S&c1:exF�X��|B�I�O�L��3�uਬ���׀
M*B�	�We@����j�	!�g�_Ȝ��'�b�IJ	�F��ࢂ]�H�v��	�'b�2E�"G���R�IJ�M�����'�D�'j`��K:Gp�XH�'�T�i��Q�@!ƍ�%Û�>�>D�'B:��GC��X$�+0�է<5x� �'݊xs�	eI��ŗ/�
ȱ�'�ȝ��M�N,)�cDB
(&���'P�!��d
ta��1=���{�'Q"5�FG6�HtӡDN�9��D��'a��o�w�耈Wƛ?(�Ԣ
�'%�QA�-H��Ժ�Ք�Q	�'��q�8Cp�x�dZ�M����'��!�)��dQ�v╏F^���� ��b��ӯ�P��4�ڤnˊň�"OXY�	��L�Uؕ+=�� ��"O�mz�&U�8����L�Q����"O4P���L�#�P�)q�A�o���1"O2T��"�)K!]���M�j\92"O�a�'�[7E�(�ۗ��I�t�ӳ"O2Ⓜ��f_d(c���O����C"OZ1Q��$x���rL̄C�x�(�"O�1�OSj.i�֌�(`�`@#"O*��S.H�}�ع�7��gOB�V"O8x��FY^��(8P�̻& d�"O6,:�ǟ��墥SIF�@�"O��⭂s�:�ڣL$�RHd"O� �ROY�X��l�pl_�vx��B�"O�K��_�!����"Q�6\z�æ"O�9 ����"@h�6�:A�"Oz�%��<%�Y)��:~���D"OT!U�+1��y�p@D�`��"OP-s���03Cy���:[�9�"O��3!e���
�U	�4Fz�+�"Ozͳ��q����sbX�?��E�C"O�Ԓ)�C��3�D
�~���Yw"OtUC嫒�H��Y�2��zL> ��"O2Mѓ#\�R�^���ҷ>��ٕ"O~B�kփ9�\A�AC~�0�P*Ou;"LL�!V[�����
�'�0ıRǞ�,���/�5}-��9�'��a��ޥt��!�
���	�'���QG�	�4![Tm�2G4\�R�'s�X��ѝ\�ڌYd�_;S4���'�(�C��@�Q`$F*�x�z
�'�z ���0g��x󍏸-��$�	�'��"	1���P�`龹
�'iV��%�T������"�X=�	�'�A������P�C 5���@�'��0P�����ɳΑ�,@9j	�'шM`B)БH��(�hX�-�"���'.��w��As ��3�d���'�� d��6l�#	�-��mK�'t����;j���DW$';ʡ��'J�|�����س	߼�|X�'�F���£�L����J�� 	���D�^](4R���� ��ْ�P%t��'���j�X��I�,� ��{ ؼ��Io-���(؛`�.i�!�,ER@�I�9���!��V�i>�OҗD�R4ET�m(��P�
�G��`Y���X.t|#�W�4���P9C@KG�I9fb̭9�<:��I5&�����Ȋi���2D �S��ISR�pl���6_?��p��N���e
�� �^�ӳf'�OZ��3&ƽ	/��X���	�����G�f9�r��ōqP��@��	:EBj�[��+t�J�H��Ԑ�X�Q���T�]['��7��%sG4�P`�
����#=��}m*a# M�=s&u��-��Ǽ����5�P��ǒKԊ(	 l���
����Nt.�a@#L�j<I#�O(��g�"� �L��S@;1DI�%�j�����gF�$�q�S9T��u�t��D��+�B<�A�ۚ��	6)���㉐ryr�"#.ʈ��o$F̸L�t+ŵ ��<�L�z��p2�<���pѬ	6~;la�' B+�@�`�''����&�=�L)`�|���<���P���v��ד8F�ᓱ�fp�(:�Pi�Sq~"?����E������A��(OL�G����5����Ov!�O�s��%�`ߣd����\�!�g�	�}ܘ�y��3V��`*ÓBj�r�� T&����+#�HK$�-#�4  �L���)���	@�g�ј�nQ�O��@��ְxQ0�ņ.�1ȲGC�� �
O��z��dF�u-��R��z�	��x�1&��\���]�"�2�$�������2Ze<�r] 9#rB�F�� s�]
����D��t{0��d�N�
�:^
�ks$G�kˬ\����[�x����91Kf����J57@땈���g��ɀz L@'G���P�k��|�Q����ȃ|,X �ǈ�	 �X��B�ҳ�Q�h`}�����#�Jq-^�?mI�f��&��S�����)� ���"M�0Kx)�.ԭq��(�/�/�d�Z�5�V�Z���˟ʧ^H̨#%�#+��G
5��Z2��^�m��m��5�N��O��ZP/�0aW����#��j[��&N��&eY){<.����o洍j �1cW���Ɏi\��v>�$H� ��i��ya\!F�)��'�(xf�HST����5-K��פG#}|�8QD��h��X��]0zI~0&�\G��c��:̪lqA�.Y2=2j^�hO����3*YXX(�� �`{�r2o�jǶԓtL��'���'Պe���p���C��UP�]R���_ڨa�,D���ү �uOl�� z��ec+D�L��Ŵ.�V8��¿Ԛ����(D���ṗWU�m
q���T�(��	'D���#�ۤe-(���=��e��$D�S3�t9<1���@�^|āB��4D���A{A<@�N��d����n4D�4��J��)D�\{� ��-5�	Eڼ�z�O�s�O8���7�تI�ĂV`] h�b�'���QdX5b�p�ơ�nx�SV��@�E3�>���>d���B 8�N	�d��� ��[n�<y��C�X��rd�O.<�E�J�W�:P�uJ�D���ң�'��h�g�6kT �� 
�T��TDAc���!]t�z۴{�V�p�OT5Z��z�.�ZՠЇȓ6�PaCI�7n3p(sBۅU$��=�B(q'�H�H������]8/���Z"�43����"O>�hs'�g� �1Aa��g��U�֬B1{�(��PZyrm�r���� :
����Q� �^���|�!�d�[�n�D_���t ]������WM�сO����;�"�4�Q��!/��]��)��aK�k!\O>ez�D�|���j�*�\Mv�9'F��R!��
��{X�i(���qg| "�6��tP��џZ�aV�ξ����=�s��A�x�A'2�����Ȳ9p�єO�8�y����E�H�%j���'v���s���n�
�b��c�Ԥ�%�ލ>r�ؑꖨ-�0ifJ��ZtQ>���w�D�QU*�5'�\��Y�[Y2,B�'�$���250i�NӰGv��Zd�ca^q:sC��M�(N_��4l,ړ*�̘��Ϟy� Y6�]=����2���� .�0�`�q���s��,����2�L&�O.�)ώ+r
��VAW(�n4PR�'0���-��U�Ք'QH�"U�N�@�+�������	�'�vh闇�$���{''��}丨�N<���N(z��Qa�=�'O�<"�AR�+X��5T��i��v���A2l�� ��р��?\�b�Z�����I3~���x��L<�(�j Hq*�D
}8W�ah<�Z�N�X�f�C2#�l9��+W¨!��Ł�0?�G��,u���J�9��q�Qj��� �F���*�*p���]�/M�|��fY�Y�td�ȓBE
�B&j�@z����t��ȓA^��,K�s�r�`���F�\Ѕ�(�A���+%!�� �j�E�����'�2�����Ѣ�1VE֌W���SV��)�#@�)�`\!W���RP� ��ox�+t	���<)s��ч�Z�m��k�?��|�΁�i�d0��Oq4��
��	��=���׿|�ȆȓMc.�K��G]q ȢE'R�)��:U�h0�F& ��$���}hX���1P�y�D�'h��&�3/����?:3a-b�֥hO��l�\���&�X���B��M���a�%�r���C��uY�@�'n�ח(K����"ONIZ3��X�܃�"X4�x�k�"O�(�A�G�zoH�  ��@��"OD0A��)ptAV.�lI�"O�\�a�[{Lp�G�A�з/�!�$фE� �Æ΃�U�)�/#V!�Cjz�('��+/�HD���d�!�� ���V�ב$22Lc��܁Ix��B�"O�TYgb�11�aH��Ů$c�A1�"O0����]��p
�D�1NUi�"O��ҢoN��P�GJ�h��s�"OHH3fD
	T!0�:A�Jb"O��G��	-`�A����":>Q��"O�%)G�Z����%���Q?���D"Or����� �Г0G�28p�"O��`���L�8�Ԡ�g��K�"OV�� �\�FP�"e�.~��8h�"Old�*Q	]���#J�{�@I"O��M�)�m��[�6��"O��[s�C|K�,�iْw�6��"O� �G
8��c�)�~)�6"OV��1�T�/��D�A�v���"�"Ȏ!siE%3�fM�d*X+|{�y��"O�exA���6'�ur� ��8�^�H�"O��X��[2ER�hïId`&�
�"O,U�WD� ����c�DV�B�"O0\a�N�;� �v+	�
D2h:�"OvQZ��� f*xv�_�P��D5"O�Z����杉��I�Fp��"O2�JK�z������a{d�:�"O�Yᲅ!xd,�qc�4b�}��"Oʼ��m�2*��H2��wU���"O���Q�)^�*0�5�ͨ0X�U"O��TW��`�e��&��TB�"O\�(�n���)#6kכZ�B��"O":��%w��q8G-�0;���"O��)��͏o���kY�<�0�"O�)!�G�@�}Qj��D��]�"O9�s��;k��xG�8}�1#"O&�S�抯 5�P���{~Pq�"O��y�b���1��2��%��ɘ8`B�KR�F?���f_>c���	�Tm"`9
�"�(�pӞ|;�C�	�~��i����1���O�Y��C��.E��\0��	g��Q�rb�'��C��>+4�����g�$��$ˊ�L	�C�ɲo�(��BD�'�5Pe�)r�NB�Ip^��;��O�Z��5
�*�B�	8��KK۬��@��'��]c�$�?}�O��b�CF/O�JE+�1Of���,��'>f"|2��G�!w�I�Ly$DU���[&]L��$�Π�Gb�a�����q��Η����h>V�La�aOYX�~�qA�I�)���S>��b*߁h^X���cͽ=�h�Y�E۸)�����E,z<����.�a�D�֏,�8���Ywf�9��s�n��2��K?�#���`�2��O >�Ѧ�=$�^�D�P-�|�G��l���	�K�����>x5��'z.>���I%q�� #��X�DT10�y�8-�4��`���*�)�<)�l����/R"U޶�Z&�����6���~� O?7-)K�ꌨ�KA*IYبp�$ֽ4wP��Ɠ0b��2a�P�0�A���wVh�ȓ���3��J�9y� @�S����o� [6���iC�2�,S�m�� ֺ��#.�=&�8���!�]�I��z���; ҏ���*���pm�ȓgw����A�}�$��#����C��2s���*��\���R������Y�'ۀ@��,O�l���܀3��'4�D��� �%ɶaD�:d���'�B|k�b	+����W
�<�i	�',H2WK��n۞��@�~Ars	�'p,Dz��HyRT3���mL����'��E8�#��f�����
 qQ�d��'!l9��,M�)K2�ĦV�Q��\i��� Pp�P�M/�AY�($*yRĘf"O�H�GB"r�4�V�[�����"ONɡ����|9d�%Zx&u2�"O����9��s$ �2uJtr�"O�P��Ě5oL8ci��`e�w"O�#�Ά=��-���X�]��"O�`�kG9@\��o�H��"O"�Z6��.�4��ĦO�f7L0��"O|�a�,��=5��%!	&���r"O���eپ/��M{�N\�}�t:P"O�ICVG �@��p�v��m��0Sd"Od�ȓc�<&���c�%���y�"O�k	To������D���$"OP5��J��7�R��"��G#���C"O$�����
T�R?�EPчV�w�!��*pF�&�[Xۮ%p0��0k�!�d����|�Ef��|��F@�2�!�D�,!�Νu%̍"��Pag�
O�!�Uxn�!!�J��(ܛv䎧k!�D��)����FK$%�E�#!�A_!�D?_z� ���3r����W/.!�䗱��0�g�h �}ae��*r!�$�(��a�Y<`d L�q˙�|�!��X(b��}@�w�lp�E^,#�!�d!}��!�!#�&;����쏍m�!�]�#i:`���C�
#���F�=%�!�dT�kD�2$�ҙy��'�+Y�!��=]�l㧂,$�.�Z$��'C�!�DU�E�
1�3��~�c��ˏm�!��>,�mRg��L��a��47�!�?MD,a�T�b� ���&p!򤝦��q��&�,�6�(�*P3=h!���{���g�֨z��`��JN�rf!�Ď*e$dB��_�Q�=YG��,�!�$�#��P�U=���o>����"O��1���St���U�PH]��P"O���Wq�gO�R(�\��"O����g@�F�(�x7�6#��{"O�a�'���4|���Ev4����"O�訁�/�,y`�B�d���7"O|��󃀭c��9դ�)�4HZ!"O�u�'�=i^(ˡK���B�"Ol�G��78��i�sc�!Y�N�T"O`E��؇F=�}鷤���y�a"O����s�5��J��l$)�"O�y� ��Z������DE�)`"Oŀ��]�!L-ۥD�+<2d��"OZ	 6�E	-��b%dT��"O����_$aNM�#G	E=r�;"O��Tk~�Թ�oZ+C
r�"O�}���0 ��Sр�4=��Ѡ�"O^��B=)����/`� ��"O�m��bͰn\,3���,�:mr�"OΠibdH<�"�Q��}�ȹ��"OR�$S�)�053�\A�"Oa�`��/��Jq�E0:��p
�"OB#tE��Z��!����	�-4"O<����ŀ;.q��A�#��Ss"O��KG/XU�`�[�X[4�F"O�Ћ�JX :�|\ ��\G6}.8!�$�;���J �.?r�:���3 !�d͐ƚd�q/ͫ0��6��,'#!�d�?`gdh�S/��p� �E�!���U��ɲ�L/4���!ܷ_p!�� Z����
,bWLe�G�N1�ԩ4"O^��.j8Z�b󏐱 �ҵa�"O�q��D�zNF�θ9��ذ�"O���i�6;]�i�� Z�v�P$"O���͌�]�z���:�MP"Oօ��N��nXqꟛB�*ј�"O���5��/I� zc�]/D�!�0"O*�+��F�o����@չ)�x�8"OP�â�Ґ(��E� .Qz���4"O��X$NL`�r���!`�����"O�,B��2����эظ-���1�"O���Ok(,�C�_]���"OU�!��4�$u�lѠW�
�RD"O>|���ܞ\bX��$[�.�BPj"OLɪBE� y�A�(Ma�(��"O>xC�M\��s
1� �S"O�eHCNG�"Hl3�	^�X�.�r�"O �8	E���bڻ/E~L��"O��cu�ʢנ� ��ߚ
E��"O��
S>Xo���Q@Z�*�"O���Ā�qy�L�8$ �2�*O�`�B@/H�d��QMǞ~��)y�'�21�J�b�܈�B-ݓzX���'!�T1��	�[ :}����=y�v5�
�'(���"�Ph����gV�a�'���-L�$����̸~��L2�'pjE	 DχC&B}�2AX�$ �	�'R�L���L�_!j���#�o�"8`�'�Ptڠ��C��H���O���c�'��l�����R:�HI��O1q�:	�'	�X�g D�]���Rʉ�)��H�	�']9���==2�����ClM��'�4Y�F��%~���kG�T�'P����_1*ҡQ�R�/4<`�'�`X0#K����;�E�2��d��'UY�U��N�z���ݖ#=�<��'D���<nbi##��%,,yh	�'�>�F]� +��z�����'�*��&J=>��qӧf�"I,D��'CZ]���O� ILd@�CL��J��'P }iG!�>P�� Qr��4��e��'I@�ۤ��:t�`��Ǜt���H�'58�PE�Hk�����3 �b�;�'�~�(�Oކ���BY��'_��8��]�ux�蠀������'@fmS�h�,(���Jђh) ���'�2[��ڽPQ|8�f`�'r��e��'�8� � 2�nbуG65J�Ͱ	�'#�ȩ�,��r�K6�P�'��t	�'ך��#��t1������
� U:�'���Ð �N�d�v�J%S�$��'S����݉@ �lنdM5F���'ތ�"p� �=V1�׋6=	@��	�'(ehӠкvJ!�AV:>���	�'[R��`"(������+�ʅ+�'BL 3C�D�ݲ��9YjN��'�rhbf��4Dc�Q3�AC�g���9�'
�YH�*�'��t�P^�0���'���Δ?��+S��VG��;
�'��|����$VgZJ��ӪB��c	�'dH�V���}��g���BфQ�	�'�@��g�$=d������p@T�[�'[6ݰ������@s��x�F���'��0������B��8�J����� ����f�3(��VC�DP�tY5"O�rĦ�1w|ꑻ�cL�V,�u"O��N�v��'ȗ=}-(E��"O��6�_�@y�A�����*Q"OzA�O�=J��0Њ���[�"O�`������s/ۿ94d��"O`d��
,�[�o�/N���"O���O�7�`�ĈV�E*B"O&M$#1`���H�ߢ.�Z(P"O.,@��P���x9T�o��u�q"O<#۲+�����vp`  6"O΅�,�+G���8�	 4�t��"O"�2�`XL?����ǣ1(� � "OH���L�n���Rt	˰w��sW"O��25KG���EX�H^!�P1"Oz<����Q!���f�łek�m�"Oh�z�l�D2r����X� K&"Ovu�Ʒ9��(��cA!@�:��+D����V�-�'���2�l���+D��X!���|���] �0��a?D��_9�49z��ׯq��L��y�-x��K�\hU,İ��ք�y�W��p��lZ�g����R���y" K����I_
j�&8��X��yr�.I�F�	�h�%d� -��Ս�y≗E/b!����p>��X�߹�y��J �H�d��%g�>]�O�*�y�lB9d�p#F���4�|yQ���yr�G8a��&��dh|���
�#�yBX�i�Ry�d%_��T-�r�+�y��1e�:�*�◆C�h�*%d
��y"�Ec����qF�d�ټ�y��O�t�6n�k��e�4� ��y�O]fq�l�W��&$]�7��4�y� ����*d����E( N��y�ë-d��! Â7�������y��G����aĤ�U�
��yroIR� (�D-%�-c�)߫�y2��,�P��b=z88ID���y���U�s�(�	s���p��E��yeY3�ތ��(I�|L �F���yr�Ak�N�YҠ�'��5 ��H��y2�Uz�ܚedX VM��`Beˀ�y�i�"(S����>UeF��+U�y�AC�f!�s���QfVx3K��yB$Y�-�l�`J~z���u���y��_�5a�����x��Y���yb	J�J�$�Q��n *	c��ɑ�y�J:]뢅 !cJj`N�5��ybC�C؆�*�n�T����U�9�y����sfF@	���=JՊ�Q����yB��76�;SFԛ/>4�0�i���yB�΁hG�L�U ��'�Rax�'�yb�PiS�"$���h��F��y�ʕZ��D ��1X���.���yB�I�nT0�䥋�E���N5�yBDm�ֈr0��hz�p���y��T#����n �p��3�y2Ke)
q"v�B�8(E�W A �y�D�	3�(I�&�0�l�ِ���y"cِ/A��y7.H
}�|�Q��y��A�L$]@C�،Jx�H�7�]��yrF�R̀-�0 �/��\�A�yR��3j P  �|9�õSy�$�eP�ybʒ!v P  �~�<��ꃓS�#Ɵ�݂i�qh�\�<ɔ�x����ŞN�F	�2�Y�<aţ��,���FeC"-�\͹IR�<��ct�h�p�� �n�!f��S�<1f��y�P��6W�5kaO�u�<���ȸl����LZ9����Zs�<Irψ*�4���8]2,;��K�<� �ۏ�F�b��A�����G]@�<y���XA $#'d�t���`�!ZH�<2'�Mfv3 �����b
G�<9���~&Ƭx�@ĚKe�Y!�O�|�<i׫R;{h��r��E$|E�el�r�<!6!�b�p�q�%J���8r	@j�<�4+�>B:���c/juX�kGb�<�W&6,$64�jR$��1����Z�<�aß�LtS2)P4�\����DC䉺S�Z�	�/��r�S, ~C�)v��t���H
u��p�g�Թ1�JC�Ɉ)+�!�+ݚ*z�C�k�+{t:C�	�lk� 3�6�Z0A��ØE�B��)^J ���u�Ɯ��@_;E�(B�I�oڜ��4�Q�kY�t8$� �+�C䉩?ؐ Q��?�I#*ҫ19�B�ɟoI\��g�3d��҆Aл!6pB�I�[�D�D @Z�&�{�&57�VB�	PL~���:n�Q�]�,B�	�u�Y��J�&�,LqB���C�	�>.�Q'U�Y"ɰu)¾J�C�Ƀ&蘴P��*������"T
�C�I��ek��A�S����tk
�k�����B```���6vӔLPe̌ZN�+�K҂= �[R�Ϲ!�!�� ��Q	ʝ��=i�̄5+�:Q""OX�Y���E�������g��Y��"O�Hq��Φ]L�H9��њ*���b�"O��(��ɜ@����͵(d�M 6"O2���+*��hH�ATvh�E"O���qZ('����fH2{7n%�"O�b��G1D��LhƌE/L���"O ��!�K�/�2iX�*�%x��iU"O�@E��iV�ǉT>[hU��"O6I��v�~�Е(��pO���"O(���NO��(�Th��D��"O�����K�xfSGG�q˞�!B"ODX�`��� &Y�v��q`5�'��0pn��eL�R�*E��,;���F� r�Ì�x��i�Ɩ�b�4��g�O z^w���
B�iΙ)�*}CB�L�vf9�ǉ�b�䘑2���$���d����5/�p��F85�tԠ��Q�W��]���>�QaU#d�P��I��f�x�b0u?�y�7*B�X��'�|��2O~�"�}��b�bLQ�CA�u��РCCP�'H8�)�b�N�S�O�`�X�nD1�h�{�����+�O������![�1��K v&�Zbɖ�ѲC䉃D�z�a'�#���B�.'��C�I�AX��A�˕)T��ys�IG�Y!TC�ɎY�$�Rb�_8�$Bse_8�"C䉬5�0���	�7E�L�u�҅|�B�	'%:Թ�7MF�!��H�є��B�24�:��2��A��x���,��B䉘�3��ÖTz���<YU^C䉡6��`�cM�*	������
�HC�	�y�`4JTȈ5ch�s�G}�C�	29��I�ǂT������fM
�C�I������ �:�\����*B^�C䉿GS|���L��ߊ�M(nC�8d� ���K�V�8!��ڞB�I�d����%�%t,�q�6;�C�l�D��"��U��a�䊙@y�C�ɩ~f�����7��Q�h�8\��C�I:S$|�e�s8tyz��ǘC�ɕY2�S��
�
�p����!�fC�	[�޸�,k�,��h i`4C�0m2���w�X�82�`?C�	�{�^X��낁	E�0-�7i�B�ɂP��Ŋn���I,"��B�&QP�i�O�#�T����
I'B�	�t�Xǆ��;�4lZ�oZ')C�ɤ:(���wA�Lf(�R��=@.�B�	� P���aD$,\2¦�50�B�I}���iBgҷ�!JfB�	�"���F�4m%��o@b�C�	%<|�1ua��P��гF��+�
C�Ʉ~f� ���[�d��Qa��\i�B�ə"���Qō�F��T�K�;@�B�<g<\bU���d=3�����B�I%bѤ����I�i�be���-4��B�	�z��t����b�:�I�I�i�^B�	*`t�P�S��&q�Q	C�Q,�C�ɜ	�~�xP��7i*J�A�^C䉏	"�� ���cT��U"C��"M��L����-����d��;;C�	;u{��фF0'b�����Z�C�I#�t��p�ۜ2X�X��N�5
�B��;q��u:U'�>^�NA@���:%�NB�!>�@�����@8���"nT��ZB�Ir��1�"׬_0�` �Jթya�C�)� ���PSJb�c�4��A"OT�i��l������L/ d��"O$Xc�[(2(H��K�u����"O���d .TǪճ�E!vH���"O�)[W��o���A��'
=:E�2"O|�j�&^.;��u30�e$�e�"O �NI!��r n�:E#�1{�"Oҍ�PÂ,'�B��}ȨaG"O4]9��$���#�L-���"O�\��[�D��,�/s��<��"Ol�a�K����(X�r������yBg�]D88�
J4���$-۠�yҡ͚"W��;�OB�7~�q�y�aGj��.��5���y2x�LA�H�X��T���yB&��� 4��A)��o!��	$@hЬ�Z'��;�� MV!�d�%-ΐ���X��Q��}�!� pGr� `��9n�
H1�DT�7!�S�S��Q�M�ʭJ�nF/QD!��΂Jq*�P�i�q{�!�.ZhU!�$<DBTT�pl�,J�n�bE�^.!��A5AҖ�k��N�X��-*�!��h!��K�P��q棎�V�"]: �/!���H��i�c�:h��RL�}�!�X	C �@�*^�px9�iݷ@[!�D�gcH4��FN,�%��)N!��
X��U�_*d_�h�ta�.�!�D�!�~����ͅi}�uI6� C1!��ǘ�
��f�P b}��X� ɗ/"!�2jShq�'ӓ	h��+��2I!��\'U��4�S�z��Q�τKf!��@�}C~���Ú��.�BC.��0A!�R��n�p !�?�D��f�-Q?!򄖟W��0��o'�*Pc�)��S�!򄁞?��p2�a�<�� �O�!�D�:����5E���"�S��Ww!�	%� ��H�Y�Fi�#�x�!�DیB�F�����W�X�7LCaS!�Jh���B�� Z��!���>8!�D��nŖ�3A�mb\!H�y$!�d
�7��5��#YcT~����@!�
�S� �Ж ��X�<���E�d!�4T��$3B��#��
E\/c�!��[ U����CN!L����Q6�!�dŖO� �S�ݲO⎤ �Ϋ�!�$�$l�P�����
pnh �̆�!��h�
E�����h���UIQ;t�!���{���1���g.ҙ��A�`!��̌3Z�|��B7�D���a�&G!�ȔM-�eGτRvh�<!��P�Zx� AABϮM7���P��.;!�$6_CF="�%b��P�4&!�M�Ԅ
�nJ$K���3�KV�vb!�ټbL%���[�|���*i !�Dk�V�<b��0 j���!�d�#C�T�%W	���si�$}!�׋v�h(�Q�ϼ}�����!��Z.�� ���_�᪔%��e�!�䇳0
��h�k�7y�S�bU�NS!򄞎l�y2gb
2Ba:�AQ� ���dQ1��c�lط09`��PBۻ�y�I
m�$�9�G�/����l\��yR˃6"���d�0�ցK&DK!�y
� �؃D`ٗo��� �ć�2�<XRv"O���$jIg��	��F>\��f"O�`�J�a"lx���9;ԅ4"OP��+*B�j��(��AT���"O$�f޻P64<;�G�jBXia�"O��!���8v�9���м%Anx��"O"�r/!@ X�-53F���"O�)R-�W���b޸X�bi4"O�y��9�(����^MR�A�"O:��g�y?� ���K�!J
���"O�) P,έR�D����8l�
�"O�s��ۼVR`���E/>D��"O�+����"�V���O-�nyi�"O2�D��65_�9��ӹb�Ą�U"O�X��Ė0|����A��q��"O�����(W�L�K��M6 ��Y�"O��r�勲";�q�\64�|k�"Oؙ@�hZ"W���cP�"h��E�"O����Ԃfs~e�$&\�{g~�a�"O^��b��?{�ziS兗:H��˗"O���g�^�e���p ��*��w"O.���!�<���#4,��m �ab"O�Aװ�ȑ�0ʫ[^�xe"Ob��ΐ `��Zg�B/+��p�"O��`��Fo���(�,)h�sU"OV��ŀ	R�$�c�3<XX��"O�q8G�F�7��1��G	H��"O��#r�E�1�N�A����]�d"O�0�l͎^Zh��!�ѤR۾|a�"O*!�!,�6O=������L۸m��"O<H�% � D�H��Γ�
ìhsC"Ofŉ5�M�I���m�2|�:��""Or��5�2&�m�@-B��-�"O|D*F�C9^&Q���Z�~��e"O�5Y��ɉ>�XPS�+ר@W���V"O�\����3�l��e
�$g@�i 2"O���V�®:�D�3�ȇ�i����"O�y�%G�#|ea&mN��� c"O�Yc)W�j)	E� %a�&�)�"O�(Y��?��9 u�����,��"OX!�U�2w��H��V
^fB!��1ik��̀�wJ6Mcߢ�!�D�%{�JQs�%��B�@�T"C�A�!�$U+�8��4n�q��D�O�L�!��0_CȄQ�ȘF�������%�!�D��|8 �*E��JEҒ̆��!�dM {=<Ó�>Tmn�3*��8�!򄍇,���ÂE��,��*3gUJ!��E�"`ak�h�30�x��@�0d�!���>}����دa�N���	�z!�dߴwĔ��S�w��0!B�ja!�*	~$M�#�ۡ��;�*W!�$�P(cE��eѬ5��I�6J!�$�;C�.U�5���d� !4bR�#�!����+��ř8�!؃�߃a�!�4��t�EN���|b��۬,�!��F���I���p��UqO� c�!�^w����t�\	2H��R�R t!��Z;\�� G' N^�`@�V�<;!��&nڐ��ڷy\:a�"��-!��=Ғd��G��M������?'!�$@�Su� K3�Q56hV��r�K5�!�ÏA1�ܺp��%G��u�+-7!�L�X���1!AP<R�r��G�Rg�!�� ��I@"ٜcLxA�D�?�պ�"O��3c��^4�ū"A>:�PȀ"Or�I#���T������^�)�p"O���B��9&"���ӎ:j%��"O�tVG�S,�9��/��H� "OH��f Y�j|"�Q�)I41��a"O �.�wƴzv��^���"O�p�3��7!STE��31d���"O�ͣe.&�zp�S� :�!"OF��7$��i�Ⱥ�M��B�8x�"O>��v�Bt��p��.�,�%"O��G��#/R&�S#�W�ƸX�"O8x:3#��8$�H���<a��,��"O��X�!˽#s|4��׿xR,��"O��ѡFJԑ�"C�1����G"Oz0�D�)r3�@3���X��|��"O�A��+�b���)�>5q��""O�[An߀�
��Ǜi�b�"O�}�G�[�G��|�. 9�r���"O�8Xwϑ�_<P�s�G�ʂ�
�"Op�"4iI �4u"U��v��c�"Ot�#��N�=QL�k�	��H%C&"Op�p� �,����gS�;J��#%"Ox��Tl�a��}�Q,-VӦ��"O�\���W�-B�k�>�6Ix "OH���B��R+���lP�\�2�Б"O� 3�֥^���vK� ���"OP݃ad�z�q���۫o�$��"O��a�   ��     G  �  �  �)  )5  t@  �K  �V  #b  Tm  �x  ��  p�  �  �  x�  �  ^�  �  )�  l�  ��  �  ��  ��  \�  ��  �  l�  ��  M � � p V �% z- �6 �= WD �M U �[ :b xh xj  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+��6\�
�<4�d5h��'�B�'���'	�'/�'�B�'�TP�`��!a�dYq$RB�x( �'���'\r�'5��'w�'H��'��MC%���g<���]�0�AF�'-�'��'#��'
b�'���'#~H�DJ:%�^yc�[�U쬐��'_��'���'���'��'�B�'Q
�rՀA47�(Ӵ$�=>/n���'r��'0��'Mr�'A��'%�'|��A�)M\Ȱs���a8|���'��'���'���'[�'2�'ł�
��;��=GBJ�i����'�B�'b�'���'�"�'	R�'��i1�n�?�L�'�.<�f����'��'	��'�R�'�B�'�r�'�@�`�B �~�6��ǁ�U�Y��'�B�'���'�r�'O��'2�'��`�B��WGd0��%|��<��'6��'+2�'62�'Qb�'���'8���F&/s��A(4B�1�%��'[�'��'���'�R�'�"�'U��`"c�P�P8� �Ńw�8���'���'���'(2�'$��'�2bM�%ָ0q0M0@�X&-έ,���'\��'���'���'�B6M�O>�dͳ_�`u9���4^�}r�AV8�'��Y�b>�z���瘝 C��rs��i�99�E��^� �O��oW��|��?�Q�952�b��d̔��&*�?1��MO��y�4��Dm>�������sXT�0�
L�VeF�˂�̕(�c����Uy��S�:��MB��v]G�\f�[ش0�M�<����Kw���?�m3Q�D��	��F!�X�$�Of�	`}��ʀ,r�F<O��(�_�S��kejC3&�	Ie5O��I:�?	a�;��|R�-�`�P��O�]F!: �y�,͓��� �$�զmp-1扉��Zj�{3. ��.H62uj��?aV��	�t�S�Fٴ(��A
���N4���������O\q���%9�1�\u���9����̨aSJy��[k��(ɵ��=v�ʓ���O?牟uhq�:)�J�ƥ�m8�扉�MC��i~R(d�N���,غ�$?Z~e��'ש/d>���H�	���QiT٦�'��K�?��@�V8]�|��F��mK^�SE·@%�'O�i>M��������$��7"�0������={4,�>Y�\�'r46�=G�����O\�D)���OP,s4�5ز�r���1���vdZr}��'B�|���� >-��N	(p����ÞE9���V�S0������^H���e�ړOZ�Z1�|�d�$����@�B|B�S��?���?y��|z,Of�oڑjv���I�.��6�$;ް�������x����M�J�>Y��?9�=?��+Ӭ ���p���Za�穈)�Mk�O˄����z����wYNcC꛳�p�ͥ6I de���I���I�0����
��7!%�0V�D�7	��?����?���i�H��ȟ��n�e�ɘUl���h���Z	���S�4�%����ß�(P`Ymn~"f�[���Ca�h���z�ֶ�N�ȐJI~?	N>A-O�I�O��D�O��ɖ�C"�,e3r���a��م��O���<a7�i4�aC�'���'��ӟY ��`��jx�q��߼^���z���̟��IN�)*f��_1��!�	/A��5x�[�3a�	�dd��:B��R.O��?q�j0�d͹Z�����Ǌ3�HLږ�ޅG*��$�O�$�O����<���i�+��|u��&�)��j�����������ڴ��'P���?ѢGG�e�v�����
!;�%E�?��m��5Pڴ��D��J$`�c��d�A�v8��;>I��4����y�Z� �	���I�����0�O2|�`���,��
G�)��	��d�LE����OV���Ot��T�$�����%n���: d~pٱ�T�,�*]�I���'�b>5qu�צ�MČ��L��tJf�8g�Ȼ[��͓
�d�۷��O���M>�/O���O���f�d�U$Y<�TQ�Y��<��ʟ���FyR|�t\��"�O<�D�O�Pz冁=i��M	f�1F
�h��J(�	&����Of�XBt�џ|yɵJE�dj���	6?�����.�T�#gS)��',���S��?a�/�;rڭ��#� =�@�vo'�?���?���?Q��	�O���1oni��(Ͷ`y4�{�A�O(�o�3Q�������4���y�g8wY���(G;���u�̗�y��'��'���ـ�i���"l�~�1�՟��w!�$T4,1�wU�+����!�d�<�'�?1��?����?��@�wJ��Ĉr2Y2�A�*���٦��$�����������gKCr�ZA����!ud�9"�&�����柨��Q�)�S�7H��f�Z#O3$@��BГg	2�ߦ	+.O�<Knֹ�~|R[��H$��	���X�`�<3@H�#��ş,�	؟X�����@y�NiӖAS��ODu��j̀)�h1�ţ	�Q}$qa�*�O6lZo�0�I�H�'�`ÈݾT<�pP�A�%iL�ժd!J)	ߛƛ�4�6�R e��/]�S��� �ez"fB�.���A]!;��+G9O$���O��D�O��d�O��?YȔkĘ�hǯS����R��ğ���ȟ���44^R%Χ�?���i��'�����J� $I�(t<���y"�'��I�F]0@mZd~�+�������H[,yb�O�`����ʟ�$�|R[�L�I���I�(Jde��2a�@�tÆ�;�ִ�ů[���	Qyrmr�j�� ��O��D�O�˧9�D����j�� �L~\���'.��?����S��DȜQ�,c3AͤK� ��EɁnK��Տ�5F�d�O�i]��?�$�0�Dψqԥ�+�����o�=gq��$�O:���O ���<�iz�JP!½!Fl)�w�;e��u�!��:r�' J6M;�ɶ��D�O�)0r����aQ�-l X9����O��DP��F6�&?��F�kGP�I:�dlL�|e�TK�v�bP�`,�yrV�`�I埘�	͟���⟘�O��$k��H]D��!c׳1��tk���ɫ<�����'�?	A��y�e\=2e�;�:����!�Џ9R�'�ɧ�O����R�if�� >��rEd��G�H��w ��]��DZ(MD��[�� �O���|��#���� �ʃLV��+�%N>��!A��?����?y(O��o�0w�1�	��ɨMY��(ٛyІ� �m^8cn��?�@\�X��˟�$�D(a���w5h�ħ��j��u'5?�gIJ�%���4ޘOHD��?��B���y"�&=w�萇�,�?I��?���?�����O|�SiE������/}U�e ��O0$mZ2���'��6-"�i�!��C�2!��m�ì*������f����~yB�Q������I�(��C�T%Fd�����]>�0�
E ��U'�4�'���'���'�'S������}$��.�R��T��ٴA�r�����?���'�?��j
24A������;o"�:�#����؟\�IY�)�Ӎu>�9��A$x�A(q�8xFE�2��3G4��'��E,ݟ4�@�|R\����F
	Ab�iTI�AF-X��]ݟ���ğ���֟�Lyr�u�vɨҮ�O���¦�P��L��&y�ҙ�S��OTdm\��h[�IΟ��	�����D�~�+2�M�%U�T	���.SR�\�+���RE���>��*ix����Ҝ]}�<S�%�.F�F��t���P�I��p��K�'s:h=�7�7y���.[-<����?��Hƛ� ɔC��I�M�L>)�BD�C�eK��U?h?�xRa�T��?Q)O6@s�r���+(��C�:]�����Vz6*XZU!��<F���@��䓾���O����O���"cfm �N\v'�𑑥Iw�b��O�˓;Y��!ޢ�R�'W�T>)�W�3e�Ĺ;��<; xH��� ?�PZ������ '��'Q���0��^���3HĿ9���eJ�;�f��˝j~�O(��	9Ua�'c��f�L(s�`���K>��V�'w�'���O��I��M;�o�`S6�a1��<k�.$�����[��u���?	��i�O���'�OP�^�>�����( Y�P(�!W^��'�LS`�i����~m�S�O\�:����E�E,� �f!=JCv	����O��$�O����O2��|R��_&&n���+�(oS��Sq�I
H���eC2w\��'!2���'�j7=�f��t"D!Ml�=c�����%s�a�O�b>�2���=�mDT�uM�w�ڑ���[�zA�1Ox]#@�\.�?�n:���<���?����%�=p�
A�K! )+Pf��?����?i����$A¦�Q2��@��ҟ����8�J�QQ�I�JD��(�"AK�g������h�eW���IŹ%�
��1IS��sK�$	��0�M�&��DKw?���:�I��#�;z���` * ��r��?y���?����h����7(�<`�2
�� (zѲ&�IJ�d�Q�$E�D�ɔ�M#��w'��C�*��]K7�̢u�X�+�'�B�'��)��]F�v���]�u�\��3)( 2�ƹd�%q&�[�5��Q���|rU�,��ϟ��	ğ$�	ßD@�Λ� Y�� E�3VDz����Qy"q�Q���O��$�O^����ɫ�����@�gO�ѡ4׽. f��'G��'�ɧ�OM:e8v�^ M��tX��0��pß�k%����X����q�D?��<q&J�u�N�+�K�"z��=��G��?���?���?�'��DQ�Y3�����q is"��E lA�!D�| 4������C}B�'YB�'��, A	M�@���"Ք���(����f���g��,%�4�	��R�e��,��%���Un��LI�6O,���Ot�D�Oz���O��?�Q�F�	�J����#�v�e@�ڟ�������4�&��'�?��i��'b��y���}����װ	����y��'�	�^�t�n�c~2���z]b�e�d3�U+_�)���Xh�~I�I�dz�'���ޟ���ȟ|��N:0{@BȌ-��� +�=7�M���x�'a�6m� �$�Ol���|"V&N�[�n��d*�4o��5KV~���>��?�M>�OxJ�(�*�����O/W�:B���!\��i����|�a`��l$��Aa��s���
,�ld�%%�͟��IП����b>��'M6��7S������Q�0EWS��\9uͽ<1`�i��O�Q�'�� �I���8�͔28f�Yg��G�b�'�҄��i��iݱ9��T�?�Y�W�� r�����=n2�q�E��rޞP(t7Ojʓ�?����?)��?Y����iC�^�����,�{FrEr�ߒuBtm��U�	����G���H����`&�=CDV(m��g��?����Ş��Y��4�yB�A�>#���Wd�)�j����T�yb��|U�a�	�xD�'Q�Iџl�IU���Z�$ɌD��/� S�,�	�����ǟ�'��7M�BG8��O�d�Wtڀ ��%<ޝ��lY�h( ���O�$�O֓O�Hsg�̡��E12	�S�,�瑟�ba:0��LXo!擿0��oAП|P�B�/�t "�iP>�l���ß������	PE���'����f'�#k� ���c�HȠ%�'M
7͚
1^~���O�oS�Ӽ3��$��h0�K[҉�����<I���?���J5�u{�4���Ӗn"�d���S��%�ִdI�8��,��o�`��,��<ͧ�?q��?	��?م��� Ƃ����g��5L@5��D���Ґ���	ӟ�����%�@����qc|�0N
6|��ǟ�	y�)�*�<  +�/�(Њe����Pyq�K����ٗ'dN�Cń���"��|�T�x�F�J�&��a�2,б���C �U䟔��ϟ �I���S@y"�b��)�J�O�d9$e^�z@�yzV^({[e��7O�o�w�|��	ğ��'sd�BC� �.�yF&,d����і8��v�����R��TH y����mۄn̻-l�;��_?8
���bp������Iğ0�������2K��ݢ0A���/q�KZ#�i�	˟�	5�Mk@��|j��9ț��|RG\�(	}i�< �����l�Vq�'L���4�����V����&J:mB���P��0�L�C�eԊa&(��v�'�
'������'v��'�R�ӣ�=��5��Q�q d�'��\��:�4I���I/O����|2ワ$.J0���T��j� ^~��>i������F��|���|�2�I��V�h��@uҦ���ƾ<�'���������zhP6o�=y�R��#'�2ߤX���?1���?��S�'����H$�O�2��]!�R��1p̕���D�	՟�s�4��'X��?��@�UV�����#V���Ղ�?I�e�R��4����T��K���/O�m)q�͏�hJw �k8�T�#9O�ʓ�?���?����?�����O>�\�8C�� CU$��C��m��\f
h�	ş��	]�Sşd0�����,V�̼��V)������Ζ��?�����Ş)�"�ڴ�y����Y�I�r�c�ݣ��]
�y �.�$U�I?��'���퟼�I�pDXxPFg�(Į��I_3�Q��֟��Iџ|�'a�7-�ր��O0��ŰX�� "&G��P�،W�-&�\�쨭O �D�OܒO=ke�0fpQ�Ѩ��e�ЪR���ԧQ4f�Vl,��'`�l���<����.bv��I��$:N&����R��<��۟���̟�G���'f���ҍW�:���E0���C��'�p7MW�|;���O:�oZm�Ӽs@�Y$I��;c#ڿ2XrxɇD�<����?i�����4����^�%��O���AVE,��*����![<(�ӛ|�P��ٟ���ϟ�I��+�'�L�L��%x�=��b�jy�f��$m�OZ�d�O���\��ތt�v��6`H�-��D�%�4cW��'���)�>�zDsW`�ek�|8#��p�l�i5�I�uV˓d^�����O�AO>�)Ox�xQ��)x�z)Kg@b8�}9GC�O����OZ�$�O�I�<��i�~q���'
d��O�_�d�8V#ʠq0���'�6�<��9����O"�$�Oά3�C �L$؃F����3��@q�6� ?qc��9�D��V��߭���&RZ�C�%ߟB�|��4�u�h�I��I����I����#BǎV����@�˽R��1$ߪ�?A��?���ikD	S�O�r�j�>�O��w&S�>W�aa�Ɔ(^�rD) ���O^�4��a��o���el���B]&/�T�H�/�8�:�0ӥ\"3/��	X�	Xy�'K��'Z�'K�q�Q!t+�8+PJt��Q :#b�'��ɪ�M�ׂ�8��d�O&�'���)U_���	��X@��'�2��?��ʟu����n4����	#X��(��Q�+{�}Hq��* ��|�ׁ�O`�HJ>�t�K�{��ːg������?a���?���?�|2+OR-mZ��`!8��#Dt�Ŧ5UhdQ2*�4��
�M��ͪ>��NR⊙�'�<��3Ӟ�P`����?I�b�=�Ms�O���nK���L?�HB"B�'�^�2�V=aȌ�"�l��'���'{�'&��'�哜3~�9��!�8��aB�I�D�� Y�4S�����?������<Q���yW�^�
3�%� �N�k@���w2��)A)��7M��ɥ���!	���-Y	/Ű���#{����3
�[_�	sy��'E�FO�,+��6�ψ]��Q6�N�8>"�'�R�'Q�	��M�W��.�?���?af�W'�֬�4& �A|�i����'#���?�����za6E��H@&ڊ	ѦD0x($�'+��Ԅ�;�x���D�џP�R�',5�TI��@��U��Ȯ0������'���'B�'�>��$XL�RoРʀY�F,]+]�@�	��M��K0�?q�x4���4�x�P��C�R��6���W���>O|�$�<Q"��Mc�O(����Й�z�� tqh�
� }��#b웋�l�9um>�$�<���?Y���?���?)2�	/͈	��Ƙ1O��7`���d���]�1��}yR�'b�OfR�ƎMAdTS�"֩:�Z�"��0H~j��?����DC�xY�%�%�C�8�6���;�(�94B�P:��$�@8���'	B�%�4�'-�
ƨ��jƁ!돴y�P��'���'�����T\���4u��LB��`=��`�#�h T)��)=��̓}<����O}��'22�'��yB�ה"E�Tї!͡�����������R2�¶w��!�I������@��b����+��<.n<�R3O����Ol�D�O~���ON�?3'��8�0���7.�f:�N��I����۴b?\m̧�?)0�i��'2Jt2A��id�̸ �Z7ze.a��|�'%�O�n�ʇ�i�Ɍ�L �dL�{>�b C�I��9�u��L��0��<�'�?	��?1 g6\&�Mq�mJN�����_��?I����DĦŠ�![cy��'W�*xr�A�Ⴡ.R��[`�%IPX� �	ş���d�)rE'���('	(�9c-VtFX�"��L�� +O�	8�?A#%������A��	�dL���4H�d�Od��O���)�<�d�ixV�f�"jA�%�K�F��-	Í�l"��'��6�:������O���KՎ
X�P!JU�rj��:��OP���<|��7�/?��'X�X)��wj*˓)%`SF�]�� po�	�M����O��d�OJ�D�O����|�W��o^����1�"�ض��b���lŞ|�b�'�b��t�' �6=��\���G�z���6 �h<�(���O|�b>%�DEئy�_���9`f�l(�#����0�f�0��&�O��J>�(O����O�@A/ j��,I��/*��д�Ot���OX���<��i���z��'���'��q�@F4��x*��� 
�,!��$�S}�'��|b��\�XT�g 
h��LJ�`ĉ���@.�b���oш\1�t����\����%l� ���Y�N�XDГ��70�����O���O��:���b��	V\Y�H��P�(����?)P�'�^����?1��i�O�.�6���&g��p�DJ9���Or�D�O�]�mӨ�4� 1Bn����l�v&Q��E�B�����%H�����4�����OH���O��D�c�6�yC&51��E[��]!P.˓	���g?�"�'����'+H�jү��t���5'رz� �ʹ>����?�K>�|�T)�
{�Z1��+Z53������n4p���Tf~���j��I�L�'�剆@�6)¥��;��iF���:pJ!���L�	̟��i>y�'
�7-��8�<������������"�/�`0�$�a�?QbX���I����I'`°!rCI�,�SU/ʍC�Px[@#�¦��'5�B�HX�?�E����w����gF��\���ȃ�(�H�`�'x��'���'���'��1�.\%���k�����&9�?���?���i&�Y+�O��Kw�$�OfP#ʘ+]�fHX�lĎk�Z�hcm7�d�O��ԟ�@"u�i���� ^D]kg�؀t�@�sRl��=Tl2$F7vR��~�	vy�Ox��'���Աٖ�jb*�F�ԑ��2�'���"�M�M��?���?�-���3�N)��y ���u iS矟x�O`���O�O�SKz"��Ҡ�5���ԁ�0T�M��"%�:��*?ͧJ����E�\��h�\餽�@X����s��?����?y�Ş��$��?�(boJ��Bԑ$�Ӭ���h��� }�F�d�_}�'�,�A���e�]� M�[�����T��r�mզ��'�TQ��?��^�XȤIK���H4ꂬQ!�h1�w���'��']r�'p2�'k�S0qh��\ vl����Ss_��޴"yV�+���?����O��7=�b�s����|Ԭ�[& W�h�J4Ѧ+�OX�b>%�g��覽�?��02#HI�
�K�$ޡ0�θΓ3�����@�O�BI>�)OR�$�O@��pF-]&9ۇOۭq�0s�/�OJ�D�O����<���i�v�ɗ�'Y��'����lϯ3r������1���"���HV}��'��O��	���G<��C6e�H6�h���@��oJ;d������k��8e������
�E
c�at��yW�La��U�h�	ӟp��ݟ�G�T�'���'��6EhaCu��:�D���'H7�O�J���D�Oؕm�P�Ӽ��Dޏ|�B�ʠ\'*Z��O�<����?���HΙ��4��DJ�~,T�{�'|?�A���04p����bTe9��<�'�?Y���?)���?���/'�����-UW����������,A`r�'B2�)6$��T��L�$O��r�.F�BA�h�'���'5ɧ�O8H�sՃ#�U25���(�v����(ؙ�O��V���?�3E �d�<9%с>�"�j�)8L!; kG�?���?���?�'��d̦)[f�C��h�aE��j9b4c�1u��E�o�Ɵ�ش��'�6��?����?Ƀ�[�>����YSM�ҊZ>�JA(�4���K+B�$�����O}��۸V�l�R
ռ5Xt�E&���y��'���'U��'�b���$L� q牕^ ���ҁ.�,�d�O@�ĕꦝ�a}>I���MSM>�PG�&o�����L��Ji-k삵�䓪?i��|ƥ�0�M[�O6ԑ�� �U�憎i �'���b�;`���?�6 "�D�<ͧ�?����?91(
?.qM�w��<?ऺAa�&�?�����Φ��ǡ�Ey"�'4� ��A��%�\Y�f�)��[I����8�	`�)r�"*J�~�HX�VeA�f+��ڰO9h�����@�џ��|�e�+A�H�vg� �a�H1NyR�'Tb�'��^����4z��\K�eR#He�<�4�3I����/���?���6������l}��'��-sq�Ƥ?[�h3fCR;VC�!fU�������'�h��e��?�c�P�ہk�5|��t;wA���M/t�P�'�"�'�R�'�b�'���w��|����	N��h��TX޴QJyj��?�����?	D��yGEK!;*r�h���&JZ�B#)ŀx���'ɧ�O;Hӱi��I,eABuh�%�"�Z�z��JL��T�&[|< �'�'=�	ǟ�	�ı��k�,:$X�P`
u��	ٟT��ß��'^,6��-ʓ�?a0"L S�<"&e�	-%���E�H���'@���?!���_c���'cת����j�
�@��Pi'b�5P�&Un��'`�F����b+S�6�"�oJ>��7��x�	矈�	�hG�t�'¤�	B��W� ����(h����'?�7�\�<���Or@o�O�Ӽ�e�L5^�0�Ǥ� &�� I�N��<���?q�HL�� �4���I>@z�3�Of�䒁�I�PJ��s�P+���Q��|"T�������	۟x�	��4�&Β.r	j����%_�:�Aw	�Py��j��Bǁ�O��$�O@�?1UF�*m�D��kJ�v7�:#g.��D�O�7���6��1���<DC%(���n�v�d��O��<'���'L��� &,��"^�~�8�3$�'j��'o�����W�T�޴x5Jz�� �0�Q·'a��駡M�10P���N⛦��x}��'���'+8#�ȅN0���BG!o��K���������Q�,�����	����:��e������g'��ȕ6O���O6���O��d�O��?�j@d�I�H�Z�v�� �l����IٴBz��'�?I�i�'8����B���x{wa����@ɢ�|r�'��O�:�葶i��I=hR��=��qs`�ޜ�L��ȥ���2���<���?1��?��&�O���y@*<A�l�'(P��?�������f`���������O��$��=*n<�e
wzD��O���'x��'cɧ�	���Ł��%3�F�U�L'(�2XA ���Xb#���S�(bF�H���
�����J�jx�bS���)�I��(�	П��)�Gy�aӼ�8�#�'v�n-a&!�A��9����#>���OlTm�t��fW����4k@CőXau���˲"�mh��M�<�I�r�.tm�t~�$VF��4�J�)�	b�0��C�Z|&���T5LR�d�<����?Y���?���?�-��y��KR�zq��y���;Z�hT�tm�ܦ��BNԟ@�IΟp'?M�ɳ�Mϻ`V̀p��P�O�!�"�Ҏcf�
��?�L>�|��F�M۝'�0U* G�CF|+'�^�'�A�'r�1%��{"�|rU�L�I�Q$fUh��Ŋt�W�'f��CGZٟ���$�	wy��V���k�<I�[0��F�@���*V���a ���>����?�J>i2��8[e>���;��q��~f�5w��aǓ��O���	uL�f�8Ĭy�
 	i)�Xyf�ܩr/�'���'A���۟�@���n�D���\5�=0���͟`�ߴ@�U���?	��i�O��(j��u�܏J��H�A w��O��$�O��)��s�0�4��t�ǥ?�Aq��-=�5�� u��N�Ay��'Zr�'+b�'RFʄ(���2��.��xP���@*�ɐ�M�u/�:�?q���?�K~z�2W���ԅ1x�l!�֜>�z�TU���	���%�b>=�`K���2,[�2���9��,7���Ka�)?�s�Z\oB��������D@&%�P�X��eDD 2r�٥ �<�$�O����O�4�l������f �I�����Bvʟ"\xF��H�B�x�J㟼:�O����O8�č-"h�����-�4��O$rr����u���=}0��s���4�>���~b$����n�:P�T�C0pOt�I�����˟��	؟8�	i��)\S勑�wP�F�-0��j��?!�vH�f�H����'6�<��'\ ��q� 0P$���1O��D�OX���}r�6����< N�2���&
��ݛF晫�,�!�G^/BN҉�o�Iny��'���'���T�;�T@փ�?7�6UIa�$:���'�	�M;⍄�?���?�+� ���+ۮ#�� i� s�hy����R�O���O��O���	ȚᚂN�1'� s��^�6 ����uS���b+?�'���Ė��`��� ��,G.pI��̺*�b!����?a��?a�S�'��d_�)rAmE�~�i�D.J�-�p\kC��T�Tt�'�6�;�	�����O�1@��F�\j]�`dƷ7&��QU.�On�d��
4Z7m&?��qBU���2&�L9dp�)�8��5���>��ϓ���O��D�O��D�O8��|�P 1m��E�.WB����N�9)�& �5m��'�R������;A�Tĩd>R٢��
E�9�I���&�b>e#1m
�u�S�? �iso�>*�l����>�Q��;O���G��?��<�$�<�O����CND|k#��n�����o����162�'��O�/�.�Ir�T�d�`S����s��O�|�'Cr�'f�'�p�1�6@RL`��� =|�5R�O����Z?Ŏ\;�C9�Iؿ�?i�c�O��˕
7�l;Tk�4�$�5"OH|��n:r7H��
²&`}	U	�O�o�s�VU���|�ڴ���y�j��o h�5N:���cf)I�y��'SB�'�F��i�I�5��	B�ԟLA'��gbP)��P�,��QJ��=��<q���>+>��Y�m�4y֌�KC�ɽ�M��O��?����?!���VU��D&V�q2�A�D��l��?�����ŞC��e�Qf�rY$K$�V0#����M��Z���,X$-��<��<�hC?� Tc�`��+�l�Fd�~��IٴW�$�3��7#�q2f�K�
!^T���
{~D�c�D���d�Q}R�'6��'�@�b�j�q�v��Ӊ�=�,��n,�v���� F�2��T@�j�S��M2�K��T��k��
�X;���Ro�|��I�?;���Ճ��O�xh0�	2,����ߟ��I��M��W\���s�@�Of�8s� �D�1w֕s����)&��O �4��kPCh�D�"Na�G�)ZD�kD��F�%2g�My��	q�	fyR�dl20���٩P�����͡C��XYݴi��q���?����򉎏!<|�[f�M�@��	�P�	����O(��7��?���/�3��+����]��L;h��y5BԦa (O�)Y��~Ҕ|��N�`i�m�t��1y���:��Np��'<��'���\����4	
X����X.���e�<��Ч�¼�?���{\�����W}��'{������'=���(�$8���ѷ�'���F''�V��4��M�6��)�<ya���\��dE��sw��g��<�-O��d�O���O
�D�O�˧(?t�:!�(} �S`M�G|[3�i�$t
��'d2�'T�O`B'`��.ͣ0:����\إ�S��2��$�OT�O1�f���ad�x�ɴMd����&yC�Q���X!��	*M/�|�w�O��O���?Y�6�څpLM�^0�IC�`ߴ$X�Y��?���?a+O�o�8hӦU��۟��*[L~�-�����aVcë	[�?�Q�$��ʟ�%�X���W�Qk��[4�W)L��P�P�/?�h�j��y�ݴ5�O�0-���?��o۬ 1 �k"��+O�@��1nW��?Y��?����?���i�O�a�%��״�xf)�>?3�(�$"�OP\m�2g�.���ܟx��4���yg
ٵ��9�#A�?T�K4mO)�y�'���'��ً�i0�	U��ڟ^�YeJ
�Rs�@Ȱ�9T�>����,�d�<9���?���?���?y4�֌A�E���P�~�@0sM�����٦u+���꟔����%?��ɹ"*];3 �^�|�J��آ2� p8�O��D�O�O1��ax����v�!��_Ҩ�ha��	f��7��\yR%D[�L ������8q�sV�śp�����ڊRɠ��O�D�O��4�8�4��o�'d���3�f�$��*�h|J����]�b$fӎ����O�$�O��d_�H����jM�'�ܑ��j�8.������j�x�y�8�z���?�$?��ݹZ����w$W4���'X d�蟈�	�8������	@���]Q� \jD`��1e�H���?������������'C 6-'� �Mk���j3Y��=0��R�A��O"���O��ܴ$��6�:?	@d�<B�IB�Y8L��ݨ� hѣ���$���'82�'��'0h)��گY9�a��/�D!(��'��P�lٴUb�����?�����$�fmQ!)YB�����f�4a@�����d�O��$6��?i:PI�8e����#�!�fH���Ŧ�d(�����1r.O��|~�&�4"��Y��1�O�+�2x�ѩ#��Bٴ7��ܺE��o2���`�
5���;#��-�?���f�6��C}r�'SLeK�A��|�-I��	���"2�'���{@�v��|�d�fO���<�G-� .p�`�M� ���0F�<	*O�����`�QH4�N�p� FE��S~�o�/I������|�	c��t$��w� %��E�O��L�6n� elݹ��'��|�����ʛ&2Or$q#�
W���I���(S`�[�2Oꨠ���?�2%?���<�/O�Tg@�� \l����x��B��'�7�Ğv���$�O���5:ة�p�O�p���r@���qY��<��OX���O��O�0*��H�,�d��Z�T�&u�s����/�,x�l���R��Iџh�3l�=*�H��^+�|A07$$D�Soԋd�jѓf	�vBE�E�p(�4~2�()��?��i�O�n�1�(p�A�Y�$���OOl^��O���O�(9Dw�J�H��s��?��d΀�.������t��m
BGn�y��'���'�"�'��9�xsF�òE�޸�� )w�3�MCcaԭ�?����?�O~���W�4zr-љy*~��V��y���\���	ğ$$�b>e#�L0� �!��B�l{����Js�����
2K8�I��>9�S�'�p�$�4�'��e)C�߼:}�����I�B��5�'jb�'i����TU�LQ�4!A"њ��f��r��'�ZHI$eL�6��b��L˛��DLr}��'��'+��ڱ�WQ�D13L�1���J��6�����JT�ޏ0��)#�	��T�fH�h�KF��e�E�4Ov���OT���O,���O��?�b�#��n��@�X
2��0)��� ���H@�4"%@�O8.6m"���"lnX�x���]����%��_o:�O��$�O�ɗ�	�7�5?���B�2�G)��C�ҵB�B��I �T���8'�D�'��'W��'�29�BEӿX��! k̶
֦����'�^���۴*yj]�(O|���|����7o�p�˷i�Żc@�p~RE�>���?aK>�O����&ݳ/B���c+w�0Ex�K�_�^i�úi����|"�ʻ��$�������5p�R#�Pw¡�Vݟ��	����Iڟb>ŕ'
06-��*����$Ȱ`�dr#K��F��r���O������?Y�Y���FiP=�#BZ-x:}(��T�$�r��Iß�bY���'���*�O
)O��2�	�a�6Ts��w��hv9O���?���?���?����	K�rm�����q��L�^��s$&k����O�O����O�����D����q8�e ��ԥ��e��n���IޟL&�b>��II¦�͓!�45���!%Fh��D�H`1ϓAX�r$�O�$XH>�*O�I�O�9갌�Jr��TI�+��+A��O�$�O�ı<��i(t��'���'�&{�EQ�n�6���fu8f�_l}��'oR�|")� zW�X҅ɍ=^ ��ߤ��D�zd�SU/U�L�1�@�{��I�&�d� �Ę�O��c�ö�}	��D�Ot���O�D'�'�?�4nW�j�L�5��� AX7�S��?)g�il��R��	ߴ���ygj�:�:�ze��,n��[� �y��'��ɯx�
|lX~�I
���S�:��-Q�*�Rb����A�������|�Q��������ϟ �	� ��fR1g$l���tjNd��Kuy.k�@t�g��O����O����D�3�xdi���Q*j�2H�'����s���p�
�Dn�D��?k� �!N�e�0ʓ*��!p#��O���J>A+O�E�� �(��|�ǛoJ��L�O����O���O�	�<9&�i(��PV�'J�,s��_=؞᳣
U0y��X��'��7M:����D�O��MTbY�畧t�M(W�R�J��@y'ʇ��M[�O(����R�)4������,[?�\����0���3O��d�O�d�O*�d�OZ�?U3�Ϛwm��Y�LK�M;(���D�����ݟ�ݴU����'�?9��i�'��������҂�!z/:���y��'��I�"_D�l�P~R �YM�\ �9�,QR��r����ğ���|rT�(�Iԟ ��؟���	S��e��L=�ي���� �	ay¨g�p�#P��O���O|�'oo�A��OBK�f�%N��:K��'m���?�ʟՁ&�ΓNS����B�� ��QsBܤ:�z;���|"S�O����H���x����V�`�3H�"�D��5�%��H���!�l�@C��Wwf�)��B*��z�M���К���?;�j�Jg�7ze�jF�q�d�ٓ'HM�l���*�HO���ιm5�ș�$�%B�8�2>�l(�!��ȷ(�*y�(��ɋ�B85��S5)H���P��!}����'�!�ƅ2�#�99����(�'BP(�r�H��r�(�bWΓ�C�
��ET#a�\)���)x��Tʋ�n
���u��B��}K4(�w��%;�n�	#3<$���#����3��4*���'�����&�d����x��� L��,P�kR9���bb�Μ]��&�h�	ן\��By�bh��	w>�P�ř�I �O	�K�^l�-uӾʓ�?M>��?����~�K��&�̳��ŀsJ2�����d�Oj���O2ʓ9y��XG^?u�ɝ&�P�����b5�zGD+/5T����$�P����\��LaܓtlpZ�ᇔi� �LF�2�lП��I@y�ꇞ6�>맂?)��b�	[=��� 'C���`dH9�'7B�'^Z�Z��$�?u��
��@g�H怟
jż�zU�`�X�_�rU�ѵit��'f��O������Q�a��s��� �c��9��������X����OW�Y��FN4��	�4_��} �i&��[��s�r�D�O�韄p�'���);��W��":2.ܐ��Y,�\���4^��y�����O�k��F64:��8��τ`0� X즵�I՟<͓� ��O�ʓ�?Y�'p���f�1]L��q�GYA�$�ܴ��u�`L>���?���f�P��}COX�gu���̦I���)ЯO���?II>�1 �`q��cW� aXcCO��bh�'<�����' �	���	����'0�y��cLT�Ȕq@`C�<���r� U���꓀�$�O��O���O��P����T�~9����~~�թ��WTᲒO��$�O��ķ<����*2�L!h���hC�R���:��R�\͛V]���	a�	۟���;~�v����K0R�@&ղB�����b �<��O���O��Ĺ<Y�#I�����*˯r$�5�#�QG�%2���M���䓆?��pD�>�U`b@�1e�&R��	������1�Iʟȗ'�@"0a'�i�O����lࣵ�ԑx���f��O(�@Pu�x�]������$?�i�� ֡��g�8Fg��aD.�
DHmCu�i��.�V\:�4Z����8����DF�i�xպCj^'��L(��ԑ%n�&]�4���qK|jJ~nځ/����OёZ��1�	�	6�GQ�$nΟt��Ɵ��S,���|z�O?2�n|��R�)0'M�jۛv�'�2�'�ɧ�9O���˭7�,�[�m@���T�l�g���m���	џl:������|����~2��:?�F0 gD�2~P|Q��V�M3������3?����~rm>,��e���=tG�`�tR��M���0mdx�/O�e�O �O�aa�mʹM�(��!,�n�HP��+�D≑m"�b����]y�'ӄlHƅ�gvh���Ԉ'�
���d]���	C���?i�'Q����#�=�����  �H�2u�ݴiʊ��<9������O@0���?�j��i|�mz�DH1 5/m����'y���Oʓ;m�HnZ�7�4��'�σ2�~��3�@h1H��?���?�)O�KA�O��5E+a�5\��p�EE�E���h��p�^�D1��<�'�?)L?��p��G���X��
�t�!&hm�`���O���&ex����'��\cβh���f�E
� (a(��M<�,O����O���������������X�Ļ� �>���4������?!��?��'���T%	���b̚8Rpx"eS��i R\�|8��$�S�S=^u
qY���+B~x�Q���NI7�X=*�lZҟ��	ҟ��s�O�N�C�ne�&�J�@x�a��Jw���m������\%���<��Ytq��Y�6��q
�����s�i��'!�.68��O��f�OT��T)L`�, �)?}Pտi)��|b��~��?���?��%���AC���Q0_/����'�7+�d�i>	��v�B#��Ӄ��<�R�ӂ�G� ��-�O<�����?q/O���G����!lS#|�B��c� ?-$�S��<���?����'��䖨S4�+DF	1cE85�Bɚ+����U��$�O���O�t,གG8�ڐA���d�2���C�8X�Υ��V�$�����&� ���4�'#^�9u�Ī>��#&G�c�u��j*�D�O^��?Ѣ�[����O����Q.2���u$@�xĤ�bA�Ϧ%�?����ğ3�'�A�r�X6U�dDP! �N�H�9�4�?�,O&�d��$ɢʧ�?������ph�lxvA��&����}�>�'�H�	wy��O��R]�t�� ub`��GI;\����H��&����������?��u���*6�<�� )W�K;������MS���dR;Y��Af�G�9�Pt{u	Y�i�*��'�iz|l�ky���D�O��D� '��2CD=:�l¬]M �
��Ik��K�4�?���?�I>��y�'���F�*�L ��)�-,>��
�d����O>���I@�$�����K��0q��Q@����%�4��ulZџ8&�먟��O����O�0)����Kp�)X.B&{9yǬB��9�	YM���L<�'�?�O>i�E�s"��	��ѫX����bs��'�BW����П�I]ybE��M�$H2֦Y��T�Pw(�<K�>1�� "���OT��!��<�;f�2%�C�/4�����M�P��8nZ�$�'W�'��\����/�����%P�1j\�QA�)?����؜�M�(O��$�<���?1�~�$��
c���c�-K�Hv�؂{IZ}��V���I����I]y���!ꧾ?��#%Yg"����b�����CK�]}�6�'m�Iޟ�����\�хg�ĕ'���1ƕ-Pu�A�T�Q�hR�Y7aӄ��O��m!��X�Z?1�Iڟ���Wy�)�L	:Ĕ��$��$z�O����O"��άw`�IYy�؟T�ӡDțm��q�j]�F|�Ʒi;�	��h���4�?���?��'	�i�]؇H�*������Q�8�5Lp����Ov��B8O�	��y"�i��|' �t�Ӧ^����E@f��Ac1�6��O����O@�)�]}�U�;Q�B	�� ��'�����G��Mc����<�H>1����'oL\#�Kюwq���Ƌ2!R���b�<�$�O��DT)=��\�'q����|��e(�kS=mLl�� ��sO,XlZ��d�'�$�����O��d�O�e���K�B����F ��f�`�æq�ɡP�
@�O���?(O���Ɗ
wjF�<\����X�<p{�Y���f�Ė'�b�'Y�O�f�;Ajԙo���.E�Tƨ�����*\@����O�ʓ�?9���?�FJ߄�bX� ℗�| ��f~�]��?���?!���?�(OT���D�|"t,�8"O�x�r�'�*H�F����	�'IbP��IП �I�Nƈ�	�qFE�!���'J4�b �-��1�O����O0���<�f��2R�S��@�1��
�yनܷ3/F��2ŉ�M�����D�OF���Ox��W:OB���Y`,,e$E�G��1�J2��h�:���O�ʓYmH(A�V?��	����5�����'˾iΈ�HQfF�Z�ڮO����Oh�X0)��D�|Z�����l�74��=C�V�caH�s��J��M�.Oȸ�QbB�������8�	�?�s�O��7���@D��A��L�ui���'RI
<�yҞ|��� ^� ���i�r��_�V����7-�O����O��i�}U����J���ӄ��:� ℎ��MSсD�<�I>q��4�'Nn� R��s N2n=��Y8i��i�iNB�'T"��1U����d�O��	&lz����ǵ"�E�t6�-��F�W&�?�����p��}���ᑫ�
	I2���ao�ҟ�j`�[��ē�?�������/�T�pc(OL�qrƊ�}}"o��yrX�(�	�%?��V*Ɣ|8���8&窰�W@όl�`�BH<I��?�M>A���?i���$����	ĳ.>Ȣ%ԫ)�V�H����$�O����O(�=޹�u=��$h FO�e�D� ��K���xb�'
�'r�'��`��'	���R�U?6�z��¨+T.QP�#�>���?�����Xȸ&>�r%/�?�PiCM���֢���M������?��'x�j�{RB�.:�P��q^�F"��VF���M��?.OviY3F�]��ٟ���*:�:�����c���@�L�c�̛I<���?Q���?	M>��OER�0(�s+V�!�%,Ġ��4��d��/Hh%mz�Os2�OL����2!�][�*Xۀ̎1�Fdo�����	4$��	I�	Eܧo�����/^�{K��Rԋ�?�o�n���pٴ�?)���?A��j-�O��J�%�	�8q�)WnX�3R ����"@��$� ����3'�ё��'@,,T�D�0F�L�3�i��'�B��\� O<���O>�	$� Ab6 �2M$��)֭��6M7��G6aF��%>!��ڟL�I.H�z��0-�����S�{���Rڴ�?��d� D[�O��$3���°*�Né4ʽ�]�m�:���R��s$��h�'���'��O`�'C�@�޴�O�G���p��|�rc����v�џ��ɸ4,R����oA��V��)�,��1�����'^"�'��V�������4���N�C��1��DX���d�OJ� �D�OH��9|���ʍcų�%��tmb����])N�LH�'?��'�rR�D��M��ħG�h��0e�1KS,]� f�i[W���	�h��TF
�o��X50Q��I�f߉0|��%��u|���'kV���"��'�?a�'8Q�\25)��@1��:�Ė�l��!&���	ʟ�ASg~�&����
�8Eے�>Qv� �̀�`0mZgyr�� 0� 6�S���'/�de ?���R `������"��,��IΦY�	�����"Z����OIX\h�OJy�����m{�`��4P�JM��i��'�O/�O2�$B�|c�-,L�H9�̲m��dlZ+���?���$�'�P3��01hr��Ɨ'uV�`� S�'i2�'�l%h`g �4�8�'��=8��:px�hA��<���ߴ��'���f��O.���oml�.�tdH��c]"yt\o���J`����|���A����`hY��\#6�X/b4�'rY� ��ȟ���ey2@S�H����b�ԗuX����X�lk:`��#-���O���Oʓ�?Y�U�%����8S�`��e�V��t3 �[d��?����?9-O�p��]�|:� ˟dp����ř<<l�M�U��A�'�b]�D�	����	.Uc�����b��8���g�63� ��'���'�Q��R%���)�O��Z���)>�6Tb�M�t�Q;1h�Ц��	Byr�'z��'H��'�哱SrR�	�˜9��	3r���c;�| �4�?9����5�:��O���'E�T&�/S����#C�	"ՅA
zwl��?��?Q ��<�+Oj���?q�p�C{ݬ	�N3<�
$+z��ʓ#;
�f�i���'�r�O:��Ӻ��� ux1����>2�{�ئ�I{tw������"��Gv�� �,m\��a��H��6�4�f�lڟ����Ӳ����<q�$����f��:I�t���ȡP�O��y�'�F���?y�	� ]�����Ɏ�5ڲ�3�'E�'ӛ��'?��'v���r�>�)O.�����H0#��{���6��$�8r��x�v�$�O���˴P�?���ҟ����d�B ��-��O��	�&&�Y�|�ߴ�?d�5=���Ny2�'i�Ο�����8׆Ӽ1��	1�$d���: �����Ot���OJ��t���o�S p��������af�U��	gyr�'��I矐��՟\�E��
?���٨_-|`���Q*)Γ��d�O����O����OdȪ7i�OV��@�˄��
W�Ўn�f�xR��Φa�	�����H�I����'����۴t�� �̱~Īer���UF��'[��';"R����X�ħl�����=xԥp3�Ť%,"-A�iR2�'o�OIy���
)FpI�.J h��tBX�z��6�'e�'�B(U+R��'"�'�����`).T�Ǣ Vp�X2�"D|$O��D�<��NA��u׺q����Ea��Z�$g�� L��v�'�Bl��"�'���'��D�'�Zc;R��ǲ�d0�4�B?p��Sܴ�?Q.O|��)�)�

�a{Ŭ��|���o�*-�6�Ȩl �7��O����O��	s�i>���A��z{�=��͝Bc䰫r؛�Mۧ�'��'���y��'����$�:L�F���̥UH���1�o����<��	���d�<����~�a�i��W�^ Zb�m�9B"#<ɰ��T�'�B�'}��ⷡ�46-������P���o�4�DQ خ��>Y�����sB5_q���c@�,�N�1��W}"���'"B�'mbZ�hr
� �u���?�� �[�iǼ d���O��D#�D�O��Y�31 EC��5�je����s|f�`���O���O*�@0����2���bg��7\R�A�ɨC�f%��x��'��'n��'ۘy��O�m;Ԣ+�<�r%�K3&��Q��Y�\���T�I�����|�H��Iӟ@�ɠ�͉5G�%K	6dc3�C�Q�q��4�?1L>�������$6�'u(�c���q��qy¯Ly�j-�ߴ�?y�����,��&>��	�?�c�mߤ�%b,�6/}�aW$%�M��2b�5��.��i)�ȸ�i�3Ċ����܏pI�1ٴ�?���j������?���?)�����;�l�!|H\mEa=7ڞ$��i��_�D*�&�S��J��\A��b�� ���*l7�<8��pm���Iʟ����ē�?!�ԩi��ƍ"���lɃ���"	�O>�I�4ϸQqs�E�%{�	c�k��A��8�ݴ�?����?�����O�������6��l�����\�dT xA�7�ɲ�b���I������>�Ą�v��g�Yx��̍�zL��4�?yD�"wl�O���?���&�(�A΋	�Ε�K�k��hvS����<�I�����X�']�ՍW4�F��t�����x��	]%~c���M���� ��0W\�pa*�zpd���k8ҩY��=�I�"�"�	r��i�����d�UP����A�.��0���Ӎ)�(�S%� Q�x,���ۖk�C�3fM�%Ǥ愉�B��#$��$(�	����ؐ˯68��-ƐX��x����rP(��L��,E�҈[�HHҮ�H��+pJQ�%� 1�V̍����i7�A�8���9Q�g���	Q��|�\8�'*H�?�Y%�8�dL��v��t��oE\Y-
����&`Jh�S���
hq���Za�-KQ
����R�[\��CR��'-�i[##�="�I��T�*B�vj*�̉��C�p�4lA��?K��[�>Yp�M�5��´��!&�`���4 k��m���<d�ҝb��J
%NL���Q8��#�$�OD�}���M���cb��xTK�,2Ĭp��g��S���a��B�@�0*K����I��HO���@;8A�x��j�;,�Sg.}��'f���@�d���'A��'��w,����*�%�g�� S� �+��&Htp�Cd�O�����ߥ21��'Z���#+ �!�,8k
ޱ�N�;SG��� Q�+�O@�j�	Y�����RD���
�a߀��CC�Uz������dF/��O�ўpp�"!�h1a..,ތ��%D�T���W.��L�	�}�m	0�!?a��)*Or�Q��ٖ	�:�p��1��x藯�9!!��Z��O0��Oz��������?��O�ZT������ �Ĉ�he�؉��~��B�ɜp"N���Hۦ0r�M�(`2$C��¹(�,�&��8�Xj4j؞����-ê�&��(r�X+��)�`���Op�=�"݁ ;�a`�,ٞ6�̚�Z=�yb�^���Ek�aKZ=���"J�*Θ'�j��������lZꟌ��t��p4�-D�<�2 j�2Q���<y������	�|J�e����&�|���U<,8���=9E^tC��#O�Mѣ��.1����2hT����k��xB@F��?�I>Ae���uc!��V^Ę �Ν4�!��d�������z	�h0�=\�!����m�CG�<9���hD�3����B.扟{�ع��4�?1���i�59Qr�5"#&DFIܯy���C��F8^�2�'�JA��'(1O�3?���	�{��L�⥉�/+D�s��Qg�$�;��?eó望Hz ���KpM1�	-}R5�?�y��$�-Z���з'�ft|��Dg���y2CÊL��k�\?a2IX�] �0<Q��	kw�Hæj��<��Q��YO��ڴ�?q���?��(B/"Q }���?��y�;E�&)�g�bE��C�/.B��l1�	�g���U�|e��ò�AzDs�cѨ�qO,���'M����2���3q�ž' (P�$ſ'��L>�7�B?�N���Q�`Q��@�)�~�<��f��^6�e8AȪ/(�A���x~��=�S�O(.Ѱg˃�^�ŁTi�FJ���l�=V�0���'���'���s���I����'B������ۇR�jy�u�;�h��na<�Rm�X$"X�q���F�����A�A����[ "ljkE�6?c"+�
�$9_.>��!�O�8f�\��ֱn�6 d�	s�)D�\��mߗb��I�v���f��('��9��'L���T�l��D�O�l�P쒊xR��4GڏAF` ��O�	�2s��$�O��S(��;��q�����G��ʕ���?��x2gr�d��Q#`)��l�U��UHvA��p<���B�`&�� xE�я�]E���oRZ(p�s�"Op��6��s�hP[���$E�4��O�nZ��q��S0�Urd�&%^^c��*2���Ms��?�˟��z��'ʬm���f���)&hO<J�	�'��kW�T���T>��H���#/l�P+�j>(�)�OV���)�ӈ�<�;��A�P�(���F�.��'��Q��ۘ��O>��2ˇ4K��e�t�E=�X��'r�eq`��6{���\75�u�Ó$葞�F�E/��X ��P&̙��C�)�M���?���o�D Ed���?y��?y�����a�@�����`���I��'V�9�ϓX-��!ܾІ�E��<5Z��=�PNYGx�Q�-��L�%��M*Ya�FHQR̓]q�)�3�d��T��h�T1Q�r]�4��;�!��U%_d4��r��X����&ɍi~�ɢ�HO>��4	�/g	��0��W$Ѣ���h�
�B�o�̟8�I� ̓�u��'��<�.�K�K"M��xs mUYR�X'fɯ[�!��9{&@9�M��b�ܳ�@s^%ON)�MOy�blTҎm�
f�п���'�xa�&J��V)���Yz!C	�''��R-�,@��cA�2%d��{�y�H9�	�~�~$Zڴ�?��v��b�&{�RLh�J�;�b8���y���?������=�?9O>�voǁI�����N?;�6���	F8��A�,�I������^�bz��zBB���d�2x���|H�Ġ�@H�r�`Q��Y��y%w�q�!�(}8�5AB!F4�x2bj�@���\$C+�<�$;r�`q�dŤev�n�����Y�Tj�%�?9P��( ��c&�9%l0 G���?�>&�)r������p	&e�	\.8�*&}�h2�7}�X+�O�L�����A1���=!T�l��>�"DSΟd�<�j7c�=G��#�ʓ�dnY��aW^�<�.�"����8 �qWDR�������iO��``�)L@�ʲ씂N���'���'��qѢ��'���'�r��y�G:cHH�WM]�nލ���6-޲$�c�o�}����qC����|���>i$�|��B�=7a�S�[%�rm���=b��p��-�d�P��L>��`D	�D�J�F�@X~����E��?!�O����|����@�N�||ʡ�Bi}���юd!��B0^	$)���=qplL9��ST����HO��sy�R�L|���㇌Aўa1"W�m�|q��GO�;��'mr>O��ݟ�I�|�7�#j�F���Y�e9��9  ńY������I��['/��q�*=p͎�}�"���Wf<ag/�)}zp�5�Fs��`
�A~�\�	t����qj�by�d��4*�0� D�`��2=,�AQ�R!ODX�sѪ(扞��'~�j�|�����OR)�0�D"o����t�=�]� ��Oj�I4�x���O瓳X�`��7�d�z�a��L<� ��啟��x�-����'Xfe����cHy6�F7{�4��Ǔ4��%�	J�I�}�� ��/�����i���62S�C䉽.���A���"Ĭ��#Z�DL�C�I�M{����@N~ seĨ>��3^m�%[�p#�iD�'K�ә�����}�,G��:^�� �d��.E����O���f��Ob��g~�Mʕ'~֐:���;9��K�����@J#<����UK&���E/1���[�CO�DÊ^f2���� |F��Y���)��/��KX!�� 4�򕆖�m�����-W9DaxR)�S����QC���Gв|�0!5�i�B�'��Ĺ���A�'���'���w�c0!/͠4�sOM����󤅊/z�y� �;ovR$2��͐:�� rG̴��'/N���3�l�I�W:
����
O���J�y�I
�?�}&�\�w��iq��z�j�tI�X��4D���$�q��@va�[��-�� ?y��)§*� �`���p����23�ak������?���y¾�6���O��SB,ȍ��ZZ[Ѝ��XYP�<020��a#�R?q
�:EL�z�l��F��6��C��> q���6 �F�Q&�@%�ū���O���� p�����z�xq�6�^��J��"O��bω�	>j����(w�p� ��UW�U�4�iŽi�R�'�)*K7}�������J�
���'��$�$���'=��,K�R�|���AK��тY#\����fZ��p<qt�IR����!��m��c�`	`�DY��\��	�g��d!���)�ب0j�?23��qpF�r�!��\��͚Bl�xzdk#ţW!�$��Q#��C2�SQ�G�B`g�%扴rQ�h
۴�?!�����L8���K7^�h��7vl�	]��b�'K�� �'�1O�3?!�ώ����'�A�YŘr��t��?Yc�ߥi�A��ߒX�(����3}�N׿�?!�y���g�$IV�"6�C2u�|��3g�4�y��ϼs�n\QQ$&p��Pe���0<�鉡`�>0��"1��2'Æ,G"�ڴ�?Y��?�-� CF|0��?����y�;2�����6E<��"E�H*LԘ�y2)E��<Q��8��afl	�HӸ���$O`�J�Ԅ��qD$`�ѫ�� �[bA�� �4�<a"A�џ�>�O6=��۬Y�qa�J]b=��"O���֎��c܌|H&@�5�Ը2�������5`/���7o[;zy����iT~h�9��ԉ|����۟����<�[w�R�'L�	�4e�ZIɰ�R�]z�#v)ךZ��J�O����ؑ]P`Q�NܴU 6�[�G�4!�Dؐ]>@����D<%�,y�.�*�L�à�'/��%U&BB!��n�'�<=ؠG���y"�2��p���!�F� d���'|�b��P*���M[���?!�`�)�+��D�6`��
h�9�?a�'ϢU2���?��OUX�
����3_Ҵ`�2&�V0Jt��g�>l��	�g�P� 	a��iִ��t �\��3�;O�I�2�'��'��	[ҧO58�NX���L�z܆|!�'����3JL'5�8��ڃ(p����'7-ȓ	�QcLB+~��X`	Mx1O����K�)������O���Y�k86��� A�e �0B�#)"���?�vĂ�?y�y*��ɵS&���@KE��jq	�|y�'�������S�b
0�G�TO�;H׷)��'�����o�S��ᰄ�F���
Y��AUq7���d�<l�ċ� �-i7��?l�%��'�HO�W�m����nL;	D�����Ц���ҟL�Iw��)R��ϟX���������B`���/�=
P�ن=�n��E�l�ݶ9�牀?b(�v�9��ݐ��!]�x�ԒAM<<O��{4B��crm���d1��.�I�����|R�� ��hx'CU{T,�$��?�y�a�M����	��P�F%k4�ݵ����}���Xa���_<�����b�4e�׊H3�ѐ���OF���O���캣���?��O7�}a��	�0�R�3'"��k����x�����b�@���Lit�7J��	x
�'���zgI�yl�h �ڏ[�r$�aݢ�?��3�LL[�`�]��H�g$M��m��P��a� ��ZHB���Ϝ�Ѥ��<q���I2n�ȟ����2yF=
�i@|�@���μGRY���<���������|2Q�M���'�S6E� I��9�mC�AH��$@-O����$^.g܀�#�
���I��e.�xr�̎�?�N>�үN_,�tSq��9.��)�A��l�<!%�@�c���6A�(�s��c<�ֺiJ��1n@B�r�o����юy���7-�O��$%��HП�ڂ]H������5ipxf%���	�}����IG�S��Oި1Q�U�1�~(�1��Fȋ��Q��ɔ'��?ŻDl��=��;�ET#��{��*}����?�y��d��6A��� �4>�����y�l]'eHN1q��[�;�L ʧI��0<���I �n�[d�X�Xް���ݭI�:�4�?I���?��ߓ@�,�:���?a���y��oa���u�	����̜�<�����y�(����<鳦��|������ϘO�TbծEFܓ,!�!��	�����T�3S� �S�	��<��	ǟ�>�OT��GoR:#SlRc�94�*�(e"O� rxSb0W�$�A]�s� L�ѓ�T����Ӥ)=�m��+��sW�J�4�Tz�^�����I��h�I�<]w�2�'��	ٛMFT��֤_�>aD��gϟ�p�8�H!O���fP�cN.��M�7u� a
P�!��P�c���CE�ѲzV�m(6�ІwK�H�7�'����H�:/X�'G<�R=�5\��yb$,�n�0�����,�1�K��'n`c��+�e��M����?�@D�.Z.��h�SQ�\iسa���?!��J��p��?əOh.t�������0�B}�♒wvD�#�����W&yXRH=�D�8����];g�xR�ÒOv�x��$�?Q���?���n��}x�`�.Fk@�G%�6L�.O��<�)�',=�,�Y��i�PgZ$���S�E��.�#q��z�H�	�y�Y�`TDA��M����?A-���Ygf�O�)!A'"�@�6�� |�����Or�/V�P��8�|�'	Ȅ�V��ň�L�ʞ��M�J�"5�S��=�c#E�f>"0�!N?y�P�OrT
 �'�1O񟰵�a�<.k�|� N�LM��R"O8��eƟ����9����?�����'�#=��Ԥ\�x�Pf#	E����p�e�<Q�
Ͽ&�j��hS��A�JH[�<IE�Y7]'�<�#ꕄ{���'��@�<1��vA��8�>e�D���DJy�<����� ,�����(F�4Ɣu�<� [�q쎝�0ǚ'��y�q�<)��عkp���hYi�N��v
�D�<Q�LY�< ,9#��#D�-<�TB�ɷL�^=��%�%)-��FIZ�Xz6B䉁~x�j7%?G�$ W�ԙ_�FB�Q�^�R#�w۴Y��a��Q�
B�'Qz� ��"p�ppɲfVOgB�	���ɱP�6�A��^"��C�	D6�[q��^�f�G$���C䉿�[��I�*��x2c�&m�C�Ɋ>r���0_��c�̜o��C�I�Y3h���n�,Z/�	*�I�H�C�ɝf����R)θ|VZti���p2dC�ɱ_hk%b��r(�2��{�8C�	,$�Έ�@�)r|\����1�jB䉵v��dѕDE	0u,9hua�y:B�M1d<i���9E�����Do@�B䉍7�Pi&�;B�ۤ��l!�B�I�TS VXMI�q.Hd�vB�	C88�@#��v�	�#��1t(8B�	�-�� �Ӧ��\��S1c�:"B䉽:pR���U]�(��A�1��B��4���'�]�~`�pBiϋ-^C�4�D���6!��$���7y!�ȳ'�a���}I:�`�@4i\��^��x�ؕ�ܗS�%�q�R0�y�\� �H8SiD����`!��yB�܇dq@��U̙��E��Ȁ�y�D?I0 1n�&H���Y����y�Ѥ ��5� 圳/�ډP�����ybcS�줬�ӫ�7TA�²K��y��i.�'�<)Fx�F��y�l��H~b�Q��|�Dl��@B��y�7D��	A�S5|\�qA��0�y�g�3=�4c�O#z���1�H˶�y�m.O �jamW�"�J|l�y�
M� �|��¯�'��l@�P;�y�kE&(R��V
jqzҡ��y�ʖ��e��A=[S4���L��y���/L�d8��3VD������y2��5s9�P�E(FTp���9�y
� �9�C�*��Zg�,w��y#�"Ox*��0`*��ꢀڧZ��( �"O�8�'L�Qp�0x �ʊ_�b�Y1"OvEa�n��i������N�9g��1R"O��q�ħc����o��za�%"O։��}
h4SnR=`gR�a"O��*��rK��� ��J�kK��"O��a*R���Ap� �L`�z�"O��(���]�t���O, O<)��"O5�S��)�P�2&IȞ��q�"Ol@kU��(Am�F�ʍcr	�%"O�x@g�� �A6�Wh�*� T"O �Y�
F2��4'˔@*y���'D�GIʭ_r�� �q~�qb�!3D��j�Ŏ�`�dX�+F
b&xI�1M%D�l9��1\���c����l8v9�-7D��`�mR�\?<�,��^��5�4D��)�� �<E�xᤌ���N�C&1D�\2ri�3?b���ηzb�d�e0D�L��C�:���u�J)Mr
m�r�:�OM����?5ԭ�c��O�� #�8Dw�@�D�hh<1%�C��,���*�2ՔA��Lm�'�\i���/<`��~�boU����#2ᕒ:��t��	�c�<��MW1Z���b�ؔV��j�J�۟4�EhQ�)��m��>E�TLM�c����qo�3H���J��O�!�&pU& ��B[��\�QI6���	ieJ,3�F&@ay"ɪo]9"+�crT{��tڀ��V�<§,l���$���'��4�iHB��ɺ=
�'���he�@��Lt��ўm�L̓RnHQ�%�1�u��O���&ΐ}�Y�U�'��Jߓ\ͮYb�L�>I�D��/g�a(���*f*eR$%�<��f�������8�7�۬����cdK:���!��dQ�<L�E��HϴBx�J��H�^(������$�Ǌd������k���T�'K�ɡ'-�H���Qj�	&P�50�~�1O�Z�OR��p�Y\%�b�IB�a�>Ȣq��2f��T���K,�졄�����u��KW�r��B�A4�(!�\Y��pMA
';*5@��2uJZ����9/���>�� a�3s�Yp1-QR`��K�!\OLl��<�剫U��pooK�,[��� 8o&�YCg171F��hѢu�n��n"�Ӓ/�4�&U�5CS$J���i!B�{�dL�=��!ԿA:6�E��N̈́JjFi�kN�U;,a[[a C��|�Fh�gV�5��`X%�6PD�Ї�	�>L�hH(� ~�<�s1�� g�q�[?1O��{�O�R �7� /7���!� �z1"��JRв��ƚz���e�m��i�U4Bt���Q8|�8Z��-AY[�#U�3���ɝ�U J�B���5��U�2�H
�\��RT�c�;/h�5��{ ��ʰ�Cr���������P��V����ְ;U���΢ʈt�g��?���U)t�^�[PH�?�����кCb/}B��4�z����t8y e��9��'��q�7�	O �3��;l�򴙇��z|�0��`@]�E��-_�9�j�����X����IAJ]ax"�#�T�5![�P z���N�qb�|��Xr^�3�BU ������' Α�'�+c��|��gl�4^��$ �ak�}��o��t��$1\OU1C��2"�P�Vnʇtp8�`�@@5s��a6�/e�}J�cQX$��)^��S���:u�=��T1JY(�#���2�Ґ�9p��IV��!w��c�P5Q&}e����>271O��� ��xr DQ�q�S����7-�!u�e�W鋰/	0Qa���J����56)��3%Ձ,*�awK�CG6���FV�d= ���;67��r�l��dTH����䖁c�hc�x�ׅ��f����)�h'�ɢ## ���9�̩�!�]��l�'dй�f��kZ��J�*�9m]���A�;P��I�Q��I��I�0$�2�d�obT59�h�:!+FDG
	SϦ��"NE�C���j4�|Z�%xmRpbgoG�C�,5� ߁T>�H�'�����9b$�3S�˙w�8|�c��01Y"N��?y��5|��(�	���T����q�?�*����]��@�� �yl9�O*��%k�."]�\8!��A���h���-`6� �MߧW��p�ϭvY���޴̪ɻtJ"�?����c�YDu*9��(ԕ[ن�	?{Nj����-!��pD��?Zz�B�)=:x���N�Vt�)���
�? �������UxH(0J��״
�̌����3<��ɏ)���[�E''�ʰh%�P�̧U�P0�}>� L�C�V�R��A�E�`���jP"O~���̎$�zRo��-pk�m���JǛ�guf�؆���n��b�?�	����0��+c�Λ�f���H2L�!��3p�l�k�G2Ҝ�ƯI�$�zU�.�]06!;�+ݙ*|��K6�O&��1	��Obd�'�?Ţai ��?��P��'��(*[#I\ �k�`��� ���WMb����e~ ���o�%�~2M�*�Ї�IѼ��$"z�(��\���'���U�F9Jd�&*����V8���*j>)2�o�z�G��)x�8g�ͻ�y�ř�6�ƀ�va�+%Z��Qj� Jڜ�h'b�,����p�b�VY����w�!�M��Nm����I�,e�
�:�'�=�"�D�]n����Y(�l���3h�N�Y��n��{򄂄7T��bg��TB�C�Ź�0=�7M�-j!�RTg���o�~A���$�:���R/k_�C�*?�X��#�8=�@�`�4\fb�@�h��f��G��>ki���m��r���2�$0�0B�Ɇ;�d�s)�2H�*}���)J:�l�'DV�ēt�G��O�Ђ��Y`HBv�I���4"OhШ�M�Q��a�$]�E��H���:��5��'/�M��Hڶ	�L��y���דC���pI<���Jج��f��o�%dH!��$oT� "�F���43ƀ==4!�]�V������ j��pO�f!��ՈUFR�Z�I#�̉b��Q&~�!�˰kV�ȡj'I�&�x�#س5�!򄋥R���pc��!� %z��Q�a�!�d��VdA�ƤD�[���c�A !�!�5V��4{�ՎF�
�P�S+&p!�$O���Ի$�;�������!�@$8pp�;pl�cb�џf�!�F���=��G�ye�9��QX�!�dţL2����>X�t��ֳv�!��4�t��B4`���צ�7q!�D�?Q��R�Ѐo�L@�FSw�!򄃓:�d1FE��������9|�!�X���0�G�+����ˀ�@�!����Xh�G�BȞ�2��O!�D�7L\�x��*_+���h�+Y?D!�d���0	���Q���x�+]�~�!��#"�*�ছw���ۂ�[��!�8�I��̺,Ąx��� �{2!�$�PR<��e�G�z$q0*+*!򄃔�������z�ڥHN8�!�d�0h_�,e��̨!gm�%Jm!�D�	$��y2a"t���͈�PQ��{�E����*�5��s�8�+"�T3F����e"O�)���%�
Aٓ���E�*���8}�W���O,A���B���ˮ%�fuH��ݮ
A
xz��ފ)H��}Bu���ظ�8�I8q�4�[��'@X<ibGװ/R�s�o��Z�dĊ��đ"~d-H>ɉ���S�H:r�̓!`TZ��X*>�@��=Yi���Dmt$�����'���g~��I /�0���.O}}rc�22b��'�8�&�Щ�.i����[y�L��4OsNa�g��<ɰV�u3ʝ�F�0r���B%c�<tI�|�`"��!{x�+�I�}mp�r������N�pe�[� �.IH�#�[���"O��RE����U����C΀����/aX����|r�����xn0��5b��4���03	"D�H)�m�;{q�!���d�J�3 ~���' $b��dģ`�8���bX�b�
@�a�!�䀣0�� ��S>S&� ��V=3�!�\0@$t�Cu��{q$���]-!�ވB��Q��ʴb^z)Vo·�!�]2[�QɡH���l쨃��,`�!�U�
ib�����@���R��"!�� b]8��ͦ>�0��ML�HŃr"O�QbtKԫC����nS�n�@kS"O��Zϋ`�I�U��
0}Ba�"O�8֦�)<�ȱթ�2��<��"O��jb�*p��``�i4rh�+ "O�EB�,3�(8�&�P0V]0�)R"O Q�aDC�,�#��;V�VY��"O�d�`O�^Eܜ�����p��r"O,�@e+N-t�:-��Q,S���f"OYH��7TM(���m��U����"O��j%"$+ɞ �w�I#8��U�C*O|!ʠe]�4d�Q.��>�|��
�'뼶NF3H��l�%F�aq��a
�'�f8he,��OdV�%���&�	�
�'?rL�r�4o�<H�)���8 C�'k�U�tAI�`�ʭ��#_���'�>4�rb��;��|�ר�0a�'4�	�cO�X2t��'E?�, (�'��pw��q�J���BH`�'Ov��(K/i�i:e䘿�<T��'�\�H�T`L	  �
#��@�'�R�Pd���hS��v��{{~���'�$3�ǂ1	H�0��m��Q�'R	�cϗ���S��a��H�
�'���!�E�H Q��KJ ��'p����Fb�9`B��x�D���'�N��n� /� t)`��#��Q�'�����'u�UyT��0@i
�' ��ufQ���Q0�b�6'���'E�e`��A�ud\�T+��T����'"��cRMS�8��_p�u���y҆R�[�^`s�.�r`�%JKL��y��+@�nU���i.nq��/@��y�$R&}�^���\�Z�ؔ�.�y׉Q�^�p��4R��D�y���H��H� 蓫g�Y����y2�W�\B���.�p���.Q&�y"��8׶l����s#ԥ�y�G,T����\�@�@R� 2�yÛ@^j�+�9���AA)�y�E
.����V �� y^=h�� �y���`�(�Yf���,�nT�ʃ%�yrk
r�
���[\��x�4��g�<��o���7�V'z�� ��r�<�@��=7�䔠�i&A��� ��\r�<Q�(N!o��"@��#Yxy���G�<PCO�O�\�9F$��paȀN�<YpK(��Xc�D34�S��	R�<A��V'.�2`��K�?`�N��flI�<)��-e��T���A�B�8��bF�<�@��S��	�G,q���a�F�<��)J��xBiے\*� �D�<9V$^�k$ҽ����M���v`ZD�<�@H�o���ʏM�F0y�o�}�<�0�зP����jÉ,
�	���^�<r�D�(}��F&{l�h�+^�<1w��L9>�Z�&O�R_�� �C_W�<�T	�|��I�P�������G�S�<alT�g����v��12���4��N�<��˄(Tz��zF��.�ݠ�a�c�<�BNI#a�V�q �� &v���X�<��/۲E��F�/#��3�d�}�<�D��z�@Y
�n�>����VF}�<�u㜱6��(��\�(](�� �A�<� ���!͈;ntK��]60.��07"O�Z�Ȗ�E�vyz�蟹s��q"O�1�v�&�$9���q,���"OJ�%@��.���`צ^�%����Q"O���Ε�9Q� 	v��r��;4�Ip����Mm�H5h
5kLЙ�*�!�Ĝ<?BV�"�O.p�Y���¢C	!�j��(��=Y�E{�鉹0�!�d�G�a����{nV$���˪vA!�D�~��J�㗯S^2h�(K�g,!�$Ϙ��5��S�&{�8�(�z !�܆X�Z�釂��7d0]��	�Q&!���-
�)9�	�*E��3&�%!�$�7Th6a@��$:�*feE24`!�F�)C yS'��l���C�->F!��RI.أs�ZRG�M�B�8T!��0r�r 9G�?b)&�IeO"�!�$_�-ްy�&ԒP��I)��ߣ �!�DVv��(u���Z`�R`��q�!�$�mkh��@�^2OxJ�z֌mq!���!Vv|-9 �A�%p��"!.$�!��J�� � ��I�@�tLh7�X<	�!�D�A8��X� N�s��	vh�?�!��߻W:,�Ճ�|`�@��
#j!�$̡E��u�!O>��d��8`!�$�p��1s� H�`㨎^_!�dʺ@��Չ�C֗I�h�p��JI!���7X:$����׌�T烄N%!�ʁ1$��ŕ2|�d�y�l�4&!�V0���H¬6�tqp��5w!��ϒ6ª���4C� y� �]�lm!�䏥iPR��k��ZD;��>e!��\�{���+��q�V0�dςgY�䓠>ma~r�qt���sM�.Nx��q�Y��0> �"}blD�9�F���X�B���:�N��y2%�p�X[�l!6C(�H�`:�O�C��O��볫�LOj���Ž>���'/��	>E;0�I(c�V=��%PT���>�b�|�mȢɦQ��*P�ȓ#����UeYva6����8�X��	$��?��"�#M𢽒�B��%�Q�ii��t�c E�N?���'Z���E��DD8�(�o�� >z���'�����SES��B�u�iÌ{�'��zc����X���G|�q{4a�b�i�"O�y�"ʋWd`� ��,Rڌ�C�n�'�"}�'ʰ�y��G/c���IWÇ��a	�'�6�с���K�d0��KЬq�
�'N:9�TE�9Ħպ!n��,��'IdѪ9�p<���+V�a�'�Hl���N�O���� U:A׸8��'�"�[v�S+M&M{2$B4?.� �'���X��Ѹ;Ni�QA�C��)��'@�᫑CE3�n���ڌ@���	�'>H�;��ɪu�\˃i=��h�	�'���b��.������/0h�1@	�'�p������^�
�5(ښY��'�Hy0�A�v�0Y�UA/z��ؙ
�'�A
�+̵�F�r%��!1X�k
�'��:��Xq�����)e3
�'�ڨ��LΒ+����X�Y1fP��'*���E�M�mt♂��#z�t��'�� ��%N.2>�����u?,�h�'<���7����rH%|2���'��	��L".Yf5��B�l��M���� F��5����V��O'� �"OV*E�;*�n���*g�����'#�$E�����Н[Ө�$��g!�D9|�e�Fm��+�d�hPMӨ1n!�M�mZ�*���;�B���Лe�!��y�h�եֻW�4��/�@!�䝧OGЁ 1��5e�@��@F�!��Eb<�l	�,,�0ϙ��!򤐳6��U@�5�"��=}�!�Ă7�FE�v ��?����k�:}!���hz�q���:}[�	��m!��,m�X��܊'e�iO�=e!��7��Z��n&p�+���5e!�F?;�dUX�� D'nE�-�!��D�F �Y1o�	D�(��*D��!�Cv̘�b��nd>��6
��!��~F]��I�`d*qr��1b!��*.����&[�uD��XE�ɗZ*!�d�9`ޤ�AO�;I?�0@F�1y!��ǈ4��XP@�>��Ԉ���=�!�D�O��Q��G�}��Q�!�V�qJ�����b*T!!Ȯ �!�D�.Y��e���[.��ұ�\�L�!�To�5;G$Q�H�0��*�{�!�Ǎ1g긁�[f����2$!�7dH �B��8.��֍�
�Py�B�p��@�m�t�P '�։�yr"K>� tRe
�)t �0�*��y��"Tք�2`�t�9�5���yҩ�#k��	��Ǳh����u�[��yb�V:���8%hB�5hH��샜�y",U�@d����u�Y+�L�y����H��G�~����yRЭil�@��	z{BU�`�ߧ�y�@ߢZ\��H���>2�py�����yr�S�&�l9w�7G�@S���yr�D�w�%	��=�VV�.1|���.�jĤ	�r=*�Q5�U2L��ȓJ�:��J�_|��sp��/H�&ՄȓL+��w���.�@���.e�,��T谨�,T�A�8B�h�3!���ȓ
��#�3<�l�br��:<�ȓ'��}2��݈zL&��O�in�D�ȓpi��kEP�x���&�Զ0�0\�ȓ!k���e"_�q�8Ë�0z�P��ȓV?�B�.J5_� �"t�4}C�U��Q �̩te��A��=b�a�
- H�ȓ|��aPK�Vg��	7�mת���;���� \�\U�I�΅�-[p��I<����h"�e����>�\�ȓ8~Q�ì0�����
�3=�2���9������68,a�,w0�����S ���9��I 7gӦNĄ��	a�'��E��C��&I�W��n�^���'����1@�����6(O�X�v�
�'9�t����&a�*Mt�H��BК����)S��u���ʝU}��ȓ+���萞M�|��%�Ix��P��Ѩl��ɛNy�`�C��T��]��F��{�bȪn�b���ϨyVń���-Y�)��iR.\�H�4�ȓD`-��].^���h4�5�☇�_���1��VU�F��?[�|��-�p�f^ e>�h�V,u�x��S�? ��B���?@m7���.OH�4"O���vHW�3�z�E/�046R��`"Ou2S� Z���Boөk,����"O�Q�F�'S��)Qm�m&Xq�"On�J �%W�1C��9Xt��"O����Ƙ�<��5z�a��N@���"O�x�(|�n�J�%HIM�"O� �a��8s�r #CCBE�'��lZB,V�!�Z@�#�Z� �zŃ�'l �� ���R!�E,^�J���
�'���	��ϒ0�&[�dǷ
'R)q
�'�fd�đ�UƼD�2�A� h�$�	�'���1`�2eٚ��V={K	�'ӎ4�E�@ȝ�@���v� �'٘���C��[�^�{@/%�r�[�'z���U`ڥ�
�'�Z�wp��'!�L�c@�.�p����j$�X
�'1���P.˓x���U��P���X	�'��k�F��c�V8��Em̤��'+\�а�M�7
h�:b���9Id,�
�'zh�R��4a��ĭ�2���
�'���Ye�Z(fnd=�D+��y����'@�˗d5o8�L��6�:�'��ir��/
ظ��L	e�B�"�'˰�"���R)�Hՠ*����'�
�<F 4�� cY�MJ:x	�'qt��g�Uq ���.|���	�'��AQ0���'��'�I�#�!�	�'�N��,G!�@��k,-o����'�D�0&^>f�Ա���Dl�A�'�*	�$ :LO
4S@�+�����'���a!��n�1���������'�ʰ��E��u�O�� �'�j����B� ٠�&-5
��D��'�����$�lq��":
!�'���ԏ��K9�����<-h�<P�'6l�R��>��6V17�\)a�'3����m�
w0Xi���/%�z���'i�͑t�
 �f4�C�#m���'2r�2�F�j�i���<n�Zi�'&�iX7H��T�#dE�<"�8�'΂��5I5nr�`c'�3:P���'zF)���޻{���S��4k���'R~�Vi��w�T$��`�:��J�'3<������;�`���B�d��'�,��@$J3ex���=B5�'����U/H9���B�a����'�l(��۔BoJ�x��#c���'vN���g_m0������.0=��3�'��<������P#�ַ!k�"�'��i��nO:`���`eN,�9�'J�)��ĺBE��ևծM݂�r�'v��"b�	>ML��u��L�f�p�'�v��&/O�&P���� PK2~��
�'�6�2�Ad �SCS<���'�r�腮�.8Z)��@��g�V�x�'�l���_�|f032��!dM��I�'qd�Y+[�S�l��B��
V�"��'jX=[�:w��|	��Y<UFV��	�'���v�A�N�3J�M�n3	�'���'Te
.` �o��{�nU�'ʲ5s���h1^�����\�3
�'�l�B#Ӵ<�<]X�kX�~#f��	�'�vLPSl�	Mު	�ʔ�qI�}���� ��ʢ ׂ�^a�7$ܶw�D���"O^ԁe`�*��,�1���w��P&"O�)aEĤ*�D9L\�`Ǣ�x�"O���$CP�gnbTy 놎g⚌�V"O~�AAa���Y*����sl`��"O�T0��2d�m�b(~d�$��"OHE�#�ޘj���S�o��IR�"O��v�ŌO�Z(�Mǭ?RL "OD嘦�H_.��b׫�82J2��s"O�ۣυ_JZ ��N���]�q"O
x0$	�)!ʮ�۔������q�"O��r�]��!���\�(�ִ�r"O�dQ��3b. �4%�z)�B"O|�ˤ&T�Ȩ�v�&�j!"O~���>kwB5��E�=%�ur�"O��C��*d6� �
(�m �"O��3���m���n6�#"O�Q�Ƞm���#�H7w����"O*�ҧGK�F�P�hF^�#H����"O:�S�,��? L��$ʉ4"FJ��t"OJU"LӼ�r����-k6�B2"O,�����T�^11��[4>!V�"Onh`Av]x<�AF͘c�� �"O���''��)J��$EǳlYD[ "O����+��w�($x���(�@<�u*O�5S�M"��!�ܝ5�,��'�2��v� �<g^��b�9k��Y�'`��y�S	����,�@(�'��`�W"�	4RH�1�+X�:��2�'t!����x�QV�Z�@a*�	�'��`�p���wB(�إ���@$��i�'^ӅBo�����Ƙ9��4��'��,Am�<�8�Q��[�@.�
�'�:�S�g�`�j�kq�� 2���'���b�I�/`�`���E�;dp�@�'Mxۢ�ım��Sa�G~�x�(	�'3dy���¬>���n��jvv���'�D��L�U���A'��d�tȳ	�'�1`�fW�N�Б�w-B�q����'�V�]�R����&H�A���@	�']�d��&]�Hx���׃
�GfdX�'�����d���(��GyVԘ�'d�\���/B�4Ӵ>�ji8�'��H��oT$�����?_��ч�\8�,
�c�;����5�����ȓ ��{Ԏ	�&�`����*��@�ȓ_l���gت3���� hަ(xD��h.M�A#'�X'�(v ������]�a#E
Ht�y3�&7h$��5�R1so�9�0�#$�_$I�	��0D�Ր�ѝ#c�Ļ�I�@` ��ȓ]~�I�ꛐ�L" Ћe8��s��CT��5u<��W뇄9G��ȓ�L�C�3b���*�a�>Z�4�ȓId���"˩gI�Z���:6�U�ȓ
	@}Q�%� ���r��:4T�l��<���g*D�ĥ)`���0fv�ȓ53�������d~�� ^[�<�AH����Y�hߩhQ�DӁ B�<	h�&\��U��]�s�����{�<1�Կ|
��"�*k�X�h��r�<$bW9cɜL �ѝEzL�C#Jo�<��MH5�4[��B0=4�В��j�<�$ŀ���$ �W#��x���h�<� ��0��ۑl1���i�up@�r"O��;w����}2�>�8��S"O�t��i���0�B� ܱ"OR�cw�JA�4���8�P�I�"O���aM�$�Q�aB�/����""O� @틦���#n-_�H黡"Od��(��P����-ɤ;I��$"OD����
`Ҿ��JD���|	�"O@� ��S�~4y��M���ɔ"Oڕ��/V���a%��"OP�AO�PPdY#��)g`�(�"O�yZ�I� ��`[��6hT��C"O<9�Q`�#�nu���='�i�"O���f��NЬ 3��Y�z�z�"@"OF�"���DśЉ�;��a�d"O`�X��]�$d:�I��#�d�x�"O"��Oؕ0T�10�͈�S��m��"O�|:r'��]� 1�'��~q���u"O�ݰ�� Z�6��6N	�`Y�Xr"OJPT	�6@���[�VK^s�"O��EBT��UZ#B�|&�$�"O�T��� 9�N���D�4)'"O�$�! �?8�\�y��@;Y'f!�C��F�O$|H)��>N��lx �����	�'���X7��A������Ǝ��	�'�"P� &W�8X�hI3 g�J	�'Z�ui��: �L���"~YD�ʓq�H��-S69�q!C�&}`ȼ��v�y� dW�Iњ@����(7\e�ȓz�hQ�g�`�J)�
0un�ȓc���A0���p�պEϮ=��͆�	2��wF��!��4��.>���ȓA�.��v�YT��A��z�ŌG�<�#�A&:�xIǞ�b��e�D�<�%��P�~�%���0�J��Ɵ��'aɧ��dJ��u
��@Ws����  �!�dȯi�x !-)`*E�c`D?V�!�d-������L�d�¬q6j��Q!�D�K/���,ͧD��`'�
l!!��*%BEY�C3Z�&m�� :!�G�.�&�w�э#&��:��Ͷ2!�d�E��%��P*M��b[�~ў�D�I��4��pr���<�#��k�'�a|B�ςs\dU��D�;w�h��(��y�ɟ?j�t 'f�k�t|rp�@�yB��|��|� �ʓRg�d0����y��R&�0@��Έ�?�1h�,�yD�G��<Z3@���:��ÄQ���=1�yR^]^ �
�nE�Z�`M ƦѼ��'�ў�Oi�ԑ�)�,�`qzE�[�T��a�r�)��È�[!ZM�s�Kd�,������0>)SÒ�^<1��D�vP�͌J�<�h�Ysj�z�5'<b��0*n�<��͋�����'|�����<���m��C�IT�)Np%8�ɋwh<Y�ڸ`���b4L@68)�F���y"�X�Pe�a�2��.3 ųꙄ�y*
	$�.�	!��Q֜A��Ƚ��'�az�JT={�
�ׇ�7���+�Δ�ybа�8����.��4x��˴�PyR���t��ĔJA"��%AR�<�ӊ\�>�(�G
�> =a��M�<�u�V��Px�p�I����`TGy�i>��<�掝�h�@���M5�LRp'�{�<� ^��r�Ap���R�7f�Q�]�8E{��)���}���Ϟa��L�c���!�# P�(�&�@�z����O!�ęw��;%d�5$k`�{��Ǻ?C!�d(��{A������N
H!��$ �x�sC�:�´�Vh�9!�UVo�����N����1�!�d�*J�:�c��זwu*L�c��2�!��N#� ��%��O����ue�N�!�DҐA��;%	��[R(3�Ꞿk�!�$�H�<�����;1�]`�&)�!��X�^Te��%�O<�M���ѕ!!��J�tt�Gτ~��|�qG	@!�$�g;�I[э�}P�}�U�1�!�8`蜥k�j̦]0(@!��f�!�D۠?3`�d��J,)�g��'Pt!�d�O�n��]��r�#�.�=`!��K�"��+ŬU�vCGd#T�
�';"�$�%�|�DYf�H�'���#%>�� �&M���x�'��걪������+ֿ9�����'
��!K>O�@��C�.#� ����xB��Qج�#Ѩ��Hql�0���y��
�ܼ(�N'QAV�Iu��yR�ߛKM���#���>���+�쇆�y2J�%~Un�@��A�^s�l�r�:��>��O(�s0�S6dD�a ��RE���""O$y��9;,qI��9=p��c�'�!��7lV�]zB����|��1��_u�Ii��(�0�c�))�`3u�M h�E��"O4��mA��lT��߯%:�a�"O�1���즙�en� c@���@"O�((��P9 ��@����q%"O|�Dɕ�F>�k���%{(�B7"O�%���-q�
���j�	h�}Q�"O��s�)^-cEv���α]�t��"Od ����(8t�Z�ϒA_R|�t"OP0#'-e%ZчLܢ[W��e"Oz��t��#3q��)S-E2�"OFa�7-�<U��4)��?8t,�V�	h>�1h��0;��1sD���� �d6�S�''��v�Iq�Ա��}�朇ȓw�X��R�ǐ5J<\���{��!��)@�)���oݰ򡅿A�.(�ȓp@@����T ���#e��A�ȓ}�2����h�*iK��Y�~_�ȇȓ1��d����7k�[�}�,X��7v$`u"��6W� ��'��_�<r�'���Á�T3�����Mp����'���0w�Hp��K��If���'�0��_�AH����ǗJm�܋�'�L���fA1��x��P� �Y��'��1s��;!��j��>���i�'H�-��ā<EP�X�Ïb�J�'�4���'�-jݸ�9� (x��4"�'ϪI"b�����4a���w��٫�'l�~�)�' 	:�%Ǩ�[tE5n� ԛ�'r��XeM�̸,�6������'EָP��R?N$���ku�l�Z�"O�]@�l��sͼU���
���rD"Oؼ����[~"�Q )L�g�Ne��"O�4��M��A��I��>5�!�"O^ �Q�]:5w�tqṽ�;�v8�S"O���&b]Q�V�j�A�M� sS�|��)�3� ��	C�C�L��%pF%��I���!"OF��ЧEI��1�~�>���"O�%�*����]ѵ�Р��D��"Om�ԏ�b�8�c�#� up\8�"Ofq2r䎌vN(<��`�<�"��B�'��:��uBD�#�L T;n��$�7�O��h�tC�f:Z�0b/Ɯņ�_V�U!$�Q������E�mL�d��w���h�B�������
�EbQ��C͜1�H��j�9g(��J�P"O��Y#
A:J̄��@�fi�W"O�y@D@�U�p�rA�&N�X�T�'B�'6+��S�v�X�ZW��3s�Nȱ��'$���tŁ��R',��e$�9z�!�DVO+pɋ�,�G؊�ycNY�F!�$/uD���G�"t���LIk�!�)V� ��&��!�z��jG�X�!�dĽ%�h��&��)S�vY�"H5,�!�O,D�u�`��2l��Ő� Q/:�џ4E�T�;j1�)�G��t�~�ʧe����?q�'	2e�"�A@�aK�gA�z��Y
�'=l(���`���Q����ֵ�	�'�@I5b�&JP&��d�q���Q�'�*��4�ݹ�~���f^�y���'�8\�1l�?W�4��I[
\!���'xz�Q�@_� �RC�� W�؉��'~Ř��^�ǳ�$kA/�^�<Q��V��H��G�	��jS��^�<a�gͨL��!����fT�02��W�<����!`:�%��M�61GRm�C�CW�<I'��|�8A�e'�5q3F��h�Q�<�U$@�L �ݩ�)ʳ/�	ۃNX�<�b �+N��ш�i��2�W�<��):N(��� B.t�܉�&��Ux��GxD'�P��Gɘ<P���*œ��yB�4h�%���D�K��|�S!5�y�b�Bg�PJc��C?�`aC�Z�y���#$��U�޹h�̡	��×�y��H�jF
�j�́�l��  d���y�i[��ꜱ��._�t�"J ��xB�9HP���z�||9��I{��t���ᧂ���r'p�йZc,D���GN�$:9%O�(V	�Ã�+D���p��:`6,�Q�T�� `g)D�Њ�g
a��������k<D�H:���=t�P���^1&��9D����L�u�:t`$�Ȳ\P�Q��K8|OLb���/��/�"�R)P=��H&K4|Ob�ф���G��$��ďoU���O2��k����եB�fwB�R�ˍ6X�
�JfH1D�𪶌^?5u���!k�
��c�/D���rC}��P�f/<����S�.D��а��o=�FjKh΢qKn-D�8�N1.�!���Y�l�(,D��
���Z�4���"x[Bz��)D��i���&�4,��M܏�� ��"D���C�$@�-�W!ږ?��� �,D�)`���Ɖf��po�!�=D���b�Y�F���R�&"Zd�1��(D��z0a��r�[��S�C.�sŦ&D��A1�{��5��E�&E�����"D�XOQ��tCf���H6�	�'�"D������Q��ͦe9Do�A���0=�t��1)>�i��Ԫ�]k�@�z�<� 6y�p�	).~U{�@-)��Y�"Ot}!e�Vj80��N��D�q�|��)[*X�`�dc�$I!FO�yL0B�	�4����V}�<�Վ�	�jC䉻5�	PRM�5V��������C�$9Č���s���T�53)dC�}-��d���`���6C�-�*��͉42�4�4CE�m�`C�	k�����ho�r�ñEH>��D&|��87��[5�5�T��8����ȓ>������r"�8+��GM��=��V]����3�t��pB�,'����&�>MsӬW.A���֥1�����r4��@��R��A�Hx���q��8��>�2��#��l��+6A��x�^�a5�γC3�`Gb�sbd�KE �}�P���*�DC�<1�PY�U�;|JH]�f.��7C�I#<�`�rȚ?�KA�F�*���"O"�ٲ�ײh��xCq��A[�!�"O*����*ɨh���\:Wl��"O�� ���mI�[5׀WF��x�"O�8���WL���K(=rDJ"O ]��˓�#�d����
�g1��J��'�ў"~�e�$2E^}�Ҁ�<�@�1A�P(�y"�O�K��PZwÓ9�����j\/�yB΀� $]��%�=^-Ԕ��)�y���wB&P�B��(�8Y�uƒ%�y�8h�h���P�W�QbE��y�W%QB	��(]I��!#��"�y�2���)�b7@�PX��L��yrL��L���ⱋ>iv��h�E�&�y�U$ܜ�yv�-��&�<��?ɘ'n�i��ዪc>�K7� Or,��'Z��x#l��B�>��n�~2}��'j2 B�d�-uh|*�a�!���'����D�F�m�hG����B�' ����OǪ�v#�<�"�B�'�T�g�Y�/����O� b]�'���(0n�x�Q"E��ma~�k���2�^$��h�#4�8�L�J�j��r"O�#����䩐j��y���S$"O�,C	�J�����E�����'"O��rv�V��p@'�s�l*4V��E{��T�U$+L��I�5h��,Ɛ E{�O���͙.
t;6��{�2��
�'��y-�$0��x`蘰}��	�'��!F�b�&��P��>nvRih�b�'���	�ƙ�X���WJJ���'!D���g�L�ZLa�%�J��I�'j��s��&%��es6�� >�|���hO?��D�:S �0��_�Bٞf��ȓ,p� CB�ɠ��,^.��ȓ@R̭X@DխG�`+�&�ktbmD{�Ot��)v.N&��V�W�u����'ء8��g�8�f�b�#cΐW�<QM��ai�,RW,L%���{�<��`L�i�R`;"gʎV���0t�<�S���B�c	1h�\9�#Fpx�4�'v �7I�0o�,�P�v,I!��k�<12���w�(�ӏU�F�D�
��o���ϓ�dH��~����Lզw�h��ȓCO����Ó:D=y�ʣ|'f,�ȓNr,�q��_��X ���
J�!��S�? �EVOX�0���b ��uv��R"O�X���0��D P��"]�5"O%��͛$#z}�S��9~��%"O�D�Ee�'`Pњ3(	�5u,<'"O��IGm��$�"�� �y	��2�"O��<mTY	1�x��
�"Ob9�D�*^^���c�0�eʂ"O�}���uu̐���C��S�"O�q���ۦF׸e�D��T6\�e�|��)�ME}� חd\��X@�I5�|C�ɔ$��)���:b�!+���p7�C䉟~T��W�.^����n2?��C�� dd��F�K.^d�P֮V��P��F�"�"W�
���(�s�ñs����	/��Y ,�n�x����T�ȓo�H�����N>�͙r�\�(L�i'�|����A�k@"ؚ�9��:��C�!E@|[c��b^h�{�ˋ�Q�x��d'�*�ԋ�*�X]g/�w����0�8H�sd�^�Pb� `�艆ȓ���sj��a����fOH!�ȓq��5���ƧyV�����2a�.���+f��h���R���/!��ȓg�2=�w \*����*8��t�ȓ#��H4 ؗ@֨qQcX�"��-�ȓ#�Ԑ�&iV�{�^�i�M�1q�؆����"JCv�Ε��c�V;^\�ȓ�	y�k��[ޤٹ���,�ȓl4R��GI��8{�E�-ED:��ȓ]m\�Y�J�B����F��ȓf���ԧ�H%�=)Q��M�2��ȓ=�40H�)�/�D!١挌Z�d1�ȓubX�-�!��Ȑ�TT�$م�#�mi�o.lhx�����m}�H�ȓM�^aG���3���xf`���&��ȓ\��bI9�t�b�č86䁇ȓkMܱ1bF٬.w� CJ:JM�e���v�yI�<Od��1�]�	�8��f�P�Hg%� 11��&˖�C�,��ȓR2j̑�l+b<đsHZ|�̆�<�z��#�()���`����1�ȓ<2�H��'�q��e��8p���!`"���(C ��� 8_H�r�)�$ã\ �LZ���L�ـk��yB�ޑm�� �cn��+��	�Њ ��yRfɣ:�*$��B�'V����-�y�C\?g(Pu2b��wȲ\��ϖ��?�'xJ�a��Ht`�!Kȍݴ�@�'����E�8P�E2��ˏ� Y��'}���A�E��`Q�(�:����'��M��I�2n?����[U^U�
�'i�:%��*�de�6(�3�E��'a��Ϗ�?t���vj� �2-��'��M���?^>\;Ueݵ��b�'M8�^!^�FU�'�z�f��'�|�`wEG-8�^�W��w02�B�'h�{��;	窭�d�l�ⴃ�'�.U��̌O�(��˘�4.�	
ϓ�O����N�bÔ��E%�>P����"O�H�5O�x��*4���VGHԃb�	R>yp���-0��f�1�<K��#D�Љ�c̚PM���c�@�p0|<��"D��Q���H�6��k�z6B���-D���D偡icb�� /)I�}���+��w���3� \��Sd�,�0��OW�|~"@��"O�����7��EH㨏�Pq�#�"O�	� J�����%�].Sa���'���C	(c��������B�;D��)��!*�d�q���t?��w*OX$���"Np�6�Y�\�q�`"O�0�� +���!�O�Ty��c�"O���V �o3u�7��Dy�Dr�*O(]A��9dj҂�	6���
�'��0"%�[=Νx�1;Y0�2�'���Y����k-8M��Mŷ<a���'�8�x�m�<��D�l�5�@\�ʓWT��@�x���Gƒ���]�ȓh�����&=�ru/�<t��ȓs���s��fh���>�i��QA�AY7.����E�â]�m=.Ԅ�/�kD(E�?��a��e�/��-��s�e`�ƞ��j���j�-i��ȓB��S"!	�,�����G�>?o~���09°�1t�6,���ضu�V��ȓ�v�*"�L�E�ZEɷ�]����ȓE��� �%��O&4��E$@0�����M�Ly�m	�	�
)�`��s̀��"4��2 [��t��1͍�b��ȓKĵb���qA��ѤkUF���W+��x�*
$ު��ݞVw�A��@�LQ�$�
8Cԍ�Y}���"O���J�V��	��
(2^�q@"O�󡭝+}>h�VN�>�H���"Op�!��N �@���,Y",��11�"O,e{�&�X#���JڵS�T�a1�'��Ih�r���#W�����8��C�	�"�����"tk>����K/��C�
7,�Y�R�-�
�Xf^�E�rC�I5l�(��J;�5��'^C�	5s���`�
[~eȂC˖PBC��.]��i���%}�H�	u�DMZ\B�8-*&�P�*�^�0��^^��=�'sZN�@
J9xeBL`��C6N����Qw(4���یGB���2NO��찆ȓs��0s-Y�8�� ��dG4N�ч�J�4��D\ ~8�g����-�ȓ$�밀�^p2��Ѓ���ȓNZڼ�@iܢ~�����]^�5��!뾍j']�-��{cS�*5��G�0�EB�(���ҶM�/7ՀT��Mk����/��;Kɹ$�� {��І�}=�����0Z�K�>����/C�$9s�^���Qᡄ�<UOf`��ph`�`�Ğa�yQ#�Y�� �'kB�X�d�$&���[�`H�j^���'�){�	�RBBa�nޅg���x�'+��B)ˤO�LТ���a+z	�'S:|  %á=�Z�A�W�V`�P�'�Fy�ӝ>��M� ���"O��B��b�:h"N�-�B�z "O`4q��q*�u  gƯ)�Y��"O�ca�L�g��0�֣J�.k�"O^���E8~��Cf �N�4�G"OR�ٱ/B�H<5zQg�8UJ�)�"Of�!�9<�|�:#�٘D�)؂"O��z����ٲ�A>�X��"O�mcl�{x�R��ع`�p*3"O�T�gղF�pm;�O�<�p��',!�� ���s�הq�Za)7�vT� C2"O �H�(/��%�F �|,3�"O��" 
d�K��O�b�����"O@`�q�%CsZ!6c��it�x!�"O
�����-<�QD�?XevtR�"O�M� c�!H6N��V
�7S:��T��D{��iý@���$$�0BH�ԃK�<W!���-���A�'6>?.����B�!�V4������$19L�|�!�D�	�8�v���+۲H ֪�+c�!��ܲ�jfF� s�@�����}!�΅* ��+Ti�â��@.x!��V�[��Q�pWk�%[!�Dׄ	�N}-���SN=&ۼa
�'�y��O�/
S�֬��	�'���G����@ҋ�Bl�
	�'O�\
4n�=0�iP�@�Uc�'���BÌ$�|T��(��0|`P��'ƺ8���;BP8�bT�#f:qP�'29�F�$[��:ٙf�B��
�'�ʤ�&#Շo@�� ZJ���
�'�L ���
��m��-NZ���9
�'����D.Ո(����� )��ib	�'na*4�3���s��kD��r�'Nذ�I�f�܁��KYOi��']\%2ҵj�*�{�)� �=��'5li��
�Z6����ޏA���q�'����Q$�,D2��'n�.��ݓ���/�z�!��@)P����1`�0�1�"O�A�%��<߼ ��@�W��$��"OX�9�݉Ϙ
я�7 �n��4"O��������z��`�"O8����6_<\�b�@پ���"O�,1`���*t�xt�C�`�!�"O0Y���=$��A�V#W�*��Ֆ|�P����K�
|2'MW�E�0sfJר84bʓ�0?) �5u��brj�3��8j�B	I�<�t���5��0�b�/9E䔰%�	L�<�*L�w�А��i��IX�V"\E�<�$N]�l��q��+O�
����^@�<���Q�d�:l˜}l숓&@�s��UyB�ONx`E؉W�Ȥ@��2hI�qsN>q
�'o(�0!�`*}��\�V/�I�'�a~bM�'�����A
-A楒En��hO"����\0���wo�� M�����$�!�䁔k��8[P��6)E(@���U6�!��0v�"���|>Z�� �{}Ȇ������/�fgإ�#�A+?
`I�ȓ<o@��b�u��@a��]#<:�t%���I�xV���iI�ZD� ��S>~B�ɯF�t0@D��7v�����N�g�>B䉼E�-A׍b�q���
��<B��e\`�s�˶a��Ҁb�7d�B�I�<7��Y�aX���Q�Z�C�	�X8��ӡC�\���6B��"��C�I_���%�B�de�[s�ԗZ�C�	OCL�B%W�(��R2M�,C��;@�X� ��i���[�-R�p��C�	�& `��指]Fe;Ŭ�[]hC�	W[�԰բ��+��k�B�)"�B䉀D�x`fϗ!�� ��=��C�q��I��Q-Pΰ����v\�B�	-[yx-�3��/>�e���ڤPoJB�	�a�,�M[♃U�Y�#$�Ox��� ��遊�
?���[�H"Τ�1��'�ў"~BC6,����O)��M���ͦ�y2-Q�b޸����M)X�@�Z�M��y���1qs`<��M��S@B�b!�\�y�%��lɀ �Ս�"I���ѧ�ݥ�y2Cw>X��썊Bڼ����
�yR�]�W�*���䎭?��Hg�=�?��R�ӫvhT��v̺@���y���3Y��i��	u�'r&0X@HJ�g�t8q���g�*5��'}*U���)S�%K�D߷^����
�'"�-�2�\O��p��N�O�=1
�'��Qm���	Q�B�K��8�*O:�=E�@ǫn�\�� Ƈ_���+����'�az"N@1�,�p3C���p����yR�D�M�:�I�3p�v@��y"D�;L��J��Q�}�h���ۙ�y򂌅nRą�t4	4m��y�E��5��y�+�:[*
��3����y���a� ���F�L���G�y�*�9\����!���ad���y��&�T@�(��/��ۢ-����?Q�'E�����^��!A��S6�����'���@�N�_7����a%� ���'�@�j�1U=�����>g��
�'�4A�Dg�G�1G�H�
d�b
�'P��SfI	!�&u�Q"��O_�T�	�'pe#1gV��)�G��Hr�9)	�'J����H�y���<����'	>B&(0 *�<�AC�)HFa�'ạ9�¤8v�|Ia�J3/�%S�'�-g �2���P�*��O���'2jl��W�$���g5���8�'
b��N6	���ǁ��*�z���'��9��H�-f8ef,X�8�lh�' b1��L.�����ҵ,%t��
�'���ӱ��,�r()R��+8<�J>���E�d#E�_�h�F��EG��'�T�d.�t�eE%c~�26��.��(D����霴x %A9���f$'D�����OK���G�
)�p	�c�#D���ӡ�J�Wb˂u,%��"D���3�#X�rɑ5)�LQ�p��4�O��!�bS�=� ��E"�/y�9��IX~"&�`�\@p.[&H&I	�y�hR)l����"�	-$+^�����$�y(ߙ��X[�*T#{� ��iB��y�b�>U\!�A�ɟ��4IDǆ��yBB8��m�u�@&uh�A
$���y�L�
� �y2�܉lք�bۭ��<A��$A�a��蓨�8��ke$J!>!��7IZD��%�)P��1tID!�D4u۾Q�mX)�,�Ѩ�;!�_!��[����UB�m?H�!�$ҥ@M���M�{��%/{�!�d�4Ra^@��m��(�ȡ�S���}!��L1g2�Qf��bN��3�+ܭ(�!��L(CG��#@�D�o�< &+W9�!���D�S�θ2��h�J�2;�!�
�Qf\!��^b���C#ǉ�!�DӘ-��%��*.] �{�oN�]!���B@���'�N$;�r���7*!�D��F�pb�	�g�*���B80�!�$*抉`�����|B�K,�{R�|B���qY�]"9�F��3��{+ўd��3� ��3�/X,Fuv���h�.�t��"O���q�
v^����cꎬ�C"O��J�� E��Y��Z� px�"O�Ik'ŏ�b�����1&�ҭ2"O�pg"�'a:8�b���1}�´��"O�9h�N�8g�^�i$�Һ��CB�'�ў"~Zw����љ@�	&7Yz�хi5�y��Oo��4c�:*h�m�&�7�y2%®��`J�<5Kޑsԭ���yBd�h��%t���x8�3/��y��v���P���V�H�B����y�8$����甪P0$�`�	 ��=��y�+�+?z:��+��BԾ91ѧ��y2�F'h�� ����<�[��(��>��Ob��H�oRrњ`"J�����g"O"e��c�x��c�5w��a"O޹��j��.<07�N�"��-x�"O"�%��h xb�0l�n�A�"O�L�3�0s��Q{V�l���i�`�'�a��D��)���%Úma���t"ʜ�yr�S:��Q�wo�k��"��I��yR�BM���f
�]�&�`'��y�� ��� �^�L���������y$�5GRD@��E�Da�UE��y2�P2~�d���Ӓ7�vY�E�Q��y��"��J����(,#��)�䓣hOq�%�����A�2Q`�1;�5��U����	1\N��p��M!5t�y٧ǐ'qQBB�	�[ZVq���иr�ʈ ֎NPJB�	Wޑ0DҬ6ޒD�G��[��B�	�e(ģ�N�������?<B�B�ɣQ$����b͟l��$Sw�I>VՊB䉸F_$��bY%Iu������u2tB�ɪ>}��eh�/;Uz���j��j�`�O��D?�6���k�L�e�c!��_+gT�� ���8?<���I�!��/�${ �K�_�Hp�q�!���)ٕ#r*(X�j�((v��t"O`p
!"�J&J ����&��+�"O�xp2��cF^�bOb���Y�\��՟h�?�}2e`��3ݰeK�M.�}Qa!�k�IZ�����y�[� X�70�S3E�4�y�H;i�H����.8*�}�@ �yR%�:6�r�[3ň(+�"r@���y�/� b*��̌�.l�����yҬ'`tV�L�-#�hGNL9�y"�!>����.E�2Dn`3G�1r!�$�c�	j�Y�6G�d��ΣB�!�P��wa�xQE�*"k}!�\4=�h�C�ܱv?ZXӂ�8l!�D�r,�"&�;n"��	_!�d�{H�$�R�>TxQ� 'oW!�dX������.1[~d��n7h!�$�*k�2<�7�U��x���ӭ%Q!�Q!6C�QD��M������}2!��:l�d�'��5r@��2�V!���)q0��4dǎpj�9r���-n!�$��O銙���|O����oR w�!�DF�d�N���ק2����j�!�d�+1\�Q�T��n�Q���.w]!�d�9HA0�(@e@�R����哪pX!���ò����H�MH:dϻ"�!�$ѭ*���a%����a����?�!��
�{^XiS�@
���r#7Xp!�� �=��N�^	���Tm�8�,��"OPmp�&Gxh��b%�Y���J�"O�mK�@܅w)f\ s�I�t�j��"O읠��71m&��G�88{\9hs"O��`m��f;؀k��( \l
"O(HA�-F�Y$\ᖪU1`AvBt"O�`q��#�`3ǈ^ x���jS"O>�KROРd��/�b}Z6G@�.!�:A�,�Ɉ81�O�f�!��:��0q�"�7d�	ǀC�	�*����M��05�-hC�I�^F���e�
f��ꔅٻSS�C�I�^������)�����G�f\lC�	�9Q����u�Y�� [�@C�ɰy�!�+-^���S4nR�e�C�	�ZՊ���#��戱��*eƴC��C�"�g_=T��zR�_��NB��n�PE!�G[�n�z����JB�ɠU:8)Ȁ"��Z����2,D.��B�ɐU��	H����s��d�4덐�C��a`����H.N���HBC��,K�2�F�U8`h���R�C�b#�(�̗�s�䁑�mѽw�0C䉛�� �7������� �z��B�v�1wB��6�X��� S5ŪB�	>M*���p��M� ���i�%j��B�:!?̂�ęA�,u��Ǌ�C�ɰy,�5*6hËB0m ���PI�B�I��!���U���%P�O�:��B�27�Da��#�[�d�h0mP�z}�B��+K�����[�R�rP���8 �B����4EFF��LYӇ
4%�B�ɿZ(���B*����ƥq�rB�	�s�~��& ܟ2AFu���^�M�fB�1"�d1z��ޓ0ze��.��B��/@������"x���W�f�B�q*��bլ�<|�9k%�2so�C�I�/��;�)U,v�Ѫ���_<�C�I�bd�r��*uS��B'_�NC�I=UD�c�)Z37���7�ޅ�ZB�I�#���jTI�=��T�e`[=،B䉧a�����E�detܲ�i�$�bB�I;�m�Peӌh�  ���E�6B�I6���A��1G���C�ʸJ�TC�I#a(h��u�R�}�>D��ǅ[�fC�ɨ)�H$�":�����!�C�	�"iԭ�&�7c�N'_���C��&x�^A4�͔y���@Ϣ~/zC䉖5��tK7��	��M"PB�B�,R���5 Gu �<�'��(V;0B䉀:��#�ZFy���Y�kg B��6 耀�CƇ.� �@�ڷe�B�I ^�D����)^#��hV�� {�B�	#�t �$̈�+j�HR$�6U3B�	�Cn�y�LO
GR���N�>=2FB�	�U�)`e ��\�a�P�^�u��B�I�u 2��^��x�Z�̝� ��B䉁fR�lq郴��YE��Q��B�Ɋ
1�̊�i�����Q�`[�C�	� �z��mG�Y����i%2��B�ɟ����A����,�$	5|�B�	�e�����FϤĹf(_�{g�B� N���Q@������ uEBB�I �.��&O�%����2�� 9�
B�)� ���ϭ�Pಯ[�B$�5"O�ɲP�+wp�<ږA����yK�"O4���E�2r�	I ���dC��'"O��9�'^'��ˀn�:{^�]re"O��	��M"Y�m�
�4\嶵k�"O�a'!R�l�0 B���mZ$"O4��)֊^��9�(Vl���"O��zS��u�X�ѣ�M�A�T�:�"O<�s�hR*)���Æ��!'D,`"O��0�O�*�uq����uf�� "O>�lZ/*<� V���"�"Ol���jM�T �P1�V�$"Oڭۢ˚�z�0�H�nI0�V�8�"O�$ r��sҒ�ِn�_r��3"O|X�A�(G�����^�����y�gCCr&U�ҥ̑o"`�����y"�L&(S^��R���fPJ�����0�y" Ġq����Ae�\3f�8q����y"fT7`�¤@�L[_��7�^��yh�
�`׍.�����N��y����(ÂH�fr���2|��mh�'Ƥ	P%L	<݌���]"r[����'a����f� Z&����dP�pdx��'�jA��A�錙��$uB����'M6���Ə�@0Q�� �#�t��'� @�.�5�}J�GɐN�ؽ�
�'L>A��U;BBtbp���v	49
�'��
!�ӧn ~Dl
�'�@�ڣ-��>�������z�= 	�'��a��
"y�蕊Я˥B�pdS�'��`���O�q���&���&F��'.$����M� � �G�$D"���'����	9�J�y�m�	��"�'TDy���O�!�OU����'����cĝ:C��LHG����	�'�0���ߍX�ɩ�k�r?jP��'N"�'U�.<�Ыk�	;�4���'��2���E��dbR,� .��1)�'Z�i�`�RF>��­ �'\bA*�'����f �d���q�\�����'�tB&ńwf�ʢ����2�'^VDX��݌Z�l����2�*�`	�'Dę��ᖎ��1!�Up�ݪ�'�L���C�X8�&l�Hi�	�',*%�g��1���sI?8�<1Q�'�6�*���%/�y��ʯ<��Q�
�'<t�$�� J���<�.P�
�'Z� B�63��*��vV�S�'�t@���H6aF�}ؑ��=�����'ΖhÖ�ڠu��-r���@)�'��(�@�Âp"�J���f���'���ʝ�'��{�:6�0M2�'S��*���`�"�blT?,����'Q��zU�U�7���8��0s�I;�'ޮ}�Ǆ�>l����ʯ'>a�
�'y� b���2A�Vp�v.L#Cf��'��)��@iI`�-���Q�'����D����"�B�X���`	�'�4�2�H^��;AeW�O)����'�N�#❦\��1���Z<$I#�'|NI�IX�]z��b�(Gt6�1�'c�t����By�LjA�M�=�|T�'��iڢN@� (���Ȓ3���Y�'��X1Ǩ����	�A���D��
��� ����aY05C�f���x4"O����w^B�+Pa�&  ��"Ob���
W�@��A�� }��)r�"O�`�%LUgE(��G�ӆ>��� "O��3��G��"\kE�&E��4��"O����Ȳw�P�����\�@(�%"O>�Yjނdg\@q���4}��!٦"OZ��/�9@��X����t"O��i]R������=���"E"O�H
��3*�̙p%�#U� Hx"OT|h�,�� �X	���Cɀ��\��F{���-ph��U&�!��T��2-�!�DV^u2�1#H�>�L0p�@@#�!���s�&�;f��f�L�%/�{�!���x� (��H�o�����Nĭ!���q�$9}J|�':@4�g@�������p�(��'�J ɒ�8O��t��G��c�6���4���A��@��!�?�xh3�LJ�",jL:D�,�A�Yʈ��an%d����c6D��C"��o:����Z,)�ps��>D�X1�؍cW(�"�Y;O ����0D�����][NT��m@hh�Ь�<�
��v�p��Z?�$�;��S>\qJ�G���h�6az���(C �[�H^5;�~C��4c,��%4��l��!�?5]R��ē���S�,fչ�#8 v@��`��m"C���q�CH�9a>*�s�b�@�DB�	?u` jE6_1
���C&�.B�'Z�D�T���m��щ��BdT0����h�t�>%?�"ǍA�>�ҽؐiZ�{+D�U�<�O��'v
�W�� <p����J6-�d���'�Pt��/`n�8���E5�L\���d8�'~����'�
G�	@Rc)�|��ȓ_�1��7n�4��IF�A��܆�,�©����~L�%z�`_G䍆ȓ��ȑ"��p
���c♄ȓb�e�p*�%&��f�Gd&0�ȓol�ͱ��J
t� j�KϹ���c��?,Oڬ���X�!8aU(A8vԴ�b�"O�,`"*�,�2�b! �1h�!�K�_�<�Q�Q�=OL|S�+]h�ў|��ӄ�zt��e�	fГ�DʀC䉱8'��+��F��*@BF�r�T��?�{R�	�'7�ppRN=�0<�0��%	BC� {Q�x8��g�܍�DZ�L���n�a}��G5{x*�B�#��X���<�K�ؖ'Z8�˶��(��TO����c�@��y2ʉ�������@�  ��(ިO0"�d@�0��0��"Kr��p���e�<�Q.ؐ\{��b�"Xs��h��W�<�bJ�()X0(q0,�4��X�SR�<y��	�V�f��J�T�Q�C�v�<i�ȗ5$��!�e�!�0%��aSo�<yt�ٮ�v���X�q�J�:b.�l�<��� � ��I�i�����h�N�<i���,2r]�tC߷5Ah�����t�<�����L�2���_ͼ�%fKX}"�)�'4Z����*���
�f�!,	����[t0�z�鉌0[de2�ě�r�u�=Yۓ{=\Z�j�"j@�3�ĕ�)���M���R:I�#�	ǧn�q"/�~�<�����B��N`H,��@�$0�Շ�K�`�Ѱ�)kp���m�.*3Ь��	\�'�8$���J�^(���
X�j%8�O�-�O� A@��!@�*P�RDȥO
�43O���J�S�Ov،�Q8��#5�6v%����'����B�7$�$����v=*�(OJ��$HQ�b>�@�ݣ!*���`�8ud��<�O�`�'W@����/YV	)%�	2���;��yy��'}x ��Z+.}9�`�x��Y�¼i[���O���H��)��u�׫�w@��z�'$�$����5$�1Ȧ"�@�"@�,�(O?�$�/�Ɂ
H�
{fY����?!���g0ڨ1�@<i8��Cʻ)���=O�i��&?�"ƣL��U"O~�@����EM�5)"�M��9�$�O���o�g?I�.ǲgB�������T��8���9�y���2Ҋ�`0(G�NZ �	7`#��$�<�H>���ɬl�d�y�G�KBPDsc�r�C�	r�e�EǗ�l� ����
ѧ�ē�p>�'�
SK�d�Q�P�C�ƞu8��$��'njI��d�%�f�I�^e{`�m�<yT'�(Qgx�"'+2Ƹ<����h�'� �F�4���3�h���`�N x�E(���yrÀ8�L�z���8S���m,�y��Va�T|�Ѡ'Q
���u����y�kX�/��i�̑#NA%��6��D.�OX�VZ<f�. ������P��'��	� ?>�B�+	d8��`�⎧�rC�	#Zb�ѳ�B�9(�����F�0"=���T?=s�B<Q����(}���P��"��F���'*JV]�U�#m�ƅx����( �H���F{r䐋`�Ё�'��=6+��ɥ
��HO��$�MSmX3E\�_�q�U �#,�!��hT+�H��{p�pwOX$��hD�ԩ+}!��zU�	 �b�ZG�S2�yr�B�PV6��c[(�Vl��A�y�l� %D��#ӌ8"X���O��ybJR�$
�9,�&���V����%�O� �\�O�h$3D�L�
i*�Hc"O���Ξ�G5 �����,t_x���"O�D��͝<]f�R�o�>1�R��"O�%���A�m12o��`08a�'Y��OLԨTM̕kJ��!N__��@�"O���'bD$s�tS��D�(f�s"O �r%�53��1ɖ�H)f$��"O�)b�	� |�`�P�u`��X�"O��{�$�
H�b��a�à2?v%Ӈ"O���	��gi�ۅő�mB�8���s����j�E�4�D�CR��sC�m!��M�oj�b�rY� pW⇤�!�Z$��Ձ߭@���p@ԡ~�a}ҕ>�E(�I�
�(�o^�h�s����?�/O����(l�x��/16�d�r��:]�!�DWPC.��#-h(��֪N�D&!�$�v���ۃ��\�"]�	��IhX��&
Y&�P<� ��j\���e+!D��Q�O@jA�pF#>-R�{�h)D�sugM8�lR�˄;&�h�H$4��C#�,U�����S�p�lC�h
E�<�¥�B n���$�>A�5#Cc�~x�TExB-\&U�͎�&*�,Z!����y�V�c�MX�Q5j��mS��y�� 8�9b�\�,? =�����xr�ii�i���߻>��mc��I1&X�6Y������'�v�>�w�ۉP�	�B�гP�@����'LO��#zyr��L�19�`*`@U�:!�'t����	�?��xJ�ܳ$��,S ���D{J~� �����{���W�ΌN��H��"O��p��� ��A�-�TyV�R��	}�'��ɳD��5@5H!Q�dis �N;�B�	�g�V	B������,�%h�B��rI�]#��N1)/X4�+�.d�B�w8�Y	�A�e�L,��F�X"C�ɉT/��Z�M�E,��j��"<q?�S���Y�IP���gR!P����T"���yR�F;/v|`�Z�_�*��7�=�y��)�	z�����X�Q�U[b[0��ȓK69!p�"��!�s��M��%��R����R��$�^�� �*a~�W�P���7
�xth�l+d`�c$D�L���:B��h�G��2��5S�$0��{���';wҥ:U
S	\zp0�"�:��ȓ6��4`�d֜\[��-��'����J������p}��;� O�"��w���1eU$f%4�Cר�J<���ȓ1p�D�5���+��%;:�B&"OI�e*
(7���$υW&��#�"O�8"S�&��р�0A����u�6D�X8��%U��PR7��I���S	5D�,r�J>"*  e���礜o3D��u�B�t]�,ID
<#*f cqa,D���WN6����U��/T@F$y�+,D�<d��)V���*uC��u��ɦe(D�`Z�I�
&@��5�m޵+�h'D��
T�R�_��)#C��3������$D����H�0uziƃ^_��Q�3�$D�Da�*I �H�2f�F�{�~m�B%"D��xE��C��qD�@C���Q�:D�����	B�|3v�
���Y��8D�c����%j��҄:h�A�$6D���� ��(QhU�w 5E�� �5D�����X��NF�`iz���'D�ԛ�&�6d���9���j+ qj J8D����F�agJ�ԫ�]���Ja)8D�����Wak���I��7D��sv�L�y�| �_#Dt�"�M6D�|�ԍ�0*�v��ě�Ql���63D���%̞ R���vE�9a�@���1D���w�� k�`��f@W*3��,�'1D�Ȫ1/J!�q�2�Ӡ}w����3D�PqQ��$S���x�+�-Zo�0c�,7D�����<V�Pi0��d<�dF #D��(��]�!��3��x:Jx !D���w��8�LR��9����<~�`�p
��]�#
 LOt��6MB/t2���I�� 	Z�BT"O��* ��2 �ɴo`x�"OEp-P�R��@�l{^���"Of�J�-ѽ�Z�CT[�[�i��"O��b("��Jc�_&P+qkP"O�Ջ��V3_�c���z3"O�`�n�o��U��d�7��8`"O�p{��@'H��́hy�؉"O����(>$���ϐ�F�$ڑ"O�i��W):�3�O\�1�6���"Ol�C��"K�q�7nJ�
���"O�ɐ��U�2QP���D�$��6"ObP�gL�u���3NBxvv0�a"O��c65"��Ȋ�PTy��"O�0V,$A���Q��=^^nĲC"O*M�匯Q��Y'�VATq��"O����X�b�jhQ@$�,X�l��"O� ~�ۥ`ƘF��a��	4$`��E"O�؃�?zt�t�6�D0@�"O�4��R�a�2!8�T�}�@�R"O�D��H� ����S�C��$q"O┐���i���K��Ǔ/ߠ��#"O�J3"�3Bhl��Rn��n�"p�"O��p�O�Y��ã �>&�Źp"O4�r��Xy-�I��6;�P�"On �e�N7k^e{`ΡO'xXK"O��DB��:�Pggø0K��S�"OB��r��H H;�L�+�J�"ON�� -"אm�b����*U��"O�@2W��gT)3PԳH_�}	�"Or��D��5�J`�5
�+f9"`�"O|��p�ɒA�<�P�V�W<lX�"O,�	]���l�1�s&��p"O$%�(S�k�ҹ�MZ�ic�0�"Opm��Y\�;��S7o�h(�"O����A����"G)�)~y���"O.Uڶ�m.�����g��E"O.����Z�k��X�2F�N�h��"O��`��3�d����Η9�b4c�"O�U�0*K��\8Q�dI�A�,���"O>��F�*kDڱ � �:YxhM�V"O��iạ̇̄
�"���ܴfh��a�"O^U���%4�ᆛ�[Z�Rt"O���&�g$� s���R�$�{"O>5�&&} hu��L,2�j�`'"O�����X��U���G����$"O\X�6�zW�-�R�P[�"%�b"O��C�M��1O,�
�I y���S�"O��EFN�$��&FPT�x��T"Of����M/��c��0�H�Q�"Ox�4nƧc�¸�C��8�l��@"O��� �U�"�@$����B�:1"O���n&F�h�h�>v�朲�"Oܙa��9z�0$�g�X*�	@"O4E	��L#�6aY��T:Eʶ"O���KȨ[Ѩ��3��m\��v"O�xh$�'K�(�+f�R���"O,��a��F����(9<��0"O�m�S�
-Me� #2#(��U"O��
�ER�x @�Ԗ�7퉠�@q���S��!D�](x*Z5���/+��B�	5md�%	bn;���i��P�f�!�`̡��0}���'�`X2,B�\-��J��[��U�'�
�+�n�<d�@\Y�f֛d�*�+�"�B�[��ĔWm`�YV�",O-���m��H[�.������'*m�ECW~� r�CĚh��x�ǐ�y���O��TԠ��
O�ة��˽E�qy���8����T�dD�)�2yGη,�8��-�S�sx�I��:A��[��6=HB�	��r�U��]j�SFH�,u{�q�G]��ðֹd��Z�'���v�M~n���&�ѿ]>1���^�,��UKw�Sz�<!�ތs�Z��4�)ADp`����:R���0w�J��Z��7Il�oڽ℩�)S]ܓ"�P�pT��%|�@:c!�,nz����I�c*��F��8��=YB�"��s�`P�h)� *|�5��a�WL88Eo#�����tJ��j��H8O8W�1OJ4:B��S�
 g� �Z�J�����#�D,�9`���	WqFLI#�@�XD�0��<�!�F=Z�&����Qe���a��{�n��u��+m��IՆOcf�JG>\�2��!�?��3�t���$Y�CC�PeeK�~P���-2D����(4~Æ)*���)\���a��(��t�g�##��I�t�ő�5zɐZ`b/�I�bPf�"3n�\�n�HE�����L�<t��!#�'d�+��]��8���N�3n
�y�"��*�b�����`C&љA#��	ӓP�X��&�	U7Vu���[
��'�j��DA��v�A�
v΀s�J�+O:�T�P� PH�u�	����reV�!s�4"O�D���K�o�$��sN�
az&1[��H'Z#�Ę	��=��8����g�X���n��d�b}(-k�1�l�́{�А�!�x R��'��t�Q�R��E�oάn�>��掟��]`E��+����6�n���ѡ�i�A� �^�_�qO�������u�!V8s���J��n�'��-��/��]�؉��j��<�����	̞�\�(�IBL��ٻ)�7&���i��'� �n=�p=11��0w�(M���C�b5�d"�BlyM�
є��ɪ�\䫕�\�H�vh��O����@kĽ^��j�v�N���L�$�IS"ON�s�;i:�V�Ѵ8����#T=3p�K�fӍb�Y�S�ً_>D�o"u�p��[�����/�yG,,���A1+��Hn�h�Ǣ���?� �	)cj!�N���@}���ӑ
%��(�旰��#q�7J):�@�j� �P��3�Ji���|��2��!9B�S+E�n9;'ϐ��O�ز�ȼL��Ŭ\�=@�u�P�̝u���{!)�-59q	f%�2;���H4b���ʲ(����Ĕp�Q��N��bc�`@eO��2��(Z�����Q85$\}��IL#��"I�*$�x�㑰J.�tfH�N�t���wh<���0df��x�.ǌO>��

F�'�Zu�& Ԝc��D{?�`�+)�	�sCv(����+q9@T�B(�.$!���}���R(R�O]H�'K'_L�7��(�:-Ä�d�p��<AǤ�n_H����j��]�M�d�<���]8.@���N{�0y��:@
���%���R��M���<c�� 5����4,�UZ�4����v���1)��-A<�!M�30�l�JQkB�g�N���b=�"��64�|�R.Hl���!���%�x%��,�I�x�ɩ��wF�xC�-��M��Ii萺G����@�8O��B�	�r|�5�˘t	�|Ȇ"M����J�A=]��G�B�$���(��I5 ���	�aO�IJv�Ih��C䉺o��6f´-ٖ�
C�
�$�����J��ji>|�2��1��z���)��)�E�Ȁf$DX�p�H��p=) ��\> SrLܢ�M;Wl�>��PFF)x;�	�V��v�<9![�ݨ!r�(Ӡ|�:�Ӷq�N�����l�i0|G����6~��ڂ%�8��[�ٶ�y2I����q�I�(n�^�iG���x9�!�]$���'�>�I,�����N�_�t�q��{�C�_�L�'���~YhP׬Y����D.y��|A�K��=�d�k����ɐ��do���0>� �^�^$��*dJ`�¾kM(�r�GZɖ%��Z���$!V4K � � ��N�QDy�	�[� �F�t��#`�L+S!^�FN���ȹ�y"O˿|@1��9H��xiq���y�E�E(n�j\��m���y�嘗bW��*㋃�Mf
�k�)��y������c�E�,�H���f֭�yBm��K��|�`('5V��h� �y��̀~2VD1��?#�@r�]����'C�r��K1B�4 ��m��L>�S,թN�$�IV|=)g!g<�s���;tP(�U�yB\�*�◂E�"p�C�G �R��D�.p-v!PϓEn衔�e��(��\�E��U��ԣv5�CƁ�j�!��U�^|ظЂC�
�]�w�^H<����?���(�OL�f�\��3l�Dy�#�>5�E2Q&O�a��A��5q=��~zDM�5 ]& cI'k��P���G�<��*���Lx&H�#e�2��C�����0nχa��-Rvi�
:h�h&?1zV�x�Ѫl�X�wfP�%��j ����?ك�Q���=�ɸ�NɩN��<A��$R�Zh�@l��螀���A��@���~e@9yD`-q�V*��U�^ >�?���W���;�(M<T�t��4 ޛS�M9�
�p6i��k�6{����&�1$�̋b���:�[��BqЉ��<��]&o���.�,_��x�G`½��c?�$�D�$����%CL޵��.4D��yw�S�+6$�	��W�Pc��$-�tA4]��Bs~t�+U&��CԌ��~�#M<Y%�L�X�� *1�SQ�б:Q+�m<QhB{.�J'�������9oC&�
�g(vw�p1JM�#L���m���
�EÒ����@���IIz4���_qD�
ۮ=�4��!R�A}��� ��U�ޑ10"Oȍ��B" /�L	�eQ3f.)�"O.@0�Ϙ��bd[U#I�li�@�E"O� f����׆1��+�W�U�c5"O�Q[6l�"#�a�n��C\t�rw�'Y��ˁ����ɵz�$����}˲��d�	�6C�ɴ3��r����S�*=@�)O$L`�b�8P���Ne�\+��S)p��a`P�_7�ҁB�&�BB��=�6����
t7���b*:d�K`�S=���e��!��L����������ا,�\@���/4���U�U�)�B�zo�uN�^L��1"�)�6a��D���f�$~dڠ��̓&_���M�}n�L�%Z��	�>��1/W�؂$�vO(h�B�Ie�*pZī��8p�O:J邏O�,HG!�9L༽i�"�f���Q��R< ��t!Z�+�Xm��g+R�jQ���B�|`Ȉ���v�T��B��'< D��>�gϟ+e�Q9B�N_��� �`h<a5$���<�+���,8���@�-TG^)�Ў���T��
�{4��s�ٯD��H�AɅ�z�牯E��T�w�	��~�ΓGk
�B3�0\��д���S�"Oȵ�#AY�t� �A*(�R�	���**�X�!� ����
ܩ��Bjx��ɀQc��
�'�Tx�fW?i��!�	X�fv.t��oDr�O,|��Y�4#7�Ͷeݾ4�5��&9:��!D�\�'�H|@��)��'8���C:D����|m�Z��ț �����9D��(�@/`�z%k��P�yP�0�E D��#f+O�?��ip�ѳ2 (D�V�!D��ÕJ�*�8����"�H��+?D���B*�1dn���C�ub�y�6�=D���`F4[d��Pc�
���p�<D�$�F�R!Z,ڥ�4�F=1,RPZ7,)D����-�N�� ��!T��3�	'D��bSK�n��  ��<K���$D�<���:A�J<(�ȑ)_`����m1T�P�t�"�d��F� Z���"OΩp$B�(g����x���"O�XqeN9]5�Eq C������"O@�8U�(q[xm�_9(�� #"O�$[�B�7?��01v$W@��Piv"O���f��	9kzy���O�x��"Od��#��a`Ri�b�;N��uqW"OH��#dJ$u̰S�R
�
9h�"O��!�R�q�,x���La�� �`"O����ę%Ot �d^�E��U�W"OV��$�4�r���Y�BK׌6�!��,�4*V*�*U�Z�Re�+�!�dk����D٩�6liG�A�h!�d��L����q���h�pp*�"λg�!�$ķLt�P����{��5 �=	�!�D\�tnB�A�:L3��ZN��!�D�5q�Z���ݯ 5���EN�R�!�䋺	̠XJU�J�d2�y����b�!򄍼G&yZEN֥B2D�o�e!�D�s�y�*�/w���YA���h)!��ΌX����ŏ�LA�]�U��!D���g�Ɩ7���^�t�2��U/z!�dߝCK��i�)�<�hm�č��!��v�1�$g/U�̐U%V�|�!�d�2dCD@���	,e\rhr�KA+�!�DC�J�J��ɪ[Db�2S
E	�!�d��9����V�JHr��c��]�!����Hf�$.I������+�!�V�b��R���\"Hx��iJ�k!�$��rY�QI0/���(C/H!�,sπ�)�@E(M������,n!�B]}�E���xZ�Y)���b�!�� &qS��̸��� $�<Ŏq�s"O=phρc}bU��A3m,m��"O �f�&*�}��)Bl�1�"O 1��LT`�t�5l�J4�%"O�x�*P�X��]"�b��I�Ř�"O0��b�X�eX�9c�Z
�lt��"O"���Ŭ&��B��T��9��"Ot��7.�p��X�I
~pp\Y"O"Y���ʒv�(��!� q��q"Or�J e�3z7��V��Ujx�j"O:��4.��a��<�b�ŭ0���"O���L�A�$S��CV�!a"O�AbZ-PX82W�S�J�ؼF"O�2p��n̻�
�1�| �"O\�9aꎩd�`����
��)"OX��ɏ�{M�ZA��;���P�"O�`�f�LC�1�Y�}�^%
1"O���lD�؄��!W2"���`"O$�'�P�q�$Q���R�ĩw"O0��fK�NՖ��f��@��JT"O��BA*O4��#l���d�;�"O�8"HQ(_�: B��P6r���E"O�)�h�)Z�@L���(+�Z�"OZ�����sp���T�����X�"O�I�'K�@�F�[rc\7[�Ԡ�"O���p�I2�@)$�.`���U"O��QD�I!T}��^�$�:鳣"O���qjS�:0��6�Z�\����"OL032-�!
DiA���6�\��#"O<�k�b��K���0� 'SO����"O��� 9�z!2a 
�67j@3P"O�1��o0~RS	�c�|��"O`-��锫4(.Ջ`g�*M�$�"O��91!�=~�������N�f��"O��@�׏	���*S�+���T"O�%�c��U��QP!AؠV��\@�"Or���*��w�	�$"4�"O���Y����RNE {��"O�{FK�i����®��:��#F"O��Ro�]���� �
3�H"O���L���P(���56�f	�"O"]Ck�%�L1y��)$�2�ل"O<�v ��\\���9��S"O����h;��9(�L2���[�"Ozy@�h��j�D�`���9g"O�@��*��$8�A(�.�m�H��#"O�B7斩Io8��-��s،b�"O��:v�_�T�ġ����+�n�sG"O����*���A2P�^-��"O��)���2<�hsD`Đ9�L�[T"O����=`wp����B$w��Y�d"OX-�CL�7#���A�X#.ǒm�"Ov��d�����2��/#��q"OLdJ꒳d϶d��F�5���6"O�к&+h��;��D0&�.p%"O���UΏ�j>��_�ɱ�ՔN�ў<���9>k�>���!Po������;����*1D��6�۴*�����C�6��ɸ�Jkӄy�eXz��O?7�����EK<!%��Y�{(!�,k�V�)�%�8
x��3$ӧD����).g�i�O�0=y��]-^w�Xq�Y>u�}k���G8��Q���6� [w+������V��9�fhS�K(q�!�D��BH�a�a.E"V��q�$�ΑR��a8����V �'E@��f!d`�'?��;q`����H�b="��]7G#�Մ�S�? ��ɠkSt���h"ǔ�k���ɳc��*ag
�&uD��O�`���B;Ubf ��y�m�qwQ#���40w������p<id��"����cקlGvh��L f[�)H�	C̾��ǨW<S�J��:rI4(6��D�azb.ű
�J\+&�*�E+����dP1Q�S��>�܍h��҈i��i�<y1��_)�(��P zЌtd �d��C�ɓd��H�����D�B8�b��i]d)��&`Baq�J#/��d��Fg��P����@�	�-5�21GV�@5���t��V��/��"�35M2�xgf'&��\"��V�
o�v�S��gi2)	�K����\�H��,k�i)�={�vm2����,��͑�Q�qp��?��)и$ڪ$���G�AO��I�/ީ\�V�H����o/@��^;���-O��h E��z��z��Gd�|y��V�Z�|���)��XvTqR�=E�<!�`�8[��'M���TH�G���[q�5 x:��Q�B6@)����'+bL*�I2'òA@�/�,.a܅J��%q�J=KR��������F�*.n6��fL�םJ}��e��c���\��p��o��:���˧�>�O��S4�7~z����cO8e�gɱ�X���0�a�� |�}ax��Sn���'���)�CH1�|��$��d�`p
���T�#�> �e��gH���id�^w����U��&�3tn294x��O2%�𯙢u��u�	�dm�:�`U l)dL��	��0�n��'�Vذp��L`ɧ� G� OfL��G�̣^*�0ZC��6tP�b�Y�Fw|��O��`��D��pA��h�8�@�d�4}y�HGl�8��O�1��hC�|JeȐ:�
HįI�O�:`C�r�<	�� �q�f\���U�ܰrMτS� l!���l;�A�'��XD�,O�( �Vm>���l_�-���5"O
}�rO���\�%�we���P�+�4����N')VZ�H�!<O\�	�f
�B�x��π'�P����'���c 	�.-�Y#��P�A�\���EF�:^�����w�:q�',�qS�jӞ Ȉ�UI�/&����{Fגz�u��Z�T��I���G�	%�p�'��_{�t!G[��y2��!������:%�=�7,+D�T�q�
X8[�¡[�'[R=F�,O��1�@,2��N]�yE:���"OhոF�
d�kt�+p>t��֍9gD�6gкC�ڱ
דS��(�T��w�t��S���&\O@�J1G^+��E�!
w��1��:0Fp {V���]~Dp�"O�D��@����Q�=��d�Bvu��	S�Ox�>e���]_�}2g���S���2D�6D�������TSA'� J�QRD��(w�1�J4��	o��~�éI�rY�%��0G01�g\��y2�T�r� i�I��c`r�@Ff�
�?qG�e�
�&'lO��9����B�:��w抱x���AD�'V���N#C�Bb�A����+�!d�������yR YjrJl!���$������(OȘqp`٘ꈟ��që8,�B��$遃�N���"O��bg_ċR������A`"O�E��̙��Uk����GLԩS�"O 	ʒ� ��������f�xR�"O��kN[� �F�[ōҟ;�}�`"O*A�wgQr3*�A���?t��m�"O�4P��  u�(u��'I�} 7o�to�pG
"Q�:|�
Qq�q��'W|P�G�&"&��2�N�4��'Vx@�$,�>F�Q�#�G�/�.x�$N��X���K� $=Sz$�H�&O��yB��c�(49q�K��2)2�k����O�e�� ,{l��hP/+|M�Qf�yP�L4O��xh�v��/02��'N����]C:4��Fа;k���.OT�P�D�����J��#��-+W�ő��O������!LB��F�ī3���;D��+����E�p�@�N[�<�y�hX�4�<b�2⾵����(�������K<A"͔7qS��)$��n��4��&�g��tjR��4\�!��@ʲR�45Z�Ě) �� ��X�0R rB��*��'�\1t�Еw�ҥ��(��U��J�����@]�*7jO�FXE
��H�7]����-}�z�����!h��pc�ɼ�xB�O��@#�-o���p큄��D�-�$��RC�����91������D-t0�գ�F+5_�0
2�y�(�0k����a�..��)����>G�<��m͝�b��"�x���KL~��<��,t>�;�郳`=&,�2.|5���[n��1�Jn͌X`��Q-\�$�A�Y�A��ȆL�6X�����<� r�!2��*sf��`���l1&�'9�ĉ��Jl�����]b�H���ޠ������ѢmT*,%%ZK�<Y�d`�]����	.Ļ�#�@�<!�2��a�iB���	`��W}�<e3ghB!Z�GK�]� Ly�<�o̍~����N/%0P�I�������	nD�'q�)Y�%=v������1pt	��'X�Ā�L�5	�(�V�J)t��`��yB�J�v��t�ƥL�O��y�/�f�Q3J�S����'�L��O�<��My� ��s�$��4�\��%�+O�ջ�2�3}�B�cd,Ōqr4�'�����x��vtP��ՎL.4w �sunV:Q\$!*�G��[���bS�'���q� �V�8�Q#��a`0\XϓS�𑣇�gj>HH�'�,�rf�]:&�*�;�mQ�^�a�'r>�!�)U>!�J�������zJ>��������ӈ��%��!'~��p��ڕu>*��F"Oؙ8��5|#~� O�� H�@���U4DA�R�(1TBD�g�d��|���C��XMf�R� �s%��D�!�蕁��H�uKd�ҰD*A<l�P��]���i�&�O���w�O�P2��B�?��@"��'Q6��c��<��T2�3O�Y�`�1Z$�a�D� s�+�"O�����\b�0��OǱ6f
���<��ݾY�HG����Pt���T�׾s7ƕ��]�y�D�Z�4"�@��^'\}B/[�$bN��e�!�ۭ�(��ɪN�㢋_(��Bq
�i#�C�	�T��a2�*΢F���BmS�[�TB�ɗo��QVb׺Bz�CҬR�'�8B䉒_{�]PT�L�!�ܴ��ǍG��C�|&��y��Y�vD� S���C� AA�T�� �= .�z�H�e*tC�I#%���k�1W�Ӌ�60NC��3�"��ř���!��2{C��%+�eʱ�C7X`&$�^Y�B�	����W�@�i� t����(C�B�	��	
�ǘ:m��������B�	�˾�90j�	i��i �"R;"�B��	&}X\��?<��@B����B�	N�t�n�/b�Q���i��ȓr�hl�e�B"G�R8��l���ɇȓ{N����*O�ab���Ԅ�ȓ3A`���:����L-����9B|9�&�D9���g�I;�*���Z�ĐסZt��O[���ª���%��oȀ���/��x��^ՠ���K��
Q�U	@]���ȓ��C$�_�!�L�A�#4�D��!��(wi	�Y�΀Y���xɸ(�ȓ-�
]�T �	���Vڹ|fZ��ȓ)*DB��G
.M�5�̶;�b��ȓh����O;4��D�$0z\��ޢ��`���c�Zq�a͙�GX���p��ud.�UE�99��XY��}�� ����c!$(��9Q���ȓhL��c�4�R}�!�_8�Ze�ȓ?)JE��θ:Um�:놀�cB�����S�M(Tڸ���Ɍ���K�E=[�O=o�C�6���h�Io�6���')+/�C�I�aVv̘0cǁ@~uZQ��0M7zC�+/
Hl�TN�����صJabC�	�.�����ͤW�R����{�B�	#r`��Kd�_�e��D�&I��:��C�U�%�[�.4Ա��L%xuC�]��7�
l�A�VY�t�Ny��'�L}y�����{�B[�'T� P��Q��0�v�OE���JE�H�%�>P�zb����� ��Y�F�Vst<�w����7��]?���>��4E�=�0|Z�E�XG������=-,��Ɯ�-�ˈ_�T����%2���)§��dŇ�Q��e�!�[�"(`���3RW~��6c��p0�b9���Yi>%���,F`Ԍ�$�;(���sF�M���jf��Y@�f'ő]}�,&>�}é�00�|��b�
�nh �8%�ڗ0���Y������,k^a�4��;DNXb,Ѣ�J̀��3w��	"E ����M�g��S�'��PQUh=)d&\�0��Y��m�Bz�M)#��)��O�3}�*P���q�[��f5#w�Z.�?	������"~e&٣#�܌�U��l���ɀPg�92
�'g
\��"�
���}j�*7H��y"�U��()0)��"�0�$E��y�ǈ�%���� �@�f� "B��y���t�hibB��:�n�b�l��y�o\�S�� �d`��Z�Ζ��y��I&O�QC�T�PD!�W$�yriP�Rkp�#PO�GoȤP�^��y�ŎW6�ÆE8c꩘s���y���|E"�'f�����yRȃ9(jf���K�ؕ����ybl�,����2I�-�jY��c�Py�'�-j�$=ۗMQ�o�$qz�@�<��ҸJ��]kfJ�>C��Љ�T�<���owv�X'f��#�pٖ�P�<AR�+/��v�[�'H��Z�Q�<)���0Lʹ%��eW�U�P*6D�N�<Qu�Cc%n�I7%��-=r9�nFa�<��X�2�-�S�%��)j��Q`�<�ы�R���(Q�CL�	ԃ�Y�<�2J��i��t$��
Oi�511��U�<�$ �%J�l�v�	���*�]�<�a@�@����+:�L�0'*�d�<Q���7F�P]৹B9�e�Ŋ1f�B�	�ag<}�%�]����#�D�I|�B�	/j��#c6Yu6� ��0�B�8�Lܛ�$G���������O̒B䉣;�b|�s�@�q�tt�E�A>h��B�I7D�\��#�J�^� ��C<.��B�I1d,��@�V�MvL8�uc��.{�B��.8$�� ���En(���$Ҁ��C�I*"Z��@i�}{"�X�AN#�C䉜JyȀ��h��RS8x����\�B�ɖ	����2p�e� 	3?�C�I Ӧm����iNܭk�%�	-��C䉓� �`�Iȹ��v �C��"T���`O�<�����[^M�C䉔D}�i��\<"�XH�vB[1��C�I9I`����J�g[�x�)!:�C��2��L#�`]�MB͡��
r��C�I�Y2+F��^�8SAF�)V:��'m�A�NE	�x��h�H��H��'f�����L�8�	cCP�E�.5C�'��q�����eF� 0R�:*_z���')�h�!�J
93����n� c���'���0m�m��y�@�V���y�'���KehO�3朹��F:; 9A�'���T�K8*FXD�҆,v���'���eW�H���bC邷T��3
�'+rx�"�)�����T ���r�'4�2���l�(I+6�ߍ_����'U��Y�a[:!@�+YT����'���3�@^��k����`A	�'�6�����O|�t��;�1��'-�ɠ/�%8�yP�nW�;�<���'�cSD�w��\%ޔ0e������ �͊A@�T�ƨ8CBT$67�`�"O�s���)R�j�� оa")
0"OL-��5 �J��N�
=��JC"O��b��%p�����"#�Qp"OA��GK�0�ݐ���zl�"O�hr$�<0i�U�H<["�X�"Oڌ��J1�0B��$ZP��"O<i�	@�>T�e�(at���y盇jLt���� ��h
0���y�N�d��pY� SG�v:gA )�y��q�J陲�
�2�^�����y"g��^���˘�W�)P���yb�¦���A���N]>��A�م�y�(B3��,*���>*��A��y"�_ a`��{�DI=V�����Q��y�J��3L�0�BY�`��a˜�y�ճ!\�(����2G��yB�Ϳ�y������,)dh�1֨�sRÝ�y��	 �%a�@H�, h\Af�0�y���M��P��	�8$�����y�aD�E�f�80BB�6j��K
�y�&�7hܤ ��e����pxW� 	�yR`�,��4���+
0��e�_��y2�ˊ~"V<����U���9E�(�y"/�$H��R�U� �����y�P�46�PAifI�L�0@E�ȓV����G��d�f��m��p\�!�Ũ�en�*b��?[E&9��uV���g�(@��rS��N�<�ȓ	P��"�]&F��-���֤z�D	�ȓDHp,	�  �s!�i��FHyz�8�ȓs)�t*�%��$K��Xc���G<��VkF�H"�`%����ȓl~,i��n�
�b�4�ˆ>;)�ȓ�&Yq�#�lA�@H+�$�&��ȓ	U\s1(�IQ �+�·{��}��goJ!��`@�F�I��Ǳ'"�B剐g�"i{dO�iִt1a�& æB�I\@H�4 ��,�XhrS.7�B�	�6#b��NA�f�P1萴.>�B��R���*��Ƞ$�7D�]f�B�	<���V�DY;���ӛw�xB�@�(�&ַkՂ��A P/Y�lB�əQX$K�cT?$���-��B�I�e�jl�W�W�#����V�T�t}�B�	�g���ꔧB;�Ї�*��B�I=etba{2c�Y�"�q hR���B�I.Z$��zv��$/��6�.<�C�ɯL�D�4�C�j�5*���DA`	�'�$l)�nȶK�E#�! tdY�	�'��\8��ɟG�f��Kt��	�'}�5z�'�*k N���N�2�
 �	�'�,=�OD�#��VP�SdP��	�'~����aI���f��R궜"
�'`ZEN[��^uL�2-��'�0��b[�n)L̐%���>�h�z�'+������8�H50��<XD��'����A��-u���/## *@Z�'����e��:ԭ�+��$�t�>D��{6�D-��|�cmũs���Bb:D��yP�Uv��@�"�ƎiP��+D���͇c�V]R�K�$VXF|�2�*D�T��A�gT!q��_�~�:�	s$D���	S86�f�afd�&pM�2c/D�� �|h��<8����KS�u�:�1 "OjMs���\cd,���!?��Q "O���Ѧ[�r���T)��|pg"O���BZ�(�PZ��84�@"Oܠʷ"$j��5ڒ��ܐ��"O�8q�Ɂ3d��x�����Iq"Ol�Æ�� @�$,A�w�$�"O\�I���9�p4��J( �6�;`"Or�y�Gˍ{�$x����H�N-9�"O���3A�,
��)A&:	��p5"OV�3JR�H`����G�Ľ,�y�JZ�6P���̵L�>��%��yB
]cqj�"s��Z���eH�B�<sZ$4�̍��ʝ�K���P"O��Q�_�Q�p�EW���� �"O֝����?C�j������@H�!"O:\�'��.�����->@k�"O���Y	]@�H0q�!z��8`�"Ol� D��!)hu l[f
@Q"ObIRp��f���hw	��Q����"O�E!&Y%��9R��>�d�@4"Oplsѧ	�. t���g��?Ƣ�ò"O��q��v�21��֊9MD���"O&)0�5 f!⤣�0L�Mj�"O���4�� ��0h���J6����"O4����ΦJa����[=)>��"O���A�ݜh��$�#�ۛ/	H-�S"O�yS�
Bn~<5����sd��d"Ox���
M����t�IM6���"O��Iec[��\���IK>����"O��`R�G�<��L�G��;���a"Of�×�P2-p]��H@{{�m�'"O��0�-ޝtЄ�ѡ��_hƐ
�"O���J�+�r�bN���)J�"O(�ÏS�^|���&�e���q"ONYЁ��h���֎��
J��"Op�K��F=cpL�Tl�h]R� �"OȘb��{5,1�M͍/3���'IN��s�N2lP����M�:��#	�'��h5��9H��y��<W�Pa�'_��9�/�0�t��<��
�'����"Ӗa�,hK��[�C>:�3
�'�(�#D+Y�]���0>� x!
�'��8�"�<i4&��I�i#�@	�']d�P@E�m(����R�L��'�j��QC��w����A�*M��S�'+"��p�-E%��+Q�U�5�:��'g��a7F��g8Erqك:T�%�'`��jw�
#P�&๠��.k�'�0�H��	�*�n��#�VeY�'�JYZ�F�tX�H
����t �'y~l{�'�39;�a��P�V\r��	�'�� ��*~���*THĄl^��'\n$r0kĩ\����X,"H`�'���3����N1M�*x��7D��;Ƌƙ�zIj��Ǩ#M�ݳ#�6D�\04(�8��-�A���<���t�9D�Сg�meX9�Jc��,�ӭ��y ��cb
�#K�<��� P$�y�K����"��EJԙ�r�Ҷ�y�b@�[�v� �I@�B8 �����y�GΫ\���"F�H Ȭs�I��y"iX�b��d�����>���.ʛ�yR"ԝe��	���E�����C��y
� ������d�p�'��1R��x�"Of���+�A3PY A퓭_��7"O,���	E�j�$H�E%�5/.5��"O��d��q���Pd��#E aP"Oj���Ӏ. �4�w�7'��a�"OJ}��BM��p����P�_�q��"O��T-�EY ��<z�<�U"O 3�c� ^|�Agk&KΪL�"O����@+2\IF�@�k��u:�"O�%�w'
:����2
v��l{�"O�-��Y0�S�Jh�`"O����GT"^�P�2Í�3A����b"O��{�g��:�&�y��ʦ����*O�y��JG���b/G'H�Q�'�ܠ6g�F�b��%X1Z���'g^�
K.'�*�`ܘ=���K�'�f�bI|�<���Թk� !�'������s��İ�E�^gB�*
�'����f�d�"0amY����	�'�bպ�KU��B�X2���V�Fl�
�'�jx�  ���   �  C  �  �  �*  w6  *B  �M  iY  e  q  K|  3�  �  �  �  �  ]�  ��  �  ]�  ��  ��  ��  �  O�  ��  V�  ��  J�  � � , � h �! '( ;2 	9 L? [G �M wT �Z �` �c  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+q��62\���<4�d5h��'�B�'���'	�'/�'�B�'��x�.Z ?܎Yf��0d�tx��'��'���'�"�'��'���'�nY�5��B��0��g��ծ�pW�'l��'C�'���'���'���'b��i���8��}��dK�� �C�'1��'W��'�B�'���'���'?�%�����غs�9
lk��'A��'l��'B�'��' "�'O���ek�92�lu���D�+��'�"�'\�'���'��'B�'�n$Q&菷U�~�
�"��]x#�'���'��'u��'�r�'���'� �H�N$!��y;�Ã+K�f�0�'���'$��'dR�'���'���'�Fx-Q@�蒠�6/X��o
�?���?i��?Y���?Y��?���?�Po�^}��� �	\V�p�'F��?��?���?Q���?���?!���?auj+2��!� :D�|Hʗ��!�?	���?���?y��?���?���?y��ь�����/�&8CTtꖢH��?����?Y��?����6��O����O��DB(Hc���$��[��$�E/U��b���O����OX���Ov���O�!lZڟ��	�P��H���L�!�"��~�-O���<�|�'��7m�?3�p�)2N�&g]��*ϓ�Zφu����,�ݴ�����'�"nlr�q%�E)-`�����:�r�'hr��iw���|bA�O��)�t u=#�h���	W4+���<�����4ڧk���j���=3�6[��
b�,Z'�ie�,��yb�i�ڦ�ݛ,���d�!&�;$,A�;�R��	ΟDΓ���	�^46m`�t�E`�p��%]���2��t�P�p 2Mm�����'.�8bG�C�8 z��;1I�(R�'E�O�I�M;�˛C�Fmv��'֏el�C��:6\ui����>����?�'<�ɯF�*Iɇ��<Yެ��Zn��?���><�ޠ�|��+�Oܠ��l��|���B�`([ LK�2O�0�.O��?E��'Lt��ӯT�L����L�6LI��y,|��,𘟌�ݴ������V,ws��c!�ΗM�k��� �y2�'�r�'o��b�iD���|2'�O��!���N����!�6)����Gb��My�O��'.B�'���_�v� 1��k�/2��GM!n��I��M��aɐ�?���?�M~�<�t�*phR/�J���ӋU�>\�`_�x��4��6J9��	?K��S�%��"�L�;��C$$fx� ��= ��:'h0DrA"ŕ���<��*�I�rd�,�d�>F#�����fM�Iן��	����i>U�'�v6ّ��$��c�b����ѳp��h��Ъ%����Z̦)�?ѕS�T�޴c����n��b�bR?#�V@Zc��&r�^x�f(�6)h�7m+?Q�)��
���)���s�=�f"�|�Pn��hR�鷢�K��ן���ʟ��I����|����B】2`�M��O+ �&�3���?y�Z�F���~%���MsI>��_#L�x��Lՙn~=j6b6
��'K�6��ɦ�/a���mZs~�!P�FO����	$����A��TǄ�U%�ݟ�@Y��4��4� ���O��R�'X`��Y��X��C,�M>��$�O˓�����,*2�'��P>5�n�|Ot$�rd(y�8����9?1sU�`�I̦]�O>�O��ucr��X��3b��)G�D���&u�@(��P;�����{S��Oα�+O�T�4�Q� ������W�K�~���O>�D�O���	�<�T�i%��d�Q^S�D�"B�^H����M��'D26-+�Ɋ���g��,aG�֏%dݫ��ɮ|	�{�FҦ���4xɰh�ٴ��dhVѓ����S�?P���e
�g�Q;3��p����۴���O�D�O����O���|R�ݻsA�\S�@BE%�kB
�vK<k���ʟ $?��ɓ�MϻD��tH��(I'����S�f�I��'����$���tET?ԛ�=O*D`��͖7NF�k�>���S5O�h��$:�?1ᣩ<A��i��i>9��>G���JeF�}꘡R0�S������,����'��7�í3�`���Ot�DS�7���v�6 �Ed��?2~$����Ol�n��Ms$�x�/&|��Y�
�r��H�:���'{����FQZ
�O�T��#3��dQ0�?��G�	�dTc���*d����'�̫�?����?)��?Ɏ���O�mY�ڥ�p�z"����8��Ԍ�O�Mo�p�p��矠��4���y���c���׉wTP�[3���y�EoӘ�n��M��f ��Mk�O��³Fş�s��.�R���Z�y:�$�N�,˓O�f]��S͟�������|��#� ~l,���Բ#Z����Eyrco�N0�&$�O$��O���d�?!>��'G!�Uh$!J(��'� 7�Y릭�L<�|��F��'�2YC�%ۆ�"��͚���ȁh_~�׼5=��I&>I�I9�M�)O���,M00Ҝ3���#MdT	b�O��D�O��$�O�ɪ<���i�j	q�'wZŲ�$�W�n�jqh�,�rl�`�'7�6�3�	����D��͹ٴ<����7���8��G�Z�XT�"�z�. ��i��\�Xp`OD�n �iq�)�D�~�� ��c��PZ9V|��*A9bT�0�0?O
���Oh�d�O��D�O.���Y�� K`��b�X]� �C��Z�Vr��$�O����}	�ln>��������Wy¬L�zr��TOاW��Yd�\>��6m�<iC�i��7=���A�q�
�de��KG�P�A�p�R�ߌ/�h�1 gؑe� %
�+���?���s����uڟ>���O��8B��� ���3v�se�\(6v��d�O�˓&%Z����d�Oxm��?=i��Z��]Nm@�d�$	o���OH*�t�X����ūݴ��O�̄1��!G��BJ�_xP"�̝C}Du��A���D�ٺ/�6�T��?��Ӽ˕�S�\BI���e8X��Ȕ��?a��?I���?ͧ�?�����Pצc�j�����*�B2TV��d�6������ܟ<����]�<z�4%�@-�"�7B5z�C�L�7)��!R��i�P6MA�$7�.?Q���7S6v�i2���N>�HD���j�2�A��յl��6�<���?���?A��?!*��e�(/
����
~�4���[Ǧ��!��JL^Y�	Ɵ���/���i>i�i�%��([;ь����%"�Z��@U��MU�i�z7��<�|���1�M�'_"�"�oQ�k`x�IV��e���<��h�5!���_��������4�'�T��d��?�%��!#�D ���'�r�'rY�X�ش/��Q��?��N.\:�cڎx�a�%�,c��	�OL��?a.O��lZ�Mŵi��	�@��h�e�)5A�KuL��V�>?�抩�9���	W~�jmݕx��'U�4�I�x�P�`&S*�l�CQiշ#;�����P�	񟈗��)�O���O0TҴ�����c͌R��%AQ�O �l?Q8|��	����	ş�����w�~�Ɇ�oj6e� �ԒR�:���'�j6M��3ݴN�ߴ��D��.�@yJ��6x�d��e�V,��f� i4���E�O:�ĄҦ����t�'��'��'R ��*k{�U:��""�����V�Y�4!�(��(Ȼ�?Y����"��.��E?<^jla�*�J��<2ѩA�y}���'ɾ6M��	X�43��>Qr��P`�Ւ���fR~���,r�H�(?I2�K"Z��������'�8Ȋb��gh}Ү�5�*Hڥ�'���'������_���4|t��*�dZf�
1M��i�h-�v����x]H�/ۛ��$�ty"�'��fk�J!���	"��=S�#G�uw���K(m��7*?�"D\�C���+�$ehݙ��2ar�}pc��>%XȘw�Yj�D�ǟ���ڟ����Ii�'�\��(��|�T.@�7�҄p���?q��R����_��D�'JB7�5��ݽ\�����a��`����Qמ0��'�<��4h��O�.�
2�i�d�5��KeoǉBe�l�F�I�.�rŐ�I-N��TK�h�
�'�\��'��'c�'gd1R��6C���%��Iה��@�'��_��s�4.z-��?Y����)]9��	��+���"jIo�������O�7�Q_�|�Ƭ5Vh]q&:ȼ,���9n�U�ЀV�'r����d��`�U�|�
C� V����O��ج�vb�1�I͟��	៴�)�iy2�k�� ;���P, hq��ԦO����LK��I��M���j�>)ƷiR��1#��#"i*��U�L����!/|�R�mZ4-�n�L~��̶"D(<��n�)P6Z��Q��W�c�Dڴ%X�J*��<���?!���?����?!/����F�`��� A�Yl�.GB�7��x��D�O~��/�9O��nz���`S:L�3�!�#Po��P���MK±i�NO1�d9B��t���ɢ!,�z4(��ZJ*XӲ�����ɩG�@]�%�'�x%�L����'w�x�t��x?>��w��$h��!�f�'=��'�Y�X�4q�����?���Y��r��œ9XVM�RÌ�a�������<Q��?�I<q���)�2���E��ZuiANA~��J�咑��W��OP���	�W��L��x#�RQ�H5�.���#C�^��'���'����QEP�^���!ݥ;�b�! ܟ�ڴh�
��,O(oZL�Ӽ����_�H��ȌK:)�7��<�׾i����`���Ѧ@~� �H�(hWn�2��`DE��I�E(��i�x��d*������ON���O����O��D��/�� �Ac�$��I����wJ6ʓG�&N�"��ԟ�&?a�	�x�~��Q�O'�:��0c߻G���ʯO")m�*�?aL<�|j�l�6���� ��^�N���,<i SȈ����Z�� ���)�<�OʓV����9d����R�F�n���(��?I���?���|�+O�DovCF��	u�Q������$jɜp��	,�Mۉ��<����?��44� ���E[3v�X�;���&���M�M;�O�8"��?�r֌4���� �[���<!)����G]�p� ��s?OL���O��$�Ob���O��?{�HZ�Q,�C� H�H�&/�py�'��7M
�5���M�M>9⁓�
���C�y�RG�#�'g 6�Vܟ��S�H�R7M#?	⁍E�b��p�S�my>��
�`k�d����OՑL>�,O&�D�O����Op1�d�V�ߐ�S�!h��{w��O\�$�<1��ib� ���'o��'s�S�/7DX #��#����]�hF�$�I&�M���' �����O��``��<�F���ȓt��	e(	
���Sb��m��	�?�3�'��a&�pr§��u�x���D�\�|(#�#�����ğ4���b>!�'�6�Š����a��B�@��#��Ox��̦��?��S� �ٴv;���S��*,�C�ľcȬғ�iM2�E�(��5O���O�A}�t ����)� �p��ǳ?�����ϖE�79O|ʓ�?1���?����?����)G�|��S�XL"��R7v1
tl��?b�t�I˟��L�'|՛�we�P�� [l_v�I��B�0��RR�o�ioԟ<���OAli�p�i��D��f ���'����U��y��ě�z{�e���{�O���|���!�y�E(Ѻ^т�)�M�P$�İ��?����?1/O�oX"ެ�I����	��vT �F13k��*<p���?��^��	�4Rg���'��43�hLQ��//1�\H�E�!�\^N��M�Q2p��|����OB����+ E�C��w�֑�w�
P�����?��?���h����س7��8�.�G��H�2/�����¦Ey�Ĉ��d����M���w��9;��F�$ᢱ����,����'l6-��M�I+�t�mZK~b�H�,����ӵC���e!F7�ҹAĊ/4�'�|�Z��Sן ����D�	֟ �4��?@�ʅГ�N/}�l��[_y��g�Jmj� �O����O\����$ҋ�,٠�@�*o6�[U���s2���'�T7m�����ɿ�H��Mj�햣0 �C�O�TW�C�C�u+r8£��$+B��?�F�c�Oyb���v@�c ��,���AI�1	3r�'���'��Oe��MC����<�׾A�RUB���}�������y�,t�@㟀J�O�oڋ�M�Ǿi�d�'\�İzׇ����c�ƖZ��&���[ª�5Q������f�p�f�:��1�Um�#$�f?O����O���O����Oz�?�h�!V)=�P�g�B�(F�����$��6�MÕ�z~�feӸ�O:5S4��N|pU���ڒO�@qw�s≕�M����&��(�&��hj�MR">Z��s%�(�\�2p�_ 6���(b�'X�m$�Д��4�'��'���Gg��K��@�%`�mTh��v�'a_���۴S����'2U>�He݆	[@�)WU�P�H��!�8?	�^�4��4*��A"�?�s�A0|���QW�2{،ht��09�,8��>u���|"a��O�1JN>Q�	���	7�X�iv�B��ܼ�?Y��?���?�|/O�(n�0Y� ��R��V��(�I��	��y��-���<�I��M�����>��i[�E0��'_��9�h[�/�M`���O7���06-5?�rȂ�z��I݀��3@9>qRbH�,��H)���2n��<��?����?���?�*�"]��	~�!��_t���������� ��Ο0�Iԟ@&?=�I��M�;:� B��?g\1Be��W���MC0�'���O�И���i$�D�Vq��K���3R("�7�ǐ/o��0��([�v��O�ʓ�?���~�ViA�^Na�"���<E�Qy���?q���?I*O�qm�4�2��	ҟ�	y�.���G	,`;�H�+L�<�?	�S�(��4hR�x�Q
'J$�����҈�3e�<���JA�у��ؐ~8ғ�����y8@�$Ƙ`�ʍH���ud��E!8
���O��$�O��D �'�?���)��rgĔ y~��HF���?A�i�LX`_�|�޴���yW��0'VF����
�fV1=OR��; ����O�6��H��7�<?9�fG�1JL���uf`h叞�EO\���H+�,EM>�,OD���Op���O�$�OW�:К�b��Htl⨚ŤJ9������jd�����ߟ(&?���0rh�
��ݠ�&T �m�0C��b�O��lZ�?�H<�|z2��G��\�0��*8�����'w6U��H���$�3~��ȡ��'=<�O��x�D��� v��|�Ы?n��H����?a���?���|�(O�~(@��F�'$r��V���kfᐟx?�u�'�p7�7�� ���F�}���M�!B�sG�]���F���R ӭ �bŉ۴��J��H�h�'o�v��|��N�~x�h�FO47�6̻FFW/L�D�OD���O���OD��)�S,�I���#�l��TfL�����џ�����M�fS�D�i��O%1F�<A�\���"_�C� �R��/�M�����D���}ћV��0J҅�x��i#��ʠstQ10Έ�K�����'c�&�������'b�'a�8J���.���㐻kpsv,Tk�$�fT�\9�4��@1�OG�'c���wt=Ӧ��9$՚�{堚�v&���'krW�؀ܴ)��]�l�O$��˒�OH����.�)+��ذ��/�,��4�Z�iq���GZ���S�i�b�_{�ɂ0�By ɟ�|��I0$��.Y?���	ԟd��ݟ��)�Nyr�d�D���K�yD }�^-������bΰ�H��6��_my��i�n���啂#���'�ȂF�Ĺ�Hf�Ȱnڕ~Z��m��<��,��!����>4�-OpM{w՜A%�1`A�٠�e��>OX��?����?���?������Z�4�Ha!��);0�d@S���um� ]�-�	D���?9�O	���yW�74�bܓ|�f� �G�`��7�矀�'~�O,���OjPz��ik�dʢ��1�#�ܿK�� $Ɔi���Eb����Hr�O���?��^Ą��rf�Y���1�O�S�p�b��?��?�/O��lڊLGp0������I/��BU�SW���h��ًa?V�?�\�DaݴJ��x�hI)zB|ɲ$D>;o���č��yR�'r!�#..`@�\1\����S�2�T�l���]�r�������a�^�i%Tܟ��	�����՟(D���'��x�Ó 5# �A�8/JA���'�7��r�J�l�f�4��4a�BX=E`D���X�0����O*6MO����ش,Op�4�y�'�4D d�?�Q	� t5�A�9)bR�;p��`>���<����?9���?!���?�SɅ�Ls$4:ъˡCC
��G����dC�����ߟ���䟄$?�I$4hp	p⨗�e2�#�n�#w?���O�`lZ��?iO<�'���'N�Ct�S���!v-���[7禈r/O�dX��U>�?9"�4�D�<Y�Y�(�@i eꝔF��}�!߲�?Y��?����?�'���T���: F�㟼QP*��%��HA���Q�r�۟�ڴ��'���}�����O6M��w�X�(�,_<u>X�CM�R:Ќ��mv���	՟0CE,��Yly�Om��;)�D�	�9H�A���y��'9r�'���'>B��1]n�����0�R���jXd/p��?�Ķi�Dq�O�" i�*�O�����`ܴ�æ������!x�I��M˒�i��4��Rz�f<O$��ظS��)�DZ�5�uh&�X>$}�d2s��?��@4�d�<���?)��?�v� �X����U�ߦx� rH�?�������(T���ϟ�Oo�䣁Ş��V ��΃�P<��O��''T6�QߦA�O<�On�����0���1��w.n���(� x�&��4�` �?,|�O�ɗC\0+��왶�;�N�� e�O��d�O���O1�xʓ]?��Х����2�'W�^p�F�(ܜiP�X�P:ٴ��'�^�N̛��mZ`8� �@6ȝ�U�ףI��7��˦qz���}�'^:Ga��?����d�s�J3�:��׭��zR�8O���?I��?���?�������~�Z ��%q�iB �V�lںs��y���`�Ie�S��I���k5�h��P�7�1R澡Y����&R��s��%�b>���D¦��9+�+��I� �B7MwK�,�@�%�P��O��yO>�(O���O8}p�jD�_�z�`KȔR\���(�Ol��O��D�<QP�ih�`�EU����+�
u��_�_��Q ��I.`<��?��\�t�ڴ"����8��0�D�±ŏ�Z𶕨�FF'���'.���wl��,D�b>��'N���	�$)j��צt|�e�(ɲ&������������z�O�R!I�.&�xZ�(E�r�z���׶(�!f�>ĀD��O��DOЦi�?�;FBIb��6!�x;d�@�����Oj7m�)n�R6'?	T�^�	�����HVX���հb��ÔC0&���N>�,O����O$�d�O����Ot8�7*�x˒�	��|r�ϭ<y��i`�Ԃ�U�\��V�S۟Ƞ`ɐ82n�B�zn���IK��d Ӧي����|�����P	_�Y����2�"u
�d�7 ���N���Г}_�p�c<>�O��L����3��ʇa0�������?����?���|�.O
qm�)N�vp�ɝc�rQ:��܊F���DHDʨ��	��M���<����?!�4+�J�jA�����p��� V121cǫ�*�M˞'
�)FfH����9l��?I��W,\��iG)~���T�Q�>��şl�	��<��˟���|�'Q'��H�ܩN�.pУ�O�O��D3���?���">�6��:����'��7�(��[�"b��zc��28@�AvN1,��$���4zƛ��O��ca�i���O��%&
a�j�k�䙫x|�r�ǆ�C��H���N�O�ʓ�?��?��G�VM񑊘=�T�+���!�~����?q)O�oQ2���˟8��P�Da��K�h�GGP�r�P�X��F���d�b}�f�����Q�)���K�@쪙�������n/X��$>���+O�ɇ��?Ao&���T�X��'�3��$��&ԌFz�d�OX�$�O��<�$�i��!B��Z_<8�@�h�'gS�T�r�'%07m(����DB�Eې`�,]�IK��^�T8��\��Mۅ�iB� �v�i���/\��-S��O2�)�Δ��
L�7%�ش�΃}��mϓ��D�O����O��d�O\�ĸ|Z凁�Y��#qŅ�?��A:�d�K:���|&��'7��O��ޟ��i�qYCJN9:xx�Z�3YF��?�۴�?a�O�O�4����i~�J�U=���Fj�� ��l	����Ro�\����t�O���|���C������ :`n��,�r>�#��?���?9(O\�m�0j
�	����Ɍ\�7+�X�+����І�N��$
���M �iG0O&�����?>��tj%�;��xC7O���I�lP:���H�0����?�r��'o�I�I�cJ�EQ��(89�����*$�����ܟ�I�4��k�O��l��@�㎨{l����R7l��l��xA�O��D�ʦ��?�;��U0��_>a� ��� �:����?!ߴM	�v

������xJ������+v�٩�&R<$�Rɔ9D=<Y$�(����'���'��'���`
�k���Ń] L�|a�[�\1�4h��x��?Y�����<�(�>����N�/y$P�dI�V��	��M���i��O1�����AI���{F/��x!S@�4`BU����"� �/n")BP��|yҋΧ8����@��� � �D�
0�R�'�r�' �O��Ɏ�M��![�?��牦6"G��+=�:�l���?���i��O8�'�D7�P�U��4߬���_�&�`T��GW\��qZ��MK�'���J�?1�E�S���d��Z���4�``��C�<`&�4
$ӻ{�$�O����Of��V���'���\������@�p�Bod�I`�������M���A~� k�T�Ol)�Q
���(�H�EG�p0`��R�	0�M�ױ��tΉ~ɛv���R҆4� zXb� �zy��:����5�\@�d��%�?ٗ'9��<�'�?���?Qwj	��aPa��(p5X)`��%�?�������)�%��̟������OMJ��]��u�Q�j)�UJ�Odp�'��7����l&��'j��qA2��2y܈Y��	z|�ē�"[&��J���4��t)�"픓O��@��a�H������x�%����O����O ���O1�8ʓ|z�&-�-�, Jĝ�88F@�יyB<D���'A�ee�&���ODtl�%s���7�9�h`��*�{gh�+��M��Ύ�M��O���K���ɩ<)���-tN,��5��w�}ps	��<a/Of���O|���OJ�$�O��'#��iP���,Kv�p3oMI��ѓ�if�ђ%�'m��'D��yҏ|��Ζ� 2l+	^�iP����C�4,umZ�?�O<�|R�):�MK�'Z�m�¯��FF���G!��O `��'�
�k�%Y۟�K`�|�U���ܟ�D٪q��r�� ���*�g����쟤��hy��t��X���OH�d�O�)v��
-��=:�M�?�m��&;�����Ė˦�Y����O���ԅV["@�&��<Ge&H�'�D@&�B�m:��g���g�՟L���'��ӆ�W@ubus�׵h���Bg�'���'Mb�'��>��e��D��a�)�"�C:=�m�	��MSf�2������?ͻ�˥@�*�8u���)C�ځϓ|	�FA�O�7
K�\7M(?���)L���i:���@�h
�?W6�r6ǆ Kk��K>Q.O����O����ON���O�T�@<��,h��=|��q��f�<9�iDƅ�D�'@��'p�OAR̲Ek��԰1�Ĉ�'�'4z��?��6��O(O1��A�S" �VKf ��!�a��d�aH�,bn��n�<���!$���U8����DC%G�����K�8��#�P�)N����O��D�Ol�4������)��'�/�%&<i�쵢���T�	�0
����@}BgyӒ\����1�ZB
�h��<(�~p��JǄP��o~�E��`��+�O�W ��YX�#�/[P���R��ɿ�y��'���'�r�'���F7x=S���:�)���>T�˓�?��i!~���O���k�p�O�)�!B��>��I�ꂆ�H:`$\B��ǟ ��ffKo��s
�� ��A<Z�� 3Hy��ҥ��
M�6�$ל����D�O��$�O���H0Q  �2���OeTHB �L�T����O��,��V�ڎ R�Iȟ��O�|2�Fތ[Ќ�zB�^)Q���1�O~9�'ո7���'��'u�;Ƈ��c�r�@�УL��%c�0<V�|��#��4��@���\��O�8���I�8"I����q� ����O��d�O���O1�f�&
�V��&{���p��
�-$�����$	���'ODy��㟼�O�En��d�4�cC6j�n�jV��f�@Q���M{#G� �M��O1�Ș��
B�<Q��>d<B�;s�5����<Y.O
��OD��O����Oʧpf�q�d�ƷcՂ�[�D�/myN��&�i����F�'n�'��OlR+n��ΌG�"��SW
c�t�ԋF9�mZ��M���x��$B֬G���4Op��Kވ_�|	h6שy�Pa�d=O� ��T �?�w+5��<�'�?1�e��3O :���*~>��
�
=�?Y���?�������¦}�5E�����IџHj�'�#I�Ґ`uIՃ�.��d��e�
��I䟼nځ�� �~�d��6����K,p@��'i 8���]A\6����d��Ο���'bR&a�5�*-�w�N�>�P0a��':��'���'-�>��k5ʔ���YO���Ȕ� 4����$�M�Sm���?���ޛ��4���`-���Ց�,�:4���4Or�nZ�M˄�i�ؑ�!�i|�	't��-���O��y�/�s@$Y)	˼X�q�q�\�	|y�O�'���'_��)0�B�H0HB�њ�˔*5���/�MK�,���?I���?AL~��b�i��� !,�"���i�xy�[���428��� �4�|����\�f��?K^n��k�$�$�jiq6T��D��\�e��/�b��m�Zy2-S���IX0/F�3�d�	sj:���'���'��O��	<�MK@%Ή�?ae�4j#(�� [l}�vj�<���i��O���' �6�To��yXB,�k�1]���f		b����	����'"�i�F���?�Zf����w?�`�ή�R�S`M�$޵�'��'�r�'jR�'����*�G�A���;��Q�dV������O�d�Ov�n�6u�p�O���'��I�u�Zh	�|�����J��~�BO<!@�i,V6��^e0�y�R�I���Z��+~&��Q�*����F!H�YJ4�b��'�~�'�Ȗ'���'���'9����Ö8Xn&���4��:��''�S�̨ٴ~�D����?Y����3l�^��<2���X�JW�� �����Uj�����|���<�h\`T!�X22��>~�X��I�;q;������sy�O�ȵ�	���''�qs��F�PJ��4���p��'�2�'�b���O����M3�LM�0v�ms�A�*J`�)r�C:K��1++O`m�S��/J����M����j�A���/Z��TA�I�b��6.c�J����n���I��L���N���
pybg֥"L�k���^u���q��ybR����۟���ϟ��I۟��O�1����x(����H���4Ix���� �O<�d�OT��:������9Eq`��#DI�)��L�׉P�d�T�������|J�'��֬�+�M㘧� ��	t�E$��h���$*zHY�;OPDG��?��=�$�<a���?�ǔ�&��A�H�.����.O�?����?y���dH��%h��W۟���������P+U���k����� Ȗ�Z��7��I�Mk�iP�V�9�mľi@<�%���P�J���m����^D���A�� ����C�O�;�XF\̡��J1 1Ȩ�6�F`�[���?����?����h�n�DU�\D5s�d-@v@\+�F���䦑s�3?)ֶii�O�.<���3b�P:Kj���ЯJ�W��$B���Sߴu,��'_�gT�61O��$�!��`8���,�G�H2�u!QK4�~����2���<�'�?����?1��?��S�k+���r$�*��cw���D���[�}������|%?�+a�����d�78�ti���^�'S.O��v��($��i����I�A�6��fg���c��O��A�/� l��	?U��9��'��u$�0�'%�ૄ+ٴģ��e�����'���'B���X�� �46�Q���T����"�'T�b�Ұh�/`�TA�$��$K}�%q� }��Ħ�;�"�J��9BUQr�ɴ�S����n�^~&�N�D���.h1�G��.��E�Q�M=�|�h�A�yb�'�B�'&"�'�2�	@-Z����%Ѻ�K�o�?1n���O������$�m>��&�MK>����κ�Ҍ�
�{��O��xx%����4���m|��ڴ��:��`kө<���aa.�� �։���:�?�c2�D�<����?���?���I6r}J'�ԳL�8�H߁�?�����d�-�Ӈ՟x�	˟4�O?
���끰����`M��O��':7���4$��'l��M�g/X9���j��Sr�
i��I�*Jv`�կO���4��<��9X�Op�J��H8d!��rO��G��O���OL��O1� ���*H._B ���l�%�>��h��U���T�h��4��'�>��CX1�H�ڦ-���5�ԍ�6�i�L7M�p7M$?�g�2٨��#��D�=�p�8U���M�`$#��y�Z����˟���ퟔ���H�O�L��g*\�;�*�c㠍0����N|�<�eg�O���O����d�ݦ�]�f��q�ȇ:
J
5���\�@|�شJ�&�"���R��7�b��8��Br0�$��y"��Q(j�t(�C� I��`�Vy�O:� �"��q`ę�`��,�\1�'���'}�Z���ܴp�������?���N�Y�ꌻ;z�p���N�66&�q�"��>YӺi7�6-�j≹{�X��7�җS|���1�� $������9u.^�"~А
�B+?��$F������?����,�R�01��q��I<�?����?	��?Ɉ�)�O�u�b��	ʦp��>\�L:7`�O�mڒ~�x���ٟP��4���~�g��<�d��p4^��#���<Y�i��6��O�dKw-`Ӭ�u4r��i�����jʑI�P�
��g��TP��^9����4�h�D�O��d�O���=Ub\�"�d��R"�{W�8%'˓�����j��'%R���'��=�3
�.C^�B�Q	Z.h���O�>鲺iD��6��	ɡN�mr��ˊ*��СÚ�k�D��!�&M�,�h�N`�pA�O	�J>�(O�L��m�J�����	i@50�A�<���?���|j(O��m��6v6@���v��&���)�N�
@�)M��� �M���F�>�6�i"��e�ƀK���'�4�0��p\P���
�Ga�7�&?aE��=��)'�䧰����N�*i�s��:O��K�#��<����?)��?A���󉚢-��Q��"[�����Caڠ�D�O��YȦ5�!o{>��Ƀ�MN>�&N�:U
��s�B�h>�!��ڵlb�'�x6m��)�<eL7�!?�&_�U6����;󔴣Zat�0Ζ (���O�	@y��'LB�'�ꏶ
m��sG��l�.�{�M>�R�'b�	-�M��A����O˧#��%�5���7
�,AE��8�O%mڷ�?O<�OD�Qh�$G�.8|�D*~�1j��Fi�����i>��6�'_|%�L��O�xĞ����C�M���p��ҟL�	ȟ��I��b>��'o�6-V�6z���k��g6 �q�<C������O����̦��?Y�S��Xߴ�ؐeM(�.U2��S<=Ƭ���'S��J�{4�6��ؙ2.TG��$)Ly�B ?Q�0)%N>BަA�f��y"U�|�	ӟ���ܟ�����ȕO���!�M�(����x�D��w���˷��O���OT�����PԦ睊k�(�[��K�{�0Y2���GU�(��4K��֩>��i+3�27-�|�u�-r(�����U�%�P�K1ni��"7+�	KB�{�	Iy�O�"�;T�6�X��`f|e����/��'�b�'��ɹ�M��E��?���?�GJ^�q^ ��ԫ,�d��A����'W��a�fgjӢ&�C��Q�df�*�(*�e�A�6?9U
(n*dk���G�'c)j����?�r�T���!�l��h����3�Q;�?1���?a���?!����Onu�V��-I��R+ �vIΙI@��O��o��h	�'�*7;�iޡ���V$��Pp��?>��Cp� b�4}��o�Ȫ�g�Z�"}}h��柪RV��k��q�`��ш��`��h9��<ͧ�?!���?)��?i���5H�T[�.��f�4�������ha��ߟD�	؟�'?�� v�R���
,\bIM�5�ΰ!�O`�lڅ�M���x��T��� 
���R�vV�	��1�@�f��u!�I?�b��d�'�BP&���'���Fl��.]p��τ7� tQ�'�2�'�����4^��۴K�-��m�D	�OJ%�Ԣ���!k��̓����DJ|}Bs�Ʃmڴ�M3������j2Î4��¡e��J<�t�ߴ����x>������OB��]�2��JI�70Z ���$�y�'�r�'C��'+b����
�p��'K�'eF�"B n�@�d�O����ۦ�P�Iyb�p�>�O�Pc�Ɨ�D��Bd[9`,Y���u�ɞ�M����2�K�-�Ms�O�P㲦G1n�L`� 9#6�*�^"iNS��RQ��OF��?���?y��Z]$�4�P�"�l�Hg�S%0bh���?�*O`�mZ%�'��P>y�m�yb6�C&"xBx�3?�G\��c�4��xʟ�5�� O�֌��L/����� $�x�M֨b`P��|j�"�O��	K>)ԋ��H��D24���9��C7�?A���?���?�|:(Or�oy�y���8p'� �H�vK�QS'	�柀�	9�Mˍ���>��i��lWF�����@!�4Bv`lӠ�o��]��Lo��<��1����� �X*Oh�1�HX�gŒ����*��<O�˓�?9��?i���?�����1b�9�E��� �5�S/1�@n�=K'j��	⟨��g�s�8c�����$�?u���MB; �t��s��L��!�O�O�����A�>�P7Ma����g�$F���m���gp�8J2nD�Lf��r�ILy��'�"�Ε��5�e� �9�t9�߮I�r�'R�'U�ɾ�M�񡌜�?���?��_&���;f,��S���'E,�v��v��O"O~�(�V�x�D-�� ՈR̂ةE<O��$� dtx2���Pn�˓�j�!�Oj���fH��P�ݶ"�v�����T~Q���?����?����'�?����?�)�(�����b�8!��D�vmQ�?!��iږ��'���'l�]�l�i�咅�Y4z@T,�!�X�=��$���I��M[g�i򩎹d�F��؃��%���$z��#U�G�6�Zae��\�ZD&�h����'���'�Z֛&�D="I��q���+"%Ѣ}S���Mv��?���?	I~Γe���
А5�T� %A@t��#E^�L�Iğ�%���"�zR��z2�H
l��C��A5	S �;Ю> �ʓ�4Mِ�O�d+J>�(Ox�0��	+J�Y2�D�:?�<qr��Op���O ���O�I�<��i�^�1��'Z�$h�ib)c��Ǻ�#�
�=���Ʀ��?�4Q��i�4:�B�i�T�ʇ�@�8��8�l�-.z�i��6s�������������/g�S��Փdlׅ*G����$C�0���P�x�X������	ߟ�	՟��F��<D�X,��^�':-3éΑ�?Q���?�3�i��1r]�dKݴ��I�8�+H��4�[�(X�%)����x�"q�V���D��czӄ�K�(���,��9s��`��}������4�|�D
������Or�d�OR��	�\hP*�^�j`(8��ƭt����O����E�.s��';�S>uS����/:�j-"�Ȇ�:s�I%��������S��lA�z��a��?	��9D�A�0�V �
R?2����u^���J���k�	�,{&RD
R�pbe�t(�+)���I��I۟`�)��Wy¤c� �32	��bG���������$;�����O�!oZ]�W��	��M�K�q6!R�V�gϦ�ڶl��2�i��h`ֲi�I�9����O�xM�'Z���h� /ТeI�dZ���Z�'��	ӟ���ڟ\�I��H��s�����ݞ)�F�+���U�^�avNq�H�R"5O��$�O��������<�jI3�P*�� ����-|](A��4ye�&*&����<o��6�g�X2sg����bfhK�Q8�zF%q��� ��f�r��j�I`y�O���&(=b�/�ɚ!C0C*J�b�'�r�'w�
�M�W���<����?�K�<�Y�C��'��Kd�����'��L��dӊ�'�$��G�|�[u�B'\r��`${�H���U,ĲD�X�	I����t��O��A�s��E&4f���8���^<H���?���?���h����%wfha�j�+n�!!`B[������Ǧ#��`�ɯ�M{��w����U��
DZ싓*��P�Db�'5l7��˦Y�ڴ�:-�۴�yB�'���x���?��e��5�\H��Y�2W�`�w#�9r��'S�i>=��˟��Iʟ4�	;I��� ��|��/��!�ݗ'
�6�90�l�d�O���'�I�O�ܣw�(E�����ފO�4��vE�}2�m�j��Ik�i>��S�?Q# E��Aqa��^�tX�@W"m���h�iFy!J<]��}���Q�'��g���ihګ>�vU��ڀ0��	П��	ߟx�i>y�'@f7MF�?ST��]��\����M�e:i��LYD��Dʦ��?)R����4u�ijX��׃H�<6�2�nƔq�.(�"��8]ڛ6��8���
U��T&�_����SEM�
���k�f���W�c���I����I矘�	ß��r/��qs������L�P�Ӏ�V�?!��?��i� ���O���h�J�Ov���o��* ���n�q�e�X�ɋ�M�w��jVN���M��Oz�1���"v$��bF�5��D�,M�~�(���"f��O ��?Y��?��1g��)���R�H��55B(����?�-O�lڭ?a����@��X����k�2l;��M�\I�k��U���d�Y}�Ju�8���F�)� *�Ӆ��b����9j�H|;h=%h,ى6[�w�|��|b��O��O>���Nv��3c�ԣ-�%�'CP��?	��?��?�|�+O��m�(4��o̶|S@�I�(Z�r!I�h�џh�Ƀ�MC�&�>AѴi�0���üvŰU{��V�[=� �d��O86-	���6�#?9�a@�mކ�)׭��d��w�>�Ard
r���q�Q�J��<9���?����?a��?.�
�s��0J�:s��$��Zs(Gߦ�z�A�矰���� $?�����M�;iD
e��T�+d�P�7�H�n���c�i"�7�Y�)� "L��l�<�� ��p���f�g�����N�<A�iD�FkH�Dʫ����4�@����9�����_;���H���H���O����O�˓52��Cߠ���'/֋R�b!
�-�v���K㬊��OBu�'[d7��ڟ|%�pj�D�>��a䛌/�Q�1?���ַR\��a����']Z��$���?�QiH!+�)B���Ӟ�S����?i���?q���?��9���8#C$
�����\)_����M�O�Po�����I��Tr�4���yW/I%�G�#��a�P넩�y�&x�ȥm��Xʓ�Ʀ��'��9�p��?1Q�&�X+�H�7#@�x�)�
Q�Ii�'��i>u��ɟd�	�x��u`l�%"S'�zj� �C3�9�'Y6��6���D�O���.�i�ODk#�����T��on�aKvmLv}"*o�l�n��Ɏ���53+�!�D�b8@q��ayH� ��̡8�ɶ���a�'<p�$��'�^��!���Y�v�7R�"�'y2�'����S��Cٴ`)���sW�-��*
�o@X�yQL?�P�2�u��6���jyB�'˛��'b��ach�!aM´�T�?���:�"I 8i����l�� �h~���9�@\k�����T���9o���T2O���O��$�O����Ox�?�1�T>y��*�������� ޟ���ß��۴v̧�?���i��'����A��<#%$��Ѵ������'���+�Mc������՛ƙ�Lr�\{��Rg�!n��%���2c��y���'l&�|�����'���'^�!RuJ:Y�H tR1�䉺��'��^�@�ݴ=�֭
��?9���$5�Cp�tf��eٖv�ɣ��dM֦уܴ�?qt�铝7J�`��F�gy\�AP�E9n`4�ɳ1&!�!�6��擦cJ�l�k��(�e�0^��R��cY�H��ߟ�����)�cy��m��PK��D�^W�<��+�/	�2-�C�-e�L�D�O<�nd��8��I��M�t�ʟ5�̹`/Ч*��QAA�	:�F�'�Xɡt�i~�Ir�^8�w�O��,��s��]�R��`4i�B�!̓���Oz���O����OX��|�qMͅ>�:�7��jP�������V��x��'����'��6=�
���CӦ+�p���	k���g��ʦ��ܴ�?�)O1��a[��v���$g�����r� O�6B�?N�9���'�$l'�<�����',R	3�F�Fܫ2��@SS)ޟ���֟��	ay��m�6�D��O
��O�D2r�#G\�8�3�����ۗ�+�	����O7M�O:ʓs(���A,M36z󌐩t�
5�'�f4�OMjq:���-�̟:e�'���@��J?@���vN��:.>	��'K��'���'��>��	q�>D���,���Y�Ϙ_cq�	��MÑ#�1�?�����4��)�w*Z�V�>9zao~<[C�O���q�h�ҕg�86�!?������ܩ�p`�)]�9��}Cwj֜'�ҡ I>I/O�	�OJ���O2���O��sY�l���Cϼ%Zl��FA�<�պi:&��B�';��'�����	�,�`�# �UJ.� $�Aky�'ᛆ�'�)��_�t911f�OI�Z�����HVb\:>L�q�'$fQZ��D����|�^�T���M�x�$PY�.�+d�R�)ϛҟH�	ß��Iȟ��Syq�����O���HP�=��a��8R1˔,�O�unZ}�I��ɣ�MKҼi�b�ѦB��M��JoF&a���#bՆ���i��	d��Q`��O
q��N��@T��37���=t���b��e���OZ���O��d�O���*�ӤO�<!��8	�Բ�ᗼ$E���P�	 �M1��|R��x���|B�4@m��3%":�z�p��$�V���ٴ3f��O�d�i��I 3���c�D�2gF�s/9bd�R��?p�g�~�Iuy�O�"�'��P
o���6�^�)؀�������'��ɜ�M�ANɷ�?����?a*�X�i%N�u粸�aUq�HM ����0�O�El�M+��江(Hk�dP�p�n�f�� 3�&�6/��ML2�p�	�f��i>��Af[=��I�7!8A���.D�a1~�ؖ@֦^����E��d�5��`�w=݊�Z
ui���.��TX�-����o�8�%�R7B�G�� �E� �UBmБ��O�8`DHI!_��$rs�Z�FHVQ��E*e2e�nO�� S撶b �A��U;Ԯ��C]:q��R>M�2�kD4E,%A����&
���ڥX�< P�N�'�0���&��jdM?^�c��B	ܯL��D�Ђ��X��3&�?)�8	;W�E�-�&�#Ff��s�*,�d	�y���"�>�-O�$.���O�d�#M�8�"�۹{'Ĭc���k����#���O��d�O��+�b���7������̡V����6 G�7�<#��i��	֟�$���I֟ 2�q?-،Rh\*�� �a�O�>��'��'��Q�,F�����I�O�[Ս_e�Tj�Ǉ��D��EƌǦ��IX��ٟ��ɉ����=� $}�"�m�]���N<E���iN�'��I5<�
����d�O����(8@�U�E*�W�Z {��]�a(U%���	��@xЇ@v����$���Z+0,K2��(]A6}�fC��M{/O�Eۦ�D�)����(���?��Ok�/��	SJ�p��M�AG���'Q"�Ŵ�O.�>����Rt.��S�n� ʙ8Yh6m��A��m럘�	֟��Ӓ��d�<QU�.L�^���\�u]�3��3�&���L���d3��Οt{d
/G����6��q���M���?���Ie��9�_��'B�O0��iQ9��U�E�Y3�BE�i�����O�P�Q+}�П�������hT��X�r竇�h6�hb�直�M��(�H�"]�\�'�V�X�i���'��$S!����K�:�$��%�>�H�$���?)���?�/O�qʱ�� d�@�>_J�8��CP�Qz�|�'������%������dz�'ì?������u���c��'M��&�T�����oy��'vv&�Ӷ-��z�M
Di�'*Mഐ4�a��˓�?qK>���?�����~�ݵnAШ��jǖw�顳K.��D�O��d�Or�A�h蘥R?����n�Y�4��O?�	��A4�� ;ش�?IJ>I��?�6���?yQ��e}R��{&v�rP�ƱjW@1������M���?1.O``D}��<�s��8�`Č	Kc㗭q^�p��
9��<��A#�?IO~B�O�
����'g��x��
B�DQ�4����Q$n���s��Ia~�(�d��ae��N���C����M++O>�3���O��%>�Oc��Шs�Z,;r��,o���M�G��f*e��7��O���q����}�i>����3B~L��ɺ:���j��Mk���?���S��'R�ЍZR,��ѢӼgɞ�����)�x6�OX�dy� 
&��O�i>i��G?�&&�#rDH�f���h�y�̦���H�I�������Mۢ�Q�4�Ơ��F�o���㇞ɦ!�ɼe��Ŕ'�L�'��'�*x�@�-b)�xƧΖ"�;`�"�d�"R�1O����<9�n�45y���<���SR�E)̀���O��d(�	ԟ��Z3T�"R
���P�Rǔ�[�qlZ�%��b�`��Yy��'vR�KU؟�-s�L޽#n��	�ʊN�&k��iB�' �O��$�<� ͦ�[$閅l��;�c�L2�p2�2�d�O�ʓ�?q&��9��)�O�2�#X���=Z`H����{�k�ݦ�?�����w�'$����$�~t�&��3coI��4�?q(O��D<?
ʧ�?)����}E��)7�@�N��b%�/"���&���]y���O�L O�61�"��8M�L��J�/P���Y�� A �M;Y?Y��?�A�Ot�u�ՕM��ix�E
��``W�i��	�,�ɱ��'��禡���W�j{J�"��	�o¬�Q��oӚIaFM�ɦ������?i)I<ͧF��M���?�L�f�&`���i�i��'��|ʟ��O��Hƒ>#� :��1[��-�w��O����O"牉W���&����p�}�蠃��^�WO"$h�Ⴡ6� 9n�ן�'��r����O���O��q&B<`X��x��������A���T��"�>1.O��d�<9���'̙���\r톏9�4����Ht}ҡ�y��'Er�'r�'�剉9:B�#��!Vx5�1��y�f��������<������Oj�$�Of�Xcn��J�D�Y��6��t�I�W���O��D�O��d�OJ˓9T��)e8�깂COB%���b�T;D‌A�ix�Οl�'yR�';BHD�y��ޅZ64ʆ�nު���'��b�H7m�OB�$�O��d�<�cA7����֘;'C��@2�Z�Kf~�jݮ �d7M�O���?���?ib��<	-O�e�f����-��B&^��y��c�y����O"ʓ@���a�P?i����D�=f�TG:<Z,��"Z&����O��$�OЙr";O���<9�O[<5yP�%P�d��iتT�lZ�4��D�|°�n����I埨��������;gC�)}�r��V�D�i���''P$0�'�\��<i���bA�T��S�/܃]i���ȓ��M#'I��i�v�'�r�'l��O�>�/O����J/|T sf��1	t�#��֦��Ю`�T&�X���&��I���0?������T`8���i�R�'��˝GlR����O��	�	h�������Z�E�'�6m�O�ʓ5OZ��S���'p"�'hLrrN�d��4��,����AD~ӌ���eThh�'��	㟜�'�Zc����|�*Q�ä7%���+�O� (!?O�˓�?9��?�.O<U���Y��!��L��������>�����?���Ә��'&j��@#Zv*�A��<i*O��D�Oh���<��I�@2�ɑ<O�|L���/% `< ���]0�'+R�|��'*bN�/��ɗ'M�p����#C~ 0ke@�>���?�����$��q�$>1Q"��j����6f��$ѓ��Յ�M�����?���0�^h�{��I�f�3L����B#�M3��?q.O"0��D^B������4�"�j�$��W[L��sO<���?!�h��<�K>a�O��䋑�D�Tm}��F;G�)��4��DH764n�����Ot�i�c~I�0U�uX��Jw���S'�M��?1&���<�L>���  ��bc������q-�L����v�i� ݛf,r�.�$�O����|H&�t���������<N�(IvL�1���޴O6$�Γ����O�R��G��� P�[�u_��9 m]�7��6m�O��d�OTt���CX�ן,��C?�Ղ͞?;8�(�a^4L*Be�e+���%�Dۓcr��'�?!���?i��ZQ� �N2m�8��C��'��'|��J&8��O:�d&���ܴ� m �p�f��+��H ��BP�$�1aa�L�'��'""Y�02�cɉ�th:�,!N����Ou�|��}��'��'v��'=h������B�P��RŐ+ ��}��(��y"\����8��py�`
e4�S8=���'�^�8X
�j�f[�_�^듻?������?���N:���EP�,@3 ��I8���֥�7�( 7\�T�I����xy���$~7����F��5Y����ܖR����L�ᦹ�Iv��ꟼ��hˌ�	t���!"f��he�Xz��S+1g�V�'�rP��
�����'�?!�'*f��R��5O���w�ԆLI�L�T�|�I��`�I�g#���f�	GB�	�&�ře"���,�w&HΦ5�'oPY��y����O�r�Ou��2{�u��	�F�` 0G$����lZ��0�	�Z����~�ILܧ8$���c�ݏ)�0��'-Τg�Ԑoڑ[3�9��4�?����?y�'[?�O��0Wo��6�>�x��*��`��O��q5�YG���OzrA8�H�"s��:I���Z4�`7��O,��O�lq�"�l쓊?A�'(���H�{�-��X��쭪�4��t@��S���'���'��l�sIж<�yv$�����
��k�,��� �~��>������c�0I�< ����֜:'NR|}⮝'R��V�������[y҉IAd��H��W��stkT.)<�� �Iן�'���	ן�!��EL���RȊ�{d|��wE� �H�	my��'S2�'���;F|�O������~;}�pz�M�Oj��3ړ�?!�)T��?��aĬ yj��1
"^�� p,��GV��'
�'$�X��a&���'!y�M�rnY-AT�\�oH�I�Z1kӾiўp�ɐK����	韰�PW5�e�J�fջ�Ф^��4oZ� ��lyR��=+c����k�٣sR��@���ƅIc!Z�O��d	)�L��'�T?!����n�0A8�N�t����FhӐ���O�P����O��d�O��������Okl	+/^D�S�L	H��h�`	�(���'}Bm%�O&�>iH���:[0��d�-L7�KB̝"�K B�s��cG� �|N�i-�
��]qǀO�DP�qpKV(hF*i��*�Ua��
pI�I�T%Y� ��T;R�Z\��@�ץ��By��j��H�9I��!$�	dq�I�&^�<���{��_<�H`�%\�~�������X14�P�<@�����$#�@�T�3�� B'Y�j��!)s��DdA��	���e���A��hI�(C��\��A9Cж`����?���?����d�O�擓R���#���W�<2�D��o ��Y�B�5"ā��;U"؅�FG����O������H�@�"�$<ߠ�;�j�y�lKcL� L�����9�衱!����x�U����Գ��\�������y��d�OL�=)��DkB�Z4�S(r��qQ6n�(�yR!�;oܖ�Y�H\�R���q���'꓆�LJ��'!r─h��:��I� qC6b��'zB�'p����'3�1�����ڱY���+$�݄'t�7��3x��G��[t0�i
@�x�C�g$�Q��h@7qN� ��i����.��6�|y���3E��u��CnD�	��'D�{�P?z� p���ߦ?�z�y��'W.�3�:V���8Տ9��ě�'��7��^dJ�i7��f�����ޒ\e�<�B�y��	�0�OH
=)��'2x��AL�,�����;(�rЈ"�'}���$a���C��G�`J3��O��n����D������Qل���c���	�0�`�(�gJ�5 ��Q$Yq�O.f\G��7b�,�%�1!��́J�<A�K�Or��#ڧ�?�q���n*�ې��U��,��%�ȓ�{�ő-��Pr��11��	�HO�ștBʸD����1�ȭ6�,�Ĉ���e�I���	��Z��G�֟��Iɟ����}�a+х+,ze���Qul��W�(���ɑV��ӠM�+�<b>�OJ�RPLk���
qA���4�L�7�����O�HIC�3����N�8��6v��0$�O�QF��yR.O��?�}&������(�FuS&�ާa�8���9D��Cwo(s��d��!�)AX�:D�*?1��)§m�vdAP&\�=��ݣ���'a�V�H���2����?	���yB����d�O�"4�,�"���w�4FОx~���Bb�)"��z�͝�w
�q��	�-P���SHIu����W�s������B4	�J�P���-�i�牵�"Uh��
�cj��Ə���9� �O����O����b*��M���4��d#/T�iu�sФ��]� ��i �"+���D�<)���"?��'g���R=a�@{q��sFɄ�%�r<O����'�"?�܁s"�'{ɧ� �加��E���RE
V�����')�Q:�Bj�_��d��C���4����p<��Iݟt%���M�6@݄�ġ߹ U"�R�G!D����/�=7�DH�B��4^��Dy��#�@iش��-A@��8��MrvLӗR�$�<����QS�f�'-�?U���O� �CٚqY �aH��pV4�B���OT��.��d#�|�'�Ȥ"�T����)�#&)[�M�����+�S��t@�y�EV1X�Y���;�bħOl����'Q1O�\Њ3L�3[Z$3#&�.�13@"O@ӥDa��u��$�!5�$=���'�,#=���W(@�8�AD�(�
S��I\���'�'��RQI�.Z��'T�?O'n���x	P#��*\�i(�G�\�1OP�I��'�t���A�z>�$!R�Ɲ5��x�{���<�f�ųUb8�It�;�&��V͙$�'�.���S�g�u5����΅��J��QE��'V�B�	(�i#d(�4 �<HJs1�����"|jC��L� ��cs�A�� B�ci��;�?A���?��'6�.�O��$c>���˕8L�Lj�JZ���@ �
��pB�	 ~�k5�X�ɻ@O�$i�e;��K5&B\�<�g�6�*���$:*��#�O�H"A�V5�-�B8�}K"O��EK�9b�iS�P,?�$���$�S�S8���i��'�0ˢ�E3�D�V&^�i�氱��'���9lnB�'���TsW�|��Isw�ad��\@�Qf�W��p<�E �D�X%j9B6�P�Q"����G�#j���	�AaN�D(�d¡p����Y2e��Hó*E��!�Ĕ8P�le����F���r
R�:!�$KǦ�f���hM���퓚{12};�g1�əv{�e3۴�?y���	��E�B"V�	�p �L�Nip}���f.��'�@����'O1O�3?A��7�Б wk�$@����E��V�=���?iy�%HNc��S����Yc�b'}�'\#�?�y����	<d���Q傁kcx9Z���y"��,�P�Ν�n����[��0<�F�4N�rAXS��[��5
�� f��P�ش�?i��?�Ѫin����?i���y��7iL�)��9�PaHU�	o��dp�y"��<���gy�B
]7?�L�����<�`���5~I��O�a�@�$
���<� ���>�OR�a��!���'(�K�<�6"O�=h��/B9,�r`F>!�Z����i����*1�4ڣ�BjXK%C�o �Z#�͌<B*�I����	�,�_w
B�'^�)ǐWTE�W$�k���C�_�N��FO����_=yed(ҳA��]�\-2�*�a�!��=y;������z箙&��>G\x���'�"�|��'�B���-y�>4�6��F��AK��P�J!�P�66�]�c�Tb��݁�Ζz�1O4 �'���4,�RqHش�?1�\v�$��F@v ���w��5q��a����yrjA��?A����ԢMD����Z�N�<�uB¼I�/X����h�d��	.�}P��
�H��f�Ɉ���L<Q�J ��E�r�x`K��'�L������a�[]�n0[Ө�� N<(��_-�]�c%�.6��
d)ѩ9+���� қ�]�W��<��@�b�$�jD^���'A=�'.nӎ�D�O�;v�	�9��q@���v���FQ[_��I���џP�<����<i8l$���خ$����Ѭ 5�~&����E�;Pg�d�t�*�F�2iR��ΐb���R�k�+0��Oz٣��'1O��`�	 )R��M1����4���"O��x&�Y/WV$�KV��R��E�P�9��|�!�I�~�@�#u�'HС"V�S<<~L��4�?���?Pm��
zT�J��?A��y�;W��y���0��c�$��j�y�y�����<iG. 09�/@2hs-�/�U��N���	9QPxeS�������3*�!o���<�s*����>�O8,�HJ�c,ؘxRlͭV�hp02"O��e�ݒV"�P����xp�r������ᓘ����'=����ꞼOk TB4���}�	՟P�I�<\w���'���#\��S�J�P�j���H
�mGJh@�O&q� ԍr���C�a0C��-&ܨ��1��R��j����b��q��g����f��5�O$��ա�9Ybq�6 �m�vQ
 "O��7��n����AR�s�(�*�u�O��Xs�i��'�yȦ(� ��L�w 	B\����'��d	x��'���F��!�&��fg�i86|�`q1s:Z����O�a�jS��'��A 臶����"o3���N�Y��i�k�(m�u2f)�p<�c���$��WJ�Q���ѧ�Qa^��ǡ(D���(�!2�ޝ�È-N>����2�P޴)m0lH �r$��8�
��^��<��ţ.���'-2�?��V"�Od�Ӏ/�P�\da���k�H��� �O��ć�'j���4�|�'�~�b�&]r�-(�
W�8�~�K�D"�9�S��=.������?��㶅_]���O����'�1O�xC��$zB*q��n	29_��"O�8���E�1R~�Ň�
O�웶�'�"=1�Ê�0@IWD�Y��tQ)�'p��6�'���'P�a���+9?B�'���y�f��qΉy��L�7�"�s��?^	�'��\z!�$glџ(`Մ��"�)���TsDS�m"[r�^�(D�qAA�B��>1��AV���$�`֘qn!u��E��%�Lfum�
�M�g�8u��8T�������h�&E2,_0��%�N�BJ�{b��OT��ʜuqʍ�vh�1�4���فy��I��M�%�i��+n����|�-���
p�\�
4F1�m
�xs$\3��-Xp�jG��O����O��ۺ���?1�Oqjܠ��	��u2eh�b�J�`��ܿ�BKaEW�a�Ԥ	��IT8�hr��� tR���/	�
�qǭ�l��p#!���=9�̀C��x���
a�Bْ6�BXդs���	�?�5�i�Z7M0�I���OC@��&������� �bLK�'�X�i�.V�P��YpC�(%�B̒�y���>A�yҙ�Į��$���}����o���y��T�t[ȼ�� �4|
�<Q��N$�y����f�N��kZ@R����)�yr����++��?)�a�t)�.�yR̟"��m��Dؐ4n��4Mď�y���<ߢ5�FK74��-`�����y"�"w~f�{������C�O)�y"�,��I�S���^V)��_��yңܿ7>�%h�T5m����W�7�y"(UZ{tX@�ۖk������y�����u�\$d%�4j�)՝�yBNr���3�Y�s ��0����y҆ʹ0A�:eHȶpFf���y��tE��x�A��	�Q����y��+w�`�q��c����� �y��e�y����`�~����:�yr��)�DY3�I�VȔ�Ӡ͛:�y�c�w8��g�L$oͩ���yBo]	��2񨃻s�&�j���y-q���B !6��l�7�ԏ�yB�D�
���5��@�Q.�yb��;Dj$a�cK. �,�ъע�y�eT7LK@0�͘�u`�䀴����yrGτ1и@k�o�.u��������y�٠r���O��g�@�E�L��y�63X�x"0jk�NX�U*�y�A�_j���w��!��ʈ��yB㕋9�6 ��_#j<T��u���yB7l�.���n�>h	,����:�y�
͖}<vu��8����
I�y��� �VT3�]�6��z��ߏJR)R���3�g?��	ή0d��k��0~���# �H�<	��.ԱUaK w���Çϟ��a�@_a}�	������~g�٩�j���=��������_���l��-6Uذ� b�쐅ȓC�脲O�^�#"�D5s��0�?��N�"��#�a�1� �"��x�aّ�Y�<� >��ܪ_�DY���b��1��BXh؍�=����O�Y#�j�64��B�%>:��)�"O�a��/�8i�&'U-��&�'2N�Q��tX��j`�����sm��d��|�B>�O��T^d�Iюļ.M�Aᔊ��""O��ǋ�=S��PP%��K�l	R"O<y����
4%���D��U���J�"Oj��q�J���APE\�Z����A"ON�	�͂�a�<�B�
k�L9�"O���e�#՘��̅2�z��u"O�� �%D�uL�؁��#:�0�8�"O�Z�O<�D���)f�(�"O�4(� ۺ:�V]`�`֦}�y�5"OH|�bb@��h�B��\��)ð"O�5�ro��a8���O�GU|P��"O� �t��L�D��L�/Q�e�"O�x���P��Tk��]f��	i�'TƐ����<-n���[��`"
�'ւU�'fT�9 �����:
���
�'�*��O[����3���L	�'�&iY��������x���'\��JG�@���n�4l2���'>�ld��O8=J#N��c��	�'��7hǊZ�(�i2�;
��4 
�'0X�,\�^6$�s�hP
���k�'?�Ey�@W��ʘr�G��Z��X�
�'s���w�P��æ,�$�*42�'k`�
�4J����ԓ{=`�(�'j�1���-:4>�%�مj2�`�	�'OhXb0�I�pM�K�A��dP0	�'Ȅ4��"ހ�f@4��._����'���zp�;ET!U�C�V�b1�
�'gN�j$��$(��[Ĩ��N���S
�'����1S�<uDm`��HB���'ʺ���îs�t��w�M�58�Y��'[�\�
��V��
��^�v�K�'��Q�*Y�%�В��S8�����'�X�9 �I�K-�M�Q���	�@�X	�'&ܘ��ZO܀�XPb�|��qB�'z��fH�	޶����%w�Z��'c��9�k	>�<h�ፁ�"EDh��'	nx!5`��Z�PA��,�AxA�'� ���K�LY��J�t��'��}�4� ��h�Cw�+hn@��'V�c.�	��`�d&^��]��}�$��আ#���lA��nC�	�wx���2D�g��_�C�/̆؈���9��!�ujO> H�C��-Ė�1c��{�U��&ۢ01�$[��7�����_�ΰ>��ԎN'�u���טS���!��G�Tz�$A�ּ��	���L�C�l�"�e��KFvИ���uN��b���/�)�����I����'WF�) K�6��'�(�'mٮ�pU��>�&��Ȑ��ܩ��!�>a�L۴ݘ\��bQ�L�~�QR��Y��	��D
t#/�3�Ix����9��N4@��ɷDC��x�_1hFP� �;���ʲBJ#s�Xy�aX
�#*=�OL�&ēp�� H��T�I�\)p�')���DA� �JlfJ�>���G�<��ݠCfNj�j!-BA�<I�E�/)��
�g�*y�+D�F~���\�kֈ[1��"�&K-��ɑ+[#05j����E�<鴏�L�9چm͞W"!���J�H��P����	�| �c>c��qC�Zd�a�+R'5��4B�%<��1Åی@����`R�F��3�)~��HT^n0�)�tB*�UC��8�9Iҡ*r�H�ቪZ����H�
�@�#�O� ���Q�@�j�=��c̾�&0 �"O�����
(I��]�Kk`LRq��p�@Kй����$♲�ȟ�	�"G�
�VJZI�" � "O4��&lY��Ы���q����u@R�hʆ��'� �Õ/����Ϙ'O�u���Y� H-9j�KHf8��'G�U�q�ʩW��@"�!��M"��V$���:E���
,���$���eIGj��%G|�˄A�=B:ax�-J8V#�yb+_$R��4 LrU-^�r���G�	�j�ȓ:_*a���;���I���U���J�JΕ�Wp��ӭ:�*$�ȓ>��Eh'�&��`��HU�9�Z��ȓT��8 Q��#!����ũͦ$
�}�'����M�6$S��3�eq�(�5B��a��O�b����"O�0ۣ�
ڰ� �� 7p2i���}Z��	%h_���A���g�A�A�
�9�� �]���ɟ<�X�'��=MqFU[��A�n�0��@�fL����oE�E^��a���p=�֌��w�@l˂)�?���CL��	7�,�fbӚ����-� ��&�ֲA\�Aȑ� )I�I3n�3R�ؖ$� ��|
	�'؄tj��ůMG�I��CJ�z�B�MI妵���	S~iKPGJ�u*��PZ���DZ�~�R�Q�w���X��ɈQ�(��Aʩy�����'��A��$�V�t`ܞl���8�!:Prz`��a�mGF��	�w�!�&�u�g¡1��$8���<)�
(sW̩�G≃*�Y�To�`x����∁.��ɀ"���&�<�$T��F�NN���FZ�Oz�8��DR�
��[f�Ϳ{�$$���c�'���
"�۷HTxf=�\kH>9�À5�|�'_RQ"U�=H˞��t�YoU1�-ь	?e ւZ�Ae����_%�̛�+ �OTXS'�7U�jt`"�
�]×O�7��z�	:�FuT���AM�z�	�źi����w�(�����;ɂ�2�q� ]��'}��cC�FA��3��^���eT2�Āj�#�� ���O��#�C4�d�����ɍ3�L=�1퍃E>6����ݛ~���䌁A6&���O�x%*�7]���SCJ�S�P�xQo���?�։S�X�$�9#�w5�I{!"�W�';ณ' C�]��Yш��P8BN>IQ��{�@�&;r��?֠s�`,2�� �E1�nPK��\��|���JQ>�^���'�򨑕(�!~��q�e;LE�g..?��6xBf�Ȁ�E.Ur�d;�cX�y"l��l��Γ	4H#@l��;}� �p��!�*J��u �"�$���E�۹no����EG5R�Ia�e�>yG�l�*�1�D��r�����͙%hf�H3�ѧ*�Rg�;���]�H|��ص�ݍw�.y����}��6��3X;�����/��GǾx��T*�ͨo&�CM7n���Z�, O��
$d-\���'J{�*��b��XCR��l�R�2
��".�9*r�:�O&��A��ڐ�D�8L)r�	w�>!Q�^0R����ğ\z��L�<%?Y���v�	�e��B�>8�"n#D�����>=t�J�lޅ� lNh���ɳw�xݴp����~b���K���4�r �c�! �"�?$�x���Ŵ3��y��ì_� ��BE�^M9�����y���q�4��㉄<�R�pA��>.���D@(�O�����)�$)ߒT�����mQ�Q�n�����J��:$��ScRL��b��A�0����+�	p��X�N�Q����DS0]���{�۶>��ҥ�'4�H�Ѓ���V!Yw��3$���K2*�
5|���Zi�Pa�.�V"X�9!)T����{^2x�<�S�%��S�� X���\z�<����7�A���$km��;�Őu�&oe���?�}��Ԝ=�������Z�����x�<�̍�p� �SE�a�6IH�h�6�@	�{�^5�s�LX���I������Ɠ"�朙�I�]�=�A	�#MW`�H�oϛ�x�~���H�T�_��`w�'��<	��U�ۘ'q�yZ�(@t{X�2ue�_���#�'Ή�sd�3;��#P�V� M>��#Q�����O��2�Õ�hI���dQ�ɸ�'�HHBK���(O�=H|R�r��K�axr��0w"��)��_�Vg�41��Y��yF�,y~E�F`K�`�>�pVȂ5it���'�2��F�R��D�5LO!b���[��� ~i0�٬3�p1"��5#�\yA"O��R[�3�5���S��Hj"OȰʳ	�=s��sc��{�s�"O�<k�b�����$.$����"O2�0D��0V���%W1m�%B�"O~�2A":8Hђ 5NB�@"O�%+@� � �Hc�"�2���s�"O�)#R�ڇ��A(c��77ED1�"O�� ����&���Z���>5`H� "O��#g�گ4q���<o�h8"Oh�CR �uV�y�ڧ\���A"O��XI ���ՠ�7x�v] �"O� �"3f��8рދ_�؀��"O�}��h�xU�PpQ��%YÖQ�"O��(�D>[¤�a�4�(��#"O�=9���7�,كF�Y��P��"O�5;�g�:DH��en.L�:�"O�;g(ü{|0Y�U��,70�5"O"=���? ��c���_4�К�"Oހ!@L�x�:݃��kA���ȓ%�d��I>8���� >�|��ȓj���p� A�b�\��c�J2����*��"�Ӧtց�j�JkB��0��Pp�_�-���b򇙌h�ZL�ȓ?�Ƽ�F���(��ځ�4M ��ȓ}:�TDIܓYG6�W��c}�̅ȓH��HeM�M�l��ȓ2��ٚC��@�i�4옅+�d��7J�\j����򨪴擺m��C�	!y�bqP ��(I��xa3c�mhtC�'.NHP�E�Η2�V��ga�$�C�;Õu��:c�p�-�4�J���'�\�6f��Z-~�"�*���I�'�<9���"V�X\cGCD'��đ�'Z��`n�b����ʍ�lc��
�'y@Q��ٵ;��Z���i��Ur
�'xZ��6"�?�����%`�����'i$4{��;D�h0
�,K=��Z	�' �� �iI�Wj>lS+ʺH�`y2	�'�80q��L�4�(<	׮ծ���	�'��hsO�[�� �-F�Y�l��'��UUhQ1W1<q���4t��"�'�x����4q$��đ#tB���'��`��C��)�L�g�J�nVu�
�'�j�ғ"C�A�4��C�
b���9
�'��]*�D�(Cfl���F��YB	�'����5#\	�������=��'D�x��^�QD�U��<�
�'�9SV� ��3t.�<t����	�'���#eı>���F��gX&��	�'��p�0%GWCL�!�팉h�,���'�@ē�+:n��%� Ƹ�b�J�'���i�f��<'0,�D	����	�'��X�.�-Y"ܽ�3�!,Y�	�'RDP0%�X ;�6���%8%�6�	�'����P.؎oj�`R�bH�"`K�'�%�ф���\�� �F��t��'�=+P��h$��b�)|E�q�'d<ɥF�f:U�5�ʅ
��!�
�'<������5��6w�K
�'2t�%�5w�2�M�}��y	�'b��v�0I��!��|d�l�	�'6�}z��X1l�.5j �S�f�4��'�(��G?s�$���L8KP5���� ��H�%C0m��UI� U_����"OH�h��ۍ^a ���,�bh�"O��:�gS�{	Ĝ�a�_�+�1"OD)��A�=Mcr�c�i͉"ɴj�"Oj1��nɸ*ݘ ���YZ�8<&"O��=@D9��I�7�H]ٴ"O�a�e, �gv(!���#C��� 0"OF�{�/�>Ø5)�ɞ+����$"OČ�!J]�S���"ń���"O0��F�� �2���s�x�zr"O,đ��.��AAAW;1����7"O����^L�`L�s��(`�"Op�J�k�B	w�x]�a�Q�n'!򤕀<-��жm��5����r���5!��%
Y(y�� H�d�F��.��'w�KBV��p6nɂq⨠
�'2P��pq1S��l�C�'jzG/S�7���c�6g��t��'B������ X��Ǥa6m0�'�R���9d�3�� h�օ��'�^]CB+ٿ=~�s)�,� t��'�졺��?~� |:C'T xRt���'��p�0u�xI)sDƟ^����'��	I2�@e<�d�r��*[�4i��'����'�+*��̊Rf�� I�Z�'9h̡�셒Lg:EӴ��FMs�' cG!/	�H8���<#V����'7`��M�T)�8��O�6-�Q��'�ڼhT���0�P�DȞ;֍ӷ"O<�t��0#�&Ŋ��M;�4�p"O��֎�,]�uS�J�A��"O挹���l�΀��nVd@z��"Ol����y:�MB��FL�"O��`� ��~x�Yp*�^���"O"�;�ٴ*pڙ�w��{°!)�"O��2c'S4L�� rU�"`��ѧ"O�����<�� �޾\�61��"O�	���Q�������8>��9"O���j�VlH`V�O;*L@誇"O�`�!C)r�S�J�(��IT"O��!�_`� ɗ��J�Z�"O�$c M��l06k(��y��"O�)��%�<&����c-�:��5"O�C��
C��dL@Q�`��"O��&�X?��#ҥZ�v!(�"Ov�U-Ԅ,�x!J���>(j$|��"OzY�"BH�A����-aT �t"O8�&�P�8����ˏ:Q�=�"O�� "	Ӧ!���q��R=I��"O���qN�����L*=
��"OtH�'�,#��9�')p�8T"O�I�FL�L|�[wH	}�����"O&�:Cۥs�+���i��@��"OX��ՌJ�N�v����ё�2� v"O���$�=���{!�˪^�P��%"O�����N�/g��bTDڂl��m1`"Ovi��(�2f���[`Iʯ�ha��"O�P��L��N����ޕM>�P��"Of����tB6%�q�LT@� �"OQ���/ x�����:=����"O4�E
U%5V�e��`�;�$��"O�u�g��L9$��pnފ ��$��"O���6Mכ@��r2Hvs<UB�"On���§q�ĭxlד%X�ʢ"O� $�3�i�>7G���E_�\M�T;"O��0���"`1��d��2~�j�"O2����"`�t�h D�y(�La�"O�9�>g29P�a���A:Q"O(@�Q�X>s>������*6���	�"Op�����)�$��ە=�Ȁ�"O�26'] ]�zT�#\{J���"OB�H����a�#E(4Fѥ"Ov��c- 0l��1$�.��2�"O dh�o��?�聶��A�`�×"O*İ��"/*ё�Y�E��X��H-�S��y�O������W7f�d�'9�yjĈ'ټm�f^-4Z\l�4/�y�#NT��y8`�L+;�t:����yR��;|M��ӡ��Cg���\�y�]�I0%I�`b�X��J��y�`Hm��Y+U�
2���u�F�yb�>b.��p�@|r��`� ���y��N�g��x���v6���k��y�I�a����G�@�Ĥ�Uf���y"�)_@�-PË��m�f��V����M��4丧�Ol����O�q\��r�`?=�*���'��[�i�u�t�K��ݣ�
P���/qs(���O� YD�)N��i� U`|��K�"Od�SQ߭0P�� �.2q\��X</���X8�����)����W���.q���M)lO��JM>IӮ�u>���"@�a�v(9��M�<m���X�"I�*V�6!�f
@ܓ��FxJ~r�b�;z3�)��"�{��8{ͅz�<Iu"�++}е�צW8e���rǏv�<��KI�:�N�¡˃5�F��y�<��I�Kyty*Q�,eL���s�<Q��O�Fk�̣3��P�2͹2�T�<�f.ߔ{{�ݲ�2=���a*�S�<1��1�DC��
^}P���j��hO�O����dI.7�@���JŒ�t"
�'^��Qg 
��֜`�6wd�k�')��!

�~����"�ҟ[����'�z�#�R�R�n	XG�ܷr� ��'d���v�Žs�Y��B���9 �'�|�����f� Y�!��!��'���`c ^fk�h�X,��'��ܫ�E+M��QbL8jI��K�'�v$a��(�M��-��]�f�ѯ($��Se[4\�*�P<-���uc-D��0���C����t��\D1"��&D�L��h�$���6�]M�� 11�*D���b+C	
�,�Ӯ�Q��؀J.D���D�1�~�+1i J$1	@�/D�A�����P�cU *D��G�i�`�@�*�!�:�K��(��<�C͖;y�B���ǌ*���CagNF�<qE%
I"P$���	��[�DK|�<!!�
}0H��Cӂ(EP�{�MHt�<�B�
S�rr d�&N��!��j�<��� �6��rE�98n �
�c�<���8F:�0b�������h��@c�<qc�N�7)"�B#�F�}.�����`�<!�+ݳl`�*��՗|W��8u�P_�<�)�%/��8�k�8_���2�b�^�<�a�  \�"��H4`)��:%)I\�<�D�C�a���f�vB0:�!I`�<)�EP�o�h�
7o���j���u�<�7�\C�����Q�sb��n�<� &1xQH��_��ᗍʯ��Ļ�"O�iC�A4	�������m��@�"O�][Gaڤ((X�J:-�<�3"OL �Re�j1��B@�Q8^�̨
�"O�Q�����Py��
"�\�˦"O���$�-aP�S#L'�p�4"O�dR���Eb�$�ʏN�Lpp�"O��1ド���	��D6ZȁU"O(ura���hS�����n-T�y5"O<�5���4x�L�p���O)d��"Or����F�<F�+&�O���"O\�wI�&�(��Ѣӯ8�Hi""O�
�ܹVE���c����#"O��t`�@�$L�#�Er<���&"O2�(d�$c}�C�F'p,��c"O�1��'M)	{84c3k��l�@�"O�uH�o�,_*m�/�xvh��"OV����\~< p-L6rf�M(�"O���1�3�tA�ʍ��l[�"O 	�֍á޲	S ɛ�w��<�&"O�,RclP�M����N L����"O�����zG�5y��G����Q�"Ol�Y����|�&�zU�F7 �r"O��ٓ�:'�y@N�frY{�"O��I���r"��`����K	��k3"O�TS���G��)��Ú���""O(Tb��|���j
�x�`"O���\C���`��m��h�p"O)ǃ��F��1���m�"OP�z��ŕQ8 j��@�[ȥ�"O�Ȧ�������#ÌB�xɶ"O�0����=|ހ�r�`�z&�a�"O�-i�˛�Ľ�D��(��r�"O��؂�P���h�E��
��؂"O�᪥č�wS�=0���:)�
TXa"Oޡ�W�W�q
F�R$�)�(�h%"OA�3O��KN�����`C�xsG"O�e��/N�@��@���f.�;S"O�q���2j�t]j�	 �=�"OPM£�Q�\��3�&�<��d"OR	K��,��Xa��?(W$Ii!"O&u�!f�<Z���nI�l\B� �"O�$Ca%�u7� �G.��]�4��w"O���K	(t��ҍ�h�D&"O[���$����mB��ey�"Or�`���?8 �س-ǭR��X��"O��1�菮9���уm/U|��s�"Oސ	��[2��ό#Վ��U"Of4�T�3�U�̋8$�yC"O��b�)B�Q4�~�`"O
��0(+MBe�1O�'��x��"O,]{�cC�O�0�SD�"o��XW"O���!H�- C����̀�94"O���,���+�f��(Z�"OF�Q��Ȝw�(A��iZ;�Z�"O���&�<j�lbj�����"O�h����gq�Iu�	.i�	u*O��*���%�D��AΦAR��'�H`�GꚺM�@��nX�7u� h�'�"�PPFF!mH�t�3]�Y2�'�iPcQ$R�bM�
 T��i��'$�(�'��e�$q#�b4$�9�'�,-����<�$�3��N�L
4�b�'�FP�7�Ō'����ま<��ܚ��� ��ͯ~��(s��*n����"O��kFb- ��B BT�YR+�"O"���6�xq�`N	MR ��6"O$A	��2�"��2.��Oj0�Rp"O4��3J?7�2!�d�J�A\�$Rd"O"�Vg����|�`�$X�\�"O�4�6�̬&t��y���n೤"OjȠ�g��<&8�g�D�h�ठE"O�p� �݂I�Ƹ�FF�����"O4@ ,Ķ~N�P��"�+�^��G"O��@�kQ!Gf��a˜TZfq��"O�}��N< �X[4뛟I,R�"O6�yD.�=�}���I񀔩��9D��aGC�kxb�K�m�`L�v�4D� 藃Қ�А�f@�w$D1�g4D��"��|�Q%fI�򀝈�!���kG� �'��&�p񕠇��!򤁝%��m�s*��R��9A�n�!��_-Z8���� O�N�9v���.�!�DP�"mF �D���/��df�ٙ!��4V�#��ԠSE�t{7 C�T!�I���A�c��7)�A�'
�"O=!�D'GKz�J� ܉.Z�p&�2.]!�$W�O���Y��
D��W��<O!�D���)@�ƫ X�ȷj�"_!�d�:$kf�
'I�W�J�+��%\!��
9G��#�BM��rE1�h��Q!�8c)����n���U��"k!�F�v�L!���*$RȺ�&<f�!��,�*WM�#]	|�`d��']�!�$��Y,z���.ׂ !�]�%��!���?��0DA�f�ڵ�V�%z\!���3��Y�eo](�T��텥Q!�D��#���G(=�6h�dK ]!�ե��`#�/G�8�~HP���"&`!�$Ksj���#��@M��/��ea!�DY�$��+�A��N���B���d^!�D��[3N�*��5b��L�T-�2*�!�$.����%f�!�U0O�!����C��s��Q4OeܕP���Sj!��D9�4��S*P�xu������`O!���.oYP��B��q���sa�mD!�$\��BaD��	Vu^��w��/!�!���#��e��wfn��J��t"!�dڨ�h�s�^� ��8�A��4w!�DCs��F���S͂Tz�M'�!�d�'z/f����Q�
	;E�$Z�!�$P'I��ZU��LpG<G�!�dI$
i� H��
��$�A3@�>!���Ac���g�.��W�	c�!�Ke���BF�H9W��1z����Xl!��W���,��;!������v{!�䈪d3` ��m�jn|XdM"}A!�D�+^^$<3�@�"m]�Y��N�~�!��DG?Y���]�#$�m�FdY$k!��Ҋ��PB��_<7�8���'1�!�$�V�X�ҭ��u�y�@���Kv!�d����e��?" �0q���E!���e%�-1u�|�������%D�!�$IP�M0��(�n��#��wx!�D�'h�2�`���LѼ-R���nk!�d���űg��_�dm&fۀbP!��T�&a�vi�i��	���*o!���H�� �C����ud�*j!�� *����S vB�9K'�[�)�H�W"Oh��܆�섢�H�/#����C"O(�p�gҠ_;��G8���:E"O
%�ժ�1K�myae\0dàɉ�"O q2�\>�~T�A�И/�����"ON�pr��:x��p�_�^���"Oa�sNC�)�R�A�@�7+zT�Z�"O�L��I-�Ҝ��̋�;i8!��"Ol�����UQ�0+!�1d�~�r�"Om:B�R�]��{$D<M�Ƶ)�"O��2	�
<�X#'�W9q�U��"OH��j��bx���w)�@8"O��2�&żs�Y9sς&o>}Ha"O���o�v���ط�@5f��)w"O⤯���8M���ؒQc�`h�"O8EeC��e��a��[!YQ�)�"O��چ*%�B�@%�_�6촜'"O��5��$�BܱuJI9N�>ؘ�"O����&�8qj<�/�1 ƺ	0�"O�Hk�`�T����Ө5аh� "OP���oY�*=�$o�)]�u�"O�=���Y,����QF����"O��.�I�1fh���A^y�!�[��` yvhͦ9X$�3Q �@�!���B@�b��><ZL���3�!��
��Xq�6�TN����b/A�%�!��G_ (*� ��-�VIۆk߽Q�!��D}�ȱ���78wQ�Ф^8D�!�$Q�������6�`�b#�!�$� +����(��t ����!��[�iETz�BW�*��q �Z8RU!�$J2NA~�1%���߄�XĭW�ct!�D�)���P#,���0�Nټp!�d��8b�}I`��8��&LPv8!���/��������u&@T��4!��C�,Ѡɏ)�
���O�~!��
�,,������tB׉՛!�D�%�$ố������k�!�D��/�T� 4��s��C(�5D!��1d�8�R-ŭ1�bE�ʵD-!�J<>����$!q�j8C��z+!��BG���S �V0Q2��Ro!�䉝v�Z!{*�jdŪ�@�aV��䎃ft\T:�/�`"��3l՛6�0B�ɚ\�j�*b� >�4�1��X�+IB�	!o*8Q�a�A����`��8"�B�	'8�L�y2D�
{I��(F��N��C�	�	Lt�S-�@�q�LC+}�C�:P���
�M�xw��I��2_�C��0{��C�	�:]�L�񯔢WE�C�I�[��U�sf϶5�ڐ��&z56�O���� $F4=9��?<�B�fצ.�!��"@��L�L,(<"х^�g�!�Ĕ�W�Lq3��A	��
�'�!�䖉Ә��G�T`��d�Jf!�_k`pxS
����
��<M!�DU�^�28�.�!�4�J�I�=!�dE�f�N��s�+���z�"M={�!�՘O���� cOF�c��R��!�$���X�I� )�$�
��!�!�Dvwr,�jR'=��i��Oǀ9�!��V�H� �	M�dݺ!)A��/�!�$Ͷd��	B+�,(�t�[���F�'�a|!["� �9(8d����ą��y
� &Dԇ�&{69B�ZR38�E"OԄ�tN�������cY5K��a��"O��:�ə7_���%B� ��T��"OB�(��ׅB�X5�t�����*�"O�B��	����L���R�"O�C�I��|���ŕ+|��'��'"��>y�'AF��XJꔒ>�Ahg&�S�II���OiL�a(�)ry���q�̊q�<a
�'ɶ죓�J� ���RG	e�Z�C
�'�v�Bcʙ�g��q���.�:
�'�07 �r_�qCE�/O�Z���'�`�4�ϩk�nI��֑J�ʤJ�'�Z}��A�9~&N0��
�Y�6q��'�T�h���l��zsHՓdQ8�H>�������Oߨ�ە�ȀV�
�Ӈ�d��a��'/J��7�'D>^�[��R-]ђ�C�'
B�q�F`+I�f.)e�2!P�'k�����*|�8���g�^
���'�!yƩ���e�P��9�''�X��1(0��G�Y��t8�'>z�%)� 1�l�{�d=R�}�������O���>�IP�|��`���-0�hȱ�K7D�����3��`e͹����7�4D�pI��?7dZU�d#
c����M'D��'c��6�t�k����~�~�Df#D��:�%�~��01�7>�j'N"D�ؚ�R9,�¬����8�`Xs�2D�DB�׿�n�d`Q?.�tLs�1D�t8&�[J�xh�,:-P�ؚ/$D���0e�=Jit����7qW �8d-D����
!Kti/�!X�l��+D��cC���&I�ϊ	>���'+D��c�N�Nt�"��]�
���&D�<ЗU7+�j R�D�$�8��#D�8a��99ئ���]�s
넌�ON�$#�)�'62�����o�f`�wdȫ9�����'n���2�-�D��ǎ��~� ���'Vn� a-�;O���2D�
��#�'����y%R�r�����V�<�fb�G'�L�R�M�|N�P�F��G�<�AdJH�̙+D��VD�XJlI@��\�<I�iȵ�L]��kА+�t2t����x��W�S�O�bV��"A���
�i1 �����"O��	���0�d|�E� �j�Q�"O`���`�o���r��ݢ,H��8�"O�劰c�vP�i�Vn��S.P�u"O��S0M��Z����,*D�"O8}q��V$�4O��^	��'�"�����#\hJ��\)r��y�I�O<�D�OR�d�<+O�c��`Ԇǉn�h���_8@ �Y��#D�<�E*G�<�NLP�Q�
Rsc"D� ��L�,�9%h��ʼ��!"D� [�C��uQ~@	�
։.��l2�!D�xʄO�1Y�T��R^Nuz�M,D�|13�Z+u	���i��xDb��(|O���yrO
�YLν�A&i��H�C�W9���hOq����J^ �q����8>�|P"O�q0ƄԬ���d��ĩ�S"OY�&l$:����+����"O�xDD�v�6 ¤�P(��I��"O��)􄑶�����ډ|L�q��"O.IY���,E��6f�'�"0�"(��0|�Ao�8w;��bC㖁[�ɳ�*�q�<��O0&�04����'�o�<� �Q@�۠W�t��ӑ{��%@ "O�ĳ�$�`�|�w�5zj�id"O!ؑ���"�.hJH�v��tA�"O�h�gI��
V1�*�=і%�c"O$�Ʉʜ�u�\�*��m������/�S��_]sʨҠl���r-�B��%!�$�;H&���F!%�8�Q�
�u9!�D�u�R���E	z������L5d�!���! R�Qag��]�L�)]U�!���?,��J�N�-\����F�!�d¦g�T@1�"��:	�mE8$�!�C�.��ᣄ�=^5�6l҃�ў���y��Pyb�ښo�]� lS'�d�O��O8�}��+�J� 5/�)f�h�"g^&�昄�#�L-�d�Or���@�	ͼ�F���U�����ꕊ���/X�n���b�G�<!��P�O��fک	a����C�<�SA��4- �����p!��@E�E�<!��^�Q��SW��@Ul�A�<I��B<h���J���	ȁ�T����'gɧ�i/�	�O�N���)\�B��L+4G[WC�ɪi¨�Bj/t��J�MZ47��B�	?V��c,[����S5a�1KvB�I�;{=� �
S����A��:B�	qPN�G�hHl�e�[kPC�I�� �AG��Nbdz1a�Z6"��$q�$�q�	?j�D�V)(�j9�d�/��4�O���À�?���
��8�AV��G{��)��=֠�R(�?!:L @͞�}��O.��"r���:�`�:H��)a�!�d�M@|�N�+�8r�:R�!�D��H��M��@K�+n�ȊtÔ1�!򤑢D1�l��߂$Z���D�חơ��%���Ac��1~`��n�u�����*�H��%�ިi�x�Č�x�C䉱W�T��s��8~�jV�5y�C䉀;��� ��!Nf���Ob�*C䉡W��%���H�h7ܣ�Eݡ��B�	������_��L]�]�C��h�	�[(6�ty��V%m��C�I8S�ʉ�	G�5�����%^�qhJ��ȓ
K1��L&V�*�"��#\�h��X���xc˨Hd\��WQ��eRdp!L��	�wKHm�U��Z�j8a�PJ� ԡ���~L�-�ȓqj:���N�52�	��ۊ#ǘ��{�yb�� �xX�b� I��o����<�Fꇾm���% �.y���	Q"D�|���V�o��x���].���1b!D��I��JO���!N� �&�f>D��*��	�\���G�g�JQC#)D�P�b�ē�0Lq�"�!�Z|�eL&D��o^�n������� ���/�I�<��aϙj�nH��ƷP�ΤzԪ�D�'Ra��"�RF�$1tL^o�J[�����O�#~BC���@VlĻ炆�'�T����{�<��L�3ytr2VO@!��e�b�<qw��`pԈ���	�ø�Sp��g�<iVo�#\�&��v"L���a�<A%�=OL��@��ŗ2��0�t�^�<���7�&� `MDHY�e��Y�<р��  ܡ��K���V��V�	ٟ���C>A���)]�2b�W`�ajq�3D������0
�p�mI&g�j�Y�L'D�� ���#F� ���S��ؚ�B=R�"O�T��	֒@x9S�g9%�Ty��"Ov�*q�
22|�8�`L4nl�=�"O8�4 M9J䔥j�]�x�8%)"O�i@G]�{�:u�[�O����"Oƴ 䀏��D�H -0i30"OU^'Q
���ǧ�+�n���"OPt��	@49�:U�L� &����"OV�y�cQ>jl�hRR�@ ����"O�9I�E�#�8-����k� �+�"Ol�˙ f{�Q�gL�h���!"O�9����K�<� -A�����"O���ք�,_@08��B��<�1"O�p{��B�]�@���dJ��9G"O��q���#���E��^@ax$"O��Qp��� ��,�u�ɺO>{"O�����]�)���"Fܐy��
�"O2�A�D`�J���"G��X��"O�Ĳ��zĘ}��o��1U(y�"O�=�G�B;ZOR��p��6vG8�82"O�P+5�Q�!OHUJv씓{0 ts�"O�����n�y�R�ǜJ5�G"O�]�ԠM�u#�ċ >R���p"O�MKנ]�/ٚ�hq�@�s=��"O S�@���(	��ܷMʀ!��"O�Lz��&s$�DC1�\�w�&���"O2��P'X#�����<U�6��D"O��[Q��u�f����ͮ<�I��"OD��AO��X�.�1 4p�@à"O`2%�V���DY�9�����"O�{R$ %���C�*.�5C�"O�(Z�gC�Hu֍�ա�:X��`��"O8�Vd�/�����m\i�,�W"OVt1�[T�VQ�*@�k��
R"Oɐ��Tl��JV��`�@�ñ"OZ�b��ٳ�L�yCҷ>t�:�"O�z��̈́S�j@!�>54Q�"O�!H�]0��K��0n��њ5"OܐY�����B�OX�k�ry�"Ovͣ�@ ���œ����"m��a"O��
�����LH��ˣ*W&�(S"O�`��܃L��Ĺ`eǦTV����"O���k�.&����$0����"O���qE��w�x���`�U���;D"O���H��DҠ��ψ�c���a"O\H!�<<p���ytmQP"O~�(r!P��åM�E��u�"ODi�v!�y(r8�u.^��xr4"O~�!D�?|h�v��=0���"O�YÀ$�*p`r���b���:͢�"O A�
�
�f�C���" � �h"Otܺ6��:L�+d"�Q�,�"O�s�^�G��=�V��[��ͱS"Oh��䏁 U��1�`�3�D5r�"Of=ѠU:8,t ��/Z��6�a'"O��1�AQ rP� r%���g?�4�"O>8bql�(j��;��X�p��i��"O� Jd�̼S^�X���{�Ɣ�"OL$"�C)%)J�B�l�b����"O�U�V*	�*=R�ڴFS����w�OS| T�
87�P�C ? 6٣���y��.-��� �!lv�81HN�y���:�Z���P�I����)���)�OX!Ȇb��
�%[E患1]H`�"O� �`��$��eJ���GI���yv"O^�i֋	H�`�s�(�`a�"O�ufGUxl�tS;d)"�Qd"O�Dc�� �c�D����s�@��"O���� �?�b@@Gű�JdR�T�����l;�҃2�x�
�f��D�O�˓�0=Q�پ/ �L�΁$R������}�<�S�.}�<8ptΝk�Q!F�|�<��#�8A��a�� 6-���Aiz�<�`$ڎ)�P�p`�%����O�u�<�#���Y\�X��`Z$��aQ���wh<�UO�u(��@BޓQ��-Ё,��?9.O��d_�lì��u��%J ��'I�K��'a|B	�,�f���*���r�'�-�y$_�T�A��Ą ;����¡�yrP.1`��h�*ht8� ��yB�T�?x)x�P?�Da@��y"3sJ�@�ꘜ~`��X�$,�y���-�D�QiR9+	�$�U�� ��$"�Ox@�sb��
�b���5����U"Oȧa޴Y�h8$ �m�����"O�ͫ��� �p�+��ʂ�2 "�"O�\K��E.[� pV��/]���Y"O�*�1�| ����w�;Q"O��Zr�\58��D���["O�Tr k�0���d#�P*���D��r��W�D ��dY^Ȩ6lW�<@��	���y"�?/���G�5"�0�v��3�y�'�pN	鐌C�&i�ƌR��yr���h���}9�3��y��JpI��Bi������y��N�˂m�Cڀ��q�1�yr��W�L,s�F*!x��pjS���'@ў���<U-҆F�ЫVa΄���*ZI�<Qu�ہ��N%m�r�{�f�n�<q���i�f�ŖXJ�-��g�<��×�@N�ۢ���9����a�<�`g�Dv�}�ݐw�I�ƌr��G���O��:1)ǉGK��CѢ]O�(��'i�,
�[��	���0�DBJ>���?����O�+'Jl�*DM� �l	�y�,	��Ӑh�7{P�aW�D��y�ɜ��Ʃ��k5B��q��*�yB�i�bY�uk� q��Z%��y�� �P���ŏe���0
�y��H���	��Z �tH@���y��"'	(A�!ْT� X!�D���d�Ox�=�|��X�aA���
\�S/歙 ��y��[$���J�XO�B�7�6�y"���id���I\�5�G�ѽ�y¥Bd4��pK�E��Ɂǉ���y� �6+�f%�s`��<�*����y⤔�q�@�:7N�5D����]��䓖?���d/d���!'���P �&
��yBJH0�f��f��CWi��!�y�W*M9�a��dƼ9O�}��ȝ��y��[���#J�+�@�`�(�y���S!����R�/�>��n��yb�؎t2�q�M�.��Xib+���?��'j�x9c��n\<t�R�V�P��	�',ք��h��Hn�{"��T	t-�'$��+��O
q�NLQb��/L>J�k�'��t��cY7|���P2�H�R��I�'_t�������za�۶I`l�
��� |hpu�MQ���+
[�B���O��A��
�v���mu�J�)D�l������}xg�S����)*(D�h�����r�^`h�H�=�Sc2�����H�-J8���`��m� �D"OF4B"έiӨ�Jr �2V���"Odc�4
����c�ɑe;l��S"O�t���[�=
��x/�'$��ag"O��I���)������l��r�'�!�D�D����$˸j�(����l�!��8d<�  ��E	�-ۆ�Ώ+>�W�l�<A��@�O6e�UbSj � Z�aSo�z	�'���SQ 
�c�|�!�ށ;��Q;	�'cBEJ�	��|8q��£1#���'r6�1�]% ���	�Ro@� �'\�����yY�i�AĜ�^IT�.O���ě���U)��D.�9RU�J�7*!�d���0t�b��6U��� ���Q���|2�'���'����+ϾjO����I
gT�x��V�s�!�DY�-x\�h�{M�IiE�K?D�!�ă]L���G���fV��
+K�!�ňx�D��@�/DV��p�ʆ�!�N�
X���mF�O�4�x�4>p!�Y�?T6���iC'{Ji#tEF!;[!�$��O9�����7M�������!�dH�u��tphыn��ʵ[��'�ў��<Y�ęݚ\+PLːq8�HтD�R�<Ń�-:�!Kg'D#�i�!b�e�<)���ez���Ӭ��' b!��'�K�<���r�)5犊;�,��DB�F�<yr���U��4JE)�^��E	Wx�<i�=a�y��a��V��c��L�<�u 
V����7)�/� Ȑ�!d��hO�'Q�pB�PixR��jɅ�%��ܚ6�(�h�)��I�̇ȓZ-�ip�7p��E�>/C*(�ȓ���.L�o�����H�d��ȓeR�1�͉/N)IWf�7��9��h<w�Dl�FT�F���H�$��X�<��NĲ)���u��l�WeT��hO�}���i�Ò(7>
�����(�Մ����4K�*O�]:!E���Q��N��i!3�V��8�{fjͿz���bs��$ݚi�f�W���_��Ą�$l��cb��fՠ�HFMV�@0����M���١��&b���� �Z�-Ɩ �ȓ�)�H�-q<q���ɔ��?Y��0|Z⛫K�C�`@66Խ�hVJ�<��	AR�ƴb�L�)0�.�j\�H�ȓ�&maሓz���g��̇ȓ`�`�B��z����$^ �ć�D	:\ui�O�$��I" ֬��l�p��&H 7�"$��d]�z^��ȓ[�&���9mT�Q�j�0 *e���D�r�W�-�J];��24=�h���JH#���.XG:-+���Ht<�ȓg��ly�F7(���!�ARօ��=v��ב"P�$ �/Ԡ]�F̈́�RF��@������ �Y3NEv�d9��3�U)d�H�KԩJ')�����*+D� ��$����I��SԠ��0�'D�Pj0��_���k&oRz9�؈`	 D�ԃ� �j��ӵ��;��t�C�	 �����*ε��/$z��C�)� l��gՠN�fYH���R�UP^���	v��Vn_!{T��G�]�h�Z�$;D������)�B��`��Ӥf<D�(�`H�	$4�1d!� /��,�B�9D�@��MǲVb!�r�O�u�<ZP#$D���DÃ&o��,�6�?+��܃5h!D���q��,&���QTa�0/�,i�� D�lh��ˣX�!�ɟ�,����1k�<q��$-4I:��/�!�b��S�	>`�0`��B<�'�� ���	 �6(���{���F�<��̝g,�ъ���x�@�k�.\�<�L�3`�l4�p"�3[n`[�IZW�<�gδ1����B_LR���,H�<��F�k|J��f)L�p��EC�<��;�}�U��L���kv/[gx���'et%��f�$�L��"Fԋpb�)[�'r8`�(՗�x-�2�К��� �'X�)SD�2�Z�*� h,Y�'hD�ń�	p4�(�U���d�'nf�x��<���!w��~ٶ��'Z�p[�h�3N��uZ�͗*y��)�'2�8���0I"��
�/C�Z!�
�'�H����# ��IHj�	*�ܹ	�'s���pcY�gV�8b�It��I�
�'����nY1GT"3	�%�0̙�'<n��B܇ϸђeM?~�q�'��x��"'.�����ԃ;^���'����S��F�� Y� i���
�'�
̸$%�NB��C���d�,�
�'��VB�2x�[�h@�h����	�'�p�tąD_(�)C	�6wX0�'V�d��BN�rM�AbT�G6�;��O�x��&@22�dT�T�:It��"O�Y�Fو�~mK�B�LNP��"O��$Ȱd�V�S��N�8��"O��'ڥP|.�ZGI�|68@�"O<�˦`_8'�!3�'0l.�E��Op�XĝcC� �$/A�j�0�ˀ�<D�H�fn�:O,#1ɀ�c^:�z��<D��7�&�9C&b@�Q�$	�ǌ<D�ܣcˏ%{=<]�!K�%��Ѧ;D�0���2X� �b�<3�AE=D�3(I6^��	���(^��� =D���$!]�k��qC,��k�|L��9D���5�p|�s�öd1F�9�),D�h��͙)g/��Ȧ���Dr�@�58D�T���c9hI�K��1��i���8D�`�w��/Iz`*S�P�&�~��F:D�h;1�@���
v�M%CT��#�<D���c* q|�xRF�E��� F�O���O���<�O�"���Q慵z/���I�'x:��!D�А�	<<p$�O�4��p�!D��B�Hm��% t�#��#�B>D�dl	���q��-_!?Ej\ئ�:D��낭ޞQ�`��D[����B�=D��r.R�8
�xa��.n�H���/D�Xi%)N��!S�P>d_�y���O���O`�O�3�	$r$�sD��
xN9qr�� ��B�?u�f��G&��/�*a!i����B�ɄMے�b%$8��Y�1L�C�	;G���Թ2�|)Q�!ǖC�IJ��X��Ķb�Ј8&� "6�B�	�D�P�:Nf�ɦ��
�$B��8T'�(�ELw7x�: ��8!$ʓ�?�����S�π �2�NA$tP�h>}B�|�)�b�f����J��l)ˆ ��wy0C�.5�T˂�
/4L2Q�T&	"F"�B�	i|���֟j��p W"M�=C�ɰi���di2fH��3Eŏ/8K0C�I�uH��C�E�c��)E+ C�	%3V���k�]u\"�)�, C�I�
Vq{��O�`�B|0d�3���O �=�}�	Fk�e����R�{ch	N�<���ޟ=�@����Z�>��aj^�<��!��Hp W~�v=���X�<�IǠU���V�Բ3X�:���I�<��-f^���3��D������D�<���z���ѵc�O��Q���e�<!�B�{�tY`�@�cB��!6G�c�<��'E#K�z$�vdԭQɶ�*r�^T�<�r��j'`�v�S�@��bAƜX��n���OAd�� o�B��S�n��\b�
�'�����A�2%���P��4i�N�z	�'�Z�Ru�lf!���)A��Y
�'V�Q�&#á/�01@�@��8�Vq��',XL�C����	V�в7� M>����I0wL�� U�N�
�Ą�å]&+�!�Ӄ M�\@ �ʵ]�b���	X�	�!��A��$/) ���[�!�F�:_t1
$�KO�AzGV�!�D�h@�(a%ċF7b���eW|�!�Ɠr��P���܆u�4��ھX�!��x���D��N��D�h ���	P��(����3��%Pta)V���|Vy0B"OTd���p(��jӈÈq���{�"O E�_4.Y*}���S�S֛~�<ٓ�;n��1�Z�+�&�b�<Id�+m�Ti`�+%���%*�T�<q4�W�������5�2}���	V�<f'�Zqx@ PB�SD�d����N�<y�l�.a?h����$���J�<�q-ԣ�<�b�I�tH
my��J�<�ѫS Ijlq���\��pk�F�<a6f�?Kh:��r��>^0Xa ��l�<���_�
�t�P�W&$!!3��<��B Y��<���<5^�\"'@���lG{��ԑ�x��O�KlB�ku!ۿ|�LE�3�8D���Fc�V��`�K��O{&��sO:D�YF#7ypD��@��&h��+Շ$D�X���Q/FE��F�/1�$�v�#D�� ��^�ϐ����	k���ie	#D�(S���-A�=�j��fJ���B,D�(�kF�E�t�pf8M���0F�O��D<�i>�DxBe_�dޘxP���R%�(�AQ6�y���<�=J#n�P�|�R&�)�y"	L�()V�����Q�"�_��yR��>�l�f�A�w�8!ׁ.�y"G��x���h�-L�zO�[d,�y��\�)��(x'#pg�}��L��yrb��hq6P�c�g��͚�	��$9�S����lp��W� ��yCB�e@p�0��$D����b͋h˾�	����g2Ae�$D�`��H� @��h�I�T���hև$D�Q3�>I�$�R��<'>��'�#D��0dH��Cj�5�r������7B6D�HV.��hĴ�"%f�e�<���&D�h"�ԣ#�e��ҕR�Q+�-�O�=ͧ�O�m����H�r)[��H�6��1a"O� �R�%D�*�Dɱ�D0�>up���Ɵ�D�d)�*V,@9�R��D�� B�Ý�y�`\XK����5l����&V(�yB
�$�5id�������D��y�g�1����'`5�@�4	��y��"=��*"$��[�^5��ӆ�y�IN�V5���'`�(n���i���y��U]6�����"Vn(�镏��O
���O�b>�b�ψe��td�@:�Hi	O)D��P�ԵWp�e�J_�`�8�!��3D� �����.�2�Պ[�E���rm,D�P�r#�=>`��Q�m�Eܸ��J,D�b��YJF���ϗ X�r��&6<OZ#<y�Rf�H�⯒(l�p�F Dj�<�"�īWN�!"�H� TP��X��f�<�m�:zN$,�E�YO>\uKr��c�<	�È�=T8���ƗiZ:���a�<	�	��D���7�ߏG������G�<�-������v��a����F~�<i�Cߟ(���F�%w�!#�@�G�'�1OV����#�z܊�(�`	�pJ"O��%�=bl�� ��t!�̃�"O�)A�O�
k+P	y4/�".�,1�"O��: $���H,R�CD:�|���"O�9�Db��c匄9�(��'�DP�G"Ot)ffE>G� �ӤgN�0J a�"O&D��)bV࠘�Ɩ	6AS�"O�q� .�4�EB^�1�2"O@����0-���
0��K�<�"O���b4^J�<3uH\�+6�l2Q"O �АB��Od9+��4��"OV%x��Ҩ:�,�&g�
l� I�"O����kJ�8��f.T���P"O�,�7�B�#��a�!�� |BV$q �'*��R�nF�f���a@�:�d��&D��HbLM�A�\$)$��S͎ [vf/D���'��/(�p���Od����.D�@�q�ŬUA�i���L	�v� �.D�T��G�&��:�eJ�4��{�+*D�HCQĄm��Q茴:��ܒ�*O"H��,ąV�0H�Q�2�X"O�%� �����fI���"O ẗ�OײhC�e�l�DX�1"Od��A�L�X8��s�S���k "O�8s�G�SՄqa�cL�XE�"OhI�4� B�0��B$T�6�!�"O
	��NH�N�y{��C#:�<\+�"Od$���tEV��/"�R%p�"O B�_J�x!��I��:"O��
3	ډ7&@����-�ni2`"OT�GlV;\��)���@�:=�R"O�,�� �l�Q��p�Pc"OD����U�j.V���k�?r4��"O�4����  Ѱv��f�W"Oz�ό8�T\�D�+GL�z6"O:(�rثm� �x�&�r7vh
�"ON-�QAϖ*9�p��%��KQ
��"O$)2�Z�-W���*�<s18��"O��"P��'b��1�''�N!>���"Oz�b�½F'�Y�#G�;9���$"O�T�����?;,�Xg&�)_6��u"OvPx�&�,�6�A�� -,wB�"O�����ւ
�T eP:5WzQɣ"Ot媃I
V�x�	�*���"O� ���dm�x��@3cU�~zFm�"O�( ���?
����"a]�Kv�ç"O�m�L#
��` j=Ҍ��"O��8̊2��#�/0=��"OIpg��آX0T(_�S*p�+�"OP�{!���"z�E��>"��V"Ol�+��ɎWD8�.>k�E�B"OB9h#��	t�՛��LR5���"O����nɼ*�rp�"�AZ"O.ɰ��V�k�4R�*L\(�٨�"O2PY �U�C��D���&"x��"O�z����6�cB�L�!
�"O�9��d
�Ȁ5F� &���)�"O��"VɎ�K�.�Ӥ�$����2"O�P��&S��$Hj�V����D"O	 D��M�]�T��L�
y�r"O�Xc�K��c6<c�n	!*%�B�"O�@�C
�s����Q+g����7"O������x	�aY')I ��!�"O��+M;H�4��6n����"O"�IˀK��Ie��^,R�"ON�d�4D옽�"��q�P�jF"Or�-F۞�YŦ�� ��y�"O ��^/aa�5�gе��eQD"ON�2� ��C-�pЁvsZ�P"Oz{el\�Ai�����a��)p6"O����6̨\��Z�#�d�Jq"O�P��J�=r�d�`�ꀡSy�H�"O���S��63��P�J��Py�4��"O��X��ɰm�<���Y�$rri�"O��2�,4G?�t�4�L�_���$"O USv'�W�J0��Y"�Ȅ�G"O�S�	�	 \�h���_����"O�m&NF2⪐ѥ�ߟY��[�"O��r7�I�)�.M���/;����`"Ovr��&��l)4�Z����"O�!���Os`�
�$H�r� "O��1A���X}�f�S!mHĻ%"O��tLB�'�~�S3��=T��"OxԁM�Ơ����jɪF���y�E���(�A�	.�X��gO�y��H	w*� �ۡ�Rh�v�]��yb*YR��ш]��:� ���yr��=.��s��P!�L`2Fm��y"��'#� l 1��u!ȵ	V<�y���(|)�! ��n��2�G��y2[�(|�����T�~��4c��ە�y��ѝX����{�Ԡ��C#�y�ܧEF��C F� �6�j�k��y���tSҘ��KM�	1bi�,��y�$�Yh�|���Ơގ�BTD֍�y��Ȋ$p,��G�C���dA(�y���Z2z�@J�?����� �yB���
% ȱ9x���n�,�yB(�"3e*9`F�Ҳf*6r�$�
�'��j�f�g*�Z�G�N�d�;
�'4��P*ڊp�v�+��<J֑
�'9蘁fh�	V��	c���A��

�';�P��+g�*��=:�*�'�re��
��y�U�T��F�x�'��(P�ʁ)�v!�P%�o�����'$�)�#`� .����A��Vi�t�'����$�]GR�p��;�^1c�'2�S�c	�T9��@S�S�
L����� H�eP�$X��@�:��"O^�:���J$R�dZ�I�\��"O������~*�:���T�ѥ"O��#bp���ă:u⮨[�"O�e��������c� �x�"O����ʽpM`H������|t�U"O|}�oϿ*��T�AN��IR��7"O�4j:f�P��@7Ny�u"O�$��Ɔ(�HX+�$��v$°!�"O��(���+���&�G�v�Q��"O�-`u%F7;6�X�$�E19��"O��`�g[`������l��M�D"O��r��I3m���ӅC(cO��!D"O��2���+u �+��ֿ�2Ds�"O���-�&u/�p��ԏH�l
"O��A�*M�j��s��5D䠻�"Oʅ�g+'�J��)�a���v"O }�F\'B+�Ś���#$~ެ;""O6�[�)��59<lk�%.nl(J�"O�-��m%Y�2 ��zU�� R�<���c���*r�8evP�NU�<I�aȍ��B�rkb��@��,n!�Xi�����!l�hIDI�al!�$I�@���X�l�ee��y_!�d��N4:'Nt�d�ԙ U!򤚧/�-�d�F79**4�3���=!�ў!g����o����'x-!�$Nj��Dcf�:e���2bԲRp!��|S��
f#��y��1	��ш�!��?c,M�������Nҷ �!�dP� ᚄ�5�[�A�>{�K;D!�d���|����L��t�l�0!�d��tn����x(r�+wJ��u�!�ů\
�̀@�S�+���I���i�!�D��u^�	ʥ��+(��X�>�!��&12hy�8r�
������!�d�(Hv�C��9�FP���pw!�D iY.���KW4Y�d{E��hr!��J-��h�i�*u�+r�[�)�!��(^2E˥)]�	���8����!��(�$
��X#2��X�d�T�B�!�$��4���
^ $l0C�7|a!�d�����Qi�s|���"S�}C!�	@��ȳ!��F���u�ؗ�!�d�c�@�S�N�x�ZL)�h05�!�6&L8,kQ�ȝ|��U	w)��h�!�D޼l�6p:c�'t*MJ�jX�]�!��]""7�����<>b6ذ�҈d�!�$V��:��$���˕,]:H�!��˔y�mi���FYn8aUe�Qv!�$�3|�~����{W����d9@!�]�6=���כC@�H�d�2!���0��AL�m��Q��͞�!��[)+��0P�d�2�9�6O'�!�$\�r\�wc�)2u���`_,�!�D��eL�D�b�\�'q���ñ+�!�$ .6z�֨]�s�b�(R�3M�!��@��qǄ?-��F��7k!򤟚}�@tj!EOr�pe�	V!�d�l,��%쐁u(�K'W�N!�D�1i�^�'�9p��Yh�.d!���<�~%�� Z�F�I� Gɕ7Y!�ĕ�N�&����^�]���k=i�!�Ā+�p4y�b�;S����[,6!�� P�Y'mT�(i�A4�z�J�"O0�A���	N*��R��U��x�R"O~(M[*�<1���q�(-R�"On���t!���cf	`�4i��"O`$	'HT#����֡w���r"O
dzA�J�^�,x1��i��"O0ȓ完>"�JP�*��Es"OB���I#V^�(i��sG�� �"O��St$�P�F����2a,f+1"O���b�N�V��(xq�ϊf%~4�F"O�	��L"&NJ(�O4��{6"OX8��FK�6��9���+�P8�"O|i��ª.=`4�F�;�$��#"OLI{�H�����̕ �$��"O�|$�S"~5*=	�`:�Ġ��"O��Ӏ�
<�tM����(��"O���B>#.�=��#�1�:��"O�}h%�ȍ5L<"C��3
�>��"O@���N[�b�x��#B�rހ����'8�O�-h�-��iP�p�q�M�H��|:a?O����	 90f����0@+V�[�@n���Lb�	�`,��ʈ�aC���5.� .�FB�ɴ@}�,[�	^,sp
4�m� |��B�	�<�pX@����?��!k�oI�-��B�:+"�Ђ�F1&��A�afB�]w(C�ɏpV��[E�HA�0�����j*�B�	�k���A@˞�P#�۴_�0��ʓ�0?A���=��A�E_��S�b�n�<��T���r���7�H�@��f�<!�E4v�,����'��ᒄ��e?����$ɧB�h[�蓧(���� ֱB�!�D��00zehT)�!7�h��*��,��"=��9Oٚr(�l���#6h��*>	�"O��f �f@չC�ԃ�
<"O\qR�@��L�ڷ`�:q��Is���	:�~,z�Z�ؑ�k�<�!�$��L�`�e�	�1�ށ{�*��!�տR0SU��<f�F�P�K�!��Ŭt<��T"B� �Q�D�0�!���V�����k�3St�ur7J4z>!�$בO<-���2Y����Ѫ�2
,���Os������/ 14&�2��C�"�p��āʡ�yrlH�Z�0H�Q
�H����`���-�Oɒ�e�(<=�p���$
0�t"O�d'�v`�8�f��$��ʗ"O`,Q�M� ŀŢ�11� �5O@� ��Ʌhry+�N�xR�ݐ&(5D>LB�	�?(���c�~�9�([��C�ɐtlI�Q@�$4�������"EsB��.XT<U2�'��9�j�P���eb(B䉆#͠�ݜ��˅��}F�܇�I*!�h�S	�L�x�
����C��+ �$�@����>�1!�e�7հC䉔��	��
<iv�P:g	���2B�I�<.��d���z�+�]��➜F{J~*��S53N��3���HP��+NT�<��JШ\:�L� G��>�pI�1B�L�'_ay"O�$���P�U�P�N��M��ԟ0"<��fX�=px��䆥f�6��-�G�<fj�xjZ�csڜS�|����E}�]�4G{J|�r6��z��s=�h�r@Zz�'�?iW
	�hԔk1.M9cZ�	�:��W����.K�*y!�f@�S-87��<\��hOQ>]�F�ݹ ���*۝A��X��3D�� ���0�ӵ��h*��vc�]��"OA���\�.��� ��F���"O�@����5\?J,�2�]�&E �b"O���B㍏=N,y� �.Y�XXS�'kqO�0�˖�v
+7��Tb�	ޟ�E�ī�*���	paQ	��y �����y�u�䒐�ε8��Dk?�y2�{�-����o�%Y��M���$�)�>��M��[��̹f�L�U�6I�$oGUx���'
�%8��Z�"�|󗨃+Yy~Y��'D���d��, ��H��1W�@I�	�'��(�%�v#>�Sqf�<@�y���hO���U��bH4�cϏ0hV�{�"O�[�"|�rd�� TK�B�"O`��-N�~�E0�y1!w"O�(�Uh�;-i�D�aW�wwt��'��e��a��@�:�)12m�=������?�w&�)�N��T|0��YT��P8��Ez"��Xy�{ѯ�8*��c�!&�0<q���U�dG���fcH!u*�a ��E�>z��hO���f�6;��*���i`"O��+u�[�T̮��m�.M�� "O
d(�����Q�U�P42��S"O��J7$��J�$�9H�w~���"Or�S�aʌ
;��	F���7����"Oh\��Ç/5240��!�17��×"ODx��эM}J��AI�έ�"O~��uM�\����4��MXq"OP����8 �&�8��� '�8�"O��q2�Q� (���ֵX$\�A1�;\O$�(pa^�f&���G��*'������v�<	��������:�����v�<yt�	(bsL!p&�'{�V�[��o�dF{�N#	��Pգ�9B?�8���Y ��'Zў��<+h�^�����u&�	�5"O�M�QM]�n��)I�L7^#^@�v"O����'	�x�"6�ߥ;�d�K�y~��'R�ギۣ.��$�i�\հ�'��}p@��44ޅu�T%	m�<�'�^I���1�5�kW�S��y
�'��mc!�ˮ$JX�`k�
?y�{	�'��A�#�PdE�)�U������'�^qScB-$�.����ƴ:��H<����!���J�
j����fi��u��^O�H�� Y��H��D�nnB�ɉ6��iG'r�0A�f撕&��܄ȓG����M/��]���Զ~���ȓ6�,�pqE��0���6G����'��Ey��	Ρ!*���խM�L�2�k�<�O�%C/�s_��*�KKuBʝ��dk�0�=9�5�d�-p��Q�ŚnL���ÇH��d?�O �3 ��&���OB4kV�1��O�����7 �!��W��dE��C��O�!�$:M��-#���pӖ�a&�(�!��ߖA�B��w�ɢ<������f�a{����5V8Qx�F�f����Sx�!�d�Xk AX��� ��HK��I��O�=%>��4nǡoÜ�S g�9_���p��)D�<����Q��`�B��B��%D��3!,O�~�d�kM/b�-�gB$D��+�ѹCd4���P�a�t,��'}b�)��"u�|�[ �J�[��Ī�5}9)�����O�I��Z�����L=b��\��"O  ʷ m�$���`��E�>=j�"O� �Г�T�Y���[�J6z� �"O:$�u�/[Ƣ��+[�J�"O���`��.o�6���k�I��qR�"Ol�8��~��y�!��4���ʔ"O E�w��eL� �g�r2�"O�CbBN�M\R O�6if�=y�"O��&ÞH �@�2BrB� w"Oּ�SbԮK��P$%	�WZ���'��$��PAH�jԮ�i�d0�����	p}���S�JH~��G�\�p(j��P/G�n��"?Q��	�L��-�d�;k,2I�f�{X!�D)h=x!�.Z��|��]�!��q��(�4��g+�
K���R�3u>iD"O��@�K�=s�ۀ%�����d7�O03�K�)�����ΥxK6\��'�L�����`��`�BI� a��1�/1D�XA`(�06�4�agF8?�TI��3D�� b-�����3t'E.`��	P�&1D���hЪ�i �$|����$�,D���r��X�b�Ӄ��Y@� D��{elBTp���.u����3|O�c�d�A�H;�(Q��?b��*�l,D�x:r��s�:�Ɂꓝ\�t�#�=D���N�V������S�!�8��:D�|�s.C�	Ϧ���O����
%h$D�|�Uj����O��$�O#D���P�E��,bEm��X���(&�<D��93N�,]�g��d|b"�:D�<I&�J�WX4��%~D�s��8D�t����#�`"�O�n��Ak�,#D��C�K�c����bd߈\��%���4D�\0��%u��=b%�G,��c��2D�ċ"�ɻ\�X�uG�;,|�2f;D� 0Ag6��q�d焠(C$�"O:D��'��Z�e=V���Տ4D���4�K���)Sn�=��i�N1D�l�%O�?jV�O\���Q
f%1D��y�=�z����� ��g2D��#��LO��sw�W1	^(�a �0D�XIed��m:��R�{��Ab2D����'X�
���a�;v�d�(�.D��1�e�>l��2͵r�����,D�����li�����"2��,.tbC�	*�M��M��V:Bi � ��>C��c2ʵh�.�*LXޭ�tM�N�C�I�9�"����M���)�7�ܬ��B�I5J�K���6$��ڢN�u#�B�	n��}3&�P-Fe�PX`�؝��C�	1S�}u�_<q�}B$K.3��C䉃a�����g
)�e��ܜw{B�	c�Z�bTИ8�j0�#�)��C�	(hՊTA�&ۛ4��U7:��C�I�N�^%�2+�G��P+r/� hB�I5+��q�sMH,9�u�IӁI�BB�	�]�AK�*פ{R�CE�L����:&�Z�F
�nn�B��ƿq7�8���@5m2ȈrěJ�!�dԖh>,����,+/n�� iAc�!�bK6Mf�4]�A�P�!�$[&7���¤W9k��%�c�GQ|!�$W�+�X<�g�R�*g���W>Z�'����/9�i��䌆_�Fh+�'�NdP��҉q��-�a���U�z��	�'WT�Q�xlܠ�Т�}6�E��'��xfh�!��`�E�ԘC(u@��� ��
f9�
����͝Q�%Y�"OV�eoɯ
��u�Q��}Ӽ���"OV}A�B�I���K�oO����"O���A�]�|K
U��(U j��=�5"O�)@��v���G��x�"Oz��pbY���Tŀ$pi`"O� ��^,S� [ ��![st���"O�<���sy�X@p�
3p���W"OҼ3b�|����,L
�,��"O�]�^�0�h�C_�e#^��G� �y�H(���#��U$ĄK d���yR��<�� g�	7�j�d�ҩ�yR�AN�"X��L<y�|B�M���y�LC~	�m�V�I�"���`$���y�����	���58,X ����y��-��iج
�4��4hY7�yB*՗}Y��A�3R�𓭔�y��EP�P)i$�M�5�h)�b����y��V�4m��d��9z{����K$�y�I��
�(��-b���yc�5�y�&V�	�p��1j� Y�́�7�yr�ƤR֖!ۧ��?S]�xd"J�y��KF|(��G�_;E��OO�yR/�,��#��I�B���x��ˋ�y�gW+�h���YF���A�ʤ�y"��*m�V1ʧ�*�������yb)M�z��V
Kx�zw,	��y2$��e�d���`��E������9�y"b4j��4�蕶KR�TQꂢ�y�f�!U����ŧۡi*0x�hA�y!¿V� abY�{f�( $��y�C�:�� B ��{�t���	��y��X<�v�2+�%Z���Ar�-�yBG�6iX0ȶ���[e��&A��y" �*�����CRTjZfɇ��y�+w�$2�+�K�����y�		�x�Ȝ��CƚA� ]��^:�yRrW�0����=G�@���Z��y"�Wa��92��A�?Ǣ��R��y"
�2<�*T�2��5˲��y�
�6n��r�֯_�h�yr-�y��
^���/R��C��Q��y��Ԫv*�D '�E9v�����y2#�9Pv��dR�O�$���*��y�k�(�q�V w�MЁ ��y�V�aQv��a(�/=�`+mȢ�yҫn0��〆X>8�8�-
��y��G6HT�3��TIV�ҠBJ#�y��ȵ�q�e&ז+2p�V�y��Z�=F�����;�� � a��y��#>��PCAk�]q��z�GD��y�K^�vxbD��ń�#*���N,�ybď�a��)�e�9nP��2'��y�DF�~��r+��d��8�j@��yr�E�D
���ń�"���!I)�y2��*X�<��k�_w�@����y"�ն{tpB�P���Y�,Q��yFG��J\KC��!@[.���Kޢ�y�nW7v�0�+�N�!G����F���yb�����"���~��"���y�bC5ݞ�+2�^&N04��ڄ�y���!U����W$��N��̩!��)�y�D�22xp�5�Y6qk���n��yB���1��N�i��ޒ�p=����s�)��h�� ���%I"�Nz���<4�0�I"O���#L�؈�Q�+���
������*��c<��}���	����Ξ�yW�@a�F�<9�(�z)иKd+	��~ �
 �����ͺE��� =.^�?�'[����.o�ђ�e�Ƣe��'W�a�eΖH<؈1&�W�*�����bV�D�d�g�p݄�I�!�,�H��(��Bv��m��󄁩��"�m�k�aB蒠Ts�a�a
�4�JaQ��47��B�	%,���0`�k�~8��#%��Oz  pG� #�l��K�2e��uC�/c ^T8�C=ٰ��$�j�<Iwf���Hh�����5�*]�5��rk�(��E�j>�\HC�R5Z~���O�h�gFӓb�L��Z;n��O��HVgn� ���,e���E��9:������p��ܯ^�|��Č �عqt-�o4`(�����1�牵!�͸���'I��R��D.�έ�'[q[�0�)�	ɂyؗO0x���ݾ$��4��J�Ș%�$O�ܸu�C&���B+�C�X���d�T,��<�W˟U�44��1��q��YX�8P�g��E�h �H�U�!�EEM�7z2�F���7��4����<n���8����|m!�X�I�|7m��q�-p�\sU�I�?<�	r�P.rgay���,s�<�����X�HP9��>��и/���Ԛ-S-BP(�$ڦL��.��yLC�I|$<�����<��K���K�D���CZ�'�Dd`��	'Dx�Z(A��T"Hˤp���:�3��'��U٢��i��5oE�v�rsl(����]��	�z��s��p�h<���x���'LU�2�O��qY+����O�ƽS5�P+��Ȑ�"�9ˊI��O$ձqI�q ���D�8��$M��f��sR�;ʌ�(Ac܋��OJF�0���6ݑ5OH�7	T��"�(70@ߧ7�B��+4a���V[b�:�>p� j�&�*m���!���K��'o����KZa�<ҧ�T�>�f��qK�	��xh�N	���<�V�/�7�Q;$#L��t��6��$ X(#z)��� !r�He�K��C��RRG�#��)�'<�8ȳլ�U2��d%]�l$}�K>�T���m&y��=Y�RhHCL�˘O�"�j7�[��BD%��0��êO���G��-]���'�IzdE�j��1&��(@a��P$FRN|��۝Ae4����O�vXYpJy�0!����ʺ���$�?��"i#=n!�$I�����$�;x�y��V����9H����oQ6.�s5AȚ�����zy".UƼ۰�Ԩ-�j�S���K�(�ʤ�B��t�
R�Omp�0�)rvjV�5qĔ��+��G��d�0#`�``�(
��ɝ_��Q��I�**� �b۪fI��j�`P�K-B�25	�	y]F(�f�4V˘Ћ����̈�tIG ��p��4��J�'�~�ȸUʴ����<�E	ѝ;�`��B�q���߷]���!C_�3�<`�ߐ?�u�}��/��ɚԨN+X� %c-��V�����/`JpC䉂ztb0�͙�rat�P�t�J9�GGցA݌Ma@�F@�A'˔�p=(��8}���#�P�.�Z�*�[ :#
���GͶ%a{RD�tR���v��">Q!k�BM�����Z�����02,Ԍ�P�ڜb"�'e\�)�A6��Ol�2M^��49��⌅z�=����@gʼ�a�I�~'ZP�dB�1�O�r�""O��s�`	��f�B�
�[�OV��W�P�5yj��d�.`� ��E�����'ҔG�����&�9�F�8��|z*Ay��Ϥ(�DE�ݴ/�%��F�>(�Ha�@ jTDĆȓ?t°A`��+oi�P*��_3d�s'�cV��6��D�y�&к���(F��(�P>0w$�
5dʍ�a{�N�P��l�`ղT�p-�׊��6d��0I�p��V�� ������'U�D�e$�m�(uK�?	Ŧ��,O����O ���2|1�Z*BFтM|ʥ,Ρ
�~Q�mG�l`$��-fX�@�G���N���D�B+_2F�~�p���)r �@���D�>��#�떎t��:'B��h��d�9o �L�Sd!o�`�rW�ˀ(���Hɔ��E�>��f�ԁm<����G�x~�ӧ)̟�Ao�r�� �<���D�mX�D4�`T�[��"cי�M��I�"���M &��/1B��!!��=v���a��&d��3��:,/�Jt����
���4mD��L����[�A�8O��p��Y��![4!��O�nih3�K	w��|�!�/3tU��Zh��v��O�B�Dϑ]S68`V�[�aゔY�'L��C�g'��O?5�'&\l*��� �z�fl�G�'z�Ѣ�3� ��i��J>�(4�t�̹M���rq�>a6�s�b��d�- S�-`��� ,�*%�!�d�%=DZ��R�]�T�Ib�H�>�!�#LǼ�(ǆ��;�t�&H3i@!�$��}�8�b'K�P]���Gj!�$�80��(��ܙ]��%��c�*1T�'��5����i��@1��D�z�d��"�4I!��_�p<���Ֆk
M�'���U7���1�+����c��u��mL/&�\܋g�C	[���ēfڬ �6�C�}4�M�NG�/J��v�˲l�8��d� FEfᄢv�x]�#Cېayb,�B��&�,�2�`�n8�G�
&�!dI?D��鳠Ȫ_�1"&�W�4 ��k1�$��Q&|r�{��D��5q�dIvLX_ሑ��J]���O�Tc!g*�'#�r%Ò�8$̍�Lݰo�� �{��6G�zb?Oj�"e�>8z��2�@�M͚��7O$���G.���h�� �����U�P��U�E�&��D2�˲hLC�ɿd�0t9��ۈf�
���T�q�t�ʢ9�M$\OT��u� 3-,���NB
+y^`!�'+�<r��+"pl�Q���]�M��Ҷ,#^���'����-%�V���?-�4	�����0{߀Ġ��)�p���T �7}}�Y�Ú!D!�D�'�̽x��И.2v��eT�DI�
T� ���{���P"|���Ӈ ׁ�xB�C��@l!�䐳d�N�H�&.�|�P�1)P�M_.H�
�xd�ia"��J��ؕi�3��U��8���r��N�Y>����&��xɄȓSˀ����U�%V~8Z��Q����ȓb�A� ٱ�4�$oM�"F1�ȓ#�tʦ�U���z����yr��7L6J��1��M���	G���yB�Ü%����窞(Ct ᵢ��y�'�2�����I[�9�,�kE
כ�y�k3G�ܰ#��2�*�%���yb��h��Q)ɡH�eQ�4�y"�ئA:&�Z��� (��|���G��y�λ_GH�H�*ɖ&2��b�^��y���y�2�B&H�#fE4�eӱ�y�i֣D��� �b;������y2���х���7b��z����yj���ȓW������7Sl����H%�&M�ȓ%>��Ȱ�#H�\P3� 1�!�ȓX�V$�doɭ�8sWE��b$����(�Q�/��:��>~�H�ȓ_�*���c��]�L�bGU9Oj���7>��'���`h�lZ�LKz!,���/��4&Րj}�D���� �����x�A��.]@>�B��\�
�ȓ_;����x�E�a���6����/jB䐴MʂA)*1§hǤ_�Tt��K��أ�jP�V�"QX5��.xԨ��z0P2�ՓW��Ux��[�� ȅ�l�p\��JS�C&N �Q �܅ȓM�I����/��'��V�b��S�\� �(�
=A�xBR͚���x��h�x�A�dٙeX4��C1}���S]�f`���A#u&�(tֺ�ȓY�x��jU=*׺��Fb�(To�h�ȓ���1��Z�R�k#�M�`�,Ň��*�9��4`���"����P'����c44�P#�_��@z�*/}S�!�ȓ!�P4sd�Ȓ��%�É3AzU��E8�(��	!t�@T#d�z���ȓHEj��'J^�#�B��UE�?�ń�S�? vE@!n�^��-���+��lS�"O�P���C0P�)xeL�M���"O��ѧJ�#D����²+9�\#"O���v�"2t�P�b�2,>qh�"O��B�o�UX�Xg���WN��"O�k��M�`deXS��:��Е"O��,E/X�����gX���{�"O
���!{֩b3�"yƅ��"O���k�<;8j�0�c�I�ك�"OX��&)�:���q◆\�Ɂ"O84	��9��ܩ��\}�U�7"O&��cJE�W��)E�6IT�1Q'"O���Ơ��<<��J�4 O�"O�lA���~3l� �KV�1,�|�"O���z���!	C,#���
D"O���;0�X"����є"O8�0��8$�} ��^	'��	�b"O�PA�K--�4I9���/�84I"O&,Bwo�r	<@xb�/`�4*O\�C�ٷX�4�J��� {�ޕ��'z"! ��#����P�T`'ر��'��#�j�y=�ب4��0XF΀��'�bB��:����#�T+��]*�'V�L�5��!A���j�#n�9��'>Z���I1C�,�[!�j��<r�'�p����+|�*<���>P�|��'֌ ���)X���%D&D@T��'�9�V� 3��s 'V#'��
�']pq�@j�����2Z6-��'�:��v���b�@-�fk��)T��B�'�0��d�4��y��͍;Qƪ���'��m��)@w%x�`^'N�	�'�n बؾ?,q�����݀I	�'��방"�&ɲG����z	�'r�D�'A�;�L��@����	�'�=��c_"D>2,��/�\���'����,��u10�)􏃕_���'�n�
��W5MV�e�C�C�T��L(	�'� [WŞ�UMH@�S)\*v�S
�'Ln�v#. ���&�.r��z
�'슱[�MT�G�5��n���bi��'kB4b`�#$�\ �PJ�P�'4 ���VT��m1Vm ���'R��g*LZeTE�����A��'�",�Q"��X�[*K�V�D��'L�,h��ɮZX������
O�!�'�D!�l��� ?�A��'��a+�� IaL�ZM�6��' FlcD��!��1Q��D�9����'Xx�Qġ�*����@@��3Q
��'[2���ًRb�|؇�U�{1ZU��'����&�2S.
=�F�ο	����'Kx	�W�!W(���"C	���
�'游�u��-R[NP�U&�U�Z�	�'�)0ugY,�ܡ`�52FZY�	�'=�1PġD}�d�V#��.�E	�'倭1Q�1-��T[���Vx$��'_���S�$Ԇ���� xj�5:�'�sq��d`Ip�!��Ȫ�'��!��"R>Ei)0���.N����'��Hu.�"@�� '���@I�'8��`�����W�EM�C�'T�z�D�e�X�9L�&O�fm��'���+J	 ���hňMnA���� fC� M�RA� �tջ���"O*٠��{�8 Z��e� � �"O����;�����C�0}A"O*���D�#T��MQ��@��y@g�'RС00�<h�]Γ!��x�1� �f�\�@� H8NI��Ͷ���L� g�Fs�9g_v��<	S���eZ~�ـ�˸�h��H�rm"X�"C��L���"O�+�f��r`�D�t�ܰX�lep�Q�Ah�UWfd?�F�����	)FĹ��*���$����bC�	8`�ٚp&ߩ;��%P"!�3#� �"�m�m��J�'a{B(�80��q3��5�>h�u���<!�I�7�&@����1���C��
4�q�L�p�T �u���y�'^�-�����#����MH��"����'�i{t�����==񟪀@�OӌD�b!�B�4�Z���"O�����/̼@B��	8�.��A�>SR0��"
'!����O����&��ņTc0c�bT9|�tهƓ8j�8���R�(<
2o�'b#�k�ƈ�8��ayE�á%�2\vB1,O$��LD�&����h8�-f�/��<��eL
k?�5!-q�x)S&�YSI������*d;��3�i�d��C�ɛ)ϖ����W� (���	:�c�8�dS4>���R�X�-QrAQ���(G�j�X��+LRYH��D�yb"���U��;SL�S4&Z�P$�Q�a_�21�c��O����Y�|aӍ�*3lR}:�C,&M�L4K0D�(!dF��"���ju# LN�X,�<�&kՏbL	�"-,O�ؓ�K��K�Θ� �\���`%�'���PU�K<*�&%H��G�Y����_��R!BH<�2�d��5���6�6�x&�G�'�E0Ɯ-8���҇+8�d�h���|'�\@"Oʱ{a�K�vLA�غu�j��O�T:�#�����h���c0�eݘ���߁cc�؀"Oj\�i3[j�u��-O"[������R @���	������	�0z����̯�����L/��Ma�H��2�H
�#$=hU��
��ٳ	�'���0�I�;%�-���$�FIZ��$��&"�R)N��O�U�ː8G�c ��$�b�'C�J��YSP���P�ʩ9r͓eߒ=P�eʘ�ҧ���]$n8 ��Cq�A.xP���)<D���SB
�vM��n
����0�>a�-�4q_.�����EX����*#4e����ڶR�ȥI�B9�OH}��c~��2��-}��e�fg
�m5d�Ƌ�:h]C�	�޺�a���~��BD-��~~b�<����Ԯ�1G ���O{�؈���k�
�5�[,^�����'a��Q�!�_sT�T�<" �&��F:��g�R�B�S��?��
�kl��2eF'EP�lX���i�<�Q �tl�Q����A �40&�c?qso.
%:Q��qx�d�D6v�(	YP+��_��	9f'2�Ozaʇd��N�y1�Sd�5�w�]/5&� r���y��K�F�2��`�ӗw^���.ڼ�(O��+E�ʹC�>�È��R߰ՒD��8���,�C�!�$û��b׈ޫ-�aa�	�:2�+AiQ�u��ʒ�>E���8מ�B�T+T��D2��I/���ȓ$�0e�!n@G��0�P �8	�2��'&(�$����zr�F<��%���ϬC��-��M����>���
Un6M��A.��Sm�I�T)�*¶P�!��QKeĭ!�0��O�FL��'����M�o&��;���?�Y��'���� 97����0��
�'>�!4*�5F���biRd�����'x�qi6��`�$���O�Jm���'w|�[sӘJ/\�w��<��	�'�<�P�U�=�� i�36"�z	�'�ZpP$��1EP�@ՂW�~����'*<`��_
�0NC�m����'��t��`�- 2B�(1���oÐ!I��� D�31d�U�H�t�3�Zx�"O	��c
l��b�C�%��)R"OX����%��;�cPR�΄�"O�5q��L+~.`!pAEN��3W"O�dxDdأ ��h�A\�b�ĲT"O�d@�3L� xh���4����"O���F��B�ԂQM�+U9H���"OpI0ף��î`/A�P��-	�y"撟/��(f'Wbk������$�y��\.%]�%+T�]�I�Ej؃�y�],=נ���J��P
bYô!A0�y«��\,N}(S�D1B�bq�k#�y�oN�\@�f.�'NN������y�Lâ|^���f�3D��0���.�y򇝐?���(ҭ�?�t��ɂ�y�>')�4�F����K�ƙ��y"�ȒKI��xu&�I���l[��ybN��}jt��e ��B��8;wGD��y�Ӫyx��&T82`�l�y"�T qY� �)$-,��E%J�y��K�:���V�$Լ���!-�yr��?!��+�fD�
K�ؘe����y���n�݊��ăxق����3�yR#�	I9��)A��n��_/�y��<���.@�ʺ-!v���y��߄Q��� UZ���M��y���i�ȭ� ��G��5	E���y��h�|���g��8��෨��y2�V�p�ڑ�d˔� >D!����y�O�C��s�	�i`�ۖ���y����q_��R!I�!n%���h��yB�H�B�����"b��h�R��y2��3>�ȹ!�l�u锑k3�܇�y$��)z�q�"�O92"Ή�b��yB
BQ�=SE*ǔY�&hPRB ��y�F�}׊�pwf��V����&ㆴ�y��Q�4�� ���D���Z�o�3�yb�T4�y�DU�L䘀��'�	�y2,I�-�Pċ���?�lh� ��yҏ� g��P�$`������y���wT<�Ǩ[�}vɺ�eA��y� T�$[�	ԗ	7���Hߗ�y��T�Wl޴Zj@�YFZA�E�A��y� u�h ���Z�c�FD��3�y����������^��ˣ���y����Ȅ�,�� X�9C���yReE�JHb,�1��q�����K��yBJ�;N<`E�q�*zcEʓ㙶�y�Jק$Ǵ���ڂp�8 � �y�!��+_�P�hpY`F�y���R�3� ^�AI�x�7�.�yR`A,s?>@�0��6l�H�i�-��yR��F���,V�o�F蜆�y��Ɣ�i!C�(B�r��W��y�k� BRC�``���"+N��y"@�)8H�򲅘�nT�k��P*�y�cN3��=ʂ��q�D�%�T��y�$�\�����	�*>V�9%E<�yBb�v������bt�s%�C��yRGɁJ��`�߾d��(at$��y2%��D�t��A�_����8�y�1;8ԙ��oG�Vi��P.���y�EIP�.�P2l�8u�$b�\4�0=a�d�=Jp��[�(EܼjqnȒmkmjƮЀ����_�<� �,zƃ��!$�!A�Ƌu�Rܺ$"Obm!Ǌ-7�H$�ΗW�t2c"Oƙ���<�h�ul&~*�	R"Oj��a�v�t�_�:�	�S"O����Ct�$��J�!�2��#"O��0�!J�s���!�I��p"O��bg�T
܈�CU)���$�IV"O�Z��K�[��H�T(砱��"O
��[!(C���GK�W@lI��"O\P�VN� 1Fr!�)K)>,�5#2"O�@T�
�;_�Ƞ��,����"OS�U�]���W
�#�2W"O�@G���rP�Y���<�&�(��'y�ov��#�N[��|k�*�>bT@�v'Y�1�y��	 2gh>E3���2����[C�${�����	78���'>�ю��oO'fg2�� �ua ���g�|��pjfá�y&�-~|$������tM�oB�%�B �e7flZ�醓A�vM��O�,�!C��O6���S;'�a��E=l�6�J1��p[��,�e���
Q�
�ӂ�O~��H0/��ۖ�Ue8	�ڴQ�����r�Py+O�?M����`:�9��h�(N�HՉ�4z�=	��ڃ{��IO�3}�O ���m�?]�.�[V�%<�$ �ڴ��"~n����)V�Ixb�Y�bP�vtB䉤h�\���'b!h̹"FʲW�dB�I��� aˆ�m0��p	ǅ][LB䉸^g��8f �A�e��X�B�B�ɏA;��3�&�?hV��g�T��B䉸��q%�;o����7-�$u�C�ɰ
q\(Z�V1kq��B�N�K�C��R���g�NGJ@	%E��B��=s2�a��0
��"�9���d�0E\��J�uK���A�P/!�$]}Y��1щ{8�x@��֒r,!�DB�~�|���&E�,���nZ�e�!�$',��XyFȝ�1�CI�3U!��"g&�jA�֟@x�6��"�!���>x���[@�{Q�y�`C�W�!�4�"�UgE�[GV!QP�O�!�=K�����ӑ�
��p��~�!�d]=2@[�#� #��=k@�GB�!�$� |�>��/������&  s!��%
Ĺ��͂�p�z�J��C�!�C,dM���TKA23ؔ5�bCE�!�$+�����X��YDb��!�d�_�tc������%1!
e�!���~����ıB��壳���!�d�64z|jQA�bk$�YC�Ӌ9���B'Q�hP7O:2r*!r����y��܊1䶜��E[>zP�*�]�y2$�>@���wB�mO�ـ�$Ĭ�yrGX()\�Ճ��űX�D�³a��y��ӎF���yՀ*J��G�!�d��Xy��a[ ��[V�\	!�Ė�n�~!{B	�p�b�î$!�DE<L�P��ȝ!d�|D�1@.N�!�%k$�$Śx�t��;�!��W&k�^|;��P	R�ToV�g�!��˔] ��·K�X��Ō:�!��73��\����/�ީ��AU�`�!�$\)bd��0��T��#oYZK!�4 ��u*�&_�r��l�����U�!��B�7��2:� }@e��8vx!��C�ql�m*H�rc�Qc*C�w���߳Lx*=Ȑ��pF�C䉋w+6m8��D'vh̼jPd�5� C�)� �X��$�"n��4�b�1D����"OBy���N���z�aF0C32��"O4��&hҹ2�n8� ?w���5"OL�CW��n���k�H]�~e֍"O�I�&��� �v�ʜ>�\��"Ov��*��������`q S"Ox�0�7lA����1H��"O��Z��?jHa��nB�w20XK�"O20�c_�i��`Rl<>%ve�F"O@-PF�ԯ$�2�2�֤
#"�83"O8�� ��M�<�)D	M"-
�Ͳ"OR��u%A���80�G�-�ވ�"O��2eD�r�>T����-Aߌtx"OpU�n�4;E̬ڀ�X�!�܍��"O&� f1:�b�2%L	-�|�C�"Ol���,�2�*Q�����d��"O���������Re�ċq��M�s"O*�0�LY�X�(@e�`u�I�"O`�cׅ܍�}�s��q�=��"O�����V��>���B�l,D��"O��獊+{P�Ӧ�>i��*B"O(���4`�������n�Y�"OH�Sd�yL	����:���"OVb�H֪r��43���}߼x#"Oy�bM�@�p�"Z�X�v	�"O��Z� ��}J������.���2"O6T9a'��|.�jA/V'Eb�=�2"On����&sn�rX��&�*8!��i� I`6���0¦�B�%W!�$M%h1Jq�@>��`dU3Z7!�ā�d�{� '��5����P!�ҍ:�rPK#n�@"diAR�2�!��,�fQ`r��z�����ӏ]�!�$��i>0!3��������b�<]�!�d�>>�P�q�g	�a�P�YToc�!�lm@䀃 ��.W�Ԋ'A̚S�!�d]+"�H*X�:6R�JB�pd!�DXH�t0!�c#څˠ ��Rg!��p��f�v}0t�5�E�,\!����D����.\�N�{���B�!�@T(N����w�Xġ�-�<x!��_�h�X����P�3	.)M!��V��-�w�
0$=dXa���W"!��Ұ=c�� W�Ǻ%�J���",!��B&n�F]w��+�p!܃j!��ܢ:`Zq�C)�<P:�S��ԞY�!�0�nq	����HO���S R#�!�ē�R�4����Fi(�zV��2'�!�[�<e�h2�N�EOj3��!��<+ v�{8���
��Ql!�
a�ص�B"�T��5���ɞ&W!�2}:`�IqL�({���P�J�q7!�ޝ*#`L�whM,A�P��Ş}�!򤏒b����AS�d���r�!���&���R"��M)��X6B!�&+z�Z%$Cb������/!�$F/&|�}��yD�q�֥�j3!򤛞Bp��+E�z�]�^d)!�d�9ij�
Ad2l�
vI�X!�ě�TV�ݹQ��,�$\+�!�i!���I�64s��W�w�n�JC� )!�d��8E@0��~x�ٲ�+D�(�!��(-B|@�!��%��8s*V�A�!�߷[��@��p�8��L�!�� ĳ�EG� Z�����Pz��"OMr���0�,�r瀗EJ�<"Ob��RB��q�$�Y�/LP2DH"O����O��p #�oϏc��{ "O&0���ܟm]��ڶ��V�Xqʁ"O�Ӧ��~�F� �'^�v�G"O�Ԡ1-P�������q�>��"O��+e���maZ�Q呰J�Ti��"O-¡��i�}�vF��5�<��V"On�@aU�9���ӄY n��v"O�R�(�Sx� ��i�S�>Ԙ1"O��wOt���P�iqv(($"O2�j2)Y%H2q�);v� "	�'GT\�ԭ�&�Yt� /4��3�'����a'G<t�q�c���0&�Y�'��r���'��"	2Y�X��'��5��I�5�땟�(���'{r�jӆ�,b�j�) �N�|�F�
�'c2�;�/]��&ɀ�![��:��	�'��ZC	!K?�����61$U1	�'����C�7����N��~�\�	�'v�(���D8�kw	\o�H��'� H��g�^X��+ס�i�"Ȑ�'-B%	S�j62R�e̷w�~!r�'p&���M�?n��DY%%�~�
�'~|2��$E(�d���4��9�
�'����L�HV��C�D�'�����'�~���M�������('�Ɛ��'H�]�D�hrT��5*���'4�A��@rꀕ�Ԅ��>�Ԙ1
�'l6<Ұ�
v�Y{�;Z|��	�'�&;p�V��T*��.��s	�'
-���1=F�J�NG�~4MQ�'��L�#n�Y����k�^@(�'���"�C.J�Y���b����'�^T#ҩ�����놁�b�aq�'J�`�W��W9f����T5B�
�'rYE ^���G_�LE���'���C	K8_���)���Ah���'�������[�td��儙8��I�'$p��)�i�N�P!��Q`���'��3��T�V��mZeƝ0rx�h�'�*�i��̮""rŹ�ꙟ ���'�V<��W+�����b	r�'�̛b��]v>�(��S��PMh�'d, qnٺP*�'��&�6q��'8Ԉ����O
���v�X�d����'S��W�W*u�X�z����.u��'|��K���1k�H-z^nl��'{Q�ơ%!6�ȹ�쌮n��y��',J�1v����AQ�X�P�'Q����$5V��S��񈉹�'�hh�CLB1z}���S���+�'9f$b�4G$���Hx,s
�'Ø�[s��r`�����*��1��'�L��N�z^��A0,�Ԝ,��'�<z�.Q?ꉢw-M�!����'9�K�LW;c�%��A
���0�'�h)9�X/)�>	³Ëa"h��'�\�'�T"C;�D�2	�U	��	�'��H��[/ Ѱ񚵈�:R����'���2�̰:B����	¯A��y"����&�24F#���&�y2ǎ=;2Aq�6z|9���y
� �}�����Q���̵s�%a�"OV�k�F	�B�ZP!�Tx0"O���/���2	R�e4"3���"O�xy�Hޘ�d�F��`$�r&"O��
��a�W$
(�(` "OrY���Ln��)�@�[�:��m{�"Ot���J&���#���R����"O���w*�6��,����, 
��"OL��a��� ���[�
�-��"O�AaR�D@�ࠧI�[ҭZ�"O�A$%,z�՛�e��I�"O$]��o
v��3����6���T"O�(�PdՈ�4��e��o�8i�"O�k�S"	�
	5�H�"��Mx`"O�A��ɂ��e� \+][n��"O��N�0^�����nBVa��"Op��ᤏ�<T�F& �I/��2�"OPpQ櫃�O X�6�
/)b��"Ob�"� G�x�t��&��j��p�"OޔA����eV�򲥖�N(�"O,��v��;�P05� <�N��"Oh q�kO
L��T�W=o�T�"O�4q���9N�[���B"Of8��g�����âҨs��=B�"O�}PcMȾ2aP��٨Z
���"O`؂'"�5m9��� ��� ]X�"O^<���*��!��/R:<�ic"O��)D�1RT��ƠR�0r"OHD�   ��   �  ?  �  �  �)  5  L@  UK  jV  b  dm  �x  ��  ��  ̏  ��  �  ?�  ��  ϯ  �  ��  !�  ��  ��  �  �  ��  ]�  ��  ��  9�  � �	  W �! ( e/ b8 �> <E |K �Q /R  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+!��6*\�c�<4�d5h��'�B�'���'	�'/�'�B�'���U�W9��m��Ʊz�0�b��'���'�2�'��'�b�'�r�'���k��.Kªa��͎ 5���Ha�' ��'���'�R�'���'���'����
F	�>]�&ΏfEP$�b�'�b�'��'�B�'�B�'O��'�$��zm@|XpjC�6�D�'��'���'v��'�'��'�"1�)ֽⲵpa����j5�'���'���'t"�'��'��'�%؇�Δ*��� A�B4%
0��'�R�'��'o"�'�"�'/"�'�f}�b���Xs���]��X��'iR�'���'���'��'W"�'g�=��'��"��	�Jw���'���'j"���d�'5r�'}��'��u�1� (iL�\r6e �t|:\���'�'H��'J��'ZR�'vr�':h(uC�=��)��G-P�����'��'u��'}��'���'u�'�;+�'HhufUmzn��`�'���'|��'���'��'p��'�J���R�h�����*|h�p�'���'��'���'h2�h�x��O��"�q�R��t�T�)����G$�|y�'��)�3?E�i)�ZT��}G��E�ɢf��<G�)�'�63�i>�IΟP��fL��,2�j�>LX]�� ՟�����Z�]E���Tn����O6�,�3�=��)DK�I�T�J�yR�'��D�Ob^�'(P�,Þx���BxHl8c}Ӥa��d,���M�;(��j�L�'���	�"� w�8�����?њ'.�)�S'���o�<�C];�NŊ4��6L��g�G�<��'�*����hO�i�O,���=pUl���*П��ik 0O����F��f��֘'p�Y��n	�G�PSuj�p�̒��\}��'Q";O���\�s�(�����ڢG�_c&�'��\��H�����VßL�v�'8�	��b�8�tKS�ćc$��K�S��'%��9O��"��8Q�D|
��N�5�`Ab@5O��n�/Dz���V�4������ňY��L��j�0�1 4O����On��;�6�=?ٝOx���?_$��)S�Y�;� �E�]/_�z��M>�-O�I�O����O^�$�OАqU���R����G 9?E����<a5�i���!B�'x�'��Oy��Ql>^p�1(�%O�!��H�AZ��?y����Ş(�@C�.YX�!#�gʼ�p�MK�_��8S�{��d6���<tg�?^:u�"I@  � ��TI���?A���?����?�'��d���\��
�O�|��F̵`�f��p�B�!�\�u;OYo�N�7��Iݟ��	ԟl���w��m�t*�8~��1���
&�Umx~�DX?c�p�nܧR�B�=������_���S���<���?���?a���?9��4�
5?�I��H�����cR�'��`Ө]��3�����]'���W��s/�$iA�v_��Pm@N�	����i>�I��զm�u��+�,4�!O�;�y
l�/<��@�'��<%���'N��'���'��9�@�|�.�k�n�9��	�D�'8R[����4z2����?���I�caPA/�8@qI1��}��I�����O4��1��?9���x�P�i�7��Y�Ѭ�,���s'&��]*?ͧv�������Hxt��B��p,�qٳG�����?���?��S�'��DϦ=�T
Qw���#:�U��^�3W4�KtU�Xߴ��'6�듛?I$&���	'�X�2r̹P���?����� ڴ���.z���'����iJ�pt+�/R����Ӊ�����IyR�'�'�'bS>Y��	-v��R��%[��S`	��Mc�Ǝ��?����?�J~�p{��w%� �6�Y?D�L���
�\��p�V�'��|���h�>D��<O���'/� �;���L� |�"6O�a��m;�~�|�X���Ʉ�	�`�rB�^�4�ԟh�	П@��Wy��o�@��b�O����O�(v�U]@�Hs&���R�!�!�I�����OB��%��p���a�W�qt��rUl�"*�ɯ��a2��5Nvb>�ir�'Dv��I<~�Q���m�Œ��N_��H�i�mޟ���͟�F�T�'U��1�\4F��8�N�Bo�]Ғ�'XD7��>:��˓ZZ��4�$�/U�t�0�0��ֲ(x��r5OR��O~�$��tP6�=?�t���i	?(��I��E�Du��%M+�D�J>�*O���O���O��d�O���f��W@�f�֔a�������<�G�i��l���'���'��O��nD�.]ԺC�&�rȰu���Dꓸ?i����S�'PTz�)��0)��q��_}�00�-�@�M�'�0a��[� �6�|�X�H�߱wb�9�EB� l���Yğ��	ן��I���`y�h��M��,�O��2GcK��>�Ƀ�ޕv\>�p$��M���i�O���'���'[�Y�kۈ����[8�`�F� #�|׿i��I#�<�c��Ojq���� �58��1pt�!��ӌ"�(K�0Oz�D�O���O��$�O��?mK�������Q� �4@I'�������(�4D�Ҕ�'�?i2�i7�'gV\�S�Q��<�#��Bx��|Z�M��|�Ah]&�MS�O̬ȁ�5hrN�hEbO�@z6�i�/ЂB'`U��'z�'��i>��I���I
jf�Q��Ǉ'���"�@]
t�v��Iԟ�'{X7-�����D�Od��|���)> &��7�U���St"�u~�A�>Q���?�K>�O'�z�!\�BL�E�(f��Ѐf����P�i��i>�*�O��O���f�0lT����-�^��#��Oj���OP�$�O1��˓B��&�W0+b��"`�eА
����'/vӢ�D��O����Aݚ��7�L.Yπ�[0��'h����O0��7M6?��W���� ��˓KJ��sb�:-kLLs�(S	N�,\͓����OZ�D�O����O<�$�|J���I9(:��t��t �Аm|���VB���'H����'��6=���$N&-��!Ā^1 ����OT��1��0\7-~�$r�bLRp���ǄE�!6R��mn�` c��|H��?�d�<����?��n�����$	B��yP���?y��?������1����矤��ϟ�SE!F��郁�E<�CKS��7y�	�����X�	7`(8]��eƾ]��)&+� ,n�|��K���TX4��|Ⱜ�O ����"JJ}gn���މ�	ԘW%b��?��?1���h�������p���{j��� $���D�ڦYp�kMRy�gӶ��1[F{�Β�DP��!���|���џ8��ޟ�P���q�'x��#�%�?1i�_'l��@F�++x������'}�i>��I̟��I���ɔBѮ]��xH��ǜJ)>�'h7�$>����O���(���OJ�[�C\0>pM:�(ç3�;�X{}��'��O1�4$:�)G�x=�I"M�J�Hš��Ar
�ZԈ�<!���@���Q�������P��U�71��QAAH�9V^�$�O6�D�O��4���h7��J݃+l2�\"��f�F-Y�0����yb��a�O�5�'v��'!���W�bX��
�Q�Dh���9H�b��ֺi��I;{� i���O�'?1�];ɲu���ފv��U�DD��v���	�D�	џ��	ܟ���N�'X�D�Q�ON�qڡ�2,Ǭ����?Q�����W#����'��6-!�dY�?d��rE��`L1Ӆ�;��O����O��9Iz7�??Q�&
+F�xæÙ�z���#gi�>	�Q�r����'�d���$�'��'u�a��1@�=i�kWqh�Y��'��U�� ܴ9F����?����򉗠�n\���"+��*���.6�������Ox�d&��?5R����q��q鐥�J�`�1u��#UkD9�i�S���|:bn�O��I>��� (eˑ�^����+5#H8�?)���?1��?�|�(O$`m�Sν)��Y"�&�H�^j�Gsl��'i�6� �I"���O��'hCMmL)j��]�.�>,i�h�O&���z˸7M7?�ІV�T�\�>�b�͹Be��R��v9���e���'r�'���'���'D�ylЀ��I�be!��=�@��4l�2����?�����<y���yWΉ'y@�^�D�����*�E��'tɧ�Oʎ�鷹i �F�(���N��	���P�BԊU��Ā(1���� ,F�O��|��K��r����OҼ1Jý^t�b���?i���?I-O��oZ�:����럜�ɗt�^�
ΔI�N�3�- c�6u�?�w\����|�*���V�����-r�Oخ����' R[4��:w$P�	���������	Q�'<�B��?C��zT(�'��+��'�2�'���'�>��	�B\�����E�cT�Zgc��O��Q�ɍ�M˶�� �?9�<��V�4�
yԩ��[M��Ke��|pB�2O:���O����nKb7�1?AƠO7�����z�@�0磓dRT�¡Hۤo�<�'�Ė'�R�']��'���'C�x��!�3�rA��!ͭ`���#EQ����4
�K,O(�d>�S*ZH��{vdR�b�̄�TXE�H%��O2�$�O��O1�le�P+�{CB(���[|�^l�"��JsH7M*?q��%�,�	H�IRyRnمk���{�۠Xe*E���X �b�'�2�'A�O��I��Mː�K �?�9_n��q����O:�y"�k�⟈��O��d�O���0L���Ə�%�I`$�4�Rh������|Ҵ|[L�?&?e��PԺ	��)=-�,��a��.1������ ����I���Io�'Xa�9ic�	�U!L��h��*@���?1�� ϛ� Z�����'K@6�)���Tb�)2.�5:�XjՎ�3^Bz�O����O��Рv��6m%?��y�Q4��7v@���D��6?2(�qfÙ�?1$#��<���?����?y�%Ӻ�(��	�Ij�<@WB��?����DWئqĥ�vy��'��S���|��#�<D TQ���� �F�	�����$�IW�)��+���z5�źB�:��*[{�`� �K�L�k.O�)�?a��0��2+)���ˮ��1�倎���d�O����OL��)�<1Ÿi�r�3���,O5��R"�zc,գ�gǭs��I2�MC��"�>���XV��nZ2n2�a񲬇�]Z����?��Ś�M��O���ٌ��I?� Τ[�#�6_�L	"��[B)�YR>O���?i��?Y���?����i�S��0@�l�JK"���!��Bmp���ş4���s���������_?0�`�FV9J4$(5�3�?����S�'~�&]�ܴ�y�/�	��=Sr�pČm�b�y�L�>%:q�IQ,�'�i>�I�Sްaa�N')~��$˒��N9��ԟ(��ΟȔ'�6M]��p��O��dҀPLl��#m���(�:AN�=3�*�ȹ�O��d�O8�OX�v�W~\L��/D�?t������@�_�� :Ta%��>��aE� ���K	���^�iw�%H�L�ޟ�I�d��ΟPE���'l\�%.�7i�A�wA�o��u�'��6�י\�&�F���4�p4�Q�Q�x�𮔌*լXX9O���<AG� 0�M#�OH�S���Q�P�N��e�t.�����:�F��,՞�O���?����?i��?��n�&X5jC  "�@�����Ad��S,O$�mZ7>lf��⟬��Q��=���X 1����˦"l,ڤQ���W�S�'/�x� 7��
V4�d8�"-���aᖙn�d� /O�����?���5�$�<�d-T�� [�a�o�����?q���?q���?ͧ���U����Z�g��5��)���L =%�s"�ៈR�4��'B���?I���?�PD�Uf�SW*|���E�l����4��d�#�t��'��OU��VB �y�H�7q��k��J�y�'���'�R�'9b�)	~[�����@�'��c�2$��D�O�F��m���DRyrw�t�O��oH:OH��أ��_^Q5k0���O��4����{���Eu����.W
}�j}P�S�6���k�%?�t��J��^y�O_��'IBBŭ~B�����h)���T�B9R�'�I��M�����?1���?q,�f����Q�8�j<�儮	L8���Ts�O�d&�)��L	]�e��V<Atr���Ꮵ;�� !uA�4Z�d�S.O�iU��?�n0�$U|�F��U���V��X� �F�5, ��O*���O����<��i@|� �&�7O-D(�T�X�1��ckm��'�J7- �I����O��s��Lls�ȐEH(�(�r�@�<��Մ�MS�O�q7'	������<	�M��2�VyIp����#)�<1+O�d�O��D�Ot�d�O��'=�.p��(�Y+�m���8e�h)B��'�}����?1�����<QA��y7�۝f�C�'�'���@��3
�b�'~ɧ�O�P���i��3a����(6�d�H�_���9�d�'I�'�	ҟD�I5lz�%C'2�&���Hz���ϟ��IԟD�'l�6��c�����O����5P��7&�jQ�%e� jn⟌�O��Oz�O�i�a�4P+��`�N/�xi����r��X�ld�r3�SX��S��p��O_7<�|� 	%����ٟ������	ğ�E��w����\8R:���#�*j�ȀS�'8D7M�?x�d�O�o�L�Ӽ����>���B$L�B�U�����<����?i�:�dm�ܴ����~�:p*�O7�8+�DԹ��DR ���ǖM��Gy�Or�'K��'cM�^�TܷB�P����I���M�W�4�?���?aJ~
��G=:��Dæ\���e�-n�L�{�S�d��Οx'�b>���d&3��pK�m��ݠda�Llu3��IByR��k�~�,8J>A+O 	Ӷ�,z�.��A�8h�Tl����O
�D�O~���O�	�<iw�i��t�W�'o�����J(R�BE �IG:PLX)��'0�6M3�	4����OX���O6t��"�X_T�XC$T������}s��4����~�p��O��O�bM6T2���
^]B�1T�ަ�yR�'�B�']�'MR�I	(pX��1*U#:%HѠ@MT�E�����OD��ܦICM>��I�M�O>��`�">L�
v�B	$I���e�9���?���|ꢄ�,�M��O61�5�ך�b��i�;	B��i���(J�b���'��'��i>5�Iџ����d�iW�3n(��3�Q������֟��'7�6��а���O��Ĭ|�3AW�8�b��㝸L�Չ�%AW~2,�>����?�K>�Og�<�p�Ϲtᆵs�iڕ-��4;bfN�6 ���i��i>m�0�O6�Ox�6 �b٠���Ⱥ9><�0��O@���Op���O1���7��6�˲�RB!���f�:4;��N�'N@��'cr�cӰ�\�O���9�pQC 8��	�3Y�'����OB��jp��F�Py`.�S�mp�T��P0	l�e�)�;X���Ey��'�b�'X"�'��[>9w�ޞ}��$�	�WX����ل�M�#�?���?A��t�j��.D��U�������@4k���O��O1�~ȣ�z��I�6?�QP��N�'�P�bK�y�B�Ie���rB�O��O|��|���g�dI�/�`������0QD\
���?q���?y)O.�n��$���˟4��e��2S��S^]��G�>����?i�W�`�	ڟ|&�B��?�{�!N���l9?a��E�9`~U�i�v̧>av�$�6�?Q��n4�iѧ�T�v�b=�scߧ�?9���?���?���9�5 q�R��\`���	}�H���O�EmZ1�4��':6�8�iޕ���%�d��j�[f&�y������p�ɆO��o�u~�)Y���� ~�V�Y�l+h�
��J�W�N����7��<�'�?��?���?q�!^@�(i��݆>������XͦM9��؟l���x&?i�I��`,�wɎ�l��z��X�-<��Ol���O�O1�@Ղ��ϔZ���(#�ސ:��mZ�	�)�b6M8?�����`:���\��qy�,ӽb��[��]a0���)���'���'i�O.�I��M�DJۊ�?iPK�+��Icȝ�9 �(B�c��?�U�ia�O���'���'����,"PD�#m��l�`ɓ0b�����in��$O���P�O[�h&?��ݞ,6$�ɂ5VDL���92��	��IП �Iڟ��	Z�'JՊ���G\�k���	�I�0٘����?���{+��e ����M�O>AB��-B�,x�	�
d�!B�:���?���|�s���Mk�O�(u�K7]�TE�7O];'Ĩp��`7nۖp����֓O���|z��?���k��z$�C�~QX�rp��&��8���?�-O<��	 �l�D�O�$�|�����k_�e#f��TjLq~��>����?iH>�O�d`ĩ_�y���U UP�: �4�AFH�= �(\���4���S����O0���HK�q(jxHc��_������O��D�Oh�D�O1�P�e�FdD(+C���ӂDF��P$��5L���',"``�`⟈�O���.L�r��p�ܹ%�x8	V�ҌyQ�$�O
p�m���wdYg)�S#hZ4�+�����مL>a��xyr�'�2�'�b�'>b[>Q��T`U,�X@��:D1�WΘ��M��/ť��$�O8�?�����uG_�j.Z�Ar��������?����ŞS��={ߴ�y"�W�y�ū �C:]]��Q����y��Ъ
C<��	��'F����ɽ"�>��g��� ��N
4�����	ޟ��'�p7M�y�����O����NAL���>�\|��a3
"J�lh�OL��<�I�k�~�)d��(C�Ԥ�A��`C*�Q�4�a����g���N~��O���sV��ϋ�5��M�Ҧ�vz�ai��?���?9��h�������@�$�b��b'���nm�Ŧ�قK�ByRFn�L�权 ��B�,C8��h�G�~Ԟ�Iܟ���ʟ���֦e�u'B����
�Q"����i��l����-�E&�`�'���'�'W��'���ծ��sW*�0����zEn�s�Z��޴_ ��*O��$*�i�O<��Kt�������zv�X}�'@��|���DE(@.��G�B��,��G[4h��c	5�MS�Z�8ڢE��O��<�d�<�E��IL L�s`�<q�ꀄ��?9���?����?ͧ��D�֦�Q��ܟPȰ��/.�d�2�܈A�,��e�L��4��'����?Y��?&��l9&�*2�On��A����6�y�4����z�����̸O�����\z���-�*Z"�]Á���y��'���'�2�'Or���iVJ�jE�4�ȴ��$�	�����O2��Gʦ��u>�����M�I>I&�V}��,�P)%!��xdB�����?��|�!H\�M+�O���Ԥͅ4�ݹ�Oގ�����]�XP�'��'b�i>��I՟L�I9T3��
Aɛ�	q������d��hyR~ӠECsM�OD���O˧,v�a�hN�OU��9��E��<�'���?����S��F~rq��쓜&J�ږ��;<�`<�w' h��ƕ��t�d"�D	4@����+�88��:1C,h6�$�O���O ��<�@�ilU�U,7n�N���)�@%Cbᙳ]�"�'�875�ɑ����O�H����3��;�B�=3��L�#�O�d�`�6m0?14	� ��>�"��32���W�k��l��x�P�'���'��'���'��Do�]C����P%{��,2�bQa޴uq$Ĉ/Ov��!�	�O��mz�!K��zQ����� >p�9�ʟ���}�)��ry:�l�<IAi��n>jU ��R:���r�K�<��cS���IU��Cy�O2�Z�cv@�I(^���E��O���'�r�'4�ɏ�M#T/�?���?��W8H�49�1@�+Hj�:bh����'���?������G�^���lZ+4{�T�'���EA^3�F`)�)�6�~"�'������Y�a�$��<P� ����'�R�'
��'��>��� �%���$	�|i�Lϻ����	�MS ���dX��m�?ͻ��ͻ���L'�1I�Y�y
0�͓�?����?�q^��M�O�|���܂��7���DJhyad��>A6mVő�`���O<��|R���?���?��x0�u�-z��mJNV[
�١(OL5oZ#����Iğ��	�ğ�둪�\G�9�d Q0z�\y���J ����O��b>rc��b��ѱ��̢,�P�qB/E�n�*FHOyR�GI�]�I iu�'���,X���f&^ɚl�bFe����Iٟ�I՟X�i>��'46�qzn����JQ*n	�Gj�%C-Hq���I��?qEY�T�	ny�
�
��SfY(�p�@��#��|�@�ik�	6�lli��Ok��$?M�]�CN����A�%rb��ìSFWV�I�t�IΟ��	����	\�'�v:F�N���f�#cx(��?���%��,��I�MsH>��NǿC�$�(��ߌ'c��[b(���䓇?Y��|�qo �M�O(���� .�e���0$�)��M� ˓��~2�|�Y��S�x����0�6\�	1�d�׫��b����oR�����py��c�Z����O��D�O^�'VK�L��#ɗ%�1 ��O�y�'����?a����S�ꀄ��kצ�% �hg�X� ���Q��؂T��Ӟwk2cK@�	&+�43�ʿ9Άв���!�<��䟈�I��P�)�ky�LbӔ8Zh�(q��r�Ε8K|d3�@C���˓LV�V�$�U}��'�ҡ�� Bk���үE�0�t�g�'>��K0������!�Пp��t�~��cW	D� ��8R.�<9���<I,OJ�$�O(���O��d�O�˧h�aT�_@o:=�b�Y� ����i�lݢ"�']��'��y.r���2|���YS�F
}�pФm��0�����Of�O1�Ĕ(W(w�N�	�7H��2�M3�,�@�n<n�n牛!S� 9��'�v�'�$�����'TṈ'�۝W����t [\J5���'�B�'2T�P��4��a���?����h�����^=�VZ%S��0�bD�>i���?�N>�4�ü+$`A�C
Ib(�УIt~��� <�u�4����O�a�I`�⥙�%o����y��K�]�h���?!��?����h���D�P��p�ɹT[=����g�.�d���VM��|����Mӏ�w�84�aRGD��InEdhb�'�r�'�Rm?7����֝nQ`t��?�d$(Vg�2�=��#��Qr8��a�|�S�\��ϟt��ݟD�	�����BũBh������lD��h�Py"��hQQ0j�O��d�O擟������m��G��	X);G���"�:�'Z��'�ɧ�O4��K�J��~¸�A�%�k��!���ϛ�N�<�eE !'���p��Sy�H�D���2-�b5@1������'���'��O��I�M�`���?���� S���D%��-��O��<Q¾i|�OT��'�R�'���A(%��gE�Hc��45C�ɳ0�i���<p��|h@�ONq����1p@�C��gy��Y~a�$�O<�$�O����O��.�0{9Ƹ9�@ �^�.�Q�~�Ꟗ�?a��?Q�i6��\���ݴ��^�����!��h]�4h%]20�d��M>i��?ͧW"m��4���פa~F\9sŊ�c�&����%V�}(����?iM"���<ͧ�?y��?�BL�>���F~�Y�0ϐ�?��������[��ş���ϟx�Oں@9�@",��Y�Bَ)��1�O� �'���'�ɧ��R���a���:l>�X�iO5#.E	R�8O�*�sї��S�q�B��G��p5��pd&�r��3'��R���ܟ�I����)��gy��tӘ��#�l8Lp���!"����U��e>&� ����a}��'Rd�&ʚ$ c�톭t�<'�'v�G_3�����Ё���	��ě~B�e����]|`��p���<�)Ot�$�O2���O����O
�'x���e�=�H�x�+�Lxj�Ÿi��M���'�R�'���y�'o�󮋓vU`l�,t��fjȰrW�u�	���$�b>e�g�@�9ϓ|�| �/I'J�<��Xy	���o��t��H�O�ŘO>�,O��O�L#��6�xxi\	|��l Ӏ�O���O��$�<�0�i0p��]�\��pz���;��d�>Kq��?�pY���	|��f*����Cv=��,�� �'�4z��E�Y8�P��t�ڟ ���'��9�N�,HEԄ�RO��&*�7�?���?1���?���I�O~�u��Fe�:î�!db\3uM�O��mZ�\���	̟|�4���ygO" �-ڥ�E�AŰ���ә�y�'
r�'M�(��iU�i��Я�?9 2��=�T�
�ņm�(�.H�h��'k���	ߟ�����	Dj��E��,(ĉ/tVE�'"�6��/p�p�d�O��d/�9OН���'W����"� W�by%
�I}B�'�2�|����W ���+E!G��0Ɂ)�<BNHl��	�剦$�e1��'B\�&�h�'��Qp�cϳ"�H`�j�4#\�S�'U��'�B���Q�h��4"�,���>��t��k�,4�be����� ��������o}��'L�wL�A(2N��-Kƅ�X�!��qd�"�������M�j�i �I��|4검�;\vĐp0-���
�9O�����sK* �1�P&̈́�x�E	8.T��?�P�iʶ��˟�`nD�I�����	1*P�PD#�4IV�L'����ԟ�\k�$mZN~ZwK�Xk�oÊx[б�gABm��
����]I�pyB��T5Ȍ�Oȉ[n� �\�h(��j�4H�� +Ot���|ZF�_�(E���T��0�jP1R ^^~��>1���?�J>�O �U*��"nqT C��Q��r# ڳ2/ޡS@��8,�i>�h��'�%�$Se�6�T��%h�����@�`-�lrߴ/��q�e�X�<e���S)�Lx�^���Ă�M�?��X�<�I����ɔk��B􎸑�̋�[ �%��ٟ���j�Ǧ=�'g2�[#�|2.O��ӣ�Yr�`���~�ڨ��=O���=a��#K|S@'ՙ�i}֩��t��A�<�����O��7=��#Xl���"6�&�x�j%��OB��?��i݆t��7md�� �%o�x/�m[a����taKE3O ��b���~2�|\�ȗ'��pP�M�A<�7M�V7.��Ók+��ꑳ~�����p��-�@<97c�(p�*�c��H��������Ih�I��k���*��%B dY.n�j� Ur�����#�M#%�����P?Y��PT�9E�W�p�6��D�נM�8��^" řsLQK������}�����f�#��	��M��w=@-b���/Bj��	�!�7*��i��'M��'���0|I�֓�`�
�l��iغ"�����'/t���g$O��Oʓ��O Io��%�Q�B/�?"C�����޴<�B��(O���=���~ͺg�	}�$d+��c0�K�O��$�O��O1��$9�OBH�N8�Gd���d��Jt�6��[y��4��D�����D��
��� ��_�bԻƫ������O����Oz�4���>��I�2�OW.a���G�lH�,Lv"��b�~�h��O��$�O@���4Muƥq�c��z���0ՠ�@�LE��r�V�S,������J~��nL���D�3�Q��@ҥvV�ϓ�?����?���?����O�z4�vh�RGjU�%ӈE]xX��'���'�7-�U��˓S����|��C &�p���$da�Q�&Zc�'�����b{����֝�C�`�Y`��0�\��F�N�KuM�۟��|]����ӟ��	�� �Ɨ/�Pa��ɆW�4��&(֟���pyrr�@�`uC�O��d�OZ�'�r �o�p�VS�僣sQ���'&듣?����S�$��f�����P��(1�D'9 l�j�b��x�P���T���0�B
A�I&��7�Q� �����&������`���\�)�gy2n�0��@Jh8����`�bf��"����O��o�B�����ǟzGF�)
� �bO���a��J����I�n �l�P~ZwP�X0��O��̔'[Vi��+ՄdN5"QO��2��b�'��	��8��џ��Iޟ��Is��ႌ?{Bt1��A�v�z ���`[L�6mR������O��D#���OXlz�e�MY�o��X:�H��xؙ�&UƟ��	e�)�S
X��0l�<a0��=@yB����VE<`Q��I�<�gϰr�N�������D�OX�
�q���s��2�(UXE%s���d�O����Od˓|/��lk��	ߟ��IZ)*
�)YF�ۈC���B�	ʟ��O��D�OT�O��h�n�lnP���m{"��*���%Z0���#w�ƥ$?eKW�O��dެLs�1�e�52$<�2�
�T���$�O���O��d:��K���1q�T������	Y�`�S)Ʉ�?�E�ia`��a�'t��i�`�O�9�(A�%�Ի'N\<�Pe1`�`h��6OL���O���C3ph�7m.?AG�"[x��)Me���u
E�l���9@�`�ڽ'�ԕ'��'�R�'y��'I 0�!9G��K2-�5�.�/��B����%b|y�'M�Oc����A�@u�#��)��8�bɊ4{���?����S�'_�����G�&+�������:|�̠B.���MS�Q����`��r��*��<�铰�P�� ����s���?���?����?ͧ�����Ec@��ܟ01K�{39 $��2fo̊c���I�M�H>i�H��Iܟ���ӟ��4H���q
�(��j��XHq���x�8�lz~B!EN�2�S�|��O�gf��!��d��'�6(�fX ����y��'_��'B�'���)��* �ݽn;� (��ԚP/���?���i��r�O��~�(�O���銋4��E��.�)#��+���O�4���:��J�.�eꥨ�b��ș�j�
|k��̟0U����n�Ijy��'�2�'��mQ���1s�Ez�1�N�,T���'���/�M[������O��'JuV�b�ʎ>涔�en��h֘�Γ�?iu^�D�	��'���J��7�ٱ/۠q�Uz�,�� �L#v�޴��i>A���Od�OjY�� �!=�l0ja�$:��A��O4���On���O1�.ʓs��&,����uAŦqf��� �ޅ��t`1^�4�ڴ��'m���?�"��x@t��5f�4^�⸉�^�?���5���ٴ��
!p���į۠<���$��.\U�'J��'��	՟d����\�I���IZ�d��.��c��1Q�@s��3$�t6�ڿZ�˓�?9����s��n >�����Ϳ�B@5eYY���OΒO1���{�"iӐ扣�<ŹT�I�~������	3��	�K��4���Ob�O���|B��FP���u�L@�Q�UEj�-P���?Y���?Q.O*�m�2'"x�'fB�h�h0휱z]:��ѯI�t>�'V�>Y���?�J>ia#�<g=�����7>l�����r~b��o%� ��i�ʒ�n�a�',Ҏ߯'5��G�Y&f�h�#�c�R�'���'���s�}�@�G11wn13�U�7Cʜ	�M�ԟh2�4Y������?qt�i��'f�w�p�V�F��r�"`U�$�<8��'U��' � D�fe�����݊$�8$���m2H8���tc@`�q,[���@۰�|B\���	̟��	����ԟ�`�K.���u�$�0ЕGxyb!Ә�� �<����'�?��+0�0t���c��[�R������Ij�)�(4�� ��[¤;TA|��z�Ҵ�zӺ��'�lЊ���g?!K>i+O�Q3NK-j���C�\.$���E�Oz�$�Op�d�O�<Q�iS����'(����P��ણ)5����"�'7�!�$�O��':��'+R��.@�$�w�Y�O�A�p>>Zʩ��i��I9p������O��}$?����.����B)u��ʂ�"�,�Iݟ4�I����I�t�	y��a HPgn�Wv���1Ȇ�/�e:���?�4Ǜ���.���'~�6�,����l̘��F��A����)E`�O����O���/)ݴ6-7?��A��	�c���2�)K?' X@+V$^�?9
*�D�<����?q��?�K>`�\z�c�n!����G���?1����Φ�X��xy�'���=��U�v� k� q�LP8{) �ǟ��O��d�O8�O���jt��ِ. ������B�Q7�|�F#_@S�m���4�l��'(�'����T P��0�Dě,~�Y�b�'���'!��Oc�ɬ�Mk��d���4��G�
���H��*�h��?���i�ɧ�4h�>���_1�|:��P5�xG�ǣl������?�����M��O�D�����Y��@�+�9E�����`��w���i�d���'�'h��'/��'*哶v�,��':�2����  06 J�4	�a���?q���䧆?���y���8����%�C� ���G�u���'^ɧ�O����i��$�>$�X<�u��xk\�`��?���ŃqW����S�O���?����t�2Z�|�G+��xD�d���?���?-O�l�
;�
����x�ɂ چ������/����)Է:���?�AW�4��ޟ�%�8z)�(8y>}qGʕp;<l٦m7?�↔G_F��4U��O������?aF��8+��Q�E�E<I�P��,�?	��?)��?ٌ���Oʽ�Ƙ �\���	*���R)�OȜl��1���I�pݴ���y�h	�/�kF�$[x���,M��y"�'���',$� �iN�	^�ndC�ҟT�cT��l@�a�?4�~�Y�l,�d�<��?����?1��?1G��<]���`�\h�`o�K�`�'S6M��{�����Ol�d!���O���Bg�P�q���f��8���UK}"�'�b�|������p0�d�Q�P[���}���D�iw�d�P�b��7�<�Q�5_J�:��%e5���s �f�Xi����[�F��&ȷ
B�e���0($�P���2y�,���W-J��	�@��o��|9���"#%zu���Z�,T�rc�K�A���B����?yS�?�&E�t�&��	��ͼ%�8y��Q�D�%��=>x԰#h�*BO( cS�T�[�r�C��;�>�B7+A��[���'
۠o�4~7��"ХY�o>Đ)e�оH���"�8|��T�!�	�X� ��f\<�D
�y-�8ãE�k�2�Cáʌu�p��BRӦ�(�NߤhgM�#F����&�_?�M�,O�*�D�O���91���X4de���6��.��K�� �I�'`��'�☟�8���]���'���$@R�L�v���i��	ҥ/b���>�d�O�D~Y @��(P�L�$E��D�ս+����ߴ�?q����ݪPH��'�?���TnW��b0q�J�
V���BL]K�'-��'�R` �'�'��)�qk`mse���vy�*e9�&������e������I�?�ۭOk�
N��L�ǧ�8�N��f%��B!���'��� �O��>�%�}Z�<�㣁8V�Ċ���O@�ه�j�8�D�O�����T�'W�I�7�`��㌌נSu�J�<�*�Yߴ_��P����I�O�E)�CK��s�jɾ.��������Iӟ(�ɾ5�`�O���?!�':L�1
�%�e�\:-��4��mN�������'�R�'a���2��(b��T}%�|ڄ�x�^��˟w�b��'��	��H$��X�,� 01�/�ؔ����9��R��4�<����?����(/_�j�c�P�1����tL��rI�>�(O���6�D�O���ƺ*8V)Q�c@5O&�����(y�4-��5���OJ��O�Y�D�A�OT���%P�)x�1B�L�P`�@�ݴ����O��O����O�s�P������4;�؂4(��`�^	Ⓣ�>Y���?����$ȴHk��'�?�`�W�k����Q(6A�p��or�f�'��'�r�'��8�����{����[�M�Ět�Yf��&�'C���@��B^���'���O:��(P`Є`&���0*4s�.ݛ �4�D�O��Μw4⟌��A&(:�M�K��q�_f�X�l�D~e~���'��'|�䮯>��~��@�勍�vC��ض]+A�}lZ՟��	0.���?Q����(0�d웳o���F����?��h��M���?y��6W���'���#���8�|0A��Hq঍mӈ8V#1�	n�'�?	�h�wj���ƃ�wn]A�NK�!	���'���'�,Y��J!�4��������)�-��!E�!a��A7k�`��%��V��'B�'K�)E7S\!���! � �G��{�H6-�O�Y��[�i>��z�W�ĕA'�ī ����	(ҎQ�H<������O���O@ʓV�,}�"��v�tM0&�� u"ܓ�I��_!�'�"�'��'��i�=�����r�Xe�%���T+o����<A��?����D�����ͧ|z��F�=:tX��>uz��'2��'�'3�i>M�	$ �T̀�E�g�l��f�:�J�C�O����O����<	0K	��O1��  5Ps�\�4\1�o�Y��v�i*�V���Ity�O��~jT���aQ�}�R!�=cR��!�Q�	���'��#ǎ&�	�Op���Z�j�"�!c�́�$%Z9KK\u�g�x�Y���I���'?�i�y�~�J	�!O�;3Sr�i*l��FD����i����?��'<9�ɋ/
����@3�lH�R�**��7ͥ<I���?�����ܴ��M�H� f�����v�n��(����şt���H��yʟ�M Q ���}����-}e�4��Vq}2�
�O>)#��Y�=�Yb��
�N~�q%���MK�������S��>!�C%]�ess
��{^TX�7�W�]�����D�'�DJ8��%b NR�3���{VC%ț�'�DCcV�@A��Z�d(�I���T:�eU*/Vݡ l����+��Q�'��'bW������ !����&�]v���8I�l�{I<1��?AO>9(O�U�QUkQJ��/eE�r�Ol���' �',�]�x�I�(�t�'S���0'��PH�ٳ�^8hG��m����Iy���?!/Ohʲ�i!�1�r��PpF�󏏲w%�J<	����O�+!
�|���_v�Z.K�bd���ơX3\�Y�i
�O��d�<1�^�	�!y�ty�� Z&t�ٴ�5Y��7��O���?�!�����O�����kLV%�^�
F����!J��'�Q��z�*�ӺS&���7#�d���J���Ћ�c}R�'���Y��'�b�'Z��O�i�%��A#4��s0m��C@�a�n�:���<�e�l���'DUt�cG%ŇtS��7ݽXA��o�<O�����4�?I��?�������C�<���õb���=�q�<�
7�O��O,�O�s�X��=::�!������e��$,t��ܴ�?I���?�R̮b������'���5���Ip$ĢB��ժrbE�z���'�'���<9��?y�����2�L�+/����R�r}����i�b-#K�O���O���?9�쇇a)�<K���&I��q�Ոׁ7�'��Y���I�����fy��1wv��Eo�#%�pX�N6�Qz��>i)O����<a��?��� jelϯO򜀕fˠ5x<9xWl��<�,O����O����<ы؃����q��Y3��S�
l8��_$i���^��	My��'jr�'����'�9�A�^'ZOb���"�Z@�U�R�c�����Od�d�Oh�?t�y(�V?��i��*�&�*P����W�9ä�A#�`��d�<���?i�'��a̓��Ɏ9<�`NxCK�TШ�Xdd{�0���Oj˓��0��Q?��I��|�S
��86���ZFl��aV�g��p�O>�D�O��T�L�Ĳ<����d�]�,�(5�6�Z#S=*Z¬��M�)O��9Ca	Ҧ���͟0���?�Z�O�V� �PX#��ǖW|~��UÓw���'"����y��'B�	kܧ,x<��'0]��Wӌc�ڜnZ�����4�?���?)�'G��	fyB���^�2�2�dӦ��|��úki 7��9���O|���OSr+��f"���Ʀ��K�Hz�`4G�6�O��D�OD�P�(_}�V���z?1���1.�Px;RCˠ`h�
�]ئ��IJy�GD�yʟ����O���ױFJ]p�d �.^%s�,� Pz�n�,��`�����<Q����Ok��P���"3OP RH����5��I%x���	���	柈�	ʟ��'�З)^30��F�&��q���M9%8 S��'[rU��I��h��o���'Ɋ� !�z�%��ZW"a��A8?Y���?	��?9,O��; 	V�|����,(��h��1E�2��B ��y�'a�X�|�	ޟ���,Qi@�I�YP�T�bɕ��O��E��4�?���?i��� &�^��OXZc,-Ё�ޘL$�!��/&}$i�4�?�+O2�d�O����)����O��	/��EJ���6E<P92i 7`G�7��O����<���]��S͟@���?�{]�_���A��Pb�I!`fQ�����O<�d�Ox��=O���<q�O���[AJCr���S)-{�P�r�4��V�b(��o�����	۟��S&����TU���W"�@��fG�1J\����iQ�'1R�'��ޟ�}�(�H����d͖^���葩����L���M����?�����V��'	����Չx�\h�1�$���g�r�j�AV>O�$�<I����'�\M���,)��b�I���\�3SEt��$�O>�d�:VgZ��')����I��Z��˘
>%�rk�6S�enZڟ|�'Y�=阧���O��d�O��ZC�٩��dR7`R�o�H�D
P�5�In��Q�O��?�+O��ƮX�㠜�b�r�k�d+W�����i"rI�yr�'y��'�2�'�剝*4�ɓ2��O��!
�*/O�"���E����'J��|��'Kb���6�'3�]�B��^��k��'v�I쟀���ܕ'��U���i>	�&f@�'֜�ƙ;A(�4��d%�$�Or�OL��O��7O�c��',N�!6�[,��P��C}"�'���'����ؐM|�ǝ~"��Ip'�c��X+#��*���'�';��'��hip�'f�ILʽ3�nF-in��5�=2Dmm����	by�
��&�������꽛Rg� d�p��Ue�$��U#�N�I�L�	���IV�	@zc/��OP0PXA�ʊQ�Q$��˦�'[�(K��z�8��O2�O���S�? Vp�0�T
`�5	u��"̄x �i�'����'`�'�q���
4+J #p��ф��#7�`M�v�i�<� hnӄ���O��������>14k�F�z}��,�!V+p(�rFR�nf�v� ��y��|��i�OT%�陛y���cF���x����Hئ��џ`�ɚc]iK<���?Y�'(H��8!Q8����#"�`�0�4��l�"��a��4�'��' Rp��V����c��V�x�#��w�8��ҩ}<�%�d����<$��آ}�� �A\����V�R������ ����O��d�OBʓQu����摰LȌ��=gf��$E��bm�O���:�d�O��d�5MjR9+&��
�� nb*4�f5���O���O�ʓy�����4��`��I��R�k�B�W�N��EV���	C�'��������#qͤx �L���朷P��݂�OP�$�O$�Ķ<1vl�<q8�O���Ʃ
�u��=`TF�$p =���gӺ�=�.O\��.}���[���������j�$^��M��?����?AS������O|���B"�0�z�0��ڐ{�z��qH�a�����'P~�C���TX8��J�Vl�B<'9�|�g�i�剦/���ٴq�����Ӑ���P, \����\��C�b��'G����D������yxvu�ÎҦI<P���M��.�?1���������O�V�qZPΘ�H�|�[����x� ��rQ��D �S�'�?YQn� 7�n�����:x�$�c�Ø���f�'<2�'�6}ZU�?�$�OJ������ED�P ���N	T�j#<�	.F��b�`���h�Ia�$mhq-�?�*��Q�7f��;�4�?�c��c3�'r�'�ɧ56"B�$���f��7�-"/Q3����~1O��d�O��D�<#BNs8H��e��uI.�"��.4�V���$�O�O
��O��0O�8,d�� d� j���0GΟ{�1O�d�O �d�<!!�M|�)��[<����K��UB� HkR
ps�'���|��'��l����H .�t��GD����jj)3��I�I����'č	v!2��i�������,�j<b�(J���En�p$� �I쟰!=��98B���'�Y�cg98�`7-�O���<�b��h"�Orr�O(Bܚ"�^�u�\t0�e��/��B3���O\�dC6��'\Ō�Sb[�0Ԁ�@P�+~8�'�2�V2���'M�'{�4[��ݔ�H�KW�&fk�I"�J��D:T7��O��)e��ExJ|�A�")=x%�v,�؇G��=ƪ��M����?����r��x2�'��҂��9g�| h�X+qa>�O6�DW��H��f�ȫ:t�'��4"�oZ��	y��F��' �W���h��\�� C@��J�0g�'5��'�B�p"<ت��yD�u		?$�:�o�ɟ�$b��ē�?A�����[��AkRh53oI�	X@8�y}	M��'r�'
�I��*��R\����5V���'�+>�ؖ'��'�b�|�'���H2t�a1�LD>��u��?e�6lь��$�O*���O��Z���f6��AX��J%��u�aC�,\�e�$\�����(%������G��>Aր�]���V�O8�V�z"lu}�'Z��'z�	�HUO|B�Q?zA5{�����4����BɛV�'��'�B�'�P�3�}�A�u����Ќ`�r	��&�MS��?�)Oԥ!� z���'F"�O�0��h^��i��P��,�>����?���^��4Γ�?�,O����n*r�q�ʕ@��q�0�ŀs�7m�<�5�3,�V�' ��'����>��:����AS�$�6P��NB+�F�oZҟd�	�B�B��,�'q��-�V$�F�\3���~h2ͰG�i� D��|�t���O��D🬑�'��ɸ"	�1���F�(��*�vtt��4&&͓�?�*O�?���1;�H]�`�	&����s�˛'�|)�4�?����?9"���Sf�	Uyb�'��d��
>�K���g*5���'L�f�'��	�i�)����?��
�!1GS� >@�˕��\ ��i%��\��p����O���?�14}�aJD@,3�MӲLʡt�q�'�f��'P��9zx�%�`�R��F�O�|�b#
�Lu���&�J�6�BXI�'eVaq&M� Rf��/&���$[f�ܤq1�@"`�dՈ���Wv~5�v ֒6;�p �'��_|f�v��3O;
����6R�9X��E>o��mS�"݄cV�`"��k�4R���-sC�f�_��,��&�(�(�a$�	9t]�[4��)Gj�)��H.���g�M6k�^YSB#X���\Pw�D#A6&�*W�E��Rhq�C�y3f*\�<�=+@�',B�'�b)i�V����1�d� 6y����R2'�Ťj�R��姐�w����'MY�'��Ax��,]����!ݺ@ʛ�I޵��-�$����٘��K�&у�l������O���-��`���^�fp�ɓ@���`�
�l��`� �,7�t�h��Z�WK�U!6M:�O�A%�$I�L�-W����@�19%��$�x�̀&k����D�Oʧmh�����?I�r̸$��,}�}�@�6cnmp'��]M�ʥ>uVĒB���%��Ot����8>�h�s��k/�G�:XU����a�/�e�Mǟ"~�)� �d
P�|,�U"V�E�*��+�%�'e����O>�S�K�U�n��v�̀8��d1šC�8�ZC�	�~e"���D�G�\h�U��yH#<a�)E�ݼ2+�Y��ƒ�CS� �?Q��X� ��U1�?Q���?����.�Ot�d�"@~\t�ʠ$� ̂A�Ό ����<؝����T����	|D컵쓄4��]�ҁ�����9R���W��B���W��I�G�,"9�oA�=�2��>�dm��ܟ<E{�T�t1a�P�*�� �F�	Z�`�$D��f#�׀C��,��!
V���HO�SvyRE� F�6�I�TRl �k�� ��z�N�����OX�D�O�e���O<��y>��i�=M�BJ�%*T���:GG��S���mV+�h%#6�Vux���FJ�0:���"���W*r@��,��tC�W�R��t6��Mx�h[��O����(ݴ�*0.�!��1�� �)�Z�=q����{ؘË��\�=iW�H�!��KԎp2#�B�}L���!����X}�\��{%�\���d�O<˧@�6�"�Hɶ9�B`j@!Q㎐��M��?���?�5$DtڄN�$��0���)եt:���!�m��ɑ�b�0Q�ؘB�C>�l�v��[�RU$>��pR����Ā�!�\q��#�h�0,����8�ꀀZ��dzt���W�)�D"�O���֦�%�>��Ai\�D	$�9U�'LObى�h 09PyAʗ8;�<��t7O��;!F�����	՟��OP�}E�'�'���Q7jK�rņ-k����p ��DC�B�T>#<���I�y����
�Ew���ᣘ	KM@������O��B`�ݧp �y�E��rt:�`_,���D;�)��Tj�OӉ_Ԕ���U�#N�1� ;D��T
T9�� �3n�6�p�d.o����'H�y��lݨ{f��q�����?�3BU�l&��`��?���?	a���4�4pp�	.)6�<�' ]�I#H�%�O���"�'! q���/	�<{�͇w�TH�'_��i�_�=bt��2��ցאp�h�@`����u��H8D��B�q+���;+��=@��5D����m��`�X��f��eӷ�HO>q	�����MkFţ\:|����; �9T��?���?9��?���8��?ɝOX�\���?�d��;]�v���t�Y��E��L0�|	���ÀGp�T��.�	��	��SY�|"����?�����h*���=+�6��̓~��ȓR(���C F�"���`��g/�ȓ<��=��AJ�%�\S5�(�:��7�O���M٦����<�O��u�4��b���5D�5 ��&�*J�"�'#rn�
K��T>��!葭&v0�Ň3��s'�=ʓTm)G��Ē�n?�I�����˶Ē�(O"�p��'3�>{����y�V=P�.�����./D���CL O#��
'�3z�[��?�OFE'� �c��!�� ���$�@�k�'|��ʔÕ��M����?	+����C�O���Ot9
��@>iP��S+�=� ��MU2w���$5�|Fx��e\r��'���SG�*^�&���)�矨�ǤŦ
C���lC�&�Ԝ�gψ�zHZ|�	i�S��?�ҤFL��8�!��x�n�z��N�<٥�/#|���MgZ��B B�'\�#=�O����"�7]q�Lk!G4>��C��'"hBL����'���'�2w�-�i�Y'PpΥ�U�:p��L��d���)�O�Y��֦i�h#)۰lL欣�O���'�����(!���A��:l:�'L	a����=� �tbY�T�ҥX2��ӣ�B�<4G5>�0��qkb����?���"|�4��'A��)��y p����k6,� �n�2�'.��'x���'^�4������'�r˧R���dH	{PIE�ݠ�p>�#��uyb��c����e��({��.jrȅ�I�X�h�d�O�]��S�d݆A�����=��y�#<���O���<�)z���9T���7���_E�Lh��@�<٦h�r�H[�L��[�F�#�<��W� �'5��K���@���O�'_�����U��Ƙzw�X*ed�12�W:�?����?�6�� �?��y*�^P[��N3Pl��ζS7J�)��	%#���j[�%�.$���!9z:L�Ҋ�W�'�0x���h�� �Ux��C<��KG�$	���	�"O�@Z�.�����h ��`qd�'<�O{����glV�Ԥփb�B�p�"O��1�N�QU<M�t)�#�tA�"O��p�&���={�;U��|p�"O�����C
���מV��$`0"O�hrb�&(��mQ$��i�D�`�"O$�bb� �6�dx��i$���"Od)�"M�-�P�I��5�P���"Oj�)�FH8W�v�l��^��!�"OT���Ha��dfZ�8lv���"O���+��lk�8(�"C	o^�,�V"O�l{�*F�3��/�!5B�tXT"Oz�r�(��f8�d�(P��!�"Of����\+@�L���$S�yPQJV"O��%G�X�<�b.��mU�'"O�9�,�#k-�� Kd��%"O^�[�)g1�� �MX(>BB��&"O��ҒHL0)���X��ڃ,�TXr�"O�,�d霞K�rP��&۷t�ژ�P"O� �/ó<����}��!�Q"O"���Ƨ6�������.���3Q"O��S��Y,����Ɲ:'��)�"O��x��6yΥ vK�?���X$"O$�t*�1Q�j;'wt�"O�k�؂=�T��#�J�C"Ol�	� ͥb)B�I�ҭ{���Xt"O��`�RO4@ѻu`\�2��"O�賡%Ѻ@���Y��P�Ы"Oة3p Ҭ}�>\`�g�(/e�!��"O�%#���:xI�8�R�Ѭu�ܥx2"O��vDJ�t몵P��R<"�~�[�"OD�À�XD��=�6�
J�����"O��:��[��Z����B�|��t"`"O��)�Ǟ��4ͨ�㉡1���Y3"O�L���V���BA������"O
L�6�%.�I��ʐJ�|hYU"O0p�g��Av��(�,Qـ ce"O��1�(ګ<�l@:�N*����&"Oh$��܎C�n��3-��<w:�A"OQç�3=�T	�0F����Qr"O��y��ׯ*gZ�q�,D??~fi�"O yb�	f�@���sSĽ�U"OX.@�G>�0r�cاjMP$h�T��(B����=Q���9��!��j�$*���c�Acx����@!�?���Y�}ڝy��4!j*`����\�<���_��8��gR:
����V
�n�'� ȲS�^��h�&ݨ�A�T'���m,1O
=�4"O@%��IOP��ʬui0i�v	T D6��t4�)�矌{�`�7u9�Q�R<3��0�h0D���wɸSS����
�>w � �VM������R����ۺ-#�p�υ}�l����H�4%�|R&[�'�´��^�(]X����0���Fm��j;�Q�ȓSGL���`�xܑ�U��$$@Dy�B�WO\������&m�c��R|��rh.�!�RJ�)�w��>}�M) �/(��a`%$� ~b�"~�ɾxX0�a��B�P����"&�C䉩_-��x�-�#v �,��d�A�˓l�ȡ3�'��-s��.4H;7��{��I9t�H:��݆�I>���*��u���l��D�j�DN@�fF}R�˚��>u�s��N�t%���DN���0a+��T���J�Q>9��'�W_�}r2�?�}�������Q�S�O�u�塀�-丰�'dĈi
HtäJP5^X�
9��)�矜�jW�G*��i�"p@��e'$}R
D60a{
� �up�f��+9��j�+%�z��0�O�}�`� %P{L	����Ά}�*6M5g����\��	��Z�P��|R&Yo�R)��͘�1+R��*�0P���a7N,=��F}2"D�m��>��qbV�[�+W�K$rm|���."�Y�2ܡ�bW�_�#|��!��6��j�@��& �V��C}�W�O�>�s��Ǭ=8�@���O�6��@83�n�#�PP�ӧ��r
��Fv�Y�n
�mm��j�����yf��~Mly�GD/�XY��!����<*2�8���x��liffT�D�a�D�3�Fq�d�3D�8��T?h>J�h-�#<�� [�C�I>?���sF���2�<�Ѥ\(_nB��?YX�Ӯ˾yO�y���Ȁ��B�	3t��Bi�"�H<CFJ��S�rB䉠"�p��Ҙ�2O�&ZB�I-��`i�Q(]�� e�*B�	O�HY!�eI��u��盵Y� B��(i��q(����
�P�C(Ŀ>|�C�T�vQ��%�*��4h�)��C��"W�d��[�&�c���q�$��"O��'�1:}d(qV
O+Ҏd"O�9k$J�|`��
�����"ON���0M�\����"�ZT�"Or��ɍR�����/~�La �"O����h�.+ظ��L�;>x�� �"OlxU�^�����! 5��!w"O�L�m�$����E�-,��9q�"O���*R���T"$&��G|�h�0"OtIP�C�J3Ly���U�ra�"O�Tc ����aC�1N��)�s"O��A�O�`@���3����"On]@p�
@
���F��aj�"O���E
8E*����n?%�B"O�hK�(r\
իH7Pe�a��"ONc#aL&	�@]D�Q/FMYr"OΤ��]r(E*�)Q�?J83'"O����dŎ8��x;���F�b�"O@0'�WIs����O	;���I�"O(�9���_/$�i`���c�"O�-�� �bK؄"���07TK%"O�0�bA^�<�h�<��ɥ"O4��#J�D�>E�Df��.a��X�"Ofu���O�A�:�Ҵ$�x_^x�s"O,��W�Pq�LH�䣙�`��U�"Obuh&K��J*����] ;{�p�"O�r!OQ�-t5Sgڗ\�x�4"OFY�@�]�t���˺u��zd"O�4�4L�IV�Z�/_<�����"O��I� ��R�*�;P�O�3���HS"O���� �3��X����{��\	@"O�P��J�L��9�Ta��1��h2��
��Mk&�kPd5�3����zAR)C"*T�d�e٠�$i���DP�$M(��a�$�"�kǆJ-�:��S���.�� 
�+#�HZ����9�z=�fk�37q��㉁?���u욯a���(|B8E"I� #�4UBa�=NB@B�IN���XC�TO�.i�D�$���'��}��.jA�ه�S2Y��	Yg�eY2l��0��<�
�P��ǅP0P��a�J+MP�����_O��6R�������Ӻ�C�OLAb&F987%��%5r�`d
O0Ӱ�4YY�Ց�nį��Z�� ,Ja��Z��l�Z@���J?��b������D���f�	 0 s��'�I-RPҌ��J%2�����2	Ϫ7Z�U�"`J�Hޥ��)�禡�p� Kpp��fި��6$9D���"A��@;
�2C�=���""�>�W��}�|0�k7<O������/�,��B�;�D��Q�'�&�;ӯJ�u�� (�R�&d�1"5셒�:��:4�H�
5N�"Y�@A?,4I��C1�J�eH���*Q�?������1�$�ޭx�� 
ф-D�D����H��ʒj�.~&l�j�zx����/1���`K�"~nZJ��aZ!�D�p6�|@�(��$�FC䉪?=VH���;>(�����-�T�]]^��ȝ�ސ��䛹/Z��唧+�~�rP��=.a}⬄���]p�I�x'���cOҧ+�� z�cO�O�,�Ɠ:��U�EC�3q�2C��App�Gz��G�=���'�H��}@����0+�y:b)�3/F���ȓz��ڄ!�2��z��[�8`o��9[���Sj�O�S��MKf�X:^�	Z�!ՆS��I8�!�]�<qH�2IFR1���?!4@���cy�̗
d�~���'J�D�Ռ�~0��F"J��!�
�'�v�2%��Xǒ�HA��;q�,
�'q`�A߅�Y����	�R�2
�'3�U3+P�S�yrc�Ŕ2���
�'q|�@P�����T�3m"=�n�	�'���� T�:@�*��<*�"	�'9ܵ�!�ļg�v�3�&F/p�0!	�'��Y�W��'>E�9ٕ���ti���'��mq�D��.�԰5�� k����'��A�.�� �*���+�'�J��0+H>_��9��Q( �@���'ݤP�vm�]߲�b.P8z\l!�	�'dx�c�.H�E����$g��	�'�Ra���O�a�j /UbL��'���ѡ�Z�'�.��4��=RE�yדOd"m��>��MD8Z��A%(�"z�`!z��y�<1g�͔h�J9����|]�1�� qܓ*Ȉ|�Ѐ9���N��S0\F�	�N10]@r"O�dЖ��Zh�M����h� ���+Ji�qO�P���Y�|��������	fF��צ*D�����ݒ7��ؑ�Nvt��$ǚX�9�>�OHq�fI�i�L����:���J��'���A��6?�L�q�Tę��ͷZ� s�EF{�<!���Id��p#ɴ�<񖪑u�<Q��+RHD���lp�(�q�<AbM�52xLa�ӄ6˰lPrdLr�<�֌�69w޵���8"t@XF�AX�<��,$(e�ɋw�?T���1'R�<!#�o���k%��>6�f<BT�t�<q�@N�wT&� �cD�h�
̙7�x�<y��G�qV���58!���"s�<��F�UW.48㏎�xB���Ys�<Q&�߉-��B0|F �P��f�<ɰ��:g^��G�ԭ}ڈ�h�f�<���ʌk�(��H_	  3�a�h�<qe�V/�Ƞ!3���5�Nպ�+MO�<�oӳ�x=����0B��$�Q��c�<9���=A�L#R�Y'���e�\�<YG	�v� ��V�ev�#��FP�<ɦk՛� M��Ì�@�!��f�<�UL�)��J� 8]b}{���}�<)�7 �@��ըM�鸡�M�|�<1�K�,c����hm�X��`u�<I�'_"8���#˕,m�!����r�<yT(�0
�x�
�'0�̠A�^o�<y��A�jv��>
��(_n�<qՂF�D�0�H[�!yԮ�h�<�0R� �2�0"��T�M�Z�<I <s�j�8E�	q�`=
HS�<A�ݱ]�
aZ)��D:�X�fWO�<���R^�'��X�b�a�r�<� v�iǮ٩����/R��J:�"O܅�s.ܱ?;�@gOВ<d���#"O��3�̽9Sj�(�뚡
Z8=QG"O�ڵ$�=����<0����a"O<��
�	R����qH)��"O��B�:K,��ʥ��%o�iSW"O�4���.\	����dax1��"O8H@5@[�p=���^�	W\�8�"O����3Y��9�ω	q�]ZS"O*��_!��j�iوx�\<h�"OZ��a�0U{�l#�(A��rM�q"O:��	���TB���.[��` �'I2L�g޶,&4q#��v7p�:�'�J�h�l�.x\���%u�<�
�'H�N[�c� hQb�JB�x�b�'s�@%�;j*���Ý9Kx8li�'T�id�<�(Y���5-Ȅ��'�
(�����@7�SQ*\�,mMr�'Zyӳʆ���T�u�Q��~�A�'x��SFȵt�Liť�.E}����'/ 8��%;����[	I��-�'��QJ6�<[+ś�B1H(Ni�'�z�d�b��@2��uY	�'��0F�܂X�ʵ�	�'�	�'�\m�5у/�H�t��2(�ȁq�'�@�3�ۃG/x)��f=��?D�,{0��k6lh��F	�(���1�@0D�l��@_$S�05��jZ�B�"bI-D��C�-���C���5�t�K)D��xA&�"_N��Z�R�`�:t
r�<D�c�@�Ny�F.��)A
��V� D�
6�ƃswvt���L%e��A+�:D�t8'$M!:��"g���V,��6D�;�E�#{ ��WJŎ6G�4D�L LɳZB����-�1c)�=	�*2D��0�OA�R'�"��f
�i�`,3D�<;#�lV�8��K���q�/&D���b+M�H�����El��d.)D�d ���r���B.��,Pq���%�OR�����K����.�8o
���M�<��ެ�pEC߹ ��x*`,_R�<�5�H�g�Z,ɠ�ٛod�邑��b�<���A�:I���>-�9��kC[�<) ��-��˶]O*,HR-N�<�db�br�X��F�9(��W(�M�<I�ܻh�L�q4F
�]rD����L�<A���MÜ�
6
� ��B�JE�<q�؍o����cnE�\6z+0Ō{�<ѷ�۽T��
�瓵M�[�/���JѰђq�F���*ǲ�B��ȓH��2d���Ht8�JIK%Q�N0��FȄ���h��>�D��@EQ�nQ8$�ȓO���;��>�P��&�_08��ȓC�ӄJۄoÔĢ�N#�����Q�d�e�W�V}�XR��B�G��9�ȓ��3�CԍM�vd�p��z|�ȓg����OP�@�Z��7HQ�TޢY���� �q�� e��ц^�X:���ȓ��$�q虴5�zhC��ͣ$��e�ȓZ��"�+��3(l���ͦC�pH�ȓD����JR!WV���o�	.4t�ȓ/8F�ۆ	��QBF͇��؅�I��~"c@< ��.O������y҃�̪) � �:��` (Z�¨O��D�� ��WF��X�D�L�N����e"O>�Җߨy��\�|9��OD`Ez��)Z-T�V(�!�ĿAE�j%N,!�D�/�`f��u�X���@1@�3��|�gZ;�.M�*�|3\��*�yrKX�hk@���F�s��X"�.�y���l���'��=Q`���n��y��Sn�f��G��22;t��G�G�<�I�(�v��M�1Q���r�<��gU;^�Y�t��Q�X!��Oz�<���R�B��,:��M7+�~uN�<!vJ��Rt�Y��h)�ԍ��\L�<�d�Q�;����W##��R7�G�<Q��a*�E��i�
� 3F �D�<�%-��lRA�G���{��um�C�<12�U�y�a��;�X�ږH^t�<Y��1}�7IQ����#Yo�<�5�i�F�)u�B�
�F[v�<�F�'��2 �	.L��&�Y�<AEI�)UD�;�hQ�v�I��J�S�<�� >Wb	�B�ѕ5Epu�vF�x�<q9�89���`K^5��l	x�<���v��@�o�`��XkUc
v�<���è#VD$��كw�~|��j�t�<�6�ԥkz��ׇC�*s�
f��q�<��8%�b�F�ĔdRZvaFF�K���O�����X2"f@{B�̌G5&��'xBq��i�!߄1��ɉ�pȤ�
�'֠SH��W�BhѓEN�lb��
�'�;B�#	���Y G�a2�Ta
�'-ԸQ*�@��|��$!X�|�	�'�����L�Q�� �.^7^�vy��'|�[`l��5�d��oJ�"�Խ�'�*�Z��R)�܀YC�� �����'�,�i�)�)
�"i�7!8Z��' p��V�G���0 ��\���'ͺ���ˍ�}��`b0_�h����'ֆAd�E�@ގL1����h8�'H$E:%J�.�2�:FB �Q��1��'l�����Y*���yi\A:�'��(+d��&f�%�kw>�z
�'���Ye51������>^�܈�	�'b�����2�s�U�rhC	�'��ԋ�"ҢE����򯎣��1	�'^����K;���2���{�(�J�'F��V�S�^�����D�,�
�' ���RL�=Yzހi���=W�P��'����҄8�֭�6*ˌ �4�K�'�<5�'��<N*X�B�P�r���'?6��Qw�YC3�ʍ`$$��
�' 6Eh� dxș�U�ϊ��ݻ
�'4H�:��Q86>��CR(��s��a�	�'��}��g�/N�jUK�K�}Z�K	�'풉�K��^l���D=v�v�C�'�J��QӸIk�M3t���p���'[4��g �
i74��sn�#tw)
�'��L�gphfK� ����'$�EZu�K8(�+�"���'�%�穆��
]1����te��'O��ϕ�|ʪlգ�Fٚ�I	�'�h���GW��-���	�H ��	�'".���,��N��USA��#&ț	�'�z���2o�੗	}ܖ�	�'nj�{�F��K��Q�7�^���	��� �����D�s�|���Տ�* ��"O�J�[1Q��Iv�͠Yw�i�"O|� ��>���h��y��S"OI�����9c.	��X&2����"O ���e��!���R�n�@Y"O�ta����L����j� �X "O�1kT�S?p�T�*�ߗ?�D��p"O�,p����Uz�
a���!��"Orlq���j�剋�M�t<��"Ori����#�\qI�H2�K"O�	㓍F'�����: X1�"Oj��w���&p0W'əb؜c�"O�����L.�4�GGǴ%`�yxu"OzM��IS�-s�[A'>G�a�1O���$�� �T�vtV(�U�^��!���K���B�b� ���h�:h�!�Ď
�#���g�"�AC�#�!�*�u�)R5� �C��Ƙ6�1Oܣ=�|�ף��+��B��ť~dz�����K�<I4�EV�����\��h	��E�<AcU�&�q�M
���VJ�!�dԔz��q!�9 mڙ���Or!��N�0���Zu�׍v��!��'x�!�d̕}��sTj�w����Db�!���)>6�x���%�uB�� `���)�O��QD!�3/�R�YD���C���G"O��A9D�)C����U�w"OB�)���S��)=�,�D"O
+EM�!E4l5��>��,Bg"O�)�@�� $���ƃO��	JG"O )�D
ԏ2J��B�fݲ����$"O��A �+F8�)QHJ�=}����"O�ԋ���S� �R#��
3���"OԐ�DG[�&�6<����nq�T"O���ӏa��p5:�W"O�\s����y�d�ۣ|'���"O���I�T��RGFمy �%"O�3��ۣ��52DE�������"Of�R��.�AdéS���"O:ԃ$%Q&y�Q"c���� �4"O��9Wi�e�,��p��Zm���"O��b�aO.>f�ԑ7"�3h	��"O����/Һ?(��0c/S�kJޅC�"O��#�>�$K#�\�I��
e"O�z�@��Q��x#!��_�"̠�"OFa�l��0���`i�.foV��p"O��9F���� �o.8�"O�lR !�.C@��E�G�y �:�"O�x�')�>9�@�͵z�6�7"O&�J��=2�Q��� `����"O>���D�&!!0m���4"O����6�HXVL��|p "O&�ۄl�eb��qk�=9z0蓢"O��`!@�Z��� �J��O
5� "O ��B�A�(�Y�ܸ&��X��"O�a�8����BB� ��A�"O �����&҆�������"!"O����+�(��Ո� Y�
�&�a�"O���@�D�{UhT1�o�	l8���"O�|{ť۝d�p�XBoE�T7�\��"O~�Bύ5V��uXp-̇B���(�"O�J�X��p3��2EPh�9#"O*���K� k���±�
LF",�%"OvH EA�y1�|�2�Y���Daw"O� Փ �E2|eb*4�)6�`͒�"O�!RlD��i e$�0rQ�"O��@cP�D�R�q�Yu�p���"O��X��ıg�5(A�)��"OV0kp�ٞ7d�I��j���b3"O,u��n̍:c��C1@ʅg�t�1�"Ot��,��'�,{�,����u��"O�1��+͸N���S�%U�
�(h	 "O28���ܙe�,��[�q8��Iu"O$Ѻv,
*E�B`b7"�H%`���"O��ؓbؚn��X"�W�N�b ��"O�T�ӡڤ,xX
W�ӘI�l�A"O���է�=ںh����y����R"O�I�3�J�^�$�����܌:�"O�y��"
;�*���������"O�qBw��n�NQid����P5"O����S�Qĝ$Ɯ
M���P"O��k�O�dT�X�A�`X�u"OvѲ�@�+��Y�w��>gԡ�5"O��i��nJ�hڗ#�-flA"O謈�C�*U=������Rn��"OHZ$)ݦx�Ra�cA�bvh3�"O�A�G��	tv�Ipd�|r��b"O(]��&��{Bt�����PH�䈔"O�}����
3�/P<4!S6"O�)��_M�ؑ4녧=�p�"O
����0e��	�"@N�i�`�E"Ov�3�I�=�nP�.̇@��"Of�kT�_f>�1�,Ⱦ#׬�Bd"O��)4-J�y;(t��?#�]#"O��$�L��;tl��b|M[�"OB)x¥¼Bl@�
�y`,U�"O:��G���a�.e0�̀�|S9Z�"OL�ñC�����['خ�N�[�"Od�y&j�^)� �v�ߓ-}ȵ9�"O��١���*�las���9�QQ�"O��S�g�)�Dr-4zͲ���"O�	�F8i0i�U
ͅ��x�"O���0fԶ��Z�/�ߴ��"O
���L���8���ͻ"�b��b"O,���K�r ,ٛƭ;C�$��2"O}�3��(�l�m�y�"O��x��	ll���WK\xPX�0"O"5ʆO��,;��"nH$)#D"Op��K�:^D�=k!���|ڤ��"O8�c�,�#zx��תԂ`����!"O>�X �5_�ftRf
K$S<"Љ�"O�	�bB��FU2�46Q�G"O<���Ý*7�a���3y���2"OX��ȏ9RkL�3��CZ�$��"O�Q*��A�k���6�S�{�m2�"OH��W�
"&�:��14����"Odd蠀�/&��b��E�%��1��'���3�ݝagH��FܓU���9�'m��j��^&�2ջ��$Y�k�'涰�H��_{J@�aD^%p����'a�����{�X<{�eI�uM5	�'�>��G4B�\���5|�؃�'��])T�]xHp1�б_�����')^���MW�@�ܥ3@i
D���J�'v(��ċR)�|҇�&?�n�1�'��m�-*��7��jc�"�'}�0PC��>TqF�0p�W�e�0A��'5� ��Q�j��I0Sf_5aq�Л��� �h���}��Q-0�̄�q"O|�y¤�	I粅��d��N�e"Or����¡#R�����	��"OF43�aS�^�P �G:7J���"O��cN)�p�B�FUW�8��"O�d�и	�,\�P
,E`@��"O���v-��f�[��_���"O��)tKI+mD$qrW�	�8��@Ӵ"Oxy�)�5qL�a��Nmr.� �"O(��wN-������� y����"O�!3B�';�R�@�Ax����'"O��:�G��QA ,W+x�,���"O���AO:X:�T�)G,�Q�"OvP0��3{Z���\I�U�6"Ob��PD۟�x�L	y�n-��"O���/E2�2�kW�G�*4Z�"Of͚ )Q:-�E[�
��o�X��"OJy�l\��^�ӫ8�0��"O�����|�7nv�`1��~�V��ȓnM>�Bw&>n�sKɄ}��E�ȓ8!�  ¿?����n��7��y��%�(:v���o��| -
	8��لȓuUPT�'  �-8X�����C��ȓrJZ8�3E��
�A�^�����ȓm ��;��Ā�4�T$��JHA�ȓ(D� �����4��13 H�>�V)��W�zPH�>h? mP�e�q2�}�ȓa�x�CG�-+����"`�=Z!z��ȓ	�h��G�`��	�1lE�k9�}��[�R�N�I\���u	%r9T��ȓ^��4'�.L�C�̠c�Դ��%5v��� �Ƹ.1���K4�8D� bFbK5o�E��(�C��tS��:D�h3&T�i ]#��P�qJx��u�5D�P��L��H�Ҕ�ҹ���P�`0D��u��^_>|;1�Koh,�R��"D�(��έq:+��:!fj��#K"D���f�ea�)�#M\���'�$B�I�V@�|�w�ȍ\��b�_���B�ɉ:�c鐑d��e馅��hB�o<��LX$X�� $ݎAd0B�	:rsV84��b�L� ���[�B�I�<Z�H�J'8�-҇*��K��B�ɮGnFTX6����1�BF��\
jC�F
δQCo�:`.����ُA<C�I8U��O���I����`C�Iv3�|b�˲?�����B����B��A`���f�,=����_�n�Pg"O�+Є�7���� �ma�@c"O�e�w���&Ru1��
2�����"O`���͎�@1��r���B1���v"O�q;w,��I�2�0��R37�Hy"Or��0.	�G.�&�^�T�@�"O�:0jC#4N���l^�ߘ�X�"O`XG,��I�m9�	׬�\��G"O>��g�?�:�QI\�pҜ!�""O*��ʹ6��}���S����"O��r#�
�aܾ�Ir	���p�"O��+���V*n|0�mп9��X�4"Ox�0���?�2�+�$;p PD"O���3	Ö<R=k�h@�.,.��"O�4�r�388x覈��""O��ƃJ'Un|��
��@f"O�`i�J�
.��|��!�k�X	��"O� ��Љ1r�L�j)G���E"O΀�+@�#���瘭clBMQ�"O
Հ�J��0����h�9m]�A2��}>�$ �<٬�X�F�������O�=E�@��Ij��I$J£:��ъ`e�?(!�D]��ܜ{�
E�%�D���@�/b�|��'kD} �!����0�Ă�+�jh[	�'^2����B�\��-��@Y�'��pZ�`��f����
� ޱ��'5��!d\�D�x�x�k��z:��'�\��F��	W�`Ca�8EP�z
�'��A�S^jqp��8�C	���y��ږ,ɤ�0We��$��a�
D���>1�O��+��0`K���dͻ6E
L��"O�h`�C_��PlʠEҌu(8,�"O�M���T1%� :PN�".�8`"O� yԅ1R�d���L[�l�N�jW"O,��閅B�8�t��j�Б�"O �,�u�dl!0��9\i�<��"O���GE�qy�9t�(��+v"OV���A]UU���IG�P̀=�����@��,�5[p�EC�Yn ��q�>D��C�4:Jd�X��9R�[ !0D���āW�n�HY�'��[����"D�,X�	Q�*��q�E�Pj�<#2�<y
�(x,��!EZ(Z�x�E/�c_����=�䁢�c�}��0n�.7��?q�b!̱[3�
�{�����/!wq" ��b����S��u�.�aGb�\'tE�ȓ;I�$�ׂ̦vc���R.M�/�8���(���2A$��3!b�A�Y*��]����$�7~J�����O�~Նȓ+zR�S�]8i\<Pc7�ǧ��ȓ[)��g�R�cZ|�"��"o˺����Je2�΁�do萲%A̟jt�l�'�a~2��+���̅�x��C�ާ�yR�m8��\u��D�yr쒶� (c� � �X�c�-�6�yr��D�
��A?��#�R:�yr����1	'O-�  � �ǂ�y�c����3�W�#d|u��nA��>1�O�X���ױ>N�%����ٺ�'mў"~B1��.|�P�A�+����寐�yIF0fGv�"�
����еJ���y�mەv`!�MڤvoP�xU��y��ނ�:�y@�P8��eB�6�y�$M�Qy��q
Լ~�FXE���yR����@��cU1g�əW��?щ��S�j^�3�� ~/�!+vC��%�=�ȓݚ�H�(P�R��
S��;
GtĆȓZ ���^n�Err)�;*�.؅�F�R�*s-ۜVex����K"=���g~b$\;�i�ILlY� �?q���T�$�kjʝ#�����F�{f�مȓ
���(�l����� ��U�h�Hv�׮,�ѓ!�F�^�����W�����5�V�oX�a��$8
�'n�)3FL�ލw��'��}�	�'2��p1�U��8$�Ɂ2�$	�'7z��$�}4m��nK�|-�͢K>����'u1O�`�vLߑ:N�J5�R�K�*�(��	`�Ow�l���<�d�Rگs加 ���!���*� د3\Pe�֓�� {�"O$�RvhB/�!:�B��pv��""O� �yó`�!����b�*p��;A"O�M��^bƠd����9T��廦"O��P��v/d� �0^�j�:�"O�2��
WXJ�i��G�k��uYC��~�OP�H3���:B���h�Lދa���D�vFp��9� \�sP�q!�T�H�mcG"־-������Ca!�D�#$x�&D�4�j�����!�$CPI�r�S4[n�kc+0W�!��;i�V�0T�wS.di� i��{��חaI�l�T��zZ`���'(�'Ca|2BӍ
�6�h����B�O��yҭ�0.���ffD�c���`u
H��hO"��D�! ���@��M"!n� di�6
!�dK9'�x�2�%�,	>��iZ^!� "eVy��T�_���0f�1F�}�,�'���p�ApI�!P���)��0<5gF0]�p����C�kx0��D��hO�?`b��)��K����+�'wgH@��/6��S&ǜw�{3B
�6��ݗ'Qa~�\ j�6�I�^�njD$ָ�y�O��j*�1���޹(�H�I7�F��yrlј,+�p���q'�P�F�T��y���7s��Au�/p�ҹ*ǅ�hO���ıs)�U��(L �AbFn��8��O��=���ḇ�B�+�<�aaC�62w��U"O��+��L>_����/�^���P"O�8���OV��	�v�O&n^��� "O��J%(�8}�=� �G�tR`�[�"O���*[?D���J�1.�b6"O��1�V��P�#J�	M�"	�"OT6� �V|����E�L916l�<	I>�N~���`�=4�xA���C���@$-��y���(��a��P�Kצ\�&@�,�y�o�(�i2��z����ȂN1D���##	�_�`	qK�@G���6T��Kv #L��UJ�A��pJv"OpJ�k��c�^��g-+_��� �"O�x����O�r�*���I��"O2�[䭗�F� y�C-f�nm0�|�'��L25� %��$� �9)�t(s�'B(E"�jѿ-#�5x��j �Q�'>�@yBI�t�*$A'K��_�$��''��j���<���F-ۯI%0���'��U@��4��ږdH&p�*1�*O��7�)ʧ	�.��7�]�#\q�D
\ƦX��p�j<����Q�x3���+s<��ȓ�J%���߳
n����� v4�ȓP�P��GL#u>h馠O�P�.���B� Q(헾~��`2���p��ȓ|�)��� d/e �n/wF�@�ȓs*asa��+�p�G�/D<��'�ў�|
��K�(T\9Yb�8f[r1q�FAd�<a�H�$h�@��qJQ	#ۦ� rBDW�<)��L�
��L�"	��
�SO�<��iPl� �����d��Iyb��P�<q��(J8�X�j���e2f˘M�<!�f��m�p��bL�>c~�s���K�<Y#�ދ�Z�b���\l����ly��'52�|��ˢ8���8�+S��7�O�U�!�dļ��\)���du���XA��'Eў�>�r�$Q� mn�ʣ�W{+�<��/ړ�0|�c.ђ.����υP����^�<QWI�:� �T���j���Q���Y�<� ^��v�
C��SDɌ<�x�h2�'�󤟊wj0	�E:�@%HD�d[!�N>y��!ȭ(�t�HɊj!�Dťq��٢&��;4:\2	T�E>ў���S!��U.�Y?�����<����hO�镽H��}�`�V�|���@�`ՂH�!��%2,��ƭ��O�xS�NZ��!��I4��rM�<P�D d
8�!�D ��(�B���z������!���fa��c`@��Z�NW��!���)<tp�1� ��~�B�c��Z4%!��P>騰�M��z�OW�	o!�dս2�@�QF�
��z�섾ZO!��?�HL��'uF�� +$,@!���(��t,[/s������7mI!�d4Vn�$��8Qflu�f	V�*�!��$%/��A헧!X�����I�	r��Z����䜬=Kl�96%�)vv���]]!�Ą�7O(QF�_�G@@,sM0i!�$�T�\	��^�+�����X��!�D
�m��h��aZ�:�ǘO!�$��;�`:�,�}b�Z0TJ!�d����x"��c�|ԚD$���!�Dݿw"F\�B+l��#dcK)^�!�dY0r2��AS���,�`B�K�1�!����8��%�.��=Q�Ã*!�$ط#�RDKQ�H�j�"��։۞v"!򄌍wb��Q���ikj=�sH�.�!������	FG�U��E8��y��'1O@���5���h��V�H��"O�I�"�F-]��=��L�vq��I!"O�A[�	' �L��J��^1��"OTE�B_�Y'�P���@�d̾1��"O���1G�8K;�љ7��){ƞaY1"Ob�Jg�W4���	���/��yE"OD���-Y({�Pg���h��8�"O�-�v��L���l�%4���@"O6�bV��]j�W��?6�
��V"Oა��v^B�:���cq(�ʳ"O���'� ��G�<X�@��"O������e�������4��p"O�P���[AҨxd��a��,�R"O]I KW��Ѫ�F�Jӈ�P�"O��3�`�^�csş�nҖHs�"O�����p�x-SFą�.m�-�%"Oj$�V
G:㎙�D_3GZ� F�$!LO��ʄ)ϪG:�03��1�؀ZF"O�|�s���"��'I	Lx�$aB"O�dp�É%�h�!!��Hh2"Ov�H'��] �Jr��7�.���"O��[�jI�4U�`���Ñ�ܥڗ"O�%8e G�ahf��` �Y�����'��d�o����I��8�q���.�!�dN-A�p��%PS�h��]�w�!�I6Jh������t2��Jc��z�!�$ã3����S��81��r�"�3!�Ş}��agO2R���܀E!�dcF�pN��qα���I#v!�D��_�n����n{иEf�~�!��v�h� ���/jx�HT!�d�2c��\�vfX�w��[scC�g#!�$N�t\�A��Ib�^�HB�	:`
~�k�LAE���c�#*;2B䉺pz�5Z� �#4\�؉�� �C�)�  [Ώ4^��C���J��"Oֈ���DJ�d0����`�E"O����P�qAG��Uޮ�z�"OT�5oL� ��9ՀPTrfX�C"OlezB.��PJ�+�j�p~�x!"Or�r�F�?W�V�Y�E�<`�"OU��*C6"<Aك��)��j�"O�IҠ,0?j @	&LX�SV!Q�"O��u
�
sn��נFU
2�1�"O z�E��1�,�m�=C��"O��S�����Y��K������"O�Iӯ���|٩V
�(^��p�"Oz,ڣ�H$�X���4���KF"ODȁ�@�YqH� N�h��"O���I̦'�xTz����4��"Ox��A�Q�B:T��`Gi���T"O��0A��.�\d+ n��KXL<��"O0iZ��A��Bˍ^]�K"O���:v� �x�K���HY�q"OXX���/e�iB���:�dГ"O��f(\5вt �&D3)�H��"OdD���_f�8'�2%T �"OYP!�.f�*��@�(eIt"O��A��S7:���UN�Զ	�*Ov����*$ylp��
G�X60Q�'l��Q$'ܲ5�Nɶh���v��'��+'O��i�}񘘋�'ZโT䎧X��+b]�EV\��'@� ��.@���� ��Kzt}�'h����пC���)��2E>��	�'�VY�Ťܟf��iWO����U:	�'̐�×�γy:��ʶʒL��'�>�c�i@�4����`��d� ��'���)�ό�j.�(3���0D9I�'�:�*2ʃ/0;��%�
�
�'��H厙���E�2(�.X3�u;�'���򌞷M�d��$�U��'�abBgLb�~��D�:�2x��'�lq���s.��Q�J`�z�8�'�x�*��(� �DfJ�OF���':�p`d!�1���Z�}�J��'�����ۥ:~�,9�!�,x����'��1�1 ɳD�t�E�٩q	�:�'ڎ+�䞨	�9��R3
����';�0�R�T�Q6�ȥ"(^ ��'�J�5(�J]R�)%T�'����';�c[�IQ�Ł+�($+
�'W�i�C(�2?F���À۹՛	�'h���HܪG��(i�D�4��a��'c:��`@1v�8��6L� wL4���'u�A��L�"����i�H��d.�#9lT2���x�$����0(K���ȓ*��x�%�1L���q�ß7z��;��x�Ǯ,FP�# <�-���\DBDE�5p |� ��J����ȓ^�ޘ����Q�Y����c@ m���.u �jtφP����CGu��Y�(�i�J�#zHp�U8e��T�ȓ�܅���H�k��X��36.X�ȓM���2cD��V@��BB�P(�E�ȓ]�� �cp bR`O�2K�m�ȓ~�$�B`�l��U��)�F�ܠ�ȓ9�j���
��>�!�E#���ȓ|���"�HE~
er��G�\0�Ć�S�? Z��<_����ƇI\�$�7"O��#�h^,��&��;?��"O��g�\�	oh�de�
X�B\)�"O�;*J�:��H��ź`F`�C""O`���#� � @��c6>F|�u"O����NĶ<w�<S`l��'$M*b"O�]h�d�N�^e1��«pjh}A�"OL����38���d�=K�ʰ�3"O
��t��Xo��6�Y7o��p�"O$���L1V��1��L��E���f"O��0b��&)�,q��ů|T�"On�ñH��7U�%�V(B1|��8�"OX��DD� �"5�b�Q��
aI�"O�T�EҶ^ج�Y��J�z� 5A�"Ol�C�_w��C�	�8����"O�-�Ө�.��y��R�A�d�x�"O@|��*Y�qmjaA��Ntv!�'"O��kuK�%
"|)�)M�"b<�z�"O�YCt��"6zX��"�ظ�f�J&"O2�qe�͇��qL�2�T��"O�quj�4HXz�am�06j��K�"O(��Bf�uӠ���+�OY�[D"Ot�q��.D'T!���Ã_P�P�"Or�HE�"u�����C��&6���"OI��!�4pJ��k�U�5N���"O�yx��^0�*��'��6"ORXx�h¶(��5�iW�'Z̀�"OL=ҴF�)%)6	ဃ�M�2�s"O.�f�L��@4�`(��16OZ����L�������]���i'D�L��F��hG�����ϕuTU[��'D�t��o�,i��L�ju:��1D��`��g�-w �j���-D��x#N�%z�M�Q	�d���C�e+D���׭��D�p�R�T�W��XzT�,D�x�r$M��D��үG [�D�Y"�5�O�I 0vƨ�Ɲ�,!BȖ	�*˓�?Q	�1�`	�KL&^1\���`����,�ެArE \�T�!%��)�`\��1V�� &���*�ёSJN*[(�|�ȓj"���	C#Y���u��g ��CG��J��A�B��Q�K��ȓ9�~�e²	�u� ��	vp��S���A)�C��u������!��Y�Pe�,�Hp�V�C�nN�Նȓz��@{�^2AS�`s��!]�2�ȓ��m䌜 	ՠ��1�3Q	jȅȓ!�8���k#�����O�:,����p|��I���@Q�m!�o���4��ȓT�
�
��_�0���G�,Z�T�ȓ	;�0p��W(�\p���/Y�r4�ȓ2q*D��,ɝLF-8�l3V��ȓL��h�����}[��[ǣD��X!��d)���a���Z{�c�@�+�:���"8�K�"oJ����^�t����  L=��'s�e[\i��d�""Oj�1��Lc̽YP4S�:A� �|�)�ӆ"�;�&Tx�B�{FFm��B�49F:��Qf�=�����h�C�ɨ��-+��V&CwBpʗ-%G�C䉫X�H	���/m|ر���ֱ�C�	 H�l ec�9A��u �!�C��8�  �"�.n4���ˆ 6C�I47Β�5��-�,d5$M/ Y0C�)� p���z��$b����7P����"OPKtO�%�\Р��G��H�`"OPR���)�zQ3��.]¼�"O&e
V��X��DB���M��]�B"O�0��@�^�!��i113�	q"O�i 5e�*o�6i�"�P�j�H<��"O��AK�*g>����r�f�c�"O�l�7�r������'q>�P0"O���7D��R*hy(R 	&E2�Ps�"O8������Ud��
��ɶ> Э`W"On�%��T��"D��m�T�"O�8��ėo��4��R/^$`"O�tF�N�N��^43I��c��'�R�'w�dǱO��<��Է/��$��cK!���2����^<>�j�2�"F&��h��D�֦N�z%@P$�5�\�bvn;D�`���l������?`�3�:D�x#�	�$j#�Ȥ*[�P"T�6D���Rg�$}���8�'��~��5y�"D�h��x^ݛ��=-t���* |O���yR�H�F)���lD/Y�\��'�y�@��,@(\��>N������8���0>aP0h�t<����%"Nusq�WK�<	'��LnQ
�iΧP?4�c�IS�<�����Ҽk� �'�pc���O�<	ć̐A}Fx��͑]V����)�b�<I7��W���	RDGh�F�r�]��D��ݟ�Nh`��)S���m�C� )�m�ȓ(�(�N	�4��T� �$�֭�ȓxp�a�FD�e����S,��=񈬅ȓ�,,�'@,o�:���a�#����"-�yIQgO�-~���1d$S���m;�@���S�N!xL�w��1��a���� �K2V;K�5J�p-	T .D�X8Ą��l���#cO19���2S D��1�\�I�@���L��q��K=D�|s	��=n�0����2����W ;D��آ%^
�­���QD���p.D�(a��A8(���ѸX@t5b	*D����S	-k����O/GGX�E�:D�@{G"�!}K
5����kEDe�D�9D����(
B��)KV�v�"F�4D����\ג`I,W�@�a5�p�!��Z�@BVAI���(q'���{r!�'F���#�0*ʵꇍ�s8!��NR�\�Cw�K$T$�A�4�B<{�!�D�nµ9fe3<`�ÅH�!�� \���/Z�)r�IƝtw!�����i3�\>X�~� C	\�S!���)Vtvh�E�7l�~��2	��Py����KC�*�5*�(�[��E.�y�n^2q�*���dF�M���L��y�3LD��Xx��r�E��yBn]0xP��3��x�Ը��\�y��I�1��X`��J[(Щ��D��yr/�<JՆe�n˯Y��X���
����<Y���~��ar�JB癰�`�Ȱ��_�<�#@�lP>�c�&�-u�A�3/EZ�<Y")�]��P��M'G�B�[�PS�<�1G�2S�AC$��3BiC�%�h�<���`��f�T��kŋhh<ѱ�N�mc���Bξ�t����H��x�hY��^Mk���/3���&��(8Q!� 6#��4�9:�E��=A�!�� ��'��9`�bVu�2` �"OL=�pē&shB��t��a�b���"O>U ���*U"B��'�"�b"ON��GČ�>{#�Ph��'i�
U���lJ6A�_5����!]�مƓGȊ������V8*���H$�"��'��Q��o
�c�*tS&E"o�+�Y�<��=I��!1�˩EXn��P��U�<��"	�4	xnG&Rޢ���+�U�<��������,��s���T�<��	U�D(<qm�$+�T)@��j���Q��J��,"ڝboĒ:X*ɇ�i��T�)7��KpDՏV�|�Gr��8C�py��]�7�	h�J��fu��O�����fL<��N6jhx�A���y¯�$%J�I4���d\PAhq�Α�y&��Xp%n��I�(	[�.��y��%`6�=U��D�D㇫��yb���T��"Êj<���OϦ�yR�?�h���L@�]�,-x����y�.rP���Ѥ*'� !�?����"㖴��+ �X"��ŽyOzu�ȓ/�ʃ ���0 �;b��8�ȓl��;��ϘT�t���k��c�
��ȓ�0I���rԪᲠ��8����ȓ;E$X
Ŋ�mS0���i8�'� F{��4Kq����LT�0�Ö�U��y�l�K��0�.��L�1&a��ybD�	����6o�<�h�I�����y2��r����7�����L�y��
_)|�Q�>�� ��D\��y�G����  ]�g��늎�yR W2�ͻq
[ 1���<-�!�ߖ|v����R�<��$@;I��y��	,��÷	�$[;*S&!����C�	�]t�M�G4�@x���G(C�I<|�l�#����-����CƄKP�B�ɮ8���Dl��.Mtm�Bh��]{PB�I�U�Q� ��ua�K��W)<B�	��ftɁىY�ڙ���vc&��ȓP?jT��)��P� +$ȥ�ȓ`DqAC==���vG��T+��ȓFp`a᠁��W���G���~�ju�ȓl	�H�$~n�k��ډl�|q�����٤���tE��	��1\5��0�x����ʩgs&�R@�U��x�����B�I�g��jG%N�w2����D2����mHpl5��b��(�Q��"OdIR�ν_d�P��CR���B��'��"��b̛�&�gw|0���>L^!�D�L�zl��9xj"ٹ�(�8c!�K2�f�sbf�"YE��fǴW!���C^\��UK@ra��E&7�!�d\Gľh�AɄ�o&$���<�!�$�0`R|��J�y�DY���-�!�dάY��-PԀ+�q�7H@%�IM��8�5��X
M��9��$Ӥ"D���ф�%U*v$�K�0��8�G"D��Cab�OPM�#JG6�z�!�n=D�p�T?-iJ���._�R豆<D��q�	ɾa%��xq"�=aCFYc��;��z��̋#�%K�lHdÄ�p�F�8ړ�0|"�g*^$y�dʈQr 3�ALC�<�ƯA��8+��S���\ �.f�<� �ٲ����P��0T��"OJ���$��GfY�Z��\�"ORt��y�Ӈ� D����1"O>Ȩ�Y9	A��
AaT(B���r"O*}�aa��C�F0���G�bD
E"Of���&
hl]�p/��~��V�\����KY�U����@����FN����?1��	���ZV�.#���[���5!�Ć�[��0#Eo��-��Q�/M	3!�$ͷY�3G��k�m2Q蝖V5!���A��<	�nʩW��(7��&B�{b�dW�;����0EQ Q��P��eѸ&!�¦�8��&�e3VuXi�k�̟Ї�j�L���)9渺�/�
)���$��G{�����7V��e!��0CR1��	�+�y���j�D!�����5 �p�I��y�@��,���T�vL�h���[��yU�j�
��[�]J��7J����<���$�3�R0*�V?��yBF͈.!Y!�R#>f���vG��k��E�QK� �!���h4Y��`1" ��#��3���)�'4��e"�;bp��:F"�73@����'ل`+�M@�LJ� �fI$T�I��';HY;֍�&E�Hp2B��j��}�'�
�ذEۖ�D$��xA�$��'?�@�W�T4��Q�S�)r��'w��ElK�~�v4���/&1���'tH�Ā�0�PBuj���#n�<�d�R��ZAb�/�W4
5��g�<�SS�Sb$Mq�&��v���B�g�<a委'tl}��F�� �+6�Ed�<���Q�"�(M�aɽ2�ԴۂMSf�<)gi�&~]��!7�Q2<op�CgE�e��v���O�F-�m"j+ؤ�Š�li�eS	�'Ӑ�Pw	>#�4��t�X�b)l��	�'5��1���3�N�!�&`�`��'c��'t)4=[�,���i
�'a��7�R�	ř2Ǚ8it&�s	�'�h�ңm@'H�L�B2��b���Z	�':\�퉨^���{�g�T8.��(O6�=E���m��9y � �`��̹���yB��5NQ	�+P�	@���)ژ�hO������`B�d��*���'�a�!�D�$X�$
�`R�鸬���ؗ Y!�$[ W�rX9��"؞��ⅎ�!�D�)T۬�Rƅ�,;[���b��Y�!�$��R��i�CΘ5PR:�0�O#J�!�.P�@+Y��$�w� .a3�'�a|��M!ٖ�A��f������ �?�)Or��D��
�x���Ֆ/Ch�I���d�!��ݵV?|��!O
/#>�s�3 �!�Z)��M�#M F�WEڦ(�!�ċ�=�N��G�V Q�_]f!�$��"����ʎ'
pb7��1B+�O�=��x �������9�	��F���(D�XQg	ٜ����C
\�ia�8D��{��g��8��y� 1��"6D�0r M�$*����'�0�(@�3D��I1痈�p�&I
� !$�?D����E�x��Eh�8\���%0D�8���J �@@rg��#�, �.D���Id��@{���2֬��"9D��[��.z�,�f����V��O�C�əs�h�v�_�2϶`�	�S�<C�)� �����Y�N�h��Z�l4�PQR"O1�N�)+��f�ëwu��(v"O�r�Q,gq�4rvb�C���"O�<���7!��ԛp"�~�-��"O:���/
�D�t����Thi��Z�"O����@�8L������P;c�zH*�"O�����b�Ex4�	�P�V1�F"Oh�9�m��^h�p��2	��-s�"Oܨ�@�:�Ơ"-�t�aC"O�	q�̝�7�&�ځ�f�^-Ȃ"O(�)#l
T�80�Y�C��
7O���� թP��s��-_D�z�H&D�쁓O�r>Rlb5��<E��p��#D���
 7@��9�vI�:6�`��"D���$�M]H� �$��-\����?D���ЛO�t���J���9!�=D�<9 ��Tz~i)�C+#���4n<D�H; �	&����m�09�E3�k:ړ�0|��/�0�<��%5�NղD�z�<	fӄ!`q�eaU��Z��t�<�Q�A��h�W��E�(����s�<�'C�%azLB�LBd�JKq�<��ߋO�LԚ�f��
��$��ME�<��C�T0|����$6��	���C�<�3/��:DJ�h
�.1��F��A�<YRm�>3!�![G	�,ߜ��PB�<a�Sz���so��E4��"�B�h�<y�G(3Z��
�"nU$�b�<����~�$��G��m�b�a�^�<Y��X�c&r��E�Y*ɲeOM[�<�p/�2 MF�P�g��6HR���*�Z�<��ד
yH���D
�2*`�ѲCZ�<	p�B(u�f �2$ 9�f���bUq�<�ÍO2D�� ��7Ń�A�i�<�g@�)�`���)�2+ت��e�<Y��C�|B����V�(�dAH�<�ǃ��xz�l�2b�|1@/�i�<)$�6�rQ��T�`�NH�v#��<�%�ė	����$AA &2����o~�<���G	%X`,JE�'(x�@H�FU�<!U��9
�<��!CEH����_y�<����d+��)p��T  9����q�<�H���Fa�H�r����
Mk�<	#) G�I��Ȁ%=�ɐ��b�<��� 25�`�3 ����H[�<�e��]P~t�ԫ���9�l�<���)\!V�0�*��c<��h��n�<� ѭL>H�j&a޼?�.<p% U�<)S�@ Sr@Mѣ�H	f�34�R�<Ɇ`̢&Dt%1B`�j�H�+P,�O�<a�B&��J!��x����NS�<�`bO؜�sm_�ZTT%�'t�<9P��z���a7�T��9�D�s�<��ʋ���T�@_=Wex���q�<Y
��Z��%
�;;�m���n�<1NQ�wR0��#�33��!�BD�<��K�;~�r\(	3ń_�,f|��M�؄��"T�n���D�CZ�Ʌȓ"�D���G��0�%��a�VԄȓn���"��
0��`�Um�x4��5����H*
!�U��2𦹅ȓcPXM�Ƀ�*��C�>]/p�ȓ=���jbhZ0UL��bB�I��NL��.Y,�/)�M��H�/a�}-!��  ����D�i캀�uJ�I����T"OY@�"�#T�@ô.V�J���{D"O|H�`�.i��,Nw��}p"Oxh���\�S� �J�" �"1"Od)4��TO��2l��U�ؠ�"OhV�2(T�2aG��e!\!��VC�<!c�6v��4ف畱CF�$�o|�<��#�5��Bc�0C��
%h_x�<�C�(@�\�łP��V(�SIUu�<96DS�5Rp��iO>4�vHe�v�<�Ǫ�T<����=`��Eep�<i�kţ'��C��ɱJ��dAg��o�<���9 2(�)�� -r`H��i�<�˜�
�Bm��Ɠ{�d��
�i�<)թ��DJ�d36�ȕ$��m:S�~�<�)Wh ����I;~��A7�Xw�<�W��hbf�4Q�d@�f�<�R7j�2�*�4o 2%ۦ�t�<s��%��䑣�\�VohXJ�	Cr�<�%�" /܁"�� �^�:U�o�<qa떼���Z`M�r����	�@�<	��@(�$�"KR�� `�E�<I��.H~.t�ҏ]E`�@B$FC�<1C��*Xt�Z�`T m:�L0�t�<I���o������:s���k���F�<�Ʃ٘3�ԃ� �a�p��4 �Y�<!�AV�7l�z�/FOy��!��K�<I�+�
=v��"���*����Jc�<�sL<q�-��M�@B�!�ō�F�<�։Å[�]�`��!EDl���<9G�[/��t�M�8b�T
�A�<��iڻeF>E
 @OZ,�y�%X�<9 Ϙ
GD�P���1�8����~�<�W���&�2L��IR��OA�<�t��3\�xXg7J4����Q@�<AR+�p�x5���/�PAa�C��9VL�ْlЪ^��P0@@(��B�	� v+a���`������B�	�H�&t���:�\EK&+нt{�B�	>H�`�*���liF�%�#BZ,C�ɑ8�P��@a��)gԉ��K>
{�B�	�e��FI��-5��b���.D�B�I�k�B]K��'�D,S��@�=bJC�I<e��J�G��r�TyV�^�6C�I4	�8�Y�Eb,E ����`8.C�ɏnȢ�MVi���ի�<z�B�	&<3�	�D�A�4q���f�%I,C䉓<����.B��8j��D�p��C䉕!y(@�D�\m�A��!$�C��S�@�R��W��5�s�J��C�<!e����iA�F�t���.U^�$C�	�z� 5���=fYF 5�6��B�I�_>-2���4�$�Ძ��d7�B��5[��i[@�&O�����O��B�/I��Ae�U�T���C�pm�B�ɼw�q/�!��4��V�bJC�-^��ar`$>j��p�<�C�	,��1�rjΌ���)S�[ �C䉊`��i��Nw������}�dB�	X�� P��Վ0?�@�aDPY�.B䉾P@D�0��C=����ϐ8H�B�ɯb��P�cB�C��ݸG��})8C�I-H#pk!K�e-x���ɒ])�B��-�(�ӆ�H29~��#�'ƒ{޶B�)� �DML�2L��4��F�ZQ�"O�\c��CM��Y��M�@�(�!�"O���`ūN�qǔ�Y�d���"OYh��'g������Q�ZR�"O���n gs"ґ	��Q�B"O����. r��b���n%��"OvAc�a�'�Zu�)R�8����u"O�`9Շ�;o'","1��f����"O��r1k�*.���R�]�2����"O��ef�)�)��,]�P}�"O�%��F?�j]�*fM�"O��ʣ��x�ԅ��E�<|'�%�C"O"�yr�:3�ssD�K�
�"OB䋡
,�r��Ud�d3f9��"O��
�`��6ͺ��%�_:��"Ovkf�]�^Q�@�O�,�8��"O �S�$B�5�ڜ�.�U^I%"O����'��e��� !��!��S2"O����]�v�^xZ�Ʌ��<���"O��*@G�D:�z�F�TC8�x "Oj����/l:l@��-��B1"O��`s%@w:v��-\+2�c"Or +��b�h��T� �p�"OV�S�#W.6&`2��!wk�!��"O֡!W��3����&GA
�õ"O ,I6��]O�bV�b8R�Y�"Oz������,(!!�%E6`�X�"O�[�I�	�v �Ra�m�`u��"OZ��6`�GZ6j�̔Ȑ�"OУa�ܰB��Q�N��t0D�,�amF�0��Y�a�\R9�s3�3D��	Kq�\[�o�� �U+V 1D��[ǦԄzb�@G���+��c�#D������-U��H�`�}���UJ=D��A3�
�K�Tao�#��� �@1D����JQ!68��k�N�Cz�(Iҍ/D���3FH�f��2�OB����C9D�p2�f	"��lC��d@�LH1�7D���3╳h�`�GI�=	�x�i��6T��@�ם��	j$aC-'@T!�"O�I��'�<G
�9' �8Or�T	u"Ob݈ŭ8Bj.����V,xw�Di�"O}�e�C�xia��_d�H�a "OfI1�''rg�p��1{2m��"O�U�"fW�Y���ANN�]��P��"O�	�H�7,|��"�+Ⱥ��X�6"O��j�гesDy�)���d��"O���B	H7 ,p36�̇kqX�0"OP9`��M91���M:j�x��$"OX�@u��V6>%�FAԮW�Ј�ȓe�C6$�	�0�� $  ���`�l�'舾X":ɳ��	�|��q��M���1���J�8�	Ȝ:��ȓ ���jAl�F<�.�&2N9�ȓe�>��I�!��9�A/�����s�`<���ƬF��tj >P�2�O��=�"�h�5Zu()b��I4�셃g.GU�<�J�ITT��'�#��a#�g�T�<����Z����	��rQp�����QX�$Ey�&�@1��ޫYH J�m��y��߸g_�!�ł*NQ>5�w�N�����hO��~D0g�O�+∢�#5�Θ��'ֱOD\����t�ֱ�B��ۜ�@&"O��q��6fF�d:�#O�V]�"O� ����LN$Y}�4��
�-6N�ˣ�i��d��:�aB���g�.�y�A�>t��D=�$�<��'Ή'ܛ��S�*�VD
t��(����`	ϵ�yrn��:��XU(z�bHX`�2�p<���$��0Ex���O�K�P�@\(A�a~*p?9��CԔ���Z�S&*1I��^{�<Ql�� y^�0���&+r[�5�t�<Y"�=B��D�B���pX���x�<afI67	�U{�*��� ��d �. �`r����OZmrc�U�5�YqTƕ�U
�i��"OL�@l�R��!��G�j�� J�O>ꓧ�=A�A�Ha
� pdM�%H��^z�|�@	6` �	`ܼ��G�_lP�*e�6+����脴u*|�փ�(+��d�� *D�(�A
�*�:�a�G�<{��)Ԋh�֣=E�ܴ	�#3��/�4H�!�O�p����hO��6�$o���JPlH�/FF����a�0��e"OԨ��J5� a:%��;��t���d!�S�'x�$�H��=Љ�����E'2���II?q�GXy<"4F��{hh���J��0=�5E՗s�1���J�Q�R�2�MJ�'n"�}���%?�*�a�T�x
��zbJ��6(����^����b���T��L�r �6C��R�'w�D$/�*MZ5�D#�pj��
��C�I�f����-ż ���T�	pؾ�'5a}(ۙ8�@qy��ԅr��Q�&��-�y2�K�~��h�G
�9=v-�f����y�*�����j�%2kP����\,�y��\=D�t�d+^tlR'����ynа&&(rm
�?qH�[���7�y"K��u9�5r+�01��,x%�A��ynQ�96|��eT�]�0Hj�R�y""W��XDi�nR�JCDe�D�� �y�E�/E�����o�"Fj��1���y�C�����S��l�)�A���x��|f�����~�(y�F�a�tB�I3.��q�S��;��U	�rf�B�M�ё�ۃ4Ï��#��B䉦V,@A�e����*Q!�h��gN2�IZ�&&y���Śjd��ȓ|\j�zUc�� ��ÂM/J^!��i�Ty�&$��XR\k�LIh)8T�� ��xۣ��)+ph�3�))[P�ȓU���J�ى��0�g�#v���ȓK,��sQ"A�r��)񁘞.{���<��ƥG�Fw�������X��>1�a�ڔ|!aCY�E�����u�{0�RD�A#XP�=�ȓ�J��F�+�0m���F�q�L��ȓ��$�����$�F���5�4�ȓ&[@{�@�d�Fa�m��O�@��U��8�6`�0Lo�� �%_�,*�`�ȓ*B��e�\������G�n��̄ȓ�$A���[ 	)2���J�>���ȓy�hl����2T�Eha�_�G1���N_`T!�A
!L�> �]9R��؆ȓ#�b c�*M�'�L�cHQ�_[��ȓ"��)ɇE|�P5��'Pr1�ȓLP�lx�h �Tm�`Z�j\�+�n�ȓe��D�!�)�A�%bC0$8���]2T�0eF Q[f���O�iC��ȓ[��1#�O�+�,����ap��ȓ|%�#o��@7��OP�ؚy�ȓ+z��Ą�#t����I^�s����S�? �t+���<�p�p%��B:� �"O���f�Z�f��Q2���;Y��K�"OR �7�O.
�"��(؆a�~܀"O�Ej�`�l��D�ֆž j�"OH�X%NR�)j�̛�c�d�#"O��AF���^��+�aTp(�"O�L�F��4J^T��K@�c=܉B#"O�@�gMǖq�R	N$
+:a:"O�,R&- 4s�;�(�$&�M�V"Ozɱ5�\�#��X:5I�b�<���8LOfaj�gZ��Ⴂ���s�x\�"O`�SF!�p1�8��c����D"O��S�L�TW� M��%�@u{��'n�tS��(x�lmI��X� ���I�&D���T�.nn�"�)�8D��=�v):<O�#<9T�H�^Xa�u� �_���ZRn�[�<q���f�,2@˕�!F�	S��FX���0=� #Jc�R�e��R�<ݹ��S�<�F�_�8���W��*ߞ�Y磘ԟ ���s4r\��&�'E�5��WF���XW���f�� <���Ģ�*v),��t"O ̹�A��$&�a��#f}X��e�'lQ��cN�gvT����&x��$9`n!D�(�t��;�L-"#^�}�05Z��?D�l0Ъ�9I�
�w,������"D�@3�"��+�:��
Z>Fz��2'�+D��RǢЌ|v	�v k��R�#D�x	ύ(m��ԛǥƘ\r���"D��S'	�4,f�9TLƹu��%҇sӜz�)��)c�!��:A�þwG6����4D��*Rk��	֒ܪ����9��+�<�`�'���H�

��|]�f�]��~2&�Jb���#X q�� ��>a@�7�,}�i���=�T�'����`�S�0��j�Ö�b�]��'Ѫ��C�Ұ}�U��ݨRR���'�����añ�����F���������'
Ni�7 ���D�R��qO*��d�Ct
ر�"�1ώA�����5�a|�|B��9�KRTc�9:�J]�yB�9	Af4K�3H��ag����$�<����?�G�"'!�IG$P ��S��8D����� ?%��Cp'��y�HxK7D� b©�-݂=3�ˣY8�r!/7��G}��OP�?�X2A�:B,��S'���_�j]y A��0��I�*m���'�~����p�� D�꓁�'�Ӷ~�qO��@��M���j��j�\�$"OH@:����fE���7j
�K�<@a2�'�	f�S�O�.�h �.{+�`���>;�i�6�'Hў�0Q�@�}j��J�Ĝ1��0ɗ�s��Il��O�Ƀ���:��hƟ)��Y��'a�V��t��k\���
"�O>�8�9�B�OC�I&;CI��	Pu<H�c.�8��<�����'�6ţEڳ/�آ���!c5F!�ȓ_���X�&��EO�M2(M5��Iw��'��T?����TR�
�F	�6�d���@�eE!��P=�"uAt'(;�>�	�i�)�?��S���DAd���e�ȘQ�JE���[��!��r.)X��8��m�b&ٛ>�!��8#lq�Q�@.Q�8�ITlD�|�Q� D{*��$�0!�1b�RQ�`	E�F}pT"O�t����&�μ"k��*��E"W��I����r��>2�tH'�N�T]�ų�E��yz��(u��&z�`D�utp|�ȓ]�툓�0���b�.L��S�? ���O�F%�1��`�MRv��"O���%	�'1T\�+�/�� r �q"OPtz�k�w�tA��%?��yv"Oԫ��<>�m#�ݯ:r`�"OšAj�U�~�c�A )tQ04"Oj�
C.���T��/�	%̡�"O���ąoN�Q��X��r"O�=C5gp`����,G��(f"O�a�mѻVc���Ƥ�;#˲p*�*O�(!`KJ(Ь�ȑk�3�i��'b����G�"H<�!��ԃ5����'���K�V��!q*B�-yl�H�'r��A��^�0ODK /�#��ĉ�'�P�!�j�:T��nT�	2v�@�'��я���UlȢnn
]p
�'���aꛖw���g-?k��5I
�';8�"Ӆ>�vQW�V6��'��7�_"��m�1!�z���S�'\��r&�#d�X�PM�o� ���'��i����*StR��ܨ��'!R����M;(Zթ��D
��aQ�'U�e�S���E[*I˦"��}<�y�'_Nl����8��YK� _+(@.�
�'|Tĸ��*�\��ۥh���
�'�$|ktG�)4�@ذD�O�c��� �'Ć�tM�VJr�AA�آ_0n!z�'�,#�
�$9`H|����Q"P4c
�'$�ĸW��_��eP`�%z�hi	�'b2]CQMO�X�Q�G�ƿ~���C�'h�k���>�b�s'��/wL
Ȱ�'ؐ��&�@M8�H�lж���'`,y$d��v�*]���ʩ׎(���Ĕ8|�* bS+];gf��-�sV��d�*j�T��4��w�Q���N��y"�S�vF�y����6kf��y��D�b����J��D�`�@�y8i!j�r�,�:@vH����Й�ycD}����⋻FG��7)I�yr�I�q��i��V�GN�2׬��y��|�
1�Ǭ�2.�%��a��y"	9}H�b!L�j4�Y�����y�:*6�2���48Z�������y��� ��x�H�.`7D���Ԛ�yИ^����t��4��́B��yBh��X�L����/�p������yr�٩o� 0Yщ�Lި���ø�yү��F�])FI��D���Z�j�y�ፁI��p	�N��<2���'�I��yR��:�jH;�OG7[	"��s�I�y���;WvLԳ!uHLs���6�!�$�1%n���K�ر�$�%6�!�䊽(��'gE8�Fp����,�!�^Zd I��pn�\��H�e�!�D� `?�ݒp �,!YNx ��Z�e!���-V��ȉ�J��@�a��q�!���rxv��V ">����R� �!�D�h��*���&}�q�ͣq!�d!(�Vd*�D�N���B���a�!�$�5R����#&�U�d=� o�!򤋡:&�uwnX�Z�
,�����>�!���n&�.֢b�`H5�)�!�d /l|���"a|��r�L�'F!���W���+��� ��`��Z�< !��e;��gł�5bz<�'��m�!�d�a�ڝ��c��gf�)O�!�� ��pAnM�]�d�H�]�hzZa�"O��r�B�=��i��>}��3d"O"��P��?��u���H�hU��"O���¥�CN��#cì*����G����7u�����
=K(���l�,oO���u(��=�!�J1 ��%�g#� ���z��_#.f� +�
R�	#/bQ>˓�:��rbP"(m��	D��':2�!�ȓiJ����/g.0)�h���İp�j�0�Z��"�O�͛���T�� �Bճ�T�t�'�V�X�a�����-}�eGE0:�l,J&��A��ȓ9��S�"w�Ԉ���\�(��<���@	Z�0��C�:���ma��ѼQĨ]�/�u�H��ȓ2)����� _��Z�k\�-6�Jc��i�''Ppb��t��̔�',2�p@H�\Y�F�9D�d3<�kD�`�褘�!ڶ1'� �c�1DV�|�M�{K �y�BRf�Tv����0=aq��q�M�(��e�	�+���e�2j�"��Uo�9�fC�!N���rc�ӃH���B��Q�Tc��+���W�@ʔ���H�f�Җ�I4ƞ�X����!�j��"O��HA�T��hH�@Y�:�z%H�K�,N\s�,�~�����I9#ԈmA� V56�V�)B��81�C�ɣF�b� �S�C��q��8vyB9z��֙,���������E���6��C��=Mm�m�뉹n����R��CI� V>Z4v��"䶙��X�E�!��JM��|q���e��+��O�ek�!ʩ->,�s��%ʧAT�����2
M����K�E���ȓ0P�<��j= �H}sp&�^�$SeL1.�~�;b�4}��9Or!� ڞ\q�)r쟃F$�b�"Ov���2���!��V162Ƞ�4O8�`MMW�`�	�d.�g�ŊM����ǁO89��I�=pd��	A3��us�5]V�" ��H	���gl<D���2���1��Ȁ"�����U���=�_�б�b)-�H�м2�؋D4���Fk��}	W"O*-���3EXEP .��H�`�yt�iszs�(Ck�S��M�A�ٴ��yr�8&w���G|�<�u���|��,)6&\���Ug�z�<Aӫ���������Q±[��v�<�J��U��5aWË�w�L����m�<�G �(C�T�puˏ�J�0:�a_j�<ib�� b����ǅ��00��ȓ��y�+�?M����,���A��!����af�-��@p,M?nXB%�ȓo\v��� iw|4�& M\��ȓ?,T|�x�ӄ��'����}�j���1�
�pE�=E"���ȓ/s$�Ӏ�)~�kCȏ-Q��Յȓ|��t�w�;w,��1*K�L�,���:�5�`��R���A��,�lu��REvh{Q�L�C$!;� .xy��.¸)�À�5' z�R^�l��MFi�<��(W#.IJ�e΁,��lrv��}�<q�x���zdY�$�d�2)�~�<	�!��}� ��B�3��h��i�u�<���\��ƍ�/s��}S��q�<�����!
�i��+��7�Hi��"O�C�K�����a�%�� �ر��"OH�8B%
��UC&c��a[N0��"O��� �7|^�9c���%``}�#"OM�&=ِ 7
W�}p8R"O­����X}\� �Q�p@����"Ojq1 )K�[r8(��/�$9��C�"O�d�Y>6Z$9ӯ��"$�t�2"O�p��9pQ
��[0{"%��"O�5K��)y��t����G$ �%"O� &X��O�y��Mxգݶt����"O���p���@�?9��H �"Oxd`��܎t���逇Y���X7"O��"0��������2��Pc�"O����cN�fR��O�p�f�[�"O��	�o1�X�MƤF@�u�dP��j!H��a{�ÿ)Z(K��f\�I��
�9�p>A��U䦵��OJ-i�-��h2L�ef��C�	-k�a��V�IS�ݙg`��<�&�k3��6M1O$�{Ǎ7O{`��e���OsĘ��=M ����UӈY���ǔt�>��.�S
��0�.�+��	^=
7\��P���Y���(!�b�%�g}�LޮPl<���M&4��h3	����ٜi<����9��)�'HF�@(bjڰICȈ:$��5M:�n��	ADY+V�ȘR�h���)C8�����ݧNu:,)�!T���rA�k�D�(@���/��Od�B�"eǮd0R*uw�,*��	t�Ș"�ϡTlC4�O"°>1ֈ��B��E�f"Z)�p{!LN�3�hD�f�ٶm#��Md�Ÿ�M�h�Rhku��l,�c>!��Q�W�,�a��eiB�� 9�I�l���䘏8���f]9�C�&��s������	��75 �9�:C��-AA��1�>��'���k��Q�Cw|1��G�)q�O&	�C�;I5Ĝ O�"}:ցʫUD%���;G�`�fP�c����e� Ҁ�+ġ�k�3���$mz9�I֤q~�tva��f��'������Cg���Y���I[w:+� &h
b��լ��T�����X�2�^�
�֭^Ψ����Y�t%[���H�E����=P�v�H-v� ��)OB��!�X"`����
�v�0�A/4�	Y$ ~�A6$��Y@�)���X�6�џ�YԦ�
*b�|����mvP+��!~�����1X�* �F�$%�"�g���G�dQ� ����+hS0� ��?Q12�Zd�%?IaF�`�"|J���e�tY# nWx,j טT>��a�l��nU�G�ãux�A��dS�
�tap7�:W�PGF�:NV�$�@E��RG:3X�y����~2����8'ĵ��R�H\: �S��2,t���)�2;1@��m�D���?��N�?r�J���$#dp�3V唖*��gQ.�bY2��cVJ]�"	�z�j�M�!ax�E�׼k$�ĕ\cʌ8v䞿'�(�PT�Fx��@� E5BH�c,��"�ͻKq�h��gVqr!�&ӛ,�Ь�$�φyzby0w�Wd"��r΍{�'<<���
1[(|��e_��b���D � 8�����@�w#��[�擊:�(�c|���䜢�7M�gq�Yғa�b���sD�!O|̉6�\�;�R嚰�V�U�XX�·�i���냮T�l|�8È�S�hС[?IHs�ǫn	&�j��N5X�u�Ä:;J �p�P�g�^���iW(<1�CQ6 �v�S� � o,,�j�NY>F4
U[�HG�'�<���-S����Q��x�s��Ol��b������fe�Bw�e1'gRb��{b'pu(9q6(����b��߀I2`�@r�e��IG'.a�1��#�'��D�:;kt�@��':D4��y�ɍtH�e�g�|9X�XP����'	���R����$��[;2�b���*��)A/`L쫧o/�d�OY�t�"�$��x�4�J��f؞$�$�F.N64�z�e�)L�*��
�KxrԂģ*^��$H�O�j=���.O40�R�'� ��Jv����Y�
��ߣpޤuJ�E!D��r�F@"g��g˝G������Uh
���ۂ{���'�� �1�M��x���Ѷe\R� @�*�bޠ)���LV������8��P ���B�>$qԀ�
]J*�l!^f�pP&~}rIĒG�`�c� 1S�	
`��/�HO���ߴe�R��5��	q����r���RV:�	>j�x�X%�.��%��hDI�
"86��/9G���A����cю��>)`/�t7VК����̊E��%���Ay�E,8�� 왅]\ҽ(@�q;N�ʈy��h�ɒq&��؛U�J�ل�z��b3�ҋ���� 60գ��imfUj�!۠pμ�ObAR!��vĲ�0����y�σ���Y!si�mfx�;'iB�p>�1����� ���8��)��Z������ُr�6�'�d��CGư�>qB`��<⑞Ī��T�6���Y� J)P�z���k/O0���-�#RH�\}r�*�
��#܀�j�m�����<�h@�2$[�\��	���?�4$����s�Q���tNL�'�24�h
A?Y���Y첨O>���$�I�F�g����M�M�LC�	�j��H�u')fn,̩w�N�<�x�;@%[3��=��S�O:J�r�kK���*#m�d��'�f��Bb%�D�:�/�d���IK>1�oJe����d
V2D�$I �<�I�	�XW!�Ӝ)R��CǤ	bb�a?�$k�<a`���J����$���Ĕ`@��k�<���K��!JE��
�P$��JNo�<� �#Rϟ�!��8��E#u;�u�T"O�P	�ϯ"��=�d�N�����`"O�ڔ��=G&�5��n�d�pUK#"O�UK�g�rيA!BM �{��u! "O�� �]�0J�͛͆�dG$��c"O$=�Gd�!"5�	��O�lN��KA"O���b�~�Z�*�GV.��"O*��4��$&"V�rH�>ga��"O�aa"#����)r%ޅ|�`2"O����Q�E����W�Ҽ!��"O��Ϟ�	��p��.�Z�˳"O���e܍9�F�KE��rzB� �"OJI)��@p����OadDp�"O���+Z'E��+�2nL�
"O�P3s�׊pU��K�FK�5��"Ot)� eV	GjԌ����#FM$�P"O�l��ϔ�jX3�ʌr��U"O�1�1A���Q�Ӄ/���8C"O <���L�/��E�R�ٲeW�,�7"O<豄d&�\{gܽh%��d"O�ܘ�d�2�>	I5l�)L��"OHɶJH ��8�F7D�0�Ȳ"O���QQ�"1�,Q�*�8<)\��@"O�h3�CTz3YH#�ĩ�!�$ �9�d!�j\�r.țz�!�d.R����w*���p�4)�!� �P�p�^�WX,Bs���r�!�d�5r� س��[;TxsE�#+~!�$H�V4�XQ���s�}�`Η*m�!�Ӿ���AM]���C��5�!�b`R�P5��MN� ���_�!�d�	\<ç�W�*��h�!�4!򤂛l��P��͔r�浰��H�h�!��t*�y��FH
3����1R�!�$�w8�h)�M�	>Fd�C"�"2!�DP�L(d����qvD�@L�8 !��_XE!��78��Ik*�1]�!�Z9s�A!��^�0�A��<�!�D�I�x�V$�'s�d@{�h�*P!��ʳ��-�'��{؀ݙb��]k!��U���Ĺ$]U�L`1�Ǡz!�d�-N�*����ڔ$'j���e�3GZ!�d� `�0P�����1�\#J:!�\�<��8�M�#��!�!�	�J!�d�?�^L�7H��:J��S���)�Py".M08�a���Y5�T9�2�@-�y��%p��gM� �`��E��yR@Ѽ}�hB��2z+B��'���y�¬G�0�1+�"B�d���M��yB�ւn�n���иBR���W�C�y�	�?o���T��+0i����'��y�&d� m`6D\1�YK����y�.ݝ+��h��Q4z�����C��yBh���Yq�QD��p����y2ۦ����G�=�V���ߓ�yB�N(�Qٲ���#��M1����yr
�`j������W��Ŋ���y��?E��uV��>EӮ��#䜓�y���5eՊ��7AE:��C���ybe������,�#�6Q*3�̦�y�)�*QӢ<d�Q-h�L��"���y�+I�Z�Z q!��c`�g�-�y2l_�S����ރd�]�1���y�#ɖ<�&��Je,Fl�q��y
� �q�z+�]�)�0!I���W"O`q�aЋ\��\���!^��`�u"O ��+�AP|z4��q��k�"O01�+O�6���xe�֏�Ұ��"O����A�$j�NPa��=>�����"O�ukA;$�"�: �*`*6�k`"O��i��×C6>�Y0
�. �Q�"Ot�1�+H�P�p�� �cRa5���U@ۉ��:xǖ��"g����QYwϒ�!�d"P�j�pw�BRd�@I�n�5��5*��FN�I�4�Q>˓u������7�X��D�5)����ȓ6������V�AtbӯD���`#��&��'K%�O�UjCE�y���rE� ���1U�'�@m���ÂV�����7DT�t'��K���@�[�J����9ӆU9"�$iˈ�x�Б>�T�<iBBP�8�L%�c-8�GԤ�)�Ю[N�	SV�R{P}��(�^�2��
;%��I�R`(!�RjT� ��'��L��|[	��iǰ�&cG9NK��b(D�$���S !E���.�7I\9��Ȃm�(5p���L��|©٬^�	�SL�� �pp��0=9�,[T��� ��?��'��.&����?%��<��CAC�<�4#�^ ���A�K�����e̓J��ٛ�l�M6���B��q�2�1���;@l�`� C�ɸ%P� `�k�_S���R$�pSP���́5����%�O���3?`� �[��̢�h��LI��0�~�<��H1	� 4��^�4��ŽQ.�[��E��)�u.\OLq� ���'�PT��a�h��Q"�'�`�� ��`h� 	�� ����w�4+*���OŎ��9�ȓY��T��I�sm`�
lV���>1�B�j9~�c�E�&�(���&��UY0�1&�k�����"Oa�����D)��"��m!�P�*�-�q����)��<��陶&�Z=0�қY�;�"r�<����6�F����f�F��a��<y��+A<YF)$\O4�81U>a��eR5�� +��m���'M�e�/�L����(u��� � 2y�ģD���y�L���跨�%�dKt	��(O��WB��"}ƭK�Ȕ��҉]�.��8¤�y�<�R��$��!�ˍm'�d�Φ��@#qO?7�a��Њ���-1ni�0�JE�!���*�6�<�xM	�$�4�B�ȓ ��%:j����T��L�ȓ�p� �O�n�8+N�dD�ل�$��9����&7�B��!n��e�ȓ!
������\#��%�>���+g�pK��qpx�d�J>}p���k����3d*�xCȚ;4���j^H{�4l�a��e��m�����"P�'���e�ư[.����d|pCC�,���ѲI�G^D���,�(��� [ x� Ĺ�٤H�dԄȓ����"Q�#�������;�ȓg�8
 UZs�"/W	1X�ȓmCּ�c��&�\��#�N�3��ȓh@\�Q��3����E\�_` �ȓ/h�i���u�4��&j���ȓ|�Q���8}%���m�Yc|E��2H�Y
eL�]�0�`��V��m��#��]�#Ԑvm	��1:Ɓ��*�H�cQI��G�t�[���%Ңp���8���K��o���s�m�"*vbԆ�!8�B����H9w�Vm�:����P!S�گ:��4%�$F��ȓx���k��_(:�H����gl���h��
M;\@�ժU�xC�)� �a�a�ԑF�j��/дSp���p"Or��AY�05��5�1fr(�"OV�Aηr��K�(`�d�w"OTE��cʈC10�@i₡�"O楙!H�<� Q���U3Wt�|Z"O�bp!�� "[%�X=Q�R�i1"O�����h
F��c'ھ/W�C�"O8�d"Su��d�֧�a5����"O�%�+[�\^��UC�7C"`)�"O|dQ��F0�Hl�DƬ5��,+�"O��ڧo�:~�H�H�dW;�c"O���􎗗RV~��!�OJ7D@:O�ɪ��s�*0��N��'��K����8�'�d��C�A�bT�H�j]SM�Ē�����Ht�qu!�S�EX�\!�f[�"�5a��Ҧ`�B�l(�x ؓ~-��%N��z�a�Sq��3r@ӧH��\��N�e�9�m��:ْ%R�"O�u@��?����u�D���I�8}�k�6��q�@=����O!Up�	��pAh�B��D 7;a����Z8*�n�%7R����ӡj�r��o��W�U���*�x�
Ƌߜ�2a;�DY2�&"?A�c�2X��t��I;�i� e����H�A��Xq�I�M!����rJ
�'N�����5��	�RUD���.��S�Oᠠ�R��b��P�T�"m����'�~iAV
^�3=�]��
>�ti�ǜ>�V�Oy2z�⠟��}�f�4ޔbSᖖ$���iqd����?92�MoJ���ㇻj;@5#�XW!�h��	�u�̼HT+�/;����ݹc�j�E�bQ,V�����0y�%�p��$=�:ԫffE�
m!�$^�6u�A���\/�����gN_2�ɹ_>>����$�Ԙh �Z7g�`J�CL*u*B�I>hF��&�����DMG=���4Xbr���-�$k��0���H_�OHh�)ג$.ҵp�\߈��'p�`5L��LM�H��LKC>�G��Tǀ]�ĤK V�$�tD�����IY��06��jұ�v�P�0� ����2����ʇr6 (��e{��25+Lx��d��a<�ip�g:�O�H��Q�H���*���Wj�Mt�I�'��T3�&&z��T{�iUϧ<����:KK���`k\�.5��ȓF����D@:HX�/�y,��i��ɫ-O�#@��)�:��"ΟC���F����P�ɦØ�P����L����ȓ����­��)B`�Q�Q�J�+٨��RD<-%�����|��-�Z�'��	��a�=:?\�� 윹+9�<���ā��CN18��!�T��-���vK�HNڑ�$R,$}�ŸK�+j����'�f)�#n�U�'g$=����w$Ts K�/��q�ҥ��;D�`:4���`�����U(��4�",fg�&.�SE�BC�A�!Bcs��@�"�O�ě��r�Vm�t��I�Lk��l7�QqW�'L ����5e��Ћ���s�RyΓL�Hk&?�0-zs�Z�*D�"h�Ȭٓ"O<Qr%@Rr����KP02�f��V��{ �W|����k0?i��
��p�cסcl*�
�m��PxLGq����$e�/@Nr�	�0|O"�:D��F�E@��F���ʇ�")�,:4,�5�B� !��e�ܽ1Q(��J�Gz�o=�:u�Ɋ�<�$$�Ŵ��'�l�ض^~�i���L~�Y�S�kg�e�'�Џ.�̴�@��!<�2ey�����2)M�t���-o�� ��̞��Ё�a	ɧ-&��I���]s�����h��B�-n��� Lv���
�M��a�˘p R��2D���5	�Y��)�'�V dgV<4D_��M�1��B�R�z��|+عG�L�*��M�b���ϻG,hh�ŧ���Դb�CC�xLv���'�9��Q
��pᖭ�I�b�ȣB�r�8S�>����h	"� F��-ڸ=K���I�\��0!�" ����A�
P�ax򍇈
�y47OP��t��+�xUY���K���룎۾{���JWw-��t�'�v#&h��g���sc~8� K�41ǆ^B��D�`�xC�+)��O� ���.��csh^�w�L�+�'��TqW�"~������ѦWX,���O�G��?|�4�O�>m�S��%v���0䞺uhX�r3`>D����6N����i�=-{R��#�>�DZ=,yV���S�? ���td�N���֢��!��B"O�p�BH�=_���� B���E31"O"��b�<rF�i����
�D�"O�| ��%N�h	��( ��0���"OP�飢	�(�0&�9� ��"O�m#g�m�Vdx��O0B� `B"O~U�E� �)����S'�"]�"O��
�Śbz�a*$K�b���iW"O�i�e��mL�8��U,}��j�"O���&!.Ȱ�@'E� ot���"O	��"�4I� �:��=<`��"O��)�ȗ9f�V8Q�B]�=�T"O��� )&(*�a��FV��t"O:�{��ϣEצd񂯉hO}ȗ"O ���P2_Ȑ|�R�s-,qC�"O��pd��&�rp�gM�'Er��"O�}˕�[�=�&���D�"O��璏8^�e�(S�IÖ"O*�����L��Q��҉Y��,9�"O`�&��0F΀+#BH%���d"O�5�k�;5�:<q2�+� %�`"O֝�g,�3����Oژ���R"O�u�T����d��Q�ɠ	Ep�;�"O�4��ɓvƪ ��h�3|q"c"O�%Q��"f�ɻ��W�|����"Ob��V�����bT�"����2"O���&��1C���rW L��k�"O|��� *1�4����)��a)D"O�H jÈ��x �тY�t��"ORA�Ҷy�Z ��Q�M�L���"Ot1�r���2�Z1�_��	JW"Ox�J$dA�V>Z���m�D�FD�"O����Z$ۤ�붎Ѿz`Ƚ�U"O5��*,#.݊$k׮W��;�"ON��*B
ɨ���ʟ	a-��)�"O���&%�9�*�w�J�(a�\Y"Oz �`G�[f@�iQeXF�hs4"O�l�B��l^�0��Y�{N�,3@"OZ��1���g�8�;�`υ����5OD5Fj�?D�`�Gl�"IPD����I*F��EX1�!�ȁp�
֔YBvB�.|E�G�	�p��:�h�/tB�I&/��e��'����D���P%H2B�	6mg�RA%��4� HR9<C�	$I�V$ö�M+qT@p9Wd��6u�C��'sAN-Ccm��i��eX%Y�H/�C�:Y ���MS�Q�/�:~�,B�	�;��l"DȣK���̉�n�"B�I�f�Bd�1�:M����LȤ.��B��MnV)걫T��( 4$Ȃl��B��2u�pH$mB*k�0e��fC�I�9��]���O�l^���gO�,�ZC�	�iX��ѳ��"��B�gèJ�TC�	���i�a�;6�a����k�^B�	�Kn�`x�JL�{�j!�v��6m�(��D�v}�-@"[�LAj��?]>�x���*�ē�xz�D5�)�ӣb&�V�^�t4���@E#o���j�H����?�)�'+�腘�k�pS��ză�	I�doZ=�|I���S4���u�_���rÌ�R7^A��H�P��0|�(�nJ�h�Ȁ�YIV H�cB���'���@��>a�M�r�#�N�x�Ju)3�aܓ�hO�O�J��R����0�lCY6&��'���ŀIl�0CS%ƣW�̙��'o}q����\�܀@_�Q���+�'��4;�L}��B��U�H�pk��� F����'� ����!~U.|��"O�ب�	hP��uʆ�AS�9�P"OX4R���HSN�b)��%>����"Ol۴f��o���b�͚C1.m�v"Oh�
r/��Q�<Ӆ�� 1�Y[3"O��)1eK7y��"Ѕ+xJ,�"O82� O�_HLRË�9�U�"O�93
�<c�hu�F˓��52p"Ob���ݎk�A�@�1�h�ra"Oz�	�l��~����Ȩy)F��"OFT;��\�9@^	�d�/<'0�*�"O�MHR�X�5���D�8�����"O����*�İ�E��)�TY�g"O�a����e`��e"��%��"O��������<�g���Vt\�CD"O,*!,[1^�āj��j�P�v"ONE��i��\LE�tB�2�h�P�"O�U��h��s�Н���� ��� �"O��3��"*Kb @�+ܔ9� �"O���_0��+֧�V6]y�"O�=	d�2[N��#��Q��2"O�Ճ���7u�e@�*ό]F���"O<|��(��?�|%r7�Ĝ;_��;�"O�L@wHZ��~9q1"��W<-pp"O�x ǭ�-R���׀S�U.<h1"O��&OK94��RD�٠>�ᙠ"O~��pbX� b���n�L3�"OF��d�ȍ��!#?!)��"O� ��ۘ�xhTl�O�B�"O�SgCG�Y�u*�[8d��"O@ B�恤s ܽ�`����"O��z�D	zO<c�`03D�� "O�}xaMɉ;/D��;I*�ɛ"Odт�I��7���Z�R��t��"O�
�n߂b�ȓO#6�|�"Ol�ag2X�<��!��/�6��"O��Cd����� ��#{R�)�"O�|��ӪRP1f�����c�"O�\Q6�Σpє��rʁ��"O�聦A�0U�=��hZ	g��;�"O�рPg&0��1�����z�02"O�уS�3^ S�#�	J��%��"O�A���*6�<aա���,���"O��F�Ks�y�e.�1�u�g"O�ٻ�_�6�T��,
�*�D���"OP���|t�E�s�J�J���1"O�̺�����t���!7��K "O���L��;���AB;��q"O�(��Ҥ2;�Xڠ _�
9 ��"O�僵��eF�UiV�U�yb`i�"O��)Si:1�T�kwd�w���"O�5��G*3���2T$�u��"Oh���ϷG ���D�-i:��"ODI��RSl�͠RdY+��i�"OFU�t%_� q	EA2��(Җ"O�@B�ꈓ2!�(�ԍ�x��B`"O,���) &�{�Lυ2�2$�b"O��#ǩW9	}p	�`�#oH�s"OVԁ�D��h��B�";�Y�"OH̳Th�"n�zP�#N��Rx��"OT��옓~�u�%��  �@9�"Ofpp¦��	W��&쀀)Y����"O��3�ǚ*h;h|B)�>9��b"O>��6��z�h�@i�8m;8h�"O� �]�H��N�1����#�D�6"O�pX��M�I�,��"��$y���"O�,X$�4@��yS�V-`h9��"O��mG��`Y8#
���U�6"O���Ei� ��� q��6DF"O�r���'�8���@&S�6��"O�1�f��J��xBdE�d�����"O�qT��-d;���cK~�H��yr���-���oJ�m���UG�yr�	�4W^�J��\� ��UC��K�yBF�7^X��SMP�gxbb�D�y�kM�XA�h��_�(gj 1�AX��y�&��Q�e=o�\��]��y�b�&Y�&iU��7Zq�H"G�	�y�"Ռ#DV�+�M�O�*eC��߫�y2��S��ӄ��M�x<���y��4��Y@�͎GU��D
�yZ�={%��,U"dS	��̈́��،���G>~i�iqw� #��ȓ?�t8�ʊ��I��
�n��ȓGC�9����)K��H� Ո�Z��ȓʆ�
�*�MU��������"a�ȓR���P)�,cl��!^0�����T� �����h�h��t�ȓ���a�ȋ{���a��..D�p���V�xܡ�IЬK��:s&+D����� �do�M{��M�BP��@�*D��ɰ��V�؀`�+����<�;D�x��];\�.��p�+ ��uct*.D�P��$oa��G-.���BW���B�ɊpY�,��
�b�"�CfG����B�I�-�\(���">-�Iɣ����B�:Z����6�@>���0�����B�I�b����/T�^��{�-I:^��B�I�N
�)�',�V���31��5�B�ɳ_6��oʮ`�%A ΏGlB�	lᶱ�4,����aK��d�B䉔Z%)�#�b�U�$A�9#�B�	{rE�L�}r|	�SO�!"$TC�ɢc�Шgʙ94�r
R�E�	?hC�	�&I�1j�*r��d�։i$�0��"Oؠ�"b�)BO�L�կ��9�ɑ"O��JD�tb�jA���<�r�R�"O�aR�O��8���*s����	Xd"Oh�	�N�h�*���9��4�#"Oh�""8���s���(C��h�"O�����Q�,y�@��Mx7"O�Y��X302Lx)�,��}^�U"OV�2��p�-q�a�Y���6"On!���W�[v\Zq"ݱ`l�d"O�3� �45��}��U�XR��"O<�1����p��9�f��7"Oz�R6@�t�(h�v��$V�����"O$��0O#���i�G�2ֲP @"ODt�h�"�p�B�`����Q"O�5��$�Wt�@�$��>P3�ሔ"O?H�J9��nU( ԥ�"�0b!�<H��B*30j�%���#w[!��3wABu�F7 ^
: &/P:!���lx���q�0RY�L�����J�!��Q�ap��@���9G:���S�J)�!�D]	2��˟�T)>M�EGy�!��+|��e*��H"���õd!�	&�8�Ȣ��#n(��1@ªX|!�� ���� ,@�4�2� ���0��"Odl8�o� ��=xU�	�*�`��"O�͠ ��q2��e��tS�"Oġ��+�mC���8�,��r"OZl:BŶa���FN�Nr1c"OV)�3`I,� ����B�3"OR�Ǆ�$a�}����)�v,�"O�Ya�Š�\�5Q�m�f1J�"Ol��JЯ;B�B	��J�d"O"��ǎ3
�1)!��P���W"OD��RU����&}�b�"Or�QA�S<��ً��R�i����W"Oθؗ닥yv� Q��T��Z�"O��훷9�b �(́�@���"O��x��G<�y�CҸs�H�"Od��6	G�?��	s��7�N�80"O\E�P�U�ܰu��*�̰�"Oa*��s����-��:�ND�G"O6d�"��)i�hLj�5,*Q"O�tb��/�&���".+���*�"O���Cީ[��TX���5U2
D"O����e�^��9���?!Nh��"O��XƉ��/�R%"N�aCR�:w"OXE[�hC$'�j���o%��a"O����M�;O������1v4�%"O\�@�f��F`ȕSt�9K�H�v"O Q��b��Q1υ,re+&�y"�I�V����ٿd�ƹY�*M��y�BsԬA�LV a[J��eV��yr� U�|�'��
Uvr��-���y2�%j �����BL)j�8Q&N��y�� A�ݛ3	�xמ���I��y⫘2}��	ׯ�;�Ҝ��N%�yb�A&mn �8��K8��}��DJ6�yB,�M�� �%� *?�|X�oE��y2��&0M�)g�C81��<�g��yr'�:���6K�<;RfF�y���4�01���ȴ����Z+�y���ovvmI�hE/ ,��!�
�y")Q?j�v@�a�L
�;sAɃ�y2MË0�1b�
�C@�h����y�M� 6��e8bo1+�*hL��y��(%��Y�V��3G�9"Aũ�yB��1�G�1q��ɔ�O�y����5x`ba�]�Q=���C�y" y�Lh�¡�Y�8l5���y�jQ�j\��F)�@������yB-�)x��5X��2J��h�`���y����b��G�=;]�5����=�y�f�Y%�mȷ�BL�C2��y2����AqE �zx��!�'�y�`V�w������0p��ڲ�!�y��8-�hh@�
62�����&�y��ȋ :��W�M3��
l��y�@���u9��H�-��|����PybM�� �*5"��F�S%�K�<�'�o�!x.Ec$2�k��m�<�7�¼mNj����	pF��ףG@�<)r���5����U� #���-V�<Y�Ǝ��n�C�cW� B�EK�O�<A��O�1�p�KVҞ	9�N�<)$��$� ���#�� Fa�e�<Q4�T�׌�x�)�vct�p�a�<�`-2�����^eD���_d�<� ��J�B>F# �K��]�1�l��!"O�e�֢Q �����Na����*O���dF6R	JQ"��T�R}�
�'R��K��λ)�j�H6E��N�T�'a�$�   ��{m�NHW�<!����SH�eIvcE'y�D�#�$SF�<sB�|��5���	�[��_�<q�A��]B5a�U���H���W�<��$�{���C � ����a)JM�<�q���ugR��DK/�lh�!�R�<�U��	J�V|�@��:>�Z�H�n�P�<�7�Ć_�j�90`�����N�<��C;J6�*��gV�����J�<��K����~|�D�e��jE��_����jѥi��i���r
 ��ȓZ��0!T�˔"t��h���?� ��!cvD��K:��ݠ�A�)B�ȓ
.l!7j�(a:��Tc��<�J��Z̰q�d�F�\���߀_�0��F��� �G�^d󤍘��y��^Vp��ē?[�e3���?4�r�ȓqiD(��1>�h��4 D4eXXɄ�+I<��!��/�:%ئQ`*L�b$Rmd���J�jɄ�	-0���W�g� �[e�	�{_lB�	r�@�j��ԕ+}�i�Ǝ�n>�C�	�/3.ب���?
Sz�1vFz��C��*N%��0a�"P�}PD�>f��C�ɬ@:X���+f�P���/x�C�	����z�ɛ�<�+d)�5w�`C�2� �7&�i�����5!tB�	� rc�N/0����ǘV�>�I���V�<d��aݝ��+,�
.� H"A�' f���� W%X�H�BI ��҃\Z�hI~��� ��hA�J<�(b���(�J�2e�YI?	G)P�u��AiE�֩�0|:�!�0 9I���I\"�:��ܦa�F@�'�R��#�Z6�)�'������k����F��<b���勄)���� �:l֝�3�����0�Ov:e��I޽"��0Z3��$I��q��n���#b�N�ѓɗ<�O�q�FD���ۿ`lDL؆��T���sB?���'cRmxf��I>�	ӋF��lR.����N_~���q7�[\>���&=�-�alƜ:�d��b��4��N�c2��y6�|ʟ�=�Н����>�(�+�%�����x :l���өnQ<Q E�K(g	CK��<>d���S����u��4�d�S/��U[*�A@(A�TͰ�h�"O��҂��]U��(a���]!���"O$�K4��W=n�n��(M��"O2�Jbn�!~bMn�T�5	�#D� C���5���\�-�x�rO!D�$Îͭo���� �Ja$u�>D��Ap�×t��c�ժb�VU0#'D��0�˟��b]���T�9�KU�9D���ӈ��:�|�"-��py�Q3��6D��;qG�2	�&�{1�OzY�1��?D�h鷀�&lɊ%��hٲ��i��B>D�(�vg��s��Y���Y�={�%Q6�<D����KߞCv8�Tʘ9PҌi2��&D�<����"h�A�ŬE�(I;t�/D�P���
	nrm�qG��aJ���"1D��C�
�*K*50��O_H�	fn-D� qV�̙F�4IS��zW�$��c8D�$K�g�y�<tC��?�U`S 5D�Xb��U/=�2<�k-l�@v�1D���B"�^�*MK�-�p��M1D��3���J߆�:�Ĉ %����J;D��;��#G�(�8�C,39�
��7D� ���޲ys<�"�莔 t4D��8#�ߠU��9����f^f[�=D�<(���a��!�!��P�V���7D����>(Қ|�Ԥ[$luT�Ť2D����!W�B���A�W>{$�#�+D� 4DĉG}ޕkǎ�,L���AG"/D��K ��4{�(P��E�ot 08gE,D�̣��m5�v�B�k���xg�(D�d�d�@*/M�<q���$FB�+b�&D��h��	]"5����0LS�!��($D��i��M2L�>}a���|���t�!D��+�J�n]K�M�bM�VE-D�(+��	[��k�ǝTD�5�tN-D�L��E9�;`�*K�)х D�H"��U�$����#��A�yI?D����@�OK�ЙgEٛ8���`WH<D�\:��:LDK����R�����@?D����$B�Y�jK� �Az��RD<D�t�EW��8pd��ހ�ra@:D��*���sX���ЂP~��	e7D�h#oS�V�D�f�	�S�dC䉴"��1Y�R$	`M@�A�x)�C�!/�@xy!gDtX*��Q�yR�C�I��@h��#<n,�۵�C�30�C�^U��x�ʏ�(��ӧ�?f�~C�I��^�3�\�#���h^F�|C�	v�j(P7�� X.ڬ�A�o>C�I�Bf"�q�I a�L
f��"� C�ɂ6����F#2�����T��C��2c#����jU&��WB԰|��B�?s��)�ˉ����ʀC�I)
�H1��=+� �%΄[�@B�ɝPl��:���.P�zt����z�8B�)� ��s�d�?h�LH���/CZ���`"O��[&]mʠX6́=3R�4��"OB��+ �y��q�P%WM^81q"O4�J�JR�s����1+�$yG,��"O`���ҷt�0����4���@"O|�$M3�T1�*N H��`+�"O�)à�	:E������ɫ[���b#"ONA�"˘n8�uZA�T��EP1"O\a�
N��Y��LZ V�޸�k�<�ĕ��P	��Z�b�I�OQ�<ihR4b��8t�0_q0P1s �E�<��#�u�"<#C�σ�L�A�B�<q��
[�V�j�V�W縰I�G�<q�h O�}�'e��f�f2%��l�<�$����1n��W�I3d�^�<����Qo^����8�%k�B�<i��ܩih����ĒurQ!�&H�<9f�G*-�Z�5�Z2�DAw@i�<) ��-��8��n�&�H�-@y�<��D�[(�!�χ^`֨h�/^r�<��G�
��5*�6l@���g�<�R+d�0�"Z�P�pᥣLK�<�MG&����Q�Ll�<	��	��	�W,I�W�>uʠ�B�<A�z�6��СP�@�N��łt�<��֦E�n���lH2Jvd��L�o�<��+�?v������E�Z�1��g�j�<	�F��Bm�])rͮrht��#�d�<Y'�9R�l}!���~�TM��_�<� z��`kQ$8��Y�]	!�].uw0��'���T��)'��g7!�Z�e�����+:����\3#�!�$^'f$X	�GE%P�ǎ��!���E�ҙ����G4౧�R&t!���w8
�'��Nd�H�W��hK!�gĴ���3AcRY�fFN@!�D�<X�`����a�naad��Z!�d��,k�|KV,(5��
P���9A!�DX�!y�m�D��*�!�b�*!� <|�J��>�Љ�+ۖF�!����tmc�c]<O��4YPK� 	�!��i��	�KB?�j�Q�	��#"!�DA�.��`��~�R��5�Mr!�Q)O���A�E�/��U����A�!�d4cMp�!o�3���-�<�!��C܀hK���<�|��"�\!�T�7/��7!	�v��1d�J� \!����8�JՒc�4U)�$}7!��Ɓc����°-d����*I�F3!�$�=7i����f�;[���	���*'!����~��3CE�u�hء&	��j�!�d�� O�ڶ��g���ѨN �!�D�B���t�_��|��]�!��:z�TA@6%.I5v@p��"#�!�$�)4�c���}v,=��F�^�!���8K�쫲խwuԽ"���&	�!��	���+ 	�gk�tR4!A�]�!�H�^)��ÒA�4?L����Ə�!�� P�Q�Ԡ�($>���`��Et!�$W)q� �����|tO@�SR!��RBX�q"��>rh�y ��N�k!��u��Q�'!B�?��	�B�ԧ1!��>:�"18B��P�JA���_�7f!�$W���)灇�J�9YQ��;!k!�� �4��'V Ēl�E�I�Ҏ�s�"O ��g�E���p(@]>1�hL#�"OT���k�5=���e�M/4<��5"O�*�6�z!��N�K(�XP"O�e[�ǂ�X�lɲ@$+vQ��"O�ȩ7�%�ҍ��E*>���"ON��_?�<���.��U�"O����B:l� 9��`S�n�zD�@"OFA��H�*���3��_�>��6"O����g�X��'�7q�8�@"OJ�� ^�I�$���_2P�����"O~�#	��^�P�F�r���C�"O,|G�ǂ{LYh���8b$H�"O��j��%�txq�տ%���"O��3�B�2f��(cD�[!&��v"O�K��h|
y DSy�-�"O������2j߸�����&n� 0��"Of �g�͙;�c���.Pz�鑇"O�I�%�3� ����`ي�3�"OtQC���	�|I�������ؑ�"O�E���
 }�`y����z�¨�W"OVpbqo�2\ʨYg� n���s"O6y!�!�.#A��c�#](8�����"O�}O<��h���C�kuZ��"O|bq�U?��}�����\N4�F"O�}�Ң�\�l)D�
����"O0�+҄V�QJ1�2d�(VQ`��"On՛�"aڲd�����(��"O�!�tl��]'qk��C�=�> ��"O09e@��k���{�B��\�h���"O8$ʐC�V��他��48�>5��"O�=P��o�.Q���5+��+A"O��w&�%͒ {��K�'4��"OV[�[�0Sd�pV�l̉�"O,���!TN����V4��r"O��ч'��[������R�ij��C"OjAi�*Gs���'Hï^�4�S�"O>a�� ��!a�W�3��4CE�T��y�HX'2�DY�Bђ)��u�s�'�y�,�b��}PV#K^
�Hd��y��܏l�1�P�L�>==��$X6�y�h��J��u��E]d�Ձ��y�	��Ai�u���>>7�i�����y�Īe�DR���/?e�qQ�bK5�yB��TG�� R
O;z��2dJ��yrF�5�M�ɑ�U6��c�y�΃�-$�xc�KB�x�h}��)��yBd F���w�G1#��j�JW��yb慖J׸��v@"#��}�ń�y"��_�<h�$�ϨC<p�˄�ǖ�y�9k�0��i�V�Ʉ�]�y��,��]	�
�Z� A����yrfԐw�܍@�C�VKHU��':�yb�g�6��0�șK�KB���y�
�O(a�!-٤���M��yr@�_4��s���t�)�r��y�\��,��rd�1jG���솨�yN�9wh�ʅ	�f/nh[����y�� �-xc���6�fL�a��y"g@�x~��@�@��| v�"�F�yb�̉�x����h�"��3퍻�yR����>`ˤ���Iط�y���(b��]�#�V<G^ISA���y�"!��,I��I�t�2��C\��y
� �:`,W=:�rHC�,A+*�ȍb"Oح�q)٬yU2��pMV�����"O ]�G�ŤkΒQʗ�'�q��"On���à_W0\����k��8he"O� r�@36��7����D���"OJ�SE�O.����A�W"Z�f�"O��EPQ��-!!!ގ,͎���"O>��"Ǚ�q(Xp��@' ����"OJd��e�<(���O
1A�c�"O��s/�7b���3�`P�U3��#�"Oֈ��R#T��P`�7L̰��"O��@"#��x�@$�&6�@��"O�e��M{<�Ҕ�-x�4"Op�J�
��팑 �A�=Sb�aYr"O�L��B�K�R�I7A��a�(Yc"O��d#ݍv�@��`
A@^6���"O��JL	xix��0^���"O@d�˞�-F((���UZ°�5"O�<��c�H�xEH���0D�pK�"O�Y��D�H&L� (ǰu@>h��"O�\��   �<� E5_�xH3�ǀ>�yB/B='�BtŇ�I�8���+�����ʎd�fA�a'��O �c���4:x���@) �F� S"{��E���Ț�~"⇙��GxR�\�~��u�mL+ R�i��R�	NVi�W�w�̼F}2��ti&��ĕ'{4ҍ̪�x�!��F�'�V�0Ê�z��a�-c[�O��:�슎2E�����D�'h�d�(�2w�N����90��+�8;vY���B��"E��c@��ħx@)�V@,@'�Q�_�ES���l��RԂNv��ӧ����`���2r��K$�����F(^
"�$#�Mѻ I�	;�k�j��OC�!{��LR}r`H�Z�Z�i1��\�E*�+���DƱ4/���4�װ��O� 2)�u�Y�k�H�L ���>9 G!�#���4�DS�"��� ���'pr0.B94�\�ȁ��y�gn�%@��)R��o|���!�v��A*�M�7�H�q`�jxf�zƄ �G�r��E�T������	�7���8���C�JJT��i	"2�<����T�LY��''�ܴ�`��Ua&y�p��(D:Bȍ�(�OJ�*�/̓S�LTjB 1�4=�	�'p��p�D؛z*g��$7	.q����4I����gR"t�Ls����'q�l"3��>	A*GѼL����^�:�x��R��$�O��
�L��׈�|�ܱ�u�X&��� Dy�<�G�]Z�yjA, 	������R�{ �d�Q	�m��ɚ�H#O8�#����HU�|���%E���1iD�l�>I���G${0(L���ԼtLP�f�3�O�PF��7qW�,;��� �␘r�>QV"ӕ@>��	Q��)��|��J�d%4c>�W#˓b�pmX��3G�l���9D� ���\�-8F%0N�,R~�b4J�h��=��T��	h��~2$V�nø	�̡f����Ɉ��y��O,[:��LI_:��uـ�?��#ќ(ǌ���c,lO2����Q�y�\h����W��@�%�'Є(U�
�\�8�n�<��I�ƙr.�W�P�{�TB�ɤo���h(0��@g���0⟘�CBǀO��-���ӾCr*)�w�[1+���p1�"O��Bc���9��qC�1I�*L�F-0\����]��"�g?���".2P3�c�/*s��r�Vo�<�Q�K�\�M;P��%^*r�F�`�	�Y�Q B�$_+a{�?w�j�
"d�z �0P���0>	��r8n  ��\��YA��8d��3͝-rc(��ȓI��u*��ީ_����J�}�B�Ey"iԟH��qF��GQJ�@)G������!��y��5
q�4�e��H�ƛ��yb+ߣs���:$�PX�r�a��y2��R�r��GC���¢���'AZlq�N}����+�f��<B�K��B��Ih6�9�����.*#*R�)�	2żI���[7�h��r�`��� ��T��H�*a�LM�I�6���	1S�.ђ�-V14��O): �F+�*R�J]8�E �W 9��')�઀�8/���5i��K ~�/O��ҶbU�d�"��M��|�A%8AnTt�	٩��`��u��\�ae�8H�"�����%0��35���&���>�7��7ET !�1�\Lx�JΎ���+��b��F~�_�Rw|T�土��Ė=E�ތ: ��YR-Y��Idid*�)Qa"���Qs�(z�.�V�I�X�j���5���� f�:ʓPv� ��1 S���pYC�4ttf\zOU�$Z(��"O�(�-?h��ٗ	7D���0�Q�`�V�^=%���GC�F�iȿ@�	"�Ϧ>1��έ3��<xv�5,�@ +GM~��i㏉�=��4��iJ�+0���Ԯ�s�����Ȓ*����v�����_uF�"?q���%-UH�B0d�p@H��g��X�'�"D��eU)Dܕ)'���<Ha�Z�H����_g��CS�S�*�����@���C�
P\B�[c66�*)�.���:����9��ן�p%�K/"±1p�i�5��ĳ�g?l^jH�E���:�.,;�O�̓��ԃ�_ {�h  cZ�'��Qh�"�O����0��bO��"�t�<�l;�#ۊ"��`���IZ!wL�YH��b)��D�g	k��-�6a�ڟ6���S^�,��坾{d᱃��*� ���xQ��S���9�����C�fQ6���d��nH�`r�ǃr���pu ��	D�����T�^�)�����d��n#V�%E�t����#@~��;C��Jm�X�t�&�~%*��'}�h)�I�88��f
�E������QDP62X�E���!<Y�$�d�rNe[c�^�$ϔ�;&��0rV�Z~����ՆH�0؅�	�$�� �wKp\��2�τ;d/�"�B�y�H��刯D�R�;��d �IٷԚr^�SF����'u,�aS*}���F�$:D��J�'n@92#/ν����'�ޤ��"�/�j-Z@��'����G�*��bP�V"����ѻiq������{��(��ŊH�z�Ӈ�L�w���/.1��(0����M��9|���JW�]~�9cc� #)Y�}8���;��t��K13~ �
� ��M4M��x�0�!x�i�f����"|�Y�枀q�(�֪��s��9�G
i��%S���*!e���^��pL�S�B�I%R��\@�¤i�~���KT�'nX��I��6�(L��O�}�NR��ey"��fd��su/��X�����\���U�PbP�y���1q}�x
�͓:8-rał���'(pxJĂ
*�ax��5f��8�ӁN�ﲵ����>�y�!��[����@{��Ԋ��yr��X�|��w�.MgN9`�O��y��8 �Tʔ�E� ]($��y"l�=]U0����9=�bipW���y�F-0��|1�h��7�R5��P��yRi�M�����"�����Ί�?y�dЌl����|;��7�ϸfnޑ2�C�%�a{ͺpF�h���O��e
8%90���N6p[���p"O�\��_871��!PNІ@�1���DÌ"�]��E����jM�)B�K� ɐB�J5)���"O8�j'b�6X���yV @���cсҭs(p��>q�b#�gy��ް4@�� �G�dkr�Iqꝣ�y2�D�Mzt5B�@�%�� ��kK�{J0��V r�hA
�iktȪ�x/��P�#Ϲx����Io4�а�n߼t��$�(�>��U�_�"!^�Q�K_1�!򄓲=$ұ�2�\�o�Rm�����qO��x�LT�r���1��i�"(����5tPYw��'s�!�dX�%!ԩ��k�$h�`�DL׭[��-
�B�(��Z�D�|�'Y$A���ҏ޾p����#f��m)�'�ʤA��'Z��0+$'�SL�|1ň�
�a��i�3�0>y��܀�PKV�s)nx���A؞�z3���Mpx�tG|�ѥX�/�h���!7mr��ȓqP�]���b�1 Da�,M�?��âh�"B6��	N4p!�@�LOD]0%�Fz�<q�&�LV�ԑ�P�1G�\���u�<a2�D;^k���)ݺ>l�)�g�Wv�<�U���B����DZ�l���(�s�<�ǩkIz �q�Z!�ӕ�Na�<!�Ő�~�hb3d��"���2@	j�<QP!��`�49j���9B�lDZ���L�<� h �"@�!�����٫Z�hʅ"O4i �I@�]���8����"O:���	 ?~1���2D��w?ʉ`W"O$� W�7�<���7^�Je�u"O4���jЀ[Jlp�sɳ+b #�"Ob�r��	�=���K�/����t"O�%��RHu0�@�%%Ȁ�J"O���($'�1Y����^���"O��(x�p����E;!h�\��OSb�<�F�
�7�@�1n����G�<ٖ�$
���ퟙl׆(6��f�<q��T=/�bL�b�	�F�ܻ�CS^�<)G�R2�!D�)
%£a�`�<��R<#C���Ac^�v��1j�X�<�PO�!e�*S���d���b�R�<�4��-��UPtd�R`�i���N�<��kL/:L\�`�?�0��RXF�<��ǋ�{�"��%K�!w�T�1��v�<����"�^����B"�m�u�ȓ��:�� ��i��"�$ǖ��E�dt��E1�n��S+P>f%��R��-��Ȍ)A��hjP%�sFf`��$��@�đ�\��	r"�ڦFa�0��t�ܼ�S%�8�c�!���ȓ�v|B�. <�r��23�z�E|��5����Z���Xd2���H��M���>D����.�9T�B��.3��!��Njϸ��CĔ{-�B�?ئU��ӷZ��u1�m�#�DC�3kT���I�PL�qC����b%(C�	3T$�%���)���N���B�	�W>�<!Hm;�%ʝA��B��^�h� E�R�J���F�_�B�	��Jx�B���PH�N�B�əx���sM]������,+�R˓m1B�<E��-��(1̕��\�"�"Y�ڱ�?��<�S�OQ���m\�z H���M.�bܨ`��O����8,�B"|�A����s�NTNU�|�qe���%�x�aE_s>��0`ݑ��y�'��><BS�2����<8JC�2��La��?�) �øo�$ ""O8�æ;�Q7��L�:�:�"O8v�׏xꄋG��rN� A"O"��l\�zu �H׀�1�fB�IP8�L���<�Rn� x��)��#D�TGQ�X��)��+ܳ	�����N=D���-�[��@cj�3i�J����/D��KdD�0o�1�W����(�҄�.D��Hhҁ^�8�G��6<s�Ɔ9D�̙���ɪD���5It.LBBi7D�l��-] 5`to�(*�A��0D�<떫�7������}��Iza.D��SC�:�ԥ�0@F�Z+�)���(D�,��"�S~�]���+n0X�%D���wm�'`kp%8�KC��4���!D����.��b�����B�	�����*D�@:E��^캀�u%�=iL���E'D��́k�4y�\���+d�#D��;�C"H��	1�� ��q�M=D����k�Z�~Ţ"c�3D��	I��>D��A��C �U��#�7{��
@7D����mʕ)�N�b�MC8��I#�`:D��0aG� {I��+q�_1E�E�6D�������g�"I"�J�+:e3�o3D���D�Q4� ���ئ�*A�`2D��U�^�"�\���<h�)('c*D�� �H8Ə��Ib���Wg0`��%�"O�\9D�9B��8�f̅U��T*"O��c�ė�>��6�w���Ҳ"O�����7��9K�㏇c�H�S"O"ux Ă!o|h`��"ĵ$��1#"O�E�r�� g
$#T�%�DI!�"O,���0�@�
 ��M;�"O��X'ʈ)VѦ�yb�Bى�"O����KN�fj,\�qd	��:�Z"O�1��@�=+j��@d]�8k2"O�DÁn� g<��9�CU0MB
!Iw"O���b\�*l> x��L+g9rᰰ"O@�;�-��/`6,�QkC�9�@��"O�m��kZ
G�00�0��-J00�"O��Zv�͉1������]f"O"A`���4Ǹ�Ү�9�l��u"Oԇ1</��O.X��"O��2ȕh�`K��X�ڰ��"O~ �@I�Y�4	RQǹ*0FthQ"O<�������Q� 1����"O�u�We��*���H�G�5^����"O>-Z�k�<�� ��W�R�4�w"O���5��P�Hj0��'x�`�f"OLh��T Ev0�#G:1W��y�"ODћ®�C�xMx�r̹�"O�}�,�,����\X�Q1"O�-��̭i5�-*[e�B��%�P_�<���$2jb�W	
��āR�.D�8C6���Q�4�A1��1XE�(ȃ�9D�8��M[�T�$�VC�Z[��p�b8D��w(�`8�e�S�8>�AH��4D��R��Ș�ȁ�`*"
�U��G-D����nB�S|<�0�
U�3��r +*D�pP1�	`��5)6����m)P�-D���⋗G0ĺ��`�F!D����"�� �2Q!�M�|�l�C�#D�{�5�H��&��QZ&K/D�t���׍_�2�Ac���V|���+D�p�VMֹ:y�A��	PC�%q5'6D�,K �T�Z�Tq����0	�f�5D��+#G�'��)SJ�.&���4D�D(��D�>��|arI 9I1�H.D���֩w��+V�ܰ�$d`�'2D�4Y��G�[�ڼ�P��c��
&#0D�����7�&%! �m��iۖb,D�D+ ��b���@*րBB�;�i,D�!� �=~�������g�(D��P �� $�A�K��,־��B�;D�Гd䙦St�(��&L��&D� "�ʓ�!@�����%o�"�B�"D�H��� M��q��^/TG�S��?D�t�ǭ�@Ȳ����+:��}%>D��s0!�I->d�ق)���I��&D��y׍����S�� =*�� w�$D�� G�#��1�ф���K>D���u!�B���iROLp%��M<D�x�!�ϩR�橒�)�dx|��n>D��.��yRZ�@��$K� Y�f'D���T̛�Ū����>�:�0D����A���l# I��T�C�� D�
��־,K�T�	�91QB�<D�,��B��I�g�.!?��!"i8D��悀]c�ݫ��?��lI��7D�\xU(ĭO�D�+��<��w�7D�� z�ďx�!9�ǂ�x�PdA"O�P���6�R Jcg��0��a�"O�U1��ٓ��X��fY��"O^��� wN��,� @m��#t"Op�e ��5l
��+�^���"Or���H0Z[��R��Z2(��3t"O�Ms���0�jݹe� �n؜�#�"O.�����9<ExvF؎o��TH�"O�8ĩ�u��[�DM�i��� #"O�ɛ�-ˊ!�r�۪)��`1"O�bt�A�1Kڹ���ʓ%�����"O]҂�+U`�l����)��3%"Oȡ@��7b�$`s"�P[D��i6"OTI1R���T��B�|���"O���c��>��9���5�`��"On�f�[����I�
�hX@��"O�� H�-� ��6)��dB:��6"OF��`��2Hv�a#��=B��iZ"O�`#6�ߚQ�����oº:����"O�er���05��x��+9�ޝYA"OhW.�IF���-�4v%���e"O��+VJ]�_/"M���$Q�"O�XHQi��*KXQ��H
R���t"O����w��E��[)��=�"O6a�F���ZU��'C1� ���"Ov"�"�!}�e�  �$�tl�"O�x,�t+��ǂZIfT[8�!�ҏ7��#Ԭ�>A�!��ͯ<�!�܇p����iS".� ��ׅ�!�:5!b ���]�4��c�%��'$Բ��ʲX����I	�Xvl��
�'��9�+P����:M����'ҕ��C2���K"2�T���'����A�936�	���*�6,��'�|ʃ)N2��J�ɖ"rfy�'堘Y���G���g������'c��ǭŀd8aq抉��
�Z�'���;2a�a
y�5/��T�.9�
�'
p�a�L!6��{��F#��
�'�h�s�ыc1x��� ,�B��	�'(rdRE���������S�I
�'|�}8҈�-+�ڤ�'S�!��@�	�'`�
#���a��<��Dq,Q�	�'�bm����Pm���p��'),J���'P�q�fhI=�� � ]�|��'�]�'�	�V���١d���i*�'��H����)'@�i�.m��I�'%¨cP#�(6�>[(��w����'k���M6+,����ѷh�uB�'�12��ϛ2������ڤ�	�'V�q�.�af-�D����~���'-��4LZ�s-:� ǌ)�0���'{6�rqF� 0�!�D��9)� �@
�'M��R��,V��m��a�<�t�C	�'\���-O Zۄ�H4LG#
��@��'�4ʰ��^�i�3.�}H���'04X�5.�	R�nx�g�V)*׎	��'ʀ�J$
D�
n��(�`M�%�-�	�'�PR'�â[L�����ž!~�s�'�%��!�+">euMA�&"}h�'�H�ʵ�/)vؙCSw~pz�'�F4��݄,{���e�DL��'�ViqT5�6H���U�6����'�dB�-���5
!'섥���� p����+U���D^k����F"O�0G�`+dU��DZ;Z�D�b�"O<�Xd�8Mf�,�֣�v��p��"O���kL`J�|9��Qu��B"O��QЄơu���Y��`� ���"ON�����N���b&�X�~<X�"OT���I��
�����j��!!�"OE����\X�$YT��;c�6R�"O�]"��C�<uk�3:�d���"Op(;�����"1 �*F_��U��"OL���C�?#>F��bÝ�0ĭJe"O���O�(q��1��"%����"O�GN��ˬ��� 0n�v�0�"O8�*
ɍ>$���pB�^����"OJ��bA�*Ǌ�Y�.�!gѦ�8�"OL��3���D��	�Ѭ��z����"O~0G-�
Z_z�k7�'c��L��"O½p�f
�|n�&Ǌ(6����"O���� ,~�1B�%�%Kl~�"ONISc�ǌ'�\I2�T�,el�Q3"O�d���I���q�6Ώ�e����q"O�(;&�+F�L��+�r���c"O�����B%_��(�Ӓ9Z�ȣ"OTLK姕�X@l<1p�]�$Q��hB"O=ZR)�H-љ& 6ך0�B"O�E{��B<�y�% ��q9�"O��+�̗�T���oP�a1�"O��"�/#�2$�#j�<,cH�j0"O��Y�Ē�s���e	S�6���CD"O:,��-�f;8����=:*	�"OԴh�L(aӲ���fK+Y�p "O��Ҕ�7\Ř!SP�ұA:4�zu"Of�qTeY3\ވȀ5��0yΰ@+�"O��c�)WC��iJ�$Ū[����"OԄ��*�"�����#џ'�"X*�"Of��fe� �=Ec��#��p`�"O$Q@C��)=���\�)�V��t"O^��� L}�6��T�O�?���
�"O���M� Cl�c�"߭�<5�4"O��j ҫA��,���سkX�Xن"O�|yq(��"��}ȵ��?c��}��"OZT��ʘ{F�$��^��`�"O�̣э(��m�t�D�T�j\��"O�,�F�$��h2E�!V���"O�����?�P����']�`�ʗ"O�����F�a���B��@b�i
�"O }���?�Q)�I�C��!�"Of�@�"��~�6���I�F���0�"O�p�S/)8�6)9ba_�hNyJT"O�p;5j�+[� !)S`H���"Of��6&��D�qi<bE^� �"O�T�F�� +����H��Lx�"O�sB1S���0&V�%�B=I�"OF�2r	�2�V@a��Ϲ{��ದ"OB��A 
  ��   �  C  �  �  �*  _6  %B  �M  iY  'e  �p  @|  %�   �  ؗ  ۞  �  _�  ��  �  _�  ��  ��  ��  �  K�  ��  R�  ��  D�  � �  � Y �! ( 2 �8 +? <G �M \T �Z �` �c  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+q��62\���<4�d5h��'�B�'���'	�'/�'�B�'��x�.Z ?܎Yf��0d�tx��'��'���'�"�'��'���'�nY�5��B��0��g��ծ�pW�'l��'C�'���'���'���'b��i���8��}��dK�� �C�'1��'W��'�B�'���'���'?�%�����غs�9
lk��'A��'l��'B�'��' "�'O���ek�92�lu���D�+��'�"�'\�'���'��'B�'�n$Q&菷U�~�
�"��]x#�'���'��'u��'�r�'���'� �H�N$!��y;�Ã+K�f�0�'���'$��'dR�'���'���'�Fx-Q@�蒠�6/X��o
�?���?i��?Y���?Y��?���?�Po�^}��� �	\V�p�'F��?��?���?Q���?���?!���?auj+2��!� :D�|Hʗ��!�?	���?���?y��?���?���?y��ь�����/�&8CTtꖢH��?����?Y��?����6��O����O��DB(Hc���$��[��$�E/U��b���O����OX���Ov���O�!lZڟ��	�P��H���L�!�"��~�-O���<�|�iӸT���_�6HF�Z��
/��A( �C-)l�	9�M����y��'�����"қy����g2-m��Z��'9�훑u*�f���̧ca���~�6DI�o�P�YfJ�z�����ND��?�*O��}2'�X.xȝ�����\����X�jƛ��!��'���nz�]8�"D�O���3CmX1'�̻%��՟����<a�O1�i��u����9o���3B��\;�슰�"����<���':$F{�O����>��&_*�xk��Y��y�S�t$�0�4�4T�<��f�5KQ.z��N����	��A���'8��?y��y�Y�ЫIX�cHp�s`䆵]�>L�p�6?1�T�q0�j�'T�����?�ѐpI�Q�Z�$s.qR�����D�<y�S��yB@�#�B�a4�Iy�Ą �y��l�ƽP3���b�4����T!�#^��rd���k�f!z�$�yB�'�2�'߸r��i����|��O�x!*�m�E]Z����gA�4HTb�IBy�O1��'��'��ݥk�, D���-��H�銙r�ɽ�M��"�?����?N~��JGX��7h�|l��q�V!{CҠ T��2ش?1��(��i� ��B��;.��q��ѭng^��$,��[>�w���~����:3��ɓl���S$��	-Ix��P)L�9=(T�I韬�IܟD�i>��'B�6-�<>���F�H���#��,ƚ@(V"�%����ɦm�?y!R�4�ش�&�}� � J"l2`sg 3ܼ;�n8f��6.?Y󎟺�*��#���}��]	%�� ����6�� 	0F��I�������h�	ڟl�IH��eq�i�@ۺ,o�	��*B�S�A��?���q�6-1��I��MCO>�T�������4�)�x(I��-N��'L�7-�Ӧ��b�x�on~��I�@;נ�'m*:�B�MO؜�� ���P�VQ�,i۴��4�`���O$��>N���fo	4˖LQ���h�����O �����V�'�r�'@RS>���D��1���]O��q�1?�7S�(�IƦ�RL>�O`C⇒TjZ�iQCǩ}��@���-6�<	ꇠU���d��֩�O�Ġ)O�ѐ�y����e�dDIW��W�,���O��d�O��)�<�u�i��	cŇ�F�RI�%�>����	�����?Yw�i��O�D�'K����DMfu���J.�}Q1E�W`\6�즭r6�\Ӧ��'@`�o^�?U������K�)��$�sH��%��	Ϧ��'2�'3��'��'���?.�ҘieȎ���s��G�1��4,��)/O��?���O�!nz�m�珄2j2����/\�`�Hq��?۴4ɧ�'�(�4�y2�9!�1��,��V|�5���y!�9�4U�I�\��	�M�.O�	�OBaj��V�=@����́�CF�ya5F�O^�d�O*���<��i����f�'��'���:g+ƣX!H"F��G{����dU}b�f��l��ē1���Y�ala�&V�@�������Q~�o��p�`�@�-��D�ںc6��Oxi�@[����㗬�D�l[U�py����?����?����h��^����1�x�ؐD��t������M�G��ϟ��	��M��w�n���;#�]�����DQ�'�6m���Q`ݴm�(�ݴ��$�zJ��'V�x5�F�%_�pW�K�a���1S��<�ҹi^�i>���Ɵ�I䟀�I�j���C���i���"�Ȗ�rTT�'�.7�M�e�r��O���1�9OT�a�.v��($DA�[������D}r�q��l�=��S�'m��|ad�Y5͠�!�ɒ�ZH�"�冤u��%�'�$�*�I̟4K�Q���ش��DD�E������@��l���N�8�8�$�O��d�O��4���<_����	w b�?�^�p�Q�������8�y$u���{�O��o��MKղi��}B�*�'�^P�`��cҬQ��ƛ1O�����L�#(�k�ղCN�OcP�=� d!�%Ȋ��2�� ��N�l@��?O��$�O`���O���OH����Ӊh�Xh@֊�i�QȐ��~���D�O���Ԧ�#�*�ݟ���ܟ�'���"*P1H%����(_0,p5H��K��M#.Oj�mZ3�M�'�@�ܴ����Z�`ٳ�ϙ3Z��G��y�j��qER=�?i���O���M�����'"�'��I�wa!C�f|��X+W�^����'vRX��Z�42Q�����?�������\e� �LM�I�Ҡ1��������?A�O��$l�Z8oZB�'Bq����H�lRs�� ؘa���v�8�W��a~��a�=���'o��Iğ杘}8� ���A�>�@�bЯ^�+��q�	���$�i>IQ-^A	�4�'Q~7͖;h6�q�ƨE�c�phUF�41tc�<�����?�(O�9mZ|�jT[��88r��4�Xyp8���4mɛ(ġzě���|K�-U�9>���~�qi�7H�%�A�ީr4*P(��K"��Y�����4���,����d�O`X�X%�,Yz�vO�,`�ĩ6m�����>_(���O��i��'M4˓�?ͻ:��dcF� �PX���x�+��iAj6��Ȧ)���O�x#��i���k���vm�4���	4��O��č0b�q�LSJʓ1Û�P���ޟj��O/R�L�C'�*`r6�xT	���Iϟ��	AyR|�L�o�O�d�O:��"
�0��5�ti�40T.�O�ʓ�?	�P�D��4Tϛf�rӀ�z0���paA;Br�\
 .	8@R��'���Ta[,
����Oͭ��n�$���?�0%Qg	x4�Sj�^y~Рw�N��?���?����?��	��\�ɹ�ztIc,�/X�0 �aE�b��ɘ�M3Ca_�?����?q����4��/U�`@փ�	~�i ��\���Ʀ1*ٴC؛�
մM������v!�<��t���Y�B(��wa6K�BR:�0�A��� �	��M++O�I�OP���O���O��)\���@I���TdC��<q��iA2���B�b�'����p;��'��M�%^�
�S���	=.9�g�RH�U��vHr�Rhm��H�B��l^O�Lhx��ͽUl.�&,�+ ^8u8���|PSmؼV�)�Iy"am��� kj@2�B�;f �\���ƨJ�d����?���?��|�/O>t�I2p���=^̱���H�U��rB�}�Ĉ�!�?��Z���I����4Q��BD Iz<��TiUjF���l�?�MK�O�m��P���J?e�Xw�IGp�x�FI�&*nxӢ�C��yr�'�2�'���'���Ӆ6Wؑѧ���MF��;�O�cP��d�O��릙��)�qyB�o��O���R���Vƪ���"�~�p�X�i�I�MÕ����眒N��&3OF� ��H)'Ģ(Q����Zl~�)���S�,���IZ��P���.}��Ryr�'R�'jb@Q�w�
�;��^�z'z�`���i%2�'[���M�6 ��<���?)(� ��vF6���G�0}iVH�7����+O ��e�v`'��'Kly�G�B�"��C����,�ʰD�k�(L�"��~�O��q��<~�'a�-³"�l	��C�ҹ\���$�'��'�R���O���Ms�āY ����9Q�*�:�L%�ƌ�'7M0��*���S�Ar ��"2�å���`�!
5b��M��i芁�Q�i���v0u�%�O��'#� AQ .e�\(P�mYmB�͓��d�O��d�O���O���|2��Ʒu\�$�5h�?0G�Ź񧜜j�����y"�'>"���'��6=�"Xq�W�$'�!S�]�_�U�D&J���͒O1����!q���I�s0���ą�Π�2+�:1N��ɿ�H���'�¬'�蔧���'�2������r�\0��4���'�R�'�"]�d�޴X+Y����?����5h�a˭b|`9��ƻ�C��<���?�M<)ck�?<x,�'�^ 8��:���k~RN�p���&c[0Y-�Oj���I5Yd"	2m 4��Bk@��d�#�i�K�"�'�r�'���(
7�M;z���s�[�6U��JQ��\�ݴL�$����?�q�i��O�N��3%Ba�Ei${�E�Ȉ^~�$������M��m�M��O�I����S���QŐ���ԕOp�ac���C�z�O���?	���?����?��Rqa��P�*�1���H2�),O&�o����T�����j�s�Q�	�=}�p�R��pk�����N=����Ԧ�*���ŞK�\+BMïzm�Xfo��U�������-O�u�P��?�0�>���<AF�Ϩu��7�<q�|9��j��?!���?Q��?�'��$���	ccm��dƇՐu80���;UlX��럐�4��'Jʓ�?1���M���W?N82.R��2�(p�	�#ڀհ�4��d�!_,������������� c���%Ɂh��,	�Ɓ�'��'��''��'h�P���Qd�(8�!t�a�R��O���O� o�u���|.�� ��4��$��hN�u°�й+��O\o�
�?�(��lZs~b.�� 7^8XsIA"�Ju�e�՘~��"Ɵ�!b�|�R�\���T�	̟p�`��^ٞq2��W4_���x��ޟ��Ioy�`y�\`�B��Op�D�Oz�'`�z����)+����ذ\���'�Z�l�*�O$O����`<I��ц{�$x���h��8G��<)���G
�7z�z������O�U�K>�c2#�JG`�7Rp� .���?!���?���?�|:)O�Hn�?af�	1���_خ$��C�!H���vCV[y�F~�
�d��Oao�m�h�
�D�x�n�1�
�J�.$�޴�?q!�_��Mc�'�"*D�}��y�-��� �I�ƿE4�ݪ��*cB�!0Obʓ�?a��?����?Q�����-��\�sH�'���7%����oڢz*��'a��)�¦睙V�$릆_V3"����F����{�4"ߛf�'��)�әY�Dm��<)@ON~�N�%A�D�{���<ɧ(֭@X�dW?����4����җH��M�#�I(t�VE0o�%;���D�O���O�˓\����/f�"�'��@g%��"�؆W�:��fO�V�?	�S��ڴ=����' ��*_Jt������"SBߴy���-(N��@o�#W����|�q��O��S��?�J�C���qH ��%��¶T����?q���?9��h���dZ��~�������� vI.���@�qړ%VSy2�m���]�YO�y�7��~z
q�'O�	����M�ǿiJ�OG��v��<q����de�\�FI��g�����ae��]F�T&�������'���'Z��'L�0jpjўVf�-�Y�Ԛ���ݦ�S�J؟����%?�ɬV'.ْ�Ә���4�[vd�X�O�l��Ms���>���,�N�Z(8�C��P�T,�¡\.MZ��d/&?q�E�O�*��]������F�
|Ke�#n#�l��L�v� ���O���O��4�,ʓ!��)��y2�E#��uhZ� �5
��y�i~�㟨��O��m��M�Ӳi>ΐ�����"_d �'T$m����	xț���h�� �3,���i��^�����t��K�톰^�Z���>O����O��d�O��d�Oj�?9)"lY�N4�M],&H,�W}��	�BشJj���'}�6M0�ā<\��D8`@��w�4��59�
�'�h�4՛�OX����i��Iy���'���v��䇙�f�-b�Qq���{�	Ey�O'��'�Nޑc���</94��ҡ9���'9���M;�G�q~�')�S�>s��9��N�Cpj�+E�U�c���t��I��M��iqLO��#O��I��
�P��SF�ԋ];�p0��(;����#?ͧGwV��ԇ��>��ñ���)G�yЂ�҉O�"�H��?1���?Y�S�'����?Miڈu����F��8��r��
�˓d����$�l}�Ns�j@z+�r�9r�L�dߞ�֥�䟸lZ8eܘ�l�p~R�E&9��ӱo��	n�#BJ@�|} `�[ -���py��'�R�'���'("[>A#g�S�L+���|ɤ�'!��M��&K��?���?YJ~�'盞w������:d*�jV;^�� �{�����e�)擉G��m�<����h���!*�Z�&��ˇ�<���̀�L���+�䓔�d�O��d1(�b��1B"���I�?�2���O��D�Oʓ["��C�V��'�bF_9 ���K��L��X��Сx`�O~�'-�7͍� %�pz��Ead��Bϫ$)*���8?2F�\�� �	�6��Q���䏶�?)��2U�� ⭝�|Ip���Ջ�?���?Q���?�����O�4�&��+[�%S4�Պ2r$ԃ�!�O��oچ҄���ğh[�4���y�Β�:�Nh� ҆ڤ|c�Ō+�y��dӄL�	Ԧٸca�ڦ��'ޠ\aSdL�?u��*���и���	���aD#i��'��I����	ޟt��ܟH�ii���?�v9�נ�6]~����<A��ie����')r�'��O+b�'q�,q!1��}�Z�0)��-6b�	�v��O�O1����m!a��*��<&>p�2�	~@j6Ϲ<����+m��Dؼ�����٣s~���C��W�|؉�n¾(���$�O��D�O��4��ʓ2��*Fd�2�i�p��L�#uRl)�#��y"�wӐ��­O��n��?��4w<@��:��XS ��B���P"�M�Mc�O��⅜�:�'����T��6F��������d��0O��D�O`���Ox���O��?�@�G�#F� J�{QыS؟L�Iϟp�ݴN��u�O�7m#�D�PDn�#@�;{( ��G�`6t%���4T��O��0���ig��-!;��؆h��O;T��A����D(`�@l�CK�IIy�O���'	d�xov,��f����k��K2�'"剣�MK���?	���?�-�z�s�C�+\�!�,�~خ�U���q�O.nZ��?�L<ͧ�J�2=��3%*���BT&��\� "��06Q�Ѳ-Of�i��?�F�?��U�+V	 !@�c��+@��]S
���OT��OH���<��irjB�$�h4h���B"���A!I ���'��7�$�	���i�.D�3��'l��"&'̬lv�z�aŦ�ܴl�Q�4�yr�'�81c#���?5��[�S%�V#T��%�
�DM�P�Ghc�d�'q��'�B�'���'Y�,�@q�� LLq ���X��c�,ţaD�O����O��ɶ|Γ�?�;.gH�	������6�K�p�z��0�i��$�>	��|�����S럹�M��'q� ��˷�P�Y�ł�j���'M��(�͕ڟx�v�|�]�X��֟�� &�I��t�ȼK�j!n�����Iß`��tyb�z�ZP��O����Od���hͼ��IR���"t����&��2��d���e�����-�Z���K�~}<� � �w����?i��͌�\C���d��n�C��>��Dmc�4ڣO�!t���E���@�$�O����O��d+ڧ�?��JU$OT��X1�ȘY&,a���?y�i�,	s�'mB�u�Z����d<��*ñ(`��0.�!UVf�Iަ5�ڴ�6�Mʛ�2O��$��	�0���L2�  ���Q)C��P"�����J)�D�<Y���?Q���?���?��DÙzАPcR:F 楫�+���$Wݦq+f]ܟ�����8&?���.rkd���Bр3�l�B4-��sb�(�O��m���?!O<ͧ�b�'4!
-	Pf�scr��6I^>^D��㨏Ge~�q-Ot����?Y��<���<�R���sބ;gJ��_1�	�pi���?����?I��?�'��DSݦ!�be��<q&m��S�)%%J�k�~�kW�z�4�ٴ��'�j�rԛ���O�7ԗ�x�€ͣ-?H��b� a��g�eӨ������"C��,;��YIyr�O�G ܶ@��������Y8�fO��yR�'�2�'{��'�R�)-0zx)��ʬW! 噃iQ-)�Z���O���VϦ]�sas>��ɹ�M�M>��ǓK����2O\�A�bߩ|��'�6mX˦)��i�.o�<A����=��
�}ڨ:AhϺ>(��Q���+@���H!������O��$�O �DЩ�"t(��{mtزF��E�r�D�O��n��̄@��'1B^>� �R�P]^QL'i�XԐ'�$?!�]�T�ߴcf��l4�?m0�
�I�Zh�v�	6X�xa��s2 ,� E
l}���|�T��O�HIH>�,њ`��k �^�7$�Ay�'Ɂ�?Y���?	���?�|�+O�,n��C���#D/۫v���`A�/M��1�Ϟy��c�n㟬ɨOlZUl$���G�
2-Z|�Rh��uΕ@ݴכ�k<$̛v����N��3*���~z��S�Z��]����2�v	���<�-O����Of�D�O��$�O�ʧ��ko�t!��<K�%3��i�~����'��'2�Obb|��n 9���7��<K�9�)��J�ƕo��Mkx��T�SAU�8O*1�S�[@i"w!Nx�*7O��ؐf���?��g*��<�'�?���ɣA�Va�5�F@�� �?���?������Ҧ����_yr�'W��$��A�~���`+=�89�����f}"�aӲ�l��ē����"�A�]� �,��T9J��'&��r��_<r�`����џ�`��'���Y��,0�&t�V�VPƤ��7�'��'���'��>����gl�$X1�H�g��1���cƥ�	��M+���:�?	�)ɛ��4�F�R�H�A�@�<_��s�3O��lZ>�?9�4Lf��ٴ����D_����'?�<���Ʊk`�rgG�N��ru�*�ĩ<����?!���?����?Q����C��!&y�O
��d�Ʀ�"g���t��ß<'?�I�p��i�[L�$�!��rK�u�O��nZ��?1O<ͧ����I���ւLZ���#� >m� +b�$�@]�.O��Q�엉�?�u3�d�<9r�Kh���'#��g���JgCK��?9��?y��?�'���Y����П�D���zD�a�¤�7��V#����ߴ��'����?���M���u�XKgKB�P�t���`F�,�۴�yR�'/,�b��?�
Z������E�F�еPZ���R�Z��Q�ѭ~�X�	ğ(����	����J��'K����0m�<&�h��
��?���?�ôi�I��O��z���O&��U���$�H�*��E[.���n�k��;�M�g�i%�+�^��f<O~��B+#Eƕ1��]0TBmP]ufy�b.��?qE!*���<����?)���?`jO�#b|�J��9��y�3�?�����S���Wߟ|�Iޟ��ON��Wj�
�@����������O��'o�7�U���$��'g��qd��/w���G��%K�@ց�U v�N���4�b@���0��O�$��L��" :�*A(��\$��O����Of���O1�.�9M�)]�%�Ri�u损|�R|�#胺z���R��'e��e�㟨J�O
�m�$3��A�NǖB�=�2�`��YPڴ0���LУu�Ɩ��Q4G�C ���~B�AֆQ��xS��k�˒��<���?����?���?����?1�⚐3��N#�,� �@B+ir\���-՚t�y�����?���?��i��'�2^��N�K?�K�CM�Z3<\1��H�?��426�U"��Y��y*���d�-S��7mk� ��k�q#ݨԩD�J{�a|��W�PK�"��@�	Ey�OG�dܯ)�:ap�$9 ��ji��'k��'*�I��M;����<I��?��lť"�HK�ܞO��bT	���'<��BǛ�Hh�x8%�����,��x��@�02�H�?<�'m�B�5�JT��,�7��埲���h�
��Φ@��8
�zP.lA��Y-Ӣ��O����O���*ڧ�?Y�ẺeJ���͝�(r�Ip�,�?��iw���&�'��k����]
^q�I��@�0�d�2/�J"��ğ�m��M�d��MK�O�A� �%��SMU%\	��+�7�:��*^UWV�O<��|B���?���?a�I�*Պ ̅�3�b��Ǭޥ{=|=�-O��n�&�,��I�h�	X�s���yp�(Ku��d��P������D��aY�4np���O�Ji�'�L�`Q�5�*>΄� �#+ ��*�O�	CE����?AU(;��<�SF�5�0�!)�'�j(Au�;�?I��?A��?�'��d��ө�ޟp�ZV�lk��lұ�cC6�<��^����?9�]��pٴmۛfAj�pɡ�ÖC�^|��&2�M!��
Y�~7|�X�	�	�d��3�O������;:N&h����*��� ��C=9�DUΓ�?����?����?�����O�
812�N�G��y!��H��O����I`d,?	�i!�'�̭�d挺DdH{X{3dPK������,��Fm��)X�k�7m"?�d�g�? �������<� � �@��v��;��?��- �$�<�'�?����?�%�+#Z���򂀾E��0��͜ �?a�����!���ڟ�	��t�OT�����Z�d�p��ϟ1W�T@�O���'��6�Z�%��R�����d\�9�b,;F������.W����ĵ��4��D����̓O�d�'D؉��!sN���U&�O��d�O����O1��ʓÛ�Ǆ�-ޔ ��B�]�fRbG#���Ң�'(2�v���L��O�o�:|x����i�3)��t1*C�En(���M����M+�OpX@������<!��׎mEl��!6g������<�.O��D�O~���O����O��')�H!�.�
�y)`	
�xn&s�i�R�QA�'��'Y�Om��'-V%2���aO�帠ϟ�N���o�"�?9H<�|:�!?�MS�'H���F'׺@Ä�W�v@ !��'m����l��k��|�\� �	˟ ��ፊ}".�9S!�n\�(H�F�֟�	؟���Ey�wӀ���G�O&��OR���ND�F�.5��� "x�#�%�I(��DP��H��ē�&i��h�TȊ�JS�e����'��� 5M��oȹѳ��������#�'���1O	h�T��牌�S;�j��'���'��'��>��r\��Qb�5�ι@B�Қ7yB����M����9�?Q�&㛆�4�vU��E�b�dę׃:,�r:O4=m��?Y�4Ns�4�ش��D�:,����w]p��a��WD�|�"�-���S/.���<���?A��?����?ys��>:!�[G�8)vb���O�6��_ͦ	�E�My��'��O^2B�)Oxpn�bd�� "b�h�h�#��F�O`O1�t���k���uz�/�>R^2�ܮ`!�����<I�J~����:����d2h�t�P���#m�b��������O����O��4���#w��А'��^�^:����!8{������ry�jcӰ�p�Ovho���?��44���"c[�[��	�����$;&@��M+�OX�˗��$�z��?����
*�e�B��.�5av��V;O����O����On���O&�?��b��z��h���sG��ٟ@��ɟd�۴l+"��'�?ᴶi[�'H|{p!��1�pj�H�$�9+��!���O���O��Ԋ�i���/���͘==�X<���Q�hTr(�߼�����䓙���O>�$�O���r�+.�e�1���e��ǟ��I~yr#i��
E��O���Oʧi��8@��'��i1.��T�d�'��d�6k�OO�S"e�މR1m�4t9���r���m�n<R�] ���AׂX}y�O��Ib��'�B@����"�٢��~���v�'R�'�����O��ɼ�M@FXOA���$�R=$�nU���Y<u���,O�oZD��!�����MKe��5��P��\5C�JM��o�Rb�i�2d ײiO�IK���%�O��|�'�ީaOS�X�|����U�&��K�'���8�I�`�����Ic����rX$9DI�B $���T#�6��+�.���O�d"���Or�mzޅ�B��/@�|Q��Қ^n� �N �M�յiW�O1��,K�Cp���IZ2����K��48tL�<Z��.>D���p�'ʹ�'�������'�2	�3n��M���LR�if�'\"�'lbV��!�4qL��z��?i��r�}�rhU�r�����oڃ	��`�2
�<!��M˱�x�%H\�b!O��w� c�ֽ��䞤2-�p;deK�~#1��|��{#��$ǸP�v��ƕ4^�4��A�žN�(�d�O�D�O �$"ڧ�?)4�>j3@Qb7%\\(ma��?w�i������'#R�l����'X<x� ����w�h�0*�H4Z�I��M��i� 6�W�`6$?�G�h�f��	�ѩ�B�
�+��٩%���I>1)O�i�Od��O���O�P����;OO�r�ܪ
��A�	�<ҾiHĸ���O���.�9OZ����Խ>I�5���Ӱk*�Б���X}R�y��o���|"����Ƥ� Lv����2Ԓ���T�n���a!V[~�]��y�ɮ6"�'���R�nlI���f�:ADGB�_��H�	ş$�I��i>�':�7�hf����%y��g�N��a󪚀h�������i�?9�_�h2ڴJB�i*�`�j˖ Wb�1(մM3�	tK��b�֑��`�(��	5��$�G��߁�c�'%��0��u4aC�ko�|����������I�T�����+�,,�����:bHQ�`g��?����?qb�i�dY�˟�8l�џ��'��I� ϕ�b$���B�A��ъ �8�dĦ9ߴ�����MK�'#Bʘ?��h������
�8� 8�P�Jϟ8z�|R�|����Ο���GN= m`G�[d�C��<��Syb�dӴ��1g�<����i��S����eP�5���8.@�Ɍ�������������|���?��(�4�$�a�ʷx��qa�-P	4ƶ�Ѧ�����D�� k�	?D�O�)�0�U�?������Y5Uh�H!q�O��$�O���O1���a�V��>W����e�\�9C���Fm��z%�'YR'pӚ�;�OZohن�YuI�]��@M�n�1��4%��6�'n��f?O�D�3J�����b��w����� �:0O6�1V�ٴ�r�ϓ����O|���O��d�O����|��2DJ⬒��ښ7�dJ��6A���U��'bR���'�r7=�8	�bO�9r�$LD�w\�<�p�[�	*����|��'�JQ���M۞�� �Y[tfT�CɈh5인Y����;OJ��l7�?9�*2�D�<���?�D�^4%�Q�e+K2t:��H(�?���?!����d���I�f���X��� � ��D%:'��H�)���`�2�	+�MKS�i�S���B��99=��0(�G;�Yi��p�x���𨳐Cи%2�bV��Oxdj�L���BWƎ&�t\㥍C�=������?����?���h�>�$U7{��80 �ZbĜȠ�K44�@�ČҦ%���8?ɰ�in�O�.
�4I8�AvA�.����*^�?�ܦ�!�4;e��-J-%�V5O���I+�����'3I�h�C޶sp��)A W�u���ʷ*���<�'�?����?����?	P/IY�!���@$���[4C����$Dߦ���c|�`���X$?�	���J�ٸ|V�au''1�3��D�O^7��X�韼�	���-S��)p(���Ɯ6���͜oؾ��P��d��&�9��FN�IQyre��G9
̃4��halLq7�WlR�'T��'��O�I�M#F�ƫ�?7%�g��`3��]�wʂ�@��?��i�O���'��7m���Dm�^V���Q�D@s��őp����	
9t�7�%?��%���I��ҘϿ��-�i�m����Us�BV
��<����?���?Y��?)�����[1vAٲ�@y�fԈƥ��$HB�'��n� R�4�l�dM���&�t�T�����"G����u���A'��!��O�O��k�0^�f��d���֘5#�$9PNL0�zEp��� G���q��'�� &��'���'4b�'�(\�A∂8���,g����'�P�Tbܴ2ޞ��(O�ĵ|��$�E��}z�
A��N�8i�~�!�>90�iښ�3�?�"`N�y�TlP�9����(n�tx���H�>喧�t@I����|bn�{`dS�NL�7�rh)!�W�c���'�R�'c��4]�T�ߴl�$�����>DTh(@7e�:�|��taʪ��dJզ��?7U����4)d���+��0ًCJʳ*ઉ�U�i�x7�_�U7m:?��K���>�	+�Ԡ����Q��t��udX��y�]����֟������I����O�P8���U�Z[ވi��[��C�mӬ��G�O��$�O�����DH���݃@N6p�pE@�W����e���$���4>���5��	ɓ}��7�s� �S$n�XmHB.�7�6I�p�P�ƁU %��i�D�@y�O/X�)����O ?F>�x4o�1<�R�'���'�剩�Mk2���?a���?���� ��Y��\o>�Ec��H���'��� ���gӬ�$�؁�/��Y��H[q�<E0@It� ���l(hK+�|������O(���D��3w,V?6����/[�BՒ���?����?a���h��ė&%w�M��<t_�RV�[�C�\�d���=���KUy�sӌ��]�ecέXcK��W~p11�@�a�b���M��iS2Q8~�����X1Q��0`���眠a�J]�ri�2�>@����5WuF&�P����'52�'�R�'�Q�4��t쀰u���q[؉X]���ٴ�f�����?�����'�?�D��
|��+Rk��Y���C��"�I��M���'����O�� �e*�l@�e�i࢜HfKZ6��B�_���r-�*j�
l�	jyb*CV{��kU�×[���T�X�y�����\��̟�[yBxӞ9� O�OjP6L܏���8 ��er��>O��l�S��t?�	�M���'�L�=_p�;F�Ĺr"A�1G�	l��0!�i�����e{U�O�&?	���K85�F�L	[ڎ��@�=��	ß�������Iʟl���Oc�\;�mI�$f�I��J%W�0��s�'���'� 6�xp��kț��|�b��۪lb�O�!vP����*2+O,�l�*�?��7���n�W~�b��a�R	�CKZ�!ĩ��PRTq�G�ӟt0$�|�W��	��	؟�3��՜`=`����0qS�I����Ify�Ge��0����O4�$�O��'J(�X
�V:�L�!�3k�u�'��Si�FE�O�O�S�C��T�탚wq�yQ�ǂ�rw"�8����z�ǘEy�Ok>��Ic_�'�|(V`�q�V�%��0
!n��'��',b�O:�0�M�瀋�Tb��U*"�(9�p��7��P��?���i�O�p�'��7m���Qk״o�B��f�<���O�7���6M#?�2/U-Q֠�隁���x�ɻ% �@�N��`�<f8�D�<1��?��?���?A/����I��bܩ)d(طG���!]��D�C���	՟l'?�ɻ�MϻV�x�Ԃ�'��H�!oT�R�d�h��i�^6��|�)�l��m��<I�h�
\C@�^��&)��<Iq��5	��$��䓈�4�����L8Lx8E Y1,�Ęh�T�/K����O��D�Ov˓Z�F�H�zA��'Cǂ�i��p6��,s�h��$b��s�O$U�'��6m�ۦ1�M<��̥k�܄p`��Dd�DOZA~� .zE�}�t����O_�a���1�Nų\�]���i�x��[����'��'�2����J�n��L�p	9���43�`�Q�^��4ufr�.O<nZK�Ӽ��T���*���+c� ���<A6�i��6͙����&�DĦu�'ˤAB�A�?�
b�K#��y[����R� P� $� 1�'��i>�����T�	ן���;�vQ��$E	jpH���� >��ȗ' 7�G�V]�d�O>��$�9O���⥖�aD0p�B��it��`��[}"�aӴlm����S�'O�L�� <i�5H����|+%@Y�<�ZH
�)�Y��ɳ ��݈d�'�>�%�Д'p*@;��({>j�H�՚8BE$�'A�'�b���U�|K�4}  ��8,��@g��a��I�!��:~��͓)0���d�M}�ijӪ�m�M�%���+�(�0��ݸSJ1���k޴��DN�P\P���øO�wNqe�X+F)�Ir� ��a��yB�'�R�'0�'O2�IͬW��$�6e��:h�NZ!Y`���O����Yr/l>e��6�MsI>��DY� �!��G��ZE�\�{H�'�r7m��I�	;Z7-3?��DʄLR��w���I��'��� ���O0�J>(O����O����O�}�V�X7d��l�r�Z .Ŭ�2s��O���<)��i۴D"��'D��'���U/ݜu���хL�M�a��I=�M��'�������0Q�a�cA�O�B������D	�E��(%�5[d)�<�'x����%��Kt�����=NZ�l�H�r������?���?��Ş���֦�pDС&iQ6Ĝ�tTb���훲b�'�7�=�I���DE�EA2쏕�`y�3&��\�6�Se�=�M��ir刖�i��$�O�h����ڴI�<�Vl��]�B��&��3E�iZ����<�-O���O����O����Of�'&W��X%� ������X�h��3�i/.dKB�'���'M�O�@u��΋�'|��t.U�n��a#����,�|�l��?�H<�'���'H��H��4�y"f��Hs��@H�w����f��yRG������k%�'��	ɟ8���/xv ��J�=L��@�Y*]���	ٟ`��ş̖'Wv6����&�D�OP���1t!x��������P$`�>����O4,l��?�O<q�FK)[���h0J�2v?t���D��<���4)� Z�9NL�3/Op�)��?�q��O���s� �Q*Ď3e��;�Oz���O8��Oꓟ�ä	U���ښg��Pb�]�k&�R�o�)^ˈ���uDMğ����	gy��y��Z�q��K���4Z�
�
�*��y���^�n���)�ܦ��'�
��H��?�"ލ"�t(�7+Z��Ha����.a!�'��i>��័�������"'�ܱz@NM*LaN(ТJ+^�@�'��7���:TR���ON��5���O,\��\4z�D�3�^�&S��T�Tty"�'|J~�`�A�M���%�;\@1������ݣB+����d�3;����O�˓d ����:g��TI����d�VLY��?����?���|�,O0�o�32s����6|؀��g\�C�5�ca �Xǆl��6�M��F�>i��i�d�D�v�s�g�e���P+�+ڐ��ь�ze�7�2?a�BW3Q������ܿ���WD��Ř���.p�ȓ`�N�<I���?���?1���?!���@��p����0�K	[Q2ؓ"�,R�'�B�k���@�5�H�d֦�%����d�8P��ӿHy�q�5��ē���k�O��d"E����w(h�̌`6�(hEN��sg��f쪶�'� �'��'���'K��'�H��f��x�T��3�W�
}q�'�B]��
�46�nm���?A����Q�D��pb�� ��i�#��I�����������S�dj�)7�p̉��Ƿ3װa�R�A�`���pc�R0N|@��Y��S#H>�m�u�	���F4]v�(���]K~��I՟L������)�sy2-m���)��ÿD�Ix�� 8�uW��>�2�^���x}B�u�����:��E����F-`�S���ܟPm5K��oZL~2�
�KĨA�Ӡx�ɟ����S&X��Z1BŘ[X��	`y2�'}��'���'�"U> 2
ڴN���k̆692��E��M;F![�<����?)H~�9t��w�0�+��`�M�b,��<��mc�2�n���S�'D�ta(�4�y�_3�T`��KT܅Cp#��yb�K�&ZQ��;6�'�i>��	`�`�x�d��6�X#
޴+٨�����Iß��'9�7-�-]����O��䑗Q���A�ml�ja�ԍo'�P��O�m���M��xb��M0N�"eѡ/��1i�Չ�y"�'eM��8kZ���O���?�?9���O(����
�o|�Q��R�e�l32h�O<�$�O���O��}���+t�}�@�2s8th�d]�� ��#�> r�'��6$�iލ�$� D�Ȁ[���L�P
e�r��P�4@ɛ�os���P0�vӺ�	�$�$�&Q��$�Pv��A�?46����R'��%� �����'���'�R�'� �+f�m���h���BX`�!]���ݴ(z����?i����'�?i4[=T���:��%7����-����ɹ�Ms%�'߉����O���X��pi1*ȣ5�ɹ���8:$���B�	��剳"��0V�'\b�&��'�"�pR����7�.����'qR�'������V���޴%O�;�bך��VJ�&�҅�`�Y$��3��7��v��[i}bCh�&��	��MS�F}���{!m��0�lEb��ɢ1l|�n�x~r�Y&�X��ӻ��O�+�d"��ցBa՛#�^�fL��Ot��O����O�� ���d<�7̒M"nY0�f�P�� ��	�M�`���|J��}��V�|���@��a:W�ǗK�����M��O�l��?�SO�v1l�b~ҋ�=@@0�"�ͽ~i�T�����'>d���蟌��|�U����ʟ���ޟHx��_�j�2,,��2��ɣ���ß`�	dyr�^��Џ�O,�$�O��'i۾�B�C�2��$�@ܯ#���'Ք�l'�&��OzO�3� 2��!Ĵn����\;5����㓊W��A�C/;�P��|�s$�O� O>��j��%�r��.۱S���R'g���?���?����?�|:,OԤoZ�$��*�Z|>�i�nݱn�D���HßD�I�&�#�R��>�u�ih�p�3ǜ"�ly��m��$m��O�7��>g�6'#?�SN�k���C������D�k~�b�[�m��$�<q��?���?I���?�,���*<+pb]�@f�_,�<P�Gɦ�s!�쟼�Iџ$?�����M�;4��8ɇ�̫\x�h	�lށ�N�Av�iYT7-�^�)��\���oZ�<qρ����҄�:5s^�l��<Q��X�/Nf��T��䓭�4�6���.B�li�#ض<��+1��8�~���O��D�O,�?����q��	�Z/�E:6�
�i"�Є��`��[��	
�M� �'G�' ��h�L�:F�*D�&#�$7:j���O�U���8M�ո-�I�?$�On�
[v��F�D
h��I��S>B���'���'�B�s�a�qB�y��8�h��D@ -<�ݴi�)s,OP�lZB�Ӽ�g֊*��TY��۱@L�庇�<�f�i��7��O��	�o�n�EL�᪶��T���/߼�i2N�� �bЁֆ����4��$�O$��O��$��fyi�����6?6%At^�vp�N�6��7;���'����'�R���U*B�
-�Ә9���>�v�i�<7M�O��F�t T�=w��X�K�{��E��9Q$�Ä*؉��$
&fr�D��w>�O����$R�S�9X��V(C=o�����?����?���|b)O�o�f����	1`J
�tŔ����0�R�a.批�M��b��<���M[�Tc�<af�]�X@ʭ�gJ�"�l�/��M�O��@�����w�X��eHBl`иJ�E�,�2�'���'��'���'%����n�����f�=.��x���O�D�OBplڌC���':V7$�$V�\�ED
� ��բ��k�|��<��i��7=�ȹy�`h�*�Zi\8��L�0�0�Ҫ� �JIh�!��(ɸ�$�1����4�0��O��
5*
}ɕB�("u���ǏÐ@�j�$�O�ʓǊ�?9��?�(�H|s���[7��R"r�ȤJb�����O��n��M��4����0S$�*zO�2t�Dh����e:D��z ��O[�i>)���'���$���Sl�}`��r�iʲ'TXP����㟰�	埰��ğb>��'�~6�_	o��q��۠n%���`��>(R�Ʃ<�ǳi��O���'o7�V"#��,q�)�;	���-�,�Gq������B~6-#?��ۦ1��	%���)`�t�3�K���r�*�y�\���џ����� ��ȟДO�� ���=H��Ē�o�7�
) �gӀ�)�O��$�O���$��睥=�h�̀<�Xa��m��� ���4?���'�)擰d��m�<��H�:����mA,'��s�kY�<��Cۯ��������4����_��ʇ,�X� � v��S6D�$�O����O��=��VIƹK��@I@$��@��3a͂�8E&�h��VU��C�����lZǟ�'�P��йv��5j�h޹�LS�O e�����+��Qf�G��?�f��O(�1�a�0,�t|��̢a`�B���O,�d�Oj�$�O��}���L!hA� U"iWܵ��AI=q:��I�^I2���$�ɦ��?�;4H��0�F�k�Vѩ���ʰ��O���pӴ��KY�7M&?�i�;y� �)�^ ���d�؄R��aw"�!K�p�M>i/O�I�O��D�O��d�O\A��a�9���V�U0_z�}�W�<�ҿiOƠ�3_�,��X��
�h�pl��4̸M���`�T���P�4��ߦ=��m~J~*A�;�^�9��\����07K�(�t]��ˆ_~2n�0s<���?��'r剅��R�!Y l�^�J!;��%����d�	���i>��'��6���{�(�D��){���	�{��Y��D]7!���ۦ%�?�V�\��4ܛV�'�\�jT�2
��薭 ]���RG�{�����`��#�V���9�p��lI�R��E#P�2D����3O��$�O����O��D�OP�?��'�Y!^�r4x`��hq����Iǟ� �4�x@-Oz%l�I�R?�1�F
 -�nmBG+��Icy�G}Ә(lz>1��LA����'OH� ��th3���:e^��KՎ�	��x��0s��'��i>��ퟔ�	�8�YOK�=*R䀠�U
���IڟЕ'�6�!7����OR���|���7I`,v�*����C�w~'�>���iV�7��O��~���!34P�����ą��N���l����;��������';��2�gۥ
"XH�T��M�'�Y�w��ZQLӋy
�}"'.�g���ئثш�ye�1^�>��TL�E��[��|Rn��|
���̅धB���O�J��HQLhpc�ҝ�J�KǄĸXBޤ)@ə/�A06!\��}k�gK��ĉ��ci�H`"��߲Ljn���̒Hn�q�

;h�&��g`D ?�:�����6}T�q(���1�^��,�E�ݳ���(� �#nW*+���)�I�!RC�9�GA���QCA��5l�� 4�O�@Y��:D�7Z$��ZC��>�*OJ��0���OH����^�>-��Z� ;d��W#8XÀ�3���O\��O�ʓg֬��W=��tKw�{ �S�@O�Zഅ�D�i����X&�\�����TCQg?�!M4vhT	��F�$sQB@n}��'�b�'剶3ذ�y���M�O<8�:R�S3�*��+��j�nZǟ�&��	ǟ�#l�d�S�? l	�m:�J��K��I��R�iF��'�剥SO��Ү�����O���O�y^�\�G
�9�Lm��٢G*Z\&���I�j�OCS����)�	!��[D��:�M��e�3�M3)OV��H�ܦ���ȟ����?���Ok��p�1�BL�^�pQ(������'��h�4�O|�>�ǉ	�(;���#H#i2r|ЍqӸ���������͟p�	�?y!�OfʓVLK�-yޤy!F�4\I�e�MS��Y�?&mYT~2�	�O�l��)JLv�E�F��lňQ����ϟ����	  ��Otʓ�?�'@�P`�蕍	^r��[�pm"'��̦��f*?	�/��w2�O���'�R�Ō�z�{ū:(��$Z�ꚯ/7V6M�O�}� ��^}"S�4��Iy�Լ�Ī�,�R$b���h*�Q���G}���,n�'���'wBY�4q�G���<4�J�"�$�s�.5�$X��O�ʓ�?�I>I��?	Fb�7S��a���>4�Q��e O��
M>q��?������ ���'+�0����w�*0H-�S�ao�@yB�'��'�R�'N���O$]�R�ǭ�l����߃ 98e��U�$��ԟ���Oy���3X�>�'�?�R)J�Nɚ�x���&,�"�+�`�	M:���'l�'���'�h���'��1®O�ˀn_�/n��!�9j���i.��'��	6f��[O|B�����@H7'
�L�LA��ӛ<�N8$���'��M���'|�O$���1%��BA����[�D�-Y$�6V���g]�M�DR?����?eK�O&!1d��	k`)�bN�ըE�տiG�ɩ(��5�����'�򩶟T�̍c�`q�gC�`�N��s�l,
g�̦Y�I����?!�I<�'gnRy�@&U�Xi����J�B �J��i��'1B�|ʟ�d�O��Y�I'��1B�]�ū���ܦ���\��

��K<�'�?a�'�Ƞ!!���z��2q�V8��P#۴�?�N>�GV?���iZ8�����VH�QC@(a �O�zc��<�*O����ȍ_����cF�.�Hd���3 ��<�����O�����$FF�	�aӀ;Ǆ|k��NBظ˓�?����'Ur�OJ��)�B�4��p�ƚ&�`��i��+�y��'��	ǟtBv�_h�UA�(Y8M�QG�5"��wn�Φ���⟌�?Y���P1$�&�A1�,�2���k������	���?�*O���B�N�'�?Q���Tc�`*F�Aq�1"6J�)s�����O��>��%��b-7LQ��W��fu��j����<���`XJE�.���d�O�����U�3G� �������-�h}@�x��'[�	!F5�#<��!q���d���!�h�j��Û'JH�l�]y�,��7��6m�O�T�'u�4�-?�/��b��X���S���d)�ɦ��'�B�':L�������=���򋛕k�IC���M�	^�ZR���'�B�'9��%*�4���a�$�/0ǀ82p��6)z�HEA���۟`�	o�)Γ�?��+
r������6P�����bś��'x�'襃��8�4���ĥ�,��OF���$��悰v@�ԛ�yӦ��4��s��'W2�'a�OƟ{q%C�'W  ,�a�@���7�O�iۖ �D}�[����|y���5f�і~��A���Ɠ�yؤ����DA�r�$�O��D�O&���O0ʓE�"5P�ă��H+�`O
5��p��d)I�Icyb�'A�	㟬��ݟ���*�5-<M���(�
��f��k �I����	����	ßP�'�x��@�e>���d��O�j��E��8s�51)bӌʓ�?!(O��$�O��d�^�ȼrd �p�ՒKc����1.B�}m�̟P����|�Iry�E31���?�1Ul&e列(
0���b��-pb�l�����'�'�"���yrP�00G���1�~d梇�US���O&�	��'[�����~B��?Y�'#cj�����U�� ���N�`0R����П����0"���'���S�6�4���*�!$2�1�nM%\��V���r���M{��?�����^��ݖJ�.�9�f�<R�Nh��J[9+�@7�O������:OP���yb��U	��T���>iN�8v��0����
OX6��O����O����K}r\���J��1۶�2L��*(!�d��;�M�b��<yK>)��T�'���ru�M�]��e;�Ȗ:�-��zӢ�D�O<�D�]�2P�'���ڟ(��z��p���>��N)^do����'t�j�����O��D�O�`�KS"&��DG�<Mpp!eF����ɈP���K�O���?I/O������e�����ȿv�L��d]��Rh���'5��'��^�@�Y?��p{���q"�M��d]_�,�*�.�I%� �	�8"�,V�l�ѢₜO�����%׭
���myR�'���'��	 )p}��O�,�ZPhX��y�e)K�`�ؑ�N<�����?�����(*��Z���勤K��k�]�i�^��[���	Οp�	oy��E'{�$�.xIU�QPg��AT!ġ`�9�weW榹�IQ���)D~��=! �
+`R��c%�f�΀0�)��)��ş �'�:I���#�i�O8��ExXA�Ċh�4��ϯ
k�D'�p�Iޟ �%fm��$� ��!|�H�ʈ5�����Л������'m�,�dv�@��OT��O�`�Z�H��Z�7%�$�oռp���lZԟP�ɳ*���s�IU�g�? �Ų��2�0�yF$N2W�r��5�i�xJV�s�����Ob�d�t&�����,�L����S� B��f���ݴ @���䓘�O@R  �?4���%�A0�6HYU�T%#�r6��O��D�O�vĎN����P��Y?� C��~���2�J'~�)$��ʦ]&�<��t���?����?����"?����1*�M�T�@τP&���'��]�4�0���O��D.��Ƭa�jL$p0�����q6Rt��Q� ˅�h���'^��'^��*6�  ��p�E��f'��q���%���}�'��'v�'a�� wX)�V-ٙTha���yW�\��韸�	\y�B��=Y����}�E%ЇZ���:DV�l6t듨?A�����?I��ZSZh���K�{3�N�zj<h8�Ǌt�$�A�[���Iџ�IZyҌ�������#�)o��𑳰
%o�$A�n�ןX$���ןP�D&l��O*P�ǁ1~��8WDۖOth�K�i�r�'���@O�]�H|����z�AB���u)r�X�\[5�w�R8/��	џ��I��h3��x� %�|�� հI+ ̀�G�~��ƒ,��nZvy�ǩ0\Z6-Z`�t�'��D�%?�5	��c8E�Q.�}���VE٦�I�4�6�]���'�@�}D,{0
݀c@[�*"4��Ԧ�0�*F	�M#��?�����v��8�HY��*ƞ�^u��j�>q��=m�)x:��?)����'𬉀eC�&]선�o��{�����i�����O��d��Y;�5�>���~�,�X��=Z��g��BL��M;N>�qE��<�Ok2�'�R,V�y��X�U*n�R�	�Z<7��O����Am��?N>��Lv��aC�
�-N�bP�S8:�i�'���c�'��ܟ�Iϟ`�'MVe;"��l�p�B�S�_�N�@��O%#:�b����J����	�=���3��H9IĂtc�	ӋO�9q�������'��'�r^�*������*Ԝ!�8Ɉ�H��Rs�/�5��d�Oأ=i��?�z�"�)C S�N�aH(@�a�\�c��p�P�iaR�''2�'��	� H+H|SH�#
� ����z���4B�f����`��H�ş��	Z?��e˛caj�3�E�/i|m9���ɦ��	����'����2�-���O0���$�%�D�Qr�hQ�g�<+.̒��$�O��sM�O�O��
z.����o<X��!���@d7��O����C�<���OH���OZ���<��O���D�T�_��0�T��-Kn�nZ�������""<����J�<���Re���$��<`2C |4xHj,7h�t�ѬB$������Od�+�Ɔ+�A)�U�i8�-W"O`X��"�GvN��ү�>,� �c�:w:��5;xI�zSt����5i��1���6Ś	p��&3&a߃�*��wD�2(3��ґ�\�#!.m!/Нp[�|#r��"����Sa�	�z��F�<4�}�[�7	~�H��Տw �8�p�hF.y�%�٢si^Z��uG@���O����O�8���?�����X�
(���f�1L��ѻ"��/\��s�G48�=��R�u����8�QJQk��^�+Q�dZ�I
F�4�R�u�t)��?E�*	���Z�M*�̚K�'��Y�lY�e��ɡ�ǃ���Lۻ�?����hOL���4
�xp�ph	�tK��Q7$ D�����2xe,t$5E��a3W�<�Ɋ���<Q3E�����p���TH��a���ڴ�_��ɀU���쟄�'0{��!V�T�*� M���߳�M���Bk�j��q��R��D��d�6"\Э��Ϋ~k�-�a�<�б'H-^����Ϟ�5�����'�bxa��?�+O�4�ІE�	�!���0��h2��$#|O��� �R�2t�Y3$�*
sDi��ORPn��Z��;�m�=H�Nh���J3<ư�I~yr'.5����?9-��؂���O���ɛ>H��+2�`��mKT��O^��(ǲ�q��S�T��i�C(�'�򩁹���`�E4������@OX1��+9�9����H�0��V�Ǯc�l���	\�0��}�>qG����j�O��"�tN���ED��Jz���(O��y"��]�$((�ݯA&6(�C$���0<)�鉥/:��I7�����6�س��A�޴�?���?����5Kؚ���?����y�;$-��q&n�bQ�u8�˅q���3�D��W�d�|AD*�aZR�g�;����(��lC�%��FT�R�T7[���	i�0���|r�� g��+V@-�#0<\d����"08��L>B�^@��"�A8$��	i�<	���P�@���ޭh�� ��e~n4�S�ORbY0���:�ֱi��Z�g��p���|o��c�'�2�'��xݩ�	�ϧY	ucC��/Z͆�K`�G���9� �, ��A��n�#4�^XHϓ)�x�He��*`�H�JΎ�\��T&��b�.3���2d�> R�a�.UR� %�US�b������������?9��tc� ��m U�1P��h'���y��Ř"�TT���t�@�S����'�x����F)l�l��4�ɾ&�u3�e�R����f�0eS�a�I�<�����$�	�|
$�ʟ�'�� 0A�"HS�}8��[([0(��';��،JO�~�l��ʃ45�E��e��p<�.��<$�t���4���C#���<ލ�6�8D���"��1���Q��"MU|�X��6�dcݴf�1��$�2&�d�C\�z��1�<1Ƥ��y�f�'�?U����O^tQ�$�5�8u�Fo���� ��O����&Y����.�|�',���3a�1>'|9wj��V�>�
J�$��h8�S�'l?T�8�([Bp+f)�{�ŤO���'�1O�>l���]�BD�2u`3(���"OJ0����N<�����`���A�'��"=�fD�g�D�z��23��T��� nǛF�',"�'��x8�-XR�R�'�>O��	�_�X�c��2A,<C�L�-
81O��"��'t)r��]Vl{��N4P�0YX�{����<!�-M5@La�a�21*�%S��;��'-�%s�S�g��?q�lbfl�	n��C7e�$��C�I ��S�(4Y��*�@:�#<?y��)§?�����W*]��mA�ō�x���,�-&������?����y��`���Od��!�5b��B.��/��'�� ԭ0�(W�\�-1R]�%��`�,�ƇN,e*C���/1�1d#S�.y�q�,��J�NI���O��$̮mj�C#�7�F-�R�5g�!� -1_ƈA��J�V� a�e�Zc�1O���>A�۸<���' ��O�2�5��׫M�^Ar�؃l�b?O~`�$�'��:�0�Ұ�'��'F��1 CH�jp�� P��Z*Ǔ*�H�?Q�����e�So��1��}X
�i8�����O��O*ESsL��dfl]¶Kں-()�g"O�u�`�kLι#�+I|(�OJ�nZ7KB�D"�`�
L��Q��Xc��b+�3�M���?y˟8�cu�'N�� ��Ҳ6�zKDᇴjQ�SD�'2I_�rp�T>��tH�V��͑�$�-�re�OH9�`�)�S�l0��2��.J���x��V�8�d�'�(�������O+dm��������RN�f�	�'n�H��I�9��@��IЬQ�ÓG���|�7��b�ܣq�ԅ�͒@eZ&�MK��?���sl��� �?����?阧�#G��8Lxd� ���Lv8�k`ژ�'1�Jϓ+nX�{����o��@��#�Cr8Y�=���xx�(3gG�#d*%B ?��H�#�z̓<���)�3�$J�ue �`�@�0d�����
�*9!�$'=xT��Jp� �3G�͔R��I��HO>�D�H�`��0�c���8`�.V��,VOΟ��ȟ����uG�'L"4��YSa����ޑjC�x�F�D l%!����4P�!w�K�ah�P�u.�	h�ܫ3O�!W���`d1��I
%Ȉ�7���'��'���'��O���W,ʥ��Tn�s�2�H�"OliJsHC?lX��l w�j�4��_}X�����M���?��c�iG�Mc��U+PDA��j���?�'���
��?��O t�BŊF�'6Y
1�|X�e"!#
6���![f�*Ԛ7�Ky8��K�K�[iF��1�Ї��L��d
�tJ��`E�tj���
��x��H(�?�J>�ň�Tm�A8ֈ��~K���LX�<��=ge4G�ń8�`�B�LOQ<qw�i�� a��7�Jqn��JwT�y�gގtqV6m�Ob�D.j��ğ��������!zU��&X��Y��ٟX�	&t�R\��X�S��O
l(PE�-(�f����ݎ=q���!�>3�������V>`r"~���
UBY�P�����/�o�D\4:r��ɑ+@L�kA��nw�}�= �!��kz��t��\ъQ��k�� ��=ͧM���tA	���	��.;*�>�ZwHؖ�M;��?Q�&�����?A��?ᚧ��pdA�)�ř��"7�$���#��'�֔��HW�#Ƥ�mc�e3@#_�L�=��&�vx�� ��,�F��g*X&.�x�å��I̓-�x��)�3�?�$`��9B���
�*E�%�!���_#�����PXf��v�-C�����HO>I��U�a0����+#�����PA��+v�ʟ�������u7�'��>��5�dI�
�>�q`���H�B��1�Ĉc.!������ �@���
<�@���E$[=.)+'�\��*ߊF�T���b�$bȉ�6��A���d0�O�U{��S9Kf���@��̬Q5"OH)(�gG5T��b�����C��d^z�2�x����i��'��dPäј�d�X!aU?�F���'\�ֱr�'��I�-�j�Zp�Y�Ɋ9bw�fӜ�P�#��s�8���VD��q�'�-�q`���~|`f(J%D�cؕp;l ��!���үZ��p<�A�ǟ�$�PZF8l�5YQn�?z�*D���G��������9J}C�)�l9�4'||���L�x�΁��Ń��U�<A�k�D�V�'b�?	�P��OD�ZУ$Dah�@��:ֶ�Z��O��D�Qa\�D+�|�'�"�;W��,�p@�1yX&�;M����:�S��`L��6@>N�T0��P9�2��O�	� �'
1O��r��u��-*�"��I��X��"O��#�*P�		����#>��(��'~"=aL��r�Yq��Y�v� ��)W0@�&�',b�'��aYD%�(Y.2�'����yg(
${���(�5{�������z��'�vP�EM׻C�џ�_(��']�+�qӣ8:C����"���3�#9�Ջ`�!�	.�E8�7O&��4뀇I�l�s0�X}Z ZG%�ش�?Y�C�?���,O��U�r�(��&ɯ&��4x�[=��!�O��%��0}�����Z(����t��Pkܴ|��v�'��6��O�˧��i���d����Y� y��WK���?�؄K�C�O����O��NȺs���?��O"К񊓟t��`m�U��x�cY>,��aH�	�:z�y�.Ek8�4�t�:3�@��5@��oP\�bC�B�!K�8lo�U��c�2B�x�LA�3��� �I<V:Ua���21�����b�F�k���p���$-	�9��<K�#ѱw��L����y���	;�n��(O j� �e���'N��Ә'�O^NH��L��Z�pB�W_����'��U��ʖk����ĕ�'dfL��'ȽJ�HKl���b�$!���'P�;�M�� ڜIUKNN��b�'����D�xς��T�MA�x��'��"&��S�ȝ��e��D�j���'̖�#�JZ����kvkR�5�@�'.v��sI��d�m�Ba�:@��8C�'��uj�b;��S��D����'\e�����
��iѨ�;��S�'�)q@/Z�K�6!�׈R4� 9�']l]��������f� %��<��'d�����üG�� 	E������3�';b���� 
)�)��^	����'��1:!)Z�x4�d�d�i�`�
�'� ����G��!�f�V���'�"��v��N���[��X�'�.�WLD��Q	
ARd����'#��eL�9����V�	9D��}�'�|M��NZ�\�Va ��܍>b	�'��`��F���$S�M'����'v��0�F�t�V�9n"j�t��'�P�Z!A@��=�W�Q:��Y��'�Ș��Ôn�h��M�5�"Y1�'�-Kc��(R�.X(�,�=&p�`
�'����{�p�'�J���	�'c082ՋԦk�J���cQ?�Q	�'�BD��Eʀ���
.b(��'vra8��A�$��ri�'���'������-C��a$�p�h98
�'L�;#����Ypf��vla��ռ7z�Oj�}�'ui�u��H��9�qL]54^zM�ȓd|p}�fE[�d��S��2E���ɵo^�E
�'<� ��S �����\;�	X	�_�l�5#�>	��I�8;��ED�1s��(2��Rn�<i�	��nE�����c��!oh��?(�mBU�2�'Gq��0# Ag?8
''ܚ�]��S�? �:�
cUN�	&F�P��$C��ͣW����=���O6��EΏ0$� �`o�wn���"Oƈ�d�Y�Z�	`�ǨA<�����O\�1w����>1ufUiJ���tbWHņ��7m@l��l�'�8u�s���o��!��lJD��'�X�t�4b
FX�t$�7jEnt�	�'���5�� #��JQ�@i��e@�'��ᇄO	 t�H`�dU<D��'w���A� �D�ˋ��2���'�6b��E >d�H*���.�v��'F8M��A׏(��d\��ht�	�'" 0�Ǚy��q�bo��[�rġ	�'�Hz���+O��8��@��X�<Y	�'���	�K'h��P�*��Z�ޅ(�'�v��4
M3)�V8�pė�N \��'�t�"���u��#�,9�y�'A�V�O�W
@Dk���)6>����'���x�J
!)��1�EH6i c�'i M���$_��H���^��\��'Di�U��b������1!j�m��'L�(adAHE�a)Tn��*|���'2� $F?Jׄ���B�f���'�� �e�&E�Q�E#�nX��'Fɢ��SU��H��I%��=�
�'d����%v�@`ÑD:s
�'�V �G&��GR܈z���(z���(
�'�20a���(PP�0ɳ��i{���	�'�b���H% 4�k�O�h�ʁ	�'1� �O� �����D�\����'�l4AkV
D�r%���X�Y$�A�
�'�� fh��t�~e�7.�$CX6AP
�'V���'m@�b���b��18G`ܠ	�'��Ij3@�����3�A�1�ĭ		�'@ě��Q��1�ƅȼ*�����''��PW/�3D2�MI�E��Ęi�'<�a����@��y���xmr=��'�  *Q)L9���u%��Gj� S�'�H1�p��p�$$�p�Y@���*�'ݺ9Jㆄ�r���
aDU	a�][�'�� �E�M�VZT��U�2�2	�'X��Qj�D�l��
A�IH&)�	�'ޤ<@����k�`H0��"@D�a�	�'���[i�8���W��9Z|��'�.X�q�H�zF,L��`�7DU�	�'9��A�ƍ!6ʥ��4[ �0��'Jb�r2�A�W���`ǃ[�R���'%R�9�nĩg4�a�IوB���'i���Pj�.p����Ǐ��}"�C�I�&�(�`���r�)��Ɣ�;	�8
`�br���矰۰>!��O"�a�ΉP��oQq�XR1�	9{x^d��$*��DV���`n� ����.�'"�!�$3m���vНP�ZTM��]�	�?�5���_�D#���ەo�"Ё���6?RFd"B'9\!�d^�z�0t,�;N�[��X�5��u ��B}���̺�����yb��J�$��7�OtҨh����x��N��m�AfԙS5H0�ag7r�c�,�lV�yՃ%�O��&�L?{�`���p���+��'n��k0B� ����>��+�;����3�E?�v�	�$_x�<	Q�� 	:UP3�S��P@1��t~"f�|?����bm)�#bs��T���S�!s
�q�'�Bp�<���}��`�Mߊ^z �����.Z����Q�Ԓ�H�
/fc>c�X�0kr�F0�qg��x���E9�x��kB�w����#bƍA�@��c��z)f�:g�(=*v�X�o�9�KQ4�H,���ּC�9���Z�z�I�b6��X�O� �̲wN�)�x5����+��EK0"O�q;Rd�#}�����$���`*@t~�ލ"� ���U�lԨ#��J�K%�xKŤM4pl��G�e�<y'2�2% ‗�#�@Z O�y 3 \�<a��� |Ҹc>c���Q �Y5�X�j�j����;����%@���B�Q�����A�^��` �>�:[�`���bc8 0�y�s���-��H��	���!�Q̚�?�dM��O�0����+zU��P
L�D��h"O\|Ӳ���X�lI�%I�E(>�s�"O�����9N��
�d�Ȁ"OyʴI�)Yp^��n�)R�9
3"O2T
�E�5��1�L��Y3�i�P��j�L��r\̙�B�8�0|�gF�#sR@����J~���,Eh�<IVhD�Dq0�`G��>t2Ĳ	]�E�K�']v��-��((:��O&M*A�3hP����Bɠbm.Y�u�'V�2��&��	۰���N��Ur ��c�>X0x�a�M�����(��y2r)�,�8��қ��'$�x@�ә�Mc)H/�������u�x]y���!bY��2�͆Qb��:@�D8f����rN$D��`�����횤�?2i�,������f�K�=ST��*�%�����H��(t�1AI%>��QD��߼ G��<\���.Ɂ
�BP��`h<1�k�������؞h�`����.6@�WハY��͈DޮA~���pk���ٯ;�"P��c��/d*�I42��FHJ�=��-����v"��DK�9���'<O�D#E�I=R�ѹE�ݒ�VT@���\\�"���?�^,jwa\7 ��]���Pr�.">a3$�a��d��g��^�\ ��aO`�Z�L �'a�<єR�=��p���]AX�D��/(*�[��
ZcT��d��;j��򆪂��a~"�]a
*�u��.2:0颇Y"��E�' :��ƨ�,�	p�M��JpB\����N̪�!V�i�`0TiC"F0h����C�̤ԡ��=� �{����	�Uφ(��̓5�7����Upl����9�0������	��<	�nE-O�^�JG7 ј���QPx��X�JF5$��ɺ:p"�:�I�!tL��@��:Kw�C#J�X�G˜�m�J��pO�d���9��dV�+< �K��,̴�X�a�$��'Ĥ�a�f~�)�(Y�h�� �)����s�-EW��cD@L'���C�f�$��Pp������dX��Ԕ����7Mn�s�k.k����'��)���8�)��q>���ٍ2�n-��wޱ�dƅ�p�up�ST���%9D�L[��G���f��m�$�#�k��Q���4h�?,�m��^D��6�����-Rz��'ɠ%3$	��H��@���x��'I�$1p�/`
� ��ګ>�����e�%]����*Bl���� �Y�q�?����LF�{�l�C%O�B|�u��	Y�����,
��O�C�"�A5�
/~�����x��!B9è��ɑH=��Bq�Ɇ3��(3��Lp4�OְSbK�B`h�9���N9�t����fi���ؽ�-��A0T��'y>����Oy����I�7Cb��p��S��?�c@�;
�y3 �^n�'�����T
�Ж	�XG��N2�!�Yo|
����M?5V��D��v��$�¯��.��dհ)�$(h�z����e�L9�p�c�ͯ2��h&��#,�S����|����!&Fe~d�`b.�K��ТF�{H<H�\?�5 �'�1o���@�ĞV�� ����'���<a�j�MK�Jg��*��x��hh<�eK��}��}[�#	/�! ��V�E��h��'@�C�D��Iז��U�	�&�jϓM߆���y���&�~�O3P:5���"�y"(*�X�� �_K�1��씩��[C�����doW�m��\:��$	��}Yu�	�y�ѓd�YC�#=V�-�lU�Z����'*�*dZDL���/ޠL��E�	�'�Fe`7.,{v$��Ȃ�,���$bUr�!���?&�d����*���hN��y���"1O"-� OK�)B�� !H�t(���"O�r�)�-���j��^�`��0�|2�_�h�Oq�,�&�0��]��L�
q�B�"O>���9�BbTkœtfF����͊U_0��DA'�h���)>\���!��Z&#��BF�
�,��eH�üEr�O�����3ye�����ɛ0�*I��"O� �2�$��E��4�w�+)���1"O�ɲ�g�>o�$3g�
��2�"OL]� e�bO�#��-h��L
�"OBI5ĽAZ�3!�Шa�&t�"O8�X� +&��t�0d�6w̜�I�"O���gYl�����ϜN����""O�ԡ��Τ!n�!�)O�!�"�6"O�i1+�	cp��E�K�kI�T)�"OlD+M�ll��gG6,r���"O����f�gR��^�8$B��V"O(��읮u+8�2BbX�r�"O�d[B(�-~�F�˶ �U�"!��"O���&�'k��y�a���:���w"OP���\�sen�����r�ʥhV"O�	��΄�"{��S�<:rF�c"OhURnx&P�*��xx��u"OL�de"&��6�W�/�����"O\���?�zL�#���kЀ�U"Or�����	r����+h�=`q"O�H��m��	&ݠ��J�$�� "O<(�Cţ\큡�ǸB9v�U"O6�A
��7�*m�Tj��Q)4�y�"Otha�}T꤀#(L�Pɀ"O$��P�^�+K�2�ȡ�FKZp�<�a��"6�����B)i^K7@�P�<Ydf Ti�D�!Q�	����J�<�t.�\<���(�\g���5OF~�<�"��S9��*����9fT��v�<��揟V�D!D�D�:���2#B�p�<���@<1��2E_8
�d��.j�<q���25�4�w�µO�vㆨ`�<y��1��	�2(�/9
����F�<����ic4�3�ǧV,Ա�Y�<����N�R�Q@Aj �z��p�<A��?h��"#!N�<���BB�o�<9b������sf�5u�J%��o�<A�d�-�T��"&.|�m�@#�i�<i�)��+	VM˰��9�ё�	�q�<���T�x���jN���`�l�<��
�-=�tur!��=(��A��<q��D\�0-���]�`I�s�<��Ɗ�.Gf���G�6+D��*
v�<�1��� �h�p�A�:ƾ!�"HMr�<���	(�u�rYl��(���X�<YG��-#�x���#�z���"�p�<�4�U�_,��8 ���8��Ee�<�s⇫c%ju!��@�ƸM���c�<aa��N�I��lX�W:>�`�Kb�<1�k�8ՐH��݆+��8yr�O_�<!b�3O��\�gNV��<���aC�<	rJ��	��i�g�
�xqJ�����f�<ɕ�_�H��R��T �i�<�%l��b��L2��D�&� pG-�i�<��Δ=M�@��K NbNa��"�h�<Y�Er��Do���1)c��e�<��6D�d�kE{o��U,h�<�2�Ҋ[?8p%��E� ����j�<i'���m}l��cOɊ%��5
n�<i�˝�7��\���TY��d�g�<Ym�$]P�d�7��2zD�#U���<���ʚi ���%��jK��B�hC�<����^��(@#kY�;Ĝ�ʢ��z�<����p{B�j6�����TM�|�<��`����S� �R�A�*B`�<�  �b�Mм?�>=q��;[C���b"O�Y�N��N���!�+<b� �"OP�Ч�Oz���C˃H}6A��"O�y�Jܖa���A��_��d"O��z�Ȗy�)��ڲ(�����"ON��#XwA��⑦��U��-�yR�ɖE�����`Dք��F���yR�
"jd呇.T�g��Lه�)�y�;��IÍ��b�3'��2�y%��1j�Y��Х]&��Q`��y����_���4��s#�=�����y���"1�a��ǔj{�Y��f�y�D�s���R@=cφ�jG���y�GP�-��5劈[6N\4���y�`�rOm3F�Wdl=�V���y2HF�-|-�׊��^��D�f�B�y�S6�����ݟC���a��y�� vۼ�P7n��9����e�̱�y��Q�z�K�E�(c}�d僗3�yrA����/D��ڬ)���yr(��^<� �Ѝ^�*�v�3�y�=hڐ=��˂��TP�l���yK�7�c������$j	,�y�@��^�^�7���`����e��y�*�S���S�F�i�b��㥑��y���7>�S�kקh�lL�-� �y��"�.�Igj��UF�}!g@��y���X���!3�ոD?d\r����y��a��`J��׏8K���R��y��61 rPk��@/�thZU
^�yB���F-2)����U�Y+"�I>�y�@V�yK��Zc�����yr�ߌZ0		S��;Tp��C^��y��� ��`z�Z�b�]�ф��ybc��&ݸ��D-#���Ѷ��y"I�>	:�P��L�� $����I��y��#
	�A���tf[Gf��y2�B>�D	6��HfԪ�'Ο�yr,.\H��"���("b��b�	���yҫA�F�d�W' �d0�(1��'�y"��v�Cg�WC��`�
��yb$: ���1��Lh��i��Ê�y��I�B��(ִ0~�#�I��yR,�;FX��e�Z�� �ũ"�y"GL�'�,h�!-�) ��"uK��yb��$8g�
hJ��#�'�y�c�Hf�����)1��c�?�y���8v
 ̉�.W''�6#҈[��yB��- ��bF_5vǼFq��j	�'J�r��I�L��
J7�|]��'|duK�+a*2�#�|�:tb�'~JySfEbˢ�8���p�=r�'m�h+qBΖU|�(80'ͱQkL%0�')�p�WFR�hyq�*J'J�u"�'B��pjׂp2�@
W 4\IA�'��)�2D�Iy��C�*���	�'��|r�H�#���`-��)^��	�'��͹t�0H Dk'/�+�$(�'9<���i���蘘�0��"O>q�q��#p���dg��y�͹5"O*h�F�?r<b1  <5��"O��፱]Hp�#e��0T2�"O��tjޗF��aqSD�i�|�`s"OP�FG�5hr�5�ѥ!Z���"O� ��j!'�`
"u���I��5"OָsƊ��_��L����5!X]kw"Oz�0t��\��<�'��W��a�"O�1)&�D\�����&l���"O��3SdȰ4�Z������"O��bfQ\2p�_��hME"O�M�)2����(�l Z�"OhnFOI��v������&�(D���7	Z�h���3�	F��yBd�'D�SW�@//��Q�ӡ�*1��T%'D�P�f COn1A�/���M�q��z�����d^
N.�q����D��8c�J�H�!�-���e��@z�8賩M�#!���'
�#��Fw�	�VZ�!�d�<29ny�Td��0��ZQGT�N�!�d�4yT�`1����ش���4/�!�ªt:��*�K��&����d�9$�!�I�*j��r�bC<%&�!ƈ��p�!�$L�m�苗&ߝx�P�gۛM!�d�E��)��� ���+L(!���wy$����ƚ�:(����6�'��F�iDqOq�RH���7d�y�.U6l`1b"Op��H�Ep|x��,�w��%����IܓQ��I���L��2����[u,�xSG�<?�����-D� ӷ�F���a����΀@��/}����p>�o�:l0\tsp�M:m�,�%�^U؞x�T�|r�_�OA�6m���A�*	��y��f� b0��e&	�ò��'fb�q���� PL�48`!S�Hr�P�3)�y��2�9	$GD�8�2����yL���@;� ތzK�i�R���y�ԃ���"N�	<Pa���yrɏ�j�\��G��$�p�劷�y���|�]P�W�(�8)J���y�D��s��[欖�n�8������'ў�Ԉ��W�kEB	sF߁f��!�F"O�#��]q�ԥA�DH�B�1�"Ox�A�fȨ#�p��7����5	��>D�DC B�Fd�A��-*rD� >D��4&�� �У�lp�C�;D�����ƓZ���R!�4jz&��B�'D�tѓ�K#k�=�%���2����!�$D��)`E�J��`;�FP�:b�!D�@p��O�`�n��$E*`5(	y�� ��xR�ҭk��A��J��Ïם�yҏ͛%FsQ�ߕ���%Y��y"�ցpQd��U{1l��B˴�y��J�1��'��6z��0�K� �y⦁)C�����,m�\�ڠ�ܟ�y�Q�n���h����ś�CB��y��
�lbt*r��<�|�x',F�O\���ߺ��t�0zph�'��!�$�9&�1�$�*�42�/Dy�!�$�'S:�D�qď0��Iv��G�!�HuW�}(����Y�P�C��V�!�ć\�`���a)� ��0R�!�ErR��b�̚0y�� $��(�!�Qi�0�M�C�2��W�O�i}!��7���1�摀+�T� A�G'L}!��b� H�AqUVŢ&��Q!�_��H`@g�z�n�6��
�!��p�jD[�( �T�Hq`v�^�G0!�^�m�0pӀ̀�wqLA�Ц�t!�$0\�H�$oP4'^�S��4 R!�� N� ��"��	�&֘<��!"OP�!@��$c`0�#f�a�tȢp"Oԅp��$9�$"�k�Z��`"O������x�n�Rg�-]�V���"O<�*W�_=j��xGNs+�[�"O\�0�E�7� g䏿Y�� �"O���H�'� u���7 e.-�%"O���3��O��yУ�&a��i�"Oz"�C�.zf���%�"O�5�S��K�Z�&A�t4�I4"OL�3�#��h�����cU;%����"O<H1-��@ԞC
���a	�"O��g ��q����n�����"O��[@郐7x°�@���~q(�"O&P+��F��(�J�G	fy�T"Ot�� -S����ޜ9���K�"O@�0�"-�<�rWL�	y�a�"O�ĳ�L<�*3k�E��Ԫ�"O�:���;���S�i�>�@�J�"Op�R�k��"D��"��#�ȼit"O�ܚWL��8�D��5@��U��}q�"OP@��`'2wv$�`�T/�Ta�"O�i��˘k>V�r���f*v(@ "O�\��"�!r�T��m̸M"�y�"O��@���7nk�5�6-�LB�S"Oz5`E]Z�{5�D�D����"O�j��O�8����,/j�Xp��"OZ����������<s�"OF�(ga]t�.��>*fʐd"O<|Z'm��e_.��&,�?c�K$"O4�ڡl�#_�e�W�TxJa3g"O�
f�Z+h��x8%���fq."�"O�Š�&9M���I3`�t�"OT\�O���������!"O�|��!��+2���"�zѪE"O�4�&R�z8�P�p���h�~���"O��A��%hvk'���f�8�
�"O:��D��9��<Aa"%Y+��Qa"O\�)�����Q��V΄��"O�Pe�4�|���l��yQ^݃@"Oj-[���9���i�[?Z�k�"O�!��H�VдG���v@��C"Ob���Er���)�^�-��ٙ�"O$M��R���Lڗ(�ҭA4"OP���HG�Q���P�Fo���"Oة�kĈj��=�4�˃��	�"O@�C`Η� �|�Ѫ����E"O���N)h�>]QFl�B"m�W"O.`� ��#c<�P´ ֙{	&�A�"O$���S%�����_/#�Ruy�"Oƨ!�Ȕ 7S(-ѓ]Ty��"O�9�ϗ�V�X� �m���P��%"Odp*�@I�p���Э�+}*YP�"OH��a�:?-\1Q��HQ���f"O��x��FGz����e���R"O0���ׯj6$�	����>!�L�"OJe�k:��(#��A��# "Oμ���JI���BL��Z��ԃ&"Oj4��۸Bt�3�	!C���"OZy!����~5�3�ٌm�r"O8�0�Y�-l(e�b�G3\r���"Oni� �?@*,��B��6g@r�"O@02���iup#�ѢWK0MS�"O�횔#��sr����I�5>4�"O� ڰ�@XT�0�aJ�i��87"O0�A���A��*D�-=���"O�-��mY�dU�8´/Փy�(�+�"O���%Ė]�X����,a�* 9S"OZ�@Bn�1��l@���UBX�S0"O�Y�  Q�fw��p��U4��"O0�
�Ð�uT�P0�,ƍN#|5p"OvUk���
	_�t�aˉ:g\H*�"OLX�p�����q��1j��1"On���@�|%r�it\ ZP��e"O⤙�MK��A���Z�0C��"OB���H#S��Q�c�}%=�q"O�T[��>�
d
�M���X�"O�ГQ�
iox	�� a��5�s"O����'.���z�j�7�pL�g"O�0�$�C�KFZ �� ��b"O�%᫔�7�.\z0K�r�x�Z�"O�Y��D�*�����o,����"O@Q�5�B7�T�O m��@v"O�q1��	x���Z@hďg ��"O�%u�2Dᩤ�����܁�"OPHQ'��	?`�t�wFJ�2h�lBr"O���$�ȭ<��r�R�F�DӶ"O��(D�X&U,�Q񆝌)6R}��"O0ma��D���ah��}.���"O�鹁��K��ӡ�5d��P"O�l9p���IA4�34���u��K�"On�SƋ�k����T$6�$Q��"O��p-��/�l����# ��<:�"O4�8���,XZn�(�\�Y3"OZ):�H,�ƭ�-�[��aAd"O� ����H�i��i�8��"O�� BF4?$�����l<� "O*���F���A3'��=i��ӳ"Or�iWdE�S\���TeE*J��+�"O0�1�㛋���X����b�L|3 "O�蚱���su����߲R�z��@"O�PVM�;2�l5!F�C,_��A�"ON Q��.}��2 ��R�� �"O��Q	�n������w�0`"O��&��:&�ӷBS)N�l �"O� cE���Dl�!��N�%��"O��7G �r)�e����ne"�	"OЌa�����r�
7`�:@"O�{�̃g����L�$2AC"O��ᡔ�6��A���lH��"OdT2�b�
##�A����$7�%Q�"O�8P�E7 �@�D!��,�ؘ��"O&�q� ПOư2�I��3�"O6D&�t����'H�=����"O��Yvۂ`��D3����~�V��#"Oؠ U&_�Y9�颰*�
�~���"O��0��*�P9�c�цz��rG"OH$�S�1?�ڔ�'B.N�T"O��8�ܘe�n9�Da�P���8�"O���Qb<yH�9��"ў����"O�Ɂ�I,9�UA ��3!5 ���"O �J'���e'�|zU��;l��˂"O�wn@>QL�q�pA��g����"O~H�%��!(���u`���T35"OޜkB�̀���:��P���ա!��Y2Vd
Pe-y�T�Y�"�c�!���D�J�c�A�J�6��S��+?�!�d�i�2���h�W���w G�"u!�� n|c�)Ä,K��гgL��"Oޱb6��	Z�x̹7'@.@��{`"Op�
��ͦ}-FI��ߊ�#"OL���{J�H��4h��0ڥ"O ���!=�:� �����2d"ON�!E�� ����4��&0��<��"O�!R�C�>٪l��H�l��  %"OV1C�ꅯT��� h8kB��A"O�@���RJMJWFA!(N(�+�"O,q"6	Ҍ<�	uE^�m?�d��"O��zB���*)v9��s�`�"O(�sK�p�"�Gi�/��,u"O��ض&΁J��Q3�-£\�$"OV�:�)t
p`׋� �@8E"O�ps�f�9
fHx�)��{O��"O8!q���88��p�Ё�.)�"O�!BԪ�*A�E�T�b�b�hf"O��5F�)vER#3	�,O�d�"OL@&�4gX܂�MЧQ�zL`�"O<� �枇0F�"�nO�C��۷"O<�:��C�[۞P0-ʼ$+�ŀ�"O<�؃&�)(�baa�,�$	��d�t"O�u@���j�8,U-��v��u[ "O�9�bBA�v�#���@�����"O�0kD�5?W.�d$˨9���"O�Ś�+V(\yP�H��*���yr &%2ܭ����:9�f=j�lL0�yr&ފV&��!m�,2zP,��+^�y�F��%�����#<,	K2n��yO�.\gRP#�V?;����6��5�y���.�2@���1. �X��y2H�`��ң"4*Q�Ř ͪ�y"i�nq����^�K4@Y��ڴ�y�g��u���Pc+[1I ����d�=�y"	=f��I�⣄2F���(N��y��@��ruS��W� F��"ħ��y�`Oɨ�Sw�~I�xp Y��y��#�
ĨTŀ1x�ؑ"���y��W'�}r�΁k�:K1����yB� �`��1��\�f/��W�ħ�y"ˆk�<�j7��d�p	٧o�*�y���0=b@
ŎZ0Z�X��A��y"�#p�1QRhQ�d��2W�T���xB&�29DՈT��\`j$�W�+kr!�aGh�+����s�j$�Zu!�Ě6�J���"�7<D��K��F�!�$� q����k�	 ThZ�`X�!�ɤ}Jٴ	G0)� ڧM�<�!�dL�x�Q��$�10 rx�DbX�-�!�N(~P����10:�IP ^�Bu!����
�Aveޒ^������v�'a|�ˌKu,�ӡg�:.��Ff�.�y�+�"F��lxd��52�,��j�yb��Z���6��2�
#���y�2t1�B�"l���ɢHЅ�y�C��AZ�a�W���Z���\��y�k�9A	�]�e��P0�*���yB%	z�9S _�
5��!V��y����yhZ!�A�����ȍ�y"�]"D���i�7rY�� ��y�)�����)ED3z�H!c	ط�y�
����/�� b���IP��y���$:�t��X�"��<A�F��䓑0>C��F�jy�ԡ�a� �Ȱ�=T�� ��B@5��xK����^#����"O���dj��Eh�=�e�# �91�"O&庀�C�f�xA�QJ��%��T"O����O��F�iY1JG1�L�V"O\Ո����̱A�h	+$��ӓ"O� vd��8\�hH�/�����'.�'����>��"�?�|=�ݚ�rQ*�#y�	A���OP����ИP:`���	5u�T,��'P�+u'�e@�� ��gh�'d�y;0E �?��y/�����'c���A�=>���Ūjyr�'�$$���\9i�$�*:v���' zM��e�Q;�E`$i	�b�'�L��T�ȗ#�҉�S�µ��M>9������O
�L�E�=zB�<@R��}!�8�	�'�j����::p�1���sʐ	�'E���CE�iv���.��d��d��'R*(�1�9��e�'@V11Мx2�'P��[�NΒ2A�4�	@�*��]��'�ZM���X/�$x�H%���	�'ܽ�ao�$[���M���08����O���>�B�Bũ\�`�� �&p�2����3D� ����	�~�P��1lQ���b&D�8���4i���F�p���A$D�ȩ��Տ�0t���N]��G� D��[$�&%�r��6�M���4D����I��.A��V<N<�P�1D���b'
+�~�:a#ׯVt���2D���3`��f* ��t�Ҫ"��3�+;D���A�S	U��IF��6J��@��5D���+�<����a�ݜH���H`H D��s���Y%���B`�y�$,ِ�>D�DSfA�N/�y3E� V<���%0D�@+f�@J��k"DèQ)9*C@:D��㡭��!32�0ӫ�%Cep�O�O|�d:�)�:�|l葤���"���D�>�"���'�u�A �Y��8��Y72�9R�'����#H�+@��Q �w���'!��á��<����'B�g|r���'�8���
켄���o�H��'�|���6���/��j���xߓʘ'(�P3�`�6�)��Kƴa�(I����?q�����"�����PSii�/�? �C�o�BE���^�� �)�!�D@�v���C� Ҹ������]�!�� v��d��'GcɌ�{�ʃ6�!�$�N�.��!f�*TW`�Isk�7D�!�DL����z�GG�j8�)Kªܔy�{2�'��	������	��NnT�i�L�\����O`���O�˓��D%�I:A&�e�t��5,u���!3-�B�	;U�`)��D�W�.11���l�B�I�f��'�>b~��:d�L	C��C�I�������:u�j�QŜ�b4bB�IP°tEV;D�0�`ږ��B�IDnLQl�� �&��_�
��D�<Y�'�|��#�s�[e�ZF�KK>����)X�^��u�`#��k��p���I�!�D���Ԝ9�&�&��ҷ�ʘ�!��<Y�Y�%�R�:Z$g*[�!�d	l疱�	���Y��ɝ.+7!�D��度H�"��`����R:!�Z&-h��1�X%m� �	�G�>d�ў���S�)6$s�g=�F�37��S��B�	'j����*C1C&A[�⊊y.�B�)� z�b劘4�h�h� �NRr,*B"O�����$�2ag��@;f	�'"O�k��%Co�q5f�_.�Is�"O��˧ޒ&l���Z)Lp�6"OaY���,2ҵr`��d��jB�.�S���xH�P@��?ڔB�Zf�!�DW�8U7ώ�p�� �!�[-3u5ɐ
�8
A�Ġ�9-!�wӬ�e���:�A��g�!��q�}�W���.��0$N�E�!�D��I��!�IȨ4���#�+�!�� ,�ej���:M������
Zўȅ�ӛTb �f�Ŭqz���V���Oj�O �}��@2l�rؙbU�b�*P!xɇȓA��!��%^_|�y1_�j�쭇� ,^�sGAϑ@i���$�ڕD�<�ȓzI���"o�>X�"mH�<D�ȓF-}����)J��UKr�QpNq�ȓ1�p-��ʭT�޵�� iB�ȓ����A+��B(.p��W�^����	hyB�|ʟ0b�0��bݹ@�&�)%1K��e���7D��@EŧU��h��hA�u=��e�+D�<G 
���HBO�*� ��2%*D�d@bY�5"��+W��8��E5D�D�����5��G�+I�6T8��4D��Z�BA��T	�A�P/ZL00A'�OD�	W�.����4nY`��74|r�O�����.�-�V �8������'9*�IX��(�0��v� ��6��3���X�|i#���2LOB�[��'ra��x��{�˘�y�!��<N3�d�a(�p�	H�!�$׼X�xؓ3�^�P�*�h�"s�!�d��YΒLI�,I�s�:���E ġ��%SH�O�7�(5BcҚw��T��	��2��O��X�<0TH��C�I�s�xXa�"��J��B磒z��C�	�m��$xnԻ`�n���� \LC�	���!J�DǙ-jV�����C䉪t���	��]^|  ��6�$B�I�?�E+jN�M]F�@D����C�ɥq�Vm��Ė�q��%���Y�t���7^D��U΀3 ��ÒA]�'�BB�I�f�l���H���	�"ɩ9��C�	1c���)t�:Y�p� L��C�ɓsKD�� �nt^!��3ϚC�ɳD9~ �'ȗ�Q�p*D�;w�rC�;�P��P�*�.�P-޲�l�1�S�O�F�S�R�X��a����f�¥!2"OZ��2)�,T����B�jX:�"O:����$;!�L2�'
�l�� ��"Ov��6�	�G��(�$�crh�3F"O飦��2,���%^5�Iq"O�<�v���>�8�Sbԙ �@u��"O�B���r�ś���te�Q�	Q>!
M4e�]� �N�h����q�<�����4]��KY!y0ei��@�=2��"OLp�a.=6P�����&� �&"Ole�]�4G�R���R!D,ч"O�lp%�H-(�t�H4e

J��"O�ܑg��-.�D�B:i�(��"OP����x��A$�>�J 2�"O�h���3v���V�4,�}J��|r�'�
�'J`��vb�0h�����ˮ""�����xL���^���`�a��+W����S�? ���Ǎ:���#@A�l}^I�"OjH�g��#a�xP�%(Q�-�XT�4"O(��w�8��1[��	nU�i�"O����D�!Ih�HH֠O��т"O���C��&~#�4ɡ/�nE����"O�bi�1Mq�ђeD�n�D "O D�T��>���D��0*a"O��{���^2,8q,O.~��I�"O���'�B�o�.4�"��4*�|QB"OHX	�k�8W �X�!�ޒ��ٻ�"O���4ˊ�sw����W�h�2p"O�Y�ao�w��VI(��.I�
B�=M����g���F1����(d4&C�	�_�F���"
8�8}��M�6f{C䉱��|�D�N(�L��1g�1��B�I,��ꉢJ&�B�e[�J�B�8��+�O��l�6���N�5�"C�0�����V�tS�G��l�C�Ʉ�d��0�K�R��W��]�B�I
`Ä@1gł�c�ҥ��hM�B��3U\:A�"�R� ��͇r�B�	23_z5aК�!���ƩM�B�	�>7��t �u2�-Q���F�$C�I�N���P!IҾK^����c$j�C䉮\H~,K�-T�_��A�)o�B�	�F�f��dE�j��h�rG]�w��C�	�R
�E�0��6�@Z�j�#��C��oMМ�@�S^�8�J�U��C�ɓm7��b�۴[ .1��	����C�		{]F��A�(�&�:���"qЀB�ɒ$ē��@ ܰ��G�F]�\B�I4?CFl�&E� �v��DkF'(�B��}hx�3�ڋ<'j����ś3��C�	�I6|h��8x6T8e�'b�BB�	�ELj�;��׊w�\��
�DW0B�	�}<�0t,��1K�i��`A9Hy�C�Ir"f%�`�Y�j����@x��C�,N�L�!��.Wӎ��e��B�Ɏ�����F���%kW�83C�	�k ����e���;�хn��B䉙,|l-�1G�?��ś�ЮIm.C䉲DU,��g�ۙ}��,�*��B��B�	av@��Έ��J��F�q�|B䉆q���*ƬÀz�.�����Q�C�:P����A��
���
'��^�C�	�Q�������
�eF��'HC�)$��	�W$�6?��樀�<C�I�t5�"w����"��D�!9�>C���|�GE]�+�Y#ĥ�2!VC�I0�\H��G�r��Dr�^#S��B�� [k6�AIY��H��ۗGݸB�$Z�^p!D��2@���3��]5��	�'��"���>�H�!��A�W3�D	�'4��b҈��:H���դ�� ��p�'Z�US���&0��R�*S�Kn���'d(%H�-K�bwR4�+C�Ɣ�Y�')�@r�[ =$B���*� �H��'� a)�R?��i�G@�,1���'y���鞽;U8E1���S����'ײyX����h4ps͎�Y&�c��$2�	or�7C%XL�9qS�ƫRt&�����<AD�)r�8R�ތt+�)��"M|�<a�/�<(��pC M�z���l
yy��'0Y�ы[4F
؍i���[�-���� P���M�>�e��2(�`%�#"O�aI�#S�-=��$��!T��P�U"O0�j�kJ[(4���gy�8�"Ob��,��\ٔJ�1l~��p@"O<)�צ
�N9�)��C�xq��_�H����4 ��������i�e�����O���0=�Ǭ=� 1cZ�X܈�b�M�<A�'�b4u�6���P1A"�E�<��%�8v�� G��d�L��jx�<)�%�f%����(w\��E�Kv�<1�&Z�p�����a't���@�Pzh<�v��}(Q��@[�X+��Xv�=�?�)O6����4ʘ� �F�wcp\V���'3a|rR�[n��������/��y�#��B��]9�OA� �1p#�y2%�� /��2�	�nx�y��d�7�y�k�+c��ҦǼc"���Ō��y�	GI��a�W�N�\P֣4�yJk���@Ϧ5�뢇_,���2�Oft� �H5�I��ENt9�!�!"O�R�f�yA� �dc�$b,;T"OdI�B��_��l bT�(Ʃ�&"O��@܊[ɸ���@�3U�b�3�"O�RB��:E�q�#��X�6q�"O`,3&�,8_J$�Ə�AЬ@q�"O*(P���.-> Tk�ώ,q�\TR���|�Im�ďI9~[<]�B��G�����+W�y�'�3��\����DiȀ�+�yY�THtA�"Kb�Ũd���y�o�W��ɚ4�Y/S�޸y��Z�y���
gH��e���L�0 Q�U0�yr�^/:;�)�Al0V�H��̶�y�K��`�P�x=$�|��ФI���'Fў���<ɠO�;*H�@ɝ�%���wJ�D�<9�%T�P�����5u����UA�<�F�˕x���ŨԆE+��c��|�<!��59��T���?��A�b&�r�<y7 ����C��}��PZq�	d���OO*�0T�O�M$�	��Ϳ\/B5S
�'V@8kU�^�L����R]�a�I>A���?a����O��P�Y0x��������*!D���"�<{[�ઁ#����:D��QU��-%��|:c$��F"�B�,D��3oDI���C�	j��њ�)D�TI4$ҹ0������̱1\Խ���%D�DĂ˳@�[��+�X�˧!#D�軀@�-%L���%�	>|�L��<9��hO1���Z��ªRɨ�c<��e<D�p��I]��0���˰= 	��;D�{ ��;�$�e�J'L��AP�'6D�|�"b�Ls� b�H
7gܢ]b��0D��CM݁V��h�d�/j~y�v�/D�$
� 2Ei1"D�r��5iԌ.���O>㟄�<�w�\5>����JŇ$�RQZ!��D�<A���D�QņT�MÒ�і�~�<��#�����mS5G��a	a�^x�<e��/iҥ���JN"݊c$w�<iQ�Cp���'x�>��r �<Iã�=oi�0������hk�П<���n���Q@�E�r�y�D�z�̄ȓ4�=*�A�,k��!%@.xX�ȓ�(���0]5rgE�%K\����x�1��Gܗ���⦐�Q��ȓ�]!�F]������̦|_ą�S�? (h�%�N�B'Bu�q�ՊZ��("�O�������`���y�1yw+D�X��ي2'��0E䋨~��`�I'D�xq�F^<GT� R�l�S���I%�&����T�AT��0s�0(2Wm�6if�2"O�`����kDD�d�8)���*�"Or�{ӄّD����V�J���R"O�\��nº<��y�ARCP�D"O���a��CB�( %d���'�!��	_���AI8,��Lȴ
�/\!�S:�	��ǌ�c`(ʥPџ�$�$�O�p�тG�|^����K�K3��	�'v�I�,\ 8��4+W�+z�	�'��-��Ί�4(���F��'`��'q��z���_-D��W"�(�'��x�D%��D�b�+t��,O����4� ��0�P�N����@0��<�	�<���ÉdbL�`&i�7���%�H{��^y��'5�O:�9��1�gKZ+L "��K#"J0�"O�x��)� i��	r�p:@"OJ|Rh8��Z ,��\�Vų�"O�񥞵I˦�10ꆗe��5P�"Or
b��V��(2ъ�ͪ!D���3��`����M7:�e�f�=D���&�]�I���D+�'&��3��<D�� "K�|4�`��9�Z8�)'�D*���'�[ÅY�@�X�	��6�c	�'RPD����c�f���Oɫ2[bXk�'H�p�T��	�c���+�Q��'_I D��"#���B���v���'�����AN ۬���㑬Q�	��'%�C�� F��C�-ޤ�
��'��i�҂�<=�����]4�[���)�4aI����|͂p��M����ȓ6��9B0�L=K������;����4�P�%�;��DҲ�Q�|ڂ���:tb,q�+WB z��ΘJ1������0�p�آ7�*,zA�U�<���H<�Ac�9�.��pɀ��x�[�l�i�<�W��%^r:��3�d��`C��hO�'�R%��:a��BpmQ4l���ȓj�ryӊP ^��J!�N�Oޤ�ȓcd�*���n��8���Uv(��#���(��Ԍ5���RU+��ȓCT�� BW�V=|�(� _Z.�H�ȓUʰ� d-
�8����M L!���F�8�@�]�MY�Oͳ2��0�?a��0|�򨗑|.ƀA�I0 ��Fx�<iqՆqRUȷ�M�t0�EZ�<Y�ۤ}J�s��{bB� 5�]�<��N=/-r0B��΄\s&Xc��\�<їHF)2�6db�&قJ?�4`l�m�<y0bD8ZD��'琪9/.�8V�A�<�U�H�0r�*� �T3�0��<��BC6��0*F�]�;`(�ð��P�<�J�5+��Sb�'��l��V�<!2`�:V��Y�hU	M����JS�<�D��0x�@������T���1��c�<�p� W�D%z��6 4}�$����T=�=+m�*p�|�@�&����7[ʭ�7��>&t�C
�rnŇ�%E\hC@/v���d}䔇�Q\d%P�����};���i��,�ȓ`�L�f�!R��I�byvm��S�? �=R����S�X<�^0��P����h��k�#$��
o�;@8��g�;D����P�c׬]K�a��T҆\(�,'D�<�.�*;}�E3G*�@���"#D���G�^.C j-���V����"D��*��K`��q��B@*���.D��h�� ��5��Ĝa�H C�+D�db�b�;[B8õ��DVe���<I���1A��ܨwI�ж\�_�&�Ԑ��o<���[�#jtX�e&+�,t	֥�o�<�F�E>ex��I��:���(5�Dm�<�ሿڈ8�FF�ul��D�JM�<16�@,�(Ыǉ�ܡXT�V_�<yg۵$4���F!�x�dm��C	A�<���ɸu:>\���QI��E�{x�(�'6Z�rb��h�2�;�aW� �J���'� Ph'��
4,�؃��t1�U��'Qh��Q[	-�
\����t����'���p``��jTC�(�f��'.(�rG�H��8�a�����:�'���Y�OǊT�D��(<5�3�'�v,#DMG{!)��vF�c�'V	�� �$	NE��oP�{{����'�0 F���*H����	ok��I�'�X�` T��vH(�'�`L�k�'Z6e��,{��L�M� Q�(p��'d�ibE)ׂK��6
�-N��@�'!��1"�h��MeI�E+��	�'Ì�7��
 �B�)�(�=�� �'*}z�n��}��ف�쌇 ���
�'�p�����5��/�#B����'VH�9P�ۓTs|��H����5Qϓ�O�����ŤuL���b�G�@YZ�P�"Ov�c&��]B�i�P�E�(T�"Oh)��3-���ZP��PH��+�"OiphB�m*i��\44��S"O��z�[�I@e�g�9Q�>0�A"O޴3v*��US���D^� ��\�"O�,�ш,X���%2���"O�d��[$$!����+ڀKij�"Op���*��),�",�F��!��e�
����]�<��bL�~!�ęf�F���
K�����Cq!�׋E�B�P���5 i�(���k7!���4[Ek�F	:Ă�1n��h/!��1A¨1&�PP�X��+�)4$!�DAS� �kek��`L��s��U�@!�$Vˤ�� �7��A"��B4!�Ę f�,ZՀU)K��d:�Eݕj%!��&� P9'ٮ[�����I��R�'���'@�)����O�n�����m_�1����5N̜{!��?"X�KR.��p0I-bq!�D	�;9L�Q�m�	t��e�ӻ|g!�$�$���-�*	R�Ұ�N�i�!�D��6�<��W!�43��y�F��b�!�$�5P��m���)��U�!�d&H�8b�N��U��ֺ�B�'v�|ʟqO�c��&�4��
�66��"O�r�ڛK��)���A3f%X�"O6i�ƈQ�kٚ�@�jA�u����D"O�-#2B��s�zE��j�P����0"O����M%E6L�p4cڱU���cT"O�a{2�%+��ܳC�:8���;R"OX�$M��Z�@��&���kи����O\��;��3� Px��jċN�	�ƭ5���j��d�O����P-���RQf[�##����  !���'&Gt� ��N�g�N�I࡙91Q!���n��k�UQҀ�!F�.=!򄔖_��� &΀�4x�)B Ɓp%!�D#y���J�c��g"�5;R�@xw!�dK#��ܹ���1���F��-�!�$�1�r��� :��4i���}��'�ў�>���j��O�fa�A�D�ze�v�7D��A�`nHD�g,I<xRI�2J)D�$`�F�(N]�"�̉Q����9D�衴mZ�f�KB$�m?��۴�6D����V�en�b�)4�b��v,4D�`Zrm�@&\!A�F���Rf2D�h�Q�t���Q�6o<���(.D�P+Wi�%T��*���|�Y&�.D����$*N\�b��=P��c /��9�S�'����L�B���d�BJ�-�ȓzeBEɊ�-A��M��L���c�*P �e��[��C�<��y�ȓz��u�����4~�GF!Rq����3fI���(�*�z"!+3�'� F{��d		����M\�W�L�p�a��y�@ȗk�y���:�z|�6�V��yB�4�
���1>��i�&n�-�y�h���߶4�v�c�'
�yR,ݸf��;��+B\�LBl� �yB�I@����,m��٣��yC�'�zY�v�}U>��d�۷��d<�S�O<6x��!3�����W=5t��
�'+�%YU�W��I�Nҕ%����'@D��1'�1�X��KȚNz,1�'4\��a�ШW�IS�UNd�E��'��x���	4�<Sr/�	u2��'�\�BG�1"��!n�YW���
��-���L
���B��ZQ�(#
�'f���K�/u�m�>h��q��'�(-cA��P���`ӀL&3+"��'�PM�Vg�.v��Z��L�;-��
�'��E+�'�0XBڔ[%*81���	�'T)r�K���'�/e��|�	�'�1u��-y��\hb�W��}Y��hO1�J�O�JY���y��(���&J�P��'�&@��"�O#u �,P+�<��ȓP�@U��G�1s��P��)^�����Ųs�ܿ,���0�>
��ȓu�))�$�<�h`��%1��ȓ|��B�
O�Mw(������>��ȓ?�hsj�����Q�-�2c���ן��?ͧ�O����΄�5�2��&I�����"O"@:C�5]��� k�.�'"OL���n�j5�L="� �2"Ob�8�
�2B�
3鄲Au����"O�PցT�c�L)sp'^�v��"O�	���M N����&F[H�t"OH��_�H��x�R���*U��Q�PF{ʟ��'^2%�ujF�[�F�NF.cj�$��.H: @�_~T���$5����#�I���b��u�&n�
3h؇ȓ!�l1s�[��)�@M�5Kj9�ȓ>���A��/r�(�%
2HGP|��1�q+W�3ͮ��o�YQ�}�ȓs3���F#J<O@U��*Ѵff��	k�����	6;\���+M^��a`��]|��B�)� �4�uH��%����`�u�b�����\F��ŧP��a�#�ư%���у�y�f%x6�i�Pjшڌ���`���y2��+a�\+R��e��;aJ���y哻<o��H���[��qkw���yBGB*g�TDr@�ø N��/Ǌ�y����/��P�AC�lBl"���y�,�1#�H�y棖"��`wF7��O��D�O`b>�ദ͔C)��+��+����"c:D��ce��%%�
��A\�!�~-1Ɓ"D�t���awh���]�:۾���3D�H�G㞝=5�� a$Q�<jƁ� &D��X���ӥ��';xZ}c��jXRx� Fx�k��I.������/=��R����y"�D)
t`�C �/�x��S��y�d״?p���,<�k�)���yr$�O;	�g� �fQ�N��y�ǺV��ɻ�0c_��f�@!�yҏ������(�A8DA��yr�_�w�ZԳEN=����D���䓗hOnc���T�Â� X��D8v>N����&D���3��Ti��8��	&��sc0D�ĘT'�o���u���P���2D� B!��.je��Bu��2����L-D� J�\�^�Αpa)W�I �R*,D�D#�س5�\l�Ħӌ�� Tg)D�p��c�1�l��CD��O��  ��2D�Р��_3M@p��Hb�P�k�g1D� p�j��!����҂�!E�<	�q�0D��H�f�
D�Y����ʲ�/D��xk_�XQb�3�y���.D��{AbƂD&��0�%����L-D�����Lh��D�0 ��&"��yD� D�p�BON�=���D��<:?T�`�o><O�#<)��6 �s���&H`|#�GPr�<�a��Z��	6�Ј�d�"��i�<A!ں7��mi�hW�Fm��GO^�<� �ܡG�h���f��qA$F~�<����p�e�X�H"�Ls�<!G�L
[=<l1u�R�H�ʼQ���c�<���M�8�ш�B��q���_�<���׍H�1&'H�[�Q�^p�<I�hK<&NP
rY�#��@A�h�<�㌖D&�P�󥁐c�`=ɴ.e�<���&����d��,�� �g�<� ۵"[���P�?(��R��[g�<A(y��:��I�@��*
�_�<�2Bb�bPۓLܑ/�L�Z!��]�<1b/�4�A�(��h�y���U�<7*�%���:F�_'o^�uKh�<��!������`�<� �D�c�<1t��X�^@ےdO�N�Aʄ��`�<�&��9nb��ee�(
u�@���Qx�<���Q�JS� ��!8�Z�ˉs�<�hD�2��G��(V�1���k�<�𬑰d���@b�((�g�i�<�; NI5���7b��T�i�<�ƨ_�����N�.�\�@sIEb�<����cNt�BC(-4��9�(Dx�<q1�. g�$2K�p�9a��i�<���
{�QGŗ��%i���c�<)� �;ˀ���\�A��x�A��D�<aw�ôx
��ȿ:"tI���j�<��C��D��C�/�2+���I���i�<� �A�T�����y��A �ih,��"O���eF��D��A���҂M|	��"O����o��EJ� ���ݺ1IV1pc"O��3��\4f*��1�ޢ^9,�P"O�	8�,�W$���4�@1��2�"O�ب��YЄqF�6*�k"OС)E M��x(�҅R<=%��	�"OB�h�O��F���bЄ7
����"O��P��3�:8ڇa�;um�%"O��B�ӌ)���JژS�Ȭ�C"Oz<�`S?�v��$�:g����"O�3�uZ��Ԉ� |�ܜJ�"O>�+�mU?B~1�!�
;S�� `"Oz��"9�੢�Y9"�.aQ"O�	CW4;z$+E<�2�$"O�K`i�PVP��i ����"OT�-T,Πhp���ck��"O�ę'�ة}�`��'֪&BR�"�"O�MH�%�#0`N��'��U4��"�"O�=��e�0b6��s0��Pn|k�"O\�3�H�,p��1���|���b"O� 	p�9!�U�A��n�1�#"O��q��:�`}�BH
G�Hm[�"O���r퐠|���%�C��r�T"O"�u+�.�J�����p(i"O�0"�h�@*e 7_��T�6"O��
P�}V�,Ke/L�9.�Р"O4$�eŧ0�CrMR*���"OF��1E�'Jv��Elڒ+�ځ��"O�q� ��� ��B�Ѣ"O:�&��3l����-�D�t��"OjIۗ�F2�ZYy��
r����"Ob@r-\���ѻ&C�3\o�`�"O�h7�Z�]�J�-��rr �"O�f�Y.2�,���z^� `!"O֬(�>n1�a����^:�X�#"O�ݘ!Q+�tx"�̠SV�:U"O��C@
��=����ba[3'��mZ�"O�A+fm�U���H5�	�-j6A��"Op�&aɝ0d4���4.�U�r"O�Ű�%غ>�".O�I��u(�"O���w��/�6 �Q�9w�
 ��*O`��3�W)@�0S��X�PZ:��
�'Tb)a� N�Fd0Y�HX)���
�'UJQз�ц�~�i�D�T�z��
�'�Y�0H1=S�i��+�K��L�
�'攴*#��r���('�N���
�'�9 �\.���W�Mn\XT�
�'�&�5�M� 8�) E�a�D�
�')^����\�I�@%Q$dL6R*~1�	�'P�ͲwU�����#.�;	�'#2��e�9.x�(�9���	�'�F�0�`K�M;F�ѱ!�n߮�X�'����B�5GuTb��O$gт�Z�' IcZ�#���dc�-9�'�"����T�D�6��(��c�i�'Y��z3 [�b��ŉt(E&��9	�'�hK48��AX�b ,(�ʨ��'���r����X�Ė&GZ���'+85HqdK�/�lJ��|4, �'��aQ"F�AshO�Y�T ��'i�5(�T(M5&�����h��	�'} H�#k��6cdXt�H�^
�q�'e� ��N(�F�ۃ$V
�!���� >i�`�\�l����#t�D"O�,R�N�Y�*%AEߺ""�HE"O�|Q� 5L"Ա0d��;Ȁ��"O윛1�/K$h��O]d����"Oz �tE����Pt΂-M��c�"Oq� ��W��A�t�Xw��aC"O�]9��u��B��3b"Hi�"O63 ]�2�Y�Q��<�~�
'"O6"��%gƼUp�C��je|0�E"O�Iۃ`�6��1�#>\y�� �"O��!p'S<
�����D��T)`"O�Y�Ch��~A["aҹ$���P3"O���Z>^r��!�4�|p�"Od�h��U�w5��r��}�+ع�y��\)]q��b�fԉ.:�A��U��ybL�73��,��Q��E�c�U#�y2�X�%�<��s蕂N�B�	�O0�yR�Ʃ9�I����Kx�q�+��yr���>M�du�A�@����`�A�y����E�5p�B_��d	ޢ�y��S�<�<�:���'1�И�ϙ�y��+P�.��$n��{,���Ğ�y�I"z�	���F����ND,�y�$Dv�Zg[F��i�tK̪�y��-�j1��W8>L��{As�<�G�l20��qi��3�D��k�<�5dL"� �RAڞ:��� �a�<�ć۝k���fi�����_�<�`눦6��r��_�~N�H#D��Y��71�lZf(Ӌ$�����4D����Q�s�d��?C9B���*O�QJwc �!�c� G;(�D� �"O���d�@��I3�̾{p1K�"O�I�a�0
>��sfG�(n:�"O&�� 晈;6��I�KL� n��C"OPѳ���<iiFYe�ϮvX�"O���C
�B\��)�i�~KR���"O��V.�4�&�[3�L+A�T*c"O`Up6��A!�\2��.F5�Zt"O2%`�cP)[d�4�G���C��t��"O��2�fڃh�r�2���"O�QKr�  \$tI�Yvp��"O��k�K�?�m���ށN��G"OFa��j�����K\	 b� �"O����n�;4�<q�D�[��Y�"O����,%F���h("���"O��mK�y��;�H�mP� �"O:�)u��A��]h��KY>��#"OLQpV�zF b�c�Y'����"O��ZĆN9g<ti�)�>���"O�!%@�d|��tǗ%p�F�jp"O��ӓ
S>�Ĩ{���OI0� �"OH	@2דW�(X�����$�D�"O�*���qf�����;$�JT"O��C͆4�z����B(
�P�v"O� ���F�jR�''޿5����"O|ȋ�i׹<��&,E.3���9�*O B7D��%x ��v>>l��'�,+��
�\�,1q�m��={�B�	�"έXU��7DP���FaİY�B�	-S�4���|al� ��5��B�Id2V�ӡ�"�D�jvME�)�B�I#8>^d��_3g����#N�ND�C�ɢ*�|�Xu����L���!�lB�)� ���Ў\��FT1�J�Kv���u"Ol5z�G�]8 �Ӣ�	z|�!P"O��J]#!��:��4d�`ˠ"O�]h�ȡw\, �C
�(XBd%�"O\���CK�o�Ƶ��#X�� I�3"Ox�s �ĒR��(ҁ�7�2��e"O�����<���Y'_�Ntl��""O�P�C/	�<��H�Q:jD��3A"O�) �hCP���)pU�4�f"OP��1e�F:��C�<B��K�"Oݠ1�Ȓy�^�J�h�� ��b"O���g� ,�\��նSB���"O��҅�͗(�"�I�&�a�b�c"O�@�c)����A��)$�uP"O*��!ω��Б�`�t8,q+D"O�HrB���4�*pz�U�M�)�"Op\q��(������%7@la�"OTu�#��<WH��A�&�C�"O�H�P��,"I(=�&�Gnm` �5\O<c��� F\ΔDH��)ls#t�����-M�Y8�h�'<E�=a�" �n ��	��ē)�tT�X7�L����22��+�"Oz����Xj��ʂ���D%*1�%"O�k©w���3$�����i�"O���Ř�(�s@_�n�PH�"O&a�Ƣʄ(��� R"�>I$)w"O��I�$[?&2�����.=J`�!]�L���{�dIy�,�;+$���$?@�B�IxI�D�$ܳ�B1r�n2��B��0�`Yz�K�P
ŚW΄;'���e����'p���>(��Y
�h�����'� a����-�,�sx�xCA�	T��y����"7'�2Y����I
�yb���\l5-�1�<�R�M�y���4^��``UVL�@��D�O��=�Omh1��ށ	�B��┑t�՘	�'(�0�OE6J�|!3��o���'�8j�J�Z��`�ҋ/m��	�'	�ݳn���r�g\.g�H��'��<bF��;;�yB,�����
�'�~hz��M9)����tL�<k���4�6�<E��4��X�q���ap��w�^6�b���V��Ṳ��tw�ɩ� 	�,�� �'w�~����'�ġP�D�*�� �ti1�yd��LlT�W��%3��S#m��yrf�%�P��O�
���ɓ�y��d'O2И�Ӣ5 ��c(�YHhY�U"O�삄J =\��jw��8��"O4!��폝'�t���?q)U"O��:�	� %�$MX�E��7"�p��"O�bq��Jh�-��O"b�1��8lOvIf$�1ی��R��0_�>�:�"Oq�7l]�r����(ԓ�l��"O�+ql�8b5��\�	k�lST"O�0X���� �ah�@�&n�Pg�$)�S�S�H��$�'�Y�u�L���d��-w�B��%7=D�ic$��|`VѩǢ̤V�$�<�˓;���aI�!k�����O�X~��mZr�����ɾJe�̻׉��L_t�M�*T!�B�I�i��'��:o�N9Q��'R������&�S�/&7��Y��M�t� &��c�^�?����đS��%.�0U��HdAS=U�OȢ=���+��F�F���9�,��;��:�P�@G{��Ʉ�n�}���\���੗)W�!!�� *�is�C 2v�a�C����H��"O&ݡ��1j��u����Q,����"O���'ݘ!㢝!��ĳ&~�0�"O��ą��&19��P�ep�ِ�'QqO��b7�#*{�I5�����I�� F��-~�<쓶�?2�̴Q`+Ă�y�˄�}Bh�; ��U�E(nN0�y�DM���}*��TS�B��m�:��d/�>ɕ(ȉ#PdH v�w�t��!Rmx���'6�Q#$m�5'x���ȗ|��
�'�n�9�̏���g�S<�-`�'���bN0N��V$���
AÓ�hO�Y��I?ߔ����L�N��P��"O�8%��	f!j�x�)Zm�J�t"OHI��� bJ��b.�,�x=�w�<)��3^z�<�jI�>�h�d�@X���O���6���*�O���0"�O���V0^�. �&���RDKe����x��I+G�R$�ǃ��rf��Pօ�
f�����?ړ3�"| d��X�*\��O�W�D8�O��=��Q�Y��Se]�wL���im�<@ѕ<�&��/2za��)XQ�<4i[���Ț����X�J֢�P�<�ǆ0&�<X6��9��%όF�<�4%֫_�
�Xm��\5�YK�Ɨf�<��Áx�:�$�خk�d�@�DDg�<	G��r��غ�o�d���h$C�d�<��MP�u�r	�e�"0��KS�Md�<E������9i[�|@�U!H�i�<�e$3d�pu���Y?܌�l�_��p=��l�"P,RW-��@�����P"m|!��-2ަ��@M�\f*M�7*ڿf>!�$�4��!!d�YO
��'G�u�ax��ɩRW$tIv�)/\�P�0Vc��E{J|Z�N]7
U�Q��Lt����g�<ɥ��q�!�����l�z�&a�<�g傆(�ĘB�Ol�p�S~��a8�X�0�����1��_F9xfl5D�)���J����!)�L�]�&D��C2*,F4��f�� �,"�M%D��s@�?��ئ��\���)��!D���B�Ȅ`�>���<����� ?D���A&��F��`3a[�L�D�(7-1�$=�O8e)v
�Y�T��I�A��@�b"OL(⧏D�t���i!Ņ�oG�rE"OͨG M�T�uX�L5���"O��Iӳ$f�Re��aD��"O���$��5�]���SF�ⓞ�����)�'P@|+��[,Xz��"�H�n�$`�IQ<��Z�J�{�v�Oq̓�yR��˽�����N���qP�ոj5����߰?QK�o������B�jQ����'�ў�'g,8lZSC��h���EA	Â	��z�r1�f(_ɀ��0�C� �]��aB2�b�_?t-Ճ^� (����Nܓ�2�s�	 <4�"�R�H54��ȓ,C�8�C]2p��!� M�wh� �>������Ĺ%���%���v1�e�T4�y2, �u0Z��e��2pt��'�Z��y"NM�b�)��n�c[�RP���yRo�!πAC�BQ�\2�=���۬��z���O�X�;�a\90צH1��?v�PA wI.�S��y��OR�(��o��o࠱� Pp�<��	]�^�̐;�Ȑ��oZ2�y
� @��Я�`7d��2�E�]��`�"Of
�
�v]��i��?�"���"O�t$��?�D��"�]�2p�t"O���EJT���e�B�<���"O�� �h��N�����/_2-�"O�i���,�N�@K�8�X3�"OJ�(�(��Ea�t�G͇8��B�"OV�P��E�a�H�`D�R��D@4�'B�$MYM��
���P
T=��GQ��	C}��� ܮ8�*	(k܅)d�
�"��#?����9�bq9Bh��z�n�JP矋D�!�DW�a�j���B|m��X���Ik��(��᳴�}�`i�7a�N�T<ɴ"O٫���$5`�̢7K�e&q�V�$4|O���qIS�z8�$M��1J�ٻ�O�\jf�֥����Ι+�\y�V+�q�<���	W��]�0��?I���@CBw�<1�HĘ=�µCY;4��d����q�<郩�2nO�q�G�m�:�C7̖Q�<�snHb!�G�F�I�f�L�<Q% 4<����%�\8e�^�p�f�]�� �<��B�#�l����� aωZ�<�
*q��5��D):}&��S�<�c �.O�B��i��;�Az���S�<)&���v���c&C�Y�V��M�<��d l��C��W�_k��j`q�<)d�FA��ɰ`�:,�"B �j�<�`iR�Y#b�[���q\z���Bg�<Qd�N�t��U�l��B���|�<��E�843vE8&HS�dx,(�@�|�<�#,\m��M�
=k�
Sb�<��͊6��Lx7�L���z���s�<���ܓ����h�6k�P�eK�e�<�W.V�0" /]�ءRTa�<�Ũ�:@$���,�$py��F_�<�,�%-�@�c�%ӥgth���_�<)"N����X�~�]�%�@c�<ɱ	�^ �h:G��,�������a�<�`o�{֤x4��e�a��_�<�&'�t~�u@`�sJ|�� ]�<i�ٕrv(���0O������V�<	q�J�4�����FF|�����[�<Qɯf�ze���Ϣ}��!OO^�<Q&�ӎ"�٨�Ϟ� 6�y��[�<qc5x���E w��E&WV�<���4&�AAԧ�Rf��$.�I�<���G�.fV���'�sB��Y� JC�<�B���J��	�F?\�03���@�<�V�Y*w-�q0�f�^)z]��IF�<��@*n# <q�%I9c�.����@�<!a�V7Bbl�t��7\{r��PGD~�<�����ؔD^�c�Ґ��"�r�<���.Y�Z@�$�A��h��Y�<�'A��v��t�R�������E~�<���Y#)���'��[�6d�ՀB`���� C.s������A�A��$U�/y�tEo�vD|,�%c0D��pTm
�%�!O 	�U�L;D�`!q��L��=��n�l���Շ4D���7M@�!㢼qc�7d��H�p�5D�h 3F�+\�%�Pʗ&@��t��a1D�(Y�nK�@�\���KI��m�6�,D��Y�A0F�B�G*`��m�b�!D��� .�]_�x�GG:R�����!D�����j�Z��@�ŦMg�M���"D�� <�%Ă&9��@S��PR�,T"Ol�'�ɂK_�p���f�X��"O@��f�.i�-u���t�[�"Ou�'��1zB7��>7-5ch<D�p�d�Z���P��F)x���4� D�X�w`ZJ�6�{��P�eh!���?D���I]�2Gb����<P�"g�?D��h�ň�G*��k��H�<)���=D�LrV
�;�j��3J�-~�8Y� �,D�h�6��G��x��ɉ
�5�tC+D��J�;�D i��ҿ7��H���,D������ �l��A�ʔ�DN-D�����E�@!�{���`9D�`�!��f���K(1KxT��4D� �7A>z�dx��:`:���*0D���ׁ���qr��@�PP�E��1D�`�L�
��d�/R�C�`�@#D�|aE�T6[U��y�cѨR�FoH_�<!�N�-�R�8�K��6�ȉ��_�<�p���	U�t�TMԩkI�qh�b�<�c��2lݾ-�E̓�os.i�b!FX�<AEڸC(b<R�٪]��ђ��O�<I�
@�b��\�%ګ%E$��E�<�%�ٯ����WbZ�r���KR`�h�<�	[n�<x�e��lT�i�0� k�<����I�fA�5��G�p��b�<Y'�J
Y|���RA���A�\�<!E쟒K���7R9�N�j��C[�<y�n�%Hm0@�Ζh�T��g�Q�<����SJ��p �N�n���*L�<aŇ;M���Vf��L~�u!�L�e�<����t���U�J�DMPSa�]�<�u�����'�J��z1��[|�<����I�De��0x���Bn�P�<���[�	�f�t�W�5b��S�<Q���7QVh3���$.�H,2ap�<��ƪ
K`�r�N'4�F�$�l�<�q�\>O7����TV�Ԭa6�Ak�<�ЅՎ
f ��̢lv΄�QO�f�<a� +>�P��L�X��H2�T�<y&�=8��rO/tA@�W�<�r�#Z[\ոf����-�UI[L�<���=t������;Р��L�q�<�v.C���Bd+Ĕo����g�F�<����1O���)J�Q2�A��F�<1�^��miA�R�r��q�`h�t�<��ˎ�F(��.��A@�����~�<)GBZp����=�^=���u�<c�
_E�ń�tХ;�%D�<�φ8wV������  �>����F�<�Ŭ˨J}��R����"i�ت }�<���&M����gE����b%�z�<𯈆D��rl��Z��*礝r�<�׎^#1cFT��K:;a��za+�i�<�CN���Bd�� Wm5��f�<��H�V��cA
ʊ{6�4l��<���U#	φ�@�(��i-d",z�<��H�:I�=��	4�pxA0!J}�<��k��CZ1#ӏ�dp^�#�$Xx�<���$wɰ���I�1e~�\�b��s�<ِ%ҁ$�R�b�造h�l�$-�@�<��I^�2U�܃�a��K�6ɂ��B�<��ˑ(�Jrf��lS�0��Ww�<Q���L��i!(H.F+8�3!�y����Q
O�H �T>O� ,		�/�|�����D<4[���"O��x����Z0�%�a�ϑV3J�2#�O�T6@�s���E��}z�E3�I(�%�;#ԡ�#�Q�<�2�ξt.��{૜�Jh ) ec�5-���s�b[���d����?�'R�1jdM�6j]Ju07�\�y�p9�'�"���ȕG)�y���MC���F�B�JĔt94%�2D��	(S�Q �>d���bZ�;d���Dſu|��q�[�=n�$�eO�WtI e���n=�ĨţgC:C�	�k�`�uÆ�z�f����
��Ob���L ������A7[3h|�偠.��3���'f4�Lpg�Y�<��錸zZ0�W+۴'��ƍ�?�ڸ{a��2{��Y�`"Q+h����O��A�O��9U��=Kk��1BOLT��L,x��q$��8a�� ��*S�ƠY���B�*�CV��ٰ<�#)�{�����:WK��U(ax��A Y�TL��%h":�F\	C��?3�b��T��eC����1�':T;�㊗[�*�s�Ȋ\z�њ�y��^���@÷U0�P���"��~ b��ܫq�~���C޺;0B�W�V�����,EA.%�rCګH�P`�*��f��2�#�?��!�gy"�U:���qw�L>E��aY3%�)�y�� z(��iB�a����"/�4��V�
}��"
��ٰ<1e�D�#J 0s��H�;��"��Cx��r/�P@�Au$I�6촥���K-���"��V?UF����B��D�E��w��̣���),�}�(��J�p����O��x�2@P�m���J�)J$Q�(%�˓[�>%)��3�dת��r⩃25pj�c�H�I���N����{��	E G��q̓�6a"��6���dw�'n�lHэ�C�S�R6��5M��:�1h�HI�}�t��'ptK�L��i��y"�!��X`�]�{�ҤF�O�rFqO��G�x�6�K
�rEn�9���9�h���A i�VI�f�Zh�B�	�:i�]��ʊ�L��h�b^��5^���<�u�^��<� �$�S�zǰ���"E!7�|��֬��R*z��Ai����ٻ���Ho�}�iB�}��	�u+��m�Z `���C�x���O?�Y��^0F�q�g��0`���gb�Y~�X!`ò5j�O�2I��G����9�����ǕdZ�@jV���D��?�p��G�2 Gay�/�$褐#f�h��QC-��2���Aq�Ί�?���N7�ȼK~n4i��)ǆ^30+�E8�Iٙo�Y(��hE�vL��c�~��؅a��(2��ܔ������ǣI0��4� ��U���)��O�S-���ˌ}T��S��-��"ж��)G IU@ �&����O����ƁM1i�☙4b�����q �o�����h� hl��ȱхW�.Hjp�� ��)�����eB�-�t]A���r⬐����>y�kJ�%޴C�������=ڧ34��r����`��Ƞ�C^o:%���h)C%ć���|���j�0�q��,'<{��D�Kޡ��t�H��P�ñk\��<���'+ܤp�	�4�li���լ^dar�G��9eC�v�����Z:S��<�����������a����L^�@�!�j\�<u�	N��8��	� ��S��Q-�΄Ӥ'̺)���K�,(ҨO���	L:Hqژ�h۾a����+qݑ:���	K)�J�(ɘ|z����)�r����-&��ҧ���a�D�GiպO���g�:�~2���Ť� )s�!0�Pa2|��IV�-���DK�@u�=�r��([�I$[�z�㬙U��8�CA��#e"��Z`��B��y1 `(�N�1R%
͓��N*�T�O����+�P1��4c�lk1�2V�\=��B�#?��܄�ɫ'3�e�#��/T�3Rl
�X�%�t�*{ر�0�D9&̶8�% R؞|��϶9��D��Ń�U��C@�%��x�#6S*�)���<qXt�Xwh��r��&�*@+��5c�h��'��"���"x�&I� aHf|�ҫO�s'�J�Kp�V�U� �[w��]�p�	ٮ5�\����k
�l����	�a}2�ö$)��o�=���)n���zSn�O� ����"�ژ�vH��5�Ju�t1��$��äi!�&sL"��P*V7x������Ybѱ�����u�h�j0)^	�f���^�)��Eak���``L&�O����f͏Ln���a�+��пi�Ԁ�!)qܓ|l��Ф��;[|��������7�MA+���k!��8	�!�D�%d�����
v紁�1�)Y�	�]t@���܌k�@���Rr?�����[���{�H6'�U3F�25������fm,8�U�'�����S�dW�S˃Yg�Y�\Np�J��Uf^5����ݪ9��`M���懬�, F{"(A6k?�  ��5dW�?�Ą��@�	@\�q(�_Bt1���m(�E;� c�d�@#�@�9mʥ�ȓ;���n�=�H �b���͇ȓ}�i�2`_"lP%Sǋ�"��a�ȓC��h ��IWR�qm����E�aR�ܢ/rm+$e��ni�c�d3d
r�S�'O�dx�2
�9'刵��'3b����J�J���[$4��fb�2'tԄ��{�Y�9mHc?O�KcZԩ��9�T1�DO��Bb%̡e����H��Wy.�3g�!]� �	�����E�D\� ���2P�^��	0��T9��|�Tz��	i�(�<q����/۱�yB+֑at:���۾Y�:�f����|��YhW�"�)�Ӥ)��48���x�,�ԯ�=M�L�>�b����H�Z9P6IvC�2�\v��;��5�	�9��A��L<)j�%K��Z�,��>��=;���<�4AZ-Fʖ㞢}���ìb�.L��؏a��x�r)J
?y6�:�'����F�.R��t�`�/�����O(q������=1A*L"lD@Ae+&��X
6 <�O$C�.LPa,�z���t]�a�� =��`S"Oȁ�"��$=;���
��A�T�Q�ɹ3[2����S�8���㖫D0Q�&�S4 $��B�	&>��I�:8}� ^`p��&D�k���Ӫu�tDb��wo�0���VB䉂H�ԔyDM@p!�T��)�%e�'�D����'>��A�΁�V��]�/��9�'U�LK�ح�P �!ȣF ��'W"��"*�<���Z)DR�'$|��F-Y4|���J� ,B��
�'M���iE 8UL��)�-����
�']�n�|@�pF���.���A
�'�@Uĕ��0\8E�@�	�'���f�
 Yֵ�'j��`̈́	�	�'�(���HѢ8��E��ɘ6gˊ��	�'�V��A��/m��}`@��+X���'�~aV(O�#���T�"&tL{
�'�R	�a��&x6��P�T�Od,�@	�'c�azcW�$ڌc$?g���'�%�bnZ2Q���!��УF%���'pl���&KDi����Z�M��-��'\��% �F�j����,1`j���'���h�ꅀM6���@�A21
�'�*���I\�zP��x`����'hh�	Ѷ&q��fO5m$��'Z��L���T7��~p���'g8���Z�k��H�N�I=|PK�'���q�VNi�� �\�K/���'!Y�˲XFI�u�+���0�'���2�g4<�����7R�����'���K���X�9��Vx��	�';�S�O��!��$��E��D�p��'\����%�HQAD�:iĽ��'4^�*�f�%��`�d@=��c�'�h�2fʓ<s@8ԃ&`B�*zb�0�'|�xx�m[�`�Fe&$@�}�
�'�J,"4	��T������zH�	�'�L�"�,&A�M��>��`	�'� y���S9,x�J �S*|�n�#	�'�4Y�.ۂ/[CG
� �jݸ�'��=�_�@��ܓՌ[)�T���'#b �1�L�����(}�X�+�'U���"��b�AH!H%p�ɻ	�'�J��C.��	�ZB̕7���'�u�d�(qR����
�?�jL���� P4Y���z� ��*�4�c"OX���Q|�@�q�gOF\�"O����'(4�P��
Dn���"O��Q��k' <蝥x(˖"O���0h�;A�rQcPjS�f"�q"Oh�M 0��4;qIü�f��"O�U!�FA�����x�(���"O�;�E������p�P<Ye"O�i.E1��"`��i��(�W)��yb(V�"�Q�p%��eG�P��*�y�#F>]O|�X$��k��daY�y"��o*�q�����q�	$�y�G�:����H\8�jЁF)���y���9S���@ @D��yˉ9=��Hj�A�u���h�� 
�yb,G}m�|����m�y+�j���y�DQ 	�:�+� ���@�2+�?�yR���+��9)e�Ɋ*�Ѳ��8�y���L@��$��_�������y"�� N>x,&�81�� �y� �R����&h*��r%�6�ybM��a�z�	�,���
�M�0�y���001��j �ɩ�Ht��^!�y�)�.L��7n���qvY�z!��� ��&hI�Dr1@���ڵ"OD �uDJ��n�rF��D9TX�"OfIA��G�n����@�9]B�5h�"Odi �%�_f�5���6I 9ht"O���S�	V�`���[9���"O�`�����l�z=���;4jjM��"O�D�q�� ����'�Q:���"O4���FصM{��V��Z
<�"O,�abHKs���`#fA3^D�9"O4����|
§�?}T�|:!"OX5붍��*� S��φ1��	�"O��a'L�V�8��wb�
#
��T"O��0�ٲj�����U�_ê�y""O��y����/����"��g���"O��.�in� ����2CNԣb"O��Ґ��c�H�Je(G� ��"O.�8���! ���*�g߀2�"лa"O���1��9{��i�R��jsL�x"O0�)Ba�w�l�X�+;hL��"O�В'��=w
A���!N�q"O|�yB U�Q�µ���ОJ�=�0"O(�{�ѓ�乢� K�0:�� �"O8Ȫ�.�01��ba@]�u=� R"O�4�۪,K�l ��Q�8<)�"O@���=xTD�R��W:,�h�"On�z��<h\^�iꁧ_�`�"O�� ��)2�@��>	�$kD"O�q����?_�����G�BZ!	"O��rU	,��@y6ӳw���Q�"O�}��b�+o<��oè>���	�"O4�z�BO�-L��ò��1(U*m��"O`%���%k&�fI	2�l���"O�HJ���l4�2aȃ��bIzR"O�TC��0yQ�z�
��-�t#�"Od��r�ћ~xd�G��*d� Y�$"Oָ*`'��vY@�E�m�
��"O�x d�\)��$�"����2"O��Y��AE���n�B��5h�"On���a�Q~z��5f�Z��<�q"OX�
 |*B�B��[�(�nq"O� 
�����a_Z�I'
I:O����"O�I'��Q�D(�tlF�{����"O�D8�j�*��
_ �qR�"OJ0�R*ܶr��H9���&	�J= v�'S
<��	��S��Γo� L 5�ز ��U���O����ȓ;�
���_�4/�ݢG����<�gٕ􆕒)@.�h��U�P	S�=G�aaI�,���"OTp
B�I�y� ��&�2��¨Ŧ#c�(��Ar?q��ė����	�(�"� � �?��s�)�5Y��B�ɄR�Z����w���k�n�T$q	���/e�h�)w�Y�4�a{�d�$g"p���`���B�ʋ��<a�c��f��<ʂK	 N2@ )ԪB�L��,2��Yq됷�yb"�A�~e��� y���S����!|�̻�#��)� )DIW� ]��ș��+��\���(`V�mӣ"O
ذuFG�48�@YV�D�(�6.�^kld�Cϕv4d1I�+��j��� *�xEI��84�U����S���Ɠ���4o>1�D�rD��:kʽ�u\E���C�
�(B~^���<,Oғo�VfU�3�;^v��A0�'WbA�C�U:]q���"8��x�oū?�<��Ff
!Ap@���	gH<�%(X�s2��V�HI'D�9'	R_̓I%L�w�\��U��g�o������!;H��d�Ň�m`7"O������N���D<��l����N���i!Ď�HCz����8�Q>˓?��$0v���� C�7R�R؆ȓL�.��u���v� �Ȏ,#9�	�'VR����	 ?����I�6�2}bT�4�
�{�O������d	*��hS��=�%s5B�AP�w�D�M�а��'"��Oǝ}Qf�7�T�YK`���������*�S?Ct4�0���d���1�̕�X(�B�IA��Z`cP)2��a¦a�95�����N�����ӵw���@�@D�I&
Bz�C��.70��ʴ8d5��P5��ix�BV�!��<�Ԥr��q��'X��a*U�HFx�d:-��KJ&(��ؒ?\0��	7]��-���)�!�@/hjX�Ɂ!"Vq9���x�ў0"�ۅFpR@�iD;$��
R+�v�-�P��Py-ߔS,{���u{�����?Ya%³q�pa�g.}��)�-�D��4fѪ}�	X�a��NB�	K¾hj��ˎ0ӄ�1q.�Q4*�7]|��欏�v����I&0�q���[�dy�c��Kr���)mL�Q�� p�T�
��?@|nA�%!ԸI��5$��Y%kJ�z�����X���,%ʓM�^�	�+�O�v� ��cCk�65���ϥA�Ʃ`��A�yb��j
e��J��-�&��w!]�a ǢV,�P�Tk�<E��{��2@�O>i�~:cV�#�:E�ȓ��)�d�
V�;��P�`b��%�0x��];�� ��	4S��|I6Ū�z�s'냝'8����-|��h�->-�C5e9z��4���V#����'`�q��H
`�ҹk�7J��d��gh�Y�F�H��ЁȖ�R3�:���aÕ�
�bU"On��bEX����F ��P���,S�<���_h�S��?�d�
��d��n�q� ��$�EE�<���D"02�[zZ���/L�2�f���+P��p=��N;��h4H�!8���I4�^}x��Y��=+ ��I��3���sPk�-m�DۇFC��yҍ�My2�x�M�-y���#ϔ��y��,�e�w@
��HSJ �y��N1\�RѲ�+�� rU;���y2o��{%IQ��ĉ#Y(�
���y2���m���Ƒ'��r6�A(�yb�ͪ��Ii�CN�*hF��y���!26����:�^���_��yҏ�7V�0���"<>�����yNA
E�p9[GE���X��Ѭ�y��fyj������������y
� x�:��UEBXS(��%f�A[C"O�i���0t����
7�9��"O,�9w��a~��1���7.��S"O����E�kA��02���hj���"OF�yC�O��@����i2 �b"O��)�$ӿ8�Lh��)Τ�v8)'"O�pQ��>P��-P���v� ]r�"O���5��{R���(�*�Г"O
iE��1��L=(n� ��"O��'c	"����E�(S�`"OZ� �ɥa�금�Z'8��aH�"O�!����8�p
׃R�G�B(��"O������<#צQA���x�|e! "O�ux�oߍ�.=�t
@�҅1�"O���ѦC>b2���I� ���+0"Od9��M�faSëQ3AvP�U"O�Y�7��M�P��ɗ!cHFفG"O�mz�IZ�hab��'H,���"O������?xP�;�$�~0X�V"Oh�+5��& ��=iƪ�;��!�"O�Q�L�&S�H ��pC�-"OP���1 8a�TM�DVqa'"O~����Œ�@!��˺2;^���"O*\!���(l�h��6D�]F~
r"Ox�'�3�ƌ�a�϶?$zDi�"OХ�!B��@$#���ΩH�"O�ЂvC���#f��2R��Ա�"O�z��K�g Ir���0���"OH�c� �$F�FE+�\<`�Px��"O ��&��'��dT T���ӣ"O"�K�#������C
�0x��)�"O����ō?!��z�L�v��iʰ"O� �)w��p2s�F���,��"O`,AtJ�s�fX�e�؎D���"O�Q��'���R�J`�q�"O����Ĕu�B����' ��xQ"O���eD�M��|r�$_W�S�"Oj|e�CT��L�0ZQ�83"OF!�R��ba�=���Ӛ=율�w"O01�a�Ϟ�Q���X�-�2�k�"O�-jpف/�����L��&AD 0!"O^�PE�(,j��Eʑ�qZ�cS"O�	���m ;���gJ�p"O�l�j��76�#�ǌ�^����"OƈQ�KG�8�Rw� z����D"O���͌=���)�Rh��"OjtY`푠Fb�i��<Mn�!�"O6�B���Ij�	C:R_��3u"O b���-���a�BXP�"O�h(����'` ���W3�x��"O�a8�D�N4�<����5N.��"O��0��
�/�0��-M�7
Rl;�"O��;����]�H�갫ʿI�ԌA�"OHH��D��=@y�ə�`��9q�"O��#2�$H^i���#ZZ����"O�l7K̝L�3�DTF���A"O��3&a�4�&I��$��9����5"O%ۖ(��kF:�7�Y՘��"OPU�t���d!�,ϔC����"OV�G¨x&�z뎶k�`PH�"OxTr�<x���z��Q<A~r��G"O:�e� �jlj�Ɗ�S�b$	G"OD����r�R(��dҎG��A�'&�y0�X�r��y�����o�~�E���)T��5 ��� j�P0�Q/*�t��E����k�"OPm�^�F�����ʰ�Qˑ"O*�ki�Eپ�ա�4ug"O�ze��0B:� �t�g0��"O�k'hU,�*H�e��O*�1 "OX�5̃�+bl�aB�A�p%�He"OH,���Wa۳O�4*vX��"O*;��D<_ |`֭Y/��E�"O�ضd�+\��c��Z���9��"O֭���ƈm*,�d��7�nt��"O�I�r�Y�-��H�#,�Ӫ,	1"OP����S^H�)C*C�G̲ ��"O@�D Aff�Z�������S�'5�Q-�2��ԃN�Ʊ���O>�����3]N9��y����c�=�Į�а)c���%(|%1� ����I�KQʧv������t.B�%�7N9\fX��hW!� 0Xa��y�@ƥ<�t!������ �EŊ�pP!D�|���S�D�$�dS�O��\+k�̫��Oy�3�"���= p�T1w|��˩O�� 5�A+����s�N>ݢ�.O,c�<�(!���6����c�e���u�ا$��[�ƴ<E��?i�B���L�aN��H$!�1j;P��FĈX�Fy��>%>O�ΞuC��г���6Ԍtb���1
��N(�S��Ms��ߤUO�m�����wG��s��S�<�AG�"���Pa]�jl5�D�<��� %3�hda�6hn(4����|�<a�� N�m:�K�6�D\�$JQv�<���%<8;��4�ș$er�<P��	^�r� C�UB�B�z��j�<�#�7Gu
�\�OB��r�L�g�<y KO�b��U1�K� X��Ȃ�d�<	G�~�ܸ@,_�} ���GCb�<�a/�z0R�6
��h"� �V�i�<i��i�tA;d��Rt�B�g�<�p �?:�J��%u��"�·I�<�����$R���<�� pS'C�<d�WlQ�q�%��&�т�F�<���2w��$+ch�	H��0U�n�<�&�"�,���I�0D���-�m�<�v �%7�e�DX�<�(�M�<y�36>�`��*��4��$��gT�<1/@�q��p�L
>��Z�
R�<��l"��P��
��0���O�<f�65r���3��X�d�<�`4m�D�iZ�7�nl�V`�Y�<Y��_;X�r�b�_�M����!z�<	FQ������C11&�3��t�<Q�H�Ft�,ц�� \���c��W�<�ĵxq(�k5�N#v��[r��T�<��� ��D	C�8v�����PM�<�蔋@ Bi�v��2��0��`�F�<�p��,�����eN�z�
�]�<�DnTO- <�Tg����%�n�<�1�%@T��u@ϟX�B�4D�t�<��dƥ(����jݗk6Iba�YG�<�/_5�LtٔFUV�Vh�u/�h�<q�JL�[�4��bgNw9*H�r�f�<��"�pPx�#��6|Z��f�<y�$`ɧG�	TdX#Fm��&GC�	�H���a��"|,��u�V�!h�B�N��i����7�H-X�BT`��B�	�Jڙ��)�>{z<*��\�b�B�	���y;��ώ���p�؆h2B�r�ȔC @�G������V�8C�I����5�@B��X`#/�C�&��Yy�ќ!���j�nZ�6B�)� ��A�+� ,�tz���*��e�2"O�= �j�*y/^1zSB��,�Iu"O$���$T��yGǪ7��iR1"O�lJE�8fY��E�A��x�"O*�S�h�0r���#�-ն\���2�"O�eYW����[�@�谹�"O���p҅j%�Ask��r"~=�"Op�4D�-Z�ri)#��)=��(q"O�e�b�6�4H�P��JW"O~t�p�J�`:�G[?)���7"O���%�[l�3 HT��n\#�"O�[օ<$0�p�#)�(w���F"O�{bNݤX�*] T�V"v�5a�"Oƭ���ˎ~h�Q!!��Ш�s�"O�у�'�@O��� ƌ�Q�p¡"O$�@ ��4�p�i�d�C'P���"O��䛥!�,�!D�f�,݁�"O.���A�C1VB�)6%��"O��҂C�37h���߬R5F4�6�4D�8��
W�=#Dmk�A=pr���4�4D�\��b�?lv�g��A��R�=D��8���)Y� ��- YVe�O;D�d�w�Y�ІP2��*`��Jg�%D�h!�(I�4d�C��J5j�sB9D��;�J��N!`�*0*�F�!�4D�$��-�0 q���"͆2U�X<2��2D��A�Ǌ�P�Ӧ�Ĝ9�U�2D�t
���I� ��;jZ©2D���ਆ�U�cW'_K��px�H1D�xK��1t�a���Z�g��d�U�-D���VG�#/+Y��(�f�t���',D�`��!"�X�o�o��3s�(D��!�Ԏg�	�i߆\��H��#D�*�j�:56x�9#��/G��!2� D����鈂S���:�J��>TP?D��0u�@�s���h�@�8J�4��n'D���P�2p�,�$�ɍ(�ihw	&D�\R"-^�9����,�/w��y��0D�<��BH68��5E��+l�6�,D��(��D8�����
[A�A`�$)D�|J�m�$TZԃ0�M`�h���*D�@!2H� tT��ҁo�3-
P�p��<D��C�ȅR�D��@�$�^��=D��Cf��>0`���oVI�,��ă9D���R�zH�ݘ�bV:,Z
H�$#D���#�P�5���I�f�yC"� D�� ��-�xYÒ�)V+����?D� ��.D2L>~0�	�t��lI��=D��$����)Ӕ%A��!��.D��@	a쐍�щ̙Ld��Ʌ/+D����bW�76���I^E~�9��)D�L��i�v�4j�3�B�3sl<D���pKI�[ $ݱ�(Zi� 0�Q�-D�L�bܳ�Px�B�`B�6�,D�[#��?\F��Y��ܣ@��i��/D���mӖH��I����qW���q";D�P��.AU�L���Q�g:r�ҳ#7D��@v#�z�f�"���!�@@�'4D��Pb��� 닚Ah�8�d=D�Pi1���1�j΀L~��@�5D�4bd�|��b'�f��V�(D�|�v��p(�K��@�~��x���$D�� U �h�0x��k������>D�,�œ�>�X��T�]�Z�:�k'D�� �4�FfW�Gb�q�P�6�~�"O���A%r" �Io�ȭ��"O@�@����Y����`IݷL�Fl��"O�x:���5V��xi�!�FP��0c"O��tB��{VcG�
?Q:��B�"O� U�X�I^Aڑ/���}[�"O��S�M�WR����m��
�If"O����b��R$��7�TG"OJ-r ��X���㨛�>I�C"O������'g�$H`j�:]�P ��"O�9�`��0��d� *��\"�"OF}{�`D�KF��B(ˊb��`9#"O�����V, �����l���ea�"Ot��taXiN���D�|��"O^��Q��6�:1�m��P��`�c"O��BvF007�$д��S���a*O�̰D��_(��A�ř��� �'�t�x�Fʛ��4#.E�NH!�
�'1�Q�%I�b3�/L*2�vT�	�';����3:�q#EL�5��!��'[���԰\�<�+�C�1�����'됴c�䛖?v��5D1q�hk
�'E�@'�CK�8��^2%>�{	�'����,
�REQ�,ϣ�LX+	�'%ҬSA���!�R�Bf����H�	�'�R����:CFe#V��LE��'�z5�u��3\*����I5���x�'\���M��)4�����4` ��'N<��K��K�Y E/�+_�͒�'	���WZ�H�d�^%Ge�@�']�6$/Z4�KWc׿�((��' ��H�J.!H���FH��>h��'4��m� ���~"�9�'��t�DC�{�&�p��D��j	�'ǀ5#�/��hph(��L-*���'`p���j�>����ޠ�0�*	�'����"Y %z3�ㆁ����'Sp����"E�8��0F\�x?*lK�']�m!���RT��w��#B��'5n|�d�2N� ��1�H��p�'��ũ�C�lX��Q
�k�'�Q�#� u,`A���(p Z5��'	
�!��G�$#��)�'��j���
�'Kr*��N�̘0�p>��y	�'��D`Ӏ�l0\���m�����'Ry
Ug�F�؛F���j��49
�'�B��%*��M�8��fZ�2� �	�'H����V�r��ȣ��^!+�.�8	�'W2В"Ǔ�X��@��(&xpɫ�'���8p�׀W�b; ω�����'����q�P����Ȓ�S<�		�' �U��A\+�1�7".Z!�5��'��a$̒I�b�����GQDu8�'8I�G�k�Je�d*[�T �Q"�'���0�ꋘ\E�l�S&�G;��!�'���S�	�/�1Y�
ӥD|xd��'.d���,ڮ/�I��g9Rܲ	�'�R���>L�� 3+Z7*)i	�'r�B�hUJЙb�ʏUz�Pp�'3l�`��	ht|���N�G��	�'��p1��D�!(�QJكE9�e��'
4�©�9"��,X�'��]��'�6P�H��
"��@��%����'�hp�ŲP��� ,�
������ P �b�A8�=���� O���@"O����W&�x���~B(H�"Of� f��hz@���凈9�ݛe"O�q!����`R�IQ�5'�I�4"OHـ�/@�vIͻ��L!)��)A"O�Eh0��=����%g��a��]�a"O���Z�F����%FT;�j�K�"O	��(0�ڴ�_���"O��j��mir�c�C͗����"O�xB�`""���50��A"O�M�Řb{�y�é#m�T�"O>�� Y,l�VA�6�[�s�$�"O.-�� �p="�"Ҩ߶[�^	�r"OJ`S��% ue\Ӧ}��"Ovi�	�a� qYE�Fˈ0�""O
E�P��ti{u��.s���d"O�)�"�G
LҌ<��$ٲd�z|��"O���u� ����s$[�3�mf"Ohi��.�54�j��B�.0��؃"O��V/U�i�Btb�K�B(0Xy"O�PE'�;E��`���85#rp(D"Ob4{QJ	9||�E�΀���p"O�1 ����؄L��B3v��`�"O(��F��H�J����$\���""OZ ����,�,<s�ш�2�Q�"O���"�=V��I6���f9"��"O�)��n�fv�R榘�.Y3"Or�b��@l&e����2��K!"O@�ҕ   ��     Z  �  �  A*  �5  �A  RM  �X  �d  p  s{  �  �  �  ��  *�  ��  ��  �  Q�  ��  ��  !�  e�  ��  d�  ��  m � > � n  �& - f3 9: �@ JG �Q L[ �a �j �s �z -� m� m�  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R��'��:�aɤ,��`vcء|�~Id�=D��Q��ˌE��z%O/Fs�mQ�7��)�S�'XM0�UhR: t�3��UU\`1�ȓ���q���*T <Ia�?c�ؠ��3�� �W���TCԺ����d7�-{G�0R�
Ը��̳c����N
��
����J��8�2qz�=��wYu���'R��r����e�4݅�u?��+Qœ�M@\
1�W�1�؅�h�eI�*�~UZD�����ą�T���Q�dD������(m��ȓ	��Rr+���<�Aj3\�Q��I�}Ru��4y�v��`E��2�b��ȓ2�,a양^�d� �N>Bņ�Q����$�Go 4� ��@>j�ȓZ�X��%G�,�Xd��غ"t�5��W# Ct`�A���X#��rg�-�ȓnV�yC�U���x6k�[K*��ȓQ^@d�p����sVl݁oVr���b2X�3SMD�=f8a!���t�ȓ0����I�<�XXC�
�Q;���ȓ�"��w��7+�dȘu�ȷ���ȓ;Ҧ ��B��IT��(��D�꽅ȓ9قu1�f�y_t ���7v��P�~- Q&�Y�F4���-wq�(��@֚,@�ϔ.���V�`'p܇�l;��GD8!�,�w-J*�هȓ5��S5!O�tk���f�<z6�ȓ~t�i1C�M)><)��EJM��{�R} �L�j
�*3ѢM%r�ȓ"��\��o_�4�WbD(l��@����<��;-o��P��&>�����C �3�^�A� ۤO��X���ts�*R)G 0�pHb:�H��?y
ӓA��Pq�*K<T��@e.�'�r5�ƓydI��C� uj���� �A���'7�	P!H�a�������far���'?(��]0:|��F��6��
�'"2���a܋,��aCN��
lL�	�'�҆�;V1�@&� |��TP�'0���"#�"�d��e���'xv%;	�'��$�߸s-V�!K�I�����'i�}�# )�j̓��_�@2< ��'��p`��
(两j��0=l��'Z��)�� �K��{S�L�@�u��'�J�#��D3.��i���ՋlG�
�'�x��&d�0:Ȗq�f&I�a�fԳ�'�\1Z�M���h #L�	a�9a
�'����'�<�,��#��I�*(h	�'�X��7gNa]r(Kr��F^���'-����;�t��*ԑ6Y0���'���t䖓e����FD�y��X�'È�r��4f�� Yu�
~�Hq��'�$3`�W��б�1b����C�<�AW�Zo�h�5˞1M�xS��z�<����6 x�y�� <�|���d~�<��"J w��@Z?&�HP뇦^z�<�0!%B/���� ��X�'��n�<�DD��c����-�{���1�E�<����;-i���g��n&�pT��H�<)f�<ؠ�h�s���sb\F�<!ң)]ݬ1A�m�$gn��P ��f�<� L0�i�3:���b1o��O��郢"O�A��M��]��8�-k�l�v"Ort��
D8g�\T��̜�f?���"O|��V$�9m���a��%
6�ɱ"O�Ī��$$���2���D�l��"O��)�ce<H=b$ٲ+�� �"O����Ο�t+���%�5}ò�ڗ"O��4��M��A�#J��t���(0"O����*ٗcJ��p��d���s"O
�5����6�h8Wo���"O��A�&Jt�H*�%�"j8	��"Of�->5���Th�hC""O��w/�p L��g�
M�$� "O>�`U��c����g̈7�v|x"OƜ�� :�)�k��E���"O$��0��<,��H=�� R""OX ���9^�H\h`Ȝ4��xIP"O���!�Y5�`��D	�6��V"Oй���X"	"m��AI���"OV��Z�SA�!�Bs��"OМ(�F�����*<���x�"OΩ�X�ޙ�4gW*���Id$PU�<�V�O�~�	�d(	�3Ѱ�Ɂ k�<vCʚQ��ݛyu�#Ak�i�<���<&�8a���yf!0���@�<yG�t���b
�S��U�<V�['g�Ȝ
 ��Z̐��FT�<�Rɝ<Gt$�#͈[Wꭢw�v�<��G%)�޽�5�ϊj��ⱍ	v�<y��0E����i�{��pZ��s�<Q�W {�j��B��y�>(aFU�<��Ɩ�5�"D!������ÊW�<YGF�y{��0���8�ɡ�i�<YU��%"
Й B<!db�hD�e�<���;1A��ӑ�ɸ�@ݓ�JI�<!��Z2q�@�D�$I���p�<���
�T'�ٓ�Î,B똙��N�i�<�	A�sP��Sũd4����y�<! �v����L'��5���O�<q����BB���j�v�"a�K�<��#À:�Z`��dݙR
RIȕH�<�e���#��8� ,��`q6��A�<Y"ݧS�i{v
�D.t�B�NA�<!2��>$R8�'Qx���
��W�<IB�֏}�j9�X?f���JB�Q�<��ȏ%ҭ���O�d,�Xc�r�<�e˔.ta�'��!HvZ	��S�<QP�_�K�B-�W!ٝcD�y��GL�<�7���v'ĝ�%�ΩGwRB�	Pd"Lq�J�H���k"�� :��D�[Ԝ�yP�8v�T��:x�!�$�'9]�a qHС84]㷯G�	�!��[��� �fK�56Ͳ���H�!�$�����P������p��܇r}!��50cX ��!�=;	��ZUM�g!�D�%!Z�u�����)ԭ��>�!�D� w#&4��ȯ�t��D��!�$��]���ȵF�? ��ٺE@S<!�d��Qj�%�E��(f� اF��X!��	O��C�A�]i��q�H�<�Wg"��u�ͅg:�T��g�o�<qGO�1�؃D
߷2�=���j�<�b�l�N�L4`B�Uç(�f�<��Ά�!�������8XN� mH�<� �s���Z|Ä�R?T���"Od�ڳhL�,n��֮	&V�&<pW"OX��@�3�����n�,T�Bw"O���w,K�]�P@Q�,жx�2�PG"O^�B��D�L}�,>����s�'���'��'�R�'���'���'��Y�̊b��D"a��?�@a#�'���'��'��'��'���'�F����)�� 	�!�3r,|��2�'�b�'"��'Dr�'���'&��'� x*4m�<$��B�i3�'���'4B�'t��'2��'���'=��I���B��q	�-����M)1�'1��'���'tB�'���'���'?r�
c�KX�<��k��:��M�'�'���'��'E��'���'���'����g�6m��@��եO�A[E�'��'`��'�"�'[��'��'I�0�� �w;T�S�+��I)���'b�'���'�B�'-��'#b�'�m� \<~=3�
;��c�'/�'U��'W��'���'���'!f��HU�1��}��c_:�~���'���'!B�'W��'���'���'�ˆFQ��Y��L@�8�n!�e�'W�'���'�"�'���'���'Y6���NL-+�V�z�ɑ���#��'���'���'+�'�"�'�b�'�\sD�&d�c�\�e�l��'+2�'���'7�'���|Ӕ���Oҹ��ܽ�6	iT�S]!b< ��Ky2�'h�)�3?Q�iTе���z��,�d,����,�C����d����?��<���}��i�
�b��\���یJ�4�����?9��Ѫ�M��O6�.��N?����\ ��Ȩ��͞3�p�+Ql<�ޟ��'4�>�-F0�l홗M�rXP٘��Z��M�&�m���Oc�7=�\�{��͝Z���O��8�2&��OX�d~��ԧ�O��D�T�i�󤙑D�D�y�,W��y����v���e��z�g)�=�'�?�A,îu@�,k�^%l�p�`����<Q/O��O\�mZ#7�(c�����	��[���z��h�n�����ݟ���<y�O��`0��$�Ȕ;��Mol�}Z�����	�J�z$���(�J����ߟ|9�
 OD��4@��Z�&�Wy_���)��<	d��Y�0|+F��=$��xpr��<��i��X��O�-m�}��|��kĿ�ޘ��-p� I��+��<����?���A2f���4��$>���'�hacG
�u# ���۠"�]�D�6��|�*O���H�.��Eu��YR+BT]*Mᄞ�48ڴ(u�q�<A��d��s�]�D��:L��(�K%A����?���yr�&zs�T
� �y� x ��R��$Z�BQ�������U&���?i�o*}�gy�� �&�Ƞb�1V��/�1+"\�\�'*�'S|6-V6c�Z�:���#�ڇg�D����6s^���U�?��<��?)��L;�b��Jr�=�Ƅ�)��y��_��M[�O��$�����)g�����h)<a�6��7�TP��i�D�IFyRQ�"~��n�?b�� w��" ,�	�S"f̓�ƣ����$�¦$������q����2�)�@��0�O�<�O��D�O��ΓL�66�9?a�� �G��~�P!�VǞ#R�訉@�Ox��4����?qTa��:��Ab�/�h<n|�WA��<�K>�u�i�ꀺ�y2_>ia���b�"MbC��\F~�D�"?1V�����|ϓ��O�� 	B	L,C�T,�f`E8I2�1��'@LPJ�M����4��������O����I!H$�q��;"�R\�5l�O��Of���O1������H�+�N���6�LT9դ�
i�`���'��keӜ⟠3�O�0mڣ!tz�x�N��Br �i5���,Z�Rڴ�?�iS�M��O^<��� ��H?)8&!_� U���q��2���bs�Ȗ'zb�'G��'/"�'��Ӏt�>$��ň&h8x֙��fґ�Md��?A��?YH~Z��Y���w[���gg�*N����2J��tM� ��|�,�l�w�)��]e��l��<yW�^�J۔$���ƇU�u����<��-�"mv��W7�䓂�4����
2�\a��d
�d�d�i'j�e�6���O:�$�O0˓l*��
���'���kx�i!�$K]QST@LS��O���'2h7F��q%��J��]�u�``QkP�L���1�h'?��DY |��*`��]�'d���D���?�!�&E*8"���$��9r���?���?Y��?�����O��RT�=Ft>��d-[�Abfh���OoځT�u��̟`�4���y�OFW�"�S������92EƠ�yB�b�V�n���y��㦍�'��(B���?q��ڿ`	h��f�*	[3х��e*�'\�i>���ϟ��IßH���}�$�r��u�$�j�N�j����'�7�
:n��O`�d+�I�O(�`�ǹ}�L!�@+�R��J�Q}b�i��mJ�)�&��Q�P?������K�H�%��`A'!9?�ta4;����D2����dX�dx��>6��\�4jZ�f��$�O���O �4��ʓ��F�
�� �p� t�E��z�̘ �I��yb�aӲ��O��m���M�d�i/��jfnș;�Z�A�8���vMWL����O���#�H?o1�����{�v�N�� ���AL�Fy`ek��תRdnH2O���O����O0�d�O��?icFkK�M�ѡe�,���{�\����	ޟ�P�4'V��'�?	��i(�'�0\c��>Zv$jU���x� Ȓfn#����	��|:���M�O�ax��Cb�\]�`*غd�֭��ǔzRt@�� �O ʓ�?����?���./�e��\��	2�G�6{�H�p��?i/Od�o��3Y������(���?=��5��T���@"Y6�T�bT�0|P�n��I�M�ӱi�lO�Ӊ.��E���n��x��'g�6��B�ؒ5p���&M�Gy�O]����2_�'10r'��;84`�̆.cՌTy��'aB�'�b���O��I��M��T�)*�]��ӗC1�8�R�RLPxP���?�ƳiW�O��'ئ6��;�t@{�� N_X5r��E�Q:ʱo���M[���M;�OjL��d�����<��e����LϺ}�|5�r���yBZ�\�	ߟ���L�	��P�Oז@�F��$|
h)2k��N���07)o�6Ԩ���O`���O��I�|��^w��wG�h��֙	D��@�9H�P�sd�Oh7��q�)�	��4�07mg��XW�[�rh�Ss@J�i�^t�v!q��*w�<7��G�	~y��'��
dڹ�p�*����p O.Aj��'���'T�ɚ�MctF��?���?I�B�TZ4 ���	�i� ��s���?AM>I�]����4
���3�$O�T���d�����X8V{�	w��cb��p�l�$?�C��'�l��I,,Q$Hi )H��3���RMX0�I��0�	�d��x�O�"�*e1��q�ǚ�-�
 #o��n"�y�Tx*���O��������J�i���4��+y�5j�f�\F�<`����L�I���ݴi��uڴ����./Z"���'��X�/>2,�wC�{���.9�D�<A��?���?����?a�.($R iB��xT�������Iڦ��/��h�	џ($?a�	�J6���� ��L��Pb��)�Pd��OH�l��Ms�x���h��gPAcdC�$���#q-(��<)1U� �	�H��J3�'Ђ %���'��L��l��F�\���iə��\��'�B�'�����t_����4d/���,.��z4��{Dy����w�V��k����d�h}RE|�^qo��M3��;[ϊ�e�ڿ�Q�X��9QR���-�'�bͲ�O�?q1r����wk*�1�)=C����gD����'�r�'/��'?�'Z��T!���7B5�Ű�*�f1ۖ��<i��͠�a��d�'� 6M#���s��p���r����.��M�=$���ݴ@���Ok���b�i��$@��)6\���h�fU�q���#�l�:Q�I�f/����?q��?���d�H#͒��2�S5W�1 Ql�O��$�<��iKFD:�'*"�'�哣>[�I��ªTQn�ze���	L����ş�m���S��)#F�F���	��w�bbƇ��x��Qj���7� ��_��:>�"O�o�I�B�|��򁀓B'�0����:H ��I����؟��)�My��v�l	�U���|, w�U�5=�a��J�N˓z����Tm}b�h���jM���,Ð��8N�1���ix�4g5��4���Ó��<��'4�˓Y��{0K�;I����@́\m 8ϓ���O
���Ov�d�OP���|��;6N<�R�F<�����-+��-/gC��'�����'��7=ﰤ1���4�����Tް}Ғ
�ڦ���4;f���O�~0���i�����F�z �ƸO&��rT��<��ĩq@����K�2�OP��?Y��V>xx��ѫ
2�x��'%������?	��?�(O�nZ=dD��ǟ��	�'�D%����bZ�yǊ��x�̸�?��_�$��4����=�$�2��0IQ �J�L�#A�m���9��zF
(�~�&?]Z��'�~���y�b� �g�����N�6R�la��؟<��런��^�O.Ҁ`2:�ڒ�M:�u�0�ιO��e��s��O"�KҦ��?ͻ5_�,a�GZS~�+%A��.��A�F��F�j�ZElZ�ƴ�o�A~�*��C"-��%*	Ô�\,n	�7Aí[
��AS�|�Q�P�I�L��ȟ|�	۟8X��'K����Y�^���H�VyR�iӠ����O��D�O�����C�p��MȲC�?�fy����=*��'�ұi�O�O��WC�!e`t)tJ�;^:�Q��Ί��|�RR��(�eI9'b�
Y�IUyr�[Ol�ԣ���8��a��+��'�R�'��OW�I4�M[2i��?��l	&y���ǋ�9?fq�R���<Y�i��O�M�'3v6mB�uQ�4h,u
��8u���a�A�:�(��re2�Ms�O�<bD
�
1N5�������c�ɀ19��#�EJ��E0�2O����O���Oj���O2�?�a�m��}6���Я�:X��az�kZy2�'�7*����M{M>�������J4i�y�*���J��>����M�Ӻ����T�P�����oԓ�`1���ͦ8���d�?�d�a�'5�h'�D�'�"�'M��'D	!���b��F�i��'�2^�4�ݴ��I-Oh���|�S��1��� Wi��~
����SM~�>���i0�6mh�i>�ӗ=O6�Kt�Z�麼qPI�$�8��sEC=/�d	X �Ky��O�<�I:n�'���1d�c�(��{b�q��'B�'xB���O)�	�M��fW�+��d:B>1Ș0�5,$$@�����?�Q�i��O� �'�N6͛�+`�A��]�FȒ���ҤnZ��MS"�@��M��'^`C�j�(���|��)� Rh``�2m��hs�+?:ī�7O�˓�?��?���?a����3X��� ���Yc��SaC�d�o�8{<t�Iޟ��I]��ޟ�j���˄��2z(N%x�`ݫ]l�T�L�F�eӎ9$�b>-�p�¦�͓�Q�G�Y�:w�͢R♱{����zԪS3'�O��M>Y+On���O$ z�d�8'/�5��
M�ZTr���O��D�O��$�<��iB�{��'3ﬀ��&׾/�j ����v^B�za�dkyb�':�6��O^� 蜁#��]�C�T��H�ol�H͓i��xTL�mTI��·�?���T=+�KZպ�p�'&��p��Z�x0ZQ2�ז?`<���'���'�r�'~�>��I2L@ʉ#7�,:VŹ�bV���	�	)�M�M�*�?9�N��f�4�m;�mP,S��c�_/�$�Z>O�n�MK'�i�p�Ȧ�i��˼ ���\�%C�m�w�RTc�L����{D���y�����>�]�<�	ß@����������Ic�c��Da���H{H����TyR�ӔBW:O��d�O����d�{ؙ0
@�+Y��r3��CŌ��'�J6M��$�b>�� �K�a��IJ�k�^8�cI;+v���6+����`녱*����&[κK4�>ɔ�<�'��Xx�51���r6.�^���'���'��O��I�M��`�<Ʌ�-$���tO�5hv�D����<���i��O�ė'sR�i��-ϙ,f2�2aհV�D48am��(��Y;��i�I�Z�����Og�'y"���8 㝱np�dd�9�ԡ>O����O��d�OJ���O6�?�G�T:zNR`9��0jt��)�-7?���F�a����¦&���@,�?JHL�cI�m��I�v	�j��M�Ľ���'V�v�v���� 	ߣ3�t��$N���|�*��W�>4J�2�'�T��'��6M�<ͧ�?���?��&�1@��)(���
s�x�D���?�������m�#�x� �����O�%�w�@|�J�f�/c4>�h�O�̖'�i�1O�S�g5�x��k�N6 �d�V	4���xf��@���*?	����@�'V�Ӽ+���()#El�@�F��V�W��?1��?���?�|�-O��n��j`�[B��qo@�;
_�U�n��(&?٥�i��O��'Ǜ�D�0U�m�%�Wt�q��;PI�6��O�d`4�xӆ�,��z����OXѪu�U�+���S����	Ν ��u�"��?���?��?I���)�Pܨ�qD\�Z�r�B��%t��m�"~���ΟX�Ij�s�(�������[�U5ڥ���эmb��C�B "J�i]1O�O�D���i��$�e�(X�pa
(0^�R��ܗ4���ƕ ����y�˓	V��W�����r�ԣ{�H��G�\iĈ$�՟��	���	ry��xӰ�`���|�I)P}t1�Mǭb�d�i��
1A�4��?��X�����%�8@��۸,Gd�7c���L�d=?�!j���i~�a~��ۆ�'HL=�ɨu98�+5�q��W2]>�hR$�O����O.�D�O�}�)��H*N�l�)�q`�?Q'2��@қFe܆��� ��?�;Wy��G�ъ{S��9��(3,-�`�v�j�X�D��U�z6�=?YK1>2<�iY(~!�0�&fS�����!P��/O�ImZ^y�O#�'H��'�R-�=��}�0��%�챐�OԚ+���5�M���<����oZe�s�D�§_�B~T'��D�.���������j�4��Ş&
V���ĕ;AqP�K��8(q��:k�Ph�'���x��D����`W�@B�4��U?q9� ���;'� 2F/ޛ*���d�O0�d�O��4�`ʓ'���(��l�R�ُ��%�"������Ѝ�+D����⟬��O�mZ�M¼i8:]a񆐐TJ�H:0��X�hEٿ>��F��pѳ��	N_�d���1��׾8��	�P�N�N���8Oz���O����O����O��?]��>� �ಯ��?� ͒EnNş��Iȟ4hڴMl^�ͧ�?��i�'{U� ��04j�	S��1EN�q(�1�Ǧ����|�5�Fβ"�%?��(�Zd�@�JXa��I�&�x�A�O,Q(H>Q-O��O�d�Oځ�Ĩ^$:2xT�CE��O>B�i�A�OX��<)��iJ�tk��'"b�''�2h4��uM�`����"'��3��|��i56M����M<�'�z�㝪@w�TP���jT���@�8?���t�ߔ^6��'u�����<2Q�|��P� �@��6Z�`�ゥG�"�'r�'x��T^�x��4z���sa�z�M��Ԙ>�q�u�S�?��-����G}�t�$|��Z��c�Z�k �p���J,'��.f�A��i�"�ܟP��&��h����+?Y3��:Rr����HY]Ŵ-)&�A�<	-Ov��O����O����O��' xl���D�r��A����X!��iG$�hp�'���'񟮸nz�킒�]:A��c�߄D����6�MK�i��O�I����逼+��6l�X
�f��,���!"� GX&��U%o���K�"j�dB�	\y�O�R�ڜl8��K��92�h��h��f52�'���'����M�'�U��?I���?iEi��9�ݑr�\�R!^���'0�o��6�m��U'�lq��5_�� B MƑ	��g�o����.ldP��]z�d��zB��O,���Ae���AJM�&��P��ղv�8�����?����?����h�����P)vT���*? NH�*4���d����S#Dɟ �I��M���w����-�'�^	 N�3E�h�@�'z���eӤ�l�pA��mZ�<�q3�(:W��X�� ��1�)��sA�EZp%�/���<�'�?���?!���?!e� ��0Zf@�n�vA���H����ͦ�K/��d��ϟ4'?a�ɱ��@R��ۺ7ۈ4CgO�(JIҨOV�mZ�M��x�O��T�O"�Bʇ1ʐ�2� β`y� =a8|8x�O�e!��D�?��b9�$�<y��$G�
���_�E�:\P$ ��?9��?����?�'����e�&�V˟!㮐S.L��)VY����џ�Y�4��'>L�L��Jgӆ�mZ��B�$jߜ!(&����E�m�f�faK٦�Γ�?��mΌ*����~~"�O�) c��d�5��mRx9�.�y��'9b�'���'�r�	�52�F0Xč�ZBgbߨ+q����OX��m��n>��I�MKK>QQK(T�$���W�����H2$�'�D7M¦e�-9��l��<��%��9�a�f�8�H%M�jE\	#�%����䓌�4���$�OD��P��T��Lε1U���$��Yw"�$�O�ʓ0�����Vb�'��R>A"�*9�x"b�H"�FI�ѩ(?Y�T�H�ٴaI��j.�?ŉ�"�Ձ�ֿ;y�dIԢ�ubU�g�o�l���O��?��/�d�#��S
Z�D+�%���-9.��O��d�O`��<y'�im6��LF	bFH���@�4l��j���>�r�'R�6�>����x�����S9�&�;���Z�,�H���eٴ=�����4���g��{������_̜ ��
4(�xdH�ʖ�bb"�Iay��'���'�b�'%BZ>���ȗ�Gr�+d�
������Q��MS	��?a���?9I~j�9���w��Pf�E��P���5e��i���a���nZ>��Ş&�plZش�yR��|sR9�T+P����yr'��J���OybQ�������'�FtY�M }�) �S����r�'���'�"]����4g�4Xx-O��DO!V�n	�b$[�6.�A3k�WA��X��On mZ��M��x���U۔,�~����(����Y�������E0
/1�����/�ʢw��,�`B£(�ĝ��)@�L%4���O��D�O��,�)�Sf�9�*��2b-	�}K�M��ly���U��OFn,O���՟T��I��֟�<s=&M��Ń<����Ǯ+�l���Mw�iO�7���F��6�{���ɟ`Dx���O7&���
_�P�Daz���?�,���z�Ay�Ogb�'b�'��A4b_�m�G�E5*�����e�.��	��M�$k���d�O���d�Ҡ�k��� 6 ��ч��;+�9�'d6�˦	ϓ�H�~�(�K"�:9�B��(�y��C�~(��`㝟��t��v�B�g�JylY>u�L8�cH��=iw�1��'�B�'��O��	$�M�`���<aS��k����5�W`�����A��<QĹi��O�E�'�±igH7͕�
�P���;��@���#��퉳t�F�	̟�p�ݠ8�T�=?���տCЏ;n����B�/���1C�<����?����?���?Y��4��� �	���E0d�%�C	A��'u2p�t s3����E���%�8���2\��!�"$x��	��'�����f�j�p�	%"p�7�s���"_�Y�j��>�j���l�:��i0�M�`����M�	By�O�2�'b$vD�8��(��j�a	��'`"U�(�޴_8�+OL���|2���N!fX��
�'���:7�[~�F�>9�i��6��H�)r �=IAF,�0���G���^�R�B�!��1?�'/���$����rj��'�n�,��Ռ�-y����?!��?��Ş���Φx���y�'�Īb�F�"'�lJ�{ț��DTq}BO{�h��(ݝ >�F@։0�&9 cJ榉�۴R7����4�����
?R�H�'����Gb��,�:=�|rA�?f0��Xy��'���'&��'��^>�:�.A�p#dܸ$%ʟ��a$fź�M+d���?����?I�'��9Olnz���H�8�����+��ł3��!�?q�4YZɧ�R���ش�y�#��.��zP ��X����u�P�y���#%�	�_�'&��Ɵ��I�)sDh����+T����w�Y��՟x�r�̟��'�6D�Y�Nʓ�?��I�:��Z��ל+P�*� Ķ�?�+O���By��'��� %��%����U�)1>�8�	̜h����OJ���#ʵ����f����j4����g�0�9�QaƦ���H�����������	̟�G�t�'�`���gX�G@IC��Iq2���%�'>�7��5.)���O��lO�Ӽ�R	Q3T��)�E��o7�Ik2���<A��ie�6�ͦ�������'�ht����?j�h�Dg`�k��5�҈`��'���h�Iꟼ��՟��I�OZ�OW�|��p
�b�p�')�7܈9*�D�O��$-�9Ox\����:X�d&	"i�/�F}��b�Rl���S�'0�����*K8t"��O�Z�ph��I����'��e�M�ޟda��|B]��b2��=ir�P��?QI�i��F�����Iߟ�����Shy�r�.81��O>I���·o!����[9�|�����OXHl�r��<�I��M�C�i�&7��:"�`�hfd�;�Z�q��?�@٥�c����� Z 쁬uL���(?a�'Կ�Q��[q��a��[$)�pz�*�<���?����?���?q��mJ-q��� m)>�jp�E/)���'�R�`�U�15�X��ۦ�&���`k��N$�3̚�+��E�����%V�^<��O��	"s�i���)�� Ԅy�YO|�����3:p"��I�?��d>�$�<����?����?���mKp��fI$�pl��?����J��%b���|y"�'��	d����ߝ6�N�rgJԮ4<��`���M�'�i}�O�ӹ5˨�bEN�P@��+�ݑI���[3�k��x���ny�OC��	��'�t,�@��*h���9�LN�|$l���'��'�R�O���4�MK���:[��P�@�]��ǌD�(�T|�+O�@m���]�I��MK���+��K �R?�b�W���t[�F�cӶ�i��yӖ�)��Sa��|�-O�m�ʺ`h�)Rb�fr�Yp�1O���?���?����?	�����gG���1�!(�zSe�I搨lZ$ �d-��ğ��	@�s������k�E���J�g>���KF�V�vjѵi�
6��D�)�Ӳk�XqlZ�<YqR�e��Q@���y�h|c�N��<i����dǷ�䓔��O ��ѽ%މ�`�k�X�k��M�`V&���OH���O��@��F�Y��'�rm)G *�s�VW�����_'-��O��'�(7FئU9N<فHP8*.�(��Wd���CJ~2��8w��@,2w�OR����2:ES�r�8L���.�����(~�'n��'nR�՟ 
��
�&h���S��@�P}�ST�P��4Ul�y�'�X6�;�i�q(�A&6��xU�ہO�>M�$s��z�4_����s�:pQv�uӀ���y��K��4�N
�%V� U`�+=D(L�Tg�#����4���$�O����O���֣E���
 b��/��:AE��8��˓C���%��yr�'�R���'&�q8p�I�Qz�\s�خ!*D02G�>�շiq�7E�)擘`ZB )A�^�ZX�a�BR����H�a��v�!�Q��O���M>a(O�U6L'0AT"� �D��!�O����O����O�<��i��5��'�4 "g/U5@�,�#��Hr�B�'�H7m2�ɿ��P˦�c�4{���R�$&��BV��(��#M���3�i���B�6���OJq���NL�j��a�)�
ˤJ Nݵ ���O����O����O���'��_"��+��"����H��I���Ɍ�M�2c]~�"d�t�O�9
%����!p1��|~I����c�	��M����D��Is�撟�sT/��l&�@biZ8m���Jw�_�9���^�M�4<�d�<ͧ�?i��?��^"�j`��Дh(E�T�P�?I��������:Dl�(��ǟ\�OFLŰ���6 c�B;V0�!��O�X�'��7��A(H<�O�J�kt�P��ÕI��a%m/S�J�b���	>`��O�	5�?��3�d](^��8�j\Ėc��Q  ����O��$�OH��<y5�i� ���\u��b�gRVʠ �G�y��'"<7� �ɝ�����}�G�Ǜ]�Dd84��kOjM8��'�M[��inR���i���]YD0��O[�\����.Ց[V�p򁠗�2_"H͓����O���Ot���O<���|򖠏7o��d#KT!bNz�"�i�)M;��E lFr�'(���d�'q*7=�<e��dd=\т�)C3��l+�������4U����O( B��i �;j=��42k�XQ���5���1�$��/�^�O���|j�HM�T�t��4LA8�a�
 3��i���?����?A*O��n�NW�<�Iӟ���w���F��U3�	�E��4�}�?Y�Q���޴��v8�C�D$�@�-�`�`9��N��I36}`%�A��*�b>E���'�t��'>%�<��8�N�fCJ$��(�	㟸�I���	w�O�Bg�1{S&�q�Y]�����1}!d�dm������ߴ���yG�˦8��$�ӇD�S��U�F�Q�~"�''�FN|�����{�x�q�PK�(�(���]�Yq�9�D�^�GSv�r'����4�����O��$�O��dO�18��c���8G�y�&ʙ�u7~ʓ=ћ�+	��y��'�����F�$�;#j�&B���tm��
z�ɩ�M#�i��O����Z�Ӆax�b掍����gc�6l4����.+�	�m�j���'RV�%�ԕ'�����:���e�7l84���'�2�'����^�<��4'
�T���Y`=��4hS�"{S|d̓+{���D�]}��n�,AmZ�M���^@�c�A?5}�`r�J�Z��X ش��$�� �������O�G�Y�Q�f0�0��� K%`����y�'U��':R�'�"�IKD
x�LL�<Υ��� |��$�O��D���YX�f5?��i�rQ�D
t �ZZ�!:�C��Y��Y��D�&��M����o�H��Hl�l6�e�����@S�lk!�.HrR�QU��?}�M0�<��'UZ�}y�O,�'���A��6��%��hO��(��'�RX�D��4B8�Γ�?)�����Kn JN�/Q�Ԅ� ��I	������4�����O�����C�+%8�s"b������A�K�v�Q��������H�8��pF�Ox�3���Nr��A!�7J)F�E�O���O��$�O1�l�|r�&��O�>��FC�~B�p$MC1��E��O<�mZt��%q���Mc�e�3V���c��*/��i��N:Y���j�
��d�r�|�	۟��B`�C�dd.?���ʧPl��'�ě.lHi��<9-O���O��D�O��$�O�ʧOV8p&'J�Uܢ����ݎ�Nڦ�i��C�'b�'���y�Ev���dopy�	�HS��qU�(#JX��I����I>���?}���N��n��<� �<����N�ܨh��q�!rp2O�H��Ȋ�?awa?�d�<�'�?	�?2j*Lh@�N!t�x�c!c��?���?�����֦ys�0?�������F'S<�,i��ݿ2����C�>�e�i^7��n�I"Z�����s1�!kEÌ�I�v�I� 1W&�4 ���>?9��1��Ĝ=�?9���%�� z!A��ް�4�V�?���?	��?���i�O�1Ov,���ƌ��Y��`xr��O��mZF��A��f�4�0��ě4O�,�����B���s�8O�Loګ�MCd�iG���i���Od���<��D�1%��qB��.�l�"u�^֖�O`��|
��?a���?��aܔ@�f�x<}�4�9�X�/O�(mZ�S�������D�s�DR��ťP�ó���U�ָj�����@ަIPݴRL�����O���aڍ<�.� '��#�*���Ξ(4c�!�����$�={i������O��{"H����Q�i{*-�m[(�DmY��?9��?!��|Z.OԌo�Y1��	3!$R����*4�B&H9D*~�ɮ�MS�⎷>��ie7��Цq˥�32fV"��-L���;��
$�$l�Y~��\�*�p��SZ�'��Ѿb���G�N�Y��u���<!���?9��?y���?���d�/IR���p�JQ���'�?�yR�'��g���iӑ���ڴ��1���
��.b�
�N^!�"�@�xl}�`eoz>��� ��!�'d⍊���1t�;�P 8b��ïJŎ����3m�'��i>�����\��Y2|:��VNu�DC��r4`���T�'�7�����O��d�|brG�Ԉ��
Nyxq��LD~Bʶ>q��i��6M�F�)rc�/�p��%DՂE���)2
Ϳ56l��P8B@��4B�៨2��| j�C�F5�VLC4/��#��',B�'���4Z� �ٴ݂]�墕�.8*��Å�iO2��L�U~�fӬ�PکO�%oj����i��d����i��'2�P�޴9=���vl�f����L�2d��$�~BB��!�Ľ���T�6�~,��Ǝ�<(O����O����O��$�O˧7l��Ȓ$I�4���9�h	�'+,mX�i�~��V��	Z�'&��w��Y��CR�,)�=b��R�>�Ν� H|�4@n�
��S��".AӦq�B(0���!��!�(aj���Po�R@��O�yL>Y(O���OB`��`�v�xC�Ŏ
D�4��O����Op�D�<�Ĳi��I��S����c�(�:�iY�r�l�h�hG:^�I�?�R��ڴ"���3OT�0�ldqn�;y��|zww�L�'������#�����ԁ\؟P��'W�A����2�@c�N����r��'r�'�2�'�>A��+3�T�Ц�Y�T�̌3%��`(����M+�n���d�ڦ��?ͻ���� C��]mXZ��@�0"]ϓl1���m�0n��R�vs��F�b�a�O�|���)B)�h� ��/O�0 �!�Q�ny�O���'���'i:㢒:'�\ <��ŀ��<1B�i���ؤ]�d��C�SƟ(g×�\�.��w	L���P"E�P���������4H����O��X�$���7$Rh�UH+5���굪�L��y�O�MC���?Q �$���<���_
q����;PgF�Z$�'�B�'Z"����Y�x��4wb�)��:���a�/��@I咥c��0������~}Fj�Έn��M3#���]��A���G6%'(�	�G�;���۴���Ԟ$Z����'��Oe�@�{	��ud�Z�8W��j"��	��������П��IB�'�X!�gA���mzF�Ö}�r ���?9�FV��a��$ �I�M[L>Q C�u�jd�3#S L�2� &-32�'x�7����
Ux�ns~� FN��̑�,))W��Is/��O@����ݟ��b�|�_���� �I��x:�莰��(C��X�.�Ґ�G�����ay�eӊ��f�O�D�O~�'n�8�P��K�D5����%�=i}V��'�p�|�ƣqӄx&��'!'����h��b.��%5�`8r��0@����Wk~�O*�(�	�VU�'︈����2�y�
S�&� 8���'�"�'�b���O���*�M2튚M�x���!#z�����w�����?�p�i��O��'���D0{� �X�N�L:��m#`H�7M����A�ɚ����'��Z����?����-�3 ,L�X@ɀ*5��h�<O�˓�?����?���?�����)ߩ��U���^0�s���xhzUn��K�,��ǟ�	|�SǟdZ�����΃�x;�L�� Q��c5���(�)g��9$�b>���^ߦ�̓�h僧	1~�(@�!m��9͓z����ӧ�O��N>�+O�	�OrUy�D�=$�.��u	�+t���O��d�O��Ġ<�T�i�P����'��'��\���Ң�2���퟊A�Dh���k}��r��`n���ēF����7%�92:�1��jm5�'vdjca����� ��$��'�8hASȝ�WB����@���̓�'�b�']��'��>��	���
Km�N��gC���=�ɳ�M���)�?m~�"�o�q�Ӽ�A,�1��	���,@!��#���<A��ia�7�Ȧq�����-�'�FP��&��?2��������ڊW�����m�=h��'��i>�����d������3B����V8W�nux��ۋ/]�ɔ'�87�U�!�X���O��D<���O>��� �&Mf4�����Hђ�M�y}��x�^�m+��S�'
�<8� �!OK�.��!/ɱ
�<�+W�T���	�c��P'�'#~m%��'*��27%w���&��e~�dy��'+��'�R��dW���ܴJ 8J�����@ΑmL�|`C$�N��&�$KB}�f��o�M3e�
�P���^�<�Xz�J6��iߴ��DI�Qp~UI�'��O�_�DH��Ķ8��ݸFJ�wl���?����?a��?Y����O�Fu�q�Ы�p/�
߲� Y������M�����|���6�|���xc�%�"�S8ym!�NADJ�O�$a��i.t�6�(?Ap�W�6-zl��FM�s"�8��G���B�O�1O>�+O�i�O���O�����Lh:-���HB�����O&���<9b�i��s�'���' 哉v|&��̈́�a�c���[)��O�����M3��i��O�S��.Ls��A%-�D��
Ԓ:p炜(���p'?�'7R ����jn�B���^���(��"y�@����?����?)�S�'��D
֦���A�
)��1����GW�xa G-vTf���ݟ�ܴ��'.�J�V�C20��r�(0N���iȧh�86-�զaj&J��m̓�?�a��J�8�ɖU~"G�QwHK�F�{��,ñ
���y2W�����`��ԟ�I���Oo:��FI�J�"�b�Љ2p���e�QE��O����OȒ����L��睾xIDiw˚�2*�[�,U�4P�����M#B�|�����'@�#�4�y��cn��qI?��˃Nۖ�yR�����	�<��'��	韴�	*?�l��f,:v6�rP��	>cn���ş��I���'S 7�����D�O����
%�lM��1b���邞,�����OlHn��M�x���`7:P���\0�#)���y"��5�J�	�� 	�I2?!�'��D���?�ֈS��:M�v)�fm���FG�?���?9��?�����O��Ia�9�fY�C-��xY��ҷ��O6yl�`��Ea�6�'ɧy�LX�U^�,��:s뀗"�|)�'5Z6m^ۦ�2�4A�v݊�4��d�D���'%	����w�U	ReO5K=`yB��0���<ͧ�?���?����?�6!�6&�.q �%Jp�$�%c���\ۦH@x�H�Iџ�&?�ɊP2F���c�a�hQC!�q���a�Oto���M[%�x��T+�}�*8�dV!d�|�� N:V�إ�B�����^�t��g͚�Ox˓X��Lqq��/�H}���I$�Ό����?����?!��|:(O&5oP�D�	^s�A�A�Zܹ`G�]?扽�Mc�2J�>�P�iqr7mH���B��$��Yyf�ƹvX �#/��3`&�m�i~R�)|����p�'��6�K8,+�!�G
�XH�a�C��<���?����?y���?A����F�\b��*�̢@�"N����O�oڒ3(�zd���|��M�Q<(z���7�����	�>H��O��oڿ�M�' ��#ڴ��d��v*
���Я�X(���_lD�ȕ��?ё�%��<ͧ�?)���?��hѮ�. !�
����p�ئ�?�����H馥ʄAw�\��͟�Ou����"�M��t�����,0��O
��'��i% �O�S�K�Ĵb�hTҞ�P�d06���m%i�X\C�M0?ͧ_Ӱ�D� ��+,�y@�η�-yԉh��+��?����?��S�'��d�ǦI{�A�8y�� � �H(�88J��<���~����A}�Mo�@Tx�6k0h�#�E�1�<��"�Ŧ�ش+<R	q�4��dXjjl��'��S�s`�l��Ê�S��->Lɜ'��	ş �	̟8�I˟��N�4̓�K��퉑1*�Ȉ�Q�X6mi]��O��:�9O�-mz��+GC9r�
��	&���Ѷ����M+b�i� O1��sr�s���	��N�8��_�F4I��]�[�z�I�-�)���'�!'�0���t�'���� ��LѤ��d��<2��'r��'	R]���ڴa�m��?��f]����]�&�����ͫ%�%*�"�>���i�B7-�F�I1+Ŏ�x	� ��� C���2������"�_�z!*��$?��'7���	�?	$C�y�I��bφT�V䚐`͎�?���?Y���?����O��!2gFDU*��HE����S��Ov�o�2A�6�M����4�.���޵#d�C�鏭}�&<O,Uo���Mr�i�ܐE�i��D�O��ze��Ҥ-,:v��!��Ztɠq&Bt�P�D�<�-O�	�O����OL�D�O�t(�/� ;Q��@b�p3��<Q@�i&���'X�'L��a5�y��'D�A�G)Ȇnl���2y��V��/Pt�jٴ	���Z���O*�t�ҶtY�`��*���89��Ɣ�r����Ӌ�%���)w�j���L�Z�$�<�-On��@��^@��!��,��X����O�$�O��U�"�H��<9ƾi ��w�vt�'�G�,���hʞY�a�'*6��O���|�GQ�4��4Ư�Ig�Ez�"��eQ<0�H�UQ�|�rh�
WX6�c�4�	�O��t�OĢ�b��l�v��! B<#�]u�܇y4xU��?i���?����?�����?�F矪#��5;%�@<(F`@�%^K~��'�6M1,��O|oE��[W�M.|�����!܈�aI>	�4d/�v�O~���q�i����Oʴ`.ԫt%��K��%��C��K+sS�
�3!R�O��|z���?1�O�а@w�|�L��3BT(��@���?I.O��oڳv�Z��'y��O���K��]�|��c�6h�m���R�yb�'Qz����n�z�$��S�?� t�2,Ә��X ���3�Ը AeG�ªLp���'��	�?��`�'@�E%��[�H��2Ң`X�����	������	ȟ`��֟b>ŕ'�26�ϼ"���
@	�E�d��C��!w݄��������4��'�z�Q���T���o/c\|��0��,>6-Pզ�#�f�u�'��@��M�?���\$����$P�T`�����<��0O$˓�?���?���?i����I�p���K�
��.-&��m�<hmMg^��ş��	T�ş�K����pn$-szp(�Kӄ7.�dΙ=��i�~�O�O�`�
��i���Z>tY@A)a���.���+����W�I��
!��O���?!�Hi})]�f	���M;��,���X�	��x��]y"Mt� ��6O��d�O�0���>E��%� p�(�`,�	����ڦ}��4{�'���G�_جq١H�<<�t}9�O�YC�C�8:it肢�iߟ|Q��'���y(�8#~!�1	@zV��86�'���'�2�'��>��I�ch�1
rN�S�>����ܕZ��e�ɲ�M����?�� ʛ��4�l���_X̚� ?F14��23O��l3�M�ҿi��ɪӽiq�I�~0b���OJxX�w]>"xĀkC
��$��2��E��Uy�O�b�'C��'�	D� z(�
�E1j���]�w��	1�MK��>�?I��?1L~B��t.��&I*wD��r�	9�JU��W���4[���`4���N�@[���U�mª�A���9=6@����V�	$8�z 2 �'�0�&��'��-��MH�l��+
��5^�t�I���i>m�'�6�S�V���d~���j@�l>ru�B̘=�����M�?�W[�d��4ab��b�R)D��5�L%
bI�"��Z)P3��6m4?���V�[K��/��߁��nǟ0lp%I�mB^F��r����֟��ԟ��I۟x��概�}@�L�A۶"��8DЦ�?���?i��i�:%�̟plZ@�	�7�5��G}���KtĊ�GU2��H<	��i7=�n9�%gv�(�T鋀��=2�<�1�*L��g �>���#�䓇�4����O6�ē�u�^c��Y�9p��"
��t��d�O��
䛖g(L���'mrU>�R��,n�L�s�!R�:}�g&?1"W���ߴcțF�;�?�"��/&:I���p{�Yp�FW�!����e�S�N����|�c��O�՛H>��9v�8 �A7���2�[��?����?���?�|R(O$�m��_c 18sgL�TW��J@%T��|��#�CyR�`Ӯ��J(O��$�1h�%S��B��d�'���f6 ��]k�`Pܦ��'�IQeg��?M����0`�7�1kPEڲI�\��3O*˓�?����?!���?����	�U�-�ըŮK|��`S��XHn�n!�	ßH��Z�s�8������k��tNR�fm�k9�I҃���Ҵiɮ�O�O���i��Ę)y>x� t��*��4 C�Մ%�d�h������5�\�O���|���a�vXq�� 3����CdX�)� ���?	���?�(O6(lZY���	ş4�Ɍ�,@�E�?���s�HO�|H���?�F_��K۴j~���1�M� ?���$v��!�R�F���9Hz��ڱ����c>}�1�'����ɫ6I��آ 
<D���Q@��`����	ߟ���؟��Iz�O��M]�#fnH�DOA=2jY(�bCx���`Әp0S��$:�4���y�jl�|�Gw}�X
Ã�y҄gӂ�l���M�Ä��M��O�L���Q����-�.~���E��p��J� �O���|���?!��?��ux��`1��'BM��k҆P-}B�J-O��mZ�Y�h��I럀��c��̚���2�Z}Y��K"���3�K�9���O�1�4���OOl!bv��!X3hT�2�߳ Rm)"�X.
3:I��O�:W$ձ�?1�O&���<A��ǧT�qP��ӣLD����W5�?����?9���?ͧ��d�ߦ��V������$yK��@�ᑆ�O"t�����Mۉ�I�>�Ǻii6mX���٥�\�[�rh9��ςF�	�H�����n]~b�SYktI�|�'��;��by&x
VbJ�J5H #Q�<)��?���?��?!���kQ�cZe���
���J �
)k���'F2/i��,zw=�>����'�C����mtB]H��Z(��������t���w��)�3j��7*?���"�,Kbk�^0R���h�i�2
�O>��O>�*O�	�O(���O��7�ʓ,�|�Hv�ιg"�� �c�O4��<�U�i+H���'���'��j_z%i0G�:*U!"a@�e�P�x�I��M�f�iMO�0TަL�3�M+�l�i1�
�*C%f�DT�h1qj/?ͧ>���d֞��"����C�E� -�%�2E�? �<7�'?�'Mr���O�I �M#U(S+/+���N�	�-#�!\b[�����?	b�i-�O(l�'�6�����i����n=�M���%.w�	oZ�M�'��M��O����@ޕ�"H?	�gMMɒr�W�-��O?u���<A��?��?���?�*��Q�g.p&u�6�%5]2`��զM)��A� �Iş &?%�	��Mϻ	�*��Ӄ��R�1�A��>n4�&�i�~6-g�)���eo�<Qs�� ^ �0c�
��M*h̔�<��3z���$������4���$S�'�$�X�'	x����ݕH�r�d�O����O�˓{��H7�y��'�"j����(�>~�Bezc#H&H��O�0�'?�6���1M<� @��^�ty*�OB�-j��@�����X��<y1!1�ӏX��!��B�D�d~���^_An-�W%N��x��Ɵ������F���'�� Bs��8yt��ᦝ�[x�8���'{l6�Z:�I$�M���w�̭���H�h�ԫ]L*fc�'�7�Cͦ�b�4wp�ڴ��$���J�'�$!{���3�2y�&Eѥ6|	rn2���<�'�?1��?���?�c�'*��q*�o
�P�����(�9��$�ubWmm���Iן�$?牟z*�8rNJ����sȗ�S8ڬ��OZ�lZ<�M�f�x�����@��N8�1��1^HV��P����JI�¨z��r�O��Y,F���`Z?F�r�8���z�,1��?����?���|*O�}o�"���I�7��z̱7`$@CSF�H�I;�M[���>I�i7m�ʦ����3O���+ާ� U!W�1?d��l�R~2�\[�t�����O��ʀ40���V*b���(��Γ�?����?)��?����O�䠈&R�;.LS�KI�Om�	��'e"�'��6�H����O�l�~�I�M�� ɓ/��+�i��\@*u�L<��i<t7=�J4ʤo��.���IS�ǱK+*�����+��eh�P69�l�$���䓻�4�f���O����t�f�A-Z9n��q��O�)�j�D�O6��V"�(E���'��W>��Q. @�����8T��Yp2f)?y�S��z�4*?�F 0�?�I$�
 (f`	�.�C��A����D.�}��©0����|: �O��H>��(�@%S�h��v�޼���S
�?q��?����?�|Z.O�m�*^����UǁWS���'�B(f�LP��>?��i��OZ��'�V7�
K |ܓbm��)Ӗ�1vɥ�>�lZ�MS&��e}���'2���m��?%���� ��L�v ���ؿC
`���4OV��?���?A���?9����d��UFT��!!T/Y;um��7*����� ��p�s�p�������}ˎ�)��4T�~*�-���i>�O�O2��F([��y��DK��٥LW5�t��Ë��y�aL
]�vu�	8?9�'��i>%�I*�����i�z"��t�7T�D��I�x����'�L7�θO���O���99��5�w&[�R���Y<�����$�V}�i�r0m��ēzt��Ќ55\��i�)�/{(�<�'m�,ړ�P,[�R@��$�P�|��'��2F(FND�]�.�`_R����'�b�'��W�"|r�\R��&��>4JhJ/�9��N �/@����IԦe�?ͻw ��0w)�5��)�(�&�X��?y�4w�����"=�h+�O�5��º���"ȫx�"��u�[=
gN���.�OB��|���?���?��*a���ۥZ���)�� 8���+O�}o#CJ��ݟ���m�s�@�r����,��^Z�e�@�L���O|7M�D�)�	��i��P��2֐�ЅkK`<zЙ�f���	�,�zT���'0'�@�'�<U�1d�>����˗��Z��'�'F��'�����TW� cܴ,�������aj�؜"̱���{m��K�zݛ��$t}b'g�n�mZ��MS��A#dB�b�	WkZHU�D�`k&!�~Ҫ��R�Smܧ׿c7�Dh@��ʴNث&RjT*1���<���?���?���?	��4k�0h#N�OґPs��1ck�b�"�'�|�L�R�?��ܴ��K8X�ru!^0���C��>�$���x�fs�\Dnz>!ÖI��crh�I8 ���B�:N��d��N�/�0��W�A3D*$�dL�����4�����Ox�DL�[d`q�ɍ?E�D�#�)���d�O��u��Ɓ�����O{�̺���96*�����>>Q8��O�`�'�:6m[Ѧ�HI<�O������K���V#6��(H&�O�(2K��P���4�d`B��^�h�O�t�Íe���wŃ=@L�kRO�o�7����������d	�
-
Mð@˟h����MS�2F�>���i�p���hCV�R�B\�/�Vx��dj��l�$`Ĵ�J"?Y7`K40�f������R�(�㉃�#h���S$R�$h��<	ߓ�p�Ip-�&z|*����@	��i�B�t�'���'/�@lz�����5|�Ѹ5n�8Q��ɻ�����M���i6hO1��P{si�-\���^ي &c�o����R�D_4�d0e3Ѱ�+�֒O ���K	01��q�� jx�y�P��;�ax�i���ђ'�O|��Oh5�a�O�D��Q�q�L�cMt����7�ɻ�����ݲ޴2��'�i�s��g¢9��_��e`�O�E3R��0��1�?�iʱ�?���Ofy9�/J�\o>��Ӧ	(��C$"O��CL��4���>#��LzR��O8�l��f�^1�	ԟ���4���y�
T���Xz��߫G4LzG���yr�n�R�o���M��OT�R�)�'0J<rwFZ�?	:���d�:����?$D�bgl��5�'"�	͟@�����	����ɨ(����)�+Tڈ�:��7w��'�47�6���Ol�D5�9O�`��ޜNēkR�p�8`�3�Au}"h~�&�lڅ��S�'hH@I�ل�D��d])m#�����_�y�'�F$�%�ߟ4�|BW�0r�i�w���g+Q(S�zu�0.埈��ğ��	ݟ�Ryҏr� ��3O��@qc�U�Dݓ�� �g�4��8O%nZh�m��ɡ�M�i�T6� ���`)֊r3|lcUD@�h��J�g��:�x�(痟*Ջ���i����Bd���_kt��(U��H56O��$�O����O����OF�?�s�H]�p��2���-R�b��3�k������4Il�q�'�7m>�$Z�~�X�CTC$=���@a�<3��%��	����7LhEң��X���� M�x�D�q�V���9m�6,P�'��4$�4���4�'���'��R��=�	�ֽz4� S�'�R�Aݴbb|�ϓ�?�����)��C`��d`�t؄𣜰F������T𦥫޴]㉧��Ws<t��lڗB���GB �p����U�f�y���!����y�-\��b�T�Q����"Dur8����`�	���)�Siy�nc��#!޶-���v�@28���ܺ+�	�Mˈ� �>!��i\dQC�k�5?t�(��������M���i~��٣�����D��AF�(�����"!� "ԠW8B���C�Ҥ~�0�cyB�'���'���'��[>-�À1rb�憎d�5�Q�ӓ�MsE'��<���?yH~�:��w���dGر W)+�O��$�@!��p�lo���S�'nV��
��<YQ���lz�a2H�^��I�b�<�W�V���������4�f��ٔpD���Xw����o%?�����O����OJ�@�6fE��yB�'��,�vk`]��o��o|���a� �[��O�)�'�d7�OȦݩJ<i��I���n�0�bhs��x~�Oݵa�Ua�%�טO*�u�ɵW�B�?;�L�N�?]^�� �]�X22�'��'v��Sٟ$I�H��BL�D� �J�3.�;�Sџ��ݴx�Ty���?�@�i��O�.R	�rY	�+Ĩ+B1�"�5�$�Ԧ;�4�?asAA$d�'��(P��W�?iPT�ȼR/᩵Lژ-P�9eK$��'�i>������	ޟ��I�#���C@Cy�4�&B-6��'-h7��)�ʓ�?	K~���[6��R$�^n�Ph�v�l�`��S��ߴ:C��=Op"}2%�¼D�:T2q�-u˴�@�B>j@p��t�v~���6|���Il'�'�剂A.U�ȚO�b�("%�[��I�I韈�	۟��i>1�'(�6m�A���֍&�Yؔ,�#J..xY��_	d8n�d�Ʀ��?qdQ���ڴ&��'X��P�� ������NC�0��yʕɗ�/.���O\œ�K͖����k��ǏN�k~����-�MX�p��du�P�Iߟl�����П���(]�iq�9tO�.X�1��!�%����O�l�u,���X��4��$�T����8�uJ��G�r�':�I��M�����N0>r0��O�H2���%q�J�J����LU&߿R��(�� ��O���|���?Q�wN(�6�-^b��%��J�%9��?�,O��m�)^�0�'n�R>�x�HF&P�L��KV�(�r��)?1`W�tX�4Lj��9O�b?�i�@��FذI^'$�h2Aɚf�6j�/��~��|����O6��L>Q�\G�؋)N���T��DP:�?!���?����?�|�+O�m6M�.%��J�'$p�$�p�<v��Bs���x�	��MӏR��>�жi)��wo�#yK
e �X��l���j���dϻ9^��@���[!d^A��ԓ~*��N�15fᲷ��2=� ��uf��<+O��D�O^���O����O>�'P;�M���&��'Ů	�����M��hI&��D�OF��t�d
���5Z�� f�=A|�KB���ѸݴgÛ�7O��S�'߸%*���<�@�Y2�bb��U4ҵ����<a`��?*�$X�����4�����3J���C`�� b�c��P(_�����OR�$�O^�p^���� k�	��H1�Fњ_q	p�B��$��Y�T��T��!���*�Mְi��$�>���R�x��L�2��0/T�2!�Jp~�e�aN���cXƘOz��IF�/��e)�1��n�_.x;3d��?���'���'��S����j=�D��EJ�3+bBUNݟ�@ڴb�n,�')*6$�i�)�c��<>����b�C�8E��,n����4���p�8�e&�K����C�:��C�O��UzU.�1����J�f���e�	]y�O-"�'(�'�Dˁm��+��/zl��X���1u�:�M#p%��<���?yM~Γn�4�j�)<}�")1C�D��At[�h8ܴb2�&�;���9��0��n�2R5�-�`L�o�<_$�4�e��ܘ�y��˔V�Wy���@th�G�I ������ѹ?���'A��'��O/�	&�M˗���<A��5N^���C��Q��0����<6�ix�O*y�'�X7-����ٴA����J�f���(T�L��p�0!PM�'�h��' H�?��}J��}��i���+���Ъ˝`̎͓�?����?����?q����O�B�uGH��a䀍2
� �O����צ����(?qd�iJ�'T(���B�Y�8 C��'@vp4`%�$J֦����|:�m�#C$�'Tx����sk���M՚W!�H��ȏ7u�Y�	2z��'t�i>��	��I�<�$��� ݩ@�&��pHI\3��������'7m�"e��˓�?*�DY�3 '+�d�R'ׅraP��4���ٯO�m���M3�'�����ƈP$��Qb��(^�0�H@��\)�!l�i>ur��'
�H&�4X7�ӵ&�ƨHS�	�O��Zc��Ɵ�Iϟ��	��b>ɗ'I�7�&9¶T�s�Y+�l��#Ϭr���y2,�O������?��Z��i�t�? ��6)��@%R��E10'�S�JΦ��ɲ?��(F-?y��	�M�n�	)�d@��!�И����"��
�y_�0�	��H����|����x�O�������?k�@��5X̤�U��M{T$�����O�������̦�]�Y���Ig��AeBEb$�;z|���4r�F3O�S�'?@FPV���<Q'f��\=�2��M�$}�o��<��O�5��D׷����4�z����LP��;��4��a�1��\����OP���Oh�pɛ��ڹs�R�'G"��2W��i��:�����"'�>�G�is�7�Lr�	"!�>8��IV�H�1s͂5	���c�T%�F�
zj� N~���Ot�H�H�e;��	�LZ*Q��Mp9�����?Q��?���h�&���*���@ş6r��I��G��$�D�yj������ɒ�Ms��w��Y�7 �'�����;�^:�'��6���u��4
t��Ϛl~��;�V �S�X��h�X�x|�3CO�5�h,�&�|rS�������	ٟ�	ğzd��

��9�p,� !Ӥ@9�Lry��d�4��2e�O����O����$�9U|�Hd���i\ؙ���UJh��'�@7�ɦ�J<�|"զ�%�, [�H���Ъ�oU!%�ȑs�.C���d�Q���k����O��-$h��Hֻ7���tE&�<���?!���?���|"/O�mZT�e�	.?ft���-D8�!ËR0#/��	��M���<1��Mӕ�i��Hy�)��&gx�te�@�����嗺O� I �O�]g)����d%�i���!R�Ȥ�А����k�f���7O����O����OB�d�OH�?ii���<��HI�vi�p!��Vy2�'��7��%3l��O��lZg�5� �R��5&a΀BjD"Z���͓�� Ѧ����|B�M�xM¨�'rր�oD9s�M���Z(���K�$�N��ɞ��'��i>A�I��T��,;�I�N�9�:l� ����I�l�'<6M�*�˓�?q*������^6�:�AA\�������8�O��l��M�'���
���#�2k�		s樻B�A	w����ˇ�%��i>U��'c�)'��M_�fy����gٴH���$�I�����ҟb>Ֆ'��6�K�]�pPK�̝#���Y���.l!x\ޱ�$�OF�m�N�{n��r����Ɔ��w�`4)����M���Vy:e�A_~��a��u�H�)���(r�D�%���Ҡ�ݾ���<����?a��?I���?-��aJ
;>����jG���ȕʦɐ�DAGy��'��O�Ra����R���R�`ͩ�6Y��C!5x@dnڋ�Mk�'�)�Ӎ{��*��f��u֣T�-����pl��m�JE�>+���V�I~y�O�l�]�HU�E�G0��рO�>���'��'��	.�M�!�#���O�@CR�*U~�{G���̀�K.�	���J��p�4�y�S�\�p,դ(X�ݫ�%��0%|hb��=?�WA��y�� ^ḩw|�Yv'T6pfdu3&"Q�;��q`P��N� ��>uJU��
�&�ࠇ�6mV\�!V�/ք� ���8 |����(Af���� T�q������O����e��&>"�b��ܲ,q�Q��(UԺq�|�W#UU��)�M�v�IQ!b�eK- +$������xł+V�Ou��s���?xQ��
T+v�J�[�@;s��Y@��6��@�L �vi�Ðké?^�}�eR�l��V%>�^LZ"��&J�a�eN�bA���NH�	 �C�c�d��EԠ{�B]kD
L�i�HE�i��L;kuNO����O̒Ok��m�*(�'	O�K�����׷���'t˞'Y�	㟀���`��ʟlA��hPYZ�ǜ�F�x��+�9l��'���'mҖ|��'lb��?���ٍ6T� $hȮOK�Ja�(!2n��?A���?����?�QÀ��?%d�*8,�s�a�;,o Mӂ	ϭsћ�'K��'J�'J��'D8�����M��d��s3LP�4V�3`ȸi'Gt}�'���'8"�'�|U"[>���5E���h�M�pt�Ү��yߴ�?�L>q��?���$�%���f�M_H\��ǎ��Q')x��D�O����O��م��O��$�O.����L��u$�!�&Tp���v>�+��i�I��$�ɘ֢��!�~JDf�.VƘ@#�߾N�*��t�E�	��؟��m�����qy��O��i�q�B�[ ��hh��6��qӊ�D�ON��V�|�1O���L���'��$a�]o���ij�l���'���'@��O-2�'��Ӻl~f�[��
 ���=B#���ܴ�:%ȴ.�{�S�OCBmU00f�`�RO*�iO\%e�"7��O@�d�Or�P�l�d��?Q�'����ƃ�!5P���B@�%ڔ̀�}�ǁ�Ԙ'F��'"�"c&8(�Ɣ8Ga�H�U	X7M�OZݹ�(X}RQ����b�i�Q!�GƲػ���/�
|��>�%��/���?���?�,Ox,굊�4?JV S��ݿ~p�c��(t��D�'��˟�%����˟@����^{@I{��X$Ew�a��� Fh��%���	џT��ty��A��)��B\�	0�]�O8k���}n��'��'M�'��'���[��Oj�2��N�&�ꗮ��7!��z�V���	�����Sy�̀1P��'�?	2N��H�7��.��E	�J�9`N���'��'���'��ycF�'!�Bp���X	Ir )f�x��@�Ц)�	���'�$A���~*���?��'h��R���p�J5Y��$;��i���x��'w�d�KU�O��������d��n�#�kU�
�|6�<� �W97����'���'��dj�>�q�? \I�h�$H��	��L�W����$�i��'��Л���7����hց�%[l��4@�no�7m[�G��}lZݟ��۟l����D�<ф�F�lbY��7��i�����RÛƯ��s��O��?U���?"L\����"Lh�A�ִ��4�?y��?ivm��R���Ry��'����j�`)�fbK14�Nus��^�#��O4$K$)(��O|���O����Ɵ5������a̺�*�A�ߦ��Ʉ:%B�J�O���?�L>�1O̘�!<ܬp)s��*U���'U�Az�yB�'gR�'-�	qBBԛu���ZE��/�|:�KvD����<���䓟?���Z���R���o(�}���&�ڜзK�4���?��?�.O���aB�|���^��x�_�k��8r��͗'B�|b�'~r쒘��	Jm�TAR���F�� j4�US��	ޟD������'(!�S��~��Jm���$҂}ڜ=! �ߡ'�xqe�i:��|��';�؇'�>F�Y�u�©X���������צ�I����'U�*aB>��O����F<��B�8��Y�[ N��̙��x�]���I�p%?�i���M��}0t	K����i!����EӲ˓hPHㄼiC��'�?I�':��I�?BUj7cұ�`šԭZ���7ͧ<����?�����ܴ;ܨ��4(S*En�Ԁ:Nn�o���Pݴ�?���?��'n����dM�;�Rh���u�h�q �"_��7-�O���O�O�s�L���� !��� 5ڴ�Y�e�=���"�4�?����?qC�޷)牧���'P����H@��
Tpr����(���'I�I#@�<�(���I�p��c�~��sl�U�HA�n��9��ao�꟬���
Ty2�~R��K��2���c��L��!;��O͜�9s� ���v��?�)O�����D��щ�:f=z�0ŀש?�N̂ao�<9��?1�R�'g�cԤB��܃�D8eJ�B�&�?"0n�b�����'hBR�h�	/'؊���x�`0�*�Iʲ�Q`��[�<Un�ʟ$�	f��?����8)�����! 1��H}vAZ�eK7 d�H���>����?	����{Jna%>�q�Lѩo�����N�)�hU1!�1�M;������$Q�{C
��/��f��@���)D�{��h��Mc��?A(O0IR�`YN�ɟ �s�as��Z�~���3!�"*p��k{Ӻ��?Y�"������'��1��ys��]��5���ׂ{W��d�<���Z�&U>����?�[�O�L3С�&	���N�5�n4���i剁&aT��&�ħ���ݺ���n�H��K�)x֍x�!c�~�I���O�D�O����S����m��\3E��?Q�@���͸M�,6-Y2��l������"SC܂x���J�2=>\�Ƌ]��M����?Q�����b�x�OO"�O�Ղ5bO�<6�93��> yq�i��W���w%����9O��D�O��$��XA�fn 
��S�%"�oZ�l�'����|�����Ӻ[q圼	 �*��
�m���sr��n}��J(s{�U���	��IWy�ÄB�tM�B��^�@�a�7c
�(�"7�$�OD��O*��?�М!��Ν�d�����-=�v���/�+�?�)O���O˓�?A��C���d�(j���H�f�1`Z\]	�lԻ�M����?9���'���D0�@ܴrjn ����$�0�r#�4b��i'�x�Iryb�'��y�Y>���$�,��ci�H"X,N�.�>�a޴��'fb�'*�aA�����[~�`�eF�/~�P5��@[p�Xo�ݟt�Ijy�K �?�����$�kl��s��z7@�R
��ucT��'���!R�n-�	q�SGj`d,n�X@�@8ѣ�ZR}��'4��x��'��'PB�Oj�i�=�!�/~b��㯊7�Y��@fӆ���O��i هT�1O���A#j�}	j^�9�R�pָi�j�aTBu���D�O���⟚�&���00�S�L�!>����P��гܴZ��|K��?�*O����I?U^~� 5�� `��pqm�Q!l��4�?���?y������?9�O< @���0.p�C�D
���(�#\~̓0�����O��	:_:<��n	�\�.H�Wm�h7m�O�9���<YE[?��?����1O`q�E��^�! �/X�L��	�lr���>?��?I����dצ0i�ŒBF��T��l	�O\?K�9���l���� ��C�xy�n
�/*֌�Ɓ��M]j�Xen�aL� �b�'7�	����ҟؔ'>�DF�k>�H�X�B0��2��+yY@��>����?�H>�)O4� 0E�O�S���&*Yh�Y���=T�e�@[M}R�'B�'��	;Q-���O|r�	ڪv:5�.�%�~��Q��*11���'��'c�I�2�4���D�I	�5��A!A��@|kq&>oЛ��'~�Q� ���=�ħ�?���a��!X�@Q�o�a]&DtDp�hyB�?�Ҙ��ٟ��y%e�+/�2䙵K�T����i�剚7��l�ܴ0���ן��Ӭ��䀚~)��ׯΌ1�H��jW���Ɵ��QfO�Ot|&>�%?7�$i1"y2��7�����	�	���CʲO�7M�O��D�O�i�b}bU����o�\���+���;�����_��M�$J�<�+O.��"����e���R��m�Oǵ6�|�#F�0�M����?���wp��R�l�'���O� ���B��B)H��@G�~��S�iXBX��K��}���?����?�BA�>@����^'|�T�B�
F9��'M6����>�)OX�d�<���kR��)��Z2oڷO�
�!%UO}R�����OJ�d�O0���<9�%D�{�|᥌]z���'-ɰ5x�]�Ԕ'i�Q������8k^����j\bQ�"�	�AC�|��e���I՟(������Ly�L�.)wn�S2��8e�O�X�1c'�)��7�<1����$�O���O��72O�)�B,���Bc��
!j��4!����ПP������'��ɸD�~B��`(٘v��(:��+B�D��9`Ӻi�2T�$�I۟��I�u\�c���*W4�@v��f��{�I�����'��\�FD������O���|!����;Y�\��e���L��I�@}��'�r�'�Ұ��'��'��^�>�^�`r��L��2c��h�i|�I�a�2��4�?����?	��!c�i�1��\�v<EPl�LyƕP�~Ӕ���Oޝr�?OZ���y"�	�g	�R 
3$�J�:�/ˤ]�vBM+Q�6��O��D�O.��G@}rT��K�c�7z���wH�#nP9����M��Z�<�K>����'���x!.�RPv����Hc�@2'd�N�d�O:�dW�4���'P���h�2Y�$�k�1�YY§�5E�H}l�ݟ�'1Ș˜��	�O�D�?�h����z�<�1b�3CN�4	Fe����6���'j�	ß �'kZc���O˻%����T�'��,b�O���$=O��$�O&�D�O��$�<��l�m �u���.��tSp)ˤn�$�1R�X�'�S�\������=��Qp�F<|,�̑G��+@��P!��q���IܟP�	ڟL��yb!�
2���{���1>Ȱ%0碔5�t�ٴ���Ob��?����?I���<�w@?
zZ��(8ထ���׬w!���'��'<�^��Kq,&����O�(�Ө	7ZJBT�V �5)жj[<�6��Od��?Q���?q�.Z�<�J�Dʃ��[�T)�,ؖQ���s�~�"��O�˓b���Q]?)�	�t�6k0��k�j�91������*B�zD�O���OT���/f�D�OD������kCt�8AFè'��cjQ��M�+O�<���m̟���ϟ��ӣ����4M�.��80��͓1�j��q�iT"�'T��'<���<���$���v@p���a�x�9-O��M�HC.%���'kB�'3�$��>+O��k�&A�:��hʅ�N��A-oܛvn� �yR�|����O�DRdNW����c)zK��-��޴�?����?ѥ��&��Idy��'^�ğb�����/��k��Ŏ#ǱO����$�O���O�i�ׯ�w���w�8C�l��%�զ��I3H�� �O���?)O���Ƥ���8 >� #�MA�P��Z����>?���?i��?-O�����ū�B�ãǖ�W��B҆,EY���'��Iן�'���'\2�ϊY�Ń��5��T3%�#�4��'4�	֟d����Ԕ'��Y8� s>�' SD%� ��/'� ����p�ʓ�?�-O���O`���s��A&1���s�ӓ<�)���P�R�m�㟘�Iߟ(�	Jy�ňz���'�?y4"��8E�7h]]�E
�bL����'��	��d��۟���f���f?�҆2Ml$ b�t�:�Ĩ��M��Ɵȕ'��5`C`�~���?��'~�t��7�L�G�t|�r�D�z0kQ\�8��֟ ���|3,��ĥ?��a�b*�8AT�����p��mxӎ�FV�hX��i���'+��OӶ�Ӻc�dF*P��E�!���`�������Hp*d�D'���}�w×5�H�����)��7����c� �M����?I����7W�L�' ��i��)%��%o����7�p�t��>O�O��?)��*2(�R��Ũ3�K6%��M2���4�?Y��?х��Gz��hy��'��I�(�Z�S���&��Q*� ��IQ��'���*u]�)����?��OK����ń�|����h��p��ڴ�?1��J(���syr�'C��֘���� U�U�O�.�E��Γ�?���?����?.O~����?5�44�C�]*5���i��W@���'��ڟ��'���'kҠ��07VUcb��+�P�Ӓ��
T'#�	ǟD�Iɟ��O)���0����2�q(�*�Xi�q�xB�'�'7R�'ih���'#t������3� n��ّ��>q��?i����dAt6$>u���3O�1�����l��D��M����䓾?���C*D+���I,[ԕsO�Ie0�
aI.M&�7-�O����<AhA�Y�Og2�OK�E9���{||8��J�
0~�@m%�D�Ob�D�',Mr��/���?ͣRO�9_����썁hKP���mb��˓f @[��i�&��?i��9(�Ɇ;:���H�*$@���Or�6m�O��	�6��5��$�	;���1gR�MCP�KA�U6��1�xAnZ��	՟�����'������@��<Ǩ[�ʐ�r������O�O<�?�	  �ʕ!��:򎝂�	��8p�4�?i��?�ӥQ{��O*�伟(�%ˉN�P��W��4Ug�@�6�c�`�O�ݚM�G��ğ��Iʟ�rBC������ɞTn`p�����M���3���s��x��'�|Zc�2E���8��u�B�>	h��O�8���ORʓ�?���?A)Obd��$4C�k���{;�p� �D�IbL�>9��䓮?1��b�� ��C�Ɋ&4�¸+#�Y	T��4k�<q+O(���O���<�c��:��i�m�މX��)_�pz�h����|��O���x�I(i�@�	�e�8{A$Z�Xh��7�Щ����O��D�O��<�w�I�#��O�^ ��!oM�LU-.,�rb,f����+���O����-$����#}�@�PȌ�C@M<f,�T�0g���M;���?�/O�t�2�h�埔��P�NL�RL"`�&�"'�X?�8H<���?A���<iL>	�O�mPu���j��0�%B�L2���4�?Y�������?�(O��)�<���.�Jw��_ш[��R:8�o�ş4�	=r���h��8�)�CДs�T��hE� �T	"�72J�z�n���(��ȟ��S��$�|��89�n��T�#���d���sԛ��43U�O��i*���O�Ȃť:��m��`��
�hqC��������I9N`l@�'��� �v�d�#�JÜP�8�����c�2)����K����&>M�I<�ɬ|�0E��ɒe��{�� 7�P�4�?�����?�o�����'�@����j��t��N�J�P�EJֳ��DԊ61O@���OJ���<YCD)�������N�q�Jр6ײ���x��'�'��	�4�I�G�br�	:������"#H�I��b<�I��(�Iry��'z��Q��d@��	��NB���m٬FY��B�i��ş�&�p�'���+u�I��Ms��
4]u4q:3�Z8+�A�l�~}�'�BY�X��Id�~�MY=y�:�	�	#B�1��ǃ�M������׻o���5�x�jE�$c�,O�$&X����į�M�������O(��R�?������j���2%���HF1[�G̥�I<i.O�sӇK�K1O�STݪj��#x�V��cɴ6��O��D	�<;J���O������?��:�n%�P�Y����QAW�f��Um��4�ɾ4,�"<!��/�'�mb��?]���P���	�M�An7�?Y��?y����,OP�'Q����.m�ժ�8q��ictl���?�Sݟ؂Ǎ)
F<T�õ#�j�gù�M����?��h�h�.O�ܟ�3z�8�u�^���I�&g̙`~dm�T�$\To��%?�9�@SnpH��i[.��w�
���<Q�l�#Rpe:
�'�Zx�ա�$+ �}@c�[����:דU�T��n (m��1ɗ��TXni���TXf�!ѩMO(0 �c��p<$������Q�  tV�h��Č�`0�`R���t8Db�P�:��d�V�]'C-����`F)�re�iJx��d�
�f^�"a�U�[` �I�0sLD˕�J8(,��l�q������&n��Y�	����c����,���|z��U�h����l�:Y��a�a@Ly��=����ㄈH��?������	�Y�i$���>I!�͉>����@F��<B��)��i�&#�>dԉ�N �9Rޕ���D�'���؅���!J�ѩ=����yr�'� ��b	��O��XK�52�z���'�6Mȥ����tEQ-a3j���$�0��D�<)�I��"���֟�O�Y�&�'�q�n/2c�|��x�Z�'�2g<%�d�FK�A������O�@��d&1J0�!�(Є[�8�ر��I4>kd� 柨s�X�����_�O׈aP$��;W� "g�����T�J��YD��Oz��<�'�?��`H�+� �-�cwɂ�}���ȓh��R�.�%4B�( �ױ%w ���I��HO��H'$�<i,���+*J��	{dDIk}�'>�B_�`Q��'��'9�w�"ȣdL��0�4�a�B�m0�1�莴l�x�C��O�hx�e���1��'�Bm"���0��H�)vΊH6�خd(}��E�O��tJE�����LR�!�&�E0Y �'��|g�S�����-��O�ў�R�/YD9����-L����8D��L��?�\��)��{P��g�;?y��)�-O� ��.е��(Jq*3L9�P�JQe��(����O��O4���պc���?A�O%Jik����Db�"z�L���Dې�x2'ʜ�]i���g���*�f�!A9�]Ru"�3j:����15��#�!�=bFa{���;���M�m�:�c��U^2�����?y��$=��%NNz=*@+�	L���X(_��@B�I�a�JMK�lM0���Ѧ�]$0�c�h*�O@�	>z�TZ��	6xݢqZF� LY�E���a��M�	㟠)@�������|ڴaT 5�ܹ��G^V��u��4r������u��c�&�)�H���0l�#Un���+#M�)�� ��#��=�4��4\�DQ��+O��
��'�bR����I<H�@�23��M�+,��b�4�Z@��n�.b����)�_xB�I�M�`�W(+6�$C&G��)L$)����<y����_�*�y3#�7Gg���*�I�&B��8���A��-�rHS��f�C�I-��x
C��%K�f:��L���C�
`7~�;��GL:��A�)�!�� *�CQ��?_�H��c��l�$"O�(iVi\hX��K�$�2��"O&�)vk�"��l���&"���(s"O�����[��a��d�Ҥ�ʕ"O>tKFh_X�𴣵�J&4-ۃ"O\]�P#Y�4�N�H@�� �rh�"O� i�dϭ.�,�(�X0��(��"O�pX�N�(��Ȳ�Ş�P� A�"O�`���Lޘ`��]'e�4�H"O�@�Bb�j��XtI��8�|5Y�"O:]C��m�����e�(|R"O�P��50�s^�� $@1"O���f�R�5�>��C悲X	r�j"OF�c�k�Z��P���+h�i2"O"�ⵆ1h�
r3��L��KE"O`t�ԌJ93�ԓ�팚#LE�"OT�!�i�-0��)�W
�+_��"O8�0�l �J1����S�"O0[#�X%4�^�!����1E�hs"Ot-�K�:Y�4�kc�U�fX�"O��w��14���ztF+_(��G"OT�`���U������U�9@�%��"O.e�0�2Ρ��C��\��Ĉ�"O��p�#F1��Al�I�HX�e"O�0�ۈ�Z\9R���*B��ʄ"O�`P4#S�hV­��OC�M��].�y�
�8x`��/Mv˶jքX7�yr�J�a~B���Xm5�<��l�-�y҆\�(�B8%HY��Xǁ\�yrH\�E`|y��2�����J�y"��Y=X�g+���Q!f����yb�Jj:t���U���]��y�	�lm�-c&�ڧI��T �-��y�˓2Yf���E���q��y�)Y�td�@�Q��=-��{��V<�y���9D��Q�%���\���	Q��y��ޤz�u` 䊀r�DKp���y2���~��T�%j˞��T#��y��I�l��Պ�Z��1o=�yB(^v�z<�sG
�t.}�U`9�y"�۸F��IE���(�r�el��y��A�~��s�J�/(��tB5���y戅�<�sB�,�<�T���y"���>����f�r�����p<����&�qO���t���"���+�%}g4H�B"O�-)$˝;�&ip2kW+~ZP ��^����ٌ-�b��|�䫝vgF�j����t��<�@�Ju�<1�kY�-ತ�l F$E�q�dY/FY@�J"� N8��#fȿR�����ń�HR�7�O���q��`�9�LbH�3PH�KT�є��'(ڄ�0?A$�¢? ����nOX޹	���x�'cȠ�� ;�:����7����O�Q[��1q3rڦ�L�
�f�'n-4���d�.Z؁�0J�	y��h@W
�O9⦍8O#t���&�&4%���g}����o}5C�i��o�*���I4� ���@��X Q�+>?�y
Sʛ�SZ1 �%Reʰ�'JN8j�P?7��/%�J��
t��F��r㯁�(�b4���=�O2�j-͛nX��oъs�fx�Ul�]�>��Jڼj{�:�g��?ّ�C{.�����R^���ME�HMiԮ��OQ�L[��	��^���E6XHLkЦ��S"ku!��%�f)�Ӎ#)50$�
�'B��ЗM;d�� �\0e��X !��)=Y��A��Q�Nr�Q�e�%P����#&́�&3��Dg���
'ʓk�`4c��S ź�;2�Z�J��D��
'l���V��Y�	X"@��c�����&^$
*�%b�(�V"'*�m+�&���|�Z�� o-�c�b>�K!�T_;��ç@K���3S���77�����CŴ�85FPs�zw+�H��:P��� @��7��p��h�J�v1��p��O֠+w%Fq}��	P��̱�M�k�����M,���#��yHV�V�M��y %�>��8��捅`�x嚌��*E5���}�0���O�H,�Fj�1?��m�0f�r 0�a �\H�2��זw���OX�p&�ƴ�ywɕ��.i2���d��fR�b�b�<i�/�'S2Q?a� �=jLl���n7��&Y�@ܡJ>���	P�3[��kC�˭F�r��w����艀G�m�V$ X��N��(�>�~r�I�%����C�Dԫ�J�2W�b%t�U'�N�{�@U�~-�-q� F �Z�s�╾Dթ��D�7=��HA��:z�du�#�";��DNV���'�]s�+	�p\,��SDF�{bz ��'�����X 75��Z�i��?�X��#`/М%0�C��O�Ⱥӎ�}?a�MO�Tu$�z���0�Q���Z?�'�g�j�	ρ:i��c�E_��?y���P8����|�M��m��V�BL�3�MP�'��$ATM+���)��ؐ<��8��܆r�����!�;�����Nm)U�	��	�'^^F�݉m%�@C�w�*�K��O%un���I��4������@&�t�>E�T�F�))�d�T� ���s�j� 'Q��Pd�X$
T*�p�� �I�e�D`�'
L��&嗧 �>��uH��z�����'�,%�t�7���dT���q@��:��ӣȄ�)~ ّq�\!T\ա��y�*�+��=YإQ�e�'ԨOX�G�?��R(����Y+z���!ky�ɓ4b0�K�<28�@��VW�6�^>f>`��>��`�ת)�2�1��	-n�<���	�aiV#*��a�)��I�1|8��4@��0�I��}T�ÏÚ
��X�C�g~B��k����(UX]i�"ٿ[D��H�~K���7�BV��]�E!
O�"e�[�n�Xs)�l�頔��p<�DXm�,�0v�vl���Y���Pa	)�q A✈eBB�#E��v���煐�J�$�X�	��	#C����$��C��=���A8#��5 v�ɖ�1Od4C��Фp ��8G��H��1Ο�X�(�.���D	�]L�Z� "@�`C�ɸN�| ��
�	F-�`�d�\�7���r�"m �c�J�FΕz�!��l �W
)�'>���gHK�X>���Ta 	̄��"Od��ň۰q�}Aq�\�90M��E�:L8M�%pN�+��$����O�.b�(qe���[�$�s��BZ�h�{��5LOR��c-�tx�x�F�;Vܐ��D�<aj�v��DΈ��h�-���]������T� i�����V�(��)�8~�qO���m�ezJUH�U���O�Z�K�=;��rޠ�Dt�U�*�!�1x��a/ܚ�Ĩ�v�]�V��I�q�r�1�>���O[�h�¢��$�L�k̘֭G�P�0�'��j\!B��aQsN��*�MH�yrF��n��l

�ؾ ��-�6Eg8]a2˞�z����RP�EQ�v|�Y�&�x刀Sv[�����O��cf�T���s"�h�V��㉻i�B$
��ĉ�r�����E��|t��bFO8�!��5����U�՘K�=@ '�\��'�,d; @/�)�ӠF� �n�>$~8h�5+έu�fC�C2�` @Q�M������Lj^C�I/C2�5J5��|�ـ��;�FC��%
�����CH�C��Ⱥ7�	�h3(C��4K����CE���թB6k�B�	2O������Z�<�h��3u��B�	$;�����8��1
���&i��C�	<n�.�YRlܳ-����u�ڳ^��C�ɬI/�Q�	7���{2`*+APB�Il���D���(�,�x��
G B�	0c�%ʲػ>�h�0��-:C�IzpM�%*k]T���GP3>� C�ɛX�t��s�Ѻb�.�ハ�VC�	4`���L r�ԙ������<C�	�z�T�]�i)�E��c��B�	?|�F�:b��+�Ϟ�c�C䉝nCr�㬐�xx�t�W�6͚B�I�c5"X��B�v%
��ՂR�|�$�F8tz��' ��	j�����#v<	�hIh�q�aƁ�y�O�
0�ꔡd,�#i�R�١�ԓ�y��|�L��둈.D���虨��'9S���?-�?)Sbэ[;t3"�3���P�4D�L`Ȓ����Iv���K�'ǟ�y2rbx��]��~Ҡ�)c��&LI�:��`�����~��5eB���� �HC�	�LbT��DhG�2u���'�����F�)L�Q��k��_�~�ĮH���e(�*  Lߪ=�Hi��DꁯZ��	2y�撟����'D 48q���	�t�$��r6�ʊ�dB�(L0D�OQ�2+�R��:�6ͰC	�'Y��j3��)!&8��k�?�0YҝϘ��i����)"s��>|����ځk��H�� �ا�:t��7�ۃo��� �?W��N+%w\��f��=!�Q��t�1g;qa���'Ϣ���B�=�ȩ�$�;q�8��xX����O����U������J�9����9[��B��O��+D�f��$�r�S s9ᚰm^�fHD@(�M0)?���>�(�Tr�I
�T����D�f�δEy�M,�D�~
SN�^��0#�l�R`Zaht��4�Dm��I1&�vM`��D����F�R�bXh1I��
��P���	l�8���T>y(�I����p����?UR&��;P���ar����0z�C䉆s\�����ݒ6%��C��L���	.熔i���Hl��6N�;*�D�9O1�j@w�تf��i �P,G"<���'�T<�p[�<��-YB>9�0��;5@�%��kΜ?т���8��h���E��O*0�O%u�Xpc����5�yI�剕Pa:Cs�S�g������ɂ��L��U:v��T�)��A��(�����ئ*Ɏ|���t����M����ا�	��d0�`@@A����e���
7��y��
<�\�ȕ"Of��D�S����[Ѧ�@�� p��'L(�Ȁ+ɾm:9Ad�
 3�v����yJ?��Վg���P��?3��)ά>%N�8ӓx�|ÔgW]?���,�^�(��<~�*�΍�2P<��6U��ϓV�̨�g�'�D�wi-f@�*gA�?�4@Ӎr�l�(�����ޙZ����S�<Ҡ%BV$�u����(]�:Mp#>٧B�@��� K��ȅj@��&�*��8S�L�J0�ˉX�b���O�m�Ն&u�����
D8`��aH1����4> �=�l���$� h0ܹY�f˜ �]Kf�ߔ!��Ü�g��IR߷`n�mY�*�"�����禥"��!QO�� W�ʊ/�NUA��S�%jL���ˈ+�^u$�OҼ�&#Q�3�X����+�(l��"O�T�� ܗ(�ĕ���Fz�!��	;l�x�a ���0g�-a`���@����ȓCHh���J�pLБE�	�����9
�閯�:jL 	 ��:�4��z�6��� ��{Ծ�x����E`��Ql�Tp��ǫ�(�x��C�1��|�ȓ��I�� �FS�8�<!����"E�	+��O��B�ܝ�yr�T59}n@��쌥z�D4crAB��y�	��0�`c��fD��*���y���1���l��cS�Q���	�y�痤2S��q6i~8����I��y"K86�)��J܅�d���@�y�DIS^������q�@�K�#��y���!��(��C[/oՒšAf ��y�� *wx9�t�H1d�*�q��6�y��_�n��&E�D=�����,�y"D �*0��P���<Ř=� �Ī�yB�K�~D
uL�41N�P��y"�Xy���� T8_�r��)�y��Δf�L0�k�8Vb4p*w,��y�.�(>^ֹ��Ԉ�5"aU��y�ϱ=���-�0E�rͱ0c���y���np���O���mI��&�y�BA!~�|��#��u��Y�yBm=WJ�U'�(���a=�yRcH�b��Q���N�6%$��y� N�I��ٰS,A�^�v�H���y"ϙ��ޅѲfW�V�RA�7ؖ�y��Bs���	[�B���l?�y�,�0�
$Ђʄ�ZT�����y��1?Vl��އ��кCX�yR��a��Y+��	�v���ԇ�yb$� pޚ�J�	��n�S�L���y
� И��(� -�=Kw��:\�X�"O��Ó��7���Rb��O�>hs2"O>-�"ͿM�D��� �`�;�"O�ɠOѻ3~9!c��-L��m�0"O�LKA�� x�x�!o��agd�H"O29�ׅ^�0R�"A�՚d`|��"O�E�'eܢY�:�Ag-��qs򤰤"O.�1nZ�9Ij�:���H�"O4@u��$Ed�	*�e�x�v,�d"Op�a��qB�2�ᑹ��5�a"O4�L�?��a� �9T��B"O�UX�F��v�V��Woۃ{V ���"O����W�N�{3�]
E#F9��"O:�zTK�B1Z�c�ylr�"O\� #ɋ�'pm�DE��1���S�"O�xX�ˌ�}0�]C��Նv�(�u"O�����?��H@�B[��-�f"O�T1ԏ�	uM������4�a�"Of�S�]�-���*%�0*��Q�"O�uy�l��E��E/^�4u"��"O�}3u�_"Vd��#$\C]���"O�M8b�Zo�q)ǎ�62=T��"OܙB�+8����ц{"�\*�"O\��)�&.�]�1hڏe"U�v"O�Iv-O�U��=��D��s��2�"O�Iz���
�H<pt�̓\ Љr�"O��p�G���A�鐴�"OP�A�A��m_
�y&�V��X!Q"O�4��F&�щ���>p���@4"OFи���rĒ%o�#b�>�B"OL�7�g����W��� [3"Ox��T��h�Cv�ϝX����"O�\���!�e�GD`�)�"O�P�̇,B�ʳǓ�v��Y��"O�4!%��e��6'ާ%�����"OX�34EWT�A�HȚ+�؁�G"O��QW�C:Vp��F���"�!6"O��0Ѫ_�H��w�9k��2w"OrL�P�	�бs'���\0^ثU"OJ��Q�\�{�<�҂Kߡ)�8��e"O48��V�7X )��i�@Sf�A��|�)�ӎBL�s�3@�@"G�Vb���ȓ�z��a��yĮ�>$�ȓ]�03a��U��ᓧi�d���ab>�R�e�V�a`�JЁ���� R�y�ǚrxXY��G�~�q��w|��7X:�*@&�D���]��
!|�`lA=%Cf5@Fmɍ���-fH}`g��" 8�C���w>N��b6�1�����-�5@�&N)���ȓp��]�a�Ɋ/j"	0��КE�ԆȓKn�����Ϧ͓�/�=�ȓsG|��Q
5o���YV�Je�t ��X�x�0vƋR��S7�8&�\���@)<���$�� ��5�J��.܅ȓG�PȚx6�S��v9*E��6�&��Ř�#�$A�Q�.$�d`��&�<!�V�̨��x(��=�)��;������#ai��hQ
�R�섇ȓY "H�'抓�&�v釾Y�r�ȓx��;�/���]��ʓ.n�1��-���@篖�s~J�)OӧQ�ɇȓjE5�3n�p�!��M�����(YM�D&�г��Qn���S�? ���KJ�@�r��g͒O8\KF"Ob����D%: �Q��,��t�8�S�"O ���U��6�q�,Rp���1"O�Xˆ���`�q�+?RZXX��"O"�i�GH�HHS2�5(A�!"O�� 4"�;(n2��_
4�j=pr"O��鱄E��3G�_�X�,�zA"O~�+��^�O�n:�G˛W�4�`�"O�y��Gϱ6\<�5LGH����"OJ�C���
�41�H�6<��Q�"O��yC��zO�x��
9T��"Ox��M��I7�}ˑ'����r��'K�<[��T����O�� �b�(*D��ke��+�m�̉J��jD*D���&��"���(?K��!S��)D��2T�\�=Z`�c^Q���4D�h*E�1<I��E��S��k�N5�$7�S����څ�	OEz4���ݿ�N��ȓ;�6�R�X�驁6)� U�ȓADN1h���;,���A#$�/vq��ȓV��u��(ֈ{�H}���P��!�� 6\�s�A�b򔵰��rC�ɠ+���V�MGl���ї`��C�I�6�}��%��Ik��N� ��C�IBdZ8�ë�%t� ���E��C䉔+B�#�\9!D�*Ʀ�\>�B�I�VXT(����\{lHg�C�_g�B�	6�J<#Q�W�y�J	2@����B�I�Bu��8tF�[\<����&8ŘB�I�f���b@�"9���
ςw�lB�I�z+ؤ��/�!���uN�qb�B��4Z-P<+�Aˊ	��/Me�B�	$�4YI�1 
��G��X<�C�"g����ʋ�w��������;ͲC��g�lH�S�s��\�&��l��C�I�X]�x�Ek��"��HL%6^tB�I�'	2q�c�w��D B@�\�jB��$����&ś'4��F�8�FB�'_"Z1����0-9*k�L[�<\�B�	o��p%&�\�x����<�pB䉫&�򈚦��-}p��7�� ZU:B�I�K�j�U�H$=v�	G��P�fB�	<��!�	B��.��f֥\��C�	�;�BTs�&���j4!bHڇi��C��2\�PD�dB2���چ�W~�4B�I?^�,�P�ޅSG�H3�٫WMTC�#^
I�C&�'st��4
��S80C�� v� PY@�ݠK(���C��,WP=���N�_�eS4��U��B�Ɏ⬉7���zC2���Y�",�B�	�3	�p+f+�(j��(#�[�|�B�	OTp
@Z�ax���j�AF!�dB=~0P��.G:&g��J	_�n6!�D�Y���Β򍒶JR��b�'��$��D!B� ��2���A4�'a�M�d�ߍ1c �Y�G��9!�T��'k��1`L=e>:����՞���P�
���h^8q�:X�ը�`���(,�\��	�
v��u,�>��ȓ6�b�Ӏ�\�z_0 w,H&�LD�ȓ$	��w%I-1�ɳ
�s2l��p�E��l�6��I��iY�6��<�ȓ���z���5n�Y���P�[�"�ȓ040��G�?Įi ! �&8 씇�S�? �cp�Թ{\t�8#B�C�H���"O��K�A
=)�ԐK�I�e�M�0"Of	FO1�4P��FL=c~�h�"O��(S`��,���S� �Q"OTqJF(�&`LR,���ʻ@;�x�"Oh�� �C�<��eMK�?􉐦"O����`�}4���N��a�����'ޱO�xRE�@a�92'�
��]�"O��ZRDY��*�3�4L��"O�a�R��5`�(��P� ��Ad"O"�!�$�(����p��[�"Oj�!&���r�xع�]*@�
lA"O^@��ˈh(���\����"OZy��h�b���3�M�Ht�"O`Z�̈)FKr���ިJ�Z�"O�Đ` �	?���ʕ�_�ZB���V"O�@0�M��LI�p,�W!�%��"O8��&���0�Y�f��~�Q�"O������W����$˃�+ȉ�"O�U����>��)�	ӈq�H��"O��IfNG)��1����|�N�*�"OJ-�a�J�uax��a��Xˊ���"O�9	�*�z�t�M���"Or��s�M��D7�����!"Oܭ��A
j\�m'�ϽAϾ!��"O24�F��*M���85��h��"Ob=!ī�6�	�	��N��[�"O<t��kZ:����D���1d"O��k���)���SǕ>�d�ȓgǒ�@�Ϗ"i�@a%g(^~���%(1�����l
��I�>��I��LZl�CsO�.7n���
4�"e��}ה�Y�-�l�b�A��Z�R����ȓ3��tYKؖ4�9@�C�����=�$���F�64�Ā�<�8��ȓr�22��Q�u�(ib&�-Bq
%��?��ȓ��[jh�b��wY�ȓ�d�!	6��k�͊(C\���VU`%�bA�S�����&
�Nq��y��)hG�ՑC m��]!c�",��w�z�֏K?SY��J5"�^�V��ȓ?}�E(3F�*��������B�]��b(& r��<Q�S�ث,:�����ׂ;�j�PA��8N|��iǍ�F�<�%f�9���w�ϝf���@'c�y�<	�9Z:��6��O
�5� �x�<�"��d��P�a�7T��@A��K]�<i�IT#İ�2�L�8]p���W�<iuf���<�ңjW�Z��� ��~�<a!����ѥ�#P8D�"2�S@�<Q��=l �e��/�(=���z�<�CB&1{Q�#%�5ߞ��`��_�<�V�A0�D�(c��c����1 FX�<�6�Y2-�{�d�7d�	Vʏ~�<1>��K�	�1eA*�q �y�<���O(��@�a�(W��|a�$u�<ч��+LQv$����xyyU�m�<�4'��0Ip,��x7q J�g�<94dĚD4���Q��>L)
0�V%�h�<�bN��W_��h6�O?6�PX�jIN�<�2���Q�v�c���#w֐���FH�<)��#�6p����+�\����Y�<���1. `y�C�RNh�o�A*!��ҬLVhy��c+d`�-*���G!�� ��@�$�8��1��)Ԥ�8�"O|�i�k̆J���C#V�'�bH��"OB����4���`� 	�S��!"O.l
�G�o���("J]!%� �"O��KD�q�!2��[�]ĐHw"O�L�U �2�=��a�I��Ԙv"O^c`l�$t'Z{��H��X�S"OF�b�h߶B$`���΍4Q���A"O�����I�5z0��RN�1oO���"O��r��O8w��ȃ��/G�tj�"Or|��C� D���2L�pԜ�b�"O���s�ԲS��|BQA��yK�"Oژ�f��n���@�?U;z��"O��@�E��Wb2��v%ÂA*�X��"O�#�iT�Sn��#E�\=�p��"O�UX��/0�0��QDTa\Z�ؕ"O0�y4���,�h�mMt�b�W"Oȼ�"K�2��Th�6A6T��"OP����/G3����,��H��"O|����r�赪�(c��	�"O� `� B5|�L�Y�&Έb��K�"O���DǨ����^���)w"OH,���74FJ�vj��X5PP�U"O8����a�z�c��-)�k�"ORĳv��
o��Ѡ!��wF��"OJ9����
��3
��o����3"ODd���):�pD�6I��`�t��"OrA��T0	*�����2$�H9e"O0�!#C�eDx9�aKƟ]�e�e"O�Aࣄ q�|�&j�	>Ve��"O� �l�|���8���{���c"O����#)��C�S��m"P"OJ���4�0kp���tE"O¹Ir�<l8$�	�̈�k�I�g"O88�V����i��E2D<��"O���w��K>%�7�i�UJ�"OMPԆ*�t����2zzLa�"O�zGr�^)�GA�c� "O�qj'��`�&i[R�[ib|e{S"O��򕦟Q��Ѣ�_$k�j��"ON�*S��|5l��RÚ#(��r"OF]�̍�ƢuS�T�c����"OJ���"+p�2'HU�{�0"O�!�̞�0	"T٠��j �!9�"O�eA���.�����'
�u�. �'"O6�hf�)t�
�u�F"{)ND��'���#a��C7���$��	��|�'��\�D��n���
I��|{���'��(��&Bur ȵ)ʇ~M搀�'Rĉ����?h4���v��3�'Q���s����E�0Aq�f1�
�'b8!Pb� �M;�X�`+�7}G��'7긒�GF���UiM#-ehq	�'k�����62M���Ef�+G*�0
�'���u熺T�2��`�K�(�@A��'=�!��Iˋs��e�2�'j	�'�m�U�e� �9%����'.(`�4�Ɔ ���I����,v)��';�!��פ;��X����6,|��'� �����,g`85#M�����'��򫘅+��i�c�:�dj�'�� Bfa܋L�z8�v��,�u"�'�D8HuK�VPZ�rV�δwݨh0�'��y��7BFDP���<vޮ,
��� >� $�"���'HB#�V�2�"OKg�$V=�� �-C�1�2��4"O�0AC�[<�)�%b_�a�����"ON��U���5�P��qQ*�""O���AJN*,�@a�r���e����"Od)b��uN�� �PZ��"Obm��.��vD|��.E�	@6IPP"O���#�H�^-�<r��_$*=h"O�(�F��_E�a�"�6I���"O�5��J֬(S-{Q�:* ��"O��0��]5:[(��M$G=�1�1"OĤ2��:Z���@|���e"O4X�Câ6���K��ȳ7~��Ӑ"O��XCݺ��0���N�Vc�q�b"O܁ �`�{�e���[�2b�1��"O���Cƽ	�f�"��2t^̻r"O�X��[$��a�F����6"O�iKń��Q���s�$��]��I�s"O"��+ >��3�$V�$�w"OVyم�I�M���
� ]����� "O\��F�: ^H�1Q�Z�fh �"O"��#q���t�[����×"Ofx���H�j�y0 %7Re����"O�i�nަ0o�p�i��4Q�C"O����E�&�u�G�C9Da��"O04�PL�I�Y�0��1A؁c`"O�)P�&��A	�e.F��P"O.�H� S760��ǲ\'�
"O��(U.S'��� P�<!�"O�84 �N��9��h^�9�"O@x� ��2%>-�����&��"O�0�C��60�$9S��~��г"O
P�h��0� H�!��$"""O�1��¯]��'�.��y�"O`�� e�-$�2�)WdL��4Ia�"OZ���GUC��puB����A"O����W(\ΌA�
�S��da"O� �O�Eď�l70� ���"O�h�dMS.�b�z���zy�5�"O8�mš-�ȩB@K����mʳ"O&�۷"�5'h,��
�1�f�p"O���'�o�&JDǒ�8̰�q�"O PJf� 8�:EO5OrA#@"O�5"��q1�x�ţ��Teڄ��"O�HB�Ǆ1)-���1-[�-L8Ԙq"O6s�O�=S�	�7��-8|l�"O�zGi�j�D���*7�y��"O8�Ѵ��J�6�vǘ��Ի�"O�
3/�8s��J���p�V�a�"O�1Q�k.6k�LJ�Ƽ+�6t�b"O0���+'!bej��޼3�dT*�"Ol�1W�ɨ~R�<�GT$Z� ��D"O^��Ǝ]�)��i��������W"Ov��ue/^xb֦\!����"O.I$�����J�ʹPq� k�"O���CɃ4��q���o�ޤ�f"O~	��\	i?<���p���B"O�e�?�4��͖ �<���"Ol�C�����8RbG�_%�!��"O��Z�:=�L�9���7���"O(	�5>�j�A3͙#<T�ԩ&"O���D[6a�*%�"X�SbX��"O��t��2D�l��`B�[0����"Onl�e�I0.A����II6#�\C�"O� \Hz�`U�k�`���2���"O^�h�P���4��M�d�Dp�"O��, �i��T9�Z�<D����"Ov��wIF:�L
��S	2B�F"Ojt����	Wc��P4�0��:�"O���"C�w��#�Öw�N�%"O4�[��۬��=P@#�0F9җ"OX����=�D��#��f X)�"O~�q��Af4
	�s��?Pd��#"Ox��C�_l��c�.�''
�����c>e�d���x�d`�.�\ytЁM:D���&iԒ`σ
Ǿ�� S�y�!�d�2!x�r��/ �d`Ѯ��0��'�a|�d3Lcҡ���7��-��BU�y�ImD�II�Ϝ>y��p�c�.�y��ӈ/�<`q�C��T0c1.��yr��2W6l�[���)�l������y�WR^Q���2?2�B˔��yr�M2S:��"��	�
� 3aN(�y�A�l�*�S�,��eO(҆� ���0>9`P %;@m���6��̨u��d�<) �
�N�JUDH�7���v�_�<�� {ʦ\r!��4;�\��d�<����~4x �Y�Fo�3�Jx��'5��H��ғ/-� Y0Yȥ�	�'z��T����^2z�ɋ���$3�O���M�;&�H#��c���5�����2BtXz�a˭;d���#�O!�$_�d����$
?'Pʑ�5gɼ�!�D�Du��٥�U�~�N06�ΰ$�!�dZ�:e&����2L_�� '��x�{��'��I�m�j�j��ȧ�b${e$I�3iPB�I�~�v1Hb�0"Z�9s��6�0B�IO`	Bqn!/<"0�C�G�d\�D1��]�O��2H���ږ�];�i�g⍭o!�D54�f��w�þF�R0H�6�!���#��x@���r$�Z�/�!�d�8���z�k�&a�xݙYaصϓ�?����d�#p�:�/�SN��EQ2 ~!�J�T�Jͨ��W�\�t��f�`	!��]�E��!SmA�v0dQ�-�!�dt�N	��3s�@�k�A�!�Σ~R�rvi�&D���8g��*�!�A�\���(��W�pؓю_Z�!�Ęqk
�p�f�v��Y�e��<�!�*_���"k��U��]`��܄?�!�$PS����6A�����	�M�!��ͳ"�E˃� �+V�5"@�!��$w�~����VVP�a��&}!���5�ȴcE��:r.V,q� �%k!���[���J#�Z1'-�5�ǜ53p!��Ćc�=�D�?�<A�"�	6d�{�Q���L�HP�c.o��ܑ���
=_�8�ȓ�
�6$+t�h�ӧ�օd�nh�ȓ��u1����k) d�S�Ţѩ2D���r�� �4�BQe�l ��l$D� �4�5$1L{�7-ʀL 5�<D����E*wd�4�p��I:D�t��-K T3 �R� E�af�
��$D� �T(�D�6M���B�d�^�pp#D� ���׈a�=��K6�]�(3D�tH��"$
r�� \����>D� j�`^-&)��́y̤��b�<D��
iٿ:�F��4&^@�>Y���;D�� h��34*����l�?4�^I8�"O�5����%Ǡ�pq%H#_Z!�"O~P�RB�Cq���qĄ�pL$A�C"Odz�c��p)q�Ӛ-$� �"O�1c�B��w~��uaFPp"O����&��x&x#F� �,��S"O`y�!m�
W��C�g"E�I�"O���U'WqN1� Y>GW�ű�"O��qCɄy��(ha���y��ڵ"O@5�G�1�MH�	�f�򈢲"O�ͱ҆ɭTa�X��gŊ`UL���"OJ������څF�)X*�Qg"O|��t-IW؎�b�D\ L���j"O�`� A������"�u�:i��"O���eA?��6e�/F�v`q�"O�(w��X>@b��D�d{ � �"Ou�4�)G�5�,�$
���"O��)�� ?<Ĥ�	�#c����"O����$ɇDf ���hڍ 0��{ "O�	3k�k��q�h��g @��"Ol���!
|
���d�R�̭qQ�����!V�v@{U���6�����a�4C�	<<��� A͟d���%�V�C�	�7/A�F��B`�)H�
VӲB�	�}sԁj��\	�Qʑ�� ���`�@�xdʊ$��C��F�-���D�:���h\�A{e�W"�P�ȓYuƩ+A[D�^i��)�I��4%�ԇ��%;��0a�N�V��}�5���Q�bB�I$i�P��W Z�p{Ul\�J�b�?����ӫ��yg'������-�'��{b�$dd|P�F�(-��9�!G�_���IN��8��eT&sgbd-40�`��ѭcUB�	.1W(�!'t�e�VI�"S����<?	s��v���0�e�6XR�W^y��'{f�KV�t�\}[��ѱF��UK�'P���C��!ub��JA+ �+G�hA�'�����6����%_(�,��
��O�d��G�1�b��5�ށvk�U��S����	�6�R�A�-�W���ɤ�ť8[,B䉡n�b���1�l<���&cf��$$?Y�n�Rnj}��/ņK�DpQ���t�<��W&H��u�d�(��uSFk�<ѡ���SԌ�T醋z��5QFg�hx�dExO�5�C��D���sD��hOjʓ�O´2�˃Q{6`q��T�5=h�_�Ȕ'waz"& �O-Z��U��B����[��y"�U�7u t��nC|���C3�Ԗ��?	�'
�$#������})��D38���'�.y(cʁ�X�����8'��p�'c��ٓֳL��d��fD�1���3��?a�y�(��*���+B/ۂx�ިsCɀ��O�#~��gL�>̌Q�;t���s�z��M�̺�Z�28Z�l�M!b�q��/D�8P��]	��L�ǫE����#D������~�0���	�-E�i0��"D�4Yъ�]&�1Wfć`AXDF!D�TAu�Ѝd��	��h��^N6e�č4D� �@��6}?*��H�/�K$ �O��0D{�O"���'���Y�s+�5 HA3L>�	�A�X�Z�F8x�b��d�ȅȓ*��i�,5���hw����\����bXA�o[�JD tP��Ғf ��t�$D��X&E[�2?x�C$�ó�*\�d7D�� .Ys"��>!��abbŝK�p���"O�,�Q��_�z�s@j��Q$"O��+ �:@h�J�,[:z�,��d�Ir�O��A� �A��D��"L� �'w*e	���%�ջ�� �\Æ��'(T��q�?��� �S��Y�'��]���T��แbN��a��'),�c�DATG�D1�	Ħ7�`%��')���-].+f�@��.j(���d>�"���j���E�&�\!p2�X� "O�f.À[㐄ɰ�� t�n=y�"O<���<�� ����]; ɓ"O����!�B�(�����	7��zc"O.P���a��)1gP�g|�(6"O�Us��L#_:�Y2 ��f����"O��qH�x���B/C�K��'"!�D�t
#��2{���LZ!�R�|���AZ���A,�5!�^�V4҈Ȕ�B)�du��+*(!�� 2������u�Fi����.w!��z�N���'ߗo�~�3P��?�!��+m��}��E�g�Vz��Y�S�!���\��(3(:��%XԈR�zl!��$L$		�!���9��B�Q8!��
@B��E�Α	f�h��Ļ+W!��Q�F��ƊL9fW=9p�H�	!��El^\���W?bTr���`ǀ^[!��,�L�s�]=0���#;�!�D��J�tp�Q�ď�a����A�!��N�����J�^v�U#�L�n�џlF�$E �b����V�B3Pzx��cҪ�hO���i�!E��c�C*XF�����!��>8�P�ф,�0.���N�h'���'�����Ą
�F�h�ů5W�e�e�'�!�d��=����4K� .T"��L�q6!�$U'Xꚜ3`��;="���u���x�!�@/Z�쀆����8"ś�z�@��?��|���4'�J�sT��P�
_�����D<�'Z�8#��N� ��-	�b<ܘ�ȓ}�]䂅!�d��U�����	�<	���#o�Eɦ#����Sp�� ���j	fL��ؾ�2`�p-]�DjBP��Rw0%�1�A)(�L�I3*�2xb$���;J�ɡ2�������GV�
�Iu��˟D�?������R4�P�gC�aYU�`��ԟ(F�tIG�--���̊�4jx���E���?����%*���%F8���Sh�3M�����r��B,KN�Y�,�b�> +��؇���VY�2�F
$�U�����?B���9�L��%�]�{L���aZ�b�M����<����32;�E����l�vI���ny��'j��b�	^���f�\x{��$�O�"~���#�~��򪁌_{�$��
�i�<qvė�A4��ab�Dq�c!��c�<���'`��/q�~��2��t�<Ag�W�)�H����'\VQ�S�g�<Y2�1C$"'N&�����c�<1FA|fh$:p���",<��'�]y2�'�B�K��q|��X���*A�Q	���5����re�:Pc��L���{<a`A��I�H�YV+[���9g�N�<�P�]Bn!�p  ;c_�@1jQH�<�FZ%*��݀���9mМ�V�F~�<)1ȝ��x����5hǤ��V�Yv�<� D�԰Z���@ �0"J!��"O��q� ��vt�z�F��Z��=�F��ȟpE��	�.g����5�Q3���҃�]��y+'t��X�!�J�e#�E���y�����k�醦H�����Hٱ�y��^-Q0`M#��J$BFI[����y�ϖK000Abȥ3s�8s	��y��Ǻ��!5�T#$*�aз���yҌ�$`l�BP��!���J6�)�%��g���Lȕ<!���]x��P��V_���U+��0	!��\�nqf鲒�^7RE���J�$y�!��:����g�a3]!�)pq8�'��l�+\�P@j����>��z�'ޞ�k�8`ٺĢ``-] e����'�ў ϓg�v<����w��mۣd>TK�=��e��˓'\/w8���۶7��ԇ�T��)S��5I|��P�.,(���iXN�(�A�v�:q��l�Z��ȓ������(�i��\({P@4��>=��+7K���C#
JZ=�ȓ<���;���a��tufB����ȓ �M�6H�9�h �d�۝9�.؄ȓ��E6Z�J!R��G��4ȄȓYv.�3Fŉ@�:�����	r�q$��	V���(C]�k�L����!"�L�&�"D��eʆ;Re�,P`�
��x*UL"D���*�������@ e�'B$D�l�d�atR1��ìd"��C"D� �*�:��c��*r�@��ì D������im��+�BC�_\(�7�$D�#$�'o�l��C%U�d9��$�$�O�����hb���!�#O�dY�� a�!�@��Bp)�"$WP����_�M!�d�t�2�鷢]�y��B����r�!�dȡ3��a3H���d�ɦC�!�E�gh��]�Nm0��@�:�!���YNq(t,ۗ����*?;5!��uG�bW>_��p��^5/!�ď�vM���a/ T�8 �7=_!��	�b_��1��A��dd� \l�!�ߺ_v�����C�X���=q!��]�[��z1/֧'���h�/�R^!򄒝l0�ĉ��ؒ$�NP�p$Yq+�}��q���p�f�SG��#!N�B4��OZ�D��'􌘛wTFɄ��퐜"�n���'�Z�(�A��,�����I�z���r�'�ax�
C�z7 P$k�>y���PH���y��.���-_�o0�#��%�y�k�1����I:�@�@7�ʋ�y�6��<��ڌ68�5h�K�7�y��ɚ8ؖ�s7���/0�b�G�#�?yI>�������IG��\��	32�x0P'j�-cfC䉟jev����Y.&F��0�\6��C�ɍI�F��&aX�wx�) ��]� B䉉\��i��f@�HB-+�B�	B�.|�I!r(<�:�&�F�xB�	 e��x���/+����,ݤm�NB�	�B��lQ���="��������B�ɋ1Z����?r�D;����B�	�.'�,{�L�5U����ϙZ�2�$��I6>���R3/�!��s��
/<U.B�I�X:*�xSEӎs@��`jԯ2�B�ɖr����aE�;�X��$��B�)� �� ���&  ������Z�T��4��p>�9�k�1�PC�%R�N%���5D��Em?&|	`D\ryء+4D����IN�Bt��3[zi�u�O�=E��$���xI�Q�¹q2��#s�ЛS�!�dԅk(,"�A��$+~�S� A'w�!�Кg^��D�:��I{���
�'���Rj�q���[���YvZP���D8�K� ��g��=U$��FiJ�~r%�I|�����	P(�|�v��.e�#ס��^��B�	:R��t�XQ(E�R�6TLC�I�5i<¥mW��<�[R�ћ6݂C䉀g7�1i����	I6� ���}xTC�	�p��3�G�Y9�abc Դ>�nC�	�r���j��x�ވ9�͵)�T���7b^ze�Ch>	Ñ���ee�L�����*4L��T�Zf��2z[�5�ȓ\*4�j�-��:���f�(P�J�ȓo�*H�C�܂ ����Æ�PAL���x�$ۆ���]r����Jb�,�ȓT�!Iœ�a3|<��IEML�ȓz�T|*Q��� �r4�A�݋a��5�ȓ,n(�v�4D��`��ET �dI�ȓr.0�'�Ή'�������{b���ȓ9r�� В<\�l�POg[T�ȓ�RɈE�^~��[�-�=�n��ȓq	�z�A^���k�)]F�(]�ȓ_?��$d܆S� IG^Id�ȓ�: Xw(�fu�Y*A�6yڽ��Ie�'"�]�`�_fn9�t�G5h��E��'�N8����4�D9�LD#*�V���'�X��W P�Ҹ��V�4HJ
�'�Y#̨~�Pw�G���y���g����E
0� J��y��M�2L��㥡�?��p%���y��6*t���珖n*���߰�y2�^�!<Ȍ�K��e<8Q8����y)MEl����)\��]�դ�y`�U�U�1J0R
Ta_?�yB��CLf�B!�ĆX�\s�H���yb�_�x�4� ��:s�������y«�;�l�x�C!2_���允�yr铭=8�e锨ִ<�����&��y�&(��\��I�;pA؁��8��'az�CT�}�@�8�(��]@�1�-O#�ynHA�a��/D4����6�A2�y��ρy���%)�ҵ�����yr,�nl&���gp�XFh���yR�&h���[g�N�an��ӫ�y
х]���H�χ�f.�i��ʖ�y2(ýu��*��i��i#sdձ��'Paz	)p�P�Ɲe�hL��n
��y"F���Lr `�3a��
QD�y�0�����욵p���8`��:�yr+�2�4��j=d��P��ڣ�y2�!	T����"ѰaO�u�&(B��yroSz�x��!�/"`b�a�mG+�y2GC,N�di��˕�����$H"�y�@&�HAa��HPfh��P#J��y�� 5,/~<q1��PR�Щ�)�(�y��I �<I�P��K]��r��Q��y"�Y��R�׫6L��p���X(�y�Gԫm�rcHҲq��{%F!�y���(}���R�\�J H@-�y
� �-��`��ijz)�eQ�w.��"Op-{����+�P ��)m�H S""O��y�ݫhX�04�����"OZ�20�ےWBj]㖪����'"O�+1,ƞmũYh8 \��"OpYkP�9W����� ��ۅ"OB�K�� �C�9!���)�B�(v"Ol:E�<7�X [&�"����D>LO��P��ރm^�Y���  ��M��"O��q�]��θS+�&Φ��'"O��"�
L��2��5G��4rf"OV� ��i������
)u�� �"O�5ImC<��R�f(8	e"OU���(i�B����9�DQ�U"O�I��l��/a�t�EK��E�Ґ��"O�Q#�LQS�Z`�j����A��'�r>O~�1C�ھ`��9�	޷/�<@H#"O����1o��A�t��m�����"O ��F�R5-��=� � e��#�"O�/Y�(s��9�-��qQ��"O
5Q⧄�$ߠ�� O�<�yQ"OT��RDҦ#��EH��������"O$j�i_�3,�a���6!��щ��'�85���[�"��,�/=49�'r�a�lG�rf2�h�=w:��	�'��t�4M��V���ZSCO**&�PC�'�h㶁��W.Tq�&�r	�8��'uP�	�@�#24�� ǽn(�L��'�rMѥ�*�I�W���T+�'6H4�R�R�y:Z�;)�� ��#� �^�e2��_{�a����+��B�I2!�h#�Ə4P�޸`��k�FB�Ɇ ���fe��j|�sө�?�DB�I�U���R�ڒA.�q�&'֌)q>B�	�-�`$�!C&4�����!
��B䉦B�>�C�!]�>0�H�E�*xI�B�	:��8�ǔ-X.j�ǪF5�C�/ �KE�͆s�D8�!�)[�B�	�����$��"��VB�=z:�B�ɐ_�Zը�� ,F�$ �럂<=�C��>\��]�"��4�#TE�7:#�C䉨#���yc!Z;�`p��ƁY�tC�I�z�2���j@�c}��rG�P3
�
B䉵�����ŘGM\���&�f|���?	���?��'6�~�Y�F  0� �ЙB��4��u�j�QgG~�!���e�4��*��HZvd̸<��W��� ~L�ȓ[����"H���Qyɛ2T�n���C����֐��Ip���K��7rĈ�U�8D�,��ȭ[����fZ M{�(���#D�t�H)1ժBfY�H�n�#�&#���Ov��>�+C�+	y��E��<X�{�� D�\x7"�>`Y |(�$ �G�&h��	*D���DoS6b���;&ȈR� �D(D�4���~��8c���@�r&�%D��[V���Ki�Q��Ņ����D�8D� ��֘L~^!a	�c2����,D��t͖�-p�P�C�jhd�0h.����G����		�䘑��"D�<��1"όUl!�$Ru����$�-s������
b!�ʵm���K5B�Q�Z��w�+Q!�$�mi,$)!��nQ� ��:<!��0I0�@&��08 Ud�<V�!�=�<�L��I�P���P�!�� &J��J�)Bth�(Q�9X�3��'��T6eX�H4\��"�N+
��-���;D��)!����I����5Q/�X�c�8D���A
4`�-X�O��JКq�8D�p�B?]v�ZF2j�P��ѧ"��O���J㮀$R�]�q�Q��H$�+D�Xr!�3�&�c�õ/��p�F�)D���MW�lB�4x��Dh^"Ppv "D�����
#xyF��D;V,Ru�u&>D��0�ֱe�fIXsf��	�Xĸ+)D��g$���,iQ�0u\�I��(D�XPWM�j�FM�a�v_(�ҁ�$D��a�jJ�L�e`� J�H����<��	vBH�#\8��fdӄԤ���I�<Qb�ҵ�7-�h��! %�hO����Xn�0 5��%���C"��]K!�ā'����o͈@�l��F˙�-�!�$��.v��JC�S0�
e�'�]�5!��˹t�m�р#:uhwH�j!�D\�%j(���h̦"@$h�jQ"z8�O���)���Q@nd�2�˰�� h�j�`a"O�Dx ��JP���Õ7�Qi��'��0��IT�|-�R�'`Y��r��<�M�B�Õ��I@T�`����d��b�h��Ť�
Y^�� ��WфĆ��ß��bk֌9;tir��9��IA���ȗ'Tў�>�a��H�s7��Qo�_��<s"�<������(��IX��2oT����O: 0y�"O��Ŭ�!O0x�����1v���"O�y�$'�
�ƥ�DF �t2���F"OᘱD^A�N�Y���9�ȼz"O�D��lY�	�FD��7g�8d�c�'��$�IOH+ѡ�0X�����/ln�X��D{��4CF> 9��*'��p�e�J��hOp��	@�i0��!�f�)4*A�� _�:2�O`��<ђ����}����"OR0�	,QR���D��ȥ	3"O&1AB@Y�^@�A�F
+���@"O­z��խb��x1�ehM���'[�,Si��\�.I�b��x@VB@Ht"�|��'�O�v馭h��P�+~��¢o�x"ą�g�'  U[��Hb����}����r�'KP=3�� ;:���ʶ]'����D ��M�%끕Bj��c�*8�|t:U"O���:*��+�eH�G��%�2"Oܬ��̙�=�Ptb7�� �:hI�"O��j�/6�
�B!
H�dU�ɳ���q>Y"�U��0��1dP&Wǐd ��3D��RQ�R'}�F�!��M���c�`2D����X�eJ��Wɇ�7�~�@P�,D� 0Fm�s�X�u�
;P�p�6D�`K�iL�,�>QkI��)�@�B"�4D� �G��H��[0� K*��3D���BB���0 �0lƻD��q!>D�Ԉ5n�)I4&��!�0�����!D���'�k����5M�! V��<Y�~�&\���ǈg��I��q��y҈�z�\�����9*�X��ҋ�y2B@"��]jN*~�6m�:�yR�8r�j���G�f���h���y������ ����cb)�y���c-���DQ(tV�ac�hH(�hO.�𤒘>���4�,>+*d�ux!�$(�*����ܷD :����)8�!�� 3�i �0CeQTֽ�$"O�}i@�_w�<�Ӆ�w :M�"O.�S'�����Ƅ5��E��"O�Qf��F��MS�����8p"O:D#UN�#;�����D�4b4���@"O6��N7t�����ӡ]��6"OR�I&�-V����/�&dA�"O�S@��O�����8�>-�q"O6=jDG���B�]04pYj"O���BG�	�x�qpb"B�p�"O�c��ۙrch�@p�J@j���"O��x1�s�"h�r��,�ʓ[�LF{��Y$J�𸗃 ����9C	ȴU��D�O(���O����O">Y���hS��(&� �����e�<i!�C
�֖��R�Q��[�C䉛[O�|Kr��m�
�rS�:�C�	<o���-���xIì��<~���Ofp��醤HYҭ�r)&]�`�HӦ7D��bX��ue�/k6\X$n�O���OB�O?9se闕h�Ro�S�tБ��l�	����	��x�	P�'�Ѱ �W�V��&n����'v�R�
�1V��2��'q�v���'��)��#��إI�h�q�l��'"D�F
�c�%��+)R�`�p�'�6���Q�?64(X��E�X��
�'VL���E�=�ba"D�o�l��)Oh�=E�T���S)ĉ+q�;l0���VdW!&fb�'��'er�'4��sW A2g�h]R�lQ���1G�:��0|2r��.=Y�97H�a��9�c�q�<	�_Y�=���G#E��l�FEJm�<)r`��5CBHRa��!-8y��N�<�O�7{��Չ2�U�F�P���R�<�wX�猉\ĺ 2*�w�<A�E�Jc�9���	3����%B�W�<�KN�[��U��1U�<��*�[�<�bhZc��J.	�1[�:娇Y�<�SfX�Oe^! ��XN�܀J�Q�<��ʟ��l���ݽCMzp��_�<��%�p �r�'�<�>�7�t�'�a����=,�&	jd.#t�F�a��O2�=�}�3�H2�A�o�l�l#l�d�<�fO�)[Q)3(u�S�#]f�<!��H+v�T���Me$��3�j�<1�KG�����K7�<�Pb�f�<QR+�� �4���G�;�����e�<!��&]\��B��9Zx�3P�X�<����GV���$&��8��+�^P�<�$m jb�+B4P�-���ҟ����S�Ft�R�b!"�;�A�Cyp8�ȓ2��w�8;V��Qʂ�s
���itfq�E�?7t�$M��X��E�ȓDD�!�͆`���� B:4> m�ȓRSЍ��X1Sq~ #`D �pلȓ1�����䈧vB��j6 W�F����ȓu�.�R�H͍����#�V!x�
̇�b��L���W^U���O�m��L�ȓ$8�Qqn +5uX@�fe�_��A�ȓȪe+��MH�psc�Ԭv�ц�Rh
��e%��	Jn��@�{����ȓjIn`�	P6 �� ��\,Z9��xl���Mݛ|� ؚ^礥�ȓa��H��νfYh����m� ����R�L^��<uq���/F]�-Ro5D���D#��u;���*S���!ڐ/5D�� �D���H�,=�����d��Ä"O�0'L�? 咬�ק��x�� &"Oh����ɳg��'g��N �� �ICyr�'1�������2��`d%��_�R�2�"Or�
c$6GY���CϾ-~pyJ�"O��@'Xኔj�$Y�:� "Of5��ȔP���㊞.���[�"O����.Y(P^p����I�T�p�"OD�A��Ú�p�P%e�����"O���k��Su���`�Ȝ	<�9��'�X1HU�H2N���dDR�O&D�(�P��li0 �@2w!JP��A#D�9�J�]�(1��*OP�c�+ D���fLG�s��R���(�j%�C�<D�h�A��Je�Kd�:_��"�:D�0�G& ـ�3�n�),Qz����9D�p��!@&�j��&v���d�8D���&�!6,y�����o���8��6D�|z�eܽf:�M�b��f����=��0<�!Oy�9P���b��-��!�b�<1�_�^A�8��6�zd*@�9T����i׀2���/MFt\Ly2�?D�T��+v��˰���Drq0D�h!V�J����1G�|����.D���D"|~�-S�gݚ%�l��5h7D�8����hۖ-��d� [`EА�9D�dx橘�H˾𠔥��M�� �u 8D���V���0 ��%f[�<��5D�Dx�L�/N8�k��ڦ5c|�"� D�����ƹf��U�Ø�1t�*ӄ9D���H�Ǝ��i�� l����$D��K�c"Oj���$��h��=D���c'Z�"�⦭ΌeJ0�B�.D���0�z)6�`�͎' ܋3�-D� �U���V�����(7������0D���ڇ1���%�&G
��:0�-D� V�m��F��-y�|S��,D�4��F�'I2f\�p��.㘼�3M-D��0k��H%zH�4��N^`�i"g7D��9SfU⢵���J�s�R��5D������C�0��S!H�K�b�i#�7D��)�%�#/:~P��M[�r� @�w�5D�;��ҋI���J?Z����5D��3.^�gE�8��g$f�42D�\��D��TX1dZ::�H�h�,D�tQuh�3,����Q���I\28�UL5D�$s�䞙I&�A�g%ĨX�l�@s3D���WɎ7{P��sK��l�P�*0D�$`%i�����S��� X90�m-D� ��J7|�f0��
]�TY0Մ0D��(5KH+p�0e�@�Y#Z�"틗c/D�ث4��]_����K�e_�P��!D�T�J�-�N���ʥvT�Q�`2D��Ţe��C�%�@*���b 0D�`�5�R?@$��Fk�:� 苵D+D���7$^�9Ũ�"�'	&>�^]���>D� ʀ��Z!�a
jF�`�@-xO>D�p�L�;X���=lZ½2C:D���U%ˠ7I����MS��jw�7D��2"�*���3#�3�jA�Ê7D���0A��`� G�M���6D�4s���6)��I�Z�؊s!D����JΚlؒD6�t�Q��2D���ؓo��)�RA���j���1D�� D��sE�#p�0p7���Q��y�U"O�p	���9�qaօ9s,Aq'"O�93��-����q�07� �"c"Oآ���hD)�,�5`�.�c�"Od�jTIg�'�Z
px;�Ñ#�y�@Ȫ.Yܵ!��2��5�SD&�ybB" ��G'6.z6])#�2�y�"�H��.�6��3f��yB�J�oS@|��g�J@���y��B{�&��_��tx����y��Mm\�r�J;lm�)Q�y�D��d�5K��e)T��_~j�ȓ?h�H�A� Բ���E�ڨI�ȓ+��<�3'ڴ�(�qe-̫Hr���ZK��@�-G�z��3g
$)Id���_C�H��X1�P� t���[:.m�ȓ1̌17)��4�E��ǋ2`�bX��4�<h�@�L�y���"���؇ȓk|1�cj�Ĭ!�,��	掅�ȓD�t�c��4hX&,i��v��ȓX�$ô�O�'�"� �쀲Dך��ȓ��0�É��J�%)U�;aP��ȓE\�m[�k"�MP���MZ�E�ȓ+F��)�#�"�k���f�:|��V7l�u�خOg�-�0�-�t��5��4	R$8RY�G�Υ;�����Y���ǋ]3� ��NN�@9衆ȓ�Бv� p��5��a��V�%�ȓd��)�Q��&��h-�}ԅ�:5h���K�Yܐ����N��ͅ�6�h��]4�=x_c~Esw"Oᱡ̅�B��iqV`�iOH)s#"O����L�b9����8B\�"O�T��l�T���&/]�g'���q"O\(����V��d�V�W�Ƶy�"O�`��BO���1wo^=z�����"O,-��&�+6�*�@\�3֖�CA"O܌�#�ތER��1O�I�bL�F"O8!c�	�!���s� � ��%y�"O�M��)�o�|���\����#"O��Q�4hx��	�$�A�"Oz4J#kj��͠#�B�%�q��"O�y�_5vbX�SIN,(�@���"O,��b���Dn (�P�ۤ�~hBp"O���v�4�R�Ӆ�z��pr�"Or�0
X��'� �Μ�"O�yS��7 ��@���3F�\!`f"Oh���9�$q�[�l!�C"O���%�C���;A��'݄���"OT���f7Aw�M��B�g��b�"Oތ���^ .��|��	�w�P��$"O��{7c�x&B�c
�	>�P"O.p�t@�M�Řņ��4�<��"Ol0�S!�����r��
T�4"O@S�qO�����[��E��"OL��w,_�#�F���	x��B"OZ��!�S+&e	lˎE��`��"O�I+�B��y�EY�j�,!L�`"Or�ر�ΰ<z^Iŧˠ8{
�B"O(�ɦ��-:D�:���(H�t!�"O��iF-ŉp�da��g_����"O�l�e�]�Sq��+cG8%T�d"O������/!0$�G�^9���C"Or���'D�3��r%��=�D@b"O� ��22e�!V��Q�R5}J��"O��r�n̽A]�M�&�}X���g"O�xC*.�$�x��&[Tz9#�"OXp� K��+E �Jç� �"O,Bw���{^|`�רQ�6d�!�""Oʕ2T(W63�q��$��3/X�0"Od��!V�Z�Z�Edr��"ORq(@��w��m��DQ�5���9C"OT�Y�5���8�� ��a�"O�D��q&��Պ�GkJ]*"O�A�a �B�>�TC8�i��"O<��� P!T�\H�EB��NӴ��"O�A�C�Z�N���Z�ȵb"�A3"O�T�5�S�H4���C*	@��G"Oi
�j[���9CQ���s�j]��"O���qh�����(6�I�"O.�;d��!~n��
`.	�o��<G"O�Ƀ�E�o� �9��G=!��$��"OT�Rk��P.�У{�RVp�<9P�ӷ1%�;��޵}�Mi�%p�<��l�:8�x�;+�}��Q��T�<q2/��]Tj5 �"ϯ%X�)�N�<�3�ǚ*�=P�(m�>�A�kFH�<��e�9���`�K�f�2�o�M�<���.R�uJ𬟝!hl�j�~�<��?��T0�͘i�|����e�<A��7vg���r�W�yV9CEn	]�<ɥ��Tf�A��^�=���"A
�M�<�����@ƃӘ/,ѱ��G�<)BEMQ\�y2�-"j��!!IG�<�g���C��K�HM7q(�(���E�<Q�*-	)�D)3 �>m:2ؐ��El�<ya�**"ʙ	C��X���<ɗȼl :���g$����hc�<��J%|W\9��Y�:�㔃_[�<y�BR�S�9���B�:hKQ��[�<q�gT4~4 P
�ˇ�}��ف��M�<��D�5D� d"�F�X��SA�<!���5\��"A	�Qv��g�|�<Y�/ʆT�p�K���,��u#1D@�<	G.Ŧ
ά(
���H�.ia�<Y#� 3���r�V� �[+g��[�<y�c9,��ͨ�LG4�R�����[�<i�i̩5R So��&��Tx!B��<I��� ���	�U�rtDig�<�go8y^lIɷ��,w ����H�<A5`�C6~h��#�$+WJ�#K�I�<��.�qP�iw!�	#����%�Zl�<Y%+U�@3*x�`ɱ'�@�<����� �PJ�	��p��q��Mu�<�7HF�R-R�p������V�<1/��*�Ұs�C�n�<=�eZmy���v��J>��	=q����G/�<e����<�S�G���$�j�cۜ�S�(f�����H�8�I�bC x3���t�G���	��p>�Co��A7�� ���2T� �Ơ�R�d.�S��	�>ᷩ!/���񌅓ښ܈�-N�<i5G�, �"E��zed�qV�#Ⓚ�\��%�.��x3� 
��`W"O��bEe[.�Qj�+��L�P"O�E2`�,U��%���Q:H"D[`"O�Dӊ��9�� )wF� "O|�g��K��D�Pb+�u�'�	_8�(ӱ�͸ �l�:T�K�`��;�7D�� �q��k�U;w��(��u��iQў�E���A�a���Ĺ"=��AD�����>���<I���Dz[t���nJlB#c�F�<�rG��9q8!�CC
�#&h�� ����P�=a�Û����'S��	��:@�'*
MBلȓN�l��/֧

v���]AJu�d�'��O��|?L<i��yi<���D6�v�#3K_�<e'�h&�1�&���u˂��~�<��!���zg �,%����#φ}�<�%ɜP�F��C`']!�x����t?���'$��t ����K$�X#V`<	��(`��� ��de��#��"\}��8�>��G�Q�� �to�:zP)Fz�'(����[�g<:��ա24�	8�'gdq���Z ev�W��7�%��4��$1�Op�p��0t��h۱(?Pz5�|�|��'�.���fS��&lC$��Ĉ���1<Or�bpG ��>9
1���cE��y�On4׭�	��3�¬Bv��H$ˏ��>��'�	J1K8d��b+��SLD9�S��Py�F�o��U�P��*YxZeX`��\�<�N\�~�JC�޺Q���{5�X�<!��/��e��
N�Nj�X1�i["fў"~�I�j����k�A��f^�a8J���>��@���.����f	rf���0=	N����<^����T�r�
R�7�O�O�Đ%�C3�l���	�={N�;d�I|���i�*!.��`Β#$��Y�&$Ä1�!�d٪>I���Ćl��cG�ў<��ӭa�̫���L�@�õX }�,C䉖!�05�b��2"��(�Ⴠ�UIC�	%J�����hN�\�".˱3��b�L��	��![Q	rn��:�Ȭz��B�ɹ|��+��� ��{������O���?�L~�+�^@���^�fyp�qt ��]�(m���t�O���F�ΏHQ"�#��ۯD�p|��{"����<іƑ��:	>R%P)h�&t����?��A�j��\�AH9	:n��q��x�&R�{6�g�Pe��1h'O���yB-��l�F"§Hk��v�Y��y���
����CE^�U�����T"�(O"�'���d'P|�9QD Y�BdR53} !�d\ql�+�*
6�zQ�7���!�D�?pj���D�%!ފ�#�,I�n�!��?dQɃ���!H�Ȳ
<$/!�D����ꧨ�c(�!�^2OA!�DS�K�$d-�M�y @W/q9��x��8�PJ,+>��6mB�~�(MC";LO��O���Ϭ4��	�Ko���U�2�!���:�L+��D�Mm©U�L�9���3���(%��B��^Eʀ%WoB�8e"ON���O�mNq$��4��+�U�D��'��}h��h���	b�@#�4����N�J��\P���m8",#g��`�V
O����X�J�pT#�*|c�����'�������(P�@c�ġU��@�/1D���*��Q�b'B�My��i�L1D��P4	�wD�݊�C�,/ܼ�C�/D����'Vg (]Y��E2e&���V�,D�x�V!E�H ��A�4���&D� �B�ƨ4�D��K�9H��Ѫ%D���Kр/iv	#ݶj4QY8D���SjG8'H����/ip.=��N4D��	�ǝ(������A�X��(p�L2D�� ����^�`]�v`�<EZ�@��"O��c��I�G��0ȳ��pH�� "O�<�4Ξ�K'4Q�#��]H�)W"Or�i���v��Yu Ǜ	�cg"OFcE!Z=D��ѪQ��=@����'��	V��R�^N�<p�ʚ/��">����,@�ΩÓ�F�6*���� 1%!򤖶y����j�� �З��I�5�S�OJ�U�!+Y	t8\X�' WX��'���4�۳(4bIx6�
x&����'��d�,/KP �5`C0t
�(�'f��k��^E��#�I�4�]���D9�S��I?S�53a"�;\�&]@�㉤�ynI+S� ڳ���jq�a(c!�9���p>!��� /��ZQ�(gT,hǇ1�D5�S�D��O����<�-�fN�I ��8b"OT�2���(Ue�/z8 ��x��$IJ�'�0y3��	��q��߄5u(�')��`�&���P�I+l~��ˌ�;�	V�4MQ�g-,��愙��T�v���yb�6_(�)�����А�H�?�y򋈝f��h �K���ݨe��1�~r�|r[���ʧ#�t!�枹v�0[�͆�npB�ÌK��������#7ޅS&EY�_�`��FLE�p��L��?�"5��"�L��&S�[�� 5Fw��B�	6w�JL
7N��J�����l�=���q\L�q%˞Vg��'ʛ0�ў,G�T�i%��s���a0b�:�뇯I��c�'�4݁cm^��m]`�%C#>]<���2�S��"�# GTQ{E�" ���؃J��y��Y�R��v��%a���� +�5I�v�=qF�i�����C*Q��@��XӬ�V�<I�L�dS@ SUgR*�2]Pր�m�<�ざ)M�<,vL�����a�<����9�4���$8��3.QX�<Y�^7f�였"���	�2�i�<�!C/]�*R�J���H�`}�<)S��>Q� �B�����u@2Hֻ�hO?�I?	>��g*r/�|r1�C�	35�� P�Ž.g�@��^+Pp��P����d�����eN�3}�ak�(��0|��E8I�c�FH�p�F�H�'=�xr�4>�$�JF��5gjmYN��yr)żo� �V�ʥ����A��(O���$�M
,h!�,L2=�7�ޙ3�!�D�>a��hh���9����C-P�!�}���h�Έ-Ҟ��˳z�ay��	,k�A�HZ�PeK���9��"?�q�?�'�X,1&�@�9o�����ڞg�l��3�t%�W��M8��R�;���'��'U�?��WN	L�8����ǻ<�|{&�"D���-X�I�.�� F�[`h�
�%D��� �"���N� Vu[5k%D���t!<;�0g�׺r.�IG�6D��Zud�,gd��k�?n��$�*D�(�ʟ�����)�4d�v�z�C)D�@xOT�\���GK�c�R`j�m%D��4ł�R��`Cg��CNPz�-)D������S�|��ՃS$��ׄ,D�H�bA�f�T@`өT�<(��+D��gO�	�a1�㍣��q�6-D����!~��3��Ԯp�a5D��P��ŉR;�b�C@���%�5D�����gX���6"č'��QCH?D�� .�A�狒d�| �D!ɌP]\�"O��j��%

�u�� �@?rq�f"ODp�M�/"��w�H(78�@�"O�x���58�n�IE�ۄ(0� d"Oޘ C��P��Qǁ5;�U��"O:M�u��\�Psd�E�jH
E�f"O�D*��J5AT�]�׮�f@�q�"O��r�)Ƕe�y@Ӯ�,c6���7"O�\"Trf塡���1!J(J�"O�`�2��0�Y�P,�+T����"O�M�c���*
�u�$�ƈ��"Ofp�fj��D�fa�IH����[!"OF�ҷ�ē�pxPM��Iz���a"O���_9�"��#H8+�.r�BC�<!T�W��|�;`�8_��Щ���t�<)gE]�p��QׁU�t�h�7��l�<i���#Fʨ���'d����o�<�t���f��q��%I:\��)�k�<���34=�� �^�Z���i�<��\ ?�j�8W��:
��Б(�e�<���D%9�|��0E+�� �$[b�<�ԀB7Ɛ3C��&gJ��#a�Ra�<i��޲~T����ޥ0�\�3GOw�<���Q�j���d�D�L����F	p�C�ԋ��3O" ��F X�KyP��<��%�on��r���Ҩ3r�RG�<�"ڮT�Dd�O�B�
���g�H�<���ԫ���c�R�D�Qe�Nm�<��/(<買�*vf��7�j�<�qW=�NpR�h�!u� dV�e�<y���+
�l��-��=o��І�Ay�<Y��٭JA�Xx��4H `2'�^�<�W��mZfL�`ԬH���#�MM�<�A��h�������{��-�AK|�<I�F��&�t�%#�5'T�4k�JQ�<��G\%2[J��S$�6��!�$h�z�<�pSr����R��4��A�l�<	�+ѶtU^12��ߋV�(����Ov�<Aԩ�pv��R��A��b�����q�<���J���\R�M'<:`y�@,�h�<1���G�2X�6���9�D�sq/�i�<)q��d>�M���4X��K��M�<!U�'>Ѩ����ȖAEhȥh�I�<9t�Y]vԑ��_	V �+�H�<A�m��
E��&I�:i�1�eB@�<9ń_4v`�U-��;��[��@�<� R5B6=���1,�j	p�A�<q���U9��u��h^�0� {�<	4��# NPQr�,d�� �l�<1��&<""�E{!ŏ
3��-�ȓ!m,+U��yW$����Y-8�؆ȓ[��iI�/X�O�M�Ŋ��!z ��ȓZ�&���b�v�Jy��ʚ�U����ȓ17B����ȟ��Ia�F�!���ȓ,Φhx2A�'�%JBOQu^؅ȓ88<K���<�)a����ȓ?�Z(�G�����!���]TX9�ȓ?WXa�)T�#���&�LN@|P�ȓ B�L@#gͣ5�=[$��I�6�ȓMc�K�&(1�j@�#���P���u��+��H��ԑ{������6e8�9/l�9!���3.�(ąȓDo�� o�'�i�C�I���ȓa�ڙ��A�w,hDP� �#�܉�ȓ5�5+�M�5`ʈӱ 1bhh��S�? ���iE�;g@�a�m�,= L� �H�p+1��� !���1%�*o��H��G�[��B䉏��U3���"ؠk'ł�,�찠���P^,�O��}��a����*N)S������	[��Ą�3T�A+;�JAz�$�`���l�q$|�1���J��{��I%od&x�!o��D�"�;�%U��=)��tl��:�!�O\��ri�
|
)��|b��U"O 0J��φ����Fŏed�92��٘8M�dX0H�/�h��A�gj�
�)��
ϔz�\$�1"Ojћ����[�b  �ި$� �����>\^�e�U�&}��?�g}B�:,fb4��.��=�p����(�y�FH^������.����Q����M��+0&@�e2|O�|�3��'��X�D_�!$|qF�'����E$D� �b����Љ�KD�X�dq5C@b_�C�ɠa��£m�|�@҅�@�++���7�0@�.�G�D�J�V�.��k2��'H��y�!V� "�pq��e��x�0�Y�y�m�5�* �K�B�>���ߛ��'>�$��&Qv�O�ވ��͕W�n��HN�.h���
�'C����HʾzgP
se���b�J���O��:��Y�|q�K�l���a�mN�(�lp!"#D��;ׅU�8w�<�e*9�2�I�&�rXT�G��Z��|�%ˡ-�FE�T+L�-K�b�ć��0=�Uf zj������,�8_�����˅��c�<D�ԫ��l�4�4ˉ<:�E�S�=�	�8�uɓ�<8+Q?ycC�ނT�(U�%L�`�J��=D�ۅ��9��hhpgF
8P�(f�T3ZD|��a�>�,k�����/dFD3�j:WK
�JE�S�%�!���z�zTc�G�1N!��.�8E��-F6p�~��1�3!��O�.�y>p��i<l��<���8Z�޴x�GI���r�'�ٺ��K�'�Р Q�ÏL����J�.��@��:j]� "ػdH��=!l݌0'�D�5I&>(��I���0s�L�?�0��������G'��,F~���`6�	
.Aj�� W�aK�>)A�@T�H@���艒6���
�A�\XU�td����0As��Oj��Ǫ0IHS�	�'t	H5�҆;��5�R���;�X�g*�cZE��ڢ(G��<��OA���Co%}b��7hBd`Ã�7	���$��,�vć5;4HA��K�uC��Aq�A�iAlp�フ5��O�8`��fC� a�K^�pW*��$F�$RVd�g��IY��xY��ș'�v��nK�z��0$���-pQ���"&*���NƋE�8�iN���`HJ�BR���'H\X��K�����5���a%G.�Z5�ЬB�iMT]z��h����,��.6�(Lc&-Al�<^��B��6؀��Զ�upb	�83D$�j�h��8�K��ğ/O��pR�'d�Tҥ�QF�% 4�����]�T��Y��n�'}���Y��J�X��u+Ŏ\��`�J�'<����ڟ.�B�F?[Z����$�0�@�G�z1�í-M��O�2ǚ�۸��S($2P��>^�n�
@A��J���Gݒ[��Ė�����_r�%��!
<[�|�Z���\��`�!L��u�W�R%8���II�u���`B�q$��?K��]j2�ć�0�� l<�Ð@�CW�ejrї.�� j2������0=Q�bǶ[�T��"�,{�#1+I�b@�@�>,J��2G����D��
�]�
@ã��.y�Ak��-�)���6eX����j���*�U�ay��ˀr:��&��)v�ߢhک�喾Y"5�`�� [s/Ё7�\�2+_
,�����26��SZ�\x�t$��y�`��y�nQ�,p��0F���i^���H,�)����"
��!�>5���E])%ђ��hAK��ӑ�ߝB[܍�mȨ:���d�=>���@�)+�=��n�ֵ��C�~�N�T`�q���M�s�E�"vnu�R9P��w:�"�ժlba�ܹk����&�#)eR���F�5������Y[�uH3/��p@}(��_�,��y��1��*ψp�"��A��4��&_����p�(��Iͧ
@m�t���1g���PH)ι�ȓn�j�R�bR5����$ߍs��<����,Q)JE	%�M�F��P��a�S�Z����.�>y%	_�g@\��sG�"K�6L���[���ae�߹&T���g�=^_�A���$-fxqraT8w��ەE�yl�h�%��4x�i�Oh��+s�ޤz��觋&�i8�aBO���1ZT��u����i�uӱ'�~��*�*"�T��fj1�O����O3K,��� �Q�P����\:� #�ЙR���A�t�y&	ä@��$?%*��T�m�I�٨R�L!F�#D���d�2]� H9��	J���� �^�Os1˵N�#[J���-��	��c>���.?�d#*\u�a�Q�('�b��U��P(<�D��vht��ԈV9b�^���)N�nZuq��G�I�n�3��5�O�ez��#Xh��&��1h,���'Yl�,��&�r}
� a�ӳ&�d�	��6V���B�O�=+��0>Y��6��A6�٤oY��v�,I�C;扷-i�#���w���2H���r�Ai���5D�p
pb¯&��"�G_<D��i*3�3�I:L`
`�d ��^�>�" DJ��P���+�h���#D��X�J�w�)-��P�6��]�z4	,9Ҝh�O��}�M|��:4+:�����ț�<켼��	�"������C���h�H'_��xS�"-��O�@�e
w؞8SA��;!ℨ�p�+-�4d�� �I4]
�
�E]~R/Um�0
5`ʺ��D�(�F�B2OӾ "ɫ�@��<�sLX�Y��)F��?�@�Z4=��{�N]y"��l��,Cf��V�i��@3U���կ�f(h�L�8�!�d,hD��"T
H���P�>1��F���bU��ڤ��̃�Ę�-��$i�ᚌN�ȹv�FN��z��~����'S'b��I߫|�|Ԛb�K�&�jh��P��?�Wo�,*���C�&lO4�PG	!а�@d(��cu�pR���09�@I!ĻX�L�l���1�Bɱ��b�x�(P���G��%���"1�B�I%��H�	/#v�;B��r��}2)�r���
�C#p�g	����@�I�/"t���9H��!VYZ$s#לOH�:@��&ta|R�Հ� ���'f$݉v"�:W
ݛ2�� �3�Ҟn%b�ɳ�Q�,�A!pK�.3f ͹�b��?_c���!�(y�֘�g�͸
*����/�	�V���ɡ�P���ԚrZ((�-��>�i���(~�A�e�L0����L�W�d��BR2`�$�'��ы�O�_q`��!)_i99��j��@�UGf���cђ<����1�U�^ul�ȁi�o6���|��YW� '� ����C2l?�����*D����N+�\mcm��A��I�"��L�n��B�U�5��0t���B%��T��)�D]bÍ������w0��c��L�@$Թr�M"��'FH�{��''Z�l�Hcb$I��N�D�j�c��?� ��Ħ��C�� 4��28�ȣ��?-���`���͉�	AY"@����#7����?i���:#�C��<��M�V���,N�P�h�`�U+$t�0Fl4U�q2G	@'H�"b���=q���	+p�(�J��a8�� z\��V� ��	���!B
�\)���,����GG���2�<��6��-T�&|�f�E�<Y��Ю+�l�I�.MA(�1�BG?i&#U)K�|i*")O��60k��g0V��D�&����V��qa��&|���"r���s:Ĭ��I�bh��a&�3֦� pG�s� .
<�{ulu��ҁrC��'�Zs��P��G�(:�:@�7X�X�s�l0ʓ�@��'�Q��!)E&�Z��4b�"'�u��Sf&x�e�q�<%%��H���0�)P�e\R�(2�6D���7� i#�Ч�řZ�XPie�5D�L��i�*Ұ����S���5g3D���'.��Ua:	RIè�@���2D�(
Ң@�8�P@��)5NdٗI*D��$��7$8<�s�]�4����%�O\��(�H��l�^�aؒ�u��
�'�ڵ�BB�:mٰ�ςB������/b<��I+S���A,�.�>�醤ڔr�C�I<+�py���:*X���Y�RZ����<�A�򍍍y��{>��������4Y��(��D��Ҍ~�[�cZ��S�&a� 
 �˙
�hx�O�&5x	�Am?}��3I`4�R"Z~��1�J�6�$��#��Z�=3׌=ʓr��!�A�*�	9d��x��ST����F#^��0�;�P2V�(�h�OأeA�[5D-��"�[D�G�A >Q���䀟.B�ʁ��������ee�9I}^��&�ǻ@EF|��"OvBB!�T��y����7G>Ax��Oڭ�	�ک)J��s�aZ$1��`�S-,,� ��o�z�L����'M�q�o��<)p�#-(%+4c͹�D�����C�$ƛp1Z�8�)���0<��'����"#�=R��)�#K�Q�'8�[��d�!�^ �D
�s����D�-�n��e��.���3�'�XQP3���ݣ�[<�dx����C�"����>�Ӛ
��z�jM%p�^�Aw!�87D:B��!'��b-ܷr$:���A�@��p�Ι���?�)ʧ9��A�Ғ"*E���*��9D�c��>6 ̓ �`gN4���7D��rTǘ4vE�P��/_;�6`y�I3D����HO���-#+ݢ\e�T�q;D�� 
S)��
�B�L�2)z ��"O�A��F�q�� ���3)"(�"O̠1c I�DO:l�� -x�v�Y�"O��  ��:u�񯃂i��=�"O
�6NF)y:Ĩ{�#I?5b�h3"O�@��D��v�E g �z i"O�}���?.�V��!+���"O$5K�e�[Jt0���o�9�3"O�0[�IDD�h��#.&����"O�\���WX��i�F�H1���{�"OҜyv �5R�RYu.�{�ZQ��"O i�C�n~0,�n�)b��͸�"O�dB�Ɋ"�lݡ��8%U@�"O���$'A��/aCf���"O"�q�NUH�x��c�۲h�F`8�"O��$"�R��m��m׫=��I�"O��qB�#<�LdK�f�>v���"O �A�"�~�c]����"O�� oO+J��ґ�D&QӘ5�C"O��Yw�5O�X����;n�$ha�"O0�qdԺo]�u�0�v��"O�Yʴ�N�m��i!g�;�X�A@"O�` S��I��8���N�%��ź�"O0�+�����;�!@P� IE"O��sG&=��[�S�V�@|)�"O \Y�#�=OX�Iģ�cߢ��"O�9#���y���Q�a����"O�� u�/���vb��v���q�"OZ��ƛ�LVFQ��H)�*�B"O\�����8:�B���� O`>��3"O�u��B�~�td+@-PW��I�"O�5�B�Ç3�>�� lH�(]p�Q"O(� �+R%heB�%��9c����"On�aF�K�Pj@x�TJ�3�lͣ�"O���l�=>�у�����"OX�ۣ��"��Ā��B�z�%"O0��*b�`��<�C"O�Qr�e?F�Ddq�"�����j�"O��ǣV�/��G��f�4@��"O ,Ȁ�C?{���S�\.o�"�"O�16#dY��E��;��qB�"O�t!T@Z�m�8!{�g�kQf��"O�z��!IzZp ���_���u"O(]���ޣT��B��_5mE@@#�"O. y��Q���5��cU"OnX$D�~��XB���]g2�ڰ"O�mDC#%�H�hGLȗE����"O�ē@-�0X���& �<:ѐhЦ"O�`��#Gk�y"u&͖Rd��p"O��0D�\��pQq�K�!J�p�'�,]y�M��g��AB��(0�v�j	�'d2՘�H��ؒҳ:Q���'��=i�n�)Z�°�Ր6f��'�V�c��2MƖ�i@K1]���{�'f�����`�d��d��gͲ�
�'����%��>��ᛓ�\�H�\	�''r��50C<iz�
��FV��;�'BV�Ӈ� 3���b���h���
�'��y�G�T�*��!�P�Ģe��9`�'� ��A�8K��؀G��P�:�'j�Չ�A�I�l��Gh���`��'��X�r�Q4>�ы�f��A3��)�''8hqA%ßj�D�1��˙���)�'p������h$k'�������
��� J����_K���QM�m��(+�"O������%5И�1K�%'��X�"O*Y;�CÐh?����������"O��U�&)L
0��p���"OA�nцv��\�bZ�(���d���>����!P�%M$(�6�ވb�B�	�?��������R�ޭ]Z�����H,r)4�O��}�WF̓���>�Vx�6��m2|p��/}�Y(�BŔ~��*�K@����m�	@��b��"XG�{<	0�b6b�Ry��ZG�����=� j�1]�v�����O��Q�(-�VQ�BH�|k�5�W"Ohr#�#�T]�EGH�f��{��$�,=����L5�h�X���iN2m�TX0 �N��kU"ON��a�1� { iE����d�ş1��I3�(}b)$�g}�̆/kި�vh�!�����F԰�yb�!.tJ�Ќ̚y���M;��AD�J=�a�9|O�ܛ�HVP�4� SH��v���g�'f U��N�"R��(�ɮ	� 9��!V��a@�Y>��B�I�o��Ā���+Mʨ��w�⟐�.B۴�E��c;"���8p)S� \N��DHT#�yb���C���P�1Q<�D3�B��y�H�%p��tDo؃z�AT����'zݰD�Hb�Of@��ޢ������PѠ
�'�.��T�P$~�W�ʅg�x�5NH�ȒOpٍ�Y�(��.�!����A�����23B D��чI�B�,�T��5~j�!��^x��
:@�|r��=O*~M���t�͙5��0=�DW8d���*2��t���4IΎ]��+]�Y;6�:D�`�b��-et����"fUyJ6手%re�
ׇ.�Q?]"s(@�*� P�v
	)Gp�uY`k4D��eO�1v�����JzX,K��ճX��08C�>I�]i�����Zm��	�-�dMZ)I�n[&8�!���f��YJ�	ʙ;P�c�M:,��P�I��b���i���#l�i�fh2Om~�SG��?/�x������?�����'�qY�c�O�'�vТAM��:�����.9�qxG��'>(X6)C:Z�AExR�*Xx`ˠ.5N�,R>q�����O�\궈e����6cקb�~���y��g�f���I@e�O�U��*ɃM�n�ơQ��h1#oЄn��$�dmX���0�M��
)��ټ�q��>�ċA#�/M"�����,͌ȳA-}���6���I%d(�	����Z"m�P��6\� U`S�v��5`S�	pyӅJ�,�9'�A���' y�KSwL����ǶWq���A�]�:�A��o�'>R�6�Ͻ'�$x����)��*G���
��ѵ&�<�V��bO��w����@ �X�� 03��Ͷ��dK�k˼!��?��L0wD�-gU�O���E,�ݎEC��1~�}��nI�]Ĥx9Xw^�4Zq���D���A�$�X�H�}"Ɇ;W&�|E�4FH��p��0N�'30��2A�.$f��zю<�Q
S��-!~�2���-�t�>)�;B�%)uO��yQ�4E`�,c�BB�	�+x���ˑ���k�&ޱw�&��Ҁ���$)P�Cc�k�-�|��`�J���'�R�wgM���UCGg�|2�l�ߓtv��W�H7�\�+�K<da4.�*�DU!�I�}�P�+��"g���a{B F�BN�z�f
�i�xx���O�4P�- �H�2�Z��`�@Ѡ��
�I����xqхԟ�rH����4+!��� {lV��P�-�����Ǣ\s���&E�
W*t�"(Q�9�~(��M zmQ>���R���Bc��:Pw�y���6y!�dX�0��A���2Z�H):�.X	U
�m�O��b�@ܲ���qO�:�:DǄ�
�O�:^6�q���'��jǮ�;zB�O1u�@���'_�R9�ӇDo؟#��U�!��9s��&g�:��4�W���gM����­�g��!2�z#A��'�)�g"O]���F�,�|����C�2'��q%Y���k�	iހ>E��m�VO���Ee��}��]����y"�+ڸ��J��l���+�d�'34���@�S �ϸ'>*�IG��	8 Qp�$�0(?�%"��< �qs^*,O�-�ǁ� x�rd�ۊ���K��?���d�Xa�%�+yH���'� �BH-�X�'��R�f^�/B`(�k� iQ�9D�� ��*�E��^���3��B	-��	��>�G��X��?q��e�h�d��T��/ ��  $%D��!��JN��@J�7���B��$D��x3��nT�P"�m� /��zs�&D�Q��l�q�v�?;0��&,��dSG̓��a|��ؠ�A&���,��.ר�0>�FIL.r�N��8��� �L
_��Ȱ�%/�J���{>d�0�C�G���'�"�e�?Y��#�rИA'ҧ{N�Mr���j�r�ZW��X��ȓ�f��U�0|��0bݞ�nIJ�kG�ZO��g�>����O ���ߤQ(x�JR�!y\Hq�'$4$���t}�i\�,��d���R�[ �a�B���?ٲ�(4̓U�:lO�a@V�A%*���
խAK
y���DP�@��<�g $?a�
V�#�$ui��`ݹH��A�mM����F'Y>� �/#D���%I��	s�ĐX��A�^�I�$��<q!�'��;	2�針�yW��d<̲ KI?Rq���R�y�x�\Eh��)'����`J%h����Մ@Rƈb*O,����)RY	�}B�����O�(��ċ0�p=AVA�L�j,�r��-�Mk�IpZYb�@ʟ]��H�m�����PgU�e
���u�'Ab���]�y����ڝȍ{�JH>z�P�ZbK\�zG�	.UC��C7b�?��� ��`�Bݑr���ವ�j7D���#k��~�P�%m%p��D�;����͐��?�vB�L���C��~�@%ȹ?q�?�h��ï��N�lL��莌l�>9#�'v`t��i�	�r�̖
w���c����0�s�Qq��\�Pg[>;�ly
��
�=FU8w�̗	�Ń[��O�����D
FL���Phh�� �k�q�'�S	�?�Ņ��&�0�&\4}q4�����N4�<чK�.T4D@`θ�b}��c�{���RۓA��-����H�vL�1?�m:$�] Tq�@a00O��3a��D��B�
�`��ʲ8�y2d��b�e�]�b��ӓ�N�^�~�[g"O걸hJ�~�mk� gc]��*�=�q���<h��TC�&���э�n#��v�A���w�F��2�2yG��x6��j��H��'�м��ȉ:\L�o�� ��D`4�ˉa��%i%�Q"3:R�k@J�A-��X��X�U61
��?9:��Er�G5(%�@�Y�f=
�����#MQz �?i����rxrB��<�@G'+: �ai�<�Ly�sFů/���ba�`��+�O��>kL̚2�Q?��=ѷ-��y��Y��m���yZ���>�� �	�k����y�s��d�iۀ�D v��s��_�c��^���'%ѝr4�x���F�<a�ED�D���(��;`)bV��B?ᶇ�k���a��2B,�B�U�oy\��&h���*l#t7m�� ��r ɇW��I�L4��¨@��D��\�>9�ݰ6�(c:(x���Z�¡��#�My�������ɜO��;�	�%�����!܀H�H�<���D�N�"~J�� �c>����/<iT����\�d

8+�#I��	�"m|�q�+U���5�ʎf?^B䉰-��=���MK�@���3�*B�Iu�<�QwƠ����2Ʌie:B�ɇI\~�*��D MUV��䃝V�C�	�	h���/@a����8dP�C�	�~{��:�Љ>>ѹ��^�4�p��$��y��!2H�7V,�A�#E-f��z�fI���xb �� 8� K�"��p
���O&�XW���[8�>ݸ��V�72�{#;2xl�P�%D���Go^��;U�T�ND�������׬(yg��f�>E�4�@/U-�Z7fR4L��F �y��U*
.�*�۟QZ���2"���=��CUe�)F�axl"!��	���_�N�Ā�h��p?	 �ײ����2�ݡ��HŊU#u.rPQA��/�C�	.g���2CA��r4p����Z혢>aVLʼ/<,bpj'擢:UR���(�KdYՆ�W$�C�I*s
�r5�2V�c�e�b]��	+C����h޲/��S�O%��;��ܹI�P5��@�	�:̈́�Hq4�"FNW� ��yǈ�;��x�O&�sΐ	r�q�
�HV�����2X�&)�Q���$H�4��I�ƈx�JO�6/�����&=�	�C&�C��)�@��E�+��A�Ęx� ����O��Y� ��0��>1���#+�8�kج8�My�l"D��P�ܙ;�h�V�D���DK3o�<9���4➢|� `�@�EI�M
���2��joL�B�"On���&0zT�8�)*+�q�"O~�j�ރ.�8 �0��O���Y�"O���a@ݬpz�y"��Y�%p!"O�-���1_ʕȲi�HI�` "O�1@��]�T��iD=un؀�"O��知&�B�+2���LG�((�"O���w%R�r]0���ۄS醰�"O�ѣ(��3e�y6�����"Ona�`��f�\9ԧ��h�As"O�	��
[P��7��(�r�6"Ox��
3�(��d_"�2���"OR�+2�в."�X1G"�L8f��w"O�I#�]�=�8c5KB3A.X��"O�Pg����Ѡ�+݄(�d��"O��$�X�~0��ϓ�9�t9�"Op@���+��"R��#�T;"O	�� rA��+�O�ru4,[�"O� #C�K�M����1+U$`o���'�y����l�h�����**ze��'������>Z�A�L�2 ���'edlp#'Ѩ" �X��b�$����'�|�ؗHǺ�r�������'�<h��ߕg@"4jr�B�ﴼ �''y+c۽Qa���|[z,R
�'{,1' F�}����o6c��x	�'pU���*�����C�P����	�'�b�� �>�����,G�J����	�'�d�rU�I�G��xH�a��T�X�:	�'p�]�j��j��T�qE�{*���'`*����	T��A�W(֨p�����'|�r'�#� ��fZ�>vh���yR��9yv���!F�'x|�Ir�Ë��'�|]����!d�X!Эܟ��B�'6�@���
�L1W�OO2xy�'�:M�ՅT%��t��G�{|�
�'�r�p��]q�(V%\�!(  �L���'B�*ç��q��-N@�����s<���qm����DV�z[e����0|JGA�>z]���OԐ7x�U��E2t�$��o�F	q��%{�X ��ӷi��i��I�`�$�P�T��74 L�5a��`���
w>y㇩Gl���BBN�8���jϧ0|�r�f�(&p�?O��𩉑R�J0卍�pF��U	�|�!����S����'at@��'K�B�kU#Źq>�1JB��,⾈�T�=V4P�Y�y�'M1�,�r�I�$$Lp�kB~���>��L��&���ç1�Zi�c�-�e:E�S�s��'�N C��T�OH�A�OQ>A9 E7��I"lQm�DHT��Ovt�L�$���N�"~ґ� Hl�bt�Ӫ:�n4��� �~�@V#{��O�>)p��͞	N �̏�SŜ���"0D��U
��W��DJdk&o|Z�0�),D���a��s88��,� 2�T���,��9�O΍Jt#�uX48#�Or�(Y"Oh1� ǒ�c����P��`<�\C�"O��!ѧ8�r� [$)��"O�,Y��#��0x�.��)�c"O�yؖ�V����I6/͙X�P4;c"O�qy���$	��1z�oU�$}�9p�"OD���(4�QA� s�慲%"OI"I�b�6գ�FA�2Y$T�""O���R� ?�i9��UL0@�"O��9j��(@�\3�钾�Vh"�"O���J�=@�@�*��H��!;�"O"���,:�H#�ְ~:��"O��كa�/]���k\�T�I�c"O@��#Ƨe��+$G�l)7"O�dÖ2R���
�K;*�\4�0"O� ��h�f�	w��5*,���SQ"O��ТmV���� �4+N���'��`�U˘!�HEK�*��V�0��'b*�QC�ؓI��J �]99���+	�'f�qI1/Ūo�^d��'��*��H�'dr���˃2�v�QG��� p���	�'�,�{���~M�V ͉�hH	�'�Ԡ"��_�6=����^�p��'����.�2��qa�R���b�'r�-Õ떖���a�gT�{�x
�'����a(:�ШA)�!E5�h�'����AJ�%\����B�x��'�2�qB�D81���W� .��i�
�'�8R7`��|:ta���B'6��
�'�.�KNw�Υ��R����	�'_�MeO^��
��4�Љl͈	�'=8��'�s�,,��jû	1��	�'S��1��S4P r�h4�H���E�<ya+ʯF�xؑ �Y�	 ��A�<�!�̋|h�"	K�vl9֌�a�<A�cѪD B��t�<X#�	S�<���
^2$e!f��SA��)$i�R�<A$b�1}�p�Y$��=k��	ɐ�
K�<�7���R��$��=B<���jn�<q�틧W��+��F�����֣�j�<ys�z�(���4�]�Cg�<���U�uHb��F@��T �)�Yz�<a S��j=�T`E&jBz��&)Zy�<Ia��LU�U�A	r2yy�B@~�<����,�t,Y1倠Ip4ab��`�<�#K�r<9�4#�����x��B�<��m�!d��%�����-�<�@���A�<�d2&���Rd֋P��Ի`�KB�<A��T 0�L��'� ��$�E&�A�<!E� �C$,JJ�Z�XԈ.s�<�D�$��<cS��(G���!O�k�<�s�;�R,���X��P;'Jq�<yaEЧ!'� Q�៮#4F�q݌�y�f��dln��ۡU�>%�5G��y��8(��"�(H��@�� ��y��IԔH���/���4��.�y��O3{���b��V����œ��yB(�4M��T�-�Q�$&��y���y� X�4�	
Of���I�1�yB' $p�qqv� �FĐ��$����y�BK�u��!���&D�r��4�G��yrL	�%A	��Ά��<ei#d��y�-�Ȕ�A^)1g�c�@T:�y2oIB�e�E��&��(�;�yr��??�:�`�G��ʝ�t�6�y��A<,��(w�ψaݸ	r�Ǘ��y�+F���u�^RൃƬ�y�Í2�H�!�ō�X��e��U��y�Ƈ��t���M�N��i���;�yҥ^(>���6�ƩE���2��ʙ�y�ˋ�.mx�a@�=� �`�M�y�HN/Q�܍򔫛5��!���y��Ȃ ���R��۪.Vr�J!H>�y��ެ_Gt��`�'tܹY�X#�y2A_�g����-W��P���_��y�Cϭw�DӞO�x��$.�y�/�4�P�1�/M�6�уSJ��y�%�f���S@�5�~�p㮁
�y��+lk�}�@�1x���G%�y
� lԣ�f�(I�AӥDG	=I��y�"O<�*у�I�RՀ"Wg�B<�"OmѤ%�c���� �$�,�q"O��dd�!u]T��� S�" �sE"O��؆�j<P:��CF�:�R2"Oqg��-����S;)5�1
�"Ox�B���A()���>C�lj"O}	0dHi/vY�m�73X���"O�)b7㊄��y�D��i"O2L#2B��`j�KWP��e:'*Or�7T	A��)r���B��\��'g�������d�$9d&���'�.i��B�2�H��[�5%�8��'�p$ٖ��Sw��k�名.�*�Z�'dH �I�-J��ٴ�hh��'��xX�,�6x{U&�r�d �'�����Fڷ"ۮ���d�'xj$��'�j�0!�Y�`����	K"oݲ|��'�hpQ4g��x��9z�g�b�H���'��(e'��5�N�P�T�٫�'-�!���< �z�����)N�j�0�'��a�I��_�n��G�څ�حr�'v��Ko_*'��h��(� cz��[
�'�ެ[��؛b�J�	@�l�:��
�'��3��J�H!�D��f�p9��--��e�I�b���y�M��k��Y�ȓ/���(Y3V�҉�@ �1l��Ʉȓj��7�]�L^FX��*-l�<���	�zse�sO�m��F��@H\��*�#0N���@� �) 2L��ȓ=H��)�㚏i
�1�k+��X�ȓI@��b�X�m2�J�A$f��ȓ(V��j��BO7�a�i��;G���W�>4zՏ�yt����B ]��	�ȓ|�Ja�4�R�a����U*�L��{U�9�B�S�EH
,�ք�"|��Q��\�n�a%���G3Ry��g�(��ȓi��D:`+�{�t�!@+���B����ii�N>�x谤�>h]�B�>� �!�,�0~w��9t���?z.B�Ƀe"ةQ!cG+\�h�g�&d�2B�	!Fn�2����ZI����^�"B�I� ��S�o�'q{�=sqnԧ6ưC�I)O���2�F�(d�����P�S�xC�	��k��[8��dZ֥�$0vC�
"٠Ĺ!�9���Kf�ק-:C�ɍ
C(�xbh��{^T�3�c�RsC�<!��8���9o�D��U�Q @�C�I�Hb�@���)d���j�	>��B�2^T�}�o�	�ƫD��zB�I�9���+�+��7�ޘQ�� -{n�C�I�#nĔaT�޲���2Ѝ��F��C䉢&�ta�D�\���]--JB�4��	3F�=J��$)��M�C��%P!�\���}$��H�$��(��C�I�}Ռћ,��!Q|�C�?msJB�ɑ6����29�PX��	KR*B䉑<UT�ի��9�(S��L�0<�C�	f���3��<Ϛ1�.�C�I�-�x��qbߖM����Dd�lIa"ODcg��%z�(�����AO��y�#�5f�u�� Z +�U�2
��yfӪ�����FK�x�x�81���y�#�9<fT�H�G.wZ=kʖ2�y
� 㕥̯[�D�ьPb�I"O�� ��^�_1�[�( 6��:1"OҜ27B
u̓���=)�@��"OhT4o��>\l%i���o�
��T"O"�&�\�<�DHA��4���q�"O����c���p���%=�ֈ��"O��'�m��tǅ�4XH�"O�pѪ�>0�5�QF̝Vx.P�3"O�x;vC�<��D�0w@��f"Oȸ(Mɤ!Rb�Q�FŉE<	�"O�u@����dAhkP��x�"Oh�{�b���X ��BI����"O����Cp��X����'H8V)	"O�)���!� ����l1��SU"O %)C�-n��PE> &�y�"O8l���^ l��� �h�*��Ђ�"O�i3t�>I���1��*,�J	�'�+1iZ/A
� �æp���`�'��@��dӧ>=`�ʧ+X�~ɣ�'ن5����;�)T#�Y��'� ���U��=�@!���� �'}��k�G�20�BS�Ł^�*�'��� �ei���3���	z�s�'�E���<n.�҅��6{:=��#܂D���.i�@��
�)&@@��ȓ^��q�e��f�4���@st��ȓB9���S#��`�:��J�KJh-��Az�����0���d� �ȓ=��@����<H�獁�P� T������������V!WN;f݄ȓ\T�2� v�x :$D��1��,��,�*���t���Uͭ}-���vx��U�M�5����	U�g����ȓ,3��.�99G���$�x�� ş@�<9EA���pXV�*Q2XW`~�<9 j�;�b�3Θ��x�[�c�t�<�'��:=f�*�%F0uY.�C��F�<�*�)<��Q��-
4�8xD�B�<I�hU
[�\@�AY�f2hPi�dK@�<��~� ����W�
��rϋ@�<aR�ԿjT��Cև}ºm)A�He�<�c�¦*Y�����i��)��,j�<�0�
pHr� �/@��4+^�<�+Q'|�\ 0�I�D:z�+��V�<�q�X�]�d$�J��HP�#Ff
V�<�6�jo����M��k��Z�<ᶋޫ��)�N�'q��D{�j�z�<Ƅ�F�@A)%_%4[�#���x�<�b�Ό	�T׏��Z8�t-Xw�<9�M��1Y,jᔄ�Rp�<!f�8^���J��	 �����Vl�<Y��AS���Ǧck��M�d�<y�#�N:���-´e��y[���U�<�P��Jv0@C"��	E�%3w˒O�<���C#�T9�6S�h��)�ĥMH�<�V��p�lxW�5�t$��F�<Iu�6�(��"B�'���c�[�<�e��o�&\)v�� ��}I��	Z�<!�_�Nj��V�
�"�e��&V�<1���H�Z@A�Z�.�B�O�<���ս8]��ȕ@S�Kᄄ{��M�<i�    �