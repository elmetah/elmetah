MPQ    4�    h�  h                                                                                 ��C=W�������[��!&��2��vS��/1�T�*�Hq^e�U�� n025����$w��b�!-�V�#�&���>g�FĺaQ[Y|���R ���0v�z��j<׺��x�h�w�U�K���z��I]׎�@1)��{<p̠8�S�T��d��ՙ��w��w�Da=���"U������moL��Y�|��=�׬ݿґ��Mï�W������9��:f���g1@���|���j��=��bK�7t�p�2�9̋[Up(��A?.������<�2�/���iZL�vq���8�]�b����As�P�ܲ�Z#�fY��(@�-�,���ܸ�B�[51a\z����qc%x-��s��׺_�T��H0����w)�2;aO�:4��=�ʰh�}�����(���&�H>�ė b
s�����	�5�,܂�L4�M���z��\�8��>;���,�F����bV�z�����
2����ɠJ-6�X�uUT�����L AL�~���؇؋��K��e�Խv0����RS���ϥr��h��ݠ l`�j܂��ă�V���w�K�0����8x_��zG6-�0��tQ��dV�H��E����C#[Rz���N3��67��w�fi�WBa�g��D%�{Bg6~Z�\�9��T�Nk��7Nx���P|3�R�NX�/7�I��s�.��ZƤ	���b��1�W�2&>uid��!��5�>?��q>�����رϢv2WV�t�̩g�t�C�1��FmiP�� (�Qs*�1W�ljy%�V��H���V`9�)�L37/��Pɑ<
�T���"���I�]�e�:h�ƕT�>�p
�L���?N�d3��j]�V(�ӳ ΡhH���/y�QC�"`t`ޙ-�vz:�8�5����($�=�ky��Ryl'����,!���=5�̣�Dʶ�`�4ŵ$������o�B|s� ��������A���S)i��8Ulᶕ��N�N���J�^�z�K�Ѯ����z�D`4c�"lC�b���H<��m��6ʁ��j��`l�g˂QV��؟�@�?8����e�r����>�g����&p+	�.E�[��{�;��M�ă�����~��9sL���|u��z�rW�2$��>V�� '��6*Z��y���_�������*s=�����eV�.(f�ٖ��g����3�mꏳB/^������F�v������J��Tj�RNf�j����$m���b{������`Ѷgb�<��ܴ�
�G�'�>��օ����ؠ5�g�J�6'��t����:QNN$)���"��p,gm*�<�BP3��IYwJtWS� =�G@�`��8&�P:����u���P	*�(<P�l�aIpl0���F�?;F�jLE�����p&¯Y�ou��\l5���p븼\��O��R+�n�z�G�8��H�ݟ�9�hv�a�f�p1C���T;��M�H�c��֮�̀�f$���|�_��=
1�ZIM��k�x8��-��򍲵4��'��pVR݆F!���+��T�c�{9�@�HBh��$U^b�2 h��SH_��u?�;��GT]�����3	�L�%�ô��	����8�k��t��1��*4���R^�TlY¦� uf �R0! [C,�XZ>6�C��=k4��B�A�b+b�NC1,���M����5�cЌ����Ue��aJ�K�=��¼�:��k��6횶�Mq;�����{l�v��N��]Ѓ�C�1.����n��B�t&GO/��㒹�h��M�Hd�CbU�0z�G{�/�]������������dpF#9r�7�%�:��%��Ф{N؛%�p�-���5w4�F0�ӄ�q����^}j���ڭ?H*<�XX:$�Ri̔M�Ň�,Vc���h�Up͑H��J�8���#��l��� &$Ϫ�M?��b��ûO�Y+��{\��w�P¬6!��i/�j�9��1^��Ϧ*4'�ls��_��;�,[��ӥHj�� X�c"�U����q�����w��bXiQ��{��'�����4v4�����d-AV�];��m�N���QD�s7�ګ�Sb^�� ���줫�E쿬I��;XO����R�n��0���h�,����ΠIT)�dz�����!*5EueĲ&�¤�����מ3��|� �:�Bh�%K�Љ	~�}清��!-��0���7ӓFғHչ�{]�@�)�W�+Z6�9K�</�<;�񻫦WFs�����n��i��皀t���t�WЏ�ը.�ê�9�]ZzJ����	����}��v��c�SZ�%����~��ۼ'2���{� �o��=7�p tT7�r|�/���c�ZXX��l8�0#=�
�ƨ"�۸����5��B�`���A��^I���ŗ�`&
+_�#�a��VY�Дvv�t�ṋ�Ap6����L�TJt�`b� ����痤޴sT�G©�'�{��X�3�ZUQr脑�E�����6�n.Ξ�6�2��l��_	:@.��,l�F�-�VF��y��F��O$P("t��:�&v|���o�nK�h�P�5X�Vo0M��2�E��:~���5����k���%hWVۀA�7����4MD!u}��rf||�Q�Sm�Ԭ��{,�{�E��2T\�Gδ�#�qr���0�|�g\
�b����Yj�ah|k}梆�~��@��ﳝ��q2.�Y��/`�t��Z�_b,)F��E(�;��0�ҋ�H�Ƣ,�Gu�H���SJ�Щ�m��OZ�t����1(��@���6�wV�)�����0�%���DML�j(�Kg��Yqj���t画�Y½p�04���/�3I"ux��2&���&���|mc��	���v@{���l.ʮF��3�c�1���_��~7�b�$a�?#�����:ʄ����ÄS��v�ܥ�F�H���Gj�;@��T�)�����\UsE�	��g��g]nv���P���;$�{�ȍ�f�O�����A:�~;.K������<\�}�Z��Yr�pϴ#<7�����d�
�̐�l�huf�j��<Q����eȏ-F"�4�I ���a��o�'>u$|�^	�*�oV? ۉ1�_v�4K�2Z�J&����V�[/a����h�71@b��Bd]��֑oҏ�()o��ݶ>��x�C�DxG��wP�\T��x���.K�^a��}�Y���E
S��"Y�d7x�W�B3�����G�@j��W�/����^�iiU��x������g�uC�P�]C��"�h���2:�,*,��
_�9'N=U+6��\��;T��<ͥP/\h:��~Z�6, ��S������AC��Pr"��U�f� p(���G+��W����/p��\b��zPF�h�-����	 ���̐����k������r��2�ϋ��m��X���+�!}��69@(#PP�! �>�]� ��s��1�O�g��Fܽ-�4?ඞ�a�\�p:}���	�*�ê!h{�b�#z�
��O��lӠe_{���`U/�T�6�� �A~�:�J���F'K	ݧO~wvQL�`/:���+����ݘ��l{�}j�(��t� ľ���~-�r p�U����xz��z���-�V��<U�؜V�d�X�x�#v0�WbN���q#8�G�vf��͙�c�"B�D@�B�"�Z��b�t�7��u k�V��?�x��P��=R;�t�VڡJK�e��.�l��%)������ЎWg`&GGd�չ�h�.>:�qiS����c�Jp�22�t2�gh�C�D蒡��Pm(���*�I��G��y`���6ӄ�娞f��`�x�g�N/#�+�<E;����~m�I(&IeNe������
�aL���?� �.a�j��^(_2� ��:À�
��Q~``�Eޔl�v�X38>����0
�FM5��hl�2���6!��=�Y-̾���1d��D�$�qdr����D�B��B Y�)���ڒ�ō�S)���8�xR��B+NL���c�yކ���Y�i�x�8� D��x�������^Ǥ�:���:)������a��s�}�����Z+��Z��j�ne���u#�8w����&�K"��p�[�h���r��#�ľA�<���y��є���K��|�F�z9�����y�ǛJ��1���,�P�d����'G�Jǥ=��3���ɶ�f�;i�Q	��Kߥ3��6�.*^�x�L=��@mv����s�C��T�\rRɘGj�u�_*��<j{퉱�c�ǈv�K`���b2�Nf	��EYS��>����ྪ��F|P&�gn6��t�u��ՋANI��ZX�ǲO,�+*aPB+�;�M',w��S�y@���4`�xU8A�>:"��P%����L�А��w�p'?���,�?���E��L����.M5&��XYIAu��h�_���<4\C�5O���+}(z�@�8�	���y��C�Pa�p\p̔����K�rH�`���}�W��@$&��|�M�8Zj1@��Mc�ܓʞڨ��h7u4AЕ'O�$Q.�R8��ӌ��a�u�>!�9/loH��A�^��� #Cӓn��]������}+T���ּ|	?%=�����²X���>]G�~�>)�,#H*��1�o��o���!�uA1n�|+ ���S�6l%���~�k3]�ǽ&��=�ԉ�u,iEc�H�E�Ep������(�������T�i��`t������Gsk��5�1�MLm}��9"��Nv�O�#���>��C �%�~n��;�G�:��҆�V��T;F��d��b��jz���jk������9N�T����x�pa�rI��%_m(�`<-�?ѹNӤ}��l��`yՄzw�B�F��m�b�H^x>ۑk��<�7:�}�RD�锈~���X�c����rp�>H�J;JiS�yɽ��n�p�&9t���5�z7f�/OI?~s\ێE���16��i��6��� L�h
*��l�~/_c]�;�,w�:�AH%� s�"�>՜�qTpN����r���w�jX$�5˖��'�j1���C4�F�|_B��A�\�]�_��&�?:���MD��7L����b�[� ~���;��T*���II��X�_��~�nN�u0֧����/�?�{*��%8d1w�{�����5 ���)���ڼ���p=qZ����:@D|��w�Ф͗��-���E!h��03�[�2`cF-�	�q�{x��פ^˦<�th-<���7�(����ݚ�����O�!�5�6���$d�Jjr�I��8b�]5�6����l����N!�Q��SuO1�<aR~����bp_֧��M�U{�+�to�Zr��6��dB̕��6��+�$�e�������������l5x��ћ4"���M^������ W+z,���V4Í�X����n�����'�M L�2J�7�b}���*ޗ?�xsO���.��6��X�:�Z�;�þ�A�'�=6���I-��4P��+_�o�.�hQlV/��sHF���y봸�wu�$1-z"�~I:x��|91�oPa�K{�⚫�X�X0hX�2(x�?O��D.�������~hǒ�ۛ�\74���-D\Z��;�wX8QBpm��������{q�T�L�Gi�#�WrZ70BΏ-��
����p�Y�l�h
j��4~�e@��T����)=�4p�j"?tR�]�Z��)��yE�*�����>)�X�,�p��G��6J��ԅ2��������+1c�@����1|tV\>�������竃�����xL#���Fa�V%�$��(���O�k"���x��.� "� �m�%����_S�m>ȏ	)�ac��.Y.%b���R_c
��sP뎲g:̝	$��l�:"y�vrr�n䷄{��>�R��
������z���I��(������פ E�H����*��_nq��Dr�~�-;?]��C(f}9Ȥ�Y���~6���]���>�\��Zf�Tr�'�^l�����G��eJI��B�h��jW,Eι���*�4F�X�j����w||p�o��>P|���ŜyV:�&�lإb�46��2� �J�@����]�[*풪<��hk�@}բB�0w��U2��.t����PJ����x�!��}G�X�+�mT'R�����.F��a�$}|��Ӿ,
�DN"48Qdr��W�A3������@%�r�o���9Ui�|�xd���������P� 9�.����'�,e�����	Z��9�0_U�c<�w�����n��<95/�b����Z�V�ر�nO'�銥��A~�VP��P5Hf9�(�*�b�?���3�����c�\�2��u47��-XrC�$Ɩ�U6�ұZZ�\P���mg�2�]����sʦ��}g�8t�M(���z�>V� ح�s�q����1��nP����4�P!���鷏<ҩŔ��_��3���K�߰����
���Ȃg���h�N��U
@��qd� w�o~���-V���K$W��^�v�@O�N	�ʌ���'�^��S��l���j�S��O-���v���mq��槃�\P�x��z�W-���wV��7.�V̠����3?C#�.��#}N���/e��~Ef�o��$���D[x�B]/Z�t���^��t
k�(P��P:x>P��R���h�m��m� '.����Zbj�mY0��W�&�85df��`>5K�qĺ�o6(��]�2p�tm�g�<C�wΒ�q�P(]Z(�[�*v�e�"��y�A=��}��㣞��Z`�t*ӂN/�����<���,�zy6QI�Me	���K��4w~
x��L3R�?���)��j�(�d .5>�T���Q�jQ`��cޏ�fv0�z8�(G�Q�"�!AZ�,l]����`s!J��=��;��̞ʬ���~$��uG��9-B2|� �r�8���Ս�gb)߀�8��[��ZN���K䃔�:�A��D�5�s{|D�CF�b���iU����'N�,˜�e�p�ւ���@�x�TY�����uȉ��<e���t�~�� �&&��褼�[)ZS�qµ�oS���?׫x�t���)����|��	z�5Ғ�ESԴ�5�6���,x��ݰ���R�Ń$=^��B���de�f���������|3�U돩1M^�o؜�p�Z�v�I��΍���j�T�ˊRD�mjs�e�����{�bʾ盈1��`K.b�WqAVq��A��]z�>�qy�;�pԛkk�g��O6݁4tiN�p�UND`���q흂˒,�D�*܃�BY.��%sw�߬S��?��P#`K8\�4:��N�+s������^} �Թ���.p�m��3�?1� �L��d���1&���Y�m�uLE8��%|�n��{\~�qO1�z+x�zDZ�8mN#�u���/���a��pg���~؆q�"H\0��D.���j:�$a3�|*�D�3�]1��Mpfܮ|�#���C�d4|z'�(�Li�R��?����F�ꔵНq�9j�AHx�]��^ex ޳���8���l辽����T���ַM�	�
%��B��k��ӏ����G�����T�'��*�a��� ��z�4u����� �
�N6�k2�g��kN� �8������,���C�X��G��8;��\����������/��s*r���I&g��՘�TÚ���M'�p�-����]v��~b���]�C&����n{�d����}n.���u��-��d�bK�qz\w޼�'�D�݋���گ�ʘDA�p|��r�޼%:�-������F_N����<�E���{�O�wq�F曛�HĘ����^s2ڑƉ����<2�?:��R3���B���c�J`��Np���H�J�P�T(��"�Ve&Ù���5,�̻�O�X�Yr�\i���.6B�i���mKg,��d�*�Z�l�c�_���;�L/����H��E �f>"��wn�q�`��D{�m�%���X�\�˱g'[>����4�
Q�¬ð�A�i]�6����uS���D
7�U��5_b�* :*�"���;�ƭ�KwI�WX�N9����n�}�0��I���Z����V+��A?d��a�v;�5��b������ڗN>Ḿ������:�ep���п��s�Ʌ�L�!�
�0�g�-�F��KI�{�{D�˦�=䯥�<Q���2c�qz��뿜5n����y�zJ��Es�����
�*ǰ�XS�d������]
s�8o�_���so,�5)S��$����~t����Η��˖�&�ɰ?��t��rrjI�e���
M��mÛ&K(����w|w�e����G5S�֨m�w�^��]B&��9h+�}D�WS�V���T��@�n����B���L�nJj�mbX>g��ȗ�a�sJ�7�_����8X�a�ZKF����|O���G�6���TD���@��3_�Ĩ.�m�l����c�F�3�yF�j�2��$L*�"j�:SfA|t��o�s�Kv���eXsؤ0�@z2��;�𙐁*���Ai�=V�S8Xh���۶��7��;] �D��ʜ$$`rT�Q��}md�2���g�qz�V"�T��G<L#���r��0�?H�s
n`�K7CY�C�h�Ȯ昊~Z7}@dΝ�ӣ,gA��w���t����U�p)��eE���-�ҁ���`
�,8%R4�幵Jl�Q�����j2c����1��f@+�#�,o-Vi�N'E����&|���	�����L�Q�A��c4�����h;��)2�s���0b�MN}�);"+���(z�������m&�	d���c�Ȃa.�5��?��c%�3��)���p���-%$�B�5A'��p��)�i�/|����������<��~�{�u����rP��|��o2�R�E���1�=�4K�nl]��d��9�y;Z4�����fXC��Y��w�y~12�H�H�{�[\��Z���r���������X̃ɒN����t8Nh��Oj�a��>�i
�Œ<F�X��ӥ�;����o�>�>+S|,@�`�{V5�n����m�4Q1(2�J�B�J���S[%�����Uh&E�@�C�BZb����>���^������xE%�����GvՎ�NTb٩�Q_.A��aN��}7��|
I�"�d�|9WA>3����v��@�:�������tPi�Vx�[����S�+��PW�R�(7�^?~��3+,�\�JJ�U?d9�2�U������la�IW�<C�m/�} �RZ]����7��?h��饧u�A�M@P�/�Kn�fj�"(qj�}���M��Ӧ��,\K#�p8DtO�-a��?���п�Ҍ��0��UW�h692LE�kApȎȲ�!��}BS��l(Y��/>��K ��Cs���E�g��}J�3�#4T�ڶ�x����9��s>� ���׻����K<G���%
C��=�S��#���B<U夙�d� W~�� �ؼ3HK?�#�E_�v�P���ve�r���L������>l�=�jx�O�*�}�4������h��AX2�x��"zy��-�ɲw{��v�V��G�V�9#�L?M Nķ��[F�}2Lf�-L�h�����|Dv��B�[�Z�0����Y�%�lk���H��x�v�PͯAR1U�C������.�oƵ���(A�� oW]v_&�J3dMP&���*>0��qB*�*�iC׃@k�2�,�t�uOg�3C��p�W$oP�Z�(��*�ڞ��AOy֤.�lH��{��`j�@ӝ�5/uJ���1<����t�I��e����2�e
Su>Lnˆ?B5$��jn�N(�O� �W��ŵ�SUQ���`EֹފJ~v���8�R:�"�Y����TO1��l��q+!�v=f�.����'�t�šK$<�9�V?��N!B�00 ���S�ڈ�q��с)&�8&�����$N���惯�߼{n��"�+D1�����s�;ꩤ�4̢�{ܺ@J��>��8	��sS���M��̐����`~�e^S�H��4~��a�&����_(�[D=F���J/��4�zr��o�;�J�����|��Oz/�ђ�E��_���%�'O���<*�ڄ���y��@`�=9q��}����3Rf�_"������73���$Y�^}����	���cvӶO�)��{�T�Z+R�] jNof����r�C{�ٯ����`"�b(@���I����>�t֖cY�+�����gdV6���tX|��aBN?.���=:,��_*W��B����C.w��S��;�X	�`�\8w:3:5��o�%c��ͬ�8Ю-�p����2Y�?��O� )L��Ҥd�f&�ܴY�{%u��5��_|��\�߁O�ߒ+s��z���8(�f�qwX���b�aO�p����C��DH A��+:��v�ET5$��i|����.Z�1��mM����N<ڞ�O���4�p�'���G�^R�UR�0�8��]����9�"hH�Q�.^sJ� �D����+�S���+g�IJ�T.��ֲ>�	��%��H���M�N���ɩ�����Eo��"{�*E�1胜����F��u��u\ ,ОI�]6"�I�"��ki�ǳ��M���z,�"
�>"���r����ƌ����|j�|V���������������C����'��M1t�ht��L
v��/�Ijд0-C6P��z�nVƽ��< .B�Ҝ�
@
�~dId �Zb�LDz7?��щ�������
����)�p��r?�%3��ָ �u��N�"�I��N(;w���F��ׄ��Xܘ��^nF��!s�p��<M{o:���R��4��&N���c�)�yo�pI
�H�~J_���/�b�Lګ��,&m�^iÀ�@���g�O��4�\Qc��!'�6��i@�΅j����^�b*�$�l$i�_��Y;⌃��1�H�� ��'"����R�Hq�p\�ߒ��h�K�-A�X����n�'�k����4'&���D���QAggW]lw;�m��5��QDR0�7�C����bo� ����=t���o�}�4IP�X �+��6*ni�0L5�����
b�1L�~�dK���qM���5v���d��o�r��gs����:��D�V1c�ڵ����L!�\�0iM�(�vF�x�A�{�jך�V��_���<침�-�9��C�n��PH�����U��ŭ��ko���H��=��ex�w��.(]���s���9���9������S�� �2�	~O�#��L$�A��j�'��+�t���r�hh�@���%�l��!H��.�2+��,�ׂv�N5.��=m���^�������s=+�������V��w�����E�n�[��Rܪ�É�L˓J�֖b3��Y_��uShsE�iº�����X��Z�p�y�W��A�s�F6�ޤί{�c�U��_z:_.��+l̏'���SF��Iy��\�� �$gGv"���:.6|��o��IKq�u�a�X.�U0�HI2���B�e�{����Ŧ���h=j`�ѺB7*8�8F�DҸϜ�,mp�Q���m���ӵA��1�T�G���#��zr��0��Vcbk
~ZQ�&�QY;hM�K�<J~�(�@�ʳ�W��x���s�qt�<��Py�)W�QEYZ~�H�.��"��;܌,s������J�F�J�(�/�|������]1���@�u�'��V� -	�J��|硔��1����LY���<�X��A�,s��Ƚ�� �N�L�^W��C�$�"�q���M��d�U�;m���	�E�G|����.�(����c@�p�i#��h�P�r�$2֦0��,���߄J���4�4�i��V�9��?�p7�L�������{�ͣ_Eg&)�lE����ng2��ش����;u+ӗ9�/f3m�9�#� �~,���|��64!\��,Z\�Nr��f��,��R�̃��]���/N�h�m�jM�/�$��B���`uF�4� ��������o�R>E�|g�	��vV0ò�"2ॐ��4l�u2��J�6�Z�r�O�[ e��vh���@��;Bճ/�d7�� GY��3g�^׶O��x g)��O+G�q���T�������.<W�a�G�}�_	g3
��)"�Ţd�.uW��3����L	@����?�e�*���[i��x���������]P���Cqzټ���`�,�$���1P�98UcU\��N�5��$/<~��/-�'��Z��]�!�O����4����A�+�PC�H�F��f�	<(,�6������rƮ�!\�3M�k\m���-�o��Zr��KiN�g�U%����c%�2����&ۆȩ��ʜz�}׭��_(��@���>�� N��s�����+
���4�n�S4�������m��H�b����(Ҫ��Q����������8�
�]����ɠ��;�D,U�)���  �*�~�+E[%�w�>KZ1��Pv��E��? ����}M�>���#l̥j�
���T�o�f�O��c���(a���x�;Gz�`�-k�����m��V�x�꼰���#Ǌ&��N�贌"����f�te���S�D��_BS��Z`�%D)���&k�,�����x���P���R��Q�d���6Zt.�L��;��H�;n�W�X1&�|Ad����9Ȍ>+{�qz�c��;�^�����2�	�t���g9��C�=ϒ���P�x�(�m*lS����y(t�3��?.�w�0`%��Ӹs/������<���bp�o(�I9?�eIt�2���*t�
.S�L�d�?��}j�)7(�� ::�4-c��ܝQ/�P`�Hޅ��v�sI8o��=3��7�׈lO/l��S�@! �=!x���ʢ�S⠀$w@�CX���B�� �M�nXu���f[�)U��8�^6���N]�B����D��7���0@����D��	�ؽ���M�_��a�"L�*,�L+��Kc�n�� &؋�s���'�ۙ�e9��ȗ��u��»&�ln���[_@A�go`�%eS�o�I���j
�ѥ`��|�%|᰽z�x������*�=�luã"F)�=7��&���RB��\=��ٸ�}�"f�!	�b�g�|�3������^X�t����U�v�Cj��Ƈ�6�wT�	TR:�^j)Qw�"۟m{�1��tv����`=_�b���O��q�����>��c�����O��Ufg�,(6��t���̦�N:`�k�8��\E,��*�J B��c���]w���S�D3���`��&8��9:�����ny�<n���>Q������pX+��M��?'���9�L1 ����&�+�YZ�7u�$�9�r �W�{\�>fOg&+n_z��&8�7�������.a�Op�Is��(f�'�eH�/��3�w��� ��$��b|`��)
1QXM�����@�	y����4���' �B?�RI09���S�?ꊖ���p=9��H�r�tU^�O> T���������A�sfc���YT�J�֭OS	PN�%n;Ӵ���ɜ�ʤ���/���7��Wr*�C��>ct��$;hu҃>!� �Q̞D6�6}X!���k��]�.���Z��:`;,:��9���V$��O�6�%���sD�W=��.שֳ������xJ��5󹚢rM��Aw��~Dv�^4QY�o#�CQ�v��An1G������oI�erL�9��d;2�bA%�z'���@�za,���e:���2|p��<r�S%�ň������N�n���x�	�&Fyw.�F��������3�y^iz,�|А�+�<hq�:	J?R��b�9+9�S�3c�(���MHp��H7��J� ��
%m����A#&7���rZ��u"�4FO~��c\�}g����6L<i�֚�%���zk�yd*�.l_�i_4cp;��s�K��HVf2 Ċ�"�d�-x�q�1�z�J�c�-��� XU����'�����$54bac�M�	�|�A��]'�?����L�s<�D�vk7Q�ᗐbʜ� ��%�Xq�1H$�XW�I�e�X�6ֿn_t60�~��5)��G��@�id�{��l�H�:251�p�KmZ��M��{ �����:Q�������U�iĊ��Z�!Ϻ0���#ǺF>N�X�{�yh��n���.�%��<��V�([��'�C��kB$�x;6�08� 6����� ��k
�{�ᨚ\N����]����uVU4
��j�%b���S�_į�{G~*���$0����8�f_G�\o*t�c]rh����>�F=��ﮛ��v_���\�G�6��e�5	-��L� �#$^E2�?��L��+���M�,V�.��	����m�n��̡��<�~n�LGyJ`�+b�औ)z�e�s@*�{�g��X��ZA��T,����!L6�Y�
ҐŎ�q<_���.h��lp�ę�mF�ɠy�����f$�� "`��:	&M|�ko!��Kl@	��VX��j0�p 2�3�妯c���Аw���0�	9�h�l����7����-D�h�ZU�h�~QSB)mگH��C�g�C��TH�G:C�#��frk�%0s�`~K�
�f��O0YVR1h�@��~:�@�'ܳ	,6]�����1)�t#�7�K�)��=E"��cm�w��Υ,�<�[����i�J"�zZ�J8��`�X�d�K1�@a]~�"��V����.$��=��y��0U�L�T��7���GV�0��H(����)|W����Y���"�Y���A=����^�m�A�	ڞS€����.6<��n�c[Nֿ�<��C�c�N�i$��ަ+�7ه�����e�2��V�D�]ܑ��ϴU\�k/���%��@�7���b�HS1EB�0᧐@�j�7nb'�Um�ȯ�;�B����
f�F�tD���,�~'n���;����
\��KZ�/Nrg�N�����g����)�v�?�ꃾh�Z�j�bn���}���w�F#��{�ˠ�Y�͘�o���>�K|�7GԖ�hV+��}r$�K�4���24�J�	����.([Qg�M}6h�ҏ@��BP%��?�g�[Z��w����'5x��S��Gl.���T�G+����.7�a	l}�L�$�R
?�9"ż�d#�Ww.3 W�,9 @V
�î�2�ʗwiA�ax5E}�}������Pͨ��^�TZ�=,}��	YK��9��EU����X��~���&�<���/�'� Zu��o���w#l�]��A/*pP�xZ�A@3f ��(����J�C�Ɖ" \�\�d��f��*��-��I�uxb��2;�B��W9�!m��^4�2����a�Ċ���}�z %�&(�����>gz 	4s���;��|�ܩx4�E������������*ⓒә�����,Z߁�t�ڨ
���ȳd��g!���U�Ξ�"�o HrM~�f���l�2�yKuΊ�;��vw�8�����D����*�oP݄�Gl�-jn���ཛĪ%�����^�������x�szo7c-F.��(|�h�V�����ds#��5C(�Nz9�]%��f�ۺ�b��ND��B�5Z;�`�̏[09k�^V��Dxo�yP��R'��1ȡ6�Ű�#].�I��k�.��p��V��WS[�&��_d�J����>&C�qհ����jy˭6��2�Ht��g�R�C~���PY��((��*��uݳqyL���=�����Ҩ�`�n���S�/k�^��'"<1����CjQ:I��Ye:���MM��m
	Q\L�`?U�8qLj$��(K�< U���,�v��QjW^`{Mހ�avA�8*m�X����4ֲܩ�ol.M��![~�=�l��*����{�$���y���}BC� E�f؉�z�~lN�A�)��8\��|�N���|�X��G߲�3�Յ��$��Dg���	�r�)-������ ��<���)����n���i��j�^�F�S�V�.e���ΦE�e��C�&7���_[zcD���ǆ ��ĪƬ���eV�� ,��7��|��Sz%JU�y�8�e�����]��	�P��L&�6yi=�m����51<f�L����7RZ3�y��^3+�8F��f:v�� �����mT��R��)jS��K_��Q}{٩���؈bS�`X�b������1���.	�>��r�L���=����gZu�6n)zt�I�A��N5*���yմ,�4*M�PB���9� wQ��S�'���`|�t8�H:����w�m�/��`Q��ѷp�+�hx?��o��OLl�ˤ�{x&��Y��	u}2@�+�&2�3\/�O��+iP4zUf�8�ܙ
���ů��a��yp8���-g��C�H�_�Z���,���$�p|�N��$��1�'�MO@���Rzڔ^N�ԊT4-�_'��&=��R�*��*��n���7ڝ� �9Y�HI����{^)u1 �ٓڐ��I�оN�����QTdȾ֨�	��%)�����Dӳ��h3���{ h�Sc*�����I����W���u�4`y�] b� �?��6������Rk�Axǩ�w���O�u7�,��4&�����
ϊ�1�Ɋ����2D�@vX�DG<��R�Z�+�3�,�Pr�h�M�t���.��v{/(�xh�*6�Cl���n` �3�N���bM�������dV�Sb�Nz�.L�V�K�̗��q����{�u[|p�#Br5I %�x��L��Ыg N���MzҨ�o�Aq�w���FwU ������e^d��ףN��A<��G:�#�R��@�tO؇�F�c�G��/Lep�}�HR��JU%����G��:��9b&!3��рf�~� -O�F��.�\Ƿ�W
�6Ri�*g��C�Q�T4�*{sl��O_�O;�l ���H�� �L�"}���-~q@�:�"~�^̖�u�X���'y�-�d��4��j�����A�R]�X���}��+�1NG�D��K7�~��x#b%�w k���s����.�3`I��XXV�Xֺn�n��a0�B���� EX���E{V�d�r�g<L��5���9�����(����kC���:�����j���䋍�f!Ta�0����zF��|�{�Fא��rU�`<"#��#3��������\�󘖲��;ޟ确p���};n�6Ꭸ�a��$D�]����(�ND���W�C��=_�S�Op�(oq~]��N���,	��q��������t�>r��ʊ��]́����ț�����?���ŀbW��l��5���чň�H�^���n��G4+�0���p�V����D�~�{4�n�ok�o��9ssL8��J��,b�
��A���8s;�B�py�"3X��Z�%]/�֩-Ϫ����6z��eGI������<_p��.C<�lBp�4�?F�ĳyW^�cL$$��"��x:�5�|%��o�k�Kgy��~X�
�0Ը�2�j���ݙ�������d��h����I7 E`��MDHە����cyQ�om��I�	�m�⾱��#T�=G��x#��rƐR0.U.�T3
t���
�Y���h�č� �~kk
@��ѳ$ ��G�ޠK�Vkst�/�F��)E*E�	j�~L���#����,�$�ϊ����J}5?����e����Օ?_j1Oj�@��?��Vze�"�I�O�%B�[�k�k�qL���2��tl�R���z�
�a���W���6���"<b��YUM�:Z2�KM�m���	m}#���>#.�o��p�cv�c�_vӎK'̉Z�$h �&^���+��Z���?��*�G��}�̉��O�Ыfy������:5����"oE�(��*0��n]<��!��jv;�y�/�qf� ����>�HyV~"N��Y^ͬ�\�ZR��rB�f�Jm������3��ѳ�����h�g�jCy��p��:xȖ�dF	�����l:K萇o�p>��o|����1SV&%/����Q�4�z)2�z�Jm$l��]j� �[]檨�hW�@�MuB˶��������/����T��,xvJB�,�`G�
l�p�T/��"k*.2{�a_��}hY�?��
�"�"�Ӵd^��Wh�3z�@��E7@���=[��ͥY�i|�x���x�G�<|P��x�yEg�G�y,Q|�9F��9��gU�Z^����%p��>�<��/c���\�Zn���!��ϛ��v��8^SAjH�Py^d�<�yf{Z�(�UT������-�d���H�\�#�a��i-D퓼����AT���m��(�Yc�2]���n �ߛHʒ��}�>c`<�(*���R>�<� Ā�s+��϶
��Wj���`�4%�ֶ�g+�#am���E�
����h���7������8�
T\��n�"��9��:#Uv���]% ��\~���W�����K��꧶ 3vR@|�:��6��������-�?%�l�j�A���R��'��!�Yu��R)?�H��xB�z�-*-!�D�c��أV����gA��#�fm�iNU�#���"�N�f�bL�yȭ���]D�\BI��Z$��RD����k��Y�x*MPLTR�{W���q6��l�.�f	�Ɠp�Y���q�hW�}y&`@�d��߼oQ>!+�q0�7�[�!��>�S�2y#�tY>�go�Cy���h��P�(C�*b�ݎ9]y����=hR�)�-�`�W���S]/����r��<l����{�e��I��]e��h8Z� �*
�n�L��?�����j0�(�w pƯ*@"�QN?Q�; `��{�-v��8召�s�g}֍P��l�#�H}!�g�=��_�E�4ʘV�V�R$� y���M�B��  m�ؤf��掍�@)��Q8��q�wB.N�07�ǃ )��-l���
�_��D�������2A�|�*��Md��I(��/��	1��du��*��/f��hf��0�e�S(��)��M�{�&��!�+�[��O�]�;��0�����CN]�`�[n��%(|�z�;ْT	;Ԡ�Ǣܦ��y�����>�&eR���=�t�.1���_�f�������32�Ώ���^�ќs��� ZvĽ�:`Ŭ�gT�=R0u�j�tɬ��q�CV~{�A@�*�-��g`s�b����+�l"���x>�=>֧J@�\K�׿g��06I�1t	v��ܐN0X��!g�nn�,	E{*ȑmBr$Z�t^w�5�S��i��`7�F8ȫ^:�Э��<��`ј���$��>{p�hWニ?B�kL�(V�5�U&�)�Yg�u8l �h)���\j]�O��+d�ez���8Y��%&���vŊoa ��p�9��R���HH�C�8��m�Y��a|$MH�|����D1�M
�������4hQ'V�s8��R�D3��%����ʝ���9V$�H�=�`~^��� ʶ����!���K�)<���l�T�e�֣��	%�t�/x۲�)��Z��n҄�)��op*VZc�PX������u�U��� �m�:�63��S�k�
��$�3��2�԰.9,p^��/�>������Lm�w�<�k�{xv�ߐ���c�����y��kњ��lM�F��<��ȋvvw�꿗��h	C�����tn���n%��,Ά�u�7�կ=�dq�{b76�z�Vf��۪��Vۋ�O=�U̘0��p�/r���%�K����$�F]�N����B��C�\�Kw�j�FR��4��iih^_B�2�����6<���:�qR�ϔ��+��sc׆̲�jBpzgHm��J�i�����g?�wp&+ɾo�(�!?��8,|Ot��ŭ�\����6��iQ�3�����HY�*VB�l�8J_j\f;�)��/H�[� �.�"�����aq{ax���i�Y{&�>@0X���v�'�\k�?�4�7ƌ�����2Ax�`]��t�6�ꦣ�)rDc�7Ś�y�b��� &H�����'5����Ih�X�p�ֵ:�n�,0}�C�
2��{����n-��dd�=�b�k��5���TXs��>�9�D����e:+��7��+�2�_s��A�_!�T0:����F�}�7�z{����C�M���څ<��{�+f�ݗ ��
���F�n���=@�v���<~���h2��d��N��ІĪ��]|���$�1��V��f�ې��W�S�_����~��\����f����A�0P��VMt�9�r^$��	̼�'�=���P�,�8�c�Ҁ}=l��m5����¹���� ^���ɻD���U+�Ce�V{p�����n�)f�ch ���LS�|JV5�b�9�
��F�Ts6��ˣ���ȎX2>�Z7�c
���h�}�Dz6un�������mv�_�Z�.��l}������F�߂y�س�&$�^�"V�:�e�|`�?oW�Kb�Ěr�GX_[�0� '2���\E��א����@�����hn��"T�7����w�D�W��u^��Q	UmP]��$��]�K�%�T��<Gpʢ#�;�r!�?0�F��}
��콷�]Y��h3�~Ƽ�@P��?4�S���{�~���tY�v�A��)h�E��ԙK��mj���,$������љ�J��#{#)����V(��<�1���@�<��{jV�7�:��d�e���6iK��;BL*
��-���is��׬����w��������������"������UM��[gm��'	P��U���.��X�+��c�Z���;��Ӛ���~$1��!�8�=�-�ڄ����Ú��m�9���b��a�@�]XB���2`3�>E�b���unXq���%c�;���efĪ������z~NQ��P�g�J\(*�Z�Qrή��=�#������,�y�`O?h�cj��Osd!��E�1��F/��1ir�';9�5o���>��|����5V!�g�3S-����4�}�2��JHZ_�O�d9#[�����h�@<NBFh���yQ���w��^X���`��x1���G{gGbNr��TN6���Y�.-=#a��_}#�TZS�
5j�"{
�d��W���3u���qN@�Y����7�̀;�i�νxk�\�s'|��o;PC#Ô�YJ���T�,�=���H�At9I|�U�(��B�tN��v�</��/�'��JjZɯ��T8��?}�mꞥAQA��pPdf�7��f�2�(]9)��m%�9N��?�ґ�\�%��\�����-�[���䲺�%���6���xWf�T�2���Whc���
��}�"v��1(�J��>�( �sF�*�1�y�2���˜4��p��L��~�9y�m�`�	��ͪC��r�N߷����W
�:�)-�,墵XUQxd�� ~a$~�<:l1�ب
�K�h�1�Vv-��u���	>���x�%�k����l��jd~��z� 26� ѓT���Y�;Cx��zeD�-��zɞ<��>�YV���.���{#�9�dN0;��L���@�f�	��N0��L1D��?B�M�Z�_ʜ�	���Mfk�"'����x�)�P9�*Rs���_���R��.���!p�� z��+�WI��&;��d9��
�C>36q��э���?x,�	2T`�t�g
�CtVS��-�Pϑ�(^%*�|}�i!y�q=�ز���p��C�`V`��	t�/a��M-�<��31M`mIJx�e��(�C"�_�
���LZ��?���4j��(�
W ��r��C�,7�Q�?�`�DC�v�5v�� 8�9���v��k�h�Dkld	��!q==R���`��ay�1��$(/U����B�A �,ؿ�t�[����)��8�ds�r�iNnJ��C[�˘ߨQ������,TD������!����E����}Ժ�����j�����_k] ��ؼ�u���a�L�e�>�4;!{�-�v�l&�;�K+[�	c��b����� I/��R�[N%Ѷ"��|2;�zM��/J���;�=���{�NVް��2�A�Ɗ,=�`k�i���k��f�'��sq���K3Mʋ�7�^�!h��
��&��v�������g�eT'��R�gcj��
��9۟�z{���ʅ<���xs`��bK4��������d�>����-��y7��gPfg6$99tD	��w�eN+���|tz�)'�,$�*CevBMg}����w���S�/��*N`�.�8�f}:��r����	ɘeP��C��x�p�7'�1�?��@g�6L�ܔ���j&��>Yk��u���)�B����\�O8�d+_$�z�<8�]@�H����e^~a;NApnP�՗݆8��H��S��5��^$��|1(��D1b&�M�Q�5�Xڊi����4�1�'�nx3p}RZ>��7'��ׇ�`�W9�KH
��]^�8 �ǵ��C�?�����5c�T�#�֞B�	a��%����J�Ų:� �5O�Ө��Q����*���ow���	�M�uc����/ ���5��6��(�ɷk��ǟ�;�_Β��Ev,]y�*��g����(ߌgA���[���䶚��z�p��l�Z��A&���(���Mn8#�Ti�����vqߐE'�Р�EC�8ҟpn�y��]��l����vɓ�jd��lb�n�z��м�^�K���M��v}���pr+0%�>���1��r$N�z<�+�:7Ew'�ww9�F-qi�oB!��^Z�z�����\�<��:z6LRf_���2�$�fc��=���p5q^H��fJKξ���m�8���&U���N`�����SX3O�L+\=���m*6���i�3 �V���_�J	�*1�-l�X_�E;���\o�H�� 1_"s��վ�sq���K1�T=��*X�)��8cQ'o�t���4�u��j�6A���]X���*B�!��D>	i7�9_Қ=b��� �d��ZF��[�����I<>X�I�ְ&9npV�08��%�����Ν���d��@�]i���5b���o�9�0��މztqEߨ�����:b�V�B$��F���zׅߛ!��0էЮNoFOj��_z{g�׆m��('��ַ�<X�C��8�*t�w���S��[��������m���K����Ьܵ��˫���]W�R�_�&�@���6��p�S�����~����ą��
��C��wȔ��$tU�r٢]��WL���P�� E�_��IѨ&���CC�bb%5������t�~��^���$�,�}�;+󃇾y�VV����N�!_n�����2���yLn{�Jєsb�� �EH���Y�s1��&�g����XM�Z�Z�幖��e��V�6p�!���Ou)(6_fP�.�e!l����jAF}ys����k$���"�!Y:���|�(o��K]���FpX�0
��2
v��7@i�Qj��H�z�\��h)���=�o7�_�?D�}��+�vY �Qd4�m�8�?n:����v�T��G�#���r|��0�X��
jL���YX@h�a0�D�~!.�@�h�ZhQΖu�Vy�OFt��J�<�)�]EE9fԴj��l��cQ,_��,���aWJ3�(6��������uԕ�881�z6@2���V0*���C�6��{���fL�}�(Y�*������1�ت [sº�W��TZ5���"�ҵ�����p�o�A��m`�)	�j\��Ζ�1.G6��檌c���UIЎ�|����$�|J��٘H`��~`��aU� D���!.�Blυ«\m���!o�qݐM췒�!/E�a��X���;�HnS��f�;���2;�Gd�%g�f�TV�%���~r7~n��:b�"��\C��ZH�Tr�"'��-���������҇(w���h2��j9��Nd"�.f��?F��>ތ�U��[���o�'?>r0	|S��g�V�����|�'4ؠ�2xg;J#��F`��q�[�8�^8h��@JOB�9���zΑ���e��¶��\x�k�bt�G�#|M��T�]$�Xh�.(�a�}���u7"
���"Va�d�7�WH;i3pǇ�=�e@�1���Q�8�[=+i��x���n�L���P�p�ï����~�/TB,ǅ�Q�!<N�9�mUH�����v��΃<jLw/��5�X�Z$}�IͲ��F��}���C�A��P��`�2k�f1+�(=�����,s�̽� \R�Z�W,+;�e-����J��7O
�ӏ�6�����O!�2T6����ʈ�2}�&Y�u(`~����6>xP :��sa�Ϭi̞�>�ZU�4[Z��{QG�ى4�Δ{�����9�=�쭌��R+��˸j

ۦ����">â0��U,}��E� 	�~�׮�+��cP�K�e��AFv��,�l͎�U���
ݵ�Cl8��j��ׂqn�[踷����O������\x7�)z�z�-��@���S����V��Z�강Ǧ#3�T�L�N�R�:䄔�f��#�/�r�?��D���B?Z̻^�ᯏ,�k۴��Y�x�&�PTTiR���擡����@�.� z�|l�ϧ����EW�"�&�dt���Z>[Kq�Ƌ����ʩY��2/�dt�vg��CoI����P�/j(yz�*Xu��D)�y�tӈs'~w����]`���$�U/�[�(�S<�Y���[� I� �ekX���n����
�
BL�	�?&Es�j5�(|I� ��] ӑ�@�Qd�`L��q�yvR��8[x��wM����C�JXL'l�0K��*!l�_=J�{upʎ��<]$ci~�� �+BT�� v�������;����)A@ 8-Q�m"AN�ɟ���6�=�#W�fD���|�D8q2��C��:��v�`V������d�8�{�?���Z��{�H�w�yE��Gne�Io����q�J&H���#[ˌ~�SIG��|�[�Ny_`�V���Nz�h3�|M�z�~e�
�O������j�b��밁��\�����[=�l�٤���f}i=���$�h�<3h�����^����S���v�����9�"�gTBHR&z�j�\���X�y�H{��W��7��;�`�Eb��_c�)��RY���h>�c	�]/p������g�j6��t�8���N&Y�סP���[,?�*�XkB(��꺣w"!�S�h��=`��w8�A�:-��M�@�(�T� A������pD&����?kB]�L���k.�&��7Yƣu�?-D>�^���W<\��@OӀ5+Z��zf�Y8ϊ[>w���@m�av8�p	P����R����H���n�oc�X挵Q$�|�Ď�
�1�U�M�0��PI����eY�4�1'�v5.k�R��-��r返�v��;� 9�H}����^:�K @�9�+	N�Q�ߑ��py�T5[֙�4	�O�%Zj%�e����69�g���`�L�T�	�*��*���,ݞ�~.�u>O*' 3`�0D6� �ɚ�k��x����:�l�&}�,�{��%�Z��)��;�ߌ�5��m������܎��?��)'kp��d)������O�MIJw鏶W�S�3vlg/��V�[.�C�A��}Xn�6M��}�n������{��%�d�F%b-�Wz~���e�����k;�����p��r�Ӑ%\Q������|��N�cy�^3��J`��>w�'F/v����ܟ��^U�"���H��[<ԉ�:�oSRA���%|	�c�d�@=p�gH�R�J�R��v���sfƨ�=x&��	�%�w�����n�ROjU�{N\x&��(O�6��{i�̅a	�g�#�*��lKc{_�ռ;ɬN��N	HBѼ 0S�"�d5ՙ�q񡏀��h�O���4@XA��Sp�'�J��c�4N�y������A.2�]�:�Es�z]�'GDyϥ7��4���b6^E ��z��=��p���YIw�X'BQ֫2n��0�ƙ�@���q���x�,�0dRJ|�X@]T<5�Ċoc�|[ڹ���XOzw�؉�:�͋��0��a���U�����!ؽ0p�]���F�vU��}{5���G��(���<� �{���t/���j	�dq�����얡�r}���N�L5��g�/�1[���:]2�o��^�^�{����O�n��S2�䯙	x~�E^�����}����h�ҀY�H��t,�}rTA�����2"�sq��Ì��,
��tـ�iB��K	5u��8��R�^�@R��Ը8t�+7i�9��V1~{���t�LHMn��o��D�jA�L�w JL�bz����N�|��s,~�L߀S�RXh��Z-%�ӎ��n`�zSS6knG�v�o�
��D�._�e.�*�l�0��FxuUyh-ٕ���$"L�{:u%&|�do���KX�(,�X�\�0%Q�2�!2�[K��୐��N���u��h���XZ7����D�����7�T�Q�omƊ&�Z���S#x��T4��G�ў#�)pr�cZ0_�0�/|
��{�m��YB�BhT���z��~|�x@�Z
�u�*Iny�1@��t����7��)�E ���ϩ�c���ժ,�1�m:��IJ��M�� ��L�U��U�1 3�@͛Ծ��V�<d�ye�������������L`?�#�O��Bx�L��{^���&������"M;e��P��������km;��	�C2N�_���.��_��c�����␎�E��:�d$9�3��*��S�����"�(������}�
� �>�W�|�,��h���4Q�E���ᓹ�����nN;���]ț��;��\����fzѤ`�~��~���jy����\^YZÅrӗϴ�=<�Y������⒴�֚�hMOj��a)�s�i,��g�%F��g��s����A99Jox��>M�}|���|�V�̉�6�7T4��s2�zJ�%����4�ʛ[A��jyh�m0@:xxB<+�����G4f� ��1Զ��x����}�MGX`�(t�TĤ��N.#!�apN�}�?U�;�
+Y�"1�Xd��W��s3k�傘*}@B)�/�k̼Z�6_�i-ijx����i7��M~P�����s7@�
!�,�*7��9��OU$C�4���j���kFf<���/4��׆DZj�f��+���c1���f�AcAPJ�R�-d6f�C=(�`_�� �/+(���H��\�f�R����-u�K��У����Ү�C�����J�x2n�s�ͻu�0�g�!�}dJ��(�	��O�>ӨW �n�s|Vi�'I���v�ܕ��4�K�vv�4N��74��>���1������A����ƨ
e�3ȟ�6�=pI��#�U���6 ���~͒�"F��KႺ�'v�O'����O4���7��X�p�
lS�BjZ�L�Ė���V�|�J�c͠y�xR�vz[��-����n�t�/V�Ĳ�x�E�P�u#N�/�N�r�IT�fַi���u��O$DX�B��Z�7ÜLأ����k�fh�jJZx[C-PoRe��"ݰ�=��.�}l�׈6��O���I�W?��&�Uzd��N�@a>��qAf����3�"\�2
:yt
'g@4Cj\��y�=PE�(��}*Ӎ��Q<y8����UyU��>^Y`����?�/W�g��D<�d�i�6V5�I �ke&,�����򑜫
u�YL�B?��a��j��"(7� �q����hZQV��`�X�l��v��p8��ĘVw� �l ���l�g��!��a=��̖�*�	`���$�ÛJ@��lB�
� 1������j����)|��8�]?�h´N$i�h9�Qo�ߞ|ϮA���D���������jr���{#+��>�bi{�sAb��x�U�e֪�2���21�B�e�t��'l�%֎l�$&�����Nc[�/���O߆lR�ĖK��Q���l���#��|h7=z�m��+b�QT!�s� �	�4�#��</g�wp��"+�=[������衫1fx���)�D�#�P3�r>��^��e�$O��\��v��4�K����0nT]UR���jp���7��${��M�;�N�`�Ab
&7>������>�&	ָQh��4�(�GgF�86��8t���̭��N!���2��[,Z�*9lLBM�%�w���S��Ϣz��`h�8=�:����(�c�t��Q��0��O��p�4�����?���6�LX�.��=&��lY!r�ui�Y_z٦E��4\�IOng^+Ux"z��V8���v�!�����a�B�p����ˁD��Hy^k��6��**�g�T$�'p|g���Z1�M;kE�k��ڀ�\�@�54Rk''��)��RT���������e� �9F5H������^�J� �H"�Fq@�5�E��l�����T��)֔��	 )%FD����0�}���u6���)��@*g�5��$}�G\��/Yu8Te^� �3�+Y�6Dؘ���-k&�Ǖ
0�f�a�l,A�A� ���{��Č�I)��(ܢ����,?�װ-���C���10���p�	2 M$|���#B��kvgj�U���*C��W���LnxǬ.3�Kӆ�n��,NY��6zd��b�?�zY���B������ԩ��,���a>fp9dhr!��%7���8.^��N�l��[:��~��]�wm6GF���T��:K^P^�C1���|d<��:pɆRQ��` ^�Z5�c�ղ��Zp��4H��JA���Q�ә�H�H�/&�����o�R]���O�DV�`\����P>6��ib����k�$�@^�*�(l�(�_;B�;ĬK�N�H��� K�k"i�W�t@*q,ri���|�J|��O_�X��-�n��'en���C_4�iьT�8�*�A���]Λ3�`������D��V7$u�<Hb��4 W\Z��@���b��$xI��sX�Z�֦^�n&�O0�ݺ�[����JV�S�g�$d����S7c�*�5ؤ{ĥH���ڔ�C�_-f���Kr:Ϡ��]D�|n
���х�,�!@�`0;c�
HTF�h��{P��|r��ʏ�L�<�u�����=�����g��NѲw�5�'�_��,��q�����"X�!�Ҫ&�]����5r\���v���8��)�SMP1�}R~q(��:��7��ӕ��-Y���`tG�Yr�� �bS{�mk_��!�GU�=0㨔�Ҁίi�XU5P	�sV1�-A^�����<��mS+R5���TVb��0Oo�玓n��t7�%�L��JǳjbU�������zs'c����V���X��GZ������o�pQ6f	��Dg�Ŋ�_��_\��.�=l.�hĠ0�Fs�Xy�L�O#�$	�-"�j:P��|�o(vkKS^њ�1�X��0@.2 �j�핝��vG�~X����Lh��c�s�7ߏZ�pD4��a �O�{Q��m�Q��u���΄"Sx�To.�GAq#�Јr2�0��$
`�5�H:�Y}�h�~3�u-~�p@�7���0l�e��'�B��t*�Z�2')y��E��r��������]g,��b�O��QCJ钒��n��j|��p�����1;�@h{v�	��V�n�k����W��L�����W��L��w�u��!����g�֪��5�p C�����z�"�Ô�E䶸��ͺ7G m7�	=�����N�.�|��\ȼc��*�K�}��.�u�e$�sU��}�N��F����Ղ-���)ܸ~ϻ��R��ni��M��d�����E��h���w�qVWnI��3��VB ;�ݗ|�fU\���f���x~����͘�\y��Z>k`r�,��6n'��=ꃦ)�=2��p�hh�'j/����g��eF��l�B)=�X�[T��o���>(�b|�VIԝ��Vi��D����?e4G�2n��Jٻ����J5C|[���vZhC�2@U��B�<|���ؑ��렛�B��!�q��xb����,GӼ�`9T�﬎�
.C�a˯�}T̫�_

� �"odJ��W~��3f����@�@�J��G����ih�^x<� �d����5:Pt����m"�Mg��6,=v�����24�9Z�rU�Q��O���凭�Fޘ<�R./Ϸ���{Z�w����FP���V����AVXP�4=�(}mf�{W(����:?���I��Ї��-r\�7��MԲ�f�-0h&��vغ-q҉��~~�(W��E_�2�Pq��%�K �~տ}?��Lyx(��l��ɋ>.b? �S�s��$ϢH���ed���z4�]�q�S�2�������7�}���P��#U߈ͻ��d
����Z���X�w�&��U����I� O��~�m�}����;�K��:���v�?��&���s���a�6�f�+�5ln��j�/P�'���Ѵ��WF�Ey⾪��4�xm��z�G�-�K}�O���V� '��nA���#i����gN��B��"些�fѾ��8��DD3A�B5[Z������k�b�k�8���[�x�TP��R�t@T̡]�M����.���2�x�E��CW�G�&�G�d�웼��S>Jq�u`�GLf ��I:2�ֽtE_�g�PCe�t�Ԅ�P ��(���*Nƃ����ys����R\tSp���`�:��Z��/�B��ޥ�<X��Q�I[�pe����$��k�
P&L��?\&hdj��(�&� �^�汵���Q�1`��7�gC�v
�8��S��٧�8���_��
l5���0I!"MD=��̱�Lʄl��Y($�=��*�aaB
�r �+P����
��6!)�*?8c�	�c��N(�#��lq��d���K}�Dn����9����-¤��"���=	���ܜ�u{�P�1���q��M	Ų���e[���ͿL���g��&���|�E[�ͷIv��GH����I��ÞL��������|��z�A����$Ԍ8�+����_�F������	Ԋ���=6�����<ZfsM ��UD�ޱH3��3���^z�̜_!�����v�18��pŘ�xTx�rR�TjK</�rq����s{���ʖ"��	!o`ߛ�b�ú=�X��5w�>�	�����H�,C�g���6��0t����H;]NP~��\�Z�,uE�*��B�`��wX��S�:��Փ�`#��84X
:u
��b����(�6�&�t���b�p�co���0?	�D�.�L�����E�&���Y|`gu$�Jz �T�Ky�\V'O	n�+PR�z�38E�1�֪mT���>a�lp?f��&��IY1H4.ֻ��pYՇ�B�g$9]�|^h���1s|M���܆��������4T��'���$��Rk�(og�����l9���oC9B��HP��!^�� ��n�a��Hq��g���Tk�֏U�	r.%�A紛�������ƒ�Z��������*�g蠫��byA�tQ�u�	��1 i'P�&��6���?��k&o7�w��a�ԜK&,�*����x�������}�c�>�yFU�g�w�K�D���!� ��X����`��4�M��O��@���;vb�@V���s�C���x��nSq�Z�U�g��@՛t�d��b#�Zz46�}�p��Z���ڇ
И[pTD�r�z8%��sܮвsoN������k�"�(Rw�d�F�
@� ���+g^KRƑ��e��[<
�!:�B�R��蔛䁇���c�����#8pfN�H�t�J����,<���䝨�?&򒺾�JG�R���O`T�1�c\�j�^r�6�ii��f���3?e����*�)�l��_��s;���mmcH��Z f��"�&�O��qgbw��H�Eg�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�"ڜ4/z^�.&�7'm���n|� �5OA����s���%D��e&�=7<�5�����P ��P%�)��D}~��(�c֡6��B�����M�J�%�VI;����*b2���E��Y �07�G������o�
��y5�&���ps&�==��JWS��f���)��'�|��&<��6R̦�39݁�x�芔� ���ߖ�Q���` ��zR�K��)�d�ǉw_��?bO���~�˳������5@���v��3l����T��D/��E�N�V]@�3e5e��=2�1^N��_@p{5���F����x"���E��+�h�����J��#��	��K��5�x����&3����9@�"x����TɂrD���I��]ⱆlT�ec��N�!�W'_�f�oBY�ޡA��48���CN+�3�H`�q,�0�c7��P�(�X�xD��k�5�*��d\�) `�n�i�q�gz��B�`eU��y����D�g_��� l�_Ʊ���3D��'�U�@I�-��Q�p-�R�52`��M&��ej��K���|�~ȯ�g���9����8��jR*(Ϣ�%|X,�΋���+��G�]�"�ks	k��H2V���B<Rk����:�i��vVs�5DX�m��&�U�*�
Y}c����S�8k^ l[|4�~�)��0��O�,�x�b�h�k�� �tr�n��|���EwˆB4x���>#
n��i����}LS�9�E�ӗ
֡����5�z������J�7���MY�pW�,�kM$@�ǻ$���q��E�|y��"���k,Ƈю�:�ĵ\��Bi�Q�g�dHh�̜>}�.ˀb�J ���D�����m�bKk���Rav�`�ཇ��\���ߚX��%�ۘ�4!*�nD��;�W�xBrw�W��Y�:��%�F���r ��j�#~ ��k�\���:��A��mL���낚�N�p���6V��g١��C�a��"�"���9�H�&��=�Ld�	�O��MaP�)�_W`3�i1�t�;�9<�8e��7��v( px��Z"H��C�`��;��������sL-4a�]V7?"H;��m��A���;9ro1��5�k_����ښ���Q�0�������JpMӮ�����C��/|S�w��L-����Ҫ�*��A�Xu��I�ɞ�5�Z����A��g�����<mPV8�(�%"Q��ݠ����OV��ڣ���V�@�;Z�[h�Ș��'�\��QՍ�����(��,d���_}��%�Y��k��>B�$案� 
�K	�#;}R�B��%O��N9~{W�k��K<�
�<
o�5J�W���d*��Y�pW�0�\����
��2�1̚��4Q�d��	|)�X���>?��@�.��15�vt3�_�;���*��U���O|��Jc$���v�&�T$���
�_�N�W]|�n���l`k&�����=�퐪3�t	i�r+��S|3��ت�ӷpE��ǯ���~@��dr�(׌�;��+t#Zpo�١3��9������gF9�9(P�E��i $Z��̃Q�q ߏ^j�Q=g&�pg���]���Fަ�k�_�0s�X�t���&C��8h��W�7π�X�!�s��D�\ ��W2���Q\M®����Z����Q6���q���S׻�.�M]{;
D����5�'����J���?�L����,�X4�IUu'f�C,.�yO����$�w߼�9+a4�	�������$��.2�Z.N�V���FI��ͼ�R�*���k�Q�鎦�Rs{}��ESv�_����^��q?�<#Y`��u-�	��n����h�`��蘷��Sz6%z�k�4B"Ԟ#M���
��zd�V�O����e揲@�糹B��-�T>Mo�n�Μ�~�~+J�o��d��R�� o{i�w�*dӶ���AY�K.ݥ��5�EXW�ci���[�Y;-U�:9{C͆�DX���y�4ۻ+��ɴ'Z��P����C�Q[��^�AT�����}^C�6P��=uձ����ABC&���ċ]gg(��.lq�fe��}�CUx�Z��m&}&Q�C�*[!���CI%kz����
��I��v��������"t��#�-���>@�uw�^��뿯bn��/fބ$��F{"��Y��o���g^�P�Cl�qpP�p�ė����Y��a�/�0(����a�/f�bR�ƕ��g���a��J�A�������䕅��}JiK5W�ޤV��_E�^�ӠBi2�w�� $����C �l�.��j_�:(d!�'��\��E��9?�|��lAr�r��,��u�)�l�/'�A79�J~��<���#w�:/���p�(���4�}b���� ��A���y����\e%`�$89 �w��.X�� wt�E^`����Q?��z\�[������2����̺Ƕr�Hr&Az�k��fC����e+�~���<�����+A�̧���^:X���Tb�8���"y&sfQ	�E��.�*���x����2��s�f��{�VV|�).�k�;m@��_�<��P �)Dg�{�Ƨ 5 ��0-����U�����ƈ�(ƭʤ�|d�ye� �O���.��U .��'M��&XJu/��������rQG�%x��C��<&�]��T/�h4�����g�6K�	J���m>�<@���JH��x_��LĖS$��ҭ	នN���
��Z̴V�t��cz�'U�{W5�(a�ǣZ��W�ɑ8��c��h��K5�����QQ��Q�,f��墧�\�������J�.�+�a ��X���S�$s������U|�oJ��(�g#>\����JbU�����|kڗ.RS�����:(�q��2�k��[cI�5�6$t�l�n9�_1�qv�T�GM�C�U�H�nK�3L��*�o��g��)/��Xϟ ���KUA���ǝ��\���%Xۏf?��XE�3}�'��L�I�F����?M|%Kl1�RW�k��P�w���?��sD��h������c-.�-��o�ל�۔AQ�V:������0��`U��,�����}ϔ�f�Ti�)Q��{�Q�����_M*5'o�4*��yf� �Knq�x��S�hLB���aaqS���8 8���d�Ĺ׽�-�N���5�g 實%R���x�*�\��#��R��_#��^��Tg����K7��x(�,�<���Et�9Е%��g��l!d�����g��A��1ͼwt�͚X���lN��ב����/�A��~�	h���=c���2�΁~���6�����r`�(��ɵ�_��}��&m�'�,����r��6��(T��M�x{����_�=�}��c���5�4����J�+�	f�}M5PZ�}��0���M�3B������!���z���s!.��`X�?���jw T�}��<�pn(aQM�Z�6a�4�j�ש����yO{���]g�Xy��K�6ա�9HH��g�[=����1jW��ɻ���m���唚�](eJ�g�����x>�"�3v�����b�ˠ]���"B6t/�$�.��[7�m��X|:�~�O��]�.hٛtB|DC��e��97t�<�>�!W�ȸ-�ґ+�D�~�9�	!�����<x����<,�V��y�7Iqb�D�!���Aמ�~惯�����J����৙�>��z�_p��H=�u)�����M�c����"v���v����{S{R4�3�lA��w������▂Ț��� >Rv����,d$,����2N��jqy��Ӥ�..�'�0��ty��:~����QU-�>[��)�����gk5y�{�#WkK�a��Fu�S[DCT�,��8e�O���`72��`�Օ#�XS����)uʥ�@�d;-=-���n+��`��"�$q��[Q��J�7-�1m-^�>�&s�`������$�%?����U�̉9qk)?�J�5��=��(��5YX������7�����2¹�� �����snC��ϓ{�&7&y�&��2c�ʻ��~�ynop�S`ۤ��m���I�ˀ_i'�W�-S�@��L�-�3�b�����ݠȱ����Z(��X��"���� ,�K��Z���gH{�f��eoc���Z"K�ɇ���4_0,ӫ(|aL �s5o [�t��@� z(oI�]*
�y~|� y!.��Na�u_P�nt27,_�I̻��X���ɚ�P_#�$ŕւŘ��ҩ�SU�7�j0S��ћ#/���V�uG?�4����]�> �0!6UJW���fF!o���m�kB|���{��M{ϟ-������4�3X�������� ���;�������@׹τ��#)O��h��p�"�_r[bd��$�B�v��UDZ>
���4�����C����w�;狧ߤ�{1I>ؚ#�5�PQ{o�S�Jw�9���������/ݲ��t�|eC�W͘ ���>*J'b����ᩏ�C�eva*F�|7g��6�6�?v3�� �S�QZ�W��ZZ	� z�LP��m<G�?㥈DN���r��*���Kڥ�Lzށ��
�� �=���d������g�^M+��T�?jX���k"��<x��G��1���Pg��<� ���Ե-��x�4E��q�9&͘����> PQG%S�)�	+���Z�#;3�$ͳ�0�ɟ��Ȟ��T�'\�(�=�Z�t��q�l��Q��o�x�H]��|}���v��8+(B��S]B`*���@Y��VF�x�%1]�)o��p�\B����SDoW�4,�[
��\8W�]�P��_ ��?�Hh��	�� [�;^�A�١�lu��5^�v/�h�w���`�L�?YR
���z��2:5a����$FňmBI�ՐMܔ��['4�����s�<�	�=Ŧ���K$la	Զ��)�J�ª�I������sx>�O[�v|����j��,�."�����:�q����@�>!bv0��[B#�������Yq���Ô��H0�]uԝ䖝��I��ͅ�>k���b����(�J*|Ou�'�~�FbU�o]��nq�w����z*�2�,�/<����g����ݥ�Öw���|�-��|�|6�Q8,j%�����)�d��)B��8���zz?�2�Q� D��p�#s��=j�+-��,�:��s5��s��c�<8�e��qs�+�X���$}�Ƅ<6s�9 �F<d�8�b]����)omӒ�Asd�T-ʏ2��䪜��ۧ��~y�6Ft�`(S6��c�؎�uU>W^?/�t���l]�e��C6"U�t�4ܬ��g^[l�C�T�pnꏢv��/q�Y	���M�0ӝ�'Z��s_��$�sح�^�ݿ{J�f1'w���;p\���JG&�W�V}�o_c19౺g��w���$���!�el�#��%��_�΍d�	@�Gp�Mk9](���l�$V��-�<�S�R�
�{'FG�9$��~����$����\�J��w�/���m�؛Q��|Y� W�v��T�Q���eí$�:1핳..6� a�E������	z��[,M;��iв� ֿ�E\�a�Z��<�HP4�zr5L��@ˌ��+�K��t�^��SD�II�̅�;��{Xd�n�*�ba�Ԧ��y�PfoOE��.Fp������
���s�K����{�M|�.2op{�v@9(_��)�]!{ �x ����Ue��he[����(]�d�yC���z�Ì5U>^B��'�
&�<4/����^���M�6G�n��է<Ĳx].h�/�4|䤁^����p	h3^�K�,<���6�� 2A��Jݖ��\���	�7�N� ۨW�Z*!z�l��_*��̡{{�ӨF8ǁ���뇑�Ǎ�1rh���5J����:ܽ�9�
z��w��������VJQ"	+]�5�l��L`��0�z���O�e8J��p��|\�G��(���"����'�LBM�����+q(5rq�p2����jdI=�6BF�����g�_��yq��ٶ%�C8�Q¦�K��wL��s�����=��!/�.�Xm*�����Ks��߶��5��\O��%vdfPX���}Q����4*I��$g�����%i3�����	�+��k�����]��T������c�p��\-�* �� 1�|IQ5:?�EU��2$��p��l�A]ܞ�+.}�zif��nǇ&VٙnF؞�7�f*�{��3����`f<`�K��x��ΗF��T��a�%���V8n�$��|����K�Ο�t��#3���R&�T�V�jh��Ms��&TwR�5Z_�g^Sh�g����)�1-���,��	�]@�tRrT���g�yl�?��Hf���;A��q�+s����⽪��S<�F��Z�e�{$!e�f�c���rum��;���	B�ƾ����~��#�aèѩ��U��q�M������O�z-���[�-6�R�G�b�cXC�0m��>�P���)��6+��h0�qtbb%.Ǳ.�tF+{hr�����Q������EL��@�nt�l�J�LU�aiFN��-%���w��3�3�Χ �[�[W���c%ؤd�9HZ�z��/�(�I�G�]�p�<��2�cv	_�E�8�^dt�ĳ=E~~ϣZpؔڕ�%xP�a�3����9���|=�VFۍ	�o�6��8"�a�qʭ��/jKG���{�H$�X1E��d�_*�ni&x�YQ��ɢв�X�$Z��ɡ�9�6�>�s��~!@:�3����>
6�tJÌ8_B���.��8�~]�3c֥�x�&��at�A��y_��g��Pd��J+��h������ῴ�73x�5�vjQ��b2��4��٥�Dj�)�wފ�v��Cr P�2i�Q��#}DA����U�Yέ�֡j)�����Q�j_BY�rd�,��q:�1����N�1��欚G,M$Y�iٞ� �+�:��w`�3���4����������e���]@)���3�y3�D��:#���PD����ƅNd�F@�Pe�dҚ٬1[὚�2P{r�^�Th�?Mkߕ�޷bt����h�:���N�*W��b�K"�:��>chp���l��9�HFx�8��t|��gZ���ҙ�&��"�e`PBN��b��4��C>M�c��`�֛��n��%VN�QF3A�`ó�� ب�9�Ix�}��b ����p���Ïu�h^�V�3�F ���7:Tp�AO2�]R�p�u��:��G��PF���O����|�l0�/g3� �r���[\���}d=�Oa7T���`�]��}�)r_�Ꙫ\�t��o��:�)��1Ҷ��m��))\4nQ>���.�z������.SW�0m��ȐtC��'Hc��,).���_��U�б��a�z4o� ^��M5����}h?�L�j��K#ݥ8��d�ٯTծP�L�8�=�j;lϫP�|������5:�������L�	T�H;��߻�R����W��iSJ�V��5�^�z�5��~c�S0�c*a���Zk���l$�5�K2"}0Ύ�O�<OxQ��k���=q�W�g|��E�Ɇ��Zhx#����{
b�i^y �f��#��E���
$t\ξEn#]��i^Ҷ��7�V��vO����,%��M��Mp�7$w�#q�c��<��1��>�:,/����m1_��3��:���m���C�V>��-��8�J�*��gԊ<d��Dk�A��{�ƷT��&������Ӯ�	X�3%s�i�=Z�5�3��+���DBr �Iєu�:jN��xV�0QrI�i�td~��h�[���:�w��7PL�[�˫>��K��<�I��}�8ي�LMa
a�"9�y�v=�9LI&/��z�y��(�O���ay�令��3V_���;�ȓ<a8���� �O��H>!��饴;@�t�J����L6C&;��V�4gH�;ym0�ڙـ9;���.$�tg��*���|纰��}���uR�p�$��7���ﴱQ�SN\(�S
��S�����p�Aεƀ�C���Q����-벡��`��mز�V!4Y�.��2���t��X�2D���𔤧c;V�O�;c�5h&6��Y�,����Q^VA�A��(y������g�}��H��a� �Ռ�B����Q\j
����}{�B�=0O"�N�88WGw���
�֏o���Ъ�@�zd�r���!�WL�\����}$�*1�k@�}GVdU�J	֘��yզ1'����7�]149v�bU��ǂ.�9:�I^^��8��S%��#�W�����4�B���i���]e�{wgj�|�&5lE�i=Y���*	؆�r�BS���HOD�h�Ʒ�h_�vX¿���@��]r�<ו@ń�y3#���B��~C�u*�0�\�½P��뙒�?Z��8��&q�a\^��=��&��G���J�����)�kG���+�s3�Pt��q&,P����8�/uW���$��!�AJs���%�s�@F����OM�`"�7�v�B�}��>-�7�q� x��@N���M�F!StB%W���':5��a9*گܜ?��0����u:�4b�U��?'�j,���y8%ٸ��s�ܽ�8��]@󅙎�~��CmR���ۣ���Cs�Vs+���-����B	���t���1`��d-S(��d�7���%�H�i�qz�r�Y9BҢ:#�Y����z�h��M?�V➏bSQ��B�&3��U�T�7a�
��8t��.XL����U��� �s$i��*ĳ���WA	�G.�������vW�S^i�=T�N�;�5$��� C}�D6�)n��k��C�='
!lP�h��֛C�$B�y�-(TG��m2�^�ܼPx�u���⏕A��u���,w�$��������Z�@��)xU�b�����;��z[�YE8��%^�������IIvF0���ёDb��3�� E�ݐ����u'�^QР�_7��p�U�E���"��i���t�~x^m��CJ�p ���t$�A={Y[B��0��W�9��ߚO��EE����J��U�8���W��_�er�JW��4V�MC_�-���I��Ew>q�$i�P���l�ń�w�%_�=d�J��Y����
�9����\l�%"4����A�%���;'�6�9���~���쪅��ܰ���e��� n��<���-�]�N� i'@�oqM�'��Ce��$荢�'q�.�  '�jE���2U��z�[~�+�b�Ѳ�"����g�����f��H"�z�J���L�N!�+�lԆ6��Cd���cm�W<��X�w�����b3��Ը&�y�Z�f��E�0P.Xi,�@���k�+����s�}�o{���|�k�.DZ���@��_��� ��)�m{��8 �P���'�`�U��P�:s�����z��,G�yN��I����uU�9^��'��&G�/HNu�0t'�_qAG_�g��l-���P<֬A]��/���4N}��pM����	����y<�	����4βj��r��j�X�	�i�N���ۺ5�Z|�$�B��\���c�{�;���ۧ�S+���虴�Nsh�m�5\FI�H�罢պ����9W�ł�E�A^Jc��+������؂h��Թ�������K�x�J�o�H\iA��B����m�,8/�޴A���p飊L(��Sq�J�2x����I���6�*2�Y���n_�Nq&�<����CJs�����KL�RL����*)�=�FVq�/~p�X��L�NK�Tб��G�\��%&�f�C�X�8x}��w�no4I�18�6��ﱮ%�f��b���60� ά�Z������f�Z@�Ğ?lc�j�)�-I������m�QGE����@��;/�B��,��#��e��}f��L�����+���Z��I�@*�sѳ�ִ^L�fNO�K��xC���]7�f&�a!P&�f�8@���c�i�H��_4�q����=�_SkR�囱(q�z�2������3R�r_�'y^��g��h�������%,D�/�#tdpr����g��l�\��Z����ARf.}�t6����g�h孀�Υ��/B�<A�����������A���{u���1q�n�IࠨN�"��(�ۡ�e��84Ǡ>�mnF/,���"#!6d�M(�5M�E�q�ӂ-�c�*����ﺧ����.�ƹ��-`nP��B�-����U��Y8�3�?�s<���'�*�8ԇD!޲�`㹩Oj�j'b�-�ρ쯽n��9ML#�6��r���,=�^�{������`��y|6�07/�Hn��g�����f�1���y����թ6}�J��]����g6���.�(+"���e^:�PQ\�P��]�Y�"��/��{.>2o7?�+���8�OY!P��r�$��D�-�e>I�7$��<�IA�ѥ0�h4�����A<�D�;��@�ֹ���Z� ��v��b�b�T�VaMg��bJ�p��@e���H-��_3���łχOQ��fQ�>���*z�p�-=UԖ�b3���ţ��$�Ҭ�5�z�4Q��+L�R��43QQ�Ő򑊬�ȗ����2�x��Q_ ��QR�4��A(�d�V�����[�����(�D�#�4�Z091#y�~_:̮W�l�xQJ�>��٦8�wguy�B��7{K�X���A)S�'TX�$|���S�Y�7�l`d|��e}SL�U��� �p��d끰-��n��{`b&��P��=��Qb	���[���5�-e���cy�l��{b�������y�
�9��k���Bg5g�Og�kKt�Y$R�yy���q�����`�9l�̹���Ǡn���C"����d&�y�����2�?��n�.��n_�S� �v�������{G�iד��݅�@�������k��֍>^�a�Q��zZ�
��6r"[��%{��PZq�mg���fk�o���c~"��j�bh�4��[�p|#a�#�o��ut��!�K� *�QI�x]
1�|k��!���S��%����7ܓ=I|����v:᚟]~#�7 $u�/�2�L�����М礬0h�K�#��Ш���u��k4L�a��i>�_�0�̥U��W i!rY�>�]k��!�XV��{~(�Ot�ί�B��NsXb��������T;>;Nz{�P��P���i2�ܧ�b)���hJl���r�<�����v��U��k>���� ������ʃ��#6�hp�W�S�+J�>�#�:�P�+o����}�90�:�PW�e���b�6�$�~e��&�B���w���@*�I ��]��8aӲ��e&�*��756dsN?&���'\��WC�
a��z�L ��m�3d?�(D��ӑ"���VpX;�UîL*���v��ް���2'���3c]	��>^���2djG`�PN?�Qu1���������n�׫M� b)M�����1z|xsE>�Mm��H�E��  (c%����K���ZUҟ;�y��c-��6��N9螈7e��N�(��4Z���[�l/�>�r���K��iѧ, *�Ăf���8��}�JB���1�wYk�jF2ˇ%��A�oEMs�mƟkS����X[��A\诅$g�D L�?6=Ph9
.	I��[����/����l%�f5�v�Lh�}����!��Y��Iࣃ��5?X�:~X�k.�q����D���[�'�1y�Ĕes���`$=uӸ6���<�a�\�K.R��n�:::�����jD�#뗍�#v,�Eםl�qw .��'�S?�:1�#Ó�y�v�Nޭ��h4�XKX��9���bQ�ãɎf(�0����&�v}8�&�*�����MB�ѡ�
z
I���Lr�}3eBv�O�%HNJ��W�|�؜s�
Q^�ou��Z��~�d~b�j��W��9\b�n�	褂1}�E�
d����kQ
�\w��V2�A�XsZ���B���D�����cߑش`�GX�մ�����EdWC`������ߞ�Z�}�1���p�
%�K��z�6�m{#�.F�~\2�]RRvF����z���N��}T��a�
`sl��є�F]Oh+	�jX���w;�q��RxA|�����t3�4�mh�t��#�"Ś�x2OfT��W�H��J��m��2��j?6�>�̈G�x�NH��@�_cN�+A���:&T���u�DG��L:��z؂�D!	���VT5$S����*w��RҮ���PU!H�*fO_~�or�6���<��g2!���r��#��'��߅6�}-�� :��.�t�M�K��$Չ@�������-�4�HS����b<��C��, ���b��y⳦����<0](�b�sǫk�t������p;�豯�`���^���@�m�V��J
�h�lB�a�ENO��-�v��w���m-$�!8�[�b���c_ud.~P����z�(5�0G@O�p�]E�j�c�@R迳��R�t�i=��~Io3p��̕�_�!	aX,�ʟ�ޫ{��=
5LU3�Q���"f6� �ۇ�g��/d�1�EW,{g-$�ǥE�g�duaai�,�S9��/�d�.$v0ɛ�7�po��1t~ە��-����6d�"�F�=B�o�hO(�d�:~=�c
=ِ�ǯjo����yY?�ˡ�MP�2����)S�䍎�[�h��	��/��j�q��^w2s���W#jO��w�{�v�3�J� ��2#W�����D{м�I�̌�c9��8n��`�7|rу)�d.Y!!?/�+�+_�1��/����P��f�_G&vYY���P"+Fy2�qv�3�j�4$R����
�����7�@�=*�-Wz3��l���_�D�e*�BMN���@�I�e�������1�ޚ�rv{l&Mkҹ*��O��ޱ�9�(�@h(EY�Na��$�Q� UK�Km�`��b��1��}�Y9��Xx�#���ƀ�i����������te��Nb���y��}"�9σ�����G���g4�!��Nn�,���Z����$�Ti�gN��y4q����CK���ʩS#�T��O�`�2�s�G�7�P`�z)�.aS_v��L���C��dl�-&�n�7`�� �d�PϗQՍ��nϛ���-�x����L�cI��IJ/Ź�HOκr����1��z7k̨���5Xz���~VY�|올���z����#Q���m��$��:�jn�b��v�i�6&���)"2�]ػ�<���2
n��{SC�	h=��=`��>i�n	��b@��Y��h��+��րȴ���P�:ZʞV�{L�".�դ�����Zd��gK��f�go&�0���H"Γ���j�4����N,!|d�����o��t4M��� ]2�I8�a
$��|��!���5�M�� �7�PI�����z�9��RGp#�WO$�B�EĻ�BE����ȡ0V
�����#�h\�9��uʑ�4�����V>��50$U��T³O�!�Q��Jk%R���{�n(�Ϣ\@�b������X��늙����J���o;Ag��u��:�|޶��)Ҕ�h}{�e��r�"��������Tv�.�Ug��>�,���$�6�������Odg�j*���t>�I@#��AP��Bo�[�M��9���c,���5�$�W�9e�#F�5�����y�&*�Ɖ��d�u��J6e�+*�R�7j�76x�?9���C%J��D�Wv<���(����LST2m�;�?�&XDqXU����� (��H�1L}���)�:��W������%��5)�^{^���W՗j�T�c��Ļ�|���x����מ�� �o̡7�b�D��x�&�E*��@��z83 S!%��;���t�e�Z(-;/�������מ;NF��;�("�Z�Q����&l���v�Y�r`ի�k�?p�7�����n8ȸ��BO�����Y�FE~�%T��Pox�n��qkƒ�SG{�җ�][���\[�Q�
����g �f&?)ih�"b	�Ю[�g��d�9�\�6lX�5�[v�,Mh9�b����ZYu!.�[vȣ���5����-��I�6���pfB��'|�W%�s��b=(�wI[�n!a�u��~�U鍑�- f��U����6���r��v�_~�мR���.�뇻��K:�/2æRN�a!v�m[%[�,旧#�
�Ӫ0q0bN�WFHSgxԀO:��eZތ}��A���~�b�a��Km9*�<=�9���b�~�o`�+n��w��$�.��*'�#���<]}��j��ђ�N�w�|����U_:�Q{�]Ș��(�)W����� [j�Z�?�iQ�I�'�c#v����Z+���,��4��A����:��\�pj8�����l+�h���_}C� <�|9�F���8��]r����)�虒!�sG�YO ��2����L�H�Tߞ��`]�ƒ"���w)���~cC�-I�pEq�߫���*�F1���p�$����z�XQ�:꧑���~i�]�i<F&П��1��������Mc
��B��t����F�Y+��X�cwh�K����A��*�o��d��{��!�$m�v����+�����L>2\�͑H3����7r�mL02ݖ7?ߘ�>-�yGՀ��ӣ���I_Py{�ɰ��?TP�u=�,G%�L�"��6���oZ�!��G�L JT���O�]����m�׮a̠z��!��Df|���dI�riJ��ҽ3�ճ���Y��%����Z߲g0J��mj��;/E��s�M��#���jԼ�p�M-t���UN��n��b��XC�Oyչ�Κ�M��F3.��pj��0
�kbi�ǘDt�-"�c��>��yo<����������@�{���]J7/�9�9at�cN\�-L��v5w�������N��[�*��uO�cldOd�NDa����*&(¡�Gm�[pQ��bI�c��X�l�n�e5t���=�:~v��p_�ٕP��Ma�t���h�!=�\��L��F;�C�o�ʴ�J/Q+��һ){�
�$_��E&LgH|��i-�x�@( �V۲��N$�J�蘶}|���s~(m��oZ���6�XE���B���u����c~dc��<�? ������ȵ�y��dˮ�)P��YQ�Q��$��q���8ؾ�e��Nj�H��0�2�W ���临j|2Dwe��vz��b w�2p"֗y͒D���v�|���B����������Q ;Y�0q\������1��
��X Z�QtG�Y���C.�+��ޓl3�5�4�P����9��n�,�2�O@�^$ᚑ�3<������?D��G	�N�@��eY6���'K1��%�/�{Yl)�n�����â��p�5�fhՈ?��\��׬�S�Kɝ��-}������T�*g�9�rxѣb�;D���(>��.��_��voe��N��+�{���
�jf۾��n`;�ؠ<���N��'3(>`�)�</^�=�I�:J��� 'W�w0���u��V���5�ͺͅqI:��=�h�l����y��u��:�4�GD�(F30�O�\9УTm7`Cgħ�mf����\=r�}��OTg�T�)�g�%���Q)91^�@�,\w��f�����%84�c�T#�)��n��n�a%z�/2��U�T���L�W���S=�𽱓g�#�<��R�U������A��`P�}��5"����ʻ���j��K
.��lf|��������Ȫ���8�#jB��ϒX�|H�n���ļ�^�7�8�Mt�f�	[M�H"͢����R[�-�ދi�d�Vc"�54C����+��E��;Zc��g�C��k���lKW�ҷ��0��O���x����k�%��d=q�^_|��Eg*k�2��x���.b�
^��i�n��me�
pEz��
�T{���d�j ����ҽS�7{(��=^��`��,�l�M_���"$�,rq��}�������d�,�x|�~����G��ͱ�A���TO��
�>m/��pC�J��-�4j�ԱJ�;�k����B6<���8�X)�L�\���!X��O%z��$Q��2H�t�V�+U`�Wcrgs�ѻ��:qr�{<��C�r�LZD�~�ԇ[L?�41:�A�����L�t$�r�(���`Py���Ό���ّ�3��a�P "��2��:�9���&v<�w4����O}.�a@u��Oz,3�ꁲ5;ޚ�<�Si�;��H�jm����h�����O��N��J-y����ޘ���*bnSCZ��������붦�5
��'0O�bN�[��t2��H����~i?�sX��{R�h@%���J�����o(ay�.N��-�����w���t�Y[�]�z��cITd ��FC��	(�P2G2B�p��g�.cb�6���J�CtJ7=1��~;4�p�2��U�d	aJ��щ��� 5=��Gʓ�9�K>��-���G\ʙ�/�( ��i�{Y}�$�NtE+���S�Ji�o�����Yg�V�Z$F��U^�"�ߕH~x1ߟ�h�!�6V���x��B�)O��
�V�d~I1*c|�h�d�E�\Nu�-@�yˢ��Ss�P�:,6�y�_�&�����MXa�#ٷ��Z�j=���PQ�2��m.3*�	�jAnw�\�v�k�@� ��+2U�͗�vD-O��;	��V��G�'VRE�)��ѵe����Y�1�!�2�]d�1M���������NG��2Y�T��I�+x����sI3�N4�E�|m�\q�QÉ�8@g៦�3��^����WD(�l	�NГU@�3e^��҆��1�׾���o{�0w�Èҫ��߁���#zg���,h�њ��8��DP���K��t��D��3m�o%?�o09�dhxV���`C�[���9��HS���e�JHN��'� z)�/1�+���_@1��}}��5N��3��k`�Ҭ���l�2I䍓���0 ]OA�\a1�`a�u���Ԩ2֐͊��:@Q陭M��)�����u�p�:���G���F8�O|�!��fa��g�{��߳P�7\��}�bO���T&6��L!��F)^.��Wi\ܮ�k��&�0�j4ƶ��b�D�)W�n���Ɣ8z��i�����x�m���|��{�F4�����ȂJ��8�U�x�	`E�f��%���l5'f̢iQSj��?K�nCݑ�ܢ�l�@���É��a�8'�j'lv�N<|m7�����!P~�<�P��O��L��	@;0H�w��˒2R I��C�ai�ɖV(65y�p��f!�I�jf�ֿ�kcϣ�H��k�u�l��1�ύ�#@0��
OfI�xk�����ky�O��B�C=e|!��E�$����x銝3f�
S�iʇ��R�ڳ��7E�7a
���H�W���zO��GҢ�U7 \�b5�%#K,��M�C\��$�/�q�R��w{J��p���z,O�у���Y����E�&+Z����/��>2B��ծ�J�]C��B����5��� k>K3�g�b���3�Y��Q�8ӚYX��b%_O��ƭ!+^�9�+������jr��� �x:V2` �n��ur� �n�~l� ���:���XE�L���7� �pq�e��5 ��c	�v����a�G""��s�b�9��}&��W��#O
�ae���K�3�
�)�;�q<����O��N�� ����3�H*�8�U�Z;,�����ō�NJL� 
'; V��/H�[m���څ�/9��������Ђ
d�OB禲{���g�a9p��q��O�!����tS�|l�?:�"�!�~:��_�A����h�ɳ�w�L{�E�\E�L mD�xV�i�����
M�gK䛤�3��%�����2IV��;ϼ�h}·�����hQ�E��-v(����ۗ�
-	}���嫰��S���Bo����?
� �0s�}gP�BZ��O�+�N.�cW3��؀��
��oY*��绬�Pd�D�N�W86P\FZO�m� �ˏ1�b_��TdA	qu]��I��\�������1 B�v)�f�n	���&s&�4��$Eϣ�F��E�o���Ok�����N���_]Q��4>���&�DB�O�=Ũx���S	D�Fr ��S�`l�4�#�����zĶ�ɿt��@�uvr�p�f~��L#���.\���>Q�a��Ĝ\/��P�y�~��Z4���ؐ�q�^�Mt=Q�s&�RƇ���@��[��k3$��s�"t�{&� ܓ8}��W�*���W!ATs����E��,*�+��M��0���U�.�8��E�P�q:7i��Df�!:7Mr�I� ��>g��'&z9��qڛ�?���ƿ��r.4N��U��9'��,c�;y$�s�zY��^��C4�f��韊ƀä����/.��Q8��mF�X#�"�TR�W^ۈz�܆(��{�s���Z������)��Ñ�ѳ�`��-x���V���YU����Q�~~z�z٠�B��$#ɵ�(z?��熛@�G[!�B��Y����TS���#�,����s�&��/���&�'�� ��	i	*���W2�AN� .rJ�m��7�W\wTi ��w�;���/D]Cb��D�Yb�N��0�����'P/���� C��E����3rT�*��V^�o>P�7u�-�t�Aw��������.~=�o���Wﻧ�s���jx�%��BXd���X��[�V��Wo%`�b�}3��? cI�.��j�$��ɕ��eW?�o�"XZ�ӂku��Q^v^�$(�մV��%�Qe�"��C������o^���C� apecK�y�-��Y�Y��˫��u0]*�^�2��f�wa�J호���V"J��f��ٮ�7`�R�o��K�J"WC��V�_�1���a>��w'�$�-:����lLa�����_gV dV�#�~�Y�9T����Z�l�)�g�A��?ݪu��AQ;']֭9�~����Ȋ�\e���I��E��$�ؒʉ�S�8 B-����fnŘ+�ke�ä$���3�.{ ̺ESqֲ�jt�8z1.*[CQx����fd�:f����Kg0H��Ez��&��k���+��E�+����2�����ܯZ��vX{�ơ!yb87��]�Vy�!f�EY.}�#�O��Ц���݂s@��򴽲{���|@I�.i��R�@0�V_�����<)91�{w�2 j����%d:U]�?N�K�����2?y�H��$��ã#3U5��R'�Ս&M^�/-N`��pr���G$,d�ׯ��� <{D]�0/��j4�.���/����B	_�w�"�~<�v}�?�$Η�����(���#z	���N�"�_w+Z�7�'V��x�����{�L1�=!�X����}�-�@���|h>	5�'���Q��e��q �:%Z�)��z�B�0�J���+t���Gz�m���yz����~��4��JА<���\�)n��7��:^��q�z��G��9����jq(L�q�}2}&?�<mOI�q56�ҩF�Y�C�o_��uq��_���OC��=��K1��L=v1��������/�pX$�F��|&K�!�6�J�l�d\fOt%mb�f�iX�"�}��r�SV�I7�s�[�ȓ�j�%`8B�g�����{�Eap�?�R�"���0�����Wc�:�j��-����l0��Ql#��\e��)79�GyhT��ؠ��J�} +f�&aǞ]�ِ����.���**f̳�Q/���!fs׉K�"�x��'�/��9�af�}�K`8��[�@��..܍B8�v�C�i%��/�R�J��r���S�dڍ�IR�Cr_x�^�GgqkR�6��}���",��:�45t	���g��lV��������A���3=t�M��Lc�2�����w/~A�i��١^:���Z���a�`��V�[�3?��L�'��(c�ɪ��7�âm�!�,g(���[�6i)�(��cM��պV X��͂R�_c�_g�J�~��Pǟ�����X�PO���R5�Д���3����̾��������!��`�թ�aKj,�����1�$n��Mс�66�Z�߅�����c3K{=�w�Rb��҈����6��H��WHӫg��ݐ*us1_w�^�d2����ϔ�&]=�؞����X�b�m��"�Ɂ��a�us���]褐"���/7�.���7$���7��]�5O	��CS�)��D���e���7	s.<31���}a�-"]��F^�D:�J�֞95��AR��p�'��A_iVf���Wb������v	�m�V�$�$�e�ό�L�as���<��Dhp#i=z�S�'�>�b����Z�w��z�$�0��>R	$�3����튱���>��wc��E� <WRٵ·�d9��0���pZ�_ް�r!��ɬ��YlP0���y�q#:���`QJ��>��)^��]��g���y�a��̋KL���;,�S���T�t���L�����W7��`	����S1��^"t����d��-���n��W`灅�$��"�aQ�������-s���ۗR���k���X��G�Z�@����_n�̞`�k�H0�5�D	LQ]���Y-���>�U�L@�˦�Y���~?���U�L�n��py�;��&�L(�{
�2X.o��+��o�nDݰS��Ā�c'����� P�i�h��K�@!�!k6̨�y��>�֒{�e���b�Z����mY"�E]gR�`Zv?g�T-f��Mo�x����R" 	݇'�v4t��`xB|��g�h^eo��<tFR��p�� ��gI
h6
6�|�!#��m���n�C�$7���I�
���l���Ç#�fV$��+�WPʻU��h�i��0�n�ѐ��#�)��K�cuϡ4�Q�r�X>��r0v��U?'��!��=�c�k������Z.���$2�����ɼUX�����_�����;S_��o����N�4�,��)$hhA��7�r\�7&	�7J&v���Uy|�>�1��������҆�*S'ጇ�<OO���A>ۀ�#F��PfHMo�)l����9u3��5��-݇`���E	eX)�G��UQ����*� ۉ*��\-�wP�e��6*�
7��6���?�t�U��&�W��o[����L�z�m1,?x)�D��!�G�П�e�C��Z*L�����ޕҙ���I��V_"�R|,�^��_WjM)��5y����K�����EѸ� �װ: ,R��	����x�Y\Ec��2��ͭ�!J�_ ��~%HQW���� �qZz�x;�����lǒ�b������x�����(4-�Z�Jȿ �l�l���S��j��= :����I�����W8�]ǁ�7�B����*�Y��F_�%f8f	o
�:�qk�Ƥ6�S�1K�)9'[�������u�!�!̀��H���x	����Ri�<�
��o�O����'bB�X�d�M�	&�N��ۏ;�Z�
�W�0�6V�,LC{�.��m-ǈ������]�9�(b�hHJ5��P�=�ܽ7�R�и�jI��ӿ��s��`�J��r+��̽Bϔ��'���ώAx?���d١J }�z\����/��j��š�����i�����(|:q<��2��l!/I�6�RGv���s9n_��=q��!�,UC���mO�KacELm,��/1k�2���`�/�RXT����Kf��f����yU\��z%�ڠf$��X�f�}���f@Igò������V%��[�O���h��u[#�o�d�R[��<�51��3~�c4�a�ٴ�����D��LP�ς?�c�"�w1��y�C�����)Ͽ9P��c�?���2���v3���܅���#@xϼ���Y�!��S`Z�A��Rj����?�J�>��njh�MJ
6#�)�l�h����0Zv{���_pv�����Rw6�#���)H �.go�u����1lB��nE'ջ֔�g]j�Ҟ�+�����z�"-�V�7���b(�ˢ��]=�"�<�/��.�D�7�������J�O���p�E���tD0�e���7���<��Z��`~ȺQ�O�����D�/�钁��Kڝ�,�Ξ�#��� n�\V3�����b��z�c��ü*�Z̭���_�=q�Ym ��>��u�뼞Np]�=ge;���ŏ�k����v�������:���R�z�3�6��"�d�~#헫�W���ğRZ3 ��RƩ���? dfX��9�����lNg��|�T�F��0�z-y,�:���~�wQW�c>����%Jgm��y3�P���fK���HZS�sT*��R��Q��Q37�c`v V%lS�gث�����Zd=a0-%�n��p`t}������Q4�ɺ��ӛGM-��!�N�"m����D�,��Nκ����M/��1�k�?;T[y5�"���|mY7G����y�������칋ځ�^R���rcn�ϕɭ�hs�&�=ٳ��2e��Fy� ��n1V�Sbỳ�!�~!�ȍw�i)�B�o�@j���[�5wA�*�F�_f�s�7��4%ZI�����F"m���b���8ZC�zg
��f�K�o����5{'"YB��ׅ4���-][|#)��u�JoBp�t��1�]�2 |N�I7D�
(o|}�!0�k�����~�0��7.g�I��ڢ��$���#`�$G��DwQ��x�V�F�0D�ѝ#l#q��9�u	�#4����[>���0�eULT�2!�^��Pc�kD*������M���a4l��h�v[QX4'��؄U��|���@�; 2��b���������y-�)Ah�9ױd��r�\/�oF�D�v1kU��B>�iv�6 L�#~����߃�����F�������>�U�#�k�P� ocsw�<9�$ŋ�+�73�t�Y�v�	e���x ���:���*����wv�k��=�e�T>*�H7)��6�aw?��9���y���W��S�����^�LU�m>Tw?%S�D�0�4���,P�|��'Y�L<�����BY��V���<6�4�A�^����t�jZ�}��\�#V�����3&� �}G% t]���h8���pxE��EP�d��v��{ T8 Nn%Um0�U>�m�Zg�;5;��������`Qy��Q�i�(�}XZ������ l���U���1�4�J�ۧ��}��+5��Ġ8-2/���B�g�CЊY�5�F�J%�`S�$o������ �q�S���6IE[L��\��_˂��� �2,?c(hK�
	��p[����i��YklwaL5���v��h�Ov��8���Y�3�Ի���>5��B��0o9��/��g3����'6Q?�V��s�=Y�W=�KB�;���a�q?���錙�(%����!���ߪ�Ѫ|v>+������e�.�bĻe�:��g�%Q9���kv�[D=>�+̧f�ВLq�;���,H�$iW�Sԟ�E����k��� ���Դb8~��;*>ut�y��-�b�BdoĲns�w�z��Q�*f���.�
<\P%�I0E��_�����wA��|sg��>|�~؀Qzr�:���o)�7H]�_�6ޙ��?���Q�#��{#5���?p+o-J,78��5�������>m��8J$��s
�+��.�}��<8��{HkF���8�Þ]��o�QP()�.��Q3�sf�N����Mצ����6\�:�`���a�/��2�ѫ�Cl�4�/n�� �**>���1"�;p��!�ל3z������͑:>z~�+�]^}FeOI��{�.��NX�tT(
l���(˕��WF�t+XkwG���q�A�������ߖ���%�@�Nm�����.۠�ulŦ��2��*����Ԯ��V�/mK(X2��U?���>���G��i�Z���̅�_o���P��;�T�u܀-G�	L�#�u)f؎,�!���+�AT����Ǣ�)����Eu��%��6�!Ԁ�f[�;�#*�rC�Q�z�sqܮ���UQ��0Bߑ�	�������J���M)	������m��7�k\��}5:t��Wz�w��d�DȖ�#(h��R3�����Z�Ň���pV�H��jWb-A���;씌��K���¼ݰn{[Ϫ�@�?�.�!
�mYyp.�=X����og���+�å�U��Z��wÉ��8R�3�@��S�+������"�n�W7 Z�*R�����ʳd�E���Ѭe������аƤ�'��7K 0��y]�F:����}'Q�>N��|:Z;�wg~vydd����K*�����mSNe�T�k�b��b/"�7:1`�.�S���|Wϥsm�dN�-V Xn��d`�� ��89�q&Qvj��\��$W�-Ѳ��iH����y���T�xg���޸���k�XmŞ�5J����P��cYˢ�� r�B�����7	��<�W��j�n��Ϧ\��h&���Y�2�9���ż�ځn"��Ss���9b���}���]�i�z�� I@;ʦ�7F�F��[��ְ���p���\Z�`���TB"^cy͕��Z���g{^�fN[oVr���"�����n�4�m��~��|��֝b�o��td�(�N� �f,Ih^�
T��|�	 !��Ac�ȟ�!��7? �I?,�+Ĵ�o��C�#ڵ$yy�5Ի��N����
)a0�p\�.��#"z�iܵu��74�c����a>�V�0T� U�.��1�!�B�A�kUF1����.��"�ΒQ��'��XL���C�������;qWO��k3C&׬ �J�V)#�h�WI��sJr.C�� ����v⠇U���>����G�?�T�^��F7�K��%�������*>�7�#�P�.*o���}xw9�n���v.O�e�����e���e���3E���Hw*=�&�H�l���_�e� *307���6G$
?i�$�s�����W���ͻm��	�L�j�m�(?ֈVD�  �%;��=t#3"h�x�tL��8�Y�N���Ղ�������ڈ�^ ��K~j됽��E������L�DLܸ1�+��5! ��g/��t�:x_�EAh��DZ�yh� ��%�4Ò���>�dZX��;Fcp�&C�����ˏ�k����(R��Z��S��B�l�����f��N����o�`�g�w��p18>\Ձ@
WB3�@���YN �Fu0%��D�Vo�O4�ϻ��Sw���[���\��E9'�� �?Yוh��&	,][�y���+��(Sl�.5��v��hB/���t\�?-�Y��L�����5��
�]�[y� �U<z搠���i�'G Sԇ/ys��2��=X�y��	a�cנ��9��E�]�,#'����f�F���v/~� ���48.՛���<�:���T�đL�v�U�[Uo��\� �S`���(q`CÇQ�H���H��԰�	�0޼�`�q�����Mb����{W*/�������b(��o��	n�w�7��^�\*W��?YL<���ۚmȄ1G��D�=w�I|D�[�/����Q�#�8���>)����0��ފX?�mdQ
��W��#�mǢ��*+ �_,8g�&�y���yp�p�8��y��+��߰�n�}sq�<Itg�#,F��8/];na�\U)°v�B�"sw4�:��b�:��]�x���f�`��@�R����p��TC��c젛��l���w��ZЍ1p�D�[�zQ�j�����~��]/FV.o�V]�O�3�I����C
��T��Z���qF��+&@�XGk�w������0A{U�ZU0�]3�:e�QP�m�������� '��7h"2��5�x^�Ű��g&�m|j�2�?�>]�G@���+����_�];�3m�O��T�U�umb�G5';L�j��f�k؟n_!�h#�|��T2g������ aŝ���J3���!�of��\�_�r�&�� �D}$���ߓ��������z�$��v��k����K�M����T�F��-I�D�-�5ۚ����b��TC�#����'��v�妱��!��0:�b�ؒ��H�t=�uRd����ݩ���V��T.*�@Я���Jg/f�i�Wa�]BN�8T-|Q=Kw����*���~�[�`�ڥK�c��dt�o"���h(�FG��p���uuc�O��;��3}t�z�=<��~�;�p�'y��v��l+a5��������=����_N�v�Us�䘸ǈ��5�/�Ol�f�{���$�ytEV8��>.�i]Ψp|��0Ͳ��{$��8Ԏ���/�ʋ�~X+�J����T6����C�B"�u˥N �A�~���c'OF�oZ֯�|��;�y���ލ[P�����@�
	˥�P��T��o���j�J��;x�2���ߥSj�fw���v�564� ��=2�����D8mP��ӌ�#'�r��}����� ��t�Y�*���[�(�1=�u?��������/�GC��Y�(۞s�8+C����3�
4�Xr�������\r�b�f@�����3@.#�IS����qD�$w�|N;_@��.e����J�1�`��3��{����(|����L���N���e�h!U�˸$�A/���= K��}�]��{���r��Z/n9A�x8��k^��ƈI������a�@(Ye��N��J��Z��:'B�k��3ko	����@�N�׹3X2�`��Yl��7XI�`� � HA�7�8�u�_\�-����2͵-�:�
m��8��q��u��D:�T�Gt-FcFO�����gOgJH+�wZ��J\m��}�2�O�	�T�+���d��fn)ik�p5G\�ZY�}����UP�J�3��) oXn(�^����z7"�b�&�� �>`G��+ȇ�j��32��N��2S���ʘU�Gx���qU��`���Z5R|���,���j
��K:�Lݜ`�;ѐ�q���
��;8��jrq�����|x��������g�9�}᜼7n1	�[%HR�F����R���24i�вV��5d{�&��/�u���*9c� �s��k+�4l{��&�IC�0��O���x6 J胖kx���ٽ���|�T�E�G�b2x���^^W
�P	i�6�ҝ3��:uE�A
��YzVܐ������f��Qb7���m�����,��MD�C��$�T�q�ð"������%=,�>Ѯx���"��%�q��s��:[�>�1ˠ9J B��d���ᕴ�5�rk�LĘr�+���~`�|�x�%�X�?%�b��T��,=��?��[���s r�����:�`w��k�'~r �9��3~@�"��W�LC:�_؟��L��9뢍�;h3��̨��������k�c��a�T"���-!{9��&�F���P�,EO�r�ap?	��)3� !�<�;�j<������]��� ��I���H��h�N�;�����#�5_LM_�2o7VW�-H[tm�\���9�r������slں2��q�������pm�_�4;���ɴ���S%�E�
��M���	2��JЯA p���ɾ�v�z�R��xԡ��[��i�m/y#VX�h�E͉�����ěo�(�/��'O���"V�'�;z��h��0��|��Q�� ��~i(в��03���m�}�J�y������#�CB����W
�r���.�}r� B�	O���NY�W�jY�k�
 ��oag��z�dJ�)�y�nW�Oo\1�Q��qL�3}P1�I6�T�d�/	�%�x����ay���{N#�1+�v��e��ţz�B���U�o#@�j�<�����2t[h��&|*y,�n��]����W��o�&����;=�(��Sm�	/�!rK�5S����?I<�?ν���=�#k����@�gcr;��׬~o��z%#z�J��8u��$����ć	��`�P�P"���BZ�ݜ̣dq z�^��R=<J%&�����D��$���/k�6��1�Ts�w�t���&c|�e�8�E�W��=��O�!.�s%��|#��w��ּtM�}��:��︥,L��~q%����#�̹�M}jN*�"]2Pw'�|7��o/���H?��\��L�z4t�U"T�'�O,N��yom��k�����Z�=��G��|�o�Փ�6<�7�]̈/q�4��j�<^��2��	�f\�i��<��P�F]�~�ŭ�H��φ�����	]�Nr�ۆ�}ZȽ���\�͛����7{~!��gǟ0z��j��4"l���h�8�5({]�����nm��(x��a���v�a�����J/�.+� �y�����i���l�ir�e���[TJwR�c�m\5���F��a���xd7��jO� 5�o�(�%�qs�2�1u�c�FI�j6��NU����_-/q�s=�CO�C^4�D�5K��L�+�����m7"E�/ʽ�XK������Kэs���ݝkX\��%�&f;�X�;�}���:UFI�І�7�;T"%�R�����D��L���&�m���*�2<����j79c)���Dk-�3��S��$JQ�T��|gِ?-����{׺��#�1Ƙ}�`'fv���%&���cl�	�*1 ��,���:f�Kjh�x�՗d���2e�amh(�2�`8��vo(ĵ
�����ν�F���M���R���tX�F���뒯��g�R�r_�~�^�&�gX+p�G�}^�g$�Z,Gt�{�rt0Ө�!��gm�il\��&��c�$A���Rmt#CT��3b���q�1/�<pAmE��P�yT��~Y{v_��V��qV���l��nn�(�b ɱ�⠊�.m:S�,����46�M�(�z�M�1l�=��[�@���0c]U��u,�������[�����P~`�����,�%�33>�!�?�*�,���&���b�!��p`T-��>js'��c6�8@�n�m)M���6��A�fH��R̼N{dO��Y˃�A�G�s6Qy{ bH:6hg���Q5U1f<�E@�����u�R���]��)�k����t_("gt���վ��o˜Rn]Od">$�/^Ҫ.��z7j��T���qO�'���BƛplD� he��t7�2<�؂���ȴƝ��,ҍ��Da:���
օ{-���R������Ϩ�<�V�.��*:b�U��.v�=_D������k�w���Ӽ���}��� ��s]p�O=!qT��iX���;�ۼ��σ� �� W��wR���3��\���&;�e,f�~����c� 2�R��Ϸ�v�d�n:�����fr��Y6��^�� W0�Oyf�:L�8FxQQjy>��l%
~uggr�ym6��aEKs���B�"S��VT��:H���KF�%6D7.�@`0�0�TS��%Y��<�8d7 �-_-�n'6'`.r9��`�	�(Q����Lқ@$-ڸ��"1���{s���X~nH�!�^�kv]���^k%9���5�b�30���}Y�,��ś1�:;���'4��t���+��s�n���ϏЭ�Y�&����q�2_z^����zىn��S\���BLڟ����G�i#K���@�a���%�/2T�d�������-:���ܰZ����T�\"'Vø   �  R  �  �  O*  �5  ?A  �L  X  zc  �n  �y  ��  ̊  D�  ̜  �  Z�  ��  ��  ;�  ��  ,�  ��  g�  ��   �  f�  ��  ��  (�  j 	 � 2 � "' d. �5 �= E L FR �X pZ  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�xR�)�S�y���u䐷Y�m��ìS�4C�I
Nԕ�d��Ų��G ܜ{����p�qb쐪a��1r�a���ēc}��[�.��m1����cC
QV\��"O\��G(=t�,ya���:�0e�' �p��Ü-�Q�� �t5��&!D�<�F�8NԲ4�g�Q/.�|ZVK �v���R�P�V�Q3m�$����Se��ȓ*�.a)�%�54�����͌i?��S�? ��: &&<�tHp'�H�G���"OXui�JU5m���p�G_[�xHS"O�(p!�#Se��N���(0�"OP�HE쁨3�r�htn�@�>-sE"O�YP[�8c�i0OY_���)q"O�LRAH�%/$&�J��Lh�r]�"Ox��S���C�l�XD)PUݤI�"O֌��T��X��1�CC��0Q�"O�|����)	 ���@OH�-"��!"O��;V,�=g���JA�B�3����"Oh��3Y�,*�Qxc�-Z�t��"O4`� �3+��EA��}�I��"Ox0��V�f� �
��L�P���C"O�h2��Ӂn��<�#%	l��a�"O1Y�#�3��� D��|2�Ȑ�O��=E�$�(�̥����%VHjD� �y�-.Zxђ�A����7��ItX�8s��A�1�"��7��r�A<D�ܩ7*��!�y� �|�Xh
.&D�D�Z�D0F�VH��`�8D�X��i�"~�䠅l\,@�
(��`6D����k)Tp"`��h܋^�@m�Te5D�����rVd	�bM*b�1�s9D��hSB�x9��c��?3��`3֊8D�	Wo1Y�L����G2 ��D� 5D��2Q�1Q�#��'kVq Ã1D��Q6�^��p2dD�#1c�1D���� A�ds�k�$5� �!�<��2����-$q��Kc�X:�Re�ȓ%y�|�t��:x� �;tP`�ȓ~���ƨͳ>�p��K.IXZ��'�ў"|�A�&�<��3\BBש�D�<��'W-�*��5Nۨ%�J�q`����=i1�� q�jT	����
�t�1�B|�<�&H�1Z��`#'L�
6X�jG�@�<q���X{�pW�H!%�>q���~�<)���kv]�Tg  ,���-J|�<�7�ׅsPXӷ`��H ���an�<a�͉�%��0s�Dv�$��%�L�<�ኍ��rU�-��pu���d�{�<�֥͹�
�G��.�j��f�Jw�<Q�-�#h-������E�$���Oh�<90�Q,9�(���# �ZL@��Y�<��MV�0�\�8�HԪ��u��T�<�4ܱoF�cR�Ӳ����G�E�<aCP'o`�ĩ�-�����n�%�y"EJ%㰱HB����LU�ͬ�yb+��"�e�r@H����"�GU�y��l�"����	�`�#���yB���H�+�fN�M�$xbV��yR-P7D+�l寅�bh.ABG�	�y"b^7!3�����#�tP�a'�(�yO�)��Lc��)o�(pqρ��y���.�`qD� %�m@a����y"b[�7"���k�4D�e������y��Hb"Vɑ�c[,3�>(#�(	��y��ki𚂤#f��6���yb��<��9u�^pp�� &�X��y��Z�F�p�I� �f����.�yb+ܥ%.�<�W�MY���
5A��y%Ϟ#y0��Y�KT@��"=�yR!�,M��a��4�	�B�y���M�\0 ��h�����&
�y��ˇh�@��HW�_�"�s���y
� ��giѩU/̼��/Qf���"O���2o�&K��9C���Ĺs"O*��熗.T�Qk6��*��!"0"O�AP��L�:������`�z�K�"O&9�UH�,$��kCK�s�`��'���'���'m��'�b�'��'������G����X��)2U�'���'�'��'��'�"�'���
T�B!٪a��F՝LS�ʅ�'ZB�'Rb�'O��'���'YB�'TXm ���/�b!`�ޯs�>8r�' r�'Z��'�R�'�r�'���'.2I�d.�9���Zt���O��E�V�'�"�',��'���'��'���'�l,�C�#PL��_%~�
��'���'�"�'���'r�'�b�'�x��%��K�TP����&��=k��'}B�'��'���'���'�2�'s��ʦgҹy&�q��M-�H<j@�'e��'�R�'��'0��'�R�'b��7M�pXf��ԣ]�{���.�?���?���?ͧ�?q���?����?�#��d�]�3�G���P�db���?����?A���?����?1���?����?�q�Z����c�C8�9C]��?Y���?���?���?!��?i���?)tI�"�U;���ju|i
�$�?y��?y��?���?���?Y��?	@�\���;Ge�g6$sS�(�?9��?����?���?��87���'R���3�r�RtÓ�LcJ����
ʓ�?!)O1��I��M�ČFm���K0M�;>r�%	&4���'�6�6�i>�	ß����&�$i����;b�d�៼��� �(	oZI~26�\���E�)�2�H����<%���0�aL:D�1O��D�<a���P�qO晀��f���ʔ��/0�j�o�o1�b���g��yHZ�`���e�+C��-[�j/F���'�D�>�|�'�!�MÜ'	���WkK�e�rPb���i�9��'��G�$���i>!��1T$Fd��%9���2�Dſ'y��	vyb�|��qӎ(j��Y�Y d��[n���CB��j��D��O����O��IG}B�(Kf  �t���}g^h�����d�O�H�1�B�vO1��L��vOj�� =I���K��W�0�ߕb�ʓ���O?�I��b�[Ƥ�;��E@b"O	��扲�M���t~�GfӖ�擴n$� $.MxΥ��%��J+��ݟ��	��@�,^���'��ɒ�?�� ��	V�&8��	��k�"��ъ�A�'��i>����@�I柘��%)ݴ�p�I�s�����D"����'TV7�C�&�ʓ�?��4�� \��Uj�0_���I�	ؒ4����FC~�*'�b>�#�Y�e���!7�=��a���rtd}9h�̟��Q��B�GVֺ[V�x��<IF�oc�Y��^1�e�ǟ�?����?���?ͧ���ӦQ��O�d9T�]�x>�#!*I8y�l2�֟l��4��'�2�v��tӺ�DJ�H2����
�&z���D�e����d}�p�ɘs��DHr�_�9�dp�[w2R�O����q�˶[^�X ��/ ��sօ�h�	ß|���\����4�J��L�'��2B��_a8��=�?i��?IԲi$�q��P�t�ݴ���䔻%��;q�� Nہ6�r]�Нx�'��O8(���iQ��n(�y��T"f,چ��X���&�ܓ���`�Ry�O��'Y��+LQ� ����,��:w
�*b�"�'��%�M۠�[&�?9���?1-�*!�@�!np���a��B�s񚟌b�O����O&�O�SI�jŁ�9{l,i�"L�>6i�ĩV��,\oچ��4�����'J�'i�5�a���>]�e�<�u��'1��'k2���ON�	��M���j�,aa��"�x���Z��.Ox�nZi����	͟D���R�^�Z�(dO&���VI䟸��>54l�[~Zw�Z� #ԟL˓-X4$�6`؊W7��j��^���̓���O����O<�$�O�d�|Jt��t���􈓠&�:S�\��G��s���'&����'�.6=�Ypf�S�'�8B�	C#3���)��O��d�c�)�ӍQ�]oZ�<ْ��<Y�n}�A	�!'�(�R���<�խݷ�N�d�����4�.���b$*iJ$�%�`i�@�ɵ��$�O����O��t֛���O���'��NϚ1�f��i�:D�-�f"�l��Oz!�'���'��'�f2�\tx�8$��|v�a��O8��sȖB݀ؓ��7�)��?����OHI��Oʯ@[X��ň�>T�(����O���O>��O.�}�F3��r
�_>N�Hӡ���	�7�vZ�m��'t6�,�i��0���cw � t�n�hw�t�`��̟�I;x��	lp~Zw�n�x�O��!2&�gв����x�8Ђ�A�O�	Zy��' ��' ���yG��&~��i�u��:$�P�p��=x�剭�M���?����?iL~���� xh��]��)[�Je�xaC�Y�l��ҟ�N<�|�%"�E5n�i�,��4�PI1C�A�`~��U�Z~R� �&����5��'�剪U�q��]��=s�J+����I��	�(�i>��'�D7M�o�R��-P��*���}�� �aV;O�8�����?a�Z����ğP��4}��`
�AL6��ez����k6\J�	�/�Mk�O�ur���j������ �)�)�.���ʶW/w@,�=O����O&�D�O����O��?�jB-P*JDy�"?����B%���ԟ��4fn`�x-O�AmZ_�	&b4H3D�Tb���ٴ��7�hJ<���?ͧs���[ش���PP�3�\5<�P�t��(�\� ���?�C)5���<�'�?I��?�U�I�|)
��˥���wmԷ�?�������%�ת ���Ɵ�OE`�
3 M�e�t�	񪕳=`���O���'nb7�D̟�%��|�@J#$I���� �BJ�~t��
�&51�!_���4�� 0��y%0�O��+R�QX0�'�)J��#D�O�d�O��d�O1���$��6�kP,uc�n���
�던��Y�FU� 8޴��'���]���ז
�%���C(d@ͩq�х�z�$}�Ph( k�B��fP��a�����.O����lL�Yȝ��m^�7.Lx��?O���?����?����?Q����	D:2Ց�Oڦ=�r���ⅶq�"�nZ�pb�Y�'&���$�'��7=�v�:'�W��������+D)ij�O~�:���\�- 6�v�ЫZVYRGj2�ـ��p���%B� �0�'��'��I埌�I8C���%��"j���@�/Ԃ%;��I�����ʟ��'��7�Me�\���O��D�SHq�!#X����Ǚ�eՌ�T��OunZ8�?�O<ɕ&���4f%Jw^0y �w~2L
J�\d��O,��d�B Ig�� 4gŇmB�h֮�%B�'k�'�r���P�"/
�<2�|I�.!*zB��R(���8�ٴ;�R���?y�i��O�n�2s4P Zi��G��p�)�hZ�A�����McE��M�O���i̦�bG��*����e
�#���@�b�OK.�O���?���?��?1�6h�9�LU)fIz3��Ć/�D*O�l��#C4p�IП��	q��П8�����o�B��R=+�b��3c\%��d�O�6-\�)��� ����S��x	B� @�@"C5���Q�љ8a�ɁD�jPIS�'~'�X�'N�
�R�7NHs�`NBȼ0��'v��'7r���U��ٴK]�)�U���i�DJ�N�6`��%Ɉ_|��@�F�V�$�Sy��'}��v�4Ƃ�	T�J�LV�c�ia�KP:�7(?!�Œ/GŊ��#���������B��B�Q�����u�(�	�D��֟l��͟$�Z��� c̨{�IE���,�T�F/�?9���?)��iL�R�Њ�4��&�� �\r,��T&O���06M	�ē\��6�x���Z6-6?yrJ").F1Hu��/I5䘚����d�4�"�O���L>1*O��O���Ojt�g�Q-)-�0�4�'*,V̺��Of�D�<��ivNd��'e��'!��������;IG�(I0��#E(�:���낄�MK!�xʟ�����p��c���-VW�KE�^><k�aH���a��i>����'�t�'��H��K���!�c�qYD`�� G˟L�	ܟ��	ݟb>u�'J7����B@r� ש�h=q&.D�w#x�ۣ��<!a�i$�O~=�'��7�f]�x��	��ZBm�0e�����+�T���'f��𤆎�?)�6T��"c��1�ݰB��>����&ku�@�'���'��'
�'��ӾY��m�S����2�L�3�F)�ߴY�*d����?�����<q��yׂ���L�Bډ?�e�s�YB��'y�O1���S�Cl� �	�d���D
�w�$�Yp�@PJ���8h��'�$�0�����'>\�{�擑��Y�g
17��Ñ�'LB�'^"Q����4>�.��*O*��� x7�そ4^X �&�C�[,���O����OH$&�cǎ_(Jɤ�@�K�=��1%*?ɁB��+����a�Q�' ���D�?� M^'$B��A#>�����؇�?����?)��?9��	�O$�b���x��0Z�!�_��4����O:o1�6T��ޟ$�ݴ���y.�,.����r�A��9�&i���y��'���'C�ՙd�iH�i�Q�f(Z�?����6��t��>�~�s&I*U�'��	՟��	��Iҟt��%/^ƕ�Ed؍^`�ă	9���'�6��7&���O��&���O0p!���j���P�NƶV��EjDcPU}��'�"�|��$�Նc�)��)�l�LX��Q$UDvL�+�#��ɂG�TU�A�'��x&�@�'��\*�Y�jf�(ib읐LMF�R�'c��'�b����W���43��@��bd�ػ��<i`�2�"^$b��A1��"s�V�ě^}b�'��w.y�u�Y�o~Fċ�/�M:�����#A.��<O��D�6(B*X��O6�I�?y�]'�H�@-�&B
��B�VI�^�����I⟌�I�D�	E�'@�F���5� ��,�"��"��?��C�������T�'�x6m0��'�h�c�M�>Z��6��
`x&�4�۴*a��i�$��4��D�'�n�U��@�$=���9���'�W�?QTn;���<���?Q��?�$F�<*�qa/��AKY�WK���ٟ0�'��7m���O^���|��΄</����؅ ݾ�J� �X~���>Iװi��6-�K�)����7@�ŀ3�F!£�_�.yK6`��tV����- ���`q�|�I��Y!���#@;|�}P�F�=*���'r�'@���R��2�41h4��.U�;��;Dd�g0�m��
��?��M�F�dQy�i������++T��v��G�ysf�m�d�n�8<��mm�f~�=+@����}�� ��w��$q��9���U ���9O�ʓ�?i��?q���?���I[�p3"L�Յ�8�`=q��8Z��EoZ�tи��Iퟨ��w�s��S����d;-�&� �*T�&UhV�Q�m@���wӾ$�b>YZথ�kQ���,�� ������%��ϓ.˶x����O�]�I>�(O��O !(S�	�,X`��bZh�bd�O����O����<Ѳ�i�d���\�����?�pd���]�z��%Q������?�'Q��ڴL��d!�Q^H�a���R�9�H[��Ix��]���>Pc>���'
P��	�W_N5��f��tcJ�ⵌ7P�4��I���	�h�	^�Oa"E�4����Gk̕���C�_�^�b�hh�ᏺ<I6�i��O�nh���'��t�m)#��=^(�D�񦅘ݴAZ�v$E���֛� ��C�z���-խ~�Xi'cO�W;���m�?7�<�&�����4�'`��'�"�'�ҽ�"�b}�"�E�~>LU0�]���41b�����?	�����<��.$=���![�n�+0lF�<��Iߟ��I���|b���GƑ�w�~8�&���3���&\;l������V~�oͮv�B��-��'��ɚ9�:u���H��0,��Fe�4���韔�Iӟ��i>u�'|�6-�{���d��S�
���QAb�ሕB}��Bݦ�?a�W����ɟ�	�G~���D3g�C�$;g�\+�$����'��$��CQ*L~��;/f�	���ӽ+8�J6H�� I͓�?Q���?���?Q����Oq9YR�QT/٠@�B�`թ �'�2�'I`7�J���Oh5nZQ�/x�Vp#�(ڽAB
Hc'(M�F؊O<�ײi�67=����֫t�"�^�歐vȅ�
�	��8���M0�J��>g��O���|Z��?)����Py��6�2əFaԕ6=&�:��?�*O��m�9=1� ��֟`��[�4"��'i�G],2�h3�Ţ����x}2�'��d0�?U׮����ɺG�O,��áʥq����V�{~Ҕ�����Ο�IÒ|��A$%�\�u͜%:@
I:A@�y"�'���'����U�� ڴg2Y�@R�%FTsEƱ2/ݕ�?��k�V��X}2�'B20��Ѻ1�y�,�#.S�#$�'��f������]�1�
����$̕	Tpڷ��g�JA
4�Cj�ĥ<!��?����?)���?�(� ��C�,�@BUi �B�%Ҧ�CW�EZy��'��O��q��N�
���7�фw�Mk��ѐ3c���l�H$�b>�s�F����͓bap�Q�JV,�@��B�9l����$���+�O@��L>�*O ��O4�1@,�]U�u��+x�*.�O����Ob�d�<)s�i�>A�W�'��'�&�� �B��\�
�%ۤ�u����a}�b�.��	v�-h��ͩs�D�}v���A�o��=�Z�@7k�<,���O~
+�O�̹�j�̸��L>l���W�UC�����?y��?���h��NB�E���B�=il�Y#�Do�>�D�̦����M�����'�M[J>��SdG��1�qo�I��`�'���<A��?��H�p�4����`3k����ArLJ�)p���A�Oƪ�Q�Jü�����O��$�Oh���OR�$��k��u�J�2ZV-�������ʓ2���,��,R�'�b��t�']�P��EMB6V ѣOÚtj6�Rf��>���?��x��D�ҹ
�� �ŪW����'g��"F�P)���b��C�U�O˓p� ���H�8d�Z$�X.0�dYK��?i���?)��|�-O$ymZ�d֮��I�&d�6a��I醍���5ڤ�I4�M��d�>��?	ƴi���k�nU�+)���D�/�N���`��6���;��h��$����j�3���'Z�D�aj>G��k1:O����O\��O ��<�|�`�(^T"p��# �*]*��:�?���?ѣ�im�q[�O��a��O��WL��_�Ձҥ�{\5y�k^@�Iɟ8�i>Y����%�'� �*ֆ��;�(�R�IP4[#�8�f*izlU�I,E��'y�i>��Iӟ���*MR�LXs��=�f���#��Jp=�	��'��6m�>~���O��d�|R�ƝJLl�Th2��f�~~B��>���?�L>�O7<UХ	�X�hE�BBΒYCd��V��]9�D����6%l�i>�8b�'є�$�@K�WRhش.I4Y�8��b����	������b>9�'�7M��J�h�W"��*�ݒ��ݫ1l<;�$�<��i��O���'��o�T9�un�"��9�򡔺h;��'xrI0C�iF�i�Q�5/T�?�rU����⎟[�PY#A$�dm^a:�#f���'�2�'b�'�b�'��S�aTʀ�T��$�.��q���㦡z���ӟ��	���'?�����M�;���I�h�k��ж
�
+�M`���?�N>�|�r���M;�'�z-E�ٮd�Tј��^�YĴ�+�'���K&�̟�՘|_�0�	���Ka "%�zHf�_�H4Y�P����8��៼��Py��`Ӯ���o�O��D�O�YY@'��&���M �f����>�	���$�Of� �D�Bz|�A��U ��� ��O���#�@����Ƞ#<�H'?����'6�l�	,4�<�0�	9�  ��A� ����	͟��	ğ��	j�O�b.�7F������G�T<�!�$\���gӨ���O ��Φ��?ͻ]�씊Ū޴3�`�ɋ )��Γh��v �O47�ό1��7-6?���� ,����Oi�? �h"%��3X����f�da3&�D�<����?���?����?��-K�*�p�0gI�T�T���L"������0�nԟ���ן�'?���n
��{�nCpC��F��9����Oj�oZ��?QI<�|r�"!5��Q���_5���[fb�&1���Rp����$��4�� ��w@�O���Z&�ȳDt90SA�J��4����O��O����O��<	B�i��eq%�'����%n�:�@��H/�ਚ�'r�7�#�I���D�O��I��m�sA�h8��KN�Vfb�FQ��V����57����'������,X��(	$gĜ�@ެY�D�O`��O����O��d1�S i�؀h�˩m�Tpq$[�}j(��ɟ��I	�MK�E�|"�0�F�|bh��� A!Th(�ؼ��
|��O��$n�����s�i,�	�q�jt�ǍD �I1��ê 4�#r
[~�rN�F��Ey��'��'bjҙ*����Ó�`}�OǾS���'��	0�M[�j ��?���?�/��<�'[tt�P U?R�Z�I����,O���y�B�%��'t�:@	�3bA�ͫ���<7��[G�b���;$�y~�O�\����s��'�x�0s!�'P���/Ef�:(*�'	��'�����O��>�M�BAX�IxLL�uo��(K���-D.L1���?A��i"�Of��'h� ��\�)���J�@G�ы�%�:S�2�|ӮD�4md�J�� �RAE���O$�HvlC�P�T-���V�L��T��'��	������ �I�0�It��MD�U�ڰ�.����!�oۗz����͐v��Iҟ<'?5�ɷ�M�;�֤1Č�Be��
$@ȔQ �����?9L>�|z��G�M�'�$�%�6?�l���M�K����'@� �s�V������|B^���I���K�Y��@r fO�i���oI���	�(��Wyb��Јs�ǩ<�!,�)Rl�y��A4,�1��8��O�>)��?QL>q��Y�PD�j᠐�8��Ё��E~���7�`i�c͕�F�O�du�	�ڢ|��Ա�
 �h8)s��j���'�B�'���� ����y���1<� 9Kd���l!�4ce�".O&�o�W�Ӽ�jH8>:��0��$I�|1�-��<��i8�6-Ҧ��+O��E�'B�<�"��?1)�E��h���'e:�+�`�.Z�'a�i>��	��$��˟��IE�H�g`ȕ]�
Y���%3k���'f�7m�:u�&˓�?�J~���4�xǣ��a6�ljTʊ�2�bU�7[���ٴV�r�x��$,�Ku��U��5&8��B��5���{�aS��� V֔�#�'*L'���'����� ?�4<@���3���P�'*r�'�����DS� �ܴ=y����g�B8{�C�m��Y������a��1����N}��}Ӣ��I��k'�./� c5h �`R�3��J.t�Eo�X~��H�+����S�;��O�g$�X����5���Q��y�4��y��'���'���'����Vz�b�����0V�,i�ŧZ�k�d��OX�����eaVI�my�cy�N�OB�����!D0�<�vm$gc>	# $�x�ɒ�M�5��2����M�OF�K�^�<�
!�ĬrW�\x +��}9��p��ؒO�˓�?I���?!��Jr��L)K
��#�W�o���ȶK�O��ģ<���i~�1��'b�'��S�A�ְ#祐�i�����K�|������MK'�'剧�)ӭƠd�E'O2j�"P�
�a�6ݪa�ځ9SRq�d��<�'m��ē	��#�0̀���2 �Dm�0�؂)'�����?����?�S�'������z���+5�\(���j�[G�ơ����ҟ��޴��'k�듃?�&���r,�8i���G�4�?1��+���Aڴ����(8�M�?Ֆ'@��i#�Uẽ[�F\Zh��'��	�,��ܟ�������IZ��N��Q` m ab��� �d�N��6�@�5!D�d�O���=�	�O�ilz�=��E�N(� �^�C�������IB�)��5,2Po��<YbK��DB s���G��i����<�A�	0"�	I�IPyR�'r��=\�@d�$�������'t��'��I��M�G�C��?���?�0�?�tej�KLn���ň��'Ar��?i������ijuO	�O�@�� �{��'�$�����Wi�v�-�I�~B�'�X�Jg��P<�`C� ^}�\���'`�'��'��>��I|���k�2�p@KG��r�I�I��M�p�\�?��a�6�4��i�
�hnūcR=�e��>O �n�=�?��4]�
l�ش��$=�i����n�`#�di�h��(�-'}T��?�D�<����?���?����?�v`K�4�25�p��6�y�cѳ����Ʀa:Q��ʟ�	ٟp$?�	� �^��b���l�q�_�R<A�Op�d�OƒO1���dG;6V� lJ���(�K����3#�<���/
=>�������ߋ9�
�ET'7��L����u�����O,���O�4�J˓/��ãM��"��zԚCT���i�T�8�yҀf�p�X�Or���OJ�o$��+ �N�o]3��8/m� ��b�ᦅ�'���C���?��}���%I��𩙀��y�ea.�͓�?����?1���?	����On�a׏2��k`%D76>�HڢQ���	��MS���|���T��v�|2��}�*�X�&'������"COx|oz����Xdc�,� �2�� �m�S)B�v�N8�6������&�?9��-���<y��?y���?�7��`5���T���>I6��A�P��?����$Ʀ��gD�wyb�'3�S!	Dp�p#�S�P"���y�L�`�ɖ�M+6�'���)1p����D��v�17a�-h&ӆțE��`K!�<�'h �d���)ؖ�q�� � EVf�>k��mq���?����?��S�'��d妽q"�I>/�4CףÐK��AP��f���	�L��4��'H.�)͛Flɥr��h�@��]f�a��*�"����m�@s'Hb�R�^nx���$�0/O�+`�_�G���z�0"�a 3O�˓�?���?��?����I�3X�(��6{�V�`�o���	n�9��ٗ'"�	���ݠ5�,g�T�Aʲ �$�Ɉjb�R۴U⛖L0��Iau��ڴ�yr�;D�@�5T+�N��Vč��y]�D���,kD�'��i>%�	'_Z����/�m�<踃-޿}���������	ɟD�'�>6�8jN�D�O~���x��[�)@�3��w-L3G:�裪O*�$�O��'���s�Γy��e�$ŔD���P�'?�6�B�>��k`AYJ̧5����X
�?Q��$�a
sgL�:���	M�?����?����?!��	�O�(��i�6<�z�3Ć'�^�� �O"YnZ�o�ڜ�'φ6M2�iީ��	^�3(襻c�*�a!��|�t�IҟЩ�4uJ&=��4���N�|���i�'K��q� �	f�ص����X��k>���<ͧ�?����?9���?y����F@q�W�U�ɱ�)�����m�AhN��|�I���'?u��-lZ�<�%�&k���3�
N�s���.O���`���$���,�c�P�
� !�4FOH⮠�S��o��� ��PAC�J%�RT`��Ty"lJ&`�~A#$ڪ~�F%q����r�'��'s�O��I��MU���?Y��U��`��
�2(|"��c\��?�$�iR�O
,�'���'�6-D�J�(+'D�gRM���� H������o���.���E���>���
�N�Qj��K��x�i]+���	��H�	���	ܟ`�	[�'�)�+,;�`AqӸI$�(O������J$�`>�����M�H>��Aͬ`�m1��	'<��kr�I����?i��|����M��O��,V�:A �V*(=�nN6~��;Et$���'��'���'Q0<²n˦q���c�L^�dӀ��'��Z��cܴ,��e9.O���|ʢ��)�^�C6oDZ͒ �<����DԦ�X������|���6���yf 	�M!l#W��(@�
8�h
J�t��5����?��?�q�<��L_�U�����4(Ĳd�]�l���Ov���O���I�<1$�iq��D�$5�@㖑L2P�D�&@ ��'�|7#�4�p��'!bIZ�?6����H�Q`y���m�R�'�	 �i��i�A	S��o*-O*q1�͠9��D���[�wl�t�;O���?���?	��?�����	�R���s��=�>���B)5Ǣmm�k��1�I�l��x�s�0b����!�ֈr����0�`�za�E��id�O�OS�����iq�$5-�LѢ�V�֩�Ui<� �D}��\�l�OB��|��E��1#�Nؽ�yk&+E��n���?I���?�(OJ�nZ�3��e�	ƟD�ɃE��l�� N!hB% 3��$�?��V���	؟($��Q�'@�/�b`!�Şp<�#b�)?�BHS�x�D�͖��'Q�����?�`-.bY�Б/���D�)����?���?y���?��	�O2|�QF��DHq+DP�<
���O�l��uEl��'�,6- �i���)O)GB�Q��24��lf��	͟�(�4\�Hh1ڴ���D7�P�'HyD4IG���8q��e.a`1��g$��<ͧ�?q���?���?	�j�8xL��k����dy������ЦmP�����I���&?�߶���HҦFx�e�ˁ#�$��O����O
�O1�������oT����H��m�c��z� �G�<��i�`a"��������d�$_zL���Ȗm��[@���r�T�$�O��d�O��4���U���g�2Og���J������(2���aX�G���q�d㟐2�O����O��d�{%��ZW��d���p�Q1Sv�xa{�"�FŸL�����xK~��R�T���+�Z ��(T3����?���?���?����Oa�H�v@&Ҡa�͆J4�|Q�'��'�B6V�x"�ʓ$Y���|rĞ�ek�=Q@	"������E�';���
�z������e��#���'

8�r�D�7��1X�k��Xy2�|�[��	ğ����pAs"�=S|����1hc�,C�̄ޟ�	Sy��h�J���O��$�O�˧`h���X.f���F쐱J�zu�'����?	���S�4�;v���HP�$��Ы���Ѣ�F�:V]�RU��|�ҡG�I}���ao����T��Ĕ� ���I�d�	ş@�)�Ny��vӠU��l�!}y��h�'\(F��b%h��ʓA��V��g}�rӜYy��]�u�6�rAH·޸Z���՟�mڣ|!��oZA~�M4}~��S�'�I�:�,<��/`R,K �2P�ry2�'�b�'�r�'�^>�;q��
�B$zW�.PA�q�����M�(��?����?�O~ΓoǛ�w3$�H�gP�.�ؑ�F(A�jZ�\7�':R�|��T�3iߛF?O� ��� #�$�5�˙,�|0jd=O
0B�� �~r�|"P���	���HP�R�����_��P�cş@��埀�IOy*}�F\�F��O|���O��$J�X� Aj%�/$Y�h�R�>�����$�O��d ��^�{�0 :w� <������E�Ri�	R]�R�V���M~�娟��	�Z��qZ�iU�b���2��������ퟘ���<��T�Or�A�G�����ƒ�c����5^�t�0���O��Y����?ͻ_�Diī�W�����m�D��?���?!ł@�Ms�O�N�j��S�q�,�A�� �����A�5�*q$��'��'&B�'#2�'���rI��za�g��d�(d1�R�8��4sp>$���?����䧕?iT��44�]��l�7�Ȁ�t�������X�Id�)�+gӞ���lUco���4GD�Y/
���hӺ��'!*t{�@o?QM>Q(O����n
��b��Ї�=~.��t��O����OB�d�O�<�0�i�谳��'���:��ԨY8 XpS��>/*�I��'(X7M'�ɬ����O��D�O�4!�k�u�̱:s֕�TP��F��4��S5w��01�O��O|W+D�t���[���8L�<��w��y2�'��'���'�2��"vL~�)6b�Q|Tizg��:}���?�d�iPC�O4r�d�6�O��Q�֦Wo""zJ� /�b��O��$�O�i5,v6�-?�;HP�d9פ�騰�!�W9<�6@{&���?���#�ĩ<����?����?��(Hj��@q���v�5[Ce��?9���DƦi�'៘�Iϟ��O�$�+`�R*~Й�񢔚X��(�Oʅ�'J2�iN,�O��-C��
���$\$��&2 ��2k��+��mK@'?ͧ#U$�ā��1�$� "ھR���XS��"}�������?���?��S�'���Gߦ��5iV�m<����Ņ�uJ���H��d����4��'��듐?iũ��C���pL�M��Z����?!�1�(,�ش������?�'ͦ�GW#)Dĩ�F�[<Z�y"W����ߟd�I̟`��˟��O�����N�!�l3�T<>�{
r�<3��O���O6������]#Ev�U���$)�SL�Rе�	��p�I<�|�b���M�'I�X��*Gh���S# �zY�'�r��j�� �0�|�Z��ß�"��J
<�J����I�I
JG��ퟰ��ޟ`�Igy҅f�����O6���O�lȱ�I�W�N�!�Ñ5Ub�1#/�������ON��1�D�)ea��S�`~&��P��"ro�I��� eL��J~j"���l�ɔ,��}��J��"r�d9�Ş��H��П�Iџ���S�OTj��f��IRm13DJ�q�B�-���h�
d u��O��d���5�?�;
���sHG�/��@PᇃD��d͓�?Y� ��/��&���P�A�lq���Ј
LȔ@͞'Q�$�t�]�5J��$�,���T�'���'�2�'��l����g��b)�j��#Z��H�4��P�/O��$#�	�O"�����b����-άn�c!OAk}��'�R8��)��
`z�4�ڲo�� tl ���ҡ��-F��	 rE}���'��Y'�t�'��x��ϵa@�H�k9@�FDr6�'X��'�����T��z�4&�={��Y(��SW��^���Ԩ�T��͓>,�V��\I}2�'H�+e�jD��A��f5�5,�@�����,4rV7m5?1�"�S��)>�S��!��g�MHY�!&L�	%t�`BEn���IşX�I۟|�Iܟ��%��6�zy�'J+{!�t�ԝ�?A���?ֶi=f��3[��۴��B6i��W�'72h��ខ��5*đx�c�V����	�P�{��CBi"��ņ��d���P�რ��E*L��M������O����O��d�(}
��0&�*���a�ˊ�FX����O�ʓ3j����>B��'WU>i
R+��v�x���	N�MzH���*?��S�p��4]@xʟ�Hk��D�:��7d;?��V�?�.A�A���we�<�'�~�����@��sG������q���!���?����?��S�'��$�U;�O�F�V�#�����Ek�D�2���'�6M;�I���l�I�w�� �}�'�0�P=�����tl�TZ�	n~R���8���t�� T�f�9�d �` 5�F'WP:�	Xy��'�r�',��'U�Z>	��@�p��#�K�w��Q"��,�MC�&X��?����?QL~���'K��w�K�3��`�'��|j�ڳD9�?1���Şrys�4�ybA�I�^�,��`�	#c���'K���@㟴0��|�P����ϟXC���?�j�8e�߂o6t08��S��l��ş���Jy�FfӼx�/�<���4��W�B�~)r���?p):�1�-����$�O>����;�t��4�!6b!�!�4YF��C���ŉ�!#����|Z�i�O��y��{���E��4���g�V62w�����?	���?a��h����I'�܅�d�BO����+���$[ۦm;�	џ��I5�M���w0�� �g�10�={Yy�BE@�s�h��4���Ox�LIڠ�t�(�~º�*`��T �p���f�Ӱ����U�,��H�H>�)O�	�O��D�O��$�O&4�SɌ-\Z��D	�|���Ƨ�<�мi����#�'4B�'+��y2O͘ $F��D�u��I@.�@h���?1�v����OY�4K� �P3/0S��@`���k���9 AS�2��I+R��s�'j�A&���'�vdbs�[!�b�J��L'o�V��'��'�����$R�lR�4'?����P j���?wVNl�6DI�Tj��x��OC�����R}R�'���'�j�j�U	L����͓hE�Q�W��*%�Ƙ����!���4�I��j �5�k��<��']�*�╫!<O,�D�O����O&��<�|�ge�8��%r�I�O
��A'S�?Y���?Ie�i���ØO)��s�\�O�y�N*yyxm{c(E�Z�v��@'�W�	���mz>�p�ɦI�'ڼ`j��ЅJ �"�/D�#�8���oF�3�
A��,b��'��i>��I���ɡ_�MP���\��Ċ�3��x�Iϟ��'��6M��T�r�$�Op���|B��1휜 V�L�V�@�9��Y~�>9��?)I>�O^�r�g۴w�l�A!k�1W�"��6U�����i<���|�bG���&���T�C��P�Г! +Ĝҕ�H�p����`���b>�'��7���x;0�5ɉ�fOjA	����	���O���D֦I�?�U�4��(v�T4�C�Y�TtD��B�{����ßd���ئ��u���Tv��<�T�.6x|�rD\�]�zX�G���<�*Ot���OX�D�O����O��'2ᮐH����!cL���I?e(ݨҺi�jM�v�'8r�'b��y�a��..�dJC͋�Go�5�Z�5r�D�O��O1��x�/i�B托)�b�p
�	�$�"f�9L�I��0�@��'h��&���'���'�6��$�\�l	�D0q �,B]� �'l"�'I2R�tQ�4[�~�h���?y��5:׉�vm���dPY�9�R	�>���?�L>��^=?�D��-Ӡka �B��n~"D۰A�&]�g��W�O�"A�	
WA�&ar,"G)X�c�`4�g"�?"��'���'j2�S۟@3�
X�vT�;pl�v�)#�D��$�42�҉����?Y�i��O�ڎ ߪx�O؜�>٨������OD���O� �umiӖ�Ӻ{�/N��Z�MJ��
x����"x���"#K6�O$���O��x0	 #E�����c���֒��!�4_��}����?i���O�L5[�cH-r���P�*��>���?�L>�|��ұa�4��@��7�u��dO�&6�	�B���S�����(�O����u��
C��+ҫĄҩ��	��M[���*�?9��
m���)�8���s�bP)�?a��id�O��'B��'&'�
(�)��D�'nVꭐ�c�s��Ͳ��i��	�-y̕�E�O��$?���4ڐ��
J~A~e�H�3,���O����EO��P!@S�[3u@�=�F��(�I���3ݴ/��l�O��6�?�ȧO��BI����N�	X��O�D�O�iő�7�;?��b�:���
E͔Q�
'{̸AKѼ�?�l0�$�<�r�ޕLgʠ��?���sJP��O 9oڭ1'0���؟`��h�d�H�`~*�nO�/���FV%����\}��'���|ʟ
����rMf��%g�`p���,~^�[�Bc�dؕ��4�^b?�I>a�'] x�b��ۡ��Ձ�� �?���?���?�|�*OzYn�	@Pةo�@����Z�ǮP��&�ܟ��I1�MCI>ͧ$�	���UoZ�OL�eۑ�
'3�l%Xs��֟��I0���l�h~Zw�5���O�l�'���@�a��4ʑk¨Wv��'�	�	��0�	ʟ��	T�$D�y�6���aV� ��� E�[-6�6��(w4ʓ�?�I~��$ԛ�w��d��+�;v]l��+ѕt�)d�'9�|����?��9O�A��*��}����cRrM�d��<OD���Y7GЭ�T�ɻ��í	2|�J%C0�ޝ@)���j��&�Fhj��Y�iwD���0u�T����
��ȱ1�1�0F�  R���5Q�/W<X���q�Sf?�FM�?,Y�� ��%�%ò'zy"N�i��0,J%��)Sƍ�BB�t8�I
mՊ��lD�$Q��@�o=u5�����V	-�l`�c�j�N��%²=^�EqY��@x��
�@KIjR��!ߚ� 7f�1�0�U("
IJ�i�K�,W�:��GL�A�:Q�%��P����6�]�E�,���;> ��KǨ_��M���?q���{1r� AGTZ��!��BC�f�'�'1�	���<�	��~{�#[
KH�)S����^6�O�$�<�qƃ�<�O"��O�~���P��Zaҵ� t 0�hS�.�D�<�Ix���IB3{ֲ�q�A
"ז�����yP�v_��T�+�M+U?��I�?�y�O��BJǚ'&��	%_�Ia�i�副�0#<�~:��S� ��-��?�� ��m)�% 4�M[��?i����0�x��'��XѓLW�cD�HXb<���:�~��}���)�'�?ѧM -jd�bđlH<A�&)�
U_���'S��'���Y!�+��Od�D��4r�nE�G4R�Cn�x!
�
��4�I3h:`b���I��d�ɺ�UQs�X�:<�x��T*6���4�?�� �'z�Ob��:������ �ށ�P�~/Yye^�����+���$�Iȟ��'dȒ��S�}�|U!��� -��Ӥ
��i�>OJ�D�O ��<!-ON��e�׺d��܋Ib֑kC(�,1O����O���<�)D�D�I�N�����T�6��&+��쟴����ly2`C����-;m�d�A��T��[-�82 ����|��ǟ��'
Ș�D#�IN[�? ����oǄf�d�Q���p/�6Cd�`��=�D�<�SHB�l'��  `Z� ࠃ!Ȉ#<���l����I\y�G r��������xR��^-��8c�
�"un�B��YJ�	Uy�$��O�S��ީZ6Dܡ�ND���Ԓ{6Z7��<�F
��"��&��~
��jT��`@Mȸ5<�-хC�8~��j�'tӢC�	;!:B�P�&Ϲ�X9P�'ց|47-��9�`�m����	Ɵd�����?�ʒ�5��Q��Ԡ$�<�T�m�a��'vl���� P��`�E�Уyk��C��n����O
�d�,Q�$��'������mby��iF����d'P{��ml�E_�'����͟��i�a�r�F9�Ж�]�=:������X���q^��q�O
˓�?�J>��F ���q��%B�)�cѰ�B}�'4z1���'��I֟(�����'����
CF ���f
<Vz��XW�;$f����O�O����O�!i�晌���F���.	����*S��ON�$�O����<�bFS�V����6�n4��d��RE2��`�M�*O���<���O��d[{� �E|��83�glb�A��O̮PV�T�'��'XBW��ch���	�O�8#��I��|�G� W)�0�h���Q�	Py��'�R�'�.Y�T>�@��H*%�M�@���H��T�b�oğ��IHy���[�"맒?Y����#��9��4K�a��~�D9��B9Ɖ'�b3O���R�$�?�s�H��:H�C�mSd s���<>^q�i_"�'��O���ˇ	�z��ySaiF5Uv��#��妅�	���;��I}���ON��d��p����������q���M+���?a���S���' e04�M���#MU�t�����oӦ�8���OH�O��?)���BS
X��D�$G�@�%W�/���:�4�?����?����3D��dyB�'D���=B~̙�b�<����`�ǵD6�O���Ӫ1��ON���O
�)�
%da܅��Oo�l(�ceΦQ���%в�O˓�?�L>��kl&Y��ᇶM��H�>o2x��'� ����|�'�2�'���YNM�bVH�
�.�nuB�����.�ē�?9�����O��Ӻ��	U+t�b@j�<�j��ϋ��	Gyr�'eB�'�I�X���
�O���Ƞ��c�\���O6.�n|Q�O����O��O���|��	ZiX�A�x�s�=J�m*F�xB�'��BH�\���'�����pdX�����"4[�l��0�	cy#;��AE4Y���X4)�4��ȟ�L���n����Fy���9"r����$��klFĈv�>�$\�qe��qq�'|�	����Iz�s��]>lV6@��˕�ְ��Ń nq�6�<��!A�s��E�~���z����@1���q^��w�.K���s�'k���?���(Y�O���Mk��'1&Ѱ'�����S�[ئ}�!럔�	ޟ,���?����ɐ'
I(b��D6S������h�oژ,��e3�E.�)�'%�@Pr���8*S�%q�'"�d����i<��'5�E�2ss�)�H�,3���8�x�'!�)�H��s����'n�+�n9�i�Ol���O0���I4XaĽr�B�U�P�&FT��9���mX��K<�'�?	I>��-V����Xd.HY&�SL\8�'@@p�'H��ݟ$�	��$�'��q{uAܚ�B=���s��X�Q%E.W��Ot���O��Ov����5*�:k�`	��_$bҡkb����?�/Od���O����<Ag�Q�R�	���$j�-�5i^B�`���,��۟H��[�[y�
c������ЁWb��(dMs���V_���	�����wyrǂ�m��8ā5I����@�	A`���2�Z����	�D�'���'�n�[��'R�v/"M@%�:杀cׄ1���o�����|y�K"y �t���klS:kNL��Q":lu1W擽	Ӊ'u�əy����	F�D
fˉ�;�uв�|�P|�P��J}��'�����'�B�'�b�O�i��J�l��7 ��x�,6vm��(#�fӐ�$�O�U sLүk�1O�� x�ΗE�􀀷- �B1�N!m�%W���	�|�'���[��'g2�
�c��K1l�q�FY,M���w�ift���Y2͘����p�%N�$_R��C����oN������$�	�k��ɕ���:}�F�2�|̃�eK�/J��"d�"f��c��y��ʝ��'�?����?�Rf�2М��4'�+\M��2�*	�`*�6�'���xĩ>I.On�d�<A�����3
�ԙt Yo�`j�PN}�,:�y�'�r�'���'a�3cfԘk���1���a�2K�m�%c���$�<������O��d�O�i��x,��A�K�JM�f�$:-�<���?q���&Ra�DΧ$����I�1�ȀС�k��ش���O���?���?�DJ��<�C����5;v*#����hR*y^���'�"�'�2_���F-����i�O�"���8Z��b#��T�!� �E�Iuy��'�'���K�'@�i��b��@��Y���5e2��3bf�H�d�O6�=1Nt��R?A���<��-<�Cr)Ĺ0t��"�D�ҽ��O����O`�����'��',�ɉ�w�^X�#M�'��x Mџ.,��^���U�@��M���?����j]��=� `��Ql�Q�nM1���:#���R��i42�'�:���Ojʓ��O����ÓA�v )���z��42J�|��il��'�B�OM����C{d���LFL�\�B�E�n	F�l�\r��ӟ��'1�4�A�i��
%y�P)e4?��	o��x�	ß�ɦbU���Ī<	��~���j�L���(���������M����E��?��I������j����3ƘM�����*z���۴�y�I�'#��zy2�'\����ؔYd�Yi�B�g���Ѭ��KZ��{���?����?!����9O�l+Ѧ����A�# IcJ삢��8l���'@�I؟��'AB�'`���2�J5s%��?3����"!֌y���2�'���ʟd������'2p���%l>1�D�Z!R,Ҷ� !o M�j�x��?�+Oz��O���@�O���5x$���o�Bh����(A~�nZ����	l��oy2/��D�2�'�?�v����s�U�H���(�ٙ6����'��	џ���ןd����[?I��D�FK���㌟#TeDe�T��⦅�Iߟ��'b�a�L+���O��F�x{I��Q
t��P[�L� s���%������C�j�$&���h�������s#�F�lm}y��ӁaF6��V���'7�t$?q�d��..XdQG��UN5hC� զ��I˟�8�@�$��}��F^�T\��%��0�p�[1E�Ԧ��F�J�M����?Y�������^�p�,�!땼	� �!�"]`��l�M:�	r��E�'�?YYy;&�I��Z�u�#�c$L	nZϟd����PY󪄗��'5��Oj%)$d޽6a6�
�e��-�X����đ��(�O����OP������h��7׾a9K�c4lZ��P�q�ډ��'5b�|Zc.�,QA�׿:��[�(+J� �ӬOYۀ<O\��?����?y-O��i�*[6lo��2W��z��$2`�� R�Bh�>!����?)�{�\���C�DB0�xk�)�����<i,O��D�OT���<��"m��iZy@8$�\`���B�	�'�2�|"�'�R̎(:B�$'Aĉ�mR5Xl�[��	G����?����?q-O�!#�VM�q��%o�CV�w��/Jfn �ٴ�?yH>	��?I��<�M��fDǇ� �����;j[9�Ԍc����O\�`G�Ts�����'��dE�pXe�'�ީVjzS�"
�Y��O��D�O$��=O��OX���!_b�X��X�9�X����C5t�6ͫ<Q�� ����~Z���Ց��#��YL�
�����~�j�EmӲ�D�ON�y O�O��O��>1;�L�)=�d1ckϫD�|a�!kӞP�7��֦a�	��l���?�Ɋ}�LT,6�;rꞘ)W�A鴀�!T{46M�PZ�*�� �Sߟ�XDM<n��2*ԶE��i"A�Mk���?���M���v�x��'��O�Q�ኄ	��D* �Z.B�҅9W�iH�'*>�yP�,�I�O8�$�O�t(� �1��1Y�C�����զU�	5(0|�8J<����?�I>�1h�н*���%:R��閛"�L��'�$`z��'������IޟЖ'�fIxb"�'hy��3�P�ծԈ�kF'ބO����O��O����O��ڵo��o��-[��1FZ��8%
c����<����?�����$�e��l�'z�@)4�`!pͺƧ,��X�'���	~y��'i�p�k�&Z��8��H@�2	&Ϳ>1���?I�����5"F�%>�Z��I-�pr�	t(Uf���M+����<���	%6�9H ��(j�QT�{Ԃ6M�On���<	u!_ƉO����5V���`g�@*a���v�I a����'p��ܟ��?��\��:gbF� ��$>L�2��'
��%%���'{��'(�d_��]+Ǽm)��
"�U�.��Mj�6��O��ExJ~"�	Y	�v�*�*��EQ��lӔi�0�	�I韸���?A�M<a��I�>�bf�J2Ԕ���ͶX��l���'	���pH��F�V%��/i����i���'!���OH��O��ɗ3�J��bi�)1�}��j�w4�b�$z�7�	ßx�IǟT*�N˱cT�$�KTJh�FmG-�M��Ry�q���xb�'�b�|Zc����@�)�d�C��L�d>�-��OX���d�O��ķ<Q�p#�8At��i�6}�U���:�Δ "����O��$�O�O������Z78��$�%N.~?(Ă�Dpӎ���������~yr��(��S�u
�hx]p�1f�s���P���џ�'���Q�-��!b\�N`�\AS㓴G*���'���'�RU��z�.�!�ħ3�Μ�tG�H�=��W�r#,���i��|R�'�Q��0tnՒ=���P��6 $� d�P��OH�ɐz����'P�toՅS�NO�Ȫ̋��_33�tO��D�O����~*��R:��D�,��M:�#[�E�'��tr�<E�O��O�&�	\&�i���<"P[\)(1��m�ğ�� �#<������'�.Q�`N,�@���O��?��j�+7��"�ϟPt���I'��ݪ�C�Ib�5����OB�Im��ׄU�J��a��M-C6��% ��vQ`�
d(�
̄d��⅖@>��V�P�V�ځ��J#W6f��",� �DX���m��]����)	�ۗ�A�o��18f�ܠW��i�SB��g-r���y͜�����51����D�{�F��<�H�bB%.׍q(yqS���?��?����.�Od��u>�!�B�h/��!��TB~����ߴ-:6�� ��	J��*�"ʐ[*��d
�=% 3c�#i��P3s�3������6*-���D��I�0+#H�
Lܸ2�'�I�V&PMQ6��$��&/�^��P��O��d$���'��,HS�Y(M<~ �V&~Pa�' ��MU3��B�Ȏ�N$��2�yR'�>�)O�@q�NB}��'�차��* �icP13��b��'�� �V B�'��	H19y҈k�\��\Hc(b�\�xR9��8��	`A��ڤ�'�4	U$��DB�1�%L� H����A��-�E�V
rS~��� A)�p<ɇ�����	Oy"�>-�LHұ�бb���b� ��'�{��Z5$�PpQ��&�BhA-� �xBCe�&-�N�td�f�6#�;�=OF�?��A�"T�4�Ig�dcFo�'N�<_x�@�c@2#� 9��@8`��'+�����͋��Q BQ��T>)�O�;R�W7
�}�� �/I�2!ZN������=h�0�C5��J.�dG�$I���hҦJU��Ĕ�é�;��I+--R���O@�}��b�MzdF?јY`VdWx�i�ȓ[V^��H�rv�KÆ���(��	�HO��և��G��يb�ڇr�9��^}��'���ճ6���C�'�R�'��w��|� ��8U�*�ce/\آ$Q��ů,��9�K�Ob���	�1��'�@�V��� �������˘�M���Aqi�Op�AS	�����y�����Y��X��ܬ_^�	_r�j�Op��������I�_\mQ�L8�H!�(�/dC�ɮj�ڑP@�Ukt���f�4-�z�{)���'��d۲>|��r��k�&ƀ.ʄ�Y�<D ���O��D�Ox���?1�����P�{�����c¨�@aJ1<�j%�T�8;XѢ"�� :s�yR"%x�ȉH���1
 ��%�2��˄I� 3��8�dg��y�)��"
��U�]=��dɆ�
�ry)���?y���%��#~-�̓B��▼Jt�f=D�5%��y�����k�X���>����$�<��Ē����'��DV�6TL!��}n�c���1!wB�'���'�'�r1�ʥqw�	4](O� �"a�)pu��j>Q�7�'��Dh� �1NA`1a�/&�1w♄]��CE����qU��D@џ�z3��OP�d�<Ѱ��9Fi�'��/_K�p���<���?������BM�5C`a�-I��ժ�oдbO!��22�TE�)cn�< ��<A�f�\�'� ð$a����O˧[8��p�akPmO�K�(	tDB4O��=B���?9Do���?��y*��ɲnezU��#��Ȱ�+�{V �' �-�����G60:��p�L�$��-⅂Ɂ'��'M��	P�S�'-�8�&<2)��҆�je�ȓ1��Y���{����c�����	��HO��*#b�3n�� qTm�V���Ab�˦��IΟh�ɨ0q�#I�ɟ�������iޑ�N�tG�,��C#��;7�ɐ;�"4`��@�Lf���¢@SD��|&����͔G�&�[�q{�Ja�	�=�P�K�"��L�� ��'V@�>�O�|���+L�ر���h������֦}��П�PM���Sҟ��I��	ݟ�x"�ߟ3}XL�f�&��;GD�Lh<���}��i�C�ПxF�d��A~bh9ғ<�	sy��ɞb|9T q�-�k��u?ΥH��Q�A�2�'���'f~��������|e�D&u_�՘$
��}����&XT�����V0����B7�h9;FN��pf�x� �b<��Ƃm���8F^��r)�Ǔ�9x�(�IN��,S2�׶9r�Q,5�z��H�c�!�dK�<u���f��P=�9�SN�Uh1OJ��>I�AY�0���'���$(Z��cS˅+�,<hF�׽%���'�nd�!�'I��'[BU�oK�=��OP�ąX [����Pk�����'�ڬ���u`bi���J�g-�q��nH3\jP7M߷Z�d}��IBv8�`�A �OX�df}"��W@x<��DMx�XM�M�y2�'H���S�mDy�$)�X�ppҋ�ja�hO1���ll��m3�G���	 fo�.d
���4���ձ8qHqoZ�x��A���ݤB���*<�tmч�S=w_�}Ӓϔ$���'��i��'�1O�3?	F���t[�tf�ɟu��ɒ��E�$Ԉ	���?�h�Ìp.��gg΂8QQP��*}�OΜ�?i�y����3R�2i����^H�x�?�y�
ހ<�r��tHήJ�&��e�ܠ�0<ab�)� ���֠ɄK�"�����z�f�����	֟��I�kV�0
Ģ�џl�	⟔�i��b!�W���:���k��5G(�@�H�Z���	~t��)Q��ڜl�b(�<1��XH��+<O QaN�/{��9g�֪r'����!�	�p'����|�P1\^��%�/I�	�P�B��y��]���q��8T-Pʀ.��]@���8�s ���e$���$ �dH�� V晙{ڄ�A��O����O��������?a�O5�Pp�K�[�lܛFG2�0И !^�dD��'�����D 
�(���=ŖLTaG$f
���'
c	�2��񃰆���ܡ6B^:�?���?����$�O����R��*ePԢq�6M�lj��;D�����O�����)M1���v6�ɥ��ļ<9U�^�Jd���'!"��>�(�@���?`2�@�d��N��'PT\���'A:��E9"���a�Or�Iv�K5J��\��&%`Z�u���'���1b��d��']哅��9Dɠ=(��!$���ǓJ�%�I����ן,�׎tv�Ѓ /YVoZ8��_cy��'I�O>1p��Z1�����)�v���=�̋�4V���g�J�m�z]�lU�@mϓ����󙟰qc�2�D藄
��D��7D��rA		QV��:��ɑ&�@�(�6D��`G"��H@�)8��E�|�ZX#4�2D��"
�����D�_�hXc$�2D�̱fBD?z��4�A͈�\`�8��+D���A�K����N]M(�l<D��J%�M5 �(�80�ʿ�y�d"/D����V��d�6'�
8�y�Rc-D��8��M+���hCJ��1�Xe+D�LC�N���d��D�>>���� <D������!�:�,سK1tՑ�7D�p�B=u����tjȕhj:�!��3D���@B��� �3��*s�8�҄	3D�P���k�l;%J�r��u�e<D���QoΆ6��	� �3j��YX�*(D������$���ΈV"l��A&D��E�� �z`��HèE8� D����0�<1���6T�ᱶ�=D�4����4h&>���c:*��PA�<D��!#oT)0~v]!����o$ۗ	<D���(�>]��K="��hp��:D��c#�8e%�$9��Ƿ+���f�7D�T�wN.( Xe
ı/a���0D���H�!3zQ��h�71�-�&�.D�8C2a�-=KL��eǀ� ����֢9D�����Y=71Θ���:zk�"D�,B6��^�љ8H ���*D�����ǉ
t����K$��ى��<D���P/���vn� I?��c�K6D�H�cNق]-HH��J�jR�9"''D���6���MTp���b
V()�s2D��p�X2԰)���k�́&C#D���+W�`�rIh�兴(a���	#D���V/Z�B�Pp�?Z�(tg.D�X��ñ�X��F�j, �)D�����M�R`X}R4-B�_"I�N(D�`z!K<� A�-Kr�&����0D��C��ɇ)�`�s����q�P�R�<D���ԡF�0�8(r�Ѳ~8�+�k<D�8'�-$O�ـ��R!w�X�*&D�$(uo?WS��D��'U��;7�"D� �V��(�~��À+��=:7)=D�0�æ�R\�ɫ�@ ���FC<D���oA�P�� �SO]���'D��	�G�;5�X)G)O�68�AH$D� �%��@[����DZ,��b�=D�� 0�ZU)�5Dɳ�.N8(���"OTE����d�6�{��қ&T�b"O��Z$�Q'��IS�B�t^�)@s"O�ݸ@�вp�,��(�*C並"O�}q�&�tPAf�Z�"Ƞ�QS"OʍZ���l��銤�ġ@��|rt"O�5A�7h%>`��U�g�l�#�*O4Y3�޾71�i���	-66��	�'��ݣ��Ц`'R���jS�E�
�'�Vy��(a�^ �c�X;
�'(1��C�&��܋��p���'�P��DA�|Y�=�S��!,���'7N�+D*�.T�rq9�D��u|,���'W�m�&�U��r 1�͛bɎY:	���ɂsb.LH���t���f�K�<��kK	 Ѷnǅy9D����J�<!�@�g4^�
6���[�Г*VR�<�W%s�c�P�h×�QO�<��FK�	�	��F����M�<���7Q�2���OU�<��� SDQF�'ME���5�h�y l1�$�S��<$���"O��D��<&� }�2�āE�,`� ,D�,�#�	�e�)��,  ���� �<#�:x!CN�D!��J,z]��e݅-�Hd��GݓsQ��ö*�>L��":lO�b�L݌-�<u�1�+X>�ʕ�'�p�X+V&��6@A6a�Lx(@쒛>\(�G��0�y�Ӱ��Ƅ�29T<ѷ�@�(O4A��Ҳ�#}��)����I"f טR}`���
�f�<��!�{����@x�Orp�7��2+7ɧ��Ҏ<r��������0Y��2dMڷ�ybF�\YLp�#7��sk:�~�J�$H����'.
ѸSHU1N� HǔF�j��[
1�Ѭ���M��l3;���%��r�q'ʒ�<���* ��Q�U{��Y�A�R�'L@�F�(�>i��+�1M^�/%���z��:D��&� s��=Ҳ#�i�
mH��zir(r��!��S��?I�V;u������K�p{"�m�<Y"I=�����9j��!Ml}R�F�z���Q�L^�`�gR�f�	�v�K,-�ɀd�~>0��'R$҉𙟌K�,�5K�e� g��lL:)�d�%D�L��M�c}�824)O�V�,�I"KĶ~Д�qV'�!G�����@f�\�Ƣ�#>��0����(5azR�`r�ܐ�I��y�j�	��Q��aK���0���y�N����ЂBG"n���`+���'����+�=�$0����M6?�U�@S��)��Z:�!�䙇� �����g���H��R�Dp�Yxp
��n��	�h��"|�'?t(a4Ï/hR�c&�t4�@R�'r\�Q%#C=_�DU`����j�ƕ
��Q:"��%KU�0>1�\�֮�C�5T {'#}���awɛ.���ӑ��x!p&
2�F!�Ί'���K#i<D��aBD�G���9�o��F����d�<扞B���䧝"L�"~Z���=���$ Ϛ��p5�x�<	���k��<��m���=���ݳT������Q~�+ȹ����/qR*p�Å�7DjL��=d�C�	�#h ��u��"$���ܬ	BA{�Z�ljRA#�O���[�l�5[¯ >��8��'ي�� ��z<��'f� ��7g���F�%&�j
�'�kQ��
�ڍI���͆��y2��Ŗ%�D!����D�; +ȨHX��j�nM�[����"O�y��ї+��%�!�S�"�1�W"O�\ZT�1��(2V�e��z�"O��Y��34��12C���yq"O	j��=$�2�	�	�d1�"O�p3����137�T�K�J 3"O� ����ӌy�����6t��h"OF�ǌ�wD�`Q���>
�ѵ"O^��a�44��33@J9$@��6"O�<`Ӏ]�����Z�n����"OFY�A�5� �؂�5j��L�a����yÉ}���'���k7�N�{�gY[ߐYדs)��[J<a��(�f�a��� M+�Ƀ��@?I�#�p��jر|�ay",��R� �q֊�9<є8�i���'���2�D�g���'$��f~����7'���uF .�����Y(<�⌱n��aO/%���MP��N�<AI�u ޖ9sk�����`R?�p���
�Ol�"	^V��"O�T�6�^&nH8 )q��,7���7�_5�zD���V��0�^�xU#���M��W�\��[���v�U)V�����N�,�jS��>�����4US��#Ք	-���%��ȟ�"D$(Y���$��t���1�G�WF��O�T1O���C�4��X$�����?��f�,����,��>;j��!![ ���'=�O���"�?�fu��M�#��� �j��"P��P�����s{�瓽 ;*P�"�'�x3�O4q���D� )����@ҒNm 1���'�R����DyBA�P0�0@[�|�� !b�( R�Ǚ'l0U��%�0L�cV�U���3FC��	�g~"g�e�T8��I���R)�� ��g�¤P�#�<���I�+B�FQ���萳
��A����1	� չ�A�T��FP=Tz0��B�{�$1��EU|�`�T9�FM6E�U��� �fy2e�$��ux���gض �I^��LSB�|�  �y�>pC�R,�j-PTC��R��I���W��֘kvy�dI�M˖3Tx�4�G�%�<A�&�O����
��O��JU�,qV�5(ѫ�zN.�KJ�Dt���FjX�\ &,��X����������ֆƲ;�D|�'���&9"�lˎ%��AĶY�hm��'�v�*�o�/�>̐Ac��Z*O��P.E;5���ԏh
ѓ��xR�_���#ϳ@�ʤk���#1]��7U�p�IR�h�1�;]�I�d�z)��!h��[S��ё������
Yy�'�����ʸ#�̱���Wa䐰q�[�ݮ�9��
l\�pB;g8���fXTa��.��I�r9��O�cE�l;��M,L`�����5�
l�2,�b�O�)��Hj�B��h��d+�b?�W@Z�7�ĸ�|�SHJ�w*Ĺ�A�;����҆ԅ-a�!�A��5��	�K�A��7��ir��>rpL#��åz~$�h$OL)1��ar$�$m�\��C�rĕǢ��M ��ە����=�,8r�z2�>Ld�e�d��Z�d�m�h@�!�/ߚG#���H� ��$�s��R�����QH�J�4:�P�k5��	E�#E	�D,$���	�N����cG¢��1R���Y�a�P"ʹ~��-ٷ�Ujn�)�Q�ؓ�`ׂ?ԩ�O���@�Ξ9V���8J	�!�'B��DJ;f���Y,1����­�\v�b�U��`��nO�ٔO���wG��K�<�cK&��}ҕ���h��J�>������\�&D���@�%\�$�� <y��ɇb����:�����ȉD
�GhVW[��d�z�"Ђ�����ǆ��� :�{�@�
������J~䀈 ����T(=�T�'T$0�0�A��%3�H���GDU̓k���hQ#}G2}§@��w�ŻB	� 4�s,�<�a{BHϷG� s����Y�L����E�}�s{Z���w�<ڄ�	!SN�L�D��9�:�{��nވi�`C�_B���d	D�g~f=A�LНI���Pm����
ܛ`�Z��IFkT*`F�2u��0�ԉk3G.�wIh�H�ػ &��r.�1���ϓ}��x�W�~!��c]�p�:4�O��@REך a�tj��:O"����$U�a��zu�[&JZ��hte���$Q�׺d��M���6�:�$E�!B���DK(l��H���;W�x�ʧ�Aަ6�-�i���'uz�"��	p��ɕ\	�U��L�'���`'��wL�U	�X?Eځ��dؕ��+�H�֔a�Zn�&��ǅċKY�� ���)�:D�'�.d{2��i��9i:E��g��J�d�p獦R�HB�̄%fؠG|RKY�,���K0	Ș��Ox�+0����$�2���V���>�a��7n-2�A�>�&����D� 4����R��ΐ T�!y����O�$s�1$�ˏ�D.^�4�x"���5�T��'���EZ��E�g"j�X'E8�ʰ��ə�ڔk�	D����b`Q�+88B䉞�v ��BU�>�qB�&jrB�ɓB���qW�Y�o)R�ɻ%nB䉏?|J�P���F+L�K"剋Kl�C��:~(��W=�����&y��C����Ɓs֜@A�X�B���:D�L+��C�e��5��e�&1݈���M-D��IC&\�>0�E��2!:�╁*D�� hYkV�]-F�L

s�y�A"O�LR!�M�ȑK�
ٕl����d"O��IcHM2qG�ة$DY4z@�{�"O�8�7�֊,��L�tcP;�xܠ�"O��h1��2>��tc��t�L�"OD�z��F�H,AV)�~�< "O��C$CV�̅��i�ʡ��"O��H &Kl��Ig�N�w�L�)"O>ihަHPB��0�C�y� 	+�"O�=y#����+��g{�=	%"O�ai����
|���Q�8m61	A"O:iSə|^@E e'>zP$u�"Oj	�n�!-�|D�ϞzQ�EKf"O�e��L�H���#'dR�Ej|=�"ODqx�a�S���#Z1;Gx�� "O��)��� ��M��D� 3TCP"OP��b�ݗe���1���"rl�c"O�䓡g�

�Ɲ؇�Q�al��"O�HA3�8A)ZQ��Xh$T���"O�9����2��ԓ��3��9�"O�x����/	���l�n��9�e"O^�)b�B1�|9�AlD�p��	H�"O
�7�W7�HA�kN��� ��"O�az2.U�n����1@��9ȥ"O<P
m�W�����$�$�#T"O�i���{4$��(�.{жIs�"O,�f�_�Z�X�PG\<�~ �"On�q'&�-`jQC&�%���!�"O������H�G�xf��y�"O�!A��2��J��5���q"O��[D�ΜvL��*�B�@�d�p"O�@�c��#�"�K���!I�� @�"OJ�!�-
�z��຀eېe�N���"O��H�e��|���E�\����ZB"O{��	` T�g�	 �~��"O�yq"��$@��%�;�`8E"OhIPA��ZN�MJa�Ԗq}p	rT"O�e[!G�,|����A�N6m|E"F"Ob`�C'�YxTr���aaXh2 "O�M`�i�2^�|J��+S�A��"O�)���S�?�\�	�fP(O���"O��ɐ�F*7��3�KWIA�s!"O�A�  Rɼ�z��ɪ)F޹�s"O�H*�̑	,���GO�&g�|CS"O�虄��z�i�#�wj�詖"O�B��1w��]/qwj0�$V��y�h��t81�En]%h��H��yB$�`I����ŧ8���q,ܕ�y"
R�n��`"�g\�%F�8�7� �y�a�V��A�O�L�r�
w@^��y���1@�#�n��Cr�k�&��yb��'9W�| �ۗkyA����y��&,����r��	.tF�21.��y2�Ƭr6@u�㎁/9��)�C���y��!@��H1�i̅<ښ�z����y��ի/�t���-״
�`9`��7�yB��"4�}arN�s/�0Yb�Y�yR�?;��̄�7�rtc ��yBd�8���e�-���X¥I��y���-`X�C��U�u��p+�*�%�y�e��t@r2���m��p��"�y���(S�mڕ*�/�vqÅ��(�y�┐-����p&K 8m�U�֨�y��ށqK�K�Ӑ���҃,�#�y
� e+���5(o:xJ�K3�|�0"O]!�9Q^<��`:_HY9"O�4V��o���r ��{��,�"O�=y��	�i��R��(k��-R�"O�,A�H�Ktl����?���id"O�#���4$�ҭG(��x�"O�qKB�Z�� 3�M�~�><��"OH��f��9g�X�`�Ą�"OF��C"�x�d��A��kcp��P"O U�fB�8@ܹ��F�Ab�A	"O��bm���A)�ϩY[ (��"O4��dƂL���0b�W�oN���g"O�*��Z1��j5Z(5�"O<eʕ'�n����f�mq��W"Op��"^�`��#\oa��"O���ˍ7/8��1e�xr��hV"O05XDkP�+A��.V��HY� "O`l G�Z�O�ր�gk1�4uc0"O��A�X�`�:�7a��j�pZ�"O����:&;:��`Z�4&�'��OȈ�v�J!n	��Ѵ E�>t��"OU�G/T�R\zd�'�5{_B��vEH<9vj\�E����U�*����!�\�<���'?�35c�z	�����a�<) (]��;@m�Y���0D���W�Z�.��)��)B,~B$}y�*D�p�G,Ĵ���M �*��(D�XHŃ�4 ��P�$*$���K�(D���7�I<�\���8Ns��(r�:D��%/������e��/r^�8��.6D�T"��7��A���_�o&vU��5D�𚳀�)=��awEI�z�;&�1D��@�`���A8�d�8O�� P�-D����ꔻH�P*G�Q�=g��1$�.D����W�"x:�
SHO�F^��Ō/D�<�")]'��`2`ډ7�)���.D�4��0��]h��يΪd�`(D��j@�n�!aǛ�x��d�,#}��'E4���㜌s�(��6��.$tƌ�'���u�����hp��/!܂�
�'ň�!ʛ�2db�ôJR%g٪\r��&�&����S��]�M��P�ꅾ#���B��i[� zA,�� 8�y�ˉ�I�A��Q }Q���_	�y"��
D�&���l	v�	���4�y� Q)�����bP�!��q�F�&�yb���&pt���m� �F��'�yRIɃG�+KY/E����6Z�B�Ɇn��%8�eN8�!#��&��B�Ƀ�2���!�&p��)?\B�I$n�&-�d�-\�<����\��B�ɑN).���)�Z���F�(,~�C�	�	b�L�A�Ԑ&P�	!���7\hC�3Hx��\6+~$�6Y�5 B�	<s@�:a�S�Ȳ���
T���C�=�@�!ɗ�Q�=�)��#e�C�	�RZ(I`L��e�B��D�͓U��B�	4LA� ��s�(H�a!�;|��B�	�q�4(
4
� kc�0�S�+|��C�I����� �	g���)6^�!�DΣ~�l�
s@�?>�����i��!�D߉l�<(��f�;�&Ei����&K!�$�>lc�`���,|x�i0�ר{V!�d�%�e��Ƈ��>�R��2[!�� �}��Ю�Ƹ����Z��"O2-��NU&02ub&�O7X�4�B"OF]!pʜ�[���3��'t����"O�8�&$ rQ��hg$�H�2"O�XQ�H���HmρG�-1��'!�OQ(� A�6 i�LP#��3�"Oh3��if�U�""�>bf�r"O�,r�*��8�����Z3ZTj ""Oм@r�P^[�Ԫ`�YlՐ�$�#<E��2'��R-	�,F>e�UL0󖍆�q|s'�R�:M
8��CdD��'S����I�Xu�Ex֥@1SI���f�H4l����$@��y�i!�U�
ΉzA�����<N�L�
�'82옔iW� 	� ���ǅ@}L�"
Ǔ�HO�+���<j�MᠧM� �m��"O�4�tDI0,����a��8��;�"O�iၕ�u^Zu`E��<�^d�0"O��A�H����$M!eu�P�w"ODLH5�ѽ.9@ͳtC_�fh�ࣵ"O�%k�jNFu86�R�
�����"O�E����C��(Y�+A1��IbF"O$��Ԣ��P1X� UA���v"Ol�;�䏇mxl�A@x�"��"O�ՋE�X�X�8�em�;|Z`�"O���'��#u1��0�,�;@�z,)�"O&P𗭍a���h���*��ZU*ON����9����Ǚ0@{�
�'p���?f��y�L�2��'V0���ݳ7 �<��m�I4=��'�h\��1�4U���� +�|��'�:�;�k^�nLs�J�=y�&�Z�'�Ry� d�I��K�o��mr0��'�XR��֮��-�`�=Y@4��'Qj����9Q�ll�l������'�",��#�V8�o�%�$r"O0�H�M��+{���F���
$�$��"O�%p �PB/��`�/�+l��"O�3sM�4lD��$�+zN�%B�"O�b"kW��jQ�
'Ol %A"O�E ���O�H�����h�z�"OT����<8lL8Ǆ͋���#U"O: ȥ��|��� �#Ws�����"O��g@�7F�E27����x!"O���6D���6�"g��Z~, ��"O^4�a�J�@�8I����<t{N�("Ol锯ҒAY�@��U�D0	!"O&�3��� 8��v��%9�,�+�"O�A��gֳ0X.Ĉ�i�m�1"f"O�EZ��Il��1�!�_�Si�Hk�"O8M���MNhx��U�3Tiq#"O8]P�"�
/)4�xPɖ�E	�"O����� :�@�a�P6��kf"O$��3/K�}�6�(�Âs���"O��BV�՝nO��ۧ��Bس�"O� �g#@�|k����h�H�Б"O܄��@H) RÅ�:~�L8�"O>�w�vj|�0*1`�L�V"OU�g+�V��H@�ANzp@0"O�9$�%/+D��쏼67����"OH̓3CM�m����#%/b�""OJ%�k�2DLhx�#��	�0c�"O(����/=|�ЁlJ�Ah��s�"O�4;ǡ\#�X�B�ӥMY\e�@"OX8���n������LR-�S"O� X� uHP*���
���c��0"O�q�2�
f�$�aG��,�#�"O�$+���0��V`3A�\�#"O���!iT4
PHs��C�v�St"O�:�B��Tn�1�AQ�"Ol�#�E�~ȸl`G�ʤ;Fl "O�Գ��Y
kD�	("M��XC�p"O��Q��ϩ��My���F0 䛢"O
$hC �&XpjG��b��E��"OVzwA9?x�K*��i��l��"O����(D`w$��� �f�As"O~��e&�RQ���
�B���"O��q$�y�X��;��0��"Olq��_/$̀Lx�FK��\Up"O�5a	�U&��R�H�9)�,�Q"OdY�q��=R,��^r#�(k�"O�`��ض'�͋���$N�IP�"O��`��9]������	;K�D�A"O@�@F"���(���8-4 4"O���Я�!?Ӯ��"K�k��9'"O���mȀS5��b�o�,�lEA$"O�p�`֘D��KvOM!v�=R"O��0�ȏ�d��X��ԇ=`~���"OȄ���$�VH��'��`��C�"O�Q�D�,f��Ճ3�=R`"�a�"O�M��'_�7;1���}Z�!��"O�|2��f�vp�7O�OK6��s"O�)If��&`�
�	�P8D@��C"O���J�<X	FN
1�U�"ON`�pՎu�B��	����"On����+�v�K��ҕS��#$"O<=����9j�:;�R�"OؕQ�B�!"�b���Z
��J�"Oԁ�ph;R���y ���FW�t3A"O�xT��F |�I�6#E����"O����(C2^xaBcgK��T�v"O敹t�A!,���G��/k, �@"O�	)�k�3@v��(w�U�u��-�`"Ot㢨]�F���hծ�X�+Q"O��:�d� �@�����8�"O �2B�4#��caOMj���B"O�����Q�$A��jN2yJ��@"O�([�*��Q��ߍ./D�)�"O�X��.Ϋ+,mAW��&.�	5"OШ���T4Ƅ:��Be�M'"O�� H��j�BK�'���"O��V�f�Eb��#>����"O&0�#@�	!�a�1Ɇ!�m��"O�	j� '�t��ɉ�x���"O��6FN�j�2(���_�=��q�"O&(r���6��T�;¶�Ȳ"O6��L�!jײ-��ƃ<��|"C"O�Tb�nD�4Jj�$e=Xb���"O��A5��93��g�ςCf1"Oڐ[�%V 3G*�Y�eǯn�^m�!"O�P�%�@3S��ѡQ��>V�D$�"O�,�&����0!̸/�䓳"O"Qq�g��l����o�<<�Z"O����'�.!�N`+���(X4`�@�"OƁI�L�8:�h�&*J�KJ�B�"OBI #��8y�(�s��*j8�tW"O�� �
浡�h�JTL�	�"O6L�W؂y-ȡ��9��Ș�"O�|ipd� OZ�͛"���B|�e!"O� �q�� /��@�ݪEKH�1�"O�Y��Yg�vmVOA�t1)� "O�}:���y�p���M�
$,B)�r"O����f=	SR4�bJ+|P�z6"O�t:���(9x8p��aӮb\��@"O��:B�ǂL�q�f&Z�"h���f"O�i3�P$��BU�,vz��"O|Xcd��_�3&��[<x��"Of�`#�m�t�C�D��"On��
A�<*N��v�1$��p"OJ�(#��=t&�s��ҝB$���"O$a`)�D�p.J�!sr���"O�H���]5�:�an��dlb�#"O������S"�E˂Ï�|P����"Ob�YP�R�Bs��Q�3nN=в"O��!6ψ�z�*@��
8~S��"O�����	6QB�d��ɍ�@:Jt	�'[n͊�,�+PU�y��^*'��8��'�EJ'��y�����"$
p��'S�!�Ve�<���g�/�����'Kl��A�(�rܙC�<cr�8�')�ĺ��N\%�eH�-&���')�0�7�\ug
��Hȥy|<���'�
��7�Ѓ����'�ܟnM؜Y�'ɺ) ��͚Y����M��z��/D�,���7�d�qa��"q��-D��!�$�.�4���L���u�5�=D���/(�����E$�E�;D�T8fN�*sʤӡa·-̬� �=D��q�%ؠD��Y�J*�l5��:D�̰�`�/�����k��a�Xu{�8D�h0Qo+8��T�èJ�z�x�i��3D���m_�/�����;bR��0�B3D����ć)j���r&;vD�1D��Sa��Wql��G�����q��<D�苠��� `�G26f|hБ�5D�:ơ�&^�E�u�i\��o3D��4��3e����G"X6���.D����/�63�|��DDZ.�T-D��Æ�Q�a�0p�CE�|p�r��)D�(r����m��M!p�p�,D�DiS�:V��ipk� 3!��?D��*����v�Ѕy�m�6~��=���"D��Hd��~�a��1-���c!�;D�p1����=�>�b!Od��R��7D�0����$��$D?;}��"D+D���B0���5M� �0�v�=D���l�)VeN<)�9{�E��0D�@�!�
X��	#�"!��M��i9D�\��mL_� ��� r,����6D�l��.�&t}롉ӿ�%���5D�H2A'oŞ0X�敊8���W�9D���oD&n��j¯��a��!��6D���Q���UY �;��O�<��h���4D�����_�:��4�M8+����U�>D�\k��ɔa}�aq��!y�K��9D���H��V�� [�eׂ[H���E7D�d U�	G��a87b����)`�� D�lHa�5T�|u$�32\���-1D��j��a��UX�g�/"�B�;tc.D��H�F�=$�:�y�͑�l�:$�8D��Y�Q�U��B���L�2mY7D�����K�b@���E�˩p�TM@�� D�pH�ϾX0�|�����OGDL���� ��w�2�h�i& N�~m� "O��aկ+&1dl�([&/��-Pr"Od�@�̼t�X-*��L/jn\5��"O愨�
K�-��	(�,��b�8c"O!xs��g/��3Pm�?"5fIZ�"O6ݨ�"\<�(�q�f^���Y"O&A��CE98�̽KP`�� "O�)"��.-DࠖO��9,��`"O�h��̷Q�\��Q�	3�y"O��r6��.��q�@L,mZ�"Oj<����Y��%�Fʾ�9��"O6T�Ŏ�=.�	r� �2S�����"O��B����Y��@����B�"O,x0Ýi��J�h[���]j�"O�m��@E&	~�����#~�\�8w"O:0�Ϝp��r��f��<��"O�1 o]�W&1�҆��B�����"O��Gj�4�A�ř��2���"O�1!��%��Ұ�,��e��"OD�A$�:Z��u�ˁp�4�C�"O�CE�Y�Ɍ��]�C���c�"O*p�&�Z��>�GD)�d+���3�S�)�)Tt��iV�N7�m�'h
� !�îmH�a�c�y�>�r�(O�!�dQ&B�XB$��9��l�eѢ�!�D�L��$�L�N�Ҍ����:!�D�7s��!�)�$(�i��O�C��'}ў�>9���-�z�X��U;F4�t,&D��v$V��Z��TDΣ*��.<O�"<��ɣ.��E���ļ��sF��Z�<�6�ϳu�`� BiN�p� 6�W�<au$�	 ڞ��f�P�jE��S�<�) �L������<�����Q�<�����6ZVPj���1i�V�� Ps�<�F,�'A�4�`�)��bN
t�<6-��GO��bI���#p��{�<�k.6��l�0^d����b�<�e�:6�V�ag,�=�̕IL�H�<QG[+��	�v��1���sQ+�E�<q��r��8���bV@l�FC]E�<��&B�ju�.V;O4����A�<!0C�.Uؖq��cG1��qv�zx��Ex��B�]�T�@FkZ,T�L��#�&�y2�J�_���5�	�M�ٙ`���y���!o��(!CѠj�x$q��>�yr�'HN![�A�:\~�
 HO6�y�Ȼ����	*>8�cP!��y"T:̑BV�֨;,��NC�y�ȫ<[��h$�F �x	
���=Y+O��I&��h��E��'�B���Ԗ6��B�#���ԧ�!+T= �v�@B�ɢ�`�N�6z���4,P��B�IR5�-�A?{�"P�5G�jx�B�	�=�8�Q����	��ݺV��PݠB䉹Pl�С
M�L�޼(�D�q��D>�S�O����5��s�����۟;��a��'�\[pÖ�~2"胁����z�%�	k���%�v0��9	i��垑j�jB�		���Ch��Jl�0��B��C�1l!��2�S/w%��!��_0C�	=sV�i�����R�.�3`�LC��1X!�I;�B�$;���·'Ǖu�HC�I��M��K�0iu��#
6p��D'e��Q(2.�`A��iE�����S�? ��#��֭n�b�z F�#+��!ZD"O�����Os��922JK�	l�	�V"OT��I�:��R�M YH��"Of�q��V 9��	�Q@x��U"Oޘ[��M6WH�����?v���"O���uǽ|�p8FZ�B1�%{'�'��$�=l<�%$��vH�sqbJ%Y�ў�����M����3��yq�ĳW2DC�I0�pk�d�%6�E2��V�B�	�-������L�$oh�2��L�p��B�u�~p�"!�7�T���Xc�bB䉮Okd�a��Ǐ�z��wo�r�d�O��"~��OQ+(LҩР\>�>�b�G+��>I�O�9�V_<.���0�[���E���	l�Ov��"��L/A�`�L��	�'7�l�C�ޜ<�Xȋ@G�"?��`�	�'�^-PW"��,��7K� 8��z	�'<�5+��]I��A�h�1"��ȳ�'����
�t2L���&ЦH00�'�P��Bc��1��1	 *�c	ĥbM>9�����t���R��N�|���t&�y��$��?�����^�b+R������^�bB=��"O�Ij֋�j���R��{ʩ��"O��X��V�J��A�;
 �"O�e[#�L.��!;0��*�6]�"O�I�'ǻa|(���(�g���i"O�-�tI4G�-���&�6l�s���O0�}��N)�LR��6��߮{n�G{��Og>�EM��'�Xg���P�'u(t��jڸ	���ψ[)���'{F�c�Z@T����X�S�0`
�'<^�`�*�H�A�[�J_���']�����SD�@a+�V�d]�
�'�B��*%� ��7X%N��[���'�?Q��-��5���G��	p��S#V�<q@͠8rb�e͘ 7,kІBG�<1O9�nE��*�����.^�<Y�$� Z9�|+!�H�'[�EÂ��Y�<yA��:�t�rȘ�Xm�h�Ԁ�{��0=!g�A(/�\a����(),p���s�<��� 2�8��&G�]�h`�q�<�D>@�X� J	_f:���$Qu�<�P��:TR���7��+&	vd{0�Z�<��V�E2,8ۇ�$\Z��6��T�<��k?(�|+�o�W2��7�@T�<��i�=Ĵ�@�=��@A��Q��0=#K[o�����j�V�%�T˖U�<Ɇœ�d�����!F�mf�-�D#ZT�<n	�]�+��}�~ ���t�<�p���c�^�
Q�<��4�BX�<I��{�P��'���hu�U�<1�͘�=*�uA�ϱ)+�]h�A�G�<�l�k��d����19��a� (�G��0=i����Ԇ�`c�AOL��S!�\�<���kޒ8��/��v�s���Ux�P�'��ej�+F5�ă <GN=*
�'B�(�B0��ɹ�f\�0hhș	�'A�h���4N=����2���'��i󧟟m����ƨ^Y�h{�'v�!��'�� V
��,9J>�-O��$��(R� g�ŷ��0��H�=!��,Ιk���= ��%��k�џpD�t(4���h�(Z�r���*���y"H9a����/��V�|���/<�y
� "���P��MIԋ�u���""OP�V��/9��3,��g\�S�'U���"ڜ�6*	|pQᅔ�2h⟌F{J?= !AW�,�~,�0*�8YY�c�0D���L�$$�qW&����Wg*D��P�n�*��(�u�1�⑫TB(T�PY�JY���B�l�Z�
�"O<�£�)1?B��Ah����z�"Ox�����V �� *Tq E�"OD�d��(e���O��/�^�r@U�8��	F�V,�1��7���@A⛬m��C�Il6�Up�ͤ+T@{b�.8��B�%�u��/�T�Z����*��C�	�5�*��NY�� IMvC�ɵ^�:P���Q S�����W�C��uƚQ�Aɘ�h�b�[����%��B�� 2�����0um��r�5�D-���͚��aq@�I��� k0D�T�&�M�	(��G�Y/��aA�<a����'��@�'��L�H���'ȶo>�A@4D���@lǴm0���ρ�a� �ԅ-D��*w�UUT޼{A��3i𜙩u�)D�hA�o����CQM��,:� 
3.#4��c�F��zQ|�8�nM�&�	�O���'h2T��g�Yxz�c/\:Q�l1�o��pW,��uu�|���	9�V� ���4�	R�����,*���@��ٺ�'�-!0��s�4D��AĐ� ��!���C215n�R0j1D��ڑ.��YS��򅕁^VV��e/D�0�U��a�tm$ ӃI���1��.D�x"Ui�O�ؔ�7\�d�v��<�)O �O��K~���"��=��*�$�j����?Q�'�b1
0��q��E�-�3�x�C���hO?x��_=��@j�I2z�aSmHly��'C8@��(�7G:|�$�	4ȵ��'KF�����-X ��� .�Ь�	�'񂨡@,�4Y츍�pL6s�@���'f�y��]1�hrH�/�谸Ѧ%�O��	;Yl�����& � �P�_<�d�O��0=��D�	%"�DHP*�b
�!"��Gx����f�ɟ{9�ӓM��֤��{��p��ex���	�fI0�T���gN
B׈B>`����r<���'���G�T�>��p�qlRF�<�r&̼9xj�P����PP���B�<Iv,Z7#k}���!�X���[���G{�OD�O`�3�aZ� ��*e��L9��`���O~�D�OP���7lp����F>p�V����D�zm�{"󄜽5�✠�)��-�` h��?P��2O-�3h)?f1���N0���H��'�!�$�RF�����+�ؽ��셽QG!��Y�n�A'A#6�0h.׷M/!�>7�B�[u�]&��٠�ّ;��{��_!_�d����
(�؅y�cНu!��G,T5�<�!*@1'LF�Yp��V��y��	�B� $��
�&h��T>{�C��7FƮr�&?le��!g��{���I~<�C��87ڱ��&��3kTbŊ�x�<G�XI̬
���S?�ԙq�Hp�<�gbW���cԠ�)B��a����q�<QT-�,w��i��ߍ)ծ�c�)�H�<��O�
Mi*���D�?`��ab�A�<�$�P#P@S�i-���� �A��lD{��)�65!vp�G�Ȼ0^���-?�C�I�,��X��X�J�p<I��+
�C�)� �$�"�L�z�d�5B�)z�}��"O0b!eA�(' �r4���Hg6`��"O�<���Üw�
��Dc�`��C�"O�����zOj�9%���au�p�AOH\SpED���tJ����;z05�`��O���=O>����ƤL��:0KZ�*��DX"O�)a�D�Y��2��Ӯf�D�1�"O�S�L6~���"%G[ti.\@�"O*��a`I�:����ȟ�OZN�y��'-ў�Sj�'�3TnΞQ`x(�Bh���
�'�����r�&:����"���	���y��(Y����p̛�44��kD��?����'v�$t撿F��!���
.ƴP�'m�0�[~��,Y&� 伥��'���q$Q�s�P=8!�Z�e���'��8�0#�&-����0��P�"h����|��'81OXy���8y��r���ة�"O�]곪��w��s�oœul�h'"OޡC�f�1d����Ht�a2"O�y`�-�Zf a��1U�dc�"OђϜ�3�.�B#49� ٵ"O���ͬj���]�
�h�v"O���i+@wx��% Ik�"O��;��+s�֕� ����i�"O����3F	R�$Ճ�T�"O�p�o˝b�0Ű��*��x�"O�]@2o����|���A?�4l{"O�$9%((;"X��Bi��[���w"OR���H1�T��Ú?ϒ)�
�'?��s��-W)x��@l�a�<eq��?�������i���:f��Ö�Ƀy+J�OB�=�}����!hR�k�"��a|�@�c�F�<y���0�v�y�H�
?B���+�X�<A5D�x�n���_S:L���S�<��l��h� �!K��䈪"��O�<)5$�!n�ѳD�Yox��TL�<٣��b��sOTVN�y��_Qy��)�'R���SٯfndD��R����ȓ!��3��Z��H3e,��!��`�ȓ(��j�aW:�"��ӷm���?Q���~�vϗ?^:���*f�>9{��V�<!����N�$\��IH�.%L(���O�<!��u���:��7���R�Q�<���n�^�[7�]-&�¤�2DCyb�'l-Y���i���D�P�4���R�'�JR"C�3] d�1��R�,�$����hO?)Y�1�ؕz�@
;4U)�z�<�d��tȐ+W-ZL` �a�<�T�:ÚyW
]�q�@GO�Y�<���J+~�yX $Ӌ]�ru��'�m�<Ԡ/y\�!�Nǣh(Di�	�g�<�$+�!d�*��6ϑ	U|f�ؖeHg�<!t�NO^ �	�h�
�N|9�'�N�<9h�,3�^���.�>�y�4/QJ�<��oN� t�Գ5����
�O�<!���.��QZ���0A03��TB�<17,Å$�E��R�]��y
&�[e�<i���9?���Qf�/L~Hr�B�a�<�SD[$�.=�	��F;�l �/Rd�<y嫞�\�����ڨ����F!�$Բ]��ݱ��Hk��e:GL̛Dџ�G�t��'�������Jc����X��y�J��4�b�/�$x>D�!,B��y��X@e�G)M@�p��FF�'�y
� ֝(�֍����b��>v� p�"O�x#����y��ע{��x@"O��[W��49����"�& ��i��"O|����I8e
J8S�O+x�������O��}�'!�5SG��#+V��S��1��`��'ӌH07��^)��8J_�H���'R�Ĳ�
ثh�T�ƅ��=\�q��'�f�iwj�<z��SE�G �բ�'ٖ��"�A;�����ǝ�*�����<��yr�Y:#�㑊,F��}�OӀ�y2M�h<���oX�9zy�&l�%�hO���.o�n���oGYN!5��6U!�d�"�Z� ,� X�;�*�'k!�ċ ?:���m�:��E a��3hR!�$W0z��GP}���q��R�y2!�^�)�聂SY5[-��!��O�v0!���~ع�흷$�q�/J*�!�$� P���hB�ڔ���1$O_{�ў���	�e�r\����L�X�`f�9{��B�I BI��rNV��ac��[�L�B䉗lܕ��<6=�����B�I�3��Uԏ_M�0k��-4���13f �pC�+n��:c-��|<x�ȓ|���LX"c{F,�&��p#&͆ȓf�֘2&#���t22�ϳa��؇ȓ:T�QuI:�츤I\
\q�x��%��̐���
���Î#���ȓZ�8���V�'צ���X_���Y�Z�#�&D���\�&��Da�d�ȓ7�* r�/�*r���b� �`E��1Ð<qM�@Np��T�g�ͅ�!}�-+V��K!d�*�֌�ȓ"�6����  2u#��v�P���v�dp�3LI�I�X�ꑫڞ*�PA��wJ�����!V9��0��R�����ȓ%�������TY�G&K�
R-"ړ�0<�&&ֺ,/�͹w(]�
��xpg�C�<A0M�p�N�kP� ;�t�%�UB�<aW�[�R�"��2��:�D�B��}�<��JؖT�.(�ţ��D!0�gd�<�e����&�|{��-_`�<!�)U�[(��y𪇈1�n�ۗ,�e�<s�}44*pDZN������[�<�FM�	�(I�F��-W(��d�P�<q��Q�t.�Q�g�+krL���_r�<�ˉ�Vh�!D�, ���l�l���0=!� ��8@"ѵdSj�К� f�<�aN�l���B
Y�2ׯ�k�<)��^$b���ˁfnrБ�j�<��jΪ���������cD`�<I�"��8!����Q֊�@�<��H0]S�ݓ�.Mgd,X��B�<I7Dٞ::�<�t,��0�9���FU�<I���0fz�82��Ձ�6��H�O�<	go�j���RCͼH .uZ£�r�<Y�A<(-�\�Gȷ&q�mz���h�<)�1+��$h���2]�XM�n�I�<1H�
���B��K�K�<Q���(��lC#���.}�d�q.�L�<�uE !�X�ґи�H;�͓ry���o�'_8J���e7�-H�h��Y��)�'�����Lpk�H���%��c�'��i�g"K)耩ю�$d@Q�'������*`"5���[v�K��� �4@Ä7.�$Ցtm�&A`"O�Q���{vd* ⚒Lβ$��'�T0C*�$�`/R�^�U�v<%��)�'��q0b���  d��fg�a�j��'�jÙ�U��m�6NЅ(M���	�'�������#3 ���؄KL ��!"OR�S����(\�za��A�v`���1LOr�ʂH[���3�NΑyL���"O���C��Mk:�е��$o���"OΥ�B/��T`����АOSD$���I~�8� ���n�Nh��+�h ��o=D���p��_� 
��*�, �s�%D����0p�F�s!�*:Q � Vh6D�ȫ&.Ô{�����R���v 9D����B�Z
􈩠��DT� �G7D��*�� U�|j��R"�yp#7ړ�0|Jկ�/�Tm��^�}���
�ǃf�<!��-/�
�Y��G<#�\`aV�m�<I#�!Dv
!I��H���:�B�o�<���ѿJ�Z4��&5,d6�7�Aj�<A�/�x^���á�(C�cc
�c�<�Ӄ�<�!1�"ʚ�kǅ�y�<�!k��@�p�埛=�J�c���w�<��FĀ1�~d��ހ(:��@�r���Γ!��mb�ꕏY��D�"�3�ج�ȓ=U�(��O H����M-nXQ�ȓ~H�-���+``2)�'#d(��ȓM��x��� �h,�f�
�}��4�ȓ]��G�|�`|#Ō]�+P �ȓ_	.l1r�Ҵx�S� �Y� �������gJ�I<��"�՘A� (�ȓa���XP��Cw)J*AJq��?��Y%]!�:u�!{[ (��_ ��bf �?.��59׉%�)�ȓO���1m��f���Xv�E>B�lI��o \�Qԇ�@ Y��n�N�	��B��0�&�"5�Va�b�>J��H���pȉ��0���[g���`e��g(��8��;���!�Z�$�C�I$���҄o��`+�ř���&MfC�ɺ	bA����f�6�ش�I�7*C�ɉ]vv�8���
c߾-;��]�n.�B��Z#��� CD�*G�Q�]�.W�C��xJl�t�e�r<�L�3�"O�`	�C�B�f��[�8�ز"O��z%ظ��ݻ��	|b�qc"Or\�$�z�)�BO[�dy���v"O��k%�O]p�̑��Ƚ	�I�"O�8i�	F =�P&�5	�r��"O����j&j��m��+O��H���"O@m�&����ݠ�+�=g�p2�"O��3F`8	�LBŉ�2b� ��"OJ$;�����rFB̾n�ܨs�"O̵�Ҍ: ����a�,#}�pw"O��H�a�@��IFbM)�"O�,�cS$%��E�u��<;�1�5"O���We�/�r-�����'CF0�6"O���6�:��J�v�i[v"O�e*G��6DS�H�K�����"OT�X��7��%�'Y�z"O�m ��(i~��S��sX���"ORqI�*�F�Z�95��'%��6"Oԍ�E�Lc�����`t�e��"Or�@Q�"l(�#��g ����� �E1R��!�����<�јS"O�0����FjM���?f�4m)"O�����:Bni��aE��$��k�<b�.2"깱ա_6K32h��p�<�A�	�su�<Y� X� �DD�Љ�o�<YΙ���8˖JŦ ����e��l�<ye��Y�*V��"~Tf���ml�<Y!ĂZvјŅU�N����bA�h�<�)O>zWr S3̓�\H*� �oYh�<1�-�>�
�sŎ�67@�h�mOK�<)�"�Y�b��X5e��@(�O�q�<�3��E��`��FE"i����`+D�PӰ�� 0���B�Gʊ��F�)D��zAE��/Ă)R���x�
T=D�p�&��7����p�6;N<Hp&�<D���M�N���3GIY�F=����';D�h�A�rN�\#�&��t���+D�0���K8lخM��?4G2�0��(D�t e�
�F�)$����Fّ@e&D�����.'e�`����+����/D���l�
��8s�o��R� 9�"M:D�\(���c�TH��.�(wy�T#�b,D�P���U
�� ŀ@ ��(D�����]�J?b��gF���:�RgG#D�P�`�S(nTP�)t2V9�R(4D��Ӏ�G�B.4cϟ����ũ2D�܀4��=IV*i�C �7s�5���.D��3Ę�a��ad/[7"�=˧F7D���M�r��3%��QY�&2D�<k��@t$�f��0���S),D�D����4: ����O]�^�@�	/D�l�V��w�&Yj'�
{2$̀��9D��Y��,Z��m�󠇱V �R��2D���c­t�������%��0D�p%P�:��)f	�fD���f/D���cA5$�j�)�Ƕz&�5zb�2D�Hz��D����AX9:킕��"D�����ϲt�$\��J�.y��1��#;D�(FQ�6d�3�Æ<�'#�Z�<i�&�PP��Ɯ5:�Ե2V-�[x�pGx2⃂ �VԘbOcc0iJ��yrjkT�d�D�E��h�&�+�y"��$���X&b�Q̪�ʅ4�y�CN�3.|Ĩ�)(Kd�<�"%�yN�/U6�P��H�/�� Z#�.�y���bsءۤ���%���P�̊�y��6	^+U,  �����9��x� |W����W�-�X{�	Ɓb!�E�>�F�A*]4I|��B�D�U}!�d��dT:4��r<v(�
sy!�$^�u�l���^���I�x!�d^�*����2�A��EQ�H�&"!��I�~.U�H�cd�l����2�!��2]�d<*�bY.nR0�X��T�!���`_P}J�D��B����E�%�!��<VG� ��ֶ��L�'�V�;*!���	&�$3q�[�%0��"�bޘ!�$Q�%�j�t&�<>.���O֖1!�ă�i �H��g�'%R�7�N��!���8%����� .�:p)��E�I�!�$�X^@�1�C<s��p�(ٞ^�!��])��<K��z���aAݟ�!�D�&��1�NG��priT��!�ˑ`
�<3Ro
����Y��ـ7s!�� 1&C G��x �)��8��F"O�I��!�2F*LP��|��A"O��aj<��R�
M���(Z"Oƭ�r�"�*�h��M�^i��"O�,�2��c�h�\�^͌���"O􁺶c�PJ����T�xq� "O"X�6�Cָ�Pc��Ҡ�!"Op��1CVe�2BV"@_��y�"O�p��X0��#ab	=IS�K�"O�ab-������M<��k"OF���8{�9��Ϫ(�Ш�"O���N�4 d���pB��%�p�#"OdH��`2���#k@�a�R�˅�'�!���%9�4I���`���1��ٳhg!�D�'2��	b+�!x�PH�"A2\!�d^@��RB�L�5�,���!أ[^!�dC�x�vD��_�u����UDL/!���<�l�v�Oa�^�a@� e!�d�e�B����?���!�I�D*!�dץ3
�H�ŉ0Z\qj�ř�9!�dS@���a�xl|�J�Ø$@�!�$+&�B\�M?�`��q(�;A�!�d;�>)�O�v��$b�ݲ �!򤏾���
x#`��o^�u�*�B�'��Hy�A�]����R��=滋{�'���U�X�aΟ3M���'�(H��B���+��P�_N0��'H���m�%4E��P�T(*l��'��}���ɴwV��@GҸQD~�j�',̙Z��ǵ)��m	Ă͡^��)��'��a�#(O�\�#�8^�N,{
�'7��뉗M�hY�A	:G�&��'�ڍa�(0Z�A�2O�)/R53�'c&eq%k=xd^|���J+�A�'�<q�� /"s�%�(�O�%��'T�PQ"�N4$I�X[�f��Ĩx�',�IE�
~ȲuH��[�V)�'��2%)�Q�d���9��Q�'������*"x��O�y�*O���!/�T ����ɤ\�X0�'z*1���6�6YCGf��JP�pB
�'1�E����F'��y��֟KJ���	�'Z�����h�	��4Gp�,�	�'������� |�$��E�� D��Y�'���Q�����j�LX&Z�t�'�&�HT�X�2t,�WKߋ|U���[A���G��I��T�Պx�89�ȓ-�J�G�p�@Yf)@P�Y�ȓcQ@������H�@[\�i��Dm�� ���mqW��<>��(��
#�gb�a� �61�C�	��p����
���֌Z	D<B�6|��)Rf  S����&*�b�JC�ɕu�M�����S�*��tjU�u 8C�ɳz0N0���$Q��Z7�0+�C��=;z���L��"ӥ]�f}�C�	7j/��11��`K^��⧝�&�B���%j�B���c#�	��C�	!C�`U�d,X%D�e
n���C�	9������7ɸYd �3
C䉢)�N�P ���{�Ɉ�� �U�0B��&U��E3�G�JL�t.�A2!�D	�tx&I�`�\�vW�
�!�D+IW
���G�C������C�H�!�� ����
ѩ9�F<�2G44���"O 1�7���4\�
�%�����"O|-h�EۥC��L��㐧+��0��"O�
��О<ڼz�L2���"O�l���l���Y�L�e�����*Ol1 %ŪR'L#s�A,SzF��'��8�"��
 �Q!I*B��A��'"(q���S�Z >$A҂�8*x�J�'��H��N�8�J���+({f���'��mK�N >d�����ğL ��'⊉����� ���A����'dVpK��@�
�Ԓw�;��Q��'kF\C���5C�8(
��-� �'b6�ڰꑲj��Eb���y=���'�X���>d�Hj�g�5x%�܋�'�
,�Fʎ�z=��dôi�p�B�'�,[��]�TnBl�dIWx���'5���T�p���!פ�B���'x���ۇM$j ;�õR<�b�'�^lB��=w��cmыO��T�
�'n������ g���*LSD
�'�(0Zd�I��¡���ZO>��9�'*���Ȩ$�����_�H�%X�';Z(c�E),�F])�FA�2b|�i�'�|����0c=д���D=}���y
�'F�� ��
���K�w�p	��'jVTYq�$P�zc��@����'5�0RR�
Yb�I�r,�=H�#�'��TS�c;
Z��B` �#����'�(���X� v���.����'-p�Q�Q��dQ��[�&�����'}���I1�	� �͉%}5��'Ϭ$�3GC�P(�b��_!�b%8�'K�%�0a&�@)2-�C�D���'!�L���Zo@a`E9^f�:�'Dx5E��"
&��MEG@�-b
�'N���jR"�*�i�5>=(��ȓ�6}c��	=�V�jPE�X����R3�� ��Pށ�&��af|��|�:i����*S��w�_�[��Ԇȓ/,��ߨLB6Db��Ѵ= (

�'H��t�x�� ��ؔ2�8D�xZ5��`�:v�\y2�����6D��A╇h�RљV��>3�$��4D��x&E�i�ء��)ȳBd�0�/D��8p�(`��Eaqg��1�hy��y®�Vqh��4�$^�Τ�����y���F��d����G�|�(��/�y��X�Y�$�5����2��7�y��̓[��-jʅ�8)�� �,��y�C�T��ZDg)7��{5ȅ>�y�f��2DC�iK2���j�J��y2��:�Yӥ�:��H�dT5�yr�=����QN�	cj����0�yR��>���H�HJ"��O�m�<A��_#w6�c��c"T 9�Rs�<��`d�l �dE �G�v�P��n�<�3��`���._�Yn�``�Ln�<�r*J�_��y�枇}F�pC�Jp�<q�_���P/� n�(
���P�<��d\�@F|���f�o����^P�<ɒ'�>�2�*�=�2�lw�<���?������X"乓"�H�<��jۨA�U!Â:*dᩓh�D�<� �-��cV��y �lq�0	�"O2��H�:F����'�ڰ'r`��"Oօ�*�N����r���3<T�"O�`�P���x��Q
h���"OԸC6c��͐�ek�;[ҝ �"Op�9�������\|¼�%CF�<!�N�mJr#f�Y�,��x���LE�<��/��#Z��;D�K(����e�<1b"p�R��$5eJ�bC�CIa�<���C4R�ЃZ�r�M#p,�f�<�q#�0>���6��"iʲ��e�b�<1���5:B�9�
K9��c�#@`�<Q�&Pi��5�'͆0�M
#TZ�<�#��%v�6L0���[H��d~�<�N^�8���Yf�u.$�ąMy�<���8O�:3@EE�EȎ�ȡKy�<�c	*hdΘ9���j�By�p��j�< JZ/JU��rD��/���j�b�h�<���� ,6l�⧤L�_�*X:H�K�<95&�|�\а�E�B����S(F�<A+�+K�
9 �M��"�ʠ���D�<�++�̪�	'FSrݹg�A�<f�^@e+� [8v�v`Q@[G�<A�/�sk�<����v6�����}�<�Lb��9E�B�f��}Y�EC�<1	���3c�4{��*�,�s�<�
ƱLO��a��qF��r Cp�<�$�E�:G����6��ڠg�R�<����'F�y�\4X���XF�P�<ɐ�A1*��HBd#�4{V��L�<a���,�h���K����L�<	�h˜a�)��I�>�"���N�<���B�I�0Z4g����w(�p!��ؼ�"p�1`�HB�CvJ��f!����NQ� � �nG�svgµ;Z!�$��` �1z��N4H���f�7�!��߼Nqt�xG�"jͤ� �CM�S�!򄈎��ق肔<�8�yP�Qs�!�$��r�r�%E�7���0�E�\�!��1�H����&�D9�AH�9�!�H�K�h\;aoس�d�{F��!t!�d)8d9s�C�Cv0-�d2\!��Q��9��yu��qw*�5>!�$=j@&`��� "B���U�åA�!�$Jw�9�e��P�� �G��!�$Ȕ?kJ��4ƂS�,��$MIA�!�D]!-n5����c����[�?q!򄇿l_
��*�.l"M�P���!�D�]l8A�Cd�sŮV�L"!��נ_��5z��'�����\�x!�DL�"��q��e�2�q��Ȅ+�!�ƕB��0u��C��|Xf�ֺ�!��GP�J}xCk�b�ި����>�!�d�(�p���hXX~~,�r�uy!���()�!a�Ou��0��'{!򤃦>�<ٚ$���R^������l!��Im'N��8P���qˎ(`d!�$_�|r�и�GʻnK�-�4�V�+&!�D_�,0x5��`�PX1 	N,F!�R�^�0�E�G�4�6R*!!�		q����� �G4�|�R��<!�٩^�0�8�LQ�1������
7�!�d�3 H��97%������h!8!�$Ѧ^p��c⟖#B d����)@.!�� �pY�`R�q�,9q4C@6;�P��"O&�@�L�#�84�)�l��"OظJ�ȎYF�k4�A	=A:�"O���d�Z�I�I2�@M� �,+G"O�P��:sgd���h4~���`�"OrrAc�4Ş\Z@H	�p�@�"O�h�A��<}b���%�7�U"E"O���H)��ȠǤuٸ8{"O�hA7��U_� ��đ*�����y��>�2�kB%����r�HΜ�y��9yH�d���(b��o��y�@A? "ҙ�4h��"�q���yF�&f3���6`޾oM�)J�&�yB �ڨ`S�K�b�޵Rì��y�J̙4�4��[4V��Ie]-�y��-V#�!�rgGD����I�yR�W�|VƄ 1���K��-z�Ə#�y.�*�Dq�!b\�G `'��.�y����,d�X�m�)��:�J��yR�G8k  Kw�޶7� ��߈o�!����U�Cc��h�`��j�!�Dђ0��Ec��֟cl�9�.�"e�!�J�D��9�"��*k4k�l+�!���"=���L�"�I?O!�$��|�\�Q���u��)�
�P�!�����!�p���2p��IP��+�!��1A3��j��FT���4#�]]!�dG�֭��C�F%G$LM!�dΩ���J�e��^�4,㲣ݔ&0!�䇈HP��� L�h��ktb�$X�!�d�.p�\�
��b��`��"�!�D����7�1��9��@Z�>n!��A�����B�W�f��S*
/>!�dű^�X`z4$��k�T5ZQ��t�!�\�!~����@MYG���g�5!�d�	�&��4`Y=_-*�S�ژ%!�d�n����4����
�� "R!��V)&:VĐ�C�b�0`X�&b!�ܢ�ڸ0��@����@��W�a�!�d�|Pb�r��]�@�~�r����PybOF�
	p�K�O�Bn��ꣅ�,�yB��J��;��
h�Z����J��yBiXI� %��ʖ�D4���I[��yR�^s2����A��4].�y2m� '�P�q�@U�S�J����5�y��W"B5jy�q��]7 ��ا�yb	ՄxN � ;Z��`��N ��yb$Ϛt�j�˧�	�.���h�
�y���<3�-v��>6�p2�é�yRZ�B�"h��O��&u�E��.�8�yr(��l���уKŤ%*�h37f�4�yr��C� m*����h`$L�$�y�ȝD�,Q�U�J�����f	�y"a�-E����:ChÃ �yB��$�ƏQ�3��8t�
8�yb��5U&�ix5		//䌄s"����yR��0q� n�� ��ƙ�yr!�\��]���'Z��寏��y�b���xA�'�ݚTyh����B�y2�_ ��= v�?��a�m��y�
Y�U����K�9ް{"���ym�M6��K�c))�R-��&+�y�L	m]�\p�V9t<Y��O���y��4Πm#f
�=w��1%�U��y
� �����P�9h~�rA�셁F"Od(ꁍ\�m,THz��ѓ4��*%"O�1C�L_:�tU��-�-"�p�"O81â�B5X�xU'�jl�r"O�X���ܩ�jA�ƥ�'�A
%"O"�u�OS�"��0y��{�!��	;<@��N�(.���l�8��y��!,���"�� ��Pd�ֽ$>�B�	pd#�Jl�	 ��R�!�����S��(S�.{q�C0h+'���=:(�R���${�jM�f�*F�ф�Y�Rp1wk�4a�<Py#���DD�ȓ6�����N�N���ؕl�d���'_R�kfE#6pz�8a�D&!R��4�hO�SG�H���X�D�[ct<�t�J�W�ȓ(�4la����Q.���!5��Gx"�)�3�S�?��S5���EHCd^D�<��Jm�`t"�(C��&'Ʃ#Q��G��'�N��J�+K�N�C��؁=�65��'8�8S4ğ�~� -��ɾ3�Xܩ
�'id��pi�(4�H�w�	�%LdB
�'�h`�Ԩ���4��fU�g��I�	�'�`,xd��.pg��#��J3�\���'Td��h�?6����F���'t�i�V# &U���8g-�!ƌ�I�'�)e-�5~��=ʖdM<Q��'���N�Ā�a
1{c����'�Eq��� #+�0�P*ñq�th��D*?a��)@3Y�P'��HN��2n��K
!�Tk!\ey�&�(eF��vj�
g�!��5GR�p`�D(�Z��QL�?X�!�D�V}�BAs�tL1��_.s�!�'$�q[)V�	}�$���"�!��
l�f R�"рt����Tʀr!�$�#D/����+
;[� ��$
�Ee!�ņi�=��M	Ep �k&Zj!�?.hM�r�F�kRz z�ѮXc!�NHTaHq`xP���JD��2O�x�%�oh5�ޡ.N��""O�|YD�6��u@��zV�(#"Oz��Dj�u`a���	0�n��3"Ox���S�:���`4�D@�X1C$�O���$

c��d� n㶱��o@-�!򤎖,�<�0'쐆s�����G_"�ўt��Ӵw�Tp���d#4i�nY��C�;�E��8G��`���֘C䉽+)�QhAn��3;H$�O�#(f$C��L�z���m�<�D,� ��M��ʓ�0?y��L l,���Ui]�QtX���NeX��Oz%�'N	������|���"O $2�-[�:�,��Q;�,HB�^>u 4J�l�@D�s��7Z}�aL%T��r1�H�u�"�!3�;&�2,��<O�㞐��I�~W.y3%ŗcC>�s��۰�R���1�$�0�8�PA��)8 �UJ�
��f
Ob�{W�ѷ�t��T�֢0��M���n~"�'01��8YqO	X�X��܈:�:����':���z��=��H���p��Rdr"<����?U�#! ��鲲E�$��1�F'�L$��d��*-�.���)�uKx���c�>Y8�Gxb�'��l���&/�DJ�(@0I�����'y�"=E��+�HT��D.�� (�P$�R��y�`3Z��if��Kz�\�^�nM���@�f�<�~������T[��#{� �o�r���֧� �m�ԭW�V
Ir*�CM�i�"O��X���<5���h3^t�P�'�9�'�R,��/J$>���+šE�z��}2�'`Vͳ%��?.��\��#2ǘ��&�S�T
U:%������=g��	IR���y��+/�$�K
��luLt"U�I���<����OHK0j�gf��B�[e��`4�'�d�.�����U�r�l��9�0?���Ŕ�T<kV;{Ü���l�'C�����'iiNX���)q�Q�Q��&L��z�L��&9O�<;Ԍ�H�P�Dyb;O�#~�Q�&H���J���KWi�	�#�y�c�;n���c��,ԨI��拚�?�*O<�Iɦ=�O��I[y�
MP��-|s<]�0�K{l�|r�x��z5�ħN�)�Fe+�A���HOX��$Ѣ_�zxhcg�R<t\�3T<'9���$0��IFd`���&\�1d�5*@!��S��a�C�
�
܀����_=�	S}2�'�L���m�:��nS�}D��	�'��X�5�L7<�*E�D���y�e1	��Q=?����K`j�5K3x
!��[�Ee��9>���!땶4��'���H����˖"p�&N�R�����m7!��Ң5�x���AήG�v��A_!�Ă�l�\�Sc� !���D�X�t!�D�ed̜�'��X�:DؔfJ��!�ϫc�R$$\�zn�`9�
�c�Q�8G�tg�?9E,��O� �	���M��y2�ڥ�0\1��.
f\Q����yB.T#Ar7$6Ec�b�>�-�
�'v�F$�#}O*�I���62��1��'o�!U�G#q�[���`����'�@�Z��.���Ԅ�<f��1�"O��!g
)R��� �ڳP4A��'�Q�lh '��?�|8W�Ҋl�4!�	"D� ���ã;� I@VН|)2�"-�D�S���OT��1�Ư ~:!���70����'�6�T`��������z>5[�'n��@!�%J�5�5��=���Uh<Ym#`���S�ӛN��4zjB䉙b�R-�<L���Q�'7����?�I�"�aS���b���a���5q 2B�I%~X!�Q&�>`�'��d�pB�9��,��-�(ٴ��GS�=��B�03�f�A(�QmN}��.��B�ɓϖy��� &�N]�5FO'.�B�ɀ&�
��!�<\�09c���H�B�I qA�E��I��}&!Q��!x�B�ɱ��)����8D�k�GB��B�	�Rh�IQ�K��\�x�R��GC�t��p�����Dh��ǙS�B��̂O;2XIG"OTu�����  $�KUKE<+z
u��������(x�a�>��ku��$"�B�	?zW^srÛ~���[r�V �4B�ɢ��ٱw�׾qK��S�)�NB�I|<1U���Z��8��D7���m#kݝBm�U���!\���'�ў"}���Q1�~� q-�Z����S$�i��Ԕ'�Z����Y�~���i���03ДD��'�ʕF
O��5D�0pެ(	�'��t���tC.�9%f�>R�^�q	�'�C�!צ��JS��?�
����5<OXh
��ԍ%�lH��:ZwEj�"O�aRT�W����s
E?U��ˆ��$\O� X���a��E��}�Q�/z*�)�O�`8�ϭ1#�P��m��5��#~�<�իU�.Vlkp���.��S�I@�<9�&M1yĺ�s&��8]ݠ}A���d�<Q�AȦ~,�\�5J�O���6	��<y+O��d�<�|�'������F�7�9#��O�n��Y�	�'�&]��5.]�Kŀ�^@�Pc�Of��$�nL�+���lC.h�'�W�x!�L�	,�R2�̓=T�@p%�R�b�!��>&��q0�L/0� �bY��!�$�!$*�嚷��I�E�g��3�!���.�Z	�"��O�H��!�<l�!�$bиŨ��ʍ$�~��g�4!�$����
�A9�����q�!��G9b,l��%eӈO܀JEAɃa�!�Č�=i�у���^ �=�UA�	�!�'l���r$�	9w� �6��
u�!�42��X���/\�L!d��!�dU�v��8QH�F�Xu�b��,�!�d�'x-��"D�oۘ(�M���!�$�5r&̐�ܥ=o6	��k��/!�d_�h��BP�G�L�����1!���kԐĉ��хt۾��$J�*>2!�$��HG��b�n�	҈�Q��.j�!�Ą�u����%�.	�� ���F
P!��ڐ5�p��N^�a���XfLĂ/9!��8qf��!1C2Q��\�F*!��șQ(�l1�ꡣ @!��\�s�xف�W'�h����$!�$ˀq���BS'f<qc GH�2!��+}�l���6Z�Z�� ��>�!�%��M����(<�2��6ɋ��!�$D6D�%E喞qe��+G(��F�!��7H�z��?r�1��g��X�!�D�`3V;"�£�P`#F�m!��Ď`Fđ���B�h@Pӏ��p\!�تxy"�X1D;Q�Д����(7q!��e���&�6=�I!�t�!�dʲ�`t�D��7�X��-ʨ{!�DL�d�LT��H <n�Ȱ{0N�?	!�%t�&0Cu���
D�!��έ0�R]��C��O�*�[��H�@�!�D�~�<)2&牳��X8$M3�!�d/&�XMK�˔�.+Ɂ0I<[�ȓh|�ZE�-t8��(�@��R) ��?�b�AcA�pY�GD�23p��<�P��05<n���ɇ;����Vv�Q�$D�QÂ�|�2���@�1-uP̅�;nI2� �8\���i�$�6`�ȓ@�M���X�d�^Y�%GU7�x(�ȓK ڸ����F���E���N�����w��aTK����5��n��*m�ȓ2<+U���nG���gmΐmX`�ȓ5�p�#�!&�h�	QB�)K���ȓ#�.Y�NݖC���@�!C�H�������$�)���@�7���M�\�8��J'29܄fN\�N*�e��G�ԩ�f�"�z��G�8���;}nL�0E������$<U�ȓP�,l0�&�5d���r��w$N�ȓd�J�1`�N�tb�p%-8�L��ȓg�Z�g�1�� @)�OO者ȓ!�͚�O�4��'S�5�f��ȓw�(TCW�"�4Pb��`�� ��t�^�A��0�8��K�9����S�? ���e��AX1 �)�2��P�"Ox̪&) 9�`4�e'��!�$ AV"O��b/'4�D��"%���G"O��	H&+3p��V��s�Jze"OZ)�I6(�j]�� ҥ
y��I�"O"�� ^:~^@��H��#mB)""Ol��Ԃ�.0�Q�EN�7Y6x�"O�y���	�{�t��w��=|�lX��"O4�-�&��P`�B�6��d��"OB�yw������@�:0_|L`q"O
=�O^?6?|�IF�C24ܱzc"O���t��0�0(��8RE�)W"O�@�dCSf�^�@7)�Q?�$A�"Ot́������)�� 0=
(*&"O�i�kJ�i���y�Q�1$��
�"O�8�G/�\{�ܨy�3�"OH�7�ȇ4���.Ө	�l�g"OV8 �A��X%�D
fn">�@� A"O\)B�ܡ$w�ATjҼ��S "O�YBC�v.�q��,����$�5"O\,��X�i������;Y�3d"O��hìݐo�9ô&St"Oc�B-d�T�CU` �w=�,xD"O,���Գ2,�qK3n\�t�n���"Ol�є�x8S�ݝ�� "2"O(���͘�m�h��BK�<��ݒ%"O���C(yS�����Ik����"O�� ��ّdT�A1��ۻQI�,�U"Ohܲ�L��+`��Q�\6xkBD3P"O ��_��И��H5GI�59"Ov��UA�~�b<K�f �q�R$��"Oh�X�F�)�ᥦ��&��B"O�mY��ژ&j�)䄹A�@�"O<+@��3Z����r\�`(�"O��`ㅐ�%�>�Q���$`T�1"O��c�
ͬ [���I��8j&"O�E�Ø�=/��S5(����9&"O�A�2Ŋ&{���u�P=hw�A"O�|�`H�L����PS<-��"O��(h��V��ɹg�S
Z,\�0"O:���-�66Xf���ȍ~�H3"O�a�rI8`zT@�`%��|�jQ"O�9+�Ǝ9�pC6mS?f�����C�d䐋{��9O~�C�O@L� "�-TL�z(��'&��R��>�����,ldi۔e���mFҟD�i��C��I��I�~*��6W�Zʀ���ңA�z���0	�m?�'˄��i���'��)b��ۜ*)��	�f��E(��'U�V&X��=a���xp*��6�vO
�P�U�/o��Ҍ����ļ����(q����ȗ�N��q*�m�<��Q'��F��ˇ��)��c�P���O���D�џ�A'>�Gg���&�g}�t"�0{/����(��0��K}��4g�J��;tF\p���=�M����Gf䩺'�.|O؁�����1�D�2��8��do`�NT~yB��)i��!t���?�qV�]u�FM�&�ý$-J�;o;D���J/­+TG�:M�PѺ1�V�B��Y�r �>y�J����)reO*操��ܱQ4���*��3	��!�,<LlXb�J�iQ�FF�f�����$"l��t[�0�T%��p��3H����De�F�P�0�k��џ<�"��`��CM�8�D`�'�d%+s��?�9��
��t�	�3������_�p�f��
��L�1���IJ]�r�>���Z;1�Dz�Kd�Y�G�?����P�-6��|*Դ����<<rႆY� !���k�R` šL�L�8e�~�����jćRΈ� @� Wڵ�7�~3 (�ēt�.L�6�<L��q����.�J��	�P��A\~��mY7��	n���`��'o��m��_�p9���Ə�8Fy��S�? ��1�-	��8�S�l�X��8��ɚaچ ��Β�7�ꑸ�R�̹	���AJv��%^�>��|(��K?~�5
�O�p22)����)�m2���d�O�]qGe��IK�|�A�q�(�K�qVrT���*Q�-WHm� ��(���O��y�-��W�6Ě�1!�nԛ�����s�L�-
3�4K2��n��	�Xw�X!�0��+�nG���$����`X�Z1J�3%��%,�zr��F�F	��tJ,;'JS�^$�����#��,{�H��w�<��D�	��X�Ggx��D,X�8��Oʒrv�$ �fNqO�B�I��&*bɪ���,{T����OB�%��7q�fy�Ƹ0��9F��GB�@��w<a���!��!��ьK���W@ɰqV	n 5�$�1i Ӧ7�� 1��@l�!���y��R#�S�AJҜ%���e6������{�
��R�|��HXn2:���>R���u.ǀy����Lyb�H�?���M~2��銷��Xe�K��L�F"�`���C��|s����umO#u(h�v�]�Q>8 ��#�Ď�f�vd`2*O��!�/'���3cZ0 6�Ė ����(5{L��㩉��ճ�D�R��St��.>�!�d�I�2���iO��RӬ�!���_2�2 ���5=���@x�!��I�l�������38�b�) n�x�ȓ55`���':S�arI�A��ȓX["L�2��	���A�cr�ȓ_<�T��	:�U�vD�)=�H����^Ԙ� ��-���R�	+{�$���R���Z���'nfx��E�%l#�<�ȓ'D��SBM(NybUkBJ��X�b-��J+��F�����\kŇ]�ND���dA�lT��9u��x��A	 ~���u�)�ŀP�,#�$+&@��K� �ȓ=�
9�re����� 
bQ�ȓKӛԂ�ZO��J�V�.�P�'��x�֠֟N4����@
�	2���t`��,)Vԙ1ի�!{s(�#\��IS"O~��7*���];�HQ)m~n]�Z��C7M�G���%��|*7j߽O"�Q(S&����A	gX�@ �&6M�'7́��&��<��'�.5)��c�>q`oϟ^m\�����}�E�}���@b�`�!��"���� ���[��Ť��)��\�,���S��e�J2Ȓ�X�%�`(��@��G����i��u_HǬUC�&�`$l��~R� �g��bv�g�-�A��E窈 �>�1b��Li�cH68>�p���%�����I�%���beL�C�P��QE��m	�b�b�$��t��S>t�f�O�E/��'9�`���4%-$
�2V�F�� ���,�1��O��b� P/`�f�H�� ��@�l�~=rD��7�<E۴��|�"��N�p��)8z��Y�O|�>��I�2�jex�n��bH�Q�F���<)S�VE쨨j�h�"X��i1��kq*��ƶB
�b�^M�0� ԪŹ"pt$�'��1'�%:pqS�Qe�T�1�ț�s�FT����5���
��u��9�b|��%�|��ƀ�k1�>B�p��9n�a�'j��X<>�C�D�o%����Z(H�k�ҍ=�^��&�XB<JL���|2�X�@91��[�ՔsɊ��FL�S��#P�	�F�$"����$1�=SC� (�Χg�1��e��G}P�z�
�x�@�<q�J��y�B��$B7�U��Չ&|����+H�bc^4yH�0�`�.8]h��t�B�6�>݈P�^�}��$Y"n�= J���	Hm�<i��X�sc�(;p$��,�s6 ���wf�2C�Ka�:`��O����-@X�,ӧ��NAб���)�Oҽ��I�^�
�
v�W�n�,�i���#6��}®�g:`y�&,Ҝ˘��dR1#G2DsS�L��t	AN �ў��lH���8!���$4TR�{�f��|�QI��I1��S�DT&�N8�2�H}�<�����%!A�g#s�G���l�hޓܚ�)�⑲Ctڑ��D�V�OZL���&�Չ��Ӻ
�R(� "O��!F�P��A�阝$�z�X���aa)�Qlޤ}���	"��00�3�4��#�K-|2	�T@���	*!�~������?펍i��G&C֮XBf�̽�t��S��u�th"t�'A��H��%��Q���5 ]Ë��_�Vxl��n7-�
Lz!�~J�i4b	�'NE:4��	ҍZS�<)ԯ�Z�J��)�a��hc��k?!v*�K8[E��yZ��'�"Lڰ�� ����j$t�@9�N�_j���"O* "���u��P�]0O��J#� CѪ��Y�x��t���1�O��3F��Cy�H�]/�u*��`ح8�"����?ٳMȘ[T�}!� S~YgiRHm `��E]�1Ԕ�u�,M��性X�#?9�	�bw�ui�E��7f�Y�D�Sw�'^���w�a֐��oCp�b�^$�`�J� dY�ᡓ�/�����/��Q2a���K�d��� :*�������$�.�TxSޒ�~B�_�[Wf%7�CX�S��l|)E��nJbD�3e���C�	��*भT�V�jVN�uB�u�Uo���⢊�>�z�C��m�Ӎ9�n�k�]�X���_�H4�Bs`;O.�9;�6�OdM�0
��(�Τ)mEy$Ҹ��NågW�"��~�f]�s6�@HW�'5X(�"��{�<�K�����X��D��]*���$���~�.�
aZ��YGD�w`�
�C�+3y�ȸ2�ɟqB��ɁjШ!ڑ �A�F�Y����ʓlF�#���.5�H�I5E>|Bh��<*�OC�X�`�' ��AN�|\��c
�'Cb@RR�*-h <����,kYܜ3$T����ޟ%��uY3�0�'��q�'�L��1��� �vl@�k�i��'�D�(�d�!g��}�P�S�,[����CJ"�O�ԛ�O���0<Q�)ۘN���P�G�|jVa�Se�Y�<�c�R(Ny�0N@N3� A`�Z�<92��O�x���bH�0�V��V�<14H�	Wѐg�.�JLD�L�<� �#ތ�xao�	+�͂'�S�<�����&��A*�(P�����!�p�<)�Oͨj$���[�b���g��s�<`�G�R�v������<����v��t�<��)��)��a�+D�޴�Y�<!�@�T�#�L�"A1^e`!�T�<��E1B�%p����x��
y�<��!X�h'�4�a�S��24����u�<a�h��a��I��l�&�HPa���Z�<��>sG����ǉ���9a�
VQ�<�G#�.5|jt�P$�0&D��� �S�<)��Ԃ1��ɻ#"�J0n�ks��N�<�!@�:�hE���O����OED�<�S`�	aL��GI�_R
f�@�<9�o�%Pv��1s�N�9���fʇh�<�� �>D(H(�&ӠOc�ɳ%~�<��b�=H����j�d\�E�y�<��E�-G����5'c�x���r�<i6��[��Pp�/��Q��L��+�k�<� *�9=-�=�u����b�L�<ї&��	�x�rqH�)������d�<!�Q�N���-�L��#p)�c�<ib�F
'����J��w�Z){cLf�<���9T���Cǀ�Oqb����o�<�寉�F@���Z�,�i��_h�<9��.;+�]�����%�u��j�<qǊ��R�@�"7��KAl�<�'G��cw>(�C�ٷh�x��b��R�<� ��_?�B��,n�[@`b�I�<��"P�9��q��Ff]��!!�X�<Y��\?:�v����R�TyQ�˔P�<�M)}���bN��w��8̐g�<����&���A\/�h �&�]�<�� ��)��s%b VzJ\�a�IM�<�b�SC��St�N�Un=�cIIC�<�jRO\�5��C&{@�h�B�Xu�<y��[+#p���uNڝP��9�Il�<����6<�7�E,~�`1�Qgj�<نKLR~�j�
�L��=�uN�o�<IƂG�V���1��&��h�Uɐb�<�WŃ�B` Y�E��Zz^���n�X�<!Ǧ�� @s�Y+X��r�FT�<� l��QnC���1��Sذ��q"O�Y�w���F������³z�.�r "O`|�R'80�jE�g�:Xޞi� "Ox��d�P*PH2��D�(���h�"O�A���E7��j�c�>��X2�"O \��i��v0:&��CD%x�"OxD��)C"Yk:I��M�$*��6"O� "�I�RP<ȩ�Ɠ�()V-�S"O��Х�ψj)�pJe�ű.d]@"O~�)β^����$,��I5"O���Ł� �<�0��%c{�rG"OX��'�c͜Q(�ÊcW��"O���p,O�f{��4�|�D"O�Ԃ�/��U�uz�M��U݌�z�"O�)q�
�_V�= c�(s�����"Or�a�E�4K�|[��-|��1�"OT����EB��a��kU��k�"O>h�A�[�Yh��%�ʨ"O��"��]:�8\;VD��F�x��0"On������@C�C�!�iu"OE�5�	f�@P�`B-8X�"O�e�D�\�j	Pe��2�D(9�"Or��f"�mଉ�Bꃲ��Q"O�9��ߊEɳ�
3{l	)�"OPa���@.����H�u��]Rr"O�\��AP0|,�Z�ݬ��@A"O���W	��h&�2��Y�Pz��3$"O���$Ng�`RAD��LpFD��"O�E�cȑ�AN�%A�!I"X�"O���яŐ)U�Q���:�c�"Od������UK��١8,�0�"O0�KV���wH\cg�H�?����"O���!�Q�H�B�^�2�X���"O%�aָB�8ٖ�Ҙ�"Ov�HU�š{�ыZ=6I����'��Lap?ED�=�T�2�D	�'��bb.�o�P��ǂ$g����'Ld r�Bؕz����?(���'�� �_;'V�|����--�`�;	�'����g�ɺQ6M��i�� ���'5��B�͟S����)�*Â���'�{��[�f��$�T�D�wvq�
�'g,@�Հ�v��{�׌i��< �'�L�K�3)d�S�]�3�$�'_"��b���{ѲBM�:4� =��'3�)��Z!��C��$�n5S�'&����O>6rp��Ŗ Ҝ��r"\?<����=E��'9��8U�5`d���mX�H=2�
�'��IÇ7��5�4�2Hm�p��D2tl��k��0>�3���}���I��4+q�R��B؞��6��\-L`C0�'�^	v��8
�Z��
�Q���)�'�p�9���cB8`��'�+W=t-��}�J�Y�vĂ�g�Z�O����Uk�c	>x����Q�>�'jbl��DS� $:̛3 ��=/�j�f�5C ) `�>���>�ҠH�KE,��FTz$�h��u���g�Q�)�	�)$bU8�Ȟ,+X�4�G`C�D�7�-	����勛��=yrBPrir�:��)_'1�jH�G���TbI���䗨\-pb�R���qo[N���1�`զd�a���E�<���*�rX�+� ��iR� 8Y�r�n�A}RO�.��2�J�'*���.d�Ԁu�"|1�"L>5$�B�I	"�pDEM��ƼH�IQ�aր �+�7^�`+p/�>i���\>�)�&;�	/]5�#��ٜU�m���`S��?'̘'fqR)M�9:X�Y��Oè8�fOR�&tzL����Z]�l��l�,qB'G�0>�s�_D��]��dDP�Dٺ�˜p}�Z5'&��Jt*V�X�偡o&
��j���3� X8K��C��=1�]c�b�p�"O�H��K�E��rQj];��")��h� �p�ɑ.��]�����"��'\,@��H<�v�ԥ3��	ؠMY'JP�9�^\����wg[W����%�[�"�*0�@ <G��R�
\d�{�[� !�#�^	�p<�ꝸY������2��Pp�Z�'�ԕ˥n��.���xP#��z�)�
]�E�b��cW�B����2S�C˪=kn�n<IwF��Mo.��&�J����V?i#�7hx
�o�t���+cߤ2Dy�A'擿Ax���2G8T�у?/�B�	2<քw�M?�8�뷯Ěd�a�G��Ĥ�aߥv���LD��ýM���K�O��!���-F��q�w�Q�<��'"]X�M����o��`YRrhX�gH�ъ�`?�V+�E�B= � OtA���,_��`��Hߕ� d	��I����O�X��d1�����5kZ�(.0�Ij�Y�*2�5��&J<	t�ǧP�D�gO�!h;�=:���x}�eJ�y�Q�A\��ۑ)�([��3V�)O�Z}�������(o�!��=<eH=�D_9� x!Q�ى&��ę&����G!	#�L�S��OG�I<O��9�'R���G��6"�B��7hJ�SS(Q"~�MX%j���O�E���3'(��2��ڣaą#�BA[���
����2˪d@�9/j���a�T�`�)W�
FH<)e�֕i!� `�(���&!�A�<!��R75Ƃ�)k��u{�m33�]|�<ɓ�����P(�'7-�@� �H|�<�1֮Kmt�
��hNĈ4ǐz�<��΃�\���+c�Zb�U���@s�<�́8#�~�(��VuܤS�Ij�<��-	w�0Y[��=��ȇ��S�<�'bKPU>-K���=8���L�<1�Q�2Z�/� ���qg�H�<����]��șB6��*SI�<�NF�&��1�1�&/x*Xz��G�<�҈26)�%��X�?���C�}�<�$I�V�`��O%U&�� I z�<���=WaVIK�!�er>�Xq��{�<��"^�W*2�+Ў�,$�#�}��B��܁wqOԁ;uk�[N���X�<�d ��"O8�5�-48x��N�E:�a��]��(�@�8M�$��|�C��*�gG		(��m��Vh�<p���l����J��];bF���I�%JՃ���g�W&����5A��2o����q�\�5�D�Y�(����I�j�qq�rZ���'��13�ƂZ(Y�vd��Y�*9����
?��)����'`�
�y创�O<3���l:݇�F
N%x.r/���ʄ $l��'��+�ė�XW,�O�>eppꀗ%z *cԥ(��Ġ`�<D�|Kt
<����k���t��!a\w�ė�>�ZS��y�3��\p�R+�:X9�����ԳD����D�6���d�<��Ph�BM�e�`bw�YH:���pJ�QX���/V��K�	�M��%E~R̂�_p�� �Z��(�s�̑�xX�]R�!�/.�C�Ɏc<T��E%<0p�ݙ*��>������a'��(��S�Odb��P����m˖Mͽ(��X��'�:����B%�칒T���ӍyBK�������n��0�M�(1h(E����o TC�	� �n%rQ(�k�!AF�@'/�
C�	Af��Uo��(<�2A/C䉰8�,`����N.�s��2x0B�ɖ.�u�փ�6~��IHA�

sI�C��)<@P�A�{LЭ5Mɼ&�B�ɠp��l��"oz:o�G��B�I�56Y��썫>�J�c�C4+�L�'|Ɲ�#�DG�S��G8BP��5�����D�;/��ȓB8؅#]�x�ᄄ+�2�H>�a�)�:�|�<ADI5g�������;Z����3�[I���Pωt�? `!)��A�2���Y�\. p���1�֓A�P��I-)Zya��W���zB�/��?y�E�Z�zP��)�Ɏ#\0P�ޑ2��|"��}!�dټqq�@�A�wz�r�␟5剕IO���A|�I�V()a��I�����th*fz,8Y� K�V!�� ��K0߹]iz! �W�>��9�'���r�K��"�R��O~Z�끢#����u��鑯D����V��,'����� �ḣ��=[i�����Z�x�����=��̣�'��ѻ� ��{�h�E~R� |�u�a~xe+'�΅��O���WY&����'͢Ţ`��f-ș�T��<+_�A�S�ǭ�@*�Y؟�(�`9{���F�es��+�J�<��a���ﰟ$/��$۴�@����+ùI~y��a�+������Z/�y�j�D�Ε��j's��L㐁޽8����'U�,���eڅ	���%?��U%���*�ƝKp$�$N��(9P�W�6b���Dˇ)��e�c%�-�Nx�6J��.%R���=\�T��'x�d����X+*�E~�h��Z58(P�ł�1�ƌ���7��On��  �����'(��k�|:�����\,Ťd06�V3*�X���HX؟`���y2֝J�HԆms�,3G`�<QW�]�R��Q�켟��c�;P��ʠ���Μ'���cs!R�x�6��l�?�y��]��� �R'v~-�0(�'w��I J��E���!��c>Q��L�ayb�V%�}�Bk��iaּz񡞝�PxB�u�v�{ ���y�q�fLD �Aw(W�DM�� Hp�Ŵqa��J��i��9�:���1���HF'Q����6h��m�ȓi��T R�K�w%�LyW�~|B1�ȓx�����)5���.�.'���ȓg?4\�&Jc!p-�d\�чȓq�MB���#d0�����k���� OX�+�LI� M����J�>�*h�ȓ9��pQT��0Z�h��'�$���Ve��s�&ҟ8Tl�����b��ȓeL�0�l���%lСGmY��h"�{u$O3� �����"TQ�ȓ�xŪ6m!����ȟg�@��)gr��hb]Lݺd	P���ȓ~������Lo��aA�,J�x��D �"��'b:��F��,��ȓt�\8[�)��s�H����#,Td��k7��{���7I�Eb�^ذ�ȓ4���A�N�7{|d2��P�M�ԭ�ȓ�Us�� CT2�C�*!�ȓJ�m����ހyQb@W�,���J���Aܠz����o��5��e��`S]=��i�+���"�ȓEPl@��!��gT20�V�̎��ȓA��R�f� R�("뒅*��ȓa~�"&�c�2a�`bK�5�ȓEɄEy��֜u�e9�o��L���+Ǩ�@���a�"Y#i�-3CVi��=O,��� ���H���X>�ȓ~�:@X`bְ1�|����S������� NϏK�lлՋ�+�~��c����W͆�A;�ً,�0�І�\:����R�'�t9�Ώ�|��0�<a.N6{���0E+6Y��V`̓zf�@�a���m���eD�x��ȓ|l�:�-É{.�S��U�
�:@�ȓop]�"oN�dD{���)\�P؇ȓ�JИ��O�{fDJ��ܤpsP	��?w�U��OUF�9����ȓ}~P�k�l��G3rHYSjI&�����E���2��!��uX�ԇȓQ�
�B7	V�m� �%V�VEL���+�T��%�):R�Y��-r�]�� ]��2m��@���1���H��ɇ�S�? 2��CѰD���@%� v��U��"O��7�
g<�U��G�ƕ�7"OB�`���fYvɺv+ ?����"O\I��j��|X���8@5"OL)�*Ȇkᦕ��$�U��E��"O\@��(w}���K�~���'9�zO<)p«�ȟ�l��֣`׈�rLY�F�����O��Y���+`˛&IY���)�O��r����<u2E��`O��Di�G�)?���4S�ɨ�M�s������<�Ot0�U��=O`J�c��K��h�ώ1X���=���ن%�]>@ ��/�rȨB��aT���T#�<�1�J�Si�U��M~��閟A�M1�A�	-�̑1���H�$��S�`���������>Ɉ�H���&���GY">Ȋ��>QgG�r>��r+.8�5/��(O�e�ܙ-��	�uP� 
$��y>�+f-��|M8���ē,I�<�An�<�F�O�6 �� Gy~��)J#G�r���q�H\���`r(�X��$���{ɬ<
�ǨO��*&�ԈT��t��FϢ*�.�3�"OPT�V@�e9R�0��U�)�6"O	��b+3�D4��#t��la"O�µ��x~aP�`�� �"O��g��	J`�ۣ��C��I�"OرH�c��ip-�	=�uB�"Oج��&ž�
�l� ˖�b"OD�j�����@�Y|����"Oi�R�t?t�A����>�2"O�}23j��Q�d�oެ!�b�"O�YR3�G��*�#F��"G	FD��"O�m�a
ݢd3X��5V��!��"Ox�{f�)$NJ�m�s��=B��7D� ��  g��*d�ä,s�e�T�4D�d٧�ȱ	��Q�ÆCNN���<D�,P!���4��Yy0�T�y��S� D�,;�K�<�)kp� Dt��v D����T,f��A���&1�B�c+*D�L��?!�ip5���X�(%((D�T�G��96�I)��݂]ېY b�)D�D�.�*���i��ߺwv�룠"D����[�p��]����)1v:Y��D"D�@x4*�45v 0�b���L�j|�GM,D�$�T��
l	~dxs�(t+f�C�6D��p�Ĝ
â��c�;Mrah�G'D��x�-�`� <A�� ��cխ"D�(C0��!yL��@"�?t� � �=D�DA��x)�v�Y� �)*�	�^�!�Ve	F-[��i���H�K��[8!�D�I\�Z�ϧ#ɐ�yB ��-<!�!D���d�ΣeŔd��o�H*!�D�7X�*���n������!�P�D�����0D�,�X΄2=!��N$>4	`�.
�~c8��a���n�!��-2�\8ץ׫8�t,�C)m!�D��;��ZsD�'�f�P��ؼk!��Zp��pȭ%�Ĉ�Sj�J�!�$�<�d�`	�]����ֈG��!��3p�a2��Ӡ/�j�x6�%I�!�T�� s�UM�\u3�&�	�!��/T,�AiR;�����D��Py2�X_,�"Cm��8�:`Q�B���yr��B�,��(��7����eC�y�ܠ|�is+-����')�y�)q ذPa��=)h5	�-�y���N�dA��̴$�f����y�mΦB^24��� �wT�`�g��y"�]�H�:5)��&��괬��y�LԈy�5�� �>��|a����y
�   �E���
������*.D���"O�1���6��)�^7��!%"O��s�F�9Vl�2$��n*:=��"O��SAL�H���� L
&S�"O\e%�\?8yB���Y(R(�q�"O��n 0 FU�OςO��0e"O"I��f<к�.Zo!� �"OJ���,�T�Q��ٌX����"O
�!Č[=bT�9R�T"\�&P�"O�\b�G;.���6h
	33f�[�"O�%b��]<tD�A�dG�:#w
��"Od��f�4ola ���Vb�mؓ"O�� '���j�s*�:1[�	y7"O�taֺX�X�3��]OY�'"Oz��������5HT/F��H%"O$Xkp�U�(I�h���4��"O�-R"D�%�����ʶq�ܺD"O�HA`k'&;��7'�"0���`�"O�A��C�X���Տr��ͺ�"O��� �̾p�ޔ�d�)ul4]�"O5)�C�$]t9��)y���"O8�P�k�#��{��ӿf�`B�"O�8
T�ߺ9մI0HU?z6��"O�Q`3��d�J�R�ϵzq�i�"Ob\	�H�G:�5��d�F���ȱ"O橢$�D6F���k��i!�/M)3M!�ė�[�=1,��s�ԡ��� p>!�$�"���d%����G!�!�DK7.����Xc¡�2�N3K!�D� �:` ta�p\�Aa5�8�!�d:bq��9!�8;��%I�Mƙ|�!�� �B��L(g���aN�1�!�$3^�%�4�%������2�!�o���a��tP*�(	$�!�d�X'��P���}����SIm!���p�k�&y��8"�Ց=O!�M�%P���0`v�U��S�rI!�A�Y��a���%Ü���x0!��	~�6$;6�U�)���{�m�B!�$SC�88��3�
l���֚/!�U�1I�M���.e�r����D�!�;�ި�@h�3�CƤ�6c�!�*	B:MZb�Z���Q��b�89!��$|{�)%!��y@q@q䑵)'!��t�(]a���.@D��T��Ws!��A8���"��.-�u! !g!�$�up�(j"�#'�X�0��T]!��U����%C۵u�Ѐ�P�U!�D�+gs�Q�¤X
]�
��4�O�,�!�FQ����@�P��qyD�۔�!��N+�Z�P��M|f�r7!��P�B!�1��~�T�V�8!�D�������&U"�A�+�^�!���Rm��zg ���x�*�7V}!� <����h��HmT�h�*R�F�!�dV$�� )�,�D$aS��F�!�S�_��}2� �'/�0���	o!�$P�(���ѕ�M�5�a�M� _!���JC4"B;Ow�	�֥[w!�D�d�\(uDд!^8��"Q08!�dV4f��T��F�@��*�O�!��˻S}\��@I�&��1jW��;!򄜢S�9�B��'&���j#���{!���?8�$���#ƶI� ���K�	L!�� �1rQ� 0pi9 IK>a� eӀ"O��z@E?G���X,��}S�"O�����M�m����a��%��͂�"O �h#�T#ƶ��%�Y˖̓"O��0v�ۦe�B��u�Z`�p"O6�g��c\(��Ym��C"O��tk  Eڵ�L�)_*�2"Or��ץ	'T��Q�Z�}�@ T"A�!�Z,E�|��hUaŰ�B�ᛴ\!���$^{�+��P��o��9U!��#�d�`$-^O���1`@��1A!�d��Aʕ9��ǟpܰ��싼+(��*R��I�L׷:�,YC���yb��D�|��#���3�`�q$�@;�yBG�4!t��)���B�s�R?�yB���8̠p��35���X��y%ݺ$@3�`'2�@9[���yR�"O�Ց�"��}�����
�y�F�� ���#��E4}�,m��I�.�yBH�kW�E ��?#���dN�y/�&�J��Ɲ!#ʰ�ġM<�y2��_��|!�"�P�+���1�y⪌�2O5�c�\�f`lY�dܮ�yrk���"��M����Bϔ�y��ڕ���'bCaC�D�8t!��5.�TI@�ʒ�T֌�q��15p!�� �Ƣm��n˳fI� z2�?<!��`�ޙbg葨21D��qJ�q)!�$ޒ��L@�j�(��[@��I�!�D�m�#��D��r �ݹ�!��F�N���M|��E����X�!�D�h�(�����x�� ���*v+!��	�f�{p����� 
O�Yl!򄑏9��k���+ �r�@R	;:e!�E�!a������6�2��	�a!�[F6IV0mh�ER??�!�$P�U�hg�������e՞T�!�ƫr�h�T�rC� `KE�!�D�Y����WH.x1N�`r���!��/UEY�J�"+7Zl�`�V�_!�D^�R��E����Q~�p����-�!���1B�s���"yl���eY�2�!�DP�u�&|���Z�xj�1
��>L�!�$����m���B�ab��WZ'HQ!��8BX��х��V�5�]-k@!�$J� 1FUj� )*;,�#�� �!�R�-A�\r�ڭR9d�) i�(�!�Č  %\���	��W�ֽB1nU�L�!����r��9�M�>����w�U�!�O2}��p�Wi����Q;�D
z!�ĉ&"�ASPiRv�����կ<\!�dC�X� ��Qa46��ӓd��kD!�dEN���W+K9"��]*�$�+i'!�&r�]a�I�~hEZG!\<j	!� D��D��>�	���� eY!�dQ�5/�њ���"l�x�cW4bZ!�$X"��s��S�t���(=!��
�cr��0��O�O@�E�>-!�/]�t r��B�"0 ��џ*!�D3k|�1�ª�&1)��+�� �!�Dɷ����,=
Q�Q�G�!�$ߴa���Z��/
V���
��\�!�$ͣ<d<���U+u&h����\�RB!�<�̥��!T�=rt��(5!�� ��t��W>�����8M��I"O�\��S�$��D���
�g����4"ODqh[Y�]�M��Wm�����x�<)%��J�xYd9NZ���$�q�<aF�� "YelN�dr�����k�<1Սފ;��]�#�#4:���@D�r�<�HF"0���z��]�8Ma�i�<�q��V�p�k��k��ģV(�b�<�%B�PÖ�C�^1��V�<)W �4?zS *�<9�5k�O�<I��^��cvc �.LT�
  �P�<�թM����L�R�z=z�!�H�<�5M�(6�D�to�T���E��j�<�t-J�=:���R�B�!��m�<vgߞ���hU�h3j�ks�DA�<94'�����
}6-XH�s�<�m?'ި �S�Յq ���i[m�<��

I0�oO,:1ޑ�g�~�<����4=�d����Ϧ2���$��x�<��!    ��   �  G  �  �  v*  �5  �A  M  �X  �c  ^o  �z  !�  R�  ��  ��  b�  ��   �  H�  ��  ��  F�  ��  %�  ~�  ��  ��  ��   �  c �  � � �! * p4 �: �B �L kS �Y �_ �e  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&��Q���I�8bE!�۽}�6����>:�!��P�K�`U�1� !�,Q�~�ўx��)� h����M�+����&�R�z����p"OH��e��%�>q��/�*S�����A(4� A�'��ޙ����3J�Z�H!�OR�O,j��I���a�)� �|-�"O�Y�C��"Њ�ÇC�@�"OHh��ϟ�P�Yɧ![�T�T1BO��D/ex�5�qL����eoĶ+!�ʻvBPa!@��P��NF0�!�d��?T�5@�Ή���\�D�Ӄ8!�Ğ?ZJx�mN�`+8<9�	�,K�!��\�'d��Ǎȼ&���r�I=�!�dR	�n��*�-Of�����L�y!���H����%�� !,�D{S�QMY!�$
-t����&H gl,�rao۩N�!�D_� <�9*��j��0��ÃO�'�a|���10�Q���§'R�A �Ԩ��?!�'�J�r�/E�3�v�(b�Ȏ,�����D�~�O t���B�nm�Q� �UY<��'_(���.V�d�<���?0a��O�O>\F��O4�a�7V�`�v�S=6˂��"O���3k��d\$��ѤM�wY|DR�i�����Z�H-pu&֌3�2�8�B�%JUa{��C�jj �X�`˩2�`�����G#!�Ĉ��,d3a� �+�2xЯ;7!�d
�)i�4�q�	)����'��B�!�@+.Q�!o��Q��9��n�0tf�IB�����2 �I5/��x�Wi�U�F�:�"O��f	�)��)cQiMV�Nur"Op��#�Y���,��H,)�|��1"O�x�7�V�a�&���HB���"O�m���E�d� ��#DHj�"O�e�Q��m�\Բ�G�_�Q�A"O�5���G.m�
\ ��?c.m�"OQ�胱Y���	`H�/�V �P"O(M�Z�*BX���/��tc�"O�J�D(�lA0�%A!���"O $�2I
7b��ˁ$�
�R �$"O�`G��$��b�O�^5��"OΔ��%Ŗ6����GB�-�	�'ӂ�p2ɜ�#�*`�ąz�p�*�'�!�%oEgH�����9KZ���'TԊQk�$H{�A��ăs2DaK	�'yR	K&�Ҧ�!g'^�q\��*	�'�.��w+��	��5�'Ă�b>�K�'�b���(ŐD�m�E�^�T�H��'��u b�I)�~` �KZ�,���'�V��"i��+��CO� `�'�`)!!F9c'li�'�DYb@��'4��c �K?Qy!���K�̖p�<�ԄS�N;n�hE
u�Z�!@�]b�<Y6*� TT)�vb��@2�PV�<Q�j/\��6N�v�6�{$��U�<٠!"�H��2bH]f� 5�PS�<yA�d�)Ӣ�ק^��ٓ�χj�<٠����v�ɕ+��l4r����b�<���S����5 �;{�Ҕ{4�	U�<Y�l/��st��Nr(�p�G�<�R-ص;Π���G�캤��F�<���K�Hi�)�\+�z�jDY�<16L٣��\"���, &p�qL�m�<�"n3v��)��k�r���"LN�<�#aKM�H�'kɏ9]
��g@�U�<�#�U�Wi���(���� [�<�� 
���)�9�ȠA��Y�<� ��jrF�,JOX�)�4=Tf��"O�=;���>�1��ZAn�z�"OШ��Qt�A�r�_�'\TI��"O��ɇ!��R��T�$]��c���yba�)v�Nɡ�C��.����6����?Y���?����?A����O����O��B���>�ɒ��S�
[��B�C�OV��O���O���O��d�O���OJaC��ƹGBD p�f ���U�OF���O����O ���O���O����Oh80��3dZ�A����O��(�d��O����O��D�OF���O��d�O����O����SZ@�>t�y����O�$�Ol�$�O����O��d�O���O�f��g����n��T'�l���Or�d�O��d�O����O0�$�O ���O� b�ٗ���W�$#U���OJ��O��$�O���Ov��O��D�O��O�Z�6-�A���&8�f��O����O����O"��O���O2���O��
T`�$;�&�t�
򺵲%��O����O\���O��$�O����O����Ota��c��5.\h��.��R9q*�O>���O��d�O��$�O���OX�$�O�e�¦�?����,�8�pl�Ѥ�O����O����O����O����Od���O��A�
��@)"\�#��$'V�T�7�O����O��D�O��D�O�d�O��D�O�L�H�1���X��Y�t z�B�O���OH���O:��O���Ǧ�������F���icFパ	��]�ả���O$�S�g~��cӘ�w���j�IW�4t��#D��%P�����Mˎ��yB�'>0E�t!U8K�� �Ï�,Z��k��'2�9����8�'9����~"ҡ�9l�0�0I���,��$R}��?�)O��}j��SZ����v�U�<v�"�H��2�ƥ�٘'�	nz��)ܭ���KW�E�_�T�K�(������<�O1��xӆ�ɀy{ڴh���O�4Љ�	��>��I�<��'��,F{�O2.^?Q+�\)&�ɟz�&+a��"�y�R�x&�`�4=]R��<��ܹ�2����:��������'�b듵?����y2[����
f����/�J3:�S �=?��ȕ˦`Zs�'���DZ3�?��+P;�`Q�$xb��r����<��S��yb!ʐ� 8#E�
&OC�\B���y��i��q���`��4����ԣV�q]pltϊ@��I�PL]7�y��'�r�'����i����|J��O�Ɓ#aU�*E8x{�G�m���Xx�Ily�O��'�"�'���N�2��ЈJ����I��	�M�@"�?�?a���?yH~r���"Iy�͛�D�L� � Q�s�L
�Y����4@
�x������rm���]��9j���q��D�S-�#D��P���W��O6�hH<�_�`�Ѣ�-�ʉ�6(@�>a�`Z��쟜����$�I��Sfyrff�j-��6O�P�q��D�x���ȹ�)��6O umN�GS�	8�M���i^*6����Y���JȂl�&��  �M��'�X!Y�.ۑ^X����_��'�u����vM1f'��0���&	������;O��D�O����O���O��?%r� Ůu6^�)�L��ԉ�'�v���Iޟ���4-'d��'~�6�,��Ջ5/nu;bC@�Bs��Ps����N�$���ٴf���O
J�)#�iQ�ɪ?\��c��9~�B�#�"c2�`�!�S38n.|�sy�O�'�r#T�J� ���&ɻ[��D3�ӊA��'&�I��M���<��?Q)��x:WJ@�9S���WЮxBF��P�����O��oZ'�MK��xʟ��A�ԚvA��PnͿB4z���*�N��P���)��i>E�r�'��%�h��f�'�6�@��-#�۱�T۟`�iYn���)�ayBgg�$�f�ɽ�xUp�#�Z,}�I �PG��?�M���>�i]^Ѓi@�����Å�+��aԣe�4	lZ22t�mZ]~�I@��8�S^��I)�F�Y� �Z(��C6*F�i"��<����?Y��?���?�+�P[�n��#�QSa��H������-�v� ?i����O��7=��  ��;�ҥ��bA����������z�4q艧�O�S��i#�d4] �!ۡi�?�dh;@�L�y��d�7��8��$ȒO���|����)j��ѾNf��#�
�$\���?a���?i(O�Pog�I��|�ɅR����3$:��Ҳ�B�@�T�?y�X����4FK��++�
� ���	ڼ4ʃ�7s�ɚ3
�hrh?o5�P$?iH��',�T�I=$���]�6�@ԃv�II����ߟ��	��X�	{�O�rb�'p@d�
����pC�� f+��m��� �Oz�$E���?�;������Ւ���t�#�@�����%|�(�l��H�m�E~2���F�����Hx�1)Q�Ej��
�-<XX��|�Z� �	���I����p���{_��+��ю�Ҙ��!]myBmy��	Z�F�Od�D�O�b��
�__�$�#d�	�v�QT��=��H�'��'O1��9���T;T�� �āS6�ླྀ�*\�=��7-�@y"��V���������5&�ٚ�'?Y�Ή���I3t�R���O��D�O��4���nl�ƨ֬y8"�>e�����H�Ң=1�k�x�Bjz� 㟨�O$Uo��?�4:b`�Ac�ΑwH!P&A�{��X[���M+�O��2eM�s�4����� ��s�M*g�R�`�HJAO�d��;O����O��d�O���O>�?���Ɗ�}�t�0DN<@�x�%��L��ϟhs�4F�r9̧�?с�i��'�d��ӊfmp0�-�*^�.r�'�:6�ʟ�i��c�J6�<?�'�J�ɸL�0��á#D�7��=Q4@�O�HI>Y,OP���O����O�ep�5��2��ֱh/�h��O���<)B�iP�Tsa�'���'n�SG߮��W+�'X
rY3���9�\�H���=�M���'����	� d�>l�D˔�i��a:��Sf����U�1�޹9�l�<ͧX���d�2��bURp9��~��2�c��F%����?A���?�S�'��d�Ʀ�+��P�7�Uy"��{Vv` �@�.Q
���՟���4��'m��
Y����$I�(ub��Q�h��MZ�cU3y����r�t����x��[��0������+OvqVg[J�(B ,Y�'zi0O���?I��?q���?����׊mL�Y����lÐ�b�@��-&�m��PT����D��m�S�P����#���/'~��C�ǭ�԰�WeR�����O�O�I�@�I2#�`7�h�,�w㈭#���xЧ�č2��l��:��Y�$W�J�z�	Iy��'~R�̗8\0qPAň*��Y!ek�3��'W��'��iu7m]<T8���O8���5��=�IF�t8n1��E�Jaz⟈x�O�1n��?J<�G��'Ŭ�6��#2� ��EY~m^��I�DZ�"O~B6��OZ����T�K� �5X`d�r��\��=?J��O���O��*ڧ�?�EP�` s`Ӣ!"B�Idi]��?��i<� St�'���o�4��6ot�˗L˾!B��x�hʹ
����M��'l��@�7������`�gJ�	�[��n�"˅���䊚�xh`&�ȕ'�r�'W�'n��'Ҋ��� �q�>�C%�;bgt<�#Y�<��4nfj��?)���O�E!��Ӗ\ܠ�7�[�,�s�.�>᥶ic���"��Iͥ�X����$��lBD�CE��A�1@?{���-��gM�Oĩ�H>/O����.�v����Y0r��䋴��O����O����O��<���i�)S��'�(�D�jzl%���2VA�ɸ��'I�7�/������Ħ���M�τ����ra�Sb�m�ǯT�4�rĐ�4����*����'f� ����Nʝ~�DbV�xM `օ��i��D�O���O,���O���1��2?(��  �+<�{�'U|p�9��Ο�����M+h�|��U#���|b�(:2�"�"G@����D[^v֓O����O���z�&���A"Jm��m�uG�0�\���̡t�R!�&�'c�e&�,�'�B�'���'`N�r$�
5I����#�DW�n����'!�X�,��40x�=��?����i
RvU�B}rq��h˳�����dS�-P�4X����ɑ�{���x�i�<u��q��F˭5g�K���+w��擴,���r�tBE��[',mLhǊl����I����ן��)�SFyl������	�m�$wn�d�1D�7+�ʓ@�f��B}"ml��]���,�V��U`|��q���i�ڴM&����4��ăQ� ��'W`�ʓ�b�k��Q+s�]��k+��̓���O����O���O��Ĥ|�⅐�-�x
0D��?�Q"Q�ہ>���F�B�	ʟh%?�����M�;��
P�W�zؠD��]�`=1���?���x��4�D�3I��6O Y�2�G�|�,�2M�s�"��b3O|�	ç
��~��|bU�d�����b��=Z
�ږ��1L8����䟜����p�	Oy��f�v�t5O|�D�O�Pi���'J�aR�ě�;��h/�I#�������ܴj�'�4�5Ā�/Τ��yݠ�O:��ŕ�|Z8�a�	б�?�am�O\[�,]'��:��h(��Ќ�O��D�O����O"�}Z��|�5�@D�hւ\8�,�4I�������&A�������?ͻ"�n�l�~a(V*�G�H��蛆�zӜ�n�K촩n�i~��T�-�v���B���������k�/&J :e�|�[���H�	��d�	�4�0�	����C�Y�l�{�#�Cye�"��w3O�d�O����p0R�oY�
Ja�o��'k�6�@榭KJ<�|ZCD��}�6�8'D7+t��#@(��E:� j��BE~2�P��v��Ɇ
��'��xK�Ѥ�nQ��!�'M!
���H�	�|�i>	�'�27��(�&n����
 t��Uk�M����Φ��?1CS����4Aڛ6.s� e�V/C�d�8܉k@2C�q#�GL�s��6Mt���	.n0���O� ��"��g�8T��bZv�L)�S��A��e��?����?���?Y����O1P�c��lz�z�d�'�'��'��7-��R���O�(nZd�ɘt�qq+�>ʴ*���.�j�QO<id�i2�6=�@��Reeӎ�2�$���<L(���Y�@:�c�f@(EP��A�����D�O��D�O��D�2Ɛ1j㇟\�J�@ퟁci����Ox˓hH�FP�c���',�_>���H_�<,�4�v/��d9d=�F�-?�]����4e���j/�?��S+�=_J�jC���+I�x�b�V�>�0L����6������L�P�3�|�͖ ij��Y�Y?2��mQ�&[���'�R�'���4[���ߴ5h@
��.ZȜ��B��TƆ\�C�M���ċ¦��?�BP�D�޴KFN�:�U�v�x0��.��o���s�i�D6���j9r7"?'b�y�t������� ̔f�T�ۨ���$�"[��jA0OF��?����?����?����iڟ}rPaX$E�&	4>�㵀�T���l(XǦ�'0�����'2�6=�
4����x�-�3I�9}Y��+�@��n�1��S�nX(PnZ�<�4ѠC`��цS
jS�����<��i �Ȏ�䓓��Ot��V.�N	0c���5c#bG=�����O����O��TL�F���'�B�[�8�`����p�q`'I�C�O��'�h6B̟�&�
���
�0�	��C[Z�9tL7?��χ1���uh&��7�����?�'*W?F�����I-��C���?a��?���?ю���O$L�&��5f�\R�C�-�(�rf�O�o��:Ӛi�':6M1�iޑ���w�h���MW�I��X:Qf� r�4^��&)r�|0��%o���J�(Adb�|\C�IX�mI(�Z4	E�NW��X�������D�O��D�O`�D�O����G��q��k�b F�2�#ۊ,@<˓��6�/���'����'V\��bM��R����I��H�;��>���i��6͚i�i>���?!��D%_�E1� ��>�tP#�76uT�Q���Fy2�#����ɗ~P�'��!}�0��P��nX��ۄ�͓u=����ޟP�I��i>}�'�7�L2A��Qb�� 	�䔨N;0��%�ߑI�D�Ӧ��?�T�`3۴^E���oӴ AĬ�hn��i��ʍY�B��#�6�)?15@$"A������'���g�Y~��� &K)t�L�gk��<���?����?����?����ۼk�dmp���U���@c�	]B�'��C`Ө�� �<�g�i=�'�x[d���
�ݒt
C�v�6`�!�d�O07=� �(â~�`�Ud)� H(=k"���`Ɔ-�r���M
���������D�O6���O���D�<-PF+v 9	�MY%;�����6�<!��i�P���'1��'���"C�p�Z��4a]��֤ד~�o��ɳ�M[ �i��O�',RVp �-�S�
���K�	!�p�¢DE�n�:E�Hy�O���I�Sc�'q�͂��C�����������'���'���O����MK�� 1�>��'�:�ҽP�G�Lxv
���?���iN�O�X�'�6�U$nM1D�/�.�(b��;=\Tn�!�M��H��M��O A���.��b�<�r�G�rH�	��$2M�<	/O��D�O���O���OB�'q��a��,��(yE-�^��@a��i�,����'��'��d�nz��!���5���J�3'����M��iK�O1��A�tӜ�Di��T�%!*2�u��Zy��	�H-b<2b�'n�I%�$�'Sb�'Bn2�D�t;\��N�h��#��'e�'R2Y�,��4|�����?��9)����ĩ8"@8�G�8}�5ۋ�c�>����?	ӗx�!��w�h��2��2/d��!�Q���$
1!dN��~ӂE%?��5�O0�d�A
�ݙ�kI
jE���S�X���O���O^�$9�'�?�r(U��^�	��Ta���� �?���i�d�!�'%q�>��)q����U(l �\��
7$�	ɟp�Ƀ�M�&	���Mۛ'a�)
)1�����a�KW���8�[/>��K>	-O���O>���O���O �j�_�H(�!�"��D��+�N�<�g�i~6���'�B�'���y����&��'��f�芐f�o�4��?���5
���O�ui�K��r��_ LQ IĻT��F+�<� ႂF!��	@��by"�T55@6�q�˾[LR�j��עO�r�'���'*�OR�I��M�f��'�?�H�C�ҠI�HK�3d��L?�?)Կi��O��'���'�R6�[��x� k��L�����I�{��𫕄c�$�&�f�+&F�?m&?i�0b��!P�Hb��p@G\�Y�	ܟ$�	��t�I����	L�'aBr5�6=��Y�ʀ5N�FD2���?��F��%�����'t�7�0�$�:E������)@��8�kv�'���ʟ��g��l�X~�k��n�豓W�^�-�v�@���]��"�^z?1M>�.ON�d�O����O:�R!������&�960��Iܟ�'�D6D]Q�ʓ�?i/�
T�*��}j
dhaV�}2�ĸ��,��O����O$��#��PࢂO�S���!bR��*2��07��r޴�i>���O��O��S/S
a�HdO�L�P���OF���O`�$�O1��lΛ&hU]�l��!aTv8�:"BݢB���u�'�Co�B�̠�ODAo���Δ�wEG6���H)H�$h`��M��I�)�M3�OF�;��
�jA��<��`����`�̛G|�87���<�(O���O:���Od���O�˧,TBt�e^y,�;��R�Pz�=���it��'���'Q��y�n��NݞSo
���4c�U�ťW�mZ��M+�x���B�;G��3Of����ʣK�  Y"mP����?O�<6oG��?ّ!���<�'�?!'�\g���ft��A{�"M;�?)���?���d�����R���@�	��0� ����C`
�j�ph5��c����	��8�I��ēe�>u�&�άK:tAZ��޷KwE�'�t��\�1ط�is����I�'�2J)r�"�̓&?��҃����'���'v���D� ��:+�����VG�}�G�t�ٴ�x���?��i�O�.F�@�޴p��=`>��q�K�70����OX��ۦ�צ-�'Gب�5�[Y� �7f�0��Г��x��-
�1�D�<I���?���?����?��c��CJ�́�c�+L��
e-^���_ܦ��T韌���`'?�ɼ��9�Ŗ)� U�T�ݜ!��۩O����O�$�b>=x�$�YY�H[�aJ�]�*����"j��n���'<.]��'��'����(yu�'�U
0A�����Ɵ��	����i>�'��6��KI��D]^�Π!�C�)A2�A�F& /`����٦��?Y�V��I����ڴfD�R����A��Ũf��+!+��h�(K��M#�O����BB������w�^�@-͟Y�p%��4I)�hx�'�b�'FB�'���'��6=J�`��e��#U�H�y��ЂD��O��d�Oڼo��m�'ђ7--�H�Đ���Սh-�� ؑ[ T$�`�	���"��}o�C~�� 5bȪ	�g!�i~>d!Ҁ�J0f�3W��Q?�I>�.Ol�D�ON���O,�d�M!{�x�HѬ�.k�p�����O����<��iE�E;�'���'2�cgZ1Q�$���f�5$�r;�$����M�S�iDRO��m��lrC��y`BA52���ж�
�w@Py�O&��I�'�b|b@A�O8ij�ǀ O=�����'�'X��OK�I��M��ɕ;s�,Z����CUH!�w�b4Ľ����?)��i��OU�'�`6-��)�c	 v�rѡ�Ɛ6l?�Qoڠ�M��陬�MK�O%Ss��j�Ƹ<!��ԵG�B�K�&�b�h1����<Y,O���O����O~�D�O��'zS� ��U8RR++Ѩt�P%���M���?����?�O~���	��w��ԈA!�G�� �c?(ԨM��)�OZ6�\�)��� mN7�~�h�7�4
��͓�k�����Ӣ�x�\��[:[���l�I{y"�'t�J�z��g獤'��؈B�ȶ_��'c��'4���M[t̛�?����?YU�����;��ʏ87\�S���'P����vDk���$��zt����9zd��f+���I�G�H����!"7��'?��t�'.���ɐcN$�sĔD5&�	�e��HǎE��ڟ �	П��IX�OAr���8�H��p�@'�T�X��`�b���<ɤ�i4�O�.	�(�6�pm̶W8V}�u�6iI�d�̦��޴T��(�<.<������p�\�l��D%���=���0-�z���䛛@D.5%���'L��'���'L��'p��U$9�<�b�i������Ty"Mo��aqC��O����O����<z�R�r3`�5�,t�-D�9n���';�6�Ǧ��I<�|B�Ŭ6�B}�Q���O�vr4�Բ^��٠�T��DѤ�Lͪ��P=b�OF˓G@j��D�ݟyqʨ	D#J�M�F����?����?���|z,Oz�m*��5�IDȠ��Si�j|�	��>q���I*�M��rJ�>��i��7m���CQ���,�̝���ּsdvv�Kh0Z�lq~BDX�/�V���;s��O�'(� �܅q�*XB$|�/��y��'�2�'�b�'���i�V8��)4i
��aŜ?lO���O������	��)?1��i��'gl���]�P�Y�MΜOJ�$���6��O�6=�Y�W�r��0�T	㱇�[jf(
4�jp2TiG!
z���"�䓈�4��d�OX��KJy���#h�?x`�$H���90[��$�O�˓u���.\;<���'j\>e`gI��f�P#͜f� ����*?�AV���ܴ,��� �?�[���/��І �+2S�=F	J�5'<�In�m�����G��� �|"�ڄQ4T����
	)A>�Ҷ�W�!���'BB�'����W�p��4_쨚4 ����cpCA�����vO�*�?q�9�F��M}�e~�4qA&��5S+T.g�*�å慠.�6��香x�$_��i�'�N͑B�G�?�åR��d��
��N�3&q���j�ؖ'yr�'8��'�"�'��S�N�$Y��_BdE0�L�/�,��4yc��S��?���䧪?�2��y׉��.6�,����/Bi Q�r��>s�6�צ�(K<�|�uh��M#�'7<0�j�5$R�!2S���-?��Z�'��9K������|�T����ßX�K�/F�çI�1��M��ڟ�I� ��Zy�JjӢ%��d�O����O6�����"TD���Ej��� #��#����	�4�'��y+d�L`�QI6ϋ�R8���O�$c���+����;����?)��O�[�NM�S@�P� �<v�!s�h�O����Ol��Oޢ}����٫��RG���C��zX�AH�����C��R�'+�7m?�i�eQw�`�ưҤ��9��������46���.d�@�'�dӴ�t!�7���\�C��ʲ!��0�wg��	B�tq�����䓋��O�d�O����O�N�l{X��Q(0�r��rE����P��+Y2�'���)-Pz��Ц�/U���iG'�%Ni�'�v7��ۦ��L<�|b�jLk�b�I�1x����2򰱃� C!��d�w�hأ�� �Z�Od�	�	�#�f�(�*�:_�����?���?��|z)OĐoڬ]��a�I�g�	�Vo)��Xy#��HӘy�	��M���$�>���?��i%�H	@��:���Y�[/A&lL��"�6k�f����q�;W��=�i��(�p�*!�R�0&�"l�;B:O��d�Of���Ot���O*�?���m&@]��c��x��k�d����Ɵ|�ݴ~f`�ϧ�?�лiX�'��!��X�,� ��&�%cNm#�>���O��4��	��uӼ�O��� �p`��\���x��M��!�6=��ȇ�~"�|bT��	ğ��	۟X8�G�����C|��9���ʟH��gy�&}�F13�˺<����iK�F5y�+���|�nT�%���#��d�O��$S�)
懇�~�8�0�(�S$���،a~�8;�߀�Ms�^��i���4��� Nf�`b�G�{{��Pg�N):G����O,��O���)�<��i4~�s�E*z�⎇<*�[��R�WYr�'�d6�%��8����O��M���|�i���P�N-�7��O0<nZ�^�޸n�s~��QF'� ����č"cxr��(ԣx6H�Ѧ��(#|�d�<)��?���?���?q/���;ь�5@̂�3��^>G2�d82��񹑭�Py��'z��\lz�)"ժ^�[��(�և	6 Cq����?�ݴ�ɧ�'@�J��4�y�)��4&8�)�
!L�x�P/Z7�y� B�����	��'����H�I [>��PaܯZ�D$�'@�40d��	ȟ �	🴗'�6�k#����Od�D�4Bf��ǅ_� ���"%� 	���a(O���}���&�� rHީ+���{��G�0�2�!8?q�f�`��0!ajø��'m�����8�?AD'�(%2�Т䞵)����BY6�?Q��?���?A����O�]�'ߡH�������v8B���O�%o�d͒y�'�26�:�i�;@!�=T1���7(Ҡ������s�XJ�4.���e�h]�PihӶ�B-ht�g���"�#m��D\X�a_Na�J5�S����$�O��d�O��$�O��DܯJb 
�g������=�J˓v�vbW(_�"�'"���'������Tou���V�6Z�2�%ad�I�M+ði�6O1��Q���Y$s�J�J�^�p��k�1:j�D�·<����.0������䓲�D>��,�d.W����j��H�gA���O���O��4�Hʓ����- (�*Tq�Ep�eʯO|<��䬅�y2�}Ӵ��	�O�|n�;�MC5�i�Ve��)�MX�U��/=�t8(�%҉�����A��"T���j�D�S��a&��O/ʑ Iֆ"�H����i�8�	ڟl�	۟`��П���A���WF�hQ�E,w&a��-��?Y���?I��iФ�ZbS��X�4��Z��!C�f7pq�xi�`	,H���x"r�� l��?ѹ�ڦ�Γ�?����d�5ˣ`B�Kr���s��KO�x����O,�N>�.O����ON�d�O�`��'�f��a���Hw��iǪ�O��Ļ<��i�ޠ��'���'T��� ���67�I�@8�l�6b�I��M#��'C�����O$��A�]8V>H���ʲp.|�0��ߜ�&t�u�G���?=���'Dt8$��#A�6_Vp�0��
��H@Ē㟜��ϟ���˟b>�'�\6�Y�C,*�S`@X95d��%Q�b�����<yp�i��Od�'��6��k(Q�@��"q�6�Q�x>}m1�M#`֭�M��'�"�8 �!���)��ɻ|��lR�G��I�(h)Q��
)���	fy��'2�'�"�'|bQ>�ka��K�$���,=V����f�F��Mcug��<���?yO~Γ^ћ�w�Va���H�� 0fh(�,�bu�4�m����S�'[�^�h�4�y���4p��B��*	 `�%���y2�-(����I#^��'��i>	���7�d�V�E�6����e��VL����h�	՟�'�7�T��$�Oh�d����+�C��@K�90�R��C/O��dc���%���PB�)�=�h�,}i��b<?Aĥ�0jT�h�IDp�'}U���E0�?1 ^�A���9$�N�4�|��̐��?���?���?َ���OP����m�Z����ˈ	�p0C!)�OV�lZ2Thv�S��&�4�@Ei� ��5r�%�3[{�Q�79ORAlZ�M��i����ղi.�Ig���R�OB�EKo�t�w����L�q��q�Qy�O��'r�'��A�L񐸲a��/ORu����c��i�mڻ�t������IP�s���3lۨ(��9s��6_�,�Ê\��������ݴDp���O�����,�K�R<B��X��
�bN|F��eY��SD#8bB�Vw�ILy��Q7+:6A���3I����ښEQb�'mb�'��Od�	��M��E�"�?! �C��F, 2�\5Q�A��<!��i��O��'D�7M�Ʀ��4'�XcO�#��Px�4����aeT�B@�N~��ҷ7P����OKw��-S��!����#�h	[�Ð/�yR�'�B�'d"�'���)�3��Bk��R��a9��P-��$�O^�d�Ŧ����E~y�
zӤ�O�\"e��P�f�jan�"�X��@Ne�ɼ�McZ��ɜ>�F7�8?�sɇ�J�$�r��	�~ESf��2DSR���O�`�J>)(O��D�O<���O� f� J�T��QIV�:�b˔��O��$�<�Ըi>�:��'<��'��S^?�53A��M2 �Z�EI�$�C��	��Mkһi�HO�S�Ƽ�:D�	?9���y�
]�}�$9�ŋwh<���k�My�Oqڽ�I�m|�'��ٙ����H��I�ML�mܺX��'��'�����O���%�M;$�!���Ƌ0o�.E#C��#��(O��o�X�i���1�M�DJ�� @�|��S!vi�T�#����6Dh�u3v�o�n�#B�}y����T�)O�DYsi4!2��K�d�is�@��?O���?����?9��?9���)��?�����9- �ʃ�G[�^m�1
O��������@�s�̸���#pJ\�/�	Z���=2�b4Q�@�2R�����O0O1����z���)� ���%H�z����"14Ҽ��;O�q)�\��?�C$�$�<	���?�,�}��QT��<����#��?���?������̦��`L^Dy��'CDD��`I�´$ؓ�� j�kC���N}�i�Dd�	Y�ɲR-��
��+O��� ��=��T���#��&a{��L~��l�O��Q�5~6D@t��D�����GϢ0x���?��?Y���h���D@�}xh��CI�%�8��@S�9�$�ަ�y$��Gy��i�4��}�
�A��"�.�qMY�5����:OD�mڝ�MK��i,¹�W�i<���W�����O�<�K2�˝I>���P�Y�\ �uxT"�h�	dy2�'S2�'���'��+Y)*ah�`�g�_�&PA����=��ɔ�M�B�A2�?���?�K~���m��s!�B��8��cF8{8>��6^��!�4{:��x�����	T��4pE_� ��%) �Xa	a��J&�	b�e(D�'�D%�`�'����r�ޟb%���G��:Q��B�'�"�'!����4Z�<��4�0X)����$;���s���0N��t!���1���B}2|�҈�	��覂�Fm4�� 	�F��P��}oN~�"C�&���S��O:g%��	�j����'`��|��,\��y��'��'���'����!�8�A�%N����TfK˓�?���iKL9�ȟ<in�]�8U�ΜaA�B�@o~��dF�cc �CM<Y$�i��7�����2w&}�:�����S�ό�)��cPb��d@bB/U��ȓ��' f�'���'�r�'nb�'4��s���D���TN)X�a�7�'�2X���ݴ������?a����	�_��9��n�4P���) ?~��I��$\���*ڴp̉���^
�j q���/�����&̼.������L���z H�<�'=:�D���r�f��&�XІ�6��ir@����?���?A�S�'��dY즥A���@ D� ��-��8e�QeS>)�'S�6�!�I��������FF)^f���B�O���ѭ���M3�i�:�Д�i��I(_cd諷�O��)�'�l�� ���ݐD&.��m6�a�'����� �	��I�T��]��� -���s�)�"�z��f.Ԗ6�	U�:�d�O���?�9O��lz��r��r�k��@&�>`Y"X5�M[ �'���Og�s0�i�󤞬	�FmR�&�#e��`�����&k�%���R�O���?�-�4m"�h�}z�k�kB�g������?���?�*O>	oڌ7f����ן@��0U�8����U�-h�Y,�N �?��Q�$�޴W��x��02X 1���Y��f�����)l��6F���
$?A��'�
(�� b3�<c�!HPm�R��;�0�����������p�O�"+-`���L�HԪ�Q����i�X0c���<���iN�O��֫��r�H�xtM��J&������M;2g��MS�OxA!�f�'�ꁨ ]5֨J��`p�(�1/��Or˓�?���?y��?��hF��15�T-}B� ��탣-e�1X/O�1lڒQD}�I�����|���|z�DI�~�hTK�(��%����$W�q���S�''�^H��n���*����j�XEo²K�@I�,O�P����?�%�;���<��EچU]PJQ���ł��HW,�?����?A��?�'�����Y��՟PXG�53LB���*WXq0!��şDC۴��'���yW�ƫ�O�7�ԼKEi��Ϲ�U³
gI�#Db���(|$�U/㟲=�I~
�;��k�$��;�
�S��E3(�|���?����?����?���Og�� ����R\cv�B�aP�	�Q�'	��'��6�=5��'���|r�Y<�x���=X�
%�v�W'`��O�n�!�M�'�����4��d�]xꠠq�O2m)����$̚A!͊�?��g8�d�<���?a��?yB��,@p|+�GK�}b)�3*��?	����J��ɪ�b�П������OˌSaJ#	�0Y ���6lR��O|Y�'27m�Ѧ�BK<�OD�z �W<k���t�lԊWA4ɞ��b��7C�i>UsB�'�� $���%�G�"d���`J��9��N�����؟��	֟b>�'��7�Hi b��?hCؤy��-`�}[�a�<Ys�i��Oʤ�'I�7��4�e�«w᲌_3 � hPć���9��4a���ڴ��$��F90��"��ʓj��������m�&&�Z ���d�O6���O^�d�O�ĭ|��O�V��j6JWgD���r��>z�����R���'P����'W�7=��R���9	u$���C�9�╻��J�}(ߴH#���O��x�'�i�󄖖R=��u!�5��:���'&?��0i�]p�Qhn�O���?�X�1�G���(	����L��b����?���?	(O�o�+t��Y����h�	!2�Z�n�
�u�a�[��^��?pR��H�4<���&��˺=t��3���8�PPl��a���
Q΍* ��3=��Q$?�"`�'��}��B�,��Ԡ�NX����0Yl��	���������\�Omr��L��R�i[�!����!\4�"e��ݡ"�O4�$�Ҧ��?�;@,h1!s��U"�H7eJk&D��?Q��uR��`�%�斟���O#4�醝�A* dɋB�<��� ���Oʓ�?��?a���?��P�2�۱F�+�6Aq���($z�/O��o��VF1������	W�S���i��hRv���F�Q�Iن�"���Ԧ%9���S�'? .� tչ�M5YM��1ĘW4InO�Ak@�c�]���O.�IK>�(O|	@E],~��q�F��sNpda�OP���O�d�O�	�<Ie�iG�'��\����a:��� �gh=#�'� 6M,��(��$��Q��4l`���%Po ���-J���"�EPi1� ���i���A�u���O�q���Λ�M��<zׅ����	¤�%>����OZ���O����O~��=��0S�Huj ��A�z��B̔aF��	���I��M����V~҃qӚ�Ol�s��[�y@ G���-떤�z�I.�M�����t�,F�f���P�IM!X��x`��F0L;>�Q�ކa�����'�l '�������'�'4�.l���v���@�BtiG��-R�'>剞�Mk�E�e~"�'P�g$��h�2o_ 	����(f2�c��� �Müi3�O�S��=2`}h�m�{���1Ɯ�2%��tFl��O�	+�?��M/��@�J�~�H�M� OĆ8`�$Y�����O��$�O���ɣ<Aq�i�<��R6��1%n��|�6Ty�"H���\ɦu�?Y�R�m�)�`�0��E]�Iwc�Y)�}�ڴI��*H�.��P�p�_6EU���~*@�ʳk��x�Ck�3w'Ɖ��f��<�.O����Od�$�O��D�O�ʧEO~a�!A��ZXd�@�ܣ�X(�i*��:�'��'���y��p��Ε�Q����.7��,��� <C�qo���M���x��E� N��v<O�Ż��C�sH"�y��֯'�����=O2�����?
.���<�'�?�A��\P���A�RB$9�K���?����?���D�Ǧ]��c���	��dJ���RؤI�c偏;�
�Cm�g�~o�	 �M�g�i5�O\A�alC�~!�Ya0�&X�@1������E^@�41`�m �ӝ@�Rm���#�iьh*����ܜ> -QeŞ���I���۟,G���'\�a�����g�,|s��7L%đ#W�'Ґ6�K�Wo����M���w�	�RCڦw�P��O�K��Ai�'���i�V7M� �b7/?��Jȥ\������01@q	�.�EM, Ag��;c*��K>a/O���O��d�O
���Oʍ��`�p^� ;��Q+g%�<	$�i�����'�r�'��O�oE�F�R��e;oLd��F�'�J����dӄ�$�b>�#dhRu#.	Pv�ۓ;����dHV=o�� R���Py����Y�M�ɈZ�'�剃ܚt+QW�nY���8��Y�	�p����i>	�'��7m]�z��d������L�����Q�8�D�Ϧ��?�S�,��4t��Aq�����^�PĤN�X}�]*COP�Je�6�/?yw�=u�b�i������a��,j$���ˎ�`��d�<�
�qV�ԡ5nեG�P���-��/O���m���=
԰i�'������7l4P)eG5%&����)*��Φq��|����M;�O6My#(�8sʄh�q(J�N,�v!]#!����4�O�˓��'��P��-M'�]�& U)^�9���9��my��'R�Ӡ5�lbௐ�ND�!#0	]&o���$��I��M �i�O�ӂS�
��S�ܩ�#J��(=8E�	Yd�"��hy�O<~x��f��'Ŏ(�ڈ^j�Hw�	c��!��'�6-�&N.eS�lM(�N0��JKd�2q��d�O�����Y�?Y�\���ɚI��= #�� ;j�!3$�#�.-�I��M���K��M�O�1GGS���d\���i�6���x��0��q���'a�{r�OB�X�D��W���q��0DL6푪,j�ʓ�?ى��y���W��2�-/x"�P���Zu��mZ��M[�x��0|�v5O��T���%$Bi��\�|�l��6OR(�F"W��?���/��<�+O$��&��({(����*�$�a�'X�7�^�>�d�O<�$<�V�sR�	�P4�)��GZ�	�J�p[�O����O�-'�, ���>wǦ� v�B6��Ё�F3?�Al~���P�i��������'
B�C���4�sbN���J��l��P�:���i�'k>�G��3630�I�i՛�蝱<�剫�Mێ�w����Gƭ������'f���I�'0��i�6mH&qUf7�&?i'e^�lr��I��$�.� � ԿEՆ�36�� C�qH>!.O�?�$���23��bž)JBXj�O~�l���s�<a���Ox��ARC�s�f]�!�R�Zp��`��>1$�i,7m�|�)�S6n�@��DJ&E� �t,�#꓉D���'o��-��V�|R]�pZ��D/n�n��6�d�JP�1�OLn�Aly��:Ғ��#�b��B��q�,�I/�MC�2�>�&�i��7��ݦ)xC�\�g��1w@����<Xb��E@�Im�t~�`ݮ5�L�S�x
�O׉?rl~�!��ۛV�j�YAI�y��'� �I�c"2�I�B@�TA�(���'���'�6-�;=���MH>!�PTX;�ɟ�@����Ӊ'�����FŔb_�ƛ����L&lo8ḵɜ�\�|�3DC�C�Lڦ�O��O ���'�N�{C
M�<p��!LZaچ@I���^æ52�ʍiy��'���:��KE�г�@�3J?�U;�C<?y�[�T(�44w�Fn5�4���� H��&B�S[���S�#��)�g윸(i���d!O�8�����#��O��H>�*P��Xu�&Ώ�c:��/e<���i����  k�QH���;e���Q$����'Y"6�2�ɕ���O8и�����Rd,�ڽ1��O�Dm��b�Z�l��<�OQ�l S�?��'3�r$N/1 �tQ�=h4~��'F�	џ���˟p�Iǟx�IJ�4"M�-�$Y�!�ɹ�$� �L�,N6�F�6�˓�?)���!m��CgZl���G�6 ��಍�tC��mZ��?QK<�'���'4��zܴ�y��
�M���y����D��"���y��̣7@��*b��'�	�����*Jw^�	�O�$IK2�@?gz��	ȟ���⟌�'^6M�L��$�O|���TRq)��4<]}k���
`\�*�O}m(�?�N<�#(]�xo>�0+�	0���*��<��)�H���<q�z��)O��)\��?I���O­"!l�1�p�h�n8�.1��f�O��D�O���O��}*��'�J�X3�E�3;���D`Ͳd�((!�"���c����'A�7�(�i��s��������FV�9�,P;7+��� Bx�:mZ��m��<a�oC� ��U�Ѫ�5gubъ���Sp����@	����d�O2���O��$�OH���|䎁��dLJ
��cޫ$��ʓ&'�f����	���c�Ӟ:�Hph����)�ص��oS�hh
��+O��d�O��O���Ob�C�Jʡq��NDܵ��J�d��G�� ���9`�(	S�AУOQ� ��!�N\ ru_*o,MԤL�n3��	���~\����t���ߜ
�P�h�aĐ`�f+Dm\�Bk=H3��,n��he��H��E�t��]��Tr��UP�����RUbeɔ�,�ḎSVjq���'8h �*B�d��T@	���q^>Iz"�\3=ʝ�b&ɲ|,F	��d��)�����"޼
J�j��E6��;��QE:}
�!ƬHD�����Q$?�)��(��
��f�F�R���< �!@��&b���%.Z<o���G|h�C��Ms�a��s�FEѓ�P�/���z���� �&^�x�	[��ޟ|��-^Z���Tp���H���&%�,ӄ0�'�b�'�2T��H&����OVp˱L!1G��*7R���O��m�IR���h�	�!�Ib�D�qL1Iq'_�?�v���Y1h����'�W� Ȕ����I�O��쟆�AEǗ��ȖJª8sj(s��R��ğ����&0��?��O��)�U���R�t#ŏ��l�$�ٴ��A�W��ho�<��۟��S����Ǝ@�1h�%y�� ���aь�Ʊi>��'��Ճa�� @�4[f�Z���fg	!�B7��0J�JToZ���I����S;���<��ə�'\����_hӰd���Z�U9�����O��?m�IC~l�d�,[�&���(~�A�ش�?���?Vʝ"L��ly2�'��$B*���iZ�v���#Ty��OX����>���Ol��Oys�Q��dY,����-bca�9�I ��ʬO,��?M>��O�n����uYh���F�����'�*� p�|r�'���'7��-�|�k�*�� �0E�I-��ܱ��	��$�<������?��Q8l�C��	;<	XhS��P㔹+d X����?����?�+O�����M�|:�(����E��2Ǥ�+�.���q�'�W�t�	ޟp��9VL��QBU���@�&���AK�-�'7��'�R]��C��>��)�OUSCV����NK�iذL	 ��e�IJ�	ǟ`���dcre�=�tG�O��UxgM�&t��S�צ��	����'�
����~z���?��')gr�؅�آGLu��e��bx����xb�'�Rm�$�b�|؟��քl��I�uJI�;����i��h��޴�?����?��3��i��X��J�K#~ ���F'>�U���uӚ�D�O��;��	b�'0�da&,J
�z���T�=��Xn�<Ɇ�3�4�?1���y�� e���4�ȸClr�X��Z��z��&
X� 7�(&��d�OF˓���<��9���CL�<��̀�(�d�zLR�idr�'��IB�O�	�O�����c� V����!�
�7Y��6��Oʓv�3UU?���L�I��
 A�->IB1 �f�.<��z2-���M��'��葲�x�OL�|Zwg�$x�#G <�3GƦ�R�OT�#�m�O`�O$���<!��\F����V4����o�J��C5�ǿ���O�$=�I០��.޶!�¥�rRft�w�ŸrF}�a��=R�b�$�Ivy��'SXX8�ݟp�(!�\3�$	1��)jf��r�i?b�'�O����OH��$$�#˛���;5�̘ �CB�09VM��Z��ē�?Y)O���R�6�˧�?1�f�&RXLx�&g��G�Qr�� �a+�V�D�O��d?6���ʱ�x2D8\����aUF�;���e�t�D�<a�O�&�/���d�O����6�&o���$������ ��qkU�x��'@b�6 .P��y���LR ~0���g c�D��!S����[S*,����l�Ih��byZwG�4[!	D�h��1x�!y�Va�4�?a��_ώ����u�S�')|�)3��n	1o̴tҰm�`��x�4�?��y�'o�����㏪_��D��aT�󲄱�
��
\�6��<	n��OZ���g~�(w�}I6�w�l��6Hr�6-�O��d�O�5Yi�<�O��%�:`0VJ�;N�~��$
�<~LL���\�B%���~����~R'X�g�����K#�HH5玚�M���fK�|�+O��O��O=� ���'��6F)rP@B�@�R� &�xO_;��d�OF���O �]��U�	��"ٜ���'6s ��p#%[��'m��'��'l�i��aá���Aa�/�ʴ�i�z�Ĺ<���?�����  -�'t{�a��J@	4*�� )�>P���'��'��'�i>�I?l�1��Ņ�+1(�E��a��E�>��?����D��v$�H$>9�%��eU��@k�XL��*�6�M�������4����%����Q�hRp�
�m!��[��M���D�O�@Pd��|����?)��&έQP*����j���Z�"N�����'��py���z<���'`ب��N��[�|5���i��	�D��<�ܴ]���<��9����
f�F:���X5��� 6���'��g��7�r�~"���.���h�<Ը��2%�Z�&��4�M{�!ZAX���';2=O��f+�4�k�]~�!ŉ5X��Bi�`�֪?���'_�'�TZ>}�O6��9c恼#!�h8��a���
#|�h�d�O �$�}@b�S��>a�-Db���څ���ef�����i&1O�d��A�[���|��ǟ��a���]�|�
e��;wL��Ӓ���M��'��}:Оx�O�B�|Zw3|e�R퐾Av���J�4oU��OR$� ��O�˓�?!���?1/O�Ƞp��X�Ɉ��#%<t	�t���x0$���I�����py��'���2g�E��^d�\�ř�W7��d�'��	ڟ|����p�'���s�-`>U�w�7=W:H@�ˍ<a֊�a�)r�~˓�?).O|���O��$fg�d�o����� ���î1|[��o�ԟ$�IڟT�I_y�̉��ꧺ?��GO�MQvqoL$_����
͒F2���'2�I��0�����J��v����c?��X<}�>�;� �;5��bK���ӟ��'���B�~
��?���j������aR�=�gd�`�0h�S�������6?\��Iq�IXZ�I�)Z$h���� iL�zqRߦ1�'�~x@c&tӂ���O&���<�֧ug�T*m�<9����1&B�1��"�MC��?�4K�<��?���ԸO��A��K��-0���˚#� ��ݴH	��r��iX2�'���O�ꓵ�MX,�X���JG�RV�
�l�6�nڷD�>���X�'b�D����%$Lx�RY%JE��k.t�ynZϟ �	韌� �����<���~��;�ux�� �����n���Mk��?�����L�S���'"�'e�4R�,�4裶H�0K�v �FldӐ���R���'��I����'�Zc� @e����X +-��[�O舫�4OT���Or�D�O�d�<��	ʦ(�2�"rf�T��a�@��V�hJ�\���'��[���I˟4�I\7�Q	 �
�<�['A	�(B���r���'62�'F�R��Jw.�����A`$P��Lz�ʼ�B@�MS*O ���<Y���?��J���$&z)��с�Ԕ�s�Z�!�t� �S����ٟH�IQy2�g�q"����D`ӌ��җ���b� JN�K�4�?a*O�D�OF�d����x?YF�Y;O_����P@�Zh0���e��ڟ�'}0U�Q½~r��?)��n��SC��=�������rY�@�	��d��Y@l�IFy2�'_�IڀV��LC����
�9�|���Z��S���6�MC��?I���X��,)gd�r��H5t3r���6N�<6��O4��<^�D�O����O�F��m�/n����Uf[�Ci���شi
�:�i?R�'�2�O�����DZ�R\:y�5%J����h^��llZ
}L�Xy�'���ĕ�+eE��(X<|��)�l�V�.�oZ�$�	��!Oֻ��$�<Q��~�"��ڐ��/A
w��
4#��M����D
��?A������I�"ظ6Z)<�ڀǁ4]��,*ش�?IdF�>��`y��'o�����*� ԑ�Ay��u2#g}y��L��1��?����?Y��?�+O�� c��_��-`��YZvh;�j\*=1V��'|�����'}��'��A66%$����K=t)pZ�jW�D74ᰛ'k��'���'�V�Xytѷ����$�Nxz��Ǧ�,�se���M�,O��ľ<����?���2�8�O��(3�&l% I��	��Q���ܴ�?���?9���D�=�t��O�Zc�T���Z�(��@a�k�پ��4�?Q+O����Oj���%$"�|nZii��b2N[�vi�Z��C)y7��O���<��kǴ@{�؟��	�?��3��A�<���f������%�����O����O�"�;O���?��O���: X!r<�Z�h�3H����4��dΏkRrLn���	៬�S0����~Ij�BP4��)�����
����?I�]i�q̓�?q+O0�>A��뜥m�,�	�A��#z�����LC�mLŦ���ʟ<�	�?m��OFʓ@�1���N�!-�z�S�S*ر�i9���OJ˓��O�
6v������p!KX��7-�O,��OT0Ks}�Y�,�I\?!���]N��X��\����K�ʦ�$�S�u��'�?������� �AN̽��Z.ǚ�YPj>�M����|T�S���'V"U���i�m��%s�L�K�%�3 ���A#�j�D�d�rW�<)���?a����](x��["NU%c�y�W��6TzQAn}}�]�p�	ny��'���'9�0iև��~	�� �%cr���Cۻ�yb�'�B�'!R�'��I�F�vP˞O�d��'�,m?�P˷�]��۴���O���?���?!� ��<��� �)4��7S�(x*&nT��4Ѵi���'�b�'#�PJ>���V���;-nk3G��$��U� *t�Tn����'���'���	�y"�'H�dQ�S"�|S`$�<ʎ�c�L$/����'�W�|:Uٓ��)�OZ����n��d��s���⁗4+�p��Ma}��'�R�'r���'u��':�֟az�l�3o�l�1�ϭC�����i��	�"l��ݴ�?1���?A�'l��i��YB'�6�&�F���@Ejc�����O�;&:OXm�Oo�IU�l����p�X�*���p�߳@ݛ��Y�R�h7��OL��O ���m}�R���WiA�g����`Z�f�vЊ��Ǣ�M{hz~b[������\ϖ�٧�׊�v�`�A6I�N����i���'"dǷ6�2ꓙ�d�O<�	?|%"�Q�`�
\u����pIi׿i$�P���P�|��'�?�����B>�:H�*��Z���Q�����M��%���Qb[�8�'+�U�<�i��9���"�>���d�-���D̸>ɣ��<A���?����?�����$i-��ѡݟY�2wʋ2;�����"�a��֟��	n�֟���j~����(��v�
s�LQ&�;U����'Pb�'��O-0ZƂt>5�e��0�����h�rH���/���Oz�O���On��`�OjQ��^;~R�}9��X�$��`%XR}��'�R�'��I(JX\xI|��._��٨�	9,���$�UG�V�'��'�B�'4���}�.��n`�E2�lÑp�V �󮚛�Mc��?1*O&x:H�w���,���n��9�,�6~���`�@:��N<����?Yg,�<�N>�O^��s�J��.�y��Y .'Ę�4��� �3�v}m ��	�O<�iW~2'E��tٲE�y7��{1� ��MC��?q �_�<�H>9��TO��t��m�4;:���D-�M+ӭ[Eu��'f�'}�$�.��O8x���H���׵;�]7�7�ޙJ��d4��(��̟H,/T�����:[��`4.�,CB�o��t��ោ��n� ��'@"�OnP���p�xp�`�@6Y#e�9w�J�OV���O��dY.'�\�S���:3���PA�+ F�ho�ʟ�I����ē�?a�����C���vM\R"��~��\�".g}E�0�y�W����ş��I_y¥�*�j�VÊn}�$pG�E8Nx����6��˟�%�T��˟�q��t�f��Fʖ6�Б�p�](K-�b���	����	zyBh�4wI*�ӈ0w��I6�����S�\7D�O���&�D�O��dɎ%�d��Α�J=�#�P�O�mi7��3D���'���'Q2\���l��ħPϼ ��=.=2�)�J�K��T���i�Ҕ|��'��×� �B�>��ʫ8����E�_H��B���	㟤�'��5��5������+��f	O�;�ej"'�"Kܨu�'y�'�J�g�O����VrQ36N�z�,q����)��6m�<y���{�FI�~������ta��M�J��x�$��
?�h��Am�2���O��PF�O0�OF�>��vK_
�)Qu�%����Ӌl�"t�@���I���I�?�HN<�'@�zE�����QFe�Ӄ��kE.0A!U� �	[�Ş�?a�oX�����%�%PV&�9���qb���'��'�~�Ȱ ,�4�l�'���i��׍0�r��'�B�Y$�Aڴ��'w������OL��O�*2�����[�2h×.�	v'��l�џ<��S����|r���_OgA��L�^��TKſ	#��Y��Isy��'
B�'�"�'fJ���,�zQ"u����?���vNA���	͟���<'���a?A3.ȆX�6�����6L�.a2��Xڦ�"�$?A���?������=zX�ͧ^�2�����J�� +;pܘ��'�R�'R����1��S�?ծq�b(/j��x���I�>��?���?���?�k	5��鲟ؒs�
^��9� �#f�� ���L��5���ON˓{~��$�4�aN߂ Ā�A�6᦬�mjӈ���OJ� ��p����'��dO�
J���e�C�R�Ԝ��ưA$�Oj���O�IB��I
�B�BL����P�c`�ѦE�'�~�R����꧓?���Y%�	,��%�ŉ�;~>L���>e�6��O:���V%���}���#_g
 ���EG�uM\Цq���Ο��I`y��O)2�'��I/F�~����46$J�%.@�O6��)�ޟ����NN�#b-ȇX��i见ݦ�M[��?٘'6����x�Oz�'�:գ3%*H���R.e�
iQ�#�	.��c�����H���\u
8����QO�q������A�ش�?��1��F���'^�'��B�9T�#�.L080YD"�ݞ#g�	ڟl�I�Ĕ'�<�)W�RPgq�Ҹ&�0Q2ILr�*O��D�OZ�O��d�O�-#��
�l�S*U�� ��.W�1O�D�Oj��<�R(���)A2Έ5p6�E��@h� ��	��IA�I���ܴ�2�D�ӨÃ�z��!�s�ZQ�']2�'"�Z�4Z�"Y��ħQ��ۇ*�$]�>@a LB:$;�8���i���|2�'��ˉ��'q� [BN�
��@E�C* �;�4�?�����$�:rP %>��I�?A[���nk�8����;Kg�iۀ�����?���tN�QGx��� ��)��z�~ YG��Œ5W���	�s�l������	�� �SRyZwQ��vm�v��cQ$�-?���ڴ�?Q(O�S�)��}�J� �j�F]z'�mL�vJQ:<X7��O��$�O.���k����؃�!��������әw�����CX9��?I�^�|��ʇv��c/�,d��=Kq�i��'w���#g�c�d�Ip?��ŀ�_�yX#��1�� �(�T؞��ß���IDn�B�G�I���Q+�fDJi��4�?�s�M��'��'�ɧ5�Z�EHUɋ9`���"�ٷy�R�*��$�<���?����򄚑Gڪ����.H��h�3M!~Q���_��x�Io���|�	�?���fB��F����A`�>��4�*hc��ӧ���+~��T����'Q]yE��-d�⭊'�3�=�ȓ8G A�Ī�0qB�W0>@��"e#�I� �@���ΓL(������b����"���li� (_��5P�Y��"͓'(��6$P�R�J\i�J��'O� �2k�<�P��T�"��-R�/��L�pV��&�J� 2D)W��A�a6pw� �a.
.�x���OY�cQ����@��&��@)Q�@�c������5$���>m��"�&�[j��,����Ob��ֆK��n! �\�m�]#�۴���]>�1���?_(蛖�J�h�cQ�>}2�� ��Q���^��ڝ���˝O�.�B`��DI�>c��a[��o�������|���'�(5j��?Q����O��
��N�WZ�1�ѾX���S�"O�IAָ�c⌕6}Ђ���h��poaxr�%ғ2��{�ÎOJE�
�#g�I3Q�\����T�Q*_0t�}��ğ�I��]�j7����L�"8sB��b��M�u!��z����O|8�E��w�1��'9,P�ȩ�����@wif-�L,s#��O�a�������p���{���+'BbS�B�
�������D^� /�Oў�Z2��v岉S�����ݻwo8D����A�d��t��*��e��K"?1�)
.Op8Z2<
�ȵb�")�)�@ �,I�v7��OX���O��dܺ+��?��O����wo�/fY6,aՇ�1zf���nD�N��}�cǀd0�`��'�4��� O��f�:&i� �#銨`.��ShR8Q�$�R�'g(����E�u�����MP ��Hɨ�?����hO�⟜8@�M($��‽)r*8Y1�,D�����!c�: 0AbL�8�p���+���d�<�� ϕ�	�����T1jCn%����4v���s�G�T�IŊ�	����'B,��h��+E�J��`��"�M��m�A�6��iL2*L!�OUN8���7#��01�dY�#���k���q��ؐ���lti��&O��:�'Q�^�l"���@m�i� s�:��/$�IA�����8s�D��Q�ȧ^|`0j��#� �ݴDĆ��&�3yF�$��3BM��͓��D��5�'��\>q���L� �֭���\p��Fŕq�l��Lğ8�	��`��
*����ū(�?�OG哆pJ��
#�6��	Sd�H�K0��'<�5ZU�-� ��h1k�>�JPj�.b�jdC���#ydx[Wj5}�&M��?a���h�n���*K�*�1�g]���3�A�D�!�dQ�Ss�beg��P󢀫��@U�ax�/ғ`�ld8�D+x
��҂��y��Y9�V����џ\��O6L�2��	�������]/[�iW#D���u+�!���q�C��fe��i��W�srl8o�g��#:F���E?M��� C��Ƚ��ד O�<rG�׌ [�}��I0�I≴VO������4CYXʥ�٬a�2�1ݴ+�副T���4����:�	W�|@E�
�}Z��'",�C�	Cg�H�%u¦`�c՚B�T�C����O
�O8��4���3 �鳪G?O�4*���<"8���?����?���6�$�O�����0L�v�/o�j@�d%�� zQ�ge�]�~�FY�ZT�hN�RV8��Cȓ��`�fƅ��>�+T��%�����c�,���µ]�bIQdM�5
\�@���'�B�6��O��d!��1i�p�Y@BԋKb���a�6Cq��#�ēJ��u͓��x��y:ׁV:I]J��HB�)�/O&��_}b[�8B"���M���?y��^����(q���1�����1�?I��N�Jhy��?�O�|x����'/^C*��w�&(�g�΅&v^���9,B�P
1@|�;S�4�\�p9OF�U�'0�X�����O'�H �GTM(2I�c`w�<��Ɵ��?E�d��+
B<�`F�G����6��C(<I��ik)�.P�1�*T �EB�2Z�Y��'�ў"~�)�D�(������BM��(W�<qWI�7qe��MΧ�X��/_W�<)2�T��,�8�
�E2����GL_�<��L�q:��ҕ!�z�Qwc�Q�<� ��ARCD�$�h���ބI~�!0�"O ��7��+
}�҇�Jy΍0�"ONHC�GV�e���;�Ϲ2��xj�"O6���d�0m��eB7w�n��@"O�(H�$�F$h����պ�"O���p��[�&�i�DѬV���"O���B�ZR�bq��Y?r=@�"O����L�BT�+t�Ȱo�D���"O��[d�ПE�)�S,	�O�.�(A"O\:��Nk�!�a��I�H��0"O�����D:�!��¯k~��p"O�4 a�33Z�W�7ndu�"O~��4���< ��+�`��mx�"OV����5bN�]iAd�z~pi��"O<8Y	c���C�� ����"O���7���J�zCI�7�"%�"OԲA�ǓEP�bAB�	hȺ8g"O#$�P�q@p-�TaL|9;�"O�A8���qh2�O.Az�qw"O���q�^�#mh z%� aԠJ�"O����J,41�K�lW�v���'"OD�8q��7�h,Ɉn��sp"O�՛��F�Y�x)�e�եt��;7"O��r�L�0�T����t[`D d"Od����N?i��A�U5-' ���"O
�x�c����"�%\6$�@�t"O�9$��L�fU���ɖ:���a�"O�M�'�'�M{ƀ���H��U"O�݈5,ߜ++go��m�ȅ��"OҸ�L�T�����-8~$�sQ"O(�3gP/�"�P�o�3,iT$��"O��1`Aut�ܩ��1BH5�F"O�P8�僕z^.qA��*(���"O�X�c�`�,U(c Q���c"O�)�q���0=��`���^��-9�"O�Q���u֩�4!Mwc �"O򧠆�	fp��"�^�~Tz�"OL[��,R�L�1��kjL��"Of4���W�P��=Q�Q����"O�k0C!�r��
�W��1�"OVX����^|B9��M��b��!A	�'P<[uT$�X&Hק �qj�):D�(ᶏ� �N��r��j(�rB3D����+U1<�j�@�Чae@ sĩ=D�,����9�TEP�kY��J�:D���Ď�3W��0[����T�T 6D�4��W9"0�Jrퟍz����	3D�����A�!l��r�]��4ԨF�2ړN7h]#P�6<�n��5�>n�	�w��%?�fC�ɵn��(A�B0�f�^�5$,��G�L7h�R�{���F8}堸���I|U�/\��C�	?p����N�pƔ�.�a���	n�X�"lOh�t ڋ$�V�c%�܇�D����'�T͐D�WӦ�yAF	�	#��1IȜz��R�5D���DIۇR�&\��J���1O.�FzR듊(���1�k�#~n�4����y�/�1|(qR��K76d��C߷�y"�P�[������G�Iւ��ā�(�y�J<)Z���$�	R���ªL��y��	����M�w�-�w��5�yr�\��$�ˇL��ZS�lI  �y�CҽJ���s΁.IO��'$ޕ�yb��#��%Y�JS��Ri���y�/��a��aZ�ؘ4����5�y
� �-��KÆP!��f$"��l"O6��e i���dɃb���6"O���U�ANdZ'��V� �3"OTIC0�H8` ,p3�٦0��y�"O��Y0 C[{��' �5��=��"O,)yCȘ�X_��#6�4%��)��"OR�◭ۺ�a �B�"N���"O�(�t��8���($�QlҀ"O�Y��^�*���!� �R�"O�Ur�(��B��T���L�f�'�R�����4i��3ǀ�%=�L����P�!��^���a�PK�n�"��'�pt����3Op\��Bϝ u�i��Z	^�!�*Az����ص>^0!9�!�V��O$�ZB*4O^(��nΣk4x�;&�)��@pO���R��Z~K�J8���#��z\�qOjM:T�̭=]R0:�C� .Y��צGm���S%a}"�S���'O`b��7D�y�<�P�Y4Z2.�HG�;D����-�j��9+si���>̙��y��1�&��6�V9+ۓ|�D�D�Q80�bP��ą��*���N�{�d�۴Q���N۱0S2UZ�/Bl�.q�ȓm�40�"N���W���V���<Qע��R���VM1+��>Y!D�B�/�� 1���$`EI)�.?D�к0d�V�#
yF��Q�k�; @Fh�����YS>�_�%B�bՍ��<a4N��}U䌆ȓ
 u��Z2G�`0�Q�H��Y��Q5�3T�a{���g1���G � �̴9��ބ�0=a Cmn�<��o�)@|�V��"��eS����Q��k���y���-�)�1�\�yef�SgI�Ә'mv,��gH�W���r�.9ҧc*,��ϙ�+��]�ĆW/���ȓm`� &�Ҧq�:��%$�7�Rh� dz8MZW_��!B2�g~�M�np.<�SL�
+4
h�/�:�y"B�y�d���!VR�nl� j�#\�0���H��Yr�`�'lOzLI��/BQ����K)\\�r�'�H������t��Uck������ 1u� *�3t�a)�"O�5#	�9U�pX
R�o`\���S� gp|�V��X;��D���9�8H���IqR���c��y2��d��Q�D��F����)��+��	FK�O�|�J�d�D��O~�1������S�۩Y��3R"O�%��$�2U"}� n�)�X�
G�	3�%��� �퉴.6�B@��x�"��SO�%l�B�1;r������ �0�7����C䉷1
!B��NH �냀B�J��C�ɏw#tq�`�~��x�0(��
�HC�	�p54��t$T�7\�����'C�C�	6~��%��JS���X	����'�ЈIPc�:�(�)�
�0}A�'�Rxre��/>r@��*�=z��R�'�f���G��ؠ!ᄥ
1�%��'�R�xB�6z�)���1P�0<j'/�L�����P
]��y2Ĥ,#��ɣ������Į^��&ᅦ�\�ȓvF��lM�FSn͊V�@��Ή�+~��c��2a�ƌx��
��?)��8����1E�=�c�ˏ2<z�"&�'�ݲ#�'}r�ْ�(�BGa֍b&�����3I��)�4h(͸��?:H��9�����%�d�='��`2(���8Mۀ�O�z4��q�fP,fBY�ɶ	���G��a����0�U8u�֔a�'��KT��"�/N�L��kLۦ��h���V���a���O�E�D!��rx����z&�qa�"\O���U)���̍��4*N��Cw�:Ų�Ð�U|\6�Щ4�,PJ�#O5����c@%��<�w)�d��u��H��O|a���΅��܈�M�LChPgb��- /��д��D�q.f	�U
ӓ��Hq�i�	�$��N?I�'�T��LT�fr��QD��A߮]*��O��#�ŉ�HM����}�Ԕ?UAql��<��0`�p�$[�v7-â1�A��,gQ�D���4F�˞w�>�[g�˟_�|���"L����C�5������]����]�L��OL�p�]	4����[�|iZ��	CʔB���7SlHw�+��.[�  �{m����`�o��(@�^ɲӎ	����"B�s�����S�? Ρˡ���A#v�1��S)e��;$��X�
)Y�j�Z�'J(���1������un���p�W�f9Ĕ�Fɜn��Y��K;KW~$kK]�*�x�J��V$��2](������"�#9� tt�0b��J��M�'�X��)U� �}�"�[`q�%C��6\�9"�J�	59*��w���W�bu�caj�Ő%E[;naA�㔺\��x�ݪoŎ�Y�@L���)�c��ƭ�R�ȹ�ą��x� 24�Oލ�*%�	�2�.�B�L���� �JX�F)�tQ�5�D@ށJ��E���tU�T��>nT�sEI69/���OdQ�r�S�
1O>�b�лDhp���	��@����G	�G���3(����p�g��vM�"H�5�8Ӏ� ]y2ܙF4�vH+�i�5Մ�m���r��L�����.Ғ� ��3ǌ��'>��3�6r�nU�����ji�شY���D*�=h:)R��Z�gJ�R� @�p�$=˔)�w)<}B�D7��(Q��B�'��P�P��$�1،0i� K�M .����N-B"Q������ �B+O���@# �Q1j�S�-����Ƹ���%`� �R�k?~D�+�^�g7<P ��5=���Oԟr@�4yr�3��S�E� �Q�cu�)�CM<Z�8�R$*�9T�ȉ|A�Ƨ�O?7m�4/-�-9�,��`��y6+Ô6��I���+O��I�)ȌL����;:(@<�G���p������T�|���O�)hB�I��J'��W�,OV4;�F�o�P�z��^=~5��N�h�,P�&���'TƬ�#J
�z���`�)נx�ܴU9ĉ@�Rqu|��ł�(-)v,��@���iU��9��'�hQ��?��Жjײ^�5�,O��!b֫(f���P�Z��2�=b�f��f��!=� ĩa��բE(ܜ7�L0��Py�O?����"��W�+f!ȍ+�:��-=��x{a)�"���ڵ
��0<4m#_���1v�H�
��-x�g4S��C����>����m�9+��mæ`�,B������x�43�`�K����r�'�Mau�E����i׿s�Ub�g�(7\6��C�O.E��$K6���p�m�-}z�dǟ{�u"wg�J?!�+��M�4�]/�.ݳ�b��}�vPƧRG�!��"]� �Bc��`X (�X���%�:9�a"�)�'}��Ѭ��J���0#y�A��~I$�[ū�wqX��%k�8�
M$����c�2<�ay��(���@����tT]�e�E��xB�, n8H�O��h��M�KӞO21���'$��p&Ζ5V�pȇ�K�ةH�j D�����\(5T^ģ����1qUA+D�h)����~yi�aa	KIh��(D��b�#++�8;THX�����D#D�4r�Q&E[
�s��V<dk�Mb1$4D� �q-�!�쁰�:'6n-��)3D��x��M�k����)ݘSL��%�/D���cX��6�f�=u�,�c�a;D�x
wh�,���D�Q!�b�i7D��R�LF8^܆t�gdđ_+�q��)6D����Φ��ف!���/�U��J5D��IS�:^G�Lka����N-B1,8D�$��͊7T�Q)�%�� 񺥮1D��je���?
��c�H#|6mKT�+D� ��-�8
(���a!��q�eH%,?D�81ԃ�ʸɅ�,8��9$n/D���D�ґyb2Q;�b�wV��b&k+D�|BHӇ=�lJ5�F"d����37D���n��K]ތ���<0�����3D��ڀM�-%�� Hת��~G��u�0D��( *�a���[��#��k�c0D�� ��ڃ^+R��L�[y��y� ;D�,R��x/VP1���}N���#4D�ɣ/�>�����c�j A�(/D��i�F�)R��4+�E�->�N���-D���.L�\�x�fX54�J��)D�XR,"%FPyf�/ p`��)D����Ŝ�$dˁ��FF��-'D����k�JJ�e�FA�USv��1D#D�S���`A��P��!eur���,D����q�ЕO]�B�S3�*D����ܐx�8�S!�Z+���*�'D�x��g�n�y��)ׇ(ޘ2n7D�ܡ֌L�zN ���_���j9D�$�f���Dz���r�؊~����5D�� J��B�\ @ �K	�K>���7"O@`��E�Bp�Hz���T*"�[w"O>��$dK /�����dD�/�H"O6x��.	*z��QH��H��Ia�"Ob���]C��6I=/�F�k$D��PЁ�1S�0�*�^&,�-���$D���S�3^^��b��']�4LB��>D�d����:���x4�C�*�p�z7�:D�<{���=	�+�}�8{9D��	'GA�,<��'� j�9D�PjN��G�Z�j�+�8~¦R�9D��dV���� �!�x���6D�أ���-&E�R���4M�(*r�4D����C٨/ ��`1�"�bp��1D�<�2��"2����E�?�(�1C:D��#
�<9�x�S��i�JX�e�+D�t���@��, �Q�Le��z�*D���Ug � 3j�`t!ҥ��d�-6D��
�@��:��=2��Ψ�����g'D�8���Z�Nq3���1|�N�0�(D������(L(�t�iʲ: L�
�e(D�x"ga�9F��a7%��J�.qA�"*D�T"ޥ@��9�3��a���&D���D��g��T�:�!f�$D��(T�Y��� �%�_��,@Ä/D�d�i�(P�z!)sI��� ��h3D�X�T@�*���D�Y(Wm����<D�4�u���Y$B�
&�|���h7D�T�!h�/�,ەi\B[�AUO"D��#�'�+/�6�kao�#��ewd:D�D:�E�!�rآG�új��0`�#D��@n��J���ÿz��	��#D����-�+|� D���0Cx�21A!D��b��7CdpAK��JT}97�+D��Y���7@�ɣ�+�lH2	x�e)D�\��A=pyT���T:?�1��(D��ga�P��f�Q67+��H�#D�$�P���b���hr/�;		�hb�"D����Ň1I�����:�
=�"D�"��FC`�u(Cj_,U}�(© D��
WkNW���3ś,"Y8D#b�?D�P8%��&�=z����B����<D�T����*�0�z���7]�0�-D�Xk�"ۻq�Rmy��R>����� %D�,� �j{�Ѷ�2ZGR�%D�D���,
A��F��9��B'B�hO?�$�A�2�Yd��cEt�d ��!���$�\
�PS�G�u��C"Obe��,� �5���%��`"O���V#�(v	,��#�M#�ViQ"O�`Qg��/V�,�ǃ����"Oj�[�nߙ3� �b�A�����Id�O="c7��>��	���&+*�3��OF�s0D\0w�L%2W
}N���"O��9F���u�̉Rꀠ!�hI�b"Ol����<\%p`��
�&�!��"O�a;!���v-��V���0J"OV1Y�σl�Bȓ��
�6/P؊C"O&�0v,Õs��TbK�0-��""O��pr��8r#�Ʀ[*�	�"O�Mٶ�$��ce/	�?Yf)
r"O�p���%1��㔨J��`��"O�U�ð+m�I#W�Z�jq`�:1"O�U '���pz�&0l<��V"O� ��2��B��hR���et���"O���=L��0� �46�ҙ�@"OD�i��6���]�+v:UiB"O�q�lS1MJ�����,W|�Y�"Oxa�dY�pd������86e�7"OX-��Hڹ+`,��/�� �"O�(�tSq��\s!���)��"O:����M�,H�@e����3"Oh��c�f��ӊ�_y\�2"O���tm�p2T��ë�"W�(�g"O� ����?g{�ț�� �T�"O�K��(���q�Z�Hɪ��S"O� q�HMh_�����m��XӦ"OdY�lT=//�4#w�I�g�0�1�"O���P-�/tŉ��]���ae"O�0'*G�>��P�?w��	+T"O\K4�+	6�@�ϐ�>��y�"OT<*a��=8xHz���/u�r`��"O���\)5�����!����"O�i���5$�l��/��LPg�'��'�y�@����p���{�l\�
�':��V��ndh�"�	�#7v%�
�'��c ��1DwjL��-!X,L�	�'p�Y����p�|1"� ��n7��9�'��d3ΐ�5�hă���7���+�'����R7|z��c��.y�s�'i�1sv��;�P���.�)�';4���GT�1�.�R�A�E�$d��'�(���0oX���B�<D&�\�	�'��atM�����Ã6ö�1	�'VJ�����\f��b�#?/=֙��'��|����)�j������7Հ8x�'t1��J7.����Y�*�>�)�'�&E#P�ƙL����Mה/ֲ �'/��ucr��ꑈR�&��(s
�',�3DH�0^lکсL�,T��
듡�I�}wBL)�dJ�)o(t����xB剟%uU�t��ó&کa}!�$�a���IQ����j}jĢ�
�!�d�3b�`p�B��&-�ܐ����n�!��/8��:#B ��$E�!+�!�9D��HQ��@}�Ȗi�g�!���J��ځA�+`8i��NV!���*3�\���3|D\m�֯V`!�D��k�>���L�Y`�1q��^�9\!�D���s�kNOA��F�^8y�!��<b*��	@C 4����)]!!�d!G�,l�!n]���H�k��]!��A��B֭5~����IT�P�!򄎟J@C�Z�z�H3�K(zKQ��E�$@22�� )$��/��@�dˌ�yR��1.��mW�|���ٹ�y��K�/C^�YR̅/V�B��ꃒ�y�hT�����LB�O@��R�:�y2ǌ�tX�c@R�: y)A#��y"�Z�{\8x��X�7z9"@�K �O<�=�O�.����%>�`�¥&v��i�'ܸ�9�ŋU�2Uab%f���'�8��R-�����XI- �)�'�l�9`*��r��(p	�u�\e[�'y�]��DW/��ˇd ;n@��'l�\����h�.�q�AW+��TY�'+|tA'�7h�"�����pZ�'�@�R�P.����������� 2,H�o��n�{���-����"O~!3ՅVNF�0���)&*l��B"O����E�hnPm���F&5��"O��b	DL���hKH�#Xq("O�ݘ$ J�z0B�䄌C��C"O�y�b&�	Ԕ��0� �f�X!S�"O���4�>�H�b%�R90�E�"OM��B3�t`�O��
��h�6"O��H��8�x8
�+F�H/�\��"Oܔ�T�I,��0h�i�4�0��"OH,��
�'3��b����1�"OpM�����8�"O�+��|��"O(���Ae�<-(�װb�\�A�"O�i��*dA ���Y��(�`"On�z����BIT?�4����~"�)�'�,�-�DC�%����sf���W��	ʤhc�\ Qf�z%���B
X0��hW�p�h�1��̫�l�ȓ%�(�JSE���)DHӥJq^���F�܄٦˰v�4y�BG� �D�ȓ>0��$K�1�x�4�N� �ȓo��h�9��+L�E=D�h��!I����RC��I�i�� D���$�xX�$9e���x�[`,=D��j�"_�| ��) ���6��d���:D�,�bIB2��!��oH^��p�+D������C��A�m\.zFB Q��5D���"�Ƴ B�;a/��e�J�C�
4D���@�Z���2�'�.0�l0D�
�	P�'.4H`F
L\���`3D�8[f��9$�ػ� 
�%;�9	t�4D���vG԰~a����	P�yt�?D�(L�DW�Y+�e�I!<@QF�;D�<����[��RU�֣9�b%?D��!ꁁ[3>E{T+ѷ_����':D�����?OYh�M��Ac`	�@�#D��X��	�.<b`�t�	��,a� �!D� �6��A��kΜ?a�*��9D��QqNA)%*�!�F��`�4dQ-6D��	�jX9 l��8CD��X��"8D��jB-�[�8q;֫*Y�꽳�m"D�h@2o���|�x����*����� D�0��N>�,=X`i��
3���D:D����K�a���G&K�M'�񋠬6D���LځIHV��`ɒ]Z� 5G?D���Ή�F���:(<Ai5%?D��9�"�lF\�p���4���J>D�x�d�#7��#�0*����c1D����)�d��� �e���0D�����˓�40�7 �;��z�//D�T��$Ҿ	�ABе&�| Db9D�d�G
ff)1%J�ΐ�9D���DiJȪ�(D0 ����4D��Z���++ܠ����Î����.D�<�CΞ�v z!���j���K!D� #�>M{��+���� jH���n;D��c��]�xIH�[����,��Q�,D�D��..Jd�P�2PX3po?D��+� bv|%�PiC ���E�7D��@��%H�XD� 8{\��Jsm4D���s��#U�B��/˝c(R�XF5D�8�tO?`֐��(^nZD��.D������sh�i(J�1-����c:D��#G�L:��ac�
	f�
��9D�� D������ON~��ɍNs�(
P"Or5��I4p���βB�n�E"O>���$�/G���΀\f�,��"O~3f��6B�(�a�L)b�*O����M� �� ���,�Q�'��T���9ij ��e�2J���B�hPN�}���kC�$+�DC�	&[D�qu��K�\��1l�+KzB��X��=%>���s�lʮ�ZB�I�+�~��u?(X�q�"݆<��B�I�[{��󃈙y,��T$ۙ61�B�7<N�ұȃ��=�&˃n
�B�ɲ546�J̸ׂ"��A��׌9�DB�	�8Q�=�Q"W:C}b�p��B
K�2B�I�&X��L
R9y$$�	TBC��7~DHi�`���6�S'V/_6C�I;D���R��̩M+��R��S8/��B�	1@;������-lZ�8U
�>btB�	�� ���;}AP9�&K�W�nB�	~;$`�M�v(\�AP˼n�FB�	�0�A$B�&S�D �FΖ2
��C��,$%�%�QNZc��P�D�Qq�B�	C�� '�wc���d���B�	��8����B�NY�B`6D�Pk���q���Q֭Ŋ��(yf�2D���%`��\��8�f��9ܪT9C%<D�B�B�5(�x�lG|z
=D�\)AC!$|�E��Ԇ7�m���/D����H#u�����O��p�왵D/D�Л�BC34��ɫs�ڿ|�d��2D�� ��O�/ł���&�(�4͹��0D�<���Y;_��̻b�U�9� /D� �A!���M^6*�
�a�,D��[��U��I	��<?����7�)D�����
&ZcR}A��Z.�D��L-D�9��K�0��cf�/Ԅ%�@,D�d)�C����$�A�P�l%Q�=D���N�J#�[�j_�ux%q`+9D��V�R;B�:Փ��b&�ɚ6D�$�T@\�9����p��a�d5h$�&D��W���-=�ePӅ
-���!�8D���˜�]���w�͚4��� �)D��X2$�!����
g���n(D�d��O�z���ׅ�1P}2t;#&D���Ġ��3�j�@��@�����#6D�`Jb▏~�&�R0��3m`�}�@5D�H�P���L�x�
R>�i�co-D���'%G.!��A�󫆊���ڄ�,D�Шף3Q	��FD;W	�����(D�(�Ï?#��\�F㖽7��qF9D���@��~p�̨�
�2P���`7D�,Ge�j0�`��m6�-I��4D�����!�Ub�A�n��qp@2D����bJ�Xq��NL	 bR�P7�-D�l8AJ@3�� ��ɒ}�XUB"i)D�b$�/5�<)y�E�*I�Txנ(D�$!��K>@1�tG�s�P�*R`&D�P�U�A xZh���9P�<�&�(D�T�p΃w�ؼ��)�&|xҘ6�;D��3�HU�s �y�DN<O����f�4D��9CM�K�ɠ!��<�:B�(1D���Ā�~x<Ї�ܿF�$@��h+D����%L=z?��A@�[U<5�wn-D���eӁ&�1�7�_�!��h!�� �В�h�&��A�O�!uLѓQ"Oڌ�� ��8ɶ�^QeLq6"Oxq� $6Ia�N�W��|
�"O�5��K{���pm�M�>��G"O�,(G�èLeN�RQ��+y���"O���倎�G@L�:�	�2 �1"O-Bg�*��0�D��$P����"O��eCQ5��Y��"!��髀"Ol�9���
�ܸ 7�Ⱦ3����"O|��@�Ij�h$E�I�q`!"O����6~��#坦5g�]��"O@�S4�A�[���z�#*P>@c"O�\b��1��yrB�$A_N�1F"O�%;�!&��9&@Zz�V"O�� 7��6��#HY}I�ҥ"O�Q�bk�@�������=2�)�"O�œ�B73t�	/�7*R J�"O q�L��]b����$�*P��5"O�����?	Bh��$�7!޵j�"OX�n&EN�4"`$&&�r"Ob�����(p��Es��#%�`r%"O�x��&Ӭp�^�;U$��l#"OU����/��,��iV$�@)�w"OLt�&���1	�s� >t�ٳ�"OJjsH)/��!PFQ7iv���"Oj4	3e���)x��s�
1A"O�\,�G��bt��,p�$��"O�� �&"��4J
��J܊�"O`�����QMx���D$!|��X1"O\%z�%ɬjL4}JVa�< `@��"O|�[��;Rv��7"EaШ�S"Op�[#K�?X�$�Qbצj:nɁ"O>��4�J�Z��"��"G��]��"OFq�r��=@���cb_�^���9�"O�5��F��")���KՋx��w"O�|p��J�o�t�Q����4�e"O����	7�Cu�W�c*�x��"OF�ÓB�_��!��3y����"O:�!C�K "?T��d�������yB!٩a�bd���� S�I��ώ��y�)�;�|5�Y7�%X���yb�I<>K�u��k{\XQ��y*�
XV�����qM�a��H��y��C6�����n���9��м�y�Y����@�ӋiB$u��V��y��W��(�B�>[�U;7j���yJ�t�h��/�b�.(S��R��y��ܚJB -�CX�Z���k���yj/m�ء��N��{�@B2͓��yr	��E%j�i!��PB"�"�y��Q?Eh2x2�h-R=�Ə��y��=>��+T
�� ���
��y�#�gD5I`(!����j��yr�2f
tP�Jb�PD�ܧ�y������F�D�	.��q�I�8�y2+�!F�c���Q?�A���#�yb �u�V��(	F�J1��Ί��yb��G� I�V��9>��@v ��ya��U\����49�� &@��yr��-z�:�e`�1�I��X$�yiF�
�L�K��|l@S@^<�y¯X}���5`�r;8�˵C<�y�H%v\	��Jȼ?��"��_��y2o��K�("�N�2���q����y
� i3J͜o�n�䥆s����"O�lC�c÷/ ,���G>���F"O�U+��	��tb���$��"O�-� �A�d\���\k� �P"O�]��m˱9�iSȏ�h�:�"O����ڿC�Z��b�Ր9�R|Ѕ"O�X�H�}1�}ss喫.IP!#1"Oxhz&��M���eg]�'.���"O��#@�}Ԉ�f��Y��`@q"O��0�X G���7�W�	�؉
t"O��ψ<H��@L69,�u�T �O�=E�d�\�e����!WBRTk'`�*Ui!��`d�X�2j޾X%¡�a.ۢ�!�s�E
b�En��2���6!�Ğ=%���� "��]�b!)"!�� ��$F�m����`!�$U�b�r��+F&c�f��e��>i!���!d��0-!^���A��q�!��@:�I#�O6$�H�	��'�!�
$ĸ��pe�*��AX��=$�!��^�����&�U��ͻ2�	�=�!����8�;��C4p�C"O�xy��'� ``BU͊1��M��'�Ԁj�mH.󴘱 �Y�f@�	�'�r�6��*e���6kE�L:�'��qz0I�(IE�PV��~��ِ*OR�=E��F�=ot-�g��b��4�&@L:�?�����4��AV(Q�dy^�2���(��؅Ɠ>��@���<Hg��0��zP5)�O~��8�O$�)��/@��z

2�Ա��"O��.�5u�tPS*�
{xY�u"O�T1�a�yf|�QN.PUrЛT"O@˶!A�n+z`�tĄ%.����[�DD{��,5��!�̚�QO��S�/иd��Oȣ=��H�ö&�*�`RA�07Zi��"O��B�*#o����b�s`d�s��'�!�D��O9ށ��'I8��X�E҈vI!��b����Dc��)��p s�_$y�!�$���d�8 @ԃ�:�!�D�* �0�7HZ�|h
�$B�!E��'P���i��X���"
9��LarcP�i�!򤝭/a�IrVf�6�ށk �W!�$z����OP�E�^��$�P�k4!�D��&:AصHf�K�6#!�W��4�+W@�PH	��d۝�!�$Q47c����oޮ*����`��5T�!�� <�i�kӓ3y�0���( !��0q�L�t�:��,�r���=���â#��t�V	ӗX����5a�?z%,C䉴#
�򅋗/j� 9�QB�\RC�	<$��6�	���}R�� �=�B��(p�B� ƣU(jPV�xTbٻ(�C�$QD��a�
-�$PZ�Ř
' :C�	N� }���٬I�����6��=�Ǔ]�& ;���,��u���:>Y��,KPaR�b��0]�zE��0s�8�ȓ.��a�0�%��i���)O�R]�'7a~R(�a9�Y�K ��s��y��M�R��%�Y'Kg���%��y	�8&�؁�1��@�O��yBa�CA*<!b�3z� X��* �yBm�*T!(��f�B�F�( �ք]���xr�h���kf-��An�ܩ�KS%+�!�D�'eD��rB�+fJ4�q�.�B�'Ha~
� \`i!([57����Ձ~v
"OBۖ!�:��!ҍJ�g^(p�a"O���n�?L�5*V�I�N���4"O�+�g��2�B}K��_��C�"O-
��=4�P9j�'I zS�b��'*��R�̳&�ʚ#s��'��o:�O���d�%6�vU�C�Y�=��хb:
��f���Yu��4�ΈJ�L@7 ���G=D�dV�L�T��􇊏*�T���>D�xC�.����G��&�(��?D�(�ŁZ��v�@��&�(	D�!D��if#¾S��4qw���/��P��C%D�8�JT�1k�9@�\�6�x�3a�O(�O���>�3}��4(w^�A���n�,����yBD�=��t���f�(���ҩ�yR�Cc����ʛ�bM(�Q(�1�yR��w&u��K�0�v9k6��9�y�04&�!�Fs��u�M1�yk�hr��Y��9��$�婁��y�(��?�ZQ�	�'7�d�c���?A����c�@`�je�,s�D��Pm��&�$��	 $�d8�5Șm���T"��	\C�	 ejPp�Ҭi���2G�B�ɏS�45��)$v���B�9!�.C��K� R0O5j�:����$]&�C�IxW���W@��O�0�b!�	�[��C�ɞ6��XC�$�4 ���W��&�\C�ɽ}#t�j#Ԋ.�ȕ94 ���$�<�3_ ���`�~�^�C���gB���t�2��#.XE��˶o�Fd���h�D��B�?uh`dYS'I>�%�ȓVO�(+GK�	$- �i�N҃�օG��e-2�����#@��!��@��C��83���x�(��B�8�j&IG�IɄC�	�a�$	�v�)*��k��߁F����e��<�4A�mDDp�AM��[D@���5�$��MB!6����Rp���ƓsP���~���W��F��'�:���P�hZ��ڥ�,����'xa��5M��X��L�&Ur��@�F>���hOq�4�p	��V���ЀD �|����w"O������/�� �C�CZ���Ӧ"O��F�F5��ѫ���!!#x�`"O֙����2!w�C�(
�!A�'���O� ܖ�a��{A�T�E�-]62�' a~��ۆ<��#�X5YL�j0�N��䓏hOq�Z�K�jJc<��`��L��,���D8�S�)�9\1��Ĉ�N���F�\��r�'Y�De��)p� �3���U�x�c"O�·�O�rw�b���j9>�"O��C�EI&�@1�Y:F.�mJC�	���?A�$��k��Ȋ�B��i��K�<�yr��=��1ڀ��P�)����Pybg�c2e�W =^�H"��n�'�a��Id�A:Q�ʤa���,~W���'q( �'_!d��1��`I�>���Z "O�	�F��/c��r��ϑU��h�"OX���L�0m6�CvƝ�>����1�	|�O��DQ�B'J\4�S�	�I�V��	�'=�,��-7�xak�dʈ3��H�	�'C2�2�(Y1��̙7�P-1�l4r
�'�^a6�Y�]�G#��/Ht��	�'�J(A�_��1K'��1p88J�"O��H#'*�uS.�1v*T�@"O� ��2�V�2�dѸF�x�̱*U"Op�s/Z�b���:){����"O���E����fD�
"x�͂�"O��N��A�yf�<�r=�6"O��[�&O�K[4��0Z,<���Q�'d�kg)]�<j�1��ڀn@�;�d7D��R���偠�Y�q�8��r�*D�諃n��k�DBd��&( )*��4D��J�A�	'"Ne;U(T�+��%��4D�􀅠I#g���:5�רlo�Y¶2D�XY�מs�N�"�ɔ;.�iZ��*D��3"-��,�cU�sh29�Ҡ'D�l�db�k���H0?�M�#,3D�,�QlKm�j|�2�P�T�m�rJ1D�|r0G�I��˦)��t��X�Fa$D�|��������K-�x�IAk"D�lɂFH�M����K��<��m!D�$�c�\��H���n8:�d�1 !D�t���	�VA��&����H?D�lk!��B�Q�Չ��"����9D�� ��+������>����1D�X2�J]#�FӇ��4;6<��j1D���@�ߓ)�<��@Vvk6p�d�$D�p��)�UV ��,T?�`JG`8D�Hb�	�	G���W9D<���(D�l閮��C"�){5��I><4J�<D�Xr���Tnx=���Q�/UV��D�;D�d1���'wa���`4��0�8D�X���	&;����@4 ��Ր8D��b�]sd}҆�B6@�*Y@�2D����+S���SA����)��	.D��� 8p�>�����NG��"�+D����c�5\R��B�]>j��  �d+D��Z�¿5�F̺�[+|)�p�p .D���$۰	�zX�Y]oĠ���*D��	q\�'2�M�4���2e�<sp�=D���t��m� �F�_�8S^��5O D���GE��b�A�asw,t��+?D�hA��s�<��Pg@9N����*D�007�֫7�x�)���(}ҥh"%)D���ۥ/b)0ʀH��̢��%D��i�.A���q����\PFE$D���9`�J<�����3�-90$D�Pr���b��ґ�e�za�c�=D�Xz��ު?���{"% ol��0D�y#F�!�����ؑ`S����+D�[�mja�HU�a�0�P�re�B�	�+Fq;�"Õ�,�"d�?&�jB�ɹ?���G�7E=�2�и9�"B��?���#b��H�KT�B�	�|Q8!�4��F�N ��%/f�B�I4X�tU��NKdV���̻f>�B�I�E]�RG�p�Q�%�-DU�B�	jO���%&��n���kxB��m�5�r �uBր��K�6P��C�6F���m\�eR��`��$��"O6�@ҢΛH"�Z�g�Q���f"O��Х�ٯ-~|(
B��
K\�B�$/LO�������,ɑ�'�}v����"OLUp�ײR$��ŖPX~�F"O$�`�D4)�.��u���0I�5P�"O���H�Od}�b#��7;:��"O��W��m!ԅz!c��d�~�1�"O��R��\�D� ��*d|�d�D�'��� ����G>5~q�a�Fs\ŁW"O���!Rj�y��I�"*Z�И0"Oj��6,�2r��HI�)W���"O�	 ���l���[���_����"O����&�����;���c�0XC"OJ}`UJÆ܀���V�JD4�"O��;��� z��`��\'9�`"O�����,���B��]Ҳ��P"O��PEgPx����f�$��ѓ"O>���HҼlh�@�x��h�u"O���#M�6��Y�x�x�+T"O�`�@ޮ~���������"O6e����i~`CqD�D��hR"O`	��eD�L,2$�����H�D2"O*����֤��N6�}#�"Oj)��F������^~�m�r"O���b�4� ���F��BW"Obhdi�-��p;v��w6�P��"O0AZ��8S,�C��;c�2!�j��]���^�-nd0R��BV!��%FS�Q�cA�l���v��G!��$�|�S 
�a-�p;�쓨XJ!��şi_b�E��?'�	��mWO�!��?7�X
��ۭA�$��-�	R�!��E��U@ԂՌl���̆,i�!��%�x��FOZ�	Φغ��� !�Z�=>U3�h��`�HӅ@*!��
)$�D�7ij���p��g��}�(*�MD&LnX��g�I:!HxH�<D�xQ�,�0$��R�ŧa�x�k�l3ړ�0<�ƨ܅����Q	F����͚r�<9H+p�b]��d�:w9`���k�<���&�!��8X�u0���<�&���0}��g��>����b�<Q�E\&�(�FE�cm��3.X]�<�W� �:Bd��� �$}���*Ԍ�}�<�U�M/G��ɉ���r%T�j7'�A�<Y�Ł�{�m����T�\s�Zr�<�c������q�O�W>�a�D�S�<Y�(J>Vj�0��#|�`��L�<���H-Pk@�+E��=�h5�QXO�<�M_�>��D�%[
��I�<��ŝ�pլœQ�$B��fH�<��iV�LAE�W,�	K����h�]�<yv#^5�!е�"%�f�¯�W�<awOHY�D`e�Jy$ہ��Q�<Iv��"��A�-W�:���A�Q�<�%'��~�2�f��z�`a��@TJ�<��
G&h�Hy�6�ك9 FLz/�B�<���҃]���7�?��!z��A�<	��A� hX�R��9bB��)rO�e�<q���`�aa ��b ��u�c�<Qu���L�нP��ҕ(k���eLJ�<iRMB�Bi�� dW7E�d��I�<�w$�r�rG��,��b�&F�<�3C�~��J@�C?#�y��O�����'���Y*@�#�CԞ��D���y?�{���-dT8�J�"��e2R�4!�d##Z��#�5�H2È$!�d��(_2�Ƀ��>��*%�Ѥ;b!�d��Q���r�(�rو��ÔoT!�ۯ?�䵪0R%&�~��2"Oz�uiU#1�di����$Z���u�'K�2O*���B܂M�nqV�7���3��'��)� �%H�+��d����7��ɚU"O0�3EL j��X����2����r"O����v6%��S�1��"O���!�ۈ0�|�0��A +�\�"�"Oz)@�L��A�)C�FH�yt�1D"O�e�0�2cI8Ѹ!,��v1�G�'��i�eN�;tQj���A4hxV�/�O��W����@�=��T�w���Y����"�P����!?��÷�/�"m�ȓ.�LB *O?���u��UF�t�ȓG':y�a��h��D�����.��$ �-xS��B��)r��
�ՇȓF�x�c���o�ڀ��Ň�vhX�ȓ�
�c1���O�d�v�V4~`d��`�'�E
%�#+Ţ�P׶1@ �'h�2�AX�D�.��&L��y�B�)�'��`CU`����%����p�'=����ӟ+G4��	�r�UC�'��q���t��0��oR+l�ҝ��'��q���
Y.N��Ԭ�UC��b�'�xl9���z���"	��؁��'�����Z�"nv�Ps#���}���xb�ݚl�b���H9�2Y!U�H��yb��$���s�eמD����C��	�y�C�U�2��C�"5�v�3r��$�y�S71���s���em1��!���y"F�֌<;p�N�(	�rA���y�&Ыo�h���¦	�<x ؊��'^ў�O<䥺�͋9���&�>�L���'䶩��?]_�dy�OL� M����'>m2jT��NQ�&�'D�M9�'"� Sr-�O^jPu.�),��	�'i���Y\l�۱	Y�����'��!�C�'�Xy�O����'$�I���M<,0Di"!��2�|q��'O��ICR6$@8M!2��+�������'Vax�(wW�5("&�	Y.ٓ҆_�y���;!FP��l�+T�@��e��y����up4x���5JJi�R�[	�yҁ��p3F�L��fs"���y2� �8$!e		ɖ�kr ��yRI۲@� ��c�v���A���x2�՟E>�m�ye6���C��F��?��
���a�F=v��x�b$˝s�:ԅȓ3�R��a��=V��;�G�.C(�ȓf�($�+�l���'�C8��ȓ;�!!2�T�)A�p񎏙(2t���a��J�*Θg�M�钞R�TA�ȓ,�|�f@\�r�l�3ណ7]�xE���2*���A�M�.�:�2��P�"4�x�'�B�'��D�C�S?W��HׯB7<)�E��'�h�F�x��(r���e�l���'�T=P��݂*
P�n��X�Hj
�'��p�l��9�2Q� 芮~Rn��	�'��x &+�k�p�7w�&)	�'�p��VOV�S���E�%�03�'��y�1F�	�8��S�I	�Ll����$�5�5�c	�A�Z��^ǔ-�FT�l��ݟ���*�t��/ہ?���fꋦ/@,C�I�-�<��������1�o}�B��X(]�Ѥ��Zp �+FH.C�I�y�~��wOʡk�Θhŀ�6<"�B�I4Jm�DD�h�<��b�qA�C�P��`:�)��eYI7�A	~����:��t�� ���a���Q�J4P��Μ=E����|��'az"�EXa��:u��_�xQ#���=�D:O�Y�k�ch�2�*��ϐ��ƛ|R�'�az��H�:���O�T�eS��^��yC��-��
H�G}"M�*��y���8U�ɛ�iѶO���[��?��'������k.Z�4GAǪ<������O����p��\,4Ö�5�+R"C�	�?���j�f4�P�k�|�O��$�O����==�0�*0�к`ծ%	1O=.��O���M�Q� ��S�ygԭ�HE=wS!�D^=l���8[",��-�3Rh!�N-|@"&�(f�$U�p+�dE!����*[Ы\�mt1Su+�t��{�'��I G(�z�"
ߺhFiV�B�0B�	|�r�xE#�skތ� "y�.B�	2T���#�I�wD����[z�"�d#��C�Ġ��5A��Y*���B[R�[W� D��0s�(�� 4��/*.����=D����Q�Ud����M�6��}���:D��(�#ۄb�d�C�N��Au:�O��>3�hd�W�V ��C�E���x�ȓw�ӵ��U¬@��B��S1���ȓ\O�C`!�"��
��E� ��؆�6<�Cr
�`�0B�G�mT^�����}3�_�v䞁��Z��1��z�`�'�9h"��1���+K�L���v~BOL*r�����u��H�AͰ�y2�&'�֭���N�l��F�I��䓪?y�����c�F-��*�;d�t������yҩϴ;_(Z�[�b8B%��%�6�y2��Y��Qf��%p\�g&���y��ӸO!T�ጅS�I�\��y��B�UR�2�a#�D=��߬�hO���	�"
�L���3)�QFځ�!�d�=H�DdI-�&7x�I��_��!�0,���L�)�bܨ���XX!�D_8�y�����%����J!�$��\D2,�sh@;7�~�b��@��!����z9��z���Hă�"�!��iv�8*�=<�j�	C�Z��}���K�Ƕ-ˮY�2�4��Ũp$/D�X3B�%�F� ���W���Ħ1D�X��*��p��6T`G�/D�<�u	_�h�W�Vsf��a/(D�8X�h�c�~�Ɂ#U*=`�M$D�Dٲ.C�A��Z�钢|�P�ґ� D���&�;V.\��Ǔ5J�.�!
1|O.b����$�@�����T�,@r��-D�<��d�	Kp0H�l����H /<O�D#��2�x�Q��R�`�t�pK	�� C�ɎX��<���z4%����=yJB�/2�(���n��<ճ2�W��8B�I,*���2d�Ɗ=��8��.עP�8B�6Ir�k�o>�qI��ԑ/n0�=���?灋77Wz|[0��n��F+4�T�Ș;Cб���J.}�M`T��ɟ��'6��4����U���50TsA��7��ȓu�e@�A�!����C�܏\t����Iߊ�
��A���� G�S"6�م�
I��*�.� kp+�����H �@*eDN��}ic�S�5M�`��g�V�Ƞ��r�x�8lԇ�*}��NԈ��
/(0�(� �'
NfP���� | �#��*dD�5+˞�w�d�P�"OJ`b�FD���|���A�\)·"O��J�ѿh��Q�U�;�&���"O.�B���'G�@���� =�ʩ�"O�{W+X㒜��J�O��a�D"O��G�<��R1�M�l� �r�"O�q���Hc�%��@-�c�'�!�D]�1岉8�c�(� 1G��!�DUpyN �c͘�m��E��f�6�!�d�.R<�� �n�L��1:@i!�P� "v�qU��+�ȉ�ƪK�Sf!�Bb���A"�̡_�-0��Й>�!��=u�[�-�K͜,���)w!�DБ:g�!�g���y����@��s?!�$�B"���%�_�|�����	tD!򄋦 d���g%�1.���r �׃�!�-�5�p�O�N\�ҫW"R!��A�.I�I�>*p�|��I��!��6,d�bg�(\����ȃ:O!��ܽK�ژx1ぅ!W���4���b�!�\*n1���_�&��̘ �V- !�V<\�،ك�M�0�Le�wa�=~�!��' .���&F)f��qh+�A�!�$�?dbt�A�ε1��U;�HV�jr!�M?U�<Zs���W1(�`�V%@�!�[u�����#�-$.��4h�7d�!��^��Q9eρ�jb���K!�$�7�^p��eߣ7���hH#&!�ƫ�2��D�K��F��q��V!��ޮ7���jтS����GA�_!��%?j9�tOB��P!�F �%�!�䋜HR�ᙳ�ի��U�wMI�F�!� 1	�a���7v��)�ꑔ`!�䏁a��]��  "a�eB��)s!�d�\�x�D-NeK��9�ʈ[�'-���5/!��uт�T�'��L�
�'�<������j��Q���!?�8*
�'�L�8laD�8+X7/��
�'�b�"!mH�~�!�ӣHaډ��'�4@󀦙)^W�����A�740h�'��� �� uCt���� )'����'FB��խD���A%D�Q��a�'c�$ಪ_�?o XCO�!T�����'�������9�v8�W�P��D��'�V q7[~��uDhV��rAa	�'۔���2j0x���V�w�8*	�'{���/�}p�1j�jU8vg����'��2�e�/C��� ��=�:�'� h���Z?v-d�cI��<wc	�'s��5������IШU�2����'�툧-E�h޶�CgIR-3�`�	�'�j@҂�ǫ4֖d�֏C#2dq�'���0� �+F�B�9�"J�.�L���'A^���/��w��	�0%B<4�j]0	�'�,��r���vI�X��H�A�>�Z�'6�$pu 4c�����ʓ�2k�(��']�
��ϐ\������[^�D]H�'FV�H��-Fc�Y	s�Y�;�l���_��xBvLT�����%D�1��K-hD�B)�g̦�`qb@�:�N���#MRl�"�+@s)��qoe�ȓ�FYpe� :9
��#�ͻJ�	�ȓd{H|�$bE*��C���3ˊ8�ȓW�l=r�EMd1X1��.4�����S�? �-��7�U(�M*W�|��"O&]� h�*o%Z���W�T�&@�`"O4�����}NL�ң/ 91��	�"O��d"�$��-�O�f��S�"Oȵ��� JIy�@:{�.q��"O�Ըl��I
f���d�O�>a�@"O���f;�:Y�'�Z-� ��"O�UB�n�ހ���Ïk�4��"Ox���j�����)�8L�<��5"O��סs	�����P
Dp�"O������p����(!�He� "Ox��CR5~�r�GĲj}`�
s"O`h�Wd�Yh�BC�6MtTyc"Ob��"��)F��	A�ֳj�|�"O�	� K$���CG�
���a?D�(C�Gҗ v��h 僑t0^�ؗ�/D�,��rX�V�)%��X���.D�0p6/�>EL�5�F�Zh&pn,D�8��K�jh�T�� >!)��(D�d�C�	�!���CD�Z��|��*1D���J"���spȃA�X5{k.D���w�I�lPgMA�ErPq	�+D�@rP�4+$��СjRw�<	Y&D��C�J2� ��·^)��a$D��D�5��|[����X�=Z�h D�T��~��\�ҩ���"J D��CF� &`������ͅ+r��B�>D�DA�,��P�f��ƈU s��h�1G;D�x�Ї�eV��fǔ�{A����h6D���VeB�.d�p��oѶ6a�P��4D��3#����� �N	OВ+3D�@�aĒ/}��;��o$�Ya�k0D��w̝.@����)���YzD2D�H����
I��&��0 �pc�3D�T��*S��T�hRBQ�v�"��1D��:R�
�e��P5M#�y[��5D�4�w� �5��q!�Y�z3�ժ6�/D�xqq$��}:}���UBR��xCK)D��P4�%�x�D��T4��
(D��؁��b�y!pLўYUV���+D����IKd����1B�PX�p�)D����=v-�c�/S
l�.��C�'D�H`g�)�`�p0F ��Q���8D��Q%�S/s��X���7p~��Vf6D�Xa��	N!fD�o	1`x!�2D��T�M�:�f�F�>NI�0�>D������!��fL@R�8�R�"=D����
?H>!�t˜�;W(-�!��y�`�H�k	�V��)b��¦]�!��,Ch-b���=2���N�	Z!�$'i5���>��p ɢp=!���)e6d�5H�T %��͏p!�dGzJh)G���kըy��ٕ3t!�Ă+"���r�v�k�+��]W!�D0� 51��c�N��ūY�U�!�D��ga��pH��}�,�w�Y!J+!�����4��/;�dQ`e�KZ!!�d�C �r�����q;%�Y�:�!���?F��D��$-�,����.:�!�]�X��X�b"�u��ih���l�!򤗋E��}B�fA�6�&���͋�=g!�d�T�Jl�f��-p��AU!�9Y�l��A�-I�2�#B�[� !�DR	Y'���C���p�3�h`�!�� ���D�5=����H� [����"On�RVJɆ1U���Q�0ipV"Oީ��#�41f����G%9 H"O�=�u�WIL��
pk�:�!÷"O�(���ѭ)Nʇ�<"��e"O&��[�&�R�c`ɉ/I*��"OtM����b�R��B�\���"O�T)r�0}���R�ȽD��Y��"OP"7&�%[���\���Ze"O�+��O�G��RbD�\,B"O�,`w���Bs.�A��M�#7ji)"OI��,(W�Ζh 2� "O����h��Y�\�+��Ѹn^��r"O8l�#�J��-�$�I�;�e��"O��y�)��4�����EU��t�1V"O���P$X+|�RU�: �����"O��Y�e'6:h`�O��ih<�W"O8��	܉]�����4�qU"O�C���!��!si�s���)�"O�u����].�j�NP�l�R�+�"OTɳQ�B 2���J�� /,��� "Oz���@  ��S&�̰n��`e"Or�0VB�k8�)i[)$�$R�"O�����vՎArFm�H Pل"O�ek����SV�r��Y�A.��d"O A��o <uAV-�QC�; ^ݫu"O6AgɣS��]S�"@�st@��"O����#+���5��L��l��"O�����I�~��!ͽm���[�"OX�:�B�0���
D1K{�<I"Oz�I��)�@pؖ�Gg��×"O\m�Gɋ�d}�M@�iش_��a�"O�e
֡�D��Aݒ�i0"O*�����\DN���@���``�"O��
 *I(@UAF-Q37�٪c"O��	�Κ� ��A�K,q�c�"OZ2%�j$�8p�ҍyʀ
a"O�`�#ʛ: �k�C�"K�u:�"O:1��g�@��l���w"O&���i82����Y	r|
�k�"OR-a+Ik������P��-s�"Od�9S�����#%!M�Ф$p"O���t�W)Sgt��Ņ�VE�v"O��z�)�~�ĉP%�R�`�Q�"O�P�# �Kf6�;�K\"�����"O����,I(��Q���@t���"O����'1d}�枓3�*ͯ�yȒ;aL�Xg��"�#����y��]����4!���,��RLQ=�yB�\/>UZ�(��Z3% A�ں�y�]�Ya5n	��z\��%�y���!nx�(e��)n
z��SIʒ�y�C�T(6���ũc����B� T"�E+BFbi�&,�=5ԐB�I�_pE)���m�V����z�B�1y��Ѓ	XcV9�U@�QN�B�ɞ(r,3	H5;(�����A�#pB�y��	R'K[�Y���02#�'p`B�I~�~����Nl�p�Mڱt�C�I�D#�D�3n�35�H�;@QC��:ڌ{C����T�W,Öe�B�kZ\%3�,7LQ�x�OA=�zC�:�N샔�L(���x�D�.	C�I�پy�󩈢@�fT���
'��B�)� ���Be��t&��"�<:v���"O���`�%>���� C��0�V�$"O��R,�hab`��s�����"O�u�,7J}bB#/�PZ�"O����lC0H^�p��S��$�c"O��Z�]�v(�Tr6n	� .鉣"O:��,X�1
��ˆ�Q:q�Xa"O��g���a��mQ.���"OhA���8���A�f�<?����"O~��w#�Kĉ��Yf�H�;�"O����Ɨ�V����`U)J-q�2"O�D(�%[�1�BԪ�	Tf=Zv"OT��e�/XR��������"Oh�Baۑ ���aQS8V�P�"O4�;�Bd���1HF���:�"OB�K�G�y�ɦL1=����`"O0�V�̟Ps���3�Y�x�4�J�"O�,��@۶P)ؼc�C��x"O��9�ɒ������ƈ�W.\E��"O��%/$3�@��Z�BL���!��7c_�0��E|H�� �6;�!�Q�~������K8,��/A4�!򄄭
v���/͢h RUʴmR�&�!�䞡n��-b����4B�+ޡW�!�d�<��c*V<f�@tkcm��n�!�$P;$
r	PΔ���s4l�	s!�DӺAQ�yH!�^�l��9aR���M!�dY�C\�ƈ
&l�ڠ �-�-J!��6_�@�iC?��I$l�*O!�4��AjћI��D��	<?!�âZp���$�ë$^L�g��+d�!�DO�:3J�q��I�jX�kL!�D�X(��hb��_�(�;���'$D!�D�J�`���鈔m�PC$Lэ>!��I6h�xd!L!?�m� �!j!���l\Vg�>*)�E�B
�>!����֍�Q���J7��n�!�ĆX;(��Bq�h ("�ՙr3!�B�6ذ����Ż/��I���/!�Hm�4�#ũY�g.�e��T�vC!�$O�R|@���:�]�B��Y�!�D�>?��,[R��0J��I�%fr!򤒺2��p�V,bd�ڗIH+`9!�[(Hرs$��`��$B.�"z!��"��={��^�B���!d�I�!�ܟL���aT��"�n�) ��30o!�dǎ]0��F׬7��a�ˑ.�!�D��-�p�8)p��p��ˍy�!�D��G�����55V��r�NO�(�!��15{��*GK�%2�� �M�N�!�%z�A۱��j�j��cC�{�!��@�
��'O�CT�X7bR�{;!��W������ړl�f��/�K*!�$��tƠ]����}Ş��mI�1�!�ĆoU��;1�@�B�����8�!�=m��8�;,����e�ə�!��^��1Z�+�UQL�"�'0�!�dP:mU����,J��\x��)w>!��	�H,@b,D&"6�5�!�ŖR��e��K�Y� �w�+	�!�D�nz`�0c���fQ�t��q�!�DʱTɶh��G�I���a��>?�!�$Z�CG�HCF�F� -��!�,�!�OW94�z�%ׄ o6|�B6X�!�� Z	��[�A*�D�&�6I�G"OE �k�m�"t�&TnC���"O.5#'�^.�X���* <2F"O� Z�����:�-�ruxR"Oj�mֲt�N�!��$1_zy��"O�]�ҡR.1��K$	BLLH"O�`�U/eƐ����I�1Y&,x4"O���c͊<Vz�e�[�^p�h��"O�8ڂ@L���	�,�2F9�"OJ�r#�XY������kblC�"O���I4J�X��0��C��XR�"O���ۨ?BUK6�8j~`9t"O� `�Ό}�pȉ�dK
ov�pa"O(0PvdK[!����L&*/��A"Ov����މ35��!�a �% j��"O�ɭ�^�,;pM�e	�S$�s�<aU�T9;8��*�!� _xh��� h�<Ɇ��
B\Рdc�������d�<1S& 
g�*�)2�7v��p��/�k�<���%|�l��t��5m��6�\�<�	,H��s��ʻEF�u�__�<��n�d�2@�;_�͐B�X�<��[x�(�ԎU�I�q���H�<�g��=M�P��JP���T�D�<a�*:HÐ��j�<� 4�O�j�<A��5Z�D}�"�{����Q)Tq�<	�%B�A,���dJ֍"�#!��F�<y	J�
�^��WM2�ԙ[2@�<٦ϋ���9QYq��U"q�Ch�!��[�T�k���<h�v�pIi�'v$p%�*$����#�L�&��'��x�O	�)L6�CQBюC��Mj�'*�E9j��3q����  9=�!k	�'��8Ј�3GPn}���_:���'V
��䉜s[�m���۫&��t�
�''��ف�Ϯ:K���l�da�'���a�2;������>��q�'�
���݈	3R��7����*Y*�'M��x�j��U�)p�����4��'���r$���,�c���
j4�@��') ���L�_X�p�$gʐK#�e*�'f6 ���GI��r�Õo����'�"�:%�(x�}�B��<k�āS
�'7�<ӳ'�;GDR�����M�Zm�	�'�z����D@hXs�	M?�<�Q�'�F�ȳ�Ł^��Ȕ#�k�A��'�p̫g�AJX���S_r�QA�'�M�B�	pe,@���W��J���'�nH�/+4�@q�����)��'��K�l�Ԅ�sJv����+U����	<3�uq#�671��5��+'��C�I�C��9B���YG����a�+&�D{�����h�e"�E��q��dJ-]�N��Fe9D�H�7JfQ�X�)M�4"m�T%6D�D��S没q�N� `
1��2D�� Ӌ5����z��2�a<D�҃�#�$�Is/9oh���%D�0���T*cjh�S	��N9@wa�<��M��K�'CW��={S��)-��̇��w~��^�~)z��c��d�pZ�$��y��;T=�xA�lȌe0�A�'��')�z��F#sOn�jÑT�6l�b�P&�Pxҷi����4�S�$�RD�D�O��y��'ў�S���'�`I�
�4\��Q�I�҈�8OPHEz
� �rq��%��!��ԯyIZ,���;?	�]_Mɳ��.1V	Z7d�?V�`��Ƀ��'A@��R�
|
ջ��
�i)�'�@uy�L�E�ش0�(F2��I>�q-f���O�L��t�S�Z����¡�~��,K Ob,�@�$�̙�So;C��RT��7����#RGVR�N���h�
� C�!�ߑ*�L	C-S�(�t�@D�0�P��ȓ�T�S�	Y)���� g����'�)�� A%�Bm�2�J&E�;��}p�/D���O�5$�K�@B�!��1Ԅ�����I4B��a�O����4kE�l�B�I2NW��&�M�@�viH"(�!d�B�I73�8j�f�+P.���D9W3dC�Z�k1���,����Ɗ1R�B�	$y!\���*�1��_>5�C�ɩ}+��6B��(K��v�4C�I�r��ęeE��z)̸ۇM�2�B�	..R c�cY�S�ke�[�6'B�ɧ�"h��Fʬ$�T�Rc�D%B�I~�*���4g�� IɺV��C��1� ��oկJ���y�%L911$B䉫5FMc#w�8��6\�B��~�m�w.˽Z�t谀�݆������p<��(I3���)�FB���["
�Y���'�h�* #�<2�)p��@�'���7斌k/�"Pǚ)Wd�#�'v����N�-zM��o�#\LX�'�lXP&�Ie��aw��YO�!��''v,�v��R�q&�M &b�
�'V,�����^�B�{��.�p��	�'\B��g�W3D��I�&����'�A� �Q�(9�i�H��mA�'=T�9'	��L���C��
�p��	�'�S��*CTz�&��1����'6��Wi�4K.hH��h�8��Q��'4
�;��}UX�	&6�H����C�zPvikT�@\F9�3e%Gd�V�)���1�z�4��ڱJ���1�.�*�O0kC,�.3г�a�)3 ��(A�'8�N-$�	83J	>W�+��V� �ȓ.��%�(ڼz��Mb4���Iv�'��x���1 �XBĢ�-y״����&D�����+I���0.�t�tT2� &}��)��%Ӱ�a�[Pdb�L{�U����s�Hണפ5��l�p�D�������5D��:����6Y���A�NFn ��4D��ɇ��!��h!J��^�(��0D��9�d�U�(��E�d�͙ �-D��� �Գ\��g�,+��c3?��Q��ħk�)��LQe.����M�1�Ňȓΰ�s��6���APD��B��@�<I�
��b��SQ�R�B��ܓ��<)ܴ1��XGY�S�RQ'K^�B�.����>a���	_ކH�� �j�� ����B�#?�M<!J|R񄙞
^l�h�IMK����y����-mGX5ƦZ!L�h`�v�Tцȓ`����6���!ɉ�%�*�FzB�'p1KA��9�Pa�`JB�+�Բ�O�=E��ꄯm��;��@�%��! ����M�'i���v�Bt��h���w�@��'�(p��&W�Pk �@'�
�k� J��hO�ܨ�Zy�乹�K	T$��B"O����ܠeWH|���Vڌ:�"O� 2U+���0A��R㕰X%:%�P�D{����?�Fm8�:,;8�a��8V���)��]��#oF U&G%M..̑W@>��#��U�'7�T�D=v����S?	n�t�O���dУ#�Q!d�$��sfb�s��yB��>���P��1����q�sā	y B�	%��9����"�2�ȧH�,��C�W�^}kƬi74���ޔBYC䉛k���QC	�h��p۰B��J�C�	'	�3�,	�{��I5N�7m^�Fy��s>�k5�	�E��y�$P�~�Qo��d� C�I�Z���v+�`�����+\t�b� G{��df�.+�4sQ+ƃ�hl����=	q����I> ���z���iI�l0 �%)΄b��@�'/�d��B.W��BDL4������?qI>QgD�<,=��Z�f^�y����2��x� H�O�p�$ϾjY>m�!�����O�˓ɸO����ĭ�O�B�x�,�ŐA����x�fGqY�=����`,��T-����')�	!�$�#l����m�7
:8�B՞BN!�G �h�`�<h\lD���0�1O�l�)��?T�Xl
�N.�$2��&�C�ɱl��y*���73����G��*s�C�[�&�q��"n�(�ֆP� SxC䉣R`,UƉG�Uh%�A�{ph��6�O��Bl�M3��I%2�#�~�����>�4�j��b!�=(�F��Gx³i�a�ā��Q���36J�4	i詁fJ���yR�Ƥ#j�0��K�
BFqi�M0�y*��	�\Ŕ'n�UYQa8�y�V#��A;�e�>T�`�[Q�.��UX�� ꌵ$+�u����$D �f>D��q��ΞE{�X�g�6=��� �+0?1C�	H�'�X1#B!ؒX���ydB��TG���}��|�~�0U�`y�a
�xFM�$��y��h#��t���O������E�̍��$�7{��ˈR�xR�UR�,��B��o�̸�VBђp�H�$�鉇{HF ��Z�?��T*"hXDc�x�'��>�ɴQ�N�&'������+�xC��,U�dN98��w��2ml#<�ϓ)[����@�� roW��(��%�����#ϳ`9�!P��pc��'��}"dI3F�`�v��P(�@�7o8�yBĊ:4j� ��HQ B.��)�̌$��'�a{��#U����Fg߮8��ʕ∪�y���#`PS �5��\YI���y��	gE|�ŉ�	1-�DyG����y���6=����3#,!�Ԕ�V�٣�y2�JI�D:�"P!J�r�6�yBN�p�4jG���q�ï�y�E�YZ=+���%_wP�#��\��yrCƠ�r��ʔ<z~h*�5�y�X7)�蠺���x��8�
&�y��߄N؉�T+����l�d,1�y��ޔ�����ʏ�	��$`�����y2��5�4���1��mÈ��yr];R���J'�!?��8bI��y2�R�[��`���d��@Q���yR�ؘ^Fj`/�
^"6P�0`ʭ�y�&�P�s� H1g�F���n���y��	6t��b� g�� G(K!�y���"��Y���`�iٖ!�y���!^ÀM `�4ҩ���T�y�B��H�����	53+���a$�y
� V�"�kI�h�P  ��1��h�"O��
s��f("����Z:���Q"O����j�~i	���<zs1"O�D1t��-j}�%��BV�V>���"Od	�aE�4��p��a�*F�Z"O��`��N'��T����R��"O�\���ܗ��'�6:�m��Qp�<�t*ѯB�!1�/�Iy@@l�<i��A4ቒ
�S���Pt�]B�<�Q/��l�Jݡ`-oDVD(��Pt�<�e�Z-f6H
Ň�L.aۣ
�l�<�!��'��`��M�H���{�l	e�<�2@I�S�H�{'��bDxxKc+�c�<�c� ��ܹtj�5Y����I�b�<٥���w�r!('"��6��xIbL�^�<�P�T�_�B;�D�+��i�I]�<�6�A��	"�
�PYlh�th�t�<)vKZ�l�59S��r�x�[ %�x�<��e])o��HV�_
�vG
t�<A�
��S�X�3���CF�<)7�;Y�Ee�K2BJ$d���_m�<��J=I�vm��$4 ` 
g�<�!��u�(t	��5c8��Ki�<��6P���!Ʀ1Z@�	��n�6U^�q�C-��]{5�#|P�<ђG��Zh�� �[�pH�ˊp�<����/n4l��,O$h"�#ŀo�<YG���|	��<�\Y�#�j�<󊉑��(w�R��P`���j�<���O"\��J�~� ��`�<y� M[�x�9G�m^.�PS[�<)�a�<RdWR�m�h%A�b](x!���w��\k�CE<%���`���9!�Dz���#pk�7�F�!F���<9!�DT�T�Y�F��v�F�í^!�B�PD��/Y�o4x�uJ�`�!���+L	҃��P���	AD�!�D(��l(rO��v�Hr��Ƀ�!�d ι��l�(�I�Q�t�!�d�I/`\Cٌ�� �"�!��3$���eF���%�"6Q�!��Y�=N���NG�*�֘�Z+O!�du^���F��7v�)���B>!���#1�DX��R�p\���c̘x�!��%3,p�V��a.���!W$-�!�ŮZR6�8�Bɧ:*:�;���h�!�D��+rب,4� ��a�|B��u"Oj8�W� >�TѲ�!Ctu�7"O�)��A̩XN����G�'G(|�I�"OҼ���3Z&��gU���:�"Oz���R�� �Ӽ���"O��0G��$L������s�z�
�"O��)�b�3S.�#��F7��`�"O\y5�D�2Et� �z�D@�7"O�92ah�/s� ���Q���q��"Or\a*[	��U`����:TQ�"O�IА��xI[�Բ{�0:&"O�چ��LLڀ���"@�:��"O	x�C��H�8�J�U�ıb�"Of]�TD�0�������xxLDj#"O�(0���b�b��!hR��"O�8��D1��тe�/0���6"O�5#�E�5�Ƒ�e���*r�"O�"��B~0*�3hC����'�NX�c��cUX�� b�"��	��� @@Y��Ҩ���{v��_�H�x�"O�<0�I�I�2��Ц�}� �8�"O�1z!�ý0�=���8}�ZT��"O�u��G�	(y�'���B�"O���EY�$[:i3fD�!���"O��E�,c����Ԙ2섙r�"O���8�4�B"�|�*!:e"Op1R�C�h��"& X�I��(;�"O"���Mڕ4��IX���p��"�"O� ��G� 6�N�zFnu�Jd��"O���#��)A�	ꕊw��zU"Oxk`͊0%7V�8�I�wi��s"O�A����2	ʤ�`H
tl�8��"O��J�B�y�`�(fE��J�QZ�"O�,pƏ�?T�a�@��*v�>Q{�"O̴��㒴v<T�"W.�A���"O!��@�`��պpdY�:���"O\t�v.�C�h8����#;N�c�"On��ը��P���mٲ)�[�"O*��iR�lr؝��,X�b�i�@"O��iƄ�8L�FU����?l�1�"O2��4ɒ�`�hq�Ձ� ű3"On�3��T�5;< �F��$�n�6"OpAZc�X�h� �v��$��g"O�=�#��,t*J��VL46�N��0"O6��C�7y6E���B99y���"Ot� I,�D�$�Մ�Z��@"O��"�AJ�"��Yn��)J�S"O=��aЉ5�`)�-FPݺ�"O*�V��o�ѓ�)7��a�"O�XR�C(W�V�B�h��8L%I"O0��f�:i�g�;M����"O~�0��cX*0I�:¢��Q�O,�r��2�?6�N�s=���O X�� ݘ� �H�^���i�Dp ຕOͻ�?��� Z��`�Gl�;(��Ղ�$f�e�/���Y���d]�U�u Nض0ƈ^�&X����P�I�����J�5�H�:�KGV�2��h ��jb��֥��%uh)sH΋�a|�,4f�:Щ�2HZ��C<�����#� ���'>�{�hLp�(L��x�I�5��d���X_��q����W�VB�,���YĩQ�+�m �o� p���ĝF�%ڒΛ ��!b'�����'�O���0Ro�<<��HJu嚺|,kߓUR����aA0u��6R�~�yON=N:��#l��O�4%�7�Z���N�ܣ|�'h���SA!4�6��n��v�<�a���Z&9��p�QH�O���Ruc�3U�CV "y�����IH�V=�3���1�0>YVԔ6p�9Q
�=9���ˍ�g�Pe9�M�����*����N/5�� 5��n�	/�4��1&N!�$J�9����	
S4tI4�ֱz��g@�"o䀐`C�E�b���
�8��ħt���[�!��W�b蠄"uBԅ�I%�;���0�5�PK�:TYE�4�D �k�X�U���|�+/�g}��J��=Qm׳Ϫآ�$V�(O`=������*Kf��jݵx���'1L�k技����qa�O�Ik2��=�>I!ٝ�^Ir�&U����e�B�'��8�LNE��>�@�*��{`�Ҽ1�h�	�"O8d�p)ӡp�nzT/N1^��xH&���>2G-��F���8�>T�d��w�X�mסH�HA(YW��X��'���yA�[�
}C�ʎ.@���޴<m(tR�[#j�L��%X��	�X�U�=��ȅ8>a2 ҕ��,mۮ]��V8�d�)��T08ZA�;��M�⣕�1�$��a��t��D�qEA�6�0=A�CFt! !L�w�� ���R�'ZT<�nBA~)�'��8�%��@�0�Y �ŵq$pe�e&���J���A�<A���5Av��2�2#��$����*$�"AC��(vV5#��'/F�R�6Dq���}��1a|5�o�>�F�C!�);\C�ɘ!1h}�&�A���c�i�v���	BcV�Fff�y��:s�
�q��|
��D��c�P�nAd�����F�ּ�qM:�O�s�nG7o�c� �'�
+�P���
ßRk�tIG.Ο��IԌ~�$���'�L�f�Ԝ=u©���"�D���D�U��<K�*8�҃��}�B�0JL0F�V�B<)(���A� �E��M�ȓly��Cg��Y��0�"��4���!>sRy��a��q)Rj�o~��'�t�'B�l�����/e<E�O���/g8M�@��(�T �A6<�`xC!�ZX��%�R�K�c�r��W,�7F�1��� (Ϭ�Vmg���,|��<H�CC�)#�M�!�>���k�ȝf80��OH���:�p|`cń�+� �I�M�C�L�bv��BlU���P�Ж'[h�0��O�L��<Y��;UQ�TZ"��?0ՀL��C!eD�cee�$2.�3#�H�I:��	?WR�\JCR���OBL�"ėIo�۴�E��}�4�'].��.R81e���'@l�@1g@,~	��&��2N ��sOJq��i�,=	f���Y��'��F�	p̓?92��tF�'F�l��4#�dҴȦO��B��G	%ļA��gg�4�1�)�<Y�$�hA�Y5(��Ԩ�璲��-I��:����'���TX:5��O�Y��m��C���g��&����6~ٌ�8���Jw��Ǔ^�E�'��D���$g0x2%�e!5z���ZwH�:��c�`B9+�<��"n���rH.l��D�BϦ� 	rF���ht��K�@&�TZA�Ѡa�|�&�j��`y�bϦ�:�[�P�EBJ�]���GCWB%Qu)^�p<c�<tY�դyG܄�2��
���j�:;25����Y�����a��(����C�R I"��u��@)Ŭ̜�\:�W�BA��\�f�zDӢA܎_��R�A�"J��*�ԌC�7C����lkP,��Q�S�D�8\j3�I8]�N�5d\�v���f��'n�	a`D�XD�q�lb�*B&@�H�D\G�'Ɛ�Mި1��M�SC� ��m�3���P��2j]�89L{��59Ô�3E�)3��I�S���m�Ì��Wo�Y��O+A?�U��$߾{i��HS&<��2��'y�Ճ���W���x���A�8A�UkX?=(�7��ʡ���%M�~%�w'�7m�Ɓ�ah��O��QΓ{r\����;�>IBꁤe��0�C2�O�5pb��J	�Q�SD��`1��3�gI�m�d 	�/�,}M:!2fC]>2v�$�&
�v���4O���G)�S8@BX$�p@�]�]�G+ޢn�ޣ<�j9CEH �� �Z�I�k�b���՜\�h���C�dV�`�D�pDH���5O<�x��$APaO?���5/T��L��
a��Ô�R�yisb��;�RQ��O�'X?H�F�D�Ǩ^:����fV�se�H��IB:�0:Ef��H`rk�����>��!�v�py�嘘P�6����9�`aW�ǑdQ��Q�钫/�Q�;<Y�A�!�ٕdoZm��ʫ���"���Ra^�$����K�u�j���T�Z�0���
�SN�u���9V$���mA�*��Qu(�5Tp^��C%¯]�t���AT��I���O�n���A��R�ƨG<m�d�r��RWkH�0E!�e'��"�l�z�*˧(X$m��F���z4��!���͚�e2�G�b#|�'�L�h�%�5P{R�+"�G�À0��
Z�Ī;$�!�cc�bE���9��h�>|�*@
`�*���"O,]��G?^G~�M�J�L����
^p��%$�%
�$ʴ�O��)'�b� ;B�F���uz�j�9Y"Q��#Uh��
����K���.ؠ)kT����V�����& Ux��(�
ԷN�qx�4�Pv�7�d�r��
U�H�Y8uN5�P(�E�FA0G���v@ĥQkTŇȓNmDU"2�ڜN��d���;{4T����% ��ѹT�L�2��wEl��?�$W�E�� ْHv�1�R�k�<�@�S��-����B��t�F"L%'>�D�}���h���l"�D��HO 5X�+ֿw���r#L'��ap&�')H�۠�!�p%a'%���-�aǒX"%���ғtV�ԛ��'o����W��U��3ي((�����.9bԑV@�8xnQ!I|2eE��[����A.Z��8�6D[G�<	�T�jT5�c@7������B}?)����iU�'}����!~�8�
ï�6P�R�p7@ԩu�!��'N�Au�ŋH���0�M'��'�ċ �YX���#L4�P�C�8Y8���I7D�,���Л��X(�C�T8ā5a(D��p�ˊ��݀��B�QUHI��(D� !4�_�,��@3�;>y�1+4�+D���H7�1��o��S ��(p�(D�(r��� �0�2��>.�24�v
$D�p� k����|�B�0!c2�Qq�7D�\� ˛!T>�#�N�H#PAX�?D�\BV�ZQ@�
p�C�A\��� h;D�t�0�ٿDQ�ֆ%0�zt
��-D�<���\;A�j���<	����k*D�p��W75bܢ6�`��G)D�b7EY���O��|�:6�O�<� 2���f�O'� "�ӆ8$ �"OzH2����D���OU�] 1b"O�T��e��>�t���Hا�,��"O����+p�x��2���p)"O<q��E?�j5�Ek�k�޵S�"OŻň��ىF
ōz��Aː"O(=X%拦0|�k�%2�(�8�"O$���N�d����Aj���ҹ:""O���'�%.����`D�vl�<�F"OR�c!Ö��hWj�,lC�h�"O����lA�������\�8p2"O�- ���<D
[QҁR�n�q"Oj<�Kӓ=���ag	��(<H1"O&+Yv�)E7�pQ�"O�QT�Z� �68R�J�Gr4Ћ�"Oа*�� �ePl�d�)2f\�3"O�,ZS�����+�'52��Kv"O:\+'nǰq�ٛ��ՐM;���P"O�i Vg�p7�)�c�)K�	�"O�1��*N%U/���ɷH��e;�"O�dc�(B�%�*����Etوy��"OMr�/��h��	G�2��+"O"��Ӄ�"��`�'6�Ч"O�b����$d;u��5/����"O�� �DU�i�~�W׫J𱹧"O�y�n�L.,�"�AƨK��$�p"O�q���C<6���%��?v�s@"OR$����bhp���Pd�j0"O UKQ�%�VIQ�kO���2"O��JQ�U�
n� 22�������"O*��4��,x@�)�-�b�J�5"O�5P�
�-��8a������2�"Oz���+K�0��B�z�yG"OJ��1kٿ/�XL�Qj� A�ɘV"O@�y��׷|k��qWB��u`�"OB�z���}d����*��T٦$��"OrЖʚ�c�*IB���D�"��c"O@$�䍺-3V�ʱ(E,'֔!�"O�52G�1(˔阠h�<?+����"O���d�L�_m�)!P@� 9��	v"O(i�*R*'4h��f�,!�xZ "O�X!�U�i�ءpV$ݫ~a4j�"OLu� �F�A" ���T�0PJ���"O� @�͘���8�@�"�4a!"O������z=d��dR-9��Ȑ�"O��ʴCҧFΆ�EW-@ �"O�Đ�N>J��S�e\�^�$	�"O����8!%J��iP)>޹�d"O�u�Q�q:�-�H��*r�'"Op�Re@��|�����t��T��"O��˔�2:����4[�� ��"O�l5�]�q�z� 1��2���S"O.�����	HD�!0R`�3s+�p��"O�$⑈>�Z�P� �#)�ɠS"O�� �Ɔ&������<o�R"O�DJ�ٱ?#@�R�G����"OB�[�X92 t(UV:M�����"O��(T%2��d�3Bɔ|A$"O��"F��B�ֹ�qH@9).:!�"O�<Сk��p]<�3�
�
���"Op`v�@��p,k���*;�D��"O ��ԍ>(��)h�(�"B0D�"O,���j0M���Ш�%D�ʰ"O��σ2 uID��E/~ŀ�"O� p-�a�5F8:p&@�`��6"O@�؄CV]�� "��&eX��R"OJ�5�O%]̚L2�U-_n���"O��A3C�ti��]%L��"O�\���D�
���GG%���P�"O���F+ξ~�����x�  r"Oح�`�+��BUR�����"O8�)+���aK��Pk�"O�`6�^%��T�0�^084"O�5{ԡK�Xw�%�ꒋY!D���"O��׎Lh�����[�,)�蛡"O���f�J M�>Yҷ��v88k�"OЄ�AA�پu�O�h�vի�"O�]!�OM�.���3�NX�0�T�"O^����L7�l��&�H=�>�[%"O�a�<)���Ж�!{�(h�"O�)H���3�fY �0]�Z�� "OޡJ�mR�E�bE��gQ]����"O���F���F��(����D4
�"O��I1IN�UT�H+􋍧%��q�C"O�m��jXp��S�*�)��H�"O.,�� �.M��ka)]�zs	��"O�D$g�/WZ�'�&\b�t8f"O�^'w���+�FT��	w"Or����[�V����bQ?'�jx�u"O4��'��!'nD�yRf�<�Z�c!"O��ad�ыd�,\��%G
��u��"Ovi��H��J	��W%9��H��"O��r�ӌu��)�A̤FdxK6"O$�{����}���%oƻ-X ��'"O��ڥ�

f�n�㕮�&8��#�"O�e�r��ؔY*'�]�r%z�$"O� ;�"	7�P���Y��Pf"O��b�.��d��bK&j����"O�X#��Q����u�Ȃ�~�Q"O�p���S >!B䀕:p���"O��v�� ���D�D�7~�D�O�Q�g��?�H� +�|��O�����].���$��1>� 
�$t�A���?F-X:�py�� ۖK. ��'�cшa�C(7���X�����p����[N�u����O�蔠�>&�ҍ��P��l�H��V&Z$�<� �>Q���'`q�U�'Ox� �� s����#�(dl�L �DE��) gh>}"�~����:����rt�(x0Q�Jx:�%��_7,��	3D���
:Ƹ�Q��ɹN�N�!��O�t��s������V4�S�*}�����#P=�5bɢ-��Tx��Y���=���ˇU����g��	���*j#�2��$k��x �j�#H�ʽ��>��5�gy2'ҟ����K!u���1��U���'���.:�a	8ҧ�%:� W��`��F��'WPF�)Ѯ��vh�)��VL� �@�[Z���&D
MƢ3*i�0e����[�	��x8y����y�Z20R\|+�{Y~��	��y�"�#�I���٦he@�b�ݼ�?12�%k�u�vԭ#���㐂����Ih��1���	�"�.˞��w��f�������9A4$�wM�O�aa���a(��&jFq(�s��[�D���N>y��>�D/\�2�T �Iѐ9��!ƖZ�'`h��dou�cR��Z�)�!P�H�X��@�Y�v���p�'��t�_X����)ҕ�v��Rdۈ_�T��$�0'�P�Diʍ�(���hb���:%���Q�I��$Q�"O�X��I_�Phղ�B��>����5_��!pE,*+�I;9�|u���w}q���ΧnK�U�ck)N�l�	���ͻ\�b����Z�)t�`!T��>�Ms����~D|����.���f��c��}�w��)B��_r~� ��n�'P[���	:S�T]���\�q�l}X�B�Y#L%1�A;�|Ъ�O��2�	"�I�o �(�ĦO9�$e��I9 �T,FyB�#j���Ϲ�y"f�8�@�f���8C���0w�tP����-!G0ԅ�S�? Buа��"$C�*��]C:\*�'ԇLn"�dP�=�Q�I%pVE�p�V�&Aq�]�c�Xab�Q�O��yҥ�K�
����ٕ	�+)P�v�tyWҠgn��e�wp5
��|:�f׹b]2b�����	��9J�ϗ�_yy7,�O|�i��\
69���ʹ?B�д��=J7�!Y�	��$��NѲ���CY��0=�2LKiԡ����c��<�T��K�'�ZD!�	D�2��Y���FYE�f��b�\l����J�$L�`�L%7w.�z1m"D���e�Ǌ%����AhK�_'�A*���O|�`��	�����RhF��fG'���?�b�� ��9p7DJ�P�|`K�f�	�R�t@�f�O�pd��"�:xY�ue��7�`X"p̙�p��ɰ��YR,�y�/'͌a+�>O��̚}8qO��r��>	��#ɏ\, �34��/e�|�'�\P�7�\ʞ�X��A� |��~�b���-�������G��E���7��*�'5�l(B�lx��0��3��H���i���ڥ�Z���US���驖(߮\����2��@鰡\_�'Ra0`봢׀s
b-���T$Iv@8�Ǔ_�	�lεV�(����>e�B�4������.bu�mAu�*�:`X�4^�B����Ϻ)�F��5����7�-�I_F���ᇃX|y��_=k�:�'5���G�|�@i���i�&hб@�]���/�Hd	x���ng�(���/ݸ��6�X�E�&���'�2�K���)�I�哬d��s�R:G�X,9��_7X4�J��X<>�<�+$K#��Y��-g��ãoS�E��l����L��(�8Wa�<K 	)�O�x�6/Z�t�h�挶�J�`�FM��@��.V`�X+��
Ra�ty��@]�f�x����B�0�O��Z'1W�l�QvɌ�z�6x��Ju8�Г5FX'6 �����*E֜�Y�L�.'W"!�!٬A"1�CiA�L���"��S�@��b$��=�����O��(Ҭ֢
����4�N'�y�#*���
�Q�@k��Y)��I
�h����Q���bd��9F7^� ��g*�)��خESv��!�ֆH�,-��)V�	TQ�`G���h�I�H�r��A��	qz��1�6�L$=�Z2x�̴*C)o�B�	��R��M[V��Pi0IqaM�+7!�XRr&_5f�ĝ��8�r���!���@��b�$�7�8�B���>Ip!�'
�|�v,\Z����ӈ��u5
��C�%m��7�ܿwv)K4�ǣ6�t �tMX�7���;�g1A�t4ΓNҊJ2*�/)!�Iá1g�t����"�O.bR��*��}�Ј��vAly1$@{U���j&�<��DFj��'%@�<�(.��O�e(��:sv�����>�z�
Ód؍�CD��v��8,O��QR�@�)� �Y�`������cH�&`�I�	�h)�Ώ+3�g�(H~���΍�-	�\���o^
	�Op��M9ݸ���ˡ#V��He�նN�&����$B6,�C"�$�HE�mS�h��}LIc�����K��&X�lT���O��t�\�\���UaZ0��铄~���
��9/QԪ ���:� �K�+��R��<"�cB�����2���I��l@� �g����(�B,��S������86������	���T�Fܧ# R|9vE�}�p�P��4�]*" %��*#|�'9���hG'��X1���d�4`{�'��,
���J� �O�>m2�n�Y:Ɖ'/B$z
u�&9D�d��ѹoF�#��
�a�3)2}2�$  �����d��*EȵQ��}5��*x$�	�r$3�O���+I'X�@��E��$QV���l�@�ʍ$�J%�x�+�+Z�r��l�	2q� �`�/��O���%��#K�x�0��$.�13��[�eV8(�y�C��y�b\w�X$!G18�|��Ï�~R #5����Ep�퓡0}��Y�CU�Wj� c��+g8*C�	8o��ĩ��S�}��B�A�01��'�,8y%�ed�5�ቔ3�]�A#t�D�b�3����ÁnT<�X6�J�N]���`B�0��eN]�5����'���*�>
:yyt�	�B:�	����'V�.�q��+�S�����t1��!�*����B�I7"�*`w��U��ۣ?�ʓ|N��v�&�)ʧLAї��	z��.�1>�H�ȓRq2��ʐ�@�$(�&�ܤ_��}��\�N�B��K>%-��
�ǆ����ȓ7�l�E�N���r��'@/]�ȓ \��@7�8�X���,S d�ȓ,���"��P����w�	�H1������W/^�<�h�p'�#�̔��z����G��W���p�X�Z)����-�vx��'U) ��kܱT�!�ȓGd@�;���c�ʈ�dAǱCϐ��ȓ�6����ɨ|̔�[ר^�&8���S�? ����_�_ި����Lp0})�"O�[W�גP��s,�}}�8Xg*O%��*7<]vl 
 .���{�'���3��6�r�����%B��`�'��x⣮(d "��f�ġӲ|��'Kz�Xw��<Gւ|�щ �:]�	�'�@XЁ��M��I�h�Z��
�'h��:�UsVܹ�c̅~b��
�'���;sCȧR�=:�a��k��=�	�'��3��Z�0�戢���l�L���'�
�)� g�f]H�Bɖ)�p�')t`k�h4L>���`�''�tx��'�l}�	<I��;���"���#�'4"m��,w~RpȢ����:���'�TJ��ʎ@.`-2QW/s��X��'����!�J<~� qA,�wk�yA�'�a@�:c�ݑcG 6���;
�'W��j3 ��)���;49�	�'�t��������)�0U����'���h��-��-P1��0��=;�'N<U�b ��t��4��-|�@��&.D��!���$_m��%f*HȨ�
.D��s G�gc���$C�8wN�ar�3D��Y�E �TtHl�šRqH`r%!/D���GB��ҩ*q������(D���ai��3�lN�� n$D��S�B�<"v�xU �Z4�ӫ7D�XsY�1*B�
��ˤK���'>D���r���"��`�S��54�0��?D�d�ԬJ�w椡��T�G���B/6D���&N,����4�FВ��5D�|`�ߣw�蕙$�m�:��d�2�ɞj�$���B$��gh�N�c�Pd��BN�A�%��3tv�Ek)>D�`҂���Q��
�$)�m9�#!D��si�;D�������
}{R%�v�?D��Q,�V�̩�J�a�i2�	<D�t"��B ^�^�&N�KD��=D���N�l �M�U�D�N�,�{�:D��A�J�B^��TG�iˢ%5D�4�����v`T%R(T�PHg�>D�*"��%	�R�4KS%	��|:2*;D�Dstf�kX�u䅴,f�}�֥�<�V��(HE3��"�	B??S�)�ȓ<O8��/��^I��z�>t�E��o�`��m�F���Ⱞ�2���K<贌�"9�\�JD͗L{�-�ȓi[�,1v(�{ m;�aYvrza�ȓ��e��B�/j���LA�q��Ex�N�?:�� ��O�@] �[m4�)�G�q�0C�;O���V��z5�-���0|:taQ�u�f1�'�ʠT9�M�VIa~ro\A�p��6�:�T?7��2�p^P��I�[��婁$EXϖ��=I�#�S�01�f�^�5���3O̺&��˓{�г����E9&֤�Y��D Ǯ���dO?=rm
i�OQ?�q�FΰH�@�Ph��Or� �`�Gh��h��ӥZͪ�0	E?S��}�oD:w��\�Ō*}��t�2����� ��w
�;����X�!M�>Oȝ{�F�F�rh͓ӆ���X���B�<ER��� ʓ}���ȓa��p��I�<�~P��/#<�x��zc@�k�@6v6�$�f��Q��4�ȓ��@�$5ָI)3�ԏP�^��ȓ4@���RM��,�ڌ���@�V$舅���qF�
0-*\#��A�>���ȓI�q�$�$P���w�}�:؆ȓ?آ�r�.O�Y׼��L�C���S�? Tq"Cnذ0���Ɔ{�aXQ"OhЛ!��$4��֥�@�̛7"O.E��jȿlͶ�r"e�	<�~�""O
ŢT�^�j��`w�&r(�0��"O���וf�8z��>�du�d"O��s�S�d�Дh����w�v$P"O$��!��	���F��"�"O��iW6\ѐ�R�)fi("O2�+��W)V���*!mɠ[�x�Jt"Ol�	7 �anU�d򤸹"O2���!���(tA�*́_�T��q"O��˔L�7[�P�6�[�d�J@C"Or�	�Aq��2i�3�Z B6"OL{q'�B1�I�m{F��w"O
P�6��5g���PD��oJLѧ"OU+���;��i�g���zA|�"Oj�{��^������̬S^��"O���W�� ;���5�	<ZN� �"O��Э1jKD}B�)�$ao���2"O(���
<;����h�QO����"O>��/��(����ҋjX���"O���oH=h�±��H^l��ԩF"O*�K��.�z��1��"O0i�EMƈjcHi�SE	�6��ܩ�"O0��#NE�@����z�%�g"O��1G��L�t ڱC�#r�y��"Oٛ�@չ&�FMiQ Z�X�a"O:�Ѫ�!:D�����M��ڇ"OA�A�2b,�\�GM�5$�
�"O�J�g��`�,���5�"��&"Op�Y �߂"��h(��
�V� �g"O2�����i�2�f���@�#�yo�;�-cO��.4��UI]�y��T:%����Ƚ.��P�����y�e(6b^�s�[U�Hd��,�y�MC�r�ah&LP$}�(u��H�ym�1:���ic��D���@$N-�y���4Ĩp� J��@�50���	�y��k�ڼ곤՞mZ��$���y�M䂖4���*PO';����ȓ4v�T(F畴 �J����+�p���M��ŢDF��- �]Ҳ/�#>�h<�ȓ=:�m���V4��H�j
�'��ȓq>!i%�@�<8u҉r�̆ȓ)����3*������z�ĸ���� ���(��б4W=�d��V`(�-������� p<��ȓEwNA��a�Z��i�&#��:؄ȓvM ��A�B�A�(�%����@��ȓ%�-y��B�|�%c�����0K����N8%�,;5B1tt���wʠc�@�+�0�j ��8�0��ȓ\e6��&lߧ|ΰ���L8X���
"�Q�Sm��f`LU�$�@7."����S��(� � b�WYװ(ab"O�5�tNF�_l��Qw,�P�l��2"O���4&(NFp��K�+�8���"O��	�[�r�J͏�n��"O�9;0FLJ��-k�̍&:��AS"O�@�C)4h�qr�f�X��!��"O ��`W �々�;g�b��"O
%�0�Э}������N.|A*�!W"O�T��.\	؞P�BD�	a��z�"Oh�"#b4>�:���"Y�B�,��F"O� Z��f� �Hs���5�LX��"O�t Ӆ�eh�U�g��-�lH��"OpJ7�_�WR1�´qNT���&'D�x��O�^M����5Z�r��b)D����SY-֐�t4%��x�@*T�8yٱAE��"@D��P>b�:�"O��!*1OP��d
�\% �"O�"`EE���5#�4��"O]@���!���N�8�0��E"ORͳc'^M+R���O��i�"O&��ӂ/�h-+t/A��X��"O���Bi�%:GE��dI�c"O�v.�0�T:��W���9"OP�R�f���i�d	|�m��L�t�<�,O�'�l�p+�@��1�F�p�<	�d�@=ڌI4N� F�tq�k�<�)�{�e�Eȇ"�Va��g�<I���L&P���/���Q�C�g�<	�Ø@�p� �G�WY<� $�}�<)�<P��;#�<p����w�<�Ad�$�V�*�
�. �,
�mw�<I5dA$f�|4���|���� �Lj�<���Y��(G�V���Y�4b^g�<��7T���9�f�� �0p/c�<1�h�Xy����:e�PDg�<�v��t�D`�d� �D��$ƪ�w�<�HI�1�	s�aIMhڔ���r�<�i@�T��.�=�bAK�I�c�<Y�`S�R�F,��kGv�ɂ��J�<9 A�7M^8�to�v�����DZE�<Y� ��i��r�M��A2��B�<C�x H:��%Q]�JY�<Qs`�!R�:��86�@1�W"�z�<Y`�[-r�������?�*��N]x�<A���%���eH�-cTZ)Sр�q�<)шV'&
9�a`�g�Lzf�n�<�
��~��� o:H
����h�<aU�մL���+�f��)�fdCULd�<�1E�"�S�"��P��KX�<���U�P�ij0��_c��9��~�<I.� � ��*9���Nz�<94Ô7U���r#@ǜ"B �g�Fy�<�� =a=D��pD�{f���r�<#�W5U:��T�ҖZ���c�<q�U�>�8�A
��G~�lB��{�<��M	T0�+#����D,*���y�<a���U�Uã��6f����I�<���*�aahS "P�Al�B�<� �1EV����ào�rQCs�X@�<qf�sz�CGX�ZF��A�X�<)�� �����Y� %�5�S�<���'�tTG�{0�(�h�I�<9�-*Yy\@9`�M�T)x���yrO�nY���F�a0�9 �G���yb'�g؈tI�ǘ�`��������y�fT�z��9RPՍK{�q���y�'��wgP!Ã���Kg�$iG��/�y"D�+;�,����@FL�2�5�y2!�<�@i�fR�=h���ъڽ�y��P�%̄M�c֎.L�8�料�yr��<Q�H��@�C~��i�a���y�ᚐ}�L���cZ�y�N!��y��H���!��@�H���h���y���*�0%صL�?��� P�N�y
� R9
so�*�괺b�V�VZ�Y�`"O$�#�*��	�$�x�JX7A>ꩳE"O�I�@�B [)��׆�;�9�"OƤ(fOH�+��4��2+̱��"O��!v�«ZI��DdD�3@zq"O������z����� 2��9�"O��sdеHZ��C��[�?�����"O̍�2镰9�Hۿ$,�#R"O`- �>H�rI�dL�>L1�5"O��HP���`4����ݘwni:T"O�(�R�]
5�\rWɎ~c�ث�"O��Ѓ�: d6����l^ ��P"O�kq��
>�R@��lΘ7��ܺ0"O�����?'L�c�D \��� �"O�|���9;���c3jC�)s.��"O�	b�� �< ���Uu���W"O��êӠH��TOԮgi\��"OR|����,��+� ƣP���2�"O0T��O"{XlPd�Y<R� �ѳ"O$�d��&���s�(��K�����"On�Ht�3W� U1�(�	^}�d�7"O��U��'���:3H�m�ؙU"OL�!rX�S�A"p!(H�t+!"O.�C���*0;��M�-3 "O^-Y�C@� U"�n�82x�K�"O���Q!�dM��P�=s�"O �:��ܻ=�T���لj�41�e"OR�K���q���@$U2l���"O�	� R���	B��m�!��d�*��5͎�)��Bg��<]z!�䙯z�n���`|x�(��''q!�d�'������ҕBb�a���&3!�ڇ8�$����RL���pƓ�L!򤓶G�Jd�%c]:��ht��%}�!�W8{��E��Ŕo���Y�É�a�!��!Mq����EX/}��IqR$_�l�!��%\�XLWˈ/	��-�G��
v!�D�	��4PB�ȝ �t��(�	2}!�$��YoB=�reB;����'AI
!�	�g�v�ۄ�H5�Ly�g�T�!��:(��k�L��k�6���kG!~�!�DEZ6\ܸ� �: �P�6ˋ�A!�/b� u���56�\�HD����!��Z2xb� =0\�pKT��!��4l�,J�m��f9��wo� L'!��ʕMh Yւ�P�ȑ�m%!�2+���EB^q�3��/f!��\ӍȐ�ܡIQ j�!��U-_�L؁��!����z�!�d��Ld�j�OM����Qf���':�	ph��A��-�Q˞�W�PIQ�'�,�؁�${!r�Q!#?a�j����<�@w�[�(AYH���$Rvi��&��(s�T)�xP褉�*e�Q��i���*��?,�x0觢�g����,�&�>��~$mXCeC�y2�ɐL��K�	�a'ܩd,\.�y�垫3"�q	�h׳U�b����-�yNJ-�0xc���% �JQ�U��y�&:Heh��י��-�GZ��y��z�������� ��S��yR�P;3 @  ��   �  C  �  �  �)  �4  J@  �K  W  /b  um  Ew  �}  �  ݐ  !�  m�  ��  ��  C�  ��  ��  l�  ��  B�  ��  ��  Q�  ��  ��  �  	�  � 
 @ � ;# (, l5 �< ,C oI �N  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t����'Q��y��ɗ~�����˛[>��f.#D�����?�� [3?�$� ��R+Q9!���B��@��[�r� `p�O�a!�X
tP�A�����i���
�+!�Fd�ͱ3�Ʋ}nd�2�Z32�!򤐞_ے�j��.lw�I�P
�*S!�D�P�	Z�*͖`�m:�H�D@!�=��ܢ�'ͧM��r��T1!��Ѥ���HV2<梅k�e�!����9ysN�@<���C�=@�!��	;�Z�p���|נj�]9/{!��\�j��!�c���lB�nz!�DԕS�`����NK��` �H�Dp!�V�18^ ��m(+>�PI�D�"]!��[zR ����J$�ɩ�MN�?�!�$�p��1e��	*�bT�M+xr!�T�+����SJչB���I��I,7!�҇ |jxK֩�9%�y�VAUj(�O�A��	�ת��d��nE�\�b��*"B�	��PasB�V�I��,�B�		0���aB�U�7��PQ$�Ǥ^C�	�}�����,;�<�V���XC�	�*C2͐@HZ 1��#t��� v�C�I%v䘬X�͚9y���DÄ5nC��<�L=��)�>�)@�&�/1�JC�	3u�j��ܻ+3B��bFL2=C�	��� �-��(�^���
�B�	�Y�|[O��ft�p�]{��B�I;�J��r��>P�8Pq�-V�>��B�	�#����%��%6|��̗�a�rB��:T�`�f�Su��Xu��,]�6B�I�)����U�8�m�񍝒p� B�	&C�8�D�e�$���(9� C�	:��	k�4%�� �i��JB�	�z�~h!!�I8?���1ׇP�`C�ɛOtAY2�Q�"�~�3A� ȘC�	�J�Jݰ/�E-�u�XS�'��c�nQ�w�$DCu"�t*d�ʓj|
`{p�-E�P2R�P2gi�� ɶ!y'iĆh/���ec�l�T�ȓ���@��2"
��P��.v�E��-C�x�D�''��`�Wg��oc��ȓ>'x � �
�w�`�I�G��]���"��d��aK��(�)�5d��jc�ݷy�!�D�S�6T����*aY2��C�N�0��DF�ă@�06��LQ�,玁6&��y��p	�y�f��(B\����
�y���8�2u*0�K) D`�HԠ�y
� ��Z�M�=P2]{ �Jx�}��"OF�ICmS,n|�P*<aXl@�"O��@�) |"�89c.ùN���"Oԩ@@�Z!&VUrw�P�;�B-0�"OztHԅѩ@F�¯Yo�୙�"O�`+'"ɎZMLe�C��3���q��']"b�TcPI�.	f�BH�M����1D�����^&$�t<����8�@���'.�	a���0�o�i|�,��G�}����?�O:扇A���hQ�)�ȩ�g��-_�ɰO|�"�˽o��5�PM=M$�]�����<���0��=)8
DТ�!d��7���V~lC�D� "�*3SG�ѳF!@�l�JC��n�lZRD#�`5[�8�:C��Q��􈅠V�M"i�P$Κ.(�B�I�M�`��C�A9_��� �
{!vB�	�_��ղ�`U4L=(�oE�B�I�:S�,i���`6�Y C��|�����>�6kϘ{C�q��É�����HA�<i�N\� j��ÄA��e$�	��O{�'?-S)���.�(�ƞ�/@b|��d!D�L#�X�Z�4C��\9Z`Hҵa D����M�'k�����C y����" D���6�	�N��b",���
��<D�DÖ
�"��8 Fp5�1v);D��je��!�h1�5%Ҏ$�Hm
r(%D���-?"(�xX��Z�ԌЬ!D�dHET6w�$@����@��L>D���"�`Lرt�M?�R0�7@=D����Ȯ<�*�b�̐:h�|S�:D��R�͂&���+�M�kCȡ�2o8D��p(B�;.FXe�~�ش��/8D����,Hh��l�'%8�LJ6D�h@T��_0>}3��G^R��ti6D�Ls2�������Ӕ-��A��3D�8�@J�"Xl�	B��*�H%��	1D��4a?%�r0�S��j$A&�-D���ń�_��u��m��"�D�8D�d��.���ĈB�
� .�[�8D�� e'NO��↬ͦA ة2V	)D�X�b_+;��T�����N�d���(D��Ð���	���ǉx�
q颤#D���5�������  D�<��ソ:��2c�C+N>lз�0D���$A�0�`mpt���0]d��$.2D����ve�@CU���}},�b�;D��¥e�-A/�0�F�P xJ�#�F7D���MR+;��Yx���0�!��4D�Zb�ӹF$��W
��;gE�)5D�̚�aU-/kB٣�5(	JWj.D�0r����E7p�z�惿e5(�B0G1D�����M�/,���!F��z�1D��x�]x��D���P�C�1x@�.D�|��ӧg���Q�[}pJ���9D�� �)����q�W�SE `�"%9D���#��704�x�������Z-$D��@�$��V��¡h��z �I1gC"D� I�f�O �:tBKֽ3	<D�� c���3n����U8��v�;D����j�)L*�����AF�;D��*��Ln �|��6P�ӳ!.D���!��܌a������]��n9D��J���\^�"g��/f�AqA�3D�(Rw�'�8��E�f����E 7D�� 4�P'�3>p�PT&�~�P�"O���A%�@Z"O�-XU�݂"O�×��9V���j\�z&"O"���� %C� xq-ť].�,��"O�p�+��`F����) �wX��f�'�2�'�R�'���'H"�'��'�,��P�Ղ8�.dZ���䅢e�'��'���'g��'�b�'���'�`��^��*\�P��uZt�'��'���'���'Z��'���'�r�T�ƣ�����F�,"�f�1��'��'��'���'���'���'�j���AI^r��'n "^��{�'z��'��'���'aB�'���'t(
��C��}�����~����'C��'���'�b�'���'�r�'M&�k�E^0B�6e��Y�=a:l��'I��'���'���'���'B�'6Ԉ�vnʆy�1�0͟6^�Y2�'�B�'���'�R�'���'��'��E9��ȳ�B��JD�xx�A���'2�'U��'{�'8��'rb�'�U��挧z;@�k��կ:���3��'qb�'Q��'B�'-��'��'��x�I۱A���DA��u�P;��'�r�'/�'�"�'�"�'R�'�,��"YI��$��-�4&r�-���'7B�'�r�'�"�'���'x"�'9�ȱ�4H=h�F�L����'��'2�'��'�mxӬ�$�O��S�	�[)Fh���Fp�f�xy��'A�)�3?��i�\�犂3F[�ei��"c�DU�2����DIȦm�?��<��r�"���ȶH��хj��?���!���?�����Mc�O^�Ӓ�RI?�x�΀���U��E�w�,4H��7��ş0�'��>QH�HqP�dc���4L��ꖋ�Mc�l@U̓��OH^7=�.9�Uށ}߰�#���'8�ZT`@��O`��i�p֧�O���Yv�i��$ˬXX��pD��&U�A�DC5/��t��a��dO6�=�'�?A3nS@>h�@V͉�2���PgJ�<	,OȒOv�m|~b�������8��������%-�k�G���П8���<��O(�E���@UHơvm��������I�W�X��I(�SV�IHT�qc�,Q��'m�����zF+ey�[���)��<�	�q'lh̝I�-h�QΓlm�֯H-��D��a�?�'|_���1�F-�,9�Ɣ&&�*d̓�?����?!e�Mc�O^�>�
f
�0<�e��k�*�����w[�O(��|"��?a��?��g	�L+$�C�;ΐ[uCA!QS`1/O�n� T�
��	��$�I]�'C�a#C�ym��GG��J���T�H��ϟ�$�b>8��۫��xx�O
8���Ҡ�D]�`l��ߕ&��$��'�'W�	�qu�0��h��(����N%+��	ݟ��	؟��i>I�'Zj7�ݙ$���䙙:B��:)ͅ44Q�a��.Jd���黎�?y[�h�����	&�u �	/`N��C�0KI��q���Ԧ)�'�,��K5�I2���)8Я�� �4�i%��L��@�"Hf���Iߟ ��x�	ݟ���pEɣAz����Γf���HM��?��?���i��}H�Q��0�4���$����vr0��K �p�t\�I>����?ͧH�
�4��D�6a�t�kD�K����p�ķhJ,������?�j9�ĥ<�'�?	���?��H�}$�l	�)�-XUc
��?1����Ě��{�������ğ��O��}��c�tĨp"�[�h��d��O�h�'/R�'8ɧ�I��t�zQ"��v�0����I�#`����Hf"�9�
�<ͧ �,��]���M?���p��.C<��h\?(Ox�p��?����?)�Ş��Tݦ���ЦRz�)���Ow�9!g.�2K{a�	ҟH��4��'b<ꓥ?1.�Tb�0{R���g�H�����?�(�����4��$�5̀�z��t��G�����k\�3��&����y�Z������������������O
������l,i����qӂ��š�O����O�?e����K�( C��+ъ_�R�m�Aͩ�?�����ŞD�@޴�y���Mvf���Q����J��yrg��`��������O<�Đ�gа	x�F4�"�1DM���$�O���OvʓQH�6��&Z���'����(��E⓭�Sȸ��j?
��O"��'#���4'�����k��^�� ٿ<����-L1b���|�=&?	r��'y���!,2��%g8��Ҡ/B� ��%��������(��H�Or Y.���7	Ņ@$�8����m"au�|�Ȥ<�e�i�O��X)�F�J���7{p��m���d�O:��O�L"�Lr�@�9�@���|(+r�E)ydt���E�Ԭ��I�4����4���d�O$�d�O��Dŧm��Ht�N\Ӟ���	�� �'�v�ӺM%2�'C2��$�'�=E�Zp�
���H�H,�j�>���?	N>�|j��(�d��r��]H�i���9��48۴k�	�v�̀Qe�O��O�ʓNX��HfE��:�K�&-x���?9���?���?�/O��lڥ<d���Z ��0�&�iVP!��I**�t�I%�MKH>����	埤�'pz���K-��p:���i�Ka�B�>�&7O��z)���'X˓���{�? �P3g��D�3%Z�1$�D�u1O
�D�O���O����O��?Q!��"j���P'H.6�L]���՟,��ڟ2ٴw��*O�Yl�`�^��ȗJ�H�lt��T�dC�%���I���S�Q�NmW~B���yD�9Ӷ.'W�ɑ1O�A4Z������qb�|U��S�������\�G+�L�PdC�N�F��LZG�� ��py�*t�pQ��O����O0�'x�������I��@��I�,�'#�듢?�����S����T��#�N�r�,C�`� �(KuH�"����<�'I��Ip�ɓ_�ԸA��	=B��)c�*G�O��	Ο��	��\�)�`yR�~ӂh��4w�j�Ώ5O|
:g/�������O�aoZ@�9��I���BؾfHu����$J.��eޟ���)�(oZ~��	R	r`�'��DЏv�-�4�K%02\�!*�0y��<����?Q��?���?I-�
���Hw�����'_>҈���M#��0�?���?!H~Γl,��w��	�Rb˕4�����ī�
�0B�'��O1���p��v�X�	>���xĺ���!Q�p<s$%f��x��G=a�b
�a�	|yr�'�2$m�2�r�nĳG?�@C'��{)���O����O�˓:囖D5�'2B�9�:�s�b�6�@�Y<!�O2�'$��'��'b��u��
@t�lݔPX+�O<�q���=�7�-�S<�d�O���c���X��})&�*��(x#�Ob�$�O���O��}����񴄚�F*=s��J*�Ԝ��Q��IFgj剩�M#��w���ȶ��?�ȅ�uN�;��Ø'�R�\H�$����'�����?���NԜ>��,�ŉ��mwr�r��$y��'v�I��Iꟸ�����	PN���&޳I;�Yhb�
1K����'��7͗4W����O��9��q*<X�g��E,�h'`�,OR��b�O��d�Ob�O1��`�"�#~ y�d\.T\�#�ǭ6�7��]y�jO!,l�������T2(�1ҩ�#OL�I�"Y��&�$�O��$�O&�4�Zʓ<����#Y(r+��Rb��q%�
�&��)"V�A��y�yӂ㟤1�O����<�v�� �:S�&}M�Y�k��U��4��dB�ZZ������^�����^�%�)©�$���;@�)V�D�OL�D�O�$�O��D;�(aG&��B��P�@�֪�,���ڟ<����M;���|Z�Z��|Ɔ�P�^q���bABm"���Ji�'����ԃ-}v������ T+���˱�ݑtʔe��Ԋ	���j��O��OD��|���?y�[U����.Д^����eѢa��\j���?	,O��nZ29ry�����Ip�t�V"�؛  
U���z��ݧ���W}��'���|ʟ:y#����g��@䜜�*�7��7Ij��s�+�i>�0�'(V�'�HG�H�a�~�2��ox�maq���T�����ٟb>��'(R7�P�ӬX�������
Svк%M�O������?a�[���	�6� ��Fg���@®�2I='�i��iW��.oB&�YP�O�z�'�IK��  9v�C�N?V���'T������	ğ��˟��������ڡ8�#x<�5��D���7M\�"&f�d�O��$2�9O��oz�	
#I� (2��	H�>�(�`�П�	n�)�>#�5mZ�<�! �g�����i��upn��E���<i���|�����䓖�4�J�D��X^B�aF��<m3H�iRAܤk�v�D�O*���O��<�֋���'���B5z�0x/Γ�bl��%T�O��Oҽ�'�'��'�������+uŠ#��)!�O<�	T
�<3�7�Qo��+|���O�U �HY�MQ��X:~8��H�O�D�O���O�}*�G7F����˴�AsC�r"ҽ��ƛ��-?j剏�M��w'��P�v�t��D���l��'�"�'@� C�����@�߳[f��J®d崭#bg֤0�&�WB\O��&����Ϙ'ݨ\i4� 2f(�ũ���j��t��O$�n��L��'���	J�
"����N�;��Ԣ��?:���'�2�'�ɧ�O����Z��T1����#�x�r��"���^���5�E�_{�"Hi�Ky��H(�ڕh�g���`�YvE(�0>餿i'����'fP�C# 2�Z-S��L�]�|Qɘ'��7-<�Ƀ��D�O\���O+K�.��l�v )$a�]��섿L���jܴ����>����':(�����>Lm�d�e�U�-�eK�˜<l�D�Ol���O����O���0��:B5�'�W�V�n=�̔)\�F���ҟ�	�M�����|R��|��V�|��c���t���	���&X��4�|��'��Ot�xx��i+�	�29�lⲣU�%��XAkF/,������.?��,��<9���?q���?�� �E��I���wO�ɂ��Ν�?Y���DQ̦��t��sy"�'��Sq��TdH�R���ǦY�*�����I����	y�)�wπ�&o��(`L٦fBl��d|������ŗ�M�WX�擊*��9�$QL��9%/�7	����$$�*�$�O����OR���<�5�i�X�����{��2���84�D��5c*nR�'��6�4�ɕ��d�O��xPH�18���h�f�\z:�G��O ��ΐGD�7"?	t(g<��SUy
� d����<Z0x��&B�q:���A<O���?��?y��?���򉀨D���C�H�`V��]�I�|�oZ�>���Ꟁ�I@�s�p���P-U��l��c�ĺ4�<0�oЮ�?I����Ş�a۴�y򆞏G$��r旲6?������yR��*v|9��䓹�d�O����?M@��1��>C�F�{�� $P���O����Ofʓ^s�V�7z�"�'���	&[�>�f���]Z<��������O�L�'�b�'R1OL@�蛫{2T��	��p��c�Of�P�ɏ=��7�$�݆�	ퟌS�$�=���%P�eUF��H��ϟ��	ߟ�F�T�'�j0[��SpnzT�2�Y�o��P��'ת7�D���O���ΦY�?�;a���f��))A�B/�4H�*���?���?�抔'�M��O�л5�S(��$B� ^o6�*qC�JF���jH&P#�'K�i>��	ޟ������	8;�^,x�R3[M�qq��-\n��'��7mY�Tod���O�9�O�p�[����(J�37ʛ�,Q��O����OڒO1�n�K�JE�o8�ٔH\�W��y*��E-b��6M�@y"�S�?h�������'��>!��5(�o��-4 Y[d�'���'�����]���4:`)���uMJ�DcI���j�/[�M�F�I��:�F�dM}��'��'2,t�̧�x�0�W3�p�pB�ТPɛv������HQ>��}�xY�Av)`pcU�5!����9O��$�O�$�O����<�|�U,��P�d�5��"�N00�C�#�?���?a�iV\qd[�$��4���Ș�%�Ac�B�L@�|���H>A���?�'��}���
�h����Y*<
�lKu͙^;BA��1���D�6����4���D�OZ���5_b��!��I޼���─b����O(ʓNH�&E�/|r�'�Z>iAt�؉lh>��adY��[�5?aS� ��n�S�DbS
-t%	�X#P�7�R�N%6���c
.`'��ضV�擌(��c�H�	(	��y����=���z6�:������T�I��)��fy�	k�`�OU1w6F����q��.�^��O�Im�@�$\�	؟ C�MW�"�&�:��A�nQQ �����E��mZw~b��	��-�'��dGGpţ�+۫}�F}�1*X*F�İ<���?	��?��?�/�2��V��4�����ԜU�8�``D�}ٕ�F��	ğx�b%��y�#�V:Qk�G�r�ڐ���ڭe~b�'yɧ�O�%x��i���L�`+Z�B4�V�vr�1��U�O��(d�H�J�'��'��	��<�	1N���0�K1ڠ��f �&p�Iş��	֟|�'/6��-Q��D�O.���	/���A�794��`��u�>���O*�D0�I�!p�'�

8���CMV�^b�p`���@9=�Δ+N~R�i�OĔc��Eo�ؒ�#A�1�X�����M�@�P���?��?���h���
�
o���5�6�vk����d����%�ϟ���9�MC��w�5z�a��X�Yp4��e�X�p�'^B�'��P.��V�� �i�V+���}�Pl��Ȇ f�@�K˒Z6L�O�ʓ�?y���?����?��p�y�1�E�R��'B�B�#"�ny��h�hl ��Or���O�?Q�Vi
�c��8zb#A�]a���)�����O��d(���@)p9|:�i«`N�U��N�L�f�I�ay��m�'vrd�W
Mk?�H>9-O���Vd�T�$�0���*��!���O����O`���O��<Q�i^�e���'8Ӄ*��"���B/hϨ�ڒ�'^66�	�����O^�$�OD�#'�-(/�l��fY8�b؋�7}�r7�(?�a�@����I+����y�L��^p̫K�D�XĈh��	ԟ��	ٟ���Dy��Tœ�y�ĝ��*Θ{DQ6�fD����h����M�2G��|��0M�Ɲ|b扽\�B�i�gٟ%�t��i����'x�U�!V�U�'g� �D8no`,�DK�Z�`��6+D����=	�'*�	B��KLXqZ$�h���iÂ��T1Gx�!x�~L��ɥ<	���I�,z�>ѵjD� ]����F���ɤ����O���#��?E'���Z ��a�Jŵ"²Ѩ�K�q��Z "\��,O�I��~b�|2IOk:�qz"��r���%���'��'9��4V����4c�^�C6A�&N��hS ��H�(pQ�N��?���h���$LA}��'�:т�,!�`�s���(P�b!���'��\#>W���� �G��X����~���®y���/�܀���<�(O����O|�$�OJ���OB�'�j��3�Ar�Lu�W�
�!]�U��i�FYq�'���'>�O�2oj��/�2�M�)���FHȶ(� �$�O��O1��8��
gӤ�2,��hS�q�.�q�O/e��扏6�X���'��&�������'�D�١�ȑu]ʤi���:Bތ �'X��'MP��qش�f0p���?����Aq�咶��-؆(?���P�⌽>q���?�N>��OǸ"����nO!j�Ȁ�DR~M]0��!�i#1�t�{�'���3$�йQ�K�x��j+C��'�R�'�B�S۟�X6�(ve��9��@��ȟ�p�4S,����?�T�i0�O�NaNHU.Ζ|jք㑆�"]����O"�d�O萁�l��1�$�Y�(�?� �a %�.im�x�dC�w~�!�l>�ģ<ͧ�?����?I���?�狫���+5���e�u������S�	s	�X�	�&?Q�ɘ�Ł�႕�zP��ڜ)�xM�O����O��O1�ܣJЕ'qN|�5,ѐ[�=�e�.:��6m#?����16����I�	Zyr�M6�VxP��ޚ o$,�ekü@��'�"�'��O��	�M�����?9��
L҈��Q�"��N�<�%�i9�O0�'#2�'#@��2���j�������CK�2��Düi���-��PX��O�q��N߄�=  �(t�Zt�u-'o���O����Oj�d�O��$9�Sv��Z �y�$����V���	蟐�	��Mc�IT�|�l��֛|2�W�*㘙g�O�,>Xe��E;�'~b����ցu��6����ե
�x+a���AoR%1է�����'H�%�������'���'��Q�a]<|��5)��VA�ޱ ��'5�X�\*ݴ1������?����Ʉ�4]v�����!����Gט`@�	��D�O���'��?՛t�Lu'̭�C܁̂�	ȽI�ʤ9��ؚ9;��|�c(�Ob 2��}!���,� e��ʛz�jI��ЪA�J����?����?���|%D����-O�$nڟ'=`<��W�k��<k1��q�XLu&Cy��d���O���XK}2�'���:����glڥ�"��/�~(���'��J݇7�F3Ob�$;Z�ưSI?�I�1y��q��1#�za�I��5���_y"�'���'o��'S�_>}K��2Q��iV��\��q���K��M�����?����?�N~��V\��w��9s�m��� ��8e�x4��'Yҝ|��� E��2O���A�+�
"�P�
P����3O�`PI �?� �&�$�<����?�t
��B^.��2��Eu�P����?���?i����Ŧ�c�E��	�tS' ˡw�B%x��D$��Zșu����ɟ���A�I�"�bpb[� T,��AW� \��X�s��=5A��J~
S'�O��@��]�����F2���Ã�<��]0���?Y���?)��h�p���'f5���ZL{"$�����Y!����
ffş�	�M���w��A+㏐%]��� �U*pq&�#�'~��'�샧0�����k�\	����7XD�Q��!Z]*��;G.�O ���ObX���1S��r3偣#B�jᒟ4	ߴ7�&�(-OD�D.�jt�`+��@T��I�%��:�2�O,��O��O1��x���D#]H�t)Pb_�F>���j��-&5�%�<av�+=|��D��䓿�D�?v�Xs�䑫g����#�����O@��O��4���5��F|9�Ie�j�A�k��/.�r���o��f�ča}��'�R�'ޜ�Q)_o#��؄�&A����&�+&/�F�� �g`�7$Q>�ݽ^:T��G��X��0#� ��y:��͟t������I��	o��Y3h�[�G�9��lAf�.�����?���L+�F������'�~7M2扣�f�Z�̢7�q�̊�|xޓO����O�	�H	@7�+?a�(	/,��VޒFpz}�r�X�)�T�AA��'�ؔ'���'f�'�̥�3�N�p�έ0��������B�'��ɴ�M�f���?���?	/���pv��1Dd�Wf߃tT�
域��O���O*�O�S	'Ό�`��2&j 1㙜&��p��H�8�R	1��+?�'pB��ė��&3�����T�V�P%IC�9�B�+��?!��?��Ş���Nަ����Y�'d���G�M1Tk!	1,�ŕ'�*7�9������O�T�V�L�,��ɁA�ޜM� �T�<��� ��M[�O�Dz#�����<�dB��;QL�ك-�WcA�@c��<�+O^�D�O�D�O����O
�'h�l=S���C%�0��.o�Sw�i^���6�'eR�'��Og�a��n	&�UK�%�:�<J�
F3F���/�)�Ӣ, B�n��<AUDF(@�4[u��+	�ʰ�tA�<	��O3R���������O��-%M��!dMn�l��m������O��d�O˓?.�VM��H��'r���7�y�ŐAPf��nT�|��O���'���'X�'��Q���jy�l��BK�dz �'��5ӳ�Y�%C����3�~��'���3��	�{��t#ݮk���g�'�r�'�'��>	�	�F�����J�M)��vK�4pd�	��MSW�������)�?�; ��!զ�/v�Z�I��v�����?a���?��%�;�M�O��|���i 8�ᛖ���t�r�"��0��I>1*Op���Od�$�O����O<�(�L�.Zq�Q�3b�R`뗌�<�e�i�tQ��'G��'��OEr�U�5��(���RaX�I�/KW@��?	���d�г?�}0�*_dEK�[�*Ђ�]�J�40/OlA���?��5�D�<�R-\M� ˁ(�;�<Kbą"�?����?)���?�'����U��j֟�mЩI!�������"ecΟp�ܴ��'�&��?�)O������nL�ܺp���"^@��1`ٗXp@6�$?	1g��r�n�	����kW(\T�Dx$户z��|G��<I��?a���?���?ю��$�-{j�t�h�E�tmF&yL��'��et�n�7ϩ<9��iR�'EĘ�	�����!A�=C�B�|�'��OWF����iu��1��� v<�T�ڪ����V�A��$�˵'�#�?�H;��<ͧ�?���?y��3JY��BL	\2��ї*�?	������ѡ��Yay2�'��S�@� DĎuI�A�^�^k��E��IПD�?�O��0@fEL
e��F]�z�N%k�o� ���c���=!�i>�Z��'��%���l�(t<Ѐ����ca�5e��ٟ�������I��b>��'�7M�(L�J�;w�L�?�%oY�9��c�)�O��o%�k��l�>���e�R��'�F�]�t��A�T�X���?�sO^?�M3�O��M�W�z�I���Ā �l��tnޟn��X�Tk��,�<���?���?!��?�(�L���zmkҧb]�ӒN685o�a�@�	�T�Ih�S�(����f��*ӄǥ#���qR���?	����Ş3\ҡ�޴�yRC�"T�4�2��z<S�Ͳ�yBɵ/�n��I15W�'��՟��ɴ��* L�Jz@�81�]�33�<�������ݟ@�'��6F!����O���%@V¤#���1FQ��Q�}H���x�OB���O�O\�U�G�N�B0z�OQ<C2�u����`�
�ҠmZĻ;��I��`��f^N4��kQ�\�М����������d���@%?�I�%0�u�	���<��i��W������_�
<����M���4�?1��-�V�|r��y������+i�"���mӂ�yR�'���'?�uaW�im��O E��eZ&�
v�LY���u�N�F씐�W��+7X�O�ʓ�?Q���?i���?Y��`�@hȣ���Cf�r����m`��/OV$l�7W ,x�I�����D�s��b-�$0+@�E
R^�x��������O���#���ϐ@q����
��#�R�t��7����U�lӄ��'`��Ώo?	O>/O�IS��7�b]
 ��7�.�3��O��D�O����O�<���il\I�b�' �����l�bQ���f��	��'��6�=�����Ov�4�δ'�ͥmS����S|ɞ�a�l���7-'?ibƒ�9���)��䧲�#�$�'$V~q�Q� ΦD�����<I���?����?���?��dk��*� p��H��J[܀�9��I៨!�4{�z��'�?���ia�'� ��kS:B�:5��� ��X�|��'k�O)&!�i�	�=�d�%�-Xߦ@���L=,p��UR�8�O���|B��?Q�M�(����ޫ+�X��Q��9X�-����?�+O9m� '�V��	ߟ���m�Tc�:5~!�+��X6�h���$�k}��'Ur�|ʟ�Y�#�ه,����CL�9z͜<�`ʝ5��U��y�\ɖ��D�JG?�O>�j�q�^�"�N86�!3�B	��?9���?���?�|�)O0�o�X	�}�E�>AP��)v�֧D�ր0DYGy�ly�*��)�O���ך]��L�D�z�L,�A�
�s����OjEY#�w�\�;��(����x�O��4kWLE=�f��ӊ�9k���'��	k���rh��0���pǌ�t I�S����Ms�#�����O�?�����Æ!�=���H�^aM����k�(�?�����Ş%A� Cڴ�y��ֵ3��t����!��Ly�ʂ�y��ρ?�t�I���'�����X���f�؃,Ă{�F�;�a�T5� ��ɟP�����'b6�U0B"��d�O�dP0(p�z�n�.T�8��`�P:OV ��8�O��d�O0�O4�l�M<$�+4�݂0���撟@�WmX�:5�q��(��*:0����r0��_����U@�8�U`�I�㟈��ן��IȟP&?	p�f>��ɵh�V���ʓ�R��X�Jp�I��M;���?A��<՛��|��yG@��[��fjE&��Z%��(�y��'��'�����i����ON��
���vk$@i���lȟh�Ƙ�bOZ�d��O�ʓ�?���?���?Q�$w�����?J�4$6(Sp�(O� lھ9��M�'�R���'P�]��$��Ը`#�H�!�"�>Q��?II>�|ʖ�	$Y'�)HZ����� ��	e1x�xqOC~�N��`����$�'�剧IUB0�c	;	��My��D�;����	џ$��ߟ �i>��'D
7����4�$܆l�j�OE3jp:�!C�W{C���覱�?��Z�t��_y2.H�3X��4�S�:L�7�V�l�4��c�i����Z��B�O� �$?���*u�\p��1>I�P�w�2QȐ�IǟD�	ɟt��� �	}�'?����쏎l40�(a�]�;��	���?���l��É���$�'it6�#��=|0�M뢏?%d����zГO����O�	�q�6-,?	g�5F��:�E�k;��@�uOxxsd��\'�������'���')�m ��S}�U �^�[�-CD�'�S��c�4r�6����?I����Z��|��k֠OX��)r�ɀ����O���'2��D�w�0�����B��M6xA(�kM�"�x�
���4������b6�Ob�`�j� ��p�D�Ɓr�R����O���Ob�d�O1�,ʓEk�Int �THC� ���D�z��V��pڴ��'����?!�o�3�(�)��8V�J�y��R�?�z�ʸkش��$L&"ub������2R٢9�r��A���c�A;?���ry��'�r�'���'5"Z>�t�G1kB�@F	y[���D��M�� �?����?�I~Γ���w��骵�*�A��&�7 ���a�'�|����ƿ(ݛf5O� �w�Z�\C��؃g��r���5O��H7���?yn ���<�'�?��M��hᨡ���z��Ȏ
9���'��'��	��M�"C��?y��?yt Y*���!* �^<�4  ���'2��?�����*�x����Pz���w�.x���'�&y�l ���4-�����R�'��q�͹SA���CN�u������'p�'�b�'��>��Ɇ$ Ċ��Qh��P�4A�ɣ�MC�(Z-��d�Ħ-�?ͻt�PT�0��'m�~��n�&I�@Γ�?�)O�T�3�i���x�zl����ZT�7���i���ȱߕz6�İ­Ķ������O����O��D�O<��)8f��T�<|C�I�R ֒ ���F����5�2�'�"���'JJ��LޥQ�4y���v6��3�o�>������O�B�3��3<di��P
/D���.ׁTn�h@W��Umڹ]¢AO�yyr��E�� ���|��i*��ν#�2�'�r�'X�O��I3�MCc-��?�F�']GJU���Ƹv8���bnI9�?1��it�Ol�'�r�y�`��f[���/Ll�*8��c��j�L1�e�iH���!��u��ڟl���.���z-֡�F��	�L�$���Ot���O����O�7���O�({c/��aFڇāx�1�TH	��d�Ol�l�ƾ��'Y
7�&����,����	��0���1O���O>���f47�l���	7X+.�ؓhC�&+�DR��҅8k�jg)Y�<��"v�	Jy��d1m��r��V�g^y�����4�޴[H�S(O�į|��,��?r!
�����q��Ii~'�>q���?II>�O�����e��>:��cV`ʈ2�v%�,�I��J��i����|2爷�$�0��L9X\Uj ��*��bg*;����4�V��O��8�EBuLDh�Ȝ����B�e�?!u\���
Tr�
d�^�D���c&�)W����I�!�GҦ��'�����lr/O���%<��"��E0l ���f1O2���=Y�f�8u�(�g��	ޙc����'�&$��A��	؟��v��y7g��f�Aʵ*�ejP)�K�{3�'�ɧ�Oo����i�󄇁\�n�(��IVj�EI��͋?����鴰@�'%�'Y�	ɟ���+<]�uE�Iyx�0FX2b2���쟤�Iߟ0�'��7-I�v�����O��O�w�����⊩� ��a��D��,ìOv���O�O( �,�~M�=��N߫+K�yB7��{�Hݘ"(��$.W�S�#/�.Aş��E�Sn��I�%�@��ԟ�����x��矀E�d�'|��9%�ǺI�z|Sr
R�n�b� p�'��6�/KF���O��oj�Ӽs��ˠy!��s��a�#���<�������a�7-=?H9h��)� �9h���0�F\��j��?�$�(J>�)O����OX�D�Od���O��#F��.oD�I��\�c_�&��<��i]>���'�"�'���y*�DB9�g�c�$�A�d�7PN��?����S�'j.�8C�۷s����J� ��h��˘*e����'.��t.��|�e�|"^�
G��{�
E�,�qgS"!��L���������hy�u��B���OF�bs�U M�tq�IL�j�DEZ�O�O.<l�^��S��������0��<(,Ԑ`��S���T*R!��h��<m@~B�ȎLΌG�D C�8ĸ`Z�p����)B������;��q��ʄ�o�J�h�㟶���b�l�dXY6+G�*�9� �-4iHF�N15&X����>'�*3eԈxӄ��B"Ĺ@� Y���{�'�.�Q/�66�n�rLV�.p�\jF�;H�:�cn�#�<%�CdϨl]Mc5+�<"��Q�OQ�2X��*�D�1\ߊ}B�K�xK>Dңď(R�T8���.:\X`�eA!7f�8B�N�y�@�lsN�"ǈ&N4��x7�Ӥ-b�0)4��z8�k�C��Y�Nዦ�ճ_���'	"�'��s֎�>a(O �Ĺ�XB�o�>Y�X���Q2!lq�`n)�	b+�'���	џ��������c�8��	 '@�kM��4�?�F)�4e���EyR�'�ɧ5���a��{�m?ϴ<���G=���^�i�2�O�d�Ov�ı<�����#u獴Hp�H����X��	h��[O}�T���Iy��'���'Ң����U�\p<0��T.���9%h�3��'�b�'��U�T���K
ib́���F#�4`�fU�M�(O|��%�D�O~�d�^���I�vfh���)
�Dɂ+��dq듥?����?�+Ov�W�V�D�'wf��&@���Js�
�G���9��l���3���O�DWWf➨;!�9NR��$�������M���?�/O���e(�X�t�'s�O1�dQb�9	��<��nD t�r�Z�L:��O����
d�0�'`���e*R�X�9��@MϘ�lZRy�O����6�O���Oz��NQ}ZcT��
s.&���EHm�.���4�?I�+���b�	�L�t17w�,<ڔ�g���n�.[�6��O>���OP�i�X}�Y���gl�^椋��^`���^��M�4�Þ��'����Z/Cq�<�C��#��к1Ȕ�n<bLmޟ0��ڟ��e�G>��$�<9��~ҁ� @T�����M P`��F&��'^���y"�'A��'V0���QD���N��z�n�2��gӜ�$�y�Nd�'*�	ğ$�֘��8`1DB��B�Ѐv	� �\��n5zM>a��?Y���~�? ���p#[*mp�#4E^#��p�`�9i4�I`y"�'��'G2�'b�H�CA4)���0%�	0Ҥ1�
�:�'�R�'Y�H�qe������R�T��#� ��	�C��M�-O��$<���O���Ͳg��I�n�J$c���96j4��ޖ.�D��?Q��?Q,O|�I$ǛM�Ӹ#~��B�z�\˗��Z�T@�4�?�I>�(O�i�O��O30���ꍪh`�T�D�?a�t�ߴ�?a����8
��$>����?ט�EN��$I��_R:����2p��O���?�����<��`�Z�����|x��O<b&��okyR���7��|�d�'}�$%>?Q[Q�r�
A�.�F�Ҥ�<)ۛ6]�|�I۟��N|�J~nZ xI��*��C�D� M�K+<6--s�����O��D�O�ɻ<�OH�t!aϔ5k6�@YQ��;.^���>I��u���OH��F�n0����H��q1Rϐ�q~(6��O��d�Ozt*"��E�i>��Ie?�` ���	���83��ؑDeͦ���r�I9����p��u?�q�-�>L�f���7��+�0@o���i��Diy" �~��Ҍ�#Vd9(ND�`<i���-5��OD<�%��P���X�	Vy�-U�&�����G�}�x��DſN,�i`2A+���O��"��<�;4���K�Ő7R���G�	
���oZ՟��'��'a�Z�h�1c,��D�Q�'aesA�B Wn�a +F���d�O���-�D�<ͧ�?��dJ+��j��L&��!�սB��	��I���'%N �$�i��|�bQ��Ոc��1r�gA��lZ����'��_����|�������Y|�	A�:h��4���iK��' �0����J|�����n� �Q�ޝ2H��
��ԐW�|i%�x�'���'���yZw�V�I�
r%��������|�c�OT�䘃3v��O��d�O^�I�<�;c�.�r��e<�Dᵏ[0!�m��ԕ'#|���DH�7g�����;�TE��#��M�A���?y���?A��B(O��7g5@�b��1�r��σ�V�R	ӫO>qra�)§Gl@ ��oWg��Ĩ��J6�aE�iB�'���5��)jI�8��'��`� �����j���2g#H��O���~B���~�I-D���w�ֹ
eb�K"`�M���v#��2/OX�O��Oh!� �U58���$�[��Nu�&��Z�Ik�L��?q��?1-OL8�P	��f�X�P*e] )��Ǚ� $�L�����[y"�'����xe8`�6!�#�Ẑg��~w���'��I�����dyr�'�0�p�ߟ2�x��PFhYD��*���iu�'��O@�d�<I����qEH�Z`R�$JG �c�>	��?A�����n�4L%>QB%��ɱ��ޛ%������Mk��?q+O����|���S�Z����jZ���*Q�5@�7��O"���<I�O-y��O���5&�T�!>�*��<�r�Y��[;�ē����O���3�9O�NH�bҼ)B�o��k�<7���R�T�P����M�[?��I�?y��O���&�סMW�Y��,\� ����Ƽi��I埼�I<�ħ����y�:_#����B1��̳+x��8����O�D�<Q����?-�Pȿ�:����D�08�J̩���Z��b>u�ɲ$p���AAn������Qw^��ܴ�?1���?��L�'��IKy2�']����h��i@��T;�X=c���	��V�|�i��yʟ����O���-=�t�&�kb���GfU�D�j4n���Ё�iL�����<�����Ok�&2�Ѱ�#"U���g3�f�'�|�'���'	2�'B_���%���7Ŏ�С
�5&���B��:>�a�O�˓�?�+O����O���W-�txiƮ�?yΪ�����$�ı'<O���O���O��$�<q2��Jr�i��
�ZABb!ؕ&&h|��H9͛�Q���ITy��'I��'4�˜'f��nM*N�X �f�=?ߦ�)��v���d�O����O�ʓ9��P?�i���CI&8h�a�U,�@-x��#�`Ӵ�d�<a���?��,���?��'T�����N^�&Pc��L�
^���4�?A����$޽ ˄h�O���'���+�2�T5�$�6w��bEޣ$f*��?����?"�I�<9���?�%c��8�ز��#o�d4+r�f�҆�8�i���'�"�O_��Ӻk��
p�Й����3��H�"�ŦQ�I����Ph���Uy���^�nx�1�
�@Hj�8��'G�v͂�FkT7��O����O�iRj}rT���S!ű	v���QǄ`��1�I�M{��X�<a����8�ԟ��`��
�Rx�"��$ȶ����M���?�����#�P�x�'Or�O6):7��<J%�� S�=�lZ��i��W���۟��I�O*��?�z1�'>�@�9���7	�p*d�$�d
�����'i�̟��'hZc�ơ���ȃj�`\��j,��m��4�?�MF�<�-O"�$�O���<��C=��b�(&uR�̑	B�@�_��'�Y��	��I og(�y#D�DE���V1fܼ �%?���?���?�(O� q��H�|����}q�p���P�$i�&�T��}�'�X�x����P�	"@���60sfhB� ��_����ʳ\�&�#�OH���O8�ļ<qQG"G�S��lB� 0|��.Yj���(`_�k�$LI��i�r\�X�	ڟ��	�4���~���4-��I$�˵|lJ �R���M[���?�.O�����Z���'�"�O`҄�@�">=:��\1��B��>���?���XH��?A*O��;����,1���� �$@��7��<Ye�\~K���'���'C�D �>��UѬQI�`�)iJ*�`I�tŊ�n�����	?G�&����2�S����`��'@|U/E^p 7�]%��m�ß��Iܟ���.����<�ϒ�C~��P�k9���kr�������>�yҐ|B�	�Ot�i��\�P��� "OG&e��˦����D�ɞ
v"�{�O��?��'*�ū��"w�a�SV����(�4�?I,O�u�:O�S����Iܟ��CO���N�AS�&;ry ����M��w.�l*�T�\�'�bY�X�i��@$�F�gl�m�,	��n��v�`���DH�Y��$�O
�d�O��D�OP���� �/��P-��Ɂ;]�������\���ZyB�'���ڟ��Iş8�Y)\��E���u�8��%OSQ���z�'"�'�2�'�s��Pa���ꞌ,0���4n�]��!5�°�M�)O���<���?���9�*�͓Yuр�m�@�HEB��l�׳i!��'���'��I�SuR9����D���A�䣌% ӰUh�"�$:Xd	m�ؕ'2�'��b&�y��'���/F~�wJB'l�� �%�&��'��]�������I�O���⟜ɵ��	j`4K�d�-f&��4m y}�'R"�'2
p����?�8�j�[�t��˜~,��5�{�X�j,���iuB�'Zb�Oy��Ӻ��J�O�z�4g޳D�|p���PʦE�	����bp�8��ԟ\�	|�'���5������\�KsnylZD�$E�۴�?y��?���t��yyB��?����#O�0p2І]X� 6ξ��O��$�O��?�����n�C���)JI �����:ߴ�?���?AW��?.���Fy��'O�d����0(�_�蔱�aJ3Λ6�'"�'��m[���I�O>���O�c����+�����
>��!3�AIզ��I'��ڏ}��'�ɧ5��<$l�bGo�,$D���+�)���QX��<����?����(�2�%~1���.CA�d� ��~쓇?)K>���?��ŏ�n;Mjӥ[#LRq��F���<���?����$*q1ȸ�'R1�R��yJBqb���T���$� �	A�	ɟ�Iq��E��!f`�x��2$�LC-�U@\*�O����O
�Ĳ<�h��}a�O1^�;"���K��9�n�l�\5K�Ku�&�d5���O$�D�	q��;}�d[404`�N+k`� PUn��M���?i-O:th�-�X�S��T�S00���2��҉��9�b�P,}����M<y��?A`��3�?I>��O�ucP���;>�8"�F (�����4���(i6|LmZ%��i�O���T~�n�,}�(]1��P�\[h��mˈ�M���?�afK���' q��P�W�M/g��$�&�Ӂ�P��T�i`���U�����O ��:�'�T�I�*jL�AŬQ�-��Ar'�*Y|���4�����䓿�O��<�줊�J�g�X� � );p7��O@�d�O2X3e�n��?��'H�$r
X |�Q��nv�v��ܴ��x���S�4�'���'Ȃ��B 5��ieaS:'���5�r�j��V��a�>���������_���E�NΥD�Ȣ��g}��+ip�'�2�'l��?�F%��2n�+S�#���C�E۟JUr�%�d��f�'���]4O��ԣ��($BUHFN��Xc���'��	����	̟��Oa~,�6�*�s �*�\�H�a��`���gT�T�	r�'��	��\�.T�}�lc���������Ē��D�O��d�O����O����E�|z�W��j����ܐ��o��nS�@×�i��|��'��;��OZQ�r�� '��x�E Z�]���CõiL��'��	+�*�"��L���O���΁X������P� ��؋��M�Uu��n�y��?����Ʋ�R�F�T?:�2��R6Q�)�ҹiZ��'O`A�C�'s��'���Of�i��8�&�3�*��1�S>�0:�r�����<	�j^��ħ:��)@wl]v�\�䈚�@? �nZ+1���IӟD�'���Z�T�'�� ���6O֢5zE����A�� �>I�BT���O2���&k���Ŧ�.��5�׌s��7M�O����O�ccn�y�i>��	֟l�b�1�fа�I�V�t�*����'��u��yB�'��'k�S$�
�� �d_4c�괁avӄ���������O���O�|$�R (΂	=Xca���&\ͪ!�x2-ߐ��d�O��d�O�ʓm��A�I�$�5�Qi��d4��K�����'���' �'���'
�X� ��*3u(�y��O!N�Dp�t�� ��'��'bBW�PIbd����i[��u�1OL�>z�Ly��S����O��d(���O����H��I��Zl@�/�f���KЁ�?����?!���?�/OΈ(ь�X�ӿ<����7r���s�@�(L�����4�?aN>y���?9B�o�v
nZ��XJ���xSa	��h�lZ����	ty�Nʭ_
�����N��A�TbB����P�jb�t�D��D�����1?�T#<��OQ�����ޝ]Z^��ϐ+Dv&�ش��D�R�,,nZ����O���b~
� ���D"ƻ_TXz��D���Ҹi���'!p���)�S���=:u+]"�6B�/e��6M�j��oZ͟��I����Ӽ��'��e��F�Ģ�
@lO%>�n�0Am�2�Z��	Z���?�!���n��	�<vt�V)הC<���'��';�����'��O��䭟4&�5h$Ը� �x:���1���p�c�����,�ɰw�M�e�7�-	0�k���4�?9W ʴY�'�b�'�ɧ5�dņP[� L�v��m����������/�1O����O��D�<�L��^E��\([{�̣'�йL����&�xb�'���|r�'��nͦz!��k��.c츩F�G.q�v�y��'�rQ���	�1���Y��:� ��$�ްс�#H�En�֟����`$���'�� ���M3��8�U���u�h0���DF}b�'5��'&B�'���r"V>���9Bi��`�Ӝ�T��6C�gT�ܴ�?K>9���Cf��'NPI�eR�]#��[F��b����ܴ�?�����d�����%>5���?	�SJ��8>����b�6`�.0е��:�M���o[������i��HR%_�)�(��O�@`�Iڴ�?a��f��m���?(O�i�O���z�q��s�����
�Go|h �i�r^����<�S��  -��^d"-��
�k��$�������*p) �H@�xu��ӧA�0�B� 1�D]�V�K%-�`���D5}Dr��֠bن$r�D�zcl�s��G)�����N/1�4wG;i%F�21ɓ
�hА���"�� �*�:�|���X)�2H�H�*��H��8p� ��>���*)���,A	��)�f�¥�VL��[g@��hJ�����������^w;��'D�i�3+ژ�8�dP�h��YϛR̈́��3k��"ʵ��ǆq�>��F��S�'sr��Q�F!bi,�x��.Woɚ�b�����Z���E�(I��i���"�I�,�viB��<^��� �;$�2�c�O���'ړ��')�lyW���Ɍ�
aE�!�^��y�QB�$�y���.TXp�a/A���'��듔�d�\�L�'"!ˋk�:��DJ�~!�$�D1��',����'Q5��!.}��u� ����	��(y3sM�6,��I	􎚭zV����.c�n����ܳL�6��D�	����$?���K��0gd�<��ɖ���d�O��IU*-{G��[%�\�0O0����<��s�68��(T����܃?�������Ëz<��3�C��S�P�:P�Ҝ�yRR�T#fK-���ORʧV�	��g�t[��Ʌk�H������)����?9Vm�N_����h�1_���S��S>���	N*k���������҄"}�d(q���M�H�~"5�7_G�ɛQ�S�{��P6�C�D�t���'��>��	3SU�	�V �P���W�4J�VC�� ���*QOܔ*�4I�
�6<2��v�'� `WĄN�L�j�m[�=,�i���>)��?15�#o������?���?�;2��9�A	s�i�BA�T	<tQ����{�5�C�'�$fN�����Z�jй����dкS�)T+&����I	�|8u�'̜e+A�f�g�I6u��jA��4$K�E�\PTj�O�6����i>�F{BW4|%6�m|(��)�*�y�[>B����/�8"%��������C���)�<��� B�0��ؖkj=��ԩg����2Έ�?y���?��!����O���`>M��0s�|�4MV6w2"��ħ%@�axP�̅y���T�'Z��	@�&@WH���
E�p�ȴ�5D���!'H\5��ɐd�ЛU�2����#aRY�5c�O8-lZ��M#���'���7꼁��J.�����A
r� C�I"~�n8!e���E4BD�@�3&c��1�O�˓i��d�c�iT2�'�P�!AB�FNX�r��F�|x�'4be�w���'��ɚ�u1��pǞ|"HR)d7� �
ܩY�l�X����p<Ir�D�B�qO�Us�变�鈵 Tj���	˓1���I矸�����{�ڻ]��y+���R���C�fW{y��'��O>����z�������  V�]oc<��+�J�{բʣc������Kd�L`��hO?%�Wŏ�j�ԘP2��mP� sM9D����
U ��[�Bն?�T
�/7D�4IY������so����
G�!�$RCl��r¸#\���O�L!�$N�z-@���~R�)A3�:q<!�D�,���
��U&�h@Dǐ'/!�Ӽ[@� ��+�v0F�ڏn�!���i��lϲ)�������B!�Ě3I�� �J�L����_�!�� �ju"V�xٛD�X�W��<!"O�p�IM�@lfSR��<�d��r"O�ק��A�~`���Ѥcr�܁�"O6�c� �9���9u���P��k�"O�h�
ך\%�!B�*S��D��"O�r1�I,��
�>��A�W"O�٣��^�2�t����Ә��	X�"Oe�� ��u*P�R�� o~�"O� ��b�4�Mb�n�$���d"O� ˥�G8��kƲ�I��"O\�C�#�, �",�p'�X�"O��Q��X�'<��K՝y#��0�"O��
&l	,Z)���<Y���"Oh���] v����KX�&�����"O��ന!]����^%�-á"OVșu�I�f#��@���$�rA#�"O��Q��C�*X��Hp	�x�"��"OB@S �
1�d{wFͅ?�q�u"ObT���2��M�M6\�����"O"-$��IZ�� ʎs}�b�"O�Z� nh&����X!!�ɋ"O*p��-1��4*�� ��!�"O,��A�@�M�0�	S�����g"Ob�� ��D��1w��#O��Q"OVPC�ɍv�!Ój�\�D�3�"O�(㥍W�+}8�a'D��d�����"O�`X@�[{��ab\�2k*T�"O,��#B��Ul��SaF�W6"U"O&\�� ݙi�� QՁ�q
���#"OȑH&B��ow�P�H�2���)F"Od��C
� �	X@�F%jAz���"O�-���Tp3eA>L�� ��"O��ZC*H�W�$U#���-P�6�?D�L�g��	f����7��-cBH�)>D��
��Сo�0wQ�����FI
�',�����4}T����f�1s�0�	�'����æZ�7�<Xq�n Ry�p	�'������GB�yTm�/;Q�(S
�'<��Ն�.�M��Haq���P"OJ���גjn���
�1k_���"O4�ˠʚ##l.���zT�=�"O���S�-��XZ�1E<pY��"O� �b9_~=�d`�{�R�Yg"O�YA��%���*�`&l�T�)�"O�����,I�.�3o���,�"OhD��Qa+����C��"��C"O���5I�Hdpi-�2�p��"O
M����
2��h��Lۼ\�,�{�"O��Я��WB����fղ1��"O(Ȋ��D�Y���1щ�2^�b�"O.�$�$?��)C�/׵C��܉"O�Z�8ĠR��MF�4��"O�	�0��Xf�`;PcϺ� ,��"O��Y�꒩0� ��b��LU
�"Oe��d��&�Q� d�<��"O�z\��`�.\$I�(��F��y���^@�̊A@�Dt��A��*�y��-}�^�9W�А9d I�� ��y�*��$8��j6)>��w,���ybO2X�D��.ȡ9�D�C����?��Oŭ�<j�'�,<���8��!����Eoh���6��t��Z�B�/��9�䊗�|y0k�Ը�M��-�G\��<E��4,W�aI�ޕ[t�����
:ݞ��?Aç�1SP����dw�d�Gǯ7ʨ�5M�/" >�ɠ~�~�SB���p=� ��`J�3��ժ�U�3(�ǈ�9j	��y�8�0��^�fQ�#� �7\ԸT
��q5����5%Bc�8D��*� F˄Q[#�ߋ2��7�j�  4L�1��h!��>8#��(�"C�)��E�DP��Y��+o����ӋŪ�y�l_N��z��މt�����ӾNO�t㐣���JS&l����Y��M��E�v1�0�\�eu�h�bI?D�d���L�D�6\9r��_x�igi]X���I�bӵc�Ja���ΰ6�xR���Vܔ���	s����.'�0=aČ��f}��
�5���ð�.�@$���{��d��N�1�<C�I�K,�Hѷ/e�
�����0�O
�����7B�0պ�ʝ4=;p�P2��L�RY��+��y^4�T�E[��i�ި5�y�g@a��0���G_;l0����"{ PD+
�+�|����)���"�� 4��'D�A8���<D���F�{ӆ��CX�$�䰡2-ȳ/q@Y �
O�����5�&0��kF���x���nP��`�?fU8uş5dV��� J6�ɫ/���b�?mäKض&i�1�a�ހX(�D>O�4K��-w�xD�8er�`�!$����ԭ�4ǌ�RKBA� taQ�K�J 
�'z(0J".�����	�e�zJcb)z��Rc[LZ�x��k���v���µdF��L��)�S�>�1��Ie�p�3z�S,�F���Ԇ�
C)a{�ݸO	t��ĢI�A��Jw�I�.�،��H�.���H��4g��.� �(�+D�++¼)���M�Co�� �ʱ�f,�+?�;��H�'VHj�{��� o9v����Гy� y�eJ�a���0�k��/;<��I�wަ���[-�f��2�!�i>1���ɠf��a�Cb��Bl�@�1�<QM���'���E�a�
�kI�P�p�s6W&A�0�h$��4��о�pd�P� ���I�)g�8��oS*�i�'NJp�Ce�X&TA�"$~�<H;�{�捃ɟ0ACզ�,z���h�2�J�Cf�'. aU&�ق�� ��g�h�խd+B���%�?I�H-rr�']�AC���.��	-cF�)�E|�lIRL�'�f�?Y�GM���'���Q� �0��[C.��y�.����)�
�W&J�ud��c�088���I�,uC�G�4#���Y��9\�>�Aۜ�J�y��>S���o�>fp��f�W �r���N�FN�58L�i�wA(<��Z�1�$��fO�_��`	�t~"Cݾ(7���:(�T�4nS��?�v]��)�c��҈E�3.��x���h!��"�g	f!{�-_��.mI@"�8 ���Pj�7X���¶D�2b�-e!1�b�L��S#Ӳ:���" ޢl�T����.��H���2�y��^�WR��ƣ?��!3������ys-!	l=��g	c:�x���N}8�誖KB)&p����lhn�pJ��*9$�`g?Kb�ӧn�m|,�C#� �Ц�Oq�̀�ڬj:���v*�YU���o�l(<���!p����,�r����,��<#HNߟ )��Z�oA�ݪ��A��Ζ����X�R�Ih6D�,��@�A)Z2A+a|bR/
Q�XU�R	G�ȓ�b�6P�H�ahG#jAȼ���%�sw�$�#)�*W젩������ə-����w�BO�(�D�#8V�"<a ��s�X���瘥v$RT��qy/��4f��XʇfT�ɣ�E2 �
��[�%�}j�I�|�Z%�:��1#j�k�]��c�n�2��W��;s"�!�"��i�f��"�y�&61ODQ�u-��8P�����d�y�EEH<���?�������<�������3�ЈF��r�����G�;O�.ĘMm� ؆�_���x�d�JvDa|���2�!j܆v�r��DD��)�01��ȟ>UsvM�H>�����vL��!W���x��C�(������G&c�8��'\1�1Fx"ΐ�.���I�FXp!^����#\�4}�t�I�k���q#���g�\1�F×����BL?�p=��"�Cg ���a�jX�h��!;�"-2p*����휠v�D~Zc����)�(˂���,�>h{�'�(�KBU_���aRΓ?P���'�TD�� L=&e<�q!�I�Şw0f}р�52(�āY"IX�݆�,G�6pb�@627����-]0@n:��e�̔l-N��	]�/�ZN��4	�J��?����ܙWȡ �'>\H���d�1O>]J���$̜{�I��\�pȲu����B��AymJ�nM����>n��+0A�WQ�ԨVl�Ry��ɕ[g�9kƇ'�xy��Ϝ��\�qΏ�vq`}zfd��X����?�O��T����]�u@V�^a�3"nE^�yB��d���iń0���'��|Ѣ�v��Q��c>�Ls�y��V�.Mp�O4�����2��"�ӑ���.8��1���6S�����퉅n���3���D�a(�(#KM6�U
QT���i��%L6��2F�6�	'���}����)�- 2d�?���a������+	D��(˸qZ��\O���<�B�bz���7x���)@�1c��ԟ�;(���rd���z�����4s��D��S�NI�aP��jW-��'�R��Ŷi���RR�P�3؜CKM�a���H��e%d:��	q4������OΈ��*� d>��yR�b�? ����F��J5EJ�[��=�1�٬Jx*1�?��	N'�HO���(A�yK��:�A�h(�Q)W�'��\�DB�B�z�\�	��ج,�nZ�(��P+Sc��[x�(�O�&Z���*�cI�^�Tqh�O$��6f6ғq3
�ZV�����q��O�(����+�~,�+��6��m�򀄒:�!����2<��7�L����S�C�d���Z�G���	�>��S��>հ��Í��]J<�<�ǅ���=�D�ӏ{E ��WKi̓`�r|xR�ʂM�~��_�c�x
B&קG���
+1��z�F�$l�S�ПܱX��օW'��7�Ke��-nX�QR�ҋS���-����'ӛ^w�λe�� 2G-?�����b�ev��Y3]�"�?�'�^8�CV�vH�z��h�F䕓�d�9e�D���+�S�n�vyB�1Oz%��*Z,V(��7�U�g���lH�I��e�
�@Ld��n�6)!�1lU������Zȟh��Y1QC��S� 	)�����ft�4S�d> �'��P��-m��u�5@X��<�Ó,i�Q���AB����aW��(EX���1
��*�̞n����.�%)������P��%�&�ا�O���[��ȓ>f�ۀ픸BϘ��I�`�	�	1�0	a냗0�{�ϼ>��|��Ѫڏ�|GGėX}tpw"O�`�q+� ���(��ՙ,����� �Ud]�s��5�>E�T,	�z�0P�+�#5�,��C����yR	��z0���0�.+pp�`a�0<O��0��!�1�1OX�P�Jd�@0���1��p�bOY�Th�\�(����H��}P�Z�T�v�ˑ�"�O*!C#,ӒT|� pjE�=b��U����R��d�I̧j��i�)#�N����.�&�ȓiv-���6;\ru)��8;c���'����VN	�S�O�h�x�.K)F��YU�_h�Z Y�'���q��W��Ȼ� "�`ʏy�S~az��Ae�����$�FsNL�UjP�<�S*'\�L�ꖃ��b�h�Q�[B�<!Q��B���	���
sFFh�aoX{�<A*Y	j�>8�2,(m\Ej�B�n�<�W�1L�=�D*R=G(���-Lh�<�֩�V+R4 㐷{:���4EAf�<�s��~+h$1�� kl�2gE�^�<1垲,���I*�ɕ,Xq�<�Ў��\z��Bc�̨��io�<�%�	ajT+��8�0	�u��i�<�Z:.(���ei��%��B�h�<	���]jq�ٮ)���Ŧ�m�<)�n�
]�XhBE�Y�>� Kn�<У.jG�zvg�$^�� YR�W`�<A��בl٪Y�E�y����c�S�<�u�����0ū�C-� P���R�<9�H�'��� � ��N�kV��J�<YE&\)LM��솛G;�@֡�`�<�u'��g���k�K�p�l b��d�<au��
F�Z-�"����vE�0.�_�<9�NM�=$��KeM�='�!Ă�W�<�4���iN�QE+˄^ͮ��_�<1�A�-d+\�S���n��1�u���<Q� �L�V=뤯�"��4 �m�B�<��狛Q�����#��B�<��
�@�<�T�� f����Dt��l�c��}�<A��ӗK�,uQ�L�2k���CbJn�<9���1�t��h������2�k�<y�7G��xBPHٮ8��a�@i�<��ϙ"�������OR.�@��c�<�u�Z�m=���\I��h6��e�<��	�K�uRF���N���l^�<�ϯK����w
�b%�qSlX�<��o��IZA��R�jZ�U��B�	."�2�Ȥ�P�>�V�C`GS*�C�	N�"�*R�_+d�8�����B��/Y ��0E��pBP��6�DQ�C�	�+��Ν��ՙ���A�XB��:%r�k���;Oi&���!ða^HB�)� �l�a��z!���qsD"O�@��O GX4<�`ږ���Sf"O�I��O+9TpaAW!M� � M��"O���@\H��	�}۠u�!"O�9�`O�S��)��H4m�@�"O�e����l�hbaSU��"OL1��1>�� (�=�����"Ó�nB�|Z���� t��!HQ"O*�	,ؔ#��1ň1^"��"O�����0s���˼z]�]1"O25�.[c> 8DF�\l���1"O4��� �0��6hެ+c�y  "O(`��ʄ3NS�%ReV�oKTtH"O�9b�f��!K���,H��P�"OFYc6��D�HH�d߹P��4*e"O*��3M+>֐*"�ĶQ� |s�"O��"B�ZD	:N˥���;f"O&Y���en�:���g�^��V"O")k�I�z�:@�ѠF��8��"O���݇>�BP�@�˄%ٌ=��"O��J�a�%MjPp����E�C"O� �3�ºU�u��/Gs�je �"O<�a��H���3��}:�r�"O:}�W���EQ� ���,�PhT"O�xpE���X�*�
�(aՓ�"O�H�- �mT�=��R6Lp�� "O�6)�l�#�(�%�n��D"O�T�Чي�2i�F�B�]��@�"O�({�P'�T[�ژh�="O�L*5�ӘXp��:�"��c�D��"O��@D��<�e[�G�H�¬+�4OF��b��S@͆h���l_�a�!�䟰�,�af'G)��h�j+Qi!��M70Gv�;�G_+4��S�T_�!�$��|��]� �L�B ����)�!�d_�PJ��iW ��Q�.�B�3�!�d��F���c3c�p�2��"� �!�dK <�!DZ a��v�O84�!�$� ��uRf&S�y�3��=je�B��"f�rL8ì^�ı��oҥ6��B��p�z�6�!z��Ur3M�##�B��3p���v&��BO6&J�B䉲xT�=�1�.f��Ů>^�C��7�cd��[�X�� Ȝ&@N�C�I�I�Zp&��tR@j��z6zC�Ib���f�ZM�$�HGZ�S�zC䉦t���\�-�0؄��=vDC� &v�ʱ�Z w��B%*�8�!�Ù_(p�q�u�4 r� *{�!��M l(%j���hL�����?�!�$
�]V�hP���y��`�d��!��q��hC7��:�M��#$�!��W.�F(E�n�tr'�ې1o!�ٗ`h��BR ��9
���B�]�W!�d�)dlV��4 XC�P!�$³-�~�Xs�o$�F�^y�!�8^ne���M�� ��ԅÕG�!�D��Jh2���'�9N� ��g��J�!�E
3d�*e��h�r);�!�č��8`�䢄�*�hQa���8W�!�d�94l��-����[��L%�Py����I��G
P�T|��)߸�y���)Z��x�cV�Bd�ᒧ���y�F�H7Hl��&
�:�.��
��y
� :�z�KAj"P g��2����"O�}��L�?
�����Z�b�B�"O�逑	ߊi,d� !_ex�p"O`Aa�2`]�C�/�T�q�"O\���D
�$�9�Z(\D�H�"O����%l@�c!�S�s+~�"O��0BR
`ĆXa�Q#p ��$"O��q��M�~��5�_@À"O�l���?!_�$;{��+�"Od��fmZ�eN�<����
R���"OZ5*�ȏ%�^�`��	���D"O��1�Q�tdZ�R#t��%"O��ˏ/t��U�.A
O�.Q{7"O�q�j_�'���u��Z�9c"O�@h�@�ƪ\h�������"O�x�dMS�F��Sr�Y����"O>���� 8T ��Bb�:��"O�(����.R�9a!�{e)�"O<)Y��J�Dbc Øp �x*�"O��ZBN������%l9г"O�p1�F��f���I�� �e�R"O�����	l5�S��
.(�7"O�	�-ǢFQ���׭�7�&T�"O����J�+`2�
�,���B	p"O~���C46���ʋ-v ��`"OB�	����Z���KQ�k"O*<!�T�Lw��Y���-Y���%"O��:��ϻ/F���BK�4h�|� "O�0�Q� k'�ѓF���6����"O�� T�����Y 3�QzIa"O��zD�7h-�8؄lĀ"[�0"O
 �3&y%X��u��u5��1""Ot����FX����k�(|�p"O�m� H��ԺA�G]c T�3"O�9�2!%At��)�%^����"O4�ddOc���BI0G젅��"O I��@!i9��3�@�fl:���"O�9KЄQ�"�	bP�)T��q�"O�ѧQ�+�Je0����l��"Of���b� ��h5cC-�`��"OD�5��*,<^��$B�8���yT"O��Rth�|ȼ,6#%v@Pt"�"O؝8qS6c�N�z�ᓮ[2T"O�0a��w��ҡ��	H�Н�t}��)�'B�� ���ga�Q"U� >م�#����Sc$�U��LS�W�l�ȓ@�<��dHF1T��K��S�b��|�ȓP�H�s�MSb9���嗱8(���ȓWbA�4�BDª��G�8c���Gy2�|
c���b��H��A!+h��K3�u�<��.�,=϶�b��OƬQs���Y�<y�7G�r�ˬv� a�EL|�<11b(V��1	K�L�]���Z}�<y��ݷ	�y�T��=�:�A�L^N�<��N�6�J�՟u�0	 -Zb�<y'�u�� ���4�����Ea�<I4fE�9�����-V��	�0M�Y�<�r�N�,Θ �`�L�t]�h#+T���P�7�.�k����V����(D���t����\�Z�%{V����#D� ���Y5T���"
4���SA"D� �q瀉 ��p�*¹)I2�+�a$D�l�`c�PH�@�O^�\>DI6a>D�1�&_|L��]|�:��H<D�� �hc���5{Р�r 19���&��s����ᓻN��1QFc�=]�� 8D�D{��:�\��$aFNt
�s�(D�T��E�)?pɒ���.W }��(D�� #��.���"���PPU�+D�yO��AJ�jsOɂ(��JA4D�gⅥ ڄ9����w��Q�5D���CQ4!D`#&�F.Pb�ٴ	5D�Pk�Y��.죕�wL��(�j4D���p(�#]���'lB�,����V�%��-�S�'B�0x{�	�x!��I�O�b�$D~2�, ݒD��3�H�N�U1 B䉷eפq�$K� �Τ8�Cڵ)*�C�	V��4���	�Z����NՅ&C��/}�a�H�"U��,Aѽ���*O`�r�R� ��K�G*Hx4T�G"OP:���6�����M�UD 9q�"O��0 ���B�{2��u0i�g"O���CV Zva�-PL�B���"O@Y�r��}��8��ŬZ�I��"OtPٶ.����qR�� ��T(�"O\Yض/ūIT����R!z��Y0�"OT�*��
6!ULa�AY 	s8��"O�1Q�$����Q�"�0Kt"O�3��sztmKӏ�r�6��"O�$� ,Z\ջ���Gڴ�8�"O$��E��%y+�
�J��ʈB�"OTl����5~��AToW�@��"O��q��~鴄�P�J!s\���A"O��"C�*'�:X�b'Q,��"O@�Õjǯk?�I�ċ�4��q�"O�{F��&�LHPw.O�C^�R5"O�@�(%�p����.S_20�$"O���Pe� Q^)"M�=O`���"O��H ��Dnj�е�ʶ_J���"Oi# �j)��"��!!
����"O�10ը[�tn�	�
6N��q`"OT@�1�ʖF��Yڣk�cS�(�w"O�\���I�����J���HK�"O�t��,� H�t�S�Ɏ�/���"O �d�ʟ`�q{��N�9� "O"��k 8+�-! Ե!�͑c"O.�G�(��Ё�EV-5�B%k"O���!d�#c,�1�7yz����"O��:VG�5@V
�q�_ 8^xY�"O>l�G�+s�l�C!�5$VPUC""O����V�}�R�@��H�Tf�t@�"O�9��i�Q�d�E��7~O:3$"O�Y���������q�H��K�"O�L�t�|^�IR.�>S�YC"O�8z���/��m�F픚�Z ��"O8��a̗�t�R����&�˄"O|���EG.aH�\++�?�l��f"O u2um�i���FJGd�T
`"O� ��hZ*)A�1���O�E�j��c"O0p��
N4&�*d[���#��sw"O���H�4mQ�P:�(4\W�x�"O�4q�a_�u�l��D�"��Ӱ"Ox�1� ��3$0������NY�u"O�0x�P���v�S76���С"O�)	�		�ec��XFM���:9˥"Or ��A���̰6�4qoݹ2"O��r5�1�x�ѣ�wJ�`!"O�Qp���	�b�i8�
W"O� �M*�I,	�[�ˍ�lR�af"OJٹ&�K�y*���B
�\h�aA"O��2�A^�q~����q�4���"O�yj�,�:&��z�gCf���G"Od���#��}�E��O�-X=��{�"O�)Ɇ聋m{�`.՝6XU�"O�ay��]�p���խ��W+<�rR"O|��`�)5h���L�u
��"O0\Bp&��KMl�#S�?Xd�ZP"O���/W����!�#X6p�T�[ "O y�e�ҵ�2��@�!��
<EZ!�DZ�o/��R��U�TW��y���	2�!򄓭# ��@OK�1xe wv!�D��.���"'G�H���� �!��т4FpEXVb��a��}12��#E�!�$#m����V�z�Ź��:�!�D5�d�Q# /nkB�aO��!��3�Ա�Tl	i8))��F�P�!�d�xe�D@�a�8\&}����{!򤝓��qCJ��ID�X�/�";�!򤕧9����閧+��X��W(D3!�$T/�ƴJe)к!D�a�Ȇ)!�D�	>��}[���;��`�E=!�d�8
�$����%5"|�!�I;Z�!��(h6v�Pe �7!� ��	&{u!�d)3�H��Le�7*B!��_�C�p�At��Y�nA��1Oy!�$�{��)���?|�HK��[�v!���QT�I#v���~[��2�R�n!�d�?p���y��/\�����a�$�!��Y�!|^�Y���)}�	#4�^�L�!�W�	�^��s��1-[*)D��f�!�0w�|�y�c�_��S3�Q�!�Z�aJ�a��K�L�\qc��$!�D�gTa�[,2����/�w�!�$ѝlSX����,%�,,��kFQ!�$ �$b�7���iS>Ԉ�J�R�!��\!&��Э��wj�ТU�_�p�!�dU�,��P��*�&=M�=k�	�+j�!�,�H��O()3PQ��>K!�DB�_w�h	��H#{p�QfX�m!�$QlFz�م%�5wI�`��$��!��*I�ija%���6T��J��+�!�$ɉ_����S�*��<�B�[<+�!򄄧P�t���bģi�D�a�^�b:!�dT��z5����w��U�r,!�dV�3UN����+(Z&P5��2 !�$U�0�H3ٔ�2�p�^�@�!��*����(�/=|��B�=�!�V��	k��A*^� X%"�7l!�DՠU���P�#�d �f �%[!����`b���dJ�e��<�!��6��!��):������U�F?!�S3(�ЀZ��^�>��I��ƁT0!������Sw"Ƿx���ެ	~!���+/]T 0�I�N
�8��T�fk!�$P��4rV�Îz��U87��>^`!��%
K�@���6�h�mZ�w�!�����ؒ��T�%ޜ�q��8r!�d:n�L��H�6d*xFЩE~!�D�0z]9`��7Q�����2�!�!m�`�s�ˤx?xY�3�ӅH�!�DBY쌘D�J�>�:��r�@(Jz!�DK!�)�[�9�x��A?\�!�� ���/� +r��b�6��@�"O����7_c�i��1�j�"`"O�-�D1|��y)�d�7E6��25"O��+T�@L��$2j'�H�4"O�0�"���40 킧�����Р"O
!��$���(�9�$ͷ~/��V"O�ݪ%���z�2L8�I֢2:jP�s"O�$�d�[l�"|���&6H���"Ov���B��<5h�!�,��N"�ibc"O���7���eR���W���J�N93"O4��`fX=8�fZu�� e,T�"O��`4�5�*�sf����X�"O�d�r	ך0����9Q���7"O��B«�w�B1��	T�����"O��K2 �P�h�1@�\�c���'"On[v��"�B �v��o�4�	V"O&d���1�8��7D��I�"O0�2��͝-�0��ꉲq��Y;%"O�V�3�.���挦%�L�q��L�<I�ڠ4�H�bʤ&���0�c�I�<1 �3"��H���%�F(�F�<a��A�F(�J����k�=��C�V�<�ԁ �<��R��S��i3��~�<�Rßd���#��
D[���E�R�<F��(���a�-Ӿv���B��h�<	�Ɉ�@+�0�I9kn�m�b�<I��ӬBP��N�A0��se�_�<񄨚�p�f1@aL
G��d��Jr�<Ʉ`�EUb��wh�o�\�m�<��w��̓2��lݔkS��S�<��3Ҷ��aLΏ%;�2�)GU�<1���8G��*
\���
gO�<��JF�>���K�cn�$�{TN�S�<AS �P�$����b�AQIZ�<)��Z-[X��@DD�M\�AH�T�<��3zDi8���%���^L�<q"��B��t�6N �N�As��L�<��I��Fe.��Pm��y/H��玐F�<�s��1k����F�5J��ْ�Tm�<9D�eXHuc�i�1@�Db@��`�<�A
��uX�㓎��6���q�!FZ�<���j|*�gE1e�&�A�$�m�<1R�*�|���;��p� �O�<��Đ!�>�ZL���ʄ���K�<QQa͵oz��]4%�U�s�XK�<���A�e|��q�Kz8��+�D�<9��W7m>.x��GF�~� ��+ l�<Q��"��m�#���yDL�e�<��D��<<!ڣK�@���C1mU[�<	F�C9s��%N	S�±�@E|�<I!뜔DMc�Zw�v�� �q�<A1�ʇ({�����Ƀ-�F�@!#CU�<	$c�y0-��ѣ2�}�E�i�<�@�6�PY�W��!W-�ؐ�f�<��IP�z��k2�ظ40ft�%)�H�<�p�
�xR������P���Bx��'�6�2�M lZ���DO��F���'0 �`���	�1q��A�Ku<�J�'��ui�NZܾ� $g�Z8"!b�'F��-�7�RL���I�;m��s�'%9 ��_'}���.[6��s�'��[�oF�;��x
c��
(�<C�'��|�q/�F�:�R��(�H���'e�4�qBTbX�`����  
	��� ��� R�Jl\�4$�#w�~I�G"O��K��ɵ]��,��ʤ,�.�8e"O����L�m<<��/=,�"�"O��b5�ԩF����s�ɦX����"Onʷ�<[�Z JR/�-5"ORYb��	2BHy�+��Bx�"O\5���,?6�0�9�<`$"O��!�D�j��tIپ��`"O�ш�Ŧs�XL`&�'h-�"O�ĩ�F�'u�d!趥�t&��"O>u��ՙw1C�+�@�l3C"O�b��`+��P�Xt*iف"O���ծ��7�1!��!eZ�!	t��+�$*��D,
�rx�8�l�(6��Ȅȓwٮ�bs��tf��G�M�	�|)��&4x}ۇ!�$!6�BE*������E�^u��J��m�^łՅ@�sB��ȓT�j�����x䖔�0�߮XH��ȓ�L4
�jR�>$�cGn�%긄ȓ{�X����0��9�R'֞19���N��e�`[��ܥc%���N<��S��Ã#��h�r7a�:G�هȓ^���pq���)�"M���܏ln5�ȓ���µ@Η!-4��A���U���ȓYq|I8�����x��B̖eۘ��ȓ.�^m��%A2+h�h��J�;hY,��[��92J�o���0K�G����4=�pЄR6�ܱ� $L��\<�ȓ�bD2���2y���EN���G�Q����:]@�H�o֔Y����.�䃷kD�0��A�J3.l�ȓL��b���ʔ�f��(�x�ȓS(����S�c&X��@�8@L4��0
��/U���1����=������hO?y�bጯ[��� �MF	4��iu/P�<����a��;��_ �<ii.�d�<���)j�lY�N�B~<��Qk�<I��.&�~��(X
~�ޠ	���j�<9ᬂ�%i.�82 Â&Sd��T˚d�<���$\��'$��6< �b�<9�6C�e��K�_����Yi�<I���Wz2����|c�S�DA�<��/ ��2�<�L���{�<���K�(�lC�T���t��}�<�FQ^��p@���=	*q�<�a�տ*�������\�(��g��p�<a���q���rѠI R �dDj�<y�i��b@�\����Ǩ �F}�������H^4_�-�/�!aD �ȓ��sCeB>Cc�P��m��>� �ȓ|��aC��$fR���C���jGH��ȓ�d���ר>��{���V��܅�$�M)Ũ_��,4Kr+���ȓ!z�$�
�K�C�.�^�����G�JD:V��NdH��э�:q~���%��x��ٶ7�H�y���5�\Ԅ�2�88��S�F/:�S��).r������H�D o3"��ՠ�`ɘ��ȓ!�C��ׄT���I�1�H؇ȓN��)��
96��y�B�ԫ	e�ȓ����'�L!q�)�n�"59H���n~��2�`zR��>x�t���yR�q(X��E �,��7C&�y��U!����O��vrax��®�y
� N4�˅F�P�$B���+�"O<��a�q��r�E��<��M�"OVq�4@���XQE���x%"O�uR��@/���;3�]�L��"O�,�%�[( 	1��j�l�"O��A��_4,D�u���3hm�Ց"O�m�$G$BB3�V)H ��"OPAc�A��4ٞ�"��L1[���C�IT�OTV�"���f(�ʠl�lԳ�'̔-� �=z�Q0����} �q�'��5�@&�w�y� ��	)�4��'vl�C�AC�L�T�'�[�&����'���t��	\A��S� ��HK�'��L g%���q	G����i
�'U,�񦒓e��+�M
R& �	�'�f8�MR7D�![�Ȣ��p	�'�<�r���kx��I���8MV�Q	�'�z0� �Jx�!���+:�6Hy�'OJ�����V��]Q�E�.X���'��@K��)|��}�����*t��	�'�D�Q!�����P�W?-�ԌR�'kvE���\�1��myw�8�'�2� P'��R�l�V����<�O����ɉ�*��,����b�]S"Oܰ�bdV(7T�!��(��]��"O~�c��>�<E0u
˞k!�����D.LO��`c
�`�Ƒ�AID���.�y��9C��y1���:a�X�3���y��Z5D�R���K
 2]f*3 B���O0#~�����i�1!%�Q���S�<�� A0�ܡ �BC
�^t��md�<їN�Ov<����X�����^a�<�`!��#&��{�eג�^4�ш�ߟ����Q�D���%;~E���K�
���'�a~�K	6�C1��m��%IH��ybfY,��|�Q-��`�"lk���y#ؑt����h�?Q&:M�.�y�gJ)o���j	 P��H�����yRG	;|Dz'+xJ4��J��<���$G�R���sƠ�[��{a^�!�d�*�DH@��ٜ��\����}�!�����J�6�l��"B�!�D�o���x�k�
6�|pI���=8���$���i��&T P�,83��ى�yBf�eh��es�����Y��y���V�(%z#K�(�8Cb��yr斿.��|;ѭ��L51"���?�'bn��A�	�H�4�;e�,!�����'a�i��60��]�@�5F�*��'7B*�&�+`����ei�F�'�c�	I�(�n`Sa���1�| 	�'i0<X����t��a�a�@	�'̘9 �Dr�H�0(�3]����'5\�H��;�5����^1���?a/Oj牲&LT�{ffϟ[��(�2��9��C�	�˦�9��Й�\�#@�ưK��C�I�5;��	�@Dd)x��� ��C��/ ���ݸ\�8-���E�pi�C�;���1,��yPঁg�bC�	 D?�q�w�ҽL��Iy�8_B�AQ��iUd�"h��0�.Q,�tG{J?�j��ز��T��+ټ���� D��²�B�(2(TA#��-@�ڱO 4�QcǛvu
�'�)0zt�pßE�<� 6x e$Ʋ���(�ȏ*h���4"O�%ڃ[�4MV�"��:%�L���"O������5�v��%!K.R3�-�A�'���ҩ.��HÁ�#n�jth�#�q�!�X&9I�,Fz�Qp1PH���+�g?��7q��So^3*�JȘU!YS�<AVg��6{���E�f���ɔH��0=�4�	tNuz�F]�Q^dE02-T|�<Q&%ͮF��u�ïs��{g�Wu�<��J�]���hS"�k�
`��L�<y"$�d.�Ц ӡ!���EJFA�<��mʜm��L�0{���`�E{�<�TgҢ88�M �Z:?�DL!��v�<YT�1u�@óL?;�F�X��Yr�<�����*eHQi#BD6 t�����Em�<q�,���E-\�3�Hpbq�<aL�$�r�qG[�UuĹ�!Nh�<A7 �o�6�jpO�l,X�$mL���D{��i�
�����xb�1jա��;�C�I�3������S�|�p��/�:8�B�ɝ'��aE�;���]�y����F{J?ݺ��D:w�&���"#:l���'D���DcOX*v�7b�>D<��"D�d�w�_�O��I�CMR}��䀂�,D��T Əf�2	�e�flb�س,�O�B�I�1�00�7� ]�P�d_�s�TC�ɔW����/��)Z�@�#ɟ2^����)�I�T٢+"#R!DP�;�D����B�	pq�	s�7f����z�B�I�D"dl��W+.�ЁkH=�B䉔:�1���]�
�2 G~��B�/_o��a�cy�X05��O��!�$�|�O�1X�Ê�9d�1 �`\�Gۚ  ��G��	%k�BJ�y`TNR-C\�	(�n"D� h�I0��*�A�p����!D�`�Q,,hX ��ˍm�*�+�*D��Rl٭"����Ө�c� �G�'D�1F��8D��R"�I$F��H�w�'D�$Id��>)2N��'�C68���`Ch%D�`��Y0|�SA�G,I��pX�f�O��=E���O;�FL)�A�p52�ёd;]!��=\H��)#�r8���s�,�!�D�r���:@톣#-�x�D���$z!�K+�"I4Η�x@Պe`]��!��AF�`���M�{L\B7�ӛ@|!�d@9+�8�L�R��פHLy!�D�'���V���fx@!S�nh!�Y�pN���ˁ=LU�PFT7�!�$��;>< kѩѣt���1rO #1�!�D@�B$����2β�p�	2�!���!=v��� �t�HA�V�BI�!�D��i6d*�(��ε�A�i�!�d��� ��B�`���+�,H1�!��BH��3�ߌ��Z�[�!�d�k
��a�#�S��P%
Q�U$!��.AyB��У�*x��֎�9�!�,�H����\qV����s�!���Y4�26�_.Z�Z�/�!��
�6��9!f� [�4ad�ӻ/�!��m�!����0�,d�p�p�'��Z�'��~�\��.f,Z���'�����-���yr�[:���ʓj�]���1'�F}�3(H�B!���$���'�ª4Ή(�N�������S�? ��3�C@�� T�"��^D5�"O�)���
�<Ũ�[�"��H��"O64qA�c$�i�pa�1F�4 2"O"��ĺ]a�ĩr�6X�Jq���'�1O�%�c [��d
!�=`+�A�3"O�0�H�p�#ꌑI+�\��"O^�����U�g���q�2"OT�3d�$�*���U�t4��sU"O\ a�H���@�̖Q�����'���@&��ȓ�r����CI�kB�I�(�|�;P�Ȁl��#��- q�C�I�~���ITm��y��d�P��(T"B�	�L?n$ "	H&*���jd��Z���$&�n� ce�՝1E� A��ck�!j��<D��!�O�<�n����;KÈ��;D�X�3e� ��I5 �B���@0�3D��"�T�W�y�!e�J؂i�4�>D���(X�e%R�A1b��C��=D���pA� '�V����Y�3���e�/�Ob扄E����Abj9oE�:\���$%?Yw����D��N�,~�4�z�B
n�<U�_#]4-(�/y2���!�@�<�e�mO�,����Q�0�{ƪ��<	DE�^m�@R�� �Qq����B�y�<���M�c���Ls�L
�f
`�<9�k�((^����"Y�:3CQa�<�e&G�+:L���1"�6+Rka�<	vI�9(�>a��dD1��,���Of�<!d,�}��@ ׫o��A��h�<)'/ۆn��V/M/"fh��v��a�<i�lX<��XbK��\F>��a�W]�<Ap�K�d�Q�K�" <NX���O�<9B�;S��!�ϖ&���"�R�<a��f{��gi�X��*���P�<	�a�)���p��6H��SF�N�<�W�J�&4�u �����!�«�B�<9��3L?�m�@�L�^`s$t�<��0��x���x	\���Yl�<����D�ج"��ه[yhy8�L�g�<����8tB�Z�E�[/
8�ѧ�f�<�6��x�b�
H�cq�W�f���ϓ{��H��L%"Mnl���N~v�ȓcɘ��d�
���B�)wD���ȓ#�h@�H	��"s/ۦV��E���OP<lk0�U�oҌ �֢��B䉄OTb]�S���t����'iD�B䉦X�P���0O�<D�s̚�F�NC�	�Xbr�)�W�(}P��D�XC�PC���i�
�'ji��C2&� C�9c�D�z5��`�z�8����Gz!�ēr�n10��n��e���X�+T�{�|bOp���T#Pt�e s9�Ie�'��)�'��"t�✈Щՙ`V���'�A#�p��|Ң`\7\��ͨ"O�911/K�1�TA��h�� )D����5R/���% ��.��2�%D��	�& ����'.ض�"7�%D�$�F�o)���	�/���ڋn�!�Ĝ>z�q�&�[�[�lE2'a�$y!�۾T�R2���cN�Ј��o�!��!|,,ac#C�!n9.E��� R!�D�'����'�%���cƯf�!�$�"Z�:p�%�L�R������0A!�Ќ?��ԁ0�*V�`A��i�;!�� �TP%,�t86Q�f� ����"O��{Wډ`��0$g©T�h�p�"O�E�mɠILij�OzFd��"O\2k< b6�bcL�*gy��#A"O�5��c�/E�L\+�A��v]��y��V>=��h�ؕ��=�@@3��
��y�ʒ��f���́.�M:�ϊ��yb��H�(ԣ�b�z� �ã���<���䏳i��=Y�m��O�1�1��P���$O��R�U-����r-�|�q�"O���6Eݣ)#�t�u�8j�h0"O�峲͟�}7�hp�+Vht�]c���*�S��/Ud]�0cP�B��Q�0��n�!���}P
=�b�B�)�<]���U9j�!���|6�L���B��Pڵ�]!򤊿}��hP�>^�\Ȅ�xZ��)�'|���Pf"<��A�-��Zv�$��'�X-z�hF�X� ��R*$0��'=�A�����O�&�jaP M>2�ӈ��+�t`�6���a�H�Qj�)%8�<!�"O�XGƖ�%�<`"�h!k-vI9�"O�=��H� �N�t�@� ��؊"O�t�1-�N���!'�8 c���O>��ـ�v��%*�:`F�@��Y��!�d�=�Rq�s�'8Fl�p/��!�P��!o��T?��%.�(M�Iv���8�M�{Þ��h��h)e&D���l��M�Q�Q�FH���e#D���B�~���y�Â /I���Q�"D���H13vT���U��4-q7- D���"�M3\Q,��Q�F�)2��W
#D��0C�Q��*Q�K�l ���vF"D��@�g J���22
&M*����O�ʓ��S��{rˈ	>ꨴ	3K7�� �'�/�y���n;����'XD������y2�ܦj!,�yI	�,irMà��=�I>�D��ZO*����=�����"��y�ŞN�P9�B��d��@Af��y"ޭ4e�PYa�T�x�@Ѩ����<Ɏ�$�BNu07�,�� %cѺ_!�D΢iCn!���,�z4�a�*!�\�q��!�(X����M�y�ȓ&ʈ(B�Pz��L;`�!mhF�E{��O��0�W<&����">,Щ
�'�j�b�3n�"�L�5�VT�'�������L���PѢю?6�+�'!M����%� y;pdƔI�+	�'�5A�L;T��I	��D�rQ��'�p���	��C�"��S&�E�^1�'��X�-0;zQ���@�\��'U��kV��Av���jL�aq�'�"��:,��
ѫ]�}�D��'��J�+�t���a�|̀DS�����?v	`UpE#�)kh���Fw�<����;O@L���j��,��,D����S֭�U�[,ue���f+D���Q��D�J0�kZ�E�Έ�#(T� p0%�+f����6��$ZN�a˕"O�]���|*�q!��xų"O�%�@�&E��M����f~���"O\C�`ſ!'�%q]�^}�hb"Ol���A	�c�VMǡ@,ɘ��&"O��R�T�z���\�_�Ҩz0"O��
�ȓ!v®�)u���@c"\�3"O� `m�Fg_�'�v� ���'s �PC�"O�\r	��H�R@�n�S��y�"O$����s6(uq!�V�bXpI�$"O҈�PC6,��mQ4F*c9: �'+ �I��C��$X"�ߏ&+(�
�'X�vo�S���`˞��e 	�'�j�#'	3S���.�0d`܅ȓP(�2Gc��9p�1{�B�����N�����܅v��9 �(�
o.�ȓ0BB�j�`��@�$L�*��Vuh���gH�:U@�  Be]e���ȓ*�ʸJ�9� �����+�DA�ȓINR����J���񁎡[�"���n�8����֗w�|P��8��8�ȓ $J�У"�9l��F�Pb/�܄�~ZB����Lg���"G�Tpt�ȓ���(4�����-��0T�1��
��j��_� �3��@u�ȓ��mYԪ�H�� ��+Mp-�,���2�87�Z9"|Ң혽un���N<��5�ն_o��AF�ۀ}� |��*��u�Pb�'�*Y�"��NIj=��{�ԭ����&8��g�¯v�jl����Y�E4s�Y#"H�!�ꕄ�3f}�DH-�Ѳw�OQ��$��B��Ѳ���F;`�"�*"��ȇ�nЪaڼa�vѲ�`H(9�e��mt����B0��\b� �&D���Piv��C%�-.�~�2�gd�`L�ȓg�T-�2�X�F�p��k�2D�ȓaB�27j�i��]��A �F,��~�t;V
Ձ'�	�t��5�����J�)��%��|�e�Z+Y�ȓ#(�� e�/wdN��w�ۻ0G@܅ȓ"�ث�fųn8��o�9�����[�P���B]*�J���g�4=v|��ȓ@t�E¡�`�����,.�"���Dh\SF���Ļ����ΑG{��-
q��T�:-��'�8d�Xj��<a�;dOf�&/V:{J,�#A�y�<y'`
M��T���6L~�rQh�y�<�gI%��.��g�9V��t�<�6@ڙ#��R1y���@]n�<I��R�cby[��]cq���Ue�<�O,���7A
JQ䕻$o�a�'�?���Y= x	s��ު(�=�@)D�P �r�Q���\��@�%D�$��[�c�jP�@|Y��##D�h)�ݱ���wnǧ^xd�+��,D�`��X'e�P���$��$�%A7D�j�I�E���Q4�ڼP��k��'D�8���׫NZ�L��̉K�P++D���P�A3N8��
K41��� �(D��
��xjf]q�ݥ}�̀�'&D��L$T�.�C�V
��9s�/$D���vkV^ݘ���͒!_����H#D���r�[e0U���͠N�8��7��O"C�����	�-�y��R���qg�C�I�T	�(ƻ �n5�-P�h&��%kw��d�R+pԢq��?����~juc-ؐY�	T!5��3��W�<�!M;e�2�J�Ա[�hÊU�<�vf�r���җn��,����S�<q1�G�U���0~8� $`Y�<� Nq�ҎV�]�0=[�d�V2`�+�"Oę{#h��ɒ�Js�2
�����f>02�M�gP*��3"I�c�E��9D���t�Q/�yj�
I4��Y�7�5D��#A*��Q�P ��
8����'D�X���B#>�,�1� ����9�S*%D��IӼk�o�nEB���j�Ј��'��}��D���V�+q!U�]����'d�Б7�	�Kv�!ɕ*R�WW~ ��'hd�s�&� $̪@HQ>O�)�'v��YY-=ԁ90��^�L`��'�J�A��Þ�t� O�V�f�B
�'���xvoĽw�Hi��e�2P�20�	�'�\���}i d9Ө�g�(	�'��wN�S�B�ChB�`9��')����T�=$e��A�ʔ8��'>*`����=);d�3��
u��Y�'[>!�tJ�4��C�B�pX��
�'�l0@4/*���+D��?:A P0
�'���2O�l�@Q�iʩ9�t�p�'��쓦��+�P#D�/�.(�
�'7��j�(�	 	��)6,ϗ\����'�4U`�cR�b�-�%)�`;d5��'[�$g��#A�A[Lðo��`"	ϓ�Oj�-���@��'0��<c�nOZ�<	 O\�e��֮ h����]�<�dBH����'�6%0�# /V�<����)Tkȉx#K4F~p�v�Q�<q�L[�e�@���L	�t`RK�<���]�D��g��Y�EF^o�<���n��Y��C�g6f�QF��lD{��I�=Xr���A'�<���ϼ3tЙ����@�R�G/=Ȑ7�ƾ^�u8�'�ꬸb��WH�9������C
�'n����ȵf�E`��N�wgH�	�'�!h���-XH�#�;y0�X �'���p(�'������I]1+�'��=0�8+o��ҭ=F��P���ybY�iZ�`�By��R���yR(�J�����3mJ,�*�%���y�/�^�����̪t�4����=�y��S4\V���w��V18QIV��y�T�H0�����S�����*���yR(�J�L���]6x3�@K��y�M�?C��bn��n�f\jD�ē����$#Op��4'ՔJyP�s�(�
-�>�Z@"O��jvCǪz j�i9K�����"O|�;w��$l<
0�_�\�N���"Ob�ɒ�;\/��`� R	�(�2�"O�2@�Ď=G�1au K�Hs*0�"O< ��`B�xz���O�gεa�"OB�飭� 5�~�[�e�Uk����"Oرj�C�	�r��®�;y��x�"O�)�iJ�p	����L�57l��`�"O����̑猄���T^D�au"O0=��g�h���+~���t"O\,Q5J˶Mz���`��Z{�-��"O����ת#���C��.v�Ȗ�X>�Rr�� N�z��B�L�k����0ړ�0|�$M�4r]�YB��
:>m*��QU�<I7͝�؂�ha���DJǋ�T�<�f͈�T�T�6G�0��q�#Ax�<��#�H̊�b�#O	:�* 1 @@�<��@)Y�l�	ׅf�$�7�y�<� �A`��JF���/���K�"O���k>���΅;L��l"Odt뢭�J���H7���X���s"OB��!�y6V�1х�ql�8`"O�rBB�Lz�J1儵1��S"O�a�ש[!��G@� �赩D"O��"MI9H8$��5�� �p"O�u*���vM��[�j�zXc�"O�Hq�!Ei����r#�R���H�"O^�u�(
��i�a�Q��!�'"O2�i�(]=H�l졒�	�X���#�"Of�FnZ�<��PU�$o�H="O���� P8��(�gm��W��C"OT��_�%��H��ɉ��q�"OxT4�� \A�,�s�M�*��m{P[���'�ў�O;tq�PBm� x�&J5@��h �'�D�c��,W�P��&�	4���'��<Ѥ�A�x;Ҭ�C�(E�I{�'��)��:�t�B�Zh,j݋�'~�P���(D�����,�2X$"|�	�'���4�6�$�p�"TB�e��'*�Q2u��"6G�Cg*R+�@1�'=Nq1ť^�a8���b��5��"O�В��� P��׎fo���$"O���iT[�(�&�7Y�|�"Of�8h��$��A� a<X��"OvX��������E�N&�	P"O e��hEk<�Ҕښ� -y�"O �	W�Q�%	�����\�g�-��"O�=�C/6"X�)�A��U��a8"�'�!���0�֝Q�"ɖi���c�!�䚲{O���4�µ P��!��i�!�$Z2'���&�4��XH�.]�!�Ā�m$��s�O�Dvf=����Y�!�d��%m���v�U1i���CbϘm�BO��>4��$j7F3|~<���"Ot�HEe�%����vb9en�{6"O���ITW9��HW8a��q5"O:�1V�<\!�4G� Tj���"O��@��F�5G*��O�d���R"OZa4cٖq)��`���VG��w"OrTH�c��a��M��	+Y8�p�uU����ɼJ����p�j�@HW�įE˰C�I�R"ɅM"���D�$i���"O��a�&�W���ϙ,MxӔ"O�C�T;=B9�HN�FTl��"On�S�ċ)Il��3f�v	��;2"O�}r�ڸ�@����M�y�85��"O~�����$i,<в�#O�Ĉ�"O���v��6L�ܨ�BJ"`b�^�,����P��$�V�Ob(s��F�Q�zC�IT��P��-oX����|�6B��/;������6X������PBB���4%s�EJ=6asD�>|��C�I ;F��ZRp:�e�-qQ�8��"O����*r��0JP��!k����k�OJ։
S�Ʌ�yТхx��I8M>a����D+*$�!�E�*K6�Q���q3!�/X]��u�V� 7��i�.3!�DH�m�Xu�ɽB,�]�$�
�!��T�!,N9�D��P�z"NF�Bs!�D�xȪ��M4w��䑣f��^ȡ�܋A��C1��� 2�q�`@��>gnC� ��ay��\�^d���°@ꮑ��S�? H��ģ�&�m+b�րc�2���"O��i#���� 7��b�th�"OZ���E���KP�8�m�6"O� ��G�#o�`�f/�6���c"O�l/U��I��O�\D���B�y��*R�����M��X�C��y
�8-9��a��֫��2�H���'zppf�f`�kg�׮/~�y@�'��	�`�&D,�XȐ�*�
�'i:��Ь�)0�I�&b��
�'�Lt{c���du��Л5�z�	�'�jX�𫊃|��������lWZB�	. n�-sW �9&� L҇E��^�<B�	*4̀e�2��3N���1b��8�B�I�&q�	�4��$ be9&/<AC�I�Gݘ��F�_*���L3x��B䉘�<$�l�	9lXy�6�I�C��C�	5y�� 뇣J�Gp1p��1oxC䉷<��L1�g�N�*��L.t"B�.�d1cT��f�K�`��1��B䉲m�\��̄S%�܀"dɈm�bC�$m�I�r+Z�,MsbjA�2f~B�'2��R�!�F��^ر�
�'��i���l� H	�ĥ*#
�',�#��@&d�Hx85�ԡ�J��'9��*�["��4܀d���'�T+�j�u#�Hx�-�.u���'^�	���9B�F��lϫ�P�'�q��-�9s����d��'�����"Z�b�敐1JGN���'z
���na�MX ��	���K��y҃ɽ5�K�AOH9����yRM7ZuR�S�M��l��EV(�yK�'0&��܂̫�jB��yb�8.Bx���LF��=�L��y���7@���"��/�ޜs��y$�a������T1VS�=lē�y�c�7_��ЋG0P����Ҡ��y2	��+�� a��W���"�I.�y�ď��T����'��=b���yBMYy�1X�iȽ\E�h#��N��y2 �(Ei|tQE�B� i����yB�J/W�����������1���y�'� Ҙ����
� ����R��y���:L��!)��U��P@s	��y��Ɔ4N���ߢt�� PaK���y��h��p���<7vXP�0��/�y򦜮R|�h�i@,��s�����yȆ_�b��'ɜ�4e>(je�����R<R ��PR/:<�7�H�^��ȓ*s��LY�L�M���kLXD��z���.L����s��&D��t���X��Q���Wf���a\��U��%��s�'��2�����B;XU��(ψ`���	��]w.��g��هȓc��d�$��X�xs���$��5�ȓ>	��Xa�	bHT �W,��8�b��Ӱ@O�Hû��B݆�%��%*A:&� ����ц�!aj$��6��}x"#�>.8}�ȓU@���q ��0eT] ���7p�P%�ȓ-��hqR�[����&�Z)}�jl�ȓk����Hb=���1�
�#��P��=��p�F�A�{��ų�Q����S�? ZQK�*�.+����)cЀ�d"OJ��͂�Z�,I+S�Ѱ�J=b"O��:"���=��`�R�=5,U��"OPvK��n�Â�G;H�`u"O���3v��Y���+cR�D�"O�K1d��7���w-"�m�Q"O�@��^�z�h�� �o���$"Oz��sI�d+"�a��U~EB�"O�|i�"���lQ jC�)�d�"O��)e�o`v-Bj�q=l�s"O�(�G[6���#7
�bQ���"OL1����G�������3(���"O̬�t��>~༔s���8J����"O
`�˾c^�܈` �1�B͂1"OnaH,¯H>����lF x��"O�!�_	v����(լ�U��"O6���I';��ݰ@�T�<z���"O�59烑>4t�z"��W_�B "O*��FN�X;dH2-5.�y"O�	���@�EBlh�-Y-F-RѢ"O���e��Fn��Hu���$,��"O�AT�WT�x(��bltq `"O�hKs(Q�@�R�tB���	�"O���Ջ5fdNTxe�óG�x�T"O ����Z'���f��4~��1"O6< Ef	����BUlB4}rx��E*O(�0��\�ٱ�̟�0@T]z�'@�=[��-Aj)�g��T�Ź�'A�Hpk���MY��(����'>�HjE#U�ЩY&_6�:% �'�t��E%B_*J<2��R/�}X�'�v�rg.�;-��)�F�䮡#�'iȌ�6$����Bp�|�t��'+��b�JZ�+b�kw��=r:@��'��zq�X�)�9b�\�N먈��')�|�㉱Jh$�A��Q��)��'�f�hDJ]i)�|s��OX�Jm��'�`]���Ny�L@B�;c�`<B
�'s\\��.H�.����E笔�	�'�[�l�;nn���ݥ����'��I�V��&,�H뢂��T�tC�'^<Q3QK)z.|9�rcF�rm����'��$��%����+�#A�����'�(Es3�%��<�c�@\iA�'�$U���2������1��p��'H�Q�0�-:F7�, ���y�{����W�кfIا�$d��'UB�B'f�{E"P�@lY�~f��
�'��I�Wb ^Z�h�P���	�4Y�'�=�'��%������ �|,�'F ������HR�M�JP
e��'���㱥�6uN�j�h\�?��ŀ�'	�@���I{�݊�D@9�L��'���i lȣ&��8FcY�2%�ܢ�'C��#�Ď,'���K �J+(�hL��'�T��@`	>/$씊 ��� �*5q�'��A��Z�Jv��PM_��^|)�'��Y`M�-bcdԛp�"c��K�'|p�ď%s���Ѱ�)c� ���'��h %�P�脳�F
qH��ʓ-����� ��F�iJ��E1�4��0�3va�yIB#fK$^���ȓ?�ɀP�R�i `H�=����&�$@K#E��W��r)^�!5��S�? J��vbρbԜa,w�j��P"O�T"Co�1Wb�b�JX*'в�i�"O� ��h׮{6l����`rt"OP����6~���"+�D��"O�� �H��a�X!(�0��`��"O�UyW�X )<�RP'X�h��4:A"O�̺�GEv������4u"O���I�\��%$��lf(��"O(I�-M|4�ɔ��m�,��"Ob��VN@�6�6L������d"O���+�`eH��ä`8��"O��k�N·f>���cZ�:`X�
&"O�x灤|�d(�p�[=8�<��"O�y�aE	U�|�ɕ�-��9��"O@Lz�BO>-��R �B.U�l}�"O�)�%jс ��aS�MH ��c"O�l���F�]�ޘB��F�[�4CP*O��pdV�3֨I�QJ�g�!��'wB�XԪ
�d3��ڀkK�]"��3�'��K�K�
��%�W���R�����'�|Ɂo�6�B�bOfx�'�ȹ�sG�s׊Dr��ɡ�h� �'��l�p	/#&����-]��s	�'���KtI��x|�8��W�.5r	�'��H�I.P��-����7t���'�t�bs�P�d�,1c�~���'h�Qx�iLG�Z�'!H(���k�'*���ڗ,�`ݢ��_$f*���'�t���B	5� �z&��W�xt�'�L�n�$w�젲R�ׄLY�A��'|�t�sjFs���k���z ��'��@�U�	M'�)�V�B/ ��9�'�|\!�� ��$R&`)4z ��'/�H�QƜ#K��ez�)s�N��'������=ATp��HV�� �'�@]A0�C�RM2@��B�;~`��'��]��	IL�����0����'��ii��I�2��"��X�r
*1��'�HE�`�W9O�q�E���0�j�'�z��:���m2�2L�	�'�D�p�#Pv	P��v�J	�'J@x�p�V�>���sgԥt�����'-�T�s�Oj���F� � �V%�
�'H���H�x	f�����B
�'ڢ�Z�ᐢ#i�ʕ�=G�^t�	�'�lePv�B�(��q5m8BԲ�;	�'���8�aF�Yh���d�؇AA �{	�'ج�r��9}L�0���3y�a	�']����bV&[�y�Y.u�b���')�AJ;W����쁐f���X�'�b��K�SiD�˓�R��@�	�'z9!u�6j֐�H�(�	p�p��'<�=�ǭG&O��+0����I
�'BU�s�����aH�sX�	�'iT�)�C)
p��"f�#�h��	�'j�'��T`�����fdb	�'�Ĕ��J:�%���E�V���P	�'�"��oZ������ܖF]��Z�'�0�h�
�RK��`�
@��(���-�&`х#�;$-J��.8,^8)c"OD��E�_CN��S�L��JS���'�ў"~��,��逗!ڣVG���̂��yrD��J> t�%,�	J��9��F��y�*�<s���D�'l�D2�`P���xr� <��͊�4:��L �f�Z9��"O����S��i4�Ӱ7�qT"O0Y0ヿ&p�#�Â6.�U"O`i#"^
vnR�����>V�	e"O�cqfU }H�L�|HX�U"O��ذ$�>8��QcѥO�WcD�0B�I\�l���^���􂟶o��(rEE������ 	�K�:�D�D*�7'r��%\Oܑ�O�<XT
[��ʨ���T(b�T�R`�'#��`a�Y)�4�^�E����b�!D��9�)ɲd��%S`�\"M��:��=�D3�S�'RDh�?
���I�蓖μ�Fyb�'>z	�C��C~���b&�y�:e�y"�'� �k�����C��?�n ��4�Pxn	Y����gI�*$:����=��{���EM�26^�Jr
��r�3ۓ��'�$�HW��L�F)�@���T���'�V���88�tmi��	:�R	c
;}B�>E���
���"�Β(����q�āp^ �'��~r�Q�UD���$13Xӌ���� �yR�'[.`����5�n�cEO={��q�'̱ca�ǧw�bl�� �l��'5��öG�r5�}"��Z:oǰa�'ʉ2���=_,Q�d�	T�H@N<a�����*�܅���
�"�V��.G�!�DF`4 �2v��$�8 )�Q��Oj���1=���) .��o��p�WN:5���]��H��E��B� \9JE�A<�*i"OX�2��ϧ0�<���f_�P��pU�I��G{�O �U��@՜`Ӱ��EÒ!R@z`�'d9��hٓG�l��w��9J�6x8�'�r�b%�A�uW�8�w�R$"�3���z�}2�Ǆ�\�@��xQ�u��!��D8� �!������	� �Dy"�|�k�Mn50��Gv4e�`�;S�HB�I����DhŭS�y���".���=f�|���'�.�WJE�rȀ%���
LVZ�	�'Y.U��g0F��x��`ر[�x�i�y��)� B�x�rd�C�����5O_#O@B�	?
�-C�"՜E�������n`5�`O9t�'a`#}�'����:e)RNq0���'�"@�?.d�uJ�ǂ�� AV*��y�C�;b�B�;7H)~&HS� ���hO2��%>�'��JM�]�C�
�L���u�2D��B�&H0��d+�E�* J$�Raa/D��Oَlc�d e�V�u�*�2?����	h�`�N]]�|h���z��IZ؟�z֌��C~b���υz���a�;�IT��ħ	YPݸ�&p��C���[�	�ȓPP�k`"�L��QN͏KVP�Fy�!5���Ċ�q�"��5I=0*̒ ��-�1OP�'�Q?u�U !v��(P� Dh���8D��SN�d����!aԠF��2�N"\O�b��r�E�}\:5�4/R	F�Z rph>D���@NŁ ��Q@�P� �#�8<O�#<��a�0c�xA��G!�P���hOp�<���L�<�\IB	�=��u�ѴB�O�=�}bWj�R�&p+AƜ�Q�@�g�d�<a��H:p�68S 9� �-u�<A׌�<:��s�͐N��L��'��dF{���[���E۽\RL�Q+�:|3T!5D��9�)$*(��#���r_ �;2�%D�<��G�`�؈��-"�@I�<	��%*��]y�Y�F��8�AǦ�'�ɧ���� ��.�\�*E&L|�t"O���d7Lδ!(0 �ա�"O�p��KH,4�P�z4ٌ>^4��""O^�s��c�����zD�`yG�d2\O�1�A���f��(&����xb�XJ��
�@�|dm$ѶE�i�c8���ɜn�KfX�]n�!;R�N�3��O
��\�A�&�H׈[<;qly{v �(�!�dLL�α����"Z��  ��!��%8ڈ�񌂎C-�,����~&!�M!'��q��mB��w��0�!��ą+D��a�FƲ�\��a�!�d��G���b�@�R���e��(�!�$o���YO��Q��ű�À�X�!�Ði�j{rX�Y���	U���*�!��n�q�܄<ʼp��+��D-�O �R�  Tvq�F�G�Fj���g�']VO�txDm��s���cq+�=G�(��"O*\A%�;,����
��FFZl)Pቜ�HO�� ����Ȉ�$YR��o��B�9eGMY�C۫_����Þ�b��>�$iPH;���vl�g�Ժ��O#~�� �#��h`��3K���3�E�t�'tўʧ�J�a`�^?p�A �d߽v����	m�%H��ƅ /ٮ�Á�΅��u{!�)��<{I� �`�۲��,!vf�@�;��!��=1��a>��d�T�_d�U`U��<	��?Y�
^%q 8h��ԛY�(@�ĂT��4�<� -#�@���R
���y��h�?i���i*K�,��q�#%EP�<��c� 
&���Ņ,v:H"D�^O�h'��rGfĆT��Lqc!ު0�.t3e	$D�0�7+�3i���D	
	����!�y���|ra�="*�ti�B[�Yi�-�Ah<iJ(���f(�y�{2��&���a}bʡ<�K|2M?��g���d����"���eK�?LO���UK��K����>^�kb�1�d3�O��Ċ�;��a@v��:J,��"O��+c���qt�C=H�䭪�"O|d�T�E���i��(G:!�Z�v"O�H�A�/�.q��(W�Hy�|"c"O���6�Q]�bI��e�&2a� )��x"�)���]���� ��d�2�ɞ"��C�(.���'�L�Q�� 6g�V~��,��'ª���oX�">�+�M�J�'�0���� ����)�.p�р�߽�y��B1�z���#�lX)Ŭ_(�y��8~Q�%I���	�]�y)�?:����	A�������y� ���KE(�0|�.�d`I-�yBH�R<�#FΝ@Y$���9�'���s&a��8�Dd��Te��'ߚ����K�.k��b��)T����'r�iө�VAt�{��.I�
�'������/[�ʨk�G���Y	�'+6���e��iڱ�ɠB:(M
�'��up0�Q�,IV�ka��ImvL��'}����O�x�D����?,R�
�'��,��l�7
�JM{P�
6�B��	�')T)x҉H&F	6����W�~��9
�'o��Bn�3]%��C�X �)�'����ꉬh�C��	ːp��'���A��X�׮<�U���
ZT��'g�6<
�HP�\�y>Q ��� H9�F�
+D�pE3�-�q�`@�"OZU��%�D嬘y�:���H�"O���bX�Lu���©�a�|���"O���B"U��u�F�+gN��"O���H\&�H2�Eڸ&T�8��"O�=!)Ò!qB�'wl<U��"O��D��cL��RBj[�r��"Oܹ!���	|O�MنhՄs�V�z�"O ]bQFH�s�R9����V�dB�"O�91b��'O�Z6�N�a��@{�"O��L�91�h�K�^Eb%9"O�4Z`��(	s��CP�%!9�i�"O�ջ�MƯ�v��A"3] Pa��"O���Dj�$@S��3r$�P"O����G-C��p&���>p�[�"OfL(��J�!�\��f$u���"O�ؕ�
in���C�ѱm��DKB"Opܹ3���K�*����ˏTw�}	"O�pB_�V�ZaCK�f��2�i��,ˤ&�m���.91O*pb1�5wQ,�㵃�9YQ��H�"O�A����=GK6Ih`�7;�p���"O���b�[�lX6�00��%�I�S"OLH��ȸ� !+6�O7)����"O$0z4HO�+�r���d��"O�����9W�ȈKa�S9�2�"ON=�j�L�n�3�&6i����W"O��Z��ܔoΠj�䀑xЎ�"O��R��0,ƼB�C����"O��kc/X;��\	v�Z<�����"O@Ec���6	�d�G�Z5�q�2"O�����.L����p*�G��mS�"O H.m�fa��ܪBː���P��y���J�T��*!2$.9�`��;�y҂T��X��Б7k���Q�=�y2! c X��"D�~�8	�``�y�^X�m�1�=Y3.PJ�,%�yL�K��yI�O_�^ ��k�ċ$�yb�]��,l��̒;O��A{FL�)�y�`Ɓ1�� �!�2FvM��a_��y�AΖ��8�-�_)0�Ԧ_��y�ϒ?g`<���,Pܼ�"���#�y�':d ��-Q�$49Q���yB�ğ	(�H�[>��z�X?�y�l��e����+
�,l����y��ͩ�������ty4JE�y�o�)��L�Te"�lt����y��߇2�<p���J1b��;k�,�y"�Q?��X�J��:u`@Ҧ�y.��dH��@�?q���'/�y2C%�Rq��c�3!_��߼�y"�b��-��MO�h@�a�K�I!��]�L�E�1�L�J�e1bIU�^J!��D[��cO�m�L� '!��^�*��dMɒw0 @��n!�$� gR�`A@
�=|M��J�!�D	���{A�p;�B�O�!�DC40�B�� ��LL�����!�!�T�Gf����v���8�
7<�!���
<��֢R�u�P�@�c��7!���aV�H��Z�6�JL��%E o-!�٣V�VT:�H�%Z�8�r���Qa!��R�GՂ\��Y�$Q8�ǣ�)�!�dʳX���ޠ6@��z��!��u��Lh�/�K|t�BCK�92!�� ��с���^ƈ��$�&Wh8h�"O^��'���QPh��&������U"O���Ռʮ"�J��+	Id�s"O�}���t8Lъ�
P�d���"Oj%J��?aP![T'��c"O^���ȁ"� �Bb���1"O�	C���-�z�j�$w��y�#"O��2�F�=�.� 7�ӆ{���c"OPHB�ID�
���8&I�/r�@��s"O���V&�$���P'�0��"OBi0CA.�~a�!͊:ń@"O*Ȑ��`���{ܬ�	�Q"O�Й�H�r�8��&,�k���1P"OJY�� ��a�H"Q��2� u-�y"���F�!J��#����k���(@$��%��O?���y@|��'c�&$�`Rbf�.9�!���Sǐ�C�+z�;2�uC�$�:&��i�"W<�p=a����gt�D�҆j>ܘwE�z��h�F!zP��S���$Hơ!db &Zsʽ& �?@�Ɇ�@P:\���D%e���A���L�?�!ԛ,��\�C���,-�c ��#e�E*��ݺf����"O<��ce�^�6�;�P.n>I�1b�*?Z�x��.�<!�IH��~R �Y�<X;u
_�QTT�c���yR�^�w@�q�g�B����ˆ��?iW��>~��ˠD���'O�m@��~~2�]20u�H�ze�H��g����=�f�_v.K�3Gj�d�X�[G�M�$�˳R��I`�|2��2P��Y���y��<3�m�2�V�D�])5�V���'��̊�@]�|.v��0��@��z#40	p%��G84���g���aŪÒR&���I���r�݂-W�8	EK�54�	Aa+��5�R�<��'?#�<3 ʗ'JF�'|@��@�.��	�C��pi,�!�I|�ɲqk(�1���|B"�/	�)2��fȄ��R,ҏ�y�`!�(���,�&�'@�mS����Tbӄ-�Pq�J�uS��Y�h���^�(daM�5�@D��";޵Hq��ڦ����ťO� ��.ѨL��(�.N*���"S�&5��b��?���	�!49�1�)cy҂B(x��}�����4``�>S�%�)}����"��sL8@"�E52Ɛy��ژ(��1��%hN|sc`��]�)�'270Uc�B��c�6 ���C'��Fr�
���� v�S!,�Ɯ�DƖ�(�!qu���$=�"+�<��$U3@\�L~�=I�	J�I��X�W#FwL{g��xyb ]]��q`��E��)+NZ"��҄gj\uA2c� ���!b���?�2e@��5�O )[��x�a��]�yo�p�IU?f��'n�`�@�U>�J ,�#�E�G�O���d��#�ȬJsc�??ژ���m����>1��L�55�#<9�B	��"L#S���;��iO�R(���I40�@kqc�K��\��(��a*���. ��-�����07�0��7O��"��K��O?��ĩ�30�t���$[�V����/�9M���l��A��O׽��gܓ)�d����������/�L�'CJ�@�U�`D~"Eޭ΀B6ヷR3��t���s1*�kTa+b90l;ϓr5&�;�!)ai(=����?H�5�@��<[vHIJ��2�� � yv��i�h�KIZM�`$�wx�#�M@uE{�E��S,(��E]_�-���k�ϑ�rH��%D�JTV�OZ�F'�	Q���
�'IL�J�*M�o��H�-Ѥ\��� f���1�
&��S�O������:64���q"�L�t�9��q �X�$��x�F�9�RX���J�<�+�H�?��dB�(_@��O�#�p<�3#˦a!�eo�}�p����O1�d
&a1\O�0��Ҏ(���2r��+���c��ȣ	(0�a
�(��xR'�@0 �QrX��\��B���hOݡT�ЍKt�����h�9dv�d�1�@ f��z�&��~2g[� ���	�Ea�!RR���PX�{V�Q&:��I"$� �"�~�)��,F"N|�)��
�B���iE�!,�i��h��'h���F�9^ �m���I�P��O��ˆc�(X���!��\4�  �K�?�̟<��EF�
P�4�G�����Ӈ"O]�B��|��e�w+�T�"�R��Q�->��7o}�
�H��u�>�!+n웄II$3���"���!��ȇȓBZ���D6.�l�%�j��+���(~�TP���G�cW,��F(�~yR�2��Y%��9�I�@� ��8}� $;��&\O �ڱ$��̒��	�� \չ�bX�¼U 6���fP���Ԝ9*�I�@2�w�JL8��K­N�8q��kCN��'�e�V�1�IЦYKh\kr���cd��p��i�1D�l�S��=z�X�� �F�M�>eۓL	�5��ԫ�'#���C(w 5q��,(4&�"��ڼf�$�J�B�A��ْB#�!#��;L�*r( %a��y��Vi
�n�{�e�%M�7��ȓ R�� 
�$v��)�/˓zO,
 �^�LJ�G����d@b?�Ґ8N�<�We(?!��H9���W�S�gh}�6A�b��\�t�_�U�Ј݌&_�8���O*+�tjv$g`�2 	2j���2 {��cԀ�0<�gk� mਫ����,�$ PQ!�A�o
���, �Y�VPs�ݬ4���f��z&��[Gl��PK��G#H=H �G���UOĭ1D��<8�4وwG&}THA̜�AR$Ի�zBxh���$�ĥ$�>=�$��WT?��wK,���(�q9ڡ�����mqJ�*�'�hZ�#͡z��Ԑ����X1�xB5�&d9��w鋎���Z5�pJ�'lɋ����)��''I���`���xq��]}
D;ד5?VH�f��� @�IBSNy�d�(S���#j��C����>��W�S�4RǓH~N c�lM�(���6�<67��<�m�=50 ��T��2����؊����$>%��h���+xj��A�J�����{8����@x���H�
X�����
B\D̀0��d�Ѐ�@%)oҺ��%Č	72�OղE{(�	�ɊQ ̵zq�]�=���
�j1
��B�	�:;��C!X�90d�"� �Cy����Y�:�����)����><���O@�����>{r�	�+}��P��$P+G��9z��Է�azڞ�Z����*�[�J�[�[�2�����d�8!�1���áS���rc��[�D͆@�ra�e8������iƮZpl��ƃ�$l���i1�ɤm���B�	�K�|����h:�@�N|��Λ/���ƅ�K;]�eE�+䔙"�.bY<��ėb��	f��u�N��W�p�hf�fZlQ��E3*w�QE�?�����
dP����O�q3K�s{��
����[l�u��"O��7uˬ�R��A�}DF��3C�	QU2m'�K�@
��'�iq|  �>9�/����xP��*-y1	�V �� �S&��rt�'� P��f�0�5�4�ķV��	��K�n�	� ��wڠ-2Qȟ1�ҧε@*�0�Cf#񙟤���[�\��7b@�y�V����<A4�_� ��C�n�8a����D��­� �,>��GO \1��ԡb&ْ��]&0�x�YP��%�F	:��"`� 甋4g��j5C��i��aha��7u@�xF�Q<N�l���i�r��VbF4w�����6�N1HU��~*�[��\�+�~��ʂue�hJ�B�8�|�G�ɋN`�4�fiV�v4(|�Ca��yq���tF
æɲ��FE�S�+
�E��]ͺ���9R��
y�����OH�'�b�Ѓ�P�
/�h�w+J�"��7+���0�7*�Y�zlH��#m�n�l�D�O|�@��W�1��	>���`uˑ��P�=s�4��+Y��x��I �䜛�aƟTZh���Ή 1��q��T�8L@5�4J�-~j^����io��Z6�Ihx�hX3d׽k��@�h�`�Otٳ��K.��G�=��O��O�͛���6:�����a�@y�'R�Y����}�vl��!<J�lE[��ֆu�H���Gv<a��ʸ:�����ř?�N� ��e�'����+YVV��|*Ҫ.�LFάv����Q+j�<��`IZ���#�+<#���@�s?���\�ZkV�1�=}��Iɤ$ L�S4.��7��M2��k�!���~����F���	�#�Ot�'�
Q3CG� ��x�m�=���jŀH�h�� C ���?1�-��<9��  JV�)n廦��9u2$��9$�d��-�'�|��6���r�2��F&%D�IU��)d�t��o;�	8G#D��Zs�д*:�9��wP����:D�|yaJE'n����$O�@:��R%D������]�pM{S�,^#�`��)D�,�Wk[�QB�@���W���p�I8D�H3` ӆ[��Uؒ"�%W���"&�8D��'���-:�+&�Ȥ\6�t�%M7D�dJ�@2���Z�g�"U�$�T	3D�P3��}4�p�7S�<0�(��3D��s@ʃDP�X�w쐘1n�)iD�+D��;E��u{2�B����cl��!C�"D�P�lͽ�,��"��<� �Y��?D�ئ�[�L���)-P���?D��y뀎)�.�(�L]W��[!D��)A��f)�	��OWrc� �h!D�� 
�7摚��Ŋb,>���1�"O:E{3fH�����Ɛ�?����a"O�,"Jۿ&XH;�%���Ft�"O.���aǢd� ����]��Xĩ�"O��EJA/\����l�39�x�7"O��� �Z-0.���&�T�t�1c"O����@F�#��K@ϥ(�j 9�"O�B���q�<a�Β�+�|�yU"O�	i"�L#���`tBդ!���r�"OV�S��\��-�`�A[�"1�"Ov���B�26nLK4!�1����$"O|�'!MĜ��T2}���Xe"O\� �!�)"��E1��ܼn��T�"OV�
�m�j�N%dHʖydh�"OP�ڃcI�<�LM&�c2���7"O�ţF�=�����&6-�s"O2�$ �m����&H*3����"O�D@���PX�fO�-HU�f"O2�@�˛�!.��#�)~��"OҠh��зq�� 5��q����"O���u�>S�4l"��� L�6��'"O�u�N�^�\u���'El�ab"O���M/6�ΰ����jD��Y"O�a;�@R�5f��Ip�</�*4�d"O(�UF��G��L��aX.�"l:1"Ony�E�w�N�jP���X�ֱ�"O��0@
H�pt;Tϝ���Q"On���+�����	��*YP�"O�	��/WR��P�A�/�	P'"O����
O��q`C�ED"O�
��/��d�4Xl��*"OB���ɝ�"ٺ���A�8�\��"O:� 5�ެI����&IP�f���"O\�)ȪJ���#{��Xc "O���KX$2T���%�(�zt�G"O��r (	*H�عظG����¯3D�أ��	v)�bj�|�:x#�%D�<{@�qS���F�0���G" D�L3@��%���h�m���y�j*D�̣�hW-E��0s�E�;p�"D��J��[)M�����C�uQ��E4D��֭V�Ey�싞_�I��6D����bdx�bէ9�D��7D�8p�d��rm0�*� jnt	��)D����T(G:���� ,OV��i&D��q�N5ۮ�Jc���X�A� D�$���[���= �Ъ]O =#0@:D�@{�
ǈ gLyPl��m�*��3L9D�Hᇎטf��at F�%7 !�v/6D��*p�/`ϔ(ʄ�ű@Z顥n;D�,y��2aBf�k�K�7Mȼ���%D���k�g��Q�퀂Mg�h"'#D��؅�]��*,�q/_0G��$��2D�<�VGO��b�btk�$�H��Fi.D��"d��&�d��!�X GE8D��Ӣ�f�����JC��*�4D��V)
�h�t��,ĥ8��2D���2F[)T�N�j��4�ȁB�<D�ܩP���u(�Ÿ��W![����`'D�(e��"Rؠ����U���5 +;D�<���]!t�r�{�h��h�8p�'D��� �V�UK�9�g��)���A$D�����ݼh	���aHR:
֤s�A6D�Թ��3����Vm�	�X�6�5D�� F�f`��L�\���;XDz�"O�`3���'����䌜2dNiy�"Oz<8�$D�=�0�!MM�/h�Z�"O��z�M�-jL� -� 8��� 0"Ox��SB��YW�D�#�ܽ;�Xpq4"O�H�p���2x(dkW�r��ԛ�"OH��5������(+�Z�["O��Q�'Љ��|�u
=FT<%��"OL��F�:9�l)�
��x�����"O��SBP�0��@�&I�ٰ�Ir"O�M����"p�	S�H�P$����"O�������k��q��-�H+@��'"Ob(���#j�=ൎƑt/���"Oډ	�m�(���3aʞ�L �"Oh�T%�T����5ƅk��=�5"O�I0���F�ArGE��o�
�x�"ONy�@cU8UN1��⟹$��mg"O(Q�@d~h��7͎N��i 6"O\0�ʞ[[��AT�̔$E���� b������Z�)�矸[�H?~����iݔV'zk�`%D���S�g��\� %Z0�1���v�0jV��W��p�'v��PĠ��7� ��s���v�(��>U` RlB�^p��X�9X��q���+-�����<�y�!LHUK�jF $�̼�f��'���1�)�G8�����S=�@��Do�+���c�M)�FC�	+K~^�)pF�87T�	 f�`��Dg��k̨�#�<����O&p�dƇy��B�P�GJ*�"O�(�3�ӟ��mK�鐸,2R���'�2�9q�52�����K��q��O]���:p��H�\4ȩ����Ctff�[�� o�6����U$2s"9�)ֶ�D��N>1੖7�L��|�<�f��mZh��g%O� .^�7(XJ�6�
%��W�Ҹ�:I~BmV<"nI	��j>�İ E�.��Ub9R��R������'2Ш,j�DJ�,�$�J��i|h2]���S�xø�iP��5(��W���0ǉ.g���HG��[hM{Ŏ!����YlEk��L> �˩O���ȬNn��1EL��<������FJ�Q�� 4���V �('u(�5˩��EҐ��<&�=['�(SQ����4zH�k�$n�Z���\�=�A+"ϭ}*Jp��~�PX�L�b@ �Ԑc��kB�5�<Y�#�B��B���K�<B����?�Í!��P�C��n���w��F��D@��\�v90��vL͂x�hu1�*J���
��}g�*v_j�b!�LN��?9����N��]���%�iC�K�b�Rb&�a��Ɋ�j["��\��`�!_%-f�]%?㞰��	3��Ī5
��Rd)C��<I2V�_Q�b��,}��d)ձ@�s��F�$4�$�� �4&|t����@ux�cb�'�$ Q��Ѓ\�H�q��/T?:���|���V:0���'4���
�Q`�z-OԤ �l\� �BG#�7V��w�0�"��=�	4�}.D���b��:��ђ�X�8bbd���� �#��(Œ��S��vy��� `�tJ��Y�$9���	��$�H�.���G*��qw�,�we�\[`:2H^�_<�('ǩ<9�IH�z�r@�L~�=I�ᕌN��,x�⟂+� 1�p��iy��E�|�@2���a�'�4�����l�����x���B�g�OQRpA� ����<Qҧ�J[FPq��Z�\ҾP� (�K�$�:aIֶO\��?�郢8��$�$?�	�=Z��3�̥~����c�d�'�xYҢ��Sc���~"A�C9Q��X qo�;��!FdQb��^,u.*�",H"�0|J�l��0�����	�8qG��,�	&2���k��8:s�S�O�Pyp)՟E<�1N�")Fz!���"+NRq��x�P�b��@Rg�5h0&��e����ݼܸ������p<!�b�2��
�f�aa�px�
V>9/�8�a/\O���O�i�Hz��L�}LX�'��"1D$㥌���x���e�P�Z�&��S�@Z�����hOt5�d�����A���y]�}p �R���[���~B�����m��]�q@B�ZV��%Mצ"�x�5.��!�]�)����/O@��x��+�t0 /� �2�����	�����6y
� �!��m`���x~1�Oj���I�4�Z��Ϡ9()ā��L�O�D��f�A���0PAB8�̽*��� �0��9>����uN�7zUXL��f�L;츣Co_�\�u��;k�>��B�kU��\,EH��䤕��A�ː�H�Q�~�h$/T�� �>��k��V�D�LIa@�py���Z7�'��b���0b��e��SH@��&J9\OF�2᧕ꨡj��
'?ςl�
�1W�:�� �
BD+p��7��$c5�D0:OjH��nT�_����N�v�J�ɒ�d�]/�T)�Ã�w����/�!���f���E�+`^���I��`�rᲁ �^j����<"D�K��"t�|�薊� W�&����q$.=g*V�k��p�R�< L�G�� p�t���<�;	6��&�̑8>`�g�ʺa�\C�I k��Ó�L�1w
����w"��f�=;`�dC�����d�Ha���)�f�8J�`���e�+��q�f
Lj48g<\O��r�A҅3��b�w���x��#�F0'�������~�N,8�	���w�CBeE�6F���@�(.�|\�a�6�Ih;"�6�X+.�!@�O���	ǰYɈ`9�h�)hg$�B�A�emn���]'P�(���'���(�`�?rfY��I�_)$�uH�0��3'F�$��P�	�_���3 O=wnIʨ���HN<i� ��(}`�*��r����l����Q5� ��gFY>N���� QI�g퐛za���DZ��it�_4@i�A����	��	/��	:��)-6aY�%D�h�Fi�*?Cr�3CoÀN�+Q�$�^�"�<Bw�2O>0#�B-k��p5I�0t\����':8b[�BN��'��U�����ʴ0�1 4�T�Hs0��RO�Q��P�@:D �5�z�aԨR�Xt]�H�TAՐ8R���Ƙr߰���2D�@P�
S'tݾxk� (����2�I�)
���GR��OQP!�o��|*�Ѯk~��a�8�Ѐ �.�g<!��/u���0��@�������T	~	�8*�	ɍ@�
�'�`1�N������d�"l ��Q�S�
4&�+|џ��c��L
4�;���_zs�x��9r�	��+��)�����'��<����I�DH酎��l�%
�l��4<��gξy@6h��"���'̐q����cI���'O ��M�5	��)��ų"?���'Y.�bt���j�A�1NQ����ĥ"}�"6��
�	��s�>��$/��;��>N1*qkW�K�)��CDy������=e�h� �B
� x�pH�噀j*�KFI�
a)��'�H0Wl���X��	�$�����#!�6���L4u�˓@����`* }r�\?z�9��!�@�3��@z񉎦	"ȑ��Q6�X�-���t��'�K�@%�tdϩ���Ȑ�Py��S9�^
f�iu�IMC��n�0����Sg�LZh������C�
<�~R�B�P`�P��b�U=V�#��/%���Y�� j/B�'���˃�i_Lc�>A���68����L���iN����跊Xnla���ə>��<[�
�|���ɦa2�ҦYl�xJ�$
$���@S��U��-��\�A�$�Y�(�ChĠrM(h�d&S�V������C2J$5��lH��>!���Od0c>-��*ud���B����-l�\�����>�1��Fm�8@%Z�7#^Y	Ǣ�]��
55e^�Ҳn��0<9@Gܷ\�2س�l^�2v T��B�����wӘ4��yd���J�>PLt ����|(!�D�=k@��W`�� b"BL�$�Q�ԓf�P=fpZ ��ѓ`�J�V����*��'���y2�G?h�H(�,˰B�T�p�K� �~0e^�	2�*�S���r��$���Z4S4$����. �B�$dRP��`PRZRw���TO�(�ND{H��I�}5|�ZF�:#fP���H��"HɄ|7lѕ��,+�4r�HǠ/Ǽ!����VH<��¤M�ځ��}�(K���Y�<1�
�9H����"j�4�pΞx�<i��a-�����Y�/u����z�<�
�a��i�PM���N{�<1& �
��Ds�>I�Xy��|�<Qd��evqa��,
va$e�|�<9��62و�aE�èT�@�$Uy�<Y���v��P0��N_n	�3,�r�<�Fi�=F��,��W�Z&�zud�z�<�T��e>�̓k����2A��x�<9R��<ʜ�ӡ�ْ�@���u�<�Rh�E�������PE����� s�<� &p�F��#�E@6]�x�h��"O%�i���B��!c��(J"O� 	� Y:�!�QeڔbN��&"O~Q����t-�u�ȑZH5�t"O�̊�K[Y�n�s��2}da"O��2��4\�4E酧�6[f�x�"O�;ҥʺSu ]��LB�rCT��"O0�SF]vﶁ��KN(^��A�E"O|LX��IѸ�*��O}��#�"O��j��\O����ٶWaDX��"O��pR� /�h�2B/MQ6J0"O���$��T&\�s$b'����"O�sݣF:�$`ߒ��XR"Od��%�ͧ'6��	`�Z�h��4X "Oh��UJ�<n> �`V-�!{�,���"O��D"��mB�"�$\�@��e"O����^>Ċ��;rl�H�"O�APӬ��.�:��Z1e����"O�@[5��QA�&)��:X�-p"O�|*B��E@��Pn=M�ڑё"O�x�F�N�pҔ�Y�����"O�q��KG-Vӂ �V���j��з"Oh�󪛩��$����1:��TI"Oء�Ņ�}��r&m�jH!�&"Ob1���%_7��Hҭ[�p��Y�"O���c�DQ���I�L�(y�G"OJa1�OM&�
0k�I�5������"2��!�BՕ��X��H�0�1O�h��	�)4�49��,.�L���"O"��ӇD�b�]@��M�P�"���"O�ũ6h��e�PmJ�_���"O�����{��pW��%���S"O�0�+
���) I	T���W"O�I"f��-f�[�	LTd��`�"O��`�.�1M����X�r�jL���I�t��m���)�Y�L�P���o�D��s�_��pM����O��S�rJ<a04
�� x��H��# ��%��@��W� ��!��Iݞ[$V�s`��>����������	^�����Jc�	��(�`]��MЅz�%�%Ě�@�Jͻq��YP�g2]C������H�@��4��cϽ[0�V,�4��Pk�Ky�q>�A�ȿD��R�C��K��I{���T˂�C,O,��7͝2�0|ʅ�C�6��mÀ!Z�J��4¶+�(\9�Ih(QS�(�.�Q>���i�	F�+g�MK���;)��RDNж_�b0�bf�4Dl�d�b>xր	�a��C�M�l �БJ�g���
 �<� �����	�)b�q�'�$\h�bU��"x�16O�H�姆�VD\)���O�jm����-g��0BB��#e��'��z�/J3 $f�3B&K!�0|b�!�.2[���c��3ܾ�h�g���*���>w�8��[Oy��)��I#z��A�U��� ��.<���$�W
�5P�_�h��2�t8�����H�Ahk�O-)�nǃ~	�����Z&�$}��0�S�S>�ʝ��S�{��I��!W� �s����3m�<P�
��`�OC"\�A-��Ɇx���(6k��b�}2���)��O��>16}���+C/X�`"�(%���(O�����d�GY��AF+E|�*�"O����Jb� 1ғ�/O�4�
f"Oj<��M�h48�v���1��x+#"O�D ��*�$y����9O��W"O�4)�8�j��A�1Qo�|�a"O��*w��>�(��pʌ�w��ј5"O�PS��
�=Ӧ��vi2Q��9W"O�1 ���bΈ�����+=n�r�"O�#�G>F�
�yQ��)o�]�"Oj�
��W6��q��f��0��"O��j�ݸ+�zĨClD�/D$�Pa"O0]c�B�R� �uKԡ"��iF"OT���#	,��W��A����"O� ���$��%7R�"�X2j����"O(<��¾rօ�G�$F
��"O�Ɂܚv�H��8M.Vyz4"O\	�2a_)K�P�ٴ��1{����"O��;4�G{Db�!�
��qS��ґ"O>\��D��]���0h�6:s�c�"OfH+��>]!�E�&S�o@�u��"Ol�BC��Y���+�Gʏ7��Z�"OF12���|rl�
X�쩷"OZaRt�ƶ*PE��fN;�Nh"O$�)�C8+8`1�@ʤ�^a@r"O�@���zp�]��-����"On��B��B�V�y5��*xæ��0"O��ʳ ��Bq��[����"Ot����$�Y�a�%K�0�"O�`B���� ��Iz'��,0U��"O �����A���3#��R�h��"O��҆�Pt9�ER;~6��"O` �Y�jԺ��ӾFP�=��"O��� �]�4�J�n®F�`��"O<�����i�SlZ�t6���b"O��S��V1�"��p�M8J9Dx�"Of�(CR��僳�OVeZs"O���O��=α���Q�
�P�"O�$!f@W[��=9���=�)Sb"OjDإY6}�`r3�N!T,�1h"O�9T�Hc��3�b�{�2T��"Ox�k���6�"pG�'7�j�K@"Op� b��:�aS ��;�6���"O>1�`HGoPtu ֍�< [�1#;D���M<r��Dj�%�(Pm��+F�,D�\�O��K"^�A���F��<↥)D��2��c(l`�U;<�J��DE:D��8�'ש���!"�)�N�5�%D��c�mH�$�Ut�&�0͊�B%D���u�֐VjU[�o�:�PP��#D�P�ʏ55J8�*�/���<@�!�"D�,jp ����Uq�H1�;D����@E3a�v\�p@R�}�ٰ�f:D��P��ѽf�|���GO,(��=[��8D����a��4���"�%]���p c6D�|�#E�K��raQ=�z��C6D�Hy`"�o4@E�uˮ�0�f5D�02�F���Н��EG�A(x��Ї=D��zg H{\�g/� FC@ F;D�Ta�b��~������/j!:B&D��Y /	;T��#GH�5"�>�r�B$D��K0�L�z8��I�']�x� �"D�	�N�w�X�%VqA,�0�"D�X��bȪqX�M���G�(�9r&,D�XX�I�(�	P�#��Ki\=)��+D�$z҈�0p)L�0��3�XՐs<D�H)v-H�H�2p��.ϙ.5VUzф/D���"�Բ
�(Ij��ٜW�j�!Q�"D�X�JO�I
@ہl͋8ܒ�
Tm?D��k�IK�n	�IďI��'n D��c�qD�Ia���4mZ\l+��"D�H��65����Q�O&Ț$�-D��CZ�Mvڅ��:qdR��2@&D���Ʈݓ pʀY�͑n�8)#�&D�,Z��8g[4���J:0��Cc�$D��1��rn��٧��<J��@�/%D��h�n��0�Į�K�Fe���!�yRʕ�� 0��;��!qs�ϛ�y
� \��-��2�9H�UH�"O>$�N;Nyb0�%1��"4"O �qg��q��Y�K�lwfxE"O.qV���H�Ԩ�j��6"O�!bbl���LY3Q�X�R�!6"O��J@у�ȱ�Ч�B�D��"Of�"�䌔�B|k7$"@n�"O���L�L�D� �47����"O�����'BP��6bU�x��Q"O�٣f�
x�'�^��%��"O&�[�cF�,���I@��Y7"O���@#�/}&=:�'D&Q{L�G"O�d��.G�U�%X�Z5Q&��"O�F�]Y���d��Hk�"O�x�t���.ࣀ�S�D\�"OB�@ ���}�Fm	ÏU,��A�"O�h�J��r�\I�p��9r��)�"O)�t�� D�EACH�rZ4�0"O ,cCD�	<T���[��p@
�"O�����:;�i�B�#R����"O�`���@�]X��1G�ٮnO�@� "Of`UMߒ-��yr� ���"OVA���-��Y��4|���"O$�M��f��#ìX�ȈBA"O~�	1�43(j��1"�(����"O��/�q*��pq�>mm*,��"O�(�I�?�H5
��^,h����"O�e*XX`r�`����Y�g�""�!��nC�q	�-ߪ7����`��3>�!��;}d���b#
��@�1ʛm�!�D�'�:���dI�R�xk��:!�$	� �[�˛� ��|�Q�G�!�d0h	D�F!�h�IE�!��9(0�8`c�֊W6��Ƙ z�!�D
�(	�����If�����!��0V PG�����@�$���!��S�K3�����b�d$�%ٟl�!�à5�gC�r�6dA�i��f�!��X�iJ.ѓĆ�f���IS-V�!�dA�M�ua�̛�A��q�'ܚ\!򄗣"����(E� ��!G�*O!�D�a ��[f�ϱI�<M�
�!�$��kM܄�Q%�`�$ر4X)0!��T"0�T8�n��)���E�%X$!�$��2���Ԇ�<��uKŋw�!��&
�ą���PQ5�P{��P�k�!�$�f�4S���R3Z�J��"r!�ʮPQ��a�i��P�e��+>!�Y�(H�xi �G�Lp��,!�d��=Px�#ށ4n�� %�;4�!�F/9	�B���J���FB�!�d��*6*��"�'^V��H.!��[4Ur�!� c^�}E2acp�M\�!��Q�X���K�n94E��m!�d͔E����
ơE3���C=E!���<�q�C��.b�s'­E%!�ď��P,�/��� �`�*|!�,i"��2E�֒|�T��!�2;e!�	��@�r�M�0��<�7g@�!��W'f�0Ҳ�S�f�*u��/[ !�d�a.�S��D�@S"@1�i�{�!�ĕ�dQ�&�T2xRb��.!�$��y��''R���"�@2�!�-%#nt1g�m���0ţ�*�!�� @͡�����nY4Ɂ4.T�6"O���X8��@��&�I�"O�|�U�ݦn�ډ�0ͰCH%�2"O��Qs#N�"���ǰu2���"O�u	���e���p�/76L��Ȇ"O,%�n�|���mD�3>��s"O
�r�:��x����eE���"O�-��W!�
@�r%_1/���"O�<q�S��tH���z�R5YA"O��A�In��	SÝ/Q�i��"Ohp�m�[�P-���j�`4�p"O� ib���}�BY�_�lds"O4Y��±>��2bB
� ʤ�c�"O����m�%s�nqx�a������"O(%���^J�d�G ���P�"O�K�H�:u�%�d.��u��p�!"O: �W؁�:�C쓄c���"O4U�&D'�4� 7�C�!�ڸ"�"O��	�#D 1F��`���!�l��0"O�]��H�|����xb�a"Or���i `!"�g`�j�&x�c"O@ ���@ E����ŮW>V�<�'"OZ�ьJ�1��`w�N�s�c4"O꘻�G�%@n椊��1��@��"OJ���݂y@FXK�9��L#"OQ�L��~�:�nRm��"Oށ�HZ�%���C�<t�K�"Obx���W7�;T�	3J�W"O�P�HN/Q���{�oآw�J��p"O a�$�t|���h�]7��"O�d����>��n�Y9�֝r"Ot�p��W6/@�݉�$�ΔB�"O������'���P��(rZYpQ"O:$p3��h�e�w�����x�"O����e^�c����#(0��s"Oܰy�@N�LE�ڂ��u$0!a�"O���r��,#	��!��
����4"OJ1�� E�r�1r◀b`�d�p"O@2b�JX�~("%�=~p5`�"OP!s�ՐeJ�UB���= �><��"O��XT��J[n]�Ѯ�d��|9T"O��t��o��`��9i��yF"O��@��0h�@�ң��Q�"OVD3R�M�f�&�ɶ �;����u"OXX�N�I�Q#�͂�n�X�"O�	�G� j3f�*�m��>��m"Ot���萏cH���6'��� �a"O��Q�D�35���+q�Ԏ#�,�&"Oܵ '��!���a#/��B���"O ��#b�n��D���!!�V  �"O�ᄡ�3�F�A�-�$8�}�f"O�	~�@�`ul��1|If"O �:D*_1}�h�K��<e(��:"O^M2�([
4�� �')(�8�"OV�YE���w{�I���P��a�"O�k``�N`� S��g�؝�T"O�q�s
   �P   �	  �  A  �  �'  `/  �5  �;  CB  �H  �N   U  b[  �a  �g  .n  rt  �z  ��   `� u�	����Zv)C�'ll\�0"Ez+⟈mڙ����8FT��D�@����n
����=QK�4F$�|��p)AG��b <9� ��f�~���=FH��'�������*��r�����&1D�``$Y�� ��VmN'>zAfg�=Ya�	H7���� �������/j�q���
u;���J�4^,>,�5͌�:����	$~P��2�",25�۴d�����?���?��j7�9iu��:�H��ýj������?�q��2!Z�Y���I
Y�j�䟜�ɽ1V�]�t挢kɾh�Ċ#l�2,�	3�0y����(�IN�6��S6@��j�8��="X"�(���6��	���4(�����<��V�9>~D�A�E�$~Ʊa'e@I}�3O��<����ē*jp�Ŗ�D�=9�aԏr��������Iן������	����O��nX2_0v\��b�@Š59�
P��jd�ҽl���?Y�4�?!�#���y�]o���LJ�c�g������V�d��aR*��x��ézF�A���5*��@��b�*��]P�X�H�h��&.lӺ�o�?�����;f�T="}$�1��0|&Z-�R��|�:y�ɔe�ɫ��u�Ƃ!z�8YHBb�֟H�?y���c���@��]�|����ѭ�?9���0?�%�A�>s���ĝ-s~�&I�b�'A��'�1���a�/M����f��W�"�A�X��G{��	�&O�R�t�2H�XRUkZ>���$5ړ�?���?��F�?���?[� <��!��<U��[��O~��?q��?y���4 �d��@(˄]��@��#��� mZ>H,p��Ř[��4�$�6�H��8��Ͽ�cV���C�T�aP��:4H@0!�+yJLB�a�#1����Q��O&��3?qgD���zD�=_�|[����t�����?E�\~v]C2�6A0�k$*���R]�?	��4�P��	�@0PyI"�՜&6�m��Y�(���3�I�%~�#|��w2b�C,a\�d�W$�a�^���'VdڳN9U���Qp��'�d�8�'2������̝xK��tZEJ�'�Q ��X>
Ѱ�b�/Y�?Ȩ��'Yƀ��%=��a1�)�:����'t��c*وm���*�3��|S�BYlpGx��i��Js��×.�W`4��l�6�.C�I�b��s���X��'��L��B�#}	u#�#`����̉� ��B�I*�����ɽ[h\h2cƐ*ޢB�	�CKV�V�K)0&�1��i��B�ɸ=q��;%���� �s��R�w �˓y ���Sm�mX���>n���P"Ń&B䉼Om���,ڣ:�j}�A+����C��M)��Cf�	\a��qVF�}ЂB��+�8B`�9�XHB��a�C䉙{[f	Av#�u��!�#kذXH���D���'�DX�w�"L���UGK1P�\�R�����OB�d�O�Q!�.߼UZM�3�Z9a����ңj	P\RC�L.	jYr�	�'0����d�� G��c�ߚv��ᢆд?MRy��% 4v�0E˟)�芧a;�5��x�ɠ�M[��i�N;t'��׭ζ/r��#��o�����D{B��L�/���6�-	<�e���,9��b �O� ���t���Z����\�`@�#�'��	by�n��=��O&��,c��zPo�l���Y͐��C�I�0xby�f��a�@�1�fP�ҒB�I-i �MQ�%���?c��H�"O��BA�u>�ئ#A�D`���B"OhL��J�r����e-zV\P�u"OV�pL�	cd���"L�?	ߒE�`dӎ�O,$���������OD��<	v�1j� [V`�W�D=z������) 8A`DY1&��M1��(������ē;t6�
�}	d�YF'L�<��Ź`�xҖ��GUu��[@��E�'E8�'�D|�w��
idh*#'ݯN:���i�ʓ8�~��E��0�I͟P+%��A0R�h�<�\mt-Yɟ4�	Qy��'$��_��00�W)�|���R�#���'Zv6͛�a'����?��'[�]Z�N�?�^Y�EC+(����`��y��'<neJ�k��&T�x�c��/7�Jui����x�����E�"��O{����I�5��H0
�'��E��dJA���I��J�&n��?�S�'�b��&� lm�1�f�8<6�H	�'랅��P�)�]��7MrH>	v�in�'vj�jv�<�	лdT����؍"�iۗ��5WmRW���	ޟ4�I�|�N�C���v�^] ��Q�w��� � �M"r��}ˁ�9[G,h��M,���,s4+ù}�ġC�����PD �	F�x�B/��d�A��0��O(9��'�����ha�G��ds���ڈ##�7�D�O����
9g�$� ��2����w��L��"D�O��
��
2lD��-��>T)ٴ�'r��cq���S�OJ�Ӌ?ຉg�0^!rAI$�pF�ɭZߔT����S�iiv@��ȣ[�jI��>�t�f�ޠ)�f<�)�']������3)�\Q���&�F5�'S��:��?�K~���4�E_bB�#�@D�1�̚����䓴?�	�k�����m�=%ldUQ�kѱ=�V�D�m4�' ��Y1B��gh�5)��Ϻ	�^��4�?�,O��A����$�OZ���<ѳ�8w0fMcV�"z"�� ���O�܀w�H�Vq�xb%$DÄ13��݌%�-�%�dv�cG�h?yR�_s���|�<YB�q��D
`�7�2�� mڟ*�4�?�Z��?ݴ���<�':9�!��ǥ(T�r�
!Bd�fůO����<Q���O�50�,]�4��q�䋡�B�Bq�'�r �>�/O�������<��=�NLRJ�L���F� Y����?���?y/O1��EbEf�6<"Y��튪T�(�åeS�ݢ���8�pt;ƈ%e.��EBHSH�IKȧ���s���-hȴ"����,�LR1_�h���	�%F�i��A�(�uۅ\2ij���O���O��,F�D���L�<�Q#Mɠl��2o[���=�yr��pp�d��I��gZ�!���O/������']剓�P� M~2���+�d5����X+P��ҟ��')r�'+���$`�0e$O�r��,&�t(J$�з~o ��!ـA������*��k��S��W#���@ �!���a�q6�5P��O�<�1����O�հ��'aR��@��E[	UG:������3b⬣��<��O����(�&�b���� M��Jq�0�O��=ͧgqb��@����>.�QHŪ���?9*OJ$��U�9&?u�O��a  �7V��L���hM�IX�'�)��LI�.��:v����WF%1��јG I�����Ө�+��Eȵ��� v@\�;v̝�ю
.-Ө��&�D��o��#��(V:�Q����qY���'�r�����?)��	�O�I1D��7g#���K�U��LK��!D��B�AP��	��K��|`4E<ړ�?���	�\d�ܛ�F�RL�L)q����4�?I)OΘ�������O��Į<��G?3�͂Sk�aJ�9�LMK��.o��e�&��: �e�C~̧��6�p�;bF�F��rA�8��%��C(?�E�0!.<�|�N>�!��<9��`@��܊�F�̟��'	�=���?����'�Π�̍%V���5%M,�~�S�"Ot�� X�Hh����a-x�C�'.r�1��|�������@IQ�v�(d��!�+6�ݡ��Φ�Işd��yҘ��FMH0���(e8���ǚ
d���R�^��� �#a`MA��3��[p��z6L��f�2q�ӛ��M�����Q�$1�Iϳ!9��ch����ON��t�Z�%N�A�Û�J�^��h�T��'1�'�r�9O�(��gF(�h�6菂.~��F6|O�b�<�C��lxp1c��Q0y@ɳFf'��O}���K����� u�84�`E�=V� ItH�>1!�dɉG���2��fS�xن��OI!��·9NL9	 a�1N5�e$N=D,!���Ԍc���{,JE�w*�X�!�$�z�i���X"Tň`��}�!�D�?7b�Q�Fɭb��MiħA�ўp� 2�'U�*I� �W�
,1爫����ȓ1��h��T�@d|��C&lTz]�ȓ=NF4���)�`�1L�,rlA��8��I�A/ ���8i��M�.O�`�ȓ(a�1�Q�LD{�(�ˊ6��=��[N9��ŋ�k`����K�J�R��I�T�B#<E���MC_&��5�G-S�u�F�(J!�d_�/��`+�L%IJ�th6�աE!�DY��n�y�Ūo$U#��$!��1W��z�G�t�~}: �ڼ:�!�đ(n�eB6�%��})�X3w�!�D\�8=� �&p����� �e��I3(g>���O$@\�#��>p�ub&��a�!�� �uY��ؼr�p��4=��i�"O�!c�GY�@�� Cv�X��i�@"OT�kw���*�7*':��"O,� %���l�ؑ��fÉ,ح���'�&PP�'�T)�@&�D�Q@R��wJI	�'�X����ǩ\���z��5qh�	�'�0�(3��-gf�`�T�)$��Q	�'�^���`���踇k�y^X���'��9D��d���
G��u����'�0d�I33��}ö�وir-r��$s�Q?�°��I��m���T+	�P��.'D���IPw\#b-�2Й)"D�PS��"	�42WG���+��>D�D�6�]*'0`"�	�mӤ9�7�;D��H�gU\��ƫQO�4�/^�!�� r�&��udO�8`nњ�g *8�����O?Z�ޮ5�J�ˆ���{��tɇ�v�<���Y��0���m��X�h�<� ��W��p8�nL5X�T�A�g�<���,H�aJT��h����|�<�6cT;Y�"�H� R^�P�����u�<a�Zr�Ha0���'���y���qy�j��p>9em�;0� ����-�L�h��Kk�<����� 
���*0Gz��/�f�<�C��*�(�iu�Qh�
�DAc�<����(06m*�c��<�zIҧ��^�<1�D}�b��3��3n�,ʵ-@Px��1B¿����D>��z�(Y���ի���yrJ� �&�V`�V7<��B�-�y2�D�?~B3��H3M#��R&�=�y� M#ga�U�#�Z�M�!NZ�y��J�g��E�T��)a��y���[���G�Qa��1�Oܙ�hOT����$Y���B�C�A� ݱc��&#2�B�ɭ]_�� ��#Uo� ��,�'�dB�	'`��a���hԦ����_�'�B�	??���f���nNȀ"Gc�Fe�C�I�lG@���h����H[0bK���C��=q���3��[�38�TS�O_-c+����U�"~�Bb���4����Ǿ(+X=W�>E�ȓL>I��	��0��)��&_;x���z�P�u&F	i��rMܳiR	�ȓ �tY�a�S1����.�#�ژ�ȓs�p�b�0br*��t�ٓ(��4�ȓ�1a�ƙ="Ќ�C�Id�65�'	v���D�,�Hal�8U	�C��x��܄�j�|��3Ɓ:+�HP�B>����ȓ-�u4-q���؅��;0���P!�:���Z��� ��A3 R���\7(�a�����	@��0W����(� y�1 Q���{�[���Q�8��>F(��cA��vqb'�'�&��h98�1*K&'XB���w�����@��@��-G9L�bS�U�'��H�ȓ+ԅ�Nғ|r��'�J�"2��Ր�J3��%d�AC�У^ΊHF{�f��ۨ���sRD��&�`�"�%�1=��ݹ�"Op�!̑v�Zг��?f�X��q"Oh�Y�֎{_M�Np}��@"O��i䎛�T�d8�2?{��Ҥ"O�MSA�>P���t-� {���"O�d*�dT�Z	QGo�k{vmAV�'�ȭ����Ӓ0Z��aQj��O����W:��<4-B�O�$l�T��m,<�04��S�? ��g+4ok4��7�~��"O0����Ӷ�(y8���r��u�W"O~��%J�NM�X�g̘8ֲ�i�"O�s�
�8r>m9�Jk$���T�4C
'�Oꭋ7B�#��<y�IܢY�0��P"O.}���lˢh��A �m��"O���O�A�.�s0�TB$�+�"OI��!ܯ��:��T����"O4�3��2z,�+U`��':���'�(���'����F�ѥ&ܪ��pE���${�'�!���e�� �e����x�'�$iq�E�F�֑��!L�0��'x8�w�fku��(Ī��I�'4�y�hN�Z>�K��Ʋ��Z�'���R��3En$@צI�p3t�����9Q?M{G���x"�aڽ]��,zH5D��i��i�NT�Q��ig��� 3D��Rς�y�Z|&�N+��4�!�ď�f�Ru��_'�P�d�D'
|!��$����b9"��+��]�4o!���#u�n�#t�L	6�J5㱊©xdR���O?)���G"٬�ʃ�?XaB�e�S�<	��hT�4�Î�4M0U�D�<��<a�H����	vt�fj�<��������i͊NZ9q���q�<i!㋦g��	b��R�0��Fm�<�Dg�"zV*Xc	(Fb�8��c�Ry��S��p>	��C�MW���7'V�e̴0��AY�<!R�O�e�Х(��T��ǇS�<�7��Iy����=JԮ���L�<ٴ�Ide�	q"ϐK�|D:��d�<QqS�h��0ɇ`�	.�L ZB�^Zx�ܡ�C��<�AK��k� ��SmB W-��8�!,D��P˛��b@�c]�-�|$0C"5D�j1'
@>|P�B�1~�Aa l3D��a&DC�"�^�xE(̾�°��;D���rEЬ.���H�y�t�P�;D�p�$�]������mǂ5`�[ѭ;���tG�d�Mexݰr�E�'�L|��ϔ��yb�\/]��1���_/m( ����y2nҳ3��5㢡�{4���`GN�y��W�^��t��J"B�\����+�yr���M;��#T M�Aq��rF!�y"Kݽ��p�U�18�=S�Ӝ�?qg��x����"��2��t˶�!�cPЭ�`�<D�,T��$��t�K�i̩�3�,D�sSGQ�:��=Y��� Ԟ-cM8D�|�Q��O� <1�C�"3T5���6D�l5��k��@���E�m�Pա�o3D����ǐ��ԃGň:=hY7f�<����z8��X  �!k����B�ky���Ǥ7D�(�P.܇~�v)1�@�Gd��S�a3D�D�B��he*�zB��B~*a��1D��Ѣ�X�6$�B`T~��v�0D���rHC�&�"7�Еg��pE�/�Om���O��Js�')$�A"͓bv*���"O�
�LM�@�h��ػ;Yʰ�B"Ob@�s��6JS�,��H�U�`q""O��
3�>O�Iш�!�l��"O$J��C)jbX��s�@�-��݋�"ONċG��d����a�t��1�l�~z���sƚ�ⶫ�$�H,af�Py�<�g�'�2� Q�� xg�x�*�|�<�>)�=���=W�	2d΋{�<� �M�!��:h�ڠ	U�ʡ=�*E��"OL�d1�x�YU̖�����R"O���`�MqT%:��K��(i���'��*���S ;ͦ\ ���?F!V4���@}�����ʵ�N�Bˎ��b�A!9f�l�ȓ�v�b�썊'�&x�5��`����ed=�� �(����"
A�I,��ʓK�TZRD�6xg.�)��0I=0B�	<4'��7G�9?
\�1�����˓bՇ��	!JY�"J�9��H ��)C�C�4Y*��� ��uo�YEA�
H�C�I�Ze��0]���Cg�,k�0C䉪�@Ia��ʯi
��X�ROC��'g�*x�cc���ϐ5aj��$O���D݌{�<�B#,��-H���3H5u!����8� qH����%�-TI���j���xe�M�#J�9H򮊯�yB
�y���`�3s�<���CU�yRI��K�ԓ2Y�G��ԘH=D�pA%�w��RM���$1�=ړc��F�b�R5��q���Y�������y�.�,�؉���X"%8��%��yҧB�:���w*�W�nֺ�y"@^�}� jP�~6���Ӣ��y�mޱOt�0@&"әv"�x�E4�y`]3���1�)b������?���^����P;A	ܤx�z��e7���$)!D�Hi�+�n�lAy���HEi:D��3H;&=�皮	��%2S�8D� ,u�N���'Qc0hrgnH�SG!��)V��EC�$	]:eÚ�J1��$9��t�SE��z���� BD��L9Ax��=f;��%W�P�2O��)O�X�g睽q$���C� ��^ *���<����?y��R�"	0�����H��b���a�+s�Q�����΁�C��IV�i�4�"s�Z��"Cb�<ru$͘,�5ӳ��Rũc��0!�jp�$-Y�@��)b�+9u*���O�b>�(Wly& P�,��{�Pi��<�+�Bӣ*ڛ �tj��ե�j�'��F{�Oh�˓Bi�K`l	Km�x3�F�S�Hԕ'}8����'��S��O���'���ʃ�%r� ��Q�
nnA�"�'���X�Ěb�Е��?\(��5NI�O� �"T�U=jz�,�A� �1���
�'��U��/2J�0�˓�w� k�-9�'b��RCc�o�bBrBu>V�͓67�!�	쟨�䧭��ɪ��U�a��vu^��H/!��T�W(⤀%C�#�|����c.�O��$V����bڝ@���ʒg߂2�s�-��Y&"Z��qEg�������d��_y�O'n���4r�K��Ƴ+\�@2bd���Zä�-`P��á����I�D�s��#�Z��i����r�9d�Ԁ��� �aV��XB-NF���&��qV�aWIX�(*��x�����$�{RT���ퟌD{2O�mò��)^�N=h��C$|��2�O(͈D��L�&���تzo���d��O
$Ez�O��]�X�c>��Q�$e�/qL|�B���C��[�4�?����?�+O1��X���T�v�i@��!moj�mo�S�\��B����9\��9ȍ�$Tf���D�2
�E`K?5�������,��@�r$AL|p2��`�'�b���h��5B"#��'��a�I{�����hO�#>)�@.��T�3&��dkgrx�0FxrD��
����С˷aߦh�F�I������	�If� X���JH�jN#߼!�� ���t"OL!����4aBP	�
~&�Y� "Of�x2�;[����D}d�a�"Ol|�"eVk l)�dתrB��5"O�I��G��Г�6s�ʥz7"O2�Ц	�� 4�rsc�.�J��D�*��O���S7$��lٲ�Y�fD��Q�'&�� �+A+����O�]�"���'���)��$��Y���&ci�܆�S�? txA�NJ�e�NL!�cM�N)��z�"O
͊Ӡ
�<~љD���|�X]��"OX��Fۥ{������"%��!hʯ�O��}�r��h�Q�͜c���z�H�2�^��2��P�� R�DjPJ���X��%��]��P��G/{�B<�E�G�[3F-�ȓ{���(af�>9���Ĭ�� ���Hj�A�	qB^��lO %J͇�%�2�Ȑ%8x�� ���w�H���O��3��'H�� �4$� ݩ��MIb�0��'9��8��ǵ.�6 `OG�:���8�'�6�y1!ӛM[�)��N�,���'3�)��\�y��	�4��K
�'��h��	��8��I�.r����'�V]!%������RH�[9�q��'�`*eN3/@Z՛RQtdy��'R~ Y%���]�b���FC����'7�E��$zt!+""[���q"OҨ�V��&M��P�n�^����p"O�<��b�&	�aʄ�"��Ś�[���	�@'��|����.w-�W��R���pt��u�<�a�N!�
����M�ي�' |���M�O<Y�F0�S�}�x��t�3�6m0�
�11��f��$ӱ1��S��'����#�77��t[ա�/*��q�O$���1��I5q�"�'u���9���< ���V��*N\��"�ڣ��I�~��s��yD��+Z�p�C��+��}H�&X,E���'S��'�di8M�<���p�Ӄ�J����q�e�\�K��'ܠ�#N�4X��3�'l�~�+4��%f��ڢ#M�^V	��A����O�O�`�>y4�i� �ꂥT�tP�892ᗔ#��I�/O�i��>ن�S!lp��ʢ.ޑ?`�kq�G|9��'��� N���<���y~�g�Y8�!Qr!����e��4����S�t�ҋ7?�a�-�'i��Q d��H\.a�Ca�3'��������
A�)�iL��|^Q�5��eR&xh͇l;~p�I_$aH���f#�ᆞOS���Q$�y"M��}8
��7��4N���1�M#���?�N>i���i�O�����R�ɢ:�1yD�5�d����?������O��S�禽Ga��_Ly���2 �(���<D��`hUp�D{1(�*B[����#<ғ�p<��ˏ	(j�Q�V͝6�8Lk�(P�<�&�A�>�����!dJ�Y0�E�<! ��6V�
�1���Vy� ��~�<Q��i��ERt��>A�EI�a�<�&���e�H(��[�/c�Ȱ"�F�<!U  =*�i���;k�h��jO�<9 �F�LT��J(��_R|A����@�<y�"�({�p�+Ƥ׆i�g�|�<�m�TuΙ���"K�|L3��z�<!��J:t5u+�I��؂ê]�<Y��\3{*�!r�A[�@�L��F�W��޸�ҢO;b�B�+�24�Bɂ�n��#1��/H��āW�(S��&�O'o��ċ��Cv) p r�M5\"�S�*C�&��d�ԅ+c��@=[�
d�R�?bW@�'�d�)��Y5Q�֡�6�F8&lZ��!�t�F����R5�d�a�ڑ/a�'��{�͛�h��m�U�$Uh�'���1�ٵ�����:��l��'�d��K��z���ie�[3?	Ľ��'f��%�F����z�㗾D�6���'�p!2T�|��Y�^�r|�ѳ�'�,�vI�B�^�`���$d�����'����U�O�-HsL׎h�t9��'�*��'đ�'/�C��
�Z4Y�'����U�� z�8���/��	��'|�,��"nt�U+�(��0~�|0�'�L`s�q�����KK�>�<H�'���XTk](O�J����M`,���'I���뎘.!�`Q�SB�4��
��� ���"�>P`�����g����d"O&!3�ZQ������)��A��"OlSU�M)9�ّ��*�v5��"O&�٥E��%�8�:�B '�Mڇ"O��j3_���kE)q��R"O�%題�1O���rsGC���k3"OH���,-~�(��@
óP�T�	$"ON��׭ޛֵ򡆝�� }R�"O�� F��� $� �^>[�&Р"Odh+�H��,l �%��ʽá"O�4cЁ��@1X��VDU�m��"O�� ��,(6�b��FLb��s"O�c#�'G��{hP�pa�"O� �%EF�wݲTK���� �T"O�i��잎3�npc��G����&"O�0����?�vL2ԛ7����"O�� ,�-�L4+��Z_�b��"OJ����Дq
�$�@ �S�z�j�"O�J��	#[[N��5�^N�i�"O��!��-�&a���׫ l�T�s"Ox���܇RV\"�n�@2f��"OΑ����; Ŋ��/_ �#"O�i@DI-D ���i!D�@ظ�"OZM�#ȟ={>P�(�@<r�� �"Ot�1爷&b�(�OT):I�9�"O�42$#@�h���5l�,2 >���"Oh�(C�ρ	ժ� gj֥Ix�t{3"O z#Ά��;�(\ #����"O��QB+��4��q6H�-�ph"O^�A�����@�E�!~�0Y$"O�xH�@"���S �N�2�"Oh���� r|	S-�i|��c�"O"���+�2�(c�KݘJvN���"O����0�t;Qʉ�,^L�"O��Ѳ��2,4�sH��HjV�s"O���ø:j�=��fg.a��"Oj���
� �`����sM�@�"O*��4�҅(�@��E��mLah�"O���S�T-}-���/�?mS��"O�4��ӾJ��8��oN��"OH�0�@56^�q 읠k' ���"O��WM�%+�ʛ. ��C"OZ��'��/}FH���ޚ	:}#�"O�)e'R@޽aq,�ߊ ��"O&�ˀ-vA ,I�9�D�V"O$�Ǌ��[���"��Z�[�0p"O���Ȑ}����Iu�`�`#"O���d�5j�bR��n�ڸ8�"OL|KC	�p�ɲ�c��@��"Ob�C�E�bY��P���0�G"O�dZ���~�(%ɒ	L�;��D�T"Oҝ���l0`ѥ����"O�ͱeg��r��eȝ),�"�b "OJ�Y��ǃ�8��Rg̨fX����"O�-���V
\@���O�A]�D"ObU�p,I?=#8�u	�;|��a"Or�9Ư�dQ`�2�A}��Dy�"Ox���0s�`��慃.�d�"O��z�G�O8�!R����N���"O��Vʒ�h��}+eG�GX�)�6"O��a�jT�`���/u+DH�e"O1���&"�$�豍WA�^U"�"O�r�J�h��a��EЎ5
�"ODiڧ�U7-sJ�R�F�8��m��"O� Y��!M}�p9R#��rA��"O�%s��Xh9Ȓk@t7�Y9�"O�h@'K�>!�~��bjR�RĤ""O�P)g�Y	l�*�
����̚5"O<@1֪��@�� R��Z=Qኔ#$"Oj9�C��vM �"�F�9*��j�"Or���c�d�X#f�"p$��z "O��0��u,��
e�"�aBV"O�����I.U����O H�X"O6�������Q��)�q���"O �2B��	U�ْe
��8(�"O�)�֤Ƶ-����� �4�F��"O�����#8���#�&2im<�K�"O
����wK�M;4`T�\�e1 "Oµ�t�+o��I�	��s=H�	�"OD��4a�4蚶![$ Z�0R"O�I�AÉ�7���3�YU�dh"O��jp��>rsh)C��p۔QyF"O��Cl�%c.uy��M>d̬��""O��:��k��2A+L']���+�"O�1���
D����Y��	`"O�U:1d���a�^A�z`r"O�QF��ic�ep� s�l	*�"O�5�4�Brr��9eF֟�P�u"OZa�q
��,4���T��H��"O޹����<K�X����!�4��"O��5I5�N�	���-.�4�R"O�L�V�D�L�\�ɅXAx��3"O`��wZ����N�:�*-�Q茯�y���1ծ�h��=YY�AH�9�y"C	�?�8;��V-ް���Q&�y2n�i Ip"�	``=��(���yB�ǣP`X�2��� ;�W3�y2�H<��!z��c��A9F+�2�yRK �􄣦�ưlc���E�§�yBc� �*�R�ɖe .�0�
�y�֔�R�`uC�3�h�
�h��y�J�N��-�TG��W�������4�yҧ=D}𝣰��!&����`^�y�ǈ:A2�� ��E�*��xk%�%�y��^�gD�Qnϒ.W��Y"+��yb(�#m̂)R�
J!5����te���y���;@���w��%-�RK4�T��y"OM�!<�0`%W��e�`�Y �y��T�g�K.I�ܘ뒏���yZ�i�wO��B����!J�&`����'w���RAԦMO�k��ث#�8�'��c(�7�����`�� bY�
�'f���n	TG�x��ԅeov��	�'\�@/³*�DAC ��bR�	�
�'���JvF�u;@e��'D.����'���u 	�7����D@�2���'(,���Ď yf��c.n4)�'��5�t��;3��Y	ׯ�gvB5��'��c��Ͼ@��1cfǑix�Y��'1�B�ՖLH8���5_��z�'��Yh�K��	�F}����[��	�'l<ԣ0��m�*|K�
C�MqH	��'h$p&'�9qv�e���W
{����'= 1w(ǭ^-��ņ�\�����'�����/F�;����M�&i��'�F�@GOʵg�F{G^,IW����'��1��dX�qzg�I�P���r�'�zq�mR�mN4�{%U:K�b�Z��� ���e����)�hP.O����"O� �Vz�< j��֮bx2h'"OF(��nˀt��<�fMѰ&nܡ�G"O���!$͐���!�,��r�H4B�"Ot�8�'ږ m��)�e�Sx�sd"O�9QG��4Kु�ȫ;��he"OR �4-��^�,����#$����"O��Ir$��k��ɵ���x��"O�I��x)jV����¦h�?�yR�¤es�}�����D��+ �y��3shNyVN� ��2��J�yr��A;p����=N�� %�� �yҨL�p�FO�� f��*D�I,�yKT-
� 㒉z	P�jc+�0�y�jٕL¼����F�k"�"#���y�l�>o��E"�h���:a��(�yr8)�������pHi�
��y,ũVb��J�t�5AaI[?�y��ݢuŮe���g�T%р��y��ő0QH��X4R�㰁��y��	���I����\-&�����y�G�ww��8����d^�c�m�3�y2�?&�:	�GI�
q
��SGϷ�y��J q� ��):D�	s#�yM��`�	^X���ᓓ�y��!*(���F R�*��DG��yB'_��X3�ɍ�Z��!��yR@ѩ���Z�)�z�����lX�y���bzv���o�_0�� .��y���	z� 	���,��� `!��y��ӣ|��15/��;�nus�i֮�y�*�M	� R�<hj%)g�
��y2%K"&�hp�ҁa"P�����y���Xؔ���SW��f�,�y2ʅ�+�l�R���QȆ�9,��yb
�\oN��sbɇB�� ����y2��'^�je�W@P?7*����@W �yɂTXB��^�L��L>�y'�,z#xj0��F;�ـv`�yRl��lE� �BL�~��)1b�2�y�A�[�@ `�T�U���wO��y"�I)��k�	٬Lr0hJ�+Ԁ�y�*L>p�l�2%`P3K���	��Յ�yBN�mr�%c��<��!� ���yR���[l����.՟i.�飀aݨ�y�]�n��xp'؝s�$�)����y2���-͞��r.^i@ڍ��.�yBK��D%fL�@�ۧfDu���B �y[�5R�� ���^`x �ӑ�y�m\�{}>�pS��-�`��y�#R�@��5v�4�1�/�y��o
����o��%���y"���-�D����f�� ���K��y�7n�Պt�]?^cb�:���?�yM5��q2��/-KNy;0Ȅ�y��'J|
�`LA#��i �Ǩ�yR� ��2v�ɗ�@�Z��'`�-���
��0qR���C>�qN>�Qm�"!�XIZ�c��1#T}�T@Eb�<išR���M �Pd��(��G�<q��Y�d��,��/CW�l��F�<9���P�����~����$��B�<A`�à+VƄʑIbU��Q��^�<i��J���2wCс!!BE�ĉZ�<��+�n�j=p�I�ȩ��+YU�<� 6��`���u��X3�ҧw�����"O�q�䑀9X%��B�p>L��"O�M�r��$$#��f�V�l$@�5"O��[�g
�E���Ha"�7��Eb�"O9��B@8��#و��C<�yR�څL�qc�e�����AQ-��y�(ӣ_���#��K�1�P+̂�ybk�Td����\�U<D��
��y� �54f ��9��,9Їս�y"*D�i�p�O*.�̰�B��y⍞�x`�4�3d����e���yR���a���$�0N�r���N3�y�#���n�I�Jk�jVhO
�y"+_�1.ve��l��D���9F��-�yb((S�D��d@�u�D�*)���y�ӕ
�(�PLG�;��t;F�y"�� P���V�պ|��b�B��ybm��__P5+B���3�DK��ט�y���%1��c���n̨�Tđ2�y�O�qcFE�����0�
��I�yKH��ؠ��̜��x�ꋈ�y�}u�*�A�h� �����yR�J�^���s�M���
DȈ�y�F�TG�ٲr��+tXZ1��	�y��ؤ7p�z��z���/�yr-�S�.�@u�K7w�,����4�y⡌�`��t����=J�����ͮ�Py�J�]1�Iu�H�'������y�<�Ae�#a��ekGOt��Sl�y�<�fI��뢩�b�l!s��J�<���Zm|-p`ˁΊ��B�J!��ڏw��{�$M�`��="A�7)!�։Pgj����/e�F!���{�!�_(qYX�'�P��<@6��!�!��a�|��q���dW8a��v�!�S&N��Hb����tL5���f.!����Pi����b����ꄍB�!�D��X$��N�J�%Q��\9_!��ѹP8�MP"i�	~���	�Oz!�d�`)�!8�!K�B�Ԓ#B��o!�ﶀB�*4���r扄?h-#"O�x�d�?����ś
S� %C"O���Ě�!� �@��A9,�9�"O,@�G�PIf��p��)R�d�x"Oň���55�|�v�B�V��Q�"O���Q&[	c��Xj�%T3-��`��"O����뗂QFH�!fX;Z�.<��"O �a-��N� I���>=�r��`"O�Á@��J���W�t��tx�"Opv�Y"�R�"�)^ͺT `"O0��f�$F�1���%E�:��F"Ot�5'�Pd ���J*:����"O�p��C�B1����`[�z��QQ"O�2�,١INAAPM%ܚ��"O4�B'���N"��_�B(�عf"OB͛4̚�#8`�`�L�T +|�<����M�y2�
�H��0����M�<I�ɜ�}�4���G8,M��C4�H�<�d	&dic��K�ap�QBW�Yi�<�toV3S6	��BlfjDC�n�<Y1IZ#Q�d0CE٪s"�Ѓ]l�<� ƀ.2#H�*�̒��l���%�g�<�v&N�.Ǿ�&@��.B,��`Y�<9V�r��Xr�5[����L�{�<� �(����<c���ţ�OR|ɐ�"O�b5�ѫy/p�	�P.a��;�"O�Y���H��1c@���=P��pG"O���6�̵hU`�Q��$#�,Z7"O�-(Q�B�IPN�!e��`9�3"O�<��M(oW"Qj�A/8k��#�"O2�3���3=ʜ'`�w�ƌ��"O@-�Ù5`w<����?=D�P�"O��yp�61t���3@��S�"OVQ��K��nS��
s$��-פ�s"O�p����$E�2��=l��kE"O����h܈a���x�0A�&�1"Oa3�	�d��[�Ā9��0�!"O0�ppE��.��D�R�B/	�~��"Oh�I(�)�V����Ç)���'�8���HX�V�B÷��*Ta,�
�'�0��P�Ʊ!7D���SgR��'��	�AU�B��{æNJi�}
�'nd`��1bc�Ah�%EJA��'����w��2��u��E�4UN�U��')���G/ٞ1L@��$	�S��,z�'�"2.Ԣ-c2t����� #�'�Z����Q3�h����M�F���'Hq��ɕ��h�I��� ��'������<Zp�`#뗙ɀqB�'�,1a�/Y�Ș��΁�?K\���'0R��W��0��5]P��'@���.�;b�6tH�lʰ )J,��'���W�51.�!YÃտ S�i��'%Zy�"�O^���)t-0n�V{�'l�9�#hl:
Sr�|��'���"��ɐ]��@�.LX8�'�>�XS��	c�=�#�Y=þ�
�'��+"IU�C���c�F�|���'��3�.�7Y
U��Ɨ>�4(�'��BIĊ5��L㬓7�P��'�H��QEH=s%H5�6�Z�'r��p�$H2�r5aR%f�6�q�'U����U�A-F���ڎ����'�B�ɀA��3*���R�h8�i�'��d��R���B�gI� ^��@�'}
-��M��rj�=��G
1�8��'N�Y���{������`�Z�'�p��(B�XC��ЁF*7T�i�'��ke�ê[6vp�f�Y/=���'����'K�� %��6���'�^L�p����Z$���;�����'������L���`�C̖����'��5�Hӭp��u2�Q� �B���'�J�I��q>�8��H�"H��}��'r�Ia���g��䙑ĨW�J�'`0!`+��@���*_%TC���
�'S@h'��MVd���M؄D�
�']�\j��_#���k���K�vt��'�]#!��I>��h��a��<���������&L��C�9�7.�S�<ɐ��tp"𹵣V�D<*��&�W�<��V.K��#C�-m�4��g�Q�<i��
��m�ԨC�}��-h�Fk�<���� `�Е�sAV#q��H4i�e�<��dL:2��`����� ��P�]Z�<�!�M-Od���`�� Iv����W�<i`T��&�W�J�"���.l�<!��ٿY*�x���6�X9 b\d�<� *l����f|�����'l��x�"OЈ�#%|2�P���Am�`YG"O�\�T��w����t��8\����"O� ��9X*aE�Z�w�X�9�"O�X9G#�7Q�\;`��(j��) "OthPa�]�#m�y� �9%~,�6"Oj�H�A:U��:wĊ-�ذ"O��+�Ƿ"u2�a�ɔ E��l)�"O��fk�! x�XӪ��$�|���"O��[��J�r,z�P#jS!8�F�S�"O��C�O��!o�9 �&=h��"�"O��ȃ	�,��n��Dy2�p�"O��������Rx!GmRmeb)�"O���B�(��(��-؆)D����"OM���^�9��YvԖqS`"OZd�&��M��]�4f�8�m1�"O�ly�_�cm� a����2&���a"O�]s��υ}Z�d��Щ*MP�"O޸j���9�Ա�S�!(�"O���m�#����)ĕnf� ��"Oh��7���� ����w�$8@"O8��I��	�b�{���v� �"O�e�$ˊY^����m޸-�UIR"O@�Z��Pc��&�^v�@�ˠ"O��s�
�� �{U��9��"Oج��h�U�ݺ��Z+���1�"O�a���X�X��qn�4�SS"ON�6��7��Q��[��|a�"O
��)+�4����(@�K""O�y� �w�D0ţ Y�K"O�L�IP�2��b�0}P��"O�8��֦}���3B�2g���"O�)��D�'���s��(9Ap R"O��H���jp�hP���	���	�"O^���1; 	SE�.�Nm@g"O,�a��w�h��N�*k�Hr"O䱹��1O����� �NР�"O�\B#�U��������@��"O��d�;�-�!`�=&���"O��qT;Z���m�t�b��"OR̻5�P2W��u�c�.EV�!�"O���+T�@��I"Z	��{E"O:L	w ��#&�18�c½ov5�R"O:8(���*M�P�R�c��+y�=� "O�����k�H̛� �^`�AI�"O�ѕGT�8Uܽb��VW:��"O���Ĥbo�`�Z	����l�<�47.�R@0���?#l����f�<I�_��-�a%ۛ5ۢ��Ql�<)Q��`��1� ���S~�飯�f�<��� 90w�h!-�5[��SAi�<��Ԛ
;��/I�<)��C�M�<)2,߀zeh�bM3�𽂡(�L�<9��^�xz@!,4��p���G����J�Xti"'�,m����ٿ��݆ȓ/�\�(Ƃ"��Yh$�38L|�ȓsC�0�gͩ,��Q��	F��Ąȓ�J��lK�0�``���0%%h���*p:�B�ge�Ȧ���c��	��"O����k��z�ʏ8#��P��"ON��ׇ�]�j���HT�
HB���HE���p��Dl�[Tǌ�f��'?
���G�e�R�R%X�i�dP��'>�pc��dZ.%;UÔ�.��!�'kz,[���mJ.�ZU��(r+�4���� ±@�>C��8��_!8�H!s"O�8ғ .s�HM�+�#�v��S"O�T;��;Q�L;0$V#I���b"O�l�A=1�&t�6 �+:�r�g"O�!gB!���z!��?z6�}��"O���f`�N�JE@��*V
��B�"OJ��W�G�4�r a!��5EeL���"O�=������ؐ��H�(�A��"O^�QrO4*e�|H��>iZ �s"O^�2��[�T$�t�&��y� :t"O�p[D�9������@[��cg"O�5�s��`�pHc@�5i�h�"OB�[�S�:�+eT��,���"O����j��4^(PB$e�-g���P�"O��8�E($l �j<�^�l"O<�ԣ՗kaΥ	so;B��� $"O�	�2n?>D%�
_p�<kU"O.�bfNϪ	/�!H$"i��Is"O�@��@Igt��A׿#�\}Q"O��1b�R"�H��U%X�� �"OFq���5!er�As��6"�0I`f"Oh���i��R� >[���C"O�!h<
Ȋ�'��=M���["O<��"f��!e��䆃&�J�
�"O��4�AG��QEd�Z�x��"Or��un%N@JU��l،ܲ4"O�S�P�8�R=2ɂ�M"�0��"O4UX��(}���Xuf��er�q"O������F�k��R��wjBn�<Yq��;	ip�؈�v�X6*�A�<�"�9!�a�e�W<vFT�+S�q�<�@b"6k��0큷��|t͕m�<����- �8d��'b���,V~�<9��O�,Ⱙ:�v0�cX|�<��`ԢJX�h����0v����$Ad�<ѣ�ău~���ER@���q̟T�<�Х҂/�P �S��
zJ��.FN�<�7ǂ�_��!K����0�A7ʙP�<�4�5@��31�"0����OSL�<Iը����i����	WD�tu�ED�<�4L�
.�A�5�0x	������<��L�&H�2�V�Gt��	�<�U�L�h4����?x`�HWg�b�<�'������A �V�~,z!&U�<q]i��F't8�=����]D!�d�=꼱��͕{��z�1!�$�4{�ja�4aX����2C*!�D�3>����',����ʉA%!�$�&�Ш��+���J��-H!�$�`.V�cWˀ)x&�Q�	�A�!�ٷb���u*́l>���!�,?&!�dV>@�Ba��,aK��)�!X�|3!�܉��=P0ǉ�,!� a��y!�D��z���ŉ0
	"� B:�!�d�`��h�3�r;t䔂�!�A

�-�s?L�Щ!1䔜g�!�D�3et�E�? IR���"it!���>	���*](�y�m�`x!�њ#��@g
9M\~��/
pY!��M�\%�PJ�J�*L>�ң�A!�dܷjY��y���iEB��rGK�],!��<j�\8�D�!wZda�EU�}t!��
���E	d���@կ�!��-�fe{�LB�(��*�L.p�!�� ��+dj��pq��)f�	�j���3"O�5��N��<�񉍰�|(X�"O���c��UjXu:�)��O��<�"O�4��T��s�Pt��Q"Odu0"��T-8�Z%��f��ٖ"O6쀲�
�?��tK��:a��zt"O�y��gc�8��G	���7"O�0��(]�$+��A��� yp ��"O��z2��b9,ɓT��U]ޙPW"O~�RJ�Y�̜[�#�?e��E�"O���$����ּ��B+�����"O&T�� 
�X�aS&�޼59q"Obq{,Ϗf�� ���z��b�"O��Ђ���l��r@J�&�lpH�"O�gB�s�P�b #� j����"O�I
g�I
ega��?Rr�Z�"OM��Է�Pa�� .!�&"OF�� $�9p�m2��>�@�9P"O�\�(���X3A�`,"XI�"O*)b�I�U��y᧤ԯ!����"O�}�&K2(~��3�#�L)�كt"O��jq��Q2\�q��MCu9�"ON�{��˿t���s��Va2$��"O��Ѯ�;K�$`�ٮT���c�"O�h�S���X$ �A9�=a�"O@Ɂ'爕���bA�I4&%�qC"O�( ��:D,0��k�T�5"O��8��3=}�y�E�Q�K�\�x�"OdyQ��­(�,�
#j�$�A�U"Od�3HҘh�r�Z�_)~�4ӡ"O|񢶍��֠��@�Gic�]��"O�%��?r7��j6��;C_$<
�"O��[T�G΢��0
ۑc*��q�"O��r`�M?��Da���S��k�"O�%����#>�hB��.��d�"O�9��!לXz,i��]�p�x��D"O�����_Qr��$(K�%���sS"O>��n
%�
�se�����P�"O"L��>r�|� �$�j��x�"OPPH�@�	y�4�VE��\��pB�"Or�HE#\+��hȢ��j��4Qp"O&-����UPuC�%g`)��"O��aA�Cp��xaÆu�иX�"O�H$��?{.ؐۑ�A�0���e"O<�Fk�m�d<�HA)���[�"OXDYwč9nKP�*�Ǜ���bR D��x�R�-,4U@���9�1J�c1D�X� G��7� �3��e�D�JT�*D�`���ϴEs��"F�.X�d��GG'D��h0	�1Q��8�Gġ<�����?D�$����5u��܈�HC�=!��y��>D� �� ��K��uqPe��\9�-Br�=D�8����r���ڒ��J�ưz�C(D���d&�]5���󨒍Y8��rf�1D����Ć�m*��!Ԅ���O4�=E��I��
��y��C�6
��Br�ެ�y�aG�%v�=Ðm<{�P����yB��hRVe3c�Ǟ>���%#S��y���ۃe�~u�F��yB��v�f�a�OٽsaBh�Nϖ�y"	(؍X@S!"��U�0��u]!�D)Iu�ʅI�"5��+�Ȃ_K!�
��9����QЫQ+O�m,!��[�z+����Ee�$��� �{!��  }�v
�9,��=K��W�rي�"O�q�r���3�RK
�2i�#"O4��vG��P�J�+��Zu���e"O�9&��f&f��Ҫ,�&m �"O�Y3��b���7�ӛH��u�C"Ov0��eċ[@�Ģ�d�8a	g"O�0�Ì��4>�c'�0��(8t"O�ꦋ�/O.^�G&�>X�5�"O��RGE�X���d��<��`"O��������B�/|3:�p"OnP҂e�$��qD[�����"Ox�'U�N-����c\�YS�M�"O����M����@!S&�$��"O" �����4�>*�_�t�e��"O&��k̻,��w*ܞ= �%��"O��9�78�z�`U����QC"O�	ӱ��wP���QiJ
s��"O0&�8������8�2��ȇM�!�D�>���S�'� ib���M=zN!��ѓ"!��A��l�0w�
�}!�Q�ldδѷa�+X�� '�	!�$G<guμ!!�\�R�Jq�OC�!��0]�@z�K.�T��7BF�!��Y�\y �8�DĿC�2�87��'!�dM}����J a���2��&l!򄆆*` ��wǅ4T��gF�=�!�8J� x�c���Hnj�1�kϚ�!�ĕ�v�x+0k\�0���ۋ�!��b���a�MC�W�R��BH�!�ȳ!!"���!�����̶
�!�Dҡ(x��åFE-*|���M6]�!�	�[��iˠk�$y�H��֓1�!�ď���СW@�$~���ҥ�e!�D�d�����
��C`OT3w�!�$֔`� �P <�$��r��+�!�˖+QDݲ�oL%e�4�N[�d�!�Ҧ ˢ���h��nu����]!�䊴����[!_ZL�Q�մp�!��75F1:$^=HC�� ���, �!�d
�v�$�D10��H�^62�!�D�A�h�Ys �L<P+0+�,�!�d*I�3��W$?���)���!�+7}�l��J%nڼ<Y4HU�9E!�$Q�::�a�.��Uό��B�I�J8)��Y�7�(5w�G'm5nB�ɋ-�!B����"��e(�#oBB�ɝl52gL��6�PQ��0l>�B�I	u�ݦ !��%��(F��B�d��YX�kJ4ߔt��M��
C䉻t٦��3�3=�` ӯŏs�$C�	��śD'͂(������?lf$C�ɂb�x��ܿ5���D�#TB��|��4��(W�2�X	�Fr�>B�I�7V� ��C.Q@
Y�BS�e� B�7P�aJE/�4=�� �EMy��C��=@IBI����V���cg�+7��B�I�f��� �H�$\̰r�ml�C�(X�ĹBV @$m��u)�(B�rC䉆6�$�Pg�e��=�A�ʦnȀC䉢d�H���"�iӢ0�	WVC�I	<��l��@��~P����bJ.C�&u��8�kA�Lؠ�	�	�B�Ʌ1�¤�#�$L�E���BȢB��3�v����
�<��)T6U�C�)� � �N7\$�Ѕ����	j�"OH�iР�0L��3K��r�"O�uY��ט|Vu�U,��2�zY�V"O�MqW��($����6N��(M�"Oj�3b�� &�(1�w������G"O�h*��`$!Elح�xI"O�QzuG�)yH:��b�&�&<�"O^ա�K-V�6�I���=���"O�L�f7M����q�۷R ����"O���7N�B���\72腠A"O0�b�
��\k�Gp%60�"O�Usf�0V:ԸcF�4G���B"Ov0(cM�k��Tq�*2] �!2g"O����Tq�ptJ���]+'"O��8V%�[熴�B�>6�9'!�V}��U�d@+}.r���;!�F"y,���k�7J�q�F%I�^Q!�d�`���0�L��$�#�ǌsT!�Ɯ~��i*��L�K����a�R�jT!���9.J%��FR�;0�P�L!��Z�KS��}D\D���D>�!��B�F@xfm�JPd�+��A�l�!�$^�j����� 'HHyئo�M�!��C�"�r�����uG��x���+~!�	<#�������y:=`����}B!򤍂g�N�`p0���"a�!�!L�n�t*�|�mA̅t�!��A��
X�' 6i�ĝ���*�!�!?��� �~���񭟍?�!�d8����BHG3��!PF�*Uo!��\�I�h��/<^����^mg!��<S��r��)�~1���n\!�d�W����R��<D�A8� ��1�!�Dք\��{Ԉ߁g0Dɫ�@�*E�!�DF��Q�QJM�aH��8g��1	�!�$� Iٲ��-�	kF"��նfP!�$�'+f�%��n:M�v<[!n�k-!��f�Ed��:Ͱi��M�M!�Ď9y���W�̦B�b𢍂a�!��o�EPk ���#A
u6!�$�RFi;N)�L��	?O�!�DӠ8���D��%!x���� 	&�!�$ӟ��N��8�d!��9UN��"O����$K�`�j�/��t�� k�"OXD@b�V(C��b�֣A��p"O`��aT�j�B9��۶|{Vd��"O�P9O9Gr�qd��~��A"O��{�"�-V8�M`Հƃ1x��!2"O�؂�l8|�5� S�y�]��"O��� �ϖ���b�����z5� "O�(h!��nx���	m�4��U"O��ğ0F�"ڑg���x��"O�}ڄ����ixE(0}��p��"O�rQ�
?Z*�arg�%y�����"O`�CׯK�=�2i�Q��:�"O���ə?q"�v$�6?�&���"O�<�7*�shƴ:�a��}e�Q�"OH0cs/��Ws6��!��7_���"O���b��c+��ha Cr-DM0"O|@E�C8A�&��/��:�7"O�m(T�	�� eIP�ҍ~8��"O�(���O� l���{B��e"O@l"��+sL����$T�?�R� "On\�( <h�x��RBʰk�-
#"O� �)B@Q����Ba�9d�4�ru"O��� �V\���Y�oX�i�T\�0"O&��ԁ�
��HS��:!�)і"O��	�hh!����"P�d"O ���n`�`.��%�v"Ov���9d4�XB�FO;u�e"OBP���:>�43u���ِ�1�"O:���j�~�@�k�B���8�"O:1 !c�=�v9�FaG7A��5��"O����$�.ج�k�eY ?�ĉ�"O*�S�o�T.P9�$&�����"O\i��;0��x��o�E�4"OR0�ֈG?#y��'!��S�0P*p"Od�yE�ܾ{�8�A�@֑��zT"O�`1GW�b�"����?$�x��"O��be �5*�YXs�=Y75��"O<������-RWS-�R�"O���Pח���CD��%�_�yb�ջf�~���*J�Z ���yr-��A���T��?��1���y-�V`L=���@$B�V���a�y��B}�$�"Q*��qٚ��L՜�yb�$sv��A�'�1�����B�*�y�Ā*M<�����)���ɠ%ӗ�y"�È',�q`�¦1�,@��N��y��X�+�Z [�E�T�\���+�y��-}6<�1��Pn�� �M۾�y�9#ɜ��1��"̤�����ybNS 5`$8Hإr��`ō��yB��PL%OZ��`ѫCK��y2�ň&��⎄)&����]&�y��Ψ|����'�?N�Ïƣ�y2�����Mj���d\�S�O��yr �<A��ۼ3�@����y��� ��`Z�M��l�u/O�y�N��>�T��q@N�k @�hKL�y܎�h��Di?T���ybk�>B����qmН*n<E�v���y/R23��ep1/�+1V�J�Lě�yrE��1�=�rJE.���NT��y�"�&�x��%���	�.��yrIљ��Q�G�!��f��<�y�[R8@W�E�5YvO��yR���I`d�Y���,���+/�yB;{8ĉ����Y��Z$M��ybg�8�V�
�j b�ĩ�K#�y�g@���j�]B�&؉�y2���2a&e2Pg\�e�D ��@�;�y"�Z55�$(Q-�(	�(� i �y�3pvٓ@��x��� / ��yb�ɺS�,�8����nu�P����%�yR�A�P۲})Ђ4h�l1�q�_��y��BM�2	psb�!`L8��%�W��y�@�8ʚ�BW�ړ"j��xϕ�y��="��Y��
��.	������yR�E/o[J!C�hɽH�*��S���ybn� u��p���W8AL�	�U�$�yBd��O��C0��:|�m$&ޏ�yB�?�0dRi-�\�� n�yb!� {�0���KpW� ��,��yR�M0j,V�	�`�	0Ș��6l���y�c͛V*���&���P$!k����yBć�>-��o�M5�<bvNR��yb�^�K-�l�l�����0�y
� F\#R��(6���b*C�~k `CV"O:��r�H�c��2��͊b_��"O��+��
*X�,0`N����g"OT���� /�yCq��/� ���"O�0X��ܢ7��!��O[�7�j�!��O�2�p�RP)³0��I���ӧ�!�A5Q�)`d��JeZ�(�<u�!��W�N�D�	6��XH�;f�_l�!�Vx�0��_�oG�3�(G �!�dܿ��5�R��+C/?�!�I�Mp4 5�W1n�X]i��ܫ(!�$��I�4X�B�y��}ٓ,�_$!�Dˊ�Y��m
[n�xB���!$!��E�?x5J�-�"y; �X"���E5!�� ~���3�z8֍� ���!��4�m�T��,{���솂F�!��((��a���PL8���?g�!���<1
�:ʏ�s�8�(�ᓵ�!�>}�z�v�y���X�j�%!�dڇa ��v	��g�D��
gc!��v05�� ��6U:�����F!��\���c��g�) ��E!��\蒝�� ̃n̮}�f'�oE!�D�?��<	�胾:����d��6�!�D�'HH P�ӄv���r�F6�!�$^)K�x|��L�%>s��x�H��J�!��Hݴ��c�2mb^���:N !�$��&#���"�Q�#z�툴דl!�dσ0 T�CcXY����`F��(N!�$.��Q�t'K��X@�G65!򄏄l��ȁf�Jb�t3�BU-p�!�DX�]��}*��a��h�G��� !���0IFR��r�}� ��S�ă=�!�D�L�����$�8M�(1Ȅ��7_G!�ά�(#�V�y���tfзZ)!�䜕_i@	b�ʃ�#�r�Sd`��e�!�$�A@4��`ß�dT���Po�m!�$��	p`���Y�n������c�!��	twP`�D�ڈ�A�Wc�!���^?��S$C4Er����x�!�Ē�h	��	>S[�S�X��!�dC���z*@?J���teBh�!�4v�41H2eU�&����d���G�!�'��Ĩ�C�6��2Q�!򤐌c�E���\*/�v����D+!��	�>�����_��^x���׌(!�XN݊� ��"�&4�t*?�!�ܶ=EN���j^��j0I]��!�$�&[��$�s�V�9!�P����?"!��T!e0zS⌐���f� )!�ۄR���Q��K>#x)Z���D!��7b�,���BK�f$)��	�{!���g�}S�"�&� C
��f\!�$�74�(��˖i�	X�H�Yx!�Ğ�0��/ހB�Zu����,�!�M"�t��⅟	��xK'�M< �!�F�G�rE�󪗭w.�|��nŨ �!�Ě�p�Đ���3�\�;H�p�!�d�3v�I�@��!	�`|G͞Ts!��:}D��)ЬN���x3�@1�!��
���E�ȋripPh7�Φ=!�As�Ա�p-��L>��`UE�
�!�D��VB�"a�Y6��9���#��B�I�Q�-y B,Qd]�/��B�)� Έ�s�	-fC�=�₶q���4"O^��K�� ̻@��Eي�;�"O�|h������p��
;�*! �"OH,�a��8�����N�^f"O����%#��	��&\�,�
z5����\��ŨIN�f���!^�R����PLt�c*>=��k�%U�� �I��!�G"2�u��陬P ��[�Z�	S�)]F�逗b#��M�VB�_J����a�+&��TJQf��Z�d�*�&4�P�3B������m.@�%�![�}��E��?�7�i&6-�O�'&���ɒɌ�'�b1C�oā_�p�br�'��|y���'S>��D�"�XѲ��}�,ܫ
��M�D�i��S�q^ ٧��U-�A���M�~"T, �6��O���|�$�K�?���M�W�HN���Q���j�������|d�d�X�	z���d�bO��1 ��i����S�h��C��%$�"�I�ǐ�2��7-�1 H��g"Z<����iK�������H�x\�K|��=L�e�WAA,(	�B�r�� o�0�2�$�ܦA[-O�Oi�s�.#�m�+9�$l` �ZFR�yy��	UX�0�Eh�)q-����N� �a�3ғ�M�r�i��h�]�!"LY怀<?�Px���ܜ8��4-ObAb��s��D�OV�$�O;��)^�\�"��K�	<�X\��/Z�!>09�f��;��(�s��2a!%�?��P቟T�2�2�.�/Y��a��U�.Hd��m�w���rA�\�PQ�c��~��Ō<-0�F���Ð�Z;z� oA�	V�iӣ�>��#���d�ɺ���?9����D�)Pn�"6O+Jy%��t�Q�����Ղ/�B����!;����g��\�ڴ؛V�|"�O<�D[���ހ+���`�b�f�4*���}�%`@̟(��ҟ��ɿ�uR>����1�rE2��L !B����ɘP�⭚-Y�N�,��c.�:�B40櫐0~���@;UQ�DW���R.x!*��p��!b��c6g҄F�a�$��?�ʘSeǆ�Us��	�}2O��?����8��X wfC�t@����]�=A���@�i�R�L�IN�S�T!N�Ϣ� C�^�J�zة�݄�(OУ=�O�B�D� ?�� �IT��	��'�H7���-�'��uB��>yJ|:ǭԛ&�V��$k�qb�Y�喾s��dj��'�"�'O�er�G;�V<�vLE���q�|�d��*w�|5�S���KQ0�BI�{�'90��cQ�N�ru�T���q�T ��7;���#d��fP�	�\�BC6��� :#c�9��O�����	f�$�,�B�2�*� �:M���ز+�MnZO�L��>�DZ�j*�mЏ��3���8�iV�k7�|v�r)o�̦�RA,�gf��Ԁ�u����������RB	�;x��	`y�O��5��'���i�E��Ն�Zu.%�9�G(C>x��M�h�'`��4��H��6*�?��O����ʤh�d�?M��s����r(pR�i^F���Ǚ^/,�u�7<�E "�ĄT	��"���a�

�:���K2F޶
�L5BмimPA���UK��J`��d,���u^�6��dx�,I:7X�U�϶�|�Igy�'�f@���0�$0/ЪU��+��g�v\m�A�	�?ɬ�L���p@k�{�*�0��͜C#���4�|��'L��� ��5�=�v�N�<�ଋ�rUh��5ت0���@h�N�<�#O��h�m�25΄�!Je�<�c�+;D�e�Y�X����&�_�<�@C74 �h��h^�\l�aL�u�<�6 �!Y���P��T��8��J�<�B E�1��[7��).,��fE�<��n��d��S"�(�x�h3�Rg�<9X����נލe"BE���ùS��C��H~�YрQ�
\��
b-߿l<�B�I�8'��e�O((�l��#4�ZB䉤hR�]J�`Vv.b̸1��]0FB�	;`�vo�0_�N��� ����C�I�|Uඇ�]6�4����<�C�WA��e O,��a_?"rB��_vFěE��#�Kr�E��C�I"F[�XS���0t�� ��%|��C�	�g<�v��+}jj`�ܕo�C�	$|���q��2(��V)	<HB��w�@��+��A����&���:B䉏�j��֡Y�\��m���T&u�B�	�G
	J"�L܀�K0��I<\B�I�=Pny��`U<h�`��!MJ B�I-n"�����]�!HP�)�kĦAv4B�	�D3���ҫ�-:.x��?9>VB�!��h�&[3R�2�J�,�12B�	)�N4�Ej�?����NB�	(�*���l���M*DC0C�	v��L�	��{n -���9@fB�	9P�m�&�ʞK�.42"�W�ya[�-���{���$G8u!"l^��y�)DK�j<�h��,��|i�ǌ&�y�e {8�p�ɛ�!�<��O �y2�J.xyZ���r���-�y��&B��58�/�~���)Ϫ�y
� �C�ȏ�Q�li �$��(LD�Zb"O�9�!F9' X7E9&���"OD��Š:�,(�ᬃ*-9��a�"O:`�!<2�� ���D�("4� $"O�X�'��.|+��/�@L��Gz�'��`y�Tm�X�'c{n����ߥ ���$M�E�ڽ06&Ԡ|�R�'(�镖R��[�Oӭ	�V�@�� ���'%�F\���_6Vt:� 
B$��Fz��ފTGn\��I�oX��
�I��)�e�B�(�9C��^�n~�)g�ØB,p��dNnb�'m4�x6M��"�������*�d�b�$+d���[��"~�I~Y
}{$@��D�0G��8&����¦YQߴ�M�ɛ�O}��� "�� ������Y?��ٛ��'��i>�8�&H�,�I���A��W�(���#Ù`�J�s��HiB�0R޴@p��A�H*D���Wܧ��^c�!���h�6��E"u��3�4m�f�"�K�Y��1 7��Ǧ�[w�_�ZA�U���\c�ld+w#�f�R�Ƶ �P��4m�n��	ӟ|�.O�D�sӶ��@�^�q�p8i"cI�j�B"�O���+���'?�Ѡ�ǒ
�}��
68ز���D��m�ٴ��O��N�_�^Y�5mRg��ݨ�+]:jf���'�*x �bёt���'6"�'0:֝z��oC�t�F��D����L8����<B�o��&p(8�-�#��`��O�DԪ����-J$���̞`D�U դ�7]��1�ɩJw&�X&�Rd(��20S?�o�W"�%���	K�Ci�i��f��? ���C��?�ƞ�?���Ei<�gyR�'���0���Ɖug�-�f�^���h��I.,�v�S�䅖k�Q�c!��M���:E�i�6�:�4�����<�퀬/�v�Q���� � �E]�����?���?Q�"���A,�J�d�K��K2�\
X!�r�W�,�p����P&ky��6�ݳ!���(ڗ��O��� ��)�\q�� � 2���`F^�꬀s�.R�>`~�#�I׎;:mx�i�'����D�OD�*ǪW�6�l� �+�<{���3*_�>Yl��t�'���T>=��D11
��E ]�>��-�G�#}��)�S�>���RT�Z�$��-�A<
�
���M���i_�ɗ9����4�?	I|ʃ��#U�*��g�R�S����e&K�< ��Q�'�b�'w"��жi�~�S�j�?$�$�:t샍��ti�O
��u�Eh2qR�a���HO*D��N��`�e;愊���)k��G�K�����I `~��@1kV�~z�8���#kL��qd��O����l�Ҧ��sl�3(fHP�H�#�ER� ���?qJ>	�S��?9-�>t�d���RLƲ4�'�UU8� 3ݴ�?��4M�(��L�P���x5�ʱIn ��#�z%V�앧�䋟�W"��'q���\zf�m�`���N1v����Y��<3'0�aN�	[q�Pؒ�
͸O.�d���b)	�r6$�����I��i��L a��b,�T$3O�In��,�s���	Y1u�
�R@&S�)�v�XѤ�>%+&�'��-�P��0��	�����O`�{C@��vYq�？ �	ܟ��ICy��'s��$���0=��H�B��P�`���I"�M;��i��'at�'GQ&�XmX7�`�Xš_�1A�qT�|��'����� ���   �  B  �  �  �)  5  \@  �K  PW  pb  �m  �x    �  �  K�  ��  ܣ  �  a�  ��  �  ��  �  ��  ��  >�  ��  ��  .�  q�  D�   U
 � g �# �+ �5 �< 1C sI �O >P  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4��'d��-1fA�r#
<���`@�4��T�ȓ=�b���
�8s���>h�D|���P|�Ң��)O'�Y� HY"3�8B�I�q���j i�3D���"�W�! B��2��=�KV,!X�IR�d�Wp\C�)� vd;c�OG��A��Y48�(��"O�H�c_�ev�|��jͳU�z��s"O��c��.N#8�g�ÌO���HA"O��B%��,V��Q���ب��`
�"O����;���o�et�I�C"O���s&�;����V_�E9��'Rc��a�C6e�h1�&�FQ*���d6D���P<�ب���p�$�s�	9��M����H�W`���m+(�$�۴k8�O>�	in@��B��4&	�e��Lq�0H��O��Ip�V�US�`U��d���I�<y%�5�S�{j(��R��16�����@��C�I�G�|��+�Ui��Q'!J�
R�C�ɫXe	Q%�
�Øq�!��X��C�	3H��H�& G�C�& �k�HXC�	'd"�q�H� �c1k�#}rC�I@Q(`�?n�!9�
�^�fC��/V!�Y9f�7Td�(z��˦SN���D�>�a��$��d�!��X���x�ŐA�<�֊��Pی�z􂒿Ha�����z�'�?��&���"��A�a�P���5D���&�P�4���P CP�j5a��>D�\��%Ϗz�\逬�=7W�0@�*=D�p@����`z��]�\d��SV�/D���qfܪ6�Q9�ܩ���/,D� �E��k;��lT �L��6D���hA�| ��%`Πn�n��g(D�(C�� O�N�x�$��w�`��%D����oS2sn��b��vH�)�uI$D�HZ��O�ct��8~s2�`�#D�HP���;>�5� �f(���b D�$���� ٔ�9�lB,fr��<�!�䘛B����qꚩU�F1R�N�<>�!��E�f[�QiVI�j`A1�>v�!��NH"$$�ǩB>��J���!��.f�=2v��;>$�s���,�!�H{����$;X-���P�!����������~��JZM�!�\� ���XU�q�X�:T!�Ą;6����V�$��tJ�dӑX�!��Y.5��pbԭ��P�D����W�z!��U�h���0�TU�0ԃ�#���!򄌵�Z��aÝ/u="�2&�G:n�!�B.Cż����F+8>YPeφ$�!򄘖lU������& ���H�Q�!�D΍h,r��7Mi���o~!�d��Dp�<S���K�h9�DJO�Pm!��(*����p��L��T�PFK�N~!���:ct$+Ǥ�&d���f��Ev!�G�k�f-�Ć&1�<��wd�2~X!򤄵a�HK �۳tH� �`�i�!�F�N�\�F	�qKz�s �΃l�!��G.�M����f9d�@��>�!�ў_ �i�+�[ּ%*��̩1�!�$�+C3�(2�G��	`�H���!�d�X����[	�гu�_1?!�ܱO_
i	�k�Z#(p��
f !�$�32�tj�رWD��jS#!�� �"a�k�d��r��O�!��Fi�`�`f��7$9�5�0_k!�E }�z�͜��)��Į$�!�d�p���*N�\�&l�V��~9!�dOm�$��#Ɔ
�p�֏Ӻ�!��j���1�Y:zF
���#r!�� $�EbW�Sgl�V��k�"OR	�e��	dȐ�fD����E"OH��&�[:<�n��w� r~zxɁ"OZJal:I܄���� ~����"Oz��FaJ�W8��teo�%��'|"�'���'���'Y��'er�'r�<1`��$/jl��¿.�0��'�"�'���'���'9b�'��'��-q7�V9EHH��"��@�s�'�B�'�"�'���'R�'���'��0���H.]�E�|�f�p��'v�'�B�':2�'b�'���')>L���i��}U�93>�@��'XB�'��'���'�2�'4��'VzT�w� _b�rc�_5$��\�S�'("�'���'���'I�'���'&�AYs��;={dQ��"	�:����'�b�'[��'�B�'Mb�'��'��\x��ټ**<�b��7eӸ�j��'%��'oR�'O��'b�'���'��.N`����R�
�1���'��'���'���'gr�' �'���។B����$(��6�����'�'�"�'���'�B�'�B�'d5r�Ɂ$�z��tf��fΖѺ@�'���'\��'��'��'���'�](��LA*��\(0iz��'v�'UR�'�2�'
��':2�'xV�s���3%��ҖE�!t�8	s��'���'""�'���'�bno���$�OtDB�����1�������dy��'J�)�3?��i#��wߛ=�Xf��^1��O	��������?��<��#ظPrŃqtP����9��e�'V򤌃v*���hͧ;��D�~�w$؃p^Jq"V#��o�&����\z��?�)O��}
�щ?��h:aY�(��app��5(X�v��͘'`� nzޝ�BC�"�B�D }�:$���ɟ`���<��O1�4y`��s�v牝�x�;է��ڰ�aG])r�R���<���'wԑF{�Ow�JZ�w��)华!CKB���ω��y�[�(%�<
�4Y��<a( �'�ޙ"�	�)4�����A���'�0듇?!���y�Y�X�'	�8pVG��{��zTk$?Q��`U����Vm̧`T���V��?1R�L>+C��!���=yPmR��G���<Y�S��y"OQ
>ڸ�G�3��Q2�U��y��c�x��b���jܴ�������>.f P�/��.�L(��޴�y��'���'�~Yq�i��	�|�'�O��2I�< y��BF��t=NBN�Iny�O�2�'�r�' �'ѣ�cՉ�2=�h�zR���M;f��0����O��?iZ�HF�;��aѢ�$�.�r�f�2��$�Of��7��i��f7̑ &@ˇ*U�q)J�}��L�`Ll�(I�'P��z�G�F?�J>�+O�<�G�Є�2A#%+� �p���Oz�$�OR��O�i�<�Ķix(\�ܟȚ�H�0'y��.���ꣂ�|Jڴ��'Μ��?	��?A��� Q�
���� $#�ypQ��z��ݴ���Eu$���ǸOg⑀E��Xs� ���mC�L\�yB�'�R�'�"�'_2��^�Uz��24�##추�a�3]����?YS�iN��OH
q�ԒO�`�qH^����z�$��r��� u�+�$�Ox�4��	�%l|Ӽ�-X��f+�CM���!���
1ēe���I�����4����O��%/$b$2P�?Y�b�X%FC	,����O\ʓe��AЇ(��'<�Q>y8�cP�3X�l�0$R�J�D����"?Q&Q���%��'|Vv���(����d��.�g%5����b�*��4��PH��t�f�O�����Ø���@H��`eȄ��OT�d�O����O1��ʓ1웖٤�Bm�v�� y�\lYd#Q�q-(\"��'u�+e�z⟸s�OZ�DD{�RAr�b/D�fL`qR�D�$�O����e�"�P�@���k1�S���H� ��}�m#�������ty��'���'��'��^>���ЎXrv�j0��/��NK�M[���?����?	��$Ez���J9ly�5k�oQ�lP|���GL�7vn���O�O1�$��s�o���I�%�ĸu��A�h\�7N��q�	�[G�)�OF�O��?��^��ԊZ-�Y��/ϙ�����?Y��?A+O޵o�:`�.H��ڟ(�	�@~�y�$�@o�ۥBL�i8���?F]�L�	g�x\�%q$�C8�fi����`���'?(��!��%�f���$a����'l�M���:�+׆��"V��p��'(�'UR�'T�>��ɍ�zXhUK����H��eG�N~��I��Msȋ�?��3��v�4�h�!$Z�@�@�1Ӄ�.x&H�C0Ob��O�Ğ�u*7�:?Q��	X ��)��^���#��4r҉�����L��M>�)O��O���O.���O0��0�]�>���X���>��9�M�<��i8�Hu�'��'f�O��Bs�8 0��ֱg���
	O$ꓴ?9����S�'W���kPiY5B��ɡ�(>{��#�&Ã�M�'R���3��56�d-��<yvf�(`�@����*m1@���Ӈ�?A��?A���?����$[ܦ����<�w��@��|���^�]Z�96`�L"ܴ���?�X�$��`y0������
t�>x4.�v�,!
0�i
���Ob���N]�����<��'�� �Qbɐ�I�j�[�-�=(N��{?O���OD��O����O�?��I��z!���LZ5G����"(�zy��'�7�	3>����O��ny��/@�>E�E�,c��9@�GȰQ��&����؟��w�Yn�\~��O�n�ɓ��~��@W�ۥi�V���ޟh��|\�������䟨�'+I�j~�YB��ٮ��FE��<�	cy��kӺ@�D�O���Oz�'O�`�SP�Y�pR	�-�wn�P�'���?����S�ą^�|�������Q+�/��}]��\ZԱ�ܴC��i>����OJ�O<,�d/; r( ���5����O��$�Ot���O1��˓��V��4Xf�0%ʓK��;��(j�0%Z��'�R�n�l㟐��O����h��c�`�"�
�!Ӈ /�h�d�O@!Zvld���a�,x���?q�'Z|��7HK�d[^��Ì�59��y3�'��I�p��ܟ��ܟ$�	l�4���;��Y�F$�8:�48RE��h��7�Qր���O��$0���O�nz� �F�"H*��ᮊ�
5ph�M�����?�|�'����M#�'��c4É3,��'X�����'2��13� ��P��|bR� �	џĨĠ�:@�����V@R(�ߟ������wy��f�̘@�O����O�AkPm��	�D�!)���a9��(���O��D'�d��'�,c`��H@�4���U�0��I%��H*���Ϧ��|�D ��H���C��&Nw?��B,�vp��������П@��H�O���\�rpʐ��#/�vA	�K�g�(o������O���G��)�?�;,��<��!�a�̉�iC= 3D ��?+OX0� nӲ�|�Z�S���<kšJ L��YK*J޶�K"͚�䓚��O ���OZ���O��D�"?�6x�RA�"K<x��l��AN˓=˛� �g2�'���	Q42��t��hϘTc��$���'E��'�ɧ�O5�, Ȓ�H���P�ό�^�&R�� 2��v��<4���d�����sy򆃹u-|ɧ�Y�@�w�}P��'���'�O剂�M������?� ��$�ޥH1��"��)s�5�?��i-�O���'��X�{�DՒ�(s���{�>xY�ֈ���l�w~�e�=[�����$m�O���[�<洜�WǕ�?���!�#�yr�'&��'k2�'�����wV�<�D�}�DY#��?X��d�O���OĦEAKy>)��.�M�K>�R*�� �����Ӥu�Jȫ@G��䓵?���|�����M+�O��:!ϔ�m�kFE��r� � �3
V��'+�'��i>���Ο��Ʉpz��Z����sz�9ف�г50$�����(�'�V6�z����O��ĸ|R3G_�ʩZP얭xTZ����_~�E�>���?�H>�O�X�:�Ȓ�_T�5����,F�b���,E���ۡ��4�p]���F���OHmX�&.���0Ǉ�6cuDm��Ob�$�O����O1��˓J[��eի}�AhE;f��8�e�ȷ=��l#��'��
i����{�O4���4R��s-C,��,�3�ӄt\�=�d�۴��9&�&L��'=��˓?h��yc �+L�<��Γ%`�$l͓���O���O����O��|�ŗ�~@Dfl�4>F��ҧ���ᛷ(���'TR����'	�6=�`Ȑ��0^mʅwJ�:f�i�c�O��$<��M�\�7mu�lPG�	`%*͋b��>^��te��V��9(���Po��yy�O�㋹C�rA�C��(m�@q�2��	��'E��'��	��M�2%߶��D�O��q�Df��/�8���IV�˝b&��0��Od�$�O�O�T�3iПP9F�[wNX�9\h�晟�p��\�#�xl���RF��	۟�*a�%S�p��G�����ـf���|�IΟP�Iϟ�G���'N尴`��zI��A*B�|�'�'<V6�I6Ѧ�d�O>$n�N�Ӽ[��)/xmcw�	i`����Q�<���?���
Q؍��4���p&�yR��n�L%��˞�QYL`p�̍N�(�4�d�<�|�<�"�D+9"$,h�!ЏjC�U�]~��k�*YIr��O����O��?�j���3<�t!��Q�fN��fa>����O���.��@�o%P,y�3֎2�X����`Ւ"y��c������O��)L>	*O��y��t�{We�n�x�+�'�D6��>A��d�K�i�
��n?�)�嘸e?T��S禥�?i�Y����韠��@6�sI�0(��a$$5��`ևJЦ��'��@�EP�?iR�����w%���A��9_P�2�+m���'�B�'�b�'��'v񟰤��ᚮv? $��d�#v.�c���O����O��m��\���Dq�4���jёu"�5�成��� S:�l�I>���?�'&Ǌ�[�4����ztZ'`+.A4�P��&H�VTxQ����~2�|�Q�H��ٟ���ן�A% �so��Z@AA|�d���F�͟��	{yHj�L����O����On˧8Ո��� ߾W���-ؤA¬�'�r��?�����S�T���7���#��4.���so�'txySΒ>��Ȭ<�'x����K�I�tΊ��흺O�̸�HZ�J�U������şD�)��Ky�+u�z�b�
��4<�����0�P�R��:���O�nZ_�(��Iӟ�(f��&e�^3��ӗe�R���#џd�I,znQo�o~�I��W�N��'��� �@"���!��J�(݊0���:T7O���?����?����?������Y��j�%N�:[HP1/t���lZ!����ɟ��Iq�Sɟ�:����V�@6{����L��F��eCQ��?�����Ş$\j9:ܴ�y,Z�d��	`��͔��V����y"�� g>�������O����)k(�bЊ|4)�@lP<!��d�OH���ON���^���'��'�8��>|��yA
V��<����$Qf}��'<|"�V�>�����Ҩzؕ�)>��䛥F8�8��t��c>YZA�O��$�+`ޘ��gV�D��VB�"�B���O��D�O��$'ڧ�?� D�U'�)���0GLX֏�?�t�iu*���'���`�4��7	^h02g�*<���q㋃O"��ޟ,����4��Ѧ��'�jd��SHJE!�i�����V�����D����4�0��O��d�O��ճnKT����m��E�g�5@<�˓`��F�ǨRb�'&��I�!��ٚu+��+@�e &�'���'ɧ�Op���dת}w|+i:_"A┍�5vu���<�	'd����]�IsyB��W�p����6�܁�nN? �R�'���'��O$��&�M3�*_���Tśu\f�2a�U�+�2�@2�V��?���i,�O�q�'��'�#�&]
���BZ!<�Թ��*],b�(�zc�i��ɫt���@�����I��@�]�R�� ��'�l��w��I�D�	ޟ���Xy��I/2&���$�_8^Of����M�^�R�'.�gn��8��;�H�dN���%��1a�4�։H�J�C�J���_�I쟔�i>݀���Ǧ�'zL�0�hY&�Ե� i� 6l: �����ə��'��i>%�	ƟH�ɶp(DY"�0pn�R5�@�P���	Ɵ�'d�7��. 8�$�OL���|ztK��mUhd#���?{@$�%	k~Ro�>�������L:a�}�7�G�l�޸��k�*�Ȥ�w�Ұ����<�'O��$[����pX���(���#���0��?���?��S�'��B���Ó�<ui�;����E"���	ן�*�4��'�ꓜ?��%�$A�����l�:w2���
���?�k��Ȃ�4��$P�V�4��O��	2�$�{d�{��(��IP�i7��I|y��'�"�'�"�'W2X>5Q��"X���	���G�����	?�M��ٗ�?����?y��d�l��N��S����s�Đ �ص{T���OJ�O1�d%�Fiӄ�	�;fb]i�O��>��c«ϰ6��払&�4��s�O�O�ʓ�?)��Py�C�Y's�yI�{�����?���?Y+O��l��`����۟���>6O�|ʦ`���	��&��H���?�eY�|�	u�E�������2�@3�&^�;�H�'e�݁��{7䅘$��dB�ɟ����'^^�0S�ӱ5�����[����@��'�B�'O��'�>q���@�Jt��nˠVH8�cӭ]����)�M DB'���ᦱ�?�;	$�����7ȊA���3RtP��?����?�#����M[�O�=:������8��3��߾V��}��JЌ}��'����0�I�����������"̪첆�@,G�RQ��OC�ŕ'��7��sy���On�d6�� ;�Q#�/ɅY0�"oL+�
I��O����O�O1�b5q(E�f��E+�#A�����9��6��^yb�ح-rʉ�������	@��<kV��Q~���!F͉w����O�D�O��4�pʓ	p�F삭��؍6��<����4���b�gL�
$r�i�P⟘Z�O��d�OX�ā�Ze��BFJYn��G�|t��[E�f���/T��	0,����>!�ݖ;N٨��٠�8�*^R���͟��Iٟ������O2N8�VOB�{ml8"n�&��M�b�'�b�'�V6���sP�	�Ox�l�t�"\�c.1WQj(ZB�B�Rb�(�Ioy��;U�6��l!�FP�#-¡.�V���F�> ��ص��"(�lUJ��~y���]z^	�e��E~Xm�w��;y���rݴ~�\}I��?���Ƀw6\죠`�T�xc��s�������O���%��?�K�o�8h���!(v�m��CB��6Hz������B/O�3�~�|�:*5y��T�цI�*9)�B�'�����t�'���a{���1+ n������
=#�%�?���ݟ���4��'vz��?�E�HjI&�cL�#+�ŉ����?������
ش���[��F�������hP�������Q�i,�n�IQy2�'�b�'b�'0�X>�Q�Gn�ٲ&D��[M��Ȱ��M���ƻ�?���?K~���7��w%b �M۱!���9�!�#��$,��'�ɧ�O�P�j#�i4�#GQXY�+�S���I���g��k��]��A+�O���|R�tY�����o���jΐ�`�� ���?����?,OL%mZ�jp1���$��88�*�b�ϗ�R�t�AO��9n��?�FW������T$�`*��ה��E�ª?�v�Ad# ?��EP)����ٴ˘OX�����?96�R�h�� ��.O�]g���S�!�?����?����?i����OJ`g��IŔ@�"Ĉ�X@�%1�A�O�	n�FU�����@1�4���yG�Х���46^�r���$X�b�'�b�'�b��-��֘�@����:��� ��!�]�p <��b�0�8yl,�ĥ<�'�?����?I���?�p �5��`����ܺ���Ā��d�Ǧ����ݟH�	؟�'?A��5�$�I3�	Z�Lu�B�<#M���O����O�O1��{f��W�P ���׸:�|�-I�.��7�/?�a�6!T��IJ�Qy�V�D�uSeC�Ff�Y�r�K8o'��'���'@�O��MC��7�?Y�
�*n�h	���V�!r��bG�3�?	ԽiS�O�i�'���'n��ӡdVv��Q#��������M��kֱi���:d6��$�O�q�z�.˝.��8k��<l�h\J?x���O����Ox��O���;�';Ţ�\~Ϡ�w��g8���I�d�I��M{�/��|������|"��4k��{5�ޫ_=�`��J�'}�����F�R?����ag�ZwW  ҵ���| N�s�e�/s�4�x7�'Ѹ�'�������'���'�����Dn��:C��EFf�$�'<"\�ܙ�4!�z��)O��|jD�w.IXu�<
ݱ�Mg~��>����?)I>�O�
t�5�A�T�H�n�
fR��s�@_��HA����4����	h��$�(��$$B�hER�}̍,��c�-�O���O2�$�O�i6)��8"Я�<���i-�Z2�֍*�T-RW��!v#��i�aU)%`�	(�M3I>��w,�I�cԡآo���2*��!��"�۟@�	S�nZ�<!�Aߖ1Sj;��'����DU�r��Mg\4�'����0�	�����˟��	H��o�x��a�/�-�J�eW Yͦ6�7��˓�?�O~Z�����w[�@9B�Վ=�@��̞80�Tċ��'��|��tI@ ̛v2O(����]�L�@�ƈyR�Ēs3O�M g+��?�''�D�<����?A!�H�miH(ҧ�M�\��xdM��?����?�����Uʦ�b������	ğp����/?�~���;7��	"K�V�F��ǟ�I{�˞5r�h�w�,l���8��%��Y�2M�q4��M~J��O Թ��5F��@�\3���S�i~.����?����?q��h�����`8]�ǈV��KC�)480�$�Ŧ��eO@ӟl�I��Mk��w>\����(�N�pK
\��)c�'���'����=��V��В�׺~���Ƀ6�p�C0�V0Y<m)��M�+w�O:˓��OVp����$��C�E���1V��P3޴i�ɚ��?���O�ѫ�?k@j��D��5#Zީ襎�>��?�J>�|J� ��h1�&/ 7qΞUz``&Bpu��ɗ��򤁁 @� ��Zڠ�O�ʓ�J%2gߦ2H�!�m	0�pJ���?Q��?y��|�)OrEnڴZ:q�ɒ_C0�K@B.��I��I�/I()�I(�M��/�>���?��>7�$��BV!D��8��ȁ�b�*�-�M��OX��DH���(���W0l�4`��%�Y���3&���IV�d�OD�d�O~�D�O �d0��U�ݨ�����2��o?T�	̟��I�M����|���4�6�|B�P�Sn�pb(E�.6Lp�e�@1I��'�b���Tl������+T�Ta���J��Լg��[%�Y�_�����Ot�O�ʓ�?���?Q��f�q��)��-�$�;�z�����?9+O.�nZ@j�h�	ٟ\�II��O�] c/֦J6�#�KB;���m}��' ��|ʟ*-@ԃ�]ح��N�m����^=�YCb!ך(y�i>I���'[�L'�2Ӈ�%�H��&�4B
�tJ���Iß4�Iɟb>��'�L6�8}�̀K��"=��۳��8A�ptN�O�������?�_��I�s� �@����p�~���˟�&Ԗ'��՛�i��	oDw�O��ܔ'����K؝4�H��	C%nĥ��'����4���x�	����^��$�X��2dò�K��ˑ�O��1!#�TǟP�	ӟ4%?]����Mϻ:�4x���3�uiǻ�Ex$�R��<�?�|�&��M�'e���'�J�W=��U �7{6��{�'���x%���h���|rS���	ПTX2͝���#�!�@�q������՟���py"�m�����#�O����Oر� ��4��Ր�	�V<���<������O���:���:ra �p�a!�a&��Ir��p�����|z����|�	�s>.�C�%�('��yt$��c�@4�������՟��IY�OY""�n�X9�"�<�ՓG� /B�}ӎܰ��O��d���	�?�;'�8u:eML� �`�ÈY�̓�?y���?��	��M[�O�Ȉ[��R�9�t�0Ή�g���V�fC}�I>�-Ov��O(���O,���=vl�OL,X<�\`J���@U�4,��b A��X�����$?U���C��3f)� �ԙ�?W,��OD�� �)�*}��À�ϲ!���^��"�����0	4}�'8t�&�0�d�|rV�hS�*��S��R�*�}V�jf�� ��䟄�	��OyAiӈM����O� �!]��(f�!0���G�O��m�Y�I|�	ܟ`�'��Qc�f)_�*��V ��
�l) ĵ2�����SҦ��|��ʗm�����K4P�h�9C�&j�`�K}�D�	ӟ�I��	������&ũ
lxi%f��*~�ِড়6�?����?)�i��mОO"�l�ȒOȨ�W'��~� ���#GⰠ�,��O��4�x���{���3�P�� \�C�a	�7��\����/=�]1$����?)#I+�D�<ͧ�?����?�ġ�w� h�K�@������?����$֦������\���ܕOl US�C}.ruyE�����O���'����?�	�C�-�<�I�h@o!4l� 힚`
��ÄAM�D�*Ŕ���OSǟ ���|2,J8&'*Y�h��0���i�k���'���'���4[�ȋ�4�zty n�0��*�kO�I�X�a`���?�����n}��'~b��dB#TP��Yd�)qaB�z��'I�
[��F����5TD����+q)�	bX�m�`hK�J�FJ�#!Yz�	VyR�'���'	b�'4�[>��$�g���i���W�h�����MC�M���?	��?�M~����w��t*&Ë,E�G�	4Y������'R�|��D@6Sқ�8O�c�!A�x������'Y��Y�>O�[�	��?�e�(���<1���?�* xp�A���ys�U�3����?����?	����dΦ��蟄�	ş�)#S7�j�!Ə7�:a�@^��D$�I矜�	I�	�b�~|�m�*|`��&����!T��@��\�MC���y?���>	XR�Ս.*�e��RmV�}*���?)���?����?a�J �?qbD]�q�씳lވp�-(b��?�ƿi2<Q�'�b�hӤ�O�9�h�x�D�AxL�b�Qg �9OT���O��Ď�a��6�{����	;��h��O*���u�
W�~�+�!,��E�e�i�IayR�'m��'��'��O�:@���#�;l�*l�ʛ�9��Ƀ�McQ.H��?i��?�I~r��5�b�H���,H+�,��ōH�\ҁX�@�IğL&�b>=I�d�@狞��U����E.Шm���|�)R�'6�'��AvȨI�$� ��l���C�h-����۟��Iߟ��i>9�'L�7�16O��Ĕ�p���iۓ`�lh���YSJ�$��A�?A\�X�	埜���vV�5XxU��S�$�ș���ǦE�'���"g��?�;f���w�4��Dm��=����-ǅI̚d;�'���'���'�"�'��,��bkʲ!����(��.�Ȑh檲<a�K�Ɓ����'�X62�$����"���b���lY"��O��d�O��S�0��6+?Aृ=#Uܐ�VIɟF�<H֮פJ]��CBE�O��aL>I*O���Ox���O�H��O�����M��b��  ��O���<aƷi���cF�'���'��ӌ�<\�W��m��6J@�0&�8��IΟL�IE�):S�6iFL��:^��`04��3u.Y!2b�&�M�C_��g��7��t$D4o�0��a�ׂ�ti����Oh�d�O��I�<	Źi��Y
�A�jdf��ČM&���ҥ��0R�'��6-4�	0��D�O�t�%�N�F��p��Û/��B���O���:x��6m2?�Ӫ[r6���*��A_4�J �F�>���Տ�yb^� �I������|�	ϟH�OOv���C֝Y�6����]�oMr���gӶi!��O��$�O����Ϧ�.&��X�
����R�nU�A�`��ҟ$$�b>U+m�ڦϓ1��jv(1f]n���JM=D��f����e���%�`�'j��'��蠨�eh
�c� t %��'�r�'��V���ڴK0�.O�$�:ؤ��1��.i�X���bGL�x9�O����O�O�!��#A�:�R4�[�6g��9כ��h� X�k9���n%��'k<rn����@�D;$fܼ1�gX݄�s�����՟��	��XD���'P��R�&� �4�ش,���i��'ZR7�,����O�m�W�Ӽ;� �%0{ְ��)G�!��=�ǋF�<�����ǈt�6 ?�߳z�b����KI����)�� P"��uO�,C�v��N>�-O��$�O��O����OzE�� ��C�@ ��X�����f̾<���i��h�TV�t��I�����V���X`�D �9;� ��������O��1���QF�$�Q�%L&K�ڰ�늻#k��)GOp���ws���'ꒁ%���'LD���+M2o�\��!]�0m��q�'���'4����dY�H�4<@��Z¦DZ�2><�`��YX�����m�&�D}}��'r�I&���m������H-��T�צ��'0��x��	�?U���w��4��]�hN&�'
���d���'���'�B�'���'~�2�`Ef�+
d/�42�y�BL�O����O�MnZ!P��S��\�4��o���&�T�]>��C҆�pf�m	H>A���?�'�2��4����zq8d���6j���y0�B8RD��G��~R�|2Q���ן��֟�ɔ��:I��9�d�ڗh�(��OΟ���@y��N�d#�����	՟8�O�p҂ĸf��H���}T�	��O�y�'�B��?%C��_�b��q��,z�ؒC2t���i�W,핧����h�$�|��X1����B���3A˫E��'���'2���[�@ ڴYPi�$M
�B�LY��O�!'Q�5��ʊ&�?!��U��v�D�}2�'Ӹܚ�$��(r�P�rN������7�'H2��*����(��*�7�Ĝ~:W�ٵ3P�QS��U0ޘYSkD�<+Ov���OP���O����OH�'�� 8��M5<�5���@��+��i_rE���'@��'2�OA�`��K�C����G�E�2�ASջ&�p�d�O�O1��	IB�x���)� �����$g�v�f�#hD��;OnH�T����?i�f$��<�'�?�f	�+lSQIA.e�@��Eֲ�?����?	����Ѧ��W�H�	��4�2�_XaGH�V@QϘq��b��I����o�	�EO�`��	lbd13�O9�J��p�z��$J�"O~� �O�j�.����)O ��Z�ꈸ:���c���?q��?)���h������.�CE!����i�B	/0~,�dD�%�ҦS��,�	��M3��w����V�d���#]�[�4�'�RS��"e���!�'<�}���?��D�v�X08�JB�.�6��Qe�	_0�'��I̟X�	�x�IܟD���%u���$ �2 �h��� �*��'7H6mִ%&�$�O��d �I�O��
��ԧ�RX��X ��<��Cj}��'�O1�Q�ÁM�����X�<����Y���𴈱<�ƇL�b��dӢ����Wn���+5ha��b�B�O����O����O�4�Zʓk��vA1���AV0b���&0>$)"�]5�y�e���|X�O��D�O4�D�+fQr3%��.V横��6���5�aӊ�W4X`�E�?�%?1�6/��T�v��~����]?Jj�	ş��I͟�	��P�	P�'(LNq9 FοyP@ 㗯�5Q�tԢ*O���Ys�v>����MkN>aqgEq�z����6I�m�bj[D̓�?�.O~�{g�z�\�w:T�CV�b����)W�d+�e���#��O���N>�+O����Od�d�O}!�'џ./�s�f�y�~�	��Ol���<q$�iĔ�#�'�b�'��ӭr�HH{q����H;dL�3p�~�5���\�	t�)��	:�X�{��U1�j|H�L_�z,p!c�(=�JM�*O��������|2�W�&u�=@�T�(�FU��̗sb�'Y�'r��dZ����4NDt%���7��(�7��@5�=�B�H"�?q�T����$�|}��'W���kȯ}��J��]?s��]Av�'��+��0)�����n���t�~��/��X?�ȩ%��q�l��4�<�-O��$�O���O��$�O��'l��@���BPK�9�^,�3���M�A��6�l ���?���o$�r���?��Ӽ�w#� ����TN�=]���H�O� �?	����|���?�P���M��'�x۷h�R��s�g]�L��'�VP��	���y@�|�U������D��H"�B� �]���ᤕݟ��	���jy�!z��p,�OR�d�OT�J1e>56ܸ���:M���%�	3��d�O���$�N@�lP14�R�~�${u����ɥ~��u�+F;�$?=
q�'1����r�PD)e$�'z��p�L��!�	ݟ�I�����n�O��*˓n�ʑ	�*&yƸi$�ݸ&�Үt����֤�O��D�צ��?�;e���D�$��`2铢w{�͓�?A,O��vgvӢ�C�R)*�����C�O!
~)Iv!�8�D�Y����������O����O����O����)��:�K �XJt��6l��ʓK\�+��[~�ٟ�&?�	�K_&�s2 0q>L��aԝ,�Ҵ��O��d�O�O1�Е�`�x4`Q��H�K�K+'r,A�'���2��SVKOTl�	RyB� ''吭ٓ䂶G�f�Q$l�~b�'z��'��O�剮�?y��͟ ��g��i��X������$HП���4��'����?���?Df>La���fi���Qkvcލt�v)�ش���ٍn7����I��q3Ɂ�c ,a�oŢp��Qq�2O��Ċ��ʵ@T�96G�܂2)��0����O������(��!��iV�'ɤ)�4�	2[ڡkp�@�B\}Q��|r�'L�O��+��i��	2iJ2u�P������c	@e�.���)�$�<I�bB_��~ Af��H�X���ͧ�O�l��w4T���џH��N��2I��j�f�B?��9������}}�'H��|ʟ`p�6�K3F�$��C���F�ҭ��G@3�s읪:�x��|�,�O��K>�s+�
�rN��.�le�G�^<Yr�i^p�3���td�g
Ĭt�p�% ��9���'�N64��*��D�O��֧_�5�h�+�.W,�����*�O��d@��7�%?�k!��Ay
Y ϲlH�#�>�dX��Kޏ�y�\����I�/��A�؄V�z��OՓm1����4�|���?���O�7=���JA�,	��r�
R�5�8=[��O`��)��i�P��7�|��J��_)h�%�$}�I�k���JQ7/d�ݐA�T�J�Rp۔��2_���R�
p�	��[D�$�'~��A�!@�=o'�B�	EA�` Bg�//n<R5�_5j娴���9B��R�G.Hj���b����GO7Ah ��V�Q�����<���B>H]"0Ɠ*$8�Q��d���$�"w�"3V/E�A�P;u(�̠ܲ-au@R�&�3��H�(���ls��A��_%Ik��i��+�b���EY>�>�,�Ty ��VqT��'s��,�|q��Y�6��]�l:O��)��.��p۴�?a�!z	��jƼg,ِ����U���i�|��'�r��(qOB�˃��2{@Y�DfUu;��2�ie"�'��I�~��EZ��*�d�O��)"`\2)�	ٟ#�n��E*ܡ5�U$���	��T{��g����t�P�;h�9Y�5~����P�̼�M�/O��r�ƦE�	��<�	�?=٨Ok,Vu��ye��"\H\��G�#ᛶ�'��֙'b�|bT>�S�? ��
�Q�`(s%Uw�A ��i1��a��{�l�D�OB�$�nu�'��	"P��P��H����ЯZ���4n�1`�"�	�O(r ,̤'���s�^4��� !K�9��۟���&ߤ@�O�ʓ�?��'��U�"ڴ�Er�)L�&4�J�}ҋ���'���'�BM�6_�����I[�2�!�ak�i��7�OH�RTƙr}�Z���I{�i��2�W�N���'�W�,�x#��>��kE���?��?Q-O��&E�6 ��q5̓2�y�R`	R�`�'�����%������`�B�e+�f݉E��9!�-�%�$�Iϟh�	vy,ۻ��Ӌ\�<�i�*S�	o`���>)�7�<q�����?y�{�yX�'y`������z�)!�	?:���O$���O��ĸ<�d&@�E&��😃ecI�Ry3$B�_�]��J��M�����?������>��nD={~Hm�Ęk��	5��ئ������'�:j�̾~��?����Lt�'cǫs�&����ڿKKZQ�Ӓx��'��Gݐ*��O���L�z}[�f֡M�T����;�6�<�!Gݎ:,���'���'���>�1;�ZQ�(�QT4��A�J�@m���I�u����?Ɍ�-֗\����ᅝ{� I�Q� ,�M�vl�?a<��'��'����>�,O��� E��B]��K�>#�F����Ԧ]��/�h����O�R���ɲơR�[��S���Ȃ6m�O:�D�OZI��P�i>���H?ْ��r<}��ŤF5��#R̦���g�	���9O^�D�O4�� SpX��G�Y������-*�l�Ο�Jn����|�����VXxY@��s(�!#զæC�����x��'��4�I蟬�'�D��рʮz�rX��h��3�SQe��Od���O̓Of�Ӻá��x�� ��]�"y�%fH�1��e�ɜ��9O�$0wc��8��.�-|M�8�a 1?x7��O���!����4�'��|8�4�����K����q!Բ̰��'\��'��]��%$ �ħ*��X8`�Z.�������4��q��iGr�|�S�����*��*��u�vs�jX�#�����i#�]��I
H���O4�'A�\c��h2L��P�ňȼN�Z-�N<y���,���] 4"���BƉl�`���P��7m�<�b.X��i�~J���b��x�{V6��d*G�tQ�$gӼʓ�?y��29�O���MK&RE9�0Cm �w!����BҦ)X���M���?���T�x�O�Z��Ԡ�x�L�]u�\cFJf����O��.��?�I�P��⃩�ƕ �@�<r%��
��M���?!��(:�E��x�O�O���Ď�t�Z��#̜z���5�i���|��'��	ݟ��	�֘?T�X`W��`nZU���Y
��6��O���̐k�i>��Ia�'6�E�Oӡ*�
H�CZ�,tK<Y�����?�(O8�$� �ʁ�V�W�a� ����'s���ꢎ�<����?)�b�'$�d�MXJ�@&�!
q�4��c
�͛V收�'=RR�T���p�)��Vi(1�����S|���e���9�I��p�?�����$)���ˇ(�	a�� 
h�� G�!���?/O���Ϳ]��'�?I�[�\�jp�Ӣ�K
�(���!����d�O��4�
�%�LP3�#��DӰ��0��ct�s�z���<���C���/����O�����E#��H�N�tP"�K"#�:���xR�'G��>K��"<��{*y�gC
ul�@V�:Ij�oey�B�&RE�7�~���'���
=?�愪@!t|�v��

�ES Jঙ��Ο����dL|���iBP�Wc�
��lk`CE�Ul�ɲشe=Ш����?y��?�'��?�WM�`3~x��)��������wh�b>����`J>�Zwh�1o\i)e̕�-+�X��4�?1���?������4�'<�o]�C��r�BMA2����$�s�Z7��OP�d�<�Z?�?y�K݊e�Ss�Fi�`I�_U2�1��iy����*O���O��O�\D�A�$˄9~1����iЗ	�'��W�(�I� ��^y��66�Ti12H̋Y�Llh��+A�B!jS&5��O$��,���<�;+-�Q!l�T(�e01�,J@"�l��8&���	ay��'(�$џv����n0�+��L��iY�'��OB���<�@��)su�͐+؞Cï�i��ʠn�>��?����§ci(��O�b�"3�+@K��A���[>O�V6m�ON��?	��?��*�<aN�\j':���4�C���*��dӊ�d�ODʓQ�1ˤQ?������S��E�Ί9�8��H�-_Oΐ��O��$�On���&n����O��$�O���<���2pJ�1�8�(1$��6��<Ӄ
	��v�'�b�'��d�>�;k�>�Yr�� d؅�`�&u{fn�ǟ0��`N"�-��9O��>�D
�M�jE�Uʓ�I�(W p��q�i���	���I�?M��O��A\0�L �P�Ҟ��	Q���<3Ǜ6�^$�y��'��'���*[ ء!�2*���&'�4,d�l�֟H��ݟ��Ԧ����$�<A���~R�җbV�q����t�d�S�+�M����$�,k��?u������� >�$/���8�2�sQ�i"+�;ꓒ�d�OP��?��FT�	���[�a�\�RJ#.`bi�'�\��'2�'���'}�P��׍E)��Y��Z(xh+���i�Z���OR˓�?�-OP�d�O��L:F��a'�3M��5�����4T0�0O����O���O���<��-A7y��@�}��prbܿ�25�WE?
�_� �I{y�'O��'�R��'��|$�ȼq��c���Yw�~�f��O<�d�O�ʓ@.��R?��i��pTΉ6&ʰI�:��:�$x��$�<��?)��G���OJ��zJx)g%GB8*M��풋&����'�RX���
�����O2����)AD�7H����F�/{q�X{w�Xs}��'s��'{��)�'��	���'����J�a�x�V�G�Qz��mYyR,�\7��O��$�O���Bk}Zw��e���l��-���#a�Y(�4�?����'��	bܧ��t���K�	�茘� U��am�->\5��4�?����?9��:y�IDyb�~����݇H<�y@��FCN71l�D ��0�Sޟ�r���q�z0Ȓ�X@�-�%�X��M����?���1l�K�Y�0�'��O��x�IAYĩY�/R	�P���W� �'�
Ԓ�O�)�O*�D�O�a��nZ�VO~|��j  Z�`�� �٦I�ɥG4X��O���?A/O����<�kq
Jp�	ˆ�8qJ�	Q�U��i��q���	P�I۟$��yy��	_�p��&Ր\��
a`�T_X)�� �>�,O|��<����?���8T�𥉗�~D�bk�<>o@qT��J~"�'F��'��_���U����4�Җ.Xy����'j�$�"�X&�M�*O��D�<����?���*�$�OS�T��ZJr�[r�N�%�"���O��d�O"��<�U��H��˟Pb��*9���š+;|��T��5�M�������O��D�O�@+�8O�����`���É_;�bv��5}�B�cy�$�D�O,�y�lQ:�Q?y�	ߟ��ӏ�R໡��-)�Z��]"�CX�����OX���OXi�4O|���O��D�?!��cH�I��yʰ"�xS�d1Wip�x�q���;��i�B�'�"�O��Ӻ�b��3Q��=���B�yrB���l�ܦ�����ˣb�����"���xs�ˆG�J��N.~b�7�@6n�qm������؟P�����$�<��fW+p#J��rI�+(�~岥�P曶O��y��'���'��4��ۈF-Fp���y6%��"W�YK4�nZޟ����D(bK������<����~b��'�:	k�j=r�]����M+���d�x;�?9�	�Vgӎ8��K�|�R�r�UX�3��ۦy�I 6k�X�O���?�(O���ƒ̛$ҕ0���gO���\PcS�L� �,��X��՟@�'k@�qv�P��Ґ+�x�C�,(��I
�O�ʓ�?	,O����O��$�f�fc��d����"�3V��,P3:O�D�O���O�İ<��N�J�ɖ(O�>L#��V�>d�:�b����fY���	Uyr�'e2�'��1
�'��=�S%%����Ȩ1��Ec��qӨ�D�O\���Or˓9���PT?��i�i5��Rp��*Ə�C �b�D�d�<��?�
Zϓ�?�'4�D8� _?�
5X�^>�p`�iVB�'��%/	 <jH|�������A��҈�i��H"G�Ɯԉ'�R�'����'G�'�I
�Z�^��M�^�\8�0L�_ћF[��(�.�M[]?��I�?�OJ`��/�:n�1iQ��=-�`�ֺi���'X�[���%�'[V�J�1HnƑ��)�86867�� [��$nȟh�IΟ��� ��'Vys�"� 8�8�z������mӂ S4�B7�3��%�S��� �p����%-f1 �+6���Mc���?��� mZ}�D�xR�'`��O���Z�p�4@�#���@,0#&�i��'��Lџ��i�O���O��XӨΟ_Z���@���!�!�k�����jSJԣ�}r�'�ɧ5���/ N��аM��y@!����B�5���$�<����?����W'�t��E��1�lJ�~��gb�W�Iş���l�	ş��	�@�s�����z0b]#��@�l\q���L�I��'-�+�oc>���e	�,����E�@Zl�FA�>���?�H>����?��@���?����?C��%����v,-(F�Ӧ[��I�<�	��ؖ'c��[U�%�鐠D�FXXe��7^:(��PJ �<HR�m�П�%����П�f�`��O�P��ӕvؖP��䝂�v�As�i��'��ɱ"�КM|2���bK��f�pRœ�cC�1�)'�'���'قE���$�?���)9��̻EF��I�,=�q�b�8�u�NHBQ�i;*�'�?��'`��IQ{��*p��1zא�O�-F������OT��X8t,U�C���Z :���r��i
����}�^���O^�D��.�'��Ӭc��ԙ�,ڕ(�B�p�D�9@*�)�O��$"�)��ٟ����)ײ̨�kݟJ�,1�"��M���?��z�P����?�)�*����`��-^�tZ5
Ub��_��rQ)ȹ�O��&>e����4�ɶx����b189Ƀ
ȯ^7@��4�?a�CI'Cz�	�����OJ��7}R���>~�EPO3S
���"D��ē���?Y��?a��?�%�{�4���킋z�>���	
�� ��?���?I����?A�'Ԕ��F�i���ӤS>���4�,U�' "�'52�'9�ʾ/���=� h��g�iM��ұj]�vkNdA�if��֟�'�L��Vyr�ٲ�M��i4V��w�S?)XRl�c�KF}B�'�b�'\�ɬu����O|"a���H\k�V>6�f�Q$��P���'����&ϱ��Uc� �o��qBk�+yH&}`��i3�'O2�'��ѣ0V>)����4�S+�� �EM���0��)ڜ��}�M<�����Ђ�i�u�/�!�sS.�C�P֔
�M�/O�js(�ʦi@��"�������'����H͓r��d��ٴ�?���|�d�Fx��Dǅ�1&^z�f�&(<$`SU�X��MӲ(��̛��'���'��9��O�1Ve
-A�H��r�I<8��3@���c��4�S�O@��Vi	�떁�	:z��Y錌?��7-�O0�d�O�=���w��?9�'m� �i\
~��)��߁[Pc�}򨕖��'�R�'�"��v�ٔb�.� ��E�P6�t���$�8^f�>����ˠ��.$�(�+� ·X$b���g}��R'��'7��'@�R�|��.�NeV�fī^q
���L�����}��'��'���'� �X�
�d�ִ���V3Qz��P��'s��'�"X�l 3������/ܷD�*�S���T{�̣S
��ē�?O>���?� _|}���.I�;�ḀS+���b#	��D�O��$�Oz�i/4��C��T�K6e�J�q���l�pu��n��C�\6��O�O���OȬئ��o�����7I?vi@T�I$S��f�'h2Y�8K���ħ�?1�'g���� QB�ܲ��%[��5�r�xr�'�R(���O���KSl#˖�,�H�z��R�-U�6M�<��̕�4��vƭ~����T����a�F$H��2���J�:�x�+j�n���O�\/�b?f\�?|�Q��Ɵ�.�jrEu��Eq��O����O���韠�S��ܜf��`�b-X����&R�q׆7�R!>R����埜*#�><~"d�u$ȥW�LM*�����M���?���U������?�.����� �`I�P�X���.�
�ب@$ͯ�OvY&>M������%b���p�,�ZA�\X�Da�4�?��%"(���$�'W>i��M�C^M��Z!BSv��l�A}�Ɋ<��'.��'���'�r#�	 �U{&M5�0�b��#�ѓ Q�d�	柼��@�I柸�+_�P��ҭm$b�a-U�o�
}5��'ʮ�yD�%�)��.Q�J1ph� J�8s�aƬ��y2E��.=! j�5bŻ5!��'��Ղ�!" 0E@�I��W#d��P�\(� �B�Q���pr����<�ֈ�.q�l�N	"=��� N�b�p\s�gƋ'�l�30�3��@U��0Mg^̘�H8}��TR�&��?���8>���ƭL ov:��AC4 �(}��a�R� ܛ�$,cμ�w��9o�!���=���t.�Z�i!b_����?�J"M*eqrH�#=\<T�(�%���SH�4n���xWiܫ0Hv�������,`BP[�e�!�	0@��ۦ�c,�N�S�m�t�7�ӑ[_�<�gxdJ�'��4y��?9����O��K��`\�*b��&�����"O@U���ϐ +D��BcK�Q
����'�x#=��L2v"E"2D�N/j@��F����Iڟx���-�8���)��0�I����iޝ��	8�̩���@
v��]۠AR�y��r^����:�Lb>�O|�K7f��1�$j���R���"Z�d.4��O��1!靝����ΰ�Еʄ�T�s���E�4�P���D�*s��O�ў��ƅD>{�8�R�؅W?��'�7D�T�K�.cc�dp'(�%0���2�4?1�)�+O��ZFh,m�ܐ�j�?��|h ��d�T)���O���O��D��;���?a�O
LU��gT��ZhW�N�c(�.�p9&�]2e����$؈3A�)A#lp)�
P�R�d #��z&KO؞xd��!_����N�fkPAb	Bf}��D�O��=1��dٝl��[Î�(&W��`�'���yOU�@R�`� Ț�6R�BD���'ɬ���AJ�Y�'��o�dH��U����7�r�'�<{`�'0;����RHF��"�Q����7͇�<^hyÐ�ݞ+���sc�Cc�x��NBr���ɉLQ�)��i�D�P�r!Ň��\e#!S�p<�$�ןx�	HyB	��h2 j��X�8�`�� 2�'��{�P*:7��I�lS�s���N��x�.o�PB�"P�C���# BQ,l�d�#=O2˓yp�}��V�8�Io���'h�%�.F�|iW�B�t
"�����b]��'���0&V�Z)�)A��~*�ʧ~A�a�	��4T��j�Y� ЦO���5�'
�թ	ũ���$9�t�\�y:u�@MS��$M�w�>�v����4=M�>)��]��e
0i��}H��I��h�Ɠ\�� v� p�`��n�d�DD����HOlp�!��X��"�$x�6����Y�I�����Pv�PL�柸�i�7��Ol4�;-�,U)���uY��[4"�ع؊yr�%h<��� ��h]�xD���M��:a��d�D�ȝ��	�`�m�4��6�i*� �S� ����L��'2�]�)�<�u�}��$��TsHeS��:n]�\��'��X���	U���f��Q��y�OTMFzʟ@ʓ7��yx�rӒ��t�ݨ#��TB�'�,T�M��0�iE ����R�'j�����!X�t�āX^Θq	�'��,�@i�w�.Q"�FS?PQ	�'�x�����:����N��=���'�E�P�1Gf�K$%��:ݬ���'�Z�*��G&S�z-)-׻G�P	��'��,9�e�8�%�&c�/h�f�@�'���y�Ąpf�`"�4_ې�J�'��mSf �$P��p��CC�e�����'��!K�T�0��ݏ�*ؙ�'�Z�:s��=b�0R�o�~�J9�'�"�����1uHf���>o��h�'?�n��$>����P�Z3ҝ��'a\]¦��lK���Y"t`��P�'9�I�3h̋Ih���DeTX h�'X<(�'��Lx�� n�1c6���'ʠ�#�F�P�^���j%\xQ*�'��(�U�u�rM��W�Ss���'����#�
U�p����P�^0��',��GG�]������ T�B�'sd5⳩NT3���D�γm>4�'+�0q�ďwة����-���8�'J�U��M�u��ww�`!�'�J�#��H�\hx��F�>��I
�'��,��&�<Dȴl����i�v�	�'�Ny;�鍴Ul�X����`zn��	�'�Riz%�F�P<K�m�$[���	�'ְm�f��j�|s4�HOЂ�	�'=z�1�
G=���ԮCq���'��$*6�0{�����ѳ=N����' A�DB=0��m{���$9D^%�
�'0�-2�C��Gۂ+g���
�'0��b�%�4���	
�m `Y�
�'�0��_("LXg��Z|��
�'�ܙ���A�:J�����M3z}K�'%A�a79�jH�B$y$��q�'g��j�K�fj��Зqoƽ��'��t1�����Q�����q3��	�'�`=33H�}RP�:g!�#3#���	�'����a�4j^Z�1������"�'w(0RW�C_p��H!&�α*�'�~��1��=K�lZ�P}��'J�#���Z��kU=\�]�'�p��GXa��Ё,�1p8)9�'�j�-ڸ��Ȋ�+�IH����yB��x��2�]�0� %�A!�yҀ�}�򹑒�\�+u��)��y��B9qnY�f+�'"�"��QK��y��U<1$Yz)�<�PQo��yr#Կ��4�b��L䪁�ߢ�y�	Ý>���|���:����yrE� Y�8��ơͩw��� )�y�˖�|+S�9�pY	&D�;�y���L��uC�J�6��*� ��y�E�O�]� #����ʸ�y�יa��4:c�мk�P�8��  �y���+;X쩳��b�bՒ�����y� 
�ıa�
�O,^�I�'Ѳ�y��= �B)�`�-F��C�����y
� ��7k��nw�|�V�L.D�)#"OJ����0�2q2�`] �9�"O��i���=	��D�����"O�+2�C/7¸9D�ԉ.����e"OdW
� �:)��������"O�z��I2Uʽ Ge�h�fA��"O���
Ҿm� ��%τ�Jd���"Ob���͇-�F�+�۸_7$X�F"OL4� �42�Zy��nՏLH�V�g� e�����Tw�>���3����7�,v�dj2D���]�.�F K7 N<-�T���S"vʥ��nr��e��~��ݡ>h]����lh�b�)�y��@T^=2v�Q�/�h1��] �?I���!g���p�'jc�c��q��5�`�� j�����^.-���>b���&����l��thY����y��(�E䅰
��xke`�o�]ExrMT�/iة�YD�>����39��H�bٰ�����(D��K'�h=�I[󆑃zz^Q���3D��1,K0tp�7�8H�%i �7D��� ��a��H[7偙sc���J9D�`
Ӎ��=��$���Ӭg)(]�7O5D�Tq�e��E���Ҙ5�����4D�ěA#�|k�ЫƫR�(��x 0 >D������n�	`�N�S�Ԅʠ�1��O�W�Ĥ� �Ы(�p�F��.'����B�F#8y�<�y�,�!m���Yգ�0`(8T���)e�b8��-ޟQ5���'d�^	��Ox��5��0�P��zf&<�fO��%_>*BnV� R��0�Ao��P�~U������`�@za{b�ǡtX���jW�QUL���$���<Q&jV�U]\��a$�^>n6�܊h{���nES�d��+�y�!�d���)XedDx
�K���&-��'p�u��$)�q9�˘@�O�,��C3 �+��Β3�|P�	�'����@j�,l䠅�)��hjѪ>�6\(�ͣ�l��FRI�g�dV!o��,2�L*Q�(��0&_<S�'�8��So� �W�6�上Rɐ�e>���'ed�1��3O|�:�G��G�쁲����8��P�0Q&�⟘  �l�Ѥ��1C,�Y�mW�n$��!�.?����h�{�E[9;�p��jQN�j#��q�Z���zmaB+D�F���%�L7"�Ƚ�4 T����7՘b����,S �+?�EN�?e(x['fR5M�\b�(P~�<y�:S��!��M��Y���i�w~R��6=�"=:�+ʪ��']�<9˟�-a�G�y�N��J�SZFP�0�'��!u�UPm�r�6P�@�"��B3+z���
DQ}N9T�Xҍ��y��ؤ�RP�w敲,�H�Hd��
��Oz�
��?�ɶS��S)TOx��X�*ˋ}���!�呿QU�T�ľŰ>�A�%U{�uZlHE��u��E�ayRiX�%I1O��*�eA�A��4qѡ�&�~b�H-�	��÷n��P��o�y2��-�Y5,۟`��՚��	��d@�_	z���YrbF�XΟ��+�k7�4E�:6���(��2{����Ro8��#�k�J�&mQ$�.|�$����D� 9Y�L�y ���kR�M@���e�p���D�4�lf�@�v�	��+��s!K�&R�69���!�6r��@@$k�#v�Q����R�18��6 z��8d��j
���䈯���pԆ�q2���O�*d���UM,��,#�Zxt�@�O�9)�c�
}�����o��y��W�x�`E@AG	'}�xJWn(�y��F��n4��eK�#"�)㺼��V+C9Rw��ژ5YN�pW��M���#s��?o�*��]9�EE�-�J߶X��aH%� GT���I:�O8�v�� R�y�g��Ty��R��r`a��dpV�SI�w��$GA	gޖ�
�k�.[U{��I�w�R)*1)3 !�1�v���i�֢ś1)���	�P��B��Amڼ���#k�A��§1mФ���àRJ�;�j�<�}��'����*@�S�8Mb���
���h��>+8��6xZ���Ê�Vz��³&X�3.�La���:x,�k�w�4��Hº[V��@��#��PX�'�ʡ�� �]d �e�G-F�,)I7��
���Az���c6ʚ�T#J����!O�d!�a�Wc,(K�w>-Q�J*A1��MH�i�Il�DB_�M��gd�#�E:�I6S��taP!פ\��*2F\�s�e0GP'f��L�cl �B�Ģ<� ���@��dY���*٣=�U #ቂJ�dp9T���)۠�1GºZX}㰣�/m����ʑY��~���-Wo�]"f��Iwt���D'V��p���"6���pO�x�@t`ɟ�I:�*� ��`�p���m�+e��Aҵ��dW���ȓar���-;!?��C��y!"��I(Qr��+�\y�f�>:��& ��	)�y���`F�?7S,��@M/2�)��,LOpI��9B_�tbNB��5	�-�19�����\�$ʢ<Or<�CD\0O� �I6%Q���|�tN�e	�I-X�Ye��nPL���޾'n�b����Ξg�ՀhA�VJ����O�9O�(��B�障��`G�{�) ��i�\�!�+M�wQͪ�g�ALF8S����
�?��#������h��Z�<+1H�-_�"iS�"
�K
68�!��ӟ��g̓�����'L����A��m"����,y���A�}g�On�1�-�Y�@��K�I�^- @`�5M�LH��9o��e�?%?-��!�)	2`�:W�G�E��ո�N��C0N%#E���~b�ǇqJ���Q�� �IH�,R�^������m0͐�2FR�B�<�0K���� ��t��0��?!!@)���$ɏc�&��CHν�h鱠_��1Oi뵨O�Yc��:ra~��	��i��9O�L;!�S�x��$�"�V�d�;�D͔S�:��s�Y���mcaB֜G��m�?�sH��?h�("gBP��OU�u>0�����&R p"U
zqT�[�sӀ�=�OW"����Q2վ��$�L;{�6`�v-øL�
�DXI1��H��9�,l9&� ����胩;ړ.�ƥ�I�Kێ0��i��a�D�x}蕊ء �|���O�c=��C��օZ��=J��&�[<��Q��H/ p��q���4Q�U��5�l(�����t�D�EX�S�ǖ�i�^���C�2^$��9qu|	�N<�r�%9��l�K���q�բ�I��K�m��P�R������VNU;���)��h؝�L0落9�@@�V��1����ۋ{����Ka �pGL*J�n���GX���䞸d�G���B!xK&D ��)����.a�r�g/H�CPd�I�ZJ�.㞄8�-g�g�D�3\��=�e�܍G�q@ؓ+�<�!@ϓf��zPP�4�|Z�E !Ϯ�I��`)��g2>�(�CG�$9�8d����>� �7X>T�Ӥ/(	T�#P�����Ur4�IB�nձ�_�^`�F}��0�!��ݞ�
)��l��x�6^ą�E&1��!Y�'��1jHL��"`���$1�xH�p�ϸg������V8���D
�{��<Ypgv�	�/<T�(�Aj���[���s��B�I����Yg��
zc�8E�(yh��Ut�)�u����S�O�� ����d	a��`k�=�'grM( $$&�2`��!
�CGF�cH>��)��F�aÓG�F�]0�Ԙ��ʼ����3F� ��в��@��hȂK�0E���Z40x
B�	;l&Eг�ʮ+��M8��O�(����$���v�@���ƌB���Q��:��x�;D�P�d.ú&6�Hʤh\��1�c&D���l��od��`V����R���#D�0�BT+=e �ꡋ�4��h�A�!D���Ï�.�q��#Q��� #�g>D���׀J�pa^<3D7C�4xc�=D��)�JI�<ؚ(i�Ӊaw��s�L=D�HC����S@�C��ό?���V�<D�h�AL��,��1��T�~�Q D��K�A
A�m")ϛà�p�:D�$�D�̦,��Q��%D9N�I�.D�� �&�,b­(E-�1a�x$��m*D��5ȂC=��F	�>y�eҖ�&D��y�	]��{�A,�vUk�F&D�<�6a�"�8������Nc�h�L>D��8h�/&��H�e�]
Mzh��V>D�`�ի�t��ػ�LV�sD�"
0D��I  ��'�lم�+CX�r�/D����BH�5B)S7�^L��<(��.D��:T��	~z!T.�X��X[� )D�S*�=6�
�0s�Oon���-<D�8��+�o���{���.8���@�9D�|��ؓd<t��Y�F�!$�6�!��T�Ʉ��Bm[�L�~�㷂68�!�Ĝ�2�̄Y��Ǯ:��3!���!�Zr*D��ꜧEZXRgP-�!�� ̼�h�}�Y�e9nT0`Ir"O�,��[!Zti��ŗ�NK�,��"O��BÚW�e�=C���"O�E�q��o�\����˔TUQ5"O�a5�F�l�.,�v'¼Y\�y�"OB�8"N��B�J���SH�YH"O�$XW��,��  'b�l,
��"O��IV#E;�L[� P�Pv
��g"O�i2W�J�v�Ju�@���0c� b�"O�8Ѓ�0oؘ-J�:L`PQ'"O����[6+`���
�;��"Oؼs���q��&�ΧA�Pk�"OV�!-!f�)��9U�H�r2"O�f��?�X:�BϭN����"O�%"�P*Xj����r��Q�"O��y��Xx|Q�lŻ+�t0�"O8rb� :R�(�ʙ&�Fq)"O�Z�&��;K��WJ	0m��!�@"OhY@5���"8*���� o0b��W"O\Y�g��'P8���2'JP��"O��Z�M��R=���U+s@�H��"O~q�eg�:���z��?Q4�U�4"O^�	�W�e��- ��Ԩ#��yKq"O
��t�8R,�iɡ(�P�j]	"O|�#s��t��#�l��ak�g)D�4���Ηj٤]; ��V5i�j%D��("���D�}�7J�3�~ܺ��&D�� �gX70�ά�#ܕKq�3��9D�*�{,��;e*�45��HrFf-D��#�
E"1I�Ö�<_�`hwk*D��b�F =���A��U�Ẁ �t�&D�t��(x�lH,�`𪀇%D� 9Ũ��6ZĠG�+n����O9D�P��Hd��07DG�f�^�87�7D�0@�k�7���g-3L�q�D�4D��� )���r$j1shz���0D�\�$ܡ0�(�k�h�*�M�.D�ܒ�If��a"�D�0���`��'D� j3�"y�MA�j�J��0R�/%D��� ��,o��,Q
N�s���C�b"D�d�D���-R��eC�1Ј �"D��1�^6j�(y�S@ޏ*W��"D�xp�J	H�He[U�I�Z��
=D��	7���I�,�I���d<���$�<�hO�S�^H8�5Fݷ&t���lC䉬M�.��$�v���Q �N�dOHC�	�)�X�*��uE�ӵ+�� �"C䉅j���2!	)��D�0�Ҫo��C��.H���z�G�m��գ%'�U��C�			T�� ���ҡ�³,�C�I�9.&��"��p2Z�2T�@k�B�	�V�~�P��ј@�B�◪��5{nB��#�d��H�,i��	���pB�E����!`î1�N���`�tZB�	�%��ၕ!Ety�D���G���ĉ/��#ҡܲ����@!J����d ���8�,�B���q��x�<�� �X�F�&@�_[�H���A�<�JFI�2�p%M]�<6���Mh�<��EP����m��)6Ȳ�LWL�<q�`G�[�	A�M�R �8
�HJ�<�Pf�'�^��'$!@��(7*�B�<��m�.@M��hQ�R�vD��Q�Cw�<i��ؔ�����M=����\�<� Je�2���y����p�_CN����"O����;N]T�P�M�3u�Ă"O�D�tAP�H�Q�c�ųL�@�Yr"O���̊�� TA�]?�j<�3"O�PfD�in����C��J�C"O��{�a����b�ѧs��!"O�y��c��O�ܤIԥ��~��$"O�Y��C
:b�z)��G2�8���"O^x!��@ ��\�R��S����"O, �4*J4�<`�ώ%ʼ��2"O���m�8&���ۢ��0_�̱2�"O^��'��.k�X��NP�+��:�"Oʔ�傃XN@%2��Y�ܘ��"O�煣k<�0f�֣(|	9"O>�#�JU� {���2O]�5"�"O$��#D��4��+�J���P+�"O�Q���)�%�����/��0��"O�,��B#Yn���������"O����瑯'x45�f�G�q�PxW"O�;ӣD�,5���F9zs�P@�"O^���L�Y�0�2�n��w"O�M�d�V ��E ʺPR��W"O�e����`��M����a<����"O�B%"��z�rXC�Έ�BM�c"O�͘b�%UM��p��C7��d�c"O�Ui�l�z��҂��5u@	��"O>�Ɇ�ߺ#�(�Hlg���B"O|iP,�
.��s�f�>H�eK�"O �qf'ʖe�5*��X�2���V"O�dl��X���!����"OB���P���o�k�dd�4"O&%�S�B*��f��_~���&"Oέ��)��M����-Z�Df,���"O�x�,� @�p�ȱl�ir>��"Ov�8fN܊���1$Sd��"O8���b`���	�w!�$Q�"O�Ie$�2�r1�%�	<9�:�"O�U��eذ��i��p�6�"Ol�ɣc�&]��bg:{<��A"O8�;�)j�p���6qI�"O�x ��6D���ЯD�5�H�"O 	@��R�Uiژ�``��U)w"O�i/��< �肤>�!��Hq!�D��1� ĩ�e^��	�	��Bf!�*mdD��bQ
|�$]إ���<s!�B�)��S�+�\��5�����!��˻)z(@�%�=���ғA҂�!��O*=��I2/�l��<�Ѐ��H�!�DK1tp�DyÃ�RjM���W7!��� w���B!�6\C��7��}C!򤚵8�a�Ɲ=8�N�K��ݱ.a!�_�m�F�sFM��;��p��Ѓ4�!�DчH��n�dlH=�&ը	!�D�C�*A8s��
��hS�B.�!򤟃-�Zp)%�׬s�Ţ��8�!�G���`�� R���	&�X(5�!��T�h�8�,ǮG*�0▃L=7@a��Ob�5���)��eѥ�.TP��S"OF��G@��
�re!�)N��#�"Or͂EE��+���(�L�X�Z"OJ$ڑC� s`P�4Ɋ�RG"Ot�qf
Ȁ[��)���a�4��"O�1bw�.�`�T�ם`H��p�O���d��|��(����+�&p�I$E!�� \5ކNn��C��80����"O�X�1M� ��ݫv�̈́!��� "O�qd��t ��'SZU��a�"O �s�jG�(�x�/{�䱱R"O  bG������6W���"O���H�JB��&�4A��ٹ�"O�����X;L�*���E���I+�"O��b l�Of�h��&��4�dmS�"O0�tE�"���S7F�D�.
�"OjX�ߕ4�̘�߉cK%u�!��8T,�0!K�l�Z�K���3�!��9X����I'O��Z��J�6U!�D �g��cB,��֮�î	7\$!�$N�n.lxF!J7����A�ζ2��{�D�;���6&�UHPi�2�H�	�!��C�D��0����Ѽ[�J�Y!򄅠�xx0� \�P�J�C�$�!�1��e�p���� "t�6�!��C�*r$]٦!Y!�2`��hSd�!�$#XS������ -���I5-І*!��ߎY�	iC* �x���ۀ%��md!��酣7N�d E+��C�!�D<~0r�;�G�8��� E�j��IU��dAF�?P���(dj(��C�:%������_�1��@%�`O��dF�@%�{�cI,��h�jI�*�!�d��M]|��f�8���4��-Y!��Q���(��G�$�Q�U�R�u !�d�9Tpi3`E�f�x@[���d�!�]p��D��Øe|�xX@I�G�!��4���!@��Cuf=�QeW�k4!�HY����D�]�E[���gR+f3!�X;h��)��U4{?$ `BʼL$!��-�F��1�Qw?Dxq"
�V;!�đ�e��U�a�˨H�䌐p��-RN!��I�	I�8ߌ/:r��"O�&�pB�ɉf��D@���:{�&h��(e2B�	�`׾|��ǚ&.��y2�@nOB�	8`��x��JQ/@��#A^`SRC�I�{^�IД�X�X�`�
���DC�	��J��k �Q��\�"��x�C䉬Hz�)�HXh�}X�/qF�C�$C��(b`��Kܙ\���d"OjA�����!����^�Yg"O(e�D�K8�lA��f���"O�� &�T�~8�E�w�����<�0"O�i*bjN<5��K#"L�����"O<L�&���3�y��k
�K�4D�V"Oʝw���x��`��JO��I1�"OnR%�ݽBI�mҕJ�c�bȲ"O�����s��1k��N�H8[�"O|I(��=�JDZP	�a�|��"O��x�a��Kl@���NB6�}b�"O����K���)��\$����@"O�S蔠i�����j�,Ug�Mk "O& �/d>h� �dטi����&"O���ǻ?��{�	J	�H]&"O�i�aw���0��ɲY����"O"��
�\��U��Q�;�\1:�"On��w�ɉ����逝\Ϊ8�"O�ȪSIn�Ā��蛸Z��t�u"O�X��K�yO�I���C�0�vE�"O�)˕��H�;�3[z xP"OrH�N�5i6j���^s4��"O� ��2�́�N��C􈝾Cy�W"Ov,p&l /WF��H��.`F�Т"O��c���$D�e�7dɐ��mr"O�Ź� �P[r�Z����� ��"O�;
_h�, h�b�8#����"O\P8���*��$�$�j{��Qd"O���t�N��#=	`���"O޸����'�=�'cٮsR��"ORDS��.�H��� {ĦX��"O��'�M�{2��jA���z!"O����фqW����C{�q�3"O�t2E댶O�Ē��ǈ$�x��T"O����ҙ0�xԪ�KG�.��L�`"O�Eh�JʂR3l��F�#��y�"O�Uj�4���g'X&�H��"O|���/t��ĥ�%?�����"O��0է�:h�p�$��!u�͹�"O�ER4 [;	)��Z=}��k�"O-��*����*��	,�>L�g"O�Dx'@��*�J�W<��\�G"O���3�+�쁱@jP#�ntʕ"O� �'�U�y> ��o�8���3"O�(�E���钎<�l�A"O����)�	|����<i��a"O$̰�%\5>d49�L��RI.��"ON5� H�7�$�Q�-p��S�"O�1:�	1DBԝx� �d@#"O�$q��@�j�n\�!ҝ9����P"O��V�M��V�K�">���"OZm�Ö�k'�9#��y�.!#�"O������~�fk���ĉ��"O.u9���cv�]s�j�'�IC�"O�i�J#7qdT��ꀓ�X�p�"O��˅	�F� �ʌ���<��"Of]z�#,����I�y�\�3"O�@K H,<̌L� ���;e"O&y��	�\�b䔧\�,�p"O��C��D<^�ڧ"]�J�l�'�� cҥ �.���%��k�y��'kTd!�g��Il��*�낁i�`	�'�xP6��v?���D��9S�u��'��ͳ� e|��tm�2)+�ui�'@�l@�G^?@�򩰔�B�&�����'Pڬ 4�^m`SPJ�͢�'�2�À��i��B�[��"�'�} %�	@�j�2��I�c�'������r��®Mr���'�b�aG$�U)M�#�AC*@��'#���	�F$���4�QGWqK�'zjD�$ꓸ*��sA��8R�-��'�> �H�),�Xs�39�0�'�� Cqg=~-���"t��
�'�|��� �hd$"����/̱K
�'��R��,Hw.$�%E�<�DY�'����v���(��IR��C�r`p �'���A��%_�LC��[�:BZ�
�'�"��J�|��1����4���B�'J�]2�-�^��b�L�'�����'�h�D�\�*{0���JT�Ȝ

�'!8蘵 M#cĶ=�&�݉P�6�P	�'aHq��?Z�6���E�H��3	�'UKM��
�J����\�8<@q	�'e�SプO{�%I�gE�c�B!H	�'��|���4�La�g��o������� �1"�ļ"^X�i��o�<��"O��j,0؄h"&K��P��"O�㗋�\� �9&�SV�P���"O�y�k�*\|*qG�ΛRײ���"O�$3���l�.�ȵ����0)c&"O��ap.<̀}!R��!S�hi�u"O���h���I%߱'��=s�"O
�:�͂�P4a��K�(}v�V"OB9�M�z�XY���62uPu�""O���L2
�lc�F�bx��ab"O��%��'U*��U��`����"O��&��%=	�HivIֈ����"OĘ���!/�����h�+ИT�b"O�Y����d����Ðj��Pص"O����\=g(��(�(J*%��Bs"O|u��EL�i�*|(b�7KɜH0�"O�e��e�3�����X"w�,9!"O��9����X� ����y҄\+q(d���&í2�Ձ�J*�y�FA�B)f�X�<�.�#d.H��y�ь]pf�j��:�LA"h��y�L � hw��)Lb��1oA��y�Q5w$4U������ҁѮ�#�y�c����'ξ%%�a�D�ȓ(Fe�Q�
Q�A�ӀM �͇�Sf	�u	W�L#4���:K����t�����M��{����b/T�k�>��ȓw��d���vJ�l���)��ȓFc���6AܞDͤ�!	��Uv!�ȓc�p��8l��Q�D���6���ȓ[[�}�&L�Z�؅�TM��V1�ȓ0��Գ��}ӠT9E�I=B��H�������|��M�G�@�#� Y��O+�]`F�1m�&p��+BՅ�ao7m�&��REIY��M��K�,����V��u��� ��ȓ�`��1#ܙT�fm #�Q����ȓg������_İ}�3aњ7�Q�ȓiݢ�.��k0a� �R}ib�
r�<9�� ɞ<��ˀye�h��
r�<	'�@�YYT�ZpI�J\�}��%
n�<�A��GD��`��Ӛqq�JGj�<Ye-�m'�L����8��@��N�<�i� ���)�d����P��M�<����'Q�{1	
�l��0!�
�G�<A0�V�~RU�u���r�\��pK A�<q��.��qUf�$!��u��y�<�& U$qp�TY��tb98өv�<��1�V*$/�^i4�$5ÜC�	�nZ�b�[!<�(,����"�ZC��n�Ĉ���x���Y"�\B�I6^�.��rHsQ�}x+@B䉧S�m+�-� W���[d�	[Q�B��/9�h��X�u���%^�B䉣�Rx�FI�^�^����Y��B�ɍ^y�sc ޖqh��B�V�B�ɐ,�<DP,�(/�MZ���;��B�ɫ�$(q�ɎP��i�kJ_p�B��z!Jսvc�5���J�t^^B�	�q-�ɲĂ�0�r4���ĖM�C�ə<$����u&��Je-�b��C�ɉ3�0�&���Y�fԋ�iШ6�C䉐�>m���O�"�L�RR�*c�BC��%�	�v��s��Sg*s��C�)� �5)�玩 76ܺRۙ�^��%"O�ؐ�C�RP`���Yz��a"O`�cg�#FDd<r�N�m�
��E"O���ƫ!�@ұ��*��)B"OҰ)a�ól_F����%�T�w"Op���H<�Y"s�)\H@���'�ў"~R6kR�lDj���ހf<R� �
�y"�Ż%����AM�F�����ù�y���(�J4�R��7��p�i�yOX�밤x�ɺ8��qp�C�y�fŬ����<U���&� ;C�I/Ih�換�(��\R�	M��&C�	��dz.\5Xª����εh:�B�I�8�4��eC]46��9P�P"�C�	<Iٜ�3���\��6��B��~��H��,��Z��q��/��B䉾r��|x��  vBDh�X�U�|C�	�Z�:Q����(֋�*B�Ɍ�*�80a>M�ZUC(��F,*B�I JƝ�䦒#*�k��OFB�	+$Q�%�L�D]*�Uؖ6�:B�I�:�p�b	�:6�b( `��=4�C�ɨr��x��$��&Ւh3��H m�|C��1C]�X�����D
VCHr-^C�*&',Iɷ�S�{*�t�b��� �&C��=f!.�ذ'�m\m�?,�X���,Q��!*=���x��WH���?	ӓ_(,��J�
�Ny�T#V,I���]t,�S2�̒~����"݅i����Bl��;���x_�͈eeX���;���ԮI�^���j3�'[�v������Jr*݁2�|��t�D���Ab|=�6���L��M��E}@�ȓsf`��gB%`�X�#�JB�ȓ/+Ȉ�点/AhM�3%cx�م�1*"@å�
+f�=�$���&9��0ŀH�T�	! Wh<�2%�4~
��ȓ-�P�kXky���U
G�e9J���`�R<��J��5j(z�!]0i]^��ȓh?�Y���_�LաvBL*gU�ȓK|>�;e%�r�:1z��%y�|��ȓN��@sNӭY��9!�'�+�.y�ȓ��Yq&�z�����d��A��C�����D'^z���DA*��ȓir�����&bxDɈ�`��x�ȓOz�`�
S�{Nd�DO��SBNՆȓ*��|p��ʈ�@��A�C*cb '��E{�Oa�Ɋh)v�ڒ�B�X����'�S��C�I2[l��� ����!DB͊C�	�#
�f�٘=?�h���0�TC�	�"��a�e��D�z��+f�ZB�/=Y6͸g�����Qiܾr�t������������a��z����ȓ�0ɣ!@�=C*6fN8X��f��q ��3YqK���0R�,�ȓ{r4�P�w�0��D��#5$  ��J��xz�+��G9����)���\�l��FI�ea���mH�d��ȓ�&�;�Ao���ÖL����ȓ��@�d�K:p�&)C�H�hX�ȓ? � �QV.�� )ܥj����ȓ=�Fy��E�0uwX�JF���U���Sy̔��(I�R��e���]�Eк��ȓc`l��W�Ft�h�L��S�? �A�NS-D��8c%[/fTY�Q"O��i��Y�^���
h8��a.D��1���^��9��%�?b0��i+D����GV������ەs��s�+D�hyu��$:���/͏Y4�U���*D���g%_/���3rKO�A���4�&D���P+LG,,�RkξRG���so'D���@�U
Bm(�k���޸�P��%D�H�JT)�&�b�R&1_�i�sF"D�8�rd�@��]��I�&Y����2D��QO�E���+�-L�ii������O�=E�$CF�/ېu���H\�d�҇&a�!���+Q�>�I'G�#��x��&�<i�!��(4a���B��@�d5�Q�˶K�!�� _����sx
�@$n�J�!�$�!T�͒G~}�Y�dϝG$!�$ɰ��܂��y���"�g!!���K�:Qʥ�<0R��Ee�0l!�����A�v�W��$	W#�6W�!�Hz�9C�e�M�`q�"��<�!�d�{:`j�]�|Ur���|�!��F6p�XɰdR.B��4���U��'�a|bBV�i�q[0(�J�,roO�y2�	5����DC*V�X �a�-�y�,M�;?�)���R;L)%�dI��yrIB�>>�iR❲2z���Z�yR-�0*\ce�V�F4�+��H3�yr@�(<�D��VG�-~����y�g��g�f�I$,ɺ�h$s�� �y�n�Xo����3iI0,�'�y"Ǟ?��a�K�{)>��d�+�y�&�%NMEzA�V��(�����6�y����!]@5��OƸt�V\�$lS��y��L� U!���q]�C�'�7�y�b��Ay��*��b^Љ�lX��y�YOɨP��)�[:��Z�8�����8�2�PŎ3(5d���O^�{6����"O�t�DK��(n!����n�X��S"O���"�:�\5���Z�uy��'��H:ËB��,�Pu�ُ,���w�9D��Jө�7
�4j��W�X���#:D��8ūA>:R4���)er` �*D�8�l���|I����&gL�b1�3��=�OҠ�E�F���\�NӰ*("@;t"O�L;����r״H��E'$� "O�I��_�0Q���@�'\����!�S��-�8a��$�(C��D2�`Ȝj=ў���"^DUi��\ N�p��d+��T�C�I&ͨM{�`��̑�+�0A��C�	��I���T;Z���fPjC�I�s�~HCCʂC+b䛖�
E�bC�	�v �i���@�8�=<�$C�l���	U)ΛT�X�႒�U��<���2,3��ʃ-�FxqćP�C��B䉎��Ig��N���Q)M�B�$C�	;{ft���$vR����V��B��<y��ys_?$nl�hD�B�	���� :b�f�k *DC�[�eS��T�x�(��T��C�XC��Hq�I�"�^�o�f��VŞ0\FC�.m�$��@�B��5a�� �~0˓�hOQ>�x�B@E+�!s�B�<���0�b.D�IeF��@KE���&�ٵ,D�( 4�K
d ^���D ��8@�&D�� L+��Ԏ.��8� οL鎍�s"O�	��<)�j�� �s5*1�"O�[�n�(Je��S�I��J7f=��"O0�S!��)pHMiG��/
"�jdX���'-���>���@�u���T�@�����WME�<y�m�$46�P�����qb�Uj�<�`�C�;pJ�<����H
o�<q�H�,�ڠJ�"eR���Xi�<��^F��`�����G(-+��N�<�%
�(`+TԹ����X��8�ӨNH�<�E�E����ݠp�<�r� [ȟ���8���f`K�i�>Q 
��N����ȓF��e3Dh�(6���V���*�ʤ$��F{���$˨m�z�� �I���z҅���yb��xn�+�`��k�t�p ٺ�y�!�,V���'��/1�M#���*�yR�Z�UW��1"�V�v�2�)��լ��D$�S�OҪ=Bq�ôRm��ç�v�U+��?��O�TH L� c��|`ՎZ�$���w"Oz�sr��$3)F�#�	�BtS��'r�H�U�ʌWb1����E�\���"%D�xS4��4iX� �%o��'I$Գ�i#D��H��Sk�b#�ɟs�\p��&D���(�� yBFĬC)��c�f/D�x�g��NĨ�Y`n��Z���۷@+D���s(�!�X�3�DbH���'%+D���SB��]%�E�7��>q�<���*D��r�Kn�\8��*�r?8#� )D���A�E�Xp��X�e5/]RA�Q-(D��WLӾXH5h�mQ9?���w�#D��;�I~m���@!��p(p��L �OD�;���IԝK�<qs�A?B���'��E{��D��3g��e��ȯo�0��0i�y��P~h�a��ƟR��9	 n��y��\�*�� �ǅ��G���hG�Q��?I�'*8��bm�	:���xBȝ�!ӦIS�'�z !��萡��;	g$��'���1�@��7!����ͯ|O�С�b�)���A4X�bR�̸k+:`��f�$�y2HA�q�RA��pX�Bw%�=�ybO��*�!��b[�(S�E�hO4���SM:q`� �
d<�Ԫ{�!��Q�^�fI�cEMeP�r`ˋ�!���3N��xG$���&�j��D/~�!��y2�0�h�J�`	!')D&e��y��D̀N�����n�+7�BU��oP�y�|㟨�?��y�P7Hyx�-�#D���.@(�y".6)�nh�Ҭ�"R9J$x�$ߗ�y"�Tz8А����ְ�@D��y�@�1~^ʡ���!#�x����y�b&xl�Tҕb`28�gψ��y���J�Ȑ	�E���P��@��y��1-A<ݑ̟�=VD����B���>a�Ox��iR�>�]��DW)`Z��b��&�S�)��h{��C�ò8WvP��Eԩo�!��X_Y l�"F���D���c��N�!��0	u8<Ä��`$�qԌ�!Jb!�ۥKʭB���:�T�k��m�!�����#��0�P�2a \H!�>2J����F���*3�btB�?6~��n͸B�6!�ÄN>>��$9扶S���i��[=H4qC1ͧ'i6B�ɮDnT�0 �	-[f�iv�&HMRB�I�w��qJM�Q�� �o�%(C�)� ��d�����F�z�4;�"O
m�[!l<�3���k�t��"O
��%3�Y��c�x���u"O<�{�D�7Y� �٤L�q���A�"O2%!EB?V(�c�j��f�(�"O����D	$�	A�	�<e�&X�6"O���
ÌQp0hΧT�q�"O.�8��W�.!Ԡ����C�f �"O<t2�Ǔ4[D����� GæAڠ"O6H�u�F�1�x��� O#&QhZp"O�THĄ���^���F	 ?��d"ONJ�gD�%�|���ߟZ`��b"Ob�a! ��|�Z�#ā��V�>t��"O���΅9"��K��U�#�*�R�"Op�qB��	e�̹�Dg� @��ܫ�"O6�QTl�0Z�$*��0d�`��"OȘ �*r'��R
4y����"O@�z�m�&M��"�C�lYbԫ�"Ozi�C�F!l��<q�ˍ to�Q"O"��AO�O8���H��tO�!Ö"O�X��$ٗX�f,	��T�6�-i�"O������N�����
x@�K&"O8\��o\3M��h xD���'�ў"~�'��9�H�����Ey�'_�y"c�h&ܼ��C��` §f��y���o#��B3N�-P�4t����yD	<.�R��ڬMmn(�U�϶��<	N>���	eG8�QXȴ�w�O�Pi@��8D�����3oZ !��� �ř2�,D�`��g�#Iv�Y3H�30��	��(D��@G'4 �"yIq
71\�p*�#D��*�/-g~��u��<i���T�+D���@��yઔ���ʡ��<����Od�#�S�Ojh���},e�v"�9������hO?��ّtT�ib.	</���hC�G�<�c��\)��UlķD��e�Q��h�<Y��
l� � �	urr�+���c�<��� kq(]kSK��T�Z�KV��[�<��[&n�p�CCM�	%�����T�<�V�Sy��� 1g���r��S�<��U�8�hE�d��,@G�U�<q7/�H�����Ñ�P�8ŋ��N�<��+�ed�QH�b�47Ͳ�c�F�F�<�����|�ڀ��q���@L@�<�J��2I'���^��m�P�Yb�<�#��Fd񬕫93���e�Z�<1�*Uh�n)��&��bhXa�<2�������H�a&�����`�<9`O� $t���	�J����XG�<yd�;p�"�	��H�
��u��D�<A4f�zNd��� _֌����[�<6�G f���p��N��A�n�Z�<1��V���h����\�2r�Yh<i�#��>�8��Q�0�����?��'�"�s�¨B8�W-B�"�`U
*O�=E��MA�nxB��rb���q�$�y��e^,���f��yvN¸�y"J�?�����&I�~m�������0>���J6}C'F2I�.�9��Z�<����vb�k�ݗ u�<��\Z�<9��įL]J�B�(�a�I�RAHV�<qu��(�틵%��+M���
�Q�<�E�B�t��hX���U&|]���T�<��OY"8�6#k�?~
�a�ƧM�<� a����*Q�ı��]
2�٘��|��''��(?i��O�AI��W5y��T��Qs�<�P퓡��p��,�-o͊ų%�n�<�w-A|_$ �$� �X��ViFl��b���O��Qs$�
a�N5Y�jB��	�'�2y����<��8���\��i��'ݔ5�UO�NK�'��N6��Q�'�
��ψ�,�T� �X�V���'f��A�]�Q'h��7,�*?ה��	�'� �1�[��P��38�	�'�fQ�F�ŴbgJx�& A7-��ŉ	�'�d�����67L��6O' �ꡒ�'<��I���"b���#�dK�C�-��'p�S���
/��Q9*�|A�'�����_%8=L92�C���8��'!թ��ȱa�$-��g�+�h��'Ԟ�	�F4 _"�qw�)@zl���'Q
q*[���x�3��I���'����A^7)���CN�/C��+O����qL��	BET�et�da��@&@�!�dЦ
bTj��--n�����"�!�K�f��������9b]��$��O��P��U~"�^�&
$i`� _qX�cJ��yB�Q>����e��H"�dR��R�y"�
AP�X��ϗH��u��AD;�yB�4Y�#�_>d� � ጰ�?a	�'�X��k '@(\��Է0\n���'�" B�nF8KE��c��(Q�T�'{Bd�cb�4�� i�+8:�l`��<ayX�pc��iK�oK>.!�D�v�~a�r'�0$��	��NY*�!�݉	��
e�1T��1��m��J!�$Y>u�G��V�:�X,W��	D���!�_�g�}"�`$�ظ��$D��
�≳��ɗ��w�����#D�� �K:S�}�#�b�XL؇7<O�"�	�D����C!��.�� �f��z�dC�3T����D�1��h��� dVC�	-1!A�����v�!�	;��=)�'H�]��FK��D�� B=>�|��T���s�O�&~Vl���T�p��[�X!���Y,B\��s����E���`���s�gI��񣃢jc>��ʓ�&���Nͨ.IȒ�HvL�B����A'�&Z�V@{U�D�\�dC�I�2�L00�7'N�{��A�d�|�?QJ>�ȟ�1�

'A!2<��������pE"OF��%���3���%`�+6��J'"On�(�����%�@�#H��Z�"OZ��BhUrU�@��m�m�@�|bY�D��'>X��w)E���5'��'ٴ{�'uZ�I�J,jzҏ��M��P�'f}
"d��_^ȱ�f��J�����'���0q#[�#X�i 2�š{��*�'*�mx��7$v �9f���}��	�'�� v�Z�2��T2��Ŭry�p�
�'L&��� X�N��5B���t�.O���ص�p��o�f���oK�"�!���g"P��d�N�c|9顎�D�!���fT��"4ty QY���!�ʡF% ���A^2xc��H�O٘X!�V9���r'	C'�n�j1�ޱZH!�2J �3��Љ�:�"牘N>!�Ē���%nM�[�
��tHm�!�� r�)��	�6>��PfI\�O��5P'"OaC�gR�s��d�1N"�ZȠ6"O����d�ƌ�2�B<+`��"O^X�QJ�Zf���DO�8/n��D"O�XZ��L:vy  "��1���I�"O�0��S2<�(�`�	�R��"OD�k�n®9{��qK�'�"�p�"O\�!c`U'�|rP���t��q"O�ؚ Ç#a�6��,�Y78�q"O�ܩW!T(	��٢wJ3Q���"O���w�|@��`Ʈވ8�4��"O��5b�N�yJ���v��ub�"O`�AO�7!5bE �i�)5F��"O,�j F�T<z��2H�2f޼K�"OFMYkE>N�C�-c���f"O|��dUҌ�eO}CR�p�"O��X�-�0+�!ْD��R$z���"O��pC8}H>0cT���"Oʑ��m��S)�Eb�(9�m�"O�`�4��8�6��â��3�$�f"O8�Xb���S561�� ۟<�F-!�"O&]y
ɝBהQ�w�]N��
�"O�0�S(�gWPh�;-��"O����;ZiA��_���"O��B�C0�8ڇI\�S�9�"O���ef���XRr�/�v8c"O����[� �RD��&Q�A��"Or��E-ݗ5z*�r�M�52���"O$���R�<t<��,�:2V�"OJԳf$t���� ��:�ma�"O,��@H�2;x\U��V"��"O�9i0�
Y�5`3K�*�����"O�騦#�#�4�ԯ��8�&`��"O�\�ͷX4���櫐K��,2"O���Q�"�X���}����"Oށx$�VC������b���s"O�u)��bt�G$�={b M��"Oƈ����$`(����D�.��"O����He��q�5f?pmJ�"O�!Oڈ<�*�y�_� ��"O\-�D��"�jAl���]:q"O,��!l�9��l�4,��n����"OTU���m�����T,l�-�$"D���2�^:�Lq�T���!D��!2H�(48���0JU/QR4�S�	?D��!��_�,�l���ԯ6�f�B�E;D��6��>Kƭ�&�ӫ �$2��8D��[!�Î"�^�Õ��N�Ц�7D���t��|p�-��^[Fr��4D�x�6��3�:T��hƛiQ�-k�B%D���ͥ K�b�E���?!�dX+ށz�`JV�B`�퉺^��'$�OV">���͜j.V�c��U;&�u��ǆx�<9��H�\��─�4�T���*�t�<A�gD�`�*��y`E�2$��ȓ l�Ӏ�?�dH9�"�'j�t-�ȓ6ݎ��� �=*��a�A�T�%��7q���"��I�A�Gˉ�7�����D	(�̞ ���bsn(��'�,��I��8á�?�F��TcZ�xB䉉m�|�q/@&�p81��?F	B�	 ����SW�S�v�!Ǆ.:ǶC�I�G4���ovh@��D�#q<C�	9u�$�g�*��q���-T�bB�)� Q*���BY`�\�)rpc%"Ot�R��8�l=����n@��W"Ol�rK!h�UA�8o5����"O�@��3d�~A�a��-W:tk#"O��ӆI�O��ᩓ�B�6��s�"O\��`F�����E�i9� R#"O��$�,�hH�W�ŻG�Qj�"O޴鐨B.l�����X�j%��"O��2��%���ɳU������$"LO�����N?<�zt�. =���f�'�!�d�:�&��:_�ތ#@��K\!�$�!���;f̂�H�� �6�!�d�3<J��d������ڝp��yB�I�xlj������;UiH�c2�C��d_x��c�E�Z\���b�.7F:B�I/P����"Nɜ_dsdJ�.�<˓�0?�Ƈ�/1'�����Ik+|�8%H]�<	��M^� �H%_T�tȂ~�<�nG�[<ِp��.}ڔS��c�<Q�'y5XՃV%����́�[�<b�Ѓ'��a
'�L�*��,A��B�I�(���jv���'�`svf���B�	�c�*�+�'T<Q:Pr�ᇋPF�B�I=y�����^�F�ǿ��C�$V8$ �A��=;�F����0�ZC䉱<���1�Ύ*`��h�ӆG�C��09��țI�^���h�	B�N�B�I8k�x���N9��X�C��|{B��'������*�	C6*���B�	�$�n�����(RRx���_5F�C�I�	�����ay�:��^���C��3������p�4��6\+E+nB��kP�A[��ި6!`���e�(K,B�	�l!l`�Z�p�D���&�*~�C�I#V�.�rm�/ <#2.��"DB�	e��(�p�
�	�,��iB�I���z��Ն{q�񒕪��%g�C�	 w�%��$W'hG�	����>��T��K�d���W�2�b�D�[��C�ɻs�*��g#��45�0��Y����ȓ�n�[��=�np��mK�k^f�� ����7�Og7xT�I��?�����{�
9�É�O'ڝ(��/��l�ȓIfT�s-Т���3��2B�¨�?����~���[!Z���e�VÁfC~��T�')1O>!�h�1G��qRK��Dy"O�`s���#%���ӵ*��;x���"O���f�*7��؆�X/O���҇"Ox�R�̓&���&�EXL�1"Ol1��� B��Xjb�*T��"OJA��%������-mp�"O`,#�K��X�D����Q�t��q�Q[��F{���F;pti� �V�l�Z���=�!�dV�J$to� ��Z���*qh2C�I��!�SE[0J���G�ʛRQ�lD{J?�@Pß?JUVaRpiP�Y�>�e$D�DS��Q1;h���+��C����&D��z�FϟQ�����=u�J8i��$����D5擞V�*����^��A3`(��w�(B�	_�dj�THl�Iwa�|Z"B�	��t�"���|���^�, B�>/Ubq�GL�$�+#w�Lj�'�T �v,�7\P���n��(�'�l�G�ٜw@A#ץ��`x�x���� 
0�F��H���ӌa�Pq��"OL�2�$�1;�@�9A,�+x����"Ord�3iA�R�^]aWeבY�:(j"OdI�t�N�7�Ƭ���Ag"O�M�VeCr4�Qd�s�ɦ"OH-����P $30c��pK����"O��X�X>�ج�!+N=�H�"O�]xB�2w���QT�<m(�Q���	�@pp���5������L�ʓ�0?a�%�201"!�7��BkנeX�Y�ȓL���р(9�:42碔�'RȆ�����bH˚=�2-�#o4(�BĆȓM�������.���x��B�,F��ȓF6*AcǶC��K�Ej�JĆȓD�� � F̾�x��v-O�}az��ȓ;���s`��8�����~H��ȓf�k�a�0u�8<���Â_�2�ȓ2<А��E;Y���BS:H���ȓ`	��Q ��^ۖH{p��?U�\��TX��Ko�Z�"�nД��1?���#@�G����]�&�ȆȓqSvћP�^$0S�t�DJf���w����b�/k\��M:,�����]"�ɸ�F>c^�����8r��8��]���[�� 7�z�Ս�5~�x�ȓ޺=��>��9�C-�&��=���S��D�/@�,�U�L>"V܆ȓY2t�i��E�j��� aʠx*��D{�O VU�E��bl�#)C�1�H<��x���q�������4ryw�U��y"�w�B��g�@�<e����y�Ɓl j�g��!*v�4�y�b�h���ޕ�	��	�yb�#�����O!� X�M�?�y�L	����ჷ3��$jU��y���+c,n퀅����"��yR� ��I�϶
���h#����y�)��"70�qh�v�"����y(�h�l̩'�
l��q6놥�yb/�:I��)P�[�W+���2��y2��N�@t����I�mۢ�;�ybE�����,�>ٜ��q�	�y��Μ%�4=���/[R s�,���'?ў�O<�� D��hI����b���'���`d%�n�B��J��T+v��'���9F�@/Y:D��q�W����'A���gB�z�pdמQ��u��'2�9�G)[>"lvAq@lF�~xh呎B�)���W3����Ԍ��S4����
΅�y��I�|��S'���&!��yr�B?1�N��3�Ĥ+!\���n���yRG	F-{��!9F@Ռ˖�y��*K�]�@M�;�0y$`Ý�yr��HF��j�r�̱pE@�&�yC�<6�z�2���e�T�Q�^��hOT�����m���`%��,Ǆ�(��\!!�Ĉ��i�Q`�J��Q�$�,G!���PFмp�[�~ Z)I!�Duk�(�a!�
n�|�PJ�7@!��)L�\�{��K���`&*�0V8!�D]$3�J(�Ԇ�	��x� ���GI!�I
~��- tm�+�$|j�[�MG!�ė$ �t	�pɅ6Z�(�J*7ў���ӆEx��!��n�x��1��(�.B�)� X)�������G���I�u+a"OTH�rN@�S�����H5�y��"OTt�"� *�t�JA(V0w�@�"O� ���m9���!\�L�V�9�"OF�G�/M����u'զDn����"O�{u��e
���aނ5i��cd�|r�'q><+�8	��Z2jӀ{L���"O&M�R�ʨo�x�S�i��?䤹�4"O"����ԓ!���:R+[)�v�Q�"Op� �5_Ϯ`XR	ݔ�Xlj'"O������
K������ K��R"O��k�aX$7��3�,��B�6l鷛|r�)�ӱ14�Ԋ�lX5	��x��Cd>�O,�=�}�s��lٺ��@ȕ���7Ŏ �y-��p=
k\�#�6@F�$�y�"�fBd��T�SF���č��y���Hl������L8��A� ��yR`X-a^��A�>Ț�à���y���"9�Xx2f_�5���  �C��y.�cO�AA�ٍ',ڭ�W�_��y�<<����2KKdL{����y&T�m� �"� �F��1e��ybK��m�V�����h>V�;3�J��y�́�m=̐a���,�R,��獸�yB�1PnQ�����\�b�̓�yr+ȼ<�R,)�A���bh�� ��y�C�[!���&��/F{<�y�gK��yR��Hq�0z0H�r����c�N��ybM98�r��]�i�Ā+sG��yr��/���Е��a@@Q T���y�.�,.3�E�󠊢"�|i�k���yr���r,�0���\�s��I#G�y���7�J@H��]�iAG��y�d�9^��uU�ɧE�(,��B��yZz@��@!�IF���AJL�a.�-��x袀Y�.ɥ=��-)B�
���ȓr�z�`��M�
��ܐ�n	H	�T���2�-�	Z��q(q�N.,Iz��ȓc��H!h��>bꌩ���m����ȓ�6� �O�:ޅɥlA�2@�݇�B�B��Qc*�|��鞛d��Շȓ��i:��\���!f��Jx*U��i	FΎV�H�iw0��x�ȓWِQ(%�U�K�P��I� {���ȓ)w��$���JD!�'$�>���ȓRX�`PS��3g��M۠�^�'�$�� K�%l@=.j@	c��R�V��ȓQ�Ȱ��35;�{R,�<T����a��)�6����}����$B�]�ȓ#:b�#�`���閆5D���C&�|����T�fe�N�
��ȓ
Bt�ht͇(I�4��"��j���ȓuƉ�)~�h�����%�ȓ1�� ���ca�M:� �$��8��c]�i�?�=���S�>;�=�ȓ.~ YvY�,�1��^� ݜɆ��m��nG@8�!*��+��l�ȓ�"J��)�|@a��h�` ��:,�x
��!e�:M�6����}�ȓ	���R�aH"Ь��Ӄ�_[ֵ��(E�=R�J)���g�
p��q�ȓ�T=��N�,�dUA���w�=�ȓ+����4ZB�pf�_���h�����{2�U8��(o+S�I��S�? T��фئwnz`��^:�Lp��"O�̨�����|po��r�X9�"O�Z$(�)!/�T薧ܶNk�xb�"OF�v��@�T�R� R>#_��&"O$\
S�K5Mr��&o�>j��+"O��bs䛑��u��u����"O�)�&+;���T��:mwz��E"O8��ӨV'�ݺbl��jV"Ox�!�P:@="6-ڷ*q�asD"O�̓���\�$-cEeŰo����"O��r ��-������N
��b�"O�̢�-JX̎Ȼ��g����"O�-�5�5V� P��te�X�"OJPB�DѦO������
I�0��"O��ipGG�KϺ)�˻9d��"O ��q��>?K��"ĕ*�BT3�"O�y"�������c�,�X$Z�"O�!�I��i�^I@GCT]gYSE"ONlJ5�D4�X1��ōQM�"OD�I ��`����������"O^�����
��UQ�`� �r���"Ot@"V�8N�((tA��$8Ay3"O�칖���Z��t��o�U����e"O`��m�D}����#T*�P2"O���	Amz�]��ن]FL�[�"O�=A�H�?���k��D3��0"O���`�N��@5��'<*��8�"O��Ha��mQ(������~��"O�m��聮Wq���&��a8���B"OT�+��(EP�I��(�#)t� a"O���V哅P?!�F�
*6��"O��'�<;��JE���d"O����:tsʥ���9� ��"O�Hb���3L� �Շ�>\8��"O��ʒ���T+^���gۢY^\Ir�"O���',;A�lq���4 "��u"O��o��E��U�a�T�,>����"O���к01`\:��/W=��"O��0���2?�D�@.X�<n�!�"O��+�⅛�*`C��U�F���"O�t�� ŋMǞXP3H�0bڔ�pG"O����	zH�Q�E���C"O�}j��ˣ7Ţ���fz����"OS��W�U��p�G�NR�\p��"OT�c�
��+&菨N�jd��"ON�*��ܥn�>�Eg�%o��ĺ�"Od�h��&,���P�Z�!�:l�*O�9�'"Z�`=�&�7_|)R	�'�r�+Ǧ	%��!QRk�,3� ��'\�\�BK%����1Ύ2C��h�'sh�Q�
K�s��\AQ!
�# �
�')�x����9n�pc�Ҋf�T�q
�'����.(G�@�D<$QS
�'3f�r!�ڍ%K��at�С���'�dhІ�2��LQ�ߛt|$z�'�R�K� =>�a�딸U���$�`A��+�伣3�M�x=&X��pK��K���D���E%ϰ��%�ȓY6&�+���y�8yċ	V�x������b�b�Ȩ��������4aht� ,^h�sRDO;x�>���s!�p$]�n����Ě�:%�}�ȓ"+�"�}��]�Ǆ0� �ȓt�$�y�f�8�H꤬υ-�Rh��S�? 0���_�7�R��Ç�AD,�@"O�;4ɂ�Q2�@
�B�Y
^8��"O֜R�D�E"z4��ɕ[�d)�"O(�X�c���̅�A���"O���"��Ehx���o�o�̡�"O��DN�*�V2�N8!��R"O��[cG�M��S&N
>DB�[""O8�b�)֭i5 �"�[���H+�"O�q`�C٦-C���p.�.H`^�Ѕ"O��#��F6�I@1� �{���c"O6)��	8��Z��Y�
�����"O�5Q�E�VB�3��آ3���"O��@��C�.�4 $�/V�B@ �"O\�+BHʿ1ؠ�f��0�Z�C"O@�KW�ҝU\P
@%���5�"O�= ��Y"CO�@2gd��a�N͹w"O!P1cڟ#�|\1�J�R@���g"O�cp�^�"+[yrjù6���ڐ"O��z�E��V?���ֿn{��2"O`]��
Iu�ip��[b�5�"O���kd5h�me�n�A�"O��[w��A�8;p�̽��8��"O<��T����(����e��[�"OJ���";�X��W	Ĵ;!��"O*|��(74J�d�Y�;'Nɲ�"Ot���G�T5��D�!Y��0a"OL�ɰ�G�o����_�v���b�"Oh|q���Y>
=y���9ڄ�Q"On��1m�
V�)a�A$q�j!q "OH�[g��m�h��5,�)@�4Q�""O�)��-��l!&��q�"Oh�1$.��s��9cE1I�fdh�"O������D�!Q��1Kv"O(죁㔺yA��!"×�/��,j�"O`�#ND�9�:1��ͫl����S"O��c���Z$ހj���*,.��"OK��Vy���EF!0�`�7�;�y"(G'a���C��J�?N)�J���y�,ܠaJh:�M�"r�ԽK	1�yb!��6)P�L1\��}iw�͕�y��զ-�,���+�`(��S��y��ւ
������**�Գ1�Է�y+��\����)�)��Q:��y�I[��p%!eP(��*�E���y��cM�y��O�j��/]�y��R:`����h� ������.�y�L�k�iZ4hCn2��@�%G��yR�={�e{��W�s=L�PhE��y��\�%C��b	0m�F�[��L��y�,S
mD�{孛=g+>���߲�y2 �SD��
�k&"=����yBc�2ܔ��0�*_y"L�@�M �y��
P3�HI�L�\v��aP�ͧ�y�⊔d��R���[K�0XS����yR(�;�t�8á]�K�	R��	�y���Y$�@��9@ ԱHb���y�Nq�9UN�8٪�����yB#M�9)��$��:��)�A�?�yr�`J����!6T���=�yb��5J��]��M~k*�����9�y�#� n�d�S ��x� H�rJZ��yB���`˂+�%n?�0�#�7�y2Ɏ+1|ʈ9�/Y]�jAYP肴�y��&R�N�����h� �)�f��y
� t;@(��y���y�K�#˸��P"Op�p�B��z,����E�`P�Us�"Ovu�Ql�>(\�	�eO�b%*�r"O$�e]4'w
 ;%l�1���"Oty*�'ޱ%5�q���єH%\���"O��ذ��� }�rL�%H�!"O�є&ʽj���	���,W�jr5"O0,�CN$\�t h�@�J��S"O�հ�O�i'��DϞ�edi1tP����� �` 3,Ҋz-��#ǝ3/�����2?��c�V8S�;R���(�v�<A�!TGE��f(;A���0B�Z�< ڸCz���;�Io	^�<�ZU��t��DX�e��Y1�Hi�'�ў�>���鞗x��y���Ƀ�"�(�*D��#�$�lH�U���<�p*��'D��X)�:oN�ab�)����	%D�D�$(�.���6���ыdk0D�XB\Pn�[���x~���Ǫ/|O�b�l����B���r��[�eZ��s�,��hO�6]�:��`�ă!g�U��nU���@G{J?mAt$�$b�b��=p�Dy#�ΖxG�<E���PT�R5�׬%��$�R�نx#���?�ӓy�F�10*��vx8�N�_�쑅�N
\QtbO'X�I��W$u}fh�
���'�]�d�G���)�4j�i/xI���hO*%k�� ؎����0�x!���D=�S� ?u�d��L�%9 ��07D��C��#GP�q��@{��_BP���Ix8�K�j^$6hF�� B~�`�d,��p<���7��A"G��s�Π2�N�j8��O��z�M֯U�`���ڦI�@Qa�E2��hO�S'O"Qq���0g4���"� V��">	U
c�,F��HT����T��GӖ��a½�y�#�U���2(K)*���P�K��y�
�(�a�#f��n�F-���0D�"F_4��Y���ƽc&,��*0$��ӷ@��39XYB�FCb�Y4�� �yҋL��r���nl��������<���d��|�%��"mf�9�mZSNaB�O�L��KڈYN�%�a�L<��L�5"O��P�)O���@#��/�L��u�'��OL���@F�)�Sޖaht]�؄��H8��	�(��)�'�b�B�Ʌ?|P-�ק��A��ͪӮT�G��C�ɉJ�� +�o�4+��AD�z�֝�����O<�(��6dS��Y�&l�ɣ"O��Y�n��nF=�F��::x�q4�O��'��<�|%�ޫX����C*�<��tF�j�<YTʕ 7�Y�"l�6%���	�^�6	в�=�)��<iF;B{^���E�0<^�b�Fc�<�	9
���$��%P/(9פ#��x�`(S^��A7$@��J���=i3Ȁ0R���'�`Qa0,P�y�hhȆ���X��K��;�S�4��)�~���W	l|�)v�׵�yB*�\�)8���%X��k7�y���~�V�&酠

,��e�	�`����oܓ��O>!i��N�Tlp�Ӂ��o�Eze"O.l��רB�(e�GKR�S����Ot���r\�R oD�|��p∑�'�Q��D{*���wR)!t�K`j�s�8�{�"O�}P`+��ADOe �4��i�����2
ڜ!P, >%�`QT���b}a{���`��7�TK�H#a/��h��)�O� q���6��̄ᘍ�F%6}��'�8���#v���5"5< ��P	�'�0��%�ϻ
Q�5
֤�67�h8Ȉ�d.,O�р�J) ����(�`�
�"O�򒂝�T�^h�ɏ�0�~�I3�$-LO���%�΢WQ��ptB��H���BOP<�K�(bC��0Dc�;r�Ɇf&D��
^
��ؑ�Y$z
�Q��%D����H��-�l��-��}��e��&&�O@�oO��A6
��{��C�M�;�R|��hO?��稂�k����s2V��N#D��qf'�5,�0+�@I�rD� D���9-hp���j�Bs���PC �O4�z�X�k��5^~ex��\�5c6��"Ox4��7O9`�� ��-AD4c"O��0f	��EI�ٻy,��R�"OD鳕kB�E/Z5���E5֥�`�'�Q��R`�eobuxsM�{7�a��)����}Bv
K�	x
|j��N��C��N�<i�-ޥ �bl �A����3���K~���:�'{�� ��R!X�hA��B3*NB�	�)YB��TO�A
T��]�:�B�I�v�L0��:��չ�޹SZ�C�	��8 �Dӱeg���E�fB��N���*�.꤅���<F"B�ɼ)Ƥe�ƫ�rX~���\{�C�ɐUrN}��\�B�
�s ��T�C�7l-������m�1B��&@�:C䉤���a�4)�yp�-A�%�#<!���?偗�ͷT>a"���o PЪ��1D�T0"�/AR��!zG��F�P�HO?�u3���G�5A���8�J���B�ɽqn|��C�[�������	'��?�tk^&Ry�3��Ԃ26����,W�<I�F�v�^�+��b���Cn�DBў"~��-Vt�9T`F5`�����[$d�|�O8��d�r2H���J�q�<��#F��D"�O~��"	Y���c�A2+��-���d����=q0�x2�S���s��_��}Ad�����O������B�%�E)���F-͝4��(D{ʟ�r����-x4�"x�&\	���|F{��	Թ52��cD���f�6hY"���Dnў0��)`88��#�m�JQ:��;Z"<��32<�2g$�;M��q� �K؍�ȓuu2$pt W-�v	�͝�%UX�C���s�𫳣y'�-��;a$L�g`<LO"⟌��MD�i*x�zMU���e۲�z��̓��>��	T
n��:�m�'֘�q z��q���'b���;J���UF	"Ǩ�"��_�7�2X��� �1�"G�4	 ,���U.:?j#<	�'Eў�]�s48ۄOS�Y BhZ�e��pLC�I�Ѫ���*:����b[w8C��t|FI��%�3��݀��^�_8C��<7��	�ɇ	���S�N%�C�	8� Xr�2��J%j H�C��2��t6�I�T�	�uh���'�`�0B�w �E ��L6"d�Ǔ"�H#<�`��^��ܩ�iK�U��]Q�j�V�<!����=�u���ț���z~rOS~���l�5O,v{,A��C��:���"O"���\P�QlU;'ڢ�{0"O.<3�8 8��R�*F.GsFP�"O��0�^4qX��7�A�t�ze�"O��+4�
l��� �<q��9f"O� .��&�e�ȈU7����"O4��&cɛI����9S���cu"O:�:�W:H�N���V�o�@�"O����%�H����*5��S�"O��#�Q�8h�������`E�`�3"O�]R���x�����!�n=�Y�"O���1"B�2��@�"pZPQ�"O�10*�$�C��[,��7"O���Aq4�Lj'�8kD���"O �Q2��<#9�`;����>\���"Ot
�Q<L�tmqM^1����"O�<ۡi6j{\U T�EJ�j�t"O���(	-���N�/:E�a�"O��8��H�K��MR�@��.4}P�"O"H�m��zX��4o_����"O�A$��;p	$��5.ƐB
�A��"O�I�����2 �VG�/�2��%"O�1�V�_$%��T���M. �ԡyU"O�\����4���9`��&v�,رC"O����:�iR�ȗp$U�W"Oz :���:�=cņ�Kx���"O�1gj�
]ְ�E�� b<�"7"OTْ6k!M���b@&ݓ%JV9�D"O�5�',Y�Taz�yd��8&�i!"O�8+�.M�Oκ����^`���)r"O�Дe̓:l�z�"�<w)��I%"O.��Ǩp�D`d 
�BuĄ�0"O"H+߰��Q�<��9�""O,l��_	7�N�z'��8&=RT"Ox����I�F���cҲ1�� p"Of������!���JRLCrѾ���"O��+�Ń��Rh�cʇ!N�"�!"O
���U���S��F`!ۥ"O�5"�A��>��9��B�59Tx:"O�����DC���k�  9�0e"OR��֯#�T�"CR���P�"OĠ��X/f���^�
E���y��p����nH@%ɂT�p�'Nqk3+�4z^F�%�E�Y�R�'X��vD�*��#u�܀���;	�'���bhG�5���d��sjH���'�*�C64dP�eg&kR����'�rѳ�-�-8^��5��1o����'�VlX��רqt(ܙD�E30&���'8*ti�"Ļ4^n�A�T<)�����'�i�uȕ�0z`�� �Э ��up�'�"��!C�+]E�H@ť��1�(da
�'������Кb�����]�"�~��	�'��X���@������Ɗm��	�'V���VmZ#Z��"�[[���'�V����k��B �0��x�$+D�ȗi��}8��U��6u8!{d*D����*�"���N%y��:DM*D��`�#S���ۇm#+1f&D��ٰ*�vb0��J�1G�5�b�;D��H�]�����F�ظ�Rh6D�S�dK�0bf�xfCG&c�����6D����IU @�Fhр�SZ�9Rs)5D���΀�.��P���XŒ����0D�pc�͛*i��)F#dz��1D��q̏	Ee 9sn±v�(�@�i3D�X�3	]��D[���,��%�� 0D���*m�� #%��G@���2�*D�@9V%�c�Ke��Y|��ɢ�&D�� ,y˖�ǾMLę;gDZ�.���
w"O�U�� L�A�B[��_-<����"O���ŧ!k�5ҕ�Z%TN�P"O�����L7=�|P��o�$=��F"O%(7��=t~U1�/��~�(4"O�D�bD�8�YK�&E��
"O��Ѩ�P>�b+�t��x�"O�a0�15l��S��]��:�B?D��ID��@�r����66\��PҮ=D��"�L�n�4���S[����;D�����U&<�#�#_���E7D���0,�"-�@p��oQ�+r¹��2D����*� Φ��Ϡ[<���P#3D��C��V��݊�#��*`�*B�0D�����B~U�f��HC(�u�/D���%*M(,J ��Oʥv:��t*O��H�]|0|��$�ysjy�"O8�����Y�L�@��e��Ui�"O�!���b�PVY�
l|�/�b�<	�K'v�<��g�[e�$[e�]�<�weǹ.���f��R�|�B��]�<!���1y`9�HR	�:z���W�<	��|�l���� $���G!3T���ce�;�.6*�"�$e��R!�$m��mQwA��H�,t�*��gA!���\<UQ0MQ[ܘ0 qOC�3D!�Dޑw�X�`�
X���-%v&!�d4KŊH��ܦ#�Y��p�|r�O?cd�UH�i���	/pm���;�&|�'�
U1 �B�}�m��M�y4L�*���^`�2��(�b4Hq��O2�e�V ��3E0�IB"O��h��L���j&H�122p�so��$l�D_�g��}��~� ��}�sVf7ø$�T�C��y����Ա�+K��!��A��?Y�����̨��3�0=i���54>����ʹ BǄo�����$xT�:�,5��0���8*�XM� ��\�u�ȓd�2�J��L� +�+C,ףz!��?i�D�wƀY�5�͘��O�6�Js�Ъ�x�PΎ!�N�A�]�5E���
�R��bP�U��x���Eʂ���o�|,U
���Ky�:��8��U�/ܒOp���]�kOJeK��J0o��J!"O�) IҒ~�$L�6�B�����'�,5�WH�o4��1�[���,�2tx��>�q�
)S���(A.$q&ԥ�f���RB�BBZ4t�!�E�/?t�1`�oܸ�r�`�'73
p�ғ>ɥ��8Jdr4��O¹����.T�'%ҽ��.�%)�uK�c�((���%�@�Si�:��O�@�+���dȔ{�D�Q1v �ӓb� q�!����`��!nmjB�>E��o�ج��oĎ2��č@�o�����M�[�D�O��C�5�r�{�ƍ��	]O��&#��j�P�����"�r�।@Ky�^�d�
��A���{r�*Y�̊1+�!D�| ����d�-?�U�!�̊��)��)�@���B�;�Hᵌ���n01��Ɔi$���0o T���s� _�stL��0� �����bK�P"�b�Xb��>����B&g-�!�'�(�	B�l�5Y�i�p�L�+��'<��	L�3�<����Z,^�H}
E*ˀE ��
ӏ�)x��ٲ�h�$W��p$P��|�&��:8(�$[eK��K��s�����Q񇙫Y8	$��b���+���)��*	{�PQ��)3��.�*ĉ�����g�,��	��.�
J!�� �H�_@P���	�&0�(B��'����D#b ��T���%2�E�c��W�� 2�FA�K�az" �*GU
�`C�\�y��
�#T������jW� ���;����%��M�4%#t$p������̛����hOnD��݈��02���*9�Jl�C�W8q���!0BG����/r�PQ� EZ]a�tb�%J@<�'��=R��Z`���?A��đ}8�Y�cE8}��II>=�t���B�@�DS�˞�z5����7}�@<9�~�}&���eo:U��,��W/L���*���<���֊X�(I;�� �^��ٸ�*?��cQ�V5N����G��ړ�.<O��T����;���1(�X����U�	��к��'T����z?��@B�n]L�J�� �\K�h�4#�Ne v9w�L�c��I�<І��	+Q�O}�-K��p6�4Ѕd��Qddʒ86�GC	�<�᫟�@D���>���nE'"25�N/�(���ORd�C�!z�(pP�Oީ�t$f����-�,�O+d�н0H�=0��QW}8�"O*}@��E;���& �u3�mr��OЙt��6 
,��q�S�|�:�a�'H�x+�`R;�4�'��	`��2�J%�G��"����	d�x���?���Q�(ĔL��� A��؂�l��W�H\��d��}�`L,��3��m��L7A�S��K���~'l�>٦�N$pV�!�H����W�-�La��/?�Ղ0�Vh%��ɕ�U�`�Z��,	�48y��'F����$��>�,-�b@ةbՎ��O�HQ���{tVq
4�A�WϾ5��@�u
����I^hq�$�9^�09YF��'�Px2"0fn���5n��ˤ%҅G"�?i�F�	^�x�,� Xa`�����eh���U�@��[��AV�;֜;C�%eRA��nD��x���H!RI;���:v����;� ���pf,�c��L}b�HYw�&�`um��7Ǐy��i�!D��[�(�e�=	�:&�9�OvA�G�!w,�$Պ��Ë�n� �oWu�z- ���(2�Ƞ�a�2r�r�I�l�X���F4b�	�)[D����pS�j��[b�=�u튗R�R��#�68�̄���[޾PqՀB-2��mْ/ܫ~�j�hUM��f&�2�'�V�K�#Ʃn��<��I�Tb>��v�Q#1פ�{�FS&w�z�ēm�B��[�0d,I',�Wd0푶kС2Ҡ��e���r3i�	�̀��B�?�t!%&��@Jx!O>���C��\�����q�У��,L��ԼG�~�Y���6>��q�B�N���F����w�Ȅbr����J���U	W?���	�W=����*#��p���)
�f<0�9H���K!K2 ��� JG��<���?�~�'�U6�(�i�e~��1u�%+G��m��A�	М��O\�`fN�`�\x�1�12�6�sA�fL�ѕ�1�mZ�M\6Y���xVG����$ӛo��
�,Ų�0<���Y�,Xjƭ�[R�)�2K��<���$dڴ�����0+��	�(ɰX�(Pz�]>�B�Ģ'�V��cIp����$��V�F���:G!�$ۻGߒ8`�N ��c�KK�ǢmJ�$G��)ȢbA��u�[�	�����|Zc�����D��`� �,/��e�	��j`�fl�x��Z�LO�j�e!S��<P|��N��W��4�v�ޖ2�|�c!�{}��u�'\ar����ڇ'(��G%�j�D~��͆�6,a���+{�T�O��\iT�E�s*H YAM֓ �����D�\�O�ɏ�Y�|��ȍ7_�RH�b,F�6z�h�t'?����mn���ɼ>�oĦ��|
CG�_����m�k�~�* 0Fz|�e��ݴ��9�hQ��,�D+�4�*^�+���� ����xD�h�O�=��P��P�M���*�F���tA�+(����k!�s3���aR��T@E';r�ݣ�>iߴ���a�/	���$ ,4ũN~�)۲��/[B��	��4�p7�9�O�9�2����a�y�`�҅`K�!�liY��8��Fb�B@T�s9���d�!@���ƪH��$��$ő<�џq�"	��6�����M�C;���c��Kz������o�.]jt#�D<����	�WR\�"3���6h��h�}�˓{Ԉ�+J 
	z�'��yC���C���'݀d#7޽ )�����Y�ӎ�9�S߄l3g�
���)(PO�>*�8	�	�(yA��'V�-Z� �oH��I?DZ]"���u���<#��ɓL�*i�晃� �:��O��9���f T�c=��3�R)��Q�]�qq�!aF �M;����	�����
�>��g~��G�$�j����Cf�j�⡋8�~B�T��,�WOy�d�PS\d���m�1���ۇ ��i�Z���(`�Z��
O<~�m���'�0p1�^�h!��V��$X�O�7-Ļ�J��� %�d�Ȧ�eJ�>��C�Dcbl�3��Y��H�'��J��@��C38`Ro^�1��˖f��<}0��Ҁ$��'3�$�e��8u �1�������%��d 2fCgv�p��ɡ[	(h"�l��"a1�V�����3���C��?`VH8&"O4�kԫɀ>���dl��~<�uR��O�0��$e	J��I��}�Ѫ�;P��q�F�7� 1c ��S�<��eɏ�  ��#ä9����$+�g��G�J{\y3�V3�0<��mU�@4j�s5��.N�	����U��, 7eJ6VF�4�(C2@Urr��)3��5��"O!���@������;rj|{�&VP'�� r��$���}:p��
D�vL[7��I��h��)\�<a��7%˜\�dh�nԺ@��Ryb��8��U�=E�����9�]��$9u1�y�V��!�y2`�D�P 'Ωh���r��6�y���H�xp��o9�}��h��y
� >P@�'�-V�l�Q�K˾D
Z\p�"O]`#��_�X�� _$��"O ��ͺ-����	�#
����"O���U�V��ґM�)8.,���"OLM"�F�|	f���lH+(Mѧ"O����J� zV-ôl "(7�|�"O��0m�C����(�C# 	�
�'<�uH��-8ZY������'rh�HF&��3Td��'����'�����?�R8Z�"
�ׂL
�'�M1d�]�V����N�:�d�;	�'��r�U{�P+'d�,<"��[	�'^}�+��t}Ib�+><���'F8ؕB��Xs�G@�?\���'�ps,
 K!,[���9��	�'\���F��e�x���8��2�'����F�74��'F�>{?�T��'��X�ņ��H�͘��|'ޑy�'�U����h0�tJD\�Ԝ��'h�š�f��0�9�
�^��z
�'�L�ۦ�fy�0kOـ���'�X�����x^(a0	�� ��%��'���8��܇t^�! v�8`]���'!
��ۮ|"@�9Wf^ uL�r�')�8�"X L��l�o�	r�'ܘA��6� ���Keɜ0��'�ܤR�X�B���!��]�L ~��'4��[D�p��T`��rl�E
�'��-��l�J�xi�"(o����'���k�NR�|8�Q�5j�?[M����':A�M6>V��eg�G/>���'���ZDH��zQ���6�6��	�'�m;/��DQ$�:(���''��B�S�{#&1�ӌ�(%�*qi�'���x1��9�R�X�Ň{�Q`�'E4xH�*��A$���$`9��'��(b��	܈Rő�gT�H#�'>J��c���'���al�7��7D��@R�PL>���(C$c���Z+7D�Hk��/RFd0��(s�L���5D��K�$�5'\|�)�9S�`xȓL<D�\���>w�>��%[(��?D��K�ۊ?D�!����p��Ģ&D��i�n��Ď� ma�<1��%D�ܳB��<�n$���+dqj�HB$.D�ԁ��:C�p�dB��/)n�zh-D���}a<E���J�h=Q��4D��b���@1DD��eF8NrQI�5D�PY�Һ��a��ţu�(����2D���a��*R����jU�5��0D����h��5 �uh�/S��r,J��%D����	q<���C�WA�`ɸBM D� �7&�t��BtJ� M[HSË5D��!0�fh��Q�Jdr��2D�<��.i\�DΊD����u�$D�H0dʠ6�<<�T̮?�(e���0D�P* ���*@� ���:�$���+D��*'���+�H� #+�>�P�b�'D�tH�����Z�ƃ�j�\�p��'D�ԉGьR�8%��Ñf&Q3B+"D���㋃_���͉+�!�
�n��a� ���a�u�!��A�WDJ4���O^t���B��!��C	b�����,I8�e��[�{|!�� =�lÀ$��!��b�'Z��a�"O�}�C�K�~�zW
�am>H��"O�iI0*ǸKkz�SQʅxF��!'"OX���R�W��[�^� ���d"O���ą.G�P��I�%��K0"O�2A-gZ�@tK9]���zR"O�Aa��V6p��E!���{���Z0"O���צ	!��U�``J.\y<��"O�"�B(��x[��יiT�h�"OL\�穁
&���b�;�I)�"O`�զN%��Q� !k�$�A�"O��qA	�֤-�&��'��=�"O� ���8��l�"MK.Y����%"O̜z�ǵg Ly��X�#b�$"O6�r��P�DKH.txA"O�9F�<Yv�2u	�%��x@"O�b5�AZ�쭃bb�ZP"Oh0�g�w�5ҳ��?4(
�3�"O�P����}\l����B�?�(P�3"O܈"��֞�ȥ�� =_���:�"O�\S��3y�Ȧ���}��t��"O�X�5�ސP���XE�g�̬S�"O��F�V�,�Z����:�^1*�"O���%�O�m�̜�ĦO<5��p�"OH��6���Y�j�ôG�+K���4"O����HY�RԫqhN3{*��:"O$1r��"��Q` �2�	X�"OLQ��GO([\� ��ϻX%��"OP0 @��Jt�ŉ�Ǌ$��xbS"Oδ��()9^>dQ0��N���I�"OPʥ�T+�L�Q�G�1D��"O�}�#N	"[Li�S�."�����'���h

�`^��K+4����A#�v�9A���yB��,E�]��K\�|�4�z�m��O�%;�,�*[�<0���IԢb��!)H��\���bX2�!�$Q)m$Ԥ�f�1t���&��"�Ɓ#BJVpV]��F��'���p,H6W^�-8�'@@��a�'�@A��@�c�ވz�-�y�����Ti��2юa�ӓ(A�z�.�$�|XI�92+r)��	F���Cs���-F��q/��-f�U���Q����j\`�<���^�,���FY�:_�ћ$i_�{�*��8��M�����
�|qc 	�Qe�Tദʃ�q��Ww<��a��wq�9k�� h-��[X�����#�:�'?���xːx� :�ă4i��"P*�96��*���B�!�܊6sT�H�J�W� �(Z�ǅ�`�T!e�YQV���O@�jB*�2���'t��Y1!I*Y<�AW>'�|��	�|�K��&w��]���{f�Ԡt
м\D�ds���cj�x������9��t��K���5�x�lH�sQM�ǍQ�D�j�J�X��O|��g�x�$����g����A
�`��� 7�<x�q��n��l�7�1���N7�S�O���ңg� )`%CCi[�/2~|�Ǐ�-<xB��"6�����!a��	^��D�N����;�^�x��
���4̑/C%ڥ�'E>����D��ϸ'fK�$�$| $E;��]~`�,O����m��pGb �I�b>URP��8]�����XU�@d�E�ֳ7|J}�j��$���	8n�$� �G�:-�B����5% ��N��*w� +o@ �$G�81geګwP��'����PF�Z�L���[�u�$�)s�'v��� ��MHt9 .0t`vÆi�<h���j�����ǆ��k�RЫFX��|R��<r|�p�5��Un��AN�^���&/{⴨&� �%HMm�|(�d�&y�D�Z� ��^���!���s�� ��gܓT�~��d��F6����&k�����ɑG�t`��'�Zq�E�ćS�n0�Ph��M"}�QA�4s�^LX�ǲ�az���K*,���+�K��}3�ϖ�����¡@���\ZU/[�}q��P��|��m��n��\�%�'8@b%D2�hOe�O�,/�zA����Ɗ�Fs�#��ؐ�dhB�.��$�1#��h��%_Xa��O<v<����h�"̃2
3�?q���
$ڈݰ�h"}���=� bDڠ ݱA.<���N�H*=�� ǥ�{;�t*� �3��
�n�`��G�J��5�ġ�"�I�o�>��.�hE��"b�91��6r�$ ��Ň;v^�jP2&h��I9qJ�h�*�3-z}h���4"����mU4;��Tx��'��I8A�N�n��Q�0���44���ݭ{��G{��6	�̲���M�'f}�P��!�Q�w ԁlf�$�T�W@T�mqOq�΀�c	ۣK�Ba��]<�d@D�'��%�$iB*�]�O?Y�e!�|�b�kc �n`#�Nl�<1udD8O�`�1.Ӹä[��sy�Ɇ�O�`�,�I�H	�D�~� !W3D�5�����z�o��8��,ׅ�<�H�A%]� �PG�n0x�ɣ���5|@�O�N��O��y�K�w����`R<5�:eB��½��O��j7+��hI+M�h٪,b"/�$����'ѐܰ�M
#%�yZrPX��X�JS!]��,1.�"��=� =lO�-�"�ҽb���BէF��Ir��H96G�yr2Ӵ`��K��;�X�O�F^Y��K�~L�Y��M9�	?'�ѸfL�}%| �
\{��2J��p6L݄��3яءV��%��!�f�!�$G$0����8�l����6jblR�͎OK���c��r�L�@ö��L��&R"���g?��?c.� �٧&\x���ͰQ\��(:d9���|�^	z_�@��D*0xiR�y�D	��F�,lJ�� �p��W�P948�D5��3焚>3.�Az�&��??����	�h�J�q�N")�p'oX�|�N<Y�董 �&T��͜+t����O���j�P��Ó~�D��#��U���ɑ�ƏGK�]�=YG�#�6�#G"�'������?%���;�f4ת� ^	8��Ff_�nq$�qq#��r�!��B�Q\��2��$��hId�əT�>�z��,eZd�
�Ft��i���) VHٙ�����9O��	mn�Hc�Ɠ�h��p���yc�\� ���_�7C�)��C� 1�(�E��\|�1��"Y]:��'�����o��"���'�&xs3�S���4+�[L~�
�fgTt��	C�@�Yض��iRx9c��I�D�`�˒A)D8��O�]�b�NT�Z	�} �sb��=��K��#
b4��?yd�S�pƄ�yʧ1@�;��qux�sӬ�)P��a��BɉTE�09w�7� �$�U-p��t3b�]�F�8y��$�i�b��E$���O;h���E����Jfj��Gr���'C�����o5N��UO*7�4k*O��(1�ֽ5��T0��P�O�HDx�)H� ���b�eK�/fz)@�'����(6�0�+���+~�p%`��Y�P�O|�P��Y���P� H�H�˕K��:�Va�7/<O"�3�n׮��'sf��3�Ŕ�����W0��''�8<RP� o�j8��K�mS 6b���N�2BGZ����P4��D�.�dQ9��k�D���~��U7@���&DU�c�h�� �� �y",P5,��eްh���@ �Ϩ}� �'Л���:��#t�>���ǃ+xJ�ϻ+��˅�O�$f����������ɹ-���V�;�4�S�M�.]Ǆ�8 -_9m ��[q	3}R���w�^`K�B2� pC���T������R!p�����f9��G\���b
�H����adiB eL�8ұ
��E�:5!^�E�>42f�Y8�|r��0H��|�@U�q20l���� ��B�W���l����+���q�`�	�TI�02u�	TK����`K������UK���L��L��`�E��+A����JA/���1T��mڪ�n=�OT��ѦSpɮ�E1���Ea�%5�`i{GaP�A	�`G~bŜ�N&����h{t�;~[ }JFÂQ��l�n�>b<ym��H�dP�O���d�^L���$>�#w�	)u��_�0��卒Y�<��+�2�BpgY�/m�ʓ!��$ۄ��dն�u�a��t�F�R���x�S�ч T�y��D��p>1ĥ�=a������.S�Vt�O�`~��i�V�+Qe>+��'!Br7����I��E�-&Y4e���͟77������<�Z<3$d�AB(��B�8�̑ӅK�)Hh4�I��;�'P�➘å�=��t\�x�1r�F�?�f�9��M���O���5	F%Mf����!���A�B�5� ��VP<�yB�E�QV8�&B**��t���~�b6�Ha�[H���&ՠ��W���<^���jD�o�C�ɺ!���+�ƍ��l�"�N�w���'4������z��	��l��d��iXp�Q)^b�����-+�,X�E |��q��n�� ��ȉ7��6����'��|��WX��A��pǦ1Ӌ���E�x��P�/�]�~\CF!׸y&���jN�Y��B�)� 2�H��Ǿ!_\��.Sx�ȇV�xaE��4k�qOQ>���G �!�(�,+���R�7D�b��
<w�V�;f ,���ɔ�'D�Cd+޷m�쐕 ���}���+D��ʆ'��z�8����_|��5�'D��%�T)W��Ŋ�Պ.~-��+D��:�-��W"Eshӣ|�hU۳J4D���	]8?�r!�e���	Sr�&�.D�PDF�4̥���@�f�:A!*D���u�
�ԦՑƋ��Y�MR2D����fG=F�����_�%L����#4D���愔>J����b��)rp�/D�(�Pŝ6	�PU8&�.�2A�Gf,D� ���S.H]�"��b�� ��b,D�ؠ�H^8
�yTl��G��̡��>D��"A�˹Z�\xK�֥&r�(��G)D����ք5���!q��+g��� D�Q�dA.C�Z��6��"fA �5D���E)>*2� �(�,��C�3D�� ��X)6K4��rM��8a����:D���%��a��I�%�^����:D�\w
�*p�X���a�q�м��6D���Y%��Er���"�}�����yb�M�c�a[��ۀ�*Gk=�y҃��bL��(��qX���w�@�ybh�)+����rΐ�j�)�F-���y����Cxp*��ޓ $H��V3�yBO|'��+��²Bz��ec��y��9Ud��� 	FJ�(d����y�m���!eN<
��X�C�T��y"��4D� ,كƑ�l�����'�y��K�d[����"K�fH�P���=�yDI)Q8nz�-�F�:1Z����y"J�-
�d���$G�H���ݞ�yr�˒{����χ;;t�����>�y�dP}P��1��
2%�����D�y�/D���f��3J�����W��y���W��y�B�ߕ8+�������yo�)pk���׃A�M~�Z�π��y�I0$���g�
:�L}����y�mK�OUXdy%`�9.ςYa�̋�y�뜑0�| Ĥ[3&��C���y"E@J.h�PWi�3R���KM&�yBf��x�s �\8[CV���̇��y�KW�t�PL�0mh�^��A&��y2��P8L��1OQWl�"����y��βh�� RFJ����h���
�y��Y��R�WÅ�&q�ƁQ��y�L� �p�R�n�!�m=�y���'����VQ,����h���y����r9�CS�;�� $��*�y"�;M���뗦��Jc X���N��y�MģvZ�3��РNrE��E�~�*�E�c��'Θ' ��qգ�		�L�:$�߅�z����W<(����$��ӧ|@ht`�K_�ga0yW�#Cy��v���p&Ӈqt�5:T�0����u��4u�� &�;=�ٗ�9Z&�I[W�Яap���\}ha�D�ג-*d���eU�[��h;�:~)ѲbF:]T���6C�ԩ��	�|j���'5���k ���:R!�E6��xZ��:�xn�C+&�`�Ok��םK�P�ь&���FB�L�hUx#�+	�ɀ�AHyB�͸4�a�$I�yH�$V�ث4�ʻ�f��/OZMHr��<+����I���J4��a�V�qc�ϥr��I���}R5�ͥ>�șG��o	�zC�4j1'ȥL�J2r�CĉN�dC�0b!�%L�H1�$���~���G6J��� t*3�z�G�͈Qx`��ʍ@�@5{��ԟqO���v��H��`!폐^)�����nv\d�?E����� ���C��{($#%�4E`� ��.4�0Z��� a�|1WH��T�S �6D�@ R�L�.�"�ˑLQ�So
$˂h'D���b�,ڈa+f$� 5綰�Ra'D���Mō;��1�EO��'���ô3D�0YU�2&4&k`��IF�(a�k1D�` �y�-��j۾yV�;D���@�k�,�Zc�-F�L�c>D����
�u!Xaۦ.�"���J��0D��R	���f��"z]SR��yBD[�X�D�+5�ܖ�:ػ! Î�yڄ<�Č��-LM�}�m_"�!�Ҍ7��IQ���|�l�q�LX(}:!�];i�0$�q��>&�H�k�(!���bϖMB� ��@�#�B�^!�D@�5��y���ߤ6�B-)��B:
!�ě�l�@)�b�w=ʽB'�r!��ӕ?l�Q�I�Ĳ8�@�Q��!�\9)���CDA�_�:Ti5	V8�!�$COC�tiG�]���kĺ�O�!�Ǧ7����DF�\y�ȑu*W-]!!�$G#̝s��][����F�7�!�$�-s�ڔ ��X�lX��@���2�!��Ϥ1������S`D�,h�%N�J�!�d�g˰P� _j�" /J���ȓ~12-�3f��Q���8� �S���ȓND`��ߧ0t�<@���T����/k晩C�ݍ<�^(1ʛ�mQp]��T�@4p�蟬_eT�����Cl�ȓ5���S�]��KPL�/N5V|�ȓx݊���*E�Zy� A�,K*q�
$���f�(րN .lR�����"\2�0��~�V��cɅ�}'�Y���HK�̆�"��X1����}�x�[�� �u
��V��0��J��"&Ή{#(�G����!�%ˌ$|>�;r��T�؄�u�*/��q�d��B�.ZB�	 $�t6�[	Y*LQ�)�0B�	�>X�A8���ĥ�^6�0B�	�X���Tg=�y�S��E jC�	7KL95�m�<� �P�a�8C��T^� u��64 �ˍ�rB�	;'�݃�gS�5#�b��17�pB�%*��8{ƌG�J7�a� �̸5qdB�.e��)���\��xs�ʅ0*B�I@�� 3	�;|���QG�6$�C䉓	D�(
'�Ǝ|�8lRÿxDi�"OĹ���'1_Ҕjr��#&����w"OjIcW�S�i3��ٴNY8�JZ "O؉���VO�)B�,e{<	#g"O�T(T�u~�]��,[�e�Q"OF�fLQ�Q�0QC���DJ�0"O�i�R�?T 4��GP6C>�U �"O���oء<�F���ɨU�$��e"O���`f�t#�����i��"O�4`1�[�P����ǃϓ�f��f"O!�f��C�( TƯa���چ"O ��M�F5�ip�%��s���"Om#���9�*��O�w�:"O��CB�|7�1�4c	�E���"O�}�SgD"�rQŢ�KN���"O�ur��G�r%�&�H�2G�0�"Or4��lP�i��顥@�E-&�""O��8�䒁���ʦ��D�,i �"O� �̡1o��g]�@0w�A��\�9c"O\�Վ����TG�A�!s�"O�t��*T�~�rٓ3�F�]m�0�"Ot�	o)^�S�E�SSܱb&"O4-R�`¬K�����o�"*3�=��"O��C��% R�ı"�M�Dz�T"�"O����]�A����r��GA���"O(�Q�'f�j��%#F~/�ؒ3"O���p\�f4���!�vh�'"O�Y�� W\�l�� ?%���V"Op�Y�NT//r����ȎIVu�U"Or1��ߎo�X�i���v�C2"OH��פR�F���GD)X�`1"O� @*â*�H��D�J9z��X�"O�Q��m^3|�((�Ċ�Y�6��"O�`��'D��"C�>^����"Ol�W��T�^]�`�#�D�%"OD��a�Y�N�h� 7h]�g�Ċ�"O���S ��������O���C�"O�C�ř�L�V�pqH�{�l��"O�aQf�V�dߨ��MƳ�(��"Od��Ӎ�"PV�\�웑aV8��"O@��S�͛&q,|��iL	��Ъ�"Op���
��/V�}*f��I��E1E"O`� ��6��l۲bG�X�LQ�1"O�cc�]95H�]��d@:9�pI�"O���nh-�u�^w)�Ixt"OV%z�K��B��2g�ٸ(���;�"O ��vaE��A��y�dݻ=�!�E�;���WO�8E��U�$�3q�!��۽z殘QѤ��:ǈQF���!�Ę�; ^��5*X�'`~ѐ%V�!��#|W��c�L��@�$ݪ��1!��*傐�`�$ ��ID�.X!!�$G�!p�T��+ZM!uٖ/���Py�g�0aL�����=w�� �ܣ�yR'�."vܼ�@:ߔ�A�I؃�y���d�4}�"�ڢ/���6-L�yb�7@A���G�VOV�5�ڠ�y"nK
�\�uA a��ᣐJ?�y򧑰~TXxq� ��W�=�����y�(�"y�Y��C�P `pq�P��y�"� J@'�DB�c1��y��~B�ȐA���4 ��)��yG/�� r̝֠C���j��yr?a�6��pgH#r�
�sf�/�yb"E�mQƩ�7�ϱ2S��Au�*�y2� ��ԋ�J�&������y2��		�|并��J6E�5�Y��y"!�}���C_=C�歩Dꞛ�yr��(���[����o�8�''�y2������G�%d�
<1���yRȈ~L��*�D�T�8y�&oY�y�d:���!��I/��' ��y�ݠ/(���ab�=BY�b`튦�y�&*�x����Aњi2�%�,�y�p,�@��f@�2r4�'�C"�y��K�"�𨢱N]�#(
\�I�yrΆ6~,r=Q'�Z�+�d][0C҉�y�h���¤�7����۠�y�M�b)Уů7���7"��y���C�:�Q��V9M;HTs,�$�yRo^�R��;�K��C�PĉP�P;�y"D����@U,-B�m��@��y
� FI
2)�B� mJ"�A���#"O�e;K�<~�h]2�2�~t{�"O"�@&��,q����#D���a"O&q;�i�$l���?��8�S"O� @���H�b��&&��A���zd"O` mݕTKDp. ^��T��"O���W��V�:Y�C�2��|�"Oԃg�ʄ
��YT�]��!B�"O��ᔧZ�1c���hִ
y�8�5"O�����S��Iqh�6{v�-��"O�<jvjϝ�r}I�l�KZ�	[�"O����m �mڂu[��@�\<"=I�"O"��t�?gk8���b�4!�E"O�1��a�)r�� ��Ԙ��("b"OR-�t�ça�r��V�_�x���"O�����;C8��4�	�۸��"O<M�3M�"��2�&д_��Z�"O$M�C'�4y���U܈��"O��� �&i�`�̕�r%��"O�-p1"�TF�h��ԲF��Yȥ"O��AE�1Avjl�-�$V��"O&D�aOJ!�0q��N>"M�QX�"O�Q�GM�q �%�!H�-���"O$I7�11Ŏx�aK/���
"O~x�¦�&.��� ���5 ׸�"Opt�Ť��"L��(ӽ#��ec�"O<�t�<N(��DI��B��)��"O ��F	�,]T��y��\!V���+�"O�����4���ph�J��s�"O�l��ϔ�}!���@&O�D`���1"O��RG'�\N~HK�˟�~D�P;e"O������7�>�J�[(�P4��"Ob�B`ES�y��c���w����"O���բ��6�Y�r/��V^�|"OИ[w���?��R��VP�z3"Ou�ˏyv���&e>E���w"O�к�g�*h���f"�f1I�"O0�S��!`j<p`��@�vH�D"O�q�P kF�M���YH�&��t"O"�i!"kύw+�40��~�2��t�8L�@9����e� �(�ȓ{�,��u�хb0`��MEh��	_<;A�?`�!#UE�.u���ȓ	� �qUO�u�zp�tn�..ߜ��ȓT���iڠ������,W�P}�ȓR{����O9Z�¸r0Ǐ�FG���3��iJr�
kqX���D9TeHB䉫|��(S�AD�Y#F�bB�I%>V�$
�fߴ΢09�@4EB�	Z^4���"��]�x��c�	C~�C䉶-�:HQnY���f�z1�C�	�O,������E%b ���L(+�>C�I�&��xg��T�\����E,"�>C�I&j}�j�'�6�����0d�B�	�	���j���3E3^��4c��P�C�I8g�|l'n�J�H�ӆ�_0hGLC��-=΂��g�p:mܾlфC�I�F| �E�PG�	�J��R\B�I�*҈���.x����ZD'HC�Ihg�a�o��4�\��@��prC��G����3o�>����܃JC�	�Y+|��qf�(C����5�="�DC�	��8Zc��\{���d�ٻv.C䉇e�<�jpn� �����h�<6\�C�)� �I��j��t̑;e!�1@""O���fD�3�4!�u���>
�+"O� sCʗ+��"�Q�}�n5�"Ov�É
R�4�._��L�0�"O�Y�B��j��.��.����"O��#�   ��   �  @  �  �  *  �5  EA  �L  �X  �c  `o  ax  6  E�  %�  i�  ��  �  G�  ��  �  E�  ��  K�  ��  %�  t�  ��  ��  =�  ��  ��   Q	 " � 3! ) 41 �7 6> zD �H  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C��'��'�ZI�`88y�)�3���y#���'���<���I6�r/��{�rD5�S����t=^hg)a�LU���ͤ_�!�� �!Ʉ�P'^r� ȓ*T
T`��Z��	j8�ە��4:Y�}[1�R�I_�p���0D�|z���Z�	���)_P�T%-D��z0C(OUxPSR�П%�p)8vd%D��Z�Dòc{,���ù�4)��%#D�y�/��@m�(R��͚'0%+�( D��)�+G�XX��ѯQ�|� �!�p=��1j��#���"k�p�&��U�'�ў�!czؑ)�j���(�Q-L>��
�'+��*3�u���#��X�>U0�%ʓ��	2ʓV�ɨ��,PJՂ���+=vf<�ȓ)��bǚ��!C*T���eXP?��'~T�	ă�<'^rIa�l��y�t��'[�+�N�dq��C-�!����'��\z�E�"1���ń$ >�!��'���ta�!s}����J�d�yq�'HTt�M®@�����	5���'�nM�%�� Q��C������(�'
�(١Z��I"�S�ud�{�'�>�sB�ۦ��*_-~EY�'�@#��W?UB�a�6�޵jb���'r��H� �C�2���2j�8��'#B��ը�%�6��ĨГZ�t3�'�T���0� 1�C�ĔB8B�
�'���A��j��hF`A�>>D
�'Z S���&h���`tTy�'����v̏�F���{У¿IC����'���b����2r�\z���>���!�'w�����-<x�'#2E��(�'����P���y)
����ՂY��a�'��s���H���d͑�H�a
�'l 1��8��-A�)	�'�"���+�؝���	o����'�� s����W�8xyB!��9��'�
Mq]�
}�UO�Wi�ܠb�j�<����܃��Љ�Ҹ���Z�<�Ѐ N*5�waC�*�
�c4�	W�<q����!/�)�V��~t{2iO�<ɥ�-O��Uhs���sG+�@�<��Ёcm����҄{ӆ�Ida@{�<�B�]�G_��qP�D:,�Ԭ1S�w�<�P̔;+�u�e�F.:"�$'`�G�<D�^L��t�&�O�E7��sa�l�<9�^� �h�N�� j�XՅK�<���YR[�$ҁfK%{���� eP|�<�"+��x�����ƅ�p!qz��u�<a���%x��a����2N��3�J
[�<�D%G�y�Z��5bK�8�`��G�Z�<�@� &|�d-B���D;�@DT�<Q�69D���@;I��<3&�_G�<��C?*�Ҁ��"�:T�p�&*��<9b"�/+�hd�>l�,٢pYA�<�2R�zD�� S��<>b-yg!�y�<q�+�)0�[�7y�A;�K
~�<�C��*�,%A2,�wExݢEώ|�<I�,��m��S3ŭH{�T�&Kr�<A�	J@_"��q!]�~���ӗ
Yo�<i��T�|�D�A�(�r��|�5Mo�<a�ß�>�2��G�p
t�D��i�<ᥦ WFp�̓#] V]Kj�h�<	B��:(5���U�����9��#@�<A�A�n��T��fir�<9f�X�0�n�"0fC38�y�*Qu�<I��<B'�r���y(0	{D��f�<� Ƥ�4��l2%(�ʀ6R��5bU"O
��Ċ�>1D�8��ѝ%�R�:"O𘛆�J�a�(��#&�*W�A�"OtA���A��(!'�6Q�d��"OP
P��IU$���0)��R��' �'R�'g��֟,�����g岽i�m�4�@�
;Fm�$��ğd����D�I�����䟌�I��`���u���7��R%��" ���	�������$����t��ܟ���џ��	"	J���$JE�q�����B���T��ΟP�	����ԟ����������|�ILؼ�B�݄5
�q9򉙾O�"��������ɟ�������Iٟ������I=F�N�B���N�nMS��y2�����	��T�	���Iß���͟@�I�wM��32�<;sE�ֆ��+��X���4���\�I䟨��� �Iϟ��	*��ih�!V�u����gj�I1re�IߟP��˟��I�h���0�I����w4Veir��[`��B,�98�Iɟ��ȟ��������㟸�I��(�I>M/�m�0���`��2k������?����?���?����?���?���*;la�E̗�5���=r8�����?9��?	��?I��?9��?��A�X�:7���[<1��ð\A�����?����?����?����?q���?��{�
����1�vhA��%����?����?y��?����?�µi�"�'��X)��C��A��(Ge�<A�����p۴O��5&K�8e���1�E�o���;b)S~BAdӼ��s���_�&�˓�Ț\S�:�� H�m�I��L�4����'��I��?᧟�qct�]�)b�'4�p��$�Or��h�n�b�ҥ+���(� �-~�3�cN��5�E�2�M���w��I�&��VԼ1��X.=9:H�"�'*24O��Ş
P�ش�yB])j���Y7��1/8 Hvo�<�y�;O��Ʉ`�ў�SşP�c41�y�!h#��f�B�<i(O��O��l/aL�b�`��H7Kf �s+�쁷BV��)��	����<�O]��������!O��9���X��8C�xsc�>�ӸCr�^��Ѯˇn�،�u@�L��P�D��qy"^�T�)��<�C+� �w I8.�$�b�F�<)c�i-Th �O��nY��|��,�5D��� �HxC2��r�F�<A���?)��)g���޴��$}>ѳ�'4ׂm��� mH��$�(��8�8�$�<ͧ�?����?1���?��C]�h���"��߀z�����*�.��Ŧ��u
F������%?��'\B�8��K��;��`\�J�O1n�M�Пx�O��t�OIZ�QE�K8r��b-P�j��J�Y�L�D�'#6��b�I���$����8M$� H,O���	�W�
!��iE�OWDx�b�'oR7M��I���e�)���g�]��	��MÌBϽ>!��?Q���R��PW�Dh�pb�XT��(aI��M{�OfQ C=�r�<�I��@��'B+|gဥMNI6y 8O �����~���1�I�+$���S$+�.��?��i�&��̟��n�l�	�r� �@�%�~瘑y����$y8O>q��M�'v?.���4��C9# ����ڙa>�+
9d��S$ʚ��?��:�D�<���?Y���?Y` �wT3�e�(d]�L�W.
��?����dW�=3u�ןh�	��O\t��ա'lfj��%����a��O���'��7���}�O<�O�~%�E	
P��j��̲������פ]Ь1X����Yd�i>-���'�f�$���U�B�G2QѤ%	dH�r�	ȟP��ӟ���b>Y�'�7m�"��|⥫�3 >T�)��25f!���<qT�iZ�OL��'S7-�K�'���Q"ǆ2d��� ��w�V�m�4R�tm�]~���5'�����w�)�;�H31��.�E��c�����'s�IL����ޟL��g���
�4�{��޴o$�E��똅��7�Z?S�P��?��$�z��΀�ViP�ص��c�bTR�>$Y��٦�9��x��� 9Z/��5O�lB��ő,߸���A������S>OT)����?i�;�D�<ͧ�?Y��7
j���D�)Z�y*Т��?y���?I����d�Ȧ-�uO�ҟL�I��@ĝ�8g��@W��m	4���q��t��ܟ�oډ�ē6�Sp�G�#P��5o�b��'C�H��˱�2�
��d����
��'ӆ9� ��  ZH�Ǣ�����T�'��'"�'��>A��?��r�W�"E��:����T���I��M+Rn�����Zæ�?ͻ`L	�a�(za$]���;oP�͓0�Fl���n�~V
�o�~����w�>���( �����,?d�	 � W�g!d�e�|�P�\��ǟL��ǟX�IП����+#��%��R|D��K�py�G}�l$*�O���Ob��󄓎rZl�CĈF8F8�8���͔4�h��'t�7-�æ��J<�|�f� ?U8DXh#� �Ɨ!D�hkR%ë���U_������O��Y����r��,��Ȩ��&8��*��?	��?���|j*O�o-Lz��I0�ĀBe;���P� R�3��I��Mˊ��<Y��Mf�i��k%��G� ���3N)h�����Mƛ�:OL���?p��''��"�{�? �8k�f�������!��p�6Od���O�D�O��$�O��?)RF�LQ�$��"�2�X��ß$��ҟ `ش@о%�'�?q��i�'�h�x0��7vX�`�HĨE;�y�|��'��O�9նiR�iݥy�N�,��͠V��i����BT=���Ijl�'��I[�x��#�i��<\5KZ*�Ex�}ӰP�`̨<q����i�� x��ϲ)�$���� ��I��d�Oj7Mw�|�t�	�P1���T@�-���:u$�Mתq�%U��ł(O�	��?k+�D�l��&�HܹW\!E�!����q���$^�����K
�hن�9<��]�'=7�+�I���l�`�p��ci4qI&j���`��On�� �V�Z6�:?��Ni"�'#jfʓHӂ��Ј	:̰���a�"���Fy��'~B�' ��'aP>�4K��K$ֿp<pp2���J�@�l�$7ކ��IΟ��I{�s�\�����G��(��-,�!�����
��?����Ş>�<0��4�y�#W *X���`�G�i��-���y�%H�	'~h�I N��'"�	柜�ɽ,j���Ɠ��F@��/� ;:fx��柬��ҟ��'ߢ6m�5q"��D�O����1k
}zr��\;�HX
K( 㟨éO�un�	�M�b�xR(�B�v8ɦ΂8�(�"@�9��ĝ/��b$�_5x81���"�r8���s(|1�I��5��!�� �$�O8���O^�$:ڧ�?�ׂE�n��}�%^>3���f���?�Ծi�`��GV�h�ٴ���yw���0@T�fʙ<ny���sK�8�y"*d�<oZ�M�����M��O�8Y�'հ��בU5}�Hߋ6���!�Qz�O���|����?A��?i�� >h��/�oU��z�,��5�B(�)O4ul�1(>��	̟���u�̟T9�)	�|DH1E		�4���T��$�O�ox�)�'�l�Yaj4�M��M��=��=��ϖ��:��'��K�i�����Ж|�Y���c/3:�ђ��}��R�C�Ο��I՟��I��SvyrGv�J�S3��O��dD�m�&��c��%���9���O��l�D��w:��ٟ��	ן\�rb� u\���	}�p�0��8�l�l�n~��ش6�������O��F��̲tRB���g���p$E�	�y��'&b�'@��'�R�	H��uB��"�T�%�98�ʓ�?!��i1���ɟhn�{�ɼ&�h�"2#Тa�@EDH�3�2�'���	���Ɋ1�p�n��<q�O�h��f��#J|m�]�4�����A�h�q� ���O`ʓ�?	��?Y��
�
�����X��D�h~���?,O(mmڸ{J����<��v�$�[.jW�Տ��i{ ##
M����ZG}""m�$poZ��S��$-�HH�7d�>����FZ�M2��`+϶u}֭�T��+=��F�@��3�dEn�Qt���î'���	����	ݟ8�)�Py��eӴc�9���A��(iX0��BQ	N�ʓ1r���d�X}��d�T�jF	��b�!t́�@P0i�D���jشf3�$��4���WS�^��'@�ʓ3^�%�0
^�\15�%㏰�"�ϓ��d�O��D�O����O���|� mR2r^���`AO���Q�ùh��hn?-�y��ßL��F�s�ܰ���s�(�-q��(�ޤ%P�@�Jw��&�y�	$�b>ݫ������ΓE^t=�%�N&@B� �?��\�Zr
� Є�O��I>(Oj�)H���	HS �1�59�i��I��MC���)����O��d�J0$��3B��Xg���+�	:����O��D)��1@~TE�ǁL�(�k�"�-Gt��)8��9PP�@�[���&?a@ �'����	;3�u�%� )|x�@�D���rx�C�I'#y���d�5Τ��w�]4�zA�	8�MC/����զ��?ͻKu�Y�$���P09�m�cJ:�Γ�?����?i�̏��MC�O�.�iH4���<�N�-�X���B	c�&d�u/G������O����O��d�O(�D͖.���E�ڍy�$*f���!��ʓI��)��B�'���'��y��P��PnJ�v t�p�+�>���i��6M n�i>��S�?%)�K]�*��p�Ƣ�w�4�P��C/����k�ey�CA�#��I�u��'&�I"*���$ȩ�V���̃$y����ڟ���֟,�i>��'�6mK+��DM��uY�k�'F����`Y2���Ӧ��?9�U� x��F6�X̦�C!iن=_XH{ecɅZ��t�&G�<+J}m��<q�OМ	��B󟖰�'����w�<B���g�l�22���#l�T�'���'���'���'��\�%�ǎu�
��B�40,PJQ��Or�$�O��n�>nH��'�`6-*����i�Ih���+2�u/��Н&��bٴeE�6�O��� �i��$�OЙzs�F�q�r�B� B�/��*�TpZ�>��OR��|����?���3�H���(X:|�CW��[$�h���(s|X�*O�mڗ7ux��֟����?���e��eX�m��c���e'ф-��	Ɵ��O���v�(%��ǟ���I�h�xq�v�;#�Dx���"�(���n�� �'��4��̟�|H10��IʚDP�iq��� o��'���'��O��i�1�' �	�M��F�L�^�&��SY�4�ǡ���f��,O�hm�}�	���ʪO~�n��*�-��韍l���r�"�Vp�ڴ0�֡%\뛖1O��$	�R�xh���{���S�? �lj�GWJ-@��$���S���Q@<Or˓�?i���?A���?a�������%�"U$h�f��2����`�oڲ>�X���쟸�I�?��E�jybEx��Ε/D�fU���K%cp���[�T�^�D�O��O�D�O7��`��!�v1Oh���	s��m*�X�b�a+�8O������?y6�3���<����?���6j*$�d̽��� �_��?����?�����Ӧ�P$Þ֟�����\:W��={��J󈛓M��m)g,Rd��9��ɭ�M[��'��'�z�J�C�6?��0�1	ɀc.:���O:U�A�E�9��t��*=�Ʉ��?��
�O�y{cA�W��8X�B�]D�9�*�OL�D�O\�d�Ox�}���JL�����N�f4�珔2M4q������ն�R�'��6M&�i��(�ݜR��p8�hE�x���(|���	���	�Aט}n�T~Zw�x����Ou�q��!H�Bn�YW<p�h�4[E��|yB�'���'��'&BO!'[7��Y����/>L����M�oT��?���?9J~Γv�tZmj�r��U,߰0S�L�b�����	Y�)�S�TjZ#��MwH4�pC� �cb�)	1��C�5�'f�ሷe�$�F�|�U�$��`F7:�%���_�{�*��ş(������I��SMy��l�����a�O	p��l<j�HA�x�B��0O�nZM������M@�i�6�ש;�HX��K��K�\H�,�6�2��0m� �~�@�e��P�>���6���Qw��S�������IݟT��՟��I�����[��$����~�`���N� '�h���?���|d�֮W���T�'�V7�?����|�z%kӨ� &�h��ٻ,��O��O�ɐ�	Ӱ63?��Q�R��5G��IcA�-��0���9�?AQ�9���<y���?���?�""ǗX��|�t��&Ψ�򠐻�?���D�Ѧe��Ƌ�����ş\�O�ZT��+���[gC�:+tE�' 
��?����S��h���	��A�3/�X镆҆h��!� L�VT��]��S5�\e�I-�p��c�B��c�IO�Ƥ�	ן���$�)�S|y�Ej��Q����j�xHXw�*@�h�+�"����O��nZm�2��IƦ�)r�[�"t֔8�a�V���D��?!ڴ Y6lC�4��d'k^����u���:�6�	ގ)	ni"&$	2\j������O���O�d�O���|R2lT�1x��냩]O��㖫�;����V�py��'�����'�P7=�P,�٠�"Z>����E���<O*�d�O��O�d�O~��X�D�v<O��U�{RJ�*�E+^����7Ot�k&�E��?��
"��<���?qQ��+C��6)� =N1zb��?���?������覙�G�͟0�	ٟ���- �n��	{��Y+��Pm�I��5	�	�M��'��'��p�&�.t�Htg>��(��O��(�(^CD� b<�)X(�?Q B�O�e��o<7bj�'��0"�!���O��$�OD���OP�}R��g(ʐya�Wa��q���­�4��fk˭.F��'�r6m-�i��zFo �G�`Y���~��a�ej��������ɏ��lZo~Zw��q��O�0���ˑ5݈����l���[�`[Q�IOyB�'"�'f��'���6ly����߬Sbt�!CJ3/A�	��M�cM�?���?9I~Γ3��S��_(�� $'RphV�z�Y��H�4 s�F.-���?�Ȁ�vO�6|� ��"�X#�q��eI�I	F��b�'ߒl%���'��$�5Ɏ8�h K���}���'��'�����DP����47jT���I��LI�F.����I`����Fx���TZ}"�'��'�
1"&Nʦ0�d�Q��)�V݋��B�S������[�*��C��)Lh��߱Yc��L��w כr� ��wex�8��ן��I����ڟ�������p!K�+ڢ�Kn���?9���?�"�i���ۚOb`tӴ�Oҁ����*G��Iơ+����n=�D�O����ON̠��z�\��X*�)ڀ=��hz�,����q��^<����R���O�˓�?)���?1�o ����ȕ�c��*Cn�A�%���?)O�$l�M*@|�	ȟ��	E�DD��	�0�ūġԍc�ȝ�j��	%����O�d!�4���čy�$K�A�8fi:�GK�1V(��gC=�h�cj�<I���
��)��:�H�i� S�=G*�$!��Ԕ(���?Q��?��S�'������ɄI�]���f�S�d
(sӊ�fi�'Ͱ7�9�I���Φup�\�/\0�	��.iT>X#C�C'�M�ӵi�D�Y׾i��ɜ.�0���OQ>p�'/ތAUc(� ���(ډ�aۛ'1�I㟬�	����I��|��e���
X��E��Z�_e$���?8��6�G����$�O��6�9OЕozޝ
�D� jۨ|5$V&��=���)�?�޴.�ɧ�'DJ��޴�y�$R�b%���� 	��x�*Y��y�/֤,��-�ɍG��'���������ZB�Я�|b��l,I]�	ӟL�I����'�6m�*A1����O6��¾ln�U�C�Q�g��+E�U��"��O�Pm��Ms��x" �e<�QjP(� s��DoX=��$P�L*��Ŭ�0xP���"����zP��c�Q�P� �WIP1O��$�O����O��$/�I�-j���O�<�E�u�p5dOL��Zű2��O^lC����러Y�4���|λ\rd��P 2	)f����Ѭ��4nZ�M{t�i�t��0�ig��O��u퀡���� �bGL�$w����!�B�L�T	�V
(��<	��?���?����?�5��+:�����G�7���Ҕ�M��^�AI���Iޟ�&?牺(��YX�φ*%��q��nGJ�O����O��O���O ��5� ��7�{LQ��ܩ64��bYzM��r�n����O�5�I>�,O �醂�u�&�1D Έ t�� �<����?���|�,O�m�4_�H�	
F�<�e!�e��}�G�����牘�M���D�<���MS�iT�X	�AL>e#���| �[�+ۂ@͛֓�(��f��0���o�A���e[�F�9y�8����iֹ���}���Iğ8�I̟���蟌�)Iʬ��n�*zB���
8�?���?�e�i0d�'P����4��9�D
��:����fH�y�pm�s�x�Im�f%nz>�%���e�'v���ّcٮ�
 E܂Q$���L��_Ֆ�ɬ �'��Ɵ��������)��T([�.^hy��M�!� ���ןX�'*6M�����O����|җ��=�n��2GO�i0űf �d~G�>�r�iz�7�i�)J 
G��0�)�jS�Ap�iUkȢ�D�g�T�-�<�I.O�)_)�?��G0�$=q�&AӳM�P�rP��*�=~r����O��D�O���	�<���ig>��Ħ�wh�
׆ȳI�HQ��׵Jn�I��M���>��i��u��� ���&��*BEH����~�b�m)b� uo��<��so��`l�\z(OF�����<s�4��}�5>O2ʓ�?��?���?�����^?u�d��F�1+˦D"���!�f�n��c(���՟��	}�s�P�����u.�%��ܺ��.���"a���	�UKM>%?���Ϧ��+0�1�K�{��j�$Ù����%h׈�O8��K>I/O��$�Ox�$��$/�,��d��:i��hPPf�O��$�OV�$�<���iY��1��'Gr�'0��[ဂO���K��sܕ���d�}�`��hoZ.�ēa������>lƤ��.�xB���'x��K3ӆ��������gǟ�"�'���	!�O:��P#j!�+g�'�2�'�"�'��>��� &_�I�t,�?^��QF�1!j�9���MSB.��?1��]�f�4�.�(g��<��DsFmփ0x�1O����O����v_�6{�D��9p���wfB��@ �$}t��b���`9c-��<I���?����?����?��0��� ����e)�������]�ua�՟��I���%?��1Q��P��߃Q/*��v�ߺ䒽��O����OғO���OH���	Q[�H�s �gn���0�	�T�QK��?� �$�⁦�O���J>�)O���完%fTE� J!Z�ژ�)�O����O��D�O�I�<�ļi6�T�t�'���*8�vA0�	)~6혙'��7�0�	���$�O<�D�O����E [b~ؘ��H8v��SR�C��6�{�`�	��R�H��%�<������e掯 |���0A�	o��d����<��?���?����?���$�]gmF��*ɬڅ_zR��`�'i�'��7M��5�i�Oam�q� ;O^�0'�3r,��� ��" $�����0��;�0�n�<!�O^�Kt,�!4� a�VCt:�蒸E�r�H@�	xy�'_�'�CT%7.`���N�|��]�@	���'^�	4�Mk�C��?���?�,�l�+_gi+ƞ7P�,��AO��"4�����D�O���!��?�b�=d����󧎠Q'�;��B l���'R>u�)����.�ޟ�Y6�|��W��$�pʊX68D��AM ��'��ϟb>Y�'e�7�ĸ���j#�K�i��xr��h������O��$�Ħ��?�3P�����H"ap��ϋ;3FM��b�!p����ƟX	5����uG�ώ:4�db�sy�M�S&	����G�~��#��ybU����ǟ��	ݟ��I���O�"E;�`��S*A�`�� �B0�q,{��,�e
�O�d�O����̦�ݏ-��$�FDՐ!ĸk�ꉪ7\��ڴ$ޛvD ��U�o�7r������q1��LI�e�:,��f���(H�`��b�Iwy�O��+�y#�eA�M��${.�ȅ=�2�'���'����M�!Y��?y��?� Y���И⏜W]H�����'���Xɛ6��X}%�຅"f]E+U�փ]�<�F��	��$ �J��<��U�䓟�0����r�B0w����P�&E��@�����Z�j��Od���Or�D&ڧ�?���'�� ��Ʈr�Ĥ�"�ڲ�? �i����u^��K۴���y'F1J �e��"f7������y�Kb�,�m��M�a
ٯ�MS�Onh�2���FI[���Z�_(7���
����O���|���?���?y��p���b��Ay*t+�I�^e��2.O��lZ?����	�\��b�s� ҃M�ͮ���̲c��$Z+

�������3޴E)���Oo�4�ҭ��Q���Z1��@�>��oN�"���X�.4���O�tN>1/OT���玨Mz��1dǒ�/XV�+��O��O����O�I�<�i�����'�p�S��[/j����L  �5��'��7m?�I���$����!޴]:�F)ؙ&�u;���Q��!A��'Z���3#�i���lh)�O��&?A�]77�)���D����F����⟜�	џ��I��`�	f�'0�$ a"\�tƀ��DB/v����?���K���ՃU`�I��M�L>��,���h�K
9�8���Xʉ'�n7m����4�� o�e~b�$ƀ b��C��"&�>9��S�_��#�dE�?I"�:��<���?���?q7��:t>T�;\]�1�QƤ�?	����N�M���ȟ0�	���O�Rv�>\\i7(.e�d��O~��'Jf7m���L<�O��Iȧ����ޕ��-?d�B�)�|ҸY[��5��i>!��'%�l'�zD R�Z�`���K4�^�X M���	��ßb>5�'Ŏ7G�~ ,e�dn��OX�V���a�� (˓5ћ��dp}�{�e���v94P��#U=��5BA���sٴU�!0޴���;9\���?�˓(�T�c.�`q�8�������̓��d�Od���O����O��D�|���0i��҃�}!0�����<k2��.Y[x��'�b���'�87=�bJS�]*���*T��P*f��Q/�� mZ���S��!8��m��<9�(�<}S��U)��i�D�0�+@�<�7e�8R���Ԉ�����O��d��G��\H�AJ�b$^�)7`��
�v���O����O~ʓ%_�&������'7�*�Z�Mx��+b�<H�׊4]��O
��'z7͓Ѧ%�H<�PܑQݪ����9h�JPX�+�F~��2rC �S�%WҘO^��IR���p;�q[��G&:l�Rg��'Q���'���'�2�i�O�D�p�h5��/s^�C��ܚ%�\�$Ӧ��@�ʟ��Iן�&��sީ㴮F�f t�hF-�%R�<��4U�V%a�
=�6s��IǟlHp�ڀ@z �X�V�I3��Y�`��3兂Z
<ec��|U�x�I�����ޟ`�	͟|��%BțCy��h�-z��[;�F�X�D���'�O@���'O �AIb� �I�Y���zk���-O <m�4�?Q�Oʧ�2�'9�e�Á��f��F��z��A����+O��[����?a�O'�D�<a�N�}]P��΋^l��EV$�?Q���?9���?ͧ��d�ŦMV����ZL��+	�[�E�q�@��才�M�����>����?Q�R)r�
�%��acN>j�:)��ͼ�MC�O�];� �R`�/����EJ%� �i{�e�'E�0XJ�3O���OB�d�OL���O��?͚�ڦ8��H�M-N,�!zTL@�x��ʟ��4dg�-O`nZ|��:|�]r�˚>y��Ջk%,��O<!�i��7=��r�	wӖ�w��@���س~ʴr �ՑTʜ���DV�˞�$N��䓐�4����O���8 ��d�ԣC�$ ��0[����O˓1���ڣ4��'H"R>e��\!@YDF�D�Vɩ�6?y�Y�ȣݴLu�vH#�?����$^�b��ՀR�KW�0U��x�n<�doQ�_T����T�R��4PA�|��	�~y,��#�?�J�s\.$���'���'����]��2شd���s1�6��#n��`YfLC�}��p�'��7�+�� ��D����c�YJF\ј�t���I�2��7��ަ�YV�����'��80��?a�UW�HAU� #�Ma�؂�4 �bl��'
��'R�'R��'L��t�`'�2R �����}��@�4/�l`C��?������<����yf��&����t���Х��%ʦ 26��Ѧ��O<�|:� ��M[�'��P�N�$�yQԂA�����<	s�Y ���B0�䓁�4����Mx���w�� k�T4jD�O�����O����Otʓ95�Fe���?��gz�Z4�S�.r
��qe!a�la��N�>Y'�i=���*�Dd0�i�B�L�X7��gG�1;����|�n8��O�c|��$?��'v�����p>|:��H�4�,��e)��c#~��I�$��Ɵ��	u�O��B�%~�  b�� nm>��E5!"
i�,$���<)0�i��O��ڷO��ң�		Q�pAyB�ծ�y�z�8mZ>�M�U��+�M�O��R�D+����bI�@-E�c���
�$�yή�O���?i��?��?Q��P����fQ�B9V����5�$�,O��m��h���	����a�s�Y�@�#��@��P�6e(š��Q��V̦�b۴9v���O��5�`W�1���ZPjT�͹7r`��g�n��i��	�B�ן��v�|�R�|0��L��`c8�Hʴl�����Ɵ�����\y�BiӴ䨱��O��7-ihx˳K�(=M1�:O��l�L�28��
�M#&�i��7�D�-H��Д�' ��3�	�6�PP*2at���N7����>e�K~2�;Z�h�k��0|X��uEN�*���?���?I���?�����O\5R�ΐ7��,�$��;T���')��'{z6Z�h�2�gt�f�|��0(�@ej�I�t!�"+Ȣ@-�'��'aJ�;iۛ�2O���&׺��&�"t5�5��ڢ �d�i��ߟBǗ|2\���I�\�����ȲGR�H�b���\#t$�q+�ş�Iby�ln�LUR1	�O��O�'}���9s�L?1r�d��Ͽz퀨�'J��Z웦��OLO�S�"�<��&�W�9��
"+2b���("�?�v�ʈsy�O%�P��*#��'��8�ő>�QRBM\h�I��'w��'�b���O��	��M���!H����l��K�Z�b'j�q����?��i��O8�'^�6�0Κak��[�T�p0hպ8N~�I����Ϧ��'ϲ]qVM��?�4^�$f'],�B�"Q!�?��1�r�̖'^�'�"�'���'��S����(iJ�j�D�y�ꁵ7K@�:ڴ+_�I)-O���<���O��mzޱ8��M4X=h���)ь]�>������O�)�&=��l��<� �݊��˻/ǘ��(�>X��m�d2O��+pLK��?�U6��<���?i�.\9��r�+�'}$��	H��?���?����������	a��^yB�'�pM+����%�U#� �8.�(y�s�^a}��'�|���:���B�� ���!��$�&!,t�b�
�FdB��X�Z��Cd����][�=a�'�%�R�/ЙV(��d�O��D�Ol��&�'�?yƅ� �4��ˉ9'�LH�m�=�?0�iPBd8�T��k�4���y"�FmAA4дN�QQ	ӓ�y��'s��'fy���i2�i�9	H�?�aT��)�[�W.W�z�6���s�hy��'�'�B�'�"䙘\�Fm�̈́)a�E��ɌTx�I'�M#'З�?����?�N~Γ�Y)u/Xl}��gYR�[�P�x�	֟`%������!�J�^<��q�T4F�0M��V�hĬ��%�<�4M_����������d�z�\1b�Aן._֩1�惞q���d�O�$�OP�4�˓B"��Ö�S��ړ"�T1�[�29d���E�G?bow�|�xS-Of���O�7�؟3�c���r^H�@P�q|D�z�h���	̟8K���3>�dQy��O�'�,MM����	̃H�d�C���y��'���'�R�'g����{�*�Ů��cv�MPՀ��<U��d�O��֦Q���
syRbc��O�쫒̀��x�ZW�KH�p {.�~�I�M���:�k���M��O��{�m�0o���5�.{��(@m�<I$��[��Z�ܓO�ʓ�?���?���th�3�ǤP^����N�)u�� ���?A,O\]n�y�µ�	�D�Iz�#->۾<� ����E�d-���DKv}b�'���|ʟ����c��h-{�)���iҭ^=���"FƲB���|J�c�O�J>��.o�$�&'
�_ё�-B�?����?���?�|�/Ob�n�?�E��J�,/x�yT�
�tP"g*[՟��I�M����>��.��)���أN��m)��8q������?����M��O��ӣD���� 8���J�Di�pi �{W�Չ�v#��<A��?����?a���?)��-��K�W8����)
�(�C���Цr�/�����I�$�W��'��7=�Nxp���&��	��O1���D$���'�ɧ���'�B*cs�f?O� "`DG|ܴuن+CY�N�:4Op�ō��?�%�-�Ĺ<y��?��oхn&�8	�BӬ$8~,�@E��?a���?�����ۦ���Lߟ�	۟h�'П\n\��v%�m��[0��g��g������ID�	-Xx)za�GJc��B&C;n��r��̓~v&$�K~��B�O2$����V��S��d8X��#�S���<���?����?����h�H����~(yJv��f۔����16������e��I�SyB�oӠ��]8sd���@��a~E��o��`Ʈ�����ԟ��SK�ڦ��u'j��a���&Il�(\Гk�.�>9&��a���$��'5b�'�"�'ZB�' <MÒ���{����D���
n�2T����48�xQP���?!�����<�k�/XW4��wK�"M@=(Ĭ+u��	ן���a�)�Ӣ)uX�DƘl�S���	�쑡�O�1K��'.&سG���a$�|W�t�T��$���Β�a��U�� ������Ο��	ڟ�uy�gq�pT����OL�p�<	��q�� H���9O��o�w�0��ɏ�M{��i"6�.����Ub�1��O��y,�EI�~�������󑆅�8�$[gy��O��D]�Y���RD�*�B��REC&�y��'�b�'�'���)Ƌ_2zI�&�ƻ|X(��D�>�f���Ov�d�٦)��\Ly��Ӡ�Oz��q(�!|n�m��Ro����X��-�Mˣ������B�v���C�P�{���fW�&e��Y�O� ���b�ǧF�A�R��d�xc�7<R�����!�Ӈ-�r�#����E�:��oC�uD8x�_�q�N�8�.�<!���tǋ�=|x�	�\�lԚ �#늳PB�$IJ<9�F�?�L��Ƞw��c�8sh�ҳ*Ԫ%Z�<�L�8"��pD*3�z���$�(g֘�+b��>[8tʥ
�� ��hs���1T�]�̩j�8x��H�))0 Y� ��>I��
&����2B��=35�ǣ~�h�UoA�'�HiB6�f�# $�<g�V$��l�+� ����<>�`B���¦]��۟$�I�?IP�]��9���x)t����ē���F(��'8�Dv��p�jX`��Z�&i�yl�Ty2��2En6-�G���'��d� ?)�/�AD̹����`����a�'�$舏��)ڮh�ȵy��+M�Ű�nF� 6HV7��O.��O��	j����Ы��\C��$+gCB�I8`���M+���W����D�!2X�!��,X�M�� �z���i��'�O�^$O��$�On�ɢ�uQAڰ(EDqk���Zeҋ}� ]�'k2�'����Xt���h�Z�K��Y�O��6��O0�cm�K�I֟`��F�i��(���5�*�cԢ�/�(��C̩>�D��l̓�?A���?�.O�ժ�C >�`�K�d��R���Yݖl�` �Iן�$�(�'�:�J�^L�2)��۞Pj��'@S���'N�'��\�@;dȞ���d��B=�1��ùhL�Фg����O����O����D����S�>�2P�'�/@�1:��%&�t꓾?����?�-O�1q�Us�S��n���.I����-�p+�4�?�K>�.OH08���L�a��+�;4�N ����sf��'��V��� Ɋ�ħ�y��q�� �}pW�RV�|� �]�Jm�����xQ�x9V�.�S��JT�~���H�W򭘲@��MC+O�`0�OԦ鹭�N�矴L�'>�i�!�%k��a#%��#Bz�4��Dژ�b?=���'��6.��1ֆ���JrӶm�U���]��������?�cN<i���굉��+-�U(���p)�L+��i�6,)�����PJ[J�BH��Y�8�`�#d۬�M����?��^3�h�C�x�'<��O���A�M�(����-]H�H����(Q1O����Or�D��`�|��DC<P�qN�4)Z��n��H(3����d�<�������Ъ�z
T��%�6#Ò�¤�f}�׆u�'b�'H�\���q̕�L`��:gw"h�Յ��^�ҬO�˓�?�L>���?1�cY7�@Ș�)50�>�3@��F\�H>9���?����䄖�}̧
h d/Yy�8���@;|�lZCy��'%�'0��'�6��d�'e4|�@��^y|}�+�,m��a�+�>I��?�����$�9a��O�R�̵Y��t�EaҮvj�y��?e*�7��On�OV���OT�c�,-r����0���HԢ���#'|7��O&���<9r�97��S��@���?�҇�G��M���K/gB��%�����?���7� ���џ�P m@�f��sK���9��i�	w�b`+�4�?y��?�'��i���6���hZ�dy��,��쀗.sӤ�d�OnuɁd4��N�'y����w`�>h�B��5f��z@B�i��2��>���O��������'*�I���+7�B�SzHX�$� ��$�ܴC���Ћ��)�O��C%����B@�&���)@%Y̦�����P�I�@���O��?�'}*�a��>5��ж�G��Ժ�}�� 5��'b�'�"��/q�z VF^!5��MqCl ��&6�Oj��F�q}2X���IR�i��+Э�.J��P��@%� ��>YN����?���?!)O�RP,O��{1�1��=�tiȄ'�b��'���H&����������^��z��]�t��$  	�L��qy��'��'��	� ���O�P�i7�ùOؼ!�ej�:�E��4��$�OR�O���O�Q�����0�g�'w��,�#�2_��M��>y���?-�M{-O^p�Gq���'z�]{k�D��y.�o���Kr�t�`��$���Ob�$]�z�㞈ppKX>	R�!
gb
�`��,���s�R���ONʓB�<����'��\c��0�É�ƍ���:3L<+O��$�O����*@Abǀ%{(z���ʏ'tQ��iI��r|#�4<^������S����G�>�k'�?U1�鰃!o���P����֟�{M|JM~nZň�K0m��P�JG��e>&7�K^8�n�����	ϟ�����|:FlW�{Iڃ���$�9g�/ar�F�'U��'ɧ�9O���U�e"`����P�����A���m���ܟpz�lP.���|���~R��CG�2feX�,
�Zfl�+�M����Ab�3?i���~2G#V�
噇l'���su��M#�'z
)�)O\�O8�O���_�v��c�\;0<p2CC�X�		��c�4��My��'��aYp,�,�f�ذ�_�(�zUJ��Iܟ��	U��?��'t�!��-��'�6��Ǣ�w�
�jڴ{�J�<9�����O�9EH�?5����F5��ܐ"樅 �i� ���O��t�	py�l�<�Ms�
�X�0��G�2s�]��n�Y�	ޟ��'��'>#�S��<�ЈĆhsU�A�av:0g��Mӊ��'[���O�\��lZ-��4�T��K,�e�V�i	2�'��	d7,�JN|����1'��D�U"��?�1!�,�r`$�4�'-lԒd�'�O:�)Ǌ#��`��޴hy���
2�fT�����C+�M3qP?]���?i�OY��Ԋ�Lk�� H��\+��i!�;9�^��	:��'���-�I)E">��M�Y�&4�h��UJ�h�u�I�����?��L<�'1H�:4�Ю;�ls1E�*5�`)b1�iH�8��'�V�&?�k�0��H5'��q��a��� �i3B�'��F`�)L���FS(>����4bRDA�oQ>��''R���.�I�O
���O�hz��]�B����/�!X��q8��J��I�s��E+L<�'�?�����]5n/�"�Y�}���Aր��,o�㟠���|�����'��ޟ4[Ah�M6($R�W��Z`C�Y�T���B���+�	�t�	�NxĴ1&"�
<��d�5,Ekt�As��|b����qy��'5��Xݟ<0�ը�		����*ʂg��eh"�i���'��O:���O<��`EV�p�����-{P�h���B�ҝ��b�����O��O��J��XvX?	�I�-��t��Х|�>�p#���Q* ;�4�?!,O,�$�O���ŻK�i>7��?E|�;B�_v0y�Cä{�f�'�Q���Sퟘ��i�O����4�1�E L��p�5$�(f	B}��'2�'�*���'M�s����Tk���qO�	6�%�W�T�<�lZvy����	z6��O��d�O��IPA}Zw�ЦA�82<��F�k��T��4�?9��Cz�a�(4�s���}���~%Z��%X�n�����˦�ȕ��;�MS��?9�����Z�ܖ'��� ��1�/E�R�>�)��� Z�hu�i�2l��'l������P��`�`�ϖ`ބ��`H	8��5(2�i.��'\�
�:�����$�O\��?E}8�K��ȥJ�4�R#	�p�$6��O��$�O��=O��������ᴉ��/N ��H���)�edD)�M��(/�iGP���'1�_���i�b��ߐCL�s��݆U�h-�v�>"���<����?��?A����d�"c-�1rG�Ng�xJ6��,f��8�b�c}B[�$�	ByR�'���''��I�NU �T�z�N��ild�i��E��y��'�R�'���'��	�cgXa�O^t�#��j��K�=o�hٴ���OD��?i��?�2�Ue}rhV�$���a����hcH��M���?����?+O���ύD���'��Բ4$��Rq�_�#$
,�"�h�d��<)���?��e�PD�|nZ*"Ԝ0X0L�.��!�߫-�|6��O��D�<��UM����|�I�?s��J�nh���w����G�P���d�O����O�%;�1O0��<Q�O�
<ф�͕V�=�E!�miތ��4���I�
�Zeo����՟X�S�����["n�7l7@ɓY�z1K\��MS���?Q'���<QV?�Idܧ`��@�2��r3�G Gi��Ikӂ��"�U����	ӟd�I�?YѮO��$�́$%χeO>5��B�M{��*e�iָMB�'z�Y�L����PR�H�#g21��,zA���`J��ie��'.N̚L������OD�I#K���B�%���'F��6�)�dXu��?���������~5ЀmI�XG��Xc�GJ���4�?�E��bh��|y��'�����֘.wЍ����@�O�"��7m�O����2O���O\���O���<y���a!vT����iE����S�,��!R�h�'��R�l��ϟ�	;L谌eI��XXTRC]$��Kb���'2�'��W� z�g���24�.��w��K��5Z�ɭ�M.O�ĳ<	���?�~�̓ah�\8��\k�yw�Y j�����W�������Igy�<#�'�?1�P�t�PT�g�`ȶ�#o�V�'��	���	ٟD�� `�|��MK͆�J�$/�/#�x��C
ئ��	ɟ��'����&��On�Ʉ�)X�A��pD�cŜv�0%�������Q�"l��%�d�'��|�1Ҭ-�=�5�N�b�`moZ[yL>Y�7��v�D�'��$�0?��Ҟ;Ia
S�E"|R��Kɦ]���Xk�n�p%���}z��I��2��ΐ�����]Φ!�s	��M����?y���$�Z��I*�R�=�5͑�X� Ql�)���Iu�A���?�Rf�&Fʔ�����~kd��D�R�	�&�'���'@�d�N"�Iȟ���۬h��A;��+��%b���o�T��1R��O|���?9��+� Xä��4�>�B OV-�� g�i�^��c�D�Ix�i�5��͐;���&�2+��»>QЂ���?I)O��D�O ��<���~��
f+��+ؼ���/�$gP$*��x��'QB�|��'PbLK�P�z�)�	=4��%��g��(���'��	������l�'��s&'l>��.�d
 �"�n�y��2O�>y��?YO>q���?��(��?i'�wZ�aPD��H�<� �3(��D��򟼔'�Z���'2�)���̢�k�( � xs��	y��o�ß(&����ßlXfet�X�O���a��"��:L]<b<!��i#B�'��I=C'Px+N|���2alܴ7-��QT���J����#9҉':��'sR�r��'�1O��̋�$�ɴ�E�N�ԲV��&�Q�H����M� \?a���?!*�O�T`@m@ UŖeQ��S_@a�ѹi��'
bܚr�';�'+q���g��P����wGN�.^��	�i�Y�f}Ӯ���O��d�(��']�?T���H��m��7$���4t̓�?�.OH�?a�������8D}�����]�D���4�?Y��?�$�(��	xy"�'��	zr�`Ӈ�2^`�P3�gθT���'n�I;x�)*��?q��z�ai���#I�$=�7%�6���袸il���$'�ꓪ�d�O ��?��R��t�e �
&oD ٳ����i�'�t�'���'F��'
�X�C�͟d��8y�AH�Mu���!����R�O�ʓ�?�,O����O@���C�X+��s�L r�♣.�N���6O����O6���O��Ľ<Ѱ���'k�2P�`�:!�Ǚ)t�	�J�$7h��Z����|y��'&2�'! �y�'�޹�G��"9�}&� t7�X�Ѡ�>q���?�����A?���OR�W"<��,"W��M�n�2x�>7�O���?q���?�1��<IO�<�gF�o��P�4DޑO;�H��uӜ�d�O�ʓeU��sS?%��Ο�����"�V {`2��ل5B�s�O �$�O$�D2��0��?�{��J*Uqr6F�2�Δ0��l���qg�EC�i�"�'��O���Ӻ;@�U�����n��n��#�Uߦ����hȥn����Ny��º*�H���*1�H ���+CΛfmݼ�Z7M�O��d�O����k���\��a�L��PA7�G+l���	]��yݴ��m����Ϙ'}$	&ey�g�8j4�=kaiL (ؐ7-�O��d�Oܱ1E�O����D���S�C	0�b�rS"'6��@𔊝��'$�i�ge"�	�Ov�$�O~H�F�b:�pz���Y[ܑW����m��:(�P�M<����?!N>�q�? yP��>?���y�)�di�5�V^��c��%�	ϟ��	ɟ$�')+TdɴcV���7��=�x��+1B��O�d�OZ�O �D�O4̺"ۚ>t�)�+��+���D�B+qO���1D�.�:"~JT�?i��3!�P����$�i�<q�;���1��5�����aXk�p�LQ�`lU:\�h�i'��I׊�TN��n�c��?9C�丵��%3�l���cJE?XI3s�J�UǤ,�#N�HS~���)+RD�6��?��H tdEqW��r�ǼYڵy�� F���'$��E�|����fp´�B'U���F��68Y�.	6r�����L�`�<�Γi��1祝�3��x�h	�%?�]�	˟��o@��h����^��	!�%�2��)�|�@֚$Bep�\�
S2�(6GUv�ĕ�|x�ˠ��"Jq�E[s�d�EZ�,��Ä_�FI` cӂ(���qHO8��R&|�	ҟ�D���')��"᧓&m�0|P"_97��ك�'eNY ���.ezt�	�f�$1}����@���p��dǫPlj��7h��\~fq{�.�7����O8�	;4�������OB�d�O��4�2nϵ��h1�Q�
�f�E�#;�4�"�O��Y��8�1��'��b��Ŗ&�
ӹ!�6ii1�skɀ��'��hD�FC�g��}�N���a���V�C;,t��e~����?�'�hO��3��PJ�~�H�5k�Ԡ2"O*�0�kV�.d�(A�J�C���x䙟�����?5�'�(�$��	�T<Zn�0=�ج�� Q-h0���p�'���'�gݙ���(ϧl�H��m�]�]ꧏ�U��xsD�L����l�<N�:�h�1�1#ǊO.i���r'2q�aPIJ�E¸X����b��F����vOJ������ j��&���|�	W�'_�O$|���S	^!A�$,^���"O��wܴI(<��^�P�\��r��o}�\�|�JH����OHh ��A4|��0D�D2���Ⴉ�O<�$�=�j���O��S�Ku@M�@l�"�(a�iBߦe�)X�Xy�N?$aȶg>O�ܠ���*�\�`�疆y��6mH6jAz$I��@q��E�u��xr����?����ߏl��aA�� 2�Ƭz��#�1O���D��= �D;&K�Fd��bF8�!�MӦu�d�O�e:U+H	!�,��`�(�'�`��Qh`Ӹ���O�˧O����bǠ2u��MlU`R��!�@��?Y����h)��^�x�r$�)q���P�T&���5��B �k"½
����f���NN4(� � 0��z;�f9f�,�x$���^6��Xfmfa`�'�nDK��?1��?�������glBa�"��e��ߘ'���'�(d#�����X;��<�t���	9����FK�Y؂bD�ML,�����M���?���&P�ȓ�?����?Q�Ӽ�cˇ=��jEOO�~��#�Q�'��}x�$H�����t�0L�n�U|^�ۧnN�>ʪ�2$�|�k������}&�ty�bQ=d
���� �9!��[Ο���lQ`Ο�>��?q&�/4�){"AU$F��A����(��xIK�t��(�#�/6��YA�ޑ���z���ɱ<�@�7Z5
�2IY|_���$B�Y�<� @W�j2���	]H�P��o�|�<Y����LG m�U!��<�^|��x�<1���/+𴈂(�.- t� ��r�<��"�����aΩ��X�+[l�<�EbX9o��qr�)��h�@��<鳬����@�#��%��j��]�<�fE�bN��d�<A`���Ly�<i'�?:�9��*لR6�X�su�<��eơ7��rA�tF�xV�[�<$e�
lD�p� FH6J��TŁT�<�7�V�|dx5( �~�*]���EV�<A4h;tM6�iT�ϕh=��@�G�l�<1�G�o�ք�u�В,���Dh�<I���c��x��U�K:N�j�N�<!'��BRV��"(ёEa����/�J�<�u@S�s���9! ���˔�KC�<�ca�JpX1uMɨ\Oj+w��B�<��j"1��#�Bߍ}�$�����<q ����Þ�7� % q�<�Wj��5�\����t�4��W �n�<a$O'>���3A�Z�� �BdPj�<ASa��p�veH�i��N��C@d�<� tz��,MV2-xE��_��x��"O�`QWJ�E��L�'���@�6U T"O�����U�>hZ%��<N�����"O|��q�ڼic$l�.^�wC�l""OZ-�����,��x�"Ҫp6r�U"O�a!�%�$h��h���-V����"O2���ֳ`ڊ\��E�Z@���#"Od��wLH�hE����A%w���1D"Ov��ڑV����0-�|���c"O~@�p*��&H���С���N!���
6���*E�\"��e	�48���:3ɰ�0��N�u�
��D·�yB�8@�,t��瑚u\�l	����y(�[�9p��	f-$=�C�K��ybIv�)���%Vsf�&芤�y�햳,�N<hƌ
�TD[�ꅚ�yB�G,h���Y�K]�FLd�[��yRը�%�d®C�B�����y"k��(�����h�'fƾ������yr��$4��CͰK}�1C�M��yҍ�{����T�̊KF�13���yr�Ĳ|p����?nP�����y���RӐ�r����F���<�y��s�Vm)���}��1Xb�.D�l{|%xq�C^���]'�y�iV>tЫ3&S0J'�`C�J��y��O=F�X��	�:NQ@�#���y�ÀI�DD�d�M��AB�!U��y��x�x�{��ϽR�m��N�8�yB��!^�P	��vZ�Р�i��y�.P%af2�+ �_�x((��yBeʂx��*B@V&
�/��y�ʕ�1<b��r��0c��$�j#�yBj�  ���U����L��͗�y�;ɜY1jȒԦ�-4�މ��m��f�90�EhǬ�&a���2���r�4z�48����\'ta�ȓsV�}@��ɀg�~�C%�G*,�����T�)p
#��uSc��JՀI��njC�Ǚ"��1��\-H���lH�j��\�� ʱ���ȓe|�!���S�9@v�O��t�ȓ	�f�1��ޒ"��:���h`h��ȓD�t49�I�y�0�1ҎJ�[^`=���E�C�ΈZ+�� Ș�c=�P�ȓ[������6�rL;�HړH��܇�	 mG2y��'H�a[���_�V�R���P DC�'�� ��i�R&�!��(uB��L�,�Q���m�V.?13�.,L��f#?�81A��@ �v�S�O�z�!@*��$#�� �%����i$�V����{���'fl\�����~D���dŀ`\�L�$c�D�H؞�Y3H?.jP�bǌ7<F�p��O���	)f�O뎆���	�_]ƌm5z��� ��K) �$�i�ʝ/�0����9V�AΓr�΅��.�"W	P���鄟=�}�'�L E�>1�.������*U-�H!�n~I�bg�-|�r��d�/x�b�I1Dh�RN�>?�D$ B64Sh�ɔvj�#<E�d�ٓ@�2����a`9h�CԵ�hOn91v$1�Yk�A���8f�8�)ԋTA��L���&�"��3��4�]�J�����*v&��?E�4
�7Eȳ��_-pQ�qӃ"8!�ҬXȭRF�0&���$.�!�Đ44jHZ�?>{�P�0��6!�dưl�r䓑B�Nf� �@�Pv,�&��$ʁ$���,b>c��0Be3?LL�sG	3�X 3g�#��p�e>� ��[Åب�Y��"�,0�3�Oٻ1T����'FN���)�t%-+ �
%�a��Kyl�khXoHp�'��%�?h"�����'8U��'|� )%�P3S%ޭ.�MN�0��OZ�-\���!6�Ol���Դ)�r��53���E"O�z��4���;�L�L��ph$���3���*3�f�PH?�3�I�1��3�߶!��As��W>|I�C�I�5��C��&A��`�n�=~�R��5|�LRT�1�O8�q���,�dYW��<��5��'El� �$ʸVW���O����2^�<��Ft�8l��"O�����aR��5@�z�j-�ј��0k� �>���0���y���e���a6OX�c�X,�w"O ��`��#GL8�FN��k����:.��2Eߜ�	�!;�3手c��c���	.�q�����#�|C���g�E	��63�@���"d�d�)�X�t��@sc/!�OP�q�F[����J�`��}	��'Ҳ� ��]�%��OHe�G$��5ј�QAL7���)�"O�9p"��X��j�F��z���U��2=(jհU� ��T��
-7H�F=cR ��"O<Hj�c�tp`�z��_�U�J�"O�"ѡ�����C�c��>��d"O��K��F�H�r�9��\d(�[e"O.8���ݼQexբ5!�?K��"OR�7��V:�x�O�G\��;�"Oi `�Ql<!Ѩ_�'F��"O���'A�'T�����A�`b"O���A�JH�hF��w"O<���1^k�X �����9B "O&�$O�SN��34�	=P��%�v"O�}Z�mH(g �A�E�/���p��'��C�M�8o�	��2p���<|�2���/!�B�I&"cp��b� ���<��L�*��eb��
*��
���1K�5���MF�$U�#�O$�t����P����Ն��s�P6d"5!G�}����SiZ�x��y`�L2����g������|��8O($�~&���a��u�\:�`ƷG-���L#�ɡI�+&A
	K<����I�0M�dx��-Y���`���d��� E�|��ѐ	���=���2�XZ#m
�7%�ᡢ"�5�|cg鎧1ڦpy�Bܦ�z f�k��S)=�����b�ʵ��J%
�s%��=KԈ$�� �:p�t$�if�X�B,Aeڑ2$z�>m!��hl�,��
'bp�������O�o$��'>z���܂~!��x�Pu���ږQ�8X��J ?Ֆh@��p���.D��,Ԉ�.]�]�6���OF�3j�2�>�rT�vB:e�V�isV�$	�'j`��FX�,XJ�04oŬ�HOt��DE��1!.r�"�0��!R@
�ԩ�� +r����:f�랟o�/<0T0��ZQ\��'͔u��L����)R�%��q��M[�?\Oje1��!�}SbdH� �J��	�(&� <0d��<)Sgk��̈��'@F0��pW���c�:�^��b޻XH����>\�br6[p���F�E�k�������7cԴh�!��_���Ѧ͍=?��{5JU���dޘ-����O�|ʢ��	osƵj�wHL��W�X�^���[�_X�Z���O��#3,�H0�����pu
��C86�2���Oj�pŬ�(3*i7Uk���2NOw���0�J���$� b_#`��sà�H�Q��A��Th���Հ�' ��@�1`=T�NC��ߊ��}B�i6�	:T���i���l#0�Y2��O`Q�Y#��q�A$N�h!�%�1ea�t2���p=��DH:pm�\2A!�)B�hj��$@J�)AW���H�A[;X|�S�K����~R����p��q�nX�����ܠ/z�)Ó�hQ�F�^�d|�� _�����4�C.�Ȅ���Ó[	|�QA�o���c��<�cBEW���Ur�����F"�TESu�ÐN9���N����+`�ؗU.
���>���G�k#\8ET V�H��h��>�l��R�X`�I˨9(ڹ�f�b6|Ճ!�\�:�4������f��#b�GX�Ȥ��EӘY�Z�FyR��^��M� �6(�>�McG
�V�r�k��eK�C��[}�U�@h�-Z�T��Q�mQ�(�F����
SxA31�_<YD��g�?X�a{�� [0������o@?z�|��}�Ǉ��O��C�@�0���=@������<3����Ta� ��/�<����-�V&
�����zU�Ti�D�t���چ����S-Y�F�ԡJ��-ؾ���i�f!)�LVHଣ�#�
�|�n,��[C)WU�P�r'��d%��Gx���;I��`Cŭ �2��r��#�y"��/�dA��lV� ���R�4�X��E\Of�
�{*�Z�+��J#(��N�7�L�T��tv�+b�p�!�D�7w� �ah�1u
 C���   �}����8��_�A�@��@%S,!�3�F1o�X���(n��%B�d���ɘT�Bu��7h�,!�]�w�,��e���#<���p�ܦJ��I$�9D�p
�S.F��D�G	h���I3?���,R��a��E�A�x���'ʧ1;���S��;�T�`���[.���#�&��B3@ �6В3��1c=h�+0�)C ,;�hy�g�(Dt���@4n�q��kS+`�J���h�u�w�!��u�=l]tU�Wb�>��!F�1�`���M'\O����@R�x��A=�����'�X�p��o���pL�@P�x�'L�YtHe`��ęiTD��C��y���A����ׯQ0 ���@!]���I� ��8�R�D�T��3��r�O��x���Y��]�W)5��%	�'E �CBW�Sx�ٷ X�?��r�'_��r�A� �)"Hǜa���S�'�$q3q��WPr�ױT_F��'D]2�i�p����6L� |�
�'*�y��	(vc��t����	�'< 9լv��I�g*��,�	�'Ӵ ��� h�ȕ��0K�
HZ	�'�� S��^;mȐ�(�!C)̼��'t,
VO]�Z�֩�eF��3�@b�'��R�,J.0���KtF��0�H���'	�t:3*��L vm �,�� ވ�#�'<H�q	ͤVB�k��̦i} z�'���`���ZH1P�B,^� ��'�����!�"H:�0��Z����'x�	�TJL-#�ZI���OZL0��'��)�t� k1:كM�|�'�� ���Q���5*1��)tHZ9�	�'�&��B�ĒtDڸ	aJ�` �Ѩ�'�� j��nP`<0��U�<�'��!R�
��gq^3���?L3��J�'�6z���X�N
dCۅEƺ��'���Ѣһ^�hѢ��	E*���'�Rd��S�"��mа�F4.]@�
�'S���a�v�>(��n�<z�
�'02���/Z�> V���]� �T���'l�����C�K`�H9��
���DB�'M�aXf��~H"`�Q�z�FDR�'F���
��ڄ����l����'&`݋�@�.@�`9��6<�V\R�'���3C@:,�1#��|;2)��'7�a U�H��I�T�t�����'r$�똇W�轸�A �[��x
�'��,�D(�F�r`���XM��T�	�'C�EXb�&<?N��wꃾH�����'C���vˀ$V<xTB6�g���'0t(#�m+1겴ҵf׈0�:�	�':|sc�|���ĉC#�
d�	�'����V�̴%��ҵ��G��y`�'fL�6OZ,H�1�d�E@$$��'$J��2��)k�����;�JQ��'�6�볌�w,���@P�%�""�';�T#oW�V%�Gc�Ɩ�S�'�R��ǆ��f���X�E9~�D�z�' ^X�Or	��#���*<��Z�'��(�fC*@F����Q� ����'��|����	F��D�mֺP���	�'`�[�j��Hߕ|�&���'�"�4�ܖ~��X5��4%ǐ�(	�'�R8{�g�q��9a�Bޡf�T��'�؁�!n#�l �P T"sL��z�'��ت�(�v��J�O�q��� �'1���ɏ~�ع��4c|�ɢ��� �%q�E�7��|��d�9yä�b"OPM����2,r�SD���U�- "O`���Qy����pQ�4��"O� b��o��҂��t+\aab"ONa������pk$,C$F�۔"O���
Ęo{�Ѫ����2t��"O|E�}�|���Ԟ�(PѰ"O.�e�-OG�}P�GL�B̭��"Oh��ZD�� �e�-|����"O��J�_C�d�de�Y� C"O��Z��`�h��b�9 F@��"O�ƀ�	1��@䐉�Nܠ�"O�y�&V1O�"b���z}��W"O�Ђb�=~D�A�a�\{j��"O.EJ��&+��]��ʆ�\,xP�"O��D,Y�[$ ��dT6�0�"O���g,�*И@�B�E8��R�"O,d2��0���p�NS$n #s"Ofiy�J�9u�HP��_�wԜ�F"O��ha�Z&o5�@ȗ厅��4�"O:����sa$u�T�F;a�08S4"O�m���Γ*f�!���B/� �I�"O�m;5,Y ~~�"���f�̹��"OL��5a��
���2���x���""OȨi��3	�x��7��Co���"Of aV-��E�T��Nγw��B�"O�E�#�k�Pd��[0n%`""O�x�%B�
0:~A��C�'R�)"OBl�WL�j�
�3S �89���"O�3�N7(6�MB�n�3Ь٧"O�`��+?�Б���ԙ~�*��"O�l�&dߚ-	�MhBY:
l*m'"O�c��	yhQ�DG�}��|��"Onq�H�Pƞt����'ba��"OJ���o晙�#�"U�G"O���åаM�Y�qH��@�r�۴"O$LY@�C8~W���ǌ%�ΰ� "O���T��7�����Gg�$��"O�Ѐ��Gg�y�(��`�4�B�"O�����B&�8�V��v_)��"O~9��T>8P-pQ̉�LZ�i�"O���vfk�������q���1g"O�˟0U�����i
�!��%3�"O^t)��O��i1&h�p���p�"O`� aM"2 �	���·|�Ј�%"Ot���L���{2�ώf��)Y&"O�A��N�(R�CсE�l���B�"O����X�.�p���`T�[|�I�V"O�4K���Q�ހS` Ϛ|nP"O��[ѯ]?O?�m[�Pv�d8�0"O�LZ5��Z|[ *C�Qeک�!"O��X�iX1O^"X@�Gɳ`���"O8�!��� g�� �V8Аih "O�x��.}ѠT�C�e��4G"O�,rb�-�p(CԀ��_d�81�"O�4kŨ�,��C��@�\���t"OhycQ�Q�hF�:à �@Kv|�C"O�la�?_��b�oU�1�M��"O���gNE=o���"�N�/N�	P�"O�|Ke̬y�@���	=E�"Ol(2+P�̎�8G,ӟ#8 -�""Op�a�$@�P�Ӭ�h�2�'"O���C�1S��}�� �s�i� "O��ie�?XL�SK(=�Z���"O� T��������͜bM�9E"O���S�W�YDf�OI.L@F"O<�2��g�,��&ŃB��s�"O ���(�;?����E�J�eI�"O�Qy���b) U��)��h�"O(��q�o~�	Zv��>%�T��Q"O�$▁�Cg8�E)  {�b4�"O��s".u8�9��2�� �"O6�P���4�!x�ɛ�*�,�D"O�,i#-�0jȂ�IR��A�D��f"O��
�òz��h�e��mj� ��"O��E^���{���.R��b""O����n̕N�D�A�/	>#nJ	`�"O��`�?\���%�ٺd�����"O"d�##�/X��e��  G{�sq"OB�0D�sةS�K�Oh0h:�"Or]����:jFLbD̙��v���"O�)�d[�E&��yU�?�r�cD"O��J��= ���6	��`��F"O�ѱ2셑_\@a˓)�H]BDx3"OҘW)��,�L�Ն�J�pd��"O�����ç�������P2�=X5"OLz�,D7	c�H�$l&�h�"O���W�=F}{&��΅�w"O�%a%1�����	g�p��"O��S(������M�`K��av"Ot��K�]и�&63MN-��"O��3b֥%��q�Ď#1B��"O��i��B! �2���$*`����O�=E��X#/ψ�J5f��jЉW�S8�y��_��\"	�?*�	��yR�R�CL��jƺ۵A�
�y�"�0v�6 ���q����5D���y�%-�20�paJ� ��COS�y-V�#�403�\�mn�����yrE�v���z�kX#���h%��)�y"��wl�PW��2S��c]9�y�+ESK"x��
�1�����y�`�&�"���F1&ZFd�m(�y�\�`OJ�@b-x&�yL� �yr�ͽw�Ȭ�!���o�������y�+ CwdC7�epb���0>�L>�3b	�*IF�(��F����KG`�<���-�"LQѳBy�sD��Z2�C�	�EQ ��ClWB@����>�C�ɷ%�>h��f/ro��a�*�+L��C�	�Hں�`ă�`ºq��4(�JB�`Α����,L=DuB�96�B�I+3\*�$hR,��E��7հB䉲�<��#C����v#��<[�B��%4���O�R��)��-JcJC�6j]�=��<)����%2�C�����#f+I�X{���
a�B�I؟@�oÔ6J K�F������(D�h1�ʊ�>p8�퀙I�~��A�$D���*D4vv(�a�^�&P�3�I$D��R��׹t[�epC&�/ z��V6D�볪P/1FA�@� �O^d0�4�5D�p�t/L�F�^�B���F8�5�4D��F��=Cp^���b�f�T�M2D��Ғ�[xt�v(��RY�T�k�.B�	D��Eq�A�z�d����aʌB�	) tD%p��q]T��F�� @XB�I?���C�\CxP�'��p�C�)� ���O��7z�iQ�MӬZ@�b�"On�`����|�)�+ǦB�ՠq"O�hrP��r�Q�
ĳ��b�"O�!�.Z�8u��C���b�B�[�"O��Y��T�zBd��E'd���"O<:w식��8�W4I��
O�7-� 9��|����q�jp�'	
�!�d7LM$�� ES���.�h�w"Oʩ�7`�c���F�3!MH�"O>͈����
v��r��Q,KƳiLў"~n�����t@�5B�a��=f@`B�	��6"s#�2c1�!��8� B�I�v-�`ѕ _�?h��[,w B�IN�tl0�.�:MQ��GD�۠B�	0L�,)Z!�U-�����@��hB�	8�j˳�J����{"��<y�\B�IuU�|K` �*'�A��)['E&B�ɻ`tL�P���e��J1n��w��C�ɗ|�tu����[T�b��s�C�	/0��ڧcE�ww(q�Ƥ�+?MHC�	�1�8�J'�J�j`<E�#�'jC�I�z�rY
A	M�~vĸ��[b9�B�I�>?�1G��$�&yP��W��|B䉔`��aR��9f�2�á�I4C�I >$<AH���s���,WmDB��^����G   T�X�jH�,f B��5/V�0V��}:�0Cn�:��C�	���r��E`D�C��ER��C�	&_4ƹ R�˖�,�Qu�B�	3XUB�І�ӸQi�@�F�(1�B�	1.��34%R)z��(Я�6��B�	>Ob�c�s��8��.U�hB䉄G��Sn��wܱ"�K�4,C�	
�&��ɋ=tIh[s��=�B�	�1 Q:����p��e�$Ͻj[�B�	 uJ�d:��\!���Q2E�
J\B䉽pӸ0!@�L�d���p"�Z�T��B��r=�dꞶ �n�Sf#�3�|B�	�a��8��I��J�dİE�5;yZB�I�_��T���'��臮�<:�B�	+0"2�ۃK@�Q����3Ԕm��B䉢�$����[+`�š^��jB䉫8|!1�I_x=�y�o���C�I�~P6�ks�Ru���i9�C�	�#xY��a��]BwCY![����"S���Q(J&T�8��o���<	�ȓl@��z�$ԝ"�lQG M�%�ȓX��)�իĀ!�X��Ո �Z~r �ȓ+������
5V������ YH4��*nN��"�<׼=zu �\���W�q3/\�w�t����?r�V��ȓ����Bos��̳o�*ˮ��ȓyb�h;ĄQ���@�Є^�M���ȓ�҈`���9c"�����Sx���ux�"A�E�\"t�Iւ1�ȓF��-؃���P�S��?6��h���S5F��>��
��Իh9J���{�B���؃<�� �,� �V��ȓ1�41��َ&j5Q���/�HA�ȓZ�A�FݧJ}�b��"�����+���Bճ)G� �7�X���U�ȓq�X5p��B>L��$�e?H4�ȓzw�SKӟ^ު��B���)����`^f���G[���vꎋL�^���S�? �4��,�b���Fj� �~��"O��s -'^sĐC�B:t@�;"O�Pk���i��$
ʂ�~�I�"O�9[v�_'fY�&cA>�`�r�"OFx����t�29#qB��U����"OҀ��ݷg9rh!�!ү?whm��"O(��b# )8�P�J�vqġ �"O���	�rԲ1k���-|�^�`�"O�X@fH_/`�V��&����Eʶ"O&�f�I�P b ����GP腢�"O��XG�ѪPdƍ[���q:���"ONEb��Xn�:����)sQ�|�"O��[�'�On��`�� 6~���"O�	���;-�|��c�U��Q��'�����N]�}B^���g}��9�'��`�O��N�6EXQ/�,$m�,��'{�H��õs)jdS�a� l�B}R�'�S��[,hP3R��
k��
�'<,���	��P�a�Ah��p�	�'��˥��*�z��!��RTp(��'{\��P��1&��1Q&Ɣ����'`Z��b��O�`ً��˧��X�	�'�(��@$��_�l{��Ks/S	�'���3&釿ӒP�eC��}�����'J�H��Ѕ	���[Y�n�B��'Y�� βt�;r�[p]����'̬�� ��4�DBKf�|(��'td��BX�g�,�S!ָ_���' �Y#t�E/:@��4%3?�
�z�'�P�SƖ#c�0h2���;$�x��'2�IɆ
�<+���;r`%5�0E��'s���#l�$�pp��,�`���'y��C��4�
�nL��Q�'����͓�,�����=E�8���'��� �ѝ^�\\��D1�����'���+u��P�%�W@^0!�P�+�'l���院EfVH���AK(��'�Vh��%S��p��-7N	��'j��@��Ȑ������}����'�����Ն	�
, P��oj��'��1�TlJ�vB���0j�0mTʑ
�',��F��bV�@�@ѵb�ݣ	�'�v!9TEFr����ǁ�W4J
�'S�Lbb")5j}����K�a`�'�� a�b�\�����B�@k�'ڍ����DС�@ҿlJ^I9�'ͰA� H��k�L�󃜫5:P��'/K`ㄊYRҀ�-îF�(	�'���Sf��!�E�q��
DP��'x �S�E���a��;"�A:�'=<�R.�?GJ��!�%.�B��'k�I�h,pls�!�$T(���')���aS�	]�@3a޽J�pY��'e�q�s�W`�@0�C�%�b�*	�'0�h�"�M�?���R��&4���'$�ygdӧ-�fl�gZ�0_�P�'��@����Z�Ȳ�9ժ�:�'�|��%m	9+/^�;SKH�-iT�H	�'���a��x�J2*=NS֡�	�'���0�ƾ<���k"E� F'ty��'���*���)�!�FF��<@�'Ѫ)�sW� �Bt�9Z�'��LQH��(X^0�b���3[Rݒ�'��L��I��P�y�U{#FLj��� ~���Nݧa��� �ܸz؎�yU"Ob���F��%(`P_��a5"O�l�WoK��4	s���M��$HB"O�Y��ɵZ١�F	��|Ju"O�xA�*X�
$uZ1�[��Д�B"O�L��cT�vS��
�C'7�f��"O�9K2�^;bz=D)ϱ"�R��"O
���Ύ.�����*t�kg"O��sA��5c=�4�r�*�q5"OVT��
 �z}�1�L�ge0��"OXm@���Y�.Q���S�i0���"O���W�	H��J���!@rZ��B"O,+Uo&4��x�6�0@���7"O�Q�G�2MD���/N�Sؒ��"O�)g+�� ��@h����C"O�M3!-C�Z��qc%��S�Vu)%"OD�pK -9~�t��	N%'�<@�"O�L��+�E�4�N[�8�P�Y�"O�I#B�:"N��2�M &�0�*O�ͪ�Lۗwf�Yfᐐ)@5��'
2������/�0�8�W"`hy	�'a��9tK�(�x��􈂼1O��:�'!�MSr�K�(���Q!BԴ( ��'���KK)$�6�#ݥ }�9��'`�|C�OL%|���)5�� ��0��'�z	b��*,�6�dV�)G��'k���"L9/|uKdƐ�n��'dz�"�ސ@��c���m!�'88���ȷa�*��P���zXP `�'1L���#�v����x���`�'��̓�$�F���P��oq��Q�'~ZP�� �a���Ґ��`����'d�	p�*c��!HU�'�d��'�j�c�T�Bw��k�/�Ɓ!�'$h��b	<�� ��O�T�t���'T�X�	��?(Q�t�YS��@
�'x��į-.[�}��@S/�p�	�'��3Ā�pk|P�f�K�f���'4 u�s��Yc��Q�"K�:h����'��e�AFPkP��|ކ%�
�'ڐ]����
�
4`��W�>��l�ʓA�L�i�NI"M<��c֏֗"����ȓ�� �Ó�NYk��@U��U��")L�%�ӒS� 8��� ���$�N	#sW�e������*|��	��Gp�3�m�0(�av�êQ��J�B�T.ށ1�0��J%~��D��wV.,�T�j� � Z�z���Y��ɰqk�4>�����K����! �0dO\�3$�A�9Q�8���8dhH�&EÃZ]�ؙ�j��1�ȓ.�L�h��>u��-9Veю	q�5��m٤����:��0����#���ȓng)ôꗛn=���陕)��Ѕ�HP^���®_�����RF�5��vȘ�h����m��Eq�
Z9;M�ȅ�f[&��O�8IV����
dq$نȓG�BI`�h� %��� ���C���~P̔�R$N�r(��V��:?W6E��E�`y���!#��EX�I^�3<0��ȓt��[��;kJ�K���
M���ȓ!�D�ӖF�6n��{�FͅD��=�ȓJ$0,��K~��3�`��[�|��ȓ-|��K��,����b�j�\1��S�? `��H�X`�Ԃ�N�֤��"OHY3��P�vf��§�z��eY'"O����I
gŞ�����@Ph��"OD���⊸_l!�bBT!pT:��"O�yz�"��м�#��K�H(�]PW"O�����ij� j����\ ;4�'c��`@��?EبЖ�0J�*��n:D� ��!�.~1\��(�7<0�1ړ�0<y��
ќ [3�Z"J��B�n�<U+�*c;
y�7�/��%`�D	t�<4nU�=�d�h�*�!�4*%em�<��Ƚ{F�X0��;{����b�<���CX�qb�3}>D@I��c�'�b��!$���sT�^�D�(p�1㜴94C�W��٤���e�����ʓ�0?�F�D:#�,#��� ��x�c�a�<1EE��	[�	u�<&A`SA�R�<ya�L�(Q��߲#1.M��L%D�pSkE�7ۈ���]�)��a�'�-D����Bc�ꈈE��*z����?D����(�Lo体ff�:\�DɁ&�(D�\Zu��Xn
��7����Agi�O�B�	�:8�0�""&����O�JB�I8U�H��jF#qs��x7n�z-�B�	�E�ܬ"�7@���@��e��B�I�a�1���E?4�(�A�e�3TfC�ɩs��۴Z1tF���h�!$4 B�	2|5�A�Ó=~�8W�"HB�I�.R�}��ˁ�X�PP��e��o��C�I;b��-Y`�,)Vc7 ��C�ɧ.yrԈQ��u�0��BRpC�I�K�B4(4�]<W"�1P2�8��C�6Gʰ�����|�v�R� A�s�C�ɴ
����e�C�Z	L$���=� C�I%�nH��<`�j�A��A�k"B��(�u����dn\�1�a_>l<��O`����2����1�R�uD��g�!�$�$�Z��v����){��\
`�!��Le�({qэ��d���s!�䏥S.`)r�g�'}ې �d�+z�!�dC��(�6s�X���Ń4�!�S<O�@�H4��1Z�x��[�Jo!�0z�K�2:}��E�У~��D`BS����	�y�R������ft ��e�@TB䉑qs�Q��E���:%(ЛfQbB䉆4ٮ�z��ŝc�[���A�C�ɢR�:\���s�)pрAm�DB�I.	�:� MK�q��U B�,F�,Jw�W�hm�}��-�B��*�*��'�J*R�:�H��I(h�&B�	�D��s���'�Lr��,�C�IW ��N�.J���&��6JB�I)sI�8���29 ���:0�&B�I�(wlt����/��`��ۣ?0\B�ɔ N	
���.w�X�2'J�0�8B䉘E�P)`�Cƍh��q��/��B�	�e��Dw�?@=�^����D%�L�nP�r�)�'�Η���;�� D�|�Ҋ�J�b��[�l(�a=D�T�Ђ�����أm�0�\��B;D����i�9�*��fO�;6,�`�7D����Oh\9���	�N@�-��7D��S�0�����C������)��x���A���/g2k��K�F�Q:�I(D�� ��'��q�~�2��A�dר r�"O�u�ת��@��j��E��x���"O���Eg��Y�����)�$�r�"O���K����b$k ��P�"O�Ѻ��X 0j�Y�SO��E�"Oļ��nؓi�Hak�,�/u
��'��O��}��v�ȟ�
�.I���W�f�d��ȓ<�&��R&�6��r�ОL����}�\��Eb�;'������O���ȓ{�!�A���O�L�*T.Z� ��i�ȓA�� ��B��I��5J���XSv���z5�!�i�+�$�Ң�Qnz��ȓ���)�@,����$�	X@��D/p4 A�5��I��R5�Θ��f��u(CdG�D�I�@B>qv���ȓ<�0�ib���f8;�E;���>x������T�J�υ�jQZ0��'A��9@��^��3-K0V1<��ȓ_�8 sփǳb��Q�ϣ,����ȓXk�` ��J���G�#^r��ȓ}v��Ivb�+8���a���!�ȓ@v��͓�z�]�daR�<�P ��1��܁ ��Y��B���Ad���k�0p�]�"�2xIwLO����ȓt��p��F��V)�=A&a�_�����F�B�B��[;̾$I�芰2��C�	�ore�D��8v2a"���1^�^ʓ�?��|�i8ǩ���E� �^:}*���W����4X`7�H=���
��E�!D��k�K�\T6i����#)����%H?D��C���7������9i_���a=D����̭=����V��/.��P�>D�@�R���$�tʃA�&=@&Dɥ�<D�\[��Mܶy
%ႄ	"�@"5�Of�O��S�g���b����C���C�T�]!�W�&�j����ߗU�$}��_�VE!�_�>�P��%�$nZt�f⑍9'!�d��h;(�W�MiY㴡�*}!��üR�����E
-�2��s�!�䎭�*�S��ʧjF�[�MW�X�!�D�h��!:g�״�b胍�?�!�d�p�X���*�0PH*��K�A��|��4i���#��5�+~L�	`0D���aˑ����4-�J�R=q��,D�����dY���x�Li�t�,D��)���#DfxB��͓]r�|#Ջ8D�`)ن�"�Iń
�m9H� �1D�\��eF\���#�L%o.$��;D�`�N�\��8���ZH��J��:D��2Ϛ%5�cOH�;?�ih5�2D���aC2y�T����R�h�Ã�1D����o3 h"��y(>��EJ0D���ģL�6�F����1 �����-T���A�\?wް��n�-z��"O��p���1�nu�C��X7ʈ0"O����O؍&Z��a"�	�E�|LЁ"O�J7��9�*X�� �t���0"O}PփQ/\Ў��H�=G����"O8Ј�G4L�`����W���t"O�) ��q,��k�)w�n�IC"O � �g	�>�����W�b����"O��;Ί�F�9@tj�0<�|P��"O�s��N�V �G�ҷѪ	��"O>����\N)RgZ������"O� ��xS��Y瞔Ȥ�ŀL��,X@"O�â	�b�����A.�`Y "O���7��+1[Ԩc&ۄ���0#"O`a�!�1�¡3v�ޭ>����D"O��JB�![��i�D[�N���X���3�S�IЩ#�M��i��QC4�b�o��D!�䍁�.��R@�a4�)�����?�!�$B,+�,0 �b3B�8p��:!�D�P�� ��j�0bu�D�N�!�D��)�B	��ҌJ	h}�7�y4!�d��d�	�[JvtH򊟺V !�DX�M�j�i�m�<H�a��J�-�!�dƳf�$\[T�@&�΄�ɒx�!���Ω��h��P��Q��&T!��X��IJ�p�:9����-�ў ����h�i�
}�r�i&0A�C�	;&Jx��/8�
�+$�ºd=�C�	 ,D亦F�j�x⣄.}��C�	�V�}0�)�,��=y���c��˓�hOQ>5�6�ż.Ծ9�E[�A6�KV�<D�`�ahC	.��$�ã6
�G�.D�Xq�剶9�l
c��9
v���*+��~y��'0�O�8���51P��bmFJۺIH#a>D�Ģ�jY<_B4H�ˇRژU��>D��hf�QKo�԰ׄ(Gq�!Q/<D���K��|�%΃;~�T��n?D��H``
K���`��G/�V��;D��H�lX�T�2m��E�`$h�ff9D����
5��ƍ�#@�D�ˢ�7��B��]�'��К�M�2�T$#�fTy��A�'ς�+E��|<�v�&nt�8��'ހ)��X�d��a�&�<d��(x�';Ɛ��+E%@J�镮նW�F�i�'�96Hĺ
i��P��S�F��r�'��$C6��+�n���Ϙ�Fa��7���lW��jAF�""O��Ɛ~�xb0�[�]O�}�E"Op}�r��-��ܱuf	�߆`Q�"O��%KԘU:H��" "���B$Oq��'�%.͛�J1�丂�3D����܃}��x)�N��]Pn�Y32D�hh��� m�<��O�����/D���#L�A.5B�m��]���aC ���O"��Tq�P9@�d�
I�	{.P�v!�בtG�)���zv(0��;�!�dP+0d�\��Ql�� ���e���d
|�R)��l�/k���!��SVV�$9��ܟDF|�,7�,K�kޟ�L��dbȶ�yb$�8[���s)���h}�d�M�hO���ɚu��Up��������1d�ў$��	0RD�pR�Q� b�M	�l�8r~�B�I��@S'S
vh��x���+Q>�B䉘d�~h6(۽HR��R�d��B�I�G���{�ķW�$��ҩR�j�$$�	J�$�V��k�p Q蟐p�p0�#D���p��X�`x�� �c�qs7�!�S8>��4)ɋ~A`$�b�Y��d��ʼ<	�?��DRqf��Z>N�`��i�d�ȓy^~m��φ�M��V�̙8h�P�ȓ3����PA�>���;D�;0^Xt��{���ej�29<�A3�n)lJ\���'��pS%��b�F�
�-�|��'����Bf�I��1R� 
�*#X	��d ��0bB�V*����RD��}�x,��|rƧ� �� ��O_��`W�әW�U��"O$�r�&@�/�,��G�8f�f<�"O@���˘�w�2�õ��b�Zu���'=1O `z��)D;�US�՚f�ɣ0"Oz-�q��L� �a����`��"O@QA����j7��%k�"Of c�%�th8�S�	��U��#"ON����
������!5j�إ�WK�<A����1�LM����8����LZI�<��)X�C���@��&8���&�F�Ic�'�1OHL���^���	�T'_�'k�(kT"OPŐ�(7��E�V�p�r��w�=D��#HE�f����v0�`��OƢ=E��*%A��ulݑK~�a�o<l�!�L�.�<(��������7@�!�����1 b�O�`�P󫘏K�!�pbda��ݜs �X�
��q��C�'T1O���Iܼ`E��0��e��"Ob�D�X6L}�5b L��W��3"O�t��cP�}� �X��F6h"�D�b"O�\��!��uA&9(P�ńhP���"O6�a�F��̝��(�jUPM:�"O��))V)�~9��aI´�F"Ox\ �Eލ*�8
ǅ�`�)BZ�����,
�FЙp��+bN�K��Ǧj4C��&RnX��aKE�p�*Do��:C�	�`���t�Y8�t��шϤ(*C��+<�hA�r�?X.�����"k�����*�	�!�f�q1h��^@a%@_|h�B�	�VZ0qPAM̷QsT�sR�"/p.C�	0
����,�5� ��sL�,�8C�ɿ&��h��/���d���q�^C䉍x����#�*el��^|=�C�	5n�YWhE ��)����KG�C�	�ʡ�VIQ a��Is�m[s��<���.V@r<�Lצdո�c�� D�t	@�L;FQj�k�hz@��1D��be�_e�l��K�=LK�1�*D�L82�A-p ����ˡO=D����^�:������u�;�#:D��� Ő�U ��dF�?U��H��8D�Ļ�i�'�(!���%.`���5|O��!?���34x�I�W�A�5��iR�+i�<v
�5(:��@�V�UhR�����h�<)�.߈s��e�$O@�%��gD�cyR�)�'bexa��D�W2�c@䔖 ��ȓi����e/��d⬽�VΒ[^h��7����"a��Q��h �W�-P̈́ȓ~�n�P�IS�Iε���P*#*��I]�'f|T 5G�Q���aL�'@���
�'��� Ά4�Rؠ�ɬ>i�u��'�P�3��-ݒ��c��2��+OR�=Y���P"�2�	c�M�|>b��񮔺9Q�	ǟ$���I^�O��0��ʡM�"�c  �!w�u�	�'��Q�䊁"ڞ�2��ʍ7��]
�'���9���:���.�.C�����'�`T�X!#h%��:	8���'�Nxf-�t�Xԡ\�8EV��
�'Q�e��}? ,�aB�A|�e�J>����i��A������3�8ȑ`'ͪA;�y�	�.�j�k��:
��WGXr��B�I 2bD���ĸq�5)v$��mB�B�	���e��$�B}x�6ȑ�y�B�Ɋh`���Ch��
eJM��y
� �`x��7qF0�s'�<	���; "O�MAc�E>jf\�0T&G-\�@E�T"O��cc��!6�/˃%���1"O.!(b��2�|qDF�,��0w"Od�RC��7�93��;ir�+c"O����>{q��"[������"O�A��D��P�b8�ա�h^�(��"OU2��!s�ޙZ0�ƻ=cxdx�"O<ik/ּ<��So��JV4�*��'p�I#z�0�A���cS���ee	�IB��O ��ޝ8�y���|��C��/v!���5?�t�`!�c쌂�� 6!�D���(�$�ޗ ��j�v!�I�����B�8J��d�!��{�!�*�.��T�8��`qE+�C!�DӉ2"8��˚�*��S�I<w<!�D�&ܽꇋ��.[�P�B�P�!��R:�*���ER�Bp�h	��S�!��	tYv��ӧ������]w!�dL���J�W>!҈��Dg[�qe�{r󤟧f���	a-�Hc�(���/_�!�DC#.�M�p"@@X]pt�;$�!�d�6�@��w�W�h��1�R�6�!�B��L� �%��zn����'��!�d�8%����&�B�"e��g�G�!��[\������S�X$���J�B�)�'.��$"���`8���ZC��K�'�$�Ů�.�|�P�'P�:�����'��@��.�)+��9��©+� E��' (Hw�,h&�h��R�&����'?(���j�%�TC���$p��P�
�'�FH�)�G3�Xp =[�b�B�'�,�g��0ՌD�'�E�BQ���$�O0㟢|R7��1C����<�
��w�<I��Q�t���f�S-����o�<�D�]�U�n�k!�.$C$L��s�<)2�ɖ,�\��A	+r�>��'�d�<V�A+Ktx�Q�l^�����C]E�<i�X��&���S,JA�y{��C�<��(\�3����Р(j��HsDA~�<�J1	�P*�c�\0.��/D�<���1����,ՠU@��{�a��<)6@��>B�Z"��`�{���t�<����:܌�� _�D s�r�<q�H�!ZB��cAg�`=ȴ��t�<���f���P�D+�8p& �p�'?ᡃJ[	s*�աbhհ`�$j O$D����a%!)��(�搂_� �F$D���P�@�Q%z@)�	L�v�\�@vJ"D���թV�7<y3�B�?X�J�R�?D�ɇ#P�^�#��JuԁF�#D��d% �V����� 5`6��P�>D��a�Q� �PqdkT(��H8���ON�D ��f�'�����BS�-�hC�n�Ob��
R�'!���d�Qڄ_=ul9�G�ڟ[D!��2h�@�ؓE <�@
 I�!�DZsĥq��� %�ih�
Ύm�!�$�w<I�c"�/Ae.8�
�z���Py2�'KH�yFi��@1R�Rs��_N ��']��i5�=LYLP��*΁U�Rl)L>�*Or�=��PQj����׷<#���EZ� f���զ��r���1e��> D��7�� D+ɑ0NйU�v���� �J���X ���Eͤ+�ą�S�? ����޺_�]svȊ9CW�bP�|2�)�#�^4r ģHP��b��'�8B䉂?	��,�-~%<\B���eB�I�5lL0�6��yp���C��:O�V-sIA%O��d�p��%w�(B䉭C䜬�
�}D `QB�P�B�	�Z��5Y�*�6��4k[��C�	�#��\��I��n�Lk��G��B䉙���پ ���� �rǆB�	Y�rB�	�("=�ǜ�H1V�O&˓���'���¶%�R��S�f��ɢ
�'5t�"F��2��y�� =)��lY�'LL�w.M�H!3!)�PY�y��'/b$H��DH�Xf�+}�Ĕ"�'�\����:شm�bmM%ab�$��'y,#Ga�l�@H�h �X�\4�'�V�yWC�J����
ȖKW�\q)O��$�<���ԟl��A���3w\ R�Ľm�^-�V"O��0%  �jz�ˠkT$rD3�	t�P�� ��m=~D(��J��(m6D�p(GBT�l5>�Hb^�R�&��3D�RgJP�_RdH��^���|���<���'.Pqǥ��ڽshM{m�B�I�a�t�K���vpX�f
�����#�[(�ɩgD�R���Oal�ȓ ����[ �n��1e�S����ȓR� �j��
6��vٸU���>A��J�c��D"��Հlc��ȓx?�1X$� M��a.
�jD\`��b�0h��Ĺt�􅹇�߰kj�8��w�eڰ@�gY���`���PJ���L��1aE�b��y1WΖ�@}�l�ȓت��d�<v�ܱrb˲����ȓ9H���H&P�����Z0 O�H���� �)A�PG�,+�� @�I��2�0�*ƩDG���G΃�G��U��=����EM1Ku����W�G�$�ȓ�§�z	F9� ���B�" �Mʓ7Z�Y���O��̆ȓ6�,YS�^j�P@�u�.���z<�(��c�6i�|id&2H���c۠,H�/�&q	R �ǯY�}T�)��{�D4�ըl�J���F�@8�݆�m�  �TآA����E�%:�z��ȓUd@�∍S�i§��|kL��ȓ|�̱Q�-�pb0m��	>�1�ȓ��5��v$��`��)�̈́ȓ����'b*�]������Ąȓ��I@sLSp�\�d%�_ETd�ȓE��}a�C�#�(��`@	C���ȓ;*�)e��z�v�Їj��IӪU�ȓN�����8�t}`S��:5�*%�ȓv�\5q��č�
`�
Q�g����v�$��A΃ a�v��iB5B���'#a~�É�!y���@�� �A�B��y�ϋ�����Ģi���-?�y"DY�U���3thZ[�e:�Ejy�ȓ p�P&�ƥ��5y�|Q�i�ȓ\��� ����\J¤�%k� p ���ȓ3�p��S�?e��4���Q�b�n��ȓ&;X����G�O�p��sj�2Ȇ=��W{`�#TC�-B68C�,�,=B��ȓ/���hP�ț2��{i�$o��L�ȓ=n\�KޝJ�����!/����S�? ,��ꓓ���o�n}n�"O�IZ�e��Vvz�G���p��"O�,p�/Ӎ
l�I$��<g8�{a"O��IaM��.=��I���$��4auR�|��ɰ
!�VU;70�Ԫ�FA�NI.��'��Hr�k��@�v�q�\�? �u@�'�n��5O�s�}��eQMO�qY	�'�ԙ;E߼>��})�	B��
T��'T�T��n�dQ ���B�����'r�$�7/�8"8�Z#�#	��	I
�'<.�Cp��4�~��7O�)W[qH�'��}!/���W�F$&k���'	����Q�x
i
Wi��-��xJ�'$pi�!˖S)�E�c �V;~Lp�'��q��).X9*c�7��8�
�'���R�!=v�
���C�@%��'G�9[�܈p�N���Iҥ<�0�r�',� A)�uK��ӰFŎ4�ؽ�
�'���q��'2�Z5���3j���'ɨ�z�H�>UŸ�[D@�/��x�'�.�S ��2Cd�j��"x�l�I	�'�^u����|�tDȤ](X�ȼ��'�l,�1�V?O��T��Y�d�R	�'���q�3nOjA�F�YY��j�'⬠VиA�VaJ�J1T��	���!OʱAF�a�B��b�L:	��lÀ"O
S��2�x�x�!�)j	��"OfP� �4e�������b|��y�"O�����Cc�h��JR�\ʲ���"O~i3§HA�2�肉�3�����"O��d�[u�DjH-�L%ɐ"O��3v͜��xP��>�J� "O�)J��:4������%�S`"O�au�g��u���� �2"O(���MP��1��W�pS�lzb"O�:��ǨS�.��Rh�<=�Eq"OX��IM,N̬U���\.Fͣ�"O�ᙲ�)S�SW�C8O%I�"O�@J��]I�\�S�E"���a�"O�-h���
��[uBN�	��v"O^���.)����k������"O��"i�Ku� 9s�97�,$sC"O�"�$��]:�t�fAB�+��u"Odx��E
�Z�x̱�iN�b1�u;�"Oʔh�C@cx�#��K=l0�"OdQI��J�+X�\�e恌x�\)'"O�9�#��)�����U�d�|���"O|a����n�<9���'ct��P�"O$�ʄ�L�؉an��?��Z�"O��\J&l!�Z9{h�ꡬ���O�#~bG�E5+2�#�"H�m��HӣZ\�Is�Ƞf�:�6�QI�~'@Ԑg+D���1@W�?_�P*!E۩sh*�y% 'D�H��MVC��́�,X:nw08:��%D��ڂ�Ѽ.��9A`@�c",>D�س�X$wFb����)/��׉;D��!��ҭ&"�M*r�[��8�qD9D����K\�W�2Hi���$},y�UF7D��ر@�2%��y���]{�����8D���V�T%N�t�oƸO6P�D�+D��[���ƌᓆC�y���-D�$��I�@H�G��V�D��*D�H Sc0 � �0�*PI~4z"J)D��ejP.��ȁ#O�n�C�!D�� �y��IGr���	tҹL�q�"O�@	4�,{���Bެ�µ�"O��8+�2�(���,q��)�"O���'B7�ܒ�	�FԎ�X0"O^YQ�n@
q|��6
4R��u��"O9�2�ٞ%�vM�S���%�n0��"O�����@2�����ɰ3y��"OY�Ù������ɂy�tX��"Oа�E�*.O�i9.�E���B"Ov���@�x����,K�4djp"O���|��1�vLR�	 q�E Aj�<�f�06)����/p!�Š֫�[�<t�
�՚A�	�\��!WO�Py�*G���� n�;K�<�Hv�K��yI$QB� 	 ���֐�U�N��yc�7O���@�z��1�3�y)�	� ,��ß�#�$�3DJƯ�yB#�0Lq�����j�p`�pH�y�h��z��ei��Ha8}��Hҹ�yr���Y=d �`ƏK>����d��y2H
�k�V���yh
� w�	��y����e\l��PF�j�%�V�B��y�m9v�ڗ=],�X�Ԭؤ�y��W�p�t���7Ԇ�p��5�yR�A�jv� kW�:3�X}�`N7�y��	��G
*��*��Q��y�G��W������F1m8:�ȣ	A��y�'֜ .P��Ʀ�'c����b�L��y�B>\l�s竇�T�hI�n܃�y�F[�7��* `��N�n�+FmW�y�-�&���z/ь�Z\�&Nʛ�y�O�J���X	l4 :Q�I��y��ҷ����)��D�Q�JB��yr��r�<9{&��)R;��`$��yb��*dX�07�G	~�J�"w�yR�D&0}V��@ƁqBe����yҨ֦k?�p�]�}C���R�آ�yr�4m����C�_pf廂��-�yR�N�5�ԢSAP^Exb +�y �e�q�"��	P�Ё1#���yR嘼$�l�y�)_�������y�Wx�I�@���~c��5��y���j(������"y���r�R��y�c�(�d�zG���lF��� 6�y��5����e�2bU℣���+�y�L]�f�L�B�`�_&��M�#�yR�)J�����aP� �+A��yb�ˬ@r�d��5�7��y�NΫc;��A�1���V�*�y2�H�f$+��)�� )�`ф�y�U7/=�3b%ÐQ�R|�!�#�yG�&?���ɧ��2J�rQ�A���ybK�v�H533�Z?&"��A%�y�⏣U�p1բ`L�PI�y�b�l�����Yo>�����y���`�<䍔X�t|Y�j��y�OˈN�­ItÞ�IC��x�g���y�聀!�`=�r���U�{DĀ�y�:DY,��� H��=ASOW1�yboE
?�)�U�<�ty9R�]��yo&Lm^q���ދF<UB皀�y���n�x�r᥏�kz+A]�y�f�N�1ҁ͢dj8�d���y��6cp�c7��;2��r�̄�y
� �Cs�Ñp�Fl��&(x`�p"O�Ѹ2D�-_�P�c�0kc�{2"Of�;c[�*v�r�@�C��B�"OT��DG���욂�@1Z�L8x�"O�:�B
h�p9�-٢D��ͺ�"O����=�)T����T��"O.\W�9�xT��+ �*m �:�"O"����O/2$Z�k�*Q�%_RŠ "Oh���B)��9Rj��?Zv�y"O�1� l?�)`1LZ�Q7��"O<E���5���8���E�xa�"O�`K��P�8����:u��b�"O�Q���rMrG��_}���"O�x��X�I����Q�ߛJn��`"O\��Ո\?�Q�fl�4=��M�`"ON�y��~��Z�6��!%"O,d�`���#�\qt!��O�����"O&!vBM�}&z�:R���@@�"O���a"5�1ȉ!~<�"O&�qd"���
(y�Ɩ�$�t�"O�Y��DX�ޥb&�I�^��	�"O�H+6,	?++�T@�)qY�A�r"O)�AfB���$��B�"�H�9�"O}�6��rBl�"�p��E�"O������XH� �-i�r�P""O���84vH��ԭ��e���:W"O��1�N�
�� �L�s*VA��"Ox9bT�܅{ ���	5># z�"O�`˒
V��|3`#��}~lM��"O�xkV K�P!�`��Z=^��l	�"O�}�H�O&�@#�+.9���"O\�arJ��%Ж�ֳfF��"O�r@�[&F�,���)b��"O�Y(�Be�Ր�b�JB�y
�"OD�I1\pj�j��ʾ<"���"OJt�t�H��z��Oܮ�-(v"O��*3ň�^2�����:
(�Pr"O`��fD�h���C�@hBJ]�P"Od�`#�
U_<��]09+>��B"Ol!����K���{Go}$�,�g"O�qa+��Es@�4���"ONU��S�9��A0.n0��"O�S� �p�6X�f�M�D� �3"O\������עB�@4����"OT��A�\P�Q����W��p�e"O&h����RLAv!A�¤�"O�8���(3�L�:uރv!v�y"O����j�j�z�U�Y�9g��Õ"OV�{B�G�0�`�����z^���"O���A���nr"�KP#�;qe~U8 "O`mXv+��(���Ã؇c`%��"O��Rh�.�F��K{G�)�"Ov�20�*����A!E)B0���V"O���7;����`޴��T"O�U�7+�=i���"�Z� �"O�@h���M�ܹ����'W�1f"O����֫;��qqS&J�xB�pJ "O4l;�B
�D����+]2Q
(8�"O8����"����W�zVn�1"OH<�R!�ݮQ���Ϭ)\`�"OlL�3M��N���Ȩ�R�H�"O05��d����aa�$)˰"O8�9�뛕* �lX#�6�ĴA�"O���7	�S�p��-v�ά��"O� 
1�&N��H]�`bsnȭ0~�d��"O.�jR%K�LX��Y3�;#s�i9�"Ox�;T��O�X�1O�KB�;2"O͛f��,���äE�K'đ�"O�Y�!�[,>ϼ��r%E
�!"O�9��m��>�~PxE$�9�$�AC"OX�aj�<P����!U��b�"O��XD�Eq`�8B�J/-�pH��"O��2]����膯[� ���"O��ă�*��HP''P��qQ"OJ��7'żx|ąɑ&I�3���3"O�}�F��J �⦢\�.F�4j�"O��ar@^,�pH�!ڶ�T��"O��I��ּ;�����i�4f�}xf"O ʴ�A/�T�K�&� O��H��"OxEb�HK�B����'�޵�A"O���n�"	�v�[t���W���b�"O�U���M�4�W��4e~<m�"O�!u���"�P�!Z�v��b"OЛ����N�
��8L�|z"O�	��̚�����@�}��D�3"Oz�� �̧}�|�&��+�>ɡ"O�L"�JJ����Ê�/�i�"O0�³M\�i��P�V<��� �"Ore81O�>�%!�J�-�4%;�"ON�k`�.oSF��\1U�� �c"OTԀ!��U�`�C���2�t�"O�A�uk��t|�9�^7��pG"O�\�F� �8QJ���iN�:��e�t"O���&G�?i�6ͣI[ 
\1U"OH�a �U2n]\� �JB�6�y�"O�<�5�K�]���jg�ɕr�
�;�"OL=�
�"B
��I�O��,2C"O�%�����Á*��_̐P!�"O���d*@I�d�i�k���KV6!�dA��� ��4w�������!��J=�@���]
VPPu;a/�8!�$^�uJޜBw�-�%��zKB��'��D���T>�qz���
�x]i�'�
���G�v9ra��<N䌸:�'��!��3_t�p��Z�G��:�'�N�����4���ܺAʹ<��'�֌�c^��}����9dct՚�'u�%�E=�Vpir	Ee��0�'���B ަn��E�I�-r�\�#
�'��	���Ň"��r��Կ=���

�'�8��1�X�x�b�E_=^�]�	�'n�5R.m��A��j���X�C	�'[����Jֿ'V)�ģ;vq�X��'��Q��g��T��E�:A��<�':��+��G*U_�ͨCbeB�9�'�HY�!�'= �RlBP�*��
�'��@3Kɶ_X5(�/K(|ܘu2�'��#��3��IB��	t��	�'t4,�lΉ��P�e�?�h}��'��q��z��b3c�'��z�'K B �N�&�t1"$�US?�-�
�'Y$]Q��P����:}E�а�'�R��S��10\!ʴ`�$cJ�Y�'
j��F� O����*�3_m^9!�'xF��C-�
���0�(��܉@�'/ Aak*u�<��%�q �1��'��uR�jT�FȀCܼgcn�0�'��]���H).u�4F	"r�^Aj��� r�W앞%�	��Z�8�8�r�"O�9����42Z������8V��$R�"OP�r2C�<=>v���u����2"O*�c�T K�T�p!ϸ��a��"O༹E��*W�y	� � �t���"O�0�Uf
�*=>�s�/� qg��ː"O�qKq�� 1;ja�o�6zPF���"O�<�7�ɖz#��q��!7ڵ"O.��(֊X�h�'� 0n� p"O>�*3�ܻ#P�탡%_16���"O�1%kId@��}2:%��"O�P��) t{��B�Δ�Q<��"O Q{�kǾy:D@��ܱ`���d*O�T`a�E\�� cP�ϟ]�(9�'��� �R�.hS@-�(�(���'D�Q�هH�١7���&��0�'!��W�>�,,B��*/+�D��'ɂ�$Ț@�)z���Q�Xa�'|�!���
_�|�
\�=����'�<���"'��ծP9��	�'�� a͍$v�n(�$a��8�R`��'P̵�0�[
5E�ts�NŸ����'%:����&%�6�c$+�(����'ŘY��-��]��Lx�
 
#��0�'��QV��^�񏛦 }d!��'R q΂'V�䨩��Y�Xx�B�'�pX�C� �.x��J[-&ba��'��ٓ��֕v� U�w�E �,x@
�'����w(̍?y��[�y� �y�'2Z��a� !A��ͩc��l�@]�'.�CЏ;ך���"� 8̜1�'����k�<o���m��/g���'O��s�dS$/fش�qg��&�Fl��'�L����]�(8��2����
�'
A�k�#x�Dzŋ�=^F
�'�h�Q�	��i��`���)K�'�l�pŮ��wL�A�n[LYj�'�ryZ`
�L�H��A%��_�*�'�v�ƕ�p,F�[�NT�)n}��'#��r�$��a�z5��/��0��'��](d���E��m�8�'L���O�_�l�b$`ɮlo��'/<���܅r.8�9���^����'*^���C������@!���3�']2с�I� 3�H����1w�T-H�'Z �j���ebؐ�oS�i��C�'�>���
;��TY3�@�y�H��'��Mx�W� �ʉcS�x��L��'L��ۀG.o�$q�G�^�w%�M��'��e�&��7SPB4�b�O�u�ܥ��'�yx���]�p�nƃp��r�/�qOV��Gކgލ�B�
&a 50�"O����V�#����t�a������c���A�Z�jvj�
$���P%��y��Ą�.�D9%�X���#%�H}�ą�d�P�
�.��I�v�-��	N�'׊�Z�憎F��,��-D:R��Yiٴ�Px�II3_�)�ⅸ��уTX+�yB	�+;�Y�$�¸P9�I�Ģ�y�K��#`���O՜<a�Q�O6�y"dJp�(Ɉ�� 8�t �j>�y��9w���A�$��_O�B�I4 �f��(V*]�(���F�<��$��D��L�L�����s(��[��"D�� .��h�a��Z� |�t�+�"O����H,�L����-�|���"Od�3BS��ܭ{����n��b""OT\��'��p��I�>����g"O@�BVa�5�Z����j�ak�\�L���2O�a�bؕ$�bNO&� ��������'�� �"�&v0b�1��C
�C�'�, �ѯ��G( e�b�Ǯu�*���u��B#` m$�*%
	tC��Kg�B�<��gK�W��L�So��k7���W�*F�v�3�)�矤�g�[;$/.�2"G�I�����*�O.�O.��7閉@F$h�]�z�F��"O�	����!��aB*�����"O�E�󆀾gC$��P��
Yu��P��	d�O��<S�M���A3��$x$��'E����ٿ	Mh��h!n���'W�i�d�KN��y/(E����
1�$����H�Pi�%ՠ$8x���2���K'��F1��M�:6ąmIܓ�~���O8Y	��M�1�.�b�F�E$�(���v�O�I��.�>O0�]�b��*5�N���'���(U�\��b�iu��zY|���'��II�|*H~j�@2k%���"-�2�����l�<y ��X�D ZG#O����Ee�<a�*�:v�`���*���xե\h8�h&��r��Ū�
�`�͌�i�P�8�M2\Oftۈyb�ER��p������pP�P��y�/Хn�4�U�ěDj�	ܺ����y�T��'��?%C�{� �`�	a��Ѵ.M�<IaI	�y0�K$��;Rd$OI?1J����'l����A(Fl���.V@.v� 	��ē-���۷L��T���Ǫ��L��o&��<��yB��K�,��ac�5Q���G�߈��<9Ҕ>�'LF`�'Rt��ǂIU�A��'��A55�>!��U�	��X��O^���<��}J~��͞�N�q��,����p�Zx���'����0F�Aź���?.<��2�'Kax�dZ@y&���i�:u4�$��)ӈO�R"�S�_(��i�?+�BZՏAh�<ɔ� cÄKR��v:���ȅ�<Q���S&[�����J��	! ��6����$8�'O�cw�ǋ=.���G�T��`]�4&C5����H��J4oZO�����a��a	8�ˑ�E?	:P�n�"�y2aV[K�H��LA��z��
��$�<�����ħ:9�$��K�$<nd�'�D*K#����g<�l -�Xy�m�v:�kEF�=�?a�����i��R��d�D�}��� j��)��U���8lO`➀�u�� ��Y
QD��?P�Dh)D�@��dٜm�����w���D�I�O��=%>E� 4oW�ȘD/�+W� U �G,D��pIђi�p�{'�=*(� �)D�,Z��s�D�XeX�gh^15�'D�,�HѴ?\�1�6K@��%���(ړ��	b� Q4�x Ί1h���9N�x��6G�y{B��	�d�)�0SglY��1~���M�vD�ɧ!U�4��܄��g�$�z�P��hՕZ���Tl!!���;C�r��I�~���%��r!����-��&�0B���aĄ�.!��4j�y�u�aS����jծQ�a{��$�1<,�U�H��H�Y�
;or�y�|�2O���aז0]
�"��8����"O
��d�o��Q�+�}����A�'kў� =r�CS�@H�-{T�Ҁ�$"Ox�RQ쀲/�"�a���;P?��S���'
���>��B��.%J�̡��^�WD� ���?�y�i�"Kd��'(
C�<,Y�������0>�7�%r�����o@.����Lx��Gx җWq�%�!�X���	�����'ўb>u GF�]c49#`KR1@��]�l$D���t���|��M�r���!J$���<ҊRM��i�fu:���!n�<	�E�@�.�9&������������C��=���Q2���V��<Y��&�ӖRp�3�m��t�(e��=ܞC�I���:G *���J�$z1*B�ɟZÜ�"E!,Aޭ')��Cd�B�	�yt�0�E'���d���b�$��/aF�e0�霚<���j�%A�^B�I-_xJa�w��7|�4�z�!һ&4.B��jy&�J�A�b��Bpkͻ��#<�ϓy��9�(�6Vs8u	6�\���W�-i�+����4BU�3�� �ȓyC$�j�$�	2�ı�"XW?��=�M���|�/�p@aed�1+\����_E]���%"O�`�5r�`DY�#=^���W�d�O ӧ�gy���9���K�
W�D��$���۷�y�FҬ#�f�h!�� 9 @(�e`D�y�Ε��$����I:$0�%K���y�� �p���Ĵ0�R�	E���yBd�+�؁K�JA-"e@�e��ڨOH#*� �a(jas��rL����o�j�<)�J�dz�P�����4s��j��d?YH���O���!��aaɿAn��E%Cq~�B�	:�̘3E��u0I�`�T�%��D���Լ*S�rg�K9@h�� �r=���U�b ����a��$���8�x�D��e����6���	B@�ȓf�L�20�B%V���/	���A	4``V�͊ �Hہ'QW�ԇȓ/�v�z�OZ�q"4}���1m̈��Px`aꦡ�u�ΠÔ�&Azp���U?l=8U"뜹�sO�'Da����;��qɵoD&�"�+F�"˴8�ȓg�6e�4oi��b�  !k/T1��h�Ԝ��B^��vT*T����$̄ȓv=������M�&�� +�؅�9���t���kcxp��&~�݇�$Ȁ�[�lI�Y�-����
���ȓI}�ps�GU�%3���SO��	���0V9pt� �F����u�ȓmx��ز�K�X��y�EU�O�(��ȓE�A[�,dV�aх�>A�f��ȓy|,!k���:�l��Ǌ�� ���ȓ]�ą�
ۄO�2) �
�FSڜ�ȓ,�#6H7�ZPb�j����<&�q$!L�@�R����([p��ȓ�6$���̆$Zp���C�0�ȓC��� �<d��Y!K�*.0��ȓ"�H��ǭ��V9��gᎰeRẗ́�j�Ǐ�wP6�裢�(�!��W�.���)��7��eЦð;/ZQ�ȓ@��Y[�n2{��H�C�_��Ն�}[`����)��Cuʉ�;yN���6<�+wk[u���KW@'lX@�ȓFFZ��BюTn�k����C�⑄ȓnb�(u�q�|�3eĥR�5��S�? B)�$��*��4��młJ��y�t"O qE��*�`+�^��س@"O�h�#�H6'\�j�`J��vX��"OXR�K�A'&A��`�3Ԫ�1�"O�ɂ���6sʢz�Q/���"OFsO�8����aO����!�"O�4Zr*��n��	�$A�,b�D�"OzX�oW1pE��PW�8[@P�U"O|�)EcC���Փ�mR-N+@I�"O�|����!u�0a)7Fl����q�!�$J�b�+��E�n]P��-~c!��֔�qfϋ*�areL4P!��T�iϺl���c��Dp�K�)�!�$�[�f�h�'���@bl�?u!��/{�ڰ	0A3���Tk�(d!� 6ڌX���Y붴YF�Hn!򄚥I�b���f�=�.E ��ۮ`Y!�DK�[?�9�PG�$���Hсߔ?!�ܕ(T�`�X�e�\�CꚜK!�d y�;�G��t�$f��H!��	:1:��	�<��I��UJ�!�Đ�1Z*��! ܙ1�,<��HZ�!�!�׾N���a�~aD-��1]D̩C"OL,q��; �(�tҘ�c"O��������3!�d�� "O���sCT�
N�`��9� �"A�i�<�L�-��[b���)d���k�<񓤍�Zc�!Z`�+�FSy�<IWF��'��b�(��#�Cc��{�<�C%I�|9IQ��q'�t�0�}�<�EmUx����'��8:.���h�t�<)����<�8Ї��,N;���w�<��1d.����Îc <i�K�<�@�����Zߝ�@i!c�<�5��1|�C$�t�e[7�UE�<�rEC	CRi1E��0r2)�5�	F�<��h�1V��D�)K��L�y�<�n�T�L�9C�Ofe"D"�`�y�<a,�p�&��g���U��f{�<YR���r� A��'G�A8P�/D����@Iڀ�v�ȁz@���3�+D���Q�/M��4#�BV��s�&D�L� K�3 ����Y�E�$�*�6D��+�\�@�$�#P���J%g.D������z��G��|Ⱥ��� D�|�����is�˓�#d����E D��Qe�cTv1&�03�J 2WH<D�0ۖA^�b�p(�L�Y^���>T�P���u�LS���U�\�W"O��c(ߏM�L=�A!W5l.!�"OHbq�9(���φ�Q�"O��IrB�'r�P)�.\c\� "O���ژ`H�=�F�.{~��i4"O
#p��9=D�A����#�^L[�"O���r!%re	�eI�;x�\�"O�H�aD,\~�q��Wi�z<��"O`�Z�k��4vE(w��y���7o��0y��y\��!���y"IZxݻPTgN�$��y��Z9k���#C`�Sx4:����yR��g7`���\^1^к��Y��y�˕�X��t�t�]�}�����E��y��b�VH�'̂��J�;����y�jT�{Ȯ���*A	v�$��u��y
� P�J� ]#0\��t-
�f5�P�!"O�������d�w�_�>�lQx�"OF�b#�
!h6��c��f��P5"O*8�e�/V eR�j&���"Oxa � ֘p&H����Q�%�""Ov��@��*C�e8����`"O�h;�@S6����i?��9"Oz�$'��H��Բ��K�<���"OJU�kM�b�:Uyw��	$eB�"OJM:��9#��hHS��8��m�a"O�\��
L�
c���W���c�Lq�"Od�e�+�t� ��;5��hY�"O6�{��(A`{�B�*|���"O^d��!�@fИ�����b:؃�>95G�R;�|2�GA�ȟ=SP��	T��t�WB�}t��"O��H���y�ty��P`�X"
�6����'�H�R��ИϘ'����;UT,I�䍚�I��x�P��*TAA3Xs��(f%�8�*�%�L,�Ug�aP���]��ш�A��12�e[�@�`D���"T����͕h�R��1��q�q
�3Qe8�p'��z�R�@q"O�yᢃLy�>�)��9���jaV�L�d��b�@d��+��pY��D�4J52Ֆ�rķT������ybB�5;ר����\�L�����Q,�d��m�(�?٤a޳z#��HM~�=�!��	ԌdQ��:�Z�s�C��8�Q�:s��	��0��5������Ps���r2�Qî�C��H #��}4Tc��?fH8ʇ�=��!�Nԁ�͌y�epa�����Н$`�����v�j0�+���y�̞U��a:�-k
���K��Đ4M��5pt��(��(�G5ҧ<����4�c� �U�����'�� 3L^H؞|�g�;B��%/�Jl$��c�Z%NxJ�3t�O\XBsi'���� g|��ܴ4�~�Y�m�8�L!�^�_4���q�Ծyv� "�
O��^l����d��j���p��՟zs��v�KR�F�Y�6l^��WGl����D5��,�0���iB~�Z"�>	����	4#�L�)1g�<�6H�'��(�!$FH�H�͏�h�|9rl0Dj܀�i�����}&��e!� sj�L[��Z�^�B�$$�	�M-j�P���+r	��*�6U@QC��Sver�Bj�e{�� 3x���'2��a�iX���NޕN��m�Ǔcy�AX�"�:xR4A�G��}"@{m\6k�}�"U>8���k��-D�Za -#�~����	��!�"4��Q�76�P
S��qx�+H����xF�ǄD�� f/�vh���"O�<���E� ����#�[/,Z��*��J3>HL<Z Hύ?��S��?��֔9pQ��Y�%��$�z�<�g��?���0��<��q�q?)�Hj�f��G�+LO�ي���8��zw�6S@L}��'����t(5Z�I�X�-k�Ĳ��W�D<��
c!D�(��)J�e_�a��R�Zh�rÂ!ړ�$e��D9�'#��1���1 �T [~{�1��1.���HO��ea�V�,��ȓDCԐ�Qʞ�:��	��O?xh���u�=���WwF�鄡�??z4���Q�8@�e��}���yT(-cT��=!��ֱ�����۬d]4\Qc@Z�}ߠ��6*ڸG�!��ɮ���EA�6�ٚ�醘[�#���J�DS0�4�?�'���pr�'E����ƚ4Y `"�'jr0�%E��{�r��ek�j|�8�! ̸XQX���ǛX�dU���4s$�h���E���1W�ax��!��p �.�s���%�i%FTi�1#�v���`�� �*ĕG�\��	l���!B�1�άh��Q�I
�j`��q�(O"s��­�?:�B��f������O]j��v ;~u�ܒ��I0  j���'���쏴�8�LG�4S�O�k��XsA�	�/�|���S���'-�r�б��2�y�`�%�#�^�2 ��£P��d@�1`H��{J~R��O�&��EI��%0idt�q�Z&"2�=d��p#�}B�D�u��^�D��a����>���	�B ��$�6cE8s~�'��4�f�E9r����4Glp@ �#�~�'N�|��3w�K�/�n�Qe��6Q�H�"6�;u۠�²�6lO�	Sǎ�U�? p�1'l�9g�@T���SK��Qu�W�q�4�{f�J�B�H�`u�٘P�l�)W��e�pc��DQI�������Z�F�|�C���$-�#?�3����
�K<�I�V�i�c'�Ȫ���|�H�
/�$<sz�8�l�#^�n�����$bYA���UOu��Hn̤B�HD��A�D�ޭ9#β>I�J�
\��.-}��4��&��,�%����Εk��K�K���%F�_����ݻ�����Y+Pv��j1�
yLE�f�I���1(�.oZ���H�8��#Q�ZҠDQYw���)CO&}�� ��6�uA)*�tʇ��4�b�1���O���,*k4���GZ؞Ԁ !�%yM|�E�TZ���6��K�-����XfJX�EωoZN|�p��}Hx �%��M#!�ʋ���8��A�7�W�AC��H3�����#?�'΂�\��-*�l&�Ix�hj5/�"N�fp0@�I�z�"������U�t$�K��T����	� ���O`��	?o�q��R�U�D���S�|��`O�T�>��5�>�}ҡ�]�%�j���e�T���PSt=����8��5X���LV����j��"�	Z��܁RI�X�	)�s%ґ5��d�W`>Y�1 �=].qc+ #�u/��J�>����(h|x	���xo�K���c8@���A�� Fڄ�AH?��;M��T�7�[P��N���DД�O���E�60�8��iJ�j� 	1��C�����,)�X4�5Nʏw�5	_:�����~.���;x���C�ȝ<oj]������'[N�vFص�}6��jy2dӋ�d�b�v v��[W�����S��ы���9�L9���2"�F�����=)����T3<�n��$�jW�Iڃ#�2)A.�e�'V�^̰4��$V�f�D�VF�g���ؕ,�JBpѐ!V?�� �%��%�5��!0�$)D��q��x�8�������0au)��Xy��H�*^�^\�M��P������۞!�:y͓\VD����=3�����̙Ӫ��	^BtA`j;p�h���Q�">��	7�G�"�+��G:n����'Jк���(P`)/۸hK���^�PtF8c ��${�P�Zv��;Sc,qEL� �\�e�"Ϧ���K!�}�Ӊ��nC~-Z����>��';��ňM�,���JSw�|F�DȚ'|���^�?����\W������I����"<liVO��~�q�L�]#�(2�i�.�!fb���Ϙ'zį���L��/"@Z�'�5����B��k�#���H� ]��L�q�<u;�dѐ�'0,�	j����U	��l�
�Jr�x������?Q�Zrh�i@�C�&��.k�<�D-ME�fm��.Ӿa[���g(�Z�'���dmF�O<�8���T�h8��у%��0�
�'4�Xx�)�%R����Q�
�M�T�	�'���)G�tpj���50�@��'6șr�f� &��#�ġ5S>]�
�'��i��!��Zc4���({�H��'��L �LK,�� ժ�+pwl}Q�'������d�^P�d
_jM� 3�'���G6&,<��Y�Yv���'?��y�e�>�P�rc�ǈO#\s�'!:�+ש�01T�zFk
-D��Q�'��P�q ���DH��k^���'����$�ǜi��#��l �1�'�^p/�d�Ht��搀�00�	�'9L����&r���`X	�ޤ�	�'�A3�(/_�P0�7��p�	�'|�m��J�VϘ�
F�(-����	�'�<]�D�xf*L�?��H+�'�轃v�٭���u�y����'?��P-/28p�:e/ƹp���'�mx�cQ�}Tz����?�����'D԰ΛqfPiw$bt(
�'�>A�B�/*���q�I�MI��	�'��z��n"
��@�\#:�2D��'NbI���9�8��ʄ�?����'`Ԡ��[�M�����F�+_�(���'�h�C-`4�H���>I�����'�0�(��×Q�Xp�׭��I�6��'eԌ�G��	t�e؇�1�2��'I0)c��]�?m�aw抪	�4�'ex5{R*�8!^�c�A 7|!��� ��Q9@��x�p�M�"O�T@��(7 ������A�9Hp"ORyV�W�	��󃍟�Y��"O�X�6@���	��@�8>=1v"O`�р���X �C��;ZF��"O0�����X���3+� lð"O޸��핏9��y��Ѫ
�ttp�"O�L�g�S>(l�����ҍum�`k"Or<�G�Ś}��Q�ê�=.�h"O �Aη ����H�WN(�"O��)��H�����h�����"O��"��&A 8�ӳ�¿z쾜+�"O1[���j_\E�4	�:�
y�7"O\�;G�6g؜��i�,x}�t��"O�����(	����HR"2q��"O�`d��jg(���ʩjLf(��"OyB�Eяt�
�!��($"�9��"O� j����D&�yu�$
��"Oe��/��yHR��E��]��1��"O>L�V��E�� @�B�x�e�w*O ��"T&:ނEqbGH�,K��S�'y"5@��T>|Y�Ej��0%��̆ʓy�tAUi�	�|�1��?_�M���$$�B�A�K���V�س��]��-��-Ə 6��Mʭe)P��k<�Pւ �>9���!H�ڜ����h;7#Ȳv�1NL���ȓl^�9p�I�P~8(��.B�^0�U�ȓ;|�)�$"B�`��0�UJ�ȓ���kf �	F2�SU)Ve�(	�ȓ~��q�J��Hh>�c�fTt�ȓZB,�+eN�%5�©�T�yJ����X���#�:q��24�Y�R��d��L�\���:m�v`rAOC�"��ȓG���aW_~�䃁d��(�&�������WEܡM��e3�iO *��Յ����r�*�g?έJ���xܲh�ȓ)dH���K�7��j�#�#��x��v�Ȅ�@Q�� 
 �]QY�����l�����8�Pu�AX���V�<Y�
:P�A��@4F�	q3A�i�<���A�[(���u�R=Vo���P�Ed�<��i�9Q��3B�9Y����'A�Y�<��B��]̜,1�-����@ �Y�<�6@�F��p��Љ&�FE�",�_�<�1Oڞe�2���M�w�A"v��Y�<a��(!��}�D`��8�~�B�%@T�<���(p
9x�ı1�Ċa'}�<��W�!&�h&'EIv]�4�_r�<᧪�:wj��u%߇����s�<i�/L���C꾈�#,Z3u�6e��1oP��W-\=��!ڡ���uy�܅�$|�e@���E��1�Y�v��������7��+r$���Y#BńX�ȓk��S$	9n}��� ��l��ȓ�4�"�d�����iΈJ�F!�ȓT����I_"=茌�G/�19�����eb0`aE�i�1;�K�(�ȓSI:쩂�"gT�����]�ZL-�ȓ�v٠��˞-�2 s�iT�K�4T�ȓi��\A�%
������N	|��ȓH#�|�d؊>+䬚1K�>8��ȓ
d�!��j H��SQ�]?	Ej!��d�h�!ԧ�)ji�IE�ɣi��ц�S�? \���,`r��c�_�X{�9�"O�X��G�Nf �:vc�8PV�U�"O��z4K�E���{���'�Ll5"Od���"yj��y�a�2P�j�Sf"O�����F%� [���L�"OX�d,��p!b���Z�hc"O�A�EL~��}{0�X�0�����"O��Q�j�Q0�$ӆo $q�"O<kg�&o���#я�
Y@:(�"O��9D�]�C�9���,G�rX�E"O6�j���4�jC��hZ<+"O��2��M�T�C�+�<][�(�"O:eC'+��:��Ȇ�±��H�"Or�0v�ϷO��8ǪL�&�B�J"O: h��+Y����R!t�D�AW"Onx�3A��D��5��ޱY�"OhrQ˙�|�B��H�+��$3�"O<��@�/<5�ԇ�0������>a��0b��1��ȟ���wn_f���s$�J��yP"O����,�4m��q^�PB��i4.�Y��D��'��:��N��Ϙ'�z�R�`��(�^�x�����%�Gw��pۇ�U�"�܌��b���Y�fy�&�sD���!��0>��\��F�	#K�$����l�'�Nh����#�<��n5��	� UH��R'L�Nd�(��E�;�!�:�F-s0�H5~F��R���V��I *��y�&�oBBq�!a�O��x[e1q��	s���,��ls�'�(���KB0{���┗z�Pt"
�]�*��^.@Q���%��g�;�0��I��,�)$��3�d����9�$1A𫎓l5F��Z��"�Ȃ���GH�/�ea!�(�O��Gxs�� ����!4Љy���	}t��AVB��j�� Gf��|1��[U�$��kM-3�,�ؑK�U�<Ib�B�N6�]zя��0z�ij�c�Lyb�>���af)�h4��� ��K��Y��G����O!�ʓeH$D�Gl$lO*�#B��~P2xX�ښ���b!�;&b����'�Ҍ`	���M�L�-"�+BF���pH�!�e�4`�4�JBብikbt����w4�QlD�݊��`�z����! Sy"�G�_�u���\�T>�B�#N�Z��9��9p{�q�Ǝ;LO��UJ\�?�:˓m���a�{� ՙ��ι:t%��FI�z���]���O�h��1J�u���Y7 ��$��� w��y��'q�&���I��w��	w ��J+j���N�:����: �����ߪ�L$�p�wz���̄���|r��3�lx��
C�'���* u^�}#�
��c�(p�ȓ*��(� �5v 3'C��9nl�Ey�f�/���P�C�O`�y[c��y ��*6�ŵ"�x�B
�'�4Q0S*K�Qa0u3�iP#��P#0��\H��S6��)���rqDLd��D�b$�l��#'�+D��+,���x�	��*K
 A'���`00oO�@IB�'��l�S�F	������[�`Eƽ	�$Â�Sa"�M{��Cp� q�x�i��s�bPB"O��0�(�T�
\�`�H�"�d���I�`9H4���Ө	�F0�
(SF��[�ɕ�G�B�	ȁ�r��r�);%+P�"��C�ɋ�� I��ET�L�bb�9_B�C�	�`-��q�^N�(yٕ�պ�jC䉚�Y��O5c���*ǂOt�(C�ɚ%�����K˖æ̳OpB�	�;pU ��!8�N���O=FB�I�/�0a*�Q1l�
���+ʐO �B�4'r�����?y���tOU ^�C�ɕ>=�DJ�	>���z��r��C�
����O'g^0 w��)t�岰�
�a����ڥ����zb�@�!Ɲ԰<A�iG�w��H�L�Hi��"7 *\(���-c?L��`c2D��̘�@*D0`U��y=2H9��3}��4�tx�"h�g>� $�V���0�!�W�9\��K���@S��2r�qO>��l�~���SĠK�95���׋�<��'qbH3e�E�g�ɶ$��!!��i��:qj�MȒO��!�E�Oʢ>Y2 �v�F�I�԰b~���@Xe�Q ���GZD������P�:b�ڻ?�xA�&�.>8�r�< @����$\�k�ژ��!G���]�=�
�Ò`WL�� p!$\�#ב��	7`����x:E���΄%�pX1�癆��ȑ����I���G�zⵇ�VN�q�e�:L���,��,�`�-~0��.��gL�ӧH��|�vJBCv� gKC�#*��iI�l��G+Jt:CO2�3��_L3x�q��ِR��"�ʖ�T���'�6�����.n���'<4�0�g͌/a�A`Ơؾ-�����0}���B�[D؞0�s��� b�<d��C�ߦGx��{�ۈ"�Q��S&.ȿ&%�i�O�C�/��R���ه䜎Nlpm ���Od���.N?&��O%�)b�\�j��ڐbM�,�j�;I>Ѱ"͢-�h��>�W�r��M�$��spġ��K�>�'�
�B���.-}��I̒�lAsg��?L�q�K.�!�H-U��s��@/m%T��&��=<�^�L���͚fyz��H����:?���'!d�9�%_�& ʰ�rƂL<��O'X�nQ����L�}c�L7f��,��6}�l�l�HeI"�ɄB��\��79�~=����6t��dG@���jG@xȜ��!��� ��1�B*Ev�����>���ěj�\�1)�6�b�'�Uџ(R�G�u�ʴ�u@�2c\��'7����?8q�͋S�ܟ\=�m����Z���\@��1g2L%�'R|"��	�7��� �,�"m�lD��A%8(q�@̂iU�=e�ӏ�yB�6��12�I�p�p1����Za10c�! �p�'n�E��M~�=��")O" �%n	�!�v<F�P��ѕb�SB�񂧑p4�Ձ,e�|X�$Н-��!��E�a{r�
�Y�Fm��ѫI-@�p`�����ObM*5%�:C�*�8�C@Q�ȫZw2�A$	w^웃,�%w��l��'��}��+T�O7�$��p�0(O<���L�%`f�	�C&q�����	 �7@��6�˗jj����l\�x�!��U|!�M�E�VdQ�ya���T큷�X^2f]mڀ7+f�;�#2�3�I��>|�ƀ��@���AW>n�fB�	�m0�!�,d�R/42�rAI�0�5x���SJ$��Iu��)�M�!K��qd�V�"��$W�!>B�j7��O��`�$� ��0�t�r�`V"O���C��7����T�`���剙[���
���;�D�I!
� �&4��AC�\y<C�ɫ}e��7�I	z�<�q̲Jp�C�ɍr���b� ���u�%��{�C��s�܊5dؑY�e�ą<b*xC�		ȴ�2-�6[Ǭ��a�
�"C�I�Yoz43V�ƴ<M�9��cӯ|P�B�� %D����2u�(�s�Ǝ:p��B�Id�X��䀻Z��BBIX�i$TC䉎]�<�c�i�c��C�!�;�,C�	^�(ː��Mۮ���-��$�NB��+��04�� x����^�B�	#u��e�f�޵����o�zzpB䉷c+p�g�D/֬q!�QB�C��	P��s��lߨIR��#֘C䉸 Ҍ���,�3V�� 2#�Z)sjC�	c� 9��;IR�h���.Q>@C�I�2�L;
f~Ȓa��7YB�	�Br��"'H-0�Z�"��2<>B�	�T��荐Y���qG��,��C䉇Ǣ����z�*w#�a��C�IU�L �$i t�%a�C�_����>x" ��/�Z8nB�FM�J��݉h�]+�.Xw��B�I�gޚ�D��:#�!��l�3.C䉔����*FEA�g^.{��B�ɇf�ƌY`%��<G=�C�R�#�C�)� @���جb-��fǦ�-�"O�D���?Vtt�z1+���@��"O�q�@gJ�L��"�G.'�`�P�"O�hPP�U�J��a��n�z!a�"O������r\�����Ys�4"�"O&d�&#bh�ʆ!VpJ��"ON���&�#-�Ҡz¡Z�Yh���"OXTb��&C
����aƔ`Ibi�"O�SS��b�������qC"O��IE^ ����*ty��c"O��Z(�-v_V��O�8�x��"O��/�(4*���!���|X�"OV��@Sb�,��44<M5"O�`��7e%���
r�tu�3"O��A� D�a
�=��05���"OP����U*�KU�۬�t �R"Oڽ
f��3t35%��.����"O��ʀˆ3^�:<x�C��[b֙��"Oִ!��Z^����՟x��X�"O���aKD.kk�kӃSl}��"O��z3�1DjY�v��7!�:5c7"O��P E�����{�9�U"O�E1�#Q��(sG�.S��<� "O@�3�g���^��B�o��x)�"O~�C�O]�~2�U`uǏ�x�nMb "O��"E� ���"�#�Ȃ�"Oֽ2!�I����'�I_�����"Oʕ��CH#L��tRBF'~����2"O<��V���Ȧ���J���(�"O��u��7|�h ��	{�mIt�O�����=]��>7�J�t�.$�v&D�ry����&��(Y�0���L�ɧB��$O�-�$��PAҀa��$+A�H��$�
���{��i�2�(�ٰOW���T���=��Ff]?���=E�	�>d�����HȞ\i3J�J�B�K��� e>M�D-�� ����B5��E���tܓ^� �Sgmڥj�F �$�̗b��m$>�j�M�aR�$p�k�13���\�D����)Q<�%���M�)9�O哠eS�m��(˼8�0}�3�̼o�XR&>}�G�y�ҵ��Sh��l�w�_ef��C�>zJ(C� e#ʨ�r���?u�h��JJ�B C䉄] �݊@g��g��< �!"U�B�I=W	n�S�-�@�88��Y��rB�ɺJ=Pu����U���Ç�7(�TB�	�D'|=P�#��ju��K����vB��.�$c0ے=��Mȫ!]�B�	�E�Fp ��L E ��b��m'&C�	�9�y�G�/�����)D-8�C�I�[X��a�I�c��5)���A��C�I�\YK��__<�a���]�4�C�I���9���'%K��Ƞ�P�O��C�	>	DEr�A�3vv.E3�d��C䉯�y�G�"� �ò�B�	�v�^�x�-MP�Z$��,8�C��Z�^	#�i��V�b���a�FC�ɬ4�-%�� n|V5pm|�JC䉇��D��O�d.9*GR�;8C�I�=]2A``���}$�9.��l:B�I40;�a���˧�� ��,�#B0B�ɍm�6�hQ��=B���C'�OR�2B䉴%ظT.�"i�|h�N�Z��B�I�{�Bd��Ʒ�Z|�%�	G/�B�	�w,�噗/ٗ8�h1vf�
��B��=q��i$*L�>$cb�R!n��B�IM�`QWD�B)&�� �B \C�I�F���$Z2����BtC�)� Bٻ�	�@����m���~��"OBx+��Нr��LY�M��wȊHy�"O�X:���9{�u�E��pbb}"O�d�獏�VOJ,�o_:1S&5Z""OHDZ��>OY((�6��3*n$�"Op���H������bǸx�X�"O��BC�T��Q2�*ŏWh�,��"O�|+�l_��Ҡ��e3jӂ"O���bk�=",:�C�-��{6<�"O�@��bX����K��F����"O�ȘǦа_�ʁ��@«��ܣ�"O���ϓ2�Re뗏N����"O̽A��ʙ�b�
�/5~�^��U"O�xP5��")\��#�E.o�$(�"O��RӋY�]�"U��N#!x�dB�"O�U��K T����l�T1� "O�ٻU��0��KafN"s��q�"O�hb�	Ab����wRt@�"O�H�j��J"4@��,+�l���"O�$$�3r�P�'�֚E��D"Ox�cM��d���ǟ�4���!"O|��� �}a4���f��6��Q�G"O���$��3�nD��0R�����"OTk��Q@��굋\�4��嚱"O�y��j@;��\9�	p����"Ov�;��`��� �B�>��E"On`�A�% ~�����MSz���"O��pʔ|�R`��M;K��4"O:!{�T05��I�fڣh!z\c�"O�,�5 W�0�j�Ę�30PI�"O(� g�٥(Q^X[��P�X�ِ�"O��+6�߱ ߌ�Qr�T�9��Jg"O��㕭�*`�q&�ɢǮ�X�"On�� 
 <y���9������2"Or�1D ~����DN��X"O��cb�T�fX2'�ɪ.����"Ojœ̓,+����RĈ:Q�"�+5"O�}�$[3p���b�H!q��ze"O"���R�r�
P�g�\��|��"OySB��(S�*�{ �U�ST!��"O�92�Գ8�����QN�$" "O|
��4d��01� l�6I+�"O�؊�'0��u�g�ŘB�jو"OdJ����n�*�bRUm�1�"O���РDJT���ѽ:_U�A"O�ᐫI�
�4��:XNx��"O|5���K�@Ϭi�n�7 A<U0"O�)p�ɩ`]�e�tΏ/����"OȘB�ȑS�d��%�j��{�"O�e�W��I��p�&*[���4�`"Ob�T�̯^I�y��Ȭ)��H��"O�u���M"e# ��T͙���՛�"OF(�4DW�A�
0�Ԭ�8T�=�"O�)���
sNR-���&~i�� "O�E���t`�I��'A�}j���"Oε�(V�_OX= GD�!b�X��"O�������lh�#�<W�8�U"O��8"��za� ��L�,���qs"O�}3�kŔZbh8��JeO��{�"O�YA���)\� ��^f�"O�P�r���E�tt3�5d��h�"OH,��O�9AF�����{o4���"OP�F�J�����N�9|t�e"O��Q�A��i�J��1Xy��"O� ����"�C������
 U"O��+�?+i��!�X �X�i�"O��a��.Ap�#�G
3`��%I�"OZ���F<�Dg�-S�5��"O��⃍�D�|��OZ9`. ��&"O�Y:�̏�<ڀ�cE���nJ��"ObIs�����z�M��!��	+U"O�<۴A͍eRN`9S�E�0��r�"O�4m��Tݨ��+L�(ي���"Op��#���Ar�P�a1�i+"OL���䍸2b~�q%�O�f�:�"O��J���=_t�"F��z�[�"O���#��-4'���“0/ɖ(��"OZ%*�l׎8u�H8���%;�p���"O���w�}�U�Ff���"O������Ba݉e�֔��"Ol�*�9D}.3��Z�Bh+�"O��#!��@"@ȉ�h��b'�IQS"OX0�co��v��٠'X~���8�"O�u�s�X�V��R�S3q��0bv"Ov$�BΦF�"��̈��I*F"O��8dA@RaZ-S4T X"O !�� �?^�P�J۴>D�lQ�"O���%�	S���N�'�p�"O�8�r�j��5ZQ�ڈQ*����"O����,ɋ2@�]C2+G7!PT�1"O:u�A�ܦ
����W�}e|�A"O��
C��hҪ$��c2�v��"O��s�G�|D���c;KͲ��$"Oez�.ű%���YǡA=zД�Kt"O"=�0���~
���N�-����"O�\K��=3�v�xa�U/(I ��"O�uԇ��X.&�9ŉ,<8���"OX�S��j� x�+\FH���"O��Wm�o��`Sa�}�L��0"OBx8���/�L��tHO�`���Т"O(4�Wj<)�\�t'��p�H�K�"O�	������)�� MNj)q"O��(��WB뇅ǨEІ  e"O|<@�;#؂�d�<n����"O����bG�%������8�r'"O [�)gF���òY�,��"O,�	Bݞd�B,�#��J���"O(��Qo�8TA�UY����G��M��"O�U�2��\Y*����o�M��"O<� 	 b�4[��[��@��"O�p�3
�5P�ᨰ��,�\t��"OH` &�
���xQC�4"�P�P"O���p���bs��7/�L]�"Oz�H��S�y��aE��"'4�p"O��b$�52��-�vE��th��r1"O41����"k>z�� r�(�"O�`��� EV�q[4��|�($��"O�1��-�3N<�� ؒMtdi�W"O��j�	{P����(to��f"O������8sB�̉c��"C��Jr"O�3��rO�A�c��D���"OJ$�R�̴N�D�Z�cH}�Dps�"O�l ��S�-��(EH�F���"O���POR�j� ���TE�!�"O�{֌�>�n�%��c���ʣ"O,y� � 9�ZD��a�rU�Pa"O&�ৄ�/�<m���B����"O�eS�A�cx�����6��-+�"O� �l��j��IX���&`�d�"O������F��4x��L� T�"O����8.:����!m����"O��S&'P)#�� wJ�w���{�"OH�Zv�@B��ڳI�-uqЅ�"OH�z��#��2T�&5�4��"ODQї�G�S�š1nD<V *��E"O�<k"���@����bތ<`"O((�wPצ���Q3��1�"O��8��
z��]5x����"O�M��44�X��I�d��i"O�08��Cr���(C�b ��"O���� �1(NҌ�������#"O6�ybd>7=nl��
0{},9�b"OP�2E�Z�Ov=�Cɘv��"OHt���0n�	���I�
�Pɛ�"O�xQ�q�V�0�(�~�Ȧ"O�pa͑�0�h�(�����L�8�"O����:��e��<	s|a"O�Y�A�=�z-��dRl<��"Oq�h�^n$u�p�����"OЉ�(P��j�Z�a�+�4!�"OV%!�&щ�~�����h"ȑ��"O��;1L��s��IJc �\� z�"O�e�2��RUn1!��F
���'"Oj���Z�X��pm?|���`o�<�πc��q�E��2���x$.�m�<��(ڿp��J�a�M�*�òBOk�<���KN|PQ��L*Px����Ta�<1S�G02!d�\� .�:���T�<�Dç6t�u3�+3���� �][�<�Ag��A`7��?�`)��.��<i�ꒋdך�q�A��S������z�<1r���d��,9G�K?����hVx�<����$h�uKɼgc���lBk�<ieF�,oR>!x��Á+z:�y�@�g�<aB�W�x���6��ִtp�{�<iv��"NuBT��/?�l\�%z�<�ꄡ,~m���6L�NPAB�t�<��*CD6q��hA�RBv|+���r�<����+�jEx��ўw?؀QDJOE�<��!˰q7�UBE�����ӳF�<�f`� @  ��   �  B  �  �  �)  5  Q@  �K  3W  Ob  �m  zx  �~  ��  �  &�  o�  ��  ��  >�  ��  ��  ��  ��  g�  ��  �  x�  ��  �  R�  '�  � 8
 � I �# �+ �5 �< C XI �O %P  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4��'d��-1fA�r#
<���`@�4��T�ȓ=�b���
�8s���>h�D|���P|�Ң��)O'�Y� HY"3�8B�I�q���j i�3D���"�W�! B��2��=�KV,!X�IR�d�Wp\C�)� vd;c�OG��A��Y48�(��"O�H�c_�ev�|��jͳU�z��s"O��c��.N#8�g�ÌO���HA"O��B%��,V��Q���ب��`
�"O����;���o�et�I�C"O���s&�;����V_�E9��'Rc��a�C6e�h1�&�FQ*���d6D���P<�ب���p�$�s�	9��M����H�W`���m+(�$�۴k8�O>�	in@��B��4&	�e��Lq�0H��O��Ip�V�US�`U��d���I�<y%�5�S�{j(��R��16�����@��C�I�G�|��+�Ui��Q'!J�
R�C�ɫXe	Q%�
�Øq�!��X��C�	3H��H�& G�C�& �k�HXC�	'd"�q�H� �c1k�#}rC�I@Q(`�?n�!9�
�^�fC��/V!�Y9f�7Td�(z��˦SN���D�>�a��$��d�!��X���x�ŐA�<�֊��Pی�z􂒿Ha�����z�'�?��&���"��A�a�P���5D���&�P�4���P CP�j5a��>D�\��%Ϗz�\逬�=7W�0@�*=D�p@����`z��]�\d��SV�/D���qfܪ6�Q9�ܩ���/,D� �E��k;��lT �L��6D���hA�| ��%`Πn�n��g(D�(C�� O�N�x�$��w�`��%D����oS2sn��b��vH�)�uI$D�HZ��O�ct��8~s2�`�#D�HP���;>�5� �f(���b D�$���� ٔ�9�lB,fr��<�!�䘛B����qꚩU�F1R�N�<>�!��E�f[�QiVI�j`A1�>v�!��NH"$$�ǩB>��J���!��.f�=2v��;>$�s���,�!�H{����$;X-���P�!����������~��JZM�!�\� ���XU�q�X�:T!�Ą;6����V�$��tJ�dӑX�!��Y.5��pbԭ��P�D����W�z!��U�h���0�TU�0ԃ�#���!򄌵�Z��aÝ/u="�2&�G:n�!�B.Cż����F+8>YPeφ$�!򄘖lU������& ���H�Q�!�D΍h,r��7Mi���o~!�d��Dp�<S���K�h9�DJO�Pm!��(*����p��L��T�PFK�N~!���:ct$+Ǥ�&d���f��Ev!�G�k�f-�Ć&1�<��wd�2~X!򤄵a�HK �۳tH� �`�i�!�F�N�\�F	�qKz�s �΃l�!��G.�M����f9d�@��>�!�ў_ �i�+�[ּ%*��̩1�!�$�+C3�(2�G��	`�H���!�d�X����[	�гu�_1?!�ܱO_
i	�k�Z#(p��
f !�$�32�tj�رWD��jS#!�� �"a�k�d��r��O�!��Fi�`�`f��7$9�5�0_k!�E }�z�͜��)��Į$�!�d�p���*N�\�&l�V��~9!�dOm�$��#Ɔ
�p�֏Ӻ�!��j���1�Y:zF
���#r!�� $�EbW�Sgl�V��k�"OR	�e��	dȐ�fD����E"OH��&�[:<�n��w� r~zxɁ"OZJal:I܄���� ~����"Oz��FaJ�W8��teo�%��'|"�'���'���'Y��'er�'r�<1`��$/jl��¿.�0��'�"�'���'���'9b�'��'��-q7�V9EHH��"��@�s�'�B�'�"�'���'R�'���'��0���H.]�E�|�f�p��'v�'�B�':2�'b�'���')>L���i��}U�93>�@��'XB�'��'���'�2�'4��'VzT�w� _b�rc�_5$��\�S�'("�'���'���'I�'���'&�AYs��;={dQ��"	�:����'�b�'[��'�B�'Mb�'��'��\x��ټ**<�b��7eӸ�j��'%��'oR�'O��'b�'���'��.N`����R�
�1���'��'���'���'gr�' �'���។B����$(��6�����'�'�"�'���'�B�'�B�'d5r�Ɂ$�z��tf��fΖѺ@�'���'\��'��'��'���'�](��LA*��\(0iz��'v�'UR�'�2�'
��':2�'xV�s���3%��ҖE�!t�8	s��'���'""�'���'�bno���$�OtDB�����1�������dy��'J�)�3?��i#��wߛ=�Xf��^1��O	��������?��<��v_$#C�d�JX(%s��'R&C)�����ţ����~b���?<�6h�����gHӈ��'�rX��E��y���Bh�5s԰�/�;
��nZ�'
c�������y�)��y���kDaQ�1����(B�f���'�Ĩ>�|�ꎳ�Mk�'-�}q#��~Lm�@�q���<�'�4�$��hO��Ot8���Q�#S>,����2-�&<O˓��^q�v̄�'��аD)e߾e�(���f�dBY}��'�B9O��F;�(����% 0�vEQ��%�'F��V'dK���^̟`K��'Fv���/O�x����ںF����sT�@�'���9O���F* �i"8Txg�X~�Ӣ6ObPl1�n����4���׮@�5$�@f�]/ql�[�5O��D�O���,W8�7�1?��O�T��^�7�|h��ǍC���3S�œd'TlqK>9+O��O^���O����O�}�$ʔwI>��v�J1�T��<q5�i}��a�'���'��
=p#�AI���0���r/b���B}��'�2�|���N��3J������ܫ$��yA�����i �ʓ�\Ȼ�ͼ��$�T�'���B*�%��}����+iq�� �'��'�����[���ߴ��R��^qҽ�rg���	�TQ	��h��Vp�6���]}��'xr�'�<�T-&ʂ��E,	u��2���m��ƒ�Љ2�<��d�i������Z!&Sn�+���)~��6O����Ob���O����OF�?i�wk�/|
	:���|^P�D� Fy��'r7Mo�I�O� oZB��/� %b��j0��[��U(u�&���I�擣E�l�@~ҋ�3Ha���ah�1¼<Ri�+I�޹�fGI�40�|RW�����	ڟ�{Ѕ�H_��z7��}��pK�*�����	jy�.q�e�P��OZ�d�O�˧;�
�q��P���X!	Rc�0?��_�������$��X�"��&�?���+ԚLN��EjY�4G��������4�����gа�OX�)�1(�$jKԂ
i DRt �O����O���O1�j˓:��X�bN(q�P.�[�f ɂK]I�2� ��'�҂f�d�x��O*�$J�L��%���I- �� �%5Y��D�O�����m�b�}	��Bk(�S�Db(�1 �"j�:ES�����IXy�'��'8B�'�BT>}j�%D�	�˗��sIt5����M��H !�?i���?ь��t��.߂��4`̇�;�d|�Wc��4[2�D�Ox�O1�<��Fl�v�	Rʘ]��%(얍9a��Ou��5Y 8���O��O ��?��c�0���F p���WaI�&�N���?���?�(O9nZF�v��Iǟp�	d��i�̯T�R9�1����E�?Y�Q����W�p����mbb��ʛ7$��'�6��Ǎ$\H`����̟`0�'R�$�q��</��K��������'���'���'j�>]�ɬHXQ�Fo��zT�V�:�����M���ʶ�?�� ��V�4�p�cC�3C� ����E�bj�>OT��Of�dL6:�j6�*?��l����I�xSҥ���
�D��EL�$�O>/O�	�Oz��O ��OD|�&%�Roh�yg�Ϡ�H<ж�<) �igF�K�'��'>�O� ��Y�*�hF�8T߰�[��ʱ*�|ꓐ?�����Ş��sj4��&�ɿ#C�� �W��޴"�剼F��jp�O��Ov�"����f���Bje�ǀ��P�����?����?����?a/O�1mښ/F �	�;�~m�E@�5��81t嘕���	.�ML>�'(����X�'<yhf�IV�K�L�;��>"7ش��4�yR�'ubhӇ���?�a�Y������� ސ�S,�<J,�����3�hK3?O����O��d�O��D�O<�?IdA�g1�l귅72��qJ�Tyr�'�H6���=��I�O��oZ{�ɵb� 4sr�I�|��aa��j��L'�T�	�
�&|n�Z~R��!��IRH�*lX�b�l�4@��Xө��@�Җ|�Y���|��� ��K�{b:��B��##��̉D��<�I\y"$zӮx��E�O��d�O��'$dȨ*C��$���B�g������r�O���OΒO�S	���Ї)P���[6c��yk�����0�>9lڭ��4����'��'O��[ቚ5�jp´H5n����r�'�B�'�����O���M3d皓,*�p�A� N��� ��
O�R8Q���?ӹi�O i�'�W�� aX"vJ�Y��
F�C*��	ӟ�p����A�'M@֩�S*+O��ң"v.������ �0O�ʓ�?A��?����?	���IX)Ϥ)�E̙9O�6�z��)l��o��4Ȋ)�Iǟ���r�ǟ|����7Ƌ�=��aCͥ�U"�/���?����4a��k}��9O�����T,32����ǆo�q��<)U��K6��D�8����$�O*�D�qr����He.���X�{�h���O��$�O�o����G%2B��'�Z�+�iS7*t�[��R����R����^}��'�2�|��]�w����_(��Y��16>4)3��k�$c>MZV�O��$[s�:i�֠�27P1���9����O"���O0��?�'�?���ɭA��X"F��H��Qk�#ƛ�?���i l�R�'n�Fo�d��]*/F��4,#S�΄(��,%/���󟰔'�jmJ�iC�	�2��B��O*F@�����Ϥ�k@e&)���T�Lv�Ify��'r�'���'�R��3n��p���� {�v@���XP�2�McB���?����?����-��0c�D���ɬqV�h󔌎�U/\��?�����S�'rZ�\��So�Fx;!���w�*��ʠ�M�aY�@����%|P��;�$�<�V !�
2$��uh���fO�?9��?����?ͧ��ʦ��!���(p'���r/�}Q�f-�26�[��4��'M���?*O 5�"C�2,��q��[�P�5�̙B]>6�)?�B��0E���)��¿�N��}����(?JK�! �F����IԟT��ܟ���_�'H���R�M�iP�U��Ǌ�V\���?��r8��	Ё����' �6�<�d�I����uXz��Un��~rf�Oz�d�O���1�7'?ѱC�K^�#ť!l���C϶y�t���E��|$�`���D�'�R�'�J ���3����b�j�tt���'C�X���۴,�I���?�����W�}�0��S�`�T�i�jS:(�	��d�O��2��?ݨ�n֘l'x���[L9�
��*�fa�Ƈې�N��|���Or�(I>��ѢH-.���n�g�Z�Ib&<�?i��?9���?�|�.Ol�'W")�&�ɦ(00�Wg�]���js�ßh�ɖ�Mk��J�>q����;�GZ�6�ؐ�^at�,O�;�@r��cx�; �˔by�-��S����vaO�*�@��D��y�[����՟8�I� ��my�O@^a:��V�~
�-(���%����}�L���O����O�����$����]�q}n5�F�ԁ.hذtg�-0PT�Iӟ$�b>a��-���!�9s<  U�<cb(0��I�5������5`#��O��SK>i+O�)�O4A#'�ӵf<r�aG�J��4"`�O��O���<�u�i��I�$�'er�'h�1�e���^t�s��m\85	���f}b�'�R�|��Z�j1	��ڂ@��P3T������%�l�x!�l�:L$?�R��O���ɳ�r�'��qtX����/�$�O<���O(�� ڧ�?)Gz��`� n@�J<���DS��?1��i�da3�'Ub�nӊ���s!��!Y
���)�b>*�Z��ȟ�	ޟp�D�����'zJ�Ǯ��?��F�ȟ0B8�#��B�Bm��(R�wE�'��)�3��!;>1ڲ�U�{��<���6���B�����>B�'�r�I�+���#�WF��կɣ_��e�'���'Oɧ�O�!K��ݜa�ԑ2��]��G��^��5Z�|��+�A2�����3�Ha bF��zw���#1�a|h��l�*�O���s�W-�$ f�}Vd-j ��O��nD�Y�����H�I���jcd ��IH�E	4 ��
9nPn�G~"�F<<���ӄ?$�O�W%ܑ�|e��"�8u ����y��'4b�'A��'�b�iĵ4�H�)��Z5�.�0��)*VL�D�O��DܦA0��j>��I	�M3M>i��Ę��t����0-���O�����?���|�Vf�.�M�O�23f�7&����pE�)*�g]${H���'��'���������<�ID�pK��^3sV�����'}v��	�d�'�6��rm2��?1/�t�X��9.wBi���V���	8#��H�O.�D�O��O��q�v�K�!��/p�N%�����El8mZ���4��)��'�'�TQ�E��M� 䁣*��I�`��#�'i��'�����O���?�M����.8O�� q���)Ƕh�7K���P����?a�i��O��'}@Z�t��8�%�O8j��l a��'|<P�i"��/.Nf�П �S�? �lk��:�PvhX�66���?On��?Y��?9���?�����2S��䍘�J��z� ���)n�on��I����	}�s�(k����Eo
�R�DA�!^&l7& ��F9�?)���S�'G�
���4�y�Y�'@���Q\/XR`�v���y�������������Ot��C�l,��Pul�*0t��0�V�z�v�D�O����O&˓eu���:�"�'0RL��d�;��Y2[��9tAЙH��O��'���'S�'��M��A�2Y6��9BnW�0��S�On��rD@�s{�7M-�>����O#��J+<sTQp- K}��c&�O<�D�O����O��}:����iR�G�4�a %� �7t���y!��Y����'�67m?�i��s�H:`����ud͍�P�ʷ�t�$��ӟ����{�4�nZI~�#>�����C�`�r�6�R,�B�׈,��L2L>�*O��O��D�O,���O��7�?4`��i�Q���ʱ<���i�q���'���'�kg��c��h�G�K�ѻ��Op}��'���|��ԉ�:P��]�D_�r�!)`
I
t��]R�i� ʓSHҠ{en��$%���'��1�S�,��ۧB��oNd� �'���'2����Z���ܴo�:P@�k�@��W��n��$(�0:��( �X,���d�J}�'4��'�<��b��	�T v��@�Ef	:˛Ɨ��uԢ�Q>�D9C�
�Ba� �ũ�;h��������4��͟����O�$�ARC��a-:�BU	T�{�@����'6�'��7m�3R����O�ili�T̈|�"�R�fUG�݋�I$�T�����:�	n�t~B'"<�h�"�^O(&B�!j����˟���|�R���ڟ��I؟�hڦ.�>���%26T`�e*	ğH�	Vy�Ө�ͺ<�����)\ �(�����@��������	�����O��'�|R�"D�(��ǆ�r�Y�`��'/���X@Ď���4������9���Oi��p��ݡ��߼�`BԨ�O:�D�O��$�O1��˓[Z��ĝ2�9�D{<�����81y�@"c�'{2,iӼ��p�O2��O�\�%�HQ�ܘ�*1���>�D�O�P�T�s�F�i��(��?9�'1���耞�����a�ip�'�������T��ʟ��V����{��``�K��9��2RA�`�6-�9s�|���O2�d9����M�; $0��cpx���6*���R��?)N>�|
b��2�M�'�pA!�'(O�ҽz�oU�lp��P�'~���	�j?�I>�,Op��OT�(Q���fx�i'ˍ+o�b���F�OJ���O��ĭ<�$�i�t�5�'h��'���y ��,q^�q���Z�R�R����K}�'��O��귩���p D��t� �����`��?a;`U;P �G�=`> �՟���B0��aZ��̩�t0�Bi�����I����I㟘G��'(N�!�M��4�y5��Ȁ�1C�'P6핎J�,�D�O��n�B�Ӽ�oBBǀ�Ȁ*ä8{�IW��<!���?���Y��iܴ��D�&r��a�O����"��<}�bPp�n�0D�<D��|�^���I͟��	��	�̰�̓2T�p��Ɠ?����R�ZyҪoӬ�Z���O����O,�?�aF��T[P�q�i�ZHE���d�O��� ��i^�XL��h!���|��L���٪"diz��r�$��'�Vx@j�j?aM>1-O����ƌ��h2į�5[����)�O^���Od�d�O�I�<��i��T�'i"�۱bP({��(�'�$DY��'�7�9�ɉ��D�O���OPAG+z� �3���_=P��{�H6�2?@��U���?���1+ENs�Q��eUV�<P��lu���Iџ��I�t�IYy���G͒o�8���* {4���
�C��'RDk�T�`h�<Q��iJ�'�h���ǵs&��^<p��C�y��'�	m�<Ao�e~r�Ƅzv8�Qb�6�9 ��/BѢ'��|��|W���?9�+܋3��P'j�1$YfI���AJ�'�~6흉/���?�-��ĂWO�e�j���X�I&h�Ɨ�ɭO��$�O0�O��?l}�m1�h̘]�(x�wJ�����փ\*<���o��4�~�q�'_�'��5P�"��Xk>̑䊃�{X���'2��'�2���O��	5�M[@��&m�,L
gOי8���/jF~�#�@S�������M����>��Pmb5	!c���,y�ㄇ�q;\I���?�5(��M��OP��c�4��I?u{���>R�\[v��5~}p�"��m���'���'���'�R�'���!%
t�0%˅�����@(��RشD�ֽ����?i��䧹?���y��/{u� 9Hj�δk�+�${R�'ɧ�O~,�;V�i��$ŊB[U��+�1!��E`����t��P5��3�s��O���|Z��5XѠ
,Ka��Zb��p6�����?����?-O�4m�^�X����\��*"0
��î�2QzDjG/
r��?��U����ȟp&���G��|�TB��~<N�Pl*?��
Z%)J��ش��O(P����?�aع�D<+�٘pu(t���?I��?Y��?�����OV���p�\�k��ɑ��@��O�-m�IV8�Iܟ`�ݴ���yW �=o���$�qR��`	:�y��'B��'L	��i��	��:�I�ޟ� ��&�'W�$@P�n7:gG �Ķ<�'�?����?���?w��@u�$����1e�j�'@����Φ9�K������t'?��I�5%�l �ˈ��r�@�JA�A;�a�O����O�O1�*a�|�X�%�+�8`�V�7#5|7??逡^�ߊ��@��My� {J�؄�S�U�eJ��P2�'��'��Ob�I�M��fB��?yQ��<!��A�/_%LDxk���?9d�i*�O��'���'*₎�V,.``!��.Ȝ-Q�oH��X4H�ic�	�!�:�s�O�q�X�Ψ&��� �ƌ�D�4�2��^���O��d�O8�$�O���)��1�uzV�Y3�L�G
͔%bT�I��	��M[�g	�|��!�&�|�H2.�
,˥��5t�r4��愥9��'����$�Y4����,�Ə��%=\$��͊
h��I��
�o
�S��'׬�$�䗧�d�'��'א�3��F�my>5㣅\�.d�!A�'��U�Ta�4^�n�/O��D�|�" �04��Dh5�˞@2x{��A~Ⅴ>y���?aK>�O�T����ϟ �� K��^A�L-l$P@�����4��L��=ub�d �W\��9f���p�D:���c�I�
���O����O(�4�RL�ckՅ kF�N��FeW�3�L٠�A�&o�@Xb1'5S`��0�Z�@!ٴ�䓎?R���	3x<�
�HGT�\�R,��n��I���z	C�%��?y��;�H��y+�sܭ!�D F�l���Ϣ�y�P�H��ҟ4��ǟ�������O͔�����ub�s&6 %|���Oq���Y�!�O���O�����ZΦ�]�t��I��X;&�� �T�v�R�����'�b>IPc�RϦ%�#v6A���^)U�倴�/]��͓ZZX��Ŏ�O���H>�-O,�$�O"�3���	R_V�#��|�r����Ov���O��$�<Q`�ir �q�'���'�+�
o���MCb1����DXV}��'��|Ț�@�<	�l�7�^�G�
���ِB"���;<���艱�<��ǬMyځ����� h�C M,D���O"�$�O.�� �'�?�'P-U���׏�����֞�?�4�i���`��' ��n�6��]�H
�l)�M˶iC�.I~t(��3O��d�Oj�D�3j�6M"?�e�K4��]�V,(Rʍ1
�� cu����v4&��'�џ�rfR�w�TXfaY��p�$?9�i<Na���'���'T��*vl��B��@�ƀI	V褈2A�k}b�'��|����2G���Sh��6�8`W�gq���eL#��	!\w�����'�,&���'Zđ�A�eah����G�c��@�'���'>����4]�<��4 �Y��o�>� �����%�8<�\�j4����hy�4��'�P��?����?����,@aq��a˴b�>J�FZ+^>4��4��~��i���)�"�k�9���Q�J�k~x�r�9O����O����O��$�O��?(W`_�?����%��a�6�Yd�U�����Ο�ܴN+0�Χ�?)�ic�'4��@��N�gb���-�J�(�d�|��'��O�R�:��i��I�.`�ҕLL-2t���[�f`S���]��D)���<Y���?i���?)�э�:��w�_=q���S�M�?q����d�AZ�Fß ������O�"|��lD�����#��o���
�OZ$�'("�'�ɧ�I�=v8c��M,��U��li�6��6!
�o�ԑ➟��^��ŝt�8(B�V
g���r瘢I��,�	� ��ҟ��)��Zy2m� �"k�57[���B֧IJ�$s$�ژ��d�O�`n�P��\��	՟��%H45�\V es�� r;~˓r�*X ߴ����p.<:��uY�ʓ��$�aa�
u2��#�ߔxz�����OL�d�O.���O�$�|�v���EPL�����'��X#��p���D�3�	؟l'?9�	��Mϻ`���>Y@�R�ϊ�"Z������O�P|���iW�$A{ �e�##T�W+N)�����^�$2\�Q�z��OV��?a�P�tqEE˅424��F�?�������?����?i+OtQl�kH��۟���
*�����
/.����׸X�h��?�`[���	ϟ4&���b�9j���ܠo�Mf9?Y���2�´�ߴ՘Oi:����?Yu�ܚqxZ���NL�hGx�ҍV(�?����?A���?�����OV���3.혝���]�䥱��O@9n�X����I��`#۴���yG��0XG�X�.ܗQ6~\���� �yr�'�B�'��T��i��i�5ӧ�T�?%�5���#�)YUc��@���z�.U�@��'�������۟T��쟰�	�y Y��	
����!��x���'|7-�6@�˓�?I~:����#�D"��q �GS�V�i6_� �	Y�S�'Ք���	�8�k&�IH�H �̎�i�:��)O"Y #���?��&.�ĩ<q �
1�qS��`�����M�?���?����?�'��D��MJ����9�ÕA�괯�)T;�U��bڟ�"�4��'\듓?�*Ox]��/ƻ7><4yũ�1V���
��6�+?v.M<[�$�I���'ܿ#RiA��zuqB�FbD�%"��<!��?���?����?ы�㋟q�a�7oU5�lが/\2B�'�R�b�p�0�;��� ��$�P9V@�	Q��	�dG
Q)\8��T�	��i>�K��ۦ��'V�U�� t+����k&�kA��!o#���	U1�?��G"�ĵ<ͧ�?	���?9��_����Ǉ�LҸ90� :�?Y�����̦1�k��\����O�a�M�;�n���.پw��U[�ON��'B���?���F�Rp1w�S�|�,��GE+<��ax"��s�E����������|r�D���pI�zfB������$��'���' ��S�y�4��}�DA���e��`���L��0ꕷ��¦�?��P����*v�p��ۘGb�`�.��-�IΟ�bŅQզ�u�۝F��ly�j�2jeĵ���(T��iӤT��ybV�X�	ǟ`��͟�����O�$�������	��0�����Mj�Ia�O����Oܓ������]�!��M�0�r�"AdE j,������'�b>)���ܦ�)h�-Zģ�#.���B�
5`ΓD<N=jb��O4d�J>A*O���O�qsb�L�9��
�A�]��)���Oj�$�O��Ĺ<!�ie�S��'�b�'J�Ř�ƘV��)0$�?ED�hB���VT}��'W��|BEW�xs����ȍv�����d���ב�R�� �g��c>�@��O��$�+uh�\���L� 玱xgE�u���$�O���O��5�I�O�͠���O �А�S	讥�����l��CCh�OV�m�Ea����ԟ(��4�䓩?�;)�(�� E���刨o̢q��?����?ɱ�І�MS�'*$KQ՜Q�E2���4� ���a'�W5 +
d���|2_���I͟��I�l�	ϟ��"%��L{fo�,Z&0���ty�q�H�#5!�O���O����D��ؖ��i��d�;���/�e}��'�|��D�ڂ,�|PX3eU�n�F�q��?x��u!��i6�]~��'.��H%���'�� �� �G1nL�A�F�tn�ѳ�'J"�'����V����4L"r���TX�*��Y9\�����q$0J��=z���Q_}2�'���'~Y�ː�K����Ly�X ��K�<śv���1�F����t������'K�AQY�� ��
b3m|�P�I���� �������V*J@�"&��?mF,�c�Я���O�lZ[�|���(ݴ��"�r�sQND*<�0U	���2�� aJ>	��?ͧ\�4sش���H��j�K����E	X�w��B��	�c���?	�� �D�<�'�?����?� ��!1�  ���
M��y&L�?����d���1�ޟ���� �O�j���Ĕ��bHSaI�e{u@�O���'�'Mɧ�I�7c�: ۇH=&�|�S�?�|3T���]�Z6M�}y�O%�����u
��Y�i�>��e�BB�u�mh���?����?q�S�'��d�Ҧ-(EֽDgjhQ�g[�q�|� @݈څQ��l��/�M���d�>��|l}	�
�:o?�iF�[6B�4�����?	$�R��M��OιB�N���N?͠4(H=W�}�V�ʿ"̢��� o�@�'�R�'��'4"�'R��<v�q!P7�Pa�CM���ٴ\�����?����'�?yհ�y7�x�B�[fA�%S��(#"*��'ɧ�O�lxh��i4�P&K��0��iN����r��PA�D3K���'7�'g�͟|�ɯ,:ZP�`R��� Q��_V\���ӟ���ɟ��'~�6�F>H}J��?Q�+@?����x��H�iV0��'>��?����e~�k�L	o�9k�W��� �'��0r��:wa������������'jq	CV)>����sPJ���'��'{��'8�>A�I�0y�|j��f�T�{W�H��h�	��M����*�?��f���4���	�$DXR#�&�����=O �D�<��k��M��O@0�ө^���IݡkϞ��c�o|k�OG*nF�O ��?q��?	���?�Izz�RSgFq�]�G�U�E����.O�}m� b��!�'f����'���{�b4;n��p�A�C�D��g�>q���?IO>�|
Rl��H>�dJ��S�n�}B%���N��i�O~~�J �����|h�'��ɫ&�~���$$��D��t%��	�����ʟ��i>�'�7���*]V�$�2,jlC�/�P��O,Fv��Y�?�Y����HyR,�1Lˁ˔�ۧ���s@�9�kK��MS�O�)"�����F*�	��BY����0)U��
Jh�I6O\���ON�d�O"�d�O��?P�b�"ʌ���`]>^��)@���L�Iʟ4��4W� �̧�?���i�1OPݡ�֥^ �i��J�'V"H��|��'�O�֤0��i��	TYh��-�2�����؜*c|8�G�y��D/�Ħ<ͧ�?��?1�@�bA!w�G00����?����dA�my!�Qyr�';�#���9�E_?5yXQ!�HP2B���m�Iڟ�?�OʮɲA��WX��Cv�
�C0V$���!�$4�u"
8T�i>Q���'�P�$�D�q��nb���&�9b�asŉ�͟����������b>�' �6�֥u����a��b�TMS�F<��5��O$��A˦q�?�R���I�Yqd�Q�h���43p`�EP>�Iٟ<k�HӦ��'g�h����?5����DF8\���䞹e�JI�0Oh��?I���?����?����ؿ3�L�	b�H,�%����>���n�	E�@��	����q�S���a������Z���&!�+�P���I��?����S�'5���ߴ�y
� lH4��a�$�z�dų3N��4O���䪀-�?ic�4�Ġ<ͧ�?c$�+)�B	�C��c��a��Ϻ�?���?a���������-�H��ҟPi���#R�r5�>X�첐�PV�$�����q��䱉�0���㧅��<�a��A��##��qI~�&A�O��9����pQQ�����ѱSy`�q�g�O�D�OP��OX�}j�aQ�uH1��8&��)⁞�7~�yI��ӛ����>A��'1�6#�i�Y%��M��*���:3<`膡w���	Sy�n۱eƜ��S���o�t��y���;1�T�n/R�yӋ�'ox �$���'(��'���'���'���PU��Z5���4J�]���]�ܴaѤ�
��?������?9���
�t<��D���ȴ"R�>z���l�?�|�T���~Z��I���~VƝ5H(380ˣEI���D�,;������'�O�˓<F�uI�#Ȝy�L��Kud9"���?1���?��|�,O�-n�$jL����sqdiq`�6E��Щ@�p�I��M�bš>���?ͻB�>m���&Vݠ���X����.���M��Ob}0p&R���T��4�wH��/ѿE�A� �M�.fYӚ'�R�'�r�'x��'u�JQ�և��M�C�C�Il�Ж&�O��D�OJDlڞ�Д�'
�6�%�$��_%��+��zg�����LP1O�Ģ<Y4��(�M;�O �JT�M4aϚ�yUb�3�@��BP��L;�U%T�O�ʓ�?1��?��:%���A��\����F%��;��?Y,O�hn�����@��R��	�Li(5Q�P��AV��.��d�L}R�'M��|ʟ�L�5+֛~��A�$e� ��d�!'ˤt�Bղ2�
L2��S��'�dH&�� ���s�j��A�o�ȁ��ܟD�	��H���b>��'�6�J0(`يQ,����y��S.]���B�O��dB֦Q�?�U�t���5�����s����!:JB��П���hΦe�'@�p�B�\�?M�����a�̓�ZaCRh.nBrm�S7O���?��?���?����)�6L�L�:DK�)=)n<�Ҡ��{q�ln5!�h�R�Z̟D���?�ӂgI֟��Iȟ�ݬ0Tne ���&l�,�qp
=ap�L�I�L&��ßd�ɲ3��m��<Ya&Y�J�)�E�F�Q2���<��+�T=X�������4���A&��# @�+�LQ�eh۔\����O��d�O<����AW�u��	П�;gl�(,����ŨVZ���+E|�x�����Ih��,Li��b��ҫt�P C3�;/��V���"�U2^��O~Zh�O捐��%�t*F�Z $9��FW��9���?���?���h�\�D�D8�R����N�
QB�l��T����C$�Hy�n�Z��]/�ֈj0G��dL؈�ؕ�
�؟�'�a�i�ɍ�uY��O��< קB�O�������Cvc6�Q��[yr�'�b�'=��'"O�6�|���_wS�1�%�[�c��iٴ	,�+O�d/���OL0
�ۉ=���3pn��W�`8�f��b}��'�B�|����*=��	Q��1v��p鳨�O���e��$Q-���!�!�ԓO��w��h�7�U���ˣ!|Z����?���?���|�)O�}�	������
C��zr��/m
tLz!%��Y��$P릱�?��Z���Iܟ0���Yynq��4Ϙd�cG~�!"�������'h@A�N�^�O�W!\7	ĞL�c��)%�2E��dY(�yR�'��UHr#� h��5�Aɏ
l�t ɦ_��I*�M�R�Vv��G}�J�O�u{��	0D�C�
��
B�:���O��4�d`�1�eӠ�j�i�)�/�Qz &�)�|�R�-R�z��Q��iyr�dӰl�-�%��.D��`����d�ڴm�0����?	���IŨM>�ӵ���ru,� z�ɢ��$�O��3��?}i%&Q�M���S�ߐ(�Y�'�N�V81�dF�:;8-�����R؟��$�|"F��oF,��j�u2������x2Ev�:����\�`m�]�"�>L���Ҵ�?V��˓?��&���~}R�'�Z�3�z���)Ҋe�v�Ca�'���L�M����@+�^�i�ɵ<�7H����\��ذy��"����<�(O���D�\�P�S �ٰ5���W�R�Y�6�l�4�d,�'�b������B���x�#�+t�:���&3�����؟�&�b>- �oG¦Γn����C�ͽw�,y#�*� 4AB�ϓ<T\�ۧ띨�P�r�J#W�\4��c�&H���׌��!#�d�L@�r�f$X�L�T� ���l�� g���7�E�Oi�4*��ϥD�^y��ǰF׶��W C�h�Ь�5Ȓ9%-��UNM$��am/����fƶ���
9Z`��M�iHy�R��;z+��A�"3��8���8iP	fÐ52�&݀�I�6��B�[�*4)����^GH�#�'(DEh�ŝ/��=A5F�5^0���V� r�IBACӉh�t����C(r� 1D�D(�(&��*>�� �f*6x���\������M���?	��O�3����2��
��#��Yқf�'�'�r�'4"����!P��� c>�bLԂ��j����'$�P�sӣ��i�O ��� ���+��*��bhY����0�]��4�I6S�q�?��O�֝�Ʉ0m&��EA� @YD4��4���O�'{�n�럈���x�S�����y �Уw�9g��:\m���d�i��'��ؒ��'��'��>� ���a#�vx|��%[j����i+�	��n��D�O4�d�l��'��dT�c�͸n������F�<Q��A�4 �J �b�i�Of�����x|T���&P�Sڐ������E��� �	:8d���OV˓�?��'q6��6�y��c CڐN5�D9�}r�Y
 U�'�B�'u�[�0�A�B	�1p ��8��tO�7�Oh���X}�T����z�i���'@,0J(��7_�fz%#Q
�>ѤE����?)���?9+O�<�6 X	5F����ɒ�
���@��'��I���$� �	��$�W��:ڜ$���n͠$�5�ȁS�&����ԟ8��Iy���"�H�ӂA\�X�0�P�3Vj���fX���Iy��ǟ��������(�컡oMX%TLSW��*2f ��'[��'�P�,����0����O�+�^�fٖl�]'A�ְ�GJզ��	Z��ԟ��IQntb�R��<ZGh�I�&�K���7M�OF���<���Ô&k��@�	�?B���ÒE����J��(�!�͕�ē�?Y�/��}h�B՟�<S��+Mp8�)�ԞH�@�C��iK�I� ����4�?y���?���q��i��jW�2��C����`�`B�}�(�$�O���p�"��nܧ/k�X��܊$D��Iq���y�t8lZ�:�eӨ�D�Ov�$���'�	<�&�d��D�6�;�m��H�jeSٴ�$���	�OJY��d�3�ȥ@���e��h!�LѦ��I����	7.z�92J<�'�?i�'��0#FW�3��݁��@�!�&�k�4�?�K>9�\?�Iݟ��I���0s�P�!�M�ḫR��𫔋�M���m���b�x�Oc�|k�i�p�(�ʅd'F��Q랊]�hO��<Y��?����D��$wz�����}e�/��`��\�ǟ���U��GyZw�z����C)�l{$��C�!Bܴ�?qL>��X?��� ��Qb2�e�kV�� M�,H�-�e����������?����DR�<��GB�@�= �h�)����l������O�D�O�ʓ?*�)`���)ж"��)1T�xX��*O<�7��O �Oz��|����Ӏ;4�!�Q�9'->`k��z�x6��O���?�%΋�����Oz����kl^�O��D�2K�*-����w�мT4�'[�_�����=�Ӻ�V�	�'-�񃳦
�F��I�#j�ʦ9�''i�F$z���O�r�O���h�%@ �A7�mc�*�,\��l�vy��'o�%�=��is�E���l���l_&Q$�r۴Q�\<j��i���'�2�O4O�i7S�����I�=�� ֪� 6�m����	ٟ'���<��s�r4s��ī��(qV��,�H�1�i�"�'�b�9�O���O�I�p����B ��U��m6��OP�O���<���?���T�դ,��ıI���Jg,̍��7��O��$�w�i>	�	E�I�I=�����gװQ��i�9$v\��M<����䓯?!.O\��(C@�5s���4H�-+p��@������<����?�"�'�� 9ix��ݼ^`��#�)5���b߰�'\�V�x�InpJ��'eVⵑ�BN�S4���Y�o�00n������v���?�.O�ͩ��iL�T�2aU�RO�9X�GR���K<�����O���|��W�y�E�Ճv���c�AX|�� ��i��O
�$�<�T��e�	�B��Z1g�7L�]!`��}&7��Obʓ�?�Ѥ�����O��D�kl�(x w(ϛ&�$�Zr`�Q��'L�T��c�.<�Ӻ;խH.b��k���4��l�G��Ҧ�'�8��'sӼ(�O�B�Oj6�
 &<h5��j	v}фE�";d"�m�ğ��I����.���<�(��&E�ީ2�C�)]���2��M�E%���?�������S��I�$<D���M|��|�Bg�#X:��u�Dx����'^��`���2�����H5���b.|�l�$�O��D�v��'����,�ɍ?���4�R�e�%A�@�U�l��4�?!���D�p��O����O�M�c^F�8�R��:7y���`������0h�HO<ͧ�?1I>�;W��Q��h�����u�� '�`��By��'��'
�	.]�R��B�)[1<ѩ�jҐ,8h��d���ē�?	�������` �+���f�);P*t'�i?��|��'k�	ԟxq���x���υ%�l��k�i�� ����ʦ��	؟(�?	����D�0���*	"^ٓ�!D�+^�}��������O����O��<�hEU?5��*	��Do�)p���1G��[s�<�ٴ�?9,O����O��dR�ET�d;}"(�dĄ�A��_�c�R����MS��?�.O��k��r�D�'�R�ON��2�!� .�B��rJ���GA�>���?9��+��$͓�?����?��OB���B�s���ƌ�5�&I	�4��DܛA���mƟ���Ɵ��S�����J-���M�Z��Ui%�(g���A�iQB�'bF��';h��<q��D�ڦ�B%QQ"B�Z4RP�2�M�ֈ�J)���'���'���F�>1.OF�`�$ϸ>jR���K��'�H��n���q��b���Iɟ���^���?y2��!]�F�kN)s,X��F΢h��'�r�'*r�Q���>i/O��D���c��[�J��HG��W]�s�|����<�s,J�<�O���'&��;� 
&/�v��-��_K������i�R�;�드��O��?��i�)34H�'(h���V˙�h�,u�'0]+�'�B�'���'8�\�سӗm���{��̲a�� �ȩ.2�®O���?�-O��d�O��Č�|�IF(��rD ����r{��63OX�D�O|���O����<ar*��t'�)�=~�.�cQ.���'�@�I�v_���Izyb�'���'��b�'��K��� *��$xdH��U��4��'b���$�OL���O��h׌8r�Y?��i��PE�+O�`�A��*�ޘJ!msӊ��<I���?!��\UbI�O�����@@�%�b�WL�
�mΟ��Iqy�l�~� ��?a����0i��g# ��S��G� (�N��a��ޟ<�	�x*��d�ȕ'�"ҟTK���%9��4�Ĺ ʆ�	7�iH剰?k�MJ�4�?��?���5��i�{��ڿ'��[�U�}R|Mp��vӐ���O,���(�'�q�@e3� 2��s$׉�Dyҥ�i�bىba�R���Ov���,�'剿
���"Y�Z�YF-��F���aش+�l������OD�_ FG�}S�CJ|^�ī�*,��7��O����O(4p�Ŋ|}]���IQ?�Enc�܊,@�t�SnĵV$E�'��ɯ�8��|Z��?q��8+vq)��څ{�պ��m�d�(�i��!Z�X�����O�˓�?��5i��{@^�N�z��	_��m�'��1�']��'X��'��U�d0�+��� 'O���xp �\�J��O(˓�?�.O*���O(��׆_;�5` 0=XDڳ��),
��������	͟L����'��tYp�u>��#�D�S�-˥hD>M(��0�r��ʓ�?�*O����O��$ʙ]�S�W��[�m��2�>$[��	����?i���?�/OB��@fG���'V��"��[�5� ��-#qG��AMyӶ�$�<1���?���4�=Γ�?��'w2���_�TfѪ�8)��a��4�?A���$����O�2�'��c�!hW�l
AK�B����I5M�.��?Y���?Aʍ�<����?����$k��lԭ�0�X�A��0�!�;�M�+O8�Xt�Ϧ���ܟ��	�?��O�N�u l�R�i��u�l��^�k���'�.V��ya�~���O)V���cs�Z )�������zݴ6��hhW�i"�'�R�O���򄂅�)��AN�.����e�==�
�nڸuT��	����۟�����b�@!�6 �9d��։G�RlT)G�i���'�Ұ\,�pY�̕'l��O�$k��IJ0$GO��HTJ%�i�Y���~��'�?���?$���2�0e�#�W,[4�!�.)�F�'��E�>�*On��<���S��]�,0¤��揋V^*Dk"|}2y9�<���?I���R�"� 9����<���`���3кS`Ms}�_����^y��'���'��y���8��H�Ek��&� v$Ҕ\���Ol���O��$�O^˓J��5�J�D ��f�V�d�� ��񻀴i����H�'���'��É�yb��/?J¸Q3�D��(Dhۄr�B7m�O����OD���<9�I�����X��@�#IH�v��1��+=i�6��O��?A���?�V���<��?�t`T trb��&��[��ͣ��	>x���'�b[��D
 ��ħ�?��'|r�@�i[!�Z�А���.� Ԗx��''�����yB�|R؟܌[4m|-8��d�<�hQ*��i��I,�h�ݴxY�S��������WÆ\jc�Q$_4q�%ǯQ1���'l����O>�>��� �y,�p�J˨3، �&f�H �gaTŦ���ğ��	�?m��}� ��|��B	!ʐD�@M�Bl�6M�?�T��9��1�Sڟh�AϱD�&`B �%����H��M����?��ZKP�ǝx��'���O``�%j� g"�x�*Z2x��i��'�h0A���I�O����Ol�R%T���qB�N�.M��*�ڦ��I�@I�5��}B�'�ɧ5V/Ӟ^ ����'t�`"�7���*7#<��<����?����dW�rJ�1���K'~بӇO3Lb�{��S�Iޟ@�IH�	ޟD��H�H���6+W ]����)B�ر"i�A�I����ԟh�'gܠ��j>is�'|��ġߝK�]��H�>����?�J>���?�����?��&Fڪ�P	޶��P��d��
�	����ޟP�'*�i��l?񩑶Ll�9l�4M\̋�%ʊ2n�m���$������H� On�\�O|�C��θD��e���F�¿i���'5�	C����M|���¶�ɛ
9���!�h��<�D�^�ĉ'���'�DT�r���?�kË%r��}kEn֓$���vgd�b�A�� QҽikF�'�?��'Q����N�6ĺ`���R�@岗�7��듫���O����sՀ*}���'��J�މ�ųi�0pJ% vӆ���O|�d����&�擦�>My�b�<,�|X�G���:M9�O���-�)�֟,y�T
S��Q���'#�<D�A�Ɂ�M{���?���L��1���?�+������(�ըB�W\��;�!��#�&��R�G=�O'>��I����	�
��)���ݜY������E�DX���4�?Y�Ș��I���i�O4��3}��%l��f�F	Th����Ĕ=���䓦?����?����?a�͚=<���j�~�>�ذ��Qk@�A��?����?����?�'� �HR#ǣqc��)�
m��J�4h���'k��'���'�"�	���6� fFa��l���7���l�<�Q5�i���'���|��'��IVLr6O"��X���݉ ��y�n�e:���@�	ȟ(�'��2��#�	��nq{��B�l`�!�_
�hYmZ���Il��/�Ԩ�~��N�P�z9�@�݋�bS�n�禡��䟴�	�HZ��^��^�h����91�i�_i @�P�R�n�l��Ɵ��'�����X�b�$�5zv9��T���ժe�i��	�@�5"ܴBF��ßp�S���$G�ROzM8ꂰyF�,�ʹ$(�F�'��o��O��
M���ٖ}�y򀞹F�m�i�j�r�o�����O������%���	-�p�%L�dgZ�Z�*W:5�8��޴X�4Dx����O�p��gH<V�E�*P�(?��{�������	�� ��@b�4�}��'��D��,�� 
C��~Ԕ�
�ӂQ0�O��d��O��d�O�C@�PU�z�G��t�y3l�Ħ�I�m�*u��}��'�ɧ5fJ�",�>x�`�˯U\��Z��	���gF1O����O���<�qcС.�5Ps��y�x�Q'�H:Q]�*e�d�Ol�O��D�O��B6�Z������$-GX�#�A�s�1O���O���<��#�rZ�	�8'�L��"�=l�9���)kM�'��|��'�!W������
�l�g�5S�P!��H������	ƟD�'O2Բ�*�	�zl "b�{:�LS��,c��Lo�՟�%����՟L�%-��"p ��@�C'
U|=�T(��fz7�O����<�$��L�O�b�O` rV�I=5��v�X=/*0t�w�6���OV�D�����O�����ȳU|0x$!t��nZ~y�l��	R6l�T�'���!?�6H]!_�̽yp�?]�da93���������* 9�S�'x?n��7M]$�\��5�/&L��
�#i���'�r�'��d\��'6%��ѳ���]��8���� �p�i�ŰD�ޏ嘧�����F��`��C6���R��n�埌��ڟ���MJ��X��i���'��$�'�ҡ�LZ8kټȣB��5��MDxB) �	�O�$�O�H�0�$�X�%U#:2�Q���Ʀm�I( =�D�H<ͧ�?���I4q�Dт!�<t�PД�;2�,�;xe�<����?���?��>6HD��,�Dr ��nA={xe��BZ$����OD���O��OF������.\�s:�(� �5o���n�<x0��>�'�*ʱO�bbK�F�Fd�Y��2Z@���U�z!Ҁ��=<}���CW�F�\��=!�k��C+T��EKPc��i���i�t�F�U�,�r�*^�IN���BV��\�rA%=��5y�`>0;LՐ��>c��3P,S�}}�1bpEYC�B���G?	��Z��̆<��I0"_�J�@��L���< S��)���K���6,�[�π���p�I��|��|�ς�� �٨v� ˂>-�u8[��d�O�@�&�Ą!���ԪG(h�Z	�3�����Q>i�3)^;B��Ѐ��h(hA�R�H��0u�H+3���Y�^���Ӡ�M��N��J��ɑ�67�ܥۃ�+o�b�O�K��'�r��P��X'E��PTNw N�0�7D��(��V�Hm 7M��d��,5O`MEz�c6Zl5sA�/o&��E�`<f��?a��X>�+Q�-�?����?	�Ӽ������;��PJ}S2&�g)���̴>�pn����|&�h"�M -���G�&	�̙BS�X=	J�p�T�y&�ف-�q��'b�mP�E�j��$'Q�P�"Nԟ��'I�����|��$˼)yn0���&
�9�1��4@�!�ů,5�!�&�=A����V�h�����HO�SDyB�ڛi����▅j�^!�q�	Q�p����^t�����L���Ț^w "�'3�	� a� Ȃ��C�F'������_�<'`ё"Md؞�2ЀK[hHb��0���Y4�Τ3�j���g=6����ۓW��$#mf�`�/�5SB�������E�'�On1c��7P��t��ɏ�}�n��"O���f �k8��b� �\����n}�V�X�N@�����O��A�"�[N~,z�`'d�t���OB�䋞l��D�Oh�?l:lT����>t�n���G[���aF���m�
h�a*A���R� O�3��N����mэ4V7�܏i,��1�Þ�P��C�P��x2��?�����d	`yT���� �@�Bf_X�1O
��d�G/�4��!8�^��geN'_S!���Ѧ�BL�(ja�'
FZv�� h���'a�|y���>����L�x@r�$�:&�C3�<"�b|I�	Y�<^��$�OZ�Z�H�c������ |�T>%�Oq6��c더r�zh��c�B�]kO����ʌ�`�Ũ�m?��P)�	X-��R�fO;&m����I;}�.͞�?D�i�("}���mWt���B V����1���N�6���'
��Q����`�j�/�7LF�t�	�b���Z2�#'.�����m$p����Mk���?�؜�PՅ���?���?Q�YZ�Y�vFm�`��yV��F@�<Ęc���5�P��p<� �����Ň= B�8V$�oJd�*����Ր݇�I�xȬ`R���g�p,����:Ɋ��ş<�ɣj=P�)�<���!!vIC���4j�x�@ GP	'��\�
�'S��[�@��e�4}P���6-�OR�Ezʟ���*@��\H�H�����%(�N�@"O4��k�EȜ���Ɍ��9s"O>`0��Jq���b3f �I�"O�� ��"Q&���5��7Y���CD"OZ��EMb)r!����?  ��"O�m�QO�^J|�1�D�O�
�3�"O�܃�F&C�~t��J j��z"O�)��D��L̻�i��$IC"O -�P(V�47��uiQ
�|��*O�Xf�6{��1�B!����qb	�'΢�b�C�}��� �A\����	�'qH��"�!M����8FR�A	�'�������6����!���th��'#�PQ2Ɇh�����$.�ZQP
�' ��Y���F�(��i�?(t�A��'�Phs�욍#}2�΅�
{xl��'w�����;Wu�![V�e8���'��5�N"yT6��!U����'���0$���g�ĕa���M�M9�'�`�W�0۸Y���ۚO��d1�'�~=(ԬO�" �]@	;�'�<���Ws����%V�NRV��'�X�//�H��IC6>���
�' �U*wXN�:����46J]�
�'�Q���J�a�(F�4��A�'��۲d�j��������I�'Oӡ��r��Gg7)|��'V�	��S�(ܼ�!Rn����'Uf�OĲ$��E�~���`�X�<�T��/y�n�2wOKg��$B�	Y�<!��P�$T��!o�:@D(�dBS�<�dB�$�к�珳I���rT�j�<�s��#l�Ȭ3E�($��  �\f�<y�l�3(�Z�Q��	�erj�V��M�<�G��p�V����ם;h����M�<єMV��B���gȗAG�\��H�<	��?�X)�ul̹V!x�K��]�<��$>K%<pa`�58*�+p�9T���fǇ�E�B��a�TZf�i��1D�B7���vY�TD҉1�����g1D� r�IŅF���W��"lrd� �-D��	 �I�nch0�C�Z-&8�;@*D��[��9iЙ�0�'
�t١��:D���5�Ȩ;S��c&��:Rgha�5D�(Ѥ��S@�(eȳ(��<)�3D�(R�Oܬ!�.� �D�)C�N|��>D�T����R�Y�S�A��c�/D�ظUk�'q�pd��f��w(�32 D�t�g�I6q�A,�� �@��=D�Y҈�T
�10���D2q/<D�\��	��y����+�<�1#-D��'J@�N�N\�1Č�'�~�!�E?D�T��4&�9'*L�Jt$B9D�49'�̭!�m!�J� i6D��QR&@�ˤ�R'�ƖJ�`��f1D���s�Չ��LpcAO�Z��h)��.D��z�f�1o������<6����k+D�� "e�,����-Єv2NT�'<D���+��{�+Fk� t�%�;D���$B(a��E�tË�Wp=Z��%D�� �b�&v���(��G�}w~��"O�pZ×�5���.qlx�"O��y6��=�vD����Q<����"O*��"��/9�9c�B߳"Z�ئ"O���Q���v��5'`?����"OJ���&_Xz$#f�0fl���"O� �Aܺ~lx�����s�n)Sv"O��Z�#�~X�z��@�h!sw"O��y�$C.XA��0d�A~$��Ď�Sk|3s�HD�O|^�3�#�� 51sȐ41���'k�$��cʹV}0|x����0��9q7�O�o0��+U�xb����B$!��c�A�@�x�w�<D�8��G��p�@?QB�@	���O��0o�ԇ�	6�( �TC�4�<�Ї��E2����!u����$�����@]��B(i�E��ÀLZ%�2D�����O{�Z�Bǿ2R~��@6�
�Z���8��>R@a�=c�բ䡊��$	�� D���I�Y>4⯈�NTs�D,D����Ȱ��Y�H Ntsvc>D���`��aVpe����#9��}��b<D����R�q��X�!"�?��T� 0D�XQG$΢r��:��I�ܰ��,D�dZS�4?2�*	T_V��P�,D�T;�c��
V�%�R(9Y�X�2**��S*=Q�x��*K�G3VYE��iJo�|�B�(,K%��aS���y2�����2 ��0�Zyɗ���. � �Z,j��I�X���O��̐�8�"}je��h����O�Y����$�����S�x�)�af��-A�h8�b>e.��ۓGR,����#u	�=��ջ �ไ��!�5thN�R�����M� ÊH�)�������N�<YP/4�b�Ă��5E��WeH�1M��Q�e�����铁$>�q���S~�8 ���<�Q"O��`r�G3+`����e�5�"�n��x�I�GE����O��0��4^�pj���,�0my!�|B���p=y!G��,�)��>{T@�c�Y}~�bB7x
����	=B$��S^�R@D�X��F�m莴�q�"�ɡv��]��	.��r�;}��Y���I�J�?Q���?��'��	��W$s�FX+`m�$��g��!\�D1!�']|(�NH�	|
8I$J[4t\��*O6�i`$0�
AI��*�(��P�j��q�����Q��G]��p���r�L��'+��j{��5-�ɪ�'Uvuh�fC}�T:L~j�j[*���[��]j3#�TD����#(��_�@(	5�ِX8��X4�x����0c�'ڡ����Ϙ'��4��&ʝ�:UX�Ə��2�ȉ�Z�,jb��`�C�7�a!u�ϢEj��J��C�T�{�� &2z-Y
�}H�)3�,J�R�N,`2�ԧ���'�Z�{1��@�H��8��Ѡ2_���'��}#%#�5��ys��O� ��'�d�����'Ş�m�?s�XĞ�x�
�0F�v#���y0�L���O�HmPU�!5�����3j�6q
�,O�@��MI"VDѓ�JD�b\/�B�+C7Z��ѐ�R3$S��It�U�c %�3��>#����BA�U��x�#�=7*@"<��N�=�r��g��p̧��(�GӾpi
	�끾y7�%��P�������  z���ɽDc���>b���l��{q��I0)�f~ph�+(Nv����0�G�2{��Aq�G��X��3�,aƫ@���%9+!��	~���ڳo]�Iq��BaG1 ����#���V%��c�;0>t��9b��طgM�	�@eO@*�n�V69��C���$��,U=Va|�.')�@�RCA>��ݿRX
���f�69�J�Q�-pAX�*��ت��h�妍*1�>��͟�O�;������'Â+I<����;��=;rJW���{�G�%��y���ѣ��8σs��a×HI$�A���U�S1��2�gI���Ĉ.�D�8�'T�NPl��A�*��)�G��Bt� �F9_dy�v��"N:��;�+L�.���G�7J�[��f$��J2GD\�ٷK5o�!��)���Q��\�F�P�VrC�M�f$��>���iL0(u� 5 �4i���U��^F�T�F;2��n�%W�褨�sM����
R�a|R�W�Ր���ka�l+��%��m��#K�%[b����Q��!��:��L�U�m)���x��� �m�P��6�r���$��g� ����6$��8�B�Ӓ$jP�_>�R(�-	"Z
�,{�Q�F��~b�U�R@ĳ�N\�uC-;i&Yq�N����*����DѰ�n"�'"x����O\�Q�a�M��a`��}����"O`���U$~t8�)�Ln���F�'���RA�W�#�	�C� \@�O�ap��z��a��� Z�>��S<P�(1P�n��0=)�	;�y�Z=o��P�?tt�����:i��yI]�<�g�D����'j�(�r�z����b��E�'��H���nb��R)#�P(�y�B	cQ*'���_ �)���?��<y��;ֽ�#�2ۨ	��_����hךw��U �j!�P��s�'�	?u����Fa���=&2ar�W	���in]� ��g*W�"7�1On�С����I��*�6{��&�*)�兌6^ �H�?�FE�HO2q�r螸U��-�EF��+�@H��'�Y����t��Cire�b�@ n2�;tE  ��e�Qo�#ReJ�ɣ/
h EzBY8Y`�Y��D��Pʴ��$2j�pS�\�s; �"����]!3!��G�6ђ@nR��������[~Դz��F>w4V�SG̓I.\\�<QCœ7	�\]��O]��j�qCk�ܦy��<��#��qҭ�Ԥ�+�͠�D�j��3)͚
���{�j�,Z�d9�b�D�.cT���Cm�26�K  vL�[��IE�3���##� fτ��M���T?Ys��S�||��� �u������q(����"�����\�DEN�����8�=�%���hO��)�#A�38p�!��nH�>OLq�S�l��Ϗ�FjF��(�#7a��̄�hO���稁�Q=.���-��Y���>,y����"տ��؈��[�@���/��<�R��'��8e�X�h���s*$�J3�|���[X�� ��j��dax�8^����?d�"G���P��2�޹4A^��B�	=��!
-X�k���,<��3�=�)��H>z��+J<�@�4h(R�yȅ((PP�"�W�b#R����M�а����qҼY�o�Q�N ��{2n�*D/��m%���R�V�.�iS��!�J��R
șh�h��j�Vy�I�;܄�)�'A�a�G\�x1��3F��'�\�Z�D�u���D�D[p$	v�/[(�p��4Tz�9�� 𰁊�*G	�@A����A�p%G}rWN~��m�'E�
i��j��xr	G1Q5���E"��;вq�`�͹k�2PO�R؅��+C��$W�	�,,Qb@�_#(D��$��*ϸdd�c�?`�q�����*!C�0�n��W��L3���%J�#���*f�˗C���S�O�4�� J����1�RC�N��b�'CZ�j��w�P�%� �E���*J>�!��z��(Ó�<J��_-@`�H3öM&����Lk< �r�
*�Nyx�FܵDRX����#k��C�ɡ�f))�m\�YpN�1�CȂ�@��DY9-cB�$P�gH1\d�[�Ώ�p�(9+a#D�����,�DlSF�8t�`10pJ=D�l�P )'@1�T��%���Ճ;D��B� H3�F�E-4�xKC9D��:F���;��d��[ 32X̆ȓb�r�z3�\�2�t sBR?Xh4���t�B=x��}UTl��oT"�Bp������cA3'(<�'Ț�\J*���k69��#��=O�$�5a��)/؀��0�i�B?��=���@a���ȓO���()�&9�N0����2Vf����:̃s-J� Ni�5�Z����T��qa��^#aR��CS��~�H��A�JH�����	�q���g�����k�\�I�IQ�E: ��W�+S�^��#�j��s�T,n��C!+Z�=�ȓ#���ޏ �Vų-��J#�A�ȓ6���%���tg���m�ީ�ȓK��g�L殅"jX/e�i�ȓxc��5�% ,(`uX�rc$���H��t�M�*|s$��+`� ��(�Bh���S+p���ʈ�pb����Eaph�`;t"�xp�ˣ+�f,�ȓyT��U�ؠm8��Q�� :�BĆ�z�ZA�
�/:o2�A�M��L؄ȓb׌��F�ޔ�\|y�D�#HUJ`��S�? l���f?	c��#T��M^��HS"Ojc���3�L����7L�h��"O�	r$ьr����3:��qR"O�EPNI'(�z��X�r���AG"O�����D�]���A�,g���"O�ԩԄ�0�p�A�[d�J�"O�$w�V�2 �q Q�l¨A�"O��+r!R4>M��2���]���8D"O�D3)�&� ��A��%�9
�"O�t�Wj^WP�yY�)[� ��I��"O:Lpé�5Q<�P�Q �6���"O�ta�*��1��3���&���jG"O ��Ůs\h�g�ȉ~�R�ж"O�Ր�!2�P��g�,}P�AS"Ou�C�/ur;g�p� `�f"OB-�#�J�p�(�92e� m�V�`W"O�e)6k*'��Sn�  챴"O�X[�ɼ/�\��r3\���f"OF|k$�I������h0���"O���������C���5)�|Q"O����mǢ�SׅNԸ3�"O��1�y�����^$P椐��"O��0BFQ��z���7�(�"Ol��$��*�~��"̽A�b���"O��#��
mĎ�$�U�{D�P�2"Ol%p��U ,�Qr�O�;&� �C"O
��2J׾n �l*��&�1jt"O$� D5A�H!��C�8�2��%"O�������"㚥v���9�*O��2� z��+�*R�O�՘�'� J����L}:���l�p�vE��'�2��mf2�e���F�42 PH�'�h����U�w&P�r��nEI�A'1D���1�G���\Be`�]�:��fb$D�\��9'��QrGҟ.逅� D�Ԑv�U,h0,Zѣ|��T�"�!D�<�`��~�b�{'�������9D���d�6 |�� jԬ�0��2D���r#�E)���#?!-�m�aF3D��rUd�D�i�m��FŦe���<D�� �ĝ,���˙����(�B<D� ����y�Iׁ�
7�~)�Q�8D��j��1�lp�3�U�M�JՒt�6D�<��L�GF�,y���v���`%�4�hO��!yfiipHB4
�ma��ZbC�P�N��6�U[yh[�S4K-�C�	!t�v�����/%V�M��^�dC�$E��9[r�B��襏�=B2C�	&�(����3�|�H$	�1A�B䉪7�"R"T"�RM����T�C�45b��'�^u�A�H�t�fC�I��N�3�.�hذ��E'T]�C䉊��Ua�	y��¦��6��C�l�8�8�ܥԔ`A�_�,��C�I$>��{ħW�&>�$s�'��$�B�I�6�x����$	+�d��e
j]�B�I4!��q���hv������9H��B�	�8��i�G�)��ؓ3���Ha!��ʔDΖ`�$�5w�v�8�v�Q�ȓR�x�0e�w�8�X�bµ>U"��� j�I���zZL�u�D�l�&L��^tXp��] ))�d�D�ΉCru��BWN�z��_�}�����=l��5�����9B�:H����oE�Y����S�? $��	�z�	KG,
2:��`"O���#�B�	�@"�5wӆ �f"O�� �IH? �@`X��(A�,Q0"O0�s&���*� EH@�љu��|١"OV�+���?�l�Ä����qB"O�����B˪�Y�-�;@�
 +R"Oɳf�ظc�g�9�$"O��x�(G�rt���M�\����"O��7��b��yz���?0�ؑ"O�I�� b��9��,�<��"O�Mr�E��(3.Hk�ğ��b4�0"O�e�	�0.1 yB�؇8����"O�S���U�(rƖ��I��"O��rՅ	jYHX��2)�q�G"O��Q�׎u|.Z�$1%jj9�"O�LU�PJܹs��Ydl�2�"O`ɠ�Y0C��(���ʵz��cg"O�T f@�-F6��$���Z5"O~�j���bo6`��cݶu���ȕ"OJy	���x�d�x�� �V�� "O~YIǪ.3��Q��:d���#�"OH�zĬɣw�����7C�h�X�"OF���UA-�H� �ˬ\ªA�"O!�BEĜt�vp��
�d�J�@P"O�U5"�#G�.p��)�0xQ�"O�e �qz��Q#�"l����"Oērm1';�`�
-}�P�`Q"O�4	D�6E���f���D���"O�-�S�[�`)�v&����	�p"O�1P����p�M�E�$���QU"O��C�L��
.�6(�R"OpCL�n�-9�*�%�*�p"O�\"d�8`�����N��u��"O�Yq�j����L�+~ܸ��"O\�X���>A����M[5l�cq"O�p���ǏP�e�Ďrd@��"ON�p��P�!^��pg;X��Y`"O�$��R`��(�d�ȆGOhi�"OZq��("��f.�!@9:�A"O��	&�!8�1����{x�8�"O��q�ià�6�RՀ�]C"O�YS$�Ҟ�t��OԘIZ���"Od�ѤؤP�vd�􍘵k�$���"O5��ܰ�ޔ��&H����"OLa�Ά�w����Ȅp�,q�a"Oh����1д3�ȗm}=i�"O.y��@�7����`.L��{�"O�ei� A:;��8���O��8� �"O��z\�C~�(���=��"O�dzv`@2n�9cQ��/�l�p`"O� ���ys�[o�#L���s"O��`�);:�+!�W�[��e�v"O�4zDE��J��1 2��Y�vЫ�"O��{a�U�oEș�b�?Oڲ��F"OH��IT%g@�U��f�*'"O:UÕ]1y�
��Ơ����t:�"O(*��~��P
шB�*
�`���'��B4k	@�b1A��Z��=�w���b!�7�\]Y��]0/E�m��I��X!�D�0ɨ��G��t-�]C��L�!��ۀh���`�)�T��ˑn!�d�9Ol�Ҥ���Qp����aH�|V!��*N�<��(�kD�1H�g�5?F�>�O�� w�P.^}�f�1Eq�5{�"O� �YR�.��w�T��]���"Ol����b�0��G �8?��""O�D�T�����8V�p��V"OFXR��.m���I�rJ���"Ot�X��:I�����I:�h �"O�@p�g� )�*��c�_jNZa��"O(%��N�g���s�Om;T$�"Ov��e�9��c��Ϳv-PD��"O��ɵC¸��D9BI��C�<1�@�$NH��@C���1! a�B�<ɐ-f�����	�ߘI��gRA�<1K�x���C��gh��x�j
D�<�v�ۏqD����J�XJ�0�d#�U�<y֬ǫ�.Y�g�.��-"s�R����<Y�L�.��rƋ�V���AJ�L�<Q��1�̭��#$*��e�G�<�5�[��1ɠ����aJ$�[F�<�6	ٌmL� J3�7}�8�a͘A�<�!����A��ʰ�v=����y�<a�M(z�A�gL�*u��Ho]`�<��� Wj��yf٣Y�`xaˉD�<q��S���8x�Qi�C�]��\���d	{lA���-�,2M��_B�b@юY��[��K�r�3�'pra7C�b7���爛�<J�N<��:���w���R�~���o�s�d��C-n-z"���O�F)�J�i��> �����(�, �t��5h�ՄȓK��@q��:W�*���Q��=�ȓ ��@��BD+W�^n�p�x��'qd�xQ�]�4��cC�x@� y�'=�8��@"�&��ذ=Z� ��'�Z8����n�@�lU�d�ⰺ	�'\�.�u&��R5�
'Fr9��'
�Mt�&\��Ԭŧ9��H�
�'���CŦl�<���11�T��
�'T�m�d�M"+�~�d�4s�^d�	�'j'��rP��4`�6�b\b	�'����b�ln��C�Y�/�'Ŧ`P�F'X�K�DO<0��1[�'���`�Q&�4��Qjȓ.[dqR�'>�ICe$*k��1Qk4�VH��'b���'�9x��:AĲ,t��'�d��	+�^�З��.Y;fL��'���SD��"d���C�zє ��'r�d�����|KR�dGѩ[<t���'7�Lsn(	Cdu*�DE�!>"���'��x��2�8�A���+��<�'V�
G�, Ҩ�(���*�h�'lB�"���3[\��L�L@��S�'"�9� өt|M�a�E?ґQ	�'�ڙ�bM	0z0�� c>>����'.�E��
_6D4ڕ*]5	N�S�'{��,��
����恔52b�B�'��c���0�����J	[b|l�	�'ڤ�"6�1^��|av�ψ&�,)�'�BH ��>E�
�ե�V��'b*kM�� ]X�2��&Zd��h�'68�s��!j�ބ`�)B|���'J�pB3�(��GoK74GF-
	�'�zͫv晰�x  E�2W����'TF���.C!z8��G�Ȏ� 	��'k�ASD.}�8i��F�@���'ˎ�	��̥o[\��`K3@}�L���� N����#42�D�6��:I�X��"OHDY�/.Q2$19'`ЧJ�DХ"O���gG�����C�(3S"O�lx��
�=��H�RLT�����6�y�sL�:T�O(b��P'��y���*7�՚6�\�%��j9�yB�
�q�
(�I5 =� ���P$�y2��)�"(�3*�q��=˶`N��y�7(4.p�E(ؤ{���S�Gޗ�y�.�4q��И�@�?��kM�	�yR�;�8��ڭLNL� t� �y��ϖS4Y��fV�X^��k���y"��:0|!�R ��}��R�D��y�e�?-���:���e��@�w�U��yj��^-����e��+a92f͆/�yG<j�� 6�
+#G��QE�P��y��Ht��kbnд> �B��yB+��J��i� �Ǜ2{�V^��B�I_!ht	�FԷsG�H��FM�d�B�	�x��)��0!�F�B�F�V
C��
7��=�w��?6Q)�Qn�)f
"C�	�P=R5:�M�7,�>�����M��B�	�p�݂��?&3<X��I��ɠC�Ia��R`L5p0,j!���o�C�;�^�s�m�;3xr4��6~@jC䉻 �T)���MS�-S�9yz|���&ԙ�	�
� ��`ȅ�{�J����Мyb�ȭZ���j�hL�j�N����$��A@Z h�`P�� m����\!	��M�v&��r
أ5�H�ȓ7�nɳ��Ab��$��Ԅ�A��dI5*�p�l��	v8 ��G�ޤ�T�R2��℅�8[jІ�S�Lu�!K�VD���%�.�\<�ȓ}D�*�jָg�xщ5��q�Z�ȓ/�Lui�] ~��!ITŽO����E�L�h���OIzH����∇ȓX������	�1�B��4: �ȓ/��jG���?Ԅ�b�0j����ȓ3�N���9Mj��	�z�Շ�5������Z�a֞9В�����a�H��xQԧ��`l�����y�Be59��ʒ�I I�ʥ��VM�ܣAĕ�LYZ�	�Z7J���ȓ;���15.=J��U���8X�ȓn��9H@µd$	��ߙ<ވ|�ȓYqf�걏Z5~�@�pv��g�z�ȓ�$��M�j#zL���*vp<��P�8�0׎W2l]��ʦK�h�ȓN�V�Km�x�����N(蘆��Ѐ��~V��y5�I1�L�ȓG�.9�#O�T�ș�iĨ
;��ȓ++��)�
6+��P9DL�	SKh��e���Z���r{����d��L�ȓ���K LU/��l�@O^�[�z�ȓeJV�نO��
D���uh�3I���ȓ���G?<�V�p��ŬJj,݄�m-��6��5;��b��v��фȓV�̈�-УX�
`��B^(U&x���_������^��z}�����\��]�ȓ_���+�*'τ h���e��A�ȓ"���K��O
f!k�O�@s�@�ȓ7z�4`�CS�]����'h_ {� �ȓI�&��B�?v��4邓V̄��S�? ԱBa�I�p-��道@F��"O(��tO΂h��(����>pD<�!"O`�S�)_:M<�d��+P
6=PU
5"O����NE��i�!	��8�c"O�I`�ϙ�H�,���G�/R�԰�"O�8랔v�\�¥��}��}�R"Oz	�q��>.����X[�`S"OJu��ɸ>���SCP)yh5;�"OV���$��H\��q�"Oق�&� ���шO;({�͹V"O�4XQ�˩AW�ZB�4om ���"O��Yf�ɘ/7�u"�g	�;�hl��"O`�iA�1E���I'�U�l�C�"O�њ�*¼X�w��;n��h�"O2RT�8$�Yk�Oް	�>� u"O��J���7U� �D�^�x���"OT�����
 )�VNP�J�nQZ�"O��UO_Az�QC�m���!"O�%���E!�Bmx G�-�rݳ"OZICR�N,.�
 �<|�$ HE"Or���¨a�h` �)�Q�z��W"O�@8jՒ4t,��i��AH����"O8k�hϒ"�ri#�ț)c�tyf"O~X:���> �i@��a�ּ�"OJ�C� �ftY0-�/c�,�w"O�1��b�����>y�J��"O���	�;F\�r�)g����"O��+�;9{��"dO�?e!�PJQ"O�
�]�(���F�Te\ͨv"O�1 S@��^18@�C��&/\2Q�"Of�{7���b�X`&׆vI�l��"O�yCa	��bx�D+F ���"OX�K��@I�ѱ7��?)&]B"O`5ڵ�8ws�+"�U���0�"O���&!)�u�q靋hx��+b"Op��m�3V8!���\�p��"O���P ����Z��ͫXN�-�&"OٱP�]��L �@W2C=�q�F"O��J����n�P5��/L�%�g"O��)�@͸�0|a�I~@�@"O:��!�V�$�րB�= ҥ�a"O�h*UM/��M* ���)�6��V"O&8Ң#̕xl�[ GE�2��A�u"O�,)BϮwiԑ�e�@߰�!"O�4a��+��  "#Kf�8k�"O��Kr��?����ၱV�☻w"O�E����Ac�(�U��'�:�3"O� ��	ؼ`6^9�L0qP��u"O,I���U�������CO��7"Odt!d�^ Tޠ�P�$g����"OB��dGQ��-rtaQ�CJbTr�"O$!/�^�1�.*��#"OD�c��7)��� BV�L�P�Pw"O�T����S�ڠ��"9@d�ZF"O��RD�@�Pg�h�@&]�W
�)�"O�[���:hZ(bt���y�5"O>��‗ kvd��ĕH��9�"O�IB�S��LM�3�<pG�ɳ�"O�08Ń�$��#���`�)��"O�A���.}��kb��pP���"O*/����qR1�M�2�sq"O�@ �+�>T�����r���C"OT�p��G*G(���U� ��"O���(��5�<�˲b�"Zv
	��"O� ΥH�������kU�$XmB8�"O�w��[��͐C��1[D���"O��Ipo���6U�E��0H���"OBx㵊��o\����>���!"O\�hƈ֌o,�! N	�p��,#�"OR��%j��oԀ+��
 4�Ƙ[��'�ў"~� 	Gu�A�e�	"n�@,I.�y��F��!����"-Jvy���-�y�M� N��D�PFǜV/NT���ߏ�y�c۝[F�\����n����^%�y2����5�n�~�C�!�yRnγF�X��uG�*w����g�C-�y�]�s�T� pj�89��	�ч���y�(ø5��u���L�6�T��	֘�yb��c����J=6�����U��y��rv��1#�Ċ0��� �a��y�⒕Dq�S��ǋ'�B��f���yr�S�/���' 
�"Tr������y�LR)A�R= ��ʂ������yb�ר0$"@2�Hі`�|���3�y��S�4���\6r���	��y�O�>�|�`�j���1�D�^�y�%g�� L��T�*)�A�;�y!S�(r!�� 9�
���y�oY�KN��QLE)~��cRBŞ�y�hS�X�P,�f&P�!��Y:&!��<���Tk�	U�=�`�i��	#c�O0����2\
}x�AL&hUh�ǜ B�!�d�6w�xl9��ȆR �Sv����!�$��C����M5?#��B��#{5!�T�+�Rj��Y)7�D�@��!��G��٪�C�/&�bj�5!��:de��`�\=Kf��0!�$
8�D���T8<�s�_	{�!�dг�"�L�,7T	C��J�!�d�BB1uC^�vF��cgρ {!��C�>��4�##4��Vg�7[!� C{�  v'օG�>%���Q�pV!�=|���ꍶ}�4�y�G���!�W>}U>LJ7�S�N���z�]�\�!��2��ܨ�"H,*��}[�+Z�!�ą3f|B�B%̙�#�
��&�c�!�d� )!��A+_8N��'h�'#�!��3C�1$�>`���f�!�d��{V��  )�^R�� E��!�dX���X�t�T�N81��a]�<[!���(H��!A�Ȏ#6�`*B���5Z�',ў�C~2���)�<��6(�9��G�M�yRM��]+΀���6h)�7'L��yr�˸���ˡC�\<d�HW�_��y�e�[�*�̂/����VEX��y�- >l�<��E24R��5l���y�E�'�h(�ĩ	��a;r
�%�y��8g�P{v��*5�X��nR��y�	��r�x(7L��ykA��8�y§VMvh�P䛉	���pF޴�y�!*]��������J0���y�. .D���-t���q���yrN��?K�rg�Χfи� ���y�L�S-ލ*6�.X����O��yr�Jnha w�W�JC�!��MF=�y�KK�I ���@���̎�y�)T�0#f�y���LN�){1��9�y�(Y�T��]���-�:�[�jE��y
� \I@F�Ð��3�K�Y<~�2$"O�Q�*�	-͜�z2�]�)P�b"OhM0�ER��v<1tn35�d�"O@�x���wC�!9֍&>�x��"O�A�dC�<JV8X�o�EG�""O(���!!��0X��N@�4�R"O���qd�&5�2Ē���.:*�ث�"O^U�t�P<6�i8%iΕu�jպW"O�A�%J-̅��'�%�lt�R"O� K�fزe������bI�ٵ"OδT��x��ɰ�A���@ٶ�'�ў"~�������iuj���a"'��y�!uB`�X��δy�����y�FK�LYpG� |'f�D�yr�O�#"����P?G��C���y��O-�h�L�*=�F�01NA1�y��V�𩙕�9ٺձ���ybL�,%��˅A-@*������y�L6Y���k1I��t�K�y2,\l���#�X4]<�T#�y�i�eR)3�!�,<j�pb��8�y""��/�zl�)�
8D�%�v��䓝0>ѕ&O!Oz �ԏ+!(%c�Â]�<�QT@,dk�m��<�JC�L\�<q�^
LD1�5ǖ<�V|*�$[�<9��L���)'h�>}Q�	��K�S�<Yu��KĸT@�;)�I@�UU�<�"N�Ȩi���D��R �&KBP�<�@���WMnl�-T�]Lj�[���M�<Q��ML�)�Iͨ��a#p�YM�<)P*G���	Џ� "V���hYc�<15"�#!먬X�
�<}"��� LD�<�姁ܴ!�'��f�=j�B�<)����Z��ճ�l*h����G�f�<Y%A1v�*� ]"���2��^�<�nYS��)M^b�,�Z�\��Fy��Od����K�9��K!d?K����'?��� ����B�gϓ?5�I1�'�15BA(d�~Y�֋O?�@�ϓ�O�\�GbќD|�d�R'N'Wyj@�"O�z"Ɯ;`u��tE�pb0��"ObUb2ջk�zL���`e���J�f�<��\.L�x�"ō׳�°��X`��w�(i0��9B�4���U/>��m3��.D�<�&��P<�!!0@X ��Ex�-D�lړ��*+�5��'��ȴ� �	s���S�bXX(�J���n����Y�	��=�ç"�^88V,Y� <��dg�2

�ȇȓ[����	�t����60ݢ܆�^E��� �90~�At�I�C��<��gk�,!��ܗd1�q�qʂ�f1֌�ȓ2��ѫ�O
0|�t2�Ǒ�*� ��\���1���v{4���dǊG�l�?�	�B��R��U��P�%.�8u�u�ȓI� ٕc�5��� �A�N#���s�}J�FQ�m��2W��?M��Ć� ٴ�{p�� � ��_�hP]��yXF��գ�Hj�=�����05��o?
�3n� z% Qm�.|�\�ȓv����Ã�P[ލ�	�����ȓЄ���Ab�Eђi��f�!I�U��D{���;H �$���(qV��E��35�!��en~�(���a]�	/�t!��3]������, � �()o!�� 4��n�"�HE+s�HZn�Q�"O^�X���	��M®�*��9��"O��iR�s�yғ-�]��Q�"O���>�Ĉ�!�e;��_��'��>�7#�,H�*�6ؑr4	FV�<q!͍kՌ,���D�^�Sg[V�<�C�GM5*�I]�
a���m�<��B+M�z�T�D�F�𔛱�S�<f�@��yh��E�0��E�K�<!ǡ�k�K-f�}k&+�h6B�I�r��	!Qeӎ
b�3G�����$3�h�q���]&��G�N����=D�HȤ����#'� V�N���&9��8�S�'3{D�R$c�-��8R�G��ȓ9�8\	g�N�f#�q�N�=!����t_,�#v*�#|y�ф��͘���\0-#�l3I�V��N�^f�!�'�ў�|2G!"e^Ĉa���-3LGe|����Ia~"������	�^�Ρ�t��y�D�$"+Rp�Q"JX����D����<����mm���C
�.�h���~�!�D�%��\�W��p���*��9&'!�$�����p���&=fUrWo_�.w!��R  \.�W�ֽ@ڴ�� �~D!�D�=K��ɂQ��r�x�2�.P��!��R.iC��!����5˘����P�j�!�dE$%� �5�Q�9�,�2��s�!򤂋2� ��,��<��d04�ӀR�!��l�6��5��܈��T�8�!�H��bVk�.T�:��U�R?b�!��1+�9�NO 6'�պ�F_3k~�}╟H�"�ԍO�Ir��p"��*��'�S�'H��Sa�ݱB�����
:ф�`�d�7�B�zhI7��L��ȓ�$Y�Q���	&���띖/m����R<��*�8@@t�K�iǊ;��X���c�<��Xu
��-Kb�t�P�G�\�<!c̏-� ��A鈽z�(t0!D�Z��hO�\����r��L�8`Cƅ(|��)o����ǘ^���� ǈ,,���]ΔpIv͜7O��ᘒ�H���D{b�'5:��]�p�HP
L�s�2�'�
�!KT�E��d����^��'�"BC� <Z��CI�J�H�P�'�h,���߇h�$�
��5�v0�ϓ��'C��`���༨c�O[��M�2�d8��s�r�Xp�G�Y]!{�
[*�2Q�ȓm�
�*����N!�����0fep��ȓ^��1�r%S�l�5�֭��J����B�t �d���|�ص�ҁ�)s@�ȓj�����
U3<�^$����T��ȓ����Y@\�pAe��2BZY��8�0� �H� E0u�6JL���Ԇ�Ip~2&l���ˁ�thx�&����'�ў�O�>�y���ep��in�-x�pA�'Ƣ!se��#��i�������''5��Gؼ/�l�#t�ړu$X��'ǆĩwӿMd�!T�NY&���'S�q�%�ΌC^���G�c�1		�'U
E˄��*E�,�[dl 'V����'G������<�jʘL��d�ߓ��'�0��b�L?��b�Ow�Y�' �Y���<v$��tJq} T��'�HA�ŮH�c��)�4�Ԍi,��J��� (
���&J��A�/T`R"O2�h�:3Y�!,Z$P�B"O\�� �2��T��iܠX"��IB"O�tE�`i���e�ֲ@{"O�I�&�|�U��A�0�"Ol������D#��;� K��b�"O}9!AW?7���Â��`X�U"O	�gB*�����+G����"O2�J
��Ctp`�Ӆ6Ј�"O�a�1��?�|!��=S'"ቷ"O� r�����$�0)��x���"O���u��o%��:p�^�1	�"Oֽ1�K�+&%KT�6�)����#�y�aDhh��B�V�)�\�e��&�y��c�@�Q�_P�(�$���y�����h��
>F�`Ă��y���3��jr)����y��t�f]cT��
-���fb��y���3vɪ�'�&���/B��y2-��bAHXRF$�!uҭh�"6�y""4A�@�,] x��F����yr�"0>4y�`�;���A�yA�v�J�ѕL�8p�����?)���S�&gz�2�=J��t�����ȓS����b��Nju	�N���L�ȓc�
t����TFhY�7Z�J��W���
EgP�s�ڈ{��(mh�'��It�)�O�ra�Q8K�������� �"OZ�A ��1��i���[�`pB"O�5h�F<8����Q�E�0b��6"O4���F5�ZQB`ݎG��cR"O�$Ȓ�	�~T�
��"O��sŠ�|\� `���9���J��'S�)�'	��͡�V;]Mr H�bF�Vv��	@�����8z��Y��]���	U�.�I�D&D����DJ?��Z�A��zu�h	7B&D��q"̒�/�m�.��A�\m��$D�l�D��*F�����C��r����'D�8���6���� ��� D�0d�3Έ�K5�ԺP����8�ybH�+l��3�f�R�z= �S!�yb��#E����kM�r-�� ��y�+^�k��]���]�J6�M(�E��y�\��X�:�@8�2��&�3�yR(@�#gV�A��t�Yƌ�?�y�aW�D4����^65%�L�b�A4�y򆏉8��� Ã*�V!����y�Վch��Y�r���Ѧ��y�C�$��͠���b����nV��y҆��y��d��T#��1�0��y򥊡R�d�:0i	.=i dY��y��H�� ��]�d^�EI1��3�y���32�3�S�lu��E���xB%��]���x�I [� YJ�E5��O�4�s�[�]׸m��$�>6�,�Z��F{���
?^��h�1.�4G���i�,+/!�d�p�i2�$� z�(�X�f�<U:!�d�7Q� 11v!I�p��A��B�!l%�'�a|�X�q��i�����0��/Ã�y�%܏	�B=�OJ}H���$�yb烶@oZ�I/ѐ��P�$$��y� �n��A�nZZ뜜Q�
��y�ʸp0j1r�KÅM��1:��G<�y"̚	0�`u�D<��3����y
�  ��f�6t4�(餦44�*��p�|��'����0?�PϙL,��>*�.�$dg�<����b���mS�E
�P���b�<� ,59��$���3{F��*УZ]��}���O�$�KՌ،}hJ��R�Y�xa��'���X׌�5}70�k5D�:@qx��'���Fj��	��d/��D�3j��y�aR�J7L5�⌎C{�}x ��y�H��-�1l��;R6<r�gZ$�y��Ft��AQ��׾CL
�j���)�y�U%�̩Aa̔Ll���Cץ�y2eR�.���y���5�&xA�h��y��L$n�:��kH>��!�����yB��T�:��q�1H�B��yB��}��ɳ���yz`�	3H�)�yB�P�oX�8�c��w�By�g���y҆h�J�-J�%����CP$�y2���6A1��]> ɶ���#J��y���tRċ�LA���`qě��d/�O@y*�ިA1x��@�D���"O� Rg��a|��s.D����*s"O����Ij
Yz4�C<i�uP���<�Iџ��'24�x�(�Q2�Rqn˲^�a"�'��I�#��!=!B��!�O����'i�)�f���~pm�Q�G�j��[�'k�`�W�+=aTL���A.~���xBה�<��k��b
<a2�D�yO��82�-[�nl)"g���yBF��%�4��/+9�0p��9��>��O������{��	uC��|AX�z"O��r���t�t��a��/QN��"Oj8
�_4l���M<�!Y7"O��K�+t4�@!qA�Z���W����I�7���)%^eU$�#�R#S��B䉜(&�J�/21Lp�R3 ��C��.l���ѡ�96�	DF��=�$���O�c�,!��V�~�d��n�eT�5�0D�ܙWG[	9`,�t"U[�����-D��`�P����'.!d1���+ړ�0|R��U�uZ4���&^�c{^EQ���T�<yW="�D؊����rِ)���Q�<)�g�"22<�'���2���`d�<�w��(i�P	@Aܰ P��'&�h�<ah��%|��V/�|-�"O�<i��يS�2t9Ū�'�v�1	B�<!��O�\����N(9�����y�'�'r�S �hـ��F�:���&	(ƴC�I�P�}I��Wi���%dN�`��C�||�
d��5LKȔ(2rcPB�	�2 ��Ğ�%��LZ� V #(��O$��h���^$P�|�b�:��ꇈR�`&!�E$U�r0p���tҴ�����V!�y� 4
0���el�t��#q��P���:K�|=�G���C^8�Q�Ϟ)��B�Ɍ.|����m��ʖW�FC��m#ڥ����&9`!��.CXC�ɡ=|�v,���pgJ��ʓ�0?ID���t��egM4g���@�z�<AF��,��!U�ȴ&$0l ��Ts�<y�n^!:�7��+��	p�f�<�tF�s=F�S�
D|{� �v��j�<�x��ϖ;�h%�e�Dp�<Q�L'kV�s�P�V��l�U�<�'�ʵ;������@O֡haL�T�<� �A�ւ ?���pP)#�X��"O,=yB�� �si߹~�.D�"O��h6�ҋ ����^ ��}X�"Of��r�E=.�Dp���
�y�ЁC�"O�X��R>� #�G�&Z}�I�"O~��R�S1��'@N<fj<ٶ"O��Uር?���UM"d�����"O��!�Γ�k�X�ST̖|��i0�"O*	Ӥ���CK�<۔��"O��  ��/q&Jƛf�f��S"O�����,����'Ъ^��%�e"O�a�_������z�B c�"O�ؙv�_U_RI��%B�0d,��"O����J:@��@RׄN36
��"Od�p.��D����t�M�s,($X�"O�]	�%G��hsf.2"�t"ON�+��C�xp�Jl�$3��� "O(�L+\����d��bt"O4�D�B%@�TspLS�"Ƅ��"O��k�(]y��F���А�"O>��f"��n�RM"7��4�2�0�"OZ�I`e�
�$�0M��X"O�TPC��(�N�s#@S�?W"Rc"O`TZ����+���R6�I)T�Xw"Ort3��U11���fMOm*1��"O���g--�.��#m7k�Q�%"On1�%,�� 0�aC둙*{b �"O�z���=pY��I$z��ܨ�"OȐs����u%4�@U��S����g"O�m�@�ã9&P��'I��M��"O0E��'�M���G�QҶyp"O�)�3�MA���u%��_�v9�"Of�#�aB(3�A8����}�c"O�X��@�J$��a�X�b J�"O��1rKH� Ax����=/�h�92"O�hк}7ti(쏰{���	�"O���V�[/u�@2u�%K��h8�"OH0�7"^� �\��j�*��(��"O�Pa��]CԿ\j��Sw"OHq�ƫǇl���1aB�ng�aJ�"O�@��$HB�BYAUs�*]�q"O��ZT  �[+d��S��{v~��F"Or���PC"��Paːn^�r�"O�P���1Dڦ�Q�eM7G���"O.Iz���z����&��2���4"O��z5k�:G�Vy���ތ�)!�O�V�pDYQ◴&,&���l!�U�3��u@�c�3;}]J� �!�D;*���e�N�fc�ab#ꛡ=���DZ�:�d�/�*�D�_�yr�шQ{�L:���9-�%����y���(��Q!���  	ᘷ�*�?����'P�lrů��p��S��[$O]���!�;D�������[���c,�L��'�9D�X(�a yd��	��X������2D�<J�#\�r�TՂ��W;�=�ï/D��f հn��l��ն}Z����-D��pA�8ʰ��!��l���6D�X 2��(d�lh`�L�:x�L1�d3�OdhA䉏8	:A�'���g��̒ "O����hE�J<x���?���"O�I��Þ�U����}�T�&"O�0���f��(�J�y$2|�"Odt��0�YA�c�7\��TS"O� �H��C�)��Q��"S�P:��"O������!t2�P�@�l��(""O�(����xZ$D����lQJ"Oj�R��R �;$l�!���C$"O�����+7D,��7��I�V�X�"O��D�G OԈò@"s���4"O4q�(\�l>Ma`�>c��Y��"O0��eH9�Y𒏔�>�܄�"OX4�i��2���re��>� ���5LO����/熸�c�>>�D���'{!�$O�#��g+�'o������"5�!���&� ����7)}舑P�IZ9!�DTVVA#ad�;<������S�yB��&.6�p�h�^Q��ڷF�k �C�� x�'��ZL� XpѵQҦC�	�F4��͈���rE��.&�ʓ�0?yeJ,>qi��5tAFXGǙS�<�b�Ԃ<�0)eh�2%G�ăE�y�<q'ƕE�2D���Δgf�԰B�Xy�<9@��:B��l�3�P�kP���V��j�<�ANεcm�����W�`4PX*h�<���U�5b�X�V�0� dA��V}�<YP�F�F��D�*T �u+��@O�<���5<�� �/X(lI�A�s��V�<Ak��-֔qa�I�	V����r�}�<�K��[��4��
Z'��WHE}�<��!R)k2�m�m�&&�he+Ё�S�<����F��h:p ��F�j�<Q��X�Iqg�A2C:d��� �~�<I��I5A�d�sb�7
����l y�<�r,ƪSh����'Q2h��y
E�t�<�C�!=�>U�Be��ofF�Q��e�<�1P
,x#��,hF���mId�<q�e֩iXh1Q��]S���p�N^�<qӽ�����^`�!*׿.�tl��Y0�z�MH%��U��U<��/�p��@�Wo��qs�<�5�� p���.\�f-�!�n�p��?�ӓm↹�R!�<b� ��e�h��}��覄�F9[$F�,��%��XR̡���Μ �st��j�܆�\�pdIC�� ��jqNV&װ܆�H70�ڑ�E��s@��pU�d����!��!��}��$�c��>G�d��?���~J�G�Jj�����́gP�k��s�	F�'b1OL�� ��F�̊��S���"O��'J	�XT��iH��c�"O2�*D���(ҥ(ۙ{r�T��"OP�g-* �\\!4M��m��Q�"OrhiΕ�)��@�a+$*n�xs�"O���Q.X.%�6�3��ͥ\TryK�"OT4�p>rTt�F��G��!gU��D{��)ĹK6QB��?gi����f!��Ɗ+u�qR��[�m����Y�!�]d�qj���;��e�S�G^��O��=���9�w&�	GC܈�Lتc�,��"OLP�h">��h�3����a�"O�K3�T<z*��Q+���G��Yy�W�4u8�v)]�>�N�3�ĸ|@!�N$4]t��UN��u�TM�<qW!
�CB�m���v��2@�PH�<��lh���2G�=I�"a�Bn�<�� U�$]HP�J��'Mz�y�Õk�<�t��<6P	$�9I��	�@�i�<� ��+Ǔ(!QT	1��a�9 �"O2��e虥dVFt�S
�ht��"O�j79)�q ��-+�\��Tg�V�<��.�1����G@!Ŭ�zT�MT�<A�l�Ҫ�a��!�@-��(R�<q7FT�t)��LH(�cC�<qe��(On���e�
,b��C"~�<	)�&g��]&k��9 �|A�|y��'O�h!��.s�zP�+m���c,O4���5�b�(g����@?^����'�qR�LB�A�Y�f&�*R2`�Y
�'4�\�g�O�S�N�X�J�4����'3�!�� �,����R(he��'����`ÙRȠ[Qo�)&a�p��'��U��O��
qF�Ya螄">Q��'"<��Ϗ����K�\�P�'�����썇A%VtB�B�3���{
�'�����B�D8�d���W���'X���O@%:�4}r��6d����'~��Sag�>Q�A!���N>�A�'��Ue�V:�أ�99h6��ȓ+������>�P��a%C�� ��ȓz\~$�$,�m��d�ݭ�ڬ���v�2_�je���4�Q�{�~��:���r �t��c@@A�m^�'��`r����oµH�i��@q��' $�gC^j��q��5�Ju�	�'P��@PE�lnt��̑���@A���%�@��2�G�V��t��!BP~��@�'�!�d_�]���SdDS�u���2@��M�!��ڐ���R"�;C���!��h�9[S�*
��[�D�!���4N�FP�D	$��_�!�$n�����&�"\�t�s�(��!�Y'Q ̩id���$!rt��!��-�䁨��Ҫ\2l�@�ڭ#�!�D��U6���#Vtܸ�Ư
�Py�F�&��$�AH2+�vi��Mݫ�y"NI�(��F�4^��@��yb�j��y���3tґ�����y���v|^;W�Ȕ$�&�K��!�y�N2걒&��n�� "��yb�U.RRL)�!�%~(�a�BS'��'�ў�O����fk �6��E8�g�7_���'��`�u�2�
�7��b V��'��]X�,΂�*eśT<~|C
�'i�'+֮P+`�����N�4�:�'��dq�j��Y5T=�EKS�L���(��)��`�i��1P�B<	���ȓ&���y��\2>��ȳ�c��B�bnE��y ��b�,�c��R5�q���y�G��N��	x�F8S���)��y�*D�qw����N<�Y������y��W"IR\��n��JC�8U��y�OB(A��<����*B��X�/�&�hON��	,�
�	�}|������%�!�<HJ,��TH��tn����=!�$�>`���v┎_Y��h&�\�~�!򤓰?�"�R �H* ��T�CF��%!���n��c��B��hYsD�> !�D�#��h�F�F���J�R	!�D��'�P�qD�]$.`��P��e!�$7=^��ђ 7h���F�\Hў<��.	X�LB�cJ��!6*!�"B�)� jL�6JE�% yҒ$�eM���"O����B�65n�x�C�-x�M[�"O�h8V���u�� �m�<Ͷ�ړ"O\C+�k_��3ċP�uɠ��"O����M_�+���a���6PȔ�q"O�����+m)<��gJޫ)L�؉�|��'��*����-��P����AJt!F"O�qA��5�Ph����WD�h8�"O�a*�lT� �m�Ċ�#h�h ��"OP�z�ǈ�2i�|)��
5 �[V"Op���L��l�U,�#{غ�"OvT����4Y���	ǬV�P�|b�)�=XBNX��MF8A�%�Fo��P�O��=�}��h�����jsBΩ< �1ip�<�Sk��$� *V
��3�@�戒o�<FC��x�h�d��sƄ���l�<)�AT�L|.��2l��N��5:�-Rf�<q'��0i"иqɉ0��Is�'�L�<�w�ɝw��	�gj�fSTS��E�<YF�."��Y�BO��N���Z�m�f�<�vΏA��pkņ%e�1��Y�<�T)R���(&���Z�B'l�Q�<iA��Yg0	�5;�X4��Öt�<i����p��pnN�R��@IOt�<ɲ�g�0�)�iF:B(@�8�X�<��JY�bʽ�l�5%~�x��V�<�1`��d�	�G��I�� Ug�Q�<@C	�$@"fç����6OK�<a��;[G��CQ�֡F��h�w"Q�<��Гx�e�aő�X�eX�(�g�<���ҏOP���"2F�)`��e�<���'*�"D�E�4ɮ��`�JZ�<ɡL
&LE� ��b�J���LU�<�BL]k�j�#�^�R��P��y�<���SG�DE���R�� ��!v�<1��(c:ɛ4i����2&Er�<Ƀ쓅��p���c|b�6�d�<)p-C�[��c�(�2M;083u�CH�<�(���L��2AʵH��%���Bm�<�VBX�X
dS �+���
�f�P�<	��	8W��ޥ&��A�%gK�<	6���R�fղWL"�h�ꀀ�E�<i֌^:�`&c��	��I����E�<�7�5F�Ӡ��?9F�r���B�<1�.ԗ(���ɥ /t�0��I�H�<Y�NM����x��J����U`�B�<�D��%t����%G��1SJ�<��M�=�:��3/�09;��%��C�<13+�*S�52G�C5�I)��<��J6e;"�h&�Ѿ�qI���z�<�` E_O*�s$Y�2�I��hx�<I�H��$��XBMS�1�]�BKr�<W���j���lM4<�8�B'��V�<a��[�`��P�I
:DL
8)a-�i�<��+E��Mq�N*v��)���a�<9$�äYb@Qh�_:������g�<نGW�H��͙۠���@ Xe�<�E$��L���yU���Z���E�<q�Ó�r񪐭�.�
�JDC�<�� Z��e��&��7����OZ�<�c��>Vyɤ�تUkF-�!'@o�<Q��R/$@��aJ�H�#Xk�<	� צ>��{��_�?Ƣ��O�h�<i���J���˒��;<�R �g�N�<� dɐ�.�X�x�7gJ=�@��"OZ�˱-��89�PBW ���a"O����dZ	9��#��4ȜQ�"O��y���.P9��e��q�� ��"O�� �Gm��1��g!�j�;�"O&�K5�U�@�y�/U�b�10�"O�t���I
q���>k�n��C"O0��QCUH���n�sH~�1�"O�Ib�M�O:�p��O0,=��ː"Ox��mMG�����>AF,�"OL,�g��2z�aW�A첨	#"O�uQ��;2���Z�B� Ҹ�z5"O��S�'ܨv��ӧC(v�$+�"O�R�M�C��S�շy~����"O`4z�É�L�
QP��<o��@g"O���V�Wh���iR.B��<y�"O���!,��lW�=ك)˳�x�U"OX �V0;�<5�����Eb�"O��{���y�\{c���S�D�$"OP5�/�q�̀�N�~](p"O<�"#ƛC�l0�K�`���k&"O��
eؒ ���`0jO<}�Q�"Oh�q@W>�p��;���D"O"}�%ȅo�d�pN�ݦ��A"O֤!�/L�bc(�P/>o�&�"O�T�ƋT2�tY�����x��"O����K.��� %×z�hH��"O��1ʝ�nh�	f$�^�T�""OlXӂ��V�K���/t���"O��)�gZtud%#�1\F��6"O8��^ $�P�3'��#� ��"O83̈#K������˖A�@��"OpK��ڨ6hL����"��d"Or:�`ѹ@�1��JY�0���'"OH�˥�?L�0���)Ǭf�\`"O^m��
 [DdEk�FRp[ ���"O�97E,XM��[��?Z�M2V"O��ª�/4����F+>~�����"Oh�s�@F�ADU����H�@,�d"O��jf,\,]~U+�/�:��YD"O���GHl�|� �J-$2�	�"O|�C�䅊J���*�hR3a��0�"OJ��o��7$�b&�(���"Oș��6�&� ��U�w�#"O�����B�~!ꉣ�h�5�>�bS"O��g̊��K7)ç6�fp "O�H��I��U�a�'��g�N d"O���/@xR|Ayv�&����w"Ov(	2.ү09*�reN�~��y�"O|@�@�1��*p�/9�HK�"On���S�-���r��V� �иt"Oժb`�;f2� c\9= ��"O6����[�0x���h�*	H0q�"O<cb ��i�l�˲GҼlb�Q6"Ot����Z�����g�<tQ��9�"O��1b�C�:z.૴%�"r���8�"O�q�(Vxؘ���_�Y�y#�"O���`�1�,K'�C�8�Ɓ��"OU��ʉ5Y����,U�2(
�"O
��T͉aG&M����"R�Y9�"O��;U,��=d��a��>9���"O 9�M�_q��@�O�W�xA"O�}F��^X-ۗ�6}�p�a�"O��nǚ2�ŢWχ%!����S"O� ��e�?o$H�BD�K�*�@%"O"T���M<���p1��D"OT<�f�X*D�@xJ$'<����"O&��$� �9���� /��@�"O�	�l��>θ��6��*��pR"O�9@c�ÔJ����#_�9�Ȱ��"O��K��]3W���Plլ/�\e�&"O��P�ʅ�<f6�᠓9?{Rm1#"O4Y	D*M�x��`r]����"O��`�j5Q�$�� �̲���"O�hÉ��uF%Ӑ��c�
Ic�"O�x��#Ư]�� ���/}��|�!"OV��c��3g����r��8v��%"O�����O���؆d�p��� "O@���1�j,����u��AI"O<+W�X-y�J<�G��+N=>(s"O|@�
��4вQ[D��!c���F"O˥`�n�z�OךNz�+"O�a��LQ*,{�1Id�tjAʴ"OV����A.�L�D�׍,vzlj0"O�I{$&��4��� ���q��1F"O�a�Ȭ|��,�7�Öe�*�۱"O�Å�0Ҷ�8b�̟>�����"O%�$S�l��d:wl�a�"O�1S'(�N���Y��7]t YZ�"Oj\��ꗿT��(���	<����"O^�9���=m�f�:�,��*�I�"O��$
6ڢ5c�A -�h=�D"OX���ĬǘE�wɏ7�v@S@"Oj��a݊W�A򂁄z�e�R"One�򯏷Mr��Wa�v�vd�"O"���A��ڇ!npdx"O� ��i_�>e�T�Aj¥Wɨ8"OJYC�!��F���uIսȶlcQ"O53�)A�=�e�bHɰR�9W"On�Д�ɷz� �c°'�Y�"O�����<49r��Ə'Q�< Ѱ"O�\���]N(@D�~.~	(�"O^ؖ�M>h�	�F�G���\`�"O΀�EEF'!~N�0F �p�8���"O��;�_� Q�TA�=��r"O������W�Bt'�� 'ŞP+�"O�h9B*�U~��0 
6�:��"O��pA�ɖF]̱��!O�yr��s"O�U��f��k���d�4��"OD-�Q���<`!1��(D ��"O��6eJ�Gm*�G��h�ZX��"O�5Ѵ�ܚl�
��e#ę̼��"O��R�̃~<����
�M�бx�"OUA`\��L�p�(Z�{����V"O��b%�9Ԉ)��h)iw~)!"O�	�������N���"O�Pue�l@,4q�d],^����"O�@I�h�@Sp����Y뚑[�"O�X����I=&t��%R�.dkt"O�D�G�DTx�8�K�,���17"O�jV �������F��m�B7D��i�Q�'2�E'A���m��3D��[���9��])��@6lg��
3h6D�L��j� 2@�p��!�"��L1D��ڴf)�|��_�쭸��!D��ZVAY�01�@�kΪVH��?D�@�%��,rjz�"��!<�
�s�=D������C.H�@D�	K(���+.D�� 
q2$h^�Z�����^mt�9�"OP�S���&��pk&ICYp�T"O���n���r��H�GEM�V"OJ�"UbÓZ�̍pPȅ� 4�h�"O$�g�O������_���7"O���e	7>�l�Ď�*��A0"Ovth�	o��|�p)N/j���"OF��%��	H��CF�����;�"O�|R"F�d4�a� C�X�p^�܇�I#k9:�y��5�fy�kV</����d9?��NJع�����g�X�2w��j�<A�&B	=��|�,)u� V�WP�<���AgU�#�eE�i������T�<��H�&EnѨ���]p�t�O[R�h���Ow�)�W, H|�hS�����	�'�e+v��
_��Px�,T���X	�'�mVK]D�����ǜ/�4P��'����1�ݿ\��)�	9T��Ա�'���A��J�h��*`�O���	���'`���C�O�$iZv
Q
B�̭ȉ�$,�S��nU�(��)I�L�W�� cP>��'ў�ON�����G�(���T�|R6؁����(O?��4��H��H�>��UX� �+q��O��ĆN�r��Aĸc��!��'�g̡��Fl�8@C��~u�B��6�j���6���m���a�M��A�B��C#Z�MX��!�F��tCW,\u��)�"V.H�$q�>ى����BƗQ���r!n�/��(
�����y�,A�y�6-��,�xy��;�HO4��D��P�-1`g,�k�V*B\����ə+XTR���#.��,���ǻz�\���,}�(L�m��b� �Z9�����]W��DF{���M�����4�ע�"M�8���	6�D5�'t�<���I�	ӂ�xa����ɆȓER�&ɓt��D�0�ʍ~����_<J���`�9B5�X2

^#RX��%��MF&+����#����ē/�A���J�\�Z�����b�'"O�����0�$��hQ�WA@
��'Q��C�Y��������R\BL�#�(�O �	�W�l4�#C4T���\�s8C䉸u��(�q`�0Z֐UPǥ)6�0��d6�	2�p�k�� Bp�y��:=�ʓ�0?��\�2��bT��p���K�D]�<yc-Q�6�i Վ��}�4��bH�p�<����=)n�p@��Qh�h�r���[\ў"~��v�8���E�T��T� :��B�I
.W�X%c�<�d�8P�	v���w}��d���O
���a.%HD���A:&M��s�'�����#�Z�����4��R3�%
Ҽ�=E��'�B �B��S����pF%���'t���Ƥ�!:H4x�G(ޮ}�
��bO
�Z!��,.��˵NR�0�'��MB@����D�
ծ ���<�60�$�
�y��LD{ʟT��È�\�b\�r�6N�r�"O6�� ԣǢ�#���bK��A�'��A�ďbP��cHN�i�����n����=1���>t�b=�'���\G�uJP,�j�!�$�)�")C��T�o��a���y�!���O�A��Euf��rF
[�:K�Ҧ��s���	��6# ]�U%����1����]]!���4W��eKC9Fo���CB�5J�
O����װg��	��ί�}1��'�qO"<���%��`�C�[^����O���� ���a�ػm��d䊗8�*�q�l(}��'(  g�"!��l���[�m�8L��'="�St�дE�V�Ҁ�^V�� ��D7,OƽX�
){�|�򰏖�YG�\��"OR�1�攝s��}Z� �UKr=Y���9LOm�'��8G���@��XR@�±O0�#�!I,������hd�pI�"D� SS�_��L!��@upT��#D��y3-������bL�$9bDC��,�O��-9�R�����N�ʴlU�te��hO?��U�͊p�!ӈ�0(�^����#D��������Ic� �3�BT˅�/D�t�w�_'�,� q���5D|̨� .�OZʓ��u�e�=R�zT`@)�$P��"OvAq�"�]>i2v��l]�e"O�Hg�ΎN�09{$�ӳf"��T"Otv���Tc_:�b�1�� =ayb�If�Y*�"Ф�0˛(?1�#?�C�"�'�*�SV-Įz���p�4!���yT*�ɘ@�WX�H����'��O�#~� ,5��Q��
�V��BgIN�<Yઔ�:��,�v!խ}Q*؉��e�<9��y� s�%���QZ�DJ^�<�6I�/ ��Er�G[j=� BTi�d�<�#u{VTY�Z8���Ӂz!��7E�R����:M��qP'�f!򤜶>��\���O�=�ѻgEC��!��õ+"l$3���)��D��$�-Fj!�D����q��]�,�&�I�~V�@D{ʟ ]+�-s�jda4	����q"OĝYE���p2�Px�P�DPN�����d� g|x���8L�n�I���k7!���u��4��'[�쑚�L���i؟�v��(?L2��a�U�6Xe��"D�ԉЂYܱW+T
^�tĂ lK��hO?���=16`P;��*:�0�i��.G�'�a|b
��l��-{U��t��H��	߳�~b�'U�p@�Ϻb߮h�fmQ�pAX�y2�O��XM<9�&L?+�$�A���D�>}J@ka�'�D�d�E3 �~@��o�W�B8�e	��O�=�O��9��枺&��Dɔ���Z��A�OH�=E�TCB�w��KY96�Z
����hO���$��t�p�)0�=ROB�b��P�b9�|��I=oפ�X�cڽ(��Ux �^t�C�əF��BTƋ$|&�M 1�86�G{��9O(��Z&!�J8�PM�70�� Z��'�O8�kB�����!�|���p2O��IdX��S�N�V�ڌhr�� X�ሠ�,��,�	r���y��L�B?@�p�ҋ&�i1���?!.O����eB(PB���%�2�#㏀$`�p���hO�n
< ]�䪇'1�H��3$�!�D��B���8(�sBۻH\�<`�"Oԩ� Ƴ>����6O��p>�x��"O�9��׀e'�,����2<8�3"O4q�FFѰj�1Bf�ЃC|��aO�i��աSW(�bA¨5�I�c�G�<y1�%2l�ѱ�N�|ݪ0����G8����ቓ���  �B�LX����B�	3|�j`ԉ��18�)����4��<E������i%A2^��q�$oǸ�y��RiP����F�
 �Ar�D۠�y��D��Yg%֓g��P�E�yR'՛C4����� �u
FT!�d�<�ĉ��߷c!b��UG�*>!��  �C�g�6�0�ˤ���Sp$�cp"O�	�@형���b,υz����"OT��Aԭ%RAy�_DEp��"OA�dI��2�tHp�M!az"O:U "@ѓE(Fx�J�MVN!�&"O|)ƍ�7^���W&M�Nʠ#�"O�)!(W*V����ΐfI=�c"ORDjΎ������"<�`�'"O�X�E#1&J��� V��"O�y����Z��%{B;bk䍓�"O61�ueHT��
\�ge��c"O��A�-�_#��!�H��D�6L�"O}`�?�&I��FɳO��i�"O��#�^s:N��&�{�4�(�"O����*.*��A��4"O����LН7��������{^���"O�����)'֕QeS(�*�"O2���KZ�t�8� m�RB�K�"O>0�0��:[�X��l�3G4 ���"O$����M�E2�y��{���"O��bv
�	7h���eB 7�b�a�"ONi�b_�vFpi
��nv���"O&i�U/g�h��	�K��I�"OH���C��\�����P}D� "O�Qx�CQ�l  \ӕ��$S@��"O��'M�?b��06 :�6aJ�"O��A��r��u�G�L�[����"OL��b�W�7Z���/�#����e"Oj1�rH�-|�J�c��3p� �3�"O"�f�L�&t4%��x�D��"O\h6#��^7L�i�
��-�R<�5"O��Kf�;z.������e�<��w"O
�c '�QZ�{ע�6��{�"OvH���Cۈ8@G�S�_�x]AA"O��"� .G��m �AM5(�6��"O(�j�+A�)>��5���[��9�'"O��c`�SJ��E�@�	}�x	�"O�4�fhM����ӯ_Kt y��"O�9P���[�*�h��� 2f��d"O��#�����Ys�׼H@&S�"O�!2��7I�lB��Z�v]��  "OFes���s~�!C��P4tXsA"Oj����8&V��K���g��0�"O�Ka��?ZaTÕZ[|hʠ"OF���DE4�b���OAC�"OF�&`J�.y��;w�z0��"O�4Y'��	+��(�#�/��أ"O��H�?(�@�c"A�NA���"O:�0�D��0��!9' � �'"Ob�p�	՘ln!�VnF�2KdQ�"O���Ɩ�I@���B엮V� b"OؤB�eL�x���r�ڱ~N*e"OḠ�ō&*DYq�51����"O����8r�:AZ+�?!Έ�""OM9LӼC�� ��3��9ru"O>��af�;[���bm0I5z���"O��a�
'�X=H�̂�����a"Ov%ㆌQ��SGJ܏�!��{���f��4,<|��b�\�m�!�D%%d��{��D �uZ$��-�!��0a
�o�.u�)J�i�!��p�e����9X���{!��y��ʳ"���A$���f�!�d��d�i�ƀ��T$���,�!�� ��d-׺,���SP@���l�q"O��Ȁ��5z�'���qL��c"O
�	��W%����!!0���"Ol+`��'4=����S8��R@"Op2�j&A�@U2k�\,D�"O��K���#_���`��$eh'"O�-�`�@sr�(�'ڄ0���"O�	ɰߴ|����L�
�ļ D"O4k%�R\D ��5+q���I�"O���(�(��9�*3'"O0�mÞwEfe�6�X[p�"O~�CnG�� �M�!�"�"O ��B��7���!ƛl���*""O�=�2�ƀ6{��Zw�Ъgܐ�ȓ"O,]���M�2�`�o��?�t��"O�ɫ�	,[�
�a$z�^�(�"O~��D'L�^��)P���
���s�"O�c�U�Z��|�v���:��MK�"O�U*�fX�/�i�o2)x���"O:�Ԯ�LȻ����i(c&"O�t)�NQ�_�B��_�
�m��"O8KR����(ТϩhW�L�1"O�� �"�8<�H��ҍ^�i1�"OlyiѨ5Eff�`��1G8"$Q"OJ���H�<�R��Ӄ� �J{�"O&p*a�&R.@`���2�d�3"O�q�$��2,:�Z @��� F"O��TE[&R������66[L}���'��d!���5��v&P-�]����s�T������6D�DH�+\1�
(��OY*@蛲5}Q������`0P�|�BJJ ?a�|s�Z�o�`HqD\s�<�fKd�j�"m\�h����7aڢd�XyVM�-"��a�'��>�ɛIq��0�Ĵ��ՒG��B�	3QX����F 8�TӶl�lr��dX�]�|,ҳ�M7n�����N1>Z1���XL�Q�T4�{�0�X(����3<��Z�e�F��1�b�\��!�C"O&	���V���Yi6B�l�N����䖈s�&pr���/U:��>���3���[2�ɆT#l8B���vW8c�O��ȑj����c�Z�Tp����~���`޽$����|�A� ~���KJ>���^�
�.q��=|�[U	@Q�<J��nej�$ٮ�l�����X��rD�ْ������I��Uc����i@#_k�D�w,H�w��!C��k�{�k[�2������ "^j$Ȥ@K�H�.1:X�yQ�V�7E,�O�1�"JC�[g���I�*9* �IV�!@�hAeeL�n2�}$�8c=H"<G,G�A��m�@W1�L:dN��l I��Ɨ?��-�T	S1z��(�Q)F��M���X9g� u
f�3}����z�Z�C�ң9њ��gԀ_ZH̱W��:E�$9&��]!T��4(�5$��C��-��X(q4��H���84�(Z��$��G�t�۠�,��$ސi�N��Û�,� �ц �M��Ɍm1���je�Şc��l3v��l��7���!Z |Yd�g����2���k�a~B����rU��=hdra����Z�'�����!T;�d Y�]�R���M�J�	h�d��g���&\�qc�<�O�I�$���m_FɄ��(r�ndK�i�����ŔL�ʘ�l��b����(�<E��$�(n�}��LM��EGʔ�0<�0n��fo��L>�$�C1Ly����t��`%�L�I�0��'�i�� ��5�ϸ'B��s�D?�
8����r�� �
��q)��O�X8�O#N.] S��
(p�x��ڔ{Ď�!dS�1���DJ=`B�0��T�S @!�)RN��!l��1H#?	 ��K��l��Ο �SP��"\�s�پ7��8J�����t(�	�������$��@�(Wÿc���c~B8y�-+�Ȍ
�0|J�P�:�jw�F?/B���k\���ꁡ��s�z��В>E��k ����p�@���o�Q$<���>�s��0-�\�>�Ofxإ E�mD��:W�}��x #V�IC�]6j��!:��ɇ\�9��(��1t%C��9lsF�P3FY2��=��'qL� �X1��=3�o�O�T��I�ZQ�� '�Zs̓ZP��7废x����L��ЦO� � �Ǉ۴8���'�#TbB �	$G����m�-��OL����o�*ViF��D.�9T^=�� ��z�&D�<�c�U����>=6@�H��k�FPg�*�5�O�-��(��Se�a�Olk2�Ё~��2����I[20��)E�2i&�#���_bB䉩����Q�$o�xL����<@�:�Ɏ+&}��#>>��B�T�IC��ҶY;(��#+^`�4'��|�f�yP.ۜ�j��0?	�n�%;4��ӤDm\л��ԡ	���F�H"�8Yb�F�=H�P!�oc�<ɟ�O$L�qJ�v�6	��%Q�F��6���@�q������څ*1^�H���\|�8��FC2b"�HW�^� �����GK�)h>,�fB��<Ѷ��.նq{C�ʙ;�&�����|�'���%@ڴje�pq�'�&:HY��́�_T0Db�N=
�ʒE���X��Et(<�%��Tq�K�.�W�<q�4hR�\X%G�?䠗�W�,tZ���(�"����߃t�b�'`b�l�����unv��p!в����DG��j��C����xU�,
kP����v��j��Q����@���~�x�11v݉jV@�-�$�q�j�.�����X�.D�^���h�=��Y�`�'��I���
�P���\@�$�6�B����Su
Ժ��<G"$E��i�����V-&��%*A����d�2eBiyVF�^-Ez��۽-�ўxC�,��TP����AVD�@���o
�`���F!C"/���p��w��({V�R�m8,�Ȝ�WرI����$\��`�y�
�x��͠�.ˣ+^"n�u� ��7�Z�l��"e���t�JR�z�����,��xg�)H��i���2u��4p���/H� �5��⌏��19�L�m<�9��F��t*�ظ �ޑ�\��&���;a�W���!��Ԙi6����~͘��X�v�
��D��@�.�Rv�'�*�z�m��"W�Ր*7�x��Ҿ��%�4fʩwH%�r�ȅyr6��`�Jb�d�L6���������<`T��0H�7Y��#�dĥv{���է+]��WJw���.�]|���eQ�2MX���FTh��Y#�.0Z���1��c�L[�ax��V$\7�����Z�s&Ɇ �ybc^�s
@�k1�9c�``���\5�	��|��M�Y�~K�"SZ6����b�&m��c��1f,0C���9�P1p!hÌ|�2�#���7W.ѱs�Ճ�?����P^4-C%r݉R�`�!7�9'��X�R���B"h�f��6T�m�*��D=K�B�[�/�4�l���]6$8��F�`c!��޽q�a�R��qp�_�@���IU�z�	�+�ET��fK�Tp�����K��]M8��NW�sY�!. 	��ּ0����\���������ڢ|�'����;;�DmkB>n��
�OF���jD�}�d��O����i�1�R�#�K�&�f��Ü�a�Zf�P���Q��F1�p>�a/��L�hAS���|�l�R��dA*;�Y��a��H\��-Vl�ˀE	-���G�6�*֢Ԏ�~{F�)+�!�ƕA)�	r�?��#���R�dX�O�7�ЭGx\	�!%0}�f��^��B�w�	��kM�tĤ���ՐI$�T���Z�)����[
Li���-��ycDϰU�*�ٕ v��Lb�i��i�3?s��p-���샢�lZ�&�g�' ʩ�&��
�|@$>剦�V���zA@ύp<��Ѧ��jxըP�@.�|�hT�b�Mh�G�>5H�
���=��䅞zD��@uʔ+��I�>���ɱ��X��'�6p�W�H�&�hƊO�dmX�5�2x�G���a>��`��c`挛�別��'���qW�i�h�JD�>)C'�/)K8�0Ÿ�e���87��Y؇�҂�>���	&!�έ���~~"B؇HJ��s�n� U�t�8�@L3����g�i�̅!��>�'��k�L�;���Op�)�T����'i?Z�S��O� �픆g^2A�)O��BP���S�i�L|z �+8��
u�T�J^v�s��9p�؈�C�(R�J�����Vpe`��v�u�b!M�d���Ѧ�$��0����Ш;�4.���'z����������{�*���A��O�0�!�	C�M`��)�_Gp	Q:}"�s��"�{�i��^Er��8���!	Y."}�E;v��3�@�>�3j9����9擾,��٨`K#?�Yk'C���vB�I� ^�b��}(���t/[�]���I�a�#�l&y��S�OWx]!B�Ĵ40��-�g�`��'�:���� l܋�\��ޑ�O��w#ɻ)���'����-Y�$a��jC��<���!�h��D.w^���ƍ��t	  K
P��Z�5�C�f�7e�"�¦� �m�*��R�)�6a�=�Gi��͸O�F8R ��
xt��R鈸]0*�
�'����gT�'�A�1҃g�R	j/O��[&iG�ȸ�(�`2���T�\$3�m��� ��"Or�ࢊ_�]����5,�,��B"O�Xj�k�i ��3:bus"O� ��#�'l�0l1�iH�U���Xc"O��j��׮Qƹ"�Ɯs���5"O�4Ysa��1�t���ǝzv�"O(}"IE�G �Y�C�r�$��1"O�)�%�'ƌP��#ؙt���B"O��@@�6	�K�1Y.���/�y�ΦNʘ��ъ��V��ط��y��դ�'FO�E��\�Cm���
,�Ur�Q66d\D��/qXQ�ȓ(<ա��]2v��lI��A!�\�ȓd��hS�%)LY�B�äoU�܇�C|T�C�m(V���*䄕����ȓ�D� DEƵU��t1�΢%�
���+2.t
��h�8��&�S���g7�<�&�*w�����]��$���l�����$���f�P(]�����6�H��]�-�neA�-�.�V��ȓ���#�D�zA���V<\$�U�ȓ!،x7'D�^�<E�%s+ ��F��X	���lҧY
ฆ���A�֓�U(ҭ��f�ȓ�=�$f��5� wB�0�����2ak���2M6qvbI8O(4��)%���e�S�BB��zC ��{���W#n�#��W��9x�膏_��ȓwz� :6��\
��&�V8*p�ȓJNr�Y��OR��6��srH�ȓK6$�y$K[Z�����4��ȓ���ʅ��O�b�C���>��ȓ+횒��_�ђP	��K�:���Vd�Q�"h<!(�����&|����ȓ nV9J5@1c��@"��xq؁��F���G΄d�~��e�/U`ņȓGN�Ը6$��[rX��ɗk)��MZ�5q$���b����*��)F���Ay<(���0/hL��#�%q]�ȓ
��i�T�Y����]�:��ȓ)�& P���|Mġ�%n�� ����k�ޭ�b,J�)��\��2��,��N����Л2pkCM��{L���ȓ!��$(�oP�r�js��/O��-�ȓS~��c�]�����&l{���4=��9�ǁ5ɢ�
r 	�#j^Նȓ�,�jp��c^����ٜB{�Ԇ�R�y4j���R�#�7���ȓ
���UBĊr�L�c%¯d��ه�`ߚ�	f��"yT��3�e�]�ȑ��`t�ӆYD��d�OQ�� �ȓ]�Hy�u���VL:���-�(q����:OF�B.�0\N*@��n�>�E�ȓT����O�+{[r���;0�Ї�]��p�2E��
�X=�¥�*~�����ݻbM����� ԃ8�}��K�iI���<���MV��i�ȓf+��g�C;GN<d;ܗzxY�ȓ��$sC�D�����@G��	�ȓGV��.^iV�2�
� ���~��]0"&�qj�X@��hh�U��`�.�J�GZ"��:�g�#��T��$�N0R K�#k�>(3,���|�ȓo,��,�,V@�� e��\Q4ć�2I�)�5*�5,"�:pi������R����� rՋ�N
.�y�ȓ�xm������S���?j"��S�? �ՃU�L,}+� J`���2`�i"O։�uo��4p�a��#^��"OX�a�B^-Mr��z�o����Z"O|�U��/=&���P�NV�Y�"O���V�A���x��G^L�I
�"Or(yƪ�6d9����* 8��C"O�M��Jq�B!����-�R�"O�����?��x��*�:0h�$�"O~qe,�v��eiH%uS���F"O�e�2�ϱ1�6��+��<4p�T"O�;�&� =�Ex�+�z^��iT"O���������'/[(�zc�-�y�Z �H�G�/m�MIӅ���y�K��:PYG�ϭj�3�m�2�y�ͧw�ܡQ�a�+e$�(�@�Ҷ�y��<�	�eN�gI<1h�[��y�r�:u�A��im���Ҁ^��y���St̚�d��i��i3�Q�yB#F0R��A�5��	Z͸Уp��y�MI G���#)/l2bĲ��C�y�a�85���Q��/X��&[7�y��J�|�V=B��^�m�M�y�,Ǥ3ڂ��@��4��������y���L����Û+"�9B���y©ܛK�a j�t@
�C�yr��3&+f%A6�ê�ZY���G�y"��,`14�h�e�#^H"U�V��yr��<!$q��a��������y�Ǘ +Jt��� ��r�ʒ'�y2oݎoB�Vz�+�!ƟXz|���U2�"� 2�{�A�le��ȓg��r� H=%]M��/ܔ�����ɿqQn�rң�䦝�qҴv)�L��@ϳSrR��v#D���%��	a�>Њ5 ��PRXB�D Kʚ8e�P�أ|����?J�>�#�ϘT��@0,D�<a��?(��p��∁P氙��� wU��b�6h*��'�>�	�v톝��E;�I�7LD
YNC�I 9HZ	��C��^K3K��
�n��U�#�(|+Q��7���$u�<�#�%�n�0�S��֡��{���;t-JAiІw�|����'ת��A��NxtZT"O@q�ił@��h3����Z@ڱ���K1��R���>Ea��R4#��	���8m�����Ț'�(M#�OH��4k�]]H<����<4��� �%;M�����:��I�|�V����(rI>��/ހJ�,��!���P�<�'J9MNqV솰7�"�.�O���df�t4s#���I"���CYj����~�$1 ��K
�|�p �D�	Wn���ǈ�B�� 3|�&9�TE:Z,��s,�,��`qD닢���d_J��B�WV�����;�"(�J<��a��D��B'��f�����j�'s4�sc��5� ��|J#C,1:f�*7	�j��)i�*צ�`��a�-q6�6�W>'�R��C���)§=�:�J��ձ"B�*��MX�Y�����Z;2�|Zw�X�+�L��-� `�OTհs�^�1����n��&�Ȍ9��˓<T�YZPhZ���g�KL@҃&I��F�q&`����D�'�HdJF��<�8�O1��I*�B�Z).ed^�s�8����.�H�5�S�BR����ɍx�2��s��+C\*�G��)E�ԤO�� �0.[��I�8sv�p��	�A���lQ6�B$�#�H%��jP8Nj��	�S<�ze�B-fC0x����M�J `��o�&�J$�70�D��\= F	����S����y�=&ߠ��V��:b�����O�r��%�&�$���+6�v$r����X���
�Q��J\��;�B$-vt%?�X2t��X��"k0o ��"H)\O��J'���?A"	Я���@c`� ATt��6f_�8<JiO2� ӓe1��'��o�D��W�G�"Lsuj�)Y�:��$�?`8d@���)PfH�<��a@C�˯\���.0�,�F{k�%k��ڢk�a�x@mA�d������n�&XR���':-�JܿK����çv4��s����9�NuY5"#����8e?:��S�ՖW!�S�O�� �QX3���6�b�C0q򯘄71�%�8 0B�>�3�$������$�?;�N��� _
��I"���[U�G�~џ�y��.,� m���
����A�4 D��bː�H��y��Q5%	Z���֪(�Z�c"�\$�"Q�ǯڧA`���Ix� 4�V��|�dL21^���7/"�ؔ��7�ў�2��M�Q�,���i��G��0K�m\'w�� TOC7G��'v��tw�S�'��y7�	1;v��r�H�O���	�s��8��gJ#��S�O��q��鋸A5��:��?n���C2"OV��d��:,�@r���)?��ȲqR�sP	�0��Z"�F�r ]�=�������$x�E��c���}���'�:��`H'��t��GN#_,�r��]�FT4;�HO�{�$�Ւ|��s��#��/j)�����r�*�:EJ9�:`\���6�'}�����l�)�[&���^k�����ʔ�b��d d���'K��j���)+0�8S毘�+.μ!
ۓg���ՅD�3B�����>ex�B�e�-�8݂�ӠT��Y��'�F��M3ORy *�$��Ts�{�Ksy�	Z�▞n͖e���@���\�_j`�G�\�a }�ŏ7G8Pm�R�FvH<)�a^�_�D��'�9^����p�V�V�e��	�(���%	%bM�;yvM:ab���Ok,�"i�ѹ�
,~ h+し#�!�L�*ϖtW ����%֟:�ʌ��,�v$-�1\Pv���O��K@�	b��8��O
�[�Æ2&P�pC��R0c��%� �'�����,+t�$�{`�\VX��##��10���O4^���e?�FO��dg@]��j<O6� pJʽ9u���@	w��t���D��[c"l�� PX���������A¿H,�2���_z���	�<h
x�Bȅ8f��х�L��q��	�Q(5&E�sֺ���(������`@��VeZ,;G-K;L��m��	�Y��<�]��B��6k
��:LY�oւ?#�C�	p�ڝ��O�C-ï=&��	W]Z��d����1�8��CB�����gB�	Ȕ�摟�{�3ǔL�H6o<��B�H6lO��-4Y
�b�$�d�\�bG��^A�[妓�ty.�b��>bN�(2���/+�ax�ӅD`��t�׈����e����'���u�_���l1���o�$|� 8�F�?[j�ySg���9qwm�9op���q'v�@���y|I��"�
=��G~�c�|��ػ��i�4�tٙ�,ژ ���Q��m�!�$���Xɓ�V#Qc��*��	2"\1`t�čTЮ�B���lC��A,�]�������UA<C䉲~+ ��(��_�\�����y�=�����y��|�'x��
����;�Š|j��Ǔ$h`���0�ɸ}�@t0+��&�05*��)p��W΄�p��,xr�'�qc`I�i�	q�,�H)�O�2tB\;7Z�O�"���8=T,��'�����kp�b@����	����'�n�IC��/�uA�dE<K�řS�&}��i�" ٷ� j�%.�m`r�ݼ�$ț���a�$N�x,�1h�g�a���D��"���Ĭ��D�t��f�`���۫A˞�'����_�R�����_vr���W�wp6Lk ��x{��?�U�RZY���`�!�d��0����H};2bn](��Y#$@(X��e2�Oܔa�I��*�7 
F���Z� �t�ރ/��>v�Ⱦ\ r�'Gh?�f4n��)0�K����:�%�r��,�FB��h����a���&=�[��%�� ��>��D��M{ҌZ.��{�6�`4��4�u�j��T�𗅅�vITE�#N[���O$�0�Ǿ..�A�m�a���v���g�.i�l���C)�M��Q������-E���g~�Ï�W䖍8@
�b�)AW,�~�,� Q��	�0IXy�ʜ� F].46\'>�b�֎/�U�gȨ�j���(#d�������|��?$���:��K�>*4������a��H�0DJ�p��O_�m�*���,�4�:��H%5��8���+"�Y��	�h�X��*�3n��SmB�+#��3!^�QÖ>�W8Oh�=!$a���ۊY�V(�Da:���Df��&�Q����+�H"�� �)�;j�h٠<*<�9GOD�!���d6~LG��w2��e-�6��$Z�qވ�k0��.��)ڧz԰H��e�
�j;9��0�ȓL��x �'��=S��'�p�OB�K&J�1G<��6�� X�gқg�4�
���L�i��I:m�ԔJ� ǳJ�nP0ʜl���C�%Zl�|(�Od�aяڃ1� <���Н3R����I���1G�Yd�'�t���w�H�c�Vm`���S�? �|��,$�2A�W�[�^*��ÅP���$�޹n�qO�>�"��S$����Ï�H&��"O�d��j�,w�ň��ʠ"Or�a��ҠC�pRW-܏2	,*D"Ob�h���u�hi3,�:!�dq""O�di4�Ǔ8e��b���"d*�"Ob�� #R�z���l��(�&}H�"Oj��(Z�A:EЂFK�I�:0S�"O�(1�*ɭ@F�CīB�|�F�e"O
����B
�V��T��.^�X���"OaH�Snp�	�Yt��{�"O�t��?E	ĕ�Z�eC�8�"Or� !F;*�Ȝ��.�(M�HU"O���CB�@�����N�!��)�Q"O����f%�U�G��j�4�r "O�@����$�:d�U�Ր}P1v"O��p�${2���1_f[�"O��vc�"�x��S�"BP��"Or��Ŏb	*�[!gU
G�Q�"O��.��q"�YçG��kE��9 "Ol�Rf(��1��П@6���3"OR��HüC|THR��&��EI�"OD�֢}�>��M�2����"OB��'P��HB1�RF���"O��K�'��wo���CF׻a�F��"O\�b"�.W&=B�ˌ�'�]��"O��RTn]�lUb8C�œ,rEAB"O��u���r������,\8����"O���S_  ���BOǎ�T"O,؋Q�J*QD��%[�tD�%"O�Å�	�H=��ū3�8��B"OR��NV�[Y�;eH2X�=�"O|����i*��a�|�"�PC"O�y��R�r��8{%V=�0��7"O��1f(I/p� a+�恡�~��"O:=9�Ï06Ҧ�SG }N��3"O���3N��A�*��ņX��"O����(�A�Bȁp��&lPe�W"O��臜k�U�w��#]��A"O@��h��;��ݏuI�JD"O�a)t�
�J��Ip#(�>6�Yy�"OD���bn �����HS.��Q"O�	pd��2�6��ଜ	Y�>���"O ��#C�(|�9J�K�'�:\�b"O 8�C��]%(DR T�`�0H`"O,�0���$�A�-��	��"O�q����F!p�tCA	W�P9P"O"l���O+h\�Q㔹{޴�"O�u�����l��a(4Ý�$f�Y��"O�h�`��T�&��EhE0�"OH�h�mI5Z'$���S�wT 
@"OR���Ȟ��H�����ED
��#"O�9S�	%]�2Pb��H�fh���O�,Ⴈ�A�S�D���	
|�krK�?�>��$�_<T�L)���W=&�V�$����԰z��ف��߶A���3�R�!�L	���ݝ-�iĎ͡=B,q��S�%�f��qLQ�WT��q��W���XbIF+�!ae�ֺ|y��+�8�# Z�"�6Ix�O�!��a`��:��"�K��VU�6W>1�O�����Q�(���f�F�2����y��M�ӌ��^S��1������Ot��ሯ<nn���%�G"�ZBGY�z���+O1��J)��8qCbۈ`$\�"Ϛ'.o�鲤ȓ7%�ɼk�������N>��@��]T~�yf�Y�]��lZpf�<�U��9f`t��I�����Q(�'�JlQ�wEI�L��6��n9����V�~V��,!jr��Sn)�!�sK�*ոqh�*K1+���醢]�?��B�;��?�\
ыV�,�#&���wL������%�:i���)d�� �1�����,y��,L��F�94��y���b�K���7b iR�%D�0��Ɗ<�e�@N
KT��3b/D���Z�k�p1/H�s�ja$3D���E癑*]l�ʷD8���u�-D�����:6�r7�vt����+D��"G��3G����,h��)&4D���eN�9��X�C�<;�*DV`1D�x����y����혟��Q���/D�쳣e�=*Cr��ㄔ�<����p�,D���p�"0 3�l�=\i���#.D��ZuO"Æ43牕�G}`�#�>D��X�C�f퐍��N�� �X��;D�D���G=(D�5qtV_��S9D�0î��k�&�ڄAR)[U�k!h#D�l����p�=).�(U��إ�-D���Ab��6@��VmC$vLb�$7D��AĭΏ
<.́@l��> 4�3��*D�|r���!���VÞ�^:RI�5�'D�`ѠNBdJ����j0m���"D� @�W3"p\��%����$iB�>D��qs�F�୉2�BL���e:D��P�f͊&�ر�����;�,.D����f˯r7��-_��{3%(D�� "��:� ���f�6}�:�8$C%D�lc�������P�E-b���$D�tc�fM�����O6�����yR퇦^�ҹ����_��(xrM_��y���_��r�U���1���L	�y�O0(¹F�U� �4�`dK��y�헬]r��Z�.�rGнJc,O�y�Ԏ ����䀬l�6٪G���y�7{��a���?f�$�I��y�D�A�28`So�a"�+�U�y�Ok�pu���Y��^,*&���yRE���~�aH�	O��]�QEM��y���g��azS��#A�n�ډ�y�/('�~!�d_�;�p�eb��yҦG<=qI���	j��dC���!�y����=�qA�֎�hiDGM&�y�a&R�DX��Z�Y�ɟ��yb�ʡI+�rd,9¥L@��yb��9n�`Y.�� A%-���y�AB�"�X�%�-����y���!]�E�o<cx��� �yR*U���B�I&-˂k��G��yBI�&-��E���*�6ݡ���yC���Y�����-[& \��y����m9�����K(���(�
�y���N��[a#	t��)3�M�y���
,�`P��WXJ�X)T+�y�AVs�	��*��H�V�駩Y��yr�"0���U��l�!3��A��y���(�托��	�0����/�y�d�=I��엶x�x����yB�E�-ʮ0y��_?�z}���y"d�7E��M�`��dMPd
v#[�yrA��	�2�X��KX�J��6� <�Py�:��iK��۬� "�AV�<AǡQ7��X����7
��*�DM�<a�h�9,|�L�eO��M��jE�S�<i��-6�D���Ò#y�+!��{ !�Ć!Bo�����.�z�g�Y!�d��[[��h��"pP5�UFD�[�!�� �๡��6#������tVΕ��"O|ب���7KL�0*H�CX�y;�"O��c%�(L�"�Y���cMf�y�"Ot��N?^�X+�,E�T�7"O|,)�E��dH���R�S4kmpdz�"O(�A'Fj�� ��'̀Fe�\k�"O�q�O!���A��	S-�|�B"OT��#�c�j0b�e��#"O$�`I]3VxQbG/��t<m��"O����A]�G�h}����d���"O��8<�)��KI&-�����"O�=�-C]6r�I虶Q�$��"O,��a��&9�8��WI˰ �0"O�\�o�`VH��kA�!��)@4"OP� ��2,��قSj�>t�Hp�"O6��E�#.�x�+�Z ���"O:�rD�)d��j1�T����R�"Oʼ;�%�k@RQ��'��	x�"O����/�9
&��h������h��"Oڔid�f�D#��;9�k�"O��* N�?"���dܹ�� �"O6��LӦs�X�0�ҡp�� H�"O`����f �l9'`݈G�����"O I�5c��.��x{ o�;(�|�B"Ob�IMA�o�j����K��d� Q"O�`ZV��1,���BY�EYΰ[ "OR`0p)��.Ff���Usn~�d"O� xc�B�`E�4��FS&]^N��U"OL�1sG�s���H��0x�["O��Sf��8zP$�Da*����"O�9!�/KbG<��ƌL#��q"ON�$��8���U�O)3�~���"O�F��>v�2��Fa�0m���E"O� "��߬^�ڵ�$bQ�I��s"O� �3͞���=�a�ӹ|���"O�����=W��D�v@V�|��Q�"O��[`_�&9l-:�EC�#(`1"O>u�d�V'Ĺ����XV��V"O�!� bζ)�-:�SD
�!�"O��2�k���J�`�1BcT �A"OD� a���m%E���0G�Œ�"O�p0D䛝*���
��-F9"O�҇�
/=�`���C�?L��1p"O�P��d�J�� X�y��S�E��y�`��PI!���,}[ ��3b���y"�N�4l�� �SL��x�É	2�y�'�2��(Y�ȍ�G�lу��y���p�P� fJBF�jq �;�yb�7eb�
QN�5�Z��'���yb(s/ rr���^P�QWFF��yH��y�������
R%fY�Q��y���"9�������Z-B���&R�y����#j*��2�N�^�>P�5���yϞ�c��۰�O.[��a�N]��yRo�]�I+�	CU�k'��yr�A�@�|ٓ�n#R�
����(�y򠌖=�8B!	<Yi�HjOF�<!�M_\���"`��,?��ڴ��T�<���M�a�z�i���jހ؉5��S�<�� �v�l��dmW�_��L� �W�<)��ÔK^T��r��>�J*�K�<a2iֈ_��!�! ��G�@p�f̘m�<q�K['U��E��.ڨD���dk�<i5���*+�풁׌O�� 櫌i�<� T���"];��5��A#�����"O�@�b�T���r!�
���"O>\@r��HO~�)��l6��"O����,�48�<*��:GX�4"s"O���qI�\W����!��z��%["O��0&�_���݈Rq��{3"O�� 勁=5��I1�ejc|%av"O���f�B[��ի��ZUVc�"O>�+��[` ��E�U��M�2"O�T��#���9(D�(V޺��"ORy��MSWh�HBھ]��p�"O�V�@�=e�H;�!�,� ��%"OČ� ��X�Uj$`�&�2JQ"OR�� n@
D+R�����w�`��3"O0���+e20��g����qٕ"O���&��h�6<��`m��䋳"O0�� ��d�@�6����[y�"O`�qo�O�6	��cU?f��;c"Op�؀�X4v�۠!*i|��*"OP��H��7�qi�iV�O L5�u"O�IiK��A���U�s�@1�E"Obkp�2^34�yR���غ��s"O60s�gʼX,fL��@̔���X2"O*��e�30��x�Ǣ	l�)�"OB36.P�>����Co]d�Z���"O�i���$#��@�lܛz��A1F"O�!ٖB�&�j�;��X�v���P"Oذ���18-�$���̨"�
xau"Oe�S�RB�6�*ǯ�#e�,1�'"O*Y�q�9LT"�����6App#�"OF�*ߙp�<���T��hC"O|���%>I|9����1?��F"O�����<�]�a�08b��c"O�T���3)��U"D�9���"Oī��]2/�x�(�@��Y5�eK"O�]��ETl�Btb�K�0�I"O�)U��:t��92ӎ�C�rM�W"O �@�#[c�R�ɞ$G���"O0�����A��p[��ۄV>�Hqu"O����H�
L�M�cF��~*��2�"OΉAԬ� �DP@�]�fy
�"O0A���!#0���g؎
g���"O�(Bao��>z4�JChʊj�v12v"Ob@��z�	K��t�!"O�L"�H��F��U���0o�x�f"O*!: "øT��9�ː8'6.��"OD@�!X^�q��	^'J��"O���Ca0*�0�0	�U��0xA"O���] 1	�H�`B	94�40�"O��Jp̚V���ۀ˖F�(��"O��{Cf޻>�����J�>�n`��"OD��.<s(y��M?/rfJe"O���B�W�-a���AH�)LA���"ONy��
�}b0�&��dA��#�"O,�z��O3/��!򇗗}j�'"O����ƫ6��C��	�JO��ڲ"O����
abtl`2Ƃ�f/$\��"Oļ��rK�X���a�;�!�d�8*�&y&k�Lb�`��W��!�Q��T��iR'X�da����e4!���_{�(�B�
)+/�I����?"!򄙮8@�4�6%�V8�` s�а
.!��-hRQ�#B(	����Ph-!��2KJ��WЂH"�S�e�=D%!�� � ��نo)|�!�B�0gU4��"OT�A��8h�Ͳ��A�(�"O�m�����#!�}���~$N��r"Ox�AQ匣~�b`��fM\�J�"O�� ���$�4b��м
�Q�"On���   �P   ]
  w    �   6)  �1  /8  p>  �D  K  �R  -Y  n_  �e  �k  9r  |x  �~  ��   `� u�	����Zv)C�'ll\�0�Kz+⟈m�R���ɼm��D�	G��P�Aç%�1bFW7IH�x�E%0F������e�X��!x�-���Dm:��\�$�Y�'i )p�
hUѳׇ�#9������#N� �bC��!iǄe+��C�F�Z��D��*��
��p�<`g�W�mxt�bT#B�+o���&i�Le���џ(s'U+ST,�ia$�9�M�U�ɜ�?����?��?q4'�3!����\!j`q)�ƅ�?����2�ꃶi��Iޟ�b����$�O�L����D��0�ȇ_����d��Oj��c}�\���ɤ9]j��~�8��-?�P$�"���ch�N[
 En)��	�<)t��@0j����!;������v}r;O��<)�kV�ē��d���T�T��j֍i^�Y��ʟ�������I���韔�O��./�9:��E���1��Z�Q�҈xӲQl��?Y�4�?R�iv
7m֦��۴�?����?� ܪ��-��1��۰Ua�����#�'f��h��:?��3&��%F4�YG�r�!���B��#�e�j�l��Mc���RJň>� ���҈5�j�����6}C0�B�x�6 ҌQ�l�&�̈́]_tQ�!�ʦ������mz�6� 囹�ڴ%����Y�<���;6"K���I*t�&g�}j�4FE�V�sӠlۆmI$1�D�Ń@&{��9�
�7u�4��Rs�L��o�z�^aG�5��mb7�Ŧ͸۴3Z�Fj՝m��ē� |��+�L;z��ͪ��\�B���� ۱<��h��'�n�"�hƚXgYC@�EF^���'��O��J�U& ���V�S�p�\�21�Z�["@�Φ��ݴW֛&�OM���8eN��J�i�
(�"FʮQ�l�����~[�!���Qw�'�L��w�'er1��`Pel�5~9V��A\_nh{�����Y��ّH;:D��(�<�G~�J>�jD��'1
r(����$U��y� ��L34!B!o�	/کh�
1�c޼��ɟD�'R�@#Di�m�(�a��%}�"5��?������(� �9�J:'X@�	VJ�2�f�#�'y���G~V��� 
�
p+EH��CLb�DV0K>5�;$E�D�o��c�Z��!\�j��ȓA��`�2훊?�-@E��iU���x4�6�R��ܻ�)ѠoM�ȓ3ؒt3�	�*w8P���H�s�R���*j������s���J+�?`���uZ�#��G�Z�.���`��X$�������#<E���A��=xph�|���豥Q��!�D���MчN	"��E8���}�!���q/�R���Q���h#��!��?#4��bÃ/
}z ��!��B�!�$�5+�H(�4���o���U�U�b:!�d��Oҡ�`�֧6bf�aC�q"�I�%`$����AlH�ǐ�LDx�C�ݧ!!�DўQ��qp�M�.AVZm��b��\�!��A�k#R)�&��r4��	"�Ć�!��D�9�`ԥo-H%�я��`�!�$Y�R��Pi�������`��{�z�$���O@5csk�
���+e�^*�
ع�d�O���/.����O��$ޕ<��(�Ai�3��\�1���ߩaB�	(���B@�>6����8O�ىU�_�:�&%����<���bD,n����.�vd��$�:I���?9�[��B�4H����'vL;�R�2�2�C�N�)p�A+�[�����'�1O�pb��B��@�M�>XXd�p��d+�S�$,�OBp�I]�)!����eM�fA t���'���<ZF��o#�D�']��?E���A�T��a(A�-�e;à
_~Bg�)7��=E��[�=�P�#f߶k����k[����#\��e@�{����]8�(����m��)��)Yv���}�>���OX���c>��3*��a�����8�����E2�$�O���D����D���[`X�y7�	�h�J�'��>�D�Ҵ�. �xJ�u�J�d�<A������TW��с�2gD���1��R��(��q����H�Rn�8v�|FybۯKv�S�4K�̤�/Q�;�X]�g�N�rᚷ��;$�R9����������NE۲g�;O`LL�2�S��7-WAyR"J�?�����?��3���&�\�I�d��6�2E0���?�,Oj��8�3}j�1Ym�l���!.��A��2���զI��4���|��'��[%%�HU�GO@�T�2$*�k�1�nu(09O��D���B�3��<S%��N�!lD� O�IR���}�����C<���w�է$!��}r���ܪ��H����K�Z�Ӥ�'����dR�T����) }��	Wb;J�!���Ɗ�sO�&I��<`���[��'<7-?�D�8m�4x&?�@�� :����A�АAk`�O˓�?I���?��b�r,ss�!S���E��� �i��U\����WǊ�(��6���z�%�K����A�X;l���p�(X9j R�����v�1�M�)��O�Ha�'�B��QGj[�R��`��ʕy�|�
D�4��Or��d;qh���(!��9�jӱ�ҏ�O��à��J�(A�b�N��4�'�ɳ7VV��}�O���|9^� �:O^"�������O�j�����;���T.B]���X��ԡq>��π�8��-�)§�P�,J�R�T�����(2Ӣ-�'�*�8���?�M~����π�ɢ=����bi���䓘?Y	ӓ ���Z��Lf04*Rh�)�.lG2�&�'@��h�6/��䉦i��B�l�4�?�.O��Q!��^�$�O2�$�<� $�Ii�~�r��s�� G� k�H���1��	K��*+���ɟ|�I4G� �#��~m��$�%v�h�Y!��+	Nl�闡{4r�sD�(�O�-Q�U25O� ��!�I�-��������I"3%4��	æE���	�?������,	�#G�;G�e�ç�5�>�� -���~��
c\���c�,=�+�^�?�����	iy��'����'&�ɈWG���L�#���+ӅV�v�D3����	����	py����k�Թ�d��9*���W)]�r�B�͐�\i91Q��o�)q֭*��ja��aΚ�7�H�2�AN�K�|3uBU4.���J 	N�Ht�$��&�/��O�$�GVN̒A��NM&���Q��gmB�'2���$§���2��,qY�4����f����Ln��%��#�0@p)� ��%�̻�4�?�*O�5Jb��}��\JP�'o)��(ɅC ��<q��?���Ԝ�OV�0��c!'��D$�pr"��5Niޑ���[�z�p���.џ�`d�8YQ4u��Ȟ�`� �q��J�0�u��06��52V)U&�E�lֹ�?1�����w� T���S,P���K3"�$T�'�b�'YL ���$otlA�[�a3�����2Ɗv��1`�YR�$�����?�-O�=9R�V���&?��O�®��?��|@�	])��)r���F���'�v��J��2h�yɖH�/�~���0��=����[��E 8��}�#h'?1�OD�Aʡ�@BjŰZcX��?���;��F�� ,�!�'�#?�i������u�O
�n�4�b)[��fy�X0b��x!�D�V=������Tat<��� m�џ���	M�B���q�X'��� 8�Q"��i�B�'m�Ƕ^Ќ�(��'�r�':�&��Pa +3���"(*l�<�C��)q��@�֦�fb@�qTc>c�h	���8Y�R�2�Bߞ
>8�ar	� qf�V
��MCa�ɼ n��|�<�1�J��nLR�Ը ��(�$�
��4�'Fn�Y��?����')!g�Y>����d�^0v�R���"O(\1�I'e� @��i
Il�a�W�����4�:���<IÌX���!�c����`��.E�`���?y��?������OD��a>݊vE�P���;�J�uo���ӶoCPq��E�C�Jd;�dĦP<����,p.�EJ�Y���QC�L�q�p� �c\�->h��H�%px��ZS�'��m)C���~�x�A�)ӛ..uC�у�?����䓢?����'�¬� �@�#d�R�3cPp��1"Ol���J#Op�P
�k^jX�I B�|r�aӲ��<�ɩ�~�Әu�b�H��Q3�t@1"��[��C�I)��9��ɐT�d��!��; C�V�µ�6(��5+�)�S#�w��C�	K��0�j v��Q ��4��C䉵s�
�G�'eJ��Ӄ�m۲C䉽B��|bQ%�_��ŰV���^t�=)�@O_�O�F]�0�Ȅ&��<�u�ը�2Y��'�nIБ*�+xL�̩E+\9���1�'��U�6��1P|{�-_���̓�'�ƈ	�(,�%�_�A�'] ��d�Q�eؖUJ�&�3}v\��
�'��(�gGτ2�����./v��(�� �
�Gx���_)��t���(5Uɣ)�9$B�B� P�)yfN�+���!Ð�8�C�2$��(��~��{��O;fsB�I�4����l��/��C�L�-��C��7w0��L� Y����X0�C��66��cҬF�:��q۲/&_�^�e>���	#p,m)���؁��J��5�C�)� �P�#� �/M@	0֊ T���:"OH Ȃe�[�����Q�o�8	�"O^t��f�w�T8��p�n`!$"O��� #  t/���v��j��f�']�]��'��"䁀�F=$�R��	�N���'�P�2���$Ax���$�G/Dԓ�'����ŕo^�XAABǣA�>x�' 2��W�/t�i�Xi
��3�,D�����W<,��8��a\�9,�D��)D�(s5k�/ ��u��M�����*ړU5�0E��GQ K��!�<D�<�Ф�y 2P ��.J'9y"�C����y�)B�X�	�NO4B@\� �/�	�yRc��t�T��%L�7΍��!�d״	���c4�L-"��ħE�d�!�\BFA
�n�1l�Lʂ�X�ҋ��O?	I�%�J�0c����D�͇v�<�r��5�����Xx ���2e
p�<�S�U�Xiģ�
f7�e��&c�<�e�`��M�C��cp<!�"�Z�<��f�(j��=kPl	�[�lH�r�G^�<�v�Y�)��	膃�@�v�*`y�Oı�p>I�OG���Zq��:Y��tZU��[�<��#�!["b	�C5Ugdء1#�X�<�G�����q�/N&��I��j�<�4GҥW��%ȳ�ʁZ�;FJp�<Y��	uJ���F��!� �ac%Uex�$��ʪ� h���4 �R����dzdc�I$D��(���Bg���᭄_�D0`�#D�����<0�t����i��?D�Da�ɂ|��K�V�w�����8D��k5�U� ����+FF��7C5D��!�ֺz�IP @D
��rWI ړ~˼uE��/�3)�<Z6�5
:�aF���y2���:�n��	�%-C�5����y����GMPpJT�V"RE�dP�ó�yb�� H�e�v D�N2^4�d/��y��%� ��s��Z݆t���y(:hO��٧m�?VA�tq3B���?yT`�������� E�d��Gձ|�xR��)D��35�<N���*S�U�apDl'D���AޭJ���*C.T=#�@�rH$D�j�gV�nS��B0��S�ع��!D�,�1�?OJ���U�(�L3D�\Z'��8X���FO�@"rQ����<A��d8�8 ��څء�(��r��2D�xkѪ5u��  ����(���3D�$���<I�x`!M�R���)r�3D�D��, t�Z��B;����2D�xqR�R0v ���15�X����5�O�y 6�On#~0\���E�;#X�P`"O�I�䚼mu`X�cڸ3�N�� "O�Kw(!	�[��\��p�F"OZ������������UQ�"O�(���F�X��İ��<=�TkA"O��j562T�j"@�l�yʐ�1?XD�~��K�~���iU �N��i¤��<�Si�>;�zt�u�	B�8dy��v�<)p
�%]����JšV/|A�&�t�<AB��$S���(W/��`0I�K�w�<i�L[�x�d�s�N5@��5s���g�<a�0;��Ƞ�jͯ踜�HP۟�H��3�S�O����S�?K�����K�-�~�3"O�QX��ܵ�r�򩒆���j�"O� x���x��M����76��p"O���NG:O�h��Æ�5DP��*O�@[��
�@�!��A�5����'�Y[t�٩U��	�����HK,O�d���'�m��'	�^�th��Ӣ �D��'�Z��4f�)h��N�|e P	�'2�t#G-E�UfJi�s'�w$hU��'�](�쑍A�������zͦ�`�'Dhts�f��kנKs�ۛr���B�*���-�!׫�`!� C�Wp���v���"�)B3L��1	�h´�ɇ�=��A
��B�xV� �f
��C��i��Y
⃧�&ZK�PO�,e��Q��d�7��3�����J�;��D�ȓf��5(�L#kĊ�Ru�C�-d�D{�M����hpJ�'~������t�@C"O�tC�Jh�̙V��'\�P�+C�<Y�e��@u���4�pYxp�M}�<yC�Υ/LL� %��2$�#u��S�<��+C�wШJ�Ù�r�jI�Vz�<� �¬MiVGٺ��a#"���
�#%�S�OPpIe%Z(�̢&� �?X�:�"Ob]q���\q�j���536��;"OH5@��Q  x�w+�_�Թ��"Ox���ޭ=���0׌��g^l��3"Od�b�mٜ ��(SLϟW[N�i�"OR�8��h���u�$�|}��P�\b��)�Ol�����ΨR��l��� �"O6}��B��;[�<cP������d"O�(�n�'y������*}����"O`�  �,�V�g���E���`W"O�ec&G�*F"��h]/|l%c��'��ؘ�'6�8s�� 9��a�s �����'`��#�#F(�\���9{�p9
�'z
�"��i_~�*�`W�cƎ���'����4��(Y��R�-��cP2�r�':��`$HN-L����	U�)V�u�	�'����EH�=>��!"��
�V������C|Q?��CS�pȐU�DE�,'@����5D��֏�h�%`�OE�n]�Ӌ3D� 	��0�	p�-˪R)H�`3D�2�lQ�hA;��)�b9��,D����j^�cp�u"�D���ac�.D������)S����'"��b�C��Ora���)�'#�(X*f扛,0�N�L��ܻ�'Єt�RA
G����Õ��RE�	�'
����׸�M��Y�1R	�'=2D��-��o�Y�ܓ	�t���'�RM�@�� F�h�`�cW�oB`��'.(1��+ӯw��p�4괰B,O h�3�'dfJ���+i�����C>,��QY�'�07N�4��U���+����	�'/��,N�`Y�� .I�$���K�'Nd���8X]��p�g_��y��'��)a����p���Q���.��]�c���K�N��djՈ�j���ȓ$~ДYT�I:�Q"�r��݇�!���*d5h�ѐ �7 �Ňȓ���{&�q�<k��N6R'�a�ȓM���!�ɗ(6�a�C��I��Յ�M>tI��֦X���&-��4@�E{�(�,𨟬�$.�D謙@���o]�,��"OđJ�旻 �Pc�ȑ 6�a+"O��v�A��0]j3��+b�8q"O� X��T)١"dh0�e�)bq["O���FT�y#6H�'+�l4�#"O�)�E�F�e�V��$e̞A�Z̒P�'��I����Q�6Ƀ�ȇOx~�##Z�r5���F���H���X"�`ġY�]E����>�tQ�$/�<]�Ӯ��ZS����\ ~��soA|{J�#�])>h�X�ȓA�t��	Ji�)���fX�U�ȓ}��\ �ٛw�Y�E�ݡ'���'� ���m�4[�$(U��Hg��i��ȓGR����p�9Ǚ 4����):~d
"o̖g:��P0��L)�ȓ4�0�N\�(�Q�ѧE���ȓJG�3�Y (d�|����F��5���'9�	�O�՘�o
7 >��)RA�6B�ɾ9�$ذ���Q�pɐ�>K�C�	<SJ��2� ��FHM��,4M�C䉽,d.�8Ѓ�n�L�	�a_Y��C�	C�T�IRH_2�"�"�}��C�	�M|ja��l�!x������ l$n�=A2��`�O;.�Zub9���)�:�c�"O:��sm@X%��A���j!T"O�(G��� �qoT�k�B�c"Op��7���YXxv��X�{"O|t�m��;�ju�L%0���Rs"O���U���`���S�*,G4 9��'�DT���S ~�Xh��#F?$[�`�}BȄ�-6�lE�ȸl۞�X/:��"O2`{�bSגE��*	�~|�Z "Oz�ʱ���klzt)�&P�X�"OPi%ϔ��|���M��LI�O�iY�y\��C%��[s�i@��O��z�^��:��>Q&��+V��֣�?Y��q�D�T�[�w7����U^�Qc��U*B�����?Q�n���V�IHQ��tk�A;�e�x�	�f�.-\9��*Y/w���9��4�)�d|�F�A0_��&�%�=c�����Q��\���ڳ�д	eHq#�I7ʦ��OZb>�#F�Z�s9Bp3ȕJ���h���<	�;�`9�T�<��l����&vDY��	���$VT(� 2�g� <��Y7/c��I���y���d�O�ʧ|�:���?A⮆�4Ŝ���16f���"�?�S)ĭ~�T� ���iH*%�����-擥I�|![��Ɲ9̼�	Fd� �R�	&b��`��.F�p���3�H|�O�D	�go�6��2"�\&bo0e)�'��j��?��O�O��I0�t�!�M�F@f8���Q)�:B�I(W�1�D�.���1B�;*��=���5=& 9!@F4x�Ě4�۟}����UyM֏h}��'W�'��?��2	f$n1�䚟l�b�K�L�a��=|E�u)�(1�v�'��'2����I?T�Hۆl]��5�7i��$J��)Y�
%��+��)6�	�3 I1�֫Q�@y��@�i�*�T���I͟�D{r2O"�ЦEJ+�U9�@;�� �"O��aA�V4V�C���C�:<�R�'+�"=�'�?+O�aq`�ZNGZ@+G��.�c��rRxM	s��O��D�O���ۺc���?ћO�h7@�!Ȟ��f*��7"�qz��ѳi��
���V��I8q�<37�#?q�b�`�{�g�	.3��G�f���4YH��<j<Ya�	4�V��7w���րIl�X�V�)_(�$;ړ�O4�� ���\�2��R�y��T��"Oa����5)N��b�M�U�T�X��4�?y-O��Qf��O��yF�?��#���	����,�2�dYKy"�'���'=`E���N�v}���Iʣ?��0�Ņ񟤹��*�vAh��C�_���� �Y��̅ 8�p
p&Ρ7e���Ӆ����6����ab�$">�@��ӟ���O̧��h֥yՠ���&�9#�t�'�a~�$.Rf�� ,��?�h%6 י��>��_���Θ�?��y���N���򰢥<i�N�: �VI8j�X>9�0���?���)@��D2d �>4|^y��
J�O��I kiZL: �h�, ���Ńr�6�C֟�b>�Սг`Rp5���/��)&Ce�|re"��nNY���O�TĀ��](�H�E�4'�5��Ч�/y��$P�2O�U�`�'�������S�? ��)7Ú8i�ȴqE��H�
mr@"O��牛�!��3�Ɲ{���C��	9�ȟ>1j�P�� ��S3`D�1ځ��nJ�$�O��i���aX����O"���O�5�;�?��"
zU�q�a�\�x�����Nzt�$�'��B�Y@�x˟�\`�f�%J(��퇫'P��V�������O�eE�8���k�?#<���9w^��V ���!�#��n~����?���?1��8��*�ϝ�4�$0���ө=�PG*OP(`�iA2~ȵ:�V�AB�	b��f���Sٟ��'O�q�,��v��qd!�-j��	���U�L�i��U�8�'Ar	qݍ�	��'1��#'�Y#`	���5L� o�����Gi�2�"Bl�L��%�'�n�Q��H?�lU�u�D-[t�������Q���j"��&�',O��˳�'�Lah�a^�h����F�a5�$R4�'n"�d/ڧ=Ͱ�#��Lu%J%�ܡi��a�'�:M(W
Z<j�E�W�N+�v��*OVDl��<�'&B����~B����$⋔kh	�u�TQ	��N��?9�+��?9���?��d�:�f̟A���@��a���ݖC���5��0��C"Z�����х�C� w+�9t	��B��T �bm��n�j��6L�/�̢g�I�aY��D�ONc>�R�E��H��5�I%M�p�n�<���0>�&Fك_��ݙ��ӥw�����@x��3(Oq�5eW��Ha�'ڿ^��W�����O��D�O�?��'�(#��V&`������Ld�0��hO�� �b��N���V:h<z�3��$G�s��'ɱ�.0�7!h܈�p���C| 7����'~�H���<9QA�Qc*�y�k��}ź6�.̈��kN� C�0}BG>�Iϥpj��:�,������0NR�\�H�8I�'\�>�I�����6c��d[����ԱX�.��'}�'3}���ɭ��)ǀg��dA��4>�|d[0� ��/���	���(�l˚m��%m�pؠ���?�6�y�D�t�d��vk�A�&(I�"`!U(�uR�!�3��-��$�#T��D�?��M�QR�L�捕Wgдb�.D�~�˷���|ΓW
^����?as�]P�����$a�%�������'J�0S�O~u����Q�k�D���7C���˯!���n?)r�@e~ʟ�Ĉ_B��);���x��`&�h;D������K؟�s�x���aI�){��q.9D�����0amT�����6~0��r�|���Ov�On�D�|����?��N��ك��
%Ⴑ1� W��`�nZ��L�Iqy��'��)�s�,��3�֌_��̋�R8)�����"O���Fǣ{B*�����'N�y��s8� �#����.��ʙ/?�yP�,D��j�a�	^�n5j&jɦ_�D�j*D��RQΙ/�	�����X�>�"�'D����c��`��R�
� _N���&D�x�HPvY||�v��>zL�Y�8D���"KW%,>NY��Ʉ��Uk6�#D�P��ܯE[P��>�<[R�3D�<z���%�������*�YS�1D�,2d�L;g>�[N̈,0D�l����*CR��ҷ�XecR�:"*D��� ����lha�W�~!+`�'��/e$���AE%p���?����&��Q|*�j��W�By �eS8�h�3�#��D�~�թ� ,D% � EWک�wo��c��ac\��X�4$��p뮸����Xh�a[�M��ic����AV�+���+�Li9��+*���@R�N�i�j�Kۉ\�'a M��N�z�(��@�ӒG�0�3	�'R|�Ff�(*`Ypjÿ9i�T��'�t�ŭזa< ��B���'b���Ս[��Y�G��mJ&M2�'q�@�׀ѹ �Ab+�!0f�{�'T\�ե�	o�R��0���X�l-��';���a'M�"@�0���.J�`��'�Ҭp��TL�}�⇆7=��
�'�z����@D��u�R�8�*��'����q�/K<>�j��2(���S�'�U�#��C� ��+��/�^ً
�'Y�x�����n��y��E p���Z�'|���� U��6�F�3�T�����  �ˆ��>T6dP �E}��9R�"Ot�xdg��z���	F�57T���"O�psaG�i����%˨l9Fv"O�U�6iʻ;�yX6c������"O��SW��|���'�X�oI����"O�(�&F�c��]x�@V���1�"O���(`��8�.
�2]$ �b"O���E3�� b��5��젥"O��H��_)��yg��\�$�"OX�hf��iUp�7GՃ(Y�y�"OLّȓ4���ht��,@He{�"O:@���n���ye%��}�j�A"O��)��ϼpZ\ȳ5���@Pr�"OpM�V��(cp��`v��$�8H��"Op�!G¿(T��k�	�nz.I��"O&|�橖?5.Z𻠏	5^n芣"O� Ύ0`W��J�3a��j�"Oʠ�s�͈#3�l�笜)_
J��D"O��`Ȝp��U� p�0�"O���$��i�f�'�ȁ9
���"O*-�aiK�N�h`F��LH���"OlA1��"x�m�E��2Jtx"O8��2	J{�Y����
0R�"OM��k��w>�0c/�Q� ĳ�"O^��>:��@!/�G�N��"OZ�Y7đ�s+�<P���8��a�"O��!g�4I"ٸ¸j�"O�tж�1T}�3�,�o���"O&�����@�R�`�ͅ�A�f�
�"O�-
g�,g���W.ڬ�Q"O�m
&���T���Hť�w�5"Oh$��m�W���2�dݫsW`\kd"O��BW%mX:u"�>���%"O h��ذP&���c`�2q�2��$"O�H��
�2>�S��5F2$`�"O�4��^�Ĳ��U8#����"OZ(��H����	�+�@!�v"Ob��Q;vB4��)۠$ـ"Ob��gҺ!R���Gӥ�d���"O�yjƧQ2������ k�f[�"O.�ك�Ǯg���D�خM�T5Jt"O��f`s~�bW�ȣ:��e��"O�h�Iy�b8�&+�#4�^�C�"O� ��-�(���h���4�`"O$1�I5rgP��`G-���XF"O س�&�UFP�ٗF9/��=�v"O�U�ׄ�=#hh�HKМwet�r�"Ol9zc�	5Y�)rL�[�X�"O��¢m�w
�c&�-�N�v"O��ŕ�a�F��/)��ap"O8����]�q�H(�Q.C�1�^�˅"O�e�E�؎baH&n@('�v�Ӡ"O����LB�&�Iq@c̓gv
ha�"O�B��/� �:bC�8jc����"O��*��K<5����%�פYv1�Q"O���G� ����('.� \^hѻ�"O(��PN�*"��)hrB�"M���"Ol���4mb0�]1G�5i "O8��u.��GY����K6d�4"Oj�� *[!��Ȳ�T�f/�쓱"O��8�*��O�b�`����~����"O��	gA�]a*(;�K;�: Rv"O0��#
I0S��pK��EGT""O��ČGet�{��.H�94"O� ����*�D�0�%[�q:P"OF��,�o���ax�*L��"O2��i	L�ʭy���0xJ��"O��ᔤɘp�Ku���@dj
�"Or�x�b���ʩ1bNҨYN�!�"Or���@Oؠ����s�<`"O�m�`�I�Eg���kM�+�֜Ñ"Oΰ��,_0���x��3}=2"O2���HO�{��!��I�t{�D8"O�p�T
�.s�Yy�y�Z���"OZ��h�̐��Q%2���"O����F�)�X9��&ܬ���'��L�fo�u��9�U�6`x ��'�I�5/��t偵M�*G:QA
�'��)�D&28�Fh��p�&Y[�'iJE�d�R@�l����4�V-�
�'!80�%�{�����@�%3A�M�'Ut���&N�l9bd����[	�'7n�0�i�(t<Dz��=?��@K	�'�
�K!!�#]&��Z���T�	�'��A"�F��(:eE݇o`���'�|4�0ᙁ/�
�aD�B
5h�X�
�'�rP�6˘^ƶ���ۦ1v����'+�1����đ#�G܃,���	�'��i�C$�Җ|JbO��5-�p1	�'��lr�쏍	�I1�(�*P{�'�(\C`�+2�& �E��T�d@c�'e��{5�T�k*"�����K�$��'Z���"�`�aA�_�z[��?D��ꠊ�8�-��c�HeZ#�>D��0D��&L���h$��g�d� ��8D�D�r"�T�\d���N<J|��2D���C�_Ǫ �'�
�5����1D��H�� �_�⤘&
ɶZ��ӣ=D��'�Y�.��%3Wm�%kܡkR/(D����!�$�M��'�
hC�Y�@�'D� ����W� ث��[�0cze�T!D���@V�QTb�;��\�n>p%K�G=D�8�l��Vʲx� V9P��rh;D��ɓ��?BH��VJҐ��٨�$.D�0���G?m,)�S�5X�9qW�6D�̲�Pa�V�����'ph�#��1D�j�j��t���	ϝg���×�.D�8�4HQ�Ke���w)N���=�?D��ۢ��sd�L�i7��ɢ$C8D���b�Y
|����0�R�~��#%8D�H�o�bc�!:�N�=�FQ��*D�d�7��0���#�K�W0}��3D���"B�!��Ѱ�L6���UA/D���W�]*.o�ac�K�a���f.D��1�(#����"O󞨋�a>D����ٞ�(̘B#U�|�dt ��8D�0b'�\��!�@��"�Lxҗ!7D����
�|!��<:��R�C5D�� �E�}״�k�`B:p�<rE� D������6"4�����0cV) D����F�ۤl��B �bj*?D������.g����䁏c�0�F�:D���W4@*2"E	S�f�X��"5D�p�s��%���:ׯҶ!:y /D�X�	ϡP��Aq�n�4$ɣ&	'D�����Ҕ3rဣ��,R����"D�ĳ!�62m�v��,Q�^�%� D�(�Pj�A[���p��		^Ƚ��S�? �x��Z�-dV�N�n�+g"O(�@�hQ�s��!�U�X=@0 ��"O@dBVdJ�UD|p
'�F��i�W"O̅b�%q�x�9 �ԫ*+X�r�"O"�aD��T%��ӥ��(_�I�"O�Uabʀ'�Z\P1�եv��""O�񒅊B�q2��W(S�/���7"Oȩ� �>7ٌID��b9<8Y"O"���nB�V�"���+$��"OtPFg\�8�BU���S�my\y�"OZ}�q� 0��ʳ*��se^�&"OX�z dY�
��!�S
�d����"O�M��@	)@�����A+5����"O�	cLϵ4M<���H����"O`X�F�I���STi��>m�"Oj�:��R
p�>�PQ��7T�@��"O<�8C��O���hW�^<F����"O|XÑꕀ	�ҥH@�:
\u�S"O~���`n"y��\H�lQ�V"O�1#�AI,��C��4� �"O����+�3���z ��f+\*'"Oj�#5m��w�,�ԃQt9�d�@"O�h��/k�<H*�c��/�bt��"Ox������P��
�\gzX�"O������/Lt�1���8Y����"OP��<'��]q��Ь+>tQ�"OEaE�G�q ��bRA��gE��"O��8�˟�id�0Rw&�}��! "Oʬ*�N�={�¥���G!��q "O�]2���$n>,�p��5n�BQC"O�4��'P�gul�{�MI1� � �"O>pphс�����a9��u"O�p�Q8dcb�*�mU ��"OH􂁀�*Za^�헁|��{�"O��y䑅Z n�8Å��Ʉ%��"O�x"�:K�����8]榔�1"O�<��瑄N�4�
�E���"OP�WI�KrlH���*�:
3"O (��%kb	aw�][��c"O��Jt
�v��9j�`ЈC��S�"OZ�HbL�~�L�j���4�P��A"Ov�y��ձt@\��"��2m�d�ZF"O�)�a���n��A�DN��J@��"O�0f��/H�aP�L͟X��"O�p2�$��d�C�-��a ��
�"O��J֩[=m��XՌ
k�2){�"OF��v�ο����C��BQ(�"Oj�XW�X�w`f̸7�]q�P���"O���m��r�4}O E��"Op)����<���pf��}�*I�"O��&IK�lvV\�Q�ɪx�D�hA"O�!H����(�s"��:[&r$s0"OF�����B�0\�%�]1sP�b�"O {�A��P�e떦!,ʰp`�"O�����	��t�t��=��D�"O�Mx5��.xq�$)N�SS"OF@a�Ȇ V���֭.lpQ��ޑ.W���6���p�֘5��'�Ф�7�M�b*3�F�+�xz�'n@-q�lJ�8"J�cE��&�2$�	�'s�X`�
0ah�P¥��Q!n���'�B�Z@%
�n�*�Jf\��3�'� $�ڪ4�t���I�}J
�'���3�zڰ	��V>LJ S�'����f�#�ܴZQ��VA�AY��� �����q�������"O����_5"�ܤ�怊�k����P"O�H�%T�/�� ��%]3#2�
&"O
�a�+�"=�!·���p"O*���a�l⍈s���3�X8�E"O�8[v-� ?н�N��#%؅p"O��q6!����H���h`�S2"O�����6E`��#Z�\��qɁ"O��i�a�*F�aڷ₱{E��:V"O�M��I���	�V�� ^:(�"O>${q��x�r��DJ�6��%��"OL5QQ��6X%��W<cW��*OtPD'�31��+��D	�'���d�SI�� r��C<8'.̓	�'�z�y�͎0l��1;^��'"J� ���)~$�32&Q�B�')R��'s�Th�@�Yqe��'�|� $D�*������"�и[	�'v����� ��T(�j�.@��'�(� �;,g$s��`��ѻ�'4ԣeE-e%.�f����'�.��7gH���g��>?��a�'���[U)���	-у�n�A�'��	��ֹLOBI���X�Рh�'����R�Q Bܳ!	s��`Z�'��y[R��9�� �ͷh�E�'l��+�|o��`ǌ:7�b���'��<�Ui �@Pн +ê/��H�'Pr�r�n9v���&fV�?!��'[�*&�
��Б3c�!����	�'�ڨ8���}X�A�d¬ QX���''
 �fǓ6QR�y#�Ι.���X�'���{�H�wpp�rE'i���'��Q�3��L	�M�]�6��J�'�������13�*z���e���'�!�,%KF�1S G�0��	�'�dP��fR��e�>w�h���'`�aq���h��kR� :��	�'G�L��M�#b���!f�͎���']���!E���ഈ1I_|��
�'���Z�*_�`��q��8}���'�ڈ���`�򱣱G�)p�XL�	�'��$F��X��F�%d�,(��'�2�[�T4�P)(�ǒض���'��`�eoF0@�x��ƫ���&�
�'l�|�T�n�@��j��	�{
�'�¹d�՛"��h��̇k����'�\�J:/mΔ)�	P��~�R�'HrE1��S@��3�iZ�qȘ���'��<�e��@}��ꢄ��;�(��'�`$�N9<U��4R���'�������o�ND�Fn�=���'�:YM��V9��h6 ��}L�Z�',�ɀ��'5�5�f��rp�h��'�!į�;�E��M�S��8��'�8�dĔ&�����;GT��'[�X��ն-?dH��"F}��j
�'����1BI$~�v����1z�l�k
�'2Tę�d^-P=8�D�.j��=j�'�����#}�H���[�c+���'����ۮT�n��f�	 c��r�'�qDLD�<jD�W�I,fX��
�'�ڤ�g� I�
-��-I��
�'�1�Jܲ'�eۡjX�r	��8��� �I�F�0<^`8�̎,�p	q"O����9n3�\9d�Tk�8���"O���2��۶�Z�gY��n��C"OR2R �+
���ϫkL�]��"O�q+�d�"'1�#��̭q�@U��"O�Yؕ�O>�V�c�E3�8�Z�"OȨ���=�P�ȃފ*+zd��"OP���xv�!!�Ԩ��ȷ"O*��w��2Q�X�D�&Ռ��P"O0@K� N#w��JAB,Hl	s"O�����^:|s\R�� ��B�+%"O��S��
}�JaQc��r���i�"O�ԙ���?J�Ȑ����Q�\]3�"O6�(%ߥw�iad�ۂj..ݐa"O:�a,Lg��ӱˌ-B�U�A"O����ᙇ����;�>ɠ"O�RQ�G/GJd�7	N	Kx�"d"O�3���2k̈��d(�@c���"O�Bo%&��t���{��DZU"O��)��$b�(��������"OH�QWI�mXtaEC:���06"O�y�'ֵ➡z1K�D�A�"O�t��+_G܆ī�c�nD��"O6 �*[#b��(�C��R�h��"O�����-��혡BZ�d"<pB"O~���n���ұ#�#6@r�*e"O��@h_�0�}�W��΄�a"OraPNQ@#wBVaD�b�"O�3�SҸPO�9`�C�"O��pU.�@�T�
��6I�$�%"O�<)�
I�m����`d�A�"O��I�n�V{IC$c��gÌlPŗx�@�)O�z���"�r��Y�_�H,���$�0?�C8����U#)(��ڡ��Q�*xдn���x�"�31����o�K�f<�Р���HO�4K���X`J��3�?�������=*��}ID �%y2C�Iy.`�+�)l܌Q��#qi7mХA�v�3���Jyx�S��M����)���6��>�Z�1�.�<H�"�,�Y�#\� ��qy����?!F�B�u��T����Q���W,��LCS�^J/X�]&q�a|�Ԃ(l2�9�#6
1U�p@��X�@�Kad�h��p��A�L��"f�S|�c�`�e���!O���'@6��N�V'��	���<
��'>���/�*s����̈́�D�����6D�ĂƁ b�l<��(��3����eC�	"��֓b(8W@٠yX6�}�����5�ـ��MB��ے�l���{�����̞.z��Q�'F������aJO�蠃#�`�bE�u�Oٺۋ��F�P��q����_�8��� xQa{�c1~��'ڭB!Hwc�i�\���jY/W�fX�S���4�F��2�'���� ���M±�ʅc�ր�}r鈃u��8�OC�T�D9�2זk��z���� V	L$MQ�S�!�ч���8�ǃ�5��j�F־	��-�@� �<�[W��6�d��'�r�Oa�$�s 2�x��O�W��4�gEL�!�䜙�-�D*�6tm����^�Θ�Q�͂$B�ieKǆ;��`���n�>a�B�?�Y��**`T�)Z4�K��� B-�����b�J۟	ܢ|�R�C�FF�l�d�����%ڧh5aB��P�`�x7��#�ة⡄���'�<��5�V+^!D���f '}�F]'>m��anj�B�$E=�<� /D���g"4���F>`0��e�N?Ѥ�Ũ\�� Ʉ��O?�	�hi�����H8�@�[U�x��B�	)NE�� $�ѩx�q�p���|&���O<0���RuyLq'>c�|�w�>"2�]�����9~*x�#�9�O�	{�Ν��X�	�=�Ĩ���Ug��)cd�i(<5C��@f	{�D=�d�˔��S�'�D�`n��pJ�>ݱ�A?/F�X�J�} �@N=D�� �Ip�ngP����l����#�O�q9��͜�1O�>yp�L#�l�6��_I�]Cs-9D��{��ڧ)(D�u��6��@��9��-�H����oٮI+c������R�g:!��M��tѣ��5ٌ���D�*!�dׂ4r�і ݘG�N���Ob"!�۟E��}P�K5B.�`��F/N!��O�8v����➿�(�#��\�!�d'j�-�T�-&��1Ƭ�52�!�Ăi�e���`��A�eɻ�!�2��-�p�P9D�(Q�ˌ�ZZ!�!d�%y� �4�0Y�5A��LF!�$_=X���"f��;I���MKL�!�d�OD�85�C6O�ұ�m�I�!���YL�	�4�"7Ȯx",�!�����fo�1M9�d��R�!�d��H� Q���ĦZ�|C��p�!��+A�D� @�"�ʝ���m�!�ٚ���x�	V�|�vd�p���K�!��FN�(��W�o@��΋�{�!�Γ=r����Z�Vj&��5C�7!��ň!��ΟLv8q��N%~o!�$V�(�������gN�۶�՚7 !��A)/>Ń�������>*�!�T�D�$+��I�y��`��f�B�!�P�x��b��~��#/f}c�"O���gI���0-];g1� "OT�+�ß����R`ւ��&"O��#CM�
��DE���A��"O���C��/��<j�dX�H9�L2�"O*dqؘW����E�T)&~m*�"O�g�W��$��?��qi!"O~��ƋJ�,��[!�c�Xb�"O�m�����=!���;��je"O�5 �N+���	��Tl?j�"OR�*���+�q�f�ڨc"�Zf"O�BGo��x-�$��!��q!"O�Q������e����!�lR�"O����M[S�����	;'��d"O���cnS zf�S��ߟt/qa�"O���ė"�������СK�"O|�R6�ޔW/�q �LK�t��"OL��R�p��x�'�� �Ɯ�v"OF b��Π�t�(��b�`�)�"Olx:EDl��ESUj�D���"O|@�@�S:"�GL�?�Pj�"O���$	J��|c��G�n���"O@I
�5���x���tN���"O�1i���S�0a[W$'�у�"O�ApŅ�T��8��ش<p�"O��9��6��ԑ��.]7��k�"O���s ϙ.*���d޶\G����"OHi[%�[6x��Q�d�q@ZՃ�"O�RMB�!�(KJ*B��q�"O x�t�11�R�,��7l�Ak'"O�:C���:�ƐR���2C�ʐj0"O�1�4m��o&�<���M,q@"O����c�'�.M�k��Jk*�"O*#��ԆN�b�k҇
�U�.;�"O���'M��[�F��C���ћ�"O u2�i�+���#V�+�1��$̅Θ���)m���ytk��>��'�U+ hN��)&
�q;��;�'�t�q%ޘF|��U���V��'Kt�Hd� ,u�X@��+L`^{��� ��PBG�$r�<+5 �=�ZH"$"OP�"�F]�m�uLX�&���c�"O�1���͡3�����U��x��"O4�37�KB�]{N�j	��{�"O���� �	��3���|����`"O��c���>�<��	L�{Ռ�J@"OF��w�
V5�ųIv`�]�"O���
�	��<�$)X"W��"O��h"�E�E_�3D��":J�)�"O��Ǟ�j��Ta� ,!���"O��XR�!���J��ɪe�0�t"Oh���(��f�P��U� R��#"O(���I�X&]{g�Ǥ0���{"O��rO*g���{7��0���U"Ov���3mJ�
B�4R9�P[ "O�5ٴ��~I8M�a'@�H� w"OfiZdL�UJ��e%ÃY��H"�"Ov�Ƃ^-�PI[�={��E�"O,Ӫ�Jn5s��K��A��"O��YoT�@<�
����8A�9G"OP1���P汊�A��`�ِ"O6���Ōh�J��t
�&u5j�I�"O��+bn^9�qr��#�9�4"O*��˹o* t�'�s�+"O�]��� $1rd:@&ظg�FiC�"O�T�D*P�B��#EN5�fPa�"O� �ei��(0Px����
����"O6�`�R�V�rH§b��/j�X��"O.�G�4_�ʍ��Svh��'�fy2$A1f�"]��H�&�<l�'����͐g�Թ2���":�	�'��0� �&B6�`��F���'�(-��͍��Z��J�BXf ��'М鲤d%qZ�*�"�D<>���'B�= ���N�A5�V0BfiH�'䤉J�J�-6�
�j��8��0��'�RBI�C���҅h�.{P�X�'����r�дp�#ĸY�'�B��ĄY/wJ)�W
�*��ԩ�';B��&^�?D�����$�I��'"��[2�.x��d�*>^�H�'Y�0`c�� g�b�YQ%ր9��E��']� ��/�����3p��p�'Oĸ�$b�$u��P��7z֌89�'�l����zbf��$�(y��=�'�pх	v��!��[c�@p�'�A�iHDטQf7Q�R,�'Զ���˫p���Qb�Y'>,�C�'vPx�&@�:ry���-d�(�'z�0v���z����
�OFU��'��a�kl\�iC�b��
��%R	�'| ̈`��6��R��xCD]ir"O�5���3_��I!��d3p]�S"Op���`�
b8�˅�
0k/�h�4"O��!'CZ����p���g(4�"O�5���U�X����蝠J�`�"O�2�PU5`�F�$����"O�E��D�$��]R�t>P"O|�&E֩�V5�P%K�U�@ b"OT�:����D<QV�Ҭ)H�%
"O>1����k��r�M�C����"O�ɋG�_��� cl\X.�e�$"O^����:'�|}rE�c"O䄫��
=<�u�ꋳ^�<���"O� �-@�GۺRh�y�6��mB��u"O�xjF���6$���	�Y��"O�}���`�uX���,�zYC"O:���L\�}�2;��@�	�`�+�"O�L��V�B�(���#����S"O^����C�`%h��~��d�5"Op�A��. G�ȋѫ�
�\A�"Oz`	�o޼n� S�d��u����"O��qCNΔ/e~����+;D� "ORq���d'xu����P>���"Ov�K�-��I��2���7*�S4"O2y+��Ϟ_
�峠�ܙ+ˏ��y����N��ԣ��
G|�QZ��2�yr�L2w�2�܍:��I��Η��ybMǐ	�rd�VE@�+�"Aل����yr��
Ob��R��� 9���o���y��I����O������e�%�y�c-5X�0i� ��	pb�1�y�H�sDta��(����4ʂ�!�y����}�� @%������y"dӠ�r��dn��[�y+v���y�@�^L�9�4��
X&0�s�A6�y�f�*Ҝ$ "�RL&��ꛍ�y���� 1��6x1�a�À���y2e�(�p\�p����4�p�'���yLP#_���G�C�
�Ȕ���4�y��Pf�V��e�4*dx�����y2�H)��DJ���+؂ezAH��y�ō�~�2�d)S)�t�A����yBMЧ0:z�	P�0(��S��$�yb��E�aR�[,�|�Seɹ�yR��xh�!�nČ+�*�s�L��yb�ʯA&08Ä�+X�N��1�ҝ�y���x��9$%�=D'� �`�ӷ�y2�KNR������¦ 1S	��y� ɧuDJh�ԉ��$��'Ȋ��yҢ|�i�QL�'&1�檅"�y��A���%{uF4s�^�	'/���y2MX-Z�@@��FN̈́�av�˸�y�͘�RG@M�'J��L�țPF;�yۂT���+K�z��в'��6�yB˅
d�c4�Ү`�(����y���f���j�7*� �����y���Bw`l�SII�P�is�*���yR��,���6
W� qP���y�_�.6ԱB�;H)�!p�Ǥ�y¯@�|Z�\X&�E�T��1��,�y�ANGzL$mH�I����5��y��V*[���jյ>H�@���y� ��Zv��1�e�'K���ГKU)�y��4Ȕ�A�bش?���'ؤ�y,]��&=0!�?Ӕ�3�i��yKԣZp����4��W����'�ўb>�Q����@fb �V���R��;D��r%�=|G�1��^./F�1'o8D�p��@�q�3�J2�j�ɃL9D��BfOׁ��}�N]:;5X�a� 8D�̳�.G]&�Rp䀧O��y�"2D���^�j�
eBÉ�#&pm��5T�ԛ��πIQ�Pj��N4;��V"Ob����S��<C�� CJ��%"Of�0�S�h���7�ǉT�j�["O��ڔ$$%�q�5J�"a�P:�"O�y@c��T��5���	*0��IW"O� \��ӅT(�s�#�����J&"O�LC��R��P��`�� ?�FM�A"O�P��`H!OIq��Yu���"O$��A��<*8t�̏�!����"O�]��E�R=BD��ˍ�w�\ "O�qA��k@�)ӴŖ,ʆ)��"O�	HS�H/ؒv�^��2a07"O QӅ��X�z�pD��<���"�"Oj:�@B�"��g�Gj��#Q"O(!s������i���6�"��#"O6�#�oӂq�(H�1�֯�؍�"O�)6�\�8tU@�(�.5��a"O��	3jK�*����Qt��p&"O�i��̊�#�8���@��)�А��'|p ���Uʤ;@$�ug���'>HQH
.ì!��!NYM����'�^�X�Ό e����H�N���'<f�B(0�BĚ&FG_�x9�'�<��c+¶�4��hȶ9��d�
�'@�9@�!��-Z��#"� ��	�'�̩��س>Sƕ��� �4��'�Ӡ��-6d��5�߲��y�'t���+�Rpբ�W��$��'��)�$ĕ+]���4�HQ&�]p�'
 q� ��Kj4�6�<�&�h�'���&]2�n��'Ȁ!.N�ti�'�:������8�l�@$�]5�B��	�'��� !Q�+AB4��&�,좡��'K���N�L8I:��ڱƑ��'[^U�&�Y54��d�r ˛��u#�'O��b(*T%�ݒpNɚ*�6�	�'��Hs��E	��!�FSN
l)�'�P���e��9���KS�8!����'���Z�k�2Wx�|Q'I��z�`��'����MR�H���֣\����'���`0��50���%mY�F�n4�'a`�#c+�!F�1�OE+��Ĺ�'G��XK�n�Ԙ�(�`\���'�b|�2{��i�*��l���'],Dc�ML(R�H��ᔴ� hR�'���b%[*B�v��0���]�2<X	�'���G.A�1�4h ��#��@	�'�|������j��\�f�E|���'��
fśo{���wB��!D�<�cK@~��`'��:�*�3� UC�<Qt����Q�����t[$&�T�<y���.[}��X�%)y�*5K��JM�<1�Y�>3�aE� �=��$��AD�<ɧ�M�u#N�;7� $���B�M�B�<Јζ���2G�>�HKq��D�<��Ølkȹ�-�(pz��ԇ�{�<y@��(V���K`�5I�I�b+Tx�<�2@5#iJ�9[rz-@�n�7Y�C��&K^���+�1]�@E2rȏb4�B䉥C�P;�j�N�*)���{�B��!2i�m!rj*8�*��Ϫtx�B�	-,�"MP���
��ʶ.�!��B�'>4���i� � ҰϞ7پB��?�����
JXȳ��ΠB�\��*��U2r��]3�C��/;$C�	jR����mؼ];�B0�DC��	�8�ٵ�%KY��r$��")VB�,8��k��G�@r0�C�T=g"�C�	>:L�Sț3T���#+ǒB�)� �XR�hCOW@P!���y�Xc"OZD�&�7r���#Ҥ�3zH@�$"O���4�c
.��p%��;���1"O.%�t�^:0)�t"!���~�0Xa"O����H�nĖQ��ʧ�)�yBl̛P���et7���EF�yrd�!i��)V�Ζf�:�����yB��%�e�$W-��c0�yB��k�J����J��YV���y2�%JqȆk�H��զ�y��[�6�0�a��F��a��yrȡ_&T0�C�+B�j����5�y"o�)A\Zآ���=t�L1Q
��y�)[�D���0��a)���0J���y�V f-9�d��[�V���nڮ�yRo6oL@)R���8�I�ǈ�ye�d-Z�0�g�&|���e�:�yBF�-z��$J��I _Ǥ�ٴe�y"��ZPnx�!eńP9����A6�y��^�j���Ѱ���RU*�Z�c]4�y�"=�l@��T�M2X�����y�$Inm��#��d$����y���b�
wI�<�Z�j���y"�M"H�D ҆�/ᲄcf�݁�yF�5B|d(j���{��a1����yb䆳�@�AbS�^��(����y��@O�=�"��Z{Z(�@@��y��Mz�.��Ń�<s��jv����y��ߩCw,�8PL~� �0�H'�yҤ�3�$&'�����1~���hoNpC�T�BA�,���h��O�<��G�# |�W�*g�9�)A�<��	��':p��]�}ʎ�%C|�<a�"\�HN�kA�2�Z%*
�u�<a%gB�_*�����4�=�A�g�<I�$ͱE}�� 1N�Ȝ�-�d�<@���nÜb�ȫQX���H�^�<�dh�&)<�1��=}��!q��f�<�)[!�S&��85�q�b��f�<!Q���Ko8��RF���hd��Wl�<I5�R�R��c�	�9�5ٰ�Ui�<�jN=X���0g?B�id/Bb�<A�Ǟ�F� ��Gې�L%8�J
`�<ժ̺ �tk�Mڗ�����B^�<A�%D�v%$P��JW�qGv�붫W�<���>�����@�$�Jg�H�<����(��p� �>�|RU�A�<���n��ȹ��&���P�C�{�<��	O�B��Q��N����!w�<y�G��4w.!��K��fp�8�)�s�<1VlP ��J�
�,y���9#�s�<�B�*F�(l`���'PZ�Mi�Wp�<�t`�|�f�1ЋP"mr���0Ec�<�#	�;4|M��gSyPz}H��F�<�f�V�_ �"F�5���اτL�<��* .�=i3�Ż1���prJ]�<�L�5v����#��8  t��Pc�<i1�*@�N{�-K!B��1���G�<i�B)�x�7�Լ ,BpB�P@�<�ՂC�Zdk��6�40�4�b�<YCf_�#-�Y R�̈G�ht�*�B�<Q�jG0ViB�����$y��A�<�A�Z$ȺDK���,���G��<�[#1��Cu�вaj^YJC�T�<� lh#�K�)j8�b�ΈRy�1��"O�Dۦ/�D�P0�,�
�~d�"Ol�� �|k\���L�2z��s"O*X8U��.6L�� o�pŐ�"O���Q X�4�U[�Ŋ�rôI�a"OF���N�8����̞���"O�I:�Ō��ȓ�
�%u�j�#�!"D��������b :�x!�"D�x�`S<_}n!�&E�/8J)�Q�!D�XY����p��8�r�ֿEn�s2i>D�؁��>��A���4�-��#8D� ��DF��6�(� �Hd�7D��#�J}��@�'k��~T�4�4D��5O�� ��%l�Y0}y�a1D�8����laR`+Ԟt���0D�T����5~�t��Ԛ^8P�".D�<i���w$|y�*��L֙ ��*D�H
p��|��a�s+�)v����f+D�ԑ3�*f�����/�:d��m+�o*D��2�'�u+4��RK�Nð��C*D����=|��Qc�Ψ=�<���)D�|���U��Ԭ�(A>u?�A���2D��3�_�D�l�+^=dȩȐ�.D�<��E��Y���{'�*�I�ac*D�\����ip�]�V�����&=D����$x��c!fH�B��7D��S`��>s=����2hb8�	�F*D� c l[;]��8��Oѕn�&Y`�K;D�Pȳf �D����x���7D�TqᐨQ�f�hŀyפ1:�5D�l[��/*��I�&=���1�i%D��A*��|�ѓD�Ӂ\�z��%(D�\2���^�� ��]�2�H'D���C�;oÔZ���2�@uE$&D� ��Q�K}*=����H�.%x��!D�`c���*�Tb٧j�IHS,��y*�1�Ы�폗	�YH��$�ybGB(-�����$�����a�U�y"�8�cT��y[r1��7�y��H�i�l�
�oCր��N�-�yb�S�/��hQ�4_�<hѷ�ԭ�y"Ɍ�]��8Z���_�X @A���y�/�&IjM�� V_����W,Ц�yB! �A���	$�ˎ�4|)R���y���Y����g�N���S���y�,��Z���K�G_�K�E���y�f=%UD5�SM��LRQ����y��W�*d��I�K��CV��0�yR@֏b��t�3�ܧ:��pS$�U��y"��?Q� ��D$r��F��y��t(Љ���>8�F��y2�^޸uy1˳0`��E�֊�yB*�1���+1^90�La*(%�y�&����e�S3>U
Y�d���y��#h�9i2MS�6-�ڔ%K�y2�=1z�9����<Uy��6�y�G$� Ƞs��-JhR|i�gQ��y)��wn�J4�zi���I^"�y��i��BF�dyl������y���&��ٓQ�0Z~�t��O�#�y2FZc��$2'ÅL��dk �M��y� ߲d��u�U�+:x�8����y�Ʌ
��h"WB��&(F�IC�y��L�
{���䎻�x��2��y
� ���e��ULpKW�E���lC"Ov��&NE��*����<!�TE�P"O��
�fۑGWɎ5Xv|��"O�%�0�W���=���۵���"O�D{dL݊!����Ia�Ԍ�"O�1Sc�P�C58��K�a�8��U"O�i��-�5_���+3+��tˀY��"O8=�M��x�b`	��i�x�a"O�<��ˌ�]RPDf�H��D)sW"Ol�u��ky"00��!=�"O���U�(b�`80�!&����"O�$o]�"� :e��Xx�]@6"O�(�Q(��:���t�Цgj�ܺ�"OH�Z�H�Tg@E�a�HVP�R�"O�1�m>�@2r�V�P�"O���C�<zJ�	#�D� S�*w"OD5qD
�]��Q� �.1DHc"O�Ud�Ug��	8[#�Y�"On�XB��(}!x�H���,I�Nq�g"OHx�f>{�
����B7;'�"�"O�,�@���E�p*Z�4��C�"O�8�u����x{d �w��!"O0����	s?60s@ ��P���"O^1��ᚩ4�Lc�V/��ɺ$"Oz��L"�����-ç]�N$P"O:;2��j�`�ۆ'WE�`xPV"O�m*u�:-1�8����um`� "O@T[E�+~-��L�@VD�"O�L�#W4	N��I5̒�L%�e9�"OP.J�}Ee˭q�\�$"O�M�4�@*3��%ސ7c�Y"OPy�T��6U irw��_��ȸ"OK¬�4�!�@ 6
[���Ć��y�G��`~6���ݞ�@� «���y��J� ���0tOH#� ��l �y� ����M�(^pQ˽�y2덚oÄA�cQ�(|�ؐ�<�y�C�a\%R�LK0ȕ��I��y�F\^�a�5E:J��Hz#�y���7��11��4�nY�b�y�ʁ�#rq����+�&=J�����ybC�1����E�7-.ԛv���ybb�u�D�¢l�/1 y;v��yZ�����ԗ7ڌ4��(���B�I�b0����_rrxze Ԣ&��C�I5��3�O��d�t42��ŋy0�B�	���طLߏ���J�E�<+�B�I�D��9ǫ��{D&�����V�HB�I:D���1�+#M�h�4� tX�B�ɱ�ڸ�d��5��0(t&��6�zC�	�5SJ<x��L\��WO^�P�.C�Iߢ�B�H�Hؘ��kنb��B�I8��	�ƶ�b�j��(b��C�	�C�z�@�W�>b��0B�m��C�I�]*RLCG$ʡ(����*��� B�ɏ�-� e��@���#��"�B�Ɉg��}!�HR&�1Q��(H��C�I 7���v(�Nb9x�IĿ-S�C�ɢ\:��b�U:?e�9S A��C��?8����[�-�&�� +�� .�C�I^ji8c䀋k*�#�H�itC�ɮM�R ��pc��IPlR	3�ZC�	�b1֝���`g�H��23� B�Ɉ_ �����Ρt�({0�I �C�)� �U�#�8=IN��D��#Rt��'"O��B��kOl��vLA�R��4Q�"O����o�	pޤ��b+	��pɱ"O.����D,c�j<�$��5xl���"O,�;rƅuK<A2�����P���	ڟx����6��O�gzƄ��L?r���Ě�,����rhL�����ן|P��BxZ�L
t����B���	N%Fx�S b�`��sd�8Ƒ��Hu�����/M+rTbyQ��	ź3���B��ɳ%�Q7]e��:��ӣQ���A����5�"�'��6��ON�N��5(�T*j�a!��R�
�t�'_�O�	)ғq���3m������
%��	�M���ir��A��Fc��T%ȇ,��c`���~2��0/F.6��O���|ʒ�T�?���M���2X�b𠛗R�f9��/�+}�jȪ�A\)`v��g/�>G�>=s�liܧ�
]c;�=�1z "\p�+O�7|Z�(�4g�a[%	 ;'�A����.�h�+ܢP���|��Q�B��3�L46�ʈ��(��Xn�rr��$٦MZ�4�?y���i!R�sW�đ'6�:Ě ���J�'��',�ƌU?S#f<h��0bn�|1����(O��o�M�I>����u�I�7M��`�Ê-WƪeS`i���:/� *v䞉�?a��?!��n��.�~���G�:� ;���Y.�:�+Ԭ_�@
��Űe��&)�Lu�-36E�ni����a:|U�q��(2\�#�oY,8��ӥC[8��"�<t��I+�[?���
	�<O�5��>���Z�@�
U��Z�x��I�O��D�E�	۟,�	Y}��F^�`�k�L	~ P8t�Ҽ�~��'u��k�M�Z2���D�B�|�rV�JƦ%��U�	�?��	Xy�Yܵ3U�;jo���e��$te��!%!OSaR�'&R�'r�2�'Ur�'dpp��!\�`Q�`je	���]�B��Z��3�N*#���c�ѕm�E~J #V��`"�5:�(|y�F}3l�G�{���ʰH�G�������ՙ hZb�8t&��IEz
�Jei�� h�GS�D�h`� ��M����d�O��ʧ�i��� �D���1-�(3ht�O �=��ЯД0 �bTZ��aBa?ig�iJ7m�<Q�Ɖ>��E��*Ozl%*^�^��1c�n�9��2Tئ�?i���?�윰u�h�&*�
d��JbH���\3�U��B�&qh�@�n�s��I7w�]Y��k�D9�$Є��a��u�&�Y��_0�|<b�-(���?e_����͟��ܴ�?Y���K��!hB��B�:rU���$�����?!��?������w� QC�*�VDt��ڨ!��	A
����i�*7����ԡ�`J�xF|�!�	�{����
p��x3B�O��Ħ|�,��?���M۠��x\���o���,a�w����B�]�ڸ8�=M�`ax3gM�/���Ic�)��a�do@���_gHJ���isӔ|��j �S�jA
�E�M���ʡl��zsD��P���56jz.���4,~o I��+�M�R��TY�4z`��'g?7�J�8&t� 6#�/ ��È_. ��O���Oh��?i,�l�8,���]Lrv�#œ;"X�Gzr�i�7��O$�l�՟T�O��5�_�\�b�)�F2 �V$��>�!lOFȱ��  ��	�'�jw&�;h>���
Y l�X�'a�M3�Iscԅ�&�Ĺ�
�'l��悍?���`��t��);	�'�b���ŢU��K�
;t����'>̭���7v(�B�F�x8���� D�C�՞>؎\"�B��$���['"O��"D�6L��� ��*Mʠ��$"O���P�����b��_�ڡ�A"O������0Z�	K�E��I� "O��,���1�??Fz�#"O�@��nF�T��T�@l�㬽��"O���R�M�B-hƭO�����"O~- '�#A�~l�"M��?&���"O�� +��3��@��[��Ÿ�'�t�PCn�1'��;�I�2V���'ܔ)�͗�)�F-S���<YF�h�'��bA�4XKvA_:Xv����'�.�LO6Y�$�Vc�8J�8��'��X�mɉ�}�����LQC&C�I8�d�+�� �TEy��ǜo?�B�əY.E���D�3+B�$d��6��B�Ʉ_d3�Ĕ�D�R�U*l4�B�I=$��0�&HI��9
�	�>�dC�	A����B�8^?�ո �$o�DC�	�M����dl\\jP�0�f��y�h�,� �A��Q�"-G�4�y� �
؈$i�D�
O�����7�y���+�D�h���^/�M�s���y��߁xQ�鱇*P6[8����)H��y� � PyD��!\*<���D�yR�¤n���S`"�=�� ��
O�yBHR)H[°r�Ț�5i��A3��,�yr�4D�l�#B**2Xɓe
��yLF\tA�1���zjxГN��y2�S�*�x�*6(�8lDIᢄ���y�͑��
��ƫչLu�d�� ��yR�қ/o�M�ե�;@hIs� 
�yb�^�Lz���!�L:D������y��sQ��4IN�`��ҡ����yB�=
�D�8�gS(eb0�t��3�y��ʡ���C���$%ҹb����yBT�S��]��'�3�phB���yr�'�r��eUI��@#��-�y��ԣ]�N<���:.~ET�ھ�yRj�"[l��チۃ@�:H��HD��y&�=v�^���,2A��ra��y��U;(|u���M-�Ȍpc�Ґ�yBD޶*L�$@3f)�f������y2cB�2\0��!�S�P�J���y��,Q���Cʸ�$a:3�J��y�*F6�|M3Vʍ=[MJ�K���y�-�wc�a�j��r$�2�u��jb6��E�$��eG4�.mE{��'e�<�EA��b��"�.D������'��������<|��Ɠ�K� 3
�'͠T�g J$#���8���F��ِ�'v��K��uH���@�˭;�^|(�'r~0�!�Is�\�0ē1�䔚�'ƴu F��0SCE˗JŻ;����'�L���d�&e_� ����/߂a�'4��"�柼<U"u+���j����'b�!��ȏ ����#:�L��'v�DA_�C*�� ��^�7��
�'(nsVB_�3PNtc2H^� !��'��)*��۔+`F�c!hz1lX�	�'�@=R���lD	Q��E����'n��4�Z�y�R�c��R�Iu�Tr�'~����4�����˼,�\���'�ʴ��kF$x���2#b�9vIZ��� ����2(~�}3�E�%F}�Q"Op͒4fV|
��z%�O-Nu��"O@��T��[jDMѥoSO��(`C"O�b��0I��m�����b#"O�T��'I�����=�Rq�V"OΑ��F;O F�lǘ:���w"O��؃IĤ}J\@�X6ry���"OBqc��A�#C�끊L�,��9"�"Ob5y��w�j9����O�d	XT"OzBB�̜����3�Ƞn�ԵH�"Of����n�AƩ��k��E��"O�!�a��)�B!BFW�n�.T0�"O��h�,Z7v����V�*��yE"O.D��Ϝ1V�b����9y�j9XW"O��Z�@qS|��R2A� ���"O��J��t#�#��ԅ.�j�@'"O�F��L������3�f��d"O���b-�X2h�"j�$|�X�J�"O.����yY�݀�		U�r�R�"O\4��P�V���P3*I*F���@�"O( 2'����j�O΄Jä�Ȳ"O.�I��Ӷzܜct���K�0Y[E"O���ܲD#l��B����`�q"O6=��I8RxC�+ʹ�`	2"O�����͜̡ 'k(d�|t� "O8�;� XE
�a���\(���"O�h�!�O#Uy�pbŗ}�(�e"O$D�kQ/sT"�"
+� �R�"O�U�e���Fo�����!�"O���P�7�`��E�}��@y�"O���ukA� �>zP�ƦTR"O���?PJޝ1��NM�y��"O�tB�� 
a��d�U�I(�R�"O`�{S���12��3aX� �8"Oh��F*l�.��D#a��a"O�hk�&IY�D��/�/Y���"O��i�-
�c��@� _�t�r"O
�$%@�J�d���P�(�ޤ�$"O�Hr�S�Ah�X�c�:����"OL@�B��Gr1�r�D$�<1��"O���S��^����GO]$`����!"O�%�pe1��0�X�u����'��,1�рO$��+��E�:zT���'��=���˯q�4e�th@,
pdh�'�>q����`E�����$�9�'�L@�Аt\ĉ��͜	E�d��'�^�D���r�|#0�֒v*��'� �X�oX�9���<YL���'�e@�#�5� z��S�3�*x�'�t!�E�-?��x�`��%S�Ё�'�Z�
�jW���H��"ـX0�'��P�)8����F��d���'"D�GiT���Z�+HJ���'��U�h��'�fx9%�����'�\��H��0����̘�2k>���'�$\R���.�f�+���.?X(�	�'�Z,"`��?Ш���D�M�($��'h�e"!CU����r�[�K�Uk�'�T%�i�-1��K�K�P�Z0y
�'b:�@�-��"Ud�W�Id�y	�'�2 `�'�x; �ޟLA�'�,�g������7���z�/6D��b��P#�,X�D�:i*��2D��I3h]�upt2�BK$i#���+D�� <�2���!%P`�%�@;q[�m��"OV|�в2ǢYB�B%l��"O�$�#ШJ�v��BX�i��Y1b"O�h"�
��'��y5�I���!�c"Od\���0�L��D"�C� �J�"O V�#tR�`�b�C��x"�gLj�<a`Ş�\�b�	�1]�1
"ʝf�<ө�	&��d@�g��h�V�kł�L�<9��_9/ (Q��׼*$D���D~�<ّ�U�lϤ5����5u�jt�6Oo�<9gJO==��8y�-������R�<�7�
�#@���� Z�<�a �%. @�fnՉ(�ȝ	�N[M�<ဢ��@)Ze�e�Ӌ{Zl,��Qq�<�,S��IZ�`�/q�A�J�i�<	�� �&P�R��ۄ	�F� ���]�<ц�*Y� i�6<��T�G�[�<I�ݾ'�ݒ׈��%�r�`�T�<A'��yF`鴪��lŶ �g�[�<�g�'Q΍��A����"�Z�<a�	���ji:�lL�B"����BR�<��,�kZd�FNH�5�[GI�<q�h�
f}K'�7.����ƊB�<�]�C�� 0�kݱh9f]څ'YF�<)�x?<,k"�P�5��Q�!�}�<�2�H�'��)��Z1x�����_�<�cEċTBQ�lR-fu5�@�_\�<y���?f�N��ɚ�;
�!��T�<�gH	�4�^8;���"=+�X)V��R�<�P@G5;c�I�E
�%~���Qb��h�<���N� �� �Ŋ!h�,1�o�<a���?����%�G�a'�Hp Sm�<�ÅFG�,�#��D�CnTՊ�,�f�<y���B����eL@�JH����G�<�E sx<��5A�	4����D�O�<!�/,-$���
�#H<=��lGW�<	P�O%8�9Ο�#��R"M�Q�<���0ftq32,�?>�I#�JN�<��b�uׄ(pV��@��U��j�H�<1e/�_gp�E�hi�#�E�<��#�������^��ഈ�}�<a1��Q����{+d����M{�<I6�ȤW�\�x��O5���c�s�<�s
��v��1���2*Ѱ��I�<��b��K��:���+	a���"
[E�<��j�+:�Ma�.βW~줚�g�<��KܤE?<y0V�L�_��T
GIZ�<�&F���5-^=��8�L�A�<)o
�q���eOe)"P�N�k�C�	Hc(��"�#2q�p�ңr��C�I�Hz!SF���@�u�7�P�GۢC�	����5�� d�)��B�4E�iS���M�ָ3!�0��B�ɘq>��M$Q��;��[�u�lB�ɪ@�����aHQ�U1aO�k�.B��%FyP�F��`�v�Sv�L�>��C�I:lKpU� $]3+J���-׳-u�C�I	V!�1�*��l�(��3��n��C�	�Mdq���2{����b���B�I�]18��7`^9�d��Ə}��C�ɀ#�,��J�vo� ��L��7h�C�Ɏ4^�@�WJ̝X�fL�c_!nC�I=��0�q�E9iTi��۠@A�B�I�`[F%����o'��*p�B�)� ,Qs��$[�X[0E�(h�Yi"O��rˊ1�{^͸Q���¼�ȓYZ��/�� ǲ�0vNA?�J��ȓi��H��'g�& ��ٻ�D�ȓA����яĘt �U�Uc�:Z$����:T�а��޾?Ղ+���6W��TZ���C!PS4iR�^�����ȓVad Ⳮ�	%���5�˾Cc���ȓz�F��`��
\�oǠงȓ!���0k׷b������݁eB��ȓ�d@է�VĜ���λN�Pq�ȓ)5�s��*j�Tېƚ:jD�t��C�IA�0zf��rU�L�rZ�|�ȓXy��!�;B2j��S%�?Tie��&RTQ�fKn��Qg�7O_}��%�>�C(Z(�XuL�
v{ZX�ȓK�|� ��1n�0�iC�LV��ȓz�;���pϖ��D�a�ȓ?��y�s�"q>"�yv�KZ,9��@т=!�@�������q็ȓZ?�!�uǀJ��X��&^p3�ȓ5�}�� a�Ń�Ij0��MR6��%ČSlH�� j��i��|Y@,Eft-�aQ6�>}�ȓmɤ���c�'��=�q<�<�ȓ�9[�(�+� 2�	1
d����83慈E��7B�m�d�22�����5ΰ� ��A�P#
O7� ���$��<Z�Wk�b�@0�Y�6k�܄�F�P�
~:�I##�(Yq���ȓm����f��m�Ht��ƌ�@�2������g�ַ!p���ǥP�:�(-��BRj��$\�7��9�MY�LK,��v�d�SwmH�s0Ґ�v��aR$��N�"�a'm��7-Z`�A��?DzB�ɤTy��I���->��y�lA�/n�B�I�nK���G��:U�La���]<C�	�{N���K�?#(<)�萧w9�B�ɑ9 X���Ǝ0��a���Bj�B�	�d�F�@�o�l��%`b��B�I�a:r�c�k�+��-(P,�f8�B䉼=�����x#���fԶW��B�	7L`�M���W+T�xᨳ+�j��B�ɹ`��$�U�ۓH�)6!G+f�ZB䉽g2lY���"�"Q��㊈3�HB�I#L�hP�#��2�ElH:T�NB�$mERI��-	j2�����Ĺ<�LB�ɗ�~��`(Z���0N�6��`�'�L��G
��t���u��tX�'ހP��H�[����@��h�lm�'���wÉQ�i��?_���[�'-Ly����n�|0��@��5
	�'e�5�R0P�T��"�25�2��'�l
�_<#���n91��l��'���&�
<F��V+=�8,{�' �|*t���S��-s��� fƴ���'�N��6��l�a�&m�3t�jl�
�'}<)T��;a��{�Z�Z�pI��'�,��m���V���e�j�'`�x�  �$��a���
[�.��'�Vu���I�b�H�BQ�_	Z*a��'<���t�Z�A��2!
����'�(�cثp�"xPcS��Ԑ��'�v4#C+禙ز�AK�A��� Bm��@�=��ةV�P�Z�����"O&�"���a�|<�@ͷA����"ONA��NH>�y$c�p3F��f"O��'��!�B�����wD�z#"O� �@U,
>�33�O���0"O��j���H�ް�a`F(y���"O�����@�p�*	���>��т"O��ۇH58t��@3w����"O�+%�п4o���2O�0�\�Z�"ON�zwG��w����-�.H�쨋�"O6	���
k��5���Z$QB��"ON�#��	2K׌ ���L��|���"Ou���B'{ƪ �M<3��R"Oz�K��
l��a�G�K�"O�����]�^�)��#'��q"O��q�͛�Px#PG��Y]"�G"O,�Q�N�'je���.1��g"O��8�p:��ڲLt�チϸs!���@E��e�?-JB�f'o�!�$��k�!8ݩd��Z�\�!�D�-XO,5r���Y0�y�@�l�!򤞹k25���Х`ݐm9��"B�!��4+�8h�&^�*�0f���!�J(H����Ą�G��M!F9U�!�dW�i��,�7mB�Z➽��-�9�!�D��h���E�N�8Φ���ݙ#�!�$��"��9���'V�ʴ�޹v�!�d�%>�r�P5cB�J8���u!���~�8�6¬r���� �� e!�d�q#��� �B�W3rh�7�>M!�Ϗ��P�!�'6mf`U tK!��F�j���uC�����	5S,!�(,V2q��_
>���_!򤌸)��ݪ���]^�p���a�!�䎚:����\P\�vlb�!��/Dh$�mߗCx��Ta�4�!�K4��-xp�L�0(�|qQ��)e�!�ӆ��PD�߽�{W��	H�!�D�3'L�́��ɝ
K��De�!��ոMXdmi  � 0���@�L �j�!���zݔ��#�ʻB�xX5,��7_!�$_ |Ʈ]��J�;�N� ɍ�!�Dt������z��!'m�3�!�䂆G� �������#�%�9X�!�$w���Qnͤ�6���%�&�!��dp�1��!�&x��F8,�!�$�c�.��V݀v���&��V5!�W�e�.1H`h�	���Є̃I !�$ޗKR�`�J��w�N�K'!�l!򤜷5��ꤋ� �j%���C�D"!��@K�@p��VL�A���I�,!�$Ҫ�f��
�g?j�h�7�!��C˼����B�m����\�E�!��� pV��x3k��"U��^.$�!�Ĝ�V�)5o�\E:�C�Ѻ�!�$Q)��5{A#y2��
�S5!�$=] �	��-K!�	���!�Or����	�I��%B�`#|�!�ă�k*:L�"J�`�x��`�c�!�$V�r͢���)^"�Bm��Y��!�Dʔ���x4I�SR�\���ēy�!�d��9�q��Ą�t2�-���U�P�!�D�,6��Ұ흽6u�2Ύ�h�!�ET�T+@�� �*�LN u!�� �(��F� r�`�\��-��"O��!�@��$���Yؚa86"O>8�b�6D0� /���@p"O��9�(�m��8���M�!����"O�m���ӻs,�5�5�y��3�	���+%��<u�)�&�$���)pDj� @�7qO ��9Jb4�և�X�.���4u` �O�t���1Yf�K4�	wY�����ĦpR�Y4B�8��Hɡ��@*$��_:�9q��/uf���)�M��-���I2%����O�nZ�(�O�P��+J 5N|hPBj����E�a	�O����V�{}��hj@���d��ۤ��p>�w�i��6�f�8૱	� 9��ѫWb�4N�$�a�
�M�fV�p��	qy�O��4�x����D��d�#�9t�7L=�¬/{=,<���)z��ڂ#ܨ��O��;-�`�����9��� ۓw]P�lZ�FM�5h��=A��ncC\��I�<"k�t�|��sj��S�׮r>Yk�J�d>�o:}h����ٴ�?����il� AwJ�%����-�.���'tBT�t��	<rL�Wb��DSD�3=�#=9�4Hq�֟|�U?���I��I�eA��N:H�Q�������'{04�lZJX��@��ƂLy����-սs�����b�&����$P��A����/��H�'L1#<�Æԯ-�8�e���t�Rt�!�ܷL�Q���I(e��E*5N=)����O!�fO�d��'B>�q�3�a�&��kâq"��OJY�0��O4dlڰ'N��<�����d-+�T0�� ���HQTBѴQ�Q�P���6@��m���xiv��,uq�M�t�i�7 �����X�����$�����Q��G3��1���ox���	��P�ȱ�ٷ)ab���oMƨۗݙ+�`X�h�2n�
Š'�� J瑟@����+T�V�Ru�5+�"���a��2����LX��c�'�+��h�ūN�)'`�h��Iڦ���E�E%��5��j�jy��oӪO����O�O���h�(��k��h��آ={"	��OF��d�9^^�X��/�1T�\X���y9���	��M���?�C�i�BL�q%l�z�d�<��89_f8�a�]|��MҖ�oRT�l�ɷ Gy�1�ђI�tBG�ܯC�x��A4��a�צ`��B�AF?���i��	�C��A��]*~z܅�c��7O��;XjV���̇]��DR��?%��@��cJ�OrHi`�'-��nӐ���~B1�ֆj��h�eJ�O̬TZCN:���4�"=)1$-,%n�r��93f\�v+	z8�d�شM��i��2,ߨ[F�u/��(\���'aLĚ�jy�N�D�<�O �']�aJ&LQ>��,R H���L�.Р�ru���es|PJrCϹD`KY3�q����w����t�I!0�MV�;� ���4z�6���(9�hI:`aW=cOl��6�	:'���|��5�Bp��J�澔ˁ킒��`mZ	�����O }��r��i�ZU�eIܛv�0-���ĀME@�'�b�'��P�z��N�XLX�H����~�Q�ߴJ(���|2�OD�N"<�ik�OR;;�A��!��9�$�&����	K� ��   ?   Ĵ���	��Z�:ti�-���3��H��R�
O�ظ2�x�I[#��y�4g�Բ �I�n-s�E�_�]	p7m�䦕��4E�� ��q�	x8�Ļ��My�֠�B��H(�Qy��7U�#<Q�
~ӨP(&m�r��xp@DB4F��r5X�T�$�����1?�E���/��7�f}2*,�1��l�?)��0��0L־�iP��uy�`�OvԚ6F� ��9O��@qJ��0~
�rt�
[bZ���(��L�@���'�,��$�ȄyQ#��!Ӹ'=�TΓ�|�YՌQ�����fn��hJ�$�<�ቭ!�'���#1���{�L:�I�h$�'�Ex��|�'�!�f�N	^PH�$$��}��-��&#<���>��I˟R��X�H>C���w�Y�D���O(��{��]�Jr؉[�B��K1�=S�,�MSV�1���"<���	��pˀ�8���(��[�HI�>q�	)?n��B�9Bw��2b^�H�����<�fȕ'5��Fx"��N��|� �%�L��t��'	��F'|�1 �?�@�"<	(�O�e(����.��L8��Ev�����$Z��O�D�O<q�	�W�؜1�O�"
�j$�wL]?y�3(o&�O����*�1	�D���N`!GK5F���l~.��>(��4w��	�/^5� �O�h�q�סe�8��F.[e�0�X����M b�\c�0�'�ǁG�'�b�S�������$�C�2��ۨO�����d[3�OL���LR&����f��0��:F"OL�y��  �~�s��A�X�"Oz���P
��)�#�;(_�P�"O2��*Z��z�1!�.Q�H@"O����Ic����B	5�jS�>D���/����+-d=�@=<O^"<����.(y��-�9��Q�G�u�<�eA�<�p��範�1ZX{A	�z�<��a֋���3��(�d�J�b�<���ȃ ��q�bC�*(����o�g�<�5�fe6I�3�P"#�Qe�a�<)��ɶ,D\
�g��bA$_R�<1b ^<�~xqP�؃o\x�2'D�d�<����,�p�J�	_4���A`�<i��Vp��8�5%7NN��U�^�<�p�%i��wIBYɒ�QT �]�<qա�T�)rU��?�t���h�A�<Y`�Y�.��|�@YH:�%1�JX�<�b���h�f�;A��D	��8�EH�<�I� +2�yC�''Zbu�J     �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   �	  �  -  �  '  %/  i5  �;  B  IH  �N  �T  '[  ma  �g  �m  3t  uz  �   `� u�	����Zv)C�'ll\�0"Kz+⟈mZ�p|�57���DB���H1�ѯ&q�5��7�$�b�ی>��+�FRH XY�f��%e$���;F�FiB�'>Հ,y�'mx�a snQ�)�8=s���(-��(:0Lݧ||<Z���I<���@�'�A����4���蟺�d	�
`
�c땘,�z���0�	Z�DΐzRf��	��<��@*��ߴ+��9���?1��?a�n�>Pc�(�[\>�j��¢;����?�
�;���q*O��ğ*K�����O\�ě�a�n�AU��8C�"��%S��v�D�O��'�b,	!���C�?ٚ'9�t-K1Nz�Q�m0\�����ؗ/��2OP�Z'i��P�2���UI֥��Q��̓��'�P�2�#L�	?� �[$��)��}���/� ��O\��O���O���O�˧�y��ېj@�@SS��/m:�A�c��?���i�R6MSȟ�n�˟X�ڴpr��md�lo�Lce'������3�U1�X���J۾�HO���k6�'x S�����0�&/���v��o��@ؖ˞�x`���ڴfۛ�{��I���CwM�
P0����W�k��f`H ̂ �fyK�4c$z���� '�YP���,S�h7�5��aP�d��4l���M�V�N�0�rw�<8��1��!z]�}`pA��G^~��u�i��6��צZ���A:���v%�	Xh���M-�4�@�D����G�#`���pKJ�H����ώ�M#&�i�>6-^�q%��φD����fo��XJУӂYO\(�g�A&H"qo�����1ʉ/m���d�c5�m9U�ٟ��?�C�. �R��$�¾eu�`a'ǁ*Su���$�
����n�8�m�?���� W$�2�8�	0|�8xC#Z|���K'�5�ؽ��t2:9��(٫A�#f
�T�ȓ&�� 눓��#!�ӣMB$B剄�t��+�Xy�p@ѯ
sVB�	���'��Cf��yүY�3:B�	 
�,"
(�J0q
2"h�=Y�g]T�O�d��q�KiP����\�"2�R�'��jT"J"{Ȯ!rP�X2�X���'��:�� �ĥ�WH���
i��']�0+qo� Ub�@�7�������'ق����[z�+B	Z�wA.l�
�'5<%���hS�I���8l'4��#R��Gx��)W&��4@�T�9�%H�K�{�C��05��e%�� �\�%Iרz48B�I�c(@�ȋ~��Pi�㔣p� B��o�^��f���b�+��b��C��,9ej�j��+_%"BR�1p�C�3Z�ֈ9��0m��:�H3M��˓/=J̇��-O�����)e-ь�)"C�%��I0�F�%��̙cm��C�Il��ӷ��2���	v� *o,*B��������Q���h�fѴZB�%"�ޘ�R.#�bro͏�����9H8�n�۟\�	�)p�E���9�nek$�V�T��I������V��`�I��Lj���ƟP�'��N�zΠ� '�
1Ϝ�2�F7�ax2!Z�ː��X�CQp���~�pgN�P��rF	V3{ f����;8s<��O:�o���ء�+��s�$\�Sp��U`Sy2�i�R��)�=,�J�h������L19&JE����'MP�Q�m5��a���D�O���B R5$��"�&V�J�ã�'��I�L��u��ӟ�'��'K�$F�L*���]3�*M1Q�z0�	+.�A���;�l��9���p���M��)�@��.�)§m�ȵ��.�
J���U��j�I�'�����?K~j���h^�Q>6%(%	�9@�bI�K����?�	ӓ*�\Ĺ�Hϵ6�N�Q U-��D�9ڧHՎ��wȾ�p�C��>f�	����?��g�'P��F!�����B���<Y�'�(+�&k�|�ǃ�^KؔC�'&��@��Y�D����DK��MLM��'�T2@��9�V�kW�����@�'�,d21-�3< I��#~�r�'H\��H__t�R7қG��ܛ4�Ĳ�yB�'aH%Bg/��q�6����T/���A���x˚�Cw ����!o�`�2q���Mp�m��'p(���(c��Ш��~�q� �?�@�'��AB�'�(Dô�D<��0��'@�s&�1
W�49�A�7˔�N>�U�i	�'1���<�I�;q�6�c.�d��y��@R���\������	6$ $j�ݳ^� �)�-��f�,�� �I(�산 4^l��)W'.*���*0�"�flr��o�����?w`�*��-�FYJ�f�'M��, �����O:�u�'V2��XY�@%�JH"qO?��M���%���O���D�ilĺp�
>e�����۳�xR��O�u"���Y�.D�G�<ɼ�A�'��I6fך0�ڴ�?�����2��R,)�7�����(��kρ1��'#�Dh�:�p�%B�k��T>��O��̓�*K�.Q3T�ߍZ�����O��3�.��ڴy��A�@���}�El��aqЕz�b	NPx���M~�.Œ�?	��h�@�Ĝ�i����r��!��"J,B�	6b1,��4�ȡ	_����!r��?I���1D��`�@V�bc�z�j�-ZC�$l�ڟ��'Y6��pa�����Ox��<Ycl �����e��|y�"݌�F��"	�;�"QX5��&D q�*�>�I�o�	�$L@@h������9���E*H�2�a@sc,�6p�)��>�u���q�O�L�v��p��
�T�(L�bR�'{66��O�����O~b>˓�?�EG�*D�40fe�:d"�ec����8ړ�O̸)"o� p��x��3���{В�$oZ͟��I��M��������)��#�T@ce6ţs
7\�X=�4�	Ŧ���� �Ioyb^>�ϧ�^���%B�?i��c�,(]�0��A(�5������R�쁪V�����O���t�iY7��"B��<��D�W���D�RN��#���;R'l�6N��Ipޣ<��ݍY�
��b�("y�h;��O�UL9�I��	�4�?I,O��D�<A̟$�AU�͗��Rr��;qM�K!�|R�'� 2��̍1�4!���&{Z�����'��6M�O�b>���>){0�	/�(X�g���5'@��cb]�P�C�	�u��%f׎Xp���e���C�I-���ac�Yr�8����B�Y�&l�p��j��:0E�[R�B�I8
�Xy��U�;�z��'.�"�nB��;g�<T�ʹ�~a�f
�<�,�=I!U�O:Ԍ�P.��z�O��n���''�9��ҚE��@�EP�X���
�'��ty���	OS���f���M�
�'T�e@���G��!K�����4�
�'~D,J(/L�V+#a/\TX
�'v�H@`��`PE��?R�^�{�{��Dx��)�.���c'C�b�YҰ�ƓSTjC��%N�VH�3Μ�-�*�#�MD��.C�I�x|��`�U���E��>]�B�I�$n��ӷ�ˈe����`� >$B䉜3p�l�'+�%.�ΰj�@�� B�Ɏ,<�'�jh�őp�P&F>�o�T\��I&<�~��"�ŷ���%+�F�hB�*D}Иd���} �!�'jȖi�,B��v�ي��Y�X>~qK��E(�0C�ɲ��X��N�&n@ kH<,,C��
U�N�p��c�,������$�d
�$�6���`�K�(���*R�Ūe!򄇉v@ة�	M�o��I�V�M�{�!�����ʴ�[�ER�P�%[�ZB!�)pL}z5AQ�.�k�e�%!��RT/˗'����%_1E,!�� ;��K��C��Պ�$8�ў�P�/1�'i�PR3�����B��Vd����N��h#�c��M�le�q��\A��h�42�ԯ?�����jР�ȓu�Z�?PvN����479��@��x��8h!j��&`<QOẍ́�t���D��`����'*H�	 ^վ#<E���N��9�S@W�t�bEkuᕯ**!��+V�p�o�6�P�
ӡ��M	!��ؚ/j,�8 ��Z��XQ�V��Py�&�S�\@ё'��X�JiFؾ�ybI��S>)X�O�6I&��y�ə�]�����+�\UP݋������o��|"葬�"U��ŷ�eҤ����y
� ����,�nM��ʟ�v~h �"Oܝ�눢��£��t_:
�"O� ���4h,jO�DZ4|S"O�Cg�4�V�����cS�p2��'����'��AR��
�~Yj�a�L����'�4kr��q�Z�;�l�6Z�5@	�'���1I�'H�`�6m�T���B�'X$�$l�b�Y�#�Jr��#�'NF�ph~m��5+X]~�X
�'�`��엣G�}�ŅM=���ʉ��؉~gQ?=Hb,�d�J��"�A&d�,|xB)#D�ԣ+Y�rBi��!=3���@��!D�� u�V��@��2�da�W;D���W�6x۾���O�a��0+5D�xA5�ǄU���Bb���t��2D�܃�n�gl���ȑ�vU�0D��O���a�)����B�Ɓt��ѳ ��V��	�'=r�1�n�Вqy[v��#�F�<T�� H"�sw�H�mg�$�qO�A�<� �ep�T� 	Ѵ"�ZQ����{�<I5eН=�*���K�3���AK�z�<ٶ��
d�xh"e����"��OyR�W+�p>���WC�����^�l��z
d�<�!m�;Z~舡�Q�\,�"�^�<�v�0vo���f&[V΄�,O�<ɵ�;'�	)�
ƊV��h2S	�N�<��
�吠c� ��>d�B�Bx��Q筺����^�b��Ȓ�)^� ��!D�tr����O*4H	���m�Iæ� D�D�fl|_�Yk��� ��XR� =D��Q��4Pn���I��r�`ມ�/D��Ӫ֡@f���8�Z(���?D�L C�j��-�`gD=m0��k;��>mG��Y
�T��q[5Mj�zGHߖ�y��H4p�N�~<��c���y�@�O�n}2�B�,q��M�W�G�y��$"� �5"ޚ{U�1�B�(�yRĝ�6x��;U�G�x�>�@S	D��y�m\�}�B���_w���i�%ΐ�?! ��c��������Ŭi:6�� �Z�+�U��;D�\ÃF\G��<HD�9�؜�5�:D��B��^�r����KW*m@n�H"�7D�Ęu-Я����
Z/+�`A�g�4D���Ԯ o���i7�W�'�B��)4D�x���ۍnp��.
��"e�v�<9ƍE8���u��+
� 9k1�
*f�H��dg,D��6-�'Dv�4C΃�)"��C�.D�lZ�J 0�Q��_6F�L�PD-D���d�+N>d��蒱V�ȸ�N+D��@VgW�}]��9tH�\�l��F-)�O�3��OX	ad�8`�>�k�d��?����"O�j��.��!��c�/<r��"O��Q��4Bk��J�f�B�"O:����Σn��,�'I� �<%�r"O�,"�i��s"b!a@A�Rh�"O#p��A�r��r�2.^�xT�8<��~�$+T;J. ���)�~3܀���e�<��.қC�� ˳&����/�b�<����3���:��+G���[�$Rc�<�Ђ�2r,���4��le�W�<	T���&��6�W ]Ö��|�<Rl���P@�ϋ�@�P����@��*�S�Oʪl��oٜ$� ɜ�X[�4��"O�x��!�����)uX�SW����"O� ,I�d���Hsjȉt��8�"O�����ȇo�8�Qa��#6�ɑ"Oxh�e΅�a���	􊕙`��5"O8�X�"L-�����e��=��X����(�O"A��ÃN�0y�T�S�~l}��"O����U�;\A%�F<m��4Q�"O�9�`A�z���ǩG�D��"O�$Ȕ��K�RHh��z~D��"O�Y�ԫHW�|xU��΀�a��'1~��'�i��6^w�H8&�ֶ)��i!�'	�p#�E22V>�8�k'�����'��QG��O����ⅉ-��h)�' �<�nI�	a:YR`A6!X�j�'�N�1��r��ԯ����
�'�lL�t�B�k�^��ceF�"�҉��X�d�Q?�
rO�(�Q���α'����D$D��PB�&hL�zG�A9�>�2P� D�l�a���%��ISID@�B��?D� Jգ�9L�-i��)Ya�b8D���M��]���In��3��4D�L��%�>��z0O����O@��)�x^���^��X��荃�^U"�'�l��O�IYڐ{T�+Qެ�
�'Be��$��l�xȁ���?:�ܵ8	�'������N�BM<�X
�/���	�'����bN����h��H	<�}��'�y���ՂW�$ŘdD�6`|,H/O�$i��'���窎�"��k'��%,�}X�'?lt�B�'[G>�KbjT'�`��'c��)DNO�{N6AB���	�-��'�A	�˂�8�l��E���}!T�p�'�ܬ�W΃'�I����p ���������HE��
5�@�K�1h��ȓ��})��ѫ �B�h��L-q�����h��iծ"�X����E��y�ȓkߪ���#aB�Y�.^K�t��_�Y��D/[��H5��3;�E��DA���`H��Y��#-(�&�D{�쎯Ш��0B��M���X{���	�ňa"O��Ru��"�n�����,�>t�1"O��(��6=�(��Î���h�g"O\�w-ӱ-��{�b�"u���{�"O�͸u�2NhjUX��T�5��%�A"O�Y�%� V&"5K��߄$���'�'��������>��J��Z(,x(�S�f�4���ȓ=A���p�ʩN��T#�D	�i�ȓL쎁�2#�3.<�����YG���ȓ7�͋���ҨQ�NZ?588܅ȓ	i8�hg�S�&r�8A3��/b�D�ȓ��U��*X�#�X��#��S�`�'�p�
�>���+�뉂/������X5zd}��J>d�tϜ�S��H��R�U��4}h��`���0����Gʘv��T��rnd����U �p�q��0옅ȓn�����&��k:���eI#ȭ����r�6�ɲ(��Ɉ!��|�f ��R\���מX�̼��@�)=`�;��L�G@!���
��ٲê7�hPdeX�B7!�$�fJd���$8�:�i�c/f�!�_��E��j&;�aF�L�!�DK(I����̅�+>�BЁS�:ў+�%>�'W
��#B�B4 2�h#�ʆ?r�̈́ȓyun�* N^�)���rw"�ԄȓZmb���")��h�6!������S�? ��o�-6�%Z�͔+�X��"O$���F.©�FK�7&ۊmY$"O �aS��G�႖�{Ǝ�t�'��p���S�q��)t�O�a̜�y��Z��z���P����
 8(�y���ͩ���ȓ#ҒR!Ҟ1��i�@�nS�t��q) 5�ል�*��D���E��H�ȓ+�D4���'�8��Rk�-d�v���g�����3�T1HR���V��'1`�
�8�r����@e�bICS��"k��Q�ȓ��Aq6E�q`pQ��[.����i/�Y� �<l���R�י
|�ȓ;-2���'�k����Hx������j������4a[N�a��QAx�h�&��XqW*�G��m+b�ԡP����Ў=D�Ԉ7˄!09x�Ȥe�*|J�31�:D�$����	���C �A}*X1�e9D�$���/;|�Qү�k��d���2D�<*�{��a�9M� ;��5D��AnǴ����Gf�3a�2�4��yD��+����7��E��)I�y�k��P����tcʚ)ZlA*�.$�y�h
8�� �A/|ک�&E��yDY<l؂�kς!��t�&N��yҫ�}2��j�f-/2<�c�=�yѐj�(8a�S�Թ�J�?Qb������R!�Z�)�����"4�|r:D�أ��W3I���26	ɓ�|���4D���!Zd���,��>d>@ �3D� � J(�4�P�*�8o  �6L;D�ph!mu�6@� ��th<���/Mp���)L��C��yR�����O� �Ϩ����O��`��ԮF����ʊ5+l@ັ��<����?�cujFm\�;�qKG�n�y��O�2�I'F��mI�IBL*��@���}Ԁ�1Z/�ik�ꀐ��$����j"8z��0X|�!���R�&Gy�R��?����On �1����o1h�8��\pz �,O���d��d��") y4Tmr1Q�2q�}��<1�B�.Ǣ��D��5�D�[��\y/� #��'j�I{���'k�BͲK�U< ��	� PV�-��.(�XP��J��K��x�j�}���!^�
`��D�Cd�X����<a�)N9"�4 G�Ƽ	52Ё�E9h���c"8�JH�!�<W0օ��(��dF�I���$�O��S�V~�gO)"�� ��p��y0�`�>�y"R'5
� ���kji`����hO��F���э�tz�+�+ִ���ܱ_��'�R�+�����'���'5��O^��Y�H*-h�L 0W���$�Яs=\��G�}�J�&��j�Z���
+���D�4+G���`*�׺u��E	������A-;�ΥH M�@X��#�?%�Ɨ�ysh�6��I�i �qP�av�8�R��'������?����r��:���-d�$H�7KH���FL2D��	�鋊H���+Iغ�#�O@UGz�O�Q�|�ՈY�k���wa�u�\$WD��mY�;3	J�踤����H���?1�IΟLΧE6�\`S �8&��,��"�:���ĦG�k�PR1,�+D�I��4H�"?9��O�"�2���:��\j��`!a6)�h�N=j�A>���� 	f�ʽEx��_��?�%%Eq�P�0ð1*Z��� �?���:�hx��k�v@���>E�ȓCOHA��+N����c��U��'�7��O�ʓd�Չ��h��1�����&��(u#��� �i��	�?IńO�?����?Æ,`#$��@➆=����|����?`ܝ�d��Py�SPE�~�'gŹ�3$�L8�#�iK":y�钮�Ow�d��k����pQD��O���(��1]��㲨�/��D�c*ɪ!�˓�0?a�	�~{:��5D����elSx�<�*O��1ŋ
J���t��7B
^����4J���,����� !V.��9��`��P1�Ix%�-D���%V�E�d0H�ڕ�ne��$)D��9�JB�J�4Mrb հuI��<D�� >�xf�:���1%o��rl�M�"ORYR�»B}���-& ���"O�萱(�*Bt��#��r�����Q��O<�}����Bs,C��3ӡ�6�(ąȓp=���.��8�a�1
Ե}�Y�� ��!�ł�:XRL�īƭ;��0�ȓJo2(2�������$�#g����ȓ^���5��;_UB$`A�V���s����GQl���D�r���Ƀ3>p����&L����ō�:`����Ɣ26!�$�����c� +l� �c��?%!�Ď�*�M�D@[3����C뚈R!��?5)~P觌�K��%J3
�n!�D��'B��J&�p18 r�[џ�����M�I>"��=�|�[7`�{�p����X[~b�'�"�'R���aؕM���!I�����j#�����J5�=4�<؀�sz>�X��I�fƚ1��0i��x HK:.��M�ڀ�a��ŋ�Ѝ
��˃A�x��2�I-���d�O���Oh�S5���;�T�۾	a�A�r�P�D�Oh˓���	>?q���L��"� ���,3 ��c��|l���d�u싮Qo�E�f�[7�ʴb"�꟨�4�?Y���?�.O&�d�OX�5L�Չ�iMt�r(��)�(@���'+Q��F{� G
W����e�5d�V����D'��'���K<�g-�O:�'	���qE��i=��2�OW���d�'�z�	"�ӧ�9O�@����$I
Y�'p����t Pb��Op�,�&��OV,$?�H�E�<U�܈��ꅣ:v���5M���Ɋ�~��s�L��M�M�V�K�a(�`ABM�rn&�'t�';:q�J���>�B�`��!�8df_�mt�,�?Q�@�x���U��?9pK�$wҁB�M�bxr�q4gV��r�"}b�3}R*����ə�Mcs��#\�b|)t�Y��`���ĝcyR��9���ȟ�PA�v���f��* �����z?a5(I�T>�I4�����֟���'B�|��i`�:eo؍� �\{�u�޼�'���D�T
�B�B��GL	{O�1�p"��?9�L�����!?��y2��~��?J�(�a"D\��䙈Gヹ�?��m �O���f�J�pt �Ie)ʿ�Tcw"O� G��9_�Y;�A�31�x��xRP�0$��Sٟ,��9S>h��o��n�I���#��X�O��O8�=�OR�Aqo��CΨ��Ȁ�P�؍}�)�	��~l[ЄW�z.�z�_+!��ش���*�3����7�+\u!�Dc��� IX��h$��*�=!���yAb�1k��� Bgk�!�D9;\���(ʇU���goi�!��0�����B�ks��`&X�!��3n��p�P�R7Xtp� �i
!�$Q�'Ʋe
��K�9�:pz�
ʔ�!��/l)X5#�O�:m�=Є�ūE�!�$K
A2�V2I~�x{�"M$Vs!�dO�������@S
����O`!��Ao,U )Œ&A�pQr�
 %d�O,Q�$�J����	"]��y�E�KR�P� ,F�h1�1�!/���7DU6�W�Ly�a��C�t���"�M�DY24p$;��4(4)x=椨ԤA��o�D�NhUÀ�o���BD�O�& ^y��o�X!$������s���AG�u���Q��F�	 .���C/ �D��&��'Y�#<Yϓ 0�d3S �"O. �"��!�ȓJ�d�A�ʃqk�}��J� %�Q��Y�Q�rI�dn����B�\��@��<���a�N��S�.�����M#���ȓ �&�0k֦���C3���0�����_@Y���	�2܊$�	>j����	��sXn�
���d1��b���6�[�r��b��;�de�ȓ+��31�����6�t]$p��rX5S��|�$B#��*ʢ,�ȓ	leX*��f"u��S�"����@�2i]�=ҵ�4�ʹRFp��S�? R�)�D�."~��RfƘ�N@�D"O�0p���wK<3GG\Q�b� 6"Op �#Q�=��L8U�D�{��|��"Oܬ��V�4����Cx%`"Op���*zX>��B�%<ʼA�f"OQP���@��<;#���z���hD"OV]�C��$3���ϖ'�<ɪ�"O8x	%�Ւ9��T�%��P�v"O@���Ub��En�2X
��"O���a)V�C\����j�>CR]��"O������9���)�<\*�"O���wE��U���R�G�' ���"OhU��.J7?�F��򋝟uR"O���(�}�H���F�Np)JB"O��)gf�0L�yp���%�Z��@"OdY�t���+�)x��\	"O�m��D��l`|�k#h�.�Va T"O�@Ѝ�{e�0R"hؑI2�̀�"O�$���C�V�)�MP�2�R*6"O�ݲ.[��t��
>7�
�s�"O~��mX�r���WO��D��"O��QV�{� u��JعWmz�5"Op��^2s�J��J�RUjl�"O�!��� �"��sc˄Y����"Ov��%�C��||z�D޼;B 1X!"O��0X����# O<�A6"O��%�:x�!��eΐ\1�"O���R�B3�� fA0�E��"O�h����>���B�
��*����"O��#M�9,ԕ��)G'}� ��"O�лэU�gj���A	���"S"O2��ݧh�V #� �2o��Q"O�)�TK�]�$�O�-/�>�Xc"O���O08���z - �Iߠ)�"O!��0Y����Nk�B�r�"O�M*��Ӫ�jPY�#¤��E"O�t�mշ �r�8��+"����P"O�L��F�{%�=lc*��Q"O�%�.@z�����1{v]RT"O��!��0�b�ģ�,Z��"O�S���RԠA�FÃ�S4��8�"O������36
���"�<mмI�"O�	kUă.Q��TCS�Í��"O� "�F->�����/.g�~�iF"O�D���Q�a*v���ӛav��"O�ä���y�,
��?U��"O��.\�,���-@T kRkɅ�y����U�ܨ����h����y�DŁ HK��+jJ\Ј]��y�d�2��	xԇ�&�\0" �2�y�χ�k�`@��"R�'rN�@�9�y2GƫJ��ĉI����O���yrb�I�f���ӊ�v�	%C��ygE�td&\[BB��}�����y��}��E��*� � �bE���y�5Ѻ��ī|6���Q�yR��-��b�mtԞ��Ѭ��yb�A�\���D��r}�+� C�y�e�5�J)ЖAęc��yK��N+�y�� <XЅ�«U�DQʷ%��y�#��;\�ьȋGdm�G,���y2�W"<ـ��@�7L�p`�Z��y� R�"�I�'
=6��)�#��yb�$o��8�����3�Z�hf�4�y
� ���a�E!��#BE�2N˘�2"Or}��(V��^��ġ�'(��x0�"O��x�o�2��
�J��>�c�"O�ɡ�	��\Q�*� 	Ϛ��"O���N̈́`t^��lѰK�`�	""O��@V��hچ��b�F

 �v"O�̀��ݍ'�	��
m����"O֜hG�ЙT1P�1�B�?��Ȃ "Ov�cэF#A�j��t�K;\�Np�#"O�yqt��0F�2��_�K�����"O~4��+�i��u�0����H��"O�ȷ�T]I���q��l�]XG"O�(�#��|q>\{������"O��(Gg�cTt-a%N޴N�^ْ�"O̐:$O�P%��m�Uh&�b"O�`�T`�s���U�X){b8Y�"O(��E�W+(��L� PThQE"O��qB�I�>}j�˶�j;j���"O��A�(�w�Z�X��	R2��`�"Ov<����!X��=KGL��p0&`b"O��r*E#d/�����G,P�Yj�"OK#m�����C�?�^�"O>�$�H?аt���&�1
�"O�H&���t!(�b��S0%-;S"O����&��Q�ɣ#4���"OLApщ�����6��� �P"O�+��=JWF�1�e�	>Feڧ"O�4�4���?KP���?$郖"On�YUm���l�$b��d+6�s"O��3��Uv!y��H5�5(�"O�=4K�h�����!R�W����"O����#�3j��b��0j	;e"O Z4���D51��ƕ^cfm�"OZ2sn�pFD�:�O�CEJp�"O��{�n
�\��܊�gܭ]).��"O,�3�+�q��Arc��	u��A "O�4	 A)����!jņX����!"OjS$h�6A��K$i�6l�"}��"O m�nB:=�8h�P�h��$r�"OȘ�Ƨ��sy��P�փ>�L<s�"O�>;���bn(=�b�A�"O��`�CK�oH8�(c��k����*O����`ؿL��r E�T�[�'ֲYѐ���2l˂g�PڒQ�'�FQJ�)��䀡a���3/X��
�'fZqh��h�"�!�
(b�<�I
�'nd�Z�f�"�����ϰMK>͚	�'V�p��\(�t�ǌ³?VD�A�'�E!�֓X:
�@7�W7��`[
�'Ω��.U�u��Y��z��
�'���Q��/=�@���^�b�t���'W$� �dI�;�l8R!�0O���3�'w��eG!T�e�򍊗PFν�
�'f���f� AD��ѫ�H�F��'������\�%���H&ԁ�
�'�R0�L"FwV� ���r����'Ȗ�A�܂8�����lа���'ȶ�y"/�wġ2eˎ/4Z��'��[ATU�"�i%F�0��}
�'ܔi[a	E3+�"K��(�z��'� �j7`]�,�N �đ��z�;
�'���b���&��@0�� �$���'�8E E��l���J5D�	{���p�'��tf�K�3MF����lf}���� ����	���@q���3�(l2�"O(QIըW$r��8�D�	f��
`"O��A�іxI��� �<�\h��"O00Q�70A�}+�$N/(`Y�"O+d@�e�V!,��\q ��.�y2+@=b��!���""�
�b��yɜ8;��0��!������Z��yB`�뎤��E�K
�R(�0�y�l��Mo8Q["�D����a��yB@�#�D@��7x̠�搕�y�h6��$Z"�^�y���A�ņ3�yR@�(-p���Q�n�xqi'X�y�ؾ+��h�����3(N)�y�ܝBpf�j '�H�u����y��+Y�J�@��6"��b�Ά�y"ƌ�!&����9to�������yr`�D�ȓ4� �g#&�{A�G��y�I�_`݁�GAg,,<BBj�$�y� �#gY��I���X�"@wa�y釻J8T���%#��P���y2�ћf�.�*scM#<id@���y�� k�
��$\ANlz.��yb,O�.���D��UP2(�OC��y��
�p����� A3Q�����Ͷ�yB��n�T���!��5h�8b�]��y�$v}�s�� ����a��;�yr�^?*��55g^?����0�[��y��R�t?���d� �RXd �y�d߭K�T�g)9_��J6����y��6>#��b�G"u)��;����y¯\&G��	��)��$�U�Ǩ�>�y�D�5)��cҧ��r5ƌ�� �yC��dN�a��S�oN	���y"l7'&a� B��hh:�.��yr�N�@>�r��
&@�s$�F��y���9��,;�"H� ƨ�+� �y��@�OI�4�������u����y��:7�n�V�	┽�A�(�y���
��L���L��d	��y��Y@�qQi_�J�>`����y�F	:��c/�%U������8�y��ǆY%$����µO����%�y©��66x�k�D��������y��M:*/H�q� �F�����f	��yR�~*A���9�R`:��3�y�
W��H8�LΏ!p\v����yBF���h���z3T=�%�[�y"�Dh��𢠉q�0�T'��y�G�[�1H�V�d�"XCi+�y]5_�渑�	�f&L9ٔ#t!�$�q�x�WD��e��eqq�ڊBq!��j$��A��7ux8Ԉ�
��6f!�d/v�������,rR=R� F�'f!��G�$M���፹t�����ԜML!�_�w��z��Y ��94�z9!�'G7�Ո�*�F?hѤ.I8/!�6T��B�02'�]2�F2& qO�P'0T�������6J�8��|"�ֈQv9{'�A),�mh��yr���Ko*�y�� r�B����W��y��M�O���l�":o��U$B��yB$��>Qԑ:�E�&*T2x�Ȕ��y�h]�orhQ����R�\���!��y�
U�	�"L�B��T�*\��yb��- ��8خ
�fI��/��y
� ���6�I�)���c��ϙ}0RDJr"O�)�	�;��!��D^p��"Ol��瓣<� ua̵�J �"O�XQ�g@�hl
����y�L%��"O���b%�9qw$L��+�>� "O�����؇q���{��:8��"O����W�M��I�bG,d��K�"O�U[a�*6an����D8DP"�"O~��E*؄+>0��[Ve��!�"O���jV?x�՛���+
� ��"Oƙ3���E�>H�Ħ�<ǐ�!s"O����F
N�ԳC���1��s�"O�e8�jG�.|1�w+��n��$�4"O�Ջ5��=��ɞH�@d@Q"Oh8R�/ż`���7��.Z2��q"O��[E#L�@
ژ��_2��h��"O�h_b�8{���i9�"Ozܨň�)C��5�Ġ_�m	�hs�"O�D��/]�a��Qs�I%R�0}��"O���@��$�RF���@["O*	�,s4�����èi�½��"OL�"���,�p��0E[���+�"O��q�AP"����Q��,E�"OFˣjT��}c��Q�97e��"O�e�`��m�v�BT�̡(+$�kP"O꩘T��,y�PȔ8��5�"O� ��`��F�YC�׷q�t� "O�|�-�8���H��E� �:Mx�"Or<"Q(R�^�RmA��̄s8 ��"O�����ɑ�예 ��O��"O�d���7[�t[d	�:HA�1P""OrM�J�)V���$h����(˴"O̬g'�D � ���[s*��E"O��
e.lDj���ݒ[b� Br"Od����PԀ�����, E@�w"O���'� �u��胀
*����"O@�$D	-]"�B��A��.�"OTx9v,�:O�L���+G��"O��B��6Fl�P#�O��,���"Ox�ю�P�XՉ� �!P�yc�"O"�
����%-ӖH��T����	�y��N���Y6
X@�
=��̉�PyRHT� -<�3Sn�O��!p��e�<R��*a�=RC�ڙ?�Ʃ�b�J�<�w���.�T�����.�>�&&�D�<�$��T���qjP���Sg�I�<�k	J�����?�Ҭ��o�<i����LДcɾ�[�'�n�<�$���,�$	;�Y�'�S�<�flL�T\���� M�n��-To�<�E��d���×#ZԐB���l�<�r�%pPF��g-O��~����Us�<�S K&{�>��$ѓ;��ۢ�M�<������"�I����#�e�E�<�cN<
Kʽ�e��/B��D`�B�<����h�n�Ze-G� hT���y�<�kM�@�&�J3	�-�֦Np�<9��7w�n������ZW�ɑχc�<����,0�a0���hRpԲ�Kh�<�� O
��Pum ",���S���b�<I�%�"SX%���=a�����h�<��ԗ� 1�kŵ� �N�E�!��%95��j�(X�N]�����$�!���8%��A�dÕaun��t���!�� ��A��*8����J�U�"O�,H����r!L�ل{�s�"O0D3r��:�"�ó�E'���zc"O@�"��B�T�8e�'�ł���'"Oh �3*P�=Sl �bj��X�����"O����N�.�ts&�
<�H!"O�݂U���F��M2�(u0�T��"O:]���B	\��.ѨB�0�D"OƩ�1g�(ֈ��n��}��!z�"On�S�`_�q8��r '\�'����"O��S�s�"m��/�8�>8��"O��¢�H�}~��s��^R}��"Ox�p��M<&p�ؠ��ٕoB��Zd"OԹ�$iNJ�"Ҫ���E[�"O�J�J۔P0n��ǬY�T����$"O��x"
 � ĸҥIA�.�a1w"O�E�G�*u��XpH�7����"OX�H3h�nвI�O� �"f"O��h�K� E0�L�ٴTP�"O08��Z0��	r�@4Y�ܔ��"Ox�s/�B�.�!j�|�J� �"O�aP�Z$Hf	Aȋ�v�Kt"O|� ����M�`=�q�֝ ʆ��"ORq���ɭ0�F�ѓE�e$�TPv"O5B��!���fD8p�� �"ON0� O�N���.ǽ&4T� �"O��5@��~�X�
�D.�#�"Ol�P���6,3և�(,���C�"O`,����9G�sG�h����"O��`F��s�
���e�-���"O. Y� X;�����R,#�"O����3w���X��F�Y�xK"O��0"��[QN0;f�^
U��]�"O�)$��~x���D�ޚS$�T��'p��+7��W(�Q�H+6�^���'!(\"�a�V���㍴.$nU��'����D�
+R�� �g����y2�'��$j NT�����QA]m���[�'O�X
�KR�4b�9ڰS�69��@�'L��L[<"F�K���=f.��!�'Y�`:C�K�\��H�@W!Q�� �'�|����1�N�����FԈ1a�'Z��r�F�9��10g�U=58
�i�'���y�oO=)�.q���\�*���x�'�m���s��LP���*RBI�
�'�~C��4tJ}0�ܾ$��Y
�'�8�r�L�3$�T����>�D��'�np�[Yf:�"#��H\�R�'���b���:tĉ���B�8�>y�	�'m�2mR"s�(���bZ 2Ƙ��'�D!0+\�ځ����+��P�'��� i�?$�|����Y�� �	�'�\(
�O[���CʳW���z�':��u�#X`��3�� �	�'}��`g�00�����)�\l��'����e�O�7X(��/��&�<�K�'@#�$ѦZ$D�&�����p�<�PE�$h�|�@�ȚzZ&�5��H�<�ul@�_�Ƙ����*6l�R��G�<AAM<E�q�D&�$J�3�CW�<q�b[z.!B�uqd�˅h�<�iH����sA�;��h��˃l�<�A_�U窜Q�CFhJn�P�/�B�<�d�?q��=�&�P*&�^U�RhQ^�<� �,���'E%<P�FK�2�=1�"O1@��R�c���s��@ψ��&"Oj��e)T�QV*�2iȷN1�!�"Ot���h�^���
I�"#.��ST"Oh���O\!yD�! �"}��m�V"OLi��
�bF��!�:[��D��"O��(q�X'h�hl��l�2o�&��"O�Dh�ꕢ�0l8��"�.�p�"O@�:G�ڌ^gtq{G��aϺ�s"O���TƑgX<�J��V�_3n��g"O\�"v�A0k�f�����.���"O"�A�りTE���+	z´�2"ON�!�H\;l���B� ր���3w"O�1�bF��e�<�yQ瀣9����"O�p:`Έ%�pS�]���*�"OvA�F��L�r@��(��	8�"O4Y�ʖ�O�xѓ`0;���1"O�� ԍA��D�d<J�Nx�"Oz(�E��Z�P����J�r"O��墈�
��B��06��ڡ"O�(�մ�H�yF����,�"O����1��L� n��r}�8��"O�qx��[%���Y��(JA�=D��¡o�7�I�+B�Eh�<�#�0D�HZ懊.���Ǖ
=$��l=D�(y%�E�x��lU�F��U��?D�� @*��W��y!�$_�t�cN;D��z��6��h�����H�a�:D���!�0PQ�`O�Q�:��Ć4D�СP� �|]��)�k�B��%3D���E��@O��{��G�"��X��2D� k8tز1$đH��@�1D������)M���m',kڌ0��3D�|q�n�?!�蠢ҴD��2�'0D�T1&"K�'��\{��%\����1D���A�_*u�a�.O��m	��#D�@�E�~Bz�X�O�=��xѣ4D�X�����H1.f,�5n\�=蚌���Z����;V�f�R��=:�
D�ȓAX�|{�T�a]t��`(��4F���ȓm��9ɕ}0mj���F$B��ȓtAn|�e��v���SQ�U�¸�ȓ@��XQČD73�xHk��7I�Xl�ȓX4r�;�e	e���@1f.���v�,(W�ю&Y�x&o�05��ȓ��8zbH f�lD����(3�I�ȓl��h�MH!ft����*VF��ȓ\d��#D�y��ӓ+Z%�:(�ȓ}�t�D����}�a#�5/�A��3���9��9�: o)�4$�汄ȓv��؆jʖ"�����a���ȓay�Y�
_�{G�A@6�	)kf��ȓV "aԉW$��'�6�v��ȓb7�P�吹�� 蓪��]R�Ȅ�NV�� +E=���i�C�'q��q��d�e�K�]`��ې�ˠD��ć�_GLգ��
\��|��S�/���z֪e�`(�lhx�f/Ɨ&*��ȓW�^	j��2Z$��g�J�V81��P �A��aȏ;�� ���$��ȓs�la#��714�q�!
��d�=qԍ�v���a`1m>��S�I�v��,M
|6ܝ�rC��;��C䉡@�h�Srb� .U��W�N�s��C䉠{^��`���~>qH��MtU�C�)� D�A���&j<����H2E��"O�Y(�l�!�B4#U:m:�	s"OFHu'�X�zM pk�<0��@�"O�\��E�.tY*Yq��<[��Pc"O0e�l��|i�!�Ĉ�0=*�h�"O�"����셄�g��H��=^�!�d�r��ے���;�&U��&�s�!��Z>|
e�`.H�5�J�0�凩!�œ.0��쉺]�be�b$�fY!�d˾R�2��ӎ8?�V����>,o!�$
�)��T���U��-���	$ZU!��\
yi�M DQȥ���\�!��@�C�����MY�,!e�
��!��0�����l�F��#���{�!�ϪI$(d� mD�x�`q��K� �!�ĉ*�}B��>W\Y����0,�!�D��Hwň��%BZ\�d�i�!�?#@p��G��(Ḷ�#Z!�d_K��9d�E
^�lI��E8-�!���% �����L�fE)˽
�!�$� ���
w/o���[�x�!��05�2Ap�E1+�̂�Ոw!�DW�.��t���S�6ǲ���>a!�$��Ԩ�IueX(��U�
շd�!�$�z*��V��
�k�?GY�� �'���v
V�w|l1�&Csc��{�'A^<�4��x,1s���_EB@��'���ӭ��y ����: ����
�'4p��%$�5J� �UoN�t�8]k
�'��9��� ����+B��N 2�'��!!�Ð�慨�᎐y�``��'���L�60���C����'w�PC�M�,���eiU����'����G�^'1z@���N��*�'0F�QvEE�Op�9vF��-W�(��'�0T�6�G�"��E�ΦTr^��'!$�A�O��r�#àFƂ�y�'c:X*Q�%<���ɒ�˷@
�<��'���rO�{�V���kC4;��	�'�����ŋ�6��r�K�[�z��	�'�K�(+�Zyq��	�x�,�gQ�<aԀ�7	��$[��yG�PO�<1����	�� �;4z4���Mv�<�O.i���re*O�?N<�`�n�<)��G:
D5&=��9�Pl�<	W�̌_�d$����5�^�q�g�<qu't���!�	�O� l�f�	=�!�ZP]>�sA!Q(~20�c��!�$>x.�;�I�|h�=�s��cA!���3n��ʠ�MM 9iDT�j	!�$I/T���t'�a=XK ��!�D��1Q��R�mF�P� 9aQǜ}�!�$ٽx��������r�+��b�!���2d�D�&R��� �Z�!�$��@�e����w�a3�MT�d�!�31C��3�h�,�I��,�!�Ďy���pQ��;���t�Ѩ�!�Ą?B�h +b*T�X��D��!�Ě�j�<�����#�|��\	�!�	>X�(0j�	�*��q�`�=#c!�D� д1;������C.l7!�D=I�Rђ�׫I�[�CP�MT!��Ϩ/v�P�F�5if�y�f;!�D�/����R7��Q�NG�Z�!�� �1!W�0��j��߮`�~L�f"O��'IX4}��M(Ǧ���̡"O���r�Zy�h�҅��`�$(;�"O���&#5/�\���e6$E�#"O�`�t/��F��s�ɐO�~�H0"O��{��ٶN%@vd��К "O�T��	ɔw�X�"�B@��l��"Ov��0)�((~q��!So4AJ"OvP��)O�ಯ��8�X"O蠪�HS �����m�6t�����"O��6�Ӧ0�dm�VL�fvD"4"OVP�t�ƷN5�	���΍aO�x��"O�E�'g@
f�P�D	!	4b���"O���ƃ��n���B���7a` "O�X�mM`���iG�y
���"O00���/����b���/�1i#"O�ࠧaHPH*Pʆ#7����$"OT����<2����\3F�00"O��NK�7a��1H[���͹�"O�Q	�(P�WT D��[7>|��"OH�P�e\�n�*l��a^6h�pY�c"OP�`���VQ�<P�'{*�s�"ORI��(����R�e��Ȅ �"O�-xa���]!6�`�E�d�zl��"O�V̙"<D��$�w�4䲥"O��9%O�7���`J�"'�X�@"O��b��E+�nH	gh�ZaXf"O�֭�*,��#���`���0�"OJ(	R"�iL��SE˪6vq�$"O:�yf���H�)!���#DEbs"O�p"cWX_�$:�C��ޘ�"OJ�c� ԧc�����- �4-["Or8%��E\r-��	U����w"O^<�bX�^���
��E��"O�Й0�(�Kԍ$�v9�&��yr���j�r1�׀I�"`	&���y���6w9�6�@wN��	0�ybgל?#�xaCjV+l�D	���y�F�i(���	8g	DD���<�y�ɳ}�RI���u�������y��
	�Pl�w�B\&BɊ�	ܬ�yª
UR��E�S�
���$��y��̓(t�=��ā4�d�D�ޱ�y� �E`:�jT�('܌��O��y�Z�4��IB�l��H2C�N��y+݄]��� Ym�ک���Q���!�S�O
���o����K 'Մ͚�'��l��lM�0������h��m��'����ߵ��P�"C@�~�<i��ïS
t�x��E����~�<�烅$;����ŗ�U��2wo�E�<A1,#q�RE�e�؁t�شJ�MN~�<�5�G�en@;q+�>	9X!�m}�<�C��(i�qWo�7u�u�R	Vz�<q�o�1L:����˵H���A�t�<YQ�۳e7��D	_1{yF �@ m�<��!�"#6Q�G׈(��M�ao�i�<�l�t�.ɠo߆d�(`�d�Nz�<���
��&��Kn�跉�}�<��/TOnQ"T�q��BBR#�!�$�@K�ak�˓�]�ȱ�@̰T�!��2_9^ ;a�F<h[LЉ���'>�"��L�+ɲ1��囱a��p)�'E��y2�D�.2�(���Q%3�P���� 4��H��}��{R!>��l�V"O�-�P�D�[u��C1b*���{�"O�1�M�v� т�g�+;�� �V"O$	 ��aڂ����=Ђ B�"O�Ģ�
".�8m+����)�b\��"O@�Ԧ���E�+ݭzD�@�"O�ݡ5K�<E�P����2:qa7"O�`�u+�(����u	X�f�Ա�"O�A�ՄU@��(]���S�"O���S�D�F�9b�'��Z�*E"O��)���&~��bB�� �T�#2"O̴�j��241Jq恷<�0И"O�)�@@�>��@����@�\)c�"O�� �O�{�p���c�z��j4"O���&�4LmӆB�*8j�i��"Or����݃"�P����gĨ@!"O^����o�0�e�Yv�����"O�e`��-fWb%1G/�7_��"T"Ot��%*��qS�9�#�Id� R�"OR��H�8�8�a���M�f���"O�	��)#��\���|�|"d"O���B�,a�x��؁,��u�"Oa:wL�Ȑ����Ĵ�.�y���d�T�oH��#�y��\~D����*b�:ĭ#�y��E�z5v@��MW���WkA �y�	Φ�؉yQo��}�$�foS=�y�]�&E���� �@s$����y���u���"��}��I�)���y玄H0�Zv�Y-�|�3�yrc�'j781xEI׺b���H N�y��X�9+4�欝.a<
d��٣�y�����l1!�T�] B٩��[��y���kB�x�1��!`,��L���yR�c  �cT苠����y�G�25��s�I� ���4�H��y�(��<���{�Gճ���0b����y�_�}_ح�q�� ��L�К�y,�6|�Xz��R�x �����J��y�۲J;��[��]�^�Q�i��y�o�O��D�S�C7u;L�0�y��U�������;qBx��Ś*�y2+N��u��n��I�Ԁ�PybG ���Ɛ+'���5&�\�<���
O��
� ��7Z�lH�JU�<q2o�?9�`�" "5�d�Q��N�<)�&	�)랔���ܹ:�a�`Ht�<飡�/4����6jI%��n�<1�C~|���1tn�Q)Td�<�!�T nE��!ѻP��t��T�<Q�F�t�8������d�5�f�<)7�B��&FazR ���v�<��E�A�����=F�4h���x�<�u�d0�g���-^'^�C�I����f@;$D�M��b�>C�I�qy����H%�m���Oz��C�I���@�G?�����xC�ɶt��di��[�c�P�Z2oã �ZC�ɐ{�QÊӚ5b����B�@[rC�I���h����t��3�A+U^,C�	(-V�[P�6��͡�d��VVC�I�l\:���E=5�����1.G2C�I?V���Ɓ~D>�0�E�X�C�	�j۬|x#aN�M\2!��o	,� C�)� ��s�a=Dh��H3W�(�"O�T"Ĉ$�21j�<H;V�r�"O���c/�<�l��"i�48��"OPQ W+�%xSHY�⊋<A��� "OnȐ�(O2FL���cڋC����u"O hC��OGZ�=B���p��)"O��I�L3h���P��Y�[�{E"Ox�;p�ѣ
��4&,��&N�b"O�(c@��*2:Q)��ƿ|�qɇ"Ot��/[ }_~"�)�3=��qZ"O��K��)�([�Mq����"O�D���$38�`�'6�j��S"O���5�Q'H�h��5�]�5h>-K"O�Hc��>nZ��ʳ�X�g"�3"OLP��)WII��,[�,[{"O~L���_�,u�A��]B��s"O�%�fFD�J��h��a�'K��@A"O�1���jzhM�����T��"O��G�Mo|�ya�*C�J��i�"OB�{�LX���:4�����[�"O ����L/$tE���t���(�"O�@r�D�.��І͌�;k�I�""O���W
��!~)[�[<RS���"O���K#W�, ��	�a5�pj"O-����>T���t)�$\"����"O8����˩V,* Ѝ�yA$� �"O���i@-{��D��+	�8D�Pzv"O��Ɗ�c������]3t@xK"O,Zrn�\���$� z?H�Z�"O�ۣ�ː"���$�G53�2 B%"O�}�v�D/h�+��ߠ3.;!"O�R��MlP�f�!>�m�e"O8� q��)���8p��(Q�؈q�"O�����.3GP0���`����"O�a!�	:5ܰ�PᑻZ�t"OB�)t�vbƜ�B@Ѥ���j2"O�� "�1�H�e��Z{�i�"OԀ2���m���y���"O�Z�NA�2�$�x��Ͼ=&d �"Oh9Bc��m.؈�'Gu@|!p3"O�(�Iw�Hi���a*p(��A6D�kC�Ժd6�#�Ή	^��Ł�'D�4�Gk�'����B�<���2D��q��׌uv� �'ϔ.�M�3D���2 �[��������
1D�C�%�,ZP{�E�z!�`Q�,D�ԪP�O�2��3AL�!�X9��+D���˗�W�`!���H�B��@�+D�$	�/ơa�аRug�'�t�Q(D����>/�� ��`xh�l0D� �G@Lg�� r^�x��1Ao1D�����Y���Z�!lr��p�/D���R#J�?*|dHv
� C2� �B/D�D��E�7�P �e�4j��u:�+/D���S�K5W�4�ZR�� ���6�(D�Q���f_n�e/~F%��h&D����ޣmz�5 ��� �Ҙq1I:D���i[�)y��$E_�K��X
!<D��8 �L>�~�3V Hf�|��#'D���æ��:v�[�!ƄswD�6%T�:�#ܔO�E9Ң���� �"Oʤ��%��&jXpR'P*�8IKc"O<=��/Z�B8�H���S�&uB ӧ"O�8��%k��)&$D�xX4Q0"O� � څ"�\�����ᆺٞ0s�"O���b��(��w�0f�e��"OtIBf�RVH�P&��OO��"O6!9�ObIF@[���B⦁�y�Ⱥ��Xid��>H��0�A�]��y���T�����
�n�6|�� ��yr��!3W��j��Z�]����yb鋮uX��j�BZ�g6!�P��+�y�K�Yu�5QU�A�s���0 
��y��I�.|���E�D4c��A�E2�y2��41x����̸\�z�S�'�y�怭0�~��g���AHN�1����y"��7i��ITlڅ:�`��3$���yr,�n�l{�&�4ڪa����y�Ā
(��9ya�P�0�9�u�'�y�ۗ:��;F�V�3 (P�+E:�y�Y���RnY�*fl����y�V?')
A���@�D\Q��I���yR -b�X��K;�JUX K�y�+�MO��jr���$�/��y��;g��8���J�MP��F*�yҧ�RۄAY�G-H����+�/�yB���:=���q��8�Ń��y�耀>�1�'LǠpe��hX�y�$@|�sFh��ѓA��yg�`���ZKJ]O�����y�i�4D*:u��)�"M�v�j���7�y�E�)<�TmbNܵ.ɾ4���5�yr 5Π�q�nJ�#��Q�Py"a3�N�i�#�mn� ��J�<GI�* 5�y��F�p�����C�<1�U�����'�H�aʕw�<�e���}M�����A$Pʑ��Cq�<Q��ץ^�L5�'a�<���l�<Ѵ�G�K���Z��N�s�2�cgc�<I�G�p�d���.=N�#��t�<)t�	?PL ���(�<`�D�Es�<Y�E@�x�^	�UKҌ�`�B��E�<�S�J	B��Cg�
6��	����B�<1��P���"d+nt2a�]|�<��I���؈�Oۦ:���A�|�<�� W\���#Ǌסg����E��v�<aÁT�0z�� P
q�81Ӥq�<1�dF
|p��p*Ŕq�n,Y�a�w�<Q�)��(t�WeO�jw�)�g�\�<�t,�
p|҉���D�4Z�U��Z�<��C
�tl���ě9	`���QW�<9�&%Qm��Xn�x���S�<)�)�6j&�*���zP����N�<	��R� H��ӫpA�uXeęS�<���4a�ebE%	���ˆ�Q�<�#��*) �k�g^&=����.�F�<u� �Qp���c� S�:���C@�<���ru�yY�Ƒ�@�K�&u�C�	 6�k�L����i�C�O�C䉔q���!�Fͭa7�,�OދHC�I�uV���˲hd��
H<>�,C�
|�A��Tpb��Eż�@C���!�G�>q f�(�p�jB�	�R�`dBC�	�O�nX��.�v˜C�<�n)*S.3-���	@��^?PB�I3=uR���E��hn:����S��C䉨$��Y�4@X�� z�"G2B�|�.%�C�C&l���Z��N���C�)� �䢓EQ?���26gM�HH�� "O���dƆ|_�y�Te
;_1n|!q"O�WK/q��Ǝp�l QJr�<)��:t�c��L�.�D$�DD�<�Ս�;	�~,R�Ɲ	k��K�g�[�<q�Oٲ3�$HI�!BD;����<7$�)*��-��Y�+�<�2�KA�<!��Z$*�k�>l�b�9P,R@�<�MA�~n;s�f|B�C�IWx�<!�G)+a������1AѶU�K�t�<����z�Le� .)qU^�2��Cu�<�a˓ 
j���`m����_{�<�c�27�P�����0s���BI�q�<�Q���J[,��aŝ�uΖ�[��l�<�6�L��,m0w��X�VYyF�~�<9$KAO jPhPoЦ��Dq�P�<9ݼ1��c�� Y<�ts�#C�<9�hӹF�����&HN�)&��u�<�3k�R#���ߟv��M{#B@g�<��O�eB����]&aYT�RU��f�<���(}F�r��C&	�8`���z�<IS��08&tb�e�EM��ɧCN`�<q�m��Yk��z��@}��8JU�_�<�+��6r��"�T�����]�<q���#�'��3�<�T�HW�<Qf�R�@}X���nF�@൐�`MU�<��I�;G�� �J3a��P��H�f�<	��=1]LԠpׯU�,p罞!�䕫P��hC(ٜ%��ɰ��)�!�D�W=��R�@_�QT��XU�)�!�dG��¦������Q�	�!�_�|P\�BD�C���@�)ʲ)�!��^8�i!@ f΁"¥	c!�$
�� �A�ŏlX�Yp��,#!���0=`���&͝;S.m�Dd��I!�� k���kP�"�r����>.�!�$V
ž��dn0>\���!�)V�!�D�,)�hHT�Ϧd@��jbY R�!�t�~H�c+��2v�jf��}�!��A�T��)U�B�*��9H�����!��Y"Kt�ר�+u����ϙ�yn��$��<s���=DpZӆ-]:�y2��^8�u��W?%���q�]��y�
-��r���"v*$h��ɛ�y2Ň�|�RL $����� Y��yBm��8p襑sl��h�����I�y�g[<���Sk�>deh��B��y2OH�X�: �U��%[���(�y�Ʌ��t�۲)�*Z��0;�#Ʊ�y��O1I �IơFM1� ��߯�yB��<����$�Da����y�T=��y{�Ǘ�D�BF��y"�5 ����� 	t��83�I��yb�� �N�.��	����"�ڳ�y��+����c�$q>~z��X9�y#N�]zQB*jC$��'
7�y'O.
�#�
�c�=��	7�y�2�t����X��wg���y"���	,@uR���N�HL�qE]!�y"��~v�� f�R�oh(	�h�$�y�o�u��H'
2� �	�'�0�y�@�o���K��0yb��(B%ަ�y��X4J��d픤({�!1�K�y" K�dy��seҞU�n-ÓO!�y
� lQ��݊�ʨ�v�֠@��m�"O������'�P%�%DD�o!����"O�Ź�8MG�$��"V;<@�"Of�r�䒫�l�e��G;0ɑ"O~Pj�%iwP��@��(� ��I��P]����i����AsV�Ұ.�<`y1�[>������O�h[����S�huiŤG@`˳� >���JJ"���0g-JFײ!:sD��HOdk&�X�L>$�'9Y��9H����T:��G��G���*W�3X�4A�%AޤK��̓ti�O��$������F�oN�i�Z����b���4+0A���!�i>�$���'���xV�Q�0�zN��I8�@�Û&/fӠ6�	�U�|��-Y�t�d ��FS�P`ݴ'���"3R�ܖ'���O�'�'���z21iC�\>EB�ʁ�ɑGC�ć�&VM�3�X6,�J�i���Ͽ{��Ko���$�L�;����l�ʦ�E� C�����x������w~A�t@�4{�1�k�L�dK�(ɢ̈*%� 1 �	s��L	��?A��in6��O�#~n�-
G�eQ�������#��| ��ß��'ayb����ȴ��[?�	�%E�HO�7���'�(�O.�rhQ�F2��*E�ʘ]�HQr'A�<�Co�7(k�v�'̈�{C���@�*S��@K� �D �(0	P����X�F�2k̊��ψ�O ti�i������;,ޖt��N_�� 0P�+KLV��q�D�!���ڦ���g�ɽg������7a~���T>s��k�(+
!H�aݛfI�t�,O��ķ>1g��v���To���%��A�h�<!�  2DÔ�^�~�Ǡ�,#�� ��a���oZ_�	�����<A�����0Q)��?��BcωG#���E�_���<I�GpDX�� �h�)J<1�|��CÛ#�  `pN�C�H: ꋝ[R�"?�%&��Aʖ�#D �d�Xxap��;M�m�c��3r�~�A�,I<gd��ѦF�Fx�!�?�۴Px0�#�����Y�T�X8�jPlD��͟\�	[�IF�S1�~��P�I�A����$G���IE؟Ԓ,A�.T��[Æ�*,a��r�A��?�Ҵi���'B7-B��mZ�t���[b�Q
i�t�5���q��a��B�B��?y���
�L���:c>�Tb�)�#%�擩X:����,R7H<��EOr!�#=hX�{�
�FR2/JV��s����u�'��-�U��.-Ԁ�b�se��	!l]p�d�O���	E�����T��V%S�	�d�7�H�eά�D6�i>�Fzr�8��Q�ʕ_ �8W����p>y��i��7�wӆH�ьW�O��6�F�D�����Oi�7����	Qyʟ�O%Q�&��M���4d>�5aTk4 ��caH9j�����P
q���x����W蔻Mv6y@�E�o� ��k���M3�O�=�tH�c��OC��{S���@��̻��e�����X�Uƌ@��H	�f��x��˦;���ON��_y�����V��?�8�I��+Md8����~"�'�azR�O`{�䎖%Wj'<):Ф�M�Q�4*�4(���|��O���ʿYP�t��Z3vJ�(�LT� ��4'��퉏e~p   �   9   Ĵ���	��Z�:tID:,���3��H��R�
O�ظ2�x�I[#��C�4e��B��.�=H�n�,��x�$�#f?V6͂���H�4;p�1��\�I�$U
E9�`[*P��2A
��l�tD�UE/�7�T#<)�&i�Z%��MX�J���$[���DX���'e �jm�,6?i��K) ��6Mp}"��t�Lc��&q�N�3�jAg� ��
ry�.�OB�6d����9On��$J�)Q����Qa�dL"D�#
(6 ̋v�H���D�==�������'���D$�q��Ȫ�`����H(��%����3##�'(����Ð�> ub$��T�M��'��Exr`X^�'��E.��!���Y�P����(N.#<���>ѧ*�4e@>a����Ty�F.r��)�O�ڊ{@�Y�V-;��ΠZ�<K��F�Ms3�-}n�"<��/�G�ld"sf�|e�Z0�E9Z�p�>�Vn)�n�4�t�xEY�(۵#H��U%��0�� �'(��Fxbn��nfR�� 7{x��K��Y�0վ�a�:$"2#<���Ox�$��q�E���6[�ٱ���OB�8I<Yf�;t5���Q�I^��p��ZS?Q8�\�OR�I0K��p�"�Q�Љ�ޢ4�.���h~r��97�]��4*��ɏ1qࡉ��OT�qakHn��SӨ��
,MɁ���H��܄N�Q�����>%f߷&.T���	 ���3ǄI}R��j�'ѪGxr�H�s�NS;2F�� �%�y�n�J�  �O���Q��U"�GUy�Ne�
�OȔi�)��8�L�)�A�2�"�����Y��M�@����nD
V������)��3� ��w�?.��E�d���V�>ŉ&͚0�?A��:���<�'�?���?9 '�!1r`hlA:���`�O6�?i���ċ�	����۟ ��̟P�O� ��F���ӈ���t}��OJ��']p7����O<�O76��U��v�>e"i�%cLY�c�aA��4��(�� �̒O����>A�#��19�B)(3��OX���O����O1��ʓY��O�=�0��E�F�;!&��em)C���*�_�H��4��'-&��M� �z!��C�	����yZ����a��od��Y�a�|Ӿ�|#�틆I����O�Zc���p��@x�`�:By
�h�'~�Iß����	����IV���3e�4�I�#���@�syB6-ջZ!    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �   C   Ĵ���	��Z�Zviʗ&���3��H�I�
O�ظ2�x�I[#�<��4d�v�V��$�s�ի-h�K�GЃi^7-ƦR�4WU��!��U��) ��|�t�G�,�B�Bc"�3���uH4�,��"<�hӐ ��g�
8��b2�Yo�p��X�`���gxN�Ѣ�*?�W L0
7m
P}R,l��)s�R�9��\�S#Y%B���k\6��aqB�X�i�JC�x�+��,�k�
�tj���@-Y�x�eӋ��F�� �'��5�����'r�[%C�^:�nڠ"S��PM�p�Z�Y�ǁO�(�O�����$����u+��
��$ӬqU��-�Pp��"<���>�]B-�S%ۻ[/�,���К�M��I�)�����Z��20���3j{AM�3�8�� K4}��e�'���=�LB[|��L�-,��A' �⦵��I����!m��o7����R�ԅ1�Q�1b�0y$�	7&p���m�j����ؿW��@�GJL�T��˓��"<)� �	�f�z���@<i 4���	��i��ɮ52���E�'��Г'&թ]
9r�ږ!����yRi�'�J�$�T�7;%f�;�j��T]�aX�����2S�ɄZ��'�f�ɱ0�\P�+x��f��O6���~~B5xt�l��4��	S4�x2�O�T0B��@<L֘aI�ߧp�ڑ��Y�T������c�X��Q� `�'ApE� \E/�|� ��[�X��O�)���䃼�OHt�c`A�M�����E	'Ӕ�S�'�@ �����d�5�?�!\���ɬ��ˣ��&�F%�P�l�L�������/Q�
�B�{yԠ��ĳ?��'�de����;;ب8@�J4�|��'�I� �I�������0��w�4��e����倗>�Bh��J-
6��B����O��$)���O�]mz�IBɆF�
�{��̧L���Ċ�����z�)�S)G����b�$��ԜTDi�G�x��@���h��IE�В��$+�ĩ<����?!��1-����� E9D�	�7���?��?A����$���2U�C۟��	�hh2��^��p��0c�*a�n�D��3P�	ޟ��	p�)� (���̔�4Bx����$�5�g�����ƤXw�QbV�W� Xs���O �(wNҊr_�AQ�٤�r�t��O����O���O��}���<�F�@�kͫn'�J��3p�y�����֠Q    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �   F   Ĵ���	��Z �t��8-���3��H��R�
O�ظ2�x�I[#��q�4�?iU/�+SM�	�pMW�0�h<@P�\���j�6Xoک�yb�$6��[EBhR e���B!N�v�9R��Gu�p�i�vu�o�/�z)���&pF��'�DA�.I�$�*O0|B�99#61X��9��ϥ�̘2���5f̴ �PBP<Z@_�L͓Ooք��Jʻ�ē%ha0P8y�l�3��y�D|�4�%^�態wH�<)�k�����&�����nu���_��YX!�+)
�˲%S�?4`g�5��L�OH��O>	�/�o��z�&Qg@�:�V�<J!i �"<q4m�fWd�G�Nz�<�#�����̻��I�y��əR����5e�9J��,Ӑ-�ۄ�'k0Fx�a�Y�)��	0&Q	t�3(_�,lnڭ:��X���I6kH)2�����FG	��Ȥ���/�I2� K����P�L�L�XɆKǺ2��5`%��<�e�$�R�4KԄ��_��lb�l��P�������D���a�	%}��G�9wH|�,I^�ܬ������'%�PGx2�Dd≋wD�{�Ȗ|.5�q��	�EI��D�xrn��� CIJ�G�n����N=��(��o�O��'De�aߌ�M����9��Ҕ~+�ŉ�}��Fi�F�Ƀ���.�剄��I�1��L>���'�xb��<=�`/ݤ3*�������N��O��1�����
@o��d�x���R/!�$��#� �  ��O����<�O��c �ۜ^Fe�0��b��Pa�zӮ��g.�S�1O>�	�n,�E�Ր
thaäj�!pt��Pٴ�?���y�FGh)�O����PR��T��ŃKզ�Y�&I!lO�$�OB�dv<��s�CW�X�"z��O$H���o���`I\�ē�?������f	<#9�gcH�F���AQe�o}��U"��'v��'t^�LRC�){��U�Vn8�eA�Z�(�J<Y��?�N>Q���?�ebD�&�z����B6���
r�z��<���?����?)�O�ܠ0�Oތ��FƋKL�PQ.J*#��ݴ�?i���?�M>a��?At�J�C]B�l��Z'b�ru'[�f@R��/��|ꓥ?���?/On@B��J�D�'+bU��Oތ�8��.L�HD[RdӢ���O0�H��7�I��������`J     �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �   A   Ĵ���	��Z�ZvIJ(���3��H�I�
O�ظ2�x�I[#���ݴjk��&ֺ+�j��'$[=Y�"�a��<EV7�����4=�$>��E�	�!��l��d,)���Q^�(p��J2q��"<Y7nh��(��+S�@}�U�A��P� �3+��@8l^hy��ćayL���D(��D;W�,��H���R͡�@7`���0����D���/R�-&��r�ʛ�*W�����E�Op���G�V�~ ��|2!��'�pd�K>A��� �� ������0�OaZ\�Qe��M{�D�'��ò"�i�'��d%��o�ܺ��
C�\������yҸn��hd�� Vl���� D��2�"S��]���$
<�O�Ey�O����K�$L*{�	>0�T[��>���,�u;`�`��R��V�r���/�c�d�l\��d��O�MH�f�@[���nҼ6�$�ע�<�O�������$j���J�~&��ѫ��\��!*��p3��Ċ�f�.%�؄���q��8C_RY���T��O���E׶����Q����4k�%����<3�<�c�O�L�0�|��Q�  �L��Q�OV�ۉ���
�����ѥkdtMi��2�� y0H�ZPr�WUy�d%F1fA��4���W�\ɩ��Of�ٓ� /G�dأ�L`eh�qS���/��1Y��O���Ư�=A�'�8�y��"���1�/��U��O�9���_��O� V����D��,۩E��+�"O�q���  �  �"O<�iea�F�8x���-?��k�"O 90�
�(O\x@��D�Hks"O�虷�K�?�|�/E�b�0D��"Oz�:�a�$���{���T��t�Q"OjxP�Ł�a@�c�1y_��0�"O���C�Ι0���p�ၑ==	�"Ox\��AT�tQ́@7�7i6���"O�)�RKD�SK=Q�	
��p�"Oި��k�2"G�p�vZ:u�f]�"O�m�F�ܙn�@[���,��Qd"O�0,]��Em�)���Ӣ.D�D�r(C�D}��ɘ8QG�e"B��o1n�{�)��]������00*B�I�/�Rq�X!_��mawɞ0k�C�	8����W�������G	S\~C�ɻ9���Q�aG�Q�%�6G�$�<B�ɒb<�� à5�Vye�8B�	�Js�M'�ef��`-�' HB��wD�p%    �    �    ]!  �'  �(   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic�'��}9���p��"��hl"q�ƘRS ����;D�(X&F��;L쉰L��2�u�vF6�I)Yr�P9'��F����7pL����de�`r��ƈ�y�b?S������1bqЗ�ɮ:���1q��>��DO�g;��?�'Ҭk�F*`b�D�38.jt��'M�� ,�z>��iF���<�>��1�.A�Ȣ�kX�&a|"&�D�.M�5T����@���p<�0A�*kVP\"ǧ�#����شy�2f�.4f@E�P/Πc�2��H�R5٢��r6�;SD�BJ6��Ols�� f�mB�C�f��"}"��u�p�z@c��r����G�S�<)�Ds6����/��B8����͵"Ϥ2c��?z��$��o[�]�|�<i𭏏9��B�-�%���b�D�Q<i���/$�6d���C숋èK(Q�( A�cSI):���ɞ�x����A�d�����|VJ}�EiD��џH�G��K��X+���Q�~%a�'�$h���tFI�Oꔣ��[#u�8�ȓ>且#u�/L�4+���k���'<0֤̉�׬ �neH����U��D'8��%��7�B�ɥn�lGh ]Y��X�GI�]��1�2�푥M��{��/��!�	2�ȴ�C,U�{���󄑜W�����L6ȱ㓋 L�5��C��B�,�b�
~98 �N#{�d)p�>LOjR3nG�c��aGyƎ5���ɘ]9�R�J��]��9��ދԍ� 
HSpF�(�V�3�Nւ.&���"Oz5	B�@���SR���r�Iq��٣��z���ؗ�P�f@) �Ӻ�ƕ��ن����q��$&B�=|�-&�X-D��@S�AB92������ ���@���$�1%k*�3�	5��E"eL4LrP%c5��F��B���5�2KA)1�бcVd&i��Ag�O�&�v`��w�ʰ��+��1���8G�8\���	�3�0�ō�>7$��$��ZΌ��R���J�[�[�y�ƀ�\z�@��;�V`IG�Տ��'�Ґa��;C�r"~�#뀑/���a�	g� XCѤ@T�<!�iY�tҌjvz� ���2b�dI#�X@���H��	t��1A��96b�hrfMG�6�8C�I�}��Dp���b~�q�k�dL�6m��H��"W�'���₤�� �,�r��&
Jfp
�gzJ`��OJ�YBH�%���#q��"O�t��1*ؠikT�`����"O�;2�;nq�3�Y�+eh�2�"O6�1�Iߜ0c��8���8*u�-y�"On��'�I5*h�D�� -.J"Opm� "<.�V��eOʀk�l���"Oʠ±E�/J>HIp�L�K;�ܙ3"O��(񢌢Xp�H�m�4_!���"O�{��XR���I�n�Q��"O�Ə׶'�(e0@�ͺE��P�"Oq�A��,b��4c��XQe΀�"O� l��%/ 4�f��,H��yc"O`aH�̎��]��L�' �Qj�"O�i�bdł��a��i��3x0x	�"O� 2d?%����i��h�
���"O������er���	�<�d�x�"O6Xs�N�,���n��]�=�#"O���.��X�p�Q�n܀>���"O�p�V쀏(�&,[q�CA��p�@"Ok `Y�#�D��ɜ�s� 8�3"O�y���?��Ir�m��*gH�"Ot�`&�ߍa �<�T
^�fMv�rb"OȊ��.EP����,D@("O.���P%)=��ۥ�Dn��sG"O~XBaa��D�UK�<B�("O�9�@΃`r�!{�	D�l��v"O\��%î*����Q��2"O���u��$n?���׀))�%�W"O �PG&V���k��Ǯ0O��C"O �$"K.u E2ԯ�0	mV�d"O�i&D=(��R삽N��I�"O;�[&!����u	۠XB� �5"O�yp���1 ��s�!_�8�
��!"OW}��sL^�z�X����  �!�ʶ��؉ue�X�13FЫ_y!�� U��<qUm��e��d8�ǌ1�!�l�^�!�O�!1Zya�/�*2�!�]:Bx9aTW�T���/Y+�!�T-7�8�kC�VS��p��ϊ�Z�!�DX��:�p��K��H�ԦQ�!��7<:� a�O,i����k�Y!�d�p�E#���&~2�9@M� R!�D^5@R�QrR���y(��Ub� �!�D� %/2��VoX<V�]��W~�!�9}DyTN�1`$!�1��=T�!�ӬU���jUa��S_X%��GA)'�!�������� )AT�n=CS�v�!�DE�E���BY4��+�F�!��N�p'P��h���@|�!��Жx��L�EQ���!Ԯ8'!�� ����]d�����-pD�a"O��3�LO�vl I����1�@9�"Oh4�	T5	5�	�	�_
�8H�"O��6��&RS����E?#��c�"O��sw��1�I�2��?�@"Ob�[�m_"%�ܕ� @�(*��r�"O�p�� �+*XT��gB�+}��H#"O��ٕI�+�D3$Sf����$"O��s!ÒF3�|�'�F�M�2"�W�,h6��WX�p���ƅA�f��$aЏo��� �#D�0P���~@�9S�C�=A^���� D���p���, �4���;P��c7D?D�؉��F=�R��2��+~��3(D���A#Q�&a��
���Kl�$�B D��`�)�<H�X�B�Ms���Um(D��r��@�N����K/K�H�A�&D����� ,��9ۇEI�	3�k�8D���W!^ �C���K� �+6D��P��x��!D��/|�h�Q�2D��'��h����ւ\vl,U�/D�@�Ɠ#k�:9���Ӵ9т��,D�0Z��ЗT�+��E�v��y�'/D�)�]>"L!S�D�1+o8�j.D��se֦a����SA7D��Zi�C��M��ڃ?#���B3D��83MF�w?0����1���Ѯ-D�D:��
(y ��J�%\�� +D�h�f����ȃ�D|�%D�t�񥋝T'x�y����[�@@)w)&D�{��B�4QPp�˴6�`��:D��A�(�.�ȐIp��2K8D��;�m	C�h�6�K�D-�%3�m4D�����B�~$�תI�4�A#3D�T�Fh�)V���+Gq2���*O�k[t�2(I�h��g2�qB�"OI��!�.}]�A1-�}X���"O&0��AËE�\���޹pf� �"O����g��fĵ�@
_7�թe"O�ȸ��vaDԂE��GSx�G"O�y(V�M=V���B�B&=�r"O��z��͗DGv� A�>$+x0��"O���W��̽	G�� [����"O��"M�R��H��yR�9��"O�)�q��?Z	�=Rb�G W9&�1�"O�5h�:l�B(��� t���"O ��سN�1p`�Al���"O(�Q� �"J����.ւ�U�"OKp<Ah�a�S�0^��"O��z����C*L�(�LO>B@�"O�ph$��:��u�$&L+f��ei"Ov!'�>�.��A]�z�I��"O\pZ@"�$>f�Ѓ��7
�֩8q"O�@C`�:v^�`���(s��E�"Oμ��+e���q�J�o�T�id"OZq��O�GNu
4�Oq �"O����T�q��%A��D�9J��Or�<��Hߨ46��*صe]�x:�b�n�<�R��(���1"�	�u`l��k�<��D�tR��A@�2�;tPj�<�2*�#;���X1p���abM�<�g9������O�N�C��K�<n�%9ע=9q���:e w��C�<����n��0����=IR����AX�<�ř	1�5I ��<���"�^W�<� �U�g/�n��	��/�� "O��#��)Z�����A�HĔU"OPTbCM�% ���An�)�8h�"O�ă���4T�9�@�2��	�"O�̰ gU�a$*�P@ L1F���$"ODL; a0S"2հ��V3�-�q"Oh��D��m�f�e�]���E"O�0GN=4N�C�X�5���"OZ=h�NۜG>p\��h^Q���!"O�0�bf �'!���1�L��"O\c��=�"0`s��+5���{�"O�����X�R,�Ѧ�0},�z�"O� �&  DƩ�d��kd�pp"O:Q����3ڶh�t⁆P �P��"O�0�B�W=oj)p�
�]���k�"O���b�ݕe�f�6oG\����"OX�y@#�!g�ҡ5�]�@Qt�"O�;@�<���A�m�ntb"O���u�*>�A��!�L�2�z"O���GE>��}��1̘U�"O�1C5b.,��p�u��y����"O�sR�A*O�@��˓�9�"O�Dz�ĕQǜQaF��	f�`��@"O���i[�Um���I�n���{�"OH�:GeN��sv�Џh�\1"O�(�5E�OJNh�R�K���"O��!�e����&��\N�8�e"OJd�QaW�i+,Y慄�(ʨ�#"OVU#E���I���!#�ZB��"O��16ˏ�&ھp3%�_95(���v"O\�{�ǘ�}����j�Dv�:�"O�ЈC�X!ӎ�0�h�^��q�"O�4�P�V4uiMA��lq�"O>�Zc%P��Ӆ��M�*��"O"���� ZMn��D ���"O$c0��,!��;�c��hs�(��"O
��@)��`_z�
W�S�&V�;�"O�0A��4LG�%ʵ�=��<3u"O~x��k�4k����%��U�:��"O Qj����=�$@ؕ�?�BP%"O <yѭ2-9���W�qr����"O��ks���K*����ܬs��*�"O��� �Ϙ��CJG�lk�+"O&�K*�o���`3,�:35�1k�"O����
F�0`�낭e��Ч"Oz��uJ��~5�!�c�U�+�ū�"OЬ��.W�"�IP�]	���u"Ot	I��JvI� N� @�t��c"O: ��f[?B��`�W�%�pi��"O^���L8G�v�dmw��hpV"Op��4G��\�r5�*�����"O Z���}��lK4�:Air"O~���̙)|I�p�LЭ�*�)�"O� P��X;TȖ�c��]�9�6p�"O�ݻ��TCX���
���yK$"OZT�!�HɎy���ʯW���1"O��f�P�e%LPCh�!y���"�"O�+\�L	�Ί*<]�T$'ӏ�y*
�y�:��?�RpP���yҀ�й	"�?S��r`���y�(��׮m{��2��	b�շ�y���{����7 ن/2�h�A�I��yR%W�C��0
���:2�q���M��y2�ٮE��)�G,�P�z`�Y��y
� ��PO�)\U�=hE(�d
l<C�"O���U/��=���0H
�<��"OнFM�6:<��Q��.F�Є��"O�)���"ݖ\�� ӆ�"O�\`w [���Ƌ�_֬�p4"O��p�)Lj\�kQ*] 7Ǥ�y�"O�$y��փ,َP6#̺m���8p"Oމ��#�$�g��
!:�*e"O>���Ȏ�.�F�rQɖ;�z��q"Oz��,V,%ha�D�M������"O� Q)K���Z��O��9qg"O��e� 8d#�#����"Ol�S��$q��i���$�&"O��E�)C;��Po?/�.ܐ1"O|�9��J7z�Tի2ǜ�o��s"O\e�a��,1�����&Ѳ4����"O��Շ[�nd� ���*�$e"O4��eFǈo��������354�#"O���q�ڍb�X<tI�����r"O��3�I<N'xt��f�|`D"O���DC.rX��I"f�D�����"O�d�,�)H��F  ^�X�h�"O�
�e�e;X��7c�"]]���"ONس@��?v�H�ǂ�m]�X�"O�Sׅ׃_B}�Ve�3F���F"O�k4� M�,��-y9t	ڡ"O6-c��D!F�4�lV:5�X�1"O����2y�\�I��ȯh2^� �"O8��5�ۅ"lXS�`>@�F"O~��Ꮪ> ��A��(���;P"O"��"䙍j0X*C�ӡPv����"O ��Q�ne�T9�ը!��]�"O<�j&%&���ӳ6Wz�"Ox}i���a&��ñ��f[��T"O$s�)ɾ4�裂*M-(@Ѧ"OhEzE_�N��ea��*d*�D�3"O�0#�nK(KQ��H�撧60�"O�����0e��PKwk\$]�Z*V"O��`T�>b�Q�M	w�ܹ3�"O�p&-�(�F���A04f�X1"ON�qF��%��h�r� �U`4F"O䨉�,Y<zl�fL�8|�N�z�"O�P���:�
��3O�Y��"O��S���)4�r�C��_��x1�"O����$�=��u.���hI��"O�1�c4x��!� ���&"O�8��D h����Ď>�*�:"O���@ӣ��l?�	�-OWM!�d�J* ��햨jM4�M+&!�d�*��R�+Q&)P1�KǶV�!�$U�BmT��e��"Z�S��[!��S�^�x該#�B������Ö.Q!�DŮwD�3→+E�j�A��.o!�D�;{T|[��\$7#lL�Q�At�!�$��;M,@2�^�&p�a�9�!�Q8ך�э�2M|Q!���	w!!�$Џ{*8�3�ߟ+���wcщO!�D2*R)�叓W��t�e���;!�N��r<��"��pf�`t��B!�d$-� �B� ��zU�b�3r!��H"&| ٳ�EQ5 ������
�!�DJ����!��B'Z��Ճ��]�!��;sD��*ң�?x�s7c�l�!��'���$��)X����U �?8�!�� "�!��͞}�4�G!Cc�a�1"O����)��Űw�\?(� 5��"OT���A��[[
��Wo'�b�2�"O�=Jt�D�k��T�pQ�i�6���"O��
l�B޶���Ű.�R���"O�`�Ү�B�9u#Q�1���i�"OT5J`j��CE��bW{�xX2Q"O�r ��/u*� ��� #4��"O�h�'  k5"sAҎ3�
V"OVu"T��q�p`��TNs��w"O��W�	���D��NDL�&40�"O�h��!c�v��B���(�"O�A���2Y`vA����jr<�R"O�@q�  �   U   Ĵ���	��Z�ZvI
)���3��H�I�
O�ظ2�xbI[#��4nk�v��K�x���:�B١��I�Bh6m�ɦa����yB���<9l\=���*Ն ��&$��įH2�ãv��,�=!�C)��7M�,F��I�EJL�g�Ё��E+h�1O�q[��)��$5����^���'��SMT*Y1����DR4Ś�[6M��Dɖ'.J��L$RaX,]w;��+(t�j�B��H ���e��H�r�ؐ(
�I��<�"�C�ADD$����B��I);yxx��V�o�@�ڠ�C 5]0�I<xņ�[��>��b5�W�K}��"����c���rI�W�n��B0O��I��䇐�O����%�P�����L��d��d�'!�}Dxb&M}re�!9�`|�"ʭo�ۓ�ҭ��ɫ[��VRܓT�և_/0��\�b�%,�lZ55<���V�	<t**A���^�i��<�<]�r� �IO�����$��дI�\	ciL�r<f��`Ǩ<�w�3��P㟄��H�
n�P�� �:!�c���?r����I
u!�I���@��@�(�\;�����'�ؠDxR��d��h�f�Y&*ef${0-�ܸ�	Q�$�ѕx�D�?)1
�u@���M�?6�̱�����Pİ>��X�V~��mC�	~o���C�O0��)We�z�lI�`H�GV8k�Y�X*��V�6.c�8�6�Ӣo��'�A:TȞj(4K�3I�(�O�ᨌ�$A��O�賄���b�t�CqM��%g"�e"O�Ȋ��  � �   @�?g`0#���-�,��F�9-]!�$�*@�nUa�fX#͌�x�&�%!�D�7������1`���d <!�d4e�4�R+ʕP�1�6���)!�d�
ir�����˙&BdMS���)K�'bў�>��N�z�`4�2"�x):��A�Ic�O�"H��K�	70����CF���'rN��a*FS���؆dX�'��U�g�A&Z�x��7c�<������ �X�so�sd�)%@$i8�X��'����0����#ԉv��x�u�X�]�!򤋞y��A6J�)�P!`�C�1em!��Y���#c�_�TH��o�<�5O�����=,�Z��v�xq�"O���@V�J/��1+�>�TB!"O,�!�
π|�.� Ӓd�X���"O��ʤ뜬UT���cE�N�`I���'�1O��qBӯ(�՚XY&����ៀ�'�ɧ��N�"�
��H���w
��/��-<D��١� ?�����f�	�G�44����C^�"o� �'�R� 3��b�<�#]�����_Y��RP��Z�<9��1J.�q��"��C!z�#a�*D�|����7 9���b��40���1eg)��䓹?�ʟ������P���@&�f1���S�XG{��i�U�Ddc�T�j�D�b����*D!�D�4��JcG�..i� ��34!��D�� aAʖ�(V�K�CB�9�!�DQ� F�$�c
�5
6��S�@6O�!��V�]�����Ʋ7�I1��#!��P`a��+N
tVոC@U��O(�=ͧ�y2����%�T��v�`C�>�y�F7X�Y"E�K�$��!�n��yR�@�~.���WGK3;�X�+�l��y�jte�)PBfV(=b�8���y򩆻X�|5c���D��A�����y�/��.Y,YX��֍;��Qe��y�*V�w 4(y��I:,�`�����䓫hOq��i�ݰX��e��4M���J�"O*i��;��u8oH���T�"Od巤Q�@� vhbY1���y�*Y�� J�P�A�ZX��gX�yB����.P��$��9�d����y"�_T��qjB�9D�0�cT��1�y��Y�`
Z0�/�Xi�Ç���?a���S�q|��� q�ȴ�Ӫ �ގ&�Ԇ�+�ruӢ�_�"���D5
�C䉺)#ެ)���k��Y���fǔB�IV5P��A�Q���l�O��.�lB䉎u�2YH�H��QO��ye �r@B䉣xك�i�"������(qu(B䉃0�z�� �,n�	��\�p^�C�	*�#"'M#���\Y���$�O�����/^Ǽ����Ӹ	7� �L��'�a|R��	ejH !Ő�n�L	�Wl�=�y��S(��ժ�!�h�i����y
�lƎ<�bC��K�bQ�v��,�y�!A�CJ��%�X
lc�eI
�y���c�X���/B�܁�ؙ�yR�	(g�[g�.@��:�/\��y�-R.K�,h����<KF���y�*�Og�����-J�q�&l�y�D�(;��ȃ��Tp�!��H��y�˞%�bH(�`��`B�І��yRn�2Ud�s'�'�Xd���G�y�f��F=5�
߯/D��6Jլ�y§ 3	$v�!�G�)�,щᇇ�y�*�w:]0gG	� ��Õk���䓓0>1sJLL�v�[ �H�5Z�|JG�WC�<y��B�6PJcn�[���1�o�t�<��d�a@j]�C
H:usNHie��n�<���K{[ެАM��=x�t����g�<�@.�$�|kB�[P/�`ąN�<� n�Y��)#W��B0�Έ52��j�"O����FO��8b��D��h!U����	��:�BGm�@̘9��C��B�.-D��mL��0�b�'Z�bB䉪(pHt�C+��,��b�/q�B�I�JlhUXg#H4x�h��L�=!ĢB�	���%�C%]��e3�/	��B�IV�,H��aܖ8c$lK�ύ<BB�	zd0Д�Վwd��'�=��O ��č	^L9ka��=T�ft���	U�!���n�2,�@�ߵ;��H���u'!��ܡe���u(I� ��Qo!�3:4m"fm�̨�n�)�!�	-4��=a��s��ô$n!�� 	�<rB�@�:�\q�3+�!�D���ӀfT�j5�P�PI��[�!�dӪ ۴�"7�E�! �=�u��	�!��C�lq��A�
e*��� +�!��Ty-�A�M_f�b�c+�5"�!�䆞>h$��ʛ=��b���S�!�/ڎ�r)�&4{h�[���3��O���$
�Np0�a�@�"�E�D�!���J�P�K�zjT�JS<
!�$�Y�U� Ύ�+WĻɍ1H!�0��}`U�Y'tFRp'��-�!�$o�1�'�ەB�r��匮f
I��R�jT����3'�<t��S�eǮ4��0ղ��Ei�.P�d�0l�� t2I�ȓ�b-����	"��f*F�O.XՇȓ
n�}��C�n�D�QL�ȓ>��4�K�b'��3D$!5���V�.�� ^:O�x�Uc�:����8[n����0{DN���0mb�Ԇ�:��h� W�.�,+rH�ȓ�Rl�L�H^���E��������IC4!
�,q�Θ�	��ȓl�z`��%�S�m�Fn�#�nهȓ)����jtN|=�aUV�4u�ȓS��q��!��JP��@)ev��ȓ��h��K�����j˧=��цȓbr�e�f�C�g0 �F�P#]k�U��m)X���;QpR�xª�E�q�ȓD�M�V,�C���4m�'�bx�ȓ(�.��͐�Sd�u�I�F�*-�ȓR{�t�sa�V�����"�h��iԒ`[����h�!Jǁ�G�����G=B���,�y_������Qz����>i��LFS|���+��_��m��,��A���C�/�QG)��@����t�������`iH>'!�9��ʞ��툤�/D�H�6��*�<EH0�����UA'�-D�P1�HJ(Y$Q���D����CQD,D��B�� �`�X$��KD�w�iJ��*D�,J�#H.���J��Td�Q�s)D��"Ro��A�6kxȪ1R`&�O�����UѲ@�C�me�yhp/Z�Z�d4ړ��OD-jb��L�H��+�,%�*��"O `���&�N���B!Y�m	�"OД`�(�<z�zh�ǡ�zS�"O�1�$Ŋ&�1� V�8t"OʝJ��CJ��Ю&<�B�Z�"O�۰aw�ꔘ��	���-I"O@�
!n�4ͺ���ܘ�:M�#�'��'
ў�Oļ�)ŀ����M�S
�b��� �#sH�1�H]�w�#�9�B"OT0f��J����ܡe�""O���7	�� �  ��)��q"O��׃@55�QǮ��Y��Y8�"O|-C���";Ă�����R���'���ߡ��9����,J/N5���7]�|��)�d�T���8�	_�1�ޓ�y"㑼^.@pB��L���� #����'9ў�Oufm���\�͋��UU��
�'TJU0��ޒ{����.��U#X��
�'{:�� BC�!��KS
?v2�
�'ܤ����g��� 4X�/{�� 
�'k4\���1�x�dAǶ[���Í�'0ax���d2��x��I�Z�#H��yB,�P�P�ޜEX���a*Ѫ���hOq����w��i!p�YÖm[�"O��2Ĕ*���0q!���8
�"O|}���*{G��Q�{�xY�2"O@�	�@�<\`*0H��k���H�"O�	Ѓ*
���RAG�[��md�'�ў"~�1EƼ}��є$�#9�z�yG�	���=يy��.<C�D�k
�C���2tό2�y�X�*�ȥMT�)�6��>�y��Ģe�>Չ�& !��,x�����y��9L�J�� �Y1����y�(�����F�X=JB�A5�y��*[�!��y$�����?����S�v{ٻ�f�)Wa$�A@[�j@2�ȓH�������<��	��M�.�=��W�l��Bb�7�V��I�*x촄� �2\��枎8_b�����L����ȓ#��49���?�`��\Y�^ԇ�.1�0� �T+�2%�0`�T���	��)�a��͜P�A�X��8�?��.\�y��K�0�q�ë�o"  �ȓrR��c�� 9�HP%�`e���rz��1#DVzt�!ůs��Y�ȓ���jS`�i �`$)���F��+�\�#bK�(R@h��F)�X�ȓt�H��9&Ʃc4G��cptȆ�|y�Ԛ�L�8'h�SӅK%%`
y$���'��>��4:�N)Z�����c�O<��B�ɌY&ب���� �.��-F�B���x�r�`�+���:�lZ2hfB�	�,	�l;� _!=��`3e��U�C��:Ԯ���M�Pv�D�fA��ftC��<2�b=S�7����a �~\C��^a�����܂��[B�a{ C�I�od���"�!xt����H�HB䉵<��mIsg%+X�v�m(� D{J?���	��S�:\�U.MX,���H D��QFL�6Up�i7�xX�=�5�1D��ca�U6E!��aپ��A1D�@���y(���0%( ��q5�0D�P�Si�>Q2�j֋UlxQ��d�<�H>�
�'L��h��P�[Ȁ��Օkv�A��x�N�Q�o�Ojv!ڠ*�_N�?���~:d։%l�`��+T�"�ӥ��d�<�s$L�L�h�'�&aT� i�^�<)��M�#����gG�Ei`X�D�N�<)�nG'f�(� Cl��[%\r�'�@�<YR%���C��:���A5F�ПhE{��IY1K!��X��"em4����H��8B�I�N���AE��u�8��%�G}6^�HE{J?� ñk�<S6h`�GFd�1�"O�С�lL?U���b!�&W3�@�D"O6!�w�є^�4�Bd�W l�I�"O��5�K�%�T�$�ڷD��b�"O�����R�a���_2G�^5��$�OF����-�=*5��*J�`ҡi�=r�b0O�EY��х9��ě2ٜ9�`��"O��jj�	2f�;bwD�B�"O�,q��
?�8mP K/Xh��1"O`�Zf�D��ur��4FI0��C"OzH��'m�P���P�YLxh�"O�$볈J�~�v\7h�.,�͑f�|�Im~�e
�`��T�c �8�xU�p����xB��V�zh�B�SV��훳 N�7I!�d(J����!Z�c�t%.d����"O8��@S�p0�Q��H�Q���"O�x3qH�55=\�S�m�4�|]��"Ou�$ͯ��eyb�d�l�1"O&�4�		1�~}�NN��\6�'w�'!�)�L~'��0��ɥ�@�
&�	� F��y"�ߧIIZ���0f� aˆ�y�����Q�S)(萣�;�y�+ЍG�*-q�l�R�XM���M��yb��:T
5�$�C�0������y�)֔P���e'G�,�Ѷ�W�y�V;�h��7D+`�|����D,�O�Y��fQ5<ײ,s&%ОO�V$�0"O�0�_�g��\��M<h��`�"O.��D�,�l��"J@���$��|2��5h6az�CPԆ��Aa�]�9����y�E��`q`�Yi�)�D��Q$��y���9I^��r��3�Hz� X<�y�*�>-���E��9�>���Ɲ��y�E~}�Cě�3�.C F��yN��.^b��}D^Pq����y"�\&(mQ��1w<uI/��?����D�<a����5e�Ԩ��-�PSE��!�T({��b�̻~��ј�,��!򄛑F�9t-�##MT����!��K��er�(��a�б�rO[�e�!��-)XP�0��E)�ʍ�r.�<C!��
	Z=�� ޠA5��hӔ^���M��4���̰>A�����"�,�P/#D���G �Y�c������ #D�8��`�&>-����e̮>�p��$D�,a��(���y��ԣ$�D��&%D�@{�F@2Bh}	�n�3�M�QE=D�h��J�?p8������ "�%H'�?4� �2oI:o���h��'H~٪���H�'ya|��ߊ&wf��Ӂ�$q���Co��y�g��R��H� @��i���*��3�y���sfz� ���a����(C �y�%6g����Oٖ[ ԼRbJܦ�ybM���B�jG���V+�I�Q��yR�߮+�,�"L�G��:��Ż�yRkOi��0���̀Ft��i��+�y�̓�%+ڬ
����f�iY7H��yRnKd� �3F��¡�f.���y��h�.]��u3p=�jψ�y"��E�%s�L�n'�!+�
�yr	�8��܃!�	:��p&��y�j��-n�����V�8z�x�	�y�_L*��҈�5�@�Z���1��$%�O��d�-8�Ĭ8&�6"U��9�"O� dDzI|�|h��\	5���b�"O(QI��!&�e�FG�7f�<rb"O��C.�%3z� �GJ{�=�""O��+����_�ZV�]$U̸�p��S>���A�; 8�a�G9�d�G�5�O��uP8��`¯>�j@�SiH.W��D+�������9L��U��"�6�a�8D��r��0����w��U�t�"��4D��6��.��Y�c�B���$ D��:�ڲPM�؊`c	
,ތ�uh8D��aө�#9Y�4l��]��)�Aj�<���#}*�(�(\�w숵0w�^h�<��U��} �ϝ>2F���f�IX���OҐ�`�E�b<��'$'9fm����dЬ'?�u���H��>��'V�^>�IJ��\�'%W)x��&ޠV�@`�J2D� y@,ʄ(�PbdJ�ޤ}�A�+D�X{욇37�t���_H�\PGf>D�����W� ��ز���;cƸW�8D�L"S͆-[: "�J�Z����7B�OT�=E�dC��'�$�U)�kj(�Lg�!��"gҜH���̆&Wb�
H�*�!��:Zn�I��O$%�\���� �!�DV:wJn9ڰ0 ��$b@�~�!�D	�'Z��a�ă%Ŏر���pzўL���+q�6h	���A��+�H,ZO�B�	�\Ppəu��7p��e�:R����$�S�O��`��N�<JƸ�!E�M�7�C��Wl�x��l�@�j4	��{���ȓc��1��Ȁ�!�Zy��*�;>��ȓXġ#���l*%J��j�����^~�s�@��y��m��-N6L���ȓ`���cI8\0��p�Ҷ%L*��ȓ2��`͝ 0u��:F�I�&Z4E{2�'�$z$H�1J"@�jE7)t$�����y�C�gH��OE�|X
R����D3�Ov��
ܡq��K�/V�e86"Ot1���ЎW-0�0W�WI�lB�"O�хJ�/.��6G�&b6`���IE>)��3@T\RA�ֳs�l����3D�0K�%ʍW�8W�S�q{�$	�
�<���Ӣ�^�#����5���h.B��D0?���؏x��\�%�7d�v08�kRAy��'�����2dI�&�١+#:1 	�'����)���͠v�L�o��!��'3VhxC*�m+��;eoʋZ����
�'1r���n��eQe\�=%V��
�'j��Y�T�;�p�PR!��O�%����hO?�p�.��V�rVJ�
�}�a�Hx�<I�̌A���Ǌ ��`ht&i�<���.m&�a��+��/�%ȷ��d�<1�(�
5"2�P���QCRd�2�K�<��ήr~h�"�T�]���#KI�<95��b;��C"��Z���І��]�<��B5c�N�хi.�\�e�@y�)�'M989���K�p�j�R&EXC4�ɇȓhfh�gg����ӈ>����_x�<9��ͷ+�V8�CL`�~ YŎ�u�<Ѱ*o��Qr+'|�<�`��BX�<�%�()d�&.81Zd��H�J�<Y��5]�D1KF2v�()B�L�<�	�*�5�a�	��9d[J�<!���
�	+�.��L�0��HyB�'��c��x�0)�@=�(���� |a*BO݆�\��ր541�"O�8�gL�	�����.����"O�c�� -�V�QɄ�.����R�'T�	n�)�=qBΆ�?ST �񄁟��*�	�l�<�P�\��`�A�8��H3�g�<�Q-O�d�>����ـ 0h����b�	I��`P	�x|M�n��!�tp	$D���4E �b;�=愁�;&�K��"D�8+& %r(X�_�B��SaE6D��
��X�d��v+�gG��P�A�<��2��m�Ba?8jh@ C�KL�|ՇȓS�j��g퓃f'*��؏n��݅�i�`�6",(��˧hY��r)&�0�'��>��*V	�!��B^�^�е0�k �e*2B�I 6�Y�� �̮i�d����yBȌ�d�B�&�dT�@Y����y"��ow��mG�X$��;�G���>a�O� Di�=zԠ,c�ȅ�^:��[ "Opܰ7-�7�����b�h�%ZG�|r�'�az"� �Ӡ$���(4І`_+�䓑?��D1?A�f�D�16bPcy e�wM^�<���Z+�� ��?i���@�`�<�eo6u }B�"�����@�OV�<��/�vb��Yr"Q<b�HŰ" Sx���'�dK�P�8 ӆ��$ڨ]1���hO?�	�.���P�S�W�h4�}�bdU\�'�ax��ޜ\��x�M!-�t(��ǜ�䓉��3�SJP���Oʠ�JW G
1)�b�<!o��4{���M�M�^�q�[g�<�A䜬1�)�ɓGݠ%H2( J�<1�/F�
�p���ʔz�(У�͆D��x�<�S���@	��"]�uk�˟p��[�S�4�'��	A$��$�T�K����CY�1�LB�Ʌq�8�����~���e���L�B䉅%��@y�k G��Z��<\�C�ɪfÆ]QT�&<?��s/ӫahC�Q�v�;�e.V����!�mVC�I�qcl��@���C��1�N�'(cLC��7��`�H�8}�W�̲C�ɏq�xИ��ԁR� Ŋ�x���2�S�O<����ތf���ZW蚶gq�d"OV=�U�V ����Z�nWU��"OD��:��yq�KE�8�H��"OB�(�cB
FJH�3%��o��T�S�'��Ez�٢F��ly�:�jY	a�L<��'H~ɩ��I L�h��dĒ�^�-(�'����	��7=YYtcί |dK+O����S�L�@�����P��OC��P �h*D� -��OUd�YUN)3.�ܹEm#D��%�]�m p���*@�.m��.D�0+vN�)���ˇ�4h��P��84��	�>Xr�ҐG
�Z.�t�Y�<�"��:X16H�ON�_������K�u���O�\"ыD�YI���C��b]	�'��"�N�K�R|�Th���8X��d(ړ�y�NY'_�"]����q�h�8�h0�y"J�+e���:� J~dp���ֲ�yB"۶"��HA� �p� �"����>�)Ozd��G��e�-�ʖ��C�=D���!J]
tT�T`��att�" �ON��!�)�'	�R�`q���t�T
E���Ѐ�'k"Y��o�$���)�l����$%��.���k�X	J&"p[��Z�O|�<�炂�56�����ڜZK��Y�B
u�<� ���	�&l�2YB�U\�2�"O���cD�2)i6����&gJԨ"O6|�F�x���P�M-N�6C�"O2����
���⠁�bp�X�6"O�DȤg���Ȋ���;G`��7�|��)�ӄ'�PU�ˍmd��˷�H>�(B��,yθ�ɖ C�L���ʀG�/R�B��7�Z,�� ]!�켺�H0��C�I�	�Rp��NT�|�h	c�:]r�C�I%\��y�"~�8�@�dv��B�ɡ_ hA4��`�J��QHS��B�ɶIT��/�o�>5� B v�<B�	�Hd��l��mx8�IF@´B�,k4���� (=�T��,Q�0C�	�AB���T┦#$4,2�nY8#�0C�I�_�}��"Z$7"�ZtN�e�C�I.8;�k�)L�)�K �n��C�ɅLX���7�[�G�|y��ž|�!�䙴z���2o��߶��vD_�m!�M�;��(Q�/:���_ �!�Dֻ�R���
[ͼ%R����!��ȓY	20��@>0^"���,�#F�!�ײ�x�B�8cpvh�lTG�!�D � �"f�~*��j�!�d@�`��BT�З#FP�2)�(�!���MP�����LKx�`��!�!�NJ�0����$�n�i#���`!�X�<9�h$�˶��R�˚��!�ĕ��45RI�Gޢ`q�
�&�!�$�X�8ڒo`+��*
9B�!�H�o��
�eC3(��HY��!��������+^*�!2���-s!�Dډu�Q1���4%K�N��!��u丼�$�ؐo�h��C�xm!򤈪N�j쫇��2~>�j�@�8�!�ό~~%��ס-f�e�P%�=@�!�d�(S/���T�XIv։�q	p�!�PA���5�,V^�-�d(�.Z�!��G��P�t�L�JK�5H�5<�!���d�w�}W�TA�aX
u�!��,���
�#F/g@�Q:6�_G!�$W��"��A-��s���;G�!�*���(7熃,r�<QnR:�!�WY�����N�8h|\գ7�>YG!��	Ħ��@�[���+���Y!�$��!
`4RS!��[B�����X�!��u,��jǽM���"f팅#�!�d	^6�<�a�@�`�;s�(+�!��
+Μ�"�_-8V����	�(�!�$C7*XZ�e��-	p	�эݡk|!�$��@��j
�,;0-Jti!�M�x���փ$|���=|!�dB�4�t�@)�He��&Z�6�!��֭\hT�%���Y�-Q�nʩ5�!�$ϳ]
�Z�з�.���U�!�D�;ef�����$8d J05+!�D�+��}1� �'II��CB�o�!�D��<٪ �E� 2\H��n�iD!�d@3��I�^j�]"���Z@!�`3�H#0�؎�̢�FK
yhB�I�&e��
�.�H��K�ƅt�~B��C�f�G,q�à
DX[�B�,8{*P�R$��M0�e�r+xB�	�z�$�A�K�F�}��e['EVB�)� N���H�:��h������"O��)�-���6�Hg��	n��T�P"O�9A�HN
�u3��ݬD¤	b""OTA�@��-hb:���K�X����B"O��qG��:�R�h��b��	�R"O0�`C�؛*��1�8V�,�W"O<\� d����B$��zF��a�"O�]�f��S�l�9�A-Hu95"O��褢�.�(���F�Li�"OBura']4���=��M��"O�f,X�6�Blr��P�G�|-��"O lYW��4� ��|Ժ�ѧ"O4����o62�Sd���M t"O�5����5�@�)qi���~|�D"OL}A�n�EHƅ2E�F.*��u�"O8$�Ƥ�-���ɶg5C� ��"O$�82'�.L x@iB ��Q�"O���g���BUʂ(ƅ_����"O��RKe�`乲�Lgj��z�"ON�����2X��+�	E<Upp�"O�q��`��}�tW�qq�ѹ"O&I{����_��-��G͠jEb�	�"O����I!~�1w�V
�"P"O����,�5�Fn�]E"O��q��>i�*�X�o:]:n�K�"O���2�ڤ+�}y�i�*R�*�"O�� P��e�(�JG4�@=��"O�S��̰ Fh*R'^<E���E"O�}�ǯ�}�fb&a� ���2"O$�9�kR�0�Z��Q�_M�X�@U"O�4��/7GT=����`}(�c�"O�(��o�A��M%KӶ�y�"O��'�� ���Gɱ%s���"O½ࢊB�/�`F^�I�.�!�"O:���AڢP 9:�NC/6���@c"O�0�ͅ�-��(	�-�U%��1�"O���5.�H1�����QD"O ��EK?=�&Uj#�G|���Sa"O�� $8E̪����4�9�"O8�)u㊕y��ࣰ�I��.�D"O8]@�݌Oa�ͪ���A�>�K�"O*����L�?��1&K�q���`�"OR�@�Ӳ+�0)`s]�!�"O*؃֚S�U���?I�$�s%"O���7 D)9"�|زe��|�&ك"O��bC$T.XQ ��&d���}�6"O��b�e�2wn~lxg"5z�t�h�"OIs��A(%��Q5�N3o��c"OX�AS���r�lXC�NX&H6"OF0D��-�����O����T"O@���a�lo&(�����x��&"O6h�H;���tm�R����"O�Ɇ(ӳ>���DmUf�~���"O��FC݆L�ݘՉ�K:(��"O*�3��H�*j�Z�Iӿq�D��"O�4�5�ʖ\.*I)p�ٰ��L�"OL�їG�F;�Z���\8��"Oԁ����$�<��HF!t�1W"O�1�"R eR8���۠I4���"OB)��ʨ[�0��Nߞn���qP"Oα#��
|���3�-ܢa�XrP"O¼��kP,�-��ٖ!h�BR"Odts!�R���,Ʌ�� ��i""Ot���>j�^���U��)��"O� ��hǄG�`	⣣��Q\�{@"OT��K:����@�ĳ/C��"5"O:��i��"ul�ː��+p B�"O0���K���1Unȭ4i��"O�K&&��+���آ8 -��Xs"O(����A
9{Z�B�@�r yI�"Oh�[�Z[Bp!a(�?C-4!�"OzI�!��8��+3.˱:�H�S`"O"-	��.�* ��N�n�2�"O��E��?��T�SȀ�,�`"O��qCg�-���`�F�VL�"O0ui`�T��d�J���+�☰"O|�	E��"H�:P��'
?k��9��"O0��! �,bx���f�>�9�P"O��:sOQ���$V"s�D�"O�)*�$_�2 $yQC.����"O�	�v)؆r6��C�R�u�X��"O^��S�β%p�:Go
)$w�s!"OF����:@��1�R��]ї"O*7�8(l���En֋oΝ &�#D�4��gΨH��� �T%>< �Y��#D�8a&F�7d�D�4+��'���5�4D���#*�#qo���H�3@��x�3D�̹�)7<�`,�h64�|aiw�1D���I� %���ĤslAS��/D�\��(̄I��I#�n�wN����-D�4	���c'�#aFB�f�$���,D��Qr�M)�F�7f߸$;�X��+D��GJ�"%ZDx�E$��rA�Љ�e(D���SF�D".ɰ�D�l܊5��� D��O>,�ƝXC��:�x���*D��pCLS�hz%��I�mV<ͣE�<D������	��b�/�4}��<D��37ɂ�HT�� T:��%���8D����׍Y\�m��hΚ8��9P%h8D��s�(��A��p��Acg6D�d��
�����5&��5
:D���w�͙��I�a	��t�U�E�;D��@ԫ->���7'�qb�IZ�%'D��CǏھ!�(i��ɢ/�}:/&D�\��ꕝI_(�*�j��#@VB䉏D���rFK�$��90ϔ�+�B�	�J���� `�	'P�4j��H�C�I%K~��F��:d��G�Y3�B�	'X���m*A��j�|C�I�#q$UZb�W�}&�1	�&��<ZC�	�ob2Px�خv�5���E`�C�I�E.p�yV��&_h��Y��B��4C�I�@�j��\�FN���_�r3C�I�ަ��7�Zl�t�Ŝ1F��B�	�\X6|`��N$Z�dز ��K�B�.h�4:��Z�{�zl�E�[���B�V졻�O 4�HT�b��N��B䉔�@0����7M�:t�w�V�MڄB䉬��f!�Be�?y)L�Aq*O�͚O�!�qisD|���"O��Pa�Q�����U.ظj�A��"O� �� �/EҰ�%C߄J�!�!"OJ��(ٕSR�5ءaF��h�"OVY�b�ϡ}�n���@�$��(�"O�%�Ң��\��p�!7Q�<��r"Ot�h�ܥA�H���;q �8�D"Ohĩ$"�3��!�C����'�qO��/C&"�X�rI��1��A("O�  �(���m����2���`��'�L��'�b�٥(�A�����C5�=Y�'�9�5O.���H�9�|*��d'�S�Dʓ�]\&d����A��h���y�#S��9�TZp�� �T�/q�<���O�(�-Oe������n�H���I ����!�[3Q9�Ţ0�׌�b��Y�hc
�1�2�4��=[��2@�)+y����Ñ��'}}�'|��#H$T]��S����z���H�'�&-�\��؋&q�Ɓ��OTY��O(�	j�Ӻ;�O��36+�3I�h�b戅�3_l�[�'��U�s���hy�!x2œ!F������'�ґ|"P����ʑ!G0|�D
U�SaRh�cVh�<���E3'�$){��&~��x�b�Za�<� �&�,����׼cK\Ը��Z[�<��Ƃj7�T2���yl� �,�Y�<i�E¥BP��Q��8I����eY�<)"�ҰV�2u���\</�B���S�<aL�%����9i��;ui�P�<�f�dl�Q�v�̭8�:a�$!�$�	O�$aA���T����)��k�!�DK`I� o]�h�V�2!�!��˲=�R��Gtԅ�s�\�j/D8��hO?M��9N�$�H�BѧMڢ��U�#D�p	�Ƕj�� �φk��$�!b7D�D
�gH-�y$���G2����*D��e$Եv0V���@C�sh�ʷI)D��Ĥ[�3��(�fj�L�d$�s%%D�p�  ��sž���6M�b�r��5D�H�s�*�`*��b  �))4D��ҐD؟+|���ߞ=�
 Ò�p�E{�����pB� E�:�Ą%-!�D}���c�ϥ9��y��IݪW!��(h��d�3�&��&��N!�d�6jB>�$�&j���0���n�!���g
�51���,�rf��X�!� ���ۦ�L(x(ٛ �ΏC�!�Ԕ|�i�筇h�����,^�	s��0<�I_ʺ1Pd%	�@
��$k�<�% �/\ph�3G�H�U�0R�e
릑���/�T�d�J��N�Ť=cBiF#C�ZP��6�q��VP��G&էg�D�'��~�#w��IF��^~�p��Y��d5�S�O,�A�BG n�&��B�L�a��Ep�'��+�ߓ<6�|	����T5����>Y��	��t|p��PdY>Ti�V*�	F�!�&�>,��gڟ�Kѣ:��p�ݴ���1���O�@A#��a� !��Ȋ2�nM�'F$ы���1�����gH-0A�xS�'�д��	
��uA�`ԛ'�LJN>����~��tR	�0,U(H����ȕ�y;<\�� �K�j����RKD��R��<a�O�ܣϓp��@gٖ���9��$Yݴ��=t��ifjݝ_"�-H�	�yr�Gx"�'���X���1���ׂ!H��4���d>��UeC-Iش8O^3	�(�0Pa6}b�'SP�zg��G���ж�M�C�f�9��?	��:1�ѡp��5ͺ�Q�g��k�!�_�z���j�$�@`�4p6�N�+�ٟ�'��;�Oq�
$z�H�]��dCr$P�M��=A�"O����♎>��<k&�0,��,;"��3LO��x�
�+I}H�Sdl�(%l�q��"OL�l@�Q�dЧ�U�`ܩ�g]���I�G��ʁ���fL(�Jː*��C�)� vh���ùl�����Yk��	tX��Y��[7D(�(&m-YV8��.��1�O�� -a��� qo�; V)0! $�\�f�E�^��p��Q�H�Kc&�z��D�?�e$څ|^x�K#��2�4ъ��L�<�#�U;]l��@E�,Z�D4Z��dΓ�M�O>E���d���B��H�&�2���J��'�H��?�͟��J8jYP�dj2
M��֞~���'��&�'���3k�u�q
�͉���a��>�e*�>�N|n�?'v�,Sp�)!�U�ƍ��l����ēMj�H���؀"N@@(�nLE���Ml��u�=q��T?��r��.�
|�&g�g7�A�:�c6�I��P�p�圜`��xT����84�x��)�S�9�ؙb���-�`���	��b@>O���۴�ا�O���t��0e�`�+�23+�y�O����5**PK����Z8�D~�Gx2-�'�?��w���d�ЀII�58�Bʇ:��ȓ�6�8����+�@D���T�����p��>	��3�f�r��AM�Q9D$����
���ȓj�Z�q3�
�;fE�p��_	�@��O���G�*�(Hb�/Z��O��@u�u!(�21��/����Pe3D�L�� ʗs��yu	��P"��#0D����P��8p`j��a��� /D�dY���Zc��` �]&t���XAM+��6�SܧVJq13��};�B��5A\Xԇ�A�&	��d
��J�ふ�(�Gzr��d�O-��i"���x��2�@83�4��'2F1÷Q�h�x��B�G��4ճ
�':*��'��,}z�;�A]�t�މ�	�'��U�T-S�$�z��T�6Mq��'�p��K;3�Vp�қ@�^5��'����%�ʢb*�<�D�)@�f�8�'ˮ��D��i�z923 �iD�Q�O���$߉j�X���l��&�.�Ԡ,�y$��asCnJ57��Yc!��~R�)�'n:T�b�J"�� S�ɫb�BL��ID�k����D�Eh	�eXe�$(\(�ȓF���c�<A7X��`�Y�"�����hO���`I�/ԨxS��������T��DR���'�(��`�پJ��5#�;6 8��'� �C�Tٜ}:E�92.`x�'�*��1ڬW߆0����[�s�'��,	�)��p�왻������0>�N>!WG!�H�3��	W�F�zg��<�'�Ă�-��؆C�8��S�Oq}g?��(�9$P�-4��R�S/0�����"OP����L�o�D�������'��<�	�O�8{��H�cG���Fįw���/LO"�`�ׄJ�[����&�@px�� ��>1��-�b��$'��3��C�&T�J����8b�H���$(=��ښm�TXb"O���QMX)?�`�6nC�U�ݐ���d�ڃ��D�$@q�%Ŏ8`�Ҍ�S�<�6`�F�8A�_�$H�-�t��<Q���6{�Ѣ��
2R~xx6NO'��c��D{����P"a<8���?�$������y¯�+a�� V���r�|�"&���y��/qGF��'X:w���!gk�%�y҂�q~���T�E^F8;�N[�yr  ���3�IF�T��X٦ ���y�!H��#*�Gk�A��V�yr+45P��"@L�.D201)5g��y�̖�r��a����>%"T(J�7�y
� ���#�uZT�ħߡQ�����"Ox]9�D��b�C�ĝ-F���""O�Ȉ�,���1���N4Xa6"O���dl?��(d�9�1H!"Ot�S�Q�:��eH1�P�U���"O��y!(A�4����0�-\�r��"O�����k��P��B��zG"O^�S KF�Uw��KDIQ�?� Y"O���G0�[Ղ^��ڰp1"O:��ЯJ�j�`�Ȅ� :��՛�"O2e*@�B�\ܰK<�fl�S"O�]��!W�/�0��-ʭ0��<�"OACU�^m�Hs$���1���"O���U
Ĳ+H$A!�ю� "O�e�"���DIpӬ��VÎ��u"O�]��'�:F�nX)�+P�nI�"O$r���j��݊�)|����"O����:��H�$�)cy� '"O�b��E/4%̽�6I5p
�"O���Dbϧtd\*���5@���"OB�K���?A4ؐtȮh*�At"O�$��˩Gz&�j���v� "O.%ఊ��l�\���j!�i'"O
�§�˘24v,�hF�r�us�"OD`�
�z�`�f�C�~�xV"O���'f�.�0hӲ�&O����"O��6���e� R�-=��B0�J�<��
H:`�h�@�pN���G�MC�<��@N�?C�$�I� 3Zt�v�XZ�<�#D�>?~��*�o�1��bX̓`��s��;M
���=w�t�<)U�S "B���^�xTx�Z
Q�<����G���-�#
U���T��O�<Qテ&ݺ�`��5����f�@�<a����Ҍ��Ѵvʍ���@�<� ��&�{Ӈ� <�āp�<���Y�B5���׳*V�e�3-�v�<�v���p攕P�Ƃ�wvL�ѩ�K�<13 �/m"&P��NZn�! fN�<id���Ԥ�>p6�Q�VR�<A��9 �:��\�2�����K�R�<�t�Z� �����y�6u�4�QM�<�C��T��K��K���{S%�f�<�d��P�R���Ki081[P�Vg�<��E(\��}�D��tJ<3���D�<����$$ �X�B��r �A�<��N$(��SpC�P�� �`�Yj�<�
ߣ(Y�@��@�
�y�g@e�<A���VTllá���r�J�a�+�a�<�剓>;W����Ȟq�l@��"D��3����$�3��pVp���!'D��3`ڕN��r��Ȉ	�Ppq �%D��W"Ҭ	�n<����TB�r��%D�Hy�o��#ΚQbpmF��v��M/D��"�%K!Q�TZCÙl�^ҁ�0D���Ug�m��� A+{B"�.D���Ɠ	2m���9o~	�I/D��F�V�H	���� 	Ap;F�-D�$��+D�g1|�q����&�[��*D��������Ul�#m7ܬ!��*D�[TQ/X����.߳2��J��(D����혋u�8ys4�V��`�A2D�0$b��+]�a��h�H��ԛC�0D����(=7�yc���7IJL��0D��`��w#�1�u��.P��D�,D�� ����C�%8tY����L^�iv"O��C��Q���� ��_�`�( "O�)٤�&S:�q�`�4	���"OR䠳�!�Ψ*D�*���H°iv0#�'��	rC_�cd�rǋ�\�Lu�(���2a7?�s,[�xAXݑ�GК~Dp�+��Vz�<�!!Ö9:�<��	v �+��X�
��9�c,��A&�M5.��TrA�;u�=�"O�TQ��]H3��b�!�I�"81�䈗V�qO��#��Y���DNݫ}��"�$�)ۨah�M2D��ۆ�M8l�fbt�+l^�X�>lȨ��6�O���*� __�D3SiR�m���'��H�da�A~��G�<z�Z��O�tP�'�Q���x��-��!��l��	��a+�+f��Z�x�FV�cU�O�On��b,I.A0v�v�T�# �9#
˓]�n�S�.���|"�  !(�b�P��R��'!�$]-���@n��1�a�F��%���VhZ�[6qO�����"GƷp�`<J��m�PE�V"O�(�b��Ey��FI;d�%"�,�	��-)��L<�Q�H5>��k֮�$�f4(7��vH<9"-?ԨhI��M,Uba��E�9ɖ܃0�*�O>��d�_U�`	���R$���Q�'�D�*�K�M�I �j��aD<1U!�$�!XhDC�	�2�\u`a̞��l��
�&��O�`��J?�)�(R\�6��[�M����P+B�	6Zժ�L��A򋝷V�B�I�^�F�ߺh���5↔r��C�I����b�S��";}�C�7s!L咒(d���N�(�C�IKe0�KV��0c8t8׃�G��C�	8��{@A�� ��@���C�5kh�Iq�
6�8Y�	,A�JC�bX�{'D��q��ATIG�#-.C��ol:8P&l�j����BB�I�n����ٱ��	��ЂS.bB�7�P\[�J�1y��ce �׊C�	�H�]0�Q�9!H1�Ԃ�Yo`C�	�.�o�;FR\mKB��e)RC�	<�h�aԈ̕e�\�8dmA�(C�	�7�\̺r��t>���� ��B�I�9a���ҥѤ|�{b�"'�B�IC�b1�FG�-OX�������4�⣓�5��?M{a�`y�,�7��5�|]��"D�Db�(����Fه"x��`_��ؠ0�|rO?�g}2g+4J�D��?K񌽠'�,�y�]�)��񨧭YA��L�fD�ڽ���yܐm ��N��0=ɳM.^��e�Ee�"~}�|�0�Fpy�-��T�����|ZwV^5�wO�`��ͮ5�4�i���+ ����'�҃0�P�'��t(�"E�k��+�/��h�!���01V ��%����X��T�8'�b�qq�]�<&�=A<��v��S�	��/F�9/a|Х|3�Q!'^�_Z�)�E�]{
	ӧ�Z�t��Ј �T&UP��2~_��a��JXT��e�~�B�x"E9z�r�3gۿeI2�6��э,��ں��<I3ޱ�'�^�&��i���	�@�	?q�&iʠ$S�R2TԠ`-F�s7�$@*�K����<)��3c�D�%/ "D2���	�0��%&n�5[�*1B�d�Z����3a�l��/�!&N&�ɵi5��%s�?����u�ˢS8V�(�*��u|R��Y��(2�7u
��T,��t�D�Zӫ�u�RLXs� /L��1��E�6���׈�4r��,͐r�L�3ًs�@\`s� /q���2��G���4bU��#x����D�~��@N�|�BE����JJ,���jg��qPR���v�m��D�;��0��"H\r'Ϛ&KL.����	�g����ٓ�I�a�ҹ�N�*V���8$FX%�c��9&�:n��zg9�L����?E�D�Q�e{HQ���_�,�#�$\2�y#6g��:ޕ�%o�?F�|�UcX�cw\M��A^� �sԛxr�'��lذ%�"k�n��&�J�Z J@2 �]�1���:k�<��'��L�e� h�j��<+�n�1��Af ��VH��Ni�b�	Yol�(4��o���)�$ΐ��,3L�"ׁg��,�PC[�_���2��)ql0&H	�7�����*,1B�B�A�g��,l6� |��FQ
>ԙ�'�Qf�P�=]�6y��]x��@R�^�^�:m����؀ �	Sd>�6	�B%B�h�|t�B ��1D���h2-^0doZ�[蓦ɾ5z}
&�
�o�\��0� �?qX#V;M
R�4.
	p1�� ��!�r��fl�Ojf�j�'��nEr���n_>GAP�I���)ts���D�y�ըH+0/2�
�n� ���.?DF^��'1.h
�m	2*�W,�/.�LM���Q��0�B����铄5$|"�k�W.*Xh�#�!_d�5	W��	���Ae�1*)���]�s ���o���k� �6��j���%���'�Zh���]��)�'�)�^�n�;,�=nG��AS�V3{]���G�-��	�d��k�(a��pE����i�&}��含mV��OI/|�d�4F2a�� B�0}r	��f�Ʊ[�D�}����o��1�8�P��vܬE0wBΩ��yK1�	�5(4�����rڤM�~J�G[�X�`0
��S�G;�Z4�̌@p���%� G�.�P�C� D����Ox����<���&��ƍ�9�z	�Ѩ��[�������+ݹB�:&`[*t嘨��g�-U�ԍC� ��f	��"���-��J��'�X��w�@-V}�%��5ΆP�'`%(p
ʌ/%��Y�>Ap�T�XZD1LI�P�H���L��\1��y�G���(��2k�I�b���5���E�S��~	���Qي��c��1���A��ӱ��bL-a�¥f9f�R�9~��>`�gّtVdk7H?7*�x*��/ʓS��80g'X�|Zt{���o	n�r�@#@�}��,��G�"��L��.�
0
t�WoO�z�D�𙟜��F_�xE3Ŝ�ed��"�)h�=Y�n��PWƑP.O?��Ӓ=�1{�!K�?Ḅ�gMZ:)a�#_��8�s��}�d�5��U0@��a�C��6 ��)�J�>���X�\� �l!�	�]�(���9T��z��0az�pV�H5X�|�`g�-��(3�'W�Y�b��3b���a϶~/5�U�Z$6�����V�zt`����8�� ��׭dl�ȰgG�|��&��p�N��T���x�@A$Vu�<YW�-F��IP�I���@
u�j��R0e�,AQ)xO�pl�����y���Z�:��+�(�DA�����y".�Sa,���
�UG�������j䜰	e&+R��`h���a�Ƀ��T��E��f.����&�?h�bxc�6A��~�2K��pA���q�"R��X6�,�B+�u�<r�UZ
a{�<20&Yڔ-�+h���ܩ��O♡ai��n�B@����x�ZIZa��������
�$�g:H)�"O�=��(�"��s��nz� Z�<��bL�2�Y��`�mCr1����G=ꌺ`�B$*L,���C7JrB��*@*z�(�a&��UJ��@=0�b ��A�.O����Y��xgOٽ:�,؛a��� �:�Z��%D���$M
��s��?��0� a�qՔm�@�=����,`�vKƶjWh!��Ľq:���C�4���@lڗH̙���ne�<uK&eJjB��/$�2��& \�̌L��M��-Lc�h��K�G����@���4x���_5���A!�z��C�I%^ <d�͌7
�Ip g�%+�R]�%��&k�ΒOP�}�j<�c�lΩ�8`A�DN:oq@����Li�f�U.,*�q��;G�*�ȓ"�(@�@)-�̵H�FF2|jnu�ȓ � qU�
M��w�W� ����ȓ���Z`�zAZ,���1>�\��O�T qO,�}��l���*cx^��]�TI>�ȓx�%9��8�J�#�O�<+��n�%�
`�B�i8�P��D�a���-��A	��25b6\O�ac���}�F���'��b���1$�������Y8���'A��9��_�x�噲��َ�!�{"LɀhM�8J�MA�O� �`��;Uz�2 *�� �'�����Jҷ)]�F�ζ!����e8�*i�J�����<P��̆KT%^,B� ���i�<��NI�kw,�8򌒠c?~�  j�X�'S�&�"��(��(�&�ްDA0� `V���A�RM�Z �E��y���in�9`�W?R~��0��N��yU�?�.J��L-��K����'����Ņ<�b�E���!���(�/�F�Z-�pjS6�y2� K�n}�a�Ō0Qh�{Gǉ�rL��OV7���b�Q>�|�����b����;Q��хȓ~�����kd�P��1'�Z�mZ�bҚ�K�!�L8��b%�\�i� i�BJߎ�S ,|O"�ԭ������=ZsV��`�ζJ�	��}k!�d�5^1��Ǉ�q�M� *K"o!�� �8"��U+�RQ��r�n�3"O��� �5�TXJ%�M.0�8bC"O&�A3e�S^J	*�͕�-���S"O��FG�|�3%0�*�ѥ"O6� �j�!�`�wn��@�@"O0�z�o�;�] ��� i����"OJ�X�lO�/J8T��� ��L�T"O�dK`(^K�t}��Ͼ4��,��"O�Q��S�Fs��9��5�V�а"OT	�����ĈF��0�d�"O:U��_Nj-���y�4���"O&���N�M��V䍐C��-j�"O��JW�Gk2�9FYAR6��S"O*D��5p��	�@Kj(��"O��z�ƀ>"B�����"*TC1"O*x�
*D4�i��3"�|<��"O�a7���x�ɑ*Dd�:�*!"O�-(�k�&(���Y��w��l��"O�l�f��&(C℀7G�&�\)� "O|\h�#�b��� ,�|+&"O ��2,�7!S���
��8|�1"O���`�1-^޸J��d����"O��� ߁N��E���>��Ԓ�"Ob��c��CN^YH坫Y@�i�"O��@"�c��l�Cˏ�G��\��"O�Lv*K<){��Y���8�����"OL]�]�n5
��掹1����"O�ܢ�4�b�H���!G�����"O��H����>�NE���7BK�؀�"Oh�Q�.���d�aOF)S�m(�"O^)bU�N WVX�2��	onµ{�"O$9�7�O�J�}f�8]f	i�"O�ap�cL�5��H7gԓH�B�H�"O�%#�H�>L��Q�2)P��|�{"O*�9�+�~�ڐ+R�Nº��R"O�pF)f�ȸ�/�@�|��"O��3�R1+#1S�v�K�"O�U1pBD�FW�d���N�bx�|s�"OK���=�ѠD�ie���"O��h��O���H�U@^@����"O�dH�`ћr��lbA�N=v�\�Q�"O:�r.W�����H�;�J��"O�D���i�@�cMW�>���Q#"Oƨh� ��~:­��L�>�4��"O�Vdݫ)%��j�?V|�S�"OR�q���G��H��
zf"Ovq3"��	�,�+bi��ڂ"O������7>|�*&���`�"O�9�5�`a�	9\�:��iW� !�ě�B�f��eG��.���v���#-!���)��@�C$Y�ڕ���7!��H�����>d"YC�o͚C1!�$��6]H���JW#F���ڝc\!�@�GU>x�qo��k]>p(��!�ą+,|<�b��:Ui��+�N5)�!�䄔��ɡ`�V=,��-ΚE�!���4w�xCV���b�LqslƎ&�!���}5�����t����Gh�!�$ܷ\�Б�tȄHF�D����`!���Mt k�A�H7���u�!�D�n��ʓ)�<@֕c�c�: �!�� �2	��)F�i�*��0���!򤍴�Yy�N^�^�H�[��Ȩy�!�$V3*0��b��D&�E2�(�6nS!�� ��!��-�.� ��ڂ\K�"O�(��	�V��2	��d�s"On�� ��|����3��6~����"O\d��i�N�hr�$d����"OԹ�>�� s�D�0S��"Ov,(ԧS+eu��j"�W	�0���"O��#S��Y��$�#A+5��#�"O��	Fa��X�ZY�'"O���r�"O�x@�Ì�;�T8��8Eyv)�a"OT���Ɔ:-)�n��;f�4�"O��ycj�9	���.�����"O4�+�C�y%چF�X�.�:F"O�p�r��|碥��o�7�$���"O�H0P�Z<�#X�4��䁡"O�Ly�Díw�n�����6��M�"O ���Y�S:�l�˾���"On�1���� QJČ)(�^�p!"O�H(��2" tԘԬ��+��\�"O6<Q��¸�u�2��%�>�"O}[�a@2z��P��	�/K�*��"O�m����g�X�4�
"{��IZ�"O胣�ѦO��5`�ۖ>�<Y�"OX��pR�e����	��LUc"O�9�#�X�%j��G�3�N��r"O
q	E�G�A���# P & �"O����➖@B�q	���
	���"Ov�3��F9�~,�A&�
�i��"O�`:�[�,c��S�/L�u�T��"O�L)�E����Ϙ��{4"O��G.�)^����qM�:\��"O�5�vFF��0��NR$��"O�IPӌلPUً�ʄ"!���"OJ��6%��M�|��B�_���Z3"OT8��Mdܰ��s�ǲ-s2�R�"O��˛/@��ї�_�
KDd
�"O(|4��0�G�U4;�X�g�<1g�"S�H2˂7�l�pl\�<��ŝE��3��KM�T�
���f�<1���dk��g>1kr\�u�FH�<��
De�t��";�b����p�<ADf�5QVLK��`� ��͟r�<1����z	jE�PH�$��Ēw�<Ib�Q���X�&%��+�F�h�e�<��G3q�h�pD:$�^L��-x�<�7��!_�$�U+I*[����⇂u�<��l�ր���ռl�d�f��l�L�h�ō9�'| ���<�TiAN�',!^��Z�a�U�%��1�	\f�v}Ұ+�^�OtuF��O�q��o4;pp)`����jr"O��z��Q/*��ڴ�K�%�V�&�ɨ&���Т��L���K�'�0���>Ro���V�D̴.OJ��f�9N`�O�ۙk���L�c�:	��\*2����FH��X��QЫ��dP��d
��Hg�ղy�c�\;y�$�"%�}�Ƈ�:r��e�"��&�+r�Z�my��Cg�x�}X�-9x��e�C"��`Ä-9�O9x�G�&m�20�f��p@B��*X� r@$�Āԗt� QI�$�O���JB�DI	BiaWJsEF�O!�O�𱳩� |���ǇZ?Z�Z��R���#�SD�$I�O���hM8��P@��9zNu�5f� {MA��h�7(���'��&Xo�=�$�DX�4�F�^3:���C��Rj��
n��)��-�g1�hI�AƐyШ��^29��IV���W~8���k���¥�X�D�<!�BB�j�j!I/]k���ȗ��IqƇ�2�@��v+G��t)�N�btVCp��)k�`h�����Yq�1 �T���F�
�k��Ұ u�˹k�HR�.ٕz�����'H�9�r��7�V��j�&(�ja�!R�Rd��#b:vH���t6=��Tf�23���Ľ?��R�Y~�U�UP�}P����,*s@^���'�� ��FB�R�Za�Wq8R���O��:v��($�]�U��?64ɱ��јoӠ���Q]Ǭ�S3�-3����� ��9�NU%:�"�3����$,~%��*L��L}�S��0*�z���9�����$>�6�s�BA���N*6{P�+"+�'�VD�`��(�I��酊'�(q���zǼ��ثD��ث��E�6���w��?h���
�H=;�^tP�I�zŲ��FX�D�����)4���R���c�Z]t��;0�o	�x�퉹x����lC��9jDHEdH1py�m����9-i��s�F�WL�<S�޶t�Â6O��x�*��X,P��WM8�۰-�{Հ4�?	P/Z$ ,�P��i���̘c�	��E�
�f�L�1r�"���~B @7Xa| ��k�U�hᠯ�V� �3!�2A���������0p%J �9��S�O=�x��	�uZ�BS&ػc�Ų��ƃ~tlPJǰij�cW�\�ZU���� 	��h`@�$�d�����d,�	6f4Yu�F}�	28�!�i5�|X�'���X���6>6�p��"d�r�	��p>ch]�'�0�I�m�iR�h2�S�?:,t��Y"Ym�Q��}���n�U�M	���[$e��1xx�H�뇻{��k��I�D�9�%�5~p��~Z�)@�Q0��-.s7����gګ�1�E҉}ڼ�槈��䓄9�ƕ9`��v������7p>A��,]�:01J�y���'��fL�A��@�D��gΜM��'�کC4O�&B�Uc�L2�Keg��JC";��˗�Vp�:2|z�!�W�0P�}�@) ��"��y�f	Y�hL=e��[sM,`��I6|O5����.�|!a'm�A���c��> ��lXՠR�&�R�\���M����GB#��O�2�a�&7z��p�D�X��q��$�$�&�1bf5y��b?�0�ժe�9�Ӫj�:�e��z�L �0 �lj�G}���iY���� �),�p�*��y�f��
)\	���2A��M� �S��?q���֩���"�N}�aO�Z�$��F<J��v��0<9���&��&GڄLtL�*�DR}�GƱ;�,p�#�i�'M�=iaA��7��Q�Ϸ!,ԃun�*���(c@�y�����/�3����gEi=I)v�д{��0�3+
l�'}\����g�E��H�<����'%#� �H[%r�0�C�^��P������mڇm��I��@�1��t�o�0D���������
]��F�d@D� ݶi�6�A�-�H]+�Mг�y�L�a��� /�h]��)��w�
���'<�����W�]�N�PO?��>�F獏'�4Ec��;+{��2 %�]��LY#��49 I�#I����{@,�*���Z �Ѕ8��(��ڽ�*ń�	2�6�i��:0��"�b{d"?��i�"Y.ؑ�_<< �S#�ٺ#u
��?�v�]��\����P�<�b��N�*ĺ�k���BiOy���6R��#�#
&R0���|�OӴ+g��0Y-�ɲr!+@�xc�<�S�^)Q(�k� �>�2��ݨ=Y���<db�u�Q>�X�.� 	o�.�@�EQ4�p�ȓVݔ%��e�=4��@��#Ŷ�0h��ٳhW��#ꋅi<a{��;CL\Ѵ�W9<��a"֤�9�p=�u��9t��)�.п�MCu
�����(^�l�lK��p�<��
*^0i�C�74*\Kb�Pl�WŚLD+S*�z�}�����r�L��W�e���"Rf�<�c��q�r��3Kψ0�F�`� A ?4�x	goN�	`��~�ւ2�-Z���
+�F�7�y"5{ �u!Ӹe߼���O=�y��Ԟ=�T�pf@�f���)� �0�y�	Ԕl�`8p�;_Q�墁��y)S�,��іo?R��`���;~�6���?�I��~"o��|nmK�愂���BW�y"��H4�t/�7@�9�ɉ��M[#�Ad��Y�)m����F�%8�!��q��=��	Oy������!~��ی����S�	Y �{G��O�!�-z-� �m4<,V�N�9�qO�gQCld�{����QN�����
mk��V�&!�d���`*$a�f�(�[0�:zS2��Qa�'@�u�|�'7�rt��-�\�K�Ϙ��C
�'N�LY����{t<��=n(�(��VQ�5��ǁ2�0>Q����,��A�%G_	e���W��Q����'����I�S4ON|���@�\hqa�/ѯl�J��"O*|g�>�"���A�6s�d�w�$�8F�l���!�9����:�	��,x�®^φA�G#!D��+EL@���P�:0~��#��8Q�
L�J>}b�x����Y�)����a�ԝR>�y&�ÓV�!�� �Y"�F)a�t(�w�;i��iE&� u�$��|"��"u���F'�H��A˒��=�d*Xu�.��t��g 
��9��!�4I����ȓ�(}���s"r۳KN/T����8b`��o5hY*����]9�݇ȓv
U� ˠ/'�����s\���Ny�غ�Gܪz���;e�<RU^��t�BDQ���""~��`C�' cN���x3�\IB�
�u�n|���c�|���9�j� �❍v)\��H���ȓ,��]�p��7�l�� �F	�ȓ|��h�ML:=D��Å�j� �� ���r��z�J�@P�
W����D���� �	q"���վY�bD��S{Jx��,�Q�h�G���ȓ5P���j�*mzI�	�"mqn�ȓ2�1q��߶?�P\S��"z�dI�ȓL���Q�R�waɲ��X�EGh��ȓ�4���ѓz :�b�bT�^��_�t4�b%ATb�E���,4*�X���F���R �x��ce�,���Y�'���xT�ΚS��5�A�(�
�'��J�V3_G
��
ݦ2�� 	�'���蔣�jd��� -��+�'����qf��T�B" �/ ��	�'��X�B�3}g�9*������
�'�d}����i�<�Ï�;e`�Q
�'zq�r�Yj��8aF��zʌ	�'��Q�A �E>fa��EN�D��'�����L�\����ň>��9��'�<�y7Jʹ
ă�҆ �a	�']�`�פܛo.��УK*��3	�'|p��9�n �S,��w<�0�'�A���&[��3dS�����'o�AhG����\jqkW�p_d���'�8�)�扎p���PNޫsh49"�'�p���le�� �a�l�@Z�'?���+c`8ya!�0}�lLَy��O�z�rp��ϋ�<�A�fR���'Z��Q�|,�i !�7r��Y�'��ᢢJ.j�<��R	p����'zh��e�G��\=*R�����'�D���#p�+��J�4ƐH�'�dEz���Ta�Tb���g	F��'*�s҉[�a����v��'t�*);�'��Z׬��m�b���ɲ_�$<i�'�����;u@��"1e�Q�4���'H��BP�{�$+��V
Ji�MH�'�D	 'P� ��!�劆��x��'��"=E�@C�4f�0��>�
t!���gg6�Bs�Ocy¥�6#�����-KE|�ʣ�އ13L�X���{�xݺDT���q
�
�����O�8�ZF�?Q2��K〉\�����'I���1��M.���]U>�YR��	3�ݹ&�K�%ņ90���%��� ÝkC�|��)�q��b:`�8�d�m�����^�~m�%(�#�CJ��h�����������,k��Y!֬ɉ,
�T`��>�R�X�=�����/,r�9���4NҪa��'��	�h��Q�6,�)���5����g�I!B���t�:qp��+~W�*��<�)�'h��mA�6v�6Q�$mR�z�J��ȓW��@��3"�d\��������ȓ��0lɂp�V���ٍ �5�ȓN>�ٛ�
R�
,+�hJ�(5GzR�'�tӥ��?� �E	[�yg��'v ��`J�	�.����Hz��xp�'� 4a�f�4��`(�A�'r�ٹ�'�lKd���#6����HПǪ�	��� r��l�`"�Ѓ�{$�h�"Op<���=J6�0��"k
��R�"OL�4�Ű �l��'�#h
�uRP"O��b�ր �hb��خf����"O��btJŊFX$��C��f���H�"OVec� ߒP��P[��)E��D4"O���D	JMA��K�
�R��8"O�	���GT4:u��F}ϊ���"O8��@#�&�VI����&dv"O��
��'�貴�D�+�P���"Oh\9�jCb��5��G#<::���"OZ �c�]�0Q��fi� " -	u"O�	A'f�$-{E�ԑX�A"O$� Fē:�A��Q�`��Չ"OL�c�A�T̀� ��.;��۔"O�u���� ��4�0C{X}��"OS�&*^�P��"Ɓ.Xx�"O浑B`�2_�,�+���Ie4���"O�R��k%�ͱ��P';O�p��"O |�jIx���A>=��W"O:��t��8YÜ<i�l�+U>P���"Ox`�ע��ę�+P�x89�"OV
Q#�x�������"O �D��i���ҷ+�1`~���"OlmS��1}�� ��.p�dV"Ox�����"$����(��6i�d�#"O���&��;@�ذ��GIPf ���"O����@�6I���#���dW�@["O�@�Fd��K^�!��D�3cT||zG"O�x�u ��pz�!�<���R"Oƕ҇bU�~s��"� �O�N�y�"O"������i�/�d�	p"O�h��B|�H��%�HQJ�A"O@u˶j�>�N���7�b8a�"O.�B�&�yV�b#Êh5���"Ox͒���z���*tC�-���S"O `{!���^dꑄ�=>��"O�����#���$cEp.Ƭ�7"OM�È�2p��ⓣ�r�
"O��3��ri�+w�M��D1	�"O�e���P\�V���O�C�蜒b"O=���ڑ�����@]�� �"OF�b�4��������HՑ2"O�!P&"t�$spE>P�|4s�"O�x��iI7[]r�٣������U�!D�t� &?K�{`b\�R$��u�2D���0g�\����Y�k%���2"2D�����4�(d��'V
o�Ыa..D���f��3�-i��8������)D����C�)��mYↅ�.1bQ 'D���&��^ncf��:~if�0��0D�PQj��=�Ed_#f�D�I �.D�\�@E��WGd�w ��oO���+D��R�/N;/[>I��YQ0+D���a���7�ѝ��rPL�Z�<9І�j�����/ra���}�<�ckS=�K���d���fN���C�ə D��:��;MaPE�aI�8��C�	�^s�Sm�(J:Ł�-E�M�C�ɬ&�� ��U3E�R@#�	�D$�C���֐�pmW 2Ft3%��$��B�	%Nm�šd������F�T!�B䉃}��@��Ή|��cP��]L"C�I=3jd�򷫆t�����k�6x1(C�)� ��	�*!�j n+zy�@"Oj��s!� p�5��ְ�T%�Q"O�81파E6b)q�9(�4�kQ"O�-��.ΆZ&LT�}��U�g"O��� '�wj�²����8F"Oք�6�.�*��؜��(C"OԐq�6�yF)zZEС"O��x���!L��J��Z���p"O���p��=&f Adb�w���f"OL���A?:0ha;�c��i{�)�Q"O ��oX�]��<�C��:9�Hy�P"O�|���	O�8�c߾n���yw"O�遥��C�.T�g�Ό>�xf"O`�H�B
39x���H��t��"OX���-�68��B];H^�"O�x�pgC!n�V 	�CʰTiI"O�] GㄚJ����U��i��"O�$��\�c������)���4"O�Qy�!�'I� U���Y]�t`2"O+Í�;C��Dg6����"O
���M�9�,ܐ𭀻�|Hx "O���cD8)¤*���\�T��"O��±j�%b1<�{�j��Mf2��"O�	��i�2gbtY�L�Fk3"O��a�ތ{	�������H�8��b"O��x3+�Rw�L��Z�s~�YX&"O(�seMٖ �B�BaB� %��a��"OR=����,1�K��ŘVX- �"O8T�ՎK%Ny�5��䄨p9<=Z�"O
��ꅰAD4�z��S�+
pa"On(�S�:L����!	8��� 7"O�@�
ɽ7���x���Yf�k"O��藠
6�T��6Ep �"O4�󳮜�JIĸ�w,�+]-&!1�"O�\���\4J_�W�^�#]ó"OB����>/WN�9�,��&x2#A1D�|Js�Îo\`�˗�8a�TX��-D�t��	����d��`��1Z�+D��'N�RA�YАg��T� ˵)*D����T�2��礃�l�����(D��)V�3}�l$��hC x��`E(D����A��r�3�\�#� p��(D�����Q�i�>�k���:�zq)5n%D���1��n���
d�9$���-D�JW������-�H��(���-D����b��y�6᳖��h�hP1�O?D�$)1��2	�zLZcE�!�|Š5(?D����P�e,|��!R�d�zq��=D�t����*q̰c�
�%]��y��<D�|���45����������:D��7A��II�����[$����9D�8;���68u����3:�k5g)D�Y ��t�ְ�¬�<fQ��0�:D�|ɡ��.�t�$M��/���#D��xujɈN4ܫ��[�d��4�R� D�T;e���,c��)���cP�>D��Z�-T� �T�#3XP0�!D�8ٱ�W	�Չr`V�uzu1��1D�xB�F����U�CZ`�Q��3D��r��ڗ>;ne�fL՘GU�YZp�6D��C'O_N� �̔���M0u�0D��;��E*n��Z®ђ���@<D��Y�)���H,P�Q���w.8D����%AB��⨎<ƀ�b�;D�� �̳<����/<0V�\�"OV�$�#�p��͟�NFJ�{"O����{!^�[nY,eǖ�Ce"O��ᢍ0t_���Ae���#u"O��f��
ٞؒ��Uhc^C�"O�]�i�/`��"�HX�,q�m�P"O($�iH�E��y@���>7P��""O�!B#H�W7֍k�aUH�8Qa"O����K4>�
y:��\>���g"O�0q�	{�d�"����+xx�"O�!����jk>y�㘌}�:��"OȘR��tL�"�a��~�쳥"O�Y���[dd�j�a�!=��H�"O�8�6� �S��z���!"��q�"O\q��*�8<[�C�Tv�!!"O�	2�
;��A��c����"O r��.6r���,�>���Z""Oq37�@"zw�}@�j�p�b�S�"O���� �9�.��(��޽��"O�8�2�UWu�`��L�(7٬�j�"O�Y���E�0���O6�^� �"O>��3�M"}�N$��m����"O,)D���xAd���ǂ��"Op���E��W�L�ci��U�p��"ObD�aL�L�z���U F�y�"O�q�K^=pO<���ܲ.��W"O,)Ss�P<_�,Da�7+BM��"O�����4/�:;�տ<�0��A"O�ܺf$OT�S��Y��|�"OX�3*X!�V��EV9,���"Oz|��K�b�� D��X�A��"Ojt��3׶��AB��w"Oz���	T��pA��r� �"OHX� �ʭ6hJp�r���@��:Q"O�]�1�d��u"jv�y�"O��)!�^�q�t�����A"O�(�"D!z��i��C�6��Sa"O��ӇF�#qp��C�̿@�Z�iq"Oΐ@�DT-V���s���4)��̐�"O�M�c�R�?q�(4"��0�(	��"O��R�aĨ&,�X�A��<<����C"O��P��I�m<�[B틏7���T"O�Ԁ�F	�xW:3���[�䨦"O� b�h�1]�|H�l��)t��$"O� 2�'x8�Br����'o�j�<�nKTj1�A'۸'dD@�W�A�<9���:m�e�B��t?�,2Rf�A�<�W�Ʃ-��YIQ
�Z&�av�}�<�!�IgM����ĎC��KVgv�<QuLC<��,p�49�-�r��z�<Q� �"d�B �R`��#*T�<�`�J�rb�D�"�M���j`��_�<y�fQ��DE��F�<$�fLҤ$�^�<)�F�>���1'��Y[xE*��V�<���ڤ����Y�NY�����N�<1��N�m�4A`FO�)3���I'�q�<a�ID35 ��VKJ"����D�b�<�	Ծu<d�b`�K�l-���^�<�C矚]�TQѥMΉpv*��e,�~�<�a��,}�,����̉!��2�)�{�<�cR%/��a�"�ڼQ�0P� .Tx�<�6EU��~<��f���ybH�I�<��D�$H�H�r�®~th�G�]�<qA�Z�&-!헬 �̱� J[�<� x��K1M�!J��9Gnm�"O�Tۤf��!�̸@�<��b��>D����9Mf������x��C�d*D���u�   ��   �    b  |  �)  B3  �9  =@  �F  �L  S  FY  �_  �e  l  jr  �x  -  �  ȋ  �  ]�  ��  �  %�  f�  ��  9�  ��  ��  ��  u�  ��  *�  n�  ��  B�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�VO&}��a4/zY;�#m�����#D�D1���'�01Vo^w:,�U�!D��1G�;(�x���n�$X�6@?D�P�$�Õ�ha�v�C�y �a=D�t�+�p��xj�N9N|�C�<D�:�K�<M�N<ca��*�Ĥ8��9D���������%� .�7Ẕ��<D�L�p-��h�u W$�[Ri<D�������e��E��V).�&9D�T*� -5��dKq�߾{|��聥*D�\�t��J�9��D,~|qR�&D����O�RtN�I0�6S�L�jUC&D���f�a�R 	!�j�T���$D�d8�FD�p��a���t�L�b��&D�|��揺-����e�˳I$Z��A�7D� �Q��,YX\�;5M߾[~X}��5D�p2'����(��R�,�^)#��2D��"�V��V��7-V,�^�QEF#D�(!�c@�x��V#�FP�-&D�\:�英B>��aι�m��#D� ���9SO�ؠE�l��В�'D��x��̎j=*���?�J�A&D��Z%��.}> Jr`�89wQ��N>D��TBԖoƾp�1���HIF	!D��-�$[� ��T���p`��1D�d����S�����K�,t���h%�/D���Cn<5TP��޽2�x����-D��[#.1S���g]�?�d�Q��,D�,��'i�踰�E391`�֢/D�@�OH=�)��ƀ�M��4�,D��8V"J�Rxv&� +�4U��*O6�E��#Y���d�Ѯ8�*�HS"O�H��E�<X�b��hF�U"O�cQ�0��s�;-�q	�"O�P���,�.�8qe��N�% �"O��HE*UR�����]U�T#�"O���HIi:�֧�\���"O��[����d�@��2�"��"O�kҎ��.����o�-|�Q!�'�B��P��B_�TQ j��G�II�'<VEZ&��9/<Փw�׳*`��I�'ސ�������Щ� /���
�')�9�#�W�cp
��
тTx�'.ıRV�A�Ws��id�D�o%8���'�΀UBDE7�³j�����'�@	�W&ŬI���K���-!س
�'qPȻ�+Ӽ	��E��
.�R�
�'(�D飦�"�`5 W:�U�	��� �<(Ĥ�
N��Y��KUR��ۣ"OvtSqJݲ>,8�&��w�2|i�"O��S��^�@�
�5/ɬk���2"O�X	A� ]1앪1���
1�(��"Ỏ�F�>�`y��-��He�'@�'2�'R�'���'��'N�
 �A"t��I��޵R�0�{��'���'B�'���'���'��'��������)�/��{jP{Q�'�'���'�b�'�r�'��'�Qid&Ǹ Ub4�^�l'邑�'y��'�"�'���'Cb�'-2�'w�td(ګ6���I'Kx��G�'�R�'���'���'~��'A��'��%�B/�K�lX�5�!?�.8*��'�R�'�2�'���'�R�'�B�'�V�A���mО);�,ӎz��Ybt�'��'���'�'���'���'��Q��L1�tT�����.̋W�'�"�'��'2�'���'���'�N�Y�D�%�.A9 ��k\T���'���'	��'�B�''B�'ab�'���4��%%%�!	vMIx�J|��'���'�2�'���'3�'�B�'���X5 Y��N�3ӭ�`3x�҆�'<B�'�b�'���'���'9"�'2�p��f�_��Y{��JZ,����'rB�'���'r�'���'P2�'|�Ju�ݤi!����늏"µ ��'x��'�r�'X��'�b�j�����OtUP�GN)J|�!r�Q9���`&$Ey��'��)�3?Y��i`� �*�Ɣ`�@�,kx�С������O��<�'��A��`:�#M�Ι��l,[��'G�����ia�	�|RC�O��'J��}�f�<ܴh��FԤk����<����$,ڧ �ԝ��@^iۺ9�F��!\r����iH@��y�i�O�.�rP(�{fb��Xz�X���O������O�	U}����b��F7O|*ĩ�3"�L��D�Ew
�H�9O"扔�?Yt� ��|:��k)����� t��(c'w٢��p�X�'d�'�v7-ږL?1Oq� cH�GԸ��`�2r�|���0�	wy2�'*b>O��\"&!�2,[p?��S� W)�+ ?a��Q���NY̧Q���N�?A��W}~P�&Lܼ3��Jb#����ĺ<A�S��y��!�9c6O�3qm2��b(�y2!r�Ft�4��h��D��|2�IU80=x�h��\�* �	���<���?��-)ݴ���i>�0��U��u�3��O�E�5������K�=���<�'�?a��?���?Q��ۧJ(<�pwc�"s�h�ivD�;��٦�RM��|�I柈'?u���0Q 4��@A(�)t"�:*~D�'�7��ᦵϓ�H�����eZ�8S��@��jx����6Q�d��X�����ç&���I�Gĉ'.HʓPL�y���Ig>�ˇ��n4�{��?)���?Q��|2-O�mo�0T����ɽr]��6������部��;b��������?�+O��m��M��Ee栙�J� OӠ�Q$��B�n��+�M��'@��km=\b��I%�ӽDfk��-2T�PTm�-h�����l��j��d�O|���O���O��!�S�A��0�Pȏ�w�@��C�*0Τ��I���	��M��F��|Z���?qH>���~�6T{�Hξ'�\l`�R{��'�R������Ni�v��싧�R�(wL\K�E��;�ޑp ���(<���'K$&�0����'���'�	SE�7Z�(Y�F�*l�Ea�'tB_���4h�������?A����]�75\\�bh�n��T�FM��e��	P~��'��f�:�T>U��g 8y`ezB�� 6[�ѣ�]�&5��(��'�P��|���OH�L>!��N4
`���U�@�9�!eL(�?����?����?�|2-O��o��HH4m�qϚ��`�8�^:���PaFyb�'��OZ��?q#��xy�B 0�T�c
"�?���i" �ڀ�i]�	�L�P{q�O��/b@' RnPb���K�ϓ��$�O���O���O����|����5c���V���m�(�����ϛ&*��V���'3�����'��w�l1��g��H��I3I	� ���'���:��)V!ch�6�e�����	�7`޴JeE��N,x��{�M�US��DQ�Iny�Ob��j�� 1իS�Q�����0W��'�B�'���/�MS����?Y���?�폦z䒘���M<:=����mߨ��'A�IݟT�	���L�b`�
)p[�IC
C�]�'�|3��\,���[����ٟ�[��'��y2Ԍ���$��s�T|��'���'��'��>��	3fA$X���B&�ң/��h�ɣ�M� ������O���k�a��Չ;�m��g�s>�	ޟ�ɤ�M�+آ�M��O �i�B�RG(U���jA#	<r�����.2�P�O���|z���?���?I�U�X�a�V�h鶸�Q�Y7D�\�j)O��n/\ɸ-��˟���u�˟�ңˋ1�HP�E��iW�I�"�KyB�v��Do����S�'�^}��c�Pp�3��/� <�靤);��'Z �z�ES��L4�|�U�xc e��Il�9b��M��|��%n�����i�6��O6�4�.�ep�6��/-�BX��2%V� 4�v`O�$f�'��OV�?��47��O�|�̜`gBC��^�y��!�sW�i0�$�OH|��b���������� ���4b�.v>:ak%"ScZd0�$2O4���O`�D�O��D�Oh�?a����P)���%N�1	�����Ɵ�	�hڴ�j��'�?����;&9 â	"���S��3{������x2�'v�O>�I��i+�����w�R/r��C�YQ�z��B�_}�R�K{�IUy�O��'tK?J�镊¥`����u���'��I��M�Q���d�O��'V���ua�`t�:�I�?i��u�'[�ğ��I���S�4I��Ӱ�k�'�%�6HKr�"g�ԩ������O� �?u)1�$ˊ}���3V���;�%�f ���'mB�'y��OH���Móh!tTL�F)�J���#!H�|�NZ/O��%�	fy��p��#pUc�:��U �80�V-iv�����Z۴�ة��4����9����'��S/Ns�PC߉Ch \ �@��6��}yb�'��'�b�' �S>j�C�"�\,��*.���xY,<�nZ�^$��꟤��b�'�?�;PX)�ɏ��5#�
��7�i>67�g��֧�OTlP��i����o
���KKd'�Q#��\���A�����!�B�O���|���yȤ���F�N�⭹��S&4�v�����?y��?�*O�eo�S�Ԍ�	֟��I!#,e���@��
�2p�P�s#��?q�O(��f�J$��1�A�!vÔ=K�T(��08d9?Q�B)=�~��t��E�'0�j�$��?��ٴ�FĈ�=mpR��M��?����?q���?i��i�ONbf�� !���z$P Lp,rR`�O<@m�>[����Ο���F�Ӽ���Q��lU��m@�Mحz���<�r�iҺ7mæ�	s���e�'�`Ye�B�?a*"�ʿ#h*5#��:<vuځ�A�T#�'�i>�	���	۟<�ɷz��A�@�?V�ش�5!|�N��'��7-�'@��$�O���>�i�OX]b� r_���e��B?�9��<A���?YƜx����5w!�͡�nH"%FA+��ۼ"��ɒR+���]�QEջ��9�ԓO˓8�8�@�W rE�RVog,�����?���?���|�)O��nڧE�\���2� �d  �P[#�Ӝ�$��	��8�?�O���d��pl�%I�Р��И|�l4�f�E�Bl$9UJϦi�'
�$R�?Q�}���P�H�s�ҖJRz1q#�_SwP���?����?Y��?����Of�p����YNVHq��J2e)�Zٟ��Iџڴ`��D3+O��� �DѶ�D*W�ߣ:�QQ�HH%he'�8�����!H���mZ[~�h[�����李p�f`�Ug^�>���Z��̟�'�|�X���՟����D�D�G�=,��c"T/4B�43v����l�	by2�r�A���O�$�O��'j�z�xw�]-y���MY)�T��'i��M�g�i��O��H�eꎎO�bAx��!,�}�t�=�ʴ�4�-?ͧt$���P���*xU#�-

�V�H�KR�؍k��?y��?A�S�'��Fަ�p�[�}��Ѣ�7]@�D��9���<��p����O�űG�55�J���D4`�B�ODQoi��m�s~������Sc��H34���ǐ�Y�Tѩf�ȦG��D�<Y��?���?����?�˟�hE�V��.����̫x=���AbӨ��#��<���䧎?1�Ӽ�A�-"���֌I,A�=�tO	��?!�eω����'��$��o�F<O�;� �%+]���3�6X�~��b0O�\2ЅY��?���'��<ͧ�?�`.��Q	�5�� ���(H%��?�?�cυ��?����?a��LZ�.I . ���O��i��|��ޑx��9YW��DY����D8?���Mk`�x��@7����B�R�nX������y��'�*u�V'D�=�8݊�O��I��?�]
��_�M���&gV��)i� �'m��'���ǟ�H��5l�v1蠏J%h]�< u@�̟<[�4n�U�,OH�9�i�Ia���Vq���yZİA冡��lZ%�M��i�@���i��O�s'�+�j�LĒi��E%�	�Ԗ8z�T�2�|�V��S��`��ݟ4�	ϟ(3��K7GIFqA]�Z������}y���*���O��$�O�����dD[��	K�#G �����Y�dp��?y�4cSɧ�'q\}����i*P�0�J��N'0 B���1��'�N�BT�ş�!#�|Y�@3�]�t�Q�D'C.PZd�F��I�� �I��Dybil�:	XVc�O$Ͱqi�
e-T�0ʔw�\�`�O�$4�	f~"�'Ǜ�)f���U��ou@���C�"o�P%Ǝ�H�7-5?Y�`;<Et�i;���iʐ)I�.�j��w)F_�h��z�`��� ��ퟌ�IڟH���b�#�P�#�̅���
�3�?A��?1�i�رi�O)R�'%�'c�A��̆9�PHRX�rU6Oj�2��ֿ�\��\ǖ�n�w~�7KKv���R1U^t(j��I6J�f�C���ꟴS��|�W���$�	ҟ(��WrS���!+D�.�� t����p�I@y��z��z���O���Or�',e�AHЍav�0�!M/H��'X剞�M��iE�D ���_����n�͎I�gA��)��/7������ˁr�i>��՟4�0�|�i�i�,QH݃xK��W"]6w���'�2�'e��tU�Bߴ
>�M0o�I匁3#�J��Dkt���?���?���V�����0#�7x��%�5e`�x�	1�M��ʞ��M;�O����<��J?� �%@Ü�?�|��+	��X��6O���?��?����?�����I�,�$d;��a�F`���NRx�o��)z���ɟ��	I�ɟ��i�����)T��ҁg�V�����(�	��Şk�i��4�yr	]�e�:9q$��C�b	��\%�y⮓GrLD�ɑ��'v�i>-�I�3R 	jgꝧN� 2�S�^�b���p�	�P�'�|7݅/g>�$�O��3O�d<�!E����w�N��?��O���d���&�,2��J�]��`��9j��dj(?�"�S;I��c�i�g�'A´���'�?	�T/,���Ƿa�&]J%V�?����?	��?��I�O����X�h`򂎎��\@�e�Oftm��I\ܕ'�b�4�|%;3�.f��E���2�::"�Oj��x��mZ�'��ul�O~rL�L		���q�ViX�B@���yG�Hnm"D�|W��͟ �	۟��I�l�@�4,U2L�3#O�w��0� �WyҠe�b�����O��$�O4�������>�<�� N&A�ؕ�4��*\�ʓ�?a�h����O1�F^�~�*�84'?%�5�s�N)"��1�OL�� �?IB6�d�<s�PI@�pp�Z�y�������?����?q���?ͧ���ň��؟dZ��qn�Y7.�*�¸s��柌��[����զ�a޴I�����'LN=��h_�
�ҕp�B�=1�y�u�iL��.
-�@S�Oq���N�:�F�sE��t=�V���<m�D�O��D�O��D�O�'���~K
9�(�\��X�%}���I��	 �M�G�|Z��?AL>!)�t���,��X�U 8F��'�z7�����o;�lo~(R�3.v��f�LfO�|rRg��~B�6��)h���`��'t��͟�]NR��?A�Rp��mU������˥,]���%�H���?��B�@z�����ɔ����<]�Z�ZѬ�g�l��O�1�b�	ǟt����d��ğ�Jٴ\1&$	(���$˩d���'M� @�h�&�{u��t�]")��(ԓ�(��EW����B�'zU�gi�e�ێdɎR�#�1�?q��?���?i4GŧDǌ5X��?��2����j�)"����&�@S!R�T���O���3���զ���	^���I�!��[�O=���"���Bk�˟�Jߴ
�� ߴ�y�'��9��Ǡ:M ��O ����ܼ?Θ����i�"O���%!W%=,�A+x���B"O����a�#Czhk�����%xR���l�t!��h�MQw*]�1��q�@c�)W#*�+7��c��Ÿ��� ���d���h03@AT�2l��#�m�x��q�@	4 l���0�N�)����8�s�BS�.T�\�0o�l��Zt�C�2�㕮X�"�p�[�6r�C�-%�5�v��)�2��%-�#lC�T��CK�'B�ҍˢdY�",v�`dB�0��	�4�߽:f�����Q|^d��I�-^�m#g^�6&U �fG�PF�P�0j�qIB��ee����u�%e��N��ץ����ގ�J��	��&P�'�Fn��) l[�Nz�\j�ΉJ��ɀ�}��I2D�8��^�qO\����چ5٦�{5D��B5ʍ�R��[��U�)�S�,-D���p��*�D]S3B.
p��iFA+D��$��\M�9ѐ&Ւz��hQ�*D�DĬ�1IǞp஖�9�yQ�-3D�X�������X�!n�3%�8Z�
-D��Q��D�	w�H�K��� "%?D���V�H+DA�`��M�l��.>D��*� _/i�E��&H�5o�(��<D����k9[�i�c�ӹ55&<���?D�����&d�:�*�HR��-!r�!D����,B�HHY�M?9�έ[BJ:T���D��P��h���^02���PU"O"��@I�|f,���܊330@"O���'!,~�Z�dG�[2$p1"O %c�bY�[��$����/>�:!�b"O�ѱd�0i���uR�c��t`@"O���
S5�2d��m���c�"Of�)�,�/|x��`ކQ���p"O���s���d�xdE^.w����"O~Y�c$C�EPj���@E�>`(pB�"O��#F��>��}�7 ^S^���u"O���ۃ}�	hQ�߉g��I�'���q��EV^,��L
3�
��'YƘ��	�f�J�C���3��99�'���ao�5K��j5��1��};
�'� $��c�m� ʁHȗx��\�	�'bB�8��=�����4:G��	��� ��h��HN.��#�<Zd��5"O�x��%��2�Y���4_WT��w"Oh0�!U�H>��gGD�ei��H`"O|�A�lS1'�"�
�H-ޑ�"O���*�vq��Q���:�x�f"O��(��8J�q�$��@(�x@�"OTԋ��Y$O�\T?~�x4`c"Oȋ���F�a��k߶y��3�"O�٨7As����
�F�*Ò"O�E�¢�:P��;JI+*�n�Ђ"OX\Xo� c*lT	C� v T�X"O��DN�E"RX�@mZ=.���2"Ob<a�υ� z�1Į�8�:�'"O:M�@,�J�ӂ���̠��"O�Xi�F��B�l!6�E�1���e"OZ5�2� v�8�B#2z����"O�[�
�Ky.���C�5*�,R�"O���!a��Z�u��	6B"ObEzClʩf�T8RLJ�$]�5"O8�z�F� j���re-͉4�ƥ0"O���k�M؂x�5�K�Z��!�"O�dA�MEL[�M�"���zz���"O�x7�߭ �ƱY�i��9`��`"ORx*p�BLl��
��k���b4"O�mbw�5�>d[���9�N�Y&"O�$���^�l#K��8�i�Q"O����G�e�Iа���u�Z �"O4x���[��ؠ��L��,a´"OΙ��Id�P���;O)`=�"O�=�f��R����	O�V�
��"O�]j�G֊<�X��-"����"O"����0|(@ F\"䠀%"OI�ѥ�8\p9!vcܦJ6��s�"O�)�K�%J�RL�B�,nX��"O��â����'O�Jx8f"D���`�3��H�G*̫q�(���>D�����G"[S�q�`$ʾ,E@q2B;D��c� n�
�C#��31���P�D8D���#M���܋�B�U����N!D��a�)f�����L5Z�e��!D�|��.B%<��S�ꈬx�0���=D��Se��#"�mCq�2�V�68D��2�(A	O{�|����;c����C)D�1���`X�ܙ�b��Hж�z!�4D�L�LF����3eE<i�ޝ��.D��!�A>F5��I�-W�{��)C+D��97��=	�N�(ᓛQ�D�҈6D��P��M�o�lBfH]�A��
�5D�haT�M�?�6��3`��7p ���3D��X	�"�f̣���:Y�څ;�n3D�h`ۼYqd��2(Ŭv�Z���TJ�<A���.
-��Y�H1$5Vy��l�O�<�'�q�^�AU�ޭDÀ��ML�<�MA�

t��&9�1���H�<��ꇧÈ� �*K%���#�
i�<Q��M3��*v��4{z1�Q�]f�<Q�m�t�� 5�����P� �^Y�<�wJ�2hX�"�Tk�d%�T-^V�<����J4�A�7��3aD�ٺ$�y�<9���`�ly1���� �
��u�<C��qt�SuU> d�X�PLk�<���9M���[�|�P�Q��_q�<��	�rÌ1��6z���Q��EU�<IǦێ^�&�X6!�-���p��O�<� T�JB'X�+^��dQ�,I�@r�"O.MA�L�E�0h�� IH8Ĵi"O> ;�k�<7s �S�E
�C$- �"O�ёG�>{��a�v�Ȋ�*ܛ0"O��ڰ�8w��qa��[6CےA�w"O�]p�"[�_Yl�2�bH
^��"O��1�ϨGR$��@�E�)�����"O���"�txF�Q+ݍx���"O�ԛ��^_�jƇ��J00r@"O` !�:obzyr� е+D)��"O��#�-A+dA���nF
W�-��"O���W���qF����mh| �"O��x%OQ,;��m�AI�P�j�"OLI���}P1B��\�2E��)"O�e#����vp ���� V)�es"O�$��%�%v���Iط}z�X�"O\�i1g��&l�����^�@ȁ"Ox�B���b��Q[�w�b5:�*O��(�@&�j`J�rKx��'z9�G
�*���yg(�;�9��'��mIc˚ |�\�f���5�؊�'���P��L.��G�<����ȓh>��J�фG� ,�7-<�<�ȓC�Z�@���'?� �q־T��ȓ}U8AW�4�J}�2�S7$�2d�ȓx	���_��D�����H��؅ȓ\wvQ���ϰ�6(��'<[�N,�ȓI� S�����9@d���ɇ�^�,�3/�;B�,�Ӥh 
sHR�ȓL�� H���4f`X07ꑃlA^��ȓvn���� �gȄ�f�ת���D$����L�_�`)�B�t��%�ȓ9O�����ߠi�����Z�K�Ĭ��~�nժ�Ő�DY2��ğ1w��ȓv��Ps�!�ɺ�/	!�|��E��j%�΋{�j�``��G@Q�?�@3,O�pr���U(C~�ҽ�On�+�B�'
��'�	�R�%1�d��B�tB��+Ho���h���ܨ�G<3����$�$���<��BOf
ze���q!�X�<i6dW�L�̐�MO,K���i��TL�I)j��?�}����^�<]c���bDnA�҉�F�<AQ��3Q2$aH"��$.��g�[�A�|�q���2W ��v���x�"_7C����Ɠ 2� [��ͬaP���ώ�b�Tma$��e����ܪ-���sA�F�e�4�EN3Ű<��ν�J&�(:��2t+�M@HL:m��-D��{c��5_��pc�v�����7�x,�4A�{����C�z����Ls��Z4)Ö�y"�-��d9�K+f��X"l4��' 	�9OVQ��̘*h<l�x�ҀzBO�0�F䓦/����BC�$~���4G��h��C���0�Aǎs������9h-8U�剾}'
��=�ͪ>F����K�*n� Ӕ�j�<)�'�����&�;p����Q�I� j0�}��D�]����Z�p�2��fdɍ�yR��l亡I�#c���P����'��U03�3O��s�̈́^�5(��H���rO�q�O��`�2�~�����a�2�pu��~��8HFM�`�ej��\�b������>PqO>��qK��А%
��8;%���y��"c����S��Д�й�yү�v&!�s��97IB���C1�y�,Ҡ}�P���ɩ6K���OL��y
� <���V������4��KC"OB�bاjiX�pA��cP�� �"O �2%B�5r��1���AG�g"O�eiv@�6�ptr��ܼ55l%��"O�!��/�$l�� ړ$Zu�"O,�Br��9gL7��-hv[�"O� `͙�I��5gX�nHJ�!�"OZ�i�   �l �eO�%���"O���DGۂn:2���$H�V	��"O���o���D�n�"O�,a�[=p՜�����"H��"OR�� �Ɏ�J�(v��cҤ��u"O��� ���H�i�����"Ot��V�s!�MbvkU��Xб"OV|� ��!O��e��D�/_Ў<y6"O*%���Tff��W$;�J9$"Ol)ҕ@C)WM(1QS"	�+��{""O���T��$$ \��?�<��q"O|�36/�w�T���*s��R4"O�
�DV����1��ܘ!��)�"O* @A��-N�&���@�4AiR�3�"O.�
/����oB�b7�4Ya"OD1� ,�&OXi+�O��d̰و%"O�5���#+�r�;�Q�t�<�3�"O6H�及,Y#Bݲf����+#"O6�[�%�7Z
$#��
=;�i��"O��x�`�8@֐�1�M�/����"O�uj�/�SGl��e��>fp"O�]R��"fCꙑ�dݫz�:��4"OIHB�ޝ7v~���T{211�"OJ�{#��=����Ꮽ/�H��"O��8f��p0ѣOC�*���Y"ObtH�-V��y��ْ>�:��A"O0l�Î
 ǌ�:TÂ\��X�"O�����
��
_)tX�Cϛ��yr�3�%�6㟎W�8TSoV��y��O(c|�[a)S<xk`����6�yb�
-?��!5��s��u*a-G��y2f� bQ��G�L�p?��p��!�yb�	�@��i�P5p.�H��,��y��R<}(����7n�(��+���y�.N�=<e�wC�z�n!��ق�y��5�0i�@�qז4��!�y��V5jf$!5�S�\.�PgW+�y"`\�o@X	!�Y���!���]��yJ�>��MhT�Չ0��u*��<�y��\!����4.��)�� ��ϛ�y"@I�W��q�bַ�^������y��Ж	�f����R ӄ�L��yr�K%���@B�l�T��G<�yr��<< |���b ��.H��O�y����푅K%f8���eլ�yO��n��(b��>uU��c2�M&�ybeD ;h���� 8mJ��$&��y����V;�lC#KZ!d.��3���y������!	�0,-��Ϟ�yBH͌=bT�)�F"���v��(�y�Lنi�uB���/W�m!����y���X���#$G*f��`V�y��3=�}h���(�jZ��4�y$�*�v��B�I5�VL���@��yR��"a�x������)���1-���y2M�
N� `�o�+*r����J��yGQ�G<Z�J��Z8��0���y
� ����O!o��ia*̜0��]�"OJ��A⒞Yx��B	ʿf�<�"OT,�卐.6��=���Qhd�3�"O�J7O� _�\z��ƭSMV-9 "O��b 1 �z��'c�r�J�"O�X�ǫ�|��MRv�],	�\,i0"O�	�׉%�Vx�7���">lġ"O�a�dF1CP<� !��"~���"O"��F�"�.d��۵f���0"OHd�w� |G����Ȝ�^��,*"OB�A�C_��\-١�Fo�^l��"O4���046bU�7�C�%چ��Q"O(Y�q�H �д`#GL�r�F�V"ON ჈H�h�6H]�.�Z��"O�D��d��>ˤ�ё;�&�q�"ON̨3"�5BP�av썥�\��"O
�Ђ��s�i�Z0y��h�4"O�0�ШyQf��#t���"O*}2��K�i��()�
�^Ҕ��"O$�ʄ
h�����ϲ4Il[�"O� �C�>,]bt
�#Z0ٰ"O��k��$5����k��a6���"Oة�����c�Ԕ�𫕺&=ʵ�""OT,�Q��0���n6�щ�"O\��4�ȼHQ~)�@bҜc6()�"O�����D�*�BG>;
�+r"Oj`���v�x1i�ҰB$(�;`"O�1p����j8"5��87�e�"O~���Ži@������:/��a"OV{DO	W�b�F�8or�`�"ON�c˓N��ūs�F�
x��"O�Q3R��3n��č�x���"O��u �&n�����E�و1��"O
�#�L�D�R9�o�3���h�"O��C��I!Yl\���Ң!��\(�"O<w��o+Hy��R�
�^t
b"O8�Q0��+6칀\.�1�*O��*��X|�-�@F�;N�{�'p�eXd�Ҏs�!���1�� J
�'J������|���Ө<�V�	�'r�x�cG�X�� #���0�h���'jtA��P!�"	�Um�"��e��':���ញ$X����lU2���;	�',|��7�M�5b$8���'��-A���V�U�� �6kJ����'�eNN9YV�AEB���,��'�ֹ���|!���b-޲�i�'vص3%�hǤ���6h{�l��'m����숩 p��QŌ�3dF��	�'��� c�J�i����>`�f��
�''�R3AC�� i�@�+� ���'5� h�GHP��E�N�v�l��
�'��A�&eά"4�Q�9�D��
�'�V �$�
�V����/�&aP
�'E���K�t&�X�ҍ�>!v���'f���N�A�B9��'M�2�[�':�u�v��/r~������?HX���'v���		�A��4��[ NeJ1��'���p�܆Հ�)�i�G�0!j�'{\�I�O�<bߪ�ۇf�1G�!��'�8d��J��4>��W�8�R�'��<qG� jˀ�PE�L>Q5j\�
�'@�	�t !g� ���D�#af9�	�'�.e�S�Yhֺ���(��Q��H
��� (܀w���H�ք+8�`U�"O��3H��8HI���g��+r"O��p�SgC�EQ���}~����"Ot9� �݊!9@��ra��\$��a"O"�c�J1���P��3@tlJ�"O�	����0dj����20�Ձ"O��IR�Z<xB��o����c"O4�#D�0V(��㊤M�h���"OҨӂ�U]�F��b��b�~�(�"OdT��!�b�R���[��\@�"O��4Cbp�3'��2?{���ȓ���2�)ȩB�FX93(��-Hz���t����F�0m
��8e�@�n�6���h9����i����u�uS-r��ȓ2�8���Aĉ%r�h��8d��.@�ه��Z�ҁrQES�K�Ḋȓݰ�*�	N�O��0��0_�`��ȓ��u�w��'l9����* ���$�ȓE�=�@��>^��b�ɰ��`��OD}`�I�O��Q��%?�|�ȓj�-Ζ)�vɠ&
34�H��3��Ti���6=��b�`ės}�̅�Nk�����I���		Ɛv���I� 1)���+q��r�A���Ą�L�n��F�!+,��� P�Ȇ�q�Ȉ��CŀXƐ�g6+�̘�ȓDF��:�4g�U�1H�0,6�ɆȓK�4#��:VI��wCҮ7r���f$�]j��-�n�R$�R�d��͇ȓT\m��8~d��BT�H�0�ȓZ-�	�Bj�/C�X'+Ř`���ȓ��}�P�!Nr�J���6�v��ȓUl�����4^Ȣ���K܆�ɇȓ�m�ᮇ�<�6h�%�+Ha�|���6��j��Dٞ��7��d�4$��5:� aPV?@�a�C�
$O:�ȆȓD� %p�&X�6NZ�0C�;Q�Zp��4�fܫoܲd=��l�
m��U#�'�hd�!bN9Q1��<���',lD�p�U9p���qR��zȉ�'t�q���V�����P�{�z�9�'>�#%�R�5�xā��={�����'ي�bTD�c�=���r�\q�'�R�����-)�P�)�唝t,
���'����F�]80�6�s
��e><Q`�'Z�!��_(`i
���eA5]x���'�N���U�(G�P�B��[���

�'n��u�^8&8��eT�h���'� $�q�����o8f�X�'��X��Q8x�~[�.h�PQ��'"`Y�N��v;K��U�غ�B�j�<iq(0x�R��&�z7@���_l�<�g�����tꏀdօ�D�WP�<ipa�?z�z�*�댹�8XB�V�<Y�씘4ĭ"���5a�8
� ZU�<�'�H/Y����ώ.%�b���O�<A�D2�����OձQ��M��B�<�q̄�FMbq�w�\�����FG�<���(\��@�J���9U�ߖ%!�$ūf��@M�%g��B�c݇>�!�$���Uc��M5~6��R�e�3t�!�C�Mz�$���ͽ(�\�+���!�D�m2l�;ԆM;Ant��©�?!�X<<�d����֏kc�8ȕ�^+�!�� ��VFL!�؄i��L�}Yv��"O�\Cr
���ɂ�DYH�����"O�@�$������&C>#�0<��'�x�3t�_�5?�II��T�]Z ���'�A9�^7���Ջ��j`q�'ΘYS� _�(y�#���x�6@�'6�bt��9X�2(�L�i���
�'f�m��h�>��BC_�3j��;�'�l�;p�<Rj�Dx���C<���'g~@�T���s�$�:��<��89	�'������|z��V
a`�%8�'yPh��L,tmNɻB�L1�J���'� �h6�4���2)C�3�8!��'F�a9�ҟE�x�VJG��iI�',J�$傴L+q��J�,D8���'*N�n	��!�\!��C��0��'�i�J�-��}�^�O�0j�'�% W�V0W˦���
ǐM�p��'����%e:��d��Lpr���'����-/�@	���R�KU����'�� ��FS��i�R�D�q��'&c�!�)U&��g�/@̙֔�'�
%kԏ֦/a�Y��6���2�'��Aԧ$g}@�8�ߤ;F���'.X�� ȝKkf�3�C��$��'��(�蔤!���C� �#F@}k	�'�J��+I I��\µJ�7;�����'�Ω�0B-0t�����<�HU)�'���;㋕�¨��M\̩[§���yreߎc�P�k��L�<
�ؼ�ya/x�|9 �nޖ<�D�0��ǯ�yr�4�V͘�)�$?H`��y�]8$`.�8�fΠ_U��[��>�y�%�qh����0FHeivɞ�y2B+���խ�7���� _��y2aL�U"p�c���+Ln�ڣ��y2��D��(�[�*��M����y�k�G; 4�a(��(k<��C
,�y�%��~X��0��j����QJ�yR�@�`���3vc�j�:��I���yB�ؔ>[� �A牝Z>�������y�(P��@��CR�X�D@����y����J���s$� �X�ẻ��y��Vq�$��B�6u����dë�yr]�����OJ�W���/���y�	��r?p<e��%(���M��y��yK�@:g�Y���}�a%�-�yR�-$y �$����q�&
��y"��i�rh��j��A2y+���5�ymF9d��*Dr�vYs�#O�y�h��[��� �V'l�D�ٴ�ӑ�yc�oT�yXE��%j�,��D����y��@�_4Hp�L�c/0K�j�	�y�� �%`�jA[t>T�����y��� �F�bs�P7B����bgʗ�y�*�[)* �Kʆ�3gj�/�!�d݄Rh~��0w$�Y��Z�!�Ă >�cb�W6kl�X�P�Y�!�D�/�\	�R��-`�y:deC�P�!�$�*}�$��%� uu$��I5P�!�$S1jd>� w�Y��P�"�ڧ�!�d�"a� ӣ��7�2B���!��N!�#$ �t}��St���q�!��[?�>}��e��(zD����:cT!�� �c��A�k�dUp�I��A��A"OT�Kҗc+&�Õ�=-լ���"ODLـ`��0܄��g�H%nFlB"O.���ܓGH�0��pZ���"O�� �t�5sS��H����"OL�ٰ*F� ��Es����)�t�"OV��M
�a`6�)¬C�l��I""O0��a�m���J��?ݶ��""O�Z���Ű7����4�NZ{!�D׾#�=)��e>� ӊ�Dg!�ĝ	_f�����D��E��^�J�!�dT1<�-z�.@A'�ȶf�!�D��1�Z��Z� pK���3�!��`,����!,|ZfO?5�!�D�7���.tX���v&�)I�"O�ث��K�.�q!s�H�( �;�"Oū�h	8�5K�!P���q"Op,��̚�{
���Ə&x�Bqy%"O�h2B�5�E`B"���bi�"O¬�s��(�������{�"O*�s�P5D�����:m��4�q"O`!;�ʑ�h{��s�� 9�"O
���H!}I �wc�$F+!��
~��<f:����W�g�!���8D����#REYԂ�8�!�d�*!��|�J�Yg>2�S	dU!�D_�"�@�b�I4Y2Ĕ�"�L0!�D̗ �	���ۃ^�,�ۗ�҇i!�D��IzaF+K�e;��^�N!�d�iR��SdE�lhnqoA�pV!��4A�fH)E�4?^4���9_C!�DQ3x�:`�iE��˒��+a�!�Ā�zz��ü3[.��PV�ԊZn!��خ!���J�<5lD����>h!�$F$�21Q��$G���ڳlÏd!�$ �9K� � P2A���R6
�!�D�,T�T(���í���C�-	�N�!�ݹi.T�W�y�NP��l��.�!��B�x,(�KL)�hE�S�X4Q!��7f1�E����q'<�@�^*6R!�81$Z5�Ṗ0~�b Y#>L!�d<_x�˖,�9m�U��6F�!�$��)g�E�Q��<hj�A�� �!�$F2<���dH,��d��7-!!�D�_�m�P'Ӱp���aa��!�$JW�Q�s'�����%R�!򄉿~��`��F�2"�R ��!�ݒ42�T�@W����c��LM!�V�:$(`*]9&z@����:L!��G
>7(1r0�Ѩ����H7:<!�Ƽ��� 1�H8�bV��""!�䓁b(���'g��G���H��"!�G'
�<h��̇�ް����M�j�!��#j>� �B/ۃ}FYٖ�_�j�!��ɴ;X�G��<Ci��h%�^�6�!�3n(�b��ΨUJp IWG��Py"␽T��t*ŋ�$=*�&ߋ�y��H��L�ڤ�Ϥ^�(��T �yb˓+k�Ւw��'�n��N��y���u:���w��`Hb�R��y� @3�
\�CL�3Yv�〉̦�yRC�'D��A;����ـ`�L��y���#VZQ�is�p��W!�$�T1�T��oT`r���e��!�� Ȉ��㇈Q0Ҽ@�K�*
D�t��"O�X��*�&�d|����8)��kw"OJ��ϑk A�˘�=�9�"O^�u��3�RH��i�(9Mb�r"O|�y"1q����/W�?��"T"O�����}�n���58 61j�"OV5�I��k�*M`���.�kc"O���`��F�b%��.�:hp��
@"O�M�'	-"��+f��7CzF��7"O~�"��96�G�oj�%��"OH%��n�fM���(NP@�S"O�i��֓~�u�U�^�Oh�|� "Oz()da��-��X��Ң5`\��"O
��E �f���ц����"Ov�#��PPd��SJ��zS�"O�����X���1z�ƈ�zIB"O���$Ⱦ{v���v�Z�L�2"O>�Q���5�6�'��e��"O � �һb�t@�1�V\��"O������r�j����HR*��"O��i3HX�_����b��jE�isU"O�<��R�ʚA�`�!)�䙆"O�H������Z�����I�"O4	�P�� qč*#�I��ɢ�y҈��<H���$Tgn�!�M6�yN;DCҠ�R�W�A���)1I4�y�
�e$�	���7��L� Hͤ�y�d˫~2�i6��,)�`� )��y���Y�:%�2��P�`�PG��y��ٜfP3�ܹIp�㖌U>�y�_�*�"���B��"N߰\�`P��Y_�(r��Ƚ^_h�MO�"1�ȓe��[���Q}^D3����Q��ȓs�bܑ#MKed<��V�$`���[��`�v풓S�н"+Êc~@4�ȓ?���w�O>5R b�
.��ȓdf0� ��#���W	+���4�������g��"�"�\ �ȓ]�����!�?V���˃k�.��������k�	;�%Q�AS�Sb܄ȓZ\�ɸ��[�l$�MH�B!:�R��ȓCSإZ�!�~xݳ�B6T���ȓ_�1'��009IR_�2��Ʌȓc�����O����w:-��x��p�H5p���V���`	�Q@��e E�V`#|Qa�K��ȓLIF�#R�[
m�0�@����݇�@�PK�������
uG��q�"��ȓk?�Y��-ź�>)�s�F�[PZ���m��4��
�5k�,�a�L�[���C�"�y�W�R�y��N�d��<��BN�%�'m L�f$*4��%e��ل�k�4\CWa�7�A��%O$.M4y��RW�XxS煵c�I�!gK!H�T�ȓM)�\�CL�N}�4��Xr`��	�"�7.J	.<H�GY�U�8���&�}+����bQ�IC� ہ\�H���jO�seܲ�XE�vi�8�^1�ȓ1j�Z���x7h����1������� �@�H	*#�	�2
D(j����p�� !�*HKn(s�J=W2�<�ȓ=��H���H�dph95��?J+
y��d� 4�S�7߈Aɗ�;�z��ȓ%�T
����lP��V�j�����S�?  :!�E�<x���*�3��Y"�"Ot��"�������c�'
] �2�"O�@�O�8<xUC��;T��F"O�)x�N
`�a���8͑�"O�ѓ3�>I*��[��5��< !"O�ݫ����eބ\kE��/,HA[�"O���OV�s; 5�FI���\�"Od�QA
�e��gF(9r$"O���Jۮ/�(Pr�'_�mB ��"O|MpDE�l��f�!N�#"O�i���W�kr�Y����>��I[%"Or%Z�,2cx��W�Dzeᘍ�y�@�:l3�d�U�F� �"��T�]��y"��"� EHĉ�8v[U��䝳�y�ʈ*��J�I?l�2��bQ����hO���<�ňٯ����I�2W��q
�@�<	"%�:#Z�ԲD�ê,W
`*c�<	!ܦ?�6 ˶�L*PL0LCԈK�<�a�-�6��6��Sþ�`��p�<	nR�<��9�E��v&�P֤_o�<A�� ;�JA:��.-���Gk�<yf�!����-dN֬)��e�<�4�x� �B�U�~��E�Id�<��Ā�g#R	4 ��h��y!lZJ�<ɶR�7{HT1�J�o88���D�<�&E�b�\<y��PH��D���<�䄝�d��=��ɋ�v�� �#O}�<Y�D��d(�YU��1���p�KFA�<�2gΜ(X�@���-)�!r��F�<��R�0��@�#�'W
yX��VB�<!`
;^�x�� V��Ś��e�<���0i��gʃi��Ē�*�l�<�e��WtݑCL�d:Fb�e�<)fj�,A.5��mF�W��t��b�<a�ɥ[811��=�"<+���^�<�5� &�\kQ@H�A(Nqp�D�<q^zH�bv#̵U���ó�F�2B��"K��1�f�9rc�$Tč�VOTC�?����/Z������%���Yh<y�ՐnP�up"�^�gDu����\�<�G%HC�l���N�a�F�@���^�<I� ��1=��q�鏇_'Np����Z�<��Ӊ{�fC���w��y�f�\�<i@�@"b8����ʆP-nU�cE[�<)���w�@a��*�7�N̉�.�T�<�".�9�pU���{��Q�͎U�<qv�^�@�h]As�.�l�h�L�<��"%&C�eL�V��h1�I$D��1w쐏`t�-��A];)�8�Ej%D��"W��Vmr(� D�&*�̑�o#D���`�ϴMF���$U?zθG�?D�4�1�8e(��[@AD{�8���;D�Hz5(H�)=���B��*v(3�,/D������	9Rs��O�{TH�Ņ!D�,�E�BH���/Μ=T�*"D�(`2 ����)Fi�q����M*D��!�m��6�j�G
�
C ]xV(�O.�C��zC"�l���K��	EQ~e�ȓ]���JR��?>R ��Im �ȓ0�)9�jϡ%�2	� ՅFܔ�������ö1��yҔ
X>S�����s��D���ŧV�,�KE��^��}��-��DaōN}*�KЬ�i���ȓrU��3�M�p+��#�I�tm䀆�S�? ��
�!$�n�
���1C`0Qw"O�(����9�>ѫP���[a��(v"Or���.}��tZ!J<ZHr���"O�S�J������$�?#\�H�"O�����p3�4`��v'n��c"O�Up$LF4��<h �_�;3����"On��c���	�`�A���i+�d�'>b��;\� �!��{�a�D�O�h�p��ȓ2�2�����,�n`���=a����{k����!��Dm�%��Y�Av݇ȓ.��Q�v.��Js��Bƒ���ȓfe�,�`ΘB_ XZdd��ˢ���1��m����3 �0r�66�� �ȓ=��!�D�<� ЂAU�T;$���П�'��D��'d����+��q,a+��=�$���'F���n�+�*1qF�e3�I��'�c�Y�$61�D�LX ����']���T�_��*�E���y2�]F��ȓ��A�@AD`���yR��
3�f��1���$�lt��jS��y�CK/_�@�ʃW'0������G)�yB���R�Խ��-P%&��e�2ꈼ�y��)G��|(&៫%=��3�Q��y�!ħ#�BL:G��I�Ԥ�Ƙ7�y�˛�h��C.I<<9��
�
�y"�,m�fYId$�l�X�C�ݓ�y��O�f���)%j��Q��J�y�C&g2�y`��<75� I����y«�D��pS��!L̍��+��yÓ=Ҧ�CB� .� �ή�y��7P����ՆpR t�GG��y"��	�]�������OP2�y�!�h1��ţ��p���ǋ�5�yN��[� CG��sz5	��y���6�V����@('��91�]�y�$$�j�;1+r�ub5��<�y�b
��5z�&Jm99��\��y©æZ�J�[�Z�d�\y1��ُ�y⧓�N��9��e��I���qD()�y�'ҹz�V�z#k�42V��9%Ɛ�yb�7�؍���5\\XQĢL��y�.��/*@hJ�l�9M�
��yR`��5t��I�3=�t���U�y�O�d��z�I�ľ};f�\2�y���7EI�����M�P*�yb`܆]`�BjW�Ύě"�J��y"�� 7���a� �5���9�y2/���q�T��<Y/.-VDɜ�yb�׫�J�̭Se�R婕#�y�E�<y&2	� 'U�L�X����yB���_��Ys�G��Qc���y2b]�g�T�K���9�)顯٥�yr����AQC��CXVa�A���y"a���XܓD�?��2��yb��S�8���ܷ'�rT����y�*ِa���qh��"��4�vk@)�y�LN7����DW�(6�*�y�چzt[7��:9�Y!&`� �y�,_(z���9��
.�p�P����y�M\�u��{Ƣ�)�����y"ņ���Ԓ�iŐkO�=���L��yBi��|�h�%%^�e������]�y2��wH9K�c_ /��1j���y2��|`�pR�71P��� ����y
� ��;���X���&K΋@��p�"O��)QO�t	�yz�iG>|�LqR"Ob���ɞ(o�ұ��(�$�j "OF��f���t$��Ǔ�F�:�I2"O2�K�f�WR����R�&���!�"O��:Aā�!v�3d�	E�.Ԩ#�'I��'��
���7f�B�1�I��`H�'nH��@^�t��5T
�53��a��'�v��5:H���ş(l4�!�'�8Az��Ț)^�5�2m��T-��s�'�ʝ0%*�}�6����/@O0���'\���c�q�S�M��4�L��'�^�Ɖ�-6= T	��1������?Y
�D�|Ys�Z�W@��q�n^�H���A,�pC#�J?*d�hG�O���ȓl��Bv�4�>�����~@����ް�RQ�P6l��'J�??���ȓ|L��x�&��<�9� �ɀv�x��ȓ:�(`2��ʦ	�.a9�e�>��ȓq�p���)��V��h��޾NIH��ȓĒ0 ��T�B� a�5ϲn���!��}iqiŰm�J�KP�E.��Q��,�p��gV�
�D��2O��;�4��-�:���C���������^��ȓad�X���_�v�kP�`x*��ȓJ$6u���\�$�nHo\���L��'H��q�.#A 2���|�N ��'{�<b��8��y�Wg�80�B�	?+�$�h�#�� ��a
±��C�I�}��I�d�R/bW�������DC�I�0:\35�!rx���
ܾ,i@C��.�q�AaH4�,"ai�1�^B�ɯs`�	(�I�s� ���Nػ~.rB�	�j��@���͐��t�󇙵q�|B�I+MX CG���,Hr!�p�U>B�I-��r+��P/�x4	�:��B�	-+8��𢎐D����>)P�B�I��!��%|r�
��B�f�RC�6`��hS`	�$U�� ӪG=�C�Y�h����
�u�bD;p�ۃa�&B�=yf�@rrƞ�gBjLc����JC�0l�a�&9?NdJUI�/) �C�	�A��X��FI�
r��xR��M�C����س�(E_3l���ܱr��C䉂 �X��7/P��� A��C�I4Q���fe�y�&���C�Z�C�	�Y1RA�7c�+pMX�w�ܗA�@C䉰F��EY`@��4Y��nЩ[��C�I�3֧?̶=p�
OxX�C�	�.�h;E�z���H�ΰ��C�	-yj�(GΓa�\s�96ؠC�I0&� X��  ��K���w��B�I�d��BF�ȸV�0�M5(	�B䉵!��i��K؃ ��Ti�h�c֦B��1[��d���&Ln<[t�Z��B���zi����p��e�'%�d3VB�I��NQ�cW�-g�-q%ġ+��B�I9kŒe!
1*¥YQ��N]�C�	�0�Vq�"�Z���\ ��3=v�C�I�B�,�*!��$��K�W�B�I�&(�4[��G"��଀8n�ȒO��=�}���2��ǌH�f��0��HV�<!��M�O5�<P��)�4�ub�O�<���1;x^P��f$�<�!`��K�<� X���a�4e���vG�,gČ�"OJ9����w��<��GM�\6V�i�"O>����R���i��ۮ|I1�g"O�%���$�:��6�̋;4���_��G{����Z����iF �����f�!�$ܦ@�v=Bum1>ɮ4hݽ<!��� Hz= ��V�TP�!��*�!�N6z�}�iG�^���u�O/)!�d]"O�I�Ѩ�s� ��/ԋ!���SX� �F/
���U�!��Y� hip'�����H ��'�ў�>�3�E�"$
���-Xd���5�?D�\'MS� ��'K�G���G�2D��S!/t�1" �n���E�;D�TR��?U"�y��^�#M$�I�N4D�����P�V�X�o�I��kq�$D� ����4G<i��J�
XSZ����,D�l8�AY�d=pay���5i������*D�H���ܒP倩�"i	��P��N=D� a!�/2d<�Y�ܼl���J�6D�D����%@���+�hL���(D�t"� H�L��&ưW�Z��w%D�(ð�:w��y��O}>!�#"D�X�H,v�"�2o��5e��6�-D���ħD./߮�B6�Q�&�ٷH,D���1"ޑn|�+ Đk��[�+-|O$�D2?�b�"8�|7$�Kεч
O�<a��=h��*�MռZ&^�!�$�M�<a�F��x{�h"c�:E!�g�D�<�E(?��i��H m���a4bY�<)��,Ly���
}
�d��T�<٣'�b�P�r�BYKF�"��_Q�<q��I��J�jZ�7Ϣ�"�I�O�')�Od�)��\�\�@|S��E�0����ȓr�j��/��G���jU�&x� �ȓb
�����[i���Bv'N�Q5,��<?>� �4p	�Թ�'�t�5��u��=@��ڦk2x% R�V�8)����`2�A���EvX�cU���\��v\t���HfN���M"AZ�'���Id��DUg����]�w�U=��a�5D���E��cYB�Q�+�M]�Iq+2D����)y85b��ԔW�֤��5D�H��EB�W78URD�l�b����4D�@;�,ԝfblQ˱� c,@�rA8D��*��V<��K#�ޘO�n�0 �<����
fT���ա�R�ҙ�Cغ[�<�=)Óa!8E�i�/� {�#��D��w��A`)b�"c��R����ȓ2�Xly��#�r��������y�BT�1I^�G�,��1�ֽː��ȓ{U@�W�EZ$u��F�h��!A�����R�;��4M.�F{���<��3XG�tq`��0{���3�^�<كG�i	Tݒ��U�:@m(�CW�<�G/����a��,ew�H&l�O�<A��įo��Z�����ț�A�<A�xK�@��C:�P�3��r�<q#BY�1�C7�ۄl3��"Gl�<������t<��O�>\�q�l쟠G{��ɞ	~�h����B\���E�F���C䉟I{^%���T�*����oD�k����0?�p`��itT��m
.fQ��h�<`"\+~�p�) o§LYJ�g�<� PM#��5�؀!�O���8G"O|��*	i����%%B��Xg"O�9�ת�C�pը�*�+><br"O�˓�ǅ4�F 3��yq��{'"O�|(��
0z�<D���Ӕ']l���"Or
�+���z��ǋ��W�<�""O����	�\jD%_�@D�p"OHrt.\2_J|�ˑ�py��4"O�Hyq�Z�*<���#��L~�#g"O& ���	Z� Ѩ$h -�R"O�<[���P�FP����H��1��"O�yQtbA�C��`���=[�Z2"Oe!îӊy20����̱<PBRS"O��+�ur\�ZCMK�a�U[�"O2���Ef�٢�J�`qQt"O�X��
-=d�%zw*�)&�xQ1�"O<ا&B�VP�Ǣޕ#�:�{p"O� �b-�<�$�r����:%"OdE��BV3Kh�h��a	������"OĀK4(U��@��&E�W��x��"O�y�Q��/kUD�	��G�#�4��"Ov�eFj�<���ގK�$| b"O�E�b�X�i�:r�i�{P��"O�9���R,WVl b�B]4^a��Ie"O\,rGQ�(�f�xᄖ8]�a"O�f�1J� ���Bi�F铷#�<��nnD0&NО,�DЧJ���|Ş<ó������a�-��ԅ�'}t!@�)�����gP){H}��V)��S��5P�+u�6 �`�ȓ�؉�g��zT`S""T)F�(��p�B���H�6
��*�bG)M]ƹ�ȓPSd
e�1^|��NĥVN �����!g��.�D�9D����8p�ȓw����M�"z�h`�P�]�!���NI�lSqA�8��If�в4!�D�����[�I6AVV��E�ӳ�!��1Z�*e��g���1�9�!��qÜ�ۢ!/�\����Y!�d�A�L�R@/Q�.%��	�m�!��V��:�"��w�lв��;�!���r�����ϴ�,�c��Z,�!�d!⺰;�L ���T	�M�!�DN*؜H�e�6>�@ȚVl��]I!�$G.$(@)v��79�Jy�#�BPQ�2�)�dk�B���#��W9O���C"B]!�y2����ɐ�Ј���Xt��{Ј��SH�UT��cf�愇ȓN�������M�X�d��0��D��P�H�Q2�	�u)���g�����8h>�aCM �p��ӡ[�$4��u.A����tw��(���7��?ɉ��~�ч�Kq,��$��4Ct�jՁ�D�< ��=:@i��+�0b���g�<� �]��2l"��_��P��u�g�<y�b܄K �P'�?O�1���b�<��"G�7]:i��:r|��J��QT�<	ã�9��T§B��Rx�����V�<I$/� v5�X�^�1��y��NQV�����n~�  Ӝ!V��'`��,�q͛��y����Tb@$���Đh��� ����y�bŨN���LȨ[�n0I��M�yb��VN ����҈E:�y�m���������"m�t�٥�y
� bȻ5!O��hԋ�g��E��|�F"ON�K��K�2�yr�Ha=08�e�F�����J~"��FҢp@�M�>�L� 
���yʛ ��1�°I��b��y��m�@-��.M6Hlԡ7Ő�y���t�ƀR�%�%=\�ؑ�W��yb�%�-R��Ҕ4Ѿ!�ai�=�y�AY;vI��S�cW���1���y¦�7	���#c�(<@`�/�y�͇^���
"���_��p�gL��yr(y�F��0h(�� @�б�y�����0�+Q����n��yRJ��yf�`�����H�� )6"ƺ�y��kۆ�Rq�į>(�pJE"��y�!�*K�l��./��tp�ŧ�y2DL s���Q(�<��݃����y��D�Wm�QI��`��M0@�N��yRM��;�(�3%_�S<�����I?�y©�.$��B��M>�:A�1�y"m@�n^D��K?3����k��yr�R M���Af@	�U��X�Cͅ��y2.ӊuΈ0D�I�EF&	肤α�y"��/I�t���U�1��ZK�+�yr��$�Dm�)"�� Ӧ�؊?!�D%�e�� ��5z�P$ 
w�!��:WC��95a����b����!���EPh��Ӫ?�l �BH_+b�!�$_��4�Ⲋ�1��|�'ȣ)v!�d�)%��ջ�(�z��"��#Ov!���
��R�Ԇv� ��C�X�^S!�$C"h�x��ԦD�2�(�2��� !��J�q�th�F$�c�<�4
M�L!�Dҟ~AZm�L��
"V0��ȟ5b !�d��h�e����)Q�hH�ö7�!�ĕU˄䒤�ΦJ'|����In!��]�Io�X J�V�j�F1g!��U-D���
�9A&�+EPȹ�"O���C�Z a0��A��#|;�.���"�O�5���Шj�z���DW�Z�J�s"OL�r�Ӌ5�Ή�2Õ#}���@a"O蹲兙�ok:�R%dH,IX՛�"OV\�i��8[x���m˫26��J�"O|r�h^.PM���K��e��E1�"O�T���!�|����͢#ll �`"O�X�!�� ���K'�@�4�X�i�"OJ��L� _�6�����3j9��)""O6��Ũ�.m�R\x�kG�*�0"O�d�G�����C"%N�cr"O´*2j��IQ��Ӗ*g*�J�"O�S뛈.% *Sp`s�"O�)궉�m�l�T��+YN��{�"O�#��P�H�H%
7H^5��Y0"O>i�F@�b�����@�*r=`p"O���q�X�Ty��R̶6�8���"OZ�hƤ����Ƀ+��yZy�w"O
����["�C�ަ.u"��"O���e%`�I#�F�q�#d"O������v��QVF! Y��[W"O<D��R���B%��<Gj4��"O�
g�v���qoG�4aH���"O�M�u�G_W�\��+I�Z�d\��"O��4o�;R�e�jJ��(�"OB43�b^&�X�
�fF�j�±b�"O�Y(ՊW�j�Hb���R�~�2a"O� ��c�ď�(��W�LĀ�"O�lk$�^T4`B]���l`�"O0��ހL:B �V�e~�k�"O�x
���^F���5�ާ>� 9Ar"OX���R�B��"U�@�X#hiH "O���q�_�5u���gcWs� x�"O��x"��X�9p�":R���""OF�9g�'�@kUŢE�\rgO�m
�U�q����N[�� �	9�!�$8��(c%1x!���i��u�!�D�c�L9C�Lb~�XXqIA)2!�D�U���gE�.Ey�,`r��-C!�Ę�v沘�l��?b��i6j�$.�!�$�$�fxR$�V+-�<��0��/U�!�D�5T���*���	���L����
=,�^����.Z�H�9��E�lE~C��2 	(����7�PP�PJ�7�hC�I��R�Y&-TWhѱ�O �O8C�IN��93�ߎe�6db]g'"C�IΠ|����a&,��Hk�B��81��}"`�K�b��l�g
"
A C�I�sIPhʠl����v�4B�Ƀ\��DБ�F*�Rl�'(D	Q�B�9g��=��T#VU:��%�C䉟s����� 6+P��^Q���	�'�Da�t
Ÿ8~�t�%M��Gv�`
�'&0����+(P4��Q&T�P�'��Q�Dj�-%���J��ũ#f�T��'���@�bQ*l��-֓RA
���'��A�TNJ14 ����@V��-
�'ӆ�餦L�wL��Q��*Lk�U�	�'��u�W�S�:�Kq���IuT �'��(��tf�BKΞ<5f�(�'LȅHDE�.L������7]��B�'�����E�h�p2�1$"�	�'È塑���� �v�$\+�'3�C&(ď ͠�8��B�!$X��'a^43����u�����W ���p�'n���!���M��oT?��'k8�2�� ���X�+� �ɩ�'��|�ѫ�%�dH���	<aJ�y�'3��p������!v�@�D"���'���u��>A�}R�#�%�h�<i�_8���Aƌ�1nҒX�FLN^�<�b�JJpz��TI�91�)�X�<�%*�mR~�XW�B�x3r�(��NT�<1&���
<�v"$eĚ���n\M�<Y �T�<1��ag�["9�8b���E�<���� ���:jX���JI�<)ABnt&zp�� �%�o�<!�G��1"�L{��LS�N�tʐj�<a��5\�$h'D���Л�%c�<�u9�z��R��= ���y���[�<A���$'b����P�x>B`9�Yl�<����<c R@S��-B���@��I]�<����n��<���Z�=!����S@�<�p�σ ���1��+����\{�<�$f[�b��,A�#λ;�*��v$Ax~re���0>Y�K��`�����4�^,�P�Z�<�S���.x���ڂ�h� K
V�<a^ɠ� �-*�p`8�gUR�&=�ȓb0��ReKߊ5H��A �$��ȓX�d&b�%n���1��A��$��Vs��;CJ�}���e!6r��S�? DT����D�v�� Qv	($�|�'�֥Ǎ[<��;hR.���9�'��0dg��r�
�Bч�9d�x��'�r�&�ݒNr��b�L5E�q�'��ۡ �8x�F=!0�n�j	�'�v�C�\GW�H�ܳ��
�'�$�;����%�J�+��,��E�	�'�l�W ��	�ō
՘}�	�'�>A�ɏ$8��m�  )�|��'4 -���^�?�V9[�G�3��<��'��h��X'�`[1�_�G�N ��'��ih �Ą-����@ �@�����'�^m@Xh	G��)Sd1Ӄ��y��&>n��SgDF���eFP��y2�*e��&O��Be�X�����y�C�$2xa�"P(;���w"0�y��i�<e��<7�9��+��y¤O<b��$�3�؎?hcg�֦�yr�� �.1��Gl��h)��y YH{�D �-�J�t��yR��o�,=3Qj��4EV�j ��yrb��
�($(��Y�&���y� ���yb���xID3��E	Rm��y� 8] �Y����2�4���́!�y�i��X����)���
��yBA�z�T�*(8����F�Z:�y�Î�,�h��߭-n~�`�*	��y��>gv�2�������6�y�,jA����!H�hѭ�y2`A:!�jꆦJ9r pS�J�yb"�s�8�E�U9����RLH��yg�	�	KW	J88r���y�E�Dv�P#�}�.�x�bK��y�j�&4�fi�U��3y��r�m���y�Y��QRĎth<q
s���y"�؊ -�pk�,C�oe��QŮ+�y҇C8_|,paǭ�np�����y�M&D�0��DkB���R"�ybG�x�X���^�e�D(���y�*Y7*
���� {��B!���y2&חK�HL�֯h-l|�kQ��yB�04�Uɋ�c�@h�'ſ�y�g�7r���E+?Y����邬�y2��%]�-�Ɖ��x�D�S��y�	�=	�v�^�jp�
�S��yH���U�	&�<L�f���yB&�d���c�gB%y���y�̎O�b�����mJM�V+[��yr���M�*(h��H�8{ ����K4�y�L	#�����>-4�r���yrn��o~���N��y����f��yBȃ�H5 � �PrԨź���yr�ٹ!2Ȱ��_�e�B�v���y2�	<�6�C�@
�
��)+V�ė�y��(_�r��6d�����s`�N8�y��]A)x�*2ɐ��ǅ�y� ��+Ȃ���΂vl�d��'�y��G�3�uB��2_�����(�y#���aң��-;�t1��+�yr$�Z^}�G��P��\)P��y�mB�4���ؑ{N�P�C��y"GզW�X5�3�ìb�dLpN���y�H��@>��v��]d6�7�W�yB!��|V�u0%�\�9����y
� 6urH�p��8cg*ߘ�H�A"O����LѓM��a��3O��I�"Oh�kQNص/؈p4%�]>F�A@"O<qS'�ԭ%���:U�͂!=l� "O��)"��N�	��u�H�""Ox�YM�2U����W��2�a`"O��ȟtt (
S� ;�:yZ�"O���v��Y��1����u�L��7"O��Z�$|ԙ�o��~#�]+w"Oy*�(�2�L���c��~,��"O6�����.�ؑ���	���1�"Od�ِ�/w��)cb�J77�~��"O��(�A�(+�� BŮ��6tr�"O\u�u�Y)^�R� 3.ɮ~ָ
"ON���!B�b����wLX�=�M2D��� �A���B�V 4Z He##D�Pi��t2����g 6�R�/#D�l�5��8zR���AI-D^��"#D���5�3D���YwaF�`�B|`�&D�h�Dֽd�"	S���rB�� E�'D������&T�8�#��7p֬�6�!D�|Y�%�8��X�c�vqtY�1�$D��+�$�H�^`GX!L������?D�@R�gO�Ͱ�BJ6?��eQ��>D���ckk�Fׇ�pn�@CO��yR��v%�e�R��@��4J�o�yrIQ�j5��(�ȋ��8������y򅛨c$M�u��z�x� ���y��<y��F�V���f&%�y�Ϥ�I�(���!�!��y"����`ǧ �"��߀-?!�DV�MX|H�%A�9Ft��d,�=:/!�DO,
1�Y!�F�OG��23��"!�ǁ"��ኴP��KBbA!�D�'b{L}��X#`��ݢ�˙�Xa����b���J������Blߵ�y�������̴X��U�Ⱦ�y��L���,��%@37�3�I��y�%K8.ɑ��&-�P��埞�y2�(}q�C)�Q��X��y��T�6�D���eܙ"�(��FN��y�m�F �m��a^���%�Љ�y���Lڑ9�
��4.N$1����y��P? ������\�E�wN�y��.���[��ǲ���q��3�y�c�[P�E�Q��y���4���y�Xo.p��%F?�ࡹ�E 
�yҏW�}���Pd��l��%*�M@�y��D�=8�� �ߐ_?�PC�٣�y��ѐ}@���o�7n�"]3����y¨]�uj��Ύ�=mnihݵ�y��E�J���I��Y�:آ(��A��yRL�Q�Ӎ��>a� ����y2EԺ�,T�V�� {D #�_5�y�MI�A��R�kWL鱣���yB� (�Ĉ�닂3��}h�&�yoD	8$qB� L,��aa�� �y�bʂ:H$�+�c����ph��y"�>;����Pꅦb.�	G,�5�y"�Ix����6�M�q�F�N��yR$Y*����1�S�F
y:��/�y��9���qō&l�(=�%���y�aTt�+R��f�JXFcQ>�y�n\:_���2/�\wH-9tNÀ�y
� B�A����,��A���L�v4@pv"O0�8%4-$~̂��<<���"O����M�-߰�Y�7S:��"O���V�6CF��i�m�4�I�"O�����[5LƐ�Wcʔ@)I��"O��� �H!|��Tb���a��"Opq[5H�2c_��q����SΙQ"O�哧(��Q�|���@\�=PF\0v"Oj}I�
T�v��٣!fJ2-�AB"O��A�ה�n�C��U��`�"OPq�ʙ�L�)sd�(&{ U��"Od��0�,mJ��[�b�:���#�"O�uh��7F��S�/W<�r�X�"O �)����;���w�>�Tyic"O���E^? ��Y�.�g|z3�"OV%@A�T.!�����1~cN8��"O�)P����<�WO/V&��E"O`! �bP�2�iFC4ZC�{�"Ob�ÖfY�/�$p�@���>�`��"Or5x�K��t�=��K�BU��sT"O>���iK9�.yYa�������"O5�fK�\���T�T?>�V��%"O <��,Z!@�Dx���V=4��}��"O"A�Q�AzJE�� N�R�Ę��"Ox1��]�;�|�������4�� "O��I��g��x��ݰ_��=�"O����;]�AH�#ތ|5�"O�i����%\�̩C c� �
"O�H5I��
d$Ԉ�h�E�"O*�aa�^�����ao�?�l�"O��* S�X�p$��x�"O���a�J�$�.%�jL0�`)�0"O�!؂@1Z�`(�D��r���� "O�q����!��)�'�^���"O��3�P�H�r���HK����"O��
tʀ)Hh�b����4�d�z#"O���`?,�A�"��n;�9q�"O��Kf�9��Y�&�Hd��"O4@*3��@f�(8rf�9$<1�"Oʨ��"�A�fhɖO-:&(��"O�����/K]�qc���6�1��"O-2dܵd|�5�îF���A"O�Y�"����qbb�H��- #"O 4؂hL�s�µ{$���qt|�"O<���cOa'4��10T�ia�"O��у��|���g��t;9�"O�H��_ %�ph(�eL�&/����"O`PQ�]�+t,�H@�L11ɼ$C�"O�@��30��*a�EL��z0"O���e����hȉ�d�-����"O�`�K+ H ǄR+08����"O�u"���W��p���?5�MBb"O��z��8Id@��p�_�h����"O�dC�N�%k܎p�S&͡*d<���"On�˞�a2���o߬((�)�"Ox#s% }�� 	��N+e4�hr�"O(;��
#.R�Q
<N�`��"O*�"`��G~l�!�����P�"O��b��+�𸻴j_4�ؼ�"O@@�����L�+���84M��v"O�m�#ц[ʑ����&����T"O���Pa��`{�M�����('"O<<CR�Oto���bB�'����"O���I�F~�A�&� :'[����"O� >�C®w��h ��/,Cƌ# "O�k�f@�k9����F c$4!��"O(�I�C�I-b,S�O=$�H�"O�rD�a��U��q��i2"O^������L�9��'��� @"OZ�����mr���T�x��I�"O!�eL++��<���f�abr"O@!A��I�+���"^,�:QR"Ol�sEN8z(�ș�.��C"O��@�Z  ���z��8J�R�"O:}�5��59�`�ő�P5Q�"Oԉ9����Y,��D�*jp�	"O��X���=�(Myu�R�Z�6�yB"O`: �@���\D-�Q�*<�"O�T,�,Rp��߈K�v,h�"O��ӭ�0L��jʨF���V"O\A�RZ����,�&��lҔ"O��*H�:`��!G�~�J�bu"O�E�W�F�W���7�y�"O8=�"lݨ` ǭZ�^��8��"O�}�bfJ�y׺�HmG�h�t�؆"O�$Ja\�P̜�)qO�>����"O��[b��t~�Q�ɓ3k�����"Oȡ�nӃt��YU	ƪA}��*�"O��ǒ4�u�P�Ґ5�b�""O t�Vŀ4J������U} �Ҁ"O�a;�`U1T��q�BT(|��4"OnQ��N��Z��'�D�E]()�g"O��AW?!��/����	�'JZA��D��U�g�X�kL����'0� ��AIf���Jg�]��'��$���_6^t"0�b�O1gt��'���2AǕT�a�g̯2����'�>XZcZ�Z �J�	��i��'�ڑZ0֝q��4���F 00�D��'��x:U�~ՠ`G�QE�Y	�' ���cǾt}Ҡ�W�8����'x���_�A���r�H�d�j
�'��; `�?>����a�HWvL 
�'/�h�F�Y�5!n$kae�Dx�)�'jt���$�%e��Aa�Z98K2 z�'����+�DٷK�1m�1@�'"Z�ږ��$r���G��=,҄b�'���)�dtÃ�b�ذ���:D���C��5�U D�هM�h�7D���F�2Ű�� 7���H �3D��q&d�3m���b���IȐ��0D����d�$�@�#7e��(c\9٦�-D�L3�җ;�#�ɋ�>%�*D��b,>��I[g.�{d�`rpc5D�Py�˙s�fU��哢)k����@7D���2J��J���MB��i�m4D��C4��J �]ذ�(O�ܐ34�4D� �"�!T^��� ܠe%0D���pcH	2��m�$+�5׋.D�D�FK�2H�P����$]��F*D��ڦa�����׏3�xu��%D���p!N�^�L�A2-�p�d'(D��80�ܐs�tP3�@S�S`�4�%D������
��Qz aV�roj,�FD.D�P�sʈ,[ru#�/U�w�x�Q!,D�j��
�I�8ȩ��:d�/D�;�-P��p�ʄO![�1:�l1D��f�O
>��ICѦҨZ^t�9 i0D�� T��gOI5��
���J���"O68@WY�;G�-���I9�va�"O2��$(�x�V�ҦhD�JP�=0C"O�<`�ټE�Z�*���O��`yU"O�j-Yrx$��dL�E��ݻ1"O��!��y-3U%KA�N���"OLM�fɏ �x5���e. �r"O���:!�Y�F w&P8#"OP�Y��X�S�]�O�!c�P�"OV�k�b�x8ғ�ٙM�es�"O�\ӑ�\f��9��L�'I���u"O�qp�0@� ��%M�V	H�	e"Ox���u�\���Ƒ#��"O��3���'��IVňM&:#�"O�\���A�{� ��B�"i �"O��	��B#?*n��P
X7 R�c"O�t3!M�.�����e^���"O
՚w�� FD�e�ܖ�:5ҧ"O�@ӑN��4b
XBRKC'��(�R"OB��a��lhD4bᚄN�v���"Olz�`˷s�z�[E�]|��2�"O<5���?���	�9]�ӥ"O"|�dl�!+}��za�C�!�����"O��K�eҥ)d���Lc�"Y�u"O m���ޑ �6�{ׅZ+r�0��"O�`8#�  ��9��L�&Ҷ�"O~��J�6�"T�#�P���Y�"O�YG��
^�����E�lU "OT���gղ6{r0��b���¸��"O�]�S�+
Xd��KC$x����"Of�HU��:^����G�M[rq�"O� ��u��@��L�	���D"Oxe�#k�2},4@Ѝ��f+��J@"OP���jН2�����B+
�`"O�0b��Iz�؊�;�e��"O^(��$æ!�g�Q/]���g"O�<XUf�0Y`D�p� R�4)�r"O��qE�#��Lٲ����R"O�9y��N6>E����(@+u���
�"O�]�Ԃ�TU�$:�}��(�t�3D�����M���Y'i8�xY�`2D�8Xd�2��]��Y)?�~�3�4D���'n��i:pI�K="�b��$D���jA�!L�	%�R.O"��2i$D�tˀ�Q�*-�R������ D��HA���%ې��%U('!v�{4�>D�`��hM�lS���z'dmr'H"D�X����~5t�q'�
�*a{�'6D���0͔h�T(@f��n���'D�|�qf�13�\�#��'� i��9D�4�Boӥ,<�t�O<�P���7D����7WVvmQ���,S�X!Qp 5D���-K@`�&�'LZ0���g2D��rl��-o\���@J�3-���.D�L��ٽM~`PÆMI?��H�
-D��y��AP�B�Ѵ��x��(�3� D�$V�* �L˷�E�W���d+D�,�q�@��5��,z���*OZٚ�ꗬI�$i�F��=���Y�"O��A�i	��2�*Ҥb@���"Oj��Pd΋c���,&���'f�\��oY�p�♑��G�*`)c	�'���h�2ZV�h����6lh�j	�'�bUb�ֺ�2���LJ�|ʬd���� @(*A��
���I��ބ[ٖmC"O��)��ʥ}�0����C�Ԉ��"O�)�VG�4IJy���vҾ<�S"O� @�)e�J���#[�E`��K!"O�XʧBP�.y����I^�rs|!!�"O��( �p��5�4OS'©�"O������*~H��'X�쀀�S"O�������S�F	����(}f%��"OZ8��ª���jg�G5=�|���"O1"TG�n���yF+��^�PA��"Ov�1����
Ba� 7\�Z�"O�\��Wn�<��E
�z<��E"O����H�Vs���Y�1�hf"O~p�e�]+_w�h��唟|)�E��"O�dBU;�-;'��>?ò���"O~�W���6��L�@�R�5"O$x;�m�;}N��kX�pR���"O�i��ۥm%�؃���-GKJU�q"O�i�r�ߒ1V$\ g�{,�Q�	�'��')Ԣh� ���X��ح�	�'�8��Ꟊg�dс2�V�_
F)q	�'3.5�H�7[�������U�<��'�ƹSpR�M�n����2S1`!��'$U"w��?@��A޼M3Ե��'��i�#&_-Z@��Ȑ,E��0	�'}�D�AD���d�P�X�tez��'
t�*��57`��`�]�e8�')�L
Ѩ�*_�`�7)��
����'~�Ac��*B������7�����'��l*�g�7E� `�7@ /:D��'�@̉�Ǎ�Q.�Ap-��v����'w���FD��\r�`10�ۄi��I�'�^`3��Vצh��/Z{B�2�'F���O`R��g�U�����'*�sa ���lX*��"dx��'0���F	�s���	�_� R�B�'ɖip���b���@�B�
���'���A�ԱMpbmJ�&�	@"5��' �Aq& D=�F��ѳ7�J5�	�'�� 閏]�]Y��"�Q.�&�{�'�0�/���2�@=R���A�'-*���X��L�y¢��
�'�Fmi�X.q }3v�U�j�dP�
�'ξ r J�<�ځY�7t��*
�'�X(A1 ш)&�C��:��4�'��l9�m �"%>-)�mЏe2��'\8�Xq�#%9�Bc�<s�'ꎘ�'݄/D�9!��X�P�0�'�B�c2 ��W��@�N�B��h�',�A���2 ����#PKX�x�'o��J� {:I
"mV"E�B�	�'�d�c� Ea�(����5���1
�'�
�O�ii ��b葤,"�x�
�'���%�Z�L��c�!��	�'����;lnyHb��(yL}��'`rX����ʸ����.�Ԛ�'Y�8j�0A����']޲�j�'����Ǽ0���'O�d�
�'ټU[��\�G�$E�?���3
�'�N�x�MO	A
�`r���IRZ�Q
�'��lX�I?T�n���1����'��鋴���Fl�\)�c��n� �'xFm*�b֨^���C�H�4Td��'^x��@�+
!�DR�h�x�
��� (�6�C7~�4j��N�`�q4"Opd���h�|(*bcZ�t��#6"Of����c�|! "̑�.���"OU�6���8f��@�\=�\��"O���RGISn2|{嫋�&��T9�"OhL[�*��%��A��i�7k|��Q"O�UJ��o��鑪��7�V�C"O�M�VFF?g���3H��%+V��F"O�9֥�8(�����	�%��Q"ORT���<k<"PAa0��h�C"O>`q�g�K�����@��G�<e"O�iDf�&+���1�NȶL���X�"O6m��c�����d�:
�� #g"O�9�`kD	,ۂ�(����QUt��"O�b�P)(��a�1-F�VD(9I�"O&|qpd�6*r�(��757�!��"O,;6$�5_��6��"&긛G"O�UѴDΘ,�"�9g,��5
�Xч"O�<�4��>/���&����L0�"O��a�ꕷХK�@�<-�����"OT �e�.޼�#���'p�}�"Oα!�j��/�a��EI4V^���"Oi9�Iڞ� EQC�S)&}D�'���I�H�嘧��>�0G��G�bP��y`�|��h*D��`Z-�P�z��[:$̲��5ˤ>���
��-y��'A��,�!<�6��%k�,�F5"� �<�*�HܑD*��H7J��b��dPP#Ҡ5M"���"�Oh<�U�*N�:��(�"8=bt����]�'���#KȲW�m*5�1��F�T-A孂�q���ҧ`��bu�B�I%:b�X@#�!�5���P�:�X�C���P8��Z�mQY��,�g?��̤z)JH:ǁ�Hb��u� \�<��BQ9FWl��
���\�7��ݟ�{$%ւ/����} h��D�1�4k�fL=_����t�N�y�F�=^������
�H\5� �[�H"�| �C��$r΅��D

�Ś�'�v���S�N?xE�C#Mܲt�L<���F�,�}і)�\�BL��)���O�ơ�uK�x�V!��A�?�U��' :`�e�(�H�Pǭ��"�l�j``�'[-"��A�Ռv�v}�����O���'����&T�{���"f �@jԌS�'��Ď۝qu I����V�6IgΪw��!'�R�mq�M�
�wp褆��2id�Z� ���!��a[Xz�?�s�]��HX� �mov]�a,[�;�c��w�
U�%�<iSl5J��x(<Q��^}J\;��-.�՘ �yb�Џg��l��C�w�B��#���P���P5�q3�� U���pc���y"���.1 �8��НqL��i7nՑf��<�£tb�1�d	r�N)N~
��[�$0z�Ĭ���ZL�^��c�54Qa�FJ!c��y2�.��E��i@�AZ5x8�
�mK�%�"DoX��q	g��r��x�j��9i"\����
I�}��A���O���|w$��g�{.�r
�"::�m9��N@.��b�&�t��c\V(<���@��[�h�;_n����{?�%�By����7a��ɫb�\��K�韓^n��;�E��F~�P����!�Np&H��s&�U��#l�G��y�b�:h��#@Ś	5��h	��~��`
4h�e��18��d��pe�H4m�,��	1I}�����������ؗt�0��A�:�R���\-��I��g��g9��ǓN�0��u�	3 P�i5��Ul��E}r�]�{��\�V��} u��K� �(�/R�~��a�4��?	/h�4�`� C�	�H��Y�Ǌ�mҔ�{��L�H����?T�L�fl�(Kh�iz��Y��[%�I��OAb�Ҫ�i��5�<� i
�'$T����Ȳ��1�0-"~����;jy�0��H]2׶	�G�ˍ��S�g�e'�,��(�^ћ3g��Ih�0�O��	��O!$p��� �*"IdI�EC�qz�x���ʪ	���5CY>��'�)G��� �R5�Ѥj�X�b���9��u)V+j�*EK��*����eG�U�n�KQoD%s(���e�a�<��M7���[ �ǧ�ȃR�Py��!�^B@�
 1CxMy��M��(���6'�>w�z]�WBO��("O� R���#$Jh�
�(�~�� f�ŁK��Ɋ{���IAL2�3�I.s\��c�)C5)V��� X3[�~C�ɹ.�d49���#Lu�q����#�H��	ƓBJ9��Z>���L80p�`�$D��.�Z��ȓh���pr*�	}��)��6l�%�ȓ@z���hSos2��&a�f\��&"�|���_+o?@ ���
����ȓ2Rz'���T�L��
�� u(��ȓ/h�YV�c�Dp���SNh�ȓC�<�i�J�N�� e�
;]0�ȓQR��� YqR����U
�n���`��-c$��j���ځI�$�ȓ<�)��GInހM:p-E�Q�ޅ��M<�0��J W��	jdbYH�L���KqD<y�+	�'V���5��v{楇ȓr!4��dB-���GC@�����8��&ɤ91�!�e`B�&E�I�ȓh>��PN�9�ht���z!B5�ȓ.'<�cJ�2��5!7k�9��!��O$������]��<���O�A�,Y��	%R�Vǉ�g^��3bJ�	�a�ȓ^N�UJg��[�d����('jT�ȓ � =��bE [#:X �o�?>��d�ȓe,~D0���&~�@��f@�K����:-� �,�g�}�P$'> ��Ge��BROSF�\�p�S<3\\��}�s�5E���S��'�E��j̬���1Rz��s`X����AA쌉!���>�ȤcJ��)ޅ�ȓJ�����N
�2B:����%��ȓ{nlM�b�� %���*���8`9t�ȓ9۴u�E��$�����9,����"�'���!琴q���2~޸M�ȓTl���VJ�"G����'nI|�f5��|�P��a��w��ԋ�,]Bn����?�L��	��
gL�^�P�
�� D�|H�i^� Və�}�@��w�?D�����[����xEO@�y*�!�vO'D�x0��W9$�t�!F)��Z��!#�/%D�l(GjXR��0Xi�-��-j�a#D���2���D3VM�n��I�&d4D�����R�0L攡��*3�i�*2D�La�mJ��{eg��xָ�9��.D��jդE�������'=���.-D�dȥ��VD��u.��R���N>D���G�3<��xp��E-?䖸i��?D��c�aݷ]��R,��(��5��*O�(#���:TӶ��@ ��_�P3E"OȠ��Ҥv���r��I&��h�"OV�K1�56J���E�� �"Od��s���Q���ԋH�u�-��"O�<�-\!Prz|X�
Ƙym���"Or�H�B���L���D�4��0��"O���`�)������3�<�2s"O���F�5�*���8L� �0"O��Ѝ�l� �e��$ ���"�"O��Ӥ�]�.-*�+
|m��i�"O�1�s��q�t�آI��^m��`�"O���Z .π��P�Ո%�$A["O ��6
IjwN +�S�`�dA"O�^
���% �c�	�&!�y⣝�a-:��a+���,<ju�B��y���-@t���+R�b@J4�D�y���v�\�����0I� $��
��I�" ��*,O� �@�dN�-<n�E1sƇ��~�`6�'<�Ų2�R9W����M�XuY�O�>#h�I\<���%z�p衧O�M���[Z�'i(�v	�%^r��sA�v�� X*�Q�c��R���$�}s�B�I^l0sF�0A�" �>^W�7��g͠)(vH�[hM����}��M��,K	��u��'Z�~\cA�Rx�<��X�$�l��IW�>�
��Z�҈��M�~m�3M��rG����HOJ� �;��˰̓d���pS�'_�Ւb�4C��H��I����0��jX��)ɯp���I@�NL���Z��t����L�c���C'% �uQ
�jc�P�q���Cq�a���=�hM`�c�Zl$��wC˭��L�ȓ5� ����+�����CٶQ���RqK�{��b0�>	4�q+UJ�-�h����:��%/�4-�ZɗL\# �!�dA�M�<:VEĿ`G�Q�b�P}��t`�aPH�C�D�,�VxCU7�Ԣ=��[zYkcɂ�0ĉ��^��ǁ�=��<�6K��r��Q�r/�l�� "��F�xp��4.��M���a.6)9�
��k�@y��[�53n"<A��,�H@2���!W���JK7��6�`@�&���
O%!�Ĉ>q1�eA5�NB�k"j�����3GC[Q��`���#������(��s �� D�r��F��?����c��t�<��ꂑɨ�CP�ġ���S��.]�&���9�\4r�L��0���'�hO$�y�$�+`�N�i��-b����V�'�lˤ��7^��B�[:/j��0��
R<�ST������[
��}+)s
(h��L��kѳ�(O1�P��(w 8��ѻ D�˟�c�:6,
"P�0x�MG"O���3H�7�^dI��37��I��	�>�,DJ��D� �:,C�Y�>Q?�$�0|T B�.4Ρ�Ȝ�|!���B���F��$1T�G�X�R��rhD����#dL=St_?#=���x�4�3�4�`��gqX���	ϯ`^
��7�T#Q\X	�d�z�:�Aц�(QF�("��U����`^jT�h�N
'�>H�7k'��(���fܠC��)��
4P��1�)D��J�t!� }��)���) �ti��ID�]��ΡNH �K��)�'M0,C�<d�BC�M�:����.��(��	WJt�"�n�3b��t%��*�Nճb�ay2h��T��?2�J�"S��w�!��6<hZ+�<rTLzr��'?�M�ȓ(�8!8�B*W����4��!Q���ȓw�"$��	�����N1艄ȓ)�\� ���/"���y�EO<UF������T`O_�pmAQga�z��ȓ��h3GI|�u9e��>F
��ȓAtJ��3����q�"-�>�ri��hĐ)��ۙ6h�qqC91#D��ȓT}� �����"��?�����8g���?�Q�u��-ȅ�_s� �q2I�Ԫ�'u���A�"��'R�*�F�`奐�������6H�fX������j���J˺"U�]�#�X��E-��'���ȓ ��ћ5l΀$�B!�œ�B(�ȓkS h(�%:LHIF/ϋ%�$�����*S,E̕���	O����|�̬2��B��(�z��E?OLr��XUTq�BHG�w��%�I��f�Ʉ�%8j���i�FH����qG\Ň�IO��2�+�lնuT�W��*���zEtla�i�*;�ꙛ����o׮���!�ʝqS%@�BFf}s��v���Q�Z��'�F-򖝚@�V;h�̇ȓ5�f�i�"L�i#C3d��ȓnR�x��ܠ��!�60U�L���J2����	Jqr���eصHN�H��u��}Kcc�#0�Q�V��
/� ��S�? L�� /��Дpp
Ax��Q�"O��i�nΘE
D���85�52"O��@q�N;�@����G��'"O
$��J�"�d�T�}1"O�0r0��4��)څ*ښ�ر0�"O��C��+����vN�p/�%i�"O�\+�W�	�֬��ښ~�@AB"OMR&�ǁj�P�zB�۱oh�z"On1��%2z�p�{�cܩZ#j�p�"O"apu"ז@�6�+���3 ���"OdX�4�%&\b�(� �s�
�Y�'�y�$�9 &t����.%t�`��'f�}Af+V�z��7�ȅ�t�1�'�{� g��\��	�(&���'��d�A��P4�bd`!�,K�'8�աrc@�^��4�^*�hPx�'��< o��Nv�@���
� "�e��'?d�s׌��:`ī"J�F���'@����א Wx�6�ɬr����'h��l�2 B��D�]�dVĝ��'A�$�@'�<-�T`� �ޡ^�ua	�'�x �%��"|DꐅɜJ!.)J�'�j�['�]
#o�q1�A�ek	�' l�!���E��|��n�A�����'�L�i����p�(�굣��0���x�'@dᅞ:CED	��H�y
��	�'Cx]`��YF�;g�M�4�C��V<�)��E{�S�O�Z���'�� ; �2���!@"ObEQ$;)wةP�'��.	t�R�@��΅�=}2xYӓ&UKG-*��	4f��N�\��I$�0�Be`��E�BD�a(�^��8���t��!�6n$4��臅@� `F���.�;2�As%N1�i��1��� O̜8��I��lAr�f��>0>�`�>b�!�H*�D�`��9ghX�n��0φ��@NE��ڸ�F�y��ʧ	L�dI$x#t%?`ȉ�U7D��ٓ�E>Y^�p"'I0�r���A�O^軕%��"y�(���G�[�x��ЄB�̒�.K���� �+��<��ϖ.J���RB�ڨe�i4� ϒq"�2)b墠g�
l���G~T��N��|��zCÂzh'�<���+ :�VhN	P���
�/�cܧz��ؓ�B�v{��!��0��#6�HID_�:��ғÔ	o�c�AM���CG�)>?N��v/�aܧ��OL��QvD �B�^V�9��~LT"BL�:�F$���,m�e����!����� \6B���k��=���񤌀Et��$��la���Dmџl��Ȓ\J`�m�-N�A�@P�����뉔a�XD�7,[)pAB}i��>��j2��*�J��\�S�4Âè<!��w�X���lʌ&���a�)Q��%�}���0[,e�T�R����HFg�<�@�C�1p�D�Ve�*x�P`p��"pq�'��o^t��g�I�+*�$?��'�)}���)r\��{c�1ra*��t����?�⁒P�&QR D��D�����oޡW}�X�� S�OJ$3��I	��12�G�4�p<�g"�v�� ����h-�9+�x�''�XQ�K�H�b}�&�4�l���L*��E��ȮXk�,C����4�Ro?�,��Y�E�Z�����y�1�bO��(j�B� ��T��l��|�ȣ��S*V�@��e�=	���Y{6FX�Ē�y�i�"��[B�¯cbfQ����X]S�+;"�>�26�WH%�,�I?Q������IY,Lmڶʂ�MV8 W�B�6��䐵Vv�X�ưW�\S@�׻xD��'j�0|/p0/a�H4K:)��#u8O��[Ѫh���7O�\�ȗ�	����ض�P;�~=AQ�	y⼀�JL�Vm�x���?�V񃔍Ǩ&�Hb�'�H����@�be8X��S#h���'�S���k3��z�ԄR-Zٛ�@ް0��>uL�=5��m@G現`:V�	�l#D�|t�ŔB��り��Y�6X2�D�VP��9-��I��	� (&�O]Vŋ��xR��-\Ozl2��o*(-�� ���p?	���D�biCD�4��`R��}Z���lδ`I�$
cA�%�rU��eQkx�� |��ց�X�@1���������60d�tj�S(���휆6:�h� ��}�bGE^�VL(0dh��yRB�L
����샘f�ԡ#'�����g�5�2GV����l�n�Q>u�qk��a��̰�K�D���Zs�.D�t�`�ƃ2�t�7Jɰu�t;�O5j�`8�H�6�^�g̓=��0��16���-_NHx��RM�u�PF��B����Qi��F��"�ݗg�1"��'QP���ׯgޚ@C��qn0��'��H�w���Z�!c�� �rM��'�ĳfC��8#����Bi:�]2�'BL�ͪ���RgI�m	Vp��'L������,D�H�`�Tp��dJ�<�Y`4\0�iӺn�V�Ff�M�<DV��hmx�e�9���ᓁ�J�<�0쓃m庄�t��:m`��z���}�<a i�?Z�� ���>/�)Z�b�<Q�k�"9�y"�Y54h{ׄ�]�<��ɃF�P����6�dR��G�<A��޵s~�|z�nG��u�p$��<I��-����� ���a��~�<�`1פ�aV�0���Z}�<q�c�(�^�c��ܼ*�(0��@W�<�Ƭڷ��)2Ǚ?�>�+��Y�<�Fϕ�Od��"S�@�Q�[b �U�<��n^ �6T��%Úg��![���t�<�tiU1I9�Hc�` �YT6}[��Ty�<A��@��L� )�f8	��@y�<���95�Y��l��I۾�_�<�!��RI��b�6�"�A��A�<����P���Co�h��t�Sa�{�<�G�+`�n��J��:p��ąv�<פӎ.��@f�^��`�w%�u�<�6�˰5
���ғseT��Ev�<Q�K�D�<�,
Yv�=4�Yp�<�Uo����Q$Ǥm�ko�<��'I�y�0��l���jW�^f�<Q�N�h�����B/�Z DOW^�<�#\�x�R�� +khũ�Om�<�e�A'xDBB���&��eqM�<�ɗ�\Le1 뙢]��)g�\�<�k)1ZG�xcx4�T�TY�<����6N���c
*��	��A�P�<a�!��QS� ��e)Bˑ�M�<�3D�l��2w�K�G���փO�<Y�$�	9�nI؃�_�d:A	�K�<9�L� g��@BHW<��ҕ��L�<��nK<W$�Q
	�X`�
��a�<1�ۢaj�[6�8g���2u�
]�<�
����6Y�#�&^B�<aǡM��&��l�0B���K2̀v�<i��B�[))p%`�]��{d��q�<A�+�3
�hi�qaܰ�.5µ#l�<yL��&����A �,i�H5m�i�<���(�}�M��7fACV��L�<�uF�7f�������iI:�
')FM�<�BD�h���#0+�+N�`��GR�<�U��)$� �	�S��D�W�p�<QR��6~|����mZ�;]@�H�Fo�<ѣ园^�r�2EM�pӈ���^h�<R�T�LX�d(��W~6U�H]�<ّ,�.>�xhaL�Ɉ�a�X�<��N��Nx�􋀻lwL�+�aWc�<��dEQ]�s
�(�1��p�<yw�ą}�n��ġ'9��dK�q�<� �=Ѐ�èk��=����`D9�b"O�䋤-�k+Jp��\)�xzf"O����ƶ6������ʼB��C"O���&	�.!.����oӤ	a�"O��pJ]�9���A֭��0���5"OB����il��!4�(�p�h�"O��քI�Il@�dK�_� ,�"O� "�e��J�'.�F�� "O$�&�)= ƀ��b�.3�P��Q"O��Va҇/���r�<�n���"O<�h1���~�
,H )[��Y��"O�Q�v͐�5����B�5�4�(#"OB���{�l��Aʡz�<Hv"O��	����Ĩu���:�$lS�"O�!y�&��o�HaH#6@�0�"�"OR0��0����Vr��R"Ov�QW�%<E�Ad�xB�hG"Oi�{�H�A���6�Vؐq"O�9�'�L�%�@yPm�<f��u{t"OD��*� 3�F�x6M��\Xd)��"O�{&�^*[�d㠌�HF�D"ON�s��\7%Sh|�V���nl�0r"O\e	�؃6���j�G�$F{����"O(�"Ø w���rS� c�\X�1"O@�y�֫+���/�_䔂�"O ���/@�Q�	S �C(}D�"O(�'�=H���#d�5nWz ��"O��K�a߻Z����]=��	�"OLQ('2��3Ck��Def�r0"Ol ��[�.�bJ]�jf �'"O�t� ���a��ɛY�t��T"OP��G�98��,znM?k�ڱ�"OuH�h��sMұj��3"O~q	��Hu`�6���zDJ4"Ozၔ���u$�@pqiD�i@���"Oj�i�'p8D=���B?���d"O�A"YC �* Ǆ�<��$��"O��27��^�i ��\����"O���?!��L�$�K@�4Ҧ"O�H���/5}���wm3e1��C�"Ox�Q��
C=��C�L�n����U"OV����>y9���PACqy<�#"O`��"�D3���O��S��h�"OT��5��)�]HA��K�<�"O�d�E��j���4'^���R"O�d��B�:CA���o�/Xbe/x!��K�>�X�v�
tr�"T#:1�!�_�/�a����?Aȱ0QBG�0�!�$^�fk|�9�昣]�`�c!a!!��l�2�@�]�(�H��Aʠ�!�O1������Z���r��-F�!���<�W��6��s2N�>�!�1S��-���@7%�R����Z0sx!�D�*ޮl�� Q!x�0�P��k!�DY)E8�-��������<|!��߾uZQ1�LK��9���!�D�F�� BF�M�p�ڦ�Y�"�!��J#"Y��\�J��AOS
|�!���R%⌂��t�l�z�/�� !��>.��ۤ��1yL�S��; !�S�h@�쌉^{�9��.��,R!��}"l���M�Z\�A��My�!�$N�؈�c��+k�
�L��+�!�DSJ��Z2���Z��@+M�8!�� ��[ +L;8��۷�	b�� ��"Oҙ)�l34Ȣ��b��&P�g"O��P�%�L24ы�W ��"OD���/
�+�r�y�MˈET詓"ODE��mG�=�.�n_�7�"O��9���O���H&�D���t��"O^x�a0w��l�&(\<���h"O����ZtT������7T�\P`"O�Ա��CX|��H�;;�X�*"O�|A�D�Nl{� eFܺB"O0)�T�$X"��{�/��1��)�"O�,� 	�8򔫴�Wg96�|��)�Ӵk/L@�Έ%ݚ���Ś!i�B�Y�z�Z'�S���4��珍<�RB䉥J�`�hg�>R2�����y$B䉡>lܴ�u�_-�<���O�	�NB� 
�r0��!MV��1Lƌ�B�I�D�P��;���@fI�f"O 1��G��E`� B= @ի2"OH|b�C	r�liU5߸�ȶ"O\ �Ƥ(LL��C��0Ό�b"O����^J����ՆZ���)D"Of���^#Y�lLR N��9j�4��"O��X���=6,�i�Q�ٙ)�T-H�"O(Qс�ڨ�Fmp�8pl��V�	��� �"AT�n�N�#�.f
����������	�N�;$҉��..)H:�XA�x���\S�O���5��V�[(�9�o�,89x�V��J�If��|�>�u��?���E ͶV��2��Zᦅ��7�S�O�F�0���
&��y��،uD5��)���x�!h6E��'ʜ]��Q4�ϑ�y"�d�$���jIc"MϤ~�}��,��s��_6	bdKǠ�q�8��OGP���߻~��	�FG<Y�
�ȓEs5c���!?,���gLL�%��%�ȓ�(���_*Kb���f_a�~��ʓ2m��f��@kX�i1�.e��C�=hMJX���A�88�c�|C�I)u5GZ2�c��r� C�	�j� b��J�u^��v�(,��B���d`�EH��4	�C�<0� B�I�ikB�`�æ~1�ak�6N�B䉢*��Cs�p]ا�ژ��B䉋�V8�,�n-*��ֆV*B�ɮ~BtX`f�Ĺ8��:���W"B�@����t/M����&�W;~N�C�ɺ�[�K�+B�Ⱥ0)�Eq�C䉛HZhɳ"J�	�=�H!w�RB䉘[𹱷cŮ9�t�#B���ZC�ɝ������9~�(��/?PkB�ɔjl��
�f��	���Õ��'nJ�C��$":	��(R��A���C䉯V�e �� ��#5�4?B��)5x�I��K%bݴ�3��J�B�Ir/�@(AG�Abr*:O��B�	#(�m�P�U��!�t*ː<|�B�I�l�� qR\�)��mk��v~B�I�m*��u�U�o!^��r��=�BB�I�jU�ds��I�-�~W�v*�	�'��E�Ū��i'R)۵��Zh�
�'.(s�Ӑg��I
�o
��|�1
�'R���.Y��Rh������	�'�2l1��(ڥA���԰Q
�'���H�ˇ/>瘈 %FE;t���@
��� �H���re<	٣hMe �Q��"O�$��$ �yBm�HӃQ�tTq&"O�H9&c�#$$q{���j��7"O
(��L[,���c��� [Hh��F"O�<���%T5� �@L3E0t!�"O6�)S�E�==^�����%!?F�:�"O�8d(^/;��u/��}	���""OX)؅�sĞ��v.�?dKz�x�"O�XU(�b`P3.��J��5"O$<�Q F��]Ґ�������"O�,�5�ߔ�&���*RQ�*���"O��C����	�mq4�Ì}\����"O*�PE	��q �Y"4���&r�#d"OR5a���Y��D;�(OJj"OdH�Q��P�d��!.�髆"O�%X�ԟ@����a�(Z����"O���GcI<$P�+g	�n���"O.��5��jѪ<󐈐>�z�s�"O��#F�;��Q�Q290��I�"O҅��̓G���ʁ���F�z��d"OzD*�hU7'�2P ���<���9�"O���$甥muʐ�V��f�����"O���@aԉ��;�'2s��{�"O�(�$o��cV@3�JW�� �"O�86j_�)��iw����@��"O @���ӽQ9�%)1�Ñ-�x}R7"O����\�B�V����R.J���#"O��B�H	d4�+�Á=W��@90"O"��b'W�)�=����*�c�"O�@! ��
8  �eBI�Kt� ��"O�`Zc�L1�n�p�
��8$�E"OⰨc*[�i A�0J\��i�!"OZ��@B�(3DA;2�}"<��"O��Yq�%h	C�A��Hܢ=��"O�����Oj3v 2�@��K�6;�"O������g���B��<X�6�i"O��`�	�?��
֧ol�MXB"Oܜc�휧0�P(�cGM�syi�c"Ot;�ᚵWU`D�f�>�f���"OL�cF��p���_�-Ӳ5�c"O^���"]� �	�� �,�s�"O��`�$��wi\"��6J��@%"O�1{�EA�55%EV'F��"O�	s�+�/U%zU�"�H#W��Ѱ"Ox�X��H"���"�C�4)�"O�@��ɒ����3ŉ�?���#�"O.iAa��[w%Y6h�2w���*"O�Y��
�z�|z�AS*T&H��"O(h@��8>�CV!�?8��!Z�"Od�z���C]�t8�	P�0�r��F"O��C����2��T	\8}"�!s"O��*�Zmޝ��Ʈ��PR"O�SQ+�^��=��>���J�"O��1��! �1�Ƨ>�6�
�"OX\�J������Ƽk~B-	�"O(�*a�OȖ%@�cĴEi&��f"O�\�� �-ɦ�`p��;Ng�C�"O,�V�N(}inQ�u�U/-K@�X�"O�CM]/Z�J��o[8.�$2"OvI�Q%��U?�l�W/JF ��"OnyHP�R�x�kƺ ?(�˷"O2��G+Y�T�\C7��;,�]�"O$R��*x��{JZ
't0��"O����G��Pr�p���cH�I�"O� v ��F����a4�[=m����"On��1��6:�����"-�y&"OĈ�R09�tP&�=0��Y�"O�	)q�F�D�6�@�f�X��"O����(R�h��$�>1�y8�"O��i ���x:nM�ctUkA"O��a�g��b��d�$c]����&"OL����W��$�TBO�[c���"O!�R�N�&QBR!�<���d"O�#�
2]����� U�t
��H4"Ov`��F��I�t�s5 ؼܙhW"Oj�TO��<�bd�� �4�(0Z"Oޡ{�NT5馤���_2C��#�"O̽9FƱrQ �s�73,��y�"O��OJ�� ����аaC���Q"O�8{A e���еaݪe'�8�"Oh`(�BZ�qGU%��>�]r�"O(p�Gě�f=@��P�a�"O�)0�F�p��%blO.@jrģ`"O.E1���8�X��Eןe%"O"%�mӇ8.�:���F�0I"O��q�F�%n(�����r�H�٧"O��&OP5=Iθ	Fc]� �q�Q"OT=�CFl�9��a� -���`�"O8�s�CV���5?H���"Ox�IƟ2i�,�c�A�5.�Yjt"O	�ĭM�h	X���K�=y�"OfQ�a�,*���ɧW���Ӡ"O蕸�傳<�h���=.�5��"O�%����5 �N�=�BeB@"Oz�9aո;]�d W��'��TC�"O i0t���R�lBS&͝R��p��"O6)���_6Z`v��SjQ����ç"Od�y�m[�u�uz�
N�^�N�� "OH�K�G������"��IW`� �"O�4�Hܫ	�0�V�9I�@X"O((	W�)X0�L�� B�� "OB�@�Y'e�5�5"J3D'�}�D"O4قR逭h�Ȕ�&��f�b���"OB��gb����uP%�����!"Ort�'�
�.M�9�Aʃ.��JS"OH|A�o�Q!��K����~m�7"O�-����6P��`W�U��j�"Oz
!J��ؐ��.�J��"O�i�p��|jH�)U�X&6q��"O\�b#�
nq�w��;YCrH��"OV�@j:Gj�h5!��>���"O$�ʶ��V�$;$�h\��"ON�xU��:sT��g ю6_@��S"O�1�V��8�xI���O��(b"OzPZ��H�u� 	k �|���T"Oj��*M*���s�jڼ=#~��"O�x7��nt���&Mm�X�"OTp�Ej>oR8��'�k[v���"O@�� �G�����iQ3�:� "O���F�J/i����/,9��؈a"O9���+5�L��}�ZUkQ"O ��nTM��:1�;^_����"OZ!9G�M����b3�/N�"�9�"O�9��,H2+�Z�R�L�uMX�;"O�u@E�֝aSb<�r땬C>B|�a"OhQ
�g��u��,@C&e%ʠ"O���DaH��2Ɵ� �l��"O�@�� �[	��"�d�uѼ�U"O� �� �ސX��P��:�Z��2"ON� �L��X A�\!�"OXh��I�z��\z7��>B���JV"O����)4;�R�n�34����"O��I��P<jZ�Y"nY[²���"O�!�C�	l��=3c�J�#Ȝh��"O���D<f��*�kVf�@�""O`ɹ�'�;a����"Et���"O�l��%C%V^n����8Uy�$*�"O���:m�N�p�ʉ4Ds Qc"Od�x�L֩Z�2�Ǝ��5s@�l"O(-�n@�o\@3ȕiF�@�"Oh�3��^�	�Ua�m�U$$��"Ol� jD�� ��j�g�`��"Ox�8�G
�\�N��l�9vu�lb�"OJ��.��d
`�#����S�rp��"O��tGX���Ѩ�*!	v"O�-�l��N�b���Fy�q�"O6�ѱ!T17lD@A�Q�a�̩b"O"��J�-6�.��ĭt3\r"O��aI\��qGT �!8"OȘjMW�D,�0���=t�Պ�"OR�i�+a��X�@���>�~��A"O�!S�d����Q�g�����g"O~��áҧo	�E�T���L�y"O&ъq֏�¤H3f�(\�@���"ONX��R�T��恘H����"O�\b��0�� ��\���	�"Or1�Ud�9<��1i���G�<��"O����,%RP�BᇔRؒ���"O�(QEBrvR�K��D�*L�"On����Ў;3M�%�:�╉r"O"�s�' ��DŅ�
��x�"O���r���v>�{��G>]��)��"O q����(��9zT#� ���j�"O�k��ΏA}�X�C�'l���07"Oȸ�   ��   �
  �  8  �   Q)  33  h>  �I  �U  Ma  �l  ,x  ��  ��  �  A�  /�  ��  [�  �  &�  o�  ��  ��  6�  ��  ��  �  j�  ��   �
  � � &$ h* �0 �6 /= �C �I sP nW �] �d un 'u �{ �� �� �� � '� ?�  `� u�	����ZviC�'ln\�0�Fz+��ɪK*$ac�'b��R���|�ף���H8a�H��41As�9'��!��8b:$����V�,�C��?y��um��u�ă _���&�4m�T#��F�l���"_eڐB���!�%�q"ǽTӞ�"�O�mܺTr6��/]D�ݵ1�FA�S��Xa�ٶn$@��]5����'�nE
�,I-9J��$	�b�~���$�O1l�nZ
e�֙�I�|�I������$sb�1��
���xJ�۪kb��	ʟ�feV��@|�'/rn�&����Uڴ�`��������u��&�H	��?����D�O����L��9O@�D�<.P�w�� #n�GiD�'���q��QB�&<W��{�/\H��I��>��'��O��+я����
6�FF��"���BJ�?/Kdx�	��I쟸�	��	��O�n�#GH����K��bX�uJ�)I9��b�m���M;��iB�b��]oZɟ��ܴ�?	%�H+B��l�8�P���Z�P���JP�<�B-�Ą��uZư�ѡ��9F:��,��NM8����j\nZ��M��i��ħ}ݕ���HF�e"�Ly��a��4U�8��c�Ȓ�M+��0T�x�@��V��n�.�T�2JˇA��vj�v�oZQ���)��=}�X��Ә�fD�@j�nx�<n���M[U�ii66�B�>Q�}*���J�F$C7#�P��hT�e��{$��G8B1�E��C5Z�6�T�Br�UmZ��Mce�iټt��9YhMʑ��/:l,�Q̟*:�V	ױ+��hpn� !g�cՎi��Y1$�
o`I�ծ:<���\�=�b��&䔑���WYz���卼G�dm� �M��i����O~H� *C�|qxi8��'o�銰� ���Z"h��Ey�"Odѳ4U },Z��A�
PS���"Oȭ�6J<Jj�Җ.�bN���"O�� >��0.Ʊ	<���@"O�����_�&ܴ��)���0"O�$��dN���&Q� �BX2���0]��~Z�ĕ9�:܉$O�2`B�ca�N�<�A\�S �$P��L���Za��A�<�ƅ�>f��$1���.@:���C�{�<9p�O] ��k�'8r8�$�v�<�F�4m��ȫd&L�D��C'h�f�<����x��U)���J���埠{�%�S�OR	STEͼy����#�3��q�"O|Ԓ�����&Ý!����"OV�"���>�^y��h׌TX�!�"O�a�MO)[�䥛���W<�ĹR"O���"ǉ(�b͐#�P�1���!"O� �0	&u,����1".�9@v[��KD9�O��IoG�#D����)k�f�("O@L�cΊ�9�&z�eN�8�\`�"OIh�1�xMД�ЊrF,2�"O.��&��G��rgO] ��A3"O]���ېN�`ܡ��S� 4��u�'$��z��s�"�8�$%a��l[H��#�ܨ	��i�	vy"�'���'��ܙq)[BM.juL�,ET,�3�Ꝓ,Z��#ď+}��i�㋝2g:�?y�H^&_κ!̀�E�D� ���W�R9�7E�9��D�̕'tE��d����'��6�O��C�)-4�1��$��_4���o�<�ܴ)�O���^2 �t�Ca�O��r ͉��PC�.�C'��&�!��|j��'�$t�d�X,�mdԱ⮵����E�W����O&����y��
0(j�U �4�>���'ғ���H�XqN��{���?K�\l��D��$B ��Ҫ��	�E*�4i����1�,�i� �K�H2%�W;"c��p��I���%?	�|�t�.&B䀙�"�B��Rr��O�Iş܆�ɡn`�Ѯ 
�,	���Ԝ"���?yF�x$& B�G>L�q'N��J��mş�'�<ubV�O����[qm^��bN?/TA+��f�b�m�˟�	���7\ �ٗ�(O�Q�C�xS��{��'��xs�I!Mp�ѤBȤ3�Lt� j�?�1������ kc�A�g/ ��V�ea� �3�X���,O ��'�1�"�'��"[*� �@ώ>ʾ�96@�u���'������On|c�M_	���HR!��~Ul���]���ߴ*��|�O��V��rF��%T���׆�G�@Ly)�,#;v��z��rms� �a*ȽE�f|��.�	N"C�ɁD�ȍh���< ����e�>6_��0�3��H��=8L�(�a���ʼ��=+���C���ا��9Ȭ��tiJ6�)� �<D��PS�I_2�J�2*+�$@��;���ͦ5%��Ґ�^���E�0��Ն_�>pфdţmCf��IWy�'���'M�1�Fgڶ>����U�I��!��� �9{�l��;VB@�a�/f��ԓ��2�4I
�h�cB[�0�ðI��}�6��0�H�|�Uvm��3�|4��W<��O\��G�'�R���r2�].'�D��"�w����g�;���O����܇xx�5����,�|9C�"U��bB�O��q��a�XMYwb�=zP'�'��Ɂ}0�9ٴ��'����OU��N��#Z��r։�0,W����OF��
�V�qg�:��ɔi'Zl|�~��_-M��	�@����S".
;���Ә_x��zV�P�R�D
6o�<4�D�?]����a���!e�u~K��:?��C�ܟl��l�O��k��8@V��k�h�#�0d!�����fj��$��/��2��D@�O{`Q�¡��dԺD��IP���iW�V���gI�?i�	ڟ���~yr��`���C��9o d��JxK�A���(��t9���.s�r��F�i*��J�<Ά�
��fb 9㰃_rz`�k���`>d��5�W+7T !V�i:�Ă�>��e�IH�)grȡs[2�����C��O����O:�̋Tƅ3j� �P m�Cw
��#	o�<��
�+�0�EO/n�:!`�EyR� ��|�����ݼB7�M�a�n�
��$+(hhq��O����O����<�|���I�L���"Ϡ@�|'��q_��@��{K�\�rcŏX���4��m2�B #D��+!��eE�D#'�42�LAqOV�%����Do�'��@x2�0lAŉ�j`����G�8�?���?������I``�B�@�r�����LC�B�	T�[#g��XôH�IK$k�R�OJ�m�֟Ȕ'?LH4�-�)N*w��`x���0$���垶R�[����ן��I+{�A��%�[���D+����1���M����\�`�PQ����4��O�q*p�bNN�
�4�����A�%�0���O��؊���k",�?Q��֟���O~R�� 2�A��K8R���QoV����?�	�l{P�� p��Cځ:(�!��G���;�t��4$(?劝�â��sX����Wy"�v�r�'/�^>ٳ�����X�0��^�l�P���-�� Vcğ���ma֔���QvՉ�&�?�O(���R��܀�����Z�r(9)q��$�p!T�!%:�s�FА.S@F���S�9p�3��I�m�.4�Q��'���	�*���'��>}ϓE��]�׋�?N>X�r$��%0���u�����F݊�~������ �F��0ڧg�������t;l�(�bMR��$r�4�?����?DFJ�.!2����?	��?i�w^��Tđ�}vB`��D�~g*�*�y�H	��0=��AX`
�hR	�o���C@Z̓N�| ��I>Q���y�h�H�P��#�S ��O����<0���0�<�Oo�,���
�E��1�d*S�@$X�'��dz%�خ�ɢ�SHJe�/O�iDz�Ou��������C.���ȗz�p� �O,���O8���O���KǺ#���?q��m!��ag�-sy|E�S�5j~@a�S�_ L3��S�=x��(��'T��2�N�r``]ñ=�~ͱ��O�$��9��Z����Ң�[�	�џ�rd�]���JІ�<c@>P�ag����D���ߴ�?�(O���6�/�IY�	zlВ���GU0���Z���H&�Jƶ̉fGZ�Ԕ'I��e�X�D&�9O��{��f�4@h6!�s��&|źa�$D�p�����3(]M�Da�sH'D�@��K)����e��~�։;�:D�c2-�;"�2��tFF8c����W�7D���eZ	�]��o�8�^��%A5D��BeQ�U1^�D-ľs�fm��0ړ<@��D�4����RA�����_�-�Tl��yR�/)��L�B������;�yR�6 ��9��Wޅ0>త3	�'�h�'\�Hd�Q5�ԆA�	�'[
���J��y���Ju��n���Q�'���&M�W�؀�"�>l.��t�,�Dx���Bh]��s���8���jӢI�:B�	�x*4)I���-1��2�U:�B�	���X̜���O�"���c�"O��#f"N�Z�I#��z�����"Ot��!��FIv�q��B�D�a��"Oh�Fd��P��B1��O?rU:u_�\���:�O���ΉcFa��(�b/2젆"O� ��P�hY�!����r(ÏZ�(1"O&ْ���	��}��(�TmZv"O��e�M)Z��́`�֒�h�#�"O�U�b�E�=B ����Y�Ueb�F�'����'�ȓcd��y$�Bٹ09N���'�r]��ܬ2U���vW�.�vL1�'��!ᦌ%#��PfĐ. ��Ē�'�T)��&K�p��1�MX�iF5��'u�����͖�V�Ţ¨�`ݳ�'4�
�ִ#Ԫ��Y�8D������2zMQ?mU�՚aY���F�����(D�,�b^�����]%P�l<i��:D��k�m��a�a�[�5�j�Re:D���1�Jr�>xG�X�_;�Ac�+-D��8�-`�LA%(�t�6�	h5D���j�+���H�-ιCN���e�OHAJU�)�-:}2�̡4� ehd"X�0C`���'T���q9�-�d�+6��'x��Hw@V�i�|P��B��Y��''�Jr�C�2������!Z�Ej�'�Z-"f�L�up��+�B<��'|�\�P�B*D�b�"uÅ�01��H/O� p��'"@�"����;4HϙE�ٓ�'xb�IC#��&5�� ���� �'�R��6ɛ�v��)�`m��*)��'�>�B���xX�*AE��yd=�	�'���&�#:k܁��������y 2���X���0�&LT�h�c��S� ���3�D�2��@E% �(HU���ȓ�A���K�
b�# M�,��i��K*49qs@B�+��MAI�*�V$��V�!@s�ݤ"���!��[I��P������e-�
yWϑ�t���F{�$��ͨ�0�;B�3R�&\����\4�IR�"O4-�5���Ni�0$�e+|=9�"O�`�E���R���]#��02"O,���$�J<L�� �?D@���E"O>��F6+Ś��Ή�|>$i�"O�`�ӇS��șpc)S��u�'�ĀÊ��Ӗzܰ�p)��k��SD�899r��DJ��w$Kg���83�ٻ6�}��;zd\���ň3�f���m�	8D��%��	���N0!碟>AD�ȓԦ�0hS�v�B0"��_Lwji��. �I��l��"���qV��4	$�0�'5t=��ub�"Q-�.ޒ˗lA<09v=�ȓlL3W��I��� ��6����!p�ݪ����iW�Ց㐼6o��ȓ-[�;�A�1����S�(�H}�ȓ_?�x�����QQ4"�P��	�l���ɠT-�Yp&�4�z���䂱'�BC�	�n�z%��s�n�{V*9�
C�I�I�H��i��vd0���Ā��B�I3^��aU%�-V�^�����t��B��t=����?|75ʆ�/�B�I,f
�1�п?7�8`�)$�l�=I�dF}�O�~�7��?t������.�~���'\DaS�(	�Rx���Q<$
���'���(�'��L���1�J����'RZ̲�>%-�J+W=� ��'����1��G pӀ%�$T��Ż�'�{TKR'@��K���M���8JڈEx���Q�S�\�{V
�R!*��#ѰKIxB�I0�
Y���3¸K��>�FB�)� �]�w!��{:�)D@�ֹ�1"O�\i�nF�~��)���J^�Jh�"O�[��T�J<~����>b��l:F"O|aq$��*P@�1��N6���R����(;�O�\�e֠8ȹ��]u�8xf"O��70� K%Y9!hb%�s"O<���-�P����c^�RJ6@`�"O(�H���<�
#� *1>�!"O�Q�`d��J�	X���SK�����'�\%3�'l��@�X�]��:R�Ø%:��#�' �\��A�<�������8��'A
99砊}�@pI���X���
�'��l;u�?Y'��#6-ƮG�2�	�'���C�ˏ[�X�(� �A|��2�'=D��R�B�_�l aBL
�	��a��D��.Q?����tX��٧bJ>1Y6)5�;D��۷�U�!���6~.<9�&$D��JR!��I��F�$2#�-D��jOO,��"	�&,��B",D�4�L��Tn��Z h�Z�LX $.D��A�.Ǯ@x,�*� +#(�����O��s�)����2R/���p�Wҥs^��3�' 2d�C�H�P�l1!��|��!	�'u�����#��tZ���d�+�')6is��yrN�b��@�w�T�*�'N�#��F$��`"W�u?�s
�'�FA`ɇ�.�6$⠈Zs*�*ODQ g�'M�}��A��;a�L�q�4	�'�0�j��J�
)� +�eˬ��	�'�<�)�
H��X�cȈ��ĺ	�'��!�$�
�]�K�OG/�^<�	�'��PÀ�U�ډ�ŏC�vN�Z
�	��t�q��� t�ҥ�JG�N�:l��q� ���ۜ#Ҩ�:�&�8������}��hc���L�2���?~~!�d�!g�JH{�	Y�<PHr��-6`!򄔠k������;��� ن~g!�$5)����%V52i�'@_ў�z��2�!�Έ��[�]Ɉ���d����m�ȓm�d���K�`��S����Y��kT����Ύ�/�NY�W�H��q��^LQTBN�M�����F
6��ȓH�I�I��&t�H
p!��kʙ�ȓ`�6d-I��e�v�1W�z�ȷ��OLIH��)�,���
�.żFP�L����s�s�'�
 �W��"6,�����4��
�'B�xc��xc�`� p>҅�
�' ���ai[b蘐���oX�لʓ"t)�d�3D�"ɪ��dz �ȓ_�v&��(���Tk�$D|�E�'	\����1D��°�ՈҡX� ���@�lE S�ȡR��P"�U� �Ņȓ���{�	ғvU~��яX	h�ن�%$>uKV&V�C��除���b��}�ȓ
���)R)G-^\���I5&��9����Y6�I�|�Z���j�q�IS�)�+�C�1C�T��`Ue �]�ծ��q��B�I%�3D�RV�L7=�q�!l)D� ��$pɢ5c���r.����D&D�\*�ۥy�"D�Ƭ�e���! F9D��#��V�@��� ���8CK�a��B6ړ&v�G��S�.�P��d���fT4h�3D��F��`�rb�?J�E)j2D�l��_�W��*�$�		��I(wK1D�� F�����
E�DSu
�N�J|["O^RԽ2�t�K2��!�F�0"O�tɲ��f��
N-��%� �'$������Ӷs�����e��Gk�TZ�aÙ�\���)��-r"�G`3jmA�m��4j"E�ȓV�9#$��G��UQA�ܨG�*T�ȓ9�օ���!)����aE=b��ȓO$!�s�J�%qܑ�1@=�PB�I����mͥu�D B��:\��Jh(����a<5�@lX9>x�(S>+�C�	5L���oF�>�^��R��Z�PC�7w�<�"fX�0'P���nJ��B�I�u��m�s�@i;H�!��k��B��YB��e�s@�銶�R���۹x��D�
y���*siB�~�䡣CW�[T!�0u�z��G���F�<��f(4!�D����lzGk��_�R�b@B�st!��^���ԅ�$l�\���*Df!�d�}��B��2bm�`�Mr!�ǳN�9:q`A�d�^��3���ўC,�I�����",��Pb$M06��ȓBb��v/ң7! ,Zӈ0X��h�ȓ.�����Y��r�H�)	@B%�ȓvC�9�7OٹX�P��f�B�"��ȓ�$�!rj_�g���&E-8>�l�ȓ%�(`��	T�J�xs*E�?6\��I~�#<E��ȟ0[��9�E$X9=zлg�Ǖi(!��Ƭ�"ٺ1n
z	L����A�kt!�dУ.�JI���^�s�6=�/.!�d%��pR���1n͞���3k�!�D�]�ib�Q��J���	6C��d6��4�7�P�K��p;��?GP�O?��5���qwb �	�z^��O��p"X�h��ٱF�L[�.p�Ǵ<����?��[��LA��<I���F�; <���O��x���	f)�BEO�,{�}a����UXą 1��	'1jX s�C�����]�W�j�J���:|f�'&W�C�����*�O���*�'O�sR�, `�Lzg슃|���0?aP�ɸ	�6��e�{i�h9�L�ox���/OX ��)��|�@����A�LHn!�[�h��ڟ�BrOjy�\>e�S���W� ����Iՙg�,��OޟċRgW�L�!H�Ň�
��Y����h����D�ҍ����C�J��l<O�aY�k�Y>���F��-�j�PW ?ڧ. Q����=8�e:�f�E�6t�(K�������'��d׀.2�M�E%Q��p����!�ݪz�&�������0H	�j�'W."���'W����I�~��1�ͮ.g���-O�]���Od���Ob�ĺ<�[ЖH#��n�衸VOH�)���0����X�Ek_�X��Ql����	;��0n0����2v�ip&K O8����Q�\�|!X �TP2n��g,"�B�L7dy��	7l�_BR���F�����/�R�'cў�͓&��9�ԥg�����O*D�x�fC�RNJ��u%�1m����7�O*�Dz�O�P��
;)����iU�,A����J>0������0��򟠗��O�`�a�G�?��5娒y�`h�I�&@��	s�Tu��ؔ�L���?��J�gC�:��&w��Ѡ(��$@�ş� qJ�{�N�#"�������G���M��D@|���H��<���b�'\|I1�E�-b�1u�D��
�'I�	  ����15�ެ,7\�*O�yl���'`Fle�#�S�J���1�� r�TQ:�D"|�x�'�R�'�⬘���p�O>q��qpr�9;����� �\��%N@-8.ni*uM�1����@�V%����c�5{�r�9��Z�?I�/��n���q��ؔV�E�6�
��e�Iߟ��|�V��&a�l�R�U����U�Ӻ���?�OD��@���>�>��$�.v�ޠ*��'b �~��aP6 �iȟ;�(!�'<T���m����O��'*R�����?��T7�J���$�a3.8p��ҥ�?�CN٠X!��`U��]p��*�#X�ڄ��p��r�	^�^��J�C��nE���n��
��s��|�VLX�;�|�K7/��H�NP!ՇC:)p�9�0�֍O�AR8O6��2�'�"����,�S�? ��2oP�i^����	�>'|��d"O�T��&�,V�*����O|����	4�ȟ�t��7�JE�ѯy���R��O�d�O�8�u :QE����O6���O��;�?�`��xƄ�rem���b��bB]�'�`U��'�0`S�[�@�5Rɟ��1��ɋb<� �A�|<X���NeD �	�0��T��a�Y$�g�'� x ��~lE��$NЬ�{�OԊ��'���'�O��'(#Hi��a���~X��Iq�C�I�M�j)K���/	fT�ň�?|��DIM�����'d�	��PŊ≉B�ܼY�'�n�p�c�2?ٞ��	ߟ���ş�^w'�'�˗\�x1y��j��-���\�u�����ȕ,4���tHP�P� 1��I�h����
�ę�$"�Qܔ��Wmĺ锸����0xV����v�-��8m�8�"��.�Z-�"�y��Y�I����?�����/.f���5���;�9'�>��B�"�x�id�D���0���x��b����'g�'Ƅ7��O���{��@�A�yZ�Q�&2��\����OtY�!�O��d�O��!�g�7k@PD��>ي�mZ�|:��ߣ]&$�&b��BX"Z�'ӌmz�o�9M��d�a�ś5&�|kP�O9`��t�\��]�g�i|�����dG�5��m~�t!m��� �'H~��J�P��ě��F1t2)�I�tE{r���!v;���ѩ;.�n@3�i��ch~���JC}�ZJ��R�P+h�`�r�	óI<�'�B�':�	u����H3�)ʤV4�!��� +e����>���D2�L�>���(�	��q�i�#���?Y$�B�	x�'v=T(i�݇ ��ȱ''�7G�h�' ���GJӧ�9O<��QM	OC\x�6�3)�� �n�9g���f��t;>�O�'>5 �]=/�u�Q*�	Z�����Y-���$8��<W-�X�8{p�و&�؄�F(�)A�@��O�եOdy�>�P?�����z`��� ��s8�+�#�O T���>���G`�OĨ�O�'y��0�(����'�d}jH�,�L��S@#?}��h�^�s��T�u�B�+A)л	n|�Q�W��ZO;}R�4�ykZ��B�ˊks с��W�@%�W�OLp��>��yr����d�d�ȝ��
fO� z�b�.gS��BN��i�B%?��,�'5ݬy���!G�hIA�N}L<�	'���) w�)�#����r�Q塕4}� ���>&t�	�R	aR&@"y܂�@�
��2�h���y�m�>������6C���QmK/�M����?�.Ox�$�O�ʓ�?���[v����0��Jܙn�l���ަ���ǟ��'��[�b>7mdH�m֠J��Î�uZ!�D�;{�����#�
|��)���vL����㉰r��s$�/,Zv+Z3~VB�	�5�ZG�ȲW� kB�!(nvC�I�G���SF� XR�� EeY�r'�B�ɞ�Nx`E��p�����E׺(rB��:#(�m��
vH*m�Y��C�=rKvBǤ�����v)P:&��C�	�TT���(�f%6-�3%N�zy�C�ɯmZ�I����2.͋���pC䉆NpjQtÍ1i�H��Ba0�#?����?q��?	���j�IU.ؒX������	IHYHu�i�B�'�"�'�B�'���'�r�'��ћ���{+,�`���;�� ǩzӀ�D�O����O����O����O��D�O���g_]�28�͆�C�����V����	ǟ���ן��I���	˟H�������V/�!��j��;��)[���?�M����?)���?!���?���?����?a�e�kޠ,��`ыoD����V
=����'�'���'���'"�'d�ۆq� )���{�fpP��}i�7��O���O��d�O��D�OL�$�O���-��qI�1����gR3
eo�ٟ �	ޟt����`��۟�	ǟ��	�9*�e@ѪEʅ!!i�L�sݴ�?���?���?a���?	���?�������̧m���J5hC,C�ެ�A�i���'�2�',b�'�2�'���'�8��Bl�mU:�w`͛��{�*zӞ��O ��O&�D�O����OV���O�-�#��%sѴ���ɋpfe�c���q��ן(���X�I�� ��՟��������,�@`P�ǟ%�lj����M����?���?	��?Q���?���?I�噚<qY���+� T�凩�EDq~B�'^�	F�O�L4���V�ȭBU��QD�i@P�i�"�Èy��ɜԦ}͓?�l�e�ǲAJ s$��%B���Ɵx���$7�	�(�6m��Pja��24�(Mkv��&D��K�OR�4�?9�`$��|Z�'F
�µ��,���ء���3�����2���I��C!�	n�? 4Q`�V�0i�X$����r	����K}��')r9OZʧGv�ɣ�H���"h(0�ҵ�'|B����J�O󉘡�?��u��AA�_V�� �b�T��>�po�<�+O<�D!�g?!��	�a��4[��(]J�@�)Oğ��ߴ
���'T$6m5�i>�Bv��"��SD��"-@��x�K���	�x�I�TZ�np~"9����ẳ�E	O���I�T;}	��q�`^�'yRR���|�3�D�P-f�S��w����J�Ny��k�hӆ��?�=C%6f���5��5Q%�0Ir���d�O,�$k�HF��@�<&���!��[�@�٦O�t@��b�ߝ����O�(K�;㦒O��)�Nx�)�P��Մ^�r�48Q��?y��?Y���?.Oz�mڸM���	�V��A�e盉%��-���f]�	��M��m�>Y��?��'�)2���t��HF��>�.��3dӶ�M��O4 jJ�����)4��cޝ�1�I�C��	EJX}�;�m�O�B��TlX��LZ4�Ǯ٪#N���O����ަՋ��q�TCjӪb��(�#��j�%���1�Ψ��6���O����O��$�k��Ӻ����p���k� e؇��@ш���^��O�ʓ�O"\sA�[��3��5�dI;ĦQ���'ж6m��.��d�O��0�/]�X�9��?	��$�"j\Oy�"�<����M2�|ʟ��cԩE7�
�kBA�U��)��FP�� A���F^�	�?)���'�U$�8��	�,g�RABː<�|9q�ҟ8�I����؟4$?�'Z�6M��H��eŀ/j�"5�!g�; ���b���O��Ʀ��?��P�\��4vR$���J�G�� �g����`w�i3t6�ڂ)K�6�1?���Y�H���I���)�6����@E�%9,�q�Cyi9����OB�D�O���OF��%�p��=U��
`��o�4�G���M�%N5�?Q���?�O~Z�D�v?OJ�s�d_(?e(=�W�!oզ����t�P�oZ�����'D��4�~Bˍ�m;��`0�T���C����2ٴo;��� ��O��KN>�(O���O����0t�x �N�^j p��O����O��Ĳ<�u�in�A��'�B�'�l�X�DU�c`�t��1����Q~}�hu�F)lZ��ē&{���#NERl�!k]�kr�Z-O`���ѕQ`�ih����%+��c��<�Q��3Ű��w�
^@��sj��`�	̟��I���F��:O�,iuC}�d��!'Hn�"��q�'kz6M��25����O��mX���s	)Q,(�q�P85�X�	�*�y��'���b��٠��r���5�Y�	����%�0���@�'	`�L�v����O���?q��?Q��?��W���D)���k3��.f��e#-O�(oZ�9v9���D�ID���`Fc���1AC�Bl�W�ҥ���Yڦ%��4u≧�O3j(�ϴx��� �gǕm.�bA6=��X��^��P����2-�h��Oy2��;r��"H��5_>(+RO\t��'���'�"�'/��MӦ�.�?aq�F%xXm+A�L���2��¾�?�i'�O���'r*7͜�ݨ�o7��Pr�е69��3�G$P�� `�����'�@ɀ"��?I(ԙ��2�VZ'C�O��[uf��w�@2�'3B�'_2�'B�'�>ISIW?c� �d��~�rycs�O|�D�O��mZ?�Ω����ڴ��'9��0�Z?u��9�KUB�)뷓|»i2�6����Z�Le�x�	Ɵ��!�j�^�
�V��X([`$��*���'�l�$��'/�'���'���k��x`j�h6��H�0r�'�U��ܴ�n1���?q���� 	3L�K�NԌY䧊�c���*����OX��)��~�C��3���qDŻV ����28��8��@3Mԝ�'����o9m�u��'l�R�#�8xUE�cR��"�'�r6�ӇyV�]z�GP���G�s2*j`�O���Ϧ��?�R����<�Hu3�C�>���aU�D�\n���M�7f��M��OD}�ǀ�:�!<
t, (�&)�t%�oD�(�үRڟ�'�a|��ĳz��Ee��-xIAڛ֬N-(��'O���ᦍ͓k� �hL�`�VD�3n7/��i���H&�h%?1q��XҦ���_���9��ۨ-+t�bBH��YQ���	�cT�����'�T|$�ܖ'��'9Z��3�"K�M�DJO,-r�@B��'�2�'�bS�|;ڴh�x�,O��d�M!�M�h��*"���Iʢ�l�O��d�O�O���'�'<{,����0�d}�M�<�d��<�m��mG��'4��$F��yb�غ}Ŕ*�e�#6nmA�#��?����?)��?���e���6%��F�B�!�N�-\ڊ��\A"+r��9��O���ئ��?�'_bA�v�Re��RM�&���_����lӨPoڱ5>�oT~��+4�m�S麫Ԡ�1[���Ԍ>0m�� ^�My��'H�' ��'o����@{oVU~�S���W=��)�Ms&��2�?���?�O~���o�V�	@��֔T�B㆞i-�ې[�hjܴ}5�v�%��i�Dk�x31	�sRJ=+Q�;n�L� ��7��	�w`pi�d�'&F%%�`�'H�\B��!�J�b���-^��R��'6��'"�'�P�4��4E�-C��� �)�$KZ+,O�@�]/��;��'��7�(��/����O0��q��r�c5���a朩t��yb'LF�}@�7�9?��ɖ�c���	L����y'�ZA6&Q#"��"�&�JwE�?���?���?A��?���)6^Sȥ�5�&<X1DE߅<�R�'n"$e����'�O��Ą��<	��͆K����J/��c�ȕc�Iϟ��	㟰�3N]ΦU�uW����h�w�_.6��P��o$����'���'���'���'6R�'����G�;+k&����Z!�qg�'j�U�؁�47�^�r���?������Y�n(��Ջͨ>%��"�B�PR�	>���Od��"�4���$�9e��� @)t�b�ˍk� JQ��Jh^ R�N�<1�' �$�P���")h|s�ޒw�Xxp��_/DM��B���?I���?���䧔�$�Ǧ9{bF'DɄ��<u]���@)�?h�`|�	ԟ���4��'���oћ�ˊ3'�V�̎^�	K�j�+_�6�Z¦ݨ0GY�%�'�t���?KB�?� ��	�L�$��@�3�|A�v��O�ʓ�?y��?���?�����i�$�����2 ����+��	��7Mњ)����?AO~�|/��>O� �D��"�ƨ��5D���'�B�|�����U�<՛�O�Ш��N�{H��I&�E,G�Q ��'켻�ޟ�B�|�U�<����d���A~5`m�f��%��d���ퟐ�Iӟ��ISy2gy��-	�m�<�����(+3lA!K�0k�$P���y�RN�>)��?yL>)C��o��U	���#m����dL�J|)�2�?�B��P!�����IkFpQ�SU�HIB�:"�ى5��B�I�s����ܯ	L�(��+
?���ͦ}+��ȟX����Ms�2�O��=x�'�;#�X���0=򄼃Q�'�b�'����_�����]&=怠�S�g�r�x@�Y�*���I�Mί{4ș��|�]���ɓ}���'[�%U�����Bn^>�G~�֮F��'f��;�<4I𭗺vh�12ad�@��'�B�'ɧ�OJ�Did(S3Z��ͫb%ur@�Ε"�2�S]�pȡ�>V�Ҍg�y҉�6����Uh�<0Q ���v��'�B�'��'����Mۀ�H;�?q���3�R	�%�L/�:1��怭�?r�i��OD�'>7-�ۦ�J�X����XX����m��W]Li!� ����?�꘩[�4�iױ����X�ݓ,��t���?��1F��1��$�O���O~���O���$�'ތx!�NF��ܩqFԣ`�e�	ן�����M�b��?�����\#60����7tT(�h"��k��O(Ylں�M��'N 0�4�y"�'���`�b�f�<���@��X����>\�ɝ?��';�i>��I��(���AEDUJG��� Z� ���9�	�p�'�|6���L�d�O�$>�wa����R���Ky��Aw��Sy�>�i��7�O�i>Q�S-t����(N.s�� pqO�z�@�Q(`��3g�4?y�'^�0�Dܩ��_F��붫_��`�rDP4�������?����?Q���?A���?1(O��mZ���а7�Ŧq�8�S�F�G�B*�k̟h��)�MkK>��r��	؟@���W'^��@�d �vW �Qb̟���4g��a�4�y�'�z�ӷ`A�?u��\�t�cɂ�ǆA����#f4A�՟d�'#��'��'�'�Ә%�u[GF�(8 �kbjG� Qm���� �R��ş��I�?}�ßP�I��M��O� )x� ��]�z�Z�߭��#��i��D9�쟼���@Ԛ�l�p�ɣ,*`�C�դ-)^y�1�Y�x'ʱ�	:T�Pi�2�'I�Q$�d�'��'��D�!�ыfDȴxf9@�H��'Sb�'�(�k$P��ݴ?��8����?��*�*�X��\�0�xQj��c�6�O>q��~��	��<�	i��s�^p���D���ˁ�B3!J����O͐� �J�4C���<a�'�&�D�"�y���?�*|�f@-�USw@L��?q��?Y���?i���{�p��d�hɡ�&	���%b3��O&m�\��4�I󟠺�4�����`}�1*��GS�D�Ѐ'*L%� �	3�M�p�'���З"G�f���� $��M/�t����pR�* �6�R#2�Ɣ$�Ė'$R�'���'���'XdM�E�	~��hA@ɜ>�HtCW��k�4|���,O2�$7�i�O��9���1);|�3�>r��`�Щ�\}��'��|���bȿ�lE��l��s����S���rP2�#��ֆ��ɕd�٤�'b,'��'ʐ5r� �C��с�@_�n�j���'y��'>�'��S��i޴r/��'���c�֥!���0��)Cˬ�s�b��V�$P`}b�'�<O,<0��y6 ��@$�eH�bȗ)V�6����6$ 
���c^V�S�[q�I�ZX	�D͆#84��J�ݟ��ǟ��	��0�I��D� J3|��@+�Ha��p�2���?����?���i�|7�'��p�*c���Fm?6�6��A�]������|≺�Ms'�i���m� eɛ�����w�Z�,�H#o]<q�q��)�9+s����'���'�������'���'��(�kV����ܕ<<���'�"S����4S���'���?0$�H 8��e�ucC�O~� �<��T���	�%��O�bɑE<�b�'�L�Y� �c�kM4Ƹ�o�0����� � �����O�mZTk@�&�+���4#���?����?���������� :�j���4��Y#,U�=��8���?&���'�~7�8�I���$�O0�/�
P�j����7rAX�M�O�ݒ47M6?�;}�B�:�'r��'~�1ɔ)�7�4xC5�������Sy��'\"�'"�'�?�YW�R:=2!��ٸ3���Lצ�)��A�0��П�$?=�I��M��'}�)hef��(�t��d�[��'7��|J~�g��MC�'V�F��x�4�3d�H94YNu �jT� ���O��I>�/O@���O(���.��lf�a�5���}��,����O ���O��D�<�ֺi󨈓��'��'��P%�V�֤4e�Z�$���]y�'j��|Rb� H,�-��g�O.�J%�Ơ�?��`xRp�sjƯbxy)O��	��?�1�l�\�IxsZ y�d��]=���&�����ܟ����F�t<O]cv�'&��4c&o�>e�q���'��7��.N�����O�qnh���uJ�$-��X�c�%m:����Y��?у�i�v��m�Y2�eӤ�$lN������ I��k�?N\A�Fܨg�0x�AM�����d�Ob�d�O��D�O���H<BdV�衣^r$�-#`,L��Q�v*ʔc%R�'&��d�'n��I�+E�2:U�7��Mf\�����>����?!K>�|���)��A�g#�k��r
ޑ-
��$k���)UG� ���p�O��{b�z�A�95�1���q)���?���?���?�+O$�nZ�}��p�x�||@RGD���!��M�Jk2����M��2�>A�i�(7�G�����$^�NT��)���P�Y&�@�_LP6�(?a�玘;��	5��ɼ��䇺F�b��2G��]RfDІ�꟬�����	͟����G��h�8J�y�b�C�|�!�v���D�O�,mZ�^�x��ܟh��4��'��U��$\�*s��z��ȵ�8�*M>y���?9��U� �z�4����lU;�MO�%'�	3�&� &e��"b���$��������O���O���J�`�����9	�`��������OR˓ �V�%i���'�"�?)�#�
2d�X��Ի<��3�˨<� X���ɟT%��ݟh�;��A�ddI)_|nܻ��Q� m��҂JL��'P�� ��YD�|�ܧ(��	�pA�}�a;�OX�f��'4��'�R��X�H�޴=��YY`��Bf4��M�_��h�"ӕ�?!�k��6�d�f}��'����"��A��qs��W��ę��'��n.���6O ��A���SW��	�@'t!�'� H�c�
��W����	cy��'���'���'���?y{7��#��i�O��k<JJAM����۟|�Iʟ�$?y�	�M��'�,�J�)ݹ#�T�����gP�+žii:7�HD�II�ӓto�(m�K?7�5b���4YyAxTA^̟hP��P�l��G�V�Iy��'cRß&�ڜ9V������0��'���':�6�M��
�?���?ID�D�@����]�Uޒ����Y��'SR˓�?iڴT��'LXE���_x&m��K˗3>�b-Ov�I���8Cr�X��<��@��?qħu�0�ɝX�h��|��b ��DO��'f�'2���<Ac
/�8S"@>`0�Kџ�I�4g¶����?i�i�O���Ϸ����	U����+5�$]��Y�۴n%���T�#Лv��d+a�׹k����(9�,q�U@�Y``�ǲ!s^�K>�)O���O���O���O��-j^MC3N�1|$��n�<�G�i��Y�V�'h��'���!ǁm�剭0�b4Yu�66LnxѲf\(|P\)+O��d�O��O���O���O˦<-RaM�*U����*�`�$��PX�	��6 ��' BE$�(�'��H1`F�6�,�a��{N\�V�'V��'���'2rQ���ٴ[� m���
���!�
,J���:RȔ��>����$�`}��'�"2OJ��ć<:
����� c��!`Pʃ�[ۛF��d:&��S�����P���T�S�)F,�p�W17%�T���柀��ҟ�I��l�	hy��Ԭ�V!$����
 G&��bɐ!�?a���?��i��1dY>i�ݴ�'� �WiP�C�]F&":�L�1��|R�'��F�O\x���i��	�\�������*�('��FΖ��@�=x���B^��|y��'���'��O�3	;�E�q�	0$�tkƇ�1z�B�'��Ɋ�M��/����O��$�ȍؔ��k�������K�T|�'M��M���	i�Bd&��O�Ф2fB �f%&�#��\����M^*1@=pU������L�8��I;
�OD���ȡe�$�r�o�u�G�O��D�O����O@���˓{ƛ��[6)1����%DJ��"�	ێ0����2�']B�i�.㟄êO0�m�,1�R�NO:S��Ԅ¢EV�=۴}U�
�:!��F�����Gϖ;T���Bp�ԯв#3��`f�B=����ʩ�?*O��d�O����O����O��0��$AƦZ�n|�(�UXSd�M�ڴXh$U����?	����'�?A�iD��ݍgG�ò�]*\��p�%��R��7��ݦe`O<9���B�'xvxE�ٴ�yrd�/GQ��TD�=Z�����	��R��K_b<�	�T�'[�I՟����\棂7(���qD ,n� �Iܟ���џȔ'&�7-#kۈ���O����>���gƷ?���Arn'q��⟘P,O���{Ӭ�%����#��M�)a6��%��h�Ϧ<i��ʜU�x@A�Y��X�v��Y��yR+�PϠ����J[Q B��?����?���?���id�� �-KmG�>���[N�%l��`�D�'�6���	�����O�To�a��2��'n�qI2�˛`}v �uā��?y�i)D7m�ߦɡ�&�٦A�'�����H�?5�RF�+��Q��"2}�h�.U�DؓO>�-O����O��D�O��D�OH�x���>A��1�Ъ�8�Z��v�<���i�X����'4�'��O6�A�hX��k���%��Q��#B�d���?�����|����?)���'�I
�(�	��%Sf7U�bl�@N����DL��xͲ�lR��O|˓0=��8���/�h����t������?����?A��?�/O�el���!�	?�Έ�����&�ƮU+�v	����M���"�>����?�'A����oX\nq���9s0Z|3R-3�Mk�'��
Ɲo�� �S���I�?�ϻ�����lWZ��[#G�<�`��I͟\���$�	��<��T�O�LK`R�MG �@���Uo�����?��k����^ >'��'ޢ6�;�I!{aj���"ĀJ����=L�ԒO^���OL�dߚyx�6�l� �'VaByZK�]�pEq�ĉ"\�@ �� '�?�E*>�Ġ<����?���?�'%˸uY 8;Щ�J���C� �?A����d�æ	K�@��I���Oy�Ցs�4�6,[�-"���(O�(�'��'pɧ���'<B(:ЭS�B�Q�#+��"|ɑ%�<�I��\����?��W�'Tp�&��hd�(V`*����-H��kVJ�ݟ�Iҟ��I��T%?M�'t7����}j��q�F�r��۪�v�0CH�O�d]�a�?qu[������ذJ��4�|�:�&ʪ���	��,õ���E�uO��5��t&�x��ꄉ	�Л�B�&QX&�CC��?�(OF��O���O��D�<�'L�N����ܷj'�A��	���zݴE�Z�����?������?鐳i��B,\��I/���Y�χ�MU��'��'5�O�YԹi[�D��l���BdmX�=X|�{��\&J-��;Dǂ��	�G��'�����<�I�mb~ѣA�U:7�P��Я	8.!(�����L�Iǟp�'�6m��b)>�d�OH���?�HQ ��8kvh)%,Q:� �0�OHm��M���xB��$
�0`+Ib�,!aHc��ɁE$�Ht�:,��|*���Op�;S��f�$
�5pa4-�XM�	ߟ���Ɵ��	m�O��D�9]����� �z�Sr+��2`ӈ��So�Ol��)�?i�'o�}0p�W�d�(�k� \��x�Cƛ�"|���n�,+ߜ l�w~2.W6x_� ���~�B�	�r�n�~:�,��⅀�����Oz�$�O����O��DW$����d��F�����9S��be�V%Mt"��'�����'Ψ\����Zܐ�(bMȴZ(6�qG�>ᣴiv�6��F�)擘E��1)��n0���RCGy�2�1��K�2�Z��d�s�O`�jI>�+OXl�%�[�Wϼ%!@��7��t���O����O"���O0���<1·i��uJ��'�4t����y́ASeƈ'Ԙ;1�'F�6�!�ɀ����̦X۴� R�g��@�P�)�Դc�B�1�P�ݴ��A�F5�(���D3Ē���}E����F � gő)~������?���?q���?1�����ǀ*�0:B�:�T4�G�'vr�'�T6�٢Y�����O9n�|�1s����Q�]��t� �GwM K<	&�i(7-�rL�T�g�:�
b�	��@��~�f�a���<�Ȑɍ
��֝������O����O��$�)w��ѫ%m�b� ��FA��U��D�OHʓ*�� �Y�b�'��?��I�&Q�i���H���E��"�<��T���޴8���'3�~r����z�:�p�E�J��+r��5'�����_Е'���"���hQ�|����Q��T�_"����	�(���'�b�'�����]�8�ݴZ�D�I�&�Y���bf@�U�@$*u���?���B����A}R�b�V��@O#�z���F��w�*�ٵ��ͦ��ڴu�V���4����n�F���'u���dϮ�K6kqQL*�(��w�\�	|y2�'���'�"�'���?]hg��6C��=���09C��AjȦ�*��T����IٟT�b��i��D-�,�s7��/F^Q�ߵX]7��ŦaN<�N~re�R*�M��'�T��N�#x *P�D��lmC�k�=R7B�O��J>q/O����O�Eq�V�y���K/��j`��T�OR���O��D�<��i��\���'W��'�,���ȯI4���P�<�2��Tyr�'�&�#�ė+U�$�c,	=@@v 
�b˕oj剰$n ���T�-R>�$?�	��'W>�͓o��Az�lY 2ʂ�A��fl�	�`��ҟ���j�O�� 3l���W'b���)��ns�&p��A���O4�D�ئ��?��'2�xaA�d�r��� .��*�I�DH�F`p���o�$kXF�of~B&\1V��K6H
�j�J�m߿HKvt(�[W�	y��'�B�'���'n� F.�R&e��h��er�aλ(A�I�M�t�;�?���?�*��d�OvQf�ߢvy�dB�q�0Yx�Xdy��'r�|�����'$��(�j�*&��� $��0�e.�5W�"�c+O\�2��V��?�$�$���<!�,ҿu��L�JH��PqHi��?����?y��?Q������}�"G��FCE�0����	ʋ-�n`$�^�H"�4���?1V�<�ڴ�"�'�>dRg�99r��
��2Uzn��5�ɠ�M3�'�OO�9udU�S1s:�I�?�ͻ&]�Ų`�Q/B+�H�&�9O���	�<�IԟX�Iϟ���π X�W�Z:{�2���Gg�M���'B�'#*6��0�d�O=n�K̓2�Ax��+3f������5��'� ��ǟ��I�j|<l�|~Zw����
7nbhE"��J�g�:l0��H�n���v�	Cy��'��'Wb��qĴ��NS?	�>)`��,9���'��	?�M��ϸ�?Q���?y͟d����,'�n8��:$�H`a�_��
�O�l���M#U�xJ?��.7-��j����v�r5z�\�����l���?�3��'�4$���'i.P��xP��ɝA�����ҟD�	Ο���럴%?I�':�7�9�!��떬L�|{��S�f�җ��Ol��N��Q�?�q\�pܴ7D� ��]� �
�2`��E�i 6-�� �N7m!?� �	�
^����2�����k��i�4�^���"`�*U��Z�d��ʟ�������I쟔�O�t�+��٧X�L=IS��s��$ɤ�i����4[���Iq�ڟ���4�y�Q*'ì%S��{o1���_�"�i(�O�O: yAҵi��D�=5V�E�O:�&��F,+ "ޒ1����Ɂ��'����L��n�HA�H[�7�8�2b��=/��%�������ؖ'�6��C�h˓�?F`��nY�`��#�K ,�L��'���^[�6Kg�&i$�t����o��J�H�E�U�w-]y+� ��x��߰��4�Ek��k���ɟ	!�	S$��	u�ȆL�<'����O����O���/�'�yY�*ռXۥ�^�&���� %�?A �iǌ����'���j�⟬�� %�:�Z�F��� $�֯P��Q��1�M�1�'���"̠f+�֝��(��V-Q��$��#� P�#�]� ��E���h%��'[��'��'�r�'f��"i��-�8]�c�[�w�l)�fU��[�4@n�K,O<�$7���O���p�e�Asc�̫,r
��0.|}� z�ȹnڡ��Ş.:Z �0"��4tl�T�<+��1H�D�I#xi)O���`ړ�?ɥ-��<I�Ο6_0�x8GN�d<�,O�����X�	����ȟ��'�6-�,|�B�d*���@�B"|噵OU+I���R��M�?�v^�x��4e��f@�O��a�'HE��N|���#�
&�����1˃<9���	�W�����L�Φ�2$(U�lD����L�\�	�D�I�����ҟ`F�TꎣUu^؂����yag���?a��?�üi׬5���'�R�f��b��H �EϘT��)<LD<iq�a�I��M�i��� A%JΛ敟���8�Xa�K�}��3���V���!�L�
�?��(��<9��?i���?�S�B�o<Z��4�_�6i��G��?�����D�ߦ��7�����쟤��|b�׻{P�0Æ����U��xy�ȹ>���?iO>ͧ�?ieg�	�b��0�H��qЦO?WvR�قJ�K.��.OX�����?�/2��	i�y��A���{2�
�D�ON���O��4���<�w�ig�A�N��Z��<p�`�.f�ܙ�V�@�l�r�'G�6-5�����������b��*-���c'dֶ4��� ��?��4J����4��$�S|��C��kt��'*^���� �\��J'6f��|y��'���'���'��?5�qhP-�)(wi/�}������w������L'?��	��M��'@�A0j�?w@�qa2�kb@���ihD�$(�6���X=�6�����v<��h!51V@s���O�@�k#�?C,�$�<���?!R�T�M�f�3fb 	��R����?Q���?������E�E$PƟ,�	ɟ�*q腕/|��y�G�*$ך<�d�n�%�����T�	j�o���
`%�@�j�J􈝯�|D�'\ ���M8���d��ޟ��1O��#ȁ)^@s/NB�{C�'���'���'a�>��-W$D�)�Em�B'�U:B��I��M#AG��?��1L�f����сH\5e �����\@	���O���O���.5�T7)?��q@01�'��C������o����(!�ĩ<A���?����?����?�bB�Oq��*.���R�"����D���a�Ȕ��d���%?a���'�ބ���&�0t�� 4���ʪO����O��O1�B�!F��M�paw�Ѧ=��+5f�+B��jЈ�<@��V���@������#���`�7��ɸ�ՄL�d���O(�D�O(�$�O�˓^�F��R��G �%"�
�47���3���j]��y�L㟬�.O����Ol�d6����m�<�d��'�V�<��@�ix�I�8&Z	���OupQ&?-�;-�$X{� G�f�Ě�`�Jh=������� �	����V�O�L|�R��F�|I�p��52�#���?1��$��g�` ��'�n7(�ɶ�̄�sǠ=$92�PN�li'�<n�'�M��� �h�ݴ�y�'��E8��ϓb!^1���^Q�f(���>�����,��'���ퟄ��ߟ���!�H���L�
P����B�^ ��O:�d�<qr�i��+��'��'�S�'�Ě�̜�C°�#�A|�@ʓQ��	�M��'����S��jff�/#��7M�Z�v� {��8Tƍ�'��d��x��|B��8?��qN�MV��M��{���'���'����dU���4��UB��/�Ly���#Dml$ȅ'���?���?����D�{}��'s
���m,�����.D�5���'9B��&ě���֝�m8����,DV�S2r�^��'��!hP d'M�p@B�)� 2ydkG`]}�D����ĉ��"O��bZ"��GL�+��Q�#dJ+R�U"i��cn�$��	�"v�TQ�_(��XY'DK�7���ˢfO?z0����:9�I���F�*�J��a�QcX��s� ��i4��c,�� R`5�G�0-?�*P�A�6�(���wr�\����
3V��A&Tc�F�0�&ɒ ������0He�'�R���s��/3&QC�%Sw�ppa$̄۠� P��X>�0zqC�a��hbT��lX1� ȯ�p=��J<J�ۦ�bn���.����e���\��y:l��xú�+`�\�w�xQh$l����@H�k��eP%/־j���s��0g@� ��­9�b|�6JMF�X��3��
hFpl�2���w����u�$_0�'�ţ%�2ܛ�HH����@C�2W
�`*�
	�6�c�ŗ�����'�2�'���q�4�	ٟ�"�Z�ҧN#B�bp�bՃ���?9�F
y��?���?�5��6/� 䢵��8gV��	��?��^GF��E�x��'<��|�� B�ԥ�q���r��8�ge�#��I�3VJc�H��՟���Uy��Z0�٦6��y�"dF3���!i#�$�O �D6��<�4c�-���猫r>
-sh�%M��8�<I���?�����T�O��p�S�DC��1�Ʌ-ڮ�ʣ$By/˓�?��������F�D����ޒ� �*w�@��� �Y�������ğt�'��{�!�i[m�������4�\)���E&DZ����O�O��a����=�g�K/�Z�ht'A�:'��Pu�Hߟ���ş@�'�P��R� �	�O����/:]�	�E��5]�Ԩk��A0w�ΒO�ʓ[ p�Ex�O2a�Ԋ�w�|��#�	^k�4(����Dދ5%�mZW���'���l�<q�Ĝ"�\XԊЙO��(��&�Пȕ'�Δ۰�4��|a<I觇��Y�pPQ�a�;
�V��I%6Zl�ݴ�?q���?i��i��'9� E���q�GB�7j��J�y�J��O>��	�L6�YCM �*�ؘ��{��m�4�?���?��bZ�i!�'7�'��$��w�*���A�w�(�A�4��OuH ��O����O��rEDQ:Ѯ�hd��D��HqR��O��mGj��>�����EJ�� LN�bi�$�d�@.&o�`B)O�����O<�d�O��i��` d�q��A�΁�1���O�. �x��'B�|�S� Ф��Q�����,k���F�OI*b����П��IKy���Y�8�)}&vܚ �P�)��[�o��	쟄��o�Ily�^�~�F_67�b]�cǕ�X_�	������$�OP�d�O˓/ֽ��U?��;���ڇ�@s.xL�w���x��	̟h%���I̟L�$&�e�3B�c���5HS�G�̅pԨ\������I]yr��P^맸?����� �':�����K�2��1�@���?����T��r<�� {. {�,�Ic�'E��@�0�'�剩�X۴�?)���?��'dh�	�N�z�k&"M�xÃ���70x�	����IG <��{�Iw�'|'�tz��X�}^DR�̔�?�e�I?+��q��4�?��?i�'J���Iy�jV�~�"��ƃ$|��@pcW�p�������5��4� h�;o8�qQN�d�Ni��H�M{���?��KT�)VQ���'b>O&-	�v����Aܱ�м ��D]�h0��OR�$�O:�$�$ �������!!�d�*l���O*,xb��R}2[�P��A�ɿk���	��$��1�S/s�[�'d���|R�'(R�'��I�qM��P��<�H�p�,aW4�Ѕ������<)�����?!�Q�!��Z33�����D?J���H^����?��?9+O�E�N��?��W%ʚ�Ԥ��,@�GL�3���O���?)L>Y���?eFC��y�@�@�̍���Ӑ$�xp��`���$�O��d�Oh˓ �		^?��	 2X\)Z���������O����4%���(��Oi̓p�8E���������ìE�x�I����IOyb�N9�맜?����g�6o&�0�
���Y��$�䓑?��U���(������$��t�����.��9��cޕ�?q)Oz���MϦ]��ʟL�I�?��O^�h�(���#Z�h�+^?J���	���)���?)�����[d�H��B4f�����̾�?����ii�&�'��'��A�>�+Oi��c�5n$eҤk�&5�y�6+�O\��2�	X�'�?�sNj�Ak]�`xF��ѥ4�&�'5�'����<�4�|�Dp�L�uHP�bjl�i Ȕ)H<}R�
�OR��6���|Γ�?����?4� ���WF3�y)�C��GCzL����?!��ٗv9���D�'��'���u��7O�n���Ӱ}08qe�|�'V�Iџd���\�'Ϯ�갍9@�yѢM>����&�I!3~OT�D�O`�OV˓3���gů
�pr&�ړM��Y{���?�)O4���O��$�<�P�۵0�$��$h�dy$�}A���V,�7����Ov��;��<�'�?�g
W 0�ZȢգ�+�p�!
H)�䓳?�(O���-y��'�?��J	RnaKg��#,H�@/ܽ�?)�"�'��	�i���'"��QA\�s���hQe���\��?I.O
�ܪBpVʧ�?��yg�S0�0�Bi�,PR�≾�䓇?Y*O�<�4�)kVh�(��	{l
�+�(֜x<Ė'&��1XF�'-b3O�tT��� ���ʸ��(cmW�y$*��'��]���gG7�S��#^�X��C��������Ҩ->��'��:O��[��'f�0����j&=�����w&.(�+O�Ub�)��ߟ$)��X'74�L�F՘}��С'![
�MS��?�^�j`V�x�O�2�'��P���y>mH�b��H�*�+2�'���'(�o�&��s�������I�@ִ��EJY5A�Ԥu��`Ў���˟t��iM���|����[ j�C5D4�p�(�x'(,O�iCu �O�˓�?���?�.OJ��M��x0���󆄲rG�`3��E�Ԥ$���I۟���Ty��'lb�H=w8�Q@p��.e9PqRfFF Ld�g�'Z��ٟH�	Ty��''�%i0�{�a���F�H1��9�B����'��'"�Or�d�O��" �������)t,Hi�ƕH��ۂ�<����?�����SE��Q%>�0'�~�4M��MB.;5|}[ Kܟ\�Iğ��'pb�'36�rS�'��Y�NuHPb�X4T���4�b�I˟��'�2hG6S�S��Ӽ��/I\0��ɱ�M(�B�3�R�	���	lH8:��$�?ժ��?J����$�\(��<�{�@����?a��y�'���^m���: �] 3��s�%	���O��D�+�j���i2n����Y�ʱWZ�O2KH!m>
7M�O����O��ɘa}RV�(��&�Td�<�N�g���Y˟�%I!?.O��?Q�	FG.�@��Ś=9O��{�4�?����?qq����	Ly��'�A+V���#����B�Q���'����&?���͟���
��tå���^*Jg�Ԝ@T�	��XC�������<����sޱ	$LS�S[����$M��,`eE�<a���<9���?���?a���D��x�p`�F&�I,,�A���c 6�7�V}�Y����ty��'���'�j����[(l/�|д�� lQnUQ�Z7�ybR��I˟(��Iy2H�E����DOlPՋb�V$"/�S�	Y�BV�8��IyR�'���'�9B�'m�y��D�,$�s���@{�� 4�'���'b��'��	�1H�<���D� ��-{@��}�F���iZ�S��d�Ox��?A��?�qaY�<���yR�O5#�����+B1&�ڧ�?��?�(O���C�s�t�'���OVLy@�Ä�]��;6!ʯjKx�a�T�h��ğ(���3�X��w��'N�+pV@��=P���`^trU���.W(�M;���?q���2Q�\!����J`�'a
4T0�а�K˟�IƟ�� �(?!(O�c>=����OS��"�$ B&����O���$�ѦU�������?�8�O&�s���ĭ��~9`L��BG�F��l��x��$��?a,O2�?�ɪV�fTI��Q�J�xv#�5S4�pݴ�?1���?!�Aʆj���SyR�'��$]#S�����^*!`2cQ�b�'9�ɜ8q�,$?��IПX�	5d������	�r�5Kʖ+�P�������t���$�<�����l�mX2*��y��4�jţn\�#e��<I����<I��?��?����$J5'2l�yV�5`9f	ҭ�	-_��X2��]}�[���Iwy��'�"�'��qeD�C"���C"B�6U)`'���y�'�2�'D��' � wTxR���\dri6S_���׫A(3O2u�Idy��'��	�d�I柰��#p�Pҳ��#�,�8U��7ct,�D�MSy��'��'L��#i4�ȩ������ef�iō��acN�����Ovʓ�?���?0g��<����?)�+�O�@!ec�W��������?!���?y-O�8C��S�t�'UB�O,�a �*
'|g~]�G)ǍT8D��\���I�T�I�$J��IY��|�TD�e����D��,X,!�c����'3��(t�o����OX�d��^��'��mA����Ok��@POW0��[���h�O�����B��$0��0擽f�r5JdaS3��LQ��#h���d�F��mZ۟��	ݟ��Ӭ����<͙%!�ְ��AS��f���N5�?Q���<!����$(��֟H	�)�01��\ ���Z�4A
tL� �M���?��li�M��$�O��	�Na���%�� ��Ek��������Z��)�N~����?�Oz����IA�o�Lp%S?�����?IsH��}T�'���'��'����A���НIg�K�S����Y���Ls��'r�'�rP�ܐV��8�0�;Ո#�� ���;��`��}��'I�'��'�p�� N)]\8m�����]�(���y�U��	�����Wy�.�BL�ܱqc�ґFa���I���rM�u�|��'��'`��'���e�'�>�y�-�z�Ԁ�D�>R��9��^�$�IԟL��zyB���x���yU��o]2l ��f :]��c�O��!�D�O���A�/����3?qf)0[Hѱ�mN�����N[ӟ���џ��'`LD�6�i�OP�	ڽj�t��A���: ��=��O8�$�O��7'�Oh�O���]<@)@���<l K��Y#w���$�<1�j����\>����?�k,O��:��!�ѡ�D�J��9�R�'q�'���"��'��'�1�V Q�dX="��E�
b�H��'�V}j��i���$�O<�D��8�>Yb�RD8Dđ�Gp�N y�솗�?� �F�<	O>I����'�,љ�FY��l���L�k0T!���rӶ�$�O���01w`Y&�8�I����S�? Xx����1�l���lM��� �'I1O������'�1�J��c��;&X�	�����*(�'�� �*p�b���IX�F��昌X��Ӷ�B dx6|�'b�I�'����������'~��FX�v�����޻`��4R���!�����$�O˓�?Q��?ц�Zb�h1��:l|@�@F�jl��̓�?���?����?�-O�h�����?Y+a�2NIp�8�A��4�C��O�˓�?�(O��$�OT��K��!s��Y&���?4h���p�d�Oj�d�ON�$�<���O9�S��(����
I�^��e'N�u����t��(�Iyy��'���'����'���&���X��I+R�d�+w�1di����ǟ��|y�#Ǻ<���?)���Z��)��8l��m����.������O����Of=@�4O���O��Dh>ٲ�L�(��a�f�VRj�3��O��9rZM���i��'s��O���3V�����rMF�R���
G�RP����?!��<�:\���ԘOў�I�@��������ր��$�����i��'��O-�듔�$^�gu ����
-�(�W�3��$^ zy��0�d2������\�8!
 ���v����C�"�M����?���i	vL��S� �'�6OpHU]���c�\�|=��J��'q�'��0�ו���'�B�'t���Z�l �qh#l27���["�'��MV6:����$�ORʓ�ywD�W|�� ���Ԭ��JJ���D�z���O����O8���OB�3����֭t�+�<Pԝ�fBJ�Tp�q'����̟��	zy��'2"o% H��b���d}��lLH$^��y��';P�4�I�(["��'@�Z��''�J �0h1��4N2@�Imy��'��'���'o�s��i��٩��Կ[��)�0�J?N��W_�l�	矔�	}yb��!k����$_	Jo~]���*X��uA���O2��5���O0�$�pqO�TY���$	��c�l� <��'�"�'7�IT �L|������� L
�p�2�&�es��Ê�䓏?y�tF!Fx�Oմ��@�<�^xEZ\��`��;K�=�3*Ԃ@��au��H̀�t����Ywod�Z�q�1Y�h�k�p� �L
4���i� 3���O���OP�O��d�O�Šg�A�3��	%�HC-�;@m��i�6m�㟌��ٟ���W�Sͼ�Ȁ (��u��/a�dQD�͙.���!��݄��k��	!��>i K> �K�CE5$��}�P��Q�<�c�9Dz���u�J�I2��3��}2��s�-Z\�����8ZބYqgb�?Ia؁���X�X�Οi�(��KM�{2��(A`L9���@H�<dd�,x.t0�/��7�l�q!L@�OZNi�fG�j���M	�l����L��:a��yv��pCѵ�:�QW�P6)�AI$C�73�bU`�o� u���'m��'�:�y@Ӑ	-�9F��8����̛Z����䌅c:R<!�I�(A�xP�Bs~�K5
:�ЋE����4���3�f̢q��&h���nZ���a�����m�ɱoy�)y�I�G�����>0�2k�����M�}G�OI��t��鞛�j���%
�I,D�t�4M;P�0x��ܺL�}���)}r�3�S��\��	�d$�KaY$���IuȜ:�J��Ҡ���?9��?)�%���O.��>�Ra��B�8�����"ap0��+=-eԤXgi�
�)	ۓ<�:d��g)iWb����A�p;��/,_F-�u�߲ia{�+�5K����G�>C��Y���	��]����?I���)�I}��T�������*�f�`��C�IF��5x6Gٖ<��x��1,����O*�ytD�7^�xoڏt��p9�G9���K�K}�����?q�̅��?9���c�C��8��M!q�X����,]��]qRg�# $��v�L�Tt���?|.���&+P�h�*��F��j,5�u ���������vȆ�ɑ@r�D�O
����+^�B�S�Ȗ9���=A�j�X��3�\/'D���#L�`�� ��D<�w�K�k����أTa$k���<�';$���̧>�����6O�7-ϯ|�����	>���(瀏	���I��`A�E`� �⊆�KɎ-��S�tR?��WÛ�V��a���V>�.�1�$�$E�Fq��q¤����r5�7�'X ��C���P�P�h�#�S�x$������O��D"�'�Mc�� J(d��S�}�R���XY�<)r�	!\py��P�[����!.	|8�����d�2k b4�A��p� �h��P�$%��4�?����?�3�ڮiѮ� ��?A��?�ݰ!�4D�2(5xƐ�Bj�A��kL��Z��5*՛�:�#7M�0��O���czz�HM"xS���q��~z@�3Va s�������.�N��ԡ�b�d����* ؕ�$�cMRj�n�`���H��?9��T�tI��S�gyµi�4���-':�%1@�'Q��% CH1$�H�dJd�T\��I� � |*B�>}2D,�S�DS����u�2%�W�F
�����/3��x��M��?��?��t����O�s>	Kn����@�A_m�A��ȑ-o��y��E�Ux�4�#m
sƒ���	�^x�A��U�l�Rq1F�Dwx�x9� 6 �ŬF�/@����:c�	�m�����Iҟ���qy��'W�O���3�כ+���B�I�.�<H[�"OJa�B���P�S�ƙ(���f��k}�\�T'���D#W�JT���Q������3!�d�xP�#��F0�թ'�z"��oz4��S �&�@��΃k�"��g�U<J���KK�<��ƅ>������@�Jݓq�GF�<!5ET�c2�3V��4)y�@SB��}�<�7�<I��z�� 0/��!Pg�S�<9�H����I�
]����XC�<aT��
�5�Q� +jR����d�<�d����|�d
R�8t�5��"�e�<��i�:��D2#G[�i���� �u�<��&~���	��[�7j���-�D�<ٲ�����$LӀHjl�G��]�<�Q��%x�D*#hT6v����AX�<��/ٔgﾜ�� �H��X!� �Y�<a�_8ߎ�0 �ԯ2�8�!�EW�<A�c��Ra&@�1Ϝ�Y����t�<�ϐ�q�	3���3�jB�v�<��U�H�L�P�\#RȬs!�l�<�	��y������܁B�
�X��i�<�$�#7B��1�D��w�5�7a�<15��aΡ�Aʞ48(X#��b�<1�(3
�̀�i�1%�����@u�<I�a�CE�HQ`k�
��#,q�<#��P�0����ќ h ���h�<��"I��>����j�0xUjk�<	�jR_��4��I�Bo��6ϐl�<ɷJ�WC<J ثW6�|`D�h�<v,�+-~P9�AMY�UD\Sd'�~�<!&FM,�щ�i]�&�:<[Q�f�<� 猙o�RT��凤.��]bv��E�<yFH�9[��HH �!V�p"a�^�<�;�L��s �XSZ�F*�V�<��C޸?9����ធu�j��f��U�<Q@�G�\���$�Dy�`FMGP�<�$̢rZhɰc!�C�t���P�<�5C��K4
i�׍�=a`�`&��O�<a���_��u	����7R��;e�FF�<�S�`5�=��΄[�C��IZ�<�P�A0Fx1gJ�m�d�"'N�\�<�� >R*�����:�XʦF
Y�<�Rl )D�HV�\�chfp�aņB�<��M�96(��n��G��4j �~�<����T`����*ߒ��tp0aG}�<)�_�|Q����a�2�#R�x�<�vչ���(J�S��	
���w�<��e�$E����qBN�1��p��q�<IDcY�,P2�br/�ve��u�<�D�!w8L�baءC,�0A!�T�<�锖O�*a�KՖ[q�s�B�]�<)��ƞS�X&��505�pS�	�U�<qeΝDF���\-�|�+��Qu�<CoH�D�h���$P+*����`
�u�<!��_l/"yѕ-�Q�*Y�7��Z�<���f|�dbѸ1(���G�T�<���+��9����u�zyr�CT�<I�,߄C^h�R$KL����)�b�V�<� ��G!iH���"��!���	S�<AҠɓ��� �g�<@�H�e�T�<A�-Ҭ��m��ɼ-8`�C� �M�<Ic(�[�$U)T�#O�|<�`PH�<) ^�a��� EfN���(F@�<� �a��d˞�L��F-2y%hf"O�`q�K��`��l~L��"O=�5N��n��(F��1E]0
�"O�=��e
L*��M�-@�峳"O�|I��"}�����̏�`oҍ#�"O��q�eB�Ȁ$a�M��%I���"O�3T(9o�:ԪC�Z-Ԙ��"O�IـƘdX�@'$8s�>�@"OH��@��z�!Q�G�����"O����N,@AX��8�H�:V"O�����X?j��m��5���g"O���k�=>ܮ�Rq��"��Щ�"O�M���܁YAf�����J�0U"O�����S�XQ"�+�H�:)<���%�I�x�:�-O���bGL�g�� P�΄�NHѦ��pfЊ-��C�I(zcl��D� 
���}�A d�N���"�@� Z�a|�Kʣ��ջ����*��B"��0<)�^;:M�0�ԓ*~�x���u�Rɰ�J©�jͰDgF��m��qA�18��ۧ%�ܨ�"��%�q�'�B�����M9��.�2%�>X�[q����#[����J5D������)b�U��jE��JL �) )�2I�R�������T�b>��ȅ�T���%{n�t
��! �!h׈�-OM�C�I�|ze�")�k&ny"H�s���2��J�,����&�lm�W$P���S7��S�����T[��N�<���tC��XAax�Jz½�񭄤@�"��'� �8���~� �h���$��쓄i�Q����J@�~Gd���$٘8[H�����a�,��1g_�<>�I�q�\qXg#�=uh[s�@�O	����AIW>�ɒD�$���� �j�PX�#ޭK�<�Q��'`m¡�I"|�D�ޅJ�j�4l]��,	#}��'��Pcȟ��$��:QH�N��2�>���/�^��h�A�W%��xC��^dJ0��O�
�@��T�K�A���f"�d�0I�HV�0*�O8XiV�q"���D��|��/ k�nl �"�dq�)�BX���`$;.�42� V?)�%��0l2� �3C/ ��T"M8qU�!YcF�0�)+�J!؜��O0ғ�B?_P�Q2霦E ��q��dS"TȬ��1�=+4�3.��Q
-X�g��e�^��,��2�r�I��pp2IkƎ��p<����v�6U�O����a�"O�8�i�{�g�~�dA�?2�@�KPX	:�>�d�{�F�1��05�0t���Rd���')t�t�J�<��%VX:v�V�J<A,F1w䰁@��ĭ�|�ÇT6�O�h���Ёk�JxHå�`�����'E�4��ƍ)S'�5���P&`����dJ�|f��R���"+_eF,����O��G�"��C��u!�
ɒQQ�`H<�d�]`��S0�F�y�FyY�,O���8�2t���/�F��y�,�v�2�L~z�s��
( � U��I����Xw�DVL�-��UZ�6X����:G!i��FG��1s�u(<a�C�:0^d�r2[���%�P�Ie���k��$�l`h��F
NR�e�}B��A�%�d��� fޢU��C�_O�3�h�'
J�{P�P�4,���e$K2v�=H� ��U�k��9�3}��4������B9A��MH�ă#��xrC��]��K�<���)�"(<�U��ᏸ����K��,��I:A��,3DKT �R<��IS-m����Ðl-����IV�IA�b���2��!�U�8x�gT".B��1^��G ŵ9�\i�K� oPb�Xy�+��jZ�8�E�1zTX�J��[��0��I$80Cj�K�<g���M�ڥ3�(��5J�;Q"�qu ���(��� ���̣|�'r��.�=Ad�q�گt���	�'V�I�Ѯ؅<��@��͉��ʠ[���QЃ�ˤܞ����5n���*7�T66�Ƽp �P�azBj�qaZ	0��(�yB��	1��D� ��(i��(Y��y2�V,"9���gC�bކ��q��+��b܎��!#J��p|�C$ʩt���c�<]N��DF5D�D�I�$�p�4�3<Z&��w���~��H�O�D���L�g�ɈTt���g�8F�qyg�Xn➸�-�,6����R�л�0=���нv�h��l[��+�R~
�{"�Q8���+_*�TL�b֯NJ����P��Q��z
�'g"r�T�0hs�.'7� )Y@M��A�2O��?��kI�+ODT��+�� ����W�qSI�	A�(i��K�x�Ӄ]�,Y�d�W�OΨ�O�/L��iJA�
f4��.O42'i��"�m�L��|�%
�'� R3�A�7s�%:Yh��I�0�CK=���ēQC2	�b�>��Z�H��3�>�B
*�	:O~&�l2��Ң�b�Qs,
�F���s�Lf�>�.�7�a{�L�E5�uX�������gO�Yj
䒡�]�@�@	E|�A��X���dAy��*���$�+\��9+qG����O��s����i�~��N|�4*��-/p�ɰ	�{����5L�]�I�z�ʥ�u�]>!sT�
�g�ပ �DF���,�<q��V�yB9�O4}���7O��jS@��4�ccNL�f��Sc-��'N�ٹ��Qt�#!�yK�\ M��̸!���ɹA�����K�3�ɢgn���E3V���$`ϸ_2"B���fj�rTm�!c����i�%5���J�!��E�b��O�ѵb���O�㊲C�ŉ6�ƫts��V�'��6g�X��ļ�$S�MǣW����˄%6]V�@� 3�v����d0��9D��Y�8��+�=t�ax2m� yz�ze�I/^�C��'�|�S`+4d���K���������Uc�Xyjm����)7f�'��̚"MR�Tf�P��3�h"}��N�-<���$�����3�}�<��m^)@��`�T�M��k'F3Z��:��7K�܄�q`��pn��|�<�R��*�`h��$AFЮ�#d�Y<�g	�K������1pGJ�N�����N8\��a�Jt����dΛ0tv`�&�I�"ؒ��L�U\ax�������d�¬z��D9e���1t@ ��^=Y��	w�Be?ɰ�"O��d�_������e�̨Bי���G"'��y���x̊����S&�<�C�I�W��4�@���:n�B�+L�čQ�v���B�!�h�⁕�G�y�aW�J,8]"�I&�3��?;�V-��ʭq���q�P��tB�ɝt�Bq�sĆ<d�����Aڄ��ӃT�<Ch�s���D���5\�C2o�5N��ЋU
�[	꽄�,j�t���JO��K��K�b�DlC�(Ű,}��*V�
�	B�	�'x��F�R��M�E��xJD;��Ĵ}��5f/�'��ܒ&��v��ɣ�NR�i=>��~��R�g��J����NH1W���o�X���a@��sӊ|)�N��v�3b]������"O���̭q�sA�ڨ=��Yp�"O��Z3�˂^+4����8N���6"O�e[��CK8y���m4�\!�"O<L��"I���i��āJZ#e"O��ٶ��?�,�-V����"O�X���5wJ�QV&D�W	�٠d"ON�0�%
�H�&U�F�	���	6"OPDx @��P�B���K�"O����@��I�,ٖdH�tzމ��"OR̛r���JAb`�� KW�T@�"O^�B��D-0 x��ק"D��Y�"O�� No�*��oS0�*��"O�Ah�&��0�Hm�p��#�D|z�"O��h�/K�e��a0�d%h��)c"Orl���
P��|#S�[>���S1"O� �W�&�ҝ�vBB���u��"O�)�gC׺��]����	FHd�D"Oh�R�$ЂB)r���'RJGz:"O�ç,R�A�2��DJ ���Q"O�AC��ߍc"L�sa�d���c4"O�Z����F��X�$\�|�14"OftY�DO�~Ǽ�Br�A�j����"O6�c'+�
LN ���A�)^Lp"OΤ���'|��EƧi�8�$"O����(`ܚ���;D	,���"Op<z�"0^��#�U2I��Ő2"O�i���A|��UQщY�7uf�i�"OL%��'J�w̘��'�5CP@!�"O�M!�BP�&϶��V,��B���"O� 0��7@T��&��`��'y^N��"O���莂��GIR�z.h��"O8����S0{��֨
�u���"O�mQ�i�a!��I�G��^bB��r"O0��D�Y�1��2%��@�����"OH���ˆ;:C��QEE�G�&1k�"O��T٧}+&��t務|nDdA�"OP�3��Ǟ\<p��"�3�,��b"O�q��U:r�"��N'�����'n�+�"�/L��#0'Ѕ=T���[-5F|����T�~цȓP�65Ce�Ο$���SW�ACP��ȓh��}h2"�5v�r�CZ|�y��r\�����#��V�� ̈́ȓ���ط����x����܈�ȓFYI��[}�Xx�	"^� $�ȓQ�h��/ɝ#7�����L�n�����l�4L�5k��h���ڳ� �X��ȓ��
E�[�B(��B���?Y0��ȓB'�܋�c��,�}��P�"聇ȓ3�>| Ӄ�$)p2��$RV~Q�ȓ6��`�m��yW��p)�
K>����+�",�  6V�%�4���*:H��ȓ�*Шc!÷m �E#���*Cs&��ȓt�*��Z�K@*�A�� ���Y(����./t�L�afۙ81�-�ȓ�~��oO"/�<Y�� �S7&���,�ě��ьJ�ࠢCn���p������a�#�jq�!���Ȇȓ~E�<x���8Wxi���
���ȓi����C���y����(?(Ȇȓ@XE�&_7Jl�)PN��=�Q�ȓ>��TUc���Y`aE����¢h��$�u��PP%E".��x�ȓ?�������$5 ��b⁆.K�U��d�BH��A��2k�����>+�j��ȓO@p`���ڧ>&�[R��[Wb��K�J8hCm���#r�H�����ȓc� I��kN.>@�ӕ�H�=@�ȓ�<5�1��U%�,�D��ii$�ȓQ6�U�'��{��B�n�=��X0�92K�ɠ�ju�J�RhRA��4b,�A��O�D�H�Q+�لȓh�d�82�Z<3Tq�W.!H��ȓ`�L�ajD�G�f�(�Bˢ{���ȓ$B��jb�L�F�h9�r�O3r�X��ȓ61�XB!M:=-J�'"Ue��͇�X� ��&a���N��PPS��y�<u/�>ᎀy����@�P�<	���j�`9I�f�	@~P���`�<	����	n�����I!Yܘ��Z�<�ʗ4j`�#�ł�I	���z�<D@_��>L� sF��>��p�ȓ\I�pqÍG�b�[�._�~�������59!�%e��Cg�F0%��H���D�� �l�<1rB+ڷB�K6D�Hku� 8V�e� .�hJD�J��/D�$� %�~=X�u��p�$ѫ�+;D�`�6��� �)c���`�8�g8D�ĒSnº5��@T���x�8��L*D��C�=1��d�b�z�@��;D���gٹ3�T��-*B pb�N4D�()*I�2��|��ӱb��E�p�0D��c5N��)E21�cW�4��)�׍(D�@�$-�9fp<��k�1쵸!�&D�� ��Ԋ��3�&M(�j��W�z�"O:!����_��|hsIG�'%�#@"O�E��n��J��P�aM�hI�P"O$M����-B�X�g/K�&cn\��"O�9��Y4���ATΟ�=W�(�"O��c��Q�1���r��qN!P&"O��K7FK�$sJ�4Q��u�G"O>�D,�>w�I��IĆ�r ��"O�dɒh=*t��y���8��m�e"O�8(n���,�)"q��Б�\45�!�$�3�<���O� SH���-��N�!��B4��2>;.lCqMZ9kv!�䋩$�,\��`SՎ���KʦXl!�����񪋞&Ӿ\÷��1\i���
s��Ո�����eH��jdJ�Mܸ�>4[�Z���#2�S�O[�l�1���aT�q��k>�ٴi6�tr��+�)�禝��F�l�  rBB�	|�14A?�䅆\ ��dLr�(��6�̈́, m�J8E��I�=e6DA��'�<���.9e�
4��Ps~���E@<
�����.|>�a�B�F<S`�X=km���ns�z��'��d�E�>YqL�/���u'�%�\@s2��X��a���	�hOĩ��@Hy�	<c/���;�D�4�S-!B�Y귈J,}py�'�z)Q����2�^-xI��@�8�f�G/p-l">���ک�h����'�C�2��Y�D��j;�	�%�x��Ͱ=���³�:�B��f�¬P�_�<)@�������u���(�'m��i &���z�C%~���'�8�"U�C7l�AH�1"�x�c�O���Ȯ��af��258c��'
�DpQ��$m�>`@Ŧ�o��y�ȓG�2�2�"�5g8���G؃҄<�I��\p���H�)�Tb��a�"�u����7-���X"�'�ސ��HC�Ĭ���0v���&D^�E���p$J���e�J��$xl��'�haU#5U��B�6O�,K �T�d�D���U0:�� �� -q����ČZ�\-��KR��y�HN�`h8�!n��X~�`r�������:��y�`��--��* �2'�>I��bM�E@Z(��nY�	C����1D��!P�߉*���&F�[gp��B:-l��T�T���H���/���>�O4�{��W�c��A�^+g	��Ym(<�wdXBԑ��3Hl��@�/L����H+jv���*�=$>B��Ě\ ��+Ѡ;Vuc�(�kO�x��E�$��S�P�D�,<� �5�1Ԅ�>,V���*B*j��фȓ#�F(W��J��9`NG�|'���O��S�̅�41�mP�(Ǹ`%* ��	Nlh��)˓X>��3�
)w!�G1,v�k��ƹk�",���=:��5��ЀV�"Ҁ����U��t�5�$Y%(��F�߆;^VQ2�!I�����$V>t��6B� (�ɂ���CeF����Q=�,��ͅ|p:Rj���0=a�D�_���a�d"+M�[!*�}�'�H���"�.b� �T$Q�qb2�`�\�Eu��k�%�"k3hP���K>:���}dJA�Bڸ/@��Kڶ7�v��$�������~u4L9�`��� B�N�H�O!l�P�ӠyȀ0��-3X�x��	�';�)�j@��6��f"���4K��dc�E+j��� @���=��)�c�1Of��+�]>H�SAM�������'���b1��&�`�ˋ�g�:�1pDJ<F
D�c*A-V9��{ ��(c�$���'��$ꒈ�p���W��9;�D|� ���YF��b��0aƳc���J��J�}FR�z�I��[�⼢6���y�(X�d�^�'O�:P2Ja�&j;�~�"9rԀ�UK{�XH�Ko��E�Z���$Ӡ��1����U ]��y�bN��-�p�B6A�����E��E����"jרdd��P�^Q&>Q�"�˙nP`�s6�ٿIO|�"��Y�uT�~c5n�@����98ء�É���)��e֏!��ǉ�-*�YxG�b���a��Z�U�h�:P�ߌ �<��)&�~��XQ��C5��
�/�XXb���h��m0�8PJ�E���W �rC��& eb�3�^�<���Tg�.���8u�壄�̅z+�q{�d�r�����IĔY�y들��%h���@��a{2D����A◊-�2�r���N�T��a�A�4T5����b��w(j����L�� ��hTITY<,P��ٻ&�.ѣ��ȺN��"�P'Ut9���T�V�N�E�(�*N������Ɛx}h4�FH�Ҩ���8�
�j��A�,¬��ā4)��3��"a����[b?�_>=j�M�� ;�9�"]��T���$���T-�[�}Æ�:,Om�áJP70�����j�y4!L�K��84�6����BM��C���QC�݃"�^26S�(��`R����(;I�M�;�5޴&���c0�I<7Q��z�i�,g8ĦO���q����q��, �0��1��'^�.m��E?"��0N�d��A��'����T��ܦyYB�����$ֆB���m%�HOFXaJ�luh6iY<����`ԡUf��r�F�&�E�7d�N���O6�Zw�q �OH��8ǅ<T���Ć��`����3���A�`�~؞���� &y^zd�vꆅb�L<a���5�A�c�W��$i�<���*�	m��S�az��ѐQB�1���7j��d. �V(�G� �]�e��GC.���-��YZ@��FҺy���쓝Y2ٛq�5}�g�%?5��9�$��S� �yǂ�V���6�QIB��8��I%2�,���1�Xq9ǂI#c��gyrŚ�SO���&q�h���`%��D�9b@�W��8
�Yqw��p|�0r������q5�I�p�zE	7��b�?����	V�S�����X�C�p�����e�����g3{��T9���<P[�'��[b%:sն)�E�%j�b�ˢ��!^B����0o!����b΁#�*�p���*"�h�j:O�=�@ʔ�k+���i��)������E	�.P����;���������'�,���X���Da�S���b뇒^ riq�L�=��=���%� �;� �4t�'�X h�P�Q�<���M�'׼�����2g�'ְ�H%�Il� ��B+�j�a�O�$"���M�� ��
6U)�9���Ʌ����1�Ҟ�.�!���T]Jd���]�,��d�Q�>�?�ax""�Mr�#�U���&B����� O�z��1rߓ	�L�Q�=#6|9���._�᳦�Ճ[-�Ѕ�>�nd)� ��bn|��O�4�Jx��(,O����M�<y薔���lEssG��9Q���0��}��A� �m�'�ECF/Ӑ/�����D6���e�.�u�֧yT�PJ��7�8y�O����49��p�����s�Cj��wG 1A&���@�vh�=WdpxsO�9%`�W`zqZp��9e_��3b�����{��E��"<�'3J���cot��aЭ�5f�4��6�A�J��U(+/�0���^�u�\�JJ�t�x��C��W��'��A�f��:g/��i�����AK�}��S>=��+���~��\᥎��p<9C���+H���w��n��$��G_1XR `��9�Q�`FW�dp��!q��8R�kE����DЂ"#RT`1���~�5[`�$}�j }� h��J)!~�	XTlTj�OΨ���ˋ��>x8w��4@�Ԑ��'�4��1�&4��e��q����G�9Y�Pm��I�/~Z���������a����=:�RTz�M��w% ���8Ol}��9x��E"�H�$�~�'�җ!���SL2$	C��'LOxi���Z95p��q莍KȮ$���'����Q�ׁ{�. ���^� (;ag�t$��3���X
�Y^�<i�KV�f���+��H�rZ��Y��q��۱re�E��W�#�v�(�䂶�����M?H��eڴ$P�� @"O^d�6/��~M^̓�i��>���u	�FR�f��H�I&0��A��L<0KH,nddX��T�h�(Q���C�<y`J�S�~�3��d����~�<E:�@�"�/~���U��{�<t�Ԓ͢�paj�J'zq��,q�<���ZG<(H�U�Бl�lLX�E�p�<����v�|�J�@V͚�p%m\i�<���T�9&e��H�gu����b�<viO2��裤b@�p�q�%h�<)��ȝ������I�c��+�aZg�<	P�ވ
�|}���J���fT`�<���U�Q5j�b�l��"%�����_�<�� 	�$���Qa>_�XIЁ�	]�<�����:�)��9	9ީ���[�<��չ) L%���T����O�<���J�V�^��ɞ*枘�f%DN�<�#�	�n�;�%��f��J��_�<����F,1F�q����
F]�<��^<]�@1'� fLD�!�a�<i��M�����a��-��r�t�<1�$�
 �а�Q)-&��5Ӗ!Gs�<�G,�5$����%�ӾN֙+��p�<� ��[���}"a��^�0�kW"O�D�%$ık��&�Ʀq2e�5"On�0�kD8x?��Q,�.en5��"O��5�L�`��DK���@]�բ�"O���H�:9�Ȉ�ʻ}X���Q"O|���De��l/A.����'J��y�#�N��T��ų1�p��#��yb�S;Zl.�@V-G��0ɚ��y"�x"�,б�I�*CZ��f&��y��Q;B��]���^�(�T��B��yRn5%,�:PE�(����̼�y�k�M}@ �應W[�ɏ��y�B�:Mj� &�Iް�(�c	��yR+Z��`�$�^�9q�YC��<�y2�-i��1c��zPx ��m�7�y��V�Sm����ѧ\5��kՆ� �yr%�! 1��ڦ*��Z��R�Bř�y@��v��Y�'%ǟgz` Y�mT
�y���5D��8�&D�1 �պ����y�J�e�"Lk!c�-��_�y�I��C��0ِ���"L�{�N���y+Q(oh�dd�ŏ,P��$�]��y�dэa�8�%ܒr�Xs��7�y�@z:��˃#]�	
قG%^�y�Í ���a�ßt�X�#G�y��N [iT�� �̕t�8ղ����y�iٗH�%���	t�4���2�y�,��e��IC��9��aE
���yއd���B%��>r���3$�*�y�l�A��*Ul��cb>�
&	�y�n_�pb ڢ�_�v`�o�3�y��- �4�õ%�St\u�a ���yB�Q�K�b"C��4M<����^��yRH��K7��ƥBL[�0(�1�y2j�u��ر��L"RI�ጅ�yBR2b�(3$��9v|���!��yb�׼\��q�+�@����1���yZ���/�[ǎY!��Z�|C�ɉT�$�c�M��`� 
����B�I/�H�8D
��7�����S�~�B�ɤ��� ݈M[\D*B&�LB�Iy�N�3�cE�0�tp����9'.B�	`l�	�J�_O�pqD�K�&2B��3�$@{B�-rLB�d��HC�I�-&�P�D��m&:���+�	�C�ɑ@�0S�B�eo �2p���C�I2C�� ԋe��r���%��B�ɥ,���Q�\�7��M�v I�B��-)�1���@��ّNC�4HB�	(Z?��G-H6x��#��p@B�ɀ(oX��� ۂ����y �B��6�~�j�U"mZE��j�4'��B�	$�r`�S��ߔE�j�3u��B�I�AERp���5JkD�p��SbtB��1n9�a�gL�-��'��]�FB�ɚ|m���*�)II���դ��{!zB�I1.~H��޴{5`�$B^pB��	oZD	���BJ� -r�
��2D�����@�}G*�BLƀT�~�p��.D��uB�#���P�E(�IJ�C D�$0C�ݘ0�
Q×îa)ެ`$!D���x���A��ò6K�9q*O:5i���M����B�a�-��"Oh�I���2��a�Z��$��G"O� ,�����e�Jۥc��m+�"O]ʇ<:����nW�w��"OX9I��^�S^�	j®K�?'� �"O4�:wܗd]�y8�d�%*���"O ����2�K���-��5�w"O��z"*�-1 ����1��a�p"O����`Y�V'L�+!G�k�걡"O qQ����9�6���1"O^��Ӥݑ.lJ��SE�n����"O4za&οgK�4��N�v��lR�"OB��g��4s���� K+O�ib"O���G3��lp�Ԥ5�L+�"Ott�r�A���� ��=����"O=����t"`�􌆋O�HQ�U"O�p��M�{��9��ġT����"O���25
��{��0>�}�"O��`!H<>�85"e���9(XP�c"O������f����g��lzT�Bw"O��Q��R�
���������r��"O�����̙�у� �"5�J�(�"O>}@w*m`J�`PM��\)�q"O <��ƌ"8�Ĉ+���d] �"Ov�C�޸}t�#��$����v"OT���*�(t#��׾"�HŊf"O�yi��^��������Պ�q�"OD[�Z�i0$��!�)�bqB"O�%	c��+n[�k�D�E�JD��"OB��1+��R�`A��NL�MָxS�"O��I&��i'8����*Y�)'"OЉ����db}�ՠ��Jx~���"Ob +5'E_�E*�-J�a�]�v"O��7#N�5 f����H�9H��c"O�Q�e`�
"�"c� q9�0P�"O�L�Å�h�jl���7k$�L�f"O��w�.~����6GΑ	1`�6"OR	���_>��$���E�j�Fi0�"O�сL�W��zQ$ɹu�\tA�"Or��î[
��d:e��5C���Z�"O&�s��P�$d�ua@�R!wʺt��"O�Lq1�	�NS��ЍR> �H���"OLqi�A�Q�%��L��$"O�]��,]8��:���o�J�6"OV�i$'ܛl|H��KI
{߲�˶"O�5�t�0$�WIzȢ�U"O((2�Q+U

�x3c��:�<|�1"O�Iw�����t�ʌ?��ԩG"O6C�(ܒ: �aq����GHt���1O��=E�TO^0 �Lj��}(L��G�y�@Ep��s�*�&���F��y2�</R�DQ��	L�
����Ε�y�B�LZ�E�¤Ī� �E,��y�iϠ3n��0㓽 ��B�@��y�Ƃ4�0h&�$�6		���y"d�>SM��)*��Y�"�	��y"�6#X�@J�ɞ)~�@9�y��K�V�[���t���p��y�f5e�6|�f�(���2�N���yҏ�{���'T�{�l�AMU��yR"W>>�D �0��3m��y�Q$V��yb�Y5>���E�<q��� �*�y��'o�<(�ҌJ#4t^�Hu$F+�yB�5�]�֏�-^"]k�/�1�yBh�?X�p2�*�$z�m�b�T��y�
n�u`�
�r'8�k�����y
� RК��7c��`k�훭rJ��s$"O����ט#\�{V��!3����"O���g�hc�@�򭊶�c&"OJ�Rt	 �NQ��
�&��U�""O^(Z�E�7hH�	*QaP"~:��S"O8�~��,;�	�*>a!X"O������a> 	�@��A"O"u��hF�T�Ĉ����[>�͋�"Ot��E��*�6x	FJ���H�"O�$k�e��N��WcWzb
$"O�Uj��
7&�X�@�ܦ3��Z�"O��ЂJ�\������MuLb�"OL��G X�T��z��]2y��Yc"Oh!�p�X'q����`(Gz��d�2"O41��A&�|�3Jݪ;F [�"O�� v�@�r#�99҃�����"O� Cwm։Ut�(�V㗚�Ң"O���ϑ^w�ؑ�Q����"O���$�l[xD�g� /���R�"ON%�P`�oj��Ć�<(њA�3"O����IS����Q��ߐa�N�"O&]��a-&������@�h�+"O&<HWo٘-C�9����1�����"O��k����"���p��X�H�"�"O]0��X�pd��Xã��B��tJ0"O��;��(3.��#D�E�i"q"O�9�t��S(U��K�m�PR�"O���CKC.+N�P�; �|�X�"O0<z�#���|l�n�E�"Oް��-��)UjO��5"c"OP��,
h�u-^�JPhf"O,D	C��Y�,�k_����"O�M3E�3-xT��INt8Pű�"OP����-�php]]�-@�"O�P�1��}�D���
�"OPa�3���s�p���U�D����"O���
�D��u��j*�n9�"O��"d
�R��=B���/%��X�f"O��� �I=+CQa�h �|<�R"O�ؑ��I�`��h�"���r��"O����ŶF�Pct�ٙd�~�6"O�	�av�("PgW�b�؉�7"O����틦���j1���q�"OJ=��������;��e�%"Oi��'΀<|�-��J3i�P�7"O��z��O�AѺ��ePt��p
�"OZ!��O eY~��wF�K�i��"O��D`Z�]�z��ƘvmHm�q"OԀ*��@g��CFM�CY��.�y�I�?��D{��A(R��\I�<�(ҝ$S��5���̐(
�NP�<10��]|85WD'gfd4J`�\a�<a�B��(���C�#Y�<d��-Y�<���T������3`T��xTdY�<qb���~\L4���ٺ
����f��N�<�T�O�9� ���jɫ"Th�i�J�<��3W����'N�6��EÁ�N�<鑬�e�����M��u�h�kL�G�<1 �.u�X�b���d�3v�^]�<��)��*A 颏�/P�j|�Э�[�<�+Z�6�$���DC* T&�<�s�ٴ]`H�'��Tȁf��A�<�T.��B�U4�@�P�Z8v� ��ȓ;��'�W�4ڐ�����yx L��S�? zp��k	-0 9sbFt��x�"O�jŏI���S�i�/{�Q��"O���d�e�`�1(�5ai�e	�"O"ݑw!��Tѹu��0u���C"O�9��Χ/ݠ,sw w���T"Or	�Q��(KrQ)�р�v0�"O
���D�K��q  Qܤ]��"O��H�}��� ��8�"O,L0�DJ.;��1�T̤�3�"O�����Y�.����3��y'�Y�"O��R�I�L�,q��C8&�Q��"O�iS��"e]�(���S7Xl�@"O���"#˒_q�R�R�@"R�c"O�I��(4	��X�7ZQ`"ON�9T(4-T�ݑ5��-`��ӧ"Ob4 w ���y��F $Az5Zb"OR��2��"X����	4����"O�!1ǂ͒,�t�V�=�E"O�PKSD�Z��Gk�7wx�ex�"O.���J(Y���dS�Q��0�"O� 
��� SR�3Ã�3X����"O��wC�<v$�v���j�"O�T��JY���)uHV�Ul)��"O��$k�Lt�<�p(�%E�֡��'�"T��A�ज*]�N�i�'% ����E��Ia�`�����@�'Zt=��\�|�H�q�ޔq�rq��'�(�褁V%kE"�3���f����'�����R`Bt8��X6|�C�'隉�c�K,L+�4�[q�,���9D�t:��A��ri�h�� >a*D��B�F�؈�����N��� �'D�䂥(M�� �ի��+[
�ȓ!%D�h�v�:^Z�H�qǐ�P����%b/D������[�6Pږ��(��	��@*D����!�	4����ꐺ.��#�5D���N�[/�	�V_+@���2D�P�Q���V�: ��<HP��Wm0D��86�U�ߠ=���,Jh�s�.D�L	�쀩4,�@cv��YN�S�+D�<�v�(O�*��W5���w&5D�xCv�}�4ARV�ժc��pk�2D�\K�N�jr�Y���_o�r����.D�p���T�VU��D���P�;ǆ+D��q�����9�,��{�|A��)D�l	mN!?=N�i�fĽM
lŪ��!D�\�p��6nf`B�F�1$ަ���!D��ӆ��� ���!v�L}>	8�?D���"E?B�,I�1B��~xk�#?D��p���j}��	�pr,���>D����Ta��I���}��B�?D�8�
��D*����R'Mʔ�W�1D���@攚���A�E�2@Ϭ$�T ;D�,c&�~�68��*�$t��Q���>D����
Q�M͠Ͳ��֡i�a�R'>D�h���A;1�!*�$�^��*R�:D�t� �]�7�B1�S�O�c�Δ�֌$D�D���h�9)F�
6J���B�(D�t��҃3�\���MǯB��3B1D�@����֌bdd��N��MIE�/D�H"��Χ��- �C�}��р�*,D��5��z�h��'h��=a����(D�,q�Etи�D�ǨA�PE�(D���t�A�p��Y��ɀ�2�B���!D�� �-ڦ+�͡�	F�m��s�"OV��������+c�+ﺀ��"O,D;w�N�u�2�+uFߺ�P�[0"O�|�`�F;2.��t��$0�v�{�"O���ȓ�kO��ib��=U��
�"O�|�!NU�~�ʴj��(.Q��"O�H�F����*�y_f�zņ���AS�V�)
m�u��.!�,����Aٱ�r�i�3au.Նȓ$
P��A#Ov.5��D�,�D���t��{v�=,��乂�� r8���V��a3��& �޼Ywe 9����@����%էXD}!`���c�Єȓ0юqk"��9�^]�WDU��V���JȠQ�l�7_�Qy�
E�r^�@�ȓZ���P��� @���~��5�ȓY�\�Q.Oy+�H7�ɾ&��ه�>����f�Q����$��6+R~��ȓXǘm�7�^%({�x ���1AK���P����2�ǆ } �i&f�*q`�p��F�	`�Oϛ��M)�Ծ_B-��
���x�`}����!b^�j�RI��p/�0q� d���IG-�|���w��I�"��7g�=j�'ZD>��ȓb^6bDNQ�J\�4b�¨=��ȓQ�t�9�S��X�ٲcԠ	�*d�ȓ@��Ч	�HA���c+�\�8=��):n��5���^�P��V��qrbp��\>�D�/	=A,] DC��<�ȓn��GH͙Z�v��R��i����M��ź�I���Y����3��9��:,ĩ(Ub�3$�`h��
��І�T���`�&F$�RA"�=�> ��S�����'v�@W�����i��w�	H�H� c)�hB��X∇�G�~�*%��7p��+A뉴O����r�lDhg*���IXsL:=M(����@��N�-Z x�ɕ70���H�<��5���=�x����4 ���ȓH��U(�o�95�d]s��G�~��ȓ*�$�5bЬ!�=ge��;O�ȓ{�\pJ\;#0Ƹ�vD�
|nI��+a���r&Ya}�s����ؔ�ȓ+5f�!��K;IޤH9�[.��I�b�R� �E��9Q���{����ȓ�d�X�&��&JP�[p�M<4�B	�ȓ0~Pc��7yZ�:�GO4W�p����ر0#-E�5ں�e���)�(i�ȓ����K�s|D���&)`i�ȓM�,�Hg%�<\��qt���e�� ��N0�����U'-P�p)L�( ��M6�J6F�='$�@�8��� Y9�V�1TbHˡg����ȓ[e�-R���b��b��Խv��؄�v��Eq&]�Qf\5Q4� 4�ȓvSr��s�F I�~}je��4~�ȓ��Vh��+/Vv� "O~ip�=�f�ehN8�Mhd"O}�3�ǹx �!tF�A�x��"O��q&�&~&��R��0�\a$"On�"w&��,� �+1�ۄ"OH�#��&�L�5�+l�"O.!���m0~�;$�I�(y�5"OXUQDH#�x0w���f^���"O� F�1�U<�ҁ��HZ�X�ܻ��x2�'I¤K��˾`!��S4������'"r�(tD�$`�j$(T�1�;�'�4P��dʄt�B�r��T�����'}�Z��Q5�(R󀃓Y�Zt��'�\h O��x�	�Rm�VQ��'Y�u�*�r������Q�zP;�'ܖmRaٰ:y��4&�P��(	�')�5h�F��h*Nų�M=M��%x�' ڠ�"�3{f���@'[c�T�
�'8z}���ϱF��� ��O�X޲�*	�'(Ш�L��sc
�X�c��?9��	�'�^(w�	1>�x��eI$5�q��'{ ����D(""�dbW�<�pЈ�/�S�$bG�b������cֲ��B�O��yG��s�8I��CVFx�����yrhJ�8"�TN��@Q`�q��D�y"��^�8H#h��?1�pp�'Ф�yb�F'��t� l�"gྀ�qm�;�ybO͠+J��փ�S(=��`�5�yr,]7��1��G�i	@��y���	�1k�!ˋs,��9�M���y�K�)T�`j$��r����Oχ�y�V1���q3�#Zڢ�#'��9�Py�Ҧ6�H1�3��n)2i2"�P8�hGz�,]f:���K�^q� �F_�yr�P�*�l��ҭȻ[hޅi7d"�y2(��lG^|34IE�U�b�a`�4�y���=�z<J��F� I�T�O��y2B�
x�ԘWj�*/���K�	.�y�*ԩ!���ۤ��*�U��J��yr-�*-M褫��o�U ���>��=�y2n��A������	gG��x钋�y"��	V
8H��隳X:Xɩ��	�yR/�*/��`�g(L���1b����y�̋&vrNH��D�4pb�L��yB�0*�VM���@�� �q,�y�	�s��Tq1+H'y�N����8�y�h��;��� ��F���
�a��y"��l;�M���8�~	۳�y��0I5$}�@�͕)��!P� �yB�[.:�"Q�@�$�0}	c�]��<ɍ��_z�� N�kf��3D䂾�!�DX��u�Ĕ�xZ�	e�K�5�!�$�$.�44� oG�rI���'FPG�!���^p�VR3z���d��*��q��ty6!�3|$H�VICƖ ��&D��zf
F�tT�w��4�*��E(D� ��爉e#���`�SA ��w�'D�$)1�V(6%��0L�e����n&D�cIG�l���� ��5)���7D�x9�"j�0�P��u��<�9D��j���"-�z�qq��)M�\m3&�;D�<JT��?U4��A��ՐSp���3�<D��b��FP;�a��k�6v* ��;D��87��K�@�
Ԫؓ^�^|���8D��fOղ8 (=�mz��H���#D�4�Q�'J��+�T-<��ը�,"D�� $mF=.�N�21j��#8&l���#T�`Xs��\<�@&#ǒL	����"O$TY��@�1"Z=1��=_�N�!"OV�!VhJ3��m�Bǖr�Ԡ"O<�)��	F�Q򒨂�t↭a!"O�������� W����$$�V"O� ��q�óV\����Uz�᪴"ODx��K�'��� �c�&ypm�"O��)F"QF�����9n< qq"O�Y�-�sV�聢�:6W.�9�"O�ڣ�a�r=�v�Ăgl�D��"O�Ham�)��Q�C�*x�"O��QnF�x��A:�E°N�4�D"O�$�=�������1?��"O�Y� �8���X�@J���Q�"O �J	��-� P��C7_�L��'"O�Pȕ)�KM�E���4p�p"O��͇  `θ��
�CH�K�"O�!�bj�61`9X�fȬ6�ŉ�"O^����/G��9EEݔ|H�AA�"O�1��i�0v�x�cʷ#7��C�"O�%x�%�NH^1 �#ߙp(�%�d"O�����B���0ƑN� 1�'"OVdx��@�#������p�R�6"On��*P
�ht��g�H�@�"Od �V�I/m�҅�v�� b���"O��gB?�r	4Gƞ��lIA"O$軗	�L��2@�8@]�A'"O
M�@#�_��<
`2WzI��"OriǮ�1ɢ@�L�nO�肠"O8ii4���|�4H�H �P=6���"O�cR-��g��j�G�LL6 ��"Om`���H�%���	�J,ݠQ"O�R��U�d̐J @ʍ`=6YX""O���E�g��"׶'nB�"O��SC��y�b�;�CRZ��pY"O�:v�ʒ{߰�/d�=6oþ8�!�d��\&1 @�Ǯ4�lu���L5�!�dI������7B�B`rӬӮ=�!�ė�X��A2`J�6ن�S�G�L�!�D��&�q��I_[�&�z`��!�!�ۅ:�5��M�'�:�2J:;�!��Y����b���:��JǁPO�!��[ߤ����չ_T4�C#�6�!��N�>�
�ۢjɁNʹ�!"��!���>Ą�M�O1\\i��αj�!�'6�p��E�-svi�@��C�!��5b� ��7�J�Ap<趈�	Y�!�$ˊ9l��M��@�����n�)!��N2f"q�F���	��g�"yc!�ě�e�����/<oǜ4h�ϝoa!򤛝%Z�<���y�б�U��#Z!�$�//�H+$G���6U�ׂD�U!�H�
5&-��tv*�+���5J!�D�t \jAm���E�7�!��ҥ+�x��32 �2G��.u�!�D� -�$��!�GV��C]
i�!�ЄԹ���h+JeC�AD�<�!�@>#�á�̛!�tr���>l�!�Y�>չa�İ#>0��&ͿF�!��7MNqI�e�� �Pț�e��'�!�DC5a]��9������J88�!��/\9����-�aR%j|!�d5�1-���TY��sl!�dO5"�ܠg�Վ;��!�l!qJ!���:�F�׶J)���F�^�Fj!�d����츤�B.���TJ�(e!�$	>Ta֤"$@��(�r`IsC��`,!�$�n�A��GA'Ky��+D"�!��/	t��ì��(��,ssʒ�h!�� & ��#q�ҭɲo�r`�"�"O8���N<kؠXy��@�#H�ܫc"Oе��Ł(.�4	��-zg���4"O�uA	-�-�CIR�8�V�{0"OP�Pr�å�2͈�'ӡg(�`5"O�����L2y[���d�4
���"O� bU��+Jݒ���*3����"Oʥj���8~H T��Lq�8H�'"O�`�2�O�qr�����C��n!��+��L�.��H��Ҫa1!�$��3��
���
���!Ȣk�!�$"Ր-��jO$mu8�[pA�@^!�d�6
�
tR�5u]�M�� �<-2!�D�HZY�V��!TA ��?/D!�dU�f�"��#��Ta�� �WX!�D��]b��PoއU4�eѱk��[�!�Z��ra�U].�<�gK8�!�d��Xɐ
I#b;~�ap
t�!�D^"��AkB̞M�h�$d� .�!�dP9�t�@Aڡ]�FԊ�"չ:�!�dH'Q\M����\Թ��Um!��r;�ˍ�J���Mկo�!�ĄL�E1�A�n(�J@�W�!�ۘ0 <(#��Znl���'H�!�$O \/H�����Q]��P�I�6�!��)BQ:�3D�R'ٙ�R�t�!�ޱ	���9�*�M*1�t���E�!�_^u�-�0H�3]�	!����!��&a	dd �hK<y5^��S��%�!���P����� ]f�  $]�eg!�H7�e*�$\�f'p��tL�=c!���2 �)Ħ�x���K	&?�!�	%ՠ����7uT�@��='!�\�5�8uH�������#�WU!���W�i#��G���tAX�u)!�$��:����ϟ�{�Ty����`y!�DH���Xh
��,���`�'y!���V�B������)`,%0��8�!�Dƭ���"A�A�.��:�(�!�䞭|ި�Qgݏv�~�Ӂ�l�!� S9��Ą�O��BG. !t!���8��d�2^�Li{F�V�"!�T�Bmx=��@�8$k�Axcnݴ5R!��ժl���0�
�!���0��+*�!��?
�����W���KՃZ�!��D�!�2d��i٠3
�$z��!O�!�d��=Fls�j���9�4�ʆ�!��V�S���Aǉńe�X=���Ü�!�$[�W��lR�I���
V�͗�!�$׏K�ztq$�ӆV�����^>n�!��[g��K�� ��!s�$�I�!��X0P>���00�@��D��O�!�Dȩh1``Aѯ����ە �n!�䒝z�P=q��T�MJ������w!��(A�::�j�M6��[��Hbt!�[<����.Qj���Nq""OL�딅Q!d����$^.ܶ|�"O�e�aǰ*�����!�2/��͸E"O��QT�K�hX�Ԡч�2��L��"OA��ԝ�"���=;����F"O�=hҫ��pO�����{�`T��"O�4�c)��S���I�J/�4"O�Q&L��ҌyN&�q�"O��� ��W�4pR����sA���2"O� pफ^4��՛�o�,4WB9Ӣ"O�艥MP�Vﲭ��MC`7F9��"O�|���
m�� eF[�hyF���"O�B�B��J�`���b��Q���"OD�+�O��Bm@X`�	m�P}T"O��:���F���f��Rx2A�!"O���3���TG�qbC�l���"O@�ra'O�vF����
�V�;4"O�铠#�<-/z��`$+�T�A%"OU(W9H��P�R�����1"O�d�Bu|mJB�Ɨ5x��p�"O p�οZj��(v��!(t�ِ"O��e�Ǉwc 0z���56�H!"O�0w��1�`h�d�&X.X�s"O�T�B�@��X@���D�VH
"O�4����Vi{aX�M� \�"O�H�gg��Ե�#\����"O�9�j@>	����Nc�C"O���ʦ!m���ɠME:��@"Ol��E����	3�iPn|�Q"O���dID<9��!��]�5	ZdJ3"O�y*�i، ���a��L4�)�"O�����6}��ǡ@ �9��"O��ا�Tte�	�� \���"O`�R��j�8`��?q~μj"OL������(��zt�[=<|����"Od<�Vm�9�ē`���~!�5[�`T#��"�DԀ�$Υ0^!���
_}Z�N��H��שE!�dJ�����&C��)�y����!�$uy����$��>�h�B��}!�D�r��1�'XF)80�-u!���PJ�{�%��V?�&�F�6y!�D��r)���'�ɢo��!�D:Wٸj�F��	�&�ٳ��,�!�$ӂ{V�u�a
O �rqBc�E8�!�ק�L�U(�=�$T9D�Ա�!��гYZlkgM�$�P��b-�P�!�$�-A'�E�p&�V���@&L�?z�!�dG��d)��Z����H�
��a]!�$D	���A�<-�,E�c�ϙ$%!��@@,9�G��*/降Y��Ɨ1O��=�|V�U2 KB5���Y�|I
@Y�<�����%�P|��&S��4ٓ��<���
���V�`dܥ�4F��wɜU�ȓ͞��2&ДU�B}hD&�9܇�k����,Q�jh�чW^��ȓX3zBF(˘ ^x�K ���湅�?;l|��B��2�j��W�<E@��'oR��S�5Bl	��N��ëۃ
�����<��@	 `4��i���cN�m��	[�<i��<
��������2�@�~�<Y�%^�G%�P;qa �]�����C�<	�Q#t�!��]51�e�B�<6l�g/Z�����~HL�2���X�<a���>�h�Bң�
$�\+B�]V�<��IS>Z^���qD�w����
�x��%�\p�K�s��W!fK��8S?D�X�nU�U�Ti���B<�ycE�;D�ԐgiO`�4�k"��=" b�M;D����U9tH|Ic�Y�,$�˷�&D�P����[r,��䋕�� �q :D��3�胸WdZФΝ+�( 3�"D�`������g�6p��	Q��%D�� �`���]����i��N1 yf"O"Y���Άa��9S�KМf��Y4"O&�zpd�~�`d�\(G�h<�f"O4ѻ!���>����-ߏ4��$K"O4�T�5��5�A��,{�I�"O��؇�9	��,��I�+Kk%"O~�Z��*;�d0t�	g�Ѩ�OB��ܿjg �QRO[%I5��#�N !�䇲8����D9s�9�!�䚫p�n�)��Of�$ä��&N�!�Ͻ�>�	&��O*�9��k�!�D�p�C��|4�FnŪ+�!�J�7�h 9��Z
1Ӓ�Ʀl�!�Cb4^��󅋛TT ő' �a~�[��K�a�g*0H�J
�D��@�h$D�� �h��a=��kƣG_y����b%D���%�<k��B�h�:h���K�n(D��a���<_K����!�!?+���%"D�x	TN��d0Ii�'Z3.�>���?D���dcK-i����Uw�!�1D��ȅ
��@N|!�M�}|���0D�d�7��:':��s��ܨ4!3k!D���$�æy{Px�4�I>_ȱ�f�:D���$X�_�Y��F�	<�qp��3D���k�iF��E�[�:��t/2D���Q���L�� H�CX�L�����H*D�p�W�ּd�dh �H)+���S
=D�H8s�[�d-���}>(��j:�OP�OԩP��ƅN*V�A����S"Ob��u��hk$(���/YW.P�q"O~��@�Y�`�(�+�.NBH;b"O���ǊpL�Z0��8E5�kD"O�bd!V��	W ^��"O��{fCZ�EN.���Y�V�
d*e"O>�P�5�"Ms�� ��Dؓ�54�@u@��G;�}��산J�lٷ�+D�Phek��N�(В$�}o��J4�)D�Lh�I���H�ȌBo���4D�  T�H'W��l��	JȀ{�"0D��E�T�g��l�Sċ�*�16D/D����n��@�FK|����č-D�,���^�� �/K
5ɲ4�l�\��Bx�P���L�H��B��f�ܴ�ԣ)D��������¦�I4lԢ4K�C(D���/�y6%jfK��15b��3�"D�X
�\� "���t��	nu^!��I<D��ړ�XBrj�iUeԠUFa#u�?D��p����(�hH:7�^|���Bc#D�@��Z�+��š�l�E�����K"D���q픉!���h@�-��H'"D����\͔�BUDު\��� !=D��[�)l�(!��i�$F`Y�B� D���Q]�`�nX�M�A�$0��O?D����d����u��7W>Xͺ,)D����ǁ�_�����Z�J�$�%�&D�Ԋ��� 4ٖ/4 @ �zb�&D�� `�It�u!�A��B��#D��ʗ�;|��\���E�"D�\�3ǆ�EThYB1J�%(��5�!򤗼q�$��패&��$ʃ#��,�!��I�"F$�����E����(E;B�!�$�K��p�s{����@�a~��'��b	!�I�R� �8����-6�yrEG4f�����
���4�eW���)�O� 6���	r��)���T[�n ٴ"O����G�27i�U	��W����c"O�Q	Q�
G�$�U��8^�L���"O\�"U �$B�l��'�{��勠"O(�+6-\ Dxvy���	:���:�"O�����{���$�3m~��ʽ<		�_��)Q5�ǐY!�X��uG����ڸ��Q���,�2HHMaL��kq���ek�06��=�lɐjD���s�(���o]�v���O5/��l��b2 �
!�YTR���m�-����ȓQ��-Y�c]9
�vXSkӪ)G�x���%�� lR��5�@K[j�t�:�O2�.U�)�ő�'�,�0Mͧ?@��J��L��,�&���_�@5Vl�ȓ�8�P��2K���C�K�q�&���If��7MH=Lh~D@�ޤ(*����o֪���\Qj}���f��ԅ�P��D0�ふ*�-X�`��3F��<,e!�.�#��+�I�.�Ԩ��p�ѶO��J�Ia�ݍc]`��Y"�2i�Ϯt��D��9�>��ȓZon1[�J��`��dy��[7��ȓxW��T&�v�̹�G wy�Մȓ^{"��$N��� Ӽ
k�фȓ~_~�@-�hp��O�܅ȓ%"	8ԅ����)b��FAK0�ȓc6|�C� �:}���f¾��i�ȓP��<��Aۇ�Qpt��;>"����_N����@��Z�C���.x��@�-�D�5�B���)�&{�ȓU�� �4�ߌLi.a�%�����ȓ �~��ɍ�l�e���׽ ���5D(�W��	�2��]I�A��'D�$;�K�1rz��;,�1"T�'D�����P�d�!�ު���#�f"D��G�׊A��DS@�]�A���>D���!k�xY�$�$k[�*$z����:D��ѐ��fA
w��5��<x�@<D���Q�P� �@q	�3�����/D�(J�֭>���	�:x�}�hCy�������27��+�B�3���U��g`!�Ĝ;o��,�C�:25x�AƋ
D!�@.֔�(� �1�~݈p���Q*!�DDvR
�ZV�-p�8�#�$K!���3Xd�aT��>��E��+�!�ԁ�|���ε{P���B!�!�2�Z�� C� [.�(���N�!�dP�)]z��t�ūoV�ʏ|�!�$�X���/ѣV���ޓC�!��P���fLFkgN<C@i�#��5�S�Or�+�5z�8�Kŏ��8qV�{�'6��asND+Y>
��@�B�	�'(��4Y꼚F �'5.8�#g=D�\)b
=u�(!kO6(�:I��>�Ij��0@�	N�aW��p!I��T���X�;D�$�(К�2=��̓{�j�b�H8D�����](G�T����`�	�q��Byr�'A�O>����=_X 0��ǵB�p{�1D�<鰈NnbB�KE��V�zM�2i<D�l�F�IBO���5�@(>r\9R�#&D�����d��!�A^�J�<����"D�ȀQ�� pV��P��3T��ĉ$�$D�hу�0hf)f�O.[V|�ǁ7D�� b���E�~�B�lى1\8�a)#��7�S�'q�P���iL;k<
��AKX�;ɜy�ȓ���+�++jH@��+�6'4U��2�m`��P
F#�`{iԼg:��ȓ,H��2��T�!>�6� �PҎ���|����\m6�����q�B���v"q���4� pG��n<>9��"\�E˓IS��>�+�$P)h��ͅ�1����b_,m������ч����lM4uXVI�T��:T��P�ȓS��s��4zPQ����*Ք؆�	T�D��I����G�P�P4�N�!�f��ȓ*)�-8�� erv0�G%�yk�9�ȓ7W�q�e�V�L���A߷E��ԅ���?9B�Y��-�e'\`"�DJ���xRA>Y�.4��fF6)���5�D.�y�+Џ-#�����T��\#����y���S�n�����>S���s��0=A����bf���R�_�0�� ��Eفv�\�̓�?�	�<�X���\�<�0�Q�M�R�Zq��Xΐ��*9p6p�9��GǢT̓�hO?��U@�<$�MY��@F��ٛ'C}�ԅ�ɋ"x�`�5M��Ԉ0!�C�	7J!R���XO>�YA2G�C�	�)#R��g�ӆX`�P˕ș KV���3�$Le�ddO)����0+�
B��$8�O�T� c�1$��E�#�h[�"O�\��H ����cAHJ�-�l�+c8OƢ=�|:,O6��@j�T�-���:M�jD��"O:	���־Z�:U��ƈ%�Z$�7"OL�(#ɇ����h�'�@�:�T"O�M�1�������/�0����'�O�,ꤪ_{7zydL;���2"O<��C&-�0��a�Wx��t*c"OL�SP�އ-"�Mx���!\$Ƀ4O,�=E�D�'`D,('�R�1V�h��>���	�'�"Q�P�Fn�t��EN�*�(���'�� 9���,���#��"��eq�'�^0���%�<�ァ�l�����?�S����d��ʷjY�9�^e��yr��J�H�m��F&�s��y��@IRȹ��VꔋUޥ�y�" ��Aj��N
z
u1�͂��y��K�=��<I+u	��X ����y�MȚ&"\(���H#C�xU8�x��'1քI��̳ G�J��ST�PЋ��4�S�T;#����&Z҉pg*���y�A0�.$���ܕ��Ȟ��yb�P��� :b�	y��ޅ���%�O��TD���z܋A���n�"O������h���C���)c&�1@7"O���b���Wbp foߏV~x�v�')�I?*I*�� ���yZ�Ğ �#<����?q���`�bg��=���bAn�, 0C�Ib�4"2AQ�u����b�J<�B�4� � n>Q��AaaE,"T�B�I���!�J�{9b�/R&SDrB䉙�.�aI�%4�����&I�DB�	:�B[BD��V�(8+�BНoI��D�<��.�n������L�E��9B�}�<�fZd�΍��oB-AJ���/Xd�<y7Ƒ�\-���,Dɴ-��
Y�<a�.���x����P�N����_O�<q����@q���N��W놭P4dJT�<� �Eh�]�P�V ��ۓW����"O\4��͉1\�Yj�H9б`R"OD5��� �,����qe�b��hc"O�Q̍,@4�B�!є<Ж"O�5��i��X{n����ټiQ����"Ole� �$a5F�qAه~#d3"O�\
p��rr��� z��8V"O����Aq�e���u��ȷ"OR4�4c�;DTP�l�W�y{w"O��a���~f@��^w��QR�"Ol ��znf���.Ќ< �"O�aB7��FDB���"��a�h9{�"O �#Lɗ0x�XWb����h��"O� ��ԗGb ���L��5`�"O����	��~:r�87�V�V8΍ *O<��(��A�f�(�!�"�',��;��� N�00�(��>(8�y�'�B�
%ǌQ�,5a$�@�z���'�C!�Ȣ'r0	I���+Vľ�;
�'N��5a�"h̚���T�$���'G�u�G���|;�@k6JV1��'�\��왛-j-Ih�>�v�'��8ԇ�5Τ���΋��s�'�0L�+ħ��,�cAEP��ЉyB��F��"x��0k[>����S)^#5�?�����|*H>Q��дD�Zy@p�ُ	�t�{gF�b�<A@F�(�\P�Ŭ�!y��PC B�]�<!�%F�CF���z�p�3r�s�<92��=�ܜ�v
cG��k##X�<i��M�x7R���#�
P�~}�TN�_�<��ƃ(}�"1�#gCBz�[�c_�'E�y�(w~T �B�|[�!�&�@���'ўb>}�w-Ĕ!:��G�7�����(D�P"7D�p�DY�!E4���Z�
"D��zP�ɭ"h�:����;$L�->D����G�3̈́�W(]�#�@3��?D�2�斧XIV\��[���{�>D��J�&�g���;���	P��<D���TT"  ���d�55K�{� =D������D���,\d@*��;D�ȩ3F�4Ƕ�бb�]ݢ
��.D�H�mS,w��@z�����cU�,D��Z"lA2X��q'&ʫ����#,D����$=�:ݻ2욐} �)Q�-D��H��ɾ@���`�@C����E0��hO��$R��岶�S,u���3��1o!�$@�X4dh����"�� ��]|b!���.�8��@�9���!˝]!�M��쁚sڗb���� �ӻL�!�(���K�B̵J�|y҂�Z�V�!��yU�ٷ늜y_�x���h־%�ȓh��	�s�/Z��g���V����ȓ�.�h`/�7g����`��	�ȓH8a��A%<(�!��
EXJX�ȓ]�F�q��'%�2@�C��7Cȅ�o�"��Ń<d���(ᮐ�%�ȓ_*LTJ��S.?0 �1'K�}�؆ȓ5[��
�/��tX��O5ґ�ȓx,j���\�!{ G�2h��=��p�V�Д�H�D\�E��0��X��u���E)N(!ڐ
L2+���ȓL֤1ËM�,L̕!��0(1���'1�}ҩ��ߠ0�c�+*�$HR앏�y�Hȫ:�@@B������H�KȜ�y
� ���@�ѓYgR�A��AX��"O�,�fmg�9�t�Q'	�<y�"OZ���(�q��Y�"ߎS�}�"O��Sϟk�4�@�bxDBH�"OH�7bռ��(RDր
Ns3�:|O�̢a�b��{�c�8*���"O�	YE��. J�Rf�0R'�U��"Ol�BQ*S�2�>x�UD��,(p�"ODa)��M.�l�փ��Y T��"O�|8�͎4����c�!�4�1"O0�ؗa۞+>B�����8��l�b"O�ɐ�+��[�C�`�)^I�"O>�#��,v�4�eoV)����"On��RhP'Mo��'�A�3���"O��yBFȿp�@�nKu�8M��"O&m��-�h����S�Ӡv-B9�"O&���)Bdq4+�
E&US�"O^��c��4A���ZBB��C
����/�S�OF !òn�o8�$R`�I pHA�'d�����k
<��ҧ��b���',t��J&�2���4/��:�'6�芅Mӄ!�,\+��I1]r�0�'�� :gK�8r�����>�VQ��'Jz�2���7�Ys�%��7�dY
��?�)O2i�V�ߚ0�P�٭?�ʼb���TF{�O��'��P�HǗP�Z��c�E {����'��&S�X��|��J��ot�@�'�81����P|*�8#���kJ���'1�I8��3xf8�HH�k�����䀡s�tP����5LhP���*}�B�	�=J��8�k��M
p@�Q�W=`�B��֟\P�m��#��X�i��E��l�F{���K�^n�!k��>Ѩ#���LW!�K�}S���B�8�U-��3�!�DG�4���۴��8���_�J�!�F?^��$cO�T�T���"͠>�!�D^�	�d��M,U�R��C̆>����I(��X�cP�DK�ED�c2�C䉑MB���;��ሄO@�$��C�ɢ~ H3J�.XL6<Y�͚�]��B�	�7B��O�/�0t��
l��C�	�
��0G/= �	w�òMq�C�I#(���!@�"S���4�C�I�,�Q+sǊ-"���{t�I/{Y�C䉢d�F K�E��l`�@0��ǡ.8�C�����q�)��n����Kڤ�p�y��&�0��I�cr���A�+�L�@k�]FC�I�8��}���߁:x�҄�,|&C�=,����+{qؔ	�DW�n�^B�	�=���r���*��1��4�@B�	�S"�pbX�TW:���bIWB䉟<��q!�� �L�aEj�����D�O���u66Q���D��E@q�^5��$<�S�Otܐ0Bj�1PO��c��	` ��'&���h�9uyS��1Z1~I�gOx�x$�VGqz��s�rX�d�����69v�Te̱6A���%R�ͅ�.e����� �1��5��!r����<)ߓm��u���?t�3��s*����N�6xh���ur�Y������<1���i�5S�P+6 ]��2�
��!a�!��\>�X��cA�!��(`F�21�XB��&m���X��]�4�9��J>-�C䉵a��� ��::
e��ɢQg��� ��#Ѯ��3gb-"C�"u4.@ڢ"OH�c�O�@� [.(,J��7"O�D�E��:��HTከ@J�i�"O�!�n?NU@d f\�F�2P�U"OD�D�<F�1Z6�[�IŪh�"O����Sd>xkr��7�^���"O���	�[�ڱa��J 8���"O��5攌O��"ӥ�=��"Oș�+M��mbG�4l����"O�"6L߁b�LMHҥ��hR��J�"O\�4ł*�d���c[�pւa��'c�ɲ#��=+���W�`��lW�<tC�	�\�|z�Oɰn�~� �*A,NC�	�\�Z���ʟ�+�6��e(��"MB�	$.�X��08��`�A�a �C�ɠSL��J	)�� ��:a%tC�({n�Ѱb�=G~T�dKG<>^C�*]�`�Ѣ�7�4�sP�"~lC�ɳc���C���>{���#ß�H��B�ɵniVE�=S��](\P�B�	N�����ɒ5�Jt����B��$I�ٵ��I� r0��u��B䉴���ƂZ�:�J��Î�[�tB�ɐSc�$�a N.:� u�U�51GJB�<T�t̉��/]p�XQ��,�fB�	#bf ��,L�H�ʘ8�j�'K-B�ɼ\�����R
�|�q�S�1�&C�I��FEK��ܳ@��������(z�C�GU��ۦDˬ#Ҙ��t�-O{�B�I�q.�Tk�_DZP@@ �(7,�B�I�\�h��S���)lV���I�A�B�	�c�$	��Ё Z]��c��6��B��u���ۅ��?O���Ԥ�3��B��2���6��5H�����:c��B�	�3���DąV䲹�Q-��6רB�	�p+|4{��>:Тear�� sotB��+U}t���ɒm���H�~�2C�	c
��������@�kE6A�0C�:Tm�'�dq����3|C��a�k�� �]A�V�Ow�B�ɾs0��$Y�S	T�`2�R�C�C�I-U�*A�Ď1	�reyHC�I#�x�bD�D�%�tf�IY��B�	�R��c7�x� ��\@�BB�	�g� �
"��#nĹ t��d��C�I���AÁ7��ѩ��P2; C�	�VU��9G��&֨�c퐮=��B�I&BDn�r��۸��԰����WŶB��$ ��U���m�n�9�%@5J��B�	\�&�����Q��)�Cݡw�nB䉾�R�rB=�^��g�^B�	�4�&�����k�&Q�'#�<"^�C�I�_��́��K>AO*�ϔ6;D|C�ɼY�|�W��9''�T���άf�C��g[�E�C�-FӸ�a�rR�B�	�+6!�Ǒ*���
WO�B䉥ZrXXB��o۠�8��Ƕ7�C�I<;���R��8�5Hq�ƻ�B��2$��њS�0%���ǡ�4 �B�	�t�
 �'j�|s��� �8=NB䉤*eK���G��3a�R�o�VB�	:���qØ.x��JK���C��(~yJ!$TcF���T,9�C�<v� XX�d�%u��V%��c��C�)� �x��P)yʹ��hG��<L��"O"���e�n�nA����>7�t�e"O���Κj1��KN�����"Or��-��b�-K%G &t�Q�"OT��2Ȋ�#�輈���:�6ͪ�'�nxEKP)l�����H�4�Y�'RD]�U/O���i؁�H�)9�'�
��E-X�%�1��"ԁ++,m0�'ۺ �4�G�;8��`��?e���
�'�H�c�I�?O��1ʴo�X�r
�'A$Щ%+� ���P�R"�Z	�'���V�b�Y`a��B�l}�g�yB�ؐF5n�*�.+k�lAp_=�y�I�2}hA�F��*i���m­�y��6^0@�2�MBO�&��b��yj�#d���Se�q�Ő�/��y2Ȋ�g�FpW�	:a��B  <�y����UV*���چ,1�-�gG!�y��Gy���6+�.:�d�[g��<�yr$���ٓe��(3�P���E���yd��n@��[:(�@�9Q�6�y�.��?��y���]�P��(S@&L���D6�Ş�?QR*��mb��b�"\��ݫ�Hz�<�`ɀ!`5�\�wgфla�<�d�y�<q���l�$-�Ӭ� .���B
�x�<���gKb�8��N�Z��	:�^�<�B�,��C7�12"�(0�_�<������ͩ5o�B?��+BnVa�<1�jS;wE:�K0B�#|6r9���[�<���~.Q�O?8DE�R�Fa�<�2ĝaߞ� 5�ՎN�>E�C	DE�<�bdŏGG6ds'N�"<Xˡ��<��E�l 4y��A �P]�{�<)�ڨl�!irň�����n5�ȓcDyA� �7Q(����0�@i��`?�BK�>{���'� }���ȓDt4Ac҉�4��b�d�H����ȓKW�:&bؚ*ڔY�_�a�X��>8l]�G��l$���O�����u�(�&K�#�>�� ��YpȆȓh#�����'0�E�4���8���7����Ň�3���U.̷|e�@�ȓj z�nB�y;��蛵���r��w�@��ۖ;�JE	�-<!�Ę�l;reh&�6L�byb�K"B!�^��ňv��*�`��!�y�!�H�5'd`�Y �ԙ� ��!�䀄<bmq����*��'֜x�!��L!)�n�V�J�~~�Ԓ�%P�I�!��C%*�A��8h�b��Kа	�!�dN�x�h𡓸\�RPr��,�!��5]�4e�F�9� y1�F�!�䊥\�&�0eoT}o��l.o�!��Ά?Ш�
��^�2�����D !�d��F50uRDQ�dX��@�!����.�2lX��g DIKq��8Q�!�P;3�h��Z�O����D�)!�$�e8[�hB�}<�xX`���g(!�d�?-�v��d���O<�u)@c�)~!�$�2jH4�&kDC�,�b���v-!��]�%����Бw�Nݲ�ˇ-w!�N?2�@���D�����KI;!�D�a��٫v�	����Yª*!�A�}U�T��+!�Ԕ #j)N�!�� z�@TG_�
���á�ѐ��Y۠"O�H G�6'��8�p�"N�mp"O�؄Eϛ(�����܌p{|���"O�E3�E�JAy !@����c"O^��&��6o:��!�
l�I�C"O��#a�F7k7beȂ��9q]#"O]q�\�j������kaN�R"OT�3�DZ�x-�`HH�MM$m�"O��G�P�;il�i�N7����"O@���B��P1iU*"4ҝ
a"OL@�E(Rcȼ��(Ѓ}NdTR�"O��
���fK� T��H0�\1$"O���E��N�|�(PD�O+���"O��2`[��N� p"��1��I�&"O8-q����L����L��M(�"O|�P��
%w��Y!�@�!�D-��"O������	E(F�,��4Y�"O�@E��4r�r��e8;�("O���"?�L%�_�Դ��"O�,)#�)D�}!�d�4�H�S"O�d��/�l��1�g΁�J���I�"O��H�>~:~):��ݩ⪄2�"O��I^$&NJ�B�R�0����"OA��"Dl����F m�J"O�@`r��hGHQ�6*�����"Oά{�9
U Q��'��@�L��s"O�����g�|*f7����"ON��(]p	��2�F�.|�tU!�"O��v靚HJ�0{Vl�J�Xh�#"Ov0��ؒS||��*^<dn���"O��# MS+-G���y�f�GE�<�bI
�&W�Ls'��!B��s���X�<)�*�PT 
��@�t}6ݑu��[�<Aa,�),+��@n��hx�@o�W�<9�o�2������)Hp IiMP�<����|��"Y�| �|۔�XH�<q�7��ջq,�#q��+!�_m�<�SĀ�2,� �����PSg�l�<��$�(��2�n	�6Y@�@�g�j�<����JS����#���b��GA�<9a)��|�&���_�${��Vy�<�s�T�B$���G	V0�%C��J�<�$R�&��Y��
�� �)�	_D�<!F�v�4������u��d�@�<�u��**ǎ�p��KB����e|�<�2���8@�vK�x��웠d
{�<����6���yVO_*ej�`��^�<���6غăGL1��%x�J]�<ᱩ���h e�)D���0�.!�$^#r��4:#��"i�XUy A�ee!� [��q�U��*|�u����>OY!�DL"{�v�9���bBL�	c �j�!��Ǥ:\Pԑ�CO+a.��P�h��R�!�dY2)W�ŋ�Β�]\�)�h�O�!���c{z0�%�ą#��2G��!�D]!�&�"�aR%'���O,+!�DȊD��ӢD&q~8xb�_!�$)p�Ьx6@��:%X�!/!�!��OFTl��A;i��8@ʕ�z!�dJ�$d��qi�>�zd9PCƪn!��%	�U-$XIأ*J'	MB�1�"O@�t��*�F�&�޲�q�c"O�Js�\�8*������	�~��"O�(��hB�

N5"��u��K!"O� *Z�f��B*d��A�˹5^����"O�d���ّJ���	�-K�Y8R"O��@��#\b�hjޘ,��Ex�"O�$��� �N�Xա�(�0\�m��"O^t����q����-^��1�"O�x���. ��PĭB�( �"O.T�C���he�#�O�AF���"OB�˃c("1�Ҡm�}��j�"O�q�"����Z0��*V"O~5RAM?#�`���a�P��"O`0��`.X��7�@�{��)u"O�8buc�i���.E"3�>h�q"O�SR��MiVQR��O�x�XA��"O4uv J%|jD%��?L����"O���`%׫�0)
��A+|��-��"O��ڕ�S�R#�"6��HK�(ܫ�y�5�.�Seb�DARh("���yrFE^"X�p��S�)��� �y�H'h�!&��I�z,Af���y2Eݪ{XU#�Ԗ��:'+[ �y�c�
(��z֪��Z �F�C�y"b��?�H��v@��U����y���1ƨP�����9��(�0�y��g�H
l�w�)��U
�y�iM�4�臋�g���17�K��y"� s�-�V�R�R������ ��yb�ۤ�<��1ٙ|�nq��y"��B��|�Ck�6pT��ƾ�y�"�	L���CQ�v p�����y�G[Ț��GT?g(��Hڱ�y�C�G�6h���L+X2T,��\��y�d�7Xn�Bg���!R�D9�
�y�O�:B�����X���UY�!�;�yb�.\����g9K;��2W�y�g4zx�c!nR�Inّ(���yb�B�?4J]��mN<}2�Z1�  �y��F�(�і�#Ie��0O�y"�
m���X �G#̽C%����y�璹J:�Ą�3-���D
���y"EZ{G��"�m
,lb�rN"�y�aW?8:�Y�KO;%k�!тdā�y"H(D(�3l��"��k����y�>6�h�䇄�eZ,Ө�y`�ߨ�jR2^v�$���y��A%N�"�Ү�. ֹX��S�y�
�%6yT@Ҷ�B}� ���]��y��"�
Mщ]/t�T��"̈́2�yD��i�tI��ۿr�d�����ybc_�d�� C�Ӂ7B�������y"cӞu�l}���$4����%���y���R���D%@!0�(�����yr���8g@E��+�*=;P�
	�'.r�e!�q���d�m��'������4/����'f1"�h�'kٸC�֐u=BP�#�I�O#ZI�'����VR+��*3K��Rք�+�'�����d��**rZ�ɐH��h�'��U��7/��Y �A֍o�@�H�' �b2 �A�F���	�h�����'n��3e�,.a���ַn.j=z�'�R,J����:�gI��l+̬��'�v���E�:��yS���]n�
�'����7�N�_ބx�"�.����'7Ihw�Om¨�p�I=wdF]
��� �U(*�6��!�KL���B�"O�c$��,iw@�x7.E�5f�T�c"O�[5�Q�����H�Q8���"O�4�#�$jx�:+�Ly�Hq"O��+�3y�Qؐ�2aaJ��a"O��dȼx��B2V�mW2�3"Ov��g9D�h�"�4]|!p�"O��O�fL��E�88$�ѵ"ORxi�o�'W�t�B���T��"O|Lsf�R� �P䄎:S*(�'"O* �2|�����	�:D�("O����
�;V�PbƜ�0�0���'>tl*��_)J@����Cޣ>J�M�'2��iԓN��0��B�Ik0p�	�'{�  ㈛�9��8�b�BX�vPi
�'�6=�Cȁ$EEm�$I��-[	�'�u+�� ��4�����:�"�'�N0��@��'�v�R�`�)
ll���'�H�A̄M��8�ʜ$9�q��'M
,��=�N�Pkʟ=��
�'z&�x5��I�6��CӘU>�z�'�R��e�
	�}�Q�	S�>T��'�6��rlX98:ԑ�g�G DMl,��'Q2�҂��W�p�	� C;����'�x9�S�+FԼj7χ���(�'�<���8Y=�!���\�"9�A�'�V��rm^- �-²2���	�'�
�X�왮2��TkRc�#d��'�B9�#���&0��!AA�/�@���'�]G�B�`�ɚh�%tԙR�'�u���O, �x���B "
�'ܞY{B�F�7�>l��"G`2�8�'�j�SD��Yh.���_#5$��'B�!���5��(�qX�?�a
�'�^Ta����DI�*�F�1����'� $f+P��2a�C<���'"4`̄:>p,2TzQ\1j�'X�4�"K�F�p�H0��q(ȼ	�']0lR��"{^��RƆ~G��	�'۴=
�j�dh�$hB%�$fi��'�F��BNK5x&��!�ܖ	oj؛�'��L�5�wx�	��Ջ	De��'���¢
U�Vw����(	-LUp�'6@ 9�D�0`4���Y<m((͋�'�Z4���� X����Gh�c��D��'764a'@�hD���筃�2���
�'�E1��%�6	 �f�*L��i
�'��:��Ͳ?�l��c숒0��	�'�`�V�_����b�*S JU2	�'�8x�
B(&މJs��
!����'�n0@�	_c�j�*�h�	p���'hJi3f�i�x�2���'|unI#�'=>+�I�4��2+C4\W��2	�'�jd���D]�P� -ޘR�9Y�'Rހ��G�W�l�XG*�R��X8�'LDE�p�I�J���]�����'�<PkQ'��Sr�5:G�#^� �'���"� �O�� dl��(�P�'�ê	IM��Z�0R ����''���N.Jۂj��|ϠX��'n�i�p戳\Q$-a�D��v/�UC�'-DHF)"��x��J�f��t��'Eb�2Kɐ�衇ܘes�}��'=|��Ԯ]� �6�I�I��,k���  ��ē�G,�P� �m�t��"O����#ˍCƪ� �O�?�F���"O��C��^v"�xY$�J��8�5"O�P��9q��"��q�P)B"OL���!=����D"G�u~H�"O����'�kTDSWA�1k�xI��"O�e��#@�H��O�2�r �0"OH8�J���cX�'�^pI�"O()#�L�Ja�2KL�7ن��F"O:�;��À{
��sX�]� I�e�<1��O�v�����;,	��r�d�<����"�8B���7���*�`|�<�f�EF�t5��풳k�X���lTv�<�'bD;*nT�!JL2&	�|�R��o�<q��.ӈ}����s�D d�D�<�Ģ�
��=���HR�sE�B�<�55R��2$] �6D��y��[<����
�:�(���ܲ�yR�D�k�:�	�B#�hb2�´�y^;�� U��B�DI�a$Q��y�&a��V���AK��XAbN��y��ޗ/׾��#�JD�������yҦ�� 4�T#�	X�p�]�y��<p�4s���%��O��y�'�=&`�f���\�3�)]$�yb��)�j��u�_��a��L�y�@ɫsE���Ɗ!>k�I����y��Ia�$��e�->,�5��7�yR��>r�ܱ�S+��8�԰����yR	T�^���-U
fi�lbSx)�ȓ]����V�:T}3E�	e���r�X�"��/"���V&?��ȓ�f�d����<�A��e�]��5�@�"	܎�`�q�G��Vh.��ȓ3UR�I2̾�q���(6�ȓvU�L��	Kx�X9i�)#���ȓK�T�*�s�@����t(�!!��t���:�΂�M���3NT:*r!��O�B(�2BO����г*Κ*g!�[��%�t��e�L4�����8F!���x�{U�94F(T"F(\uB!�$B�/�2�Y�s�
t�Bh�++!���d0�uH��Z�|U��G�1�!��5S�$�Jc΁�^n����Ɛ�@�!�Q���uT$Y⏜&7{!��ޯb "��4w�nؠ���Rh!���< ��)f�Y${�����ݗiO!�dL|��l�L�`����#ЊQ�!��;D�0�h��;?J����y�!��F/>ި��]?��Ї�@;!��~�����O&�ԹBԌm4!��V/6�\4bh�F�Bb_�&!�2G�f��ē�&��!�F�W!!�$L$V
V��s㔯0^�[A��%23!�dU��Դ��-�/P]ڴ`ſ6�!��;E8�5��[0d�^ qq��6u!����"O��j$ �9�0��gV"J!��I�1� �����84��0�E7�!�D�4{i�����^��S�΃W�!��'���p�)
Sl=��'V�!�dV�R��5�V�[5DfE�H�!�T!0�b�&�((0j�ʐ#Y
T!�N`���4�I��ލI�_��!�!-�����2�RCL�B�!�� 0M��(�l��؆Ɲ�/7pbc"O(Us�ML"s��e�3Ƃ $�x�+U"Oꑲ�%Ɓ,>4m
��Ƣ6ỉ�'"O6�#V('Q�Jd�`#�	F��E��"OH��6��3Ҫy�p(��҅
c"Oh��w�"��(U���i�`""O�@����-GpQ9����7W��r8OH�=E��FӎS��Y[�IH�zE҄"!D۸�y"�Pl��8 a :oƎh9���-�yb��;|��y�$���3�!��c��p?�O��� `�P.���-
��P��"O�y��^"!>R�a7�ΝTG -���ɞ�ȟ���@&��^�r<9��PAf�b�"O�0cu��](Q���� 2�K��O��=E�.F�3��p�At�MPd���y2�-g��Ġ��і^T��  �;�y�BF�z�G�T(Y���2ł��y���,�8AI�.E<N��u�����y"	�43u2�P�T�������yB��:pdp�t���i4�w��y�c'@�K��J(f�^,�T�Z��y�� �u�εZ5�A�[ܰ�Ā��y2dӤX��T3�(T���:����y"O^%k�F�I���7L�D�q�Ȕ�y��O4	��Y�4ț�.Ll�A IX�ybF9f(���d�\*$��t�O��y"C	,u�( W�]�%?p��"Y8�yb�	��2���<���!�y�i�Rbt-9f�˧
Y4��A��y��0]�,I �Յ|L$L�p�F
�ybÏ�= ��#S�S�=!�|����y�(*X9��;��٦2|B��Gi�:�y�.�)C>��!"�2����G�0�y��ڣE���%T
{4Ҥ�����(O
�=�O���$�������R%l�X=��'��Q��	�]��Ұia�Hv� �S��y�a�+e�6���Cٔ=t��C����y��\� b,X�@7�8�+�,���?�'T�P���j���jJxJv�	�'�ZX���%Va$�9���*&��	�'�TU�PI|m���ܵM����'���L�0oW����'M/�L+�'�F��q凒K��U���P5@9L�+�'E�쪢aؽ"���Q���3�d��1D��[bb�7D�l)k���37���dq�F�=���O� �3��.��EIJSQD͚�"O�J&�O�5|����@�0d�a �>O6�s�'ў�>�9e
�.I,���˞@+�p��')�O���'��]qR퓿"�z4R2��"��H��'hp���5\R���
�&մ��'��+g_�Nm3#T)�0k�' h��E���Q`��S4�*hP�'�2=jv��+���P�،�h4p�'͒�9!�كM~QwJɋg��q�'=X`%�8@�2���c��e
M
�'e�X�*eʸ�e*�`�,��'�P��2����D��b�X!�$��'�ة�	CZ=�Q � �J	�'D��2��a!H�������	�'�(��¥�T�vD�΀�6��T	�'�:%�����f�fd����\����'���22AE	8���"��EA6� D���VE�ew�X���-j�z��q?D�xj*R�m��9�"ު$�
���=D�� ��Q�* ?$ܝ�$-Y.n���"O���c\�*C�@I��
�U�*�F"O�T(+���Ȳ*�1i�����"O̹$R���jE�D4V�A�"Oe��FT�,� ��Ԓ} ��3�"O��a��ˣ[�*��R�]4IM� "O���Dß
WH�G��F�mc�"Od�1E�V���J��� RAduP"ORL���O�y:x�D�� ���"OV����	C�B�CE��L��"OR)
!��O��)�ED�عz�"OtT�A�Z�n9A��E% ^��P�"O�����L&ֈ�I�I4d�D��"O�d��m3�y�	�����7
Y}�<i'&Ƹ4��(�A�V�
�.�C���M�<!�L6	���)������I�F�<���	�S4 ����� ٠��XF�<�%��V%Z�ۥ��=ۖ-�F#B�<U�ֶU���@ቿ"N:�� J~�<w���7��[@���lQ�m��N`�<1�/s�܁aAH@ /��u��C\�<�Qa�/g��S���aW��;�Y�<����~*~d@�EQF
⼫&��U�<���$#*8����6@�4-��NAO�<�l��Rk:�d0Y��� ���G�<��C���ŉ��5*ܜ����n�<�2(�%s8xf��-vE(�5�On�<�"G��eE6�����k<��V�Pk�<y7AR�R��ظVK�M�0!j5n�<�Eŷ\�~� ����N*R��Ks�<��JJ;e���1$�-*����EMk�<��3�ޥy��+B��I�dO�f�<Y`S+6��M*���<=�89Y��h�<���$/�\�Ea�5kT�&�c�<�&�A��$ˇ7���p���v�<٤eH�>����FQDh�`�� ^v�<�^��`ar��:8�H=0�"Z{�<)U�"W��8����:T�ԓѮ�N�<	�ٻqI���W�ȴ*+:�S��G�<�Ӎ�+fu��k1,˭ZZU��b�F�<��"	a�� �`Q�l���FA�<��m�6<I��>m8<i��Cg�<�2�J�2������
�@��1j��i�<A�`��pdX'nܶ'�HR���O�<��ظE� ���J�7��y� (�u�<�g��RO�\���ڮ6o$��#|�<I�֑B��������'0r��A�<A��ъb�P��&%]'x�8)��z�<�#�r0t-U���qzv��6	�r�<Af�å{�%��i�7�Q{d��f�<q�@�%S��k͢5�8���`�<9��h�j�s�۟a ]3� �u�<a��3�����'hk�#PF�<�!L=4얔�cމ׮Ě���]�<�eǜ"��q��߅/��h�O�s�<�qNL \�Ty�� N&��y���D�<���=�^�C�$l֍c�-�X�<!ai� \{f�F7h�9��\U�<1���)�����$T�y�}	���W�<�BK^�b�0e�cJ�cE�5)f]P�<�P���iD\�K��8l�xB���I�<Q@�FS���*�[�p��h
C�{�<i��K�J��UxgC�-6L@
C�y�<�'H�BT���b&�3zc8Ab�)^s�<� x�ؑL�L��vk�Np`� "O6���úX(	��Ø�$YLY�G"O^8C&�29o� �F�M8Hт'"On���� .El���ʶW�͊r"OP=b�OQ��؆� �X0c%"O��z�a�v�b��'b�i��!�"O��T�жP����#�@ V�ԉ�"O��%�ӓC׎��e	� d<&p��"O�����ŉg�y��a�::`"r"O0@
�ɛ%d-�I8���M%�4��"O�y:��Km�b���f��}N�yA"Of͠��P��Ƙ�cŋ�f' ��"Or�SF?ż�J�Ğ�R�:"O����/�yި�Rb��(T�"�"OJx;��AOpp@AᘕLEF�+0"O�E;Y{����*�+Fl��-�u�<� �W28��� �ӗ'�`���t�<	�J*=������X��|���j�<Y��֢T��y��S�TIN]���_k�<ɂ/ēnt�R�K��W�5�E�N�<�lP
xX��Pǈ�R�z1���d�<9`�O-'+r���@�n�9"�Ka�<q�N&ł��#b!�QH�<�*� ��!�ThϊZg�$�r@�H�<�f� D�)�L��nn�3@�E�<1�`ȊI$@(�2Ȍ/"�%C�MRD�<@/Q�+�r	��Jۧ��5�I�,����.��Y�wB� ᴸp��
�!�$
C�('�ݎ0��p�a����A
�!.r<Q�&G�s��p��9@��p��:d����o�tO�P
�iݲ8L�ȓk�2�1��#��P�0v�J�%��G{��Ӑb;�	s�Ӑ=pP��
�Zo!�߬r�,�Y�&"0��j	�=[!��="���@��-<d^a��&K!�DQh��x{"(�/3Y��g��I:!�˞?���)#[ 4� �b&k��F!�D��� ��ʾU�<��RR�!�d�4�Љ�df�[�����
�;�џ�G��!�~rq)�i�P����M��yBK�rV l)uO��B�L��c��/�y�/˙WX���6>,�(4��yB��l���z�' 9a+ʔ�Saܡ�y��Z�p�x����[�^(��M'�0?�-O� �.�~Kz!�g�L�Q�,u	"O���cb��P�7L�b���SA�	��M����27c<]�5�1��i3u��a!��2K��8�&�s�b�qE.���ֺi��"~n>��kV厊06!YG�&b��C�I���A�SS�3��(+V,�����M�R�'�1s^i�̪3a��~���$?�S�FG�#H2�f�� (<J�#��y��ĳ~�X|�7i���h�S�6�y�R�`Ipp��2f~�"" Q!�~��)�'zDt��a܎1��	����]y�t���R��7l0WsJ�s�Q�fĶm�ȓjz�y eSv�Z�[����?�I��Y�֜�WO���a�ˮhT���ȓ0<\9C�Z]{���Ӓ$��)	��O���d[�$�:T�H��BRj��0��B��H���V`*5z)�1ꔳ�DŪ�"O�kA��g*V�q�n�q#�ؑ��x�U�P���]}���5�$XB�Aքn�*I ����y��h���*��gb�H�7I�*�y
� �sDĻ&��I f\s�`�R��E���iA>�d�˔�U�@A8	�E�]ױO�������<h�)��%�]*u����p?i�O��AA��*_=!�F@����eU��sK<qǓ��@"T!�����r�Q�c�L(��	v���n ����o9��У.�Q6�hQ�'�D\ D��-9o�X��_9"đэ�$&�	���'0�Q�@cơ���Ce[�1���Fx��)Җ�E�>��p7�D��B�Y�L�C̓#���Ӧʙ�M�����̦{C��R�'��	7|2�4�A/�xdj���L~�d=�I�H��		�kC�S�L��'�� ��#>1���ĲZF1��U�$&�a�n���$;�Ov��N�G{�Yqnƅ>1��Q�O�=E�4Ŕ![>�`3	P�g�z���mY��yR�	g��h���EH��$͞��XX�4YjS���q�ݲ�@9���<Y��哕2�C���7��1
��U�r\vB䉠'���
�o�^�ϕ/v�fʓ�0?��1����)e`��:UI�Ix�D�'��y�� R0�H jQL��z��y����'1���O:����6� X�t�4G�^��"O�$"Eh]?[|6533�K%s�����'����m榅�=�O�Ѝ�5K;lb�-�OYv3�s���)�TO�'3Dػ�F�|%B��M�5�y�aRu�8��K o��#����hO���d�;�z���jM�X ��!hN�(9!��3OǞE�m3[�3T�>=%!�d��vM�����P����B��?!�dK�W� �@�զ0�8Ĺ�׾4��+}��)�G< 4�B.��������G�!��T�n@A��Vt��iY��D�uD!�ď$H7^�(�+�	rPܻEb��BOў��'u��a&`֠_�x����f�tB�IG�()[U܁`�v��� �vl�C�	�1p�(@��I�'����, #*W�C�H�6�[��8_�����\"���F{J?��%�@At���a��t@9��1�	L�	B�O�0�ZFI�5�Ab��܍h��
�'~�����jV����X���xN��D{��4H��8�Đ%,�\Tr�m��ybS����O&n3�@� P�V�>��IP�1��dY�k�D��_�j�B)���?	�ւ~���6(�}`��a#�[�<�2��m۔k+�?JԲ-+���U̓�hO1��D�L� 
5l��E	��cL���eX���� �gM>}५��)i��p� $D�t�0�_�$��BL�-.t�;��\7��x�eJ�Dκ����N�)J��:Q1��=�y�m�遢� m��(z��M�yR#F�r�b�=o�B�(��P���'W�GyR��؁G��P���s���A�2ВeN&D��YwK�J]�"��q�m*�N$D�䱐�̭-9 ��D�1Z��E���!4�l���V�+Ray5Gӫ[����T�e�<�7f�R���J fS+]��a;3`�L�<�`�W1���q�e�Ab^���SL�<Y���<�U-P�/6 �����U�!��><x���s Ő[�.��q�ˠ	�!��RY�G�jP�Ia���!�J�9�leq�L,N���g��4o���f��i��"|j�O�rEs��ט�ȴ("��* >����'��[4,�om�į� r��ߴ���d����̙$ �����6	�T��5#D�� �U�'���B��M0�e�,J��&"O��Q%�
*_ڴڣd��*Xi�"Oڬ�C��N���@#K�"�T�!"OV��¨��}T����C�u��1�Y��E{��銽<��hq��k1�(iύ&�!�ވY��,�L�24@Ó�	#���'�|B�{�]ѧg[4~?�����0=���eW3v)Xt�$e�qj�yF���y��Z7�4��Ŏ��r.lRf���yB�(jE�(��&j�n���,[�y���j�|�`I%[/�H���Æ�y������AN����t����y�J�.%#Ì<M~1�#hK��yͧ^��i�p�Y�zZ$y�$M��y��	�`�X��l��|�ɉ��y�n�666h��� {�mI�5�!��$��S*7�B�X5m�-�!�D^�Y���+�*R5�� �jʴh�!�䏇Oqx��p��-��u��"�7�!�Ȭs[ �bDE�.I���q�!�(Y�!�d�$#� ��tg�x~\��a;yl!�D؇mc6�Aq%�pi�	�Rˆ	|c!�䞎o�I��G�r9 ��)��Py�H�X�h�׭��Dl^�*�'�:�y�+:7�z����76�����7�y"�� X�Uj�/�1yF�� �"���y��C1�Aq�H ?�Э���.�y��-'&$��Ci��qc$����yb��R�p�{A�Ww�X��y2m�MX1K��Y�-�g�^*�y�c�k��! �9C+�PR�T��y���,h�l�� �-	�A��e���yB��d)�U�<�I�b"�+�y���(l�\�"��EФ8��+�y�,�6ߘ�)�a��?��5�A&��<9�ՅXp��4JNzs�����M�<����A?�d�F/'-f���0�/T�@Y"����t�E�Om�K�#D�x;��%I�Hc�Nz��E�ud%D�T�(�$1!|m	R��/_���$D� r��'B�ܩ��Y&�Q�d�!D� ������0+t
D-D��DZv+"D�#ENR4:�&�Iu�΀��.%D�(���٪i����N�
��4yl!�D��ZC\°_�hXl�{��Q�0k�z"�ە\���	$��R�t1g��'���f4�d�� �T�<iRAA$hF���e��zd��u��R�<�AGY�jM���f��p ����jEQ�<!�a�7�x����T�Ƞ�$�IA�<i��Ji��R�$�S9�T�R�Nx�<9���R��4'�� yv̠�)t�<!ӌYP���![�����Gw�<!5�^5?���f���(��� d�j�<��`�W�T�8��'b�U�%�DY�<Yf�Y�dd#L�
Q�D���N�<�����T�"L���D2/�๢��I�<����D"�c�!(DZ@�NCK�<1T�&%�:�*t�(kь5:�\M�<Y$ϖ�XS��4&�1i�� і�BU�<)�jǮ,�U0��TwT4�"x�<���B�h�:�� %"� r�[a�<�����#���� 7�yP J]�<�4�X9��e�v���P���X�<١逢`��г��4�:}Cp�DB�<� ����V7J�T$�*�"��%�0"Ou)P�B�9@�(Pe�V'-U�P"�"O�p�V�Z0\J4DЇ(۴^Y����"Oj��6D� r�p	��">3X4�3"ON�{w�;yN� �HU/9��b�"O0ܺ1��1+��YX�%W�d'x���"O�\�s%'i����!C�(`B�"O�@I1-5fN)(�m�5$��}I"O@�2� ��E �cXe�Á"O����m�k2<!Àg3lD&�(�"Oֈ W%��;�<}�FS�CZI�3"O��s-Ǚ�:���	Y����"O�q��mT�qX���o
UF�� "O�AB��{�,�/�Z"i3F"OH�ҧ"��-���RR��D`8�"OlI�`��r�G�=( ����"O"���l\���vY2E���"O<R�Lݽg�@$�B��jR�@a"O����4��$5���&�K�"OZ����_�����V��0&�l+'"O�{���8i_<�˕�If�)v"O��#F-�+�Ba�eh��!B��"O�Lȁ'(�lV �2�F��"O\����B�(0���*L��� "O\��A�,��� ���0� "OT��gĄ,�>A� !�wHjqȧ"OP� ���=���!��#{N�8�"O�ܫ#Ԩ�>���N��+��ea�"O<��k�?$ƚ�#�L
N�� S�"O�8��� �\�Q�JBv��X�"O4���鑢l�����Cd��G"O�����*c(��q��'/]t��"Ov�j�CK�����G�Ȝ�s.åd^!�$&Z�аHÉw��JD�،H!��W��\�#���8ׂ\�+Ƽ2!�ݠK��!B�ړ�v8���X �!��
D���C#K���s��?�!�D�'S��ps� ��.�
)"!DZdv!�D&6YPwIK6\��YI�!T�<!���Y&R�8�MD�ryj!����'nV!�$܂�����;e��K�iM*UZ!�$ʉpf�1q�ƄDR�	R��-u!�$�mh8��`ۦ7Xm���ɾt�!򤎫va�ӠՋp��+�i�!���kɶ@JC�͘Bw�C��֤4k!�;/�"� �Ƀyҥ�\ %�ȓ ��+�tɲ,����33֚�ȓ_`&��F�hiɧ,J�x�l�ȓWPz�ڧg�5��������u�<�3 @3%�}��F�PS� ���Cr�<�&� BL��+��s$zi��Am�<Q�Lķ,��U���]� .2��2gW�<�P�\�S5�-�E���Z� ����M�<)#&+5\�p�׍X�`��HR(�2`�B��<�&`ɡ%���'G��Y�J�!�D��">mi�'E���`��9gzh��jΗ,�N(у)�;3��c�'�s��x��ɠ{R\�7c��6�0��dZ�Z������<Mr�Q�	H�$Ԥ�B�O�OB��� UU<�pa��>�R��"O�[�Ú�z�u���X�BHR������r�L�M���X�e؀u�vPG�Dfύ���%+�0DѱEā�y�HR�$:���LӒ 7�q���-O�0�+b��C�R��d좌�T#���f誜',�h�	 Ҙ�Q˖�ȉ��'&�8v'�e��uyq̞$����ۉA{i ��Z��Uhr�i�zy#O��4Y�O�:o���1�?(����E��$$��;��q%��-\#�88T��ݟ� ~���R�/���FaЦ9L���E��)-� E�"�[i�D�/�(��	���<X� 8(�{�n����q6\ hW�\
?!N11u#���h�|�����=�E�Yo,�����k�h�90N��[���b:<O@-��gFܺ��� �$#ޱ !��1Xuh,Y���OhcR݊��7z<	�DdݕpV�.>kT�#th��W�^$b�	���OV���=#Q�0Ț�n12�$�+
�c�"���a8���J�ؠ0�Q�/i�ph��O��y���R<�� 2o�~�"�i�&z:,�a�?$��M��'�*Q9�ƚ�m��2�
�*q��d�c�S�Fd����k(!���Mg����O:Ic�����Q���$(����`�D�[^DU��i:�&��r4�K_J�U`�녳��I���*D�`�$�#�J�1��p<!�H^�L(�K�fQ+	��ʐ�3���{,�~����F�6�R��B�f���F��%4 ��툞����F�͉�dR
�'f<iS���z�WIZb�m�H<�.�5-��1�&�$k�d5���O���O�^P)�J^ @\x�;6-R�J�x�'�k��޵p���u		�����q#�mk�h�R���)�쀚��Om�Z;-)��)��22EĆF�����AH R�ؘ#����*�,~��Td���6���Yb��3y�6��W*���p<9T$M0_���Q/����
LX�Tۧ�y
�h�����!VG�0�$əH�q�^]��Hv��&T�"��[&�)
V\���$��C$�9)UA��YNQj�S��}ܧX�T��́4������慐�<qf��4��5*��K��t���ίd�ea࣑�X�hh��	ɗ|�����O]��̄g���13�O�J�,�sOVْ$b�a��8��}��"3��H&��(��Q�W�0�Ð�	���<��H�w��q�v� <<�����V��@�2�C�Z�j�K�C4MR.AT���Qq���J�0�a	�dh<�U�:l.,����DV�
�#��OZ̓V���@�[����֢��OSR�e��LXx����.:#�	�'�+�LAv�l�"�(6
�a:7�p��y����~�/Sy���D�X|���Nџa^�e�fi��u1!��Y�d�"����ҬVC����L0%2�kB;L�*�r[^؞�0b�[�2�����`E>	W,a�l0LO�LI�b+	��C&8O�P��`O�\;��a�g�9DZ�"O&T�É CZ�;��-t5�i5�|���v0�y%�OB��lΝ$]�PH *�T��'������J���Da��gt|�@��J��y;�����x�J�b��B�F�Lk���jX"��'�X�ZlQO�'O�-�cW
C�z���d�2㚹�4E�H;b�p�*i��0���"?v��IC
�PJ#�P�W�T8�!G_�'���`d��1���'�X4�a�b�d"Ө�W[*�2��D)!��)�#�ħ4���ӣ�Bd����_[3��%��ڇ�<�r�������ШڜA��1(�C��Z;�ʓkw
g�Q6�nӧ(����G��d�q3�H6Vh|Ehs�{�$�'����f+�3�-T��So�<��D�en��w�pئO��� K�#;�ړ��'��=�&�E�mxBu�V�9S���3[�ihL̚��W؞hcBM��X����w��7���)��R�w
D��(X9��0��&��="@��^� 1�"@�kd$��J^�EZ��bK3��`��iP�J�z�N��MS�IВ}7� r���8u�
|���|�Ό�w� l���O͔�f�F��<3Q-K�T{6I+O�Rs�ŷ)�^��H�b>��)_��[s'V����(��
d(VȂ��+�I2)`#|�'�
�b$;%u&�J�n�N�� }��*�@a���{RT^���Q&�ޤ< h8蠣ݍ�xBHT�\Q�5�#��.�)�5�ق~�P�3T�_�;#��"��G�*�P$Ԝ�.D�/L=%i:1�؅�I�KF� �>)�fD�v퐧A�gd�{u��GՆ�B��Q���?��M2C����A�ɪ[^Zh�2�QQ�"����KZ���K���l�I]	�� 5�&� ��w��4 �nB�I)lj�8��Ķ�D	���\��l#��r�HB�$���f>�b+�OC�� C*\�.��7D�*M�B����W�i�{l� p����Qd�

pz]��j�!�2c>c��򋉸si0`(�G�O��%PB$�耂�:��C���tDT�DM�(-��{aX�V����DľJ��z���a��S���L�aת��0<�,8ps�H�4J��PI��2��	��b����i��sf��7�ʁ��S�? pX�j�^��)s-A�R֭B嗟�3�ۀg'��s����Vq���ӛG������E��!�F��3��B�	�m�^�2$��"j�c��H�1�d�歔-E�M��;�� 3�*�3扼z1(gn�<U #4 �.!jB�	��(
G	K´X�OG�0t%�`#!�t��Ta͉ �x��	�t�D��.�w�V�@5�Њd�� ��	����*V�θ�q��֨0�b��NT�B*X����T�%��'��ɋ�JJK��Q��m��MW&,s��DB2��ݫ�j*ҧ�҆�7|�H�E�A[�Ψ�ȓU���;ʞ�j�vh°M�>��!oZr�DуE��s�^�)�n8G�]a��x6��j�"O����h�0�H�2��M�]��%��"Oz�i!�m�$�j���3W�Rb"O��ڱ�W�F�(H��&�m�����"O��J��]���"!$�P{�@"Ov��&8��ta��dt@��"OX�y�.��,��15�	�fi�""O�C�E��	g̡{�'��dƌ ��"O��t�ن+,ˑ��:~+�D� "O"����P��n�� ^�Z"�"Oj�J�#�$%[��@�` �3=���`"O�P�ǯ�)D����#�K���!"O��C�KJ�HI'�ɦP2�k�"OА��c�?Y;���E	�*؍i�"O�PH���&x*��*U���R"O��1	٧7�.���	D����3"O�� �g���R(�A�ÁԀ�k�"OY��]�`Ƶ0����>���˓"O�`�tm��\K\!��7�N��"O�)@o��@�|+�C-8��)�"O�qF�	\|�p �ՌR8��"O��0��V�}S� W�h�XY�"O<y��o�>+�J0ʴ�^� '�1��"O�� u*�]�Ľ[�OEu,"H�"O��R��-�ݙe#!1T-�"OzW�	j���Å�a��9s�@�m�<�d��9�!B�j.`�@ �
SL�<фCI\�Y��d��Oi�0�rI�<	 ͟����U�<Y��mpE�YK�<��F�4���7,F�N��`�&�D�<1���56	z���0	�$帄��m�<I�E�p��%��JC2}���(��k�<1�.��\4�UPB�*Eq�TPsG�k�<��������ݥk�̙��`�<1�A1%��iSXf�p�z�"S_�<�4����d	7��HW$D�p#YT�<)BE��[d���`NP�b5N�1%	[�<)� )����&J��v�93�C�<�姜�g'B���+]:e�<�	L}�<�f�3YA�8��1=���S`K@�<Q��"!6�JQI��Q�\y�IB�<�0�N�^5����5d���V�<Qԭe�hIpϐ5<ˈ�r&�Q�<16!�0���"�µ�X�d�<�֩\�-�����,��@� �b6�c�<)U���Re��X����}=&��v��X�<�sʔAT��r��*�!8G&�Y�<��^��]U-&�r	W��V�<�#�6S^=K�h�?A��\��XR�<a�Ç�).�ѪA�?:��r"KI�<a2FV��
8�󍊻y�0��FJ�<QCo-aVU��bm�{'�^zNB�	4%$P��SdϦ&Gp� ���;EvB�ɤA�P���F��t�Z`q·�U(B�)�  {��c�j��G� �s����"OB���B�l�����D`P�*A"O|x���e��{�+@�^�v�r�"OYH�X2g �	&/�)@��Xar"O��q0�{Y�E�nΌ@���E"On�"���}��}�� ��|<��"O-0���5ŒD��ç	eH�p�"O�5{��3;j�0w�ҜiB:d(�"O&d�jTD
�9���]N�5�"O��kP�Bs;�xRe�:ix��2"O`�r��߈g�!#d�D�Sx�x�"O�*T L�9��50P�z[��E"Oʽ��&��@x~a8E����,�7"Oθ��;B�D6������P"O�0�gdڱG��e�s$� �`2�"Ojh:#薫A�ň����F-k&"Oh$���0�Z���N�f�ԍZ&"O�q�ďT�cb�a"�k�"@0t"Od���-�00�skѽ1�~���"O,8*���]J��˷k�F��(�"O���!�zf�ceHR(_:% �"O�L�vL�j乣���2$O��sa"OX��G7l��I]5�s�"O�P 3��X�Rɓa��-!.�\9�"Oҥ3��N6e�e���K�'j�1�"Oڰb0Δ�Y�l �R�A�X0Q"O��+�����Ћ��F����"O܄�� P;6=Sb�P�v��b�"O�ͻ�JÁKF,�a�SB*����"O��C�(%_+X���ę*
�J�"O���"�ȍ6�hӇ�S�V� R�"O*��F'
������C���(f"Ofd�7c���z ���V�i{��*e"O�l�`���4ꌑ`A-Ϣ�(�b�"Ox�eKٰ�\���Ô=�p̳�"O6TJDi�2x���#1���]��"O:�c�ҖA`��d+Y�V� �[5"OZ�BbE�):�� Q�3L1)�"O�	���NG������ִ��"O"ȋ��7@�A���Y�0D:��E"O��0JǫP��٘oB�[Q�'D�`����	�F��Ō�"���#e�'D�h�SBF�R$�>K�����9F�!�$߬n|"��Աn�P�9t�ӜC�!��8���3k���W�I�]y!�d���>|G�Z�x,zR�F(�!�$ǩ_�,��5��z��]�ߨK�!�D͡P�2!J!BI�'=�����S�!�D�)z�P|a�˘?�\m�5o�6w�!�d�`y �G z�*�0N�,!��]x�
�m}�Ŏ��2�!�_�꡻��b<}��K�X�!�h2�7��uy�3��݀p�!�dŠ��$h a�nTt
'F�`�!�d�m�p���5?Dڼx��EX�!�䟙I{ܨ#�Aю.���AQ�[,E�!����2��`o�P�7��K�!�$���( 7�D�2d�� #gS,Gs���p*���$�L���~&� 2��׼uΠ��%�L[���� +�ɢ�ڬN;��F� �p9�$�?:Z���4�1!`0�'�Q����� ���$Ɖ� �)�
Ó%L��צ3H������?At�D����:o�8iM��h��_j�<-�Rě3f� *0b��b�э��@Pl� ��]�1:��U��h�*d8qfC
��r��WM`��hv"O� ���A��yE��y!��Poܐx� I�(¹�D�Oz$3UF�!1�1Oq��!��5�,�!�d��0k�{FOe�v�]�e�.�`�/�'J���Ĉ�SZ�y9V�	`��P��$/|O�����?t;�E�1�<(��B�'�����Ӎ��!��k�o��e�2q���n��a��D��y��;a��k��f	"+GBœ����:�lp�E�!AH�Kg1ڧTҌ�QTI�
c~�r����X���ȓJp(UJS�V���d.Ml��|���R�>�b��A������HE��<�֊ȅKr(B�ʑ2cw����(]��ف�Z~(<Y��ٌޠ9��!J�<?����M=
��Ѐ�M�l�ӣ�<G�C�n�>A�J>��##�%`oQ���#낌q�P�剢7��%���h�d	�0i㍐� P�*H�8�X�n�'h���@+[$�S��M����9w��iXw�ѳ0�(Tj�)AiܓR"��� T�ȟD̀r.(y2&��"l�#}pD[0X���Q�d���'��9�a��vnb)*�b�	;+�8�qO��~"1�ŵ)ȡKr#
S����/�4��쐯S�C�kRv��,�n�� v�]0`�>"=9��	7/���@F�.�8sne�$f]�f�*c�Y{X\C�	�,��+�L�
nr�����&�7m��r�y1a�N���)���xg!�,	$���F�?�14j;D� ����#T�)XEB�Ly-��ͥ>���(G�E�(!<OF���"�z���@�Z{<�1'�'�lb�)\��3ȕ˰!�!��x�4�]nh<�7�t�"�yRh��	!|�u��v�'������	a>���ɀ�k߰����P�Q4��#�9D�0����{�b͑&U��
v�<a�H�&.qO?	%,W^��E���U���tH#D���q��<m�
Yʣ��=��S£*D���Q�!�����|�T��2`+D�L��"��(�.Y1��Ns�pxb�,D����D�?��1gjK�D�Q%�6D���W�@>#̐h�#ɵP��i�!D�����)<~d�f�S0"���0�*D��	 	�"|���{\�Uõ�.D��Q�c�/6�ޕ��J��a��A�),D��;��)��0DJ�8$����,LO2�.���	����r���ԡIc � �B��4 ����ăT���z`˖�W�O��Z0kփU����͢C���%ͪ<�r�����#>�!�	�J��'cW�+��qP�o��ȖH��`>}��92�c?Oȁ�"��9)�\�"�݂/��|hE�DAax:����DZ�^���O����F
&g�j`E��{�HX�	�T�ݱcM.5��	�t$�@��*Ԟ9��Z����
�(�+��M5��Ē�iڞlib��*�ta{-�(�џlk�eI�M���Õ���LڻE���B�LU�Q�Uڅ�Ì�ē�E#_&Z�*����-Z�Ec�+�$\�A�S�˓pn�(���NhBҧ(�Xh%ÐwdT��&@ W�j��5�U7�'��0�=�3��-@����΄�k���çP>�tئO��#&N�
v����'�P�Ȃ��5}�d	�wi֗}��$34�ي(
q���P؞<saA"[dB@F�MG�@��Hޚ5��ȅfťb���ٲ�ۃK0�K�V�ĻtBS&d�\�V�AW��ya�#�L��A��ڣC����q�/��lE�!�֢��dA��@��|��,fD��P��O;2TXg�&�ք§�� 
/OhTj�J�^d8H��|bS"	R]�`JD9{�2���57'��x�s�:�g~"�T�/�4\y��'>�y�ѯ�)K�N�'7x<òC�P��ϸ'i^4cǧ�L���]��x	�'hZ$K�۹Q%F�S��z��%h��Ϻ�E�>A�W5
��?A2@C�z	QD;^<4XR�m�y8������x@�@@�#X�����V�S��q�]5	�4�����f�X44.I��e�R�����0B����ҷ.b:�uE�şprP�����}�G
ϐ4;��t�,D�$�R���	��(1���$��@� $?A"$�oC�	��A	&_ h�%�ӥTYʰ�,ǥm-xA����G��B�	j�LM��⁑Kv�
���%9�\�F�O)I�d)B��h�Q,�3�)� ̥�4�ڶ�ɘ"�76*�1@Oȱ/�57b�S&/G+]��%����h�z`#��;f�f��e�^��p=)`d�6b���#*J������Z��pe�W�4L┍��C۟{���C�50�eN@�]��B��5T#ؘ�@�E�iQ
@����J��/׮4Ѐ'�1�p�vꅙ�|Zq.�'�.���q���M�<y�f�4d�F�ccCՊ$" e
C�Un�a#���53P�@��'c6p�|�<	b�+`�+�D�7������~(<9��C(VK�}a�i!O�`!�q�^^��J��^$�f8����e�zr���8��t���_���B'ŕϰ<����0-�J�,�$P;B�R�����V�����ٷ<)!��7��Dc&�Q�'��aj�"NQ�(�U-5��@G���D-Y-�|�P���@l�<y/8�y�Hݎ&2��h���;X�p�b��M��F����"~nڵj��jB��'/���b�O�>�C�	=$�`h��S�X�����	ieXB�ɟa3ly��ter1@j�)n�"B�I�"���I5%��20��ɃPf�B�ɢ,��)���@,��� �\M�C�ɀ+Y��D��#B�@3��R6�C�?L��ZN��|�հ��C�"O$������z�!Լ[:ޡ���R�<!�k[�G�
�q��۸����oES�<��G�B�xE�-��8�.�a0�IL�<��.\�)����m����OP�<��@�F��X�̑��T(H��D�<yPe��;L�7��+��=x��G�<���Q(n��ȪgEx|�c���}�<��E��$Dn̛E��D1��m�<iRg�J慲����f8�6��<�w��- E�dC�]�QP����`�<ѳ�X��s�V�an|�v��U�<�Q�B�/.t���S�T�Lq�GED�<9f� 5��I��ޟeɔ����A�<�1�NPx� Ã_(
(�R��<��m:W<y�ĿY���!M�g�<ɢ K�S���l�"s�(qÃ�t�<��a�h8;p�5�Th�@�x�<�0+�O.�����N���Ԣ�u�<!4+�"`��S��s!H�Bg	M{�<QG��S�	��)	�H��[� Zw�<�$C�
qZ ����M��S�$�u�<�jI�9X�y�`�A&&�v�q�"�r�<�& ,B����e�;MY�8���h�<)d��>��̰�@�U` x�<A&P[��<`�L�-�JA2�MB�<��	�Co3�(ڂ�2�b�'��<ɳ�С��J��Q'`Y�awbBt�<�3&W����V��RA5.��<1�a��,%���G[�1;������z�<a�.�(  <�N��Z �����i�<�T��hR9���^PP�$���j�<1F�F� uBYx��-�f����Hf���B��2)� Kb)�>��}��A���b��U�z���K"O��+��>lZ��ԢH� t"O��W���F95ka$̵5�@`�"O�z���o��zEj��3}�MQ�"O>��bё=��X��ծoF��W"O\�h�!�-S�6i��գn�q�@"OP4B��Ɏ[!�՘��ÍYiޔB5"O�Q��/��:G�M P�P�d�K"O� dK15�,�4E*6�n�!V"Ov��&@�J����_.���j�?O6mɉ�d������E��
�n9ӳ�7���/��Y�e�����l�
�π �t�#�F:g;�݈�m�E��)p�&/�D��E��-x��OɈ��!��3hS2@C� 2�����'�A��!Z2Y�q�O�.:�'-m>i���;60x����o�%����&K"�k��/���OoE�!Ȇ"�<��b�J��z�
����h r\�T�a(���YUL����%hfً��32�D�cy�$��{P2<j�'<��} �CS*BBL���W:i����=6�nH}2^��}�
$?�*�J19GZA���mG�H��l�?��'�L��LO?�a��囿S%����	\�_ʠ�������^Ȥ��!�)�ӛX� ��g�(b@4���'QF�Y�n�	��:�)�'�v}�F䏎2�(u�T98LL���lE�� c���W��1�,�ڈY�d�Ĺ?��tqeh���0YH��ؕJwN��j+�T�H,�Wd9k�K:%H`��iȂA�r�ʬgzm�O�?�rb��2 X��Ï�!xx���ì'��)�U|���G>����@�J��)��PMh{�'D�PkgP~ Vظ� C<2�B@��0D�4��͇�,v1�2���i� .D��ǁ��<PB�A('a�ua��,D�d:a s-Jŋ�#�7��5i�+D�h`(L�=�Q��Ly� �3D��*�%�%�YSn�e�r�4D�h�G����!�dÓ'�b�Xt�0D������<��1��@9_H��A�1D��8��]�p� !��/Q��<D�ĳ�TMU85��f�4,�0!׮<D�������g�ޠh�W�U�Da�Wf9D�ѐ+�{|H�Ţ�=r�X��#�6D�0Z�hޖ[��A���Q>� �s5%1D��U$�D�`Yru�JOT	�P�0D��@����V�[�NÙ0\�:"�.D�P0�!�7|a�T�g�4���>D�0#T�2Z	���+C�7J��=D��K$��cb��1` <<$"3&=D�d��G��zq��%�Jm�p��>D��W+�<Q"UZ3H0&�����:D��+sT���h�)/6���N:D�����R)$��81D�Q><��,D�$�S��?@�Qkm2�L����(D�`	GȽ-�`�@���lr�	7n#D�LZ���9o$�Y��ޯ	f�§	.D��1�ɀz`v���"_�xd��4� D��:�	U��lK�k�5S�ָ��+D��0�[�.:n)XRE�6%���B@&D����͚9Ų� "�s�zu@G*2D���j��m�,rP��Dd1X4�0D�Ȳ$
�I��� f&�$UC(����;D���,JPUQr��#�.���:D�ܸ��8%���g�ʺz��l�7D��A�G�
hܻ����09{q(0D��7
km��K@���o-D�d����\`��iB a�X��+D��)�na^>U���,\f���`c(D�$h!F/m��@�D�`���'D�@�JǍC��er�IT�P ��+T'D��)A�W�ty��r��=xh`��0D���w�F��!�bF*Lse�!D�P�r��=ɸ����,B�-*��>D��c3A՚G�N��1�3�ĩI��&D��i KI7d�,4jQ���l��M9�g#D�4�/�M��%ٚ}$�)��n=D�`�c�hMND��n.�h��3�-D���B�)Uu�-����t�
�в/D��9W
��V=!��9U�K�/D��K�n	�xq��2*KV6��F D�����Ä�6!�vN(!چ�F.2D�� �ha�fv�ذ�p�NyPA�"O ���䁯=HrP��$0/�t�h�"Ot����F3^�bԍc�iؓ"O�`��(�lܜy6�ʠl����"OZ�aa�=WҒ�;V`T�k�*щ�"O��#��#HR@Y�O5D��A�"OERː�ja�u�D�ZR{D�sC"O��?Ӿ��C�$=��%�"O� �初
i�5q#ǅ<h�J|*G"O$�:Q�M$"OD0��H�xT���"O�%3�/ΐ �R���g=���"O:�sT,�#/��� ��f� <��"O:DD_�>*p�׏��a{���"O Y���
0n���Œ�]���J�"Or���ɢk��#��4\�l!c"OP��f͞�Pʂ�;�杲q�h�q"O�5`�a�>�� ���_p�pV"Or8����UD>�� D(Gϒ��Q"O�$H���u�m��k��E�"OH���OO�ih͚��^^�;�"O���&�U����R�E&�KA"O`�3�X;(Uΰ
�h:r-`��'"O"��҂�y��%Hc,�!""O��)-ԣ�8�%E�n��L�"O<�k��EmF�����_oBx �"Oj1�FITp��Љ�f�!W��"O`���0jw�uC#ۈwd���7"O<hU㙉q���T�].�4�"O$	:��]�:+X�{�e��O�Hzc"O6ar�X�1�n�y�ő�K�.�Y�"OD-��)%u���p����Q�:1��"O����0�d{P��h��0�u"O�}��^>!�$��7��^�P�Qe"OX�i@���NW��qRnI(���%"Or�� &.��T�'팿YQ�1�"Ol9�:Fyc&�X�A,@��"O4��a��h�<�C$�<3)�z�"Op�k1�3S��c���%A�l�8""O��
0Mݹaj�	q����p��"Oĸ�C%@�(�t���-vW��P�"O��Htd�0�H��$Dk:��!�"O���p	���sdF4bUֹ�c"O���f��� �Dޒq���"O��H��Ӕ 0Pp�_kF�}R&"O�QzDE�hV��%�,���"OL����A�#h�e,Dq��"O(i�"KHU�Y9e��L�P0"O�8ٵ�O���ҷ!уV(��q�"Ot���cɂV�^T^x���"OR ���:�Kڎp�B���y�Gs`Ѹ��]�yx �@��W#�y�A��6�<P����a�>Dh`�y�l�!�:�V��;Y�<��B�1�y�6�`8��!��OR�MC%�ɲ�y�F�iC�Ӌp��� �e��yb�*0ŀ�.�0d�F�%���y�+ڰ52�
��Z�MǄh��i_��y���h_�kgI�0��u"d�#�y�̛X����%C� ��% q(�,�y�E�y�8����=-9�#����y�<]p.y�Pc�<-���2���y� � k���#��"�ѻ��y�MݺL������l��As#�/�y�̏�" v�Cf�R��PR&��y
� �t��A�='R]� �(&��I"O�鋓�E�Fn� ǁ�c�\ͩ%"O�1"��>��-;B@�)��QF"O��w�)8�<ڀմ1�Ec"OzM3�l�6V����'B1 a�d�"O���EX�n^��I��\�@ZԹ*`"O�=���r'<��*��lH�t"�"O&��/V+�9hSJG�96e�"Ol����xN���t�,WİIYV"O�a!%B�W�x�d�׬�����"O��sM0J�Aů�*��tc"O��5������6�]�>��q�"OL�R��:y8��Vn�+���C�"O&ĊҮD;!�،�q���Pc�"OV)�hA�F@�e���͎�� "O �Y6K�-C8�x��,T��rpq�"O�|��/K8Em�0;��Ί��@�"Oz�I�I�g{��a�]�� 1�R"O�R���F��'�
0ހ�1"O62Qo��'Ǣ�*a)�b�	�6"O��˥�S3}>�i�¤9��mBe"Oͺc�ǅ	�l�%GЊc�����"OL��L�le��
 	��֐xg"O��,@6\O��2n�#	�D[�"O�U�G�K�]2��Gc���"O�A�v��2�@EsS-Q9N�(�"O���������'&8Tá"OfЛ4��O���eD	Vˤ"O�4L"z9���Sf�9C\��"O2�@#��! AD��X��[e"OJ@
w`f�ȍ�a�+�y:�"O � ������R�8ļѰ�"O��
�eM/xe�}�MY�"�@�P"O�m[�� Ɉe�͋@���{�"O�ʹ��xQ�l �5B�1��"O�#&͆Z$z���M\-^�:��p"O��;�f���!K'�-.���ybI#y
R�pB��.C���M��yB M�X��L��KŘ9���+�/,�yb#�$@:����Ѭ+*��ׅ]�y��^��V9A��ܿ | :G/��y2�*�	aקҰs4�������y��w��4Z�o �~������yBU�`���e���C�N�ht���y�%`P�*B�8m���sO�#�y�脉h�<���5јԉv�G2�yb嚛t�D`��K�B� �D�^�y«�m�Q3 ���oDq{e`ֲ�y�ǉ9YS�! ���x�p��T��yj�=U���I&�[�&�5��ƾ�yR.�� ^��aӱ��$�C�X��y�R�0U�T ��*�	�ԫ��y�$G�x!���#|����~��q�@���O.L��`WJ�'f�Ʉ�k����.ߟ��VW�,n�0��/�I�Ht&���"C�y�ل�O��8��A#NP�C`��aּy�ȓW{֑�f��	B���{��$W�\ɇ�6��Rt��6��G���Z>p���͊cK�?GjM;�kӚM^��ȓ-��(�&+R!GDxCp/�$��ȇ�5����@O�,�8��A�=J��ȓh�θ��o7&�¡'
,2W����Bt�h�2떑��lr�m�6��T��S�? 8�A�ዷd��I�[�n��@�V"OB�����P��Y8����Q*"O.��Kв0 �8����h(,�"O*MӖ΋!S��S%� Qo�uC"O|�"�'2D��1`E�8�$"Oza��=r��)B2ɘ�n68�j�"Od��¥��0���y!b��A'䔱�"O̀�`V�G�LY�7b32��"OHyU��h F���R7?"���"Ou�w������#�����:�"O�A:1�R�"X�hiAF�f����"Oh��""le�é�1.�^0d"O�Ac���,V�0��F?2��|�"O�頥\*����eB@(�vu�U"O��H �_���1�K�\�<+E"O.�p�Vv7^I�bCR�t��Z	�'d�=Y��Xr�5�E��** ��
�'�@ z�I��_ʬ���ۘ ��8��?�4�W�P& ��6I������V/@ʌA6�\�k���'o��'���fY>9��2B%@��P��%�`��Pg/!Ɉty�̀��91�M� ; �dc�
 ������
��~��UXW2EQ�` ���K�0LI�㌋jM��RCA0I���gl��t^"<���֟oZ�)I"��4��Sl���F�\!�|���x��'2�|����H��b;Y����2����Ō�'�y2̟�k��Jv��)|���B
��~�'h��n�ly��9 z�6M�O��t-���[:>�|�ǭ��J�(�Eה ����ӟ����K4��l�?KT<tP�)Հ#gV�ң�f>I�w*�6t<�+����:���H�-�F�H:�2$� ��PJĦuˀB�BD����b�	1�X��X�C�m,�O���5�'D��"��k��Q1��+/|X�H�	�l���ӟ`�?ͧ�HOb��D8��5{�A��]!\y�|�*t��n�˦�#?_Ζ��*���������Ԩ��A�Mk���4���a��O��dc�t,��^b$�����
R�1��E��2F$X@&�S��D�sB�|<������6��5�nM�4J��^Z�	,�!d=X7M6������2/�R}��C0;Hם8c����|�1W�L�CGט-5N� ��[n��nZ){�$�O^Xo��LE�ܴCh2�o�DZ:)*���RI$Q��?i���(�I |�V\���Je���8��ߌ,Q��<1E�i�V7->�S����#fI��K,Mz�D]MV��-O�y)W���
���O����O�;����_�43ҔWi��q� �$���K�D�'e�M!��	,ܣS�V�?1��/+��pj���Z `Ci	�`���q�޶4���S�iI�6�DB�ɶ~27�_~KP$��ڲ�֔#4�T��#��XBW⓪�?YbCO5�?���i�\|����O���j�hW����F핦e�d��	D�'S��q�l�5�(9��#�lj7�Ѧ=��4��������Ą ��qb��h 5ڑf�n^��*1)�6����O����Ob�jfc�|�&�����4��Ż�D!h{ZI8J�|����� ͦ2ڜ�3�a؜yɚG~�K�1v��%��7a��1� W�%%�śB�Dy=uS�N�|"����^u������O7�	8Sr��p��|(�O�g�<9M<���?�J>�I|�RAR2�<�%���QM��B'J|�<�bH&�"ਢ"[,K劐;d��m?�i�"]���W��,��<��]�UDa���o�J$�W��K�޵9�J��	ڟd �� w܆���D_�Z��0�DKC|���M�76H5PF���'�P!٧�������`��֨�jv�b�Ernd(��D�2vJ�r4���C�|����s/\"<9c�ٟ��I��M����� �ı�/V`}��9�
�6}�N��I[���?���?�+O��K�r�B�ƭ`�d8�D�C'�p>iV�i�$7mk��ԑ#MݮhY�s"-ĂXwB�`�>	礸�l%�L�>Y�"   ��   �  V  �  �  *  �5  VA  �L  QX  �c  �n  u  *�  �  b�  ��  ��  B�  ��  ۮ  4�  ��  �  k�  ��  &�  r�  ��  ��  :�  ��  ��   x
  R �  ^) �0 7 [= �C D  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�v�*���m���R �>�`�'�栨��¼`F-k��K��B	�'2B�z�� �g�-Sa��(AYQp�'�z�I��<2���Є;+fX
�'N�i�2���!'x|Y!l�Bq�,J	�'�P]q��Fd��4���B�4A�HR�'c�����<]6p���]�3���'��M�p@�^�0O�1cO~���'x[ŭ������5�J�T�ތJ���	/_�P�����^���z
Ȏ8��C�	<XMf4���7�Ȋ�>.���"O*%QQ���tKJ�	}˼�""O챪s~J�⑧ô ���;�"O8�7��6e�P[!�K���6"O^�
G��x����Ϟ�U����IZ>ˢ���2���:|�!��/D�8y��ξ_�|"ao�4]yf]2`3D�t�V��3S�:XKEJ�(�J�!�2�Ol�	��V��P�ۅL��9ҩg!q�1?���9�%�xEJt�N�iΌ!a	�*��Oع&��+����+��Vmy.�X�,��"O�����t����&��=���#��g�O�t;LH�a�f1���V7��P
�'u����K�G�|��F�څLʐ��'��]�B���Q�½�Rl��@��%��'�Դ��C\�&�������&�bu�
�'�rh��刯9j�`��
. �r
�'u(���S8,�l�A��h`1�	�'+�%��j�6pBHyȓ��$�b�'L�H�-�d��9(�o����l��'��P��Eڗh�p�օ_�OR����'�|�w*��x�zbF�2Aj��H�'GT�����j��I %�����h��n��L� G�x*"l�ȓ=�ʉ��kZ�yq�� 狁02��ȓ9sh=3�e�i���� бwC2���i�ڍb��cN�4��h���ȓ\d��C���(����w��9���ȓ
�Ȥ�B�&!k5��Hi��݇�c�:Uqh��%*�xJ���/�4�ȓ��y
��Uz���+]L���ȓ(C��ö#U%8��a��*j�� ��IE�w�b� g��k�����ԙ)DzC�I�:��d����? >����V$�"�\����~�dV�?�4L�q��7(��!�Fl�|�<� �af��UЦq���2~$���g8�D��ȁ���b'$.l"}2�K"D� �S�90�P�'�-��tP�."D��;d�*Em�\Ҷ�O�7�Ɛ)�G3D��	��p5�R熠�t%D� ��ϙ~Ȁe
7�N
nT�╀5D��I")V�C�TZ�-N�y�>ܚҤ8�	��p=�!'�n=&�Ж̝�x��U�R�T�'@ў�� n�R��1��b�3)U�G�Ș
�'5�u���H�rE�"�H���AUC-���)5���)ђO�
} ��U�iw$��Jc�t����.j�Hd�݇hJl�f��~�jU�މ{�λe>�  (��y҉]�A����T���ek�����yR�Ә.�Ɖ�+X�ǐ\2@��y��N?�jW�x\��Pp��2:����@`Xj�?Z m���X�h;D�,�_�m:��EA6@�J�J9D������8�艒&�I�%�TU�H"D������#�@�{uIL�6h
��/ D��'
��x*�iktM���8 �+D�$q�c�=Z8�2�O�"d�$�-D����O^+�p]��EM���r�b+D��pv�"%��qkuJF,9��U�$
)D�,�����Ы��³"#�I�@�%D�D��O�Q�P�ysd����8�
$D�H�T�ϤH��Q#�����
� 5�/D�(�4�8mJ�*T�G�\a�q�0�+D��S?j_L��5
ѻ1dR�`)D�p�T/η4j�,�4荝A�
��,D���a�>֞�q�i�%��ԣU�7D��F/�1�Y����C�*E`�0D���'+��!rh9Eς�U���!�+D�`@��� �p���@���Jq&$D� ��$J���� R�B�!�b D�hQeM 8PAJc�+F���b�)D�P�7cP>jH\`3&�ƭA8���#;D��J@�_��иȀ
E�Pa�T���#D��� ��B<z��C�_P½��6D��j���rl��1N�a��B�o/D�����v�T���� >�
Us��-D���o��NN�]R�%��:��(�� /D��Ƨ�>':$����+�\PxUj2D������\su�х �����:D�ԉ�J�r.��I��
tIR�±L%D��BPC2"(2`�N۟N���W�"D��:�IShW�]�"��'��(�#?D�0���KU��ЊB)<W�`@>D�,)�����K����J!��]�G(�+ #�"Q[d�'b��!�(�||�G,�1hY���ÁB!�$F���L�%'EpE���`�&�!��T-z(E�ӡ���d0�6AE�><!�]�% 	�� ЮT��%����7!����0�;������@�O�;!�E� �<�h�)9f�D��c�� !��B�N�.�c�GҮ6Y.�Ц�ۜ*!�Ğ�A�,m;�ƽ'F*� �>
1!�J�Z+��h!�X��usjG�!�dԁU�I�l��y�U��1!!�Πs2���:c�q"F��R�!�x<�U���(G��YC
�!�Β:���*�.;3�TӃO 5r�!��s �h���_/�l��n�&/�!�� "l����5&%%�%�Y+�̽à"O�a�Ǒ>|2T `�06h�b"OP�b��!L� $��ř=R�\'"O�!r�םi6�ȑ�T�@lt�k�"OV$q��(w�4���¦oe(���'62�'2��'���'x��'o��'8�E��͎�bx@@��L�Fk*i���'�R�'3b�'b�'R�'n��'̀4j�4^��3aZ��@H0��'~B�'v��'���'%r�'���'.~h��(ݮv�>���c�Y�0X!��'���'p"�'�B�'���'��'��Q������cr
?�p``2�'���'�r�'�b�'��'������k��GZ��9u�?\�`�f�Ɵ��Iџ��ǟ\�Iɟ8�	��Iş<y��V�R��Ch�>Zfz�hf(�֟p��ޟ��̟l��ߟ|��某��ş��S�����n��P�t�㟘����8��՟��IП �I������D��J�y���Jfb��LM9��̟��Iğ���������h����P�	������u��4P���8}A�m�e�����	ğ����P�	�l�I��D�I���� �S#�@��P���F���8�I�������ҟH����4�	� ��h�|y��E2|J�{u����iӦ���Oh���O���O��$�OP��._����`�.��дn�Op�$�O`���Ox���O����Ϧ�����[7��SS �iV�|����d�9��d�O��S�g~"�a���p�8Mp�����Zw7�@���&V�	��M���yR�'�v���*�6$)����G�H��1�'*b�F�W2�柟��'H�t�~r�J��4���i<���&)�H̓�?�.OТ}Jb�'�J1��@��:��YXG�J8��ƭ����'H�:�nz��+��O��JW�8W(Y��ȁN���I؟�͓����0I�6�v�89��ċ9�XhĆ�t�����b���Fmr��]�����'�x�8ց�0��æ�"����'��J�I	�M;�Wv�0���&Y�P�,�p��#��A
���>	���?q�'��I$E�J-*g��$V+���2������?���]	�Q�|����O�Q���!qd�[An�4S��ղ��h�ʨ*ON˓�?E��'\���&��#�tє#B�r�'J�6-���*�M[��O�DglX8EX��"�e�tR�'�R�'5�쒒n'�&����'��e�w�$aIg��"�س�D�^�$������'|R�'�R�'CX�˓+
�Pr!��5t(|�vP����4� ���Ӳ�4�?A�����VfT�%�F�B�����/dIj��?����S�'eI��'�bx=:J�_jl([E�o֪␂�<��,/]���B������\a/��;fN����Ӫ�a|�)a�N����O��&�z��F+W4��En�Ov�lZN��f��ȟh�i�)P�٢g�L9Ce��!q��"�G�s9|�lG~������S�6�O��m��_��s'�!mv�A5-ە�y��'����/Q�*�0&`�M��p�0X��Ɍ�M�PL�D���v�v�O����U�֑�����^�S��n�I���oz>�Z"N�Ҧ��'kr��Q��Q��� !)H�)�8��'�w�X �	��'��	����ӟ �	�b�LYS�L�.Dh������E�]�I��,�'[F6�T�W�����Oh�$�|�� ٓ��Ś��(<˘p�#i\~~R�>�0�i]�D�>A(���MRĢ�C�ȶR�V�s#V�S��t�DL���m{�h�<���
=P���#��8 �Y$͜No�Q��D�Q��0P��?9���?��Ş���˦� �i�*�<����*G$B�ᕢ�v�ԩ�'Q\7�/��)��d���)[�
D/L[�%( �ߓ�ܫ�K���M˕�ir�X���iw�I�L��] ��O��(�B<pw�ڡ>Y���@�n�H̓��d�O����O��d�O��d�|
�Ȝ0lR�����B97��	���=\���V�P�ן(�"��y�J��8n2E���e�����	 o7��)xO<�|"����M��'~���
I1u�b���@ٯx�.�+�'���Q�Fݟ���|�_��Sٟ���\�`��ٖ�S�1���e�����Iԟ��Uy�}Ӳ�p�	�O����O�	�`l[�l�"�V�ڵ���H?�	���D�O�7�u�I����5I �lS���j�<�h�8�qW
;M�P��|�G
�Ox���*� $�" գ����B�5>]�@���?i��?Q��h����M!'8D�iR�m�Lx �K�K����Dߦ+W" [y��t�J��]	Z����э6������d���ɜ�M�Ŷi�7MD�$��6�.?�7LL�`��܁I$�qѩ=RՊ ʦ
(��N>�+O���O��d�OD���O��j����)���uI�G1��cUù<��i������'��'��y�طa}���g>�� ŏ����2��pӠ�%�b>���U�Zޠ����R�U�F����B�c�媵-Thy���%�T����P��'��	�<j�׈�0c�*T�!�V���I�������i>��'�:6���,�d^20@)Z�M�UՏ�9fj��-��f���by��'g�oy��D1��Էк�I�hʭʠ��3!�L|�7-t����4�&���O<�]�'�t��� �,�0���
�+4�K<Y���9O���O����O����Od�?Y��!;A���0������"Ȑԟ��̟�@شʪ�'�?I��i6�'�n�����%���@AEN�\[�T�|B�'��ON����iY�i��AaU�Z��y�`�����i��R�R��	�' �G��<T�-Z�KH�?��S�o	$la��Ex�iӢ-��(�<1���	O"�nI�CƔ،$˕��(k�����d�O�6�D�|Z���5�A�/_2-��P���w>�I����)o���(O�	ݗ�?ɇk+��C�sTp�@���>1���t��=6!��D蓮���]Qo���I�+��� ��4��E��џT��4��'�0��?AeA�E׬�����DT�����?I�Pb�h��4�����H1o��@�K/O:i��
�.��0 e޿ޢ���3O���?Q��?q���?I�����]����$�n;}�#ء+	�mZ�-Đ����4�	^���8���c���"�0��͆s�z��pc��?)���S�'I��l�4�y2-C�|mjPNد}�֥�񫌳�y��W����ɘ��'�����$�ɸi��i����֒i��x�V<P��?���?�.O�Mlڇm��	������:C��P!W��G["X0��A�N̩�?9�S��0�4.��&�,��;
����l�)`�����E#S���S|�Q�M��F�Vc>=���'�V���x���(g��)6�ĵ���#$,��	؟��	�h��M�Ot��C4J�d�f��n��Y�a	��n ��l��b�-�<��is�O��>���F��@5�gC�f��Ѧ�����n�Wn�l�C~���= ���?_���e�/�:S��m0�X�|"V�������ܟ��ӟ��R�ċX��;K1�` Fy"l}�إ:�Λ��'"ҟ��'���	@�l�T�qKٯi�HR�B�>9���?�L>�|b&�ؿG�С1�[4	��� �MS��A��d 8Y0D	�j�O4ʓ*�0]�C�?����'�Y8]h�!��?����?��|B+O�yl�cc�D�I��H�����#ҩ��aŴ������Mk��.�>Q���?!��/�*�)V*��h7��c����
���Bq�W�M{�O.�2k�=���)3����t J6�ˁI"`�:��0T��<��9O��D�O����O���O�?����2���������@���(��؟��ش�>$�O�p6�4��?W���m^z��삓���#���O*���O0���c�z7-w���'z�� 2l��"��(d, ><T�sf� �?y")'�$�<���?���?�BƘ0IYIӏ*EK�@�c�<�?�����$�Ŧ��i�ԟ����$�O��ʕAH84Ku�i� .|R}��Oz��'���'ɧ��֌���. O�B);��Z9��5�Ğ<��jծ��4�LC��P�L�Or���ʩ=� ���A0Y-�%�O,�$�O��d�O1�<� �֣Ʌ A*͐V �-
��)���/.I�R�'��~�L�4��O���I*9�$�x�У�(�c�$vC���O���d�rӖ�Ӻ�NR#�z�c�<����IeS3kI�st��S�<�,OH�D�O��O����OJ�'Q|�����Q:Z��,I�MS.?�u��i�ndC�'H2�'��OK�Hz��nK)q�@@�'��=<*���
�-b���O.�O1��hzSIq���	�B�<*V�	.VP��'�ՙN&��I�b���r�'HX�$���'/�	�eZ���a�j�AB&S=6`�����Ϧ��C�П��Iן����@�"�Y� �ʹUS&I�g\Z�2��I۟X�It�	�4��1J� �"�<�Ťـkjl�<D�`��9S���H~�e�O������0�W'^��eD]�W��ȓO�6��k��9"��X�B��׬���� �������'i7� �i�MX%l��,y2t+w	�@8��Fy�h�I�I0��n�P~ZwK8�
��O�f���ޞ,eJ�C���/|�<��@��c��ny��'_��'���'�"M��*N>�H�OB	t&��Ӂ��	��	0�M����?���?�O~Γ41�\���Y�c:ᢔ,� u�T�Q����4zț��"�4�����ؔ���ѭh�+��)q������**��ݢVǩ<yRN����$Z��䓌��- ��
R'�����ҥS�Vb*���O���O�4�zʓ,�Fř�1%"-H�|������R	J}�b�W��yB�j�(㟈��O��n�1�M��i랠S7"@�V<��L��޵��OBv�F:O�D߻(<�9��"����?��]�c2��y#��|B1#���<.���Iޟd������ݟ ��L��S�f�P�l�EY�r�CȺ]�0M)��?1��-�6��7)��	��M�J>��B�/`4� C퐐К�B�aE-�'��7MƦU��!�x�l��<A�,�"�*Öp�<-���\�ʑ����\�"�D�����4�����O���B �8 �� =(䔓�.�$`3��dן2��p��ƢY[I�t�'y�OP�$�Ə
#�h�f�
�b�z6�5�y"�'��듙?�'G�����'R��!S"r��+H�N�H���[�.-��ZV'׬��	�?���'��&�(b��&)��MQ4dZ'F��yu)���x���� ��ʟ�'\ux�H.Of�lZ_�@��2(=#yz�1Ա!�$�c/���ɲ�MN>ͧ%3�I��MC���=d�PI�1�������K�Vdx�f:1mg��	ҟ��'�{B�T'my
� .�*��Eƚ�׉�/rՂ���1O˓�?����?����?�����i��H�lY�+M�Y� �b��s�TXnM�p�������	�?q��yj���Q�V{���bI�H��U8�
��_�����&��i�����F��6�e�x:��_f��1XW�ӛ9=���r�j�|a�j^t�r��]�Ayb�'�¡�&1����8Q�V�IR���T)�'?�'��	�M+5o�(�?���?	C�$�v����ؤn�LP��(T
���?�-O�nz������O^�)�cG2A'48�ӬEi$���5O�Ć#s�J��'	K)���j�*�O8�p�9���V�kB�q G�f_"�Y��?q��?���h���䛷<�����gf�Jˎ�/y��D�Ԧ-q����I
�M��w�,�
L�J�.�I'��bFe��'!�'��cV�/��֒�֝�bRy�S0.�5��mJ%@�,�)0�Y�J����Ř|W�4�	�����П�����)����[�~�I�3}�@�a��UOyb�p�v�i��O|���O���x����l��F�6rѪ1C��>���'2R�'ɧ�O��%�'I	!̥;Ԯ�s(V=�׃�#j����V��XUA�cH�IJyR/��obT��3աfd٠�䊦^�R�'���'r�Oz�	�M����?)4��=U�m�≝�9��F��<!W�iY�O$T�'v6���ٴ�P�oV�l��)�흺"�z��ȝ�M��O�D�a��"�:����wLE�n܉v�<��5��hyX���'�2�'j��'e2�'�񟖸��g��S�*n�B� ���O@�$�O��lZ�T,�'��7;����}p����;���k����S��Oj���O�IH��6�??��)�	:�dG�a��)C�h&�4|��� �?I�5���<i��?���?ɴ�0Z"��#su�����?�����$զM ���͟d������O󂌃����{�fO�V�Ȥ2�Oځ�'f2�'�ɧ��ݨf~�0�%��q������Cڍ���)RM�18  �<�'�F�����%���@7�H�>�n�ˀe�%�ذ���?i���?Q�S�'��D���S�IZ�y�e���Z�\nJ��3Φ��'�27�/������lӒE���E�{E��� 슾qh�
� ğ�nZ�cd�l@~�V�"[t@�S�8|�	0�l�K!�o�X��Ug��K�R�I{y2�'�B�'��'Bb[>�J Q;T��P�'ӶjFz��+^��M�D��?���?�M~���-Û�wD�	�(�ug���O���,�s`�O���<��O��D�O P �i�d@�D-�a����1�R73<�Բx������O~��?���.����W�~�!Qoɐwmz%���?y��?I-Ob�oڂ,n�H�����	�r8�zA&�8��4z�Ø�)A���?a1W�0rٴq�x�(�.L#�`�?PORи��D������b�⁣�ꏉkւ������n����9r�=bv&�^�\Ф	[�u����O��D�O���.�'�?yVGMFX��(�7r���v��'�?��i�&��^��޴���y�E�+2F]�ã_�v�l �I��yb�'���'���Yd�i�i�I� �?�"���*z��PZ'h�%sBpdYB͡H�'G��������p�I`����fce��r�}0��
�(,��'�7�O�MW$�d�O��$'�9O��b��Q3��
�!,D�x�-�f}2`v�rmړ��ŞU�p��I�=�l����?1�4i��ݙ
�� �'f�� ���4�|X��2���-O�X�"�K�~aD�C3���0�	�����dy�/zӾȣBF�O&���
H1{�j�A��>"ء&�Ov�o�c��&��������䟈�,WT��i�%AԵ��J�/�l^~�<a� %���p�O�''/>������q�m��LQ��y��'���'���':b�)�%܄���Ē�B�[�!E,X���d�O6��B�uYq�SpyFm�0�O�a����L~:�R��D#"���O>���Ob���O�EboӞ��`��K�: �g˱tK��ʆ��ܑ��mq$�O�ʓ�?Q���?Q� of��U�ݹ3�,�(G4����?�+O��oZ�zdPH�	ޟ ��[�T��B�ekX��$"�� ���x}��'�2�|�Ol2Iņa�ȭ;	Q<*9�0 ���TF�R��+W�P�%m'�N�h����+^)�����8	�M�I�����4�)�ey����5�d%đ_ �:�EZv����L�1VF����[L}r�m��iHүZ-a��Ș�  �@��#@�Ʀ]�ݴc�@��ݴ��d�-,��Ġ�����9�M���� �� �d�[e������O0���O����O����|*$
�Jys1I��z2���A:nm�(�o,��'X���'�86=��Aشo��7�Q`L�#u�~}��\ğ�o"��S�Ӥi1Yo��<iS��̀���-9����V�<9q��wS����0����d�O��Dסh�2�n _�`�i�`^)H�^��OL���O�˓\��fMb�'�2_�hĲУӨG2��cd��B��O ��'D�6F���J<qU!��h�rMs�(�)Pq�{ӅZI~�"фS���T�K4*��O���	5*�b�J�n#|%��O��[j4�D��'%"�'���'�r���H�,��D�'�\��!h�	K��9$KW�B;��q��'��7M�l�$�Oеn��':�w�c�	��p�b�=R�0��'Y�f)w�0�oZ�:m��mZ�<)��/������ڱ� � �!i�9�,xQ I�&EV^}2�G$��<��?����?i��?!¯0@���R�F50�
ia�����$LҦ1�#Hʟ�I۟H%?��O� ��ևP�8�`�ju�ӿt�P��O��$�O��O1��(V�Ϳ"� 1�$�X�W#f(�T��s���{�<���X!N���H�����T�?QP���dE�5!PE"U�ӎM��˓�?A���?�'��$Z��!U&�蟈(ኝeg<�K'� %o�
��Jo�0Z�4��'z�˓�?�4�VB�u�4e��I~O�AB. �(�"�J'�i.�	� ʢ�H�Oܾ�$?��]�n�ĩ��ߍt=������>��ڟ������	�����F�'9�Fi�R��12�������l���?q�3#����r�	%�MK>q�'�{r8�1��ەk���� |�'Y�6-�˦�39��n�I~���(+�
5�S�ҸCG$e`Rd]8$�j��6ΐ�;Đ|r^�4�Iٟ�������G�,T�*��_�v��G�X�`��_y�z�jhA�O��D�O~˧0�չf4
��H�O$����'��d��*fӪ�%��6e�-h �\�L�����=�<EKS�˂{�����M��4������6u:�OB��&@h�l�jr%'[Ӻes���OX�$�O4�$�O1�`�Lӛ��ҢP�ĈrĦ��7���w� P�l�	u\���۴��'���b7�V�@�B5�5�̀7/�$u�����6�����9�% �͓�?���Z=o��	ۍ��D�c|.Dsw�A!�b�*A%� �d�<����?i���?���?�(��Ų'�*_��XuGӊ>���Y�]P ���x�	۟�'?�%�Mϻ<%l,��`�?Ida�f���$^��C�'��#����K7+8�F?OL j�/�� �<YiSÜ<}	�T�f7O�y���P�?���%��<a���?��,��\CK� vr�{���?����?i���DD����c�˟`��韸��M��*q �3t$P�8��t��JK��U���M{t�i/�Oj�'��p����H�06��c���4{aPt<���_�S�u�͟D2�!G�v�Ջ�ɧPUصh� �	�x�	ş@G��'5\�`R�ټY� t)�i�	*�5҂�'�7��"D6�$�O�9lC�Ӽ��"��x#l�� 3G�<)��?���jy�ߴ�y�ڟ�����T���CE�)�ycc�ËP���j�ɚ������O����O2���O��$κY�v�uН�����,Jlʓ\[�F���&\2�'�r���'s^ܺS�*|��
���-�~��Q�>����?�L>ͧ�?����!YAap��t�T�M��@i�(P�/T�@+O2	�E�"�?AP"$�$�<�dITV��u�Զ:�:�Iܜv�2�'���'��O	�ə�M�"*;�?�D&tŶ�H�C��J�pIԤĴ�?�P�i��O��'K��'K���?(����D�9~�]��d�F� 1�i���:X ��(d�O�~$?��� ��97��LJѢx
buC;O���O>�D�OB�d�O��?�#I��xa��p��ɫ=��A����IΟP��4X�Rp".O��n�e�e�<�PQ������!*<Q'����֟`�I1%�x(n��<!�O�<eP'L�DL1�K�J���[��t�@�F�ICy��'���'/�杼y%h���s�|LiңҿIr�'��	��M�D����?���?�)��!q4lG�D��a	�,C��I������O~�$�Or�O��#5�v�C�YE��O9�h5RnǢI�B����Wvy�O�"���0_�1O*uT�P�	���k#j���'$�R��)��_yB*wӀ��g�S�zj�1(q���_��0��ƺV�0�$�OޙmT��F�	՟���[9Fo��yh�3(�N��Ϗ㟜�Ʉ�n�u~Zw5��iw�O�N͖'��KQQ&�ʀ#�-�I�R�ў'��	��������I���	g���G+�)5�ɱ�L=�fb`$6MR�F�����O���*�9O>mozށ�d���ywa�3xF���#�M�p�iw�O1��A�k�`�ɡ+~��$U�(}c������Ɍ�R=�q�',$�,���t�';(M� ��NY&}�C�>~'z����'9��'bS� ��4[3B�y��?��r���tHX�p(9�!�A��5z�B��>�`�i0*7��F�I:�D�K2�J�k�dx�Т؋)���>�ȘA�*S�-�H~B#��O�-��cET���Z��h�c�+Ȳ����?Q��?���h�����Efۧ�%9��G�0	�����������ry�`k�|��ݵR}�@��H޽X�D���&C@���	,�M�2�ict6�C'mX7M"?9�#Z����)͘bH�8��ɪ������f+(� N>�*O�	�O0�d�O���O�8�e�5sgtES�HąA���K���<Կi�n���'J��'���y�&��+r�ts�ܮ:0��g�
��B�'�f"c�HY%�b>uˤ@̡0n�P-�-89���� @|~���X^yr�W% �%��c2�'剤:|��`�l�-a�̹y�e�*\ �	ןl�	ϟ�i>ݕ'6�Vp �$��=�N��
"�4�V2��8ϓn���dn}|���n�
�Mk�!�$H~����,"��e��k�j�j�4��$1��m���i5������Sc��ԘB�[�)����tJ�����O���O���Oh�>��5Q��í�Z_�݀�fךQ0�)�	���I�M�1��=���H�9$�8:�n�4Y� ��1/�-S>	�����[[�&�{��V�(76?QtH�n�? ��Y���#��Pk?�ּx�f�?�A3��<����?1���?9ŀ.V����_�!θq5���?A������˦i��O����ӟ��O����)c�A���!5b���O*E�'�7mԦ�;N<�O�2��"��w�̍�$�2�vL�v,Ù*��9чʜ	sh�i>����'#{�'�x�c	�0�^�q��X�0������'�2�'P����O~�	9�Mۗ�yt45�C�s�y�BJ��)��I�/O�Mm�V� s�ɴ�M�F�J"F��@�瀖�M�z��Ċ�(u��{Ӑ\��`cӤ�E��A8�`��p�@)OVTA��P�t�v���Q�B��A;O˓�?���?���?����IA�2�R\�L̿
WօhG�qf4mZ�;���������I@�s�"�����I%���S�@�ʅ�ǌ�)�R�i`N�O�O�};��i��ħPXd 3�o� %ׂ00�G��W���0n��j��}B�O���?����~xh*��`�d�22ƅ~,����?I���?�.O4nZ8uhu�	��t�I�D��)��՚'	Bu!�	�w%���?��\���ڴEM���(񤃟[���b�*]�4���;W�����I�p�Hu��c];.c>� �'.q�I�h��$V�N�~�$��=u
M��柌�����\���?�;2V��-�&2X�[��v�T�y����aҶp���M[H>y�Ӽ��OF��X��@�X. �������T?q޴���D|���`w�h�Ɵ'Ou|���X�F����c�r	T�"���-ʈP%��'U��'X2�'���'H��v��2�`!��^�.`Г�Q��jٴW:�q���?���Z���?���$�Q���w^0����]{�d3����צ������|�'�B��>���z�/#D��r_E0ʗi���$�1@lI��4���Oh˓�v��L/^�1��܎1w:���?���?��|B/OZ�m vU��	�R�0� +���@�&��wg���ɴ�M�Rb�>���?�;��k�b#�@]!rş�X\(�5@צ�M��O`���F����.���� 0fE�
���9�	��El��9OV�$�O����O���O��?y����ԥ�$�wR�<���ן��IٟP޴':��*O>oZt�I.
��A��!��(��*���H<E�i�6=��j��j���^P��`��78} ��񬀞#����p���x����䓀�4���$�ON�$
�����h��{|R���[�?J����O"�r���C9@^"�'�]>i�p�:LiH#�?����P�<?a�^����4-��!�?�g˖��F��RS���8q7�9p,lI� )ӥ) �m����B埔H�|��R��R�e��m������ 0L��'���'����X��ݴ'�5`��)]�>`#��ߩ�@z5�N�������?A�\�lڮtcB!s2�G��l��Ѷ$���B�4eL�F*4��Ɵ�8c���1����"�<ɢ�Qc��#c=D� F� 8P9�u͓��$�Of�$�O����O��$�|�z*%K��?�����oM�-L�FI�4d���'3b���'ɰ7=�x�ȵO�9���A��Ht����ϦI�4$���O�&a�c�i>�䞺!�Q �oA�A���ąAX��,�[��B\�O*��|:�y����U�Y��yˣ,�ɞ�s���?y���?�)O�tlڴ*��5��Ο��ɶ]yr�C�Hج2�t]�Չ
�r��e�?QP\�pJܴid��xr��D
pH��f>��Pj������ |��j��j4�����:�o4,����]/ܵ��n��I��"�K<C&���O���O���'�'�?⊗�?�N�І��f!�`��*��?y�i:�%��\��r�4���yG[��P����w'�Iү5�y'u�b�mZ	�M�tLݲ�M��OB��d�����`��v�D��I$[9��S���8n}0�O�ʓ�?����?���?)��RG>$3���D�@IӣV�� P�,O`�lZ�NK���	�(��`�s�8w��,�@��3Ӯpz0�����DKʦ�J�4O���O#.H��͉X5�Fo8Qt���a/#~�ވ �W�����;]�rM�	zy�G��<�:�kުJ�l9�]�ug��'���' �O�I4�M���ݺ�?�Ěz3�k��*ouƙ�ׂN�<q0�i��O���'��6�˦uڴqz��nɿ��ȋ�O�,���l��Ms�O\�h2���r�/)�	���42B��
b@�St���:.�zp;On�D�O��$�O����O.�?����	F�ʑ���6ep1�cY~y��'��7�3����O$�n�x�I/+lm٧��^�dݸ�дg���J>��4fΛ6�O<t�ZQ�i��d�O~Y�a��!`H�0���(�Caf¨2M�R�Þ�O���?���?��j��bI��]�ՀX�<%�i���?)O�$lZ�<d]��ɟ��	_�k�2@���⃁��5>r��!iՍ���Q}"Mu���	^�)ra��*t5��Vܐ�(�#!2xME�vϾ�)/O�)�4�?���5���8:@�l�!�,u0��� �����O^���O����<��i��D�1��u��JSV$0��H`�	�M��"J�>�t�in���A��:�X81%C�E`�9Y�@�OH7�P x�D7m??�F��j/����"��ՠm�d(y'�Pz��C������<��?q���?!���?�.�@(P��ʞo4�a[�BP;-VFq� .�ɦ����� ��럤$?�I�Mϻ���0�0IxZ԰�N�������?�L>�|����!�M똧� ܵ����Z��B66��В3OH0�B.�7M֌�`��M:}��c�(��-���ί�DAّ%ּn }p�	9H����g��J�R���� )���#�a��MΨ
Ǯ��C-�ݹ`솬bZ�0ł$l�Ġ��a[Ѧ���$�5G��y"�;C��!$��<)��I�� Y,Q�<2� �  |��P���{�:5���
�BOJ���C�~�P49�N�
h�ʍ�2%��E����H�Y�|ya�+ӧ'��9�L�B��xH�\�-j� ��ip2-�'ܮ|��lCb��g�TY1�P��G�R8�p�#�c).��T�ǊZ�EX2���eg����OZQ�ӎ� MFW��/�A��dȹ=���'��'z�ɸn6�c�Hxt�S�vnl�E�K������n�l���O
�2��8z����'l�t���j�����fY)���ሊm� O��K��TFx��2=K�O�93<I� .�cL��#��ih�	/6�4�y�4yy�ٟ��S*��DKq:����O���.�sI�Rw�6^�pAe1�S�'V`x��/'���2E�Ҹ6-�2nw��D�O��$��P�&�L�IǴ�h��><���e� h�l�iڴ)�pEx��i�O�4bR*Y�\�Qcȳ6�<5)ք_Φ�������`����I<	��?��'��!�آ<��y&{~.�Ј}�唘Ԙ'���' R
GyY���)Ex��(��P�.�*6�O �k�R��?�K>��id �&�?J�~a)�O^1'�@�'��`c�y��'�r�'��'b_��g�d��@�%ߪC���"0�-���?���?�*OR��x�`�,��Svxijq&��W<����_��?y���?1-Ov)�����|��!K�wU��C�Y/O�>ā��	�0��O�Iqy2�����t(��ab*��N ���;1��	۟��	П��'��Tjw!4�
7O�8���'E��+�fAQ�&�n����&�H�'�̵x�}2�7t8VQ�g�+c�ܜ�R�^�M{���?y-O`e"���z������?t���+W'dk��MC#L����N<�-O�M`�~4����	���Y!8��A娝˦Q�',��DfrӲ��O���O� �%�I2#��OL�1R��m�sy�O��O�� Yx� �S��H2'��pĦ��1�iL��)��s����Ot��៨u&���	#h����77�ju�-�i�nĘ�46
\�Gx��)�O��P'��1zN�@�K�rު��V�զ���ȟL�I]��@��OL��?��';H$�AO��;�TA��� Cl�ٌ}cǃ5}�'eb�'@� Ǡ#�8�H������Ă��{7��OZ٩� �c}�P����V�i�ѣ��R!:M8�o�6�`���>��c_;���?y��?A.O��2挞]��ȫ��^�kq�4qc�N�A�x��'��	��|$�h�I���ۤņ'�LI;�D�o�}��ģE�hH��ny��'���'��ɣ7�B�A�O��	a�����p"ƴX�>�h��ۦ�'�|��'�J��=����lb9+�$C(L�܈��0��I����	���'�&p��~��lb�ڲT	6�.	9 a�'�^�c��i��|��'��@;qO����÷{��O�7Y	Ѕ!�i}��'=�	!l��R��r�d�O���Nh�,$
F�F�|��H{����yy��x��'knPD�O��pW�m�3 K)0&4P�M�9{�7ͪ<12$B� ���'R"�'���L�>��b�����L�/&~�4�TV��Do�����	K�d��?��D��L�����A�=��);r�S.�Mc?W��F�'���'|�d��>Y.O�e�D&B�VT��(J
�m&q��	զ�P��{���O(B"ڮi�zm0�%ȋ\�E��MS�Br�6�O����OcFH�P}�U�(�If?����([L��Em_�.���u�A��|@L>Y��?!��>�J�b��_�붙Ȥ�Y�f�`�i-�N��Qr���D�O�Ok̅2_����W��L�$�#�4w��$ltTA��Gy��'���'剻Y����I@�2�r	�bψ/x�	to#���<	�����?���UE����Y8��Op$3f����?���?�)O��P��|��؎w�`Xu#��jz�!� �զ�'�"�|2�'���"F%�âNr��P���p{t��я�4�������ɟ��'h%Ҁ /�6{<�S�ǘR�8׬�=	��o�џ�$�ė����'��'e@l�A�[�S��q��o�!5�J�o����zy�
_2Ȱ����kl�!,l(�K�\�z�Z�
��
�nʉ'�������@�s��]�	�䉁��	� �<ar���7�<AMt}���~��������] :��B
&}�`zsa�ʓ�?����O���M[�cQ+|n���J6;���/���	���͎�M����?����F�x�O�Z�sVT8t�T�pmV#VX�J2is���$�O��d#��?�k�l(�ҽ:��X蒪�"��Bĸi���'E�dU,T��)"J���#OI68n�Ak�.U�k4���nM��O"P�~���~����^�Ch���Ӥ�Y�MS�'!�	�,OF��O��O�|C��[���#P�8��u��
�^����b����My�'*���m\���]�T�ʍ��J(��	���Iz��?A�'���S�1%P�L�vlG�h��u��4� �<9���D�O�a�F��?����5k�	ۧ��"i,Ή��z�����O�㟸��zybN�R>� F�	E�U)q��p�J����Ts[���	Ο ��sy�K�9�\�DQ�T#��nM��	��b����a�Iퟤ�'��'�����' �8���#�]q2��V�[�j�@�o����	fy��;����D��kp��r��O�B�l4CK\+/��'��I�A�8��H�SW�V�5��Ł�M�["Fp�2��ΦՔ'��A��s���O���Or8�2ZT���ܭ	�ǉ�#�)o�Ꞔ�ɓQ[ �I)�ħ�j+�����*/�e��C�m�|u�Cfύ�M��M7�?����?���Z(O��*�d��Q��)=!ܑ�M�33��İ�4ebd��R�[D�S�O0�臃����N)I����EA�HUl����	�S�����|��?��Lw��C�,^�Á���I֤�ݴ�?���?qť��,��SN���'�d�#�\�0�">ذ!1���)���1Op4�FT�$9����G�<TF�\��Ƌ�k��d�a�����%w3B����O�ʓ�?��A�)OTT	P-�r3h1Vɀ���`�*O��D�O���I۟
�끚xw�59�o.gQ��(��A�$i�Tr� ?A��?����$<dR(ͧi*8�
�)S�v���2�̛K��lEyR�'t�Iş`�	�p��>�$��.):���$�+6�N�q��Aͦ��I՟T��۟0�'���Z��~"���-�50�1��"A��a� R��!��by"�'���'B�K�'w�s��ip�#XI�h�8NYt���@�i���'f�ɠ(�6������$�O����l$�Q�h $Q>�y�w;v�ܔ�'r�'qR���yrP>�I[򅧐�k���0B�(8�%L���'���p�(a�V���O��D��(ԧug�ֆ5^V�@���&Y�G�D �M����?I�l��<A(O&��'F+�
��΍m�j�3�:m^6M՝[�D�mZ䟬��ן������d�<�  �V�JX��H�.\?��I���8\��)�/�y�'+��'���d](G��D�6"0��e�W
U1n3pumZڟ�������M��$�<����~�K�7!D(8����C�M3���$��?e��ܟ��	�7qF<c���>C�
p�ܯVX����4�?!�@��<��lyR�'j���X�2�R&���~&1	�Ĕ�r���WF�ϓ�?	��?Y���?q*O�y%L����
P�Q�3
8
P��0W����'���ßĕ'�B�'��@� {��g��-@h�2�O,���O
�D�O\���O˓5	`ո<��i*v�ڡ墭@3��&Zp��A�i��I��'���'� ��� /��P�N�z�A:��7)`���'�b�';2U���`��i�Ok��7Jo������d�ִc��V�Ld�V�'�I۟`�	��G�����M�7���J���KgEՠE�,m��Iʦ��I՟��'ϸ�׎�~���?���
/J��e�L?!��sQF�1w�}[�P���˟��ɔ<��	Q��'(���h�Q�M�,^h��@��_��]��+�@3�M��?Y�����P��]4A����ucF!b�~`��A�!�6-�Ol�DV,����OV˓��O���"b�t��4��ˍ�sXTݴ1Nq��i���'T��O6�����Sd�d�G����D�D!�@@n*v���^�I]���?i�Iގfy��q�!$SA�a2D�<n�v�'fr�'^�0���>q+O~�d����af[�Y�ziP��D���j���d�O,�$D<��?�IƟ��əm-�q�&O�N��M���-�|��ڴ�?	�.Y�#��xy�'8����؄?nlR�V�\rW�4t̊�<
�p�����O����O�ʓCBV�h�&_,F�n�Hr�2'jؙ�D��Zk�IPy"�'��	П<����X�!+ĺ��;,����aD�%v��	yr�'0��'��I�;!�C�O����#�^�6i���ZDw��ٴ���O���?����?q�i��<ٓGQ�GZ\�P"DV]f�K�G�3u*���'��'�^��hf����#�eB�:-����i�)�����R�	ܟ��ɉ:�	P���A���U��7<J\ɄL�*P�V�'��V�d����ħ�?���I��%�U�'= a顢�B�\C�x��'�����y��|֟�H�,���Qh�:mY�e�V�iQ剃6D֙�ڴ|%��ʟ������S���p��R�o┑ҭO�!r�f�'o�J��y�|��IԆ);�y��`�!#d��
Q��%��gZ�oc6�O@�D�Ol�i�C�+;4(�T�ކ�zu%�tc��p�i�,�?YM>!��t�'�14�0G&q�m
�,[�0iӰ���O��d�| V,�>���~����Z�C)h%�� R����q�i��'����2�	�O6��O�]�Dφ&PR� ����G�r%�u�����I�k�\�jJ<���?aM>��t|lt��n�=)y0�ū%H�'xjE��'��	̟h�I��'�j5�E�χE�E�G��"�׉]��O4�d�OړO6�D�Od� ք�
En$���C��IBa��z���<����?Y����$���̧P�$�����\�8��f/P�{a�u&���	d�	ߟ��I� ��ɤZEN����8�L�h'�%��a��O��$�O��$�<�A�	f�O�(��@�|`�qѡ��-���z�'o�X��-�d�OZ��Ͳs>��6}�,��2/F܋d-�H���I�HG�'��\�X2�
��ħ�?1�'ue�4�skΛg�`!��(N�!�$9��x"�'Br*ۂ s��|b؟� �\��$V�{3n0:JP;F�:�{�i��)j����4�?���?���\��i�鸅�0)?^��$�̖/��9kq�fӲ���O��xs0O
���y�I��$04q���F�4���Y�^��o٧m~7M�O����O&��o}�W�ȁ��9Sf�݊���?-*X��ׯ�Ms0�B�<����<���03�
;����Th;A�����$���M[���?i��X�� � _���'���O�l�����N@HpW �.� �&�iW�Y����{���?���?��f.�Zy@�!�P��,#ěv�'٢Xy���>q*Op�$�<y��SCmܞު�����pQ�8Kv���9�	�	��Iן�����0��ǟp�'[h�C�"~��@�HD�bqSP�ٖa������O�˓�?I���?1�-�!>4A�W05��)�g�u��������O����OBʓ#t� :��=� lS(@�QX���	6��(��i���'�'�&A��y�A�f@2d*�Z�g�a����F��?y���?!-O��  ��p���'A2T8��/Q��QRL~d�l`�2���<����?���F�P̓��I�[N�S�쏼e���P�πK�.7M�O����< �Y$�۟�	�?-9a�[4w�x$ie��r\������O��D�O�ݻ";O����<	�O��ٺ�M&�Q��0�81	ݴ���[�s�<�l�����O���O~�K�����`'Z�}l�	k�C̩�M����?	��I���'8�L<a0ȇH҈Q�;P+v�R������%	ݟ��	���I�?��I]�	�N�	BLك"�~��'gЉ��ܴi�����P�S�O�&�q�9,j�`��g	�!���C�i�2�'�2�� c��O��D�O>�	�CQLY ׌�H��KQ.�	��c���M-�័����@1U�:���Ys!I�2H���aT#�Ms��Z� )d�x��'�R�|Zc�L �CJN:z��`u��]j��O�4Ku�d@6'nE�UE;�!�:��3hX�}p�R�.Z�D��C�	�O��i0FP7�hL�v��4�>!��Y6f	0���m*l�ɑ	��E���j���@Qڸ�I�0e�Np*R���)��`�'� {�\\�fjg}E�!�JR�%�aG=)�DI{B�G�*�D�ƌp�TB��؈=���4��}�f�J.Bf��`C�
�A��ь
*l[N!�W����@�˷��/ި�Ů��hضi1���/ =jM!�%�.}��m���'Z��'NBPsԉQ�x�z�Y�c�7 3�M�s�Cu��g��e�ШU��6�_�I�<c����@�ca.��04�T;�4~\N�c��c�譨�Yx�t�@p��>8 �DGyr�N4�?9���OG2����n�\p�X��	CԬx�܄�ɷ'�v�kT$��V>X�$I��WC���$�Z�&Ƒ(�-�c���(�O���	,X):�O����|��K�?���?��P,Fp������=��PA��U�&��+�!�/�J���Υ>�O11�r�զO�ZY�Fܺ,�%�b㈼z���[�L!-��(Z}���'F��#�([5O�&��b�W���y�g��="�2�'4�)�	 ��ʕ
\�	0�OJ�1K-�F��A�!��6L�0��1n�]!	���N������?�s�O�C_�� �ȏ	bDr�������/@�t#.F��$�IП��I��u�'�"���lƱKc&l�X��bdH�dl��d֠O���wK	�	#DT ��hOF���)�$�>�R6"L�
�����	П@3��3R<����Fs��	�,�t,���a���`�L*2���	Q$����O0�=�,O֙�G�@=��D(Ӽ��4$cIx�<i`,R�eBt��p']�J���1y9����ͨ3�m�N�l�J�/�kv1��(E�w�D�I埴�	�4ɣB�ş�I�|d�	D�ѧn_�A���ؓE��� ���-H
i�l[��<) ��(&J�X��M+�}� q@�RK"NT��dY��<�b�럜��$~N~@A@D�7?I\�@
�
=D�F{�	pn�Q���	_&-S��@�SGC��-s�bc��%o����,�"Tj��	���d�<�@i�)#��f�'�r\>��dӈq�P��Z�&ݪG^'
��I����ɩX�.���W��꓉-h��9�4ݟ�AQf��/�� �v���&%�����I,|��eB6�v��]�6�HcN�䦞��n�(uM���V�',�hI���?����?�(������F��)� �ppO�O|�"~Γ)�0M
PN�Od\���L٬9��@��ɲ�ē_F�JPB�(zkV�:u��+R����n&u���i��'���h�t��	��|�Ɂo��pE��TJFٙ�N'9-�\`̄;k�~�N>�Ok1�҃N�C��l�M�W44�3�P=N�C'j��
�O?�$ˋ(� �쇝�����!����"��O����O*��+�矘�%�Q�"h)h`�@3l����'p���	Ex�ܲ���b�
1&.g�$����2� ����z���	Ge�^`krOL�^�R�����?��eܶL*���?����?Ib��p���O>�yȂTޮi���ɒV�n)�F�O�[U�'!� C��:��"c��3& $8�'�E��S�? h����'&�(@6#$,���W��O&tj�*�O*���O�Y�L��yr Ć�0�90	��^�H 3d�Ą�y�(�J�	0u�^�Q�X�/�Yr#=ͧ�?����Q$<U�e��L����&�W��yR'N��F-�P��1pQe1q�S�yR�Q����
pd���ר_V���'�`�@����N܃�F5U5��C�'_Z��1�]�{|��[��
b���<Q��B�2����`̑Tz� `Iq�<Iƣ�.�z$�*�	"��x@s�n�<B�T)�p{�VL]L�	ŎN�<���}d����)K�y��=�rJ�a�<9���!���B�",�ȴK��t�<��E���H��'W�j�,,�w��n�<��Mق&�j�%`��-f�I��i�<�t�L�!��)SmR�qv�h���f�<A���9���+5��-*���P��c�<���� (��E�i�j�z!��i�<1ש��[W�|�!O�DC���q �h�<ydlL�I�h������Ӏ��g�<)�l��xvp��i@_� ����M�<�5@�XN�X2J�K��=�%��L�<y�ܑ���6���~ɺ���G�K�<EL��n�|IEO~�E����k�<�w��r9�0��i�B�E�p�<!wb		���"%�Ʃ%Ȥ�@�CV�<1`�+�<����ae`��u)�U�<�+-$���(5MR�tD�H�O�{�<q� �eR!���.,�iv�
x�<�'#��-�pƋ�E��� ��Y�<�vn> Y�t�7 ߊjI���ǊM�<������
"l	[�y�d �o�<is�lX�$FB�ps�`��eR�<��ښW#p����t�h���Fy�<1�ŋMbip�#͝/���h�H@N�<1��H����ޚe���^A�<�u�áMH�١䉝D�
��%Sz�<Â�7En��u�S�v����k�<q�/� m��\CTiR�F�j��Ki�<����!k�h1��^�*�����L~�<ub�<�Ԩ�0��@�6ǘn�<A�`۹|^�؉��XiL����@�<�D`�&���8����M~�{ b�A�<٥Λ..Uh%{s�,2+�F�<A�d�Gj�hP�!ʙ<�����c�<��K,7� �;�!��e��(���D�<��遡+*Ja�ꃮ(	��(*��<!��(U�(:&%~��|��/�W�<IDܩ*F�� �7_#X�`c�T�<�
յND*��E�|�zq���k�<Q󮃃u(��2뎊C�^�@�Qd�<1Ѭ��ax֩y�j�Y��ݢ��c�<�r�U�6;�����k�rU��j�<�@o��eP�ť֥wpn2�+�d�<���+H#0�� ����t�H�<�!��P��]
�r�q�Yk�<�#� ��$+� �A��P�c�<-^L�#�(�U�\(`IO�B�I	僇�
paX�(��&PB�I��i��e��W���C�c�5��'F@�H5�Rq/��fY�K)F�
�'�<x��\<K�T���ݱ;�J��
�'�`jɇ=�t���`Ґ~挰�	�'�0��@���� y���J������� Tp�@�Q,��b���a��$)%"O�آ@!H�2A^� y^Q�%"O��酃,="M��*w�i3"O�y�`샻P1��TE_?k�A "O�2̎�����A�ƫ2�Ȑ+6�6D�0sj�4-e|y[��֞����D2D�0�V��x.�![0�
=2�,���%�d2�O�M��H�#��!
�:[��ا�'Z��C(�>��Gs�Ѓ�۲Yy�,a���~l��R�>�	=2@j#<%?=�U��UP�| "��Q]4-B�=}�DM9��H���'tJYZ��o�D��%��$��j���Y�KxE��6 �rz�� ���<����Y�`����3�L��Q\�Zk* �C�z,p8��M|MPt�}z��F��d$cS�qǆ��w�M1�-��ar���Sx��N(��$��3I�D��N�(p�Aw'�
b�9�E J"dPɄK*��Ā�,jOJ�xAOC�9nj��^7`PDR�'{�rTfF�.@����,P9|�x*��:q��hA��<�q`�M���!U�D�A�i�S�Ӹs��}P��ӕsht"�6.�T"<-  �qB�o
�\���<CB%o�~RrCI�wB��Ei�V<�6NJ!7��OV=��F[��OM`B�T�`�nIHv΍�m Z-�$/�$f��4�厴/L�����2(2�Lc��$%9�^>�;Zq�1�������`�Zd]�13O���!t����� �)�rPh%�8��G���X؈q�4&�rzL� �O��."�&�oZ}&�ɦ��1f��d����U�p���$�<(�-��`�>i�����H��u.D�QQ�ߦiqh� Ad��_N��Y�N	5�l��'�v���OH��'�H��
���	 ��P�J+����I���4��u�xx�L�/~aȔPU!mS�}Q����)��I��mMI��8�E�֬BJJD���+W���D��]<z�(��T�io�>�&��s��Ԋ��_�,t���4aD�+��!9�R��z$�D�U�.S�� �'�Ո��O�h��թ�iU�oJ��$!��,L�Щ9P��X�+��	����$�O�!�ďV" �����?H�5�$�Q����h^�����S1k��a��ōR*�	6M�9�\�hlU�����uR�ǅ����I�T��p�sKUB�¡�SIE4"������:+�(�6�P�,��db�L@=辍��_�Q�E}(���ƚBʸL0P(��P#d �<9'$ː9�N!�"�&�	����E��)� ��D��L�f19+O�j��	+�Z����R �X�+�O�q����X����5;�h��Ɍg�њ�.�\�p6L�C�*�z�� �i���n�9����nM\�2�]�$:�:B䁏p%��s��r���e	5CX"�
S�'��~ֱ@Ůd3�(;�j�Jc/K�R�`�<I�+B�v�p<I��K4��$��L���.�w,�������q��GR�pܔ��$��$$
�E�/M�,���1�ڕB�K��o�i��B�y�p�Qì\+0���H�����O�6%���ֻ;Z����!}���h;Q���3$�DE��EyRL�a����`(��7,������8��L,���R`��{B���E��0���	A���#��̨O4�8��B�I��ĩ&f�"A�S�@�X�)ļ$�H�hiF
r�4�OX�(�iGv�$�zu	�#6����DJ�5	���a		�Lڀ=`W�L>�p?9��f���B��� UE�1�K�Sh�b��<}�bǕ.���#Eƻ���ܨYߪ�݇ĳ (1~��e0�
f������>���5Xa.}����pGp���	�:�pÕ��L�A�T��qDF��xqr��1\7��hF���8q�W<,m���KY7 �XE�.�8>�`kW��J� +Ȓ���o�9h٫'.Ć}�j��6d�_������:bBm�ã�(��=��2S�Q���҇�.��}{@�!��mJ��<1���t�y�!�N�����[M�'�R��BF]�P!5a�]��  %Ōm���	�:�D��a.ǈ0*m걂R�;����gB*Xfr�
G��F�'
���?��hQӄ��v7f!;T�B9B��A3O����U	.0���`*�4���[$�+��D$Z�: �ɷ^!~�(�0s���2�$�,�ryh����F���#Ӡ� �!�
 �2Eۣ�¯ue�xH_�(xR&C�}j(�XS1 ���� ڨO�ψ�]|��b,3�X�7�'�h3����8�d��h�<z��P��E,1,h���	C�����OI*�\ņ�	�olD1��n��/��	7bÎ8�㞄�i�-\E }a'��7�\|sQG]X�S�,��e:���qpʑKvm�=2
N�����WU��',A���#a�#[ �=r�fƒ�DSԃ�RF�8��>�������Mۤi�7j�.���5[\H%���M�'��Y��óH�x�E�Up�TM�-��4�MI�"���	�������-ʒ�TdX���<�dgI�Ť1,�~Aɥ�Yj%$��/"��A�vK,	�pk��I�BTJI�lטT7~u��΄o߆�Z�hJ�3�,�H	�Ӫ��bAT�[?:����9Ô͒�*��	ype�(,�9)���y�Յ�8%���O�8�]�|ٷZ�?����-ЕfY�AgF)w�0%(���@��v���$ۢ ���*�� n`k�� �0:a�,]H�p�5��lb Fay"I�+s\dʓS�,�pՍ�/̒O�4�C��b2FTZ�◣P��af$\1<�Hc"kT��~8aF&!F���D���uGC]�og�LS���84�<h���jRԤ�r��E�l�A��ѣ�
���R�� ��>wa�H�Xv�AS��i���H��tϤy�'+��; �̥�|J'�d�St�ݾv[.��i�C����ɶ~�d؂���(I�>�n�������i�W+�>q��	WF1�D+}b�V;��i�����:�R�+c)��Z�Z3�LO<YX��ˣ�	0�� S�B*c5��(b�~:��%kD�K�F2���qTÃj�qjyRqj?
V*�h���0H�p�OD$��9w����B-Pwi����@T *hn�1��iT�r�.��D%���(O�8�!%Qa��wC��P]���[���!9���k4ŵ�p<��ę8l&X�+�_t
ԺbfN6}Ϝ��fa��d����$�?o$H��j?6�P�cf�3}A����Tj�x�gDN�߽�t��n��� #��3���1�/XQ���:G�K?x��p��.�x �v+�b�L@�g%�7*���FxBMɞ�,���F$LE�����Z�/Ԅ̹��/`@��KU�bC:]�j�.�bˉ"�A�#��9��m��xE�u�&Ŕ���V$zXb0�R� nLa���![�Vm ���B[(4
f��4&�N�af�&�zY`4�	�*sʰ:�i�>)�b�x��D3Hq�6��S��6%���Jղ5�'���xt I�1er1p�G�S�+nݎ~�Je]���S	�dv&�"��,�|�����,6
�Abo"lO|x��N�=�+&c��VO�Y��ie�=��I�(�=�d�g�<(�D�k-��0�Z5q����㎐H��W��b�5X�i�*b�ț!F�=a2�Y�<`p�A2ʭh���b�����&gА��~L4BH�,/J���	�VԒp��T3��E���D�)���jA%W����wqNX��	(Zh�
��J�`F��'��Y[�$�%�Ba���3G�:�+�A��ո'ΔΧg��,�Pm�8�+O�L0�\�r���qj�4]�H���'3��XC���&T��@x���#�NX�(��ڛj���}��%D��"��KÓ@��K�I�h�@Aʷ�79�H)Gx"�
	%�8����>$Qt���g�_�	�bp���c��^ԁ��U��!��ю�la3�ѿ&�~@��L�J��z��C��i��)ε���s���G�M1oKQ�9���X�(%!�;��aنd�#��h���#z�
�1D��-�v`:6��v�9��1����aɹդ$2��M�z]:S� �Oi��¹r�����,�k�qZ�Ǌ�^�iW}�RQj����p?s�ȓLs���BQ���� �e�'��a� ��g�qy�C��P����RtZ���l���FO�:}Ƥ�u"OJ���V�3kP)�f�r�8�+ӭT�0j�:��",��#Ӄ�ܟ"~�I)+J�P��K#Ҡmv���[L|C䉊H�s���u~�	����"X�dC�
"�������B��%ʈ��FC�I�D�D̛��)xH��0��%��B䉅
;�:�O�H:5��*��G�B�?.��]s�g�)���7'AZ�B�	&P[<<a@W6I��j� nH@C��2Jb���5��o 6��6b[�J�~B�\3�8��c3d�b4��%K�C�I�3�4��gD�.ve^��c)^7��B�I�S����܋q�� '�@��C�	����͹eD��+4����C��:.ވ9p���
=B��!��sM&B�n"�`
Qg)�i�Dn��3`C�	�S��C0�߳;�)A�i@8|\HC�:	2 ��)N,/B�\;R&@ ~�B�Ɋm�l!*�Ep�l���ߛG��B��+&��i+"�O�e���p�eµ>TC�ɍxR@N��DZ0��g�E2$��C�>y��8q�)_!H�� 8#�бiPB�	9)�
 U�۞:��$!� K>B�	3&���+t��F�I[�
�9.@C�=|>E���0}�~�:ƀ܎[�C�IE���V�P�I�d�S'ٌ=>B�I1x�r�S�Nٹ"�	(q�ԝnm,B�	-j���U�^�rՃ2�֑M84C�	�GF4�;�([b�Xu�`)��+�C�)� �m3s)_N��iCb��(�p�*�"O~A�h�$g5��6�4_�X�"O�#s��~�� р��r�"O��
%� �6���RuBT�0 �*O\�P��	V6-#� 66�����'~��q�P�s���H!U�}3�'g�,kǆ�-Ӛ���
�ú��
�'SQ��O%:��$r�#я��	�'�J	��C<��L[!FG�}oZ0b�'�h%;uL��bӮɘ��5��u��'���`7#�1k���а�A{MnЛ�'�ΐ�d�;oA���0�^$i1��P�'���c�� @���Rd�(k��\�	�'�H3��`(�� ��ַ8I�	�'QbHhS
��9\I���M-WN���'`|eyD矺*�ih��Qt4�C
�'��l�Dh��#��1;q��i�	�'��H	��S䌕P@�ٚ&d�	�'zԙ�&ʟ1y򼅱�$��$�x
�'�(� E�h�� Ån�Zu�	�'� �
�=[�Չ�e�vI��'�l�Ӕ�:S0�YD��?d�Es�'V�ܣ�E�,$Z����[���'�BF�|C6��Yb~!�'�xA�7��6O��$��	 ��
�'Bd)#�v6��󢐯r{Dp��'_�	'_L�
��6#�=p|6i��'��1Â�#0trLjU�� l�	�'������&N��%�֘`��MP	�'U�m;U�H�O= 
u+�Vn��'�-�с��F ���'��b�`1�'H &E�%��HD��C�Q��'�V�cF�Y�^�PCφ+�T���'���$*��Y��`!���<2��'��csN۵#^�����|��'�d	��כ	�����CRt9 �'��ue �G�-c듇q|4��'M�-:T˃	j��� b��X��'��I�cٓl�4`��E�P ��'[�����*0B��j`(��7�<��'���0�/H�K�j�%�X=-�l3�'R\�ROm5drh�!��m��'�<�pB��+s`�a$D�E�(�'�<E �I&���#I]^�H�'/r|clЅGb�s#�C/Q᪤��'��e;!��I��;@�q	P�A�'!��ϕ>Hdx(�(�qi4z
�' ��[Dd�2Of�ɧ�W;g��j�'�~1�woB,m�t)�ׯ��!��'��AC6N��t�)~��y9�'�lA�f�5z��EVu��'m6D�5AL�DR���%CߛhV���'�1UC�zb ��/S2]iJŸ
�'���p���� P�G
�!T��-X
�'�Ru�MUV��Йr�EO�a�	�'���@ިS���a��k��c	�'� ����j�w���[N��h"D� ���ğO�̰�b�/HN�X&!D�`P0�� _��@�2 ��с"+D�X�f�	!;�8,�-��0��p�)D�P�F����p��s
,* ��g�-D����S�%�D=�/U�:\�(�'�+D�(���ʆE���Hv�c�z��gG,D����+�{T ��a�Ef~`ю4D�� <��թ;j��ȠA�_ڲ�g"O�1��G�~�L$б���tX"�"O<XH��C�Q��c�hW�f�i"O2��q��J9tak "ưJ����"O���ծT/����6�G�T9nT��"Ox5�D���E1�PK �q2�5ʴ"O|���U"$3���'����"Ov,�j�G<^��G]
^6�\�g"O�9�2MjsH,��b"L�(P"OPLqg��7�U�� pz�g"O2��TǑܥ�U)�t�ѥi���y�&��/NN���:#:a�R*�y�PJժ���Ϙ�)���Q%֕�y2hB� �pq2W�	W7�8�!����yRB
(�@�6���7�����X��y�nÒ|�p��#yKr�Ib���y��̌�T���ޡl��t�@D��y�!]Q`8�@.(NF��¦+%�y�X5IU�|�1�3A�6�xՉ�(�y�͘��I��B��P?ܼ2�-�y�Q-I�B���bM�y�M����3�y����?1�}S�Ŝ�[.���X��y�%_]!����p!`��C$X�K�'���s�Z'7����E�	�Lq�
�'�,8�"ռr��U���P
"��	�'h�D[���qipD`3�S�{qTH*�'o|0�1����{eZ�@:����'��4�c�+�,��N �3b�x��'�J�!�FT|����)Y�P�'�<��kK�W�d	��RT��[�'o�����;-�B�b���;M�ui�'��� �#N�8�%�U�r����'���ʦ[�9�*�<�|�!�'�l�bA-�G���5 ��/�@�
�'��͹��A.q�ք�yU���	�'�q�g-,,kj]s6�\
���'�^�B�L�n�nD�E���� U��'�֥pW��}�6Y[Њ݈�>� �'s�U{�l�az�d�K�]*�'��T��gJ�a�b�O<<)��:�'����I϶^��q��MP3��u��y"�)�!)G -
u�&�:Ļ%�9g�pC�ɹs{�9ڔ�tS(�x$�	P�,C�	>��Aj��R#9ZH�s��.cC�ZҌ�F8-�4# /�*k��B�I f�1h��T�W�^Չ&�o}�B�I3y@d��Kƾ+�*��DŃ_@�B�	�u�lpwd�7�ZdYs�A��B�ɘ3�~a�0�"2�CAD�3i�BB�Ƀ4^�x�+ďdx�m�T��r�C�	�u��@k'����a����B�I�&�X���̌�����gF4lnB䉱;F&%h�Kϲe<u(��a>RB䉙u9� c2� *!�� 1E�'mg�B�ɹ\��!sh%r�1ڀ��<��<��K�0E��&̘T��B�e�>y�%�ȓv'�@��^��Į��jx�ȓ-&�h���-d����ň1��5����@�@P^��MrՇ�;&:ɇȓc f������)6� ��E�s@`��ȓ���j����i֨�1ƤD3L�j���4�^,�F�p)�h�q��ACr؄�h�����89XH�	a"���݇�L���"�A�e� qaQ)�<#�&��S�? z�"��N��rj�`�6ذ6"O��0�Cj��p�k�0R)�@��"O�����d`V�QA�N�*��s"O����ъ�.9�2�˽h��c�'�ў@�gk�.��U;��܏^����aJ,D�쐗	��zfld��ď8�t�{E�(D��8�GTf�]2b�	qL�3SA(D�\:�"�(\���Z&�rp(D�Лw�L$8 �v�C|���`�$D���ଋ'9�,��,�S���Ԧ>D��sF�&/�t��C(՟6���ңM8D�4 sJ�>s�d��dF�zA�e��*;D���4�Z5e�	���*�ҭ���7D��zb"�)�AiBqz�聣(D��"bR�;��s�˚R��"��!�O��Opt
�9E�(=���ۢv�T"O�P�@6z��%��̂"z���"O ��8/�Ό3�蟤D�^8"B"Of�زh[�t�x�bgҜ	��"OR��c&��q���k�A�"]�H�c"OJ��P�ض
�93����|.�%��"O(� p�R	b~��с���x�Z��'���ΣU��prpC��17.� B�!�$Q�X�2�0��C?bi�F�`�!��C"s�4}�d/�!T��8�d:n�!���h�7��W�ڸ�3�HFO�C��&Px=�b��1��L�R'ƇHGzC�	A�ā)��9 ���� #��C�I贡SE�r^@�AB-el�C�I2�z�yw��
P&���U�g�vC�I�m\��Pǌ�Y�
�)�&G*#�C�	�g'j��C=O�YH���]R����>�L��X�WN�!N���؄�֚N�!��9�E���f�!�&#Ї@�!��D
#sr�j�'�/6���(�<.H!�$��4�^��3�@l�h���ľE�O<���ܨ&�(1���}��};�ǔ!���	�B$�D��\�$�&�?:!���W���"$b(M�`ņ�v!�$̌]y,P�K�eQ��c�f-�!�DְT.x�т��ICJp�&6�!�J�%(�Q᜾��0)����C�!�.�����ƽv�^,0�A!_�!�dR�R�&	�K�&��𕬟�T!�̹�$9#Fb�tx�Y#C!�䆉�Fݢ1g�_h�����Ӭ�!���$�1�8zKv�J����W�!򄋹	Lf:`攇u�^��Y��!�D2 'Lmj¥\�HѦ]���ň7�!��U5�@T1P���f!x��֢�!�D߾H �)�X !�Pi(l��!�$�/M>:��A&�*���Õ��Br!�$y� ���	�=y�����`T!�D\ mX ��Ιqu\�g��%!�Č���@���܄:��6�W �!�$Y/_5���ͦ/s ͛4ოa�!��Ƨ(� �cb�&h]ĉyV�Ѫ7�!��
�5��!��a��ID�t���@�!�D\	Z[҉�m�:/7�ūׁ� R�!�$�����
�'4yBgB�4�!�$`S�p�C���ivQ`� ����Ty4�r�a��3ʢ� ��yB)c�d �f�S!W{z���f� �y"*Y�	��r��@�D��&�N��y
� �����<<C�]��'��"���cA"O���mڛw��D�GŃ��(�D"O L�d��%-��A,Z-u�P�;t"O�[!�ƹ��U� ؎T���A�"O����O�JFK�]�)����"O�!�8	��%{��6�:��q"Of��2V��ț�Y|bH Q"O �ZW*�QiT5��� a��ґ"O.�0ס,n���*w윉P�d�k�"O�9�R#^|P�C��6$�j�"OPJ��XW�.��S���5���"Oz%���آx��5����p�"OL�r��9�D�k���M�L��"O�D��C�d��h�!�(`n���"OF!�D�X���k�A��%���"Obp�w�Uj��ц�.9��"O ��Q���13*���O[�8��]Jt"O��D&�9c����M�����"Of,����h� ��8.� 5��"O�	K�DO(t�@�+�:Q�I�"O yz���,�r��3��I��"O�((�������RA^<�8��"O@%8@�U@�X��`��M�<u8"OH��ժE;Y����n�5G�EiC"O$ XG뗋UVԩ����Tx��"O�� ��N�L�	����[�9��"O�Y�Qj��/�X�p*�8y<x��"OĀ:g��9�4���_� ����0"OV���Ʒ^y��'
�~��	�"O"����Y�F|�v��5�0d"A"O���s��?hΥ��*�DԺ% `"Oh�qEhR�0Y�SK� ��B2"O�ᒶ,J�&���J��Or�)C4"OT(�׭�P[��0ǌ�UF��T"O� �1#Q��D��!XL�;�"O@�mO*gq�yG�J�%�5A�"O�`���	�Н��� �B�d�"O�h[p�QCdx���$Y��U"O�uI�ķE�P��^*<Fna��"O����ԛ�pzb
2#���"O<d;PMЛTc�C�f�!�E1&"O�P�u���<�D|Еf	 $��"O6��$��g�����JN���"O𤉂DW�&)�p��Z�>x`r�"O�Y8��[�+zQ:�mA�xp�"O���H݇Y[�D�G���*�"Oa3T@��c`,�ٱ�5^�a�"O��@p�2͒y�'h��5��"O���v�L0%tq�0��D�B�"O�|	�퀜o��p��Ȇ.�q�"OD���Fq:�DY��h�b"O�rt�UE�x@�D<'��	P�"O���&	�q�`����T��"O����aI�#��"$W�Y����"Oz�s U�E��uJ��9h�\��5"O �
D	����@0��M9�j`"O�\Xd�Ψ+�.�c ��w�^U@T"O�aj�aԭE#��۲+�`]����"OV�8��'��)��Å ����C,D��2GM�#� 䉃�Ƶe�8@�n$D��[���j�<�&�*s>ܰ�"?D�pZb�ZkF�U ��K�6�*ܱ�-!D�Tz#�:W}�d�5	��PH!2D�p��cC;J_�\"%@.S:�C�1D�� 
)X�͓y�*D7a�*z��I��"O,��d�б	F��07��*'zr�x�"OB���Y%!>^��ń=!�Zq�"O�=��(M?~�p[�憎T �M�"OLL�@��g�=��·33���� "OtiY`�ڬ<(�b�"Dv�p�"O����D��G�
w���"O4���O<��bV��Pt�x!A"O��c3!�7 ������jm���"O Ś���{Î�!@�&ʶX �"Ot�=fg�
@�ޏ$� �:�"O��aԧ͇`O���A*eQN��"O6I�u	7�%��bÌd����"O�t	���8"u0,vh\7!�Z��"O��g�X���!'�w� �C�"O���c��*	^z���䎳6n&�rc"O�I(���P-�mcǰZO ��"O��i@=u�ӲDM6��P��"O중)�E�� Zd�
3v�8�X�"O�)E��4�ؼ���:b���%"O�d��l�&Ü��qA�X����"O��@��]nF��@ҔK�]*�"O�T�Q�<
@ܵKTϙz�6�x�"O��򆂟K�^L3/CP�.ī�"O��:�$P/ `�%ƅ}'����"O���%l��_t X!''�%qP"O@<�F��5%��	�囼S��@"O ����	��U��$ϚX����"O �a�3��-���;mJ v"O��d@1w�l�Ge�)t��{e"O���Fc�=���%*[�9Z�s�"O�Uѱ �U���A�>)|[D"Oh��-� ��HC��!�9He"Oh�	Q�B���{"D�8#n����"O����T3)+��HP��5�Pّ�"Of$Q� �QU�dk����!�f"O���k� T���8���;{���d"O��Q��A/?��3�
فS�r��"O�i3f�)]h��Щ��i4=AT"O>�h.�
5��S��|1�l�6"O"�Z6��>6 j�(�胢
~��"O��S( bH��E\;	`S"O�a��f��S�H㑆ˉ�\�r�"OHej�^�%�TA2��iB�"On�03O��D�|���7��T�"O��q���� ���O�J�¤)#"O�8�UO�!j�\��n?-�D��"O�qX`Xk���@oȜc����"O^��q�߷{U�����:.\���"O6!�@��!n��aH��_���A�"OrE�ehD<�6���#�"O(g�ߌF�H�so�t��1"Oj��%n����xP�1&���B$"Op1���=:̜��.��l�D�j�"OpHimƟ_qƕ��dd�$� "O�)e���m����`-D�#P�L�$"O�PSү�1���NS6��YU"O�E�1o�Y� �@@M�#z��r"O�ո�)^�|)4l��.ɤU����"O��ȶe��q:Vh�� (����s"OV)͋? �A!✏?��ɂ�"O�����;�,�a�D�<8w"O���0��\����� ��V,��"O�q��×�B뗏��8!�"O� �!ӢF>0k~u�eH�l�(��"O|��bb��>�=�e(Y��ƙ�p"O�+�mS�Lc�I
e[�;�4�z�"O� ����"}�<��}Y�)s�"O��FK�81d���ăb��|)`"O�h�QA ~����Æ.��t)�"OL�!�Ǭ]"Lѥ��n9&��"O>)"1́�z�P@Ǘ*[,��"O��b��R&X�`��d�d��"O�i`��&Ѽ� #L:9���"O@���B�Q��� �H�0S�*�hd"O�m��bT=;��JV�V����s"OB�{`�T�O���n����"�"O�Yq֧C5$h��3�E�jU����"OF�0
�&?T(���^�"���"O�i0�`ɞ>ĕ�q�K�x�l�b"O��q�G��'��`�"ٻW���"OEb�(�2%��H��ǩS�,��f"O�̠H�f�*���c�@��6"O� J�?t�X-H@P�G�&L`�"O���/�0�T���m�hMA6"O�-���?L�	��O���T5�"O�!qh�jx�� `
#��8G"OV��̲4$ŋ�O͒]P�@�"O^����U��5a��_;p�k�"O��� O	�7>� ���1I(�;"O�A��E��ktD���$��$�i7"O�K�W']��p'?��-x2"Of-�퀃_�Ɛ�����H{. ""O�-� �$=h�<���K_J�Z�"OX�X��@K�l)�dG�,S>��E"OF�i1IC0� �Z�!g�� ���P>�A�)���P+��Q�p�x��2D������b��xM��qU��zd-�$4�Oʼ����YJ���� �S"O�E�1� �⌳�A\*
���K�"O�H�P��U*� �|��Lr�"O
̛­K�\�r�)�*	~Z\B"O쭹F�G�}C�8 �D9?pd!3��D�O����Y�t,��#�"aTy��&Q2- ��W�q �����:�PH��.^<CC(B�I0+�4*����)��e2�� �:�"B�ɡn�l@����F\�ē,�b�B��&^�<�I.�b�2��։�h�B�ɤK[���r�]^��:Dڢ
� B��,�<t��*�6P��7�6c��C�I�{Ѳ$�І�4K���xP�H��R���y���K�D����	~�p�����yr��,lH�K4�UTu�h����y"K�xД)J5ߤI��MSƮS%�y�LB��<%"�P�s�L+��_)�y��$;J�����Eh���D���yr#�\� �\%��%��:�yb�_y��3de	0VѢ��B Ց�y�Ĩ/����*$<=
n�yR�J6	���T�Gs�X���y�g�+�
)��
�9A�4������y�H�?�dx��i5` eR�Oޕ�y����4�NZ��B�8@���y�kC&"黶�����p��n���y�懮y TA�lֲ�b�
�d��yb�ǓL���c��6�p�����?9�'a�DS�@�-t���!�I#���	�'&��Q� ��8�%��~]�u	��� ̩
���f���-W���z"O�L���B��j�;'�I�7V���"O����X�V����E\�|d��"O�D���<S�� gBT�r�JH��ON��D^0Ȩ�秕�\�����8D�D�����R��� !j�Sp�x+��7D��f�P�J�R�j��}vjl)�*O����j�%�,����#d@�|#�"O8Ȫ��п>*l$����$X���"O��f�LZ���gB4��"O8�`b��|T���ۏ�!"O�̀T��/G��P'�?4�T�ٵ"O@��*F��$@H1 �.$("O:CT�ΰD��G�����"O茺5ȏ���(!h�2-D���"Odahǡ��|`����ܫI����"O�A���wFZy!�e�.���"Oj 2�háby<�C!E�"6�;w�'����@�x�Ś=\:Tp9�B�6.�!��J8&0��g��5�J��Q��W!�d<=�y@�F1S%ĝ��gǲMj!���ay6L�pǎCl�{���\!������d�=a>nhh�kɄy�!���$�R�1f�K��(��'�G�Pz!��n Q"b�ó|���$$q�u��l� ���XpJ7�^.~�\ؓ��/D��D%�5W�Ĩ�v���Z�<�c1D���p���Y-!�b\�=D�K��<D����߹1Cl��#�Z�*Ш&D���bd\�0�����x0PN&D��BD"��Pf�@�
�W���2�%D����ё;P�y�Qg�+ԺPS�"���O���Dο3�,�juc��$D��Ĉ{�!��-���Dg�,9���+BؐK�!�d�cN(� I�.����eD'�!�% �p�� �psb���*z�!�D#a6��Ӣ�a�6��R��?�!�$�1Qb=�0Er�\}xu�P�'!��ۋTϺ��1�ߩ2��k� T�{!�	�]Y&�(㩘��0�`U"^!�K5
U�%�Ĭv�8,B�O4�!�6`wj�[���s��q��d�*@!�["A�Ű@��"���+$U'!�D/f[�xr^"[p���!�}n!���Q([�G']0ȣ��
� �!���7�,�	���}��%y�Y=!L!�����E��+k2��AH�g�!�D�7<0�Uam>�H6��(8�!��ՔE��<AS�Y�b������Ĥ+!!��9|���ڱc�!j�R�[���8�!��r�vi�����k�	�=%)!��0�n ��,C�m� ;(��yB*6ָ��MI6f��Ps'f�bO�UnR�h}��
�b��s%:�	]��tp3b����*�$Q�q�*D��p��Z���rǃωk�]h1b;D�����Y�b|�D���Km����8D��(w���E��1�&�KJ�ƌ(�<D�Т�՜n���
u&
���8�5�,D��a�	�kվ5���F+"��f��</O����x�(��h�͐"�N70!�$�.�:q
 �J衑�	!e�!�$��I�u�㒼V&r�BL+r�!��əbs��1��D�%:\@��M;+�!�� ���CЉR�XUhcm�7(h�ô"O�i�Q@�Y�θ����c3�1"O��	�$9J�,��Q�0�Ot|��E��Q��?
�x�0(3D�Ȑ�ɋ)V���򨐞���#�>D���#G�	�N��d�ΡB�<{t�=D����@��:UX�͇������<D�Pi�![_�҉õbY�P���cej;D��q�`��q8�@%�UP�ԣ�':D���
�M��[�MҴhT\q��2D�p��'�:�rpӷc R6�9�/D�X���38�tɱQ)�� ��+D�����E�L�#5>	�1iW 5D�X*��y�0Dp���uˈ���0D��p-�"]M��%e`��/D���#��kdc�&C& I�1D���mD�~��a' �&�
x�&�/D����"$Ȓ�a%b�\��l#F)D��{�g�.32Aۂ�
�ъ|�E%D�xP6˝�s����� T�gR��)D�iA�Y$Y��]�a�Q@e(�;�-&D�X�V��#ਠ7��}��p�$D�D`�Db6E*/J&�>ؠ��%D��b��,e���!e�1�D���(D�5
���q#�D2
mq�	+D�|��ÿ#����@����e(D��y��&_��a�h%k����&D�Рb�N�So:Uy�Hڬ"g����"D����FU�.����r���
Q>D�π>D�%�G��T���(D����&ށ^��Q���X�(�j$���<	����-c�֭rA�ZLCX)#�#�	w�\B�ɩ[�:8�dΓ�|�IX�aO�Z,B�	�`0>�#v�Hn��9�@NӐY�B�=4.Q:��Q
&	��I�"ռSϖC�	�+."ų��O�;VJ`�����/#�C䉮0 `�Y	qy����
�crC�IT�t��mC71ք�"��Gq�nC�	!�|�g��:h X��1OJ�C�Ɏ?j$��h��R"H0�b�)S�pC�Isx�	HAk3�@��q���O)Z�O��=�}bQe�3r�$ ɔ���j\bFmPQ�<��C�u缹Z�������ѩ�M�<����;��틃g��KQ�=�1��n�<Q��- "L�g�×8q��[��Lu�'�ax�Z�;%��@"�ճ= �A�.;�y����?[6��%ŕH�BJ��X;�y��<����e�&A�`ۃA����d�<I������]��"��OT�ܡ��J�I�xC�I�t^䝈㦌<v� 9ףG
�*B�I�c�d�����ߔH��F�D��C�I�?Δ��	�O�(���
o�C�	a��bBň� ��d�� �IV�C�ɑvb-ZqGӰW8h���׀��C�>ʖ��ۂ_h Q�D�V2�˓���hO�错j<�	���(�"��7+�!��c)���+��ZxxiX�)£�!�$�r�8����){vt��-��!�dB�l�D,� �F�YFt�!d�$�!�D�)7�"=��5N'R�f��l�!���\��Eߔ94��� F�!���g��)�Y%^�fL� �Z�6�!�DǕz60d�7@�P�r�*m�8G�!�$� =��k�˙���q�ݬ!�� ��[HP�#	|��k�.g������'��	%.V�aފ1�|:�h�Q, C��9�&Dc��+/�DA' N*&��B�ɌC�n��k3pz����9"��B�	�1�He��Lë9��u��Ƈuyr�D�O�����W�
��(?��e�p�ʨ!���U���h6��,�8@T		!�
=��q�lDY�h�Y!�'��}R�'��I�N8"�_�!��B�Y�O4�D-LO�%k���r��I��f�cT��b'"O�a���H�
ǬeH�c� Wf���"Ol�qd�֨X��<ؗ�Լ~GzH�Þ|�'n�9�Y#@�!״$TH�y�'>��`�@�&p��rsϗ=,d,j�'ɾ���֤�v9��e�%m�����y�i��Dt�8[&�ޟ3�.�r������0>i���;#$Ղ6����zP����|�<���E�F[�����N�5�d)�Q(wh<��D��D��iA#d;��Ф�#�y�h�&Z��Ӆ�Y�b������y���h2� s�Vnj���`���y��	`1bT��	O���G����>��OZL��H7 ���I=s^�k"O0u�H�=C3���3	�duVT92"O���/D��9���Ƈ_X��"O�ᒋ�(\e����B�|\�����'�!�=c�A�RNr|�*���1!����iM�?Vav�j�h	�p�!��
��ܜӢ�W�aG�5f�_$�џ�F�T � 8��"�(��ը�y2��#WL���͍�J�iq��"�y���D�hW�_Z4�!����yr��lV� ��6:�����^��y�ʄ�{#:ш�`
�8�*�`v�C�y�,T�^�����ԋ{�E��A�#�yB튛l����7�.p�.�q� -�?q��d3�'}��Ye�WP��*��K�ٔ����b�F�8z�1�C?r�.]��o��Ö��{��T����G�(��ȓ0(�]�ѩ�s���%-��=�� ����d��]Zf�:2��ͅȓg�l���<7���PN�!d	Tȅ�0�&����ӠY�ր��)��AB>�ʉ�D=�t9L$� ξ&n]8ƆE�+���ȓ\�$)�B�?�80�瑺eV�х�96��bD�b>�Y;��E�hidp��`S����/ �����"8-�q�ȓR?�8$Ŏ�i�.�:@@Q7*m5����i���ЇhH��+1�5V7�,�ƓGIFT�t^�b!R�F�Nƶq�'Mܠ�vh��QAf�( �������'&�<��n���AkVG1=1�iC�'M�u���͘B¨�h�O]�9N �
�'N؉��3�(�� 6��i
�'^��J��Īq����S	ɐ'��"O��b���
����@ =�q"O@�����2F`ѲF.C9xא�s"O��XE���]��((�0� Qj�"O`� ���\i`�sPW�3��(�"O01:^g�̥��*æc�^�T"O^����ϧo@�%���@�X�B�"O�T`T�J�Ϻ9��+���yB"O�<0Ԇ��d�'e�BC����"O�y�mY28����+.�@�U"O� ¡q� ��wmH���SS���"O���+T��݂t4h�31�'����,w��SP�H4\��!y5!�KrlSrg� 7�$Q�BGW1^5!�䓤J�h��Z,߼����+2!򤃝�P��D�$�@Bg���++!�ۧ\�8��a!�s?&�H�FP�_5ў��Mp6 ��T+&$jH����T�C�	��~� ���Yb�jgJ�~<hC��!4肈1��>V#�;�S�G�C䉟	�$e�SD�6r6�4���[�F��B�8X:F2�`Fh	��@T��,<B��n���B�#Z��a���)��C�ɮ2Yl��r�|�d�C"L��lƣ=	���}��"Aԥ%������aR��J��O2�O�$0�'�y�%Y�j�ldAF	�C@Ub�GK�yRÎ� �F�!V�V�	7 H��. ��yb�	&i�ʵQ���~���$���y�l�*��J�L�zw�z¨��yJޙA����U� e����g��y"���o�~8�w� X�(����?����ӷ��)�#-�t�ʵ"�M �YebuE{�Oʐh� �
;�u�dj]t[���'�x0R��SK��2G[h�ؑ��'2���nG:0Hd!��E ��'��� Qn�'S֮a��%P�	.Z1��'�����L-B�2�A���m�	a�'�S�)9A�)yp���r�I�'r�QR��D�%2���c x�|��'����A8����l��\�Y�' ��
����偓��8�'m� ��7rs��r4cW�+��
�'��( ��n�X\`c �~b�܊	�'�␚�_�fb���P�Ir6@��'�
h`��
+��5{G�UyS��OhqzUiձ0�S�|�9��9�?��'A�A��o�r�AV��R 5H�'�L��aY���P�de2D��'�l��5bK�N��Z3��T�@�R	�'�Z���&>� 0�Y�L�H���'�
�G��
y�cP�L�p{�'P~��� x�"d�עA�H�ąY�'� QJ5�4`�` �	�E¬A9�'�n�ʂM,a8P��҃G�x�
�'o>��.V���n�S� A�`�P�<�B��u�<�eLճY&��"��E�<!��Z �nP��@�;�q����W�<1t/E<@ �d�B%�-g����T�<�ÂRX�L!+�J�' @ �ؑ*�S�<5bG��t�	�-;��ȳn�z�<qUN��蹀I�4�aIx�<�S���/�\`Q@�g��m2�M�s�<���uTZ��W��=0uH��S�Z�<Qvc�91�����bB�0�ȅB���S�<9���T�5O��Xn���c�f�<I�F
�l�� Z�NY�<Jb�<�VfE8n
T�'��h	���[�<��V�#e��R���4���Ã)�l�<)�JX�.��k����A�<)b	G(2nf�(��Z<q��H�L�y�<�ԓ<��u�a��Mn�(�y�<Q��)Z��P��F�A 8@��|�<�R4F�X���V֭�D��u�<���!qp�,C�xM�fIՏA�!�� �)��R�;B�1*�I� �R�H�"O��S*�,����
�S����"Oĉ��Eofh�i�)Ɛgv2�Yr"OZ\{��:j�l�H�I�@R0��"O�e{t`�&?�`��jC�>+��@"OЙ��'V�a�0ag/�x'*#�"O\���U���.�k"��+1"O�쉠��
&��UKn��}d�y�"OZ�U.O0<�ҙ9B'[��I*�"O�DY÷� p�_�*�p���"O���Ɖ��i#Z�T(qݖ��"OBՀ�.J���g*,��uQr"O.�#��C��6����Z��q�"O�=��g�/PHy�	�B����'�BŇ>$<��u�Y�i�.a��)V^s�OB�=ͧ�y"�ZQ�����8�dd0W㜢�yRV��0	;�ޟlw���S��y2H.���RS���nu�@����yr�^{�hB�fԷm\B�b`�ћ��x�� �aox�&Ɗ�0�(�r�
�up�	L����Ȓ�Y���"F�,��"�j6D�L #Kҷp˜0�H�6YA�8ՠ�Or��hOq�N 0�ѯ~" ��gk��i�
t��"O�ɚ�%T4U�
ᘒ��6첸��"O��A4�P'� 1���h}܉`�"O�%� ㉺QTL���$}EaV"OfdP#D��+eh{��Ln����'&ў"~Bf��~k�`MӖ����@+�y�M�~r�T��#�!-S��`��yrlL�}�FM�T��U*2P�v���yB�P4[~����Mƨs�C3�yB��Q��a'b�W��$B�Ǳ�y�͛��<�CnՕ[X��V�F4�y���.<YG��PX� V ��y���z<BD��[3������y"�.c����RA�XxʱmC��?!.O��Of#>��"�(-s���leF����WJ�<����+K/�H�p�N�j	�`�G�<��G�c�Pusg��g�1U#�A�<���Y���� �)P�QA�`�C�<q6�[�v4��D߉ F����B�<��L��*�X�xh)�o���$b�p8r��1�X���#��$�<����� 0el��E%�7�	Q��� c��Iv�8� L�&�m
Z����"O�Ё&e,�ɰ^�R�UJW"O:�`8t�� c��R�%�`��0"O(k +Ļ2�lԩ¢�<���H���Z�i���6��b� M���*D� (ë��N�����|��(0-ړ�0|�v&,p�Li��J0>��,�K�l��LΓeєlH�'>n�B�b"�ӟu�ࡆȓGa�Dp�i�"����D��4 ��2���W�2 *H�h�l`��C�Թc� �s~Z�	<}5����j,��j�蝶]�Z�'�aTN�ȓN D#7.\	�f!�����֑�ȓ,� M(�.H
y��-�r�J4dtF<�ȓZ��!Ȁf��`��9����3'����'|a~�R,F��0bݳj���xf�P��yro��m�,����bm�H˰M ��y�n�-#�Fq�v������&�3�y҂V'kh���"M.53���y��Bi�$�c�}&u{޴sh!�� ��t�JR�uJTO@-�]�"O�e� �+R��axv�ڏ�����"O�|@N�E���_�X�T�X�"O�Eڲ���B�Kg�
,/�A "OL�2&�З]&��i_�
M�"O��Q���*h**���(�&�:�"O�٩�Z��Ľ��� P�ID"O���Ô�@/N���G� 2Y�pB&"O�P 5*^�GL���& #G<`
"OzX��h)ܖ�����?�ܩ�"OF���B��KIƅ��Υ_��%"O:���mN���aqjP�tir�Q"Oz��%n@�>``�{��c�S�"O�A�+E#D�D�G�(;U����"O�H���Y�~bbL�#�����9"O�D��B�m���%E����ћ�"Oy��%h����C��r�b|��"O@�8$j�!�� �"S2���hC"O�T` �!zp@��A5�D��R"O�5rbg�%8����'�E12��"O�x6J�;z�y˰8r�0�"O��L�&�Xd��lAgn|�چ"OvM*!�6&?&$��J>'Z�Hd"O<�bW�2�0PJ'Iռ'�0Y	�"OD����f~���AFQNuB "O�Y�m˲��=�7`׎�թ�"OpdB�\�8F�<z��۔,j(�"O�� ���N]Tغ���"�8"O��y���5{\��㓒M�$ӓ"OZ���տ�0���$�(��q�"O�����Q$x�*�IRc�W��e�E"O�,
�ʈ�I��h;�a�=C�U
�"O�E���D�X��e84�/Ta�c"O�a�	De���� l�(e�m��"O�$q��V�0�cK@%L�\�+W"O���+yI��ɷ�^��ŨE�y��TF{6!x"P����A�MF��yr��3D��dk��>$� Zr�^!�yҪ\3�0)���5u�i ����y�o	�܌ �C�qk�Ӕb�?�y2�B>X�b�xEɊ�f��e9D�7�y"+�U
T�+��G(p�vY��)T(�y���j��Bu�W
Z d	��J�yb���v�\X���	X���,�$�yb��'-e��m�ZѴ�Z�ٙ�yr'גA{^��ȣ?�X�Y����y"�v����$�ހ��)���ٚ�y���x���#Áܝ���U�yR�A�a��)�w�
!V� �c�%�y���6O먭K����e��$�y�P�,��%��֣5� "�٨�y��A�|��:��N�	�D̹�섑�yb������W���*��Q��y���M�,!�ʃ~y
U��y�J_/X��B�%�"y�L��y2b�/�0-�ၑ �đt�\��y2�<���z��jܜ̳ Ɓ)�y�؉YrXX�%ꚝ`q�gͅ��yB'F.�|���\�<S���y��>}������!�
��'�,�ٓg��["�U�C,�a�fx��'�Դb��.����d��U��8	�'f�%öbH6Ajl0N�!y*�A8	�'.�agM^����׋�i��@�	��� h*��|h8q�S��@R�"O�4E�x�|�H".�3.�>	��"O�e+v�7e�̅��/�<��lX�"O
�$���x2Ԁ��ø0��p�"O6��"Lf�"�̃6?�>,��"O�8�/��``�M�w�^�"yvX�"O@���mI�.�!��D�d`��{�"O��R�˦��0�R��2V?$��CP�P��	!:V���/�^�6�K��r�!��"f8��b�ʏ&N�����L��J{!�GW��%�� Ⱥ_|���V�_N!�$ʇ@����(q �rL�#>;�O�=���g������P+P8���'�!��1e4<ȨF-�+�T�#*��p*!���vڝS�KU�2�<��iͥp!�D�F5(1�iM�D�y7G�	�!���;��T�^�h���*��#�!��J�9\%�Զ!��f@�ex!�עH��Vo���r��F4E\!�DX�X���g_W�V��ԥK4dU!�d�`�� kf��F�ʸj�*V>C!򄘊?-HL�@����Q��U*l�!򄌆A� �Ì�,Ͼ9d`E*�!�dE/w8��`iȹQ�P�+�E��!��^6�@�1ҡI>v̊-��B�]!��L!p8�$dצD	�O�{!�āY�
���ݿx�H�Di�	�!�dO6l���s�O�'wQH�mCM\!��O�څ�«?t����ʘSC!�dAjMjE
��?{�U���P�]!���s��t�"��vj<U{�lK9�!�D��J'<��C,E 	\,��w
��T!�˽$��e V��TW���g��R4!��þf����=;Z�!�>T�!�$�7E#`���$7h&�|P���[V!�D�.K�%_|Z�zAd٤|,!�D�8�B0�� �*�H��c��1!��_��
`�L?��B�E�&>�!���$237A�,*�\˴��,9�!���))BI��'�!�>���΀�s�!���)j�Z� �U:�>��6G��!�d� ]��i�؃#�:y
���+ �!�dʮ�pį8_+��@��f�!��B|��Њ��mJ�qv��� �!�$G;C�|���<��H�BAۯq�!�D�Vc�q�qV5j�b�0��">�!�&/���1Cԣ1�� )D;kX!���Y�&���d�l�5��!��Bd8A�Aŋ6�^͙��Dy!�S�R��A�A�ޭ`����J�rc!��sv��⚭c�$<#�fS�f!�G3Cg�ܘU��2W�F���e��VG!�A:��mksIɠZ�l@h3!�䓯1z(��a�-�DĠG�(�!�d��h~쀲�A� I:�r�J�u!��
?O��;2.^N<��@�%PJ^!�o@�-c���1u�|j�%�(I!���2���?�i��J�!��Y>@�<���;\0R"O�^�!�$�/o��f���BE�@-�m�"O@aa�L�>A���b�T6��d[ "O�}�F��S0�m��B;J���yd"O��cU��=[�V�q(�X�)�"O�ɉR�W4�2���-L�f7ֵ�"O� . b�a2C�z�9T��p5"O.����¥�f�q��ںik�Dj�"O�X��^�8!Щ����?Tv!�"Ovl���戤@�E;9�;�"O8�!D�&m� �X��֪m:2E��"O�$)dnۼh�90����$�j}!� �\�P���D,]�CR�]a!���7T8L�(�	�'' ����P*!���.m_�Q#7�ƙ<~��T+�r1!��1;��)rm^ X����)�
#!��!Ke��2a�y��ِT��>(p!��Xb�+g��_vM�qG�eq!�d
	0l��C� d��y�cX!�dǆq�W�*��뗧�t9�B�I�I��,�&��(��B�xRB�I�V����>��ٷ
��xC��4���hC�GC*uB�,D�}Q C�>!0�I�T��6��D�w���/��C�	�Xu9{��W�38��1kԃY�:B�ɫ/��8� L�	3G�CQ��b��B��Z< gEU#	�6���O~��B�ɰe+����c_�L �'$��B�I V�Pp$l��:����wᝩf|�B�ɕNA��yf녕��}sC� �/��B�	�a���s����4
�Ղv-�%��B�	;M��]�#�	Z�^I�#���*C��^�:ub��
1wpd�Ӷ$�2#'$C�I�p�y��KJ�/Z&�Ia.��j4FB�əI$V�i��r�"����6B�I7]
n�)Y!Z ��RL{��B�I<Q��i跦Pd԰��r�B䉖 
5�u4hm�P���T�?uB�I~>���biNLӲ�>yF�C�((M��{$aʫ������|��C�	�@J� � ����i0M�	>^C�.q��B�ѡv֝qtN�X�2C�(�����K@�3$�1���J�C��9")�8�,[�p�3��U���C�	�k�j��U�N87�HI�&��Q�C�IVPT�E��{K�	���խc�B䉻E8l��dƑ�-�5Ȇ�Q�U��B�	��&Q�K>Sq���С�$J�NB�6s�� @��B�}5rLA���_uB�	w��l�D�Й ɔ-qp%L�;�B�	�7�̜�ӂ@P�:FH2Oo�B��2l�ĵ�����w;�Yq��8U�C��L�,ra��\������>G��C��<(�5�ጅz����&nS�	�B䉠��y1�OH�a�P=#�B��+B�|Q�B�����bI�i�B�ɀgj�U�;l�Y���+^��B�+=�ιs�nE,$��9yD�@-.��C�ɇt��8�P�^���I�R���C�I�lV����	*/|]�ph݌!VB䉴ozp=��HѾ+M�1�S���556B�	89b\,�ӁT�鴹e�M�l��C�Ik�f�U��-�pq�2)�C�ɌwTY�e�O�C*��gT>C�	�|�ݹ�[�| .����π
2C��<`�����6yz�р`�,|��B� ���4j���B�	�FC��3�x)(f�ˁBy�����.٪B��<�f�N='��5R'AR�,�tB�	�h��cN_�.��K����C�)� �YW掞_��,�u�K�y{�hy "Od�bJ�T�n������#t:��"Orq�(Lv��(��&d�H#�"O�`�S��,4`03��J6H�6"Ovm��	)P**t�ѭb��1"O6�"�
+��@;� K�^\�Գ�"O �j@ɟU��õL^o&���"OBl�dfRr��w��>D,0""O\	)a��;s�(q3B˄�f�ʡ�4D�l�6H�2�l�H�,UJ2�]�o4D��#PdZ'0�P����'����A3D���q�J�ьGo��H�1D� �G
Ď%�v�c5�Kr&aȡb/D�$��SyTܵ�1 ?H1$EȖb+D�h�ī6{ Ap���= *��j.D�X�ViĸZ��2�̆��4,���+D����
bW�5j�؇8<<d"�)D�`�TD�'M�v��6G���V��B�(D�hj�i�?r��e�e��R�D�Y��4D�p���$E.��%H�#��1D�����ȻN,���.pR�J`k/D�<Z6�X����b�j�z�;�k(D���!� SF4�!HD&d\L�'(D�,�Rg�
VPPr���;Nh�Sp�#D���F� �R�AB�J1m�H����!D����
�=�
��"#�z-�E!��=D�8#�o����L�G��-�����.=D��I2�ʠxa�ţ��ҝf�&fB<D�@{U�a(�� g��{'(�E@<D��Cˊ����
`#�5��3�8D��`6-�+`
,�Ya�@����{Y!򄖁ba����,j�
� �3I�!�$`�%ʅ�(dE���.�!�m�RB� 8a궀�L�!�č0{��bJ�K��رB�Ф9�!��\2]��,C�{˶�  Ɛ)Dn��$ˠt�6��5�(�`Se���y���?�z�f�,!W�1��dY0�y���y��h�tX��m	��ٜ�y��L.xU�<[s�Y�y/0���@A��yB���K#T�+�� x����Fmŵ�y�)w,^�@�D�6m��1�vB���y��|o&��4�݅J�IR�B���y�j6;���P����3�d����
�y2��.7�Dt�a�ƛ �D�S�&^��y�K�<BD�[��wt����I!�y���I��(���F���J���y�A�1��j���0HO"z����yb����r�"�9�<��EGX�y�,ۥX�L�AVo×^��i��`F
�y�$��b�l�Y��٦%�D$�a�_!�yRk�)*�U��8)ļJ�*���y2n�mz��11b1 ( ��m^�y�+�2N�X��չ� A���yBF޼�$����~0W
ڏ�y)G(͸0���$��|2C/÷�y�m���h��
�����y��ʁQ�"�p�%B�
�J�j���y�i�A�<����m�@���y�KX _� �G1w���c�@+�y�.f���:���`E�
��&�y);q�*y�m@0RW��:�@	�y2�D< �'�>��� �����y� ��ʀ Ĥ�2	������y
� R�"a�kr������[�0LI�"O�0��.W�P�b�1@�R�
�"O L�sm	,�mRl6w�\ �2"O��B1�ɉ4(���լB%v�@��"O����-@P�Ybe�7Rr�]В"O�D{T�O�G���ag���(��EaA"O����9;���x���$LHം�"O>�(�26�&]��	�0%0�1�"O��ytŊ.�$�#�o��F�H%��"OX��A�N�~H���)C��-b`"O�aC�- 0�� ���
b�}A�"O�Tp��֧{5V����,}�ea�"O�`Wlɳ{�e�!,Z����6"Ot1���ۧxq<�*V-،#�Dl��"O�]F�G?Q�� UF �� �"O�qc�Å�Z�z1�E���3�"Op`i ��7.�@�S��0Mi���"Ov��!ҳL�1�_'����"O��RV
[A!d�jm�L��
�"O��;&K�#@8A��I��V��%@�"OP�8T ]�W�&�ZV���]�v��"O�dG�5��m:V%&�t�w"O�Bg�.#Iلc��>����"Oh�R��
�ƾ���oZ-X��ih�"O.D C�Ԓq1v�o_�O�
�z"O�|��`�\DD��*T��0qc"O���⣒!V�7�����K�"O�p#��ݪ=a0�9�J�=@��X$"OB� ���l���2Qʀ8p���G"O�$��4U�}K���7n��a{*O�E�H*�6a"�0K���a�'��lC�e�_관JC��1J��#�'Z���Γ.���IS3�BՊ�'�Z!k�n��T�2� ���i�'М��ĕ�`��q�2��`�
�'ZИʀf�]�^TXdf�s)&� 	�'�h�aƪ֓5s�!9�G�n�L��'�4�!�Ȭ~�z1��l�4lB�ps�'&@����F�18�`#Gܓ����'�=�tU*|\,�R�S$}�r���'˖��	�[��=�uE�1%��P�'�z!H�!�&*=��`�L�(ۈ���'鄡��J
���=C�̈3$2��i�'YlK��;]9��RIS�T���': 9o�c���c��Pͣ
�'�$(��G+q�Vh�ra�
~�6�S	�'0�dc2� 	?���q3�F�}~�X�'�<S��8q��Lb�
�!D$�#�'�&]�PHP�Z�ƭIM�"��'���Ɛy�\����
�G��I�'�P��LX��J@&9U�PK4�C	�yBϙ� �X�[�K�^��$8��5�y�VN�H�C§@J�\�u��"�yRi����T∘�aݤ
���yr��������e#��c�!X��y�'ڐ��p��/��1,K=�y�� ��XQ�_�Z��a��y�\�\� �P��2��X��y2��Xp5zu�-�ni�W���y�d�!��	ɇ��[���ig�݈�y�&s�P�c��S��텼�y��D"P��!�*�M�h�A,ܕ�ybm���8�b����H��;a��/�y ސ	S�� �B�FI���M��y
� !�W+��p�I��g-@,��"O"	ڗH۵�p�I�g�p�H��A"O6,��Ӣ���牨N����"O��� ��<Z���94[�-�l�d"On���֞T�xl� �^�B�^E �"O�12AB��ı��Oߕ2�~���"O���7g�/(�m	�M�)�Bɑ�"Ol���+V�k`��+r�*I
@"O$X9�	Ē= ��&j�$lr��Av"O�i�BI1(T�R
E�i�Vm�G"O
y)0��6 B:`ȕh�<1����g"O�t��M�e[�A��I�F���w"OTP�L�Y�6 �+ˬ� ɛ��	���
5��ȶ/jLi��X9W�2�"O
�Qs�4g~����F�l5�M�A�O8Fz���юs��x�v	�!���� 
�x�!�$�p;n%XG^sÎ���*5�!�dH�#�.,����!=��|��(^�qu��,F{��O���H=�4it�ݡH��(�"O<� 'NL7�b�J�S�0k\A�"Om���A�u�d3��Q^d�As"O@�%�e��)#e��n,�9��"Ol�F�3�� +��|�R�Z�"OT}��V�5i�I�!u�h-S�"OġZ5�U/P���N T5|���'�qO��v
E2
����R��-\%�T)""O��"@ ��Y���F�5"�i�"O08b��C6�&tG�Ɗg�@�"Oxa7g�j�^��Eb�01�
4iq"O�M�r*�V�,�A$�?'�-h�O�!qR"�T�����{?z0��1D���S�_�&�R���/m_fxZ�/Oo�m�c����W&W9B9�Ve
�
!����@ a �m>ʽt�j��U�O
6m7�S��t
�yB�
��pՠI��ꬄ�_�Ty��ߦ%�d�A7�t��=A�4+�ayb뀫&#}�֤�'?�l�PjM��0<)��䌪`�8�Z�fY�{8օ)��#eX!�D�=-.8��i���t�¥5E!�䁴*2�*��W�@Z]"�`�U71O��=�|r�����K���ޖ���)�^�<1%�H%DR*�B�BR4	�*,���K^�<�c*�0ؐ�uf�'�2��D 	X�<���<WgPd�񥃞a�P-��KU�<!�D�;0��$�F0r�Rq,_P~R�O����]� 9�T�o+Dl��/<;qO.�=%?y�s��<A�p�*�b�q̈́�8�)%D��Ҁgl��y�"��BHdK�*�>	O<�OTb>˓��"�ل^���T(�r0"O���OG���%훧<���[��W�<q�&P� rt�+JC�h4`P�g�n8��Dz"/`� �t��:��a���ըOq��i�0M�hB �3�X�3��ɡA!�$W2i���C
.(����%r���	Sy"k-�?�O45j��N�Z���`�����Q2
O�7��y��x�AS�[�U���/��M�a}B)	eHt��*���0���p<y�y�G|��hD@��9�{�&	*d2z���"/�͈��H#�"�����&1���!�	��	o�'s��(\-~66,ZD!֋n�h��Y��)��B�MZ���~J�iڟ'���<�)�'*��2��J~��m���E�~����]�'*I��h�A�T�����}�+O��d0�OL�i��^j��2�A^�V�jW��(�S�g�? �	b	��N0�k� M>W�ʬ!�"Oj��	+,����R:`�z��I\x�$X�lΡ!��'۪Q�e@�>��W��ħ=���C%N.hH>UUD�kjXч��P%`'.�vpУ�j�/��<�>qד� T3��HPb���ꀕD��@�ē1�(���=
k�`�G�D	[:�[DP���Z�Sܧ�y2�Ȃm�<�i�	o�%3�CS��yR�h">�xe�:o($@qܪ���?)�Or7�n� �@�����`BlB��E�Q���^z�'�Q?�SVl�"y�ƍ�R%��"�.D�����!5�\i�'�]!0�� �$��>I���
6�N8��~�ɹt�ǭC!�B�I�5?:��b	
/Bn��Zb�C+D�B�	 r�2�X��4���`& �0�C䉠2�0P�"Y�Y�PY�D�1�R�O��';ў���F�,���V�K�!A�>�!�R=f�&,�Q��!�����ƞz�!��L�p\��#���&%@��Z0v�ay"�I�p�bYkҬ��BT��ML@9B�I�X ��`���4p4�Ij;�C�I�q�2�` �� @hBaIz�C�I 	�`�Y"���$�L=���H3�"?i��I:_�~c�B���������=AO>��DAK�RT�I�ҠB�\b7����y���
=��{w`NP�!�&�&�O4�=�O.`�F�_�?W�$���jA�z�'#�	�@jW�B�]3p�Pj�b�It����E�OF�?�փ@$�eY�A�4�D-���l�<)�A?w"l�'@^
8�LeI���埨����8�v	�u��zU)~'@F{�OT0��b�S�[<�Ͱ�o�>h\�I�'ў"~����(��م���!��_�!�ˡ�⨹d��#��\�h�F)�IM���e!CF9nLb2�G�} ��'o�$��5G�bTL�1��9
�hC�~!�䟓)�ڽ
6�ܬK���ZA�Êb�5ʓ����q�d	=s04���(6�p�"O*��E͜E�B9���E�v�9!"O�0��jɅ'(�����(z�f5��"O���fʰm��1�ɳ��P�P�@��	�%|&�A EՒqm���"X�,��C�	��r�� &�HЬ��"X+HV�C�I e�rU��E<=��4��.*����>��\29��Q���4ܱ�y�<�X@NֈS�k�txƔ����s�<U���'�^ҍ�q�v�"�fm?�H���O����ڙ,����B�DE&�HV�A�!�R)�����G �6�X+] !T����N����ْ)L��{�@�R���L%D���C(ڒ(b��"�n�<}*�$%D�(p��_:#��)���:V\�|�%D���q,��|X�@&MO�=������!D����I��O`������;-�Xڲ  �	~���'m\�����E/I����*��[�И�ȓ_������iLFEHe
F�6�쀗'��ϰ<��aT�A�FЀ6oصtb��tx� �'t��Kpg
�E�X4ǯ�Gm�*�' �ĂGL�r��q�b�F�r��'�|}�R�*g0l���:EY��'�����5(��,��
�7�;�'�*��BLM5��y�FT�8L1��'�:�s��	�u&)#�MR�w��Z�'�\+���*�Љ ���@�p	��� @�Qq�&Q�jI��,�:�\��6"O"$0�B�:�$ cl �m�䍨�"OT�����[+�Đ�@��Lg8t8"O�` '+^��a�ga��	NV1�"O���OȐg�>,h�@%?&�8�p"O�P�r���b��`A�����"O�y����<7���	��]&s�$��V"O�y`��-zp�W��6z!�Ď�w�����ԟJb�hG��H_!�_�b`�1��ڭ$n��sg ]�P!�Du6@ݫ�J*vW�l��؜M]!�d��5�61pm��uޘ�T V�SU!�������8g� =�.Մ	�!�dXL��: �ׇ>HaKӦ���!�$U2^Z�R��YYl�闦��!���5kళEB�5?YV�eH\>C�!��Z���8.*�x�'(�3?�!�Z7�i���V��Es�!�:>�!�$�.B��l�� 8�خ�!�$��N��
�iC�7�rŀ���'`�!�dB6�z��g�V��:����Dx!�D	g� d1�ꃿH��m� ,L�b!�D>y��0T�H�.�ٳ+=6)!��1k���Wb�I���R�k��|!�C)��1t >cH^$� K�	!�d��$����7�Jd/�+W!�d_+Ğ5; �.Q 0Iћ�!��,U7�+1l�I(��JB���!�d>9%4a��n�.��tA4��j!�d�,L�§��U�hT�"�!��m^}�A�F 5}Xu��Da~��G��T �L�����;>l!hb��	�yo�m4������d��©��y��O��>,`p�	
O�:��1$��yR���!�P@�^lX�}
	�y�j=
�q �/g���P�a��y���,����p�C,b
#(S��yb"�1�¹�O�hlX�:���y��Z:w��X�#��o�v!�b�ن�y����G� �f�0�H�s.��y*��p���@�*����B�P��y�O��K�R��'hܱ%��Y��Q0�y�B�
u,x��JZ�(A�@)��yR�Ί�J��q�ЕJQ���)B��y2n�I�L������v�D�ƅ;�y���m��P0��cqLIh��yB�N?in mhҮƞQ�z��m
�yB蝡=�B���$>}}��zqΏ.�y�	���P�{s ڍlNҜ���U��y2�=7��L2�I{�LR��'�yr"ʥO�d�t�C�@���r���y�*/Z�"�=?�h�s#l��yb�Nv�s �_�>���ˢ�V=�y��ܞUܩ$J�>�r���@��y�.�����ӵ�K6�}hd��2�y��&
 td�4y�HP��CH4�y�'�	{������!L���Pf�+�ya-|Vf�fIXä�4�x�'/f�`#�:A@�5)\�k�`p�'ˀe�r���B���킑YUQ�	�'3$%�#l��uSV�+��^�H��͑�'2`���,�:_���n�8Z^����'m ͘ k���
�j�J���
�X�'��	(cK%D�DP�Cݴkp���� ,!�DmA�^�e�u�D�A�T��"O"(x7Mհ%C,\h��(�xKf"O�9	q��M���xvm
�^���S�"O�b 	"8��ᇬ� �$��s"OL(i�G��A2�J$��rT��$"O�C�J'M"F(ud̗���8�"Op�ȝ�)��(P^�8�m�6i!�䍖x�FeY��O�z�q��J�e\!�$)��)��U	)��¦IV�!�%rR�	U��5,�0��I�X�!�d
6e������Y�V�|�)Ed̥'!�d]��`�����KN�m�!��2a!�D��t�cá�6ARr�I �f�!��0Z²�R��WZ
-�q�M��!�d��l�l�%с,�C$B�6_!�7G��Qx�NO	qpi��oE�{	!��.�� ��(n�Ԑ�6m�$�!����ċm^yp�!�a�G�!�!�)K���ĪH����2�Ѱm�!򄔕bI��� �^`jp�T!�$]�O�8�`l���%[��N�9�!��ym<�b��4GR�T�a%��[�!򄂭u� �uM��a[�4�W��g�!��Ҵ^
n�b�hҺq�G�{�!���<�H .�Lq���9�!�$���\��&W9o
tH `G�v�!�$^3~�y"�L�"�Da���!�dޛBt�,0fn¿`�a�6���.H[�g��A�̜c�)K����s�J���B��@�ʴ���ѽa��9��f�?L�@q�Ǐ�i/�6�'�J��a�55�0��_/߾�+��$�j��A�����|�.��U�" ������dK�;��أ"OZq�rIY'jq��R���2Ơ����O8Y��'�2$�V�7�:""�n����1a�i4��:�ŜT�<���9h�J���ۍ{��Q"�H\b����',�͘��������O��@��5<OB}	�II 	;����'^�z�ś�0��W.ά�^y	ă�`H��R}���ʁ��W8��hg%�"��D	3f�hu���)��p`�U�-k��q��U�,�R�� 53���n���c =)�B�I�8���/N�x��*@��僣 @��R��r�I�*�p m?9
�|���B�@'�/:.L�{t��dxB��m��]-Tu�B��	FyI�E�_�i��My�e�(���(4�'\��瓕5_#<1a�\:n����;{4��Qb����Ú�VF\<r��]�{(�q�g���c�\2d���h5/�}&�A��O=��!���4���B�\RBQ�$�B���P�ABP�l$ j�CL�����&IA&��'Y/L�zb�
�m �:�K�jW����[���LЄ1��)j��e��խ�_�QHK�!`��]	��I�Y���2�w� �9w�J`-�2��,����'o��с��m�}�₝"v���W�XjX���P%.$�uA���-���%F�O����oʆ	]�B��4`)SR�'B�<#��1 ����T�$�<�Sd�	�>E<�5��7>�hd��B�Fp���C�'*N}p`U��0A�D�â�1[���2ba@��� ��3��I�b�ǆF>4s�O��a#��7��9�Ө�+PV�1
�'�2�������l��E�/�I�F���� _{��L�"��t�.a���5�'��q*�@���JZ֢5P҂C"n����b)�O4��k�9R�4��C(?16-(��-"���u�/;��Sq�*�IH�P�6䚳� ���I˼��P���E@�  !�E1�J��$��68�`@�- ���mI�0 �7h�Ar�P��pȶ$ɁA��As V���	R�u겥{��X�g�I#s E+e.dG|�]7vJ���c�<kg� sU>1+a�:?�:9r�BTBg값����'���!�G�q�g��=�` E>x�X]���N<Z��I��O��W�x�3�V��������Z)�@���&�i ƅ'5ظ�M:�a~F�n� �3ul�)T�,�zB\2aqON9��O�|:v ^�f?R�RAS~��P�4�� �U�a�a	 �y
� �y�,�1h0�S6� �+��覔�8��LNp��)�2��
0JF^�����E.���u"O���0 N�(�����}rF���ɩy`�D�%�3�	1V.\�`̕.B�A�@��6
B���Q �D�9�>�	�Yh�$�{�,�.{Fٲ��3�OT|��h�;#��ktS�=���E�'�TP��0N/��'&��r��%u̨�Ռ��_�z�'*t��fi��%C���6�ݪP(:M>��]�Q��>)@w3���eVnFBA�v�<D��L4z�X��"��+�ZٓQ-6D�xseォIr@Q�D;�E0D���0BE��(`�@*@5t�����/D�TCQ�By"dI�[�Ej%���+D����U/H��0r�X�Im���O)D��[�Ag���{� �l~�S�=D�L���� ��]2EWt8��8D��z�ν הp�4EA�Z|	�(8D�@S�,�*'�)Qg�.H�0���9�O�8т♴�M�%� #�.���iL�f�d���Qo�<�v��
�
��¨�=b~��aS�'Ҝh����b��>-J�aʤ%ΖȨ� �%k�l�`�"Op8�RmK<r�����Őqޔ%��-к����O��S��?�$�F'5��E��/��x��Ohar�?�)��<�CD�4<x)Ш�I&n�r�B?��K�C�h1#7LOA��j�=m�^����M *8�E�G�'�����KՙL�Q����_}�]����`�x���l��#�h��CL�a{b�S�{f}��)P��(��b��W�����D/\Ր�1�0ʓ� �1�T�"|B��9q���ґ�*�0�J��c��U#gHM���}2����D��pei�:�S�D3�b��E-P�H�O?�Drije��}�� �n�121J�@W&פ���'fh"}�'�^��A&g�y�2�#Q2��H�'�8!����}c���	^�l���:z�x�:#�P#s$7M�,t�d<9�]ވO��t'�JZrᓅ�M�!��Ϧ*ƙX��	��=�ĢE:g�3C�O~�U�.%8��+O�4���d�	%Z;�ĂF	WC�O�@��,;��}��� ���A�}��*g�L0�	k�O��0ȵ('k,d�GN[�[;�@�ٴ�-�$�E�S�O�x\�K_� BG�N�,�8�`(G^�*	�� /}R�0�g}� � k#���nҮ�����y�+W(u����
�(m�dl@��p�J'�ٚH�hX3H���:��@Fx�/�K����$�+4�4����0>�ѥX� ~v��s�  g�)����q+�ct,�Is"Z�bj�_��\1U�[�4Y��˙l��pp�"%|O���)ȆD-XT9u��)Ng�JuN'Y"�ze�ۇH���T!��i� ��jq�g�r����c� ��2{�4s��%:��fO@���7!��9�#��.o�Qe� sA��ȓI��� �1q1��s�D|��X�����ή;G��dN�5з/u��~ω~���*ɤn!�ɦ���y�����L*4���<w
�a�0K)�����"e���C�g�'�&�2$�3I�re'4N��	k
�Vsh��2%�(�Rt�3#�6E���C_Y�Ucs/�+"b/3�O��1��GH�$�Q[�>q����&m�t8C�#��%)CH��'A��tbbJY�e��`f"�&5xؼ�ȓI�n	K�%��Mٺ �g�l���+V1^����
vs�aA��~r�/?����s��.<���&�B�I�3��Y�c��)�|H��C�U^D�oڳ6o~��p��*�b@�6
k>#>���H��m�C��<`��BQ8��9��LE(� ��[r�<��Z35|�i���\29��u��c؟� �ɣ_� (�-0�#�#O�ز�4t�|rȊ�p� 
���&+�����_��y2�Ž50dyð���z��d�.��I)I/��(�����&b�A g�38RĪ�.�l!��E�xS��ŴY'����b���!�$Y|�䰘��@Y�q��#9�!��;xO�=�%�J42���#�!�� ~U�D$�$>$h�'�cs&Y1�"O�P��&Q|�9ru���#a�k1"O�%�f��`.�p��OmD�jU"O����!EN�l�� өIR�8�"OL���\�`J���L-1J���0"O���W
^�"�z`�3RȤJ�"OJyP��Q1"�0��اOJP"O�SJ)	m����Ȓ+R�C�"O0��P�s��i�'f��3F�5ʣ"O���,��@��sr��%h��e"O����!7svraꉂ,d���"O� �l�,%)4�2�L�g_�0av"O^ぢ�0�H��C�G&=��Q�"O�Ź�	ۑ	 �d�E�Fd/�1�S"O½�Ė&P�]��J66 艰�"O<� �, @���eb˷	ޘ� �"O�9$$͘FS�i��AP?b��Z2"O\�9��,k�f�:�]�R$H�)�"O�}�� �ڄ
��'��g"O��
�(�$ �ȩ8V�_9��sf"ONiQ��V*.�LD��]<�Z(2"O���HZ�Ry|���H�	���H�'��"`eر:́�I:S����'
`@�nR�%����Un�U�B��
�'s���2��P���P�
G�V�H��'a����#Ґ9��1Tmͩ8���Y�'�X$�V��BB� Fj��G3b���'��#�s�@J�/O�:zPr�'#@�(&:���P�z����'R�ySE�2+�����xa*���'�`�L�	6���t�Op�1{�'*E���?�hpУj��d)	�'�b5R���2t����NV�����'�L<�HЄ����5�����'�n��1'����&V>I��J�'�DX)�װ ���u ��dK�t��'KTT��O R2D��	�QE��'u��H����1�%�6�R%�@��'���p��Y1U`U�FE�&�0d+�'�F�p���g�:E�ĨJ�{��2�'U&p�C��#>4���աG����'�t���M�� �h�yF���$	V��'��=YG�A�fPr�PHl�
�';&t��ߩ~^F,�s������
�'� �@�H��0ٚ��Q�(���'d����h���O �l;�'*zdc�nZ�|�mb�˩k?&e �'ʈ�fO^/|��� 56��T�
�'����,��l����ә< 0
�'G�(�C��	T�&��	�'/�Y�5��S���{��
�=_�}	�'�fubP��Yn�%�=<�	�'��D��یPh~�2���
�@
�'(�U��7h4��D� ���	�'l��w�x�G��*+���	�'��u�F!���x1ʔ�Flvly	�'�9!bG�=a^�)��ݞ�2��	�'�(JЭ�~ܹ��贽i
�'��d���Қh����a�~�$P	�'S~�+��ɏޜ�A1�WN���'f�H�&��	���P��{f�h�'_�`�w����Si����
�' �VA��1����aC�s�ؘ�	�'�z���-$�0���`��q�	��� ���j�r���b�/���*�"OFaX֢Cu�>B��N)y}ʰs!"Ov\�VL&i�B@D� kS��"O�.�i��)E���ebf"O�zQk��jB<�p������Ѱ"O.�����*��`��Z�V�](Q"O�e��E���f(9��=}Z�[�"O,����7kK��+���%R�Ĉ�"O�Y{ӯ	��������z�5��"OʌzƀDi%�iR%F�x�T1��"O�((A���_E84	@�#��e`e"Oi��GC�����$ށY��� "O��8EGǺ`��c��C�ta"OB���l�}~2��Y�!�Ȅ��"O"�5�^�
/�us�&Yc��X	R"O�����������޳>6X<�"O��I -՘'��;�M(/��A"O�	��㈵$�<�Yd��.w`�"�"OJ���8Z�I��D��(�Q��"O@�R�'N>8�<��ї9�1�@"O�`�����P�m�7$�$�Pe9�"O*1���k��Q�QϨx �"OH2��Q�Q���(ClS[���"O�łT�*g�\�Eu����"Oz�kf`HC��ѐ�J!龕C"Ohy��&�	:���q@E�U�'"O
�R eN
O�$Ye�ݡ�"O���Q�'�Z1��o1vZ�r"OLh*"�\:V8:�2�^	aJ�(B"O: �0�O*�|��	V�A�"O�M!�P!#h�  N(3H0�h�"O.�A�銷!N�L �,�[%y2"O8��ЪS^����L̳Q'�ݸ"Oȸڇ�(`�1��jRR*�""O��Â
��lb��Ac�+<|�F"O��q���	&U�E+%�+Q��d"O��P���$a�M�g�O\���ِ"O^�H�F�@�D�f)��H�J�х"O�t	���J�8)J�N�"�N]�5"O2�"�J
,�`���7rt�h"O�����Z=�dz��U�@~���"O ���	��ui���0��|��"O�RQi�:d���ە�ǁu�rź�"Ov��S-N�;�xhH�#��t�Z4�we׹=���C��=�ܔ�����	lȺ�c��H=
Z��+r��
�y�`��x�!�ت-r�ґ'�8�ybɇw�����W�}f���	�.m8�a2ʒ�e�l��E�8,bB��@9X��B��+-j6�f�=Zh;��ݠ0�e(�	�b4.C�I �.X��Ř�H@!��m��̳�M^�1
hEJ��:#
�9�|Z���_+r�c���r���`��i�<AS��/w���*�.�F��j����6�H���I�w�:0:�^័F��'��8��!�9d�*(�2U�i�ҽ�'��ŋ��ԁJu�ݒ$J,ֽb��Y@5Ȥ'[/K��Qa��*�0<�Aʆ4F4���E�lch�i�f����Fƀ�r]��J�7;:�){�/�Z�( r���ӣr<p��$q9�(0q��< Va�ITs�� �0�:���O�jL�"����O���6ϒ�'B,�H��\�"��9#
�'�J�㒧�W�C1/�4@Z-ٱD�-~4p��ϸ�XE+��h��,7�H@`�-�<~:j$� �Χ	[0�b#ʄ��?���/I*qZ��'�����̓~���zq�Ԋ{H
�y��<a�j�P.�)!H���� �v��Xi��A�H��|(&�!�O ���	{,(h���2 �@6`O!h�P���N�~k�=��I�2a��8��ӧ�O�p���^�e��'�2Eb� ��d��<�|ɫ׀,�A���2a�L<��+�G�<n!DK9}r�%}:6��}&�� �9���p�Z0Y�`����Y���Ob����I2�����3�.UX�T��f�0~�ek�DA�J���U��0?�C�Ҳs	�����Sb(�e�@X8�,�ťmJZ]����dq��)��o�d�pD�F�&D�زa-�(`SR�C�L#Y�H��'}�$YC�X{���O>-��]��!�V�{�l�@p�%D�l1�F#K�h����qu*5` g�Pm0�'��L*` OB�g�ɘe"$Z G՝<H���DA�wd�B�	�3�<Sc�	�%ńd�0Oǳ%��Q�G�6��$JB�'2�x�G
B�;�ܔ�F�,w�,C�Nu8�É���+�E;D�I�1�LQ0r�Ȕ8 C��5��I�Oqx9�#�'��\�d�0���&��T،{��3w`+!_,<���7@��}��'�B��Vn�	k9��"5/FyX�'< �C#N�/b�4-�j
*%t!�
�'&ؒ�O��}{@�-S XH�'�1�C!�	!�n����fǂ)�B�� <g��ӡ��)-�-��CO�C�IA%ԁ� ��?/���@h�3��B䉻)��ݻ`˃�UA����F>Z�B�ɞ>�� B���V���!O�x#lB�	&μ��fB@3UUʀAP�,~�n��Ė,�j�iڴx_d�°��>L2��&f���T��$@�k�m�0+.��7�A/U��Ez2M=�ʥ٦�]�!B �&FV�W"��Y��B�I�>/F�ȶEָ0�B��CG��SUv����To\j�##$}���'�@I��X�8���0�AL*k4���O�`ۊ�=E��'M�y"@iG�;��0��P� 
�'9r�aD�X�$��Ԅ�	t*�Q!�R�y��z��������`� Q�'N!�v�b�!H��w/�Y���;����S
�l�x|ã`/lOH	��-�l~��wCp���W�e��%j����?mEy�CrOn�����`�OG1���E� !���c- ��`��}"k�%\5�4q\�R�}���1\$z��꒔~ ��
�	_���"�-�$A�O?�DS�ah"@�dl҈�@b@�V�J :�xF���H�"�'�
"}�'�������>����X7$	��'~���gǂB��I��ɺ�n�	�A(e8n��U�6�,1�hl!��OL�s A��4�t���#ٲS(F��ϦO�x�2͑,а=ɤ鑭wN��U��Ox��.��Y몕[�&ǣ3>����O�]SW��l�O,^�;��M�(�&aHs+�&��s�}�	&@�H�8�o�N�O�ي�&ԮT2�"��"מ]��jF�Z 3�)���e@)"Wd �! ��w�YY@@؟+W
�2b�>���>y���V���"f��:|N�0�E�<����}�l�a�٩�n��vU�,q��7��B���O�nE�x�"<)��W�-�H�g&ɽ
���:��v�PX��U�q�ĕu�ja����Iu�����]�K�󄖶C��tg+|O
 �.o����+9t�D2@�'����3ǎ% �
 G��@ г�OU���TF×\� �x�Of���k��t����
�A]䉹���=2n�0��%]4�*wM�U�ӢQul�(�쑎-4Ь���f��C�I�l�0��`���bB� �������j )�qF<,!����j��>��(X�
�i�1X�h���i�w��C�	�s��:`W�)��
Wl�Z�l�z1G-Pn9����s�2���Q��;5�
��H���'��!�O!|O�i����T���l�[8>ё�K#i}�xǠ݁-���%SȰ?��G��0oh��1p�S�KM�un�A��� >d����n��1g ��5X��¬lق�T*E�D���"O6-�����`{R �ֆ�
U�d賒!��+ d;��ia� ��>+�>�	4q��0q?�@�3�P	;B��Y�&t{EGr�h���/-� <��4n���Ε`3���Ŕ�|F|��ӓ>~�\��BU�#�*��3-�1�p>���N�ĺ�єDO[�����O�И�h��9հɈU�(��?i� �0��D�� ��T �1n�m���ԅ�= 4a$��� �-[Y������ A�Č���6D�D`&
F
$q���%�ܻ�%5}�E��J��I�=�� B�)�ǐ��l�J�hiJڼ��"O��R���'�`u�䜶q��T�6"O `�'�MIFD�6#�,��Rt"OB:WK�\���!,I=|��pC"OJ|kb�%(=R�����Xr�"O�Hs�̒04�vM��aS�f��A�"Ovr L\��8У��W+��蹅"Or���	42b��Շ��JH(!"Op\rO�� ���df§!&-H�"OܸcҎG(�m!T�6�J��s"ON]h@�B�h�a�#���.�`"O�(����[.H,���׷/C�5�$"OD�KB��G_
̋u�V�;�!�S"O���(��<�Ł��}+@�e"O~]�(3=`���gԣAON�x�"O�Y�蕯0���9�fu88y �"Op!q4*� �q�w�ֹ)��Au"OU:%
=`)�u�Ū�>*�yW"O
�@�G�#J�d��?^s��"O�)i�3^���# �[�poZ�""O6 b�iߋ6���lV%h7��w"O�����U6e�*L�R�!O���"O�X@'���D�Μ���	����"O��1(F��z2H �P��"O�03��5x�r�6'ȕ�(��"O\��� vv���'\�rL:�"O��O�1Q���7 �*$�$"O
��E$M��u���<ZA���"O�Hs�,�=�^�u�3%�����"O
m�V�Mޘ�ʷ�g�P�˥"O��@�~�|�WFW�+��k�"O65
b��τ�"� 0o؅��"O�L�&B�A,�T�G�aP~��"O:%(Q@��l�.��o�9ej�*�"OU�h�_��-Q�/��Ln�aS�"O��ÖG�rV�Jp���!4"O�$9���!�(_�>���0@"O��8$nD�8�r�	�)Pٜ�2`"O]K0!�b�1�IDT�1;F�'�!۰�v�I��(�"�`�k�g\&'�'����F�"�f�Xe��	��'f��P�ӺE�T��X�����'b�"�K;>��M��܁9�����'���Ȧ�ƿ~/H�PB��/jh�
�'���Q�ꇽLF- �,wH0�
�':��CW⎔� 
'���	�'�fu�R�=H�Y4.����aL7(t�ԋL��1�O&T���e�!������}�thRqb:
^����
��M+a���d�LXŉ��q�"�I�
��hC�I��U���I�N��T�����Z>��O�9	���5������q� ���PY����'f��U @E>�S)7�5�`�)|��	H�&`y�H�5~����6 �0|r����&+୸M<-�������<a�"�
Ѷ��r��m�)�'=M�i�4�^G�����\/h^����d٦H���ha�	�k���)�����E�j�f���eƿ�0`�t��s�\@��N�i[d��,C֦�ZrN:� �sLU�� � a��Q�d���&оw�VA��.R���	Z>���J�7cNa�Q��9G�\��l�|;6��Ox�{��i���w}Z�M{X>u�1�д�<�ʕ��CR���^�p��4i,�}�M>��a�O�2�ö�B��:)��n��Q�	��l�qO*H���8[�&���ӥ1��zd�L?���=�q��a�Ԩ7n>�t;���77�t��b]���oox� ��%�)�S�d�v�gD���t̳FD�h�##n �C޵"CrԐV2r��G��c\�i�]k�T3Fpf�Z�hԞZ8�Q��Κ���b�(�W*��C�>��pk^/x��G�!W�(L�5h�e?q�#��"%
�WA"}��	�,g�A��]�>��XzS X�e~!�� \8�2"��R[6�y2ѐЄy�"O~����j>�`8�f�*U�ltZ"O���A�-u@���م*�а;"O\�1@�e�N��E�3�Ȕ�'"O�=�e0�����5iϮ��"O"tc��Uq`@Q��mј%k��b"O��	ږS�)�0�H�wi�!�r"O����[�_6*��E';YzA��"OT���!)�ޔVH(���"O�	���3816盳o��L��"OP(��9j�`0�F�,I�Tx�r"O��!Ү���̜)��^)u�,�C"OjXh0�L.Eई�����T�[�"O�ٗ�=[��Z�$Z�O�p9"OziRD��+�D#ƌ<f>!Y	�'Z�Y���|E2�b�,X�lA��'��ɖ�Y�����A��e|���'���q@e�
��}��HC�|�0�i�'j�%�셔N���d��A��$��'��eM^' �N�VN>b�0I��'t�t``�L��b�f�!N#na�'�T�H#�E��R�o܉��'�LRb
-� 4H� ��Pz8�2�'���5D9ET�-����D(n��'8J�bu�U*V/fݹ$A�9M6���'cĈ  i�"�H�B�H��o�u1�'�v��"ᑞ��r��]��!�'Q2��! ք6��x2�1b�4�
�'Z�8�s��X�<�%R��]	�'%����B2���&��=��9x�'#��R���A���&H�L����'`pp�Cڳ:�}�5�Z���s�'��i9��ؖ4�X����b��y�'�����:���4�ޛLV}Y�'�Xq�R�$b%��P�x� u��'6d�C��:�2��)[yf���'��@��+ 0��6JɅ!1���'/�\;qJ��&,IA.�	��`:f"O��fKH?IC��4HX�#���Z7*O��) K6  ~��s	��	c(� �'�V��!��I�E��Z�O�lT�	�'�سb	B&a��Q�����	Q�'D^q"� �	[�qDk��ͅȓ�.u���<��`e�"��܄ȓ9����bG+B�Ы2�Q=KǞ���@+R���a	�w�>����B!s�I��h4E��lZ�R���KW �=��S�N<���-�>9`  S�����ȓ�$��F@�i�⵻�D�=5�}��WB����Q&�+��;_�U��_� �4�4IXa����3&r�|��4?,�IWe�}�T,[�o�^7PA��
=�pR�mQ��ગl̈́l���ȓ��h7�F	~!ʵ

�L4�t��w,X���O;kWb}2b"�9#���ȓ}��jE��<ZpV\��a3�X��b��ᅁ�J�@��#2ix���5M�$Ac�@-W���a��]{�Z �ȓy 8�j��_�tF9��?"�<͇�0�@M�F��N�i�P�\�k�ꡇ�t� )9E(��XL攉�	H9X8�ȓL1�M�[�!Y����e�"���}��x�N�@�vԠ'��0(]�,�ȓP���r(C�Gct�q����A\t��S�? �M2g.Ďf���fز}�pTBV"Ofp�%A�*T�� �Ɵ�t�郓"Ox}��Ee������#1�xh�"O�рr'��/�ԘU�3�НB6"O
� ��6�
�*��P2��I�"On�imȍ)�隅FK������"O��".�gK�1Х�?VbR ��"O��pG�o��y"�Sf")��"O���p��v�;!Z�r
΅��"O�`C�*VF�M��LM�OU�X�W"OL�ɀ!\�I�>�`��.&>�Ց�"O��(im��R�¯3�L(i�"O�1A	>P�BY�D��"p�x�1"O�Xq�E�U~KcOI?<ަ�@�"OP�*��V�0�D`����[�J�"O�}w" azz�V�G8k��	�"O�$��d�=	!�6.Ӑ8�:Y�T"OJ�Tm��>�J�S���V�z"ON4X�d)"��Y#�@/x��7"O�Q���̲�f�G
��|��"O�� u☫6�
��b�Ԟj ܐ�&"O�98v�0
Ȁ�)F��]g��A$"O��Ya&��r�Y9� ԴEN�q��"O��)7Ò�����@N�_M^I�"OP ��jJ�L!�T��/�h>�X�"O��FM��7��:� �wFQ �"O֡R%�8`,}&/�4&	�F"Ot�k��?��	z��J�.c鱒"O)�F�T;/씑���,M6p(�"Ov�^-R�xi�ssHޥ��"OvPR�I'��I٦n�4�d�:"Ob���%�p�n �)y��Ї�'D���3�Q�i;v�t �M��ń'D���倾*���h���#{��pA7l3D��sd�͸�8Q��uxP�+3D�al�.� D��?�d��U�2D���wI�HY��D PRU
D�#D����/N�9/6=
�sK:�p�#D�t	&�̌L�r��D?�	���?D�XA�:^M��1�����`��K2D�̻@�h)am�(^������>"!�$�;{Qd�� �0W�NtX6cֱ!!�L�~���4����"ǼW
!�DN'N(@�կ�(?�$�kQ!�+�~$Vc�*s��YV�ě!�!��4S=ĥ .O,^��3���#�!�D��}�I�(Mgr��P�ԅ1�!�dN�;���b��Uc�ȣ�Ɗ3Vp!�$^2
����׈E�Q���O��z�!�(5خq&�Z� $v�8��)!��ܨMw�0��K;��Ua�a!�3H�8cl�7!���ײ|���'b=����S�*Sa���	
�'�(�GPm�����%��@A�t�	�'N����ʮe��2͌�f���!	�'�8%�a]$^�. *�&�13�D�
�'5� òF���ՙc@_�&���'�
mR2MV$�@eHC&��!�8���'Ѽ}Z�-�Zx�(���I�� �'�8H�"$M���BAI���@
�'�RQ4�Ůp�$Q@̓.KvQ�'|ؔ�P$��~(9ȑ�ϳl?j%(�'�|}�&�ˣ[�T����$iҘ=��'K���G#H��p�J!A�ct*\��� ����-D�MP&!:@��6;NL�� "O^���Y}n.�+4,�#_��Q��"O���`<`���'��`��"O��Ї�ڨ�3 �x�.�ٓ"O@���R��D*��G(pʅ"O(d0����xA�u�+Q 5��"O��cĕ�%�Ա��ɂ� {w"Oĩɑ�3Kr"��6ʨ\��1�"O��+�O#}mZYsv
]�� �"OH}�UN�}�,�H��}��	��"O�(�̍�$�X��qd�+cTAb"O@١��¶0I�<�3�$SP<�&"O�E�E�wo��R'b�L�@
�"O�bŪ�m:��A�o5��Q�"O�]��Q0\B`qt`\2�� Q"O,	���,�>@
w�˱�H�Ç"O�x��m�.nB����_<�i�"O�|p���K����a=#ܶ)�E"OZUIȆ\��iᢀ�39ؐ{�"ONYD%I-J�1;�-ޱT&�I�`"Ot�RD�	K3^(����p��"O,)�3�Z�8��X%$��=��8A"O���
�yb
�{�A�;d%;!"Oj���[��c �\	ڌk�"O ����A5Mz�x���k�"O<hT�V�!)�����w�Э��y¤�>oԈ,3SϜ�mƀ�S��_��y�:$���^,N@�� �y��X�m�����^$����ʏ�yR��-��?T͘)5��C�I)<�Ȱ��֭A�"�8��XG�C�:D���`�T�:0� �n65�C�	<0�@�$.�/��	����:6>C䉗)����`Oق6�1�+܋�hC�ɢ;�,ݳ��@ ��؄�V#nB�I==�`+����}��JS���&B�Ɋn*��)�@k�v��C�K�~?B�I%��Is��d��I ��C�I"i����Li�bϊ�"@�C䉇S�!������hӤ�C�	7hxx�	�����a�&�p!Bh*D����&T�$�`"�ڔj�Ơ2�/=D�����7	��R��Z�cK�L��/D��k�Gj�DCB��1�|@V#"D�p����$}B��1����d5D����O6 !��87�/5���8��/D�H�r�v<��
�g������c�/D�Ĩ6�ܫ!6�D�2c[+
Z"��2/D��g`Q�Wfy�0��/,�d��,D�ԡ�X�P"V���� K"�u��/D�R "�:_ �)Be���kw�1�1D�@hrL�#O^0����/7�q�� 1D����@(z��P"s�O�H�l�i#`.D��`� 9(q!O@qf���>D�0p��(��p8g!��)�`ɈZ!�$���B|BQ�ߥDu�Ń׊V�!�$��X𚅢v@]&^g�!��HS-J�!�DL�L&��iV�A�2��`ǟ��!����]��� H�7�
1&V44�!����z�i� =s�h`V�!O�!�O�r<v!벌P0�T���lߠ{!�D�)/�����"�#}t��넬=s!�d@LH���̗H�X����K�EY!�ГS�TI�-��|��"�H(HN!�� ��{�l0r�UQ��Q�:��A�"O���A�[6��c)�>cj|�"O��r7
�%V�" ���2 5�"ONI���֏
J�PJOݻӤ�R2"O$�    ��   �  U  �  �  8*  �5  A  M  �X  &d  �o  *{  Ɇ  0�  �  {�  #�  �  E�  ��  ��  �  k�  ��  ��  ��  G�  ��  7�  �  � * l � �  7' �. O8 M? yF O V M] �c �i \n  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
��G�I�&�: ު(�&�'L!�$�, �2UB�D�C�yDL0Iwa{2F!�I+=dn!J�HJ:<�� ��ܾB�ɖt\��#%ĪL�E��
r��"<���?�2�[$������8��!a6D��z��Z�O���
���< /��b��4D�l���+j�d��	Z��	Ԅ7D�x�Q�5zarD�3���X�q�4D�TW��V�}�S-��U��Q`&2D��E�*���c� ;�r�0�%.D��8ɝ� [b�����3!G�a��!D�芇�؈ɡ#*�./��1�e*D�(W��%M�Lc��v9��3G�'�D0�O�IR2��z�<eY�@;i��Z�"OH��H\�AmN�����H1�qg"OΔ!�N -
PA�!�?,1�W�'�ў�Ơ�{\�y�	A-e�d`�AO%D���F�r+蔹��Y#^��,� �?D�țufY?[���� ��[��x��;D��+t�+wz��P��P�w�-D��P�B	-�l�2�!]�%�N���&D��2��
��r+�j�'>D��Q�
�0di���W	::<�#0D�4��f�Y���E�3� 2o D���bG��Aʠ�
'g�X�<�: B D��y���?FD���eX�2��[�J*D�t�Q�́}����R շn��8�)D�TcwO�MN" ����ɨ6�&D���f+ăP�<�04�P' ��1�bh$D�Q��I�u�uď�Z|jX��� D�t;�a��܅j��#/�D��g�=D���ÄC��IC��J9h��9D��Y�@�
j	 �Y��ɵb�4��:D�,b��S��F\{@��Zk,(Ӧ7D�L:4B� �`���E��sO�m���9D�P�F֖[����!�aYH:�c$D�� )
���C�0j �*�h���"O��h�?}����`����"O�I�q���<��!�1g�6Ϊ��'"O��H�>zP~�9��� *�ђ"O((pS���Ixy���~�%�Q"O搸�&׷z]�!I��>~*��w"O�@yQ��:�^Q$ ߟ`pH�@�"O�a'�ʨl��sr�dx���"OX��G�0���L�&J��"OQ��T��!�aM� g�܉r"Oe5ɜ���Źu�[!`�\EkA"OVL* ���<�N��$.�!DRl|0"OF	�4�P�
�|��TlA	)-$�!"O��Q�Eq�� 7MƂ>���"O�0Ban�jc��a�j��LȆ"OJtj���8
.�H��֛th1"O��k��� H��j�h�:ԬȰ"O�+��ա�l-����D�"O"4Y0i�x{[�8l�p���"OT%�S��"�ԴrWAG8>���z�"O:�3�F��`K������(7����"O�uˀ���c�,!��d,�h��"On�j��@�8���� �n��=Y�"Oȕ@�ɛ��6X�#�հkz�4�t"OP0��Px'.S�]$$0�"O�h�a8B��L��-�0/o@��"O8l؃�	ϔ ���A�x�Z}�"Of�"��%����<�z�0"O ���o[�)����������h"O�1���C���5��u�4�s"O�0he�Q|��q�M"sҤY�S"O,���ݦL��$�"ԫT�RQ!q"O�D��*Λ-D�+�z��	� "O�U��H��%a�(p�OǴK�R��P"O(�c.�e��9`2Cθ�;�"O�y��&��[М���ŉ,!�8ғ"Opq�V�+t�F��⯁2=�f��r"O�!�cC�$���clNٙ6"O8)#�ɇ2��В��(-o��a3"O�)��R¦m�ҏQ4RN$�R�"O��h��މS�v9� _��%�"O��3�O�2E�Z�h7?�t��"O�ȋʽPd 9R5G 14��T�r"O~�8��|U���`�E�4}���"O~u�U��:"X�$��o��R�"ON�37����1�ؓȠ��G"O~1a%&�RF03rE4I@ ��"O<hjA�ŭ=)�=Z$��<0�t�"O��7�L	�ڭ��lC�I��U"O��CT�BA���p���-��ua�"Oh51u@�/z��)���+
�1P"O�pULS8�0���H{����b"O� �v�>h��!�	�d9��"O� 1С�&/�n�S��U�EH��r"O�����8N0|�U9H3�,�P"O�53���`��k� U-`���P�"O�M�O���� Q:���&"O�P�G��/-kR��U��q �ԢE"OEy�4y�� ��,A�fe��+�"O����#��)�B\���/d���'��AwmYvVܙ�d0-d�K
�'h���v�	&~-��ɪn��B
�'�ʍ�!�O�@�A��f�+
�'PP��+ޔ��=bAEѶ]U|��� 0P��N�2�A�e�،0M�9�`"O�	c�'��\�92�9]H�@f"OR�z�Aʪ/u�xp#�@�H8�:�"Omh.\�)4�"s/W� ��[�"OD�ࢅ�Z�} �H
��|
D�'�2�'M��'���'X�'���'�b\P�MѸx�I��R�R�0JC�'�R�'�2�'-��'�r�'���'���3��;�L�I��̓>��i��'f��'��'�2�'���'���'hr��T�L�A�N�{B)R��(�'���'�2�'B�'�"�'��'���Ck_w+�;S	��i^�lx�'�b�'���'���']2�'T�w��a�a/�D�Z�D7iUz����'���'Q�'���'���'_r�'璙b�k^�	c2���kn�b�R��'���'���'�2�'U��'���!Ji�3U�-Ӄ�	*"=��
P�MƟ@������I�x�I��t������ğx��۞�B��ᆎ��T쐳m���	ӟt��ϟ��I���	ğ�����(��,QD�Tq9P$��?Ū�b����x�IП�����<���������I��@��a��U��1Wp�"D�Q�.���'���'���'r�'F��'�r`�;d�Ȩ�jfr�[6i#���'���'��'�b�'d��'�R�X�mJ�eS�䚽[{8�j�M� +�R�'4�'�B�'0r�'�:6��Od����d\��
�0܊�g��b�.8�'E�S�b>��v��5M�9��	.�0�q�.֌�$�P�O�tlZz��|Γ�?�q�O�j����ee�!궝�U�_��?��WӨ��۴���y>U��'������\���`W��%��O2��h� {��Y,-�(-��O�!0�y���Y�� 7�I@�';C��wI,�@�TI@ :ׯR��PHB��'�"1O.�Ş<�L���4�y��ƨ2�j0�#Yp˚����=�y�>O���Ɋ?�ў�ڟ���7m�0¡o��p��X�G�O2ʓ��/]�F�B*��'yB�;F���/�p��p�: ȝ��$Px}B�'�"6O��:�0D�T��\�L-���Jg&��'�"���-��H���$��˟L�A�'���g���k���ڤ���N��3Q���'���9O"�87�A3.�����@�D\գ0<O��oZ�k�X>���4�X`�Ɲ�AZ�R�x����0O\���O��j>�6M.?q�O�D��2���c�*8��&N�a��H>���?ͧ�?y���?����?!+�	g�,�A!m»1�2�c�������v�x�d�������O��l��?�	 '��e� �Bn>�L���G۪��瘉�M;����fpӆEo��v���O����Otm��� � �m��kr:�:����'& X8�F�&��S ��n�'�0q(Or4R�fϐy°9d'�������O��D�O@�d�O�i�<1G�iO|�[��'�81ѐNV.[̉yV�5Pw4�S7�'Cn7�"��8���\���Kشp����O)	01�b!H"`7"mk"S�M��'V%Bd�F mC�lA`�S;�Oٸ�n�������@�w< ��F˥����O\���O����O��D%�k���"�Dm�B���P�U����� ��.�M�@g�{���{�p�O�]���[�ZM�`s�`�zb��͟u�Ʉ�M#׺��$�!�Ƒ��F.��);L5�@��wGV�]0��ѯE)?��?�d�<���?I��?1`A�7wFt�P�BNl8a�T��?1����D֦]���П��I�h�O�>5��]<m�-SW�N�Z�I��O�Q�'z�7��IhO<�Oz��	P�EJ
�Xs�M�48
`�:��� �Z��i�"��|"� ��`'������	>���gI����)��ş,��۟����b>5�'{�6M)1�L���mN�R�Å� ��h"�	P"�'�V60����DNѦ�+3Mȸ~�n�J��$y1<0�e�E�Mǿix.	�a�i�I9~Gn�B�ן�˓Xلȥ����^�Aт�2�6�̓��$�O��D�O���O*��|�h�E����gL
�n%�@mD	h��vl��b��'��4�'��7=�Z�ئ��W>�s���_�@�+&�Ϧ���4㉧�O��u�t�i��d��27v00��c;�A��m-���:��'r�'	��ܟ��I��`���~4j��A[�`�|���ϟ`���0�'x�6��94,��O��DǾ'q�]نhї'
��aL$�x�C�ONXm��M3T�xҮ�A��=��,��_?�U�b�ƻ��$Y¹5k0xnڟ��!��	�����H��ԁk�<?{�������ҟ��Iޟ�G��'�8�4"���|k��z>P�R�'cf6�T�Ll~���O�dlZY�Ӽ�p�ةq�F��$ŕGI�cB�Y�<�iޔ6�Ҧ�q��զ��'���HW�Hrb���n�<�7e̎DNtM۲�������O����OZ�$�O��é"F�`f�B�U!7!�X�ʓ~l�� .	�2�'*��$�'>4x��L�3*�LR�-��6�D(���>Q��?aO>�|"�=j�j���k�7�q���	q\P�ܴ?<�	� �����O�O�˓4d��C��*��@�
�)k��r��?q���?a��|�*O�an/\��I�@NJC�i���F���>��I�M���(�>���?���uB���%��D�#��L�c]�DBE��MS�'�r�ˉH� �������� &Ԩ���s^,����@	'}"T�a:Ob��O:���O���O�?�P��B7$f���sp�.� �E�Kyb�'q�7mV�����O��m�\�	�9�h����,5(��=L�%���	ǟ���2loa~Zwo�gA���h���υX�������-{�d"���<���?q��?ᇃR�U��q �G/� ��W�_��?a���$�զ�� �\��՟̗O�vؘsl{˄(�"�E'��0��O��'���'�ɧ�)\%r�!�j�N���g�ӕj�% ѡAO�l6�KAy�O�p���B��01DM�%m,yu�MSjL���?����?��Ş��d������®u��T;`
2�IbC�?CI(�������ٴ��'Ed��M�����e�
�3g��7Ty�	�P�E�J��x�r0�|� �f����wG�?y�'��t���.��$���{3�:�'��Iʟ��������蟸��]��� "T� �ehŰbߨɊ6gA�:h6�%G��D�O���+�i�O�9lz�5۔��l��13b��$$o��"�Y��?�޴gGɧ�'N�Dm��4�y��¼t��d�;H;>�r��,�yGO�M�\��������O���X+]���sh�*r	CW�<<��d�O����O�ʓ~Û����9�R�'�i�^P�2pgJ�1fU�"����Ofh�'Tr�'e�'��u���^����0�K˖w]b���'	��O#��9�װi"p��j������	�b�䨐���-2����dM�}�Iٟ��I�����V�O�$�l7
�r�c�. 0��8�D��^Ab�f���8��O��$���?�;yK��ґiUpX�3���$;.����?���?��@���M��O�n��</��S�<�&	�#gn��-Ɲ)<�A'��'���'���'8��'�Z)�u�L2Eb�}�u�*�}��\��H޴'�ip)O��,�	�Oҵ��@Mm�D���?n�i#�	j}��'>B�|���c��, q�EM�`�h7	ԿV%T����i2��H�"�B�����$���'���{C��z1��B#N�H�y���i'r�'��O�I�Ms��+�?q'��8'�H�ei4]x�¥�$�?1'�i��O�\�'�B�'�Bd �@1��W<Z���@@���@��r"�i���!>- ןJ����.�i��xqqdþH��s�E���']��'�r�'���'\�ͱ�$̴M�-kd�Ӆ-E���O��D�O��l�%�؟Hq�4��k�|�;�.�Ok6:���H���xrNsӐ]lz>)҇�DҦE槕ņޱd�2[�)��N��|cT��aCf�OΓO����'*h��A {(�q���ü8�T���DƦPb��⟤��ԟt�O��� n�]���ac��1�*�k�O�@�'�(6M����SL<�O$ ۱�ž/��yr��;q�)� A�����٦uy/O�i�!�~b�|¯�b�.�{�du^ �ń�x����`�D&K�
���ڑ�Ձ)��͙  F'de����Ol�{�S�	쟐��k�$xl�MT��+�ɟ@��#?���o�p~ZwP��ןF�^N�x�&"p�l�e�6�����d�O����O���O|�d�|t.C3S���pG�#��Z6�Mc՛fN��R�'���I���+p�
,@&�	�ᬨ���J�����|$��ן���G���n��<	�"ܼa`< ti�90��8�����<��˃E�r��l��cy2�'���͇��	�1���dߪ	E��;���'r�'-�	>�M+pO2�?Y��?��_�.$��W, ��UR%@\��'�P��&dkӄ,&������%(�>�kcn�HND�t�5?��Ɲ*���V	�/����䌯�?9bMM�%W���u�&��d�W+�*�?���?���?���I�O�=#�M/&�4��<YE�|���O@<n��E�0��I؟|Q�4���yW���숀�6~� y�"�%�yB�'H��'U`��ƿi,�iݹx]e�&�У&�.@�V'G�]� ��u,P'�����O��D�O6�d�O~�Ċ5tU`{4�ŝs�Ν�AO?J��ʓ5E�6B̘b|R�'���t�'�4̐v�R&$Au��Y��@�>1���?�H>�'�?��Q"ha��d��Ȟ.����A�R � l�	���M�(I�'��'�I�
>�D�3��7N��4�Ҙq�����П��I�L�i>ݕ'�d7m��y�2��^�[`"�{a/�x��h�,,���$W����?� ^�������]�%;�9��͊SmzUI��΄SO�M�w�P�����?�r*D:MJr��XyB�O���B����@J9���b蔣�yB�' ��'��'(b�) 6-��M��J�w�V�2%�50�
�$�O����䦕�£|>���ܟ�'��r�@�X�|��4<�>1�U�Mly��'$��'����_ �&9OX��E�| ��`Pm� (#&V�Ct�e#�@?�O>,O���O��D�Ov�
���|@T� ���=a�љdD�O���<1d�i��<yQ�'2��'�哇u�zm�F*u~�����A�*�����x��$���|����~qz �okF5�&HH'N�JqѰ�� ��1���g~��Od��ɨO��'�R�uȏ,�lP�EDG�JU�'�b�'B���O剠�McPe�t���b@#OmT`ʕ.	&F���R���?���i��O*��'F�U������i�� 7��T��`�tU��~���I���+X����O���S�? @��S��+�ޥ����C�DҔ9O���?����?)��?����򉈕Zk��#��W�<�N@(Q��-��mڊ�����ɟ8�	S�ɟ����c�E�V���PH�L��""�"1r�i�O�4�O"��K>w��9O
��n/YktpAf��2�&��b7O��慷�?�J2�ĥ<ͧ�?��ƹ[����f��Yb)�6�N��?)���?	����d���e{&���������)0':)6P�@��� �>����]��M��	ڟP�����;~<	�ĉf��X�FO�j���?	7	��D���u��o~"�O����� _=�OB��rh@;4o�r��Z)+���'���'z����� ���k{Ҡ*��-�*̉ǋ	͟d)�4X�Fd���?��iZ�O�.�SE8}�NM�G� q�oJ�6��O��SЦ�`�̦]�'����w��?�*�������H�l��ȓ'i�3d��'��i>��Iß,�	��I�@i��'�!U��;����c�1�'=�6�v���On��/���Oȴ����76�f�L�=!�h�H��J}2Op�T�oڍ��S�'J�L#sI��1�P�c�ñоy���/�MóR�����[)(�D,�$�<q��KM����Q�9�Jy�2�޶�?����?���?ͧ�����	#O[��[ �"2R�uk���~� �k����ٴ��'�d�!?���l��lڡw.�\�"�F�
B�K��b�Ig	���'ov��Ej��?5�&���w{f ��\H8�%N�5z��'���'���'0��'y����� HN�)��ΙZb����6O ���ObTmZ����?����D�a�
 ���Q�sX�C���O�R%�'���~Ӟtn��?��v����)��?y� "01Sk�`e%�C],U�t����� &���'���'���'d�h�2K�r<�`f��Pct��G�'��W��@�4�8m9���?y����I�4��M��$�p\z��ϩ5��$�O�ʓ��&�kӴI�'j��?%��nY?vzN!�'��n�*Ҥ=>��6AT���(O�����~��|�G�R>�|��Z�|��4s4B�gT��'�R�'c��4Z���4}R`-�CS�v��GK�s�T�&˞�?9��?)O>�'��D��=��-
a�d��{���s����M�0�i���ŵi����O\�/�t�)�<����(�q ��sh�RG�X�<Q(O����O����OR��<�'w�k�+��7��7%�G'����d�
��w��O��d�Oғ���Đ��]�%*�.$��Pw��S��QI�'Y;�M㑷i5�O������د0�f6m{�Ta1T�R @��i���a)s�T�$E�e��oz�Gy��'rhS�E���"�c�������E�B�'"�'$剤�Ms5��1�?	���?��JN$DN�����d��ԩ��מ��'���d�v	hӖ=&�|iF�⸹kG�7=��;�"*?Q�f��ҕ�̦.�T$?����'+�x��C�R�[AAԝ8�nI1�._pp���D�	ڟx��D�O9BE�P���� �؀�H�1�NX�m��P��O$���禙�?�;M	��k��&�����/D�;W�`ΓF����r�b�o,d�<�o�z~R�߮i�D�S|T���g�.����'b��1��|2X�x�������꟬��͟l!�*�2��u��`�!GU�i v��\y���O��ɆQ�P�Ie�ܟ�B�\r�q��/�HD�3fN����O6m�^�)�IO� 4�`�GߘA��#A�>��F �{6d�B�0�;���O���O>	,O�Rr�	�a��Y�1e"+��d�0e�O����O\���O�I�<A��i��@�"�'V��p��Z�"=A���p�
,��'��7�:������O6m�ʦ�Bv��{N6hY�O��*��E�r��PW��oZB~BmJJ����'��'ֿ��%<9Ҕa���דL��M��*��<���?���?���?�N~���(�lH�@�]>�����d� O������?I�)�'A�����'W��|�X�8�����������D,b!���y·ijN6��2���|�P�ʟ�0$N�#Qzh@W.D�c`>$���Q�X�$x��'�B%�`�'EB�'�R�'خD*q \���Xa��::�J����'*�Z����4^���p��?����IX&���˗#�)b��DɈ4M�	�����ͦ	��4&������Ol�꣢��Q�5Q#JbT8��P�>.�=S��i��ʓ���n���$����G&��`�����Z������������	�b>��'�J7m��<��<Z��V����ˈZA>�!J�O2�d@ۦY�?�V� n�q�j��c*Q�u��
���#�P�4_��� %SțV����C'q��<��@!P�����D<��9�w���<1-O����O��d�O���O��'U��Q���=w��a �أJ*b�i�����'��'��OB�e��nB�,>2QjQ$\$(�X�Ӯq&1mZ��M[�x������'�66O�p"�E'k?�U0��Z0L4���6OPt"��~2�|2]�H�	՟�p!�+#��c��)�L8�0@ɟ��	ğd�	Vy�l����ª�O����O:�� �؀�ph��H����R�3�	��Č��a�ڴh��'�J�b�'͹vh8�ӎ�,\�M��O����G�8 kX6-Xc�S�q���O.Y*1��7N9�9 0�֩m9B���j�OR�$�OF���O�}��"���"�AQ93:l��u��L/x�k�+����<���'�7M�O\�O�.�Q#q�T�Sw�}b&ߌH����]"ٴCޛv�.C��F0O��䘷Hf�ɨ�π \9���1��e��^]���)���<q��?1��?����?u#��;�Iʷj�mQ�F%��$�ꦅ�L�����ɟ�&?��I(}Թ���4����*�W��`��O�$lZ�M��x�O����O��څ��J���'��$%��,wdx��ٴCR�	�/��T+��O6�O��K���/֫k&�	� �������Jo�����ʟ�SBy2fӼ,�C�O��Gƅ<|&�r�@�S"Ա���O�l�D��"��ʟ(����T�
�S�h,��_�tqB�)WIB�> <l�I~��>	������'ʿsB(P9�>$Z��_�Ei�쁣�H�<����?!��?	���?!��T�R�|���S���7v�Z#�v��'��#xӔX��0�6�$	ئ�$���G���h\��h��.#��Sp�����?I��|��iI��M�O�B�n��W�T�"��ަ7ް(�Gc��qm�Q��p)�O��|j��?���vJ(�H�h�o���(�CJ/7\����?.OP�m�g�b`�I�0��[�4!����D���~���L���FT}��'�"�|ʟఀCÓ�Vd|��ʉ2O���1�i4����h�~�����GT?yJ>i�o�x�,(��,*�t�1�ǣ�?a���?����?�|+O�)o�0�� 0�

�6�L��'kJ(�jT�ß�I5�Mc�B�>q��l ����D�B���[¤I6�N�9��?�q͊��M[�'M�	I4E���\y�J`21��b�w�9�U���y"V���	̟���՟���Пl�O4:�Õ�M:+'�Ւ0
ƶV[�$�!�u�J��ue�O@�D�Of��D�Dۦ��4�:q�ň�_|.���ց-Ȩ��	���'�b>���ܦ͓B����ZYbx[2��R���̓K[�1ȅe���'��'��'�L��'����S�{J�bp�'
��'�BU�0q۴1��M����?q�L#���M�>6Mz�zЅH�[�f�ȌbA�>���?aH>�	�c�J�V���,���@~2��?\`4���i:����x�'�R��=|X�E���H�A/��*a(T��B�'m2�'�����ĳ1O��,~�)w���d(00�����Z�4ad�����?�2�i��O󎍞�E����cGt%�#猵)
��O����O��դb���� ͵���J�*��qЬȢ2�u���_�x�'7�Iޟ��	�8�I� ��;�q`f��*s�0Ҕ�IRr�e�'�7�7AM����O.�D��L�'�?I�ˉ��uR��h\���L3��DA֦!R����$�|��'�2#�7Y�n��u�W�]��Y`��3"X@@����9*ΰtI��[4x�O��=��4K3e��q:��񦘓-��k���?1��?9�Fat��*O�tm��5�����C1$|����*܊\F+�r����l%��	Eyr+x�`��I��ӳ�9-V&! �ѼQ�Š�O�$ce*uoZ�<Y�����[���!SZ�L*O�����aɔgZ0�F��&�=q�ҵ�>O��d�O~�$�OZ�D�Oʒ����NY#r�rd��=��u�:)��k���O��d��Ap�'���������&����#���N`��I���)�S��$�O�AnZ��M;�'{����4�yR�'y$�
�N�4���Lj�r6�]�����^^��O��?��?��yH�#	�,{��thSW�[۠���_m0�-O�oZ"%�5��쟘�I�?��S���XįЍV�s��6q¤�ϟ��'��7��ϟ$�'���?y[%�U�J��Hy0��r���U�Xq)gmF6>�p��'��4\�� �|��ѝi<�8pg�ݏ&�`=@A.C ���'N��'����Z�<��4/N�z�χ��"����xEذ$-ܭ�?����&�ĂS}bcz�,!y�եd��ɠ](q�B7�FҦ���4#�PT��4��D���ƈ��O��I��ZD���*^��2$�8��ty"�'���'���''[>u:�
�8V���g�Ə�!�*¶�M��^��?���?����,p��N�hX��+.R��[%�ΣC $���O��O1��I)��t�$�	*m2� �tc�l�x ����/G���"MYFɆ�O�O���?��w��a[t�C�����ҷuNf���?����?�/O8�l���r��	�����3B� �A�܎"s\�K����5�?��P����֟�'�hf�V�kx\,C4CC�w����ք5?A���9[�,��4_R�O�����?y񅑰_��hv���H��ÈO��?���?���?�����O$a��
�%�dĐ�EZ�}�ȃ�d�O$(l�=Z�X�Iܟ���4���yGe�Z.�[b'�9u�h\�4�ԙ�y��'�r�'��P�i��i����TY��@�?;Dn	�h�!�#Bı�����Oz�$�O����O6�$��2	��b���xf$� "��˓�6�яgB�'���)�%@�sQ"@ /s�Ab����g�PM�'��'ɧ�O�V$c`��x�P��бA��ڐ��@��6 �<"f�r�$�I^�yyB�K�j8 �0��~>1���EjO��'@��'`�Op�Ƀ�M#�*N5�?�ǚ�u�p�n˸2�Z����H4�?ҽi%�O�a�'�b�'=2��*��}J2���mE��X ��7Z�)��i[�ɘf�hqq�ӟV����ȿm���(@L��0�
I�� �%��$�O��D�O����Of��2�U�&�9���Z��b坮bG���I؟\�	�M�� ��|��~7���|2�S>(�vtKgD��"d��v犭d�:O����O�	E<i��7�*?�)T�? &���j4>c�H����o@Icΐ��?�3F/��<ͧ�?���?�`H�rfk�1,R$ID�?I�����2֠�ry2�'��ӬNE��K�kED@,��*J82���V��IПL�����S�����S0�X����wd���
 �:EG@�<��X��O�) �?�¯,���+zh��bo��Y�!) r�d�O�D�O���I�<A�i����$��I4��+N
1�u�w���Lqb�'�6�&�	�����O|]b�k_�xkB�v�Txq��O�m�<x�pnG~o�n�!�z��է#R  �f�O�8ax����!��$�<���?���?��?Q*�����4,|L�YF.���C��ǦI�`�Oɟ��I��($?����M�;:Ϛ��4g�'����JF0G�>����?�Бx����\9U	�v?O^�
��Yjf�{�iS�8Y:0O�U!d�S;�?I��3�ĳ<ͧ�?��dɱ:L���ǖ"y]���X$�?���?�����$�ߦ���n����IӟD�"Q�Y���%�-`�t�j��e�	b�O��d�O~�OR0k.)�V`�V�!J�BY�?O��D�Xu���U(e�ƅ�'a�T��n?A���	8F�R�!%*���b� V�Y���?A���?9���h�|���	">ґ����EFDi$��;C���$�Ŧ]jd��x���&��s�2�eſϨx�CR�	�"黦�t���I۟$�I�3]�%lZ�<��O�"ճ�џ0(�o�k~HP1P*8zsĝG**�d�<���?���?����?�%��a����&g�=s�|@:w����Ц��#&�������D'?��	v��`�P�tټi�@��	s"^��'1��'$ɧ���'lҤP�/� �����4� ��A�ċIGT�0�i *˓'�LR�ʿ�p'� �'z�/EB�����U�u�9ah�?�?Q��?	��?ͧ����ɦ� p̟ߟ��f��@��1 �y ��cg�����S�i>��'\�'�r Ͽ_M�AC�τ�b��2х�:P�f�iZ�D�O*Ѓ" A���T[�X�S��e�/�5�h@�O�/'�'g~�\�	ߟ���۟,������uID+��zS�q��\�#7�?���?	��i�|�OZB�'��'�,�+��%&,���+>���H�|�']��'8��i��$�?=*SNZ�DRҌZ�o��U*[Sk�����O`�O�˓�?A���?!��]�ĕ�ǈ�L(����X�IO֜��?9.O��mڪ
�H��I���d�$���y�r�P1`�)���,�y��'3�	ʟ�	b�i>����}�p�B�b!pas���5�j!�GH@l�j�m�*��d�d[�'��'&�}����Ti�C[�NI����'l��'C��O�	��M�5�0c��4�c�Q�f�@��#e�>z�8���?a����|".O����D��(r���G�2��Ħ�+N�D�O\d@��b���	Ejqhȝ��TY�l����z� ?��x9��b�h�'��'�B�'l2�'�S81O`��Ǫ8s��Q�O��̜��4{�"��?a���'�?��Ӽ%��.���XԀֳr�2aش���?�����|z��?yn��MS�'5N�!v�gn��um��V5��'�P�q6F�Q?�O>	+O���O�rWNSXa�Lc��7�����On�d�O��d�<�w�iC�@
B�'���'\Z��Q�D�|�3a��pS@�:��'t�	�'4r�'��'k��ʤ)ګ��4
�E�d�'���ȸhlU���iPFʓ�
s뢟��I?50����&'B�`�#d$�	ԟ�����J�O�)�V�*- �n�V�S���2�t�BM0��O�����E�?�;O�^m��gA"z�H�3}�4��?!ݴ��&�]�����`���>J��ه@B�A1 JR�`m�#J~��Oj˓�?I���?���?y�8=*R�+&G�$
�F��$j���*O��mZ$�f4�	֟���E�S֟� b�п��XSN�3�l٧)�>��i���D$��Ɋ�c͒k1��:�!RqG0&<i��f[0�l�K�X���OZD�K>9,O�m�/�l�,t�S�Yh��w$�O��$�OH���O��<��i@�3��'t&��&���r��h��.D=/�f�#R�'�B7M4�����	Ȧ��ٴ;���"@,������?�|5R��H
l�l�c�iL�I"!J$(��O�@'?����+3�	xw��+
��H �B<��������ΟH�������a�'k
��!U�D�l~z��w��12 J4���?���^ś�ƌ���'x�6�7��Ɯ$q4P��7H��"W�Ď+rj�%��x�4/8���O��|�F�i����Ob�	'���:1��F�^w��p�JY�B�|=���n���Op��?1���?��&xBT�A-t�ա��/���A��?i-O2poi@>Y������W�D�� &4��1���Ju�HTC���D�V}Rkk���o���S��O�y�E���'}�"��f�[�𬛇�B�����<�'@��I|��!6^v)�-]�/�p�`*���\u�I���ޟ��)��Oy�kӂ 17�ɥ40��3�N�<��p�r�K"T��$�O��m�V�?y�I�$A��;&� tc��ο�J)SESꟘs�4C|�0H۴�����E ��z����SN3�ׅ�1V��ˀ�U2�D��qy2�'{2�'���'�2R>e���J��� @���YBI@� Ӈ�M{7埚��$�O�����dV���Pb ��%�u�"�	do��LM��	�HO<�|:���M󜧀 n�rv��*g���/�7,����8O���s�]��?y�"8���<ͧ�?��L�K[���9A.�L�sk��?a���?�����DYڦ����������<��CB�Y�|��ч��z���ـLc��j���l����d��c��F
~K���p�0?4F��'��@'NR3o�h� ��t� ��'CH=��H��0�8 �l���'�"�'BB�' �>�	�� ��3�Y4e�T��AkڧA�N<�I��MK&�ۊ�?���r��4�8�y��(H$�pb�@��GǮ�ن0O��$�O�qo�A�l�k~��۷c��x��*^~��ad�9��`�S�W�z0�|rV�����x��ߟ ��ٟ�r��
-�1�]![��t�&��xyr�~���a�ǣ<�����'�?�t"�]��X�5ǎ;Ym~E[eaU"�ܟ�m�(��S�S
Rl�L�(_�V���c�=K�=�G � �z��$�D�O�M>�.O�yR�ٱ8 � M�3hY����O���O ���O�ɼ<�F�i���CR�'w؍���0SB(���[�V��$pa�'�&6�(����$�O,�ď��ݳ�PF|��s�_.	��\�v"��t�n��<1�-��DG��� �'Y�$�w�Ђ�-޹qT�)��Ǝ�6h]��'���'U��'2^��'�?A鐪e3,@�.��6'8�Ce�=hk�Ta���?IQ�iJ$��G�'�b�'+�'���r3�A� PC�N�+Q"��gj�>i�"v�&ib�&�郧<�7o�D���,/�d8�A�5L��l�2i�NH��^ABH�D�	@y2�'+��'7�>2l���M�"��Dx4��$a�*���I��MCboZ��2���?��'�J��B(a~�T�U>C�������<���$����s�����|J�'3�ZB֋Ҹ���S"���U�������ɦQ���=��D�^0���m���O���b�O�|ߒو}{���O���O��$�O�I�OR���@�<q�iܡ�ua��y��g�i�vՀ^��' B�|�̦ٕ'�R7MքoX�9��B�l�x��ek=v��HlZ�M[&-F+�M#�'R�3&�X;�F,[3�I:�B0s��� ib�H7+�;�6�Iry"�'+��'��'U>��׉�}����R�O074P�@�ќ�M�֋��?����?��'��	�O@�4�}p�拓*��d��-Q��eVǦ�`����$�O�i쟤��C=q}86Mi��R���[;�=ؕL�!c}�i��.u�P�5�_�"G�D�Ey"�'��`��2��<�"��U��a: �GPN"�'rB�'`�	��MS�f���?���y�	Ρ{���!%�%>�� ��/���?�/O.`n�?��O���ە,�$����[",@�������O���!Bюc�~��`Ȳ<���J>������?�󭀼�P��� ��kĉۆ�?9��?1��?Q����Od �v&I������]�J� c�O<n-Pvp�	�Ljܴ���yW�ƐU�h�j���l���yRon�(m�M+%�!�M��O:�%��(������$}��c%Փ(*��;����9C�',�П\��П��ß��	�1��-����F ��!uiP�<��t�':~7�՞h���D�O���/�)�O�%ps�]�HX�B'����C}"�o���m���ŞY|��̍�uPɲ�+Ј2hL�˖�K�Mc6Z��ACǟ1,Y�D=��<ل�D�OJ(��)��:���Ѕ�?	���?!���?ͧ��D��]r��矈�2HU;
�CA΄�^��6L�ȟ���4��'L��!���z�@pm��� ���9�����QO4�ۂ����}��?y#���5>��Gy��OtWM���,�.n���S��*�y"�'j"�'/b�'�2�隤F����-_)0�҂��>h���?�V�i�r�H�Ob"vӼ�O�DbŹ6�
U�aD'iL)K`Ft�� �Mk��i{�D�D$R!�60O��H4 �t���I�z�Iq`�����	��~B�|�T���	���؟l�!k�rb�2�d@u�Ȓ�k���	iyBd�Pm�'#�OF���O`�'w+2����!zb�0ۡ
�4��m�'U���?I�4JZɧ*�'0��Ѱ�Q);�R�Z�oϦs���2��nPd��4Xc��?�x��OT�O��y�%R�Z��sǩ6$��,�O`���OF���O1� �XF�F��E
�8�W
%GU�b��Ո	�p�Y��'���~��p��O8��6_�}`f�BY��q �+u
~���O̐b��d�*�Ӻee���V�8H@i�78Z�"��hP"�bi�p�'O��'.B�'�r�'��S�{Onp�!9p,���<}5��)�4@;�`���?�����'�?���y���h|1Hg햌�`�cK\o�R�'�ɧ�O-,��i��:��H�K9�H(�Gw�󤙈΢���'q�'S�	ܟ���-\-d�	D�M��sbn�� �Y��ן��I��ȕ'f7�,J ���O>�$#k�*@����` ����C�_L���B�O����O��O~��C�! �|അ�J�� $���� o�&㲕n���'3M�����+��˾w)^�[�2Ym�������d�������dG���'�\Ta(_�iⰨ�R
׭2Vd)���'ǖ7MB7TB���O@�l�q�Ӽ��
�)Y'0����9M;DXQI��<���?��0��%��4����X)	�?����[�4S��:�d�5d^��(�mx�ty�'���'�R�'�"'_4;v����Q�aI5��"$�;�M+Al��?)��?M~:��a8Ș�t���-�r���>���S�l��4/�ҝx�����ހ 씨����H{j����^�_�a�F�[	]��ʓyan0���Oj�bH>�,O�Er�$h���c\6"���Bg��Oh���O��d�y�<Q��i;j�:��'arLb����
�k@|�!"��'�b�|2�'��I��p�	؟� 3��=�t��G�l��ș�$h�]l�<��$s"��&1�J.O��i��a��N�M���`����&م}�d�O��$�O����O6�=���Z�!�6FŖe�X%剞)�H�IӟH�I��MsP�J�|*���?	J>�P'�f2�i"$��O"��⭈����O>���OL�D�#vh�7�`�T��C�^�2&�D��I6g�|�Ē�D�,�~B�|R������Iğ�	DC�)U���k0`I2y�ן|�IPy��|�P@3g�O��$�O��'/X�i£$�ha1�K2�}͓�?�(O����O����I�O���B��yڬ� ��$.v��`�/�;,�yi�hoӺؕ'�����c?�I>��"ˁ���`��/	�p��&�͖�?��?���?�|*)On}lZ<},�3GOL�T��姅�;H�������I��<'����oyR�'����ӀPV����&bs��'��FO�W�3O��S�PTȪ4�On�Ɇ�X�wf��)G�p���`4�I^y"�'?r�'V��'�R>��H��|��(�	�q�,�悟.�M�����?���?�O~����?ͻ.B`Y��	>,��Ѭ�,R����?�+O�4�����O�uS��~Ӡ�I��v�᧒�~�l��0�ף(���	�*!�w�O��O˓�?)�.��I�W	��|mj�ˮx�bDY���?����?.O�nZ�i�4E�	���+(��d�R���\M�����&�@�	Sy�gj���	x}��'���D��3��$�T�L�Tz���'f�M�JĒ�;�,۩'��	�?ac��'���ɡz�Р[3"�hZ(�(N�@����������џ��Il��&.m��៸R�@0Wq��k����ž��$�E�0�ܴI(,�?q���?9L>a�Ӽ���ȮE�����mX�=".����Æ�?Yv�i��7�	Ȧ�y3#�覥��?���
v� l�1%���AE��-�ZX*��T�cI":A2�D�<����?����?)��?q���6��ݡ�	:e��$�� ��D���3D��`��ٟ̖O�剴_��xjάO�!��R��1�'�B�'���R�t�O�Ć�!y��0ӂ�Ɵb��yѫ��W��=І��0$�I�V�^%��'̐d%�0�'��AH��aw�S�Ɇ�e�Y�S�'��'���'�RS��#��B��T�	�K��`�+ѹ3<F���DY8*��	'��Ly�Lj�2��I�"æ�Jf1W
C�<�|%����:c��lZ�<����0�fL'A��H(Oz����. ��!*#6z|��`��f�P�I�3O��d�O"���O����O��?q�v�Ɲ,��R�ݦvmt�8E"�ן��	ϟ`��4 �@��'�?�$�i��'F�H���MC E�MBd��E+��ڦu���|R ҡ�M{�O�l��	�%8���R1ƃZ�Z�0�Ȅ[��L���c��O���?����?���Ar���A
}D�����!<�J����?�-O|o��9Ch�������_�da�}��Ƈݯ_�h�3'�����[z}2d�,�o�<��S�$�ݶ�ִ��/�2VB<��^�Q��M��'ZMR�U��1���WG�	�f�Z�	���.T�:aA�c��I̟��	ӟ��)��By���&��Ɗ�,z�"!��V���"h���}��ܟ ��4��'�t�%����[:8������F��Dy7�H�5[�7M���б��֦��'�����c�?yy�^�D�0v��%�0�^��r�"p��'|�{bM��K�HC�xt6������6ͅ�~���Of��>���M�;w8x�Ί*uM�řWC�]Y�d U�i>�7�S�)�S*s��1l��<�u\L���a�
ؑ�3n��<�jΘ���d)�䓁�<��� �zw�A���[0[x�H��~��*ڴTU6S��?��ej(�Rg�X�J�̰*�	G�L��[���>Qs�id7�Df�	�wje�2τ�%_��$슌+��	K%j��J�M���ti	T?���CQ(4�f��/h���y��G�@[
���mU8X ���a��x(�A6Oz�����A웶�ę���'{�6M0�i޹�6E�.2�,�ӂ�
<Zh�&.����	ަ��۴s�t���4����F-l+�'+��0p�C_�c
8�3�T.��!7�%�Ĵ<a���ZF�Hb��L(,�*0+�P�)w�Ɉ�Mk0a���?���?!��c�e���0�_��9sl����xA�F#|ӈi&����?9��( �U{��E��t�Ո������ۦ	�+OLl(�V?�~�|2[�챶�Dz��rP�H�!��܃��<�O��mڻ���	C�T�p��>a� #W�߂>l�T�I?�Mӏ¥�>AT�iK�6����R��B�nZ�YpA��q���%9Q��xl��<	�������?Ŕ'1���w�!%�<�V+qn��U#D�9�'���V6Yb/L+o6��4�R�y�r�'��"e��.����MKI>�Y�Cs����c>r�q��7Pr�'�~6�Q����ӐK�֜n�<q�Sp��p1mח5xԡ#R�b�)�τ�x�$G������/�	�qHdYSnK�r<��r�ǘ)�#<)�iP�	(��'��'b��I��A1��T�N6h���Ar��f��I��M#'�iR�O����� ��8�׾S��t@��4���P�̈́�w� ���IX�~���5��O�	L>��$٥G�n5q���	�|�v�{<�ӷi���W��M ��`�ъ���҆��{���'�7m:�������Q�A)�;[���q�d�74��Y�"�-�M+E�i��e��i���O����'M;�����<!2�[��P0�
�s��K� �<A)O����Ƽ ���띟9�~�[�oU;[��oZ�b����IM�'蛞w��UcC��C�,T ]����d����wӀ8&��������80�D7M{�D�%�X�& s�$)LD��D"v� ��a·GL��%�$�<y��?�"	�5�MAc�q��芝B�.���O<�$�O�ʓP��f��h��'���io�Qp�۴e�T{���2G��'���>y��iǸ7M�@�	$2y�M�V�ɿ6�N@"!�I+e��	ܟ�j���(Į�m�����r �'�2�H+C��8s���X��x�S��8}B�'���'+r�s޵�(՞A8B9�&��!�� ��FK��ݴD���B���?��i=ɧ��w�^=�C����t�� �e)�'E��ieN7�Z-6�-?	s� Ǽ�I����Qe ���ѵ˒;^}LyK>�-O����O<���OR�D�O��c�l�@�0T��/]��X�1m�<�r�i��fW�|��G�֟�a S��pv'~C�l+a,���D��q�ߴl'���OD�d�'j��c�C��9,�"ܫ2��F`��j�R�`�Ц�;7���X�I{y�F
9��E�(��e�GË�A#b�'Dr�'!�OS�I��M�M���?�Ʉ
Ybb��� "O�MA�(X��?Iq�i��'`�K�>!��?�Am~�`k\�?�ά 6l�>T���GcN8�M�O�PY����t���w[�XYf+E�c�^�ZRr�`9�'���'���'M��'��$=�s�2ʤ@P��&
�>xc��<����v�A���d�'�*6�%�D˼{��0�*T�F��
��`��'�B�4|K��O���V�i
���ym�!�hS�U�����C���i{ ��şZ�	Vy��'��'2M>tLYc�=��m+ Y�2�'��	=�M�2M	�?���?�-�vʀ*�>r�!��٨-a.	��?O$��BS}rh�6n$��S��+	�#�M �'��2�@�sB��+x�� 1b�B���ո�[������|�ɹ8��4��K"~�ʶ��kA ���������� �)�Syyjh��R��:��TB�� M\Mi�F�6ox�d�OJnj�	ڟ� �O�hm� OA����R#BH&��� ��ܴv�FGHv��&�������BL�i�<!���&m�2��BC66���p F��<�.O����OH�$�O����O\�'<��Z���:6��
�B��mR�i��Ūc�'r�'$�O�	�~���Z:%��$*�]�$�d���_$�?Q��V��Oru�a�i��؃2��@�$'(df�S�EܐvW��er�j��G_ƓO���|���o��QA�L#=j��۶�S�\`�����?���?�,O�XoںV#�%�I���	���<�M�	�ٚ �j�`r�4�	�����OF��WD�I)v�p�
$�_���І�E�b�*�����M�d��|"���On�"��f��d�b�+7l��Rڎ V����?��?���h���$֙X�t���ً0�x]Y�l�;�t�D��E3�����	�M��wY��#EWu���Yѩ�<V7�ʘ'���'�n6�0 7�2?�tC�
H��!?�^]�����ld~�����5��}�K>.O�i�O��d�O����O����G�X�1 ' X'tܪ�x���<i�i����f�'�r�'��O�"�̵ZS�\X��s ��Y�d��.���?�#����OZ�95�U�#~�*�Oިd�}�T-\�#IX�U~�ؓL��a�I�*�'��	�A��!ՎW1S*Z�c!T�	ҟ�������i>��'��6�H�"����H+L1�¦E,�@5�DC��[�J��A¦��?i�P�������h�4-��"a	�(G��Q16ʚ�
NskŢ�M��OP(�#��!������w�(cT�ޘ]a�� ��%m"����'$2�'��'�b�'E񟀥14X3v�0���D Bن��k�O����O��l�=�z�S�Kڴ�� n�9p˝A�`�k�c�p��5; �x��'`�Op���i��	g� )�i	�X��K`g)u:��;��L�S�R!�{�	Wy�O��'O��<Y�\e���Q�e�0U"bȍ�z���'��	0�M{æ׬�?�Ӛn�`�4��v�mH��\�f�(! ����n}"�'�R�<�?ə�.ӺV:M����*Qt4LR�@N�y�2u�����~��|B�a�O2�ZM>�d�![jT�ڶ
	-D�pM�Ѡ��?���?����?�|�,O��n�#������kr6us�NF�$J6�z�J؟��ɝ�M��b͵<q�4l)���Viڡ-.(�4��|F�!���i�.7�C&��6$?�viС/$�)9�tKݐe��5H�l�A^T�GP��yb_�|�	۟x�	����Iӟ\�O���(��SV}c$���w0�M�w�}Ӝ��r�O��d�O*����$���]�,����R O;�yf�>o������$�L<�|B�+�Ms�'���V"�:���%H$j9ث�'�a�a�۟P���|B[��Sџ *���<s����Q�r�2TH�����ן��	ly"�gӌe��<���F����հ8�ΩquhA&~A��x�҅�>����?iM>� .Y����^�:���Č�%ʬ���x�A���G��n�����2����Bb����OF�w�xBa���l��ڟT�I���G�t�'�r4r�5%b��gB�0v �!�'�7M�,�����O��lZh�Ӽ��G�y�(�b�-b������<���?9�x�$
�4����p���C�?��&�I�~A(��	Y�'�ƓOL��?����?)���?	�E��@"á=�
��,ը}�k-Oz<oں%�D=�	Ꞔ�I_���H�!�F�����eL��M[���)؜��D�O���?��IS�ah�t ��ڀ9��8�UU�E�s�u�u�'������B�m���'��B�%+C��^ dx�lO)w���*TκF]���u�PIrq�K�T1���dNo)x�����?!�V���àr5�QU�I����,�r��sa�Ŋ5�9��/Y1�`��	� h�Rg�G	pX4��W�H\ A�'{2��sQ�]�-��,(BK�b���bp�K5��x��̅,�<؀.W20CV��ӯP��$�i�L�^�Zu���F/5�Y
���$8#��0�..]��a���V.@"�CI}�
�9cŃT�8!3��Z<	Gf	��C��=X �i޴,�R���"�����b�
=���d�{� ��?�M>I���?B/�~��]����@�(!�f<�wDO*��$�O
�$�OP˓x�X�XT?��	�{n��g<K��m
��f�I�ߴ�?�N>���?���Ӽ̸'!b,3��W�=$ � t���R�޴�?���򤎞l1F��O(r�'E��΄�z	�q#����"f�&oyO���O�U��!��^�Go]4Y�b��!I'_y�R�Ӧ��'�Z����{����O`�$���yק5��_�_��t�Ѡ�~��v��MC��?!Uj��?J>�����BJ�\,�vfچ�a�����M���Aқ��'b�'���$�>�(OP���:k��5�Ԝ+U���'���oZ�%�#<1���'��IX ޅa���f']P4�o�~��O����zB��'���ퟨ�V����s����おU�:T�>�େ6�䓡?����?QhFP�J�q���Ndt�u�V�%���'~��U�>q*O���.���ΐ��.�Pl��d�M>ܓ�W�t8�K�}�����	�l�'kn�q��RP�����>Di�Y�@�	$'�,����Of�O����O.�5e��i����D�b��:nY��O��d�O����<"��)3�)��4��1ǋ��!�1�Dl�4N$��V��	m�����	#b@z�&�*����jY
��%"U.�,X�'8R�'�rQ��B�"K��i�O(��v��?J�1�D��@h3�������A�	՟��	�\g^��=q�m��#��yÂbO�(���k�H���������'��X�6��~����?���-b��V�BL���S�^���"@�x��'b�K��O��*��@=�!�7k�ho�Jy7��7�O^��O���w}Zc��I{�a
54e�]��Q���ݴ�?���l'�e@�B����tf����փ;���r2�����806��O����O����F}�T�`{p��UM��,���
e���̩��4wP����2�I�O"��o^� ��̺}��`�ɦ��	埔�ɖ}��]8�O"��?��'��[�Cą>!ʀ�v�קq��;�}f��p��'b��'�n��*N@h�Q�ƿj�X]@t�6F��7��O���F��k�i>���Q����V����QS�����z7-�>�Ca���?�)O@��O��Ħ<Q�`X�j�2��NV}�4Z媄��x����x��'g��|�Z��/�����oP$0t�@ ��K�n����`y�'���'��	�]��$�O��C��K�[��۲�ԝWqnt:�O��d�O�O�˓���c((���F�I ������;�L��%U�H�	��@��oy�aW���v 
�#�!q���p'�O�
b<x�To��E�	[�Vy2.�'QR�~RpMS(�{d�͸U��	��������۟��'�:�0H*���O����^4q�M;��*�ȷtr��P�xBT��A����$?A�'n�r�U$�^�0�8�c����'�����B�'���'���[��ݡ{\�[��Ҧ�@�鞀_f�o�ǟ���
U�������O٢푖bĄ9��P��G�shBY�ݴ�� ��?��?�����?��ǁn�0	�b�
A��(I6��(�M����~����<E��[�[�јP��(ty����F�*7��O^���O��Zq��<�O�rHܜ:6I�?L���Ǚ6<�8`�p�ԥa�Ɲ�~����~"�x��PS$�W����Ӂ4�M��%4��)O���OQ�O��kѮ�*B�x�5M$���)Vy}�m��f b���O��D�O*��<)��-���)�b��y-�)3GꄸX߆U���xr�'��|b^���j��Q �t���?�ƌ���P7
��My"�'�2�'7��*	��Oz@�ycb��x�����C%&tQ �O����O.���<����	�O��ABNt�����al�(�fɄh�ҟh��Iy��!���0����	0<�m��3иI:q��5�Is�	{y�ON�~�1�Q�8�������#l]���	hyB�'����\>	�	۟��s����KO�J4���৞?DH�<��2���O��#�d�ExZw�^���aÌ/�5���d 6}��4���>�-o���)�O��)r~��ö6����/����/�!�M�.O�D�OT�'>-$?7� 0�KU��DĶ|�v�6%|`ӽi#܀��x�,���O��d��R'��Ӫ:����`	�tPT�"��$K�4�?Q��?�K>��y��'�0�X�,@
-��a�1fK&"^  %Fw�>�d�O���R���&����$��s��0�3!��d��7A�0��oZП $�hٯ��d�O���O�0����K�ج�C���@�9�"��u�	)XSj��K<�'�?iI>�;$0�&��"�����LX\��'�L�Iz�ڟ$�'t�fH4R��Bn�E�ȫw+� 2`9*�P�L�	럄�?i��~�.�/�8cԈ�^xQ*`�=�M{bZc��?�(O�����Q���G�TH;ŮT&�`�G-��HJ�6M�O���5�	����ɰo�0��/nӒ����%{���V� ��v��\�0���@�Idybk�Z6��'�?���©0� �"7�.99�NE��'W�ɟ,�I����o3J�'��Q���33d��G��lhaBٴ�?�����$�l�xa�O�2�'��Dd[�C�"�"�+/Hn�↯0:��?I���?�B*��<)O>��O�@P��	�9��b�i��j�bڴ��$"y��ilZ�t�I���������� � �ӏ9ь���� "� ��D�i"�'X�ә'�2�'��iɛ?240el��Y�L]k�k��6�fɂq�7M�OJ�D�OL�)�q}�Z����3��@�5��X��%M��M3抜�<�����d9��֟,:ç��B0d�2'�(H�q���*�M����?��L��RX�d�'M�OL��%�R�}�H󥛐��y�7�i��_��
�Kx��?q���?�%KL�T��t��l� !D�r���~���'��-��>1)O��$�<9���,�)ǂ[*5X)z6��A64��Ox�"�;O���O��$�Od�į<q�L�`��<*7�ɮD�jHf惫� ʑY��'p�R� �	���IVD��t�@H2穆�{���De�����<�	ԟP��ybb ;��瓬W��`*&����YcE]�^�t7m�<�����D�O��d�O�0�G>O��Y��O�+o�$Ӏ@8v콂wO�����՟t���l�'���I�c�~���K��P��H��u��/g�|1H榝��Myr�'�b�',f�h�'o��'���V��K� ��*˩?���dӪ�d�OP˓< �|k�]?��	��$�Sn� ,�Ҋ b"n��w�³wKL ��O����O�����UV��OZ�D�O���;V�*`���	�=
�I�!Z$+��7�<��Pқ6�'���'d��%�>��0��)��N7O��)�#��1�\o�����	�q^�Iҟ�����}j�R��dЧ Dp��|�  ����D%�M����?����b3P�|�'�����PH�&�S�BG
_;��C*wӪ��>OH�D�O���/�S��8�j�wOteyd�ܕ,<�1X%���Ms���?��^�X��'[�d�'��O�Y`hҟZz�@�p��!��ѡ5�i�'�)r�����OB���O��h�^���Zg)O16�����T�	���H�.2�O^˓�?�,O\���&�9�l�,t��p1ĪV-G]���_�1�d� �'^��'��X��b�a����4Ş*V�r�w�H����D}"Z���	gy2�'@z^h�H��t������G���1�M��Bsd\̓�?i���?q���?�*Or�u��|z�`8f�a{��#G�6���%�٦��')�P���I����I�?٬�I;88�U!#HG�Al|�!1�;}
�1ҪO&���O����<I��B'���P!��AO���w�[Wj(z���M����d�Or��O\4Ð>O�'e��`fM�$�8QC� Hg�$�ݴ�?q����d��=�O�B�'���� :4��J 
Ld�h0ЋC�$��?���?����<M>i�O::10��>"�D���C�4��۴��d��(�l�m���������������,j�nǄ����7l�%]b�h
��iL��'�*5��'���'���I��6�a��gS�.��иV�Əy��v����6��O��D�On�i�^}r]�X鐉J5��$�W�G L��"���M��b��<Y����:��ߟ0��T�L �����:G� ,�K*�M����?I��}ݼ��R[�ܔ'�2�O�	26J�8��Ҳ�k(�y�i�W���w�i��?��?96�յ	n,�+AN�S[V��î̿L�&�'������>�,O����<���[P�ت=`�\*���a٢Fڈl�6��O�(r49O����O����O��D�<y7da$8y�'l�*�H��0!�k�؄�q���OV�O>���O���U�r+8���<��kE/�	OR��<a���?i����$�U���'%��	r���4Z��!��U�('���	A�	ϟ��	~��:��E�Ny� �aq�$6��O����O��<)�!^ D/�O8U��C�<�(���A�AaT�zcwӺ���<��?��L�<�Γ��L�JQ�&�ˡN�4S�d-a��6m�O����<�t�&1��OI2�O�J�C��]1�Z�X�@�?�2���`"�d�O@����5���?E2DA'�r�ɓiJ�m��{q�aӀ�Z�<��5�i���?���%��	t?��)F���M�؂Df>/��7��OJ�$߱'���D=��)�S/��Q�4�U�uᢝ��m�!O��7���	�v�n���l�	���0�ē�?)�m�Q���ф����8%��6C�:�y��|"���O>]*B\�v���h�>$ �@%�Ԧ���ޟt�	�%��a��}�'	�DO6'��4hA"��Qd�R?5I���|�b�8ak����$�OB���|�? J�����E,��L�9]��`S6�i���F0:��O,�D�O�˓�?�1j̭N�%�����;{�L�'��S�|�'r�'��	L���#�惘'"J)���=�`H�4K�����?������?��j�j��S�ۇ.�����^�kcre2VE�<�*O����O��$�<�ci&��4nIp��	R��I�ã��T���	X��	12Tf���A80ȡצ]^\��S�� �U�h�'���'YBV�4a��/��'rN�ӳ�&��rk�^�T�[Ҷiҕ|��'��Ж=A�>���/0h�(;!!�7ɜ!�T�ݦ���ٟ��'���Ө7�I�O0���/,��<�T+K�su�#��V��Ly%�8��ퟀ���V؟x%���'Gv*U�W���,�#�h����meyҎ�E6�A_���'-��!?�E(E5d����E�
8l39x�*ڦ��	��h8$�Ma����OL	���P{T,��/��uQ�a��4v@x2U�i���'ZB�ON�O��f&�bCM\�&��)�䋔�x�4�lZg��5��}�)�'�?q�kH.8�ʌ���::$�mN���'b�'����#�4���'N �7�~�l8c�`ŋq��4�?y*O�-)�*X�S�L�	u?����(o�TP�O�'\2�� ��O��D�:S��˓��i�O��O؍�&&��V���eS�t��T}�)e�Veq�Od���O���<Ib�I�q�8U��_�`�.A1C,SA\����x�'���|�'��f��+��ݱ��C0`$p�ĸv��쪉y��'���'{�I�؍��O��:�g����i7A���J�Of�$�O��Od��O���aR�����<�~�!'��k�(���-�>Y���?A�����̉�'>�C�/�,\J͛K
?/���J%B��Mk����?a��t4���>1`����U�Jʐ�+0���d7��O��d�O$�Ĕ	x�,���O���"d�B�#?�I��8�Є��a.Oǉ'q"�'���H�X�������2"�0�2�Xh`�p!�P"b�VV��がE��M����?���� P�֘�y.P`!&@ _N�� �B?*�pO�;w�%�I�?��O�0��͗�+t�uņ�Kߜ���p��Vȟ�������?͔'���&m��u(��&.��<�q��Q���ܴA� 3*�e�S�O.����S;N����#gX����
i[07��O����O$��&m�f�ߟH����9�+�	����k���F�����'���Y�y��'�R�''`���gK�Z Ty��,zA��qgL{���E�06n,$���	�\�	PyZc�ڀ��B�I�"����@�i��h[�O�̳��D�OX�d�O �0���.M|�Z&(� b�Z�	��/K�	py�'�I��I���b�`�=��8�Nӄ�:0h��FMX�ϟD�I͟,�����'���ȩ����O?M&��QR�$�x͒Ł%�M�/O���<���?��Y��8Γx���
��״�8�ᄅ�/,�lL��i@B�'���'y�I�Yr��٪�����֥ ��� ��CuELz��!���i�"Q����ퟀ�	� w@�	|��ǤGyK���ML��)�ȍ2C����':�Y���E���I�O�����>��"J�T+dpW�i*t(򐌘|}2�'!��'�8���'02R���v$�˖$��Ca�D��e��}H�ho�DyB��/��6��O0��O�ɇ^}Zw����IH l��!
M�9N�%	ٴ�?��r���?����?)����ŊD�����C�6�B8�b ���M�Bɗ$���'��'q��>q(O $�WkS�I�4�c�eب��Φy�cg��&�`����m1��Ǝ�~�6s��C�'�I3��iR�'/rk��i8�����O�	� ;Δ�`
ߧqW��ej��?��6m�ON���O��Ӧ3O�S۟D�I��83 ɣd�p=#��ר���seL!�Ms��wy���bS�8�'��T�<�i�ո��I�ogܭA�㈘�Xhc��>�����<!��y�(v��j"�"��	F'`����5Kp���FٖC�I&J��q �& �6u�ьd��>g�� k�p�*���t�0QG�"@��Uj!�ĨuZ|����x�~u)t�Y� \:fG�7\�hi�oT�Hö����ϾY̨���L������V�0n��i���j�D1�¬@	i�� �
�lH�@�7�� �"�p�I	'R���������M���[�`�ÖLŋZ%z���}����3gɻh��j���;$>����<�I�� :��W�N�z� aI8[�n!a۟@�`/۞���awM� \]Vy���X��Xjc�V��mht���	���?q�d�,SbV��E+@VH�e�-ʓ\u���	��`�*E[%L��D�s ȪY~�,�vOZ�<���}HAP %?�*%�ٟ.�
x��ɗ�ē5���H�
��D� ��e<<\͓g)�ܸ�P���	_�DǏ�H�"�'�h��M��ˑ-1s D���Sa }(5�Sk��YRa!L�v��T>��|�I�*,e �l�>E,�t8�FG#C� 4(0����Ub� C ���S��?��@�0��L����2����R�_
2q���?��O�O�'/�\q��,ږ-*풦u+h�'�t��𤜊7��ڥm[�����c�����!�:=P&��N�Ԍ 2�?b����O,��,N�\�����O����OҌ���?)�jMҕa����TF�;�チ�j�ѥ�'�4�����0$\~,�ҏ
XF{
� �	�ę8I��x�i�Nw�t9f�Ɵ��У��P�(��#�Sa��	�m�P0G'�<T~���̈́
7���I�;	����O<�=�(O���3�ȏf\t�c��=I$Th�"Of�
���X�6����ʹr]�'�Q���I�<	e��;�VjU�&~P5������ik�j֨y���'��'�Jx�G�'?b7�H���M	�iʚU� �T��gQ0'F��2U@B�m���JUF$<ONY�Ʀς}�d"7�0`A�#q�
Հ1��d��`<���7<O�=���' o�("Q<��d��#l;p(C��:O�ўG�N۹`�z9s�+��aD
5с����y�@�`U���*�b��)�2@ʁ�y�J�>/O�����ܦ��	�O��m�A��϶��%�� Z�<h24@+�R�'2�-K=ug���·�,�d0���)ۆ6|���F�+`��*0�=Q��:r��6P<�����1W�1���p�I�H��2�"��x�I�a��d*�'TdĤ�@�\�B��AJ0&�k� I��

�z`E�qVu�d%؋X`~̈́�I��ēw� 8�tÎ#6i2����O�n͓!p� R��iJ��'���lnf,�I�<ΧI�N�S&EF�L6��'E��N�L�hY"er��qO>�O1�b�,G�Z���C�x���I��2v2}���&oQ��O?��N�n��A�E�����E�'��[I��v��O b�"~�	!xz�]��A�9�5a"�SPvzB��:9e�����0;�h�����3/ڔ#<��)�7*����U@�5��$�ǯ���?Q��(�8�*d�R��?���?	��6,��O�A5)���AL��>��2�%ʜ߀�ZS�C3�`YꂊR<cH|��ߟFmEy2m^��Y�`���<vy`�R�,���G]&;� ��!���*�O���<Yl�[��\jC�ݦ'1D5C�(�?���ʥ�?Y���?�gy��'�剳C�8���Q��fq�� G�,C�	��L
]QLj`�4�N6>������8�S�d\��r�����M{�
Ÿj��XԄ>dؘ�C�'�?���?a��B�y*���?��O#(��?��J�73�,H3s.@�R &`�v�d8��C��<�d"��ժ��҅�9ކ�sR��y8�d;�N�O�䈑D��� V�M7'yt�)f��9{�!��N��K��ZYvt�(Y�j�Y�'MZ�r�\�2?*��B ��S�i�'x46�'�d¬L�l�'C�S> A�ܯv����#ͮV
��������Iٟl�	�[ߒ�9 ,R�O��"���es�.��̋,��č�7F	�xؙم�
j�TLu��(�ta�=���7D��E��lnL��ӡ��R���<!UH�����ݴ4ٛ�'��{d�|z7I�nBL��r�D�B����m�S��yҧ@	/�� ���ӳ}�U��蛦�0>�g�x��+D�q⛮kP����fњ�y�/�?���6�'Q�T>E+#�Zן`��Ɵ�a�cǪ&8A�֩�u������0Q�0k���i�S��D�,Q�N�����*r�T23`R'V(��k�XO7Vc�"~��+)8�k� �>Y���j,��� ���#�� �I՟��Ij��?�A/�#��Xra��Ng��+���<Q����>�TJ�BE`�R�[
q��rjUt�'��"=Yr���p�`�~��$3��I*0�� th<��Iݒg��"��5FH���Ί}�<a ��ʔ�C���
vg[��C�ɶw%8����~0p�0��<V��Ė�B�X(���[%�.5s$i �w�!�D;/\�EA�P�ov�Hh�� �!�D�P&܃��ҖA�p��f3}}!�&�����i@l��ɺ�dQ��!�$�_�ڹ1SسP���s�D*54!�$����}3ǂ�%~�Z@��ǱY8!��e���ǅ ��9i���8	P!�d��o���1LɜW�Έ�""JI!��`�����92y�'�˗�!��G~I�2ITO�}Q楃{�!��ҙv��@	���8*>JtbWG�1 �!�-Z~����ԕ ͦ�d�Y�!�$Ͻ.Y��b��6��kg��cz!�T�g�t�c��9θ���H�{�!�dӢ]n����S�(����1K� n�!�
�jʼ�r�S7�tЫ5l�!�� b���,��&0�So��{�*I`"O���������Kr���#&ƙ�w"O옢4mY�6:�9�f._�k}�u�"O>��PG��\zZ��Ń���+"O���ݕ+26��ĊG k�:�"O��BZ*C-8	�i���썈3"O�TY���
^�[��s��	�"O ���턠W0K��W���"OĠ��HJ"<p�1�	����"O�K3��7�`B��c�4�Z�"OP	�e�Z����I�W�0@1"OZ�Za�H�3�"�3CjG�|TiP"Ohȃ���=Dڤ-ҀI�+.��Uy�"ODdn����T��e[=��Q�P"O6�yG�FNR�u��'p�4uZ����J��M:s��O�OZ�X��N	WYt��a�ɳPD���'�j$�&�C��9�`�5���#S�G n�.� A�>}��\�0�A#
�f�8Ө�#Z<�G,D��ؐWӔ��!G͒`��-�O0�1�Mغz�Q0	ۓs�X�y�b��+e�e��ˎ*�����I[Ǡ��2i[�w��v̓$b�0H��ARnev+���y�'3N&4-+�$J���ꠢX���'D4��"Nb�\HF�d͛��BE�#d�B8nm)��D��yb�,�\��P�C9B�i ��+X�Q�"̔,	=*�'��>�I�A�hy�bȀxO@@�C��=jsȈ4%��a�T#v ���0�퉯;�J ���Q/6�;U�̟&HdC䉵�  �c���9����i�6�&C��A���`w����-�sH�1H&0C�u�	8��X1�̍Y�Q�	:�B�I6P��`��_Z0t�C�(d�B�	�g�����*��Q%��KJ��'\\#J/\O��2p��*|��(���&N64* �'� "���y9�"PQ����cɄ
bW l�ȓ!��H9�Ǣz��ѣ��<�uG}"Ό�A`F�dM��LW~E�`ڃwDa������?l��>E�tꑁ<����aĞ|���A)�#�~��>+�b��}��-
s�p UEǦ �=�
]m�ɤ$��ϓi��ء5�b���D͔�H�8�O����k��&Fl5EB�\����p#�y�2�[	�w��p�C���X��JJA����"Q/F�l�?!Q
*-u�6$��	�&7�d��I�L���I�x��L2��i� �$��UP!)��\Id�݇�	�FZ�#<E����~.(��F�ػa�T �O"�~�	6&��c��}���߫K�����_�J��4xA�G�<1N�YWJ�
0�N�+ȶ���Rj�d��_�M��Iy��\7�65(@ i�䁀o^@���Tm�%��2>܍p� \�u�"�� �y����"�z�ć2k��P&b���O88hª�Z�O�P�RT��{�!s6��N�̳�'��}���Y3d=ʕ��#�>>r��'Ɗ�Ѯ-�)ڧpvNy��F+2ЇՕz)P�ȓxr���w��_�\t��Q�@HB�O�����\a���
���]�WR�%�i!��L��p?yS��dغ����{�Pyv�=p����#-�	!}�Q��O� ����H[�e��Mj����$U/h��`F�TNC�F>��ʡ��B�I�k@9e4�*��<�WIQ��Re�YIx�9s�"O����/�y�dX7w�l1�$��8���Ȇtq�(�*=Y7���n�$�¤ՁMF)��	)��K��Y�C������XĀ@ᙨ0�p1���:��]�ȓ�ܵ���U��PU�R��'*�p�*����k	�[�O���B��b���iR�]� �0�'1�ղ"�b��p!^2D12@��Ok l��!M��$A+���g�S�? �2�D���9g߆w������'��5x�� �sݒM;F�Ѯ~�ЅЩ�FFz�9�%ɔ#$��3 M�<!�}NA�~;��9	��l��� Ƽ�P0�20-�">9#	°M�<�ȈX��Z��w0,D`ӘO�Z��!��R�\x�� ���'Ij��'VҐ�R��D��0GO�c�T��l�N�K��� ����4�[�Y�ґ���� a��~���_�d�ph�LM��S -�;��U�'E��
G���<Y�Q��bGE>RWl��0�A.f��Q���DDJ�hz8qr�+�_)���]U���B�]�6c^�j���mj������?����&iG�p���k⤑�S�I1�b�),Uа����f�:a��$G�֘��	;-���'�̍q���@��A�<<h(�O�Ofܜ�Ҁ ���s�j�(�^�x�T
ԿD����v��1S�`��`�����Q��r��q��:%���)
2�O�
�e#v9�u��D=� "$��p�@B5j�#g�=CЋ�!�M�*�h���q�焧GH�Ix�y� ��;j`�
w�^�c���g3D��8Ak.U2=��%�("lLA����S���S%'�3>r�#��$-� ��I8T�J��׷|"��3E_?��J�S#P����<28	:F�]؞�ВOG�4�'bQ�T�*\�O�!��I� !5ST �["��Ŧɛ%��IѤ��`�4�T��.�L�\Yw��+_.C���/8F��>1�޿Q�0�qQl�10��}�PY�<g7��z����[��L��(���
���oX�7hz���;�O����T�Pc4�Z�E1������>;��C1��$[K[?y���a�(0W1O�Qy�w�����I��;\dp �U=����'W��p�H%3�0�s.B y��a�r�{�T�2������u�j�%b<����ޙH����O�@Da�����)�� gs�����'Lp	r2O٬X�A@�кzEr�	veS�D0 )LX$z9�V�X�xA�mh� 0AE �@'ׁ��OQ�b�"(��;r)��t�$�� ቤ^�@4��՞�P��s�B
ii��ԟ�%b^�x}9� w�  	"O�������qp7��!z��݁Z�9S4�'7��@�/�1|���9�
H��Ȭ��rEA�9O��"O�2lֿHODШ�X%�\3� �nC�LġA�0�QJ߅qS�iƟ�(Od�����j`�k�>��"�'� \���5a2Z� BMéOP�"���~��q�'BT4��@	UB<��	>(�D!��^�NC�9��嗨�T"<�+�*<��F&��z��q���ϟ�Ӡ*�Ni4�PV�%����LQ�C�z�Hi��[ e���+&���b)1�vj��%i��:�V������w��GK�:߸�kÂi��q
�'��Q%!٫"���[䎂�7��\�f�x?����7���A�w���D@+5�d<��e�@���@���_�a~���2�Z�{@�X�]Ӳfȁ~���F�Ys$ r��U��	����I�f����J�FK�/��O��E��%�t���Dl)���(Ƥ�w��-X5f��'b�q��A����aG����"�3�D�*r���᪐�Mc|� C@�2��Ā�[.
��0�W>J�U)'��(v��K1��'�f��NǦ{K���-��X�Q�'_����]>u���E�ď36(���m�~?)�o�Z�~��E��o:O\�{�v�ju�=?Qb��5��Z�%���ʨ��d�S8�x(�BӳEϔYxu�/e�]
���֙H��߬7�Э�V�ͅ ���`�o�� ���:�>�j5�S�&�N48���<�P|��e�`�'����b��x�:�jt�&/����t�Də8������,h0~�IѠ�5���CI<Q�@�1b���'������Ir�AB&+�>r[@)��Ex���#3
$2��!��"�MG��w���T�ö4.C�gi�ti�'�V	����Gkv�B�e��%���X�b�0�M��`�����C1]K�i�W�'B*�5I�N	���[ĬQ�	�-o�`��/eƭx �ӑ}��y�Р�D*bI��ɣC8(<��C����>�@c��20:���,�![؁�挒^�'U�P�׉�:�pU�EHSʦ�QU>a�r���Z�۵lA�4�-�e�.D��i�'�Nxԃ�d�}��a�M�F�ҁ�d�V��̓c�=k�#~�}H���#MJׂ���3Ph �ȓ2�����	O� n\�څ M� 2�8kc�ތn��KfΔ�Y ��J�C��|F|���/|��1�[�K꼵kh�	�0>Q�M�\��w�CCx���l	-)���i�H�e��p�,|�����X 6������>^t*b���3�O��3pi��D��M�E�B5Zu���O;�% cOG6�2풱�GN��@��T�p�!�ď�%�2��J��K��h�&ē0�YY!R���h1Ě�r`R��O�"��L|z�'�B\�T ӂy��p��@_��	�"O4��2)�=.�J���aŚV� `�!FҸjb�ᖡD�yF�)u�j4���-R��=��k��JUr��5�_
N����Z����'%gJ�"�x�5C;� � :ՠ@�`~��r2nWS�.���WT��u�����I�c�Ĭ�PH�!���@CJ��ݨ㞠#!DC�.T
<�f̆F*� nX�V�Y'1�� ����3?�R���Nϖ_\��h�'Q�|���nNؠ�uB�!t��ڗ8Wΐ�f�(Z/��Q�gN���w�I��^?���j���#��EL��ADQ
�y��P`E���Vh��at��=�7��0J,h���
�<��P�27���1O����X_�24�Rʎ6m�,s�'Z�lZ6�v5 $X�(+F�Rى��?Zg��N����"$�'���@U憵o�.����ԯs���9��ğ�����vMՇU�İ&>�0D��0΄#���0���K&'D����	W+a�*(�W杬_��I���!D�P�����U� ��`d�6U�:|���>D����V�P�x!"A�&�}3e�(D��i�	,s]P��'l���'D�\@妏�-`Taqn����L%D��0Q���u��0�gN���)�Q%D�L颉���0�Y��,1>��!D�l��ߪH��h�Sg '#�i�U�;D�<���7ejh�c��-!����>D��K0G��p�T�h��T��j}��<D�<�凑p�l�BE'c�`q��g<D�D�d�/r|����G6	����:D��JCF��yЈUZ�D��y����@�-D�Ћ�iޚw��!� %�D���-D�����R�yH��I )�##��2�+D�X��O�EB��BL�z
 �y��*D�00���&�F5�r)�,G��|���4D���GQK��| ���bu�<�
2D�d��(X(^I!�!ؤe�ty3
;D�h��	3
(bU���s�,UqcM:D�L��*C�Bh!��]�,�'9D�̪�.<r���ZR���E1D�Dh�j�`�n*5'��T���#E(5D���C�(����������B�3D����Ӿy�Ӂ�8h�����/D�<B�_�A/T�A)�	A��T�A�?D��c��A�D$|)�B��q7L��a<D��	u�ߕ$�A[�'�T�V��f�/D��2r��:���� d+f��`�*D� @KL7E�
�c KYH̘t�$D�X	�֡Qö�p2K�2.dCo'D� )��<0���r"�|d΍ m$D�$x@@A�vJP��t�Vb�P�"D�D�C���L��eI�y_t�ѣ�4D���u�I���c�S�A�:L�t/1D�<�ѩ�3W��(�d��3�X�[f,D���¤I�8Q�f�Z-s8��H$D�x��q��I��*�;&�Z r�"D����.�8Aö	��gِ8Qj۳�.D���6G�D�@U�3e�F���q:D���a�� J*�LF��d���2D�dA�/���p���52��"%0D�,��<W8�H5��/4�� �E-D�<p��\��*գ�l)B��ȃD6D���&�1mv|i�\�h�.3D�<��#L94��u��.��4L����6D������1��PgX{��ó�3D��;�G�j���K��m��a��%D�$qch�����(�^�X�S�,%D���
�[�N)"��0(2�q�D5D� Y��%x�J0+��=4��2�2D��H�@��/i�]A�O:/����1k/D�H�7+B-ɼp��ꎾ����,D��yDL�'>���Z3.�Z�Ҡ�W�<D�� p%BTOЯ(zPۧρ�xhL��u"O�����ٵ+r�XZ壋Q)2��"O�h�0H��	z	����4����"O�<+��ɘX�ha ׉Y,n�"O��!�R�7 ��S+V��`G"O��[$�9�V� C$^
u���@"O~�z�gܣd�\PGcM:È=36"OfcE�¦9��+�L����e"OV�R�&Qj�恨v�8;� �+�"O�U@��"`�P<(&A�s�Tm�"OB�P-��}� m�"�M%�����"O0L[�����-��H��Z���"O�=[�"S�%:�-��g���yn"O40����)!�tqQ�FT!oy�xa�"Oɸ i����R�F�>kL�@�"O��5�^)�DD���MM��!"O`}A�耸J,�}��#�����"O��PcXZ�y��ɗ��v�r�"O��UFSE���^2�p��"O���1��7P��t��:�Y�"O�1�$�aՕ�Vg)=��m�GʑZ�<)�ǐP	����-�H��`Y�<���M�ʘ��A��j��3GK}�<IvC3Oz�xӄ�H�.��`"�a z�<9�(Y�N%��_!�
��4�m�<1BcA-)�� B�D��p�8r�Ze��p=1�l�!��,���c�0��`�ބ�y�,��ܡ�*F�X�*P�G�V��yc9V_�E����U��5B�"��y��D�؍ C"�K�9������yoǃI)���/�*a�P̬T�蹅�;XB�҄��7����WhK&u ��ȓr�)��N�)�r��ǆ�+K�Op���߁7-�1f�.���P�JI!�d�4/��Hw G?6p�]`�$J!!��dl�����=��dB � !�$�&w'�-E2:�60���23�!��M��q�m�
W�5:��ʫ�!�$��afn�q�
=J�!���:i!�&� ���hL�0�!`'�_m�	�PfQ�"|��F��5:Q;P�d�VT�$�s�<�#��d��P�!�%b
�eHp��o�	��q��*E�]Rtn\� �����!U�xC�?U��"�/	:�"7JW C�pY�ȓq�Nq�7A�=6Mz��A�>�D]�ȓ�6���E�2�m��G�~�����
���Vg�\�@*�' �<�ȓW�jx���o`��"�+�ha�܆�?�01��UT��`iS�[�@$�ȓD���Ã�J�3z6�B�h�6k��I��y,p5��DC�%*��Fe�*�nB�z�ru�ʔ&}BDfఴA�)D�x�k]�;+D0i@[u@,I1'D�8�bl-��m��|[s(*D����d!_�,,j#T�@��,pgM%D��b��W��W�Сotxd�R�#D�L�!ŊM��K�БqXD�@
=D�(hCH�3��
D�\�� �n'D��PG�
$D�@ђ3�L�5�r�( !D��i��B��b%���L1r���0q�,D�pq�NƭJ=ةh&+��-a΀vB+D��*�O
��d�>,Ą��;D�(z�F��0����"V"�r k,D�p�V)�6Y8H�0���MԨ���=D�� h�q�!�(�J���ֽI�T1s"OT�A��8�������E��"OD�&�Y&3np ���6q�]�v"O����?�jX ��S� z�9[v"Or��`�4�)QѭS ��)���'~�0��I��[�a!j�Z!��V��(��F����ƒ9BP)�iѕFp���>�hX�
��i��}[P	߇j����2Ax%H�^�V�������ȓ=SB�{��#n�zE�������ȓ] vD�0�Q
G�n�!T�S1���ȓKR|��Qf�0l\��4��oր��v��#獋�`6�Z2坯KB8��<�	�k�r\Ȱm_;�t*��_���ȓCH���@*�%9�xW��b$�ч�9@���4閘E�e��ϓm �ȓk�֕�A�Z��83&G�q@�D��aƴ�����<mxz�q'ؐ:A�]��TP. �d,��t�$k���&�� �ȓ`��h�g��7��rE�T�N�∄�gNBR��8������Y@����f3N}��HӨod���^(kr~y��A^h��B2m�����"Ӡ�%�$D��Y5E��M�(���_i,��D�7D�XXe � w?8�_�w%��2bE7D��Ӈ�}ꂜ�ރ@>���'D���c��Z�� ��Y�p���C�	졳E!�)	���ZwK&W2ZB�ɥw\�����"Ͱ�zVJ��ZMB��O~6��`%�?�Z�H%.���C�I�Ba�����I�{MXd�Y�7I�C䉺��Spg�+X��Y	&�C�I4G*�i�D:�LL��0W�B䉪+��@��A�9�nD���4�C�	�B��5�)G�hl(�#;1��C�ɨm�F}�p��N �$� v �B�I9Q%+���G5 H�GNB�hB�	#-�LĊ�/HN��,B^LB�� ,��aQ�̍=]���s�	0ZB�	�"d�٤g�<
 (��Ö�y-!򄍕��ҏ�V�T����+!��-w�5yE+���BQQC+8!�$��0x�i
㌀���'+�V�!��ˬl�T�d,���c�A�!��IE2� iH�@j=
�Cūp�!�KՎ�z��A6p^�Sc�!�d½CY�P�p�d: A ĥ%�!�d��1Ӵd�&�Q2PQ���U�n�!�$M+��5аFɵA�H�Mϰ}!�B��ZB���MSɉw�!�d3Q��h��H�JW���%�]�!��l�qї)ܴFd=��$_�-�!��IZBRIچ�B>� �r��U!��Zo�%\�NǊ�9�L�H!򄍂�"���$#�&y� �9�!���e�Tl�#Ň 9lt����!�$/j4]�ī-B�X�o�) �!��#�����<-:�B�NG�L�!򤍓C" �7�	�w��%�'.1il!�$M�$u6i3��ҹ5���B~0!�DNFk<�����2;t��eȏy!��+lr�KwHR(�����K�%!�D�f6��m�HI Q!��X&!�W��FQ�¯X�xŊ ��o��u!�� ���c�=U��A���*��<YV"O��h�jQ�=�,�� �E�n��"O�c��(l��h ��ڧG��A�5"O*�K`���E	f�J���D�ޘ��"O�\s�hɆ/�����ԇ y����"O�tAƏ���@���zq,�pf"O>�@�#�&T��Y@'/�]f��B�"O�%��ӫb�(���S�ONh��#"Oa�e�K��� Y��!CA�P�*O�X�R�_�o���藻,�*
�'�^�h��0�N%��'�>Xn���'n4�;��C"_B���\";1EK�'
ɫ�X-�>=�4��(5f
p����d�/X׀ ��K��]��8���4A�!�Y0��0c�j�+�J`D��|�!�@'Pݮȹv�O8fR�qDN�!T!��׬!:
�"�N� �5����O�!��8B��[���*�,M[C�ղ,�!�Dϙfi���n��� �S Y<&�!򤍔yv�� L8Te�O !�^:�����hԘ!p��W� �!�]�,Ҭ����j*�+"��%�!���7z�Uэ����b5/@�k�!�DّE��}#�
��7��pi�'�EP!�$OV ����uhB�"���h>!�Dȫ16d�2+S�2�ZR��Z#7!�� &��e	�S����#$>@!��=�����B4,���гc��>!�؃@��.T�U@���B�4K!�D��EC���weR�&C��(A!	a�!��®L��,�ƌ�4UJA⠗e�!�d�?��B�|q��p��G*'!�dـ;�Ȍ�7�0I�	��ˁ�!�CX��RT�T\A���d���!�d0?E��c䑮X:�,,e��;�'�(Ā n� M�L�IX	�B���'�9�⋔�%�`�a��Qy���'2�ԻVgE,p��`�R\���	�'��)�"~�tU `i@	kV�Q@�'�84�SiA�F�@��h��Т�'���d��a����&�7Z�RM��'��9Ve����x�G˭M��`�'پm����+\�5�V�9Jk�X�'p���Ŏ/Yօ�.#���'�t��G_ �!�b恈���	�'��l�6a��t���(>��	�'�$�:P˗�0c���A!��{��q�'� ��7-իd��*� �n�<��'�f�a�CQ�Lg���^1jpj$��'$�9"1A˹E�ԡ� ɥn�{�'M|��� &�2�I��˜7�����'!��{�Gچz�
�@Vjє~A���
�'�pp n�]�i�Pc� aƚ�P�'\�E��j�-�
!:��Q�R����'�L�g�Y��j\��h�D�n�b�'=�˲-�j �V�.�h�� ��y�!�6���2��Ϝ��վ�y�
�.Yl0�{�cֶ�3P����y���?M�(�<¡��D&H!�:C�8��/J1��H��#K��!��Ø8�,<[S�ԋa �r�ZH�!�D
!UfQ(�.]�	���B� ڽ2!����D6xz���1gT(�F"O`=�Nж~M�y�l�D�X�"O� ���CG�?�9���R׌�r�"Oe��Y+},�T� �Q�C�¬� "O橫rb��\���#Q�����"O�|�$"pB�!P���شZ"OX` �B�pX����є1���*"O��jK�~��ܒ���r���C6"Ox���0B��Q���<�r]9�"O���눘g�$��*��g�F���"O��0�G��rD�	^�l�L��%"OR$���L�|��ԣ���9���#"O���կ����*7�r�"O�1f�� ��Ҡ�ȥ6� ��u"O���2�X�.2��e�؟Y�$�1�"O&M����"wd�����h�ȃ'"OZ��t��8� �PnF�XJ�"O��3�g��CG�	��ܲq"O� )�퉚���[E_T��a�"O���!@��E�|`�p��(6��{�"O>�h&Z�t:$�&��$-b|[�"O@��׊^��z�-�[�2��"O��Rq͐�3�*�c0lە�h���"O��Y�J�Mc֤r�+��|�D�7"OX��Ühp:$rV��*
�l��"O0�j�H�`9
u����%x|�"O�����(h��1c�J�^��e�q"O:�g������OMT� #"O�X���]6��[�g��u�*1�g"O"L+���|�%��aҧ,5Αɴ"O�T��dϼl� h�����Bl��G"O6l��A�T <x��A(!�s"O��cG���Ia��Y�� �A"O�� �Ĝ.'�*�jpI�2F��ؓ"Oެ��?T�4i2�K,H-����"Ohx
�N�Q������ 
 L\��"Or1Yנ����.%E�ȡ`"O��"%�R�rْ�F3u�N�1"O�\���� ~a����c��ho�@"5"O����oԍ_�0��7��>^�:�pC"O&]�'F�"61 D��8Ӡ��B"O��� �!�����׽o�����"O��G���nत�Ҫ�.��ẁ"O�Ӵ�> ��Ly2�JT�4u@"O,
f��t��5�"�M$	���ʓ"O�Qr���Y��� ��vv�M	e"O2��&��}?zUs��bk�y3�"O�����1��X�F۴?y)�4"OB120��L�$��$8{�)�"O����cNM�L�X�C�	c���"O�@Q Ț�=�(3	J�kl
� "O��
í�
s��x��{_���b*Od��W��	(�8 :r�˵Ux	�'y�`A�[�RYM�a�G�H?8Q��'���Fg��aR����G �q�'�e�!��G2̛� ?o����'.�iJ�m ��;&$Ae:��'�&L"�	�wP��1u���[In(z�'��1��8ĉ�1�R�Xo0U��'�@�S���=��Y�CR���5��'a���S�aw��BA&�����'�\x��W���ݸ��ר'�Ȅ@�'�؄`7)�1[H�xyPlԂ�xUq�'7bŢ"�ӫ9r��F�;/h$I�'���x��]9����E��0#>N8��'F�e���V;�\0��V
h/d!�
��� ��0��B� Ō<2�Y�K���C"O�	K`+�;g�J�*w�%`�8�H�"O���ҽ"��AY��-���@�"O$1�󤂐�l�de�([` 0�"O��[ƌ�e�xТ"_ �&(Ѕ"O��S�T��(���+P��8:E"Oh�C���D�Q�<�(P"O�YT	�>!D��)Sc�8yu�|�A"O~h�b݌lJ��"Z�m"-X!�$�"SX�(�ș;:�5@6�ɀ*Y!�DǛ�b��6D�/G�;5杅AA!���$+���9<*��FT&!�$����Xׂ�8p ��Y��!��7�X1�%	�N���L62!�dY8\'�{��'J����FÁP�!�&?b!�����=�6�0ł�?�!�D08�q�\����05DĹ�!�$Bf$�``��C�n�2ݴ	K�C�I���y�hY�>�2���{��C�ɡw�zd����;�T����>?3�C�ɓG0T��ѯ�?v8X���2K��C䉂*���_-G�b�mÅشC�<{`}X�%��Nz�I ��][�C�ɱUs�jK��v��|	pB�04u�B�	5<0��@hL�=����\�WU�B�I:m̬5P�T(J���X�Z�]w�C�	#"}�4d�-~YZ��&���Rr�B��&ru"��vK�
u�X���Ő+�B�I��|��g(�\R�@�,S@��B�ɭ��1��f�h�Bt��-ϱ"@�B�=)k��C0-��[�ʭ����-%u`C�	�|{� �@��i"���㑳5�LC�	(*�6Q
�+_,Z�~�0��s�<C�I8���Ȩ3|Y����MQpB�	&Bw&��p7.�D��@��*B�	��L��t �/�n��c1=$B��p�`L�6F�3�Vd�C"L$k&C�I�0�ё�cS�A)�p��+L?6C�Ɇg���F�#(-֕�w�Z<^��C�I�Jg�9�n��$H 兗2��B�I~΂pb��b�*�����}�8B䉋X��(�噓3&1���B�\#B�I<?��yiE��f?�@���;�C��
[��m���G�Q����ZXU*B�I)�8	Z�.]��LH2N�=R��C�I���9@@aɛ}B�԰u�S�aS C�I�W5n��0��<�D���*A(B�I�=�
����ż`�h�H�B�>P��C䉗"��q/81�8(�f�Q�B�I�3b��	T��U:hq��I's�C�ɟ"��U�%@۸VS.�3P�34|C�I&1+:�!�ľC5Z����K�JC�I�*��P�j�֔�� �&	'JC�	�Q1ꤊ�+�"��%�K�(2��=iÓ]��l2A�L�=��h+$�I�/�RP��j<�$\%10jI��È�/�4��OU�<�F�O�&x�%��,W�` �N�W�<��M�k�T,��L�
~:�	�M�R�<i�ny>���D�
�B]ѠbO�<�en? ފLCm�Q���Ru��M����Iw~�)Ҡv��kq�Z�!��t�s٤�?IN>�����Oe�ɷr'ph*�B͵��]x@(\�@���KW\c��,`( đ�t��Ԅ�p���ь�F'�lac�U��x��S�? ����ʡ�j陡��B�Ԡ�6"O����U�I�ਹ��5i�8q�"O�8# a6��e�Ԡ^0S�B�ӣ�'k1Ol(y�,�Mh`Ԃ$���q�2���'��}��'��q��܃��\�t�ջrҤ�9�O���JN��%�K�_��A�Ce�<BbO��Pb��!����-��zKRt	�"OZ�Vg�d���r����	��Z�"O�	�C�uP9*��Ɨ����"O�P�1���	��t��/F�P��T�'�1O�=�ǥE�r޼u��W�`"O2 (�νh�x$��ƅ�s�����'��d�E��m�'An謂�$JO��CB �$�L� `y'J(�w"OD@� V)��)E��
pDPru"O�����r�ʁ�cGT}_")KF"O���F�"l2����R�n�,-��'v��#��Wu؍�3�3$$&�A��$D�L��-���^�a�K�^���෋�<Qߓ�?�G�N#�m{6) �rӬ��3.���?��'���ī�p�)� N�1�� �'�؃��:-+��
�@Mp �'(���O�e� z���:#�&���'��$(�
�
s�� kp�]�|2(��'�شj c�?LܨP1�IA�B����V�OxD1���*2��!�� �X���'I��:����[��!\�����'����J4^v�do�Xv�i�'�@��%Q��l�.ZMA�
�'	R���b��u.��iQ�BA�i��'p��Ѐ߱��-�-�.;`���'�D�p"nY����0�E�!]���(�'���)4R��E3��c�����'� ��b�� �RA��Y��
[�'%"��_�zԙq�9��		�'��� Q�}b��V�H7 ���'q�Ё�o[�dHba��Pi!>��'՜�;�J�;T������'\b(Щ�'yZ���(��M�ڑ�to�]=�����>O�Q��̚K�91���K��%2�"O���!E��_,64�w���8�@��d4LO��c���2����Jbn"5C�"O)*�عs���!�Hڙ|d��"Oz�sgL(C_�a \�m�Rh�"Ox V��Cr��k�LA��h2R�$�O������M�0ؐo�q_RAqB�AK!�$Z-�H�yս:�a�E.ò[�!�$�,�|T�B'�)n+����ǳK^!�/	�<�ٱ��= ��x��̡DY!��XZِ!E	.Ġt�U�??!�D�C �$+��?�9z`C�%�!��X�9lRH���3~��b���q��O���2���S�N�����M=XK�'+�D[�=�.Р�"r�S�b<H�!��[1Y����w��^gBɑR��1�!���/4r��#⅗�bu.9�[�n�!�d�4H�������E�b�:"�H9p!�U	 �JIP���Zø����Yg!�$I��x0��ǆ~F&�F�e\!򄗟a���[&n޼*1� �L\.V��ڰ5w���ێ�8,��<8��;��y���&�Z��qEC6'�t�@P�8D��{���m�D�q��LP)��
5D��J�&~:��c+Y;+�i��%D�� �A�bJ`c.��K,8}��a�"O��t��!�$z�i��wXʴ�e"O:�ąB&* �k��I�h�a�p�|�'Q�Oq�$,�`ɡJ��ȳg�u���#"OL��ЃnLPYV�ÿ�J�ab"O^����S�����C%�p ��"O��@� �"�^�w��t"��d"O�؁�_�u�a�]�L� ���"O����W�A,������ ��RR"O.�:e�E uZX��E��Ł��|R�)J���B&�,#�RӠ��c�D��d(?�FLf��Dч��/�uZq��d�<�Pȇj�H(�֧M& �3��_�<ّ%ݢY,ެ"��Ȕu�$ifď_�<�S�hB�H˵o	�r�(/dC�	RdΜ�Ǎ�3'DY a�T��B�ɸ�M� K� ���s�ğ&M��ʓ�hOQ>���W�Y���˴@�V�4�[#*%���'\�6O>�!	�!~�RU�&ᄽJ&�|�R��'6"�IH�'�Tp*��9�@]`��A3B!���[��A8��@m���2��q�!�%qzH	��E"LN���#��;~xўȇ�ɨ<���A��`�����_E����-���Lj�Y�>fSZt`5B�h�T�?����I2=�V��B��Bf����=O�ў ���#d]a$Ў���+w��e�C䉦5�I����j>̭(bs��B�,V����M��Nq�f-(70^B�ɎPt\H��� y��Z��B�d1���<�|�Or�fI��,���Ʀ�y	��"O^�笜'B�(eۣ` ���	柔F��� 9�2�!� V
��a���?9/OT�O?ɡ��ǫ�D��c��		��%�3��\�<�`�NdhhX��j���+�T�<�w	�*c�5����"��%�N�<�t���`;�8P&�K�%uH(cbAL�<��(t4�g�  % �Y �L�<i�DZ�V�&�!���Zo|9�g�_�'�?Zt	Q�n�B� �^�l��m:D���D)3w��0�L;w-�Q>D�tY$(L0M��w��?k��*O��Ȑi��4�qN<{\��Ӓ"O|m�֨йk���3f����j���'LO�`��%��,��ʃn�+1���"OH���L�_��H�dN�A��lb2"O����54X�83�S�e����"O�!P�L??�,�A���vv)��"O�UaP���b��B��~	�t"O*���C�YՌ�ze���L!���"O�E@� ��d?�5'�R���r�D�O���$�t.�H�#@�l����`�'&!��� �])c�ʵx���1Aϧ	!�gGD��֊�$@+t�$�!�D�7(� �p�BK ^��:�ě��!�Q,ӒT�e�M5:�̨����>�!�$B�U|Ht��K[�i�U��BN�q!�ڤzht1��T�b��`T
�Z�!��?'��pI��TF�ГiD�-�!��"D�DX�g��,Q"(�	�0A~!�ć"�1���
E#u��?s!�$��6��� ��Tx�K�&ٙ0j!�䎲=`8b񫁺,�(eا�H�j!��7��tJ�L�FH+q%��-!��l��p���
<(
��E�ܘF)!�� ~��F�C�7������4#�DHb"OV�����*'K�a�����0����"O��n�B8���ea�f�@r��>D�L�K|-p���N�{�pc\!�$�rŬ0�g��xc:�C�FP�!��ȚF�6�Hs��3Z0���l�+�!�dH�+@lDH�#(Jfڸȴ�E�z�!��V4A�z����٩t<�l5 C�"�ў���a�<PS`�[�i�0U �E�_c�B�	�F�^Y���,{H買G 's��B�'B��5撺=�v1��K:r�B�Ɏ`�(VꙧTXF��&��cYB�%v��G'��RP)�$
�fL�B䉚_ !a�#��T����?b� �S�O��а�@�v,�T+���*p`��%�IZ��[̧��A�*)��8'I��LȔ�%o'D����*
�k���
�՟dP�P;��&D�d�.���*�*�x� �Js�%D��c�)�ʲ�w�Յx�!��6D��)�B��B�\�Ke��{��p�1D���+H�9�V�:QJ����B �"�	ԟ��IQ�fE�EL�;Hh��h�R���'�r�ӔT����:
2�B���_�bB�I�Pn5��իC�:u�0��C�	�>��HV���i�R�[�F� xۢC�9&X�,pBKЀ � �XU}�lC�I�p_�4�A!$$�Ѐ3�I���B�Ɍ	�a��O'z>tP��9>rB䉰t�3��Q~$ػFŽR�FB�I.^���`-H�lK��B7j�v��B�ɡ=���U��J�|��ɟ�%�B�	�`P��ٕ�H.<Q�_I:B�	 }H�������H��T��h��C�I�}����s�4�xȲq�MKtC�	�R����!�8N���p�W��B�I.X�fAJ0ɜ>܆!���X�0�=�çQ)�U�n ]��z1!�C�����a�R�"�0:~��b�U�vJ����t���i�#ϨQ��!�P�L�ք��@v�E�fŃ3:@�11��&�L��ȓ�$����>M��)�@Z�a��b�p�S̎�yu��!�)֘*�蹅�D�����fU ;bt1p �X7$�ER�'>�1��U9(0���ե��|�+<OD"<A')˜XT" �B�߁F������P�<W�R�>��5��FRX�pH�&�E�<�7�ٽ��t�U�r�hr��w�<�#��
�D1�M�G�`� !.�^�<���v�D�0�k�4�<B]s�<� ���jY@�#�9�bq���ox�xDxF�#X+<X�' �!*�oE��yRx����'&	�K�:��g���y� R��P21��!S28�F,�y��YŪs�R V��`���y"�ɓ��yHV&I�<�[1��%�y����A�28K�-�8		��c��yҩ��p�ꔡ���	��5;W"��y�g� ����х����PdЙ�y��}/\�+֪��j�ٰ�㟫�y���9xDz�ے����VPgLP-�y�a��0���V Mo��3�F�>�y2�Չh��,CA��H���*6����y�J�q�D1A&���,�3�L �y�M��k�V���|��Ed�=�C�)� H�c�ɣx9�m
��y�0"OP �g�;%�z� �l�,<���"O��� @��e,�M1�ȺHDPP�"O*��K�c�j�3����RK0�i�"O
h�d)�8�� #���H�I4"O�<I�
�V�0��wN�#;3�x+�"O�Q:1	�4l�ةwH7h�@B�d�O���d�>@ql�*,��	j@�xfa��!Y!��V0� ��TJ�eM��AX�kM!�ߔ�E�Dqɜ��kU
�r	�'(ԨKq*�.�~S#bU�6jD���'�L�Rg&	�2nU0#/à.��
�'�d����R�Ȭ���I����s�'Z�q���k_p�Z�G�!�^Yˋ��,O���W�
t�Z�C$���b�Ѷ"Oν���N!���ʆ�Gֱ"O�⍉>)�bݨt�A<e��$��"O$�zDH�=T C��+8�T�"O,��f��(���˦H�<};#"O���'f���Y��^��d;�"O\i�&��A�V5���3ٔ��*O�e1v*��
��)H�A��k�"�	�'C�ോ��<t��b
�
Qnl2�'gB}��E�� �Ɲ����Mɬ�k�'ے����  #l<9F�R�C�`Ě�'��
6�=iґF�� :�� ��'n$���ރD��u(��}�ڤ��'.)(���X9i���-i�����'ӶH��e.b
��Z$eR�g�8i�'V|����ҡw&�`3%� 4��'���	K�?:H�8SG��~<�Z�'o��iG
�'X�D��a�=�4�J�'$x��dE0�]��@]@�4��'+4\Ӵ�M�NGDp���J|�T�a�'p�Y)q`]�/z�������qZ�0i
�'H�P��G�+80#�ܛYY��z���hO?�3��_�,ΞD���� ��%)!$�H�<�o�y-pͪr�S�T˞�X!��]�<��a�#r�N�[��
%4X��"VW�<��OT�H� U�a�D��@����j�<A$F�X��q��/P��C�
d�<���--Ԩ ꇠ܆V�I�sD_�<a&��a퀄����(2�zP�6C�W�<a!�_&8����%M�8���II�<qq�>S�eqF#^�<��P�<A ��Y`�aY�MO8V�`ǀJ�<����U��-�qHJ�<됵P�/�E�<��Y,`�6 �aa24��YC�<��e\
�!�F���vK0��#'�|�<���΋g!:��0�ͽ���!#Dv�'[?iasش0Þ9a$�[�%B<I�:D�h���^5���V��~<� B8D�@�t#�i�t�'�J����4D�����-�HQ���G�	�qk"2D�#�o��:|P��Ԏ��)��1u�1D��C���72gʜs�שdBn}�4D��Q��Fcy�d�;^C@�3����  "�KY�+)�L�p��0��U"O�9Z�o��c��2B�R�԰�"O~�p��6o)�G�&J���s�"O���lÜ#��3�&E�}m�Q�"O@��u�ب|

01.QX�r"O�L�4�ASNd]w�� Q�.��"ORt��b8}�R��B	o�piV�<G{��� ��Yl:;�|���C�
9�$"O�$�o�K��L+Y���qq"O��#��8c���/G2?�>��"O^m�v�כ^�*-�����V@G��y�P J�Պ�#	&;�9�T�y��ߙk�ԓ#!_�3�j��F�)�y"�D�y��� &���cs�J���<a���L	R���@D�7Yn�[�؄=�!�DL���r��j�z�W�ȅ	�!��K�py�}�v��;+��mހ
�!��ܳv�x�i��	A�TId�G�:�!��s8��co�'��f�
��!�j �9�h�#��ɺ&H	;����o����-��.�"���f��xkJ9{1+�Ό��if�v٣`e�7���!�i�:[�!��o����#�#h��K����!��+P/�� �Z�lPY@	w!�,?x:�2։��|�r@��AS>o!�˨z�L�ʔn��IrW�BG�!� :rł��5U�Bh�@·]�!��ƣLd��bjGs����Iŀ8��'��OF#<Qb(C$d��(�� �1I�p:�O�l�<�ץ�$KC�|�r� �f���� bl�<q@�
J�x��$�:A��t���j�<b@�t����:Q�����d�<A�GC�u^p��A�,J{4�2ӧL{�<�BO�?di~<��Ô�X���o�Q�<�b*�8{���#	�{�ވ�w�DQy2�'�"�'TF@:6��/B��%+����Z�'�����8��A�t�7}\��
�'F� ���� t��SL8|L�$�
�'+cǎ].��K��2��}�e�(D��Q��,"�4u�r�[8X�mR,:D�P��[�"�ʭ�u��cL�p�&D��`T�H���]&On-��/ړ�0|B�Ν�8�,��KѴz(4�R�or�<�J�O�u�ՍP2Ar !Q^p�<1֯����Ѧ��/hF鈔��l�<��E/k�D��;�ִ�F`�l�<y�
��)�PU�u�_y��T@a��}�<!�"*��ٳd��W3�t��w�<�O\�~�<p��ΎO��h���n�<9�]�i������^����'�h�<�į���$�5�Sh�r�(`��c�<!�.H�x�i� �7b	�L0��LK�<���[.C���7�ܵh@�Л��ZE�<	F�31�6�2��[�����m}����%zf���@�lh����âTX&����<�d��. l��gF�0Ⱦ|�'�a~"[��x} 2 ܉IA�e�2��
�y%_+cx�x%暠Fi�����y�ȓ�3)8I$*=|����W��y�)��
Kt)�!��3���΃��y�ϊH�L�w�3�Pp��G���y�CQ��A�.���~�ڧꔧ�y� � /�e�W/�%O��2�
���O4��Fx2G�} lx��<��-���y�`����iҍaC�U�cn)���1�S�O��Y�bϚ�Ӏd	7� ��0D�8��( p�X�q� �B�T��+-D�tҰm ")����#/f�x�#+D������72"`�k�+�6A��l{�A(D��pc�͗D����T�Q-��|i�'�I\��Ty��'�X,bB&P*,�(PTm&D�� �i`c��p!6�	9���*��|��)�< �@�ǌ�u"��R�L��H�B�	�9�]�6(�?b��թ��+[�C�I'�f,�3�Ƀq�,��gdT"~��D�O�c���Ç� ]����N���As®8D�P���	~'�������l3ri*<O:#<q���*]8��Bס1UB�3�{�<9�)P�!���u���BX^�	aBu��hO��Xc��Pp�������S#�}oֽ�ȓo�8$m�h�8@
S/愅ȓ����G�*/�$:D��nJ��	��@�<r@.}��I)s��G� �9q,�F�<QTjߕh�����müLڔl�$ĕG�<�#G�a�P�w�76'�`�hk�<Ar�U�+���
�B7cb
`"扙e�<1EG��C��;���+�%>�e��/����,O��]�]~�JY�ȓ�����k0hsX�ҧ��W����w̓F��(�@��d}|��QH���PɅ�_瀍{��ȴ ����Bƻ$�����"�<:D��D �� p�HjfdE{��O��0���F@ Z@�Y�c��XJ>��S^\e��&��dj�I�DވH��؄��� ���~���R�^V��0	�'��x�b�!������_�֜	�'x鱂&�>@�e��,j@D��'�0�T��g.��`O@.�=#��D3�8�Ï�.�b9I�fΒX4Hta"O`
�K�L`�k�^�R�=#q�|b�Ir̓hτ�³���6]9�JN��}��E` E�ÌR�(�K@
���&��ȓt��;��4�\q���^�v�6��YQ$���@P1j�����G$֢1��P�z��̅Iv�ٓ������F��S'�H �A��ꨙ��:>aHC�N�t��_�QZրWiM�rC�4�]�TL<c�Lkq�	y�B�	"8��D��ą;߈q�B��C�	�0�����m��#<��p�e�a�hC�I\��=ta�O�L�@ve@!�$��@~|�
�k�̝��ƶ] �}☟��@��n�=�f�L9*�*�[p/5D�h�)�G�R��	��P������4�$;�S�'V��Ċ��S n8�S%+�:��ȓ,�Ԍ�g��S*���@��E�ЅȓB5$؆ӧ~2�̃3�$'�(P��R\�H��
�|�����˜��m�ȓs��C���)a�e�P$��gܔ�cV_�	�ʸ�����r ���K�'��}�,C�N)�=�Őb�й��'��p�E!8\x���#&l����'ZJCE�I�>�9Uk�ev:��'1G���1D���G��?�Y��'��0J E�$k&�Թ�.X�~�h`�'E-�%�JLR�þHa٢ϓ�OT9�d�0g���5�1���"O6�`m�)ZP1U΍0^ʚ ��"Oڸ�W K#3ʎj�-�15�~��"O i8�BƧp3��r�z�X�""O*�F�ǱH���j�C=V����"O\(����->*��#8t��R"O�;
+�&��`�.n$-�"OȘ.��Y�V�vώ/�$y"a"On\���@-��l�/oh~1"O� �q���_F�Bن.��^H���"OL��.�8A���͝)�Z�h!"Oޱ�i 0#�H,(�U�a�����"O�ca��3�L����2�����"O�+�I66Ǿ�%�üP��\چ"O����(9�ҙW�Sa���a�"O�9�a�@8|B�1p�`\g���#�"O���"�փ*�� ��@��%@Y��y�JJ�Z���-�' e�DY��1�yb��)j@���1sH�U�r��hOl��Y,��=��ƒ�&�T����νD�!��+7��pҍK$ 5LMQ#��5;}!�d��.�l@#/S~b@1�m�Qv!�D����q�Z'�t�",�f]!�d�$YE��� ��<�\��Uʖ�f!!���-s�>aHǬ#��MQ竘-_�!�$�		~PY�fH+C�h���^�!��'L���Ȉ[����ׄE1c�!�$�5
Mڹb��Y/�^��n�7:�!�DR�40�E�ŋ#w�4Ҳ��m�!�d]< �J���#�F�s�K��Z�!��N�/���q�n���.Xȑ*Тij!�N�?9���q�3��cU!�#�>Q1��T$jTG4e6!�d�6j�n�����)^$�V��T&!��S�'�~1�t#�*)�Dh�V��!�!򄊯6v~���K�P�4�r�B��I}џ�E��	$6�k��C�L�"�3��J:�y�l�G����,I+5A�|Z���y�m�
dGv�Vo2c��#KJ��y��T'�򈓕AD"
N�"�ո��?!�'iF���ၔk�8yp�a�4){ �	�'C�YbQI@e@����ׂʸ��'��p�adԬ�&t��*'�����?���yR�>B
Ph5��+l`r��B��+�y�&9.�����m���Ba��yb��9��D%�^nBe�e�� �ybj�;�@uhU�XY\	[���y��T�-O䥋F��(P�N�)�`�"�yR� .	7(踣� ���Y�V�yr�[�m�2U�!"��*?��0
)�yr \7h�hCA��/��a1`D'�y�"���As�܌HݐX��l�)�y�R�|b��tJË+E�)@�݆�y�	��DHcLL0%8�X�n��yR�[;e���j̟1O�0�l�=�y2�'R�z�P�/���PB�*�y�g*1g �����!���#iJ!�ybGW� -���q#�2mg���BF�y��B&H��d] jɒQ0%ا�yB�R-�lh�
݀.v��W�L�yk1|��e���-�B�p�$�*�y�*�
r
�e6�4.��f�˜��=y+O��I�+p�d����=O�~��5��w�C�I�͚���Z8Y!�@`�Ô�g��C�I�2�A��$RcN���
R=Y=�C�I�(k��!��S�Z��ƈJ	4C�#hU끬Y�2�����		(��B䉈>�q��(,fS�I��3`�B�ɸ D^qTG�.� x��G5
'�?q/O��D.�d'+��ݠ�&�}�� ��Am�<a��*6n�kR"ǔ�J��e�<�ʍI�8(eȕ�P�@�*�K�d�<1B�5%��!����$s��� ÎW�<� �)�� ���`̆�lɶ(�"OP�  �^p�ԝ3�mH�&�VH�"OY����)/��Ř'm¨R�j<�4�'��	#81� )m^6H"�R�K�8WxB�	$%`����	6a��o�wԐ��T?�u3%�x��ݨ�CUe����B�L[�iΡJ�����BY+~f!��-�ʵ�ӯz����b�Mp��ȓ#�SƢ��s���zW`[�D��\�ȓ<����!�,j��˛W X%��� 1�G΄�c?��A�G}*�ȓl�`D�LX'Ma`$���N�Oߖi����<)� X{�m��GK�G+�Z��Z�<Y%�R')_p�:��9d���T�<�6�N�P,��@�Mt�y� �i�<��V5b�[go�6"��(�Z�<���I�'Y�-Ȗ��3���HD�nh<���=s���AcQ!��A��4�?��'w���!��X�����9�����'c��K�i�RY��M���,b�'[ HQOH&�$�˗iU	tے���'¤ذ�N�#�:����0^�h�a�'6�- ���ً5�
 @]��+�'F�m ��J;X%�#u�P�
x���	�'xp(8����`|Pp�d,:S�%�)O ����^d~�H�_��89B���� z!�ӣѾis�^��r}	�cD'�!�� �y\��L9{����$�?'�!�d�@1"z6��2}�q*5!3:r!�$�H�	�A)G��"�?D!�>�U[9<~�d��J�*>%!�$V
$ &����Ih񺦌#fO¸($K��nĘ�D�b��R"O܊eŧ(ZD��7	 P>�SF"O:)iG��!�T9�U�kG�� �"O.q�e����ȴ��%
,�\�"Ovqz �ޝ ���Iْ!�[d"O�(PY�:�P|�D�F��	"O^d�w��6x����)ߌd�T�&"O���G\-2��Y�3yzh�"Ojh%��K��' 	S2Iˆ"O����@A�!�\H��$ӷ49|Zv"O����%?�HstD@�:0��Ic"O��WHQ8u��D8��؜2-��32"O������	֋Ƨ'�,y4"O�|�P�ۂG�<��Q@�����"O����S(M�����*�W�j�;�"Op`!X	|K~%PD
5/���E"OD�Ё�YU�aŢТ$l��"O�u��	h��њC�
ڱY�"O���fd�#&���ʀ:�j1�s"OB��Hiz��H�J
�P��"Ob08ϖJ��� ��>J�1 �"O,X��K�^�"�X���4p�8zE"O<�J���$� ���"B)X�$(h�"O�P@ 
�>W��8��>-gjL�"O2p��T�UD愨��!����"O�qytiO�
�p�b否NNT��"O@tp1�D�\���5�D�U%���"O@9�u����,q�(�(�b�"OBEH_�t=2�Thy.��"O⹒T�̦P=������ Fs�x�R"OJ��w���.�J�RD�O1&VB�"O⁈s��L�z)����G�^���"O� �q�d��z��lX��.}��=K�"O�L�r�?>d���F�g��T�d"O�12���A��
a�	35�Y"O��0��� [Jp*��J�Kn�:d"O�Sbg�+ctaci:s\H�B�"O�뗎��T�*��G\�ѐr"Of� � H;�0؃1�ڦ2b���"OB�!��;:~�̃��]-i�v�[�"OV$�ů���6!�R�N�>-�"O���A�C�(���ȱ� �d2qB�"O&EЧ��)��@1�ڸ1xLD�0"OZ!���k6��Nn��"OY�r���ґ�$0Ii�ۂ"O*�Q�M9H<"��0��-~d��:$"OJ�iwaߢc2h<�!�3cR ���"On�H $J�Wp�)�\�j.�xP7"O���%ǭ?���c4�C�s6�d"O"4{�O,}�z���G*Y����"O�z`�VVy���0f[���#"OĨ�CH�c@0�!&�?1�nEX"O�|���!G�X��Ⱥ+T��*g"ON5���XS���ۅ!T��I$"O�͘��{R�І	@~  U"O��ӴB���Oɰl�B�0�"O���ɐ�c��x�.��F��ڠ"OJ:�H\�H��5�Q��2�̤��"O�8�w&��QF꭪s���5�""O������^k�����W/���4"OnT�3@X�m�1�R�w�C"O�=*�R\e��j���'lm@k"O����ʤ7�@q��mO�Na��j�"O�B��ДE�$���� :f���"O�*���k�X���J#ܫ�"O��`���~΀2A��,�'"O�IC
�W�@$#L�.�>i�2"OZ�! �+q��Ѡ%(W.#z��P�"O�9�/2���;���(�\�S"Or0�Q�� �SV��4X�`�S�"O�Y0��*��%ꗿkq`��"Oh9P	ؐ���r��~�ް��"O��87oU)K�\��$mזUMV�)�"OH-�A�ة;W(�y5mK�jF���q"O&��b.�-,hAPK�(1�p���"OFd��@8òpF˔)O�	C*O��`bB�,��%s2 J�hM��'U���b
������ص[X�p�'���YEꚽ!���g%�0�s�'{��Q���)C٠���%\�L�E��'�����V�m�&|��
O9t'�,��'-J2�E6j������ r/���'���Ƥ�m6�=K��Ǒ3*	�
�'^b��FkZ+N� �a���
�'��R�تJwFP�.K���Q�'{1� �L<I:YD�	,\0q�'ٔ�-	�ox��2���!��x��'.��b�]���h�o��:I��'fJ�;���7{�Hr4�t��I`�'qJ�saa��M�])gk�-]j�h��n�(@:�^�y�de�I�4)L�ȓvi��։�-s6M�w��)��E��u.t�`B��w�0�c��^ν��u-�d�tJ�C��M��_�JM�ȓE��ۣE��.�T���_��4l��Wr�P�%��:���ZP��RB�,��S�? �q�bd��Eʲ�a`��t&�԰c"Ol�ĩJ-~�! $ቿl���"Of���Ǟ-y�^I��_�<r��"O����/ڮ���vT�L�"O��hщ�,c�mk��4{@�q@r"O�-� F^'?>zt�G1SY
�""O����ɡvrD}�4��m;.��5"O�xs�lI)c���h��]	@Z��{�"O
�	Aֵ�0ȅ�[�@VB��"O]�
�����h��l��yW"O��R�^R� =��!ߓ6�*���"O�H��+2�zF�[���<�4"O.��m^�}��p�eN�/g��I�"Ohq���:�6eYf�*� ��3"O�d#v���~��((B�Dp�XS�"O0��(m�J%jd�P�@?��Hg"O�����X��eS�+D!Y(��"OXYٔA�;`]�oN
K�d=˦�?D��h��c��tZ dR
�%V;N!�$_�K$��S��x]�Ç.!��&e��H���1n_��� �6!�$��-������,~2��8��}�!�DE<0#��+6GY9����^�!��`Fi!��������T�vB�m7��3���X��9(�b��L�\B�		Z�Ţ��ʑQt[P�
��&B䉀>0��gŉ�Fqa��rʦB�?��)�*�'�Τ���AX	�B��(A�5˳���h �Tx4�^���B�I)/�2���� ��݂�B�I�
�>��@��)b��S'��0��B�ɽi���P��8k�����ĉc|B䉉U�.���N�#,^D-�*b6B�	0h ���$X~D���mBB��qL���#Gg���&߶<�C�� v�pu�e޶���R�JZ�@$C��S���hvA$o�����ٰ0B䉆`2b�؄��2z%����C�(�X�i� �>� �����C�		�}Z�W�B��i�Uն�`C�	�\� ���X�{����t��3+�B�ɛ_���rKŮG[�=0�둓ON"C䉓y!��(�dS�k~P�b5�
�C��
,.�PDO�y�2Ix����C�I�Q�	1��ђp���qD˟�TC�	�\�@���/�[���ё�\/�C�I�jG�*�`Ա	bؠ��B��Jg�B�	������+��P[��τ��B�ɋ\��T��^5f\P�큯+�B��4�)��K1U���Ҫ�'��B䉃)tbL	6��k���e��>/��B��=���(H�b~��`�څ�B�I)��T�Q+Z�H�vɒ�M�c�HB�IM����&�	q��$I��+bB�I!�\�uH�e�|��G�^��C�If�� �D�A�i)X�#P�J=d=�C�a���@ǉ�T[@�JD�ƘI��C�	N�8CƄ��CSe��`�X��C�I�+�tS�A< Z�L2E"\�C�ɚP�\�p����3�I��yXxC��6`$n� &,�?|�$�I�@:C�I,=�\#5j�o�m�"��V�C䉳m֌HqC,"��j����C�I/iݎ��ÏS��P NS�B�)� �Ra�E@�divm�pjzܑ�"O�'���{1IS�O�1X�͘�"O��+c���́�G�,>����"Or�� M-kk��i��v���"O�MI���?�*	I��T*$�%U"O�Eza�,�H�K��Pz0e"Op0���@�ٹbIl��)��"OT  oX���#@�@�،�"O
D�c��J4<�0����rd��a"O�H�ĸJ>� Q'��*h_�yb�"O�ɂFB�/���!�F�I��m��"OH$�s/L�I�XuE�e@`=:�"ON��c�C�$��e�B$� 7�48�"O�Ya(�dLiB��|��"O�܉�]�aV��#/�DČP�"OМ[h�|�	����,�h�"O`�2@a���5��A6�@��"O��8�FX��������R#j�ڀ"Or����C!kp`Â�ȏ1nEC&"O�ȉR��Zd��El���u�u"O��k�	DT�y2���g~!��"O^���-���.�iv��1�Ba"O�zDD�Z]��2�E�.?�6�!�"Ojݣ���3<0��oȱPZT��"Ox��т���mSd-�D�l*G"O�(S��!\�t@�Q,�?�"�@�"O�PV*�L�&�"�k׶w�x��"O���cMM#I�^�J�+ϭ8�숩�"O���;2��Q�W=�H�Hv"O�P�d�4q��oN *�Ƶyw"O2p���u���	[�F��&"Ol)��	�Y�<�v��8H�r�"O�@J�I̜6:�D�@_4\�nP��"OR)Q��ьnI�A�ʙ9z����"O:�9�"��)+Ra�r�I�&b��K�"O*�j� Ռ6ds�M�'(�",*!"O�p�� %v���~�Ĕ+c"OJ� �d��w�"am�ݲl�d"O�=��ɿ^�h�J'<t�����IW���I��s�h�����#Z>
M&ܔ�y"C̥*c@�)G��iw\MaU�9lў"~�"�h����4E�Tm��ΟH�T�D~b����@[��L�p���B��v�>�Il؟�˅BJP�0�95��y��	�>���S�4
�!���g�J0SD��/;�jB�ɍ��bd��� �$L�B�~�<���T>����K-T�^ ۗɋ+@��`�9D����Ț�Og� p#��=��)�!�OH�=E�dMG/]����m:2jZ��w$_:�ay��	-��R#N2PԸ����5O&C䉙#[V%@A�ʪeaZ@$m�1tC䉞pP�\x�o_�R��)��G, 
�B��	@iP}HRC"a�&싶MF�=<�B�	�jv�q'J�#�L� 1 E�u��$�
{fL�p��73*��A��#�!�d	7V��)���ʕ(P��!�D
gi�'=:p��I�`��x�6��*W���B��y��%��J@ܺ!m<�x�NZ�p<���dY�h�q� ,*�Ҁ٤%V!�D:����2�O*#j���:��INx�(ӑ��3]
����AD�:G'6D��[�,�;T�x��/�%��q2.5D� i%&3L�}
�fS����r�=D��C��
�.�4W�N+*���{ӊC�)� N�H��*%ԠA�w`��p� !Kq�'W�1&�ԁ�'�<2��P��@T�e���BFm%D��p�h�`W�b&�֊=Y��7���D/ڧ�t��a�C�F�R,�Ƅ40���F}2���!���g�W�i���MNZf7-��hO?ձB鄡W"u��C�!rY֨ 򁨟LG{���L��e� W_v+e�Jw"!���Tv����c8A�0%pT�I�Y�Ʉē{�
�(�ř�dl�ժ��c�8M�Ǔ�(O��&P5fx2���ɩ>֌0���xx�xk%=z��1G��
*H;6-$D�B��z(`IB!�x;XQ)_h<�ׄ@Q����a�O=a.p�v�y�<a���S%z�Z�	9{;Nh��%�t�<Y������F���V=$�
Ad�m?��؅p��)-�L����''?�n�Y(<�4��,K�Rd��G�-v�4��KPp؞��=�.�}�Y��,/q(�h�� �vx���'��)�3Ɉ�[���VB���d��y��)�=2=�F*Ta�5c���LkC�ɓ�N���.�<NH��)ސ�C��/?T���W�-@(Xn[�5H�B�	'x^,��O��.sz�x� ��p*�B��5;�\9��F������V<��'Na}�̨9�"�8�iL\�n����(��x�l|Z�B,�,�H]3 *P5�6�O\����2���Y�#�>�X��NL�\�!�W9	:����������.�9R�!�(
r��$薠5�0��K2q�!�ӡ=g>���hyLE���6�!��H�K�ґ-ϓQ\��d�ÕU�!��֟~�z@�)�Z)���HK��!�d,] ��e����)���q2!�䙝���p��W�m��AD;U��'����?	�B�|�قJӧe�ha�)�.k��Յ�P�����01͎HP���#0� ��>���hO���s=��'�y���D@��I��B�ɬ`H��ɇ`
;A���i7*A�|6M"���<E�ܴ&���0 ����"��5��4PjĄ�	e~Bm
�K���#�O�����X&jJ:�yr�j�	z?	���L�-��ծ�8h���qI\�v�}�����"O0�@�7��/6"1(&$�>yt�%�O2��'��:*uv��<op@���p�O��H�C��6�k�i��-�蠳"O��UM�]#�	�IW�xl�#"O�8jg̚�:b��q��:o��q�"O�� T��9BW<$�`H� m��z�34������f��ElI�d��)kE��A�<ه` �{]x�cQE�)�n#�#���M��q6e���L	Hd'��12��m��s��Db `�>	 bB戱�d��q��zH<GDWzM�P��DL��h��.Z[�'ȑ?�3� �*-y�k�NG�=�Fu��-D�<���Z�_X� ���<^�p�5$�� �'�'��>�(W��$S�X|I��B�4'�Á�,D�L��斌�D���'�ݘZ��D� eGaxR�K�DGM�p`�#p��I[@BX��yb��SWx�F��:#�$��H�bߛ�O�m��� we�Xxp%�
Jٸ�z��Iu�Oy�� ��u;�Ի��\8Y"�8�'��y��$�{�"%�7ظA=rq{�O2O��S�O<�j�@H�/�@+'➐=�V@��'u�]1�NJ!r"����B
�<∑�'�� *�J;\^3�N׬:ݨ���'��� �}�Wg���B0	�`� vB)�'G!�޻�}�5�I�J�F�s��^-!�Օ4�R���x(fkQ���L�Oz♒�=n�lm8���9wL��'�h��G���E{���"R2d��`�'�٫�˪c*�E�,��+#�	�'Z�	�4 H�j��Cч�WYz�2�'�$,�Sܧzx�Q@	��@ �q#a�V�9�ȓ2YeB1f�5��=��D0!�m�ȓ8�֭��l�>Xq��i�`��1�̸��<C��2d�\�Z�p��2l��M�L�ȓ1�Ҽ#!�()�Fᒀ)��n
�݆ȓgau�ˮ%X0�+�6�����<�h�%'��O�F�4R' ������`Ĥ^1��i��G�'+e�ȓv���#�aU�U�j�X�kf�P�ȓ@)��ꡯڞP�
�*�GE-�u�ȓSA�l�3�[w�&9P���BA��� I�V��D�FXw�5�RĆ�	JJ��W���X9�u�:<ņ�k^��S�ӌqO��;�hֽ{�"8G�l�>q�'��Ӳ?�)@p�� 8jS��zsTC�	8[��r��i�8��ʎ3�Z�|�H���y����!� ��Fؚ�����Ƣ2K�C�	/|�<�T�T;;��E�c�0lؓO���DW�,�E�C���o��ub��&J���R� ,lni�:T��ꓣ�!�I�7"Oz����U�JH҃���Q�$�#"On�с)��+�[����}j&"OR�NN�&��t�����5��@"ORAsc-�1F���Ѳ��r�(�3�"O�=��G/-	0�v�J�H�F$��"O�8�6�5i�ZZ�&��Q��"O��S��H08>� G�|��AV"O`�Zb�\�M��-�K�	�,����'?vm��]y��J7%VB]:��5�Ҫ�y�²?	����5;�B����Ix?���)<�9O�PR��&(F0�4ǐ*(X��'s�I7Bx�%��+8��0U�X�S�9�Ɠ9`�5膰좜�F�� �2܅�cܨ,;FڊG85�'�J��E��A�^Ш6�D�5Ҙ��Ӛ�p��ȓH\��WabQ1���OC��ȓ2�,��k�^�Ʊ���Ɛ}�����{$"M�[y{����'-&/�d� "O�� �)�r5����6��ih�"O.��� �C��X�2��\��8�g"O(8J�f�/l͑W.ܑ}��"O�h�G%R�RЀĭ��3jB���"O�p��ދC�f�7-ʍ!e���"O�x�4�P0N[�!x�K+act{S"ON��D-&Y��`�$�މ)L�`��"O��J��]|��JfA�'jP���b*O�X��h>(N��Ǳ>v�+ E"D���6 �	��i�,KRȊ0&D�h`��W�F�Q-�$ZZWf"D���Gʹ�
���٩?� �B"D�`CF�{��Q��V�'nFY�P�-D�`�k�TB�H
Rl�+d Y��
8D�l�gҵ{��r��44���ᗫ+D��P%+k���*��k��A�7�ǁvD!�$��O�J�:��B,q2({p�� K!�<aҀ@�ܩD����G � e!���c6���͇y{D�a��.M!�� �P�2�v�p��ÈA�*t"O����Kar��UI�
 �I��"O�(�@�D�k��񪓇�o���B�"O��y��2J��J�f؝F9q�"Op���^x$������8\rڈ��"OltIf/ި �l��dɜ9o`D"O"�I ��8^n�K�(^{@`a��"OH���_*]@H �w���F>`p��"O��!���5�H)� )O�dp:���b��%�dk �'����4"�<���',V3#4�K�'4P�Zv(ٯSy�l��N�p�f�
�'"$Zq���"�Æ�ͱr>��'MT`�e�=w��#V$R�d2����'��D����+Lٴ\�e��%/�Hm��'\PY�Gp�d�j�#7��yB�'^x{��
ǜQbt�Y7���'���X�'��j6rI���}ɚ��'�< �v@� ��L1���k}�i+�';d!�%�S&'�ԝSpJE�d����'qH��ɩS%� �GN��e�,*�'�\)� ��g�`,�g�K�
��ͺ�'$�=���Qi�S�,Y�p�'���!�Gʔ-���.z	����'��5pY�3A7�`����'!��-ɣ;�aa��S:2Z��'��`�Ϩ 1Z���b�ޑ��'��I*��\= �2"���B� �'���0�f�R��怙BF�I�
�'�b�
�D��p���0fry:
�'��`k��?"�1�k��?�z�Q�'{��i�0�H H����5���Q�'NTD3�Ć�`�P�Ұ��}:�c	�'H�͒#(�(H�Lu���X1`	�'��ӣBۗQXP���q��@9�'�f���^�(׎ٙ@��Cc<��'��{���7j `2��̤Ao�]a�'�Du�և��u�dl`��6
�\h�']���mT0 ��#�Kƒ<*��k�%�*n�qO�=D��O�Qؔa8��K�'�	dZT�"Op�r��xt�I�e�<ue�<�g�.FN
UQ�G^X�HA@`�r�4P1�wO��QO?LO��banJ:$����'.�jUi�:8,-r'�۽ ��\:�'yn=X��91"�I��hL�D0��y��̠N$�A�gVC�O�n��4BԜ� �2�2R3�q
�'����$W�V�:��H7B�j`�4��:*NxݥO^����3?��I
����nYE�V���A^�<5&¿z�<$��&T
N��+���Pf,�˧K�0hiF���I�e�[A��2hn@I�IZ<\�az�1;��T��n?�6���[��y�!(ՕV��9� �R�<�QE� �����F̾��o]O�Ȳ�I4/\QУ~r)=�\����	�t�HƟ$��MAZ�ޜ$�"~B �ҞbI��XD�S���`�f�+z �Ƥ�N�dM�U�>�S$���G/�VXRU`����Z��'�����
B٘���ɰWo��B�ƚ�%�:��&�R?nxs�&ڨl��P���I�^��A,�j�Y[�O�u¸�Y��4G�8$Q��;LO�$��M#��DʝE%Ҽ
B�Ϩ"�0@SV��Q���QAK�@/ƔJ"NOh�"����5�W�'��Ä.�-$ �ȇȓ_&ԓ� -\�n([3��0X��K�ł<Lz�5�G37�)��0Á\�.T�k]5@޶���O#D��;u㛬(���&�[�7�Ew-��Li�oI�VӼ�q`�JxX���!�0]���pd4%�Uǫ�p>��@��"���L��d�K�C^7z��C�g1
�Z�'��q�AJ�j���"�'��#�$�y����Y��
� i��c?�p�H�:�a!�H.?��`�-4D��  H�4�]�}))��	��jS��L��Y��Q�Q������©
�t�x��
\� ��X86����y�F �v8Pf.Y�,'L ��H-���2q̀p1���<)bn�13뜵�wcWZTY�ACx�PI2���#�"�U��*!�"�xU�:�
aA�-�K�<ɤe��^�*l���۬����C�<���o�R��D!aI�OE�<�)�3%먈�욦�>�gjAF�<���T�)��kc+��%�
E2�gK@�<�������S��24z���|�<Qs�M��4`BvH��V�G�<�ש	9/�u���xF\x#c'�u�<��l�m�|#�(L	OS>��Q�Tp�<����	��Ⴤ���b�����e8���O�&v1O��iuf�/�6T�Àǌ}��ˤ�'�v�p�Ĝ�8,�(#dB)4F�5@�,��	��I�Sl��K��Y����?� Y3��ĕ�}���@V�%G8� �!��"��I�I�4l@a��~zu�T�
�h��	�{�tHA	��a�:0�Q�U�l��˓|\�Ұ�ƔUs�#?y��Wqt��3��#�9�1O୲��Ǹ��y��_DlX!�!�j?ɴLí!k�آ�ÆDT�;GNƛ��b��/<h�����Z=��� �)J+0���(G Z�ae��򆐂��!J���B�՚WT��� �(O'(8ڔO(F"^�q�'�d�82��K��Y�o�>#R�d�'��u�-�py"��-B�ӗ
L�y�r4�@ �k�DrS,G>~�ʔ�����㖡�$5�z���:Ox$���3h�\B�O\��4�/Jc��"Έ$@Lyq��p5��K�	Nv �DK��!���-(��ai�U��$P��е3,"�`���Zh�q��N�$��d�����%���O�����>NT�E�
R�+s�q���O�a��n�&U��x鳏Үh��m�vO�%/�2]2U�͕:�<��f�j�a�Rn��a���#�g��2m(�R#�.�R����"�]	6�՝�J,�+D7H�J���d�L�Y������8��eݙs$��UrL�ja��q0��;<��P�kZ�{���e�`�X������҃�F8]ƅ�6I��y簠��fD��r0�#]�i����J�lcR<���G�?Q���}���<i���A/�a�#W�8���QU�Ks�'��H4��X<j���HMP��\Y�x['�e�����3~.��/�5vG��Y�'��I)ç�m���t��,Yp�Y�ݘdGG�	����.���s�G&>05 ,\�n�nX�� �=U`X����|J��In`P� )ύT2�i�1�i�<!$�(:��]P��6>���'QF�����3��y0#Cܬ;2Vl*͟�՛�&�]pn���wm �`V�S`��l ��+UA�q[��n��x��Ă%Z�y@�O��&C�`cD�U�N,P¥݆�� �DO`<P��(�'_أ=a~BDP��1s�\5�F\\�'1�10A���Ik���<txTtX�Û��yBI�K��H�a関������&����)��s$�D(u��p	�!>�Q��[V�T9 �� b����>�T�O?@yapΌ%�H,��f�"G����'���X0ɝ%]�2D�� �	?& �Ӫ�	��A�-B�On��2O1�`��Sb@��y�B�+*�T� ���0Z�)���x��*)ܨ)����M`�"�*�XXr�p�@��I(���-a��M���5
ҼE}�K^�4dXA�F,QR����bƣ��OИIe)�7�NAAW�S�����x�\܀�#ߎdB�JN�%��X�'�)��~��r^����U�v�A�k6��D�/U5dT�!ǁ�@��SS���U�h�z�C�&�ħ&�R�W	�@���c�mQ!Z��\�ȓ?X��6'�
�� B������'r6(����'�u0�MM�S;%�q�'[���֭�	r{����k�{�͐�^�ٸvhX���&�քr*xAW'Kh�>)�e,���[�+R8:Xay�إz�Hw��+$�v���T���O�%���	����I|��
W,\"aºx�ڥK���F�<�0�(ej��c�;3$��!�Byj�+�ظ����G���P�(�&�M���Ɍ,[��C�I�x̼d�F��, �D�2"��aC�=�O���5脕8Ċ\'?����ܕt���z'��c4h���6���CJ��rR��''�7Xg<�h�*"�up����2��4x�h���R�ܙ�Z��p<��B� %I^b���Ξ(Ke��C��'q�H����1D������6Dd��A��_(�Z"�,D�������%�6A�J�TP�+D��c�B/{�����_c A��(D��X�L��xD"���'�9	0{�)D�� H�x@�ȽKxm��ٓ���yv"O8x��>R��yH��3{ar�Ѥ"O���㞗K��)����x��"O�u�w�D�>�R�`Y�M���"OR�3�`�-+�pU���
��mY�"O�PW���ڱGJVY��	F"O�#�g� u}�T�e ��t`��"O��;�^1f�ЫpM�\��]�"Om�E��^�0U+c��+�|E	�"O~=�f+߆)d,�v
�#O�n��2"Ofc��V M���%��?ɶdА"O@t1&?u��3���-.Pڍ`�"O:x�!�1B)r�*�A�5_�ap#"O����6v��,��-05��P�"OBCmBy̢g���cu�y��"O�����)�����.�EmT	��"O�h�0�ƫʪȲ�/���:9 !"O~�bW�Q=Qg.����*�.}�"Op)T��'d���ֈɋ6ټ�*�"O`�t#[�M�ċdZ��MQ�"OX8a����I�TE�;F*pq"Oh�k��0VA��	EBơ��Jd"O�U��m͕Zg��o A�"Oh��S ̈́>>�tY��4�40�"O:P��CK�E&�U@.]2�x�;�"O��Q-ЖL�����KqX��"O�$��D�;�dd�-ҥ&r����"Or�{c�����Q�ƅk��y"O���íR���7�Z�.m�uqb"O�H2�I��3Zԃ�j�'KVP,!�"O�����
�
p�Ŷ#A �X�h�,q��HzA� ��a|���$O|�(C�T�:t�8#f��0=qs����p�9c���?���[�
�����^�p�ᕅZM�<!1���(�#�%��jN(�d�f�ɵkK$��/Χ���P�@y� M��b�D��M�EbTB�	<H=�t�0�`+Z�2��)�J��T�%{L��'bT����>apJ�,V�ڜc�I�%/�4i"*WDh<�e�r�-�eG�&�Q	1����N�H�NXYz�0:lO�| 7�
f�]����:���'�A�`!�$���oMǦ-b �[�$l��tʍ�>F�u2l9D�@��O����,5$�Vה��4�d��U݌�b�o�l�j��iB;>x��t���ZΩ8(ɀ:�!�$��\�PPL�<28&��f���$� �����7�2`؎�L�hg_Aش`�A�3X�,#f,4��{ǈӓ7��Hr;�f������v�4!As�� '��ԡ��'��t�L�a�J1A�J�2-G����D���Q���!��A�$���自Y�ֽ""Û
�����/�j\[�lR(+�jA�������=Y�Gm��pYt�:�'�0쀸>j�qx�f�QO�l��_��%rs�m1r�h�
{8�Յ������./��9ۓ �"E�!�ȓ`QX谰C�wX|�*U�à>C�̇ȓbh��؆ 3,��}�T� 6.|^�ȓ2tX��0`�Lɩ0�C�[)�4�ȓ[.�q��n֩fp�T���Bξ��ȓz��\��ӻ�	p����VQ��<⠸8�E.S*��Kb�B	��S�%i�E�)=�~X9bn�.H�,����6�=�d�*�b$��ܥ'�ч�1��(pK	h��ը7�Q�>HZm�ȓw܄q����8�P}�W�!�p<�ȓQs�l�����'�d ���A��5��I�N����8{.�09!�B��ȵ�ȓ���1�eШl��`KCş87��@��S�? `s2E�7|~�$+�60�$"O�4��ۢc���EJSY���)0"O�m���W���	'��4��j%"OZ�)����;�*�� @G#���6"O(]��A�4Ff�Բ�nɿA��I�"O"�ȢH���H���MGr'ʁ��"OXz6�H9l�����2,���B"Oʵ�egO
��t�b#��:�bxrv"O���#�(��D`�W�?Z>��"O` ���,d�.P� W�>:�A��"O<��6�S 0:¢G�?9��	�"O��P��R�B%�1���
�D2T��"O��Ѕ��X�v�cw*�:D;bHat"OX�zZh��p�Z�6�8uH�K�D-!�?R*f9��қ"�``�B���:*!������&ЦLC,���*T!�ۖ%h�Ss��kQ�="��#�!�~���R�Ӻh;h1q�.O�[�!��W=�X�'�KL=b9�p��0R!�d[�'6�x�F+�U/$�􄛺(G!�D��6wXE��/���30?!�d��zt��������2!dT)y�!�%s�J�h�'F�
�z��M�F/!�D {�
tz��G<M����,��.	!�d��N?�c1�R,t��1vM:
!�d̓L1���ƏW�c~L��G D!�䓀mCY0�dnY"2I�7C!��H�
��XSa���Ƈ�(!��їg�P,��&fl�!��!�$
�BB�͢lld�P�:Z�!� T�I�;V8�Z�IH%a�!�$�)I��P'KقF�����G�8�!�Ĉ�y{��p��K/w�*$) �Cfk!�D�s]��x�+
!�$� F�0nl!�$Q3cL,!`���(*�T��,E�!򄑋&�$T���NM� I��G�!��_%S�8������b.p�3@��>z!���1c'.d��F��@�Iш8!!�$-l-�B$�y.�ؒa^�!���V�.�6?��"0���8�!�]Ү�Q�M̐n�,p���0�!��~xvu�"-� u�&��t�]�3��h��G7�H����0�,�����G�&}02��g_�B�	�*M,5ʤ��K������e�⁠�D"NOȰ�AT�ey2��`��+�)��z��	0k�	�䌋
��dDl���� �%�Hi����8!�$]&i�(8�����F�9��0�1OB�	&��2��u����.�9���� �t"�u�!�D�'D�(#Gƃ�7�FU��o� j<H"$kB0��I�8F�"|�'��!F	U����w��v6�)�'�}9A�}x(�iW��{�D�{��X�a��'�\8�TSS�ٙy��h�A�ԙ;�n/LOb�2'̍�i�b�O�-��Dۡ��9�Vj�A��'�n]���ڵB$y
�NP�q��M+�y��Еu��ekskVU�Om~�2�B�'�[�z��%���O��w,�}P��O?����3���s�%�.P�X���b�:8B�#i?}"�����ɳ}5���W���	0h��J����L���T��P�nE�\1��FE�D��%QU�H$�R�E�X8�A��0n��b���7����tO8�����'|nx�O\Ly�	Ar8(�BXN l�3�F��(Oh�*vI�w2<8�D8����4�Iv!�|��Qr�ػ�bC�	�M�$R3��,P���[���O����D� 3���b
�����O�$�BQ� M���d^���m�"Ol���!�)y��٦�ʒA���z�OJݫ 5Z�$*vG6,O� >���J�k:���]�[��P#4�'�d��їIpn�"��]�*m� j�L��f�(#��p�!�$Q��
b�c��:k��8&Q���"C�T���JB�W�'Ky��1b%�(`xv��)їka���~��U�%�	N��Q���ғ{2���g�3^����o[4N��)�矼2kX�}�~)��X�;N@�{��&D�B#m@�ԩB�f�V����>���U4�B�z��=<Oрf���a�Z�����%-:�'>
$��i��H*Ѯ^8	OR�R�O\�O@�iҢ"OL���� -�l����hD�8�"O�c����K����E�Āv?�=[�"OL܀���%&�P�:��M��"8@�"O̽ 5�	���� jB:���"O8�z1,Мe �t�e�J�1[�$��"O�-���X�ت,�* �.F��*�"O=C u{� ߳L����	I�R!�Ki8�aņ��=|{�H��;!��j�ڐ��n��ksɢ-��xb+Þj]�1�<�!j�"M|*�X�{��Ы�N^�<�J��+�^%k��>4H�Ma~"
օ((pmx��|��iP�.����<E��
��!�J	ʵ{��)��):�ǂX���O��{�5���qO(hQ�D}=H��틇'k�|���'M pQ�|�p3��$���CS��?0쨁�w؟4��W��&X+;� Mc)ɓH��Pb�'�^��'(JK�Tg��.��RsL�]���e�  �f@:K>�����>@��䇈%=�H���H�z~ R���}:����	�X}����G׀ ��(�gc]-� D��}�a�C+b�4�i��D�SZ��`��J�'�8���S��F�	ե
5(���'h�|Q��`#d+xl�D�LOi�ܫ�>�4i����<�O~�=����O��)3	�xq���a��P?i�nH�L:���������%(��;~�$)����Q�å�ο#�F��fw��1;�'F�',͚7�贒�đ�b	�e���|�ܸi��jBJ6�\���M4�⸂d0}RY�6*Z!i�mS�2��I1��

��~�",a�Ę �+��!
:�iqK $G�rC�2G�Jb@��\Z��A����H�|�#�̽#�"�k���jJ�;��G�'���k�úT ��f�ѽfWp�'V':�YQ��,�ы���"�p�=y$Ǒ~:���c�r\�G��"�L��a��:j��Z-;��=9�JI�	3�S��0ӈ��u!���-�4ώ�E P�R�"ON�!dˉ)yL9B�'G�ء0 %ĜAQ������#�|lJ�O݋ W�g�l�¨�����@+�o�9q��`��	-�ޑy�ځ:8�+e�6��B�+�� Z�	��C?P�<���.m�FD&l̉Y� ��5�\�?1	�0%
lY"�֌JD���ĵ�î�+8������5����F���2bU7s�6D��K�z:䨇ȓn�a����q]��r�B�2L�m��j>�H�(�!mm�����~p���=I`�?9SV��D��M��%���̿T�
��	X�s�!�d�O� ��U�y�Ό�TkM<k���[�� yC\����#KݰD�w��a �< ag�6џp�B��i����TՋk��R��!L�zX�U���yR��q4�W�����%�R��d\�q8b(;����)�'y�`5�5@�.i������]�P�ȓ}h	5m�){ˊrѨG�5�, �>	�Bэ`gaH~�=a��%����G�8$�9�4��|���Kr��5�� �B�M#WcB��Q��gZ��+c�Γ,6aB䖵2�,$��	��u�>�3Ǆ��O�h�0(�%N��Y�H| �U�^p�z1j��_�Ԉao`�<��ET��j�C���D���G�`y2�ͦ7a�҃�]��]�*8�T]�'w�����(�B�	>u5Tг4�8д@�����[O�l3Р�;�]%?��Pԧ<o�b��4���7�
��F�$��@�T!:�����W��t��) P^ ��n�]��ĳ$'9cǠ�{�ON2wX�2�(.O��f����'dL�����4b��C	_�$����� N��P��\\��X�)�����"Oέ�BD�$^����A�<���"O��3 �ݯ-�!J�G�G~���u"O 13��O��e2�ǈ5[d��X�"O��xs�]��JY���Ѽw8�bd"O^��I >G6���C� c$��$"Otp0� _�1nl	Ba*tʴ"Oz����T�_=�Pp� Hwp�f"O�8�qi¥����N�O�^M��"O���\Rpyrd�h���IK��y"�A�((�GN;a���q���yr�L&s����f�>�B�m��y�NTs��Y@�H��R6���,���yB�+�V [EY�Nn* �ҏ��y�I�1J�r�+d�@6v�S�� �y�咩tJ|�+!*�?z�x����4�y�G\.!
������5�i��CI��yRh�d(ZRT�8 �8U���ά�y�X9|�i3��3�f ����y2��\��IQ��e/2m�dW�y§[�nw����!�j��J��y�̈́mra�CJf��!N�y���kr��[r�E(*�Pg���y�ъAH <p�e�"+���@ ��y��V�1�D�J��X�+��͚R�J��y�dף�H5�ׁ�9=� ��Ő��y�bbG�����Z�ν���K�y"KĿ1�
q���¯l���R�	�yr�R�h\��E+�2K+�Q��Ħ�y��
�P�sk =�MV��=�Py�kK�*��tP5Ɯ{��%��({�<y�
��a�"��W��>]]�]s3��p�<�#
e�ő���%#�c��v�<A��"G�,i�6�p�a��s�<Y�Cߺk-���¨U�x�(=r�*Ҵ%8��⎬)�^!��I!2�D��#�&}��m��Z�w�l��$>J�<����:`��DGtER���R��h��lX�y�!�N�R�@��\� ��$2��ϠV�'��0�	�U�jq�Kt�O��M�'H�;~,Ԉ#���'�t`�'2�H�7
\��L��R�ˇ��xɴ��u���� n�|�g���;bU�Ds��_�W�<�i�)���ʳK�MBV)�$_l��J�;+��)C�'b�Z�(R�7�=Y .G�����t�Ͼ.n���̃^x�����=
"z��g�B��V����uq���{���K���yb�X=���S(�>q��]�d(��p��uza�*.,~����*�'����P�wސӃE�g�@�ȓ%>�퓥���N���{eDU�b;p�B�\<\`*�Ʉ�O��C?�3}�L'P���hB�P��>	�� ��x*̔u�`���>5 J���(��Xi� ϷJ��cS��q؞�Cׁ��4��@Z`jC��:��<LO"%�	�|��A"R��Or���nۥI��<�E�D�6`	�"Or�1��y�`lr �֣��M�1��Q}�"܈��ň�^�БeG�)�����:GL��"OnD)P,��j�2�#,�#7"V��p"O�L+F'����4L��p���"O֌Ȝ�NF���L�/����"OH�B2���Ti��`҈+�fL1"O�Е�D5 ,9���4^�<
E"OZx�t�P8h��rd�M��~)Hd"O~0j ��iȼHT��@��)#"O��0��;@\�2���	6���"O��)�O�Y9 M�+ǜ=��9b"O�����P�{2h�`⨩X�"O*q��H�E�������P�hLH�"O� ���Ɣg{ �Hf  �ҵ��"ORUa��4 ���aun��j�pr"O�M3�'�=�tp+�D6Nf�9 #"O�AX4dVJ�v��qA�&��D��"O�EA��Z"n����
�b�|��$"O@Z��3�B�q�Ȏy�%�"O� 3��J�໳[V�(�6"O��b�#M�6�pܩd��D�%{"O~�GlƊb�]���>?�Q: "O��R �]�A�h"J��96Z��"O��R �K�u����C����i�"Od�Y�KYD�6X�Ц��pm�P��"O���� �Ȕ����V01��"Ot$邦
 ��[2j�#3L�B"Oly��	�{�fZEJԞ\'�ɠ"O�\:��U~ z�� -}��4"O�̠!ƃr$�E���L�*���z�	�m"X��'2�%�I�,#	 �1
\�x��9��'���+UB	��zLs�C w�z	��'Q %�ǈ
�u�4���:j}!��'���gnB;L��ĒG%�k��x�'���㥉 �Y����vH:V��,�
�'-Bt�VM��d�ܱV�\�}7��C�'�Q1�L]�;��x֭B/(��5��'yr���T�_��ؕ�_�t�+��d^�u���D�$$[Pvv����"!>��F��8��" <��V�$��CR�$�b��1���<)��;���;t��}Mb�ț �93ۈ�K'��!�&"�҄ױK
¹����t0��M Iz�� ܛ ΩِlG�<�� ���O^�b������z�~j��*��+7�<B�.\/W!��鷆H/�0|��@�@Ѩ��N&f�h�Su�h
vU��_(�`jF��U����"�\�h�@ܸ�h��6�(��i����[�t���ßf���d�5�ހ�Ȓ�jR��YA��.Q�֥P��M�:�.��6�[y��i��""p�b�B�a3�Q���D��!2"ל!G(��O��g�?�ⳮ�g��$��$_/+�v���>��p�/��\��cW0a�d�ʮԺꆿ���0���=}@���>�91qbA{�a�D��)W���1���g����	��ϙp�F�0#H���)�0��AM�9�Kȸ}$4����X��������͉�!^0����� k�u��j�\�{ܨ����*y��v�E��8�2"���|L�c��:2���O�,OR�!Ѫ� F��R�Y�WL�e��"O��FB�@�!cD�Եc,����"OX��%AK!9�A���;&���"O��`u/ɍt���AK4Ҕ��"O��CB�Y=2hx���,Y�9O�F"O@ui����N�#����]1�"O�x0W�@�v�|�����^9��"O���l�-rj���]/n~�(�"O�Yʦ��"��a�S�O$8k@"OV5q�,Ѓp:<-���\>.���i�"OL����ز4�f�8�)�����"O8��f�٘Y^�8ˇV�
4�"O�T��}0~,��LB��nЫ"O~�Ғ.Ѝ~n4eH�W7}��8�g"Ot=�"�ڄ|l��ڑb;}Q2Թ�"O�X���JO6"�ѧ�G�\=�b�"Oz%hC���$�4�x���0��Ъa"OD�9�`53��|���XVq;�"OZ40��T����P��J=(v�<`�"O�Ba�����s�b�$]��(i'"O�{������5W�n�c�"O�|��
�N�b�Y��C70 ���"O�0˃jZ0R�&��	�)��"O�1����a��y;���`
d�`�"O>%CР�
�&�SU�&x�@"O� ���S>�yx�#Ĉ$�&Y��"O>�A6Ob��
�(R���"O���!��G����,&@j=�"O�t3����~�L]@#�R׊�j�'E�pj���(7Y
S啜\1�h�'#��㞋lw�$Z����.��
�'Y B�_�`�6��-u\.�s�'�����a#X�D��eL����'(�����-FĩB$��b�8x;�'z0(�(Ƚd
嘔�W�nü��	�'߸�B��ݖN��d� 9f> ��'F���b��7�Y�!i�[���8�'3z�a��.O< ��e��6fPY�'�@t�������W��kіd�u%0D�<0�FNu�|��lH)}�V�R�.D� ��D.m� R#,Hw-@����,D�h±OQ�.�^|���;otd�Pt�*D��hG�YR�MŒ)D��#*D��iC����*HB�"��%D���T,�-�Q�giLFQ��#D�hz�)��C��dM֒QI^��u.D�����.[�PHI�f �:���+D�tA�B	�TS��7��(D�@��F
)D��-z�3���b|v���%��K�LB��,���@b���7:�!�.��K�B�	�i�6��vG��4�l���� BB�Ɂ �~�� b�O���1(ٸ`�C��0'�J��70��]�0��-���D�.H��Q��+�g���"�  T�!��D�(���un�7rx\R�- �!���s�q��8ięP@�[|�!�dO�M���O�+��M�	�!��ʱu�d\�w杇e���h *P�s�!�D~���ra�U�0�2Ѓ*�6 !�d�[��}��jCJ�Z3�F7!��S�}����C�M�UH���E�6�!��P%k	��)slR�n%0(`f�:F�!�d�5$,�}K2dS�#$����E�+�!�dĬ%_���E�?#�����
<a!��v�R�x6/�V����ga˔�!�Б�HK��3k�W� XN!��$7���5G�7{Uv��N�+L!��2�s��$qLDR���!=!��O�76"l����9j�p�4��$6!��
Y�J�#%ǖeu�Va�y
!�D�%%wl��&D4Cg^��c�ֱG�!��B�����^�OO*T�0 Ķ-!��6�^�E�ҌJJ!��2i�h3�L�;~�8���9m!�H�B��e�W;j��p+�
9;�!�ц�V�+E8R��i���f�!�$�6�P�	��Q'B��ID%Wj�!��F���è�*qZ)*�c�>{!�D��6Q����YW��
E���!�L�?Q�i���?ASvA#BD�|�!��8!�ܢ���J���A�ՏP�!�D�/&�Z}��$J4ﴥI#�?�!�$�u<��1hЯ!���[���c�!�$E	=WD�[#��)�g�>�!���?�bt�eJ8�P���r!�ā?N�0����h��d_�|X!�d�<[<H!
tAc�4!sC$P 3q!��ϱ;.0@kߍ~�<3��*n�!��S�K�=s�D�QɌ1 �/ݾl!�� X����% %ry	��D�1�:E(s"O��Ar��%<�a8���"�!�"Oĸ�-Q,g�"(1��ʚl�2�Z�"O���.��c�գW	ɂ2��"O��B�fF�ls��"jY�zW�(&"On�:0(_��:�	#�J:$Wf�"O��p��ߋ2���a��C��I�"OP`�g�ܮH+������T�"O0�Ô��.lP��b\ x��!��"O�2��ƕ�Ġ	d��Z�"���"O��k1m��b�>(�DaW�#��D�"O�{4-U��!��O
Tc�ؚ�"O�a�Ä`�Z��"�M):��B�"O�$�� �i��Дn��xl�¡"O���%@���q��r"O*̑� �J�f����>.s�	I"O>��#'	2u��I�M�+p�+�"O�����P ��B�LB��ei6"O�|��g)<B2�y�._0+�x��`"O��ZUH����[���<��\"S"OR��!
9J�\0 oP���a#"O���r틆'cF��Hի>�.y{�"O*�r"�[�p�"�ҀC�v�2�Ң"Oڔj�	U	*��y�Ѳ}�d5P�"OX�zYX49�n���6�i�hϐ)$!���Ȅ0dĲb����%e�z�!�D�{wB�PV��&A��Uퟘ.Z!�D]9m"yI���S4��7�Y�?L!򤖟��Z����H	F�ۃ �!�$T1S���AE� ����2�V�=�!�ɥf�T�Sb�4��A@��@�Xv!�$� =&�=Pu��T��a���+MX!��9.����n^2��3�f�~A!�D߱+���ZD�U�^B�xz6�ė95!�$�[�n�zG��	׺T+�h�6H�!�$��=�I��E���(�rȇ�Y�!��6V��
�.E�F�� 0(Q��!��J�p��͇��*��Ag�d�!�DP�Zd��ȥ-�3% 3�>K�!��Ε3�0()&o�2,i��q�*4z!�$ڝ_n4�gO����(P6�Ir!�ېO~���' 58��(�ץ^c!�8=S��@��&i��L�VD\�d�!�>SZy3���A\2�qg��'�!�B�w���c�g�Y2B���^=3�!��Z�iH� �g�w�	!@�9�!�$!S���y ������ g�L!򤆐b�PB{ ��DlH`=!���B>���6��4�zt�T��'!���>��xB*�(�sELL"!�D� Y`�ħ�"v������w�!�X�Oa���N��2���,v!�D�#|D��
;� ��+�K�!��6c�J��L�CŪ��~�!�d̮��-h�H�%��0�f�:�!�D\�5�D Q�]�7 !�e�Ł>�!�$�F�Q��J�-h6E[��=l!�]:�y1��h� ���5_�!�Ȍ7�p!�p%�� �&� ��B�?+!�dZ�p�l���%��;�����,W&@!���V�`3�^�U釪ܨa�!�DF�vz���`������f�V�3^!�Ğ%;^
Ez�D�CP����
d�!��ܚ	�.�Z�o��G�6�
�b��O�!�� F�B���P�t�{Í�`=j�� "O�=�U%���LBBM^�q�fq�"O�a�C�P8\s�T��kģ0�.�)�"O�X��HL�"J���%
�5	�0�b"OEC�	�f#�s���k�h:"O��jg+N�Y�n�YW�'_D�:"O�dst�։:��9�l�f]*���"Oz�j!�H�x���*6�7@Irt"�"OtqXvj�2VR��X$��/6�m�u"O�H{�i�d�AF��TPH�r"Ov�[SMB���%;�V�rڎ��q"O�K$"�0����Eˡ%���Y�"O*��R/�c�Nt��_!T��՛�"O6�C��v���jE�GQ�r�!�H�J��*��]5'/����,R�hV!�dE�_p�*K��1
4	YtiXQ+!���,� ��/ݠ �����ؘ[!�D�!1��0�1`�8}{�y�G�W�!�'&^�`���YOJ�b*�o6!��.���9cF�WvQ�Qb��?!�$��d�e�f-�mY�q�PB^m!�$�^��`�L_0S°�U� !��2��ӧ*_>�r`8_��ȓ?B`��7a�%|�A��O�X7�T��ͬ�H���'�ֵx�ƕ<�fI�ȓK̥"f��N���$q)rl�ȓ}KJܚ��2.{�pX��6eB����pR^`�gBD$8���ك�ȳ&>Іȓ!Ɲ����a�p̲���1>���ȓ^�"���gڛP�P��T�6` ��SEVْƦ\���Q��#E�h��+�H�U��/Pgf- Z	���ȓ{0xp�Q�k��rs��0LE��ȓ6���B֤�<yj��K�fM�ȓu�D�Z��P�=v��a��K�p����`�7Y�EÐ��p�֙jހ�ȓu `��@h� Ua���&H'�,�ȓS�҉JeY�Y�`i�c�O5��1�ȓX3l �.R<-��CsDdAz�ȓ�f�:�Q6�f0���@�lQ6X�ȓ/F5!rl�g���S�nN�"bՅȓ��-�GTB�Q�v���<�ȓVŤd�b�
&iA�1ѶA�3C�\��ȓ^��X�wOPLsR��� �.D�p��ȓ`�����I�L`B��0CK�/=:���VĬ�"rȮuZ�+5���c�͆ȓXj0� �  @�?�   �  Y  �  �  0*  �5  sA  NM  fX  �c  �m  �t  z�  l�  ��  ��  L�  ��  ɧ  )�  ��  ��  g�  ��  9�  ��  ��  �  M�  ��  w�  �  e /	 � + �  )) �0 7 I= �B  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�v�*���m���R �>�`�'�栨��¼`F-k��K��B	�'2B�z�� �g�-Sa��(AYQp�'�z�I��<2���Є;+fX
�'N�i�2���!'x|Y!l�Bq�,J	�'�P]q��Fd��4���B�4A�HR�'c�����<]6p���]�3���'��M�p@�^�0O�1cO~���'x[ŭ������5�J�T�ތJ���	&_�P�����^���z
Ȏ8����X@&!�0��e�PPfOȎg��ц��,8�Ɋ�H���J�L
;~줆���,	�.��M>֡��X���d�*��˖;c��0T��5۬������; �ld��h�BΏ.ƆHD{��O����DF>M���(�G�?H��'�R���CW99�T� �A�4��BO<�6�'��jэ�&u�,!��$W��A���yr����1Q�TM y��@����8�O�q���b��+T.!�}���ɍ��
�:��<
��G�VM�3��L0C�I1-�X$!�BQ�O��Q'��;	#>1����6+����eyJ��@���!��<e����k��m���E@(wg!��ɾrB�#&��UU�l"a�!�D!e�hLZ�@H�E:D�3�-t�!�DG!{�"p(C�����,+5O	u�!�\)��壠���@` 8�fN��L�!�䏴7��M2���i;�D� N·/�!��;H_��Rb԰m4�q��ML@�!�Č�O@�(���[�,��-�3�!�Ċ���`��;[��r�O��u!�d!$ 4�ĕp,�Tɣ��'!�уM�p�K'nэ5��-����v�!� �� @���JE��B7�E%G�!���5;��Uz�)RH�@�Ӝp�!�P�y�"����� b��"Z�$!�D�^`��9E��.��%`3N�3&d!��"tD�qc0E�묄�&腷p!�Jˤh��� �W���盪W�!�B�d�Qӂ{x&4g)��/&!�Fv%!2'xu�1��ӔH�a|R�|��	2U\���C�'���Dȁ,�y"%¤~��5뀔IȲ|��i;��'�2"=��t���V�A ��qE=�1id"O� ��B�$�2j
�,0��J��r8�h��燾b���a⨇#M?:t��C3D�Щ�(<�ԑ�r���M��$�2D�<��ͭ'I�`[�^*VD$e 4o0D���d��|:SHڼod|���b�'�y�i
�f������ūk0z493CZ0�y���<܎b�@��2�H�C©I�Ǹ'H��d�9H���\/�i��Q�i�Q��G{�O�H�6�ҥ9]����} �1Ə<D���dؤ }h���%��.D> )����(O��'�(O`QFM2T<�k�9���i�"O`0x%J�?C�������Q��%��Ov�����f4"��Q��|PђP��#FtB�I##�$AD��
_X0i��GuC䉲�F���f�7$�h�T�V�>[�B�I�|�$rc����� ��Sy�B�I�,R��Ā_bѶt�G_�H3�B�	".�F��M���9&ǘzIbB�
��|�G��O�ʗ�w!Љ$D����(r��s�̔�b�;��"D�؃e�4-fx �`�V:T���DK=D��⦜'s	��S�'	����@ D������E|:B	=��*�*O`K1$֔9�`P��#��`��"Oh�KүoXL0� CϨ{�<\�6"O�$�"O� t9�S5`�h1�"O"����U(����z�2���"O�ų�H��M5��t	�s�@"O�,�jU%k���Ȗ�Z=:a�]�"O M�ϟ�G�d[%��|Y<��"O$���"���C���hSށ+�"O��h�H�����Vh �Z6
9aw"O1�`���:o�xY��+`�!1"OxtQ'ၱ<������䘌k"O>��`/C²9jb�Ц	{8@��"Oh��"�	_j���*O�n<��"O|���	�����v�қ/7�}��"O��kF���Ce��#� c!"O���K���L-�aBB<c�H!V"O�9�a�n *$�A���c�昒w"On4`#	\%X��9�'V�IJ�|�"O����țkz�hE��'YLpQ1"O6��H8�ȼ�AkH(cGj!��"O�`�_�4�����F�D(q��"O�;�T}�� !��EA2(��"Ox����Ply�5�S�P.����"O�A4���[r~y��Q�@̖P��"Ob�
�B�'A�Eғ�^eP ��5"O�TJ�"[ ����H�<*<E�1"O� f
��G<�ᰀ�E�
:q�"O`��,HP4��G8\�|-�g"Of<�4L�84�Y�fF�M>B}�"OR��&�S�;�Xت �{3�%�D"O� �e�/e�Q�c#ؽ��@�"O�4��nëu�M���:�zL{�"O�Y��hŎf�8P2�C҄
�fr"OBt�p*F�s=��f�՟W�8h��"O��є��d�L�(� �<�� 1W"O�E�dk�2,�,	s���$�p��"O���$�	I$�����x��c%"O��CB�0�IBr���^E�"OJ��a� l����D���ޢzX!�dS(	W�L ��ي1P��['�C3o!���%�� )4��* ����7��q�!�� �%A�(yxl#��!}J�8��"ObE����_��\8SG�:�Ly�"O����bƐ��$D��zh� �WW�<	��V4���uj	�^9���U�<Q�N\_̝j�oӴm�׉<�?����?Q��?a���?A��?!��?�"��D�-�0��n΃Qp�]X���?���?����?����?���?��L��H�E���qED3r%�y���?����?	��?q���?���?I��=k(ׅ��1G���5%�xj� ���?����?����?����?Y��?��y��H��/�7\^�w넀kw0P����?����?����?��?����?���U��T�M3U�6���	
'N�C���?Q���?y���?1��?���?1�U���`"]f�4��lC�6C<���?���?���?Q���?���?��$E���T�0`�>Ff^�p�I�ٟ������	͟���P��֟l��ß"����n�A��F'a^��i���ӟ��	��\����	͟���֟�����X��W�m�t8�V�ߐO���$h�ܟH��ԟ`�I����ş`�I՟��	ޟp�� W@S�a�+���$����Eߟ(�	ߟ��I����ß��	̟���ݟ� &4
�I5��UV	#U)ן�Iݟ���l�������� ��՟$�3� myeۄ	���ǟ��ɟ����l��П��ɽ�M���?)tA�*uv`�7!�9m��a
���(O$�D�<�|�'SD6-T(6#�-���=Bd�	r�O$fV�0�!��ppڴ�����'9r�@`�ӥK��(�֑�GGH�"��'
��0�iW�I�|J��O��.z���SŇ�~���'/�Ρ�<�����$.�'G(<�	G-�1w4��%A�
xER,P�i9��'��c��0`��wh���@���X����VT�|��'A�<O��Şr�>���4�y�!�#��9��\~s:�1�'�y�8O�a���"ў�Ɵ��%#�()ۘi� a^@�Hb�y���'��'�46mS;a�1O*\�펊g�L�`���Q�ج��"�I?����O��d{�0�'t ��,�3U���V�T�]%΀��O&��J�	��ه�?��OB��@� 3�`e����~^�p���<�-O���s���GJӂ{�j�agDيqJ���R�z�8�ݴU�*,�'��7�)�i>�QW�Cx�l�SǏ&Rߐ�Y)u���	�4�I�}F��l�l~8��@��]���kؠBT�i�QF���\���|rV��S��@��՟D�	۟H�Q��-tt	�A�*mkv���EybD}�&�C�O.�D�O�?�����:&��e��l�bLRw邯��d�O@�$2���X� Abuo� ݕ%�".%d� w	��Li�)O��@�B^��?a�E.��<�2N�\�PT� �V,��	�@�z�p0ݴ^�tl��X�,a�tY5�	: �`Y��o��F��In}��'���'v��#���!P`��g�A�V�M�l�枟|C�D��E��Dd�T���Y���^�#>�8��
b�xQ"�}� ��I�,?�L�3�Z\R\�9El��D����䟴����MSd!_]��s�^�O�e��6}���$!�<�X%yA��f��ԟ mz>�y5�	ݦ��'�2�i#�G�M�FyJuk�MAxH�Dk�7_xH�ɦT��'\�I����������4=;�UKVD�S���9��[���������'T�7��-5�����O��$�|�5eϠ8B���S0O�ZВR�Q~��>�A�iФ�d(�4�
�I�#}�=p!�Ȱ0,m��+629F�7��[#ʻ<��a��$���� �kS�Sa�ʰ*N�(�V����?����?!�Ş��	ڦUJ�@O#�u�$jl��YU
B�@E���	�����4��'84�^����J�~*�#G��W��r���nɪ6��=K �FǦ��'(!�*��?]��Ziy�^}�,��`őUr�@<O���?����?I���?����򩅞<�`�i��hn�Q&f��aJ��lZ�O�"����IH�'-���w,�щc,��.T��fR]�N�Z��{��n�&��Ş`w��*�4�y���b7^!`�d�w�������y2�-VS��		^�'V�i>i�	%���q�&y���p�	jw�	��؟��	���''6͖�V��d�O��4rUT���� ���������*O��dt��%�d��^|: J�1��P��C:?�t���y�Z��`��_̧t�J���?ق��`2�Q�/X�J0ሆ�?���?a���?i��	�O�A� ��?�*̰��K�1�"}R� �O�nZ�I��y�	�6�i��O���*K�*wO_�8���.�z��d�����48���҂L��f����Oݵ9��e��47|�QWN71\��d����e'���'���'\��'���'{�4��fM�3��q�pL��n.�%Z�T�(+ܴo(tc���?9���'�?����0��)� )��!�Pg��	 �M���i�O1�� 9cFI�>�"eB�/0�����,�4H��f�<	��Y�95���O�䓻���j���c� ��0iBL�K�.�d�O����O�4����&�B�m��(��<�x�uH�U�u(�O�k�Jk����+O�dd�mo�r.eB��ޜZ�JA��ўP������m��?a1`
��������L�� 2�B����0yAbb��
b:-�t<OH�d�O���O\���O^�?�S���|�s"G8�V���c�����I���R۴%��(�'�?)��i��'h��y���;޺uq���[�|ᱤ�|��'2�O؈��ic�iݭx@��)C�T�Α!'-�@*EMP<X�T��'h��'�	j�VP�I�穓p��Ȓ��fEx"�j�<; )�Or���O~ʧ~�ށ2�O����<�`�5в��'�J˓�?��4r�ɧ�)��@���sv��!��i�#O/j��h�@/��_���2��<ͧV�p�d���U�z�8S�ŏB�&p�e�}�F���w����Y�mCd �᎝�Vut����P�c���?y��t��v��n}2�'�`!���>�F)iuD˔����'���\�暟�]>�B5�S���I'H�0�Rl[�bT���(��+.��Iny"�'U��'���'��R>�0ƅ� O^XxQp�O�(�=A����M�G A��D�OR����[��]'��@;�F|�Թ�ۛ����	ԟ(%�b>�����͓xO�v�ŜT�TJk�-*�h��k7�����OR��H>�-O8�d�O�`��L�O�˅Ǟ���\b���O��OX�D�<a��i`f����'F2�'��!'b�_e�hys-� HM�����t}"$|�
<m�4��Y�d� O�W��
�%�+nn"��'�:��%	Do�J���(ݟDJ4�'`���݊�Ա����C���{c�'��'�R�'%�>��	�U�(�q��	aDPs����V�
P�	��M�@A*�?Y������4��`3eʚ'0m��Ś\����E0O�m�M[��i��D0 �i���5b��Ox�`�n�u�j �����YsSv�	yy�O	��'��'����_�I�/z�0Xh�g��*�I��M+7(��?i��?�O~r��8�i�#6�� �!
����Q��	ğ $�b>e)e��)B6��Ϝ�6����Ӣ�@o��#ă�Ly"�ΝJ����b{�'��	�*q�l��l�1P(�lP��N���	ޟ�����i>9�'N�7�p���9�H�:��ܸ:�8%��-�jp���䦅�?Iu[�p�Iԟ�]2fX�P�g��$'�Er�[K5�r/��)�'g,�i����?�9�����w^�c�dЈ
;�- aG!k��*�'M��'Gr�'o��'
�ڹC@۩v9�]�q��1]��({1(�O����Of=n�(x�'$���|Bcpx�qt���&��ŏB�?6�'�b�'{�i�[_�>O8��p`63m)[D�!���Y:P�8|c'�🸲Ր|BW�0�	ڟ���П��3`H�pb,y6Ɇ��HR��ɟ(��gyr$`Ӗ��"��O8�d�OʧK}&$�f�?%t PFhW#]�x�'ۢ��?����S�l�"�`��j�-gޘ�2j�(��*�#�j��cY��S�gbk�w�	
U�9�Ũ�rε�C�Y����ӟx�I���)�Soy�j��@�v��	��X��=R-��m��B��$�O��lk��.���(�ЏI�yW�)�Gpz�}2�ڟ���т	oU~Zw�9��Op�]�'��5{d+�c��v�_xi�A��'����`�I��������_�Dd�U*hlI��^����)% 7M�+��ʓ�?yJ~���f���w�����:I�(��&�f:d�q��'�r�|�����x��6:O�<�@������KV=*VV�
�?On�Y�阫�?�bE,���<+O�@�0��T �P`ʄ�_>��t�'H�6�	�.�D�$�O��� ���U5��b1i��b<����l!�������O��$/�d@�?�Ƒ�$.�4v�!�J0P��83�lR�eP`�n-%?5B��'�n	���|�IC+U�p��!i��EojC�i)�D/�>!VT9G�:R��9 �O��nڄg�J���ן�Hش���y� ƕxN��H��$K���AR�.�y��'���'�Xm[g�i\�i��@���?u�W�@�<W�$#�F�&;R`x�k�:r�'�Iß��	П��	埤�IK稬���8?���m�>zT�'�r6�X,���D�O���;�i�O6zsǌ�*a�!�T8�TųWK�h}R/kӌam����|�����gMQ3)�yK�lQ�)�*t�L�. `!��ۜ���0�6��msP�O<ʓ�xX��%A:zB���T%�Y���?i���?���|z.O��n�v��l���1����Z=�Y��_�d�4���.�M�����>��iՖ7�ʦ��A�W�vI	#��/���p��	�<=m��<��8 @�����'u���w�(m���[�k�<�5���~�ʉ	�'�R�'	��'���'����r�%F�lC��Ï������Ol���O���	�;����Oԍo~��.I������)C��3D�J>E����5�xb�~�`�n�?�
���֦	��?�%��|z���B�΋2��Ԫ�N:?�|!���O¼ K>9/O��O~���O8Z�Cv¾�D�9j�����%Sj�����<���i����q�'�'s���w{ ��d���{��� K��S�̍�'��[�����<i�O
ʧ�?9��,�2D��B�,tM��7�'��yS,S//@y -O��Ɍ��?Q�!=��;D� �G@;BιsE��vc��$�O��D�O��4�������=�`�a��NF�I��O�(���"D-ْ)�xh��'��'�RY��ScyR�wӶ�r�&�{d\��'�I0X(��'EY���ߴB.1ڴ�y��'{�5#C�<"���]�� JD�V�1tip���됋D�`;�9O���?���?���?����C�r��<�G��c�TԺs�"?��4o�A��%�	˟��I�?!�O/���y��G�Ҩ���^��Q1S�Vy�8��O���y�'��'z��аܴ�yrcΉJ�2��A���J���yBl�.2l���$�'0�Iş�I/B�T��GЧJq4P����.�y��ğ��Iɟ��'V&7�B���O&�ăm0�`���Q��T�J��)�6���O����OP�O*��E��]]>Yy@Lv���*���t�R�؟^�a��Zw�S�_R��򅧘�m�ָH� �'�VI���h��ş0��ڟG�4�'Hd���W�:n����G��L�� U�'�7��;���$�O�]nZE�Ӽ�d�����$Ò<k���RQ������şP���b���lZx~Zw�d����OL�(s�CXW�b���Z?b��R��`��Yy"�'#2�'U��'�R���~cLR���u]�|�g5 ��MKqA?����O ��B���'>�
Hi��^e�̼!F�ѪW���'wb�'�ɧ�O3ޱju�$�����+/�̑{�G�nm~h�d]��3������g�IAyb��,���@ ��.��q�7Lێ3���'>�'��O�	��M�!���y�+����f�@�������?�t�i��OH�'6��Ϧ9��4?!�8���S�4iY��@�UP���b+��Mk�O^A"�����w��ѻ�/Ƒg�F��B�)��a�'�r�'@��'���'�����������Ib�83�vL�CF�<Y���v-����T�'��6m ��ȏ#�bъ��; ��!���6'M��ON���O�IѶg�,6�!?���1s�7"�ɳ7���ڥ���?� +��<����?���?�&֬#�Ubr��)<�"5j� �?�������A�gNğ���ן��Oo(�ѓG\.\����S�Pb��)�O� �'��'{ɧ��@[�K�aƵe�1�
��<�1Ѷ�Պ[%�\�<�'\)`�d��IJݫQ�ѸZ��� �^�I ����?)���?)�S�'���L��m��L�D�l�U��>ed���(�/m��)��ퟴ��4��'<�ʓ�M�Ǐ��Y���(<PT��Op¾i^@1C�i���v�,��"�O�'8XXVhH
��y�$��r>L3�'�������ϟ�������L�Ԭؖ��f��(B���q5,X�J�7M��~���$�O��D9�i�O��oz��;7�?.����Jq @�
�?�?�����?Q���?�pA�ۦu�`�Y��A;��XI��2�4͓Md����Ot�iI>�)OX�D�OP��V�Š$�Ih�ʆ4�>M#�)�O>�$�O�$�<ٲ�iM�qI�'�"�'b�I�
��=):�jש�Z�ԓ$���^}�(n�p�	m�I0Mt�2NM31\�!� ��Y&��g6��֠�C�XdIL~����OLd���p��# �3sv�͛��N� %y��?���?��h�4���I�nu����@ !y��]z��D_զ�Ag-�⟸�I��M���w��P��.M�ҁ�ϝ=��ʝ'h�'���>J3�晟�]�)�����8����_{0�����59L5��|�X����ğ��I��@��ʟ���� p~|�!t(��0j�0����Uy҂y�Ԙ"Qƹ<q���'�?�'/T/�:�sA����D���H21�����MKE�iQ�O1���b�+�,en��a���v����!����6�� �S&�� K�l�s�	Jy�]�j��8&&ۮ�@����^7/���'|��'@�O#��;�M��F��?9��|�4K�σB
l�����?!s�i��O�	�'�B�y�͆2�� I�H|�ѡD����3�i��	DTi��OB'?M�]�R�x��֪m��-j�"G?i"��ן<�I�d��ӟ��Im��nDVQ��lM?�v�k�I
/}���?���@՛F�ܖ���'��7-1��<vώ��,�w��;��W�9�t�OX���O����L��6M{�x�'[Ϝ�0HL��4���HF��l�u��?��i$�D�<��?!���?y1l�6j�����J�!��52�f'�?�����DHȦy��j�����ӟ�O�H8Q���qF���]�j��ň�O��'$��'�ɧ��'��!�h8.�P���:z���ⓤ�,�욕�R�s����?e���'?έ&������+ݤa��F�[j���#���̟`�I�b>��'�v6-\�k1���( �l( �r��X��0��O�D���?�d[��lZ�����٦+MPDɷ�"&�V@�4{���R�"Λ6:O2�DW�u�"Q9��`�˓V��@҅۾u��p�I^�v���ϓ����O���O����O���|����v�|��bM�E��U�]A���ě_Z��'�ҟ���'%`7=���*s�]�^[�L�vg�-f]���4B�ꦹB���S�'V�d�4�y�ˇ��D+gAߏ1��Xႈ�&�y�NȺr���	.��'�	� �	8)|d�97�E�rC���RƉ�P�����џ���ß��'^7E�^Q�D�O���O�b)�-���B���7���1���٩O�(lZ��M���x�V ��yAf썗!���怼��D�b#���5�Á{z�������yzb�dP*6U(�	vƋ�$i l��6i����O���O��D:�i�-y?�)�O:����^ d�m)�OQ ������Ot%mHt�9��ߟ���4�?I+O�9ﶈ�G�֛(@ u$צ$¤���r��mZ�M���i}�p �i9��Ovi�#��Lk�e�? f �1�N/�.02Td�4��bC/�$�<����?���?���?�n��7�̴A�Yi$��F͚
���y�Wd������؟�%?��	<��1�"�V�����N�h�6��O��$�O6�O1�p�;��ҋ�T����?�|��e�	>f�81A�<�qN��-�f��ń������,5YAc��Q�r���� )� ���O|���O��4�n˓l}�F�ـO nެ\�\�q�J��pR8d⑥�)9��dq�V�ds�OdtlZ�?��4P��N[30ۚ� �����2˒��M�Oj�B���%���������_c�(�'���1�X��6O�$�O����O����O��?���(�~�< ��E=>Ġ�j�Ky��'�7-�**S��O"LoG��@{@�١g�2v���܆N͸DL<��i[87=���FzӜ�+��ם%�4�_�B����eM�*il�Ti��j�O���?����?���y���h�H�u�X*sL�,V3�I����?.O��m�	!l������i�t�]�n�d�gC�+GvʬjfA�����u}Na��oZ+��S�4�[27��a� �^�
����F7�Mq��	
���� ^��
n ""�j�I�%V��*v���8Ȁ��.)Y@8�I㟜�Iϟ\�)��EyRm`ӒUx2��X��ui�L
`0�"/F�Xc����O�Al�d��45�I�MӀB�3"L���V(Ͱ]��dy��B:8)�V�i��b�)x���֟q�0Cn�T&KIyR#[�0��T3��Uy�!��"Ҳ�y]�����������ןh�O��(�d��Yk �2�.Z�uQ@͙"+gӜ�0+�O����O�����X��])���G�<��` k[�cFVԙ���M���|J~�$ � �M3�')T�J��P!Ц��Z��Ì?�y�w���I�.z�'s��ޟ8�	(�6���P��\�x�k�r�M�I���	ğ��'��6MA��$�$�O�����
0�hC ��f�D\��b�1w�⟈ˬO8lo��MQ�x�'�[��i+�MǛU�T���8�����z�P���ҫrkf��h���pk��$O=
:=��&���8А%DX�S�����O����O��'�'�?Y&cWUn�Q4�G����HB��?�?Y��i�2���'K��b����6�� ���M��,2������	����Ts�@ۦ�ϓ��D��~��d�I�*D�oL�,�D@S_?k��@%�H�'Q��'��'���'c�LKM�]�1� �Ўd��ER�d �4V�(���?���䧑?� �*kŮ �6N��GB���O�B���ş<��o�i>U��������+V�B6@M�Wں�*�)P	�>�����}yªX�@N `�	C��'M�ɵFe��CW�#-��]��L��	����	�i>)�'��7��8.���dA2Y�4����(��}P���5������?!�X�x��� oڤ4��\�7(�0ԭ�RD�-_H��a��@Ҧq�'�|��IM�?%�E���w�8-
�d	���!�&J#�u��'I��'J��'���'���H���B]3�(�"���Qv�_c2�'o�H`�6�,���'�^7M0��\�T�k�E.U�azVS�C̓Ol���OT�d��@�^7�`��yj(�&�H�:�:0d��@Tcf2�?��:�$�<����?	���?�pK�8?IIC���
JOX��!\��?�����ަ�c�D֟��I���O��m{cKm����O,!�x�Oڼ�'k��'4ɧ�	_�u���.>G��QUi�}�� �/Q�\�֜�d�����i>1K�'tP&���S�>"��#���4e�"���/�d�	xyr���O��I8�M���7s���oʪTT�Rp;%�0u��?)�i�OhP�'*�U!���� ��@̔p���}��'��L��ic�i�ٰ@��?�pP�,ha.{�l1���[�0��%Mx���'Kb�'1��'a��'���4�؛`j\�2콘1�Q>"�t���m��M�	ʟ���^�Sʟ�	���#��h�X��ƺF$j�����%~�$�$�b>9cl�ܦ�Γi49�S�x�n�H��̓;�8��`��O~��L>�(O�i�O�M(c�ӞA�&ɛí�"A�,�'#�O\���O���<Q7�i|�4�v�'w��'�<2ׁ��y���  �9���B��$�x}ҩx��l���K�~�CqJ�^��h��M�W��d�'���! dR>+"M�Ý�����X�s�'�&�3�K��~U7ĉ"��Q��'�r�'ar�'��>i�I�</\8���
�9��=YF���*@���#�M����?Y�\���4��!#E��YѢ���m����=O��mZ��M;Q�i���6�i��Ɉ2�n�3��Op�\�c �"�&x�2n��GV&e r��u�`y�OY��'���'�r�ކN�Y�C�4D�@4�^O����M;'���?9��?�I~2�2���C�@�$@x1��ȫw\��(�43��� ��I�?O�T�!���}Θ�b�D1뚍[����P,��A���OH�`H>�.O�=
���D[���oL�9��!z��O����Ob�d�O�)�<���i�RDf�'�x�z�)g�d�KT�9l�Z��J�O plL��H9����Mk�i�|7-Ș7}6�S��ھq�]Z�'����[g�s�h�B�nu��e�L~*�;|��tJRHJ*6� ��憰zE����?����?1��?����O������/�B/��l�j�J��'�2�'��6-]%'��I�O|Imm�Ʌ.|�+�ȏw2P�bQk]�W��U�J<	Ѳi�\7=�~%+��{�
�	]�� l�iׁ
d$�e☑Ghͪ$���?� !/��<����?���?�� �K�f%� ��� ��T��?����H��-c�H�4�	ӟ �O=(�Ь[�/b���C�A�A
�OQ�'R7�WŦ=�N<�O���
��ܵ��@:��&%-�����M�`|���H%%��i>m��'��8&�[!疃~���#�Zl����C�����П��Iҟb>!�'��6�Cti�7FO�k��d�g�zp�Cg�O��DߦY�?��U��2�4?��@)�%^ll2�J/Y֮��i,7�A��7"?�`i�%Qob�IJ/���J@|�I���Ro�QW) K���<���?���?���?q)��T�	�l�X��E�$g4���ڦ�tb@ٟ<����'?9���Mϻ��E�4 Sfw�x#7N�0Q������'��.���4-B)��0O��+D� ^F Pc�6s�� � ?O� �ǂ�?W�&���<����?AC��`q�=y�iH�ļ�1eN6�?����?����[Φ݊� ޟ<�	ӟ�з��<G���1nR��XT�KJ�^����M�`�iyfOZL���q�d��V�z�P�֕���O	2(�i2>��2 B˟�
`�OR pp��L#q�="��O�l��͟|�I�����ӼC��ߞT�!��>KN@��tkD��?Y��i��1�'�'���k�ړO(�4�P�i��ɇE�z�S��J^�$�	��O<6���e@�4O&�$(ݴ�y��'W����?�c�6���P�cI`��`G���K>(O����O���O&�d�Oiq�U�)�y��-ar�(j�<Qf�i�L�3�'�2�'���OG��'���3��wq��@�u#� �@�e}�oӜ��Ip�i>a���?�!<Y����ЃD@,���OG�������byBg�1	h��I�?��'��.3sH!
R�T���&�ź4%�I����	��i>�'�$7��-�~���A�8��"�Ǥ_����������Ŧ��?�0S�L�	����
;� ��^��س�� $��A:��
i�7�-?��W"t����0�䧗�;s�G1�:��f�X�5t 5���<���?	���?i��?���d2l�BA�?R�@<1W�أ;=b�'"m��=f7�n�$���&���Țކ�I�����9ǂ�!��X1��|���N	v�7#?94��;WN���3]�P��s�H�2�1ic��O�1�M>I+O�I�O����O��R���d��¢JI[2�JsF�OF���<�R�i� P��'&b�'�S���a $U�a ���[%��,��I��M�&�iGO��1e�9�P�øer��ٔ����� �O���LHYvg�Ky�Oh����9e�'�  +�15|Ĥi��.Z�����'�B�'�B�O���$�M������P-^�=�f0X�J�5!~��.�O���Uʦ��?��P��oڼPXd���o���	!�V���`覩�ߴe�nBٴ����<1�2d0��#���V]�'˷��XB��+�����Ov�$�OF�D�O��$�|���A ̄����A���C�G�h#���
��	ܟ@&?	�I��MϻO�Z����n	Q�ʔA h0���i"�7��w�)�S#n�@lZ�<�Q�Q��m�d\�|el�r�e��<��+�$A��D���䓥�4��$F���LB VS���s1	�&Z�Z��OX���Ob�[���=_Rr�'&r�X<�:�j��T^	�E)N�:lM�O�|�'�86M韼'��� ֢Pc4�sB3t$E�d�)?91���)+�X*�O���.(���N8�?Ya���\�F�J��r،(�ԅ���?Y���?����?Ɉ�I�Ovm�r�ɴXta�A �r�>�8���OlnZ�#����ǟ��ݴ���yGNX(4�r0jT��@0������y�g��Dn�?�Mk���M+�O� 醑�"�F3>d�yç��"����" <T[��O���?���?9��?!�g�"Jv�� fhF5�r�ݢB�d`�/O�lڒs������q�����hv�(�rY��I[z씢d%F(������YشS����Oup�B���
\������_H��������U� ��>o����E�yre��v�8��Y/�N�;�-޻K��'���'��O��ɿ�M�%�?I�ȉ�D�[�I	�<_�a�tI
�?�$�i��O��'9�6͛妩��4;��`��-X9�%��	@s.H��̟,{��lR~bM�hĉ��r��Ov>a #��!��4�Ce �]���KFQ������N�4x^���K[�.\lU(���5Բ�+�f�A��u�DT����;�BA�?]eY@㘛[Qlt��ŐO`�;�F�����U��|���	("�BHחn���p���06�� @����<��I� I����B�	R�k�Kҝz��Q0$��&�2�l�3�f�[����M���'G&=ЎL��ӳs��y�IHnB�rBn�/�m����Y���A� 0�6Q�d��td����	2�\1��h�����O�D����>��~�J�~E�$E씡3�R	���'�ڋy�'^B�'W�]�7l��G:�@L	�IT��vӀ�D�;"$%����$�֘�^����I=7dLY!/�q]��3W���<a��?I����$ۙL����ǖM���S���#kn���ҤSy��˟��Io�Ky)�2u���.�q:��
���U2�%��yr�'aB�'��	s�Ti{�O�p�iQ��K��hy��9RH��O*�D�O��O(˓`�=�'�1� �17�6�F�{���b0Y���I�<�ICy�'A�/2����y��M�ix�zp��2h���X䦹�	i�Ipynބ�ا� h��g4:�5�"��x^*����i��'X�	�\M���K|�����'�.��X��+RCn0���$�Ee�'�剖}�*#<�O�(9aҋM"N�%�"�5$9�ߴ���A�5G�,m����i�O.��R~B喦-.��3�F�0��)�a���M�,Od:�i!�i>O5����'��d�D#�b� 5��iQP c�w�B���OF�$��|�&���I��q��L�5I[ЅK�l�v��B�4`B�IDx��i�O�q�%�ςW��i���!BԨc�]��%����l���gu��0H<���?�'(����%Z�<���Y ���X"�[�}BHK���'_R�'�B�֏E�� `@�N�����j\+��7��O�����MT��?qJ>�� E���\��eԲ,��'�⹑�y��'���'��ɳ4�������!�%���!W��l 4ٹ�ē�?�������d�{�J��4�˦%|���U	^(3V ��d�d�O���O���\��6��,��hߍf��)qV;n���uT�<�	��'�8�'rxm��OX��	�h|8�'�de���fT���	����vy�Z�'Q��'�?��ɨ*��4�0�6oX�pF�	?T5�F�'=�'�R�'tP�2��� �>��A0�9qOXe)Q��_����'{2^���¥_%����OH��៺<��Oj@�z�"�7ܐq��)�z�	�$��9$�b��?��O�"쀠�	Vu�q�vո	��u��4���n��@l�����Iɟ��S�������&IM�p��猴^�p)G�i��'��rF�'��':q�¨H"ύ�l�@��p�F�V-ҕR7�inԸ��sӞ�$�O��$���y�'��	y9�##��JIl�Ib��
���r�4/
j�;����Ođ9E(� )�"k�!��$Ǐ�e�Iş��I�3��ت�O ��?��'x� 7�W�m(Vb6m��v�[�}�J���'���'�����)�Q�_+ǔ]1vH|����i�R���듋��OX�Ok�;��m�����\�Q�5�U���I���&���џ ��lyra��;*��%/ĘJ9D���q����̲>�)O��$=�$�O��D�>[F������7��ܛ �W>aQ"�vG;���O`���O��n<2A�g6�5蔪�4O�8CNB�-H�زu�i�����%������t���m?A�	��b�:��0J�:n������}}��'\��'�I�}MD	B���$�� ��5�3�ֿ5P��{CE��1oZןT&���	ןH���Qܓ5��}��K
�Y�|I�4�Q�G�Eo�x��oyR�^48��?y�����A��p�s�,��S㸩��i�*��'��'A�EB��'�'/��S�RZ>5 �=����o�SO�FZ����C^��M���?	���Z}Zc�`���ڀN2����J�Gr��ڴ�?�J�Z�a�b�I�b��ph`�X qS*)�AHT�Fi���J7��Oh�$�O��ɏi}S���o��9~h�EGϞ0����㍌.�M�ZD�`�?����'������7�2�z��	h{䘡��k���d�O��dV� �Dy%�������\�=�FH�;��Ў�K�<`m���L'��������O\�$�O�=�'�M�H��@�d�K�(�@@��Ϧ��I�e�nђI<ͧ�?�M>��Ya:��$��g( тK�	��$���I@y��'��' �I%}�N�������H󠍊�+�T�i#�D����?A������jx����*hxX�F�1d�r�IU�i^�W�$�I����I^yD��>A��S������	Csd�{�\5.��?!�����4��W�x:��W2</d�����z@�$���@y��'���p1[>��	-B�!�bƆ#A��i&����bش��'��X�`��a+�DE�-�~�!���+a��&A����'j���(yq��V�d�'����5��G!�~�9�I6.�R�P���$�ē�?�)O�X�i�=����
BB8���$o-�A��&�>��tκ}���?����y�����RTB�F�	ZLD�ò�:	� �i�R[�����'�S�+_��Dk�n8,�<]��ᜩ[�6M�6N�b��O�$y��	�<�O��$�����Z��t
CK�Ѹ�j�m�>!�I�g���O���Rw�a����	��SrIY.#�x6�O����O�D�t��O�i>y��ǟ������X`nC&:R�t����Mc��?��e�T0��U?������Οd����r�(i�$�6#~0���# <�M��	����Q�x�OR�|ңܔ^oܙ�wBD�A���2O�0m��3�@������Ol�D�O�˓s�f�Cǁ�`�Z�,��V�Ġ�׎>Pr�'��'�RR���I쟰��T9���paS;j�L�Î�s�x���Fy"�'}�S����$|�����{�`1i�	T�#y� ��ӎUȝn�꟰��i���?1�}f(�؀צ��!�L��X�´N�R��H�>i���?���򄘸

�Q$>��Uj�0��E�W���L@��c @��M����?9/Op���O��0#F�O��'*`V90f�h(4���^�;f�5@�i22X���	�v��OG7O�\c"����fe�qV��.1Z��q�7��O`�̮R㬤���T?�E���I�©x��#3��M ��>����1���?q���y�����\@e*1$H�<��]�P��#�i���'F��B��Ƙ��π ތ��D�5"0��u�7[廇�i���v,d�����O����~��'n�I�$28���� 3��8�"�"U����4 ��D�'���z���?96̉&||	ᣃ�<t"�&Utw�F�'t��'2|�#��>�+O��d�����CѼ����F�\i���`�j��<�3+�<�O'��'��ˠ�Τ���ϝrm�m�	)7m�O���A��b}R����ay�5�LP=ML��T�ϕOUqѴ�B����.P�$�O����OX���O�ʓ>5,xY0FԨY m��"C$�)��ʗy`�IbyB�'��	��I��T*ĉ��������	����ŝ�c.��	~y��'���'�剒Xމ �O��x$,2At��"H=g�bI�ݴ���O���?I���?�fd��<���W����e���L�`K֐<����'���'X�W�D���ΰ��	�OVp�g�K�B��G!L����������ly��'W��'��#�'oR�O U�ɮD�	Z�עF�L�Ё�i���'���"̨��������O���Poጨ�b삿[������"E�"��'��'���͊�y2Q>�dJ%ʎ��N��e@Ia�� ��#�ݕ'��9��mp�����OL�d�B ֧u�R2�@�d\"/ �����/�MK���?�c�U~�T�(�}�6��/���1�	�
�PhL��z&���MC���?��r�S��'��KĮB3a��iB��$)�0q#}����;O�ĳ<y����'�*�I�_��@��@<$Ё�,�Z���O^���'1n��'��Iퟐ����	ǎך6���蛚(SZ9o����'� �Ø����OZ��O��kX�@n�䠄�<2G ��L��	�ɥZ�R��O���?�.O���Ƙ��Gg�O����C�!�M�[��;�Az���ݟ �I����IQy"g[�cp��8��Qj�З����3�ȯ>�*O��d�<���?���n�LA��I�f�>���AM��|Q����<q���?��?	����D
^���'.���e�".W>x0H��W�b%lZty��'Y�	��(��ߟ����P�1g� \�jQ�gG����叶���OB���O�˓d�f與S?M�� \^t2$�5`�fM�0"?N�$���4�?).O���O���!"���OT�$��,^�e��m��F(�<`T&�'X�lZ�h��Sy�Q�/��'�?A���j�͎$#��׭L{���I ��������Ο�3B{��'���'@cQ�aɫ9� %�S�[�] �	lcy��b,7M�O�D�O��i_e}Zw�]�ɑ v��3��=
��h�4�?��:x�y̓���Og�D�V�j�^0 B�<՞��ٴu,��t�i�"�'���Od����D�6��CB�J��x�C��~�l�!vs��I؟ԗ'���C�a3�W�Ax���G�1e�X�o��<�Ißs�����'�R�O����4!��I�v�:QZзi�'}$T➧���OV���?}�" �3�T�P����7��]X�r�J��0�X$�������%�֘C8B��3@�\&�!c����|������O����O��I��`�+u�x�'�Q�%�(����O|�d!�D�O~�d&�>q�� ��x����C5$F��8O&˓�?����?�,Oh�(Pb��|��Q?.��q ͬ _F��C!�C�I�&�X�	���Ɵ0�	Տ s� ��E���=�R������O����OB���l�`���#�M*�X�n��xX,I4.�v�7m�O��O��D�O�u����O��'��H�k͕.w$-hpb�D���4�?!�����kt$>�	�?	 ��cx�í�Vl���
�ē�?��|��[��䓕���Q5G����(T��
�)�M�*O�l���Y��Y�������l��'K��%� HQ�Q��!F��|3ڴ�?	���bQ;��䓪�O���ŏ^v�a�P1Bm�A	�4W�VU���i)B�'Q��Ohxc����f�tJ���ь�8��x��#�M;�K�<O>�����'b�i��.�  �2�i�Q�i�moӾ�$�O:�$�?�F�%�`�	���C~r%*�@�-N&�5����[� imn̓o��	�J|:���?��O��0��j�k�bh���Y
cʮ�:ߴ�?���lb����l�i��)���N*�s!����J�z2ɦ>yS����?�.O&�D�O��D�</6��-�B�<	��[T�Ս{�j׍a}�P�X��ay��'�r�'ބ���d&�DES��Z6*��q� �yR�'��'q��'��(5|�Z�O"�9���`R����08>�;ߴ���O8��?q���?�WA	�<sB߅b��9U��M��I�V돫+�v�'�2�'��Q��Ȗi�����O�A �Đ�rN���͝$݆�I!a�Ǧ��	My"�'�b�'͘�
�'F�s�l͑�BY�3RbyB�ٔF��g�i7��'C�E���[������OT�I 
mR���
 �����5KI�?~d)�'��'K��y��'�b�'��I"F���&�ȥb'�<�GʥI��VT��Y��Y,�M����?���JW��]�7E��Cb(��a�:d}�7��O>�$V{��/�$,��V�� s�i0*�P�/D�j��6M�8Bo��mZ�����h�����$�<��F�(�Vd#�e��g�L��
�2d�Ý��y|"���O�D�ђF;r �jX�/Y�H�ϋ֦���̟�	����ʪOrʓ�?��'��=�`l��Sr8Up͜�KEPڴ��C1�t�S���'���'N,� &���-	4�9�՝kE�m���i��7�~���d�O�˓�?����!qMG�<r|;WW#C���'�4`�'�2�'1b�'}�[�H�I�=g�<P4o�0i~<��D��E�v=hN<����?�����d�O���@�p�F�1P$�U>��z�˥z��F��O0�D�<���o�6y+�O	B,�ǆа �U	�fìH�����4���OF�O����O$��J["{ޛ&2^-��xV
�(�:X[ą���d�O�$�O��O�Х�7��䌗
iw�H��7Kh��FOL6{`6��OX�O8���Od�;a��M�N	�qFXNP�귂M8u �V�'y�Y��y)��ħ�?��'E��]9!�V�,�Pdi�(*�
'�x��';b%C��O��Ik��`!o�6Eʎ䱣�W�j鴓OrP0�X�Q�X��D�v��E�^7�"!	��!��R8"��% �*T�>|u��� �8�K�_��dYx�BU T�0��
Q�2���(�Ȑ�	,�┍�<�HU�s�� ���9	��_]d�hkP"CĒ�aU�([��Ԍ�>u����V�����Ku4(�iU,_���q�l�����!g���}�D��,Zpdx�)�րL����!ȁG΂���O����O�D�;�?���;����7�m!�d
�T�Z�ɀ�ʶ�8��ҞE*�4C�	X�s�I&}J�@c����@G
&G����4u+jܳ�$�D{��H""��^y�J�ր�V�s����'NC���)���I��F{B[�lb+�,T�[�!L��4�&D���4F�	�A
(Q����_�HO��Vy��D��6͒y�}2��%>FtU���^�,P���O��D�O�m ��O��$f>���ep�A�vj�q�"��,;:�T餏�KC��ۓ�� �oL/�|��
_�h7H`�eDF[��³N2V�a{k޳�?���`���C	�.��)�0oS*v�b=���d>��L�q��@�'ۄ I"���"D��C�FX����g�D?f�
T'l�Hz�O��;N���\����t���^T#
�`l�>R]�����2X\B%�'�"�'�t�#M>D\�i�2K���T>ݠ����4�ޑ�ae� D�X��g(�unx�c�_��N��C��ħhVp*�NT�a!De�Dy��р�?����Omƍ�p-	��:U取�8��'��"�3{�1@�
E��!��ސ�0>�җxB���
3��±#!Bx��BP���y��29R��?i(�F��C�O:���O��9� V"H=�fݾ�%������&@Y*?'U����ʧҘ�?�`�T��Z����_�fGY;�d����2hh9����%P�S��?х�E�Xz%($���z,����)]�Xĳ���?9�O�O��'h���͙�]�^9eA�W^D�z�'�Yk�!�#]^�5iuC��%Y�+���}����W>#�Q�f����pL���ޅlb����O����JD�f\��$�Od���OtH�O��iZ)e�y��(0E�\9`�L�l3U/���Rd�̝ ��Q��O���<�q˕7f�l �Q͸x�p1�"=Ҟ�*�Ɖ(�4���";uȡ��QWQ�t	��T;%�> 3��tb�$��+ן�[B����0�I���<)����D�t$��F�U�T(R���/�!�d\�bR���F"FMN����b�8�Dzʟ�ʓ(h�
�i�<���Z"}S$5s$ 
6Xf}w�'�Z6�&�'����'�B1�� �O�Q��6��R��P�Ñ�>0�8Uf�+��|�時\d�$��i3��!ȕId�h3��)����
�r�����՟B�ܕ3����v��5U��+Q���X�INy��'��O��� �t�C�H�&x:���W�0��B�	=�������/�<�0�ǒ�`�\�����<i!�5?���'�R>%�/� ��2�B_�#�`D.�9���d�ɺb����C�S�Djٓd���w!�	�ljdAL��(OB��`��ZD֍���pX��@BE���<q������ޟ���X���C]��b�F^�MζX	Q�N*NB��s�\s��������T�P5�&�O�Y%�8Sֆ>Q1T c*ۘv6@�%�؟\��I�#FB���D�;.��I�� �9VG�C�	��|%@��9�jM�&̆
��C�I�)�U,*�l�(	#6W�C�	
E/�A[��j�>LgG{�B�	oe���Ī�,�lcp-|�B�ɺm	��h@�[�V�\1D.�{�nB��N���)���yL�a2��GATB�I�bi`Ԓ�Ƀ�E'�dʃcY2��C�ɔi(��Ӄm�:1/ �Ó���V0�C�IkkV ˤ�ImQ"1�V��C�)� �t{dKG%bGp�36gʭ�@t�"O�QQh��P��Ÿk�d"O����&B�4�b��6_�]�"O����͒	D�a�K����1b"ON9�Q�܄S�n �e�*�^i+""Opu{���-Jq�XJ� �k�"Oz��'��
]��3��X��I{�"O*5�u�Y��T�E4y�����"Ota���:|��%�fR�.ظp[�"O�X��/�7"|�U�U�
�e�i"O
"Dj֓.�G +y�<�f"O:x�aɎ&f��{�� [~��"O����
Y]�2&��@?\E�"O��!�O����9۠n�2b�u�E"O,E���Ԕ9.@@k����Y_0�9�"O����HE=a�h�2aQ[�����"O<�$Q�M���H���?����"O:�0k/MT���H������"O�w�"�PQ�W"����"OBi@DG׎��c�e��T�"O��`�fK�)��h��䑈���"OP�8�R i/�,bs�E#<||��"ON���Ŷ^ln�į�B�˙%!��D�.Dj��R)r�̵�!h�\!�d^kAf�q�Ac lٳ��f�!�Bb�|�r�D�kX�)D^\�!�d�k���ŠPޕ)�c ]�!��ʾ>C>Y�6h��eg�t�2�ř\�!�$G���0�OXf��u臠�!��{"�����Id�~=��GC��!���ļ+�f�	Lj���@�В!!�D jʘ �+
~6}��EF�M�!��;R�8���F�7[z�H�<+C!���x}�eH_����ߛA!�D�<N4pIb��nq� )����c!�D�'�.<��,-jZm�A��(\!�O�/W$9�'䖆ne <rbNE�!?!��1���ǀ��-\&P�S���!�D���ޠ��蔰AB&�����9j!�^�t��*�̈=XFz��`���8!�D%k���"�jŕJ�,�g�&3}!���gi��TG�1E�Q񆁨6c!��	K
B� �Z6':��X��K�K�!�D-��m�3�U8lHV��}�!�D4bQ2A�1CO�T���%�b�!򤆍n��A3�!
;$dq��/߃3!���-0m�5�e���:��"��2�!�D
"��xz��ӄ	�^����-*�'vJ���
#T�t1E�M,~���'�}����9��0ԧA�'���
�'�:�d��	r��KF
�L@�'/~l�a+7�Lu��h�Cz��
�'�T ��S�ht`�#炛Q���	�'���xcL*I�Z���9~�D��'$� H�ˌ�2����uJ�-�	�'N>u��� %_�c"�=���j	�'�U��Qzyz�i�R(H���*� 	�'G/C�651�B�'c����p��'IO�&(�x�b�$yj�	���I�U��!��|2��8h��ʖ��y���s ���槿�5�]�^4�p�R��u���l�k�e�	ju�X��:]@��õ^��1�`Z�ɱ"�pl鑄�T���;2�6-���FV�By
��ؐ#X��r��\;(�[�鞑:���kUb�Pg��³�R���'�p�z��� Hy�D��鞓V�Z��T9���?#������2F�&ǃ�"�1VbH��3� )��o�`J��6//��=x�P���r�|�'����A� 	^F�㞭+��K�#�1�T��mD<��ظ������O��7�x��l�<'g@S�kZ���g��j�V�3
�n�Փ��f���q!/R���(Mݦ]�Ąx���Ȋ�c̛^w���������5mG��3g�ey�띓v�hU���"������(ز ���saA�aY%��r�_������)�~��z�N��P+D�W8<����
�"]#vݟ��n���A�U�h7̰PKĚQJ��Dx2B�[\n��f�HY~�#�(���?�'#H7��a�xx��X�"�\m��$1~�򁗇P�(v��c��>	��B8i����ABg��M�� �*��n9,�$5r��aP����?c���&�0��NF<tQ4�t���h&�3kk�~��YLL�p��	�@��3� K//}�T�=1���:F�@ ��Iyb�Q���!�5+[�Q�lB,K�l��G�%g�z��E����0LٹTW�mc�i��4z����J�X@��W7b�vX'O@�J����']�d��)�>u:���.6C����'����LԖxob����ŁK��$c�{��Ѕ>ؒ�	4�Χ'"��y�����r��:�m\�TzT1si�!"��	�gR��!OD2w��&(�2c��>���ͺG6,}`�m,#��}q�H\(Oܭy`��'[��0��7��'��йfꐺT�.�3킵2��x��Ux������S.Y)'��W��:�i�w��PfH�FJft0$D����')Q��]�k��+Ofu2 L|�eN��P�Xp��Bw_v	o���=q�m��q� �F���@�J��Ƈ �ea�)�;������0�z\H�aX��2�!��)Ф%�hH��Юp��d��b��E�B!I�R~���&A+��O�%�f�$5E�Љ&�R�x���rU�>�%b�*c��}��(Y1`����M��p�fͅ;�4����I[,�!j7��2d�ضue�����H�vA�"S0΀lYS�٘>�L���a'�IR.�e�0�*��Ĳ���~u[���X��%i��V+������'|T����L�Aش�%bd��"�OU�]��'l�bAOT�Y��8�,O��ӷ�t�����P��<( ���T�v�7�Or�P��ʝ� ���@29K�8P���Rs$=�u�ݭH�3d�4J�j-O^#�D޲q��j��<	�n{s�O <�a�(2"��sK��XLj�9��	H�bÃ ��H��P"+��N�	�}@���@��u�䫈AZ����2d�
 I�!J6���-�=�Q�������y�)F�Ay�aH/d�`�)�gb��o�pB����-?� �H���M�� �8�j7ʃ+-����\*[�nF�ӈ6#<��D,Q�$�aG�ʗ� M:��
�[�d�1E�<6d�}��	k�nX̻9�詡���f��H ��r���	�yd��#L�?�<�i`hW�,�
PP�'
X�'�H���_��� �B����'6� �bO4jj��7��/l�P��5P��Kv��8?��Aa膭~��m�Q"�"�J<�5�Y`�<s�O�O�+f��3�$"��z4m�U��=+.{��\!&����I>h*�O���YA�*�ӯO
0�H>YuIݑ�2`�~�B��$�G����Ș��p?)e�E�{U���Kի&j�(�F~q0�*۝������
��[p�͓|���P���Ơ-y����a
B j�/KlfU�f"O41�$#� �n���U�b��`K�
�R���i1ָ�Wd�Ol�[������D\�V: H�1��p���Cd�E'!�9��I�D�zR��(ITs\�9W�4>J��s(E�eC1����O��禖T��������p�O����D*O 8p�@L���O��R�B�t`�}#-E�24 ���6Z`���$�Wh<A��@X���14�>P0!�m�& �D��]60���h�$ RR(�R� }�Frޑ(ǍMW�ZS��  2���2�5�O�,3Ţ52���q%LY"d��1��mΓ%lT��]=J� �#.]�:��	��i��8B��y�.)��j�� �a*^�ct���3�/&�f)�O�x¯�}�>	�qb���u�j��qW#�.��v Ņ
��y���JI}riݕC�.U�3�Cmx��bdK˯O�P�X��ce��6��� ��q�� �)O��r뛤o����&���'tc�ʍ�?U�%��(�${Q����K�~i��C������I�ͪE$Ñg��uz�\��aOb��=A��#?a�,�L���	:��<��A���UIF�Z��L"��:	Ny9DKң,��'���d5�O���h�CH	{~�թ��1K1d4�'=ze0�^lb�������O����O���N�>:Qq�H �'�V-XBL���/J&_��B ѳ?+z�M?˓5��Q`N�D��LĢ��b����K�e֔!�:H2Eh�	Fh��+�(O.L�p`Z99���b"�׽@�p� ��J������b�ɵ	ԎMj��	���M?���@��@���ܿ\N��#A�����$�1u}X�B��w!jP�7�TP��W�ni�ȓ0�'��x!K�I!����l?�O�|���I���D���J�-��)`�L�.���+W�ħK�$� J��0���Q6���v�^\�I��J��aQjO~d(���,,����v4�E�ھ[K���⓽
{�`SfW#��칱�>Q0N�'��%Ʉ��,~�u�D�Ekt�9�H�غ��A@
�|�S4F�g��	�-B�P����rP�ѵ#��'�Dk�!��j5����g�+=���t�\�F��8�R�,j��x
� *Q+���*�,�H�
��DΚHSe��"z:M�"̓���D��*
��6��$/n��>�8�j� }]j��7_��MYԊ��c-a{b�N�mJ��ݾt�J`� �^C"��w�Ռ+0IlZ��$��o@�.������8�^��
��4JasW��#,� J�Nڬ9�R)�C
XZ�'�kF�p� H�Fʌy0R(�GH:7E8���͵_b$� `�LST�-�`H�r~�ʉ�(�Z�̀$%q\���C��P����e��M��A�Bk�P����M�3�( �(���M5�H$b̴zc� ��1�@)��@��v�DMV�=ntIGJ�Z�%�Cb.TdTۧ�V�4$� ���;Ir�ٙ�E˽'��Iq�76�� �)��?ٛ�M۝gQ�Hs��/w�6�]�F�A� L�������	z����'UdM�g��o	8���ӥՌ�U�H�x��'�Z�*TFK%!(�G�;^&����d@:��)�s��=�����T:7Ѡ4�R�Q��@7}�z�#$=?�r�̜L��	�K��Rͽn�����RF�"�Łi炴h�m�|[��%m��a�\�r&X�V\�Yó�Q�S��w\V�s�	�L�&l���+����'�L��t���,T�V�b����QÔ�L
�����0�l+��<�����F��2#�?��!3�$�[a|���g)������E�U;�M�e��d���$J<�T"A�s]�����&�[V�S�;ĭk�˃��ΘGx�h�93�V|c��D�B�.�YӦ�g�iH=��4�6�cT\1�!��8O6�	[�i	�ݞ�y��� >
��`��5�q{��ٽwm���s�Ȑ4���=Q���`�M�5  	4D�l"��<|�,AѥKd���¢L����3��2Tݺ�BFlJ��3�7O��p5.�_��qC`QH'>��I�� ��`�ݳ.� d���I-p'�� �N�g�Z��R&:(�Մ��?L�왰��c���t���rC�I�f'��x�(1�܈C"OF,TC�I(��8�❂<���A�6%�C�I�fZ(�hBdE!4H\���O�-��C�	#5!Fl�3'�L3Ri����dC��7c`�����,~.E�V)��.C�i����՟:dc�^vHJd"O����ECs����7W���"O���n�5���C�U�($�e�3"O��n�+_�P@D@�.w�X�"O��$aL�*���B��6�(�{"O #�j�B���ԏB��`��"O|	�(-�H�sf�VJ6���2"O�H���W,R�-���C+D�\�4"O���c��g#:�"g�l%j��0"O�2'�� ����Z�(�A��"ODE��V^9̬� �q�8��"OZap�-���pm�L���"O��!�o�Tj��!� |{����"OB[�M��D����4K@�O���2"OrMٲeY�-E҉�D�֙=BZ���"O�v���v�<�O	$�	�!"O��7�0�\�7�	SpYAq"O��I���;7���̕Z�x�%"OiH�(�� ��\)@�ژ1x:��"Od-z�FH	�e�u"X�a��L8�"Ot�Qa)R��@���$��8��"OЛu�^P>��Ї
�4l}R�`�"O
�R��ХIRr93����I`���"O��a6LF�_����v�A&����s"O:���h��)&� ���/n�ܴ�"Ob�07"�3L�ެ8�E0p��L��"OlX�Ԡ���\�9��D�v�N���"O��&L�a�F�[A�^�Y�,�&"O8|*�iY��Y��� �}3�Ś�"O�������,m���U?'��i"Ot zA���y�x���/�?^�"Oȓ��Ĺrw0����C�~���"OH	���1<4�X�E��:f"O��ɒ��D���7�%/�����"O� �͉w��8k��І��"�(�R"O\l��%P�q;���!�̨x�Ht �"O��M�s�6� ��F9D��K�a�1�4��$
H�L�&�,D���t)_����8"��J_"ā��.D�,�DN
H�&%
�HΧD[�=�`�*D�dr��Ye�ZL[b�͆(�
uk@�)D��K�K�aK�������y�iQ�b)D�l`7�Β$�-��G��0�6��@3D���"��pw0,��ʕ9w! H�U�<D����K���8xZ��Q0{��Y7�=D��13�![_�%@�#�8�rݑ�g;D��j�I_j�JA�'��������:D��y��ƑK��9�5�^��9D�`�#ӯ�XQfOY#5x�S6<D�xS��:���Di��C�,!���.D�8���y��qHkЭi� �Rs�)D�,2��2�d��񈒢Mj
 R+D��0������1��0~�$��(D��Ps%C�/|8!3Ƙ+َT���%D���/�
�&m����%*&Y�4�$D��3��Q9eS�)'*Ϸ��0� �#D��(#M18o�Pk�ΏN�p����=D�����}S�rCD�f�>��C�7D�@��Fؗ8��aN�e� ���5D���֭�:>�9�V&�mA8I��o9D�h�5J�)~F��6F_4>>8��9D�8��6e����%X��a�ש8D�(�1�[��v���4w�~�r#�:D�$a�I�"�X1�Zk��jEJ8D��)3�Z�����1g)�F6D�0Ӥ�~�@h��q�ؔc5D�hC��	�O�̀���.C�`��.6D�d ��;>���A�-��IK@��E!D����gͮpVxJd�([cP��q�?D��3+�hX�(���4�"�@>D�| ��	t�M�$��u��UC#�;D������"".2�H4��S�(���9D�冐����w$
;DhP���<D�<s�.��~�,�����xܚD�:D�����ʖS��郥��n.JX#�8D�Ā�Γ-e��R� ��5Yl����9D�HK�MRbU���A�[U(���b7D�H��V�[��%���2Ј��5D�$a6�
u��hŧQ*GIj�bbJ>D�(�)-�p��R�ۛ8�
Y+��'D�l�h�!IW�5���Ka��t���*D�ؘ�D�65�piB�IV�k��� ��)D�,:g,����ճ�cO2d�xXې�&D��� ��.Q
DZ"�N�1l4ءd1D��90��K�/̶AK(��B<D���5��G�.�b ��F�Mi �:D� H@�]*�Q��E:W�Z���9D�hi�l^92`���ղ!v����<D� ;R�5:[��Ф�P*~���/D�l����m�j4�p��5D��P�),D�a�mQ�C�r��Kz���r4�(D�L
��Ě`N|�sU�̝`�&��*O��:A/��T�bA��s��Q""Oص��#�O�-��훱T��)x�"Ob���E����2�˭a�qd"O< ��앑hv��C��E$v�h6"Ojd���Y;10�@:�N�kx"Y�"O���a@:3hT[�ß�2�T�iF"O� ���߸0|4Q0cV���+4"O&J	�Iظ4�� ��G5BD"OJYc����,pwO�"l�#�"O ���ƚ�S%�HJu��9��P"O�]��#OK��  hɗ ��C"O��R��yк�R��1���г"O�iaf��\�F�#w�?]��-�b"O���6�Ŵn,���ݴ�Ր!"O^��3�P��Έ�'�L>]����"O�m���I@m"T/�2l���V"O:%�S��'��&��+3�|q"O"-RD�ΕM��I�,�!&����"O�uK�/ߴw@,����;BZ�"O2��g� *�Đ�\�{�py"O�r�O�F�� �é�.��"Ox�� �\)``���3N�!�"O���.0G^< ��
Pj�`"O���f�Cy�l��)'e�٫�"Oॠp��$V��&%[LD�@0"O�`��0K�j��ŧAD���U"O�l������Qt-#['
�"O怊��~ܺ8����sh��W"Oޜ��o� j]�P��v����"O�T�� �*K��!�T�I�@�"O��bJ�KT4٠hӘ�n���"OP��W��JbtZE'�"9��l�"O��K� /I8�`&F�D3*�X�"O� 3w�	-[�NY�vŊ�e5Ԅ�W�%4�H)%�	�x���B
������?D�\1�h˒ ��P��fH-&���5#>D��qH��s(���3h��-KV�;D�pP�M?H�TB��ĭ!�}��$6D��(7dQS�2 Ap(H�Z�l�8��0D�T��nޣ5T�(Z'j�71!���1D��qg��<a�� ҥ�U��Lz "$D��d�6z�t�j�n�Sj��Z�8D���b�ȫ>�jA�����T�Rt�7D����	��ҩ���"@Y� ��6D��R� H/-Cli@��c��6D��s'01+ʬ�6&T	z��XC &D�L����#"������eŸ��g�"\O�b��i�ꑕt�d�qR�	}�Y���#D���e�)6�D�l���1W� D��K7O�� A�-����'�`=��l=D� �%T��4,AQ�DsZ�Q�(=D�C�i=�Bu�4,֨Eo�����6D���1�˲W^�%h1�@�6�VA*"*O� ����eR(B"�z�(�A"O��iU��!i�4`Cn��W�02"O���R�T4 �n(�3g͆d[�!4"O�m�P��8_��1i�&�Jv��"Ov��
y�"��E�bEBu�g"O����@�j]��`����:(�y�"OX��DF�@���B�+<��"OVL��厸~�|��ƷG}�\����)|OB���c
�$0&��7 �%f��"O.Q:)�E��-Y �J�g"O:�����;Z� ��@�?0���"O��D���� ��CO
VBL��"O$�`Ԇʀ6���-)I1(�"O��ǧݎ �|e����'��PY0"OX!����F��.�0�޵@�"O~�6�G��H�u�T���3"O"�⋅4;(��EhH������"O� �U��K3������W�^�(�1"O �kv�05����"�*~�R�@-�S��y���Q�]�V���6sfk�8�yK�U��=0V�Ȋ�����y�B+1���'�WӲ9P��؆�y����9#����Ƭx��Ł�j��y��i�dj�*ߣ ��h[��yb��1,T<�4� B�`�XAƉ��y��!�X-4/��9/�M� L�5���.�S�OuBe����4#�R�kP1
`�dx�'=e5�V3Qo �r��ӈ+����'�0���@�2I�HL�#+G�(�
�'�`)B��c�~倓KF�tL��
�'���Wlѻa!�@{S��j�Vy
�'��4��wd����i��e��l��'�|@ �NE�r�Ha�f��=+��m:�'��zЀ�b��h�3A�� ��Y�'j�8{�Q1j5��".u�\j
�'$�����^��1H �&p���AB!�S��?�df۴5�$��o-Y�h�D�<���^O�8��3�̌[;�T� ��H�<�� 0�$Sqo��;U| ��@X�lDy�*4�j�0 ��b��u�R��y��).�h���
����4O���yRM3Fm�d�Rl*����yr�<��j�#e.\®�y��LP��Q'!Ɍ�lB6�yr�� �=���T)d�����
��y��V�..:�H�K\<j �S��yBBQ�(�V9[�LG����$�?�y�'��egP!���	�Ή:��N*�yBc�>2���h�+�#��x�矇�y�fFq�(�����Pʶ|Rs��yR��3E���tǆ�����r���y�7��4�%E��C)��p2�E��yrǏ1���Ц��8|����Y��y"�}�)�&�Qf˼A�W���y�\�����DOan�!˚
�y2cĿ#�������N�.�iB=�y�IӸ%�0�Xd�Y�H��(
�����yr.�4x,ɇ �9:
Qh
��y�H�;W�������06 �\TcT<�y2D�l?D	IdT�%}p���N'�y��� q��:����|�]!#�2�y2�J3�ji 4���������y���r�ԭ!4��!
	(q���Py�N�X3��"3�L�g��%Ƞ��t�<	v�Y X�����Juvx��r�<��b�'jzhQ���
��ez���y�<1VDA1l�����17�4��2/a�<Y�j�L��fIJ�57@�����\�<��
�;vH)��_�h����P�<���.Zrh��3�hƴ��IW�<�'E]/�89J��j^F`�
T�<i��π;�Ji����/	 (yӭ�Q�<a��(B6T���P=B��0Ҫ�I�<Q��U� ,P���G�;��b6�B�<A���!J��)�ch����̕{�<�G�T�(�ꗘr�։a��BO�<y�A���U�B
�|��8�@H�<16A�)yN�QB���s0j}���Q@�<�aX�On��
v��8gm�{�<!6oVYvR\�ע��6v��跇�^�<A���;,a`I� J�^�愐u#�T�<� ��y �TR��P+h���"O��B���,+�
�ckŝ
����g"O�h���R�;��� �O9m����B"O�nN�[̴��g��H4�aO'D��;n�h��B�B�d_N�
��:D�p ��^�S*�A�e��|-��39D�h���%<���s�����R�1D�s1	߇>�!+��j�H�+u!1D�`�B��t�`*Z�<�
v�3D�� �mƷ\���8�!�##@u��`4D� �u	ڷG�L��pd-`H��p�%T��ä\�:?��(��H=�� �"O��Z��ҤE
<	14����� "O���a�. ���$�kV"OJ��g��7J�T�I�މs���*�"O�1zG��H9��$m�p
B��+�y�!RG��y�)��iy4�S�����yr�Ƈ�<]a#��Z��k�)Z<�yr���_��xP�"�6|���7��yB�NK "�щ7w!#7j�/�y"�G�{�����@�ly�L��"�4�y�,"ga��s(΁8�iavğ!�y2e�	qb�b���23̐�%ج�y⏗撑� c�(;��u(%CB��y2�	�`�,L
B��8< 94�S��yB�D��m�R��(Z���"�D�y�`�2}�p�*L�<&k����I�y�&њOQ��y.����U��yRD
�xA��!��- �Y��Lɛ�y�N5|�c
O>~e�=y0b��y"��re�P�G�3#����W�`�y�œ�Z�U��.�B�[�f�����'Bzt3p(غ{�p8�QDȭ^7�<H�'�����-�%f�re �.A�q��'c��ӤB�^����Ѐ}�I@�'y
i�T�~)��K�x�=��'����s�]5T� �;�Mߝ�����'�(���i�>D���bP`?: 5!�'�[R&Xt�����S��@��
�'w��8�;t����y���@
�'"���g�� X��)���?3>��'|�� ��+n^�K@J�'��<��'�t� ��E����)�4��{�'9$m*6�W�{~9�nP� \�P�
�'�4���{H&���B�:gl����'���
ўX��]�eBE�����'Z��ql�0��Y ��]��@h��'�V���e�|�p��F`@i,�*�'�b��C d4��W�x^~5�
�'�zx�T��+�@8�B��	�
d�
�'"�T�C�Ѯ
�8I��Kԅg�ԍ�
�'��A(Q�];_�!��C�ٚ
�'�i�� ȴT��)����0@P�'�.i���ȜJ��̢~ۄi�ʓ+�����A�O!��ԄD<z[,ɇȓv=����5h�X���ȓ>AX��k�7+��p٠*��&�bɆ�@��d��K_?�K�K�t͸�%2D�xs��>iJ�QE >3�LK�b4T����r>T��蕌��Q��"O��3���mG���c'��EL�A"O.���+�)	p�2`�?	$�T�7"O����׸M8��P�OO�jN��"OA;!$ʕl�)�Wo��_�X��"O� xR�l�=��	`�98��t�5"O�E��O8&���� a� ��I�"OX���V-���z�iϜ?�f��"O�	sꇨIZ��BO�<R��-;t"O��6� Us�E����b��0P"Ouʑ��^T�j��>s�HT�"O,���%R]���å�e��I�6"O0����)�t�ID�}:��"O��S� B-��w�^!^�J]�R"O&A`���xۄ���S�R��"O��T�J7�����[�l�nqr"Of �w��� Θ|�C
uҘ�{�"O�a�7N�	l儜�B)]/R�,գ�"O�)��B�@|��W��4�@ѻ"O&M3 �8e��4Ђ�֦^��1�F"Oj�0�逪pMrt�Ď��U��Q��"ON ��"Q�g��d���9V��|P�"Ov�(��٤<��#�У����"O��c�e�Y��*�
>N���
""O���u���[��M�bCǌ�4��"O�D3��2 ��9	�[�(2�[�"OZ�1��*t��pb!�.p����"O�ؙ��N/)�f��͒Q���"Of�ٱė%�x�32���r���"O���ANb��(�Y0��JP"Oi@�����=˓δ}����"O%a �̤4��S�̝$��xQ�"O~A���'������z����@"O��� !�J��Ƀkm|��ٕ"OH��P��xi�xȱ��4r>��5"O�ջ&�� ��d��]d��'�Ƞ	w�
>䬄��L�:�$�J�'�<�#��D�a���@#��(�'q��5�ԍ!�XMCÈ҈C��	�'�؛�Ҕ'~|�sw�N��Y�'���Q�S�(� ��7aD$F�(�	�'�T�����Ya���4!2=��'@�P���8u-x��w��v���r�'�N�ك)�7ɮ�f+L+~����'�
X�➗u̥��"��q'��y�'fHũ�+�?�أ���\��+�'�шu� l�h̕8PPR�C�'vޱ@��ܰ=�~�x�@�A�nPA�'�J��u��h�"�
w*N�P�03�'~��{��%�����ڳD���'�U����a�`<�EK��;���q�'�>�1ʚ��蜘�)E�7/�k�'qj+f#E{����4l�z�$��'�:!b���$��9��X�g�<�Z	�'ɲС�t`8�R�ü]�(�	�'Ȇl{!B
��ę�!ТZXJ�9�'�b�u���d�.e��%¹b��t*�'�����g�(�YFmț���'`d@p���1)3�d��
�
Rl��'#,�*���x�<��u�Y��b��'��(��u�9�8ՙQ���"�C���U7!Su�,aDݻj��I�
�'���e	U�!XS@!:�4]r�'��aY�	�I2L�r�9,8�'L�@u�E
x��ɨeA_��h|��x3��H#�-���$G[)RWv���/���
�U�|�#A���zL�ȓN�Na�Q�^�00�f���1��L��i� N�ys
���FG9�R��S�? �ڵ��9A�tޚ{�Lm�u"O$� �%�& (�f�7����"O��V��[%Di��X�0�ʰ��"O��5�ؘgi�c�O�,�*��3"O���Aa��]�j��G�A&#�&"O4��7+��M��rD�J�V)I�"O"�;��H��@i�#�wLBx�S"Ot� G��%Qn q��(:!�"O��Cg��S
��X��=@�H���"O�Eᥨ��CM��;,D���6"O.D(ĉ*�1x� �A0
�"O,"���2�(�u��qo>��$"Ozuk7i��" FHp�	ҝNh�Y�u"OtH��� ��M	WH��v�	06"Op����/B��Z1AE�8�YB"OD��`gͻ,i<9� �8B��y�"Oj-+fE��s�V�"��̈́P ���"Od �wa΢D!j��%/�1?��X!"O\����AT�ic��Z;8b]P�^�t���00�i�VN�2X!̱�]ll�?i��)�)p����'�S�t�ؽ��OA�o*!���h� �p�j��"k�}�Ą4:�!�D˝z��+�ԆxU��*�e��r;!�E/[�;��	�B-�ˍ�B!�d �k�Aس��]y��t�L�T!�țJ�4�+�9b`��Z���GJb�'�a~�똦[�"�#Gdҡ.�px�%����hOq��S뀂7���Y f�k��u�S"O:�Y2mJ*&��1J� 'h�x�"O`U`Ԩ@��|@�r
^l^UHT"O�Aӥ�?ur�ejաՀ���"O.��%G�#�(���Ӣg�:�s"O�X"D�J�>2lHR�	 +ݞt8"O�\(dM�)@�f�	�.�o�QaW��G{��霚�h��%R
ݺ�b FԊ2�!��L�lѻ#ڃ3�`�٧��}!��ċ���օYě�@X<cZ�B�I�i�`(S��>8���J�/+Y�C�	�]�h4�`-�$5��0+�>�4C䉰X�R\��i��O-l�7�ǵS9�B�,g�A3�L�(A�@��l�2�B��tLp�����0���ňA��B�I�L\[��Y"�Ȑ@-V/��B�	�\z*Պ��Њh� T�~B�ɨgA�p�Щ����0�5 �(C�I�[K^ �2��;h�r�(��^�[�0B��;�j`v��(�Fuz5�|ɠ@"O� #b�І3��ʳ��S������:�S��ݏq�$��Ď\=d�3�L �!�ߛP��	�V���hF��K'��%n!�dׄ+t�k��L* *t��ʕ^�!�$	�"!x�d�0��4d m�!�=Y�e�p����l)3B�8q�!�DF�]�m+�l���������WQ!��/1:��8�*\����M�0�'�ў�>IsBFH�7�B���ާzʝ�Qj6D����'�?@R��^�r V��� D��Z%	�gL$��j�<��-Ѓ� D�ț�GEp�I��\�SE\)c1D�Hx����(p�4r��؊
 ]S�+D�P����;7�R|����4 �1&"-D�8�
K�rnB�r'��,�胩6D��:v�2I���億'\�TJ4D�LK�*C�����M�?Q��C��%D�� �uU+�n�͸�X4W�H�"Oʌ� �$�|�8ե��jeh"O�C�ˇ�En�k!
9�ɺ�"Opi�� ����I�TI�;9?�m"�"O�}��l�Jq�d�BR/x
h�r�[��D{��נ~Y0̢��}	�� ڇ7�!��L�.|h��* �JU�p�J�dg!򄜍y#�-��ŊI|�9�'	�jm!�$ԓzWؐ�B�3Ӭ�I��
�!�d�j��d��aݚђع��ت.�!�d�0'sȔ�&�P�k�@ӗg�
f�ўԇ��O3�q��e�/,�bMN�y�lC�I�20XQq-S"� � ��/LC��/y��1�n�1gof9d�޾Te0C�ɅC�
�L�f�"<���6*OAk��7��ma�C�E�X���"O�mYv%�	T�r�ذ(ӥ��u"�"O��K���p8a�#��b=p|����ٟxE�ꀵH���i-:��S�̕��y"`W9��DDJ�7��E�P��yBlS0
0%��CI�&P|�Z!�
�y�	ѧ3;4�(�F��"GЙ�����ȓ~=d�q�N�J��P��N�AA��ȓS�±�ņ�B� u��(m����Y�(ѹ�v܁a��yÒ}�ȓ:5@q$��A�zT�î�D�a���f(�KK�m�R����V'e�y��2Ъ��VJҮ�2�9�$�)�Nu��2h����H^m�}�쐉52�M�ȓt��t�E ME�\���N�fɄ�?����T�;u&���Z�Y�����[g�i1d
F������@3Ř=��5�R�p�2���b��������dbP ĥ�%���U�sa�x��0��Yh�E����OT9ji����B���bH�[-:d����9`� �ȓ_Ila��_-}f|�����.y��Ky�1"�˕M���M�vB��ȓB3�Ē%��<\O�]��Iݝ\�$�X��M�Sܧ��Рp/�D+jY3��Gb�ʼ��Iu�'[@U�϶�B�(����h��t�ȓZ}pTx2�0@>�p���ۛn�TЇȓ;���[#��ao.��3�@��@��ȓA��kȮH��e���T�p�H܆ȓ;V��ˆ��X�b���ã}���?0L��+!�d$�$��H��D{�Q�pD�4G��a�ؽQ�J*C�4= � ��y���xvH��#�$Lo& �S�T��y�L�KYvY����B���A)��yn��4��lx��C <��QS�̻�yb�4K��0��� /$1h5@��yҮ�Kdڬ
��S=u(���C���y"��'��%j�E3f�Dx���M:�yb�Q�}�j�f-�[tr͸������hOq�\df�U��@�#��ӃP�d��"Ot�a�E "�|���O
�����w"O�I#t���","�+̾;n�@'"O���!O�)fA�d�B��1)T�IJ�"O��fg]�R��t�@�i<��S�"O�����m���X�@:\0<��"O�ۃᚑR���b���ix ���"O���?�:�p�&t�r"O�R�O=B|	!mВI�М��"ODO��I�J¬P8P�f��0E�C�)� � ���
�4�����DD����"O&�r��� d�18c ��%+���"O��hѵ"��i2 Ϙ(!�4�(7"O��V�^��pp@�?=�b=�4"O�L�������OM���L
P"O4((�x���N�'x�0P�"ON��Ӥ�+"�L��M˵X�1�"O<��F�5Sx�	I"l��-0x���"O�
5�X�ljn�h4J�9U��I��"O�(Pw�Y�.�ʜ��>���R�"O,r��] 6< ��Y,l���"O|e	GM��5�J'6���2g"O�I(a#ڮtJP�y��C� �k�"O4Q�w�H�
��T0��5d�R�з"O�ĺ�� �fI)���J��Pa"OTQ�+�>���R������y#B"O�zp�߁R!	��h�\u���'b�D�Ӽ�Ά�2�2��תJ	!�$S�=�2A:"
p��T��/K!�d_
l |#�J��`37!���7~`�����X��@@Հެb!�DT�zQ�;qʪ0��dip�7h!��/:!�Vc��[��uZ6�ĭb�!��̓e��س�@n�� �6E�{�!�$�C�2T�5,��S��BK�!�$K|��`�� �s��H��X�!�䝖{�v�yr���v����?i����۹$t�r�_>N�����0?s�B�q����"E����J�aʓ
�B�p�V����Y���	榃�[�$B��r��I�%$�r�&�ͺ;�`��$)�I.x�~l�w��q%8 �s�sV0C�I�d-<�jƈ<(̹��݃&NC�	/@B|X�h=���to[�:���=�
�'[�.���jS����K9Y�	�\���Q{tġW
�)u]�Eq7*��?<C�	(R�Z�����$�L%�#����B��+w��9��G9[]X��̓^W B�!U���)Q����t�}�B�"&��PZK�X���ɢ�C�	0��<�	 O���H~�=�
�'o�<��"��X�=�Q�� ���'�a~2%�%�Ri glҰ�J�v�	�'�H�8���.E���{��ƼBvIZ	�'Y�X�a@o��0���55` t��'�Y�'L wTҠ�WM�ۨ���'���vAF�zt$�E�m=����'q&Y�XF�aF���3���2�'V���)V�iM�$Q��:&����'���d�ä�4a1�=:��
�';��1G,�%:��:p����
�'��Q$V!ALL�I&��=z�
���hO?�����xFuE�+�}�5�[�<�''TL<��;֊��dVv��6�[U�<Q0%�$�HE�� H�,G���F�R���?içd��au/N2k�N���(�DMh��ȓF��41G��0' ���jՖD�ҵ��_������٬ V"A	�[�ra��9�J9��.��m�Τb`M(l��m�IΟ�?�����'b p`�I�U>B��	Y���J�"O�\���@�:|cp��8,k��9D"O��q�R<_i��z�f�"���(`��{�OvQ��BQ!]4a�bo΍m��T�
�'>�h�`o�.5�X�r�܋e��8���� �Ur���VrT�o*CȢ�Q"O��C�1������;�����]��?����;[��t�FfكT�qyԊ4�!��)M�H�b�,Z�����D�'�!�d .a�~� &,�Hy��a%T�L!�D� x3ઌ�x8Z��8!�Ǝ6�fP	`̍��R����7�!�D�hp��Cs�L�SC
3{!�䚎<h�Y4K
�*xz�ș�t�r�)���"��K�N�������p�����'A8p#��)���j�g�d��̻�'J`4�qOG��J�3���b��]��'o�|��F�1��
��ȦU�D1�
�'5�AAЏ��W�5����<��9��'O��:��-B���$�^��tb�'�j�Z�*�]â5��!~"!�K>��k ���`�(�f��	^�48��)"2���L;w�I���r���ȓB�,u;ă� ����o��?>4ч����Q�ʂ(���EEȚHjM��_C�[PL�BU�!�@犢l0���ȓ]q l�X7%��UТT�[��	�?���~z���z���dΗ$`sp�+cj�[��q��b�<]���(�:@�;Į-D���C�'TJ��2u�Gq�❲S -D�Ъ1F7*T���BbD�l$D�E�+D�X{��W$�nU�R�Bx�y�d(D�4�������[פ^�u�!�%D�XA�` �	���X!k;�y�p�6�d:�SܧQ�	�a��J������˛.}&�$������y�e���]�$H&p�B�I�nr�BG!ʮ #0��qb�80�DB�	 (�r� pE�	>P�����/6`B�	&~0n| �(�"�:�� lȪ �HB�I�k4�
�fQ�j�ap͓�u&2B��U5쐺�Ac_�ؐghM=#�O��=�}"Wm_
L�B�3���`�fM1P(�}�<�p(�#8��J��;n���H3��v�<Y�h
�W�K�e�g~>��d��[�<Q�� 	=�b��`��u2���	�a�<��WIj������-���^�<�#�"P��@@�*@ј�����T�<�A�C/�h���<�"����MG�<y�i� b����n��?�����L�<ɴ�ˉU2��I�dD�W�H:(�K�<�s�Q�vC*�7��JP�GI�M�<� ÔA����Ł	"����`�<�F�Q���@
c��;n\��1�i_E�<��JRp���q '��5N�A�Bv�<9Q���(�X��G)-�Є��Cu�<I��խ^�z�c����Q��LJ�<�J�!�MjWH_�q����\C�<��A�Ƅ����B�`l,�H5c�E�<�p�O�Qp����5.��l�Ue�B�<AG�v =PS+		0���{&N�t�<��Zz����*3�I����u�<Q� [��R1����"s�pˤ��s���<y'��e����ƚ�<<���o�<)W��[L}����-�X�	��B�<��	[ӄ��QT�.Y�eY��r�<�``[fXB���ҭJ4,q�r�<���;�4j�ۓNE��/�I�<	4��@;|��d��a�6M��NI�<���/5�UXU"�3Z�=C�MYy���<� ��zr�]��j4pFI͛BZ�=YT]�`G��'a��1� 	��ݯO,��E�Ƕ]����O`��Ĝ�7�nݩW�
J��-R��>�!���"q؆!*P/�6��rQ�
LC!��2�.�i�	Ⱦ[�&D�M;;�!���7���xŭ��N�R`2aEI1f�!�d���\�T*�d]���;;`�}��� ��I��ǣ܉�ifh)D��)|�Fp#ǡUZ�X�S�<��OZb�QLL����?N2�ȓ(L���g�^=\�hq��F�B�2u�ȓJ�P Qi��v�0���T�b=�ȓF2�z�X:NƲ����� ���f�8�
�N+&$`�`�-������1b�εwhn1	F#��RV�1��7�{��ݽIf�2�^.|hŅ�#�D���֊3i��J6��! ��ȓY=RsL͊�؍�"c��gVb��ȓ4��-����%�l�ȥ��.)�p`�ȓ2�"�+�oKO�0!�g�,�����P"L��`Ɏ-a*	ۀ$��Ԇȓ3�"�(�-�'��Q"�/s6�H�?���D3?c�-��L��(}���'�O[�<aQf��G�j|"�) ^
�Aa�� T���d��O�`�s#� �T���i��1D�X�׎0Ԙ��"�ظ�'1D�$�d-��,@���3��i��1D��s�?	ͮ��'����t:��2D�tp�ʃ-%�H��%�
!,0ĭss"1D���u*�I�D�+�O�8:V�5��.D��qBCK2n�"�B'H��U6��Pa D�+b��.7�L�'��W����+D�TA���5�&�)���zvNm۰�+D�XK�o��+���!숢�ja��*D�h�gc��Rڜ�h� 5lU`�;D��Q R�5�l`�ìRz�{4�5D�\9���7
���a�f,@\À�5D�Te���e��c�!	"a��1��k2D�d���%}n�g�=|bd���=D�4$��< (J���Mœh9ZT� -/D�\�(0�* ��H�/a���f,D�l�#��}Y����ֹ3�p)�?D��y�jY�4|� χ":O�P{֯=D��;@"��Q��E�)���@6D�te�_��u��#��&xrq#�7D��)�o�ʄ�[��ȗR��1Pk6D���щ��:9�%�3�\b�H�6D�쫦�Ul����3(C��Ŏ3D�Hq��:9j����3X�rD@	2D��Z�%�Ѩ�ʊ�
���5a3D�؁7�N}	�0��1H��b�2D�(��݃8�����uc��@�l>D�0k@�ږz@�8����2mୢ��<D��W��'���2��:9���S�/D�xb�������$�C��X"��:D���W�C�NF���P�N	=�����8D��Itn�)oE��cϏ�n��ȓ�f0D��pg�̘aͰ���C|!�ibG�,D���A7,��@#FB�3-�9Qs�+D� �F�Y��T�ӎ��)r��-D��"2ț!u�&U+�+S�gG��3�,D���Ȏ Bl���Ϭ��%�'�$D��p&�r` �%�
�w<H�rq�=D���`��xyz��C��  zɳǊ9D�� .,yT�NyP@(!�+�o���C\���	e�S�O�F����x�$1�%���w5������x(�X>D�3v�L�~�s�ݢ�y"P�3GP=�3��ft��d��yǟD� �'
'6�
P�L2�yR&��$>B���I^��֑��C�3����8�@@����L�Si�C�@���"O���@�ܜV�ԥ���9�2�"��:�S��iL�t�b\�`�sa�IK"�L�Q�!��#� Iel��|�5҄�A�'��'^?=�^�P�7Iʂ]l�J�A��FB�ɃJ4�p��|+R�����i��C� {��҆�>^�D2DL5~
���#?y�(8~�0���T����GE�<�2cU�";x�BǂO� �bl[�<����1 X�
�N�Y�8X#�\U�<Q��R�C�ҴJ�n� �(ix0�x�<�PŒ?B��%H�0Pw�T�Ă�r�<��V�b��H��H�K�m��I�<�Bұ*���VC�)I�m*�%�M�<i���T��:2��U���E�N`�<�l�#�~X�F��	
+���&�[�����*��1�D�� ���Aԣ�vNze��A�<qPř	<�2<������q��A�<Æ�\�R�ԭ�e�!��`Hz�<�bD�(o#�\:g�V� �-P�J�v�<Q��%b����O�
� Ay�Fr�<Q�o�4R[��3�׏);���'!7D���"�Û._&L)��.���A?���O��b>���	�<~��c��R&V?H��$�^�<)�ɒ�d���(�h�>�㑆	O�'a��@�sF�@��K�	���krbL4�yr�0��j�[� ����n���y�㐤%��q��y9��Є
[3��=1�yB�P<+R�rࣚ�u, ���/�y���/C:�N֮j��Dz�!H�y�A@�e�&ģ6�Я_�f�������5�O����Q�T�(�1�̐@LI��"O��Ɓ�4c�1�W�P*�]X"On�9��7d���ڕ.*J�3�"OaA��ˁzTa�pCY/.��K"O��K&@�+,CH��2#����Yf"O>a�a�L.�dX����>X��h��"OȽ۠˗��QZ�֪�,�q5"O��t��yz,$8�*��6�0THA"Oα��' 96�4P 
 UŎ!SE"Oz��d�E}�J�9q��v5c�"O �"��5 )��!g�#)�U1C"O0l(��*0/nX�\���2.�'8!�$Y�����'����D(Ң�"@#!���^����˓�
�F١5�Y��!�d\U�\m������KS�N-S�!��R_7>�ʖS����-ʢ(|!�$I�s���ˆ4�^|�4��0*l!�D�!	C��òK�jK ����6�!���)�b)"Sb0Nt�f���%�!򄖡N�PpI�̒c��8���y!��e�e9��8#����n^!��ӐZ��h9��Dwd��cV�!��cEI��Q+R�P`�ϓw�!�Q9{�8�⠅�7���(���X�!�V���a8��/D����E��!�d��T(^6e�-h�|UI3|B�I�$5*t�A Ĭl��0�:T+�C�)� jyr���N�DXس�Y�SQ��*�"O$�{�k�(;y���B�R`�$�f"O漓'�nVzU�E@F�U� ��"O�	17V$_
⡫B��&�X!"O,�������Ꙏ0���J "O�e��L��'7� @�I@?#D�R�"O�}"��ٻq���86��H�f��"Od�y�GF�^��2��:3����"O��G�B�*@���lX�Q�fu��"O�e�L��A�N�q"�Q�(`d�'"Oցc&G�"6�1T凣X����4"O���d"V9X:��A@Ww�9�"OJ�(",�lJ\Ȃb��(���"O����Y��|�f���M�\*�"Ot�:��܂!)�9t��f�B��&"O�ah��38����^t�<���"O�;�� x�nx���8D�j��E"O�����@�c���/� �Z�"O�}+ta_�r�ށ A��E����"O(I��M$&~�RŠ�� ���"Od�Q��(#h�ҍ]'N��q"O�����%݆����
��a�q"O��C§1�^ 8E$�rM �;"O�d�3iƒF�P])a"�]�1�#"O��wO�<r|qs��|��4��"O�M�����<~np��O�����"OD(�s+V?G̒�iDc��ʬ��"O<�AeO�lɩ�!�
?�ʕ�"O���ʅD�f����<�Sv"O�ՐW�H�<�؂� 6E��+�"O�]�c���T3��25�	0W"O��k�$
�#>���hH��Z�"OD-{#�݀\��kg�^A�P�ɂ"O�03��k����B(o/<�0u"O d�i�	s�qRhI�[���u"Or�S�H�*b_D��L~
��!�"O�yK����"5�QTb�r�Bd"O�X��ƫw��k��A�o�j��Q"O�D�P�J6S@mqEO�f�`�8"O�@3"Ҹr��8��
�,�0 "Ot5Ѧ�[�{�Lz1H�c��Ѓ"O�ժ�D�;;���g�V�"�e"O���d-��$ �1���E� "Oҩ�MS	a�&a�7!�~��e"Op�J�	�j�`��U�<m>�s�"O��#�T�n^u`w�	wXVh!�"O ����,7�������^��j1"O\(Ӆ�A�k�Hx	�'G+d�����"O$�J'B);W�����P�J�hDن"O�	x��=F���f�Z���]"O�jc"[�_Xؒ�\z���"O��)��F�6x��9W��9(��	�"O,�r"�wKb�R	���"�Ks"Or�aS��28�da[�m�*�Ӂ"Op���oY�"���$o�Q�"O(VK�S�&P8di
^V`1�"O���օ/O����7[��a�"O��bkZ#?�0��&��l��#�U>E��L\3[�x3f�o�*:��*D��
 ��J��9��A�ɆqI��	U�<�a*!!�f��5%щM� �h%M�<�v�K�8
����*���d�XR�<	�O�\ �l�T/�5�Zr�����%�,G{J?���_�9΢ܣ 
6}��
>D�� ��o/6�� 0���I�|�i�"O�R��#��!�B�[�(ܚ�"ON<�LӜ�Ł� R�m�Fu�P"OhM�Q�I��\*c	�:K4�Xkf"O������9�� �BMz�4@f"O��7��m��R�ťl�J�JA"O�0�@�Ҋ)�E�nY"�!a"Of�
��A<`���G��uv�%�S"O@ҦN5��l9�
-	����"OD�'�')�(g��9ό��3"O<����3%aҌq�@2�J�r"OҔE˺B�	kĥ�/b�L%I�"Od� �!��	`�x�qKL(cؒ��c"Oz����ۛ|	4���J��Yq��G"O�!���;NԜ�Sk��UFjd�"O&p �˛)eA�M�&����u"O(@�
��"�\��-�D�`\ v"O*E�d�R'A(pJ�͏�;��8j1"O�ؠ�Ŋffd�0�%&� R`"O�"���c@��;���b��u"OBi�p�
�2��!RC�5@�X��"O��Q���- �"!��*,�F"O�(�K�O e�v��*��q��"O���
��<0���jؔp��$��"O��c�	�!1�F�c�	E1T�̐B""O68ɤ��G�(z��[-u�a��"O�tӵcO�J����G�7t;V�`3"O��X�.�� :��WG_�dN蕡"O�8�vaD\����@�#>�]�q"O(Mj�@�r�t�	'g�
c0��&"O4�Ä��=Y���'� ���P�"O���VX4�0��T�9�ȸ"OzH��B6]�z��kԝ{�T�`�"O�̋#�#�ݢ�J��
��tCe"O\�`��R+?:� ��/uw�=�"O^��@�%rM�lbr���i��Q�"ORq�3�߃4��(1k�8^��"O��m-!��m��L���ND[�"Ou��HS}+F�c���c}����"O6)�Ł�6^ȠЋ$��w>��"OҜ�h�.|W\�(��
�ck�0�"Or�Q����;���Kb���"O���tE�,20k��J
(h%*�"O���&�EL�ٱ5A��&&��"O�<�*�5��m���ŹV!��PB"O: �4��ƴ��o��i�Q��"OZ�z��C��q!ĵ�4��"Or�{����Y�*4�a��8u����"O�۱�Q�L��|��/x�!��"O��G ��m�D�6oBx���"O@��A�b�X)��-�}8|8��"O2E�4�G  1{$��&z��e"O$ d��b`��쌨�J��"O��F��k/�8ZG�¡?�z8�b"O!�kznQ��{�Z1+�"O8-���U
&�.�+gh
NFc�"O$���� �KE\P�J1&tyC""O�p��"D.1>�Y��U#G~\��*O��"VM
�D��Q�D��Y�'`~�)b��<���M�~�܈�'�`�`�$����-�4Ԛ	�'���b�畬b�
Ż�g������'[�)�2�SR-��#�'Ɏ�H�Yf�N��+Q�O9�<Q��� ��������rqu��-�`�g"O���/ 	҈�%��� �^�i�"O�4*�D��.��P�]�CD���"OH]AƄ�W��yi�0Y%j�c!"O����a�A�aϴS�Y�"O8!�&<z�@A��+N�$#"O0���S>K6�� � 4���"O�8�@��h��Oжj�䤓"O��C�Q�*�\H�ŋ�s{ֹX�"O~)��#V�XPc��/1���Ð"OH	2��?~H����tcB"OnU�"ꕃ8~��b�ν,�,�I5"O�u�w�
f�:ɳ���-T>l�W"One8A�O�<�&.D�L���"O�S�M�x*����� G�HE�q"O���&
�/6|�b�I���hؓ"O|����Y:��Yڄe�,N�6"Ot��uC(���pK��d�P���"O ��e���9˾a(��O�B��D�$"Ov]RlU5L<��crjG�j��2�"O���pbZ�C�VE�4�Eg�rQ��"OJ	�(U�IV�!��FAf��@(�"O�ih�ᒰHI�E�2�O*<CL��"OD�!U�ƥ�������I��� �"O
=��)9�'������r�"O����MK�8H�*K���"O���A�u�l�b�У(�Ԁu"OX�H�T�b�JkS�K�F):���"OћBהX�LvÝ+"�2�)R"O>�J������X��?G���g"O���4&K�u�z)�bfѱV�hZ�"O~���K9T'#ۚV��m��"O ��B���I�R�0���C"Oy���ۘB�𸆁N,2լ��"O2�A�d�')����F�!< Y"O|��0�^�Ɓ��,*�A�"OZ|�(G�n�Qp�%�
d�sC"O���KZ/`�l�CN���2�Sa"O�D2��۝A"\�p�8?�H ;�"O@D�	����е%֩ό�"O�kB�kx��"2�8~�t��"O�%��/���U��B�rYB�"O�b��ȓn0 ��ul�4[N�sV"O�Y*�K��8��e;8��"O���fB@��� �+�� �"O:��b��'@�2䓟Cf��"OJ`���*:��r��'r���d"O�ɂCl��M�4���C�G�B�3"OL|�凑$�v5Y��$
e�W"OF����<��uY4gO�@�fԑ�"Oy��	Xe�(�����&`+dL@G"OL̀��  �0�ゞa9�-H�"On��-��)�"Ù0G��"O���5�E7�caC,/߆���"O��ТM��p9LU[R`�� �*��"O�e�0ǢOg�ٲ�D�ֽ�6"O<@�AA]%Bp(1���r�`�"O&����E�~�����mVY�zm��"O�<�7�����*���	w��2�"OBl{��ɔC����I�,yx���$"O<���#F9-gP�vx ٢P"ORQ���Ops�%#�'�<
��r�"O0�1!�H�J;d�[֠F�A45�E"Oj=H��H$9�,�`���P�#"O� 2���h�s�US�n�.Z���{�"O���'�"5Y:(��I��q1 "O ��O��)v���O��*Pk�"O��[�ꟆB4X�'V�L�N��"OlU	$��A{�P���ɡ���*$"O6p��B�,���tċ�PRQ"�"O�T���?>p���e*��G3�:A"O���u΀��EO��t�Vk�+]�!�S-���M~�\�륧�#�!��%:��V@��A���!�,z>Le�ĥ�6K� D��q���;P�
��A�Z2d���# �)�y�h�x}���g_'\f�A0�D*�yb���&��	t� ,Jl�@$�5�Py��&?^��b�I�#8Lݳ3 4T�(��7M���x��I7���K2T���D�
i�J4���2u;��u"Oڬ{׆L/aU��2cQ46��
e"O��
a�0P�"\��!E�4q R"O�y�ΒE�H`��	)1�)��"O�R��eY�@�0(�-u��D��"O�:�
������!�V!���H#"O���@#�_ox���Q�8]J�Id"O"�1u�S+�����B�Nr<��"OJ<@�\+
TZ���F�4s�5�1"O�����˛oN\�p��0lY@E*P"O�uBDf�k�����L�DhfTp�"O��c�E�V��'i���Vqh�"O����� 2U�%ʃ�G��|�"O�ͱDI:U���y����)�T}R%"O�Ƀ1�/K�=ʤ�N�*Y��"O�R@G�{�2��@�O�:o�0q�"O�,{Wm�)b"��B߂	��"O���3#IL�J�%��"]B�"Ol�!�/��1FH���dH��l�C"O�;�F��IZ,s���Ts(i+�"O�y�vJ2CSvI�U�G� �^ur�"On� �إz�hh���]�@�>���"O�4xu	G�?h�Q'�%\�h�zp"ON%�֪_�=&"���d��y��1
#"ON��#�:36,�b�@/d���R�"O
�r#� P!qz�� Q4�W"O���f�K-HQ�CϬ%�"OjԚ�P8`N��R/+�0�"Ou
v=����6g�Tl�"O�|���D7K|��e�,U�X�R"OPk�O5V��$�9`�|��'"O���S��}�x��)G��qG"O��q#���+6��'�� L�"Ol�C�L�%�E��O����X "O�	r�ȡ_�
٩�+C�B�H��"O6Xs�37 4A#
V/s��"O�D��]#{�i#�	QX_.Y˳"O����W�Y�V�1w|Jlx'"O5��@�bz���⯗$p`�)k�"O����!I<b4@�υ6+��Yqr"O�����0���@�$q�Б4"O�l	��ބ}�#���F�%�"O��Ţ�>>X�sTV=(��2�"OhjU��8�l��%Abh-;�"OzX0�N���Յ�:(��zU"O��)��&,�h��K2]�|HE"O�H����#ιK'�,�S"O�ijQ�C�)±o 1��鰂"O� <d��V�{$0qbsNB�$�{�"O\�XfkL66m�8�pn
	�� �"O8H
���)F�"{ H�? �<\S�"O�d�6�L�ZJ�{Ǜ�+O�k$"OB���ȓ3�.�в�M0�"O�(!�8'_�����++���E"O�)�CAX,UI�	)$�F<\phs"O�=�ׁ�x �$Xb#&u7~LR"O������N��	��oN�j����"OL	 �I�j�L����3~��<��"O Hӛp����c�V� A��"O��ZW�ɡ\�z ����\ͤE�t"O��t��J���&U"����"O~���+G�>`���e�[	�^��"O\�:��G8o.TӶ��']�p�R"OH�%m��M��0� +E}bM�"O:T8Pb�>O�4�ka�E�
E�"O�Ē!���s|Y�d8�$ȒV"O(�a��A*�!��.1�$i��"O���'�љ`� h�Ƃ���I�"On=�#R�E|VՈ�k�Ƙ"O�*�jX5w����,�.b��ma�"O��Gô�*m:Cl�/\��|��"O!zdO�o���x5FʜS{�P0�"O��Ӥ'�jM���#k���!"O��Q���]��(�5O��v"OڨK�C��"	��钅ѳ:[�x
d"OL���%< ��}b�!Z@�\��"Orx����b'Ƙ
�� X˞A��"O�����U�5K��8#"O0]27cA�?n�� �
���A�"OrYIϛ9A�T0сj��7�<iQf"Oj��3�B!�v9�'G����1"O�����K�u���� ����3�"O��х ��ys��H��Ɗyw��a"OܘS
1Tv4��4压Us���"O���t�4xt�A%��=Kb��2%"O����j�4��L񠤁�US2�"OFa�R;Z�� -��ʝ�3"O�a ���K��B2^�r��P"O.1#b��LPP��>Z�(�Z7"O�ت'�� f �ć��%I�"O����']���r��<��"O�`Q���9v�8�RE��B�rp��"O�(��Ho�t�K��MnJ�ظ!"OR��Uˋ]F^��aaьK+,m��"O�0��N�)q�&>s !�C"O,d��/��DT����pHřu"OvȺ'OOxr6%���Q�A"Oj�$�n�.	�Dԁ�P�"OR��э�,8@]��\#4^lyd"O +Y�p��#f��x�%� ��#�yb%��qO�'}0��₡���yR��=��$�!,�
��D�B���y�j�[�����m�	a�ԣB�A	�y2�33V$}�5.�j��)�Q�y�Z5 �P��ua8]�zE{��%�y�IP�?n)���R(u �
X��y��I z~vu�c3[ �Ujw���y2����S�g�-XM4-R���.�y���3"�:��%���GYP � ��/�y���6
[X@��iP%CX�P�̸�y�c �4��9��D�:u�(��� �y�O5~B��%��9QRH�&J����p>� �A�T�X.W�2p#$��@=�{%�'����`d���#���\����Um�	ABB�	��bG�|�Q�a�P	I�,B䉩c��4�e�\�Fdm�DC�>\C�	��8
���<�蠁���= ꓜhO�<y����.D�
 .[�by8�3bL|�<�2�I�:��va�@���W"@|�<a�HJ*���Zz�{6[l�<�`A�/p�2QТ�]�D�t�q�<�lZ�PILȲ0�L�d�DC�+7D��a Jߧ�,�y��p�����6D��ڲAm�T�����D�J��8ғ�p<AƌƚI6 4�������E��v�<IWIҭd�Jh�c��O��|j%oRY�<1쑖A��@�D��
���g%�`�<)�e])�0�^�U2.@�f��c�<��$�95�2���o � hÌ�_�IN���O���0�D+a3r��!	]�bYx���'� ͈sJ4��=�N�%[�1+�{�ku�l��DI�8��y3��85-ӱ�Cӡ�De����ֽ,{n�2&C��D=���;4�T��;��]�BJ�\�����6O:6�UB�+�b���F��q�d��~��!\�(��Иi�Ё�Te�-l���<�ߓe�й���#J�d4�GO+1����"��}(����L۸����P�����H�:�r3aü$Ș�:d�U/rM��'�&�*(_�u�tE�B�QPb! �'�TH��ɀ(S�=H�.YP�u�'b)
�N5u�y����#����'+�� VkX�^�,�pĴ8a���䩟xG��L��D0bQ�����6�W�@��y�ǳR.��!Y�`7L�؆��`fC�I�[��I��qnE��!�$i�����2?Y�']2�p��P�?f�e͞�2�q�yB�'�\i�ga+:J���o8}�:�
�'��J��
9�A��( ��)�'D�贆L��R�c�ϖ/.�P�{b�'�XC��Ϭ]�N%@q��,q�t�O�`KP�'&x�1̱!u�\�1b'o�`�y�De��I}�?0�d�9d]���� �yR��Nlpt�����ؑ��	d�DY�ȟ|q�R�L� �ku)�/�Ib�"O���`�O�tc��X�U�V }yAX�D��'�1O�3���1��� �G	L���14��V�'�a|��6;�	��c��O �$n�4��DQ�d6O�Hd��T�(��憜u�$�#��5�Sڜ'��)	t��j���	V�-Z�D�FK%D�\"�`����0�snK'F����'��Ο �IR�S´�S�[��!K���jY
���_c�<94EZ�+��Vm��-��}�@����xr�]�;�j�9��`���j0�X.�0=!�B+Q�]��K�B�^ǲ����yBϧ>5�-#��,U�Х����M��'J� �ec&񬼣'%D#A��
˓�(O�� -w�L�׏D/.1��"O`}A-و|.�ܣ�lX�9-��9��xr�)��^�:R��R�	�LUÇK��QL8��Z��D{��IП.����cNtORH���+����	|�OYVP��,��8��vD[O>qڴ�M
˓tȨ!�dG����(BM6]'h�'�H��	.���$�q���u��A���Ĳ���W��`�:m��łSj�)��C$D�DJ�ԉ��ՐDG��亥(0D�� l��Հ̢�Z���a�+{�y"O��UM	���4{�LFQ̅����b�O6D�h�ͭf���ƣ�<�N�|��Inv��1�,�:6�5����8J��C�	�90jR��z!a��k��@yW�!D��"�j�=V~R)��X7�45��
!��n��d �'O�����Z���C�� D��a�
�n����V�*S��0C=D�\;wMS������=��l¡N=D������7pIc .)�XY�-)�d;�O��YG�
.lg�Y"�,�U@E \�L%�l��Iu9��[�A 6z�>M�d�!���zظȪ��ޮr�T(QT�ۧ|n� �O�����1�~x�w*�;�&����IΦ�Oܒ�"�Q �J��h!F��`rx��"O΀[W"
����{��
�@L$�d:�S�	�/0�ū���]8�D:��"�!��sư ��(`Rb	�U��|��b��h�'�����9ܠ�l��S7P\�ȓG.T�a��<j�l��'k��E|B�ӳ8�,��W�V@b�8��5%�B�	$��u��KK�y+>�"%�M�+��ꓙhO�>Eq����❁c�O���L*6L%�O�˓R�%3�+ �\N��p@@�[.rx$����M�lx��~�=Z�!]=62�C��2���ʠ(��L)��au$C�	�\J&�1���:UcL�SC���:"=ى�T?����#6��s��[R��h�K?D�:�t눐����Z]���!D��{`��\n�U�c�Z��:�`+�����IhL����'�#���p"O�Y��F�{b�1�$��U�>=�"O��*.��M'��r���E�IpS�'��	-}���)q٫*�L�E�_8�2�?��nx�����'W��hN߻UI�u²� ���IȩG��@w��<΂�k��5 �!���ȓ�̓�B��,S�� ��9�ȓj�,�9d���h0`F��-=~!�ȓMc"�z#NR�5�6�i��m��+�Ⱬ5��d|l�Q�43�A�ȓb�I�â�F|���L�M��)fO1R�b���9�g��o	n�+��u��'�ӥӚ���,?wp̱d�UvB�ɔD&�|6kN�l3�L�-�
�d#�S�Oq�lsT!�V�b���#��D�X�3"O�a�&�K�J촴�����5�*M��"O����=���A����U�|��a"O�D�"�N�^3n@+� <B\](�"O�|�䃒�T2��WI��<��"O�x ���. ��DdML�?�(t[�"OhU�3h��nq��. �)�"O~<�ƆCxASk��[<�H	�"O��FO�~�����A7�,�"O@�F��"F��W�+v�)�"O��!s���x�*�\�"��"O�!zD%�3eBph�gFBG���8U"O��($&ݡr\,QoX�=>�0��"O*��(d�1cg�����F�y�Y^�ع��ː8��D[����y�	��| 1����`�r�/���y��rP.���#�`�iRi��yB)˳by`��K,h��PKe��yrl�uw$$���_�|�d�/�y��0j�J�fށgJ,�Ah@*�y
� �1�ET!6#4%��&	&�S�"O8��G�;;&�y �E�s`ڌb0"O"�R�H�s,�m�����5@�5"O2���2���V$v���z5*O����B,
0�����4_�ՠ�'-<�pD�lpM���U$V��
�'����Q�6\��y��@�9 ��	�']"=9c�:A(�4��,�~�Y�'����gS*iz�H�rE\�~��	�'5`a�/��T�� RBtB*p	�'���+E�S^�j}��cۉg���	�'��a�e�{@G��)eA���'-|����qp���)ΰ`z����'p�Q�DL�u�6Q���^�C,L�
�'j&i�c�Z͘T86�sBʜ�ȓCz0�2L̥�8��%Q�!�H$��@�����A���^���L0����ȓ	8�I�#)I!.��M�GK7A b�Γ:��(���{��Lk�)7�uD|����Y��U��nQ{Fė,�y���|�nر ��!J^��D�1�yBe�&GZ�z�Dz��ARtc!�ya����x[�
�q�53U��y�G?pkb���N�v�1����y2d��3�r���C~r���r���y2hT�J�(-����)hw�T8�(��yr���;�@�b�h�1���A�y2"�A>�d@�a��6Z0�q��:�y'�#�JHCs@��g�&�r�/�yrGE)L��l�q�]���i�!���y�iʪ8��\Q��*s�i�CI���y�!^�=���1^��U�LK<�y�i�#T �0;��H�\��������y�m�U���bg��Z�����Ƣ�y��GC�%��G3_�HxtO��yRJE���3��]��3#��y�O�sw(��fo� :�L�  �y� ��`���n�|�����L�2�y���]s~H���F��ɰs��y��c�d{��ֳG���'��y2+�M!H���f9�z�;�l��ȓi�`�'݃��Ge�$Y�Tԅ�E�6�K�ʌ<M�I�Ǡ��[gn���Co���tÇ�_���)e��xO���ȓ��·͉;c��r��b�0��ȓG1J��Ѝ9c���Ā5�<����<Ȃ	��V]���(f�25�ȓq˖!�.H���S#�اC憔��MN�;�"<BH�C�E(�ޔ��u�.u!�!��[l@k�Ð�ya|����btɧ�}rd{��V�Zjl��A�09P�M(�ͺ��s�|@��. �e8f��TE�����Z�Ή��_ ���K5����ֈ�-�P	��3�@�Q�Ǝt�U�d␀u����� ��4��(4v�"�zc�[�#.HQ���x0��I�8/¢������Ն��b�7�;sw�Y#FA}`��"E�h�1�W� P�����$�^���dq�I���3il�1��� WY�̆ȓe�8�#D�|��,w��d��k�<	$G	�M�Ƹ��,�}�݊�Od�<�B�X(R�!6#�MT4��a��m�<��A�u����E�L�zTb��o�<�"� i�����L�#%��7�O��y
� �4A��(g!H�m
"���"O�5��̑6,�����[/A�vd["O~U!f˲G�:�(R	?���"OF} R�D���{ eA�u����"O%9��'{� ���J��H��'"O���w�?��L!s�SOU<���"Oz�aDL�K�8yi��O�8G*��"O6r/K�z� ���/n80�"O�0��D D����'�>�L�J�"O6]Pd�]�p���d<wr5"Ozx��wl� @������"O|x��oǪmu�`�'oJ3Z�|�:w"Or� ���S�����˄&����6"O.�A���k��uإN̐I��H��'�N!�k�X�	 `
������_���
�J�$�hC�	,� �q�ǔ�dц�2R��4�VC�I(T�@A��
� R4�ۏ��C�m^a�d�ȋS� �	ybB�ɻ/K���AM���Bjס=�B�I�g)��S�>v� E��G��J�B�(2�$�"�%ՙG�(ce)Z9@��C�	/^�v�`G	\4[�L�X��O�tp�C��,
��)��CL����uƎN�C�I�t!G>2���!�nC�I�eIt��PC8	@$y��3�*C�I�|mT��&��5k]B�	/Q�?���мE��P�e�BE��O��#�.��-A�G�8,��4$��:� ��c��=�`�A��*N(B'�I%D�k�^i[��6�4��j� �=e��٨�E�l�B䉠-�R�X��+O,���\0b�4�b��	6	�ʴ1_���d3�g?�&A>P��y���L�U{rX�<���ڶb�Hi��
�G,
�fF�d��m��9d��l�h<��J�:��F�T29;v�8CK�)��{�×�6��Ȓi�L�Fy�R$m�B�Ӄ+Д�Ց�!U�,G!�dI�����F
�z� ��	��)
�O4�+�� �7.hY���3�zc>Q�Q���
���Kq����0�g;D�H�KY
�F���E�0��\h��=������E�tD�2�I�O��}��<��KX�;C��Z��̑5�T��'�4�1CO��ZV2�3� S7�����1�d0��e�D&}0��XM�Ё�D* �1!��oܸ�C�&|OhӦm��v,�!eĺX��ؘcAġO����}��K;Z��ʓ}�dkW�1�)���0ʇ�<�bʆc �"<yA���0/ pa}{�>)J�B�T߈�z3CM�)�³���*�'� �� <�3�5C��Th׋��dW؉Pv�4Z�U#d-�u�fTx&��Hy��)ڋR�z}�rj��Ff 
g�AbO��OW/������n Aa�D����Y���P���<69d�`aE~"�}ff��W���	����!��bWD�P�	];g����NcB0D�
�G>��T�
�T	�	�F�����Д9�|s$�ϛIea�t/��nW��H��C�y����f
у�y��@�px�D2U˂h	~ �e��i1��O�PЋ�<�1�1O�UR���������n�	6O�I
q)�U��L	צ�Km�I��FW.8��)1%		roa~Bֈ:�TLsE�� -��Cо�0<y�"[)O@� dX^~�mA�[H$h�i^, -��P��y��6*hW�[���}�"�0���6?>\�Ò�V�`ya�t$W�W�����K�GVv-�"�Z��y�%��7��47�1za�*Tu��$��{�BZ�V�q��'.��"F/�l���K/����'@^EA3b8����+pL;d�Մ��E��	�&��t���7fU*bˎ�m$�C�I�'��J���MJy�u�uC�C�I�!]�Y GC$5�x;�jA1y�C�i頁`����Q�!O*r鰱x�'-� ��F%�$�\r��C��@2q.��`G6D�� �I9�-��9�,:��Mr�Z�t�-sP�iS�
ν���z�i���3)�H�냮�;-Fx��"OBH�T���$j��1��2t �$ĤNǞe�"�ЈA(��O?��P rC�E�� ^�[n��%W�X�!�Jt��a���n����E�]2T��6MA�t3(P�m��4�B�S�
r>�Z� ���'��QQ��{�zx�eP�z��5h�(�J�ۤm�"@ؤ�1f@�z[�]�PgSvܙ�bńa,]��Yp�uE�=\O,YY�
٠[��C#ԃ7c�r��D�B��@�2��E�x1t��(m�<��)�Z�!�-���'Å�E����)+�O�%R�X��~B$q
 ���q����-<G���`�A2Z��Q��ۍ<�& ��d�y�I~қw��u`��Y)@z�{�J�`l���8@y�����6@HY���F!p}8xY��.��l$!ԗ=�xr'�B@�* ��)k�]0U��'��ݹ�yEѨ	��K2쏪*�s�HT��  ȼ%����O���#.��6<u1�*C54T���˖X�
�KQ�q#eL�0�b��+�=�|��$	+g�܁0 Ű_9�d7]��ß?�X�˃!'B�\�6�ʐS�*đcA`��� ���$���2dU2:Bّក%���`��Ӿ�r)!
�	�\�wbج&Ap�׽_ĘX��b��$�D�3GN��j>x����H�'XQ)���p�\�V�ZΈ@����D�g�}a�JJ(�"􋈈3�M�U�)���lTde2IE�rT�>�Iv�#f䠸FɲC��9�p�eT�8rFFo�S��	pZ֝�.����BQ���'> I���k���a�g�a&� 
�C��)�ZT�v�>QD��d��wF��h�F�����&*!!b5�Xp.�T�XD�zx���T��`�'��p2�m�(:� ��U��w
���4O��-I�'���Qq�.��va��H�Qw�=����'�`+Ժ#%d�K������:��h�CF؞��G�
�i�P�'�m�O49��u��
޼a��g����`3�X�[��Ѝ��h��d..'2��T\a˖�
���X�O�ir䣋?^^L�'��ӄ(G�|Ѫכ\Ȉ\cRK�/����!���z�ٵ�4%��L�bh8���3�q�����5�5� ƀoX�7
 @x�'޴<r���哇y4h��lH9Sx\(�(���pF	��!�.��#�T���I#r<��D�[>?�@�H�#�b<
��	�O�������U���(�hF�p9��([�>��O0��X$�@8_��jd�Y�S1z�B�"O$!��c�
Q���S�I�5QXt�5aR2:���EΌ=0�TqS%X���P[���3#ɕ7T��%A|�<9b��) ���bI8I�����	&����茤CzP�W5R���) g:����f�v]+���� �|�@�Ë��<iAo�J4
�k
�N|�
��[�P�u#��3�D�8���g�&�雵7 �	c������I.V؅�=K\��#D�� � _N�@�m��c��{ȍzA���7�^	[�P�FA��}��Ac��ʟ��:	�%��;��܄ȓ :��X#(Nuy
m!3o�(j/z}!�c[�7���7�Q�0�ҽ�6��?�>闀�R�
�)��
�"�$Oy��4��`��QK��X�Q�c�7��@rM[v�p�`��6?����	�b��#gC��I����l�.O�#<��e	���)&�8D� -;Н�D�Qz�e#U�\y�/̾�y�E�?	l~�yn^>I1"h�w�S�cZ���Wg����d�7%>���O�ѩ�C��+�d��UO���De�"OJ�F�ߒH l�2gS�+��P	Ҋ$�Dӊ)��D)���$ǥ|�T��O�	�4��ʍ�i����Ҿ��e��9�6�@�AM)�M� `ހ�x"��J`X|I��R�.�xMJd�X�y��	!N�� ����I�yB�l�U)� �Ex���&��9i�B�I%*�����|j�F(��r��B�ɂ6�V�J&�%�pu�g� 4l?�B��/S�������(�u��&U8C�I/z.��#��i�
5QD�ݒ=��C�ɝ{�,P�Ui�^[�@Ҋ%`��C���� ڃ��/tN�܉��Z�y*C�	& ���^-Z,�X���צ:(B�	gx����� B�,��!eR��D�'^�V��V�B-r�%	�!�dєvЖ�F`+W�x #cL#eC!򄕳\{V8� �Η����u	2GE!��Z�f���ʶU���B�NZ+tI!����- �a	M f�3�#�R'!�d�w�R������\�Hfa��X	!�� �H��+)x����@�U��ڡ"O��#A)�H�h�Rtᗵ�.��"O�a�0�)��ṷ��d�l��4"Oʉ�g�Տ.�Ir�AX(#GF`s"O�0��^�dK�QD`Mf;�8r"O�� u ͡�RT����:*��"O��� �\8\�H��R�<�� �"O�){� ��K����D@��lu!"ORT{O����Hz�ڗW|��x&"O���2 �0{L�z�J�f\���"O>@C�Ʉ4:h��&W�)T��$"O]�g���R�������.!�]����҄�	BbuSv��x!�ՄW����hAz1��ہ>]!�R)N�ZѪ�D
}����tB�l!�K�GM8[e��y3$4��!V� T!�$_�>��+� 6F'��		L�|D!�d�
R�pj� �b��&hB9 >!��R�ef\䁀�۴@���xv�S!��v��,C�+_;�)2�T�g!�[
N���"���,�
��d`��8�!��ѣm9�,ڱ��%�f4:QO!�A�z�t�z6ϋ{��u�c��4W!��ԭ.��M��	Ҽ Rd-���!�$ē)� l��Ǹ�,���"�!�$���U )�I��+!%ٻ�!�� ܨ�3 OҐ3�"80r�[x�!��ۺ_�J��j�v�e,[�p�!�d�&��l`�"N3D�Zz!��ic���
�"3��jت�!�D��X�^i{b��sL	� `�% /!�D�9Qw0%p6ϋ�W��q�оl!򄝵Y�֕X��+/x��+[6�!���X�$�@�F�=������ƯR�!��/8�)pR
GOJ������r�!�dּ�bT�0F��r"څA��<�!� �s�@��sGө@�Z��Ra���!�2���s�
�1�
�߈`�!�1x~�h�F��%{
�[!�3�!��C,�Ȉ�� ͫ7�$P7/V?P!�%k<�@�r�ؠC�<]��n�#�!�G.�!ⶋA�u�uȳ��r!�$�WN�4�B���|� q_0ry!�dL�qI\i�T��1���@��x!�5�N�*�hR��8	�B�m�!�DV�Nr�ȋ���nqh����>�!��s��Y���*bf�0����'��h���� [/ډ��I	�O����'
�0Cх�A���C�X���'	���0�FB�+3�hm�H��'�}�����z�ڙ�#��j�2�:�'�2z��U'e��  �,?'�(�'��\Jd-��s�H���đ2<�٘�'�
y[b��.g�``�M #(����'������Q�`b!+Y*֠��ȓm;*�v��K޸ �R �ȓZ���s0m	2�V�B�SJ��@��&^�4�7͞���q�یF�pP�ȓ%�X,���0Sh��Y�-��%m���ȓm7@I��!P�dx�v��9AZ��ȓz�`��(�}����5L��ȓU�R���9��	��OY�
PH@�ȓC򐘦��=D���0򥐳p��݇�	B[��;"�͠�'��m��,��S�? ��S�Ӗ���7"1{����E"O���J���<�q۳���
�' �ъ� J�"Y°�D]��!�'�h�{�DI54ςY�A�"q=� �'J����Κ�s��h�֭��` E��'mrD��I4D�����ƔO�4���'���U���@D�D#_B�j�X�'s�)2%f^�,P���0��"O��YĄ�>\�2�{�BS�r�D��"Oh!�Bt��+� �*yef ��"O�|�V��2��X�!?>AV��e"O�Rt�¿ �\�Y�a�����b�!�D��J?����a�k�L�ģN |�!��D�<m��@F	�6tsz��!�DG!�5HP�HCʂ�@	������ !�$>12f�
o�K��*A��6!!�� C>}15׹B�e3˕�+�!�D�UP挚�'ϋpx����9�!����L�Dl�5�$4n�XH oǁE�!�$ć&�,HS��((o8��qa��
�!�dP����r�'=H��!�f֓&m!�$\r�� �cR2�8L�$��[�!�ă=��|�0�ڽ������K9�!���vB.��* 5)�����@�,�!��ޘY��hɫ{�X���"�:�!���r9:D {d�L��AA�S�!򄂝�"�6Ꭹ��-��Y�D�!���3Jy{M
���B��~!��6~	Vu�����k��ID!�!~W!�C����!g�ؔ#O�c�|�"ӎ=��Q&�9Bž�@4��%z#謑BʀI<��1DOV���-D����&H
z�c
-�?`D�q�D��0&D=��W� ����S��VD:���)�dC�I	���e��( gl�ू4�>��0)�8^���: &V�\(j��3�g?	ƥ?/:;�$��9QSc@y�<!Z|�<�������B������Km$8Q�L�*,u��		�\x�eY$$v��s��#�����:��PN��DXJ!�U= �0�{MW��ZTȵ�'�ZC���T���;V�	�[8}���"v��C��6T*UO�e������3�S�?b\�Bc�ES�TO
�>-B�	��(�ˢ���IF�y��,F�?�4SA	�*Р���I�f�#�g?IG߄r�cB)6R��OF�<	� �Tl�A���-L��0��o�(k�F�i!��4���M��D���2�������
��m�QI�c�@��^�S�H ��4�ԝa���c�Mr��_m2�"@�D���;�U�P� �)��=#�XL� ��+�qq��:�4"<	sg�y@���AǼ!T��>�a` �
1I�Р�fY*�����'����#�3��� >*�����(�������a�����?��-�r+�hy��i�-�P�g��!��H�)}<i���ЀW�\��˶d�`Q�s��.3�&Eb��ϭ ��ɯ\b�Y��d_~b�N�[��,�$���I;M�$
�k��h�(�cA ����$��h�(<��@!$�H2(ͯVU�-{A2��O��R�eџu��pp�'opv�IV��Nh���5��)�"O�t�� cԹ�f��V�Fq`�鈶H�p�襂0�2�3�d��=1���GCPY׈A�����M�p��)��d( �B��.���6�Dd&E[�Es| �aӚs ���DЛaN5��	�Om�)��ˆCm�	 #�HT�JN�3Xx���J�qxC䉳0�Zy���1RP*��1�H,�$�'��@�S��#]�M�㓱<���!,J�P�r �A '1�!�d�i6@Q�U��i��<y@C�.��N>q#�V�A����'�+��I���!��x;̑
�'$@��KV4k������@�
��HD?�`A��I�M�����dHlh�͛(tj�C�)� �e۰�Ȇ��a�� r�2�;�"O�C�%B����
4hY�"Oj��p�	���M
��%�X�s�"O`����	q�d��	&|�M@"O�i�./	v#���P��IP"O�4k��+p-�<���I|���0�"Ov4�AϘg\ɡB�3� 8@�"O��I�1�|I��n3��:6"O y��� j4`��:]#��#�'k.)�f C�S�Ojڨ�G�P|��$��W;sni�C"O����7�|��0�	Ed}�WQ��!�Hl,��I�E���ӕ�аDEɱr(�BX^���J!~u}Aqʑ.f��|bF�R;�)�T!�/�]��
�x�{�Ȣ��Xa�g�xIx��|�y�?ʓO����E�d�|#|
 25J�BH?{+/ɺ ��O�-yGd[��#~�#!B&S�U��8t��:u�9(xb�N�U� ��O?��\9R@2x(�eP�~ٞ��ٶ�u� Y�'.#}�'���Y�ʜ(�@��ǎF��{�'�N%���ɬ3?|<��	y(���6�H��p�{�aO�E���k9�l��Wz�'m:�Yp�)-�^ag�Ӷ>���H��:8��JK؞�0��!�Du���'��: *�&
 X�2wD�� ����Щm�j��'��^���J,I\j�ҷ�0x=�*��D�D�� �2�h��ct�����2��o�#�+�0GR�]�0H�0,��S��?y�%�,X+H]h�X7o���3j�-W���b����I��H����0�|D���/x��@����s���\�tՋ����p=���.9�MiC�P<}e��#��ަ	�%ƾ,gX����:c�呖�iL�k��K�m�B!�PA���AJ(��bʈ?~��$�(jd�܉E�G*z%�ݩ0i��G�!��<HwD%��b4d��Y����X�O6��GK�
{���'r`��o��|J୘u4a�s�?bP�ѱUV�<�gŶ+Fnq��lv4����}�Td�B�6}"aJ� ����f�9�d 9�c[�A�@��C��\��U0�"O��3�NX�x�ԝ����@(�:=�����Ј�D�Y��'��>��(}���K�k�	n�X�Ő7��B�	�i�� Z*BKU��;���T��mZBMPm���K�V��
���O����T�u����3�mA�� 2�'q�=���'����Ր8rvy	4㚪tfS�"��P�s'�W؟,�t�ɝ^o�Mq�͓<S�d��P�3�	Z�M"`���rqf^r�0�#M|b�T?]�xi�����S�1P@�`�<Ie��*'B`�o�&=D�XؗǑ#VܝraŗR�\���H{1F��'RB�K���9s�ت��_;q�@�:�'�8}�A������eXY����r��'@�� *��oZ���)���F}�!��㘕����Ze�!����;��=�u��;������f�)��gĤ["bar��E�=��f�nzB���Fc��$���CB)��j��T���ҪA(��iyD���10�,BJ|�A�>>Z�$㋉QL.�� ��|�<����;[\�H1�чz*�ԃ�NYi`�Q�����a��B<9����'�V�h���8 ��(qա͌LCt��'g�dڥ�S`8Зi��.�x	je�|�)�
,�rz���y���a�JG�z������Px��O
 j���G��\p�� >hm���f�~<�s� �<r�PBn�+�#��L�<� X�(Ұԙ0����a��-FD�<�!eŵotAweK�M5t��'dj�<�§��|���"X}o���lNh�<a�J=@\�2��$��d�}�<�f���'9����r�ã��C�<YV�:���凇�n�6�Nt�<!��F�\�:�E�U�4�V�ꡄ�n�<遣�$N�L����7��YS���i�<��C�]���.ʈ7�cFf�i�<�ƌY,A}|`�Q���`��ǧTg�<�@ÜLr����ݢ[Ɔ�)!��a�<���f#8��Bg�|���9F'�b�<� B,�MCaX���Bf�	nX�Ʉ"O|I7�5���Q��@g��('"OD8����{�Ĕ�����t""O�5�֪�/R.z�:�G��Q�,Ũ�"Oj��0)�4Rr���æ]�:Ot"O�!��.�䈁�΅0^O轙�'ʾA2�!�1590�FfÎ9y�'0��"�ET�8`�Ø38�<�
�'s��AMKt����$F��l���
�'P���a��c�z�H�e�jT�	�'�>�Q"�<`��t�'��P� ta�'�(ac䇇�(y�CC�V��	�'z\� c��;�6���J�j���'rp$)$ˁ8�T�B�ϕ7pt�Y�'�,˧n�'��]�"�-px�'3.E��ϝ�F�Hmۑ�s">��'avM`	Ė����@�hc(z�'��c�ņXiTeeIF�e�P�'�<e#�eQ�?	й���+*,�$�
�'ɒyj�gךF��j� ~� ��'��� C�:T�X��(Пe��S�'P
diJ���Ek�|��b�'�
����w�ʱ����!x�'�4���]q�c���}\��'Vp�!�b�b,y�scOU�R�'Mb1LR�7��ЂS<v�[�'�:�C ��
"&�;��I3rB|j��$Z-|U�d
�T���a�I�ء�$@���,��e?K���(�e�#�y��>"��a�&�W�D� �2S"�:�y�xV�\�͞=^Ƭ�bŚ
�ybM�/}֠�x@J�=i�Eh����y�$��\dH���4%W��9� F&�y��I������R2o�<�04iA���'�>�8$I�0|��iI3jx(�u�H�y���Qp%�T?�#`A/[G��KfG/}J~Z`%�N��0sU�=O�8�$�1_x �I@�]�W�L��d
cN������p�Oq���R1H����u��z�&��1�V'b4���\�xՠ�K�b�)���~Rڗ��#C�>RX�c�"�#^D�ya1M��2%�+�O1�����`0q�Q�g%�����;u��\HvJ��qF��<�c�U>�k⮘+8Tc�AÁ@�~<���	<&��O :���uL�SU�O 	�e ��U�u��L�6��A!� Y��[6(�$NC��0|j4��_�R�!� �m��;DTF����
;E ��-�s���bXw��������j��٠��+��� T�1��֚:�f�*�")W�>���T>Qc� ]�6��p���/b�0�I$AK��M��&�>)�D��aJ>!������ ��"�&�V11l����M
�jr.8�f�'wJv\Z�c�@'j�(��A2wn��'�2A+q�S�O�r0#�fÏc+�	��1�~� ۴f%�h�aL%�)�'TU�ER�q�슑��gl�K����'�����Y���`s�'Ǐ[}�`j����S��a` �J�p���L&V�3�t�O':�n�8�R�{�Nړeؠ�c�C��D�kI�D;��Om\�pD�ܬT><i��U��P���U���I�/��٩���|ba�D4m����(u�)�5%�*�yR���6Ĕ=z���
��܉Um�?�y��Н<�Ȩ��.ݏu"Z���'�yR����x����p��SF��yH^�RJ8qa#�_"A�B���y��63�x��?Yc������y��W�)�P�;����I[ �)�D��y�'A
$���h	Q�x��W,3�y�ȅ�o����
�<YDt�@�l�2�y2��6�F���*�2A��������y�,K|�Ѳ#�=�$�����y��*D��k��J�?�U:�C��y���1�u��Z�M��D���7�y�)
"ޥ(���K��4P����y
� �|�'�\tp|���G�*ض�ѐ"O�4��V9�󑤋D�ș�"O�,�/^1^��VΈ�\\��@"OZ�Jr���7���gJ�ba�C�"O
{r��
Dь�:�"�#�d�K"O��ଌ%<�����\=5�*���"O,5:�l�j�T�3`�<�=�1"O�x�2,�.��ԘA�/�R�Т"O*�*���	�R}2G�� '���"OP��<H�`��cB�y$)��"O��;p�_� ms�c��7c���r"O���դ��^|��	`�Ҟ!Fd	i�"O�C��S�^"j�"�G��5�^@:�"O����{Lk��?}nr�j "O�:�0�4AK<]Rn�ѓe���!�N&&1|���CU�:CnX��C~!�dS,�����,X!(�����=!�!�$4#ղ�&O�6|�a��v�!�Y^\Ũ�l�%x�:��⫗_�!���	펥��o���ޤ�&��HO!�ʧx�x��ck'%��0��V$�!�SH1����)	>IH�J�`;!�H	^�0ҡ �(�	�g��!!��Ղa_��֤�'嬭 ��ع"3!�$�o���F�X�v��N�!�$Ñl�<�r�P��`�C,���!���&�N� I��Vx�A�mT�\H!�CB�s���e�
�b���9
�'�2�0��!>��eh��EW�v�Y	�'M��AIԏ麸�F)�}��d��'�:��O�}P� :�O�0��'1�M������D2�p�&��'��)%��3�*q���ѥ^jz��'��9;5L��G�<��*Ud��'q8��c�SPw~��-Q!xG��!
�'	�����b͛6�Ƅpn���'j�Ւa�D�V�@�U:׬q�	�'����e�} %�:1�0@��'��pB��*:RT�t�T�/>�l9�'�dY��ީ����c��X&=a�'@���n@ Y�)ӍSE>����'y���$Raf�(p+X;���Z�'b��W+I6+I�M[r�5�q��'�0���C�	����a����'2ؼX��Ol�-��5�$��'�\A��G�7x$J�`K&Lm�m��'c6�0�@M�8�}���1��B�'��9C�B�mf�hx�����)��'���p	��JPp�KY5ɬ�"�'�Y���O�bE��!��{K�z�'=>�#���t�Ʌ)P�v��,��'Oa��Nʟ&= U��b�w�����'yι�DH�"�ba[T��-�x��'F��g��=b�#Tc���A �'� ���lƓF�$�NM�M	���'�2t��;R�D�0�<r"x���'���5K_�)+Rp×F(d����'��!���l�i+7�� �e��'�,��V�� �iy�kKU��@�'�����&���M�-�x�+�'���+��܀}�����J��D��'�*E[���ib�r�L��N�֔��'���II#�ĵ�r��M�Q�'��;�ą�.����4r�0���� �aSa�ߨ(V4C��_�r\x�K�"O��3t�B�
���2AD+YZ�1(B"O
M8�EF�V��ДO+@P�	Ʌ"O�`�E�jN�a`�1:�.D"O�u@�n�?F"�]�q�E/�Hi@"O�y�jQ�*�	N�%]Qb%�r"O���18?���Aܿ/����"Ox!r�a�D<��3*�+����"Od�S��{S�^(u���[�o\�T6!�D�G�+",O�4��A�"%!��'E����ۡQ"r	)�X��ۢ5����̞w��Z��y���N��-��T�~�@�c��y�#,O�.�y �V�w.���7��)�yB���u^ ��)Y'j.���v���y��93�$��Ř�X��Dh��?�y��/e%��YN�X�E�S��y!K�Hu	�₨T�^�Pb&���yb�Q0`��s쒷Qx���cʤ�yBBI/Wx�%rW�I� ȉa#̐�y2��6:��ԳF�;=�hi�3n[��y�ᇻ H��ٲH�4H�4<���] �yҥX�%�-ࡊ����L�2��y�ԝ=Y|U�oӶzH��h��1�yb�π��P2�#�i,$h��M��yr.� :���6�F�]��h����y�+�(�,���	Ô�����"�y�Ɵ�[S��Y���}��Iq.Ұ�y�	�'s��]���҄ML,����Ϻ�y���T�tD�R�ļ0J����yb�ּnJ�X��ۿ!\p b���yHB$�
@i�J"
�RdJ�nK��yrD��\]��x���t�8T���1�yRcĬ8��K )�6f�QH%m�%�y�OJ� ���5d����$��y��._�`[���;.���THE��yA�?	.���C4)(�Y�X��y�k��C�X�v���(�BIq���y�ƿT� M��&�W�b�� aN��yB��"p��+�*�DB����a�yR�ߌ5��C��T^~��h׵�y�O}�esAlZ�C��	�	]��yB�� �x�0�EC�A�4 ���;�yR 	&>�DyT%�2T�q�-A��yr�-\�9[b�܆&�8��6KN��y�S��F�'��,$�X�+W
Ӎ�yb���Wv���QL�2�b����yR�	s�r�SDB�;�|���=�y��IJ�\�ƕU�Պ�,�8�y�I�#>�*��ٝ�\�K�B���y®܂4�2Ѹ��1s�
)f����y���	9P����*o�Y�IB��y��Μ���0Ca���y�b^�<������4Zt �ۡfG�yb���!�[т1$��HDȒ��y��Y�>���K��Q 07h{��Z�y��t�8���D΀VX�4������y�EG�d͘��S�L��)A�
:�y�ǔ ;�T���>_�@|����>�y�%Z��de�C+�! �B� !��y�\��Q��'Ȑa��E����!�yҌQ�HNqr�d7RBhT���?�y�
�jW�X7�՝?�1weȑ�yR
�Q��1�B�ĵ/�ɨ�hW��y
� ^���� i�q�.:��A��"OD�z��*88�2W)��q����"OL*��צ,IN]�B�� <��	"O�[�G���������=3h�"O������?��) f�$��q�"O��j���/P��C��pU��Ȑ"OB�1��P�ME(H�0%6K����"O0�q���ZclLJ��K?|p:X�2"Ol=S'+�m�����G^�1��"Oղ�I����(��u?��!R"O���&9l
�|�Tɉ?JװQpa"O�����Z�]��a��(U?2uɣ"O�p��DҺ}p������E����%"O�䲐��A�R(�F�&~�+�"Oz@3�� ZO��xPِ>`�<�"O�h��	�CZ�=D�eR"Of�Y��["��\�외>6"�"E"O*Ԣvi�;ue����4 "<��"O8 )q$֧z�4��u���� ��"O�q�N��m�vx�qBQ0�4`e"OjMk��N�Z�낡W6E�4D{�"O�p'�7y�D�B��Ցk(�$��"O�d����
> �o�op0�	�"Oz�-U�:
:UB��	S�R�"O�@y� �6n+�L��NǓg:���p"O��0�֔\���d�-àl�C"O��+"��)�b�c�@�L��l2u"O��9T�X�D�4T�/_*�6��4"ON0�%Q�6�L����Ix2X�"B"O���1�E��*���#����5��"O��;�CθW�P�bAC
<1�,�Q�"O��`���0z
�!�
3v����"O\��Ͽx�zd�7 �1kqFZ�'J��Vm��$ �KG��6�f�;
�'��ĉC'�v�ۡ$_"2�>|�
�'�6PO��U�q��/�:�c�'��z
MD�p��g
��
�'��1�`�ܚG#�	�Ĕ)|�<hh
�'4�v�ByXU0�S�p׌��'�0!��!�%.T8A��%�=3����
�']�t��b��Z'�@�/�='T!�
�'���yu��,��0�'�9��;
�'�$�{&�ƪY���� #��+
�'x��媃4nک� d�""����	�'`DUB5
�"M[(�H�������'�<����7j,�$�]2�4���'�@t�bK�S$ڵ�t�^%]ޜ�
�'���AG.ӆ%f�H�����E��'| � ç�(,���I}"d]��'ت�`"���"`	
,��\ W��y"�t[�љR�:��P�� �yb��W�N��H{�ѡ�H��y��+0�|�爊7GC��k��
��yBO!P�+v�L�'���J�D��yr��120��e(� �x�#�$��yR�ݗ@ 0  �(�2w�N����90��+�8;vY���B��"E��c@��ħx@)�V@,@'�Q�_�ES���l��RԂNv��ӧ����`���2r��K$�����F(^
"�$#�Mѻ I�	;�k�j��OC�!{��LR}r`H�Z�Z�i1��\�E*�+���DƱ4/���4�װ��O� 2)�u�Y�k�H�L ���>9 G!�#���4�DS�"��� ���'pr0.B94�\�ȁ��y�gn�%@��)R��o|���!�v��A*�M�7�H�q`�jxf�zƄ �G�r��E�T������	�7���8���C�JJT��i	"2�<����T�LY��''�ܴ�`��Ua&y�p��(D:Bȍ�(�OJ�*�/̓S�LTjB 1�4=�	�'p��p�D؛z*g��$7	.q����4I����gR"t�Ls����'q�l"3��>	A*GѼL����^�:�x��R��$�O��
�L��׈�|�ܱ�u�X&��� Dy�<�G�]Z�yjA, 	������R�{ �d�Q	�m��ɚ�H#O8�#����HU�|���%E���1iD�l�>I���G${0(L���ԼtLP�f�3�O�PF��7qW�,;��� �␘r�>QV"ӕ@>��	Q��)��|��J�d%4c>�W#˓b�pmX��3G�l���9D� ���\�-8F%0N�,R~�b4J�h��=��T��	h��~2$V�nø	�̡f����Ɉ��y��O,[:��LI_:��uـ�?��#ќ(ǌ���c,lO2����Q�y�\h����W��@�%�'Є(U�
�\�8�n�<��I�ƙr.�W�P�{�TB�ɤo���h(0��@g���0⟘�CBǀO��-���ӾCr*)�w�[1+���p1�"O��Bc���9��qC�1I�*L�F-0\����]��"�g?���".2P3�c�/*s��r�Vo�<�Q�K�\�M;P��%^*r�F�`�	�Y�Q B�$_+a{�?w�j�
"d�z �0P���0>	��r8n  ��\��YA��8d��3͝-rc(��ȓI��u*��ީ_����J�}�B�Ey"iԟH��qF��GQJ�@)G������!��y��5
q�4�e��H�ƛ��yb+ߣs���:$�PX�r�a��y2��R�r��GC���¢���'AZlq�N}����+�f��<B�K��B��Ih6�9�����.*#*R�)�	2żI���[7�h��r�`��� ��T��H�*a�LM�I�6���	1S�.ђ�-V14��O): �F+�*R�J]8�E �W 9��')�઀�8/���5i��K ~�/O��ҶbU�d�"��M��|�A%8AnTt�	٩��`��u��\�ae�8H�"�����%0��35���&���>�7��7ET !�1�\Lx�JΎ���+��b��F~�_�Rw|T�土��Ė=E�ތ: ��YR-Y��Idid*�)Qa"���Qs�(z�.�V�I�X�j���5���� f�:ʓPv� ��1 S���pYC�4ttf\zOU�$Z(��"O�(�-?h��ٗ	7D���0�Q�`�V�^=%���GC�F�iȿ@�	"�Ϧ>1��έ3��<xv�5,�@ +GM~��i㏉�=��4��iJ�+0���Ԯ�s�����Ȓ*����v�����_uF�"?q���%-UH�B0d�p@H��g��X�'�"D��eU)Dܕ)'���<Ha�Z�H����_g��CS�S�*�����@���C�
P\B�[c66�*)�.���:����9��ן�p%�K/"±1p�i�5��ĳ�g?l^jH�E���:�.,;�O�̓��ԃ�_ {�h  cZ�'��Qh�"�O����0��bO��"�t�<�l;�#ۊ"��`���IZ!wL�YH��b)��D�g	k��-�6a�ڟ6���S^�,��坾{d᱃��*� ���xQ��S���9�����C�fQ6���d��nH�`r�ǃr���pu ��	D�����T�^�)�����d��n#V�%E�t����#@~��;C��Jm�X�t�&�~%*��'}�h)�I�88��f
�E������QDP62X�E���!<Y�$�d�rNe[c�^�$ϔ�;&��0rV�Z~����ՆH�0؅�	�$�� �wKp\��2�τ;d/�"�B�y�H��刯D�R�;��d �IٷԚr^�SF����'u,�aS*}���F�$:D��J�'n@92#/ν����'�ޤ��"�/�j-Z@��'����G�*��bP�V"����ѻiq������{��(��ŊH�z�Ӈ�L�w���/.1��(0����M��9|���JW�]~�9cc� #)Y�}8���;��t��K13~ �
� ��M4M��x�0�!x�i�f����"|�Y�枀q�(�֪��s��9�G
i��%S���*!e���^��pL�S�B�I%R��\@�¤i�~���KT�'nX��I��6�(L��O�}�NR��ey"��fd��su/��X�����\���U�PbP�y���1q}�x
�͓:8-rał���'(pxJĂ
*�ax��5f��8�ӁN�ﲵ����>�y�!��[����@{��Ԋ��yr��X�|��w�.MgN9`�O��y��8 �Tʔ�E� ]($��y"l�=]U0����9=�bipW���y�F-0��|1�h��7�R5��P��yRi�M�����"�����Ί�?y�dЌl����|;��7�ϸfnޑ2�C�%�a{ͺpF�h���O��e
8%90���N6p[���p"O�\��_871��!PNІ@�1���DÌ"�]��E����jM�)B�K� ɐB�J5)���"O8�j'b�6X���yV @���cсҭs(p��>q�b#�gy��ް4@�� �G�dkr�Iqꝣ�y2�D�Mzt5B�@�%�� ��kK�{J0��V r�hA
�iktȪ�x/��P�#Ϲx����Io4�а�n߼t��$�(�>��U�_�"!^�Q�K_1�!򄓲=$ұ�2�\�o�Rm�����qO��x�LT�r���1��i�"(����5tPYw��'s�!�dX�%!ԩ��k�$h�`�DL׭[��-
�B�(��Z�D�|�'Y$A���ҏ޾p����#f��m)�'�ʤA��'Z��0+$'�SL�|1ň�
�a��i�3�0>y��܀�PKV�s)nx���A؞�z3���Mpx�tG|�ѥX�/�h���!7mr��ȓqP�]���b�1 Da�,M�?��âh�"B6��	N4p!�@�LOD]0%�Fz�<q�&�LV�ԑ�P�1G�\���u�<a2�D;^k���)ݺ>l�)�g�Wv�<�U���B����DZ�l���(�s�<�ǩkIz �q�Z!�ӕ�Na�<!�Ő�~�hb3d��"���2@	j�<QP!��`�49j���9B�lDZ���L�<� h �"@�!�����٫Z�hʅ"O4i �I@�]���8����"O:���	 ?~1���2D��w?ʉ`W"O$� W�7�<���7^�Je�u"O4���jЀ[Jlp�sɳ+b #�"Ob�r��	�=���K�/����t"O�%��RHu0�@�%%Ȁ�J"O���($'�1Y����^���"O��(x�p����E;!h�\��OSb�<�F�
�7�@�1n����G�<ٖ�$
���ퟙl׆(6��f�<q��T=/�bL�b�	�F�ܻ�CS^�<)G�R2�!D�)
%£a�`�<��R<#C���Ac^�v��1j�X�<�PO�!e�*S���d���b�R�<�4��-��UPtd�R`�i���N�<��kL/:L\�`�?�0��RXF�<��ǋ�{�"��%K�!w�T�1��v�<����"�^����B"�m�u�ȓ��:�� ��i��"�$ǖ��E�dt��E1�n��S+P>f%��R��-��Ȍ)A��hjP%�sFf`��$��@�đ�\��	r"�ڦFa�0��t�ܼ�S%�8�c�!���ȓ�v|B�. <�r��23�z�E|��5����Z���Xd2���H��M���>D����.�9T�B��.3��!��Njϸ��CĔ{-�B�?ئU��ӷZ��u1�m�#�DC�3kT���I�PL�qC����b%(C�	3T$�%���)���N���B�	�W>�<!Hm;�%ʝA��B��^�h� E�R�J���F�_�B�	��Jx�B���PH�N�B�əx���sM]������,+�R˓m1B�<E��-��(1̕��\�"�"Y�ڱ�?��<�S�OQ���m\�z H���M.�bܨ`��O����8,�B"|�A����s�NTNU�|�qe���%�x�aE_s>��0`ݑ��y�'��><BS�2����<8JC�2��La��?�) �øo�$ ""O8�æ;�Q7��L�:�:�"O8v�׏xꄋG��rN� A"O"��l\�zu �H׀�1�fB�IP8�L���<�Rn� x��)��#D�TGQ�X��)��+ܳ	�����N=D���-�[��@cj�3i�J����/D��KdD�0o�1�W����(�҄�.D��Hhҁ^�8�G��6<s�Ɔ9D�̙���ɪD���5It.LBBi7D�l��-] 5`to�(*�A��0D�<떫�7������}��Iza.D��SC�:�ԥ�0@F�Z+�)���(D�,��"�S~�]���+n0X�%D���wm�'`kp%8�KC��4���!D����.��b�����B�	�����*D�@:E��^캀�u%�=iL���E'D��́k�4y�\���+d�#D��;�C"H��	1�� ��q�M=D����k�Z�~Ţ"c�3D��	I��>D��A��C �U��#�7{��
@7D����mʕ)�N�b�MC8��I#�`:D��0aG� {I��+q�_1E�E�6D�������g�"I"�J�+:e3�o3D���D�Q4� ���ئ�*A�`2D��U�^�"�\���<h�)('c*D�� �H8Ə��Ib���Wg0`��%�"O�\9D�9B��8�f̅U��T*"O��c�ė�>��6�w���Ҳ"O�����7��9K�㏇c�H�S"O"ux Ă!o|h`��"ĵ$��1#"O�E�r�� g
$#T�%�DI!�"O,���0�@�
 ��M;�"O��X'ʈ)VѦ�yb�Bى�"O����KN�fj,\�qd	��:�Z"O�1��@�=+j��@d]�8k2"O�DÁn� g<��9�CU0MB
!Iw"O���b\�*l> x��L+g9rᰰ"O@�;�-��/`6,�QkC�9�@��"O�m��kZ
G�00�0��-J00�"O��Zv�͉1������]f"O"A`���4Ǹ�Ү�9�l��u"Oԇ1</��O.X��"O��2ȕh�`K��X�ڰ��"O~ �@I�Y�4	RQǹ*0FthQ"O<�������Q� 1����"O�u�We��*���H�G�5^����"O>-Z�k�<�� ��W�R�4�w"O���5��P�Hj0��'x�`�f"OLh��T Ev0�#G:1W��y�"ODћ®�C�xMx�r̹�"O�}�,�,����\X�Q1"O�-��̭i5�-*[e�B��%�P_�<���$2jb�W	
��āR�.D�8C6���Q�4�A1��1XE�(ȃ�9D�8��M[�T�$�VC�Z[��p�b8D��w(�`8�e�S�8>�AH��4D��R��Ș�ȁ�`*"
�U��G-D����nB�S|<�0�
U�3��r +*D�pP1�	`��5)6����m)P�-D���⋗G0ĺ��`�F!D����"�� �2Q!�M�|�l�C�#D�{�5�H��&��QZ&K/D�t���׍_�2�Ac���V|���+D�p�VMֹ:y�A��	PC�%q5'6D�,K �T�Z�Tq����0	�f�5D��+#G�'��)SJ�.&���4D�D(��D�>��|arI 9I1�H.D���֩w��+V�ܰ�$d`�'2D�4Y��G�[�ڼ�P��c��
&#0D�����7�&%! �m��iۖb,D�D+ ��b���@*րBB�;�i,D�!� �=~�������g�(D��P �� $�A�K��,־��B�;D�Гd䙦St�(��&L��&D� "�ʓ�!@�����%o�"�B�"D�H��� M��q��^/TG�S��?D�t�ǭ�@Ȳ����+:��}%>D��s0!�I->d�ق)���I��&D��y׍����S�� =*�� w�$D�� G�#��1�ф���K>D���u!�B���iROLp%��M<D�x�!�ϩR�橒�)�dx|��n>D��.��yRZ�@��$K� Y�f'D���T̛�Ū����>�:�0D����A���l# I��T�C�� D�
��־,K�T�	�91QB�<D�,��B��I�g�.!?��!"i8D��悀]c�ݫ��?��lI��7D�\xU(ĭO�D�+��<��w�7D�� z�ďx�!9�ǂ�x�PdA"O�P���6�R Jcg��0��a�"O�U1��ٓ��X��fY��"O^��� wN��,� @m��#t"Op�e ��5l
��+�^���"Or���H0Z[��R��Z2(��3t"O�Ms���0�jݹe� �n؜�#�"O.�����9<ExvF؎o��TH�"O�8ĩ�u��[�DM�i��� #"O�ɛ�-ˊ!�r�۪)��`1"O�bt�A�1Kڹ���ʓ%�����"O]҂�+U`�l����)��3%"Oȡ@��7b�$`s"�P[D��i6"OTI1R���T��B�|���"O���c��>��9���5�`��"On�f�[����I�
�hX@��"O�� H�-� ��6)��dB:��6"OF��`��2Hv�a#��=B��iZ"O�`#6�ߚQ�����oº:����"O�er���05��x��+9�ޝYA"OhW.�IF���-�4v%���e"O��+VJ]�_/"M���$Q�"O�XHQi��*KXQ��H
R���t"O����w��E��[)��=�"O6a�F���ZU��'C1� ���"Ov"�"�!}�e�  �$�tl�"O�x,�t+��ǂZIfT[8�!�ҏ7��#Ԭ�>A�!��ͯ<�!�܇p����iS".� ��ׅ�!�:5!b ���]�4��c�%��'$Բ��ʲX����I	�Xvl��
�'��9�+P����:M����'ҕ��C2���K"2�T���'����A�936�	���*�6,��'�|ʃ)N2��J�ɖ"rfy�'堘Y���G���g������'c��ǭŀd8aq抉��
�Z�'���;2a�a
y�5/��T�.9�
�'
p�a�L!6��{��F#��
�'�h�s�ыc1x��� ,�B��	�'(rdRE���������S�I
�'|�}8҈�-+�ڤ�'S�!��@�	�'`�
#���a��<��Dq,Q�	�'�bm����Pm���p��'),J���'P�q�fhI=�� � ]�|��'�]�'�	�V���١d���i*�'��H����)'@�i�.m��I�'%¨cP#�(6�>[(��w����'k���M6+,����ѷh�uB�'�12��ϛ2������ڤ�	�'V�q�.�af-�D����~���'-��4LZ�s-:� ǌ)�0���'{6�rqF� 0�!�D��9)� �@
�'M��R��,V��m��a�<�t�C	�'\���-O Zۄ�H4LG#
��@��'�4ʰ��^�i�3.�}H���'04X�5.�	R�nx�g�V)*׎	��'ʀ�J$
D�
n��(�`M�%�-�	�'�PR'�â[L�����ž!~�s�'�%��!�+">euMA�&"}h�'�H�ʵ�/)vؙCSw~pz�'�F4��݄,{���e�DL��'�ViqT5�6H���U�6����'�dB�-���5
!'섥���� p����+U���D^k����F"O�0G�`+dU��DZ;Z�D�b�"O<�Xd�8Mf�,�֣�v��p��"O���kL`J�|9��Qu��B"O��QЄơu���Y��`� ���"ON�����N���b&�X�~<X�"OT���I��
�����j��!!�"OE����\X�$YT��;c�6R�"O�]"��C�<uk�3:�d���"Op(;�����"1 �*F_��U��"OL���C�?#>F��bÝ�0ĭJe"O���O�(q��1��"%����"O�GN��ˬ��� 0n�v�0�"O8�*
ɍ>$���pB�^����"OJ��bA�*Ǌ�Y�.�!gѦ�8�"OL��3���D��	�Ѭ��z����"O~0G-�
Z_z�k7�'c��L��"O½p�f
�|n�&Ǌ(6����"O���� ,~�1B�%�%Kl~�"ONISc�ǌ'�\I2�T�,el�Q3"O�d���I���q�6Ώ�e����q"O�(;&�+F�L��+�r���c"O�����B%_��(�Ӓ9Z�ȣ"OTLK姕�X@l<1p�]�$Q��hB"O=ZR)�H-љ& 6ך0�B"O�E{��B<�y�% ��q9�"O��+�̗�T���oP�a1�"O��"�/#�2$�#j�<,cH�j0"O��Y�Ē�s���e	S�6���CD"O:,��-�f;8����=:*	�"OԴh�L(aӲ���fK+Y�p "O��Ҕ�7\Ř!SP�ұA:4�zu"Of�qTeY3\ވȀ5��0yΰ@+�"O��c�)WC��iJ�$Ū[����"OԄ��*�"�����#џ'�"X*�"Of��fe� �=Ec��#��p`�"O$Q@C��)=���\�)�V��t"O^��� L}�6��T�O�?���
�"O���M� Cl�c�"߭�<5�4"O��j ҫA��,���سkX�Xن"O�|yq(��"��}ȵ��?c��}��"OZT��ʘ{F�$��^��`�"O�̣э(��m�t�D�T�j\��"O�,�F�$��h2E�!V���"O�����?�P����']�`�ʗ"O�����F�a���B��@b�i
�"O }���?�Q)�I�C��!�"Of�@�"��~�6���I�F���0�"O�p�S/)8�6)9ba_�hNyJT"O�p;5j�+[� !)S`H���"Of��6&��D�qi<bE^� �"O�T�F�� +����H��Lx�"O�sB1S���0&V�%�B=I�"OF�2r	�2�V@a��Ϲ{��ದ"OB��A 
  ��   �  C  �  �  �*  _6  %B  �M  iY  'e  �p  @|  %�   �  ؗ  ۞  �  _�  ��  �  _�  ��  ��  ��  �  K�  ��  R�  ��  D�  � �  � Y �! ( 2 �8 +? <G �M \T �Z �` �c  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+q��62\���<4�d5h��'�B�'���'	�'/�'�B�'��x�.Z ?܎Yf��0d�tx��'��'���'�"�'��'���'�nY�5��B��0��g��ծ�pW�'l��'C�'���'���'���'b��i���8��}��dK�� �C�'1��'W��'�B�'���'���'?�%�����غs�9
lk��'A��'l��'B�'��' "�'O���ek�92�lu���D�+��'�"�'\�'���'��'B�'�n$Q&菷U�~�
�"��]x#�'���'��'u��'�r�'���'� �H�N$!��y;�Ã+K�f�0�'���'$��'dR�'���'���'�Fx-Q@�蒠�6/X��o
�?���?i��?Y���?Y��?���?�Po�^}��� �	\V�p�'F��?��?���?Q���?���?!���?auj+2��!� :D�|Hʗ��!�?	���?���?y��?���?���?y��ь�����/�&8CTtꖢH��?����?Y��?����6��O����O��DB(Hc���$��[��$�E/U��b���O����OX���Ov���O�!lZڟ��	�P��H���L�!�"��~�-O���<�|�iӸT���_�6HF�Z��
/��A( �C-)l�	9�M����y��'�����"қy����g2-m��Z��'9�훑u*�f���̧ca���~�6DI�o�P�YfJ�z�����ND��?�*O��}2'�X.xȝ�����\����X�jƛ��!��'���nz�]8�"D�O���3CmX1'�̻%��՟����<a�O1�i��u����9o���3B��\;�슰�"����<���':$F{�O����>��&_*�xk��Y��y�S�t$�0�4�4T�<��f�5KQ.z��N����	��A���'8��?y��y�Y�ЫIX�cHp�s`䆵]�>L�p�6?1�T�q0�j�'T�����?�ѐpI�Q�Z�$s.qR�����D�<y�S��yB@�#�B�a4�Iy�Ą �y��l�ƽP3���b�4����T!�#^��rd���k�f!z�$�yB�'�2�'߸r��i����|��O�x!*�m�E]Z����gA�4HTb�IBy�O1��'��'��ݥk�, D���-��H�銙r�ɽ�M��"�?����?N~��JGX��7h�|l��q�V!{CҠ T��2ش?1��(��i� ��B��;.��q��ѭng^��$,��[>�w���~����:3��ɓl���S$��	-Ix��P)L�9=(T�I韬�IܟD�i>��'B�6-�<>���F�H���#��,ƚ@(V"�%����ɦm�?y!R�4�ش�&�}� � J"l2`sg 3ܼ;�n8f��6.?Y󎟺�*��#���}��]	%�� ����6�� 	0F��I�������h�	ڟl�IH��eq�i�@ۺ,o�	��*B�S�A��?���q�6-1��I��MCO>�T�������4�)�x(I��-N��'L�7-�Ӧ��b�x�on~��I�@;נ�'m*:�B�MO؜�� ���P�VQ�,i۴��4�`���O$��>N���fo	4˖LQ���h�����O �����V�'�r�'@RS>���D��1���]O��q�1?�7S�(�IƦ�RL>�O`C⇒TjZ�iQCǩ}��@���-6�<	ꇠU���d��֩�O�Ġ)O�ѐ�y����e�dDIW��W�,���O��d�O��)�<�u�i��	cŇ�F�RI�%�>����	�����?Yw�i��O�D�'K����DMfu���J.�}Q1E�W`\6�즭r6�\Ӧ��'@`�o^�?U������K�)��$�sH��%��	Ϧ��'2�'3��'��'���?.�ҘieȎ���s��G�1��4,��)/O��?���O�!nz�m�珄2j2����/\�`�Hq��?۴4ɧ�'�(�4�y2�9!�1��,��V|�5���y!�9�4U�I�\��	�M�.O�	�OBaj��V�=@����́�CF�ya5F�O^�d�O*���<��i����f�'��'���:g+ƣX!H"F��G{����dU}b�f��l��ē1���Y�ala�&V�@�������Q~�o��p�`�@�-��D�ںc6��Oxi�@[����㗬�D�l[U�py����?����?����h��^����1�x�ؐD��t������M�G��ϟ��	��M��w�n���;#�]�����DQ�'�6m���Q`ݴm�(�ݴ��$�zJ��'V�x5�F�%_�pW�K�a���1S��<�ҹi^�i>���Ɵ�I䟀�I�j���C���i���"�Ȗ�rTT�'�.7�M�e�r��O���1�9OT�a�.v��($DA�[������D}r�q��l�=��S�'m��|ad�Y5͠�!�ɒ�ZH�"�冤u��%�'�$�*�I̟4K�Q���ش��DD�E������@��l���N�8�8�$�O��d�O��4���<_����	w b�?�^�p�Q�������8�y$u���{�O��o��MKղi��}B�*�'�^P�`��cҬQ��ƛ1O�����L�#(�k�ղCN�OcP�=� d!�%Ȋ��2�� ��N�l@��?O��$�O`���O���OH����Ӊh�Xh@֊�i�QȐ��~���D�O���Ԧ�#�*�ݟ���ܟ�'���"*P1H%����(_0,p5H��K��M#.Oj�mZ3�M�'�@�ܴ����Z�`ٳ�ϙ3Z��G��y�j��qER=�?i���O���M�����'"�'��I�wa!C�f|��X+W�^����'vRX��Z�42Q�����?�������\e� �LM�I�Ҡ1��������?A�O��$l�Z8oZB�'Bq����H�lRs�� ؘa���v�8�W��a~��a�=���'o��Iğ杘}8� ���A�>�@�bЯ^�+��q�	���$�i>IQ-^A	�4�'Q~7͖;h6�q�ƨE�c�phUF�41tc�<�����?�(O�9mZ|�jT[��88r��4�Xyp8���4mɛ(ġzě���|K�-U�9>���~�qi�7H�%�A�ީr4*P(��K"��Y�����4���,����d�O`X�X%�,Yz�vO�,`�ĩ6m�����>_(���O��i��'M4˓�?ͻ:��dcF� �PX���x�+��iAj6��Ȧ)���O�x#��i���k���vm�4���	4��O��č0b�q�LSJʓ1Û�P���ޟj��O/R�L�C'�*`r6�xT	���Iϟ��	AyR|�L�o�O�d�O:��"
�0��5�ti�40T.�O�ʓ�?	�P�D��4Tϛf�rӀ�z0���paA;Br�\
 .	8@R��'���Ta[,
����Oͭ��n�$���?�0%Qg	x4�Sj�^y~Рw�N��?���?����?��	��\�ɹ�ztIc,�/X�0 �aE�b��ɘ�M3Ca_�?����?q����4��/U�`@փ�	~�i ��\���Ʀ1*ٴC؛�
մM������v!�<��t���Y�B(��wa6K�BR:�0�A��� �	��M++O�I�OP���O���O��)\���@I���TdC��<q��iA2���B�b�'����p;��'��M�%^�
�S���	=.9�g�RH�U��vHr�Rhm��H�B��l^O�Lhx��ͽUl.�&,�+ ^8u8���|PSmؼV�)�Iy"am��� kj@2�B�;f �\���ƨJ�d����?���?��|�/O>t�I2p���=^̱���H�U��rB�}�Ĉ�!�?��Z���I����4Q��BD Iz<��TiUjF���l�?�MK�O�m��P���J?e�Xw�IGp�x�FI�&*nxӢ�C��yr�'�2�'���'���Ӆ6Wؑѧ���MF��;�O�cP��d�O��릙��)�qyB�o��O���R���Vƪ���"�~�p�X�i�I�MÕ����眒N��&3OF� ��H)'Ģ(Q����Zl~�)���S�,���IZ��P���.}��Ryr�'R�'jb@Q�w�
�;��^�z'z�`���i%2�'[���M�6 ��<���?)(� ��vF6���G�0}iVH�7����+O ��e�v`'��'Kly�G�B�"��C����,�ʰD�k�(L�"��~�O��q��<~�'a�-³"�l	��C�ҹ\���$�'��'�R���O���Ms�āY ����9Q�*�:�L%�ƌ�'7M0��*���S�Ar ��"2�å���`�!
5b��M��i芁�Q�i���v0u�%�O��'#� AQ .e�\(P�mYmB�͓��d�O��d�O���O���|2��Ʒu\�$�5h�?0G�Ź񧜜j�����y"�'>"���'��6=�"Xq�W�$'�!S�]�_�U�D&J���͒O1����!q���I�s0���ą�Π�2+�:1N��ɿ�H���'�¬'�蔧���'�2������r�\0��4���'�R�'�"]�d�޴X+Y����?����5h�a˭b|`9��ƻ�C��<���?�M<)ck�?<x,�'�^ 8��:���k~RN�p���&c[0Y-�Oj���I5Yd"	2m 4��Bk@��d�#�i�K�"�'�r�'���(
7�M;z���s�[�6U��JQ��\�ݴL�$����?�q�i��O�N��3%Ba�Ei${�E�Ȉ^~�$������M��m�M��O�I����S���QŐ���ԕOp�ac���C�z�O���?	���?����?��Rqa��P�*�1���H2�),O&�o����T�����j�s�Q�	�=}�p�R��pk�����N=����Ԧ�*���ŞK�\+BMïzm�Xfo��U�������-O�u�P��?�0�>���<AF�Ϩu��7�<q�|9��j��?!���?Q��?�'��$���	ccm��dƇՐu80���;UlX��럐�4��'Jʓ�?1���M���W?N82.R��2�(p�	�#ڀհ�4��d�!_,������������� c���%Ɂh��,	�Ɓ�'��'��''��'h�P���Qd�(8�!t�a�R��O���O� o�u���|.�� ��4��$��hN�u°�й+��O\o�
�?�(��lZs~b.�� 7^8XsIA"�Ju�e�՘~��"Ɵ�!b�|�R�\���T�	̟p�`��^ٞq2��W4_���x��ޟ��Ioy�`y�\`�B��Op�D�Oz�'`�z����)+����ذ\���'�Z�l�*�O$O����`<I��ц{�$x���h��8G��<)���G
�7z�z������O�U�K>�c2#�JG`�7Rp� .���?!���?���?�|:)O�Hn�?af�	1���_خ$��C�!H���vCV[y�F~�
�d��Oao�m�h�
�D�x�n�1�
�J�.$�޴�?q!�_��Mc�'�"*D�}��y�-��� �I�ƿE4�ݪ��*cB�!0Obʓ�?a��?����?Q�����-��\�sH�'���7%����oڢz*��'a��)�¦睙V�$릆_V3"����F����{�4"ߛf�'��)�әY�Dm��<)@ON~�N�%A�D�{���<ɧ(֭@X�dW?����4����җH��M�#�I(t�VE0o�%;���D�O���O�˓\����/f�"�'��@g%��"�؆W�:��fO�V�?	�S��ڴ=����' ��*_Jt������"SBߴy���-(N��@o�#W����|�q��O��S��?�J�C���qH ��%��¶T����?q���?9��h���dZ��~�������� vI.���@�qړ%VSy2�m���]�YO�y�7��~z
q�'O�	����M�ǿiJ�OG��v��<q����de�\�FI��g�����ae��]F�T&�������'���'Z��'L�0jpjўVf�-�Y�Ԛ���ݦ�S�J؟����%?�ɬV'.ْ�Ә���4�[vd�X�O�l��Ms���>���,�N�Z(8�C��P�T,�¡\.MZ��d/&?q�E�O�*��]������F�
|Ke�#n#�l��L�v� ���O���O��4�,ʓ!��)��y2�E#��uhZ� �5
��y�i~�㟨��O��m��M�Ӳi>ΐ�����"_d �'T$m����	xț���h�� �3,���i��^�����t��K�톰^�Z���>O����O��d�O��d�Oj�?9)"lY�N4�M],&H,�W}��	�BشJj���'}�6M0�ā<\��D8`@��w�4��59�
�'�h�4՛�OX����i��Iy���'���v��䇙�f�-b�Qq���{�	Ey�O'��'�Nޑc���</94��ҡ9���'9���M;�G�q~�')�S�>s��9��N�Cpj�+E�U�c���t��I��M��iqLO��#O��I��
�P��SF�ԋ];�p0��(;����#?ͧGwV��ԇ��>��ñ���)G�yЂ�҉O�"�H��?1���?Y�S�'����?Miڈu����F��8��r��
�˓d����$�l}�Ns�j@z+�r�9r�L�dߞ�֥�䟸lZ8eܘ�l�p~R�E&9��ӱo��	n�#BJ@�|} `�[ -���py��'�R�'���'("[>A#g�S�L+���|ɤ�'!��M��&K��?���?YJ~�'盞w������:d*�jV;^�� �{�����e�)擉G��m�<����h���!*�Z�&��ˇ�<���̀�L���+�䓔�d�O��d1(�b��1B"���I�?�2���O��D�Oʓ["��C�V��'�bF_9 ���K��L��X��Сx`�O~�'-�7͍� %�pz��Ead��Bϫ$)*���8?2F�\�� �	�6��Q���䏶�?)��2U�� ⭝�|Ip���Ջ�?���?Q���?�����O�4�&��+[�%S4�Պ2r$ԃ�!�O��oچ҄���ğh[�4���y�Β�:�Nh� ҆ڤ|c�Ō+�y��dӄL�	Ԧٸca�ڦ��'ޠ\aSdL�?u��*���и���	���aD#i��'��I����	ޟt��ܟH�ii���?�v9�נ�6]~����<A��ie����')r�'��O+b�'q�,q!1��}�Z�0)��-6b�	�v��O�O1����m!a��*��<&>p�2�	~@j6Ϲ<����+m��Dؼ�����٣s~���C��W�|؉�n¾(���$�O��D�O��4��ʓ2��*Fd�2�i�p��L�#uRl)�#��y"�wӐ��­O��n��?��4w<@��:��XS ��B���P"�M�Mc�O��⅜�:�'����T��6F��������d��0O��D�O`���Ox���O��?�@�G�#F� J�{QыS؟L�Iϟp�ݴN��u�O�7m#�D�PDn�#@�;{( ��G�`6t%���4T��O��0���ig��-!;��؆h��O;T��A����D(`�@l�CK�IIy�O���'	d�xov,��f����k��K2�'"剣�MK���?	���?�-�z�s�C�+\�!�,�~خ�U���q�O.nZ��?�L<ͧ�J�2=��3%*���BT&��\� "��06Q�Ѳ-Of�i��?�F�?��U�+V	 !@�c��+@��]S
���OT��OH���<��irjB�$�h4h���B"���A!I ���'��7�$�	���i�.D�3��'l��"&'̬lv�z�aŦ�ܴl�Q�4�yr�'�81c#���?5��[�S%�V#T��%�
�DM�P�Ghc�d�'q��'�B�'���'Y�,�@q�� LLq ���X��c�,ţaD�O����O��ɶ|Γ�?�;.gH�	������6�K�p�z��0�i��$�>	��|�����S럹�M��'q� ��˷�P�Y�ł�j���'M��(�͕ڟx�v�|�]�X��֟�� &�I��t�ȼK�j!n�����Iß`��tyb�z�ZP��O����Od���hͼ��IR���"t����&��2��d���e�����-�Z���K�~}<� � �w����?i��͌�\C���d��n�C��>��Dmc�4ڣO�!t���E���@�$�O����O��d+ڧ�?��JU$OT��X1�ȘY&,a���?y�i�,	s�'mB�u�Z����d<��*ñ(`��0.�!UVf�Iަ5�ڴ�6�Mʛ�2O��$��	�0���L2�  ���Q)C��P"�����J)�D�<Y���?Q���?���?��DÙzАPcR:F 楫�+���$Wݦq+f]ܟ�����8&?���.rkd���Bр3�l�B4-��sb�(�O��m���?!O<ͧ�b�'4!
-	Pf�scr��6I^>^D��㨏Ge~�q-Ot����?Y��<���<�R���sބ;gJ��_1�	�pi���?����?I��?�'��DSݦ!�be��<q&m��S�)%%J�k�~�kW�z�4�ٴ��'�j�rԛ���O�7ԗ�x�€ͣ-?H��b� a��g�eӨ������"C��,;��YIyr�O�G ܶ@��������Y8�fO��yR�'�2�'{��'�R�)-0zx)��ʬW! 噃iQ-)�Z���O���VϦ]�sas>��ɹ�M�M>��ǓK����2O\�A�bߩ|��'�6mX˦)��i�.o�<A����=��
�}ڨ:AhϺ>(��Q���+@���H!������O��$�O �DЩ�"t(��{mtزF��E�r�D�O��n��̄@��'1B^>� �R�P]^QL'i�XԐ'�$?!�]�T�ߴcf��l4�?m0�
�I�Zh�v�	6X�xa��s2 ,� E
l}���|�T��O�HIH>�,њ`��k �^�7$�Ay�'Ɂ�?Y���?	���?�|�+O�,n��C���#D/۫v���`A�/M��1�Ϟy��c�n㟬ɨOlZUl$���G�
2-Z|�Rh��uΕ@ݴכ�k<$̛v����N��3*���~z��S�Z��]����2�v	���<�-O����Of�D�O��$�O�ʧ��ko�t!��<K�%3��i�~����'��'2�Obb|��n 9���7��<K�9�)��J�ƕo��Mkx��T�SAU�8O*1�S�[@i"w!Nx�*7O��ؐf���?��g*��<�'�?���ɣA�Va�5�F@�� �?���?������Ҧ����_yr�'W��$��A�~���`+=�89�����f}"�aӲ�l��ē����"�A�]� �,��T9J��'&��r��_<r�`����џ�`��'���Y��,0�&t�V�VPƤ��7�'��'���'��>����gl�$X1�H�g��1���cƥ�	��M+���:�?	�)ɛ��4�F�R�H�A�@�<_��s�3O��lZ>�?9�4Lf��ٴ����D_����'?�<���Ʊk`�rgG�N��ru�*�ĩ<����?!���?����?Q����C��!&y�O
��d�Ʀ�"g���t��ß<'?�I�p��i�[L�$�!��rK�u�O��nZ��?1O<ͧ����I���ւLZ���#� >m� +b�$�@]�.O��Q�엉�?�u3�d�<9r�Kh���'#��g���JgCK��?9��?y��?�'���Y����П�D���zD�a�¤�7��V#����ߴ��'����?���M���u�XKgKB�P�t���`F�,�۴�yR�'/,�b��?�
Z������E�F�еPZ���R�Z��Q�ѭ~�X�	ğ(����	����J��'K����0m�<&�h��
��?���?�ôi�I��O��z���O&��U���$�H�*��E[.���n�k��;�M�g�i%�+�^��f<O~��B+#Eƕ1��]0TBmP]ufy�b.��?qE!*���<����?)���?`jO�#b|�J��9��y�3�?�����S���Wߟ|�Iޟ��ON��Wj�
�@����������O��'o�7�U���$��'g��qd��/w���G��%K�@ց�U v�N���4�b@���0��O�$��L��" :�*A(��\$��O����Of���O1�.�9M�)]�%�Ri�u损|�R|�#胺z���R��'e��e�㟨J�O
�m�$3��A�NǖB�=�2�`��YPڴ0���LУu�Ɩ��Q4G�C ���~B�AֆQ��xS��k�˒��<���?����?���?����?1�⚐3��N#�,� �@B+ir\���-՚t�y�����?���?��i��'�2^��N�K?�K�CM�Z3<\1��H�?��426�U"��Y��y*���d�-S��7mk� ��k�q#ݨԩD�J{�a|��W�PK�"��@�	Ey�OG�dܯ)�:ap�$9 ��ji��'k��'*�I��M;����<I��?��lť"�HK�ܞO��bT	���'<��BǛ�Hh�x8%�����,��x��@�02�H�?<�'m�B�5�JT��,�7��埲���h�
��Φ@��8
�zP.lA��Y-Ӣ��O����O���*ڧ�?Y�ẺeJ���͝�(r�Ip�,�?��iw���&�'��k����]
^q�I��@�0�d�2/�J"��ğ�m��M�d��MK�O�A� �%��SMU%\	��+�7�:��*^UWV�O<��|B���?���?a�I�*Պ ̅�3�b��Ǭޥ{=|=�-O��n�&�,��I�h�	X�s���yp�(Ku��d��P������D��aY�4np���O�Ji�'�L�`Q�5�*>΄� �#+ ��*�O�	CE����?AU(;��<�SF�5�0�!)�'�j(Au�;�?I��?A��?�'��d��ө�ޟp�ZV�lk��lұ�cC6�<��^����?9�]��pٴmۛfAj�pɡ�ÖC�^|��&2�M!��
Y�~7|�X�	�	�d��3�O������;:N&h����*��� ��C=9�DUΓ�?����?����?�����O�
812�N�G��y!��H��O����I`d,?	�i!�'�̭�d挺DdH{X{3dPK������,��Fm��)X�k�7m"?�d�g�? �������<� � �@��v��;��?��- �$�<�'�?����?�%�+#Z���򂀾E��0��͜ �?a�����!���ڟ�	��t�OT�����Z�d�p��ϟ1W�T@�O���'��6�Z�%��R�����d\�9�b,;F������.W����ĵ��4��D����̓O�d�'D؉��!sN���U&�O��d�O����O1��ʓÛ�Ǆ�-ޔ ��B�]�fRbG#���Ң�'(2�v���L��O�o�:|x����i�3)��t1*C�En(���M����M+�OpX@������<!��׎mEl��!6g������<�.O��D�O~���O����O��')�H!�.�
�y)`	
�xn&s�i�R�QA�'��'Y�Om��'-V%2���aO�帠ϟ�N���o�"�?9H<�|:�!?�MS�'H���F'׺@Ä�W�v@ !��'m����l��k��|�\� �	˟ ��ፊ}".�9S!�n\�(H�F�֟�	؟���Ey�wӀ���G�O&��OR���ND�F�.5��� "x�#�%�I(��DP��H��ē�&i��h�TȊ�JS�e����'��� 5M��oȹѳ��������#�'���1O	h�T��牌�S;�j��'���'��'��>��r\��Qb�5�ι@B�Қ7yB����M����9�?Q�&㛆�4�vU��E�b�dę׃:,�r:O4=m��?Y�4Ns�4�ش��D�:,����w]p��a��WD�|�"�-���S/.���<���?A��?����?ys��>:!�[G�8)vb���O�6��_ͦ	�E�My��'��O^2B�)Oxpn�bd�� "b�h�h�#��F�O`O1�t���k���uz�/�>R^2�ܮ`!�����<I�J~����:����d2h�t�P���#m�b��������O����O��4���#w��А'��^�^:����!8{������ry�jcӰ�p�Ovho���?��44���"c[�[��	�����$;&@��M+�OX�˗��$�z��?����
*�e�B��.�5av��V;O����O����On���O&�?��b��z��h���sG��ٟ@��ɟd�۴l+"��'�?ᴶi[�'H|{p!��1�pj�H�$�9+��!���O���O��Ԋ�i���/���͘==�X<���Q�hTr(�߼�����䓙���O>�$�O���r�+.�e�1���e��ǟ��I~yr#i��
E��O���Oʧi��8@��'��i1.��T�d�'��d�6k�OO�S"e�މR1m�4t9���r���m�n<R�] ���AׂX}y�O��Ib��'�B@����"�٢��~���v�'R�'�����O��ɼ�M@FXOA���$�R=$�nU���Y<u���,O�oZD��!�����MKe��5��P��\5C�JM��o�Rb�i�2d ײiO�IK���%�O��|�'�ީaOS�X�|����U�&��K�'���8�I�`�����Ic����rX$9DI�B $���T#�6��+�.���O�d"���Or�mzޅ�B��/@�|Q��Қ^n� �N �M�յiW�O1��,K�Cp���IZ2����K��48tL�<Z��.>D���p�'ʹ�'�������'�2	�3n��M���LR�if�'\"�'lbV��!�4qL��z��?i��r�}�rhU�r�����oڃ	��`�2
�<!��M˱�x�%H\�b!O��w� c�ֽ��䞤2-�p;deK�~#1��|��{#��$ǸP�v��ƕ4^�4��A�žN�(�d�O�D�O �$"ڧ�?)4�>j3@Qb7%\\(ma��?w�i������'#R�l����'X<x� ����w�h�0*�H4Z�I��M��i� 6�W�`6$?�G�h�f��	�ѩ�B�
�+��٩%���I>1)O�i�Od��O���O�P����;OO�r�ܪ
��A�	�<ҾiHĸ���O���.�9OZ����Խ>I�5���Ӱk*�Б���X}R�y��o���|"����Ƥ� Lv����2Ԓ���T�n���a!V[~�]��y�ɮ6"�'���R�nlI���f�:ADGB�_��H�	ş$�I��i>�':�7�hf����%y��g�N��a󪚀h�������i�?9�_�h2ڴJB�i*�`�j˖ Wb�1(մM3�	tK��b�֑��`�(��	5��$�G��߁�c�'%��0��u4aC�ko�|����������I�T�����+�,,�����:bHQ�`g��?����?qb�i�dY�˟�8l�џ��'��I� ϕ�b$���B�A��ъ �8�dĦ9ߴ�����MK�'#Bʘ?��h������
�8� 8�P�Jϟ8z�|R�|����Ο���GN= m`G�[d�C��<��Syb�dӴ��1g�<����i��S����eP�5���8.@�Ɍ�������������|���?��(�4�$�a�ʷx��qa�-P	4ƶ�Ѧ�����D�� k�	?D�O�)�0�U�?������Y5Uh�H!q�O��$�O���O1���a�V��>W����e�\�9C���Fm��z%�'YR'pӚ�;�OZohن�YuI�]��@M�n�1��4%��6�'n��f?O�D�3J�����b��w����� �:0O6�1V�ٴ�r�ϓ����O|���O��d�O����|��2DJ⬒��ښ7�dJ��6A���U��'bR���'�r7=�8	�bO�9r�$LD�w\�<�p�[�	*����|��'�JQ���M۞�� �Y[tfT�CɈh5인Y����;OJ��l7�?9�*2�D�<���?�D�^4%�Q�e+K2t:��H(�?���?!����d���I�f���X��� � ��D%:'��H�)���`�2�	+�MKS�i�S���B��99=��0(�G;�Yi��p�x���𨳐Cи%2�bV��Oxdj�L���BWƎ&�t\㥍C�=������?����?���h�>�$U7{��80 �ZbĜȠ�K44�@�ČҦ%���8?ɰ�in�O�.
�4I8�AvA�.����*^�?�ܦ�!�4;e��-J-%�V5O���I+�����'3I�h�C޶sp��)A W�u���ʷ*���<�'�?����?����?	P/IY�!���@$���[4C����$Dߦ���c|�`���X$?�	���J�ٸ|V�au''1�3��D�O^7��X�韼�	���-S��)p(���Ɯ6���͜oؾ��P��d��&�9��FN�IQyre��G9
̃4��halLq7�WlR�'T��'��O�I�M#F�ƫ�?7%�g��`3��]�wʂ�@��?��i�O���'��7m���Dm�^V���Q�D@s��őp����	
9t�7�%?��%���I��ҘϿ��-�i�m����Us�BV
��<����?���?Y��?)�����[1vAٲ�@y�fԈƥ��$HB�'��n� R�4�l�dM���&�t�T�����"G����u���A'��!��O�O��k�0^�f��d���֘5#�$9PNL0�zEp��� G���q��'�� &��'���'4b�'�(\�A∂8���,g����'�P�Tbܴ2ޞ��(O�ĵ|��$�E��}z�
A��N�8i�~�!�>90�iښ�3�?�"`N�y�TlP�9����(n�tx���H�>喧�t@I����|bn�{`dS�NL�7�rh)!�W�c���'�R�'c��4]�T�ߴl�$�����>DTh(@7e�:�|��taʪ��dJզ��?7U����4)d���+��0ًCJʳ*ઉ�U�i�x7�_�U7m:?��K���>�	+�Ԡ����Q��t��udX��y�]����֟������I����O�P8���U�Z[ވi��[��C�mӬ��G�O��$�O�����DH���݃@N6p�pE@�W����e���$���4>���5��	ɓ}��7�s� �S$n�XmHB.�7�6I�p�P�ƁU %��i�D�@y�O/X�)����O ?F>�x4o�1<�R�'���'�剩�Mk2���?a���?���� ��Y��\o>�Ec��H���'��� ���gӬ�$�؁�/��Y��H[q�<E0@It� ���l(hK+�|������O(���D��3w,V?6����/[�BՒ���?����?a���h��ė&%w�M��<t_�RV�[�C�\�d���=���KUy�sӌ��]�ecέXcK��W~p11�@�a�b���M��iS2Q8~�����X1Q��0`���眠a�J]�ri�2�>@����5WuF&�P����'52�'�R�'�Q�4��t쀰u���q[؉X]���ٴ�f�����?�����'�?�D��
|��+Rk��Y���C��"�I��M���'����O�� �e*�l@�e�i࢜HfKZ6��B�_���r-�*j�
l�	jyb*CV{��kU�×[���T�X�y�����\��̟�[yBxӞ9� O�OjP6L܏���8 ��er��>O��l�S��t?�	�M���'�L�=_p�;F�Ĺr"A�1G�	l��0!�i�����e{U�O�&?	���K85�F�L	[ڎ��@�=��	ß�������Iʟl���Oc�\;�mI�$f�I��J%W�0��s�'���'� 6�xp��kț��|�b��۪lb�O�!vP����*2+O,�l�*�?��7���n�W~�b��a�R	�CKZ�!ĩ��PRTq�G�ӟt0$�|�W��	��	؟�3��՜`=`����0qS�I����Ify�Ge��0����O4�$�O��'J(�X
�V:�L�!�3k�u�'��Si�FE�O�O�S�C��T�탚wq�yQ�ǂ�rw"�8����z�ǘEy�Ok>��Ic_�'�|(V`�q�V�%��0
!n��'��',b�O:�0�M�瀋�Tb��U*"�(9�p��7��P��?���i�O�p�'��7m���Qk״o�B��f�<���O�7���6M#?�2/U-Q֠�隁���x�ɻ% �@�N��`�<f8�D�<1��?��?���?A/����I��bܩ)d(طG���!]��D�C���	՟l'?�ɻ�MϻV�x�Ԃ�'��H�!oT�R�d�h��i�^6��|�)�l��m��<I�h�
\C@�^��&)��<Iq��5	��$��䓈�4�����L8Lx8E Y1,�Ęh�T�/K����O��D�Ov˓Z�F�H�zA��'Cǂ�i��p6��,s�h��$b��s�O$U�'��6m�ۦ1�M<��̥k�܄p`��Dd�DOZA~� .zE�}�t����O_�a���1�Nų\�]���i�x��[����'��'�2����J�n��L�p	9���43�`�Q�^��4ufr�.O<nZK�Ӽ��T���*���+c� ���<A6�i��6͙����&�DĦu�'ˤAB�A�?�
b�K#��y[����R� P� $� 1�'��i>�����T�	ן���;�vQ��$E	jpH���� >��ȗ' 7�G�V]�d�O>��$�9O���⥖�aD0p�B��it��`��[}"�aӴlm����S�'O�L�� <i�5H����|+%@Y�<�ZH
�)�Y��ɳ ��݈d�'�>�%�Д'p*@;��({>j�H�՚8BE$�'A�'�b���U�|K�4}  ��8,��@g��a��I�!��:~��͓)0���d�M}�ijӪ�m�M�%���+�(�0��ݸSJ1���k޴��DN�P\P���øO�wNqe�X+F)�Ir� ��a��yB�'�R�'0�'O2�IͬW��$�6e��:h�NZ!Y`���O����Yr/l>e��6�MsI>��DY� �!��G��ZE�\�{H�'�r7m��I�	;Z7-3?��DʄLR��w���I��'��� ���O0�J>(O����O����O�}�V�X7d��l�r�Z .Ŭ�2s��O���<)��i۴D"��'D��'���U/ݜu���хL�M�a��I=�M��'�������0Q�a�cA�O�B������D	�E��(%�5[d)�<�'x����%��Kt�����=NZ�l�H�r������?���?��Ş���֦�pDС&iQ6Ĝ�tTb���훲b�'�7�=�I���DE�EA2쏕�`y�3&��\�6�Se�=�M��ir刖�i��$�O�h����ڴI�<�Vl��]�B��&��3E�iZ����<�-O���O����O����Of�'&W��X%� ������X�h��3�i/.dKB�'���'M�O�@u��΋�'|��t.U�n��a#����,�|�l��?�H<�'���'H��H��4�y"f��Hs��@H�w����f��yRG������k%�'��	ɟ8���/xv ��J�=L��@�Y*]���	ٟ`��ş̖'Wv6����&�D�OP���1t!x��������P$`�>����O4,l��?�O<q�FK)[���h0J�2v?t���D��<���4)� Z�9NL�3/Op�)��?�q��O���s� �Q*Ď3e��;�Oz���O8��Oꓟ�ä	U���ښg��Pb�]�k&�R�o�)^ˈ���uDMğ����	gy��y��Z�q��K���4Z�
�
�*��y���^�n���)�ܦ��'�
��H��?�"ލ"�t(�7+Z��Ha����.a!�'��i>��័�������"'�ܱz@NM*LaN(ТJ+^�@�'��7���:TR���ON��5���O,\��\4z�D�3�^�&S��T�Tty"�'|J~�`�A�M���%�;\@1������ݣB+����d�3;����O�˓d ����:g��TI����d�VLY��?����?���|�,O0�o�32s����6|؀��g\�C�5�ca �Xǆl��6�M��F�>i��i�d�D�v�s�g�e���P+�+ڐ��ь�ze�7�2?a�BW3Q������ܿ���WD��Ř���.p�ȓ`�N�<I���?���?1���?!���@��p����0�K	[Q2ؓ"�,R�'�B�k���@�5�H�d֦�%����d�8P��ӿHy�q�5��ē���k�O��d"E����w(h�̌`6�(hEN��sg��f쪶�'� �'��'���'K��'�H��f��x�T��3�W�
}q�'�B]��
�46�nm���?A����Q�D��pb�� ��i�#��I�����������S�dj�)7�p̉��Ƿ3װa�R�A�`���pc�R0N|@��Y��S#H>�m�u�	���F4]v�(���]K~��I՟L������)�sy2-m���)��ÿD�Ix�� 8�uW��>�2�^���x}B�u�����:��E����F-`�S���ܟPm5K��oZL~2�
�KĨA�Ӡx�ɟ����S&X��Z1BŘ[X��	`y2�'}��'���'�"U> 2
ڴN���k̆692��E��M;F![�<����?)H~�9t��w�0�+��`�M�b,��<��mc�2�n���S�'D�ta(�4�y�_3�T`��KT܅Cp#��yb�K�&ZQ��;6�'�i>��	`�`�x�d��6�X#
޴+٨�����Iß��'9�7-�-]����O��䑗Q���A�ml�ja�ԍo'�P��O�m���M��xb��M0N�"eѡ/��1i�Չ�y"�'eM��8kZ���O���?�?9���O(����
�o|�Q��R�e�l32h�O<�$�O���O��}���+t�}�@�2s8th�d]�� ��#�> r�'��6$�iލ�$� D�Ȁ[���L�P
e�r��P�4@ɛ�os���P0�vӺ�	�$�$�&Q��$�Pv��A�?46����R'��%� �����'���'�R�'� �+f�m���h���BX`�!]���ݴ(z����?i����'�?i4[=T���:��%7����-����ɹ�Ms%�'߉����O���X��pi1*ȣ5�ɹ���8:$���B�	��剳"��0V�'\b�&��'�"�pR����7�.����'qR�'������V���޴%O�;�bך��VJ�&�҅�`�Y$��3��7��v��[i}bCh�&��	��MS�F}���{!m��0�lEb��ɢ1l|�n�x~r�Y&�X��ӻ��O�+�d"��ցBa՛#�^�fL��Ot��O����O�� ���d<�7̒M"nY0�f�P�� ��	�M�`���|J��}��V�|���@��a:W�ǗK�����M��O�l��?�SO�v1l�b~ҋ�=@@0�"�ͽ~i�T�����'>d���蟌��|�U����ʟ���ޟHx��_�j�2,,��2��ɣ���ß`�	dyr�^��Џ�O,�$�O��'i۾�B�C�2��$�@ܯ#���'Ք�l'�&��OzO�3� 2��!Ĵn����\;5����㓊W��A�C/;�P��|�s$�O� O>��j��%�r��.۱S���R'g���?���?����?�|:,OԤoZ�$��*�Z|>�i�nݱn�D���HßD�I�&�#�R��>�u�ih�p�3ǜ"�ly��m��$m��O�7��>g�6'#?�SN�k���C������D�k~�b�[�m��$�<q��?���?I���?�,���*<+pb]�@f�_,�<P�Gɦ�s!�쟼�Iџ$?�����M�;4��8ɇ�̫\x�h	�lށ�N�Av�iYT7-�^�)��\���oZ�<qρ����҄�:5s^�l��<Q��X�/Nf��T��䓭�4�6���.B�li�#ض<��+1��8�~���O��D�O,�?����q��	�Z/�E:6�
�i"�Є��`��[��	
�M� �'G�' ��h�L�:F�*D�&#�$7:j���O�U���8M�ո-�I�?$�On�
[v��F�D
h��I��S>B���'���'�B�s�a�qB�y��8�h��D@ -<�ݴi�)s,OP�lZB�Ӽ�g֊*��TY��۱@L�庇�<�f�i��7��O��	�o�n�EL�᪶��T���/߼�i2N�� �bЁֆ����4��$�O$��O��$��fyi�����6?6%At^�vp�N�6��7;���'����'�R���U*B�
-�Ә9���>�v�i�<7M�O��F�t T�=w��X�K�{��E��9Q$�Ä*؉��$
&fr�D��w>�O����$R�S�9X��V(C=o�����?����?���|b)O�o�f����	1`J
�tŔ����0�R�a.批�M��b��<���M[�Tc�<af�]�X@ʭ�gJ�"�l�/��M�O��@�����w�X��eHBl`иJ�E�,�2�'���'��'���'%����n�����f�=.��x���O�D�OBplڌC���':V7$�$V�\�ED
� ��բ��k�|��<��i��7=�ȹy�`h�*�Zi\8��L�0�0�Ҫ� �JIh�!��(ɸ�$�1����4�0��O��
5*
}ɕB�("u���ǏÐ@�j�$�O�ʓǊ�?9��?�(�H|s���[7��R"r�ȤJb�����O��n��M��4����0S$�*zO�2t�Dh����e:D��z ��O[�i>)���'���$���Sl�}`��r�iʲ'TXP����㟰�	埰��ğb>��'�~6�_	o��q��۠n%���`��>(R�Ʃ<�ǳi��O���'o7�V"#��,q�)�;	���-�,�Gq������B~6-#?��ۦ1��	%���)`�t�3�K���r�*�y�\���џ����� ��ȟДO�� ���=H��Ē�o�7�
) �gӀ�)�O��$�O���$��睥=�h�̀<�Xa��m��� ���4?���'�)擰d��m�<��H�:����mA,'��s�kY�<��Cۯ��������4����_��ʇ,�X� � v��S6D�$�O����O��=��VIƹK��@I@$��@��3a͂�8E&�h��VU��C�����lZǟ�'�P��йv��5j�h޹�LS�O e�����+��Qf�G��?�f��O(�1�a�0,�t|��̢a`�B���O,�d�Oj�$�O��}���L!hA� U"iWܵ��AI=q:��I�^I2���$�ɦ��?�;4H��0�F�k�Vѩ���ʰ��O���pӴ��KY�7M&?�i�;y� �)�^ ���d�؄R��aw"�!K�p�M>i/O�I�O��D�O��d�O\A��a�9���V�U0_z�}�W�<�ҿiOƠ�3_�,��X��
�h�pl��4̸M���`�T���P�4��ߦ=��m~J~*A�;�^�9��\����07K�(�t]��ˆ_~2n�0s<���?��'r剅��R�!Y l�^�J!;��%����d�	���i>��'��6���{�(�D��){���	�{��Y��D]7!���ۦ%�?�V�\��4ܛV�'�\�jT�2
��薭 ]���RG�{�����`��#�V���9�p��lI�R��E#P�2D����3O��$�O����O��D�OP�?��'�Y!^�r4x`��hq����Iǟ� �4�x@-Oz%l�I�R?�1�F
 -�nmBG+��Icy�G}Ә(lz>1��LA����'OH� ��th3���:e^��KՎ�	��x��0s��'��i>��ퟔ�	�8�YOK�=*R䀠�U
���IڟЕ'�6�!7����OR���|���7I`,v�*����C�w~'�>���iV�7��O��~���!34P�����ą��N���l����;��������';��2�gۥ
"XH�T��M�'�Y�w��ZQLӋy
�}"'.�g���ئثш�ye�1^�>��TL�E��[��|Rn��|
���̅धB���O�J��HQLhpc�ҝ�J�KǄĸXBޤ)@ə/�A06!\��}k�gK��ĉ��ci�H`"��߲Ljn���̒Hn�q�

;h�&��g`D ?�:�����6}T�q(���1�^��,�E�ݳ���(� �#nW*+���)�I�!RC�9�GA���QCA��5l�� 4�O�@Y��:D�7Z$��ZC��>�*OJ��0���OH����^�>-��Z� ;d��W#8XÀ�3���O\��O�ʓg֬��W=��tKw�{ �S�@O�Zഅ�D�i����X&�\�����TCQg?�!M4vhT	��F�$sQB@n}��'�b�'剶3ذ�y���M�O<8�:R�S3�*��+��j�nZǟ�&��	ǟ�#l�d�S�? l	�m:�J��K��I��R�iF��'�剥SO��Ү�����O���O�y^�\�G
�9�Lm��٢G*Z\&���I�j�OCS����)�	!��[D��:�M��e�3�M3)OV��H�ܦ���ȟ����?���Ok��p�1�BL�^�pQ(������'��h�4�O|�>�ǉ	�(;���#H#i2r|ЍqӸ���������͟p�	�?y!�OfʓVLK�-yޤy!F�4\I�e�MS��Y�?&mYT~2�	�O�l��)JLv�E�F��lňQ����ϟ����	  ��Otʓ�?�'@�P`�蕍	^r��[�pm"'��̦��f*?	�/��w2�O���'�R�Ō�z�{ū:(��$Z�ꚯ/7V6M�O�}� ��^}"S�4��Iy�Լ�Ī�,�R$b���h*�Q���G}���,n�'���'wBY�4q�G���<4�J�"�$�s�.5�$X��O�ʓ�?�I>I��?	Fb�7S��a���>4�Q��e O��
M>q��?������ ���'+�0����w�*0H-�S�ao�@yB�'��'�R�'N���O$]�R�ǭ�l����߃ 98e��U�$��ԟ���Oy���3X�>�'�?�R)J�Nɚ�x���&,�"�+�`�	M:���'l�'���'�h���'��1®O�ˀn_�/n��!�9j���i.��'��	6f��[O|B�����@H7'
�L�LA��ӛ<�N8$���'��M���'|�O$���1%��BA����[�D�-Y$�6V���g]�M�DR?����?eK�O&!1d��	k`)�bN�ըE�տiG�ɩ(��5�����'�򩶟T�̍c�`q�gC�`�N��s�l,
g�̦Y�I����?!�I<�'gnRy�@&U�Xi����J�B �J��i��'1B�|ʟ�d�O��Y�I'��1B�]�ū���ܦ���\��

��K<�'�?a�'�Ƞ!!���z��2q�V8��P#۴�?�N>�GV?���iZ8�����VH�QC@(a �O�zc��<�*O����ȍ_����cF�.�Hd���3 ��<�����O�����$FF�	�aӀ;Ǆ|k��NBظ˓�?����'Ur�OJ��)�B�4��p�ƚ&�`��i��+�y��'��	ǟtBv�_h�UA�(Y8M�QG�5"��wn�Φ���⟌�?Y���P1$�&�A1�,�2���k������	���?�*O���B�N�'�?Q���Tc�`*F�Aq�1"6J�)s�����O��>��%��b-7LQ��W��fu��j����<���`XJE�.���d�O�����U�3G� �������-�h}@�x��'[�	!F5�#<��!q���d���!�h�j��Û'JH�l�]y�,��7��6m�O�T�'u�4�-?�/��b��X���S���d)�ɦ��'�B�':L�������=���򋛕k�IC���M�	^�ZR���'�B�'9��%*�4���a�$�/0ǀ82p��6)z�HEA���۟`�	o�)Γ�?��+
r������6P�����bś��'x�'襃��8�4���ĥ�,��OF���$��悰v@�ԛ�yӦ��4��s��'W2�'a�OƟ{q%C�'W  ,�a�@���7�O�iۖ �D}�[����|y���5f�і~��A���Ɠ�yؤ����DA�r�$�O��D�O&���O0ʓE�"5P�ă��H+�`O
5��p��d)I�Icyb�'A�	㟬��ݟ���*�5-<M���(�
��f��k �I����	����	ßP�'�x��@�e>���d��O�j��E��8s�51)bӌʓ�?!(O��$�O��d�^�ȼrd �p�ՒKc����1.B�}m�̟P����|�Iry�E31���?�1Ul&e列(
0���b��-pb�l�����'�'�"���yrP�00G���1�~d梇�US���O&�	��'[�����~B��?Y�'#cj�����U�� ���N�`0R����П����0"���'���S�6�4���*�!$2�1�nM%\��V���r���M{��?�����^��ݖJ�.�9�f�<R�Nh��J[9+�@7�O������:OP���yb��U	��T���>iN�8v��0����
OX6��O����O����K}r\���J��1۶�2L��*(!�d��;�M�b��<yK>)��T�'���ru�M�]��e;�Ȗ:�-��zӢ�D�O<�D�]�2P�'���ڟ(��z��p���>��N)^do����'t�j�����O��D�O�`�KS"&��DG�<Mpp!eF����ɈP���K�O���?I/O������e�����ȿv�L��d]��Rh���'5��'��^�@�Y?��p{���q"�M��d]_�,�*�.�I%� �	�8"�,V�l�ѢₜO�����%׭
���myR�'���'��	 )p}��O�,�ZPhX��y�e)K�`�ؑ�N<�����?�����(*��Z���勤K��k�]�i�^��[���	Οp�	oy��E'{�$�.xIU�QPg��AT!ġ`�9�weW榹�IQ���)D~��=! �
+`R��c%�f�΀0�)��)��ş �'�:I���#�i�O8��ExXA�Ċh�4��ϯ
k�D'�p�Iޟ �%fm��$� ��!|�H�ʈ5�����Л������'m�,�dv�@��OT��O�`�Z�H��Z�7%�$�oռp���lZԟP�ɳ*���s�IU�g�? �Ų��2�0�yF$N2W�r��5�i�xJV�s�����Ob�d�t&�����,�L����S� B��f���ݴ @���䓘�O@R  �?4���%�A0�6HYU�T%#�r6��O��D�O�vĎN����P��Y?� C��~���2�J'~�)$��ʦ]&�<��t���?����?����"?����1*�M�T�@τP&���'��]�4�0���O��D.��Ƭa�jL$p0�����q6Rt��Q� ˅�h���'^��'^��*6�  ��p�E��f'��q���%���}�'��'v�'a�� wX)�V-ٙTha���yW�\��韸�	\y�B��=Y����}�E%ЇZ���:DV�l6t듨?A�����?I��ZSZh���K�{3�N�zj<h8�Ǌt�$�A�[���Iџ�IZyҌ�������#�)o��𑳰
%o�$A�n�ןX$���ןP�D&l��O*P�ǁ1~��8WDۖOth�K�i�r�'���@O�]�H|����z�AB���u)r�X�\[5�w�R8/��	џ��I��h3��x� %�|�� հI+ ̀�G�~��ƒ,��nZvy�ǩ0\Z6-Z`�t�'��D�%?�5	��c8E�Q.�}���VE٦�I�4�6�]���'�@�}D,{0
݀c@[�*"4��Ԧ�0�*F	�M#��?�����v��8�HY��*ƞ�^u��j�>q��=m�)x:��?)����'𬉀eC�&]선�o��{�����i�����O��d��Y;�5�>���~�,�X��=Z��g��BL��M;N>�qE��<�Ok2�'�R,V�y��X�U*n�R�	�Z<7��O����Am��?N>��Lv��aC�
�-N�bP�S8:�i�'���c�'��ܟ�Iϟ`�'MVe;"��l�p�B�S�_�N�@��O%#:�b����J����	�=���3��H9IĂtc�	ӋO�9q�������'��'�r^�*������*Ԝ!�8Ɉ�H��Rs�/�5��d�Oأ=i��?�z�"�)C S�N�aH(@�a�\�c��p�P�iaR�''2�'��	� H+H|SH�#
� ����z���4B�f����`��H�ş��	Z?��e˛caj�3�E�/i|m9���ɦ��	����'����2�-���O0���$�%�D�Qr�hQ�g�<+.̒��$�O��sM�O�O��
z.����o<X��!���@d7��O����C�<���OH���OZ���<��O���D�T�_��0�T��-Kn�nZ�������""<����J�<���Re���$��<`2C |4xHj,7h�t�ѬB$������Od�+�Ɔ+�A)�U�i8�-W"O`X��"�GvN��ү�>,� �c�:w:��5;xI�zSt����5i��1���6Ś	p��&3&a߃�*��wD�2(3��ґ�\�#!.m!/Нp[�|#r��"����Sa�	�z��F�<4�}�[�7	~�H��Տw �8�p�hF.y�%�٢si^Z��uG@���O����O�8���?�����X�
(���f�1L��ѻ"��/\��s�G48�=��R�u����8�QJQk��^�+Q�dZ�I
F�4�R�u�t)��?E�*	���Z�M*�̚K�'��Y�lY�e��ɡ�ǃ���Lۻ�?����hOL���4
�xp�ph	�tK��Q7$ D�����2xe,t$5E��a3W�<�Ɋ���<Q3E�����p���TH��a���ڴ�_��ɀU���쟄�'0{��!V�T�*� M���߳�M���Bk�j��q��R��D��d�6"\Э��Ϋ~k�-�a�<�б'H-^����Ϟ�5�����'�bxa��?�+O�4�ІE�	�!���0��h2��$#|O��� �R�2t�Y3$�*
sDi��ORPn��Z��;�m�=H�Nh���J3<ư�I~yr'.5����?9-��؂���O���ɛ>H��+2�`��mKT��O^��(ǲ�q��S�T��i�C(�'�򩁹���`�E4������@OX1��+9�9����H�0��V�Ǯc�l���	\�0��}�>qG����j�O��"�tN���ED��Jz���(O��y"��]�$((�ݯA&6(�C$���0<)�鉥/:��I7�����6�س��A�޴�?���?����5Kؚ���?����y�;$-��q&n�bQ�u8�˅q���3�D��W�d�|AD*�aZR�g�;����(��lC�%��FT�R�T7[���	i�0���|r�� g��+V@-�#0<\d����"08��L>B�^@��"�A8$��	i�<	���P�@���ޭh�� ��e~n4�S�ORbY0���:�ֱi��Z�g��p���|o��c�'�2�'��xݩ�	�ϧY	ucC��/Z͆�K`�G���9� �, ��A��n�#4�^XHϓ)�x�He��*`�H�JΎ�\��T&��b�.3���2d�> R�a�.UR� %�US�b������������?9��tc� ��m U�1P��h'���y��Ř"�TT���t�@�S����'�x����F)l�l��4�ɾ&�u3�e�R����f�0eS�a�I�<�����$�	�|
$�ʟ�'�� 0A�"HS�}8��[([0(��';��،JO�~�l��ʃ45�E��e��p<�.��<$�t���4���C#���<ލ�6�8D���"��1���Q��"MU|�X��6�dcݴf�1��$�2&�d�C\�z��1�<1Ƥ��y�f�'�?U����O^tQ�$�5�8u�Fo���� ��O����&Y����.�|�',���3a�1>'|9wj��V�>�
J�$��h8�S�'l?T�8�([Bp+f)�{�ŤO���'�1O�>l���]�BD�2u`3(���"OJ0����N<�����`���A�'��"=�fD�g�D�z��23��T��� nǛF�',"�'��x8�-XR�R�'�>O��	�_�X�c��2A,<C�L�-
81O��"��'t)r��]Vl{��N4P�0YX�{����<!�-M5@La�a�21*�%S��;��'-�%s�S�g��?q�lbfl�	n��C7e�$��C�I ��S�(4Y��*�@:�#<?y��)§?�����W*]��mA�ō�x���,�-&������?����y��`���Od��!�5b��B.��/��'�� ԭ0�(W�\�-1R]�%��`�,�ƇN,e*C���/1�1d#S�.y�q�,��J�NI���O��$̮mj�C#�7�F-�R�5g�!� -1_ƈA��J�V� a�e�Zc�1O���>A�۸<���' ��O�2�5��׫M�^Ar�؃l�b?O~`�$�'��:�0�Ұ�'��'F��1 CH�jp�� P��Z*Ǔ*�H�?Q�����e�So��1��}X
�i8�����O��O*ESsL��dfl]¶Kں-()�g"O�u�`�kLι#�+I|(�OJ�nZ7KB�D"�`�
L��Q��Xc��b+�3�M���?y˟8�cu�'N�� ��Ҳ6�zKDᇴjQ�SD�'2I_�rp�T>��tH�V��͑�$�-�re�OH9�`�)�S�l0��2��.J���x��V�8�d�'�(�������O+dm��������RN�f�	�'n�H��I�9��@��IЬQ�ÓG���|�7��b�ܣq�ԅ�͒@eZ&�MK��?���sl��� �?����?阧�#G��8Lxd� ���Lv8�k`ژ�'1�Jϓ+nX�{����o��@��#�Cr8Y�=���xx�(3gG�#d*%B ?��H�#�z̓<���)�3�$J�ue �`�@�0d�����
�*9!�$'=xT��Jp� �3G�͔R��I��HO>�D�H�`��0�c���8`�.V��,VOΟ��ȟ����uG�'L"4��YSa����ޑjC�x�F�D l%!����4P�!w�K�ah�P�u.�	h�ܫ3O�!W���`d1��I
%Ȉ�7���'��'���'��O���W,ʥ��Tn�s�2�H�"OliJsHC?lX��l w�j�4��_}X�����M���?��c�iG�Mc��U+PDA��j���?�'���
��?��O t�BŊF�'6Y
1�|X�e"!#
6���![f�*Ԛ7�Ky8��K�K�[iF��1�Ї��L��d
�tJ��`E�tj���
��x��H(�?�J>�ň�Tm�A8ֈ��~K���LX�<��=ge4G�ń8�`�B�LOQ<qw�i�� a��7�Jqn��JwT�y�gގtqV6m�Ob�D.j��ğ��������!zU��&X��Y��ٟX�	&t�R\��X�S��O
l(PE�-(�f����ݎ=q���!�>3�������V>`r"~���
UBY�P�����/�o�D\4:r��ɑ+@L�kA��nw�}�= �!��kz��t��\ъQ��k�� ��=ͧM���tA	���	��.;*�>�ZwHؖ�M;��?Q�&�����?A��?ᚧ��pdA�)�ř��"7�$���#��'�֔��HW�#Ƥ�mc�e3@#_�L�=��&�vx�� ��,�F��g*X&.�x�å��I̓-�x��)�3�?�$`��9B���
�*E�%�!���_#�����PXf��v�-C�����HO>I��U�a0����+#�����PA��+v�ʟ�������u7�'��>��5�dI�
�>�q`���H�B��1�Ĉc.!������ �@���
<�@���E$[=.)+'�\��*ߊF�T���b�$bȉ�6��A���d0�O�U{��S9Kf���@��̬Q5"OH)(�gG5T��b�����C��d^z�2�x����i��'��dPäј�d�X!aU?�F���'\�ֱr�'��I�-�j�Zp�Y�Ɋ9bw�fӜ�P�#��s�8���VD��q�'�-�q`���~|`f(J%D�cؕp;l ��!���үZ��p<�A�ǟ�$�PZF8l�5YQn�?z�*D���G��������9J}C�)�l9�4'||���L�x�΁��Ń��U�<A�k�D�V�'b�?	�P��OD�ZУ$Dah�@��:ֶ�Z��O��D�Qa\�D+�|�'�"�;W��,�p@�1yX&�;M����:�S��`L��6@>N�T0��P9�2��O�	� �'
1O��r��u��-*�"��I��X��"O��#�*P�		����#>��(��'~"=aL��r�Yq��Y�v� ��)W0@�&�',b�'��aYD%�(Y.2�'����yg(
${���(�5{�������z��'�vP�EM׻C�џ�_(��']�+�qӣ8:C����"���3�#9�Ջ`�!�	.�E8�7O&��4뀇I�l�s0�X}Z ZG%�ش�?Y�C�?���,O��U�r�(��&ɯ&��4x�[=��!�O��%��0}�����Z(����t��Pkܴ|��v�'��6��O�˧��i���d����Y� y��WK���?�؄K�C�O����O��NȺs���?��O"К񊓟t��`m�U��x�cY>,��aH�	�:z�y�.Ek8�4�t�:3�@��5@��oP\�bC�B�!K�8lo�U��c�2B�x�LA�3��� �I<V:Ua���21�����b�F�k���p���$-	�9��<K�#ѱw��L����y���	;�n��(O j� �e���'N��Ә'�O^NH��L��Z�pB�W_����'��U��ʖk����ĕ�'dfL��'ȽJ�HKl���b�$!���'P�;�M�� ڜIUKNN��b�'����D�xς��T�MA�x��'��"&��S�ȝ��e��D�j���'̖�#�JZ����kvkR�5�@�'.v��sI��d�m�Ba�:@��8C�'��uj�b;��S��D����'\e�����
��iѨ�;��S�'�)q@/Z�K�6!�׈R4� 9�']l]��������f� %��<��'d�����üG�� 	E������3�';b���� 
)�)��^	����'��1:!)Z�x4�d�d�i�`�
�'� ����G��!�f�V���'�"��v��N���[��X�'�.�WLD��Q	
ARd����'#��eL�9����V�	9D��}�'�|M��NZ�\�Va ��܍>b	�'��`��F���$S�M'����'v��0�F�t�V�9n"j�t��'�P�Z!A@��=�W�Q:��Y��'�Ș��Ôn�h��M�5�"Y1�'�-Kc��(R�.X(�,�=&p�`
�'����{�p�'�J���	�'c082ՋԦk�J���cQ?�Q	�'�BD��Eʀ���
.b(��'vra8��A�$��ri�'���'������-C��a$�p�h98
�'L�;#����Ypf��vla��ռ7z�Oj�}�'ui�u��H��9�qL]54^zM�ȓd|p}�fE[�d��S��2E���ɵo^�E
�'<� ��S �����\;�	X	�_�l�5#�>	��I�8;��ED�1s��(2��Rn�<i�	��nE�����c��!oh��?(�mBU�2�'Gq��0# Ag?8
''ܚ�]��S�? �:�
cUN�	&F�P��$C��ͣW����=���O6��EΏ0$� �`o�wn���"Oƈ�d�Y�Z�	`�ǨA<�����O\�1w����>1ufUiJ���tbWHņ��7m@l��l�'�8u�s���o��!��lJD��'�X�t�4b
FX�t$�7jEnt�	�'���5�� #��JQ�@i��e@�'��ᇄO	 t�H`�dU<D��'w���A� �D�ˋ��2���'�6b��E >d�H*���.�v��'F8M��A׏(��d\��ht�	�'" 0�Ǚy��q�bo��[�rġ	�'�Hz���+O��8��@��X�<Y	�'���	�K'h��P�*��Z�ޅ(�'�v��4
M3)�V8�pė�N \��'�t�"���u��#�,9�y�'A�V�O�W
@Dk���)6>����'���x�J
!)��1�EH6i c�'i M���$_��H���^��\��'Di�U��b������1!j�m��'L�(adAHE�a)Tn��*|���'2� $F?Jׄ���B�f���'�� �e�&E�Q�E#�nX��'Fɢ��SU��H��I%��=�
�'d����%v�@`ÑD:s
�'�V �G&��GR܈z���(z���(
�'�20a���(PP�0ɳ��i{���	�'�b���H% 4�k�O�h�ʁ	�'1� �O� �����D�\����'�l4AkV
D�r%���X�Y$�A�
�'�� fh��t�~e�7.�$CX6AP
�'V���'m@�b���b��18G`ܠ	�'��Ij3@�����3�A�1�ĭ		�'@ě��Q��1�ƅȼ*�����''��PW/�3D2�MI�E��Ęi�'<�a����@��y���xmr=��'�  *Q)L9���u%��Gj� S�'�H1�p��p�$$�p�Y@���*�'ݺ9Jㆄ�r���
aDU	a�][�'�� �E�M�VZT��U�2�2	�'X��Qj�D�l��
A�IH&)�	�'ޤ<@����k�`H0��"@D�a�	�'���[i�8���W��9Z|��'�.X�q�H�zF,L��`�7DU�	�'9��A�ƍ!6ʥ��4[ �0��'Jb�r2�A�W���`ǃ[�R���'%R�9�nĩg4�a�IوB���'i���Pj�.p����Ǐ��}"�C�I�&�(�`���r�)��Ɣ�;	�8
`�br���矰۰>!��O"�a�ΉP��oQq�XR1�	9{x^d��$*��DV���`n� ����.�'"�!�$3m���vНP�ZTM��]�	�?�5���_�D#���ەo�"Ё���6?RFd"B'9\!�d^�z�0t,�;N�[��X�5��u ��B}���̺�����yb��J�$��7�OtҨh����x��N��m�AfԙS5H0�ag7r�c�,�lV�yՃ%�O��&�L?{�`���p���+��'n��k0B� ����>��+�;����3�E?�v�	�$_x�<	Q�� 	:UP3�S��P@1��t~"f�|?����bm)�#bs��T���S�!s
�q�'�Bp�<���}��`�Mߊ^z �����.Z����Q�Ԓ�H�
/fc>c�X�0kr�F0�qg��x���E9�x��kB�w����#bƍA�@��c��z)f�:g�(=*v�X�o�9�KQ4�H,���ּC�9���Z�z�I�b6��X�O� �̲wN�)�x5����+��EK0"O�q;Rd�#}�����$���`*@t~�ލ"� ���U�lԨ#��J�K%�xKŤM4pl��G�e�<y'2�2% ‗�#�@Z O�y 3 \�<a��� |Ҹc>c���Q �Y5�X�j�j����;����%@���B�Q�����A�^��` �>�:[�`���bc8 0�y�s���-��H��	���!�Q̚�?�dM��O�0����+zU��P
L�D��h"O\|Ӳ���X�lI�%I�E(>�s�"O�����9N��
�d�Ȁ"OyʴI�)Yp^��n�)R�9
3"O2T
�E�5��1�L��Y3�i�P��j�L��r\̙�B�8�0|�gF�#sR@����J~���,Eh�<IVhD�Dq0�`G��>t2Ĳ	]�E�K�']v��-��((:��O&M*A�3hP����Bɠbm.Y�u�'V�2��&��	۰���N��Ur ��c�>X0x�a�M�����(��y2r)�,�8��қ��'$�x@�ә�Mc)H/�������u�x]y���!bY��2�͆Qb��:@�D8f����rN$D��`�����횤�?2i�,������f�K�=ST��*�%�����H��(t�1AI%>��QD��߼ G��<\���.Ɂ
�BP��`h<1�k�������؞h�`����.6@�WハY��͈DޮA~���pk���ٯ;�"P��c��/d*�I42��FHJ�=��-����v"��DK�9���'<O�D#E�I=R�ѹE�ݒ�VT@���\\�"���?�^,jwa\7 ��]���Pr�.">a3$�a��d��g��^�\ ��aO`�Z�L �'a�<єR�=��p���]AX�D��/(*�[��
ZcT��d��;j��򆪂��a~"�]a
*�u��.2:0颇Y"��E�' :��ƨ�,�	p�M��JpB\����N̪�!V�i�`0TiC"F0h����C�̤ԡ��=� �{����	�Uφ(��̓5�7����Upl����9�0������	��<	�nE-O�^�JG7 ј���QPx��X�JF5$��ɺ:p"�:�I�!tL��@��:Kw�C#J�X�G˜�m�J��pO�d���9��dV�+< �K��,̴�X�a�$��'Ĥ�a�f~�)�(Y�h�� �)����s�-EW��cD@L'���C�f�$��Pp������dX��Ԕ����7Mn�s�k.k����'��)���8�)��q>���ٍ2�n-��wޱ�dƅ�p�up�ST���%9D�L[��G���f��m�$�#�k��Q���4h�?,�m��^D��6�����-Rz��'ɠ%3$	��H��@���x��'I�$1p�/`
� ��ګ>�����e�%]����*Bl���� �Y�q�?����LF�{�l�C%O�B|�u��	Y�����,
��O�C�"�A5�
/~�����x��!B9è��ɑH=��Bq�Ɇ3��(3��Lp4�OְSbK�B`h�9���N9�t����fi���ؽ�-��A0T��'y>����Oy����I�7Cb��p��S��?�c@�;
�y3 �^n�'�����T
�Ж	�XG��N2�!�Yo|
����M?5V��D��v��$�¯��.��dհ)�$(h�z����e�L9�p�c�ͯ2��h&��#,�S����|����!&Fe~d�`b.�K��ТF�{H<H�\?�5 �'�1o���@�ĞV�� ����'���<a�j�MK�Jg��*��x��hh<�eK��}��}[�#	/�! ��V�E��h��'@�C�D��Iז��U�	�&�jϓM߆���y���&�~�O3P:5���"�y"(*�X�� �_K�1��씩��[C�����doW�m��\:��$	��}Yu�	�y�ѓd�YC�#=V�-�lU�Z����'*�*dZDL���/ޠL��E�	�'�Fe`7.,{v$��Ȃ�,���$bUr�!���?&�d����*���hN��y���"1O"-� OK�)B�� !H�t(���"O�r�)�-���j��^�`��0�|2�_�h�Oq�,�&�0��]��L�
q�B�"O>���9�BbTkœtfF����͊U_0��DA'�h���)>\���!��Z&#��BF�
�,��eH�üEr�O�����3ye�����ɛ0�*I��"O� �2�$��E��4�w�+)���1"O�ɲ�g�>o�$3g�
��2�"OL]� e�bO�#��-h��L
�"OBI5ĽAZ�3!�Шa�&t�"O8�X� +&��t�0d�6w̜�I�"O���gYl�����ϜN����""O�ԡ��Τ!n�!�)O�!�"�6"O�i1+�	cp��E�K�kI�T)�"OlD+M�ll��gG6,r���"O����f�gR��^�8$B��V"O(��읮u+8�2BbX�r�"O�d[B(�-~�F�˶ �U�"!��"O���&�'k��y�a���:���w"OP���\�sen�����r�ʥhV"O�	��΄�"{��S�<:rF�c"OhURnx&P�*��xx��u"OL�de"&��6�W�/�����"O\���?�zL�#���kЀ�U"Or�����	r����+h�=`q"O�H��m��	&ݠ��J�$�� "O<(�Cţ\큡�ǸB9v�U"O6�A
��7�*m�Tj��Q)4�y�"Otha�}T꤀#(L�Pɀ"O$��P�^�+K�2�ȡ�FKZp�<�a��"6�����B)i^K7@�P�<Ydf Ti�D�!Q�	����J�<�t.�\<���(�\g���5OF~�<�"��S9��*����9fT��v�<��揟V�D!D�D�:���2#B�p�<���@<1��2E_8
�d��.j�<q���25�4�w�µO�vㆨ`�<y��1��	�2(�/9
����F�<����ic4�3�ǧV,Ա�Y�<����N�R�Q@Aj �z��p�<A��?h��"#!N�<���BB�o�<9b������sf�5u�J%��o�<A�d�-�T��"&.|�m�@#�i�<i�)��+	VM˰��9�ё�	�q�<���T�x���jN���`�l�<��
�-=�tur!��=(��A��<q��D\�0-���]�`I�s�<��Ɗ�.Gf���G�6+D��*
v�<�1��� �h�p�A�:ƾ!�"HMr�<���	(�u�rYl��(���X�<YG��-#�x���#�z���"�p�<�4�U�_,��8 ���8��Ee�<�s⇫c%ju!��@�ƸM���c�<aa��N�I��lX�W:>�`�Kb�<1�k�8ՐH��݆+��8yr�O_�<!b�3O��\�gNV��<���aC�<	rJ��	��i�g�
�xqJ�����f�<ɕ�_�H��R��T �i�<�%l��b��L2��D�&� pG-�i�<��Δ=M�@��K NbNa��"�h�<Y�Er��Do���1)c��e�<��6D�d�kE{o��U,h�<�2�Ҋ[?8p%��E� ����j�<i'���m}l��cOɊ%��5
n�<i�˝�7��\���TY��d�g�<Ym�$]P�d�7��2zD�#U���<���ʚi ���%��jK��B�hC�<����^��(@#kY�;Ĝ�ʢ��z�<����p{B�j6�����TM�|�<��`����S� �R�A�*B`�<�  �b�Mм?�>=q��;[C���b"O�Y�N��N���!�+<b� �"OP�Ч�Oz���C˃H}6A��"O�y�Jܖa���A��_��d"O��z�Ȗy�)��ڲ(�����"ON��#XwA��⑦��U��-�yR�ɖE�����`Dք��F���yR�
"jd呇.T�g��Lه�)�y�;��IÍ��b�3'��2�y%��1j�Y��Х]&��Q`��y����_���4��s#�=�����y���"1�a��ǔj{�Y��f�y�D�s���R@=cφ�jG���y�GP�-��5劈[6N\4���y�`�rOm3F�Wdl=�V���y2HF�-|-�׊��^��D�f�B�y�S6�����ݟC���a��y�� vۼ�P7n��9����e�̱�y��Q�z�K�E�(c}�d僗3�yrA����/D��ڬ)���yr(��^<� �Ѝ^�*�v�3�y�=hڐ=��˂��TP�l���yK�7�c������$j	,�y�@��^�^�7���`����e��y�*�S���S�F�i�b��㥑��y���7>�S�kקh�lL�-� �y��"�.�Igj��UF�}!g@��y���X���!3�ոD?d\r����y��a��`J��׏8K���R��y��61 rPk��@/�thZU
^�yB���F-2)����U�Y+"�I>�y�@V�yK��Zc�����yr�ߌZ0		S��;Tp��C^��y��� ��`z�Z�b�]�ф��ybc��&ݸ��D-#���Ѷ��y"I�>	:�P��L�� $����I��y��#
	�A���tf[Gf��y2�B>�D	6��HfԪ�'Ο�yr,.\H��"���("b��b�	���yҫA�F�d�W' �d0�(1��'�y"��v�Cg�WC��`�
��yb$: ���1��Lh��i��Ê�y��I�B��(ִ0~�#�I��yR,�;FX��e�Z�� �ũ"�y"GL�'�,h�!-�) ��"uK��yb��$8g�
hJ��#�'�y�c�Hf�����)1��c�?�y���8v
 ̉�.W''�6#҈[��yB��- ��bF_5vǼFq��j	�'J�r��I�L��
J7�|]��'|duK�+a*2�#�|�:tb�'~JySfEbˢ�8���p�=r�'m�h+qBΖU|�(80'ͱQkL%0�')�p�WFR�hyq�*J'J�u"�'B��pjׂp2�@
W 4\IA�'��)�2D�Iy��C�*���	�'��|r�H�#���`-��)^��	�'��͹t�0H Dk'/�+�$(�'9<���i���蘘�0��"O>q�q��#p���dg��y�͹5"O*h�F�?r<b1  <5��"O��፱]Hp�#e��0T2�"O��tjޗF��aqSD�i�|�`s"OP�FG�5hr�5�ѥ!Z���"O� ��j!'�`
"u���I��5"OָsƊ��_��L����5!X]kw"Oz�0t��\��<�'��W��a�"O�1)&�D\�����&l���"O��3SdȰ4�Z������"O��bfQ\2p�_��hME"O�M�)2����(�l Z�"OhnFOI��v������&�(D���7	Z�h���3�	F��yBd�'D�SW�@//��Q�ӡ�*1��T%'D�P�f COn1A�/���M�q��z�����d^
N.�q����D��8c�J�H�!�-���e��@z�8賩M�#!���'
�#��Fw�	�VZ�!�d�<29ny�Td��0��ZQGT�N�!�d�4yT�`1����ش���4/�!�ªt:��*�K��&����d�9$�!�I�*j��r�bC<%&�!ƈ��p�!�$L�m�苗&ߝx�P�gۛM!�d�E��)��� ���+L(!���wy$����ƚ�:(����6�'��F�iDqOq�RH���7d�y�.U6l`1b"Op��H�Ep|x��,�w��%����IܓQ��I���L��2����[u,�xSG�<?�����-D� ӷ�F���a����΀@��/}����p>�o�:l0\tsp�M:m�,�%�^U؞x�T�|r�_�OA�6m���A�*	��y��f� b0��e&	�ò��'fb�q���� PL�48`!S�Hr�P�3)�y��2�9	$GD�8�2����yL���@;� ތzK�i�R���y�ԃ���"N�	<Pa���yrɏ�j�\��G��$�p�劷�y���|�]P�W�(�8)J���y�D��s��[欖�n�8������'ў�Ԉ��W�kEB	sF߁f��!�F"O�#��]q�ԥA�DH�B�1�"Ox�A�fȨ#�p��7����5	��>D�DC B�Fd�A��-*rD� >D��4&�� �У�lp�C�;D�����ƓZ���R!�4jz&��B�'D�tѓ�K#k�=�%���2����!�$D��)`E�J��`;�FP�:b�!D�@p��O�`�n��$E*`5(	y�� ��xR�ҭk��A��J��Ïם�yҏ͛%FsQ�ߕ���%Y��y"�ցpQd��U{1l��B˴�y��J�1��'��6z��0�K� �y⦁)C�����,m�\�ڠ�ܟ�y�Q�n���h����ś�CB��y��
�lbt*r��<�|�x',F�O\���ߺ��t�0zph�'��!�$�9&�1�$�*�42�/Dy�!�$�'S:�D�qď0��Iv��G�!�HuW�}(����Y�P�C��V�!�ć\�`���a)� ��0R�!�ErR��b�̚0y�� $��(�!�Qi�0�M�C�2��W�O�i}!��7���1�摀+�T� A�G'L}!��b� H�AqUVŢ&��Q!�_��H`@g�z�n�6��
�!��p�jD[�( �T�Hq`v�^�G0!�^�m�0pӀ̀�wqLA�Ц�t!�$0\�H�$oP4'^�S��4 R!�� N� ��"��	�&֘<��!"OP�!@��$c`0�#f�a�tȢp"Oԅp��$9�$"�k�Z��`"O������x�n�Rg�-]�V���"O<�*W�_=j��xGNs+�[�"O\�0�E�7� g䏿Y�� �"O���H�'� u���7 e.-�%"O���3��O��yУ�&a��i�"Oz"�C�.zf���%�"O�5�S��K�Z�&A�t4�I4"OL�3�#��h�����cU;%����"O<H1-��@ԞC
���a	�"O��g ��q����n�����"O��[@郐7x°�@���~q(�"O&P+��F��(�J�G	fy�T"Ot�� -S����ޜ9���K�"O@�0�"-�<�rWL�	y�a�"O�ĳ�L<�*3k�E��Ԫ�"O�:���;���S�i�>�@�J�"Op�R�k��"D��"��#�ȼit"O�ܚWL��8�D��5@��U��}q�"OP@��`'2wv$�`�T/�Ta�"O�i��˘k>V�r���f*v(@ "O�\��"�!r�T��m̸M"�y�"O��@���7nk�5�6-�LB�S"Oz5`E]Z�{5�D�D����"O�j��O�8����,/j�Xp��"OZ����������<s�"OF�(ga]t�.��>*fʐd"O<|Z'm��e_.��&,�?c�K$"O4�ڡl�#_�e�W�TxJa3g"O�
f�Z+h��x8%���fq."�"O�Š�&9M���I3`�t�"OT\�O���������!"O�|��!��+2���"�zѪE"O�4�&R�z8�P�p���h�~���"O��A��%hvk'���f�8�
�"O:��D��9��<Aa"%Y+��Qa"O\�)�����Q��V΄��"O�Pe�4�|���l��yQ^݃@"Oj-[���9���i�[?Z�k�"O�!��H�VдG���v@��C"Ob���Er���)�^�-��ٙ�"O$M��R���Lڗ(�ҭA4"OP���HG�Q���P�Fo���"Oة�kĈj��=�4�˃��	�"O@�C`Η� �|�Ѫ����E"O���N)h�>]QFl�B"m�W"O.`� ��#c<�P´ ֙{	&�A�"O$���S%�����_/#�Ruy�"Oƨ!�Ȕ 7S(-ѓ]Ty��"O�9�ϗ�V�X� �m���P��%"Odp*�@I�p���Э�+}*YP�"OH��a�:?-\1Q��HQ���f"O��x��FGz����e���R"O0���ׯj6$�	����>!�L�"OJe�k:��(#��A��# "Oμ���JI���BL��Z��ԃ&"Oj4��۸Bt�3�	!C���"OZy!����~5�3�ٌm�r"O8�0�Y�-l(e�b�G3\r���"Oni� �?@*,��B��6g@r�"O@02���iup#�ѢWK0MS�"O�횔#��sr����I�5>4�"O� ڰ�@XT�0�aJ�i��87"O0�A���A��*D�-=���"O�-��mY�dU�8´/Փy�(�+�"O���%Ė]�X����,a�* 9S"OZ�@Bn�1��l@���UBX�S0"O�Y�  Q�fw��p��U4��"O0�
�Ð�uT�P0�,ƍN#|5p"OvUk���
	_�t�aˉ:g\H*�"OLX�p�����q��1j��1"On���@�|%r�it\ ZP��e"O⤙�MK��A���Z�0C��"OB���H#S��Q�c�}%=�q"O�T[��>�
d
�M���X�"O�ГQ�
iox	�� a��5�s"O����'.���z�j�7�pL�g"O�0�$�C�KFZ �� ��b"O�%᫔�7�.\z0K�r�x�Z�"O�Y��D�*�����o,����"O@Q�5�B7�T�O m��@v"O�q1��	x���Z@hďg ��"O�%u�2Dᩤ�����܁�"OPHQ'��	?`�t�wFJ�2h�lBr"O���$�ȭ<��r�R�F�DӶ"O��(D�X&U,�Q񆝌)6R}��"O0ma��D���ah��}.���"O�鹁��K��ӡ�5d��P"O�l9p���IA4�34���u��K�"On�SƋ�k����T$6�$Q��"O��p-��/�l����# ��<:�"O4�8���,XZn�(�\�Y3"OZ):�H,�ƭ�-�[��aAd"O� ����H�i��i�8��"O�� BF4?$�����l<� "O*���F���A3'��=i��ӳ"Or�iWdE�S\���TeE*J��+�"O0�1�㛋���X����b�L|3 "O�蚱���su����߲R�z��@"O�PVM�;2�l5!F�C,_��A�"ON Q��.}��2 ��R�� �"O��Q	�n������w�0`"O��&��:&�ӷBS)N�l �"O� cE���Dl�!��N�%��"O��7G �r)�e����ne"�	"OЌa�����r�
7`�:@"O�{�̃g����L�$2AC"O��ᡔ�6��A���lH��"OdT2�b�
##�A����$7�%Q�"O�8P�E7 �@�D!��,�ؘ��"O&�q� ПOư2�I��3�"O6D&�t����'H�=����"O��Yvۂ`��D3����~�V��#"Oؠ U&_�Y9�颰*�
�~���"O��0��*�P9�c�цz��rG"OH$�S�1?�ڔ�'B.N�T"O��8�ܘe�n9�Da�P���8�"O���Qb<yH�9��"ў����"O�Ɂ�I,9�UA ��3!5 ���"O �J'���e'�|zU��;l��˂"O�wn@>QL�q�pA��g����"O~H�%��!(���u`���T35"OޜkB�̀���:��P���ա!��Y2Vd
Pe-y�T�Y�"�c�!���D�J�c�A�J�6��S��+?�!�d�i�2���h�W���w G�"u!�� n|c�)Ä,K��гgL��"Oޱb6��	Z�x̹7'@.@��{`"Op�
��ͦ}-FI��ߊ�#"OL���{J�H��4h��0ڥ"O ���!=�:� �����2d"ON�!E�� ����4��&0��<��"O�!R�C�>٪l��H�l��  %"OV1C�ꅯT��� h8kB��A"O�@���RJMJWFA!(N(�+�"O,q"6	Ҍ<�	uE^�m?�d��"O��zB���*)v9��s�`�"O(�sK�p�"�Gi�/��,u"O��ض&΁J��Q3�-£\�$"OV�:�)t
p`׋� �@8E"O�ps�f�9
fHx�)��{O��"O8!q���88��p�Ё�.)�"O�!BԪ�*A�E�T�b�b�hf"O��5F�)vER#3	�,O�d�"OL@&�4gX܂�MЧQ�zL`�"O<� �枇0F�"�nO�C��۷"O<�:��C�[۞P0-ʼ$+�ŀ�"O<�؃&�)(�baa�,�$	��d�t"O�u@���j�8,U-��v��u[ "O�9�bBA�v�#���@�����"O�0kD�5?W.�d$˨9���"O�Ś�+V(\yP�H��*���yr &%2ܭ����:9�f=j�lL0�yr&ފV&��!m�,2zP,��+^�y�F��%�����#<,	K2n��yO�.\gRP#�V?;����6��5�y���.�2@���1. �X��y2H�`��ң"4*Q�Ř ͪ�y"i�nq����^�K4@Y��ڴ�y�g��u���Pc+[1I ����d�=�y"	=f��I�⣄2F���(N��y��@��ruS��W� F��"ħ��y�`Oɨ�Sw�~I�xp Y��y��#�
ĨTŀ1x�ؑ"���y��W'�}r�΁k�:K1����yB� �`��1��\�f/��W�ħ�y"ˆk�<�j7��d�p	٧o�*�y���0=b@
ŎZ0Z�X��A��y"�#p�1QRhQ�d��2W�T���xB&�29DՈT��\`j$�W�+kr!�aGh�+����s�j$�Zu!�Ě6�J���"�7<D��K��F�!�$� q����k�	 ThZ�`X�!�ɤ}Jٴ	G0)� ڧM�<�!�dL�x�Q��$�10 rx�DbX�-�!�N(~P����10:�IP ^�Bu!����
�Aveޒ^������v�'a|�ˌKu,�ӡg�:.��Ff�.�y�+�"F��lxd��52�,��j�yb��Z���6��2�
#���y�2t1�B�"l���ɢHЅ�y�C��AZ�a�W���Z���\��y�k�9A	�]�e��P0�*���yB%	z�9S _�
5��!V��y����yhZ!�A�����ȍ�y"�]"D���i�7rY�� ��y�)�����)ED3z�H!c	ط�y�
����/�� b���IP��y���$:�t��X�"��<A�F��䓑0>C��F�jy�ԡ�a� �Ȱ�=T�� ��B@5��xK����^#����"O���dj��Eh�=�e�# �91�"O&庀�C�f�xA�QJ��%��T"O����O��F�iY1JG1�L�V"O\Ո����̱A�h	+$��ӓ"O� vd��8\�hH�/�����'.�'����>��"�?�|=�ݚ�rQ*�#y�	A���OP����ИP:`���	5u�T,��'P�+u'�e@�� ��gh�'d�y;0E �?��y/�����'c���A�=>���Ūjyr�'�$$���\9i�$�*:v���' zM��e�Q;�E`$i	�b�'�L��T�ȗ#�҉�S�µ��M>9������O
�L�E�=zB�<@R��}!�8�	�'�j����::p�1���sʐ	�'E���CE�iv���.��d��d��'R*(�1�9��e�'@V11Мx2�'P��[�NΒ2A�4�	@�*��]��'�ZM���X/�$x�H%���	�'ܽ�ao�$[���M���08����O���>�B�Bũ\�`�� �&p�2����3D� ����	�~�P��1lQ���b&D�8���4i���F�p���A$D�ȩ��Տ�0t���N]��G� D��[$�&%�r��6�M���4D����I��.A��V<N<�P�1D���b'
+�~�:a#ׯVt���2D���3`��f* ��t�Ҫ"��3�+;D���A�S	U��IF��6J��@��5D���+�<����a�ݜH���H`H D��s���Y%���B`�y�$,ِ�>D�DSfA�N/�y3E� V<���%0D�@+f�@J��k"DèQ)9*C@:D��㡭��!32�0ӫ�%Cep�O�O|�d:�)�:�|l葤���"���D�>�"���'�u�A �Y��8��Y72�9R�'����#H�+@��Q �w���'!��á��<����'B�g|r���'�8���
켄���o�H��'�|���6���/��j���xߓʘ'(�P3�`�6�)��Kƴa�(I����?q�����"�����PSii�/�? �C�o�BE���^�� �)�!�D@�v���C� Ҹ������]�!�� v��d��'GcɌ�{�ʃ6�!�$�N�.��!f�*TW`�Isk�7D�!�DL����z�GG�j8�)Kªܔy�{2�'��	������	��NnT�i�L�\����O`���O�˓��D%�I:A&�e�t��5,u���!3-�B�	;U�`)��D�W�.11���l�B�I�f��'�>b~��:d�L	C��C�I�������:u�j�QŜ�b4bB�IP°tEV;D�0�`ږ��B�IDnLQl�� �&��_�
��D�<Y�'�|��#�s�[e�ZF�KK>����)X�^��u�`#��k��p���I�!�D���Ԝ9�&�&��ҷ�ʘ�!��<Y�Y�%�R�:Z$g*[�!�d	l疱�	���Y��ɝ.+7!�D��度H�"��`����R:!�Z&-h��1�X%m� �	�G�>d�ў���S�)6$s�g=�F�37��S��B�	'j����*C1C&A[�⊊y.�B�)� z�b劘4�h�h� �NRr,*B"O�����$�2ag��@;f	�'"O�k��%Co�q5f�_.�Is�"O��˧ޒ&l���Z)Lp�6"OaY���,2ҵr`��d��jB�.�S���xH�P@��?ڔB�Zf�!�DW�8U7ώ�p�� �!�[-3u5ɐ
�8
A�Ġ�9-!�wӬ�e���:�A��g�!��q�}�W���.��0$N�E�!�D��I��!�IȨ4���#�+�!�� ,�ej���:M������
Zўȅ�ӛTb �f�Ŭqz���V���Oj�O �}��@2l�rؙbU�b�*P!xɇȓA��!��%^_|�y1_�j�쭇� ,^�sGAϑ@i���$�ڕD�<�ȓzI���"o�>X�"mH�<D�ȓF-}����)J��UKr�QpNq�ȓ1�p-��ʭT�޵�� iB�ȓ����A+��B(.p��W�^����	hyB�|ʟ0b�0��bݹ@�&�)%1K��e���7D��@EŧU��h��hA�u=��e�+D�<G 
���HBO�*� ��2%*D�d@bY�5"��+W��8��E5D�D�����5��G�+I�6T8��4D��Z�BA��T	�A�P/ZL00A'�OD�	W�.����4nY`��74|r�O�����.�-�V �8������'9*�IX��(�0��v� ��6��3���X�|i#���2LOB�[��'ra��x��{�˘�y�!��<N3�d�a(�p�	H�!�$׼X�xؓ3�^�P�*�h�"s�!�d��YΒLI�,I�s�:���E ġ��%SH�O�7�(5BcҚw��T��	��2��O��X�<0TH��C�I�s�xXa�"��J��B磒z��C�	�m��$xnԻ`�n���� \LC�	���!J�DǙ-jV�����C䉪t���	��]^|  ��6�$B�I�?�E+jN�M]F�@D����C�ɥq�Vm��Ė�q��%���Y�t���7^D��U΀3 ��ÒA]�'�BB�I�f�l���H���	�"ɩ9��C�	1c���)t�:Y�p� L��C�ɓsKD�� �nt^!��3ϚC�ɳD9~ �'ȗ�Q�p*D�;w�rC�;�P��P�*�.�P-޲�l�1�S�O�F�S�R�X��a����f�¥!2"OZ��2)�,T����B�jX:�"O:����$;!�L2�'
�l�� ��"Ov��6�	�G��(�$�crh�3F"O飦��2,���%^5�Iq"O�<�v���>�8�Sbԙ �@u��"O�B���r�ś���te�Q�	Q>!
M4e�]� �N�h����q�<�����4]��KY!y0ei��@�=2��"OLp�a.=6P�����&� �&"Ole�]�4G�R���R!D,ч"O�lp%�H-(�t�H4e

J��"O�ܑg��-.�D�B:i�(��"OP����x��A$�>�J 2�"O�h���3v���V�4,�}J��|r�'�
�'J`��vb�0h�����ˮ""�����xL���^���`�a��+W����S�? ���Ǎ:���#@A�l}^I�"OjH�g��#a�xP�%(Q�-�XT�4"O(��w�8��1[��	nU�i�"O����D�!Ih�HH֠O��т"O���C��&~#�4ɡ/�nE����"O�bi�1Mq�ђeD�n�D "O D�T��>���D��0*a"O��{���^2,8q,O.~��I�"O���'�B�o�.4�"��4*�|QB"OHX	�k�8W �X�!�ޒ��ٻ�"O���4ˊ�sw����W�h�2p"O�Y�ao�w��VI(��.I�
B�=M����g���F1����(d4&C�	�_�F���"
8�8}��M�6f{C䉱��|�D�N(�L��1g�1��B�I,��ꉢJ&�B�e[�J�B�8��+�O��l�6���N�5�"C�0�����V�tS�G��l�C�Ʉ�d��0�K�R��W��]�B�I
`Ä@1gł�c�ҥ��hM�B��3U\:A�"�R� ��͇r�B�	23_z5aК�!���ƩM�B�	�>7��t �u2�-Q���F�$C�I�N���P!IҾK^����c$j�C䉮\H~,K�-T�_��A�)o�B�	�F�f��dE�j��h�rG]�w��C�	�R
�E�0��6�@Z�j�#��C��oMМ�@�S^�8�J�U��C�ɓm7��b�۴[ .1��	����C�		{]F��A�(�&�:���"qЀB�ɒ$ē��@ ܰ��G�F]�\B�I4?CFl�&E� �v��DkF'(�B��}hx�3�ڋ<'j����ś3��C�	�I6|h��8x6T8e�'b�BB�	�ELj�;��׊w�\��
�DW0B�	�}<�0t,��1K�i��`A9Hy�C�Ir"f%�`�Y�j����@x��C�,N�L�!��.Wӎ��e��B�Ɏ�����F���%kW�83C�	�k ����e���;�хn��B䉙,|l-�1G�?��ś�ЮIm.C䉲DU,��g�ۙ}��,�*��B��B�	av@��Έ��J��F�q�|B䉆q���*ƬÀz�.�����Q�C�:P����A��
���
'��^�C�	�Q�������
�eF��'HC�)$��	�W$�6?��樀�<C�I�t5�"w����"��D�!9�>C���|�GE]�+�Y#ĥ�2!VC�I0�\H��G�r��Dr�^#S��B�� [k6�AIY��H��ۗGݸB�$Z�^p!D��2@���3��]5��	�'��"���>�H�!��A�W3�D	�'4��b҈��:H���դ�� ��p�'Z�US���&0��R�*S�Kn���'d(%H�-K�bwR4�+C�Ɣ�Y�')�@r�[ =$B���*� �H��'� a)�R?��i�G@�,1���'y���鞽;U8E1���S����'ײyX����h4ps͎�Y&�c��$2�	or�7C%XL�9qS�ƫRt&�����<AD�)r�8R�ތt+�)��"M|�<a�/�<(��pC M�z���l
yy��'0Y�ы[4F
؍i���[�-���� P���M�>�e��2(�`%�#"O�aI�#S�-=��$��!T��P�U"O0�j�kJ[(4���gy�8�"Ob��,��\ٔJ�1l~��p@"O<)�צ
�N9�)��C�xq��_�H����4 ��������i�e�����O���0=�Ǭ=� 1cZ�X܈�b�M�<A�'�b4u�6���P1A"�E�<��%�8v�� G��d�L��jx�<)�%�f%����(w\��E�Kv�<1�&Z�p�����a't���@�Pzh<�v��}(Q��@[�X+��Xv�=�?�)O6����4ʘ� �F�wcp\V���'3a|rR�[n��������/��y�#��B��]9�OA� �1p#�y2%�� /��2�	�nx�y��d�7�y�k�+c��ҦǼc"���Ō��y�	GI��a�W�N�\P֣4�yJk���@Ϧ5�뢇_,���2�Oft� �H5�I��ENt9�!�!"O�R�f�yA� �dc�$b,;T"OdI�B��_��l bT�(Ʃ�&"O��@܊[ɸ���@�3U�b�3�"O�RB��:E�q�#��X�6q�"O`,3&�,8_J$�Ə�AЬ@q�"O*(P���.-> Tk�ώ,q�\TR���|�Im�ďI9~[<]�B��G�����+W�y�'�3��\����DiȀ�+�yY�THtA�"Kb�Ũd���y�o�W��ɚ4�Y/S�޸y��Z�y���
gH��e���L�0 Q�U0�yr�^/:;�)�Al0V�H��̶�y�K��`�P�x=$�|��ФI���'Fў���<ɠO�;*H�@ɝ�%���wJ�D�<9�%T�P�����5u����UA�<�F�˕x���ŨԆE+��c��|�<!��59��T���?��A�b&�r�<y7 ����C��}��PZq�	d���OO*�0T�O�M$�	��Ϳ\/B5S
�'V@8kU�^�L����R]�a�I>A���?a����O��P�Y0x��������*!D���"�<{[�ઁ#����:D��QU��-%��|:c$��F"�B�,D��3oDI���C�	j��њ�)D�TI4$ҹ0������̱1\Խ���%D�DĂ˳@�[��+�X�˧!#D�軀@�-%L���%�	>|�L��<9��hO1���Z��ªRɨ�c<��e<D�p��I]��0���˰= 	��;D�{ ��;�$�e�J'L��AP�'6D�|�"b�Ls� b�H
7gܢ]b��0D��CM݁V��h�d�/j~y�v�/D�$
� 2Ei1"D�r��5iԌ.���O>㟄�<�w�\5>����JŇ$�RQZ!��D�<A���D�QņT�MÒ�і�~�<��#�����mS5G��a	a�^x�<e��/iҥ���JN"݊c$w�<iQ�Cp���'x�>��r �<Iã�=oi�0������hk�П<���n���Q@�E�r�y�D�z�̄ȓ4�=*�A�,k��!%@.xX�ȓ�(���0]5rgE�%K\����x�1��Gܗ���⦐�Q��ȓ�]!�F]������̦|_ą�S�? (h�%�N�B'Bu�q�ՊZ��("�O�������`���y�1yw+D�X��ي2'��0E䋨~��`�I'D�xq�F^<GT� R�l�S���I%�&����T�AT��0s�0(2Wm�6if�2"O�`����kDD�d�8)���*�"Or�{ӄّD����V�J���R"O�\��nº<��y�ARCP�D"O���a��CB�( %d���'�!��	_���AI8,��Lȴ
�/\!�S:�	��ǌ�c`(ʥPџ�$�$�O�p�тG�|^����K�K3��	�'v�I�,\ 8��4+W�+z�	�'��-��Ί�4(���F��'`��'q��z���_-D��W"�(�'��x�D%��D�b�+t��,O����4� ��0�P�N����@0��<�	�<���ÉdbL�`&i�7���%�H{��^y��'5�O:�9��1�gKZ+L "��K#"J0�"O�x��)� i��	r�p:@"OJ|Rh8��Z ,��\�Vų�"O�񥞵I˦�10ꆗe��5P�"Or
b��V��(2ъ�ͪ!D���3��`����M7:�e�f�=D���&�]�I���D+�'&��3��<D�� "K�|4�`��9�Z8�)'�D*���'�[ÅY�@�X�	��6�c	�'RPD����c�f���Oɫ2[bXk�'H�p�T��	�c���+�Q��'_I D��"#���B���v���'�����AN ۬���㑬Q�	��'%�C�� F��C�-ޤ�
��'��i�҂�<=�����]4�[���)�4aI����|͂p��M����ȓ6��9B0�L=K������;����4�P�%�;��DҲ�Q�|ڂ���:tb,q�+WB z��ΘJ1������0�p�آ7�*,zA�U�<���H<�Ac�9�.��pɀ��x�[�l�i�<�W��%^r:��3�d��`C��hO�'�R%��:a��BpmQ4l���ȓj�ryӊP ^��J!�N�Oޤ�ȓcd�*���n��8���Uv(��#���(��Ԍ5���RU+��ȓCT�� BW�V=|�(� _Z.�H�ȓUʰ� d-
�8����M L!���F�8�@�]�MY�Oͳ2��0�?a��0|�򨗑|.ƀA�I0 ��Fx�<iqՆqRUȷ�M�t0�EZ�<Y�ۤ}J�s��{bB� 5�]�<��N=/-r0B��΄\s&Xc��\�<їHF)2�6db�&قJ?�4`l�m�<y0bD8ZD��'琪9/.�8V�A�<�U�H�0r�*� �T3�0��<��BC6��0*F�]�;`(�ð��P�<�J�5+��Sb�'��l��V�<!2`�:V��Y�hU	M����JS�<�D��0x�@������T���1��c�<�p� W�D%z��6 4}�$����T=�=+m�*p�|�@�&����7[ʭ�7��>&t�C
�rnŇ�%E\hC@/v���d}䔇�Q\d%P�����};���i��,�ȓ`�L�f�!R��I�byvm��S�? �=R����S�X<�^0��P����h��k�#$��
o�;@8��g�;D����P�c׬]K�a��T҆\(�,'D�<�.�*;}�E3G*�@���"#D���G�^.C j-���V����"D��*��K`��q��B@*���.D��h�� ��5��Ĝa�H C�+D�db�b�;[B8õ��DVe���<I���1A��ܨwI�ж\�_�&�Ԑ��o<���[�#jtX�e&+�,t	֥�o�<�F�E>ex��I��:���(5�Dm�<�ሿڈ8�FF�ul��D�JM�<16�@,�(Ыǉ�ܡXT�V_�<yg۵$4���F!�x�dm��C	A�<���ɸu:>\���QI��E�{x�(�'6Z�rb��h�2�;�aW� �J���'� Ph'��
4,�؃��t1�U��'Qh��Q[	-�
\����t����'���p``��jTC�(�f��'.(�rG�H��8�a�����:�'���Y�OǊT�D��(<5�3�'�v,#DMG{!)��vF�c�'V	�� �$	NE��oP�{{����'�0 F���*H����	ok��I�'�X�` T��vH(�'�`L�k�'Z6e��,{��L�M� Q�(p��'d�ibE)ׂK��6
�-N��@�'!��1"�h��MeI�E+��	�'Ì�7��
 �B�)�(�=�� �'*}z�n��}��ف�쌇 ���
�'�p�����5��/�#B����'VH�9P�ۓTs|��H����5Qϓ�O�����ŤuL���b�G�@YZ�P�"Ov�c&��]B�i�P�E�(T�"Oh)��3-���ZP��PH��+�"OiphB�m*i��\44��S"O��z�[�I@e�g�9Q�>0�A"O޴3v*��US���D^� ��\�"O�,�ш,X���%2���"O�d��[$$!����+ڀKij�"Op���*��),�",�F��!��e�
����]�<��bL�~!�ęf�F���
K�����Cq!�׋E�B�P���5 i�(���k7!���4[Ek�F	:Ă�1n��h/!��1A¨1&�PP�X��+�)4$!�DAS� �kek��`L��s��U�@!�$Vˤ�� �7��A"��B4!�Ę f�,ZՀU)K��d:�Eݕj%!��&� P9'ٮ[�����I��R�'���'@�)����O�n�����m_�1����5N̜{!��?"X�KR.��p0I-bq!�D	�;9L�Q�m�	t��e�ӻ|g!�$�$���-�*	R�Ұ�N�i�!�D��6�<��W!�43��y�F��b�!�$�5P��m���)��U�!�d&H�8b�N��U��ֺ�B�'v�|ʟqO�c��&�4��
�66��"O�r�ڛK��)���A3f%X�"O6i�ƈQ�kٚ�@�jA�u����D"O�-#2B��s�zE��j�P����0"O����M%E6L�p4cڱU���cT"O�a{2�%+��ܳC�:8���;R"OX�$M��Z�@��&���kи����O\��;��3� Px��jċN�	�ƭ5���j��d�O����P-���RQf[�##����  !���'&Gt� ��N�g�N�I࡙91Q!���n��k�UQҀ�!F�.=!򄔖_��� &΀�4x�)B Ɓp%!�D#y���J�c��g"�5;R�@xw!�dK#��ܹ���1���F��-�!�$�1�r��� :��4i���}��'�ў�>���j��O�fa�A�D�ze�v�7D��A�`nHD�g,I<xRI�2J)D�$`�F�(N]�"�̉Q����9D�衴mZ�f�KB$�m?��۴�6D����V�en�b�)4�b��v,4D�`Zrm�@&\!A�F���Rf2D�h�Q�t���Q�6o<���(.D�P+Wi�%T��*���|�Y&�.D����$*N\�b��=P��c /��9�S�'����L�B���d�BJ�-�ȓzeBEɊ�-A��M��L���c�*P �e��[��C�<��y�ȓz��u�����4~�GF!Rq����3fI���(�*�z"!+3�'� F{��d		����M\�W�L�p�a��y�@ȗk�y���:�z|�6�V��yB�4�
���1>��i�&n�-�y�h���߶4�v�c�'
�yR,ݸf��;��+B\�LBl� �yB�I@����,m��٣��yC�'�zY�v�}U>��d�۷��d<�S�O<6x��!3�����W=5t��
�'+�%YU�W��I�Nҕ%����'@D��1'�1�X��KȚNz,1�'4\��a�ШW�IS�UNd�E��'��x���	4�<Sr/�	u2��'�\�BG�1"��!n�YW���
��-���L
���B��ZQ�(#
�'f���K�/u�m�>h��q��'�(-cA��P���`ӀL&3+"��'�PM�Vg�.v��Z��L�;-��
�'��E+�'�0XBڔ[%*81���	�'T)r�K���'�/e��|�	�'�1u��-y��\hb�W��}Y��hO1�J�O�JY���y��(���&J�P��'�&@��"�O#u �,P+�<��ȓP�@U��G�1s��P��)^�����Ųs�ܿ,���0�>
��ȓu�))�$�<�h`��%1��ȓ|��B�
O�Mw(������>��ȓ?�hsj�����Q�-�2c���ן��?ͧ�O����΄�5�2��&I�����"O"@:C�5]��� k�.�'"OL���n�j5�L="� �2"Ob�8�
�2B�
3鄲Au����"O�PցT�c�L)sp'^�v��"O�	���M N����&F[H�t"OH��_�H��x�R���*U��Q�PF{ʟ��'^2%�ujF�[�F�NF.cj�$��.H: @�_~T���$5����#�I���b��u�&n�
3h؇ȓ!�l1s�[��)�@M�5Kj9�ȓ>���A��/r�(�%
2HGP|��1�q+W�3ͮ��o�YQ�}�ȓs3���F#J<O@U��*Ѵff��	k�����	6;\���+M^��a`��]|��B�)� �4�uH��%����`�u�b�����\F��ŧP��a�#�ư%���у�y�f%x6�i�Pjшڌ���`���y2��+a�\+R��e��;aJ���y哻<o��H���[��qkw���yBGB*g�TDr@�ø N��/Ǌ�y����/��P�AC�lBl"���y�,�1#�H�y棖"��`wF7��O��D�O`b>�ദ͔C)��+��+����"c:D��ce��%%�
��A\�!�~-1Ɓ"D�t���awh���]�:۾���3D�H�G㞝=5�� a$Q�<jƁ� &D��X���ӥ��';xZ}c��jXRx� Fx�k��I.������/=��R����y"�D)
t`�C �/�x��S��y�d״?p���,<�k�)���yr$�O;	�g� �fQ�N��y�ǺV��ɻ�0c_��f�@!�yҏ������(�A8DA��yr�_�w�ZԳEN=����D���䓗hOnc���T�Â� X��D8v>N����&D���3��Ti��8��	&��sc0D�ĘT'�o���u���P���2D� B!��.je��Bu��2����L-D� J�\�^�Αpa)W�I �R*,D�D#�س5�\l�Ħӌ�� Tg)D�p��c�1�l��CD��O��  ��2D�Р��_3M@p��Hb�P�k�g1D� p�j��!����҂�!E�<	�q�0D��H�f�
D�Y����ʲ�/D��xk_�XQb�3�y���.D��{AbƂD&��0�%����L-D�����Lh��D�0 ��&"��yD� D�p�BON�=���D��<:?T�`�o><O�#<)��6 �s���&H`|#�GPr�<�a��Z��	6�Ј�d�"��i�<A!ں7��mi�hW�Fm��GO^�<� �ܡG�h���f��qA$F~�<����p�e�X�H"�Ls�<!G�L
[=<l1u�R�H�ʼQ���c�<���M�8�ш�B��q���_�<���׍H�1&'H�[�Q�^p�<I�hK<&NP
rY�#��@A�h�<�㌖D&�P�󥁐c�`=ɴ.e�<���&����d��,�� �g�<� ۵"[���P�?(��R��[g�<A(y��:��I�@��*
�_�<�2Bb�bPۓLܑ/�L�Z!��]�<1b/�4�A�(��h�y���U�<7*�%���:F�_'o^�uKh�<��!������`�<� �D�c�<1t��X�^@ےdO�N�Aʄ��`�<�&��9nb��ee�(
u�@���Qx�<���Q�JS� ��!8�Z�ˉs�<�hD�2��G��(V�1���k�<�𬑰d���@b�((�g�i�<�; NI5���7b��T�i�<�ƨ_�����N�.�\�@sIEb�<����cNt�BC(-4��9�(Dx�<q1�. g�$2K�p�9a��i�<���
{�QGŗ��%i���c�<)� �;ˀ���\�A��x�A��D�<aw�ôx
��ȿ:"tI���j�<��C��D��C�/�2+���I���i�<� �A�T�����y��A �ih,��"O���eF��D��A���҂M|	��"O����o��EJ� ���ݺ1IV1pc"O��3��\4f*��1�ޢ^9,�P"O�	8�,�W$���4�@1��2�"O�ب��YЄqF�6*�k"OС)E M��x(�҅R<=%��	�"OB�h�O��F���bЄ7
����"O��P��3�:8ڇa�;um�%"O��B�ӌ)���JژS�Ȭ�C"Oz<�`S?�v��$�:g����"O�3�uZ��Ԉ� |�ܜJ�"O>�+�mU?B~1�!�
;S�� `"Oz��"9�੢�Y9"�.aQ"O�	CW4;z$+E<�2�$"O�K`i�PVP��i ����"OT�-T,Πhp���ck��"O�ę'�ة}�`��'֪&BR�"�"O�MH�%�#0`N��'��U4��"�"O�=��e�0b6��s0��Pn|k�"O\�3�H�,p��1���|���b"O� 	p�9!�U�A��n�1�#"O��q��:�`}�BH
G�Hm[�"O���r퐠|���%�C��r�T"O"�u+�.�J�����p(i"O�0"�h�@*e 7_��T�6"O��
P�}V�,Ke/L�9.�Р"O4$�eŧ0�CrMR*���"OF��1E�'Jv��Elڒ+�ځ��"O�q� ��� ��B�Ѣ"O:�&��3l����-�D�t��"OjIۗ�F2�ZYy��
r����"Ob@r-\���ѻ&C�3\o�`�"O�h7�Z�]�J�-��rr �"O�f�Y.2�,���z^� `!"O֬(�>n1�a����^:�X�#"O�ݘ!Q+�tx"�̠SV�:U"O��C@
��=����ba[3'��mZ�"O�A+fm�U���H5�	�-j6A��"Op�&aɝ0d4���4.�U�r"O�Ű�%غ>�".O�I��u(�"O���w��/�6 �Q�9w�
 ��*O`��3�W)@�0S��X�PZ:��
�'Tb)a� N�Fd0Y�HX)���
�'UJQз�ц�~�i�D�T�z��
�'�Y�0H1=S�i��+�K��L�
�'攴*#��r���('�N���
�'�9 �\.���W�Mn\XT�
�'�&�5�M� 8�) E�a�D�
�')^����\�I�@%Q$dL6R*~1�	�'P�ͲwU�����#.�;	�'#2��e�9.x�(�9���	�'�F�0�`K�M;F�ѱ!�n߮�X�'����B�5GuTb��O$gт�Z�' IcZ�#���dc�-9�'�"����T�D�6��(��c�i�'Y��z3 [�b��ŉt(E&��9	�'�hK48��AX�b ,(�ʨ��'���r����X�Ė&GZ���'+85HqdK�/�lJ��|4, �'��aQ"F�AshO�Y�T ��'i�5(�T(M5&�����h��	�'} H�#k��6cdXt�H�^
�q�'e� ��N(�F�ۃ$V
�!���� >i�`�\�l����#t�D"O�,R�N�Y�*%AEߺ""�HE"O�|Q� 5L"Ա0d��;Ȁ��"O윛1�/K$h��O]d����"Oz �tE����Pt΂-M��c�"Oq� ��W��A�t�Xw��aC"O�]9��u��B��3b"Hi�"O63 ]�2�Y�Q��<�~�
'"O6"��%gƼUp�C��je|0�E"O�Iۃ`�6��1�#>\y�� �"O��!p'S<
�����D��T)`"O�Y�Ch��~A["aҹ$���P3"O���Z>^r��!�4�|p�"Od�h��U�w5��r��}�+ع�y��\)]q��b�fԉ.:�A��U��ybL�73��,��Q��E�c�U#�y2�X�%�<��s蕂N�B�	�O0�yR�Ʃ9�I����Kx�q�+��yr���>M�du�A�@����`�A�y����E�5p�B_��d	ޢ�y��S�<�<�:���'1�И�ϙ�y��+P�.��$n��{,���Ğ�y�I"z�	���F����ND,�y�$Dv�Zg[F��i�tK̪�y��-�j1��W8>L��{As�<�G�l20��qi��3�D��k�<�5dL"� �RAڞ:��� �a�<�ć۝k���fi�����_�<�`눦6��r��_�~N�H#D��Y��71�lZf(Ӌ$�����4D����Q�s�d��?C9B���*O�QJwc �!�c� G;(�D� �"O���d�@��I3�̾{p1K�"O�I�a�0
>��sfG�(n:�"O&�� 晈;6��I�KL� n��C"OPѳ���<iiFYe�ϮvX�"O���C
�B\��)�i�~KR���"O��V.�4�&�[3�L+A�T*c"O`Up6��A!�\2��.F5�Zt"O2%`�cP)[d�4�G���C��t��"O��2�fڃh�r�2���"O�QKr�  \$tI�Yvp��"O��k�K�?�m���ށN��G"OFa��j�����K\	 b� �"O����n�;4�<q�D�[��Y�"O����,%F���h("���"O��mK�y��;�H�mP� �"O:�)u��A��]h��KY>��#"OLQpV�zF b�c�Y'����"O��ZĆN9g<ti�)�>���"O�!%@�d|��tǗ%p�F�jp"O��ӓ
S>�Ĩ{���OI0� �"OH	@2דW�(X�����$�D�"O�*���qf�����;$�JT"O��C͆4�z����B(
�P�v"O� ���F�jR�''޿5����"O|ȋ�i׹<��&,E.3���9�*O B7D��%x ��v>>l��'�,+��
�\�,1q�m��={�B�	�"έXU��7DP���FaİY�B�	-S�4���|al� ��5��B�Id2V�ӡ�"�D�jvME�)�B�I#8>^d��_3g����#N�ND�C�ɢ*�|�Xu����L���!�lB�)� ���Ў\��FT1�J�Kv���u"Ol5z�G�]8 �Ӣ�	z|�!P"O��J]#!��:��4d�`ˠ"O�]h�ȡw\, �C
�(XBd%�"O\���CK�o�Ƶ��#X�� I�3"Ox�s �ĒR��(ҁ�7�2��e"O�����<���Y'_�Ntl��""O�P�C/	�<��H�Q:jD��3A"O�) �hCP���)pU�4�f"OP��1e�F:��C�<B��K�"Oݠ1�Ȓy�^�J�h�� ��b"O���g� ,�\��նSB���"O��҅�͗(�"�I�&�a�b�c"O�@�c)����A��)$�uP"O*��!ω��Б�`�t8,q+D"O�HrB���4�*pz�U�M�)�"Op\q��(������%7@la�"OTu�#��<WH��A�&�C�"O�H�P��,"I(=�&�Gnm` �5\O<c��� F\ΔDH��)ls#t�����-M�Y8�h�'<E�=a�" �n ��	��ē)�tT�X7�L����22��+�"Oz����Xj��ʂ���D%*1�%"O�k©w���3$�����i�"O���Ř�(�s@_�n�PH�"O&a�Ƣʄ(��� R"�>I$)w"O��I�$[?&2�����.=J`�!]�L���{�dIy�,�;+$���$?@�B�IxI�D�$ܳ�B1r�n2��B��0�`Yz�K�P
ŚW΄;'���e����'p���>(��Y
�h�����'� a����-�,�sx�xCA�	T��y����"7'�2Y����I
�yb���\l5-�1�<�R�M�y���4^��``UVL�@��D�O��=�Omh1��ށ	�B��┑t�՘	�'(�0�OE6J�|!3��o���'�8j�J�Z��`�ҋ/m��	�'	�ݳn���r�g\.g�H��'��<bF��;;�yB,�����
�'�~hz��M9)����tL�<k���4�6�<E��4��X�q���ap��w�^6�b���V��Ṳ��tw�ɩ� 	�,�� �'w�~����'�ġP�D�*�� �ti1�yd��LlT�W��%3��S#m��yrf�%�P��O�
���ɓ�y��d'O2И�Ӣ5 ��c(�YHhY�U"O�삄J =\��jw��8��"O4!��폝'�t���?q)U"O��:�	� %�$MX�E��7"�p��"O�bq��Jh�-��O"b�1��8lOvIf$�1ی��R��0_�>�:�"Oq�7l]�r����(ԓ�l��"O�+ql�8b5��\�	k�lST"O�0X���� �ah�@�&n�Pg�$)�S�S�H��$�'�Y�u�L���d��-w�B��%7=D�ic$��|`VѩǢ̤V�$�<�˓;���aI�!k�����O�X~��mZr�����ɾJe�̻׉��L_t�M�*T!�B�I�i��'��:o�N9Q��'R������&�S�/&7��Y��M�t� &��c�^�?����đS��%.�0U��HdAS=U�OȢ=���+��F�F���9�,��;��:�P�@G{��Ʉ�n�}���\���੗)W�!!�� *�is�C 2v�a�C����H��"O&ݡ��1j��u����Q,����"O���'ݘ!㢝!��ĳ&~�0�"O��ą��&19��P�ep�ِ�'QqO��b7�#*{�I5�����I�� F��-~�<쓶�?2�̴Q`+Ă�y�˄�}Bh�; ��U�E(nN0�y�DM���}*��TS�B��m�:��d/�>ɕ(ȉ#PdH v�w�t��!Rmx���'6�Q#$m�5'x���ȗ|��
�'�n�9�̏���g�S<�-`�'���bN0N��V$���
AÓ�hO�Y��I?ߔ����L�N��P��"O�8%��	f!j�x�)Zm�J�t"OHI��� bJ��b.�,�x=�w�<)��3^z�<�jI�>�h�d�@X���O���6���*�O���0"�O���V0^�. �&���RDKe����x��I+G�R$�ǃ��rf��Pօ�
f�����?ړ3�"| d��X�*\��O�W�D8�O��=��Q�Y��Se]�wL���im�<@ѕ<�&��/2za��)XQ�<4i[���Ț����X�J֢�P�<�ǆ0&�<X6��9��%όF�<�4%֫_�
�Xm��\5�YK�Ɨf�<��Áx�:�$�خk�d�@�DDg�<	G��r��غ�o�d���h$C�d�<��MP�u�r	�e�"0��KS�Md�<E������9i[�|@�U!H�i�<�e$3d�pu���Y?܌�l�_��p=��l�"P,RW-��@�����P"m|!��-2ަ��@M�\f*M�7*ڿf>!�$�4��!!d�YO
��'G�u�ax��ɩRW$tIv�)/\�P�0Vc��E{J|Z�N]7
U�Q��Lt����g�<ɥ��q�!�����l�z�&a�<�g傆(�ĘB�Ol�p�S~��a8�X�0�����1��_F9xfl5D�)���J����!)�L�]�&D��C2*,F4��f�� �,"�M%D��s@�?��ئ��\���)��!D���B�Ȅ`�>���<����� ?D���A&��F��`3a[�L�D�(7-1�$=�O8e)v
�Y�T��I�A��@�b"OL(⧏D�t���i!Ņ�oG�rE"OͨG M�T�uX�L5���"O��Iӳ$f�Re��aD��"O���$��5�]���SF�ⓞ�����)�'P@|+��[,Xz��"�H�n�$`�IQ<��Z�J�{�v�Oq̓�yR��˽�����N���qP�ոj5����߰?QK�o������B�jQ����'�ў�'g,8lZSC��h���EA	Â	��z�r1�f(_ɀ��0�C� �]��aB2�b�_?t-Ճ^� (����Nܓ�2�s�	 <4�"�R�H54��ȓ,C�8�C]2p��!� M�wh� �>������Ĺ%���%���v1�e�T4�y2, �u0Z��e��2pt��'�Z��y"NM�b�)��n�c[�RP���yRo�!πAC�BQ�\2�=���۬��z���O�X�;�a\90צH1��?v�PA wI.�S��y��OR�(��o��o࠱� Pp�<��	]�^�̐;�Ȑ��oZ2�y
� @��Я�`7d��2�E�]��`�"Of
�
�v]��i��?�"���"O�t$��?�D��"�]�2p�t"O���EJT���e�B�<���"O�� �h��N�����/_2-�"O�i���,�N�@K�8�X3�"OJ�(�(��Ea�t�G͇8��B�"OV�P��E�a�H�`D�R��D@4�'B�$MYM��
���P
T=��GQ��	C}��� ܮ8�*	(k܅)d�
�"��#?����9�bq9Bh��z�n�JP矋D�!�DW�a�j���B|m��X���Ik��(��᳴�}�`i�7a�N�T<ɴ"O٫���$5`�̢7K�e&q�V�$4|O���qIS�z8�$M��1J�ٻ�O�\jf�֥����Ι+�\y�V+�q�<���	W��]�0��?I���@CBw�<1�HĘ=�µCY;4��d����q�<郩�2nO�q�G�m�:�C7̖Q�<�snHb!�G�F�I�f�L�<Q% 4<����%�\8e�^�p�f�]�� �<��B�#�l����� aωZ�<�
*q��5��D):}&��S�<�c �.O�B��i��;�Az���S�<)&���v���c&C�Y�V��M�<��d l��C��W�_k��j`q�<)d�FA��ɰ`�:,�"B �j�<�`iR�Y#b�[���q\z���Bg�<Qd�N�t��U�l��B���|�<��E�843vE8&HS�dx,(�@�|�<�#,\m��M�
=k�
Sb�<��͊6��Lx7�L���z���s�<���ܓ����h�6k�P�eK�e�<�W.V�0" /]�ءRTa�<�Ũ�:@$���,�$py��F_�<�,�%-�@�c�%ӥgth���_�<)"N����X�~�]�%�@c�<ɱ	�^ �h:G��,�������a�<�`o�{֤x4��e�a��_�<�&'�t~�u@`�sJ|�� ]�<i�ٕrv(���0O������V�<	q�J�4�����FF|�����[�<Qɯf�ze���Ϣ}��!OO^�<Q&�ӎ"�٨�Ϟ� 6�y��[�<qc5x���E w��E&WV�<���4&�AAԧ�Rf��$.�I�<���G�.fV���'�sB��Y� JC�<�B���J��	�F?\�03���@�<�V�Y*w-�q0�f�^)z]��IF�<��@*n# <q�%I9c�.����@�<!a�V7Bbl�t��7\{r��PGD~�<�����ؔD^�c�Ґ��"�r�<���.Y�Z@�$�A��h��Y�<�'A��v��t�R�������E~�<���Y#)���'��[�6d�ՀB`���� C.s������A�A��$U�/y�tEo�vD|,�%c0D��pTm
�%�!O 	�U�L;D�`!q��L��=��n�l���Շ4D���7M@�!㢼qc�7d��H�p�5D�h 3F�+\�%�Pʗ&@��t��a1D�(Y�nK�@�\���KI��m�6�,D��Y�A0F�B�G*`��m�b�!D��� .�]_�x�GG:R�����!D�����j�Z��@�ŦMg�M���"D�� <�%Ă&9��@S��PR�,T"Ol�'�ɂK_�p���f�X��"O@��f�.i�-u���t�[�"Ou�'��1zB7��>7-5ch<D�p�d�Z���P��F)x���4� D�X�w`ZJ�6�{��P�eh!���?D���I]�2Gb����<P�"g�?D��h�ň�G*��k��H�<)���=D�LrV
�;�j��3J�-~�8Y� �,D�h�6��G��x��ɉ
�5�tC+D��J�;�D i��ҿ7��H���,D������ �l��A�ʔ�DN-D�����E�@!�{���`9D�`�!��f���K(1KxT��4D� �7A>z�dx��:`:���*0D���ׁ���qr��@�PP�E��1D�`�L�
��d�/R�C�`�@#D�|aE�T6[U��y�cѨR�FoH_�<!�N�-�R�8�K��6�ȉ��_�<�p���	U�t�TMԩkI�qh�b�<�c��2lݾ-�E̓�os.i�b!FX�<AEڸC(b<R�٪]��ђ��O�<I�
@�b��\�%ګ%E$��E�<�%�ٯ����WbZ�r���KR`�h�<�	[n�<x�e��lT�i�0� k�<����I�fA�5��G�p��b�<Y'�J
Y|���RA���A�\�<!E쟒K���7R9�N�j��C[�<y�n�%Hm0@�Ζh�T��g�Q�<����SJ��p �N�n���*L�<aŇ;M���Vf��L~�u!�L�e�<����t���U�J�DMPSa�]�<�u�����'�J��z1��[|�<����I�De��0x���Bn�P�<���[�	�f�t�W�5b��S�<Q���7QVh3���$.�H,2ap�<��ƪ
K`�r�N'4�F�$�l�<�q�\>O7����TV�Ԭa6�Ak�<�ЅՎ
f ��̢lv΄�QO�f�<a� +>�P��L�X��H2�T�<y&�=8��rO/tA@�W�<�r�#Z[\ոf����-�UI[L�<���=t������;Р��L�q�<�v.C���Bd+Ĕo����g�F�<����1O���)J�Q2�A��F�<1�^��miA�R�r��q�`h�t�<��ˎ�F(��.��A@�����~�<)GBZp����=�^=���u�<c�
_E�ń�tХ;�%D�<�φ8wV������  �>����F�<�Ŭ˨J}��R����"i�ت }�<���&M����gE����b%�z�<𯈆D��rl��Z��*礝r�<�׎^#1cFT��K:;a��za+�i�<�CN���Bd�� Wm5��f�<��H�V��cA
ʊ{6�4l��<���U#	φ�@�(��i-d",z�<��H�:I�=��	4�pxA0!J}�<��k��CZ1#ӏ�dp^�#�$Xx�<���$wɰ���I�1e~�\�b��s�<ِ%ҁ$�R�b�造h�l�$-�@�<��I^�2U�܃�a��K�6ɂ��B�<��ˑ(�Jrf��lS�0��Ww�<Q���L��i!(H.F+8�3!�y����Q
O�H �T>O� ,		�/�|�����D<4[���"O��x����Z0�%�a�ϑV3J�2#�O�T6@�s���E��}z�E3�I(�%�;#ԡ�#�Q�<�2�ξt.��{૜�Jh ) ec�5-���s�b[���d����?�'R�1jdM�6j]Ju07�\�y�p9�'�"���ȕG)�y���MC���F�B�JĔt94%�2D��	(S�Q �>d���bZ�;d���Dſu|��q�[�=n�$�eO�WtI e���n=�ĨţgC:C�	�k�`�uÆ�z�f����
��Ob���L ������A7[3h|�偠.��3���'f4�Lpg�Y�<��錸zZ0�W+۴'��ƍ�?�ڸ{a��2{��Y�`"Q+h����O��A�O��9U��=Kk��1BOLT��L,x��q$��8a�� ��*S�ƠY���B�*�CV��ٰ<�#)�{�����:WK��U(ax��A Y�TL��%h":�F\	C��?3�b��T��eC����1�':T;�㊗[�*�s�Ȋ\z�њ�y��^���@÷U0�P���"��~ b��ܫq�~���C޺;0B�W�V�����,EA.%�rCګH�P`�*��f��2�#�?��!�gy"�U:���qw�L>E��aY3%�)�y�� z(��iB�a����"/�4��V�
}��"
��ٰ<1e�D�#J 0s��H�;��"��Cx��r/�P@�Au$I�6촥���K-���"��V?UF����B��D�E��w��̣���),�}�(��J�p����O��x�2@P�m���J�)J$Q�(%�˓[�>%)��3�dת��r⩃25pj�c�H�I���N����{��	E G��q̓�6a"��6���dw�'n�lHэ�C�S�R6��5M��:�1h�HI�}�t��'ptK�L��i��y"�!��X`�]�{�ҤF�O�rFqO��G�x�6�K
�rEn�9���9�h���A i�VI�f�Zh�B�	�:i�]��ʊ�L��h�b^��5^���<�u�^��<� �$�S�zǰ���"E!7�|��֬��R*z��Ai����ٻ���Ho�}�iB�}��	�u+��m�Z `���C�x���O?�Y��^0F�q�g��0`���gb�Y~�X!`ò5j�O�2I��G����9�����ǕdZ�@jV���D��?�p��G�2 Gay�/�$褐#f�h��QC-��2���Aq�Ί�?���N7�ȼK~n4i��)ǆ^30+�E8�Iٙo�Y(��hE�vL��c�~��؅a��(2��ܔ������ǣI0��4� ��U���)��O�S-���ˌ}T��S��-��"ж��)G IU@ �&����O����ƁM1i�☙4b�����q �o�����h� hl��ȱхW�.Hjp�� ��)�����eB�-�t]A���r⬐����>y�kJ�%޴C�������=ڧ34��r����`��Ƞ�C^o:%���h)C%ć���|���j�0�q��,'<{��D�Kޡ��t�H��P�ñk\��<���'+ܤp�	�4�li���լ^dar�G��9eC�v�����Z:S��<�����������a����L^�@�!�j\�<u�	N��8��	� ��S��Q-�΄Ӥ'̺)���K�,(ҨO���	L:Hqژ�h۾a����+qݑ:���	K)�J�(ɘ|z����)�r����-&��ҧ���a�D�GiպO���g�:�~2���Ť� )s�!0�Pa2|��IV�-���DK�@u�=�r��([�I$[�z�㬙U��8�CA��#e"��Z`��B��y1 `(�N�1R%
͓��N*�T�O����+�P1��4c�lk1�2V�\=��B�#?��܄�ɫ'3�e�#��/T�3Rl
�X�%�t�*{ر�0�D9&̶8�% R؞|��϶9��D��Ń�U��C@�%��x�#6S*�)���<qXt�Xwh��r��&�*@+��5c�h��'��"���"x�&I� aHf|�ҫO�s'�J�Kp�V�U� �[w��]�p�	ٮ5�\����k
�l����	�a}2�ö$)��o�=���)n���zSn�O� ����"�ژ�vH��5�Ju�t1��$��äi!�&sL"��P*V7x������Ybѱ�����u�h�j0)^	�f���^�)��Eak���``L&�O����f͏Ln���a�+��пi�Ԁ�!)qܓ|l��Ф��;[|��������7�MA+���k!��8	�!�D�%d�����
v紁�1�)Y�	�]t@���܌k�@���Rr?�����[���{�H6'�U3F�25������fm,8�U�'�����S�dW�S˃Yg�Y�\Np�J��Uf^5����ݪ9��`M���懬�, F{"(A6k?�  ��5dW�?�Ą��@�	@\�q(�_Bt1���m(�E;� c�d�@#�@�9mʥ�ȓ;���n�=�H �b���͇ȓ}�i�2`_"lP%Sǋ�"��a�ȓC��h ��IWR�qm����E�aR�ܢ/rm+$e��ni�c�d3d
r�S�'O�dx�2
�9'刵��'3b����J�J���[$4��fb�2'tԄ��{�Y�9mHc?O�KcZԩ��9�T1�DO��Bb%̡e����H��Wy.�3g�!]� �	�����E�D\� ���2P�^��	0��T9��|�Tz��	i�(�<q����/۱�yB+֑at:���۾Y�:�f����|��YhW�"�)�Ӥ)��48���x�,�ԯ�=M�L�>�b����H�Z9P6IvC�2�\v��;��5�	�9��A��L<)j�%K��Z�,��>��=;���<�4AZ-Fʖ㞢}���ìb�.L��؏a��x�r)J
?y6�:�'����F�.R��t�`�/�����O(q������=1A*L"lD@Ae+&��X
6 <�O$C�.LPa,�z���t]�a�� =��`S"Oȁ�"��$=;���
��A�T�Q�ɹ3[2����S�8���㖫D0Q�&�S4 $��B�	&>��I�:8}� ^`p��&D�k���Ӫu�tDb��wo�0���VB䉂H�ԔyDM@p!�T��)�%e�'�D����'>��A�΁�V��]�/��9�'U�LK�ح�P �!ȣF ��'W"��"*�<���Z)DR�'$|��F-Y4|���J� ,B��
�'M���iE 8UL��)�-����
�']�n�|@�pF���.���A
�'�@Uĕ��0\8E�@�	�'���f�
 Yֵ�'j��`̈́	�	�'�(���HѢ8��E��ɘ6gˊ��	�'�V��A��/m��}`@��+X���'�~aV(O�#���T�"&tL{
�'�R	�a��&x6��P�T�Od,�@	�'c�azcW�$ڌc$?g���'�%�bnZ2Q���!��УF%���'pl���&KDi����Z�M��-��'\��% �F�j����,1`j���'���h�ꅀM6���@�A21
�'�*���I\�zP��x`����'hh�	Ѷ&q��fO5m$��'Z��L���T7��~p���'g8���Z�k��H�N�I=|PK�'���q�VNi�� �\�K/���'!Y�˲XFI�u�+���0�'���2�g4<�����7R�����'���K���X�9��Vx��	�';�S�O��!��$��E��D�p��'\����%�HQAD�:iĽ��'4^�*�f�%��`�d@=��c�'�h�2fʓ<s@8ԃ&`B�*zb�0�'|�xx�m[�`�Fe&$@�}�
�'�J,"4	��T������zH�	�'�L�"�,&A�M��>��`	�'� y���S9,x�J �S*|�n�#	�'�4Y�.ۂ/[CG
� �jݸ�'��=�_�@��ܓՌ[)�T���'#b �1�L�����(}�X�+�'U���"��b�AH!H%p�ɻ	�'�J��C.��	�ZB̕7���'�u�d�(qR����
�?�jL���� P4Y���z� ��*�4�c"OX���Q|�@�q�gOF\�"O����'(4�P��
Dn���"O��Q��k' <蝥x(˖"O���0h�;A�rQcPjS�f"�q"Oh�M 0��4;qIü�f��"O�U!�FA�����x�(���"O�;�E������p�P<Ye"O�i.E1��"`��i��(�W)��yb(V�"�Q�p%��eG�P��*�y�#F>]O|�X$��k��daY�y"��o*�q�����q�	$�y�G�:����H\8�jЁF)���y���9S���@ @D��yˉ9=��Hj�A�u���h�� 
�yb,G}m�|����m�y+�j���y�DQ 	�:�+� ���@�2+�?�yR���+��9)e�Ɋ*�Ѳ��8�y���L@��$��_�������y"�� N>x,&�81�� �y� �R����&h*��r%�6�ybM��a�z�	�,���
�M�0�y���001��j �ɩ�Ht��^!�y�)�.L��7n���qvY�z!��� ��&hI�Dr1@���ڵ"OD �uDJ��n�rF��D9TX�"OfIA��G�n����@�9]B�5h�"Odi �%�_f�5���6I 9ht"O���S�	V�`���[9���"O�`�����l�z=���;4jjM��"O�D�q�� ����'�Q:���"O4���FصM{��V��Z
<�"O,�abHKs���`#fA3^D�9"O4����|
§�?}T�|:!"OX5붍��*� S��φ1��	�"O��a'L�V�8��wb�
#
��T"O��0�ٲj�����U�_ê�y""O��y����/����"��g���"O��.�in� ����2CNԣb"O��Ґ��c�H�Je(G� ��"O.�8���! ���*�g߀2�"лa"O���1��9{��i�R��jsL�x"O0�)Ba�w�l�X�+;hL��"O�В'��=w
A���!N�q"O|�yB U�Q�µ���ОJ�=�0"O(�{�ѓ�乢� K�0:�� �"O8Ȫ�.�01��ba@]�u=� R"O�4�۪,K�l ��Q�8<)�"O@���=xTD�R��W:,�h�"On�z��<h\^�iꁧ_�`�"O�� ��)2�@��>	�$kD"O�q����?_�����G�BZ!	"O��rU	,��@y6ӳw���Q�"O�}��b�+o<��oè>���	�"O4�z�BO�-L��ò��1(U*m��"O`%���%k&�fI	2�l���"O�HJ���l4�2aȃ��bIzR"O�TC��0yQ�z�
��-�t#�"Od��r�ћ~xd�G��*d� Y�$"Oָ*`'��vY@�E�m�
��"O�x d�\)��$�"����2"O��Y��AE���n�B��5h�"On���a�Q~z��5f�Z��<�q"OX�
 |*B�B��[�(�nq"O� 
�����a_Z�I'
I:O����"O�I'��Q�D(�tlF�{����"O�D8�j�*��
_ �qR�"OJ0�R*ܶr��H9���&	�J= v�'S
<��	��S��Γo� L 5�ز ��U���O����ȓ;�
���_�4/�ݢG����<�gٕ􆕒)@.�h��U�P	S�=G�aaI�,���"OTp
B�I�y� ��&�2��¨Ŧ#c�(��Ar?q��ė����	�(�"� � �?��s�)�5Y��B�ɄR�Z����w���k�n�T$q	���/e�h�)w�Y�4�a{�d�$g"p���`���B�ʋ��<a�c��f��<ʂK	 N2@ )ԪB�L��,2��Yq됷�yb"�A�~e��� y���S����!|�̻�#��)� )DIW� ]��ș��+��\���(`V�mӣ"O
ذuFG�48�@YV�D�(�6.�^kld�Cϕv4d1I�+��j��� *�xEI��84�U����S���Ɠ���4o>1�D�rD��:kʽ�u\E���C�
�(B~^���<,Oғo�VfU�3�;^v��A0�'WbA�C�U:]q���"8��x�oū?�<��Ff
!Ap@���	gH<�%(X�s2��V�HI'D�9'	R_̓I%L�w�\��U��g�o������!;H��d�Ň�m`7"O������N���D<��l����N���i!Ď�HCz����8�Q>˓?��$0v���� C�7R�R؆ȓL�.��u���v� �Ȏ,#9�	�'VR����	 ?����I�6�2}bT�4�
�{�O������d	*��hS��=�%s5B�AP�w�D�M�а��'"��Oǝ}Qf�7�T�YK`���������*�S?Ct4�0���d���1�̕�X(�B�IA��Z`cP)2��a¦a�95�����N�����ӵw���@�@D�I&
Bz�C��.70��ʴ8d5��P5��ix�BV�!��<�Ԥr��q��'X��a*U�HFx�d:-��KJ&(��ؒ?\0��	7]��-���)�!�@/hjX�Ɂ!"Vq9���x�ў0"�ۅFpR@�iD;$��
R+�v�-�P��Py-ߔS,{���u{�����?Ya%³q�pa�g.}��)�-�D��4fѪ}�	X�a��NB�	K¾hj��ˎ0ӄ�1q.�Q4*�7]|��欏�v����I&0�q���[�dy�c��Kr���)mL�Q�� p�T�
��?@|nA�%!ԸI��5$��Y%kJ�z�����X���,%ʓM�^�	�+�O�v� ��cCk�65���ϥA�Ʃ`��A�yb��j
e��J��-�&��w!]�a ǢV,�P�Tk�<E��{��2@�O>i�~:cV�#�:E�ȓ��)�d�
V�;��P�`b��%�0x��];�� ��	4S��|I6Ū�z�s'냝'8����-|��h�->-�C5e9z��4���V#����'`�q��H
`�ҹk�7J��d��gh�Y�F�H��ЁȖ�R3�:���aÕ�
�bU"On��bEX����F ��P���,S�<���_h�S��?�d�
��d��n�q� ��$�EE�<���D"02�[zZ���/L�2�f���+P��p=��N;��h4H�!8���I4�^}x��Y��=+ ��I��3���sPk�-m�DۇFC��yҍ�My2�x�M�-y���#ϔ��y��,�e�w@
��HSJ �y��N1\�RѲ�+�� rU;���y2o��{%IQ��ĉ#Y(�
���y2���m���Ƒ'��r6�A(�yb�ͪ��Ii�CN�*hF��y���!26����:�^���_��yҏ�7V�0���"<>�����yNA
E�p9[GE���X��Ѭ�y��fyj������������y
� x�:��UEBXS(��%f�A[C"O�i���0t����
7�9��"O,�9w��a~��1���7.��S"O����E�kA��02���hj���"OF�yC�O��@����i2 �b"O��)�$ӿ8�Lh��)Τ�v8)'"O�pQ��>P��-P���v� ]r�"O���5��{R���(�*�Г"O
iE��1��L=(n� ��"O��'c	"����E�(S�`"OZ� �ɥa�금�Z'8��aH�"O�!����8�p
׃R�G�B(��"O������<#צQA���x�|e! "O�ux�oߍ�.=�t
@�҅1�"O���ѦC>b2���I� ���+0"Od9��M�faSëQ3AvP�U"O�Y�7��M�P��ɗ!cHFفG"O�mz�IZ�hab��'H,���"O������?xP�;�$�~0X�V"Oh�+5��& ��=iƪ�;��!�"O�Q�L�&S�H ��pC�-"OP���1 8a�TM�DVqa'"O~����Œ�@!��˺2;^���"O*\!���(l�h��6D�]F~
r"Ox�'�3�ƌ�a�϶?$zDi�"OХ�!B��@$#���ΩH�"O�ЂvC���#f��2R��Ա�"O�z��K�g Ir���0���"OH�c� �$F�FE+�\<`�Px��"O ��&��'��dT T���ӣ"O"�K�#������C
�0x��)�"O����ō?!��z�L�v��iʰ"O� �)w��p2s�F���,��"O`,AtJ�s�fX�e�؎D���"O�Q��'���R�J`�q�"O����Ĕu�B����' ��xQ"O���eD�M��|r�$_W�S�"Oj|e�CT��L�0ZQ�83"OF!�R��ba�=���Ӛ=율�w"O01�a�Ϟ�Q���X�-�2�k�"O�-jpف/�����L��&AD 0!"O^�PE�(,j��Eʑ�qZ�cS"O�	���m ;���gJ�p"O�l�j��76�#�ǌ�^����"OƈQ�KG�8�Rw� z����D"O���͌=���)�Rh��"OjtY`푠Fb�i��<Mn�!�"O6�B���Ij�	C:R_��3u"O b���-���a�BXP�"O�h(����'` ���W3�x��"O�a8�D�N4�<����5N.��"O��0��
�/�0��-M�7
Rl;�"O��;����]�H�갫ʿI�ԌA�"OHH��D��=@y�ə�`��9q�"O��#2�$H^i���#ZZ����"O�l7K̝L�3�DTF���A"O��3&a�4�&I��$��9����5"O%ۖ(��kF:�7�Y՘��"OPU�t���d!�,ϔC����"OV�G¨x&�z뎶k�`PH�"OxTr�<x���z��Q<A~r��G"O:�e� �jlj�Ɗ�S�b$	G"OD����r�R(��dҎG��A�'&�y0�X�r��y�����o�~�E���)T��5 ��� j�P0�Q/*�t��E����k�"OPm�^�F�����ʰ�Qˑ"O*�ki�Eپ�ա�4ug"O�ze��0B:� �t�g0��"O�k'hU,�*H�e��O*�1 "OX�5̃�+bl�aB�A�p%�He"OH,���Wa۳O�4*vX��"O*;��D<_ |`֭Y/��E�"O�ضd�+\��c��Z���9��"O֭���ƈm*,�d��7�nt��"O�I�r�Y�-��H�#,�Ӫ,	1"OP����S^H�)C*C�G̲ ��"O@�D Aff�Z�������S�'5�Q-�2��ԃN�Ʊ���O>�����3]N9��y����c�=�Į�а)c���%(|%1� ����I�KQʧv������t.B�%�7N9\fX��hW!� 0Xa��y�@ƥ<�t!������ �EŊ�pP!D�|���S�D�$�dS�O��\+k�̫��Oy�3�"���= p�T1w|��˩O�� 5�A+����s�N>ݢ�.O,c�<�(!���6����c�e���u�ا$��[�ƴ<E��?i�B���L�aN��H$!�1j;P��FĈX�Fy��>%>O�ΞuC��г���6Ԍtb���1
��N(�S��Ms��ߤUO�m�����wG��s��S�<�AG�"���Pa]�jl5�D�<��� %3�hda�6hn(4����|�<a�� N�m:�K�6�D\�$JQv�<���%<8;��4�ș$er�<P��	^�r� C�UB�B�z��j�<�#�7Gu
�\�OB��r�L�g�<y KO�b��U1�K� X��Ȃ�d�<	G�~�ܸ@,_�} ���GCb�<�a/�z0R�6
��h"� �V�i�<i��i�tA;d��Rt�B�g�<�p �?:�J��%u��"�·I�<�����$R���<�� pS'C�<d�WlQ�q�%��&�т�F�<���2w��$+ch�	H��0U�n�<�&�"�,���I�0D���-�m�<�v �%7�e�DX�<�(�M�<y�36>�`��*��4��$��gT�<1/@�q��p�L
>��Z�
R�<��l"��P��
��0���O�<f�65r���3��X�d�<�`4m�D�iZ�7�nl�V`�Y�<Y��_;X�r�b�_�M����!z�<	FQ������C11&�3��t�<Q�H�Ft�,ц�� \���c��W�<�ĵxq(�k5�N#v��[r��T�<��� ��D	C�8v�����PM�<�蔋@ Bi�v��2��0��`�F�<�p��,�����eN�z�
�]�<�DnTO- <�Tg����%�n�<�1�%@T��u@ϟX�B�4D�t�<��dƥ(����jݗk6Iba�YG�<�/_5�LtٔFUV�Vh�u/�h�<q�JL�[�4��bgNw9*H�r�f�<��"�pPx�#��6|Z��f�<y�$`ɧG�	TdX#Fm��&GC�	�H���a��"|,��u�V�!h�B�N��i����7�H-X�BT`��B�	�Jڙ��)�>{z<*��\�b�B�	���y;��ώ���p�؆h2B�r�ȔC @�G������V�8C�I����5�@B��X`#/�C�&��Yy�ќ!���j�nZ�6B�)� ��A�+� ,�tz���*��e�2"O�= �j�*y/^1zSB��,�Iu"O$���$T��yGǪ7��iR1"O�lJE�8fY��E�A��x�"O*�S�h�0r���#�-ն\���2�"O�eYW����[�@�谹�"O���p҅j%�Ask��r"~=�"Op�4D�-Z�ri)#��)=��(q"O�e�b�6�4H�P��JW"O~t�p�J�`:�G[?)���7"O���%�[l�3 HT��n\#�"O�[օ<$0�p�#)�(w���F"O�{bNݤX�*] T�V"v�5a�"Oƭ���ˎ~h�Q!!��Ш�s�"O�у�'�@O��� ƌ�Q�p¡"O$�@ ��4�p�i�d�C'P���"O��䛥!�,�!D�f�,݁�"O.���A�C1VB�)6%��"O��҂C�37h���߬R5F4�6�4D�8��
W�=#Dmk�A=pr���4�4D�\��b�?lv�g��A��R�=D��8���)Y� ��- YVe�O;D�d�w�Y�ІP2��*`��Jg�%D�h!�(I�4d�C��J5j�sB9D��;�J��N!`�*0*�F�!�4D�$��-�0 q���"͆2U�X<2��2D��A�Ǌ�P�Ӧ�Ĝ9�U�2D�t
���I� ��;jZ©2D���ਆ�U�cW'_K��px�H1D�xK��1t�a���Z�g��d�U�-D���VG�#/+Y��(�f�t���',D�`��!"�X�o�o��3s�(D��!�Ԏg�	�i߆\��H��#D�*�j�:56x�9#��/G��!2� D����鈂S���:�J��>TP?D��0u�@�s���h�@�8J�4��n'D���P�2p�,�$�ɍ(�ihw	&D�\R"-^�9����,�/w��y��0D�<��BH68��5E��+l�6�,D��(��D8�����
[A�A`�$)D�|J�m�$TZԃ0�M`�h���*D�@!2H� tT��ҁo�3-
P�p��<D��C�ȅR�D��@�$�^��=D��Cf��>0`���oVI�,��ă9D���R�zH�ݘ�bV:,Z
H�$#D���#�P�5���I�f�yC"� D�� ��-�xYÒ�)V+����?D� ��.D2L>~0�	�t��lI��=D��$����)Ӕ%A��!��.D��@	a쐍�щ̙Ld��Ʌ/+D����bW�76���I^E~�9��)D�L��i�v�4j�3�B�3sl<D���pKI�[ $ݱ�(Zi� 0�Q�-D�L�bܳ�Px�B�`B�6�,D�[#��?\F��Y��ܣ@��i��/D���mӖH��I����qW���q";D�P��.AU�L���Q�g:r�ҳ#7D��@v#�z�f�"���!�@@�'4D��Pb��� 닚Ah�8�d=D�Pi1���1�j΀L~��@�5D�4bd�|��b'�f��V�(D�|�v��p(�K��@�~��x���$D�� U �h�0x��k������>D�,�œ�>�X��T�]�Z�:�k'D�� �4�FfW�Gb�q�P�6�~�"O���A%r" �Io�ȭ��"O@�@����Y����`IݷL�Fl��"O�x:���5V��xi�!�FP��0c"O��tB��{VcG�
?Q:��B�"O� U�X�I^Aڑ/���}[�"O��S�M�WR����m��
�If"O����b��R$��7�TG"OJ-r ��X���㨛�>I�C"O������'g�$H`j�:]�P ��"O�9�`��0��d� *��\"�"OF}{�`D�KF��B(ˊb��`9#"O�����V, �����l���ea�"Ot��taXiN���D�|��"O^��Q��6�:1�m��P��`�c"O��BvF007�$д��S���a*O�̰D��_(��A�ř��� �'�t�x�Fʛ��4#.E�NH!�
�'1�Q�%I�b3�/L*2�vT�	�';����3:�q#EL�5��!��'[���԰\�<�+�C�1�����'됴c�䛖?v��5D1q�hk
�'E�@'�CK�8��^2%>�{	�'����,
�REQ�,ϣ�LX+	�'%ҬSA���!�R�Bf����H�	�'�R����:CFe#V��LE��'�z5�u��3\*����I5���x�'\���M��)4�����4` ��'N<��K��K�Y E/�+_�͒�'	���WZ�H�d�^%Ge�@�']�6$/Z4�KWc׿�((��' ��H�J.!H���FH��>h��'4��m� ���~"�9�'��t�DC�{�&�p��D��j	�'ǀ5#�/��hph(��L-*���'`p���j�>����ޠ�0�*	�'����"Y %z3�ㆁ����'Sp����"E�8��0F\�x?*lK�']�m!���RT��w��#B��'5n|�d�2N� ��1�H��p�'��ũ�C�lX��Q
�k�'�Q�#� u,`A���(p Z5��'	
�!��G�$#��)�'��j���
�'Kr*��N�̘0�p>��y	�'��D`Ӏ�l0\���m�����'Ry
Ug�F�؛F���j��49
�'�B��%*��M�8��fZ�2� �	�'H����V�r��ȣ��^!+�.�8	�'W2В"Ǔ�X��@��(&xpɫ�'���8p�׀W�b; ω�����'����q�P����Ȓ�S<�		�' �U��A\+�1�7".Z!�5��'��a$̒I�b�����GQDu8�'8I�G�k�Je�d*[�T �Q"�'���0�ꋘ\E�l�S&�G;��!�'���S�	�/�1Y�
ӥD|xd��'.d���,ڮ/�I��g9Rܲ	�'�R���>L�� 3+Z7*)i	�'r�B�hUJЙb�ʏUz�Pp�'3l�`��	ht|���N�G��	�'��p1��D�!(�QJكE9�e��'
4�©�9"��,X�'��]��'�6P�H��
"��@��%����'�hp�ŲP��� ,�
������ P �b�A8�=���� O���@"O����W&�x���~B(H�"Of� f��hz@���凈9�ݛe"O�q!����`R�IQ�5'�I�4"OHـ�/@�vIͻ��L!)��)A"O�Eh0��=����%g��a��]�a"O���Z�F����%FT;�j�K�"O	��(0�ڴ�_���"O��j��mir�c�C͗����"O�xB�`""���50��A"O�M�Řb{�y�é#m�T�"O>�� Y,l�VA�6�[�s�$�"O.-�� �p="�"Ҩ߶[�^	�r"OJ`S��% ue\Ӧ}��"Ovi�	�a� qYE�Fˈ0�""O
E�P��ti{u��.s���d"O�)�"�G
LҌ<��$ٲd�z|��"O���u� ����s$[�3�mf"Ohi��.�54�j��B�.0��؃"O��V/U�i�Btb�K�B(0Xy"O�PE'�;E��`���85#rp(D"Ob4{QJ	9||�E�΀���p"O�1 ����؄L��B3v��`�"O(��F��H�J����$\���""OZ ����,�,<s�ш�2�Q�"O���"�=V��I6���f9"��"O�)��n�fv�R榘�.Y3"Or�b��@l&e����2��K!"O@�ҕ   ��     Z  �  �  A*  �5  �A  RM  �X  �d  p  s{  �  �  �  ��  *�  ��  ��  �  Q�  ��  ��  !�  e�  ��  d�  ��  m � > � n  �& - f3 9: �@ JG �Q L[ �a �j �s �z -� m� m�  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R��'��:�aɤ,��`vcء|�~Id�=D��Q��ˌE��z%O/Fs�mQ�7��)�S�'XM0�UhR: t�3��UU\`1�ȓ���q���*T <Ia�?c�ؠ��3�� �W���TCԺ����d7�-{G�0R�
Ը��̳c����N
��
����J��8�2qz�=��wYu���'R��r����e�4݅�u?��+Qœ�M@\
1�W�1�؅�h�eI�*�~UZD�����ą�T���Q�dD������(m��ȓ	��Rr+���<�Aj3\�Q��I�}Ru��4y�v��`E��2�b��ȓ2�,a양^�d� �N>Bņ�Q����$�Go 4� ��@>j�ȓZ�X��%G�,�Xd��غ"t�5��W# Ct`�A���X#��rg�-�ȓnV�yC�U���x6k�[K*��ȓQ^@d�p����sVl݁oVr���b2X�3SMD�=f8a!���t�ȓ0����I�<�XXC�
�Q;���ȓ�"��w��7+�dȘu�ȷ���ȓ;Ҧ ��B��IT��(��D�꽅ȓ9قu1�f�y_t ���7v��P�~- Q&�Y�F4���-wq�(��@֚,@�ϔ.���V�`'p܇�l;��GD8!�,�w-J*�هȓ5��S5!O�tk���f�<z6�ȓ~t�i1C�M)><)��EJM��{�R} �L�j
�*3ѢM%r�ȓ"��\��o_�4�WbD(l��@����<��;-o��P��&>�����C �3�^�A� ۤO��X���ts�*R)G 0�pHb:�H��?y
ӓA��Pq�*K<T��@e.�'�r5�ƓydI��C� uj���� �A���'7�	P!H�a�������far���'?(��]0:|��F��6��
�'"2���a܋,��aCN��
lL�	�'�҆�;V1�@&� |��TP�'0���"#�"�d��e���'xv%;	�'��$�߸s-V�!K�I�����'i�}�# )�j̓��_�@2< ��'��p`��
(两j��0=l��'Z��)�� �K��{S�L�@�u��'�J�#��D3.��i���ՋlG�
�'�x��&d�0:Ȗq�f&I�a�fԳ�'�\1Z�M���h #L�	a�9a
�'����'�<�,��#��I�*(h	�'�X��7gNa]r(Kr��F^���'-����;�t��*ԑ6Y0���'���t䖓e����FD�y��X�'È�r��4f�� Yu�
~�Hq��'�$3`�W��б�1b����C�<�AW�Zo�h�5˞1M�xS��z�<����6 x�y�� <�|���d~�<��"J w��@Z?&�HP뇦^z�<�0!%B/���� ��X�'��n�<�DD��c����-�{���1�E�<����;-i���g��n&�pT��H�<)f�<ؠ�h�s���sb\F�<!ң)]ݬ1A�m�$gn��P ��f�<� L0�i�3:���b1o��O��郢"O�A��M��]��8�-k�l�v"Ort��
D8g�\T��̜�f?���"O|��V$�9m���a��%
6�ɱ"O�Ī��$$���2���D�l��"O��)�ce<H=b$ٲ+�� �"O����Ο�t+���%�5}ò�ڗ"O��4��M��A�#J��t���(0"O����*ٗcJ��p��d���s"O
�5����6�h8Wo���"O��A�&Jt�H*�%�"j8	��"Of�->5���Th�hC""O��w/�p L��g�
M�$� "O>�`U��c����g̈7�v|x"OƜ�� :�)�k��E���"O$��0��<,��H=�� R""OX ���9^�H\h`Ȝ4��xIP"O���!�Y5�`��D	�6��V"Oй���X"	"m��AI���"OV��Z�SA�!�Bs��"OМ(�F�����*<���x�"OΩ�X�ޙ�4gW*���Id$PU�<�V�O�~�	�d(	�3Ѱ�Ɂ k�<vCʚQ��ݛyu�#Ak�i�<���<&�8a���yf!0���@�<yG�t���b
�S��U�<V�['g�Ȝ
 ��Z̐��FT�<�Rɝ<Gt$�#͈[Wꭢw�v�<��G%)�޽�5�ϊj��ⱍ	v�<y��0E����i�{��pZ��s�<Q�W {�j��B��y�>(aFU�<��Ɩ�5�"D!������ÊW�<YGF�y{��0���8�ɡ�i�<YU��%"
Й B<!db�hD�e�<���;1A��ӑ�ɸ�@ݓ�JI�<!��Z2q�@�D�$I���p�<���
�T'�ٓ�Î,B똙��N�i�<�	A�sP��Sũd4����y�<! �v����L'��5���O�<q����BB���j�v�"a�K�<��#À:�Z`��dݙR
RIȕH�<�e���#��8� ,��`q6��A�<Y"ݧS�i{v
�D.t�B�NA�<!2��>$R8�'Qx���
��W�<IB�֏}�j9�X?f���JB�Q�<��ȏ%ҭ���O�d,�Xc�r�<�e˔.ta�'��!HvZ	��S�<QP�_�K�B-�W!ٝcD�y��GL�<�7���v'ĝ�%�ΩGwRB�	Pd"Lq�J�H���k"�� :��D�[Ԝ�yP�8v�T��:x�!�$�'9]�a qHС84]㷯G�	�!��[��� �fK�56Ͳ���H�!�$�����P������p��܇r}!��50cX ��!�=;	��ZUM�g!�D�%!Z�u�����)ԭ��>�!�D� w#&4��ȯ�t��D��!�$��]���ȵF�? ��ٺE@S<!�d��Qj�%�E��(f� اF��X!��	O��C�A�]i��q�H�<�Wg"��u�ͅg:�T��g�o�<qGO�1�؃D
߷2�=���j�<�b�l�N�L4`B�Uç(�f�<��Ά�!�������8XN� mH�<� �s���Z|Ä�R?T���"Od�ڳhL�,n��֮	&V�&<pW"OX��@�3�����n�,T�Bw"O���w,K�]�P@Q�,жx�2�PG"O^�B��D�L}�,>����s�'���'��'�R�'���'���'��Y�̊b��D"a��?�@a#�'���'��'��'��'���'�F����)�� 	�!�3r,|��2�'�b�'"��'Dr�'���'&��'� x*4m�<$��B�i3�'���'4B�'t��'2��'���'=��I���B��q	�-����M)1�'1��'���'tB�'���'���'?r�
c�KX�<��k��:��M�'�'���'��'E��'���'���'����g�6m��@��եO�A[E�'��'`��'�"�'[��'��'I�0�� �w;T�S�+��I)���'b�'���'�B�'-��'#b�'�m� \<~=3�
;��c�'/�'U��'W��'���'���'!f��HU�1��}��c_:�~���'���'!B�'W��'���'���'�ˆFQ��Y��L@�8�n!�e�'W�'���'�"�'���'���'Y6���NL-+�V�z�ɑ���#��'���'���'+�'�"�'�b�'�\sD�&d�c�\�e�l��'+2�'���'7�'���|Ӕ���Oҹ��ܽ�6	iT�S]!b< ��Ky2�'h�)�3?Q�iTе���z��,�d,����,�C����d����?��<���}��i�
�b��\���یJ�4�����?9��Ѫ�M��O6�.��N?����\ ��Ȩ��͞3�p�+Ql<�ޟ��'4�>�-F0�l홗M�rXP٘��Z��M�&�m���Oc�7=�\�{��͝Z���O��8�2&��OX�d~��ԧ�O��D�T�i�󤙑D�D�y�,W��y����v���e��z�g)�=�'�?�A,îu@�,k�^%l�p�`����<Q/O��O\�mZ#7�(c�����	��[���z��h�n�����ݟ���<y�O��`0��$�Ȕ;��Mol�}Z�����	�J�z$���(�J����ߟ|9�
 OD��4@��Z�&�Wy_���)��<	d��Y�0|+F��=$��xpr��<��i��X��O�-m�}��|��kĿ�ޘ��-p� I��+��<����?���A2f���4��$>���'�hacG
�u# ���۠"�]�D�6��|�*O���H�.��Eu��YR+BT]*Mᄞ�48ڴ(u�q�<A��d��s�]�D��:L��(�K%A����?���yr�&zs�T
� �y� x ��R��$Z�BQ�������U&���?i�o*}�gy�� �&�Ƞb�1V��/�1+"\�\�'*�'S|6-V6c�Z�:���#�ڇg�D����6s^���U�?��<��?)��L;�b��Jr�=�Ƅ�)��y��_��M[�O��$�����)g�����h)<a�6��7�TP��i�D�IFyRQ�"~��n�?b�� w��" ,�	�S"f̓�ƣ����$�¦$������q����2�)�@��0�O�<�O��D�O��ΓL�66�9?a�� �G��~�P!�VǞ#R�訉@�Ox��4����?qTa��:��Ab�/�h<n|�WA��<�K>�u�i�ꀺ�y2_>ia���b�"MbC��\F~�D�"?1V�����|ϓ��O�� 	B	L,C�T,�f`E8I2�1��'@LPJ�M����4��������O����I!H$�q��;"�R\�5l�O��Of���O1������H�+�N���6�LT9դ�
i�`���'��keӜ⟠3�O�0mڣ!tz�x�N��Br �i5���,Z�Rڴ�?�iS�M��O^<��� ��H?)8&!_� U���q��2���bs�Ȗ'zb�'G��'/"�'��Ӏt�>$��ň&h8x֙��fґ�Md��?A��?YH~Z��Y���w[���gg�*N����2J��tM� ��|�,�l�w�)��]e��l��<yW�^�J۔$���ƇU�u����<��-�"mv��W7�䓂�4����
2�\a��d
�d�d�i'j�e�6���O:�$�O0˓l*��
���'���kx�i!�$K]QST@LS��O���'2h7F��q%��J��]�u�``QkP�L���1�h'?��DY |��*`��]�'d���D���?�!�&E*8"���$��9r���?���?Y��?�����O��RT�=Ft>��d-[�Abfh���OoځT�u��̟`�4���y�OFW�"�S������92EƠ�yB�b�V�n���y��㦍�'��(B���?q��ڿ`	h��f�*	[3х��e*�'\�i>���ϟ��IßH���}�$�r��u�$�j�N�j����'�7�
:n��O`�d+�I�O(�`�ǹ}�L!�@+�R��J�Q}b�i��mJ�)�&��Q�P?������K�H�%��`A'!9?�ta4;����D2����dX�dx��>6��\�4jZ�f��$�O���O �4��ʓ��F�
�� �p� t�E��z�̘ �I��yb�aӲ��O��m���M�d�i/��jfnș;�Z�A�8���vMWL����O���#�H?o1�����{�v�N�� ���AL�Fy`ek��תRdnH2O���O����O0�d�O��?icFkK�M�ѡe�,���{�\����	ޟ�P�4'V��'�?	��i(�'�0\c��>Zv$jU���x� Ȓfn#����	��|:���M�O�ax��Cb�\]�`*غd�֭��ǔzRt@�� �O ʓ�?����?���./�e��\��	2�G�6{�H�p��?i/Od�o��3Y������(���?=��5��T���@"Y6�T�bT�0|P�n��I�M�ӱi�lO�Ӊ.��E���n��x��'g�6��B�ؒ5p���&M�Gy�O]����2_�'10r'��;84`�̆.cՌTy��'aB�'�b���O��I��M��T�)*�]��ӗC1�8�R�RLPxP���?�ƳiW�O��'ئ6��;�t@{�� N_X5r��E�Q:ʱo���M[���M;�OjL��d�����<��e����LϺ}�|5�r���yBZ�\�	ߟ���L�	��P�Oז@�F��$|
h)2k��N���07)o�6Ԩ���O`���O��I�|��^w��wG�h��֙	D��@�9H�P�sd�Oh7��q�)�	��4�07mg��XW�[�rh�Ss@J�i�^t�v!q��*w�<7��G�	~y��'��
dڹ�p�*����p O.Aj��'���'T�ɚ�MctF��?���?I�B�TZ4 ���	�i� ��s���?AM>I�]����4
���3�$O�T���d�����X8V{�	w��cb��p�l�$?�C��'�l��I,,Q$Hi )H��3���RMX0�I��0�	�d��x�O�"�*e1��q�ǚ�-�
 #o��n"�y�Tx*���O��������J�i���4��+y�5j�f�\F�<`����L�I���ݴi��uڴ����./Z"���'��X�/>2,�wC�{���.9�D�<A��?���?����?a�.($R iB��xT�������Iڦ��/��h�	џ($?a�	�J6���� ��L��Pb��)�Pd��OH�l��Ms�x���h��gPAcdC�$���#q-(��<)1U� �	�H��J3�'Ђ %���'��L��l��F�\���iə��\��'�B�'�����t_����4d/���,.��z4��{Dy����w�V��k����d�h}RE|�^qo��M3��;[ϊ�e�ڿ�Q�X��9QR���-�'�bͲ�O�?q1r����wk*�1�)=C����gD����'�r�'/��'?�'Z��T!���7B5�Ű�*�f1ۖ��<i��͠�a��d�'� 6M#���s��p���r����.��M�=$���ݴ@���Ok���b�i��$@��)6\���h�fU�q���#�l�:Q�I�f/����?q��?���d�H#͒��2�S5W�1 Ql�O��$�<��iKFD:�'*"�'�哣>[�I��ªTQn�ze���	L����ş�m���S��)#F�F���	��w�bbƇ��x��Qj���7� ��_��:>�"O�o�I�B�|��򁀓B'�0����:H ��I����؟��)�My��v�l	�U���|, w�U�5=�a��J�N˓z����Tm}b�h���jM���,Ð��8N�1���ix�4g5��4���Ó��<��'4�˓Y��{0K�;I����@́\m 8ϓ���O
���Ov�d�OP���|��;6N<�R�F<�����-+��-/gC��'�����'��7=ﰤ1���4�����Tް}Ғ
�ڦ���4;f���O�~0���i�����F�z �ƸO&��rT��<��ĩq@����K�2�OP��?Y��V>xx��ѫ
2�x��'%������?	��?�(O�nZ=dD��ǟ��	�'�D%����bZ�yǊ��x�̸�?��_�$��4����=�$�2��0IQ �J�L�#A�m���9��zF
(�~�&?]Z��'�~���y�b� �g�����N�6R�la��؟<��런��^�O.Ҁ`2:�ڒ�M:�u�0�ιO��e��s��O"�KҦ��?ͻ5_�,a�GZS~�+%A��.��A�F��F�j�ZElZ�ƴ�o�A~�*��C"-��%*	Ô�\,n	�7Aí[
��AS�|�Q�P�I�L��ȟ|�	۟8X��'K����Y�^���H�VyR�iӠ����O��D�O�����C�p��MȲC�?�fy����=*��'�ұi�O�O��WC�!e`t)tJ�;^:�Q��Ί��|�RR��(�eI9'b�
Y�IUyr�[Ol�ԣ���8��a��+��'�R�'��OW�I4�M[2i��?��l	&y���ǋ�9?fq�R���<Y�i��O�M�'3v6mB�uQ�4h,u
��8u���a�A�:�(��re2�Ms�O�<bD
�
1N5�������c�ɀ19��#�EJ��E0�2O����O���Oj���O2�?�a�m��}6���Я�:X��az�kZy2�'�7*����M{M>�������J4i�y�*���J��>����M�Ӻ����T�P�����oԓ�`1���ͦ8���d�?�d�a�'5�h'�D�'�"�'M��'D	!���b��F�i��'�2^�4�ݴ��I-Oh���|�S��1��� Wi��~
����SM~�>���i0�6mh�i>�ӗ=O6�Kt�Z�麼qPI�$�8��sEC=/�d	X �Ky��O�<�I:n�'���1d�c�(��{b�q��'B�'xB���O)�	�M��fW�+��d:B>1Ș0�5,$$@�����?�Q�i��O� �'�N6͛�+`�A��]�FȒ���ҤnZ��MS"�@��M��'^`C�j�(���|��)� Rh``�2m��hs�+?:ī�7O�˓�?��?���?a����3X��� ���Yc��SaC�d�o�8{<t�Iޟ��I]��ޟ�j���˄��2z(N%x�`ݫ]l�T�L�F�eӎ9$�b>-�p�¦�͓�Q�G�Y�:w�͢R♱{����zԪS3'�O��M>Y+On���O$ z�d�8'/�5��
M�ZTr���O��D�O��$�<��iB�{��'3ﬀ��&׾/�j ����v^B�za�dkyb�':�6��O^� 蜁#��]�C�T��H�ol�H͓i��xTL�mTI��·�?���T=+�KZպ�p�'&��p��Z�x0ZQ2�ז?`<���'���'�r�'~�>��I2L@ʉ#7�,:VŹ�bV���	�	)�M�M�*�?9�N��f�4�m;�mP,S��c�_/�$�Z>O�n�MK'�i�p�Ȧ�i��˼ ���\�%C�m�w�RTc�L����{D���y�����>�]�<�	ß@����������Ic�c��Da���H{H����TyR�ӔBW:O��d�O����d�{ؙ0
@�+Y��r3��CŌ��'�J6M��$�b>�� �K�a��IJ�k�^8�cI;+v���6+����`녱*����&[κK4�>ɔ�<�'��Xx�51���r6.�^���'���'��O��I�M��`�<Ʌ�-$���tO�5hv�D����<���i��O�ė'sR�i��-ϙ,f2�2aհV�D48am��(��Y;��i�I�Z�����Og�'y"���8 㝱np�dd�9�ԡ>O����O��d�OJ���O6�?�G�T:zNR`9��0jt��)�-7?���F�a����¦&���@,�?JHL�cI�m��I�v	�j��M�Ľ���'V�v�v���� 	ߣ3�t��$N���|�*��W�>4J�2�'�T��'��6M�<ͧ�?���?��&�1@��)(���
s�x�D���?�������m�#�x� �����O�%�w�@|�J�f�/c4>�h�O�̖'�i�1O�S�g5�x��k�N6 �d�V	4���xf��@���*?	����@�'V�Ӽ+���()#El�@�F��V�W��?1��?���?�|�-O��n��j`�[B��qo@�;
_�U�n��(&?٥�i��O��'Ǜ�D�0U�m�%�Wt�q��;PI�6��O�d`4�xӆ�,��z����OXѪu�U�+���S����	Ν ��u�"��?���?��?I���)�Pܨ�qD\�Z�r�B��%t��m�"~���ΟX�Ij�s�(�������[�U5ڥ���эmb��C�B "J�i]1O�O�D���i��$�e�(X�pa
(0^�R��ܗ4���ƕ ����y�˓	V��W�����r�ԣ{�H��G�\iĈ$�՟��	���	ry��xӰ�`���|�I)P}t1�Mǭb�d�i��
1A�4��?��X�����%�8@��۸,Gd�7c���L�d=?�!j���i~�a~��ۆ�'HL=�ɨu98�+5�q��W2]>�hR$�O����O.�D�O�}�)��H*N�l�)�q`�?Q'2��@қFe܆��� ��?�;Wy��G�ъ{S��9��(3,-�`�v�j�X�D��U�z6�=?YK1>2<�iY(~!�0�&fS�����!P��/O�ImZ^y�O#�'H��'�R-�=��}�0��%�챐�OԚ+���5�M���<����oZe�s�D�§_�B~T'��D�.���������j�4��Ş&
V���ĕ;AqP�K��8(q��:k�Ph�'���x��D����`W�@B�4��U?q9� ���;'� 2F/ޛ*���d�O0�d�O��4�`ʓ'���(��l�R�ُ��%�"������Ѝ�+D����⟬��O�mZ�M¼i8:]a񆐐TJ�H:0��X�hEٿ>��F��pѳ��	N_�d���1��׾8��	�P�N�N���8Oz���O����O����O��?]��>� �ಯ��?� ͒EnNş��Iȟ4hڴMl^�ͧ�?��i�'{U� ��04j�	S��1EN�q(�1�Ǧ����|�5�Fβ"�%?��(�Zd�@�JXa��I�&�x�A�O,Q(H>Q-O��O�d�Oځ�Ĩ^$:2xT�CE��O>B�i�A�OX��<)��iJ�tk��'"b�''�2h4��uM�`����"'��3��|��i56M����M<�'�z�㝪@w�TP���jT���@�8?���t�ߔ^6��'u�����<2Q�|��P� �@��6Z�`�ゥG�"�'r�'x��T^�x��4z���sa�z�M��Ԙ>�q�u�S�?��-����G}�t�$|��Z��c�Z�k �p���J,'��.f�A��i�"�ܟP��&��h����+?Y3��:Rr����HY]Ŵ-)&�A�<	-Ov��O����O����O��' xl���D�r��A����X!��iG$�hp�'���'񟮸nz�킒�]:A��c�߄D����6�MK�i��O�I����逼+��6l�X
�f��,���!"� GX&��U%o���K�"j�dB�	\y�O�R�ڜl8��K��92�h��h��f52�'���'����M�'�U��?I���?iEi��9�ݑr�\�R!^���'0�o��6�m��U'�lq��5_�� B MƑ	��g�o����.ldP��]z�d��zB��O,���Ae���AJM�&��P��ղv�8�����?����?����h�����P)vT���*? NH�*4���d����S#Dɟ �I��M���w����-�'�^	 N�3E�h�@�'z���eӤ�l�pA��mZ�<�q3�(:W��X�� ��1�)��sA�EZp%�/���<�'�?���?!���?!e� ��0Zf@�n�vA���H����ͦ�K/��d��ϟ4'?a�ɱ��@R��ۺ7ۈ4CgO�(JIҨOV�mZ�M��x�O��T�O"�Bʇ1ʐ�2� β`y� =a8|8x�O�e!��D�?��b9�$�<y��$G�
���_�E�:\P$ ��?9��?����?�'����e�&�V˟!㮐S.L��)VY����џ�Y�4��'>L�L��Jgӆ�mZ��B�$jߜ!(&����E�m�f�faK٦�Γ�?��mΌ*����~~"�O�) c��d�5��mRx9�.�y��'9b�'���'�r�	�52�F0Xč�ZBgbߨ+q����OX��m��n>��I�MKK>QQK(T�$���W�����H2$�'�D7M¦e�-9��l��<��%��9�a�f�8�H%M�jE\	#�%����䓌�4���$�OD��P��T��Lε1U���$��Yw"�$�O�ʓ0�����Vb�'��R>A"�*9�x"b�H"�FI�ѩ(?Y�T�H�ٴaI��j.�?ŉ�"�Ձ�ֿ;y�dIԢ�ubU�g�o�l���O��?��/�d�#��S
Z�D+�%���-9.��O��d�O`��<y'�im6��LF	bFH���@�4l��j���>�r�'R�6�>����x�����S9�&�;���Z�,�H���eٴ=�����4���g��{������_̜ ��
4(�xdH�ʖ�bb"�Iay��'���'�b�'%BZ>���ȗ�Gr�+d�
������Q��MS	��?a���?9I~j�9���w��Pf�E��P���5e��i���a���nZ>��Ş&�plZش�yR��|sR9�T+P����yr'��J���OybQ�������'�FtY�M }�) �S����r�'���'�"]����4g�4Xx-O��DO!V�n	�b$[�6.�A3k�WA��X��On mZ��M��x���U۔,�~����(����Y�������E0
/1�����/�ʢw��,�`B£(�ĝ��)@�L%4���O��D�O��,�)�Sf�9�*��2b-	�}K�M��ly���U��OFn,O���՟T��I��֟�<s=&M��Ń<����Ǯ+�l���Mw�iO�7���F��6�{���ɟ`Dx���O7&���
_�P�Daz���?�,���z�Ay�Ogb�'b�'��A4b_�m�G�E5*�����e�.��	��M�$k���d�O���d�Ҡ�k��� 6 ��ч��;+�9�'d6�˦	ϓ�H�~�(�K"�:9�B��(�y��C�~(��`㝟��t��v�B�g�JylY>u�L8�cH��=iw�1��'�B�'��O��	$�M�`���<aS��k����5�W`�����A��<QĹi��O�E�'�±igH7͕�
�P���;��@���#��퉳t�F�	̟�p�ݠ8�T�=?���տCЏ;n����B�/���1C�<����?����?���?Y��4��� �	���E0d�%�C	A��'u2p�t s3����E���%�8���2\��!�"$x��	��'�����f�j�p�	%"p�7�s���"_�Y�j��>�j���l�:��i0�M�`����M�	By�O�2�'b$vD�8��(��j�a	��'`"U�(�޴_8�+OL���|2���N!fX��
�'���:7�[~�F�>9�i��6��H�)r �=IAF,�0���G���^�R�B�!��1?�'/���$����rj��'�n�,��Ռ�-y����?!��?��Ş���Φx���y�'�Īb�F�"'�lJ�{ț��DTq}BO{�h��(ݝ >�F@։0�&9 cJ榉�۴R7����4�����
?R�H�'����Gb��,�:=�|rA�?f0��Xy��'���'&��'��^>�:�.A�p#dܸ$%ʟ��a$fź�M+d���?����?I�'��9Olnz���H�8�����+��ł3��!�?q�4YZɧ�R���ش�y�#��.��zP ��X����u�P�y���#%�	�_�'&��Ɵ��I�)sDh����+T����w�Y��՟x�r�̟��'�6D�Y�Nʓ�?��I�:��Z��ל+P�*� Ķ�?�+O���By��'��� %��%����U�)1>�8�	̜h����OJ���#ʵ����f����j4����g�0�9�QaƦ���H�����������	̟�G�t�'�`���gX�G@IC��Iq2���%�'>�7��5.)���O��lO�Ӽ�R	Q3T��)�E��o7�Ik2���<A��ie�6�ͦ�������'�ht����?j�h�Dg`�k��5�҈`��'���h�Iꟼ��՟��I�OZ�OW�|��p
�b�p�')�7܈9*�D�O��$-�9Ox\����:X�d&	"i�/�F}��b�Rl���S�'0�����*K8t"��O�Z�ph��I����'��e�M�ޟda��|B]��b2��=ir�P��?QI�i��F�����Iߟ�����Shy�r�.81��O>I���·o!����[9�|�����OXHl�r��<�I��M�C�i�&7��:"�`�hfd�;�Z�q��?�@٥�c����� Z 쁬uL���(?a�'Կ�Q��[q��a��[$)�pz�*�<���?����?���?q��mJ-q��� m)>�jp�E/)���'�R�`�U�15�X��ۦ�&���`k��N$�3̚�+��E�����%V�^<��O��	"s�i���)�� Ԅy�YO|�����3:p"��I�?��d>�$�<����?����?���mKp��fI$�pl��?����J��%b���|y"�'��	d����ߝ6�N�rgJԮ4<��`���M�'�i}�O�ӹ5˨�bEN�P@��+�ݑI���[3�k��x���ny�OC��	��'�t,�@��*h���9�LN�|$l���'��'�R�O���4�MK���:[��P�@�]��ǌD�(�T|�+O�@m���]�I��MK���+��K �R?�b�W���t[�F�cӶ�i��yӖ�)��Sa��|�-O�m�ʺ`h�)Rb�fr�Yp�1O���?���?����?	�����gG���1�!(�zSe�I搨lZ$ �d-��ğ��	@�s������k�E���J�g>���KF�V�vjѵi�
6��D�)�Ӳk�XqlZ�<YqR�e��Q@���y�h|c�N��<i����dǷ�䓔��O ��ѽ%މ�`�k�X�k��M�`V&���OH���O��@��F�Y��'�rm)G *�s�VW�����_'-��O��'�(7FئU9N<فHP8*.�(��Wd���CJ~2��8w��@,2w�OR����2:ES�r�8L���.�����(~�'n��'nR�՟ 
��
�&h���S��@�P}�ST�P��4Ul�y�'�X6�;�i�q(�A&6��xU�ہO�>M�$s��z�4_����s�:pQv�uӀ���y��K��4�N
�%V� U`�+=D(L�Tg�#����4���$�O����O���֣E���
 b��/��:AE��8��˓C���%��yr�'�R���'&�q8p�I�Qz�\s�خ!*D02G�>�շiq�7E�)擘`ZB )A�^�ZX�a�BR����H�a��v�!�Q��O���M>a(O�U6L'0AT"� �D��!�O����O����O�<��i��5��'�4 "g/U5@�,�#��Hr�B�'�H7m2�ɿ��P˦�c�4{���R�$&��BV��(��#M���3�i���B�6���OJq���NL�j��a�)�
ˤJ Nݵ ���O����O����O���'��_"��+��"����H��I���Ɍ�M�2c]~�"d�t�O�9
%����!p1��|~I����c�	��M����D��Is�撟�sT/��l&�@biZ8m���Jw�_�9���^�M�4<�d�<ͧ�?i��?��^"�j`��Дh(E�T�P�?I��������:Dl�(��ǟ\�OFLŰ���6 c�B;V0�!��O�X�'��7��A(H<�O�J�kt�P��ÕI��a%m/S�J�b���	>`��O�	5�?��3�d](^��8�j\Ėc��Q  ����O��$�OH��<y5�i� ���\u��b�gRVʠ �G�y��'"<7� �ɝ�����}�G�Ǜ]�Dd84��kOjM8��'�M[��inR���i���]YD0��O[�\����.Ց[V�p򁠗�2_"H͓����O���Ot���O<���|򖠏7o��d#KT!bNz�"�i�)M;��E lFr�'(���d�'q*7=�<e��dd=\т�)C3��l+�������4U����O( B��i �;j=��42k�XQ���5���1�$��/�^�O���|j�HM�T�t��4LA8�a�
 3��i���?����?A*O��n�NW�<�Iӟ���w���F��U3�	�E��4�}�?Y�Q���޴��v8�C�D$�@�-�`�`9��N��I36}`%�A��*�b>E���'�t��'>%�<��8�N�fCJ$��(�	㟸�I���	w�O�Bg�1{S&�q�Y]�����1}!d�dm������ߴ���yG�˦8��$�ӇD�S��U�F�Q�~"�''�FN|�����{�x�q�PK�(�(���]�Yq�9�D�^�GSv�r'����4�����O��$�O��dO�18��c���8G�y�&ʙ�u7~ʓ=ћ�+	��y��'�����F�$�;#j�&B���tm��
z�ɩ�M#�i��O����Z�Ӆax�b掍����gc�6l4����.+�	�m�j���'RV�%�ԕ'�����:���e�7l84���'�2�'����^�<��4'
�T���Y`=��4hS�"{S|d̓+{���D�]}��n�,AmZ�M���^@�c�A?5}�`r�J�Z��X ش��$�� �������O�G�Y�Q�f0�0��� K%`����y�'U��':R�'�"�IKD
x�LL�<Υ��� |��$�O��D���YX�f5?��i�rQ�D
t �ZZ�!:�C��Y��Y��D�&��M����o�H��Hl�l6�e�����@S�lk!�.HrR�QU��?}�M0�<��'UZ�}y�O,�'���A��6��%��hO��(��'�RX�D��4B8�Γ�?)�����Kn JN�/Q�Ԅ� ��I	������4�����O�����C�+%8�s"b������A�K�v�Q��������H�8��pF�Ox�3���Nr��A!�7J)F�E�O���O��$�O1�l�|r�&��O�>��FC�~B�p$MC1��E��O<�mZt��%q���Mc�e�3V���c��*/��i��N:Y���j�
��d�r�|�	۟��B`�C�dd.?���ʧPl��'�ě.lHi��<9-O���O��D�O��$�O�ʧOV8p&'J�Uܢ����ݎ�Nڦ�i��C�'b�'���y�Ev���dopy�	�HS��qU�(#JX��I����I>���?}���N��n��<� �<����N�ܨh��q�!rp2O�H��Ȋ�?awa?�d�<�'�?	�?2j*Lh@�N!t�x�c!c��?���?�����֦ys�0?�������F'S<�,i��ݿ2����C�>�e�i^7��n�I"Z�����s1�!kEÌ�I�v�I� 1W&�4 ���>?9��1��Ĝ=�?9���%�� z!A��ް�4�V�?���?	��?���i�O�1Ov,���ƌ��Y��`xr��O��mZF��A��f�4�0��ě4O�,�����B���s�8O�Loګ�MCd�iG���i���Od���<��D�1%��qB��.�l�"u�^֖�O`��|
��?a���?��aܔ@�f�x<}�4�9�X�/O�(mZ�S�������D�s�DR��ťP�ó���U�ָj�����@ަIPݴRL�����O���aڍ<�.� '��#�*���Ξ(4c�!�����$�={i������O��{"H����Q�i{*-�m[(�DmY��?9��?!��|Z.OԌo�Y1��	3!$R����*4�B&H9D*~�ɮ�MS�⎷>��ie7��Цq˥�32fV"��-L���;��
$�$l�Y~��\�*�p��SZ�'��Ѿb���G�N�Y��u���<!���?9��?y���?���d�/IR���p�JQ���'�?�yR�'��g���iӑ���ڴ��1���
��.b�
�N^!�"�@�xl}�`eoz>��� ��!�'d⍊���1t�;�P 8b��ïJŎ����3m�'��i>�����\��Y2|:��VNu�DC��r4`���T�'�7�����O��d�|brG�Ԉ��
Nyxq��LD~Bʶ>q��i��6M�F�)rc�/�p��%DՂE���)2
Ϳ56l��P8B@��4B�៨2��| j�C�F5�VLC4/��#��',B�'���4Z� �ٴ݂]�墕�.8*��Å�iO2��L�U~�fӬ�PکO�%oj����i��d����i��'2�P�޴9=���vl�f����L�2d��$�~BB��!�Ľ���T�6�~,��Ǝ�<(O����O����O��$�O˧7l��Ȓ$I�4���9�h	�'+,mX�i�~��V��	Z�'&��w��Y��CR�,)�=b��R�>�Ν� H|�4@n�
��S��".AӦq�B(0���!��!�(aj���Po�R@��O�yL>Y(O���OB`��`�v�xC�Ŏ
D�4��O����Op�D�<�Ĳi��I��S����c�(�:�iY�r�l�h�hG:^�I�?�R��ڴ"���3OT�0�ldqn�;y��|zww�L�'������#�����ԁ\؟P��'W�A����2�@c�N����r��'r�'�2�'�>A��+3�T�Ц�Y�T�̌3%��`(����M+�n���d�ڦ��?ͻ���� C��]mXZ��@�0"]ϓl1���m�0n��R�vs��F�b�a�O�|���)B)�h� ��/O�0 �!�Q�ny�O���'���'i:㢒:'�\ <��ŀ��<1B�i���ؤ]�d��C�SƟ(g×�\�.��w	L���P"E�P���������4H����O��X�$���7$Rh�UH+5���굪�L��y�O�MC���?Q �$���<���_
q����;PgF�Z$�'�B�'Z"����Y�x��4wb�)��:���a�/��@I咥c��0������~}Fj�Έn��M3#���]��A���G6%'(�	�G�;���۴���Ԟ$Z����'��Oe�@�{	��ud�Z�8W��j"��	��������П��IB�'�X!�gA���mzF�Ö}�r ���?9�FV��a��$ �I�M[L>Q C�u�jd�3#S L�2� &-32�'x�7����
Ux�ns~� FN��̑�,))W��Is/��O@����ݟ��b�|�_���� �I��x:�莰��(C��X�.�Ґ�G�����ay�eӊ��f�O�D�O~�'n�8�P��K�D5����%�=i}V��'�p�|�ƣqӄx&��'!'����h��b.��%5�`8r��0@����Wk~�O*�(�	�VU�'︈����2�y�
S�&� 8���'�"�'�b���O���*�M2튚M�x���!#z�����w�����?�p�i��O��'���D0{� �X�N�L:��m#`H�7M����A�ɚ����'��Z����?����-�3 ,L�X@ɀ*5��h�<O�˓�?����?���?�����)ߩ��U���^0�s���xhzUn��K�,��ǟ�	|�SǟdZ�����΃�x;�L�� Q��c5���(�)g��9$�b>���^ߦ�̓�h僧	1~�(@�!m��9͓z����ӧ�O��N>�+O�	�OrUy�D�=$�.��u	�+t���O��d�O��Ġ<�T�i�P����'��'��\���Ң�2���퟊A�Dh���k}��r��`n���ēF����7%�92:�1��jm5�'vdjca����� ��$��'�8hASȝ�WB����@���̓�'�b�']��'��>��	���
Km�N��gC���=�ɳ�M���)�?m~�"�o�q�Ӽ�A,�1��	���,@!��#���<A��ia�7�Ȧq�����-�'�FP��&��?2��������ڊW�����m�=h��'��i>�����d������3B����V8W�nux��ۋ/]�ɔ'�87�U�!�X���O��D<���O>��� �&Mf4�����Hђ�M�y}��x�^�m+��S�'
�<8� �!OK�.��!/ɱ
�<�+W�T���	�c��P'�'#~m%��'*��27%w���&��e~�dy��'+��'�R��dW���ܴJ 8J�����@ΑmL�|`C$�N��&�$KB}�f��o�M3e�
�P���^�<�Xz�J6��iߴ��DI�Qp~UI�'��O�_�DH��Ķ8��ݸFJ�wl���?����?a��?Y����O�Fu�q�Ы�p/�
߲� Y������M�����|���6�|���xc�%�"�S8ym!�NADJ�O�$a��i.t�6�(?Ap�W�6-zl��FM�s"�8��G���B�O�1O>�+O�i�O���O�����Lh:-���HB�����O&���<9b�i��s�'���' 哉v|&��̈́�a�c���[)��O�����M3��i��O�S��.Ls��A%-�D��
Ԓ:p炜(���p'?�'7R ����jn�B���^���(��"y�@����?����?)�S�'��D
֦���A�
)��1����GW�xa G-vTf���ݟ�ܴ��'.�J�V�C20��r�(0N���iȧh�86-�զaj&J��m̓�?�a��J�8�ɖU~"G�QwHK�F�{��,ñ
���y2W�����`��ԟ�I���Oo:��FI�J�"�b�Љ2p���e�QE��O����OȒ����L��睾xIDiw˚�2*�[�,U�4P�����M#B�|�����'@�#�4�y��cn��qI?��˃Nۖ�yR�����	�<��'��	韴�	*?�l��f,:v6�rP��	>cn���ş��I���'S 7�����D�O����
%�lM��1b���邞,�����OlHn��M�x���`7:P���\0�#)���y"��5�J�	�� 	�I2?!�'��D���?�ֈS��:M�v)�fm���FG�?���?9��?�����O��Ia�9�fY�C-��xY��ҷ��O6yl�`��Ea�6�'ɧy�LX�U^�,��:s뀗"�|)�'5Z6m^ۦ�2�4A�v݊�4��d�D���'%	����w�U	ReO5K=`yB��0���<ͧ�?���?����?�6!�6&�.q �%Jp�$�%c���\ۦH@x�H�Iџ�&?�ɊP2F���c�a�hQC!�q���a�Oto���M[%�x��T+�}�*8�dV!d�|�� N:V�إ�B�����^�t��g͚�Ox˓X��Lqq��/�H}���I$�Ό����?����?!��|:(O&5oP�D�	^s�A�A�Zܹ`G�]?扽�Mc�2J�>�P�iqr7mH���B��$��Yyf�ƹvX �#/��3`&�m�i~R�)|����p�'��6�K8,+�!�G
�XH�a�C��<���?����?y���?A����F�\b��*�̢@�"N����O�oڒ3(�zd���|��M�Q<(z���7�����	�>H��O��oڿ�M�' ��#ڴ��d��v*
���Я�X(���_lD�ȕ��?ё�%��<ͧ�?)���?��hѮ�. !�
����p�ئ�?�����H馥ʄAw�\��͟�Ou����"�M��t�����,0��O
��'��i% �O�S�K�Ĵb�hTҞ�P�d06���m%i�X\C�M0?ͧ_Ӱ�D� ��+,�y@�η�-yԉh��+��?����?��S�'��d�ǦI{�A�8y�� � �H(�88J��<���~����A}�Mo�@Tx�6k0h�#�E�1�<��"�Ŧ�ش+<R	q�4��dXjjl��'��S�s`�l��Ê�S��->Lɜ'��	ş �	̟8�I˟��N�4̓�K��퉑1*�Ȉ�Q�X6mi]��O��:�9O�-mz��+GC9r�
��	&���Ѷ����M+b�i� O1��sr�s���	��N�8��_�F4I��]�[�z�I�-�)���'�!'�0���t�'���� ��LѤ��d��<2��'r��'	R]���ڴa�m��?��f]����]�&�����ͫ%�%*�"�>���i�B7-�F�I1+Ŏ�x	� ��� C���2������"�_�z!*��$?��'7���	�?	$C�y�I��bφT�V䚐`͎�?���?Y���?����O��!2gFDU*��HE����S��Ov�o�2A�6�M����4�.���޵#d�C�鏭}�&<O,Uo���Mr�i�ܐE�i��D�O��ze��Ҥ-,:v��!��Ztɠq&Bt�P�D�<�-O�	�O����OL�D�O�t(�/� ;Q��@b�p3��<Q@�i&���'X�'L��a5�y��'D�A�G)Ȇnl���2y��V��/Pt�jٴ	���Z���O*�t�ҶtY�`��*���89��Ɣ�r����Ӌ�%���)w�j���L�Z�$�<�-On��@��^@��!��,��X����O�$�O��U�"�H��<9ƾi ��w�vt�'�G�,���hʞY�a�'*6��O���|�GQ�4��4Ư�Ig�Ez�"��eQ<0�H�UQ�|�rh�
WX6�c�4�	�O��t�OĢ�b��l�v��! B<#�]u�܇y4xU��?i���?����?�����?�F矪#��5;%�@<(F`@�%^K~��'�6M1,��O|oE��[W�M.|�����!܈�aI>	�4d/�v�O~���q�i����Oʴ`.ԫt%��K��%��C��K+sS�
�3!R�O��|z���?1�O�а@w�|�L��3BT(��@���?I.O��oڳv�Z��'y��O���K��]�|��c�6h�m���R�yb�'Qz����n�z�$��S�?� t�2,Ә��X ���3�Ը AeG�ªLp���'��	�?��`�'@�E%��[�H��2Ң`X�����	������	ȟ`��֟b>ŕ'�26�ϼ"���
@	�E�d��C��!w݄��������4��'�z�Q���T���o/c\|��0��,>6-Pզ�#�f�u�'��@��M�?���\$����$P�T`�����<��0O$˓�?���?���?i����I�p���K�
��.-&��m�<hmMg^��ş��	T�ş�K����pn$-szp(�Kӄ7.�dΙ=��i�~�O�O�`�
��i���Z>tY@A)a���.���+����W�I��
!��O���?!�Hi})]�f	���M;��,���X�	��x��]y"Mt� ��6O��d�O�0���>E��%� p�(�`,�	����ڦ}��4{�'���G�_جq١H�<<�t}9�O�YC�C�8:it肢�iߟ|Q��'���y(�8#~!�1	@zV��86�'���'�2�'��>��I�ch�1
rN�S�>����ܕZ��e�ɲ�M����?�� ʛ��4�l���_X̚� ?F14��23O��l3�M�ҿi��ɪӽiq�I�~0b���OJxX�w]>"xĀkC
��$��2��E��Uy�O�b�'C��'�	D� z(�
�E1j���]�w��	1�MK��>�?I��?1L~B��t.��&I*wD��r�	9�JU��W���4[���`4���N�@[���U�mª�A���9=6@����V�	$8�z 2 �'�0�&��'��-��MH�l��+
��5^�t�I���i>m�'�6�S�V���d~���j@�l>ru�B̘=�����M�?�W[�d��4ab��b�R)D��5�L%
bI�"��Z)P3��6m4?���V�[K��/��߁��nǟ0lp%I�mB^F��r����֟��ԟ��I۟x��概�}@�L�A۶"��8DЦ�?���?i��i�:%�̟plZ@�	�7�5��G}���KtĊ�GU2��H<	��i7=�n9�%gv�(�T鋀��=2�<�1�*L��g �>���#�䓇�4����O6�ē�u�^c��Y�9p��"
��t��d�O��
䛖g(L���'mrU>�R��,n�L�s�!R�:}�g&?1"W���ߴcțF�;�?�"��/&:I���p{�Yp�FW�!����e�S�N����|�c��O�՛H>��9v�8 �A7���2�[��?����?���?�|R(O$�m��_c 18sgL�TW��J@%T��|��#�CyR�`Ӯ��J(O��$�1h�%S��B��d�'���f6 ��]k�`Pܦ��'�IQeg��?M����0`�7�1kPEڲI�\��3O*˓�?����?!���?����	�U�-�ըŮK|��`S��XHn�n!�	ßH��Z�s�8������k��tNR�fm�k9�I҃���Ҵiɮ�O�O���i��Ę)y>x� t��*��4 C�Մ%�d�h������5�\�O���|���a�vXq�� 3����CdX�)� ���?	���?�(O6(lZY���	ş4�Ɍ�,@�E�?���s�HO�|H���?�F_��K۴j~���1�M� ?���$v��!�R�F���9Hz��ڱ����c>}�1�'����ɫ6I��آ 
<D���Q@��`����	ߟ���؟��Iz�O��M]�#fnH�DOA=2jY(�bCx���`Әp0S��$:�4���y�jl�|�Gw}�X
Ã�y҄gӂ�l���M�Ä��M��O�L���Q����-�.~���E��p��J� �O���|���?!��?��ux��`1��'BM��k҆P-}B�J-O��mZ�Y�h��I럀��c��̚���2�Z}Y��K"���3�K�9���O�1�4���OOl!bv��!X3hT�2�߳ Rm)"�X.
3:I��O�:W$ձ�?1�O&���<A��ǧT�qP��ӣLD����W5�?����?9���?ͧ��d�ߦ��V������$yK��@�ᑆ�O"t�����Mۉ�I�>�Ǻii6mX���٥�\�[�rh9��ςF�	�H�����n]~b�SYktI�|�'��;��by&x
VbJ�J5H #Q�<)��?���?��?!���kQ�cZe���
���J �
)k���'F2/i��,zw=�>����'�C����mtB]H��Z(��������t���w��)�3j��7*?���"�,Kbk�^0R���h�i�2
�O>��O>�*O�	�O(���O��7�ʓ,�|�Hv�ιg"�� �c�O4��<�U�i+H���'���'��j_z%i0G�:*U!"a@�e�P�x�I��M�f�iMO�0TަL�3�M+�l�i1�
�*C%f�DT�h1qj/?ͧ>���d֞��"����C�E� -�%�2E�? �<7�'?�'Mr���O�I �M#U(S+/+���N�	�-#�!\b[�����?	b�i-�O(l�'�6�����i����n=�M���%.w�	oZ�M�'��M��O����@ޕ�"H?	�gMMɒr�W�-��O?u���<A��?��?���?�*��Q�g.p&u�6�%5]2`��զM)��A� �Iş &?%�	��Mϻ	�*��Ӄ��R�1�A��>n4�&�i�~6-g�)���eo�<Qs�� ^ �0c�
��M*h̔�<��3z���$������4���$S�'�$�X�'	x����ݕH�r�d�O����O�˓{��H7�y��'�"j����(�>~�Bezc#H&H��O�0�'?�6���1M<� @��^�ty*�OB�-j��@�����X��<y1!1�ӏX��!��B�D�d~���^_An-�W%N��x��Ɵ������F���'�� Bs��8yt��ᦝ�[x�8���'{l6�Z:�I$�M���w�̭���H�h�ԫ]L*fc�'�7�Cͦ�b�4wp�ڴ��$���J�'�$!{���3�2y�&Eѥ6|	rn2���<�'�?1��?���?�c�'*��q*�o
�P�����(�9��$�ubWmm���Iן�$?牟z*�8rNJ����sȗ�S8ڬ��OZ�lZ<�M�f�x�����@��N8�1��1^HV��P����JI�¨z��r�O��Y,F���`Z?F�r�8���z�,1��?����?���|*O�}o�"���I�7��z̱7`$@CSF�H�I;�M[���>I�i7m�ʦ����3O���+ާ� U!W�1?d��l�R~2�\[�t�����O��ʀ40���V*b���(��Γ�?����?)��?����O�䠈&R�;.LS�KI�Om�	��'e"�'��6�H����O�l�~�I�M�� ɓ/��+�i��\@*u�L<��i<t7=�J4ʤo��.���IS�ǱK+*�����+��eh�P69�l�$���䓻�4�f���O����t�f�A-Z9n��q��O�)�j�D�O6��V"�(E���'��W>��Q. @�����8T��Yp2f)?y�S��z�4*?�F 0�?�I$�
 (f`	�.�C��A����D.�}��©0����|: �O��H>��(�@%S�h��v�޼���S
�?q��?����?�|Z.O�m�*^����UǁWS���'�B(f�LP��>?��i��OZ��'�V7�
K |ܓbm��)Ӗ�1vɥ�>�lZ�MS&��e}���'2���m��?%���� ��L�v ���ؿC
`���4OV��?���?A���?9����d��UFT��!!T/Y;um��7*����� ��p�s�p�������}ˎ�)��4T�~*�-���i>�O�O2��F([��y��DK��٥LW5�t��Ë��y�aL
]�vu�	8?9�'��i>%�I*�����i�z"��t�7T�D��I�x����'�L7�θO���O���99��5�w&[�R���Y<�����$�V}�i�r0m��ēzt��Ќ55\��i�)�/{(�<�'m�,ړ�P,[�R@��$�P�|��'��2F(FND�]�.�`_R����'�b�'��W�"|r�\R��&��>4JhJ/�9��N �/@����IԦe�?ͻw ��0w)�5��)�(�&�X��?y�4w�����"=�h+�O�5��º���"ȫx�"��u�[=
gN���.�OB��|���?���?��*a���ۥZ���)�� 8���+O�}o#CJ��ݟ���m�s�@�r����,��^Z�e�@�L���O|7M�D�)�	��i��P��2֐�ЅkK`<zЙ�f���	�,�zT���'0'�@�'�<U�1d�>����˗��Z��'�'F��'�����TW� cܴ,�������aj�؜"̱���{m��K�zݛ��$t}b'g�n�mZ��MS��A#dB�b�	WkZHU�D�`k&!�~Ҫ��R�Smܧ׿c7�Dh@��ʴNث&RjT*1���<���?���?���?	��4k�0h#N�OґPs��1ck�b�"�'�|�L�R�?��ܴ��K8X�ru!^0���C��>�$���x�fs�\Dnz>!ÖI��crh�I8 ���B�:N��d��N�/�0��W�A3D*$�dL�����4�����Ox�DL�[d`q�ɍ?E�D�#�)���d�O��u��Ɓ�����O{�̺���96*�����>>Q8��O�`�'�:6m[Ѧ�HI<�O������K���V#6��(H&�O�(2K��P���4�d`B��^�h�O�t�Íe���wŃ=@L�kRO�o�7����������d	�
-
Mð@˟h����MS�2F�>���i�p���hCV�R�B\�/�Vx��dj��l�$`Ĵ�J"?Y7`K40�f������R�(�㉃�#h���S$R�$h��<	ߓ�p�Ip-�&z|*����@	��i�B�t�'���'/�@lz�����5|�Ѹ5n�8Q��ɻ�����M���i6hO1��P{si�-\���^ي &c�o����R�D_4�d0e3Ѱ�+�֒O ���K	01��q�� jx�y�P��;�ax�i���ђ'�O|��Oh5�a�O�D��Q�q�L�cMt����7�ɻ�����ݲ޴2��'�i�s��g¢9��_��e`�O�E3R��0��1�?�iʱ�?���Ofy9�/J�\o>��Ӧ	(��C$"O��CL��4���>#��LzR��O8�l��f�^1�	ԟ���4���y�
T���Xz��߫G4LzG���yr�n�R�o���M��OT�R�)�'0J<rwFZ�?	:���d�:����?$D�bgl��5�'"�	͟@�����	����ɨ(����)�+Tڈ�:��7w��'�47�6���Ol�D5�9O�`��ޜNēkR�p�8`�3�Au}"h~�&�lڅ��S�'hH@I�ل�D��d])m#�����_�y�'�F$�%�ߟ4�|BW�0r�i�w���g+Q(S�zu�0.埈��ğ��	ݟ�Ryҏr� ��3O��@qc�U�Dݓ�� �g�4��8O%nZh�m��ɡ�M�i�T6� ���`)֊r3|lcUD@�h��J�g��:�x�(痟*Ջ���i����Bd���_kt��(U��H56O��$�O����O����OF�?�s�H]�p��2���-R�b��3�k������4Il�q�'�7m>�$Z�~�X�CTC$=���@a�<3��%��	����7LhEң��X���� M�x�D�q�V���9m�6,P�'��4$�4���4�'���'��R��=�	�ֽz4� S�'�R�Aݴbb|�ϓ�?�����)��C`��d`�t؄𣜰F������T𦥫޴]㉧��Ws<t��lڗB���GB �p����U�f�y���!����y�-\��b�T�Q����"Dur8����`�	���)�Siy�nc��#!޶-���v�@28���ܺ+�	�Mˈ� �>!��i\dQC�k�5?t�(��������M���i~��٣�����D��AF�(�����"!� "ԠW8B���C�Ҥ~�0�cyB�'���'���'��[>-�À1rb�憎d�5�Q�ӓ�MsE'��<���?yH~�:��w���dGر W)+�O��$�@!��p�lo���S�'nV��
��<YQ���lz�a2H�^��I�b�<�W�V���������4�f��ٔpD���Xw����o%?�����O����OJ�@�6fE��yB�'��,�vk`]��o��o|���a� �[��O�)�'�d7�OȦݩJ<i��I���n�0�bhs��x~�Oݵa�Ua�%�טO*�u�ɵW�B�?;�L�N�?]^�� �]�X22�'��'v��Sٟ$I�H��BL�D� �J�3.�;�Sџ��ݴx�Ty���?�@�i��O�.R	�rY	�+Ĩ+B1�"�5�$�Ԧ;�4�?asAA$d�'��(P��W�?iPT�ȼR/᩵Lژ-P�9eK$��'�i>������	ޟ��I�#���C@Cy�4�&B-6��'-h7��)�ʓ�?	K~���[6��R$�^n�Ph�v�l�`��S��ߴ:C��=Op"}2%�¼D�:T2q�-u˴�@�B>j@p��t�v~���6|���Il'�'�剂A.U�ȚO�b�("%�[��I�I韈�	۟��i>1�'(�6m�A���֍&�Yؔ,�#J..xY��_	d8n�d�Ʀ��?qdQ���ڴ&��'X��P�� ������NC�0��yʕɗ�/.���O\œ�K͖����k��ǏN�k~����-�MX�p��du�P�Iߟl�����П���(]�iq�9tO�.X�1��!�%����O�l�u,���X��4��$�T����8�uJ��G�r�':�I��M�����N0>r0��O�H2���%q�J�J����LU&߿R��(�� ��O���|���?Q�wN(�6�-^b��%��J�%9��?�,O��m�)^�0�'n�R>�x�HF&P�L��KV�(�r��)?1`W�tX�4Lj��9O�b?�i�@��FذI^'$�h2Aɚf�6j�/��~��|����O6��L>Q�\G�؋)N���T��DP:�?!���?����?�|�+O�m6M�.%��J�'$p�$�p�<v��Bs���x�	��MӏR��>�жi)��wo�#yK
e �X��l���j���dϻ9^��@���[!d^A��ԓ~*��N�15fᲷ��2=� ��uf��<+O��D�O^���O����O>�'P;�M���&��'Ů	�����M��hI&��D�OF��t�d
���5Z�� f�=A|�KB���ѸݴgÛ�7O��S�'߸%*���<�@�Y2�bb��U4ҵ����<a`��?*�$X�����4�����3J���C`�� b�c��P(_�����OR�$�O^�p^���� k�	��H1�Fњ_q	p�B��$��Y�T��T��!���*�Mְi��$�>���R�x��L�2��0/T�2!�Jp~�e�aN���cXƘOz��IF�/��e)�1��n�_.x;3d��?���'���'��S����j=�D��EJ�3+bBUNݟ�@ڴb�n,�')*6$�i�)�c��<>����b�C�8E��,n����4���p�8�e&�K����C�:��C�O��UzU.�1����J�f���e�	]y�O-"�'(�'�Dˁm��+��/zl��X���1u�:�M#p%��<���?yM~Γn�4�j�)<}�")1C�D��At[�h8ܴb2�&�;���9��0��n�2R5�-�`L�o�<_$�4�e��ܘ�y��˔V�Wy���@th�G�I ������ѹ?���'A��'��O/�	&�M˗���<A��5N^���C��Q��0����<6�ix�O*y�'�X7-����ٴA����J�f���(T�L��p�0!PM�'�h��' H�?��}J��}��i���+���Ъ˝`̎͓�?����?����?q����O�B�uGH��a䀍2
� �O����צ����(?qd�iJ�'T(���B�Y�8 C��'@vp4`%�$J֦����|:�m�#C$�'Tx����sk���M՚W!�H��ȏ7u�Y�	2z��'t�i>��	��I�<�$��� ݩ@�&��pHI\3��������'7m�"e��˓�?*�DY�3 '+�d�R'ׅraP��4���ٯO�m���M3�'�����ƈP$��Qb��(^�0�H@��\)�!l�i>ur��'
�H&�4X7�ӵ&�ƨHS�	�O��Zc��Ɵ�Iϟ��	��b>ɗ'I�7�&9¶T�s�Y+�l��#Ϭr���y2,�O������?��Z��i�t�? ��6)��@%R��E10'�S�JΦ��ɲ?��(F-?y��	�M�n�	)�d@��!�И����"��
�y_�0�	��H����|����x�O�������?k�@��5X̤�U��M{T$�����O�������̦�]�Y���Ig��AeBEb$�;z|���4r�F3O�S�'?@FPV���<Q'f��\=�2��M�$}�o��<��O�5��D׷����4�z����LP��;��4��a�1��\����OP���Oh�pɛ��ڹs�R�'G"��2W��i��:�����"'�>�G�is�7�Lr�	"!�>8��IV�H�1s͂5	���c�T%�F�
zj� N~���Ot�H�H�e;��	�LZ*Q��Mp9�����?Q��?���h�&���*���@ş6r��I��G��$�D�yj������ɒ�Ms��w��Y�7 �'�����;�^:�'��6���u��4
t��Ϛl~��;�V �S�X��h�X�x|�3CO�5�h,�&�|rS�������	ٟ�	ğzd��

��9�p,� !Ӥ@9�Lry��d�4��2e�O����O����$�9U|�Hd���i\ؙ���UJh��'�@7�ɦ�J<�|"զ�%�, [�H���Ъ�oU!%�ȑs�.C���d�Q���k����O��-$h��Hֻ7���tE&�<���?!���?���|"/O�mZT�e�	.?ft���-D8�!ËR0#/��	��M���<1��Mӕ�i��Hy�)��&gx�te�@�����嗺O� I �O�]g)����d%�i���!R�Ȥ�А����k�f���7O����O����OB�d�OH�?ii���<��HI�vi�p!��Vy2�'��7��%3l��O��lZg�5� �R��5&a΀BjD"Z���͓�� Ѧ����|B�M�xM¨�'rր�oD9s�M���Z(���K�$�N��ɞ��'��i>A�I��T��,;�I�N�9�:l� ����I�l�'<6M�*�˓�?q*������^6�:�AA\�������8�O��l��M�'���
���#�2k�		s樻B�A	w����ˇ�%��i>U��'c�)'��M_�fy����gٴH���$�I�����ҟb>Ֆ'��6�K�]�pPK�̝#���Y���.l!x\ޱ�$�OF�m�N�{n��r����Ɔ��w�`4)����M���Vy:e�A_~��a��u�H�)���(r�D�%���Ҡ�ݾ���<����?a��?I���?-��aJ
;>����jG���ȕʦɐ�DAGy��'��O�Ra����R���R�`ͩ�6Y��C!5x@dnڋ�Mk�'�)�Ӎ{��*��f��u֣T�-����pl��m�JE�>+���V�I~y�O�l�]�HU�E�G0��рO�>���'��'��	.�M�!�#���O�@CR�*U~�{G���̀�K.�	���J��p�4�y�S�\�p,դ(X�ݫ�%��0%|hb��=?�WA��y�� ^ḩw|�Yv'T6pfdu3&"Q�;��q`P��N� ��>uJU��
�&�ࠇ�6mV\�!V�/ք� ���8 |����(Af���� T�q������O����e��&>"�b��ܲ,q�Q��(UԺq�|�W#UU��)�M�v�IQ!b�eK- +$������xł+V�Ou��s���?xQ��
T+v�J�[�@;s��Y@��6��@�L �vi�Ðké?^�}�eR�l��V%>�^LZ"��&J�a�eN�bA���NH�	 �C�c�d��EԠ{�B]kD
L�i�HE�i��L;kuNO����O̒Ok��m�*(�'	O�K�����׷���'t˞'Y�	㟀���`��ʟlA��hPYZ�ǜ�F�x��+�9l��'���'mҖ|��'lb��?���ٍ6T� $hȮOK�Ja�(!2n��?A���?����?�QÀ��?%d�*8,�s�a�;,o Mӂ	ϭsћ�'K��'J�'J��'D8�����M��d��s3LP�4V�3`ȸi'Gt}�'���'8"�'�|U"[>���5E���h�M�pt�Ү��yߴ�?�L>q��?���$�%���f�M_H\��ǎ��Q')x��D�O����O��م��O��$�O.����L��u$�!�&Tp���v>�+��i�I��$�ɘ֢��!�~JDf�.VƘ@#�߾N�*��t�E�	��؟��m�����qy��O��i�q�B�[ ��hh��6��qӊ�D�ON��V�|�1O���L���'��$a�]o���ij�l���'���'@��O-2�'��Ӻl~f�[��
 ���=B#���ܴ�:%ȴ.�{�S�OCBmU00f�`�RO*�iO\%e�"7��O@�d�Or�P�l�d��?Q�'����ƃ�!5P���B@�%ڔ̀�}�ǁ�Ԙ'F��'"�"c&8(�Ɣ8Ga�H�U	X7M�OZݹ�(X}RQ����b�i�Q!�GƲػ���/�
|��>�%��/���?���?�,Ox,굊�4?JV S��ݿ~p�c��(t��D�'��˟�%����˟@����^{@I{��X$Ew�a��� Fh��%���	џT��ty��A��)��B\�	0�]�O8k���}n��'��'M�'��'���[��Oj�2��N�&�ꗮ��7!��z�V���	�����Sy�̀1P��'�?	2N��H�7��.��E	�J�9`N���'��'���'��ycF�'!�Bp���X	Ir )f�x��@�Ц)�	���'�$A���~*���?��'h��R���p�J5Y��$;��i���x��'w�d�KU�O��������d��n�#�kU�
�|6�<� �W97����'���'��dj�>�q�? \I�h�$H��	��L�W����$�i��'��Л���7����hց�%[l��4@�no�7m[�G��}lZݟ��۟l����D�<ф�F�lbY��7��i�����RÛƯ��s��O��?U���?"L\����"Lh�A�ִ��4�?y��?ivm��R���Ry��'����j�`)�fbK14�Nus��^�#��O4$K$)(��O|���O����Ɵ5������a̺�*�A�ߦ��Ʉ:%B�J�O���?�L>�1O̘�!<ܬp)s��*U���'U�Az�yB�'gR�'-�	qBBԛu���ZE��/�|:�KvD����<���䓟?���Z���R���o(�}���&�ڜзK�4���?��?�.O���aB�|���^��x�_�k��8r��͗'B�|b�'~r쒘��	Jm�TAR���F�� j4�US��	ޟD������'(!�S��~��Jm���$҂}ڜ=! �ߡ'�xqe�i:��|��';�؇'�>F�Y�u�©X���������צ�I����'U�*aB>��O����F<��B�8��Y�[ N��̙��x�]���I�p%?�i���M��}0t	K����i!����EӲ˓hPHㄼiC��'�?I�':��I�?BUj7cұ�`šԭZ���7ͧ<����?�����ܴ;ܨ��4(S*En�Ԁ:Nn�o���Pݴ�?���?��'n����dM�;�Rh���u�h�q �"_��7-�O���O�O�s�L���� !��� 5ڴ�Y�e�=���"�4�?����?qC�޷)牧���'P����H@��
Tpr����(���'I�I#@�<�(���I�p��c�~��sl�U�HA�n��9��ao�꟬���
Ty2�~R��K��2���c��L��!;��O͜�9s� ���v��?�)O�����D��щ�:f=z�0ŀש?�N̂ao�<9��?1�R�'g�cԤB��܃�D8eJ�B�&�?"0n�b�����'hBR�h�	/'؊���x�`0�*�Iʲ�Q`��[�<Un�ʟ$�	f��?����8)�����! 1��H}vAZ�eK7 d�H���>����?	����{Jna%>�q�Lѩo�����N�)�hU1!�1�M;������$Q�{C
��/��f��@���)D�{��h��Mc��?A(O0IR�`YN�ɟ �s�as��Z�~���3!�"*p��k{Ӻ��?Y�"������'��1��ys��]��5���ׂ{W��d�<���Z�&U>����?�[�O�L3С�&	���N�5�n4���i剁&aT��&�ħ���ݺ���n�H��K�)x֍x�!c�~�I���O�D�O����S����m��\3E��?Q�@���͸M�,6-Y2��l������"SC܂x���J�2=>\�Ƌ]��M����?Q�����b�x�OO"�O�Ղ5bO�<6�93��> yq�i��W���w%����9O��D�O��$��XA�fn 
��S�%"�oZ�l�'����|�����Ӻ[q圼	 �*��
�m���sr��n}��J(s{�U���	��IWy�ÄB�tM�B��^�@�a�7c
�(�"7�$�OD��O*��?�М!��Ν�d�����-=�v���/�+�?�)O���O˓�?A��C���d�(j���H�f�1`Z\]	�lԻ�M����?9���'���D0�@ܴrjn ����$�0�r#�4b��i'�x�Iryb�'��y�Y>���$�,��ci�H"X,N�.�>�a޴��'fb�'*�aA�����[~�`�eF�/~�P5��@[p�Xo�ݟt�Ijy�K �?�����$�kl��s��z7@�R
��ucT��'���!R�n-�	q�SGj`d,n�X@�@8ѣ�ZR}��'4��x��'��'PB�Oj�i�=�!�/~b��㯊7�Y��@fӆ���O��i هT�1O���A#j�}	j^�9�R�pָi�j�aTBu���D�O���⟚�&���00�S�L�!>����P��гܴZ��|K��?�*O����I?U^~� 5�� `��pqm�Q!l��4�?���?y������?9�O< @���0.p�C�D
���(�#\~̓0�����O��	:_:<��n	�\�.H�Wm�h7m�O�9���<YE[?��?����1O`q�E��^�! �/X�L��	�lr���>?��?I����dצ0i�ŒBF��T��l	�O\?K�9���l���� ��C�xy�n
�/*֌�Ɓ��M]j�Xen�aL� �b�'7�	����ҟؔ'>�DF�k>�H�X�B0��2��+yY@��>����?�H>�)O4� 0E�O�S���&*Yh�Y���=T�e�@[M}R�'B�'��	;Q-���O|r�	ڪv:5�.�%�~��Q��*11���'��'c�I�2�4���D�I	�5��A!A��@|kq&>oЛ��'~�Q� ���=�ħ�?���a��!X�@Q�o�a]&DtDp�hyB�?�Ҙ��ٟ��y%e�+/�2䙵K�T����i�剚7��l�ܴ0���ן��Ӭ��䀚~)��ׯΌ1�H��jW���Ɵ��QfO�Ot|&>�%?7�$i1"y2��7�����	�	���CʲO�7M�O��D�O�i�b}bU����o�\���+���;�����_��M�$J�<�+O.��"����e���R��m�Oǵ6�|�#F�0�M����?���wp��R�l�'���O� ���B��B)H��@G�~��S�iXBX��K��}���?����?�BA�>@����^'|�T�B�
F9��'M6����>�)OX�d�<���kR��)��Z2oڷO�
�!%UO}R�����OJ�d�O0���<9�%D�{�|᥌]z���'-ɰ5x�]�Ԕ'i�Q������8k^����j\bQ�"�	�AC�|��e���I՟(������Ly�L�.)wn�S2��8e�O�X�1c'�)��7�<1����$�O���O��72O�)�B,���Bc��
!j��4!����ПP������'��ɸD�~B��`(٘v��(:��+B�D��9`Ӻi�2T�$�I۟��I�u\�c���*W4�@v��f��{�I�����'��\�FD������O���|!����;Y�\��e���L��I�@}��'�r�'�Ұ��'��'��^�>�^�`r��L��2c��h�i|�I�a�2��4�?����?	��!c�i�1��\�v<EPl�LyƕP�~Ӕ���Oޝr�?OZ���y"�	�g	�R 
3$�J�:�/ˤ]�vBM+Q�6��O��D�O.��G@}rT��K�c�7z���wH�#nP9����M��Z�<�K>����'���x!.�RPv����Hc�@2'd�N�d�O:�dW�4���'P���h�2Y�$�k�1�YY§�5E�H}l�ݟ�'1Ș˜��	�O�D�?�h����z�<�1b�3CN�4	Fe����6���'j�	ß �'kZc���O˻%����T�'��,b�O���$=O��$�O&�D�O��$�<��l�m �u���.��tSp)ˤn�$�1R�X�'�S�\������=��Qp�F<|,�̑G��+@��P!��q���IܟP�	ڟL��yb!�
2���{���1>Ȱ%0碔5�t�ٴ���Ob��?����?I���<�w@?
zZ��(8ထ���׬w!���'��'<�^��Kq,&����O�(�Ө	7ZJBT�V �5)жj[<�6��Od��?Q���?q�.Z�<�J�Dʃ��[�T)�,ؖQ���s�~�"��O�˓b���Q]?)�	�t�6k0��k�j�91������*B�zD�O���OT���/f�D�OD������kCt�8AFè'��cjQ��M�+O�<���m̟���ϟ��ӣ����4M�.��80��͓1�j��q�iT"�'T��'<���<���$���v@p���a�x�9-O��M�HC.%���'kB�'3�$��>+O��k�&A�:��hʅ�N��A-oܛvn� �yR�|����O�DRdNW����c)zK��-��޴�?����?ѥ��&��Idy��'^�ğb�����/��k��Ŏ#ǱO����$�O���O�i�ׯ�w���w�8C�l��%�զ��I3H�� �O���?)O���Ƥ���8 >� #�MA�P��Z����>?���?i��?-O�����ū�B�ãǖ�W��B҆,EY���'��Iן�'���'\2�ϊY�Ń��5��T3%�#�4��'4�	֟d����Ԕ'��Y8� s>�' SD%� ��/'� ����p�ʓ�?�-O���O`���s��A&1���s�ӓ<�)���P�R�m�㟘�Iߟ(�	Jy�ňz���'�?y4"��8E�7h]]�E
�bL����'��	��d��۟���f���f?�҆2Ml$ b�t�:�Ĩ��M��Ɵȕ'��5`C`�~���?��'~�t��7�L�G�t|�r�D�z0kQ\�8��֟ ���|3,��ĥ?��a�b*�8AT�����p��mxӎ�FV�hX��i���'+��OӶ�Ӻc�dF*P��E�!���`�������Hp*d�D'���}�w×5�H�����)��7����c� �M����?I����7W�L�' ��i��)%��%o����7�p�t��>O�O��?)��*2(�R��Ũ3�K6%��M2���4�?Y��?х��Gz��hy��'��I�(�Z�S���&��Q*� ��IQ��'���*u]�)����?��OK����ń�|����h��p��ڴ�?1��J(���syr�'C��֘���� U�U�O�.�E��Γ�?���?����?.O~����?5�44�C�]*5���i��W@���'��ڟ��'���'kҠ��07VUcb��+�P�Ӓ��
T'#�	ǟD�Iɟ��O)���0����2�q(�*�Xi�q�xB�'�'7R�'ih���'#t������3� n��ّ��>q��?i����dAt6$>u���3O�1�����l��D��M����䓾?���C*D+���I,[ԕsO�Ie0�
aI.M&�7-�O����<AhA�Y�Og2�OK�E9���{||8��J�
0~�@m%�D�Ob�D�',Mr��/���?ͣRO�9_����썁hKP���mb��˓f @[��i�&��?i��9(�Ɇ;:���H�*$@���Or�6m�O��	�6��5��$�	;���1gR�MCP�KA�U6��1�xAnZ��	՟�����'������@��<Ǩ[�ʐ�r������O�O<�?�	  �ʕ!��:򎝂�	��8p�4�?i��?�ӥQ{��O*�伟(�%ˉN�P��W��4Ug�@�6�c�`�O�ݚM�G��ğ��Iʟ�rBC������ɞTn`p�����M���3���s��x��'�|Zc�2E���8��u�B�>	h��O�8���ORʓ�?���?A)Obd��$4C�k���{;�p� �D�IbL�>9��䓮?1��b�� ��C�Ɋ&4�¸+#�Y	T��4k�<q+O(���O���<�c��:��i�m�މX��)_�pz�h����|��O���x�I(i�@�	�e�8{A$Z�Xh��7�Щ����O��D�O��<�w�I�#��O�^ ��!oM�LU-.,�rb,f����+���O����-$����#}�@�PȌ�C@M<f,�T�0g���M;���?�/O�t�2�h�埔��P�NL�RL"`�&�"'�X?�8H<���?A���<iL>	�O�mPu���j��0�%B�L2���4�?Y�������?�(O��)�<���.�Jw��_ш[��R:8�o�ş4�	=r���h��8�)�CДs�T��hE� �T	"�72J�z�n���(��ȟ��S��$�|��89�n��T�#���d���sԛ��43U�O��i*���O�Ȃť:��m��`��
�hqC��������I9N`l@�'��� �v�d�#�JÜP�8�����c�2)����K����&>M�I<�ɬ|�0E��ɒe��{�� 7�P�4�?�����?�o�����'�@����j��t��N�J�P�EJֳ��DԊ61O@���OJ���<YCD)�������N�q�Jр6ײ���x��'�'��	�4�I�G�br�	:������"#H�I��b<�I��(�Iry��'z��Q��d@��	��NB���m٬FY��B�i��ş�&�p�'���+u�I��Ms��
4]u4q:3�Z8+�A�l�~}�'�BY�X��Id�~�MY=y�:�	�	#B�1��ǃ�M������׻o���5�x�jE�$c�,O�$&X����į�M�������O(��R�?������j���2%���HF1[�G̥�I<i.O�sӇK�K1O�STݪj��#x�V��cɴ6��O��D	�<;J���O������?��:�n%�P�Y����QAW�f��Um��4�ɾ4,�"<!��/�'�mb��?]���P���	�M�An7�?Y��?y����,OP�'Q����.m�ժ�8q��ictl���?�Sݟ؂Ǎ)
F<T�õ#�j�gù�M����?��h�h�.O�ܟ�3z�8�u�^���I�&g̙`~dm�T�$\To��%?�9�@SnpH��i[.��w�
���<Q�l�#Rpe:
�'�Zx�ա�$+ �}@c�[����:דU�T��n (m��1ɗ��TXni���TXf�!ѩMO(0 �c��p<$������Q�  tV�h��Č�`0�`R���t8Db�P�:��d�V�]'C-����`F)�re�iJx��d�
�f^�"a�U�[` �I�0sLD˕�J8(,��l�q������&n��Y�	����c����,���|z��U�h����l�:Y��a�a@Ly��=����ㄈH��?������	�Y�i$���>I!�͉>����@F��<B��)��i�&#�>dԉ�N �9Rޕ���D�'���؅���!J�ѩ=����yr�'� ��b	��O��XK�52�z���'�6Mȥ����tEQ-a3j���$�0��D�<)�I��"���֟�O�Y�&�'�q�n/2c�|��x�Z�'�2g<%�d�FK�A������O�@��d&1J0�!�(Є[�8�ر��I4>kd� 柨s�X�����_�O׈aP$��;W� "g�����T�J��YD��Oz��<�'�?��`H�+� �-�cwɂ�}���ȓh��R�.�%4B�( �ױ%w ���I��HO��H'$�<i,���+*J��	{dDIk}�'>�B_�`Q��'��'9�w�"ȣdL��0�4�a�B�m0�1�莴l�x�C��O�hx�e���1��'�Bm"���0��H�)vΊH6�خd(}��E�O��tJE�����LR�!�&�E0Y �'��|g�S�����-��O�ў�R�/YD9����-L����8D��L��?�\��)��{P��g�;?y��)�-O� ��.е��(Jq*3L9�P�JQe��(����O��O4���պc���?A�O%Jik����Db�"z�L���Dې�x2'ʜ�]i���g���*�f�!A9�]Ru"�3j:����15��#�!�=bFa{���;���M�m�:�c��U^2�����?y��$=��%NNz=*@+�	L���X(_��@B�I�a�JMK�lM0���Ѧ�]$0�c�h*�O@�	>z�TZ��	6xݢqZF� LY�E���a��M�	㟠)@�������|ڴaT 5�ܹ��G^V��u��4r������u��c�&�)�H���0l�#Un���+#M�)�� ��#��=�4��4\�DQ��+O��
��'�bR����I<H�@�23��M�+,��b�4�Z@��n�.b����)�_xB�I�M�`�W(+6�$C&G��)L$)����<y����_�*�y3#�7Gg���*�I�&B��8���A��-�rHS��f�C�I-��x
C��%K�f:��L���C�
`7~�;��GL:��A�)�!�� *�CQ��?_�H��c��l�$"O�(iVi\hX��K�$�2��"O&�)vk�"��l���&"���(s"O�����[��a��d�Ҥ�ʕ"O>tKFh_X�𴣵�J&4-ۃ"O\]�P#Y�4�N�H@�� �rh�"O� i�dϭ.�,�(�X0��(��"O�pX�N�(��Ȳ�Ş�P� A�"O�`���Lޘ`��]'e�4�H"O�@�Bb�j��XtI��8�|5Y�"O:]C��m�����e�(|R"O�P��50�s^�� $@1"O���f�R�5�>��C悲X	r�j"OF�c�k�Z��P���+h�i2"O"�ⵆ1h�
r3��L��KE"O`t�ԌJ93�ԓ�팚#LE�"OT�!�i�-0��)�W
�+_��"O8�0�l �J1����S�"O0[#�X%4�^�!����1E�hs"Ot-�K�:Y�4�kc�U�fX�"O��w��14���ztF+_(��G"OT�`���U������U�9@�%��"O.e�0�2Ρ��C��\��Ĉ�"O��p�#F1��Al�I�HX�e"O�0�ۈ�Z\9R���*B��ʄ"O�`P4#S�hV­��OC�M��].�y�
�8x`��/Mv˶jքX7�yr�J�a~B���Xm5�<��l�-�y҆\�(�B8%HY��Xǁ\�yrH\�E`|y��2�����J�y"��Y=X�g+���Q!f����yb�Jj:t���U���]��y�	�lm�-c&�ڧI��T �-��y�˓2Yf���E���q��y�)Y�td�@�Q��=-��{��V<�y���9D��Q�%���\���	Q��y��ޤz�u` 䊀r�DKp���y2���~��T�%j˞��T#��y��I�l��Պ�Z��1o=�yB(^v�z<�sG
�t.}�U`9�y"�۸F��IE���(�r�el��y��A�~��s�J�/(��tB5���y戅�<�sB�,�<�T���y"���>����f�r�����p<����&�qO���t���"���+�%}g4H�B"O�-)$˝;�&ip2kW+~ZP ��^����ٌ-�b��|�䫝vgF�j����t��<�@�Ju�<1�kY�-ತ�l F$E�q�dY/FY@�J"� N8��#fȿR�����ń�HR�7�O���q��`�9�LbH�3PH�KT�є��'(ڄ�0?A$�¢? ����nOX޹	���x�'cȠ�� ;�:����7����O�Q[��1q3rڦ�L�
�f�'n-4���d�.Z؁�0J�	y��h@W
�O9⦍8O#t���&�&4%���g}����o}5C�i��o�*���I4� ���@��X Q�+>?�y
Sʛ�SZ1 �%Reʰ�'JN8j�P?7��/%�J��
t��F��r㯁�(�b4���=�O2�j-͛nX��oъs�fx�Ul�]�>��Jڼj{�:�g��?ّ�C{.�����R^���ME�HMiԮ��OQ�L[��	��^���E6XHLkЦ��S"ku!��%�f)�Ӎ#)50$�
�'B��ЗM;d�� �\0e��X !��)=Y��A��Q�Nr�Q�e�%P����#&́�&3��Dg���
'ʓk�`4c��S ź�;2�Z�J��D��
'l���V��Y�	X"@��c�����&^$
*�%b�(�V"'*�m+�&���|�Z�� o-�c�b>�K!�T_;��ç@K���3S���77�����CŴ�85FPs�zw+�H��:P��� @��7��p��h�J�v1��p��O֠+w%Fq}��	P��̱�M�k�����M,���#��yHV�V�M��y %�>��8��捅`�x嚌��*E5���}�0���O�H,�Fj�1?��m�0f�r 0�a �\H�2��זw���OX�p&�ƴ�ywɕ��.i2���d��fR�b�b�<i�/�'S2Q?a� �=jLl���n7��&Y�@ܡJ>���	P�3[��kC�˭F�r��w����艀G�m�V$ X��N��(�>�~r�I�%����C�Dԫ�J�2W�b%t�U'�N�{�@U�~-�-q� F �Z�s�╾Dթ��D�7=��HA��:z�du�#�";��DNV���'�]s�+	�p\,��SDF�{bz ��'�����X 75��Z�i��?�X��#`/М%0�C��O�Ⱥӎ�}?a�MO�Tu$�z���0�Q���Z?�'�g�j�	ρ:i��c�E_��?y���P8����|�M��m��V�BL�3�MP�'��$ATM+���)��ؐ<��8��܆r�����!�;�����Nm)U�	��	�'^^F�݉m%�@C�w�*�K��O%un���I��4������@&�t�>E�T�F�))�d�T� ���s�j� 'Q��Pd�X$
T*�p�� �I�e�D`�'
L��&嗧 �>��uH��z�����'�,%�t�7���dT���q@��:��ӣȄ�)~ ّq�\!T\ա��y�*�+��=YإQ�e�'ԨOX�G�?��R(����Y+z���!ky�ɓ4b0�K�<28�@��VW�6�^>f>`��>��`�ת)�2�1��	-n�<���	�aiV#*��a�)��I�1|8��4@��0�I��}T�ÏÚ
��X�C�g~B��k����(UX]i�"ٿ[D��H�~K���7�BV��]�E!
O�"e�[�n�Xs)�l�頔��p<�DXm�,�0v�vl���Y���Pa	)�q A✈eBB�#E��v���煐�J�$�X�	��	#C����$��C��=���A8#��5 v�ɖ�1Od4C��Фp ��8G��H��1Ο�X�(�.���D	�]L�Z� "@�`C�ɸN�| ��
�	F-�`�d�\�7���r�"m �c�J�FΕz�!��l �W
)�'>���gHK�X>���Ta 	̄��"Od��ň۰q�}Aq�\�90M��E�:L8M�%pN�+��$����O�.b�(qe���[�$�s��BZ�h�{��5LOR��c-�tx�x�F�;Vܐ��D�<aj�v��DΈ��h�-���]������T� i�����V�(��)�8~�qO���m�ezJUH�U���O�Z�K�=;��rޠ�Dt�U�*�!�1x��a/ܚ�Ĩ�v�]�V��I�q�r�1�>���O[�h�¢��$�L�k̘֭G�P�0�'��j\!B��aQsN��*�MH�yrF��n��l

�ؾ ��-�6Eg8]a2˞�z����RP�EQ�v|�Y�&�x刀Sv[�����O��cf�T���s"�h�V��㉻i�B$
��ĉ�r�����E��|t��bFO8�!��5����U�՘K�=@ '�\��'�,d; @/�)�ӠF� �n�>$~8h�5+έu�fC�C2�` @Q�M������Lj^C�I/C2�5J5��|�ـ��;�FC��%
�����CH�C��Ⱥ7�	�h3(C��4K����CE���թB6k�B�	2O������Z�<�h��3u��B�	$;�����8��1
���&i��C�	<n�.�YRlܳ-����u�ڳ^��C�ɬI/�Q�	7���{2`*+APB�Il���D���(�,�x��
G B�	0c�%ʲػ>�h�0��-:C�IzpM�%*k]T���GP3>� C�ɛX�t��s�Ѻb�.�ハ�VC�	4`���L r�ԙ������<C�	�z�T�]�i)�E��c��B�	?|�F�:b��+�Ϟ�c�C䉝nCr�㬐�xx�t�W�6͚B�I�c5"X��B�v%
��ՂR�|�$�F8tz��' ��	j�����#v<	�hIh�q�aƁ�y�O�
0�ꔡd,�#i�R�١�ԓ�y��|�L��둈.D���虨��'9S���?-�?)Sbэ[;t3"�3���P�4D�L`Ȓ����Iv���K�'ǟ�y2rbx��]��~Ҡ�)c��&LI�:��`�����~��5eB���� �HC�	�LbT��DhG�2u���'�����F�)L�Q��k��_�~�ĮH���e(�*  Lߪ=�Hi��DꁯZ��	2y�撟����'D 48q���	�t�$��r6�ʊ�dB�(L0D�OQ�2+�R��:�6ͰC	�'Y��j3��)!&8��k�?�0YҝϘ��i����)"s��>|����ځk��H�� �ا�:t��7�ۃo��� �?W��N+%w\��f��=!�Q��t�1g;qa���'Ϣ���B�=�ȩ�$�;q�8��xX����O����U������J�9����9[��B��O��+D�f��$�r�S s9ᚰm^�fHD@(�M0)?���>�(�Tr�I
�T����D�f�δEy�M,�D�~
SN�^��0#�l�R`Zaht��4�Dm��I1&�vM`��D����F�R�bXh1I��
��P���	l�8���T>y(�I����p����?UR&��;P���ar����0z�C䉆s\�����ݒ6%��C��L���	.熔i���Hl��6N�;*�D�9O1�j@w�تf��i �P,G"<���'�T<�p[�<��-YB>9�0��;5@�%��kΜ?т���8��h���E��O*0�O%u�Xpc����5�yI�剕Pa:Cs�S�g������ɂ��L��U:v��T�)��A��(�����ئ*Ɏ|���t����M����ا�	��d0�`@@A����e���
7��y��
<�\�ȕ"Of��D�S����[Ѧ�@�� p��'L(�Ȁ+ɾm:9Ad�
 3�v����yJ?��Վg���P��?3��)ά>%N�8ӓx�|ÔgW]?���,�^�(��<~�*�΍�2P<��6U��ϓV�̨�g�'�D�wi-f@�*gA�?�4@Ӎr�l�(�����ޙZ����S�<Ҡ%BV$�u����(]�:Mp#>٧B�@��� K��ȅj@��&�*��8S�L�J0�ˉX�b���O�m�Ն&u�����
D8`��aH1����4> �=�l���$� h0ܹY�f˜ �]Kf�ߔ!��Ü�g��IR߷`n�mY�*�"�����禥"��!QO�� W�ʊ/�NUA��S�%jL���ˈ+�^u$�OҼ�&#Q�3�X����+�(l��"O�T�� ܗ(�ĕ���Fz�!��	;l�x�a ���0g�-a`���@����ȓCHh���J�pLБE�	�����9
�閯�:jL 	 ��:�4��z�6��� ��{Ծ�x����E`��Ql�Tp��ǫ�(�x��C�1��|�ȓ��I�� �FS�8�<!����"E�	+��O��B�ܝ�yr�T59}n@��쌥z�D4crAB��y�	��0�`c��fD��*���y���1���l��cS�Q���	�y�痤2S��q6i~8����I��y"K86�)��J܅�d���@�y�DIS^������q�@�K�#��y���!��(��C[/oՒšAf ��y�� *wx9�t�H1d�*�q��6�y��_�n��&E�D=�����,�y"D �*0��P���<Ř=� �Ī�yB�K�~D
uL�41N�P��y"�Xy���� T8_�r��)�y��Δf�L0�k�8Vb4p*w,��y�.�(>^ֹ��Ԉ�5"aU��y�ϱ=���-�0E�rͱ0c���y���np���O���mI��&�y�BA!~�|��#��u��Y�yBm=WJ�U'�(���a=�yRcH�b��Q���N�6%$��y� N�I��ٰS,A�^�v�H���y"ϙ��ޅѲfW�V�RA�7ؖ�y��Bs���	[�B���l?�y�,�0�
$Ђʄ�ZT�����y��1?Vl��އ��кCX�yR��a��Y+��	�v���ԇ�yb$� pޚ�J�	��n�S�L���y
� И��(� -�=Kw��:\�X�"O��Ó��7���Rb��O�>hs2"O>-�"ͿM�D��� �`�;�"O�ɠOѻ3~9!c��-L��m�0"O�LKA�� x�x�!o��agd�H"O29�ׅ^�0R�"A�՚d`|��"O�E�'eܢY�:�Ag-��qs򤰤"O.�1nZ�9Ij�:���H�"O4@u��$Ed�	*�e�x�v,�d"Op�a��qB�2�ᑹ��5�a"O4�L�?��a� �9T��B"O�UX�F��v�V��Woۃ{V ���"O����W�N�{3�]
E#F9��"O:�zTK�B1Z�c�ylr�"O\� #ɋ�'pm�DE��1���S�"O�xX�ˌ�}0�]C��Նv�(�u"O�����?��H@�B[��-�f"O�T1ԏ�	uM������4�a�"Of�S�]�-���*%�0*��Q�"O�uy�l��E��E/^�4u"��"O�}3u�_"Vd��#$\C]���"O�M8b�Zo�q)ǎ�62=T��"OܙB�+8����ц{"�\*�"O\��)�&.�]�1hڏe"U�v"O�Iv-O�U��=��D��s��2�"O�Iz���
�H<pt�̓\ Љr�"O��p�G���A�鐴�"OP�A�A��m_
�y&�V��X!Q"O�4��F&�щ���>p���@4"OFи���rĒ%o�#b�>�B"OL�7�g����W��� [3"Ox��T��h�Cv�ϝX����"O�\���!�e�GD`�)�"O�P�̇,B�ʳǓ�v��Y��"O�4!%��e��6'ާ%�����"OX�34EWT�A�HȚ+�؁�G"O��QW�C:Vp��F���"�!6"O��0Ѫ_�H��w�9k��2w"OrL�P�	�бs'���\0^ثU"OJ��Q�\�{�<�҂Kߡ)�8��e"O48��V�7X )��i�@Sf�A��|�)�ӎBL�s�3@�@"G�Vb���ȓ�z��a��yĮ�>$�ȓ]�03a��U��ᓧi�d���ab>�R�e�V�a`�JЁ���� R�y�ǚrxXY��G�~�q��w|��7X:�*@&�D���]��
!|�`lA=%Cf5@Fmɍ���-fH}`g��" 8�C���w>N��b6�1�����-�5@�&N)���ȓp��]�a�Ɋ/j"	0��КE�ԆȓKn�����Ϧ͓�/�=�ȓsG|��Q
5o���YV�Je�t ��X�x�0vƋR��S7�8&�\���@)<���$�� ��5�J��.܅ȓG�PȚx6�S��v9*E��6�&��Ř�#�$A�Q�.$�d`��&�<!�V�̨��x(��=�)��;������#ai��hQ
�R�섇ȓY "H�'抓�&�v釾Y�r�ȓx��;�/���]��ʓ.n�1��-���@篖�s~J�)OӧQ�ɇȓjE5�3n�p�!��M�����(YM�D&�г��Qn���S�? ���KJ�@�r��g͒O8\KF"Ob����D%: �Q��,��t�8�S�"O ���U��6�q�,Rp���1"O�Xˆ���`�q�+?RZXX��"O"�i�GH�HHS2�5(A�!"O�� 4"�;(n2��_
4�j=pr"O��鱄E��3G�_�X�,�zA"O~�+��^�O�n:�G˛W�4�`�"O�y��Gϱ6\<�5LGH����"OJ�C���
�41�H�6<��Q�"O��yC��zO�x��
9T��"Ox��M��I7�}ˑ'����r��'K�<[��T����O�� �b�(*D��ke��+�m�̉J��jD*D���&��"���(?K��!S��)D��2T�\�=Z`�c^Q���4D�h*E�1<I��E��S��k�N5�$7�S����څ�	OEz4���ݿ�N��ȓ;�6�R�X�驁6)� U�ȓADN1h���;,���A#$�/vq��ȓV��u��(ֈ{�H}���P��!�� 6\�s�A�b򔵰��rC�ɠ+���V�MGl���ї`��C�I�6�}��%��Ik��N� ��C�IBdZ8�ë�%t� ���E��C䉔+B�#�\9!D�*Ʀ�\>�B�I�VXT(����\{lHg�C�_g�B�	6�J<#Q�W�y�J	2@����B�I�Bu��8tF�[\<����&8ŘB�I�f���b@�"9���
ςw�lB�I�z+ؤ��/�!���uN�qb�B��4Z-P<+�Aˊ	��/Me�B�	$�4YI�1 
��G��X<�C�"g����ʋ�w��������;ͲC��g�lH�S�s��\�&��l��C�I�X]�x�Ek��"��HL%6^tB�I�'	2q�c�w��D B@�\�jB��$����&ś'4��F�8�FB�'_"Z1����0-9*k�L[�<\�B�	o��p%&�\�x����<�pB䉫&�򈚦��-}p��7�� ZU:B�I�K�j�U�H$=v�	G��P�fB�	<��!�	B��.��f֥\��C�	�;�BTs�&���j4!bHڇi��C��2\�PD�dB2���چ�W~�4B�I?^�,�P�ޅSG�H3�٫WMTC�#^
I�C&�'st��4
��S80C�� v� PY@�ݠK(���C��,WP=���N�_�eS4��U��B�Ɏ⬉7���zC2���Y�",�B�	�3	�p+f+�(j��(#�[�|�B�	OTp
@Z�ax���j�AF!�dB=~0P��.G:&g��J	_�n6!�D�Y���Β򍒶JR��b�'��$��D!B� ��2���A4�'a�M�d�ߍ1c �Y�G��9!�T��'k��1`L=e>:����՞���P�
���h^8q�:X�ը�`���(,�\��	�
v��u,�>��ȓ6�b�Ӏ�\�z_0 w,H&�LD�ȓ$	��w%I-1�ɳ
�s2l��p�E��l�6��I��iY�6��<�ȓ���z���5n�Y���P�[�"�ȓ040��G�?Įi ! �&8 씇�S�? �cp�Թ{\t�8#B�C�H���"O��K�A
=)�ԐK�I�e�M�0"Of	FO1�4P��FL=c~�h�"O��(S`��,���S� �Q"OTqJF(�&`LR,���ʻ@;�x�"Oh�� �C�<��eMK�?􉐦"O����`�}4���N��a�����'ޱO�xRE�@a�92'�
��]�"O��ZRDY��*�3�4L��"O�a�R��5`�(��P� ��Ad"O"�!�$�(����p��[�"Oj�!&���r�xع�]*@�
lA"O^@��ˈh(���\����"OZy��h�b���3�M�Ht�"O`Z�̈)FKr���ިJ�Z�"O�Đ` �	?���ʕ�_�ZB���V"O�@0�M��LI�p,�W!�%��"O8��&���0�Y�f��~�Q�"O������W����$˃�+ȉ�"O�U����>��)�	ӈq�H��"O��IfNG)��1����|�N�*�"OJ-�a�J�uax��a��Xˊ���"O�9	�*�z�t�M���"Or��s�M��D7�����!"Oܭ��A
j\�m'�ϽAϾ!��"O24�F��*M���85��h��"Ob=!ī�6�	�	��N��[�"O<t��kZ:����D���1d"O��k���)���SǕ>�d�ȓgǒ�@�Ϗ"i�@a%g(^~���%(1�����l
��I�>��I��LZl�CsO�.7n���
4�"e��}ה�Y�-�l�b�A��Z�R����ȓ3��tYKؖ4�9@�C�����=�$���F�64�Ā�<�8��ȓr�22��Q�u�(ib&�-Bq
%��?��ȓ��[jh�b��wY�ȓ�d�!	6��k�͊(C\���VU`%�bA�S�����&
�Nq��y��)hG�ՑC m��]!c�",��w�z�֏K?SY��J5"�^�V��ȓ?}�E(3F�*��������B�]��b(& r��<Q�S�ث,:�����ׂ;�j�PA��8N|��iǍ�F�<�%f�9���w�ϝf���@'c�y�<	�9Z:��6��O
�5� �x�<�"��d��P�a�7T��@A��K]�<i�IT#İ�2�L�8]p���W�<iuf���<�ңjW�Z��� ��~�<a!����ѥ�#P8D�"2�S@�<Q��=l �e��/�(=���z�<�CB&1{Q�#%�5ߞ��`��_�<�V�A0�D�(c��c����1 FX�<�6�Y2-�{�d�7d�	Vʏ~�<1>��K�	�1eA*�q �y�<���O(��@�a�(W��|a�$u�<ч��+LQv$����xyyU�m�<�4'��0Ip,��x7q J�g�<94dĚD4���Q��>L)
0�V%�h�<�bN��W_��h6�O?6�PX�jIN�<�2���Q�v�c���#w֐���FH�<)��#�6p����+�\����Y�<���1. `y�C�RNh�o�A*!��ҬLVhy��c+d`�-*���G!�� ��@�$�8��1��)Ԥ�8�"O|�i�k̆J���C#V�'�bH��"OB����4���`� 	�S��!"O.l
�G�o���("J]!%� �"O��KD�q�!2��[�]ĐHw"O�L�U �2�=��a�I��Ԙv"O^c`l�$t'Z{��H��X�S"OF�b�h߶B$`���΍4Q���A"O�����I�5z0��RN�1oO���"O��r��O8w��ȃ��/G�tj�"Or|��C� D���2L�pԜ�b�"O���s�ԲS��|BQA��yK�"Oژ�f��n���@�?U;z��"O��@�E��Wb2��v%ÂA*�X��"O�#�iT�Sn��#E�\=�p��"O�UX��/0�0��QDTa\Z�ؕ"O0�y4���,�h�mMt�b�W"Oȼ�"K�2��Th�6A6T��"OP����/G3����,��H��"O|����r�赪�(c��	�"O� `� B5|�L�Y�&Έb��K�"O���DǨ����^���)w"OH,���74FJ�vj��X5PP�U"O8����a�z�c��-)�k�"ORĳv��
o��Ѡ!��wF��"OJ9����
��3
��o����3"ODd���):�pD�6I��`�t��"OrA��T0	*�����2$�H9e"O0�!#C�eDx9�aKƟ]�e�e"O�Aࣄ q�|�&j�	>Ve��"O� �l�|���8���{���c"O����#)��C�S��m"P"OJ���4�0kp���tE"O¹Ir�<l8$�	�̈�k�I�g"O88�V����i��E2D<��"O���w��K>%�7�i�UJ�"OMPԆ*�t����2zzLa�"O�zGr�^)�GA�c� "O�qj'��`�&i[R�[ib|e{S"O��򕦟Q��Ѣ�_$k�j��"ON�*S��|5l��RÚ#(��r"OF]�̍�ƢuS�T�c����"OJ���"+p�2'HU�{�0"O�!�̞�0	"T٠��j �!9�"O�eA���.�����'
�u�. �'"O6�hf�)t�
�u�F"{)ND��'���#a��C7���$��	��|�'��\�D��n���
I��|{���'��(��&Bur ȵ)ʇ~M搀�'Rĉ����?h4���v��3�'Q���s����E�0Aq�f1�
�'b8!Pb� �M;�X�`+�7}G��'7긒�GF���UiM#-ehq	�'k�����62M���Ef�+G*�0
�'���u熺T�2��`�K�(�@A��'=�!��Iˋs��e�2�'j	�'�m�U�e� �9%����'.(`�4�Ɔ ���I����,v)��';�!��פ;��X����6,|��'� �����,g`85#M�����'��򫘅+��i�c�:�dj�'�� Bfa܋L�z8�v��,�u"�'�D8HuK�VPZ�rV�δwݨh0�'��y��7BFDP���<vޮ,
��� >� $�"���'HB#�V�2�"OKg�$V=�� �-C�1�2��4"O�0AC�[<�)�%b_�a�����"ON��U���5�P��qQ*�""O���AJN*,�@a�r���e����"Od)b��uN�� �PZ��"Obm��.��vD|��.E�	@6IPP"O���#�H�^-�<r��_$*=h"O�(�F��_E�a�"�6I���"O�5��J֬(S-{Q�:* ��"O��0��]5:[(��M$G=�1�1"OĤ2��:Z���@|���e"O4X�Câ6���K��ȳ7~��Ӑ"O��XCݺ��0���N�Vc�q�b"O܁ �`�{�e���[�2b�1��"O���Cƽ	�f�"��2t^̻r"O�X��[$��a�F����6"O�iKń��Q���s�$��]��I�s"O"��+ >��3�$V�$�w"OVyم�I�M���
� ]����� "O\��F�: ^H�1Q�Z�fh �"O"��#q���t�[����×"Ofx���H�j�y0 %7Re����"O�i�nަ0o�p�i��4Q�C"O����E�&�u�G�C9Da��"O04�PL�I�Y�0��1A؁c`"O�)P�&��A	�e.F��P"O.�H� S760��ǲ\'�
"O��(U.S'��� P�<!�"O�84 �N��9��h^�9�"O@x� ��2%>-�����&��"O�0�C��60�$9S��~��г"O
P�h��0� H�!��$"""O�1��¯]��'�.��y�"O`�� e�-$�2�)WdL��4Ia�"OZ���GUC��puB����A"O����W(\ΌA�
�S��da"O� �O�Eď�l70� ���"O�h�dMS.�b�z���zy�5�"O8�mš-�ȩB@K����mʳ"O&�۷"�5'h,��
�1�f�p"O���'�o�&JDǒ�8̰�q�"O PJf� 8�:EO5OrA#@"O�5"��q1�x�ţ��Teڄ��"O�HB�Ǆ1)-���1-[�-L8Ԙq"O6s�O�=S�	�7��-8|l�"O�zGi�j�D���*7�y��"O8�Ѵ��J�6�vǘ��Ի�"O�
3/�8s��J���p�V�a�"O�1Q�k.6k�LJ�Ƽ+�6t�b"O0���+'!bej��޼3�dT*�"Ol�1W�ɨ~R�<�GT$Z� ��D"O^��Ǝ]�)��i��������W"Ov��ue/^xb֦\!����"O.I$�����J�ʹPq� k�"O���CɃ4��q���o�ޤ�f"O~	��\	i?<���p���B"O�e�?�4��͖ �<���"Ol�C�����8RbG�_%�!��"O��Z�:=�L�9���7���"O(	�5>�j�A3͙#<T�ԩ&"O���D[6a�*%�"X�SbX��"O��t��2D�l��`B�[0����"Onl�e�I0.A����II6#�\C�"O� \Hz�`U�k�`���2���"O^�h�P���4��M�d�Dp�"O��, �i��T9�Z�<D����"Ov��wIF:�L
��S	2B�F"Ojt����	Wc��P4�0��:�"O���"C�w��#�Öw�N�%"O4�[��۬��=P@#�0F9җ"OX����=�D��#��f X)�"O~�q��Af4
	�s��?Pd��#"Ox��C�_l��c�.�''
�����c>e�d���x�d`�.�\ytЁM:D���&iԒ`σ
Ǿ�� S�y�!�d�2!x�r��/ �d`Ѯ��0��'�a|�d3Lcҡ���7��-��BU�y�ImD�II�Ϝ>y��p�c�.�y��ӈ/�<`q�C��T0c1.��yr��2W6l�[���)�l������y�WR^Q���2?2�B˔��yr�M2S:��"��	�
� 3aN(�y�A�l�*�S�,��eO(҆� ���0>9`P %;@m���6��̨u��d�<) �
�N�JUDH�7���v�_�<�� {ʦ\r!��4;�\��d�<����~4x �Y�Fo�3�Jx��'5��H��ғ/-� Y0Yȥ�	�'z��T����^2z�ɋ���$3�O���M�;&�H#��c���5�����2BtXz�a˭;d���#�O!�$_�d����$
?'Pʑ�5gɼ�!�D�Du��٥�U�~�N06�ΰ$�!�dZ�:e&����2L_�� '��x�{��'��I�m�j�j��ȧ�b${e$I�3iPB�I�~�v1Hb�0"Z�9s��6�0B�IO`	Bqn!/<"0�C�G�d\�D1��]�O��2H���ږ�];�i�g⍭o!�D54�f��w�þF�R0H�6�!���#��x@���r$�Z�/�!�d�8���z�k�&a�xݙYaصϓ�?����d�#p�:�/�SN��EQ2 ~!�J�T�Jͨ��W�\�t��f�`	!��]�E��!SmA�v0dQ�-�!�dt�N	��3s�@�k�A�!�Σ~R�rvi�&D���8g��*�!�A�\���(��W�pؓю_Z�!�Ęqk
�p�f�v��Y�e��<�!�*_���"k��U��]`��܄?�!�$PS����6A�����	�M�!��ͳ"�E˃� �+V�5"@�!��$w�~����VVP�a��&}!���5�ȴcE��:r.V,q� �%k!���[���J#�Z1'-�5�ǜ53p!��Ćc�=�D�?�<A�"�	6d�{�Q���L�HP�c.o��ܑ���
=_�8�ȓ�
�6$+t�h�ӧ�օd�nh�ȓ��u1����k) d�S�Ţѩ2D���r�� �4�BQe�l ��l$D� �4�5$1L{�7-ʀL 5�<D����E*wd�4�p��I:D�t��-K T3 �R� E�af�
��$D� �T(�D�6M���B�d�^�pp#D� ���׈a�=��K6�]�(3D�tH��"$
r�� \����>D� j�`^-&)��́y̤��b�<D��
iٿ:�F��4&^@�>Y���;D�� h��34*����l�?4�^I8�"O�5����%Ǡ�pq%H#_Z!�"O~P�RB�Cq���qĄ�pL$A�C"Odz�c��p)q�Ӛ-$� �"O�1c�B��w~��uaFPp"O����&��x&x#F� �,��S"O`y�!m�
W��C�g"E�I�"O���U'WqN1� Y>GW�ű�"O��qCɄy��(ha���y��ڵ"O@5�G�1�MH�	�f�򈢲"O�ͱ҆ɭTa�X��gŊ`UL���"OJ������څF�)X*�Qg"O|��t-IW؎�b�D\ L���j"O�`� A������"�u�:i��"O���eA?��6e�/F�v`q�"O�(w��X>@b��D�d{ � �"Ou�4�)G�5�,�$
���"O��)�� ?<Ĥ�	�#c����"O����$ɇDf ���hڍ 0��{ "O�	3k�k��q�h��g @��"Ol���!
|
���d�R�̭qQ�����!V�v@{U���6�����a�4C�	<<��� A͟d���%�V�C�	�7/A�F��B`�)H�
VӲB�	�}sԁj��\	�Qʑ�� ���`�@�xdʊ$��C��F�-���D�:���h\�A{e�W"�P�ȓYuƩ+A[D�^i��)�I��4%�ԇ��%;��0a�N�V��}�5���Q�bB�I$i�P��W Z�p{Ul\�J�b�?����ӫ��yg'������-�'��{b�$dd|P�F�(-��9�!G�_���IN��8��eT&sgbd-40�`��ѭcUB�	.1W(�!'t�e�VI�"S����<?	s��v���0�e�6XR�W^y��'{f�KV�t�\}[��ѱF��UK�'P���C��!ub��JA+ �+G�hA�'�����6����%_(�,��
��O�d��G�1�b��5�ށvk�U��S����	�6�R�A�-�W���ɤ�ť8[,B䉡n�b���1�l<���&cf��$$?Y�n�Rnj}��/ņK�DpQ���t�<��W&H��u�d�(��uSFk�<ѡ���SԌ�T醋z��5QFg�hx�dExO�5�C��D���sD��hOjʓ�O´2�˃Q{6`q��T�5=h�_�Ȕ'waz"& �O-Z��U��B����[��y"�U�7u t��nC|���C3�Ԗ��?	�'
�$#������})��D38���'�.y(cʁ�X�����8'��p�'c��ٓֳL��d��fD�1���3��?a�y�(��*���+B/ۂx�ިsCɀ��O�#~��gL�>̌Q�;t���s�z��M�̺�Z�28Z�l�M!b�q��/D�8P��]	��L�ǫE����#D������~�0���	�-E�i0��"D�4Yъ�]&�1Wfć`AXDF!D�TAu�Ѝd��	��h��^N6e�č4D� �@��6}?*��H�/�K$ �O��0D{�O"���'���Y�s+�5 HA3L>�	�A�X�Z�F8x�b��d�ȅȓ*��i�,5���hw����\����bXA�o[�JD tP��Ғf ��t�$D��X&E[�2?x�C$�ó�*\�d7D�� .Ys"��>!��abbŝK�p���"O�,�Q��_�z�s@j��Q$"O��+ �:@h�J�,[:z�,��d�Ir�O��A� �A��D��"L� �'w*e	���%�ջ�� �\Æ��'(T��q�?��� �S��Y�'��]���T��แbN��a��'),�c�DATG�D1�	Ħ7�`%��')���-].+f�@��.j(���d>�"���j���E�&�\!p2�X� "O�f.À[㐄ɰ�� t�n=y�"O<���<�� ����]; ɓ"O����!�B�(�����	7��zc"O.P���a��)1gP�g|�(6"O�Us��L#_:�Y2 ��f����"O��qH�x���B/C�K��'"!�D�t
#��2{���LZ!�R�|���AZ���A,�5!�^�V4҈Ȕ�B)�du��+*(!�� 2������u�Fi����.w!��z�N���'ߗo�~�3P��?�!��+m��}��E�g�Vz��Y�S�!���\��(3(:��%XԈR�zl!��$L$		�!���9��B�Q8!��
@B��E�Α	f�h��Ļ+W!��Q�F��ƊL9fW=9p�H�	!��El^\���W?bTr���`ǀ^[!��,�L�s�]=0���#;�!�D��J�tp�Q�ď�a����A�!��N�����J�^v�U#�L�n�џlF�$E �b����V�B3Pzx��cҪ�hO���i�!E��c�C*XF�����!��>8�P�ф,�0.���N�h'���'�����Ą
�F�h�ů5W�e�e�'�!�d��=����4K� .T"��L�q6!�$U'Xꚜ3`��;="���u���x�!�@/Z�쀆����8"ś�z�@��?��|���4'�J�sT��P�
_�����D<�'Z�8#��N� ��-	�b<ܘ�ȓ}�]䂅!�d��U�����	�<	���#o�Eɦ#����Sp�� ���j	fL��ؾ�2`�p-]�DjBP��Rw0%�1�A)(�L�I3*�2xb$���;J�ɡ2�������GV�
�Iu��˟D�?������R4�P�gC�aYU�`��ԟ(F�tIG�--���̊�4jx���E���?����%*���%F8���Sh�3M�����r��B,KN�Y�,�b�> +��؇���VY�2�F
$�U�����?B���9�L��%�]�{L���aZ�b�M����<����32;�E����l�vI���ny��'j��b�	^���f�\x{��$�O�"~���#�~��򪁌_{�$��
�i�<qvė�A4��ab�Dq�c!��c�<���'`��/q�~��2��t�<Ag�W�)�H����'\VQ�S�g�<Y2�1C$"'N&�����c�<1FA|fh$:p���",<��'�]y2�'�B�K��q|��X���*A�Q	���5����re�:Pc��L���{<a`A��I�H�YV+[���9g�N�<�P�]Bn!�p  ;c_�@1jQH�<�FZ%*��݀���9mМ�V�F~�<)1ȝ��x����5hǤ��V�Yv�<� D�԰Z���@ �0"J!��"O��q� ��vt�z�F��Z��=�F��ȟpE��	�.g����5�Q3���҃�]��y+'t��X�!�J�e#�E���y�����k�醦H�����Hٱ�y��^-Q0`M#��J$BFI[����y�ϖK000Abȥ3s�8s	��y��Ǻ��!5�T#$*�aз���yҌ�$`l�BP��!���J6�)�%��g���Lȕ<!���]x��P��V_���U+��0	!��\�nqf鲒�^7RE���J�$y�!��:����g�a3]!�)pq8�'��l�+\�P@j����>��z�'ޞ�k�8`ٺĢ``-] e����'�ў ϓg�v<����w��mۣd>TK�=��e��˓'\/w8���۶7��ԇ�T��)S��5I|��P�.,(���iXN�(�A�v�:q��l�Z��ȓ������(�i��\({P@4��>=��+7K���C#
JZ=�ȓ<���;���a��tufB����ȓ �M�6H�9�h �d�۝9�.؄ȓ��E6Z�J!R��G��4ȄȓYv.�3Fŉ@�:�����	r�q$��	V���(C]�k�L����!"�L�&�"D��eʆ;Re�,P`�
��x*UL"D���*�������@ e�'B$D�l�d�atR1��ìd"��C"D� �*�:��c��*r�@��ì D������im��+�BC�_\(�7�$D�#$�'o�l��C%U�d9��$�$�O�����hb���!�#O�dY�� a�!�@��Bp)�"$WP����_�M!�d�t�2�鷢]�y��B����r�!�dȡ3��a3H���d�ɦC�!�E�gh��]�Nm0��@�:�!���YNq(t,ۗ����*?;5!��uG�bW>_��p��^5/!�ď�vM���a/ T�8 �7=_!��	�b_��1��A��dd� \l�!�ߺ_v�����C�X���=q!��]�[��z1/֧'���h�/�R^!򄒝l0�ĉ��ؒ$�NP�p$Yq+�}��q���p�f�SG��#!N�B4��OZ�D��'􌘛wTFɄ��퐜"�n���'�Z�(�A��,�����I�z���r�'�ax�
C�z7 P$k�>y���PH���y��.���-_�o0�#��%�y�k�1����I:�@�@7�ʋ�y�6��<��ڌ68�5h�K�7�y��ɚ8ؖ�s7���/0�b�G�#�?yI>�������IG��\��	32�x0P'j�-cfC䉟jev����Y.&F��0�\6��C�ɍI�F��&aX�wx�) ��]� B䉉\��i��f@�HB-+�B�	B�.|�I!r(<�:�&�F�xB�	 e��x���/+����,ݤm�NB�	�B��lQ���="��������B�ɋ1Z����?r�D;����B�	�.'�,{�L�5U����ϙZ�2�$��I6>���R3/�!��s��
/<U.B�I�X:*�xSEӎs@��`jԯ2�B�ɖr����aE�;�X��$��B�)� �� ���&  ������Z�T��4��p>�9�k�1�PC�%R�N%���5D��Em?&|	`D\ryء+4D����IN�Bt��3[zi�u�O�=E��$���xI�Q�¹q2��#s�ЛS�!�dԅk(,"�A��$+~�S� A'w�!�Кg^��D�:��I{���
�'���Rj�q���[���YvZP���D8�K� ��g��=U$��FiJ�~r%�I|�����	P(�|�v��.e�#ס��^��B�	:R��t�XQ(E�R�6TLC�I�5i<¥mW��<�[R�ћ6݂C䉀g7�1i����	I6� ���}xTC�	�p��3�G�Y9�abc Դ>�nC�	�r���j��x�ވ9�͵)�T���7b^ze�Ch>	Ñ���ee�L�����*4L��T�Zf��2z[�5�ȓ\*4�j�-��:���f�(P�J�ȓo�*H�C�܂ ����Æ�PAL���x�$ۆ���]r����Jb�,�ȓT�!Iœ�a3|<��IEML�ȓz�T|*Q��� �r4�A�݋a��5�ȓ,n(�v�4D��`��ET �dI�ȓr.0�'�Ή'�������{b���ȓ9r�� В<\�l�POg[T�ȓ�RɈE�^~��[�-�=�n��ȓq	�z�A^���k�)]F�(]�ȓ_?��$d܆S� IG^Id�ȓ�: Xw(�fu�Y*A�6yڽ��Ie�'"�]�`�_fn9�t�G5h��E��'�N8����4�D9�LD#*�V���'�X��W P�Ҹ��V�4HJ
�'�Y#̨~�Pw�G���y���g����E
0� J��y��M�2L��㥡�?��p%���y��6*t���珖n*���߰�y2�^�!<Ȍ�K��e<8Q8����y)MEl����)\��]�դ�y`�U�U�1J0R
Ta_?�yB��CLf�B!�ĆX�\s�H���yb�_�x�4� ��:s�������y«�;�l�x�C!2_���允�yr铭=8�e锨ִ<�����&��y�&(��\��I�;pA؁��8��'az�CT�}�@�8�(��]@�1�-O#�ynHA�a��/D4����6�A2�y��ρy���%)�ҵ�����yr,�nl&���gp�XFh���yR�&h���[g�N�an��ӫ�y
х]���H�χ�f.�i��ʖ�y2(ýu��*��i��i#sdձ��'Paz	)p�P�Ɲe�hL��n
��y"F���Lr `�3a��
QD�y�0�����욵p���8`��:�yr+�2�4��j=d��P��ڣ�y2�!	T����"ѰaO�u�&(B��yroSz�x��!�/"`b�a�mG+�y2GC,N�di��˕�����$H"�y�@&�HAa��HPfh��P#J��y�� 5,/~<q1��PR�Щ�)�(�y��I �<I�P��K]��r��Q��y"�Y��R�׫6L��p���X(�y�Gԫm�rcHҲq��{%F!�y���(}���R�\�J H@-�y
� �-��`��ijz)�eQ�w.��"Op-{����+�P ��)m�H S""O��y�ݫhX�04�����"OZ�20�ےWBj]㖪����'"O�+1,ƞmũYh8 \��"OpYkP�9W����� ��ۅ"OB�K�� �C�9!���)�B�(v"Ol:E�<7�X [&�"����D>LO��P��ރm^�Y���  ��M��"O��q�]��θS+�&Φ��'"O��"�
L��2��5G��4rf"OV� ��i������
)u�� �"O�5ImC<��R�f(8	e"OU���(i�B����9�DQ�U"O�I��l��/a�t�EK��E�Ґ��"O�Q#�LQS�Z`�j����A��'�r>O~�1C�ھ`��9�	޷/�<@H#"O����1o��A�t��m�����"O ��F�R5-��=� � e��#�"O�/Y�(s��9�-��qQ��"O
5Q⧄�$ߠ�� O�<�yQ"OT��RDҦ#��EH��������"O$j�i_�3,�a���6!��щ��'�85���[�"��,�/=49�'r�a�lG�rf2�h�=w:��	�'��t�4M��V���ZSCO**&�PC�'�h㶁��W.Tq�&�r	�8��'uP�	�@�#24�� ǽn(�L��'�rMѥ�*�I�W���T+�'6H4�R�R�y:Z�;)�� ��#� �^�e2��_{�a����+��B�I2!�h#�Ə4P�޸`��k�FB�Ɇ ���fe��j|�sө�?�DB�I�U���R�ڒA.�q�&'֌)q>B�	�-�`$�!C&4�����!
��B䉦B�>�C�!]�>0�H�E�*xI�B�	:��8�ǔ-X.j�ǪF5�C�/ �KE�͆s�D8�!�)[�B�	�����$��"��VB�=z:�B�ɐ_�Zը�� ,F�$ �럂<=�C��>\��]�"��4�#TE�7:#�C䉨#���yc!Z;�`p��ƁY�tC�I�z�2���j@�c}��rG�P3
�
B䉵�����ŘGM\���&�f|���?	���?��'6�~�Y�F  0� �ЙB��4��u�j�QgG~�!���e�4��*��HZvd̸<��W��� ~L�ȓ[����"H���Qyɛ2T�n���C����֐��Ip���K��7rĈ�U�8D�,��ȭ[����fZ M{�(���#D�t�H)1ժBfY�H�n�#�&#���Ov��>�+C�+	y��E��<X�{�� D�\x7"�>`Y |(�$ �G�&h��	*D���DoS6b���;&ȈR� �D(D�4���~��8c���@�r&�%D��[V���Ki�Q��Ņ����D�8D� ��֘L~^!a	�c2����,D��t͖�-p�P�C�jhd�0h.����G����		�䘑��"D�<��1"όUl!�$Ru����$�-s������
b!�ʵm���K5B�Q�Z��w�+Q!�$�mi,$)!��nQ� ��:<!��0I0�@&��08 Ud�<V�!�=�<�L��I�P���P�!�� &J��J�)Bth�(Q�9X�3��'��T6eX�H4\��"�N+
��-���;D��)!����I����5Q/�X�c�8D���A
4`�-X�O��JКq�8D�p�B?]v�ZF2j�P��ѧ"��O���J㮀$R�]�q�Q��H$�+D�Xr!�3�&�c�õ/��p�F�)D���MW�lB�4x��Dh^"Ppv "D�����
#xyF��D;V,Ru�u&>D��0�ֱe�fIXsf��	�Xĸ+)D��g$���,iQ�0u\�I��(D�XPWM�j�FM�a�v_(�ҁ�$D��a�jJ�L�e`� J�H����<��	vBH�#\8��fdӄԤ���I�<Qb�ҵ�7-�h��! %�hO����Xn�0 5��%���C"��]K!�ā'����o͈@�l��F˙�-�!�$��.v��JC�S0�
e�'�]�5!��˹t�m�р#:uhwH�j!�D\�%j(���h̦"@$h�jQ"z8�O���)���Q@nd�2�˰�� h�j�`a"O�Dx ��JP���Õ7�Qi��'��0��IT�|-�R�'`Y��r��<�M�B�Õ��I@T�`����d��b�h��Ť�
Y^�� ��WфĆ��ß��bk֌9;tir��9��IA���ȗ'Tў�>�a��H�s7��Qo�_��<s"�<������(��IX��2oT����O: 0y�"O��Ŭ�!O0x�����1v���"O�y�$'�
�ƥ�DF �t2���F"OᘱD^A�N�Y���9�ȼz"O�D��lY�	�FD��7g�8d�c�'��$�IOH+ѡ�0X�����/ln�X��D{��4CF> 9��*'��p�e�J��hOp��	@�i0��!�f�)4*A�� _�:2�O`��<ђ����}����"OR0�	,QR���D��ȥ	3"O&1AB@Y�^@�A�F
+���@"O­z��խb��x1�ehM���'[�,Si��\�.I�b��x@VB@Ht"�|��'�O�v馭h��P�+~��¢o�x"ą�g�'  U[��Hb����}����r�'KP=3�� ;:���ʶ]'����D ��M�%끕Bj��c�*8�|t:U"O���:*��+�eH�G��%�2"Oܬ��̙�=�Ptb7�� �:hI�"O��j�/6�
�B!
H�dU�ɳ���q>Y"�U��0��1dP&Wǐd ��3D��RQ�R'}�F�!��M���c�`2D����X�eJ��Wɇ�7�~�@P�,D� 0Fm�s�X�u�
;P�p�6D�`K�iL�,�>QkI��)�@�B"�4D� �G��H��[0� K*��3D���BB���0 �0lƻD��q!>D�Ԉ5n�)I4&��!�0�����!D���'�k����5M�! V��<Y�~�&\���ǈg��I��q��y҈�z�\�����9*�X��ҋ�y2B@"��]jN*~�6m�:�yR�8r�j���G�f���h���y������ ����cb)�y���c-���DQ(tV�ac�hH(�hO.�𤒘>���4�,>+*d�ux!�$(�*����ܷD :����)8�!�� 3�i �0CeQTֽ�$"O�}i@�_w�<�Ӆ�w :M�"O.�S'�����Ƅ5��E��"O�Qf��F��MS�����8p"O:D#UN�#;�����D�4b4���@"O6��N7t�����ӡ]��6"OR�I&�-V����/�&dA�"O�S@��O�����8�>-�q"O6=jDG���B�]04pYj"O���BG�	�x�qpb"B�p�"O�c��ۙrch�@p�J@j���"O��x1�s�"h�r��,�ʓ[�LF{��Y$J�𸗃 ����9C	ȴU��D�O(���O����O">Y���hS��(&� �����e�<i!�C
�֖��R�Q��[�C䉛[O�|Kr��m�
�rS�:�C�	<o���-���xIì��<~���Ofp��醤HYҭ�r)&]�`�HӦ7D��bX��ue�/k6\X$n�O���OB�O?9se闕h�Ro�S�tБ��l�	����	��x�	P�'�Ѱ �W�V��&n����'v�R�
�1V��2��'q�v���'��)��#��إI�h�q�l��'"D�F
�c�%��+)R�`�p�'�6���Q�?64(X��E�X��
�'VL���E�=�ba"D�o�l��)Oh�=E�T���S)ĉ+q�;l0���VdW!&fb�'��'er�'4��sW A2g�h]R�lQ���1G�:��0|2r��.=Y�97H�a��9�c�q�<	�_Y�=���G#E��l�FEJm�<)r`��5CBHRa��!-8y��N�<�O�7{��Չ2�U�F�P���R�<�wX�猉\ĺ 2*�w�<A�E�Jc�9���	3����%B�W�<�KN�[��U��1U�<��*�[�<�bhZc��J.	�1[�:娇Y�<�SfX�Oe^! ��XN�܀J�Q�<��ʟ��l���ݽCMzp��_�<��%�p �r�'�<�>�7�t�'�a����=,�&	jd.#t�F�a��O2�=�}�3�H2�A�o�l�l#l�d�<�fO�)[Q)3(u�S�#]f�<!��H+v�T���Me$��3�j�<1�KG�����K7�<�Pb�f�<QR+�� �4���G�;�����e�<!��&]\��B��9Zx�3P�X�<����GV���$&��8��+�^P�<�$m jb�+B4P�-���ҟ����S�Ft�R�b!"�;�A�Cyp8�ȓ2��w�8;V��Qʂ�s
���itfq�E�?7t�$M��X��E�ȓDD�!�͆`���� B:4> m�ȓRSЍ��X1Sq~ #`D �pلȓ1�����䈧vB��j6 W�F����ȓu�.�R�H͍����#�V!x�
̇�b��L���W^U���O�m��L�ȓ$8�Qqn +5uX@�fe�_��A�ȓȪe+��MH�psc�Ԭv�ц�Rh
��e%��	Jn��@�{����ȓjIn`�	P6 �� ��\,Z9��xl���Mݛ|� ؚ^礥�ȓa��H��νfYh����m� ����R�L^��<uq���/F]�-Ro5D���D#��u;���*S���!ڐ/5D�� �D���H�,=�����d��Ä"O�0'L�? 咬�ק��x�� &"Oh����ɳg��'g��N �� �ICyr�'1�������2��`d%��_�R�2�"Or�
c$6GY���CϾ-~pyJ�"O��@'Xኔj�$Y�:� "Of5��ȔP���㊞.���[�"O����.Y(P^p����I�T�p�"OD�A��Ú�p�P%e�����"O���k��Su���`�Ȝ	<�9��'�X1HU�H2N���dDR�O&D�(�P��li0 �@2w!JP��A#D�9�J�]�(1��*OP�c�+ D���fLG�s��R���(�j%�C�<D�h�A��Je�Kd�:_��"�:D�0�G& ـ�3�n�),Qz����9D�p��!@&�j��&v���d�8D���&�!6,y�����o���8��6D�|z�eܽf:�M�b��f����=��0<�!Oy�9P���b��-��!�b�<1�_�^A�8��6�zd*@�9T����i׀2���/MFt\Ly2�?D�T��+v��˰���Drq0D�h!V�J����1G�|����.D���D"|~�-S�gݚ%�l��5h7D�8����hۖ-��d� [`EА�9D�dx橘�H˾𠔥��M�� �u 8D���V���0 ��%f[�<��5D�Dx�L�/N8�k��ڦ5c|�"� D�����ƹf��U�Ø�1t�*ӄ9D���H�Ǝ��i�� l����$D��K�c"Oj���$��h��=D���c'Z�"�⦭ΌeJ0�B�.D���0�z)6�`�͎' ܋3�-D� �U���V�����(7������0D���ڇ1���%�&G
��:0�-D� V�m��F��-y�|S��,D�4��F�'I2f\�p��.㘼�3M-D��0k��H%zH�4��N^`�i"g7D��9SfU⢵���J�s�R��5D������C�0��S!H�K�b�i#�7D��)�%�#/:~P��M[�r� @�w�5D�;��ҋI���J?Z����5D��3.^�gE�8��g$f�42D�\��D��TX1dZ::�H�h�,D�tQuh�3,����Q���I\28�UL5D�$s�䞙I&�A�g%ĨX�l�@s3D���WɎ7{P��sK��l�P�*0D�$`%i�����S��� X90�m-D� ��J7|�f0��
]�TY0Մ0D��(5KH+p�0e�@�Y#Z�"틗c/D�ث4��]_����K�e_�P��!D�T�J�-�N���ʥvT�Q�`2D��Ţe��C�%�@*���b 0D�`�5�R?@$��Fk�:� 苵D+D���7$^�9Ũ�"�'	&>�^]���>D� ʀ��Z!�a
jF�`�@-xO>D�p�L�;X���=lZ½2C:D���U%ˠ7I����MS��jw�7D��2"�*���3#�3�jA�Ê7D���0A��`� G�M���6D�4s���6)��I�Z�؊s!D����JΚlؒD6�t�Q��2D���ؓo��)�RA���j���1D�� D��sE�#p�0p7���Q��y�U"O�p	���9�qaօ9s,Aq'"O�93��-����q�07� �"c"Oآ���hD)�,�5`�.�c�"Od�jTIg�'�Z
px;�Ñ#�y�@Ȫ.Yܵ!��2��5�SD&�ybB" ��G'6.z6])#�2�y�"�H��.�6��3f��yB�J�oS@|��g�J@���y��B{�&��_��tx����y��Mm\�r�J;lm�)Q�y�D��d�5K��e)T��_~j�ȓ?h�H�A� Բ���E�ڨI�ȓ+��<�3'ڴ�(�qe-̫Hr���ZK��@�-G�z��3g
$)Id���_C�H��X1�P� t���[:.m�ȓ1̌17)��4�E��ǋ2`�bX��4�<h�@�L�y���"���؇ȓk|1�cj�Ĭ!�,��	掅�ȓD�t�c��4hX&,i��v��ȓX�$ô�O�'�"� �쀲Dך��ȓ��0�É��J�%)U�;aP��ȓE\�m[�k"�MP���MZ�E�ȓ+F��)�#�"�k���f�:|��V7l�u�خOg�-�0�-�t��5��4	R$8RY�G�Υ;�����Y���ǋ]3� ��NN�@9衆ȓ�Бv� p��5��a��V�%�ȓd��)�Q��&��h-�}ԅ�:5h���K�Yܐ����N��ͅ�6�h��]4�=x_c~Esw"Oᱡ̅�B��iqV`�iOH)s#"O����L�b9����8B\�"O�T��l�T���&/]�g'���q"O\(����V��d�V�W�Ƶy�"O�`��BO���1wo^=z�����"O,-��&�+6�*�@\�3֖�CA"O܌�#�ތER��1O�I�bL�F"O8!c�	�!���s� � ��%y�"O�M��)�o�|���\����#"O��Q�4hx��	�$�A�"Oz4J#kj��͠#�B�%�q��"O�y�_5vbX�SIN,(�@���"O,��b���Dn (�P�ۤ�~hBp"O���v�4�R�Ӆ�z��pr�"Or�0
X��'� �Μ�"O�yS��7 ��@���3F�\!`f"Oh���9�$q�[�l!�C"O���%�C���;A��'݄���"OT���f7Aw�M��B�g��b�"Oތ���^ .��|��	�w�P��$"O��{7c�x&B�c
�	>�P"O.p�t@�M�Řņ��4�<��"Ol0�S!�����r��
T�4"O@S�qO�����[��E��"OL��w,_�#�F���	x��B"OZ��!�S+&e	lˎE��`��"O�I+�B��y�EY�j�,!L�`"Or�ر�ΰ<z^Iŧˠ8{
�B"O(�ɦ��-:D�:���(H�t!�"O��iF-ŉp�da��g_����"O�l�e�]�Sq��+cG8%T�d"O������/!0$�G�^9���C"Or���'D�3��r%��=�D@b"O� ��22e�!V��Q�R5}J��"O��r�n̽A]�M�&�}X���g"O�xC*.�$�x��&[Tz9#�"OXp� K��+E �Jç� �"O,Bw���{^|`�רQ�6d�!�""Oʕ2T(W63�q��$��3/X�0"Od��!V�Z�Z�Edr��"ORq(@��w��m��DQ�5���9C"OT�Y�5���8�� ��a�"O�D��q&��Պ�GkJ]*"O�A�a �B�>�TC8�i��"O<��� P!T�\H�EB��NӴ��"O�A�C�Z�N���Z�ȵb"�A3"O�T�5�S�H4���C*	@��G"Oi
�j[���9CQ���s�j]��"O���qh�����(6�I�"O.�;d��!~n��
`.	�o��<G"O�Ƀ�E�o� �9��G=!��$��"OT�Rk��P.�У{�RVp�<9P�ӷ1%�;��޵}�Mi�%p�<��l�:8�x�;+�}��Q��T�<q2/��]Tj5 �"ϯ%X�)�N�<�3�ǚ*�=P�(m�>�A�kFH�<��e�9���`�K�f�2�o�M�<���.R�uJ𬟝!hl�j�~�<��?��T0�͘i�|����e�<A��7vg���r�W�yV9CEn	]�<ɥ��Tf�A��^�=���"A
�M�<�����@ƃӘ/,ѱ��G�<)BEMQ\�y2�-"j��!!IG�<�g���C��K�HM7q(�(���E�<Q�*-	)�D)3 �>m:2ؐ��El�<ya�**"ʙ	C��X���<ɗȼl :���g$����hc�<��J%|W\9��Y�:�㔃_[�<y�BR�S�9���B�:hKQ��[�<q�gT4~4 P
�ˇ�}��ف��M�<��D�5D� d"�F�X��SA�<!���5\��"A	�Qv��g�|�<Y�/ʆT�p�K���,��u#1D@�<	G.Ŧ
ά(
���H�.ia�<Y#� 3���r�V� �[+g��[�<y�c9,��ͨ�LG4�R�����[�<i�i̩5R So��&��Tx!B��<I��� ���	�U�rtDig�<�go8y^lIɷ��,w ����H�<A5`�C6~h��#�$+WJ�#K�I�<��.�qP�iw!�	#����%�Zl�<Y%+U�@3*x�`ɱ'�@�<����� �PJ�	��p��q��Mu�<�7HF�R-R�p������V�<1/��*�Ұs�C�n�<=�eZmy���v��J>��	=q����G/�<e����<�S�G���$�j�cۜ�S�(f�����H�8�I�bC x3���t�G���	��p>�Co��A7�� ���2T� �Ơ�R�d.�S��	�>ᷩ!/���񌅓ښ܈�-N�<i5G�, �"E��zed�qV�#Ⓚ�\��%�.��x3� 
��`W"O��bEe[.�Qj�+��L�P"O�E2`�,U��%���Q:H"D[`"O�Dӊ��9�� )wF� "O|�g��K��D�Pb+�u�'�	_8�(ӱ�͸ �l�:T�K�`��;�7D�� �q��k�U;w��(��u��iQў�E���A�a���Ĺ"=��AD�����>���<I���Dz[t���nJlB#c�F�<�rG��9q8!�CC
�#&h�� ����P�=a�Û����'S��	��:@�'*
MBلȓN�l��/֧

v���]AJu�d�'��O��|?L<i��yi<���D6�v�#3K_�<e'�h&�1�&���u˂��~�<��!���zg �,%����#φ}�<�%ɜP�F��C`']!�x����t?���'$��t ����K$�X#V`<	��(`��� ��de��#��"\}��8�>��G�Q�� �to�:zP)Fz�'(����[�g<:��ա24�	8�'gdq���Z ev�W��7�%��4��$1�Op�p��0t��h۱(?Pz5�|�|��'�.���fS��&lC$��Ĉ���1<Or�bpG ��>9
1���cE��y�On4׭�	��3�¬Bv��H$ˏ��>��'�	J1K8d��b+��SLD9�S��Py�F�o��U�P��*YxZeX`��\�<�N\�~�JC�޺Q���{5�X�<!��/��e��
N�Nj�X1�i["fў"~�I�j����k�A��f^�a8J���>��@���.����f	rf���0=	N����<^����T�r�
R�7�O�O�Đ%�C3�l���	�={N�;d�I|���i�*!.��`Β#$��Y�&$Ä1�!�d٪>I���Ćl��cG�ў<��ӭa�̫���L�@�õX }�,C䉖!�05�b��2"��(�Ⴠ�UIC�	%J�����hN�\�".˱3��b�L��	��![Q	rn��:�Ȭz��B�ɹ|��+��� ��{������O���?�L~�+�^@���^�fyp�qt ��]�(m���t�O���F�ΏHQ"�#��ۯD�p|��{"����<іƑ��:	>R%P)h�&t����?��A�j��\�AH9	:n��q��x�&R�{6�g�Pe��1h'O���yB-��l�F"§Hk��v�Y��y���
����CE^�U�����T"�(O"�'���d'P|�9QD Y�BdR53} !�d\ql�+�*
6�zQ�7���!�D�?pj���D�%!ފ�#�,I�n�!��?dQɃ���!H�Ȳ
<$/!�D����ꧨ�c(�!�^2OA!�DS�K�$d-�M�y @W/q9��x��8�PJ,+>��6mB�~�(MC";LO��O���Ϭ4��	�Ko���U�2�!���:�L+��D�Mm©U�L�9���3���(%��B��^Eʀ%WoB�8e"ON���O�mNq$��4��+�U�D��'��}h��h���	b�@#�4����N�J��\P���m8",#g��`�V
O����X�J�pT#�*|c�����'�������(P�@c�ġU��@�/1D���*��Q�b'B�My��i�L1D��P4	�wD�݊�C�,/ܼ�C�/D����'Vg (]Y��E2e&���V�,D�x�V!E�H ��A�4���&D� �B�ƨ4�D��K�9H��Ѫ%D���Kр/iv	#ݶj4QY8D���SjG8'H����/ip.=��N4D��	�ǝ(������A�X��(p�L2D�� ����^�`]�v`�<EZ�@��"O��c��I�G��0ȳ��pH�� "O�<�4Ξ�K'4Q�#��]H�)W"Or�i���v��Yu Ǜ	�cg"OFcE!Z=D��ѪQ��=@����'��	V��R�^N�<p�ʚ/��">����,@�ΩÓ�F�6*���� 1%!򤖶y����j�� �З��I�5�S�OJ�U�!+Y	t8\X�' WX��'���4�۳(4bIx6�
x&����'��d�,/KP �5`C0t
�(�'f��k��^E��#�I�4�]���D9�S��I?S�53a"�;\�&]@�㉤�ynI+S� ڳ���jq�a(c!�9���p>!��� /��ZQ�(gT,hǇ1�D5�S�D��O����<�-�fN�I ��8b"OT�2���(Ue�/z8 ��x��$IJ�'�0y3��	��q��߄5u(�')��`�&���P�I+l~��ˌ�;�	V�4MQ�g-,��愙��T�v���yb�6_(�)�����А�H�?�y򋈝f��h �K���ݨe��1�~r�|r[���ʧ#�t!�枹v�0[�͆�npB�ÌK��������#7ޅS&EY�_�`��FLE�p��L��?�"5��"�L��&S�[�� 5Fw��B�	6w�JL
7N��J�����l�=���q\L�q%˞Vg��'ʛ0�ў,G�T�i%��s���a0b�:�뇯I��c�'�4݁cm^��m]`�%C#>]<���2�S��"�# GTQ{E�" ���؃J��y��Y�R��v��%a���� +�5I�v�=qF�i�����C*Q��@��XӬ�V�<I�L�dS@ SUgR*�2]Pր�m�<�ざ)M�<,vL�����a�<����9�4���$8��3.QX�<Y�^7f�였"���	�2�i�<�!C/]�*R�J���H�`}�<)S��>Q� �B�����u@2Hֻ�hO?�I?	>��g*r/�|r1�C�	35�� P�Ž.g�@��^+Pp��P����d�����eN�3}�ak�(��0|��E8I�c�FH�p�F�H�'=�xr�4>�$�JF��5gjmYN��yr)żo� �V�ʥ����A��(O���$�M
,h!�,L2=�7�ޙ3�!�D�>a��hh���9����C-P�!�}���h�Έ-Ҟ��˳z�ay��	,k�A�HZ�PeK���9��"?�q�?�'�X,1&�@�9o�����ڞg�l��3�t%�W��M8��R�;���'��'U�?��WN	L�8����ǻ<�|{&�"D���-X�I�.�� F�[`h�
�%D��� �"���N� Vu[5k%D���t!<;�0g�׺r.�IG�6D��Zud�,gd��k�?n��$�*D�(�ʟ�����)�4d�v�z�C)D�@xOT�\���GK�c�R`j�m%D��4ł�R��`Cg��CNPz�-)D������S�|��ՃS$��ׄ,D�H�bA�f�T@`өT�<(��+D��gO�	�a1�㍣��q�6-D����!~��3��Ԯp�a5D��P��ŉR;�b�C@���%�5D�����gX���6"č'��QCH?D�� .�A�狒d�| �D!ɌP]\�"O��j��%

�u�� �@?rq�f"ODp�M�/"��w�H(78�@�"O�x���58�n�IE�ۄ(0� d"Oޘ C��P��Qǁ5;�U��"O:M�u��\�Psd�E�jH
E�f"O�D*��J5AT�]�׮�f@�q�"O��r�)Ƕe�y@Ӯ�,c6���7"O�\"Trf塡���1!J(J�"O�`�2��0�Y�P,�+T����"O�M�c���*
�u�$�ƈ��"Ofp�fj��D�fa�IH����[!"OF�ҷ�ē�pxPM��Iz���a"O���_9�"��#H8+�.r�BC�<!T�W��|�;`�8_��Щ���t�<)gE]�p��QׁU�t�h�7��l�<i���#Fʨ���'d����o�<�t���f��q��%I:\��)�k�<���34=�� �^�Z���i�<��\ ?�j�8W��:
��Б(�e�<���D%9�|��0E+�� �$[b�<�ԀB7Ɛ3C��&gJ��#a�Ra�<i��޲~T����ޥ0�\�3GOw�<���Q�j���d�D�L����F	p�C�ԋ��3O" ��F X�KyP��<��%�on��r���Ҩ3r�RG�<�"ڮT�Dd�O�B�
���g�H�<���ԫ���c�R�D�Qe�Nm�<��/(<買�*vf��7�j�<�qW=�NpR�h�!u� dV�e�<y���+
�l��-��=o��І�Ay�<Y��٭JA�Xx��4H `2'�^�<�W��mZfL�`ԬH���#�MM�<�A��h�������{��-�AK|�<I�F��&�t�%#�5'T�4k�JQ�<��G\%2[J��S$�6��!�$h�z�<�pSr����R��4��A�l�<	�+ѶtU^12��ߋV�(����Ov�<Aԩ�pv��R��A��b�����q�<���J���\R�M'<:`y�@,�h�<1���G�2X�6���9�D�sq/�i�<)q��d>�M���4X��K��M�<!U�'>Ѩ����ȖAEhȥh�I�<9t�Y]vԑ��_	V �+�H�<A�m��
E��&I�:i�1�eB@�<9ń_4v`�U-��;��[��@�<� R5B6=���1,�j	p�A�<q���U9��u��h^�0� {�<	4��# NPQr�,d�� �l�<1��&<""�E{!ŏ
3��-�ȓ!m,+U��yW$����Y-8�؆ȓ[��iI�/X�O�M�Ŋ��!z ��ȓZ�&���b�v�Jy��ʚ�U����ȓ17B����ȟ��Ia�F�!���ȓ,Φhx2A�'�%JBOQu^؅ȓ88<K���<�)a����ȓ?�Z(�G�����!���]TX9�ȓ?WXa�)T�#���&�LN@|P�ȓ B�L@#gͣ5�=[$��I�6�ȓMc�K�&(1�j@�#���P���u��+��H��ԑ{������6e8�9/l�9!���3.�(ąȓDo�� o�'�i�C�I���ȓa�ڙ��A�w,hDP� �#�܉�ȓ5�5+�M�5`ʈӱ 1bhh��S�? ���iE�;g@�a�m�,= L� �H�p+1��� !���1%�*o��H��G�[��B䉏��U3���"ؠk'ł�,�찠���P^,�O��}��a����*N)S������	[��Ą�3T�A+;�JAz�$�`���l�q$|�1���J��{��I%od&x�!o��D�"�;�%U��=)��tl��:�!�O\��ri�
|
)��|b��U"O 0J��φ����Fŏed�92��٘8M�dX0H�/�h��A�gj�
�)��
ϔz�\$�1"Ojћ����[�b  �ި$� �����>\^�e�U�&}��?�g}B�:,fb4��.��=�p����(�y�FH^������.����Q����M��+0&@�e2|O�|�3��'��X�D_�!$|qF�'����E$D� �b����Љ�KD�X�dq5C@b_�C�ɠa��£m�|�@҅�@�++���7�0@�.�G�D�J�V�.��k2��'H��y�!V� "�pq��e��x�0�Y�y�m�5�* �K�B�>���ߛ��'>�$��&Qv�O�ވ��͕W�n��HN�.h���
�'C����HʾzgP
se���b�J���O��:��Y�|q�K�l���a�mN�(�lp!"#D��;ׅU�8w�<�e*9�2�I�&�rXT�G��Z��|�%ˡ-�FE�T+L�-K�b�ć��0=�Uf zj������,�8_�����˅��c�<D�ԫ��l�4�4ˉ<:�E�S�=�	�8�uɓ�<8+Q?ycC�ނT�(U�%L�`�J��=D�ۅ��9��hhpgF
8P�(f�T3ZD|��a�>�,k�����/dFD3�j:WK
�JE�S�%�!���z�zTc�G�1N!��.�8E��-F6p�~��1�3!��O�.�y>p��i<l��<���8Z�޴x�GI���r�'�ٺ��K�'�Р Q�ÏL����J�.��@��:j]� "ػdH��=!l݌0'�D�5I&>(��I���0s�L�?�0��������G'��,F~���`6�	
.Aj�� W�aK�>)A�@T�H@���艒6���
�A�\XU�td����0As��Oj��Ǫ0IHS�	�'t	H5�҆;��5�R���;�X�g*�cZE��ڢ(G��<��OA���Co%}b��7hBd`Ã�7	���$��,�vć5;4HA��K�uC��Aq�A�iAlp�フ5��O�8`��fC� a�K^�pW*��$F�$RVd�g��IY��xY��ș'�v��nK�z��0$���-pQ���"&*���NƋE�8�iN���`HJ�BR���'H\X��K�����5���a%G.�Z5�ЬB�iMT]z��h����,��.6�(Lc&-Al�<^��B��6؀��Զ�upb	�83D$�j�h��8�K��ğ/O��pR�'d�Tҥ�QF�% 4�����]�T��Y��n�'}���Y��J�X��u+Ŏ\��`�J�'<����ڟ.�B�F?[Z����$�0�@�G�z1�í-M��O�2ǚ�۸��S($2P��>^�n�
@A��J���Gݒ[��Ė�����_r�%��!
<[�|�Z���\��`�!L��u�W�R%8���II�u���`B�q$��?K��]j2�ć�0�� l<�Ð@�CW�ejrї.�� j2������0=Q�bǶ[�T��"�,{�#1+I�b@�@�>,J��2G����D��
�]�
@ã��.y�Ak��-�)���6eX����j���*�U�ay��ˀr:��&��)v�ߢhک�喾Y"5�`�� [s/Ё7�\�2+_
,�����26��SZ�\x�t$��y�`��y�nQ�,p��0F���i^���H,�)����"
��!�>5���E])%ђ��hAK��ӑ�ߝB[܍�mȨ:���d�=>���@�)+�=��n�ֵ��C�~�N�T`�q���M�s�E�"vnu�R9P��w:�"�ժlba�ܹk����&�#)eR���F�5������Y[�uH3/��p@}(��_�,��y��1��*ψp�"��A��4��&_����p�(��Iͧ
@m�t���1g���PH)ι�ȓn�j�R�bR5����$ߍs��<����,Q)JE	%�M�F��P��a�S�Z����.�>y%	_�g@\��sG�"K�6L���[���ae�߹&T���g�=^_�A���$-fxqraT8w��ەE�yl�h�%��4x�i�Oh��+s�ޤz��觋&�i8�aBO���1ZT��u����i�uӱ'�~��*�*"�T��fj1�O����O3K,��� �Q�P����\:� #�ЙR���A�t�y&	ä@��$?%*��T�m�I�٨R�L!F�#D���d�2]� H9��	J���� �^�Os1˵N�#[J���-��	��c>���.?�d#*\u�a�Q�('�b��U��P(<�D��vht��ԈV9b�^���)N�nZuq��G�I�n�3��5�O�ez��#Xh��&��1h,���'Yl�,��&�r}
� a�ӳ&�d�	��6V���B�O�=+��0>Y��6��A6�٤oY��v�,I�C;扷-i�#���w���2H���r�Ai���5D�p
pb¯&��"�G_<D��i*3�3�I:L`
`�d ��^�>�" DJ��P���+�h���#D��X�J�w�)-��P�6��]�z4	,9Ҝh�O��}�M|��:4+:�����ț�<켼��	�"������C���h�H'_��xS�"-��O�@�e
w؞8SA��;!ℨ�p�+-�4d�� �I4]
�
�E]~R/Um�0
5`ʺ��D�(�F�B2OӾ "ɫ�@��<�sLX�Y��)F��?�@�Z4=��{�N]y"��l��,Cf��V�i��@3U���կ�f(h�L�8�!�d,hD��"T
H���P�>1��F���bU��ڤ��̃�Ę�-��$i�ᚌN�ȹv�FN��z��~����'S'b��I߫|�|Ԛb�K�&�jh��P��?�Wo�,*���C�&lO4�PG	!а�@d(��cu�pR���09�@I!ĻX�L�l���1�Bɱ��b�x�(P���G��%���"1�B�I%��H�	/#v�;B��r��}2)�r���
�C#p�g	����@�I�/"t���9H��!VYZ$s#לOH�:@��&ta|R�Հ� ���'f$݉v"�:W
ݛ2�� �3�Ҟn%b�ɳ�Q�,�A!pK�.3f ͹�b��?_c���!�(y�֘�g�͸
*����/�	�V���ɡ�P���ԚrZ((�-��>�i���(~�A�e�L0����L�W�d��BR2`�$�'��ы�O�_q`��!)_i99��j��@�UGf���cђ<����1�U�^ul�ȁi�o6���|��YW� '� ����C2l?�����*D����N+�\mcm��A��I�"��L�n��B�U�5��0t���B%��T��)�D]bÍ������w0��c��L�@$Թr�M"��'FH�{��''Z�l�Hcb$I��N�D�j�c��?� ��Ħ��C�� 4��28�ȣ��?-���`���͉�	AY"@����#7����?i���:#�C��<��M�V���,N�P�h�`�U+$t�0Fl4U�q2G	@'H�"b���=q���	+p�(�J��a8�� z\��V� ��	���!B
�\)���,����GG���2�<��6��-T�&|�f�E�<Y��Ю+�l�I�.MA(�1�BG?i&#U)K�|i*")O��60k��g0V��D�&����V��qa��&|���"r���s:Ĭ��I�bh��a&�3֦� pG�s� .
<�{ulu��ҁrC��'�Zs��P��G�(:�:@�7X�X�s�l0ʓ�@��'�Q��!)E&�Z��4b�"'�u��Sf&x�e�q�<%%��H���0�)P�e\R�(2�6D���7� i#�Ч�řZ�XPie�5D�L��i�*Ұ����S���5g3D���'.��Ua:	RIè�@���2D�(
Ң@�8�P@��)5NdٗI*D��$��7$8<�s�]�4����%�O\��(�H��l�^�aؒ�u��
�'�ڵ�BB�:mٰ�ςB������/b<��I+S���A,�.�>�醤ڔr�C�I<+�py���:*X���Y�RZ����<�A�򍍍y��{>��������4Y��(��D��Ҍ~�[�cZ��S�&a� 
 �˙
�hx�O�&5x	�Am?}��3I`4�R"Z~��1�J�6�$��#��Z�=3׌=ʓr��!�A�*�	9d��x��ST����F#^��0�;�P2V�(�h�OأeA�[5D-��"�[D�G�A >Q���䀟.B�ʁ��������ee�9I}^��&�ǻ@EF|��"OvBB!�T��y����7G>Ax��Oڭ�	�ک)J��s�aZ$1��`�S-,,� ��o�z�L����'M�q�o��<)p�#-(%+4c͹�D�����C�$ƛp1Z�8�)���0<��'����"#�=R��)�#K�Q�'8�[��d�!�^ �D
�s����D�-�n��e��.���3�'�XQP3���ݣ�[<�dx����C�"����>�Ӛ
��z�jM%p�^�Aw!�87D:B��!'��b-ܷr$:���A�@��p�Ι���?�)ʧ9��A�Ғ"*E���*��9D�c��>6 ̓ �`gN4���7D��rTǘ4vE�P��/_;�6`y�I3D����HO���-#+ݢ\e�T�q;D�� 
S)��
�B�L�2)z ��"O�A��F�q�� ���3)"(�"O̠1c I�DO:l�� -x�v�Y�"O��  ��:u�񯃂i��=�"O
�6NF)y:Ĩ{�#I?5b�h3"O�@��D��v�E g �z i"O�}���?.�V��!+���"O$5K�e�[Jt0���o�9�3"O�0[�IDD�h��#.&����"O�\���WX��i�F�H1���{�"OҜyv �5R�RYu.�{�ZQ��"O i�C�n~0,�n�)b��͸�"O�dB�Ɋ"�lݡ��8%U@�"O���$'A��/aCf���"O"�q�NUH�x��c�۲h�F`8�"O��$"�R��m��m׫=��I�"O��qB�#<�LdK�f�>v���"O �A�"�~�c]����"O�� oO+J��ґ�D&QӘ5�C"O��Yw�5O�X����;n�$ha�"O0�qdԺo]�u�0�v��"O�Yʴ�N�m��i!g�;�X�A@"O�` S��I��8���N�%��ź�"O0�+�����;�!@P� IE"O��sG&=��[�S�V�@|)�"O \Y�#�=OX�Iģ�cߢ��"O�9#���y���Q�a����"O�� u�/���vb��v���q�"OZ��ƛ�LVFQ��H)�*�B"O\�����8:�B���� O`>��3"O�u��B�~�td+@-PW��I�"O�5�B�Ç3�>�� lH�(]p�Q"O(� �+R%heB�%��9c����"On�aF�K�Pj@x�TJ�3�lͣ�"O���l�=>�у�����"OX�ۣ��"��Ā��B�z�%"O0��*b�`��<�C"O�Qr�e?F�Ddq�"�����j�"O��ǣV�/��G��f�4@��"O ,Ȁ�C?{���S�\.o�"�"O�16#dY��E��;��qB�"O�t!T@Z�m�8!{�g�kQf��"O�z��!IzZp ���_���u"O(]���ޣT��B��_5mE@@#�"O. y��Q���5��cU"OnX$D�~��XB���]g2�ڰ"O�mDC#%�H�hGLȗE����"O�ē@-�0X���& �<:ѐhЦ"O�`��#Gk�y"u&͖Rd��p"O��0D�\��pQq�K�!J�p�'�,]y�M��g��AB��(0�v�j	�'d2՘�H��ؒҳ:Q���'��=i�n�)Z�°�Ր6f��'�V�c��2MƖ�i@K1]���{�'f�����`�d��d��gͲ�
�'����%��>��ᛓ�\�H�\	�''r��50C<iz�
��FV��;�'BV�Ӈ� 3���b���h���
�'��y�G�T�*��!�P�Ģe��9`�'� ��A�8K��؀G��P�:�'j�Չ�A�I�l��Gh���`��'��X�r�Q4>�ы�f��A3��)�''8hqA%ßj�D�1��˙���)�'p������h$k'�������
��� J����_K���QM�m��(+�"O������%5И�1K�%'��X�"O*Y;�CÐh?����������"O��U�&)L
0��p���"OA�nцv��\�bZ�(���d���>����!P�%M$(�6�ވb�B�	�?��������R�ޭ]Z�����H,r)4�O��}�WF̓���>�Vx�6��m2|p��/}�Y(�BŔ~��*�K@����m�	@��b��"XG�{<	0�b6b�Ry��ZG�����=� j�1]�v�����O��Q�(-�VQ�BH�|k�5�W"Ohr#�#�T]�EGH�f��{��$�,=����L5�h�X���iN2m�TX0 �N��kU"ON��a�1� { iE����d�ş1��I3�(}b)$�g}�̆/kި�vh�!�����F԰�yb�!.tJ�Ќ̚y���M;��AD�J=�a�9|O�ܛ�HVP�4� SH��v���g�'f U��N�"R��(�ɮ	� 9��!V��a@�Y>��B�I�o��Ā���+Mʨ��w�⟐�.B۴�E��c;"���8p)S� \N��DHT#�yb���C���P�1Q<�D3�B��y�H�%p��tDo؃z�AT����'zݰD�Hb�Of@��ޢ������PѠ
�'�.��T�P$~�W�ʅg�x�5NH�ȒOpٍ�Y�(��.�!����A�����23B D��чI�B�,�T��5~j�!��^x��
:@�|r��=O*~M���t�͙5��0=�DW8d���*2��t���4IΎ]��+]�Y;6�:D�`�b��-et����"fUyJ6手%re�
ׇ.�Q?]"s(@�*� P�v
	)Gp�uY`k4D��eO�1v�����JzX,K��ճX��08C�>I�]i�����Zm��	�-�dMZ)I�n[&8�!���f��YJ�	ʙ;P�c�M:,��P�I��b���i���#l�i�fh2Om~�SG��?/�x������?�����'�qY�c�O�'�vТAM��:�����.9�qxG��'>(X6)C:Z�AExR�*Xx`ˠ.5N�,R>q�����O�\궈e����6cקb�~���y��g�f���I@e�O�U��*ɃM�n�ơQ��h1#oЄn��$�dmX���0�M��
)��ټ�q��>�ċA#�/M"�����,͌ȳA-}���6���I%d(�	����Z"m�P��6\� U`S�v��5`S�	pyӅJ�,�9'�A���' y�KSwL����ǶWq���A�]�:�A��o�'>R�6�Ͻ'�$x����)��*G���
��ѵ&�<�V��bO��w����@ �X�� 03��Ͷ��dK�k˼!��?��L0wD�-gU�O���E,�ݎEC��1~�}��nI�]Ĥx9Xw^�4Zq���D���A�$�X�H�}"Ɇ;W&�|E�4FH��p��0N�'30��2A�.$f��zю<�Q
S��-!~�2���-�t�>)�;B�%)uO��yQ�4E`�,c�BB�	�+x���ˑ���k�&ޱw�&��Ҁ���$)P�Cc�k�-�|��`�J���'�R�wgM���UCGg�|2�l�ߓtv��W�H7�\�+�K<da4.�*�DU!�I�}�P�+��"g���a{B F�BN�z�f
�i�xx���O�4P�- �H�2�Z��`�@Ѡ��
�I����xqхԟ�rH����4+!��� {lV��P�-�����Ǣ\s���&E�
W*t�"(Q�9�~(��M zmQ>���R���Bc��:Pw�y���6y!�dX�0��A���2Z�H):�.X	U
�m�O��b�@ܲ���qO�:�:DǄ�
�O�:^6�q���'��jǮ�;zB�O1u�@���'_�R9�ӇDo؟#��U�!��9s��&g�:��4�W���gM����­�g��!2�z#A��'�)�g"O]���F�,�|����C�2'��q%Y���k�	iހ>E��m�VO���Ee��}��]����y"�+ڸ��J��l���+�d�'34���@�S �ϸ'>*�IG��	8 Qp�$�0(?�%"��< �qs^*,O�-�ǁ� x�rd�ۊ���K��?���d�Xa�%�+yH���'� �BH-�X�'��R�f^�/B`(�k� iQ�9D�� ��*�E��^���3��B	-��	��>�G��X��?q��e�h�d��T��/ ��  $%D��!��JN��@J�7���B��$D��x3��nT�P"�m� /��zs�&D�Q��l�q�v�?;0��&,��dSG̓��a|��ؠ�A&���,��.ר�0>�FIL.r�N��8��� �L
_��Ȱ�%/�J���{>d�0�C�G���'�"�e�?Y��#�rИA'ҧ{N�Mr���j�r�ZW��X��ȓ�f��U�0|��0bݞ�nIJ�kG�ZO��g�>����O ���ߤQ(x�JR�!y\Hq�'$4$���t}�i\�,��d���R�[ �a�B���?ٲ�(4̓U�:lO�a@V�A%*���
խAK
y���DP�@��<�g $?a�
V�#�$ui��`ݹH��A�mM����F'Y>� �/#D���%I��	s�ĐX��A�^�I�$��<q!�'��;	2�針�yW��d<̲ KI?Rq���R�y�x�\Eh��)'����`J%h����Մ@Rƈb*O,����)RY	�}B�����O�(��ċ0�p=AVA�L�j,�r��-�Mk�IpZYb�@ʟ]��H�m�����PgU�e
���u�'Ab���]�y����ڝȍ{�JH>z�P�ZbK\�zG�	.UC��C7b�?��� ��`�Bݑr���ವ�j7D���#k��~�P�%m%p��D�;����͐��?�vB�L���C��~�@%ȹ?q�?�h��ï��N�lL��莌l�>9#�'v`t��i�	�r�̖
w���c����0�s�Qq��\�Pg[>;�ly
��
�=FU8w�̗	�Ń[��O�����D
FL���Phh�� �k�q�'�S	�?�Ņ��&�0�&\4}q4�����N4�<чK�.T4D@`θ�b}��c�{���RۓA��-����H�vL�1?�m:$�] Tq�@a00O��3a��D��B�
�`��ʲ8�y2d��b�e�]�b��ӓ�N�^�~�[g"O걸hJ�~�mk� gc]��*�=�q���<h��TC�&���э�n#��v�A���w�F��2�2yG��x6��j��H��'�м��ȉ:\L�o�� ��D`4�ˉa��%i%�Q"3:R�k@J�A-��X��X�U61
��?9:��Er�G5(%�@�Y�f=
�����#MQz �?i����rxrB��<�@G'+: �ai�<�Ly�sFů/���ba�`��+�O��>kL̚2�Q?��=ѷ-��y��Y��m���yZ���>�� �	�k����y�s��d�iۀ�D v��s��_�c��^���'%ѝr4�x���F�<a�ED�D���(��;`)bV��B?ᶇ�k���a��2B,�B�U�oy\��&h���*l#t7m�� ��r ɇW��I�L4��¨@��D��\�>9�ݰ6�(c:(x���Z�¡��#�My�������ɜO��;�	�%�����!܀H�H�<���D�N�"~J�� �c>����/<iT����\�d

8+�#I��	�"m|�q�+U���5�ʎf?^B䉰-��=���MK�@���3�*B�Iu�<�QwƠ����2Ʌie:B�ɇI\~�*��D MUV��䃝V�C�	�	h���/@a����8dP�C�	�~{��:�Љ>>ѹ��^�4�p��$��y��!2H�7V,�A�#E-f��z�fI���xb �� 8� K�"��p
���O&�XW���[8�>ݸ��V�72�{#;2xl�P�%D���Go^��;U�T�ND�������׬(yg��f�>E�4�@/U-�Z7fR4L��F �y��U*
.�*�۟QZ���2"���=��CUe�)F�axl"!��	���_�N�Ā�h��p?	 �ײ����2�ݡ��HŊU#u.rPQA��/�C�	.g���2CA��r4p����Z혢>aVLʼ/<,bpj'擢:UR���(�KdYՆ�W$�C�I*s
�r5�2V�c�e�b]��	+C����h޲/��S�O%��;��ܹI�P5��@�	�:̈́�Hq4�"FNW� ��yǈ�;��x�O&�sΐ	r�q�
�HV�����2X�&)�Q���$H�4��I�ƈx�JO�6/�����&=�	�C&�C��)�@��E�+��A�Ęx� ����O��Y� ��0��>1���#+�8�kج8�My�l"D��P�ܙ;�h�V�D���DK3o�<9���4➢|� `�@�EI�M
���2��joL�B�"On���&0zT�8�)*+�q�"O~�j�ރ.�8 �0��O���Y�"O���a@ݬpz�y"��Y�%p!"O�-���1_ʕȲi�HI�` "O�1@��]�T��iD=un؀�"O��知&�B�+2���LG�((�"O���w%R�r]0���ۄS醰�"O�ѣ(��3e�y6�����"Ona�`��f�\9ԧ��h�As"O�	��
[P��7��(�r�6"Ox��
3�(��d_"�2���"OR�+2�в."�X1G"�L8f��w"O�I#�]�=�8c5KB3A.X��"O�Pg����Ѡ�+݄(�d��"O��$�X�~0��ϓ�9�t9�"Op@���+��"R��#�T;"O	�� rA��+�O�ru4,[�"O� #C�K�M����1+U$`o���'�y����l�h�����**ze��'������>Z�A�L�2 ���'edlp#'Ѩ" �X��b�$����'�|�ؗHǺ�r�������'�<h��ߕg@"4jr�B�ﴼ �''y+c۽Qa���|[z,R
�'{,1' F�}����o6c��x	�'pU���*�����C�P����	�'�b�� �>�����,G�J����	�'�d�rU�I�G��xH�a��T�X�:	�'p�]�j��j��T�qE�{*���'`*����	T��A�W(֨p�����'|�r'�#� ��fZ�>vh���yR��9yv���!F�'x|�Ir�Ë��'�|]����!d�X!Эܟ��B�'6�@���
�L1W�OO2xy�'�:M�ՅT%��t��G�{|�
�'�r�p��]q�(V%\�!(  �L���'B�*ç��q��-N@�����s<���qm����DV�z[e����0|JGA�>z]���OԐ7x�U��E2t�$��o�F	q��%{�X ��ӷi��i��I�`�$�P�T��74 L�5a��`���
w>y㇩Gl���BBN�8���jϧ0|�r�f�(&p�?O��𩉑R�J0卍�pF��U	�|�!����S����'at@��'K�B�kU#Źq>�1JB��,⾈�T�=V4P�Y�y�'M1�,�r�I�$$Lp�kB~���>��L��&���ç1�Zi�c�-�e:E�S�s��'�N C��T�OH�A�OQ>A9 E7��I"lQm�DHT��Ovt�L�$���N�"~ґ� Hl�bt�Ӫ:�n4��� �~�@V#{��O�>)p��͞	N �̏�SŜ���"0D��U
��W��DJdk&o|Z�0�),D���a��s88��,� 2�T���,��9�O΍Jt#�uX48#�Or�(Y"Oh1� ǒ�c����P��`<�\C�"O��!ѧ8�r� [$)��"O�,Y��#��0x�.��)�c"O�yؖ�V����I6/͙X�P4;c"O�qy���$	��1z�oU�$}�9p�"OD���(4�QA� s�慲%"OI"I�b�6գ�FA�2Y$T�""O���R� ?�i9��UL0@�"O��9j��(@�\3�钾�Vh"�"O���J�=@�@�*��H��!;�"O"���,:�H#�ְ~:��"O��كa�/]���k\�T�I�c"O@��#Ƨe��+$G�l)7"O�dÖ2R���
�K;*�\4�0"O� ��h�f�	w��5*,���SQ"O��ТmV���� �4+N���'��`�U˘!�HEK�*��V�0��'b*�QC�ؓI��J �]99���+	�'f�qI1/Ūo�^d��'��*��H�'dr���˃2�v�QG��� p���	�'�,�{���~M�V ͉�hH	�'�Ԡ"��_�6=����^�p��'����.�2��qa�R���b�'r�-Õ떖���a�gT�{�x
�'����a(:�ШA)�!E5�h�'����AJ�%\����B�x��'�2�qB�D81���W� .��i�
�'�8R7`��|:ta���B'6��
�'�.�KNw�Υ��R����	�'_�MeO^��
��4�Љl͈	�'=8��'�s�,,��jû	1��	�'S��1��S4P r�h4�H���E�<ya+ʯF�xؑ �Y�	 ��A�<�!�̋|h�"	K�vl9֌�a�<A�cѪD B��t�<X#�	S�<���
^2$e!f��SA��)$i�R�<A$b�1}�p�Y$��=k��	ɐ�
K�<�7���R��$��=B<���jn�<q�틧W��+��F�����֣�j�<ys�z�(���4�]�Cg�<���U�uHb��F@��T �)�Yz�<a S��j=�T`E&jBz��&)Zy�<Ia��LU�U�A	r2yy�B@~�<����,�t,Y1倠Ip4ab��`�<�#K�r<9�4#�����x��B�<��m�!d��%�����-�<�@���A�<�d2&���Rd֋P��Ի`�KB�<A��T 0�L��'� ��$�E&�A�<!E� �C$,JJ�Z�XԈ.s�<�D�$��<cS��(G���!O�k�<�s�;�R,���X��P;'Jq�<yaEЧ!'� Q�៮#4F�q݌�y�f��dln��ۡU�>%�5G��y��8(��"�(H��@�� ��y��IԔH���/���4��.�y��O3{���b��V����œ��yB(�4M��T�-�Q�$&��y���y� X�4�	
Of���I�1�yB' $p�qqv� �FĐ��$����y�BK�u��!���&D�r��4�G��yrL	�%A	��Ά��<ei#d��y�-�Ȕ�A^)1g�c�@T:�y2oIB�e�E��&��(�;�yr��??�:�`�G��ʝ�t�6�y��A<,��(w�ψaݸ	r�Ǘ��y�+F���u�^RൃƬ�y�Í2�H�!�ō�X��e��U��y�Ƈ��t���M�N��i���;�yҥ^(>���6�ƩE���2��ʙ�y�ˋ�.mx�a@�=� �`�M�y�HN/Q�܍򔫛5��!���y��Ȃ ���R��۪.Vr�J!H>�y��ެ_Gt��`�'tܹY�X#�y2A_�g����-W��P���_��y�Cϭw�DӞO�x��$.�y�/�4�P�1�/M�6�уSJ��y�%�f���S@�5�~�p㮁
�y��+lk�}�@�1x���G%�y
� lԣ�f�(I�AӥDG	=I��y�"O<�*у�I�RՀ"Wg�B<�"OmѤ%�c���� �$�,�q"O��dd�!u]T��� S�" �sE"O��؆�j<P:��CF�:�R2"Oqg��-����S;)5�1
�"Ox�B���A()���>C�lj"O}	0dHi/vY�m�73X���"O�)b7㊄��y�D��i"O2L#2B��`j�KWP��e:'*Or�7T	A��)r���B��\��'g�������d�$9d&���'�.i��B�2�H��[�5%�8��'�p$ٖ��Sw��k�名.�*�Z�'dH �I�-J��ٴ�hh��'��xX�,�6x{U&�r�d �'�����Fڷ"ۮ���d�'xj$��'�j�0!�Y�`����	K"oݲ|��'�hpQ4g��x��9z�g�b�H���'��(e'��5�N�P�T�٫�'-�!���< �z�����)N�j�0�'��a�I��_�n��G�څ�حr�'v��Ko_*'��h��(� cz��[
�'�ެ[��؛b�J�	@�l�:��
�'��3��J�H!�D��f�p9��--��e�I�b���y�M��k��Y�ȓ/���(Y3V�҉�@ �1l��Ʉȓj��7�]�L^FX��*-l�<���	�zse�sO�m��F��@H\��*�#0N���@� �) 2L��ȓ=H��)�㚏i
�1�k+��X�ȓI@��b�X�m2�J�A$f��ȓ(V��j��BO7�a�i��;G���W�>4zՏ�yt����B ]��	�ȓ|�Ja�4�R�a����U*�L��{U�9�B�S�EH
,�ք�"|��Q��\�n�a%���G3Ry��g�(��ȓi��D:`+�{�t�!@+���B����ii�N>�x谤�>h]�B�>� �!�,�0~w��9t���?z.B�Ƀe"ةQ!cG+\�h�g�&d�2B�	!Fn�2����ZI����^�"B�I� ��S�o�'q{�=sqnԧ6ưC�I)O���2�F�(d�����P�S�xC�	��k��[8��dZ֥�$0vC�
"٠Ĺ!�9���Kf�ק-:C�ɍ
C(�xbh��{^T�3�c�RsC�<!��8���9o�D��U�Q @�C�I�Hb�@���)d���j�	>��B�2^T�}�o�	�ƫD��zB�I�9���+�+��7�ޘQ�� -{n�C�I�#nĔaT�޲���2Ѝ��F��C䉢&�ta�D�\���]--JB�4��	3F�=J��$)��M�C��%P!�\���}$��H�$��(��C�I�}Ռћ,��!Q|�C�?msJB�ɑ6����29�PX��	KR*B䉑<UT�ի��9�(S��L�0<�C�	f���3��<Ϛ1�.�C�I�-�x��qbߖM����Dd�lIa"ODcg��%z�(�����AO��y�#�5f�u�� Z +�U�2
��yfӪ�����FK�x�x�81���y�#�9<fT�H�G.wZ=kʖ2�y
� 㕥̯[�D�ьPb�I"O�� ��^�_1�[�( 6��:1"OҜ27B
u̓���=)�@��"OhT4o��>\l%i���o�
��T"O"�&�\�<�DHA��4���q�"O����c���p���%=�ֈ��"O��'�m��tǅ�4XH�"O�pѪ�>0�5�QF̝Vx.P�3"O�x;vC�<��D�0w@��f"Oȸ(Mɤ!Rb�Q�FŉE<	�"O�u@����dAhkP��x�"Oh�{�b���X ��BI����"O����Cp��X����'H8V)	"O�)���!� ����l1��SU"O %)C�-n��PE> &�y�"O8l���^ l��� �h�*��Ђ�"O�i3t�>I���1��*,�J	�'�+1iZ/A
� �æp���`�'��@��dӧ>=`�ʧ+X�~ɣ�'ن5����;�)T#�Y��'� ���U��=�@!���� �'}��k�G�20�BS�Ł^�*�'��� �ei���3���	z�s�'�E���<n.�҅��6{:=��#܂D���.i�@��
�)&@@��ȓ^��q�e��f�4���@st��ȓB9���S#��`�:��J�KJh-��Az�����0���d� �ȓ=��@����<H�獁�P� T������������V!WN;f݄ȓ\T�2� v�x :$D��1��,��,�*���t���Uͭ}-���vx��U�M�5����	U�g����ȓ,3��.�99G���$�x�� ş@�<9EA���pXV�*Q2XW`~�<9 j�;�b�3Θ��x�[�c�t�<�'��:=f�*�%F0uY.�C��F�<�*�)<��Q��-
4�8xD�B�<I�hU
[�\@�AY�f2hPi�dK@�<��~� ����W�
��rϋ@�<aR�ԿjT��Cև}ºm)A�He�<�c�¦*Y�����i��)��,j�<�0�
pHr� �/@��4+^�<�+Q'|�\ 0�I�D:z�+��V�<�q�X�]�d$�J��HP�#Ff
V�<�6�jo����M��k��Z�<ᶋޫ��)�N�'q��D{�j�z�<Ƅ�F�@A)%_%4[�#���x�<�b�Ό	�T׏��Z8�t-Xw�<9�M��1Y,jᔄ�Rp�<!f�8^���J��	 �����Vl�<Y��AS���Ǧck��M�d�<y�#�N:���-´e��y[���U�<�P��Jv0@C"��	E�%3w˒O�<���C#�T9�6S�h��)�ĥMH�<�V��p�lxW�5�t$��F�<Iu�6�(��"B�'���c�[�<�e��o�&\)v�� ��}I��	Z�<!�_�Nj��V�
�"�e��&V�<1���H�Z@A�Z�.�B�O�<���ս8]��ȕ@S�Kᄄ{��M�<i�    �