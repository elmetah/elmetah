MPQ    4�    h�  h                                                                                 [C=G��Iq������n�_�CB�g}o�������=Q�u��h���O�u��ӱ��R&�?Yj������҈lG��hԺ_�׳�"ڰ�M�4���������S?}�_���S��~�f����q(WHq9Z̛�KH2[�����
���ץkU*(��fJ1�^c73�z��W-�d�S�A��Ć��:�/�6`��U�R`�}ݏ�$Xt��ָا��]ݚf= � ���������s����T%�����v�c�.AB��9/D[�u�.�8��Et��q��jo"�Q*��[r`�%�Oh��F]%&a@Ǥ1�%oaV�v�W\:#ђ[�F<���>�~���u�s;���W�V�;p3{c�����xE�ُ�a�GT�9)��cM*8�k'�ĳ�$	��Y���S\��.�JJݶ�x�+k3P*?� ��
+7�|�اn�sN��v�.�Y�֣m��Aɉ�&g\���F�ĵ�sNC@��+I]E�Օ��w
�2�@egw0K�H�ӎ��CBm�P��jc|������ɘ?V�V�X�����(1r�iM�u��?� ^�ϒ\و�hl��P�'^י5n��٘PO�_ݢ�a^�K�!���>��Ϣ��(7E
�X:�(T�#;ó����b��)��dŎ
GJy�yi�2��x�'�D�.�0j�����z�%�'��5z|Ƕ(��e�e�l����sW���0��,�`���Fy�O�q�.�vr}f0� "Z3Qe��?;�k�݉�	���S�և�ԏ��]y���^!_R&V�>=�G[�ı�w�$�#�5����7qs�=}Q7��I�߼kI��>^��B�)i��'/��m�a/�_�!/p~d
_�;�KE5�)�5��*�}f�[��e3j�kU�hͼN��=/t�:�K���)|�7!�QoC$2���3��uDm��~�W'��9�y�:rH�K�7�ʷ�a�:9pί#���>�
��	�C;�4�]�B��Ij�M��#�>������)��ѝm�,{و�w=�3/���q�=�z<� ��!7�Dm�'i�wȇ�Q�S I�Md�5��F�)q�}B����ǌ�&��� ���c�}F���y�	��-O_��=.Oԝ�����|�jf�.�*�ԴlE����f_�$���p��Q��՘��"_-��U�� h���d�@\�dɱz��u����Ӥ�eYZ6�����P's���|���� �T$��y�¿zlܪ���@7��Ҋ�&��'�u}0j���9���-p-c@]�<"�Q�0 i�߱�uG����v�&2G!�a�R<�]P��Y���E�,j ��00�(S��cm86��vb��(�h9M-sKkp�C�"l�1�59+�y�z�bm�aL�Y}� {⃓N	�
`O�9(D ��t���gqTʗ�'�o�A�E)OE��n��˽:�QLv/��%��gC#��{0?C���$�����?
[�C79�b�1�S�Q�&����UdD��|gfI!Ֆ�1�FX��G�e����F8�Y��(
�P$NT����Y;�90SF�q��c%���>�z3��>"f	��d+ �v��l(��--�뷇>??��Z!�O2��WQ0�nsbV�}?���ﮗ��`�&��q�l-��8+d�����s���Ɯ��(�Q���m�ҡ�b�������2_�V�(�����+h֘�/��U��7�w�mo+��0��l*�<]�k?����e��x�|
t$?Q�y,^�Og��쪔�=����D�jϙG��7�#�����ѷ�Gd�#��,���-Y�R�#P�GR "��7����
�>��۷��=m@UP�V�L�Y�Ӗ�������h"[�fx�BT�q��T��uǱ�k���Z<!J��e�%�����ng}צ��-�r�昮7۬]�J-{U`��Q�^;�(��$*�r�5b�q�T�iT>͋���^�P����I�2�{�kF�������S��T����ݒ �U��Y���J�*s����5�ڨS��M�+{D�V�M  ���FOk�&I&�KA���c��6�fB��Z�!s�6�p��w-c�Y�t,�H�h�<�W�Օ�;8�-W�[��oH"�w+^ّ��ը+�:Mcq�.�Wˆ�7?5�OI�C|B!ө�=�;��(Q�F����ʯ�_�2O���1�c4��ߕ@ I/�N��M�#e��=�#��eo66DS��Ӡ��D;�L�`�a�[�h��st������p�+B�d3��ͨ碧���b�5oV�s'�%	�$O����7�8e�������29��4�P���lL�԰c%uqs���5��^��:�D'Ƀi��E��{�z�ǩ��GU�-���%�OUt@P��k{U߰��=fӱ�ҙ&W�s�5���O���8�����rZM�`���\D�8˖�1�	����K��t��1�0R�H�r!.\�{ׄ�5��|gL� ,�c����x/s��2�/B5�o怾|הm����v8�ج�%��08�q$4�ө�(\Ɂ֌~yK���tVTn�-�*�1Y�7�j���nJ��C�$�̋�ن���jr��pIe����hZ�H[����E��c����F�d���o;�<���{�n�Y��>Q��Ws߄�F�)K{��1��|ρ��`�i+=���x�~�g�Z���du=�Y\�8a2�C]n~���~;M�s�H$�'膕��i�Sd�Y1��)3EEKR�g��/��	F����[_Z)EA` d�O�Pg��?8���$������
Mp�F�i�:G�3�TK:z*�=m���6�O��+��	m1��#�%��X�Ⲕ7������f7\�|�%��'��(:J�F��u��$핼�����e��=Z�j���]��#��(�~|��6��&�w��X�Y��:u��O�@�6�.�-e��W�3�f ��D���� N��{|M��š��g�����`�<`o��p@Ð0��M�]�ѥp�5l���y�N1��1������$b΁��a�/-���w�L�.�a\��u���%ǹM�%������?#>�ry�ᜑ}�A���)|��;5-H��D���;�ӑK�Љb� �m��~
�:w�i%�l̔���h����4�
���������Z:u���k:j��\����U*sw����q� z�V�W�\�iP�#a�΃&V "�(�yA�2�߲<���,!y�n��S����wM5�Օ�M�6d�X�dB^��~C�-zU�KY��'���eF��(���j�c��VA]4�9�;[��.�X����n� '��o��kQEfa��7c`�U�O�ѭ��}%!Gs���U��V ߔ��#�mX[�|��:�)�y37���;���rJmZ�P3V���¡�5��֏X]@Gb�)�O̼�N+8�M�'������T����D�i��.�s��1���G�3�����^J�=k�� ��$��b]�D	|?��j�{Ʉa�g�=4IN�'�9��0G�q$�f��]�.ՐdXwe�������~��u&�i�~I��m$Є����|�f�|9"ɳ������J
�'�(r;T5�p��?���;�٣X*lvJ��Y��Ԡ�5	g�ԡ%O$�S�����fkÍ	��ԭ[��E���X5��T�v��n_)���ޙ�n�����E�RJ��ydZ��'���T�(�fD&����Jh�:N� L'�Iz7TP�C�Qe��v�Gkڻ�-b.�!0�C),�H�h.Jy�qi㈓Q�fk��"��<Q`���?��&y���I�N���.�e�Ȥ�r�C]tq���K�R��!�(kR=ل[¤��������9C��sj>QR��IA��k$�>��D�ݲ�)d7ǂ����SaJ�L�}��pY�D_N�c�5�3�אY�*���fJ5���3E�k����W҄�8&��qpKt'W)���!!N�C��;φ��΃�p��	��W��9���̵H�H���7�����#\4��oO�MFS>
3������[Cv���Y������1#��6�]��t����ǪǪ�ك�w�H]/L�@�
Ѥ�d� �&�r�mM��eR�V��y��Ű�I�b)d��}�G���D�������8$\����O��RRt�ȿ�����O/�t� C�8� |=t�	X�	AE����_ES;���z��ʝP����B��Y��UR3ch���d.�j��袱������˿b����GZ�Z7�ý'�!��7����XT�.�T翵v��ĕ�s�7<�抪���=u�eœ����W>�-�1@X_=<}m��%Ӊ������-��q`v��C2��a�tbU��
<��7,���k��c�P�o��mI*;�b�e�-�M���kKj��]�d�4��]�4�agc�Y�)�{��NT��
���9#��#�ۏC��qo��EDm��o�����E�l�A}i:f.nvJ+%`�sC��{{k+ݔ��6u�2[W�[9��Z1W�S��&�e#�@�_LT�ڃgg�X�I<WܬXe(	G�=�Y�3�ӿP[�P�^No�/�2�!S��ڵe�����ę'}3�#YBu	 �W+�v��'[r�D��T6����?o�![��Ɓ0Ь��O�}�����#�gI��A4&�������{o�+�� �>x�������]�4���|�?r��e֝-��u���B_`��R���%����Cm�j��Uc?�r�9o����;�4��#ǭ����F)/ūNeНx��,t���4w��j	1�g���I��uvj�;<�B��7/�I�͹��0mdT�����@:-�-_�FG���=t�����	ܣ����#�=N<P��L�9�������;����C����FB� q�G��r�l!
����<�[��@��C��R�}��x�crG�3�R�]o��{�@�(����(ҧ$�5����q�x�i�啋vK�^/�*8LzIܨ��N�&^I����,���˖Jy��-E[U�D���@JY�%����5W�S����f���* �B�)�kZT8IA��AM�c��6��c�U�!n
�˨�w��Y�D�����h^�W�sH�֝�-R�.�Q�~"s�(^�L7G�+�(Nc��M��z�2#�Ԫ��C�J�!�OlW�0;�=�c|������yS��aLO��1����c�@�C�/��Ս���q��n'��J�6Q�*�>�g���;������V�H�IX]Fj���^$��?͵�~D�Bb��]�o��<'�z	�v��X��|?�e@� ��bw�l�Ҿ`��Y�>Mpۯ�P�u�m�������d��J��_O�������E����z�����SEG�{y�]K���b�t��g�F�W���4=�\���6W>;�����"M��F�"�����M%��`���\���Q��$�'�^XY����l�R/�m����?����P�Lsx����׷����y����/�qc�*�����smVrˋ�h���j%F�?8��4V;��㮬��6�y�n��O�n*f(*�N,Y*�����)(��e$3���έ��L�le��)��Zl�ʖEnM�cЦ0����n��6�dw�{}bY�];Q6p�s�"�F����1�����.k�diF�����xw�g-��sPp=����rv�2�MIn�'j�#�;�@�s��$՟b5聿���҅S7%1��U)��HK-6���ڞ�t	A����_IKA{.���PB,?S�I�T�ק��t
�F&�z����ϮKu
í���ը3���+�ā	�	D.��#��k�����/���G�"�7oT��[����(���@�u=���b�h;8�a�� ��� ��8�4#�i�U�1S��J�{���t�vٵ��*i�q��Ȩ���eWQʨ!n�������T �����M.�~Ŝb�g�a��è��W䀥x��k'[��n�]b��p�`�l`�W�4k/�i}��E��ӵ�:�W�fbi9�\�>/���2�`�IP�\jb����8��58%'�ȝ��?~�p�-�U����}]*ᛦ!����5�_H_�DGb����ӑf�Ӊ���HLD~Eޢ:��i ��d��LW硞�K4Z�����f�:�&�'��u�I7/�j�����OU��&s�o����J� u�c6F͋�[ikyGa} q��
V;A7ËA���V��nq=y�JeR�㈰@Qw�_^�0��M��m��B��~^��-���K4�H�bJ��lB��X�,�bc�(�Ax�9%	[���.9��{��[��\No��XQ`��Qx `��&O�c�A�v%M��Z�E�0�Vg�MS�#�h[�x����t~�+�5;l�������=31�p?~W�<i>����x�G��v)ͭͼYpX8��]'<}��Z�O�O5��	���$��.�@ݬa=��Bs3���F�N� o��2r`N�S�U��B�"�L����V�^g��vB�E�i3��ô��C2]{cՋ,�w�i�ʶ���$Y��b�D�D�Sm�o���p@|A�E�7w���	X�L����bOtr�^��kB�?y;��Eپ8�l�Y0�ˬ2�Om5�ܠ����O�I�P�Xށ6m��������I{tE@�}X0�TX��)>r���C���a�ꎀkJ��Vy_��4!Ϗ+��CIAD�z?���%��7���y���'FW=z�H��^�]e���"j��aɶ�0ԘG,w�1�#�Qy0q�=o�,��f�t�"�, Q[���^^ͧჳ�Ы��.(�	+%�����+]o\����R�ao�C�R=|Ɏ[����`�Y{���P�fs%_Qm� I�6Yk���>��x��)_�R��O/;�Sae�A��Vp4�_��ѽN��5�I��$�*N�,f0X�gM3 �k˰<��uL�3=����K/�t)���!�jMC�it
���i��k���d��W�'P9���0�|Hg�	7*����/��ʛ��>%V�O����C����>`��=�{�#A�����q/�M��GV�b��~O�w���/����,�p�� �~��[�m�|��s����@���'"N�+��=,��}<m����B���Z��S�\�s�*�� ƍ���cP���eO��	y�|�SJ�|�����w5�J}�EA҂�t_�����H�&�[��a���F��{U�h�d�Y�|�`�����kX�˚���MoZl,P���:')������/fT�/]��l�5w��C�7�`�e|;�3,�us�̓{��˒��-�\�@S��<�g���k���8�kh���!�v1]�2}&Ga���χ��t�E���z,`�����|�����
?�mz�g�b?c%�H��M#��k&pͣ�εgM�/�/�߃��a�!Ys��{��PN��>
��9���~���*�q�6����K�oT���{�:E����N�:!+tve��%��Cٮ�{���/]����[3�9�@�1��VS���&�Ro��PZtP�5��g�k8IW���'��X@�4G6����z.|	����l�N����*��)XS���� ��A�����3TL�t�l	�*7+�)��bi0�߸4�ݰ��<V?*5X!,�ش�T�0�
��hf}u/���w�������^&��-�b���Vx(+��q��#'����c����j��}Tẖ�k��\���酮_���a����o�t1�� EU��n�m:�o�3"���=����2aP�!3� ��e��>x�\�t�N�������\��0�����V�1jI�a�=y7�X#�u�����Zd�����Y��{��-��C�\�G�����(���
�����W�-��=�{P��_LY:V�I��ޑ�سnj��:�B��+q��a�'�L��h]<�߸SȧY��(V9}�t�7��r
��mm�]�#>{�L��c@P���(��$ඟ���{q��xiJ�ʋQ�^jU��%�I���?����������s����?'�ȉ�U�?�mY�J������5�u!S��ً��O�˾ Fm�n+k��I\�A��c�R�6 ���#p!i}��&�rw��Y�4��>�[h9��W-2o�q#�-M��Ϭ 5".�^(��2o+�6�c�c ō���-'-�0�C�9�!	��0�;����ٕ�|0H��H3�&Oml"1ѥ���h�@ԧW/#�1�"��yB��G�OOI6l\j�����;5����QO���\F�����_�!�����Cs����Z�X�o�%'?�	�苜��w�!Xe�����]�B���y���꽽�M`ۊ����u�8��}V��KI?�{�z�F�y�S�l�I��RzFs�����G,E�%��?t6]�!'��&=�D ��1cW�C���z�=kЕ��³�����J�M�S�`��$\����Vm�?á�ل�����M�R�%n�h�>���Y��E%L������44�efO���v/�����о�u�m�4��z^�N'h%��8�a�4�����!���yA|<�*�Ene��*0��Y�|�� ȓ��%G�4��$�],��6��J{�5�fe�~_��Z':��/�\E���c����H�	r1��p�{8v�Y��?Q�^ws���F+�M��1�C~�7bЇ�ia	q�u>gxR0FghC��\�=�7I����2qw�n��	��;�T4s2G��:ٛ�|	��6\dS���1��))ĸK�J��~�9�I	<�b�V�F_ЈUA�N��E*_P�;?�b���_����DT`
��?FA�3�0���8K����s� ��S��+�R	��D<#��>��>��;c�罯}&17�O�����g(��U��u؉��яÛn�����`g��	#6;���M��,���|6��Ꮜ�0x��*�άsH�cN����W���������� �����	M�q�ŗ�gJC��~�l�r�����0�F>���`�]�$Vp���l�����ڹ�����_Ӑzئ�ռb�N�W	/�J��� ��d�2\�aح?|�/>�%¯���+?����Fv�G6}�2䛁9��Yõ5N��H�,�D�ﴳ��7��.��XX߫#D~���:���i�",�꡹'�4�'a��E}�u����uǭ�p�jZi��ķ�U �qsĈ2������ pì�T<�{�i���a�4_���Vv��^�A�g�h�ї)�=yGr�2�����wé(�ˍ�M���j�BԴ�~yrQ-p�dKć�����?���(e�icM�A��9�$�[ada.t�b�K���Ƿ�9HoSʉQ{�<��ة`��O�C��]G%smǵ��V�V6j���#b�:[KIŽp��o��̆��;'���P�P�63U�z�g��_�U&��zG��)�+��Ա�8��'w	������J�G�d���&�.�%(�'���^�3�?��;����礍�	~����������އ*�����z{�gm����H]!ڔ�U��5U����]��Ն�wQ��q}5�Nܵ�0K��:��mZ/���#I|��d���������Uc�y�G��rq���f�#?�x%� ���8fl�\�E�J�5?r���O�8��]�ޜ!��]諊�}�TqEېX+��T�}*��<_��Й���<_��O�JJjGyZ�C���J�s�^
dD_���e���&�p���R�'�@z�]�y6�ew݃���RTd�M0��,����M]yK��q_��p�f�y�"+�[QV�﹝Ƨ��ԉ�-�D�>���>�����]jg��o �RW�^%=��d[xĉ�(�����{�`��ps��hQ�GI7�	kڄ�>);�n�)Z9j�8;�p�a�;?�s��pfi_�0{���j5���F�*	"2fK�mX3��k�4͍9L�.t��'�K��V)�ӹ!�.C�5}E����f�˟���WX�i9�̫7�HBP"7RaQ�27*w(�%���>@��"���C�Y�.CS�걐�^�#�fE�{���4�@�v��i�y��wN�p/°��tP��4 }����Qm�W啡����ڄ��=�UŦ���O�ڋ�}ײ���9��S���n:e���F�˜��D�� k��)�O�?4^Z�n�|3�������E��Q�	�_���N��AE5�F�»�j���SU� 0hz:	d�'�7R��D֩�7��u�y���Zቹ��'���߭4��#v�T�C`�
�_�+�?=����3.7�On� W�N^�u�0��V��͞I-A$�@N��<3���a�s�0�w��(��p�vl(�2Y�a�E�*��/̳����,��[�]A˗�u��ܰm	���Yb��i�c�M�k�j�ӯ�Vg*'�'��!,a��9Y�L�{s��N�m
1Jd9����g�����q��';����Ǔo����e�E�a{��?a:�G^v�f%V?�C��a{�����M-����4%[�ڰ9�U1�;LS~gM&0`��Q��U�诐�gK�Ir�ܢ��X�GMNu��è)��� ��)�N����CoQ�S�ب���=����OB�3����K	�+������b�z��阆'�O�?�!G�7�0�����}�����>���-&����ݹ��1�(+!w�t�Ԡ��G���;Y�����5۲����Z��Q���v_8���S�#�?��������Z�U�b>�hEo<�`±�J�򘭭;���\�;V�eU�wx��Et5���ly���0�]�������5!j�
?�8p7�"=�0���d
��s�T϶�-*� ��UGc�������CoP��`C��9�h�=>��P�� L�Z7���5�����׳�CJ��gB%rXq��K�]M��n3���<��N���!��[A�y�}� �0{r�K����v]e�8{�xڳ��c/�Z(�u�$;X��fh6q� �iŔk�,�W^�(n I�	皀���ퟁ�L"�Ր�z�z���c�cU���PJ�r�����5M�_S���s#�'� 	T��M�k�;Iw�&A�7cg*�6;���
!dE��#pw^�Y�D��heWh
���-HD��yk"颯^*#�=��+xd c"MG�(���(K��`�3CBH�!$��M�;�����c�����7O�p޿O(�1�v0�Y]@�+�/^�a��� 3o�NA��
t�6��42:k$
;p��1%$�L�}���/���،#���`9�~�:�x���S3�ogI/'��R	�z&���Rf\9�eva��x��A��4~��g�4n�e�3�F�uBˬ�x<���y�=̜ѕ����K��Gv��,HAz�pa�וtGf���������t������aU�=7���í�W���fY��X��<ݎ�h0��#��M['�`��\U���G��Z�c�T�â����RRd�c��m��׵�+�*Y Li� ȯ��o�  ���iy/SJ ������t�mL݋s�	É�y%|�%8�	�4jM�Y�߁'�_y�����n�6�*�-KY���{�ݯ�CˑOc�$)�.�j� �������9e�D����Z��ՖJb�Ed��c��z�����a�,��˧�{�Y��LQ,msp��Ff��LeW1�)ϒ�Շ���i|���x-�+g��ũ�=���(S�2,�mn�	�L�;���sm����oZ�ws}�#S��h1�~
)���K�Ӥ4Y�Ԣ�	7P��x�_��cA��Z��d�P�?�'�̟��ӷ�S�
~�#F\���w��K느����c�`�+?�f	�C�$E#^ea�	c�e~���SR�{&7�P0�����
(ˊ\���us7��;�%�ר���I���k��4o#q,��Of�'9є7�����z�٫)���
���oc���ȹ���WW<���2p��x0 ��7�,�Md`rŒ��g�D��9����Lܥ�J�!u1��r�]�~bp�Z�l�i۪�����)�;���k\����&b�o��Rlo/>���C��d\`��؈���jf�%]�$��$�?4eْ���2�4}S[��\q�Ӕ��5�t�H��D��'�lE ������� ���~�::H��ig�}�7���p�Ԃ
4P�/�s�#��J��]Lvu�1z�:j�Q����U���s����2OB�@ k2�k�6��i��gas����cDV�ߥ��XA� ]��芗�Z"y1c�HҨ�f>�w���f?SM���i�B���~�yB-�vK��փ���[�������c>�A��99Z�[<IN.�y���r�1���o��Q��V�GY�`a��OTZ��wP�%�4��Er�VQ�0C�0#=��[�߅�|��j ����;�������;3�:0���rڗ�1x�iG@VD)�H�O78d�'��	����EcG��w��x1.�Wݢ�2���3<G=�|�_��20��-�Z���^~邔��А����;�t�u��g�rOz%xx���_��o����]�,�Ձ�wvX��,p���
����*a���m�W���|����R&�Tz�B.��T�^���r���a^�?/�����g��X�lw��聲�ׅ�5�'���|�O5�����c޷,ٍz��e��MEv��X&�PT1eß[�1{��
;o�HЎ�S�J��oyU�S��T�_)�y��D�c�������5)�مH'�I�zh�C���e�]2�����;�Y0ʢ�,-��myfl�q�R���Ydf��"ƥOQQg)��ߧW��������44�y՟�C0$]e���ʊ�R�֎y��=r
[Sr�c�����v�LTM�s� *Q���I��k�o�>Jo���{i)U�}Ǔ���\�a��D��z�p��S_�����mR5�w�ס�*Ę�ff�E�i�3�TkAI��(��)��܂SmK���)� !�\C�!V�\�ҟ�a��D�W!g98���&�7H�*7��l���%d鯀��~-W>[ 4��aQEC'�)��g޸�i���Ʉ#�	5���y��s�������t5�w��Z/}���Y<�f�� X�'#b�mRT���g���?C�X�v�!�5��s* }r���/W��G4��O�ى�u�i o�]�����I��iO@k�,��v�|�P��� ����Ew)Y���_V�H�	r1�\�V������u�
�eU#ǚhu��d?f���6�����a7k�P�K�QZ�/ꉴ,'�nD�h��>�T��K��p��f�'����C`7M_��Q�i�dui�ߓ1?b��-��@I��<���W��K�~�a	��K��v��2���a�*V��2���܅��%�,V���8܉�l��@��m<�LhPb�z2�~�xM�|k�ۗ����~�%[���ăNHFa���Yi�{N��Nzt
���9�;�4N9�tn�q����	7��co���ͱc�E�3��RQ�:��,v�:�%і C��{��e�u���Cq.[���9-��1y��SYY&k�C��]�P$��YKg��I����xuX��G��t�*�$©�a�[��N���{GJ��S2�6NK���Ī��3��I�b	��+l�u������O����m?��e!b<����[0a&�N�V}������x#�r��&�,��XӴ���+P�0�ۺ��E�&K��.��?���t�N�F���߹�_q�{B)*�>����ԑ����U4$��c�o�<��l�[�!	έ(6t�צ�v�Se��Hx�<t�|��e ������ }۩ǖ���Dj�ԙ3�M7@�����#��d��6�Ny��6-�Օ��G��a�nVi�^G�� <٣�g�ۣ�=�6�P��L������Pi;����9��R}�B�J�q��+�*ǝE��� <P��t+��^��}����rx����J]�|{����ٮK�5;(��v$�M�!U�q�	i@�x��^�ٔ	9'I�b���l�WeQ����EĐ\D�����r�U,��#h�J�u��I�5ȐJShU&�\+� ���$��k��"I���A��9cB"�6vs��Y�!_���ܐ�w�Yut�4�h��W�����-C���b""�F9^E>Y�f+S��c]V"�����#��Ի�>C�v�!?Oȣi;����ʲG���F����O㿍1h���q�@�Ϧ/��e�X�����Zs�Ÿ�6��!寑EFs�;�5�̖��GyҬZ�wy��So�,��Z�湽Ӣ�B�N�zo¸X'�*�	-i�|�c-��y|eX���z��J��c{߽����@0���u�}��sBu����<�Ѱ�!�o׌�"q��g��z|�/��fG��\���4�(\Jt,�j��R�ߜ��=�5ﵾIWO-��!���s������C���^;M�`���\��4˂Y��u5n��=o�}�Ж�R���^)r� A�ps��E��L�>�Ȋ>	����b��f�/��~�[�0��@m�8�N����!�%�8��r4g1ģg/�B��y7������n�ν*f�nY�-�֌g�Z���jX}$�n��Ef���7��k��e�����Z��q�eB�EߗKca?H�2���?�T'��&�T{���Y_aQ���sK�4F�N��E�1����({�L�i�U��k�xb�gޫ��Dӱ=��&߃�r2�*�n�b��;|��s���p&q�r�j����SP��1�
�)��K���o3��o�[	2[��mn_FhvA���;�5P���?c�%YN~�S��rH
9�+Fwe��&P�m�K&{ŭ�����	���e-+�%�	ِ-�#9e��D6� ����	�3�{7Hq4	F<��(�5�2�u�� ��y�[�T�
��VT��Ɋd#�=0�Ʇ�"����L��0�ň��&�����"�2��3{����WbM&RS*�Mi�� �=��g��M�npō��g fG��.	��0&��N���˄�9�X]3��p��lq��e�;���7��;c�F^D�0�b:TB�M�q/�8�c�uɚ�\����cy�ǥ��%�.g��g�?��^��Mq�}ΣN�7ɬ��I�5�/H�(>DXj��'�,��.N�N_N����~���:���i@���ÿ}|���u4��
�N�Z�볏���u��E&9zj�f���cZU�sz��m�0��� f��G�Z���i�da���tg�V�^��_�A�Z��b$����yL��Ñ-�A��w9���WM�s�Ē^BJ�~���-f�K�W6��;�=�*��R�=�c��`Aɼ	9��{[Nk.���Lz���X�m�o�5�Q��8��� `<U7O��cq%��k�U�B�Vl�����#�[��������e7;�<G�;�7���FM3�@h�aE����-�Ċ5G�<!)�¼ʔ�8?Q�'�!�+k��@*��b�U�z.1X��g��r�3w��l���ԤC�dW��������u�6�����ѷ�p�g#o5���������Jy��R�z]L�Y�|D�w����s�۵�k �Շ�5��m�����|R=c�h���7��&g�/�Ŷ�Or�>F�\�?�S��v%��Bl��j�\e����5u����SO�i-������W���Z�@e���f'E�X!=!Ti@�Z�%�L�b����PK�1x�J���yP���ώ��(����D���w��6e�����'WsYz#�\����em��&���V��Z0�W�,�s�T�y�C(qUk��cFfW��"a��QL�2�o|�d��!�i:�p��郇�%��އ4]`���%5uR�����_=�Zu[.d���C1�*c�q��"�sV�OQ�W�I-�.k�z}>���I�3)Pۍ����lhka�!R�iakpű�_:�R5�#���F�*/)f�BFu��3���k|�A�� ��$BM�ݩ�K`�f)f�!��Ck-����:~�\N��u�UW��H9S3�̡�7H��#7�e|�hʒ q&��@n9e>v/o�':<�CbtY�d���A���#r��P��)CN"���9�3�e�o��w��/8,Q�^��F� 3F�^�m�lk�]�º����s�Ŝ�\���xP��}����hq�S�����.٤Ў��>��8Ǆ�>��4�@��>O����<�|)�{�uB�����E������_�LͲ��K�w���<��i�E�LU��]hpN�d�?eӭ;�]é�Vi�+�����Z=ak����':s��#4!�Yd�Ty����*���#s��{s.7��v��lƄ"�u�{����C�-w�@D�<�����$�fCN��	Q�&��v�?2Na��B��*����n�,�9z����O����wJm�����bp6��']M�#�k�AU�I�78ǫ ��@�'�	�a� Y��]{)��N@�
g��9��׏T��/@(q��16��n[o��L��E�%�筂�:R��v�.�%L�Cj�{WJS� A6�j���7[C�9H~q1���S4k�&����R>K��F�,g�cI���ܘ��X�[�G�ާ��b-��d<�N��)��H%�Smǵ�1��;)��G3��(��	�]+G��T#�����8	���?[3!}����0<�K�t�}F����3֗�V�-:�&�t�����R9+�	����ؠ��ʜt��P�IA��+Ŀb�1։�E�����_�*����YI���}�P�Vo�U�F�^Ao����'q�<@���P�˲l��(e�B�xߜ�t�[�� �����йSf%ۄ�K�v�jZ"�.�R7�1�d��>��d V>�)9 �,g�-`��
^�Gˡ�)7��y?��{7[���K��| =tĉP�[�Lj�y�zq��kL���3���O���N�B[C�q��'rT��X<�+s<�ᱸ�5�
�p� }��wH}�r3/I��8f][Y{`0��et(��$����aXqI�i�����^���r�I��Y�Py��� K`�>�7��ݙ�Uzd��~�pJE�Y�ă5CN�SC�Rdg�]�� �U��
kFKNI�_�A��c:w6��3���!Z��7�w�>)Y���q�h���W�,��Bt�->VTϽ�X"_
G^`y3��+. �c���^;��s�z�C���!Z(@C�;`��O�M���u;�&�3O���1"y��O�:@e��/�>��Έ
ݧ�����6���*�!��;�?�g(��B>���)2i,�;C����t���������I3�oH�'p�%	/�S���н��\e������S��Ҫi�"�*����<�ruxPL�nh��\������/k��������|z����W�G���I��C��t��.���7*=m�����W�h+�܆m掅�2@���뙏uM�.�`�	�\a�=�������J��X�a�X�nR�A<�Y{�#�b�+0�`�NL_ �e���6à����/	�݂g��?mB<�)p�����%�Zl8޹�4�[��9��]�y�dR���n�*�JY�5��1�1�ߟ��m$'�� .������he� �p݀ZX�q��B�EZ��c<���mSv��l�"��Xv{iq&Y2J~Q"�s&�8F�')�FE1���H����i�+��檺x�*g����>�=}to�ޯ�2���nl�z��;WP�s�o����m���G�@S�<1�_)��K��(�-�
�	-О�g�_�A糧Զ9sP���??���yp�U��
�XF��O���1z��Ka�.�D�y������+��[	��`�#���0]��c����+��17��$����k(� �m�u��K�|���|�M 7'M���@� �#�nd���k���7�g>A���١���,{�]ȵ�4�e���	W�c�5�h�w�n�< \	��=�M���ň��g[�㺯�-��4إ	����B��t�
]Α�p��*l̇|� ���yͱ1��!��C�7b�X �H|/����)ɵ��\V��>Fg��5%��a����?��B�q�h6�}I��A�
�c5
UH�V�D�W-��V������h���~1<:~ �i9_3п8&�
��4F��)O!�&=0����u��-�|Zj���XU�5[sU�K��W�x�| a��?
��<7i�}�ai��O��V'�d/��Aش]�y���Zėyg�	>q���wtH@՜�Mܯm�W�BD~��-��>K�ѥ�N_����_�ܘ3��םc~�=A��9%�[�r�.%ڛ��A�����(�o���Q̷��=�`%�O��f����%�W�����3YV��v9�4#�V[�kc�A�J�`�r̗��;X����V�bj3�f0+C¨�Q�Ip�&G�C�)9fd�E6�8"�'(n���$�;��u���|�.L!�ݘSX�Mr�3����wѨ�vդ�w{:t���G�x�vP���8�A�qs�k��g~���T���ǔU}�%K����e]�u��w��w,�ʢ�H�V� 9Ӱ>p�8m+.р���|��B�#�}�:��8?��
�|�N�rB�f�W�$?��M�1gF�*��lm'�78��G�5�[���O�1$�<x��e�p	���i�5��E�RnX�T�������g�g� ���yv�l�JmiyK|T��{ᱯ}D����R�d�q��A'���z�[Z����e�\!���ֻ��5}0�,�,��֛�y�:@q�灓��8f�I"���QG����s����<t����u���`�y��][H����9R��N��,%=h˯[	�2�پ���E{l�
�s"�Q��I�d�kk��>�[�����)Kܙ�I_'�{a��g��g5p���_u�ｺ�i5����W��*:�f��n��-3�6uk�aV�^D�����8 ,K0�)��!��CFYx��X��aW�g��f�W��9n�[���H�t7����߯6M���>�~2�Yg5�C�1������94�o��#-��k@��o�L)A[�3o���x��j�1w_��/���l�\� ��SmT�Z����ڵ���p��o�w����}�Cj������w�F7?ٿ˯�_������y�Ă��O��5/O���e*��"�|���P��6��E� ��oJ_��*�Xr��s��D�z�UYtxhk\d�8��h`@�֩W�����Ƕ�Zزd���'��l���9�t�T��Л��ܠ3h1�vØ7�*�Q�[Ɵ��u_Q���(��~��-;@?�`<D�l���㉁��W*أ!WvJ2�a���;]�`^V�1֛,L���qW���*�vum�}��b+P��zIM�]k�Ǣ��6�/r3���*���fa�Y�Y_��{�N{�z
e�9
���z���1wq������I�vo@m;���2E�7����:^uv�B%ǥCE
D{���ݛ�n��F!��IA[��O9c}�1o�uS��&�Gh�"ghFTZ���.g|�9I�q���X�8�G�V�`��:�7�"�N�����L �iS�յl���y��`�*3@/k��Z	�x�+"5�NⱺKO��At�`�?D�!�r����)0�Z��}�q#��̗.�����p&#9��NfS���I+ƭ��E/��c����e��d�E�h8=)���Yy�|����m�_'�n����t�s��l��/���)Uj~�YNyoM���w��W�Э��ˍ�c�Ee&��xڜ�tF[�����������y�_1�BF(j�1(�)q7�A�aڭ�Y��d{&�N�gB�-�:H��Gt B��7[֔W���Rɣ`]}�cc=rIP޼LL�{ۻ5�/��O�������J��?pB�[oq��?����S��FaD<����O�E���~}����S�r�и���]�U�{;���O�� �(�[x$L�z����q#;i6׋�2^V�J?̝I�\<童Q�ʹ��;�P�JE���+˂�4�eUu�[���LJ ���&^�5�+$SO3�������B �q��t�k�I��
Avסc�qV6���(!Uu��˨w���Y85	�*�h���Wk���y�-9��"��^{���l�+	��c�Ȕ�����wn�q}4Cs4�!unY���;;n�j���������	OY�	1=�����?@@w6/hꍎ�!�_�[�;��6�z奰��p@;!ꈝ��=#����xF�)B������w�/�B�I���D��ox�'+@�	J��r#���ZqeGG&�؉)�p��e�7=� �����/�w��uC��i�����j�n~������eNv��ƹ�ݪ�z�)���hGw-u�6U�^�ut"��������Y=����-W�c��M��#ҕ���������;dM,be`���\f������'[��v��3��j�R#�ہT�<~Cd��'�{U�L���@�ڷ }��V���j/d<��t��2�m�~��l�:�&%M�s8���4 ��,;�xi*y-򱛖�inQ_{*�l�Y�����;��\𑠢u$�����֏6�}�P�e��g�:�Z�Ֆ�b�EվqcE3��A��u"z���{$�YMU�Q�XHs�F!Eg�1�S�ϣo��½�i�! �ad�x��gT���zʠ=xs��9��2]^cn M���t;2�sĔզ��hqZ���S��|1*��)B�Kt0S�G�ڥgN	(e �µ�_�ǧAk�1�<P�}�?z7��[�stw(���
�P�F����ȿUwBK��˭�ڼ��?-�qZ�+p�<	�\�F(#�Ī��kز6����b�;G7�i?�	�|(\��_uD 	�wbc�/]I�JB���L�����#"�,� p>�}�HC"����6��0�qm�Θ$��ڈ��=�W�:�6��H��45 7���ݤM5�tŃ�Lg�`�j(6��X�}"ò����i�]iKXp|�6l'�ۡ����뱬 �����~
�bp}��C4K/Oh;�������\�UI�3k���%..��M�?E�ג�=�΃�}Ĕ��إ�EP�5�H�4De������}�D�m��Z�~l�:��iR��>\��i�%Te4���=x�a�d�.^�u�}1���jF��0�U�Vs0,���t4o \�*��y�g��i�5a�F�*ϳVb�ʌQA�.h�Դ���(y�w��p{����w���7�M����z;�B��8~�NF-\4�K{k%��4�sq-�ר����c9�>A�@�9��$[ͷ5.`���)��bڷ#c�o?!�Q��T业�`��O��H��%K��!W�BD6V�����#�.@[7b���T�[����G\;O�ݝ<ٓ3x��fDs�C����z�pGqj�)Td.����8��'czm�ar��6������-Z.g
��`]�(�3�,/�Mv���H2���r����0{H��:�+ES�s����f/\g��k��]|��� =x���d]�J��r�.w�.��]B47z�{&�Ӌ���,�m�m��{/�|Bb�ދ��U�
��w������_�r�s_�R�2?@������Ey�l誃�+��6��5����w�OF���k��8��������p�-EG�fXET���w|����{'s���Q�� _J�X:yFxj�,C�6��N�D1��-u|��#��D~�:�'&"z��;��&�ec��iD��>+��>H0�!%,>|����y�Q�qK�$�s�:f��j"�˻QBG�%�질�Wv�0JS�P���*&��}]V�j���>RC.��=�[�[��Z��`H�g]9e-\s���Q��,I#@kF�>���d�)F��ǤQk��a쇅�_�p{}t_�5�U��5��ײ�[*���f�~�k^�3gשk����|���ܓ�+K֑�)9x!٬C!��1R��p�,R2��+(YWD��9�C̗�{H�k�7>�w��������+�4�>��}��� �ֿC�������Q��ʯ�#���4��D���nW+�ih��e~w���/�'�.ɰ���� �u���m�"偙��xu��p-���IŒ�n���đ}C	D��:��	�����������0��B�ƴ�*�jw��y<OQUU Y:��(�|M��+��q�EH����~�_g	�:?��Il�2�ڻ:��זU�z�hf�/dPR#�#�r�7�P������[b��Zs$։��'�� ߙ�V��ҦTo-V�v���W�Dܕq3�7^M���ƺfuu�F���y˹��-��#@:�h<�+|�M�扜]E��j+��pvX�52�c�a�ܰ��"V��T�L^h,�0I��lf�����m�N�]�4b�����=M���kmm���t�n�P�<��̓|ma	��Y��{�4N�^�
�X9u��E�W��C�qdL'נּ$�bo{�͂E�i��cE�:���v�v�%B]�C �o{�.��6���C��T�J[���9~��1ꅛS��&�⽛*Ac��OPg7��I�{�܎ �X�5�G9瘟����r):�`TN�����06S�6������Ļ�m3�����	\i+���������=�jۇ�f�?їY!�=����0����}|Ry���ݗ����&>�������
+r���]���">�*��E��c��!-�}��(��l����/_���s���AU�v|�e.��$U).�T�-o��[���r����D�hDk'+e�;Mxռ�t�z�����v�I�z�:fF�}6�jP)�$\�7Q�%�p�t�d�����Ϣ=T-��e� �SGϕB��Xj֯���q�#�;�Ti:=�?P�=�L ���E��r��y M�e�j�Q�B���q�/t(˃�Ή7�ao�<~dŸbi��q/H}����INr����
v]Qr{h4������(�=�$��R�
q>��i�r(��t�^���EI�	��򅟈�~�V���א���f�����Up4��4nIJ�=L�A�59)S�����{�p �TH�5Jk�rI�<A�c�Ʌ6'�*Ռ!P���&wJ4YS�/�x�h���WT���x�a-4���s�F"���^�O�)K3+�[&c2,Ŕ,���̠C.��!�Ԛ9�/;s��ޤʃ�7��3��W�O��1X��Eo�@{�/J�j�)|Q [���f���F�6�H�� p���;\tƝ���8(��kR���d�Di���*a�j����?�Uo�ƕ'���	e"��x7��H��e����$	k�� ��X�m� 0���U�3Lu�UL�d���%�)O�����9��!�a�zM�j�Ù�G�}����+�yut�-��h8�M�=��Z����W`?<�R4���ᶕ(#x��3�Mǵa`�wm\��˳Nj���=�@C2�W���ATR��ӁO,�Fס	C���LU%���[_l����^/�{����߾9��m8ᑋ߳W�u��%�c8��T4xG�E?����hy����q@�n�W(*7l*Y��\��#���������$�1��h�q�P�<��e|&��Z�ŝ���MEP�c��P��O���m7�9{߸OYh��Q�s�u�FR:����1����B,�}��i�7H��=$x��g����v�=s��ߔ��2(�n;N�pS;�@sY��A
��c[\����S�S�1EoU)��=KO�m ���@�{	#ާ
+_w��ABԬ��Pd��?�|1����o�|���
j�F�K�����0,�K���z2��������++�a	*8 �a#�$��Ƨ��ȗ���uD�7y��Z�E����(7���Żu�-��rC���] ���]3��ǧF�ZL�#]1���)�)��n��KN�s�ٗ/
�L���Ӡ؊j�㹂�DWs�d�X=�b�d�y ��,lM�Z{�~!g���%�"���t��D�Í����K]%Epwξl���ۖ�l����'��#ߦ���b¤�>"/�?�甎���;\L�q��?��VGl%��~���?������Ξ  }?=�Ȑ�Ӏ'5U�H�zDi���X�
����_�j��~�sA:�gi�-�h��͵�@/�4< ��J_���-��Nmu��Q7c�j�<�KV�U�(~s�̫���� W��X|��"�i�	a_|�3yV��teS�A����/�1�Э�y��4�D�ҹ�w��i��E3M�Y���?B{CX~ �W-מ7KV%���)��������N�c��cA�j9p�[��.���1��]��~��o��|QR��3�N`�$O@�"��Z%���|���twV�7]/8�#��[rx�w2��V���M�};�
"/��o�3Sq�eh��<l�}�؏ռ~G,��)o� �;�8�#�'�����%`�1?��+� ���.��ݎ����	3(d}�蔣��:�T�I�f�Ko��n���ޮ5Ԛ�R�a�xg4$ f_�<��K��Ni�3x]?�m|Jw��{_OF��3��f^�愁ma�+�v�z|c��뙉��ph �.�g���۶�� rx>0�M?��I��X��`�lcN���=3�q�5F>
��`�O�"�����#��f�J��>-�rE�swX�:Tz>�Ë������`w��+ݎ�WJQdCyA��
����E���KD�����d���w�����L'h�VzT�� s-e����Df�y�`k �0�6,,�0���L�y҈q��S�NAMft�"2Q='���Cd��r���Ƙ+ȓ�e���N�]Q~��6�R��׎�&�=^�[�C4�O���jSbӕ�bGs��Q�I�;Qk![�>6���b)A>������K(ak�����pV��_�w����5��M���*���f�L8��&3B��k-��͔��g��l�K�>)T1�!~�
C��l9��PM�F��	�W��F9������H���7y�c�9iXƯ�j�@>�|Q�uf͘�Ca�5:��щX�%�`#��b�G�ed��]�_�x5�`��wY�/i�(I.��R 8 �-/��m�|��|g+���+f'�N�0Z�_�)�}����Ө�di�������!
�U���ɰ���$�T��|�eO�8�ۧL��N[|�6��-����E�W����_�ܲ�4��Z����^�������U���ha�_d��R��	��R�3�Mu�˼���=+cZ������'K@��T�w����T��q�Q��R+�DA�l�A7����|D��8�uU\������?Y-H��@5<-<��˫�-��m�M�J���v� �26�a�2�����_��g,Bܒ���� �{���um�?j��+b�)~��:M�okH3����	aG�Q�:#a$6�YUT�{��N��Q
8l�9 �8נ'�`uaq,�	�{��o�{���?E|�m�֞:��Nv�%�4�C�w�{�4�ѝH��`1쯢T[t�9��1e�MS�`|&W���X��<�W7�g�{I����	nfXbR+Gt�z��AYλ��;�m�kN,���|���RSi쵢8���U/�53���B	}_�+��v��^+��Z���>�Ϟ?��!�(��yK(0��(:�)}S������^��&Y�$�Dy��xM{+<V�{Ƀ��Ҝ�_	 Y�$����I�:]��B��ˡ�_݆�.�m��힌�Q@M~��,U�jV�O^oΚ�X������`M�C�b0e\�~x��0t��G�Q$�'�-��V'�ۋ��F�j�@\�g�7����%�я�Wdq'�8���X-1 [���G*+��Z����燅��i��0ۏ��=E-�P�ޫL{���tߙ��W��ƈ�@Q�>�ZB,�q{�����ǉ�R�|�(<�U�=83��H��}��mY`�rdt�$j]̮�{�3���460/(�?�$_)�H:qY�i,��s�^�b�u��I��u�a^��C�@�q����������e��j�_Uk̒��fJv���\�j5�F�S�� �=T�.�U ������IkwjI�N6Al�:c�A6b���ů�!K��H�w��Ynu>� ,�h[�W�G޵�0-/��β�"��^���I�+�)cI�W�/���߷�'�C�q�!�Z�	�;�� s�������`�7�O��1sl���/@��/�����:���� ���:6�r�O���;���8�u�3M����c���_��� <�����J3�:��o.�?'��p	�5�h��ޕ��6e}������d�^��:s�����۬�&��6uI���_�v�m	A��?G���[E뎜��S7�z�D���&G-��z��h�t���C*+߈{u=>������W�ڴ�;%�߿Õ�� ����J�]Mb)�`�^0\T3�n����h��/������	9�RY}#�J1x4�\&C���!L�\*��m��a�@+����/���G�"�TPnm�c���Sð��%�K8�1�4ӎ� rׁ�]Oy#mu�L��n�o	*ҋ.Y���B��F�]��l�$�1��EJ��x��EezZ��U�Z�ʖ�E�eHc��ޛ~������Q�{��*Y��Q���s��F�s9S_1z%�Y6R�8[�in��W7�xtE�g��ŰAp=nѲ�惘2�1nVoJ�b};�k�s�B[��@=�^e��X4�S<ȩ1`{l)A6K*x[�N�ۊ!	�7�x~�_2��A89��'itP?��?�����j�m�f0�
%F�F�-U���hK|���k�����'�k+��	E��g#����0B˲l�*��!e��744.ufn��=(!L�uz{k�mD��}7�~C�x�{�B���5"�#��y�V�+��x�����K�15���'Oy�=x�w�}K<W�fO>�v�Ä�M
 �,K�SӕMk���ypQgl+�����_�z,$�hg3�%��]��pr��l݌�Q10�&���E�Ӳ�ݦ�dgb�&K�9�/7��Oq��Gh\�0F��lǑV%d�����?����J��ιE�}����h�ӻ�5�Y[Hޠ�D����Ǒ#�M�:�=�E@u~�Q�:O�3i��D��iQѡ[*u4�~ﰺx֟ט��d_gu�����j���f<EU��s潕�YԇI� R}R�J��ݩ�i(�&a�3��V؛� :Aɂ�ߊ�K����y��J��y���w%��m�M��D�0dZB6�{~}�-R)K1�T��>/�ʐ��(��e[c�#�A5E�9�E~[���.�ک�X��xL��7eo��FQϑ䮻�`�T�O{�~�~��%����ׁW��V؟���%#��c[���0f�Q;̨�;���JcD2&3.��ܦ��y��x]��0�,G��)��:���g8�TZ'�򉅗�Q�,�˟����A�I.�<�	�K�ޥP3c�������L ��k��f����I�20���B�u�\�g���!��;~�����j�>��]�S�h$w=]����j빵qa��A;�!�sm�Lm�q��|��a�T�ɋ=���H �	���E�r)١HT�?����b�{��l�M��p�׬��5�U��iBO�J	�m��>D���Ԃ��g���E}4�X�{TՑ��F�c��)h�q���^��IJ쏄y<��e	�Ϭ�3� 1D�Y����"b�RO���s'�Xkzz���eY�2����"0�k�,���@��y�߸qA7�)�ofC9>"̈́�Q8'r�۹@��N����U&5�������J&�]LI���	R��� T8=��'[�#���������]i���sB��Q*�0IW�k��N>q� ���)<���Z2X��a"n��U;�p1�Z_&�����A5���h4M*k��f�:�a��3y#kh���/o��^h�ICkKL��)o
Y!���Cל��@-Ҧx�H�@��
�W���9��J̍pHd�g7��C��pK��G2�%�>�+���7�z�CN)������T��>�#^������q��'������[�/wpۭ/$��d����(� �e9J"Km%9�wU��.����߾�ň�1�:��<!"}y�ߐ�����A�w���}C��x��>�*�����wa�O<�����|@���e���*8E~3ǽ���_Fa��_��8�(/����1v1U*��h\��d�aә���m���˗Yw�x�7Z�g!��e3'��)�������Te��,RM�����]��gs�7������*�uБӓxw��/��-�q�@0��<U�[��Ӹ���\��K6��pyv΋|2�(a�H��L��~��ι,��Ȩ�ԗ;R�G.m�P?�b\e۞4?M��
k#�5���)Vg��k���fa?��Yе�{��N,��
ӟ59������,���qGV(π�N�o�2�͸<�Ew-L��K:>��v"?�%8,C�^�{C���l������
^[/i9�:
1��S��&�O���dw7I��>�g�n�I��܄��X=��G�~�1!���(nd(<�NG���uG��SYL��=�9���>�q�3q�1Ò	��%+��O��L���z��qW�?G��!�3����0��u��}�sm��CV�?d���y&t��տ2��S6�+wZ]�U��� ���=����0�k΄G�u'�M9���k�_8�����ŹP�l�<���B*U;���J�
o^��W���\ѭ�������UDe��Hx�\4tW��M�B��?<���o��vj�x����7����Ѫ�d�WV��x��-��(��u{G��c�����_K�ge������D=�:YPϟULּ �f`���3�o�г�[�yӭB�e_qv'1����DW����<tg��y����Ae��}�58���rv��*]�]GW{�³ s@�~�(�a�$]�P���Mqt�i���N�}^��TI�����������S¡��%�������Uf��꼢J1cφw�5/��S��/�>�`��� �:+�뻉k2B�I4�A�9c���6�E�`��!F�����Bw�a�Y�E5���h6
W��1��J�-*�;�)�4"KY�^̥�h�+��c�d�ʠ}�
�ԂG�C�@�!� �/s�;̄;'�ʹ1���q嗒TO�@1����;�@��&/�E�_�z�.
�p���l��6)!��O����;���ӮT�.���!��h��z��~`�G�������5�Io��	'\�|	�����vt#>���e�d�ɺ2��Җ�P��_��Cۇ�G(�uu�ڬ�Z@��n��P/�7���p?�i7���-cz����[�G�~��5�d�{st����p���|a=����5�W�ͪ�aU����������/� iM��`�e/\w:�)�_���ۡ6<���nǖDP�R�{ˁE ���c'��q�LK���`�у���I��7�/u�Y�li�o�m.5��w_��È%�8ʙM4.�����ہ��y�Zٛ'Z~n�*m��Y�A)��(ۯ�z��G$I����|��G��r��euX��#ZDwZ�삠EF�c��ܛY̮�Fu�9�{U��Y�6CQd�s���F���B1u�xϴI���[i�P��P>xO��ga��K-,=i0��J��2�>nq��f��;�_�sϱ��w��Y�t䳝�S�\�1{��)��K�r�V��vL?	���T_��ASP�Ԣc�P�%?+gʝ,��eW����
��qF�/���8r��BKMܭ�A��������+��w	`���8#�D��k�B�����w0��7��&�>�z<(�k�Y�hu��heh�@���9����ͽ�|��#�s���F�	��Y%�S���L��ٍ�@����I�ˊ�EB�xpW)����s��&m�Z
� �x��M���t��g�������/����3��C^7�`�]]:8�pmHCl8y�����Avv��ӍG�/BJbA���4�/`N��
t�!�=\B��ت�����s%��|���J?V����Ԋ�}5�L�~`t���:5��H�N�DM�����>ߑ�� � �~P:�v�i�\����$�p�vE	42����ݟ�{���yu�����jw���B�U}�Qs�����䦖 M�@9I��cUiC��aU$6��ZtV���@cA�\���E�F4yӫ0*/��7xw`1d�	tMȃ/�B�£~6D-��`K��:t��D�&�Ș����cj~AP��9�:�[^F�.l�S������4�oprTQ8l\�)��`���O�=/���%����2GHs6&V�'�%/N#_��[����M
�L)��A;D�]e֣��X3	>��.��s�����zG��)�}�1��8���'_&�2�{�'�3��=+��h.��_݄E5���g3�2��2֨�~q�
}�&'�񁷻�dm�ن�$7�݁�W�&g�<��3�[˔A���{�y-�]S���c�Uw�$�ʎ���յ�y�89\��m��f�l�|�A��]ɦ2��$�d�v�z�:�r�3Z�C��?Q���ʴٖ��lY����	��@'5|	�����OW� �(��Y��\ǫ�1�!ŎE�X��T0���͡����3�9]�XeJ���y7U�����g����:Dyj����]1,�<��w�'"`z�n9�6k^e����ൻ�Y��C�0���,O�}��+"yW�q��V�u�f~�"h�Q3G��6���Y���<5�ڱ��Q�ۖS��P]G4���h�Rt�p��y=T͒[u#v���t�1�X�v->s���QE0�I���kא>��b�Pm�)7 �ǵҐ��a=�����p�_a	O�&�5�_0����*&KfI��r�3�yhk����n�uܤ9�Kw�)�p!tΪC�H~�g�A��Cx��<,�Wu9�gj�l�H?7� �o�����~��[�>����kc��|�C�fu�k㛸�Y�۵�#zk�hd�[�+�4!���:���V�Qw�}/ߐbX.�Hq� z���u�m�ш�rc݇�}ڡ7H�NF�7���%w}���e��:��2���+���KW^���e�Ղ;U}�rOb_7Q�]�+��|�i������"�aE/��k?_x���k,N���
���K���E�l�<U�NUhW0�da^Q�T3b��I2�CԵ�rꞳ ZD9���jG'i���������T��M����5=z�m�bC[7o[=�=ҽ�=ouK�;�S|B�j`�-~�@+R�<��+�~�����C��m %v	7�2U;\a®���2h�Lᨙ��>,8��Z4�vќ���m�nj�b��� LM��k�z�pX�?}c��w���YaZ�YK7
{p��Ngc�
n�9�i��VT7��8\qb�\��р��o,
��S��Er���tY�:���v=��%�C�C�e�{~u:�����1�e{h[��\9Ϲ�1[MVS{��&�<���24&�fvgh�}I/Z����gX�SG�w��� �-���Y��fNb99�rnEl�|S�OT���W�ֱ*��x3,_L�	s�e+�@��:[u����u������?S�!_��oHW0�y7��}M�������7���3�&��b�:��.?m+�~O�� �����;<iv�u����:�8ְV���O���U_����E���j��j����}RU�M�Eb3o�V��6��37�
����ؚ}e���x���t��F�Ƿ��]\_��A���$��.�`j!�p��o7b+��M������dg�Z�pئ�S�f-g�Υ��Gൄ��z�� ���� ���Ȥ�<x={h�Pʀ�L1�b�!l�����s$���,��D�Bb�4qqӹ9�}���u��Y�<�-���ק1!� �E}��>�rڗ �E�*]f{�+��;� l�(֣�$�AX���Eq�]i"i��)9�^Bg(�r,I�П��#���Ё��d�ؐ~��� ݠ.�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�$ڜ4qz^��.��?n��!�|,rn:Ѻ���p�Y������:H��{>����,5J,�1��=��u�����k�_Ř��7�7���iF3��p�ӱ�]X�k%6��`� ��}���>j�x�r#����-:-ڥ�|i����r,>N*�~LAׇ���P:e�}��*L_�F�w��Ǔص�i�L�����M}�o��a���"����)9�D&2Q�q-EJC�D��Q撋G�_�:�gq�55$qㆣ�u|��:X#G1�TF�ZZO�{�pV���g'm�p8����\*��}X~gO���T�-ӡ�	���V)�X����\d�h�dt�)���3"���>aF")���nE`�N�)z���_��"	��{�`���m����k�� � P�<�SH�U y<�qA���E�djq5�����jtjG��5�� �J��f�:�����q�SW�tT$8ȳ)�ˉX��/7��`�n����S�L�إ<O����d��-�` n��4`����}�d�νQ.t�3 r����-Zl��T �\��b�h��X��~}���Xfdj̅}k�ܕ��'53�"�#��YT ͘E���3���� �H�xX��-��VWn?O��*�"��&����"��2���� ����<knkS�S�������x̀�ǁpi���)��@dE�H�̯���Ѽ�Yk_ȭMx�i`zZ�����"�)n��G��Z=gD�kf7Q`o_�@�/�\"G$!�.
>4[v��'�|]��ko�>t�{��� �ZI�߷
�:�|�o!��IJ�D��~J�j�p7�M�I�yގ���0.�kj#�$Aq
�~��\}��OO���0O����q#++Ϩ��uC�4c��Y�a>|ԧ0��Uƛ���:{!�lX��0<k������I�G�ϛF�{�}�0�
X.�h���f�[��^�;}���~׵z�s�)K:hb���r׋4��}񉾖v�U��>��[������(���a�hp����J��t�>��#MH�PMxo]VߘFH�9������1�gݮ�(��e?Pަ�������D*Fc��q�*���T�~��er�*�߳7c��60�+?r�u��v3�M��WH~Vp�|O1LLe1m�kf?�Y_D��B�nrgЦ���O�!��Lv���B�r��y����ۦt#)S�c/^�x�P��jԖ��y�账�b}��"��,�wF% �;��P4�}O�x?�E�J=9p\͔���� LƝ%��N����g#�Z��X;��wͯT���G���cҞT���#< ({Z�C?�'  l{K�O���k������x�֬�%����8����B�#U�}%Y7C�F~Ў%����p�o��X8i�k��S@�bҰ03[mo\�jeY8>�}�� ��w?~�h�d�	R�[�9��R��`ul�O�5ZtWv�\NhdE�{B��H��YΕ���u�O��5]����B���z�E���#�a'��{���s�fH�^+=A���z��'�aG����F����B�����>,�o8z��7vx���iF齊�.~?ʻ�U�:��X���Jĺ��v,�J[�m���Kl���k��b�qIjÐ��H�H��������t��ec��:G ���!b�$����*x��`^��z�2b�-oY+n�w֑.��)	*��Y��b�<���Cu0��C�- �w���|m�a�x�Z�p.Q4����1�܄�)p}��Q��Y`��ӑ�?2)�Q�Ƥ� �5#oܺ��>�+)<�,1:�o[��n&��8gC�8�֯���+��>�
n}�U�<��j5>�F�aM8�%]$h���r)��:��js����^��0����a��ז�`�Ί������SCf[D�i��l���g1\�pH������z�O��3�z����~���]X%�F���j'��؋d��c�
����u���F#� +�j6X���wA|��_�A�h�ci�����Wt���ӸmJq��z�ߠ�]
� xN2��㑡���$]��
m�u2��(?�>F�GI���T����*_�uq���&TI��uV$\G>&L
K����x��!_���%��T�� �hE��!��	���h��!�zfU)��]zar�����m���F�7��.�mD�ߋ�NC�����5�t��wGMc��3a�ϭ$���i�F-�[���
��9�b��C18�rSf��)�?����*u^0cw5b���1�t�@<�-:��Vݒ� ��h� �zsQ�@9TZ��{J��2K�a��N��-������w+�f��2q�'�[}�Rڎ�"c��Sd4���5��({߹GF�kpJ2�{؄c�^K�Ś���it*=œ~Oi�pX
�i�*�%Ga^���e��՘=P��[Ӵe_�7|�	��C�-��/갰܋�{mZ�$X΢E?�A5�g:�i��;��6'�I8�j�s$���!�g��%!��~��߳�HT6j:~��BD�ˮ��j�{~�c�����S��p�����`yߐ���#�P��z���s�2�*�b�a��ط�_��Mj�ٶ�d�29�B�F��>NjUow^��v�`h=�J ��2�N���7D����O�>����[�����=9V�I���D�Yg�5r��/�1&�
H"�����,PG���YN[���+�����3(ku4-+�PF��pm=��A�SO@��᳌3I���r@��%u
D<�� ܂N��@�L�er:��81�fĚ|h'{��[��ҿ�8��7��n5�h.@��������fx0K�Y��&�6�����ge9]~�xj^����o��x҃��~��Ix�e�U�N(8������S@?)C�{wnT;����'�N4��3���`CI\F[� /�I�k�b! qF��v̬t)�uE~̶֣d�ƕ$͞��:�Ek���I0�Z�V�u���:���G=�wFLs�OI���q�x�g��||��dlg\6+}�b�O�6�T:e���2!�Zc�)��?��F\pjPV����~72��MO�\A)�q�n���Z�Ez pk�F��$��e뛁sP�
%� <�X����i\ψ��U,�� ���IN9�v$H5;E��=���jS;�K�k�%�����ȯ����Aŷ!�C8;C�j�!��+�p|�M��wĵ�D�P㷆�n�`�C	�D�H����_Q�R4ڡ�חi��V�X5���o0�5�S��x����9c��>�\��k4�Ul�UK���0N$:Oz��x��Z�T�kf8�=��B�|5r�E �ֆ �x��J�G�
�7i��9�� P��zXE3F�
�i���G����N��c-�6X7����d��9��,��M-�s�$�N�q7T�����<�����,���ї�ھ���9=���������	�>F�6�i��J	P\�mw��
�S�~z�kR'ߘ�7���Gব��e���.�X�%�L�使F�����M��$���3-r�ҙ��I:�_^X����r��zSj�~)�ᇔ���:"���l��L\qY�Kq�����y>Ʉ5��z��
t��ia��~"�$f��2V9��&��x���u�uO
:a�æ�(�w3��1�%�;��<��!���br ���\�H�X�iKc;�/��ʄ��~D�L������V ��H$��m�2U���9�fm�]d���L�b��c�:����A2���Pp�n�}�Y5���1gUS�!x�ӁR6���9�s�hAN�M�|)��G|�#����ءpS���]mX��V��}��zCɞG�{���8�X�i�0�ˤ'�LV5�;㈾h��U����E��Q������(�#��yɌ�͛}0��"�f���m��Bm����
AB��D�}�F"Bn�cO��NB�RW�̄ؔ�&
I�*omrtw�Ȼ��[d袅bGW̪<\Zaʩ�����1u����ddգ!	�{N����&7ܾ<B9��i1�4�v=(HV�������q�㫾��S��
�У�n�Ե=�F��O 3�U��]�{��̑���&�1�sߍ=�*B�\�M	Xyr��pS͐���ժ�ڊ�Y^�������C@��r�8���,��##I�����h����İ[5%��P-���LZH��lq	�^�
=e��&H�·/9+��o��k���Qis��itN�&��z4��8��W�;���H!�ksA��������?H�Mkv�������.��d\&�qN��Wv��5�dM�#ӹ��UAn'����>��/��?.5��Q����4�$]U
'�Vy,w��y�Z�-�� r;��4t�����|���ӎ�[$�1�/��F�ӶvSR�!8��ܚ�k�2s�����(��{Uۉ�aN�eF`$� -�����9�0�K�)���#��z_/�ٴ��B�#��ϵ���z-�L�8쪆�G~��c0<�BK9E����T��B�7N�q;t����N���~��z� ��Mi���*-����Ab�.��20e��\�WpOi���$�9;O4�C4C��D�����{[�DU�<$�'#��Pê��`2C'٩�[ݕ��NT 1�f{�^EUP�])u�pM���A��m�. ��-�V	���,�Os���lux�8���1��c����[���qwe%t�����S��I/��~�ъH�Ƕc��6>��g+mu�l�^
+l�8���i�b�ѫ��,�" ��?���i�^&cC�Ļp��������zu�Y��B�X/�0qw|��Ѽ��x��j�^�θP}��j��J"8��mBQ��f֗�^�J2�yW�OxV(�_n*�����EwG�$bPK�1+l�xg���^_��hdj_u�s��ΩK9�	��ѣ�l*��{���8�ݾ(��f�'q�`9��~���%��,����$�����g����&��g�C �U���fi����?��e���$���� �B.!ǟ `"�Eg�@��^ ��z�?�[W���[�G���6��!ݾ0���W�H��&z=?(��(�G(�+�ZԿ�p��4��T?g���Gf��X��E����bLx�����y/t�fz uE-�.�E��di�����s�x{��g`{"�C|Tȼ.�I���@���_����9��)M�Q{� ~n͙d��9�#U�ys�S���w���m���y�o⸋C÷_�U�͔��&'6��&a�p/�6W��kF�\?G8<#���P����<L8��ۏ}��	���ߓrP��*3.{ľ�|6�*.��K@f�_�;}�[��)��]{��@ `\Rͻd���[UH4��5؈��55�G�y�=��7����Uk
�ٴ'Xv�&�_/c�����:
&G����>������<1;-];��/�<�4�1��K�t�!�|	����)�<Kðᵉ���渭�K��X����'	,{MN�=��cZ71<�]~���������{	�sX��N;��b˯�����.�h�57�B��	�=����8��s|O��W3�&"J>�n+�H�HF��clG�/����ԗ�0F*�J��ԯRa\�H���ޤ�X���������/$��~� (´�qBs�2s8T��IJ��6�(x<����,_%�q�?:��zC�Y�³btKg��L3)����K�x���o"/yB�Xڷ��$K ���,���"5\ܭZ%���f��`XPu�}^|��.eI-Ԁ��q�*ߩ%�;�]1�v��� ��u^���P�AD�{).�9�c�:_ �-�����{��Q"���-�_棚=)
nv�N�<��<�}���f���!��o�#I���3*�g!���$���f)�KY�x� ��;��9�a�Ο��!�8��a~�]Ĥ��xK��l��|A�]iR�&[���5U������S�sR�1�_.�I^`��g���v/%m����,�Ȼ�*��t�ؕ���g��+lLW��5gi�R"A�fxMAt�s��B]����(ƹ΀��/}>�A<���ǉC�z���M�����8���2�;�J��(�� q�S頹�mI�',ݎ����W6_R(_(�MG�{����ƥ��4c�����қ���U���t���H;PE4��4w�V��{�3��#���s�����E2���Q!��R`C�(��j"��܈n����cn�W�M�*�6�Y�UD��!F��Yg{�x_��kă#(�v�16`Җj{iH	_g�Ķ��}e1Ֆ����(XqՄ�b���(]s���J �U���"��́�F�+IBˋ˓]�8"�G/�X .�J�7ZЀ��8���5O���y8p��DN�fe��G7?q<)ȉ���ȣ=X��<�D����9:�ԟG��n���o�#1��Y=��<�t�TBp��˳�]�e ~"~Xcu�`�}�:��؆Q�yD����>ZP�y�ѯ�X������K��|3G� &j�)��	9�2~�d'���"	�jz�w# 7v�،B� uC�2.)>����DFQ7�tN��LCW��	H�t��3ю�P�|�Y�<�Z7׌���1�-M��V��q�G���Y�h��A�y+�|�\�s3-��4������U���j��0�{@n.��Y3N�N��%�j#�D!e}�/ N	}@L�	eכ4�=�1��˚��{�`2�������N�ޜ���s�h�cY�YU���]Ԭ�5&K��b���M!�����(`�9��ixO��y���p:�=�����+�N�ee�#�Nm�j��d��H{BdA��@���� �.��M�Ny~X3��``�%<:�6��@�I]�S��� z��5�"�Y�u�o��eY�������:�U�f!mut���_�u��:��G�mF��O�С�U��=g�
������\��}Il�O�l�T�[8�%�	�?��)w���>��\5P��i�Vf�#��؍]ҥ).�7n�+�Tz�7ZpNwSyi��ěf�?ȕ$ 紋z�(����a���Y�Uq��A�J^��;�u5�m+�H_��j��WK��[ݪR��	����!�54ѷ&��8�b�j 6
�SI|��9� ��z^%嵊ٷ�X6���	��H�e���?kRY��Ĝ;zi8�V���52�n�.bˑ�c��	�coof��1�k9��lI�������A0�|DO��Ixą]6�ky�b���+"|c�E��_�0�exZM����
��i�G��+^�����E��
�|y�;o*���/3�����{*�7�֚�{ܻ�^@�,jr+M���%$�A.q|���p�����W���^,t\c��GǾ�mv�� ���<���9��H�>k�h�.EJn[�r��ԯ^܆ë�k7�������rg�k�+��b��33KX���%8��.�:)?�r�,����)��r�XxѹA�:/�����5��r����~�w����[���:gL��Q6_L�&�p���뷵�����t���k��O����aa�"��q��R�91�&�C�^�X]O��a~�U�M�
3^�&���x;�f<�XN�f�D�GJ� �����UH� ��΍p;ž��o�]�è�L���@o6V%�H��m
��s9`���=��N�#�9ڈ"f�����b�y����p;B��;�Ѵ�Z�S�Z��j��������zA����aU���'ʊH~�r�2��邎�J�m�{�V�!k�����#����G����̣5^5�́�Vz2E;���h+�%��wW�
�QC���ƻ�(��k��룴8�}�^T�G��XR&�q��BoΡv$
��,�)g�}��B��OW�N���W���9ڸ
���oR������d؎�����W�\�M��F4�聑1��l�"Dd�?�	�F�������*��8`��o19Џvb4�玂���e��z`��A������(�=�5o,�'��8ʳ�<n%]*\�ܵ:嚗g&��b8Z�=>�N�a��	�Lr��S����M�w��c�Φ�[f��X�@���r�����g���$#H�:̇�e�cf-����UF�j7�P����ATZm���1v�qn��^���=
u�&�<c�+ә�dޔ��k�RB�xs��'t��%&��8�S�WÚ_�i)!|�Ts��J*���)�$��M����Tހ�gԥz�Y+�Vq�ĝڜ�,��M�Դ��GVH�'E'�=���R��t?���֮��^L4�G�Up�'�>�,n^y�W�,�����'��496�b��������2��Z�����F7�:�{�SR\�9�!�H�?Zl�T#s�~�s��MG��@W�@�=�j�`�e�-QE{���Y��eh�Ny}�FX'�Szd��Y,EB���#���8�zRǇ���F�����Tc�M�B�˧��3Tl�s�\�b�6����Y��tŔRel� 6� ��i"Ak*R�ۜ��A�Vh.V9������WU��i
ĮI�=;����)RC��mDF�&�'!"�)�^�.�'H۔P�j�t�C,��ȷ�֕�tT���:�^1�"Pv�uC�G��A0#1�s�+����V�����?����q=�x�H����r��q�[.�6|%�9�����OItq�cts�'���e������JI�l�8ue&�^O�짡��G�\@����T�o	e��]ܙ&op�˩ps��==��J����J�������M�
��"GR̊39A;�x�Ί�+����Ζ)��r� �$�R�/��)��d����������>�u�G�,-4��0!��y�;i:���T��Q�>�n��� s�g4\y�+����K�W���S���T@[Td:���jA��7�C�`L���wS4X������XZ�d�yz-{ڟnÆ�`J�?���2�%�XQJO��^e���-��w�]h��;:�~������������~��S�!I�k�A�*��5OO��3�*Y��A�a������������O�!�;�����E�n�!��+��v�&�����EJ2����7���(neS����^�w��E��c�i�G1�Ŷ�@��4䢘���"��sS�u@��I�=���Z������\"C������uZY7g�H�fS9=o����K&"�fćJ�I4��C�C�3|�1~��Lo�t�6K�32x M�I�T
$�|S�!�E��$�����~7ě�Id����T>^Ϛ�(#�p$]�7��_�x'U��<�Ϯ=0���3�#ǆ0���9u�x744i�����>���0�{U�O�r�!���&��k� 
�@�u�cX �7��ΗƘ�̿�XJ���V�y�<�p;6��8i08�E�Q/܏�)�J�h2|���(nr�;�z�ډ�^)v�`U�E�>�'|��x	�y	d���݃mrV����?KÌ5>��#iLP鍕oy���479.&�8hM���J|\��ae�As�*�㘘������*��T���b�y��ӚW�e��*�`�7���6L�t?����%���S;W+.��*��,�L��m��?{q�D����
����X՞�=݁L���^� ޘm������:E���$^�����Vj���8g��9�������}�VX�ד7' JP�l�v��xx[��E&MnUƭ�0�<-�� 趆%��U��4�񃞖Z=�@;˙[�KJ����;�60��p����S(���Z����C.2l>k�w�H@��Q�ٱ��X����V8����e�TB������YS[�F�%�CA)�?o-�D���Ƈ]�S�4�̤c[�d�\�U�����B 4<a?��h!��	1"�[k�S��)ȭq��l�z5���v��	h�|o��nW��gY�8��p|��kg5�˛�"��҈���"	°�X'�)pԬ�;s��"�/K=]��ォa���3���z��"4��/���~��|���!v52ׅ4��Y<�.�$3�;�]:z��{�T�֯�v�![[ڷ����t�ޅ�h�qe�,�fHȷ5-ײ�5���+��ށ P�և{����b��F��b�*��|`��zb�&�o�*�n	^vwrE��P)*<�~���R<��p�_���<��I,�w�,w|�U�Ծ+Qг���)�xY�)��Im�L�u?Z�oTx?N?�Q/���#����+Ń�,MY����Ê���>�O���8 c��	$ +^0�&,}X�r<ίB��nF�&Q8vx�]@��ʧ��)���'c�s�$�;�'��|�M�}�~�sr,`�Ò7OR�,���'�C�����L�߀X7��1��9pds�-(z�(1�ϸ���/�~>P�]t,�F;�8��e]�t�5��ߋJ�
�*�~�\�3�F��k+��Xl��w]�n�GA�C���������:����m�*"���o����<�21�������9��Tvm�il2���?t{�>b�\G���p*)���y_A��~�^�T�FGur�8G�tL&�K	W�$�!�E�A��T�����&�����8ݮv{Z/G�!*�&fq����z*r���������9��⇓;�|�	J�ߧ_�z���3����3^�M�J/O��k�4�����-�'�*C*��|�b�?�CM�������۳�����Ơ10nb~]\�Mj�tbڳ���4�ݮgs�����~�@U�I�8wPJ,�g�Η�a���N1�Y-�"ÃwG��O���Ck�[��ڪ�cAm�dPr@v3z�;��(�Gb��p�6��pLc���᩽�z9t7p�=a��~k�Pp�ꐕ�����Aaz$���%�w�=��Cwl��!J{,�_���d��8 /��'��{�O�$�f�E[���d��]BiB4T���P���8���[$vW�=���R1��0_~=X�ϼ���͑6���è�B'�\�J��̆��~yAIc��i���i����]�y�P�˃�P 5f��܏<3���p�}��S����8�jmy|ɀ{�2��^�q�9L�jq0w�d`v���� ��2�!��.�(D]��k��#�'�w�!�V��Y�j��5��YάQ�N���W1B�I�IG��Z����GGȐKY� �8�+�(��3�z�4-0J�쬻ˌ�)���$'�2@E/Y��t�3兡���ʅ���DX���5�N F@#}e�~�Ҷv�1�!^���{��v��{2߱H�S���
��hJWp������
v���K��$���j�I����9�T�x��������N������#���de�$uN���0���_�[&q�\p�T��ɜC��N�X3�,S`��~1�Ҩ���I|���u ��������u�����X��b�ͺ:p5��ݷ���@�.pdu$�:���G��Fh;�O�����L�vg�aB�T���b\�/�} �"O)ޞTV s�|1��v55)�
��5��\W���a�VoZ͚.�/(�	�)Ec$n�(���l�z<��j�+��#e��� Ȭ��竡7d���J�V����yU�r9+ݖ�aUè��5W�y��Ut4�tj��K�D���Sx� ){�po���1귽�8W��jWlB�GT�|�Y�K��Q��lO��"�I�|�x	pkQH׭����`RP�z�s��i��V8�f5��3Q񻑚�e��BcF���x�-k�9�l��C�_�ι0��O�+dx�Ŀ��k����[T�s��|Q��E��!�'%`x1A��cĐ
3woi�1�҂�0���KE���
��jxH��+I?�D�������70����U��,AfMI���kG$:-qӢ����d��,պ�$�,K7ѳ}r��Z��'�	�V��	s�_K�>b��ǱJ%|`�	'F�&e���kn��UZ����B�L��&���m9�n��Q�����ʭ�ۭ�ҫq�E��� �Ry)��	-T{����ඍ�o�R.̄_Tx�^FW�gMf��܌?��\���,���ːY�t��vKAgb1�l��T�[7��8�nA�$��t��v�L(���/�ΦGZ/c��A�<J�$��GQ���m�Ep�A�8��P;�����S����m�o4�����_�A	����U���.ۊ�cI��Z��Ŏ��-m�L_V\	�ɑ�BFV��sS�M�I�+�R����V�/L;���h!⇴	���f�Qy�棼y�(Tl�4���9��}�'���y���0_է�=B�¸�,�F
���_��}v"HBI�DOͽ�N�K�W�����
�Co�5��d��[dN�����Wǖ�\��7����跕^1�r��-�d`�	 ���|�Ձ��������1/�vt��t�I�m��9��sÂ������^��x]C�]i�.А���]���<��&��$���=t�:�W�V	�#�rO�S ' �C�P��'Y��FD���B��v@^�Wr?��0�p��wT#�@Y���W��P����"�BPH���PZ#�"̧�q��a^��a=�M&,�J	������J=0k�굁5s�޻t_@&g�mO�8��vWy4����Z!���sP�� �~�{��Z9�M护��D>��M2��jt!��q��:��d�PzM�;����DF���'�/�<���a;?I���̫e����4Z�U��Y'���,��Uys�ڸH8��gd�ݷ�4�*\٘����ۥnmȎ~A��2�<�F��;���}R�ԫ��������ʢ�sY �i�ѿ�{趫Ήv��`�g`�\-����RS�����m輄�]y5zZ˪�zBF��#�X̵.�zهsX��J;b������BKݧ�TbI&�Je����"e��������v� ��@iX2*���&0hA��f.����S�i��W�ni�ծ���;Q���:�C��D�����.;�__��q�'�|oP�B5���C"l��mM���!�T;&��^��P� �uy{��^A�����,�c�L:J�����!��N'��g7!xI�P��!�ʰ�g��[����0�%��|7��ZI��Ј��a��h��_���щ�b�	u�^Ŕ4�S����K��%n� ��"�T��:/�r2^��jCQ�pt�ҏh����O�YO���S���{;l?\r\�H"{w�����6{a��숟��z����|4�'e�h'gH5pr�ܔ���V��p���Ox�z����?��Jw��+C�o��H������裏�`�����C�J����n�\}j���I���Q������G�H���2I(^�q�Gg2�X����I#��6葙U�A�24L_u�q:}i����C^ه��K`1�LL�8��z{��5�j/��X��u��O:Kï�E���[w\52�%��f��X	G/}7��R�IFwG�J�����%�����U�/�����nk��161�zs��?�Ĳ`�cqKz�ߙ-�7�����[�Q[�o�+e���0�֨��:T�'�Ӟy}_�f�g��m��?�K>F��]4*y���I�����fb�)K��TxW�����zX�a��M�z�18�~d����J����_�Lb��C����R������/����3�y��x�Ra��_��^9�g������ll�,X  ���ytx��iJ�g�QleBk�n����7FAfS�VtJ6E�\�{6�A�nι(/֜�A���`��T����Y�Ch	y�E�ǳ7��=C��� (���L3h���fm�Z,6�6��6�o(��M ������ւA��cT���6t�;s��(�M���A3P^L��AOQ�t�s�mI�3�K�܇���e�O�>m��!�B�`�u�cO0j��B�A'���l�n�"rM�T,6%���X8���n���C{�ڈ����0���P6�h���!H�#g1�����M1�����A�:սBS��n1]�p5�Z���͔���&"��Ɂ��o�d17��%]��"��/��0.�>�7S?;�����L�GO�W:��{K���0D� eҩB78[�<B'��-����l����ջ;D����Կ����
���ܞ �L�����V� ���e0b�����[��5��\]���er��J��w��Ѐ	���A�>i�p�1=i�5���f�-^�����TÊH��q�R��P3�+sŤ�@q����T�Ɖb��� K`�R����V�d�W�[)��zhͮ6�������T��H,0ͳ$y�S�:`&Ĭ�itQ���>��m�RL��g���y��1�g`K��&ʊBoS�-T�Z��/��~BmwX7v9�`x�Zg��S`~w�m�_���d �-�6�noh�`v�e�E��QHaQ�& ��+ۛUI-"���j+?�$���*x�ƣ��iyZ���.1q�M}]km��V��5���{-Y�9wY�$��-���¢Zx���Ͱ0����[� n3�������&J=T���2�~Y��y_��Wn3dS��쀊=K�@�(ȏQik�	��dq@,`��(�w⯕�W��!���ue��1q{Z˽���K"o�6�A�n�Z�gT	f���o'���q_"(y����4#�-���T|%�ǝ�*�o���tUnM�__� �cI�=�
�QM|#!r�{�����2�7pZ�I�	��n%�h��3N<#�:�$	�+�F�ջ$ҋ�=�{��0j���	�#�X�Z�hu�E4��x�!"o>D�[0��U�\�´>!�v�R�k����lk��6z�c��C������X�鰊ڟ��.�%�h$�;ⅅ�dh�ѡ�}��;��) �h��^���r�R����/�v�F1U���>�H��x�5��%�^76��I�0Q��k���>�#M�P
o%�x�9��ŋd&��O)�vu����e6S��S�E8�Z[9*�*�9c����Fb�e:"�*�ƻ7+��6�W�?:}��d���%=W�$���D~�Lm�m�ls?�sD�E��6��n�{�����L>��
4���ۄ��(���g1�f+5j^�7��P�j�'��dAq��ʡ����u�Ҹ�h��?M� vv��A�EA�x��ER�	m��\3���k �%����T�/�gZi�0;w,I�w2��t�؟bӺ�����(C�CZ�W��-lCq�nM�3W�Ռ��@cìX((��Y�8ogԁ�{7B�J/�EDY�;�FF�l%u�~U5o��߁ �
�3aSI�xq�[��\|��!$�Ep `�6?�4�hM�C	���[��Q������=l��e5"��vK[{h�;�CR��ZY��$���5%<���
����0\�������g'x0[��e�sY�����=	��J�
��aa�Rc�߀C�É�΁��2F�c��7�g���v@�U�1���.F^ �gM�:�Αç͡Ă��v�F�[��숭�B��Д��qR��XaHt�zYh���G~�Wj�-���`�_sb����ljh*@�K(НB��b�$po!�:n�vw�sq�OD�*hE܏pO]<�c�����[���0Pw�Ɓ|5���@����cQ���i`����)8�s�ô�!�ޛ��?��UQ[�5����#7�袁�n+�� ,�H�7�u�6�"�jxF/Z�8L��ٵ�m+��V�Ҩ.}���<z�|���F��8�G�]����3)�K%�S�s�OJл��Ӓ�רh�)]�ߟ(�`~��c@.�ة�S�C.JA�1�@R�_߬z��K-N1$��pv��Y^Tzs�����$�|��~j�Q] �Fg�I�2T���Q����?�v`
�Cē��"��1�F��+W߭X��/w	أ�s��A�J��+r�ݭ��/����m��B���E���X�2]��i��֯�ۘ"m�q�2~U?�>�>�G���.s��h_�߉9����W�Tv�u��G�7L�&�w��Б�!'����0TÈn�0�7���Ŏ1���)۽k!V�fX��%�VrJ����*�5�Ӯ�{�����5��S��=�N�<����M+t����՗��u��1i�-U��V�����b��C����:�V��%#��M�b����f�0+��b�^����it��a�|�`;8�ZH��t��=�;[@�4�dߝJ�(b����aUw"N]�7-mh�N�Aw�}�{XY���|[E���V��cmw�d�� �xd����(CM/Gʎp2>C�c�p�������t�F�=�I�~��p R`�1�b��a&L��-�l��9=��#�����'e�D0˘��9����/�]��S:Z{5Y$ ��E��	�/]in)���+#��^�2�?$�h��`�~W=��^~i���{C��*62�h��HBӤ��ve��2q ~�ZcX@���q�8~�؉kLy�9�˯�T-UJ4��P�&r� �͎Ij��sw���v�|m��  +2��BðD�Q��d������mW>�yk��2Y��^e(>�!�.1V��x^T��V�\d�G�L�Y~_֞L��+<\��'��3X��4A�i怊�ˠ7�Ra;i@ٶ���3yBM����U�qDl�$0�N��@�XOe��2�J�R1E��{"�!�Z���1�EM�gʗ�=gh^NW�D�l������K���V ���3�쳥�9��kx��Q�$�\�����n]�ʠ�y�=e�oNXl>�DT��S�o/��Cy���AdߜWI�Nd�3�`sy;E| �0+I(�ӛJ*} ��� ;��Cuu�0�
U���!��]R:>d���a`Wr�B��u��:�sAGm6F|UnO@+�,���l�g�e��H߳�2>\f��}u8O��rTjü�W���)"�S�I��\�&!�W>��s�ͮ�3�á�7�)ّ�n*���gzPv��f�ޖ)��釛�}}�@Z��v��t9��pp�����U\:MZ��*��il�p�5k�"�-VEH�ej��K�lF�U~?��'��� D��Q��8k��j�5��[Pk|1��ǜ���[��5���\��P5	��H�}̑�a2Rd���t�iR�V̸G5�����e��.���<*c��7��kd��l�3{%��1�0~��O��x/4��k=nR�풘�q|e�	EP�;�Qx���w�n
�oi=�����Ec�
�?&`��5��S�Ҿ�f��7DvN�&e�i��,��WM]iZ �$'�,qg������l����A�,�����/��O��;ņ�<����i�>vZ˙�`J9�ӝo�:���>"k�qb�+�v�����P���Y�^
�X<�N%#A���9ɭ���}���T%�E�r�*��DY+:�lD
���vr��?�&~Y˼��\,8R�:R���w�L����{���4�6�����<֌-9��:�#� 
a�F "�z1�&O�9��&�֦*���OFD�a)D�X&�3��U�;G��<�c�Q�
Ӓ�] I���HH� �M;;�w����׍�X�L�B��V0�HT]`m�dd�I'�9�����$�$��r0ړ)7�j���-���%P�pƱ��a�e�˴a�S�g����f���B�����#A~�d��Sl�w�̊S;s������m�ƞVѽM��������>i�h:W�[��`��W'�Ve��;�h֛`�	��ur�Q���Vc()�����^�N��}`��R����a��<�bB3����
q���t�A}+w�B���O�,Nr`$W����Đa
y �o����Fӻ��dCƅ���W���\�_H�1w��1�1����-#d 	�]���:P�Ve;l6P�`_1��vvm�Mx�т�����B@���s�����{(�ʭmG=���cG�ǐm]��'��E��&�W����=	����dA	���r�A3S5ף��4J�1���zu�&���8��@3�fr��c�E�ل\�#S�����#�.;��%���y6U��P];��B�:ZxҜ̜�bq9	�^�V5=�V&x��_���i�ޟ�^k����J�ks��t4��&���db�8A�%W�QV�Ա�!GI�sD���n���o��oBwM��5�����:��E�\V��q~dtڇ׻e��M6LG0)�VK6'�̨Mg�_f|?^�쁡��%��4��U;�'��,���y�^��]!PB�2�I4����-���D�8�CAˎ�	�G�C_��FB�~��BR'tu�L���eF�?�>s4�	�H�X f�Q ��ەܚ`T��-<}��'�ӵ`D)�Y-Z�O��-z�'����"B��V#E9��\�z]V1�hH"��)���`jvB{-o��9MT���g����ܽ�~�Ȧl������� �P�i͐e*] �jLA�
�.6��b��ްMW�)i�Լ�T�O;F;�sxlC&��DѮ� 1�t_Ilt;'S�P����?CW�}�BI.����TPk����^<��P�6uC�8�RA�"�^9��a��'D$��r��F��V�x�f��b����m[���#e%���A |��e�I_<G����ѺX�����F�f����Uu��^:��h�љ���5�9�"00۫o\�GG^V��C%�p)��������Y�C���7�0����"`Ǽ�8)�;|&Ǝ`�����ݚv�JRp�OdrU��`W���nJb�DW�VXA�_����LC�$>wG�$�P!�<7�lE�� D�_+;�d���B�(����9:���lZ�x���hu��������'��m9�CP~�QU�:�\;)�i.ϫ�	,Q�E
o�Vy��x[ ұ���H�*�Әo!He�u$���Pf�.Q�B ���E�ݭ�۶/�f�z�c�[�?�틧���������<r����H�>�zm���^��wH�+�+������̦�Ǆ� � E��X��>����b|���!xy_sf��E]�.AdǏII����p�+y�s���9
{R�'|��#.-.��PJ@��Z_�"�igM)}�{;X� ����xŌif�U�Y������
�V�>�y��<��ϰ��)�U��c'��'fe�&��/�ޒ����H�Gh6���)���7�<?X}]	�0/N�s4��Y����	#���fJ�<Y��6�[-��;�~��z*�a5�	�X�N��w�#�7Z̟��ro�J-f��MW{�b9��+ǜ8�pr��q2�B�h\��5E	��Q�����%-\��H�Ů�>�M�t�xJL9_+��N��-R��E��="_�U>��B/�xt�J�z� *g\���C�ڤ��ŵ&*��t��}b����(���qж22�푤 �IW6}� �ǆ��5_��qO1i�@��C��D�WK��L�C%��*��F��/��PX�rA��,xK�>��zqɝ0ǽ\���%1�Rf8�X^^�},�����I{�A�@Q����%$7��x �������q�fO2�I�Y��([c&6.�-҃��0u�Tx:Q0�O������=嚋X��k�a����}H�}f�0���T��ث�_�*n*|�n�״'��f7exK'i}xl��a}���a�����8	�0�R�rx���uκ�3�-y����[Ra����_Kc����mF��?R3+_<�W^.�g5D>��'{���
,m�-�x(Tt�]��^t�gJw=l���C�B� TA{�K�*�t�����Dx�v��Ύ�/K^�Aʞ!��M"�Β�6X6�>^���[�w����r��k�%('ԯ���4���mWK�,���Kl6�,�(m9�Mą�m�����c��7��[����c���B����H^P��/�JS��鴔�M3;җ��?h�Z�x����PҒ!�B�`p��x��jpQܖ	��u�6n���M�C6���#���sB�F�{Bx��V���O��Ģ�6nr�8H���g����t1�o��"�uv�)ՒQ#�SX]�D�ސ?ʵ�
"D� �.���9E��YI�]���";�z/���.��#7�z��X��!�Ob�R�j�m�#D\GpeǏ�7���<wV���Kh�q��櫰Ҋ��D�������bJ��#kw���:�k�2V����P�mb�)��z���66�1�(�h�1�Ի(��
��%�M��L��\pTT�=>q�k��&���֐�;*��δ�����<$R��3Z��ŹI���d��Ė�(՟ifP ��eR�C�Jh�d��1lڬK�ͣ�ȟ6����R�0Bjhy��K:NϬՇ�Q��m>�����d!=�g$>Cy�y־�K:&�PcS���T!�eu�����\7++c`Ͷ�\�}S�gآkA�Y5d��K-���n$?p`˚��:Q�枿Q+P)��{)��Ra-7#����y����*[�_��`��r�� �b[=k"�^�F5�xt-�Y��y���.��բ��7���w��u�u��9�nܑ;�L*����&��|�?��2�jG�]�
���on�S�)���#�����i`�ʻ��T@a�������eʕ�I���ޞ��0��&�dZ`�����+"DS|��$�Z���ga��f�o����,^�"���kT�48Ӥ�|z~E����oYw�t����4�# 3�I��|
z5%|�[�!g3�����ov��7�quI�%O�Q7,�Gy�(#wC�$>"�n����u�,��0b0l�v���X#�����8u�pz4Ua>�6��>�U�0:�U�p��I�s!�d^�'(k��.��@+�ĭ�ϸ���8�.׍%�X+4q��0�!�}>;���[,�/�����pA)蕬hS'���70rT�?���]�{�vH(�U� >��֟����]�^��F�%�_� D5�� �>���#��P*��oڸ]�c��9��R����..�K��-8"ed?��D4�M�OM�*���n���z��ӻF�eO�N*?�7�J6�n�?�r��)���ӽWL�p3�L��8VLi~�mu�k?<.D�R��Қ���j�
�ڞ�gL��������Y[����� �f��@w!^F�H�mk&j��i���u��.��\.��K������ ˻B�����J x<"E'�(v���q���J� i�%��o�l�1�d7�Z>J{;���͌C��)w��}�	���Q�(xގZ�$��dSlX�{̆j����Ձ�ʧջL������+58�sP��5BYHച�Y�z�F��;%��1*�AoN���5Ψ���S]U��m�?[c�\�2.���[ u��?��h��T	�c�[,U��W�rul.��57$9v fh(R�8�����Y˷P�q�=��"5:�P���f_��f��aԐ��h±²'�u��Y8sl��=��g��ģ�a�B��Tk@�#�#��ݫS�X��̵��C�v�}צ�B�n�.������:���<N%ķr�v�@�[���¼�y)\��~�q����P�H��.gt�V!w�lr1��h�W0��T�ubO�����=*����q�W,�bNkovēn�'�w3C���N*=N:��r|<������e�����wX[z|j#���H5n�Q[Y����[)-��.o�V���p��?o�Qp���}c�#���v�;+��,.����ë���ٞ���8���] ��H�}�d~�7�T������9F@��r}!��.�W�e�#|���;Qj�ռ����ĉR��PF���KQ-Z�����Bq���^L�l=>uy&AC~�HO�r�[����k@�)���sl��t��'&�)NM�8JKIW�����!���s�;;�~�Ź�ÄXt�M�%ώ7��;�n���8߰q'�I�P�S�N��M?�?,�.
���Z:'s�[��"��(��?Gs��:�N(�4[X�U��>'HLB,P2�y��иF�ZY���[��4��ٖ�+��j��H#���b�0��hxFkHt�/|�R�֨��Ι�s܎L�s*��'��������Q�t���`�K-�q�A%�i��������[�Bz�_ٍ��B��|��z�\[2c }��� B8zZ\٣�+8R�@��}��C<hO6�b�F��8�)9]��Vʁ�)!'��1Fs��~��Au���C����Mm`����d��&��&�C����_4+@��Z<	�$)1R�p� �G�z�-�)�	�j�4~n�]�^F���� 혹N��(o��zO
����X=�MEFf#+E��XFu_ww�à�gA��-��F�M��pEnm������������12�2��+���6ۆ�m{�]2�>?�B�>�pG��xȊ�����_������.�T?ȼu-^G�EOL@Y0���ؾp�!ծ�[�.T�(7���YNo���ή�ӂɪ�!{�f�8��Spr8O���\���I��<�G���>��Z�����9*m�<�����M�MY���9�E�J��_�-C���k����b��C����T��ߧ5כ�P�����0���b؝��kt<��1�1��a:�H���}p��6ݞi�@@��ˉpJFϑ�(/�aCq�N�I-ە�|w�w��׉)���]�j[sK��D�c}�dj}�С���87(�y�G|��p@B�1�!clD���.˵�4�tѣS=;D�~�(opN��nn!�a�#Q�[�K����=Ʋk�h����������#��/�ֺ���{���$N�E�w�\��P�i��������*����$�J`��b�,ch�)��~�h�iة�\6�Q��dB� p�$?F̠�~�cF�K�nr�����طO�y��m�]�MP�����)L6�����H�ح�q�k��jGY�ɚV�2/P=����j�;wT@bvI �.� bH2���Ȳ{D72��M4�}$��!`�n�sS<�?��ğY�~nk�F��I1��d�����z�"G�Gb�VY�S�R�+2��Fk3�B�4G���Fӄ�&��[��ADc@���i��3��(���1��3D�ov��N��@}�6e(�Ґ��1�U�r!�{���Ѹt��/�UP������N�hd�Қ
O�`�(��\K�������W�y�x칅�9Scgx ���jԂ��]�nBH�P�H���,eJ:N�Y��s��9d�uH�q}�
 ��'b�]u�N*��3w��`�oZK;��ʻI��=��� ��L����*� u���o����E�T�:J͠��J0&���1u��:�~�G3�F:O��q�2��K�gi���f���\,}�}��O�Tp���֛-��V)hs
�O=a\f^�5�8�0�ʹ/|��L��:�)]n'��P.�z��ፌ�&�}�&�7��Ȇ����F�x߱b�������U"��ө��p
)o�Rl��5�h�sI?NL�jI�=KY�ݛ������^�������8q��j�x�����|w��1^ī���$U��%����	�1�Hq?��S Rj+���i�fV^�5��Re���|��t���	�c����M(k�l�'A��h?0�R�O��x��c�w�k�����,.���|��mE�#�A�x��ڝ��-
ǣi}���E��Y^�E�� 
�-ғ�{�XP��c�,37����l�)�oW�,�k�M�;qf/�$-yBq-�W�A?���Md��`�,����M(��cX�A9�������g�9��>|�[�_@�J� y��^s�@��tkc��q곷
����^��AӤߥXB1Z%�f�sQ��+��ȩ�Pz��r��J}�:�L��E7�&vKr���I��~�[��
��>#:��"��L�eo��є���/gć?�|�3�� ����a �"�}M��(9�m7&%D�0���ki�O��Hao䒦^��3�᧲��;�	-<������o �,�a%H�§�v�;6��� 51�t�Ll>S12�V6տH��mf��ڏF�9�엢S�k��8��\ڙ���0~l�r�kU�p�_��s���;����uS�����r�E��z-��(�ADd@�2��ɽ�Y"��䪡&���V��m��NV����dh���\���.hhBգ��S�]��V+*W;��4h�����;�Q�*~�7�n(/�E�oǴ�f}�g��X����[���)�By��lN
7����<}q-B�8aO�sNN���W=����"�
?��o#���⋻�~d	��x�WB�t\�����D�R�P1�7�3�!d�+�	;���o��\C3�2�qmش1*]{vs_�>t��d�50�w����G=�m���������.U�i������J��v��a��eXʅ=�@J��TWv�V���_�Ð�[���\wX$A�e��}�l]эOj_Z+�d��1����Ih9ǩG��?Elɨ�&��$����*��1R'p͠9���~X�������KX;�=5��� �~�g��&n A��G	YV�~�e���$�������.�O� ��`E�q�
�g���z��[VqN�:H���B�m�c���W�>�,H�O�z\ƻ���,�&�+^,%�^ޠ��ǳa��/����:X������b��Ԑ&!y�U>f�1�ElA+.0�i����Cc溷�ss�:�GX{��L|���.����?@��_q;��vq)̮�{j�� �I"͸�1�8s�U� A�ni�~�­R���y����}�ö��U������'�rx&��/ g��O�7�wG7p�{N6�`�u<�d
]XW_/}�u4&F%�H1���.�	�,l��#�<�j�ү�Ί�!�J�іۥ��0��	i�^N��6ے��ZT$��չ�Y������{�J���)�+P���{���T���chk>�542�� M��z��c��mQ�/���m��j#J;�f+�eK����@�M��)ǎ�3"�q�>�� J��k��.�\A3���o��m�������)���\�{~�(_"�q��2P��o"
Ig�F6�����0��_�� q�Mh��jjC"�}��#�K$īL��,�����.k%/V�HXWv3�$��K��)Љr]���\y�%�w�f��rX�`�}{���F�]I�j��┓ǀ9%���:�/�����H3�2�r�u-̲>S} �vA�c�D��F-!��_McV�QI�oA~ٜ������ױkN̞=B}W^f�O<Ǳ������G{�!^�*��k�����6��f&K��x���N�>�a�*"�>�8��{o"�A3捵���IU���uy�7��R�sw� ��R )�w�U���1R��g_��-^}�Zgd׀�� �j�S�\�,���t<XE����gy�;l�U��21��+ZA*�uU28t�i�Ҡ?U���!�}(2/�Ay�����K����=:�XM4a�	5��F3�x����l(����=��z@�HmFb,z�����6<�4(�/�Md�0�I���t�<�c�:��è�����βƑ}��V�P�s��_U縜��1Z�3�t��K49��h���_$l!�ֶ`���'��j�Œ������n�y�M$��6�.���h��^���6'{p4*��������2�6]�HF�9gu�]f~1�S�Q����Ձb��"��]��n��$I��/�� ~�"sdm�=Ǐ�(�^�(�A][3�"���/j�L.�U7��������O1x��������D�5�eL�7�E�<�b=��ٯ�@� �q��Dm���f�֑O��2�����:���6xV9jw��*b"���NF�ɀ� T�7�ΰ��f�_ļ��v+�����"pc=w=-%�:�<��W�q����e ����R���3)`��hܞ���r�q���
@?��g� ���R� 5���d�����r���������e�
��S�ڏ0� yr�:����Do�Qݴb>�v�'�D?g�"0yy�_��dWK 
���S��T0�{T�����1D�7���`<�����S$ر��HWd�H�-k�Mn��`:��Ô�[�Q:�Ժ��<��T�-�^�������nFi�:h���w�wu�r����]k�l�)25?�?H�#��Y�w��QH��xᢞ��b��������Xn˒}�I8��l&������2�XJ���k���n�bS���N"s��@M�Sw�i��B���@p���A̻B��p���e+5�9�uS�Z�萹��#"3�szT���Z�ZIpgЁ8fC��o�f�;�F"ӗQ�:�|4����3nv|�Z��no�+\t����#S� �?I}2
	��|C7�!�||�9���H����N7��(IT�m���N"��w@Y#�uW$M�N�
�J�hF���9o�I�0ۧ+�# �#�{���O|u�i�4$x��墔>�\10�d�U�V��xW�!�?���k���0p��S���'d�·��׼��X:��'o�rxL�,��;&'M�(2�(���A���5o)�h"[���Tr����jkd��5�vw�U̘O>����G<�i�������]�t[{�/�Sc>�*�#Y�P�*�oiZ3���t9��(�=���:�����e���������m�*�GZ�}�iӊ�[e�>*�{�7�\6<nU?�[���8����W��↮��7�L�NrmĆ�?kրD� ���A�вU�H2y�-اLU��NR�ވ�
�/��5`m��D^�����9�j�I��(�:�)�����Ջ�w��F�<׃E :���\w�	0�xK�E~E�� ��� ���%�7���Y��sadZ-��;�إ�;g�����&I�`B,����(���Z�J�3]�l*�[?��P�����f���:���`8��U��B�B�	��YCr�F
�0%�����o�v��x�w�S�*Ҽ��[�I/\�� �gg��L $�?�hz�	!t[[�"�ɜq�a\kl��L5悺v�<h�E���Ug��,Yڛ��`=ݣ[F�5�a��΋���X�>J��u� �'���Ԝ6�s����U=MF�m��a����#M�����o���d��5������[vƑ�u���I�Z.�O��+g�:	!��kh�����v���[�V��qVr��2�X@hqU�x�*�H���Hv�% ��K/�q!���m��f$b~aw��e�*B�l�l�D4b�!�o�n�ԅwb���C�*,-f��/$<�Lp�O����9�Uw�q3|y�����Q����e�h��)|<�]��e�_�C?>��Q�y�Ϋ#����I�+���,=�����z���.��sgT8|���Z�+N1ư��}H��<�ޓ���F�ѩ8f�]0�ʗ��)�^(�d
s�C_�8s����l���m��cg�`°��'@%��Ť@Crc����y�S��p=�H�1耦pTr��Pz��u쿑U��& ~.%�]d��F+�/�vT.�dZ$����:�n
�Ź�n�Ȕ#U�F�p�+��bX\}�wM���7��A���i�������Ƙ#m��l��/�u�A�,�l2!oϑ�'3��Cn��?m�M2�5�?ds>RuKG�E��`]�����_�� ����T�τub''Gʊ7LA!�;���v!�!�1�[T�f �t��oI~��K��f�<��!ifa�����r�5���K�y���C��+���nߗZ��Ӻ���� t��#Q�M�5?�^�[���v��z-��͚�E��_lb���C=���M���j����Ŧ�Z�����0o�]bn�F�=�tR��$�$��ݞ����r������@Eő�(��Jv����Ua�%N!�N-����w7�T�?��3�[	�ښ8�c1r]d@f4��+(
�GR�p�/���jc�����<��j�*t' =Q��~[1�p���u�$���aj��񺱫v�=ܮKg����k#�����ʹ	6/������{y�O$�/EK���)hs�ei2���o��Ւ��vJW$fl�-z�B�{���n~-	߿����z�6v2#Ø�OBo��:x��vܵ~i�c��1��F)�|���M��y��s|�P�g�V���낥����m��C:����<j]���p��2Œ^NH9�)ɍjaK?w���v�o@ɉ$ ��2u���>XDM(&�[a��W�gW_v�u�I�%�Ֆ��E�Y�*$A汌}%122WԞ��M��+mG��Y�m��(�l+�qêy�3��l4�����|1�q�_�@5h��3պɸ~r�����DH� �bN�F@�3e~ŠҦ�1�����{�Y�<���6Eߡ6��C�n��� h:
G���S��9Ŭ�2K�I����:����N��}�9�URxv����E�{����������Ȥe췳N�� � �$�O
�K���\`�Q���f�3YLN��3�+Z`��e!����Is盦J }�"�|�H�/��6ce���P�y�=A�'��R�	��r���Sm���0��P��2N�^_��pq�@k�Br� ��}{���#��*Pm�f��]vA��h��BP���z��Z��N���Tqq8�^�lR=��&� �������}r�׎�k/���j�s�tla�&��%38y�]WÓ�J�!�3s|o���b�(d����MӘ0�L�*���}M#�#Sq�i-ڿư����Mn�<;��^���'"���I
�ڗ�z?�z���!�]?�4JQtUs�'�<,�8�y {�����L��j:>4��0�e7I�|J6�{nu�+d��F.��"Fz�l�s�R_�
ۄ=6�K�w"�sl�W�V������9�C�'�ͲM`�i�-t�O�_Ľ��vL�������*J�zǵ	�C�B��T#>���G�z��\��������C�$�w�B���uTO?�������~��/b� �Ӕ�@�# D�i�*��6�S27A��.n9��;���QW�Ԕi��Z��#�;~�z���GC^D	���J�Q۬�>'��P+��wA�C���z6��/,3T���}�^t�mP�KuF:��p�dA�o��P;�N��9A��_ű﷗��c9���;xV���>�)_�T�[R�Nك%�[|�yN3��z�I��
��������/��;�}���5��ٳu(�^r���"��)���M	�"hݫ�T���^��C]��paR��t
��9/Y����$0�²�ZDѼ �o�sN:��y���)G�ҽ$J����9DL���΃��tmJ�jW?�gV�@�_�x����:x9w�`$ʒB�t�
lH�8�8�__cيd�bޱz�p�6'9P4>�9l����S��ˊ�&Z�=�r'��9�^~6�����ba�vf�Z�A�ګ}(؎����)b 
�}�0(7b�G���4e���$)�툈i.��� �>-E�tͲ5B��z-P�[����Á��D��6&0�t���G�H#<z�7��W�����-+_�'����Ǽ���X��k�X��v�$b�_��Y��y���f��E�_�.yxH���_����c�}s<5��0��{���|��.e�Y��@,L�_������)��{sn� �������qU̑���ӈGyt�;��By���  ��	U1s_k�'��&Ʌ�/)e�1g���	G��:�W�	a�<w�P]An/�\4O�ց�1y�'8	[c�ʞ+�<���E�Γ#"�sjܖ$�?�� D	��N6fa�[STZ=�T�#!�䂢i��i�{�9��ԉ���Б�������h�$�5}���a�����]6�6yS���v���ioJ��2+�ғ��9��g�u
��-E�z���J̾W�X�G\���{t�6*`���m��S��������(�Ayq�w2�t�8u#IPy�6�ɟ���?��_"X�q��0�x�CC��}¹��K-��L�����/�~��i;/�tX ;ü   �  �  �    �*  �5  MA  IL  vW  c  un  z  e�  g�  ��  e�  ߪ  !�  h�  ۽  �  ^�  ��  H�  ��  �  ��  ��  7�  ��  � 
 a  � n$ ?+ �5 1> sD N kU �\ =c i tm  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+E������=\O` X��є	����bʉ�)����"O���i�|���mK�!��"O�d���,�d;��)_�����'����d���B!�$ʛ7(��E�/D�����  X^�HB�l���'�1D�0����30�!i�K��f]�T��4D��Q%
�FѢu) ��5���2�1D��KS"� uxf�3TEJ�;F���`�.D��yD�Y=u>v\c��G	c pp���7D�h�i@�ZT��;� �x� �y�*OT�PM�I<2(q�NIv6=��"On)� L\�O��93p.S)|� Q�"O8c�Q��4�b��P�����"OrxJsi�,�ىW�R�.�m���'t!�$:Ha�@`�H��
��ק�4I�a}��>1�IXyZ}b%� :���a�<����(�ya���84����X�'t#=�O9ص�� �@�npQ�jV�"����
�'P�ݣ6�x�� ��i�<��-�T�N��~2!�?c&Z8��d��}j6� c����yr�T*Ww�}���t���#2�\
�yB��3\�Aq��m�|8R`3�y���7y��	��
�W���A�ѱ�yRO��hݫa��%��l�CN���yb�ë�䄑sH�!_����ym�=9���bcm��1$`A���yrA\�N}����xPra�R��y��F�HG!2�f�(|�j�rp�̏�y�'���jpMڿ#?��Z�g��bE�O�`t(-O��i7a��fa\���ߧ}�dP "O�4��gR7\��SB�ڪ �`x��.�Ş^b,KE�{�|��#�[�.d���]���01���"��g��&�4Gxr�i�ў�=t%���A`H#h�qt��=nC�	�	�09�!�k�*�	�L�'I�����~� M-W���A��E� ��䄘�0=9�Bk׊kj��v�	U�Z�k#�=
���0�ON#W�S��l���h�,�0�P�pF{*�n�'��5�w�7h�����F�Y���'�:����޸1�c���<�DO>�$�S��($�����3k<�
�KL�r��C䉕A���cÐ?��ٷMʿHD�C�ɨW��BR�K�����M
�+q�#?��)3*�൐U�JK���7!��$!��C� |�%:�W�hA4����az��dMSrd�7�V�+,@5�&$0�!��֘�X1	�-�`�!�1��p�O(�=%>���ˍ�j�0�����
[�v,�e�:D�����ԣP.�yTB��xQs�a7ʓ�<��!	?;=F���,��2�!y��Z�<1f�լZ�QX���*�F	��Ӣ��xbӑf��0�WEE�@W�D�Ν���O�#~����i垼C�� S�<UKU.S�<QFf�6 N`��9�Ҽ1ta�����hO>���9=�:E
O=|2�JQ<D�|�0�ѷ
!^�:qi�-5��jE9D�� �,��F�X�`�`1G�=W�tt�"OP͹s�G&�6�XP�H�� y�"O"����Y
I���Kekͽv��h�"O�K0���	�>ղbD]�%�0=H�"O�y�k߹g�֩�BJH6���RQ"ObP�c��P�D0q�E9%��eɲ"Of���EM�a�����:`"ONU���/s�@ƈf�(`�"O���v�
0�,��b
�]Z�D��"O��B)K;��R!ռ:O��"O&4��/�4*%�1:��0Z]��g"OX��Š_�6lI��Z.MA�2�'���[�S�O��)"�
�T��4�~���"ODz7M{���1�=^Uۄ"O�8�R��w'�K�1$"U�d"O����)K��b��܀ι�N�����O�ZY���6u���X��
%l�C�	1��I�뉋x�����a�<	�C�0C��{A��\Y{��ƿ��C�	hӾ@���7Da4�{�D��C䉊�QzEM��|v��@�M�*��C䉕j�PE�Ӣ|\�9�m
>|ԾB�	<W��� �"@n���Ș`�B�I+�j�c�.P�2D�����&��B�\�@��ЧHn�)��R�&|.B䉻;4 `�Z�r�n�j���9*B䉂��!`�N,i�P���`ٰ2NB�	k%6%`��f�� S� �:P$B�ɭ_c8��g��b� $:ǩ�3]��C�	g�͛�d~|��KJ'D�C�I �t�T�*���g�	���C�	�ss��h�����a�`ƻ ��B�	1e���Λ<9�r5k!ƭj�C�ɉMW�4�J�.M+v�6	����C�3J�	��銚A�`���@�	���h�`�*%(��e{ޤ#���vh!�-0l8�` �Q��p��6
q!��QG�<�0V�T�Ai&(� �3Y!�ҥQ%��B�%O6Xa�s�B!��-�L�eDn���X7*�0�"O^q�r*� i�hp�B�?PR���'�)7΀�y���ր�?�~���'�D
�+Q�_�:��v/E'f��'<e؄����(�f,APR^���'�jdR�Hr;��?ȐM����V�<��`,�"ESS��t����0��R�<6*�b�d��!��S�Z�� LUM�<q��B�OҕG"[u�tW��I�<��le�����6�
�xӪB�<��E�r"�!H�k��ʣ��S�<	�˟�eX��p&��E�����O�<���Ǻa����Cв��=㷊�_�<ɵ�F����s$�%pj�JD%Le�<��@ /�����Z��Q�S�Nd�<1���F�q�(�X���Hd�<	pfС=�~�[Q�
!D��!���i�<yk�H��1;3��'ʾà�Le�<yKL��S�Y��j`"�^�<I�h�+�T��IƑ.�xqj2(�Y�<��+�1�5��Γ�9��@�W�<�S��%��4c'/� H9��E>�!�q�րb�+.j~��Ct�@�T�!�dWez�K�N�$xs^Ј2H���!������Q�ۖ
���ZU拶�!�� ^tX���}æh՝GF~m�T"O��,�y��3'�� <
���"OF��֌V!r��9ȵfΝA4�=Y"Or�Jp��.~�ES�Ĕ
%���t"O��J�]=x����kڛt	ԝ��'�"�'�"�'���'�r�'��'�
$���#�X�0�ұ9�Fu�0�'�"�'��'T��'\2�'���'����`$��e20lȕeP�P�')��'y�'��'RB�'��''�1�QΆ��=Q�,Y�W�~����'���'���'���'���'�B�'��7hΐS���(]H�l1Y��O���O$���O����O����O^�D�Ot���+Xˮٲ1�^�eI"5Xo�O��D�O����O����O��d�O����O��C,G�c�NH�4��=��l�&��Ov�D�OX��O����O��D�O���O�%��`�#V6027�O�i\ѓdL�O����O�d�O��$�O�d�On���O̙i��ڈ��}� �I3%�`d3��O0���O���O��D�O����O����O���!*M
���F�I�I:耊�e�O
���O6��OP��ON���O����O�|Hè�4J�.H���dZ�P
�O8��O@��O��$�O@���ON���O$`��Tv��,*q鎋ua2Q�M�Ov���O����O����O��$�O&��Oj�Q�B�KZjx���<b��)t	�O���OJ���O���O�$���m�IΟ|��"�� gL��J�<48���^���O��S�g~2(l��ĩ�ޔ^>�Z�*USڽ G�T"8�	��Mc���yb�'�n0��C۟e@� �D`Ps.ԓp�'.�i�W3�֓��̧?	�Ԗ~�Gg�2)pbTi�@�!Df�=ڐ��A̓�?�(O��}
���()&,p�`�ԛ6��I`E�V�yƛ&�۝Θ'��2$nz�a�#+�-�bt	����=t��t�
����	�<ɫO1��X#��`Ӑ�I�G���4��`� b�H����<��'���E{�O�B��`�ډq�N?xd���Lύ�y2Z��%��ݴ�8��<���,�1`F��O����J����'J`듌?a��y"[��pA�48�0S�H��1p���"�#?�thn���e�`�'til�DƠ�?�An��p0��e�U��u;�D����<1�S��y�H�1G��	�K��?��z�,��yBau�ب���P�ڴ������q<� SzH�\��Ɓ�y��'���'pT�ӱ�i~�I�|�a�OA�u�w�W&@0�s'�^=�4A
G�Igy�O���'�r�')�Q�@�~�Bu�@������  �I!�M��L<�?1��?�N~�xn^�*�������A"O�3�$=)2W�Dj�4Y?��&4��)����24f��2�[���S�a0!#^(Z�*�d» h��u�2�ם?��+��I=���r��G�'(|r!a^EA������|��⟼�i>��'��6m�M����WD �6*1� U��Q�����?Y\�\��Ϧ�۴L��4���(W�,PsH�ݲu��*ċ�M�Obt�A��������wH�&E81<��ۧ�L�(s���'Sb�'���'/��'�^��.�%DU(��\��h"�K�T���O0���ߟ,���<	q�i��'��30h�)}|�,*���njN�Hמ|��y�T�nz>ic�VЦ�͓R�r�� ����-aD!΍<��ū�A��E}��A��E��>�#�<	��?���?q��
'j�5C��^�0�ʝ8�홲�?9����B妥�@��؟x�I۟�O=`�r�G�D�<��7��-�����O��'?��'ɧ��1~�qb�����	H%C�Aq��aO�F��7�A`y��xݥ���O��ӼK��D�\�Z�"7�8(�̄RDj��?q��?i���?�|�+O�]n� � ���+����ƅ^� `hO�l�	��M���D�>A�wEh�[�/�#S8�AuH�y��as��?ɵ���Mc�O�b����[�Xy�bҹk��p�M8I_.	�6��M/O��d�O���OH��OtʧR$���%l�(�h�QЫ�It�ܺ��isLZP�'��'��Ob"m���ǱT=F}���E,4��0��'�f�~��Ǧ��<%?�;�CΦ�̓,���򣌔 1^�� ��zb��Γ<��	� c���'�7�<����?A���8��0j�']u��J����?���?�����$��q�b�S���Iߟ�s  �2&�B�dWX�qLT�&�	���O��"GK�|�ōC�"pa"�۪f���E�����H%�M;7\�� Zw@T��?y���o���!$������R4�?9��?���?�����Ofq`#F�P�v�*�W�Ii*�z���O�oڸ<%����şش���y�H�e��h�2H���M(RI�y�'C��'��I��iV��?fS��֟laBB�Hq68h�u�3F*���S�<Ѱ�i�������ȟ��I֟\�	�HS�����:8,���l��e����'Up6�ք'"��$�OZ�� �9O�D�����H6$�� ߠa���Kc}��'y|���m�z ΄:�eBFt�t��+M�r]J�5�iZ.ʓ_hʔ{B��x�'��6-�<auc
81ɈB�۳_}h�p"���?����?���?ͧ��X̦!c�kTꟀ�E+CE��Qሌ�[�t  �����T��4��'���?��?!��=rJ�pJT�m�����Ԓ\9��ݴ��DܒrK`D��O��I9�u'��� �õ(\Z%�t�a垰`( +�3O��d�O���O��D�O��?aX0k�S.��`�k� 3z8a�FIGy��' �6�MuK�I�OEn�A�N1JE8�.۱n+�S,�j�x4'��	���S
;d	nZ[~r�S�R�q�7�ױa=j��Wh��WR ��ov?�+O��lZ~yR�'���'��(W��R�bE4s�lƍZ�XJ"�'4�#�MӒnX�?����?�.� ��7㓵L��Hq��Y\	��:���`{�O��n��M�T�xJ?I��4_z>Uk�8�<�@j��4,����@[�#G�d���.�c� $�^wG2ӧ56+�V��@ÅK�,��ak����w�"�'�r�'����Z��k�4B�B��Z��H��E4@5�M�!�?��5u�&��Z}B/z�pb�h��!�����&ӀW����4�@pߴ��dN�	�������Ӱ^N>H�ł� =��*�E`0�ݴ���O|���O��D�O�D�|���#t��I����Q�h����	)���	�:k�'�R���'H7=�"hQ� ��0ч�_`�t"�Ɵn6��S�N�P�m��<Q]D��j��<'��1@��x���άnO<�[���<���Q����pq����[���H/��j�D��������	ly2�lӎ��Q��<9���v�
c��/)z9� �$U��9���>	q�iXP6��B��0z����h�/I~�k��E&p���$^2���eE
h�VA�'E��]*..
��l��N�z�|�+� ��Ctd�y���ߟ��	��p�	ӟ4E���'��1rPJ�
Q��9��)�Jk,4	��'�6톌1:�D�OL�o�}�Ӽ{���$U�汉��ǭ3Y�Us&�R?���M+��i��U+P�i��-��i��O_$���D6^�Йg�Ǘd��Ǣ�y�G~Ӵ��|���?���?��b�>|�@�M$j�j�0!�M3{����.O=o��[����	��l�	v�S��`�o�0J���1.G�(�¤�E-D�����Ϧ�ڴu����O���X��3��L��#f�P����
Z�8��O:�!+�'�?!�Ϸ<���i��"w:�!H%�Q`����}����͟��	����i>��'��7M�:t��Ĕ�]{��$�0K]�m����&�N��]ͦ��?قR���4 �V�p� ���Km��(5e��t$�Z�	�,6�"6-+?1h�&J7z�	:��.p����^{�)�r$"lO��W�C-u���⟬�I�X�	ҟ���d��4p�	x!��
z�Yi�"
���Z��?���c��K	>����'��6�'���$�u�I�;"P���w��=3pD&��������r�X=mZs~�@�\��u��B.�-��,�8#*�"i����R��P�4��4�����O`��Z�F|�#�n�/:x���A���D�O�ʓ/}���#��'��P>U�䚸���K�q9v̻24?�^���Iş��I<�O2qI���D�������H�B��$:*�QMѹ�����[A��O�5a+O��]�1��y"���$B��[��aT���O����O���<�մi,�����A��j]>Ўa�F��a�r�'x�7�:�I3����O��+�X	,R��3��\�B�{�O���?EF6m$?	VB�^���I6�!�8`���ˌ}�X
��ݴ�y2P�p��	 ��T3�g�$�!���rbN(aڴ2j���*O(�D"�S�M�;�N��G��=;�����E3Z����?�K>�|򐋊��M�'�pxv�>�yyU�Y�">4�1�'������V?�K>1(O����O��"Acʹ@��a4��q:���O����OL���<���'����?���2=���D�'Z�)��"G�;3�H��"̥>����?�M>�-@��b����@�t��x�SK�f~发:�R�c��i*���B�'\�ᅈ��@ʳ)b�U��~"�'�r�'���Ɵ|�6CH�Bmpe��S��������P�ڴcL�����?Q�i��O��P�*�X��f��l����C�ן,���O���O�`cҮz���~�l�H姫?ū2)�	���7I�}�hi���n�ly��'^��'���'�R�@R�����������ǿ��ɯ�?���R���I柠'?�	�j�z�9҄K�}�Bh���)4�B�O"�D�OJ�O1�-`���>b�CGD�o\�q�g؊Z��6mP~y�j�?�T������D8qL��u�;T�sIʦs.�D�O.�d�O��4�Tʓ��&�9�R+�K1ll�P"�8��m�F��1��he�D�谩O��o�M�5�i���� #�;d��9�×f�*mrE��*��V�������v8�D����v���_:���phޓd�p�9O���D���2@Y�)%S�m"·�G�~˓�?Qu�i��<`͟$nh��vY�B��5ĔP�v/G�u�L5%�P�Iɟ�S�p8�n�u~�]o��C�bS�[jn�*afҶC�`��J�~?I>y-OD�$�O���O���"�?+�W��L=P�E�OV��<�7�i��%��'���'��S�~�0=AC�#`�lQ勡|���G[��џ���B�)��&��t��������*���|n�(@��+A^4���ASП�h|�#�S�P\���M�����C��'���'.���R��i۴D������/.�ш�K�<ጽ��Ō?�?�������So}�'�q�-�6NZ�͑�l	�G�6����'��,�%�&��`K���xv���~� ��bυy�D��g�DV|\ �?OVʓ�?9��?q���?����J\8`�`��r���w)ɗ"Ⱦ�m/N�'E����'��6=��h��:Vb����,~F����O��D8��i��u�v3OL�B7�xx�$��d�{�:O�q�c���?�a`6��<�'�?YB�M:m�H���֐((����?���?�����D��)�BHǟt�IٟԱ��#�B̂s@ق!�b +�A�\��:8�	�����C�e��I�=;*��É�?���={�T 6�܉��|�&O�O���Xe�%���FE��b@:;����?q��?I��h�`���}���x6h e�lA4dаz�����ߦ�A���UyGj�H��=jD�
�M�<. Ig$E�LK���ȟ�m���Mˡk�!�M��O��떂�&�r�.�nYHqN�"yx@�3�z�Or��|����?���?���&0r�_�b�Lq��W�Fu�P2/O.�n��V(X=�	��(��q�S����S�
H[��(�B�7MX�l�$����O��-���@� 92�C'���[�$�0k�Zt� j
�&��a���`�'Gx$��'�j!�ъ��FC���̠O���c�'��'y���TX��`�4^|�Y���h���BF��j�cٚ5PȒ�)4���|�O�R��?Y���?�ƦRW@+��^6_&�M�E��N�X۴��dX-j��I�O��O���ղB�<���ٿf��hr�H��y��'r�'���'���i�bV�Ѻr=�d������k�Z����&�M;��|��DR�֙|2�I�Dl<�Ai���P!YĦ��G��O�n3�Mϧ  ��H�4���ғW9" j�=T��{��Rp���EA��~|�P�4��۟���ɟ4��JԙV�H��_yڲ,z�D֟$�	@y�ml�H�s6��O
���O˧E�(#��5&Ȉ��4��tx�x�'��˓�?��43#ɧ�i���Z]��Q<D�,W"5f��Xk�)ń�7-�Iy�O2$$����_ܴ�*f�E%%T�1k��;i�B՛���?9��?1�S�'���A��)��~���R��K!�܅�@
� �P�I���4��'�T� @��b�!mv	Yf�ʵ�~M��P<�7M�pį����'tAZ���t�(O,���`��3���A\�p���9�?O�˓�?��?����?�����\* -���G��ۓ)�{�*�m��e�'R�'��O�L`��nG28I��QD-���@K���b�v���O��O1���Q��w���	���E���8BΑsAb��l����$?	p��s�'.f$������'�u��/Q'ps�z��U�r�'�B�'�2T��*�4b�R8.O���(8�h�[�b�0H���"=,���K�Oh�d�O@�O8�����aV~����,7�&MC域�(T�y�ɛ&j,�S�y�jLǟ��b�!M�%*���-��!�GƟ���䟸���lD�d�'��XX�`��*<`�!Ȑ	�����?�r�it��+2�'b$mӺ��8U:82 �*Q��Ԑ�H%��'.�'�"�����8*5�äR���@�cv���ʴ[P<�G��r���%�����d�'�R�'W��'���3p/AEz�ԑ�D˽ h0$�Z��h�4f�� P��?������?�ՠ̓d�XA�LԼ2!R��!�I����t�)��l�@����,[�ٸaO�=-O�$0�-ͼ*�2�zZ>D�p�ORe�M>�(O�X��U�:UQã0H�1v�O����OV�$�O�<�3�iiVM���'�����%�쐀j����4P�'T�7m:�I8���O ���OX���=xtf�� S	7r�t��I�6-=?�UD����I?����� �L�X'0!A��� P��a�Hg����ٟ|��՟��IğP�"6��#⤘@�/��B�NdY����?)��?��i�@z�OD�K|Ӯ�OZ<��	J�~P�V�Z�Oٚ�C�"%���O��4�R	H�Jk�P��fd��b�Q,Z�V��!(`%�F�ѿ-L�䔏�?�*O��|����?y��{�Ȅ�!�#@���#�1s�a����?�*Oh9m�X9@��ԟp��y�t×*,�B%��A��_|���O� �'cr�'
ɧ�Ib��x��S4��	agi'kG��QGaÿP�7M.?�'��	y�	�3<~Y�`MO�4}� �Whݞ�D\�Iӟ��	ğ��)��Cy�de�(�SƏ��V�4
�	!;x,}���^���y����a}�JiӤ8;�H w<�A(�(G�h�� F�19شZ^}�ݴ��$Ɂmw40��'���2�Z�#׺v:��b��=.���}y��'��'��'�rT>Őw��<h2 @���8�~9��C��M{D�H��?I���?�I~Γ=h��w�޼J`�V�~�"�k�ĉJ�C��m���nZ���S�'j���۴�y��J�K�l�HϵGX��:�	�/�y�� n��@�ɮC��'��i>�I[�VD�l3�ȈJ�!S�W�����֟��I����'�7�0We���Ol��S��P����T.�Q�]�Dl.�l�O�oڽ�M�Ėx�두�E�5�|>������Ą�<?��X��ܱ.-1���`��+-p�dI��ԡ�'ϋ89R���C.���D�O����Od��,ڧ�?9�H��hP\�r�	�:p��A�?Yıi��+�R�Ȳܴ���y��y�(ً@�Ӊv��!j��c�͓��F�s��!oښ(WR�m�[~�لv�>���� ^�Avo�X����ؓ�~��5���<�'�?a���?���?Q�샬M������M�@��i�7a�)��Dܦ5ChC����	��'?�Ɇ
�Ve����2�μa�Eܺ�<�B�O(�m��Mבx���뉰S��m���ۆe�v��",ٔiϮ%;�
^����X2dӠQs��M+��O��U�~tꅉ̐Hڲ�9��R�Z�Ą��I��M+ C��?�E�BJ;�a/ִa�$1S����<ia�i��O0��'C��'��-5�,���dۖ�irc	��K��i����%Xl�$۟���������(��
H!q P}{` /xL��O����O.�$�O��-��
A�<����l����3}�X��	؟ �� �M�ccGK��b�b�`��#]�%������	�|A2 ,���O��4�L�[��qӪ�1��`�i_�"��� ��IlP�Vj�?���IK�	~y��'��'�ŀ�W������V�R��8��'��	��M��̛+�?����?�)�q��UQv�K$�@�+���Y���8��O��D�O\�O��'ZcA��(��m6A2$�}>�y�5�-׊en���4�ll��'�'��U@�`�.a�8��s}��I��'Jr�'���O��	;�M� �^ ]@�(��Ͱ$W�yk�%�*�"���?1��i%�'��>���i���T��;i�uЕ�E�Pb��p�lӬ�mZi�xemO~2�Lp�e�'��6��r
R�t�H��h�%��<)��?Q���?���?�)��!b����|���KB3��X�A���9W�ϟP�Iܟ�'?U�	��M�;R!�̻���_ђ2�͢d�� ���?�M>�|R�+�7�M��'�"��P*ޡnlA`&ʅI�b:�'����[BA�v�^y�O�o؞B@�ᅋ�lY�+�ϡ��'���'����M���?!��?ѡ�� \�a�����������'B���?a����x���c���������Tu�'>̵���=<؛7��E��~�'��ċ�F1�Ǖ*8Y��P�'bR�'[r�'��>��ɈY(�)6��*Wӊ�BAE��q�:��I��M۵��?Y�K��v�4�f��VG�/NX��q�_�B�5(�1OD���O���D�/r�7=?ї�b �I[]E�F@�*� \z���s�ր�I>Q,O��O����O����OZ<��E��i9��sF��<t~�j�G�<� �iDn$���'b�'B�O����u�0	�WG�1E�j�*��06�듊?����S�'FĘ��[���A]y�DD�aŏ/3}���'�ɉR��ޟ`u�|R��:�$�?�di�����|���#I៰�	ܟl�IƟ�ay��k��`X�d�O>a�	�9h��Ì�Y`�4O\�lQ��4����M;s�i�6m�%]þ��Æ��Kd�A`Z|(���Aie���jmƠPU�����>��(%]v@�Ί%n�P��H����I�����T�����	`�'O���Lۢ ������3hr���?Q��9w��9������%�@�v��`f����)3��V�	ȟ(�i>)���GЦ��'Q�e�&��Y6��tH�B|dP��N#eI����?!�\�<i*O�I�0���O��;����5	��9!HZ7jeJa@�,dF��<�G�i3�@�t�'���'����w�d����D�P����1v����'��h�>���i�`7m�\�i>m�S�$'�-��ĉg̎����J
v���H�+[07�DyfL+?��'om������&z�,�pjB�yI�� ͕wr�MR��?����?i�S�'��ăͦE���>Fd5
7KH�Y82 (�C*����៌qݴ���|*6[���I>Hɪ�S�"�Q�^dæ�����	��pƌ�Ŧ��'���	scx�.O�Љ �i���K'��l�'0O*ʓ��=���N�c���aY--���Fa�4�����RY��'����N¦��[q$�Z5���@m�Q�&[��4m����#��)��"�X6�j�lH� $v��ji�Q���{�x�TR@
�-f���7�D�<���?cWLt=ů��;Cl���ɐ��?����?���$��uɁ��؟|��ʟ��DLB&%��I�MN$����t-H�h��I���I@�ɓ1���jOC]넨*a�Fl��=�v	ـ�E�
t�|j�J�Ots����:�
ǠP��H8�/֐_�"�����?���?���h�n�d.Cb�pt�M�:�~	���(<$�����!������M���w}�ʧF��Q���&*��(�'*v7m�����48��\8�4���\,�q�O�Zx+a ��!]�a�0%�0��ќ|U�0�	ɟ(��ܟ�����Ļ�L6jG^H�D"/=�&�9'�xy�z���&i�O���O6�����C��"�ש~ )p�ٯl�V��'=L7��¦9�M<�|�աW�K�b�9�M�;�J�2�UJ&�c�4{��	�Y~"Xr�OL�O�A�����ӆ���$�̦����?����?i��|�,O�lZ{7���7@ƽ�'�0'����nA�64�y���M#�bj�>9�i�6�[�M2��W�ju�g��iH��5H݀u���mJ~�Vu�������ȿSF�)'S�a�"���U@T�<���?9���?A��?A��䥞�}�
�!�A �D�K���NZ2�'��}�n1�9����ǦA%�<��@�9.N\��KC���� �ē�V#t���[47�0?Q�ϛ\�? fa��"��x��������фU6�~R�|�Z����ȟ �I���ע~4j`�桊g	V��w�S����	wyb�v�b�y�+�<q����静c��-���A�4I�ݘ*�Y{���OP��'q��'�ɧ�I�~�,z7"��{ʐa��ˑ�V�ց9��X�{ 6�
`y�Oш�����x� 1�d�1���BG��1�l����?Q��?9�S�'��d�����4>�M#Qc��0j���℃���Q�����۴���?9V��lځ'�lRw�a��ŹuJ+��@8дi��7Z�}s�6�<?鴮H_`���GyҍI�id܅���:�>YCS���ybV���	�Q�(��J��~$���B�:T r	{�4����?����O_j7=�V�5Bټhz�Y����UE�X�j�ۦ���4h���O$|�p�i=�d��[j<bi݃	􁹴�͊?���#?��9�'$�'��IɟL�;'�$5-�=6Dt�!���3����IП��I՟�'�7-T�C#����OL���pa�uc%gS�54r]ࡩ��Pc�� y�O^�d�Oz�OR:U���z��a�7�C�	�Xx���� �2j�8�2����6��8�r�ʟ4���L�^aj�#_���|QG֢r ���I�l��ٟ �)�Sܟ��I�\>���Q�{��P��&�pK���I�M˴�X��?1���F�|��y7��(C'���� Ś`Hys���yr�'pr�'�`���i��O�����t`�Ӭ ��T�h��bɃ&\�'�i>��	����I⟈�ɰAvH�����ѱ~���)��wy�$f���X0�<Q����'�?a��G������J\e)DC�L������a�)�\}ذh�,��T���D�G�~�Pg��Q�)O�<r����~��|"Y�0[�M`&d��FƵ8q�R�'�2�'��O�I��M�ʅ��?���?f���7E��%��������?1��i��O��'��'s��F(*��:��.K�F�A` /o)B	a��i���! ��y�QڟL���.����qf��?\��u��E�����O��O&�D�O���$�S�6��p�G��s��9�����\���ן<�I��M3B"�K�4oӸ�O�ܸR d���ό1-�SF��M�	�MkG����ٷ��v���Q���&t�y��Ɲ*�1��e�)n��c�O.�O���?���?��h�J�B�._)sC&���G�k������?�.O�oڪ	�Z��	�����u����C����椚�upb�@:��dr}��'X|ʟ�,�w��/��Y��H�uE^�R�ϲS7	��i��>�i>m0�'w(�%� �!Q;� r"�
X�06f*�HrٴX�L�ʡH��%�Dˤ�&3�`�P��(���ݦ��?��V���	�*�ȭs����n�8	�"��ܢ	�O����:��7-(?A�dE�zq�O:�I 4B5b�f�@Q<����	\���cy2�'������Wh0+�� Ś�B	w��|��c�O����O��?������s�E��v�06��ZD��k��}F��*sӊI'�b>�����v��!0�,����ʻ���	��ɂ�OL�O�ʓ�?�'�ʨ��FĤ�E�]Uv|����?a��?�,Ov�n�?Ѝ�I�`�I�ۢ���"��d��qK��F	E���?��P����ȟP'�xrH_0A����Y8B���M>?A�ĳQ%[۴��O�.���?��+��m#�i��f2(���#��?)��?���?����O�m��N��������N����O�qlZ�@ر��ɟH1�4���y�L;Y`�i�+tt֌��m�,�y�'���'��=`#�i/�I�5dYS۟@�CeA��R��	(ؓ:��,p#4�D�<ͧ�?����?����?y��V e!�@ �&���#��W���DNɦ�4E��P�I�$?U�I�Vui���֦���ão[5S0P��O��d�O��O1��d�떺0��3�ƨ&v��@�lF�x6�"?��H2O9�I[�	gyR�O�e
�iCDY�4NJ����0>ᐶi5R@��'l��H�� #T���j_�T��Ԣ��'v:7$��0��������47͛fd׀J�Q#ц^�-����$���hi�ɒ��i���E�}�uПJ����.��zꈚ��P�K= Ub�*����.�O&,8�S;�}Аe�~ �y��O��D�O��l�'KB�'+��|���<�(�b�	O�x�39�O5mژ�Mϧ,��ܴ���M4;��F"��3�Iİy�I����~�|Q��?)��F7N~��aN�By�i�c�G�'��6��[�2˓�?�.���y��@�:!�U��o@g~e���DA�O~���O�O�S8wiUs�%0r��P
F�A� ��s��'v�L�m�;��4��c�'��'q8�S�CӝcW���i��{�lh;��')��'�B���O����M��" �
�s͚T7!;y���0��?��i��O�5�'��j�h4��@��+wx�o������'0r��s��&���p� $2��4�~"Ш��:�>��%�AI �a��<�+O��O&�D�O��$�Oj�'o&J�!��ƬkD�t�f��:Rj8c��iL~��U�'���'��=mz���%���?��EA��W
\��3Ү֟(�IU�)�,e��m�<� �R��1T���q�(\"
,<! ?O��7��?���3���<ͧ�?YG���[�RQ�e)J!��K� D"�?a���?y������£M������\��)->�>�@�"
ǮE�w�Me�2��	͟��	_�	�d�xHR��{̂ӲJ�"'��.�8��I/aDZ`�|�-�ON`I�y���1���{����/9	hP���?���?���h��.�x�6�5����ؙ!d�+���$�ަ�z��Cӟ����MKJ>��Ӽ�d��Hh�L�@��(d���@Ə��<���i0j6m��᫤^֦��'����j
"��]Vx��#���4{�#�#����$�O��OJ���O|�� 2�ʌ�6�9W��P��U��qX�B�4-���z���?I����'�?av хdJ�d�p��g��؄�[�<����8��g�)�6��p0�'T�n((Y�AE[Ƹ���#svx�������O��H>�-O����V�k:�a+a �gE�ه�'Rx7mU�Oi����,#���z��-[� !�� �r������?2[��J޴`-�fNv�u�7IĆYf�Ke.�$_�
4R&�f��7m??��N\��SC����R�d�>3J��aL���裓m���I�-`�S��K�C�^��r�ͪ"��Д']�c�6$ʓ�?���4��N۰U��&G2��R�հk��!�L>Q���?ͧ]��ߴ����6L�v岆�8TI�7� 3�mkrB.�~2�|�Z����ӟ�����<���N�R\�\2pT�T�.-p��˟ �	ly�E`�,}�PG�On�$�O�'[��A7C��T<��r�&GA�8�'���?����S��ƈX�@�@/�$w2����IĤql�����3�`��O�i���?�4g&�$Ɯr�B� '��}�,��g���$�O.��O���<�i��$ȃ]$j����Ͷ96~�Xr�'<Z�'��6�'������O��,�+E�P�٧Gq<I���Oj����6�=?���@�5����0�����a��j�+�*Р�S���y\�D��	�K�4�0g	�?��Q����w�����4D*,$+O�D<�S-�Mϻi�ȼ��k��0�T���M�{U�1����?K>�|
��D�M��'���Ҥ	�[/�}�F˃� �Q)�'�����#�F?IK>�)O�ʓ1��m�I�xhR�UAS�B������M��Y��?!��?yQ��u_.4ۧL�$k����1��'���%^��eyӪ&� Qg��pjPx!c�� g6kG�&?���"5�شT �Oq0����?Y� :� �c��^ �a��e�<��^��-0�)]�!���ϭ�?i�i�L5"�'��p����]Za�
Ќ�X��bg	&�D�	��M���i��6�Q-�7&?QU�ԒM�2e� �x����o���{���J&���'���'��'��'I��5���Y2:Tx.�{ǒ��CP���ڴ���+��?y���䧁?�#j��;��Y�NȗH�>L� d�g���ʟ��	G�)�� а�c�CV*E�a���Vfh��Fv7^��p��1��Oz��I>�)O����mA58��ʆ���be�l�F��O
���Ot���O�ɦ<A�i5D�*��'E��Î�cg
���N��.s"����'׺7M,���O�q�'�7mĦyߴ'�L%�E�ޞ�t%�2� X8<�
��%�M3�'��\V������d�� GDصq�(��	�`(��X�|��O��d�O��d�O��D8��g�]p���Sꊽ�F'&�q��ş��ɯ�M���Nw��Ew�z�Ol!ȁC��ؚ�,#(���P˗B�I,�M;S���TD`�f���B�LB�$�ӱ��?XA��Qc�B�>�,194�'L�'� �����'1��'b,5��O��m����66 �d�'��Y����4k3t}Z���?����i�w ���޾K-� SWܪ;i��'����M�P�inO���hs� �1��6`�^- ��w�����n�&��fO&?ͧO������DYVua� �+[L�v�A�WZ�(Q��?����?��Ş��D[Ŧ�*��<;�D�����KlE2��E
0�����Οt:�4��'(4�$b�V�U��H��U?�N=�@�[�_U~6���0���ܦ%�'먅J#���?���]�" �9�H@Ӷx�yP�{?i,O��$�O<�$�O����OP�'N��  b�9iڍ�Q�л"9�]rּi��'3��'��O2�d��nǄk��P�F<���!O� F,v@�����K>%?Ð��������e@tϋ�x�8۶�W ]�(�̓F���b���On�M>A/O�)�O:��!����!T��d{��2�O~���O�d�<i��i��#V�'���'#D<°FX�)0l�%�64<�ؕ�$�@}�lx�lel��ēq~�A��j�f
}Zd��q��%�'�T�����$R�գ��d�K��� �'f���֊i!�QIG�̖�r$���'���'���'A�>��I�,����x��]�alP� lD��I5�M�R��6��ʦE�?ͻ]�~�Xgl�1Y��pۀ�	c�Dp̓Ǜ&�r�&ho�-0Ndl�m~bA54�\��S�H����
@)!J��PW E�z֦����|P��柴��͟���ߟ8{�ɇt�բ�?9���V!Hzyb~�lY��<����OQ�"B��l}d�[�➒�@q{Dn�>�4�i��7-�h�)�ӻ(�� �͑G��S�"�y�h�kĝ�E��|����M*�#��'���$��'�Dݛ�I���Xd��B5d��	s�'�r�'"����Z���4S��B�Z���2X�`�xA�B8%
zD)��zc�6��_}��n��!lZ��M�IC�]�n1q�AQ�r-��-�v���4��d6�M�����O�7'E
X��� -0)M �p���yB�'���'fB�'�b�ɓ�\w�XY�%]r@�M%�JlZ8�$�O��������d+�·i��'gL�0s-�
2�@l 7�@ �1�|B�'�O��8 �i��Io���p�ͯQ���F	{���0�G�r"�Ai�	jy�O��'��Ä�r8����Be��f`��%/R�'��	��M{$n����Oʧ2Mx9����:"C���$F8'iu�'���?)���S��%F���}{ъN�S���-I����� ^� Y@g�N~�O���I"��'��,�5Û�u@d-!��k�	���'+��'D��O[�I5�M;6E2[o�y���P�h�����(T��n%����?A��i��O��'WR���_�)b�!�����=
uR�'�@;�i��ɽ��c�OL�B��}0��ڒt�^���\0/�uΓ��D�OB���OH�d�O�D�|�"%���U�DE�x�pj��("xl�7⒤��֟���T��h-��w�ܰ7Ë--�̹&��:Z�h����'S�|��D�^G�&>O.��V�[�J�S��	 �p8�7On�����~��|�Z��蟼z���_�$�k5�W$mb�#d��0�	����	yy�E~Ӑ]:�K�O����O:��3	A;&7���֪��$Dt��3�ɣ����݁�4?[�'	LmK2%���&�kѩ$�P���O�M��B��A�6�LP�ӥk���O�*e(��dB�My�@�"�P�5%�O��d�OF���O*�}z�EU�qGI؍��-�1�/a�@		��]؛���%12�'?�6�7�i�aB@▾@W�l�a�ҧST����e�hܴ}5�v�tӨ(�Df�T�I��5�%���\��w�Y���8�ΘN(`[����4�r���O���O����2g��mpw�^#_�%��Ai��S���ј(�	�������1@����I���	����*56������IL�)擨�LECb*J)?���J#-i�\�JƦ1k/OiI!$��~B�|2X�h���@;��̫��	�w-2�Ů����	��������SLy�ct�La
u��O�ɡ���0��� �
� �F��$�O�ls�z���m���M;է�%O�9�E%�=^��p�`�z�l)�ٴ��$�%.|�I�O��O���a��y�H�y���5�͙�y�'�B�'���'=r������p��$l�n���I������O����ئ�ғ�>��I��M+O>!�)4/�����ƲB+֑뗂��3��'ET6�ʦ�S*'RUm�U~&�(h ���v.�!_��PV��lfR58ǣ�~?YL>�)O���O��d�OPT�o�o6 �4bʶ���Q��O���<a��i�����'2��'��SX:>��e��~�����6�(�q�����]�)����,����Q�%L����
\l�G�&|\
�������<"$�|bl(
�8����>4�>�HdmA�;�"�'I"�'����Y�P��4#S��#raaK��xDXe�c��ĵ���?A��i��O��'N��IF��1�cʌ(3|�SÚ;��'��%2ùi��	�z��:s�O��',����F8%��W%m���f�-za���qAjѰG��]N�:cD,�Mq�&q ���d�C�ڳJ��{~��L:(��TY���7�,xX'��E������J�/��2H��oV�;u��1���!@	99��e:4�F(9��7��6 M3j٠I�@��P���p�P٣�י+���z��C"@Xk���8 %P�Y�h�*+���peX�!�0�p�<eAn�с&¾C����#�q3�f\J��g]�5�D�Q��2yy � $�4k%�SgZY T�� E�\*�X�%�8t�m�쟠�	ş�����'��C ȉ����b��>m���`�a�
��p�)�'�?��$��J@cR���Cw*dB"��I���'MB�'0`�k��>���O`�d��|ٔ-�,�^���ک>�n��֍>�	)Q��c������	�P> �0-N�]�D��A�f���4�?���ܢ/��'	B�'ɧ5�.�/YM6�P�.�;����r
[���dU�}�1O2���O����<1�A;nP�0�G�Xq���0d�)  ���זxR�'�B�|BQ��C�˄�9j��z����C� C#t �b�������kyRA��e���VN�Q
s&�����$���r��등?������$����	1+P��C@M4c�^�3G̵D�듌?����?)*O�t�u�K�
T����h�( @XY�!��%�f��ٴ�?L>)-OL�k����j���4-R�[!�	�1_0�&�'�b[�@;�'A���'�?��z�T�i�0P�๘&@������i��ty�(�2�����s�6�YS&@�C�n��@q�pb'�ij�ɁL�p�۴}r����������N�X�*A�d��M>%�fF�qj�[�0�T"4�S�'B[�Q'�
� ���$S�sQ��o�	��!��4�?����?�' ��'�"�L�����Q ���q��n��7�Qj�"|��U�H��P�\&�Z�Hu!ӱ>�����i��'�R�*^u�c���IU?�+_=h?i�`�H(d�]9���i�z쒱�<)��?9�|�� 5��8�������tTB��i�"�6?vO,�D�O>�Ok,�+�&mxף��w'3S��(_m���d�c���I����Yy����4�����(< ����Ѡ�ΜB�=�$�Ov�'��<��\�5*�PE�r�|��R*BbF��<9���?������
�؄�'�v	;��դ/�|E�pC��
|��m�oy��'��'���'��	ɩO5�0Ʌ�cOHd�sn	4TW�8J�U����ٟ �	ryrK ),���'�?�0�O�,��Q��N� �����i�?���'��'��'q4��`�$e{z˦$	�Y8�`�Z�[���'�"[�� �����O����ם�={|��`�40�ҹy�%C$p@J<y���?�e���'�I�A�*��a���KY�9 ��U?mG�&X�\������M���?������R��X>C'.=)V�[7��J6�;Ă6��OH��'ь㟤�}�S��f��x RcJ51p�q��㦱��DҨ�M���?���Z�Q��']8�b�O�#xB�e:��pAU�o�K7,	�|R���O����gB�83��6!;L=�S��ڦ�I۟(��!�h��'h��'���Ozq�t��>��E�6"
�&�e�d@$uD�O��d�Ov��ә9��{4/4I��JĈۚ,Ƣ�l�П��$������<�������V�X\���`��al����\H}�b��
�\��Iğ`��ryB�ΖT��T�J�9$�{#l���lC�a�>�(O��'�d�O��ȯ9پ@���s�l���!CD����O���?���?�.O\$3@A�|�`�)�`H�Qf��0�~-9���Օ'B|�'C� �V�r��"AL|�@�,U��Ô�Ƚ`���?!��?�.Or����w��'M|}(� �%T�f�j`Ʒ"9V���
q���:���O�dO��'��=v�5����#<� &EC�F���mZ�����Gy���;��6��k�5�*�酡�4�)A2)7~o�'h������IZ�s�֝�$�:hB	��< 
ҟ~�7�<qvb� �����~����x�����vP�H�I��Q����cq�4ʓ�?���v��O���MKBi�� �@ԋP�=��H�/�æő�`T �M3���?���JS�x�O�A��fa�,�ш֛wn�r�d�(10��O@��<L~��?�D���	� X �cݫw�z���^��V�'A��'^�"�.#�4�<����X{��Y�*�>P��2�&�4�`�F�$�<�#��v�s���ϟ��#g��!�d֯rLP�ˁuZ\��ߴ�?��i�	uI���d�'�bP��!v[;w`��;DB>n7jy
�$���Mc�c�<������4�$�d�<���~��m�ROƿZk��Kb�δ9\�j�L����d�O���-��ڟ���+lx��6�ĔF��003nLrn�]�_�<�c����uy��'!L��f]?��6ޠ0���mC�Ta�i���Y��?1�?��̙dX��ar���QT���o	�ۜ)���>���?����S([�( %>�B�C)u�x�bRE�9!�$-�v�ӎ�M+������A..���$���]�8k.��.��fq��g��M�����O@���|����?����#�ђ�R|P�E�;"�%k�l�A�����	*j"š��!�~2�(�2D��KF�;p�&�zd	�{}�'�\�*%�'l��'P��O#�i�	 cҮ����E)������pӮ�d�O�q�Q���\1O��8�aiT�\�H"�8���иi.�����'}��'��O��)�a�;�4�#M�#a�b��F��3&�K�"n�ZԊ�y����O�D�A��	�дRg]�M� ��Վ�ɦM�Iڟ��	#��1!I<ͧ�?q�I' Q�q�E�8i�)����7?����i�'�2��"��<���?��ڜ�B*�R���� al&ɀ�i&��X��O��Oj�d�<��N��C?�`�@�A�8h:9bG�iu2�K1>|r�'{�U�����ֳ��a�޿RR�E!�(�&e"n�N�	ԟl�	I�ITy�c�
��!��˟=*� F'X-V��'�ݟ8����'�z�ku`j>}bK��3v4 %cR'b�D�q��>���?�N>�(O�@1���O6	 �	E7tp�҇J�bF�H� H}��'sR�'�	J��M|R�mJ�[K�qM�*��#��W�v�'!�'��I.,��Iz���~��(�5��� �DAk l�%A�6�'��	ßH�5#���'
"��5�g�4��M�ŉ\��8�+ ���?)�p%N!`i�A�S�thI#�����A��<HI�,�3�M�*OX"��ڦ���P�����'���R��<k@�M""a�9W����4���ȸ#��$HW�d�s�t\��FM�qЋ�0�0t3$�]��M�'�ӛ��'�r�'z��:�4�t���L�4�fuر��xS�k�ɦ�*B�T���ICy����'�CN��GNZx��S�h���,6�O��d�O
|�E�GE�i>�	ϟ�B����c%�T�b �'Z3�y��AF��Mk��?��)�v�u]?�韰�	蟜9��}i���V(��K��d���M��+7���EY���'7�Z���i�y����Br�e���=e��K'��>�S��v��?i��?!+O��%.��xl�hΜ�2����Ñv�"��'{�ߟ�'z��'���V�N��!C�9ArЊ��ѸG3���'����	��З'hܭr�my>� ���Q���(`5#��]���i(�I󟠖')b�'�r)@��y��5�$����D�3���Q#م.ڐ��?����?�.O��3����?�'҇J��x��f�Mψe�TLװu�F�'K��䟨�I���h��l�X�	z?��CD'[b�ĚDƋ�/�<ɪ�������ȟ|�'�:4��̳~����?1�'�*�@`.гm�aKd):��q�U�h�	���I*�$"<i�O����b���3I�Dx<��4��dܧIL(nZ֟��I�l�������FT���Z�}b����W�`0Cr�i7��'�Լa�'LRS���}z��?}������g5��2'�SȦ�� J���M���?�����[��'��U���E�BE>��A��:z&�� �b�����>O��D�O���9�S�`{���$�6�Un],n?,�3�'�MK���?���B�r�1�P��'�R�Ob�P$����LR�q�E�%�M���?	�%z&T�S���'TR�'�0�����b	r��9o(����b�p�D�lo
-�'a��ΟX�'`Zc����QɒV}0���r �*�O�{W?O���?����?�*OrY��ſs�I�l�5;�
@�P�|���'{�I���'zB�'��K�0�vx�TfY�!�T$����������'m�ٟ���矰�'��Dh>u���,B<��b!$:tU3��qӮ��?I)O��d�O��D��D]��iq�R�b
��pM�*���T�i,��'��'��&v��𣮟:���v�H3����q��eZ�Y�0U�2�i"R���Iן$�I=}J��	l��Ț �Dt�$��XBLP��;%)���'�"P��R�AM:��I�O �d�"<���LI�J�.D�9���A�"JG}��' ��'���Kȟ��Tj�.�9��݈7`
,pt��9'���!�'����!m�T��O��D�ʩէugCĢ6��quf7TE�	X�.�<�MS���?ٕ��<��X?��w�'qlM�0C8?�*�k�bO�$�*nxQd$ߴ�?���?a��8���^y�h�!x���4-�a�h �׼��6��$w��D�O��d�O��?��ɑ<��01��*H,7��d�ٴ�?a���?I�h՚P0�	qy��'��$V�&e(P�N"7N�+U�
��VT����89,��)���?)�&�=�TC]�>�� FКL8tP�i�B�וt������O���?��A%��o��e���r3K� f�@��'�:P��'��I쟰����ؗ'PT�"�Ȫehj���L�/e����Ć�"Ǝ����O�˓�?1��?y�R�sZ��2���3��13�[6�����?)���?���?�*O|	*���|��ɟ�+�%� @.L�V��ߦٗ'NBP���I�<�ɵ]۪�'Jƍ��Rq�݁����'��'�"P�8��k���I�Očs�(��t:i�A-ص	:$�������cy��']��'��j�'�sӦ�CB�3m��jVԸ����M3��?)O�XI`H�I���'�2�OjHl�)�S���Z�d�"���#�@�>���?��<��̓���O�;x萨�F���49XɈ��3	�6-�<���v���'�R�'`�T�>��ξ!��GWEP:�M���o�����I�9�����D!��_��dIK'KI���C-#~�7m\(.�bdm�ߟ���ߟl�S2����<�!��5)�
P²�N/VՒ�!��M8a�
��yB�'���'Q�����;tP�`�*�(��
�P��l���	�� �����$�<I���~2 s��!ˍ YyJ��	��M�����A&"�?��	П��'r�����!b�"�1����r��aoZߟX9�W���d�<����D�Ok��a�l�p�I2{X��8P��V���.���I�����������'���؏L�4�P�M��tp���ӌ��O���O$�O��$�O e"Ą�'ߔ	a ��7@!��g�	.|��<)���?�����89|��'Of�{�-�&�U�h ��'�"�'��'�2�'��Z�'2�y(��A3$�J@rM��a�T0ӣn�>	��?�����S#OB~�%>9{@�P�l�8%�ĉ7�K���+�M����?	�F�$�0����ɀD�֡y$���xjGJ&h�7�O&�d�<��	�&�O�2�O��	Xt��nT,�"� WX�t�u`.�d�O��dR#�,�d/�Ġ?%�A�H+Hb� ��E'������n�j��<A1�i
�꧇?��'h@�I)�h�;r#[�u�:dj�G�*��6m�Ol���4}b�d0��9$���`Bδom`8�c�n�f7ҫ��m�ɟ�I� �S��'�D)&��[)3#�Fx��p�fs�p���A�On�O��?��I3/ˢ�q핓61�`HA��C[~ܨݴ�?y���?�����g��O~�Ļ��Iqn�"o�}� D�XMT� ׎t�OH�(D8O�S��h�I�ս)�橡�j�	ae_>�M��9�x��d�O"�Ok,�v��H��G��o��¡�b�����D�Qy��'�R�'G�I�6���	�M�%z��BG�kB��m_"��'_��|��'^B�׭ �N�`���%y⤑jԨ��J�F�'����������'�~��d t>��ǃ	]=^=HB)M�#�i ��>����?�O>���?r�L.�?���ڧ���H&@�	O��I�m
�2����I����'�p�
��)�	=

橃Roծ_UJE��d\�Bl��m���&�����d��Hg���O0H���Y=v���dX-��hhP�i2�'��ɖ/T&��L|����B� ~�p�GU�-�h��B�L�G�m���x��'��hY;6���|2ӟ�1ٶf�9
b��9 	��F\(w�i��ITT�*�4n��ğ��S���}��td�L6.t`����7䛶�'��n��!Ar�|��IT$K�6�1�fP��"Xʂ&.��,ݕ4��6��O��$�O����Z�H�������
l�$�3����Y��Hf�i:�U	���#����d˄-n���Rf�(Ԕ��B��M����?��=%�,��D�O�I�Rp(dؠ�	�D�����i��Z�P6M.�dG�p��$�<����?����lB�,5b��р6xf0�`�ĦI�I�b����}��'fɧ56�ߟH >+¤���z`ځ(W����(h��<I��?������^�pL�����R�k��0���&I�lT�ӄ�[�	ɟ�E{b�O�,���Se>(p���H��d2�if�^����ӟ��I{y�]L��Ө^�PA���^<3e�Y!R��G�d6��<!����O����OB�(�9O^�҃O�9UP����\5*��Ɂ)	�M�I䟈��� �'p�)`���~��#�K�c5�8ઌ�H���i����Igy��'���'٪E9�'��s��+6B�*�� a׉�4c#<\:��i�R�'��1=8�� ������O���ڠw�Ή�fM&,;���v ���'�b�'ir,V�y2�'tR�'
�Ɇ�8J$��(Ɨ7&*р�'��W�+�ȭ�M{���?����z�Q��]�\���d/��.�P���*�2 ��7��O��Ă�[�5�D21��%(D�B�m\�([�/@�oܤ7-J�)��UlZߟ��I��������<A$M�4��A��Xuw������(� H��y��'��I@���?1B�  ��Ѣ���M`�ڐ�?J��u�4�?Y��R?6��Vy��'��ё7b$��C�U��@i�����'�&b���)���?q�Oi@H!2&֗e|N(�7��<a�x��ڴ�?y���	y��I}y��'��	����5b2��[��=xl	7�˟Kh��S6z<�'j��'���'"�:I-�\y��Z� (��"��"w��+���<������O���O���U �%����="��D#��J�}*�d�<����?1����JzIϧ>�pI��)���0��Cf��� �nly��'x�I� �	����F�s�̒p���)a�j��A�b4��%�M��?y��?�+O�=+�M`���'!D0{w-)d��-��hٓ���Q&�r�l��<����?��l@D@�Oq�DR	W���hA�SZ�49sM��E���'
R[��8�������O��$��|��)�-@^�,�a=[��X�Q��X}��'�r�'�(*�']�'~��߁F� �����m �����Rb��X��w�}��4�?!���?��/�i�={2	�Wx
��¢�gLL�)e�$�$�O��$=O:���y��)��4F:��&M>V� -B ��,w����ԑU)�7��O ���O`�)�t}�P�D1RG[�P�>�X4� j�b ����MS�o	\~2X������P��Rg���_!j)A�� �Q��i�r�'$�Ϟ�;rX����O��I�X���Z�4RBt��c\6M0��;m4�?�����(�I!i�� �rh� n���f��x�T�hٴ�?14�D����Myr�'�͟��xB���C�<h!	�n܎?�Z�ž���?����?q��?Y/O4�(���j��r��ޯYV��b��	���'��I���'�r�'�2`��]/T�+Sm_7nADh��~V���Ol���O����O��
،��8���4�5m��K��� ��i��Iȟ��'���' Rd?�4"�Kr
E� +׾-�}����<)U�F�'!B�'�2U� �2N�,��i�O*ɡ�Y8_�.B�?O�0�����Ԧ��	ay��'���'/���'��I�p��b��B+m�Nt V�Ʊ�V��޴�?1��?1��d�r�I��?���?	��]̠��恐�$��4�Ѝ�r!2 P0�xr�'��I�p{""<�;_~�� #^�1I~)ӓ�[�um�oy�/;3f6�_W�T�'���&?���8�b|�Ԫ6 $ �r�Q�)L�rL�?��g�	 7��S"�M<��A���47-�!aq~���O^���OR���O.�d�|B�,�	f�(r��rAڀ�_ #���.tX
#<�|2���B]��~��2 � <��+ӱi3�'Q�HS$z�<b����c?!�#O�|��@B3��#���D�����<���?��0X�4���P'+�&�ZL��1���q�i��m�[S�O"���O��OkL�t3N4J��\�/��7GQ����?J`c���I˟p�'֕fF����80H���MN�7�8`F�'���'�b�'D�'�r�O8�C���)f�}�臆b�!��i����O|�d�O*�D�<���Z���[\0���{}�A���-r��IП\�Ia�	ПX�=��&PuE����i�1z0���k�]}�'���'��I�n�:-�J|*��\��2X���kc�?���b�4�?�H>����?�D�C�؜�1G��U�]�ʔ0 qm���������I
ǰ1�O�"�'�����(X�	�" �THN�q7��w_`O��D�<9���h��u���8�����!§|�<�J��[9�M/O�i)�Ɍ¦��������<%�'�L"�h�qT���J5{K<�Vը��'��L<����y�*�C��0	B��!��Φ��� �ϟH��]yR�O-�\yB�7� �$�蛪~pXhZ�gB8 �S��w,=�S�'!,j���bޒ��ө���h�C:���J��:eY��' �=����%&�� �5��:$�\��
��`l����8�T��RD�}�lрЮ�J7��)c�W�?i�p�N ���	5��$�$��>j.H���b��4{��Ew��pp��$SH� fF'&�r� �I���!��xR����@H����h��9k8Y`�D-2�vT�f.B�#�<Đ�j�:^t�J�M�%�������O��$�O��DR V�>���O�S ����.�I�
H8d⁈5���/�B��Q̜uO�Y�&����O0|	��0)��²���m�e|$Ț�bHG|��K��+���r�δ�O��q��'��Þ �V�[�KW?p��*DJ�9!ў�Dr��TT4q����i?x�)��y�o��jpBgŁK~�	�#�Y��yz`��Yy"#��d���?�,��<�P���v��	O7g��I�Q�J6tUj�d�O0�D� ,Ax�2Tg���O��!coX�]�QP6�۟k�z�<9�/ɑ/�D�2`��j�q���`�*��;R��A'�I���I5	-��d�O��?Q�a��bh�,P���a�e�(��I�.|��#��H��D@���)6`����E�	#P�!�G��rW,����<0�T�	�>���*�O���|�F!���?���?q���*��Ez%��m����D_�nY�aIP� 7�9��@�8�*��b>�d��tiTx��jA�=���N���3�aHn�ȼ��
�G	<�)�� 12��:��XJ�#\%B��x�B.� ���	韜��'��}����#�$p�V���x����F�D�q��N�vɴ1ZFKV+ƍGx2�:�S���В6et�%hUA[ �v�
:f���'��� w*��k���'��'_"�]�����]Wj�J�hX�{�ѨS%ʲ9�H����^չ�fݖ	u2�����?�=)��֔V,�a����!�L��܋��F:jƭi�ɀ,
 �g�'(��:��%@o(	���5A�41H�'�$Z����=I�FÍ��ir�
�U�|Yኝn�<�$��6����S�6̜8��Q(A���"|2��O�<ț�
{�x�8@�G�W°�kEN�9�b�'�"�'$Q�C�'�B?�>
�G�.)��!�E��	sNIC�� ��Ǆ�?��܅�	�u�P���E�+_���c�| P�@��|�De��d�ϰ=�韠�	$BI�5D��f2"$@/Y,�B�	+T7&0!�!4k�*J�`��C�I&h(�p����Lh,��T`_�.$����'^2x*qfq�f���O�ʧ|V��[��ïc��A*��<5�
`�?�?i���?у�P��?	�y*��maB O�"
���P"^!�r����	�or(�
���.
�v �P�܄a�lY  �TF�'�De(���h��=�f�U�Y���$6`�j"O8�v)Ιh��,@��X*�� ��'GO��c����%�]H8��fZ
�y�J�v�7��O`�$�|R%̮�?1��?׋Z9�&d�tψ� �i��c��y�B�4�κɘ���I7}��(�	W�j��5��G��uõ�L�t���"~������ hlA05�3# m��x���Ο���d~�����H`=��7�o�Z�+g�Q�y�'��}��϶*g��` �� i��������O��Gzʟ��2g��<~��xdi�a�d��J�O*��C�P���ّ��O���O�������?���ƒ!�r�aIݯ1F�ib�,A=<Ϛ6���c��� �i^�	��hO\� ��i�+��.�ŪQ�ؐ�M��eC8V�""�G/j["�3ړo��Pj���)Uϼ\y'.&� U��M�N�������v���7:9��l^
6B�x+QF�1!�$A<&:4Yb&�'X?Bq�K3WL�9Dzʟ��n�H�i �i����k�24r�MxV���N�²�'��'�2��,�R�' �IV0W�'|�)k�/.(�t9�r�H�8mQ�wA��'n�m*v�Q�pDZq���u�����O��-�	ߟ$�Gx8D��E[Q�u�Ѓ:D�X�e
���y@�~�`���6D�4�B��#T���WC�M�j�gi���=yƜ 8V��'�BY>�R$�ٙ=�8%#Bπ*5~�؀E�Glʘ��	�(��	y����ʗ�����)ߨS��ɀ���䆁�HИP6Q���VE�3a��I B �5�DI�6��4��:
�ZY�T	ժl�L���]��(O�m� �'�����'���	���FmU�&!��#^� �0�'��O?牗��˥@�%��ƫ	��$ O�	�I���O�[��Q��a�`�>�	&1Rɳݴ�?I���	�ڼ�d�Op�ĝ�[�R���-Y'.��UkSd�$-���&��O�c��g��� "5�B��I��0���Pj�Q'��H�#<E���SvX�qo�5V�r����� b;��?��y���'K�Qp�퉻M�a�4�*�<���'����Q�\(jH�;�h�K�l�ی�AR����K�xƪ�ZF���:����6�D�k�2�$�O�� �G �H���Oj���O�Ů��?�;Z�8�!15K��,"R��![6��21tɇ�I�E$b��5g��D�����l� ����<w���d�~=��+�N�i����,���_�s��'Th4�#@��n��5�ʇJ��!�
�'kv�;FP�,�z�*ee�&��HC�(�S�O��h
�Fw�@���*\�in�5P��I{��
d�O`�D�O��d�<6B��O��S�L��-�`�ٕ��Y)�.^k�s���}���`��C�Xh���'*�
����!~Nك#��N�L��gǙ}:>�j���~���fIE8����'���	
���J�nA�<Jb ��hذ�ў�G��ؼA?p����5*��-H�O��y�G'JYeN
k�� B���,�y�O�>a.O~�3��֦u�I��T�O12�����4N;@��6HT6�<d��,Ų7�'��+�=�b�T>��3ә3C��a��q��Dh5�5�u|�]G��ń�|�%!�_g�,p�����(OFH���'�>I�!L�J���3lK�q U�;D���B.�	`���n�Mk��`0Tc?�O,�$��)��|��	�!L4�`G�`��&���M����?,��i��Ol�d�Ot�Ct�@�$9�����Ō�%�@U�tuN�CA��!��S���'��(�̆�#k��#ъ� ��W�ǘ;��<Qa`d�)�矈H& ��[ED���#D�f�4��d@m��
�M��i����O��c�$�k��`�s�<��1O��d(�O�Ax5��5M�@m@��]�+p��5ቬ�HO��'!��� iH}5|�P�[������?�GdѶt4T$b���?��?�@��N���O��6.�r�(�dl�y^,���OJ,��'v� pp�Q#��b��@�,��R�'�ę!�hL�E�5�ա�
QC~ ��
�m��D��x���R���X���F/a�y�E)-D��u���p:�pqCƑ+ u@�h��HO>Y{�L�/�MC��x�Aa�$�EP&����?����?��i����?���$����KD{���sɗ�-���3�H�;{(L�$�F8�|#��?w8�b�F�{���s�S:4	�W��-
4����i�$=� �����ӟ����J^�Y�G�& ʔ���Æ�Ms�����*��}���B!l�h����I��hH�ގ!�䛄@�D��Ҧj#�`3�8G������4�hO�OlA s`M���@�W8X�"Ot�1gE��Y�@� 	�8�4d)�"O `�:��"B��*��0QR"O�Ġ1`B�o�|\�e�Vu�\x`�"O�p�WI"W�X��S~��"O�D �O�M�%�'��z3���"OzX���βi�B�lQ�0;,\*a"O���o@�vz�0�K�[�ܱ8"OK)��|�!�& Ԩ����y�MP$5���A�.�2�	�T�Z<�y�/&:�Hb����\�KȖ��y�L�7�b)iV�ނ:*� ���y�I��8�n��s�/H�E���
(�yrN -h��-�'�Q��l�JUڹ�yRg��H1t� )�La���Љ�y���W?0��+B�\;�A�y"JC�)��N���]{6����y�iA�G�ޱ�v��~��b딾�y�$^��`� @o�$#h�X�F�3�y�J�+Vz� J�.O01c�NE��y��N7z��y�,lLu�B����yB��0���k���6��<� ]%�y"'ԨR��JO��<��ϱ�yr�FE�3�������R�\��yr�¾$�Ԩ�RoַP���rO+�y
� t�#3BO�kc>Az4��3_4��@"Oa0��y���B�uK��@"O�!��	[�RMRƈ͈v!�y�"OL̈ŬF6'��xɠ��LZ��"O��B���r ���aGE�j��b"O�Y��dÉ:,��� [&(У"O
̋���L���gc��c ެ9"Oj��Gԩd�0<B����P"O�u�bΟS�<����M,�tP�"O�!���4^��P�WK2�ȴ"�"ODyDd��ڌ�i�G�Vq��8Of0ZA�̺z���0���"~��N?"Z�=�A&5�J��J�d�<Q���f��7�^x��4� A�_~"o߿>�l�)���0<I`F@�i1l[v��'�6}Y�/_V���/J 7
����\�]&($h�9h�����kG#|��C�	wX�;��4�eڲ�B�3��">�c� �p/���Ap̧Z�d����E�y"�Db`(�s7b�ȓ�P�H��@�$�"��'�@�l]̓P��
*S]yb�䧈�|���<6��D�ч��yʧ"Or�@��P�}_���f�Δ&x0R���Q��-E�Z�1O8�+�.�:]NJ��B�))��%��'��E�\�r-:��F(J����
	WW���T����xRa˵5����_�f�FPs�����O:L�6�ֱ_���+U�	��}�rApD+̬W�����g!�D�Wܤ��C���BѲ�
E�@���L�_2t��P+//��)���95�� {�NQ����$
��5��r�ܐi'킈Q�D<If�[�	ƚ��'�ʩ8̇�:��.����6f�F���!Y�:�8��I}��P��O~�8D�'�a��#1LY\�ش�w�"���$C�.6d1�� �]qn�� >��tH�E&C�(�b4��2��'۴�{E��7D*�1�!�-"��{����t"�:��,����{�-��ɋ���22��Woy��
���O����ďc�!�ă- �XP*�C#MS�]��� W�B����֥$�)��Uf�,+3�&��x"�����C䉳|$\��dLI _BL��t��"��h�U� B�ax�$�|�\����1��R*W�x�<��[��
k�(h�g	���p�c��0�8�4��(#����&��6A��hW�0�O�+�,�,ZE���F�E������0g��TyP�9$�,�l�<���SS�7c�p��W>�e2�왃I�<��>���}�ةW(U!uLQ�� :D�d2!"X%|h����96X$��ZS��T�����Y�Zq�g�i��QE�,O�Ȳr�+�<���+�!0&��bj�./�c��F��'�ܼrfH� Dz$��J�������'4 ��P��8ܢ�@Yi8�8�*Q2&H5�'B
��kA��O��U��HO
��)��δ���پ��Qŏ�It\1\����@=3���x`�� ��>��J���ǀ֏m���"E̓R����*�1
`��FQ�<�h�>Y�p��_�������Z�ʱ��3�I;r	Y��	���yCEԯR"�u�@�ppE� �w�D�Qb:a"v̞�����^F������%� �[Њ׉P@N�(E�E*�p<�@+Ԧ\4z�x���/>1��圁J4Bl�A��w?������M��"?�b"��4T�׾,C�ɒf�`#$�a"�>�!ł\@FI ߴw��/�0��	3	�Ē%gJ�-@U�!v�#B�Z��O Hrl h�'>�9��7��,���I?-��s�됻sa\�y7cݲ�HO�Ĭ�V{��2^P��ѝւ�SE�a��'�%Q��+�)�	�(o(���ا"�:���XNH8ip��3RN	*2 �zp��"#��'�:�cϋ�:'��z�11rh�{⁙=$�8;�D�;�%� ����wHR/ �B�S�EH,&Tѧ*�������
5\��3�jR5�0>��,]O"y�N��{Vb��kٶ|촱��'o4X�c-F`>�l���^;� {����T>��nJ>
��T�MHh)X�
7,O�9W����t�x�YE" ��sqǉQ38yH�W��b�IXyʟ �y� ��K�N���wT���'�hԮh�2+S/�t���:�Ѡ6��9R90oS�`U�h@�ۣv�bt�'A�	��ޗmx��+W�a��lH��� B�P��?�(XY�$"&�h���I(Z�!�#K%k˔%A��w�6�I3sxD�v/ -2Y<�[P�Y�)�5�0�W�(w� �̓]����˝w�څ8à�9�l-�7&�O��{��M�SF)��Ƃ<������$Y�2��q�r�9!�Ҹe�@�c"O|DP0($�880�m#W=T���W$E@�����$prd �.z�Z%c����9fzz�����/�]hr� �O:m���T��ZxX���`������j?P�6#[�m?�2+�5(^M�E��M�Q�
��Ḏ[�0`��?�����ُꑞ�R#��/�4J�?"~�����>ɑ�	5�AV�
�V ���5����^�R�i�!��ai�4;t����R���u��Z��q�j��59p7m=W<�ZD� nP�2�.�m$ў�=u;���00��AF��eR����?�Ri�*#�0=�!��1?n�X`
jf�0��I'����-]�L�@�w�DɍW��L0�B?hb��T!-�O��@A�R:H�p)��;]����AkO� Ȯ�� Dx�'�@�� �-���Ec_�`H��(OH�{�1\���W� �+c�I9[�ּ���O��\�wē��:|�ʣL^�)i։^�g��I��oA�|J�3�&�4z2Ë���Oh�:M��kM昒�
��� SеiG��2s��<�V@��B: �����ͻ5@\�^#\�<�����	LнY'4�OB�ؑ�3u�\v��6���!D�]i:1��	�v��9��I��F�+*>�@�9�Ա2�'�֨a%l�	�)�Cbڒ,�.��D�G{����>�l�(�Gjʲl`.��T�����'����ƌCDU�1��69h���Y`hš5�@#�h��E�#F���OE[$�SFB�-�\��hM	M��dR�MR%������� ֕��?���(��j�\02pC�!�1��29.&I�+� �d�C*3G;��>b��* �ɳG��RxXa���O�a�L���W.F��Ǫ��\���޼�N��%���=$Z}����tRs�OyZ��I���#�b��z�)r�O1���h��V� ��xҤɓ;�\Ԣ���qY��ΘOUb��DD��܈�e��.L2T�Oh�f��}�k�brnyn�(�y�.O�`�0�l�&�����2'�D a&�>9��aF��<�}�4�<1ڐ8$�2;�t�a�D�T�z����(�w�~�̐*��KO�'�֨���q�eB��!v� �j,���%~� P�� ��$` -��2�M��
Dl�@&GȄE��m�q	V�1�L���8I�#�ؠ
˞�B�i�)\��ɉ&?ʜ-�'�љ����i��ɂ�H���W�F�g���!$�_B�Q��'���B���zY�V���Í��~�\�KS!TD�U2���x\y��O"!��R�IT�%>O�8*�Q�A�,�WEݮd4�b�ቤ��I�'C�u%>s�T�s7��c�l�$F���(:�¸�����=� M�=�u�c�g0\)q���{�	c8L	%�t�g�.'�\(s���[?��L��R\��E?n���c'D��𒇚8�>x���gj��qo"�	�K�z���g#�S�00��Im�¼��L�!d��hr��`�JB�I�xI�T����>�! ��;'�B���^����+O�%	U"_�;]1���3�:M3�k�&Q&���.|�6B�	�5V�ͩ��-ޒ�j�C[��p�Yg�ɼ*K���`%�k��`�B��Wk��1O36���*��#LOz����	;+`h��gRP�^�I ˏ/�BQʗ F�Dk��Z�"O�y tAU�+����V/�?~�$�$�E�~� ,a��&&�%|�D�k2� 
V�V�Re�".�3"OP�`�i�h ����G� ��E.Z�q�@m8��z�	*y��0�u�ȹ��_��ڱhA��vO��O�#Q�MA�Sܧg�@�R$��'8�8��m���t�+��|���V)�F߉V�@�?��%�( �����^�n����EB`�x���¢!�>�҃�:Y��Ha&mI�`�%�_�G�����KV2JĊ��Q��_'|D;r��Zx�d{���.)��`�eE\�6�8PD��V�.�҂Q��x�աBڄ��sm�&l�1ȴ��@�H���г��tå��-:����'�2�sR�h̓v��qЎӡs͚�S J�5vd@�fk.g-�9Ѡ�eh|��Od�'aWt��'���x�ݴ1�ּ���U!��CI<9�MȩF0�O1�^=	R�K�/Z8xq�D� `Bh����$]�e����'g��*��/��8V�I�w��8�كn�H�:���Z-����ɣ.H�9�ؼ:�x�ymC�a��ʅ�.K:8ӰB�.��%Z" _�ذ?� �ֿ[��@��M¤��#R�'Amv����g�HRN|*@ ��$,L��5��*B��4(  L�<���'~-�j�#$���#��X�r��@-�8$�"~r!@��XpL#uf�;�c���y
� �`�w��:�*0�@�ژ?60u�"O�p+���X�:����_E�a( "O�x�g�-&�T5����8%N>m��"OR�zSe�;#� x��]f�J�"O��x
b��ܑp�#EZJ��"O,�ˌ����u%�\y9�"O�����C��t� 4�Jz�j��!"Ov9���f��̠�ÝL����"O��C���I���� `��"OD!���=�D;�H���p�5"O�|���şT	���#l��\�~� �"O�<�\�D�ȕ2�r
��g"O�h�4	_%pQ𒈖D��41�"Oj���H u������C�P�V"O�DsT��0�@Q$�C�z�l��U"Oj���_�{x��p�Ï�6�R�Z�"O`Y8q�J1W�T�b��'�T8�w"O�p�!o�B�Npq�(׵�t�w"O�����C�~� ��0S�15"O6�c��kMʸ8��S�4ل�(�"Oԭ8��:�����$Ԣ|�=!E"O��a��! ��9�)(��3g"O���p�'�"�6�5R�R�� "O��C�eϨ9�9aV&��x�0�"OB(��hS��.x�Xf�,�*�"O"�Q�f��Zm:�a�m�o�y�w"O��QA����|Q�b?i�\`*6"O��&^)` �}�f^���:�"O�L����F""d�0��x�J�"O����CS�����So�&o�]br"O�M8V!��+�$�Ѩ��!���f"O���#)ƒ�z�e��-���� "ON����(�	���J�m��Q8�"O�eB�$�sj0�F�v��*�"O�1iVGڑn���5�
r;��t"O�,��"W�}�JS� P�P@"Oƥx�邮0�u`득*Uqf"O��@풄?�N k @Q��VV"O�	���-|t���
0j�`��U"O*I�Rh�,I��C�bɭY���"O~�j2����$����6YG|��"O¬(5N��t���`�
^���3"O���$(A�d�`j@��d��%*�"OpT"@�κ�(���"t{���C"O6�(�L��ࢶcѴs<�pd"Oe�ĉ��V�v�Hѫ�Fj.�;�"OJ�y3�٧sc��Q$�Ieul�p�"O��� Qw��D	D�k� ���'
|y��O��=���StJ/S����'E�xk` ܍=��`��4~�e*�'��豁�@t���)3�^	��'�Q�5�"M��r�M�8s�x���'�����'��f�٢'��-k�@�k�'@���G_NL0A����O14(��'Ɛ���C�"4�D���ުN(��' ��ۇ쀦/�n���.ƖD��|��'k�����׋jq��LO�?�V!�'W�@�ɏ�n���8��:;�L��
�'7� ����0a���� `qZ	�'/�0�P��'%@�h��d������'�UT�!mb�y���4��9�'�f!4�L�tCC�)����'&t;0G� ��!�‌�v�y��'U$LQRIB�P�Ȣ���v���C��� Ҙy���<x�a�7���W"Oj��튿JB0PQ��ǰ-�R�ɓ"O�	���k��� Qv�Z*�"Ox�p F�-#D
D"��#v�v �T"O����D](e>��#.��p�"O�,ĀWV���{v�L8I�8��!"O�M1��P�h4Ƭ��H�,<s�=�U"O
��N;N���M�<m�E�r"OpTJ�fD��ְ92��6�(3"O`P�
՞6�� i�>m��ȓ�$��]�;�qÅ΃4��ȓI���سl<���b�/L [f@�ȓ{,e[Vˎ 0S5-�#�����83�U�aW}LL��_�����ȓ_4Xe���ˮ<�H �B�˧�f5��r����H��W�4��p��:/<a�ȓ"c 1��%�7f�i�4-��Vڈ���<8�B��D4ib$��Q.& �� y�ܰgj2<|D�Y�hY-t^|��ȓ:b&M �n� �������C��=�ȓ(C#��H��֠˭bXD��ȓ`oX�fU0�*���gL6��Q R����@�z�������CO�l�ȓV�B�ň�k �C0�F�A�^��ȓ0tJ�G�0Lo�����	�XsZ���_��X�kF96�deB
Y1��P��ii2A̢~@��)���
>��i�ȓiQ�[����8t�1%eZ2\,��ȓc(��Uɉ�,��WaO�=q�a��U�J�!5̈���Dš&W�<��3�DB�ن��Bώ�Hb�p�ȓh,��b��'d���&�|�z���/A4r���`3������+7t��ȓ�61'@^; �>����܏Cf����z�Н����@�|d0�F�F_��ȓWĄR�`V$zt���/�?��؄ȓw:h�`3@����k��/@bp�ȓ7Ѻ�RŤ��=b@R eW)1l����RR�R�mg��	Ѣz��9��0D��i'%Sg����kD�
X�}��.D��`ŋ��F�"aI�JF�t; �*D��@`�H	f`�C�灥"�h<X�+4D��R�.���w��/ nPhR�>D�HX&Nڦ1ٰѫ�#M�q�8��/D����A�m�H�2�P5$��!�.D�,�ӎB�u�vUR%��4��!�%D0D���q%��jr��� ��<���c'.0D������g� A
�<��8�F
3D�PF$��%�s+� x|t0�ao6D��8���I����&��7�F,�7�!D�tEL]G��S�ȬW��
�>D�����O{��`[� �N�����	>D�����C�C
vA�P�xJ�d;D�����۔[��h�fæې���;D�p���I)Czb�D/��~<��9D�Lb6��-�2�3G*��!��H68D�Ё/+n��0��EIfP0��0D����f�7�^�;!(� Djī.D��S��G�ƌk6%��Z���Vm+D�p���Կ	�l@v�FB�sd+D�, ���I��1�E�.��J<D��[RF��W��<��b�� �����>����ӥ4DD��_�L���¤�
+ӲC�&6�R$h$ˊ�+�z�	�Z�C�)� Ji�%�3����m�0ND���"Or�0��"��; �7r̚�  "O��K�< ���Z�g�����"O�aQ���8u����U� �T�J�"OnCFC͕MAS��,�:eI�"ORT3#�X1z&^��&O��8�4"O������?--P��̶[�C�"O�a�2t ��t#��&�$�h&"O�\�4�C��4yr�a�#e��}ʔ"O�x�e+>4q��F�\OҰZW"O��[Fi	b�`�0,_;`-Z���"O@	�q��l�#1  �\*}YW"O���p�Z,n8�G�d�R��"O�	�H.3L�d���q��ɑ�"Ox������n�ɂO�QZ�q0�"O�ɘa�O�Ȍ� O��/�@5`��O0��-�)ڧ)`搈����y�����JT�y��Є�q�<�@Q�	�uxN5�u��+�������D�E�ʺ���qq��U��	D����"����s�V���A�g��a:�#8D� 	���q�Jq�b��E��t2FF:<O�����925��0���!@�(03E +�!��N\�4Xy��TC��Q���s��$�S�Od��sǙ~&��b�� #�|U��'f���A�&?��4� �̘`�Q�<���)�'3�J����n��0�C�-�ȓ?��{ֈOVHXq#�90(��L�������\,�C��ɘI��>�����j�2(�jP$V�xA�lb��߀�y��&?ʉa�o�(���y-�73|d�`N�<>|��s��y�(�K���aVB�%/*����f��yr�f��a)׎|�]Q�	Y�y(d�V��rh�%w2	�5I�yr�1Xݮ�s����z����7�M9�y"!R�
��)�˜�q��@4��0�y&��m��,��k;nk��SgЎ�y"	�h�nX�3�j�����M��y���!��D[�8�$D��yr�ʂc$ࢠ�}��8�"�'�ybo)i��旸F�,E�Sj�y��JiR�0$�&;��u[S-I0�yBǅ�^[fu{UI���NĊa�	�ylG�^KȴC#'�����gO��y� ۆr��]����+`s��
Ў�yR��PK�qc��U7n 2�H2�yr��3�m�R�	2k�Y���4�y�+_7'�����?� �I�yR&�q ¹K���(��ՈZ6�y2�^#]Ixy 󬉎D	xD�M'�y2DЋc(�L�Ń}�`l�d=�y��@w�0�ś��������y�l`�t(pF�9�!��K��y�#"'��ɺ��ޘM���U���y� G�t:���*4��� ���HO�x��I��`I8��W/ lM&/�59�C䉭�Zҗ�NM��8Pe޴(��
O�Q�JƏ9M��[�K�.�3�"O<�,�ΨI���4�JM��"ON�(�	ˬ��d0�%#$�6\a�v���'0�N�x�V'>�7��(w5Ɇ���?�P3[��Pz�i�P�>a�`�l�<)ׅ֖*s�h1��m4L��-�k�<�q`7�t�5C=��	�f�`�<� �ݲ�/����0�δ���1�"O�ta���Κ�sԌ�UR@,+�"O�Yp�cT�T�Hل��68N%z@"O21��DJ�+ ��Sgƍ:+0 �"O�\�&�$L)�˛<_` �"OȐi��T!P�8��U�N蔝K""OH��@��$D�b���H�p:V�!5"O�Ds7ř�� �h�=����"O��hFlH�<b��	��W�z�Q�"O���t	�|z�1#�hv��%K�"O�P�pO�`�d!�����DK�"O� �uEH�5�Fl�t�^�jvx�c�"O�A��"��~(Є�lO�j�"O���"BW�>z%;���,Ӡ<HG"O�!qE�@KU��#�S>>���8f"O�A�F�]�p���J�$��x�"O����ձ:'��@�oY5� ��"O�� s)G4ẍ%�"���j{f�@�"OP	�u�Ó5���&�W7I�f(�2"Oh�0&,ٰA�ؔzf/�&eT���T"O���U�o�&,S�UupZ5sd"O�ػ��M�UW�D���R	p$��"O����_�Fr�#Y�r�1U"Ot:��M!g��{ ax����"O:e4mF�6�`| f�Ѯ3_d��f"O`���ĩ:Z ���D�e�6 �"O�DCS��z:�H��z�Dja"O<,�m��M��Ṗ��.���J"O����L
�(��ө��`n��B�"O����0Ϟ�iŉ۬m1\7j-D�,q�g�Ҏ�I�	T�aP��`%1D�H2W��&p����R�`!<`y&�-D�̛��8Bu�/c�
��2	,D�;���x��p�P�$$�y�e`5D�HY����y\��pѩ�G�d"�"2D�(�aA�9φp��!�v�:]
�0D��C���ey���uB�:ܤr��1D�����E1��&d�7ྸ@�/D����0c,Z$�3aڈ.�����8D�Lz�X�txHs&@�l�����a7D�l`oJv�m��)∀*$"D�hC� #-�,(� �J@:��$D���1yc�4����c��r�$D��#��!R.�ܚ%��MBL�jF�!D��¢��c�|JD� f<<a�-D��s��<j�YpgF� �XSo)D��� �̚���瑞G �졖:D��;������0"N�\֌��,7D�`1�f����H��
>��(k %8D��רŀAJ=��H�'����A3D�Lq ��+#�<1��1���F/T�8���U�]U"<btA״=:�Q�G"O>��!�-	���1g�B�w̈�0"O�4� 4'��)f�9��q3�"O�0i��A�5�$�D�'E�5j�"O��� Nȶ�`v�Vd܁�"O�ź� �ܚݢ�@�M>��"O���� ��	��9��˸51\��D"O
���Z |�!�)@A9�"O|�у�(#�HI2��K�6�"O�!p�d�D��<�G���غ�"Ox�X��Αr��s�o�k:vIc6"O�#>(�����.#,4���"O���6Ƅ-Zi���b&ּA�"O� ���ՙAh���c�)6��"O0FGS�D����o�L��0"O�d!��=2�j\*�0{ǰ���"O�����]rUz�p�/�(q��=R�"Ou(C+S�"�Z`YƎ�UK☺�"O�E��n�n9��(X}L�@��H�<�T*�8�yƫC�'Ӷ�Q`F�E�<�7�D�F�pA����<��{q$]�<q�K�2+��8����]G|�����X�<y2����Ϸ�VB�E�o�<�'��a߸��MM(���%��v�<�֏�|v�����ˡkl������V�<yƜ7-W@�K��J�b�P���$H�<"蚳]
�����<
�1b�C�<1AC�?6RDQ�B���j��iy�<���7#�\��g�#Y"��QW�[M�<)6�C�N�h�F��� a�eP�<YI8�R1�d�[OxY	���G�<�f�Se�����:Ud���@�<a���B�%� ���(D}�<iD꟏���B �*��pV�^�<!�ǰt7�#�ɞ�C�
��!�a�<���JN:\��̊�,�di��_�<!���8∑CB��5Br�(��P\�< ӊh�
`���Z�
�Y�HM�<9��	!�NUY�@�<cԬ)y�͘L�<�≘� �x�e>0Y��0�ŞA�<��|�ڡ��kٺ]`̕0����<����f@��!ꏺ8�T`0A��S�<qY�|��'��7R^v�##IPR�<���P4kM;�V52FNd3�[J�<�G���x�̐9q���I�<�ѩ^�7 ���F�
z!H�FB�<�bF�,<g!�C1&B`죕��v�<Y�I�^�Xs$m��*�� ��q�<�rG�$?�H��N����2�"r�<aK1M�Ԥ��#S�e�|����d�<�q�@
k��`Ce5x�t�J��^�<I�$̛v����R*ƴJo6١E@V�<IVo�:ʒ����upU��VG�<%�Z�߼,�Q�Y�L�n0��j�<�Wi�'��d�R��>�����b�<���l�DLxKυ1�@����x�<�2OʜI���"#X�R�`�-�v�<�bjҽzD|�Ao��+�dቤ�Y�<��MP:p�rV�	�<�̒]�<���&hv�A�g[F���`�U�<�eF�x�O�2�Дi��R�<a�ₖ,v�p��^�z<�D�CP�<Yv�ʈW�⢮��;vN�Y�K�F�<�b��Z���8be�� %�x�<�+��GWL��5"(�*�Dn�<ɗ"�$e��q����D1���^`�<�5 �;f�(1�$@�6��̒��IH�<9K�1_� �˃�}�v@꒎Jk�<!�� 4q�n�sS΋#�z ��&k�<!`�E�,�vi�-l��g�i�<Y�n
m��\����y����f�<9��B�|<�M���>�i"�J_�<a�cY c*�)9N�;��`B'%Y�<�����&��{�F�K@b
��
�'��̆����EU 2�5�	�'�N��!L����Q0Z<p�ʘ�
�'�,z��?5Dn%��ҳ����y
� *�jȉ3Q�\h-er��3"O�,Qo�fZ�����{>8�"Opy��C�5#w�!�W��=+��H�"OT���(	���ă�7&"�ȫ�"O�@�#�6K��DJ�V�1i�X d"O*�i�#
�8�R���rJvȀE"O����lޠl,	`��ܪ{<,�"Ov�x���xر�gڊ/�򝋧"O$Hɖ�̰T���@�	2�Ѻ�"O&�1�n	;A�D<��]�n�`Y7"O"lr�^ܞ`�Vn^�h���"O>�!M��]w~t9�ѨJ
��	s"OМd�)�,�@���5�4�B"OXY�#���TL-��jD7�t)�F"O �{��R�"$�
,I�b�m*5"OvɄIӱK">�c���Y߆��W"OeR���98��3v�L�p�v ��"O��b��1Lp�83����eUx K�"Oı+��	1E��ԀL� g���"Oz��SC�EJ%X�F��S\,
p"O�E�'�h��	צ�!e!~���"O��oN4j���F\����  "O:���a�$#< ���\��6��%"O �(���.Y�|���,�\�av"O�H��I= ������֯1�J\�"O��q��"a�Թ��	P/w�@��q"O���7B�]]���EjS"O�����EW2�
���f��"OP8+jU�@��#`$Vݨ�"O,ȉ0��"B�)�χ9}�"O�,cF�E�h"&DI*B���t"O4c�m�@&�T�@��l8�"O�|���T��k�*T{�\�"O��"�ІG4xH㩇�<9�5"O��+�i,v�L`�5�A�g���"O�d�@/��DG���tAG�' �Jd"O,�їK�����E�A=���$"O�\#��
t�[Aŏ�0��=�G"O6�*S�R�������6�(<x�"Or Hs�A2���X
�G䘰��"O�	rG��:а�wҔ"5"O����	�m��P	�'@�pl����W�<����7���2mƯ�(@�BL:cC�I�ҰP�'��y�d�R��H�C�ɧb�����A��D��ҍ�]<6B�	�{��%C�nMa,�)�DJ#�C��3�>`���3����dH�~�C�	�b�F�9dN
+�2��B��B䉱�M�f���C���Q��
0X����	F�'�Dh$ B�	� �
A$Vj�p)
�'�*Ex ސD�0<�ю�*�|3
�'�� P��

D��p�������'�t3�-u��Z�@=ro���',��S� �Oa��ҭ�[Pyi�'����B�w������ͱA���'X���*�[1h�q�n֙?�|�!���hO?A����;��Ku$4B�8�9�Ār�<�F8B4�59�F��箚p�<Q��� cD5p#��;"O�`�ak�i�<Y���7;"@j^�c�m�X^���9���1�-�/�pu#fUB�<��#|�! qbC$VBݡ�ǆS�-�ȓS�xeb�/E"x-�h���3�]�ȓt���O�������}\4���S�? *-�e��@�z�r@���܈�"Of��Ձ��e�	�
N�'Ct���"O,�z���ONm�
�.1��"OLD�K2&<Z3SIҖ4���#�"O�����S,8i0)�.Dw8��u"O� c�	��p\)�̓l傕"O��B�FƿQavٰr�ٺukP�S�"O-;E
=~&�a�j�HdD���"O\�W'W��v��0KT FIZ"OFx��'˓st�����/{���"O� A#.� �@L;���U�	|y"4O�qH�)3�9�h3tD�g�IV>���V#*��B(	99ι��O?��e����pP}�䜢(E���ڌP C�	(:I
��T�)c��{���r��B��Z�rP��j$��z1HZ�RB�B�Icn���Ђ�T����C>e��B� Wm*���Ɓv�N!� J�.�������L�'��'F�2�ʲb�X-���lP�Y5"O�d(w��N ̕��h�%q9��)�|"�)��T^x�A%摡9n��5��*DHZC�I,+5�s#ф7����r��<<�B䉗b�W��iƼ��%KWqxC�	(w`�hQ��@����M~YlC�I�z׮�ڂM�de�Q��F��s��D�O�ࢄ�K�/��y�Vᆟ29��m,�O��I�� u�s@)W�ӧ�9QS���G{J?��V�L�/����m�E`.�2#�*D�[&�VdT����1dM<����'D��х�Y�B�>Չ��'T�}�C$D�$�T���
����[#=S��'D���
+J�����Z�LC��S���OH�=E��'B|���ZQ���A*��w�PQ�"O|@�rfJ;xa�e	�5vO�d��"O$���B��]2���0ME��ᡓ|��)�S́�#�_�*R�Դh�'�h��TaBL����	����'ei#f*�~���댍;�Q�'D����P�(����'��ƨ���?��� �l �8d�P"�~�b	�'�(����I�\�x�nY�v#����'�Q��"Ć8Iԡ�2��m�.pH�'������j3@��m�_�H��'c��0qN۸Z�P��ՆY�(�'��q�4
ɑJ\�A1�m�
���
	�'���1�hE�d�1L��B� 	�'V8sFK�,|�
�j��-v6h�C/O�D?�)ʧ~��]Q���+(��O�4+6P��ȓ\���ס%Y���CB:	���ԟ��?E�$��'�*�pĂ�=�X�á�ì1�!�J+�z�1Ϙ�i�*���KL8f{!��:��< ��{ԼݻV�P!��+eN��R�>ebŨ�,� 9!��+�&ѻ�
�hf���텎{Jў��I��B�v�;'� �rHF����܈ !��_ >J�2J�J8�� �*��9���)�'ϸ�Y!?E�}8�-H�EĖC�'�0��
�]��ґK�kd|�I�'p��1׌.�����T/��@�'B�x	��G,ql`���4D ԙ���hO?����X�}�*�8u�@���1AJ�d�<�զp��Rʉ�+9�IU�Xb�<qa&�
�Z ��"��j�*��G�<q��F�<��*��;ήiz���A�<� �9��H�r�sb�/v�z�Y�"Oذ:�*��kd�5!�	7V�T���"O�A���K�$�e	ܓ6{tm��"O)����	f�L�J�唝pf�zC�'�!��35��=j%���S.Ah����!�$˳U��D�D��p�ڼ+��^?1�!��!R���bOU���A(��޸S�!��R�n� 1P�ďa�
�!�$^�!���4L����&�h�>r�@��!�Y�
���Z�k�"N��Q�ε���AHa�l4���m<�O~�=�}�'b�P��ZP"I����0�Lfh<)WN��{��A
�Hޛ}R�<�p�P����0>�pOȨG,�D;	Y��
P�/Z�<I�����Be0�T�'+Șe[�B䉆Ը��$�42w�)[r�\;~zC��?�e�n�$)�a*Ռni@C䉳a�}CB�U5Uߖ��%Kd���1?�&��g�rÈ9�� J��a��r�p��!��d\�;��)n�������OB���#z�X��"�Rrd	5C^�"C�Ɍ"��!�u�#U��U�_ 1I�B��;!��I�w�#J0D�8��OӬB�F_8�%˂<Ɉ���I��C�I	w?ӆKόbz
9�vO�8.�B�I2�\�ui�#3��C���[�
B�ɵIr�5P#,v� �d V'��H�鉳7@R}�d��j���ZC\�r�C�	��x(�v.�?��ة�%ٲa�C�Ɇ0u>�"���c��\�jV�-*"B䉯>t.@�f�C�@Pv
�:\f���)扱o��=R2A���\YQ��8}�O���'�)�Se���7��1M������+I6�C�	�;�CC��0.�8�C�n@�yڞC䉷ve���g'��_�p�6f��M>xC�I�l'b�E��[�<I�J�@��C�'K��U�Ɗ:+�.t'h�"O���p�Rr�[�ba� *��
"O�)��Idp�A`H��9"OPJ/C$H��I	, 8��Ԁ�"Od�`�K1�.ؒ�jD<V<p�"ORh'�Ϸ47���k��}��Q0!"O҈s�A3a�4�RHN�x@��"O򌹆�ِnF�����m�P�a�"Otq���#��@�5�'�q�"OƽãJ�H�A�#��s@��c�"O��%�I.�t�����I4�(��"OD�8.P 0?�)J#*��X7"O��sF
G��aF�_�&)J4jA"O������f40�ƍ�"�r"O�����@O����E
X�����*O��9��?h^��щ�&S��I{�'����_�$g4,�2i�9n���'Y����D��4#�]�@�R�&-�J>���0=A F�~�h�y&��UPԭDo�y�<A5/�	6�P�VJ[�J�D �r��v�<af�ۜB�2�7��5N�����t�<�jڭ-�|�TBZ?�u�� �s�<�F�&�*Y fiN�6�ۑ��U�<!$��<��d�%���?@:�2C�U�<Y��F��0�U�o��Z��Tٟ�$���I=z����
��d�pt�#@�,b��B�+zJ��`F�_B��`a��|B��n�
��ȃ/�T�YS�6[lB�)� ~��卾W������8e� �K"O&�Z2�S�
����TA������"Oĭ�a�U2��ҁnǶ8���"O��#4�S�a�����23�ft�Y���	x�`#�M1bG
�����pɞ�Q�d1D�X�ǖ�r6��R���iP8	��e-D�x#�*R5��KC�уP0���-D� y� �1g��삣�P�4h:p	A�'D� ���6*�|�p��E&\���#D��a�D�E� �"��`)(C�I
>��y��'|1O�	zsV"�%�vOV�l9���_���	'a�h(�#�Z/c�-A��$��C�4����D��%� %Xb� �X(hC�	>	^�@H%�4�4��Jݛ� C�I����"ּ'�dU���Fh�B��=|<�5�4<g0݃cbI�BD�B��#z���d��Uթ�8E��B�(����)��S���7G4
�Oڣ=�}"CbĠ��Q�����ԒT�_�<c+W�*��=�#!��@�h��S_�<9�J��l�$�j�U�C)PĹb�A�<�áT\���T�~� �Påu�<iF��+��"� P�T�M� %�m�<!0�T�Gb*�EY�U�UGm�<G��[ڬI��ۥCF�)X��u�<@.ѥv����X=x� YrE	�p�<�G��Y�q�r��<!���r	�l�<����`N`�҃��^F�X!�-D�<iA�H�|V A�rg82ގ�*5�@~�<�$�3VM���ׅ	�D� !��n���0=y�
5w��G N�U�D��p�Sh�<	2b� �ɀ���*w!DT�6��k�<�t,=<�
Z笂�S�6����]�<a�Ј}�x�då	�L@a �A�<��<2-��9tH �w�e'��|�<�玸G�:p	�4!��ڢ�y�<y�O�1�@U��� �-�E�`��vy�'\UjHA��좠�[=X�u)	�'��!R&�0!�a��̘<8Z�A��'iC ���Gء�B��>dYp�'H�QWi��C�(�3�K�]�����'��c&�z�\�JrMRLe��'Lf��&�N�����;7�.�`�'p�r.:$�"�KȐ_��Z�'eNm0��/7�ȩZ��L�"?�@Ћ�'Oa�TQ":`1�%�
<u(L�Q2b1�yrMܴDe4Ap�hv*<�q���y�U"�� �4��c����$�ڷ�y�`�'Tx�q2n݌[`������yr%��Y�$�3�J޵T�\���ş�y�/[�^@�@昑GL�|C�hI+�y2� 5=	Z��Q�%��#>�y�.��L)�ܻr&�Mzּ�%䍁�yr�

X��܉H3Ԛf���y��B"tM�q�t	T�O� ����y�Nź����ՅE6>��	���yR�V�*�ti����/;��pP��G<�y�ɒ�d��
O$3�����`�+��$9�O�,J�֭��yb�e\/{��apC"OR�I%A�+u�
0s"g�;TG`�b"O`��L��w UYs抵OB�۶"O�u����q�I)�^H4�32"OD� p�8||��,XT2��b�"O�Dp��ݨ5�(Y�L�1dܣ�"O� ��v��0��%2���%��p�"Od��� �]�N|������tl��"Ol��&�+�����㐚;Ȋ��t�'��$�����X��aqR�D�y~�UK&7D�A
��|0�!Ӂ���x��� �O)D�XQ3*&)����@�tI��#`�(D� X �H6S$.QrN�.����,D���,8+o�D�d�-�Z����,D�,�AE�4@`���
\<ıt�$D����R0Q��ɪBH�tqL9���"D��huLU��h��A�K,��Y�!$D��+�֎�"	��D�%C?�d� !D���Ũ�J�����:��K0*;D��B�AU�8�h�NM�p��ӡ+D��:tȃ3pFܱs��/���d")D�p
�LC-���C��Oe�:�H'D���`��0ʤi��?(�8��0D�誠�Dy~�� �E 	l,9Q��9D�p�6b��9��0enֱjCF�S5b9D�X1RI�U{JX��jX*E^�U�8D���2FD�VKB�J�T�u�U��0D��g[�#<zЊ@oN54�Jы  2�O��
�Fa �aDI�X��cN�6vF{R�O� �ٖ�ڷW����s��8��1�K>����	Y�:�tӄ��
F�E�d'-Y��7[�>=I'kR�_���$ϖ�yr�-G�4!#ː��i��M��y�'W?;��`�W�Z!t�:!zE���y2�ӎE�lp�ք��`xÔ�Q���=����d�5����G,B.8�dIvq!�䗢q	���F&�V�(^�V!��;]�
�q!&ܞ+0\�E!�d�O������q�Le��O�*3!�DƫA �����6tv`� ��+F!�$�w�X��5k乲�B�% �!�d�'Z�<��կ�K+ 12�/w1!�M���"���|*���^ўp��	�T(��0w�H��Y�6���6B��/{3V��S�&~7��0�⎁X�B�I�� a0$Y�w���Ǒ���B�IE�-"e�_�;E�H�i�TB�I|��` �9���&
�s	C�ɒ�Lx�a�	<6��Ӥ�M�7��B䉒��Q@�}*�Y��̃Z_⟠���<q7n���a'ƴ`���ʱ[��B�I�s}� 1Ać"PN��`��\Q!�B䉑:d@��'Y�!K���@�7)�DC�ɴ2$Ԁ���.J̀D�����>NdB�I�3�DD�`D
H�6�+��A
�PB�	�\�D�Iq��Dl��5�8��$�Op�"~Q`��,���*gd�f=��z����''R�'���JCa˺B�vp�RcQuW��z�'h��3�G�RZ����j���N�k�'`JQ᎘&sB�)�F�v��'�R-�c��9��u��ׅ,�	
�'/���b�M0K�R ۔�L M񶈄ȓ=+q� +ޚcQ�)ٓ���p��$��є����3k� 4��,j��A������?���L�л�@L� �v��q�_�{����:D��`T�Ș0�(�X�G��e����-7D��8�lJ>b�14KP?f$�%��o6D�T;�-�0���۠�ͫmp�Ͳ�7D�\�C	[*r(�l�$�O�Q��ɨ��:D���3��md�}a��@4"��q��7D�� L!X�E	�_HU�w/W�6���"��d�On��I,'�h@�A�#y�h�)�L��!��/D�+��D0F5d�Q���y�!��8�����BM��^X���^4}�!�$�#r�n��(PNU�RiX/}!�Z�\�.,��oP�ng~	е���Bx!�d0&��p�@ �6V��F�Q�Y��i>�Dx2�
S�ZB��E�sV�|qeH+�y"k[;H�{�jU�kl��������'?az��@#S9��
�(Sd�	�4 ��yB��)��Qp��[�8��@�y�KR�6.45ZՎ�!St$�H��\��yB�2s� �u)�G�^�ؕ�τ�y�F)Z�����j;<���CEB�yB㞗	 ����U��j,9̏��y��Hi洠f�]�N�j�J��y,�� �cd�Πj��5	!Ά�y"Bǻv�ք��l�P�lqچ�t���c{乑� 	 X����X �̅�����5ꕹqU�9�m�.�b���P�Vm��뉤;��HQV�ȓA�i�NL
8���`�řC9���I/$x��Z�3)�!��.�4|��`?0Y2��C�py���|<���V�(�h�(��i!���`HP*���ȓe����H��:���(~��p��w�U*�
���Hx�6�9��B��Μ�(5��B��X���i���~�
�fΗBT� ���
*Ȝ�ȓt��H�a.T֊G]j()��vj5 � �N�����
_����� ��q�5B�,6´���	Uzn@��r�x}���e�޴Q�d�M3L��ȓjd����m׫J�%�'NJ#����u�z�b��G%cH:}H1M�"[<V-���X9C���Fa.�0C�^�'�fI�ȓP�5ӂ��7z����LDq(�ȓp��G��(.a�@-L�KS�ćȓ��u��(wZX�`�fE�����ȓ"L�x�e�BE�� Z<q� ̈́ȓT��zg&��K&��K�
:B^���~� 5ڳĔ'V2����;��`��	G~R��:Xi�E;7���_�|�R�'_�y�`�15\y�"-M�Sn<)[��H�y�h�BM�U!*J�@��[��y2�����ӑ���V��QŌ��y2��/Q%z��̞	 �!��5�yҡL�7��c���~�6�㖬\��yR�O78�2TL&aƄ�P�_��y"F�W���ME +�Ќ�Ɔ��y�C5�4)�beE1.�ʹA&�Į�y2g+_�y��K�rq�����D7�y��Ɓ=n� �'@�o��P�7�*�y��Z4��E��o�`�qvj1�y҇�j4��B��B*k��Q@�CU��yb��O�	�Bj�N��A�
*�y��?r��ղD�W�vmb��'ʳ�y�GĄM�߱��k���ɒϜ2�y�`P�hsn9`�T9������X��yOD/ ̭Ǩ^�+��	�C�/�y�j�`�9�o�-J8�S���y�f�:p�9�2K�+{��]kr�T-�yr%��~f�D��%�[�R`��y2�e�����`K�� 4��D���D�Ol��� H9�'c֮�T��"KZ�	k�"O��BH/a ���	�FI��6"O\������6�J(`�	�718b"O��HL*|�(0�cԩl (�!�"O� �s	ȏ���h�蝣"��0��"OȔj��_| *��<�"Er�"Ox��ޅ�1U�B�@���'��	S�41�ߵ~h�012㌴j���V�9D�X5@]45�����fL;1[Jq���8D�d���$B|y��=xH�!��5D�0��Цys1�ٖ	�Z��4b%�ybN��&��!��Pw�@���<�yR�Q�0Y�,�w��dCd���!_����6�O��)�"�V�+Q�X\`�2�'���')a|���N�8��`�|�@�� *�y���fI��H!�ѷS��"¤���yr���B�ƃ~�((�mH<!�t|{�'*��z`d՟!�P8
qh
�c_��z�'|�I�7O�0�%���!V�.���'Ѽb��])¨m���ɏSY�e��'�ص+�KS�MK������K�`l��'$ Yen�%�F�2(�*>�� Y�'Z$�rA�?<�l��AÞ�k�I�'�p,���3,,�*@(7�����'��hKW�D�ba�]*�E �+WT80�'���3�F�X���[P�*Xs*���'���(5d���"{�0��'6u��� }͐i9s���r)|p�'�>�9�͝\������!c�A
�'�!as
�\ZS��&ERt��'`�M��Ō\u�e���u$��X�'1­��FK��
D`�n��\/���
�'�����
�23�X�P�퉢<nDh
�'�T����%#h�o}���
�'CpX3�_*f	�G�Dr�`��	�'���E��&�ps 	4aF8z�'�T 1�@e���C��(��d��'��!ِ'w���AdC/$
���
�'0ٚ�,U�;J�p���+Įq�	�'[�Ij�gB��P��	-4�F�	�'8uI�*Ej!i4)�#�r�s	�'�F�	���u��1�J��3����	�'�x<�����X���ã`V
mr	�'�ր���^zj�����!BN,I	�'�d���D�*>��8��ep���'(�r��j�B�i��\�d�,�'*��ف��	�����Ɉr�^���'D��t��=z��(Ej�	{�'  0���/��������h�1K�'�ze���ڭC�NUqV%�>U�X�q�'6j(q��O�z��I�F7N�\��'p	��o�6���
��
)Ht�)B�'@�T6̘	Z��L�E�(���'/�y�O�S��P���8o)����'͢ڂ�c��6�D,pȇ�-LO@�Cg�<,_Jiw������@"OJy�`^L�<��N�:0��²"O�]��m�^�|���`��;@.� @"O��{E"�$rؽ�6�l�\��	�'QhiۗH� �D�`��x��'��iCj�����UdH�tg��S�'�T�1�Q�5j,!�� �:��4A
�'=
�+|0�{�nƇ:�dLh	�'���[����6<ss@	4������ �}��E^|�ص�1EI<z]$%��"O�|cs��,9�0PBX��@"O@���N�4Pj7���*����"O�P��J�!h�j0b�w��\��"O. ��+)��3�
,� ��'����˱W�,��F�%8�+�N1D��A����ػ���*.�=�F�-D�pS��T�g�^�3�K�9��)��>D�hh�i�5|���To�%q`I�$�'D��8��R�o�Cd�go(q���9D�,0��(�y���r젨��2�O��}�\1 �>}g����-�q��q�'�0D��
ŭ�,!�hڂ�O�U#�M/D�|x�h0TlRm�k��v�9��8D�� �Mٸ��1଎1$<VI���4D�6a.}5���roX#* �6M��y�Ȅ���1�A�r�0C�
���yR�U�%!nU	�>pɠ��xr�m�z�9a��v/yHu��'�Z��1�~�T���0uQ����'v�I��6#��Ó$QE�$�:�'�ı,Yp�P#KD�ڀ2�O�b�<���Y�.)!�.�fa$��Wz�<Y�i_@U8��Co�0#T5�q�s�<���_%\L�۳�.9���o�<��V�U�-@`Ɩ�oؾ�z�	�_�<�@�/4	���H�%i��� �
^��0=�a�[t�%����n���A���Xx�(�'�6��4�^�44r��.�.��y2
�'��U��%&db�
�Q5���
�'4��W��K� ��a��9�>��	�'�&��Qd�k��	���?���z�'�<�k�fߪQ�"�+�Ɖ6x���'��i����|�����Є;j�����?1�{t��0���O���a�!2LhU��p�Ĺ���+��	j�� �k���ȓb���j�nm�ƹ1���z6��@����#,��S�!Вw;$���RH�3��#��2�AL��8��%h���V�q�Ѣ���>3����d�rP�6�W.l�����w��88
�'	�{5m�/
j`��!�b^����'[V�x���N�V�1mLUb����';���T�mAa� I'J�J�'��d��NX� �p�� �ÿ/����'�B	3 D̐E@�SQ*��'��|�a�����ٹP�AP	hI�'�$�JF�U#`��,�!��F7f���'���ae�4\�a�
��?w�,��' x��m�+:a��ʲ#V�=��x��'��țFh�/�D�QsNէ2w8���'�8	��C�j{ZB�ŌW�Y�'F�hz�$A=s�d@�r!�3'�pܓ	�'���P`����9�E�W 6&�)a	�'�Ĺ2j&	��2T�*{�l���'nY�A�Ñ9���@c��E9�y�'@$����	'P�"��n�ZI��'X�K�%о~=��a��
l�j�
�'�h��<�Ƭc���e�Ș�'s�]�cg݀�8䡛8P�q��'$,ś2����܀�'Е[��l�'�PDAMPw�i�5"\	Rm.�L>����	ʑCAs�%��6�<���Å�!�D[�U�蕸�Աy�*43A�!�� �P�i�2R�b� !{��0e"O�Պ�&��s��)�#Ȁ �j�'"O�]��E�$i�V`��K00W�1�r"O�I2D�M:y��AH�K�-F|""Ol��h��NI�]���ވT�X�ҕ|��'9�Oq���`T聘U`����	��wb8�g"OT)&k�YǪܑg��>g�q�"Ol�jV��?V�,`���iXSv"O�=C ���1���{�mZ#4e��"OjЁ�!G�F�vh�7l�)j��`"O�E� �T�lA+�&(u"Oވ�އh��Qc�ЈgIsc"O�s���,G�t5��	�>����s"OBQH���:%��p'Ӵ	V
E"O�\rPR�u��Zw֘#<�q(s"O��p�L��bz��A�0��*�"OZ��%�h����#��OY���"OV����>=E�q�5�ƅJE�d@p"O���E��e*N!�"�QK:&��"O^����άu�
c�,�)+�P�"O,��`n�&
w ����"ODB5 ѕQ����*�z��"O  a�@0z"8#�ǟ&Ou�e��"O����'X����D�����"O�i"T��;DHd���V�Xł"OH�Ej��|�������"r��Y��"OZ �U�-L`�АG�5W�l4ɰ"O���

"�`��%;Ԣ�JA"O����!�U��W�ͥ[��|S6"O���Up�Ft�%K �~��eS�"Or����5|&ة���� ���"�"O���fϛ[9�\Aq�ٝG�ȼ��"O,P�$�"�
�cdi���f�qE"O�`�7�O�w���h�*>��"O\�I 
�a�4�� 7o����"O}(���!�Ф�&dR�`��P"O`+5�Ooi�� ����,��c"O�tQgL8��T!�A"&ú�@"Or�SV_&���S��.�p(�"OP2o	t+�zK��M�q�"O��R�N�s# =�aI?(��"O�4���>c�
@�3�ó"��b"O<��+=��тT�����8T"OJH Sf�'Y%nlhSkP+>nE�"O�|1s,�#[���� �ݎu/ Q�"O��a�H��qQ$��h�%;�$4��"O\�:�BE|� ��z�*B"O�iS��ώX1��&A7lT��q"O�P�V/� ��$�� �0�xf"OP �#�i�,���A�du^T"Of��ǋ-M�p���Кp�Z��r"OP1@�DB|>��0*�x�'����(MlH�ˉ�t�J�'��S��oP�y�g #����'��Kg�*\8�xĪи4z�q:�'N.X{�,��lӠ��L[�*Ǭ(Z�'����'ř?@}$���*VDP
�'JҤ)�`�(XP����
PXq	�'���Y�(�\|�cǟ�R�E��''���e�*.�-�ĉ�Jf��A�'�����̢HQ:��$+��/�Q��'u�@�#R�$"  ��P��)��'v9���4�=���u~���'�|�µ��.%��c���v�:X��� �˳�J�E{�]��\�[�*�(4"O6q�� -	�t8Y����&w�� �"O�<��к[!2�¤�#���R�"O*�!�)�\Y�5��8�d�Q5"OʀgO�2�`p�%D�Vy��(�"O)4��ߨ��d�fhmr�"O"�1�*Ծi��B�B@�L�4ݡ�"O�e��� fv��E��&1 :"OT�;���MB(9mI�Z)�݋�"O��J��P�q�l��Vl��.�x["O��{��+1����SeM2t��r�"O���s�
�\� ��G�ů/�$u�5"O��G���i��zPC
�Lfz��""O|�c�K�4���xFIS��vy g"O���m@��v�2FI:H�b�8 "O@R�M<$M̑���̽R�$��"O�X��i�mpWҬ
��C"O|;0Gͺ�LpX�f�BԨ���"OPc�M!O�V��]��	�2"O��z��Qi�АG���Z�L吀"O8e�r��
bU��s��`�"O��C���';)�|�qA�<:Ҡ�V"O�m2���v( ��F�B?��*R"Op�k�l����9$S��h���K�<!��B�/�\qPǩ�2̀�p�Ο|�<�Ƨ��e'Y
�K�& jwgJ^�<�A���Ѐ�!@t�\����n�<�FS;ED� 	�o��ȶ��w�s�<��.� T?Z�q3�ۀh�0���KI�<aVn�"c`��Ň4m�B(B�G�<���m��i��,�2z���'ÚD�<�C푻'��0k$���,[h�<i��@�^R>�k���!<Bb�(Ơ�c�<� ��C�����牠~M��'b�<y3��1G&\1�U��C���d�<1��K�W�e�B��#WP�S�\f�<9�dWo����.ڕC����&�N`�<�p���#�,`��M�J�	%�A^�<��恸Mpݙ'k�4�����DVa�<�) �d��iV�%tIT�)��w�<y!�S�q9<{BLR�)>��d�G�<i�o�34^l�0�#��n�F�2�G}�<y�b�W^rQ��+��C@�~�<Y)��>Ƙ�sh�6Dc�Z@�<9`Ȟ�0��YY���A ����@�<y4L#Z�������x:&�Hw�~�<	U�YO�m������|2OG|�<�f��Ҏ��1�
�AI������v�<!pl�)W_L 1V0^�,�+fN�J�<���[�$� �2C�Q!�]G�<12�&?��0�R��+J���A�<�C�۴pS��I ©�Ь�$��@�<�\7t�d�3��L�\��5U!z�<)����5Ǣ.Y��1B�L^x�<��G�=��(�"��\�YÁ��_�<y0�ҙQq���B�V�>h#�/U�<!�
�������b�$X;FCRS�<�E�͎.�y���gs�L�QG�u�<IU&�4r�bEgfXK4�{�<)EMAĨ})�ǕYf��
�!�z�<�"	]�;eb0��
X��e
�&�y�<� ��;� ��M1����+|�<����]��mzW�D�8�n����|�<!�DN;B����K��Ǹ�I�G�p�<� �,��K��:���C�[]��"OX��ʙ�N�j�ER�WF�$Ф"OzXj.�E'x=��U�`�8�³"O�5�L�- ��ȱ�!�8>�Fu�1"O�@6"��p��j�lY�"O��ʐ�W�+AR�9Z�13�"O>�C��O(b�Vir�$Ün���²"OX�]�-Rd��9�bL�"OzȊƧ��k��������<�C�"O��Ia&��P6x��ѡ�,��"O�(�����e��r�k�N�"�6"O��5&\�S�N�yw������"Oε��C3�ڭ�+ӓuI���"O�}0�P48�pĳ��WA��h�"O�!�_�V<�E@AdZ##	�"Op���&�f4�u��{J�:�"O� VDЛc�Lt9E�%�ft�"OR�0B����8l@Ba�<*���y"O�	�Sb�'�H��G�}�V�Y�"O��C���e��2�XQ��"O�݉���|�B�N� d��"O�Hei;�6i�R� ( ���"Oب�	R�k��P�� �6��"O�<�Pς$U�1��D�[��@)'"O��0��8��Wd��jYC�"Oh p��)'��|��v�1"O��k'�1YR��j�B�2Ѽ��3"O�aZ@nY��Jy�4B�)�X\i�"Oh*�C�)�T��R�F�z-�"O���iP�H�l���t{l�G"ObY��B��h�1���(��&"OХ����*6,�I�c��	.�;�"O��R���E �L0�#�S]�V"OB-⢪�K��yb���!"O�9�Ƒ�ZD��B�!/�R Y�"O�X31��.]ެ���G_.�8�P"O֨
�V�Iva�3�1�"O��@���<SZdP���	?lPؤ"O,�C��'R	��������s�"O�����R�>���C���x�"3"O�I5�((~�+!� �H-d���"O��#'��v��U� �O!Y����"O𜹶�ҘM��p��Z�XFq�$"O�=(��_�$�Z�~+�xR"O�8R�A�#Y�z��u#H��0h�"O�����.�V�H�&h�1U"O�������v-鱀��+�`T+�"Or�ɶ��l��v�	Ԇ��p"Oda�`j[')�"u�ϙuѼ�$"O֔ mϪ�`1sm�7�\l(D�� �A@�~Q�y���V
�i���=D�@��hтN��5��ċ�s�bN'D��Bc��;�����^{\�7�7D��2t��L��H^���]�6"ZC��.;�(�T��	r��A-)� C剃DvPQ���B0(�i)���da!�d�]�8}�rn+@�8�[%!��12z����O�J�� 閼b!�$��6;�!�E��m����C(��e�!�DմL>�e�*K����� 5�!�&?�]����Fz&��1L�3�!��%UH
Q�ǊGuc(����h!�dX����sCٱw@�(���H3/!�D̤4&�Ȓ��@m���"�.�!�� r����V4U�$���'ߏf�^D3�"OBd(�*�>��Yq��oL���"O�1����1���C�Ő�p4�!8�"O9�1!�":�RxCN������"On(�C��S��XB��@޲�9�"O1K!͏+d2�8�-�<RԲ��A"Oy�R�E�0@��m`�)5"O�� �HK�=�ti�D�-> �1��"Ox��c޼SX=x�Qs�t�!"O& ��'��HE��B��";f,��r|Ur�.B�N�K�$ۊ�d���ă���f5�Q8Gd��NŇ���A`�f�@���QjďY�R��ȓ95{b��;h��<��
�XI­��e�xP"\24.��u줩��l&p��D�Ӣ[�&Aζ-�ȓK�MI��Z��p�wF�}����6O� F ےK�B�[&��;;a�t��J�u`  'a�, !�@�"���ȓ?���[�,���T1@�?zn͆�mZ4� ��{ʤ�0�$��c����ȓ'�0�D�X�0P��9|)��S-&���/:�&��pߟ	�v݇�p���2�g{�+���x~d���l-�0k0�ٰw��� �b	9���1V@ �`Ǘ�P�``Bx�Z��1�ԑ��]�x7Xx�V��͆�l��q�U��~e�DBJ8��u��HJ�,!W�s���3�z����?�x��b	z�
y�Ɯ�	�(�o�z�������  Nbx3W(�8<7(q�p���y2�� 5e��f�L�%�
� 5J#�yҧ�	D���q"��SFd9C�� �y��K��DX�'AZ�R%�b@B�yR��
�мR"g �(�$�+���y��V�*����cD�,p:I��J��y�-��x�"�"�� ���ɗL#�yr�K�O}@ �$��I�V��Gƀ����hO�O!
���������beG�����I�<I��'X!�dsMO8bH9JA�m��`y�	V�'X�ӂȌ
j4&8�mʫJ.| ��'��a�ElI�⍱7�R�m<=*,O&e;�O�O�g~��;b{�U
VF��q�J8[ Hف�yRO�.v��M�C(߹z������c�qO��Ɂ/u��v
�+���2��;w��ߟh:��-y���`aiڞM�ݙvJ<��Q����h2|�1H�։HY����7O�	u�bP���w�&=�� �4RB	��e0��m�4�����hԳK �'��T�,�(��h��!��4�\�p��y���qW"O
H����,A�H�s癝$㶸	Z��D{��I�SM�]#`�A�	}���MY/x�az���C�V8H#'��61ff��S�Q�Ԅ�[:�$뱉�p ����\�*"��<�˓$�:H��҅�`گ3�2�J�O2D�+_)�ܰ�5�����@9�"�x?�y�2O)H��	ҎQ��%!&��\ m�kQ��}���`*O�$E��R��h�*��#�>���ɦO?7M�A4ȕ��C�&W:5��!®T�!�X�z�@m�p�T+DPh5�s ��/y!���g2<a����6m���`���!�R�t�� /V�l����(i�!�Ĉ%`�x!JR��>��nŐ-A!�2JN�Hb5AK�h㶠�!#B�R�!�� ��3ks۪����k+ h@u"O��$�pm0�R�S�k'�P�@��\���IN���13$��4��|���q��\��(��w�HY4l��Hh�.�����kf�O�}��n�4y�C�~��C��dւU�ȓI�Х/�5h��0Wk�*�����M��>�z�����zW���q��(������?`�p�0l�$Y�a�C���4����xy�Éi���3˜�I���ēD�^��RFǨ
�b�xPO3k@��1"O�(� b�M�h���
��{s�����<���V�%rJ�%FƐ:�����C�<�f���_��բ���b��r5J�x� ��?�1h��e�NB��I5Ab�	�qI�DX����dæzD�BQ@���&����</!���
�\S���K�vHZ�ϐ�B�!�D^�u�*i����.Ce�)�gh���,5�O�iQ �u`R����-r8�����g�	,��'7jE*V���@⡥�~����'*�`��Ɍ��6�����1B^4�#�"�)�Ԧ����!@;�z�ҍT��y"iU�{�8�C\���#Bm�u��#=E��'���K�B��X%�㖟���'���3īٶ
o�UQCi�\� ����x����%�<Di�Oڦ2\h�/A"�MÌ�����|E�hv&;-J<0wʵ����y��S�,�x�M��5��i��F��~��'�p�'pe+��E
�d��s1�ߓ<<������n��t��l���E.���2a;��a�4b��]��)�*_'�zT�L_��hO����E� <�KSL��]
h����o�铁�>qv�߻kR0u��	����w��_�'�����O-z|(���:G�du���M5����'8���R���:�$��%M�>4@�B����Ǌx�����W鈫|l2đ�#t�<y6��$M�ؽJ���4{¹	�L�l�'sў�']Z��dfש3>0"�[l�Fl��vВ�+��� ��FN�L-��A��:q�G�Kl��w�ˎ"}�x�ȓf��y�)����1+
h"�P�O����]�a!chIJ������B�f��=�Sܧ��D�mv�*G�W{,�b5(��<*!�O�W����O-	���`��\�'��T�m>E���c��-��Üwdht�"?���I/S �EBG >/���� �	5?��$4�S�O�^M:�d[�9tp1���]�&Kd� "O��+���[Lb�@f��wGl����d?|O�M�p�}G�V<,��ทH�V��\�'�05���(3n�XXb�X+A��'�tqr�X,U�j����,!� �G"O�ѦL޼^6��0wA<7�U2r�'�Q�� t)Y�w� k�b_+	��9��<D���vN�	x{dE�V������C<�$ �S�')�~��H�)�̰�C�ԯI����V/l�ٴI��h0&���j`����Fq���]l+���&Y�h܇���?���+������X�Ep�<I#.�-�����j� 0�1��n�'���4§XP1e�K����Rj�,͆�#�pԘ�Mծ ��8A�e�Y��*�Ip���B0v٠&F&��Ć��n�A��c�|���	ik�m��ܰ?����G0��ϸW��0�Nb�<s�@`-1�
6g��t�5+ _�<� �EEٶ4�H�����v��� ��'K��'���,t�S���g����g��#q��B�ɼBA&p��<�x�A&���S-O�rJ�"~�	!�$�ꌜ'=@�qhO�C60B�	��f�2�
���j��Ll�7m<�S��M;CdA,p�`;�-�Ch��@�s�<��_�K�X�KӊM�=�_�7�4�P�aV� �@��d2c04�jB�7\OZc�x� @��)�"m���B�	dR���� D�(�a�L�dW�5U��0t"��� ��D?�(O��ΰYeH�K_�MS"�^]|Zm�"O�Q���Ʀ}r��ְ]alX��Z4�!�DT+� P�%Z?�,Y�ゥg��z��Hc�6�0�ن(��q��b�n���<�O2� � �"TJ}�g�!` `=��M 4�h�v!T�w�^�˅�I>c�͡\�,6�9�|�f%*"ZA�f��	���B+O�"=q0��?G�$�r�Ņ�urWa�l�<��/ʓp7VH@���O�\�`gRq�'�ў�'A1>�)�,̋p��A�ĳ�X�ȓv%d��w)	�A�q��Q,]��A��m�@���'YvI��I�k�\��0["1#�E�/,��#���Php���RS �C7n3i�e[�n�]T��L�>����Y�j	�ikj���
���+��ڞ�� 3IQ�I����e����@B� �zЍ��d]��=�IE([6T��4�PyE�ȓ~�N}+ԯ��&�8yc��B�9�ȓfW�����u:z c�eO '��ȓ'VnѲ��8�nD+A ��Oռ�ȓ�l	��)��B�D�:�#ϢZ��0����h#W��<� ��@LGV�5D}���+M�� I�G\�Bt\����f�C�i���D�2׼A)	]�\ ޴�!"O��u��Q/�貅�_3=���"OF���X�Q��H7S�Չ7"O�%J��G�\���E�Ӷi�1AU"O��Ɂa�[�8��f�(�D�9�"O�L˧I\�K�)H,4����"O�4��E�x�l\��JR0p�\l�v"O: k����z���[�-���0s"O�I	'#��xdH%�0�B<i�X��r"O���"<~o�P���T�1��pF"O(5�F�W[���d�Y�!�,��"Ol���g��y�`�
��Y����;�"OZq� ��r�hx�t&�$2��a &"O�]�ի!��(D'�(?)\Wb�<�AK�(� 4��Ac�p %�La�<�!ǥ9��@�j��8�� @F�a�<��)�%n�$!�
�>;L��;g��v�<�	��wc��f��3S����wcG�<�S3>��@��XLT� D�B�<IV��r?��p��A6���/v�<yS`:c5�!���P�$����o�<)D!31n�ر&�/ˮ�g�PR�<!e�J'tB�9��ܫ	�M+���O�<Va]��5V�N'b=ʝ@$��N�<��շt���:P�8�`} �l��<�g畢G�~�2¨��*M1N�B�<��W/^w�m�f�ƪ"2V���A�<х*�u.f|h��D�]4�A��%�u�<��ʎ8��m7M�!V���0QNr�<15�O�$�3�d�LrXh�2�k�<� p\���j��$Ú�e�HX��"O�)��	yF��GQU����"O܍V�[�
��HWgQ*}hni�I8v�TI���[!��2U�.%��牿SC��r���i����t�޽-w�C�.4��2��J9Y��Qa�/Mz B�ɷX��K�J��_],U��$�G B�:k�X	�L�]��9e�R��C�Ia���e=#�8P9C��3��C�(!!^�p�A��Hy��׬=q�C�Ɏs>(ۑO��\!��H�	fC�!s��!�+ĥ��%�(U�O~C䉪L�&�ð&�.^\����nU8
�,C��Q纑	!kOl#��A@K̀H@B�	�zN��kSo����'%�58)HB��1En	rI۟V8`D��(V�>�tB�	�=lX�@��.�HL�u��"O�U�4�]
*�p��aEV�,9��K�"O�IC��"Q�)S��=`|@7"O��F�B�6t-��d��r��`"O=�vF�^�J��"��V�l��"O\I���K.�})C�X���YV"O~Ȃ�HƦ+p�פ�R�v��"O��CG�w��X8�C����u"O��;���-%�ص��)ֆ8֨e+�"O�a81�]?U2��26H�:6�ʥ��"O���<A�h`Bf�:R�Xir3"O�P��*�fd�d��V����"O����P6P�|q`�`�:���"O�u$�-Ϝ1k�@�b�ƕ�t"O�!�"d5Fzvә6~(�q"O,`s��I% ��|
�.�4}FT�2�"O��b#-�0cᤐV��t8��2"O�I�G�6`�`[�MH�R˗��y�A�s����%�X�E���b��y2��#N�񢄍�Nh��-4�y���@�PL�޲� h#�U��y����eN�����Ը�h�
С�y"��Vu�ԑ����j�xRdB��y��ֹC����󥛟 *�Pa�,�y�Hȳ6Ƣ�X!��-xVD���y2��1*T���  �ɋ��S.�M�$	��l�%<�|8���,H�G��3$��m���p	ح��iP��Y*V�Rxw	�2��C�IR��phE�:>���*P�(T��B.<��A 6?9�O��P"|B l��w�\Ę�� >ҽ���v�<����}��S���%V_��R0�[?�s_�r(���VB~�Ou c��ȁ�C�!Zd{b��G'>X�� )�O8Qacv]jɫ�cɷ��!�1��#'�A�O|�#G��0=Y���$f��`ٝ�J<�Э�I�'�v�x���@~�P	���%j�.E]�y�#e��"���C��D�<�K�h�pdh�G�y:0��&C}���S:�ħO`��fN'ʧ!vq���ɻe;4�QfO��'@Y�ȓ�����D�L�^��$(�,<�$���dHWl�� {�[4��%0�`$�:�E�%D�\�dJ��"H갉̰ug�Q�,!D��{���4���̍�\���c�;D���Ч�:X2�PI��ˬ.�҄�6'+D�P)J��x&Έ�ǎ$1�d+D��yN�f�8���w�@8+��&D�p� Eከ6@�'���h��U��y���z��I'@[�=B�}��'ԫ�yBͳ��� ?����
�yBʆe�lx3`�97���PK�*�y���"�����W#d��@!���y
� ���'e�>d,}���@�ts@"O���e�:s�6��!�֮`�*D"O!����6"�Җ�ߜ�`� �"O(��"i�~U�q��Ҡ,�T	��"O&x�b�EP��)��� fк0"O�!��ɓ>A��,�%a�x@�@�CY� ��@�D�%��|�/�!c���R��'�40��Sj�<	"��	[�yjr�
�(Þ����)��	{U�)+B�]���g�3֘U0�%�׀,� �61*�O�	I"AL��O`\�&�2	*neyBOB�R͐���MZ�%���%�&��ď�&�P�ڂ�N�2��x�]�Tt��k*`��">���e��#+���ħ&XH����8c�}����� _��=i�Ґ.J=�"�׎N��K���'Yd�12�#�:y��h1QF�!i�2��\��s�Ǌ�4X]�-O�f��HK�Pi[���YNj�2�H9D�� Ѫ�a��.�b��O^�F���J;;�5�R��*"t�
�=���'�2�l'V?����'�]����2��';����iͫ�Ő��м}���8�]�8;d�E��R���ި��ci�0Y׌�� �^;!�1g�5_�=�m�.0�S�A#u~T�O�S�h�C�;k�4@qɒ)&����� vP�6�I8(@t.jF���Eh,�W���B��#T;N,�S!�'��Q�Or�`�'C7HEhA�@�ڞfZ�)kL���;x�|{G�*F��sC P z�$�8\)2�.X��؋-O���L�CgZ�LJ�A�p \&{��)�D��Ȩ$_4
�M�w@H���ɾjQ>�qM �^�J0�
6�T ����*��Im���(D����2���`m��oz��Su� r?1 �ޅ�=�V, D٨D;,Od����0m����P�FBt&(�y���@��oj���1!Їa��������ѡ&f��?	V��z��<?.�`���#�Љ�fa �6D4��S4.4y3
�'`\�����6Wĵ�.��^�Q�%��O�}9���L��@ �ř�[`^�����L���TAT���oڀU�����b�#n�!�$ VD��C���#b���1��8<2���.�:6�Z�-�b����'�F�8%��0od^��[��,t��+���ia̮�T��_��A��c�%]�k���<8Μ�1�O,���@�+�0>9�捆)���v�X1\����'Vb�'h�t`��<Ʌ�
Kyj-2��m̓ ��H:�-�C�-S����2�B��$k�>��
��Z�2ӯTM�b���jn��� a��0�F��4��:tr$Yu�C�,
����9N�r���+��L<�� :i���bw��a�<���#ӮN���v��(t���h��Ě�FE�AQ��B#�mxL-|��' �E ���-}ƨ�yD�Ӳ�ez�X_h1CH�h7��d�r¬��*3���퉨'��`%���a���E?[D�Z��ЎT����'(�ݠ���Ĭ�%9$�����TӦ�r!I�A�N�hs�ٰ']X�6i%4�(��/�78 �e�tG)`G�W㜩L�$Q�S@�Jp|�V��8s2ک���49����ı?lt�ȵmĮj�Z�r�nQ���y��/i�P�27.Ђ�F��Ǝ�4���8t�`��!+�m��l�	�I�Ga���O8�E��'O�(z&L2.�5Ad?c]Ly�yBo�bXd1 dg�<�i0���|%*aB� Q*��֓�����" ʝ�`b�%��=!E�ӘI.���c��F�Os�M�jP�7*�tw��0g���IL�'��h���Ҍ�?iEK>+B�r�H5Z�8BB��R�<)�E��Dz�(z5b*mI����^ӟ�b�ǎ�Q/���VDY��=9�Tn���)�zn|- [L�P�FҟA՞��	Ó_	��d��'6��$�VL/?���q��9|i�왦�PS�D)��Y��!�
�FШ���/£;�v�!�NY��ɾ	����u�;$hq���7,�������:*�z���Fthy��!�$͸m\��L[���"��:,�Є�f�Nz�l�eh�Q���벘�t��ē��Z3!۰G7�8�WLM�7���ɵ3zeqăG�BA�%yp�=]ƴy �X�P6h4$ْu�y㣅�2����\��=)�*\�)K�=`TH�~����U�H:S�Qq��'A�����
/R����)��t��@�B�J��ڸQ��i �[���U�S�O\�`C�̵@ؚ9��v�Z0�X�ꦌ�*4���2Of��a�ڠ��b}!�,�,r�����q��!���2'iJ_�v��'&xmh0b�?J/�Y��BI��Q3@�>��/�.�"�6��DI
!^�Uv퀈_���l	?~����0^����G˿�0?��%�,cA�w� s8f�pʚX�d��ss�'��9��ቹe���  �'!�q���s�j�60ʹ�{���!�����ɃV���Q��*t�O���B��5��b0LS�I[r�� �H+7v�Ei�� �21����H��ɣuJ�P�u����끨1 X�n|4�/�"Ƅ4p�H=�g�? $ F���,B�1�1��8�`Q@B�a7 ��R$�k���0k�$ ax��M�Zᦨ�SD�/�رq� [;H���U.�J?�����I��DX�B]"���dጎY��PkeMM� �j�0b�r TkW�ʵ�x�/�^P�I`O%*Y�P.�h������E��Yz��Q��L��vo^�YL��S�+�O+� 2cΑ')+Hx
���=*�0���9F���0�� >$Ԙ��d>uC���s�U����#W�F�s'�6@Bd$��'���%Z���vuH#|z/O�d����_D��2IU���!�Y��b`��K���(`Ie��p����:M4��i���X|��2�i�8P�����
�C�$���-��#�*��Xy SV��$��i�j�HqU�U� 1`��EA�۞�H��d�d��D6?,L�ڳ	"N��  ���YH�x3��65�f���U�Lh�x���'��}�.2�B,ϵ?���{�G[�
C�r�a�.Q��l�3o_?7~�����"1�ru��49���sK~*���`��ɛ2�K�[��d�c'FK�'|�[�j��/�����M�>pj��':p��WB� x(�)H����!։|)�!���0i�* ����@�O��I�9bDl*' �=f��
��G�`;��ɹ�����T�28��Qm�0#?�P���5.�\�Ӥ�X2G!Q�EL94D�"씻H1�+�䑓'\��D�	�-d��}��Ɠ�TAC#�N�#���j6o���PB@�)nd|�Y ����/P��܀@�%4��1��'�u #�LB(LÈ��CJI{����S*A0���/+I��s�U��ecu���%Jt݂�@�9EB�ܶWcBpa"D�/,E��D�՘Oj�����e��B$�T<ܒ�Y���b���a�aٮF�L���z2�ޯHg���p�˜)a�3!��(%U��f��������>��2A�E��.6s�U�-CD��h�'Tp���ڭj�$�O�>������6i#�)(�XL��~�VU��a��o�6�*��(���<���Ssg�C��`#��8Q�'��h3���8P1��`+�
�9T�Lكl�9�R���$y�Y!B�%�=������%��a�����Gy�������N�e�O��T9�kP�p��	���Җ,�`U��'��ᰱ��|�|�e�K�1"a���JJLɇ�!�)�'lD��3N�5F������
�$Y	�']�)B�J�q\�a�T�Z*T��'aR����p�
�it�^!s"O�H����&�s&A)4���%"O&��W�4r�f|�Y?
�-�g"O� k�B#a&���&�t��@"O�y�w.M#@$`�S�O@�lq����"O��-8~> �ĎE�!���Q�"OА� .�zP`m�6����"OНc������XG�E<R�T�Æ"O�l�`�^9}�^�t��	���q�"O�1��'i84Ƀf�X��r�{$"O`� `[?t�n���q�!"O����Y�pUj�	��HY�1��*O0A�$�1{]��N�(��pK�'+x-a�n�cf^��5IU�D �
�'�`IK��R�^�(�05��<-�A[
�'☜�ŁN)1[�5�t�̓+14�J�',�[�[i�,�c�%֥*
�'j��3�U�-i2�4�	�'s��4IN<��A�������	�'l�p�w S$ZA�	��[�$��	�'��r�ֈ����
F�A	�'���Q4�G�}�N�=���)�'Ҋ�(��^�"���@	�'5�P�Dj�lZ����N{��i��'���tZZ�`̄�+�8H��'�>ă���H��a�ֽi:�Q��'�j�t�ƭ0ij��$�h�H�s
�',�r���B�t�D��Y���	�'���������,�a��H(�Ps�'���ê��e����T�
�R�' * ��mJ�$�z�I_x��'N9R3&�
.��̇�N��:�'�L�80�Yz�u���؇A�Jm
�'R	��L��@~(\{B�(.r���'嘍�+5fSV��`fב%V�QQ��� P� �����P*S*?'ڰ�b"Oҩ"vό�d����o��$�F�h"Odzg�S#oG�eq���<Xx�1�"ODLp��=���ѲޏYO,��u"O�yx�$J����� 93hE�"O �#�,DA�P���	�f,�h;�"O�=�p�p>�P����7`*T��"OF��a�\@��!���f쒦"O"�9A%S�1�H����G����2"O,��ԤR� r���F�'Z�nCs"O��(͜�zpܹ҅.���A"O��V�ɘBC|�(��݄|� "OQ�UK��|u�yx"��If"Oh�p�ĥ2�� ;��\�,�<��"O4���!�r��!���E�Ψ��"O(�a�GI�SH���C�E���Z"O�X��	طo`��&#��(%�`a"O��� ��$�b�D�T$�  "O6���L�?��q���v��"O���-�.�����D��xHu�5"O�ps�N���ZģFP��a�T"O��ۦɊ�h�D(�Ѡ��K��9�"ON�"�D:QRf��S�T$R����"O���F�ً�� 0�34�>�P7"O�h�C ���l⡧E��h��"O,���%�2r�#�f����ݙ�"O�ə�i/���H+�4;�t!��"OH��u�Y�N��M:��vT9g"O��A�L�-�\�eȞ{5�`"O��CҫU�<P��Z�K�U%,���"O�!8�M�k8��3��dހ��"O�8�ԡ��`�$U袮��\�]�s"Ox�9"�	�!Tj��Q-�?
FL�q&"O
lr��`�pi[U�358��!*O&�"pAQ4i�X�Z�A]-j��`	�':�UI��%`�+8�Z��'%}�<���G�6 <y�&J�D��%k�y�<yB��< r1F*L
j��� ��l�<��� ��0&��M�I�LQd�<A0.זmbh��{��i�p��b�<�A�L�0�*e���
S�0y���^�<��S�^�x]A5C��X��@��ŌZ�<�`,��Bt*E�x�BP�4�QW�<9�L%c�4����
r���qƢw�<���a�%3ql��cCT-�cq�<6�3H�dEL�M��l����I�<��E�u�6Mʑe	a�24�円i�<yp�����A�S������s�<�N��0��k���^�[��V�<����\M�)RK�L<h��(KJ�<��$����h��'A�F��Q15��B�<�E�͐���D�
(R�ɥ�z�<I�f�55�.��F��>|/���GIZ�<ɡ�݀&��r���0�a[y�<�C �Wd@�RGޒa���`�-v�<�b�&X}�l��eH1Q�ډP�
�Z�<�"I�5{0ib�mT-FL�X�OM]�<y��KĴ�*1�$Y�������|�<���;xI����m��D}�<aw�X�!�*��O�r�v�sV�GG�<�*�$.����H�z<0�q��[|�<���>��%���n\̫E �~�<!�˓�G������KOL����]\�<	�D��yC�`J&��+}dM���u�<� �yR� �0Dlh��	R%6�����"OB(C�HǑTO$5�P��(t��X�"O��#j�5d�܋Re�$~���"O2����iE��h�9��XV"O
��`陎R
#P��!M�~؋4"O�E��٤���j�':u`^ub�"O��A�BB�|g�E@�G,zn͊�"O (A�����8�����R���y�#S�Wv�ra-M�Z5�Xz��E�y�)�d܎�S�AǊUܔUBB�����dU)RyCv))���u��mb�j؋K�H�эX���B�t����A@�H�b���\�O���e��:4�%>c��6ň-77ڤrŮ ${��$�f!?}���I���E}���bިq�d�8ܬ!�%�p��#�@�H�$��'e��ƢI�E�.qY�Ȏmt�oZ�L��%A3�JXZ�C��|���9O|�{�6\ ��B4c���&��Eܓ\�T��rn����A������|2�bY�l<�,+PJA�,7�A��C?��كT�U�!�H������g�rq��`]�����bMCV�r�W�L�}��l	�
/�\�O�G����1���ЇL�� � �"�@�' ���w�|��Ӯ@}4��aA�n1�]s"İwb֯Dd �9�Z�)�,�-O�� f�	n�8� ��D��_y:��w�7�.��[H��N�MQ�|j�f��4�*���l��|t�T�T/}ʟ2Q�S)�ߝ�d%\�v`C�����V��hO,I9�k�Ĝ� �%��#��R�Uj/Jp*��H�kD��OZ���̒4)܈Ä�K��J���;7V���&�ιt5��q� �dSbU��9wĽ��O��(�*O������:F�ƕS�a�¸�����L���)2�za@��
��	9PbQ>�+5K�,t ����j�0Sl� ��-$4��1���ծ�"_��zr#}2��T�s��_0=%Ԫ�CU�:��ɇ~���@ k�TDQ�䳑 �74�&�^�Q�آD�Xz�c�S���8q�
/o{P�Ր>��`5�a.MN�e褍K)w&"��h����m14����*��M!"a�lG�!q����&1��{��[?RC�id��ߑɒ#�5c����C|�ٚ�@$���҃�1{��;���Y� ��N6�&9��|���4��<���
*���Zf�5O����CΨ��'�Y "Ama�Q��ر��@�*�~��ۚe�&���  �Ԣ�C��r�SAńjE���$
h-,@e�Oz�b�2���E�fAyѬ)D���fKNaْ���L� T��z��;�ɑU��`;�֝Ñ>=8W�ݫm�bh��@��;�FxA�6D��h�H7��5�C޽c�hsWk��ef�\���\2��I@��~�n_:P�3�ɗ"���⍆�(O�`��.ߺЈ�|X��s��a�ME�ѩ��'9&�`W�d�^���ɝ	��U�`�M$g�z�g�Z�-gFى ���@&���~��G��+mHɉش_.Rhx��&.D )2e�� �d�ȓ$��d�Ŵ�P�0���ȥ��<LcPP���URi�����]�"���>i˟�QAq��t���	J"\�0��'����DW���q�EnЂ m^�	ȸ9�Y2�Rܡ�m	����O��D��'��s�N��6�jE�Wj�@��B���4 A��]h\��~*D@��K
|���DBl�{ď��L��d j�F�[4�';`E	˖8��Z�cє~�����&Z��D�c��f;�	u�'����0��5�?Y�L*/B\�2�@Ůp2�l�U��J�<Y��A��fK��R��mӰ��ğx2*�m���I�����DH�F�gܓ���f7ax�ZU��,
axr�\�(�D��ԨOvp�0��tDtmY񥃣j�ZH؂��K��37$��H�/�Y��1L'8��N�<�g�U�!�8����T�~-�ɫ�A^�aRc?qa��D6� 8"��Fo�X��<D�|�1�Y� ��9���� v�*v��'��;�+�X�T� ��ab��<�0a�x�n�4p�e��ՙ ؀�q��ð?�7(�l�j�Hď�W܉he�Ov^� �2��G�<diŁ݉U���P�eJpX�0�6)P�B�<�Y�2�l�3�9�H��<��`��K˞�DK�sȒM�4�Sv�uχ�f���sc��I8C�I�B	�	Q�d8M�Z�� �?
��$�A�&ʕ�M��	�׀�K��;g����A��>jK(�#�6u9�C��w�"p@�j�?��)3b=o�`�O�	����5|�J�&>c��2M�>3���ԫկY�	3��5�Ov�"�$�X�? Vl���E�)�j���	�*���h�'Ĕk�Z��� ��j�K��Z,2=��+�!F���T���\�r���4�yRح�f�.�r<�d�ڈ�y2��	r��k��1~�N�BAJ�9��A�a��=�*�)�k��I�?*/������~������h!�$�Ek
$��:��E�E&�`B*Tq�&���~�n
.3s����yR�H!)���Po Z�v��L��y¤ظ=;��ل"�ZF,3�L������N.����Y�6B�D#A9.�j&;D�n�GBH�,� �ĪԚU� I�q>��t��ԩg �r���u~5	�"O�pp�-W�X2ש	�{_v���T���`�8LH���+\�!E6�����P�gdS��O8X�~@j�IȣR#!���R+�,� [2,�JDK�[�n:]Xu"3�!��h�57���6�~�?��ܯ.*��Ř  �ճ��-�O�io��Zu��Ps�[�~���[���/-t`���6�u�G/���0>iqh�tT���K��"f,q���l�'���E�?���k�5=,H�Χ%�<(w(��G�Z<S&+G�|���0GT��C�5$\6�"%�-A����_�	�B��*�fB$�!�"~��e�2CU0}�P8V6DJ��]�<�q%GlvH�;@��")�r�� )�Rx`�F�dӬ�i�EZ-<�H?㟸�WCLb:03�@N����g*;�O������4��O�KK*��7D,F���{G�H�:������"�O���Ɛ�ga��P��A4����	�
j �Af�6���$>m�J�P:�E���^.	2�!��=D���
JT}���ߒ�
I��ߧ��Ɇ6������V��S�O0���t��4v8���A�K0V@i�'�R9���E��pi@V�V8G�=�L>Iv��9E�5�Óa0n K�)�>^�P���L���0��L��2-���d�Ead���ȓuQ
��G�'떍[��Q
Y}��ȓ`NLY��HV�0��w�S�X��̇�o�p�C�o[�q �������ȓ9��j&� 1�b��&h�8M���
qyĜ>=0:xI�i&����ȓ
�r��s�Z�rw�tC0��k3�܆ʓ3"<�6BT�ҒU���ѹ{����;~�b�Sō�\��T�H�_�!�$X?S."MO+D">L+��+9�!�$��PT	1P�  ���@�/5u!��rx��g[#>�$ 	R!���D���� �H�>a �C�>C!�Dg`U�p$_%1Qhy�Я�$\ B�I�Xx��S��`栣�aϳJG�C�I�d�|�@�.�p�5_4@B�ɣ��1�`��sڮ�㝟'$B�ɛDq��cŚ�RӵB��6˴C��mn`Wd,��u���� C�	�]���3�إ��#�eC�	�@P����!a��âc�$h� B䉓�^M�C�
�	k�*�P�B��(0biY��@<[��plM�t�JC�I9D�J�`��� ��I/W���P"O��Z@ȇ`t�\��"��=AL��"O���E۫hVдڲCp�6q�"Oz%b☄<���3�Z @%��"O���g�0�P����T��Eҡ"OT���*(�!��$J1~t*ж"O��i���(_k"�0S�'La�)��"OFqSe�<+���FY#IVMaA"O$�Q�YO�ށ�T��,W:�Q�D"Ovq�]8t!aE3V�J�8�ܑy�!���D�v�R`�̓Q�Fu���εp�!�d�TuG6+��Sg�!�!�D[��(�*%���E��ҥ�:"~!�� l�( ^�� �dm_: h�"Or�s���\�l)�A�N�U��X؀"O�a�nѿ9�J�3)��<���"O��U��<&���ۡ�z�$}�p"O
ድ�Z�qe@-H¥�E����"O�@�g��jI|�0�J@����"O�1��˒�� ��B�;�H���"O써ףя��lx��`-���"O(��S-B	H�p��$j�� +�"Ol	�5�O�pq�C���#�*���"O���"G�r����ro�'E�]��	qBؐ����__��T(]5,���	�K�Q`�� �:����[6u��B�	7\\fE�F �#�����OU6]�B�	����Ѭ
�Ȃ�" (T0w�C䉷BLz�	����pݱA��{6�C�6�X����اwadM�%f��oN��$],Pv�18�<�J��yb"ı9�8'��ӀI��YE�Y{�B#P
��ռ�&�E��5��k>Ek��'��hv(8RV<�Ҫ 4vk�yJ��pp�A>����CaL0s� �
-��ٳת��~r�ًVlY���=V$����!�(�ʠ#�W)�sA�؊	�V���L�rOBux�"\�助�`N�( >��O�J����~�H}9V	˲]��p�W�1*E�ǫ��c��(�%N7�0|�7C��DY��-�����ز~�2��@@n�h����I��)�ᓬ7Y�ܡ0/Ī,�X��&G+Md�r�5O@��b�E�Oip��T`6��ؼ�*���&S�� 	�j����(��h:�A���r��6�O֦��Q�āGO� `f[�Iɜ}jtM��Jp�DIg�q��0|�A��L���3�O_�oٶ�!'�ތɄ��S������rc����+-��Ԥ��C��pC�k����2ˀ�@Lx3�[��CçC�pX���X�O,����٬e3� 2.'�ę,e2���)m�$jB-��fP�X��^S��$�8P��O����%>E%>Ma��f�����M�GfN�j�ʪOr��O½2�*t�DTV>qJ�!u�+ Cψ-���E��OvB��01���"���~�f���._�u�����Hq��.��l�*���%8���h�Zw,��+v�U�P�@L��iM�w۔�P�B�>b��"�Ů1_������a���y�L�._.�d�u%��rMBAE�y�)�;~a^��@,�^9�(P��y�hK�D>�(R�Bh|ag+�yBK�&Y��Z �'}�f�I��F0�yr.��fű���+Y��ypeޒ�yR+^#������OB8�Pi���yBf�]�f���A#����bS��yc��I�0��+R�:Ы���y2�N���Z�C��8�l�REG�y2h�
I0���N��jZ�@�lҘ�y"ޱN������Eʰ�
#�yb��/�q�R@��J�"����y�c�72� X#b�	�&�`����y2jD�/}6$�d��o 2�8�ʉ2�y��K�Q�����a�!e:F����y��c\^�av�҄O�������y���@�5 ����q7@F��yr!ڸbvB9Pt�N&�Ԁ���� �y�a�wT	�*V�q�0��iM�yb�"G��9璋<�b�K��Ȏ�y��$)\��Yn^�b�P87�ٴ�y"ɕ}�6iQ���b��PQ��϶�y�\+�$�iŧ�'V��eJ��N7�y�D=l�bdB��S�^}��(��y�٣��u�5-[ �d[����yBm�[��-X6hJF�*��Q�� �y"��4]y��:��&:ږ谩[�y2��)�Y*b\+4���I@&A<�y�"ǋht�U�w�ܯ:���HP�)�y
� l��A�9L�h\���:M۞5��"OJ���*��3�D��F��
����"OB�A��64�$�*'�$`^�5�"O��HPJ��v�u�` Å���u"OF��
�;������8�X��a"Oh��#��	�� T��8*�yac"O�����O4���Q�&�`Fx�"O\ĘT��d,	��oA6QF4m��"OB�XwkN�#�*525��(Y�"O4q`�QV����ʀ
�V [�"On8� �1`�� pg�-F�P��D"Oh�ԉ��&�ܽ2sf]�Am~쁓"O�,8#�9F��E���9Q �2�"OJI����2t���#�/[I�"%"O�ݐ�!3"e��ƴ;>� �"O2���G  J�`q��Ol%D�Q�"O� ��D%!�0�0��-t@#�"O@�yqA�|�8(�0�ζ%���"O�]��CXX`ꉪ��&&�4��"O�] eQ�_�B<��%	}u l��"Oޕs�&V�zЈ�rŃ2q��C "O�$�g�I�t��F[�`J���"O.}A5 �� b�a���	:I.��2"O�s��P$hT4�2d�=?�Ҡ�@"Ol�j#��,
�i� � *�T9G"O��"��\'*���S7hZ�Vx� �"O8TA�@c6��O}I@��"O�A[T�r�qGb_�3U,�*�"On���4u�� ͼe�Mr4"O����N;k����/�1NA遖"O��k��6� �qǈJT<#�"Oj�84�5c�� z`�O�.�-�U"O5ؔoD>�*�:b!":F�pW"O��µ�H�}�@��ԧy���y�*͔)�ཡ��ܐk�X�F2�ybCԷZ�$��W��tK�9���%�y"��+ott���Bڠn�P����0�y§��k���GƋa�$��7���yr����À#W�v���_��yr�Q�|A�x���K9Q����dG���y�KX�{�@MЁ��Ӭ�y£�`�ȡP�[�
�#S��y�iX�x�~8�EDz�t��f,Z��y��
Cv�9`#k�nV~T��v�<V��b���a��dNP��4�s�<�t!π~�2-���8�@I2�%w�<9�KD�N2ӇiG�3��$Ċw�<Q�@Y� !�f��w�Pq�Fp�<i��X�(�1Ӯ���1>]$���l�܍!R(
�8Z��ӆ�O4.?D)��@d+%��MA�P(&��ƒ�b�"O<PY׭�(l`��fc��>#6�ʴ"O�!���5YS ����nf "OE U��fg
%aLe���"O
� ⓘR���(F�YYK�-��"Oܥ�s�
���8�A�"8xi� "O�x��V�p���{R�X_���2"OZ	�����"���~^<��"OZP�U$�6`�X��� Lbӂ"O�X� E7�� �6덯Z>VY��"OD3����]��K�V|,���"Oy ����CHD)��m�(��JT"O*qڶ�T�LeԨ�L$�
��G"OJ��ti�V?2��$r�b,��"O� :�
+��f���K�.u���"O�l{�`J�L,*����*ot|�"O�`���:褑(v�ְS�q"Oxi�u"�DE����	�o.�̑�"OҀ�d��(q�\p��ȇ�@�0�!"O�T�v*�:Q��$du"O~����İV#>$��͓�r"�8h�"O�E�VL��*g��T7,�z�"O�QhHM*��,���/"0|��"OvLz��W�,���7♴9��"O>�������+?I��LZ��[S�<qZ�Ao0�:�d�7 ˂��gX�<A�	RK�r��5.HZ�dC~�<A�`ҏll����.�1\���0GM`�<a��KFڡJ�,-VJѺebRZ�<yiNr���b���� �RX�0�IZ�<��φ4��� IZ�@W�l3c��|�<!dB��4���g�.
/�e��*�|�<����}e6I3���0JD�	�΍S�<��<<h������!LSdiT�Q�<���EY�<$�\�3� �� �G�<q'ϟ=���L��/w� �$��<���}|��`����D�ZA+g��|�<!F��9����ԏA=
��Tku�<i M�aU�]V/��^	�ЫWo�<ɔ�6VV4CQfę8�\#��S�<q��pk+%U<d��M�.`�~̄�#ڨ�[cl�=~�Ma��Xr6��*�D�Hm�3�A	0��z��i�� ��șSʛ*^4����E.6<�ȓ#v����H˝:¸�@��z��ȓ���Ƞf ��`�jG�J���i�rI���+f:�,�w���stؽ��VeZ�eo�*a ����"P���І�0��h�J\&j#���o 	2�J��ȓpA0Ĳ+�(R��rǃ�[ e�ȓOeX�H��؋G��l�eE��nM��;'~��5W$�Nh����LD�ȓ.Ǥ@	0�N9{�����-I�!�ȓ3����k������Nϋ T4�ȓ�N�V`U)Xm�.P"3��4�ȓ##����$S .��Z@�Ȅȓ8_6�˴��}��ׯ� �8 �ȓ|ɐAx��?L�lmzģ�?����ȓq���#��"[���'�ՔbwB���� ��;�J�Q�@.�܅�)�v4i@!�60w���u��Gk&Ѕȓa2�<�3@K�[�
��	�8J�X��_���F�t/^\�S(B3V�TA�� �&��e�X]�(���������@�4��U�_�~�f�ʅ�P�`ƶ<�ȓ=�����P�H-���dN&j%bA��o�J��Z�!
�ku�%v�l-�ʓ(`\$����E�~ܨV��$Y|�B䉞N�&�$�0xht�v'<lɎB�IV80P!c��v�>()G�;+�C�jD�t���(c�4(Q��SA�C�		+�f��[3�a�wώ)q�C�ɹg�*�
�/_#J$�}CC@��z��C�	�WAɆH�7��a�����B�ɻ'�蹃ηEj>x�5/�%e�ZB��R��W���2d@�T�BB�I�,π������
c����T�	�B�	�e�����R({T������C�)� 0��]�
w�+�B.�-�&"O�"T)Ǻ	X QP�U�;��v"O�iu� �` ��Y�i�|��"O��JA�7X5�rD� `�H8	�"Or,�.<H���pi� .�R"O����B،.�.�+&��H���"O����<�I��-ْ&�,	[�"Oje�ã��x΀\��u�Z9�p"O�����~=1"�#$>&m��"O�y��%) ���j�X'ha��"O �b#B��Fx��ֲl,q�'"O���
N��q�֪j�ܠ"O��B�^+}�m�D'��zٺ�h�"O`]{G��k�>��P&�4�4,��"OfQ�����f{L9��5^yv"O��!DE�Q�ȃ0N�>c
�`1"OV%r��-����06�`	�"O���v��/��uPf�\٤uA'"O�	�#�Bb�s7�e6ޤ��"O�:g V%Gl\1�����e	 "O�����M�Z�\�0p��M$j ��"O.Mq���4��h�Y4`�I�"O���X��x03��c��� "OD� ��&��Ѐ%E�6Ii�"O�(�C���X�@a��c�d�
�"O�D�Fh�Ga!�'!0�H��T"O�1���ŠN�成��=6SX0JP"O�y�E.D�W���(-V=8�W"O�c"A�X4F�xE��b1��B"O�I��ܓwQ~1���*9N�QG"O��c0�:P�(9!Q�� j�X�"O��)�O-.�* �%�C��b���"Oh�
\	:x�D�ׂJ��%�"O
�t
۫BdZ<�bΎ�Fe�5�v"O����	�)�4���nO�dz�ٕ"Ol�W�»A��A�"",a�0��"O,�B�gC� ��A�@�uC���"O�0Y7A^ܡ0��Ĳ%+��{�"O�m1W/^h���	=X�"O�m�3�ҝx�dga=Wȥ��"O8x�� 
  �P   	  �  O  �  �&  X.  �4  �:  7A  zG  �M  T  VZ  �`  �f  m  ]s  �y  ��   `� u�	����Zv)C�'ll\�0Ez+⟈m�o���I�C���DB�l�Ƭ���
��9��؍Qu���%��@��1�7T{�aI��R:���;mx���b�l���k��h4�HH����MC�/ F9[�������Z3��숱�Dp�塢��.��V�⟰�D�/IϊU�e��#�*,�O�5!�w�H��	=n��-�nN<{ߴi�������?����?ɜ'0��
+���C�;�BЃ$������I�G{�@�۴����O��i�z���O��uH/B�:	
pJQ������OJ�'�<�N�����'9}�a�	�<�'m���h�B�+b	���6���BXP
��y"& ,0��)�ź�d���5��i���?��K�: �bOڬ�oC�c�v�B�f�B�\��v�'�B�'f��'�R�'��T>Uλ��u�2nS����#0�ɽ�M���i.�7�Iͦy���M��ih�7�\�9�		h�ܜ�7�BvƢģ�!#���'E^�c���7M�j�P�dR>4:pu�
<�x�����T�����i�"7��9�S�?�9������Q�@B�@�`I�E��T�b�훵�M[�nW,M��l@���*o!�y��GÞ�?я���7��]X$�[�_8NP*�m� hd�O��bBD��GȈtC!�J0}(�;��	ԟ��	W̧[�
�X�͠ ��� �dU;Xb���'�ў"|�A��=Ag�	en�7*`s��Ԑ�?��D,�$ƅ-���T�{�|\���U�,�(�"�I�x�!�X2qk�X� fظS�z�#4�v!��'�,a �08(=�!� d!�:Ws�)�1[(,�ܱ]��)�'}��1���+�Alz�R �yRN����0�ToC�2��P9�/��hOih��k�y�+�6��DY΂9��B�ɔ9�BPZ��*섽p⅓�VøB�	�1�X�����)+n��It`��i{lC�I4��)���U42A;��V��|B�I�J_�4�-��!�
�s��'�:C䉪�ʌ0DN7'<���!Z�3;��D~��"~*��ڥ/;�� �@�B��j�h�yR�\���0-K^,����3�y�	��o+ ѢT�;TH��Q��yM�+��x��NV$�RE�����yB#��G�pI�T�˩	,�rЪ�y��X,M׮��` 9�� k��%��D�=~��|�&�6̡Y���)�$�aNͰ�y2�т�X�����'�N9q`M��yA��F讵#4FF�r6�)�-�y�\�OON)sDi�o"(��fX"�y�۟W��9�s���f���#���<FP�gܛV����R�њh��@�t��X��!��+�O<˓�?���?ad�+ P条V ��Z�tI;��i�<��ዖ,_�I��K�3���
M.��{���X'�2��:5�U�
6����N�)YT�1'���RMɔ�)��|�".ʓY!�x��ߟ�ܴ�?��.��9c�H'�x�Ҥ��n�H��?�	X��J%K�l?���U�s).Me�ȍBT��-�y���hO�)�ß��u傾_ײpq�@����B���O*˓T�t�K���?�(O�9O��ɠ�p�(cO˴J��Z5k����H�����,8�)���C�
��Pr�ח}�<A �<?��^�"|��%��h���-O��eR�%\u~b�6�?Y����'ژO�`���+ΙrL���j�0�*N>Y��0=��ݺ?^�`WHX!&�P��q�' �}�D�[�l�X�G��G�9Q+
����v/	N��Fy���0.;l���Ǫ4?<t�vC��y���9K��Tk����!#C�0�y�ۈ��H�#m���d2�jB�y�!�:3�q�w"[4%���N��y"�ő%h*��֨W�x������K4��xR�	:L6�`�)\� 5���ɷVh��2�' a|"�:?���92	 �	H����AD�E���
�'�P9A�Q�7)`8CACQih�AjK�x2/Q5j@��:k�E���:�,8r��N�BA�L۪0��dڔS�����Ҍ�yb/ç��R�7
&�ICh^���uٛ��|��-c��|��A�R=.��ף�/(?��ȶ�'*�	̟���Ο��b���=Ҿ}���@�K�bM�V�? �	�łGe�X�b��(�����1��_s�) ����B
�t���p��5�d�JL����� R����-����O>�'�'�����q��� RV���T<޵	�'��O����Y�&�ػ��^,<%�Z2m
}�"(�O�q8%�^�*��1�r �q�����'��	HUIsٴ��'����O�U���*YAD34��9����O���P� 6J�"pj�;QF���(&���~�V/z�D5��ѪU_��I��V������l�f��b�A%n� ]�ѩѶF��?i9�m���R�,@�sW�u"E�2?ٕ(�����|�O�b�&'Ȝ�ۀ�� ��sr��&6�!��B/e�&��Q%R`��y�ș�\�џ�a��)�-;�\b��.�~�2�]}��듏�$�}�����O<���O����yR�Ӏvʒh�����Z�e��
�5P��)�
�Y ����������1%���U!6;@t`�eؒjx]�1(�Ml�����-D��gU���c>%�S@Z�*���]8z�ēv*�x�f��,>bjmӆ�DUb�0��8�<��7�L��g�]_|L� %gI%}�F�s*Oz�=���䞨�J��Ė����g!��#N��Ϧ��	şx��4�?��'�?)+�,<X�(��X�b�K.�ja�E���A�n�$�O����O��Ş2������F=HG�x{��ʟ*���dO���T���"np|�R$��~*џ��q
�|��z�Ď6G�~���K�~>$	�k��72��`o��)�#S?%�P���%`VʡG�(yS���1�Y�68��(��'���'d�O6#|¶`)Y.z`�F�n�@k��|�<�ӧЧ^Nf58ԫ�Ta�L����w�I��M�����šo�n�%?�@�8
}��6*AA�)�O"˓�?���?	d�u�����Ix5L�CU�p`(�УB�f����ƇL?:ﾜ��I�9/De�q��"� (�1m��6=6L�!/ST� ��t�W n��("ˏ��u�剆o��d�O�E
ݑ��O�T���"DJ�ef&Q%����V���9@������@�H��,�O4-���n���y�L_C� ySSLڣ*F��Ĥ<YQ�N�k��֕�Y>E���JB	!�*��� ��P�&$��ȟ�j��8����HKxx�-3S6��O"ȱr 4+���X��H��D���S#<�d�	ƐM��x���N�3(M���S$@�c�f�0��~z�BF���3#�O��lZ�,��o�O-��Qw$��,��:5b!M>��KF��'(�L��;�!�-h��a6`A�\��}��F&����=3F �q�h@�L�b6,\[V���f�2����~�6�����(O�`p �ϝ��;S���1l]��"OZ�4"�#[����fβ?S�՘�"O�0X`kZ��%���E�`��Pf"O!�PH�
TL�9�C�^� f�ɀ�"O^s��/ ���`�!M�(@"OR��c�]��S���(�
���Y��"��1�O�=y K�y��5�G�T$lq�s"O�9%Q�&(Z�`���B�<YQD"O�B1J�2a@��"��%���za"O��L�gɶ�����!oH�"Oh�j$�Z�5#%�ޏ������'Dz�'�����5t��O�M�VP��'��88cOAe�F}�f#�Y鮄�'JPC#K��p����`��'���Ї90�l:�&^'X�긒�')�y(�eE�������#�H��'� �SA�eג����!�$1�����wQ?�� �1[�f�!7���](. ��9D�Tx���&.}�I�`՗g����wn:D����Mzf����R/p�8��l:D�<" �F�y���#(����04D��)t@�����.e9��i3�2D�0�%�?Ʋ���OU�3�h��t
�Op���)�c�0�����}b�c�e5k�"D�|ؗH�i��
A��AX�!E 5D�lx�`Jr&�i�"���*���`7D�@P�ς����-T"�&=S�+5D�l��Aˢp����(ԆF�C7�2D��EՊM��!��]%2t*��<�k�h8��IլҩAI��#4/ܦso.T�B"D�� ��0�%]�fݞ!S�m�0�U3"Oh�Q�f�Tf>�s�w���"O45C;,��I�䄨q����v"O���M���a�[�&��mrք���>�!kt?G�2����!��D���A�<1�m8(k����g�x	�GE}�<y�nB�����C�
  �����|�<�1 �L|\5�8�$T�b�O�<eGv�h�8&J��^\����]�y��T��ą��(ׄA�dᖒ�hOX�S�rg �)���)K�̭��	3H��C�o�,��6FQ�w���0p핧 ��C�,�ŉ@�ؑ3��0�� �C�	�cd���ǂ"X����A��i�*C䉱�fE��bH �͹�F�J.C�g�B�SsO�6�B�s���1#����K�J�"~
����n��9i���2 �$�J�fF
�y��CAphjE������L,1��B��
�f0�% D�2 ܝ�B� 1��B�ɥ���
2&����aFC�'<��C�ɛ.Ҥ=���YPӐ�B�nW�C䉻FE��Ц��I�R�K�N7-x.ʓ1c���� a+����J:^�\��$MX�E�0C�I�-�ᗢ�;�LU �)4�,C�I�窭��2 �|(�@#��M�C�I�I�ޅhM� ,PXC��&Y�C�I�anX���6t��c���-B\���dA�=��D&0fЕ"JF#���ɡ�U*4�!�dΛ*H�Ej����9z�]'�Py"%݂;$�\0J�W��)c4D�yr-�'z-����i�%OW�s`��y�عR��8�^	LBXК��y2+��:9��DK�0v���hO�11��S~b��L������� Y�C䉢?�v( 4�tQ��V�Կ"�C�I&Q���eԠ,��$ƒnb�B�I�7�؝����?���Wc.z�B䉂Q�"=����G#|�r��1f��C�I��P��aΧbOz�c�N������2��"~BACY�0�ia4a�Td���(�y2#�&Y�lhA)�,�F�8w ���yb�9W�𝂒J�z��ѓ�I�'�y2�Щ�����陬p�1vc9�yҎX1��X�H�d�D4�DB��y�HU6�4�2Ǭ@�V��ɐՉ�-��$�}V�|BHڄ �2!��/�UV�%#�g�y��	�Щ���ƆF�΀(�̺�y��}����B�t�6�yFH�,�6x��>����"��7�P�c&�^S2��ȓ3;�鱣i�G��Q�-Ӕ_�q��	+s����=��Y�@����1�㓮'W~C�	:R���g�޳F��l��B�B�I�h\v�!�(7u�P�����C�ɤdG��zE��~q�$H�-Te�C�I�X�B��Ck�&&�zѠ`?ղC�I1;�࢕�Z<3�dY*�kɕl+B�=�#�M�O�H�ѷ%	~F���Đ�&�b�'$%�M8^��\��K�qZ	�'�V����$�����|��'3>U���">�$�H״�|!��'���1g׮F¸��E������'br d_����`S��=%�I���x��Ex��Ɂ�2�D�C�@ZX�
fD�O۶B�I�kG`l���3ZfN໒�_2��B�)� d����S�6n�:e	��<��"O<d�� Z=���P����<c�"O�xR��D���"�$Ԡ�{�"On�����ČqRU�ΰ`�(u_���1�*�OP���2��A�7���Uj�Ģ�"Oܝ�w%F���%kS
K`�ӂ"O�ɠGȑ Du����.U�r4�4"O�tG@H4:q�E���0�fT�"Od �iA��!T�@	S���@S�'��'n�����B�Z?�A����:�1!�'���E�����i#~i���'rP�{`�$����!�:bĪ�yr�>�Ku��*,e3�EM)�y2^�6/�Ɋ"�[�M �l�����y�i%cx܁�YY�ٚ�N���hO�!��=Cy.�9$G�%�\����#{�C�	�P�1�C@�s+j�)�)��~�C�I�u/d�:f�|{,�H.�<{�lC�I�m�P��cZ���AFF0~C�ɑ�fͫ#�;@R�8��'�BBC�	�,��d�!P�Vͪ� �  h�$]�0��"~����x,4%��̺@�l�S@a)�yb��KY@���$���7���ykɳ\3��!V��sW��aI
��ybI� �q�d�_fy����ę/�yr��#K�LIA�@�I��� ȵ�y��^� � vJJ9<���*S��8��d�V�|r�3]ʐ�Z���B��8�!L-�Py�o^�����.� ;����KMd�<���p �hZ� hu�CΓ`�<�1���������� �[�<q�%N�i�`�)��'}��X�ɛnx���&���ë�}����&FE�A
�Xه6D�죐a��x�f�X  ��B)2���h4D�����M��dCN��(�%�0D���B	Cd�D�ΗJ(���+D�hyF��? ��2����Pe(D�t�P	S/0=�:���p�
����$�l�ԩE�����u��}��$D�?pE�ǃ���y��K=k?l0��C��@��I��ŝ�y&G�[^�0�[�K��yZ�ú�y�^�E�)1�B�N�����f0�y�� 
2��S�%=�J�OU��y����'M
��&����T���e֕�?�%KP�����l:�͚	7��ea`�U�?1΀A@&3D�̺�Ϛ�EJ0�#�"��Gd����=D��;�"S�A/���5I(f*D�w� D��{u��=&��`jS��>�@G�>D�ku㟵\���/8Q�T�{�-/D��z�A�}i�=y@�Y,T��x[UB�<9�R8��3�
_�Tx��<8Z���A*D�D��gf��1r&��-%x$�Ab%D�ܲà�0'���۵��-��Cu""D��r��R � w�����e�%�3D�P�P^9��q��:1��#l.�Ox�b��O�d�u�ʮ4������dT
�cD"O^�b'!M�;�&x9� #N�[D"O��B&J˛ �~�B��RL,a[ "O6���� 0���9��?U@<		"O�d+��F�H^�����F�w9l\��"Oܤ���_�J�,9YJ�9�"��hO�E���>Mlk�Ђh̖����6��C䉏a��  .ñP�tM�e�Ê�C�	M���#K8�|�I�_6B�)� xxB砍Pi]��ʅ�]Ԑ��P"O8�8��݌*+=����Tsx��"O�5�D"�=l޽���
<Ir�2 �'�\!���	J	�P���J3V��T0�dN�nB��ȓ^�v�`�O�^x�$��7ZM�1�ȓQN���H����lݷ|�2��;�eT��1H�M���0��,��?K#�-ܻ)���v V,	>؄�o|"e�tf7&�:�q�*DNRP�'#f��i%isc��&|FE����.�� ��c�h�)���yGt�b.=+͊���M��!k� �4Z� 4��bȏ�a��|�HP���B�x=2��AmOi����� b�e9u"�1hB �Y�fK
&-����l���	���Zc��
j�������jB�	9R��Z��2���A���q��C�		-���s6�Ar�� �Ι�\��C䉕E3�e����n� P)Ѓû3$�C�IBn�I�GP;�m�ej߱
HC�ɸHʦ0B�c@ ]�Y��� �B�=���MM�O) ���ٓ,�z�kV[cж���'v�����/�5(F�ӄb��'A �3ƄB~��� ��b�ub�'�
}a$�	SV0�����5[�~-�
�'JpAI����@i�S�)J
�'��](R�ّLU�XefQ�QL@x�]:b�Fx���H5i�h�1˕�$^��c+j�.C�	�6�LE ���0���t�6B�	nz��LW����aeD�G�^C�ɨ=�p�JT.ѤT� ȑE��LC䉜Li�,AǇ߾HQ�Ha4×"j|C�[96�T��;*�4Bq�L�h��I�����f~b�ϖ*\��4}2��+�-@a�O,%�J|�.I7_������<�3g#Red�I 8"��s�4H�d
]7o���]"��$o�E\��D|b�P�[�b���iۑ�<��Ў˫�Х:C�9OølqW�0�x��B�M0�}Fyr��'�?����O�6��U[-�D�a�b��x� ,O���$C\�d �ċ�6W���Z��8f�}�o�<����Z	|���@#N��s�m�Jy�!���'2�[��'3b�U���	rM�rX�ōQ�G�(����0�AI�|��Óby���F�$B���<�Q䘟- ؙ"���yb��./*Ry�a���Pϲ$9RD����rRd�A�'3
�����yr���J�,b����|Xi��� ����$E� l��!�cU�n3��e	��!�\�z"��VC2L���挷e�ўx؈�)�N9�ݓQ�7\R�H��J�H�l���<�D���?1��?A����ԟ��P"/On˄��@�?E3�\��,��<6M� m�ȓ���{�V�'��' ���3�:���p���-aR�&�$�ܡsk�
x�kU'�2��i�/g, �L��@�!]Mu~̡�( ]�V�8u�>?�s�Qҟd�Iq�'���K��:4Te�'"�����H�8!�D\#%Ux�Iv��;�b�ѰN�>��j8��|����ĒB2�tQbJ�3�,p&M�e%���r&�O���O�d�<�|ZFc�p2H�7HK	�4��� �R<�OW�i�����/��8��WՊ�RD'	㜀�r��9~@���O���3�@��`���2lBI��!ʓL����*�P�8bϚ%AUJ���āymN���D�'����	��l�� �w<�%#&�&D���ȋ }"� ���S�Z^�=�-�<Yt�i��d�%��eI0�����0\$� ��=oޕ�ȓ.,n��G�	�-\��D���*܄ȓ	���CAPXń��@T�w8��ȓ	(B��pLA 28�5��-�b܄���P��(܋f`�ha�o�O���<>&���t��G(a�b*]b��S��XDxJ?=�&ϖ�p]s댔'@lQq�4D�X�����\b��W iQ�hX3/5D�LcB�q�䥹UB��f�����A/D�� ����Aգ,1��{q΃�Yg�-S"OV��7N0P=N�e� [L�9"O]i#���h��j�d�]A��z�h*�O�}��TWr�H��HDx	CJ��ȓL�~�
f&W2/�d1f��{�
A�ȓ1F�\$#�K+� �]�n�4(��@h����p��Q�\E����T���@� 'pTdIA��|�<̅ȓ6�(��7��t顡2O��}�I�5����$��!�!�!U�R����F!�D@9r�Y{�Z,-�Y�C.!�ϯE�>��a/L��U*�Ƙ!�dM�&LdA[fn���1I�1�!��i��#Q.~he�7�_	m�!�Ĉ� �D܁E�_+u�Č��-ef!��D>	渕�-@-k۲ �!�ѮIV!�$@�.y����:��2Q�G*Y�!��
 �D�c�E�6,�z�4�P�!�D�?�^9P���p&�i!�Ъd��bs �� S��'L���d��e�)�',`\�AǥTq�Ҝ���I�e�'��~�S#vT��$�v��A�c���'�ƞx"�{̧s�D�`ꛁA�������&���'����<&�Jҧ�9On���e�� �tfӁwǼ�ZǢ�Y�b��\�l�O^�%>�[���4ۥ
��{�eh6��=P�+��D5��<��HP�3�*1�tA��&�J�.��!�i�O�)�O�8�4�>Y�Q?�S�CQ�p����,E��R��Ol�Ő>�Ä^I�O�́`��*K|�I�i�/^��YJ��'Q��JK�,�K��q6�=}��s�d���h��w�zy��蕕ɐ� dY�ػ�a(}��,�z1T9J	�:1vHFcΕ�F����O&��A�>��y���䑶"�=�D�[�H��+J�N׬Y� b�<1��n~rM�n�OӘM���߳Fv����LO�3[����Y(�	�`{��S��'h����'Ų�B�h��,rP��*������i ���d�Uڔ���"�
� �H�C�
�!��K0e��`e�� w���}�۴��<���s�̕��AM4U��@��4)���6��wy�ӥ�Da��	�q���B�� '1^C�	�E2L8�L9�����ZllB�	�t�"�h���'*��I���0"�B�	�d��e1V�R:_�T2ug+3��C䉮s|��@�9.P��kE�U��C��`p�t�AJ�"lR@<����#3��B�	����z4��m~B���k\3�C��p��y��h@�,Y����	L��B�	�u3��Q��Rf&-P M��B�I�Jrū�
�YS(��h�(#Q�B�ITH���$W��z�d?HK�B�ɪ
���cw)��.��a�A�B�dJ�B�IA����D�R������u�R��@����r%�E	?�>0�D�>���ڑ�U8�a�J;�L���c�i�I�|���#aɡ2���Yuf��̼ L!(eN�K���_s>ɡ!O�ʀ!��cR�jr�L3D�e��1`��`+uH���1I��!���:�@�����Y�bO>1���6�Z��[�Q�(�tfY�<1�m�����F�G"\�hQ� J�S�<��:��B�m���V�k'�QP�<	LE�m�<�c�o�,b��C�Ie�<iɅ����;2G�
h(C4o�l�<�D/�LhУn�Q��j�eC^�<it&��Y+�@r�!L
A'��Rr	Zu�<a���j���F[*p%Z��R�I�<�(�Z�*0�pjW1����R�n�<�߇hb�ᣥ	�����cm�<��LO5r�P9�1b�9Q_ Ⱥr�Os�<A��5w��d(�4Kj�;�L$T������:n�(٢U�s �8�	7D�� �t�K�)�P���Z�t6����"O�ur� D�<��\�fN@�;�B��"O[t��x�j	p*^�<��m��"O�PCw�4\~%ɲ�V�u�Dqi'"O
�ɑ;�r�i���o��t�w"O����E�j���y'Icy(� �'i��i'�ܪb�T@�bCL�]n�}��'��� �H��L8�c�D�D�ztr�'�j�C��I8f�hI�Rʉ/q<� ��'x�񒢑�F�n���i�,��'��ɐ�ϣ��`��E֝[���a�'-H��@%M�J�#҇�a `��'-�,�F$�.6Բ�qe��NAJ�'ݐ��獏_Rրr��*��'Up��K/���bѮ��@v���'�R!��S&pڔ�
"ed��k�'��� �Y 3��l����+u��mXL#�B��ɢ���r���ȓu�H;����e� ��U�����,&,�l�&�
�r���ȓ#}�@c��*],�e���!� ��8H�;u�e-0f�0j��q��_��I�7����T)�݆ȓxW�( m��8�`ՊQ&*(����ȓ�i���7d�`L+X+x�:���ES!�t�1!Э���L�L620��	+<��&[3T�,i�%�.
�耇ȓ`���A�5�"��ر?��ȓ`}�tjāј?�����O�Sz�5�ȓl���v��p����U�A����ȓU�d�j ���T,ȝѧ�P
��9�ȓz��%LԹJ�d9�W�0B��ȓm�A�O�&�qrqK]���0��R)j�A����|~�5*���(��dp�U�9>�L�Yd�ޠf��Y��aQ!��L7N,�R��63���*ܘaz���4(��씫K~��ȓ -!���g���ӡj�9mP��.�)*lՀ^z�L�1�F
:#�͆ȓJ�r�z�FԯJ,��@�IJb@��	�ݸ�n�|-� !@%�)3$T]�ȓz3��1�l��� �hO)jp�ȓ"\]������F h􉉧Rhzɇ�06L���M�>��M)!A?Q@�U��/=�{1�ۇR	�)���h���1�'��1i�=�t��D�.c*8]��'l!P�5T�H:d������B�'7Y
�+S8 �Ҡ��@OA.���'�j�z�$�$f��z�R} �|�
�'pTX��ש6`��"�[�v H�	�'���a��\�ծU�f�P9k�5	�''�)�q���E.�����5%��	�'<H1㒯%m���5�Fל�P	�'�|JC��z|�9��&����]�	�'��Ia !�}�T��
:4��'q�tH��Y�,DCeÉ�/cR4P�'������/L�y����(�RI�'��L�S�[fh�X�nD�6R���'��;�R�&��QR�۪�����'�@��B,j�H!χ7���@�'���	��^\�	q���TB�'���D�O�m� =!i�]�����'W|��f�T���	&�S_>��'H8��!��!<�@��v�YUڥ���� F=��HO�Y�f�X"�"Oܜ1rf�$/��Њ��PD��< �"OLhQ�@�$%�Q� ����%"O�!fk�h�T
�+U�y��"O�*RƆ�c�}���U��QÔ"O�Bł�,
��2˘H���ba"O�*�lV��FR/Q�bq#R"Or��׈[�!}��B`�Sc� "OţG��NPJ�d��}� l�d"O,�f�Wy�~ ��Ɩf��=��"O�E�
���ER�N�X�"O�U�S�^1W���th$o4�"O�8��k��VED����6Mđ�"O.�3F�ޤu:�ꁴ.K�Q#$"O�c�\���k��^�T�a�"OH�s�O�h�9�&��80�b�"O��:IS#K�����$O�\�x)"O� XT���4�\(B�S�9��T��"OԴrp&�<v�Lp��Ŀ����"O�m��
�;FKniRD��u%�8��"O���ׄ��?P��R'F�35 ���"O�� `g���B� �ƒ%i$��"O�|�.�+9�S�g��`q�Yj�"O,12k�t`Z<а��)a�e�A"O�	�!ǎ9K����,
�Ɛ!�"O���	������C",���Q5"O��`m�0;�֩��	W��.hڱ"O���E�ʍ�҇��H��,0"O�4k��$,��L�`�休v"O؝I��V������# jv�&"Ol���UL��)gG	�EQJ�A�"Op���U}��Ɣ�9>�Ӏ"OF�*�O�%1��1��oO�x����"OVԘ��>��8fo�P�� "Oh�0"��f�=�$! �F 	�"O��ia
:�������>1@�.�yB�G�,M����� P�@�
�yb	��'��!sU��K(�`TDP�yFG4�D�SE@�I'xa���R#�yR�	*B���1�Ń7P�$�y�_�e�h1!&��T}�t�N5�y���1}��g�Ʈ��𢡠�6�y��ߟn��s����ː��"�y�B�5��HWl�	�HљA��y�͌6q�x��O��@q0h��y⠐4�(:gŊ�q�Ask�4�yr�(D͊���IǍ,���+�y�(��"*]k�LQ[.�+t�� �ybN��[����6F�B��񁳢S'�y"$W~�6���ā!jp��K��yB�nk^�
O\)Z��(X�%0�ybI�%Y�*Yj�$�PF|��N=�y�GV%�eb�m؄<�ƭ�2�C��y��( ��9�a :F��;��Q�yR��kW@��	��`W�(r�$S��y"��)PrU3���\� T�w���yB�H;~��)U�B ��&���y"�ԫS�EgC�6:��m��'Q��yr�����1��&�H�J�y"� O���e!�8q4s㭉��yr:�8��S&��| ���)�yr�*�x�B��{�ѱ�DU��y�$"b���h�˭9�npP�dح�y���K�xB���1xz�)R����y
� �x��ZGC�X�%�4<DT�"O(P#FeQ���
��6E 2"O�1'&?3Z�; jR,tA���"O���	ӽ^����L�J�"OP!nB���q�X���q!�"O
�+WhV?iz�:��B�u$0a"O6]@ǥ; Խ�� ���03D"O��`��ݷ-�|S�V:�,a�"O����ȋqN���m��4�pc%"OHd�įMD�"�@�A 0R!{P"O�9�P��5*�0�bA�;*R��"O��ѣ�>>dΰҁj23ޕ�"O��8��z�<|�&�M�F�x��"OHe���B�\���4bL�wm|�y"O*J�,hl2�� ��L�HJ�"O�`��ޏ~�D8��ІU���#�"O��G�˳m(���O�A|���"O����hʥ}ޤ@�ǂ�u\�!`�"O~E�'�Ҝh�FԊ���"Or�Sf��$�P�%C�p�.���"O�ڷ�]�5�X���6Y����"O�ՙWA�Ga��GcK�`���#�"O$�G��Q�~�`�g����=!�Ig�q�eN�3��{4J�j!�CF�
����pɠ�H��C!�dS�^Ӝ�qoN�kp-��&��!�2w9�	��D�3.��+GV�(�!�K�=�P�9'F�.8%xJER�P�!��	�T(F!�>!�����7�!�d�	-`Q����P�l֭���!��Ҳ	�Xhk�V�1��`��L�tF!�X�x�8aC@�v�&�`��v]!��ǃA+r<�D��|�r}���-?n!�	$���6E5U�F9���l�!�D.L���z�Bx:�!�#N��!�$�O�a�`
? ��@��-�o�!�[6��,��Z�J�S���D�!�d��!�8�Y�_� ��,k�!��	ԁ��c�Q����P	�!�d��X>!���4_<���c� H�!�$A�5g���� �^���}V!���O/���Ȁ}�R�PbD�<K!�$ ;T:
9:��V1xv�1��� MI!�$K+9|j�RӉ5<E,�r��!�$�*9��M���^� +J��Q�*R�!�dé&>(\�%� �DkQD�
�!�ĕ�[d젉c��+;���t�K�Y�!��	��CA�,���c��L�!�dS<�l��M�f ��dBт>�!�HL8��T%җUA���Ȍ�U�!�D�z��͈��]�p���֧5�!��Z��$pJ����ysV�R�	,v�!��0ވH���e��E���O�y�!��J���Rv�=^nd�#�at!���0�X���m�6�%b��D�!�(Z�]�'ǃ�l���u씸a�!��N\`ȕ�:r�,a@�
�qO� K��,L�pc�K�\�P��d�|K\]K (@Qǌ�AJ�+�JM��y2!T�sL<�r@�u�ꬡWI�5�y"�F@8�ta�ncLEPGL��y��^`4�r+�m��Rw��=�y���ZD$��Ȍ�yj����y�!�/@4�⇘u�=����'�y�m�I%	k�j�@���8�%ź�y
� �iق�Y�~���� Ď#J�i�"O�b��݇0r�u���0=4<��"O���@DI���L�C���rd�"O��q��11����(4O 8�Q"OZR/��gј���� dM`� "OƀH�E�+.�M����#�%�"O�23�[�q]Th(QV-t����"O��`�ֶQ�%�sl�#i���p�"OB)�B@E)ټ9�5#E�d�콛�"O�}cPfG��$9���m[� 4"Oʠ�sK��i3��>JR���"O���bC�d!zǯڰ]�f�6"O�a�2G�iHt	Do�R-t�h�"O@�V��>����RNe�yX�cQ�<y$�9b�)i��<3�L%�IFx�<ApiM�4�,4��[1][<)�u@Y�<q��@�%ߘ�)��t�x���z�<�2F�"��H `D�Oظ��QÎ`�<1f���aҶ�Z�-�X� ���ZG�<�B+
:V{84�D!U����*�@�<Yh
����ؗ�܊)����#W_�<���F"D���R,�ԙ�$��X�<�vhN� �����TT8����ZX�<����g~<(Z�l�45P�QS�YV�<��â��]�re��e%��.!�d��KD�4�bj��Z!V�@u�B� !�d�M2�ya�ȇ'52�<`�͡0n!��
�H+�(����H��!�
��CP!�D�=4����,U�b�IJ8X�!���GlЊ��1m*��Ab�~�!�Dn��� ���dO��'�!�d��t�|��ĔwnR���	�[�!򤆜Y��9�2�՞X����a�̤]B!���;7���!��+J.D1@!V&�!�D��]���0�@L���ai�o!��irF��!�2U�^�!`�5!�dO�|Ǆ�����/b��;uO�"y!�$M�0�b5�eӐ5�
Ip���\!�d�;,1.�����c�~�{v��(]�!�ɘw�\%�"�D0�f`�q��9�!�[�Xwt�÷� �y�:E����|\!��d8��BU,�?x��8cY�V!�$�i/xL��ȋ�)�Y F#�!�á7��Ԋ��"��a�gV�|!��=��xY��Fm1J`3����!�}nF)H�S8`uHP���;P<!�$�~�~�#C��-��a��%ܣ;�!�R�F��_	:��ۄN�/,!�ZjZ\s�m֦toha"�J��25!�$��T0���'p�R��(��%!�d�+h!�P  @\��>q8b���!�$Ũ?F8`6�#a�dფA�=7!�$�0]�ͣ�I��Z�d�A * !��0j�2���H0X����>3!���8�h��)�'B�@�&���p=!��T
;� I����	T��ZV��?!�V3������ژ��a����!�䜷l�|k�M�(�4l��_�$�!��c�$�r�^-����&�|�!򤀣sN
p��@<~�,�B��U
%�!�D��pߠ���q�p�C�Y*!��j$���C���`��+,�!���	��d�@⌅�.,�m�7�!��"y�T���'9�D�����QL!�� L� w��!�j����'����"O�P�
�l ���AF�@���	G"O؉s�bW�;�nLh�+�>�Ёx�"O	�rF�^2��aŉ*�d�"O�(r1ᘩ�$Tz�kSF��)e"O��S���Y��#��a�r �W"O���D^�9��pc��b쮽�"O"�� ��w��q��>����^�<!Aȍ�`�s$��09@����A�<	p�Q�:"0����iR�Y8�X�<ق����Պf�T�b{�X��j�<G�U` ��4㍤&�*]4@Ue�<��ރ,_j��uf� %������_`�<A�ᑙ8�~�H��׀~R��4ȇy�<a�C'Eha�@�Ӟ%���cE�q�<��!����ǖ2c�	�`��M�<�+�?'.�
ӄ����|7aM�<��ꂳRy��(N+U����o�N�<���vM8��Q�/5���� �D�<ѐٚd�9.X�D ��d�<Q��W'�d���'%�U�QLXY�<���i���ѡ�U�9�4 �NS�<�  �uT�O�@��Ӗ�FR�<��Ss�&���L�*�+���F�<q�IG
1��H8��:
.���2�BD�<��*L$@�D��L��~0ք��BE�<���� 9e�ysTK�6n�H�2.�_�<Yc)^<�h��I�_�$��]_�<���[7t����ЂE�~�$#W@�C�<)�/�'2-:�(��1h�H���X�<��J�+��,p�BBH/ĕ@��^@�<!�bґ"Pe9���.6��ug�[�<�q'g�Rг�	�z��5�7�Qb�<��%1�6�  �L�7�d��C�_�<���ͺS���,W�c�6��5�]~�<q��P&7Ē�+%��7z���̄|�<��+1�/��]X��C��Xw�<��'U�.c�5"u�æh����q�<a�E�f��9��.kx��bF�<�͝4{4�m� C�djٚulM_�<aG�\&j4A#�/��a�@]�<!WN�<�c�*դ�F��T[�<��&)I��Q1�T�F^�Y�4�(T�t�w��#�$�Y�&ˋM ֝�M>D�Ģ�㊟F9D<+��1Dx�Q�V�<D���i��9f��� �*#U�U���:D�x�'MVd�9����FE&�C�I�=��Er3�8�$��D�:>S�C䉝@Ȃ7��9{�y0��%0L�C�ɃaytS�K���0s%� bj�B�"[K��z��Ȣ,��8BT����B�I�6ŉ�芜F���j��}�|C�	8���ѧ��>��Af�x��C䉂Acvx9᠊�u�x��.9 <�B�	�r.�y81IA�n;8���:�B�?
KHIR��.?��(��`�-^�C�	�TJ�8ra/ ��![B�'�C�ɞ+�\xJ�@�:��]�S�B�:}`B�	�tC2����C�1�g�O1q��B�I2��X��."t��ɁC�5~z(B䉈7�԰��<*e�}�e��/4�^C�	�H�D����(�=�s�M�?ӎB䉼t����K��Z�hP��^�4�JB�3G�2��ABˮ3�.� BÞ�XjC�)� ��x��=0N�� љ\KP�q�"O�qU�?9"$� �טkD��"Oz}��m�C������_75k"�t"O���V�.DV��B�:OD�C�"O����ƙq4�,2�##�y�""O��aR0FJ�BM�S�X��"O`a�tN]S���CC޾M�*a�2"O6�"Q>mJ���B�X�
i�t"O|٪��E�s��u�d�</�)
u"Oz	X1JG<n0B,�!�؃�Fi�"O���n��3X"��,H�����"O,H�P�l[~�#e,�6 ��ę�"O��K��k�>��&eо`����"O�J��_B����
	-�rQ "O.$¤J�Kz�]��NQl�&��g"Op�c��"8�\(S�	&�:���"O�=��S��EA��.��c"O�%
()S��m��lvܻ"O<�*��~_�Ũ�ㆲ'�!�"O�xh�H1v�h ����$*�"O�<2���=��C ���"���"O慐�8KNt�'o���"OB|
�,�%�&�臍�_���S"O�} R�h�p(��б9"OJ!:�.SW�<0 I%C�����"O�� r��E@p�Ȓ�!�0��D"Ol8��V�t�@�(��$�N�!d"O�r�%
�\��ٗh3_�,��"O� Jd8��k�_^�Lt "Oj��$��oM�X��F$~Y$�"ȎY�t^�{�+�=/UvP��"O�=Ap�!6�v h$�NWX��0"OR�V!��=�f���W�DɆ�PS�*��B��ڇG����B��Y"S.��_���Y�$T!�*��ȓ6���Q&�a���T���ȓAx 5�6��>!4tiI�
L6ʹ��l���*��8
��I���0^>�$�ȓAv�� ϖ��4aal��Fp�ȓn}��Ʃ�iS
5�.�6�݄�`�`�E�c�f�`,܃�6<�ȓ�:���
\!`r��9mx���=@�7�Q!'6���l ���ȓJ�!1��]pxH�#�/M`�ȓX���Rk؅����ԁ��_��Ȅȓ_�Pu�E��Q��i���,��ȓ	����fL�^�ZH����
#�ȓU��㎎�QH%�e��2�l����eC��~��qm����1�Qh�<��i޾*� sF�ݬR\�]��Mf�<�"kG�L�:��w#�&A�rE��j�d�<1���4x��!p�ԉP�z��'��<I�g��?��X`�ёPwF�D@��<a�BИL�P`�CܭD�D����{�<��A
5u=4�����P�P���r�<4���{5$��ʺ�(E�AK�<YƜZ@�����r�>���ǂK�<�2h����0�P.L��%pb(^a�<q�cɺdQȠ�၂k�L�r��B�<��֬\�ʉ��(x��QG��C�<#��Y���q(ʘj!�4��J�!�l�g�)l̓uᗟcF|%�Q�o�n.H؃d����x�
B��B�01���
,垈H���?5�C�I�4ȡ��G�k���;Ƌ\�@�C�)� |�ʇ.d�M�Rm�o@2�p"OpչG��%0���M6;���2"O2�Q� �-���<KK�D�F"OR8	��R�%H�$���ܝ-)~X��"O��pO��CV�s��q�@ɗ--D��p%E�'���z�O^��|+^~!�$�K(UZ��&��EHW.
1!�DRE2���O�C�>sfA$!�ā)2��X�A�!þ �8!�DJ� 1�%���U�í[�m�!�DFc�q�J��*[��@�k�&=!�$C����At/LNC���e�U34!�D.h�x�I�I�I$�{�N�R !�$��'�JA�b��"���#�u�!�D_�G�L�j�� �'i�"\#Rj!�ğ�}i����0����P`�=$_!�\�G�|�XT,� x��C�%p�B�	*]Fɚu*�>�"��_fB䉗0�x4B$,��Wi�}�r@@9HB��qP��F��S	B����?U 0B��L�����F�@�+@�jN^C����`�Hؔi`�0"���#tn8C�	�=@�r�L_b">��ț�{�0C�I�L�@d�D+{W��e��B�I�J�r9 E�߳R2\�2�֛Z�B�
T��5��*�&r�)�`&X%ZG�B�I#R,xz��,UK�գm��B䉌V���/m��]��G];J�f�x�"O0�YB��b`�}ʖ��x�V�PS"O8d�Q���$f�l÷e��-S�"O��أ�7Mj:t�V�Mg*x5"OR���7mT������ti^\�&"O�l:bޛV]š�.C�ke�
"O�H�T�G� �~���LO�=T��#�"O�mR�@���~��Vf
:�: "Op���L�>0��g���a9$��"O��	t/�cWLى�Z�(�ĸ"O��I��Q�C�ȱ��ˈ?�lH�"O.��D�ph����
�J1�"O�(�v�?\�) ず�]Z���"O i�b�'n	�1���6O��x"Ot�a��J�+��`Jq+�0�,�"Od���ʖ��lQ�&d�
 �d١s"OҝЧ���P��"Ԛt{2Y	A"O���5&�3h>P82��bf�e"O�Eˡ$�46ATk�ꖱ]�e�"O�pS��';`���A�]*��#"OB�r��*H��<3�E�+L��"W"O�=�A�4���bLM��QB"O���+.r�e!rP�$"O~���� �LT�ELR�yL0���"O�(�� 8�|�CDK�A"�˃"O���Ѫ�s۪u�wHT�'0� �"O�YH׬Y#}I!��G -0����&"O��(��-�\p�ְd�<� `"O��/
1� �LPCB!F"O0L�ҨJ�B �	P��Cq��"O�Ag(;v'���ό_��<�`"O����?_M��D+s�H,�"O��m̰6�4<K$�K<����7"O*��V�p�PCR�9�6�H�"O:����ϝl�\t� �4���@V"O�����t�ؔ��^�:A"O`�QI�-�ؤq��k��l"5"O� �dQ6I��pdXъ������:�"OB���͑`��3	��(v�&"O��jM�LX�X�G�S�2����1"O�Ʌ��P�0��r
R5"Lr�{u"O��I��+L��ii
�H�Y�w"O���X�}�٫ �S (y�*O
x��Ƃ�F���[C
P��U:	�' 4ep���]�Q��PӨ�K�'��phw�˕o��Ѱ�Dʬ�
�'<H��LH�!q���R�V�4%�)�
�'��MyqH�:���լ�?7�c�'�8����
���uV=,!�ub�'u���rc�V���F�ѨMv�K�'τU%�٩kj�;��0E���	�'Z4�4 �w�0����)����'���z�HH�2 e�o슠�$9D���A��g � V%�-s��D��I,D�r��ۺ4�P���	a����@�$D�D#�9\�R0r!)V�:�ؙm5D��X���G�ai`��m�=I�g4D���N�dBB�O�}8ڵ���0D��*��:Z݂��Gځ9	/D��DF/1����ˊB �}ɀ�*D��HE��!AL��A)��^(���v�(D���2,�;@�ȡ�� |I	"�'D����*��{x�Ɂ��ͻf+^�kt�#D�4��	ߞ��h�)Ͳ1>M4� D�貃�Z��T��X�t��KA�v�<�D/�Ek��ړ�B�y@.�K���~�<ҥ��W�D�Tf�y]l���Y`�<iԌE�-%�K��Ҳ9�.���+N^�<IĊ��%."4����+c �`��]�<y/6%�H���@*w����X�<�w���N�\Ai!�ʪ�x�ҧjDQ�<�fd�?k�@3h�C]h����d�<y񁈠'�\�3���eP�A�d�`�<9��®X��p[���/%x�I��[�<At$���B��خ^�4d�q�Y~�<qGM�kVL�M(P����+�!�DI�/�$<��ᖯD��1�R˕��!�䈛5�&H�F��#��Dp��D��!�DD�r��#��~,����<�!�D��Y�T�9��V���r��5�!��G�2e�U�*��<]��b��P�N�!���>�ąkÀ�9oA�p�5�A$~!�D,P��ܸ�;,R0���^u!�
�;_^e����_m:�P䌉,�!�d4Xؠ����Yu���Ńa�!򄕪g`.]YT*�)
fN}I�Ȉ2^2!�dV��Y�bK�_eN![���D0!��W6Nh蹘al+MƜ볋�P!��o�pi�l4d���=j!�ė"7аچ�Y2B(@W�`��T��'5$p	��#�t�B����X>BD��'ܦ��.*n�*d�Q��D_0���'N`% vкJS�`�P�6.]+�'�p�ID�'0�~��AO�|*�p��'UKr�_!eN13��ƺ@�\4��'�P�H	Eg\	� ��28�t`�'�p5Z��M���@o]�F��'r�5��A'�։�Ѝ\�Upl8��'���3")s�Y
�+�A�J�;�'���b���M�$��7D>�5��'Z��"D	/E� ��qݭe�.�BO>�	�S�? �	 	G,�0�f�G.Iv�"Oh�V*U�*>���&K�\	`���"Or`5�U�v���Q��8��"Ox)���ݪ�6�j(R,/Ĥ��"O�����)��L�! ��1"O�(ac'H�!A��[�i=J"�Hr"O~�9�"����j�H�-|��TsP"OJ���Ь6� ����,,��9B"O���g�Y��d���8kB�#�"O�	a��^(�,}*�E��"C"O6��Wϕe�H��ٙR}HZE"O�1:�i�5�p�{s��s� 4"O
X�3��}Q���
�d
�"O ��1��=� �B<4�P�"O�X�g�\�v�i�ʶo�S�"O �rU.�1�M��+e���q"O� ��P!f�蹳fʇ�XX���"O<���A�(�x�቟�-"�a³"O�� �J،U�&XK��t�"OX�(V���$���)�<sT��"O���
�aX� 釥D�
Y�=�"O�(�UHr�ޘ���Ļ}Cν�u"O~����D���8���\�B���"O��8�D�$q��X�5À�8B�h%"O�AQF��!���UrHD*O�3'I�a�v|[@��8g�$�	�'���k��@�l��Ȅ�ף{�4X	�'8�c'�U0En��7ɒ�0	��'�b#ᚘ{�2L� R8'/~us�']-oI�a(Ԁӄ� S1R5;�'�����h͂W�ι��R�J�|T�'�\l�J�2�P�{+V��e�
�'��D�/��{��urcI<Q;� �
�'BLh��0����C'�Sǒ0��'
���!#�St��C[�P�H�'�t)���Q%[}<qS��Vw�M��'q�lZUbN�c��,�03F;����'��$S�GM�iZ������	�'Vڀ�L)*2<[f�b���'������ӗ�L�F(�~�^���'�X�c�e��P:��˖Clz���'���(a�͟��I�s�C�N6U��'� ��"�2Y�D�b��dʘr�'�"���� =^�'��w���'�И24��<,��٩ѩm��`�'TTL1	��,#�g��� ��'sh$��Y�|��M�Ё�>��\�
�'��Ȧ"2,�tI�D�0}|���	�'��R"G�?��CAK�v�r((
�'��H���
�)'���B
�Xk(M�	�'#��;�56�8��0NN ���'�@�t*��H,�	����%L���'4F8�и%f]J�!�s}tP(	�'�" Bר� B%����]vz���'D��"^�a#|5���R`D\ �'W�0��G!1X,�c"�U�)�
�'��d�O�8zR���D�� F��D�	�'T���l�$(s�B�K�!66@<J�'��2C�����IP�R66�Zh�'���c����nt�W:��i�'V4P�O��0$��XT.�5s���'�����j�m����roά`-���
�'_�#r%ĖOa� �bh��X�}�	�'<	�VD8�6R�X=N������� ���'�/����I��!�.	k�"O�!Ȃ���Re�]+F阭g{X	 S"O�I��Gȸ9i@�2(_A���"O��`u�
bx�Ċ�&U�]vZij�"ONl;���R)��I7�֓	Ƹ9�"Op|A !��:­ɅË<�����"OZ X�*F�s�]q$���K���"O�-�CC��4�h}R�쎯 ��	��"O�᠒��N�Xؘ@�y�<hp"O`��A�X�7��a#�+u�r�j6"O<�z�O�C�B��E┪t��aB"O��H�.<]���p���;U.v�Rs"O&�Q��Ց� PbdE,,G���"O04�bB�{l`)C�,��"O�|�
��G��ᦈ�+l1��+�"OTD�х�5n�pЊ�G^}���z�"O�m��)�
 Z$J��@�]@n��t"O��fhU)2�֬$�S:DRa"O�Sb�(E�*icD;|�"(+"O|x��?S�n�S8���r"O�aS�/�����',J�`"O2��ń1e��ja)��?J<��"O���qC�9In��W)ZzA�g"O�t��UPkZ$�Ƨ� <M���"O|�$��;�D��M��lE�M�"O$�0E�
�􋅥Ǆ>&��(4"O�9� ���
4 �
'"O�%)qL73e�D��GĶ2�j�"O,����j���=I�Z��2*O��{#l(�rx@�&ݶV^@	2
�'}x�s���'����g��#�v5A�'gS`hђ0H	v��p±����Py�KU0ev��R'�f\���G�^�<Ag�
9;�a���\�h�b�o�<�D� T����2�h�X�ҧ�j�<��%J$x/Լ��� �	���Ll�<9 �C�T0D��P<���3��c�<���J;%�
T�P�T:~�T����z�<!,BvCR�� H[��xӋ�`�<	b"W+Fm6-��E�q�L4�V�\�<YD(ŕU�:!C�H�ü���*VY�<9���2a���c4&#nV ��@�T�<�v씙
����+�!J��`D�R�<ٵ�T�"�&_N�d81bYN�<A"��	2���:/�U�$�rh�F�<�ѫ\$�֩�e\�_�`�T��Z�<�BnA�llx)qQf �qP�؉ V�<a�OF�p��T���^�]���A�x�<Y�J
6RFXQ#*����1�E�p�<����}���ԲS�r5��T�<�7)�	X��FEJXT�����H�<�uCI&�p����R�Q�3��n�<YUJ@/w8�A`���0��.Pv�<�W�ΩA�ƥ�Ef_(Nx	�kJt�<�G�T�;��)D��"C��%�VB�p�<!�B�':�Y�!���(dS[t�<��F+7��8�����I���r*	q�<��ZTz�ɂ��N�	)p��g�C�<�b��f���sri�5��<��&��<qg"�$f����,r�$��E!~�<�
��!#^�6@�'qA,��N�x�<Iƭ����D�$FD�X�Mze�p�<y@ǌ|�c���y�����(Gp�<Q�m
>����%������C�P�<� 婰�P4dPqʔ�lӄ(7"O�Y�TꟌ������/<W��x�"OHA ��;j��]��"OM��#p"O��c�	�*T|8���#,rq�"O
`KgEP��AD�ԡ~��q�"O���Ã�#_��L�)�6� �r�"O��EY�\�5I bZ78KL!a"O08�!��DKy�����e���"O�h��EO�@
�� �R)4�[�"O
���ҋ2(����<>�����"O.Y#����W�,�1��3��:�"O�1B�i�$a4gց##m.�y��(3��$e�D,jpuc�%���y��+�b �$ҙs��%��B3�y��Ȋ
��I�@ޟ�D���"Q�y�iK=s�Ht˅�
t�"i�yR�ٮG�4���e͵]p�ѣ���y��X�^t�$D/s�,�s��ڶ�y�oD�p2���mr<�ūre��y"�F�C��]�� q-fI���(�yҩ��j��t&ЀeN�)��8�y��^�/$�H�q*ƛ@���	$�y��W 0B�ZQ H��
��y���k�P��c��Z�F�
�y�FB*#½���ȨqH��D3�yBeO�p��ܑ�aȐ`����2,�:�y�B"0�
�a��íe蠄��䊩�yB��d��p�;\a��� �7�y���T����ǆ����X���ٺ�y����'��W	���hpR�GZ��yr卋R��#W(��*�i����y�
� 
C�W(B��I�!Y�u:�X�ȓB例��もq�8�"L�gK�9��>l�h�3�	�IS�(�K��S,xC�I��8�@N�0����hA
�JB�6P|h����� r㬀&wXC䉦#������X�>t@B� �k�8C�	+]B
��$C]��VLc��H�Z*C�	�k�6�go-�B sT@�v C�	�G7�踕C� 5ΝQ�K
�=�B�	�D�B�8���?N�lӃD*�^B�IڦIE!xzX$��MZ�>"B䉌&2�iC���}�1qZ 6��C��N����(u�#��73W�B�ɮ]���F��S��d�9pDnB䉽
�t�ˁCؤ��Ī0�Տ85�C�ɠ$��������>��L��d�d��C��$SS��bl�8'*`�s*@,G�C�I�x0�Ӄ�Z�R�.��0b�Z��B�	#8)yk@��	�"|e#�Q;fB�	u#6Q׀��^8s�lQ�bB��"&���b	W
L�ۀ�O9J=<B�I�+��4��bQ������4��B�I�#%�<qr�*�(k�EK�Y�B�	�L3zHA�Ȭ�"���*Šb��B�ɞ1�.�kR`R�Dh*9ڄ䃸i!�B�I$#�`A������;�K�%&,=��0g�`Z����8F؍���X�"��ȓ
oȐ�vZ�4^�����vdL���T���I�1O^(��@Б52�B��?S�L�3 B�+?~�8S *F--y�B�Ɏ.��"#�f ��*����i��B�9d�r�0<�t�'`� @C�	#0����L�bܘ,@[�PC�)� n@Kw���&��s�E4?��ZF"O��P��,q�`�8O?5�r�Bf"O����G�E�vz�D�n% �"O�ƭ�UD�ؓ��,u���"O�i���';��hr�O̡$��t��"O�u0�� 4��j"�^�F�z�"O�{��-�Lr.�`:, g"O� ��Ƃ= ?��ۆ���K:�A��"OQ굤4�8]�D�œ ^�A�"O�����,�܁��M5M�:�D"O��I��L1a{�y@��_ �<���"O$	ka(�>�P�TL��%"OĤ*���pa�8��K�_���"O6)��}�A�mC�d�$"Oԭ�RFS�I)���c��?��D��"Odh8�)֟1X��7bN|���R�"O�i`�C��@�"XB����H�y"�WJ��E���uX~Q�eNΧ�yRI�-9���ʂk��U��)��d�yҋAYL��b0(���L�1���;�y��9z��SM�x��{T�\;�yb ��I�x�Y࣋7P�#tj�yl�8�������n̢l�?�y�%c#@(x���5����3��.�y����i��ߺ<�4�h��U��y��H��J�4>�([��؁�yb��1_$��R��E-�U�Q���yb��,#ZуV+�N��t�!���yr��H�*��®�4S\��ab.�y2,C~��D
OHκPx��!�y��+�z���
+B'�]Q��y���ap�,0��ߋb��`2�bћ�ybH/W ���QS��!�E�� �y� ̻ HqKR�A�L7�;	�y���m�����CH��dk��y��B�"���kB8R���1EOе�y��K+y�`�a6)-KOdy�i���y���|V2q�6
ISԩ�tϞ��y"-_�MREbBFn����0�y�X�V�uҀf�l����[��y��I�5PD��4��_K�s�N��y�+� ���ȶ���CL4�c5����y�p�VQ�GN̠�`�;YB�I�;�FD�ՏԠ=��-yr�X�@C�I]rH�y�m]X�����%� �0C�	&k�0��5��
�e�05YC��(z�$H��>w鄑J0N@8pb.B�	#e"<���Y9Zs~	
&�K&w��C�I)X�ܬqW�]0�H��+H(>��C�IK�D�9��3nZ�R�Ɠ4�bC�	?�(�D�P�$9�1ˏ:L�C�=\�mB��� @��UY#"��&3�B�	%1����FjJ�c����5*�B�I�3&����/7U��Bf�p��B��(n��Y�MC��"�Ή.n��B�	�#,�4 C����|s��Ӕ5�C�ɧ\�.���ĝ1>��Ԋq�ޒP�C�ɺ0�l����<���+�I��m��B�In�B}�4��i�r-Z��\$�B��b��rGG*yP�YtG�Wc�C�	-{
�D�d� "�-� f+D��p���S0�l�b���`�գ'D�`���Du2A��I[��p�A%D�����!y��	�i��V�$4��#D�� ����ݦ]�\<+�Rwk�x""O4Xy�$ܶ#��i�W��85XY@�"O�$�vf�"�JE �/\ ش�1"O��K�OH/����4m �>z����"O��B0�U =JѸѭP��v����I��s5�ĲCr�&�'P�t[?�F*��,��+��[N6mC�� �f�����?���<?̌�5J)ۺ�׭Է\)6��  m>� �h�H�� �$\��2=k#�3ғZ��Ph7@�~4��`шO��vh�FsD�|�©:u��(*E-��[yF��MQ����O�&>io��72R�蠈P�k�\�;�
�!��(H�������B�ęox�h0����	��ɝ}�R����!�۴�M���:4�nP�l݂U؍s��GP?���F1d㛶�'�X>Yc�oUş����=�CͭE�>l[#H�1o�N��b��sb`˧�G���9�un��z�p䅠?��OS�t�Ƅ��E_�3�ر�m�#�� p�i�=
� Q>~M��B.��Rt��$H��\c� �D���f,�`���O9��4a� ��ƟDq�4�?���i��eaȒ6�̣#"N��e[�']��	V�X�D�A2韁Sf�	����FO��Dy�h�Νld�'�uG��/
�$hV'�_/���p���Ծ���O����%��w'V�d�O��$�O�į��?1�4F����!D�:� 4iR�B #��*����gt�8��N���b$�4F��ԡS�'� �ڵ�I�<��ˑm�ϒ�dV�G�][Ub�fD��ȇ��=' f��OD0k�+�	�nt��v��:LR�JdM"w������b5����3ԛF��q�,O����>s���^��|�Qi��J��M�e[l�'Say��m�l0󏈅u�i��ꂱ|0ntm��M;J>�����)O9晐mu|�v!@�`hPdÕ*����P�Oj�d�O��X�pux��O��D��D�AYx9vՋ�
(�F}�c��$K6$�������K���O����ԙ(��Q�1AF�Q�廰��b\IΘ�*z�h%��%8��y�a�L�']b�:��MK!D�f ���Ι�mH��0�"R�dR6��O�˓�?��*��|+6,O% d 1C�ȿzl{S�>Y������@T��;��\)P��\�UO��u��ā �b�nVy���1d��ퟴ�Ix�$'�wI���㫁�~�䨊D��pr ȐD�O �d�O�a� �*,44����x��Sl!N��S�rn*`
�c��'����7 �#=	��"5����3��q� 3� �f	�<Jpi� �( �PB �˰b���۵��O�nZ��ħ�M;3�G�R��T���\��)Cfl]�3�2���5�Ȭ=e����K�+��0@��n��|2Gc�ao�u.Ý�n��4JR�$^����!���R�(��M[���?a)��*S��O��d`��Ԓ��U�b��LJ��ԔSPpyr�G����P�k�9F<��%Z�T{0�pڟ$˧�*]c[N\��9x��@�ĝK����ٴ*n<��T�$d(��DJf���+���56BǢ9#D���bI9s�tAD%	 �MK$g�ɟL8�49I���'<?7�E'�D�0 ��D���S�B&U$���Oޢ=9�}2k�W<~azu�J�
@*���E��(O��n�$�M�M>�Qjb>�P��Wsc$�+n��hŢ�1j����=9��<   ��   �  ?  �  r  �)  �4  �?  �J  �U  �a  �l  x  +�  �  C�  �  e�  ��  �  F�  ��  �  ��  ��  C�  ��  ��  f�  ��  #�  c�  ��  W 7	 � � ! Z' �. �7 .> pD �J �P gQ  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+!��6*\�c�<4�d5h��'�B�'���'	�'/�'�B�'���U�W9��m��Ʊz�0�b��'���'�2�'��'�b�'�r�'���k��.Kªa��͎ 5���Ha�' ��'���'�R�'���'���'����
F	�>]�&ΏfEP$�b�'�b�'��'�B�'�B�'O��'�$��zm@|XpjC�6�D�'��'���'v��'�'��'�"1�)ֽⲵpa����j5�'���'���'t"�'��'��'�%؇�Δ*��� A�B4%
0��'�R�'��'o"�'�"�'/"�'�f}�b���Xs���]��X��'iR�'���'���'��'W"�'g�=��'��"��	�Jw���'���'j"���d�'5r�'}��'��u�1� (iL�\r6e �t|:\���'�'H��'J��'ZR�'vr�':h(uC�=��)��G-P�����'��'u��'}��'���'u�'�;+�'HhufUmzn��`�'���'|��'���'��'p��'�J���R�h�����*|h�p�'���'��'���'h2�h�x��O��"�q�R��t�T�)����G$�|y�'��)�3?	��iOTt�#�Zyf��B�º�1x�I��D�O㟀�'��a_4oS֔�v'ۉH ~�w��6z\b�'�@D8U�i&���|�f�O��t��$�U�X?y��+��p�j��<!�����7�'u�xR�QV�HWΕu.˅�i�@�Èy��	�O�N]GL�c'`��XΠ0�$E[��T���O��s}��D�U�	ܛf7O�|�1FA%4�P,�׌}�R�*�9O��?��	%��|���
�X앨sB}�F`]<TQ�<���d:�$�⦕��'���E"��.\��#r�b)�����<!��?ќ'��I�X]l���#O  Zt%P璸;1�?��l޶rw`t�|��L�Obta�IцM{�T��I�$��0+[ܬ�,Oʓ�?E��']�zd�;a���%J�Y<��I�'��6-����ϟT�?ͧT䜼�!��fl}j�G%}�"}��?���?��a֠�M��O(�"�z�j�.oQ�4b�(uH�+&)P��ON��|���?���?a�����hW�(�&1���2�.My�e�O`��s[�0��A�̟��r"�~�tRj�%��Ԓ"�IRy��'�r�|���#ގx�n���ңl	b��P$E9|
"�iD��")J�8�ð�(&��'��9�"Z�A�: ��A�'h��t�p�'|��'����S�@A�4?crp`���uۑ���Xa��V��͓�?��rS�,��ڟ���?;J&̨Q(����i(&	ػ��<��LΦm�'�4c����?=�}���bP���AH'2��
����͓�?����?Q���?����O�X�Se�	���w�Q�͂ C��'P��'&�7�ݼZ	�i�Od��$��.��$G^~K� h��БJ��Ob���O�)�)`�7-2?�;f�D�S0=�}B#bS254�BroԾ�?��9��<I��?���?��`�d4�ꡅ��mF�UpԃF��?�����ݦ��5)�ğ������O�p4A��_�\B:�0DV��"4��O@ʓ�?q���S����/��SbHR�
#�=��N�\��I�"�Ӟ�$}z�O���?��L$�D�$,�$#ā�!`aV�@b�_����O��OZ��ɳ<I'�i�����$�?�<���-Ձ6�A�c^3nM�I���?�.O���@+��s��VX���`C�V����O(�J�jӶ��`�b#����O]}�˙�(6:l聎!F��L:�'��I�����П$�	ʟd�	u�D*)?���`R(��zy�І����6-1M�D�O���5�	�O�4�
p1A�G�uV�Hp�
ib��h���O��d4��I��.S�7-~����M�O���1����a�������ۘso�D>��<ͧ�?!e7B����� 1t����?���?Q���d要s�l@��䟄�Q�)Vā�I�O���� 
y����O��.�����Mjd"�J)#X�W���PG�3,{��"��)�S�,r�IƟb2&K�3��ߦnu�l����X����T�	Ο,G��'���p6�)_�aT)�t(��'��7�D���d�O.�0�i�ыf.�r��0%ٲ.-�8��le���I��	�Gn̐o�l~"�k��Z�?�A3‖a,ܸ
�:05���A�@!"�'1�i>]�Iܟ(�	ݟ`��6h���ȑ'�t.��)A�ʎ`�lt�'XD7C$Vp�D�ON� �9O�a��ŘAx����(ڎk��a�<)���?!K>�|2��L�QFH�4�YK��0��I���eąZ~2`D-�&��		5��'��I3Ϛ}sS�ۤP�LJBLT`�49�����	����i>i�'�6M�|���O�_x>�Q.g�(����J_�$�O�L�'8��'pB�?�X�"T=/�8��5���!h�!S��i^���F��첢�O�q�l�� :�6�D��:Pb`�0QwD|Y�3OL�$�O0���O�D�O�?�C(�?Ŗ���Ȁ&g�@�Pg����Iٟ8#�4X�r�/O�$9��'{���SW!��?��aç��O$�O����O�I�;T/$6%?1�	"2`T�ժ^>CP�0�vd�-L�&IHca��&�����T�'���'�&x�G�ӡZ�x��� ���'�P�DIشf�$�#��?����� �BxH��n�~�	�/�#|o�Iny�'�B�|ʟ@���D�9��L�Z��U��%T[T�{q�|����|������<���ƞ6��q�C���١Qh����I۟�	Οb>9�'�b6��4�B9b��ӓS�~�	큞6_a�Ь�O8��O�Ȕ'��iB�
��a���S�VC����W���'����f�id�i�	����?��Y�t�Uh��dR,�1��n� @�W�t���'b�'��'�2�'��<�(�h�+�,(U��VH�N�,]��4L�С����?������<��ӼCc�HGn����!hc�3
��?q���S�'$��u�۴�yҌS�0��l� O�k���!��y�	ȶ�֑������D�O����V���dᒿ!����_ZE����Oh���O�˓
p�F��	Z���'j���~À
��<	Zp��@�ٿA�Olʓ�?����|"@q��@�0hq��3b+�L[��'��ܘW�״�� ��������'ԜH�gc�q6��k�IUD؂����'~��'��'��>A��DbE��N���e��s�j�	��M��L����O���+8�t�˅�H	�9��))D�	�X��ҟ������'H6E�kJ�?q��D)flb��Q�C�sc`�I�X�{L�'f�i>��	ğ�����ɤڐi�2I�5p��YI�'١[~��'�T7������O��d:���O�ࡁ� SQNyG,��g�t4)��<9������O�8�҅�צ<��8rS�V0'$p��AO�_a|y�Z����jB<@�iy��Dy���(��Y@�J���q���9T���'���';�O��	��M[�LR*�?��EF2]Y��g^	�Rȓ�&M��?�����'��ܟ��iޡHe�
i�����G�#1���gW�1lZo~� �<V��Ә38�O*�G"?3  c��� ���YW���y"�'�"�'��'��	��5m}!�����#�L��?A���?"�i���H�S�p�	Q�&+���S���2��-h��8���?i��|����M��O�5)�N*^�������/\I��A��mw����'��'z�i>a�	�0�	"����c`x ��B�I,�X�	���'��7́;K��D�O���|�wm�-](|HQ��<1�,D(TJDP~�T���ޟ|%��D4�ؙWL�Gr����lV�n�XDC��N�6P�$'^y~�O��y�ɾr3�'��yb@�Ұ�X�+g��	O��A��'r�'!"�O8�I<�M��f9HZ^�
U@�3P��H�%O<v�n��,O���7��jy��'�՘���OG`�uH�8U����'�Bɉ�v�����+���XEq�̠�+4%R-�G�}z�@�E7O���?i��?9���?���)ڸ2��T�R��<t�#'e��n�6<�T�	ǟT�Iw�s���i�-ڳ����q��.g��hضe�ʟ��	h�)�ӹ%�lZ�<!v��8"���"����qg��<1Ri��h!x�D�����4��DI�s� Z��R�%8���祇�m0����O
�d�ORʓ*ʛVaق'��'SbH�;��`�3'�����m��Ox˓�?���Jh�����3�Q�~�y�'(�ɸcb)�J!"`���"F�4"��'��@y�f��m<���L�"="`��'O��'���'��>u�ɛ���I	C�}�Dy�Ƣ#���ɏ�M�ǭۨ�?y���?���w6p=h`�ȶ39��+d��
	)�'���'�����v��T�`�B�F���h�ڹq%$��N�s�*�O
˓�?���?����?��}kޅ��'�:WV��s'���Zh-O�Ym)h�&�����Ii�'.��)�/V3��$3�W�.���)O�d�O
�O1��)Jab�w�z��Փn�24ե	�$�6�%?�ЈQ� ��	o�PyRg_(q](9�Bm��ke�)�'��{S�'�2�'��Ox�	��M���=�?�F�9 �\x���	����ø�?q����'L�����I��D�$DJg<�Q�qb��+��Ԋ#�߹�"�mZA~B+� �$�'��˿�wOVF�%�U�nN�!�d���<i��?���?����?���D✄^~�L�	[%�\AB���. ��'��|�̰{���<����Q���Q��K&p�"�?r��M>��?ͧ.:�8��4����^���o�-,xh�T/���X�̙��H�Ć�䓔�d�O��O��A�FF9Qp����ϖ ڈ�D�O˓rțF�>?���'��[>�Ӡ�]�pm�a٣C����+?�/OF��O0�O�S�V�<���!�
�,��5�\�wkn�hẼw%"@� �ILy�O؉��*&x�'͐������Q��d�p���Y��'lr�';r���Ol�'�M3�.���k�T�r� 6�3��u�(O���9�	iyb�'��]7Ä�SdNS�[t0t�w�'4�j�\Û֖��@W�͵!����~� u�0��-H~�D�/�V�C�0Opʓ�?)���?���?�����2BB1S�-�.8�Б��,�lYmZ6<��	�I����Ix����x�i��S���c�R)"3g��.��lQG�؟���`�)�M<��m��<As�w?|ya#�$f7��"��<q���7j��M�����4�����%��	�$#�/%�$PEd������O���O�˓Zț�eB�'��Spq�w��<���h
B6�O���?����1�H)�����p�f8;AaJ�q�'�(pv���.�P3��ԯ�՟x3$�'y�|�.�ͮ����/ Ų����'���'-r�'e�>��	�u�|���J�,"���+�&4��L�ɟ�M�c�Y��?���?��w$J�0"�'O�<����&L�z���'��Q�x1�æq�'�ܵ�d���?�0r ܱn��0ٵ$��T�����'��N�'���ӟX�Iǟl�Iʟp�� '������*n��𒳈
!�T�'�,7�ܤeU ���O��D4�Ӛ;�-�d��EL֔S�'	>A��%�'�R��Y�.�$!�2� -c��E{fł�q*�|0`�.ɚʓz����a�O�$#H>�+O)�F�J�\;
h3e	�FT|��D�Ob�d�O����O�	�<A��i�@��'��ے���l9�Ĳ���5
Nfy�'�����<Y��?)��	0=�dȕ!d��x��e��]�-9TlY�M��Ot��� �"����w+�C��;kq�i#��v�jD��'N��'��'b�'[�����
��iHC��C�4l��,�O��d�O�Ao��9}����H�Ir�I������`P t��u��%7<�$�t�	Ɵ��N��l�K~�c�0}��=(�i��f<�%�,�,��C?�N>�-O�	�O����O�T𔤃(mM|л�Ȍ@lTh�K�O^�Ĥ<)�i.�yC��'#��'?��X�~H� �ܼpT��+��e�J���D�Op��'v��Hb@��1�����2DܐjȌ$Jbx�#\���4�61��r�h�O$��Q������cE6�²&��+r�'�r�'0���W���4L�`�4
̓l�v�y1�G|�^M�@%I�����O�㟐�'��C!C���h'�V�_^`����\���I$/Q��m�{~2H�v8j!�9��	=[O�qg��w 09��X����Wy��'r�'kR�'{"Q>��F��L6�M��P�X�21��KQ��M���6�?!��?L~:��?�;��0��,M��q����!17��0���?�L>�|�t�>�M�'���)p��Q{�DܵC��B�'� ���q?yN>)*O��$�O֐�5�ё@��`kR�fK�6N�Oh�$�OT�ħ<9װi�-���'8��'X�QE�>�|��M�2O�:@�d�<���?�N>���Z�P��/4P�HjPŉH~��_���X$�
��O�����|4r!�720��D�L�<M���{/��'x��'���sޭ[�cF$"+���c��irLBe���s�4K�.O�D8�i�����\� �����O��s �B	y���I������,�pnZO~2�
��\�'+�f���ȹq���Zam���Dy�J>i)O�i�Od�$�O��D�O�����  �ڄY��[h!y6��<�i������'��'e��y��˦M�a��.Xc���џ8�	u�)�S5�
�2毛�o�ʰ�1���Kʪ6�� c�H�'H.A�"-��;��|]��ڕB�>\��a v�ڝ��aX!DM埠�Iϟ �Iϟ�Ssy2ah�:0����O�E"f�"_ ��;�F΋d8�M�WC�O��9��[y"�'���'�t�!1�_0s(�Q���¤ZA�R�!�Ɠ��n�]~�	,����D
�"��Rі�z�R~䠱2OP�d�O����O:��O�?9�ӃF�B��B��%3� "c�C�4���cٴ]̴yp,O���8��ʸogq�BAU9����Q�F踒Oz���O�i�27m<?�2.�*��Șu)�]�T��3��;Q���O���&�l�����'��'ˆ �/��[��e�`&�m��Ab��'�2]�`;ݴ��-O��d�|�0�ԃlRf�h��P�LM�{FDi~�X�<�	֟D'��!/�HC�#yd%0�n��J�N(�b��,��3޴��4��0��'g�'�j���ĉV��QI֋�r�8����'	r�'�����O��ɰ�M3Q��GBDј�%�1"�:y+#�E,��i,OZ��,��Sy��'����f��("F����)5�<b��'a2.�Zj������$J�q����G�҆rJ�X�U�4E4��0�;O.˓�?q��?���?����)�v�*5��4T����g��W�\�oں	���'t����O���>LP(c4��A5�*�i�_����O�O1�R�rB���u4O�s@�k��4AI6`�l�Q9Of0�w���~�|�U���ퟨkq۞Hb����5�d�6#���˟���Uy"a{�4i��O���O�) �>$��ʎ�?���R�`,�IBy�'��|R��^����N��5�nM:�O1��d�6k~�C�+�g1�b�c��b(��-�< �a� 6=��Ŧn�����O8�d�O���3���G�Y�zy��m]�P�sD�0�?)�i��=�0Z�x�Ix�ӼkO �RŎ	����a���!ӍE�<)���?9�?�ū�4����&Tt�pK�'�� ��"�Һfhݩ���*�8�y�J)��<ͧ�?��?A��?� D�0^� ����=� rG��̦	a�(�џ ��ڟH&?��!=�Lm��m�:f����!.�蔗'D��'`ɧ�O|�5c���6-Z�1�`���T�DH��7B����RAIP�	y�d+�d�<y��
�R����1jx��]8G�ԟ�?����?���?ͧ����'��ҟ��f��)�Ԩ���I��r�I�ȟ ��M����O�$�O��@0,%�l!������J��
�o�6�??ɓjJ���IJ	��'�����ŢXG���f��lr�K��<����?��?i��?����OC?x3he��6=���8#aU���'���a�TI*f �<i����G�Љ!t��??	� ����bXL>���?ͧ<�<�+�4���&\bhX �:5��xmL�v��!� �?�J1��<�'�?a���?�Dmްw� sGn
�X@(Y�%���?�����aiwI�����I���O��Ы�k�I�hi� �5:Ȉɩ�O ��?1���S�DjǢ1�ݨ��:pڬT	N��vl�l['!̨���O�ɛ6�?Q�c;�����������o��j�"�����Op��OZ��<�%�ib�Ҳn�@ɚ���)��X0�`�͒�-��I��|�?�,O6����"px��C�:�)T �X�N�$�O�e�2dӾ��5��##�S5+����U�9J p��MK�����yyr�'(��'���'.�R>�g왺
�>Q�D�V�,\�lAUb��M�RJ�'�?���?Q����y'E+q�9�$
B�N<^��!A�{���'�ɧ�O�����i-��&W�M@�|������Z����	�5��)-��O�˓�?y�wf�� �3��pk䄏�n������?Q��?/O��o��)���I��|���6 D��7Ě�i4����"E"t��?Y/Oz�D#���RBf|��f��z�2���"��+���%�Fe�D�ƚ*W�MJ~�dH�O�MX��'7 ��d�ԝ�B���陞<B�"���?����?����h����N���2RB�z���{�*��Rۦm�3eJɟX����X�?�;2#z0q��Ӂ:E&�j�U+�}��?����?��g�=�M��O�^!���	 ��a��^��-
7��Vm�J>/O����O@�d�O�d�O�<ڧ��Ϭ�S��}�x��<)`�i\��j��'b�'T��y�K�=H=h��`!�:6K�E�Ό>���,��x�)��@@�!�@ʏ�@��r�N�x��xb�Ȧ!�+O��de���~�|�P��{3�Ɵ#C�Ъ�;x	Z0�����,����p�����Sy�Hw��˒��O�9��HI.g���!� �L�Q�<OH�D1��Qy�'f�'RA97a͗�X�u
�b�pa�e�{Q�6��8H�CU�T�	��"4kt�RC^LI0D�,����9O*�D�O����O��$�O��?ea�'ܚ~0�q+ �
�.4�h�+�֟����� ��4��*O|�d1��Z fӼ=��A�;��')��FP��O��$�O�5�7-<?�Hܴ2�t�w�A�=��0p�R�j�@s/���%�������'��'�X@ᶋJ2~Dl}����y�X����'��W�h3�4�8tK,O,�d�|����_�L8#��4Dy�H�t�Ni~RP�|�I��&��RW�!�!Ϭ� �΅�vހ�!ue����iY�i>��c�OOL�S�'�yc��i��;8���3��O&���Oh�d�O1��ʓ:��Έ�K��tS�n�22�,�䇎G0���[�l�	]�����O�����͓m~�y�!@	�\�����O���S^+6�4?9󤞟j�r�>Ոt��$0ν�.��HB�q� �Idy��'0��'�2�'��T>�0c�H?;,:9���8$�Ago��M����?���?�I~��?�;2H���`��p��i
�jſm�TX"���?AO>�|*�����Mc�'m|�P1�+,h��ǜ�w#�؛'��BYm?I>9+O���O��8rl$	"���'�0[�T��T��O���O��D�<�b�'��y���?I�5�Nm`F�E:�-ḺT�@x��\���	ş�'��J���$Fڐ����]6B� R$+?)��=���z۴A��OoB���?٠J�}��K���-A`��d�?��?���?��)�O��צ�&\qx�O���A�@��
z�|���<����yG��U�(L����$���Pc���yb�'+�'Zd�xƽiq�ɤ`|���OjV2%m�)4���z��ȴ_x�)-Ba�uy�O��'�b�'���"���*siͱl� ���Ʌzs�	��M�&o.�?����?�L~��1Z����E	��3�f��Z��@(O��(�)�S ��$A�� ��考ٸU/2�b�I d�d��'�Ve��ʁ�4���|�Z�� l�:K�Ȓ �5\Qdk���؟�I�`�����fy�L~��AW$�O١�HJ�>����J/q�zXR���Ov�$;�IVyB�'��%
 ��B�$E���+;`�`�Q7���)�'����B�?��P��D�we��x�$!����A�1?�'Q��'��'|R�'��$Հ��6�Q��d�&�:ԩ���O����O��lZ�nY<�S����	T�:
�VA)7h�70V���%�1�0�'������ӹK�nZ|~��³Հ 8��v�I1��)
B�^(j
t ҇�R*�~r�|2Y��Sퟌ�	��P�5�C�x� bbE�3ژآW�Xßh�	FyR�w�z0���O2���On�'>�`y�c/�sL)��m����'��	ٟp��^�)"�ߩ`j1�0���
���hi�&s�D���̇�/Ӟ �*O�I	��?)�"��1��U� �[�0���B��k���D�O��$�OT��ɳ<q�i�f�*E$�3��p���[��i%Q5RF���<�?)/O���#X=�6�Z��&u�4�[:" ��O(�	��{�2�UO���.�O����Ӭ�)�B��G��Z��౛'��IşX����h������y���+�T!��Ţc`Lڴ˗Iy7��%����On�%�9O��4ﶕ��N
,3�����
�Z�P#f�O��9���ƒ5��6w��b^��`�*����/��K�ov��HV/2MR"M�	oy�ON��B�d��RC�>a�@�Ok��'@�'�	+�M������?9��������)X��YdJ��ш�Z���	ޟ�&�0���]�%�Nq�6����>t���+?�dm
���!���Ba̧����C��?q)Ԉ,�tM��E�(�}�����?A��?��?���)�O�HY�J�H%�9�&���\������Om��?�&h�'
R�4�T��XW<	 x���K�6OP���Ot�d�'I6M7?�;U���s��`~MC�a�+���u�Sxv����>���<���?)���?���?����A4
�#�_�3�PBΑ5��d֦m�0�Rџ���㟨%?��I>S��x���ɨtp���O8H��l�'#��'�ɧ�O�BxY�eO-v�X"��!]�<�
��v�fC�<q@��ZD��h�	my��N Au��1TK�d�Z��"'D	#q��'�R�' �OO剥�MC�!ȑ�?it,LT�"U�J�n�`���<����'��Iߟ��I�<�Ff�Z�l��b��?e�hł�7�	o{~b�F�����r�'ȿ��I�e}���Q�O�kCH���ȗ�<Q���?1��?i���?Y��4��EI �B�������Bʝ+��	����4&�NXͧ�?�����P��0s�J>^�ف �+K���HM>���?ͧy՘�yٴ��6/`$�D�@9fg	����Q3<�kd���?1v�0��<�'�?1���?	C�wT�1�jgp )F,S��?�����Ē㦥��&���x���$�Om8	�`� ���X����"�����Oh��?i���S�T ��R���*3�Z02�@�V2�8�� "x����U~�O���OZX9I>1�-F�A����&P�Sl`��P��?!���?����?�|�-O�PnZ� ���`\z�Z䑶�S�4̈$�FJyr�'��O�ʓ�?�@_��Lݡ�(�bnȕ�푑�?���mbH��ܴ����*{w@-"�'���H�d{��E�s��C�%фb�t�Iwy��'.��'��'�"P>�:��V��a����#:i�,��MS��_��?���?M~���?ͻEm( [�G����˵�Z�M>aY���?�I>�|�r����M�'ʖ%��/�N$}��.[(��'�b���`�ƟȲ��|�P�����XaR�ͺI���&��>#��	D��ߟX�	���jyR({ӈ���L�OR���O���P�ΚSvz�i��E�i��e�!�<��iyB�'�O� �pY�[�X ��I�/���ȑ���@��S#SjR9��cM�S Ro�cHߟDbP�N=vCƩ��U#U�0eZB�	ퟘ���x�	�G�d�'^�!�V#e}8���DͲ='2����'��7-������O��$>�i��`���N��0�`�%;��`1�c�H�	۟X�	 q�֨m�o~Zw��pA�O{�����r������Gz ��~�Zy��'M"�'"�'���Ƨ_�hk%�::RH���H�t�剀�MS����D�O�������hv
Q�PeR�J����C���>�˓�?i���ŞB5DXh�U3%�*��0�n~���X<:J](O���B&ٶ�?yua)�D�<�q`#	rR F�o�=�`C�,�?A��?���?ͧ���Lɦ1��J�̟t���]�{x��٠�	 q�q't�\�I]�����O����Onq��@
2������(������s�6�%?��S�Q�~��N�S����JN�i"u�Ai�,r���#��{�0��ɜl���2�Ԛ��H����1&>��	�I#�M$m�g���'��'��u0
��6m��,K8WH�)'�|��'��O��Ƞa�i��i���Q"����E�� E�RX���;n�9�ɫ[]�'��	W��T Y�j�u8��� iU�W��|Gxw�"����O���OF�'(1����ir�u�	�%G�>�h�O ʓ�?�����S�ăҕa�R-�G��I��2�C�u>(5�j
j"4`K�X��S�8/"-Ip��O\̓�)�n��
�)1�B�	�M��⇽+���!�c��jy�lC'.���ܓ���?����'��I՟�x��O�����g�?t�z�aɐџ�I�E/V�n�Y~"�ŭ:����'��1I0�[7�I�Y �ǫR�]��d�<iߓu>v�3�O�pΈdH��B�����E�i@(��F�'
2�'����4��H;E�X:nn���NW/`�Rm��#�OH�+��)�2��7�|�� ���!f
hz�Ⱥ%G��5��X�2O�`��ͬ�~r�|�V�ؔ'��P�j>G�6= p��?C0��#
Óy��F�W� �2�'�b�\�Jʘ�����1@��`�ӄU^�O^��?�������Y�*�P�:,���K$~]��'��uY�"�j��f�6�I
�~��'tVTU��0,�	�e��[��x
�'��i���-?5d��@�Xӂ�(��'��7�B%?
��O��d5�i�9��Xw�|CF
't#�\���O����O<�D�� '�6�3?��n̓A3��S�"4��WL��en0D����4�ڡ$�H�')џ�	�Lתq��8
U�_�:E���$<?鶾i�\���'{r�'��a�W��+Xzq����\,���<���?H>�|b��Ϡ ����d�ܩn��)c��
'_U۴_��	3�Vp��O,�O�ʓj�ꠓHP_)�H���Z��R���?1��?i��|B+O��nZ�P�vE�	.Z����5.6��ԯ����	�d�?Q-O\��Or�Ӯ&=��{v���}��`�����=���b�`Ӻ�_�B,b�K韊"H~��;���"s΋�V9��YpÞ����̓�?���?����?����Ohr�Ҫل2���¤�ZfLJ��'���'�6M�%y(��O���#�$��b�T7A>��k�(_3�O^�d�O��@9;�7�<?�;>�n�-g�ٲQ%���� =9������t�
�O���?i���?��Q�U%O &��Wb�&&������?),O>�o�p���'��T>yS�#k�@�� Ź?�Ȅ �`3?I*O���O�O��9��y�B��.H�A3�ȹ@�ƥ�3d˳we��"�fy�O�ډ�	��';�ؓ��ΆCC�Ec#腻���9V�'2��'�����O��	��M[��<���i~Q��&�"�z0F�!i�I���?9,O��
�D��y	
��D��Q!��C	h���Of]��jw���Ӻ���r�<Y�*��p����T�"���2���<9/O>���O��$�O�$�O��'1��F�Qv�U�cN!�����i�L��s�'w��'n�Otb��y�⃆t�4����jۦ}�#�2�b�'8ɧ�O��A�i��d���YKI�7��9��F�K��䟵�j�I��6O��Ol˓�?Y��c�Xs��
�o4�Q@�]r��;��?	��?�,Oz���(�:��O����<Hk^�	�ᒽA��܃djQ�W|��O���<y���?�J>���:}0���Rd�d�����D~���?�p�`t�i�������'4���x�R���-�	C$�IÔ
۲X�R�'�B�'���s�]ئ+݀z&�{d�A[��S��ƟT�ݴn�$�y��?!����?�;-�j}�/�	C^pI9ԯH����?1���?��$�=�M+�O�A8���':�t��D,�$�	&L�	T�I>.Ox���O��D�Ot���O
�pq$�V�E���,r��Њ�<ٶ�i�.ٺ �'�R�'��O�2Mԟ߬0�&�\�>K��� �O���,��|�)�S�ƈ�mĀ~�l����0.H���A��M�V[���qEB�	��?�d�<��G2g�� �#�Xg�UsSɉ�?1��?���?�'��dX˦�+�c���s!i+\h��"�@�&-��@j����	m������'ZB�'�r��x2T�IЉ�K(���"ޓhdJ�1��i��I�x�MkB�OyT'?��1Rْ���!%��Ҷ|�����|�	ٟ��I��X�	w��W= �8�(�>]Z�zeW$X��Q��?���|�������'�|b�"՘x��l�Lt�Zt���E��'Yr����%R��6�����\�J���bI,��A��2M�6��5�O�OXʓ�?!���?q�J@�`�#�
�)�[2Ne��x��My��r�,�a�m�Oj���O8�'-����%�ހG5�XQb�)�6=��?�.O$�D�Op�O��J��0Q�[�6y���7�e��	�2�lZ��4�$�)�'��'���3~�
XS�(�0{����f�'�b�'�b���O��!�M�0�V������BE"��
�B���aQ��?����';��ҟ$�#��?�*�ye쐎0���Ӏ\��`��/m�J]mZt~��O�
l\�}��F4^	�PB���3��SǨ��<�-O��$�O8���O����O�˧DX��׊M�ki�M�e�-�f,ӆ�i+��E�'��'��r�4�h �v�,ʅ��|تIz���O���3��i�:[�v7-l�КU L�_-t�ZFI�J�@��shb�`�5@�/e'��4���<�'�?9!�� ip�ָ~X���G��?���?�����T֦	0qN������ڟ$��gC	K� �a�Y5
2��@ s�����'e��'�'�`�¢X�HZ���RĚ�<Gj���O�����C06P6M]S�`h���O\����� 0�&� �	d��,�Ol���O��d�Oܢ}�;A8T
���¬b7⟁L�T{�}ꛖI
U��'�"�|���yW�ڢ_M����	<��(u��:�y��'@B�'TDA�W�ie�i�e)5��?�u�
t��āAj߹1���it��)I>�'���ϟ(�	������\�I0J5�� �������F�'p�6��Y���D�OV��$�I�O�0k��(tr(����[��D"2��<���?QK>�|�ы�a�? L��&g��$��߈�"�z��jӐ��'�Fd!6��B?�M>),Ov,"r�6$�4��τ,|��U�'��O��d�O �$�O�	�<���iJ8���'��%�\$_H
%h7�͗GAT�'|�|��'/��؟��I����$'ɳ|��`��9RT쨙V���4"��n�m~�f��4��Ӧ6��O�w�((�� w��LF~���쌋�y��'r�'�b�'7b���]��ٱf��3j�h�qÈ|,��d�O����ʦ�S֨e>m��矜%�Pcr#�R[��;�
�Z����u�	��i>� W����u�&^�p�2H�ˏ�m�\�IH^�X���'���$���'2�'s��'�#����\5�`��"�u�'��U��޴;J&�����?9���I�7/%|I�b�7s�8��⏙6���O�ʓ�?�����S������ ��?RZ��.���Q`���5���G�<ͧX],��F�	� `��@��1���P��,��Iߟ��I���)��wy�ea��@!H��� ��0w�^��e@�=�����O �D%���O���?���
>Iv�r�)Ó�aZ�k��?���Mײ���4��$G�=�4q��O���<	#��`��S�^hSS�S��j�	Ky��'y�'��'�2Q>yC�W 7��T�'�@	w���1V�H#�M��-ۛ�?1���?�N~r���?ͻ+� �	G�O:@t!���˽q�f0����?�K>�|R�����M��'u�}cVOõ`����Z�k��;�'�44
V�Iʟ����|bQ����ϟh���I#<�A�K�f��yR5�X���ş�	syB�a�\d��E�O��$�O�qJ�l���@�+C�v��Р!�Ivy"�'�|���@�����N��!�j���(t��d���{�H%?Q�B�O6���M���7ɜ�B�)	����R���OT�d�O��D&�'�?9Gn�~B�$Ɩ-Zn�e���?9��i����'�R�'��O�[?3��5���w���[�4q��Iݟ���џȤ����'G�-x6o\Fr�b&���ID�S�O��=�g�������O��O��d�O���_�l��8A�k��@���Y���B� x%���?)���?�H~Γi�b�`�� ��`��h�.���-O�D�Od�O1��e"W�����⢎�<(�L���#i@�7�Mcy�f��(��k�
���b ,z��3��/�. I��"%} ����; =2�L�2���2��Ѝp��c��&Y|DJ �4	�-�C��J2�M��j���N�7���B W�Ek��2���FX2���hK�vi0		%H-J��4�EE�;���W���)�I"#�Za�硎5�$�S+Ĕ4�A�q/3s
�(0pB�����$9"���Rd��	s���-�"��1��̐Qfr��pO³q
�CSN�y>�|�����㒌rDFD���i8���	c �Y��)Įue��nZ6�L�SE�� F�t�U.Xe��#�4���O4�O.���O��Pb�O �!"�S 
1RX��L��\ �i�ff[w}��'���'��Ig��i鬟���S�@���EH�d|��Q��Q/�4o����%�l�����Y��`�$��I�K�&t��z%��jې�n���$��zy�To���?q�����T�
����fA��h��t��]ۉ',��'�r���'��'���;�>ա�e�1��9	�ōQϛR�,0��ɦ�M����?������U���=�!�Z���ieM+$4�7��O����$&��@�}���L6Wt�+��
�mp��v��ɦ5���
�M���?)���u^��'T���K�=��<s%P����lb�L�`��1��P���?���V.(B�Y1֠��f�h �eޚf-���'���'�XRS��>9.O2�Ĥ��q$C�!���`bJ�a�5��kw�ԒO������n�ş��I��P�!΃S8�ұ�ԵohX()�\��Ms�<"|���]�0�'�|Zc�p�G�Ϗ2$HP�WD��­O��ZV��O
�D�O�0���ӄGk���aƂ h
0ݺ�
V:){�Iryb�'q�'�r�'�Ę��N	?d�D0�ħ���A�#��'�Z���'��	&b���Oo�8�ơ�i����
v<N�+ش����O�O����O4��W�(²O�/C]��z$�_�P�ް�#�>i��?Q���򤀷n�4��O��O^������)G
`R��K�Ԃ6��O&�O����OpqK"�	*Ap�Y�Bm��r�ԑɑ(�b3�6�O���<ق�� L��� ���?AqF,�/A�~�TN�	p�"������ē�?���u����۟���b��<�xl4��)SP����i^剺]L�ڴ�?����?��'XP�i��@�^&I��p*G5N5z��d�>�$�O��!K&�	iܧC�%EC�W�D�PcԊYcD�l��Ħ�S�4�?!���?�����Ihyro�:T�n9��-�@@p�!&W� �^6muܾ㟼���[��X҃�ݫ3�x5Cg�O�"!=� �ilb�'�҂�0g�BO��O��I�\��YP�EMd�r�*]1g�@6��OH�Oʁ��yr�'�2�'�m�RP�;�R5�!�%n�7��¦���9.IlhZL<�'�?�L>!H�dz��I�i�8���� ���'��U���ҟ��IVy��,V�ܝbŎ�4uB���a'%���ku�=���O
��,�Į<�;xyz\�W�ˁ&}\5c X$ZbemZğԕ'��'BW��#�gK������2�� �-*˔��#�M ����O��$.���<ͧ�?�W�ڂrټP���ǈ�X]�&�NI+�	՟��	�L�'~^�Q�<��\v�? ��k���n����W��쉚c�i��]�t��\y�O��~j�u� �'
�w� 1�WZȦa��ɟ@�'���Ib*�)�O"��ƶ}YF+̺ddl,��� 	3�j���xW������'?�i�!�f��o��E�o�-CIw�~���j���&�i���'�?�����ə�"L�!�K1*�C��{��6;<����?��������4}f�0a�P*�x8*!v�H�m�[bn��IП��I�|�Slyʟ�`2��q3�Ϳ�JIa�D_{}RaD�O>)�c)R�_A �2�X�s���o֑�M���?��cSz�2*O��a�d!�Y�Y���閫�#�z�[�m/��b�$��D9�Z�g$�Ȋ�"�3ഴv�t�v���<{�RʓF��Sc�^�(�`��u=��P�G�Z����xBN�0����O|�D�Oh˓�0��CE\�sd�pD�D�P.���c�K)HW�'���'��'��i����D� IX�v��!��Y�Dh����,���On��?�b��:��D��,vM��PV����5OD��M3��?a���'m�>{t7J�F��0����m�D�2R��d��'�BQ�0�	x�i�O��i�;Pޥ��/]�HwLX�k��D� 7-"�I��@�'���SN<�7]�л3)ęO_���Q�B����EyB�'���@�X>��IڟX�s��:�J��y�fh��� �9q �r�#-��O�ʓ(eR1DxZw��ܺE2q-��R2h�
g0]h�O��Ā�c� �d�OZ���O��)�<�;
�%��t��C�G�Y~�o�����'ä1�����յ.b=��E]���y��ժ�M��
�!3��'{��'���
&�4��uɂa�V�8!!KW2�-{D�^��!�	�D��b�)��?1����:\�e�[3�H�v̓"2����'�r�'�DhY�h8�4���䱟�£�ކͶ(9�,̓@*�E+u����9�Sj��'�r�'����2�U����2
�xM $,� X�d6��O��rT��o�i>E��Yy��'��C[�^� �q��/9ֽ�wa$�$�ORʓ�?9��?A)Ox5K$'W4�h#�߳f��ĂG�GA�}�'��Iןȗ'���'\��@�VU�e�	w�H�4"aJ�'D�I�������'[p�&jj>q %�ۇ%�@uER�'T��r+i����?�)O����On��"54�71JpDjЪ%���#`Wz���l韌�I����qy�I��2H��?��PZI,Q��1�E�1-b�Qp�xӘ�D�<��?i��o�����ɄT��23��-D�RP�F/S
f��6m�O����<!G*��S����	�?���nT ��0J�J���iB����O\���O�}9w9O��?�O٘,K2H9! Qj��ӊ�X���4���D4��9lZ��Iڟ8�ӆ����{�ٝ&��I���9}��tjױiN��'���'��T���}��)�6�j��GF�q�`MRD�����S���0�M���?1��ڱZ���'��i���P{�b��()��GDi����w8O��d�<����'��q#!R&I�\2b
�m%�(�(dӠ���OD��Y�}6���'��	러�%l�U2��H�-��=��+2i��mZ���'�`����I�OH���O�U��N�S�L|���DuДa�QӦ����x�O�˓�?i.O����j��Nx�pR��ε�ȽÄT�L�#Gy���I�<�	��(�IKybGߩg!���q��i�t|I���Sk�r���>�/O�D�<���?Y�q�ެ�fA՚V�F ����\X��B��x~B�'��'��Z��K� ���̅�a'��ЀK���tАs+X/�M(O���<��?1�x�ϓ�~�i��E8z2���pd�bN̊�i���'$b�'0�	�w��#��p��Ƅ5�q�Ղ]�.ժ�)	6[K$����i_�Z���	��x���.��I�x�S�N�:e&8�5�fC�8X���oZ柘��ry"�ߩSON��?����E���4��� �n��s�4h��@���Iџ��	۟�g�y� ��yӟN1��	�PU3��E�tX�Ѻi0�ɏ%-���۴�?����?��'t�i�)aA��]P!�ɡ\��J�bf�.�$�O�!�U=OB��?����bR�1�hP�	��,[R����M/0�0K�4�?����?a�'��	_y�(L늭�sΖ�'r��i�I�7�by�'wY���J��j�}c
��mr*ՑT�����Ҹi52�'��M_�������Of�	�>3��HA��8� ����Wֶ6��O�ʓM䖄�S�4�'��'2ހVb|��5�AO�	7v钧�g�H�d�2&?�'���|�'Zc"zi	�B�<+\x�H�Y���4�?qO�<����?����?�����D�H�^1�qD�=L��4�'���:�w��s��?1J>A���?٢��1{H(E��*&0q"�biDA����$�O��$�OD�V[:`�6�$($���Dq��R��[O�T ��x��'��'���'d��R�'����MȔ��y2S$#1������>����?I������{gZ�'>a�Hڵ� ��c�'� 	j�.�,�M������?��(�������	%UY@�bc�=:��E-��U�b7��O@���<��ߪX��O���OI@� ��&�p��LG(0�U���3���O��ĉ/4	�>�D�?-����5��8'��1 ��&�wӚʓ~,���iKz많?��'��)� 4A��@@" ~ՙe���u���T�i��'�I۝'��'�q���A�W���*0�jvZLt�ih��#�-vӺ���O��@��>�A�°c�b�Y���5UA�Sv��������y|b���O�It��Bt�m�s��t���%cBԦM������ɬA�f��J<)��?��'�J�W}�����u�H*ٴ�� �T����'��'�����vR��{���K��J��}�J�D��]�d�&�������$�֘�G�p�{����xF�����:!���<�89�������Of�D�Op��4c��'����7����-sņ3*B�O���(���O��DK�2X��h��Y�(�2�pE� X,IA�:���O����O��0��u8�4�*`U雫7�&��Q@�î��R���	_�'}�I����t�Z�d��!�#�';��}˅�$����O��d�O&�(�x|�S��4'Y�T
��X�Kۅ���ҕ폫w�6m)�����O�'R���Ǽ/���R�R�7��� �4�?I��?���WYXe(�F���O>�)B�V�ڃ���%�
���� F�\$��IBy�G��O��F9F�����҆Y3v�S�fE7��X��qQܟ�M�3Q?a�I�?b�O2��V�@$a޸XEc?]?,�bxR%Ύk��OP��xb��z���D�� rRl�4�M�j��?���?���:��?I,��C���r�����k�F	������O}�B� �O1�,���xd�p��#ŰG�f��	0F�$In�ԟ��	쟠@!痚���?I��~Rh�!C1�r��7#7�<����'�H��y��'���'�}���(rLz� W�
�gq���2Dx���G�j�:T%�4�Iן4$��X�Z#j���-��)�x�q�kd�F�K�P��<��?���dF�s}v�2�lBD��D�J#(�<���gXl��?�N>���?��ă ��ff  ��ZW�ģz��u�<Y��?����d_�l�: ϧ `��� s2�[��L����&���	]�����ɸ+�"�} X5� O4$�K��5��'��'�b_�`Y���ħH fT��FԡNr]0��Xw��@���i��|�'���X<��'�pG%[�Il��#ؗT{@�s۴�?����D��\Ե'>q���?Ip�'K,���C�N��QS��ē�?��&_F-Dx���P�������&_V[L��\���	�&��<�Iߟ���ϟ`�SgyZwϺ,#'J�j��=)s&�.t!Zq�4�?�.O�\�&�)�IG�L|��3��K�wJ�Q+�-
�^�F�/p�6��O����O���BC�ǟT����-,]#Z��8��/̭;4d݇������:���L*EV��'gC��M��?A�}�m��d�O��	�i8܋���_�t�rrO�J!��d�O��D�O�p@�&̃{�4[&�W�|l�1��Ǧ��I�5d�H<��?�J>��M̒��h'a@J�pf�W��$��'�r$��y��'�BV�L�I�"�.@h�JĈV��� �\��A6Ȃ@y��'>"�'�'?2�O��2u�ċ|3^ ��`4O�T�ҺiY�h��OF���O���<q�^\��I�r,%�g��:�~��@�-9A�������@�����	(ft�-� `�#�$��#CB��'n�'Z�X�9��/��'F P��O&��8)���W�h�J��i5�|��'42X���'m:`{��#c(�*��ԝy��ߴ�?����$Y;.`��O�b�'!���͚2]���"$�HȔ� lZ��듡?I���?�Fg��<9�����?��t
�44<��j;0�)Y"�w�L˓���qսi���'r�OV��Ӻ���&Q�U��L�FY�d{ ��5�I����Hb���cyr�)��j>�����!!x��:~���ꅶP��7M�O����O��Av}2W��������퀫ڲ�RR�U(�MS����<Q����*���pPp^�5:�!���0pE0�i��Mc���?���|6Z�:�X���'�B�O��s�I9���t�$F|~h�iq�R�8QBh���?��?�s��rgp%pFD�D�Ix�ო6[�F�'&���G�>1+O��d�<9���`n4^�4P EL��{�V�RʏY}�B��y����
�h]B�� dI;�ĈU�y�N�*��0q�.`�@
�$�y�G�d`�Kv'�]��QU�,��O�PY6&�gp�)�%��R*ڄ2��ohH�I �E����VӒ�@��d���(\T4䙊���� @�����N2�:%��Đ�b�b	j���"H(��		�	�~��'H�����&��P�AnE�u�,`�Ы^=*' ��p�R�&��`���M�1�!Rq�τ1�EJ3"K�}���a� ~�<IeǙ42��'��>8�$H��G�Y����� D��'>�@[�D�$8th��n¢;T�Gy��ء
���#e�@$Y����i`6<���SbJ�`�f�:!�F4k1`��>t�u�f�%�I1O��d�O*�?�Vc�		}���k�7G_���6hy������X�����׊QԾ!�Jl������w�	�M0�U��
�	��X2�Ŋ���.J����O����|2���?q��?�@J�/���2'i��h� A�<SQzı�O"D��i�bK'�*��c>�D� _d���!�5H4`�`V-�
�M���'d<|łŧ�P����)��� �q�e��V��h�%��?\���"ٶY����O��S�}��*U?B��C�9;d��V�9jB䉴Q4*y+'�Z�)��L3�,<�P"<y��)JCl؍D�z�D 
8��'��?1���i�B��?	���?���
��N�O��ć�Yxܬ����-aĐ��f�F.(��d�6��"w"¿-W�ń�I	I�fYk"FT+^��r	��c ��I��K�6���j�*UX8��jE �	=$��ǉ/K�N��炷��� a�O��"���D^0:�rB�)H0T�&��x�!��d���'/I4/������6���Dzʟ����KE�i
��� �iy���:����')b�'�b�N��'V���! ��d�UFG(8�Vh҃��e 	��/_8��"4J��	ִ��$�eQFU#Ō��-��=#TLI4<� -C5��Q>�P�4�Ҩv�Z��ҖQ�'�XtCfh�'*Ɩ5���Q�{��Hг�	r�']0�� ϗ��i�K�%!#H�;�'i�jiȿ
������n��'nx���䖣"����'�Z>�B�k�u٠���
2V�F0�&���LN���I럠�	�DͲ�bރF�0 �g��S����H�x5 ��p��a&��(Ob��h��X���Qg�+D�X��ۅ*Z ��d�bS6uY�L(��	C)Z�d�O��?���]7� D�.FkC�pj6fn�X��ɧ9<(xz�eKt�@�E��D�����R�ID�%�AÓ�_1
daGߘ����*s����4�?I���I�c��$�Oz��é`�0�,% �4�$���*i ��?�y*���0W`V`ܴ0P⥂�Ζ���Fx���'��|����
�ԡ`����f��$bv�����ޘ�����ޔ�4����	���@��y�)�n��K�N�p��-��O\8Gzʟ2Q�0�6U�Ե1����T��pi�O\�d�d���`�O&���O����ź�Ӽ+%�?o�)����% ]��˥��e?�T�T_x� ���9z����w�\�}i�P�����̺�C1�O��(1쁍�|�c+q(����Ob���'�{¥B�\�q���1V,�0I3�Ƨ�y�E�9AK�4Se��b��ro�#=E��gQ�L�Z7���t�����'ϸ^� � ��ˠ
����Op��OL����O^�k>�YSD�O��Ğ=5��UAB(?�0X��a)t�|Mל��QVj�)�l��8����;_�|2����?��ݖ�:�c�>X~�9t)��~��ȓMY��+4��?�`��BM $6:��ȓJ^jH���dx[3N�>e���̓"/�O�5�%�릝��ΟT�O ��#ˆ��*�Y����'qr=X��=�r�'������T>	��T�,����W`�&�~`���&�8Q��D�䎕�B49�TD��fO~E�a�^0�(O�C��'N�>�ڷL]X�	p"T�Q2d�i�"D�l��d}��-:T��8r1H�R��>�O8l$�<��(�쥄�2IR��� A)��D���o��h��k�ă��$�"�'����A�E�p���!��@[1`�)w�օq��'F1O�3�
;J�	���L֊%{CÜ�����G��O?�$[)N���Rt��("��.i�B|ѐM�]Q����Ol񩟍B3(x��͜~�L��"OΕ`�K�b�����g����	&�HO���A_.�ueY�L����ʶ������hz7�4ۨh�	���⟨ ]w��w�����B�G��9�.���Q�'� �	�� 	�N����U�ww��VuL���?X%S�N���I�@-A�I�wr���)|O2�A 	�=P��1�dJ�^��"O`�u�\;v-@��l9K�Xs�	n�����!�B��KQ-;@���AģַG�zh;�����I͟<��Zp���I�Tͧn��D�I��LJr�K� �j��ҚLB�h5+�O��0UW���A��L?���ć�v]V=g�#�O�}Y��'v�C_�&,� +
y@��B L
<�'C�':�O�S�x �$��`���ꢣ�#N�C��B9`�x�R�2����gůx1F��3��ġ<)ueX�f���'k�Y>�Q�P Wđ����0	ʂ$���@'W)��럌�I�L#����B�S��g�8;����\A⩊!���(O�e�����L� b�i�.cÈ�a&!��^ꪣ<�定ȟ<F��  �y���Z���S���1���:�"Op:�nF$9%��0�b�#FV!(C�'��O(q ��ʺ1p��a�H����"O\�ȡ���:tѡ�κ�2\s0"O��i��G�4 �R�6��(#6"Oj|�c�ؔMw�(̕�RpʨR�"O(��G@�<@@��8z�|R�"O���H��<�� %$�1�P���"O�\xW��
O�"���b��6�Iv"O����^[�����&+�J��P"O�9R�d�~�%sA�@{" ��"OdM���_�V���C49E�E��"O���`��t�,�Z	Q.\cz$"O����jA
��`��:d�Bd'"O���g H�
>�!k��^�U4M��"OXt�wŉ�@�
� gc��wm��I�"OqA&c�<���C/S���"O��	ъ6il5��BJ1־�� "O\-(�
�/$�L$4�� L���"O.m���3$�P�8�Gץ_ǈ�"O���/�F"�3��m�V)kP"O>(j�)��5��za�ڡb56�!���Sl���򠘬Aa$U�pFy�!��"�*�;�#�(2BR�B�۹Yա򤗧5o���r�GB��U� di]B�I a@D��T� 9�℩u�ŉ%��C�	86��3�S�K���<:צC�	Z�x5Ґ�5����3(ĴnY2C�I.�&Q�W�8gl9��@F�Ck"C�IM� `rc!H_U<�����k�HC�	X�11qƂ�j��M qo�r�C䉺�B���G�n.�AA�DY$g�
C�	�����D�G�Z�MX��Փ{�B�I"+:��"Uo;�~��A�>�rC�Y�Ƒ9d��9T���`Ҡ�NC��
�.A���b>�
��$"6JC�əG�>k�^��T۵��
Q�bB�I�T�T���˭G�		ҭ�B�I�2��A �#eC"����[�� B�i��F�# ��Z�Lڂ[�C�ɏo0�
�Z>�u+R�VQ�C��^���92�����Rg�x�PC��1#_Puc�|�@M�0K?]�lC��,RO,\��`�9-ʔj%�3�0˓m���h��'�ph���T����%Q��Lc�U��l#s�'R�@��
M��8F��b�'���H4B���p�jPݷ
�|$����F�=������,b�R0��ЛJ��Y�.B���C��*Z��Ac��r��� \��� eH`8�8�<E���V`�,���ړ��C��1� p�ȓ]8}Д��bA���� ��j�1��(�4K���]��0Q�O�]���ƣ�
yUl�;51�O�u����6@R��g(�r���-���Ѐd���yb�O�>~X�2R΍.��8����(O���N�:v�>�Ga��&i�!a��$��q �f:D� &���"�.�d�šC�H	��͗ f��)k��Cb�S��?qc@"kܝ�Xr8A�4�TQ�<a�l����h�o��{�|Z��Py"��y�����?$$�E��ލ��*�A>�s�	��>��OT�6@���-BGY��q��͟˨O�Is�$.�'��C_%�
�� ���Fy¯^/�9�&C>ʧX�.T�����4U�a�w��-��;�������	¬��@����<t�0Ҥ��1h ����ȋ×>E���4y+j��(�А)�F�����Oԁa��,lO� P	���!����B�e3a)G�O�(�կ�vۉ�J;^��7m��Y
�\a �ܷc�|�1�B�:e��|"ƕ	M���k��C,v��	�7 dba[vd�k���D}BbV�K��>uIF�S�[q��k����@N'�	�dT	ƍR�_y�"|���J��`sd�N�3dMB�N�J}�!�O�>�
eN2c��E��k2(�Z5���T�S�J)DY�ҧ���m��a~`5q���([rp��2�yB
hN��W�$T2�r����D߽n�0�2��Y���r���To&��"k�>d�tCD5D���_�OB$�jbNџx�޹���&D�LK�l@-nqԤ96dd����?D��sQOل8N��E��*���G�!D�t�m��(��+��ǌ�8B&,D�����2+b��B�/1:�m�gE>D�TÍ���ي��h�P���a:D�Hb���[{�I���N$]�Ԩ#D��5
�%R�1w�>����' D� �EoJ�>�P���h��d���=D�ౠJ�0�4C��˄P�~�	�%D�\ѷ�M1p��Y�� �h4Y�g$D�l�qK�(��!�\�B0Թsi!D�0��IH�f�|h�nV��K�� D�h9��ϝ{�|�e�7G�-x�h>D��)7/NG�٪�L��=㜰KB�?D�Pu	"^l�r�[�@�$%)O=T�01T�ݡr�yzG� ��S�"O�\���>�9����8��P��"O&P�I�qND�w�
�D��Ū"O���U�Q�p>����ݗ= �hZF"O�X�	��rn�+5��=A��uCB"OQC�!��=���k�֯�P�Q6"O�l3��ϻe(HP��@�A"O�=D��?9>��7�&M���J�"O�y	�2[��)�����$�Bp"Ob�뢋��4c`�h ��
ڤ�"O���b��F�"td��+ڜ �"O"����Y������U���i�"OI���O�u�����Evh�R"OB�c�@�Y]�`�c�@�k@tB�"O<�:�C\�j���j���"O*���[3��E���G�բQ"O&Q&�+xI�L�3J�$��}�U"OBISp�XJ: �g��3NSd(�C"O&�8����T�Vd�t���9z+"O$����^�|��l���@�-�8"O��AV��!?�kF�kL^-)�"O� ��`ɼY)Dyh,C�??b�c6"O�ia�X�;&q*8@;�ؑu"O0(:���z��q�30�h��"O�(x�b0D��lX��J9q����ēn��2b�&�3��Сf8�ě$�X� �怊�T5k$���Q1�������$�F�@Eg> ���@�	ZSL	
�T�0Cf�Z	�-�C#��(��㉓n4�4H���I�ub&� $O43�(���'����C�I-1���c��)���
G@Q�;#��'[ ͙����:V��� ���%K�jj$��O�_���/��hJߓ�J�2�kG9���	nP�i�|M[`��j�$ݢ:�v�ڎ��Ӻ�3e�O��
���@�f)c��#Y�py�
OX��E[6_(XYq畊vL4�⣝*XY�E������8�4d�������0���^�ǥ��)DS8P��jC���>��O�x��d(NR��y&%�Mޤ"�i�ACE�Y$��O?7�;h응!�̜Pm��w���1�!�� |�-[q�d��p �օw*�ɺD8s�3)u�y�7K�R���A�(�� <����I+��]������ `�*b��/��@�E�\�*�ڥ+�.4�Hq�/h#�0Q4�P0��J�9�w$����q��?�x"�J#X��1��BS���Q���5D�Љփ��&��գF) �Z��0$t�����68{��+K�"~nZaɰx��-�>D�����(zC䉬Q�R�)��%T+F��2G�����`����&��Y���D�G� �����(q��_-E^a}�Bɏ>B,i�2�28y"a[+"o�UȦ�Ыd.� ��yt+2���>
�T!� �D<Ez"Xr4Z��Uo��y>pʒ�4$
�Z2�"y�4a��U�=�iě/����C(*8� enڍ���{�)���S��M��i �*ʴd;ׁ�Q�p��@y�<�f� Kg��I�����[CGuy�+M�"�=�1�'lY���L�u��5�ć��D}3�'r�]�G�������S<{b9��':I�R/�mV	aF��L$��'��1S�-wa��$A-����'�`�k���(c�
�	 -��~�bYQ�'_J	{�:3>l��F�1sP��	�'?0�5��$L �`�c$I+Y\��#�'���w N����	Ƌ�K�&�!	�':t��L) �:\�0��Fʲ��''��ЈʿT�D���G�8>ؼ�'��X�(ݱ��e��81>P�+�')2u)5��*�.���:�V�"�'n��uE-)0zPK�90����'��L��'���H�)1�*3�Ă�'Nv!����^�@Mt ��*��ܫ�T[=���>����;�����Ɣ8���%x�<Qt��p^9���"R.y�h�^�-�,�A4B.�	�B#��?��� V�'[�0,�"O�m�n�+��+��^���X��$�qOHÎ�Y����B�K��@7�M�"�Ѷ�&D��1WP�!%T=���K�zƂ܉d�w=�X�B4�O��q���4���f�]Wٶ� 3�'�|��`*:?	�BV@"9�%�O� �,�P��yR@D���f�S�t��x�Ѐ��y"���
� Pb�	d�::p����y��ǵ8�iYE�(tq�Y5OH�B䉩$(	���}��jZ��z"�-D��Q�kĹT�\�Ƞ �A_�y
")D���+\�#�����fZcAJ�+$`3D��#�F]� �.i(� #~2��/0D�XiRl�v2�5�gd
�0�j���)D����+TaNi�FN4yp|e(D�1T�T�KB�M����+n|Fd3s�%D��bG�`2,��C���Z@�7D��2�_�-��<#�BBT,���*D��yF$�6:���lוi�Zi�`N>D����;�j8
P�$X����%?D���pD�i�z��� �,{Ѽs�n9D���#��$N�`]�̜�nsT�x�!9D���RÊ�L�}���v��B�2D����C��ME��Ђ�N]2�0D�d�D�����(i�V�5��҄�-D��#e� mmn�<A����G�Xj!�䎰�X�qp��(MĻ��"Hi!��_�Jw�rq��12�2�S!�V��=j� W3��J��ɂ:W!�D0�v��C� /Lԉ�3B�<!�$_�%�� �́>G�Qbb�X/GD!�ď0OP$�`G@�a5MK��:D!�D�gp�<�R�hʆ<3���3]!�wT��f��� zd��>!�� ��"ؾ(9&�ْE
W\�uh�"Ox��$*�'qL$�"d�Pݳu"Otp2S��^��C@b�#l�h!�"Ot��d��gLb<���N#e>��Y�"O\b���4�&F�)�!X�"OL�[Tĉf҂�s�A�h!����"O:��� x��� %O)q	����"O)�r���IQ��V2��6"O�� 0
��O|4%�aƜ)m��D"O$��aE�<j�X��oŮ|��"OrQ��K2#�����U�$����T"O��)�C��(3��#���Є"O޹�$j.��@�!X�"��"O0��.]�>'�5 s. +e��"O
���&W�Fؖ�yn��]RR���"O��z��Z��:���b��*H�1�"O�0���J�v��jG�;:�j�`�"O�<h��R%xX	æS��R��"Ov��@��.ᚗ=�
�P�/��yr��t��؀c�E�>�jP�l�/�y��£<������9�����(I��y�@�|�TU���ޜ4έ�q���yRĚ���pĄϨ)�ݙ��yb� 4j���9��8 g��y�b_�I���ۘ��!���yҭ�C� X�D,Q�}��E���;�y2B"#�����;|9��	P����yB��
4*r�q��-{�<����y�۹H��	�R��w1�Y���Y�yR��7{��ت�k	�~>���.�/�yR,�>N��<�h�x!L�_��y2=ft�EBF�<N<i3$O��y�@�75�� ��-	�8z�<sbK<�ybhL3d&4�0EU/)�B�c�@��y�C͍x�� ��%�*1$K<�yR��N��h��H�M5���cș�y��ǋ:z��4*D�<���ڲ'_��yR	�+56�3R�>��j����y��yҹ�BΊaL�TX�j@���>Q�O>��G���-7����j�P~�7"O��
¡�2Fl�*
16�})"O����g�i�chA0־��"O��Qc�.(�x���
* �*+U"Of�g�Ag���nߐl��M�"OrU��h�
�$��GmC&*��i�a"O��ң�V�v�J����00��"O 13�⁾L�z����91�Yy�"OJ�"v�*��P B��R���"O�%�5�պ!�D���24��I��"O,`:��[/��▊����"Oޝ���v"~ Ȣ腍^�z�"O(����$˒��0>�ڽ�"O�k��[vӞ̚c�G8{����"O 	Au���D�b��ؠxs�=#"O��Sb���9>���H>[­s�"O�T�c�Z�k@��RĈ�"FhP+�"Oʝ�%�b�� &J؟<��"O`��E�Ǝ,��qbɛ�rמ0c�"O6�͒5u2�B���V�̭#�"O8J���"�V�Ѡ�:���p�"OVb�ߠmgؽZ@�S2o�rm*�"O��'��8�zъ��ͻ{�is�'�j���89�(yAOS�1GL9!Fς�>��B�:�0C OI�?�xع�I�:\�`�>��3� �ձ�Ǟ�~G���т\'!�ؐ�"O��"rA-l ���a�.r��Aq��O��Fz��Iݮa�~����>�.6�9>c�B䉇zd�tp*T�]��a��
Đ<3:�'����$�;,X��c( ��f���A#89!��ۚ@��Ŋ��S�)���3ã��!�$V�v��p�d
g����p��3a�!�5	��r�.�`y�a�!��D�.iZ�+�#}���y�G�.T�!��,r&�d�0��>M�}��f��!�Ă�k�"�3D��<���e�\/\�!�D�$�(�J��X�_�,��kC��!�Dԏi<��a�b]�e&���A�!�d1KP��
S�%H�j8@ Kǰa�!�Dو"p���#,+<&9`L�Am!򤐶u'�8�,�J6�;�@ĶBX!���hD�E�l̮[�)E�VY=!��OLi�v��2����
?!��UO��A3�N"�� ��M\1c!�dO84U�1;�	�5��PcQ�N�P�!���C��ȗ��`��Y�*�3�!�.h�Zū�Q�N�u�T'�,%�!��\�3#���tK��!�%���!�!��,yJAv�fE�D��gg!�Dӹ;aJescn�5�F@07��8f!�D\�"��-ǔbJx�!c���'vў�>�J���?wi�+�#)(�2 �7C0D��kG$[�P�|�h@��,u�$�rƦ-D��Y�.��3���&��c��B1D*D� A&�W��Yҏ]$*:����L&D��U�Ooʰ��G\+R|���1D����S�pSМ(Nۮ�}��$D��[�MόT��Љ *X�oQ*�P�i5D��p�O@/Z�b��4�$$���G9D��2��4K�*����!W�h�$5D��a@�)��}Q�P�hb��Ȣ�2D�P�Vc�+DO(Hq�
���Bq�$D���f.F��h-f�����G$D���r��%�� �Jr��	��.D�yQD��q����t�y�a���+D�I���.����ꕛ0�L�R�G,D����f�J��a�Ғj���m)D���U�Q�*Րs�N�Vz�}r��(D�`SG��F촹�0[�M*rB*D��!��\:�ęa ��x�3�'D��W!˹N��As�ܚ��ęd�%D� @���0��9S�5�����%D�0� I�(5��A��H�:X���>D���5&£
Va����U�Vg'D��'��K_�2�i#�M�3`&D�LJ!:	M����	�=�դ"D���D��!$��yw�V7	=��cI"D�c$�b*Dp[$gV$�h��?D�xH�c��tDzD)�M��-�z� ?D���&*�,RY�*��@�}bL��q�9D��3R�V:��_J*p�p�6D��Sđ�5\����A�]�Da��-5D�Ԑ�G�5k�V�!���_�0�7*4D��s�����܌�P��/�M��7D���A�ѶT��`�m��~3�kU!D�IǤ��|4�Ɗ�+_&��`�� D�؃��ޑZ>8� �/Wܴi7g D������ �9QD��=o�׮*D�@�tC�7���[�%�� *F��g,,D�� �K��R'KQ*Q�%��$A��pr"O��n�	D�l!�!�2[�H<T"OZ�2UI�H�v�H�3B�r�0"OP� ��%*�z��R�M�  `"O ��Jd�f��� ��v <�5"OLe�k��,&�}(���xe"O��*H�m�mA]��9c�%D�x"ÈL�b`� �aS���P�G#D�lD(ԉHQ�����G�T�;�"D��+� u>.���m�r�BDR��2D���3�ςv7�M�A�T>� \��k+D��Kw�W����G0F��p�6D���G&U/Vd"ՑuB�y���q�f4D��IUg�'q�L�a�\������6���5^)��E̍>~�D5�J�v�VC�	9�h��B(#6�p��B@C䉯a�k`	U8:�̓�oڃ3�.C�� h�xjC��!��x�aQ"c� E{����!:v�*��]z`�!U��yr�	/h�1B�f��M�L��e���y�O�Dvj�Zp�T"?��|s��ި�yB��9pJ���e�?h[l\)�Dǖ�y2�Zl����B?S���Xj���y��u� �m�8������o�<y�����L+P��=<��B�)KJ?)�!&j��$�E+r���Gٿ��q�ȓT5����+�=]Ĭ��B�ܲ}����E�pl�$�1c�N4�&
N��)=D����	ƙLj��h�5��7g<D�,���\�=�R5���f��QV�:D��xq(��%/���&%X.�T�*p(=D�9bnɧZ�X�9���+�C�,<D�P��ؔ ��i
��=I���&D�`
T���^�vy�P��a�.	[��)D��y��6K�B�iUZ.ZC��T�5D��JCOJ�5�FH��"<�4(�k?D�L2�Jߣo�4�+�R=X�!G� D�H�V��p���D�7�")Kf D��@3F��ɔ�@�ÔZ���g�*D�LPԨd��y��U)��hD�5D������+a��A�A�
Z)T���6D���F�^>v8��&RJ��`"�4D�<*�%ՏvTV઀H�=b��S	3D�`��ʎ�59�-Іk�,(�j�0!3D��ᅭg"�����WJUy7n;D�xiƇ�?Xi�G䞍q�*�QsF4D�|�c�W�j�Z��֯\<c��z��<D�\��	Z�!.Y���,?�yC�/D����	P�m1|���.�3Ī���.D�p�LF�7��l�S�ӡ:���[f�*D�Pp�JP��KѪ�`��KJ3D�țRN�Es����ֺ2�}�ԃ$D�ܫ2b0NYr�ˤ�m j��f#D���2�NY���є�Y(��%�wd!D���E� T&�ӧ�U2�0�p�$D�ܡu�[D�LH�bR�xMn8���"D��%J*��Ԫ�H5R{8\�tK>D��8� D�W�� 8c��K�hi���1D�( Ƙ��č�$�\7g"���'g<D��A�LfĘ�0���w�(��8D� R���5{b���O*A1�<�7D�����O�Y�Z���',�|����5D��01GŞ07�Y�t��bop��@5D��"jQ���H�G�5AH��uj1D�� �@	���ln ��ED�Z� �Z�"O�����j��ڋG���K�"OF�R���>@M�@�̀�M�.a��"Oz ��A[�PK^)��KՊpx�aa"O�"�+/���`֪>/yp��"Odp�rK��Hi��J	 ^��8�"OB��Pd"�MK"Ƀ�S}��"OTW'�&f0x�����3e�#�"O�8�)J0?�� ��nR�SO�"O��
��2 u���w.�/`�D	�"O$��Vˍ�(�1��욓Ef�q�'"OF�	�럡D�M`�aQ�`���"O8��3���G�<I���E�<�j$C�"OЄ���øl�8�I'i*K� !��"O:�-�T�Iq��a��q � �7�!�T�� M���Uu�X&JJ'�!�_����O�Hb̌���A&!�	G'N�úI����N3U��C�	�Z7b�b�O�P�x|���ı]��B�I6D���G��(��|3@Ĝ:b�|B�I�oyp�P#
�	y|^L�G뜝mN�C�	0��D�o�EF���ފ�4B�	:?�N��*�;~L�i�۳�XB�I�\�ҤӰ �"~~��eצ:��C�	�z�����=*��`�]��C��+j���%ȍ3�"����G)i� C�I�/�%� �]U�R��ĉ&�C�I�-��|J�Ά4*w.1�TjC�-�~C�	�1o�R�?|��FFL4J�rC�I�V.����\�s�y�C.L(#�lC�	�yq"̩$�Ѝ^\(�x��K�Kg.C�ɍt�L4KY�d�E�ͅ�)�2B䉣0�5�7�	�XL���(Z+�C�9fe<!c��ܳcx\x2Т��FB�/�̙��B�r�4�S�M^�ZC8B�	 E�$��$+�8}����\,NgB�I�u5H��'�]0���GkJ�B䉬C�x`s%_�YF�Zsi�n�B�ɤz��8��Ƚ1뜥9���:%&C�	6+�q��AM1B�x����/]C�ɭJbH�����$�j!�b���C�	�c�r|��ޗ@�l�V%���C䉵�6�H#OƁ2�F%��TXhC�I�nt@x��J6L3~5�Ոܝ8DC�1�z!�B��Jex-��I�6H�B�	)G�������a
�X�!G��b��C�,,d[���0���[�B_pn�C�	Xڦu���7F}^0dJ�]~�B�4>ؖ�hq��T����3��B�ɦB�´�3�C2��9H�E h*�B�	��nx�b��3:��
qg�+�C��0
j}@D"n+b�Sp���G��C�	L�b��@�N �(�JQNC+��C�T�Y#K+�)0�����C�	�KzvH���,;�̐q��iR�C䉕I�p����� >�ƀ3�W�~|C�I#c��H� 	�L��X�f��&B��$~��ۀh�iΐ��2��j�(C�I
x��aT�s=V��-*t4B��sж���k���!JG�ٚ>w,B䉗0�<�� ���.��@���0=��C�Ih}�b�(���` œ>(�B� o��d9� ��ZVt��a�R.hFB�ɜ_�Zh��L%g�
�Г*ϭ�B�)� �!a�Dy�NH��'ɢ4b��G"O~L��B�*{�n8+��CE�颂"Or��5�͢e���if�W���0"O\��,^�Kl�lJ�~5�@r&D�CՏ��b�(�
E������aK.D��Q�,��OxM��bC>+��f+D����c�w��!���YN$���#D��#��P Y�u#���$U�&���'D�8Z@�ƅ%�H�¤��{p`�@a)D��փͷ$Š��m�w�DxA�$D���hB��ɻ������p	p�!D�������%��d�i��|'j!D�$v��/�:�C��H�x�!��)D�D��ʬ����%}f}��#Q�ylO7NO��;#�������ѫ�y��Z"yx�ف�AW�NQ��*C��y�Fh0����T�`u�%꣉�y��*阝��iR�	�2� sM��yR��$�zӧV�0��ah�2�y�Ȍ\��򷅓	|�$`A�"���y�&��N���!J�%D��Th����yR����i&'��f���Pc��y2 ��B�.Xk��\�*����,�y���
?7T�:n�%7�ز��ϋ�yB�E�=S��[q�����2'B�)�y�#&?�-�LM�W�i����8�y��W�r-�y��l@1N�@m �F	�y��.
�}q��S4Dh��xF�Y*�y�FU=f���C�9RE�f$^�y�V�.s�=h�d�3��0�d�0�y���h�a+��ʞ��A�v���y�A�@b�i���6q��P�6Q��y"@� }@	���9l����e��y"���1&;Gve���ǽW��j�'s���S��}H�H����c�*���'�0]�3��Y�RHٵd�W(���'�����гf^��z��B�H�`���'�,� W&	�J*Qc�&H��<a�'��	�&x�  �r�(?��%��'y8��dh�$O0����Э6I`�0�'�B����:5����H��C�
u+�' ��[D�[�i�9�'�:��qh�'�nL�VΔA�䥢d��-/�y�
�'i�ѫ�.�Z$<e�s���N��P��'t�PrMI��_�0�y��"O.�:�*�>�ӡ�3h���q�"OIiEN	�f��;�eϤm��L5"O���COȳ&˴�8T���J|�Ā'*Od���NyDM0Ԩ\0�r`	�'�x��M��NH-iC�Y�D��'���b��ZW;�BeU@��'����n_ G��A�c�Z�~�8�'8-r3J_�q.�HQ�oN�Q���z�'�f���
 ')������\�@��'`
��WO$lOF�{�F�L=��'�d����5&Q(A��	I2D��'< �!��P6�X���>9\�ђ	�'Q�雵��8� m��	�/0np��'x�
����_���&�KK*���'��URE���Țl"S�܅"����'��\@�2TЩ����F�䅱�':b�wd
E��cghZ�i�IJ�'��eCM�
}ʦ���0ZYz�'����e"C�d�u��. �y2��� ��h���4[b����N <v�ij"OL��$�(2��a��H�L���$"O$���جE�܈����b�c��|>�#@���eא�!���
7�R���Oң=E�Į�$y`��-!
��5FF��!��(>��'��+L��X�!�U��|��'`��6K��HzPC�kɱ�@�C�'�b�#3��\��x�l��#>��H�'���G�%"�H������@�)	�'����RgQ�B^�ɃΉH�����'��Y9���(������knJ� 	�'�4ۑ�V�T?ҩ�6"��0�d0���y���b��8ڄ��.r��j"b����>��O��)�⊐�b����ۤI|�"O�m�e��}�X��פ�pI�h!"O��cvk/~�j)ZQf��@C���"Ou�j� 
Vd�QET#)>6)R�"Oe�$����ˀ)�"YF�z�"O��2�C�T�tY6�8V)��9"O6 ���k,�����*?���3"O|� N�B�����
��\P���C��h&#�U������:z�* ru�>D����v:�����XdҬ�:��)D��!��Ǩ}nt�hf��a���ZUi)D�̑���9��|�Ò�{�М��.�<�	�p�2H�����'�FN0D̄ȓYq�R��	,<�j�E��p% ��?)
ӓ\Tb;��7h�҈1�!P�V�ȓN���Х�-Fu���( �ȓvPt)C��*aK�9FѬ�لȓ:��y�:yt���Y�q�xԄ�3����ٿ��b�%�U�ơ��q�����<���ƒ�x	&��i]��s��'���X ���/�^a�ȓXe��b0�R�y� ��X;���'�a~�%ME*Ai�7��qag,R2�y�`3Cc�:����yj�X 礊,�y��wb|�ĉ�Bꥀ�ُ�y�BD#��]�ъ�*WB񦈞��y�	��4�x�J	=mx�7�I��yRmVo�ԉja���&�H' %��>��O��zwe7��uۡ�#o�j�p��'ў"~���L(�:���P-�����yRc���Д�^�|�P7*
,�y2�y�U��goָ��ő��yr�`~��A�͖�@��F�4�y�e�y�u���P�?���;elą�y���1�ę��G�<�X�$�E�?����}�����5v��¥�L.P��i[�����j,C�iH�9�F8�ȓN �IF�*G���XVKڬj�VD��x��D�ݑ-j<�p�a��ID�0���{~b��-�j#���	����ǹ�?Q���1�4*���+`.@9�"iA�)$D�����}�q1����6��P`$D�4�&ٴIz1ɲc��Z��!�C%4�\��q�ɕF��r1�E)h!��Ɉ���fI��h��V�+H!�?<:�L�2��	P�}�Q,A�_>!�ۙ^>��MT�*I���nړk��')"�$)�ɅK�� �C��>B>�൅�|�f�?���鞎y��4��Uf0�%��	��ў���-�6���.�&Ғex��T�#{�B�c�$T�6�
wB1�`���\@PB�)� f�j��}��hᲩI�a,�`�@"O�s�� ��P
v���RLۓ"O6��0�<V3&����%kܺ���"OV�����:� ���d;i�4%���}�Ox���G�(>f�#�cܡ[{�,����M�Hl�'
�MI��i�j�:�!��W.�2�.-M�pTҳ"ԛi!�(P����P��U��>A����Tg�����E:�,ɐMµ���2XD& �X2<�Kk 4���Id�֜���&4���Z�DK�H)t�%�����?M������Ο7�<y
 ���">rB�ɆZ�۹&
��*<N�ᦔ.&���=���V��Ai
Y���BL�.��ȓN��i�A�OBXM9ËH�C.������7a�.X��Ph�デ&�썆��I~�)+G��H�#�`���V!�hO��D��D���c�IƎHyGD� ��O��=�O�J4Ic�$+�Х��L�-g^��Q"O,X�'��?k\Z4�����<�2X�l��I
 ��2�Ċo���@��1�@C�ɑ4l�i�����d�@LރoE�B�I	h�����TJWdu�sϝ�9kC�ɂE�����,X.#�T����f�=Q�|��)Ӆ�ЇJ���	T��9Ix��?y���~Jw��2t��Ѱ�I J���s$��|�<qhM�,�ň��i�PPŢw�<�pM^�]2�(�6t���Eu�<)���91`��"�H6b�̘���]z�<Q�g 'W0�Y���ȵ;Z��c'^@�<Q`E@-,����DO�.�N��ւ@�<q���b%d�s!Ū6�~D���Ey2�|��4���4x�H��֌L�U��D�ŇP:1�!��G7O����˫@ܘ�G�&�!�#+�k�Í�o�:��g�Y�D�!��H]��!FW�!�a�լ"�!�V�k�2����W�|�򉲆	B0%}!�d��!r�M6�5�`�#�T�K�!��6`�H�'�ֽ[��kH�l�!�D�*=�lQ cR�,�d
�'�L��'#a|G�Wl\X�$�9���	f��y"��ʼ�@���Ǧ1`���y��sDzH��A���tqWƃ �ybb�Hʞ�Y,�%s��RW����ybI�Z6�a҇!L��vΜ���$�OL⟢|ʣ`)h����Ì��a;����p�<�vf��$VPJ���S�!Bk�m�<��M![�`�@� S�\�{0�^g�<	v��w>��k��Ɠl�,�;�d�a�<Q7��;ho*Ly%�i�e�G��f�<�B�3}#V(2�l�0�4�z��h�<4���B2��hgL�r]����hOQ>�)W/��m&�A�2��O�4h&� D�Ԋ3���&�� zG<Aw3D�T�"$_�����2k�	V���q�1D���+�a�b���$�5�%�T$.D�l��-?E.t�"A�kk�Ղ��/D��C%gޞ-FX3���
$	�� �,D������*N2���tm�'j�r�¨<���?�N>E���A ��0Λ�df�B��W��y�E�4%��u҈X�h�h�����hOq��pIg�CNf `o�G�e��IZ>�:�$��p�:��u�i� a?D�(��[�I��D燦<��D+>D�� d�uCY�n�|�SÓ/ /�9���'��/a� T  J�"a���bQ-[�!��L�*ձf#��1[�j�"p!�[�BTP�"Ō϶v��B��$ZўP�ᓛfqz=#�A�p�X��Q�W�crʓ�䓩hO�i�{�aȶj��r����e�Y/)!�D��a��Ƞ˂
?���kH)!�$I�He�Qc�5KI�Y����!�d�!f�A�ƃ%3�e�֨AZ�!�dJ�Sf:AK�]�}�j��ب;q!�d^	;A\8PB(K�n�9j%��nx!�d�(c&��K�'�>��хZ�[i!�č�N���F�8��0�cf�#md!�$,~y��ܻq�:2W��2V�!��J���q���t�Ш `�	@�!�$.JN��RgD�*{x�b��(O!�Dՙ]��2'��<\�`�B1N�7���H����dԲq�x����<���h�l��2�!�dG,�T	AG�?=���l�14�!�����]0ыF+?����6Em�!�$��'xy���1cސJ��V9!�!�$�[%*e $N��#T8�4V�!���%h�`E�OE��07��5�!�dR�h�<�D�Fa�*E��[^�!��F�) L-Z���1�(�:*!4!�Ă�G���`�KW�!A���w���c!�ڶ���Ƞ�̐(;z8#�k��!�Ě�i����q` �F��	�vEN:�!���Ts�|crj�j\D���J���y"�'1O�4� Aȝr�A@	Y%��[�"O�3!�Y:��C Z�I�"O����U�~�.M0�!�f�ۑ"O@D�V*�KND�X�T�HlU"O�q0��L&"��c�B�U�>=�!"O��3��	>|l�4Q]�s϶�"�"O�q�E�1B���`�C�/�&��7"OT�1�ȁ�1����R2{ p�H�"O��j�� �`��<'HR1ho��w"O���c��+���b3�˗I�>���"O��e�+֌��䫋�+B���"O�D��ɯ4֘e�kT"0��xu"O
�:��\�Gָ]+1
+��E�"O����;G�v �fI�1�n̸�"OȠKe��B �J`��07l��Q"O^��g@��v��1AdpyS"O��"�L�9��x�g�vf�<����&LOL�Ru>�v�� ���4���0�"OI#Î޳=IH��"Um~�8q�"O4DQ�k �Oy�$��ג)t~A"O����ބ����jj�ѹ�"O �S�
	��t@�F�Rw2��1"O� �P��!v��*����9�����'h�+�U�æ�C�
��.`!�P�����/D1E�n(9BNS
8!�\�YC�32��*�����H�%�!��;]���V��'	����v��#�!�dݢRmHXPN��3���,�-y8!��;���#�	T[Ѩ�+QIβa�!�M/<�%���6h]�M9���t�!��S���iG(C�2M�L0!Z�n�!�$�31x�t����q<��j��ۀ4V!�d�!(Q��C�ͮ��	(�%_��!�@�f?d2Ҫ�!|�wd� }�!�D[�8Ј�)5�����c��9\!!�� �@u��g�a��A��C;�@aE"O@��f��2�ѻ���0u0,4��"O"�XvH܉S1�ȸ���< �t{�"OV��T�4m��@J#H���G*O��Q�H�8�D(��A�#hl%j	�'��� ��5�f)!7��vQb�i	�'��8Gf�%ShX��&��h��Ě�'��x1�,H���r���`� 3�'R��s�dD�'�f�c �&�Ș�'ӖC"lI4"���kt��=hR�m+	�'[����
1C���D�7h�p=�	�'}�,1��ԅ|@wƈY�tU�
�'q�ԈǇ_6���U"�"��y��'S�][łD
F�MɆ�
!�289�'V�<s"��g�tI&�	,cL>8�'πE�D�I�]3DER$H5^5��{�'iT�����Tx4@ġ��W�&�K�'���Ǳ'�<P����8ya�'Խs6n�=����c��ҭ��'�z0�HP��J=+p�%��,j�'u�5�N6#3B�`�B��`91	�')>q+�� 
����h��=*�+	�'`��jwH�#W@��W� � ��ܓ	�'s$p�\/z���gm�?-!���'��(G��UЪ�C'c]@��'2�Y�"��;V8����FOD ��'�h���Y�`�� (V�;|8���'�։�0����d�u�+H��@��'������Ţ(�����=9qP"�' D��D�9W�:DP�(ǎf��2
�'�"�j�o�r� PM��WH���'����D�٘`	��bϽ�t���'}2�Beށcf�:�C+����'T�U�k�x���#��Ѣt�~P
�'�B���O���8����N�ovnHY�'�����kL�y���35��0k
�'�����̊,}��ɒ�W1E� ��'�B���)_�q�H�Pq
�O ���'��)�e��Я̂zʐ��Ɂs�<w��>d6��P��>)�`���I�k�<Y0��W�,)����^ :	b��M�<a���a����ώ#%�d�NH�<�ңF�O5��K� F�! �L�<i�N�;n֔�!T>��j�F�<�a��x�n<�r�I�kT !a�E�<��OP�R���z�J�0(x�CŤC�<Qg�M���ŀD�T�p���X�<1�+1}���k����X@�^Q�<i�:����ү��0����
L�<��۠]�c��F/*[�h���C�<�D<U;J$��	R�v���z`S�'�?��e�֎G��$[�,N�y�'(D�L�a�.�	ig
K�E�$�Po&D�H V��-RЦ�0d�J�C�ԕ*�+#D���d�ܴ.($��'>�r��u�?D����IN�s�}��C"o��P>D�(TdO�kS�ŠLC�n�H`	p-&D��k��E
}x��r�ͰD��b�k9D��r�a��g\�HRk؛	"�Y�3�)D�HzU��$i����DEׄDF�q�k5D��:��G�L؆ �B���,1D�L���J2oP��G �X���yъ-D�4�$ŷ����1d\�;k�`1�C*D�l���J��Qʃd��H��3D�� ��&`�^V�1����"l�e�"O��Y�E�+k����J��fM2�"O�� p��=V�z�HrK� q<��5"O��y�i05���& X�jl4�`"O�"f�Vn�p�(
P��r�"O�(�GD+\���#��@�j�ph�"O�����">���:B	��H�3"OԵ+�a�**Q,�����z���"O:=�A%ٕ^�Bx�G@<<��]��"O^� V�I�k��#�Y�4�B�"O� �S@B?���p��k��1�"O4���>"�PX	�/�;i(T���"O�M����'��M+�+V.	6&p3�"OL��$s��B5@U�^��aȒ"O���w�`��Xj�Z�6���R"Ob�r�[9���/5��M0�"O��Cc�&vwN��P2;��4"Opu���F%p�BƱ_�v"O�A��ʇ�'�V�`��'<L)j�"O<U/�^�\� �%(^�*�"O��7�Gwސ��ỊF��P"O�Š��7I�����.�<����"O�Y�F@9X9�D���d���"O��� ��>��tؖ�D@ΰ�"O\� ��<G���;P�J&}�b)�"Ov<�&�@���h��ȡ"O�u���*;�����/4خub�"O	�4#�4`L�8�)�T�v���"OXI�U,�nMq�D{�H�O܁)C!��PhK�(�Ѯ�j2=D�4��� 3����OՊU6'>D�8���E�#��T	�G�L&��E-?D���A�3E9>�{�($^�H	2�:D��yv:|$9cҮ�BTޤVj5D�܋fE�T��8jO�$)�䩛�'1D� S�/��׎h9�.���I:�O��I�.`⩹�]� o�U҆�B��˓�?��+f"p��
8pHJād�Y�J����Z�|�'(�[`�ɹ�.�=Qę�ȓ\Т4I�R�8M:%�S��sh9�ȓV��q��J>J&0<�/V�}�Ņȓgð��D`��>f���ӯ^3d�l��~��a�	���ߪ�4��ȓi��Ywh��~i �ٵ���A��ȓ$�YDئ&�v�	PI�"a�>�ȓ~����n��� 	��҈��`��Y�ƹ�1Kl�z��,�	�*݇ȓo��B�c}�����ꨇȓs�� ��"�\��c K #���������C��R;�m��ƚ�yF�I��RT�Q��P"O�A��F+r?�%�ȓb{L�� <�G	��(�$��-��Ty�ʒ�Lv���*��x����-e���D�-���Bq(_ 'BLh�ȓv<N� H��o�P!���ҁvZ���c,��2�C��zN̈ g��X}���ȓgI3�
ì>[���	�|+:4$�D{��t˙~q�9�H�����[㋜��yBcе^q�c��hȨ"%��y�����wfC���2BP��y2iA�14q򬅮M�4JQ��,�y"�"B���Ό>o*���@��y�T�~z�)B/��@4B4�pI���yb,�p���4G��=P���7a�2�y
� �(��
�@�����g9�X��"O�Xk���/o�4@	�[�eq���&"OHH�i )PY0Q��Y�eR���"O�G�O�r��g�B&M-����"O���U�	<��p�i�� *8�#"O��pu�u�US�h\�h��0�"OP��aƤH���HF���"�"Oh}�VFRh�]�w�ьu{4�1"O���5H̡o|b����_m�� f"OΉz�A���`� $d}���B"O� rfU<(Y =2ǥB)&� 媵"O�H��J�'����H-/iV��"OZH�J��J�* 듣�d�� !��'R��'f�dL/!@�h�	l#�*��&�>d�ȓ"T�rvD��=�܍ڃ�ی'����''a~�Ϝ4nd���>O_����*I&�yn�EHpٶI@'L�LDk��/�y��S�,�����1uz��p��5�ybB��?��M�����7G|K�a̜�yb%� �]��O��0��ra���=y(O���D�0W�T�"z��a	j�:C��&*�XE��H]D�I5�L	,m��O&��D�MW�0!'�L�o^J݉��ut!��_/e���#�f�X�(�C�n��B@!�t|�a3�̀{�9(͙�r!�dŗ�Āy�"��l$)�E_H�!��̄b�ۖD�8��0󦆝99�{��'�4Od���'�m�"(H����&�����"O� �ፐE~R�ȗ���|t��"O�E�$%�"wP g��>)�\M9$"OX�0�l��(�m����e�4"!"Od��D�cDx�X�)��.�ȉˤ"O��;��͘h^$��v��<�f�(c"O�����gh�pr��&��=��"O�]��m�+Y��4�= �"��""O ���cQ�2��KR�GgU��e"OZ%Zt_(Y��tC�R�ؐ&"O♊%ʴGiZ�b!E�b�p"O�y���E"b�0Q���"Ǟa�E"OD�#ڬm��Q�%R�|��̹�"O�9yO�_���EɠR����"Oj�r�
چk��ɩ0�{VA҆"O��pW�� $�:(��%E	Ly�� �"O�H�*=�Z�s��KX���"Ob=
��:q�n��D2VGH\��'�$�a��,Qg���AC��"m�'x>�hTcZ�5t̘AdD�#��9q�'+�+)5i����1�R7}�K�'b���qoյؒA�%�(	�y)�'��-ԛ9I:��b�L�2����'⠡�ae�]��B����^�"�'	R�����<|O���Ɔ�"T���'�dH����;̐� �ZO<�Ճ�'�Pŉe�\��4: ��C��0�'���B��z��ӿ+>c�'���� ��d0�
�#�=	cr|�,OV��hO�'u�Q�2�D��P�(��ټ@�ȓ����$q��!���\����i��!C.��8��Չ�B���ȓG�4#�*��Yӵ)�5R��Q�ȓ5����p�dr�t������ɇ�R�0IDM�8-�,(��S0X D 
�'���[F#�j�֐:g�մ:�څ�"O���f�<CѶ���]�Kܔ-� "O� ��.Y'v��8��	V��5��"O�!C���B1�$(a	��W��MQ�"O��@�Dƀ<�}Ia��i�J��"OF�ڔ�\?&�X�bȷW�Ҍ��"O���Ѹn�V(��сFmnx(�O(ѻ"$fe2�̐-��\a�O"D�D��o�l5\��p,�i�,�p�O"D���!'ˎ�cv 6�L0�0o:D�<��A�{,��8dJG�0|[��#D�xٴB�4L_���;���ɔ�4D�|���R(Sҵ�1�ځ����t�.�O��6X�����Y������B��B��JYJ,�w�Th̶�3�f��_�R�?ш��њK
V��3X1G�%����.��'Xa|r��5��d��	z� ����y�#tIr��R��
"޽�B���y�+�:�N�����0�:Y���߀�y2 -J��T�"�ژ1��Y �5�yR�J(L�*Ts�AF.v�0T�'"�
�y���it��&f��5*Q?*kP��ȓx��jQFM�Q9�J�+�#��5��h����r����˔Q�A"U%Yt�кTo,D��qҭݐ � �SU��>C��丣�*D��1F+�m��|�%�A�-e찁�:D�\k��>�i�w�Y,ڀA�g5D����.�*\n�)�@��K�����B5�D<�SܧY�@@	�K(.>��J&���(�ȓav�+KS=.#��j� �W�.����\)�����KT#�sy8���x�P0��@��L��0�V��"I�ȓ��,���j�0���@�U^ ��w{�m��ja��3P�X� �N��ȓ�rAv�] F� �ƫ�&�����^����
��)a����)K^�L���	t�'�����F�`�2�Ư�����'�&�����i�yD�F�n�p��'c�1�R�-t/�9�'�<�"�A�']�):�픋cҀi��*8�����'8�ja��%����s�)R�|
�'+R���H�S2����f@,I��"O8��c-˞vt'ڪD`��"Od�i���n�xha�fCV8�IQT"O>����iH x(��-|�r"O+�F-Lmb����6E�Գc"O\T$�ml��R���`���"O &ݵ]�A{5���;�O�,���ۺ�!�hZ�IД=Qt�0ړ�0|���X%/p>�{f�ȴ,��<��_g�<������u�Y�1K��a�%ܟl��I[Fĸ�vA%Xxxj2AZ�^p|�ȓ(�(�
w+�a2%�Y{I�ȓ|^�1)D��chQ�ըN�]��ȓ7 ]��B"n�y2�ϥT{:x�ȓV:�j��Ĺx*���d
 a����E��9�ϲ-�"�"3@���T��ȓ@��$�ؤ7O60نc��Q�'�a~Ү��c�N���⏥qLވ3��y�+�w.�(��O_��i���V��yR�_4D�\�)�8i��nU��yb!�Dk�M��!Z�P�-�.�yR˗q���A��a覈
A��)��'haz"��~�( �A/Rی����hO��L#mO��p5	�t�cwCF�!�䊳SE�]+�悉r��d��B�f!�� lD�D�=�a#�?A�<�b"Otm�2@�-�%8�2����"OH���8=���w��9��)"O�	5j�ފ��	�b�;w�o�<�ю�� �ƴXë�>~��:��S�<�Q�V�U��h�1h�I�5	Fy�'�p�F;P2�|�5)�?`Ȝ ;��d;�'`� ��G�4+q�* L)�4���t�$Q��D���Eh�7�D�ȓ<J>�����p4Ys
ڐdA�1�ȓXrp���:#\d�SP�PZ��Յ�Ir̓J	y��/�9F�"W�ʃ08I��k����z�2@��#X'p����Ic<񐏌 �-h5��p��E��g�Y��Q���O��XY���tqD<jrت0�s
�'�*5� ��r��iBͺ'�Z��	�'!�}ɡ�?|� @�5��!h:�p	�'n@� ���6������q��'S����茑t ���F�U��@7j-D�(����b�L�w,G$r�v�б�>D�����\2W`�]p�'�p�f2wc�O��=E�t�҈�r1��W/D$�؅��`�!�D�G��)�c޸G}��1�j�!��%b��B1@��tA��C��!�d�8��+��s�!!��Xu!�d且�Rۖlf �r���t!�ċ&#���q�ɔ@��@`q�ځ
!�$_�Bg*���BÅ*�l�RAJ�*K�!�$Ă1�N��׫��+�XQB�i^�
!��S3����-�]�F����!�$J*��R��&xV����P�S�!��yx��ʿ#��1Alʿ�!�$S�t7<��/��@�8�R�hU��'�ў�>] !^.uwt���J����q�n#D��a4\�B7��(��V,���.D�Xh��q�PLH������ȗ�+D��C�&���P����j�1�6f+D���`���VE����(�:��#D�4�o��*�j�j�ctv<;�*O)�tc:���mԈ��4��_�8G{����3�kc��_D��F�^!�D�!�Lx����rF����E�R�ўh��8 �F��v���[v�!�\O:B��d��!�N�+P4	�G����C�(^(n�se�(3D:Y8��V2 ֜B�ɬr�����ˁOwH����PCpB�)@�regH"b�n5�Mδ.�6B�	%/��l�݊*�� �L�w���O>��dJ.�Z���D�M��@�G־D�]����	�;��9'����u����+)��C䉘r\����J΍ B����#(.��C�ɭ�]C�,T�B�:쒒F�w<�C䉍�T<KQ���[`]"A�C䉯��} �	�9�D�A����x�PE{J?�CG퐄`.�D����/C��E¶N2D� ����oh�HPU+�`Q���;D�$ҁjU9), x���2�fi��9D��{p�S9r��V�86�Y��7D�<�q���(��;��T�=za�s�7D��� T���R�6>���� D� �'D�RJ�[ϔ"]�v 02�:D�\�`O��P^���� f��C#<D�����x�2(���'rfb���O�C��E��������2t���*��B�)� ��ÀD�O	���w��v�`��"O�|Zf ��7*d	�c����A�"O�,;� kU:����������"O�H�A=c���r��(v�B�"O��e��+(p��(��L:�"O�A��	��6�%]�ʴ�G"O⭰�Q�R{�MB�#ȒS�Z!��"Oh8�C�ũ�$e�s#F�5��UY�"O�l��)!����a�8x�p!� "OV�{@̄�Ao��u�P�j �"O�uQWÕ�
�%qa�-��6O80���oSp�@�-�-f����D)D�A�L�=Oftxc�W#��W�$D���Qf�����ۇ#��q��Yx��.D��	�	��'�Z% �N�:B||���*D���PlB8U�>�ٷ�� �$ʗL6D�`��J�ua �I�vR|@�P�4D�T�v!�&
�� G�H���e2ړ�0|"UDH!�sVj�2zi�A�
	g�<�b�G-XPp�kE83�!�j�l�<2&D>� ]2��F�}�� ��Rt�<��ܢY�5�c�Sk$	$j�o�<Q�D�!�f}Ƈ�B#d�u��g�<yqL�i �h�fJь_��"�d�n�<�ᮜ�JK�СD�I���H�5��h�<��e�7v�9Q�.5젰+r�e�<I�Q6%��Z�O@/
\�[%��j�<!�l�q)����J��U���Zf�<q'==�`�X4�B���"g+_�<!(�7���i�C�&S�����ɔW�<a�KH(a*��A� H#����V�<!"<HrDy��ʞX��(�+EK�<��eR#5vX���-��4s���G�<��P=)z�����5zeZx��&�D�<�c�*:z3�Ɍi��H����\�<Y��D{$��QB��%o��{ċ�Z�<�@h/���TL
�o� ���o�<Q�=TYXq��V�dD�l��"�E�<1���J��-Q���U*�p�BiB�<�懖�~����+�h�&�Rc�<!� �F�^e�U��Y\�-��NXb�<���ژd����E�!�X(�fv�<��
V�(-x�%2P(@�G�<aC�¨utqZ��A�>���q���D�<i�!� n�b�Z7R~�}�r��\�<���3T|`��/6��a!LDV�<9B���8X̰��K���Y3��T�<ɢ��S<�f�D/	Tv����M�<�%�ރ4K |s�,/d���1B^T�<�2h�&S�٠�i'ԘP)C�l�<l�	t[���ti��.)tb_^�<��&>���WDlIY��Js�<(�Jh�pq�H�0����m�r�<ɑ�4���)Q7��Ua�
�k�<�d�֖@t���I����ƉX^�<�t���.Bд���+pL<�E6T�8��F�H�H Ku�$cÄE�l5D�z�&��*���dؙ-{r%I�a8D�<@@�b��+��W�T(~4s��"D���pF_�#�ƥK��2)��#�&?D�L!a���4�RnƽL��lx� D��Ä�<�b4�?+��,�Th:D�t:���	��!�C,��`%<D�䁵$��Ap(��*%�p4�c:D�� ���7�A�b��$�?,0t�3"O�U�q��L֡��$x��"Oz�*�]B�B�W���<��"O� �FW�N_.};�Ðb�8#"OBt8�OC�Spq�7�B�i`"Or���Q|�q�&���%s����"O�l��
O�r�f��K�&bhт�"Od�I/�"N�@h����6>�:D��"O&�0��\"%��c�+ӡ#�y�e"O��g���}��u���ߑg�>�A�"O���Ɔ��D��t��O�~p�L8�"O�Ջ�N<�x��#;	g�,��"Ozp���ږ
�T<��C^�k`�a�"O��0CR��
�o�Q%�!���8D�\ p �}�h�P
W O���9�I9D�X��J�=�`��P5ƨ�Fe8D�|:b�<!i��P��а|P��W�4D���2+"
�:dOpp4X�Ek.D�P[t��"�t�B̙4�4r�-T��2&��]9v�z��I* 8��"O"4����~��`� f`L��"O�QTH�(Վ	��BN�@Jx�k�"O��"�3�^�2���0����"O|4�U W($Wj��r��4	�v�ё"O(�`��X7xn�]7��z�� �"Or���Z�#0X�2�ҙ.j����"O��'F�cɚ��BN�Vz��0"Ob%��-Ҥ5&���ф�7V���yA"O* b��@�<��M�b{��;�"O�����+�H� .^��u�"OVA�2-� �6�2'\�}[f�*"O�x�#]�,u���&��'+\ �"O��V�R a�8�rE��0|n$�"O�x
f��pw�`�Gj´1�( P�"O���K[9C6��I'�<�J�3B"O�!i��X_n��:��$�����"O�%Q����6`Qq�V,b�����'H�J���Z'�t��ܚ伄ȓc��)��ǀd�MH�AǓ&��ȄȓG?|s����4� ��MPE� ��dF.5���MSh�#�iǸ&��ȓ8�Vy�r" �:���0.Ƹ%����ȓ��H7(<j�P	h�a�U똴�ȓ`�lػ_� �(@���ҳGNʹ��s�\,��
"bLT��Ԉ�b~н�ȓ$�z���C(e�$(�AI�C�ImhlQ�`��kR���4C�zf��ـÓ>��l�a G�Cn�B�	���9��%J8U�|(Q�GE&C��B�ɻ_��a�i�"gYɓBX�B�	y�]c7.L�G�mIW/B$B��-�`t��[�3\��HuA/�C䉭f����6KO�����9d�B�	�ALr[�^����e �D�8C�I�e�x�Kֳ2�ٵ�Ås�$C䉝(�Q�p��*> �/�� �FC�I���,9���NMv���l�5�TC䉜6�]�5o�!Ycb��t��FC�O�ъ ʖ.X*@�m)C��"x�b ֤͓J��i9Č�v�B䉵:h=&IN:'꠭w EY�C�)N�FI)���l�h�[R� �C䉧o=�%+$�9��E�~�C��(�^az�BJ j���9�Iا'�4B�)� �9
"'�N�>�`��FR��u"O���ݽ�t\9��^+p�	@�"O�踓�_�M�dy$Y�W�UZ�"O�4�F�#JS�i���Ăك
�'��T
���f<�p����U�.m2�'�Z�q�?W~�d�U��$�84�'��8x����N�H+
Fh�>\

�'�X8�A�Z��2�B�`a$��'�����g�'�j�1�G	F�։��'�t����xeP�Z7��<$8P�'7�T#GB,��	�� /fL�
�'�(h��թSϺ(@��I.,��!�'EΡj�䔹"��l*u原R�R�)�'�&��Qș\�LRg�ӅX�v�	�']`P3!#Ӡh .TAf�J&X���Q	�'�����˜9���a%�ĒSsy9	�'\�͢D!BMRq���*uyL=��'[6�"�J(,��$�`��w����'Lf���d\� ��C�ꉱE�he9�'38�;6瓫5��-�_p���f���y�Үe�����ܒy���ȱ�V�y����s�xi0'FZ�nQ��"�y��Œ#wƤ����<N!�D��ΰ�y� �s�~=��@؃&^��`�T	�y�ˍ�4�vYq�2�Vt"7��C�<���G�#�� �a�ӽ_{\���L�q�<��H��[�>t
���2}qh��@�w�<�� �8S^A�f�0!����q�<ɤ��Ryx
��A�g�iH@��G�<�կ�W���c6��+^���S�D�<$���\4��a�I�FUH"��|�<��^�b�B�{tL����u�<Y�08���@�-^��e�$�{�<I4�T��Ɖ��b0@( p�Tv�<�i�3'��@rnV���cv�<"��I�� �A/��V�Pr�<���TN���˥�Q�vL�4CT��k�<�u�L!!�.m�F�)2�$RΑ@�<!�(��@�$���B�l�LRT�{�<q]2hI��(�ga��T0�!�ܑM`��C�9:�p8��&шi�!�d�!vPz��G�5��4	�E#�!򤓑>e��K�fJ���BV)e!�DO,!�PJ��)D\�hb��=yS!�$N5+<�R�h��S��	�o>!�(>��s�;r
fDґ�7h8!�܂,��};��7�^�u�X�*!��ܑJ�4E��e0yd�D�u,�b!�$K-s���hG��_Z��a���,r�!�d��f�$P3PӃ:}ZǇ=$�!�$ݛ;Z�����ŀ��V��>�!�0V��4���ͣo���qE��!��۹p�$x U�q�v=0�þ1t!�D0Y0\խ��� � ��ӷef!�=H*�2䉆T����A<`!���Z5*L�A%	:r�`q �M9D]��hO�b���؁f|d�I��]bF��"O��b��E�Ơ��Ĉ*`M��ڇ"OV�)@�hw$��d��TD�J�ay��I�j��5Ęv���f�F)ӶC�	7I��J�A�;�V���jF`�OV�=�~R!�v��Cg�3p�T �MB����>iR�M5eW	+���lal4p�-�|�<�a��t,��S$E �?M��[�gHx�<� �= �� 2���HQ�Y��N�a�i���dۼD��9O��:��x����iV�!�$�<��'t�'u�VF'w�$�:��H�Sz����� �y"�3$���w�K�1�m��p<Y��?bƼj�˙:�B���)T�O�a~"�Iw?���ΜnG P�*�vɘj��[E�<���Wn}�T);�-�6��~�<)��8}�p�Ą{s��CU�Nb�<y0L�a"�c�R�1+T�vm���t����O��s���}����B]6C@�U"Ohq���t�İ�Os �a�R�Oz���=qƁV0̰��`��=:��˷�N8��!�-_m}�*O��0�I�&��c���$I��M��'t��J]/18�ݳTT��I�ʓ%|.�$ Ñ*��peLԩ~��nV������S�2�.!�6��P���&P��~r�韲�$��o�+`�< rș �!����E2C�ɐB�~<��h�%����P��@r.c�F{��d�غ#b鈗�'>�l)�"���ư?��'�X�⡨M&'$e9�K�0y�,A���'�lu��*_���2!��b���(��d�i�O�|���W�wØ��J �d���ng��Z����sC���O�r�x,$Dx��u���=�Gj��6��MI쑍G��q�p�s�<�$I�`dz}�*������l�D2�OJ�	�썐(s�L�W�\
|�"O�
!N�:95�!��hĊ0G�4�#"O��p�׎}Th���r3pa��"ŌǬD�[
�={�\<��Ț�"O�����JD(aIe&�V`z�"O�Pp#��r�(�*δ�b0Q�"OL��A�,l  F,�L ڔ��"O����_2
�����
]0��"OȤ꠪8.�4Q�c�!�� �"O0��zz�[��ؾv/�,؃O,�h�EC�"�.�A!ɑoR��V�<iօ�5T��YCNNK�&Q�Q�<٧LJ�J�܍z����@�Tȑ$�Q�<A��G��%!D��"��s`�W�<QT����T����JT�T��hIR�<Y��@�ZDцG�]�Xc7��S�<y��*q8�u���,~�~)[�QZ�<Q���t?F)�B��;�*=����K�<��J�"� T�b}�-ƾ|$!򄗸^c���'�W�f�ĉ�L���Py�ES7٘���A�%�>��f���yb��b� [�'*�ha�L�y2�8-�(a�j�	e0�1!iN(�y�B�(Ǝ�r���+J��30@�$�y��B�	�d:���;S���r#j�yRF 8���#���/��u�Bς�yrƆ�VK����<$�Ԡb*�yr�R	,;�@�Ө$% U0�O�y���_1���*
�~(;KA�y�kK"]F���
My����
�y"���+�Z�hEkO�0�@������y��J:�҉��l¿)n���e ��y �Ds��7�`-��X�y���0��B� �.F\z���4�yr�-&�);�oҍ]#j��T&F>�yR�M�I�5 f"�^�\y�W��y�c#:�ͪ*
����0퍼�y��Tk>d���8��1p�+�y���損��dت�5�Whԯ�y
� $]�b�ĨGMZ�S��q @|h�"O�@0�W�.�lD������E�"O�j�.�\V.�{Sψl�"O�a�w/�r+��ʁ���ͺ��"O�y��CF�TA#h��h�[Q"O@�k�A';�ݘ��ĥ?u4��B"O�84L�;uޜy��!U>U��"O��iCnVs����]ڼkR"O�M3�[��j�*7c_e�R�"Oqh��L42n  rO_�{s�;%�d)LO|]��ev���GܣuB��"O��!��ƳqQ4�9%!�7b����"O%���vA<Q��Ư9D��Qv�'x�x aIj���� 垶s뾔��-=D�������"����U�P�Ȁ-:<OB#<I��4~J�5ك��;�H����U�<1ІM2H�v�i�o>�I`$�\���0=y���Fe�H	�V�q����\[�<y���.��Yh��Eڞ=P��ן��� �\���DV�A�b��(_���ēdW��K�	��9����E��u�f��v"O"�U&W<[��y�Z�䉃A�'�Q��)GC5=���@�Մ[��ЂC�,D����?]8Q���"?"ܘ(��)D�Tj�&�"�=X���H��@�'D���Rƃ 2�	D�!M� 32	#D��Dbʃ �Sd#�L%CS` D��Ӂ��L�q1��*��q�=D�ؙ덙yy:�� _d��U��$v�ڽ���)�禍p���n�[�@�Z+HL��c2D���Cڰ�$̚�!\�t,�Ĳ���<i"�'����Գ]��F �1F�2����~���<-�T�X�e[�Lj����k�I6�2}B�i��&"!�q�'��%.�jR�XrL�	c4ؼ		�'��01��:0_h�i���Cs�X2�'���
�� ً���ʸ��	tx���'=��[������ʠD0�{��'?ps�öW����(sQ:㓆�ۮ4H��ܷ�����g��N�ȓ�^�2bS�O�P���&>nd�'��	M���);EV\���(�w�2�+�ER��$ �-�(�J0�AbHh����y����	:
�C�o�88*槐���'G�	E?��t'�
�T9�1/=9+ yZ5 U��'�2����]	�|�U@E�R�ʡ��O�b�$�Ov�X�=i��H�k�j���W���"�|�<�'��X���(S������(R��㟜�'�1O?�)�˦F�����Q)�@��t��`��G{Ҍ�(*�"1p�A C��Q��G�M�'6�OD�>��i�=QxI@ġț_�-��$�N��ow~�c�j�j�y���+�M��JJ��?��'���ŋ
7���xAE@ 
�hi:���s̓Tn�����aɣ|&�̨��P��䭸�"O�q��˛'(æ��u��#��!�WZ�y�X�T�S��O�����
��Դm��T��.y@-�ȓ}�@�bO�(:$�#fS�^��(ۧ���O>�{�<�S�̎=l0��#"�.��ȓ5��pSN�Y�0 �j~���ȓY�8(㗦M;�)���B�Eyr�|�wDU3Z�td`?RsD`�-�}�<�`���4�`��<5��|钪
=ў"~�	�Fy�����%���"�ȓM#xB�ɩ3��!fAR�;��1Gn���DB�	bf�CbE��Y���>o >B�)� �m����d��#��f��"O|�T���o��}���>R��4(�"O����ɡYSbax� R-9����"Ob�Ve���{')�6����"O�t�U!�5! ���TE�N����"O�HUoʓWԍ��䋸'�����'��ѠqL�H�� ����1��8��'�Za�4�=���Wi@90(	�'��!pt+�V}.qZ
��;o@{�<����(������[%]�����[�<��+O'{��Z�,ʈFW��zSgX�<�r*��F
��C�.$"�pщ�k�<aA
�&KM�4�jQJ&>E�A_L�<�b
޲k���Ff�t"� ����M�<q�ʗb�8�&O݁��EJ�yBXV��i�-�x�ҝpdl���yA?_�}�m�.v;�؀���/�yB%� !���� ��\�� cJ���y"�/Fk���w��N�(�7�E��yr�Z"x�A��Z6H,������y��$}�0"�͜�?��Ag�ú�y�N���9ja��,G�Vt'j�y��H/.v�B�N��6�P���Ə�yn�;ٖ<�jG1�ܭ���yBḥ9��C���QkN��Q�/�yR��1gxV��߲AB�[R�Ԁ�yҎ['
�T68@�zdX�#U6�yI~.�(h֎48+TqkU�yb.�y�|t	f�P�7�$Y3�o^��y,
�W��x�X*�ؽqş.�yK��2�6�&%��-� dP�y⊒n]���p��O���P+��O�I�I����uD$YV���"O �R+^������B��F��6"O6UkP�P�4�1��/H|3"O�=1qς�P����ݚu
"��"O�T�`��^Ad]X�'��P��0I�"OڽV2%��$�2X��x�"O�$鵄��`��dC��:�Z"O:�@�E[<Q�r8at�ȅBA�M�2"O��(!���� ��ֆW;���R"O�9UJK�Y�H���M]h��d"O&��3�</\d���m��wC��r�"O��g(&P9�3�O*u j=��"O��pd'���Pl�%p �љD"O4T�穙5I�pe�F%	�_���1�"OR0�S���3�b��g䇪,���["O�LQGQ�e�b�ڵa�9$�z8�E"O�I��b���W�Z75Ζ�"O�,�0/�JZ]����O����"O�e+@�ǜ8�&���ץh���#�"O�:ֆ�:�d�������xb"Od���B�.eN�T�ŘW���y�"Oz��gN�!�`ʐJɺ"�F �"O�!)�*�d�n90�J�3�b��D"Oꔩ�O9b'�퀴�Ppf�)c"O�H�i�B�^x��-�
gB
e#1"O��!d�g�%)lOF\"E�"Ob��T
hz�K�?X�Ju"O��5��x=(i�gX
��Urc"O\Y��C�
��v��IGP���"O2`�A?:.��e8Vly�"O`��!�Fۖg���B�"Oֱz��ڌH��9y����ll�I�7"O 	��e
�M�ȕ�DQ:h�3"O� �U��˛%�����·B��Ap"O�%�V�Ԣ	�-iUL�g*~��q"O�����O�%�''N��G"O���!W"z�t���$#��Y�0��(f�&D9��i��5���PBJC�Y�(�i�J{�!��S%5*�B�ݾ�$�76Az�"]a�I3Q>˓e�&���Ɖ�@D4̊��]�lJ�8�ȓb"��"#iN��/S�~�\ �J�1���	��4�O|� �S�I�H�j2��3)��i'�'�H-Y������>����`�h�zq۱N�W�~фȓT(Z��â��Q��>@4��<A�m�8L,�p��5� �a*�F�;�����ƓA&���ȓz��+�bݶ�J�@s놔u��'oP<1)��'�*8
��X�7#�^�xp�O &����2D�8�m�;6� �k�-�T���m3�r�C�^�B��|�N�*8��@���	z�2�� ��#�0=i�-��aDu(��?�ŕ�a��K?IZ�hx�.�]�<�@�Z����r �"H��l F�q�I��D@����A����D`%��x&M����VjP��*�v���-� 7�&�͓4
���,Ƽ]�L�P����q�7�g~b��* �)P/�� �p��yrn$�hY�S-0HD=2��\M��U"�jV�:�VIA��Tc���Yҋ
�"�x����<\hJ(=\O�1�r���J4���/*���b׆�n����v��S�.܃�'�<X0�
��G�T���L��p�u�}r`\�G��������>�Q>E�s��0V�|�#b�S-�%��3D���@��%�ixT�<�tPhbܞ��9mPE��S��y�M�HX��	d#��n���P��y�H	���H"B�^׺�-���'���GÅZѲ���	�&b�솸��A����:����$J�th̡�&��wt���������f�[c<9��"O��IjD�Y����&��P�Mhb剄'���aE*g�O+�쒡2#r�b@k�f��y��'sp��b�ОB�,@�db�J׾��47[��sH6�)�禡i��F9[�,p� �������y�\U�0!b��B�= ��W��y⬞�(��!P��J�P�RƜ�yRCV0����m�L[B�jₚ��y�*��is�п@��t�"�P��y2��3~�����1�Q����y2%�>B�H]��%=va2�N���y2/�6DdP��o�*��T�&l_�y"��� ���Z�"���&瘟�y���[3��,�� �J�6�y�E�=/��:T ��,u�t �"�y� �ͪ�&��Ze0��D�� �y������ð�_�SxpSs˟�y�
�>�Swg(Υ�"�N�y%ĩF�-A3����1��y�&@sD(�EL՞-(�3!"D��yB��7w���0q�I� qEk�Ŗ��y�͓�1���B ��[��*^��y��
�xj��A/��x��Qc��y�c�v>�Q�񂅉/��(�!��y��~�<xq����%fց�⸇,D�$�qn .�jẶ��r �h�B�-D�,x�G�gwD(�w�3�R�6�-D�h(  �^��)�G�f^r|��k+D�0��N����& N�p�q�d/D����d��~��J��AiR 	AD1D��P�@Q�Og�l���u, +!K/D��I1✼�Z6�2B8\��K*D��t(ŭ=� ��4o�%^
�TO(D��y�a���ш�'��m8��*D�� @*�G�]���@��<~�&,(�"O��p�-85��������5"O���3�E�~%,�iK���DTxB"O�QbO�ʈ�%J�M�܈�1"O��EN�x�΀a�C ��x�"O��"��G�b ��
��U"�"O0i`֥ �y�u������"O؄�mW"� )�*�=*\�@�Oڌ�m (��|Z�NO ��=�$�	><�	�
�'�^(�U��3^������y:�����d׍|�r��6l7�S'��=P�EI�_(���҉��D�(C�	-[-L��G��*?6DC-�*�<�jD\����hK�ҧH��A:Q&��P�0`� ��{:ҸӁ"O��� �w��A�j͖F$e u� }��U�)�(`� j"��$��X3���v��3y45�#F߽Na�+N�~8CP�U >����$��a�Ҝ�Ճ�0�P�?6`^*A}h�|�Cĺ��Af��tB����r�'"�ɸ�,1.̨'?m$�<q
��̔*��)@t�f	�W�B�O┝�J�"~nZ�(_�Xa�C�>S��T��n$������$K*DҧH�2\�#@s��\��aG���j�7O� WI�4-~��
/�p<�횝~!��Há��J%�T�t"���	�Z�@��5�ħ7"�0�!�
ier}�&�;�qK�DԽ5���to]�G�X�cQ�'��H�B�TP��u�X�f'������"�m{Ek�	�AA@��J�U�����]�'|���`��=Q<�dy�@��F2.�p�N�p��I@�44����2/2�rdZG�d`#�9;�� �BC��fC�%yt�>&��*Gz`&n�$i�0��'�a~"\(gK�D�=E���JT���GN�c<J%� K�"�\X5 �-�U`f�U �9*��I�e�Jdx���-i�e�1n�6|���i�Ԩ�tζ�� �>p�(�O��1㒃� i�ҝ��Ry�Dk"�$D���ǃ	�/g�E�G���'�a��	�H"�ѽ\L%(�΂s�z��gO�$R?��@��Q��X7k�
y��`ju�=\D58�,��y�kC��n]2獦H�:���T���>�3B�>3�8Lc-@�zcʵJB��JB��@�"�H����) ����ā�9b
	r̀6yeĩr"hQ���DP��Y!��\7�ɛb�S:��@�Rl$ړnZ��l֏h��p��Ƭ4ئ�Ov(��R��6��H�3h��/
�h#U���/�tI3�m:�E�"@�7Pv*"?QBl�!Q�Z�e�a׌�BCZ%Ų:���&\�A�M�)!=�%2�[a��@�1hN@��m�d��"��ؗ|��d��E
�e�8������q��� � �	�^�()aW�_�Ed�X�!�e����̓�q����jfɞ�X�6	�ឹIz�̻zZڍx0��s��0Ic�:O����I�5S��˔ �|VΑ�/�8[�����#��6���䘫�A�OC��rၸj#NAX`��;^�̡�DN�O�x{�b�Cќ�h���V�0����'2�D�vBDO��aq�����A"Cm`>Pc ��%Z<ْLӻ���2%� 4�Mr�e�)� ��q!Z/,W�DR�7���X����J���f^k���#�ﴁ�t�Q�]f�y�6M��7���H�{���uf_n���A�@��k1��e�q�l:�HLԩ�'.r�s�.�&93.���h��X�pH��W�d��D��9k��	�_㖥Cci��1*bk�%�
���* ���,Pp�'�6!��Ṡa0|O�}+���:��7,�ġ��j�T�b�s�Ƙa-(��U�δK�5��;�AW��hx�H�b��%@��t8��D=��eS@� �td&<��.?�I���ͻ�l�8}P9�f�����ݿ
�B�8p��24� �
8'R�,؆���DIP#�v��Sb��lY���ɓ=[8%�r"�[��ӗJ֛K-�(��e��+"�m?x�n����I?\,�b1?aC�E&y���1j��| X��WeX�� �V���x�'Ю6�����Դ2P�� d�W�%z7Tq ��¶�Kv~��M()�N(u�o0�կi�!s�o�PF
y��`�a�%�O�"����Vܹv�ͧv��=�d�C���tb���R(ji���$ O��Ʉ.z�'�\�* ���{���5HA���%�
ÓN����ΓuͮP#A��L��k�$4���D(æ41Z��M�5��AJ��$�ш]7pL@��Ҫ�K���O�����ա�~�m#��i3��|�'?h8����hM�y��E�z��M������i��uѲ
���e�'?\\�4��T�ɧH�4�g�_�lD���)�D"O�n�E��E{�C�a���Hc�|���`��ń�Iia�|��� S�TD��ќA0C�ɂK��@�AhI$"�8�g�b,�C�ɞp��|��G�>L����c�
PT�C䉸!�. �Ë7h��X���$LC�)� ��j��T��p�7�NK��"O��B���e���2�T� H�퉲"OB�%O��|8�pb�'�2�if"O��� ���%�&�ٔ8zi�"O���QO���z��ٷz<��P"O�sbc7�m���^66(�"OF�C�JI�v�z��D:�AA�"O�۲�޵<B�ȉU�@�T%z��"O>-�R���+k�}�QI w4����"On1����N�:IZw�*�( Y�"O��	vl�ڭШ�{�@�)&"O��E�I'M�N��K��E�"O�q�Gb?�N��2g ���"O��Nк!J��K .ׯQnl*�"O�2D�K�4�"h����#LV��J�"O�ȅAJ?3��I󎐖{�v"O�Pc�)6�b���.,y[�"O�)qt��$g��� _��L��"O�D����e8��=�jY1�"O:a;W�к}p�ԭ
M�m��"O���q)K�6���ND<<��6"O���䜵)4�aH�픎Z�j�ȅ"O��I����iq���G�|�8 "Bi�<�& Ȅv��pr2�֓3�1�Ǉ�e�<�#A�<��9��g��vT05��h�<���9|H��+��)EҨY� m�<6��+)+	��L�.ah�Bh�!�$X�F�R�0�Wl�>,z�K/fz!�B�+^UX7�҅
ee�f�m!�D��',�qN��T Zw��JL!��y 5B��7S�Ȅ�pi)3!�dX�f���q!ݕ]����v���U)!�$]{�H� �QS�p��gNv�!�$�`%�В!�Z���/�!�$ȳD��r�٬M�h�]= �!���$ԈT*f�Ǒ& RM���Ȯ0�!���|�vmC$@A�B�ߗx8!��^��iv
��E��`:%� ++!��7-�p3FC�� �jE���n�!�D	2u]�Bi��>�Ӈ�E�&�!�	�L��hIp�Bq���'Ҵ}!�A�c��\K��/�R�h�
{h!��Îp�N�aΏ�$�F�ȳ��/S6!��J*�����֖ �ȭ��T2!�D
�9��
�Qf��қO�!�d.(N���H-\F��hӦ�W�!��	6q�Q��P�HT!���!�dW;O�]� M�#4�Y�`ƃ-0!��w���m2a�p��1��<!�1R����++|�����X�=�!��^�e�!���<Ze���%�� MQ!�F5'�UAG$P���cB��4!��K0Gj��.t\�ܨ�PT>!�d �AB
'W���1���-*5!�(z��R��նhx�I���ݦ>-!��^�� I��˦Vd�Q.��h9!�$�)J��cv�D�E��Ej&-
=/L!��ӗD���S��,~��EQ��[�k/!�Ā-!���b�&̎&(P�G��Nq!��-M�8����9N d�a���L!�E;�9S������ZA�2S!�ŐQ�D%��@�_�k6͇�t�<�b��8q� �Bȯ�z݇�p&�T�7C&�4q�5�,`w�,��S�? H��֨��ٲ�ΘI���JV"O�5)��Z)Qv�)6͗2��U�'"O��٢�ˁb]ĕ�q� �T�29�W"O~c��N�X�	S�_�_��81�"Op%Bf	�<��P�G��:�����"O�E)�c�N�N-�t��%%�{�"O��
l�e2��QR�� Ԅ$IT"Ol#�� *�m�a�Z����V �2����N/h���aZ23��IP���4�!�DڪGmd�*⊑�Q�
��"�[TA��R��h�	UEQ>�9�~y9�ϒ�-�L�m/A�YL���t&�@ۀ�BP:� qV�Bpz*�HG�5�&l(�#,�O�4Y�Jǉk����:u_`����'JlJbH�+�tu��Ug���T�>N��j�T}�ȓ&�mz#�W$s���`3h�e����<qc���c���P�+1�'i��铖gI�mgY�cie�Z��ȓW���p �!�����o�Y���5�؎���'������ש�t�H���\�*�*�:��+D��2w	�8\~d�`�昋D1H����ǯq�t��%��o�|���4&��t����B�|��ߡ�0=飅�#R�Z��үЬ�?`G�.>��@e� N2�AVDn�<��N�k_�x���W�L����r̓V�B��FQ0�N ���ӋH�
�#�K�5�&��CЫF�jC�ɠ�Q���`&4`�l�F`%��a�����d�I?�� n�����y��aA�@}<`���%�31!����Z|E�N�e1���A��N6SLZH�a�Z�p=iH��T�{V&0��T_n����U"IB(8%�7K!db�jգ�Z�&��Ń��BI"O�����[4M��`����Ȥy�u�D�2h[`��f�Z�lԢ|Z�ė#�v���[ @�20*�<�QB�
�P�xt�W́�Ae� zI���
D|ӧ���xRx��3I�����Hנ0�!���J0I�M"v�J]��葔a����x�2�hԴ�p=yA�'L0L��ai���q5-�d�L���M*j�(����S://���Ө�h%�qcv�$*�DC䉉$� �����~�v�`6eE6=,Z�<��"�&�����E	#�b1��X?!�T��So8'6!��ۃJ<�6��xn(�gnB7	 �c��f�b�=E��4/kNPK0;���д&��SOvm�ȓc��,yv']�ϖi9Q �+U�2y��nھ��"�E�d9����6��ȓC�l�q��ߴ
��FD�,/�b��Jf�lYuʓ;<	
]"�"X�k%VD��M�ȼ���m��E�cg�G
�d�ȓӠd9��R�5��t����=:6t��E�3�ڂL�>�z獒�	~$5���:�f��X��$r���vf�Ň�YU���H� 4���2X*����	�֙ ��z�)p��s>�ȓt^�	s��97��H!�������`�P��(ňi.�9q �*CaLɆ�aМ]I���Z�X��A�ߧ��ȓi�N��e术u���[H�#*����ȓi7�#%L?I1�QKP��~ ��ȓED�8�WE%U���vkO�|~��ȓ\��p����c�
-�b�X,���ȓ5�� #�z��	Ё� k����L}����%��]ʀaLG��)�ȓT^"�J�����D B'3� �ȓF�L���(
u\�Q"��>A(��N�Hy`��X+p@I0�;d��hB�(���O���h��1QdɄȓ,�uH���d#��b�0���ȓo���� *!��7�Pj�N���S�? ��ڦa�g,� !�����"Ot�B,VQmb��"�(p����r"O�m����S
EA�ᅕHL�Iq�"O�m�eBę��J�0���S"O�i���$=�b�!I%v����"O�@�E�JюD�`#�$)4  �"O�0���ھ2�T�bբ�tP�"O�x�%�E4�؉b!�P�{�0��E"O|���D�w��Q��JU)/׮Փ�"OZ p�V�J�\!ɕ�90���ke"OԩՃUd��9�m�U��@ B"O4���LI�b5�'�'U�cO6���,�%"m���JUk(�'�O��P*
�'���
���P�U�>?�������C�(Ux8c7�S,YN�"����d�2����CyRC�ɘq�&di�j]3@��ɴF�7���U�R���'7p�ҧH�J���i/.P8%��?}&�#Q"O�5�qC� }PHԂ���=b� �bE<}"i�$�D�E*���_)Wٌ��Bh Y����䁨��?�"#�+Q�t����,:����<L�e(d�֘LyT���RyI��(FЈ5��ˤ�ˣ(����c�OF�u�R0�!��$
]r%��:�ǒbp��`�'Z%�y�Ύ�Y�Tb�)M"M:` ��k ��$P�Mc
Y���I��)�'}{��A3-΁j���@�ŏZ*��o�vp
gn_R!���!���N��b �H��1I|�>YF� Gk�2W�K>%y�䒐�G؟���L�B&tYÄ�?#����8"�$IY���4M��� Ղ<:�I�&PhJ�"���O
\+�HX%�b>���Q]GX�bU�4gJ��gC D��r�5pMBg,��s���"�+?����4�P�"|"��F�*�dj�&�"����SE�<y�L��N�)Wg���x�9�B_?��@ι;1>ո�O9��Ar�OHI9b/�5z�MPDB�;�F��
�'�L� FF?%�dpd &�F�`2k��Rd`�S"�J�E��p��T����I�s� �õ��
�,!p0fX"��D؁,'�P2�����BT��2-�CV�wn<���l(J��`3�Ol�
�`ѐ|����SmԯM��t�I9���$��p��|[U+�(�.�ϧ.o��a ��Lz�A�Ȟ'pǼ=�ȓN_01H��8!�x����A�Wm��E�F�<�s��F���+�ѳKX:9D��;5��5hSlW�$����&��Y*͆�5��!�)�Z��L�A�+3��n�ꄉD,YY>�@rkF�S!M�L"<�"�>o^N}QFX�s��ide�C��@Za��EQ"	��b�E�2(�5f�%]C�����.�BT�¡Zo.l�E�	x?�5H�C#>i�b�2DI<l��,��6ЕiТS��3	V43r�Ħ`��X��ؤdS��{S`E0��TIV�����B^�P��i�S̈́��`%�*�		/�}Bi��t	R}���� W�F�KB�ի�8!)W�T�~8�HՎT9'rR�� �tVu��{��cb�ի�y�K.w6� r0��(vNn���L��yR$уAK*9S��îh~��s�Q:A) �R1R�.К���,zȉ$b��I�emu$(
'�w���`�.��AT8�2��V�s,�@�'�b�j�!搸0VN?z$4���ɪM��D���J�i��	�_LTe��ʽR�d�g��#=A� 8K���P`�/F: 	X��t� ont�&j@s��	K!A�\�p�iF�j��Q��<�*5r�l�:��݃7q<�*�W��!b�'��e �J�
�|๵�q��y%�܇�J���.��](�#g��W��q1���1Og&M�va���e��o6v��&NO>�y�C�B�n���Ud�&�s֮�3? 7MҭZ\�2bL�D�I-]H�J�W�v���6��HIU�%h<�ӡ�Էy�p�bd�'��i���ѽ6W�M/�ݱ��K2M'�غ��S��ħOJP����,����	49#=A�L+��i�ʞ�|��pP��t�<H!'�T�x�ϓi0�Y�fȟ�b�`���ۧ��J���ɇ��������m0��/�>p��AD�>���O�e�e���~�����W�|�'#��H�ԭa���Q�,u���P�b0zqBэ>o�؇��iD��'�j�Q�f�?%�ɧH�4��E�@���;goU&)(it"O ��`�GrX��./VPU�|�n�-RT��)� �1��hW�f{��2ҭ�z�8��"OF��� �ɸ�A+B�w���{"O� �����5�T"G�ص�Bq��"O�0�ǡ�3�Lh�o� "����"O*H�O,a�!�]N�\	�"O�[���괥I�l$*�$j�"O��[��άf��(�DMʈlV�c"O4 ��B6s���0�リ|D�ҕ"Ol�J�f�?/6�0[��^��d�e"O�Q+s��-u��[Pʹ\�A
6"O�(RBKiv��kƆ��F��B"O8�kW�X,�f<2�%�&���8!"O���ύ�X:r([C�]�D��@�"O%�VBI���yp�'��g�Nu�r"OKWe-"XH�� }��������yR�ʡR3�@2�@
%l\tX���ۺ�y򈒞y�J���/�+[�"T`��U�y��CD�L(�@��V3ػDBѢ�yR�*MD�Y�/W���a��AY��y2��5"A�0�%
%�P,̰�y���}�B��������@��d�&�y2��	xd�����>�D�cC-;�yR�~�2�*e I��%�� �E��,��a���ZMhQ҅����a��4D���dC�����]VH��wo"a�Q�]2X���N�Q���ȓsh�q���ն�v�u	�V����&AL<`a�j����ڜ{+
M���0\{��͡�b���`��z~긇�HҬ��ڹG*���tg�9Yo�E��t4B�A݉*(P�')0A!n���QH�cƂ�/gRlX��)`ଇȓI���2K�
b~�c��X+`�Y��QJ ��Zm���$
�����ȓV��!ӡ`Ͱ"^�U+&*ޝGv1�ȓ,nM��IU�N�q	�#e�Q���j�E#L�D����A�V��}��+�����I;@@Vq2��)o@�ȓ9����F,� %>u���R�md�͓m�0* ��]�4��֡�>���G}�mT�vs���eHA��)�5nUf�<a�זW�<9qm�	C�)���^�<�1,)�b��a`Q)�̅��L�V�<Ig��/(-~(#)�"`��̊��V�<��HEh���AH�
�&�:Sf�O�<���P�?��32G] BFf��R��`�<q">AX��í��h���"k�^�<)��X���3����.�	��P�<ac��W��q:p+��	��
c�<� ��Q^P��v��z%����`�<Q�튧q�<D`�O�>ey����B�<)�ǉ/?�H	Zg�(�x��Pw�<�eeF�qt�h�W�{��U�"!J�<�p�Օ`e��d�O 8�\�y�WG�<1�P�tP<�A�'�t����o�~�����OF��!aL"]��.4��G�6Ӊ'I
���{�S�'\jU8C�N 2@Q#fN�Vcx��'w ��Zq�S�O����5iΗ
hpS�L�,Qd��:ݴ?�$��B!-�)�f�ƅ/��Zcl'WA��a֠��'ra��C9'�q,ˇR�������0�O(�2�	,�3}",��n�t9�0�!����dݨ��'ў��ԩ���ЧQ^���zt8\ "OD�Q'B9�,IU���g��q"Ot��5�[;3�r)	�']���9F"OL�)�f^a	(yZ��İ
r��"�"O� ���COA%9��+�CQ�]�8�F"O�����A<UP��[3: ��`T"O~�r"��Fn&ecF���sP"O�=(S�p��!��Q���Q"O�����)�`�F�80����"O�I�!�2���u��4= @,�6"O�軰-$m&��b0�$Y�"O�H R�Z�66\9�!xF� "OtPR�Ҕ	��,�R6�4l�""ON�����:q���ƽo�0Ef"O��j�!-��lk&��QLH�SW"O\�%��z�.�xG�� 1"���b"O���� ;b��h@D͏C�����"O�M�肓
vd�"�	/⪠��"O����G�v�x����I�a�<iPR"OdI 0�M�vg~��h��n�B|y�"O�<I�n�'8�n�1F�<���
"O�s��Q^ c��6,���"O��h��ܣ[�&�C�X�[�"8��"O|�[��{܄�xs�\*xs�\��"O=��䐆1�@�ڐ�L�wNl�1"O���8c���U� ?�bI`�"O��W왴c�$��o�Y�\���"O~����G���e�߉+P`��"O ��B 8VǰQ��;@����*Ob���̄�'G����Gg�DR�'�
��d#��$g�9q��ΦZ�̨�'[4s��·(�p@ӓ#�'P����'!nx��d�#l����йD���b
�'�
l��?0;�u�S��@}�L�	�'���ф}6��򅑖3z*�R
�'1([� ۦ4
Hk��>8����'�*�f�� 1>��b��.l`<��'s��F�F�Q����"6,��q�'5��yd�ݧ*l�����<'����'f:�zC��I�)��e	l�Q�'Ϥ�p���8+]l��7���ayju��'%�=��僡[� �B���V� a�'tF`;���S�P!
e_�{i��[�'>���3k��@y�*�'\7K״Hz�'���@�Ļ'��q!��5=�����'d��A T54\H���W:H)�TC�'����41���
=7����'q8���) ��:�� *jL:�'C��A��S�	��߯x,L��ʓh�>l:`���i
����Q�^� �ȓ/�"�j2�F+���j��F70����q-�)ZS��30��&B�S
l�ȓ.�"��� ��,I�8�d�ȓ)��CB�.a,z�NF"�$)���(y��횜�j�6�R"+5���%� � �ϥRw���IQ�K��D�ȓ^b�������*,��&�g���ȓx,�	JC��8�X�Xu)ߵZ�D��#��E��\�w��|���4!�-�ȓ,i�M"p�
1?
e�f�$��ȓ%"
4�1&0Fy �bwcKO�6��ȓ*�<��lU�c���z�I�JޞQ�ȓ\�4�VMH���j5�I�l%��k̐�S&��#'�)�ÂZ�WK�0��'�|`weۀ?W�ݰ����x��y�ȓ���*�kL,O	�M�d�޴u����xg찲�
��;Դa�S���N:�\��X�&ܱs#]���i�h��i_Hx��S�? x���
�������28�t �a"ONAᲮ�xG��Ya�Pbo����"O4�� -o�<%����kh��a"O�U�&C��*yQd�DYj��p"O$U)�� {EDM�@d�HJ~�a�"O�Ȥ�\�(8}8���Xl!��"O��!3�2��ޏQ��-��"O��2��[��@(�Ø�d("l""ORhE�D�Z4�Ĝ�CX݈B"O~$����+P}��D�B��Y�"Oh��� !7\I�����^��<a�"O�,��D
b�<�Q�ʐzur,ҧ"Oxc�7+���1J� Fkݑ�"O�!��4(a � p�g�z!��"O�qkPUQXdx;h@�Z�X��`"O8����ǫl��5ْ�+(��9�"O�8SĞ}0B�j��F�G6�ɨ�"ON\��J5 �d�)̋��DaK�"OZ�qǗ��v���[�=����"O�%p�D�0���@�
�ѩR"O�(d��P�)���Y�[��8�"O(�:�5x��\��Ѣ"O�,�F��CT�R*��@�����"O���p[�j���c�{a��b�"O:�;�	U
7,9�5	��e�"O�T3�C[c�E����"OUK"Y�F�%Bq5j�Ԑk�"O8<�Eb1��<��V���%"O�T��h %>�$Xcn8�Fj$"OhY���ü��}��� �$ C"Oα��"v_䡀s��?
�0T�u"O&�#�̦I�j�br*M�9��jP"O�Q�r��1:=��ʃ�-��*On}zbL],����Y�wsf
�'H��hE<C �(��ςg^L)P�'��M��0S�h�!�d����yRK՝)9@Y����"��e@��'�ybe�(woB����!.(� 5��:�y�	�j���Ƞf�=+�8m�U��:�yR*�0���%C?v}`<�Um'�y��@�u�����U�{�x�i��W�y�A[8��� 6"ӛl��s�Z.�yb�D k͠�����l��kW����y�ZA"֤"2ba@Ԝ���ɲ�y���ro�q���\�`��|	�&ן�y"CZ\,1��M�Q�p��2a\+�y�a,7�����7I���ɞ��y�ѬU<��8�o�0d��-;W�@&�y��|�V�C��X:O{&MJviW��y� A�T�]�N���`��R�y2�U[��cE�Q�G���Ced�/�y����?�^9��"�>yn�Xe�N��yb�� <��|�v�A%�ĳ���y�G�1�l| /*>�lZ�`�#�y���SZ�Xs�
;^ID����E��yCܟ>���A��Yq��'��y�*��[t���c�,<� Q �k��y���yF��KqeٜK=����U��y��Ąq��)��^�7P������y�AS:pj��g�'B+0AP��0�yR�Q�68��4C4@5А��T��yB/ܖnB24��EV�4pR�����y2�0Vl�h�(~�`Y�"���y¯�e6Ԁ#$�w;�(K����y
� ���+�@�8�bC._�_@����"O&�P� M�y$�����˦v!��"OX\���O!�5�_	��a��H�<�0�/��C�!H���a�ZH�<���<x
 �M�r�-�FC�]�<I��p�d��m�5D��үM]�<i��,�0Ԉ��J�
���AMV�<х!��3�(�go	F�i"e��T�<�Ѓ޳&x���FE�w��{���U�<A#!͌jM$��bV6)�Ψ�#��T�<T� �tҞ�����.��R��g�<i�S4c�mZ��ƕ'otzS�[d�<)�AޑR��C� j�n�	"��K�<��ɝ!h`�`�n�4=�`�)�H�<ɀ,��?_n`�T�������F�<���:�p���>4nի�"�X�<���X<#b.y�V�\�{��O�<y𦆫q�N�4�@]A\�#q/_J�<rJ��쌻rF��!�z4[��Q�<�T�ڹcE��Z��
$�] 5�@F�<�'��0���`�䔪sO����(z�<��Җ]�ii�KC��6�v�<�g����؝�f�#��r��|�<I@�H6"��qe�589.h�3�Rx�<	u+�xI�"R�4bx��u�<ф�� 4�]:G���]�:�TBt�<��FB�%Щ��(Ǆ/�VyH��s�<y��Z]�4���Y�v+���n�<a �Y�0{d0h�/�|�P��@�@�<�&�U^�PQ-�fdj�Gz�<�'��a��=X+��q��@Z���w�<�Cp�@ՠ'�T�g xQ�L�X�<����P�`2#BЇd=.��Q�P_�<A)_;5Jzq�$e�(M�ޕ;�.�]�<a��	��4�)c��^p�a�gOn�<y�$\�}8����ֽ1.���Ki�<��K�;ƔMP��@7_&Zd���`�<`d8�0}#�fC9���pA\r�<�q�Z#-�:�2�n^>~�p��k�<A�bJ�
�S�66V���Lf�<�e��l�O�p>����w�<	WW��`�qk�,F��˛r�<�2����qI�c>~Q�H�b �j�<��+˂_h.���FF�X4buCPɟk�<q�hC�f��yH���o���#eWC�<V(ЙX�,���J}������C�<���ʳ'��+����L�.&�!�H&p�RE"��A.w�*�ku��>�!�$��)�P88��σ�|��B�J�PU!��	�����
 ��hB��;!��kSxH��f��K�@Ւ�i�<\4!�$V��}�ƀ�P�H�XEhO�x
!��JDƄ��B�yO��#�� !��>�dp��8%B�\�ʽKO!��(�f��vnE_,��j"J��!��Q=q �����Z��I� J��+5!򤎓_�0����CsAĔ�&J�X,!��տ9ﲥ5 N@�����1O!��m
�E�G�ɵ	3�<iDҏ�!�=u(]���F9�Hւ�=�!� �C�"A����™M%U�!��O�s�N�Z�eR5���� �?.!�dɭ<K`M�đU�8p$�0h!���A��pH�H�>�1� �/�!�� M�e�MF.�i���37�-��"O�mҠIƣ.X5sA)��  ��"O�5���+vl�3ƘD>n���"OD��V�H���m9D8��"O&���   ��   �  l  �  ;  �*  �6  B  sM  �X  �d  �o  y{  ~�  ��  h�  G�  ��  ۭ  ;�  �  ��  	�  ��  *�  ��  ��  R�  ��  =�  ��  �   � � � T! �* �2 9 �A �H �O 8V z\ �`  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" OTp�t%D��1k⭋�L���ctFR�<����� cE�+���+��N�<��+�7ƨS�g�s1V�85LL�<��C؇N�=Y���n R��@�<��(K> �H���"?�B����A�<Q�+٩$�2�*�%{F���**D�� P	"��)Ku�Z�5�&���+D�H��*�5s���i5.��en���(D����gR9&��J��F%�@ᆌ#D���3,�&���bf��*1b1駌.D��#�aիd�Y�(eot�zѧ>D��y��@~pH$�@���	3d2D��%%ǐGi*E�$�Vd4�;0�#�IB�����MN2D���8�HPd�<�;��"�d��M�0��l��,� GD���R���ƓiV�e�@N�(Z�b5�k�7i8)��	7r��#<�G�ω(�����<D���o�<���~�(\��`�4��y��Hj��x���ODZ�a�T9mVd��#�	c���'����$�O1ք{S+��(g恈�'�<��$m֟,z������8�[�'p*��)�E��lIb�I^0 �
�'[����ʊ#t��{�$] I&a
�'UDKfK�|���NP�FV>��	�'T%���ߔ*QD!��h>�A��'������6��^.�4�'��=��ZX�>U�`�lJ� �1�I�"|�']F�����?q�� B���8\�C�'��P�	�u��i+ M���� �'Z����ȑi��	�w-J�
��8�Y���|Re��y
�iB�L ~�B�[ `��yB�I�m��#�F���T���͸'������|� xQG�>g$eB�+�y�,g�$��U2`B&�A�%R��y���(#c���-F�,Hm�Tĝ�0?)O�Mi��O��xA3g.@!��3�"O� 
��u�^ڨ)�Č�"G:�4�q��`�O�m�%�9����Ù�J�m��'�*��/X�90��I��FmH)��'�4�Zr������l2l%zx��'�xa	�j�_��
_��x��'��1��ۃ�j��� ^#�"���'q�Z��E:GF�r"�89 ��'�D� �Ԏ"���+�V=gXt,q�'�6�b��U�^qQ
LL}
 Z�'�lA�p�F�1{��H@Q�I�b5 �'�&�ʁ��M�܃�b@�I����'�*�ʷ��#F"|Dە��-B
���'���1�ϖ�iʢ��_�<�P��'ń����S�]�c%��'
�� �'��q7�yc�4c�cʧThts�"O����E���9{FBc�89�"O�@B���H|b�g@.G!TȠe"Oɲ᧍�J�����֩o���c"O��,�3:|��/�5 ����Q"O(��tDޖ[W�Q��n�4���"O��!
^2C�E�M��t-��"O����Z�D�bI��VJ��5�"O@!�a�3�h��C�5����D"O�U�#	 E`^h���ߪVԞTS"OJ!�&�|���S5큦o�@��f"O�%[��B-!e�d��kϫ{�R���"O�t&	ҧX���h�*�=w�"O����\�-��!U/�E���""O.�ҵ�'%�)�N�C��Q��"OXy�7HJNXK�`Y,RiN-@�"O���$F E��9�9c���"O~����/e���"��6Z�'"Ox��� �}����<����"O�(#���?�2����9w1bR!"O��pE��I\5 �K<`���'"O�("ע�1O�H� U�f����"O~��7�.5Z\��B2h��I`"O����Ꜹ)���/аB�nYs�"O�@농�ROȐ��A�|:X��"O a��E,��4�w̙3����"On�
sAM.f�b �
�,�&"Oi`�G(Zp�suCؙzxě�"O��
&a���l 	�Ns j�"O��׃�ZLf��2*V-X���h�"Oz����1��$"p�Q5lL5�"O�����Y����d�!q�¨��"O��;3�@=o�d�-Q99�4���"O�x���3zZ�8�+ ��̛�"O@�� ���>����ɖ���"OP|�%[�B|����N.Dg�-�#"O�X�b��;���,؃wa��s "Oz�Uĕpp	����
SR4!�"O���$�ΕK�n�X���vE��H"O�@
҃��B ���-x,�]!"O���]!;Dl�
1��>r��D"O
#�¤4�H�@=8���`"O x��O�{6l8�/#�h��"O2X�eNi��`n�	jԽ!2"O�P	�I�/�1.���(��"O*�ʒ���Ƭ��B����P"O��a� @H d#��qf\s�"O�A"�@�<�,0���W��`"O�Q��`Q�8�4�`��F�wv�H�"Oz��1�M�r���L�7Zi��"O� �z��ž=-t��K�OK�5��"O��b2�Lr�aP-1���"OF�c�΂�c��pE��Ea�"�"O
(��;T `����Ϊ�~��"O$�gN�����b-�>.{�����'���'���'n��'��'2�'��9�Q�wH���O6�q��'*��'���'y��'��'B�'$��I�`���Q
E!��$�'q"�'�B�'uB�'�2�'+b�'��pT"L<�����L�XoDU�P�'���'!��'B�'*b�'e��'�Z�{q�Z�]6����瞧:z!�5�'8��'���'d��'@��'��'6�!zӉ�/�  'I+t�	r��'���'k�'Y��'�b�'�B�'Z�lS��������j�� ��'n"�'@��'	��'��'�2�'��q��$զ,Q �'�}
6��'VB�'���'F2�'���'p��'Hh��EM�-YJ���}B%#�'c2�'�b�'T�'n��'1��'f�X�u Ņy�  �'H��.s�L�f�'���'|"�'�2�'S�'���'���A��27��0�y&�iS�'���'x2�'���'"R�',��'�\p���W��c��+׊���'���'A"�'�2�'���'���'��+��Z7s�J�&��;����'���'��'ir�'IriӴ���O�X�4�<
|��f�%��。.��ʓ�?�,O1��	�M�����+p2m(/Ǡ��!��/{�8�'�b7M;�i>�	ޟ�c"��N<(�c�P@�a��e����i�q�i�����*��p�O�v�1��XZ�ԕ���޺�h��y��'��Ir�O��X�j��&$�bD��w>����Jhӆ�c���0��&�M�;4v���n_��(ؘ1I
,&a��A���?q�'��)�?W�NqmZ�<�w�F�<`Hu$���bk�<��'&N�DI�hO���O��
�	�(���R�Fh���u3O˓��W���ғǘ'����gê_��Pd�U23�X$����OI}��'�27ON�5=	F*��S_�A�0N�Q͘a�'�r�
�&��5;��t�J��0;��'J�t��7�X���a	�O���T�(�'��9O�q��`A9>M�A"��4,0�7O��mڝ!hJ� �V�4�:X�.ʤ��L��⑅!�򽘷6O"���O4�DҚW6M2?��O,��IU;u�j�j��S�'�ĭ�.`A�PYO>/O�)�O����O����O�u���N�~A"W	Zd��	��¾<�d�i X�2�'�b�'���y�
[a��x�Gߘ>|�Db�#X�������k�d'�b>��m�+A��ث�Iǅ'�lct��r�r���t��O7F��x��.Wﺣp�xRG�<�P@�	 ك��	�L�P�q�A�?��?���?�'����)�� ğ�h��)T�h6e�R��x��b�$ݴ��'�P�0���Gw�X�o�0!; �PB�V�TE`�#�ǉ���%H���Ϧ-�w��8�5�^�fC| P�������*�ީAv��.�^4��� &����ڟ��I����	͟d��@��W6������Nv.\�� F)	�6��#K�\��#�' �kӞ���'�С[wϙ�v��'b��Re�$R���i@@D�b���i�L�i���O�l��M#�'U�Yy�4�y�*I� f�P�J��^Ģt�Tls6����x!`�.J��/x˓�?����?���u0zh���t�ȥ
e�I�aU2���?!.On�l��0e6��'�Q>�0��1i�B��f�S�EQh �dco��	��䦙9�����|z�'^{ڼ��b������
=#^���Ǜ"
А,c~b)o�MY��'��'��7�L@b.�Pch�x� �,B�'���'����S�`Yܴ�B�)�Tnu��ƌ�"� ��3L�0�?A��3a���DZ}�+xӖ��%*�i� IɸH:0)�l�����I R�	oZQ~�⒐��u�b�	.+dɐ�X,�pHh&� ����<���?���?���?�(�b��U.N^�`3�A��b��ަ@�ޟ,�	؟�$?)�I��Mϻv|b�hɖ!�DY"B�]������?iI>�|z����M˚'
Z,3���(d��E�Q��{��|ʘ'�(�C���@���|�\���ԟ4��K�?�88��,��;7�y�$�۟��	۟�	Xy��lӸB���O����O��+� �+	l�Q���z�(��>�I,�����9۴�?�-Ov�X��AA���3�ڝ������@;BY��9��*擲C_���;+�� v�V�	2���Z���n1�A�'2��'���'I��i�uK�O�H��Ԛ1�p���J0Dǆl����O�lVC^��'m��|"��y)`�Ȁ�o^�I, ��$!3woҥlӮ�o��M���4�M��'y�b��I�$s_c:���ba���e�@��
qp�d[��oy�ab�\��|���?a���?��f9@UU([�~x�1A�j�`@,O0o!JlX�L����m�D�'�2�P�g΢��2��9]�1��^�(���4�M렸iX�O���<���Jʶ�"�D\Zï��mr�ؓ�a�@�'��X#�M"��JQy�Mn�������:?CH�aw��%#|�0��8Oj��'��.�>r�Ņ@r��'9���0G<��'u��5jT� �AŇ{�J�3k}�董*)�����	�X�ߴ"t��)}�x�3���0B�^ip���!�� A���^z6mr�l��
 xX��7 OȲ����Zw�� `M9T(ƫ)<��
E���X|D|ɑ(�O`��O����O����Ol�'i���ͧ+&��i������P��Y,vTu���T��?i�� ț��T?�F�)}[PlJ>�U�F3l�8�JN03.�P�%�"Z�2�>�y�i��6���Y�G�w�|�	�Ъv��fK`���U�8�d��N��th��'�\1�'j:7�<�'�?����?ِ�8f7vs��^'y{���$�?����¦[@+���P����0�O�,��B�$�8D�q`�Ci 0��O�T�'B�ib���'%��H%�����ؙC ��x«ɔ��@Y
���|z@�O�H�K>i�ߜ1�R"�9hF�肀)K�?1���?���?�|j.O�]nڮEB��c��:e��a9q��yԍ������I<�Mk�B�>��i1�=��ЋmȞ�A����y�bXSM{ӈn�:��]oc~�Фm֜���u�)͊Jf��JA�� ��h"��҂5��D�<a���?����?����?i,�`qe�;�`rBJ�	��<�w��Ǧ���F�ן��ڟ$?��0�M�;�ҽ�� �_@XZ/46&D#��i|6mWP�)擌:h1m��<��
/�tM[��QW���B��<ђ����a�
O��?(O*������˟�QiuS�H0mЖ1����%�'bU�P�"�V��?q��?�O+��_'oZ��d�Oh�Ć�0���%�2��*�2s���Qy"���61rt�'�7-�����?��ɲ(�j�Y�-��V9r��+.i&�'�r h�9G\��|r��OҰQ��|��'�;'ߴ�3䀚�5�Vy��?����?���h���D�7l��k�'I�&�L��%�/}-<�d즥K��џ��ɍ�M��w,�<�Ӌ��H"E��`�-��H��'��6m��5شx%>Mp�4��$��cZ`����Mu�Z�o��{L�u��Kp�%@*�D�<ͧ�?Y��?���?YQ�t��p0��B���"����'��7-� 4]���O���0���O"�h%�)�t��un�Aᚦ�FJ}��'#�|����Ō!�h� F0��+7�%$��z�����$�cH��3�iƒO��A,@� �8�Rm��j���Q��?y��?9��|�/O�im�'2�����1��zVB_��$�'h�%�Z���M��"�>I���?y�m�Z�j��T
H�����jZq�2��t��M��O�-�ժZ;�(����!�i�GB���z�{�n�����O��$�O��d�Ot��;�S�b(�t)5Ep$
�;����~�F���ן��I��M�焙�|��d�&�|� X�%\t�0���6�� ��-s�O�hl� �M�'8��X0�4���A� K
�뒃F�0� ���iw앲�S��?��-3�d�<�'�?Y��?I��R5;�b$Zf��^��j��_�?Y����dۦQ�C�Zҟ\�I쟼�Ou
���%��*y|��F��P��5��O���'�7����a�O<�O�A9�Lל4����
L�A� x�3���t2c����4�P�B��jT�O�!v��R�X����5�h����O����OZ���O1�b�a�v�C�R�f�@����"� ���2c�T#��' q��⟔�O�$��5]P4��CU��Z#�b�@�R���O�E{MaӤ�̈́�����\�O(=�s�Y6%�z��ȟA>T@	�'�����	��H�I��(��H��-R!ϼ�܁B�:Ő����7��LB����O���:���O��lz���'eVCr<H�ea�.q��)yw����`Ӭ�O1�V$�UHlӰ�	8�&�2���26A�P�ǡnt�I/�� �'�x&�����4�'����&]�\r�Ʉɀ�N��r�'^�'G[��yݴ$k``*���?��4
�����53�lȘ��)V��Ma���>���?�K>����9(�q����3��2u�Ui~r	�ڀP���J)�O͂D��+m�rD�>N����6]x��֫�cm��'���'�2�џ��W��PMp���(�<[�d)�ǀ��<:�4J�����?y@�i��O�n� q��ba��&r�P	��� ;��S�Q��43U�&Cڍq�f����ҋ�~�d/�F��Qq�� v� yѓe�$p
�$$�h�����'N"�'��'�N�AV�^�Z[|l���vV-��X���۴���3��?q����<���ɻ���Rp@�9_
0���/v��ҟ���C�)�*zԮAi���B����Dߡ&0�	� �ަ��'��x0��@?�K>i*O�-�����v��unQ�%����O����O,�d�O��<���i�����'}2@� 74D�+�i,mQ����'�b7�!����d�O����OL�ۡA�,���M�4+h\([��QUp�7m*?y��о�p�|��Ai��
�Z�P���~Y�ϓ�?I��?	���?Y����OA�$�a	�7H���!`��y'�'��'~$7m ��I�V�|��͂�������`]���ʱl��'��������$&q�敟��%�<P(�:ef��V�"4��G�7X%����O��O���|����?9��K�N ȗ���;�V���

�v�������?�)O�9o;g$��Iϟ��	z�t�~~��
¢k���i����AF}�Ez�oƟ4Ȉ���W58��T	UY�0(3P.�6@�z�3�F�g�Pqi�O�iڍ�?)��6��9�"�a��ׁ�,��S�T�Zo4��O0�D�O��<��iM65��آ.X����*���:S�7KR��'�N7�6�I����˦�gG�/[���:/�K<<p�e���M�u�iK#��ia�ɯ[��2��O(�g�? l��d�:A
�ŉ�B*-���@4Ozʓ�?����?���?����i��Vh�� �V*P\nE�0��/+*�l�>+��ܖ'}"��d�'�r7=����d��5ؘ�yQ�+&�!냁M�"ݴ�?I+O1�"�sr�v���I�-n�K�m�:O�L�/�牼t�({��'єi%� ���t�'LRab&�^�$ b�e�Y$uJ��'�b�'s�R����4'� ȉ���?Q�-�<5�@��P��OڝM`L����>#�i�\7�O�����t��"���u�.:<�X�'@@A���2cExXI��䥇�<I��'ƈ�dŐ�A*�i)4-��c4�"��'{R�'���'+���ٲG�O���N�� e�E��g��O6���&�O�pmq&�d�'�7�+�D�O���fN��3��цaz�q�qI�vj������4p��g�3O��$YA�xU+��lN�����5S���Eɐ$���&��'�2�����'4b�'�Z�M� j_!B*|����.R���琅��D�ߦ�
� ߅@x�E��ğĖO�'���0����1h֩�SJ*ja ł�_��Kߴ�V&�>9/���䟨��%6�B�����e�)'O��*��`s���(�E^�m]��H�	Qy�$�$Bt��⁐#1���b�o�Lj��'��'��Oc剤�M��	��?Y�(��rp#2�FtZE��!�?���iE�O&��'h2�'nre�-I��Q�,Z��u��n��9��i��I#�Q#�OLq����әS l ��1�dˆ	�U����O���O���O*�d&����!����S���jClR�A@q��⟈����Mk��|Z��E���|�.( ��L_��Ē׭�:A��''�����;!~�����À�2zr�8�D�G1f"2X���G��h�w�'nz'�|���$�'G��'ټ���7#zlA  &K�MKF�'�S�D;�4fp�����?q����醧���9��cIv=3A#�3M��I��$�O���>��?9��Yk4��do2~b(R�dX�]��)�O����|��O�Q�K>	���#7D�̚��%B]���Ѷ�?����?���?�|J-O^ln��c���"�OhM=����&S6�3��ޟ�����Mӌ2D�>1�i�6��A.(��1��&P]jȱ�&c�*�lڗQ���o�w~a(����c��L\��7�˰Ez��g@�Ĭ<���?����?i��?�)����A�	=E���QQ[>L��!��52��S��p�	Ɵ\'?u�I+�Mϻ	M(��p��,eh`	"����u��i;�6��O��S�'u�,���4�y�aHS��@E�
��r�z�J��yҀ�T����	���'��i>�I� v���`��%Qp���´��	ܟ�	͟`�'^7��?9l���O���Vy�H-�(�0<�� #@��Y�`�y�O�$nZ6�Mc�x���6,��d�F�Ѵ��U�6�ȇ��أ75��eN���1�� �������I>��
�`Q�� ��,�	a~���O��d�O���;ڧ�?�E�,HA�QE��LZa���?���i4.����'*�#j�"��]
h���DH�U������	+�'|b�'B�+S v���� �"C
~��$�߫G�e	�
5Hᤀ��F;&z�&�������'�b�'���'�U�p���"��Nt���G^�����ݦQ2؟����D$?��ɺGD��$���1��|ZT�D�S�91�O4���O�O1�x����/��\�W�O�4A�9���9e��p�����sJ��r��e^��Ny�dK8vd� �@Y=�ؙ��_�}��'+r�'��O8�I�MC�*�>�?1@L�;i5�� �-R;�1ST!�?��i��O���'���'r���J8R"�ɶT�Q��$,�>���i5�	?`��0��O�q�(���/r5���ޅ�f`O_x"��ON���OR�D�O��;���i�N���x18m��IF�n�R������	��M˓��|��j��V�|bA�!R�q
��XR(�q�w&+\VO=oڱ�M�'U4\] ݴ��D��(&��"HZ�/�f�ªI�X�tp����?Y�I6���<�'�?���?y@%� J���q�e_-
�ȰS�/J��?I������0�c�⟴�	����OI3�b��S���YJ��f��y��O���'��7��㦅�I��O!,��᫔$3P](�L�j1�*D�B��zy����4�~���ښ�O|p3�I�#] ���lب��g�O��$�O.�D�O1�r����T1S�PXK�+*& p�L�m�(Xn�Or�d�Ʀ��?11Q�$�شF��.^5=Q�(a�� �kE�i��7-��7m,?��I52P��I-�t��f�ץ�< '��s�����ybZ����џ(�	����	ڟ��O��Տ\�^�sĆ�D�8�ؑ.hӺ�����O��d�O�����DMŦ睨{�̘���V>�� �a�n�T��4c����/��)Ŕ&D6�j�h�ƣS���"@�κF� ��~��0�D�\2 Q��ky�O�k.c�:}y���8����  -\�b�'��'%�	��M�w� �?!���?���6R��y�g�S�8b��۬��'	,�P��o�D}&����x���cǎ�i.����7?��
oj��@w�p�'bk��d��?� ��[�h1�H�F`�9���?����?!���?A����O�U;�cR��	��:r�h#��O~�m�"p'|��	�H�޴���y��ܛu�&-[,(�z#h���yR�'�b�'�p�Q�iz�ɁA��4֟� l<��ܨq)�Y�CDG"BJ�	���&�ħ<�'�?����?���?q�iW4��E����a�r&���������b(Kԟ�I��&?�	�`����of(�J�
�/�A�O���O��O1����60SiP@�B�:׎�z@br��6�"?1&+�+-��IJ�	Uy�K�!HX��%+��0���w"
���'��'0�Oi�'�M�R�K��?�%�ۊ�TQj!�������O�����!�M#�2��>Id�i_:7m�ܦ���]�
	�@A��h{T�QP.��.$unZI~�FA�d5<��SG�'��+4"A17�N8��Kä��1"�l��<y��?	��?����?A���c�>x��$h���<H�.��b�,p?�'��-j�F�>� ��MǦY'��զ�."�1�L�>���N!��|��k��)\/Uz6�!?)�+Z70S��R<��b�4����)��@�_y�O|�'_2,��:H25aF��(��$�U����'>���M����d�ONʧC��H�7W�mU�-^��B-�'~�ꓠ?9����S���L8r?P)sī���`pG�T"��"����a�*Y�O��_��?��6��I%M�(���:3?r팤S(��D�O���O���<3�i���BU��3;�U���T�^7��٥�ڸT���'D\7-&�I���D������N�Y����3PN�
ň"�M�#�i��l���i��IYi��r�OD�OMl��� O(S��I�'��.;b������On�$�Or��Oh��|�2̊LC
Ͳ�k_�~�B��P :���%�!YT��'Fҕ���'��7=��P2��\H1Lػo��W re�@S�`ٴ�?�.O1�`��� ~���I� W�ԁ�کS��a�s❧TI��	�"�'>�}&����t�'�ޕ�^�QcFPo��p���F�"�'&b�'��	�M3O�7�?y���?)��S�.�^8� b�P�N=�����'�f���Gd�\�$�<��⊲+�2eH%�����Ig�N~�J\8/�dm� �F8��O�bu�	>"V�)�c�Cf��$.;~( H�c�B�'}��'����̓Ս�NRy)&D��>	ȍ� ���� �4[��,���?���i=�O��ݍ7��� b�J7^6|���M6)��ͦ��޴�?! ���M��Oh�:�6���\�8�ԭcB��WE�y����!ȓO���|����?���?��_-�w��%� ���#spb��/O8�nZ��I����	O����8"cę'h���-M�V�s�O&�������4�?���Sv�XpSD�;�X��N9,,Yd�ʕ0\��rt0P��O���H>A+O��G�?W0���� ]�v\�D��O���O.���O�i�<�a�id�E���'���h�f�,��x�a��3фm)��'�D6M3�	���D�O�7��O�@���Ȉ��B�9x�@�B'�n�7�8?�aH;��I �����Ԣ*
��#�1�����m���	�������D��Ɵ|��O��s��` �-L����,ߢ�?��?��i�2�R�O�z�d�OPQ㇒!a���R�>I��@'�5���O��4�Ԅs7�qӔ�UDtŀѫO0&բ�zu��SUX̲��Ё���d�,����4����O��]�&�L�� f!s -;����O�ʓSr�f���I����<�O�j)2v�4�&��7l�J6�)�O h�'���'�ɧ���
��"���%���W���ʑS�_�S���
����;���U�ɮd���-����1[p��8���I�L�I矐�)�`yR�qӖ} Ab�`����A%	XT}�t���<%p˓-���DI}��'����$.ߡf<4�Pb." e���'��͍0j�����˗����q��� 	%4�8����T���0OJ˓�?Y���?I���?����i6l@��CH4o������@<	*yn�yA|��ӟ8��o�s�������Q�a4PJ��7<2�u9�f��?����S�'M=��ٴ�y�,�MPZ8�!�lJz\�⅍$�y��^p5������4�"��W�^����<G/�P��dQ`�H���O�$�OD�ln��H7b�'�b�k�
9�V�T�J@bR�F��Oi�'�7��y"M<�b��&-S6��1"��W 
ܰ`$�~�cD+]C�s�H���O^����m�	�c�!y��ޯ2t$�+�&@�R���I��<�	�p�IE���'9�@�@�>A_�33$x˥�ml�qQ@J0(cB�j�ԕ��ͭ<Y�����?ͻ�ʅy�`כ3�����$Ҽi���@��w���|��<mZ� ��m��<9�41=����L�8�5/�V�$�F,4`��pt��'~C2&�Ԕ��t�'���'���'Qֈ��$o�P���g �PX�qJeW�s�4or~��*O@��=���OT��c��%>��G�R���:�Ql}��}���oZܟ8���i��E��90I�P`d��3c[�Aq�<������f��a��'ح%��'EJ����]�J�萢K1�ޠ�w�'���'�����[���شP=��;��I��"A6(����E*�z����|k�v���X}R�'tb�'�<����9�\��� �5��kF%�|;�Ɛ�ؒ�Y�O��$����t�zհ��ߧ|���V�S&}���O����Oz�$�O��d5�-{˄Ma�.�fF��k7�C�F�"��I՟�����MK��|���bě&�|"�rm`�?f���۳P�~$�'v����$&	�ś6���ȇ�#� d��h��d)�L�9x�`&���?0�!�d�<ͧ�?��?�d��B���^,m����`�9�?A����D��i��b�ʟ�����x�OVRݓ�W�$�uC6`L�u�
0h�Ozy�'#b�'�ɧ�I�$�����W>$��)REM VpH�S	ɛ(���b���7Tԕ�;K���֯�y���Eo�}�P��;��Q�)��!!R�'-B�'��O�L�X��E.D��ɍ�M�'�2TzT�vN��.��T��N����-[-O��$>���O�ʓ�?���L�S�~�*��Ci����k��?I�,�����4�y��'��E���4%�s���`J�)5���5Ϟ�b��آ�v���'��'I"�'^��'�S���\#�oF�WQ鹱�Ϝz�bM�ڴ;V����?���䧾?�ƿ�y'�	l��<���
�
�<}:������6-�ڦ%�J<�|J�-�1�M#�'�"lKTb��?������A?9�0=2�'!��#�����|[����pR�6UA��NL&f)�|��"�������Iy2�}�lA�5Ƶ<����4�ǀصs���#Џs�~���"d�>��i"6L�ɏf�LQB��2a�Z���oG�Z���f�$���|�$�O ���j?�%Q4˅7f������ϒ�\$`���?���?����h����ҠQ����ȍ��-y�
���D���z3CQ��T���M��wJ(�����'^Y��.L�gX9��'�6�P릍�I56�pAlZA~b.�g?^!�S*=;�Q�4o�(AT�@#o��]��Dɥ�|_��韈����	۟��"*�c@v���HV�,�n5	��by��v�Z��e��O��OZ����L)Q�	�C,cJ��I�����'��iU�������UA���R*�_M@���'C�U2I� ���x� }�b �c�Ny�'��&np<� ߲�Xxr�W�/��'Gb�'@�O;�	.�M��̟��?��g<��`1D� 
?� Di$�����Y�1�?AY�x@޴v��v�'XlP	��Ȇjx*�[l�;�hs�E��<ě������읞R�$����&*��*��Q1
�)|0&\s�>Oj���O:���O��d�O�?%X��5)�������%bՈ�By��'��6�@j����O
!o�c�`�����#�&��^���'���I��Sz��m{~r/،�x��ri�u��%Huϊ�uT����X?�M>y,O�	�O0��O�6O�AD� �K5J�$%���O��Ľ<���i�&i�g�'�r�'�哾QB�[r�ؗ�Ʊ� ���'.�} ������Ir�)��f�<�� ��.�6vF��%]7?nz��"�F/�M;�O�iː�~|��]�L�1�P�'t����F�`�'���'���DV���ߴ1�)�wOE� iޡa�ܤtPx�:eo�2��DD֦��?9U���I�	@�k�i��1�T�jև\+[7������b҂���m�'��ԚG�g�'n+,!D��D�<�R�I4)�0���d�OZ�D�OF���O���|Z�]"[��r0K�!X����Tc΍Rw��RR�'�Ҙ��':x6=��Q�:��y��m�8Pj��O��D?���82��6-j�,�b�Z)A9����@T=(��g��t�ݽ[b��!�d�<ͧ�?�i��Kς g՞Lxv
W�B��?����?�����dS�5�O���	ş����- �4CS-?��m9��H����ǟ4�	}��! �L` �E,����*;��XZ�����M�����c?1��%���7��/���0嘕v�����?����?I��h�8���9����j�x�����N�
��_Ȧ]ʀ*�ٟ��	��M���w�|q��R��� 3�ځZ�����'N��'K҂Ud�����(����>u:�)ǰD-�X�6�I�1n�:%H��F�p�O��|r��?����?	��,���Qc�<���5 M�3*OT�o�[;���IП�I@�П$p�
��X}8pvg���d�Ȧ���4C��OOVUz�W<{s|�,��r��\���҆Q3|�K�OLQYg%���?��H.���<t$X�(	���F�b���r�[��?���?����?�'��$��]�bS������[<�H{��r�tRQ���`9�4��'���?���?A���l�4[�N�5&�@pHA�^/t���4��dS=�������O��̜fH�*kX;b��ȑI�7�yr�'�2�'�B�'|���Y9�B��Ƨ"WH01ӥ�� ����O��D���A~>��	��M�M>Y���9)t��.V�)d�����?)��|���N4�MC�O1�a.'*89�5�۳g��T�V Fr��X�Z�O���|���?9�[N��2�´.b����O�!������?)*O�oJ��	џ|��Q�����r����A�q�踳������^}��'��|ʟ����/oA�rfD����Њ�w�T���O(b9�i>����'�rl%�p�@I�����ÿL�Ҕ��PޟX�Iԟ����b>e�'r�7�����5"��h�:��*1q��ceo�O8��V��?�@\����4)�}�EY���T�>����u�i��6͙��$6�!?��V���	8�$ިt�v��D2�P\"Sd\%�y^���	؟(�	�T�	�t�O'����*��Z�$L8�C�&F<���`Ө�F��Ot�$�OL��v��ʦ�7�<�g	3Za>|��J��lp�xC���MCV�|J~BpH�Mۙ�� �9�wh:�`pPp�Cy���z32O�#4�E�?1�H=�ĥ<�'�?�сՈ|B�("��`o��$���?���?A����Ҧ��L�by2�'�\]r���9i@����>$�B ����J}r�`��n�x�'m�p�v#��%W����bǣ:�BI��O��Ņ��e��Z`�G��?�`��O���B� e�(C0$@�pU�-�V��O0���O6���O��}2��r�䘓�@�g(`z�	^�����yz�vLͅL���'@F7�?�i����@C;�:�3��FEtB�R!f��4�Iᦙ��.ro�hlZY~2F��R���"R��PL���P��& 1	0�|rP�������Ɵ���ϟX3�c+@���9�g�j ��o�|y$p�~0I#@�O����OȒ���D˙H�py��`�"��s׏Ξ#����';7�Q����?�H��8l�p�뢀NI�P�Vn�2�1)A��� Ԍ\�d>\N�	Dy��8fbi�,C��� �Fԯ;|��'���'u�OS�	=�M+5�?�P�ʰm��=C���C�=j�J�?�C�i��O�u�''��'󩋙N�H83�.�af����ӕ{Jd}�T�i����N��2�O�q���.�]�\���T2 [�8�q��^���Ox��OL���O��D<�� 	�(��"+��-�v4d�ŭ8r���؟H����M{6B�|��R�6�|)J�g)	I��I�0-�Mɨc��'t������I���f��H��6���w�@08�`��B�N>�hS�'} '������'�B�'�6D�q�ۈ/���y���}Z�� ��'u�]��1�4I�����?���)\�;���B��Clú)�r�B
X��I.����O���*��?	��B�څαTn7��c�-T%�@K��r~�O[Ε�	d��'�x�dk�`a�i�&^mHݪ��'�r�'?����O�	��M��L�"&?���G�*TR�:�/� W�(r��?�׵i��O�P�'���]6~� �+�j��T�#
�HZ��?�D��M��O
U����N?�+��}�J|��_,#��Z��p�8�' ��'�r�'��'��ӮB���;vfZk����$�M�k��U�4z��H���?I��*���?���?�;d�T���I�8�l	�A[�ڸC��i�:7��O���|����?i�O�M��'V��$�
_�&��a"�2&$F�S�'����u
B��LcR�|"Z���ן��4�F��0-��d�n�����HIƟ���ʟ,��qyBemӤ���#�O����O1x�P�>�y{e�,z��-�$D0������O���2��S2R{J��֥�2xE2�9��ɷel2�2WY%y�c>�:�'s�y���A����,��1�U��聆nt�������T�	X�OO��Yx��և F�r��˿+N��d��1C�'@ȟt���M���w�hB(�&D	�[�Z	31,�S�'�V7-M�U��4K�����4��$Z�Lf^\���
Az�����h��� ��8yw~hP�'�d�<�'�?����?����?��I��dW��h�m�*y��0�����d�I�şt�I�%?q�	k8�q�&���Dnr�;�U�e��O4-nڔ�M��x��d���^Z��g �#-���!�;[s��������)�����i��O�ʓ8��M�5�J%mZb��'hY,��Q���?y���?���|Z/Oo�4a�����+���`��U-�ț`��k��m�I��M���<����M���E{P�Z%ϋ7ʀ�sѫC}\��JP����M��O�qq�+�:����w�00AՐ|�Mk `�&,~�*�'��'"R�'���'0�FI���((Ni�bN�Z$���R+�O6�d�O�ql�Ih�Ɵ��4��|
"܃#C�6\M�s�J@�᷐x��zӨ8lz>���*Ʀ��'���'���_��`��E x�:a��JF>I��6��'<�i>A����IHY�s�-�0iѪ�03f��+R�zc*��ԗ'�6�X8-���?�����s�M̺h*�����rA�!�#�M�<��*z�	��do��T�b�'	������9+j���#b=�p�r�_;!��!���W~�OWDx�I-/`�'����g���D�L�c�hH��U��'���'�����dP>-�'�|7�-G�-���W8I����g��2l��b�On�$RݦY'��S���gӈ5Z���!L=�#�:�]���㦉�ɟn�bo�<!��Vt�P �L�N,�'�!zT��"�\[qnT����[�'����I�d��ɟ���k��� J=iA�%��y��%wD�7mϽ,����O���-���O��mzށ�jؾa,����VCZ(I����l��k�)��$
Ho��<ق��Y	B�f�H;��02`��<�� N�bG*��ύ����4���C�G��Y#�L��4e0v�>̬�$�Op���O�˓_��F����IןX#�GU�@ B���"?��'j�u��&��I̟���A��8Hʶ�k6��X�� �	�U��'���q��� �M{��4�A?�~DM��9	��Ć7,^8��?A���?����h���$ʄC���[@#��᥋&'R���ZꦉPQD���p�	=�M���w�m���	09"4(�
,����'��6���1�	�o���mh~�(K�,������o�E(@L
�8��;�pd �C!�|�_����� ������	柸#�S7T�(�G:��p;��_yB
g� Y�&��O��$�O������=**��5�OZ�\��(�l���'��'ɧ�OR���  �bq��P����/$�j��j�-x���_��
��',����YyZ�D���U��@ [��(|�(�K�G���,�I�D�I[���8 K
Ry��wӺ��3i���X e-P�O��H�pa	`� ��F�O�$�O��|�,Oęl�M��O��e6)�y_���B�(|���C�M��'t��� /�>E�������4���v�P����@��1J�d�d�O6�d�O,�d�Oj�D(��O�nK�+��:��7����'�b�'H�7-2c��O~ilZP�ɕ8O
4�ʺdM�LS,��<��L%��������/N)b�m�A~R%·^P4��_�'���"�Q�$A� ��$��{��|�T��S។�IßL�G�N�+Oʐ�f�2��%�#g���' �	�M�Ɗ�?	���?(�|���HW��m"�CD�}�|D����x��O����O��O�S
DN�sע["���� "�A:���@�D el�y� �%?ͧ���D�����$����$�(�0�X�c�,����?���?��Ş��������å[D|<���!�pd�qc�n�8P��ßS�4��'g���?	Ej�[�H\	�:7��I�.Ǌ�?����Y�ش���W W\����4H1?&��v��&����A�@��y�S�0�I֟���ݟl�I���O�R�Z��D��ڒ"<@3��m���H�h�O^���O����$Sʦ�,Z0"$D�2K��b�cP�n�q�	ß'�b>3�S�UΓ|u�)QeJ0'N��cZ�H!�ϓUv��`���@&�\�����'Ӯ���Uj<��a�H�(�l�ە�'��'t�Z��C�4H�|Ͱ���?)�{�-h�ˌ���(��eIC��2��>i��i��7-�V�Ɍn7�aQ�$���&�3���Y��5�L���@�q'�0�|j���O�0��IΪ�S*޿Ĥу ��hӐ�	���?���?��h�.��U`�T�u#�9�=j�ʹIk@���Ԧ�����I�Mk��w�,�рf� T�R���$ ����'9��iTJ7m�"FM�6�,?�RJ���I��H�t�+�=�=��'׌!�ĀL>�.O��O����O(���O�P�BH��m߄!�D��*G0�@��<a�iФʥ�'O"�'���/�*\8�ӗV&����Ǭ���P��>)$�(c�O&,lZ��M���e��>9�rI8Έ�K%dB4w��@jb��yT�sm7?������ٮ�䓒�J�Z}�c�_�R� B�Qg�4���OB���O����O�˓d}�vO3V�-�N��M0��r�jQjw�V" ��|�v�$�<���T��	��nZ��h@��N)\lt�ئ�cP�(Si˥V΄�lZQ~��� -81�S]ܧ����ز2��`���*�Q��a��<!���?!���?9���?�K~���Z�� ��m��R@�<)r8 r�ӕ����	ԟp�شs1x����?�i�b^�<0
�9ݼ;�i��L4��(����' ·��$k��TC�F��(P+ǅ,M~ b�C�(
�(����_Ry>�в�''D�&�Д����'"�'@*Q3�dR'S�%S�_}U|`S�'"Q��	ڴ^�h���?�����Ӡ����u��9�n�tH�I����O7��O��S�t�[�Zx�N�2 VՈfK��OBx����g���O�	�1�?�!$��'^"@xq���8����f��E�����O���O���<	��i��
fK �5�>MIǚ[��A�`� `�b�'ľ7�4�I����ͦ����ю(�B����q���3���M���*��4��$FfL���'���%<S�2�����Gh�9H^���;	�4A@ѩ<u��)��bP3
&Hs�	��p3�k�7T:.E�a�	V�:�C��Rg�m�0L��<R�!-^>N�f���E��l$Y2��w��I��nÁ��'���W5 �6A�+N+x��UA�+c1X ���;��d�p B�F!�i�� ?�f��(I$��C�!wś��^=E�x���E�2LL+�A�Ad�������pdI�Ŀx+|����[7Q�({p�B�.t`�kwC�Up��AoY�v�>Y��	ˤ%�����r�4�?1��?�'5�O�Ըg�R4Q���
x�^lc�&�禥�.�S�O�"���2ƌ��q�[��@�떢4Dm�6��O��D�OR]���TX�	�|�Ia?9�C�%�6<��-�0����`��U�9�8��<a��?��E��p��,�%C��ěe���>p(t�i�b��x{
O<��O��Ok,T+0�z|Zuk�0w��`Q�Ɲ��ɨjh�b��	�L�IK�tϞ%���A�Ȑ3UKQHD�"d����?!��䓦�D߇B5���%2͸H�P�_�_�h����O��D�O2�%���ʚO��ah���$JE��Zb�P%:����O.���Oj�O,˓h	&!�'w��H�E7[B��A��9J��X�O��$�O`�d�<��,�f7�O5�u$@�Z�p�D[��H�Շb���&���<��-�X쓛�7�B�ھa�� ��-O؀d�iJ�'v�I{jUL|�����2HϨ%��#�Y�Fb��k����P��T�0�'��%�͟�i>7MmM=b�צ&p���E둌x��\o�XyB�X�ZRb6m�u���'L��I&?)�"Z�rfTaP.B�e�D�puh��A�'���ʎ��)�8<��(�B�}vZ�#$�gӛ�	���R6��O��D�O��i�J���@�!��d�U��b�,6
LJ�4�M�Ea������G��>$;¬W$r�Y���E�90�lnʟ��I�|�!(��'_�O���ᖧ/��VdI6_EH�+�����1O��d�O��$D�? 0�3���<M�`=���^�>�Ҭ 2�id��S7g^PO��D�O��Okl�[hY)�l#$�
&��Ɍ�zc�P�	����Ipyr�5�ttɢb?U�a@R�VW��X� '�d�O���%�D�<����}��YI��8�.%��A�:z���<���?���D�2h:8�ͧXt`���ɷJi��LíT�m�OyR�'9�'NB�'؂=��Oh�Y"U�U��1�gűl�J(seT�l��۟<��ky2B[�<����?Q"d\6�!{�LR�q䐢 �]A���'��'���'��<����8���b��tZ�݉� H���6�'I�^��¢$C�����O`�$���h���O$����.� ���s�ٟD�ɃT��?9�OO�HBtd:_8��0��^����ش���L�P�n�؟\�I��0�������©R�wA����1�f-��iU��'5�H*���>Mk�I�g�� ��˳ᖧb66mZ�LAnZ�|����l�����D�<Ѳ�'�1x���Z�t�i�H�r�vM^).�O2�?Q�Ie� �#�$��\k��-mu����4�?���?�]3C�L�';�Iϟ$�q�\�c �9�U�@��Q��mZS���q6���'��'��7cM>y|����p�  B¦q�d�$�]cB��'i�	���'hZc�qAg�
j̢Tlӂr�� ��O �C�O�i��9O��$�O����<���<B�2�匰��́B���"=:��T�ؔ'�2�|�'��-��0S*���E ���c��^7춤SS�|��'��'K�I�j��Or�¥d��U=�գ�oL4r�4�xٴ���O�O����O>��Ө���i�J�����E�!7���ƣ>y��?�����
��p%�Oi�J4T� HJ�7N������L�6M�O��O��d�OTEJ�)�I$8�@����<n��2��;RB6m�O��<QwoY#�ǟH���?�a�/1��p���-N&!����ē�?I�D<����՟�����:@�Ka�1�����i[�I$z����4�?����?���5��i���Æ�#&p����&�!U2s!Eh���$�O��9$��OZ������}�VJ�$R�j���͌5a���M�I��o�˟���̟��/��Į<�%i�_� ��G�	g��ݒ�C͈"��fXf]����#��џl���
��:t��Z��Ƞ�#E/�M���?��)<�����x�Ob�O`ղ�V�>�� �j��Y3��i;Қ|�
�~Γ�?Q��?����  (^��T��49��JU��&�'l�B>�4����>�$ 
_�T)���}�|"�}1f�f�	ʟ '���	Ayb�'
�X6���'����&'�^�DD��(�a��	ڟ���r��?Y�'{�-��п)�t�KÁ�[�@S�4z���<�����Ov��¸?5K'�B�qX�;Tj�c	6I	�oӰ���O�㟘�Iyy��Ms 9z�|�0I [)r�H�o�Ο��'��
�I�@?��kF�4�JĲGV�Cj�tv� ����?!�����5<��'k\ sa��
���
�[�j-�q���`�'��G΍���4�	g�{Jέ�� ���`�f	�w�v)&����Ry�	7�O�J.�}��EC�;�ԘC0�
���ԟ\[a�\ԟ���џx���?A��u7��5)���s��I�Ę�d�M2�M���?�eنLh�E�<�~z� ���lL��g�(Z`�����qT/�$�M#��?1���3�x�O`�ňDNѝ8�T��P�l���d't�~����Ob�$�<9O~�'��pmӋ}���E�-`�p����r�����O��$ɻw���S���>����G��=Xd�Y5���P�0�1O�����_�����	���7�Y)�Y���M�zM���ʇ�M#����x��x�Ov|ZwP�1e�u�X�dJvQȴӫO�ˤ�Oh��?���?�-O��k�([� ����X�婒%�[ E��(�c��ȟ ��L�Hy��8`X`��eO�1� +P��,"�l����'s�������ܟȕ'��0!�f>��!P:E��5�@	��>7`��>���?�I>�.O$[���O`r�($t.�XQ!�/�jj�-�C}R�'�2�'���-0�*$ J|I�F#L艐IJ�{b�8�fL�H���'�ٟ@�']
�X��'J�'/!\�I��(yeM�l��;�o������ay��F����$��kLٴa�����j�����z��R�>�'4�ɣx�
����_�(H<f6�y��2�f�� n����'� �3�oe� ��O��OP�XH(�B�3��	ッIz�mZIyb�ż`b(�=��'�
	��ߏW���a�w�Un�)i 0�ٴ�?����?9�'r?���tHc��0K�*^�^�d9�+N=�7͑�|��$�Oz����<)�wP�px�%�Y�p�iL�o �ˋ�M���?���V(�&W���'VB�O�����Uԥ�	M�h<�F�i3�'�8S�����Oz���O`x@��_Z������!%��X7A�Ԧ���
>�6u �O���?q(O����^�@t�! �K��	�-f�!�T�x���u�x�Iٟ��	���Wy ��'��'�
r�a�n�D~dp�%�>�(OJ�D�<���?!��� Ӗ� ��dK7��>8ޕe#��<����?!���?����^d���g�? R0j��9�L(��]Q��*r�i��	�Ė'���'�""X����3�d� �ŭm�4�j�'ٺt��v�'#��'9�^�H2�����	�Ok�<*�t��B�+� �"v� �V�'��I��	͟����g��Oh	���I��$��c�/L�,R�iE�'���[�T�����$�O���M�2}�h"���L-��8�M�$>( �'��'�r�����>����p�WoR u�h��υD�m�]yb̎�<�(6-�O��D�O\�)�E}Zw���(���o�"Ѐi�*�
ܴ�?��uO�X��?��B!и!��$g]+�0;��Ӡr� )���,�M�'�$��'H"�'��D�>*O*��rj
72}��e�;kܤ|֦���h�4��Ty�)�Opk�!ǜW6X �S烳:��"�OǦ��	ɟx�I�:��OX��?��':̼���V�[v���G[�Zn�0�4��d��S���'���'. i+�LYu�]�Ǭ��;�%��s�����1	�h8�'&�	ៜ�''Zc8��B���5���p����4��O:���<O\���O��O���<��!��}�����؛{*n�F��d��Y���'ZQ������l����,82�S�A��(��}\��6�n�H���|�	����Dy�ՕWV���d!rb�"@�
z��W;C%�7��<������OL�D�O�Q�7:OȺ��²S�4�P�D�26ϚצY��ȟ��I�\�'��dm�~����^9z@ԙ�-V�N�*V�զE�I~yb�'i�'1�L��'�:��io�:&�,���#45��m�֟��EyR�U��ꧏ?������X�Ŏ�gr���ÎÀP�ER�8��ޟ,��<���I��'��)��i
��͋_ڰ9Q%�Yg�&]�<`��I��M���?����J']���7��A��l�6r��a�C^8�7-�O��d
?[��<����޸O��A=PC8|��ڽ>�@Lk�4X�
<H2�i^��'��O�@���$�$8�������LK�x���J�n�4lZ4<�d�	џT��(y�"��2�'S�̉3T�F9����eEC�|����i���'���ƾV������O��	�4*`r��nF���0̃�3�D6��O�˓	x���S���'Bb�'*dx��ڟ>Ό���-t��X�$	oӲ�ċ7�l�'���ϟ@�'�Zc ֈ#�jJ �zq	�A"7Z\P��Ol�!S<O���O����O��d�<Q#�T#8r�|��[�a*�Ȓ�U�H�1BW�,�'p�Y�(���������/�+r2�fE�1W�����D`�,�Iٟ ��e�����Ry�@l��3F�b��ĔO�v��A�R-MZ6ͩ<�������O8���O�-x�6O��	��.z�~y�T��3��!�N`}R$-���'q�	�*�P�O|��KF�6�L����U'�Q�S�{����'��'���'b��u�'t�~�z@8
H�)O�d��פ��]n�Ɵ8��Syꇬp�&�x���Z@�V`G�i��a�`G��o�L��7,^`��⟜�I	���	{�	|0n5H�:�Xa@]4�Y@�ڦ	�'���Bh�,��O���Oт�,�m�ъ��RX�bƮ^%��n�������#<i���˅08va��5-����Ύ�M�̎�"����'`��';�ԋ2�D�O���d%W_�<�(ӫ 
n�pX���֦�P%E��$���j��E�u��(ߦ ��	�U�D_�9�i��'鞬'��O ��On�	�{6���d��3��q����[��7M!������?=�	�\�I����#F�	�H����3*���:ߴ�?���P�nV�O���9��Ƹ%�Vm�+db�䡡Ύ�0N�9�U_��ac.@͟��'�R�'sbV����ȞG6��I䡕�kS*�C�B.D���jL<q��?YM>y���?Ygn%��0C�AĎV�ԙA��~��(�������O���!�i	�l�*t�'X�0�0qoI�x�N�[�
Mr��'���Ky��'Jr�'9�����`IKU��=�v�o��	A^�����@��Hy�BP�#��Pˀ�A�O��5�O��I[̐1������}��럴���y�pa�	Y�Dg��
�aS�y�\���ۙE����'"_�tƫ�3��'�?i�'g�t ���>�q�G��hhlE1x2�'�R����y|rԟ&�[C�� ��0�]-UdI��ij�	�&�h��ڴ��Sџ��Ӆ���c�YA��_ 1��-��C�$����'�R���R�|2��-	�Ĺ�n��l���Qɝ00��!ͮ��7-�OD�$�O����z�
ꌩ�'ǅ�"�bȱu�6|9�2�i��9qB�'��'���d���M�IVU(�!5!EL	�l����	�Q��ē�?���~r�ͽ��t��ҺU��!���M�O>�#+�z��O�r�'�b�ǽMl� ��gJ`�4��o��27��O�M:�Bf�i>FyB��&�8ѩ�"�!L��T�����Ā,=*(�Ĩ<����?!����DW�F|��!h\�k���p_+vȭ���n����F{B�'�օ��/� ��a��դ2�8dj��I{�bP���	֟���Ay���5V���YQ0��įr���L�&
�P등?��$�O�(�R��O.<3�1��xʓNB�	B؉��h}"�'V�'��	)q5���K|R"㋰K��`�%b�'�AAA�55��v�'��Q���'T0, ̟�I�`v������N��6�
�So7-�OX���<��0OǉOB�OV�� |��t��'^|aq@J�9.A,dK�i���CyRc�������s�|r��M $�����o\�a!^�y԰iO�ɉC����4W�Sҟ��S����#P�6�:�.�mɚ�yB�1�Z�ЊEk�s��|&� 
��%Q�����ȕp��E�~�R��6����������I�?�O<���0�DPS��B��I1��LR�bC�i��HR�4�1O���E#TQ(4��%R��ғ��<:*n�����I۟�.v�'��S��\��8xx��9hN-�DH���qt�I)��'�?y��?9���F�lY�p�e�}��E½(ڛ�'V>��"��>9�]?Y�Iḩ̌O�B�A='��1� �\}v\��x�|�'B�'���'@f!8SC�8���HF���\$��*7W3'b�'pb�'�r�|r�'��$��eۄ���-T�P���K�9�F�D����O����O�ʓ|�b�Sv0�N���X�d`K'*�f������ix�	�x�'y�'����y���h���˒l�9��aΘk4�6��O ���O����<�,N6<��Sϟ��i���X�#7v��@�C�f7��OZʓ�?a���?9J��<9(���Z,h �4�={hJ�+�ε�M���?�/O:�r-KL���'���O�d�1e\9s��yq�P6��$C���>���?���м���9O�Ӡ!�r,��	�4��'�ڣN 7��<ᢊ�?~՛��'��'��D��>��+���'��9Q[���� �3E�v�m�����ɏ}�V扬��i�.���>��7J�"�~�(��Tz՜���l�$�<��'���'��D�>�.O6��Ί"����Ҧ9��@ڂ&�Ц���x�T&�T����rX�p���Z�L�0�U�m�#�i���'G2�������D�O�I�!'*��7Z�j�!��"m�7-�O�ʓVwv��S�iY!%�S���T�Mc�ՔK�tU�0d�IL����6D��
H�G��!r�_�x����4\O~D�g�ަ�zUcu�Y#N*
��a/�;�Ly�fH^�y����b ֵ �
(P�N�*s����&M]�%Z-��-�/��S�MU�U�,��&ۯ4r�-H��H�YM�Ma6��HJV�p�ݏ>y�4x��|ǰh�e�J�S�M�MQ|�
�
�g�aB!��'H�k�"�6O`\8�r��Y輩���'=�׌+&��'>�) -u�u��Đ�`-�e�����q&H����a�T	#�|����[�'�t1��
,�VƇ5S��V�AyL����D����6�h Z��G	>���4����Ob�$�<!1kآ�n"�h%��!�тOj���=G+�\��іe��q��.j<鰴i�޵Y��ىQ����V�[��B�'��I
2d	�O:���|�		��?�ԍ];���(G	䴸�nP��?���:!J 8���H�F�1�<�*���'F9����B?m��=���W�����O���S�
�Pxa���I��#}��zag�	����s�i�+�ţ(}���<�?���h�����S׃�ts�q�*�i=!��N�zX }���QQ��0p�"�ax�$ғ)#`�P!Ș�UG�8�D���1q�2Z���I��p�P��iFP������	��]&p$�a�@�=l	�R)ϙ97��3D�T�c�`��}�8���f�g�8%����VE"ݖ�ӕ�0�j4b�(�_9&���u�֥�4�"�3�$��)E�]�!$UP�:���v�$>?)E�ޟ�p�'����肍:V�191�T�cS
�b	�'��$�2LC%}��j���P'X���O$Fzʟ~ʓ6�j�Pש*>}�h�fnW�z+��H�*�x���b��?����?Aױ�����O���?+,�zgj˻��Hbp�!jy�Z⟷@�h$���6ײ���#w���tǓ�7��Y�B�^|��%�@+~W�x�he*�Մ牪WjxQ�.H�;9�-����q^P��O�O���=ړ��'�0���C	�x��N����'~JE��M�,��Df��6�ɾ���<��-Ī_P��'a�AV;H�@��n&<�V�ڃx[�'�t��'��' ��HŇA:^Y<�����LU�7�$�@��P!�2�b�����@��x��� �#d�]�ܭz���'h��	2@�=ǈA4
;k�6��e�����O�P �'Jb�v�v��Ɛäs�Ҥ�!&M˛�b��?q���S�O=P�i�L�?�dk��=f�j���O�=�|��i�*=��Ed�f���I)_6U��r�\��J�	�5�UM�D�O������ؗk�Oh�����D��ɋ�H�p�(�O��DV�@�b��G�Z�Nɸ5�i��ʧ���5,<  #lD��q�1�	>5l�WL,�Ue�OJHL�����H�2I�U�+�-���;(��2��>a�+�ӟ���j�O��32N�Y��A��c�@Q��#8A-��߃1ZTAw���S�����M'wfax"O5�k�P�Hg�՚ym��Xu�0j���V_�����d�c&�)-�R��I�,�I��O("8:s�U;lZ
0X���N�"�� k�[Cl��`�smX�\��b>�O����' =�E�FLD����D뜆!���cA����X���{�q��'���䞨U�l��K�T�����'s��u���4���$9�)� xq�kK�p�|�K��H�4х"O���Um�X���P����=@��j��4*���?�'g�4pFk�:N(�#+ˍ�ހ�v��zI�%��'���'GKh�������ϧ'Y2���
	g���̀#iH$j�o�Q<�  ��xǮ]�tƓ�b&�u�ǡ SMV؇�{î�8��܅cc��0,2_蝫��Ο��	�=���Cˇ-l+����u�B�Ʌ��2c�Hf�E��ϗg̈c��	�}R�	ek�7��OT�$N�Y�4�*q��:ad��eǝ�H�J�D�O<m)&�O���h>�S�M�Op�Oze���א2���2��,eLK �'0��h��)6����,�Rax4�� �p<�n˟�&��pv��0�@��Ѩ�*96�r�d1D����A�Ͼ�[�$O�t�έV�-� i�42R��1�)ژZ޺�2�!����<�'ؿ ����';�X>m�"�Gڟ�QT	�+rj���4F�-(�eӀ"R؟<�I9d�Yx���=N����	�|*�+�$	�2@&C�o��@��%Ec��t�i CǓV���0��͌s�gk9�)тÌˁ閅;�V��v	طpM�
v�����\A�4�?�M~�����9�ǁ��n�Zb �*dy�9FdC<\��̓�?��S��<�.Oε��K�~�p���O?��=�t�'Z�B��y��i��@͏3/�%��A�Vpj�W�]/0�6��Of�d�O��a5 �6dgJ���O ���O�n�.��T� j 2���e�T�Tc�����%<Od���׾#+.�AMGhqD\x�����F�y��!]��P�ճb�0� W���
1O>� �����1��0�"Ӑ������.\�lM��O��@�bR�dN�p��C��y�'�6#=E�$d�=�<�PU��8nN��JG�j[�c��5U���'���'�>���H�	�|*�	�Y��`�u`!���a��L�o��م��z�.�JT�I7�֥K��_�E��3��q<q�	E��U:�&F�:��!`�ʣ0�0�	b���1���u>4�2`�a��`�*D�8z�`N �L�q"bN$z 윙C�:扛��'���K�Fa���$�O����	/>A��)І�6aH�*��O��@1ym����O\�Ӿ	-���=�C̤�c�ڋC^���F��(g�x�.���'`2��I¹2cg�)sV���p~4�IX�I(�Xl8eŅ��Uv�� [�C�I;|,�
S�2V������T�K��C����Ms�*0c�-��G�(�9���f̓�n�־i��'?�.�4��	�t�!�]J��d���<����Iϟ�W�U��<�����"hb�8T�_�#N����Υ &�U(�Ex���'C�q��-Jҋ�lZ�j�����4	��D7�)�SE��C�lY�F���	�#�9a�<B�I�(ǒ�[@���C�¼�N4<����}�'l�T���!y�9"�؉(�h���'�U��R,.�@*�����p��'44�p�Oj�|90���>
T^<:	�'|	�t�LD�T�a(H�J�<��	�'�ԅ��C�k��L����COd(k�'�L�;��
�8�Zf��NV�y2�'���Z���%,H������M8R@��'Ң����	�Ԉ��dK��P;�'����Î�"_��%�d��(F��ݫ�'�*	(��K�C�R�[����B�p�x�'\H��)űc(ҍ��E�7;D\��'a��y��E:躆�`AN�X�'�|�P��!G���ECy�P��'x�,�Uσ�'W��O;&�`M��'�ę�F�.Nk�8f�Ը"�<��'�6�YA⇎pk�Pd��Lt�;�'��呑ǈ*m֐�D�(v`�Y�'T���D�ڔ�4��ĝp%r1��''&0�׎��%ڌdA�M�e����',��jD��$$l��:�Ȉ�aQ,���'�Ң��0�a�D�0l�~p�ȓ8#�DB,޳A��!�ͪ�̇�S�? �P�&�F�T�b5W�Z��*�"O>l[�&�p�]���B����A�"O�-���.Li`�hR�U>8�=�"O]J��ܔ+O�H!u`��Mؠ"O��M�W�Y��C55�J�'~\󥦊�:�p����y��xS�'A�)q�jǭ~m$��B��q^���'*��E��1�d�l?nǤP"�'/hq�pd_5�*�Jg��Qe�y�'����� -X2�'+Q�w�P���'l<�DnI�_v����F1o�T"O��"p�:np��:$�x�H�"O�1"����'A<Th�#�"m�,���"O�ay�H�L�JŅmۈ�	�"O(�㴀���
ѸJj�]CB"O�I� ɕ6<P�贤Ki�9"OZQrQi�
�����@W���"O���C%�+L�1����2?�8!a"O�D1��}]ܸs�L�G/ƴY�"O\d�SGK�<�p����y�"O �g;RK�A{��2i� 5"O�#��&ژ�XB,��lSp��s"OPXRȎ5~�웕k FQv��s"O ��WO�N0@�?Eo:-pa"O�P��E�;쌋D�E/drY`b"O��Q��q��P�@�o\���"O&ـ�D��O�z��$��RQ���R"O&��kerL ȧԵM�ȃ"O\Af�]�Klp$�"���# X��"O��HR�~����^�����"OH��W^(Z�⠘D���X��Z"O���E K��)!@�]�w(�ax"OP�0���"ꦑP��{-��E"O��k�c���<ڷ�H�dd�"��D�Y�F��W��~�Ov�|��D�X̑��g���r*�'��yW��*b�fe�V�ڱ�=�� �s��bo7}�� ��� SN�e00�U����Z��9D�(�GńG����׍l��xKS�O\1$Nв,�h��ۓ���ʕ,�F@��Q�ӄ��݆�	��.m8�(ܯ{͛fi�OU�i���=\�Pѓ���yR ��N�.(�'K�1MP���.T/�~rIAڎ�I�p�j�j �M%m�>u��"��SD((1CFR� s�졲K4D� �#\m�8I��f��(����C J8�Ր։�M�͈5O0�'$c�8(�H�`B�@�J��6&ʴJsñ<1�i�)=:�O�S;S���-��(P���[L��1K[Ĝ���?�1����İ7E-lO���G�7~�ū�W�BdH�yԖ|bV�FlX�{Ю��=4�p�K~:T���0�ػZ6��[Q�^(�̝)4�[���Q���9 	��F��{L`������PC(�(�ʽ��6?��$��8�>�ɝ(��=�ԃ��2��X�j��E:>�?�vlSV��b?�1�T�L�^���^a�}{p��OH�����1�����'x��p��{ap�H'���a; ��O���Ns�Ӻ��F Cv�U�2[�D��cmj��ۖ�Y.��s�"O����$0Z���n�DAB5�B�$A�M���3&(f��|b�`G2H� ���B�E�}�0�|�<��'��ؐ����.�&�YDh�;��d�)���	���G���O�1�������.En-�Q"O�SGF�V��#�B:I�A�Q�`��kq�Z�䡑�C �E�QO6ړ6����0��<��t��ׄr�*��뉗xx��1�̈J��)�k�!a��qX� �줐����R!��a�5� ���	�#3�	��Π<�npYcf��fA&➬3�LU�`�p��X�U��r��>�������:5�����o��A���j#��9��Y�@d�� p�5�2���3X�ԲdT�^���,Oq��-i�we��0����*.�J�#W1�&� �'ڲm���
���H�*ʮP&��"%ڔ:����垫`-��ajN
oҢL����(�O� >к�ICm0����\9jP��'�����X�8aC��ƍ8�����<aCQ��t�1G��-A�����T��{�e5Xu�Q2c�6]�Pݻ'��'�@����,"�Fq�Qo3�fiѡŝ;B��b��O�^�Th�x�,��p��?p�n��'ɢ�$�,6i��O\$k4*�,K+B����i��L�D�«�)uI��,*�Gj��ђ`� B�ıH�*��JY!�dwA�♇W�fѳ�(����g�~��X:`O�pI���f��3★S�v��>��"�,~~6���gn�� 
�0=ITF�1�VLІ0M���0T���J��i��a	J�z�E5ݫP �����'�f��)�5J	2�H�"���K�y��I�&���Bl��,��S��԰`3�5(#�dLfם	[`���6��z�t�xr�Ș��B� &���0Dɤ �*�hP�Y�( "j�7ɄM��R�F�`���� f*��2O|ⷋԼc����?>\�$����8���ID�<Iw
�P�b��A_�?��Չ`�
�0/`CQ ׳+����bO�HV���
�T�r<�&���s4��D�F"8~�����o�az�#;[�,�F�������FO�&�\-x���l�.=ɖ(!��h�Ţwq*���'��!Qϝ�bD��&�K1Z6H-��y��J3�X�@�0p��(�H�;-���a��"<���ܺu��d� ��bm�#ή�ybʌ�i�*$o��E�v5c���X.ܙ�r�S0uq�yZ�eG�q�
��e���On
�əw����jI�^S�V�8ɁdK�<1t������
`�H�>Lk�Z*7�I 3Ě��d�H_TB8�E�E-Al�OR�+�yk����Z��t���H�Iۓ3N}�4+�r�>I�� �-!CT����".�F����;B��L�L4c�S/O�'���`��ͤ4���@	�cIN̲�}b�H�S3��`�y�MH�O,IP�T>�kW��6��&O �!}T���e�<	�̚>�0>yd�4	s(���&"Ёc���0M�4��K��h"e*=h����K���n�(|���������� �I�!���1oF��Â¥iz�ɸ�GO�u0��~�(]��/��+���Y�	��5�F��=���wo�!��jLvq���*̖h�ߓ;]�<no�&8��eJ�9$�����k�h	���&��!D
���̡��cav9�P�ѝm���x��,��#<��m�[F��p���{[���&����	����Ɯ���c�c��C�	�&t�Z�#Z�{ȡڔ�  ��ɏE��������Ti�f�Q?�XP�-I��]I1eEi@У�,�Oҁ���z�ceԟK0`���HÕ�D�q1Ć7u�F�� V?/4]K$@�=W�lyQ+�� ��jW�	+|P1���3b��e(�ۆ�ߴZF��*Ov�I�&�K'��z�V8A�c�_���dJ��42�M�3`�s8����^a�tx �	�-7n�C�BD�A^�4�B�%fP`�0u�FT�D�O�0໩OD杰�<d\�1��,���"T B�I'�&r��j�����/K�9��sVa2?I��V�3����~9��%�zhDj4�[��;7K��0)Q�O¾8%r��RY����!�TJ�أl�lg�)�`F��lbA ��e:n,�t��")&�Qu �R��XY���"�j(�f:O�m`E�Wy2H6H�NݙP�A�[�H<���O@!��b�
P���5���xwܐ{9O��Λ7S������0b�`|	WC�I��{7͏?)!�'=d�d>�n��� kS�K��v��z2J��AR9@p�T���H=�zL�!��ئI+Ɔj��%�T�itd���Z���j��c�~@��Hź4�T[��S��V�z��1�<��0�N� �����"���Q_<7m̍Rg� B5+�!!�e���_���j�;�<R��Y�%�K�mY��Y��^JpJ@C�I��P֌K2z"΅���]2rO��q ��"&�prK«a�
`qH��u�¹*�hS)c?4�X�A�$��'�Z9�!��P}rk�`�T�Wi_�w��KtfG��O��W�����
�*;Z���L�<�1�E�cfY�7풉#�r���4g n�{h��{�>�x��O�C����O�t҅ƕ>)����&}���cLO����-X�m�1�qF��ąi��#��$y����s����ʇ3����˘`�j�d��8J�\xc�'bt�c�I�a?�z1jУ)�
)V�x��ݛqÞE��I9��,Ȑ[�Ȝ[��I�t��;k�1�ŉZ2l`M{��{�Z`���kv$��b�fz~@�F���DHX8V0C� 5]��A! �Ә!���i�bA�'E±*ũ�&n<*�U�������Hy*�E�L���Vj^9 DL43Qg�+_P$��h*�` �I�dv4�/DZ�`W�eA��$�L�23�Ğ&?�`�>�Ё��;�P�8D�4�T�&�/D�@pfR�?��xH��T�V��e�����;��S�'�� J<E��� ������f���&�y���W���t�	�L��I�����9�K��!,O.�[�c�$�r5�g��8�
�R"O� z��Gc�:�@��`ؒN�Vq��"OX� ��>oS:`ŨH	J��<�"OV�����c���J�D�,i��"O�9�G/�ZFv j�@�:�r�G"O��x��4�(ep�.ļG��D� "O��
�h��@�h��a�d���"O��r��d��q�M��@��"O��ă[&4��k��I@���X#"O���D�fwL�����W��Ԋ�"O���鄟7������4.  �۲"O�X9J�?U�FU�����S�f	�"O�	p7 L;5��|�F�h�6D7"O��j�eC�o��}�SdD�=��eS�"Op��c]�2��֬��j��K�"O�0H� � lu-``kŗw��z�"O�(���@�:`��Ѩ�N9�@"O ���56w���c��x�b"O��I��Ģq�HB��hl���6"ON��&EZz���!��)R��{'"O�jЅ+K�J�ZA�]G9j�Cn�<A ��)��E�fA��(��eNa�<ٖB��C���@�fͺs8hh`�+�^�<�W7�:��5[,2�[7@�C�<���mBʈA���R���S3�[�<�Ł@�N��s)��%(����V�<w�J�X��IM��E���LU�<u	c}�K�Կ	
R1��NU�<�WH�3$��: MʹFRAۇ�X�<a�"'#�1�E�}�
����Q�<R��.3f��jsA�2\�2Q��
�K�<��d�<t� �	�1��r��C�< Jרt��%1#�(F�D�3��BF�<�T�-\Xbe�ů��U�b*�h�<���)_��HևĘ!(���k�<1���6����D!�=O�@���ANi�<a��]~�Q)��H�	)rJAe�<i�OʶH,�xq��m��y5�a�<����PJv!��kQ0n6����VE�<��DoF�ғm��g� �p"c�C�<���Y���4��{D�m(�V�<ade6)g�#��Æ M�<q��!	!ܱS�j%A�6��7)�L�<١�U��X�w���DD𐃭U_�<�u��~�8Ie�ߢ!�֡���f�<� )Z\���b��+���a��_�<1�	��|@�����H�eJF��aKDQ�<�5K _$�Ժ���v$��q�U�<1�b]�E��@�ّEy.pub�Q�<�E^x��A���`�r��-�U�<ل�ƢZY�|b�ǔ;e�"��$�W�<q�e&`�(����K� �) n�<і���+d����W �b��s��D�<����b%4E*#�ɰ10����jF�<鐨��bF�D��)L�Y~��+bĕT�<�P��Q�gK&6:m;sj�d�<���;>�Fi��p�`=sBGf�<����5XE܈{�퀬H��4��GBd�<�Q	�i��$#��ޫ\�l+'�w�<!u�(n���P	Z�{WR����G�<�TĈ�w(��� .BE��O�*afB�	�ZIzh��,X�z�>�(�FMO׆B�	+�.����$#L�8&j�OfB�	�I�6�UY�[�p�	$EͩA�bB�I2d1|d�l���u�b�n�|B�)� ʤ�2��^<����L�	_��"Oh�.�Oͪ(��R�U L��"OX��LH�zΞ �@
S'$@�@3a"Oh�����0���jQJ�
;fy��"O�����2A�M�!�ďAʰP�"OPL�S��=F��Ya1��$ty"Ol�3
Ϙg�� ���+��%PT"Oz9�W�^dv�8�M�{�Ltp'"O�@RA舑��eS���D��Ԫ`"Oh0fU�N+�t �'����"O���Ř-�px"g�"k~5�"O*T��\�H�Ha�#i>i�A"Of�y�gV!�%/ZF.xk�c�>�y�ŀ�tʀ�A�U3R�VE���y2"�9�T٩&BȨ;`]c�`A��y��X��d��X�u`V���(�y�dʾ;�I�祈�?��"����y�N�YӢq
��[F8�4��R��y�9*֩h�L�%C�"���c�
�y��S&��̣�L�5�!qb)��䓊hOq��	b��8���褦_�<3���""O yȆMW=Nvu�!���d�@"O�i�c�͐�Zd�gD�;`�tXѐ"O�a�&���K�\��Ө 13*@�"O.�&k�%hu҅��'W0D��"O���A6x8၄�rH$K�"O� �4ݩ��@���B+�� 
0�IB�O
LmkBH(Z�E�c�aY
�' Q��_�h�}��%C�I&̀	�'M���)�+qBI�P�Y5(�d��'��XcI	?&�V}cGM+@0rT �'.��B Q6�D=�W+=X<��'�z�ǡ-Yɤ�"�F�6MH�i�'|�pᇀ��C�$������H �'�Z)�� �>��[��1Q�9��'	t*r���[7��X�HUK}����'�ll�&!͟h�h1U�K�
��y�'��)��\6X�J���܎}� �
�'El0���W��l�a�I��h��	�'�2�dK��xT4�Ƃ�� w0��'��8�C�x���ꇯy�\��'� 8��肃Bj���ą��nLf�'��SK�/9JRsD��h�h	�'��c�1=�*�C�]�����'��a�d �(ݮu��8W�\��'ڞ�rsH]�h}>��Ȟ�V�5#�'���� �Jj�1�M�c.%;�'��0�3J�~A��a�!W��u	�'i��E���84�1�A��I� ��'���sI��s�ܫ��xjl	8���'Ъ��k��c� g�L���c�'�1r��C�Z_�вA�3G�V�y
�'��Љs͌6�������DX��
�'^��8���Q��P�1��5E�(ێ�� �'b*(Hvǔ�o(2+Yte����n@Q6��	�"DY��<����ȓd�h�p�vu�����%x�z���"��c�j� 9潪aɚ�뒐�ȓB��	ce����9��'�T�dE�ȓ{Li��h��D�4:�@��(�H��DN�XBw�j�:� I4L�M��A_nAã��$j�H�T�Ђi�*5��U�,x���@�¼i��H�k#t��V�(��"h�S����(Ԗ_Y��S�? �%h�� �8�N�y"\�"Wj�2�"O�9A���
�`�C��QV��"OjH ɖ�nr�U���Z�5Gd��3"O�2R��\
��:� �o+�%�"O�hR�`ȧN�j%bMH=E�j��"OV�[�\a���_$rn��ٕ"On�3�+ǿ+�H�`^��N�`"O&q�"O�9��`+�� ά%iw"O�*Į�6i�VKbҬ��%C�"O,�Zp��26\�,a�ʊ�Q��� �"O�q!�^�g��	#C�3�^�����6lOB��u��&'��yV`�0n󈐋4"O�|R�i�+/
 �qaSڞ�� "O0�H�7]�4M����x��}x "O��
��H,@��1�$���z�"Ob���A	�t�d��։ѣ���Z�"O^D�A����9!d攷,��d"O(����P�kZ$���&�*�Z��d"O��)1� t��c�-g*t��"O(1� ΨP�}k����佚"Ob�bfd�_Q���� .-r����"Oz9�Gb����K��	�/����"O�8kV(ʰ�10o�7Y�tȔ���r����> DBԊ!���
?��&�>�PB��6*�<��4���&�M!C�� h&Zc��̓հ<�e�798I-Uk`��+#]�<4��*qE��9F�ғO����R���xb#�\:��8��	�R,��#���0=���� 4㠼�tȓ��AX�ʀ��y�L�L~<1%͌'xb8t`����y��6yo��a7 �ET�-2q^��y2OA)%��	#KȌ5�~i�U��y2 �D��C��� Px3� ϑ�y2/J^�EI�$�� ��蟤�y�A�^��Ay��yt�����y�&� tb�
C�Ǥ`�l #,$�yb,��U�����<V'��)����y2�Ђ0n��ӵ��4H�t9�"�S�y�E&.;l����q���`�����y2`��)�]R$�q���BÅ	�yb�3��cKT�m�`81���y�BT��
��2え6�(8�`�5�yb"��XQ��aF�[y�xK:�y�� ���B�(JV��37���?�����\B6���) (�y��B�]���ȓk)�M�AU ������H�&ք�ȓBPr K�C�3n��8���c怱�����pkD'[u��0�`'g� 4�ȓP�f�&����	�J��G�w�'U?�ɹgu��i���\B�z�
�5H@B�
�Ҁ+�����F���P�lC��4R�\��2�ɡ%?�@�a���"�6C�I�|H(	��R�	ǲԺ�͎#[�*C�	�9l�d��+I�1$�hG��i��C䉬$�"01%�B�Ns
��� ��C�I.��p*��e��Q��]�ZZC�		���t��/*��R�AXi�<C�I�Fᮀ2"H����S��<l�
C�I"ܱ[�a��ǂsREW���B�	#�E[҇F�b��s"*bB�	�#�Lp�윤5^ ed�C�<B�	�Bp@y�(�~�耐CdOw��B�ɑ~;��R��9���T��B䉹B�)�C�{8��OL�j	�C�)� `H�R��E	����w��aG"OL!:L][ƩW>��i�""Ov�Ysj�P�ty������9�"O���$C�?Yl����P:8U��j�"O,�ZC�D�9DJK  ���� "O*��v�DQ�(0����m�ػ"OQ�b��jIfm���hM�̠6"OHY#�u��P�� Pi���"Ox�:B.>t���3o��ffPx;#"O��g��!����w�LU�A"O8t{�؃*�Pa���!09�U�F"O�( %�"B�$�1�H�3rA����"O�y�#��}����s��Z�R؋�"O�p�Cᚯ<jI�b��r^�x�"O�#���q�P�$�
�CY���"O��VCʃ{�IFK�UT�H�"O���q��*o]F��k[�&����B"O`ժ�$�J�
8yƌ��Z�V���"O�d�'ȳt u�dj[4]�P�"O.� C�A� C�!iuxuV��"Ox�ٜ	V|
�lݥPW~���"O ��Q�uXL!3�%S�n�
��"O`h��[�4V�A�@$�&O��m��"O|9�R�B(f?�E���Դr�u�g"O����-|\z�ņw]�Xʰ"O
�!��T`Њ�C�]U>h��"OBH��n6�B�!��R"NF��"Ot�c�
n\�����	
�@2�"O�y�F�5�n���
�I�F!Iv"O>�#a�^�Z����۝u/���"O�aض� 	V���a�W�[�f X�"O�03&K~8L�p��P3	δ�'"O���΅~g ��6lD76�(	c"O<�pq�ۻk��يu
^ 6ݦ���"O6����	-\Rj�D�ن/�*���"O2| a��iR���虷"@�z�"Oȹ�� F�?k�5�%���� �R"O����AÁ{�yj�Δb��=�b"O��� /��P�E��L
��XE"O�;�T$UC��rlB�x���"O��*��$w�ZGi	����"R"O2��C��S�`�8���"����"O����2*x��O�e
�Mh@"Oļ���g��Z�W�>�� �"OL�v�	9v|�	��c�;��hP"OƵ��b�o�L1#�(˦(Ȳ"OV�`�	�b�p�˃��� �l�p�"O>�#�O��粵���[�^�L$��"O"�a�)� �H`MF?l��q�"O:]��֯j��`��+ț7��)8�"Ob 0��*hbn�c0뗒��d8d"O��2ᄵ
�4E�3�yW�C%"Op��%/�]�� H�fH��
�"O��ԃ��~�{�D.5�}a�"O
=Q�f���֠�@-1 u��"O>��/TR��Q�D���p��"O�pA蚝+��I�f� �y��8�y��	(I f�ϫ(�݋�g&�y�hۦ6<�Y���Ǝ��y�cG��ybBJ9A�	:4DbdhP��l�y�*�Q������W�9�����y�ɋ4eD2d$�;;��0�`¦�y�\*+�d- 2�*�A�E%Ѕ�y��Y.U�͙���Id�q�p�R�y
� а[%"V�WK��bN�%��@�"O���&��X���F���NHR�(u"ONt� @(*J�仱�	�h\� �4"O�pf��,�ɘw�Һ)V
�s�"Ob�p����˜���� PD�	"Of��q����,���7XVVtC"O� �Y6
��[3O�!Blt"q"O:yCq���P�,��d|P�t�'"O����KB$ 
��"9I�h[�"Oԕ�`.�o�D����*!^�t��"OBDHDEۊ6�E#!-�/%ƅ1�"O�23�]=��a����
�>�7"O�%�e��1⠝
��c���""O.	��JA!.��l�v��7� ���"O���J�>�έ0��<x3���"O��#��ۣa�{E��.&��r�"O:���iڕ9������G����W"O��b�B�f(@t`T>hd�U"ON-k�&�K~�B�H��D�dh�"O`E��/à/�0��%���|���"O8Г��3 �9Q'���He�`"ODQA��&!p�� ��4��l �"O*��&�r.�-�Ɔ«�P�#"O��z��Fk4����V�8��"Ot�9'�ƯP�Yqc�մ$��	�"O�Q1�G�f��A �A �bm1V"O�تw��;)���h[�"[ B�"O�dXu�H  ��Q���:1yz�1�"O���(t9�Abg@��:n�H�"O"�JB9q)^̈�!��'���a�"O��7��)l���`D�X�s��a�"Oz�1�Ă�^֖M��#ʬQ���"O��C�%�8F�6�3L�23ӠEI�"OV���H�a0������21�"O�Ѐ�cQ�Q��1�DწT�z1�t"O�Y)� )�r,��O�s��ɀ�"O�C�JA$j��C�����"Oj-��*��fr�,�2N�y�*�"O�`��ݼ0�zXȕ�֐V����d"Od� >����Uz�t�b"O�5�t�G-3�҉K
��R��6"O����쓻?>�y��ܲ}l��J�"O��wj�VGP� /Z�A�n��"O�賡o]�f���;�o�s��E� "O:�j�-�s9�E���r��� "O�EJf(1
�AH���k��x�"Od _$����^,y��(�"O�)�$� 
p|HiR�E���'"O^��͙pZ,�9q坔h��� "O� �B1G��t�6f[�}P��""O�A�m^>Q�,cp�@?W�����"O��rS�Ĺ GD����Z��h�"O����EȸSW&e�f�5)�~�K�"O���W�݉[� �$���]�Ȱ�'"Od� �әy�L`m];.���"Oh��`��tI;1�b�Rĸ�"O�9�A����Zg)èO�xU�"O�!H�a
0?�\�G�/�F�c�"Ox�c�F��*R>�rG��<_�D�"ON9���J�3*��g,A�2�]��"O2��g�����p�E,=�S�"O�P�d�Llԑ�O8w�8|`F"O&u��G������ɷ���{�"O�Y ƙ�d��6�ˍx
�IP"D�� 4L�'Z�Y�+�E�df��3�"O���U�/}ZhY'S-5���"Ox-��/�*z֐qeܾ/� ��"O|@S&�e8�r�D�2UޤI��"O
����\�|���d�
jK�;�y�@�Y`l��DO��@�����y�X"twl����[� �8�Q�6�y��K�"�T(C"��� Z��a���y�ՌyĖYG�W;�� ����yr�D���$�N��mN�ln!�O%���r� �Y���b��Z!�D�m��R��ۢh��=:�lT!�$�q5��G��Rr`����GW!�DA�J$Q#P�D�!8zU�$,ЖK�!�"[���WG�(N]��*J|�!�dԂOʔ��<o���C2�!�d�:]�ۢ�k6���I %!��I
����M �|�p���eޒ�!�DN]&t�ңŮBh���DM�M�!��*t�Ԭ���D�!]r ����!�D޺%q(\���I�",&��Q�M/�!��U��T1��C�%+�� �C�\�!�D�e%t̓-��f����%'^�z�!�Dܺw|�D�͂?$� @'�&�!�d��А�����f��40��A�R&!�$ιe����U�H��Z�5�4!�$Q$2�t�����<+N��$牙>�!��1=�j�9�i�!=�%:P��m�!��E�T�<I
"�A3k�ʄ*��Q+(�!���d���Ι�TbB�>!�!��H�M��JOՐ��C���s�!��*Z*�Q�q��;�<�3b.W��!�#�|�����wC2)�m��*�!��+$c�Q�VD��d!ؓa��	2�!�dВME�	��k(�zw��3B!�d�i��(�#��,�|�LƬn�!�\�{�$d����MW�Ђ�J[
Z�!��̕!6��I�C��d""9���Z��!���;���IP�ș�T*�-!�$�4�½��B�#.g���κg!�D�.q�({#o�Sr�q�"g�P,!򄕁>�NI�G&� �z�{!��N�yL���$Vl���f�!����A�0i�:!���!N;�!�d�
Kf�Ū�S d��Q&A��s�!��.� q0��)���9$���!�D�9q��CB�ȉ)��M��n� G�!�$ٓ|���E�>���hu�G�x�!�D�>"0����'�/��%R'C��Ze!��Ȉ���2R]f�j���9T�!�$S�c�<z�R�
<4`�Aa��W�!�Đg,�u�'=Sۜ�����3y!!��*:�"]�ClH4�py{��e�!�dX Db7�H��5�"��8u,!�$�_�B�Y?pƂl+�ɍ,!�d�&3�A��Z/a�X�w�Ͱ.�!�KG�]�V@� 2M���y�!�䋓k�ZG�Ҵj�qH4W�!�D�Lp�`�����(��*|�!�$R�]�>q�����vY�Q���
�HQ�{��4SZ���aO�IB�NIvE!��Gp;��1���?aљ �! +!��['��$'^�u_\����%�!�DUv���D��0]XV��L��!�� �'
� a&r01��f�R%�s"OX ktM�&^ˮ��S��1��ŉ"OVh0��D9n���򕮞�XE�"O 5��)�27��y����Q~����'R�Լrb\�獇�>��قd��!�dߴ�tlZ���,^1�7$��L!򄇗t��:�F6\��=�w#��1��}ґ��;J�%B�c��S�A4���)<D���ҋR���IU��4(��,>D�����C�[�� �ܥXS����?�����R�9��B�	���:�l��Dh����'#��X�?���R��8�mrb*hs!�䚀���
q�XD�6`���8l!�$!J�r|�� Ά�� ᄄr!���+C�܌DM]�<��a#��� Y!��֞fPpa �,G��t�ǈ)~M!�DY���xs�Ҏ@���3���*,K!�$�y���@R�0� ���
8!�ɨ^p$�@��X�z�0�ڃ�Č\'!�d�����P�j��;gQ�'!��A��IZCjU($��6#�9w�!�L�#(�l�ş�U���@sG�����
0^J�a�!-��
*�yhR��;@���5=z��p��Y?�f�I��+� �ȓo���a�/�2<Ig�Őg�U�ȓ@�d�I�m�_��� �@:$��ȓ���R��N���[T'J%����ȓm�`V�7����K���\+�"O�8�Eإ�R$�6c� :箽���Iy�'��D1��3Nˍj�� 3p�	O���g�'�b���۴���|YF,H��g�"���4D��+��E5�)s&&�+K�
���a4D�#5BGD� t)'�#7#p���0D�Թê�!�2���D�6�����/D�L��[&0m|l�a˗�o�����.|O�c�p����5	�2\y6nR�h%��D,D���eA	�B#H$+��Q�e�zm8��?D���$�; ��E��+P$���Y$�=|O�c���dN�98��ܰ��BU@��3v�;D�ؑ�o�R	9�&ߟYGre{D�9D���[�Y�xUlϤ$H>��%8D��5��F,0q(�*B���#+D�3��	�|Q�����]*pM,D��8�	l @t�F�	�H���"�+D�Ћ�H�6?��UX��\�)��(�n3<OH#<����IA�H鐤I"�.�
�Zb�<1�@U �����M�S����G�]�<���W:l�@Q�lY�6� E�ǋ^~�<Y�cBD�:��쇼1��Dr�Ο_�<�U�֋@��Aa��O�d"�i"+�ݟ��P����'_�� O�z��\���M4n�!򤔥&��H�P�Fz��0v�/4x��)�'j�b	��$H*	��u��������x�,�"-�z��Д?�(��#߯�yb�U�PA�d(�
ƣFZP-Q#U�<�@��Z���h����fܬaJO�<��F ���d��M� *�l�4K�ry��'�ֹ��n�3	s�@��&e̹���OD��ԁ �����'$>�A�Q�$'�,��	�kX�̊`���l�K �d��0?� j�#e��ы2疉	��z&��<�T�"(�z�h`�ĎIN��iq��z�<ɣ�"O�PŐA,^��\�@��R�<�@��%�C�хJ�� 0A�Ly��'1B�|��� ��*�F��2�W�J�Z4H`�"OL�зB�8�b ���K�@���R���'az���H1ǆ�aϬ9���ّ�y���6���x���+aՔ���h 3�yr �p��l���	l� (���y�N�=!����fK�(��,���yB�E�7Z�U)M�.4f��u�Z���D�Ot�0��?�'}�����cU�M�#��:�z	�'��Ey3L��2�q*G���y��{���hO?��s�3d��G��0T����<����L�.��F�"AV�+�k�c�<!�@͊|E�8!O �%����V�QE�<�4���u��\C6�[*f�� v&l�<�6I��0,���"-�~�p3
_g���hO�'}7��#��V�9Y~��"�e���T]^�أ�^�Ha�8�Mɇo���F�3V�"Í?���ɓ���Q� B�	55��"#
Y�����c_v\�C�	�26�h���A�Ps�! !�B�ɼ
d�����v����!̘)"�B�I�?�1K�ẺW�˒k��x�O���D:Y��qua��n9��@�N�)�!򄇼p'���f��hy��"��P�!�Չv���$�oJn�P/��!�ūmX�s�=/��� �+>t!�dޖBYN0pթ6|@�+���/ku!�d�7	����ᓚa�4YSMԡVh!�d܆}�����@>���[��vf!�L�)�0����dLR]:�
��6X�'sa|2i�Q����*�4cnV�d���������4Z#�}ab1�6��7��}2�"O���O�l��7�0G�><Q�"O�mA�,�qi.U�0�M�
ԑ�C"ORy#"MŻV# 8�r ]�i�N)+�"O*�S#b� ���nG 9��l��"O0��f�l	���عJV�}�Z�Ԇ�I!j��IsƋ���l5���hj�O`�=�}�a`_�&�j(�ƍI(]�$���bx���'�L��vM��~��	M�`#	�'6 T1c_�y��)�dC�,=��9�'��M��ޗ&�r�ɏ�<�Hq��'|�e���,o"�A�M��/਩ȍ��8�����B�M�4�	�,A�Lڇ��|>��$�z�h��׻[b]1q�8�O��I��0ٻ����X �ϩt
�C�I�x�L��7 (&=&U���?BbC�Ɏ_����N#4�Qg3\6C�	y40T1�fۼm�y��ئXlB�I%8�U���I���3g陌|�\B�I�V���f�.t��`Tk֢
b��?���	ضX��yA�8R�Kt��M��'��O2˧���ۚ5�*t�Cҋc~8"����!�؀w����'mI�������!�躥��G7�([Q!I5!���n��	�2 0�Ơ�@	 !�d�RB
�4Iߕ�<����!�$H�m� ���G�Mk�B�]1I!����~�A�◤}>)&K]�!�$Εex�[U� �c��負ɯJx!�!L4�3��e�zyJD �/-Z!�dG�O+^�[F��)&�pڥ/��I!�d�m��5`d&�H��BA�Ŀ-8!���Tpȼ[����[���.k��Ο<��K�޵�1F��L��P��"~�4B�)� ~����]V&���A��`�(�9�"O�1�oH�D2D) ��Y�e
G"O�T�) ,|���M&�N$"A"O�	T�G�E����n��xv )A "Od%r�-ʫ=��c�){]R���O�p�ݝ&(�YU�I5y���	�,D�J�GI��C�Ŋ$��aB)D�|1g�4���;Eo@�d��MZ�.)D��X�͒�[���P3���H����&D��Q&,U�pNhM���&=2��D$D�d�w̟�$���F�J6U�N�i� D���F-��f�@��:Y�B�=D����O�nQ��Afk�8}ךx�t�6D��c�'C�6�Q��&}�<X�"8D�L�LD2O���Hu���>nJ�wC+D�8�%�M�W�
AX�A�$l�&����=D����EǔX�����*(�����=D�<#�	���I�/!ot-p*<D�d�5�&��L���2�8��d.D�p��/}��X���Tk�-Ad!.��0|�靛N�`�J��Ƴj��E[	�V�<�BǏ(CL��$U%]QX���d�y�<1��j��)j
E�9��8��lt�'t?A�Pb΂O
��� C�H����-9D�`� ]�i��)R'f��x��g6D�\�p���o��E�7cU�2KD�y7A?D��Y���.�^y��eR�7I05a;D����- Y�@����^��0qU�:D��
,J�v�A�_r�K%�,D��C7�� X�!��&]<[�����,��Z��P2q�4>1�ijV3�`uQu�>D����ɿYw$���j�LY;�7D�X�⅐="�A*�46,r�5(D���G�M���1�ʋ��Z�ZPg$D��ASARI]H<�!�D�VD�Ї� D�.�o�֡��6������ D� KS"[�q�xq�F4	��5R�I)��*�O6�J�iW;9C���B�O�-��\æ"O���I��3�N�1{�R�˱"O�XA�͈i��q�����z�"OD���kCn��@a	��e_B�R�"O�5(�(ݱG*���DI�<_@��آ"O���w�A�� 9���(H �"O�t'`�AM��A�=(d�v^����j������P	�l��U�m����:$�S%D�p+�O�"��s񏛠x�D9��)D���t�N�z���$mף7�&����%D�T�w�H(m�D�Z�c�� Tm>D��A���?W�Fy[�-ԏj[�H��;D���%��?�j����M�P!v�;��X�'��d�RE��!�*�Q^1��
Z�^��'la|B'�C�p;���/����(��yo�5:Ń�����P	Bf��y���0����4K 9����刅��y�*��w�6��u�M��@00Uj�!�yRa�P �Y�G̔�y���s�>�yr�2������t�\��s'U��y���)O3i�d��u��F���D�O�����bę���%}�}�so��e!�$��\�yRF�:f��q���o`!�dY�/�r���)��^����#�!gY!�Ā�pђ��bE
?��L��AY�p@!� �<`��y0-۞+��|k'c/h!�$��\R>���R�3�p�c�j�!�� �1�ѭ���)��#�>���s"Otʅ �T��iAY�v��#"O@����)x�2�a��詒�"ODX�0ǌn�h ��NF�
���Y�"O깢�$�$G�Ĝ�W���JFTI�d"OZl��FL�{v�@D� �39���"O ��¤Y?��_�@P+��:�!�D�SU@�Aăc���*㡑"��d2�O� ���+>^"y�*�@{�E��"Op��
�W�5 �)�i<�Q"O��e��6dt&��5�ŗ&2Z�"O�J��D2@X����;^�)x"Opak CX9E�bu[3�ղ-�BhA�"O�Ei�&���48`L�&8ҁ�"O�I�Sʆ9*Y��5LP;"�.$+�T���Im��B�!oj��	q�U�r�
m���$D��`D�U�EL�k��f9J�&D��
� \1v��2CXU��iH/D��c`ڀ08I!1�Zp(�!hW�7D����O�(�L�V	+zk|!1�a4D�Шᨎ)P&�4jvk��uZt�a�1D����z����4�_z���l1D�Ա�F>ppL��*ݚr��X��1D��e�ޡF]h�у��?[ � G,D�8�c��w���QK�e�ܡY�F,D�`�d�1�N��w�+A���a$*D��9d�H�?�X��I�d)� ѣ-=D��8��D�U��j��L��ؠD')D�4�`�E�M��;�!�+�X�G�'D�l���C6��a���o�d��%D�`R-N%zl�j���`Фc�.$D����l]�w="�M�	=�8��*!D����L8jO�5@��	-��<��/ D���`�����]p J*'
L��>��H���S�q�4#��:ds
H��� u��$��1+RU��(8 �$�ɱN��!�h���� �"�HԑGKP��!�͸0ʆx�ϯ4��H���^�g!��i� ����\�Lī��_	!�D��4��۷�\�SRГA��(]!���Q�m��`�RXh��N�P!�d]�/�àb�6]M0�
���[!�d!B�]�S���{�B�bS�=E�{���g&����@1��b	3g�!�$�]����	3)��#��w�!��8O6]��:oZ1�[�L�!��L�����hA�YqM�!E�X�Ik��(�p1��������ɕ<�H�"O��8��؉�t=�4�@�2���2s�d>LO$ё�A�t���r#��5H傕�'B� ٲm?^�`0B��6<�Bqg4D����߈c ���*K���J҈3D� �f�V�*1��KÞM��CC�.D�X��j�-f�{RgB�o06��B�<����.@�!ak�㺨Z ��zP�C��8g�-�Ee
ɮ�H7X,:9�B�	R2 y�\�{p����<Z�?����D6'�zY���P�7�X�ZT�%n!���Pln�+D�(�ɱ�Y4b!�dA�&SH@��S�Ŋ"�Jτ!I!�4<e��bb�r���EJ��@+!򄒝IbfD����6�,a���n!�$� ����p �-��u�U"�6u!�dY"h'��(�m�${�9!�Ѕ!�� &�A�kN�LZ^�*g�@�f���"O��+A!����qA�	885FL�"O�=Z+UY�԰��F�-H�P�"OD�cL�<9\�
Uπ�u����"O"���B\! ���u���)!"O2����)-R1��ė �m��"OUh0��\MH���Ǖ�:���"O�l*Lʹ|�$�;#�Q�l�*�*O��H�.��&�@$��f���'�@QZ%�S�/A�:�ƚa�Pa��']��Xd�=R��S�Y 1|�	�'YN�j�	��p�Bs�!4;�� 	�'2z���,� :�{��xa�ȓT�E��Ǐ`7&���ဏy�P��'Lb���H��;VJ[9@{�!��D�e(vB�c�L=#7A�	c��AL�|B䉺Z���1�Ȯ!�B�"v`��8��C�	�����%%	G���$,߀��C䉗����
*b�D���=~�~C�	�S��4!n	
)�P��i�8IXC�	$[�mS�� "W���nF�TC�_�ī�!3z�n����[)BC�ɴC�@��@�W�0H2�AB�
(�C䉦T����v@�A�&41��A
I�B�I�+��2!�7J��م�Z��B�I�A\Ir�n��F0��A'%?�C�{�\8'�0&5�0�#�+��C�	�� <xr�
h��DɳZ�b�|C�	
J�8)�ui�/8,���E�'4ضC�	�FP	{d��[jPH3�C�C�I�'K����ͨ�"�iF�߁}�RC�	�(��<B $�n���`�
�$p!�dS��<�:�J� k����A/.!�DS&z��˧G�/,�hd��^!�dC	di�"��JZ��ه$�>D�!����@Zc���eNV�`de�!���se�a�peZ'>/N�[F����!򤒒y�>) �坡G�~������!�68������E���K���'�!��9
��L�0+�n}1�a�d!�[.q�<����Ba�`BF���#l��)�8q��� ��"�`�a�k�,�J�'H
*V8Z��lj��	�+�&�P
�'���aLɖ*MPp�W�*	�ݣ	�'���@�Y�9k���%�� �'���d�Gs<ֽI�@<.Ѐu��'8�;�X<'�N��4MD>[�t�A�'�D���'*t0q���ě*�ܨ��'�~U3�H�-b�!��ȸ�E�	�'�:�K�X_,bDŖ3��	�'s��'IQ�&�ā�Ta\�D����'�X�k��;V2�rA�2C�`[�'��e��d֫�<!��OHBi��'-���i0q�* �b��:)� y
�'�<��� �̙�����5�� 2
�'����pb��_(eb�c��!�'3��0���R ȫ�F@���	�'BL��g.K�"\2���!{�8d�	�'��z�cY�D�.�;�)l�`��'���r��!9X�\��K]7_n�*�'a����I�����h�%\ST�z�'�dI{����'��'��I$����B$KI"�@��	
BC�	�O��S��%~�"�E醍	�6C�I�& �Yt�ÍIb��>o�C�)� �\�G��; XaꓥH�wD��1"O�t��(�G�~��E.gJ)f"O�(�����
�V=#�C��3_v-yY����	/�x��F+Y;x6 ���N�s��B�+$Ք��� �8� ���(B�ɍ?z���ϖ�AuN�W!K)4sB�b�>��e��{h2��6'��7��C�ɻC�������1Sℙ7�lC䉻U$J�׎ֈH �݀��X~tB�ɞIZ��Dm$�$��b�����C�I�W�*Ȧn�((�Rt�I�o�.C�^���B�%ؓ
)�8�r�C5Rg�B�ɐw��a���2�tA�uh��|��B�I��(�L.}g\y�D�ݜ�B�	,����%�Z�<1X�D]�.F�B�I�G|�"�'JK��W�"lw����|��{�Ų@����iJ0R�}�CN+D�H�թV������w$lh2a'D��j�I�d�=���7]R4��<Q����k���C
�.W�����B�Xi�B�ɾz�P���H�y�X�0ŀ9^�C�I�KL�*��Ӛh,�t�0���xvjC��?>�و/kz�g�3}LC�	� ��j3��;��|����-#�|!�ȓzP� !��p�^�c�OӪk�j)�����CԾx��D���c�2��ȓt� A� Y4B_�e �@�VB剶2�Z���� 3�[$�\��B�	�����wL)M��y!��[�˘B�	�1��1��O �E�E)�s������O��!B�S�Y RܠD�L�c*ֈ��o'D���ԣw��Р
^9���S��&D�������+H��⎯`ʐ!Q
?D���@�1q��2g�D�R��`	?D� ���k�`��j�D�8�7D�4��#T�Yi�QCZ�L;4D�`�$m&���.خ=P��@��2D���&fT�vh���g�[;N8nDh�>D��sO\��&���bEoΰ�8p�ۅO6�O��)�3}"�|��`�0�D��E�r��y�-�>�\U��w; �i����y�63�(G,\�"�b�����y	R =8��ʙK��Y��IͲ�y�G~�Tt�5*]VH�J�.3�y��W�E���
Cdʩǐ���e���y�/�t�l؀B�À��I G H2���j�Hi��"��S� `*��E�G�&�R�DZ�B�	
1��8#4�V;&8�GE�
����?	���)�n5��ѓh�=J�D!:$�=�!�
�I�*!Y��C��Xa#7���r�!�$7r�d����+�&�b��94���;OļyD��
�
X��ܕc��!"O6�� �ŹV�B�"�
Q��d������O���)ˍ,���k]<z�XL8F���-�!� 
;v9���M�~:@ep�a��{�!�-�~����&_4��䠈,C\!�DP=}�<Pe�
�Π8�/��!�S�?�<����R�E�4	拌�jޡ�d�jlpPhФ_�U�-A�fT-8�B��7z�\Ke�t����@iS��O�K�F-��f�'s���C0�[��0�Br�E�#��ȓ
Gt�e���x\��g� A�"4$��D{��D���.������$P���/�y��X	!v�`��(<�-
f�]��y
� ����+Χ#�x���O�`�s�'G��!8�*��d��0D���c�Rr!�$G�v�VEȄ���q�,�z��Ƴ!�ў0�ᓔjP���g��)x:8��+ŐC��B�	�Ht��2��ť3�൨��A���B�	�w<�	��5A4�E�E�>��B��
m0�!����YFb��t��~�B�	-�V�b&):@���2��ΎMP��$&�	 L:P�z%�@a&i)s��I�ن�]���R�-`O�G�Z�n�HB�ɖ���j�Ȇ�[����a����C�I5�b�����u��a!hE+KF�B�I9d�
$��(�r�BD��or�C�	�:���B��d����j |?NC�I .3(<Pe�_��}��H�'y	�?�*O�c>a�
�&��]3���gJZ�p��8D��SRF9��%q����P�XQH �:D����d���[��x� `&��������T16�vy�A(�=sZ����"O̭�A-�/:�Lxd��v�֟x1!�ČQtp���Wb��l1!�d�b��YĮ��aU�r�N;/0�y��	i�2��Q,�nI�x�#�:IBB��<b��!	��ʔ�Bl�9��C��M�H���  G�� x%��~2�C�ɴn�D�E�� 
!b̪��*$lC䉧p����"jV�(^B�B'K~tC�Ʌ1T}2u�"<Fz�3wg�P'�B�I�ƌ{f�490��F� {tB�I�{�B�J���;v�ipEJ��$C�	�#$X4H�}�tU1���ftC�	3h�j�i��2pE�͆.A��B�	(w�����(xb���ǘ3�B�	1���D�=%͂�qK�%lF�B��5E�v���I�<"H�d�E�DB䉽��4��%��r6�؃
,B�	848K�	`�c7�X�I�B�I�Sr�B�b^�k�Yb�j[�B��	`���Ӂ�[�+�,�Q5G��B�I�b��1f�J�&��c� ���B�ɩ�4��`�:f&�0�NY�КC�I�m.Y
��Z � P@��+�|C�I�7�dp�B�N�bլ�k��9�HC�I�l5��e�/��ґ�^�e���O�=�}��ƈts>mZ���`|\p���f�<yӆ&���Z�FX�C	�)��RX�<I&�^a�a�B�C�.��eWW�<A1J	�mX&�d7:Հ�R7�H�<!�ΐ�C�H���F�O��$��^�<	ӫ�-,Ab���S�w��*B[�<�c�[4*@���GbG?��Z���@y��)�';���p@��Po��%!� �T<��T�pH�v�0f���r�� ����OgN����R�A5P�R�G�R°���$�T,�aI��:�(�b�Dq��$��-�k �7�Ԩ1��D�J%�ȓL�C&l�1	��%c�G��%ؤŅȓ
�8g	IC����7A�>8z�L�IX����L� ��R*7
ʑ�&K�QV�u�q-D����#��,L9GfI�>ː���,D�0!7(Mtڈ$x�.¾8�\�à*D��7	.Y, �'D�9c�9��2D�x�
{Z�T� �O{-�q��<D�x����9� �����?g��H-D�� :=� # '3�:HB1*[�o�����'/џ�'��͓P�Ny�	�W�
�s	�YJ\���p%\���E�	���LP\�nЇȓ?��ҡ�0������Ș38]�ȓz(�@&��������^���T�J��䓥IA��C��T�v�J�ȓg{H х��].Bl���I�>N�!�ȓk!t���M���p��H�!Wd�Ĕ'a~b�A){<R�˄B�E_n�	E(?�y� ށN��8qf՝B���a���y��W�p���ط(�6^�,��y"���yS�İ�掜C��K��D	�y���p� qf,��-�h� ����yr�HE^UD�ګ\Tf	���]�<�b�*�ĂP��pa2��v�<ip��J`���I'%H��lAv�<�cf�*����7���`��$�u�<��"E^*&jӒm���I�F�<�dب�j�$�0�Y!5D�I�<�Ç(e�� ��F�
�|�����<��e@�-[^�)C��K�q���ph<���N�]�>�{C��&q��� "ި�y��R�x@��S7&�9e�"��c ��yB-�\l����ÙI�^`�ċ���y�dĀ=	q��G����U'�y�T�wެ���EѦFG�9	�"ö�yb`F�^,HAe�ܤ:8� ����y2eR�b���b�/J�5�X���gN��y⭕� 	H��\4-%YkbK��y� ��\�RYh�C�q���QU�X�y)7���Q�ʇ�o�$��DN��y�O�"���4GK&�4dhd���y����&I�Po <�<����݋�y��U<1R�ypU�	�+�X�e�'�y"���B5!�׆�!�Â��y��ފ|��3���'o��;����yR������H'z�Z��ٙ�yL��D ��Œ	���ñ�C��yRHU4$���8K@hA�g�4�y�I,t�a�bߵ\o��@�N��y�.�i��;Gc�B��� ��y2k�.W8qU�C�/8Z�
�b���y�- ���*��ي.��l�����yrƘ!o��5�Վ܀t'�9*�d��yre� ���`CB*h�"���yb6��$��ǯ__��{De�7�ym�*m�.���ǸJ�>�[䮛�y�K>Yּ�Hr�C&=D��ϗ�y򦁏v�RL�ѣ� 4n�9`\|�Մ�rB� �WˮA	���	K"
�F�ȓF��Z0H��zd̓7�"Hj��ȓ|����"�ʾv�|�%H>���s�n;d�.T+d��/�+Aڰ����<Iʷr���@bϤ]�@��U����tI@�~�h�գ��>��]���v����\�F{@H�g�y]�ȓh;h݉V�İ$ ��yCGyLL��:c���rG�DK�D��H��5�����p-�nϙ8nAR��;���j"�����I�>��̸0h	RX�Y�ȓp>N�H�
 ��`�'�}���ȓ��W�Ґfh<�$�U5�,T�ȓ��u��BE2g1�����
1 ��ȓ�����;zI���ACܗ>�Յ�S�? �X��I'Jf��6[�r\Z�� "O` T�V1i�~x��A�$\����"O�����A0[�jA[�AK�T-�D"Oz��	B ��$�F�4t�����"O��7�M�l�r��s�ˈ�fLj�"O�D;��8�©�G�ճ]�� �"O�`z��;A,�Db���>�jV"OD=�1�M�#T�Պ�b֏t��IY�"O������7�ێkH���"OL\�&��'�|������"O`J�����H� ��]+7"���"O2 uE�?$�ĺ�M�^	"�j1"O8�����6tԊ��t��2^&�0R"O���N�cR��;qLφ>q��(�"O2hb� �3lf"��An$sk�A�"O�	�1׻f���'ݛ���ف"O�Ѣ�#;��2��{P*��!"O�9�Q�r��j�ݜq�条�"O�i bb��F�Q�B���0�F"O2���,Y<H����fR�^��xp�"O�؁bmŻX@4+�E����b�"O�M��A����2׊E�YgP�Ca"O��b	͵�����hE�d�0�e"O4,�gF�4��d'yS2 �"OZ��4�N�`ͬ�J%$�TJ�hhg"O4�ti�
*~D�A��B*��	�"O�T1Γc�ܸ���P�l $ŉ�"Orِ�gԯGl�t�Z'%Y�t2�"Ov-qO�S�����ٌ|J���"Ot�z��#L�a�*?NJ�(""O:��
�mF�-y�J�D����"O���e��:� ���\�n� Hs"Ox@�c���x`13�Q�:�Vl�"Ot������{b�x����r� Uˤ"Ob��֡�$@(�f��
j�j�˕"O4������ԕ�¢��	�>J"O��BE_����b��!�d��"OL�ď�ONeq'ѪP���#w"OLqQ'ҍ q�6�� �Flۅ"Oe�c�5���T���	w6h�s"O�UY�Z�'��y	7k�2FJ�e�3"O�Ӥ��m�Z���̞�64�w"O�����O���j�+T�"��B�"Or�{�c=zrʌ��J֨Yȴڰ"OޭA� �HE��8t'��E�B"O@H���4P@~������q��,If"O����CTJI�%I�G��\��"O�}('��U�$�V地^��x;�"OP8I,��b~$�C�,����r"O~ms �X��!��Ս{�A�"OnA�VLˌtR	�^�B��n��y��"h��q�'��<����y�(��@�����T�+��x�w��>�y$�f�HEQ'D�W������y2�j�3���{�椨G/��y��n@�y�.�o4Np����y��M;'�<�3懆n�����f ��yb��bY��C@M�;ͺ���Ⱥ�yB������J"��0������/�y2a@%Ƶ�`E��*�ԉC�/���y�o�-,Q�!�r%�&���x.¨�y�/��\�� 3Lء�����yb�[��W$�:'��Y"��˃�y�L�	H����pf�%Ȕp%�5�y
�  d�pN�"����C�f�FL� "OL���P�=��"��">!�b"O♙��$y�@�+B�I �d�8t"O�x��4/p�"H��5Ȭ���"O@	8�F�F��󴉜�X�%��"Oȅ�U��
���s�ܬ�:l�"O0�Y��'WK���`��7��h�F"O�]��� �ܠ$�z���S"O�(І��Dc��%���Q*�"O���ǈ�&{%�x���׏����"O�u@�ܛ'�D�emo�	�"O@��.!`^�B�K��:�>q�G"O��Ԃ�c�웄����p�"O���7�V�B��Z���
��}�"O8�l��d�҉��HT!	�$��"O�ըS������5J��>��"O��#o�6[HT�HA�Ы�Ȁ��"O���.���Z���Boj,DS"O��ҳ(� W��*�_���\�"O̱��P�80�U���M�AK���t"O�I�u!*Ӿ�Wm�K����"O�hї!|M�0�3�X����"O�sf`$~r٠&I&M����"O��S�C�����$�'M��-I�"O~��#��Xm���b�P�c��0�4"OΠ{׍K�:�1z��^��98�"O��2S
�#J�)�dY��\��"O�x�1&Þ_Q�x�%[7	���"O`��煣	����
;s(�9�"O��jD����ܪ��k]�p�"O�}��.\�k/x,8҈�#Bk���"O@�a�o��^���mD�j�lzG"O��B�ɏ-Q�ը���#Jϴ���"O0���Gڻ%��Yd
�+>�����"O�-��̅e�k��K�o�YP"O�uk $ޅ{������4�Ҵ��"O�rq���%3V�����$}��v"O�������Q�EfWk<<Ca"O���k݁UD����#Td��E"On ��Є�� �ɔ�LEXQ�6"Oda'��%ؼ�i��:&��$"O"���.Vp�h�cP���H 6"O~dB�lL*�]`�4�4P��"O���T��r���!m�D��m�%"ON=��"ܴ]$�C��*���"OHH�V�Y�T����T��Sn4���"O�0"`�ϛ!v�iĆ���=�"O�����5�0�[�儸>�l9�"O����͠I��u�	�M�̨�p"O��&��M�B��$$,y"�	E"OT���(^.�-����-\I�U"O�	I�� Fj��3��m8��T"O�s�EU�+~ơYg`Іf���"O��DG��G/vAӷn� >!�Qc	�'Xl��@�={�(p*@;�H�X�'yd�y��	.�kV�F�t�E�
�'��`��o�<����m�8U�
�q�'�������$��c�O�F[z�I�'�h06�!M�x¤(�iB=�'�F�HC��yת��"me!���y�/�L6�a ��2g�y�7Ù=�yB QY����+.F�4&	@��y"Ο0/�έԇ.@�[EB�&�y"�SȊ`��mf�}�DG�flB�)� 4u�ԡ�-�4��%Sf����"O����4B�%ꠃY2F���P�"O��x5(ѐ?��̙�A�6i�,�"O4$�cW@8��ᎀ0�
D�"O�9�5��&�8��V��a�T@3"Oޱ*���cB��OS�~�D��"O��"�`[�\2v|���K3�|��"O�iP �L.+=�A+�倴l�&�Z"OrA�q� 2�6=b�ĕ'c��24"Oı;u�\+��e�r!����"Oz=bP�
�"����Х.���Z "Oތ'F�7�M!J�t#�"O�m�g�j���ʷI	9|J�"O2i٠K�QJ�I1� �&FlpP"O
���Q>W6J���o�r,-�T"ON�⇪	�rA����:vx$Z"O�2PJ�_1�aY�˖4���2"O&��ㄇ���ᔠ�� �(A3�"O ���@�d��K���2�Lj�"O����Jҭ2��z!�_�{�"O��{ƶ�v�3�GJ�BqrS"O~����ܾYV��c�(׫9PH�h"ORx�����a����/F���y��#O頉R� ֘o1(�9����y�ߓH��X��'L�g��0�eº�y��Fy���Y�ڥj���+��ү�y�J%7$D���L� n���`�D��y2��:vD)��7����a�M��y�`6f'�]�CÐ5_�h4���yr��S������r ch��y�Ú����c	�PH�07���'�ў�O^���l�)-ubD���s��K�{�'��s3�	�M� ��@�rL��#�'�l#b�B�E��UZ�kܩ���'�dd
���)��`��DO*T�M����?�'M*Y�g��?{qZ����On��d��IE�%�
�Z2L�5�ʭ��܋l�|�	��?��}��)ԉ4���2��N4v��9�U�Ö	��C�!G�AC��p��ep��- �˓��'ў�S�QtT��e�2g����f����df��x�$���jf�!�T�9��!�n�����'�ў�U�7V<0�B�ҥz�t=��9���~O�����q���*�.��Fs�(�Ƨyqܘ��k���K��5n�<��X�i���O �=���*�9k` q���&p��]�<a��I�c��+N4 $�u ��'azrO@3l/l��5��-ո]`�H�0=��" ղx�`���	.��1�ۖ�y��� IS�Ac
�;�H��]���'Rў�OȚ���K�@��a�Ƭ�(|"�(��'�(�#fFD6$"\��@�l��R���3Ox�iw+�"}��p
"K5��J�"O���2�� ��c�f�J�X1�q"OT��4�	O�f�{�%ؾda1A�"O�-��l j�U�֍ �EnA�#"O�hc�1Tn����*�[�P��'����F�@qvh�/���C�gt�dB�	�TU��H�ꊄk��̿<,O��=�~2 ��G�p�5�(e� <���4T���thCb眅������#@֦���}}��O�3ʓ}������*+�����Kב��h�ȓxXY B�b�Ii� Ϣ$�$�(��I�L�v��fn��4Jق��yYB䉍e����D��\c̓�~I��"O� ������t�!3�`��w�,hi��I_�����:b][D��9'[]��G�>;h�y"�	�&:�Aå�X=�h���BrfC�I�C�@��w�5`��|�LL��B�	�l���x�@���
F	�M�ȓI�����p�4��E��(���-|��F�ǯwfDax3kD1�v<�ȓjT����d�(x%�A��\�"%�ȓn1N�a���(t���+ �� �ȓ]�x����z�{U�D9��N���fm���H��dbR��ȓC<,24�.j�h���;1�ȓaL��"X��\��B��U�	��tU֥rRIT��$��aH7`��=�O���Dۈ)�`�SU�@�(�8��7BR($ar�O�m�#�R�-�V]23�O��;*O�ݻւ�"{����� �7S�AQ�'H�If�$4�*W��i�CA0#h��6M�E��M���ZŠ�f-t�6eH��V�Y��Q�',�{��)���L�d��x��'q�<8��=���'q�'x����!�%�ظ�5���kb:��5\����I���h�V�Q6�eѡ���3���D?ړa۠hq�#iF����am����VuV����B�"Q< �F����f��?	
ӓ8�i���L����K%����)�\���;az]�&@A�����J�I�#R ;��`c���ReDy�)Y>ɀ�Z�#��{  �s*��X7�+D�T�v�E&\3�Xd� [���V"K��hO?���]:"d��E?$��q�F	�HA!��K�a|��P2�d�r��A��y&S�'�ў��W�̝o�M"��q�*��&�O���'����E[6�*��@C��mj	�'������͚)���
�t`���F;�S�	O�B��|h�f�S��z`��57!��C���5��	��Ȣ���v(���ا��r 7J�<�Y���(iK�4(V.��0?�+O��°U
z�92�Ҽ-�PH;��'��O��	D�S��<\@D��m܇K(�#�K�'c�^">ь���<$(�[�
�\a��
�@N���>����Z��J�×?o���DC�<i�-I�g���3Gj���L��F�@��3�O���uAQ�uiڤ��ȉ#N���"O&��qG�;��y(�&���4��'Q��#>�4 C��W��!��ۗA��C�48��]�E�M sj�!b�̅(�B�I.'�"mA�Μw��aٷ�I�)L�C�o�}87H+�P��c�% J�C�	�gy����	�0RD�r�H�W��C�I<e����c�1R5 2�@�}/��S����O�	R%�Ɖ
�����,���'VQ�,� �җ�hD{�Χi-|)QV�3�I=%�2"<���y#C">MB��ɷ�W9t�N-3�"O��rRF�@7�$�#%��s��8�����OB�}��I?tɻ�����m[�'$)�؇ȓVNdq4
4A8���hK"M-P���B<aՋђ�&m�$��%�D�YD� S���'�����ڠG�@�*�
̎0���(�'j�� ��  $��ݣ!�&1��죎�d#��T����?q,�Q˃��U�ȓ(X���An�����%�5j-���A�f+G���DH�82H�M�X���M�/z1���g��p�%R�j��O�,�-;ޭmB�|�.5pW'9D�� ��"�M�@�q�J,5 Y:��' 9�'F
H���I(N+4�z��3i�u8H>���I���p4x"߽cL<	'��J�Q��O�b>�7�V���`��L)��ERS�1��u���K��ڢ,[�����r�H-�S`0�O|�'�(�����n��ܢ��,��q)W"O��0���,R(	٤�ؓ;�t`w�r���'U��,"?�K��O(5TmU!h0�C��L��?�t� 9m�\�2ԇG�9:L�%�Ѧ��'���3���$������
���+���d�B�ɰ=i�9�Ǖ>g�T����Y�/n���]Z����t�m��@!	O!w}d��e`֟�D{���͏l:\��	�%@0y��/�B�	�s*�x6M!6-ܒ�?_��B�ɬTɊ��a��(�xғ���B=f�?��)T�j�����S�G���JWY�!��@
o6l�3�(^�E2��4i܈j!�$^>t|���	�.�8E��	k!�dF�qL��7Ê� 
E���Ӓ8d!�Z�e���$�9S�f}��KX�!�0����C�0Y�e
��?�!�Ĉ����!���B��]�"ʄ$!�P5q}�̱��Q�1��M�螏C�!�H�5�\��4�o?���Ԉ^�.�!��<[S8i�!�8 W>�`���X�!�dd�2�iԅC(6�+��ەB�!�dH?SQ�	@�`����tb].&�!�D�\���B* �v�)u@�	{!���}�ƍ�'��*% �M��m�� v!�@?@g����
�6=h�Yb!�d@�_��0�zr���e�J�v>!�$�~�t
�o/]^��f�$%!���72�����
DD�y��یo�!򤎃B��	�HG<���$�~�!�DY/L�Z���`(>^ƍ;u�ܤq�!���P��%j����/�!��^8b�8��̒X����8ġ�Ė#/6,���s��[����
�'��i�Q*�3?=��أ�[+��8�
�'XpA"$�I2B< ; �U!)��'Z�@��ǳ(�T-��ȅ=q�~�'��i{��)�։a�ݚk�es�'��Q;3�C���H#��7L1����'x��7E]=�x`�@=H�4E�'K��x���,F!����W3? �%0�'�¨xBf>6�\�k �5�8�i�'nh<J�AH-F8) ��;�Fhp�'��\8`�ڔ�4�tVl���(
�'7�؊U(^*���2��*N��H��'
J�	G�)!9��o�	H)�9y�'�j�9e�oL��j�X�,���y�'E��RF���'������)��u��'X�����.W�T0��/�m��'�"��ќp���I7�)+3���'&(��_� *(-���J�N
�0
�'6ځ����JtP�ՠ�!d�S	�'vP ���\*�N,j.a��')"I�a�R���܋��
��	�'n�!e+���5$0�^�'�B@����=(�l�PFj�"�T8X�'��Q��2�`�:�$/i2�'fu@&��!�B�	��J�;�'��@��\�f�(1*H�(l)��'���"��=4�a15&�:`��� �l�u&�?�bX����0���A"O&�����4Dl��E�&��0�"O�l���l>!rS�-���&"O�Œ6E�&��A�����h�B"O�xYII�0j��P�����q��"O�P͞	EYt���7j�l�a"Od|�Ţ �R� �s`GK�JU\\�w�4\#�Se�A� y��Ф�', 1$#��V����b�.��`�'�����%ڒI�p
��C&���'m��s�OD<E��0�R#B�-]�2�'��5MӁ'���6^�A 
�'x�#P.ח)� �I�;2ft�
�'DVq+ �,�����/m�8�	�'�
Y
��B�(���(�k�det���Yt@���<ըh���,gR�T�ȓM*=K4$�2a��Q7�2� i�� �N�E	K '������2r�Ԅ�ȓ3:l�j%�	&	�G�H�:�؇ȓ6�P4�$�^}��swM�T:*̈́ȓ�X�cUG�<;�pÇII�z��ȓVr����������V	q���ȓ,��}zg�&b��%3ƢC��ȓ$�Z��wǑ����f��;���ȓP���A^=���_�nn���k�IS�4fN����	@C�݅�5�B�Z��b���Y�@`�`����	�0M�13! \���g.���+�̬�ɗ�e�$��1ًd� �ȓA3�`�D`L�) 0)�f�2��ȓR<HP# �6�ܼz�h�f���ȓJ$�# &S/$�H$
1��s�I�ȓG��I
Dɗ�m��,�BN��k=����0����!� �)�����J/k�T̆�Lo�T���&P$D{n����,/,!��ϙK���c�e,d^�����B�Xh��c�Z�A`؆ȓva�Ȩ��ƨ q �����>xj�Ѕȓ1��0j���:\�Ñ
��R������g���	�\���=1�z��	�ͻ��Z������J9p��ȓ�V�3���\�6�z�o��0^@�ȓ=�q���̆*�b݈1�K$��� �H9���O23�>e� E��uTޕ��<�� ��G/Xc�`AŦF�iÜ9��Bq�uҳFѨQ� A���.�T���C=X�h��D��4��+o���RQHD���T{G�;��ޡ}k�̇ȓc\���0�^9]B*4ۣ/�#Xm���N��*ō˲r�@���b��e��;SH1��n�� 'ԉ�p#ƞKp�ȓF4$A�K� ��0�$oW�(��U:n9����2�"Q4�T�,�H��{Lh�2�	g��ad�%=��ȓA�\�Ƣ2��N�	�,��)������������J����bВ�X��L?4\�u�P�X��4�ȓT�L�	�˝�G-r<���ËKF��ȓ`�J�sr����k�$�qXR ��L�:4R��Ê)`R�5����ȓV:�!kJ�0���zV��6��8��/��<86,�� �Tl��B�
!3l�����n'���x#n��u�pGaV�<a2�G��Q� Sxb}��bRR�<3n߿8��
`E?6�Cs�Y[�<� �$X��öT��)����v�D̐"OL���N|A�āӄ߾%���hR"O2ͻQ�R�j�� ��2"O&��"�V,8��0��,���T�B�"O�����	l������?�|y�"O$�IpC u>��b(Z�p���k"O�e����(�}qFR� ��<:"OH��߀/�n�R�ŏ-O���i�"O^�kE��v:f3�Dc�J�b"Oz��s@�I�y��=X8���"O*xT�
�zf�3&eԇN56<�7"Ot(H��ȈL�J�2��G<3<�s��89p X����M�N�"��)_o)6�Q.Y	Y@J@* )!�/!�5���ґB:�3@h tj(�B�	�*)q�=�$��s�4��BO5]�)�퇉���p�";�O��C��
�y�D
aV8X��j$�R��Q9bI�����f�	ـ��6����
c\ `���IR�2ay���x+l1� U'��J�,��a�x)dq���Q!�la��L!o�fe�'$�"`���c
�m#�<�F�֦{Gx<"��,|O� Q��W(q���`nT#'����LV�r�"׊�0bªQ�
��kw͐��C8S���b�/�0Ik�*g�̰��ͳD�:Y#(Ѷg)!�d
��.AC��5�yc͕�d��k���6UC4��񣑝2�V(�/���.QE�S3���f�W�C�9�(�*5�L�B:�e��-P��{��j���R�֦%9��i��U�%�H�8��=��FQ�
H��^����J� cJ%)E.��o��e�}�H�-�J�X�'Ĺ�E����'�b�*���\6����M=�C��b)%%.�8M�?/4�g���x�r*�N�P)���SN؞<�#m�/C��Sp ���l�">؞ّ��H?�?�`��J�C��-E��k�E�%�̕��5dQ!J�@9Rm�;1����؄�y"�Z� �N9���J�WVe���ǦE���K�蔀]b��+��|ѵ��!\��4�@�1\�5���O=>5�݀YL�A���{ABH����#J�����)`�ɡu�"6�!.�R@��*�'D�VT�seޤy�����N�her�/�<U�E�w�]!/�^\ڴ�f�
��Q��٢{��1��^�ι�=�'ʮP��@P���h?��D�>\l�z�&B�C�*r]�7JLw��p�Y�͓(zI�g�̖��=P��n
 ����I���ãHL�/v���@@oy2���7?���B����8=���̻qx��A≄�ue���ϊ�aOT�ȓw`�4�w!�6$�<�p�C4��P7��"x�ek�>��C�8��N~�i�ܙ�v��H�Lu1�41 ƈ��	�PP�����
�z�y���ߴ/(�:���O�d�G��J��Y�
ۓ�(�vL<)w�@;�^p�=�2@]{*<�O�����}'4��޴'H~�1���,F-��� ��6s\�ȓ��P6D˫M�v���j��T�"ȩa-�ɰU�*رP��dB1�&�ͻY��0�ɒ��	`A�dϜI�ȓLƘ����A{wN�����8 �Dɮ	�ܹO>E��'g��J���4a�L����x�x\p�'��倱.Шb~��ãNoo�qc�'�B��K�_�, C�Ͱxfxl"�L�����?D�P��-�kߺ9i@J�j�P�i�!=D��ӥoG<V-lT��.� C� Lʑb<D�H�7c����L�)Xb�q�t/8�O�M�'C�	at�Ջă�0i��ݗ	A���'�>��`Q&s��6�D�^d� ���S8	i*��O�JTd�G�q��M7xh�U��'�h(q'Aа �QK#ރ��3��w �)�6f�1�����"~r�A^-y��Z��@
(���fNF��y�FV�a��ƏW;+�.�����Co`�I�j�~���M��X��H)�����Z�,S�	�u�D�D7_�m`Q�*�O
,��TR,�y��MN$=����
QI?��V��i��T��-�OT��6-����鷀�!uWBeh��	�w;\��F-������ U!tV��,$�և���̓w�|�ȓA�5/�P�G�Z��L�q��\5���@���yܦ͘1�Kt��?y҂�(d�dp�+O�x06��!!�s�<q'��!�z0)%�0c�%J"�R)tז�"�G�aW(c6n��!�>�'K�U�{2(ڕCH����C�]\x��b��5�0>��Kx/�B�m�"v�<�x0�L�X�������Z���9�����,��o��=��$�(����	�++"��3�m�Z�J�����O��d��R]\pC��I����|� ��Su�R;BNٳ�+]�B��h�&d+}r��I�V9�@(��$�	J��D�&�7�Z����?I����
I�i)�	�*��^s ��
!�'H���T��|���*f��0��F�/n,�0��7�O�m��C �<����v��0)ȥADB�.:l���k,�(pC�B.�N���#Z
��i�!8�\:"/����W�!���/�O  $�� r,j�5 �X�J��P�[�(q�a�}ya{Bnկw� �صO �tr�'���bs
�L6���Gf͹F2��c$�J_�'��\���h�z(+#�w�n���X>�9W�PO��s�\t�|��Մ�\��8/�|�jKI|�3���Л�@�AM�r`�� d�`|  @�*dAtd)AdbL&�'`50 跀��G]li( `�8'�Pm�0X3�C��6�O�P���"e�"��Ռ:1,��#�ʥp�)B���\�H�ӑ�C���t�"6/�>_�Lҧ5fGK�?����G[�Ozl�a���>��h�l��tфҾ ͌�j�+�?Q��Id���-;,�#�L�+7���CU���Bb.�'lQ>�H��� ��*�F�#y���ۃg$ғ<!V�@jH�JR�A�<����[�~p����-�����oߩ0��O���O?Pg
$>c���e�%:7�'��/֜25.�O�X�Cc�y��R���~��	SIX��KP�-a�%��*�B��Ӹ7"B�IL�.,����-�$��Lܟw/��'[�1PoY8>�Z��%�R��%;�50��cG�	w^�:�-O�I������0֕��\N`�@� _�u��ixF)��x�́�]�~)����>sh�rE�T��(OH����!�'	���!E�Env`P�T!;��������)ӯw��r활8`�����0�6�"~ΓI��=2!�ߚY;���e�C�L��q>�5۱�B��	R�֭Sh���.,Q�*�O�h���n/�I;榀�K��i���'�p�e�[n?���,PͶ��b�I=vx�t�)�W�<�0J2 Q���M�((92���M�'����сTH�OC^��E��9q�ܐ�ᑤ1���	�'�@H"V�]�\T{d���&��e�լD�a���=E��'/����FQ7
Ox��G�3�vi[�'��3�Д"���34aU �|;�'��a5�'38h�Y+`���c�[�(���'� ���u�
��R*M:x�@��'��=x��-kp�h���_i$r�'J^�R��Z����tE�R�����'����% �m� F�U����'(fH#�	Uo��q�S&:�@��'�L!{�N��=: y�S�m)��'y��ydyY�|�cN� M�h0�'V�PH�A�S�����)� �'�v�$�)%E�ɹ��D0*3���'В-�C.�h���ƒsC�a�'J`TɥE�L��I��`�f��Y�'F�XU��8 m�5 �AC/���q�'Q ��0�_ ;�E�r��&%d�}@�'�B`���7u�=pg&�5��'��p ��Z��T�r���G�>���'��(���J��j�nK*�Z���'-��S���?=tM�T�zfdb�'���d�ƶS����_�t
P���'=��ȴ��!ꉨ#��j��L��'��Hbu�� �T\jsG�5^��2�'뜕�$�N>d��@S�IB��S	�'��p �T�,
-Xk�!��]`�'��r2Aϖ ���Q@���44��'"���w��:d�F=y�n� MW�x@�'� ՀT+�9�hu۷�3pA���'�R5��@ݍ
66��7"
�&#��2�'��8�ܿ<<>�	f�
#���a�'�D���زh�pDb��' N~8�	�'���hF 	��p�ͩ$.���'|���퐮0���&jN�z�'�b4�D�&2tj�T�mR.A3��� V�"f���8q�q�X�R\;�"O�%K0MJ�"l�$�" �B}��"O 	8�G��j �����D,*��̘�"O$�P�ި)��2�Ǣw�-�W"O�E��ʼ}6ƙ
��B��ՙr"OB-赍���C3��:��.D�x����*�$��&E
�Z���(D����cݺZ#�����D����B��:D�D�(�(n����A�	;p6D�X�S
e
���,0�V��CE#D�0��Dn��Ԏ߿n rYr� D�� T T$Q"�\�XL `�B;D��P��dj�3�//��{�,D�8�tJD�]j�R���i)Qd9D�t�ЁܶKƌ�F��B��XI �4D�Ē �@���@u\,~��1��5D���("
4��Ъ@�4t%Kƭ3D�sE�H�j"�ik���4 �Ũ.D����ӟ6��!j�@�;,�S�+D�$��Y� �V�nй�M2D���i��x1R��׮?rx�11�1D�xB'��$W�عP*՜;r�Z7`,D��j�N�<[�4��i+v�ʥ�t.(D�Q�nӈ-0�l�7ڶ5B��&D���d�2h��;%���qZ����`(D��.Y�����MZ�1&Ĉ�,N!���_N"Z���<v����KնT�!��X��,�6��5�SS'O�
+!�dI�?M��b�I��>�������h�!�DK.|VE�f��k�d��W
8]E!�$�$�V���m
�Zͼup'(�-,!�dL67gH�J ,K���4�' w.!�Ιj1zz/�o*�&'΋!��ރ �x�V���c�T�p�!�d�$!s�!��݃+\J����ʏZ�!�d�<��aꆧ�yL��!cj��	�!�D��ZXzT���<bl^�c�� !!�A1]5�X$�Z!%]L���cT� +!�ė�c��<��X��r�ѣ\
!�d��
��@2�VT�>�#��8!�!�d�;�r��X�u���[i,L���ސ��B߇+��Ty֢RK"�9�ȓs��� �G�t+(ɧ�BV�=�ȓR;.�a�#μ7y��0��_
8�l��ȓs8t]S�g�<utyآ� ul�	��^�(\�)O��s�'Y�U���6R��2�-U��]+f蚏��-��;�D �"L��b�D��4�R�C��\�ȓ|�D:��X�k�Z$Á�F�8��ȓ3�l9��ůf��dAW���*���ȓ'O<�p$�"��HT�{)�Q��
鲘[�J��W�Th��e�+wV]�ȓ\��̓B��|��9@q��GB͇ȓ*�����ёk��k���B٢��ȓ#!zaY�Gד:�B���@-Jsx���$2�A��%6mt1KW�怼�ȓ^r�aYV��'&�a'^�r�h��ȓRb�����-&���H��k
���� B����G��a�,F[|؆ȓ}����!Z�JX|�Bgˊ�>�ȓVW���e)	;QdI��d��F�(��Q�h�@��72���օ�V!�0�ȓ)ƒ\ȳDH=�� sv��NI�܅ȓQ�N�{��\(s��Ȓ���42�^8��S�? Px���'PS Ց�	�^$��&"O�����0k�|��jG2u�Ӥ"O�pG�L R!B�M��Ȳ"OF���@	 �(�P�O4d� 1�"O�xCejA2E�6=��G�J֪���"OTq:��,p,`I1���~��"OL��u�]>;8Ĩ�O0FƪPQ#"O܄���S1Q��`Э�z���3"OD�x�#��*�<yr�X�H�E"Ot[�ߙ*H"�y%j�C��Ĩ"O���e��$`�լ��8��	�b"O����Y.�8�)V��2}��"O��A
�>�,;��Xl���"O���ӯ^1j��i��U�qG*�a"Oebwn_8b%ԇ��;~�X"O����D&l��Ir��4|7L�4P�����&m��Yb�N�$H�*F6&m����Q�!��$��jb,ϤqQ����TJ�Z�k��$��D:G��N��s��s�)D�|��r3,�:wJ,�O:��$�\��y�-T�\��]�Q.}AFA �@HP�ˤB_ԭq0ER6c<)���D"����T%۷�Ao\|�`��Y��P�sk$=����o^t� G⃝]�"塀�v,�;��N9@���B�aut� �\�A�R�ɴ#4|O�L1'��-�t�Y1,2�ԹC��p�����ޟ$s0n��>Y�|aWň(�l�	A�F3�ȉ���c�D�&����G5v{��C�U�<	D��Xc�*��M�����Δ��$�tK7C����o�H�B��@.�"Oe�XC4j �H����
������1U{�ĕYr���p�j��&�2�k�NƵ�M�sEXlv�z'� .O):�u�;R���fg�#s\�����"_�n�S�iz�!���Y�` ��0,ϳ�����Eܒ@��O��c�Z�h����f$]�c
� ��)ۖL�7|�`{2�#3	X��&��QJU���I7$I0R3`E;�=a��/4�t�H��[,�nr4陽dg��"��
f
�H� B���3vF�.5�x�p� �.�z$��ؼdbk@��$�)sfF'4�T���'M�!�$��Rtm8�$k� �鰥Y?O�"�z��ІeEԐ�6.��Y��Tl�Vp}xvd�o����?M�g���ş���5@� �d��{�O7��zVJE��K��+B7�DLݟZv����ΰ&)d�"dC\0C����E��=]�C��A0�;�}"�*���Ӻ<֦�C��D&��Ex���?�j����O��3#���A,���%��nĳ�G@�O��B4��CX�s�0O��n�(F�J��$��3!��L�>��0�ǳ��*�a��M��	�J�+p��BJ��2<~4ka?��x���/7��,s$
�;M�x"Oʽ��^���H4)�<����*xr�H@O�N��#�g?1��A3c��z�X�X�p�s�&g�<a��Mb0��'С[������ޟ��TFRw���'9���a�Ƣ"l.y�&(E;9�L=�ߓi�^��ËՑ=�7M 35@�����\(/p�	6�٢|!�Q7�������z8z� R�r��OH�7n�"h�ᩏ�IT�\~8�BSg�s�|�B��ܞ^�!��,Y�,��so��Z:�iTi͛]�hŲ�o��>�4�O?�	w\V�Ĕ�P�ΤsA�0�pC�I3pL���(����4ˠύ.(�ID��}��'����	\Ԕh���*z�f�9�'6�,��v��@sPc�,ޖTs�'
f�3o�9*��CRD����@�
�'.�9	nDrl����B	
�25�
�'	&���O�l���2����{
�'��0���"y0�)��m�l��
�'�:�B�̏�F�
�a��ذb��4�	�'�h��;Dg$)���(P���'� �y�-�b�F��@��:��@�'Sޭ��S�9���[ �
<2
ɱ�'��ġi�6X)�g�_*O��D8�'T�UFV�kjn��� �s��<�'u��M�1���FN
�j�~m�'�D���$->P����<d=��b�'� ����f��hѵ�� ^}�,y�'Y��ӆ�.��qRҎ�J�`�`��� Ȁ�҉ɞaC´K4K� ,�����'M�2�bܓBc&@� �Ւ��&^�C��)�ȓl6�x�E�3����`H�`��p�'�HBBC�  ɧ(���B�K�:{~$	7k b����"O`P��j���q�w V�ߘ���!&}� �S�-��C#��DG�u���yV���>p.a"N�(�� s̏�m��d2pq$c 
4��0��ɹ)��hkC��ڔ�����C�T"?������ (��$�����<���#2eR��Ɇ�k�!�: '&Yê�4Mh��L �B��I�T�����.e �S�O��4�T'��͘eCY�b��M�S"OT0��E�e�p�v��p�� }�A�95�.q�f�&��$�P�xQꗮj��A$�aB������g�F9�ayiU:��F>x1f���	x����S�� qRX��'�h�#?���V�,��(�Â:�IZ�L](�R4� 6�� FȌ�!򤛴I�x�#K
 ����ٯ=D�I;^B�P@$4��S�O����艾J����'�H���l/�"a��17)ހ� ������N����L�W:��3I|�>� '�hD����
:��𦇘X����@�X� >8�T�7��e��EU	EiꌡA�SA<i���{ўU3�� (Z�����c�ܛ���~qOƔ�e��4x�Ujf��F�b G"O(�0��[g����QL��U�
���"OP݁"��0�(�'�E*��́�"O�x2-Θȑ�1������"O~�y�%D~-��G�v���"O����m�)4�١6��AȾ�1�"O>��dk��=]�KR	��G[�(2"O�uӖ��y"��"�"�"\X-b�"O�W�7e$��3�ĵ�$��0�>B�I�����M1(lx(u�F�a�B�I�2�}k�͔�(�(��޸pN�B�I<C�e�F�γl�ș����E],C�,R��YDJ��"�چ�C0d��B䉵9t���3�.Q���hD�Z�U�򄊺r8&B�
BHI�F+D�r!� �h� �e���p��`(��v�!��\�*X�Q ���ܒu�X�8�!�d�͒�`�j\�d�̸[��B�|m!�D��Q8�F�^�K�@A�f�S?nd!�dˑ���R��6h:8����8E!�ğm��e�#n$qy��_�F!�h�DY4�P�f� |BtC�wI!�ܘ�����-sc��a���T\!�ݾ�jcc�yH��
��9�!��]�P���L�w�`��!/חa�!�d��v��1С�D�VH����J!�M�Q�0� �dșI�2؀�e�4"8!�"Gt(���(!;���3���\!�K�z����v�C����X�8!�a������rG&T`5
D9!�$	g:�}��F�<�p!Ӥ��J?!�@�.�R� e�Rs������h
!�͸8�Z�B�&5^�(�"X5@!�d�$g
4=A���/[B �k� ��T!!��2�xD�E�v��{#%[/3)!�d�8;��B4�l��Ń !�$��cR�����	�2��Q0�Y�!��t�NA*�/�.�Ƽ��eA<|�!���
@Ϧ �dhA3;�2�Q�J!�ۈm���%�Jr!s[�QK!�D8:w��P���m쑱�E';!���3��|h�N�YO�$��$A�#�!�� �U���"{�b�[c�]�f��=r"O��r�+рix����$��0"OƤ���!z��1��up�Z3"OR�Qt�]�m��܀��rTtI�"O~PP��;1-T�Q��!��)�"O�#jU,r��1Y@��` z��"O�t�B�չcE��i���+c��"O�5K��! N@HMQdR�4��"O|��R�PxQ�[�~�G"O�2�	�qP�(35�
!~���b"O�P�f鄢#C2ݚc��5�,��"O�d8�'�-�>MZ'#٨M�&@�"O�M�e���%�F�3� ڌ/�UpV"O:kG苒*��u`���(�^5�1"OF9ҐG��f���0�A>��Ш3�U�
v�6��
lx���'ˈ�i���i����q4���	�'���B&Ξ-vb��1iΕa2��I
�'�Z��C�]C�&͐F�P�R��
�'Y��Z���Fk�3M ����'�$hI"|C�VI��<�Ȝ��'Z\�A"�]c���5��;O��y�y".�'��'�vc>��$��'t� �k�ʔQ���mϵ��{��V�qO�>u)7d�?�n�a�藐Vr\���SrBT����6�|zӈ�o�'l禼@���+}��b��j�~��fN���xWpyR����O?��*48�f��27V�d�n�;Z��J#�S ��۸v2����W?�E���΀n�����+g����Lٳ>:��'�\1��g˜����.�>��#�Iu��δ-���'[�@�b�iaL<��v��n>|�n��O��I��!WA?��cH�p��y�$]��'�;�'hn8Ȃ��=D����!BzH=�V��,�
�Kd_�$��O�"� �c�LĐ	ҡn4}.^Q`�>�=���pU�%��!"rK� L�QPU'A�^�)��]�<yѴiK`��4h��1�8�KT���uǭ"��~�Z��ˠ�a��#������-E
���ћ6��U1B�?��y�G�\�K1�YQ�I�Jo�1�@��yȁ��ڕ[���&X�Ua�$�1H_����2�h�#
�, 3"���|�$�Q*�:���

�'S%�,I#C��
��HǊ�.l�t�8E�O�P85 �V�ve˵k$���ůi]l�x@�������|R�X8���?%?��7�O�W)ޜ�w��<�
A8W�>D��I���)`1���t/�|�̰Bc=D��C��t��Ӣ��2��dk$H;D�(��/}����@E��Z���.;D���aj³��A�"IQ�!GJx��:D���qN��I�tJ�x+^�a� >D����\.H40:��C4F�LX��.D���5�_�L��!�t�ۑ
>:��	.D��sG�����$o���E>D�H��@>���S�[1a�,1#�(D����)e�r�1l[/$�|�Â*D�����"5J1�T.a}z�
K'D�@�c���� �r�F�xhh�� D��KP+��`�l�;��E1� ��b3D��h#�4H֠4�rK�\��X4e6D��x�K�Ab��Z�ɒ�Wz��R1�.D��C�	ż"��xh!�V�7��I��,D�4p ��#75\�u �2�]���+D�T�šM7r4(�@�&��o�h�;��.D��s㡇�a�fD;��W�p�"d8��+D�<���[�7��0��L՛<�� �H5D����%\4��б	�P�a��4D�t�FÝ/t�S�ǟ�b�$1D��a�I��J�����$��X<�v�0D�(�F�7&�@I��e��.I��J.D����<y�\a�m�d��y��7D��h���s7����n�F=���+5D�`�g��(=�Pdq�\=>�U��1D�� �����I�d�b-��m��4;2Q��"O6y����V@NГ��,>/r��"O�#��A-��҄��f�vT��"O�9KBn�,A�ug��Ȱ�"O2��g��6U��XI��u�<�9"O���0N�@1QGKԷ�J���"O.��.�$$li0˞���Ը4"O�����S�X�A��98 -r "OV��`�Q�C���4CR	l��i��"O��s�E@g���DƯt��"O����D�n{6X�����U�"O"њ ��o ��j%�3^�V�W"O��	P ��%�X]�0��.�IP"O�"��"�0���i8:X0"O��:��ٱ`� 슗�����"O�L��b��l���ya�1x�zġ�"O�!�I8�� 㒏�S�X�"O���C����)�qA��c��5`Q"O��IY�1��iҕ+9*Q�"O:`ӗ��'Z���U&j̋�"Od]��eQ%^X���æ 4�ԍ�r"On�RsА �t 3��\<*d�%"O6�h�\3���N�"?���"O`m����&Tth�M@tm|��d"OXs��D!(��4Qd�ݗ 5~1�Q"O<(!c K'��\S�-B$ȃ"O �)ٓx�,��1L�r�\�*�"O*��C.��,)�Th�(;�m��"O YPp�˧l1��Z �Z?=�1�"O�1	��(!҅X��1l�rj�"O|�U�c�P�xU�S�ǦM�"O�y�nM7��<Q�Z�NO�M{b"OڰsQoĪ{׊I#�C�]Rxy�&"O���ՃvSB PQ��K�&���"O����!�5,j0���8��"O,��3�H
y56�)1�B<V��+"O���������Y6� �Tel��T"O2��Q�B�+Z�:B��b2���"OvY1���(R����'J:D�����"O�L9�^3ltf���痣m�f)	$"O��$)����1��ΰ���"O��Z��\��D�OV3<�vIBU"O��b���Z,pd�ą�&[d�B�"O������c&��I��ˀy�8�f"O"�ȢMD�}���yS����EQF"OV�	��B3� ��EJ.4�x
�"O�R�ݬQ�p�X�E_-�2���"O�)��>*	���]�U�2,PB"O:�@ABP�'�L� IT%m�2���"OT�	�ᖤp^���'��/ij��"OT����֒d6�P��}g� ��"OzةF�K�oD����*�ht�&"O�誢N��x�S�޲tR���"O��+W M	e��	�c'��@8T��"OU�s�^8ED�\��E^29 TEʔ"O���vlC�\��0�d��H��;�"O��@,��'$J���D����/U��y�M�(�����(�ٺ�/%�y%ܕ5����Ά�"/$�bM�y(�/*.�A ��d`9gB��y��
�1i�J�Μ�w��L��`���yjS?0Z0e��� m`-��Z �y��9�
�鳊��e�P�+�+
��yR�8v"����k@�d�R)����y
� #�mV1k���Q�NI'����"O�3U`�O�Xq@�2t`e�"Of���	C�/b��ᎎ-ޙ�"O��`أܾ�9po�	x^�e�4"O�P�0L�e��l!r'�p*~p�"Oȱi�����_�v2
�3"O4��Ҩ���.$�тI'�v��"OU�!j�^�42�Hʿ�@��"Ov�0d`����)�T�u�4|�"OtIR5�U&�2���5��"O�1�$ 7|�-ɷd�Ws���"OD4S�b޸`1�X#��r"��"O�U"3B]�_�rP����oX�,I�"O(Iҧ�[	(G`Px�b�S-hU�F"OD	p&E�(�Y�!A�F�1#�"ON����-kt�	�:)*�Q3"O�d&d:ލX��r!X!�"O��U�Ğ�+Ȏ'�8�""O�� �"O5,��@��a�q@"O������3{)�Ƈ7$�>5��"O6��cbˣ (��bg�Q�?���2"O�`���S�g���N��/h8Iw"O��ǌL���+s�*Tҍ��"O8�SN�9{�I�g!�?D0x T"Ol��Ě}Ю�
���2t��"OĨ+�P����� x�T A$Ws�<�`R�O�T�s��l���"e�!�d��ZY4��g�J� ��\=d�!�d��,�����I��ru�ɨ����r�!�Ċ6E��Sq	T�!������6�!�$����iw���J ���a�9�!�X<8l��a�'�U�,�h���^�!���8e ^,6�^�p�J&�2�˂"O�a���,bPn�y@�J2=�)k�"Oĥ�E�2�Pi ��TZ��;6"O�q�vM!jU�l��ϒ&X&��"O��3#C |Ubl1U���P.r��"O��bE�ҩ�6*лY"Ag"O�(�A��v#x}���*�d�{�"O@-+ ��!j��i;�	H�zϬ�2"OB�i�'��L���Uȕ�g��P"O�)[�F���%���Q�=e&��T"O�����(b.Xa�TfB�e�8Y�"O��%iנM�T���dߌF,	 "ONݢP�>��HB@o/ �I@"O
<�@�5�M��'"w�A��"O�	p�HR�df*��"��U�,A"OF��E� ztbGӘ(J m"O~<�1��*��hq���.)A��7"O~b!AE�Y[Ԑ��h]!l7�P�p"O��v��%s�䣳G�y�p	) "O(�9b�;%��s�N#� ؠ2"O>4S��3� %���1�(�"OލcG��,#d���a��&sS��he"O.9�b��?aX%����Z%"O$Z���k�E9�쀮� qI�"O��A��װ^���&K�!<����"O`09��4�RXx��_K~B���"Of��T�&m��i{�(��tk�=��"O@�����?�Ƥi��4Uc��D"O<�PAe��^2���gWZ��7"O��ʁ�d�*9C`�)6�%Q""Od-!�����t�Q/L!p��!7"Ot�{V�7fm��M
�T��w"O� ��Ik�:4�FuI4��=V�b"O�D�w��%��)Y�A
r��"O�@3`�_/6(��
s_(dN)2r"O��� �x���ES�P���"O��I�ZO����j�O�4��%"O�5�«
�`������Wb�dH�"O1���z=� ����2'�܋0"O�1����4� py��	8�@�*�"O�tȃ�Z�a�V��Mf�@8*t"O�]1Q�D5Lf���P{�icR"O<�zr���>���"@܋d`��ۧ"OX����[�2Uxv.�'D��0�"O��+-��8�FL��
B(y��HW"O�P��(H4�p���3L���t"OD`ɡ��+]E>�� ��6ED��u"O���	�.�A�ă�m4�8�"O�r%%�X���s��>��f"O>��d�� �����	H�x�"O��3F�!8cb���?�B""O�4��20��t�V��B�raXT"O�KS�C%K�,x#[+R!0��"O�X �m/5�r]�Ԣ��=l�A"Oֵ[�Ü�K[X\��A�2C�0��"Obو�A�8D�Y��ҷ72ZxZ@"Of�k��?zy$ �t�F-�Đ�"O� �a�][+ Y]�)K�Ϗ2�y�	P=V����_{�ْ��[�y"�OC4)���e�VY�GB��yRF�m'|]�d^�d�������yb�*/�hs�]�Z��d(w#�4�y ٛwT|��(�=X4�CN� B�I��l�" d���d�'��$N�8C�2e\����C%,F�;�LC:��C��%|��؄卸L2�[w��u��C�&M�1��-�F��E E-�\C��8�^Q��D�8rG-����uC䉀:�Q��
ބj�2-�G¨WC�I.�����@�^L4�@E���B�SUQ��!�8��a��S�`B䉯{T�\�d�>s�v�rO$t�8B��/a��a���-t�C ��gU�C�	�Jꪩ!��O�u��)CA -=�B䉑I��6΅���uX4KK�.C���4Qj! >oyЩH��D�@� C�I33Cd�   ��   �  ?  �  �  �)  5  E@  _K  �V  ,b  tm  �x  ��  ��  ُ  ��  ��  M�  ��  ݯ   �  ��  2�  ��  ��  -�  ��   �  w�  ��  ��  N�  � �	 + o �! �' </ 28 �> E OK �Q R  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+!��6*\�c�<4�d5h��'�B�'���'	�'/�'�B�'���U�W9��m��Ʊz�0�b��'���'�2�'��'�b�'�r�'���k��.Kªa��͎ 5���Ha�' ��'���'�R�'���'���'����
F	�>]�&ΏfEP$�b�'�b�'��'�B�'�B�'O��'�$��zm@|XpjC�6�D�'��'���'v��'�'��'�"1�)ֽⲵpa����j5�'���'���'t"�'��'��'�%؇�Δ*��� A�B4%
0��'�R�'��'o"�'�"�'/"�'�f}�b���Xs���]��X��'iR�'���'���'��'W"�'g�=��'��"��	�Jw���'���'j"���d�'5r�'}��'��u�1� (iL�\r6e �t|:\���'�'H��'J��'ZR�'vr�':h(uC�=��)��G-P�����'��'u��'}��'���'u�'�;+�'HhufUmzn��`�'���'|��'���'��'p��'�J���R�h�����*|h�p�'���'��'���'h2�h�x��O��"�q�R��t�T�)����G$�|y�'��)�3?	��i�&��#�Zyf��B�º�1x�I���Ŧ	�?��<���i�X�p�ޚn.�R�FO�D>����?!pm�,�Mk�O�S��K?�Af͇2m����K��CS��ą6������'��>M����I�,=Y�fɝ��Ud �M{&%�e���O�26=��H�N�:Hm�y��[^|<	���O���n��է�Oj.��ѱi��R:28Zݢb�"bw��:R(�3��$t�$*�#��=ͧ�?��&ޙC��Y�S\)��<1,Or�O�Em���b�����C�R��f
���"$��Q��o���ޟ��I�<9�O�A1���X�`,�wf�;��"����	<���U�;���B�����z L�4�*H��M�+\�����my2U��)��<��%�	|��0�K��)��i��	�<	b�iV�|�ORtmP�S��,P}b���J�.����g���	�x��5��HmZG~"1��)�ӳ@��˔kJ>L�b}�Ul��Y۰�|b\���8�I��,�I��H������eЕgB �P�[Dy�Ooӎ�2��<���䧊?1 I�D+!�e���E�Ȉ!�N�<�����,��L�)�N,�*����d(,�Ƭ��R�;Ej���-O�4X���)�~�|�_��!��������_�f�.8�!��ܟ��	�������{y���Ox(1��'�����ˇ�?}l|K�O�A�aR�'�~6�.�I-����OB�$�O���c,��£,į;��#C�&JL7M$?1��J��I*��߭iN�F����uq0����f��$�Ol�d�O����O��$<��Qv���h�`K���C&�@!���	�����/�M�իK���d��&��2kY�1\*�����
�촑P)@�柴�i>�c�`�٦��u�n�,���������FJ�{l�-����q�	{yb�'�2�'�R�{{��*mˋjm�JuO�2hk��'��	)�M[p�˽�?q���?�/��|a�⇽l�.t�9r�	F�W���"���O���&��?I��Ik�6mS�lG�H��i�Hɑ��(Kf@3%�N��|"�L�O���J>�� �5|�5z��V=u���a����?���?I��?�|�.O�l�7)�ys�Y�Bq�ayGHʾ;)H�cf�ޟP��
�M��B�>���,��SW�J�J�� #��U�Q���?��\��M;�Oؕ1"�(��K?��^'�QRD���y�%�|�'f��'��'�b�'��S�KŨ��
�bE�b��Yf�I�޴�������?����䧵?) ��y7�B9b^f���<B58-2�#G�9���'�ɧ�OG��d�i��āt��0SG�;C�%k	;�yR�3~VM������4���ĝ�p+�I�l��7i*)[���@���D�OB�$�Oh˓\��,4�r�'��哏�B%����8&+N\��ȩa\�O��'���'#�'s�%`��0�މ�H3R����O����!Z/x���Q%�I/�?%L�O����U��e ؎AJ&�j�O���O��Oj�}���u�b���S�#-8�C�G%.�l9�v���Mz�,�	ҟP�4���yG��*%~�@w-��8�����i��yR�'W��'��;�i��ɶ7A0H4�OΪ��K�`��|`2�n�B�&�HA�	By�O���'3��'?�(_3}�(1�'�4�D�c�T�J��Ɉ�M��$ў�?I���?�K~�Ch�kSA�Db�I��%[�*���ɗV� ���t%�b>I����LE�p�,�9;���5�`�����#?�U�^��(����䓟�J%7��Ѫ�ͻe�rU���D>&���O��D�Ol�4�f˓T����	�S" 0`��k3,�eTJ�����yRzӒ�h��Oh��O���,9�)�i��:��he��F�x}zӠ{��[p%zs����>��=� l@P��A]f�x����*�@�@4>O���OR���OR�$�O��?U9�.��o�Z�kʗ�'� �e�՟�����Hڴ/<h�*O>1nZN�ɇ_��<���6b����)2�z]$���ɟ�1%���mZK~��ס1ސ�dK���Z����!�$h���i?L>q(O�	�O����O�+ש��-mƨ+�Ʈ9�v���c�O���<A#�i_,����'?��'9��u�<i*g�܌@��-O+ˌ�&*�I���d�)Z��=:��	:С��gS֭	�,5��V�Y4�Ms�O�I��~�|"�_�W�m��(V
Q+S��S��'�'{���T�D�ݴ6�Ũ�af���w�ѿ;\h������$��i�?�wY�l��ԅ	�h�.8~Y����ob����ٟ�2%�ݦM�u7�V.�����Hy���/uz�H��ݹ	���7�6�ybW��������џ��	��ؗO�lHk�+�C��9��IЂK��yYS�o�Q�r��O>�$�OT���D���睗I�B �`�M�%�Q$�EM�x�	���%�b>E�WΦϓV��H7 �Eo.Q���o����t����f��X&�|�'�2�'p�ѱ��H�vP�X	�!^>� 7�'�R�'��W�Pcش"���P��?���N��!���ʂ]�VP���(�,����°>����?qL>�`k 4v� ��l
�Yf	�a~b�E�����Β���O����	��ֳE
���Q�O�|�\�Зg�	6�"�'|r�'Pb���#��c�lX9f["v� �"�dA��k�4�|e[��?�7�i��O����)E@3c�
��� {��D�O$�$�O�#n}���A�E�Pf��h�C�L&��!���:_��9s��\�����4����O��d�O��D�T�����o����W�-o�:ʓ=����	5*���'�2���'ܸ�*RkX�my�uSu�8"��ų3��>�������O|r�8 �UE"@�pg@�U92�An+H4Z1��V���t'�����H�{y-��B�~E��cw��@�����'��'�O��ɘ�MS��G�?Y�ʚ�l�x<��¤P_����?Y�i�O���'��'j�f�ahY@��Ǉo=|�$.��h�D�մit�	��2��q�O�$?��](q�����Y
�M��#���ݟ�������	ݟ0�IE��}��Q� �̤�����b#=0t���?��tg���.�剘�MSO>yq#W�$h�!�P�تuj�{qiG����?y��|b�B���M��O\ܸ?D^�u��&���m�Q#	�eٜ�[�'��'O�i>���՟���<r�J k�NT5pt�0b���v�������4�'�N7��9D$��D�O ��|R6�ً\ˀLs�MH�dI��#�-�g~g�>!��?�M>�OE�B�oϷ:Ȅ�� �S�AOHi"qd�<t���K�N����4����v�b�O�\뀄N `wX�ʧ�� �.}�«�O���O����O1���	���h��;�T��ܿ/�l�$)�+z蠳3]��sش��'���?yg�R�Hސ���,e�e��h��?��H���۴��� 䘠0��G�"�`8�oĔJ͜�L�/�y�X�0������I������(�O��9s�_4}6<hY�(k"��Ovӌ�˴��O����OP�����K���ݿ��h1ȕp���E�(�Z}�	�8$�b>�!�	���̓	�FI9enF�x�й9t���\�d�ΓR������O.��M>)/O��O��S�PX�����ud�r���O���O��$�<���i�Mq��'���'Ͱ�B  p���낯ˌ(��� `��Z}�'G�O�S��G�D��D
U
Za�������-$����B[p�/%��B�".��M_�c��jxy@�	�ܟ������˟�E��'5L���۪��	P� L�S(ܐ��':(7�ޖ����O� lO�Ӽ�4hچ��}ࠊB7 �J����<���?��O�(�ݴ��dȷ2�h��O�Z��`��lk���լVc?���`�|�\����ޟ��������⟼7Q"4U(e�E�̼�I�Bny� }��5���Ot�D�O��?Wr}�I���%&��Q�2�Ӂ-���?I����S�'}�*J� ��}qLIB1$�~ȑ3$h���M��O�PFN� �~��|�X�[���	wG���j� �a�V��h������Iߟ�@ybn�J cK�O"�Q�)
�z�Ҕ1�!G�O�ni3�J�OD�lX��.(�I���	���/q�@͓g�8�`5���U��DnO~�,R2`�`����'��k��U��
43���lw���L�<q��?����?!��?y��dO�(b0\����M�J��L�T��'VR�}��Y��:� ���æ&�l0���B��e0R!�y���u�^F�	��i>��E�ͦ��ug��:0��M��	�=��5��M-����'��&���'���'F��'/��pA����d��J2,EHHF�'6�]�Xp�4NO
H���?1����)�.
0P���l��Eb����	����O"�D%��?aJ�B��r`�Snʋ8l�mSb���dqT��U,�-=������{�|��|%<P�bN�]�Y�f��'i�r�'b�'���R��c�4(}��8�/E�$d�ȊM�st����ǎ�?A�Qћ���t}�'�V�:UV�R���Y�BƔ:�̬���'A��V#L�������gx���~� x8�@�Vqr)"�	űPh)�9O�ʓ�?����?���?9����)H9m��ʲf@�!��%����>�$�nZ�\� �����P�S�h+���#CAG�QX���%��u�ҭpu�6�?���Ş2����4�y���A��1pFHQ�<p�G�א�ybigk����%~��'o�i>��I"W��sFO׃n��BeA s�y�	�`���� �'�7�} �d�O$���T�Z��Q�
H��+�4�Li�O����O�O꡺5�"p���_X������n+x�g4��n/�g�����֭8oB��vCn�A��ҟ����T��蟐E���'q�-K���5}�H�Q�V�@.<X*��'�6-U�]0����O�o�B�Ӽ;2f�9j�f]؂b>;�)���<�����䀨N�6M/?�c��Y2��ɕ96�N4�B,X���Uk
N�'��1)I>A,OH���O��d�O2���O`5�h�֩��� �b�C&ļ<��i���T[����{��a�x�d̔�6I�0CXi�P�D��n�Ş<�$��o׀g��ra��f����Y�{�|}:,O�)+dG.�?���9���<�ͽ/#-3���>H�1� L��?���?a��?�'������x�����eA�)A�Np"bH˯Mn�d�T�4��'�듏?���?���_��+s���9���ZA틉h4^���4��D�5&�������O]wG@�-���Q�A�(�6������y��'��'C��'���M6?4�q �R�>�9�x	��D�O���XȦ}��
a>!��/�McN>q���+�Z���y"=Y���:�䓴?Y��|��e���M�O^m���Z�n+���dm�9*��	q�1��'�'��i>�I��Ic�
��p
�+.��t1T�F<�P�	֟ؖ'~�6Gr���D�O��ĥ|�R�6^�"oH4�$�PT�f~��>Q������Ud<��i���� �!B�Xe��#�
�Q@!�<�'/(N������F�4���Z��ȍ��%[>������?���?9�Ş���[�=y��3c�&�RBI�z�ٳ�Ǵt0�(��̟$��4��'v$듩?����v���9��6?�l �'ר�9��i��ɿh�����OGPH�'�t�F5.Rz��g��8��'i�	ߟ��I��t�I؟ �I{���1x��UŘ'�<���_�H���$��YP��'�2����'��7=���3UG�2*�z��#)ʵe�v��O���7��i�$}j7mi�PFB�s���shP4�!�k��9�J��=���'�d�<���?1��4��y����+:lJ�.���?���?�����y�GEVȟ@��䟘9�I��7?�H�M��X�ؑ��U[��M`���H��z�	#D2—�3猏_�����%:?!���u��#үJŞs���K��?��F�"��t���B�i\H��4Η��?���?I��?	��9�.QU��tIcB�(~BuX/^?��`s�\����<AW�i�O�N����� �#1�4'��`.�d�O��$�ON���%h���E&����)S_~E�F�M9&"HI��0�O.��|Z��?��?i�,	�U��
G<dV����R�Yl�	p(O6ql��Y� ��	��Ir�Sd��V5mQ,ep!J��[;&P�f����$�O���"��)�4��<aa�y��v��Z���a�G���˓H����f�OX�JM>�.O��a�Z�N'0���B�A��4+!��O����O�$�O�)�<�b�iь�D�'`L@ѡ
̔^-
Tj7�^�w��IC�'��6�%��)��d�O~���OJ<:�C�?rU���0�H�U5�����X(^~7-9?�C
Ғ��G����uTm�!3.Г��5��(ו8���O����OB���O��7���e�o�w&܁JU�E�����Ɵ��	��MC�o_1��$����'��ےm �R���Z\`�3�f�~�I͟��i>%zA���)�'���K"wj�(�qn�bDr�G�R/X�F-�����4�
���O����%^O� C�&���o%~����O�hޛV �9'F�ܟ�O���cu��`���	��i�h=��O���'�B�'?ɧ�	M�u�h s�A\d�����H�\���(&����d6??ͧ1��T�	G܍
����IW.�'�)ɞ������	����)�ny��x�L����]�m�mJD!���8QtJ�5`N�˓vE���DQ}"�'��HhR��JB�,��MZ�}۲)���'�2�h��v��pkׅR�/Hq�L9@QM��)����	۱T��y@g1O�ʓ�?����?9��?����I�'-0��bH� ��0�"���=��Qo�ŕ'V��I���]

�$`A3�̜sm ���f�}�$�	Ο�%�b>�f��ƦQϓUXJ��w�υD�
�!�!ZP@�e�z�\$ΰ��&�����'C^��@g$K�J,�`C�'�6����'NR�'B_�tH۴۸dx���?	��|H�
u#��~�V��v�
�?�Xm�� �>	���?�N>�DѾ4�Js�}�@�$�z~��\6����'Ƞ��O���I�;B��V��`  3���0��0C"�'A��'g��s�e`�kY+O���:І�ج�֬Iş��43J�S��?1Ӿi��O���dI�/Ǭ+ L��Œ�QM��O����O�A��e�R��h������ T�z���7�P�1Sf��8@�J�d5�$�<ͧ�?���?����?Ag$��J<���"�H�0�V3��$��т�GF���Iğl&?�j	��p�d0CKV�r��������O ���OܒO1�H�i�Ê'��<�e5|� UQ��#�$6�)?	T�\�L�R�IX��gy"�_�qf�2шݒ�t(7J�,]���'��'��O*剤�MC��.�?1a	�
j�DW@VF\����%��<9��i��O0��'��'$�%�y�g�D�[%*]�eIH=y��{ói~�	%!��=ٰ�O Ĺ'?i�ݦc@ܽ�V�ҵ%������n����������I�X�Iq��P&:Y�櫘��n�Q��< �Ĺ���?	��8ϛ������D�'R
7M.��҄�hM�#b��J	�)�,�= �O��$�O�)�,V#�7�2?�4��JY*(�UM&@o"��l�)Jv�� ��O�d
L>	,O�	�O��D�O�i�B�jn )�b�@�����O�� 9����d�O.�'i䠍�'�G�{��[so��\��'�N듌?�����S��P.%��0Y��ހ �ΠI���:vC
�SR��9N��%��O�i�?�3��L:c�(U��� � �j���2����O�d�O����<�1�i�r`Q��Ɣ|�8��˝�4�v|JG�ɀ��I��M�b˽>!�� �%I;;�`��ڽ�yS���?�����M[�O�D9�.����O"pP��ҬߪW8L���㳉Z�<�.O2���O����O"��Od�'�"͙�H�!�����9i0yC�i3j�:��'u��'9�Z�lzށ@%�9o�zͱ`��GJb]�Q' ����I\�)�Q�:ynZ�<��MK�\�ZaZ��Y�x}��BÌ��<ٕ�&���$O��䓟��O�D���� �њ+4J �r�	�I��D�Ol���O�ʓ�戙�b�'��L� h�����Ԑ�Xڅ� .o��O��';���8E�F]*��X�kN���U̇H���"��ۂ�%3��$?����'6����Y1:��gZ��j1�S����	Ο�	���IG�O^2�ۀ|꼣(�,���1��+���g�X�q���O������m�?ͻ4���	Cqa�uV�3'>�ϓ�?��?iG��&�M��O�N]�9%0�)� qv"e0����pء"�ʙ�~���ZM>9/OT���O����O��d�O+L�?W����N�=��yqJ�<�·i���Д�'b�'��y�.Ĳ!RhE�&葋��8y%+�;N�@��?9���S�'jr�!�P�1�ؽR���>�@JBi�9�M�R���J��D,���<�4���������V��1��O��?)���?���?ͧ��Y��Jw����df�4��l)�̅�48D��4�����I۴��'���?a��?�2D�>mHH �$��h�2�XBL���ٴ��˔K�+�'��ORצJ�H�´8c/��RA�x@m��yb�'���'�B�'����ǟ9�� ��߸��	f���U�~��O��$Gæ�OOyH|�f�O����H�t\�xyu
&P��2�)��O��4�y���f�v�#xx#�K�N���ffV$1�:�s��-6���	v�[y�OS��'_ҋ�='1�X�oF�?�z��A�5\��'����MC0�Փ����O*�'6���x��R�^!HQ�!�$=UB(�'�@��?a����S��mΉ�9x@˝�HŊ���B���$�蝴��֐��#w���8������Yq���`� &�H��D�Oz�d�O.��)�<!��iz��r�5&�.T�6iW��#��.4��9�M���i�>���(=�ȷ蚂]^�	�F�bI$����?�(��M��O�-ʧ ָO�l��`լ̒��؉B�A��'��	���������I�d�	R��D�w��اC˗R~���BZ	J�6m3�r�d�OJ��(�9O�Loz�yK@  a,Q���(*�,��	��	w�)��!`m�hn�<A�왱o�\��R
�ck�!�S.��<�
П(����_�Ty�O��o�ZD�x��Nk��$���^���'R�'X�	�M��5�?���?)t�Q�<*���d
of��2�k���'Yx듌?����=��y�`�Z$:��u���!X��'u��ҋ�H�FC&�	U�~��'؀���S�����`]�x?<U���'	��'��'��>i���o~\��bB#8 ����GnX����M�%��?i��2:�F�4���Z��քTO��ʰ/�j���3O����O���V�+tB6�8?yc�P56it�)�}V�X���ǔ�c#,P;��O>!+O��O��d�Ol���O�����O���o��i;���<�Բix����'Ab�'���y��]N*-�) ��(��!@c���?���$���N��s�
�鎘[��Y�K� $��<y��	gg.}��'��&�h�'(x��%t �9��;(��y�'\��'�2��tT���ٴ-ּ���Z}������Pd~�k���%���ΓcK����R}��'��I-m�8�ӂV���Bb��o"!�������'5�����?�����t�w���j�G%y���%	�A*ظ�'z"�'���'���'��R  ��6���$x�bG�O����O\qm,��П xݴ��u!��3DF��1��9CR�%�NtO>���?ͧ���4��d]�3�� ������5q|X�A��S �8�E߬�~Ғ|�_������(y���z/��0ևM=xo<��%G�ԟ���Jyr�~�V�(c��OP��O�˧Q�ř4j?��d� Es|��'al��?����S��Ș�Tp�l��N5N�z�H����qJe��8��x@^��� f�B@k�I5����3��b�1SǄU�ag`��˟�I��D�)�uybd�vqv �0BZ�1��H
BFɺ�m�C��D�Oh�l�c��%)��ڟ�C��/�Ԁr��<AuK�ߟ��I�xR�oZ~�K�,5�����A���y�f����K��T[�j� jc�D�<)���?	��?���?a+�>���ϼ|��@I�ȚW���=�"�ןP�	��L&?U�ɝ�MϻBc�L�2A���)�bf�%���(��?9H>�|��N��M3�'IP ��J�!Y�:�:�U�S�`��'�X������9��|�Z��Sߟ�ht�s��Jq�
X�,��ɍ͟��	���	Uy�uӀ�x�C�O��D�O���"e­/���f	�`M��V&+�����d�O&��=��k�|X:v苇B-��bU`�<a�I�ZT�QJJy:�c>��'0�����|z�M�`�`��)�����8��̟���[�O}��wm� q��
Ri9�/�:B�#b�V�!R��O���æ��?ͻG�@腯+��l�6
%��H��?����?���,�M#�O�N/���I �}�N�S�᙭O_��%��
6��ؑM>�-Of�$�Ox���O���O���u�D$TM�F戡BI�sկ�<�°iB��'n��'�Oj��ΙL�2�z��7-�&	;ҍ]�o����?����S�'W�t�2��]�/X�e��@U� pt�4�M�U��2�&3|�#�D�<��cՓ78���bEE�\[����O��?9���?��?ͧ��ZĦ�`Y͟���,� *���m\�JE�"�Čɟ �4��'x��?9��?y"�$�\�ã��_����٠�J�Z�4��$Υi��?��}Z��wGT�q�)R�q1��'��Nޡ͓�?���?���?����O�fU�ė�.q���d���Z���	��M����|z��E����|��
�=�ŀ�A�� �T����ճ[��'5������P*pC�֝��Bh�4q� 1;�d�bF�)��W�:uG�'Ff�$�p�����'��'$�4@�j�,EF]"�)��K�t	��'��Q�`��4h�����?�����	�-� �ZGd�Dӂ�����,]i�	�����O���2��?��b�{��i�>z!W��*���b�<c����!$?ͧ(y���B���W�V�yE葪QZ��g�	� M�\���?���?1�S�'����q��L�3 H�1�7�W}� ��I�1�I��x�4��'F\��?���Ȝ~����֩�rޖ��˄2�?���Xup�*ܴ��d�%Kq�q�����Sd%�R���� K!a2��{y��'B�'�B�'�BR>	�l�d}	j�!�,t©�a�^�M�pC���?���?qJ~���j2��wX�y�a�'PG\�*ExN�|)��'�|���@�[/��9O~AY#�\
���фՖjВ�t5O `� މ�?�9���<�'�?���:� $��Vm�E���R��?I��?���DC�Y��	��d����t��oC�>�x��+ϰ0 �	Sh�g��`�I�(�?AM;q$ERS���@X�1X%An~���}^z�L�%k�OR~	��$""fH=S����ac�p����A�!G��'2�'4�Sٟ��v���0U��Ɯ;���6�_ȟ�[ٴA:��+O�\oy�Ӽ�D�=XB��B�I����,�<q���?i�H�ݴ����v�34��P�A��E�9Q��'�X�����䓅��O<��O<���O��$��
�b%��Nu�׮T�UѨ�{F����'v�R�'����d�'ٌ)�CB8h�)���<lh�8����D�O��D-��锗|�����Df�"��+ò:p�� t���&��sB�Oĝ
H>i*O��` eV0na����#�u�ب����O��$�O��d�O�	�<%�i�E@��'r��#��I�D��h�ߒS�J���'ؚ6M!��)����O���O�j'""F��gR1X�T{��ӟ;Q�7�7?Y�՞I����Z�S��I�F��@UlU�ta��'���@i���	C8�m#���.��F�ʃ"��	������M{d�D�c�T�O�Q8F��"m�j�($�ے K��d�:���O��4��,Q$njӼ�Ӻ�De[.��xX��Ѯ3�� ΍�{Ò����`-��O���OD�E!L*|,~ѡ ��ah�����d����Oğ�������O=�-���݉,$�0P��	�(d�\k�O���'���'�ɧ�	�9M�4¶&�_�8���ϪZ����nϕ]]�����<�'6Ux��כ��b�9Y�S�0v�Ю^�\ ���%(���{6�bd�v(�h��@F�"Q.����'E��j�⟐��Ob�䙙���T�Y�������^�d�O`�Rg�.�|��E�?��'� ���ON� �~A`@d��D��@�'��IQ����v��(��S>f]�L��ؽ�M3�탓�?����?	��Ăn��nd�7)�	�"�_��Y26��П@��\�)��,��o��<� ��b_'!VDJ�Mõ�^��W8O�u0���~b�|�S���'Bb�kq-�d)l8��TcWF4j�B[��I��B�'N��)�6ic�@f*�@��@��O���'�b�'B�'˼�ȡ�����w���
��O�=H�Xva�6m�`��5��D�O�좒$�a���.�2\��M�d"O��!%bX	h�`*�[:i��YA��O*�m�	$|u��؟�(�4���y.	Ė�Y'�ȉ�X$! ��yB�'���'������i��I;	P2�ӟP!7�J(8n�mL!j�З��'`�	x�'0y��[���J�M.�
�OJ	oZ��4���̟���|�'m
���ޤI��@[)Hpb%+�P�L�IןH&�b>QX�ǥu(: Yc��4)M�2@���,�oZ ��ĕ2�Lh`�'A�' �I�QT����� ��;���UrX�Iʟ�	����i>є'�Z6M�%	��ȇ�j��g��)i�>�dn��]������-�?��_�|���������VfS�z��IېK�vt%��Ŧ��'A.�ڡ"��?������w�詢��ӚQ��r��G�=∋�'YB�'�'�B�'��l�դ�&0[�,(�I6�U9�O�O^��O�im�7���˟�P�4��_Qt��`�Ϲ"d��OBsa6(�M>���?�'l+���۴��������5]�l��۶:�������9�����䓺���O����O��D<u�@y"���b�MeU�Nm����O�˓}���i�:[r�'�Z>ISȔ2$n�c�@W�.����u/.?A�R� ���� '��'P>��2G�
,d�99��	�a�z��T�y�ƈ�A�����4���#�k�̒O�e�¬�0>00%��� 8[Z�#��O���O�$�O1�8ʓA�f���u�~P�P%�?mΔ�!
�tv��P��'T�ky�T�S�O,�D�zP4��PCX�j�p�U�@z:���O�Qq�o�R�ӺKR��3��Ué<&�U��v؁Q�ʑ�Qh��<�(O���O����OZ���O
˧9�8�qNE2r>���߹\���ѺiֶY��'�B�'u��ybLv��.�c����eC�?@�[�F�e����O2�O1� �Ab��8+�\X@!�6jn\q�oJ�,<*牀N�1���'�$�<�')"<O~�s���3π@x��(b̩3$�'Y��'�"T�(�ܴ/�"�����?q�`�E�u��p@���Pe_`:@N>��X�I���	G�1y��Җ�ܯ_6��W��@z�_��\�F�A!�M���t��B?���|��n>X����4d�\4t�;���?����?���h��ŧx�GH«F��1���G1$�H���⦉"�h�����	�M{O>��Ӽ{�m��ޢq���$0gj�Qk��<����?��"6	��4��d̙:9@�:�OOYb-Z6eR Ej%*�VfQ`f�|Z�������I�����ɟ���+Ǆ�jqGS�_h tR6aWry�l�b�H �O���OB�����)��
R��X� �b��1���'��'jɧ�OK��&�� ��:$��!^�Q	H�D��	�<���B0I���I@�	ey�Ƴ�DL�T�R	D�ĠB�ۦ7p��'g��'��O�剶�M�B��?�sd�%E[�Yj����d�R�x5c��?���i/ɧ�th�>I���?��c1f܈�����-��(0nڪ2[f �4����D��͠�'3������nZ6e%�u"0���`F��'@K$]��$�O�$�O��$�O���!�Ӆu��Y�HΠ�P��	�b���F�O����O�,mZ X[��ݟ���4��;��E`�$��Ir���Tk*�K>q���?ͧr�D���4���&A�( nL�o���1�O�GՄL"C��~b�|�Q��Iן��	Ο��R�Ȩ/�8Bk�l:��q�����	ky�t�v`�p��O^���O��'#8>��PC]'T��[���At����?��_�����P$��'	,����L�`Ә�4����u
�L^�B���J.O��V��~�|b�Dd�QcAH�K������Q�b�'���'���^��j۴!,��"��j�����Y-M��������?��&���dF{}2�'~�!�J@l12��g�~��5s��'�ҎM�	����p�tq�j��vzy�eb3���8�ąj�1O$˓�?���?	��?1����IJ1N�\��� �_��]]��
�i& �q�'��'S�qmzޕ�v`Аs>��C+_��d)2��X����X�)擟7���o�<"܂6��h�֊��'f.�ʡNO�<aS�j���	N��uy�O�����,2 *5j�>n��@z���"IB�'���'I���M��k_��?Q���?�S&�8��ybDN�6 y�P,��䓥?C\���	�$%�dSe�&N��$�Z�Vʥ�L$?9�I5 ha��4_��OB���?��p��\ĉ�D��!H;���?����?��h��5~���A+Q� �3�d�2��]ڦ9���ş,�	��McO>���p�:Dp4!��۰k.K��C�<���?	�5��E�4�����K�~ �$ݣEИ!QS��/aALT�r���������OF�D�O��d�O��$�(i����5�h�	��	+�r˓1!�F��UK��'�"��$�'�L�e�Q�+����rE�Tc�`���>����?	K>�|Bg��j�? "��׭�
ǈ�Qʑ�j�ε�֮}ӂ��'�TT�W��u?aO>�/On�C�ΐ��E���&�X��� �O����O����O�	�<AĴim��R0�'g�����)'G�!e���:�:�i��'0^6�(�4����'��'e���1Y��3)Ts�:��cR>K��0�C�i����I�,} ��OJ�l'?5��9"�&���ӏh�P��FՔ&��Iٟ\�I������4��_�'w�Ka���!�!��2ľR/O:�Ʀ��7�p>��	��MK>�J�Z&��nG�Jm;� ���?9��|:g&5�M�O��$B�˕���ֵ ��
�F�F����O��yJ>�*O��D�O��d�OFU�r�ٗ8�p�����t�8��a*�O����<y��iQ<x1��'��'�Ӫ�*xӅ���)�*� � �2.�I��<��O��d�O��O��(a�p��`��"ii�A
����O�܍vW�D���o���4�D ��'��'1��IB��
�T9��?i���c�'V�'u����O7��M��K�
\�%9 +[�B�t�U䞤p6F�����?�w�i��'�Ȣ>	�h��{"&PtR���@W:�B]����?��$�%�MK�O��	ֆ_����S����4G0��ذ#�&W��3�
b�T�'���'���'q2�'��өf���ʑ� ��`�&����4#/�T*O\��4�i�O�4mz��$/Tl�r��]�v�P �៰��o�)�"���n��<��/���t���J�� v��<���үD�$��������Ov����Alj�p%	$80��9E�U7a�����O<�$�O��3�f�C����'nR�[�'��K���6�����.��O���'G��'��';z%��+�=I��`q���%l\�q�O��� �W�An�7M�\�*\��D�O�)��ꓵ?�@|��a�g�$����O����O��d�O:�}Z����x��+u�`��D��⡙�6����T��'�7m �iީ��KS�O�48����4�8(j@Ep����㟸��;S��m�A~�&�&�@��("�s(M�r�� �gL�, �2}�H>�/O2�$�Ox��O2�d�O�ຠˏ�045��I�6g����"�<Iv�i��<cu�'3"�'���y���� ?|���DE"Cd���?����S�'k��au �o[�M����<?R�]�l�1�M�rY�����
�[rvM���΁�Si�v�e�Փ0}h8�$(�H<)QG��t�`�X��!t�i<Q�Byg�Y �-�|kҜh�A[1Ԭ8`�eY�mBc�)bS��!��"�h�x`7�	M���&Wΰ�ɣ"ƉM:������(ArڑH��Y�F����:W������B���1��F�P3�����wD��G�m��4�v�$k�8	�w��v�D P� D�Xͤ����,h$ ��C�>S!�T6#��fJ�$�4E9���4�����L�WھHR��:���'T�9�<��GVq4b�0�aZC$�6��<�����?���!�ڀc��Y��R�
��@脬����M��<��_������ ��m~��
?*��쟬i�AżTbla��,�5�,��C2�M������?����U�{R�� �
�c�X�3�������MK���?��O$@+���~����?!�'Q��!eD�p�Q� ,��CX��	Ğx��'���*`;b�|"؟LY���B8�M�V�Àv�P=�u�i��	�<n`n���h�I៤�ӿ����ܵ ��� ���c�n�< :d�9!�ie�'�
ۍ��!�ӕ%0���H�x�±:t&�h�l��#?�6��O���O �i�Q}bV�x��V�zY�Y:4��2bj���-׾�M�� #��'v��dI=~�|x��f�J�TlyV	�xuL�m�؟��ʟ@�P�����D�<����~rU*q��D�U�+�Jez7��0�M�O>ك��e��O\��'��Jܓ6.�A5(Ox�����:S��7��Of��}}Z���	}�i�Ak���<s�rp2��Z�N�|��a�>S�LL��?a���?)�O.��U�̅�A
G�W�&���j�� \������O|�OR���Oz� �9$4�	���h��s�+C�;pL�O����O��d#?��$W<��4u�(қ*zh	[�ͱ^��}�q�i%�x&�P��\*k�>aE�W1}�`]З�I����i}�'"��'����Ox���O�򫘴a<
!��G�%V+*�s��*7��O��O����O�0�P�%�	 N��(�&�ҟA"��H�4�:6��O��(?aP������O���l���j�k�THx�,��mcz51�o�	ğ��I�5�0��?�O֖��J�)�l�?!¸qݴ��d)	 �6��Ob�$�Ot�	�P}Zc��d9�ʋ�olz��K�15D��4�?����	�b�i� 2�z�H�d�&%�Z`�#$��'�H���'p��'��m�>�+O�$sG��XU���#���F��Ȧ=��Wj����O���F�fy�"�dW\���"'���#��6��O����O�$�d$K]�?�D��l�3e4Ҍ���j0p���Gm����&�D�Z��'l�'D�	:���DF�I#��CV��9�6�O$iYX�?�9�d�:;��9��#����,�*�$����~yb�'%��'��ӞA�=9�O��}K��\�_��KÔx"�'���|2Z��ݰL��i�k�n(-[ES�bk(6��O6��?Q���?�̟^�#6�b>=Ѐh̔+bQ�1hP�.-��ծ�>I���?qI>A)O�i�OJ�a�f��%2tː�����'��'f�V�|���A<�ħ� R՘@)�	y�`R�]#-sP�iS_�l��gy�O�r�~�逜z��4���̞	�������]��ҟ��'&�i��..�I�O�����q�I���hIr��;3ތs��x�P�����x$?�i�I� ,��O���H`B�L�\�S5�rӂ��a�вiG(�'�?!�'|.�Iڑ2���08`z����6ͯ<����?�֕�4��ܴ`�Q���-X,�qcݻp�>um�k��i��֟��I�(��Fyʟ�QJ���ELNY+"�D%�U��U}�%���O>ig�R�@"A���1>������E��Mk��?y�O��� *O��w����>~v�� �+4] p��>U�DDxR�"���d��Rl��(FH� ���@" �:Ȧ�o����CE�@y�L�~
�b�Ǿt@�(ɗ�9}2Ś�ps�Oz� ����	���	q���L�<ʚ`�� �^�u�%ʓy�V���x�'�"�|[��]3��Q�@���CF	���7��O:�O����<�
�\��O~��Y�)Y���Qփ���H��4�?9���'P��;H`ӪĲR/�#?�F�{�
�)�ظ��xr�'P��՟x�fo�S���'@�Ś3�ț��	b6e^���Moӄ�|��Py�����ēr^4숔ŔK����d&`�n�՟З'b�/�ޟ��	�?טm	�h"Po,ڠ���f��O��ĥ<�7��~��uw��(>yu�vk��aY�MyW�E>����Ob ��OZ��O���*�ӺSBLC�c�R1Y��/=�� 
�m�	jy¯Q/�O�Oj��p Yi���Q����7��!#�4.� +�i 2�'�"�O-�O�iNC��J�@���PAY�M�L7�OZ��OʒO�s�h��6k36�
�Yai�E��,�׉�Ɵ��Iڟ��ɒc�Z�{K<����&�X���̑��HⓍ�abĠm��<&�8A���$�O>��OZ�p���dA+2���mx�(S즕���r	�Q�K<��\�'�b��� ��$�矹)� �ÇrO|���<���?�����D��zݴ�i��(�*�B��Cp�D��M�]}�Q���ILy��'Y��'�j=� �ТF�V�Pp�#T�X��4�R�y�_�h�����Iy�.]�Kk.�S�g�6�#�Jݖs֐!(�E6-�R6��<�����O^���O�!�r3Ohm�Lٌ�M�f� � MP!O�ۦ-���P��򟬗'̹x3�~��3��=1���b	#� ��Lۦ��	PyR�'db�'MD�8�'���Ƙ�1̞8���@�C;N���m�П���Vy���o��맩?����c�,�Ҍ�oʩY�H=��C.w������I՟���p�X�'�ޟ�dY��WT���`T*W����iJ�I�g�P���4�?	���?I�'O��i�E@�F��LyiUm �l�E;�l�����OP���?O���<���TjDb<6!�\�� Ѝ�`_�V�ߓ/46m�O�$�O��ZF}BP��A$�-�*z�(��m�d�I���MC���<I�����6�ן�pE҈[����nw�I�ӭ��M���?)�]��E_���'�2�O���� 82��6O�&g=�Yd�i>W�
%q��'�?���?�b��8%���!��� 
P(� ;��'�ްXRM�>A*O��ĸ<I��K)��p|0�'kH/YҦ�g�c}��I?�yb�'Z�'�2�'W�I,a��Z�E�rX`s
Տb� ���"T�/��	Yy"�'L�Iٟ��̟�1)�.wH�|h��J�O�0j���4���?����?!�����y��ͧV{�bCU�$�A"bC�!K���m�ry"�'��������j4�t�0;���${B6U�"
;0;l��#�:�M���?���?Q/OZ�x���X�$��5�/
d�J���(ɼaC�dZ�M�����$�O���OJ�S�1O��D���teE>7�θ��gc2�D'g���d�O�˓zL���R?a��؟��ӑ�\0�G�.5�L��b�Ѡ :~Y��Ot�$�O�����|Γ���CR�  �r$�(5�@�:7�N	�M�.OD|������	������?5:�O�n�~Ͼ9Y��ŭ+h����l*���'�B�մ�y"Q���	UܧK��;֊��qt$�i��3#�(l�L�X)J�4�?���?��'9���My2������ä�D#�Рs�OX5wh�6mH�����O�˓��OQ"H�i��i����CҲ�
� ��D1t6M�O�d�O�u��(YN}�P����v?	�iđ춑	 !8��a�H���vy����yʟ����O��Dđ�@�!r��3�C�D�Rx��lZ蟸ʇ@
���<y������Ok,	X 0%H����P��2��]�W/���'���`�'���'�B�'��Z���#ɕ�Uk����4F�{#̕:�^YC�}��'��'���'ښ ɖ�F��������xF�Qr�ျm��X��	˟(��by�R����q���(s�ϐT3�U "ݘO��$&���O��D��OY�Z�#ӊ��n
7��49�.��]�'��'��^�L�s�R&�ħ`Ǆ܀�,�$^WP��A�:%��! �i1Қ|R�'0B˦Z?r�>a���6y&�����%���IFbͦ�I��P�'�p��*�I�O����La�CY�8�b�H��I&�X���ȓ��c��%����/��u������m C��);�uoZwyRH�Dz7mYw���'����7?� L!�ւ��	"l�{'�3E���s�i�"�',��'��'�q��0X�`?
���yvd? 81d�i���7��.�$�O���V��>a�  �1Pz�᐀��N�"lb���:������y��|"�i�O�@�FD)}H.l�5��'��a��ߦ���ş��	�M|���K<����?��'��	'�(a�-*���?����4��U��[U����'�r�'r�u1%/ˌQ5Qj�l�5I��5{�m�����?llh�%���	���$�֘�zĄZ��ŉO�ʐ��I6 ��EO������O����O>�IґU� j���FT�q�|y�]�-V�O�D)�D�O��J;r�K§��{:�,!�-	�YP�!���O@��O˓H��lhP1��5x�ӫD�\�Р��\d��HP_�,��V�'Z�	ӟD���8UÀ	2�Ş7�-3���&����O`���O4�-%⤘Ė�N��[
�VA� r4��iC+G�b��6M#ړ����O��'��h�V��;�x0"`�(E�,cߴ�?����?�5u�����?�(O��I4f%�a�F��v�����M \'�d�I~y����O�.�8	����I%�ݸD��{6Q����Ȇ��Mk'\?}�I�?i��O�ub�	��R��,���4Ƴ��'���p��D៉'�����I'�`�c&��@|��ݴS��<����?Q(ON���<q(O���)��-jĐG,�	jH�צe}r�Y��O1���$��3�0� �@J' ظ�@�,�k��%n��L��������ē�?���~����*Cfѩ`�����&@���'����yr�'���'�n�H�ߞ<�@Ƌ�,��HGbӰ�dR(W|'�h����P%��X�\����A�.DiF�
�dR� �	�<����?�����	T�fؚ�@���
V�K;Dz����mYm��?�N>���?�dQ|�q�&&S7��A� mހ9v��<���?��� �6�ͧ?��j�'7�8a�o�5ǌ�'���	x�֟������'�ؕ�R�H�J4����n�;\�pM�'�'/�[�X	���%�ħv��P@Т��4΁2$ƞ0�,]�r�ii��|�'h�L٫��'��e�4)�BfN����w����4�?A����dE$(��t&>����?%���e���c+K�~��0��B����?i��h��Fx���҃� oG�" ��.#�v�*rZ�|��e�t��Iٟ��������ݟ��'>�8��A�oϖ\�uH݋G~@nZǟl�'��Í��t�]�#L�	�@��LE�`p��[�M��@3��&�'b�'���2��O����6В�9���@@:JT\؟���m�la�U����3)�<g� ۴�?a��?�eH�]c�O��d���aY�@s2T��hγm�؁�+lO`���O��²v�z��i�|�Ah�F�$$�(mZΟ��'�ς���?�������"~=��+s� �*V�UhĄMW}����'���'G�I۟��UK�+Qz���� )c
��S��^�f��I蟼���� �Ik����$��T��� f��> �m���Y�Z���oZ�k;���?���?�+O�XjG�|�2�կ�Z��d�#�"��W@�f}��'q"�|��'pb��$�3#�H#�	�98�=���\X��Iޟ\�IߟĖ'T��1�� �i�FHP���N�:�� �kN��,nZџ�%�\�	џ�!Q�:����#����Y��)ò�U�NI�6m�O���<١�x���(���?!X��N�v*�8ҩC1@(`��f۽��D�O��d�O���5OL�ĸ<��O�.���@�8�|�pc�Ъ[�n�[ڴ���*��nZ��������������Ԡ��#7�ҐG2��U�7�i�b�'MPh�'��]�d�}:��!:*֕y"f.3��y�ϙǦ��e�M����?y���UV���'�H6)\�7��F@˺BI�Bcw�^���1O ��<�����'�½� �
)����K@�fmtӠ�D�O���D�L�\��')�џ��~��(��7l�Ti�Va�<n�ן��'�j�"�����O����O�(�3E��2�k!�I#�<���ަm�I,wF�ҩO8��?9-O:��ƪm��%=\e3q�A�Xq�V��#0�~���'Z�[�G�(�J��J?�ء����D�����/��Pǭ>D�D��A�Z����6DpޅI6�2��h��@H;5(~A#�'��l	#�K�
%�xQ���0�`�����\�C(M������h5r�A@*� 	��1sg� "��1!��2�z�1�^.I\�;!��<I��Q�*�1b]l2%CӲNr}3��Y�
m��D�#+����c+y�p�p��,V4��S����{���£�7_�l���C�(2�����8�	� Z�B¸4q����Ȫo���+�
Q::-�i�+,��x0�,W��|�f��r�Q��XTLA0�h��P4a�0�o��)����S���5{��0�*�j�L�2PV�"fʪ�?����O:Y{��X;L<��v�e��j�'��B�Y�"8�u�4�V�d�q�혰�0>!3�x�BZ �@�yedF�\���KӦ���y�h�zGf든?+�L{���O����O:lqv��^p�W푘?eZ `���PC���.�i����`�۟�'���?y�F�}�t�YF����`Aw���G=ځ����RBX�s�,DC������ 
�CG�PT4�@��|I��Pѩ��uH���O��S��Q�s�H}S����?�T5p��,8C�ɳ�l�a!��!R�x�,{�Q��J���?��Ԫܯz<P|��&X5���Rv�����"uF��3�������	�u��'����#L�ر5(Z�W��[0NY �~�!�0u��<:�)�A������^M��O;W�R�F��d�R)��ƚ��LI�㉕�P���������À�ϸ�I�d��d�O\�=A)OvI*��P�?��g@�i�Xi�"O��[��ɧ	N��6E�1{.�@�(�E���ɷ<��O�+h�Ś�uڄa��L ���q��T�+@��'F��'����'�b2�PP�gfG�;?`y-A#S��Eu��
x����(�Є{&2<O��!
��8�;���&�A� l�Nx]S�ַn�^�`��3<OvQS�'��U?lk�h�7/
z	,6'b ��=���d�!��qw&"|�L1a
��`!�D�.oD��`.V߲�iV*��88�t}\�Pb������Od�'����P�}�\t��-�A�$v�*���O@��'P���l߶5b�i��Y��'m>@@ҷ���DNdb���`��uDy��Q�YQ���ԁh9x!���'vp��D���<mX3��Z�QDyҁ�?	���OK�u#0\������IV�ت�'0�R���<�"2��4.{�qE�R1�0>!��x�AߘW%��0/F�ؙt�9�y�����`7��O��$�|JHW�?���?�2�U�X�H	j�o��NใW�E�#���������	��X���b�8Z��̱�ؒ [jq���a����"m0�$j���0$��ؕ�U��� ��'1O?��Q��| A���L[�ī �!��E�FV�sUL��&�Ό�G�F�\�� S���?PE"G8m8 �	�����BQԟ4��&!��@0�ڟ$�Iß(��3�u7��y�� �X�ǂ�h���3���~B$_&��>���8D�l�MծcH��OUU?��Ix��{`�PԊ�\X%�`�Zߤ�ɡT���8|O8����^���1�]E�8���"OLmy�K̉`S��WB�NmH"i�����х���͑&�Ռ�Dpdh�?d���Y��ܟ��Iן��I�m~����؟�̧G���	ޟ��6�̀S��"���,uڜ �=�O>h0P��c�)�47/�-hP�C�G<�+	<�O��'�'����=4��T�ۜ{��P$��3�y���:��A7�-����ӏ�,�yR ��GF(�y�M�Z���U�y�k=��)��R۴�?������!qHJ9U���M��#�X�~٨���O����O���Fh�O^c��'F�BE��3i=�����Ƚq�L8GyR+�(��d�"���o�l�G�?{8b,x �	�"l�$/ڧ5�,��ɅP�ht��Z%��ȓ4VqIAk�h� ]�Љ܁T��l��	:�ēyH��3�^�Ha��c������s��1��iG��'��S�h/���̟L���(�L���ߨI(�5B����'��X� J�柈�<��OV	��	�cy�88���j�ICdU��V"<E��V�9� �ۮH��=SE�k��ِ��?ٌy���'άXą�;t�#6�,ҪTX�'�p��!�۽	/+�؞w�R��U�*�`L���w�<�s�G�55�=��\$"vM���?�4$��\+&D����?���?	���|�4���iΥP3D�J +Yjjb��O�9�b�'�~EҒ.ҹ���Y	ڈUL��
�'����X���S�.rt"���&���P��{������2t�� ���0$�E�Æ1D�p �ݏG3*IBӉK)[�Pv����HO>�Ӫ���M;��Qr-�Ȁ-088��m�>�?����?Q�u�����?	�Ob������?f�4l�&�	��B��q�W�B8�|j�g�<�q"�<OVhi0�g��D`��r8��Z��Oj��U�=���,����`0^�T�O���OX��'T�V�I�ˍm
�)��" {B��ȓ@������/�̅���Ѿ�x�C#�Ihyrn'l�D7��O���|�T�ˣhu�Ű#!��uc��M�3�R=���?�N�$��혧�˔b��8H@��<h��@��-Y�W�Q���	'�'Zv��$	y����.:>v�GyR��8�?Ɍ�� ���c�ʶ:���pԣ!OG�( �"O�\�Sǘ4�x��K:k1Nca�'�,O&�p1�))�8P$�` 3#"O$8`�
e	�d��K��@�`�"OL%zr�4Ǝ�g+Z��a""O5S ^����3�J�&w�v�q�"O�X�%�c5����@�IƼ"�"Odm�B!;��0	dc�2���"O���c��i���K����LPw"O�$���Z��~�1��Q�Zl�1kF"O20	�@�"}f P��٬qY�M˲*O�T��MΖBE�h����(Tx��'���c0A!�~�˶I�3�:z�'�j=X�-�hk�ݰ��O���0�'B�;@��?"Xpy�b� p���
�'��\��)M�*~�u�U��@�'"�MI �G<3$���TB��.9��'�F,xe+=Q.�8)�@�Hd�	B	�'�ة� �	7G��Ԉ��)@�Tx�'� pZ��ӎ)��<�7 �0n�ɳ�'�h�P��X�q�.��� Yf�p��'��=����]|���jإ{CpK�'����"�6D��P�W/��nѼ�	�'9����$W5��J�CO���'���@�F2?�d�YqFN�3�����'E�����*\��1��i�*3 UX�'�z XY/F:�ks�Оv+���'�Ψk����i�y ,G�o�д�
�'s$� m@�^��T���]�f=b�3�'�6���&ǂ4����(�dK̑�'}�
PJ\��1�XX�-��'~��35L�"����Tb�%NΨQ�'��Eɑ��L��	h�EE��*�'�	�Պ�>!�bt���8G,�=(�'�<�֋վ,"��"���6I�' :p���-[۠x��Ԡ� ��'zX\i�'TFCT����i�	�'�B�	�DӮ{� ��� E{���k�'s�%:Sϗ
M��9�i�;d)�1�'a|�1e]�:r�K���j��݊
�'F��p2OzzS�Lٹct����'���FG/@�<b�D�?[S�u��'����4�*\���b%J��K�µ2�'�\	�%	ڿf;䐂䧘�+ �p,O����
�]��ܒ�d��[B.� }�P�b`.�O@�"��xr��1tZ�%�.�w��K��-D��fbS��$�`�@_���@�,��<��bRg�O9�@�`���ք8+ԅ.�ԭC
�'�ԁi�/b��a��fM( qQO��2p`����O�q��9s&H��<��s"Op���C�!7`(�G��'��\���O���C�,<
�{R-4,Cn9@L�=8$x;�&��p>�`�A�L�u�	�4p9P�c��>L��M�?X-�C�	�I@4Z�']�0qW ۉ}�"�<�W+�MHF��dۥ_2��`�ѝ)��Qs���"�y��0r� �D�Q"۫�J�;4H�)��'H$F1O?����g��p7+߭o�\`1Q��c!��U59zJ�*'��5�2�)��P"U�~���Ó@����I ot��(���������\4s)���]6w!�$���8���V�z���Q�ى>>.�>�ci���H���X�nؕR��܊T�,^�:�y��I�3���4nٗ�(�V��ǇM�iI:ŀ��\�O�681�O�mR)'�)ڧ}�t�����;:�,�s H�XL�D�K��M�L��##�`���OvrA`�|N��3&�9T�i�C�>agM&��=� �5˔�,���E�ȅ�"�i��O�E� �.vM>D���dLR�7��
^���� �+��"U�&X��|U��pɺ1�u���`�b�f� �>�4�G}�K_L�>�B�K�Y^��e�:1�e��b*ʓ}"� �J�]V"|J�g�"-�	�(�	w4�PeIV}�L��O�>�0���Ϊ1x��0��@w�*�q`��3�.ҧ��«�=\�x�
�_P4���N���y"B5eb��@i��G�P��uO�����	N#�zbl�����/b����f,�%v����+D�(�ղN�p��oK���a� (D���0��7����o�-E�6�:�&&D�X����k1n$hfh9+�@pÈ$D�A�
�>=�����!�yg�j�5D��H#�щXq�Á̵j�TM�Bg2D�PC! k�$��&,T-3��<D��BD׬>6���`$�LL�A<D�|�6��2{�҈^�.�kԮ,D�$�$�1Rh@�D�pa
�� �(D��O�'e�M��րN��ԧ'D��(��)�f��G�W��"�,'D�XCD]�"�L- �F
	�l�� D$D�x���+N�4A��/�z���b$D��h�e�l��L8��N�qo`�!�� D�D�W��=�vHے�pk��W#D���Pb�	]ޝ+�NQ�_h��`C-D�LKfT)[(A��!M<Wr�2�&-D�Ę� X0F��M�n��S��G%D���$.�L�2E�𠜍*"�bE�"D�x�)Y�nt2���2|� �c;D�<�"%X( ��՗��C�ɠ+��H��[&~ZP͂�鋑J�C䉨J���0o0�Poާ
��C�ɻAX!�s�C�yo��ӳ��o`�C�	+6����Gl�\t�`e�7��B�I�c��=�D�ׯ l��A�,�B�ɶR�!����X���p�탺U�B�I�b�* ��� �j.p�0���N�zB�#T�x�o�#���tH�Q�B�	:i Dpف�A�Wۊ�!��@P"BB�	7G��r��r�Z-:�F�=-��C䉱	E�HER�VLp(Rv�C��!!T��$摼E٫��O�C��?2=8yw%��4������+��C䉓i#@`8���yZ�c<o�B�I�l�J�r�hʠ1�Z-�f�6=��C�	0A��9ʶ'"j�:�!QO�C� r~]AC�Q;E����k�8�C�ɴ?�$`��N�P���&N�v�fC�I?��A�ʚj�T�!�O>��C�	j�������Ud�ũ2�����G�ɉWmv:��|r�dɅ�S�w%��kJ�4�Px��
R��$�E�g�9�J�d����ED�N��	�1��1c�*�,\ъA��\��č78_�<��ME)����C`r���l�P!W�E���V"O<$q�J�ho���ꎖ`��ԁ��>����)�j��G,�@��E�G)e���i�i�м�5���S���~��!A铁E����A)�wlR��RO��.�'�Ȅ2��X���]uJ"�1-#p�3�P;G�mّ.C�Px��5� �YZ��!M���b3g�y��,4J�O�����b�#|� �Y�f�Д�ė�� ϐ(\�}����j�� y<�F@dN��3j��l��,�5F��M�"~n�2"����m�+>� ��2�[=2�C��1~���d��>6t� ����S]�ђ6��5X�>��DL�I?��i���`�Lt�f�>A�a}"՚B܈J6�?� �5����|,J!P���c�hA�h%4�ī��G?}��p��}=��I�d3�F[b�"p���^�t�?�hbC�0��(��+0�����+D��bN�>q	H�b�
°Y�#~�Bۡ"�>^�K�"~n���l�Pk�	4�T���:��C䉢$j�= �N�����H��J��6ʴ��V!��&������2��(V,?D��sIZR�a}�늄zl2�cЏO�G��8%MLbL9egR�D.�Ą�#�V!"* <_�DY��F!n��GzB��!c1R�_��E�^�9���.k��8���E@�X�ȓ\ \(��6
��a��P�E�(�l�;%����@�Hlp�S��M;.&;� ��H·]�pA`�F�<i��W7Qh��*`F�$-!���0�\yB��)=4�K�'`��B��*�]��d3w��
�'Z��  ��%r2�H��.l�xI
�'8"�5�Úa�A���b��Y�	�'Fi� `��N~��w��Q��Z�'Z�{�mG۸A�G+�0O�>�Z�'�J��1��>;鼭Ɇ��5�:���';R��
��%����[І���'��5�7��;X� �+��I+(�V���'���i� .]tT3���,$�t�'��@�h��w�*iB���ը5��'f04 �>;�VDz�n	�T��'S�5#�c�7K	�`*�ƾARȴ!�'o�˧�5|��wBĉ)c� ��'f.��u��k=��7�JS����'NDM9цD�6�B���ℳ}��9CדTf��xa�>A ͂�z{v1hb�6"��@��S�<��D�-Sغ�kr��/?�|D�U&Lܓm62�j�'������ʭJ���Y&e� �F���"OP���"�(�oF_�d  �<:�qO"�I��Y�Dゃ�BV-����oi�ó	+D����'���"C ֶr��8@\`	-�O~���޳�p���Ӂ@hL͒��'��Yz�,?��ضɘ�[�F͕P��,Q#�N�<!�EA7*��c'�M��18g@H�<I6���_��5h�m�ds����V@�<yeh�0t�P:P)@1����W&�}�<1�'!APֵa0)�Ph�r�`�@�<�G��x)Y�Ң�r	��*�+S�<��ش@PՁT�B�V��3��K�<I�˒7bj���3:�.�;נ
l�<�G�K�!�½ӳ�/-W0<0��g�<yS�� boX�".�(QI����#Z�<�����ghM�B�*{'o<T������Đ���"^�,��;D�tW!��?"a�/�n�h��w,D�8!���Y�TbA���jtK@',D� �UL�nW��PK�B"�T��.)D�l�`�ׁ�8�W��M�vd���)D��bP'�1B��0�3�G>F���e�9D�,r�n����ٓ�R��F���-D�pe�6�@�B�r�y�d�*D�4��D�j!���Ύn��#J*D��g��>\M{�&TV� 6D�ة%/�
-z���K;U���CRD2D���ۡU̪�AT�˴k��I��.D����E�5+'5X��ȩQ��5�7�(D���Vjֹ0�1�B�ƪv� u��"D�|y�T����z�¾Y ��4�5D�H�G	��A�2�O��&��L2s &D�\y֍�s��%���#s� �@b� D��H�j��Y@f��S��RE�s�?D�� &M�Հ]�AP�Ո-����r�"O��c�e��E��(��	=I�҉X"O
�1q�V�%fH���7I<�t"O(]��H�!^䑒�%s�J��c"Oz��ǐ�<�5�֤S��R�"O�����F+I�L����_�{�xpe"O��Y��3v�1��$E�B���"O�1���P�~=���t7B��"O�cb,ԌB�f�0snȕi��1Z�"O@M�Yw�Ii��y�I��Pa�<�cǁ�z
�����%0����s�<�CK�3z�"z�Ύ� Ԥ�Gg�X�<icEǯ6�@Ga�'�0�0�JV�<�$�Q�(�"�q0�C�P�(��Ł�T�<y7IJ2ѐ���I!�����K�<!��	��|�!k� ꞡ!E\�<�um��!,[�Z�**�� �[�<�G)۠v~���Э>T\���d �b�<�5NȊd �A�O��z�B�"FE�<��l�����5!(�C�.v�<ɣE"���j�S8�C��Ko�<6��_y����e�2��D1�/�g�<9�#F.6Q�'��0e�"�ؠ��d�<A$��	����E,T͢�"�fJx�<�3H3{	��b��ϫg��qVƉX�<q#����䅹M�+\�NDk��PL�<��C{��ts�u����\�<�����ms��s�LMw���YS� V�<)��ًv����"I��p���G]�<� N!-Ų��!�PҘ��p��[�<9��T+Fvd(vc�l�^8�!q�<��T x>>�郯��2��0���i�<AH��D_��u+
I��	�v�Ti�<��ܢ&U |�ՠ��|n4�R� b�<ن��6[�d�Q��Iw�r-�c �s�<�w蚏o�\�X�V!��0�7j�m�<Y�i�O��)�у�R�R���g�<I�Ɲ�G�p�a�	+���!D�g�<�rm��`��y�/Ȃ+�@���kx�D�'I �!+�}|��ƙ��4��'��ݩ�T;j�tCB��*;p�I�'�X��@&}��P����41Ķ]��'� D���&y��z�/��_�pH��'@��bv�E�����HV���'���/� ������X�,�Ш �'Y�с�_%4h��� k�/�H��'�
�P���Pt$�p��M�F<�-��'B�$�`�\�Bݫ�ď�0!����'r�b��b �%���;#] A	�'�v(8m�;>�zT���%�t`�'��lskܧ6T޽T����'��F�,?�8]��̈
J��{�'����e;�F�82 D�{܂р�'*Z��� g�$y�q�u�Pd��'�ɑs�����b�ūv��'������Ø_�t,�c�G����'J-�P��i�����0@��r"O��K�e>/���p���<l���Q"OT�0��%oa�w�4k�h�"O ���BL"�l�� f ��sc"O�Q��D�h03�A�c���"O@� R�9=��=����60\���?c��@�H�:W��9]�.��ԖOQ!�Ć�He�P ��O��m�"eO$N�Q�@[��� �0B�P&���ץ�P%"O&��I�)��q($�B�9��y�O�Dz��)N�R�T��V�[25^4�P_�D[!�DF*���s�H�"�PQ�eQ�@1�|r��OD,����͉{�T�Pd�yb��36v
a�6�o�a��	��yңT+nҥ�P.��&���y�b�-T+t����N���X��ϝ�yBH%o\0�QƏ_�f9��
�y��W� �܉ZU�^:t�`�pFdT�yRdT��	A$D�W �Y�ш�y���� �	�U0ag��&�y�ܑE�*�HvbG�F�9�F%J��y��9GӼ��LG�N����3�R%�y��L"##�Dq��B����y�b�s��lSC-��s$E)�y����@���[qQ,x:��	�l$
C�	 �:�%�V7$<��c�8_��C�ɋu��(��-�)]� �u�D�\c�C��&[>��S��� �D�C#s�pC�I�qG�a�Ciʤ���?�DC䉸=p���gn�36���h�o�7=�C�ɤl����CW7
r���Ɂ��B�	<9[��"���TD�L�d�8D�B�75�l�q`L�\�� �"V��C��G�xK�O��d�<AVW��OƢ=�}
��Ŋh� ��ԆY
*+Z�*�FS�<�ƀK �N��Be��:���a�|�<�2B&�i)��F��:�/z�<I�&�kپ����N{8��g&�t�<A�f�\J�I[��V~�5Àu�<�U)F�+�~Hz��\����ggXl�<�����e���C�ͻ���s�<�$�;	���`A�ag��a�l�<���9��$�4��9L�\�9V��k�<)�b��Rծ�S������[�
f�<��v���s�cv������a�<i�ϛ��h����� `
�j��v�<)c���z˴l�5�,�1���p�<	�KHk"�BAf�Q&8�C[G�<��m;c���YUK�}��p����A�<Y��!Eu���#
�0�����C�<�7#����,�]�N]*w�YR�<	 l�2($�ڇÝ�k���b%WK�<)��5�bDk	M?a@�� d�G�<Q�)ձP
��s��L�H*��`O@�<	��I�u}<��׃B�Ҥ�P��y�<�k��p�4�;��bin)��u�<	2�÷>�h����i �8A%t�<�iJ�h$%���rMn� aa�X�<Q���Q�B!g�ةs2u�0�FU�<�Ҋ��8�h$p�����*$l�T�<�L$Pv=r�M�q�g�<Y�]�0Ҋ|��K��^��D��f�<q��7�D�,Y���@ۧ�_�<�Y�P���0���`�B+5��Q�<��L��*�eY�޲���΅r�<��Nۋg�x���N��P�%A�q�<�A�B<fmjw�ҏ?��§MEq�<)�B$k5S6EUxі��ǂ�o�<��b�0��x����L�Z�Zt��P�<�����u���޿W�l0g��T�<�#A�e���2��;|�A�6e�k�<�f٠��(���S9٠@�*_Q�<� �cC�Sh,<J�O���g"O���ˉ��(���C�ح��"O L!�R�C��!r�3.����"O*����Tc@3GLM�H��zd"O�j �V�Q�d��j�E��H��"O���5�X�`��Y�iI��$�1"O.�Q��@�l(m��'X�E��$��"OD%��G�,%�hl�% �pж�A�"O4J�O�\�(�'��.���B�"O���/j�p�9�-Ԯrt�P0�"O�%�@11&cٮ;c���"OJAS4���^(��e��I��  "O�H��j�,l������4 ��*�"OZ$ZQ�:j(�S��W����{2O������D�٥ė��A*���T�!�
�A�pɣs��X�F�25�)�!���e����/�>��E(>�!���-l����PqTGѿ2�1O@�=�|� �׌CS��Ҕ��+MW��G�i�<q��4y����e��MN��� ��d�<I�P9Kwd:��Ѧo�	�y��)=J��Ӈ�)3fE��A#�y� �	ɖ%SE��0c ���'A+�y���b���Rh��,��b����y�+�G��HQ)	:,�n1#�/���~r�'��q�Q�.�Q�r$E/�*��''Z�#��E�!�� Ҍ��IĹ�'�:��֬ӷ0V�xvN�m��z�'i�
ro�2u Xf�Qc��	�	�'���w@��&���	_G4��'�d��Q� "N@4*֊�)R(0�[�'�:}(�Ϝ)/fȃ��S�B�����'�L��M�;��D��O�0oI���'��J���h�2�8��v	�d�'^��i��ytB�򥂽C	�=#
�'= �څ�T����A%�F��A�'���e"\�T�F�B��=��'��,P���02�^)�`��ib��h�'I~�r$"�y�V]�W
e�����'g>a���	;w��+'�:g�d\�'o��QG޹j	�TX��BI<v���'kht�q��EL�ع��Т����'a9e,��/[�Ї�߼[�e��'KfL`7��eE:T��	�(qLj�'�.�:��;�.0@���B���'3�b@֠>հ�N"8I��
�';<cw`ҫ��������;쮼��'^2Q[�F S��Q0H����'�Qcs�(��ʧ��O�e��'0�2�>�%"X�o휥P`ěn�<���#Q��5a���5*�<)�rF�<�S�@�]�T��#�"N�L�`��H�<�"��#2m�`�Y�Z{��g��]�<5��G���JĦ��L�'�E�<��m5Ξ���鍏m(�Ij�h�j�<	3-]8.@��2���O�X���d�<a��'7�){	����0b�a�<yT�R�~v�0�� ťR�x���Sa�<��!�2,��@�QPbV͑䢚\�<QoU�;p��3@�Ù)�"�!��O_�<��B��\���P�M��#?����`�<�)N" �m�7���v���U�<��l�xxt�%�͒RTV�2��L�<ه*��h�[��Íg
zyЀ7T�� ��A�g�=g���"��_�]a�a��"O�Ix��a�3�lV PG@��`"O����$a��|�F�P�rE��$"O���cE7��e�r�C�P��	�"Ohț��܈^�P%��N4(d���"Ob`k�5�,�UcQ59P*��5"O�,��D�'+@4H�ЀOaR�1`"O��0�b�!w�^�sbJ+8�I�0"O��J鞎�&I���`%DQ�"O�	�?�}�e�A�%�!��"O�c�*�7 G�8�e���:q�"O�h��L#���՟.�(A��"O���3*'v��p���d�J�J�"Op,0��%�r��� ލdC����"OdEȵ� Rb1i�i�/b���"O��ia_'�`��j�%J��P"O4Iu��C��=�2hզBE�CU"O�yi �1,��i3��ME(��"OJ� �K�>��FDN0v`��E"Oȴ���[�d���#��8 �d`�"O>q��
���£o�9���"O����bة:"���H�!$�Dl��"O����E�H�;�EB�=��DV"O^��l�l��tZSKƱ�tؠ�"O���!�,BE!��P�%pp��S"Ob(f�L+�8e/ݕN>�"O�=�֦�@�8;��
x�<��"O���Gm�+�8 ����k�LI[�"O�ɺdfΌ+��i�E5ELh�*&"O�\kc�3wˮ`�Ĕ "/sT"O�Y+�#-�hP��ʘ4�@��"Oֹ�D @'�: x����V,K�"O�lhFE�Ty�W2�q� "O�Д&��т�c�>E����"O	t۝<`�t91#D�/�F��"Of�@R%��Jy�tOՊ����"O(i`�Ϩz�LD	ao�n��%Y�"O����Q�,�:�+���	\H�F"O��H�HW/XzJAR�"�y2�"O��;�	^`Q�Pbc��$A ��p�"OZ����Y��\��q�B�j��U)�"O���?y:$5����<��e�Q"O�I�A� �3l�<q���<��"Oz\
�V�BZd�:�H�"1�D�5"O��f��#39T�r��I4EM���"OV݁��\�֬� ɓk���W"O��!����4��O)L�`8�"O����QO�5s�&�cے�c"ON���GV�)���Z8@����"O�@[Va�<dP3��]����ç"O���w���:�^�#Q�.����"O����݀\%XT�T�x��2"OZ��$$_�G��%���A�<Ь�"O�}�C�<n�\�`
��^mڧ"O�`N�6�nh��Pk�BD�Y�<��ø.0 耦	�G V�{2�p�<Iq��Pt�� E;$�3,Uk�<a(I�rZ���![�0�
�L�g�<a�K�i	`�%NP�T"̽ʰ��f�<)���)2<M�bo�8'�q2fe�i�<�6�NkJ����Us"���)�d�<�q)^�3�V��3$� ��x�E�]�<%���.��d�ak,h�a($ȁW�<A����^�����T�Y�<� R��AO�c�B<"i�-L\0�"O���(�@\V��(ѡQ��"O�)P͖�F�|�#���k0I"O���"@<"B�x�C��g�-�"Oz��s��^DĈ��Q�'�:ͳ�"O��ՋL�"W|���*�d)S�"O��P���R�q���3Y�@�j�"O��WkȪ�� С\�^�1"O�UK�ّ/�LAòd*ذ�P"OP�bg����d�a�L�Z&N��u"OPcnD&,�1�	�f����"O����BN�<����0��.��"O��+"땭&KҔ��$�
���Ae"O��cS�%k4��q'͍�/�Ν�r"Oh\�tD,�N]3Ҍ�4:�!Ӓ"O�ݫ���& �	����Ȁ��f"O��IE$1�4P���!�H�r"O�m���(K0����%a��A@1"O��i�j9[��xK��߇(����"O�`(�"A�4\����=�N��"O.��`�V,T�˃J�
M�e"O`��s��Fq@�IF)�<{�c"O��CE��r�<��.).h�I�"OR�r�^�)Iꀪ�_���"O�����?}o����B_`���"O�y�B4m����e��R��"O�I�5!1G
���'=F4�c"O�@*�-����P��7D(����"O��@)6G���!"!f�"O���%L�`y���E��{yۀ"O���*M�Jʤ�Д�̢ZoJ�0"O(�H�&�4ʺਔ�$R<��"O2MsP�X=.G H�1�n��"O���ۃi���w-L^�J�"O��j;Z䱠��X>~T�0:�"O���j�52��{v�O9SJ�p� "O��#c�<wf$��j�v?phK�"O��t�Dk���� �:}��"O�sŉ�:,(,���E�a��$��"ON�(��I%�ȕ�1���y"O�	���ˏC @��D"Z���!"O@���=D�`�&�?.�2��C"Ob��BI@�KӼ��]��n���"O�+7%[�8"��pǅ&Y���{Q"O���$�4,�:,I�b��Pm6��"Oح�q���5�f����֭Gb"t�r"Oh3���ކ����JR�� "O`�X��Nj�Z��g��*Y< ���"O�-����#�Y���N�e�H�w"O�@k5��a�,�R1Z$hq"Ob �4���^]�%�����4b���"OH|�5	��J|.�@v��O�H"O���O���2͍*UF�i�"O�)�'�)�v���QdHl�"O�؈ǃ�=�su�:Ojh�"Ob���ӣ|Vȱ��Ʊm^8�Y�"O��ѠC�mM�xaܸS[DS"O>a��%@�((��m�1z@�m��"O0H6ˎ(��\�e�ͳ$ܠ�"OҜc��ƫ4x��Arj��A���S"O��J��͚$n������	pT0�"O����mJ+0F|sA�"0ހ��"O���	� 3T�pV%�,��U"O$|t�ҭ���� �!t�B�"O� *�Ig�*c���"�C�arn�*�"O^��r�Ξ�X:S�\6>*Q8�"O�w�A�Rm`���x�aA"�s>)�픒;�@RclDG��t��OD�=E�t
��:0��(�`��&��C$O� !�dCB�1��E��h$
A.x)2�|b�'�ܬK�Iߝ#�^��F�ۨX.ҹ�	�'�l��L�.]��
�KA�j���'�H8[�˧��T�����>�l8��'��1�U���Nz.����nUxy@�'��3���ΩIѫj�p��'V� ���ӽ2���
������yb��Jռe��4���Q�_3��>��O�|����Ѓ��B��i�"OJP��o^&*9�܋�@�v;TJ"O�<2į�Z�p��Eh�2!�t8$"OH�P�,;\�p�I�7��(qf"O��W��X��&�Ϙ �,�)�"Ot�2󇌚`�Fyc�S�8p�Y�"O:4a�oD@Պ��3���\�����"O�����=3U����=��E���	N�HH�Ή>�\ĳ�
J���k�%D��@�I�>W���2,
�%Q��!D�@�5�@&E��K#�;rK|���";D�`�3�
�<���iЯ
�I���<�
���D�6�':�ѵT2�Q�ȓ��hR�n�&j�.E��̋ v���?��?!2�+�(�4-��cTE�2�n8�ȓhX�Ѳr o&T�h�"Z�p猘�ȓd��=�SK%&R���Vb� qNF���pz�3M�d8Иh&�	&�ȓQ(�}�B'=!|ɴ��7����ȓ|B��Pp㋔9�հ�)�a���Ijf��'FJ���GK�!<|�	�ȓ �Y���%�x%j׎$4��ԕ'�a~���9|���ɐ'AmLjI�s��y�m��"��$@U��_��Y�'8�y��ŁV0p(�ԣA�S��i�!k���y�.���<�a�D��G�vT���y����o�zY��%?�
 A!�%D��9VG�>	��T�L?O�B�,"�O���*q!QW=H$��E�ҁ4R���IF���������O�?����u�e��<D� KsO(T㚍��AV�;^5�=D��Jt�K%t}(0,U�s{L�s� D�,QR�P�Q��-�$�:�k�*D����"Q �\�Bb�Y��xV�2D��ؔm׃c>�D�G��2Z�ؼ����O0�=E��k�d�L���Syv@��F�x�!��A5+,�pVn2rd�P���	�!�$�1l�4�S�R�~H��t�˄l�!�'F�]��fQ��y2c����}r��,CHo�H#���S� (C�A�O<�=E�d�	����V�C;n/v-iD�]�$!�-d�]c�kH^�F4�eG��L�!�,U�=�5��rxA���� !P!�$����
�N3P�pijEm]oJ!�䐉lJ9[Q�/~�d�+!�2!�$ĭu�d��D�+}Fl���R1!�$� ���q�U8.ƢYW��>&�'����8��$[�,���B|�{�K2j���?���)P�5ǖ({` ,�b��4�	�I8ў��ᓙ)`�E��FL��uy�(ې9r(C�	�N��`�;=Ǿ�`EJ�
%BC�)� �,�a��PU�!�× ��!�"O�-pS�ԷB�RE��ɰp��e�d"O�hh�ȋ�x��E�\�t8�"Oܥ�A�P�t�챋�Iƍj_����W�O��Q��ș>f�h�@).�&�����D��V�e�O
(��뵥m5!��Ρ"��A�w
P}B|I�ě4|!�(T=��Q�HQ M��jGC�:!�����eD���rd�Q!�DSez�z��Ϡd�����3L�{2���m(z��6��<S�X9��Å����0>1��
/-V�\�F�+�t����B�<����1>��Q�*2J8Hw�
g�'�ax2&��=��C$F{d���Ϣ�y�"K4;�X�G��:�ʄ���F��y�m+�0ˇhG*41��95��7��>��O��@�R(���P�$��5���cW�	Y��Bw
̫`'���樕�0�9+*�IW����K�R�òMP�c9jD�q�K�N�C䉞�ĩy�*.���3��I�4e���0?i+ĥe�L @ː@ܰ�U�@�<!�O���yhۏ?1X���!�x�<�Ì#8Վ��D��`J���"�t�<J{�Y�a��x\�r�u�'�ax2H�"4T��0��Ƽ5��Rh����'{ў�OGt9Y%��$<�x�k�v��Us�'�q1��ڈr΅�@�t>\Ly�'���{fA�WK�E��%�9Ǻ%��'hء��)C�>�K����̽��']d�맅�3)��H�cZ�H�'�|���揓��q�@Q!xE��'-dM�X*>@�2��Q�IU>��/O�O�|c>�e�+<����"T�%���p�=D��`�@�2�!Q�S+4(H�8��:D�X�ׅ_ v���뒙y�ީ�e�8D����K�w��0A�b��y)�-I�;D���q�B���ا-Qޱ��+D����L�;X�,�qs�9 �+D����A!�H�2d��qy�]S��*D�@r�O^�W�Q���� =����,&�$2�O����܌�!di��F�>�S�"O�UrE�\6�i�#K]>����3"O�Pi��߂l+
}���J)� !��"O8U2�JM2}�f�9�	��F��}hS"OaS�n�X���X�i��(���R�����S�O�,�[��4t�0�!�D�}&���'�p|�B匲5Lv��S���3�}�ȓLՀ�k�%�*��ta�]��d���4�d:�b؟'�$p/�at(p��M��Ze�(o��g(�����e�<�`Z�4zX���W62
\���D`�<��Ҹc��qb쉵{��DS���_y��)ʧpʢ�@\;l�0Ԇ����ą�0m���uaB�@C�Q��.V�\Ѕ��ev�_%x1��Vi�#,1RU�ȓi$��Pπ>,[��ޡ5�х�2r��`F?K�
Y�ΞI8��ȓ��A10��"z�:�#A��(U%��H����T�}�"mU��c�	�'���'�ɧ(�p����]�g��.޾}�"�"O-�B�A$r.␻���0|��3��|��)��Z�(`�g�
�d�\�jC���Ԣ=çc_�0�e�F	�f��7oP2{��ȓL�H���>�h���¥C�8X��S�? rؓ�JO�na<�;�k�&z���'3�dՠYp�u�q��$t|��rץT�N�!���3L"��9Eo�N4�H�[-R!�<a�|�#�ںxG6ܪ��J�.!ў����zu��2e R�G:@�� ��Y^�ʓ���hO���6)�P`�)�5y�)$kB
[!��ե��ݠ��`ɦ�8��*<&!򤕫J���$1@���$���H�!�Ě�f���`�7N���Z��P5t�!�X�ef\�@@EſiG�P*���$O�!�T���n�5�å�ێ#�!�o�]����k2����L�F�!�$���l
�H&�g�Ɉs�!�
0
pRhy�-��(����M�!��I iEj���ϪgbՈ�F1O�!��A�1�(Hw��=f�:9 �	�!�T�R�H�V�T�Q�	_�-���x�b����dڙr��s�A;d�V��!� gx!���	.3r�gd�.�*�`��̶_Y!�D4s�@])��J��
d��A�zf!�[�"��䛢լ�c��OYZ!�$�<?��8qp)	4�d�1`G0KY!��ٸ.G��醗��Hp-V�H!�$�:1�I�� Y�56$H����595!��i1��R�@̉*�xQ!SN�?�!��S	0bH!��oZ���M�#� T�!��"#K�%�P�۞qQ���^�!��&,W^�"�%G&�6�y��͞0G!�ā/<1V�
V�˭;�ޥ��$_�y�'�1O��h�f�="�FDA.�!D�tڂ"ODu���Ӂh��0�2NO�6�͘�"O<�2SM�<\��CN2F2���"O�$�R��̩06��B���"O��0��N"�3�IU�O�N`��"O�Ԫ��U:d�KXQ�x��k�z�<���Uww`��� cE&Y w,�P�<)3h-e܂ �u,��x1X=�D��H�<�hG2�\ᘑ($IV贚��m�<QP
i(J}�̠t���9FƆO�<9CK��;޶��6
Ýv�4k m�Q�<	�ɟ}�9rs�o�h�
P�L�<r`�i �!�$�-F�0���`�<	Ţ�4O�H�{��$h@�ҫ�S�<�wD�f9lp�EWmoD��e�<qS�Q��|�Ud.{Q��q DL�<!�ʏ9[�"1�ר�-x[�2Sk�a��0=��LxU\��&��h��&b�<a�J
@��PV��.a.�
���E�<�/�,8�fɡ�%V�d�`�bc�\�<頢SI��E#$@�$9l�]���|�<���A�'�ƴ�Ea/�Hl��Xx�<�Dğ17T`ŉ�͗$�0���s����`��= �M@u�����^� A���#q6`a0�̜>�e(�ɵ;$2��ȓz
�(��@Q��\)�R�@@�@a�ȓ ����˛$X[HY�3�[�X{�؄ȓ8��h�E�B\:��  
vN:8��2=��s�ֽ	6쌘E	0s̥��9��(Х���^ء��^!� ���5fL-s���GgJɉd ϝW��E�ȓn�"��?�
��/ԯP2�5��?�8�n$}��BMв����ȓ�Z�8`����Zc@'{k�]��S�(=�6�ڼq}�l��$4��u��S�? �ˇ�ЩG����f�3�jl��"Od<���
	����AI�;_���"O����C��b� 4��'I���X�"O�{T�]	� D�V!E�l�h���"Oniq�	xah��EgK)`L$�s"O��[s-@�k�DI�уD5}��8��"OJ�@5.��&i��±��*/I[%"ORMk`닩q)(�A�C��F"O~y7) �(���qv��qIlл$"O:T�@�O�Foh	#��(&/�I��"O�$�4b��I���"@Q=&��"OP"�HeQ�,RE�[*�Փ�"O�Ta��++ �ł���:m��F"O\t�VMHa`Xa��D
�`)B�"O>���!H�Z�`T��"P�u��4	�"Ol=�����-��Mc�BD7Q�pPp�"Oq+��[3hB�P%��6�т�"O0�#EѸ+ *����5Щ#�"O@��NX�B�&T���8bZ �"O��:�%��0�z`��K�:y� �"ORh	c"��1����jb8���"O��@Ͷ.�BSO5Z�(��"O<$3䫁8w�n5ɓ��,lU����"O�l�`O��C�@�y�� 0�#�"O8Ta�풯)e\��N�! �A�W"O�C�.ϳ'it4��ZN�X��"O�:7c��E`\R�,�)���!"Or(�A>Y��`+&&v��r!"OB�(��9?>���� O�`(lh�"O8 �/'	�m�� N�n*�("O�|����0�{r��.�2L�2"O�ؐ��(R2Ѐ&$Y�SȒ@!@"O�)#�F5s�Y�(Υ�p���"O\Hs�@8=n��h�������"O�+����L�q�Ϫ.��� #"O��+@��-U�M;�/̸ �~m�"O2!pEB�}{�1�P���0�Fm!T"O^��5ܓ����k�jpB�"O��!�'
.�4ř��YXr"OR̓`�F�4�@�S�!��"O�Y���d6��)A����T"O�ܒ�� 1M*���"�|�W"O��燏�"��qፘ�V,�,��"O����)L��\;��3o��#�"O���󃘟PnQ�a�+vhyR"O�E���!Fldhr��^��\8s"O���U�i�� #��ph�`"OM0B��~y���B��#�"O ���̚,�"��DA)j�6��"OF8�� �&.�EJ�E� ��hJ�"O"q(���( ��Ȁ�$=ga�i���A�O�`�d,]�
�*`�an�/�����'�y�"��Ut����(/��P�'�L�B��-;�\�h�σ�u2����'DdAg�P�y��}�wI�7i�y��'���c�R��'`H-��H�'� �y����q��H�7E�T�'ҔH���E5��`��T8~����'����HԻC�$�`�@ԺYL���'ؼ1��M�HMJ���	On����'@d��C�����K�85Zqi�'�Z$`u�Q�8�H��Ĭ'��(�'Y ���%�em0��sG�����'�}�go�.�������8x��� |u�â�L����0%@(%"�a"O�eJ�\�r)(D��M~	����"O����l��,��ԩ�%�=�� ��"Om���R��1I���^��e�"O�1��b���n�V!����x�"O�!bS�<b�dAZ�ꤕ#�"O��j�W�H̡t�F��Y��"O*���N�3U�miR��h$�s�"O� :�/A�8ʮ͒��L"2��mxV"O���ѡ���0��SlX �� ��"O*�ru�a�P�P��"�����"O �ڥ�UD�A)֙6��K1"O�xb�/��M!s�-�V����3"OHX{� �, hejd,�9ZZf`x�"O2���4O1��ۂ�����]�"O�E�`��(C08����x��"O��pQ!(~n:��$�O�!}�a"O��z��������.V��F��"O�=p�S�V� ��?����"O�5���֊|�
�F�L��rp��"O"��AȂ|� �+�#��?7<��D"O9B�E1"���&1��5�"O�1)!BԅsbM+����*x|Z"O��JB�լ�xY��C9^v��RR"Oz �p�r�:�BW._Q���"O�i�@I,'H,�co՚lG��s�"O4�귏�,����Ї�,6�AF"O��Q�
5����쇗FV�"O"���n���;�-�:����On�(�ZI�ڥy��Q��][&n7D�d	����SS�+�`���uy��2D�������K��aa) �0X����+D������g�H:1���m��+D�l�/�	-Lvɱ�*K�@��X�1D)D��ƊI @��	r�E+�ڠ@��+D���-�s
��@e�!��|jr�/�O��	�G����G�hl@��L=[�6˓�?�	����M[�lPs$C
r���`G�Є��A���񩕆[Z����=�؀UH�ـ��":�Y�ȓs��t�W�ߏ4Ό@�	7O���#��``F�e��T�a�ߨ��Մȓ?�2�Z��[].�(��!}����CHf��Q��`fJi���ʙK2���ȓ.�lX dʹo�`@�  �u�ͅȓ7Δa�K��{�$���>a��0��.׊���o�i�\�!�T�j^�Ԅȓ:@���t̓b,��ۺ}zb���l8�Ya�ɝ0=���VÉ3;d��se�p��E;fU���c@�A�ȓR�҅z�
]��Gŏ>,�@�ȓo�"���K�,��a�v�<X��>tA�_�vh�Tip�XM�ą�LC��q�JʻAl�}Z�͞0��=�ȓ-6��)��0e�0� �"T. Ąȓ- �%R�V*�b�e�[  `��+���	Aݲ6���M�'K*$�G{���,�9l��<	]6�
��W#���y�AN1_X��֔%"�tZ&�/�y��ݯ}�n[E �)JtH� &�4�y�l©"&,�UkS�j��P`�ϊ�y���+<Ӽ���cMbY0��7�č�y�%�K�ҜS�"^$lG�y�욬K��L!R�Y�%ā8|ʘ��S�? ��R'aV�M�<�s���!)��"O�Ա��4C2��:gL��p��"O�A�S@ŭ\��6�.��"O��
��E��|�Ů��(�N؛�"O
(I����y^��贬]>z �lA"O�����oEl�[E郯6b-�4"OP����	Q=ҁh0x�z ��"O��b`'�L�Ɲ钅��F���"O^\�2e�>kXD�p��v���"Odyx�Y�3Ɓr��#3Z�]�3"Oܵ�7.\T2��E)�4HT�a95"O�푣�R�p�d³(@�S<!��"Oj��*A
[FP�����V9&0�b�'R�'����h[F5�S���zh
� ����f�!�D�J3����Q���aPZ= ��l��0i�O	sR%��+Q�F}�� D����"��e�آ�H�1���,D�����k��I�eŏ#��@�g�5D��� �j;J5YUGM��\�ڲ�5D�� �U5U�
D�uB&� !�3|OL��y"�+=X(��$�5F�*��p��6�y"�0}O��P��YdnJ���%���0>�/M*T�ź��A@�N���bNc�<A!�|,TP�rˋ#y�|�R��\�<�� �~g�j2Hװ.4��@�Z�<��(T�i�������/p#�A���z�<9�b�ivp��BKʥk�L���Hz�����ȟl�).�ʁGןx����đ�I��9�ȓ���b� w��qCh�fة�ȓ$	<�Hf�R&x�b,i%�%:�<��
�غgɠ�x ��H�¼��s���b[;,���s�I�+��U��#�����B��cf��O�����c��x+�!�-3#�d�C�-4��4��L��8�E�Gdn�@"��R����5pE藚�Rd��T:ӊ���/$@�r��#�Q0��V1֥��Xߞ8��h-yc�0@�ܼC�u��:��h$'��2�(��$J�1�*���
hyQq����vEB��8W�͇�z	1V��c����D��7��̇ȓ�H8@����P0�c�36���ȓS�P��H3{��b`
8Yc|��Ol���az5t���8cR��*
t̻ �-/2��b��3qw½���z!`*�%q3���&�72�r��Rx�k�K:/�<�tm�=���ȓy
�f, (�6���3 *9��j`��J�>�-�牔,5�����l���o@c���m՞Ql��U����(�=2x2�BP�P�"J����`�2nן-}8	�񯊋1̆هȓD���(�ʏ�	�Y��oXX:ԇ�9�������4A)3��ۍ=�杇�^�>(��L>D�:�!�#��m⽇�`g��� �w�ց����
�x]�'T�	C����&��@+�b�����#5c��'�fB� ԅ�BW�I��	4m�EB�I�Y<�}ss���<̘����N!8r�C�I/o��������p���H���C�I-�0T
FnR�
vd���Э��B�I�[�(G�0� 脫�/�(�Ɠw"��(2�W�>"����X+�f�)
�'!�y F, �z�s���~=x,
��� �u�emn�ؙ��j�.��[�"O�ABqO��;��aw���<∰��"O&�(V/ʀy��p��!�$"�3#"Ol��wJݠY�i:�w�P�'"O�YXs�'-�EM:��i�OF�GkM7 Y�(;�H�^d۴�;D���`�� f�=@D��]'�	�:D�t� ��s��yҠ�ҺxT<D� ��"�8 H4�3��;6_�`��m:D�p�`ă+Z�Q9��16����*D��x�"p뚥�#(��^ތ��4�O�I�qy��1�,ΤF�`j3֣/�\B��6:	r�q�(E:oȼ�D�H!�?1��	�9e���w��x&�����9�'9a|��O"M��k�Ń�Ρ��ȟ&�y��ݦ15����@�eJ���yR��v��a� ��<Fg>�yB����gB��H�풤�G	�y�	����<��V&P���Yw喂�ybꄻz��A�M��L:����CI��y��07R�
%EX�T3�q��S?�?�����2�jW�G�LĀ�Z4�^�Bj|܄�ed$���A }�]�R��,v���ȓz�\XX��ª(͢��P�'	�H�ȓ&�D��'Mݠ��2�$&1����s�йХO��{���9�(�D`V\'�DE{����98�A�U�6Y��Bc�V0�y�M�>[H��b���4D6H����y���+z`r�8f�Ͻ��j�d��y���J
ҙ�� ��}��"E׫�yҁ��TI�}c��v��ҧ��y�Q8&a����#tc0I+��ˏ�y��.ϲᐰeN.b"�>�y2,X�{�l��jk��Gb���<���KUM;a�s��*$���U!�c��`�j�^����m��/�!�ɲt���(GǱ@�X-�v
�H�!�U
hw��%+�Np`��֥+�!�Aۢ�p������BD�� x���=>�|�+��HO��{��'��B�	�q���w U�ga�Qs�&fXC�	'6�#���	�"�zq���&ѶB�ɥ �2@�D $F�(�v��B�I+�����R�@a�!ڋS�C�ɋ:��y���%&��y�EE��+��C�I$1���L٢���Ba+�*o(nC�ɥ`	�����%/<�zD�\�F{��O&8E��`��}��&6xAK
�'3\���K ������T~kV����?�#�B*rb�ZĄ#L؞�P����y�!Q%x�Yb��E�o����V�F��y�f
�!��I�2+��qGrẆ�jI�ȓZ�䈕ߧyC�@���H
g����x-~DZ O���2�z�U.^�����e�����5 �\�f�	27����b�B�x����V�J<�C$B%$���'�a~���?Ot�����EłQ��#H?�yb�!]%��pë�'oX�jP'N��y��آ<n�H���;tA��o��y�d�� ����ل����ˊ?�y���qn��N8 r���胲��'zaz�!��a"nQ{�Ę�n	���� 5�hO���)��B�q�rgW��1�d��yQ!�d��d�ea��Ñ�1���>-!�� �s�$Wj��s$.@&d�]pq"Oڈ�AEɟX���2x攍��"O������Z
�(1*4Y�܀;�"Ob])��M�N�������Q�>���"O��(�@�1@M0}�$"֟,�>5y�"O� �S��0��xg�V5s��#PP����	5�f��e�^N�jJ��� o#�ψ�,!���C�m�"䘑�NR5�4��"OT,� mV�2͂|[�n�/BD q"O͛
�?*[Zt��6/� pG"O��x"�?=`a:$� N�j��'#1OD�R�;)e��SL_=x02��"Oа*!G*YJt]�k�|�Р��'<!��	�C�R�YSDX�-��,8��g��'�ў�>�3�	�} ��pfA�',w�����9D��eY�o���d)�Vݖ���#7D��:��J `��V���+�y��-3D�, ���!_���ǁV�\)a -<O�"<��JX$0���W.�(+&NT�<�f#ה.��d��p���@M�<aR��CS4��e� �T��q*�$
�$E{��i��8�����D |((���M�WUtC�:J��q�6ʝ�CNQ��k�lC�ɗIt(��#��/���S�`���B�I38�>9#v��� J��)z>RC�	z2�|�GA�27����-�#֐C�	�_��T�D\M��"�(n<9B�'�1�f�ūcd�Ē7���N���'g⵪e: ����ĝ3�nx�'�d��%G��)X)Qd�N?-ռ�3�'������3d$	�����8\�P�'�|�� n�� ���Z7A��P8:�'5��f)�iB�18I�$23�BL>����IRU����UƂ��&��+�Sl!�d�*{ j����dwT Z!��Ƣ<p9���61ojZ� "9�!�ѐI����ʱo���n�'g!�D_�`F�x�ƴT��BѽPb!�$��Ϥ����OJ^�Kv�A:{!���Kl4�#'J�kB����ɖ�w�	U��(�Lȑ�n���p��iz|�$�6"O�U��B�Z�����g��<cj�T�	\>����^1
(��ጮ�(���:D�*VÓ0^�t|�#�̹-���X�"$D�l#2�:Npt+`�+g�L�W�!D���gc�<;�%�`L�<�L ��,,D��X���K��� ��m1b�ѓ�(D�p�6�Bc���@�״^?�+��:�D4�O�0��h	� �0��|�^Ep�'��I}�4�4���B;�� �m�����v"0D�8�ԩ�8O���E�-?��J�-D�p��������,�=Wn� q�,D�l��H�-��,�'g��jՆa��7D� "Sk'1`X	A!F�5o��#�7�IF���<��J'Q�d��|X�C�*�XC�I3��իu�2
�(��Wӛ)�jC��*V�.�ȇ*	��1Q5N�?EpC䉵���BU�h5JC!I�`C�Iw+�mK�# �$����NB�>�2C䉾=����,�Z���|C䉍T�����Q�>�&x�g��> #�B�	5	a2�b��V�YWL�B�@B�	J��pu�@7X��a�f�4UG��� ��Y��'|����E�I㠍Bu+(D�� PY8��\���3A��=	�"O��k���VFT���b�!��"O�!�h;$�����)F4B"O|�⣏*v|*�����+TH�"O�ј`�یl=8@R�F,}h0Q*�"O��!'H��8x"�fB�-���*�y�ݣ,��\��
W=0Cp,��%��y�h
<j���"],���E����'����ÌF��~5so�A�\E��'�
��c+��a�>�RI��'�!�R�N֠T!�U>7��p	�'z��Ǣ]�U�jPF_�0U(i3'"Od�s�f��Q*a�DT9Z4XK�"O�CNT�*�����Dٯc�Z���"Ob�i��C#zԂ!��a�����"O�}�#�6Vx��qB8m�4)�3"O�8jf�O�[bTX�C��s��P8"O�,� �[>0�r���N�
�pX+"�`>5����+Y��j���Xt�3a�.D�<Y�j��r��P��Ǘ{�j�p"�(D�l��MF;�������d�y�;D�D#��W1*0� C<l�2��3=D�DkD���X��3)'qH�Dxu�<D�Ȋ�HE�B���^�AQ�M0�*:D��(�(��B� F\	�ZYH�;D��X@��q���x�HV+6.Y"e�8D��0B�O_<���k�^��I�	5D������:F~��T��"���KB� D�|�_�Yse� +ː�j�ǜ�P�*B�ɉ _lm8�@!M�x��b/ƟX�B䉦
��5�m�</�\�ۀ��Id�C�	�-��*ƥ�s3*�R�F\2upC䉂-�l��&�5jBȏ 8��B�I9O-L�S@NZ��1��S�|H�B��6?�(BQ�O�Asc�,&Y�B�	R� l!!c�$_�ΌRgOP�#s�B�	0\f����D���ÇmY��tC�.]�R�Xr�G�V�l�k�*�6C�	$h~�� ��4-ߺɫ�EO�?��C䉓&&���O�Y[vkG84C�	�	P`hj��Y�\p݊6EG�.��B�I'g�~!˂�F�F��R��4V�B�	���騇�R,	:հ'��3}{B�I�D)�IؠB�E�F�sS�B�	?���a��G}�)4�˂�B䉎J���2��=8���f�I3+w�B�I�/@�Y����"���k��	or>B�	?,�[h�<����ѨB�I)�h`�1��,}��:�+��>��C�ɽN�f|���A%MaZ��G�Y2c0�C�ɀ6���A�s.���GX�"��B�	o������0s��a�7Y��B�I�"X�0JQ�c�P��dֲg�ZB�	�΁�#�W4I�v�q'`ӐY�`B�	7s�S� I)GDb8�g�Q#,�\B��\�B��d�@�TZ�ea�qdC�	�J��	���'p7��.�$��B�	�[Ҙ9�,U
 ��u�ެRJ؄ȓ?0v�fi	*{�6�1��J^�=�ȓt)�iK(@�X�p��K��H��R|Ĵʵ�-�֩BC��[X�ĆȓuQ��/P�A���Ѝ
��� �a3D��`A��< �P�	WF�P��ey&*,D���� A��d��[���K�D*D�� ��A��K<���=a� �u"Oh|��^8V��A1����"O�P�cI]	%̼����T+f��Գ�"O^�����+bH�0��ҕuO.%�T"OV�dh
��B!�^
>F�j�"O\X:Vb�1CO0U�A,� 5V�zT"O�p:df	�}�V�q�a�T�Qp�"ORH�q�C�>0�iS���2"OlQ7����~�aOܗX4� �"O:r-�*8E�c��]+��k�<�W/o3j�����	\9�Tj�m�g�<�@�׮i���
�m�WAN�K�ϜN�<���S�92x����%^4�˓bR�<Y�J	�p-����!8�uL�d�<!bg߷̘�2VN�t�c�u�<�"�H9G��5� �>,x�o�n�<Q�ct�څ�GC�1WĈ8Gʏh�<�ro��\(�p���J+v�3v��M�<a��/��5i�J�e��%p�#�@�<	7T�.`b����r��4�z�<a���'��	���X����_�<���ڼQ&���G��w1\ԓ��B�<)3d�ks����.��-��K�Z�<y-B�1Q����L�*s.T��CAS�<	g�I/�L��S/�� pA��H�<��'�5h#,A-L,����"�k�<�D��"x��Ea B߬��+"�R�<�#�aߴ��g��;i,�K�ƇL�<	��X.�*P¬P2X��
L�<�I�"D_<��6�Tw�Ȱi��]K�<�6Iú5��)B���7nEa2�G�<�L�"�,Y�O2�AjD�<ٲ���YҰi�L/��U#$EHh�<)��;�Z��bg�$��Es��b�<�7�;�A����5��ɖ	\�<��Y5M��d���HYJY�<�t�&�ꍃ��?~�(��R��]�<1��'�0ͫ�H�8t p��[�<�`�+$�WE^�8cԑE`V�<�C�Ә�bԱ7��Xل���ABN�<�耥4���S%��\�%�"�^�<��F���xI��]��$)#d+T�@xRlM')�m��e�vFz�A$3D�ظ+�r���#1jD)Z5��q�k/D�T���3x����c�/\ ��C3D��z �A�ܬZ����&�$� rI/D��+�ύ��Q3���J�����+D�0Ps!F�}�᫵�
�M�\�w�%D������R�Q��I.C!ԩP�%D�����T/�����M�/D^8X��!D�4��qf���5�DQp�%��.4D�lSS�@A6��W-�w�ލa2�1D�l�դ�R<!'E"���ñ�+D���c�� S�ir�N�n7z��N-D�4a�g@�m���J OH���K�X�<��ϟ <+VcH�rFN[tb[T�<��螏,q>�Y�E,C1@1P�-
V�<�V��t�=ÁO�K,dPEd�v�<y��
!9� qL�@�����,u�<9�V�J]������=#\H��u�<.�&�����H����Q7,Og�<Q�$���j�2�C�_p`�H�,�a�<�f�8}ո��������ձ�y��/�"��VJQ�t���aq��&�y
� p����{���x�)��i��"O���ħK�� p�cCv�PAqS"O�xe̶�����	�%�ڜkp"O���@3TcŰ��<,���D"O���4�R�-�n��I�!�_� �!�Dʳ�0�Bϙ2�q��J�l4!�$I:1?z��IY�-,�y[q�@r!����d��$�^%����&!�D��CG`p��_@�D�%�D�J!�+b*��	ޑU	�[^���	�'����`ͅUIl<��BM))<^4�'�N�;'cC�"[�q���@�	굘�'�:)��ǃS��;��-j`4��'�d5ؑ��پ��W�[�|�"e[�'rF�d��FR��`��r�����'[��g׀J�&��$��p4����'�UB��$'?Te���+r�� ��'��T�P�'�41H��ؓc���#�'$�j��]�P:����TjZU�
�'����4�E����R�.KHn��
�'� ����m���ȴD��Ւ
�'��q+FCC/\��($A��C���k�':�HY�)Ѳ8s�5�s�D
jw��
�'��i����Dl���H�0n�Y�
�'��:UE���81@��J Y�ܜ�	�'�XảǢ���%�y@��	�'t����5^�9SrCw?��h	�'t��R*��x�؅����2�	�'=FA"tl	�j�plb$��/�t�a�'ߞyJ�	ҩ&x�2����z��5b
�'+�@@�KӕQ��Lx#νknE+
�'��PX��u>z��F!Phh�	�'d: ��OA��5+R/5xV���'�h��q�K*g�Q�23���'1$��c��WD b��L�t�D�1�'��Y�s �.�xY����!�1��'p.����}9J�z�_��pݡ�'��iS���7$P=qw��ĺ�"O
�U��S�.��3�Ra4(��"O��q�nÌpI���!�"O��1a]�@x����H׵i	0��"O�e�Ԑ�AǑ�[N2=�4"O2�1�*D�#x|�3g���'@���"O�p�h�� ?`Yc5�? X�"O���3 �A�\QR���'L�I""O,y�u�*���;&�M��1�Nd�<�?S@P���Q�P�R���x�<�񫄖l`8��; ?���!��N��uqef�>�V����ѦRZ%�ȓ9P�)h�El�
AkA%_2<��v� Q:�ϜZ� �g��x�.]����"ڎS�xp��	$D*�L��;����F�|���DSh�<��Ezr����-[�R9��+��X ��k#���1O	�Z��R�~� ��XZ�}��/f���jt�v;U���OR�=�Z����pe���\�zɊ`(Vk�<q�i��)9��J���0����E�j�<Q�m�5	h��G�%@�Y*�QBX�FybgVt~��2q%YXyv2�k�4�y2�\�[J.�aPETI�=aT C�����hO���,8���
����	D6Y��8��'��O޽H6��[�8�C�%�ft�$"ORԻ�L(=��M@f�˭A����"O� v`��/�5G�6L��� }�����i����.�i�p\T�AǇ��c���>���<Y�'��'ٛ�� {W�ɑT���-E�y�֯߫�yb�S��4��R�k�����H��p<���ĝU�jU!2���=)ūE
XBa~�&�|?��&��#T�<�z��M�<�t�^4���b��.�*0
��a�<��J��6!��2$g�t�!M�^�<	�b��(�)@��G+5���^�pjV�z����O�3���Q6�l��kƠ/� �"O�����ߜ0�\� ��~�
%8!�Ol���=Ѡ��	6\V4���A�~�.�ұ
F8�0�$IGU}�Ɂ$,��ْ&��Dm9���M��'�8ͱp�6t\�R�nL�1����'�I�e�%.��W@ķ2�ʹS�4�hO?7mչs��p�+W�49���Dњ���-��?��J>A�4G �1b�J�,x�,kgK^&|�|Ʉ���[S叵:u�Qa�A7h����<����i�> f��uH�3'3x��a��$ab�O����$C�4�&q�c[{��u��1LO�8S!g���̣lgN<���ɼ�h����Տ��P}�ce���A������������)�'Ƙy4 \6F�xP3@	ը,�.���	�<�{��E6}�:-r����h!�*Bƭ�y�蔅h��Q�\�S�]���K����wX��2���o�ܵΎ �%7D�$AãT�v��U��(R�a�6D��(1�2(�@��u�BZ��� D���"�
1�"�ʙ�P�@�1�)D��R��&��:�֏<cհ�I'D��6Ɉ:9$dr�H_E��=�D�8D�8��H��_�D́�nФ'�X�a׮5D�@'&�w��p�Eܔ
�jy Ԅ?D���Pl�$O��-I���.�"��=D�X�ōȌo�XI�m�N�xz�N&$�D"b�ׅr�t�w'O�4I#���y� (O�H�˦d�+@�V���Ł��y�|�tx*͓:�|��2%�&�y��%'���
`��<7�Z�c�U�y��עb3]KF�8zqR�۷��yBK�J�e����gX2e�c��y���.5����I�tt��'H>�y"F='o�U+�*�>�4Xjg�[ �y���1�8���14��ܲ�e@�yb���~����k�3&�=�P�L�y�B׶2�6��b\(-�F����y��Χ
�:�J�j]$��u�� �y2��0 ,|�:GY� �%���y",P�Rt89W��T�@][r�@��y�E���]�ĤV�PN�aԢ��yRD��#���(��L�|�r�3o��y�MS�f}�mZ�}��吮�yr`¢KI�Ah@GR��S��%�yR�ۛn��j$�_�S��y�պ|����#YXa�乁���y�5~�����J������y"Eʼ ��iP@��B�t�9��%�y�[8e�P5C��Y�n�
� Z��yb*O�CG��{s�M�vI��"ֆ�y��l�XQ�p�V:�e(d�Ҕ�y���J��ȷ��x�2h��hU��yRÛ T0~�q�a*u""�B��yB��=D� ��!ޭq�h�q ��yB������h�ꡩ� ��y
� ���S�M���r�R(մ�pB"O�C��Y{@�ؠ�O8|��DY�"ON)���U�!$����c�l)��"Oᑶ���VM��ru��,f�`��Q"O"HCF��a���q����0(��Q�"OD�we�7a�R��k�"Y��S�"O�`A���|�v�h1
A�#�"O^I���VY���G�V��#�"O�� �r�p����i"O
m �ꗇc���Qa�Ӿ]�������9LO��*w��B�$�F�Nf�1�"OP�����/y]����= >�U�C"O��K�HAuV�؃��X% 8n ���'o���b��2(;v�v)�><PHʦ�=D�0ɂ�I�>����'ƃv�m0<O\#<��$��O��A�aQa�����	Qt�<Iu�'2>�![��M�"84���@�k��0=!P6�\Px����?Yb1ZT�g�<�c��u��934`�4d"Q�C�ʟ����7$R}��hU)X�`ʠ#W�.]����_n��Fb����`�i�,ip"Ox*�Ȝ4#�G�V5d��;��'Q�,@���+��=�V�y%����?D����"Џ9+��&��p��\봩#D��+���*ZH�	֕^:��s�#D��
r`�'`�U)Y��j��e�?D�L[�쁖{�u��&�.$p��-=D����
�e�4AtJ׿2MJ�K��9D�L�� W�nv�m�ԋ��Y�H�B�mxӨ�1�)��ЖG՝k�Z�5�W9�lMڲ.;D���#���*I�pO�r�,��c��<Q6�'�8@ȷ,Y 1򋗾a����'�dK�(1�%3F�M%"���M��l�`�Dz�X6M�J�'���O�4q�AT+%2�{�J�OF�C�"O��P-����E�(Ic:�q*t"O��!2�J�)>�s�~/����'~�ɓh��i�%ّs����k6IV�P��,�|���צ<��X ��̓3|��$2�d�6V�\�s�K�JG"Q�"�!!�!�dˌ[�ntP�ͭR֍�oT�MJ��Ay��)b�M�0ɴ�bS�Ǽq`z�S��O�<���	&	�.��E�$	���K �QH�<�%otx��$��c/Z�8字G���d��H�*�晒d��J�H�EI����
�?y�Z���PB��2#�Rũ��=�'a1O����� ��A?����@	�@��=D�Tv�=� 3�Ý� �Rm��O^ꓮ����N%� i(Q�*@хc��&��5C)O��=�e풧>��@R�'Q0-����$(�צ����'�Q����ǂ�<�̩4�6O�����*�O7�;?�c�CC��(օ�+3*�����P<��ɝ�hglp��F2��yU��N�'F�b���ћ�T��8�T�B֙^08Tq��3�y����|�z JL!�Ⰸ�k�6�@�͓�򤨟�g~���X�EA�l�V8�p&A��ج1��+D���b�9(�H��r��*u{ʘ�CT0��'��Y���u��.O�(k��� X�9!�?D���0e *s�	�Gޤ��)�1*>D�$���^
9�X$�pl�*Ԩ�"cN?ʓ�hO�I?�%��A^6._��Qc 'DB�I�x�
! ��>�$-�th�-�S����OJY�3Hժ7
�k��E?�dJ�"OB�z�`�)64����0��	u"O�q��ԡCҰ� ��ӯ���!E"O� ��B|6�Q��ȋ<5��<�U"O�}:dw*�X��ŕ�f��Q��"O�������M����撑V��5�5"O��a��Μ~`D[T%�5L�� ��"O���Fŕf�ıG��q{8��"OJij�MʄAʘ�#U��	\�6"O�a���{p��6�J)B"O�ڱ���f��E���_����"O�a�ccR!��-�!E
x	�u"OĹ�	�$0��$��5��I"O���ɫUa�E�Ԏ�51J`= "O�ѡ���s��x.Z ? !��"O����զIxp3ã_�3.|���"O4��@��W|q�Q2�j�"O
A#RF-l�������"O����&��`s�֐�5B�"OL!��B��1�	���.$Dk�"OF5`������_+U�Dd9V"O�cs�#��`���=���"O��H��۞Sj`�h7�E �z�J�"O~t�ǅ�4�Ɣ 3G��B��h"�"OP
�N�=sC�� �#o�ċV"O�	q��/�x��W��,[d5hd"O��p����Q�����OV�#"O��ku��{E�����̀H$��X"O��Zv�P�F�ɂ&ȅ,B*�L�"O�!�)TTn�1v�]?����"Ov@#��1G���'G]&UG�Hz�"O��c�K�e�I[��ߵ \F"O��A�@�RfF��*B*�$"O�� �Ɂ b���aQ9����;O4Z���F��H��.���XC�*&�t���e���ҡ��*��5��'�\�:�O 9+��1O2>��K�'<��vc�9~Pt$��
3t�A�	�'���q*Ԧc��y@�K�^��(i	�'}�V�ށ��%��[�#z�U��'��X��h�;H��CI&����'�/:�@WIʑKG�a̞��y���-1��Si�@!o���y��W�)�i������H:�	��yǆdd�����.�
�P��Z�y���6�ܨ�
	�
7��p�<�ӭ��_NN�փ�8��8��UQ�<i��ߥc@
̹7��:v�+E��L�<���#M�-�'Y�q��s&�JH�<���0¦PIT/��Fa�E�@�<E"E�p���ȵ@�$d�ې�Z�<�4����{e+Ǯ]���z'�U�<��DЭ#� �@�*`΢����k�<Y��6(�j�PŤI:i�(8���f�<�f��퀴J�=�X!�E���yR��-M����̌�+e4J$���yB�T4հ%S('�тs�ʤ�y�GǊ3�*DS�֝NlN���E��ybN�@�a��M	2�I
�T��yR�C/����7�H?Q���ۡ+K,�yr ʈ��P�P���Lr�d§D��yr���H��4�d=0fV��y�ōI��eYDm5z�
���B��y"�
�}�,e�!�J5z���p����y�CS�Ӳ�R%*�܀�ٶ�yb�GP��y�)�/U�4�V$��y"/�1�dɆӛ�|�����y�H+z��9�W�?D������y
� D�E�њn��9�/ڳW�,�s"O��p-)~�N��g2t�"U��"O�M�#��d
�!KP��=l�YH�"On)��FǬ��Kͣm�2�v�D�M|�����@�9n`�S�C�C�� �T�Z�2!�Ƶi_Ȩ�w�E �jMɕ�6�`H����z�ɪ7�Q>˓/�>@Cǉ
)1#�Y�FB'aZ��\����KM�,�ه�E)p�Ʌ�
�J_�����2�O 
�N&u�~1��Ϟ!�ԕc��'�БǏ�z��9�C@l��0a�K���@�j�&��Gr~u(B�ńs͚�q`�(�ذ�<	!�]*���It�7�M��*���'m�� �*«Fj"��ȓy�.�� �*s|԰$��$,:���'n�|
4�'Z~�𙟰���W�+�Ʊ�W+��5,�)�.D�X�Pb�RӖ��k��|^ t�1��	"�`K�-X�c��|����D��,��V�2�A&D,�0=a� �)G��0Cb��?a�ST�82�L�t8����M�<17�U�N��h��j��pU��gWE̓�~}�3�ևpVe���&
��z��N�J/�%���'|��C�I�hR���	[��9��A�qȍI!&ԑ}F����O>����3?m�;F�y I֕=���b�Bm�<I6�6wʤP+gLY�EM�=���#d!�qK׬
�ẁi��?\O��qRO+N�Q��ˇ�>���'@�tˢ�	�	�I= @V�s1��"gJ���g�ǘ��Nv��3e��*YviC
�Wδ��>	��ղn� �q�����(�h��U�>o�n������Tx��	�"O��2�ER�1��2�_I��Mcp \� W<�Z�Ï
��)��<�3�4(�q$���P���D�<�����=���%NG�.9@m��E�<�C��.[�`���C4\Ojl��c�"6&p�&�<P�@��R�'��Rt*D�Q02x�!Ĉ��̭Ґ+Ƥu �`�ح�y��L�W:�T�C�w6,�B�Ĉ�(OL�x��U8�"}z� ����ȗ%�2QƐ@��V�<�S@5��H!��)	:6u���G�����(qO?7-ʂW��1���m�,T0eEI��!����!���N�,�tѢ��g�!�� 8�X�O9rd�u�f%�!�DT�
^��g�B�Ĕ�%U5a!򤑆>u�� ��V<�h��&�x !��ĮfB��� {�ڈ04�D�4w!��E�t�n\��@W�����FA�H�!�$�{�F��F�	y�Z����/O�!�ěS���Ӱ`|������A�!��/XVM$T��+J�E�a�ȓE�L8`&�v�P����D�Z4�ȓxM���Y�z��ؒ��%.r��ȓvM8<�GI�X���A$ L������L�T!"�� ��Op4��-B�`�V�] L��N�ON�ȓ|84]��N߶n���B%�L��Q��{ü 0�	.WY��BC��2DH-�ȓ6�����w�d F#���֡�w�<iIΪ\M.�rvlƤm�j`AF"d�<yA���5=�{e��CL
���$ n�<AT�P;�8��d�R�Eְ���Yk�<�����RR$��`F-p,��a i�<iբЖc�B���#N\��G��i�<Ʌ�W5���S!n�y�m�j�<)�P�
��I�f��u��ӳ�e�<!rh�:| �91i��eڬ���\�<yBD�X)8�1oD�� �GX�<�CHU�~@2�'��h�dM����a�<A Vl�l-��t
��ɼ5Jt��C��c`C"+fT��Eɕ2�T]��S�? 4�AGm�&f?6�3�=_��
�"OB�'�O{�fM�7b�K�2�"O�L´�)-����RM>:�"O���R��@�`�F�V���"O P�F)�2fm|�B)�.X��X7"O��3�'Q ��	����J� �:w"OFK�(� P2��@� ~y�-pc"O>�㛓�H�1MS�\���`�O<�#��D�;�f2;{|�x�Ꟶ_U	�'�^k2N<D֚D؃K�L�L����I8k�MK2A/�S+`��K��>T�@��Njb�C�I�d=J�@�����D��qI(����e�R	dj�ӧH�@Y� ͚5���`'d�:hօ+�"OZ!�J	b�����QO�mӣ�5}"�K*n�����+���ƪ����9\R��7'a�F��P$�D.9Mp����PJ�8�5&L�H��?��I\�s��|�$�*c䢹��NV�N(��
~�'�Zs�-�<r� |&?MC���s|ȁ2���
cU�Ӝ<F�C�8S"��N�"~n��*+ lvf��x��!�s"7-o��2�b�[��H�ӧH���0C�ՇA&j��CJ��N���?OXyT�F�>�\8�`��p<A�9�(q��ZR�T�#�N5��������7��'i<@moݸl՚�i&��73o<���B_Bn	S%�Хf��p#��'���6&͉TflbuDE5\H<3�����x�'�f�	�u%0����N�����k�ģ�z�(�K�)	��'Ԣ'��Eb�H�w�.` W�IT(tNA�2 �YT���d�'~B�j�&)P �%e��NDO.�H����P�b��q@R�l��M�i"r�6&�b7�)�'}���*􍉨/�@0��*ʸc�bQ�G(��@ڔ���N�j������%��Oj=�M�N+ݺ���<P�^��r�OJ}J��V����B�R���'[up`�w
�	1UX�*����0�𤘃!�6b�N��Ҋ�4+oT�:So�
��?��kʲhhD����0�
���+��8;��Fm�A# @x4��0�˱c|`���4�*�G�����qص���8��(��Ox� 8�J�[��s�� �ڨpq��v���4H� >wfEb��̈���!��<O���gצ#�Դ@!��^�O�[�J��|�
�rB�� ��U�Ɂ�ƍ��&^�F����"�4�b̧��T��G�38�`&l�Kt- p�O;Xj�`C�a�����׃֑�0�P8�7/�
^a	Fb'&#D"�bC8}@���aa�e(N@2R��aj��ō��(CaBR��B �ɶF�	Ì�)x��Y��͑���`c����x/AU�`tau�_8/�xD�pO�b�Xx�HG�Q:쉋�l	���`�I��
(��Qq6�c�թ�� �0�q�T�'%�1�UB+|ON�R2"ۢY/���f�@05Z6tK��0��E�r��G�x9僷�.	�!o�*B�Px��23V.\+�S�����c}��ѷR�vaR4F�-�Ҋ̦��'ZR��tg��k�Nłf���m6�h ���O��
3��	!!bn������C<8dl�m�%fE��(��0Уs�6�)x��" �$6N=B%��<vk�i����(�$Px#�Wp�S���*}��2 LC%3�$G�uc�A�GX���](��{��":YЧJZ��?��(�@��� u��423\���JW�k��,�h݋U��D++O�12�h#v(V��R-L3䝒��w���C��B�݀f�Y<a��t���'Ԕ�C���p�դ�(fL�m�%�]57)��Av�.>(\��'ꤥqQ�O2	�|�0��< �"�:���p�4�p��^~ҏÙ\d�r��BV�Nd��O���'4��Apច7��z%`X��t���Yh3D%a �Qrb!�
���G�ƸpPHB�"&"��� H@�|'n��j�`�1�fY�������$��ǟ5\6��yd�M �XX�o3zy�Q�UB<�(�'����KF~b<s�@�.c��� tM /�����'���#�W�D|qf��
F��#�n�����C�
*��q�'e���%�[���"�P/|���]!�qN[B�tݓ�kU&X���d�T�xh�3�A�B^V�AN��:�}��)L�H�iJ�t�`j�8T�l���$�:m�Fz2lJ!0z(+PΞ�M�A{E�>�0<�ca p�e��'��!Y�呚}�Є�$��.���Q�BR��u���J��E�
�@�����baIB�M��Ii�A��j%}�� F�����d���{�`ݶ���?�BA�z������:I;a�"D��cH�EҤ1ʵ�ř-���AR�L�����c��&�"}�vj߄D��,����REΔ��Ts�<!��ޫRI�l�5BǀGDb!1�)Ta�FFf)!��'ֺXBR��"�l�6�Oc*�0��'�.����H�*����._����'�l��D'i�Ŋ+V;CC����'��궨�u�A�M@4;����� \�IeH�6+�Ax��D�5ev�p2"O������2q~y1sCC�7lH�Q"O�p�4�MDjgB��CC6��"O�ؑ�ڶxU��SEa<R��D"O0�a���J����	u�H0�VoL�<�f@���D�Z�*�  �(�Ga�<١�ؓN1�ɗ�O&c� q�U�z�<�wSq��x��jܯMy��aҫ t�<QD�++�!��ʗ�u�x���	N�<���š\^��"g�M0*`��J�<���F2Tt�����#*8���6��A�<��D�W}�����&-�ȐG�H~�<qpn)n܋��U
4&X� �{�<�q�J+$��%E݀~t5P��O�<���0Ez�ӱ�Q8>��$����n�<��o:k"�D�KF,�m�)�e�<	�dܧ�X�{���,g�v��Ǣ b�<a��ЪYQ (�a�XS���k���a�<94��A|�`%�6�pX���@�<���ɰՀ5��B�?'�Ir�O�e�<	`��x��(ى�*���% i�<Y�睹6xRLJP"��C��}!��Rk�<y�j@2֌�����轛�
c�<A�H�\�<�{eE�9ihX��$��f�<a�`ȫ-9��°S�AQ/L]�<�c$��FlB\3h��Q �����X�<	QgB�s�~�KiX y�D�K$��Z�<Q�G��v=� �Fk�t�a��x�<)2�� ]� ��
�v���Jßa�<��J��%a���<l:�9�*�+{!�]0s1��襬X����Q�dB9
t!�dON�8��@� 9p��ງ���-C!��T�����74yʱ:5�K!8!��� ��˔�I9'I `��/4!!򄘾]��Z��v���	B$P!���(a
�1��)[�l��`. !�X=6_�a�Cݺh�r�8�.ųE,!�Q�Q����F�*g�pB�MĮB!!�Dya��؀@^R��LT�q�!��ӑ����	@Z�Y�+�9rF!�DҒ1����r�])ODZa���I�ZS!�DE��H,p1���\ �ȥ�d!�ӀU�fP����9�⍣u��7	�!�$� fJtӑG�i�"�s2'֘(�!��G�@E��%�
�|IYe_#n�!�E1I�~@��Ϭ&�N�k�ҹC�!�d�"l���E�b4��� T�!�Ě'uXԝ�j���z�X�"[2eC!�ds�YɃ)D4��ɛ"��8S�!�Dʎ&�:	��F�E��H��Oҁ?�!�D��~���r�۱!}"8"���v�!��ױi�|m�J�;m*e��V�3�!��$0��bakA��ƈ�k�g!���,V�|�4��:ђ܈cL�*!��.���,� �\|����)�!�Ć�bp�f�V�&j��]:v�!�$H�+���,Q95F��cR�c�!�DŜq��Q�S��~B
�����c�!�Đ�q?��H��>!@%
�BL1�!�$�� �Bd�e�=F\@g�F�ym!�ث{�r5k���P,\��eMYE!���B�(5�e8 ��#W�/2!�ݣ{��PР9��m(�b!!��8l`4�#�"�HXpR�S�D!�� L�������42���g�\K�"Or��%��	��$���.�\iS"O��)Xњ�p�Oek�H�"O�T끅@)gp��d$ �lf(�x�"O�e��/B.d�ɵ�Hr�d�"O.l��l^� B@Z�}&��"O`�0$����:�R�#]�5a�"O��b��4z�e:1c��o��DD8��*��I̾T�&��1��R3��)VE@�!�d��7�$2���E,V��!
8(Z�QsAb�I8)^Q>���9�+��:QD�h7�#K���ȓ= A�3j��/מ�b�C��!��������=���R�9�O�� ҄��kM�C6��?��p��'�9�Q@���V0�"v����FoX��4dш&D�ȓ>��E�����e�eG �3���<�5���5��9у�=�',j8�
ͣr	89�w(�	UT%��pA�ݪRe�Tr�!�&�L�xha�_/)P�'�<퀊��[5�N4>�ڑA�-J-%�^�#)D� ��U�E���y�F�FLY�Ή;J�8��U��|"�e1d�ICE���f���C�2�0=�r#��I����q���?�"cނ�x����F�Ui�D�K�<A�(%H�b8�sfɍD��8�7a�N̓E�����R�7��A�t�0��2��L!c$�����8&�8B��4~Rq0�/�Ik�A�
��0d��!Ԇ@��D���O���3?��V(m
�c��)cx�q�H�<����i����3#�B@j*p��h��[Պ� s�,\O�����6P��C�����'Uf�x�'�mM�I჎�^�ƌ�D�0W�����/G�O#$Q�ȓ/����J�NfP�ءʴ�>	V(D1'������+�(����5� N���F�QD���"O��z0)�CEмK���H�n���a�(��P�䍺��)��<1��W.Av��ȅO)m�Rcni�<Y쎆��Hȡ�^[�H d��<y���ŀ%�!\OzY����B-�-�鋦��Z��'^0	H@��E��L�WK,{��zե�}4`H�$���yB&�:~��$�r?<a"c"݆�(O�eX�� 8 |"}:3�،-�8w!��!��$H��XL�<1Uj��� 1R�$�M�6i�ɦIBU��$GqO?7M��Xi���u/ɱ>�V�Y3��l!�d#<mB@��@�>+HMJ��!�D@��.�{!D�-���ռ�!�H�a��l��I�&�
b포4�!�D�9֔�����"X���RF���E4!�
�x�n�[EB�1�~1P�̃� !�Dg�9�ǝw�dђW��K�!�$�7|l�#�d��!� t�c�J!M�!��[IȰZs�	o�r([$
Z�b�!�d�DX��`�1L
�)�U	»�!�dU�R���Q�2�yį٧2	!�$ـ~j:`�9����k޾A�!�ϦK���R���ts�!����!�C�-��yv@H;]~̀�WL�o2!��U4̐Y�v,��`d�y9d��\3!�װz&bL�P*͈]�p�a �Q�O�!�d�z�l��� ��ŉR��,o�!�d��^��8�JƵi��8Q�[�!�/dw8!;�*#$$��T�K8m!�DCQ��1R�
\�d�M3���(L!��ę;S�7�ֵh���/�B	!�$�:P�M!}�h@�W/�!�I�z��`;ҤT������;_!�U]jИ��R-�d�0�gʪ|g!�I�7���0�I:4��x�e:C�!�Ě"�P�է�&6Q>|�pM�6c}!�� ��9s��;\X�PA�;-ȅ��"O@t`#B�@w���IU~�z��"O AgBµ0��a�ǥ��� �"OZ�xbB��	Ԗ���g�k��@!v"O*<!DEp��t9� �h�V"OQ�#�F*c�x2E�z�z]"O� �ǩТ,U����dΆ�u2�"O�A9�$ʜR��%�!!�c����"O,ā���N20��`�����f"O
���p胀�	9���B�"O,�j0���k�����n�#a�r��v"O���'
-��d��T�3���KO����`5�+�"�VΆ�������U)�@6���gQ4���L�*P�Y�)�E�PxL����O��j��[�W�-`Q葫<��i�ȓR
X�p�Դ~��`+_�<Q�'����#��\��O�>!��b!�*ype�j��T`w�<D��R���JФ�F"�E���8�M�k��D/q�@1��l�o�3��h#�B�-C4R�+B <�����U�
�ʣ�H�=}��!���![h1e�X�:`����?����cѝt��B��/P4D~�lP���̘P�a�����lG"}4��K 6PC�	�{��u����%C��ŰB8L	|�~� 1R$���ӧH���6�I)
*w�aP�"OTV�{�&)��@�Όx��=X(�2<�9��*���&>c�l��Ȉn�f�1c@1_��\9F(�O
	���x���RI
7~��`2h,Ԭ���)����?�4��&R��@�m�Mstkp�'^�X��E1��m˵��hM�p��D,͞1�D"O޵
#/E�e����1(ͯ8�nݲ���<ѓ#К^pqO>) n��4xp��/U�s��+`#?D�8�_(m����:jj,�w�9?
��	qJ�AC#�r���A��}�O�"A�s�̳���&Z�.-D�@�'A6!O�T���PeB�&����P�S�#� K�Ɋ�P,d{�oX�����f��#��*e�5zK��aT���dcR�!Y��� (�M���B�@��q�`��$i�&�2�_�z8 #d(>�Oh�Jf�L�"cU�BA˝d�'�p��
�k�2-��ٗ=�@�R9�~,�2�U[R��FŜ�Y��5��"O�8��̕INb4QQ�Ê{+�p���A��@�$�G��b�ľk h1t`���(��d��b��Yi�_�]=�������yBaАY�|�;c�^=�~��s@O^1��k�>0���3j�8:���O�x���$��E��X�t�ȃn�����{�{�h2�෡��@�@��
<#��2f�VS\U(0�G����b��a���(�\4��d�1@V���΀�6\�@EE���O��8��]6f��h�A��,zM����35��/5���ZV'_�tF1 u��d��B�O�)gq����	=�B Xm��+���?.��/�L̃��;!�=���~�V !D��*��#=,�ٟw���Ha+A0@9bmF6aSd���'D��Aլ9J09�@�LS���'�R��$R�@�ɗ;J�����%"��B2)˂6�����$���H�J�v�ҖGu��{R��.hu�@wm�!�f�0��ⲗ|"�ʐ�ų��$�mR`t�cɔ�)����֑� �'%ς���b���w^\lx�f �	���$P�O�2
��S�ˤ-��ԎMd���	���(���Џ�>Q¤ ���D��B�	�a}"���j����`�թ[�
ɓ�lB�q` @�v�
)�V�ڕ(�
�"D'��$i�������wo.ɒ� ʄ6�0!��
��I��'���j��C���Ή*d� �2k{��u�BÂ�g��=%�|�2��>`��!-|� �5�DtAU�=t0
Px�b�39�� *b�'���#��X\I���Ջ!JJP1�ki�by�� �S�䗽�����!$>�Rd)ғ<Ô�!VD�&-R�@���'}DA��I�#�<}��G��<�c�Z�d@��[.��t�:���1;Ѹ����ּF�h%°�mx�����Q�%ľ\�6d\R�Nj"�4}R-H��:����c2K����?ٸ6 9��@�aQ�n��@�j>D���Q-�/kl�EH�J�?�n	k�&�>i�#W��HL>E��<��H����\e(5�'�yb�F7kK��B7"YjV����5&Qzv(,,O� �Qj#l\�A�(�v!��h�c�"O>z�D�-��iJPa�$!׈H`"O���ԧ�� <>�#@�S���X��"O�q�C�֦D���jb�[�;�ց0�"O�\���՝*�-*fM\M.�(�E"O�< v��OXR%��Z{.YQ�"O�#�
�bX5�C!�%-Q�"O�< �@'O6l�"@%y�T��"Ob,��#6;R�H$�͉X̐$"O��:��Hx�n|+V�[:S��d��"O��(0%�#=��"�H�k�"O(C@O�3B� �VK��R�Z�j�"O�٨�D�-2���x�,äv�j��f"O��g�?�Q1��4/��0"O��B��$���;�����L��6"O$u�7��@\T��ႈ|�De+�"OXm	 aT9��JU!e�D�D"O���ӊ�H$z�j�	>��dp5"O��z��R�F��
�L��fl�"O�*��̺wP��Q_�s��r"O��j1Èغ$3Ǣ0~���b"OF)��@���Txc��42��)h"O���*U-�y[S�� ��"OT�(���u�8�ڦ�O'my�U��"O������#+}*��F���y|��"O�=0�`�,�*�*5 �he̸A�"Op���!ޖ9�@�*�-T#Oe�B"O0ٻ�O��l�(���]7��A�$"O�I(%�۔g"�x;��1��,��"Oh�b�_�l�A*��It
���"O|h�+��jǴl�d�
ZTlHyP"O�aQ���WȰ����eW:�ʱ"On�K���V�L�D��@i6 *2"O��Y%�E>0�nQiD�V���v"Oh����"�^�l)R�R�5"O\%��ǑU���㣉M�c��up�"O(�ˀ�ȤpKء��
�u���"OL�� ޿	~�hAh�{�z-b%"OD�0��P�&i;���::#n]C:O�up��S5$W�����S�Z�{��	���4�4M �Rc�q���R�ZC�ə���qG重#<��s�A$L�DC�f\��3㞜=۴�3ƞ�C�	D4p��'b�qQm��UזB䉟7޽3F�Oi���㦜�xnB�I�2��1P�g
5�z��V�g�$B�I� v��+�k180|(�d�!VL0C�I�V0��R�SЕkj��5@C�	�]�25��
�����,v�
C�	�(� i��Nph]�D�
�U/�C�I�_H�PkҿJ���(�ĉ W�C�ɖ.+�8�"e�2]G�0����*�C�b��`H7G�2=�L*�
2h:�B�Ɏ;\j�p�S* �@�DmH@�C�	f<x���Y;t@@|0��Ƥ3���D�Y}b�̾(�%�u�{i�U�`�R�ē8�Ш���8�)��=~,�aRe�G�7��A��i?e���s=��ѵ/*�)ҧ`G�@ ��6 ٮ��$�G�̽lZ���9���Ӝ
p��%�^#M�i��jC�	]ɡ'Yn��0|��mO�1�V�R��	!.S�0pci���'�\�$��>1�l�o�p��:E�����F��hO�O�8�&K\95f�����x�[�'���rl_�L%�0b�C q�ڍ��'�����K\�Ui�I"U��T�� �'�����Ɂy��q �ɟ�Q�%2��� ��B	K ��!`6�R��R1"O`�C��	���T�5.{X���"O���!V;s��
� Z�����"O� ���ñ^�8���BX���"Oe*����ݠtM˱}9^H�p"O}�D��lFٱua�;��ػ�'P�i��\d��xb� �Ȕ�'D�tC���-n2T�FF*m��}(	�'v��k�Ƒ� 2��D��:�}Q�'4� ɷ�H
P�IiC�Ւ+'���
�'#H���kR�>���We�?8ɸ<a�'W��P�Ϭbe|T��`�78���`�'Ph��jӟ��E���1��	�'�� +��֒6�Be�1�F "��H��'Ҡ8X!��Ow�|1�˗�
܌z
�'n�9��Up
*��+���4���'������ ��ؐ�W
m80H�'�@�4+��w�[	�� 	�'?�%qaH�"�ĲƤ�/�(��'Y:��HS�F���U$ 9l�$)	�'����	�8r�Ht�eAČ^�R�s�' ���u�,L�|;5������'��쉋�X95Ɯ,��9�'���څK�:�� ���W�Ys�'�NyjF�8 	���p�Z	��hc�'���	6�@](!��-�D��'ά8A�
OT�vիsO�t�����'�����j��[B�yBĕjkD|��'^t�g�������Gʠ[�N���'J��iEbֶI���˷�I0Qh��I�'��,Y���O;>LZ''��y�X
�'�68�c �*���	�FN�D�F|q�'Z�0���j�����k�.8�Jl�'�h�@Qz�H�ZǇ�1��Q�'���*�$���I
w�\;/��4�'+XPgJ
eI��+?")]b�'s����@�L*��n�f��'��0���f��=�!�7b�Ճ	�':�}
"��4lۘ��f�C���mR	�'���[F(�'z��X���M����'���Z�'L%�إ�L�lT�'�|�PJA$V0�1��I�T�l��'8����,��8�4D�Q�U X$D�
�'��TЃE.�8�[A�\Nw
��
�'�0��!���ddZ��Vf�	�'�ڄ"$�,����'D�C�4��'��d���2x���斡6���x
�'TTj��"V� �S�S ]�	�'>��S�߂5���0�bĹ{M��:	�'��們2S_Z	X�Β�py6�		�'Ơ�
2oZ�\੓̚�3���'�6�3),,��8󢍔%||�'Lp�S��Q�T�S�����y��'&$�t��2ȅB��]-�����'��)��X�;d�ㅯǠ}��Y�'fl�DΌ1ga\�zt�_ b�P�	�'�����KD�Z�Th��hZ�]82hB�'�d���G�B�Cd�ʿ@$�p�
�'�t���Ã�v�lD�3mĲAT�3	�'Ӵ���K	^���b�N�1�'H�Pe�
R���iE"��<I��'z.�3@.�=c�x�t` �
rq��'@��b3�K|�j5j�H�d�V���'☌��h@3V	��F��F0����� �܀ѯK�~���q�F>@tm	�"O���E_�x���v��;T�"O�	AE�/1j�=pp�?G5*2"OLzF��%#Tx2"jP�/�\؄"O mrU�K�;����Y�%�T{�"O^=��უ���B�X��Ţ$"Oz�Ң �7RZ2�y�a�D�`A"OX�Q�3(n�C����+�fM3�"O6}� �18����U.ìo��Tc�"OL�J̓�78��
�GY,sh��(�"O�����V~��	���Z� �""O-� �� �t�
���E�G�!�$Y:>�B!���M:dqe�b��V�!�D�C6^Ȋ.�9DH�� ����!��%~�A��aڟ*�a+"Ύ�8#!�DS&]XKBecr\��(�x�a����P�p��Q�O*>�l�5N�@�<QoZ�7)�е�U�D��e��b�<���x���B��^�Q�=둮O_�<�2�.J~	��O�rc�W�<ɷ��Gt����׆Dkv5��RO�<�Pe�*Q����Nɧ_��{�d�<�2I�5(���)���4���rBPc�<)իI�1ȅb ~��y!A�!!�#2h���M��*Ѐh��Ar!�d]�zV�i���b˼ajC��>
�!���$�����-�1�:̛���l�!�D#�=�s�4RQ1É�m�!�N�-��x�G
O���Â:�!�D��u� "hHz�ԘEݸ�!򄖗+��aC�̭#2СQ�[�7�!�$��Ny�n��C*��K�?y�!��xf!�C�,�H�K�O/8!��QKX1��ЧIgtQ{�I^6"!�$$3��p�$o�5Z���'�32!���H��-9�f�G[ �ǅ�+!�DM		"��U�@9Lb)�c��dH!��W+}2؂a�D.~D찻�㘹'�!��UO�dM���K7	*�5R��{�!�� ^(�*UJ%'<˱��4m!��Gkb-��eK*AA.�A�I,V!�$�'^�T�@�
�@:���S']8!�d��m��b�L�L7�%"��S(:!���< @�(֛T!�${cG�H5!�$G	��%vbT�nؕ@䁝�i-!�䙐P���ҶX�d�6FW8`!�$P�}����
�$@�b!��%!�)���+&+= �i�oM�e�!�H�DU�!b�.��|ﰵ��m�;,�!�d�d�j��?_ޖ�6L@�!�D?"3n�H����3ՖE�gj��p�!�;q�.�@�P�U�p�I�5v�!�WJ����Vc�:D[��!�!��lV|�3a�=?��f�79�!�6Wy�B�I�BԻr��<�!���&��!#��.t�mQ�`���!��%�*��7u��Ba�Y�7�!���^�Ӱ��aj`T�1�R�[�!���m�����6�`mrG��JN!�D@�P6�iy�j	7J����3+L!�DG�+ɼx8p��6t;~i�g��mE!�Tx"���M
G;��Hwi�%iU!�D�:�����֫.�ZUP�h��&n!�D�O�`[�n�
�A�f�B�c!�� ,��j�)����a".tV��"O����N�{���x��_�}f�}�"OΤS�,̰6�LPBA�L�$��"O�����T�8N�)҅ @�wB���R"O�e˃��~���ڇ��?��	2"OhУu�&M׌H�醰rȎ��5"O�Ր�ˀ�Z� U�� ����d"OD�J7�ڨ
�\:�F�i"OR-cP��s71jG$*� �HQ"O�L�!bN�Y��aGj��v��<B%"O��K�BГ3!~Mk�
�:B�p�Z�"O*��Tc��q'�@p���0��P�"O"p��CA��ZٳS�\�b��)�"O���+b\�T�ňB�_X��ɖ"O���b���*0ʈ*��Q&?��"Oz�!s��>I���p��	)E3�x�"O����Ĺ>:������>�-�U"O��"n�}� ��b*ǃj�
�"Ot\�W�ŝ��!�o�9a��G"Oҍ EHFt�ZT:��PIa"Oa���={�drElĂ7�:��"Oba��8j�Ό�!L�2jB���F"O"	Ju�d��,�#͊ANШi�"O����,R&N+�Y#U�NY6]˵"O�t1�+��aU��2T�D�b5���"OƍC�.�/O��X!g@$X-l�(d"O8�&m\�1�Q�U�.B��K�"Ol�ծپ?x����1L�Z8Ñ"O<d�p�O%؎ݫc�ȓ�T ے"O*�C'D�@%0R����!�	�"OPIJ#j�(*�ZsWA;?�6�*w"O��˷a嘬	Q�^[v���3"Oʉ�a�e��,�0J��|p����"O�ȅ�1 :�e�s��4yp�m�e"O
���E��U���HA 
��I "O�(؂ě"x� ���F	ޤ��"OZ�H�HR�Vxd �=��<�"O��࣋�m�6���OU.(�HY��"O�H� 	ղiLū��� 8pt	�"O�H����v�T�kF�0GkxS�"O�%�dB�5k�"�
�
�,=�1i�"O��*���o�I�c	¶tP�i�&"O� Jw��a���G�<Bx�"O��Q���Mx�L�$Gñ� Ӱ"O�%�PA�
2��@֥��5��9+g"OV�""��#㔐X���.9{��"�"O���	�y����0-
�'\�`t"O���dŊ0��i�4i��M��Q"OX��2F����T��"��<�"O1����k�q��,Y����q "O>J�P4"�\��˖�J���#"OLA�^�NĄ��@6�؈Q"O��� Tzl5�d��6�V�Z`"OLH7l�3n76�U�
ҕ�ybI̢@����B�A�TFީ�y�*J��1�Ƙ�R�)�/C��y��^�
V|���~V�e!�/��yr�J	F̎=a҅�y
�D��E_��yb��HK��ԁ�<s�x�jԃ�-�y��s�,�pEbV�k���!�g��yW�M!�]Q����4�3����yrDM��� �b��FN��yȟ9l�V�#(َt���3悗�y�oA)`df�U�_�k�P��r�ق�y
� �pbG�F�<� 3�̓wZ0��"Oܥb��4T�R�Y�F){G�|�R"OѢ��ҷe�ꀢ&ˁG�)T"Ov4�F�ˀ~ژ����G��)�"O���	   ��   �  l  �    �*  26  �A  M  �X  Od  �o  I{  9�  ��  +�  b�  ��  �  L�  ��  н  F�  ��  H�  ��  �  p�  ��  3�  v�  ��  
 �
 � � �  �) �/ "8 Q? �F M IS �Y Z  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" OTp�t%D��1k⭋�L���ctFR�<����� cE�+���+��N�<��+�7ƨS�g�s1V�85LL�<��C؇N�=Y���n R��@�<��(K> �H���"?�B����A�<Q�+٩$�2�*�%{F���**D�� P	"��)Ku�Z�5�&���+D�H��*�5s���i5.��en���(D����gR9&��J��F%�@ᆌ#D���3,�&���bf��*1b1駌.D��#�aիd�Y�(eot�zѧ>D��y��@~pH$�@���	3d2D��%%ǐGi*E�$�Vd4�;0�#�IB�����MN2D���8�HPd�<�;��"�d��M�0��l��,� GD���R���ƓiV�e�@N�(Z�b5�k�7i8)��	7r��#<�G�ω(�����<D���o�<���~�(\��`�4��y��Hj��x���ODZ�a�T9mVd��#�	c���'����$�O1ք{S+��(g恈�'�<��$m֟,z������8�[�'p*��)�E��lIb�I^0 �
�'[����ʊ#t��{�$] I&a
�'UDKfK�|���NP�FV>��	�'T%���ߔ*QD!��h>�A��'������6��^.�4�'��=��ZX�>U�`�lJ� �1�I�"|�']F�����?q�� B���8\�C�'��P�	�u��i+ M���� �'Z����ȑi��	�w-J�
��8�Y���|Re��y
�iB�L ~�B�[ `��yB�I�m��#�F���T���͸'������|� xQG�>g$eB�+�y�,g�$��U2`B&�A�%R��y���(#c���-F�,Hm�Tĝ�0?)O�Mi��O��xA3g.@!��3�"O� 
��u�^ڨ)�Č�"G:�4�q��`�O�m�%�9����Ù�J�m��'�*��/X�90��I��FmH)��'�4�Zr������l2l%zx��'�xa	�j�_��
_��x��'��1��ۃ�j��� ^#�"��˓1O@�DZ�-�j�(u�ƷVjf%���_%o�!��E��tK�Gc��A�+��џPP����C�v� ����x �%!&A^[!�DH�h���q�u��C"Vj�It���җX�nrݛ�K�}���"O� % H �:�LÕ}�"��Q"O*��s��s�~<;b*\�a��Pcd"O�\���A)=��4`�bZBI�`�"O���4���Y������J��Z`��"O���DB-+�|�f[b����6"O&�+ ���t�ܘ�/V?6{]��"O���V�L[��As���P�0#�"O"�R�C�`���� 7��UA�"O�DT�h%�9	�kBzTD��"ORv���L����	�ƋT�!򤌖���p#�6�QI����_!�D�-D�5	�cRxml�a1L�.,X!�DX�M��r�fԀ<d^��2��#!�ӵ=Ō(`#�;HO=�g�D�!�d��y���C`Hy��I\<C�!���-w26GD�EE8̣d�»<%!�� b�y@�I_�$�(S<!�D�:��8�ri� �Q�f���!�D	{A���j�X�iUQR!�D��������J���$!� ��0��3d0�#d�1Z�!�d�)h����wP%.J0�D �-,�!�dF	T��Yv�H���P��O&bp!�d[�r��3Uƀ'M��(�b�Ap!�J=��k��S�x!v�iY!�� �hm�qV`]�.C:��/w!�D3Q�����tM�]�S�Z�K!�=HP���h5w%�1h�"�}A!�$�Y:��9�Vtxb�*)�!�D�	*4��֎].9�[� �!�$Ocڄ[��D7����Av!��U䞌��K-3����"�- !�$T�,� 8��������+#��2�!�D��2q���Q�t>-ش�V .�!򄖥G^d�)GF�\A줂�
�.�!�$����"���_^� I^��!��O9�����o)pd-	�:�'$bL�'��� �I�kH.W�p�'zX�'P)Q��Y�S�1*;�}��'�(����a�XI	SC�v�Ҡ��'!�anE�`�U��B�A[2���'_������4);�����*���C�'A�A�@�P�.�����w�ܥ��'E2ͱ�%6��L[�T�3Ҥ��'i<]�c❡��%�K��	�'�ЌK�$�3�hh6E�{_`���'B��Q�Ë�L���n�5#�6���'ܵ����H��H��c�[hȻ�']�����ȃ
���Aԩ�4��'�J��"�"E��Hs�/ ��4��'��d��C��������  ���8�'���*�)�p�b]�E��!qh���'�|�Qw�X,X�� Lϧ{�(Q
��� ��[�H�>H�lu�c6L:R,�"OH���,��(��-°b~��5"O�PA�.��_�4�fc�����"O�A�⟅�ܵ����� $q3"On�3QG���L�7��<O��`���'F��'�R�'�2�'�"�'���'6��S�%�9XV�3à��3��<Bq�'<2�'�2�'���'8��'���'2��2��BU`H��N�A ����'b��'�R�'�r�'c��'*��'����U^wb�(�`E�r�^�pr�'�B�'B�'p��'aB�'���'�@�&"�0�� ���Hg(�U�']"�'�"�'���'���'m��'S~��v��K�qac� �"}ɩ��'��'��'�r�'��'wr�' �l(� w��`'ȟ-����q�'��'K��'�'�b�'���'�n��d�J/����	-PD-(�'/��'bB�'u��'���'*�'O�T�I���|#�F�| �  �'�"�'QB�'��'��'S��'���$��V�ԉ�5�U�h2�����'���'�2�'�b�'�'�B�'�p�i �=�(��&t���'?�'Zb�'���'�r�'��'1p�	��6����A��(�境�'���'oB�'_��'�"�'"�'�Fx��0Z�`�'u:�"䔇{G�'u��'G�'Tb�'�86M�O�dR-D��UC0��xIbi�r��~��Ж'��]�b>�MΛ��P���iUA�J���#SnłA��� �Oj\my��|Γ�?i$뜁HTH��O_��jg�Q��?!��O$f=:�4��q>uH����Ӷ)A�|���v!��!�!&�zc�$��ay�퓈2|-"s!Ч~!����Ɗ36n41ٴm�� �<��t�o��$�4ssWp��2�a���D�OJ��m}��� ��3��65O�Q���K:"zX�z�ś�hkDiR�3O��	+�?��f4��|��� 1hf*��������������"�D��m!S,扯iJ��d�D�z%HpU�H?1�J��?!2W���I��L̓��d��J>l�C�![��0b�k�z�����L�!�[n��b>M�1�'��h�I��h��W�4�P�����D'�@�'�I֟"~Γd��}A�l0��)����x��(͓3���K���N릙�?ͧ'tZ���	3_��B`�B�=e ͓�?����?���M��O"擙�b5��G.�$��7�	q)V-&**�O���|���?����?�Ψx�s*��h&&I�k�&���b.O��mZ<Qe�4������t�s�@�"i"U�����.?I�0��!S���Ĉɦ�(۴`P���O[T�rưi��ԛ�V����q����x�3�'�jQ9@H�=5]�0;���Ɛ'���*O���I	+v�T@��I+-èl��o�Or���O���O�i�<1��i�Ƶ���'�"� �> ��LR5.҄O�d���'��6m1�I���d榥�ݴI���Q�g���Ɂ��8\q�23��;p
|��i��䏂\f�P�N�#|��;��'q�_���6o�`X�EW�2~	�'0�'���'A2�'���#�����9�Ӫb� ]rB�O����Oj�o�J@�ڟ�ڴ���h��a�]��`��رs�H�@��|��'̛�Ot����i��	�شHP$W�9����C7yb`a�%F"MrO�@�	cy�O�R�'���Y7j��X�@�Y#�г�e�0"�'�剜�M�p�P5����O�ʧg�N�+!�2�[th���m��������H��=
�����|2��?��ð⟠7��) ��\�S��H�R@�� Ѓ���n~R�`��xX�M��+�<���{v|�T.��v�NTˆ��zL�����?���?�Ş��@Ϧ�i�hNH�
d/�bydl�*T��
�H�̟`�	:�Mk��>93�i�
�R��1�J���=*��re�`Ӥ�A|0�6M9?��Z{�n��/���PX�R�bޫ1TR<q��@�yRU�T�I�D�	ޟ��	ޟ@�O
��F��ǂ�@#�p<>��C�i�2 QG��On��O��l����睗	� ��c�/����$�{�x��ȟ�$�b>Ya�$��ϓ,(0�yF�σ!"`����	:6j��ΓfX<�2��O��kK>�*O�	�O(q�,����4�t�S�[�N*%�7�O����O�̛v/ '+�B�'<�$	%u�
�p�̔++ìI�5dOG�O���'�7��1��~y�A�%���p�����֬�	��D���]�K#1��Q���0��Q�m���S�hK� z�p�	��\���D�O:��O��D3ڧ�?��"J�70BA*W`ռ|��@唣�?�b�i�����'bFgӂ��]���X1�^����fB�>>���ʟxlZڟ$��!�����'l�������?A�B��	���)���n��(!��J5�'��i>���ܟ��	쟘�ɚxq��� n�#%�iAwj� |)ZI�'�6M��w���O`��1�)�Ot2Q��y  ��,��b�D%BB�c}JxӲ�m�)��Şq�Q��GO��̵��`���
x����\xܴ�'����'����iő|�W��qt�۔A���1와P�z���Eȟ�����<��e��4��Gy�|Ӭ�ʲ����@�x]|E�$&���`��OD�l�����d�<����M�Q��arv(яs�p���ʟu�֠�G�;�M{�O�E듶:��	2�S��� r(p@�ȍ2�Y�ǂ¯A]~a36O����O ���OZ���O��?6�ǐf��|A�#>��$ɆƎ����ӟ\3۴T��ͧ�?1��i��'1�:g���0|��!ľ"��2��'��I&�M�3���4b�<U�����ɜ:u�9d��1X�@���	�&M�-K��'��'�$���4�'+R�'�X˶�^��h�
'e)%�HI��'gR\�<#ڴp��a+���?���	
�x�.��D� �J3D�/w6�	����O�6�O��S�Ԉ��'���Ƅ_�kbd���dޠ\��Ap���&Mk��:�O�I�%�?Iuf,��$%����	Ȉ;^6�Z��̵-���D�O��D�O���ɠ<�f�i��H�A`�;/I�@7̕"B���d����'v~7!��3���ئ��c�¨>8���5@ܛo��Ԡ�L�M;ŷi��Bv�i���(>������O��'d$��r'_#K�5+�R�7<�̓���O��d�O����O����|��$�=Vd8c�FG5E������n�F���g���'X�����'��6=缾iQNה@[b�kЉp �dJ1��ۦ�ڴ�O�"��C�i��d� ߦTK�nU[��Aqc��_	��J�����&yP�Xx����O�N�?��I(Q���p� B-p9Jġ��@y��A�℅�����`L�5E�m�	�?�@\w$�!A�OX��'�R=pƠPr 	A�
�r���'�I۟�0�CQ�4�ݴ+�&�u����'�"�*&�$P�-�B�A������ء.W��c�.5�1�����9�J�$׸{�R`J��=4�AB��8>����OL�$�Of�2�'�?)��ϻʤ�׏��T�bY �$���?�`�i��Q��'��%a�>��)�ј�a��7=*D��� ��	��M�׶i�7-��6�.?� �8��G1|6�I"w���h@����jZ%��O>�-O�I�O8���O����O���J�b,�(��ư�1��g�<IշiF��D�',��'��O-B��C��@�q%�����X%K��?)����Şi��m;�AW1�~lH䮒p$CƝG`%�'�hI2�͟�J4�|rQ�D��F��BC�=��dl����4`MƟd�	ǟ�	��ry��s�`�âF�O��*�G[#�H� {���W��O�5l�S��$�I۟��	ݟ��Rm�:\�!�W�<��)���WPh�m�G~R�P=n�XG�$�wVtQ��n͠H~�� ���g�n�z�'�2�'���'JR�'b�҅O�R������B�2x�#�O�$�O`�lZ.:f���P�޴����$�� @.<��ěӢ��
~�p�x2�e�>,lz>�Bŉ�զ�'.-K� �(�Z�!w)R�u�x4b��9	��Ir��'�i>��ğ��I���D� �[B�����M��J��`�	��'(�7�v`\���O\�D�|�	�O�y�I��C>!�4L@A~bO�>��iD6m�S�)ҵ���o�@��.0BQ項�I2_KB�)ū�'�j����W����S�|����t/l�9#�.�|9����5U�B�'q��'F��dZ��۴U�FQ[�]�(A4ay��VoL��c_��?��M؛V�dDr}2�'�F�J�)�� g��	§Ǳ4+��S�'��ӇL����t�#*��8~�Ԝ~�w���J}��ě
!���4��<�,O��d�O���OR�d�O˧$�⦭A-�r���/��9Ӹi��T��'��'C�O�R�g��Ҡc�p�J?�-���A�8�*�d�OВO1���Ռg��找=P�k�'҉R/�p�T�l�ɰf)"� ��'
N1$�̔��T�']���Ӡ�����h�$�	��հ�'22�'q�]�pXߴ-I�0����?a�Z���Q!���4ls�qV\����>Q���?1K>�F��0�.4�G�T
U����P~2�J�:�7����O 8�	�y��)�
\`!r0���D��V'��y���'���'_���8�BJ�.'j��hM7��S�j����ش&ߐ����?�A�iM�O�N�1�1 ȥpMNu��B�y��$�Ц��ܴQܛ6��,[!�F����6ğ��t���p	������M[rP:��Ò|B]����	�t�I͟<J�6`@�e�B�$R�i��Wqyr~��p#A,�O��$�O������ s�0@ph%���p4LW�X��H�'+b�'�ɧ�O� ��1M�:�cV�O��mr�i+�	(1:�{��O6�O�˓8)�1b�`ץ(4T�k��� �p�`��?!��?���|�-O�toZ5N�Z��ɩ}.����m��x��%�����N��I7�M�B�>I���?i�3�D�zE�N� ����L
.Z�Mp�c�6�M�O�h�6!ͱ�(����5{�t��U�O�q7��{cN��	��d�O����O��D�ON�D%����p�q.S!L�Х�<�,���ǟ<����M�ff��|���~��֘|b�OEa���S��5N���@йt�'x����	�C�����Fћd�^� թ��!T��ᄜd��$8��<�'�?i��?	f�2v��%��ϑ�O��ٸ��4�?����$GΦ	�v(������`�OX� ć��h���4�P��<���O�q�'>7S����	4��O�<|�G�!9��á G�s{Z@��C�h�*!��;��4�fݢ�{��O��Ł��.�XT�V�C�t��E��OZ�$�O��d�O1��˓W��Fa߹%�1/�ʄ��C�!���X� �+%���'�v6�4�����Y��=��e5�*�s��պ
��@�`ѓ�M���iN9�7�i��	�,*�{W�O��g�? �"��T�[o��B�� �u�6ON��?���?)��?����)Q�MB�Tc)�+}02y"�eI<INN�o� /�"��'[�����'��7=�t��DI�'#2�)ī�'q��H�CG�)#�4�?�(O1��-��i��?z��Y&�X�n�REP���7H(扑eD�1��'2(%�8�����'W����Ď�v&&`���x�y��'h�'rS���4P�2� ��?���2��<P��^(q�	�C[�)�#��n�>Q��i��6��O��l�����f �U�����n��(�'��EG�֜<�э�D�Vݟ�ѕ�'��@��a�$x�
�%f�����'5��'�b�':�x�e�O��K����O���F	�0�N���O�O�Amڈ_�*��'��7=���O�nZ�0����
C�iu�s��Ōm��Φ�۴o��f���U�&;O���^0I�dȘ��:��`�i]�X�"VE
;(*f9QH/��<ͧ�?���?���?�q�Ǡ?�zt��Z,h�:�Zt�����꟤��+�O���O�)�V˧a$xb&\zQ���A�'$�I3�V�@�I٦��y~J~Rӄ	61ӀIЁ{��X���D'\ ��@_~beG�-�H���&>�'��	�4�`�ƞ�M���� ,�5q����	Ο<�I�,�i>��'��6m�|V��n$��FG����:%�]G��D֦��?ّT��	�@��?��(��)�w}Z�1���2�>�"v�����'D�������?I�}Z��]��I4��6=d5��-U).�tP��?y���?����?Q����OU�� O���Zq��e��Kᆄ0w�'�"�'t�7-��<��i�O��n�]�s2|��M�r��4ru��&��I$�4��Ɵ��=�"\o�p~B���DF����<T���I�M�0d�|�RET��Cu�|U��S����	ݟ� ���
���j�!��%�U�WOɟP�Ijy��w��%�d��OV�D�O�ʧi�-��AGa����/ک>���'7�꓎?�����S���a.��F�-z}�����#���˄v�>�"�O��N�?�E�/�đ�WG�sF��>��P!� �2�H�$�O ���O���i�<Ŷi����q����&J!7��X������Q�'nR�|Ә�p��O
�m=vx�y�	I
��t��&�0o@P�ٴ=��/.ݛ����q0ɍ��ė~�tnR:8���X��L�@���SN��<�+O �d�O�d�O��$�O��'W8M�@��g/@��1dE8r���inM��'9b�'�O8�hl��ٷ��)A%��:Vg��0/�*+/�uoZ1�M[�����)^2 � 7�s��ZE�:h�h�ȃF�&�m�4dc���6��=n�C�f�	Ay�O��Z�0}� K�e�")Fe!�n	�3b�'��'��	�M;�Gؔ�?!���?a���- ��+�F� ڢ�[Cb�<��'�j�`�V@qӊl'��@��;����
�&Ԭɑ�&(?iAD�h����!IO|�'e����M��?�&jF�ErT���Ӓ���T!��?)���?9���?����O���T �a3���e +k��+���O�ElZ)���I�d�ٴ���y�Ob�PZU�K�"���*��y2�'b�'+J�#u�it�		(���Og�Ik�E�� �+q'�� ��p���t��Uy�OqB�'��'���&(,��C��=�����P�}�6�M�1�ƍ�?Q��?�O~Z�8������sa%��4d�ذK&_������0'�b>����ɔt~H�ڱ��'���Y�('~��1KG�2?a��[�F���������DB�J���O��Uk�jQ�|4����O|���OP�4�0�A��+T�?��gD0�<�c�'Z���a�"�?I��id�O`��'�B�'0r��> Ra�E�u���3�(B�NHI�i<�I�g��V�OMq����W<�tP�q�{Հ pl�S=Ov���O����O"��O��?��F�ƬYE��
�lؔI2�Pb��Ο������4FO��ͧ�?q �i}�'p�rɏ�{�����ܚ(#z,HE'!�D������|z��C��M��O� �#��}�#�I�B����Q$N8�����7R��O���|b���?��OƚM�Ѫ
T�*0� �$v�����?q/O��lZ%̤�������Q�T�ռ>$V��`�//~Z�KԌ����d�^}��h�ʰn�ʟ�ҋ���!d ,�� �#t2�]�sÍ�A�AJ ��Y��O�)��f7����\p� )dϊ�_m���ω<Z�,����?���?��S�'���ͦ� �e��q��C����ܙ���r�q�	���Cش��'H2�`盦�ԫJ�Zs��4fP*��5s�N7mɦ1�Ŋ�˦U�'HhX����?��V�_]������VӚ�z�;O�˓�?��?���?Y���	T8q��E;���j��)�F4e�n�)i�P�I؟���i�؟4���{��<2�6@�p%uF��1�`B�'��Fu�8�%�b>���h�æ͓i#��X'�J�D�B�M�+h�\ϓw��5�D��O�عJ>�,O��O�`U�j���$ȍ/Cg2LX
�O,�D�O@��<��i
h$�'6B�'���i*ϓO1����BV�6y�Y����p}ho�"dmڊ��j���0�%?PۀU(�Ӟ%���'��� �Ҩ&��������꟤�Q�'?��(tK�B�̑D��&�����'/r�'"�'w�>��	�~9c��Ñ+,��b+Ʃpgz�I:�M[���?)��x3��4���%@_1����D�y63�;Ot���OP���\��6M6?I���Ê�3� �� �Ip� 1�RkW0J��B�8��<ͧ�?A��?���?9E�ˑF0 ���A#\f�iӢ��#��$N֦���i[֟����x%?��	2�4 ���� ��Ѓ����٩O�D�O�O1��u�х� 7Gx�2$gˋp,U��B	}�t6�>?�T�3$��IO��Gy�#�q��Kڸ{N��EF� 
h��'���'s�O�剘�M[aI��?1�.G�����"��X��ᱦ�Zn#�M��Rc�>��i��6m�����E�*-6��y���W�V�pb�"^��o�|~��¦il:d��Hܧ����n�-�|�A�_�4�R�hu�@�<����?����?y���?i����%}:��c�Q�`��C���'Y���'*�ds�.�6;�����9%���&��]�2�BT.B�_�p��.�ēj���!t��iK]�7-4?��C�Ȯ|*��إ:��sS��+\�����O�]�K>9)O���OF���O �CC�z䠑C�oP(8�^��b�O��D�<	��i���(�T�<��J�d�ߎ�b]�.�$$ yK�NQ���t}��'���|ʟ����Ż��Q#a
��������!��4��i>��C�'cDI%����g%x,�hi�(]�J+E�,��(�Iџ`��ӟb>�'��6����
�apN�GԼ���AJ���A
���Of�d��i�?�vZ�Ԉ�4j�2�)�@_f�	�$ś�Q\:0�!�i!6�Q���7M)?)��Hg��I9����7쨐4ş m�R���yBQ���	۟��I՟4����̔O�ٹE��?v,,� ���g�c���)��=B�'$���T�'��6=���C��.)�B�H��d�"������4�?q-O1��i�Э{�4�	N;浂�gS�� R�ŏh@�	*(�z�hV�'\Z�$�����d�'aP�%�T+ֲXA@�C3�y�t�'h�'�W��4DԮ$`��?��c��͊f�K$v�$���gƣ��9:���>�E�i��7m�O"�l6���T�^ a��㣤zqk�&?9�Z�w;�E�Ӣ`�'g8�����?����B#�uL�)`�|�*����?���?)��?�����O�\{P��4.���i֭��$�t'�O�a�$��)�O������?ͻLD-���B�&�**��9�KM�fnq������`�7m/?���*;���iҲ@_P�`u�.Ȟ ps%�!,D��L>a+O���O����O<�D�OX�*�ԟV��{��5r�ک��<9�iG����'k�'��Oj� ơs[8�Q�E�8� U@t"כ�B�:-��Mp�P�DVH�OS�Ag�� �А���/`"Y�s�T5���O4D�P��?�O#���<��̦Nô��P�G2an�q���� �?����?����?�'���ʦ-��I@П���"�H�(P�m�ip�!���]����4��'"��?��4�?��3m��Ӑ�E@�t% 7��9,$�{ܴ��$�]�.� �'ȸO��س|����V� S\�atMV��y�'�"�'��'>��	J%^���9_�T����ɾ3�es&�'�2�'��$L�����'6v7-:�dɝ0�x(5���K ���n���O����O��A-472?Ir�
r��2�c�Nsh �C�K�@�	�0G�O���L>�(O���OF�d�OJ9����+�(	Ml��-yb��OP�$�<Aװiߎ�Y�Z����s�4��(m����MY-wU�x`Q�����v}R�'�b�|ʟ�h���w,�qq6��(dh2���i�"b��i>y���'�fu'���G(.tj�t�o�7'�2H��\؟��	ğ8���b>E�'p7m�G�J	X4 ذ;�@��v��6X��p���O��Dۦ��?Y�W���I4K��݋�j˴(���0���'c!�E����$�Cڦ1�'�b��Js�'D����RIF�1>!���D���͓���O��d�O2��Oh�d�|��"�3C��a"�
�8�HU���m����L���'�R����'.�6=�8���.@�҈��lK�3��}�gD�Oz�$,��)��u�&7�~�T�e�0�z�h�/��lYM�6Is�T��Gv��D2�ĥ<�'�?A�탏6���ff*q��?����?����DC�=rE+�� �	, �mͬxf 87�&#1Qy7�B��v��ɴ�MS�i��O�� ͘�R����v,V�/K������S��X?<<�ʓ$�S�?4����,�f��0m�|���[2N���������	����	ʟ�%?%+Dџ$�	�x*vIX�NvX�=�b�A�>��I��Mc&���?��.����'m�I���]�\ߎ:����d��9j�+N�;5牉�M��i��n�W�v��j�
�:3�d��'�2��$KM�F:<a5&=Q��'�4����'32�'���'4��{���	кq� M\� ��e�2Q����4ix �-O��d;�I�OZp`3�ʃ1P�H�!�%@(U��RC}RabӸTn��Tj��	��LCP�䎟�b���A�f��m�A^��3
2�UpG�'���'�@�'���� E��^�N§<m
�E�$�' ��'�����W�r�4H^�p�g�m26"��C��ȵwj`z��9қ��D�p}��'o��'�ҹ��\�PȎ��&[=i�Beɴ�SJ����P� �0t����i��Q
��Z����vL�|�j!p7O����Or���O����O:�?�8pg� ÖDi��W�ps ȴ�ʟ�Iן�;�4T�̧�?Aǿi��'�4th�������C͛�+R�|x�|�'��O��D���i��!MZ� h�S�͋?�&-�$J�4i�BX1b���?�SO2��<ͧ�?����?�CB?
"K�눜5��ۭ�?��������j���ğd��ٟ�O��ep���'j��}�����Od��'k��',ɧ��&)r*p��lX2�����ϒ_�a G�>�8%�є��2/y���U��-�X�K���J��32ʞ�U�������������)�cy�	k�Z�s��
�|�%�E����Ǧ��zܶ���O>�np���I��`�fFX�yT��ˣ$�y���rƟ��I�)�nP~c��~��$�}�䊈�SQ�Am�}[�/�<1(O���Op��O���O�'����f�}@4�X���7�,1�i�� ���'���'	�O��	��?����APJ��ĩ����/�j�oZ#�M3��x��tƖ��F0O�x�b��1V�����4U��� ;O#d�ˉ�?�S%8��<�'�?�e�؝0*p+A�^�j�"��Q��?���?i���ăݟ�E�<���F@�qcl��fhp�c4P�0�T���T}�xӒLn��ēVy��"�ۼw 0�V�A����'�@��*C�L]k��ןk��'֜���N;c+}��F�4'?����'X2�'[r�'��>Q������Gʋ�|�!3�z`�X�I:�M{�܏�?��� ���4�<J�ܷ;?��J�4l�%C�6O�to	�M���	D �ߴ���K�?m�)s�'q�(r� ��~@؆c^7l2ȸC+�$�<�'�?I��?y��?Q@��l�H=1�Oo���'�������;#������I�<%?���S)j�[` �qH6d�f��=K:�(�-O��z���d9?%?U+#*���h�Hӣ��(�R���mY�z�D�{`�0?Qc	�2(���!����Z�s��C��8O E�\H�@0���?���?	��|�-O�]lZ:b]"H�ɼ�na ��ތ�(��E�8���I��M��� �>�ֻi8�6��O���ɞ|Zd�� �T�kM�n�R6M=?IP���'�J�	<��ߩ*aMV�S�r`��eۙG�R�h{����ß���䟜����T��KI�Y��ӄM�0cҰ@��.�?����?a׵i��۝O�2"y�ГO^	ېه"�z[��س�˩g�N�O���O�Ɋ_>7� ?q%�F
zGH�b�B7Vs޴��`�8X�P%�g䴟�&�엧���'���'�F���KCX �yE��┴!��'��T�0cش Tf@C��?����N�BԎ,�Z4�xh��ϡP_�I����Oh��)��?�r�kƔp��4CC��Cv��=Ir��4C�r?T7�3?ͧ8S���J��?����УQ6&Q)�Ө/�6��	ܟ8�����)�vy�gӘ�a���Y�ȑs�ԬRu�-���;M����O(�n�v��V��	Οԃ��h�Xˣ�H�	T�X��Aݟ8��+���mZz~�@��3���}�q׏Q�f�3C�>��@��l��<9-O��$�OR���O����O��'z
��sJ�z�(1���ߐ1�6Mc��i��e�s�'2��' �O3��~�󎏱V���O0pyUxЭ^>.�8�d�O�O1����E�s����G�L�FG؟>�,,[h��#&�	�hZ���s�O6�O���|��P��y��_���Q�N�r�������?���?�/O�]m�!D*p������	� p�@�Ą�� ��EG(�q�?��Y����ܟ &������2�8h#E�b9� � .(?�F̏(�ڈPߴ��O[ ����?i�#�W�(Y8פR�.	�7���?����?���?�����O��`�X*���Ai���#�OԽo�6xc*A�������4���y	��s����$��E�Q	G��?�y��'�B�'mM���iW�I!Dz��b�ߟd�����'U2H���U_њ�A�k6��<ͧ�?���?���?a��6J
�@	J������Č����&d]؟��	�<%?����Tmi⭙6n��:gO�/S�*�O4�l�M�u�x��D$��rq�殛_P��{��W_���*�!�9���W�`��M��ypޓO��e^���Æ��L	�E�D�q{�����?Q���?Q��|�/O	n�y�V �ɨ|HF�cuo�4B��@��F<%�&��ɑ�M��⏵>����?1��I��q(ǩ�$�����ݝAР�;��F�M�OA$�>����d�w(^�A2��b���[夋�])�,��'�r�'"�'b��'�����sB'�r��,�6�$�TA�O8���OZ�lZ�a�(�S� �ܴ��oK��0�����Te�'$�HH�N>���?�'?�Q	۴����
"T�s�'�r/��(!�����5"��p����r�oy�O���'��,Ț �^iH�G�`A��c�~���'��I��M��l��?I���?�)�ڍ{h˒3"8*��[�do�Y嗟���O���O��O�S�?��`J����2�x��&�
�wϔ��cm?0(�m(3�1?ͧuaZ�$���U�D0�E\B���Yc��s��p���?	���?!�Ş��P����'� Z!�%�	NA���04ꐦq1@ �	�0�ܴ��'5�=�V�H��]��j��#�����;9��6-��I
�ƦI�'����K��?U��\\!�`��,�h��b <��J0;O��?���?i���?9���@$#�\I�(�;�XU#1"�?n�T\o�h� ��I����A�� y������i���5J�Hׄ�h�#?9�b�i�D�O�O�K¿iL�� �19G��˼���@/UҐ#�1O \`�L؝�?��-��<�'�?�aO�j�Nđ�տI�qP��W�?����?����d��͹��_vy��'�䣢��=[Z$j��Аr����Dj}��v�v�lZ蟌�'�v�2`����,�Z��޸�O>}�2��8	 ��!��ϝ�?q!c�O��ґ�օ�����(�3@��Ă��OX���O&�D�O�}b��:*���B��;�Ҭ���ӑzO�L(��8�f�u\B�'�v6/�i�%zRȇ�?�峆�:\?PX�6N����I����I����o�c~W�t���'�V�:`�߭�T`���,�f�|�[���� �I�\�������5S]FqE�ׂz�����+�yy�}������O����O�����D�%�{l�"ZQ�)ZD����V��'��e��6��D�K�OX�p�@/P�Dj�H�o= �'&h'X	�&'?i��,_�B��N����ε_Yv0��&g�-I�J����O��D�OL�4��n�fÔ�r���62��`��("���D���Rjm��pЫO���O��RT8�3��e;ƈɢ�J�|kP�:%m�:�*9R�!De���>U��6[����E�dd仃�'K�v����I����d�IO�'h�H�s�4W�d	���Dh|���?����K�����'�7�&�dU�WlV=��	M)^� 9��^9�^�O����O�)ϣ��7M.?IU�� gL-0�a�%�Z,&�	s&Z�
p��������4���d�OD�D�/!&�`aJ�n��  �D�OAF�$�O˓_����"�'�R>1c��W0����I�'ʰa��+?��\���	۟t%���jX	t��#b���[���5I�&�8�����A�E��P~�O3J��!��'�����J�?��)b�& 4��Z��'�r�'	����O-�	5�MT%s�b�I�e�:R~݉c��]�ru!��?	4�iy�OpH�'���Тy�R�� E�v+���0J�'�DQ�i��ɤ�Tq�e�O��'�)�&�67i����A�l�����Ov���O����OJ�d�|�7���k�")�dH�Z�|x�Aͽl5�Ҳ�?���?��'��-���4�@*N�N\D ���Ѽ@݀U9F����۴�?y,O������D �T�r7�t��
��ѳr������ҝls�H�Re�(+�iۑ_[���d�Py�O��bZ��\��DL�
��ъ�<
b�'hB�'��	��M��E&�?i��?#�"&�y
���<M�=K1�̂��'����?	���CH���#/��nd~�c@��!5�'�ȼR'N�M���$ş0�g�'f"��a�ەf�؊�M 
D�����'L��'��'L�>���[&���g��0�=[�=4l.��	��M�� ���?���M��6�4�\m[��N���o_�	c )�:O��mڱ�M���i���"V�i���>D��X��O_��H�L�
����T"eF�d`�F�L��My�OU��'y"�'}�D� -���`֔>Ϭ9�E),b�	��M�T�@��?!���?AH~*��`�Y�� "
_ ��&퇗Q�^���P����4=Лv
6���^-Gk��fkG�c�	F R+D$�Ae�I��8��'��$�0�'h����"��_�]��m�>a���2�'`R�'�B���W��*�46�B\Q�x���S��ƺ/��a�%�N�<ˬ0�������D�cy�'ɛ��'���;�
E���qf� �ֈ� ��O<����$ZCc*&��4�	����V�$^�)$+�%�4��3O<���O���OB��O��?�- %i�&  " 	��!*�-��L�	ß��4H*��'�?�U�i>�'|*�ã��pi�ïԨa��	���2��5h��|*-���M;�O�T"`��4'^�0�A��5[��T*Q��I3��Df�O���|���?9�b<�0E�X�g0	�c�My��s�)��?�)Oj�l��tll�'#��O.wBP�k�~�@S	����(Pv�M��y��'Jʓ�?�4�?Y�O�T�O�����%>5�N�W�Xi0���8SƬj��5������i��f���O\qr"��V8\�y+J7�țc��O>���O\�d�O�)�|�(O ioZ6z����1��T��@B�#gԅ��[ʟT�I�ML>ͧB��	䦽��ί~O�Ɇ͈-H��h2ߛ�M���_�n��4�y��'��e1DD��?E��O8e�AK��0�1E�nh��E1O�ʓ�?I��?����?���ή;=jl*'��#Rٰ	�$�?b���oZ��Fy�	��H��\�S���k���C�)��_�j��&�P-Y�:��7 H+�?����S�'!�D�ڴ�yb��*�$�\��:M�p*ۭ�y�N�$	����I��'��i>��(@��Ȓ�R%J���+5l�HJn��I��|�I�4�'�(6m�8@�|���O[n�a�(ʔi�-)�X;B� %t��?)�U������x'�tq�F�a�A�L�*��y��h7?���{��(�ݴ��O�>A��?iì��Wu�� ���h�R�jL�?A���?q���?Q����O�(�
�-[�6劰ƦZ��VO�O^�oڄt������4���yG���]�:H�@G[�R�	��Ǐ�y��c�haoǟ��A+��-�'R���G�?��ue�[԰�1���b�X*�iV�'g�i>��	��0�	����(��� ���$Ϟ[Nŕ',�6킜x����OD�� ���O`1r��ãF�$ ���MZ��S'Ag}��'��|������� ����+K-��y�QfԊqD��U%��;�I���h�
Ժk��'��	��}�P0�є7r 6 ړh;�;uj�O������8�rAl,X����O��	Yº�$���K%��T��d�1`�����+�
���?1(O��$ Af����MC�4ӿ�,LR��8�#Ś�����@hT��4�y��'�D��g��?1q�O��I��f��Q�C-O��V�]T�Y�2O:�$�OV���OX�d�O��?]�ş"-$�A�.�)���C�Dş���ߟ��4j���̧�?Y��i��'&�1�V���WFލ��@A���9!�|��'-�O�R�qƽi��		h�I��M-D��*��G�x���0�e� +D��n�ay�O�2�'����^�4}A���)*I���EG�e���'����MkD

��?A���?�*�Zuy�`�-*�l�k�#�3X'��c1��<b�O���On�O�ӋH�A �����Eƫ\'l���< hͲa�)?�'p(��Ó��c�pB0g(z(!Uk]������?����?��S�'��]ӦE�i��W�)�׎B�'�jl���G�E�$%�	L�ڴ��'�ꓶ?�C��F�;���O�p�EG �?��>\8�ش��d��д)��,�Vh��j���7��ub�	��O�]6 ݮ�f���X"��9��i�z?�*��= �ԕ�
��S�^�Ag�L�D�ڨ�U�޷K�*蹑f֮hZ$(*��Uiԙ{�kēZ)
W��d��\�9�I�[~�����]ڳ�]�J�Αj�āef��POӠ7��5h�|d8�� ��l�2�Z�V��1*�Ē��jWdFc��$����m��x��M�|Q^dѦ.J�b}x)��̈́=��$*�fCw���J��q*�<8C�H�&���3�0U��`�W�M����
.;67M�O����O�	f��L�"]�� �[~�H�Z��i/�a���S㟐g�ޜ(�J8�S'" ��xg)���M���?Y�Yl�a�c�x��'2��O~e�s�V&��ٓ��xG�M��^n�1O����O��Ή'��i	�b�ib���d�;]��)mZ��L��h����?�������l�ml���!
)!���C�#�I}�J��'L��'c2U��n�-��$z&�V�t9B̒�F"��)�J<����?QM>�-O��V T�.dQQ��[���g-]rM1O��D�O0�Ģ<�C�յ �N��n@ɘ��YkB���R�	�l�I[�Iky� �����jx���Cg���9�.j��	۟��IğT�'��Y4�n�����3|~�� `��*�Vm���'���'r��}B H	lg�XC�̎����Ĥ_��M���?�*O�TA��v�؟��Sl��b6iId�)� #�).ij,�4��d�<�E�z��O�iR,�'�Z�ެ�q� �{/�R�4�򄕴#��oZ-��I�O��Ɂ}~� ؒn�lH�b�O�E셀�	�'�MS*OZP�A�)��}�v�[BɈ�G�,L���d87��QJ�m� �	؟��� �ē�?���B���R�X�L��&��'~���cD�O>u�I !9�=�T��7V�t�E%ـ,�z|��4�?���?Y$ �~�O�䦟;b=@�r��6K� ��0ţ(�I�s�>c���	� �I�=*̸��D�&�8Q ri
�j�#�4�?��$]'nC�'/"�'�ɧ5�� Q�xY�BB� ;�Q�XQ�n�@����<	���?�����DA�=�4ȡ1/��:W�w+ qۨ=� KZ\����P��|�@y�"�b��!ԭ�#XT�Q­���¹R�y��'�"�'��	� �<x�O�5#�K1�}"�_2��4����O��Ox���O|$#�M������$8H!���˞� ���>A���?���� 3Ѥp�Oz���OZl���DT�i���{�h��1Ū6m�OҒO��D�O\���2�I'C$~��R�0 ˼���N1}@7��OF�D�<iD`�!f<����I�?������es�.��#�z<pD��ē�?q��h�
y��՟H4!�MX�R��j�B�3k��ї�i�I�D,��B�4�?	��?��'?k�i�Պe��� ۆ�C�$��� Hg�n�$�O�����FܧP�*E�D��"��u���8��@mZ�Z��4�ش�?����?)��B�	myB*B'@%xc�� 4�� r�R�d6&|1������Hq"���E.�W垛4�\)8��i��'����o�����O��ɦ>F�T��
����[fB�o^�6-�$U��	=�]�J|:���?��#m쨑С3t �m3.S���x���i���=mn����$�O�ʓ�?��'�\��!����w��3�||�',(t	��'8a�':R�'�S�(�uX�`m���-E*N��5�2�C�y���OX��?�L>a���?�&�P�}�z�j��͐����Rc���)�O>��?A���DR�frđ�'$ XA�MW�>���� ���9oZAy�'��'��'������On!�u���m���aD$H`�Q���������Wy�a�;Ԋꧭ?�u�V�gn�Lq7��'Lu�/��C���'��'���'������$Αb@��Ť �1��]�	���'�"R����H����O��d���M��A9:ĸ@H��;w�C�ECD�	ן��I�y,9�?��OEF�{5,�e40;� Y�`��!��4���ɂoZ̟��I����S������ڄC����SG��_�Ɲ�гi�b�'��f�'��K�O��>�z�eΨ�&��eK�U�,8��q�Z]k�Ħ�����I�?}��O��6s� ��0�#w0�c�d��Lܚ��i�B0f�'�d1��O��?���_v���j�aq���6SH��j۴�?I���?I�̀�,n�����'Z�DZ>Pg(�lO{`8A�ܔmW���'�'����<���?���Pg�"F�%fT`�F�*���a��iPR�M�
�O��O�O����֒C}�7�/[�qe�3���?qK>�����O,$Pӂ��0�{1��ꁢB�,jʓ�?�����'���O�4X�)ɹ��2��.��LX��iT��y��'x��џ�{�A�J�$ϕ�k�� @���;@ޘ�r��֦��Iџ�?!���d�$�נpGJ}���; Mxѣ��U���?�.O���Fu�˧�?aNܘK|�0�t �'��17-�9tЛf�$�O��a�&�0� ��D�`��
�.`lU��m}�h��<	��?��Q�/�`���O>���d,8�H'tB8���+����W�x�'5�	�X��"<��9���)C��a��=��M�M�x��'�!l�"�'g��?)��u��g+DY&ŭu;�=Ӓ�0�M[��?A��E-�L��<�~A
�9Ox h&�Ļa�a�,NɦepϪ�MC���?������x�O9́�b$ުD���V��;)��ؑƪd�:EA�O���<)J~�'⽪1�C��K�/S 4"B�gӎ��O�d�lE
�S�$�>�CjW�3�`0A�����n�#��.G[1Or$R�G\Q�ş�I���ʒ�Ѳ3���RA�W�:5��J˅�MS�H�	�֚x�O��|ZwX��*�k�\C���9	7�<{�O$��Od��?)��?�)O,��Fc"p,���C�-P0��۵ �4V,&���	쟠$���'�Tx"#h�T�IB���:F��) �!��W��I֟@�	^yb斦���W�0�8M��H�F!�T�ӵz,���?������D�7��t')��E8\
 ���"Ğc�,��'`�'grQ�AeD���'DJr9jcf2Xq�Da��[;Ph�a�i-2[�D��My¯]��ғ~"�d��`�4� ��V�%C0qAe����	��Ж'�i`��,�I�O���ƜT2C� \�0)�� V�Jndht�xb_���QdҟT&?9�'Q�V�)c���Vw����m���`�T�n��t�4�ij꧃?���=`�I.��ԑ�[�
+��S�O)_�7ͽ<`���?��������4��ٻ$NA
]��a�c0�(amZ4_i��S�4�?���?���)����^=�0H�pLW�o�D{��	|*�7���s0���O<˓���<���jd�b���S���@���0���in��'�뒱YV���D�O��	.B^��!�����f��$8{�6�+��Gy5�?Q��ٟ\�ɗ6����T5QB�����,Edhcش�?I������ty��'
������
*�2����Y�N8" �^$�	*��ϓ�?)��?A���?!(O"�����+"�v8d���'��8 �]?sξ��'�I�0�'b�'���$ �i����	�0�b �$ē�'���'��'��_��E3���$�yw�����J��������M�+O���<����?���u$��'��U�g"<8�5�Ee� 4��4�?I��?�����3�J��O�Zc�.5��X>RΈz�M�d��h �4�?Q/O�d�OZ��$_C�D1}B/�&kVU;���
�z��EA��M���?Y)O2TQg�S�4�'���O[����lŹ'���#�&���
v��>����?i�z�a����?a�6f��W���9v/[)bx�Y4�q�����;�i ��'���O_��Ӻ�IV(V咡��M��[u����	򟨹�h���I�ܸ��a�'L:2���	x���:��A9>Z�yl�a�|9�4�?9��?��S$��Cyb��~�D�fk��d &㏊=��7M���d�Of���O��JT�^�.�
�|	�����?�7��OP��O �1��P|}Z���	e?	W�k&�����{P�|d���&�K��m���?���?1��Хj!�}��-�	O�=ȃH�tӛF�'a�d3��>/O �d�<���5#R/�(-j�W
`�qI�Gr}"H˺�y"�'���'���'��I�&h�]���p^�K��<�Xcߛ���<����$�O����O���*T�1��dA��;�N8t��:#���OR���Of�$�O�ʓ{>�Yh�>��jrO�az��1oP�}���iE�IП��'D2�'@bNM��y��l�^!�fA���'��Q(7��O��D�O$�ģ<�NȠ,���ş���a(��L�Ht~4a��L��M3����OH���O�K�=O��'����/	i,ΈA���._���4�?)�����4{���Ok��'����*.����ǃTf(PZB�Q�C\�듞?9���?����<������?��ciۘ<��Y���ߔu�T�Rf�y�.˓c�����i���'�r�O�T�Ӻ��`��[E�"0�� �X�Zu���	��០���v���'y��cq��K�Sf:�#��r��q�FG�uD���[�v�~6��O��D�O��	 O}"]�p2C��CNpAC&)S�T+M�aJ��M� �<���?�Tlɠ��OX����s,��3Qo�y�cR8\N6��O����O�Ȁ�I}W����m?���^�*ђ��(a|����Ȧ��	ey��&�yʟ����O���^C� "�.���!±o�0�<�oןd��O������<������Ok� L�� ݜ`�r��3�ڟ&G��F_���u@c�<������T��Sy� ){�j$҃�!'=�RU拥5N��w��>�)O^���<���?q�xi�E �,�v���i��D,Q�L��F��<)��?!S;�?I���QW�ͧqr|���Vmƴ� �d�
���o�My��'P��͟����0Zs*}����X�Mۺ�a����q��厴����rH����O�˓Ur%�����`<!m>$賆+Q7z)i�,��0�6��O��Ob���OxuRw��O��'20+eg�+e 0x���A{
ŀ۴�?	����@-H�&>�	�?q+U��1a�*H�U�J�Ks�%�ē�?� �v�̓�������zZ4� �F�Z7b��,��M�+O��RK�Ԧ�������A�'���\�Na�,�t.[���L�ݴ�?!��,x�Fx��	[ #����#C��Rz��4!UY��6g�9�b6M�O���OF�I�L����ĀYL>�p����3��Q�7O�?�MK��޶�?�O>�����'G0�
5��6�-��m��T�j�����O��ۡ�ZY%���I���_d��PgA�)�V�2������io�R� ���)r���?�&<f8+�!��$L<}��#зʡ���i����0/"zb����L�i�M.�z�;�ٔ.3@���n@�� �7��������OX���O�˓`�f0�FY�K�&�d�ѓR���� Om�'���'��'���'�h+R-��-� ���+�'jt`9[`�����Z���I�'?�5I����� H'3��qԩZf��%�1�ē�?�-O8�d�O��$ոc;�S�G��	DGtTXM��Gr���?i���?�+Oȝ��k�S7s'���1�W4R�
y� GQr޴�?N>���?�����?L�|��%�,:DRرR���<0"�r�����O(�r4}�%����'���$��+�a�1ǜ�v1�X���-Mp�O`���O��T2O�O��SY�m�� b�a!���"U��6��<��C�+���~"���z՞�����A�>�j���/8E����}Ӛ���O2��'��O��O��>��,7`�L�i��ӿvo�	�2%}�P��lL馭��۟H��?m2�}�,ǀ- H���M$��dS��xZ�7�L� ���d1�$$�Sןx ��o����5!أ85r|Qu �
�M����?Y�'�Ą�v�x��'>2�Oj�J���(��m[Dc
��cC�i��'�с׆*��O���OP=��L�T��� ��J^(hs�릁�ɔ}O�}�H<�'�(O��1�H���$�I�&�- �\8q[�4�!̈Ɵ �'��'
�T��I"�^�a¨�eF�$�P�ʳ<�53H<	��hO�$ӕ(yP!(0P#s=@����´��4�"��O.˓�?y���?�,O�MXɖ�|_2P�"BE�:>Z��r`η&N$듑?�����Op�����O ��NS���ʣh����P�Rb}��'��'�剒]���bL|����K`n�rs(�"'�-)��!J�v�'NBT��'�z�R̟�	4H�J��҉	_,#��U�b6��Oz�ī<qЄS�(��O>b�O�J�j�TH~��2��42M���f�e��˓��DC�X��3?�禹JGm
6EX���Z�5{�-���pӪ�S�Z���iI
�'�?q�����^��D�z�6����).�6m�<!4�ׂ����L<���l�h�V��]"�]�f�֦����ͳ�M;���?	��:��x"�'���Af�ʃx��@�Qb��3�^T�A eӴb%�3�i>c�4�I����#���s�&��t���j�a�ði7"�'�넥ld�y��'t��X�:ݜHaG���R�.W5�t�DxRI*�I�O
���O�t#dͫ	�.��������s�.�Ц���W\���O��O�B�'F�m#R��Y2f��z�F�3=�$� %������(��ğ��I8G�L�����Xn����-�0��W�Tş8�	hy��'�'���O�9"���"��Xtg�yC`��i[��O���O ���<1�ݎ-���87�@*TɌ�MW�+�"K9	ڛfV����Eyr�'���'��(��'a�Yx�AH |�Ij��I�y��mx�6���O��D�O��V�1�T?a�i��[��\UY����F�")8C'v���Ĩ<����?��6�|u̓��iCZEH�O{b J�"�80P@��4�?�����Dӱ]���O���'J� ��2�����ѿV�h�q0O�A$ꓴ?��?��<i+���?�#@)پm�r%��_��P
����˓n��b��i��'���OԲ�Ӻ�7��^��W�#���JA������0R�
p�4;�����.��S��1
�Jݴj��q�խ3V�7�9i��o��`��՟��?���<�dͅ�9�p�B�Yu��8�"�3xțf�[��y�|�)�OhXДˁs�
���ح(�����F���I��	�Ir4ӮO
˓�?��'�P�n !ľ]�D���j���q�4�?	,Oʔ�`9O�'s��xಆ]\�䐀1�T�7��ј@d������\�͇8fHB0���ʸ$b���?{�0��I�.���/ޠ�H���i��A��A��5"pꤋҠÆ$S^L�Q�#f��C$H�>!b<�rdǣi�q�#(Z�JP�Ȝ;���ҁ�)R���fT5.�N�)gTS0�;����uV>�C�Ɂ�D^�p��;=&9�'�W"P�����_�;1�Q���|m@�ivl��P�h!�R�f"���O�Ժ�.�O
��d>�5K��Lͮi���0V"�lɗ� ��Xy@Y	C�\t�\e���O�|k�,�b��d�q#�0[6��Tbp�S1\��>x+�ǈZ��i6�ۧ'cE�?��d�ꟴ�	]yL�Ƹ��_0�*,��C�ј'��{�ʖ��,Ii�"�,�f�i�m��x"%iӄ���ā�`�``gW)D���2O.�>�*�TV���IM�$���Rr��'$�ј%像b��AAR3
�B�'B�D�@Ѫz��"�+*T�T>U�O���VJۧf�ya����w�EQO�h���N04�#�� ���F����!1���`�# ��M"�����	�F ���OT�}��,�	���=��
T�F&Q@x���-v^�:�! ,+�@* E��HJ̅�	>�HO�$�g�׹ 6v���7/i�3��Hr}��':�T-%p0��'3��'��wpT�CG%�&�n��nʞ��u�I6P1���2�OP�3��!q1��'Ƥ�$d9\���2�D�bF@���@2l'4 �FI�O��+��������?�-��o��Ym�m�ƥ˨����O�󓭵u���$�	�c�q��'Z�?S�yz��N1t^"B�s�f�*��KY�bI8�MS��eM���'��D�0BTxI�:n��\��٭�|�`�e� ����O���OFT���?���g��\L=Z��
�:��	�f��iBR�6��+B�������[!�y2'�6U�(ظ�O�p��������L���d���W��y�,��4��l�@C! m)7GHN�V,s���?a��D%�I�s�2�b����)
�	s��g��B�	�8H4# �@�O�"mZ'/$�c����O�˓.���Q�ir�'��\�B90�����ߞ]܈`�S�'9��?��'��"ҡ�l���ߖy�JЃ��e����fą$�X�`2	@Y��LJ�']P�Z�Ŭ)r���0˘�"/:8 �*e���!Z�/�I
�)Uu�!
���L9~;r�'A�7-�O��rg;W z\0�)Ω��]��h�<����?	N>E�A��cdt�0#nR�wq�\cĎX���<�S�'	�f���=��fR�q�r�׷+6m�OEnZ�e�"˅�O���OT�ɖ�W"�d�� �ܼ8S�6H�N��,Z�+"\���O�-�'
��v�~}��fٙ6�� ��|�.�"�bŨ��/χ[Դ 8F�ݶ��
>�v�`snˢ}k�]Vn�^�O�(ybC �|ZV��@;*Jjd�M����k�O��$>�'�?a��~T�)Ѱf�/,�(\�C�\��xr��%XL��aS�!�f���$��0<9��	�qf�b�ٞ4�r0s�2;G�8��O��$�O
A�s��'D3x�$�OX���O��w�0���@ߦ_0r�iT�B�k��(y֮,f(�����.�.|1��'�B��Wʆ!<��|�!�M;=\�E���&Z����@-�O|8B0�T����nSl���(!�Mg�\�>f�x���$ܹd|�O+����4ha�E��
?�d5�s�:o!�ā4�,�%��)D�|��Lk���O�aEzʟ�2�fJs�À%�bx�2H��
�LY��
A/J��P���?I��?ac�����OR�S�3� i��$�2Dd���
��!kLA�g�>�t�4"F!>7��� '�}�l���14$�B�� <7i@Qj�1R��C��	"U��a��O6��D��� �;�	%:�b�r2d�jd!��{Z�y#���_}��  #]'1O`\�>I#�P�֛��'52MU�
�z� 7$[.5|>�C@���'��8Qs�'Zr>��a��'v�'�J�C����>d�r�ؑ�"��Ǔ1'���?�0k��`qČļ����D�|8�, pD�O0�Ode�v�S�Cv x�`m��;�"O�����F=B3���t)�)��$��O$m� ,Z��Q�M0�:�����c�Ph�@��M���?Q*���ñ��OƐ���Z-6ޑ�e!
�'�j`��Ol���-jyF �A�A�5����W>a�����Y��*�V#eo�W��< �(���J?4�L�1�L���ħ ���rt$�)�6y��Ȍю��OXi��'"�-s���*���D��fZ�P)B�9ǩ�I>�v&�d�P�b=O"���O1��d�<��KϚ>`�K���&x�-�@��T��1�O�A'��m��"2���� S�S�%�u���R *۴�?Y��?1&��9�&�����?I��?ͻ!NTj3G�)P�^��bH�K��8��y�E���<�uD^<��R���($��x�McܓW�,��I�mK�BPH�"$A�@��Q6��<� �ş�>�Ov ����!�-��i��Q�'"D���b�К7�!ˏs��R�>?���)§F�������?g�i��ڙeSpT�H�q�~��O6���O�d˺����?��O�^4�E[�Z�L8X#��D�9�����xb�Vr�? P�z�£L�\4p3"G40J��9��ZnZH�聃�(g��hD"$��d,�O4��;���WOH�-5�T*"OZU ��:g��trG)��(������FM؞d�C�R,	���	ܹaMP��':D��! /S�m.~]�O�,b�$���#$D��b�L@6\�`I�i�^�
)�("D����'�3@P�1�U'u��er��?D���p΃r��SA�fK�0` A#D��9G��g5\U�"mp��3C?D�@��Oۄ�(����/hIZ,c �;D��ʒ�����ЉrcހkH`�9��9D� �aKK"�h�`�d��#Z�Hwk<D���q���+[D�p_�$̙P<D�c&� 5>IH��ѯ��!0�,D��a��M� �!���0^��9 �*D�Xr��U�L�����B�s��$D��cbO��x���Iө!긩 Vf%D� R�����C�1d�MaC	"D�4���X�`���t��i[Z��a4D�<����k��IS6�F�����%/D�|���Ut�hT��N��F.t��2D���7��
E�H�#Ĩ�����1D���(@*���0j^/Bn�8R�9D��a&$D�dn�g^Z��	�2�6D��b�+�0�1 rH d�$;�5D����n�>O���pb5r�0�	�C?D�D�	�) ����gMȇC�:lq��>D��ѲGڡKS�A;rg���u�U=D�����&YB��5�"<[��4�<D��3a��w��-���ݑiʪA�=D�t+��F�j��.*dz(�dE^Q�<��
 4��t����-Z��2&LG�<)d"�A�|X1�˱�V� ��<���8_8�U@AK��\w���~�<A��S�f�0���(��c�|�<�#現w
�����3�|�<y@�WG�d|9�F�_:i�!Gu�<)e��$r��ջ�� ~��	CQh�<�.��f����)��@�<��d	f�<ٗh��n� ;S��k�5��jM]�<q�Nٲ���S`K�
���0F�V�<�t"j��)hr�A
p永G��O�<9c��M�H��#�/>u��DVM�<14T*xժ1�'�_a��ZFO�<!�NFO�\|���>�`	PA��o�<��ۓB�R�@/�c�܍˶nD�<�D��I��,A�,��<tcs�}�<9 ��6��H�R����{�<���b��z$�T )�(X����s�<q���"�(\��
�?�t2e�q�<9���v|ڀ��I Tg�͓ҥ�j�<�ҍL>4�4I��Z�	Ճ`C�K�<a�ǜ�uX��(oQ�������H�<ipo�2X�I�&�F�<DK�%�E�<����,���e57٢cg�<Q��hg�����>v�<=���De�<�)��]S�����0�Xa�<	�&R))FH Q�I2p�|��f^�<�g��(���F�T�f��1�H�ڟ �R@�?i�X+�<��5Sa,��D��zVC�t�P�c=�ɠ�g
8��i2+H���bX�Z��E ����yr�P4"��,Z3��&%�yX�HB���'i5�ͣlL�E�4ϟ=Wa� � �W%���" *ƃ�y
� x���N�s<�8�����<��ֽ���xG�C�d2�g?��2z߮�%Ҵf�j1�eo�^���٧H�n�|m��@�%똰���8�\����'d�2�{(8��	7����U���0l�Л&�:Gϸ�=��]kkt�ϓ&�v�	$��1j8��
$��xS���z�E ���� �,�3-E����-b�ʐ34 ߟ[��MI�>����G����ζi��?�.'1�dm�AdK�:���[�K�џ��5�)a���ͫ��ې� ���MF(�
	s,߾~�-��ӻo]d��'��iX���c��a�ꁮW�ո�E�T7D1S�d�<A��Gq@�據K(n�`�
وt�T<�@�̘S��1X%l�?A>����yܓ��=!Ai�b"�PpV�-xD<;�[��/|Ly��;Rf}#"
??9�(�~ҰB;��e�u�C.!���p`La<�0B�=�b����3��h�Q�6d$|���%�=?���2�'�<�f�v�����0i��\
-��I�vN��H!�d#�@e���\�aM��K".�U/�f��^|��6�Y12��z�Ĝ�6Ɍ ���� H� A�CΌ��= h���u��/m�<k�i�Z�$�A�'�=e�l��'�ͣ	��U��*��]h��Iy�s��݄|ߌ�J�����ŧZ9��p����ևZ��i(R�fP0p�f��{�!�dɵ.#����(̛TQ4�!ե�"g�]�6J�½KM�<�z�)��b��#}�Ji�pc̎BT��)��ÈG�!�Ǔ�܈���[>g��
��ĈtLz�\��;wF $�F�a��Y";��LGyB@�X">�����X|�Xqf�0�p=�a,%�V��2�!9�`��G:0U	����O��q5�_�:�`0r�C�0���D^�`ċ��_6"4���K)�1O$!�E�Z)m���V�X�da%J0Y<���60���O��3+^4�Q��l�.��"O4����=e���i���4t`q�sO.���2D^�&[�M1E�>�4���	:�	�~󎔄&=��K��� |�l��FI�Bn!��4l-�r�⃤#�����Y/x� h�V"^"".hx� 
,a����6(��$0%�2�	����a�(����]/\������-J�٬S&��R�G�h�Ґ8�j�\ ���J�1��=�"�#,�}���b؞�"�".�@`�GΚq��{��3�ɘu��; ��*6�2ᐕ61��� �G8<� _w% �K�?*E>9����4o��p��'͸���ֽ��!�Bτ2�^1�T��<M�~���FO��M*��M����&�	�)b��N�9(u���T8:T;��Z8Q�!�d
�%b���c���ޘw-�$����*G8l��9$���1W���Cj�{-r��bc�S�l.<Rf���:.Ψ{'T*�b���Ioĝ˓*�D9V�bw�A�L-�3Ƈ�2���`���y�f�*���x�|�)�![/�=�7ǪH�nH�� ���bc�J̓w�4��cЈk`����4
�
A��^�h���3���i�a*
�Ik�9J��aJFV{�<�EO1X���H�1TVbTR��S�eT�4��P�O4Aa-V16.��M_��'q�.�ϻ2�0��4� R`V��Eݡ=�r���4
4k�,X+���HAeE?~�īQ�bÒ��#��T�V��sH@1<)2$I*��'�\Qa$
�9bC<0�d��ʽB5)�O��S�*vl���e�L��A*�-�/�`b���);�&8�`D��۳�O��;� �2wO� I��<��3f��m+�f�6H>��G�#@K���|���]�ZЈ|�������6.�ryr�J�G�a|ϊ�3@@���f&����mͶKq��K4�$T�bb�Z:^������1S>��.�r�!��#VCP��eψ�z
�B�I6i�
�p�������!�9ve��GA؍��_��0j�kF4m?��>�Yc7
b`uȮU��/I8t�p':lO0��!�.9��E)�*�>>pX��~{NP���:2��r����l��}b�0���Ӱ��3_�����/Ѭ`���@!��5\)
�i'>���O�A(�T?��+Ĺ{T�!�I�/3k\�Dk�<E��%�0>�g*�n~� ����"&ꔵ�p�ٰ?&b���O�{Zn,`�FI�O���)§�y�
ˣ�z�����1*�H�h�Ɗ��yª����㗥�f��`��	2b,ڹ��>��0k2i^-Y�!!�O���EyrE��o8��k�P$�V�� � 5�hO@"<A�
�k��}�&-ĀI��K�#�8�4����L$)RB�����D�2��$	N�����Q�	CWe^�,w2�Ⱔ�O��PE �<ɜ'54 CK#,B�T��(�ݼ�$��
�fi��?HETx�r!KX�<Qpc�@� ��`=1�,-ܮ,͓�~������um��[��� xם�E�O��������y�kլ8h
�+f�C��0C�~Y����t��!��\�0;�21N�0��ɨg���u���1ڄ��sDTQ�� d��bl�8U�>x�G"N�E� աg�	�ztLɪ���b�\�R�\�r��';�I��	�5t�����2#xl�9��4
 �SG�m�s�W���O������h��C� E�)�AP�-˝�0��l� ��5�D&4��$
�ez�4J�h� �Th��w�����b�<���(-0��9_�������$�>;�M�;'i�	�#�I�nLI��k��r�� ���Ō�d<>9�E�	C� (�%�Q������%�:�@f�E�=v��"U,ϐ[9���$Nr����!E��j��@w��f����AV�F�f�jQ	v�S>+�����F%%n�i���~Bd��2j��'�~�r�0�T�#�NM�A�D�2��B\4����V�:�A����?!�A˯N`�%ˋ�����U"[�.D<��������>a��y0"?T� i�����	4>����X��	�0�Oo�C���;�� )�����	0.��F�X��)��닎lX��w�;s@�;`l+_��Ȉ�'�M�D씪$�*���	 ��lj1M̤�yB&P�B�(�AćӔr���*>�KФA� ѡ��}���A��4�hVB@*F��`���.�OR0xA˗>����,YV�nȈOR�.x���w.X	Pz�"c埮q$��/I>o��!'A,6^���|A��9��>1Gk����!3r*�:�X�14S@�'�02Cc��xP 0t&�>z;X�3�'�\�w��%t���s֪� X$蓬^�=Ǫ}���>��$@�`��E~���o~0�Z����Z����z{������5/J��c��> �8��_��)���;+�,1s��$2B��r�,�3C�����*�3��A��a�Pc��5�T��c�J���N��ӧ��0q���'C���w'�i��(�`"O�H���!|3g�� 6�lM@Ĕ�(�bƊ�A�ؘ��'�P�%��zd��br��>����	����R�*��@��UJ�;Q���b�F	(v��#	$���R�ԃ ��\r4�F
a�a��I7�m�J<
f���O��}��j1��� ϫX���2�'��8�%o�{�(��Q�HbXt�'�*��%B��H���+��Bv���'��\��K!Q��uA3�S�1�'����招�78vЩ�.�<�@Y�'���"��1)�`HO�spR<�'�` ��@ȭ,�:��v�������'a��˴�1#�x`�H�4.���'�����k�-r��Ъu�W���$��'�����7��]cԎD �����'k���Q8w���0n��a��\��'�Y��*�	����ǕYɀݠ�'~` �C�A�aB:�SԂWޖ�X�'?D-�h��#��l ��:�H�[�'�b����~�@�z+ӟA���)�'�0�I&)7x���kT�cd�l9�' �I��f��%B��Ja#ɐ1�5�
�'�,�1EBO>>Qq��((q*t�
�'��%A`�J�jV��w��N:D�	�'l�13agX�A�li*��.@��'���)F��o�>�bw��K�Q8�'9��1��P�px�)B6�30W6���'�.���b^�w�<�e��#"�mc�'��\(��v�h{��L���K�'%��k�c:V%�ِt��?����'Mm�π�_�p����A�:4z�'�n�HP �h�T��6l �(�V�
�'��HS�.S�@��񈑩�&�p�'�HpZ��U�7��@�d�]]R|��'�@�xᦅ�B:1)G:V�ܵk�'��%�6��(<)
�J�RT����'��U��F��u�<+�GQ9IH�1��'rVI��$�~�IPT�������'�hrR ��p���HY�(��)
�'�^@�F`�~ufL�Cđ���)	�'1�$�<h����	��Z�'�z�1���C���R`� >D��x���3c!۵@Z!p�j(z0���V(��P��(A��H%#־���s��t����0H`���ͅV���S�? ��oQ�s�pAoA*P�Q"O�q��T�/, �����k���z�"OJl�p�G3l���Ǎߞy�!�0"O��4lO�y�^�ag��+0����"O:IԈԛr���9��@1%d�尢"O�I�A*�X��=sT��Di�$��"O:4��Y�C+6�k$�9Nf-:G"O�ĺ �է3 l�A��#j�M�"O��It��kZ9h��ȁgݼT#�"O�Y0s=4�#'� }��P c"O�
Ѧ�>��|�&��^�.@3 "OF}Y�� I�/��{�$�yBK�2bVhȀ&�$#�A3����y��V
4*N�A�	��2ReB���y�!M6I��}S��X����E��y�#Џ���z"�ۨ|���P̑��y�d�%Lf���#�nNXD��&D�y2��Z"|9�mLaX#Æ��y�bY�dR$�����, �C��yҀ�=@>�m�bA�n^�3�I�!�ybO��mXa��A�,^�քz����yrI�bόd�GOA�R�VU�p�9�yE}��ȳIP�PN	�ԋʷ�y�)P�MՆ�r��)JĶd@w(� �y�[��U	�mD6��c���y���8^��G5A=��م�W�y�9l@$�Iцܱ&�*���	�yª�1n�,� �A,'Z`9�	�y2n�&ƩC,��
�x8�S�S��y�e�&_P�}y%�)����R���y�֧��}*4͞�z�Z���o%�yr�F�<��hvo��[�,�P0���yR�ʾR�;�-'f3�T��EF�y" )����ύJ,Lt#6aИ�y�BOG�(� G�� G��0!s@J��y���<�$ �C �24�Y"�ǒ�y�o�*�� �f��.�B����yȒ�o-Z�ZE*�*-�ڱ�%N���yB`�WlȄҤ�U$/F죤���yB��=Zμ$9�I��.�&�#���y��
�`�9w �1Yp�p��@��yB�J�x���E�>W�= !���y\([��<c�@Č\��H��l΍�ybn��`�\����WSl!)U��yj��EDb���Id�Ii�/���xRK�vb��=N-�׋Y�A!��4W���p ߲v����N !�$Nfܰ]J`��2�T�!��Иo�nX�Ŀq'~`��G�O�!�d�./�,@�4����r�p�$�!���#\�ݸ�e��f�8���0�!�$�14Vt��Fk��PA��N-(�!�U)u�lТ.ԇt�"�Q`$�k���>��Je�N�9rM�Nur0#c%a�<���ߤ4�]R���k�# �Sx�<��O�?���4��/L�8��R-NK�<�E� Ud�H! �1����F�<4G.)�̡��!nl|`��K�<1F��V
����Rot��㨔I�<�K�c�hQɢ ёI�ƕ�%�G�<��L�\�]Ca�J��Y���Y�<ad�V�YE4�+�J�����4�XV�<Y�'�9n�d���Y# p��@L�O�<�3�#����[�u��t�z���S�?  �"ÊX	�P�a �-(̦�Ӷ"O�1��œ� �� ؗ(A",��DcV"O�mQv��jnQ�4�Y�F�D��"O����ٱW��H�hn� �h�"O��ӕ6���'B$�tc�"O�M3��6@creP2e�~����"O�i��@D,�|��r�p�"O����J�|�e�Sw�� Q�"O��h�� ��̫#'
�����"O�H���P!f����(%┴�d"O�@Id�@7-HljL 2i�zq��'f���t�H��f��C�|�r�9E�,D���	ӈ*Μ![�KW�G�X�dC=D��q�I[�riP��HH�}�F(�P�>D�<h1郮�np�զ�~+:S�<D�x��
B8��|��O9* ��F�.}"�'Ɖ��D�`�p�J(O�0�
�'�(T��� J���IT�>���'�:US��R8�(m��A�X��;�'���*�mZ�m��Iy�"ޛ!�D��'�Y��)`�MJ;$��a΁Z�<�@��#`H�
�'� L�Jԡ�)�T�<��,�0S���Yt�O�$%H�<96JݺY���C��`H\z�<���,�Ba���(��ڀi�w�<�g͕�(�` �%�8jF��ǙO�<������s�Ή$��@�G��b�<Q�C�h߄���	�zeJ�d��yRe�SU��gC�	q�0��\+�y"��_1��r�4��0-�����'kvmq�G<'-3��8*1+�'X���5�A���2�'����'I��q�f��0ɒm	;��ܱ
�'�[ ��C�
 [�䒚6q����'D I�PA���R��1��1����'B6]�BB�]b�I:F� ,� � ��HO���Ӡ��ç*��J�չC"O���'�P!n�8IQ�E� �4ط"O���-ۻg�Be�'IC�L����4"O�<�wk�9�B$;��+ 'ɚ�y��ХE���'12Zb5�ף���y�c�4�B+�-74�)2�)�yR#H�Q髥^���DS���=�yb�O�Kn�]��=u�i��$� �yb��l�*��B9�^�ȓ��?�y2�Z���˃ʏ"&���`৑.�y��380	jW�/"Ͷ�����y�F�g_$PAM1X>�
t`��x�uӘT٤��I \�bK�q"O4���j�8��uQw��q݆9�C�'6��$�	J; 4`���Mܸ�� �Vt�C�	-��8��b
��Q�م7&�b�D{����$gN����W=�DAB���yr���,�d߂U�t�`��O����A%/X��펝���c�b]i�!�P6�M�T0Z�`�gЌAV!�d
�P�jU�R��C.���W&X�O6!�$�� J(���+�c�䃻Z$!��*�\��"Ę?�������3j!�$��P^n=�[�=����#);u!�d� I���c"��TȤ̂w���u!���E��lF��J��	
:�!�$��9gB᪤�L#�z�RI6j�!�Dī���c���ā�)ĚM�!�� Ќrm�#5Gv�hv�%}�P��"O��P�m�Ľ��� I`��"Op\"� /��Yp �DFT��&"O�ab
Ù���Z�
!>���"O���`Z(4��m��-@3M:�"O@I�Ь��혽зL�c�C6"O���i��mQd�H�����"O:�ZK�%<���/����"O�=kF��,SK*�Y���c�Х��"O6���%�}lk�fA�y
�����'t�'䔄�p晽E%q�� ��y� �'ݨ��7.��"���P"�s�R��
�'�\�T�a�ظ���j� ��	�'�H��ĝcĉ��e�j`�,Q
�'`�q�*'y��9ģ\a��A�
�'Fx�iѭ_�z�d�x�Dj���	�'p��R�D_�H�1F!il^dC�'�F��yL�M�&䏰� �
�'���I@"̧NX4E��#(U��ix�'��%�M�G��yr�"��N E�
�'��ٳ����jo��a�E!,��	�'���9���>$z���eǁ:O�(y�'8�I�"kC3S:ܬp���0,�j�'�n�����#�vT���W+)�����'kέA��O���](%ڎ�b	�'k�(��S�_�rjt ��P�v�	�'2<���䝣;c�\��΀L���a�'5Z�3�O�%G 85��
-�U�'�L��b����v5xa�Ɍ"�X�
�'������ѼX(�+�Ζy� 0
�'9J�ʒOWt���i�+�:qq�'�И���Ћ&.	5�^!�@L�5�y�	����g���,-2���'�y�A�(B�qm������c���y�����|��-�x_�ͫ�����yB�O&5E
)PB��!3���E��yr�
kKbE� �4l���X�ybc\dI�Cm֬)���B[��y¡I�cŢ�[���JnL D.�y��{0�˒�L�VX`k�;�y�
*<ε��1 �dL�r�� �y�Y�n 0�F�${�JPx�e	*�yb�N!pbl8C$�!���6!ə�yюU(����-,�����ͥ�y��370Xd���O�H�
Z��y�h�C5p0�f�<s8�,`�/��y��/P�ԙ�C� kI�hR�� �y��A���Fl<~|�#v�+�y�kQ�w8�h	3�#�v�
F؅�y��G=3���$�A��E��yb��*v\�Ӑc�'
rx%�V��y��êU�샂��!y(�y$O��y���'tv�8�nX9��Sd�̄�y@�./��Xq�d��=��f���y���Nx�JVY�����G:�yR���Cv��@Y	��BPh�*�y��A��аFa-e��#0�
��y�ݶ&�^岁��%(�p4H���y��8/ĥ1)��~��E���y�gMv�6�#V��SZ��S� �y�g�5S����gnT5@L�b����y샇gҺ���͚2��\в�\-�y�
�]MLec�C�$*�(����yrM�;:��� џ'��L�����y
� �9�+�N�t[CB@����"O��{ִ[T,���˚o�rd�7"O�����ݦm��E�7��(�1"O�����+#�@�0$	�5t�E
V"O���#��?#sP,�D$	?|xV"O���7��\O��H�BL 1�a�"O؀�CkA�[��!�(@��i�c"O�YH�%Rv�r�0aօe���"O�1�Q�
�2���	q��ZB"OZ}��6X<b�mr�^1R�"O&IRa��#y��Y`�ȣ)��A�5"O�Y0&�W " ��(� ��9ä�["O\`{s�S�:��m��9���Y�"O��Zt���0O��3��
�Hz�!�"Of�۳�Ǌ�Lx ��t��"OP1Z�h0qP�z���>%�	Z"Of�{���8�^��-�*m��<�`"O�p��W?�툆��|�	I"O6�Ț,k����μ\��ٺ�"O��,Q�M.'�9*��a��"O��SH�)e4 �©��a�bZ�"Op���Z�s\��uh���m�6"O��k�6zC�q�#�\�6e܃�"Ol���E �O����7�5`�\��"Oα�m��_)А1G���.kd��"O����@&rP��g	�}q""OnT�'�Ѹ1�A�m���0!��"O�8� '��<��G5DD�z�"O���6���$-�FN�6�$��"O����ȗ�Ǫ�ф�0~y@C"O:Q�'[6@�s��ǟg�@Q�"OTAG� hIR)!Td�Z\��"O�p�u@��f|�F���P�t0�"O�DC�nˊ�#a�Q9�ĉ�2"O�,8UO҆,�Xh�&��(�2�ۃ"O��B��G!@Ld���D�;��A"O.�@��� Wt�1���%�$��"O@Y�`�B�r��2wBR�Cr��"O�e�Í�l�rD����w���"O�1i�lR�[�ؠP�T%�Z�r"OM�TȔ��Z��TDQT�4|��"O��U�ٯ|��I������:"O��r'fԎV!�����5�,݈�"O���F�8TSxU	�a�*N1�19�"O�� *C�t���b��4���"Ol��E�֧-aӂ@s4}��"O�|�p�]
�� �OM:��"O����2*.1� ޼;�h$� "O��3��.T�p�RȺf�\��"O }š��9.���1(���("O��b�J.GaM�߳<Z�S"O����j�$7��lA��?|&8=0�"O`���Ğ4v���C�Ʌz���"OV�@��S��U�����b���"O�H�be$g�j��nZ�S#0a��"O贙�읚t�Z�㤍˒��RP"O,���KϳI@>���˖�,�H�Ҷ"O ��(� c���
��
�C�vt"O�%�C΍T�|�dGa�E0"OT`3�ɾX�F�s�E�-����""O��0��B�,왳��%}����"O� !ׂ[�p7=r�  �`~~${�"OL�ve��AK� ��O��(o�H1"O����"&���w��lD8H��"O� �T�2�;3?�����2<z��b"O���DH,(*��բ�4]=����"O4�;�'��y��ًP�O4V9~�[g"O(��@"C=�� pg�gH�ݢ�"On��'�U�O*hhq�I<f<�Q� "ODi�u��0Nъ�n��X9�4Z!"Op9���+x��p#$�`(��"O�+tD�p� ��B�p	�	B�"O*�f�!s�*v�U�X����"O>�#���,Pt8��&��4�T;D"O\��FF(O<� PhS5S�F-�6"O���AL�N��q����	��a "Ox�wa�!-zb��倃���0"Oj%� ��ۚ82�˟B8C�"O�(��ǉN��i�S3�>ux�"O�E;�蒓zz�R�B��+��UU"O��zT�^?]��8�g��N͊��"O]�wi�U���QE�R� ����"Op  ���^���yc��#I��)�"Ov��$�6ըD�/Z�
0��"OtH���N3��[��}y�"Ona���ԉ(X���� �r�a�$"O�D�`�G,�� {!�ѝ?��l��"O�pH�fK{�P@���y�b9`"OR�렂ѭ+�ĥdAN2Ps���"O��dmQ����S�!���$"O2|�r�z�����F�(/w�q2"O�i3���]2�`��
�3M����"O��RA�82[�e�"�QyI��Z&"O2��שиr����Gm3<`�"O�Y8B�۔H�h9#�ϾN*X,+�"O�x;w�&�A� !�)�V"O( 0Dƛ�B1���D=)�R&"Op9z��צ���T������"O�%��d�1'��2	%�O�<1O��f�V ���$���8W�Q@�<Q�D�H��賧@�yD�+���S�<�A!�39�n����-��am�O�<y�΅/�@��a��F�8��P�<�k�+�ejӦ �}]�X8u��f�<�T�$?��Z�fT�?.5��K�g�<��΅-μ"��.��p��C�_�<����b���(юܘ]��=F�[�<j��~g֤+�(�f���ǰxC�I/S�L$x ���o>ɘʜ:%�B��:`r�Y��!d{���Z8.�pB�	#m"�9�揁1w�D�%G�quXB�_�.���A�;	�l�j#��}2nB���^T12�L�g|��h�F]�-�NB�-�Б1�#3GlV�V|$��'��U�&!�.U`!A�G�K� T��'�q�dːZ������L�I=�u9�'���Ê�G+��5%S0F�L��'��Ѐ5��V%����Q�f*�q�'��-�iD�# `�ڡn$OLp��'̴�:e��=R�j!v�ůB�$K�'U�)�ٕ��x0C:=���X�'��]����-��T�שԤ))�Ń�'���y C�E���AS���S�'�.س�J]�r��Q��b1��'8V�Kb�@[8L�n�$Q��X�'�R�R��=`O��3��ΗK�@��'z�A�$A�cnZtH�CP�J�0j�'�8�#���V�z���B�:d`	��� \yHaHG<H됭#��ݎ.i6q�q"OИZ#��"1����Co�_�J��"O~���8<��e�R�-1�g"O� �Pe�.W�,t�-ɘ4�r���"O��8 *�-\�r=��k�z�:E �"OЅ�3C�8
:tT@ ��)|g�`�"O�� ���j܈�L�]`XXF"O� "�nf�p��WI޻0�P�0"Opiq��Y <1J!`
T(�p�"O���'$ěA�l�u��6u�-��"O�Lc�/_�L��4��臻���S"O��c��~w�Y!Ѩ�.���e"O� ���{#�bc��!f�⬐�"O�M¶%�/dZ
q@Ca��w�����"O�|��L2u�����'n�\8K&"O������o�Z����Y'#���*�"O�l�E�BU�+�Q?�XE��"O�m���P�q@�*T'}3F���"O.��f��2_Ƥ��F;t�*��5"O�=8��ҳ$�Ɂ�&%!�:�!"O�	5���e�))P��z�VmAd"O��b���N�]�ׁ�J}a���N�ذ�(�U$6�+ΐz꺡��&D�\�'kX&[�����F���Q5J%D�H�X] �ɗ�P�N�:m`m#D��0)-����e���,I�FM&D��1e��P6 Mq5iD59�� �pi'D��[�k��Y�x��#%�3T�b«&D��aפ��R=��T.��X<�@�k%D���p��.Z��h�(n��&��<����Ӑ;�~�rp��J&h��CÇ.B�I,��@��G�U�@�:�\2�C�ɯ�V��
�#�`H��?���$ �S�O+ʌ�⩄�X~���럎g�@��"Oh%���&m�ikg%ٙ��P�"OfLXG*��\W`q���[���i��|"�'������OT�u{���H{v���O�⟢|��!�gy��H2A��Rg�B��Wo�<��@�L/b	jf�X.v��A(&�p�<�w���L�0���d��t٠���l�<�^�1ق$XpO��(��5Aj�<Q�X�\rh�j��;�8Y��.Xb�<1��sO���"�I Z)PQ�@^�<!e�0���"e2hC:,1c��]�<q�ړ/���J�Xc����M[�<1s��+����� �la�0��CA�<�fM���� �4=�)��Dz�<�E��>�}Àʓ�;��UB�O��M���O��M��"�/cly�A�)(�p���'_\IPB�z|�2�W>\$���'����L;f��iaG��OĴ���'�؈�Pɓ�RN�}�u��'A���	�'���ra�����T����y	�'�l�c�	ɧz}l��ģP�{Z¡�	�'��!3��T%1��0���#(�<�P)OܒO�����}�]�Kr��83�S�Q=d�9��'	�O<�}��@J���p�Q��}9��S���C����Ŏ̞<^(Q�kQ�.��p�ȓ���)W��
��X�NG�u�܅�:zHyc��9a�YF��2�l}��Q���p1AĢM���(m̙D{2�'������W�y�T��O'A��J
�'��	��R%l'0�sFN} ���
�'Sp`i���0V6m�âV�s��	���4O� �IgbHS���C���T�l�@"O�0���O]�	p���D�!"O�t���W�2>xp�"$C/b��1�u"O��5��t�@]��&<�*X�""Op���e�s�=�0V���0@7"O�D��N�����^>=�Pd"O4���l�|"� ��I��y�`�D9LO@�0!�٣*�.�j���x�t�+�"O�Y(��J� �T(�A��l�!"O�]����*3l�QƑ;B�c"O|`�g I(n2���ě\�������Od�4�O��y���^�b�h&�n��+O(�=E����p��)�
*`rL�EH���>a�O��3�T�\��A���RG:aZ��� �S���<�h�2�M�+�Lk�bE�y2!�����BJ��j��(zv!�Dˮ���'B�q}����:7u!�$ý}���ă�*`Թ���-^ў<���U�`r'%�1���ó:��B䉹A����S�(���$*�/��⟼�IU�}y�OP�R�� � o������jRu����:�$@R���"\i��!'����"OL��rL� R0�T�J=-Bذ�"O��H!�N8@2����eRPT"O0��	�#\�~�BMq)��LƼ��?q�^6�hSd�ͺ#g�C��}]F�8��x���7P �"`ң�E���T�hOD����!GL�Xu�`�� �����"OD ��P�=������'��=�$"OhU��B
�`�u8���K,�k�"O���V�,\�����qz��"O�t Eܭu�6�	w-���^	{a�'��'!bgP:}^�rF�gf�X��ܱ,!�D��?h��0ug	?^zn�#��V�0�}R��H U�aNh�kؤI�\�E�>D��S#U�I'D�(��	/ꄝ��?D�`2�kŔJӀQ�P�AI�(D���v���`�j �	�\����1D����:څ1g�X����0D��z���%* �t�1Qhv�"m�O�C��4o�9`�FE�EB�,i���, �lC�(0��`�D��h�R�h�O����Z/8�,�����!��A�P���J�!���(���01��M��𲂏��9�!�{�R!�Qh^:n�8h�����4�!���'Ef���.ܡ1R�p%�T�џ�D��ᚈ~=+����g9���+\��y��H�*K"UBQhܰI@�A �.�yBJʅ`���$�A�?L�
�-N3�y򆇣F�d�94#�rp�:W���y"�00*��棈�y.r9W�+�y�V���K��ޅ#�=�Ǟ��y"oQ�(���I��n��%]��y�%�KqT\��>�Ց� ��OR#~҇��9(8���cV�m�b9�&��Xh<ARNOlT�Y�OXPMʠ�A���0>Yv`E�8�NE����>����'��U�<yp��6ReDSsa�1|O&`���Ml�<E���n9X��%+�F\"�H�S�<��G��]���6�C�r4M1�"O���4(��R�Ԃp��FY�����+�$E�G�!fv��f'O�+P�ೠO�]C6�F�A.<�3w��N�n@���<D�����"㾸y1k[Dt@ч�O��=E�D� (蒈د�0]s^�2�� ��"O(-I�E�3�؈��I$>�*@�q"Ov}�q�ʪ]��agG)-d�"Oܴ�Gl�scl���Ԝ,���hy��'NJ�A�>!J��gF"-�PU�-O���dN��h��f\'Gߤ!�$K���{��(�X {����(��U-D�_Ƣl8$"O�9��| �=T��&Æa�<�TmES�`����X���Z�m�S�<9t�޿U`JiiVAS'�viZ��Q�<��IUL�H���%�X�|��0�O�<�2�d�I�ѦкX�F�a��E�Ih��`k!��^���Y�U;"綕�D�_���'�������x����'B�V^p�1���>&�C�	6B�QʂN�L�>��"��$*�C�I�T4L�	�g�53�����X�q��C�	�yP�8�E�M�X���V|C䉼��T[6��.8\����s�C��72~�SJ� "|�@���-E�TC��0�X�2��k��0"M9U2C�	�O�ά��B����#��(�B��)u
��[0-�~�%h���Ph�B��3p'���� Ń)����i�s��B�7]w��K2*N�P�h���K94���=����������b�a�'A�^�ыc"O��{@�Q${�(i8�F���T��"O�ȗ��z��0���C f� Љ�"O����DПt0Z���d�{r�pW"O@	�!	 :M
��QmT4{�*5"OB�ؔ���r����f��G@-��"Ov-(��v<^0Q�ľ(��Ʌ�|2�)�S�7)��"�͐w�x��ת�6p�>C䉫�"��F#�2H#bТ���_C�ɱ=s�@0¤X+=-0|b&KH���B䉅`
"�ҵ�	6Zy|�4%�
�B��=l3-�Q��(0>A�ScO�p�C��5Q��R4�M%A7��y�FڔC�2r�<��(�4R�|{E$K�TT�C�=��$����.%Xƴ��� -قC��4YO���EjI:��Jg ֚�zC�I2Y�)�gI؊2���P�S�M�hC�	/om��휘o���ː�3�C�4C��x���B�{C&��c+�G��B�a�z��3����훧��b!C䉠+l��@�l�bb��fD@ Z�B�	EJк��܆cj8u��+�D5���0?)�J[�_dQ����_٠a�EeK�<����"l��3�i�7��m�	7D��r�)�)U�J �4�ƫnC��C�5�$�OQi�Nd�Z��;���C�"O)�r�& >��BC��P��"O ](��G"hٖ��g�J�UX6qsT"O.��u�8:�|���/R9I���"OB9����9Ie�c���A��Xa&"O��g+
NH�h��/˄m{��*��',�LH5*��g� �.�J.����%D�P1�L�pC�ҁ�0cc>���9D���%k� ����{BV���K8D�А���젫�`W��&��"D����O���!*�a��l�@!�U@5D��Nϛ}[<��b@ޙf�n����2D��@��K�H�Zh�P��?<6���0��������� .�:�0`h��C�p��C"OX�:��ˁ;��Y�RJ�!e��"O� jŢ���*�� i	:\�u��"O���Ǆ�e�HLj H�6����"O��7��� �#��<)R�-�"Olp�W�4:���h�( "Oέ�S�־C����@�ҝCS��q�OJ����M]� �޾}�d!��'�ў"~Ҥ�ψ�ˆ'Β͠��c�)�y��D�h
�*T�U����H9�yB�U��A�4LQ�	J�
��y�N]�H��A���̼sg��CAb߹�y�%S�=y�Xaa���g�E�  ����<A��dR~�xB$((�\8b�����	S����<=p��I�DeDܩB	,A�0�B"O��%J�]^�9![&2���"O��m�*2�H<q�-N�=��M�"O���Ǝ�SƜ1�s�ڥv�^�H0"O���*��tJ�:�,]�e��D�P"Ob�"`O	)6����0hvpM��"O�Y��WA)�0��R>f_.�t��G����6���n�0t��h����+�y2�O�v�*�L�. Ґ@ٱ�ƙ�y�N��BH��0�x)2����y�&�%1v��ŉ�ƔI	���yR���4�2Us`�V�h��K°�y���&!X�����Ą�� �GX��y����]�vhpe�*d I���y��W�@50�rV# )��Sgk���y����}�:���HU"q�8��&O�'�yBB��`��I�oG��v.�%�y��:�h���ET��I9�iR��y���9�d�AN�M�&`@�'�>�y��?Xd�j�O S�p�ri���y2@-n�x<�q�ЯI�F-҈K��hO<��)R:��P�MR�Eu�mk�"����'zH��gCXgJ�l0��Ξ�H$��'�D\J��ϐvR�2�`æ~����'�,�0u��]ᆦO�{�N���'Z�@��L�qʨH�,R�?#���'�EI.�	���SV�j��`�<�a�>e��
G�F-m�4)��BM@�'tB�ӛt� Pۑa��Gn\���˗6
8C�ɚ��m:�@f�Z1�T�׌:C�	�o0�M�q쓝0���!��8*R�B�	�=X� V拥M�]����i��B䉽>���3��Ǯ��8K�c�;r�^C�IN�d�AF[(���TF]�#�LC�$`�LZ�j�9���Q��tQ*C�	0r��] �$�!baR��G/���C�ɺB�tݩ�0n�(#�T�C䉹V��!S��%�����H��=�|C�ɘ;1�s��<@�xQUdǃ�tC�I�w���ЮL�A:h(z'�J]�B�IO0h�y�cœRP2�)��$V�B䉎@�D���օ;Ub\pň)��B�I�-����3R�6D!FkG�I�C�	�k����c[`��J�Ţ t�C�I�4�a$	�)�F���� 0nC�I�B0�%rrc�+�X�b"J�0��B�	,#!����\"[B(`Fȕ/p�
B�	>e��h��m�!C2аԅ�$-�J�$.��V�1����W$Ay�N��S�2D���G�B�|�t�@�
'H�s�6D�$Ó�G���eG*��xEL0D�PڔfP||�I���s��p�/D�� L���O�W�޸x��[�M��;�"O����oZ*V�*����J�~�v��"O�j�kA9x���욂[Q�J�"ON�Q���Y�(�h_)9�h��"O���wo�B3(e3�*�t��M�d�N�؂dB�"392� �gF�U���-;D�`[WcN��x����vӎ�j!g:D��`�N��
a<�kn#
VY��7�O8�ɔd"J�R�]�f�Q �Q�6�C�I9f��x��ɀS���@�91���$��Jq�'w�8�HP��<%`�ȓl�>՛+O%y�������q�<�?��$�t��k��i�B1��KUel�ȓDe�MO Ӹu�e�5kF@��ȓ^�Y�B�≢g�Y�v��U����<I���b�!�G�S%vj�����P�<ц��Pk�H%�N�S�����MK�<)�'��z1�3K	Gd��tF�<�#��ncJ �`C�
�d��KE|��m�|�R�P�Tdaa��6�qY0�?D� �H��H���#��Y7����	<D�ԙ 5��`�P�ې,�6d���<D�$��ѶD(A%8��:�#-D����H?}�u�"B�Lqj4��F>D�X���X���P9�����<D�pI�D��
�T�q�"�E�)�$�;D�`5*�)A�Ty���X�2"�-X"�9D�	��
g����� 1���Ŧ-D������"�r�Fԑ�n�xD�-D���1L��{��q���ҷBȄ�� D�<27Ƽ��Q�%oܘ�N��V�,D�H�ԍ�X�ZM�ǕfC`-))D��c��
4�H��	��*!�Qd<D��A��V�@�R5���ȻT�!�d�-D��sr�&K�Z=��F;\�(9Ȣ�*D���3�a�}Z͂	mF����)D�tjrMO0Dr<�ӠcB28Ԉ�#fn)D���OJ�NmЁ��"A�(C�p8э#D��c�m �� ��@<����&�O����*Tؔ�<k�J����B�3?V��B�W�x�rf��'e�B�	��
�˥��q����UCs�B䉝e����3�7S��Yt��,m~B�Iu��t��'ڂH�i�kx�B�I�^D0aA>��Pe���e�~B�1}u2�m�x2��`%�L!8RB�	'33�(�5�رt効x��]�'��B�I5}x�6L;^�"ʚ�MݠB�	�>^���n�"~���%^#%T�B�I�c�LAi+4�vx�3��G�fB�	�zyb�`P%�s.^��0c� BdB�I&EF����4i~T�1�%�)��C䉉'�t�R�?/:�bq(љ{-
B�ɵ��0(Rh�"B$K�?	��B�8�1Z��A6M���
�4��B�-'���q$j8�Y��k�98zB��;l�ȰSUꂄL�)!�X��VB�	<a�u*�-�-X����b{��"O�H#,��x:�VF�1(�h�a"Oy�!��~�<� ���v�s�"O���ԓ?��e�4�'*�qC4"O҄�LS�ѓ�L 5Az���"O�0Z��+}l�)�ǈ���L��"O�8��A���09��esB��"O� �1�EDZyL<St�I s���"O�iIS�D!:�h���U	~�e0�'��ɒ^�M��I�r����噞'ʐC�9'~�AǢ˫b���P�j��6�JC�ɈK�조�a�&_:���e�Du��C�	�m;x$زfű�% 7$�DB�"O�iC�m�:�,�	0Oup��u"O�`�4�N�����gM:Kz�{�"O(9�e�4:�d�WG �uA�Hr"O�]`��J7/^tꔫO"��4�*O�����Gl�P�A��C�P%��'�f�z� B�<�nQ����#4XX�	�'f u���	a|�t�#GG-Q���z
�'��!�ui��lH�����)Q�D�`�'a�!�P�e?�q��'���=�
�'p~cE�ǆjb�B҂��EіY�
�'l�m������<�k��=�&Ū
�'�T�
@�'%�����	�*�X
�'PNe !/X?`���ѣ������'L(��$ʹK<i�'�ϳ�pё�'|T���>� ��b#T��c�'���q��A�A��YPb�c�����y2�	r1�$ #��iQ��ѕ;�b=Z��D�������$!�J	�x��\-6T��rAJ�G�Z��ȓ�DU��ł:h�2e��de�ȓeepU[R��i$�����N']%е��g]:]"7W)Z���Q����{���ȓ� �	��<w�B��sh�,���G{��O���$��7��qyeB�9�bQ)�'���3��L��@� �&5���'�HT��G�Qh<���(��z�'�ܭ�B���	s
.(��}J�'��l�#/��iP8H ���~a��'�h��� � AN� �R�_=����
�'�d���>Q�����2���i
�'��Q����Q?x���Ƕy�ԈJ
�'|<�A�T�_b*�"�h9�p0)
�'c<�K&�İ/�eI�E�.�H�
�'|V �!"�]�8��"R 
M���	�'/T��wJ MW��UT+*e��'�$<���m3�����6L_�M�'�(��6@S�H;�I@b��<T=�,O"�=E�T�KH��p��-���zpϓ��yJ���*`I�,'�A%���y��E���q�Q�R25B'�\��y��U���Y6]đ���̨�y"E��b�Pa��E:5�8 �B��y2	��`�T��d�	� F��v�N-�y"���U��!�d@�p���!AC� ���hOq��Đ�N�Ct=X ��k��$��"O��!���&/jeBg��M�D���"OZx;V�<1�I�'��6�-��"Oԅ;��~����'�#��M��"O�<�qE��,cyKt��d�޽�"O6��7�I3)U��ă>:R@@�"O��s"�z$��Pf#��N���bR�|��B�S�O5$�H�_��Abj��g�]	�'�4�2#�;��XѠ\�Z��d��'���#���,l`��EA�L��	�'�j���ܵ5*�wKL
F�f�h�'T���+��R	{g�*bVԊ
�'A��0�Ex#������H\x�'ў��O�$���z�$		n����'��c.��N�k�8>�,�p�"O� �Y7�~����&�!/wj�S5"Ozead�Jh9:�Ϛ�K���"O���A�E�	� x��A 6�T�v"O>0!e)M<����u/æF���!"O�m�W�Z�h]l�)0E�UJ�"Ov�Z7,	�twl���C�U�����"O+R�F�l�p�u�W�`�j�@�"O2�B@��c� �`a��>�:� �"Oh6,��	fL����ߍa�d���'��\�H�8����'3��xHr@G�!�DO�"=�١�c�it���Q��+���7?G�9��bۈ���;�y�*��5Ѧ���nFf���)���d5�S�O-T@b�XD�BM��h��o�AH�'@�ـf�ҥj�zeʤ`ٱz#���
�'3�����*�\Acםy�l�
�'62�c�Ǚ��=�eÌ�@�:e	�'����B�(A $	�[�e��e�	�'Z���wn�99��-0DQ$T=&���'V(���C�clZ��Rf�cu�I�K>���)T�C��e����$C����h��Co!�Đ�T�b�aaԕ~�h��Hfe!��"1!���ek&j�>�Rvh�"g��$�k$t��V`���T�2�ͪKb�B�I�F�^eӡYd�=s��ʟ:Z�B�IOf(�+�"S�P�"M�	E+.C�I�J<nx��F��:+i��P*��hOQ>�Hĥ
&/L�F�(Qb�rg�#D���$O^�j9�tB�Y�� �Y��"D��8u�F�(�h-�����g*O���a)5��`�,��m"4"O��*`�ѵvOXa��W7V��� "O|e ��
,CFҨ(4$�4m�,M��"O���Wḏ<8 ̹�C:c����3�|"�'��Orb��r�H�l������ �� "0D��*��a�^���B�yCR��׊.D�`���́moP8�)� u�UP��1D�,��AX"OB���Cn�> 
&(�%0D�4����96���T�"'[�@�gh8D�䨡I:thaPh�5G�v0H��5D�� �Β	��m�R�o��c�7��<�t>�+˜/Fx��1ņ�|��D��V1Nع!C��qu�4��bОDݮ��ȓ<X@K��R8k`�Cデ�:�&����,!{>�0����TA�H��L��B�I�]�����d�r*��:c�B�t��B�)'i�)���QB܈�`�+PYvB���j�jp�M�<N����ԯk��Ї�3�F%�O�K����@�9#0BB��?'_Թ���q�0�p!�4x�B�	�.od) F�W���[�jl|�B�I62M� �
�,��ip��
�B�	r�����R?PJ$!ە�Ǻd��B䉇0&�d�ƌ�6Ԩ�&�C!��B�	%r>��@�|I)��E�I��B�I
AX��q ��	�LY
u�^C�	Z�$�	�OA�U4u	�[�}O�C�	�A
���jY�p_ڠ��=C�B��$ow�`�P��0x�|@&�SwnB�	����䏄it8)���*�^B�ɖi���@�n�D���n�B�	k�Ҵ�V�R��څ
�:�VB�I �L��T�xH���,Ѓ9qBB��-x1N�@!)Ʒw�(�+�;%l�B�)� ��An�EB(����R%.��6"Op�D郢T�(|��<H�~�0B"O�]���-����� 4e�\��"O�0��gُl��0�`,�o�ޤQ"O>T�vm[��Y� ��4&,]�O>͚�/Ϊ'�ؔ�T)>�4@��E+D�<�(��z��%S�+N�$Y$��A*D��"-�l�А"� �wi�b�(D��j���N3�dC�M�{����3D�L!e��w7��� ��^�0Yb&�-D�8�S+�f!Z�Y���
M�@ٱ��-D��ÄOZ�Z�b�� -ח�$�A��-�OP��4a�4�t���{j0��T�λ=Q�C�	 	�L��S�V�(5y��@��C䉠^�P��C��b��L#!7�C䉲<	��:��/�� �KFgh�C��&^b��Е�
N�<krjW(<�.B䉒Q%�(A��#}���)�`֘N��B�I�yd�T��%A�}�a`�I�-�����0?q���!B�sNZ�=l��É�C�<�e�U�SR9I0GF�	)���6�B�<a�Y/7�>qcC���0���'�8T������x�ɒ��.IQ�Y�g D���V�L��*��Hĸ2��C��?D�6o�mt|)���;8�i{�@q�<IV�.HF���P u!�˅p���hO�*�h�^O��Z�������[�D�'�ɧ��>��c��r;a�(��8���CFo]h�<�a�#6l�����-z=0��dBM�<�Eh��}&X�;% �(b�JܺBBO�<)��
#m��C�I;��QSp�[I�<ɇ�O=C-Rx1��Ð�j(���G�<�t닔	�n�T�)^ZC���A�'a����B	��V�U�6=3�ٞ�yBnY�^�0-h��H�%�Z��K��y��D�3T�0�	�|ּ#uZ=�yRϨp*f���I>���r�o���y�,c�J��lE5�*m�T��&�yB��	P��a�2"�9�y�A�ڍ�y�(J�cmv�{���`�f��d��yR���7V(ĲR+G\P�2��i9�'#�ڔ���N5�U�E��7b��`(�'>�H��R�")���5HJ7rlQ�'6ȜX��%X�Di(Vd@�@�,�@	�'�hQ��*��R��$8��U
D��P�	�'�T��aȚ=�Bț�F��6��X	�'n��R-M+B��<�F.%Av�hK>����*Q'��8A��+e�l�����Ak!�d.�Sab�4̜��̋*g9!��2#���-�p��u�%F�Ԛ�'�H�D�d��1!�H�wI$�z�'��	3��� ��Q3�D$uo���' ɉS �Pn�D�!�0|x� ��'X^�b5F��.��`�{�Z0�'�҄ǹ�N}� #K�~���'��p��VK\
Q��H�r@�'�� !lײm�T#oR�2�����'��x��hN]o��ip�F� 4�q	�'+�Q4�oO$(U�S.{�4*	�'?�`h��bl[ծM�t����'�p�� N� *�$Kd��5i�\��'��4�p�Z,z��H%�ěW�j���'��]1���0}2��D-A#DPH	"�'�MC�/�39��"d�ĝ5!<k��� X%@��v��Q�"5l�j�"ONX�w�\9'����e?V
�,�"O��Bv�*L�<���S�]�NH@�"OB�k�AC�8툕��;?�d��"O�4P�Жo���q#ܙlϺq��"O�����J�	�Z "�L�)>���"Onq�bH�.?�MY��X�V( �"O<�s#�����b�	U�ţ�"OP�4�B�T�j#R��:����a!��#3�48j��$? �(�INd!�5�%�A+8�]�/E�uJ!�$��&�p��'���������%L!��L�4%���4���2y�f�V� �!�$��]��uӤb�H��Xu���T�!�dW�<�J��֠M'|���nX�!�䄮�d�D��wh�Y��G�1�!�dS�|� ���t���b�l�A~!�\F�J����qz�<�e�J6TL!�D�	���6�O,�� ���#9!�DD�P*D��5������bF�"/�!�DS5E���9p�ϙX�nx���	%~!�دem>��RG��j$�w�S�s{!��"��P��IGM��'�!�d\�4�a��R1X��	d�S?}�!��ѡZJZ�rBG^�:�d�Ȃ^!��߲�X��B~�� (�)��F!��KQ��M{!e'Z�V}��>c!�$S�V�P&Ğ�u���X��'/�!��Q/:�����@0�c�*�!��Q����@�7{iYa�!��$S�Ze�S��e����a|�!�D^�f�4��C��$Is(�X#�1�!���?�Z�(����K�"����ѥ`�!�D |;ƙ���ψb���O��C�!��@;Av0 xBI ;)N�a��=gO!�$J�6��� G�1�v��k�A!�$B�;F�����2�bI�EjR#!򤊖3�.������	�锝!�D@2/�DA�(E=U���:ЈO��!�D2l�F��
�.��q ��ͪ�!�$4(��G[�Vy�YJ�f(�!򤁎/�.4 @P*nr<`h�E��1�!�D��v����O���Hq�/(!�اc4�i�tG޷,]t+pO]!��
�s�T%��d-'&��˅�O�N�!�$QdPA�������盆2�!�dئ!	~�:¤��^�9WG;g�!�$�w�:q�r&J�r�����E8�!�D�1D��A�l�����J��J�!�dYz�(�� �?i�"H�VI�`�!�$�}%(�YU)�Z��_>�)[�'��,`�F/�h��,��6ݜ�9�'A@X���&�6@3���5�j��')"��ro��N�m1�h�3)���`
�'c�B���+aO�I�HL'�����'�T���M�]eK3�Gp�: ��'�=�kі�^�����l����'�	���ē?X�LI�ۘ_3�5�'ɠ= D���]r�"upD��'��Y[�(θW p�ӂI(Ȍ���'�B5c6O�3Y<�u��J˛b"��	�')��2��,]�`��H"�؀	�'U�}h��>{�L"`BN2>�<�[	�'����K�z:���WϘ�N�(	��� �	:�R6�t�p�?��"O杠!h�7��4�.��T�p��6"O�u�3%Q��X�l�R�*\�P"O� ��)O��Ͳe̖B�ʼ�B"Oua�K�dL�� 6P� -�W"O8HR3"�_Mv`�&�	?�m1a"O��HF&�H�B��7F� "O ��3&��+����Gb֏��,�"O⼰7H�����#N��R�BF"O�Y�-Z�07Z(r%�Վu檕�s"O�i�W�8C01K��^Ŭ�S�"O��EC�o`8�u��I�����"O��2�I5Sd�A�SD�)jfA�"O��.Qsh�R����E]�Q�"O�%j�C�7M�H-J0 �/<"x
"O�"2ǆ�r�ӡ��B'�I:"OB%�f��/gKD�6C��=���C�"OZY;�-:'d$�C��	��<�@"O2}*�V=_zh�ڔ��zn��i�"ONU�"R,գ����1�8���Y�<��Q:4c0T�af�&s/�4B�C�R�<��G�����Q��l��ű3g�G�<���Ζd�:|(��#x���y3�DH�<a��԰)��%QrƧg F��pi�G�<���H�s� ���dX�m� ��	^�< MK�l���"�
gG�y�(�X�<1bED'p�@��#8e�]��*O�Yy4G�?A�\�%O�C�z���"O��(�+�X2^��BU X�Ab�"O�Q	vKL�/,�}��&S�,�����"O� Ґ�@}��#q���-�y��.#a��#�_,I���H��yr���<�Ұ+����Nx9��o��y2��+ɬ��.P�Cf��*�J��y�b<�|A���5ݶY��δ�y��p��i��-�5xӅ��y��زQ_h�b��:���'�/�y��^�OWZ��סF'~�����J �y��Z5M��#�9|��IT��yRO�,4�j�i�)V�rN�����D��y2k_�$�1zv.#q��h ��yrM�*q ���$"�>p�L8����y��:�\��F�Pl�*`�c��y⇌�E�x�!2f�!rQ	V�y�
P��MX�dpfQ�k5�y2�T�?�l��g�!F[�F��yr���
�� U"�#:R���)[��yrH�,@��Q�C+G�$8���4&�C�	&7�C����|D81���ÞB�I�,ʈat#�/ے\�c��q*�B䉢$�%��⚞h�\� 0�J�T�C�	�b�N	����gy����=��B�	�
��Mj	lcP,�&���0�ȓxj���!�{���x��ߊ�|��ȓ-�hH�JJ*W4v[G��i^����	��� �f��"��C�� T�ȓX��H�����4�sf�l��ȓv�0���
����Jb�<9��[�f8r�_#�y���HWy��ȓ�6����5�n��lRc}<��m��erG!�~m�X$�U+,�f����l��(˷J�,P8��%2݅ȓ$j ��T�H?L��M��%���W8+�ޕ"�V`(�eȈߨ��S�? ��	Uj��PX��\0�s�"O�!0B2?DЁ���@��9�"OH�s�ZnnIbg�՛bN��a!"O�,��(�6h��� �;dI""Ob]�ʊ2'��(�,X e�:Q��"OB�ܭcV��Y�˥tfh�i�"O�m�t��)dB1``�ەP�Dq�"O�8!� Z�6)�4�B�Y�XJ��`"O�Q��	�a��D�r?��B�"O� ��G�5x�9��X1+<lp*"O� ��W�Z��rs�	�~*y�w"O�����3p2�u�r��kh�"O�,C�'G�WP��[Q�[�M0��"O�Zv��L,|D�5D���Y��"O�\�F�o�F�Kf��
�\�s"O~�µ$���9��ǯ}~�e"O �!�H-
:���A�;�%A4"O$�y!G�ef��g_2$�ȑ�"O>�"��py���4��1�"OlL"6�Ҹ ���*��B*bxQK�"O>EC�OC+p��)Q�Z���"O@�J����d�q.	8^�:�3�"O�P[P�N�)��t;�c�<{���z�"O��rK��8̙�W�
5{�x\0&"OnM�� c�&��$Q2h�(�a�"O6*��Z��²%܃BG�R"O ��Rk�W���EO���Kv"OF��U
W�����IUHɑ�"O�e�`��� �&!�cF&(t���"O�)��ꂰ;�x��[�e��:"O��p5-C�m�Б�@�85�5"OLRC���2<K�-��j����"O��#��W�������Sv"O�MHT"�@Fԭ
e��D�veIu"O��1H]4SO`�Cŏ�ٶ}c"O�P��b��Ч�X����"O6�Y�Ðx�@ØZ�M��"Op���y��)x��@�H�[ "O�i�㘎>tt�0q!���)��"Od�a1O	;
WL����%�m(�"Or�0�� /Zh���� =y�@{�"O����'N�L|4��p��;:����"OFH�v#��(�����إp%�L{R"O\�:��z�FM�3o�?�x�"O�j�AS*���qN^0�Vy�B"O�P�cq��1ƬA���"O~ua�F�!��0b�"TfQ>��"O@+3o��?�(,�'g��tB�0�4"O8xc!ڽ�ZIE+ƉV2 ���"Oz CGH�*��%Z�Ĳ@�XSR"O�9
d/P5� 		�CV&�����"OF��bH)0�pX�̞"�� ۂ"O2q��ڕ��=��.7�*LBf"O*�Ӌ��AY$��G��p/�l��"O@��®��
�@(�aꆿ}����"O`e9`�@>��J��() ���y"jγtb�80���0���@��?���d/ғMT��E���zc�@y�E�$-��ȓp2�}B��0�"V(k#9��g1D�0����#XEQ�τ
}��Kbm<D��Y�소=Z��i%#�1�$P�./?Q	�k����e]'c. !6�\�Ar">Y��!�O���L0Ja�|K�E�J�����
E!�ć<m��t��_,+�B��f��+ў��3� v]*��&s��L1,��%���򖟄����Q)�H�����[�M�3�R$}�� l�����>隧���l�P�°.
Y�ܔ���HPh<���̧`^�Eb�����
�
,�Mkߴ���;��?�O>��aDF/��³˰M�(�
O(7mSn0]�P�+%����	�/q!�DR�e��,B��6�$�"2=W1Oc�dF��6��t�&� �S��$�EA���y��P�ZR��(1�ŋt�N�@2�T�Of��X>'xܼ���6��AgF͎*%!�B�C�\� ��>=XDZg��+!�BO΍�����m!�� =�����'Y1OR�����'gA0�׽H��(2�"O�@�S��!JN� �@��J�B�"O�9Xt��"9t��W�D�"��e�"O~�!@���zת8=P,�
 "O�%1e�ۺ�Jh�D�[ 6��!p"O8!7G�V�T��R0B<��0�'ў"~�c�8{��@�`ƨ%�2\PD����xrν<��A��0 \�� �Oh��B�ɿK��B��Q� F8LqElY�;c&�=Y�O��	ئ��OnZ`	�{Z� ���qs�Uh�'��T��ꜘ9Q,Myu�B�	���4�c�DxÈ�l��\ڲ'
�%��a�N}�R�G� �4L���j�؅ȓL�P�!a˜�k������IV�9�ȓ��Uj5��S򄣱��<'L�'�~҆R�E
�I�K�y�VQYcHK��'az�cJ89�\�'!�%0���W��y"Aՙt �P1ӭF�d�r'�W0�y�Ԅo��LñC���jW��y"�W�	$X#�� h�!&L��yb�Lu.�u��6��݁�`M	�y 4�A�b-�-�R%{�,�1�yR��m��5x�":���jT���yb�-��q��o�+�"(��5�yB
ƹ7��jW �ȠRC��y�k�k�t ��M�w���#�X��yR
��!���iJnlB��
��OH"��F
vT�S ǴH�Y7(Rr�<���]t~��B̕t�R��V}r�)ҧ&-�u8�c�G�4��Y	8;0<��IEy���-�&���*��ꐣ��HO��p>��lT�!8ށY2�� @���D��<0�O���u�dq������4�;��H�)�B䉥i��$3f��[�2$�r���o��6��������|����4j� 	vGϟ'RT e �s�D���h���x�ϑAPHģ�J,���<�E-j�C.74a�6Eޅ%!�h���z�'�`Q"�^:�!�!�.�	�'in�b�K
�r�6���L�, Ҩ�	�'�d�؃��<?ZD
b���i��'J 4H�"��B�����+��ř�'V��ɄH��M�R�I�0�֫�m����d7�d���8����;H	�I!=<h!���T��瓡j( qB��M3SN�OԵٍ�d�L�$��1`�uc2����|��,���ybϝ�NnJ���@.��;VI���M���)��		ꍍRm.4�0�6�x��ǭ D��#��oJ�t(tJ 0��cUC�O�M��	�+�&����҅�1�%*A�
�^��x����!`�{�f�H_�L#��ր-�(��ȓ:��1J�ͥtv�u�S'~��,��ē�?��'����ա�f?��°&̊I��p���O&��� Z���B)T��� �^?ʀ��2����<ٍ��O�,|H����t�н�![�r���'���ecĎf�f< ��`)�F}B�S
�дQ�h�Z�XvoG�C�n��M���Ĉ�:,c� @�ZDB�ɂ���q�U�Z4��H��n�H��t��h��|��׳\v��hW2x����r"OFU�P�Ǔ(���`e�u�g"O>��7�!;�R�Ӡ��<�H8�"O���]��P�C��T%�<��s"Op`I�͒A�z�{ �Y4ڤ���'M�'����i��\��c���l��'0<(k�i�*Xd�(4�����)ۍ}R�'|(��'�B uX,�TEW���9��[�4��	�Z% %A`��.3;��Ì�+7�`��X���N:4�����{J��V+�4��<��8,R!M��)S�|!�H�2+����?���~��,Y�Űs�hZ@�7_S�<a�mJ �nt�⧛�/�J+#/��<y���w����q��a�ԁ�4;0C�?�fy ��=]� ��e	/Nd���>�#�Y�	�p��\b�	1�f�<� 8^�|��F���ED�W�<Q���7]
��.
�Ԁ�kܓ�y���!�Dԣkr�`5	�C�:����wD!���m��@{�I�%� �D,�Q�!��4Ej.�͗����R)ؔg�2�F��������c@mX�P��$�S�!9D���KZ%]�x3���' �2)�G�:}�>A/O$#<1�C�!nƖlqg�ɧs"<̘��|�<RD�>g�l��B�"I�$��Ү�:!���)�矜�A� ;�4�Q�K�5x��$Ej;�c�D�'����&)��P�B��	d
���|�B�=�O�a"�3���B�M���Y4����<�O?�m�l�Iݓ(bl+�ΐ�fISS�!�D�h�P`1W�%z����� !��O��DzJ?K���34�,L�N\$<U
�# `2�O��!U�qk#Nˇ(tLbJ�g3���F����ĥ�~`��E���'b"@�ȓj�~)��O?oG,4{��9U���ȓgx�|��"��2z���D
ѱ}�PM'����_*��9�Ԯ?�ԝ�b��'h�,B�I*i:�Y��Nֹ(��ib�יX�B�ɾn0�	�1M�CA<캡�ʌB��C�>h}�1	�LF��`�@�!6B�	� ��R ��Wc&D��c�J4�B��۶dЎ͇DB��T�	$>&B�I!O.,���]���]��ᔳ'RB�I5I�#��L�`E[RĐ6e��C��=�,a!LA�` �xЇ��C䉍��d��(��҄U�z�C�ɶv$B� ��V�`&<+A�Q&dpNB�I -<�@�	�$�.Y[��Q#�TB��:u����5��t Nh�*B�	*o�(:ի�)c��0���4"~�B��>,b�2�b�6���煞5�"C�I�d�\!�6
���iU�>B�I�K��1��_�R�����O��C��"u���ɦ�݊3%Pb���B�Ɇ|xl�a�+}�ܡ&ީ	��B�I�q��z�.�7��\��
 ��B�	/�J��oS�M�Ż�n�._ƒB�	�~�8���4tzޜ��C�;�B�ɢ�n��A��"U�P(��B>b�B�)� B)�-_�!���o$�z�"OV̫����2ZPĢ���f�T�j�"O�8��K�&t��h!�b��8"O�]+a?}4|*��l�h�"Oj��5,F�Br.�Y���7\�"O*9y"
�"m���f�6��P�A"O�u��M�4v_6�H���+{N��"OP�Y�`��<�-��i��π��y���1��T��D�Y�عc����y�݀i2�r�B�М�C�D��y�QVj�����Ch���� �y��E$#�j�Ғ-�1	W6�a/�,�yRFF�-Oʀj�@�)�؜)��y�ē }r�Ƀ��&8�&�ɪ�y�혍q��H9�KǢ ����B�B'�y�@/O.��+��_%q�>���6�yR�J�P�d�	`!����I�����yr'˪=mv���	X��-2u��$�yrA�_�N(0��ٶ}8T��yr �=f��Д�Ѡ�0������y��A�&�Uk��	^}"Y���ɯ�y ��,B1��bʸ�Za�)�y��C9@Ʊ�4I�*<�p�Ž�y�`A�F�*L�b�N���s��?�y V�P){�c5Ex�IíL��y2 M,b�Lk��MC��2B"K��yR"Z	�mx�I��0�B)�A@��y�/6v�V�A�Y@o��������y�F�%IHL7)3v��� �˽�y�kJ�K��u�ͣ.���'.�yR �*&p(�!ǚ�zy��a�۾�y¡�;&���Ȍx#`���+�0=)���?���`Ԗ	zN�!�T�c���Ra%7530�k�+V�<���FuZ��O73��M+7��Q�<�1�%S�
��F͏�l`���\{�<�c�T��ص�sM]/3���q�J�<�"E�-3v�U��	'C�0yq�E�<ᤢ�v����O�' �Е�5�@�<�3*˻5�bML��v4 ���<� -��`�����"+�Iy���R�<�eÉ8Ebx	�P8��C�G�<�#�I*?n�H�ia�>8S�nX~�<��	ѼWXp�K��_"�,��7E�y�<��Ot���IK�-H2��B�<)@�)\V0����<9ȼu:�.W�<�h(nf^�"�;dtTԑDn^Y�<�ڏX��ȵ
��?`�Q(Z�<��Ή(�@�Q�M�1G/6Աb$TT�<�SS�&�$x��動
bz%�b(�W�<y�B&4/�ÖH�&�� &�2D�XBd"�*;
�QF�R�<S��X2�%D�D�$꒦8�>(�auX��U�=D����$�6*�R� ^��1�S�8D�<rVF�'(�"����+v�mz� D���C�+>��jA"��8���;�H*D�h��l��'�d5�$=��uqW@)D���g@�h�2I�u��}( �2D���b�IN�i�l¡y+�ŉG0D��k�"R:^�䔂gD�%s(2=��1D��a�هf ȭC��H�9�r� D���2�?�T�#!�S�h�A���>D��2��ڬ���1�
ڼI���xCm<D�\�#�,t1̓�lվf~����!D��b׋8���E��w�|1W:D�� X�)��3_ �S󉐟HMh�"O�3���"7�Z	A�ġ@5�""O��� �̇!�j�Qc`F�k�X��W"O̥��Tf�u6V�c�� �p"O�T"�bZ<ĉ���v` 1�F"O��aB�G�EYt�2E�$8VdD�"OT�J��
�)v������K��E0��'��U(�0O�-A�M#sX��l��E�"TK�"OdBf Ҙ�z�P��U:�Z��E�	�x5=0�S9	!�e�˖m4	`m�E��C�"k��嘽�*���Qw;p6�!�� ��{���iԞl �G/~z����=�J�	�'jf%���5�1
 -�aj�O��)u I8��=%���u�P���/mYV�	��hX����@�S���C�;O�x
愗"S��hY/Y�y��6(]�%�m�V�*�@f���HO�9酢[��h��E%�&�PQ5��1s� �BD"O��4�E (Z(�r�$h�õ�'�\
���ӤY�X B`��]A.��k�9�dH�ȓ|c�m�7.`6�ቓ�g�9��i��93<����*�2���ȓV��a�� ��D��$�f�
7|��TA�Р�֞\��g
w	�D�����Pa��V� ɤ��,�<���0�6���d�L�#e\*-�Y��W��b�Ζ�\��J&2�T$�ȓT[,t��b� ^����)��� ��~"ZHE��\�|x�Й7�,l�ȓ>O�d�f��$aJ�bd��@�l���f��f��%b^�rVIźl��܇ȓ?Ix9a�H-'@*S�8N�Y���zI��=P�H0�Q�G���\`��r�G\;�@��׏p��ن�c� �؂�=����yHB���B��	rfϟ|��Ȼ4�ˊ��U�����B�TJ<�� ��	�ȓ=u*|X��"*[Z�"�a��OJ�ȓ�XQ�Ɗ)�U褠Z�Kl���7RD)w�B���Ur�G-ON�fHY�Oe��S���1�K��0>��̾q~�2�'� V
�����j��\	1)��-J� ۿ��?��(��8�j�8��H���P�C^����c�FIyr �Rv%��oN�#@���dK��y7���[�æ�ޮ�x��m�yR�Дi��l�Gh�*�VEcC��� m���͕{���B�.T65�8�sjЕh��|���+��)�ʼ{ �ިA&�����G��m���Q��?z6�j�iS�0P L��](6珙j�D�g�
� ���/Yav�ɶA�6zS�830�́��c�Ѳ!
�	)��j4��L���r�N;�	�Wh�AKe�H��
�,9#%�\7#]"t��hѴ5&�̓��R��,#vƁ3�Qs�L>l�~Y��'�}�� G����@`FU����jQ�*hL �N�Obi5��j� U���Ǆ���ذ%�
��-����-<o�"�9�߀zP�����e�<q �[%�~�ƨ
9/؆�/�#���)"���d����m��)��
��%�j�i�˸-��4�X���Q�*ͼP��Eہ�˶�(��"�O�0�НA�<{ݴ|N�L!���&"۔�i��F~K�`��H'���1⍉u�b ��$U��Y���^Dp��2�͢gB���u%��O�O�4�6�H�=����DˈHQ�K�n/�؛è��v<8x�g�Hr�4 @3j	�x��C�Ã�|�LpW���=	�bN��vD�S瀃t�ĘpQ�R)��Aa��9t����a1����rL�s���u�ȄH!���Q-k��� nН�Ӏ�L�&DA��>tN!��5_
�)��B?ULQ{v�ӃY(��3#�d�*��s��O<5���?5Z��)I}Zw�T���� 8	t(u���T�Y�,S���D�>Pz�(���#�y��	�al��dI�J����D@��n���ƍI�Lؑ���<��`i� ����=���q
�el�(Ö��(?�qO�}�4U��7z�I�4��Y��7��>\1�X��YS�:��"%�!�d�)F�r|��JѮ,���R���ZD�|� �뾬2�Gw�ӗ��.Ū,����ؚG�f3���L�!�	;�J�鏤e��ȗ`����	`#�#��@�O|5Q��ǐB>���� ��B��/#F¶�ըߪA��'����>�2#M�*�X8g'� B�
1�rh� ��O� pq0�'=���N�v��0��/T��8��^t��%G�5�?y�lS/8�Bֆ�%kP��aF�H�<w��}�����دPdp;��}�'���W��P�O�%IN&$
,@ e��+6��u��'�!�E�?Bm8eˍ� ���	�'p���}ֺI��j��rsr��
�'�����R.�X9C�d�Ge��K
�'�2��t��,(�
������:�Ts*O��#���Ƹ�(�^��VÉ��Y"t*�,;m�X	"OH�8���8,#��d�5��څ^�!�sfݴ
;����
�0��� ��x�ACQ�c��}B͏�b��p)���*��tò&��g. ��lf�dV�+��p��ɏkxέ��Aߤ1�K�x˨�Y��<���ˆ��d�r*F|���2���[��^9��j��X!@Q!�dN>_�6�1#M˙V�"%�2� C���Շ?c�q�jܥGV�D`(��5� (��U�4��­}%P;�$L(�y�S4O���g�.y�dy�,�(>M�T�P�|B���M���`���hO���5�J�۵o�.���s7�'�6���/ݒ{�H���5U4���0y�~5��#�*:V�A�%M�� HEL�^-ҩq�c�"[D��aE�,�1�n�1�����L�s/F��+�*h��
C#(\�wk]��q��D�\��y˓w04y(�J#3�9"�%\�xI~x`G������#_!W�=�ׄ�G�O>:���	Ǔr�j<IRH�i��ta� �1z,9�OXQ��$"hX��6���RaaU$R��A�a��d��\��]/�.>~��h������i�m V�	�R��ҨL��|���Q$a�a|򇓯,�2!�wA�� 
��m�15�i��D�T?^I�f��2{ڬk�n�JQPLhՓ>�f=���7a.}�6D�8#�0}���АFe�"<�(̚jg�p����wMxA�2��!��i;�:TeH��8�$!it��
�R�'sUh����O<��A J�Ș$&°A"�����h �D���On4$���B�i��|��-A�n[�H:ay�q�Wk۬#4��k2&���D�
54!�`'.6��S�K�|�H�8pC��s�"Ê�0"��������A�Ƥ�J����A�+���b�h�d@�<�B��S;��K5���DT(9k�GČdD8�R�^�b_�PiЅS�uyL�p6�A +��) ֕>�����Y��'>2��Ή���1p��#"%��8&�!�c �&΋��	��#'��V A�1k�Dj��iR�qFߎu���Ⰾ�d���?�na[e�]z�3�	%}Y
<p&oH�n܅��F��	=�6����٦B�3��Xr��K��8(�,>��I�<p��/1����G,R!�(l�wW.<���<d�9�
�oc� jB-ԮZ��t�c�M�Q���v�H!$�H��em�׺k3DT+C���)r()}Zc):D �.�7���jt�� ��uI
� ��yQ�"C`���P5�w�ތQb%�("z�=�4�
T�`p��"Y��*J>y�M� \������ $�o>�)��R
x��Pd��
A0�!���"ZJ�ۉF���$c֢(%|�V+�*�~ţ�@&V#1O|ͳ� ���p<���C�j�C�0Z�d,(6�Iyb'L�T�ji�'#��"��v!p(Ad��|�ٹ$N�u�B�	�d�� �A
H-V�He�(��B�I�21y�0f'�Hi����z�2C�	�6�<Xq��	��Zv��2u$�B��$0St��e��Vip����݈HւB��=��\�$%z��֝c�B��� ��F�"��i���-ԸC䉤t��0��o�ܸ¢��6�B��:lɂ�)0� ����f�s�bB��78z`}��C�A����zLB�;T�3ƥ�P怔��BN�v.�C��5˦�aE� v�F���$ʕB�B�	���Xx��\�I�j8&�\)žC�8R�]���#X|T��R�I�C�1Zz�CDM� ,����S=3�C�ɲu���t�U��T0��QP�C䉃,Dt� B��f�������2)��B�ɥ1^9�Q�@�:k�-yvdť	o�B�/|V*GU�o����>h��C�)� 2�ʦ��d�ā�˿xBp"OZu�&&ײW/�Q�	CBT$�A"O`,�r���}��C��CoT��D"O�,z��[#1� �2fP�T&���3"O>41P�Y�@����%�ę0eK�"O���D	����kFꉃN���"O�YM�7x� H��@�5 ʱ8�"O� YRD����`��'W(\���"Of��6#M�B�ԁ� f���S"OP�
�lO/u^9ң&�u��aX�"O�9��[�!�L��A�8��鹣"O*KF���f��dR*
����T"O�
�
ÿ&k�MhD�O���࢒"O���S��vԪ�*�cGeن���"O,4�3�J/=r�R����C�@��r"O��� �V)Z�(I۱"O�M�̭�"O�Pӵi�x�Bh2^�Wʚ��"O� a�&�%{�n1x%.�{����D"O"xZ!��L�V�P/<����1"O��r��[�� �n��,R "O@u��6C�Q9� �M�Zy"O�pz��_T`y�e.T_��(� "O$��E�R&�d9���4nT���"O@�#r�9}*��� V�nE6\&"O.��WE�:<��Xð�G�yf���"O~� t��(6Tx<pD�
yFd�"O������
;x���*K9t���"Oִ!T >���U�wM�Y"O������Lx�:��!a��Y�"OQtgY�w��o�;>��Pg"O�Y2���o$�� ��ǔ�P@"O�\hw�Ӑz��@��N��i�Ll
�"O����i�'u�8l�d�F*trd"OA�0 � I��9i�ʐ0.�=��"O4Y9U�C(Cn�j���"O�\����)�������Al=B"O2�J-4;%���KN��3"O���'�	vz�afI�p��je"Oݫ�+���mP�	�ѾeA�"O>��CKH�V���U���t�ūa"O�  ��(><��p fܻi����"OL\���.�� �c�3�.M��"O�M�����8�r��ǀE���� "Oh}:$"�I� �" O�C��L�"OT0Y$�*m����#�F�Z�J�t"O&���l��b0(X�Y_m��٧ˋI�<��Ţj7��ą��!w�QZC�r�<��?\��i�T��p�L�Phm�<�@�0� �k%LD^�轰R"i�<���:@� ]���<����O�<�"M�-�L��L���!���P�<y��\N�5�R�@������RQ�<A/�O-"�I7ҟ9Jj��.�H�<Yl��X�R�C&βP��شER�<V��[ 81�1F�|ސ��(�I�<AՏ����� `ϡG4e�"�JE�<�*�ݠ "A��))�$�F�MF�<q�-�m�dHk�̎��8�v�H�<�F�B��Vm8`��cU���f�D�<)W#@'IK�@�&w��(��͏}�<���P:;��qZ�!]�F� ��Ҁ��<��荾?��|h��a��=��u�<��!�)�h�[��Ό]T�t#�	p�<Al�<x���g�� =��r�OZ�<�  ���!��"|��kuGηD�|86"O0LҲ'�1`�<̻2e��x2�d"O(���d�T�Qⱦݴ8��:"O��Y��2;��ᆇ"]<��PP"Ot�`�o	�Fh�9�%�0{'�!"�"O������.]� �3�J:ڝ��"O Q�cT&	�&���T:�HR"Ob���A�n4�U#�!?#>:1�U"O}y%�ޟ�䄉w��85�ç"O4y�n 0�t�K�&N735����"O����tV��F��W"��Q"O�%����'b�����&"X�j�"O&�Ұ�^�Z�@D�6�\6HJ R""OP��V��%d��B��/.���"O�����<D?P\2'HO����e�<A��H�I6��f�Q�U҃�a�<q�F�4�*�J�k�B�D!��[�<9Po5x��a̢S$�Q��Y�<	aK�|ݖ(�P
��t� a[�<Y�O LW�822�q��CQ�	T�<���2%G~���)ڠY��U����y�<a�S'�8UAЁZ���P�w�<9�M��$�h����e�R)�ҩGs�<1`Z+g��M��
nT��Aq�<�v%Z
�.�Bd�M	&��Tk��_l�<	�i�`ͫì̒:�٢'��m�<1�EI�/&��
��IGF $be��\�<�Z����+��}�d�av*@Z�<��!@{G�|�S�� 5���QP�<Q�,(u]�M��h/�����J�<A��:AI�#V��D��F�A�<�R��*rC�x�E�h/���dIu�<i��0��"B��W�s�<��C�k�,ȃ�I�'����A�<9І͍n.@��[-�� Ha�<��I�g���&�N?(4���K]�<�����9B�Đ� q�T�̟f�<a��޼=-2�10'E2v20�B�GTT�<�qˆ�b���D�4D((:F.�P�<�WT�m��=�7&E5Qq���@�I�<I��ǧ	j��"���N��3B�n�<�%,�tqk��Í~�(��̄i?��ۛ|l��e�Ƚf$N���M�3F��� �@7|q�
�5n�a|��ÑU��a;�f��Q�I�"a�����=G�<�s5�.���@;P�܍V^�l��Js'�xV�Ո]8��MB<�!h��T�u刉��K�/����#~ޙ�%��`�	��>T�@!$�?D���k$U�~�rs�?i��+��X
l��m����6K��æO��Ci���F+$T�t�Z3�LjS<�~��r�F$J���fې����'l��P@Z"nz�m�4=��	�B�=����%� ��X���ݰ.����H�KR
�i�ɴ=���⎛��'��u���[
�X�V�	H}�ဨk
���@�����
䭝<��v�[�~n]1�S/�6t�kF/��$�&�:��B*�5K�n���I�
�ִ��̋"�H�b��A�.���p�L�Ʋ<1�'�l���I��ؠ�aL�$�F�ZRK@�(���Xc0�]��ȤG�(-q%"e�>���'Nb�� ��~�@��)�#�(e�G�W<
o���a��~�R� ".�5}Az�� x�h��i��,q��;�Z���U9v"GloV�	��s�xY����x�^6�?�`���-Q;!��H�4k	NԊ<����	?��#�ϥM�H���=�t��#m�z�)� ��7��=���sU�/8���?�EgB�]X!��/�O�g��'[x&D�5%g8y��Ə8Gٜ�C����R<�%&��ii�#4��8'�|��EE�-��E8@G�x�TI\)*�T �*^���ɇH�ȉ��� @�)���8AF�l�$��()�T ��"�h10�%/iZ �C�ާaE�M��">TX1b�A�!h@���#T�9�|$�C�&^��+�?�ck�� ;\P1B%#m�i��X�w�T+Fۢ�P��9b�`�G��i0�}�����mWL�pҩ5���;��̈l��4��e�=.�J+O�N̓n]T#<i$⁃Wj9!�"V�av�BW�B~��l2�'֨s�:�C�� ƠZ��F���sƎ��Љ5"O
<b�H���̠&��:`���9���Q�3͂%d"��H��X��m�-Qh�+h����G"O
P"�IT4M@�P�s��Z�ۣ,�$f�Pm�dD�e�9�g?yQ$%�������%�|��C�z�<y5'J�:�4)D��ts�"����#�S�Fȉ���'Xx�P0 �.U^Tڃ�T��i���B��pΛ��?�WmLl�`��˔<t �n�^�<�`
�5%�=A7��}*�]��*�R�'�6$�@J�u�O><I��o�\_�Ȋa΀�Cb֕�
�'�b�т�
M���+A&U'��0
�'i���.� $D$����L!	�'w�%��LW�
N�+��	t���'���a4�P�h&�!R'L��cF�R�'��p�ՉB�|��3wH\:Fe�8��'�Ҁ@ӏ�9��*aȔ8-�m�	�'1*��W.��f���P&�"g��{	�'^)���:1�İ���8^�����'��Q#D��<0����"Jsd,[�'9�Ȧ$H��#"�ӔFe�Ѻ�'3�P�P��]�n-s�HT�4���
�'* ���*r2i�Aˡ+6!3
�'�H��H��Qwz�a���%Td$*	�'Yt��7Dۦ?mFy��h؜E����'>�$�gı#(�h�ԧ�}r�a
�'����M��V��	k4h��:����'H�!8��)������o�iK�y�C�n�m��I�u��t��O�C��@c���"9���ͮw���a�,�'/`8�S��7TϚ1Sˑ4�0C�	�f�L�`Ɓ&͈l�����Q�"?���چ0	:�@fD;�		�k�,��ET� ���8�!�D�w1@�����Wg$Q�v�'Y:�	�2:�j��C��S�O��Pa�ŢG��\Zè�)�)��'���Kth�/y ���Mގ���钝>tc�������}�� Ҝh� N76�Db��?�e�G�M�5�Z?O2�cBa[�SSxH�GL[&[����R.	��yu��)P�4g,E]��xaplΨ*�P!������8b�P�c���,�1�'�)�yR�� ~�쒖n%	|p�`��-��$�5w�0u�#�E2��)�'J�.1�
F)0¤X��I(T@����bB���0w�y�h�=q���0N�h�P�)}�^U�I|�>ᶦ�t_d�B�/�h��1hDO؟�ȡm̭0F�4�l�kKv�;u�	�P\�h@��ϲ����.�2���h��$��f����O�x��>G]���O~�!D�>�bH�%n�$�h�G�<�����<"a(�#���q[�Q|y��v�Lh ם|��	��l�<J���#�t]�G���k�!��y����������� �L;-1O��� �̻�p<�OWL3��aC.A(e�(���X�<UB54�"��f%;Ť��S�^�<�s��Y]���P�
"E#���3�l�<	a�'p6Ș��^#w�ޙ�N�Q�<�+�,gm�T��燷� ���[T�<�ǍEH�!��&P�[����QN�<�O��ϖ|��)�/{�����CL�<�I�МB��V�?*����(	`�<	g)��1�Ɓ����<���J���K�<q�/�0R9.u{��46Pb�"�A�<������������q�fz�<���ȣ l�Z��.O@\�`��}�<0,9�:�km�$\$X�%��B�<�k��}��!AX%bcN9��
�F�<���L'6ɠ�ud]!K%$���y�<���V��A���:P�q�b"�u�<� (|C㤜:/M�`oƖXC&]
�"O����̂��DI�.��L�e"O�ܡ��"1r��$�l�ڨhb"O� ���6@�uKM�*�l�S@"O����@�4�ȕ�A����]:s"OZY�'YA�%��E�:.�@D��"On�z��όD�Haj��8�V��"O`E�J�%U�Ω��Ε��uIS"O�R�d+�!yP`�θ��"O (�Q-&���3WF��s����"O\�#"	Z7I7�4�`�G���p�"O��������!�n�@�P I�"Oa���sM`�	�m ���T"Odt�3� ,DEM����4r�Z帒"O�UPUHX�Lvl�tR7~��0"Oh�	��TV���E�ڀ^�J�0"O�`��m�n0IT�W)84�R"ORD�G	
� 5�C6�A #���"O !x�-��!ˤ$
�C ����"O�ȃR� �8�\(Qk�=i�\[Q"Op�.7k����)\: �����"O�pA��܏0�fT��I�&b8��"O�l@C�La��*�n�,��ae"O���oO�!1�y1U�
����`"O��Q1�Q�-��AVl�k�]p5"O�0Y���a���4�\�"뾨��"O��(�'H�Mx��!�+;]3����"O\�a3鍔+���,�H��4��"O�@��$L(�`�Ȱꆜp�X���"O(@An˳9u!�)b{��F"O��7%U�<��B)|x,d"OZ ��[�l(����͍}T�iB"O���LȳVBHkU凓n)|��"OT���&BlΩ��$�d+��2"O���AR�/�` p펼�̀�"O��+p��Tf��'�� M�E"O<�!/V�M�� �$4�F)��"O@����SY�A!�Α�6���R"O:l�@#Z={�D��2-K/n�P(*O�m� *ϋ-�H��6�\5t�LdHӓu+�Q�N�9Q),��B�(��PN�C����&N.m6��ȓ`�4�H�&#W,݃��_�m�ȓtn�C��̚"�U��%�57�~8��<b�)*�Y��A��%�0LB��䪐9q�^�K��;@��+>��ф�m�51PE0q�����$.�ԇ��*��#<�P.&&�2;~<#�j� c��@Gf�}�Q>��O���+�	_-L�6���ܯLƦ���{r��cRV̇��,j`�aeI>�b�#aL� F&��'}��RW�ؚA�N8�'`�O)B��>sb}y���Tt���j�4�?�#�G�@UǊ )���)�>:�L���3T|Ѐ��?8qN����m|4Ke�G�8+��ק蟶�����6u��)�0O��Pn�d�Pe���h[�j���S�O�p��+GF%X7h�"��#�t��&Hk≒0Fa��oŉGI��C����=�d5rT��6L�T��'��5��#jǴeF�ܴ%����	��NP����~���N�ΑxҠ�NW���(O�>%xsE [p��w��*qv�<HQ�K7VTh�%Ǐ|6~�g�l��ym:�'}BF �$۹(fz��dG�x��D�7DD�:A���b�� Ot ���	T��,�S]پ�C��ЕX����Ǉ,}��م��=>Y�E�ϞK}~���)�^`�w���,3���G��u)~	B��zv���"�ڻ~�.4S� 5�>�$s�-Z�B����|��t��-�3�"%+Ͱ�j��Q�r�B�'B��i�Y6��wJ�"��N(�t�u�ػq�&$�=E�4憡 �3C�˚0�4��#Jbl��1�Ie��~��(����_)+vi{!Ҭ�y��ߦۚ%�ՆC�$6��k�c��y
� ڑ�c#�^���D��q�RP)�"O����n��񑌀%-�l%RQ"O���E�+PJ�E�F�8ي�@�"O,�����/ެĻ�/\�]μP�"OL�0��_)}���4.ӜK�U;T"Oͩ�U��R��R.Z�Y���e"O��s���U$������ͱ`"OJU�P'���� �ԟ��P"O�H��S�1�9�g��"���R�"O@	ے-șU!^�xs�C�z��x�"Op�oT�5�<K��\-"x�Hj"O��k"hJ�%*0ɀ@�Zdp#�"O�0Û�b��5o�/
,(,1"O���'�B�̱0nZ�=/pE�"O����U`��ٳ�^���c�<ٰ�ϦUg�) �Ƃ�s�33k[E�<�.S(R��q2��2F�"�2cA�g�<��J�L���±%�J�A�'a�<Iu�=g��5���1, ����[�<�!m�]�tP	��
�1h|Q��d�A�<�b�
.Zi@��!���l���`Sh A�<�&�4d	L9C��2$�6�E'�}�<�Qk/i�1ER�j@5��!�p�<��C�gڊ� �NON �4�AU�<�t�Zbq����g/[r����M�<q�C����U)%�V;(Z��Kʆs�<1DlL�E[�`���8A�4\�d_s�<Y�*�]��M҃eR4ϼ9#G"Pm�<!��(���j��ڮl2ĔӶC�t�<��<.��$k��M�,��OAq�<S,�v�|��F�7t�\D��!�G�<��kԉ{S����é&p6�P��E�<��a�9��gH	����	�f�<ɓK"k�Q��0aZ�y�֊e�<�C`3(�0��� .6�.1��B�g�<���W� �@��L(#h��:��c�<I"N��N0�E�APB�&I�<ل�_ :̬�2���MF�q��a�k�<9A���4�r�Ԙv1R�M�j�<YJ�F*JD�}ߒ1�
��yr���xA���OLK�CD��y��E,��p�
�+1V��2c�y�m�3�%	>nx��
U|6��_�����(�5rE4�6��]ʘ؆�;3L��B�с����$"H�Y�~T�ȓG$Hݠ�E�� ��H�dǇ=R�=��~Q�H��#2�$�"��8�LІ���HH_�i�<T�@�ݚo`H�ȓ~y��C��0(;H� �"J� �ȓ\��%K���AX�l�D+�/��ȓ}L�(�KU]l�:���A����ȓgy#���ON�u�4N�Hz܅ȓ��a���'{�䅘�B�7R��p��V���j#�A,*B����A�--�̆�qZ"�PV/T�6�ܱ(��M��H�ȓ+윅"S	}T�x0���n��ȓ-~��q�o]�4mRa�G!A�@���ȓ����̋�n�Z4���>-J$�ȓB!B2���@�>q�2m;�Єȓ�@ɺD�0o¹1+��fظ��l~nPsw�҄Z�<�E� �W���g� 5�`���rM�D����ȓH �dÑ0ahtz��D!�����UL@�p�ꄮE�9���fB�e��S�? .Ȩ��D?}s̜���4��(�"O���q�J-Cv��$��5A^$� "O��@d�QfD���)D�r"O��{U��/!�r�3ċo1脲7"O����nϦ1�r	�(9~`[�"O��l�8��qH4BZ�	**�p"OD�)C�Ě�>��&ܹmt�v"O�!Q0��U�Xa��U�	ˌL�B"O����EX�t�PE�6��,��"O������T*p�F /ǌA+R"O�Й��ӀT`l����J4\YV"O\�r2lUL�q�#��d���	�"OFE HE]�ht�s≴6�z,�"O����׃l�|��b����� �"O�1�OS�2��4��X���"On���>`�r`b���~E����"ONU�TA��F��qI�`�<cA��@D"O��D*��l+�DJ�o�%m�n�b�"O��"	�S�K�2�칀�"O"�hG��. �p<bf�5ox��2!"O2�BD�G�&�V��b,[m��Y6"OXXA:`�KG�@:-����*O~5��OŹC�r���;g�����'}������0�W���_�1��'6�(UKC3TY�ɷ��U0͑�'6��#��?|��GP���;�'%DM��4a��0yWG�CGd��'m�RA�ʕ��!�� ��e��q��'#���4B�O���󰭘�^�8`A
�'�����f\+2����аB�*G�YQ�<� f�*,y蕨�g���Jt�<��"�(-4��U	��;[�-\�<)���|LZ��M���Ēn�<��@�0��bg�e�ؓ%Kg�<Ie-�
T�$�q�Dٯ5O�dF�[�<��b�T2w����X2g��U�<a�/��a���RX��@P&�S�<Y�j�31'a�3�޼fS�`H�j�<	tm�L��� �&	���@�b�f�<Ѱ��(X� �yU뉪A)p���\h�<�Q�ÈK&d"��F*/Y�-�E�Ap�<IE7ibA��n�ҼaCEl�<�Rd�s���v��"�P4x�(Uf�<Y'���V�Kh�
L��%J�d�<��I����j�B׽`nR��rf�K�<A�6�\���
�:��pYr%�@�<Y�g^:D�$2�]�;j�p���~�<I'R0!��I1��M�N�ӓF�s�<�	Bu��S�O��r�]��FI�<ɲ!�n2X0��|u C�oXH�<��Ț�2��ٳ��'Ub̴ʁ��F�<ɷ�J�+-��y@��"&d�q:���E�<	t�
Zr��5�U�(���D�<���>���'�:�)3�ID�<i��H�|���+`�/0�R���|�<����R��X ���p-��22ME|�<IpD�M�TYz5!�z�P��#��{�<�4�`�8���_7H�I�D�Bw�<!�)>�݈��G�T��#��Dp�<y�/(��t��!�pȱ�+�a�<Y'@�4<�!hR�E�TX�)B�Ob�<����;j}�(*�T�(�2��D�<������h�h��C;	���X�@�A�<	�A�6�v��T� �Dp��O�z�<� J��&X�,��|��e��C��D#"O��XP�K>7*j)�e����8�"O��b�䂺.	*4 �
�|��A�"Ob0��
����)sC��F�튲"O�%(�E�t�6aW�R��rs"O~)�Ш ���{��	"�2 "O<�����a`D� IѻodQ��"O���b���$�P�U1��e�C"O���G��z��3�I r���"O�X`� ����UJ3'��ѵ"O����R�5RaӇ�=x
�ً�"O͙�.Ť� ��fD�=�I�"O`����!,�^��3�C���"O�]�u��?5ԙr�e�I��q��"O؅�`�=fu� ���KR�x�"O�E�҄
�vOd�I��Q/3L���"O����&�7Z�0%$ן~&�u"OzY��F�?f���Lә!��3�"O�4��Ԏ)�lx�����0�7"O�a���T==��$	`H�v���#"ORd�D#2
��|�F��jp�T@A"O�a�֌�y�r���/HX4؈�"O*=qe�\SF�}���W�1V �q�"ONt�?<�6��bd]fn��0�"OfH��Ŝ�;\,(�!�("�&��%"O� �LW�%��ئ��D���c�"O訉�g	��ݰ�l�+H`� "O�X�l�4��`D-�.	پ�{ "O�T15ϖ�8>2���ڒF�69�P"OF5�Fm�'_8>��3cV$���"O4� ���EJ��K�;�c�"O��ر�Z,Hv��F��= ��X�f"O<����֒B�va�K9l��M["O�rp"�7��a��4"����"O4(���
o���D7j���"�"O�a�L��XT�#�نP���"O�qb�\�O=��K 8���"O�x3��u�V���@�f${W"O�I`-�1!|��(�.O�X��\j"O
U���9|����J����"O�Qw�)���
<GI(�V"O�����"��Py��Z�b9��"OX��s�ʿdF^��B�	�av�d"O��S��X�������-'�~�sF"O�u㕀�|x��3����!:�"O��r���7F�]�d/�'��`q"O�X���^�Y�*9��QM��{�"O�� ��BwK��Z5h�	J���"O� ڢ�o�T�Ȍ2�!�"O����n^��8$f�4��e{B"O<���'�H<xHy��ρѰQ{F"O��ZL�+u`H�Gk����"O�����ð��\�@�"�&d�"O&9AS�]�1}2`{��I�-�L��"OP��tf@ .��ktH�&i���"O~��4ֲ`؂e.��р"O�Z�䋰E�8�Y�_,����#"O�i�g��D p!y������1�"O0��޺2�=�����"O��X%`\D�pbHNv
h8�"O�U�U��p=���D �2k�LRC"O���A��O��M�tfP<sn��"O��^�H*�-��C�O� �I�"O�e��̞�6~x����R	����"O� J�®K�o�J����"a����"O��X�@Ӥ���AEvn���#"OF�`"o��_����c�9%��Iq�"O�Ii7��I�T�7�0I"m�"O.�B���8=x� ���;IJ �""Oqs�	   �P   !
  �  M  �  �(  1  D7  �=  �C  J  \P  �V  �\  9c  {i  �o  v  D|  ��   `� u�	����Zv)C�'ll\�0�Kz+�'N�Dl�����>O�9���'X(�4g�#-`�1W�'S���!�
L�t"���e��V9��͐Z���2�aݹ`���?
��R�?���C�m�� �A�l:II�kɹZJ$����^�/�l�"g㘎(Ɋ�kw����uwȇ�;�T�'���j׈�Z|@�Ӧ�ƶet �뗠%�t����Oj���ҝOF�����Ǧ! P�B����ߟ���͟(�H
k
�`SgL:2�D�
�����I&9�(�۴��$�O�Is6)�&�d�OH�P	G�`�������V!!�l�O��d]}�Z�d�	D]`�$~��	�5�"�qE�c��-[�+A=g|q����<)%���QQbȝr�Pk��y}"=O��TQ��]�*�'���W.Q�}=�))R�IT������?����?���?y���?+�d�]l��鐃�݀l�Ό�&�HR���LȦ��شS8�flb�x��Ȧ�	۴�?i��i7�Ã6V+]jQ	�IYV�"'`�s!ў����S�T�HZ��F48�d�FFQ�8a��U(��=(�óaH�ne�m��M��i ��c�I�fTVE����u����d@��
M��y2jX��M��d�8�ɐb"�|�k֤T9ِ���J�U'���oӪm�5@���b����s��U�5�%�*58�j'�I��Mk��i�.7M��B�:Ĥ�G�JaQ �	�*Y�M������-R�A��f�?�|��˓�il��QT�qӦ)nڗ�Mà�x(gюUL����Ͻw��P�dmUS6��yAn]Ij, ���ȏ�M�#G�֩�P��(��9" ���?!�(� !ӖP!�B�s��t��t��C�BzR�'GR�O3�$"Qs��x���w72����'Fh��e���݅"+!�dБ+�"m��E9~b��kE��%�!�D [��٘3MЖ3\8� FL�7�!�D�ɮ��̀�
�*�I�>�!�S٦5�%"վ�}j�J�%`!�DS�7���y�b[�4V���H^�Z�ў(c2�C갍pt*���y��JXO?�	�ȓ2�&��6)K$z"L���N���ȓ#z�<��$]~�(��0��ȓ
Nz4H߃*��bŬD�����[��P�5�����h�X��ȓ8 �`	=g����u�^���Q�8"<E��ʵe�NA��P�tV��0bчH�!�D֬
=�X@@ K^� �`�� �!��p��|+���d?��+���V�!��2Z�Ԃ�c�h�����!��7�^PiӅ�X�:س�π0>z!��>;d��(�CՊ"ž�4l_�I�*�t��DȕN���֨��ؔ�F�ʺ0P!�D[:rP(�^:`����싈#!�D��:n���\��B�K��G !�d��h��m��OG�_�j-�wO���!�ʸ%��M�!^��5)E��yRcB�7<?q��R]�T��w�ERѲH�5J���p�'2�'�����$�eapFX���=�-e���AO'�rpx%�ݺN�����OT�'ߎ���YN˼=+5M�$Q7d4��@�̘2�F|&-Uj^�VbD���`�R�'T(A��?�#�i���W^����N�18$�2_��	��qc��'n��á�M��~2�_ +�ة��ut��#+����'Oў��?�u
Ѓz�6-#����~�)��h���4�'I4e���'��P���s�xϓ.	VY�7�25��i�яB�i�|�'(��e�Y�S�O� ��v��S~vy���?��!��Ox8�+J�������(Wn
���$�mՅV��hG���YBe�Ob��>�i:��A�dlˠC$ِqr�F�/U#
�O��>LO\��gW;w�
�:�`MKD������#�h������5���	� �<�&()0.lӚ�d�<Y1M���Z����i~�Ż�����B|��%P���aP�`lI q�L��W>��S�~��"�T�vl���,�����@�^�C�M�U��I��i�K�%(ƪ��rr% �*y����{H*bP����04�ߦ!B)O4Hf�'�1���'�r�B3l64	 �
t��KłK����͟ �'
���>��F$9��*�+��*�<;�F[yB�w�Xm�r�i>��}y��2��\�Δ������C�vL]ћ'�a|��p�40ӄM�*1(t!)!*Z�Q���'���Ǎ����ÁݶY�X,@���7�x����c`K!�^Dz�	��,����x�W�DRRMS�(X/N�B����9�yB��h0�� s�3"!@�*V����]ޛF�|�_k����jt�T
V�Q�ڠ0��;U�d{��'���P�Iʟ�g!Z� �F7FĎ�����n\q�? 2�1&�߄'v�{��]�7D|Xq��>�Wpzȹ��9D9v�H��+MdM�F�� K:J��2�D	J��X��ƣ��O"�(��'����`�R��rI�RLBV�.,�n0���O ���!E~�hSgH��8��P	N
�R�O
�qeG�,�@��h�9����2�'J�ɫ	t"���4��'����O����#X�!�x8�RK����@���O@��E��
h��*t�p1���(՚��~
5N��w��I��}�d��d��d�3��y��Ğ,ѱah�0���?U���̄@�(A�n\$K�B�+?i�d����	O�OM2f�?
�L��2�;@�8š��FX!�D���N�0#��&
�Ƹ;B��A8џL������}�Ta��Y(�4C�	U����$Ó~��i�O��$�O�W)X�s2�L6us8D2䜭i�R� ���+F�T�L�ii�E���i���$�#%.#&־}�6ԫ5�@�-Q�e�ڰ�_�^�������!��c>���懺��d�# _�ܪ1iH;sm:��4<++2Hj�.���=���$:�<)��%�h���}��B'R�1hĨ(O�=ُ�ӖE	<�:U�D�N������]��Ϧ���ןx�ܴ�?Y�'�?y)�"����p�X�@�5x��6uol�$�O����O��S�'o�u���Y����1H�5�f��e�FeYR/�KWR�F�W.Oџ�����-ND1 ����:7��l(v�r�� �����
�J'(m��E��nQ����]������-��C��P�_�j��OZ� �	n�OP`�q�	�lA �-�	B��5��'���� F��E�k�@���O>C�i�r^���������	�O�����*F�=�ǉn|�@���O���W(bp����O���4�5C�~561�D)�M��B>o�z�@w�Z�?��)T�PR�4��d�M��dؗ#�e�@D�ڴ����1�K�Ex��p�ʚf�.���0^�$�O�Y�\�(�$��%�X t���$�@�	A��4rW�] d2f4Hծ�-)��*C#�O���ɀI�d�ʡ�Kqn�E8Ķc�>�d�<�Cb�3ߛ���5ܴ��	����D�k~j���L�BC��Cǁ'R�����O�!7cùf^|�(kv�� ������?Q�3L��P�R����>���J��+?��]e���{T�I�4&@���C�J��ӸB����Q��1Es�A�ÐR���b���	��%?��|�T�68��(���א��Z��KX��ӟ����4a�H���b�#xBD��td <t� �?���mK4�z7�:���V�S�����<�l�3�H�zA �$�0e��|�oG�5��Ɇȓ`&  %*�7n��E:,c����e�%)`.@�n`��!Ú�	�8��eT*d0���?�hq�g�[;H ��MNB��M��L��ʐƔ&����e׀���ǒ�|�*�Psg�shY�'axP��%���M~6x����u���uN*@�H1X��G	� ����Ҏ�9T�d����+R�~vF���G�z����!.�9@`��>W
�ȓ�zX(�"�:UB����<RU��	�-���	�I��Ӄ-��Gm$<�D �.B6�C�Y��(ݲ)�|��*9�C�I;U��0ӡKS�Ip!��@e�C�	�:]�Q!�!S4���t��Aj C�ɩ!b�������+��)x���O,�B�ɽ?��ԙGE1*8�Y�CO�2�=i� @�O��I�R��.L�u���F,w�����'����M]� T6�`�W�;��0I�'� � U�ԭa�%0k�`�����'b�Hx`((U>L��*ϼE���'
�s5OVl�{g[
D�ź
�'"��y��� M/:`��ω��V�z�H��Ex���MiA*�0�'V�A.���v�U=}�TB��*����oX?ʤ)�%�h�.B�	n���tIZ ��+Q.бf"B�{�U!#	���V�����TB�|;�q �oP$'6l*�k]*��B�I��%aѤy��9ʕ!ߨ��p3�\�h��(�O������bW����+�,��"O� ����řp=>�����i�&��"O�hp���<qP>���K�  %XP�"O.]Җ ��SP���j�j�5��"O"�2�
�/r$�q'�ɮj�#�'�D��'�|xA�`Z�Q����&n��z�I�'f, c���5=�I��G�:O�pX�'���AkC�%U��^#O����'�I�v"E>@�IzTL�DW!k�'�
�UᄍB��C*H�-�LP �'�T�5M�q*�) :Z���䉉y*Q?�3m|�p�!%�&�y�!�DC��5���h1��1�����j�C��F�� 执&("�Q �C�0����`ʈ�,	�Ay=�jC䉔s&^i��B^����i$,*��B�I3t�()4�_}��R�c+���d_-=��"~"�!��� ����O�j&N�Vo�y�Muߠ�r�.�s	`	����yr���h货Gq�H��J�yB�I4S<� �bۖa�}�a����yҥ��Qݒ]�d�^�R��p��yRM̲��1ƛ�H
�ʥ'6��$ӧ)�|ҦY4)�� @t�P�	$)��&��y��LY�x����.��qP��*�yᓬ]"�x!���%,�6�	Q��y�+R%"�s5�G�̀E�`��?�ybbD�'1vYh�h�Q"�=8%����>��"�?q�%��i���>1���i�i�<��6x1%[�u5JL�d��{�<ᵋI�QŊ�#,����%��k�v�<���F�Rm�<����B�B4Dv�<�0lM�27*�@��)�B��Hq�<!��
i��}# ���  ´s�Um�'J�QI��I<0�^�ҧ�� X�M*To��H�!�D�9)���
��D0aW�IN:!�$��:�z�0�N)e���B"
6!�DБax��$/�W{��
��I!�<t�(��A��3m�` ���o�!�$�A|�=CO˚j�<Q�"�t�2h��O?񉤍̖-G>U:���*^Ȫ��@�Bx�<AR(��*�n�����e]�%*�u�<A�A�U����v��S1"�%�SI�<9���o�`��G:L���!�y�<I�<�L��m�]�Hl�3K�\�<�"b�c��5e[a�04���_Yy"��+�p>�TmӅ~��ҵ�K��8��W+�Q�<���>�6����0�2�@NRG�<YGLǪ�u�Kf��� *M@�<�D�F7 �t�{Y
�B礗R�<A��$���z��B����[tx�t)3᤟�*���-� ����� p�V@q7D�Ĩ"�!r�x��h�%b�LL딪5D��C0R+h+))CC�<���2D�d�a�|�2,K�B+,�:�H��1D���Ę5�.$Y���+�¨c&1D����+�iw��o�:q�|rV0ړ?	�E�4��cӬP�*�$^�i�� פ�yb�@-�����%E���8'��yڬ, ����D>,A��B�d�!��E�"����ƀ1 Mг�8ro!�d�7Y��r��>5.�����A�T!�"t\dL���ך7�4���2+2���O?qi�NS��#��?CH�W�k�<�v�^1j�,�
ъ͢B��ƥj�<� @��F����K���OM"Y �"O(��L�8:t`���.L8�RP"O2���E��*�Xr�10�&Q�"O��Ȓ���D���DT�7��u]�|�p�-�O��)�`g���ä�x���1$"Of��� A$m;Ђ�L�����"ORxzC�,�X�&b؈�T�bW"O�=���/6sN�[�S�k�ؤ"O�a�e?j�)$�������'Ep�s�'޴��t�]�%�D���ΘV�=��'u�@��)�dl �	�${�%s�'>&a��'�. ��ʣ�@:Ȏ�#�'�,0	a��Tʨ�jd��Q���'hi*���Q�r̞yIZ�'Z�,)�c��p��!k�wCm+��DO�L�Q?-e�·qE���ժƿK$�$���"D�����P~
p���B�.߮����:D��r�K)�6MB�ß�T
�� c9D��#�?d�x�
�������*D�Ї'ޯ&<�I����	��&D���Q�C;8�Ě"G�:;�}Q�e�O�	Jt�)�!�P52;X�"��K*L�� �'�@�#Ϗ9�x(q�B�T����'޲�bGe��2��	B�J�5#����'��!w�_@�����('�vU��'��Ƞ��Xh�e�6��0����'XD�Qv� .J���6"��z�+OF��t�'���N]�.}8ѕ��bJp3
�'\��c2g��y���C���'9���n=���HS;:!f���'-���?a|�aVI̼91�P1�'r�;p��!��6NM6Rҙ��I�,d�D�$2eLA5I;B�:��K�1��a��\���͒�E]2��0퐛 �,�ȓllZ��PE��Z!l����a�� �ȓ}���i�+��E�@!�ş�9[����1#���#LʠHd����'W�d`4͇ȓ$��(%LUC� �!��3;p`hG{R�VϨ�����Q�Y�"ș`nL|*���b"O��Pg�U���m��k�S����"O�p�������E�Y
/��j0"O���4Eʊ7Ti�j؞}��h�G"O�����C�5d)�a)��+IT�à"O2]���>J|���^�03>���'3�����3u(&����D#�~t#1��=����a�x�q�Yz�6q�C�Q	����a��֩O x��1��j��*4�ȓ�̐����Px1c%��[��ȓ<e�f�9y̌(3P�W>6v����]6��3�^���@��Q[
]�'̆�s��L�t%D5��{�-��d�ȓ]U�h�&$N�i�,�Ӎ�M|v���R͆9���12����Rf�)Cީ�ȓ]�$�a�$A�qu�l��G�����=D���Ö=&�,1�޳8Ll�G�:�O����Oa$i��%�52�X9O^%X�"O:]BE�ڽ5��m����J�!-�!���Z��(VaX+��`
ђgK!��ى
�؁��+c����e(�VC!򤒔%�z<��͗�R�&	�VF�8VP!�dʺmWrq�Te�K-24�T'صzNў�bE�$�'e�>A�P�5(6�K������d劓�[�.���fO�o����ȓRG���ᛅLJ8�Tb�)І�S�? v)vÛ�u~�իʘ�� {a"O܌�� �oi�m��� (�)�"Op|�wA�e��PA�C�6�eR6�'�Ы�������Q�&^(LRF�#�ƨ�ȓs����C"P�&d=" Z�0����ȓXNH�Zv�Z`y�0��.�Lt���	�Ihd�Q)w0�V憟7��Ɇȓc�&|+0�[$Rp�����j�4���"dhI�B�v�������'�.��'�&���oh�UA��\�jUs���"�ląȓK�x|�$�f�������ȓjFl�vnQ&�0}�KV>S���ȓ$Ǽ%��.֋7��d��gV�:��a�ȓ4����C��W'��9�d�694���	�F�H���؈"�4ls셢�m#B^B�FW��K��eܑ��Gݘ]WDB�ɏ.�tc�a҈p���!���B䉁z���˧C����#
�X��B�ɳn���*��_<\CH �A�3n��B�	��t��
D�u,��%�i��=�u�YH�O[L1�Fn������3��LP
�'���&�M�p�j���eTyL.� �'B*0)�nU?Q���a�J�7@̨!��'� ��/K�W!R�҅� 2z��Z�'4Jڤ��1w�4��#�r��'�MsU�E���X���?!��)���(���Gx���U 1ذ����:��l���q$RB�/�թ0M�3��|���ѲiC*B��s����|^D����H0
B䉗Z~��-�8�X0��a>��C���u�B5a.`�U��TB�C�	>6��iO x�JYX��&���I���D�O~�@�8�dN~�b�?R�\@+D���?��{ o�;xK�	�@�	�l	� �J����F�V�����4�������z�A��}���3%Ң�O��qb�*A`�h��փVhD���'V�$����$ +���U�h���K�(O��0��'����\��R��կJ�e�` �
D"����Di���)�@<�c܎y�|��M'�O��'�&���`�(�j�knǦ� .O ��o�O����O�ʧ&O�i��?�h�3 L�!��
	f�!�
���?� 'I�f�T ���K��\���' ���D�'
���f�Fv��B��D(̓I�x�`�b�t��(�o	��?1u�T�&!v�I~�2KY�>�"hCx�LyR,��<у����IX~J~��O:�NI?0�̣��,UQ���"O��ZҋQ�@�t���M)W~Ձ퉋�ȟx� �c��1Z8ɂ���Z#rg�Oʓ^h�$[���?Q���?a-O�	�7r�0AE�" Pl�夃g�B9�Ad�� #ɑz�B��cH5*��
�&Q2��AM/8��S�@bɈ�a#����q�L�h$A	͟5B�����Iu֨PC%�Ƽ��<XCJ�X�T�z��	ԟlF{�9O��3��4��}�"�0pAJ��"O\�U�Q�֋��
4:���K��?Q$�i>]�ICy2�bs`��BB�W��z�Oߤc*�q��)X�1;��'���'����'+�>�f�Bs�K�!DT0
��DI�ܕ{@N_I�����*�3#)�K�'w��pH���a)@	a�GC�aZ�m`�hZ�f:.��"�V&3��z5�ߟpce�_1����?6C���4#[�9�`�s��4|���'!���D{��ɱ2��b�89�I�N)#q�C�~4�QC��}ʆA��K��{*��&�'��It�h�(�����z>Aq1d�?��X��%T:p&�X0��O�8B�(�Ob�d�O:rCF8s�N���"FOH�	�u��5�P�I�U���2�A®��O"�%���H�����L�j�����R�QJ�H�'F���f/ �2	S�ּ���܂���OL�� �S7we �����*��!�d�\'��ʓ�0?�Q��"� � <^0�I���kx��.OP�A�O,q��c���&O �p�^�8ˆ-�����-���O�� k��O��(�"-H��$NA�@�~�[Ě�-���Jt�ʬ	u+K�%nɐ1��O0�'�OQ�a�^�0��e�9�9��'q.i���ާi���:��թX6B$��j����6��,5YNl������ZW��y��ƈ�?A���������� ����O�p���P#T��2Mx�"O��(�j�	L��Y���\/;��:G��2�ȟ\UheC
(OH�wM)t3��ر��:)ɔ��3�-f ���Ҫx�ɺ&��Z����d\*�-C+���f�/#�ȓ.�� B��f@d��i�Q�9�ȓ$UXX� �*q������jx�ȓ=���`�/7���akI�8��,4
G�LҙZ3j�V�l��	�>\����^�'��m�G�$V>
��,�<�!�˴q�=����6M���d)��!�\"e&8&�.D���I�$�!�d�#td�h�W�0(T����LC!�Q�J�����;q��[�a��:7џpa��D��M���t��>n�H"E	**܆4b�@�#��'��gS�� f�b;\ٗ��}pi�;y,����©O�>�����"�E|�f��Cg��	���=E�Z<�1�[>�taK|0Y%L�?��<h��=4|$�D���rhx�U&>a2�!���VI[Xq���k�+��KSR�'��ON�d�O ���<1��sz�P�_,��Ģ���>as�i9f6M�,!��d�3e�>��R�.]1����?q���?	�����\��+[�k/���e� cʥ��-�>y��2�����F�y��DP@ᄯE����?�ݴ�ē[h&b>uJ�N�'cla����z�Z��6�8?�b�OH��Ɛ>��y2�S�
��e��G� 0V��Ϙ9D;Ja[2����O����(}RL.�X
����[&G��2q�]	Y��!xJ����'��>�I~'��g�]�t3E
{ ��g2}2�7}��ܝ��	���I��[T"Qx3�
D���C�"��(�R��.P����K�i ��K��Q�Fړ��?Q&�_�$�X�䏭M�z����E��"Eأ�Җ�Y�J���$K���"�����0���6.����e D �w��l�O�s���֫"?a���y<�I5C�#{x�ps���3`~�'��x��O�����	��L��!DԛL�ؔڵO��BH�b?�&�Tn~ʟ�^��DΕe���+Ёm�Ѱ�Gлo����j؟`H����M�<Дh�,}׆ A��/D��p3��}� ��ʏ/1P.!(kn�j�=E�ܴ��!�U�SZ���	�i��;y�(�'���'Y��҈1nA�0�Ӿ[e�@�E�;�!�mA cY�y(��c��.!�dMm�L
� Yo�|`c�d�!�5����$b$_(D,js'/g�!��F�H���I�	�z��L*#@�O�!��<hw�(2Ԅ
@���@�����' ����m:�Z�`]�堼	�'ҬR�)w��U���R�!~���'�>a;��/��qy��Y�x����'@��qq�T�x������D%vݒ��'9����	(X���l�'Wzp<i��� �S�t��':��AEP��йL]��y��t��I٥�[�v�^��c����'��P�f@��#V�-z���iM���Q+�cL��"���Rcq q Ǿz��r��	%<9Jt�H�K�O
)m�F�����~��A�ʤN�| �U�;:T����(�XkG�I~�����<��9�����|h�d ��;H��-�SЊ!Řm�@B�G�3W��c�4u�E�c@�}��:6��9c2d�B��'f��Ѱ[�	5a޴"E����GaD1����	O)�<}p�_�w�����)�'���[pK�C_ UP�н8f����s	��¶L�?�!�) �p����3��.<�5ѱ,;��	]��'.�O{�O�\�7��rf>����/`�s�{�'�ay¡L�4*�x�֢� �FT�QĈ"�p<�I	�(hK�	� s�d��4[�L�	��@��		�ިH� T9�@kA$�&�XB�	C Ph)1ƕ��Z��V�V��B�	;���A��4T�yc�Қ-bNB�7I&�8�
�<'Ś��)�7�lC�� VTf͑`OG5�ƨ�i�i	�C�9T}P��g�O�R��[�G�� `B��(%���cP$<T"f<8�g���C�)� ���ʂv/�K� 8�e"Ob�
q���M��cU#~zM �"OX-bݩ|�l�aěOV�ب�"O��XI�$?U6��p��3Epu�U"O��(E�Q�J�X⒥�r>�i��"O��" �Q7X�z���$P9"O��1*R��������$.ЀP�"O��`g07���AǶq9�]C@"Ol(���VP�+������"O���4L%0>����U��;�"O~i�������zC!�*R�2`�s"O�����J�)`9�o̚	�6-��"OI��i
�(i�T��.��z�z"O���b�;g�ެ*"��
U�@8��"O�x�t�P�X��DR�+g(�z2"OnU���κ�i�������W"O`a!�/ O.da@	�=H0k�"O��c�,E���E�X2d��\�"O��Z�	�)�@an+X� L0f"O���
�.LJ�cQ5i���Y��I�y2$�� � YS��s4��S⇃�y��'8�@�c��J_�z��Y6�y��Y�� 9Ũ؈f�N��g��yr�EFn6��t���P�����H�yҭ���1��õL�r�S G���yb)ͤG�e.�26�0P�'�ҵ�y�=+s��� 7]�anM�y(��w���҂Z��Ёчȣ�y��4^j��q��Y8������yR�řnJ��X���kBHT�Us��ȓa'�$�"9V��`�$l Y��n���%5:���c@�AWtΤ��.�P�)Q�M���0��mh~Ɇ�<B�=0��U0���O�T�ڹ�� �~P�O�/�@�[玊���ȓ4"Hb�āub,|��F0>|l�ȓF���rר��nP"�)�LUlD��ȓ���a�2�3 ���:��@�}�&��Mn�l��ALvBD�ȓ�ny��N��=@q�������ȓX|��R��59�XQ�T�Z?^_6P��|����J̏H�ܤ��N��͇�P�}7H�?3h��T O>����ȓ2cHE���J,��[6�~Ȇȓ|�>�cѡO:���CaσN��ȓy�Pp�F$��r�ᱰh������j<̼0񭉃�șeJ� �^�ȓZ�]b���+�`��S�
����@*��ݥ��t�G.ӫ(���o(�ڡjK�D���%BU�o�����t�� ��� A֝�GO� _Hp�ȓ8V)؂ɋp
��9ba�W�t��e"\���@DB�Q��Uo���
��)�C
\�j��R-0���q&6���G�4zU�P2���w֚���d?��K�ńVs�Б�$�/}��̅�$ߺ�k�)jUy�ÇMR	��>������ ֍i��Qi�P��ȓ�T�"�b!�mH���ȓ-��������~%x���!2A$�ȓz�1�.
ǄŃ��D,/:X��<]Z�
�#�+A���Y�C� O����ȓ%�����&ô�qQC'yx|ńȓN*���oٯ#_F���$�&|Rf���S�? ��B �Pj��!��(.�4"O)8V+�8|�
X�1t��"O �TIE3��|#WϞ(B]xh[�*Oh��%�
�v1�I�'�X���'��y��@=L�d��`ғ
�Lhh�'[P�UgP�B�%k�O�
j$��
�'�.0a ��]��Rc R1,B�'�`�߰T���o�-Kc��S�'<��� ����a��؏M��h�'�pX;$�Y�'��JO��a��	�'j��ID+g����&��)E�~1a	�'❫�ٵ@w������:�y*	�'��yG�^/s�����Ւ:rH)�	�'�8�2�Eޮ	�HT���M 0>����'�D����'@����_�*����'즈�s�[-0���.�'r�I��'�h��b��k��2#cRm����'v U���n����" �0b���:�'�|�1tIF�>Gμ� �"1 �A�'zB��#�^�=�h)!#�$HZ!��'��ڇD��L�1sf�� MꝐ
�'\��dA2��)3!��#� �	�'���A�h�\c^xI�m�2~$I
�'��x�1|�F,�˵�t�i	�'%�xq��J<<��"�b��^�c�'e����ؽ8����X.^�����'��#g�z�8)g�\��m�	�'�h�I�jS@�����ߣB9t�+�']0y�!�,1���yd�F$f���+�',��óG��JTs�9e��X �'�V��cQ�`��"��
�a	�'d����N�h�D�`rf��Vl:���'��UGԡ���b�M�����'	.4b&T�V�v̫b��Iy�(��'&�	�2蓻b9�T�G^*B0�I�'J���b:h |���0��'4�-	ã�7q��Q%�*,S��	�'��P1�p��{�y�A��Z�<�e%�4�����"��/���f��_�<	1埦/�Ip���l}�@�t�g�<�v�ggڸ��^I��9+c $T�*�*�y�̳tM��̩㣯5D��0�V>
w�*�@w�����5D��
��%2��٢%�#7D� � e[>=���R�u�f��d!D��3��M2B9��Q)R|�H=D��rT�A's�i�`�TUw��9D�d�p)XR�ly��'U$L�)���<D�(�C���<t��ױ����d�9D�����l�vax�GU6�tĪ8D�P�Q�ڄ
�8�ӧdM�z�p�
Q�7D����,��$���A���+{t�"6D��qĂV�4��Ѕ�,-��:��8D�@�Q�6yD�2cťW��4� �7D�4�s���B���?����M6D�\ر.�- ���u� �yX��3D�䠥b��B�4-)@
�(���(3D�D���;x��\q�if]��l2D�Ē0��ypIH�:J]�ԭfոC�� ��3$�):B��7s>B�ɢ|_�$;qI
���Ȥ�(o2B䉐(��x�뎟��y@�ꑔejB䉦��Z7�ODw��rQ��
No�B��\D]	 o=j���:uD
�;i�B�)� 歓�E�f%<\Pt-ݥ1q���"O���&�	�w������ÿdL��[�"O��ԌZ=�Zb`ŉ�2B6l��"OV���B6,d�UE��W
��2P"Oբ'H�2K�����

�ԅ�"O����J�@���l]�k��m��"Oy�A��b~y(2�y�R�3�"O�t��)�g�bd*̆>�(���"O&,(�-5��Ⰸ���~0r`"Oʩ+����������h""O*��tg�	�K�z����e���y���ĺe��!�p�\�X녜�y�F��Ht�а����b�|�  ��yc��.�\�'cܢV]D�uLƛ�y�9F�I�K��iф���y2��c�b���B8V��w�	�y�i��l{^����_3�@���'D��#�*Bw �y�J_"�^����7D�4����*d`�D�R��;j��d�4D���CV�(+��kW=}��{�#=D��HRʀ-�<���-�S���1�E8D���p	T	[+�(CI5{G��� /1D���iC$Er�h�Ŝ�c����h:D���Who�4�s�cY6�f(�%�$D� �gN��!��0g�U$D�V,��F!D���T��Lo�U�ŋ̀4�J�B��1D�p�pA�-�� TEO�\@0�*D��
�g]�O���r2��q2и'�(D��Cv�B�;�];��<[�T]	%�$D���qa�1����GCƛo`1���#D�|�v��&S4)�B�t�*t�#D�,�VkǶJ� P�& ����%'D��p� C'��}a�܂Gy��	WB*D� �����z�eN89��b5�-D�`[3A'x���j�6�$�t�-D�ز��8*Ɯ��j��h��Y��)D�<��	�$U� ��� �,Z Z% 3D����hU�R��3��=i�`�*/D�`�1�5Ԟ��4"['%#��Ka�0D���Qu!R$2`��5̐�`l-D��
ŉT�19�M�$��:rp��e.9D�����ؚ(n~�I%��)m2}�g�6D����)՞8O�t�c�D�Aq�)2D�xB��p������v��b�1D��1 � B����*�Z�L+d&/D����T�G��C��\�09D�p��&���ea�6n,�J�B,D� ��Һ�����8�1�&*D��ʔ�Ź^�,[���*ے���*D��B�m 	���`"\�)��D #)D�(R�F�G搙����3K����G4D�������3�x�(��٣ÒiK�.D�,Z �̹�j� �LKa���3'&D�|Z�;� �ڐDW���d��F$D�lB "	�9�P�X�B9HàL��yB�D�$�X"Łgm���Ǻ�yR�������4g\�0�����y^ ~����iƤ��D���yb�Y�[.�q�,K`R�aڵ,T��y�.�� -o�џ(���g��y��ճHl0� D�m� ���敏�y�j:NrT�b�Ql�h��%����yB/.+�x�r�%O�b�ԩ*��5������9gr*tJ��L�y���*������� ��p��H�>�y
� ��%�ƒT�⊖����"O���C�1L����Rؤ��"OH-$�8&���2�N��Q᎑�D"O�9�4(�	k����?d0Y "O�$z��>N��Q�D&�a���9�"O,YH�(]+S����s��!Bũ�"Ot����z�Y�"��>�*�2"OL��k�w�&0��R�s�\�3�"O��` Ԁ3��-[W��B�6��"O�QWhK/Ǝ!��#9��P��"Or��M4�z��bS�6����"OH�I���#YV
���D��~�M�"O-����3\�a�m��K� ��#"O�����##��+2�	G�	�"O�l*���3T&�pp�є1����"O8�;O�x����5.�0��f"Oԃ���I d8��$���"Oj�3�+D�:�,��I�jr
�J"O�1����h�1��A�@8��S"O�|��|��*�X 8[b"O��2��=L�� ��������6"O\���G���C�c�9�9��"O�����ʭ\��`#��>4Ĭ��"O�ڤ���M�
!�q�.5&���"O"�A"���t ��01#��	�"O��H�睥D�H�jB�L;!z�!�$	�<���#�R�/��4�&"��!���{�b3J��w@!��f�6y1!�$KNv�5%7V����P%�z!�� *kz2���=a'���G�9s!� 9r��s�ۧn����"��1m!򄍲S�Vt"1O�8!�� PF/�|]!��Z޲���k�E�r��9W!�dH�a䤘��a�'�=]͖Ѳ%"Ox �4�5z0"�c \�O�0��"O�|J��.Y(���8�ڬ�&"O�\ m͋U��<����6*�"OD�ӔjΝD���fR)1��"O�ieĞ�4��}I�LK&+�#B"O �!�&ms����-@,�ӆ"O,<�!OF�P����TvԄ�"OZ��.5_�l	9¯\�-@ S"Or��Q-6�0�E Vx�Ha�"O�	 1�C>O�$Qp�]; �~ R#"O���H�49�����BG8c�~%ۃ"O�<S����;ΐ!��I- ���4"O�ة���ve�=(�o��40�� �"Ot�1eҨ,��P�m�f hupR"O��`p�	�F�86��$%�T��R"O��2�3�,�C��=nG�-k�"O�0i�� ��Y� J�X ���"O��(Ls�;��A��9�"Oz��1����8Ԃ��_�<p���"Oѣ�N;��PԤ��Ao.P��"O��k�/�O��r��ٕkF0���"OZ��˂ �TIxu���fb\�چ"O�P	�?��!���E�^�z"Oj�j��P�<p��w��9�X��"O�z@b�{��}
oٳJ/�|1�"OZ�3�5v���.�.�\5P "Oȼ�D蜋d�L��N���5�7"O�E�5hմE�sمp.�E��"O�`�qm
:!i��.��(��"O�EpgL�r`��i��*n�t "O� Jy�T�Co���"��T��1"O�P�i�+T	�kա^��`{c"O��g��4��p��d�2+��]p"O:A3v)�5e���Ƞ��i�H��"Ox�K@�ҥtn����I1n��$"OKQ<o��-S&�SA]��_5�y�# i.�\
�|� ���yB��=���?`��tyR����y�K�O�VEy�l\' �T�Rb�X#�y�	�~�&��`m�	N��EA�5�y�&^>�z7f쀽s�		�!�$A�{Tf�z�`?P�v��ۭ]�!�DX!�@�f��>�N|��@W5-�!�DNB�@(�Q�f/Za�a�W�h�!�D��C\�a��uK�öO��!�$@�=L���e�(
�.�p�c�!�I���X��"K��A!q�G!$�!���r�k�W���M��䏴d!����La�*
�;3*T�K"�B�ɳ�Bl���A���}�&-E]��B�	�'�z��e��W;�q`�GؚC��B�I5�*�9��9ۄ���U�C�	2=?n��S�],��.+9Q(B�+Z\����c��f�����t�^B�I2�T��LӴq_�9l�1�C�IJê��F}w�QQ����3�B�I-*vҒ'ʁf�i��aҕ;,8C�Ʉz�t��BgY3�nT�U�P��B�I�d��20h����(i7֎B�I�ȄupP@��+��R�M�:C�	
@72��B�_�=�Jx�RT���C�I�6%+��د:�\1�TiR�4HtC�I�2�����b�kZn��6�ryTC�	�1c��;�P��JC-@��rB��4u�DQ����B����Q_k@B�	4$-r7b�_��� _�N8FB�I�&D��v�Y6 }�W�
nO�B�{�6�h%�A�V�ؗ�݌"o�C䉋�ap�
(e#`5�pB�	�M�<ܹ� AHF�ڼc���B~���M�7'�D���^o�ń�k*N��ˀ=1a�%ʢ���J�v-��@�p̚v��J���ӎȂP~�ԇ�J��sşc(|�:F�${G �ȓ_h\	
��E1YnؔZ`�D)W����ȓm�2	 t͏�\h�� ghH>+�$���,�`��f�6�.�����8$���ȓzf�h�"H0~�z���3!�*��ȓ(v�%@�)�&x��Q��Q8`��Y�ȓym*IZq#��J�2�0S��1g�-��+�.���ŹhS�Hw��=�������B�A?rt�Q u�$x�̄ȓR�6�[ nT�69X8��^�Z��ȓ&h.Q��gp<ʹQ�ˠaFBm��I
HH�E@w�ʘypʌ?w�E��Q:�9SQ"p�Y�c�{����ȓx��y˂'Z �%���ؑkr�=�ȓ2n�cÐ" ���Cא]�:$��(H�(��_�zN(T�E.M�B����N��=qKK��~|�a��c �U��Yd���ʈ� yPA@�h�~ ��T��i�!h�(�����N����zx�W���d!h2!�q\���L�=� ��c�V�Q�A��)�*T��S�? A����~
�"�EP�7�L���"O ���-3�����+�	(�,Q��"O�ph;�q�J�|�N�Z�"O��ⲀB(*�*W��|�PK4"O��@�
Âb.0�#�!(|��
�"Oީrr���H"�G�Q�����"O���K�%@��!��l�?���t"O��BSh �^U���D�?H<
<K�"O�-kAJЕI�����k�a:$�@ "O.�r`��� ��tkD�,:5��"OF	+R��7aXy8����XK���u"O���#h!x�xai4iL�BL�X�"OV��,�@���Y�VK�"OZfR����)�mOH����"O�����(L��Ȧ��4p��(�"O�( ��͡8�jB/zu�aC"O�8b�c�;��� ���B*���"OJ�2���N]l��"d��:��"O<M�Sl=}#50���$r@�2!"OP�Yfm^	`8Y ç!��y[!"O\P�p��w�)˵f����YH�"O���QfX�g�]�5��?�2l�W"Of�1qbސ���P#��
h"�"OEZ��D��IP��p:���"Od k�
�1+��EF"�5t�Y0�"O�i��L4'cj�z��F;=�h �r"O*$��֞gJ�q/��&9�"O���/S!M+ݺq�Z+va��"Or!��掐i'R�R�!J�-��k�"O8p� N<!��bO�&:��s1"O>C1EY�O�B�JQ��86��Z�"O���ρ�BQ.yI��c'B��2"O�����]!�@8�dJ�i%��"�"O�m�� �4~��l�Q�. d���"OH�;P���(w8��d儷�xla"O�d��B�(��	N�"�^���"O��I ���&X��H�&���jP"O���fo�/5�&p Ǟ~l��y�"Oʙ#%3AL�6�φP]ܘC"Ǫ#3�Er��Q�"^af(��"O�4ˑd��7Č3��ܓ&Q �0"O� "�\7-Nd ����:S"O���ƫ^+����4i�ȱQQ"O���%!~��`-�/jj�0G"O���.��ytd�"��	$h�y�"O�=H�e��zu��7d�!�G"O��E�\m�	)( �q�ެzV"O5Ʉ`|[VaA����
x2�"O60)sϕ1:�m����.���"Oz���6<��G�=�&�0""O�9�%�K<W��×���q��"O`�� �4<�ވ��j��G�|+�"Ob�H�-��5�����Ԋ��"O(�j��J/�y���4B��h"Or��/��@m��1@�	{���`�"O�4�'IP>(�}���0�f�BG"O����Bĉ5��q3 K-2��!#"Of]��H��I5�4*���"O^P#�V(`��;B�5�q"OjX�턞tS�I�� +����5"OP<�Z�)�����9�2@q�"O��D �f|>ęS��� ��"O��dɖ[�k��V ?�<-�"O��	�2NUz�C�O�N��qr"O�  ��$e�'+�Љ���Q v�*Y�"O̤J1Ǆ6Z������#���3c"O��Ua|��AKGՔA��A�҈qUvP���T��M��4<Ox���ɛ��,�*�(L�t1r"OrTI��Ǝ�0�(FJ־1��-k6"O��)�,+@���3,����K#"O��-ɴ��]�!E�L�)�"O�)�4	In]��$�̮QyՀ$"OT4	��͢�:Y���o�����"O~�P��~;�Ty"�ߣN��"O����_� ��36oА3&��"O� �rk�l8
}:Q��,k%FH*�"O��xe
C�vT�7M�=L$�9��"O����6oU�	*��\r��{ "O�
i���ɷe�3C�$Ze"O�i�g�H�l�|ydR�=O:Qd"O�ѣd-Š!qz�[�`��D�Z�r"OE�Ҍ� �zTJ�DڒY����"O��c,�9�4!�4�_"h�Z�0�"O*x�ˇ%f�Y���z���"O<9P�T��U�T"�2q�<m!2"O��c1@G:l^*��`~"0ܺ"O `�4�� �����i�U^���"O�ei��6zFb]{��H���"Or���M_�`0�2d!B�"O���v�:G�
���o�s �)y3"O�2s�:s_~���/�S�Z}� "O�ᐂ��+������^�X��"O�-���ݻ �tY�,^�&�r���"OH����)v�.�ia��*İ�"O��'`3D�����g��!5"O����a .��բ%�ӞL�n]��"O8�iX�2����
�Y�@����y��)r0��O�>_����r/E��y�ҽ���FԫZ��ݪ�hG�yb��z ��(��S7R8T��R�B2�y�lZ�K6��ё�Fe4��1%#�yB��2>�6$�w�̭I�d���L�y2O�>9'���&�<�����?�y�c�5������&<c���O+�y�W%֞�S��6����G`	5�ybiۜu�\m"F+П-O!K�iR��y�ϰ+P2�ު ��������yb�R�u#(T3F��H�`��'����y2iV0*��cf 
9��M�F����yR�N�~��i��7V������yRM��rJ�����[�*=�mʶ�y�$�	b�8����U5Ty�[E�K'�y����`FP�ae��' � p1�ᇴ�y2ҸIХ�d�I	b٢�ȓ�2�yr�d�I12S-U�Xؚ����y�'RL�x�*�nQ�O_��9COD�y�LX�`�]���J�@���c��M!�yR��=*���"�"O)<%:4�X�y§R�l�0�7�ިZ3�a����y�2�2$;��N��T2#�ұ�y��
[��y)��;J<��R�\��y��bׄ6�J$Ou����	t�!�d�&S)||�Gl�
tzީ��V-K�!�d$dƞ�ݚ]i(+��0�!�d��q�D	S6P[������U;!�d�3R���K�$\j�k�O�9:!��q�d�a&��7<�@ȋ"J)!��11R$R��>t�\�2�¶ �!�� md��<\��p%��>xΚ�Cd"O�Ua�j��c$�,k�u��"Ol(�`�V Hxi`!�. kҨ��"O�U���ܻ�f5�&�2}^��`�"O����اuj$�dd��]G. �"O���`�P�.�Y`U)]�k��[�"O��b��3��%)�BBmSw"O�`�,JaM�y�V(ά`�L\��"O>�R�͞*Ą���$;m�"v"O�(0a�M7/����S�� _���3"O�8��B "n��y��BJ0O��3"O,��W�L���,�"߅�e1"OxY!�H�{'��1F�ٰ}l�4�V"Op\9@��R�U`��c_ژ�"OF����ӉC�Й�rRb��""O�)yr� кP-��IC4p�r"O>u���B�La�����D�S/u��"O@��&Ɋ�CB�����H�-*2"O.p�fM׆��h�L�!>��%a�"O��۷ɱk�$�K�x�d!��"Ox��A�V�w�\�yg듾N�z�C"O*����W:&�2m��i��R�h�"O��#�@ 8�Z�6)K���"O
i�ɜ��R�g�(yE&�"O�L#���[]2D'��m�+p"O~P�E�$p�0���Վ,p"%zW"O���#Ã	"r�z!�ǕP\r�1"O$�C��)&�M#ƅ�){#�$��"Ofq�4�C�]���֭�8�dP	�"O*BBٍQ�m�qC�3k@~�yG"O� )��ۆa�Q�e��
:Ѝ��"O�0���.�n����R�c�"O��Q��~�~�@�bX�4"O� IF&�n����զ[Q�)��"OĤ�p���� �� �
�"O��� �J�b_�a�Î��j8�4"OP��!�@	�e1@��)b��T�$"OĄY�N7Z|勳��11u��p"O�J5��}\��'�9<.�8�"O��B�eI�uآ�ԁ(��U"O�����4:#B9+2"ϗa	�(A"O���(VO�D̐����f�`�"O>)�4��*��pHwMدn�fɨ�"O�;P*)$G��qչD���v"O6#�nZ*��5���=�ָ1�"O�4j!g z���	ڐ<Ȕ`"�"O��8���tZ�i��� Z��d�"ObD�RKޕ;<��d��")��W�`�<Y��}+�}����U(�Pڤ�Z�<��凴<{�@͊�H"U�\|�<�c��?E@�p�"߾Do���#p�<Yq��c� ����B�xx����S�<	G^"�Ҥ�ϱ#�`!)Q VLh<a"胠/����"C1b�dL�q#���y����bC�M@cxو�"֦B{!�$��.��h��K�::e� QaG�t!�d3�80���W?p6�3��� )�!��EmYL�0��3X��s��O]�!���k�f�� ��.xGȽ�v��!d�!򄁂(��X���!C:��u.ʷ_&!��I�Փ�c]T��*6.ǳM�!�d�<x��eߛ5:zP�-X�FI!�$? �ΔZ���7q����M�c3!��Y�@"Rg�2�r!it��7A�!�� �DbTA_>-�2X�]2L@��"OB��J*�6x����i��b�'+n�CV�L�kV�1�7�A�w�a�'��a�����Py�C��]h����'��BK�\oNapc)S#�Ȑ��'���Q`iL�>�6<�BO�/�q0
�'�|uPK�=<YƵ�a��2d����	�'���k3�_/�QԬ��cwF���'�hۥ�Pc:؉���Dcn���'��|��O�� 2%h�L).���'�.���α`V�I�4�O=[��Y�'%��$�!I́�� (�����':�{�:B�@k%��:YЬ`�'���"����r@���ޡw�B���' ���_(�3��.����f'�<�y�$A	|P���M"�`}�
��ybf��lLQHB ��xdZ�/ޠ�y"�\GkP��3I\'f�h%ñ,ӵ�y�g^���ĺD ��MjJ}�`�y"B�7�K��Q�K|��`q�ڃ�y�h�9�9�F�l� ����#�yRIér��P���!T�Xi��_��y"Qy�^�÷�T	�(�����y���Q;�8��&A��AȞ�y"@�h�l�T+�7&����폭�yBj�e� 	� @KJ��L�c��y���X���bM�>uJ���y� J��af$�3���6��y2�С���3���7%�x����;�y�.�o��@��� E�I�W@O�y��QO� �PN�%n�37�4�yr�I�"�tA ���#�(+�I��y�k�i���[�j��~�����yb�T�p�$�2�nɣ����A_��y'� j�V��VM� ��8i�� ��yr�f�IR�޴�}��ȇ/D��sC�_� �P�".z��:�8D��X�Š\������?&&�x��6D�H9w�Wu~ԅ��ȧ~�HX"�0D��)�aӂO����n�.��@�F)D�`��Iȹ$DxU�Gd������)D�\{6X�r��Mhc^()�t��'D���R�ێ3W`��݅A�TA�A�1D�
P�]��0Ñg�-Tv�2 �;D�h{�MzgdD�v���.�vH0�"=D���'U$�EI@V[���c7D��y�
�!3Z�e*�fS�z�t��p/9D�������rk��I��o��X���7D���c��1>fyj���	5�v�q� 4D���F��$#ZE�����>�)�0D���2J ֡�We*k�|%@�8D���"��SȤ�a�MA�l�Cv�5D���J�?F�B��ݠL�n�1��2D�X���H^,01�"�'� ��V*0D�P`c���La+1&S�&��U�g�,D��3H��x��	��圞=�v�$�,D��	�Eȏ]�]���vRj.D�$�`��:�J�I[ K#\ч�)D�XS��O-���78YZ Q�O$D����Ƙ�N�Fy��ƆKl�3e$D��w���@1,!`$�H�b|H\�� D�l�"�/��tc�	HG�.���9D�,a��K6w/ʐb��ل/g�CW�2D�D`�j�@n|�G D��,�
�J1D�� �9���ڱ �"  �'�X��*�"O�M0�kP�'}��S���r���zE"O���F\,z���@�HQ'� a�0"O&`#Q��-#�t3!'Y-#��)f"O,X!Ԡ�-Z�&��P�Ƴ]����"O��������P�j��r4L<�w"OJ�8c,k��ҰI�~E(�9d�8D��Å�� +��]Xe ��^�
��,D����%�on�h��M>9z^`S�K*D��`�]��H{���8%��t`�&D�t#�`�m��u�`� Z$x ��"D��t��bӄ��-\r
	H1/?D�t{��B�5~6��R��	�:D��Qw�G��T+��V�[Ȱ�@v�7D�$J���Q|A�cA������f(D�PQs��:��m"�T�_�\D �*D�<��N�yφu�DҲ�6����2D�(��aG��$����yff	�5';D�d9��k�&����Z
�$a�*:D�d��f��z-�إ�W)/�PJ��$D�`����?�b�����9�v|�3"D���$	��Hʞ�ej��>j�ȓ��?D�L""� <��:�M�G������8D�0����f�ix�bJ���@�6D�8��QM�p�Q4�
���8�$?D�T��/��}Mڑ�bǝF�H	��9D�P��I]�wʹ��ǌ"a��$�<D�
�I	v��}�D#g'D�@�#e��scfÙ`�d����#D��Q�'�)<2ɯ���p����y��:#���Я�-L�#�l؃�y"A��6�(�KI�8h�~������yB�I�"���Z�KA`exX
sOƵ�yrK9N(
]�E�9`X�9�×!�y��#Tܘ��`˞�����;�y�)\�fe�+`=~J&A�#f#�yBH�![������2%ex�p#/���y2  �jL���kY���9�y�D�l�`�	�xK%"P
�yA�<�|LA׀�� ���čR��y��� ��$y6`���� ��y�a�Z4E0�8	Ŵ5#$�y�K��zp���5��xS$,���y�B_g�u2��6Ѭ��@J��y"
��Ori1�AN�xz�ٰ�	�y��L
���D���$��{����y2O 8��dkUL	�R��\�C�n C�ɕ�[��E�6���͵AB��2p��P���w�D���M�:}]�C�ɔ �zMq�b��f��5���B��B�w9�R��O�E�r���f�>e��C�	l�Z���,��c炈X"Hr�>C䉂O�])�A�|����-��B�	# k����Ì~�JDᵠ��3\�B�I4}I�-(gʚ);|G��)ΊB�	�@s�Ƀ� �5pvDie�b�>B�I�i9$$�Ej�-l!v����O/:7*B�	Q���9�^�\ti���>mmLB��=�����2H�H, qJ
 �2B�ɠ-���R�U�<_P	ڱ 
N��B�	D�rf�ʉ�6M�]>����"O�д�ɲHUs�P�os���"O��)`�Ƀqs�h�'�:U�`�"O���",��&j"x���ˬK.HA�"O� k�&٦=�D�RJY�@�\ڰ"Om�r�0�ؐG�R6\��"O�40�șQ|Lqd$�8F}FH!"O������.=ɤ��U���(|t#$"O�q�G`� Xh�su,�=A�*��f"OԼ�:]����JQ�]��P�E"O0h�a��S]��[��"O��S��
=ft8����}+��SE"O��ȥ	FO�U�G��g�Hp$"O �SMΦ#�t�a���2w"O-���G��L�a&]8��u�"OV��,=l$0��Y�b_4$Aq"O>|:�O�0�"	k'I�Aq80"O�)��DGD�iP,9-z���"O�m+�*��w_(cRhJR"O��1�`n.�s�䒩e���[�"OF�x�N�j�����K�2Ҧ;v"O�I�0~�9Z��]�b�B"O*p��2��!P�R(J�ȸRq"O~`���5-�z�tM�<c9�f"O BT.�� f���@C֐[�"O��)fg�:PP�z��9@rd��"ODXaB�IL8Cu�ۛ�rT�$"O���.ҍh~d�� �P�&�{"O�-�$�������f�I|P�b2"OFI�S���m��K�:d�Xb"O�=z���"J)��p�
�m����"O8I��W��]G�H J��KP"O��2r�\�dB����ԝ{<xh�"OP���߽Uq&a�g	:{,<���"O^��E�Ճu�E�pk��ZpZ��E"O�xI��I<8i�H��
�Vj@�t"O�i�0E�5؝h���=�)ap"O�R�ـz`� 3��C�ޝR�"O$t�`�C3$�0��c�(�0�k�"Or�Ðo�	R&�IB*�|�q"O��JG' ��T�u@A�r|`"�"O4��QO�;ǘtk��S���"O4�U���EM�8*���6��K�"O�rSJ΁2إ�eBT�Q�2"O2�b��9�
h�׆%�&�@�"OZ�#*@�p���ic��?а<	"OX����\�^2��u��E��"O�[U)��mb�G�i���0T"O K�(i!��sUF�@�t�"O���k2)�&�	��L#�"O�`X�lۑe�l)��&��Y�Pa""O��;����y�r4�U�29�� �g"O�)����Z$D�BlF��X��"O��0��َ$��˂+���2"O�0˓���p�q�J�"q�8���"O�Y�D�ǲ}�p�����Q"O��b�1���&�S��X8'"O`|�	L�/��,����G��`�#"O�`I�dG,
�P�zE�q�e	1"O�q��'U�6�#�C_f�� ��\x���F�ٚz�2�yp��v��H2F)D��#L��=���A� 6Ɂ2	(D�X��ˏ������W�&���O%D��k�8��Ss	�$�.����"D�$jD�*?(\�`S#��D=i �4D���J�~�����!R1t6�JRC D���j�./�)jԿ<[�n?D�tpF(��e������(\ju�3(<D�� HX!P2/�}�5)p��p@�"O�╍S�x��'H �����"O���o���<���҈v1�$��"O���]�I f��tU��"O��bPO�,$�~-�F�+/���a�"O��X!���^��g����Q�"O~Љ��ӒDD��&*�hU+�"O��b�B�@#T�F���+܊�D"O����V� 3�4��fH�H�,�X�"OD܋�e\Y-J\�RfO�z$#"O����n˪g�@��&��X	�"O�����S�J��!k�EPGW&� "Oz|��I��a'B	�^�;<c"O ����.嘹;�nϮ0:p�ɤ"Or,�&��'U��5�`#I�M*T|1"O|����Y>6h ��bd{�r1i�"O
�1�V�4�F�	šϴ/��-6"O�e(3n+	,�XK[�,]��"O��1�k�!9�X�ط	�]hd=�G"O*���b¿6���S��#�x���"O��cE�����hS,j�8y�"O�A䁚<'�U��,�o1��*d"OD�֮ʟ�*{���|�UX�"O>p�Q�:�#�@�3	��aڣ"Ox�薾G����@�X�$(�G"O�}R ��\�>�21 ��/�Fi�'"O2 �Q'F�P��.y�^Y�c"O�p
 �S�l���R��^+~��l�"O���TȐ�p]����r�ct"O�8{g�P��&����5D&��@"O$[�@+��@�#F=F+$<9g"O����_�oF4�f� �t�UH"O�Iq�(M�0�p��In
�f"O,�רC��(vO��c��u�!�D�?���kJ�"�k'$t�!�d�,pm�x�vR�F܀��0@�!�R8;j%j����c�J�b�`�5�!�б,�vł��F����"�E2:�!�D�(=�|y���J8�S�_('�!��ξJ��zЈ�|�v�Y��)�!���]"`�ia���#��`pT��8�!�$�M�E��!��+ޜ�R2^:!�ҀA���r�!J��n`+�f�!��W
|�0��w
��m��A#2���g!��1e�]�`NYA,�g��B�!��H@���S�. ň��[��!�$�C��	�aC� n�~�3D�W�T�!��2a\�l�v-�9�v�PE8�!��K
4�X�p䖖C��86m�~�!�M�4��T����Y5�[`΄�ȓ*�li��h�S��A�"��!=~ȓ~180��C(z��ĴI1๰	�'���e�I��8�0�j_.yՠ�i	�',�m�D�5�vx�Pi�(� �'8��F��`4[%l�&g�M�'Ќ@%͊�,�Ԩ�%��_z���'&�<r�Ĉ*�Н�2��%G��]i�'��)�#$uR�ph��V�E�FtP�'􁂀 
8@I�(�0@�8=�(!��'��m���T:I[��JXE� �)�'���U/-7�ĐeeY�:E����'���Ȗ険Y�8%�Q�^�0n�S�'�ܑ˔f��HrQ�l�)�Jp��'���ggJ�;�t*�.ΡLa��	��� �`QfN wE�a�Qo��R�c�"OƑ��/ �8��Q�'���"Ot+B꛵�r���oD8z�Xv"OB���%��$xP��N�a��"O�iyq鞇3��JP톶Q[~M1�"O>Y�M�es@!C��'P2$be"Op9cC�:��Y0-B�.Cp�ۄ"OFx(V�/�1y�R(F���)!"O�I���x�00��IG�*x��Ҷ"OHD�fWx��A�K�`�ְ�"O0+�&�q��!R#�Ţ|y��� ��OP��#�Mc�O�'t�������?�4>pB�r2��,�|���ě�vJ:t�FζoR��0�	,3-h���b/	�x�}Z�'�5�OR�\*qQ�کV�(�IP�5�M3��O�첁�&L]<}��%��9f��T��.�,����W�)��@r�F�nG��c#�LզQ�!��O��dVuy�����VcH8j潣�÷PV
uIT�Z��~r�'a}�ß0��b/�8\��q�t�N4w8 �7���A�ٴ��O���x�#DA]7���8��(9�'L��!�a�f��D�)�%*ϑ0>dN����X�_�<���B@��*��\X2K��?!���lB�!R2Cܞ�b�)��{7���i!NI���A���q��`�t��/S�R���>�b���b���T��J��@ ꋝ*'��шO��'\������O��Bؖ,�W��� m�(PO'`��!$�)��l�D��N	�}"��t��h���&5]���aӎ�O���|�>L�Ĥ��*טP)pF���a��˔1[Έ�
ϓ�?i�*��>�@�cɇ#f�*��X8V&r��J�|��I�f0@RLU���/�3t�h�҈��F��jPQ��W%,[|q�F��}k2bF
y�ɣ����'5~�B�%�֐����6�&��%Ј �L�!��9U���'�����	R�`����_�y8R�Y�?�䐀����y��l��ġу
���q�B�7fo�����D:5l���h�޴2$v�٧��6�$�<�]ELH��'�(&��M���́-������\;�c�C�ʞ�t�\A�� �3�X�KńA*U2��`3�^�]�	��%�&�7-��A���	��lP����ʂ�,�*̺V�cy���ok�㟌��M�O���m�Sۦ��E���Px�t�S�b�>a�1ND��?ɉ���'��ȹ'�ͥޮ �4�](F;�I#I<a��$�秊��4�M�$�<��2(�)<7|M�[?���EI�&�'8�)�I<au&̾��I�C԰3�0���/VfXP��O�*��20�iO0=*�́�ʸO���;J��LAD�� &-U��ɋ:�(mZ��bi��98B�x`"N�����n�&3L��'?�X�O�� �4��Y2�=$��7�ɒ"�B`��lZҟTD��4&6eۣ��/E�4�3iMh�P��?i+O^��Q	U0��2�Ntl���(_�5��PnZ��M3O>��'�u��;_��11�E4m����BZ�w�ʓ0&����i�ay�O4M^`+���)1����3�év70LI��H�<C^�Lē8Tk��\h���$��"HLH��:y�E�t �)�
YK��}�ʵjn�B��]?m{EHY�B�F��OA��R
r�Z������^����H�9��$�����[?˓�?��O>�&_�3�� 8DH�:2X2k�O��=E�t��F�n�X�兌9�d �䔏z�� o�!�MkI>�+���O�6��  �  �D�)�D��'RY	�@J�W�>�Y�&M�%yb1��'d�W�=b��*�>�p�)��4D�,���L�Kh��(s	�%J:�� 2D��#'*˲P�
���ψ�D`ԙk$M0D�pҵ�H�F�d�7��gsNu�C�+D��EkT�2�(:�-�(�$�-D�<�G%��1�{Ў�0dP��閎+D�0)C$�]ݴ1H��@�?��df�"D��	�),ra,=
�j�qܨ�n#D�Hا�O�t�hQ��%_(��i��� D� �斚"duzM�8��0{��-D�0����q�4�pe�)|�f��I!�Z?*$\����N�0�%��?#!���y�F��eL�x 0xJ3Ƒ��Py�c�{V4��3�ӻ�Ą��Z��y�@K����@�-X�e�(�6�ybD�as8�0� Ӧ)�l�X5�P��y2�G*:���b�])�PȚ�o
�y�E�)�T)Q�V",�H�����y�mA�`tr�JA6#3f�3����y�G��]xQ�Wò��K��y�i�'.p�)�`زR\��Ӣh�=�y
� �)Ag� 56��V��4#\Q"O��D$J/	|������W$�""O�%��8)<�DB��X�{�"O��a*�e�DD���Y�!�d"Ot3�$U!k\A�`�#�6U�"O�-����?&I��O��s�-C�"O2$��"�����c��DN\��W"O���b��|_����_� t�ȓgb�؂B��-OX�۶����<���0� >6z�A���&of8�ȓ(�j����ٞ�iJ�L􆰅ȓF.�81�A7&NL�y���#�^0�ȓFW\�3
� )�'įt�"8�ȓ(�[�f«s�Is�Ì?|6����FYh��_,�r{WKБ?�ȓF��`�Fe Sd2��ҫӥ��1�ȓ7LL�%�j@:V�]fu�!�ȓ)�4j��ɕP��!f�S�oE��Fo�(;�JD8�]IëG:RBe�ȓm�"�����5�ƕ��MQ�r����ȓ98��"L�+qV���.���^=��q�\i���N����V"�؅ȓp�-3���E�Ryu`�\�D�ȓ{��r��5-�a� �l��݇ȓV	�-#�V�WJ:��Ca�x/���"ޖ�����R�z�+4e
�x'px�ȓkZ����&Q/��'CQ�x�`!��iBuaS��U�&y;��"o%TԆ�=΄�(Z�3$+���5I�`��Gd��ؒ%��e���1r�j���fW�3�k�);��� y�������.H��IA��ʇ :�ȓN$r��# )P�^��w�Q}Nĝ�ȓs��Œ�B�*����L'vu�ȓe�t#����$	��gB�s�Z��ȓ�=j�CX F�}�w��e(`܄ȓ!�$��&�D�X?̩@�X5��E��27&��Mq��I�BP2uB8�ȓE�rL�W�S�r�B�J�6�"u�ȓv�$��D�
�Nz�N�<����h�%�\�h1u ��Z�L��ȓb����փXG��P-F�����>�X2�ʔ�����䔍� ��y��UZv-,l�ܴ u�� n�C�	?v`X��"
J�"@��G�sg�O� sT�̥��F;�d�Q�P���OP'lE�"O�4{6�'��Js�G�%����2egt%%����<!��8m�>��GI�?����T�<�@�L?�AJ@������ِ�p��c�%V���dݟLK�ᗅ}h�� Ώ�$�az�KB?>�h@���R?��K� m����M�<��a��n�<�K�Ex8�,|��d�7j����<�W�5l�����D+�'j�|� ��!o�����J(X�0T�ȓ*9���1��%ej��5�S����b�,&��'�:�я𙟘AUf�S0��BaY' d�1�)D��J�
͍B�, �+��c�b	�V�+���8��	�r��|�*��+G�0g��3����i��0=� %��x�t ��J3hS%��0
a��'ՒXAD>D�,�$�@_`<D�Qb(g�����?�I(f����I�#I�Q?}@���6\��1�G��Dt$xqf:D��b ���FS
��U�N�D�;�aث��bL>1��8�gy�/�1W�@�ғ�R�J���)����y"!	�����R�ިL~�I�$�-�M�`=XXH��ןx������E�4 �ʞ+r�!�� BpZ�a�7i�� 7f@��ֈY�"O,T:%���rmtLpP�[�$?�AJ�"O���0`O�D���Ä�,,�(4Y�"O�� ���tX��3��tĶ�k�"O�ty�
ǬW��pSa�r���T"Ov0�w�O/�bAQ$���x����"Od<p�X<���� ?fRH�t"O���[N�f��Q�U� N����"O���Zcu���Q�Z:?RP�Q"O"Ē&��MX�yf��jLx#P"O@�{7H��{�.T�0�GP&�-�"O�4*R-�z���g��
Dp	3"O&<��G.I���5Fo<���"O��Ql݌o�V\�AŖ�@��"O��,X��^��*� $̄�"O��"�9w; |QwjB�= �Qq"O����$ص6�v�q��F�mpt"O<����%bb��iG��	qF"O> Q�	JBѴ����C1\
�!rt"O�-(RLG�_ЦEa�CMQ�j�C�"O�!�f��	A���h&z�X 7"O�\�A���k���Hvr���k�<���%M�	�kI�Y��I�Wy�<	�M�3~�0c�=����v�<)�*�5q+Z!��B���@\H�<a�� :��s%�	n�P�[��RE�<9�W�m�B�z#�� %�t$Ii�<	V@��*�G�vo��K���d�<��e�1k��+�ǂ[�`�9�x?A��ؙ>�'�����Ӳ�5���'|���O�P%�i1����n�1�����w�l�AED,c���`s茝
��gdB�8J>4j��*6��̉P�ϱzC, ����O\�BS�,��>Q�Z�y�ؘ�ڸCp���G�
k��W��MY� �4B��	WH�4�O؎%8e`�/h�D�(���\�NM����Q ��V�T
`����IT�0<y�CE�<D S�T3Q� �ŅڝE.����4ZS��ԥ�.�Z��[ e��@�shA�5��x��aK�R$}�`��f4�aR���x�"�H>�f����@�f���?�����i���h0+Oi��DX@�J1�����p��O����ޠn48�j�i���E�ɭ��=�f�_��G�h^���5f"Yb �a1�
P �
���Yi�5���Y&��@@*sT�����,O8���σ�&w
1`"���Y3�$��=a�A2QGA�<
2n ��#lڴp'#�s�1�u�\�d�!�F�	q>�U�ag��^{��56O��
��b���q��4E�ջV�S��8����m��OJ�O1F)���I�~���j�x�4Hr�z9|�i�'ȵD2��7��A<i�C��c��@� ��4,���V�
�N$���K�3P¸�[� b��l۰���(3UlK�|zVe܋%�
L��D0��������a����SŜ
q]p�Gfi���ED��6,�����:rfd9�����YFF���/s_r�?�=K�l���14��u ԁ1H���?1����Yv� �M�bj<c?A�C��'�T��%3[R9��OZua���_�R8�u`��<At���8L"�P:*:�GʘFъ�ۃ��!p"��h��dV��[DW�!��e�� !��Q�Э�E.��tw����0]��A�;^���y''�A؞����C-0�����K�FI�f"�OU�gꂑ7���X�.ĈCg�����Ȩ�`׼/�!���z��Ğ?T&`9�K52�������?K��j��$ҧ�0�`RC=P@���R蔙itvфȓ	��q����#BA��@lڞ1'a����u�)���q��G#Tq����/MvKq  D�4 $%M5:�r� �#�y�4س㣟����$���'m���slI�4�&x��O.j ���@��!�_�2���`
U A)� �� �@˗1D�D��o��. B�pP�]3X
$��o/�A��l��+-%F#|�Rʗ�2��AS󈇷����A/S�<qB��عٴ�\�9~�qÓJ 'v�%��i��H���O?�$VV�őf�K�����l!��G�-�ΐQ�NJ�)�0w�:	���̫tX�| e���0=� p(#oT!نyx��>d�Εz��'��]z��<����臰e�f�ks�J�3�~�	�.Hc�<�ÂO7T����((zP% ���Z�'mڹ��b�6W���E�dj�
P��C#F�"��#G��-�yb��_"X��.^�&k��¦h��M����i2���K>E�ܴl�zh&Տq��p ]�<���ȓv��jB�$~vBE0�S�ZL�@�'���5� S؞@P � �z��򤝗K�A�e4D��ٰ��9�6 �o["f蚕��5D��1[e��C�G3?�@m��0D�X�-J'�>,+Vl�6�*%Z�*2D�$�� @��W��Fa1iԇ6ړZKj8� @Ю���CC��<rw��3g�ۜb�: �"O���"	ئ2� �sv ]=B�|A��	,��yc��:e�듟h���K�B���v G�����^*�!��3�uٱ��4�,5Bѥo�v�A?,>����F[$EN�9��J�f$�s��	:��\"�D�4�х�	�/�(iE���F~<1��l˭{���G��'u(���B�iz�Ԇ�T1@%� @[o:�Y�f�Hl��=Is�Q�<ވ����TlÉ�T���)�L�ٱ�.e�&�� N��yB��!u��q!Cͽ�DPP"Ɣ%2-2ǌܔ=��Ca�OfXa��Y�|q�F�7�zq!eF,uM����3D�@Y$�8M�h�7gſMA����l�D72i�#D$|N̻�d��<���	!�F �'��V�L�2�X_������2H��bv�c!�e!���s6p5I0H�i�D���F�V���h.��f���@�G�H`f��R�B<pׄ1�r�B=sߐ��f	�Sv<�$F6��;]��a�j�z�s���i�b�>��n�+�������P�e���1� ��H���UOR����X&je$��o�<�ċ&�gy�G�Q'��D�Byz�z ���yb� L�`����j��S�z���2��4����a�0Ÿ�HN�,�`y�KQ

4���(m�v���B˿pz��[i�X �	�}�䬱S�3��'���	���C`n	�t��� �L
7$^x�Y��)Hnx��	�&0(�S4�{�6�)�@��fPF�x�.��M��xҠ����Jݖz�2#~R�)I�(M�\��dM 1<v��Dx�'(>9��Eȝ.��}.u��AK�Ά(P
�|��F3|�εIcΞ5&�n�'�.�G�,O�)��\T#B�W	Ѣ.���Q�3O��y���w�9�J�"~�Bf�ekֽ�PȀ)/�B�g
ʦ�!�̍;��I2�49Ó�)a�M�6b�,}l>�R�><�V-�<Z��b�8�vmE<[��	�~��qy��5���[ �«9G����U�"0L_�y�PIj�Ň	"�):�h�1E�YI`J�d(<A�kP=Q�uaS�E:@.<�#1b�|�'�U�C�]7��^��@	�80�F�iRÊ*rF��f"Oz�� � ��hؗ��*B]�1�uZ� �C�EqO�>��$ƛ ����X{v��d3D�,��
'bT:���Xl�R�Y�3D���ë�S�61Y�g�+@�8�0D�� R�w\f���ۗ�D\{V�,D�4a O�31r����-b�^9�g9D�h�ӅK,o�R��^�Zx�B`8D�Dr4,�%60�_�3-7�*D�l:W�;;4��i��\�u������5D���$�Uv���.I>
��)1D�T"���*7��h�I�vؑ��.D������$#B
�p���;��¥� D��Y݃Kzn�@IјF��}#v-*D�P�f��4��A�w�O�l��1���6D�RX�SN`��`��2�#2D�dq�a���AR�I�2��H��0D�PЅ�E�:8pC�$=�i�( D��֧Z�1MdPɐ�5\�|P��d?D������ʽQ�ĕ_�FH;
;D���I^!w���b��QV�9 �;D�H�'�Ð6��q+Y�z� �"7D�$�犼l~iq�V�nr(��"'D�� �j��çLZ:�DjUm�\�d"OH���M�@DIEV��$��"O��"b�l�X#�h
�gk`�Ґ"Olh+F���;����C�Ms�@1�"O��(�
�[�ex�/K�ph���"OdI����	Yg���qH�c��዁"O�M�e�O;`�Vm���19�8S�"O�\ڃ�G� ��Q�f*�w/��i"O��TM�:=��"�	L�2j�cW"O^�҅���J3��đQ��P�1"Oj0c7�[l�X�0�Ȝ?{"�Ъp"Odq�ԧs�8x�&K�\	�H�u"O\S�/P�7m4LACE�*��]b"O�8���5k�(�
ㄝ!@���"O�y��N�W��$��T�uB���"O�����S�����nJ37
,M�'"O��`t+��uܴ#vmn�vh��"O���g# �x�4tѷG�%N�V�S�"O�Bǀ|G����GQ/XrVݸ�"O���	�F�����C�'tB=��"O �s	R/0p1�Vi��ykK�1:�>�z��A��n����w�)���+���e��]��R&^� ��8,��\�΂H�)ڧ��Md&ӫK6����38�po�Ag0�ҡ�|��i٥U��5s�D�$_�@���,$��YR��s≫YI<�����<�íW3�����fy�Z�%�4��ˍ��xםK�>��Qx�F�rW���NWjy�L�4�Y�+\�ݨ��7m�?+�1f.	m��y�G����c砕�FAN�rק���DW�͸N��J�*�6�>Y�r�q$ވC��)t� l[览��^w�t��tdĦ@�pٓ䃞Z�<�Cdj��IFDhT(׽I?���O��"}��O��x�)ݐ	��8��U�P?��T�G��	��/[/\����H���O*H��e\%�P�1�١I[H�2���l_�!X�Auy��0�ɇ<g�$�S	$��P��?�,�X��	��1�`�d>��a��ʦ��"!��0|�eE'H��Ր�M�S�ʩ*◢\W�u���ͦ��a��U�@�Zç��5++�#!��7�D�j%�b ��O�9�`�y�J�F��a���iGv����;Ъ�A�ޔ/RX;tD�+K�8�k���D�I�r�O�>�ӵ[p�e��7U�Ȩ�ψ�&rJY�G�X<|[��y�a2�4��<��-�ƁړEW~���@�N)��8�M\(=Xvq���'�����K*
2��j�[�HB���'�Ԥ����.��\�RnW�A����	�'ĔY� !�@�΀HR"�:2��S�'S�J2�ܴG� �,��"�|��'Yl$������m���Z�4V���'�r0�WDӬAxD�KB[�L��'���g��&��)��$�!�.�C�'�6a懙�(t( ьB�'@ܻ�'�"8`3�6��3�n�b���h�'��ؠ�k^*v�K'�,[L\���'�d��gW	Ԓ�8��Z�Op�� �'C������P�zЙť\�EP4A��'u�m��$�#NRjp"�N�A+�D�'�����\�i����ģ=�
 "�'z�K�X	��}��#�m(��h�'[XP��l�'m^���s���aX����'*��Go�Q�3�܇Z�|���'
��	c�!u�ԭh��E���'Q�P��Ё&(ֈ�a�Mcb���'��:6o�"$F5�#�Tw��DX	�'ix`A���Ё�3@�vܢ|��'<���o�2J��Tr#�،\<$��'�t�hQ-F�$#H$�b�[:���'�x찃G��X�8�'a��
��':f��E��1�$1&e�>�rt��'��|���Ιu��ɫ5I��#����'�p���Hn\8��٥,;\x��� ��o�B�؄ 7�l>�-V"O�QQ����h��e����I=�|�"O�틀L��q�P��1��1#D}��"Ov|�EG�>�di��
p' ��"O�,q��PV��,��hE�$��"O���I%{E* &! p	���f"O>-��jV�u�́Pf�˯�Di�"OJ�p#�m*��¦%p򞉚�"O�y�S��P�x�K��1�ʉ��"O.�B�� {�AC�F:�ءRc"O!aa�2�6U��lYe�R%bu"O�p%�9�p�Kí�5��|H�"O4�h��κU]d�;�l���b�#"O�MY��K�&��u�^���ܺ1"O2	gg�,Ю]J�K�c� Ur�"O��$��< ��A���t��	�'W^�ӰJ��q��5�&��q#���'�,�3�Ё_6^��拎�8e&ٹ	�'ް��M��vb,ͰE�E;)`ب!�'�ЕZ7��M�th��(
.m �'��I�2�ͭ�y�C52x�`�	�'�~��0?3�8��&��\�Aj�'=vt+��*O�L���ߌf*֤i�'*�t a,ظa�
Pp�oZM�Y!�'��!��K�h�~P�4���>�89�'�E�g
�VY�	c���#|eD���'�v��foE#"�D�����
9:D#�'�R� E̗�y�9IѠ��f٨
�'�,��s���c��У��|�[�'�F�k1�I1f�B���"յ��${	�'���(Bۃt���j�A��e�,���'�E�dm֖���Ç�enB�`�'�`���$�	_�iu���y���4:u�)	p���o����ʂ�y�D�D�� c���{����d���y�F/Q~ e;����k���/H�yB�E i���	��I\�^E[Dɖ�y�/�}T�t*���k���Z��y`�*&$�]�d�˧�R� r�͝�yr*	�)��hC-&a<�9�����y�ŋ�nvH���/����j�"Ƃ�y��E�I ��f�*~0�3�Y2�ybKT`S�᷍S�C$�m9��7�y�	G�pp� ��2sSt��dW*�y�,���x2��e�Π�WiĀ�y2��{H�#��0�6�����'h��sk��%��!���KΨe��'�\� ᎑=2}LARc�I�Eę��'��ӱ��+yx8T"͜E�^��	�'?�E)0�05�̸��\�:����'K��8k�Y�P�_�����'�� 3F �4E��"�[W@���'_
!i!�>f���>�����'��� �Y�&��`�nP�8���S�'��'H�q���~��,8	�'�>I���a�a �ۘ}(�l��'�����L�46!�!�	��@M����'�,�!`�'^��m�&זk{�`��'�d�0c�*����6��c��s�''� �@J�**&Y�$�M<a��Mi�'��0P*��W�(�	#��#����'��}bD䥬�-vY��NV�<����K�@�"�D 
�Z�x�(�|�<10��"m�h8R��X
?���#Z|�<� H}!��"_@�� ����� "O`|���
Dm!!\��<��
�'���`���;#b=P�mʴ	<��'�������1Trf\�"(3	˖�Q
�'7"�#�j���xYd�.rXP�y�'���[��*O���^�{$���'��|3��C$_��a�ėfdT��'Ɔ,0��EP���`G4Ű���'��I�6oMg>���+�>�e!�'k��P�V�I�zt��K�
���
�'`����)Bp�)Z��xH6"O�(���f�80`�(Y�~
�"OB�hF��A����X>H�Рw"O���N$����$n�:j�X�f"Oj��$d5NiN���-M4aox�(�"O�V��~Ta��, �d��&"O����)�p��4�*v}�9"O��D��U���	$MK�_c~�+�"Od<��l��ܲ�I϶t#,�"O*��B�BU������R	�8�"O蔂��Q��h�SE��9��r@"OnM��ۖx/*XK�d��~W�0�"Oġ;7g��'�pD�tM��X I5"Ot裄'*��K��ϯ;L�S"O��1����̋���K�(`��"On��pD�H�������!?�����"O�a�"�S�D��O�A�D"O�h���(Z�}���h��s"O&%�#� yP&���Ƿ,����v"OB	q��h��`:'����0�"O@�ʀ�_
_�� �AKȩ,t�a%"O@�B%eӽdԐ<�DI��Et
��B"O�9��<�Ȥ��&�:wτi/!��N�A�<�i�CT!RN�Y��-_�!��B&[,A�t��N["���[�s�!�D�;	 �rc��Dƙ!�A�!��ԋ[����i�=f�.uX4�V�7!��<zrc��J,"A�>�!򄒭s�����k�DhE&��	t!�I�ODj�*�9fތ`{�c7W[!�Ĝ:z5���q	��+��D��lޖtE!�DZ�E��,k��خ��$�A,E �Py�L�+����'�
�Gfv���@��yr�ޚ����/W�9Q��ӕ�y���L�N��D�f��F���y�/ݱ5�j ��b��,,m3e�^�y�+�k�����*
Ai��O'�yr�$��9)� �������)���yB���v:~�r@u�I��.��y2猢5Lz��(�;U��B��\�y�л,h����G�}Ir4��K��yb�El7ȅ�����kvb�s�n��yR��g���W�H?A�%�U� �y�F\�<���nҕ	��)�,���yB��.x;�4��nT�8����sS4�y���7WN�J�F@/2	�4h�)s�!�>d�t,�Q��k�� ���.?!�d�.Z��=��h;43P�IU�
=!��A�$L	���8CD���6'��	8!���pu�}��(��gB��S���N�!�$O�.�p�x���U��!�/_��!�$(J^\,C��0ۼ|���0qO!��5Ƥ�A#K%]�t�:ը�-!�d�.}ڵG��+%����%�9A!�� �4�3�B@��]�򃁝X�-J'"O�-S��=_Ж�A�̈́�k���o0D�p�G���P�wY�m�<��Wi;D�XIQGO�U���jg`�L
va�V-D��r�ᜌL0� A!��:3�d骑m,D�pb�b�T`�رQJK3u29�,D�H��	S�(�4���!��U�hɐq�*D�PcqI��(d���|�T��Q4D��z�ɐ/;	$�Yt��#qDx�X6F0D���&���1HsC
94*p2��/D��C���M@��zr���: � �+D�����iڔ��v)Њz4�q�&O,D�4H��P�2��rGDJ�x��)D����MK>6��	�g�;r�ڑ���2D��0mS�|�3����nܔ���/D�@��H�NU���.9�q��g;D���C��zP�V�Ԟ@�*l�;D�L��̂\UdىbaN. �5(Q#<D�4x�j�)���b�:z�ِ�l;D�$��؈H �d+�`�lՂ��cC:D�|#Ƃ[f���̛�B�U-;D�<(��G=bz�Q��'r�B�*�:D�����6 ���0�/�s��Ѱc,D�t#W���](\��dV�,��[�$>D�����S0:�,}�� �;��ԛ�0D���e,�9 Z&�XwEB�)�t�V�.D�#Gt>��P�]�l�a�/D��Xb���gu� �寜;"�(��."D�0�'��8g>��u@5P���I��>D���)N��#�)#����3�'D�p)@MQ%�RĨ��"j�$qTF#D�P�qEҴGj*��k��o��ś�J D����gI�v�:��5��+����A4D�x���--�:Qkf3a��@��1D�ȸS��*VÌu���»<s~����;D�\q���S��P��tv")0��8D�4��J7>u���	�be
ţ�8D�x���w�u@�mJ�9���7D�D�g�W!xUh����|��9�Ĝi�<��*(����L+	a&Ă���\�<Y�'�:έ`�ͤZ��tZ�#�X�<��L:��ň���$�Y���S�<����0(h�H�E�1��bU�<�K��.����OS�Fh��R�<���,E�XQ��ǈ�p���pI�f�<9�H	C��e��0�BJ�Id�<y�H÷v��	iƋ��I k�]�<��և&�Q`q�Q�*�:�hD��t�<Q��až���k��x`aڱ�Dl�<i�gZ�s�逡���m�4�!���h�<17�Q   �P   �	  �    �  �&  q.  �4  �:  NA  �G  �M  ,T  nZ  �`  �f  <m  �s  �y  ��   `� u�	����Zv)C�'ll\�0Kz+⟈mڄc� 特m`�DB�6%p� �f�q�䐻"�m�|Mi+��.�c`e�	��IuJ܅b�"I�;0�4���'Y8��J��}��1c��)U����	��l%ʡ�bC� b�Ԛ�@�����B&� 9� ���X`�-��H���9���=vr�,��$�3b��4�WEXB�b5���1���G��z�*�4yir���?A��?A�⌽�g�X���`�r)X�������?��й0��F[�(�I)es2���O���؊\����6&���� T(�����O�ʓ����O���'	���O����tI���R�~��AY�8�O�牐�>�+�&�)������۴0�(��y��,���I<Y�D���ⓤ9>i�1ӑe��D������I���������q��?�P�wB���Q� �$/��5R��'~�6O��m��4כ��'=�6�	�y�޴`����'��3�
��K���{#��<���*�� �G�?}� �Ϊ'�0�W���LF�IX0�����@��m-m}[��i��6��1����u�?���lY�Ik^��5�<"�J�A��;:Ȕ7mP�K�V�i@DN�Y6��PA�,�D�tk>E�mn��MG�i���Y���` �="�5�j����B �ŷ!��7���ec�4v� ˃G�)�j��!ǔ(���@�֏�V�K� AO��Y�*M
g@x��pB��\��	�´i#^7͎Цu��\�Q�qR�,� zR����G(3~M"��ڵ��p���_|�,�I=^5��u	�"s��31��
d<|���U��sA6y��N�i����9=�6][U����2��'���'	���O����K s�I��'xD@�P �-nY�T��N��]�R�:Q"O�mA"�\�VƁ!�Ə�7��eB�"O����96��3R��-��%��"O���#ȁ1�И�F)��D��S"O��Jq΁�.?�	�R�7/��,	A"Of���Aif��Aj���j!;F��fU��~Z���<�n-�4i��	��y�5��c�<!v�@�U��y���G�]t�Ѣ�v�<�f�3Y4��*ʢK�H�!ʞt�<I�͝�3Ft(��͠q|�02�I|�<g"A�������ic�c�t�<	�mS�f�(�n�>�h�AR�����3�S�O��lٱG�;C"�,�B�:.�ʧ"O���a�ލ+�D*4��:�F��q"O(�#�>�:��R�� ���6"O0|�D�K�%���*�M&��"O�峕�O?CMh4�LZO_��z"O�ep'��8j�XaP4+�.2T��X�<�r�.�O(�LN �0�"A�C�(��"O&	���Rvސ�AaJ�M��%�V"Op8��K�3s��
0��[�Lpu"O����MD�ufp��Å0����4"OB�a�m�d�x��з��G��<y��X�!��������J�x�2O
$��3#A�O�ʓ�?����t��$0�npʂM+s��!C ���2㟿e�X��B�6�t�)��I�F�J:c�M=���� :B�rL�%�z�:e"��C,!s�,�z/�� T�ɏ@�F���O�4oZϟ@K2�žM`�V;dI�Y�3GSy"�'��	S�OO�Ɣ;� �S0	�K.Y; #��1!�$e�����.\����G*s� `P�f�Ox�D
ߦMr���ß���sy���y�2O�T 􎐁CJ���Ba�>�XQ��R�ϳ>qO>�ف� �3ܑ�&�^�K��i)��;?1*Ƨn���"|R�O�F����N�9�H@�ľ����q�j�D�O�c>��N'bhR�Z�o�J<�r$4���O^�����j�
tV�na
3���a�џ�Q���L�WMJ,{Şb��c���$2K(S�O���	k�,@@Y�~ni�%�Ҩ";<B�)M�Х+0��\�>��"��:-�B�I,}c��zu"��c��|`V�P��C�I�=��d�h^�+J�]��I!�C�	��lE�$�"V���#���
��C�	����0�˟.I�Z�ASKT(��KeJ}�Ć�d����P��*O&6�8׍v�p7�?����	<kD��"�[;����W�c��C��=
kN=xw�=T$*�j2�Y;s%\��Ӣ�O�̇�I	|%P�8�@
02��M�r'];��Ǳ*5��h��'eI��a�h�vr�'�`6-1�D�=o�`�$?�a#A�B���z���o¤�Q���OV��?���?���>׆$�'�%^��s!��� ����ۖ4���艟rb��*s�4�G8�l9��O�^b50��1eڽ�Tgۢ �8��0��	f��1.����Ox���'�򚟘�� �Ca(�!��7	rte��A%�d�Oz����T���A֫M1�89��+]2�O�O��(�Ȏ}��S�B�_������'��	$O��2ڴ�?�����iI4��Dд2O4�
���(_�0RR?���D�O\��c��Sb�z����(�T>E�Ow�(�`�f��s�k��+�\�X�OaRT�Lw�-r�Î֨��tô�F�v�t����2 L����O��lک�H���)�7<��ѳah�"X�r#���XB�ɖ$1��X"h��("Mh��[=?�N�?1��ӆ!�B%'��q�Hd��E~��8lZ���'��D�a�X�$�O��$�<	�����	���RV*Y�������8.:���\5T�N�(���)BS�	8�䜁�*4:AF�2i%~��0j���	 |�� i]�!�1��ORP1-�4_N�a���U���C�'k�6��O 0�*�O c>��?9�%Q�+� �	� X&xC�j����d0�S�O)X�V��>o �b�d]?���I.O��m��M�I>�O��	=vp	��K�d:Jx ���}�z�*L��M����?9���|2�O�B�pE��f�% ��Hb�ٽM��]����Vm�ق��N�џ�\c	J3�$Ul����J��!�X��0�F�jm��s���iږ����%5s��Gy"'�u�+��
F�d�I���0����?�b�i��R�@�	Qy��?��TI���V9`��Y��*��6�OJ��"��7<�	1��	�(/���'�6��OUm�ҟ��|�	�LF�H�v����d�B<��Xj�J׏� I�ȓ�T]��n���GC�^���䊵� ��9��=;�F�"p�ȓt��gC+7��� �[�Qoj��ȓ~�^%��(�,(��S5PB���o��P*S)��Hf�
!�XR�F{�'D�̨��9��^ }Ŝ��A*��wR���"O�ܛ���O²`��7m4��c"Oȡ�r2-lI#�oÎ+���R "O>$���B��0q��Z�`�� :"O�T�0`�Q?�=�Fni�X��"O�Ճ�i3L����-�>��d���'a��8���7$� �#CҬJ�R�8&`F�n&���Exybe+I4%���u����o>~,�B�͇~onA����P�4��8�BL+e)�1 �UY`��� ��ȓ$^p@{�;w;΅`������ȓK�^�A�S(M)0p�ە9�n9�'^�X;�)%I�de��8�$�7g_�-��A6�Y�3H�	8T�zj�
 �Ą�`�	(���:+L�" �!�D��ȓb�ڶ@�p�-Ąe4:���c�R@#rG�.��сD�ԥd�Ņ�	5��	4��Ȁ�@�Rs�� �U?�B�	8"<R��3\_�1�6�Wt��B�I	P|��VI�C�8����U�TB�B�I&�<��%o���G���a�nB��0JJ�$8�"	(�[�O�2x �B�3%"�s�����ѵ&]ZȞ�=��}�O�:ܸ��j�&�Xs��=>&�B�'r���B��J_4E3���0�&;�'�
�����p���pKԺ ����'� ���ΰs{�e��l�;i~��'14�X�+��g��C@�-��c
�'��)y�$�m�(�C�R㖝��X�||Fx���I/\��,�Aj��5�u�U�8�C�I�\�Xb��ω(�^5Ps�S�J[�C�	Pl�I�튦a�Hkmѯ}�&B�	4>�`�1v`چ/��D�P�mPdC�IjwvM۴�ʈ�&Q����&C�j�*��5N57g�{"LY n6˓R+"a�����(c�*K�*�"��C�)� ��ZĮ	�&4S�n�*4���@"O�9Z���24ҵ@$��*+�P�0"O"0kA�&?74�Kc��.t��"OP�� a5^�[��H�]Ӗ����',hP�'j�d�s��%^L��u+��4��'�hr4EY<E� Eo�bO��3�'�H��I�l#�'�^A~���'�FpE��7�|��D!#?���'8�U�ax��U�cF?��T��'����C��am��2��Q�v>����d��Q?�h�����(���L��aZ�!.D���d!��U{��sd�L�fy��K�9D��y�����t�4��"6��1cS%6D���e@�#"�U*�HM�6�~���6D��B��!�heHV"�a�
YR��'D�a�L�_�& �flG;-1�D�P��Oz-��)�'!L(��_<F��)6`�',ҖDZ�'���DրE$�"�D��:�a�'��|�P���_��,He([�<�2�[=|%�DR�e*��k��TW�<���d�]��f��ea�T�<�T�Y"8�
U�e׶O�\5x���Ry��+�p>1 -C���ʆ�ʵ��)f]N�<��+���D�χj��i�2�DH�<��اs��12EoT!,q�3��G�<)�e�,t�j�m��aB���&X�<�5�A	/���:��8AU6��⪉Wx�H`E��8��_�6�Z#\?��;A�4D��	q��$��)'��FƆ��e3D��c%�8K�Ƚ�g��,�z�"1D���v��U����C
';Uh4�� 0D���D���1�l���Ʈt�*p�Ec D����.	-gNb��P�)��SEG*ړVK�@D�$/�F��4w
�}���G���y���;>��a#�W	n�s����yr� �Fd)�R�/Pت�j6 I0�y��P�v� 
���O��e����yB�Д6��p n4L��1["�P�y�� b��q4-E�/�xҪ���?��F�h�����Ո�π20 �o�@���"�g%D�`�ƥ�� ��r�mK�F��o$D���*Q�PR���$��MJ@�J3�"D�(
��##t0�kG*�B��>D�����Do6��7�@�?jr(�A<D� ��+ʸ	��7��d���<���C8��A��ݍC(� Z'�� aB�\"�(8D�$X �M\C��Q�̡U��SrG"D� ��K4�R\�sb��{ي0A%�!D��z���n����
l�p�>D��C�!��erz}���_�B���R��:�O$-� �O� RF%���>��0.�9;v
(�#"O������A���P��a�s�"OP��d�_8J��d"�E k��K�"O����!O�/Lxsu��t���`�"O|D��%R
)pDE�$�
lO��	`"O�A�� H�m���F֌6�ځ21�	�o��~��F�I�(M@�2_�LҒ��B�<Q������0���^��� ���v�<�p��>e@ܨ�B�� :�*]�ȓ|0�y+D��~���4H��n���>	�Z$�+{�t�X���
|$�ȓ.`>�gb� � �R*Ɖ3�9�Ʌ٘#<E��N�1��lPj��r�$q�S�	�!�$\,E�ʱ�d&�����!T�
�!�� ��)��!<Bp⇭��-�>�y�"O.���cǚ2>e��͉�cw@��"O�hQ�G?+!���E�*`�S6"OVm+���6Ծ�3��"�yQ��  '�O�)��Mê2~<��E���M�"O�͑WG�d���u�I�a��9��"O����V�M8M�D�4/�@��"O�]13(�)$���AE	H,2���"O6�@a�"y�biI�N��Щ��'�.T�'~�<��U���{�e�-u�\�y�'f�mz5咽O�~D�fH�0��T��'3�m�S䖰W+��*�.!�&�s�'�t!�@%�z�ąkENCJ�
�';~� bɇ(+���ڙ����
�'Ǣ���gslr�˴'N�ڪ�+��DW�Q?�#�,ȋEg&�2�:yq k(D�|T��q���b����{	*D�$�F�(I�y*G ��:~�(b�+D�LZ���#�"t��E �)Lp)��H*D���dI�l�lE��\(W��8*�"+D� �ٝ{���4�A6�Y���Of F�)�'f^��q¢]>n�j��s�RU�����'c�mK��[���#�M�TD�x�'����'U�Y|E�@zkt8��'��3��Qp��07�P(h4u��'�.4�R��J��C+X%xdB���'�L,yk x�8-�d
e�l+O�C�'�h�����13�}��Aèl�#
�'⁓D�G�H.�� $nzǮ<�	�'�su�1Y����y���	�'@���T�O!P��52�]�v�\Hx�'�j�%���%��!�R�&eff})�������Aք�=���s��{���ȓc��A����3��`{Q��!���ȓ&c�Yk0 ��~B0��Wc��,@�ȓ[?��b	*Mو��c��SU@���cm���IB%��{`c�\T&q�ȓp��ㄭԃ^�@u{�"K?=��mD{B������8tI[�P�jy���^��"�rE"O�Xs7�[6&�i���'ͺxK"O�L��`��NÚ���P�j�"Oa�tm¾$��Ac��A{G���"O<��-�F�D̊�&ۜ��ɛf"O4P@#�$�UI��V���e���'�Dݻ���@CX���m_�� sA"/�B�ȓN0��+��J��8� M���Մ�$��r� F6T(t��,9
q��fۘ���ԈCm��HO�x�@�ȓsLLр�kW�$�Ƹ� W$?�n��ȓ�h��OY�U(�=Y�/�[��ї'�\S�I��	V�?f1ir�� ʡ��	#(�S�V)H=�1�d�^��܅ȓx�x(BC�CY Vjb��a�A��m���#��>E��4qvO٦El�Ɇ�I�:,��H@�Bu�-�s@]�k�����h:��*Yx�!CS!28}R�M �C�I Y;��H��͹K5��!E 9
�C��0l���g�.�n�PsF,	�vC䉞rD<1�j�2T�Ҵ!�&6B�ɡ	e�m�VIR=�:ܲp�K�C䉪y���於��P�ǐ�_)�H���0�z$���;
����rb�D�ȓ~�"h�"¿?�8( 'řg���ȓd���� !#y�4m�� L+�@���S�? ��R���M����FBWY����"O*\���A�p)��^��L�q"O,<�W-P�w_
m����t�2�$�'*������S5k����FR8����%(s�8�ȓxo@���_�3�H���i��B��Q�ȓY��:P�T	Et�[Wk�� ��ȓ<	�IS���<�����r�P��ȓ?�� �e��]��,�g M�!2N���9`iy�͜	�6�i�C�76h,�'�ڹ �g��E`c�!&��y�g����5�ȓ>��=����/5�TŘ���m�2��ȓr09� ����X�Ɗ�3�\ȅ�%�\5��D�-'�:!�l��ȓ]=�@P���xJF�[�N�?2���I�M��ɹ_ܦ9PV�j~�5�vHɖBwB��* ,SN�k~��e��/C#B䉦a�by�Ff�C�Iس��')��C�ɤ;�u���N=���s�� �C�	�z=ҙA�˗<Z|j��F,�6chC�ɩM����D%�16V)���9A���=a���S�O�`Ʉ)34���6�( ��'�H㗩ֳf@<�h4�
|�L�
�'n�5���T�'��l�@�^$yT�p�'TT�a̙6A�[Ã�;k+�� �'^rQ��h�lHZ ��a����	�'����HT����R��L�K�x���#v�Dx��	$5'4̹!��
*�`p�C�U8B�	r��A�
X&��]�+,,\
B��M���ޑj��=�Ph@>P��B�	
}�2	��{g����C
63ĪB�Ɂs�vL�g��,2��v�y�B�I�8��|B���2E�T�̒xc>��=1H���b�J?9H�x�w��06�CqN%%Z6<a��	Uy��'���'DN�ӣj�����o�9Ai�Qb󟮝K2H ?p���d(D!Z�t����!D=Ե��^-r��I׭\7cd��r�C�� �&mE�H�]&�����-T�2����I�f���O�b>I�����.^0D��΍�>5�xKSξ<��wu�aҏ�
aE�LCc�}�j���	����ѩe�H=���jP�5���W	9���!|�^E��ҟ���d����Z��'�j�R��C4���G!Q6����'E<j���P��R7�DO���T>��|b�N�md:]8�L� svJ��2���<Q� �D��d��߸�Z��I�>q\��A��h!1�X2 M�d;!R�'��)�	:?A!ˈ�!�z�D��:	Z�����H�<��FL�JI$�*Q�	 �e�P�B�'��"7K^�!��+PB_9���䥎��?)���?�3hÔ#?�r��?)���?�����d�%�����B��rp�_K��������Ò41�)�4�<Fx����Y/����< B����d����':z��8N��i͟��DK�%(d�����I�`��)5?Q!X������?ٜOp�Ԩ���,w��u�5	[:@=�U��'�f����2A�i�NO):^Ȝ��0A���Sٟh�'a��@�鈶2�2����A%*-@1&�9
�L�(��'�b�'s��h�������'q��Pa��;\��rM�^]���B��%)P4�ǅ��X�F�'�h� ����=y#��q\z�@�y��V쟁�� cs�*,O��+�'oy��/� � E����]��@�P�'����3ڧO=
���	�;��ZD&͚K��	�'��X����x²uZ� �!HD�I,O��)�Ir�:�~䥟�p7H�	j���s'��L_>��@"O��`�$&��Ex��T�bkz�Iu"O�SPo��8�<0��F�=}6nYX�"OTX�dI�:g����8º���"Ov�҂L����+�dĪ�۳$"O�hr��/~T���.f��t���D�+q���O6z�:�ٯ[&]���V�E�\9b�''$H)����a`ˍ�6�b\�	�'�P$p c5\�J����6qd=`	��� ��5Ђb��Qx��PY�EV"OЬ�ѭ�$}��5�2�.{�6�!4"O����)j�0u�!@A�28\P�@�΢�O��}�A�f��D�I�Jȶ�C���ZF��>��kB `�|5+@W�Z؂8��	��5�&���A<Х�gf΢44t��(��5�wL��MC���#�(u��ńȓR-��b�'@ a�;��>)�h��ȓXX�����V7q��EM�W��<�I2Q@���d
�E�R��/'T2P�lZ!��9v�䃵L� N������%�!���~���K�w�ʤ+_�!�$97vbPKa�� �8�	�m�!�K��q�����%2A��џ,hf���M��?�O�� *�[�@�$��ӏY�]��K��^�H�Q���?���\�B�˦	Ir�d���ITY�6=�2���L�O�Ș#W�ޗ3������7a]v�I�+� c�"L�1aU����!��127���4�b�LK%x��##��O�#|���Վq���CS�ӔAI��c�\�<�� ��M�EM�JZZx���.OZ��=XB8�9'CE
��D�#V���Οؖ'�O���.�P�0���rT�Y"�Q�Pׄ��:�|%��C�-Y�,yx#��[Rn��?�4�ēA�8b>A���Ԏ.�hdq�6z�y��(?��O��q#�>��y2DJ�@��{4E�41��Z��ֻ�65[㓟p�I���.}Rk/���ck�8hUƆ�n��t�!-^�C�ti�I��a�'��>�	KG0�C"�$dߔ$�ƀ̋aHx�dD>}�"}�`	��I�����pE�-3сv\��s��A'Ę���I2�N�*R���F���cb���6�N��놫�?Q�(@��v�$ɷr��V���.��B}ތ����)�$����)��$��c��sQ�?����?A^HQp�2Ad�x0��{��I�/�ҧ�9OhT���*�&�5H^�ʶ��`�T�⮃�to"T�'*�mJ�O��x��)�r��cR*D�;1��AIɸy��@C?��MN~ʟ�dSq��$@+V�9!ꈁ}�i��8N�2�_؟x�uD�<u2�)���A�R>��2D�.D��)ai��q]��h�
(��lm��4$��٪���O��4E���x��E V��k��^�Jh�&T��$�tG{��	{���g�H(�C�0P�d���"O�%�P#�\�d��SD����
E"O�#��JV�-�d�3{f-a�"O��k�#�/���"ʆ~eP���"On9�W�M����!/�5\v�4"O4A*I-+n��b���"O���៫(�h�3-:c���(�"O�L�d�9Ȁ�5+K�6"O\Б���<k�0���+ި���0s"O4�	�Y.Yt��kC��#R�0�"O^�JtM��`@ ��d͎�	�"OXh�i�>P98��ad�/\T��"O���Z�I������,{��D�dZe)«^���=�FN��<X�v!V�,��}�gꍋ	"y�QL�sͺ%"�֬k���8�C���<��*V	&��쀑=J�ٙ�K�O�J����۶_�&\
�� E���1�0I�|1���îF<�Y��J�P˷l�(�$���t�6h ��j�>i�dqQ�%�=[O�m�tc�7x��B�	X�lL{�	�<��@�K�G�hB䉍:G�H #�Fֈ���l�2�C�ɼV�
�%����9�L�Xp�C�	/M�0�AB�F�݈U:�+$-�B�;R�L���-����"��+vB�	� 	���h�1B�����x��C��qc�� �B�m'P�J��^,;ΚC�ɫTl�IQ#b�.f_��#���bC�����yPe�~ �0+g(X$�ZC�Iu���h�P7(����ɿt�B�	.7Ťd�!�ǖ������E�I?�B�I�x�Ɲ��"#A���ڱe�8{!B�)� xys�w@�����
��#"O\�z��?i��	vLQ�|�~���"O���'ď$���K�7A�:��`"O���`J%z��S��;]|�x"Ob��Q�K�y��H���7�<��""O���`bB/Q2�)BW��7�H�2"O�P�*�T|���ӮH��Ss"Oh��q�W��p�u��bD 2�"O�y�ai�4��"	�7C�}Z"O ���˒+-�ry*RF�#8��%"O8M��y��\ �ZEs"O����;O̘a�K�$5�U�"O�vH �����	��q�� S	!�F�"�Tepօ�!�&�yQ!�q�!�D�6@^)a2�ܻh�"�)��NL�!�d�F��ѱ�I�)�N�P W h�!��/�la� [�XЬE���0q�!��
t���&�lDR�b�2�!�$V�(G�pC疿u-�}�5O�}�!�d�h�ˤh� L�x8�߄�!�d�!UfV��C�^�&���)����!���*l¤��2|���h[�8�!�V�S��(7!ގES�@��gOi!�ݽr��)$�XC��ArM̞Z�!�d7D%P&�E� ���P��ս-�!�d�Jl���K�C�,��3Gو�!�<q�,أ�~�<P�fV9Uk!�D\#Z��hfA� +����μ^g!�߾J	X�AчH|�� @*[��!�$[�z���E��dj��xц�t�!�ΪU�\��&!��ze�4�ckB?�!��	T"��p�䕑:�v�jBj���!�d��d5��hM�'�q8�+^*�!�	�}�d�0���N����7��}�!�d�@2@���ڷ���D��&�!��\��H��
�J�f��	�%�!��=~F<<q�ʕjmde�I�6�!��&2���h��7&V/'q���"O�!-%�Дӵđ�c>Q�
�'��ժU�է_�� �fU7����'T�8Pe��`2�tI �)b�p��'����G�3J��Y���R��<��'�4���#�	GT!@�(��X��'���H� \9Q��ǡ��mR���'���`�Q �B�ҡ,�h2(tc�'��<�$�X3Fm�l �È0�R5��'���(F��r�NN�QV�@�	�'G�At̏/o�0���-xC��H�'(���`啪*U��PR��*#��A	�'$dɱN�"T�4PP��H-j- ���'����/7��<j�ɂ�`H*x�'v�����Ύd$����)c���'��]H�BP�@>���й`8樒
�'Y�HX���C����)X�h��'�L�����T�A��}:�I��'�)Z�	_���Q[�ɍ�|��|+�'^d��'�1_FE��Oc,d��
�'��1��Ї�x�S挐'!�
�'�$�CBDR G�PE�0h�
�d$z�'�ƥ���]���E�;m�~ػ	�'X�ܓ�k�:i'���`���;N�1��';�J5'D;k���p��.��h��'�^��Rh�3#��ʑ��,��
�'o��'ˣd��P�Q^4<�s	��� ���K�Gft|2�K���"O���a�����bg¢ ؈�"Or`9W"�5�z����>��r'"OB ��Ԑh3̨*2���T�)"O�I9f$��
��qri�+��`"O�!�(S3
�r�����T�8�Ys"O<���g��X�0�`�*�*OXH��`�\��:�g6@��P
�'Vr�fk�/=e��ҕ�?�z
�'��Xq2$V�zش2rD�=�<̺�'.p����9}���4L��.��9!�'�=@fI��yAoܘ&�ތs�'����B%��0�=4�|<��'��D��� 2�u�� (�fE��'�XU��b	����Y��B�ꈡ��'B@d�G��;JF���ĉ�j���'��Y�Fl@-��QP � ~��<��'��<�u���4@�)ҥg�h�h�'�,�sB�U0��$��g;�A�'�ju��B��BPY3ˀJ�.���'�����H;?	H5��BH�>7(h��'��u+�J�K�=F[(:��y�'0�$�LZ�`ܚ,X�X;
�'r6��L�L ��)!�S0[.�q�ʓy�xą��,���B�!������3��I�<�X���f��&i�ȓ] d@��������j�*C�ćȓ	*^�b��F�;
 ����ц�� ��I�T�%�d��MÚ����LU��հ0@�|�0��5j����N��H� �4܀l���'^�6y�ȓh����,į;^V�����\��fe�����I���G�	�3Q]�ȓ0(f��q�9,���:�냭D�"	���}c	A�E*����lH�l� ���pXe����~U�Iz`#��>�ȓH�F�`ҿ���I��׭q��ԅ����j��ѝn� S�.N#�Z�ȓM* �ЫVÜ�&Ό������gm�4���`ü%F�݄f���ȓC��ʀi�"ڠ��	Z=	�e��tڤ1��c�N��)sΚ>&��	�ȓ^m��h�0t�����>~����|�h������Y���̷GNP���:8�h�\�p�6���5r��ȓwĠx��kN�S�9�B�'x�"Q��D�Q�#�*ihuu�[�JH�ȓn���yB�VF���DL�v0��ȓ@��L��:/*���� ��E�� H%�b��4r�H�Q�1#q��ȓN�X�s�>�0a)&�FLj]��Z-�xi�\�Q�v�*Ba_�L����ȓy����>X^�j�疳>� ��*��r)�.�Yt��M�x��v��(��dݏ9:=@�=h/�a����`�uꉘo�0ĠF���q�ȓ.6Vv�7]6p��t&�A'�܄�K�B}�"L*%��SEHN�E^�Ʉ�M�\m@��2�h�&��S8΄��}m�!���"��L��G�7̴��#
���!+}��m;g�^2��ȓ?Y =÷ ��#�
\�ၙT�Z!��y�dيG��/]����_�R5x �ȓdF�ծ��r͘#kQ[�j���S�? �P�,��JEN����(\Ș0f"O2�:c�IYB(�e�q��٫Q"O�A�f�?	�B�Y�bNd�"�;P"O.X+�d�(�vDrrˈ?+��U��"O�z���<~͂ܨ� �>����"O��B��B��\�4NZ�~�V�qd"Oݚcn�X��5	b�>޾�2f"O��L�"/Ў�r�j�2����"O��``F48��BQ�W�^,�6"O ��&�ր+ D%�"���x��mP"O�y��F?q�\Հ	]�()"O��&�^ 8��m#'ϑ�Z��"O��k3+؅n�*u�EG.2��1�"O�(�k���O��1�zR�"O ����΋h�<K��m�Aq�"Oz)���)T��I+��=p<l��"O�9 ˀ+���b`i�%��"O�=IG��H�������W.Yr�"O
iQ��ÈyD�suA�RQZ�e"Of��Q-��a�(�Z�/�?k��$��"O���
�;��a�`Q�=�����"Ob�d,� b�tq�J�G|xU��"Obq���юd�$Dqīyu���"O�	�'Bۡ*�4ܻ/
 r�̊�"O��R�߷$�����o��qzن"OT��"^'HlH���Ƭm��ca"OV$� �"H`���"�_�f:�"u"O�9�6�.B�Z �eKGd-�"Oh�2����T����<;E�Xq"O�+��զ\�Υ��H�o�L��"O<�AVGq0�5���W�|b5��"OH<���#�X+dgYx8P��"O6 ��J��n�&`��[?��#�"O���o_��Q���{/�)��"O�4z ��Z���ҧ�����AC�"O�� S�=� 䂲�D2�j��"O�1�"��O6�(�bϟr�N$�7"Om���0����_� p`�S"O� p�O
Fr���U(�1Z`�x�'"O�����"R��xg� ]"���"O�p�@N�X�*-�pe�~o�Ty�"O��Q`��^rr�i!D�0fz��7"O�U�1���l%��آ��eZH<��"ONdB��ҜnojU@�W7F�L��"O��ؤ�G咐� �zͩȎ�y�Ɔ�S\ �##N@;��`h�A �y�� B"Ver�ڶfۄAJ@"��yB �%F�h��PŖe��X�K��y���E�Pԙ���,� j��
��y�H�q �ؗ.X� 0q3#���yBNθ7��H�%��`��x�U��y��� N����͙4by|���%F(�yr�(K`�}�6ȃZj��H���yBh�0�M���5T�V�P�L�6�y�M
�dnБsC�M��U۱���y�>_�D��t�@��P�ƫݙ�y�g��>}8�!ɞ5<5|�21+V���'~��Ȁ������!h�,�K>)�!
�}:d-��B>��rmd�<� ��>M�I*A��K=_�,��'�~		F�Ր7tQ�c�
;\x� ��'���l�+N�<PZ���%g��'l���$�T�IP#�gѶ��
�'\YT&�$c�T���Pv��`
�'9�Q�/��r��4 �ȣ=�<�
��� &Dq�hףdz�2�!��+ژH@�"On	&�M�-h�u!�4��,�"Ovɣ2M�1��;�g��m���B"Or��B�ڣP~��ކv�P��"O��"
�>�`�O	�vfҨ�"O � q_�3'�4��-�r��9Qw"Od�D�PF�d���앻
wLi�""O��m�m'�$�0# ^��x�"O�U��4E84�c cɐ- ��8�"O�1�1��C���Z!�ݜ@�\�q"O��ǬśX�V����9u���v"O���P�T�] \����6�:��"OP�q"+�-lf���g6��4��"O��Xd�3[�Ȝqvb�p�q�"Oм�oR�X��I���*|hx�"O~A�*�@��D�.�."��""O�u�mί����UǍ	"��c"O���2�D�K��yӰ��].D�g"OԨa6ȁ�K8����c�B�4"O*в+\�C%xqs�dǸ�""O>T�Ҍ	)ܼ���]�N_j���"O
�#���n$�9���1��X0"O����V�Wh6D�@�T�#"O�����E�`l��C�� �/!�	V�Q���7��1#�!��XC!��0+�̰��`!��b����!��_&q�Fف���uk:I�g�Z;4G!�$͕=�$��ĄnV"\QԦ�$e�!򄝺3�FDy�m�"HK*,i �V�!�$� -��V�^�eWJI[$��#�!�DZ�fƎ��-� T� 4�W�޼/!��4l�MK�E�$�b!���I�@�!�d��eh�q�5~>(��E���!�^�)����D�2V>�P��M�%�!��a�����D�x���7�!���a��,L�!ihI�n�c!��ÏE�Pt`�HвL�h��j�#v)!��d��@5L�^[���`Wc�!�$ˉW8��p����nEt5���Y`�!�D�~�ԱQ,ڰp�m@7����!���	_� v�+wOH�q��Ѧ&�!�O>�Z8k���B�)zaKF�$�!��(ꅬ�(<P-)��Ȑ�' �%��>�𼛓`V�p��h��'�\1�@U�<^U���ѳY�l@��'i��R�?8�UA M�q��'ɠ�UǘYq��HVAͭ[t���'�p�xe.S�d��x����Rj�x	�'.V�H�(�(0�i�¯C�]��'K"�A��0Y��!�bD2u��%��'�� �V��!Jޒ��4�CAV��#�'l�C�O�"��T�a��-��4�
�'���1Td^T
��c�Q� ���	�'j� �w*Н c�N���%n�}�<���jdL���J��i�͋R�<�A ̀=��!#��[�`R1���m�<9p%Ԁ���������H�e�Zu�<9B�!����6��wi��&čO�<9�/�{#Pa �Q$�wJ�<�g�E1M�`���$U�ЉF�IG�<v-3��А �P��%:Q�VC�<�(��fuR9�wF�9zD�Q���M]�<����F@0�a�@�2Y �I�C��X�<�� ��v��"#�)-%̨�LF�<� @�Pq��7D� p7��Fv�1�"O���'h
^<{0� i�t��"O8�"�"	(k?�Y ���6$�!�"O���ϐ9~�� �ַ2�^��"O����Q4 �8��Ņϸ���0"O�x0G�̹}���%��Q� ��U"O���lQ&8�F��@���t��"O$$��IK�7�,���@�NY�"O�Y�V�[6~�Se�^����k�"O �Uh(������@,F�<-�u"OU3$j��W���Ĥ�=s1P"O2}ZƆѥfGָ��O#bh��A"O@Hz�+P�p��-[�͆5W�aju"O~��f�����	G"�f�@�b"O��[�#�!L،8��2r�`a`�"O�����Jt����HŁ��4"OΈ���Wv��[�
 &��Җ"OD�sJ��%���T���dX\K"Oj��%Z�9�V�Ď^B=("O��؇���(�;�MT�kG�h"O�� ޘ+V�����C�D� x	�"O �x��9U��`Ze	3�8X�"O$s3O"Р5�4k2'�H�"Ot�:୊�O�����i����(�"OL(�2۝]������W��()�"O�͓E`��?�fL�7cܑi���j�"O�����>���85�m�"O�H�
1{�N0y#�P�*��5"Ob�S��>hO���C�p<Q�"O���PÙ0f�m
�J
9�4r�"O��k�C�%&�����/�t�ñ"O�,cv-݆�H��'EMV��AIw"O�#�)�6�&��s)�==�;�"Ol�#n�&"�z�k�h0O�Z�*�"O���6��5�L0I2�I�.�XHV"O�	��B��Q�(��3-��|�u#�"Od�z)�t�5y5#�9�`���"O�p��*�,4#1�
1z�� Z�"Ort��V�&�*��/��t�"O20��׎57�x;t�¯ij�e��"O��Ĥ��mƲ��4�	g����"Ore���+%y@8#@��;\���"O�H�-@�F���oҠj���G"O����$[R���ΜR}����"O:D%��{XD �3�S�Vξ\J"O�P��O<1M��#��2G(�(i�"O�M��� H�V�z�eG7	^�X�"O0�S�'�y+���W�
nL�b"O.̋W(�7o �#�*�,EQ~���"O� �)�n�}��#� i�X�#�"O�arGM'�����,�h���)�"O����*�8�����8f�P"OP��T ��j����a(��2���2�"O�(���]��谛��E�8�t�c"OB5�P�Z"!�^i��'�]�x���"O���5��k��,�v	�g�.4��"O8 �KBM�(��"�S%I���5"O.����M�n1"	ۑ ��$Y0"O��@sM;��<���L:$��"O�Ԙ���]�@��Cd,��"O��ˢ��
%;D���G ���:�"O����Y-'����g�-j�DM�"O��y��[:�.u��޴j�"O|9�[�f�*�srJT�"�[�"O� �`c��A& }��������C"O\��3g�3e�\([��X7Vh��j&"O�K��Rx%45��acT hv"O6e��̛(
� ÈU��"O��j�Ë�\z�`'H�m��Y�e"O51�I�4N�%�l9M��1�""ODT2�#����Ӡ=j�(4�S*O9��ʇ+�T[�FpM2�'HI;���J�t�1eŔ4���'�0\�6B:6��T�!fa�B��?DjZ]+�'�*��=	fJ�$y�`B䉾3���B�,�2anE��S�|��B�ɰ2p��W�
�M���QCаT��B��5>pj�⡯���d0G�"��B�ɺo�|2�G �@'6X�B�	�Ni���'V�.������A2ԚB��62�>� �R��P��#F.pPB�I�)I�\2�-�0�4����=J�\C�	/E<m�-�]]J�P��?k�B�I���}23��P��y���ʒ&pC�ɑD�VaM�Ll�������P� B�	�_�p1��F8�x�apmQ�z�BC�I�C��@��
�0h,nAGL�&C�I	CNMX�@�\|�p戕j�C�	�[��	IEBޯ6� ,@
W _:�B�	0k�
�gl�#!O�MT
�~��B�ɧmd��cH�?f��i��װ}֜C�	�<(8��앎c��쩓���RB�:h:+�='QV$��ՋQ{��P�'k,�c�H"`	F���O�4�̼y�'��	4$�:��H������ޒ�y�`͡[���Q�	{hp�X�B��y��A=v����ٹteĨ�uI��yB��M|�05�]Ѧ������y�M�Rw��� ��%��[�GP��ȓ-@���B(�l�8�0��g�rh��V��Թ �p�)��ȉ]ӌ��ȓd�D���\:�B�3fo�)�ȓl�v�HcIW�WvQ	U [�qr��P}dU�'��4X�zy2�I*����'�,�k��
lt%��_v�����!�h���PU���ŇU�VM��,P,Ms�W&�&������i��.���gg�duI�Ro�t� ��ȓt�KǢ�4"J:(�0��e���ȓ]]v���h��t��@�t�n���D�4L���0��Y�2��D��W�r(1��?��9�j�\Q�Ą� �@�[T(��)̰�B͝�b�fY��nB�����-U�@��OC5$H���Bې$�c(Ӗd�����
3K`m��'�"TP��^l���Z�-	l3�m��v'�#�n �VM��N�1K�,�ȓw�i3��ME�.�2�K
u?J�ȓl�.���@R�C�d�8�K�K�
Q�ȓ??H�)2��t�*��bD���,��ȓq�@B&D9��p(�L��6<Շȓ-? �{V� ^�Ni��'//�F%�����`��S�ipv�!�ì��%��ih`<Z�N�6`�r�G�V4|l����X���������FC;&��5�=�#�w���%��5X�$���f�	�-�,	����FȰ&��5qC�I�}d$T���H�.Z\|��76�$C�I'X�֔�l5#(�E�!Y�C�)� �ZQ�<��a�v��%*p!�"O8T"B��q�� :�.A�~!Vp�"O^���ɖ[>�+��R�;9(LrQ"O��S�̓�T1��t,
_+xd��"Ot���	� ܢ�%;.6��"O�0x`��"��A!a��M��52E"Oƽ"�ߴ#���a��)�����"O.Ԫ��ݵK�p9Vb�z�]�W"OfqX&ʣP�bL����WbA��"O�D�w*�%P:���O�Z,Q�"O@��� )O�mH��pF�S�"O�M�AdX��I3�P�H_���6"O0D1Ɠ�}J���g�>hOV���"O����14�XY�2�T�*6|���"O`��ꁻ{D��X Y�:#��H�"O&�I�uԬD12h�<�)A1"O��B\?,����W�I2"OEر"�12�j!��>#��V"Oq�L˹@Z�뵯��:L<A�"O:Ta�G��39j|�c B���ʈd*!�D�q|�+�$���J�.�+�!�?N~a��V��%�����!�d��5y��1AI�(M2ɓ�|~!�d�4��䧓�$��AzW�*�!�d����aXtc�x�hp��CP1!�$L�&�����^29^9ӧ�լ>1!���	-��H㮔y.���wh�%!���
d�(D0�/S)� Y��8R�!�Ѷ>�}z1��
Y�( V�)r�!�,�.�je'J�f�¼��DVV�!�DO&^h��s�O�jP�h31m^6xZ!��1L@��N�I<�x���C�x!�Ď'za�#�N�#CXP��!J!m!��/�J=�Gb��N���#��Ο]l!���|,����;�D�82jɐ@l!�d,�ݩ[!"� d�U7H�|���'wB��*�ޕ��A�8ʥ�'C(0�!��c���#��4��(��'�~X��zL���L#.rpy�'-xxr�2e��A(�o'\�F|�
�'�P@�#�̂q�JDi�)	d"O 1�ˑ�v�J��\��
��"O���nO���a2���s	�q�"O�����_֒eA�� g$*�Xb"Oܠ�
X�c������E~���`"O a1�ڋ0F8q�e]�>d©b"O�-��
�,9���%EU;G^�)G"O �cS�*P��e��M�%�T�"O��S��f;I[c��hm���"O�<�"�Z��U��FA�pÆ�r�"O�l˷+26:Yw+O�\\f5p�"O|u��^�gN\�9�꓉wʵ�%"O:�CD��#������$Ev���e"Ot�Caڀ2>�usq�1);����"O�)E@��JC����p��8�"O08J È��pPU���R�5T"O�M:IG�b?2�:a�]�f����"O�1s���W,��U�
-�H��3"O.LP��%XC�\y�IY� �M�"O6@�g%�Y�jܨ�����D��"OdyZDe� |����/�xI:,P�"O�$�����
���Α#���X�"Oz��@��î���2V�2 �&"O�	�#� Z6"ǋ��I~|�ѓ"O� N��>'�=`Ԭ�Yz��z�"O��b�mF I����TA>~u�@95"O�`�WCW���xtIĊ���"Ol+w�ˤA4}�Gԟ]�~���"O�ꖩ~i��#Bgkq8�0�"O�Y9���H�V���P�@`
P�U"O����J�_ � X�Ꞙ2T���c"O�8�(�NZج��,̽��pu"O���,)z�.�@��X9:� A��"O�ܨQ`њ+0x)�r�[�D��exA"Ot��`N�T69���2*�"Obp"�oH @�AiCmC�h���[�"Op�h��'YW.�k�k���Q"Oz\1cM��f�V��1@�?���7"O�����|�`4��!�8�"O���D僧#��mi�/B+ֺHҒ"O��9�(�q��M�/�6I+~M!�"Op�(B$٣����Aώ��z��"Ol q6��9<tMb%o�!r&��"O��1i��$X�I�YYh��"O�p	T�\�t���&ʴ\eV���"O�OGZ=�h	��4THP��"O�7 G�b��IKw�X#<hM� "O$A����#,@�xa璯^8<p(�"O0�4��9|d|E
�"M��35"O^��Q��x)Ԧ�	����"Oܱ�!�G����rfͨm�T��!"O�I9�'�2��R%�#.���p"O���6kL�R���p*he��"O�<KaD�S3��ꄠ��m���:�"O��C#�A�ne��ؖ�$�{�"O�T�!�7r�>��/۷j���"O���S�Z�&KBE�B`P�!"OJ���G�^lX��ڹ��a��"Oz�Ca�׷�DA��q�@�g"O��UDS=�ju�F�o�"�d"OԴ�W퇤6�N|Hҍ./����"Oz����Z;[F� �q�����"OΡ"f��$� �96���&|5"O�$�eA+Q�J��B��ٲ�"OҜ��EE�m@��mJ���)HB"OP��"!�5:��M�Uk��%���"On�&�%���s��3/`lEh�"Oh�
�Ry!��JY�zD�Y S"O��I!g��B�0�	G$���� "OT��o��$���iP��[#0���"O�ɋ��?+nNTʄ�
�	1f"O��0�0/X��z�E�{�Dkf"O3E�ۅ �4ӧ�Y�%�x���"O��0����R ����.�v"O�1�fӐ|���U��L8XJ�"Oz�	�U0i�e[�İ_ї"O�!؅���lM�pA�� 2}�B"Ol�Y�M4M��Pf�1]L!#Q"O.|��K*n��`[�6"�\��"OB]PO��R�n5#��,w���"O�(	��X��p���F��5�$���"O �:��V�l�9:wkJ.h�.�8c"Otu�q�Q60{Z��#�7vrH�""OL[eO�x�2������]h8m�u"Olh1�&]$��t��L�q\b���"On-� ���� �A�K�5f�I�"O̐*�-��dp:Q��?\�@��'?�DG7Dv]bUM�R���C���%R!�� ��f�B�^��rm�?TE��"2"O��Ԁ�	U��ƍ�*o9�I��"O��!c�F��dx�+Z�����"O� ���8� �t��j�R\�t"O���i8T4�aÏ�l֚��"O%8�&h�H�
T@4��4p�"Ov(@�kG� ��Mkq�>V����V"O���V�T�XD�B��˟a����"O�pKrJ��k���(D����y���;��"��T�B�L�� ��y�6Z�Eqs��=֮�B#f\'�y�-W��]����DlQR�U��y��X�j1>�[V��4.�Qq`:�y�C��Đ,R�#��{������y�P�Ix�(�"�R���B�yN5��ʓ�M�|ָ(	Sj�y��Q:R���u���s��A�b�L��y"ғ`��x���V�W�4d�&	Ƙ�yr �� �6�:i�"O�$��ˌ�ybn�Nv�� � �K���ZuC�?�yB��*`��=�vi� G��ɨq��yRi�6F%��
�ǅ�B��L����yR�ۀ)XL*�L�A��1Y�iѩ�y2 ��(���	T1Ì�q�N��yb�+��- �Iw��8��һ�y�C�[��ɳE�Hk/\,�v��y�l?nNĺw(*^�9�RD�-�y��)Ť\�'MGD�`���^4�y�bV�Vv\h�����D���k_1�yR.��[��,�B	D�\r�T��yrf�7`G�q��`;
x&HH��I��yB��$���i3���*��������yr+���ˆ*+^�s7�P��y� �[䡓t̗���m���B��y�膮�0���J�C<v�Ӑ�_��y��?>~��GA.5;>�@��y��T*�N�(�fЧ43,iY`���y��r�Uh�!�DL)e<�y�AI!s!\ jrE�|�L[Q��/�y���\Q̘`O��AH�� ̖�y��6O�h��⭅�Mp@-�"JR��yJ�(x%�ys�J6V/H��(ҕ�yҠ�=]��)�@*�;}ݨ���E֯�y��[�$+����x��h�϶�y��>�������6#p�q�W�T��yR�ƫ+c����^�{��#��G��y����z'4�� bK�U���qL�y"`�N��RA�J\h@�Q=�y�����(���^����_�y���_�L�w��"��"��y≔�3���Q��M8��	��y2�ќ>������5j�m��#�y�#��;D����W�=X��)�9�y�MS�1���,�/�a�n���y�J[�l�f�砏?)'�MY�`���y��G�� �$ا(rV�ӥ�׊�yb���&m�$ZA�\� �Iه���y��X�ع� U6!�c���y�L�� �˂�,�u�N��y���#�\����eGlX����:�y2A��Nꓨ�d:Z�Z��@��y2�[�}��%��*�0]����eڹ�y���<-��2fnZ�Ud>Ei�����y����p�ک+&�N�xTXQ �-'�y
� ���%��	B��
#.�q{1�7"O��#a 
F��bb�'6z�x[G"O��2�Ϣ%�`��a�h~H��"O�0s��M�b@+� %"}�<�"O�X@!.U>Du���f��b�b�"O.8q�E�h&@�$ωzY6�%"O�L#���\v\��� L�T��"O�I���Ѹ=�x�*��[e@Q�a"O X秇 hd�$�&���0`�}Â"O�H��D�5"~�IB������"O�ڢ,�ms聱2�L�u���3"O��s`n�N(V�j���-j\�w"O}X��moj��D�O�Kp�"O�@r���
'mĔ+P��v=H�� "O�Uxr����٥�D}D��*r"O�d���ŻB�NM(j�h�"OƘ� d�>c�bx[�T$���'"O��(U�
<WYHDx�M�  �8W"O�3J���8`�i�y.Pp"O��Icd�k��	Pf��(T�|飥"O~��핃K�p=�Q
�&,�B�t"OV �V�Þ}J��IP�N���U"O*���\ Y���#e��y��J�"O2�9���#Va�}�I1s��"O~�(1M�*U:0�5�$�
�E"O�2���"s�R�:�j��܉(�"O��A$](Fx�T��c�k�����"O���t�@
j��
dɇ1b�Yh�"O\!`��R/J���)�.�"m����"O��T��p��1m
 ����2"O��I��B�ᶽ�lC��Ecf"O�xC-Os�fêD�4�Qˆ"OR)Q�gM��HQ:��\z~Ř�"O<���+`<^�	2�G�A� �"O�yeH����٩D��v��j "O)hdB[2�J=P$����6�JV"O�A��[-*f�@��9.� Ʌ"OZ�D�;t��\[���$�B���"O�(YuaЦ;�p�ȏ�g�zMڤ"O@���շ]]:m�R烂Q����"O��sF�g��0KF]-�ͺw"O�,����T1'�	��"O�qJRaPoc`4��΄��D��"OL�8u��]���C�	�}��\P�"O4�#b�5Y�lp�Ē�Z�t��3"O*9� c[)>0�ãM	|���"O�Mq �:e��WMK,z_� ��"O�8���	�=2&�I\�
T"�"O�9���J�7�P��AkD-P3���"OƐ�e��'O�4Q�H�?G1 �g"Ol�g��!`T�1�C\�@�'"Ox��C�*.��s'R�1�8(�"O�{Ќ٦LpB�[� ʬ��T�u"O�A�QM��hP"�-X����"O�=3`/X�m�^X����"�A�"O ������aEG�1��E�"O�0�v��d?.̉sg
�=x�X�"O�[��
�"e�&�s�(�"O�iyG'0\J�]���A"Ox��C�&nS�K6�#up���"O�����j���s���b|�x�"O���D��-[�Hh�˚�pH���"O4乢H��O{0�T��F:��"Oz`�b�	6aYP��Ӯ8�Ep�"O� �����n�x��+^�x�`"O�}���ws�m�F��+g`XM�P"O��(w�������S!*R}J�"O֌z6��'3>��k�/�7F�$a7"O�M)EI�\�j`�vDF�Iނ���"OBL���t���x�<�f$� "O*�i689[�(�!q����p"O�Y�%o\쌲5���;��1{ "O
#��K����K�i�ܕ��"O�ڄ��3�q��f�?D#�90#"O�y��'i�$@a�c[�o�5��"O.M�Я 	Jj���p"�
�*D�w"Ov���ӛ'��$�� VQ���2"O�Z��[�R�l�Q�7s�i�R"O*�Y/��̝S�8��qD"O�]20O&9�DM�uc�-R��k�"O���B�E$�H����/?�1�b"O�Q��RIBH;"�B�5�ճ�"O���+��2a� ���Գ9��ܑ�"O<�;�����s�\��F��"O��)AHǕ1r`�8�M�'Px mB�"O��J#E�][թ�-�'m���%"O��ҁع >�����kN")��"O~���j�>\�㫄�<Ne�7"OLHZ�Cy��@��GkC.��Q"O����G)4t�a��B-`�"O4�@�Qau&�@g�^���ʢ"O�d�FnȲ!G`S��B���a�"O��"�g�hHF���B�.(p�"O2X���)S��pq��Ԇ|��D��"Ol�3q�k�d�.N#U��h��"Od@���3{z<�sa�I,<�Vl�%"O:���M�x����W+Ιi�p�yS"Op�;V�P=*�<T6K�#BK���"O��a#��:e�,b���+����q"O�E�� �Gz��ҵP+���U"OP5�+ֲw��3!ݣX��m�"O�aIA���f���(�E^�:tP"O�Ts��Q�"Dv�u�&+~��a"Od�i�bɺ��ҷ���Π:"O�8*aJ�:}ڈ��n74<���0"O�a�bɌ9o/M���kW�=2U"O`1 ��!A���S��$� ��"O�a5�̒9�*p��'P�m3�!�C"O���̛�vM)��_�x+���"OH���,2C.�{G;����b"OHd� Ȳ&������Z�у�"O��k@G"��i��� ����"O���$���� ��GI�\�rmZ�"O�!
��A�d���q��[�"O�Mst�;s�TP��D��,���"O��S%C^/24���^�z1��"O�dbU�P-���j0G��af"O���!�[?T��2�(C�T�x��"Oz����6_��"AF�N���C�"O�Hi�O�A�c��
PM�d�a"O�Yp�
����(��[L?��a�"O�d��ᔙ��5"�m��_�-��"O���c%5��Y6��*e(�	"OJ(@&��(����1�Ŵk����"OH(+�k��ʐ�	���}��qH�"O��s�a��J�)2K��@2��p'"O� f/	�9����J�	:.rm	2"O�� 7�C
oKHЈ�A����"O� ��2���"*�ȉtM�!g�@��w"O�dȂl��f��ӟ^���Ae"O�mX���.��Uk�e\�Ht�P�"Ozթ�i��"�$� 
�Ҥ`�"O���(��k�r�b�早[؜=Y�*O4��4�I-+j*�S�RD��*�'�E����E�EjӃ�+�<��'�*Ƭ����B�KrސT��'��ҕ�^,.����OҲdU��'~�]�s瞉9D���ٶTB=��'�n��팬l�����f�&�>���'f=��s�,�p�戄=!j���'�����W-0�e�"g�^ɎQ�'�rs��!�V���׌W(�1
�'jrm{��S'�*��Y�N�Y�'�52�L��X�p���*Y��}��'6�}3�mJ�V/�Y�U�O@���'��-@)��5�V����J�&���'��U�q��!�|=�CfMpT�+�'��Q�E�D4���MY�X�D��
�'N)��G��j�����S�~�Y
�'y�]:4(��N��)�6���Qφ�
�'�dʲ�Z9*�]J��9��	�'���E	�X�~��!��-+NH�'��wf�U���rCD�V�`]��'1`A�B"��n�<�{&�UeJ���'kTղ0i+�މ�����[�p�x�'7��3���u <X"g��!I��
�'����+��Ed�,��l�:��YJ�'�Zt��N*DP�[7�A�	nn��	�'�&ă�%�g��m�`��0ș�'�����@�a�f���~Ѥ��'����d�4�z�q��N�s��b�'����u�0	�|�@� h��`�'{ DZF	�N{x�7iF	����	�'���W�L�r&ӆ�5cDe��'z��1�l��qʰ��DH..����'��-�&o2C*�U����*��Hi�'Fh�m�
x�\hd�Ϫ���0�"O�X��&b�\ �ȑ=:�v�s"O���F+"���1jT�$V�:"O�ic�JQ�k�Z��q��;��L�"O6,�����<�f ��g͌K��`��'3yi�
�_L� 33 �,`��'�*�3��3w��y V'S�k���'V�;4�ۃIF{�*ưcD<�B�'�n���ٔ#0R�"PJ�'M�$�:�'`�8#!�Ո.�d��̯-z@��'��<2ЮA.���bD��*���h�'2�H��,+*@�{e���ԉ�' ���>nD���ɵAF�
�'c��+��K5��
%<���
�'/����K�ޑC�����1�'�pܻ�_�!Č�)AD�`v��
�'-��� ��7I�rDK�J���'����҂F%�0̚!=yʡK�'7���&n��Y0����Ϲ%tjD��'�ȤZ�`	�iY����p70 �'㞐@��,B���ޔv�D�#�'�D��f�=15��X��3S���'�(�1� =4���G%D:|@��'�*� S�D:B��)i\�.�`�'�h� �+dED��s��4S~���'�RI��CI�.�V��Ɖ����x��� ��0�M&�� �
�'��"O�<��EW�qq�qqc�G� ��Y9C"O�k�*H�I��+A�6�Ae"O	�r�ě*�,���3	� H�s"O��s H#��2���{�½H����,AS�LN��iũzl>��%�M"�dJ�GA#g�qO0����SL�A����8�F�s2�=~ȅB�O<�+�������bpO�.7�������̴9�]ڢ�x.��$h��g��p���P1&˼�)�(�+q\i���.-�H�r@J��b�`<�"a�<)����t����MS���)Ǻg,p��%}HcǤ!Ȱ�ʱ�'L�O£}���$ΆP�eE�pHƝHP�T����Ğ٦�(�4�Me���)8�q�LT;%����$#�w?�*W:g��f�'C�)�L<��/�"m7�]S�
C�iV��2��G.,�4�Sݴ]���	�i��f��e�Ţ��O�����b��w"����Ȟ�i�n lZ�z��,��'X�[¾ �2��;6xȜ`�d�,�>��%L�kl��j*�h`坘F8��:�ቯ �MC��?i����O,>7��?+x�2�ᖈ
Ұ�$�W#
����㟴$��G~R�U��ʨr���_: ��L��(O¨l����j�4�P�$�48�
q��]B��]�pr4�:�M#�|���x�g_	N��f�J_�d��NE�����4`�RĨb�Դ4��I.�OxQ�A��=x�X%R͌�\E4���"ۍ/t�}����|�%�],�ݐ��Y���*b�n6ܕ��4��j�<`�LE��(�!-:�`�DQ��g*�O��Oe�r�$W�p"�*ؐX�nA�2�")sjS����hO?�ĉ�wܒ��Eӓ"g�U�Á�(S�����4K��Ɣ|�O���W�x��	�sܬ@3'f�w�Q &H�L
���Fʊtx�T���lr.6��^�����/�3��5��'C�<�R�p�	�l�:$H�(]�o�"?i���
{ހ�ׁ]/ ��xE��𐪥 -��{AB�1Q#RO�h�伱/Q'#EXt9(O�����'_����5���ɵ���{0LH�H?�7-�Onʓ�?�(Oxb?u+ ��r���އxN$�ӥ:D�TK�4t��@�!N���zRa����ٴ9�6T���׻�M����ħA�5Z�j�MDD cGS;����=��X�����(ܲb�P�A1�O�ڱ�vKz>Ţ3a�4�0�;Q@ߦR���k4ғy¤E���R�b�M)�ɟ1Qr($��,V�;3>$6�5,��a
"��Uè��R����5�+4U�H�.��t�	ܟljٴ�?����yBj��:����N�e���f(_ҟ�?�|�K<�F����ఁހZ�pm�4��g8�	ݴ=C�6�i
xu
wĔ�I2��R���P�@j�'�R�ۢ�v���<�'�zL<���uz�u
V�M�Sg~�ڴ��;��)�!_�pZ�y'�3yd�x 2�Z�'���8����F�9= ���s�^�$6͑�f����I�A��b4fE� 3S��"��åU*����hi�E�3�d˂,@1u9���7�i'x����Z���<%?q��M�&�;E"yXW�L�i�
�-s�<�GU->$�MR��^�)��ӓ.�y?1I>�p�i�T#}*[w���� �ց`�a+D��>�~5���(��9lO��9`�  �   ;   Ĵ���	��ZP�viė:&���3��H��R�
O�ظ2�x�I[#�x3۴|f�v�J=|L��gJ�'��l� j'�6-�轢ٴ.q�$0��\�I�F�p�� I@��4��X����f$?�!�r#<) �d��&�R�~��� p�<
'��`�^�xQ��A�Μ��'?����6}6-L}�D��$�A����36�̣ln*�c�CN^y�C�ODcs�ʎ��9O4�y 
�/��cEI�6\��L���X����b�8��D�`�葰1����'H$�n��$iq��%F��P���q�'�dS�	�lu�'�����K �R�	�7
�j�h�'B,FxBDH�'I���vjƓ4�T����ܥ/I���O5Ku"<)pI�>C䆚�J�PMV�M���/�H��OT�R������'s<!��m:����)�*rY�8i۴;WH"<	s5�Fa�*�Ɏ(75Z� +|�;qh�Z�>��#<1� ?� �B����P�¦.x2�Kc��Yy2��~�'���?I��ؗ	h���'��MY|[Sj�?t"<�e8�2����н)����B�R�]v���s�C1O<� ��$����~B���p�� 7|��ukƐ���lT"#<�m5�k(:�R�^6V��-AfՈs��x��o��X�K���i��mGDq�����|y�@�3z���*��$�B�<a��"T��P�<�2k�3Uo�O�2��>R��#%
�f�>I�s\�l���I�-C��Qe�:2z���P�:Y�I�"7D���'K
   �a�N>�,OrE�h��y�ޅ"#ŗD���8c��O
���O��O�<A�iX|����'p��12���P(� z�p<p#�'�~6!�ɫ����Ol�D�O����C?[��}���#�D]���_�7�!?u�y�n��7���)y�J�1_`@2��j4�e�qK`�0�	�<�IܟH�	� �ґ��)i�1y�i٫b�� �/ֶ�?��?!$�i�ЈӞO!��r��O8!%FMy�jDbWHLD�ސr�J!�D�O^�4�b`��k{�|�N����-hm]@�Vz�<P	1)��I@��Ty�O���'o�k�$)Wbԁ��	"{A2M�G�A6T���'�8�MK&�۔�?���?-��P�B�@�
��@����8�ٳǟ�p	�O�$1�)҆,
	���i���[~�R��m�Ρ ���A_���*O�	���?�7"���H����    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   �	  �  '  �  
'  �.  B5  �;  �A  H  aN  �T  �Z  >a  �g  �m  t  Iz  �   `� u�	����Zv)C�'ll\�0Dz+⟈mDԤ�57���DB�������$)�9�R��<5G D�Eg�  !Xm�@�߶>���VƐ=-�I��~)�U2�'Wꊠ���(I��A��{�>��`��H�t)�#GJ��x�R�<2�¶^5���Q���������,���0c�Ш�aA�H���EbN�R]e�pJ�8Q���5 ���"J�9pX�q�4gn�<����?!���?a�K����_#>�xؐw)M;9
�����?�1�i�*7��<���hܘ�'�?��v���aD��[2�%��_c��X����?S��Ɉ*48!�	�fl�l�p��A7�̠$�.r�F� A(�,q(@����<� d��1q������℅�F�g}4O�㟬���R*-��'��8�Q�B�s%���Pl@hܼ����?9��?���?i��?�)�,�ݾ �j�[4?S0���%C�=m� �d��a �4(���i�����nZ��M���i��fg֌
f	�E��+ZŌ#=!v��s�O������9Ahd "%.��#0�,���[Q���EG�u��� �i��7��ԦY�Ӯ�RdK:*��X@f�z�Px�E�I�lQ\{r�t����P�[�.�s����h���I�Dk�7���޴�z욁�X�E΄��r�ZRːH�𢅮)���5C�����GyӸ�lڶ ��9s��%{Ӳ���D�<(tM�gힲE>�Lˣ.�:yע	=��i+pcϰ{�I�ߴ��/o�L�X�g���Y���� cvO���`�ϒ�d��CĪO3d�܈�iZ�dz��N�`xv�a���AR���'�O��aNIa�+r��R�
���g[��� �f
����شj����O�4�;Ć ���@+"��l$����ވF��i� D��'!�D�h��p1�`�V�#�25�!�O�W� U@�G�0�H�֯��!�$I%Yn\�PJ%M$v�&�O ,m!��JנxXҁZ�,��cl�:=!�$�0@V
�bağ^���yeL24ў r��/�NothP��'u�(y���%���"�X ��-���#�Z $~�ȓY\��CHĨ}�x1� �M�r����=�u�8l�]cco�b,��ȓo�$�D�;��\��?l��d��@���:�遌|w�!g��72��	b�#<E���שrm$<��%�"l�Lp��ږQ�!�$ۢh�n�iUÍG��\��NLA�!���#�QN+���5�F#�!�V�=��M"`�A�\ 8�,��!�d�3H"�B(�_�P�	�`R'�!�dBn&�C�Kg�PR�	C�)`�ɑ2˺��ĉ�s�(ib����0R�y�B	��js!��(&��x�Ņ4���x�悚 !�D� V�����=B�&�CE�	!�$ݘW����I�j��8C��܇/!��.q7��i0痍i���A�����yB��>d��6��O��N��B�y����j�c5��$�O�H���OL���OF�p0��O�˓�y��Z�uÑG͙t����A��0<�BnU��h�	6mz�		��M+���N���В�W���D)}�2�'x6��O���IB�L��xd6R$1X�%�<�4;��O�d�ɉ-��̣#�OhQj��ܓOcZ�QSD�2yx8�qd��*��|J��'�L�	<:�dRQ�I 1x�������!�����O�˓�Γ�y��7���6��(e�M������$�`g�
�{��	S/m�>�2��ڝA��q�q$�K�	%� =ʗ��S.P����%BU6 ���
 6`��K�� ��ٟ�%?a�|����O�����Ul�-� ��k�����	�q����ʣj1��ň^EF�?)���A(|��@пD�hEz@��>X�H�� ���3ʓW�����/�(*f�$�<0���/� �)y�bܲӈ� <��z�\j�̢~m�Y#sL�3�����yZ؋q��cr�$Ӓ�ŌBv����&0���Gݝ.�	��^:E�H�Ɠh,`�#q�&Xk�Qņ�.;-n��G���<��q���]Z�L�p�T>]EZ��D��z<��#p��)��wL$i�ā�}�ֽ���'p�@�"˲Lۀ�	b�"����B����� �ز�R����e˹v⁇ȓ���+0�ʉGR䢑\ ;�,�%�Y�4���� ����N�;Bt�
&�O�l�L��w�@��?�,O���O�����,�\���e�.�.�P��!D��� Y��&����(1���ټA'f<�}5�l�ab ����J��Fd\1pq��!XO(�"��N�/�3�BN ��On1�`�'��u�"}?8����m��2!*�D�O��(h�)���'u��1�D(z�����O�yH�f�aI�!��xq�T�'p��O.���4�?I����9H�b������Ԉ�7n�d`JF	��.g��'���r���t��ɣ�@Ը2���T>U�O�|,�@*�5�m��K@H�O�JWO�(�\�h�֖\w��}J4�U��!��F�R��h�F�e~�鍢�?���h� ���0��88�kR�N�>C�<-�iʷ ��g���,*Pq�����h��d�Ԧ�St��&���4�g#j����<�wS*P��'"�'��I�H&\ӣ��	MӼ Z�a�z�>�d���b=���P~���d
�K�d�O���O��s���0�@1I4@�
$c(,��_$7Vx+�L��1��܊rL�~�UFI���F��,$��p2��$�?�´i��Dp��Y���	�N��8����;*a�����.ٔ'�ў�Gx�)�>R'���U^��`J���$cӞ���Ozqn��(��ꟸ�O��%#�)�-9�6�kF�ܰ6#4�b�ሄ*�6�O*�d�Oʓ��Id>���_���1yÊ��&���'�;���"�Ͱu�Co�@�FrJe�5��+�.8iꁣ�"`#lR-�=r��ˇ����_�+W� ����(O�E�D�E�$�1U�~ĉ�B!j�b�'�6M�O�ʓ�?i,O��'[N�]#iL��Pe9�,G$R�%�l����}R@& 9����ނC��������M�����?YC���y�5F�F��׍ _���� B��y�kҙ���$��5mzy9׈ ��y	�T�P�Aci�!�4��Ù)�yb��~���2�
�;�L�����yR�\�k��ѴǏ��(Qk�I"�yr��(Et��� �={�(0����hO������&!�,PmV�\���Kp ]�8�C�I�
���cAL�v�j��v�گ&�C�I)ee��K��0@`~-Z�� o��B�ɣ>��рh#���7-E�B䉆CVZy�'덡m�,�`�ҵ:�B��;,v20��\9~U�aQ/us���ܬ�"~� �G��t�ڳ���:ǔ��d��yj��
��c�� 2 �c�� �y�b��c/���A� �}�i�A@ۥ�y2G	�&�����jM�
Q�U3��B�yr�ТiF����YkP��#D��0�yR�I�^���XP�_�c&*4������
�|R̀*��B	1Ea��flW��y�%Q���Q���&��0��bF�yb�_��b2���Q�.��e��ybKq�,x�5>�`ti��V��y��Η,D`Cf�$n�n-�%f����>1҉Nm?Q�%�\u��e�)]�ڡ: O�_�<��(�,"�6*�I��X�6ِ&(�C�<��R�#E*a� !�䀐�<y$)�CO�� �K�� �2�+�ov�<)A��;,4�U�Ӝ+B8<c ��r�<�1ǉ� 4E ��A�"�0�Vr�'6�1����>jT���Pe����J�P!����a��F{��rn���!����!*��X:4Xzx�,Λ"�!��t����K��>���t*^�!�$�o#��6��=܊,c��D~�!�ą/.�X�ѥ⏬-�Na0CF��&2dZ��O?�J�"x_$�jĤ�)Wԥ  ��T�<)�m�E��ҖL�Kl���k�M�<	4�VH�8�2��jT�1H�H�G�<���&6Y^Lk�� ly���� �]�<	7�S�|���pEWc�h� �\�<�F͗�%dH��B	}�̸�Uy2l���p>	��p�9����&�^����6!�� ��B�HƲh�:=�-��N$�9""O`1@cH��'K��D�E	�B��1"O�y{gǁ�3�܀��+����(�"O<�c��ҡ<Tu!@M�='��"�'� ��';ƘpP���f�{V�T�}�
�'vt�ڐ��:c�v(���S��)�'a$���G6� �vK�-I?+�%D�z@�Z>�ȍ#%n��O����g1D�T�EC#��I��E؇eq��"6f$D��;�ۻDx8c�	\�����.�D�AG��gZ��T����s�M��ݝ�y���?L&�m��[�'��)I��y�	��V��-���K��B�"�ybMŶQ�YĄ���}؆$��yRV)��ǈJ"y�Y�����y���GG���`��0�~��TeǑ�?��W�����Kr/�0d�"���a�h��o���y�"Z�I%���dC�
 R�)q% ��yb�
�t̠�)��u/��p!���y���
3J2h	�)��v��o�4�y�-Ղg�e2���^���헣�yR����l�O��[K��"�����D؃*��|B��%�:��d�CH,�[ƥ�y�HE1��J�2D���v�ʷ�yb�Xb���qdű7��M��&3�y2�/t�0-�q��4�tm�����yҧ�n�0��B�[� ��H�������>	sdWu?���0`�i��;vtҀOB}�<Iw�F�F�81ƍ�?P��h��z�<�TO�G�ޡ�2�Ć6��E��s�<�cD  ���h��
�T����j�<�r��5����LǔVT�Al�<��h�>P���@�i�n�1��L�'��š���L2R�D�Q㘜A�0�[�o'!�)Nנ��u�W�`Z,"�cҥr!�Ow�d�F�*&xǌ�9$!�$T=Sz�+�8-�����(_:!�D#�������8���zTA��R/!�J"2����� ޲�ˑ�Ͻ�R��'�O?i �PSK��3�h��q���@�H�g�<�nW:DL�	��:3�R�x I�b�<	�ǩe'��G!�8>f~+0�Z�<�VI̸n�������5K����ΌR�<�5 Ҕ!��3AW�8�bl�vʟP�<!T�Sd;p��%FhqRĪ�Qy2N�(�p>�!� �c�:��e%R�>v>�a2ɎQ�<Q'���P��'��s~�ę���L�<���� �§	kn$����L�<��*�Hݰ�� w��R�%$D�X��ł>+D��*��%-|�uB,�O�E��O�9��-Z�Vİ�ȖM��Y=�y�"O�]&�Է|��Hp@4�!c"OV�����A��ʕ�k��؀�"OB�ʢ�<M�A�O01�hPs"O
,�P�X�.�NUCb�z4���D"O�mqe#Y]�d� ��@�iE�DB��	����~27@X0e�ؠ��A�O�\���g�C�<�ǃD�2$IWS/�<Q�"l�g�<A��ןo|92򍐑K��8���}�<���ϦQ=��Q�
$����+�a�<���9̢�iˆ+V!2e$�`�<��oR!Q���'�Ļ>��Y�fEß���j&�S�OI4��Rep�,ЧO�Bc�M�4"OX`�,B�B��<+& (�)u"O� �XG��$��x3n@:a�.q:�"O��`2���ex�J=G|��"Op�rW�L>S�����;4�Р�4"O�hr�n�Q�΍(q*�� x��V�d��M;�Obu 2�ͳ
h~Y��IB��c�"O.pr�Io�z�#���%����Q"O����&	)Wb���&H�H�q�"O� �X�0�썒��[��Y�"O�UM���+͊(��T���Nx��e��"�n
���ZR/ĿW����3H!D�)�%-b%bC���dp��`�#D����⑓��C0�IU��wA>D�q�O�yz��CE�WmB� �?D��{r�6bL��$� �3�F�M=D����Ϛ ]�.,� .�
o��E=ړ
�D����`>�T! 9?Z(Бp���yG+V�I;'#��9�M�l��yBÚ5�|4�E��(]�`��DT��yR �*JB����[3"��Nޒ�y�"g��裌��H g����y�R�d2� jE%�^`r�ܑ�?��l�]������&��"bi��Bu�ޭ?۠�:��'D�l!m;/K<-�bG'[�L���'(D���HO��
ࣧ������*D�p�#��'h���D�BF�1@6�3D���-�d��ɳ.T8*��]��`0D��X�G�$E�(8c�7/r>d���<Y�Sb8���ч9I���ф9 ~���)D�(���-��Qr�9�Z���(D�(�.E.8�2��mQ�xeN��4D�$�2.W�I�,9����H)3o4D�4��j���`H���5Ԅq�g3�Oz�p��O��rԤ56�����JQ�N`x�A"Od�0�����M���_{��ɀ"Od	yV/�NH�a�M���W"O����>1���"`���""O����(!f�Y,1�Q�w
̎�y��Ξq18e(B�����d�&�hO�CD���:�h$�E�{�V���W /��B�	�\>xܪvdN�l&K̅b�V��1"O�����b�*0�0`ȶ&�8Di"O��Q��_���$�P��t"O(P�7EΤ"$9(���L�9�"O��	��0g�$8��5h@�d�'�0������Vk��P���
�2��� h<��x�]�ޅ&�1��C@���ȓ^f�P8e�bD��R�Go	.���QH�)k��L�'<�è$f|��ȓSX��� �X4X�B�x��ZC"��gt��4��4�l�q$dԜ	)J��'�.I�e��@@��68��X��W&���ȓt�Jp`G�:zG�YCc�@�oʝ�ȓP%������+'9����-�P�
E�ȓ=��,�!*F5��4�U�G8m�=��X.�8q�^�%�Z�2�"N	c�<	����}��	8
X��OR>�bJ�5��C� ,0��5l۬ļu�� ?w�*C�	�+XZ����:(�H�'�1Xt�B�	#Plj�j��G�Q0H�B`�ж|�B䉩�D�:�G_�&}ZQ��a�a�hB�cU�E1F��2P:��BV�=�)�j�OD�[Ƃ�4� ��tB��;�@I��'ۂqj2�ӬL�h�B�1�v�(�'�Hl"1�%I�@{���}�J�x��� �Ð�V�f�賓�*Yܪໂ"O� ���6j�F�� F�@L�t"ODL2w���z��p!N�C��%i��'x�R���ӡ��\C�ȇ6~�$L�I�+C�|��<E�	:�I�Aߢ�L�4�^̆ȓYҘy��!�#��؃�R�dԅȓVi��ע�$m�|K���;�&I�ȓ��zC�G�
A&�q��O�q�*��ȓK���΃6���KL,��'�$��W��*r�b���Qe��\��ȓ������S������ۥ�꜄�dC�y	���+��l
3��%򪑄�O\Ea�i`OV�26���i�ȓ�Ф���R�<��Z�+��p���	�m~��ɶR���H;7�Y��@�7M:C�	 v^�� %P"���b���<C�	*+��m�F�פ�����B�\�|B�		�;�T	.p�Ѐw
xdB剷=ex��w���%W��2��V�@�!�$[��=���XT�2`��_�ўаt/)�5�~�xR�e�px[5$W?v�L�ȓ]�PP��{lB�!�M\�uT1��9?Sq�j�E�Fg�
>ε���Nl!�����	�$��&���ȓ�2��%B&��m(�չ\5N-��!�4R#)��C��ř���3=8|T���Jm�"<E��CL8�S3�ZMc&f�rh2"O� Iwb�bT�A���s�!Sb"O���⏿E�u�r��7���E"O�s��4 _��)֋��E�4�t"O�Y�B�%������D�OPp�F�ޠU�����/<�z@!�f���'{��n�,��'z��z���B������� 8#� ѻ,O`���OL�䐠G����;=�2��	'@������!B�D`���L��I�]W��">���F?�TI��+U$ �j2�j�U*ld�eb�rj�%T1r�S��à�(���jD�$�Oc>��pj� �s������V,�<!�hp[�e8;�[�8�H���0��D�j�@%�#�"4��#%兪T�剟8	&\��ԟ0�'c��П4�I�!�<�Մ�4���: �g����ɷu"0\9 �~q `ī`�"�	!��u�O��� DCO=9�(��D�Ν�`�'d*�@L�!|���P�(L,؈ )�eB���x�}�`=&�(����%*p����<Y�����	M~J~*�O�sTAM8 �dQ���jޠ�E"O&E��Ǆ�T5"0Q�*�i��]!����ȟ�`�d�}،�ʹ-�lK��OL���OF��C��(<��d�OL�d�O`�)�O&{`B�k`�C�Ş������Q�1Oem9fiZ|j@F\�*;���O�b���G�Kf��R�D��VQ�5`�[$G萰� ��H].c��&Yt�'x�x�)6,i~��G�.��]zGLZ)-"|e��D��dX�Rz2�'�ў�� sщ��T��)�+c�)�� %���fM�'A;�A��]�S>��I��HO���O�ʓV�8"�8OȲh�� �媀����7y�ڀs���?����?Q���?9�����F�����')��DU�	�N�-���8Aa��*�haGC�
6��&#�H�'D8i�酞A��]!�l�1g=tE ga�A�Qiۇ0����E�@x��q���O��Ñ�'S h�wd�����F�	fE�yzD�'vў�E|�����[�:FJ'oH�o<R�ȓKyL��dJԒV�����Q�T2Bx�'��6M�O2�\�9��N��i���4�\JЊ����_&��B�_-�?a@���?q��?1Q�2ۦ0��U�gH8��|�Cn^�w$T����G�x��1G�[H�')bH���Rf����Y�C��8�*tH�	YoS�M8 �	�7�4���ORc>��F��d��ط�̝US�(�b&�<�[��!a�ϔ}yx����l&q��I��d�-c�F�C��1xI��	�H9[��O�4ِ�9���?�	�K��v=R-��YvJ�$�C��&��c�p�uy#�;�PC�I?I�8��p��l`�E$	�S��B�)� (������huRb
�z0��B"OȌB���B��юV�0���
�"O���m��T�A-�)�LtR �Q�O^�}��W��p�b
n�13��+�䑆ȓHg�%�F�X�-6N���7�
@�ȓc�n�A!�N�1D�Yۡ��N�F��ȓ`y��P�LyI6i`ceٱeT��ȓ!��kPck�X���/)Ϫ��ȓo.R���:p��+%l�6.p���&>����$ۊe��	I��3ΰmƦ��C��G�=��*��L�x0��1|�fC�	<�q���ɻ4��ك�6YbC��'e�L�ȀGH&3Ȫ�(���u�VC�I�7�ȳ�A�A�0��g����	Z�P�'N28�N�
f�@�n@�r��U��i�'n�d��'w��'��h�u���~?�iK ���a��7-��uw�E:G��pW-_�8�����m��O����fekA��-�p��)I0��*���E����0���(6��  ���On�d-擔6��[Hsj�󷥍�PI��0?�p�-���R	��
.ȵ�V�U@x�H)O��J  ��m�-��N�?a����^���I�����|�'������� ������JMm��	U�'�ў����ʄn��z��X�?�l�!�
:�Ɍ>�Oxb?�1��6��	{c�@4xЊ7M;?��OԂǒ>��y�M�x�0T�T�ؔY��$�$��Lk��8�O���@�,}�� 񩄒N583-�I���g�ER�B(K���'��>牎^D@��6��?Rɒ�[$DT,����U�+}�h+}�������i�h�@
�m��\1^�a�F:Dh�aK$��ɍr�Т� c֤j��q���J҇�]�?Q!��S��@��r3�_��,���L�%���p	TⓂ��:$��`��?5�"���CV��r`����XSv����~�$	���|�fL�Z���?��n?'�)S��JV�͑�a�7M�d�'��H��O��B��i�8�z���պX�r�yrc�_�mV[?t�MS~ʟ��T������8팯[c�1�ԡ�>k2ie؟�أ���]�������,P��5D�4��>`����Ĉ)���e�4ғ��'�"�'�Paɳg�~�ap��X)/�	��Ʊ>�K>1��T?��\M/�4Ys��/ZHX�
�M�y"b"F(�(Q��|{��Yw����y��Q��Ь1b�������V�yR��0
����!���Zgm^��y����X�v�֕��`6�U��y��?dZxU�0JM��Ys0���y�O�!ҹ�w�>J��5�FN��y�Bߙ�J�[fF0,�,bvl��y2�� �FAqf��?W&^�yBM9�y��fL ��g�RI��P�fA��y�n�r`���XEN���!�U��yB!��$�����-g����f؝�y�-�:��0�&��2	�6iy�����'n�}¦l�-q:����m�!r���"b֎��7a����̀>њ��͎�X��@�
��%�4��Q,�?�48��b*�8��Qˍ$,�jH�0ʁ�!0N12L�!?���b�L>`���h"�7gp����
'*���fiɓ϶���6$^lq�1�'T�j�O��&Ď��*p�c£
�ؘa�IBx�X� Ϥn��Y`�ƥC�Ĉ�'.D����a��L����FR�ZLK��*D��8�ˌgY��2A��(�l���&D�0HrKM,>� �����Ufh�A:D���-�=NZ���Al8}"�6D��A6���zV��x��A5D�X�a�'7#��;Gb 6���HT�1D�T��,˕1�VP�H�U�r��u�-D��{���Q"��J��c.Bգwb*D�`XDA�)i@�r�CU�HWڰЫ&D�8�#-�,qF,���2 c��d�#D�P���ѮVxz��Q.(d�v��+#D�� �d���K�?�r��O�9���"O�1*�c��z�����i���e"O�0q�/��Haܵ�W"z,Y�"O���ōT|�����v,�1{#"OV�K��.ঔ�vA�;����"O`HЊP�\���h@o�!o�&��"O��i�˲8�EKȗ'���g"OT����>Q�M���M8p�d�y'"O �P1��� *���.,-:x1C"O����D�n�x @��Q"O�(��$�1}-N0DŒ�N�aQ"OL�`b�Q�q���S:Z-���U"O�(��\"��� GŮ/ (�"Ox(P��I�2�QO�&2�T� "OЌ�E,R+ e�M�;�*�"O��з=l�3�^�v�Y1�"O:� ���0��V�]-O�0�h�"O,�)�j]�s>a��	33�"O��Ħ�ck"M�'X�c͎h�s"O>�S0-N|>����׆�b�"Ov�h5��0s�����0�J��A"O��9�b"+UJa�����a"O~����&��!���A����"O���3!}Luk�	̀��]C�"OHa�@Í�%]�պ��\�m7T��"O�Y�if~�u�'�V��"O.AS
��O+(� f╖��ڑ"O�E�*讁(C�W$+O�"O���P�ӧh����HQ�(�c"O4͘�JW>�<�k��/�x�"O�Q���k�8hKed�lG���U"O��B���NV �A�BJ�J��ܑ�"Op��`c�$����ʠS���*a"O`s�V�p�T���W?{����S"O`���# ���h"�t���"O2��U�R���0c�� D����4"O�ѱ��8&^`�"��>m"�ݨ�"Oz��cOC�*�$ɣR�V�IT+w"O�=�@CY8@��O
�)���a"O�l ���[�(Ĺa㛃V�z�#"On}�A�C�R��$A�4�T"OX�VF��)6��86bׁ_p�yC"O����%�GY{��X�eD`M�5"OzH1�ㅅ��A�" P�q�-Q"Op(s��2;j4��W,��G��K�"O]rRo� ^j��&��CӾy�"O�Pq�b�&E��@
!'}
"Opa����{��8�&k��^4� 8�"O�y2Vㄺ���E�?��J�"O�ev�_�d[49:���dĳ0"OV���D	)C���eش&�x��"O"�3� T�/V�C�ot ��"Od@c�I'C�	LY`��"O�D�$@B��y�e�D�ȫ�"OO�դH� ն��gA��y�Hʐ%������C���Lkf$��y2F̛X5�)1g۲|��ı�$�y�!�*n�0�Q�b�+�|�a.�+�y$��H�~YA��n\��sH��y��/}Π�Hs��b=�t"$ۚ�yrl�.�dD�QIюU5lK�+A��yR�7
�h�b���L�,��'%��y�Ws�~��&L����7����ybH�W�N�2��_B������y
� ��P2 �Yk�%���ƈt�~���"Oލ���'Y�Bq�2�¡Q#���"ON��	ڵ7��Q��Fdaː"O|�3l˰A��PS�ζ:i�)"OVѪ5��%,iR%q�nT�tc���u"O���Z!(�� p�+�%��)�"ON�R�e��jg�X�
��V�`l{�"Oxq�J�g�@���5��Eڐ"O�$��>���ףĭ$�b�H7"O��* MF�G�u�5h�o����C"O���#�P~ ,�(4�ͮ�HT�"O�T����-��,�t��O��mE"OZ����ւU1D嫒cU�t�$�s"O^����1$��y��A~�U�"O���g�A���{��
�{F��"O�������H3a��"CV000"O�U2�^�>�B�Ceꑑ\2�x#"O����P?lq:5��O6��"O,�����(�J�RL�5Z/�X��"O�hR󀑴C\~,�jߪk���@"O�չ�f� Bh`��)��7�LԘf"OvK��&-v�:���9�B�8�"O��'��OU\��ՏFK�483�"OpL"��)+$T�z��:@��z%"O:���$B1eAZ��6*�p�<�[�"O�T�t��|t`4I1�Ƚqˮۂ"O�\Z�\9CA�YHUO,Wa
%3�"O����ރXb �@.�(#�(�"O����GZ�v�X�C�Q-Ӛ )a"O��O1�>Pr���W��)"O&ؚ�ƋZ������3|�p���"Ol�A�k՜W��G�)*��â"O�a���rWT@T�&�v%�v"Ov,���a��D�o4!A"O�Ɂ����Qj�
wރ>C�-��"O8�)g��*\%�
@]:���"O���"NF�gj88��Z�k�ȩ�"O��BC���a��8@��* ���f"O����n�n��'��Z����"O��!��h�T1�G��W�д �"O�l���B�Y�<-zD;��	C�"Ovy�B�X6&	�5��#�P���"Ot�#��U��� x�̯F�-�v"O�`���G�.!0@��8'~�k�"O��n'��tcl�)s��q!c"O�h������R��ǻBB*��3"O�D��Eՙ;L�X{egՉ)4x��"O���'��Z�2�[�^�=��Cb"O�$qC->A�5�C�(F��p�"O�����2*H��$�K6u�t�K�"O�M��EQ�q�5�2ۜl(�*O��'邉=C����b�W\+
�'Dv�r�E���gI�!xF��'�vu�q�ջ�.�" !�����'�F=j�M�-W�Q���ދh��j�'�����=u=�q�ʼft���'��% EQ�ڍ��mޛV��Y�'�����@�_�fe	��P3TZ�-��'˖C�
�O,���V��B��C
�'uR�ӂ��'&��aN'�r����01펩Z���h�Ϝ[
�'!^�ze*�.
\�BqnZ�\n�@
�'��t� t��|����&o�Y	�'HD��V��?fLm9S��F���� @�`�])^2�e�d�c�"O�ȑ%�3�L��PТy�F��"O�<�t�L�a�pdM�|-:H�"Oz$�bO���C���<��B"O��p&�=��RTEʓy�T�q"Of<�b↑4�"���M]���	S�"O(-1��3$Xm���q˂��"O�d�-���3�ǴJT>Hh�"O������3*��b�l�wD:�`�"O���4Hú0��I!�K7�[�"O܌#0�Ӓ�(P�@j݊=�p4:�"O� �b��`>T�J-8@���"O��9e��5�Af/N�W*0q��"Ol!�CM�d�1�/	�D��s"O�1���V�AmF,���()�x���"OnU��)���i�(��M�"��"OH�C)�-Q�N�'R�<I�"O�%�W�� 0H��r�&�\�"ODIٔK�m0��Ci�<Y�v��"O��V���	�vD�3�ˢ9���p"O�t ���+}�R�S�~�,��a"O8�Q�˥@�2a٦�FH�\���"O�8
��$*{2s!�^1d�h�H�"O��y$��
3��*���/{`]p"O�+�
SUt��m�T"O�!v)V�T��y�3�[0-_* �f"Od��7���P6>0��Ù�;��)A�"O��Q�X�(ȅ��	YΜ�:�"O8x�bW [����@-��,�C"O�m�u`�+t�@�MN�fL"ZR"Od�wM�-ilts���X7J�"O�p����n��ِ5mT��H�A"O\�j�BU5��yUꎗ8�h�"O��Xu`�7 �|R��4m�ѩ"O�@{V�U�"��"Ā���Ѷ"O�!6mַ��Q��%�<��"OP(��_g8�(��b:�d�C"OBm���R=w%���1BE*z2:TS�"Op�aC&P�>�"�hG���x�+�"O���0��2"(��2W���.pPI�Q"O��R�� W��q�S���h_d��"O�p"w
,{�6	��ϯ,Zp�:d"OT4*���Z�ֱ0�%�}Qp=��"Od�(�+�M_ �q$F�>���c"O8ݩ� �%q(W-I���q����yr̦V�U�Lď.���k�G�h�<��P��j=R�.�C4�x��.�i�<y�	Ȓ�\9ȥG��AP�Hq�<	u��*rK��p�`ƪӒxy�-�o�<��R����'�V�h(��ۂ��n�<y1`�g@-�B�<�L ���h�<ё���3U�@��J+���t�f�<	�H(p����X�<� �1&��y�<�'�2
L `�ڢTa)���a�<��JX�����ݜ*I�"�_�<�J�li��pbAN��QdI_�<�#.sZ�a�⠘���XQ�Q[ܓy�Ԭ�ЬE8�����'�,�%��i�삌i�P1%��6x0��:$'/D�@�b�:2j�ܑ�ئZ�Z}Q�!D��`�o�Tx�a�G����*O�l�F�O�{�YPB�� �x}��"O.�q `�0ā�,@���2"O����G��С% مq��`""O���t+�v������| �*���y
� 0�@fH� Le1�Ŝt�B��t"Op��%�d�"���%֭tߠ:"O��X�ǔ��h����#!�I��"O��pB�� E�ڔcD������E"OX=��M��/ڶ���*�	J�q2"O0-(u���R"��8
��2���Q�"O8���M�g�.��ЃZ��) s"O�p�'���?���b�CP7la�I�!"O�}C���+,I��HJ�xE<}��"O����c��|;�Ua�����"O*@��oX�L��\�.�&l�ԍ9"O�y� iƘpQ\�"� 2T��=+�"O�yzF!�	G�t$�W�� ����"O�iچ��|�\�Y�BJ�r��Ȱ"O ٗ �%m#�8�@C/5l�L�X�<1��R*u�豃޸^>N���c�\�<2LR�G4���
�9�4M�t��`�<צ�!?�\i�"� �<�qS�
G�<iǠ�_6�5,���2���c� B�	�%X�eҷ��;_� bu�E?B�d�p ���4.�b�X<'0PB�ɸT�
@:r�˦q�L���,.gA�C�	�o%HX��}�p(@�tŘr�'*l�0glI:Y�1Rc��OުT�'G��#UL°ilf ��JNL!X�'�<�K��aϖ)�5�ȸG��9[	�'G0���&zdd��M;L4�a�'VF��Deڴvqx���H,B�T4��'�"�)uG�� ���cW0>!8�'�-c�/�k.e룁�"����'\���Ǉ�5c7�@�F֞XR�*�'��8z��X[tU�h�1:���'�@�G�?9(�W�ܜ7�!	�'>���V���r�6qj���1���8�'�X�aR般Q�Z��рNP萫�'�\��E;ޖr'�9ox�0��'{<y�e&��T Y�HW�d�ʼ 	�'�N�cc�m����sǎ�nV�Y�'���a`��J�����Yz���'rT]��&X<����	�O$��	�'�z���L�}},��-_ L�Q��'���%��z��a����B)�|��'��K�E�l�`5�`%)�B���'G^xU`;�l3&^2w���q�'E�D�"�$CH���,m��'^.-h$cW�^�~)��d�4A�0��'Z��D�4�� }r���
�'A�8��h��J��f��o�Ȩb
�'��r�N^�)�`X�AB{�(��'B�Y��'�-u�8	��쇷p�^���'��t(�hI�65
�������
�'֪�r^� j��S�l�����'(��;��D���]x��1^��}y�'��t�d,��A��AcF�\�����'ͦ}��
Ì���!c�=Pzyc�'O8��ߛaU~��E犢is��'�|1SM+-K���䣊�DA���ȓv��z���1yǰ��`�B<h�lЇ�� dkTY3p�`L1N�Af����a;Q�БTH1�u�͊s�D��s�9�6I��Ĳr@�-C�6���W�����À-;�j)*�X&'�T ��E�re�p, 5'a��I�#j@���^+l�3`Q��-a�.��{��͆�S�? �D����SH��Г�T'A�|��"ODt�m����h����\���b"O�QQ�aוe�ư�˞&~��s�"O�h�1�No�p,X�#�
#�tX�"O.���h@^L5xc�.=���*`"O�IBFb�4DL�yv���tY�5"O�ly��/��Ԩ��4��"O���W.9b�2��L�=�D��b"O i��b�#' �1.@�e��-�"Oހ�@��J|z�K'l�gN����"OZ!q�.V4;�<�"cbTa�F���"O��ѱ@�8$��,�GE�X��m�g"O m�6jI<I��1۰aF!EW�bP"O���dc�v�� ��02��1"O����6 �������$*�2"O��ց�M�ʁ	�̓(#w�p�"O4a��GU!e[��c텦D�|0�"Oܽ�b]�yC61�`e�
a���W"O�!�M�y�(�if�D�J4��"O҄�3b	��D4@b��Q )c"O�C4욃f�4���I�J��"O��2��ɹ{�ZM���*jR�# "O��#s�^�tRRX;DK%bj4I"OB��1BU��Pacr��IM�@e"Oj9�*ީ'za���q��Xr"O�<)Æ �,��	��]6E_�p��"O^X�'�P4+�YABL|���"O
X�t�%3�-qUA�Eʴ�P0"O�Ը�m^76�L��'V���8�"O�$Ƒ�2�z��� �K>��3"OP�;(XXH4[�E�
pj��"O.�s5��	��)���T��1#�"O�I�H�U="9���/ߴ�s�"Od�#Bd/�:]��0<���b"O��0G!��LE�|�ŇϥP0h�kt"Ol�� �ȍ��(��d�!	7X��U"O�US��_V켹V�MR����"O8Q+l��:xX��"�$��v"O���7ꂚ��1�D�P�J}�8p�"O@�W�S�<����%6�4��"Ot�H�	 V�d�H ��9bf"O �B��⺵�眃�J��3"O�P0��t�U�U%�2!�֘��"O��)ňr,$+��7P�H�7"O>9c�dw�~-qAj?Q"ୢ�"Oh�r��؆h�tE+�(I�pau"Oez��7N�#T�Y��`�3"O,�i4��1.JQA�M+I�b�� "O"����Y��@K��	�e�na�3"O�xJ�2R�ah5�
!k
�E�g"O�t�AdKj�t��왕t(X��"O �2	B�~*�)I"E��]b��pU"O�C�F]&9�j욲ˋ�d=���"O�0�AC-pcr�� ��{|=�%"O�8��)M<0s�i�@�r��1�"O�)Jp��1f�*7g�.Y�D���"O���%K�{D��@�E#��j"O:ؠE�)R,�p�O��Y6�(�"OlQ�`��{?�l�Ä�y%�t�"O$=��^7��!󇢊�M@���"O� (Q�&wH2�1&��2L�@�"Ot�����~Ā�v�"B|}�"O��Z���Z���X�`X����"Oj0:M�	If1��cU$,_hI�f"O� xl�@�f$�E��Q�TB��""O�͋B�]ۘ�X@��f�YH6"O�-�����怙�S(�&}��"O��9p��3`�@X`��2;V�"Odm�4��(BY��^=+mH�!�"OJ���D�h_� h�N)T9T�u"O0X��'�%V���4-]�<34��"OTA��X�E��@�F,1TŐ�"Oܘj�)A2{�D�hV�T�2P�ȓblܱ��!V��P�%`ڿF��|������щ6���y�eć.���ȓ2H����.r�$Tw��n���!Ӑ���Ѐoa���vh=8�`�ȓD�H�!�)m��8a��A,	\���ȓ7��BR4�tY�SI�*Q↩�ȓ{l�;�հ�ĵ! M�R��(�ȓ�T�����;��Ȃ5C� �ȓvǖ���f	qx�q��|9��}����$�/q�*컷mҚ(6h}�ȓo(d(�KĢ#��[ ���@�ȓh�����*r�2�AC<�ȓZV|�[DE@>L*�jd�@�j��m�ȓCx~���d�*re��H�� {T	��04�Rp'�����S�/����+����U�N6]|��dO�0ʐi���"��U�V�s����TeL�T��-�ȓ(j��h�M�n�&�üi�*х�7v9p��S��1���K�$�ȓ]�2�tp؂H�i�c�`�ȓU�V�cCJ�1m.����Ԓ/K�e�ȓq�Q�!��~#�M��A�Bh��V�( #`bN'G����1�Ss���ȓڂHRĬA�T�HP��Ї��i��Z�$���(�+��Y����4l|���5<T�D��`�A��!ɚ���1�R�3#.��کP�A]-�Ɲ�ȓb=��$���ȳA��'��m�ȓPQ���gA+TR0xs�Y+E)��Lx,�FTq�(� _t�ԅ�K��֌��d��s��
L/8���P�8��(� ���"CTB��ȓ_�`���/*w|��񃀟1i�d��,�. Pv郅E�H���K��*g����;�Tt��'%%�`��B_�-�Z��ȓb���Y�A�0-���A6#����d��i�F:(Z,J�,� p*����Yr*`Q�&�y�V*�m�m�������giԧ_� ���x��5�ȓw#��s��m�`�R�� )�Ň�n<$�'��5H���C����ẍ́ȓ1X)�P`Q�y[\Kfƃ�v�*u��@2,iz%O	, �6���f�8�d�ȓK|���¥�~����A��`���{X���-��d~���!�T�0�ȓ*� �SkU,�0�"�A1Dh�ȓ�֕3f�Ɠq��Yp��96���l�N))�g��03��h\+`���XΤw�3vX�@@�̞=�p͇�q�έ!(5	�Jq���`[.�ȓW#�� 5�3��XPwB��,uL��jy�Xe�X �ə!�ׇ2���=���K� �Q��j�:�b @�I�\�	�g��A����?9J(x[�K`�C�I�F^ȸy�A2pQ�Z�I����C�ɐx�7�H���}��,9i��C�)� n�@1'ZG1<	�1Ĉ2v����"O�zG��gj�Sc�]AFL�G"O
��K�FIl�ۂaS�*<��G"O��@��	6��lx �-����"O�I���:|�� �E��J$���3"O4���ɕ 2D�PnHP66��"Ov�
 �1C����mp'V��"O��� 6N{��r�e�BL�!���+~�٢�d�nc�T���T�!�d����s�-�(-]+J˚$���ȓ<Fj��q��:#�P�j�犑{�*@�ȓcl�{��oT}
v�]�v=�����!��Np&e�$�@�2�d���!�p���~t�t������a���ڥ�wf3.Uj�	1j�:>w���gF�Z�	�(j�z�*�K��J[a"O�7�^��@L��`�o�̅ "O��B�*!�Ip�����s"O�U
4��^(��7Ξ�E*]!"O�Er(���a�'k�)d'�<K�"Oċ����V��j }d`�d"O��	��
g�P��D�ñ?=*�q�"OL�zS���G���(�=;���"O�q�F�]6�u�#R�B/�%�S"O`��֮�k�yCU��Ы"O�{�ʘ/Q��7��<_�٘"O�E����4�L�G�	�kSV���"O� � X����#��8:�t#�"O�����*{,�P�ac�?p̕�"OJp����$�d"`�1
�$�&"O2�#��$]����vR�}�h�`�"O8ȓ�d�#�UaQ������	7"O
I��B�I%Jy�`�C�A}x���"Oz�e�?ÞM���L�e��"OB�O�	�5cHXԖ(�"O��	\�t@{�j�
L�ʉ��@� �y�#ֱDŲ�;',�*@����y��7�X�� �f[ ��f�՗�y&�*�T9*S($/?d�a�́�yr����N{��-)��A �,�y�I�'u���S!�H�6�B��y|�@�\(�J�KF�nK|�a��5D��!�lL�f��(��mD�qz��ZHB�	�7�2H��%C||`�ch�5}2�C�Ɏx!�͙�gV�g&L`��&"��C��;qu��� ��F6dq�k˛��C�	_��b��~'�@3�Ŋ�RlC�Ip�b�*�C%s�p�!�J `C�i�� V�@?���W!��U�m��'rz�S툼n�()7ŏ4���'4x�1�g�<�8<�'�A!u�,A�'l��`�F�?� !�J�|�����'x#�!uA��K�o�Lb	{�'�B���1S�L��ECT'�m�'�\x��Q$״̳�
��Wu*-��'�z����%:h�B�ՖR��|��'9����C�c�Z� �d�;%�Ex�'����Diو@���4e�n �
�'l��b�-D�oݶ����оeB<��	�'�jw&�;h>���
Y l�X�'a�M3�Iscԅ�&�Ĺ�
�'l��悍?���`��t��);	�'�b���ŢU��K�
;t����'>̭���7v(�B�F�x8���� D�C�՞>؎\"�B��$���['"O��"D�6L��� ��*Mʠ��$"O���P�����b��_�ڡ�A"O������0Z�	K�E��I� "O��,���1�??Fz�#"O�@��nF�T��T�@l�㬽��"O���R�M�B-hƭO�����"O~- '�#A�~l�"M��?&���"O�� +��3��@��[��Ÿ�'�t�PCn�1'��;�I�2V���'ܔ)�͗�)�F-S���<YF�h�'��bA�4XKvA_:Xv����'�.�LO6Y�$�Vc�8J�8��'��X�mɉ�}�����LQC&C�I8�d�+�� �TEy��ǜo?�B�əY.E���D�3+B�$d��6��B�Ʉ_d3�Ĕ�D�R�U*l4�B�I=$��0�&HI��9
�	�>�dC�	A����B�8^?�ո �$o�DC�	�M����dl\\jP�0�f��y�h�,� �A��Q�"-G�4�y� �
؈$i�D�
O�����7�y���+�D�h���^/�M�s���y��߁xQ�鱇*P6[8����)H��y� � PyD��!\*<���D�yR�¤n���S`"�=�� ��
O�yBHR)H[°r�Ț�5i��A3��,�yr�4D�l�#B**2Xɓe
��yLF\tA�1���zjxГN��y2�S�*�x�*6(�8lDIᢄ���y�͑��
��ƫչLu�d�� ��yR�қ/o�M�ե�;@hIs� 
�yb�^�Lz���!�L:D������y��sQ��4IN�`��ҡ����yB�=
�D�8�gS(eb0�t��3�y��ʡ���C���$%ҹb����yBT�S��]��'�3�phB���yr�'�r��eUI��@#��-�y��ԣ]�N<���:.~ET�ھ�yRj�"[l��チۃ@�:H��HD��y&�=v�^���,2A��ra��y��U;(|u���M-�Ȍpc�Ґ�yBD޶*L�$@3f)�f������y2cB�2\0��!�S�P�J���y��,Q���Cʸ�$a:3�J��y�*F6�|M3Vʍ=[MJ�K���y�-�wc�a�j��r$�2�u��jb6��E�$��eG4�.mE{��'e�<�EA��b��"�.D������'��������<|��Ɠ�K� 3
�'͠T�g J$#���8���F��ِ�'v��K��uH���@�˭;�^|(�'r~0�!�Is�\�0ē1�䔚�'ƴu F��0SCE˗JŻ;����'�L���d�&e_� ����/߂a�'4��"�柼<U"u+���j����'b�!��ȏ ����#:�L��'v�DA_�C*�� ��^�7��
�'(nsVB_�3PNtc2H^� !��'��)*��۔+`F�c!hz1lX�	�'�@=R���lD	Q��E����'n��4�Z�y�R�c��R�Iu�Tr�'~����4�����˼,�\���'�ʴ��kF$x���2#b�9vIZ��� ����2(~�}3�E�%F}�Q"Op͒4fV|
��z%�O-Nu��"O@��T��[jDMѥoSO��(`C"O�b��0I��m�����b#"O�T��'I�����=�Rq�V"OΑ��F;O F�lǘ:���w"O��؃IĤ}J\@�X6ry���"OBqc��A�#C�끊L�,��9"�"Ob5y��w�j9����O�d	XT"OzBB�̜����3�Ƞn�ԵH�"Of����n�AƩ��k��E��"O�!�a��)�B!BFW�n�.T0�"O��h�,Z7v����V�*��yE"O.D��Ϝ1V�b����9y�j9XW"O��Z�@qS|��R2A� ���"O��J��t#�#��ԅ.�j�@'"O�F��L������3�f��d"O���b-�X2h�"j�$|�X�J�"O.����yY�݀�		U�r�R�"O\4��P�V���P3*I*F���@�"O( 2'����j�O΄Jä�Ȳ"O.�I��Ӷzܜct���K�0Y[E"O���ܲD#l��B����`�q"O6=��I8RxC�+ʹ�`	2"O�����͜̡ 'k(d�|t� "O8�;� XE
�a���\(���"O�h�!�O#Uy�pbŗ}�(�e"O$D�kQ/sT"�"
+� �R�"O�U�e���Fo�����!�"O���P�7�`��E�}��@y�"O���ukA� �>zP�ƦTR"O���?PJޝ1��NM�y��"O�tB�� 
a��d�U�I(�R�"O`�{S���12��3aX� �8"Oh��F*l�.��D#a��a"O�hk�&IY�D��/�/Y���"O��i�-
�c��@� _�t�r"O
�$%@�J�d���P�(�ޤ�$"O�Hr�S�Ah�X�c�:����"OL@�B��Gr1�r�D$�<1��"O���S��^����GO]$`����!"O�%�pe1��0�X�u����'��,1�рO$��+��E�:zT���'��=���˯q�4e�th@,
pdh�'�>q����`E�����$�9�'�L@�Аt\ĉ��͜	E�d��'�^�D���r�|#0�֒v*��'� �X�oX�9���<YL���'�e@�#�5� z��S�3�*x�'�t!�E�-?��x�`��%S�Ё�'�Z�
�jW���H��"ـX0�'��P�)8����F��d���'"D�GiT���Z�+HJ���'��U�h��'�fx9%�����'�\��H��0����̘�2k>���'�$\R���.�f�+���.?X(�	�'�Z,"`��?Ш���D�M�($��'h�e"!CU����r�[�K�Uk�'�T%�i�-1��K�K�P�Z0y
�'b:�@�-��"Ud�W�Id�y	�'�2 `�'�x; �ޟLA�'�,�g������7���z�/6D��b��P#�,X�D�:i*��2D��I3h]�upt2�BK$i#���+D�� <�2���!%P`�%�@;q[�m��"OV|�в2ǢYB�B%l��"O�$�#ШJ�v��BX�i��Y1b"O�h"�
��'��y5�I���!�c"Od\���0�L��D"�C� �J�"O V�#tR�`�b�C��x"�gLj�<a`Ş�\�b�	�1]�1
"ʝf�<ө�	&��d@�g��h�V�kł�L�<9��_9/ (Q��׼*$D���D~�<ّ�U�lϤ5����5u�jt�6Oo�<9gJO==��8y�-������R�<�7�
�#@���� Z�<�a �%. @�fnՉ(�ȝ	�N[M�<ဢ��@)Ze�e�Ӌ{Zl,��Qq�<�,S��IZ�`�/q�A�J�i�<	�� �&P�R��ۄ	�F� ���]�<ц�*Y� i�6<��T�G�[�<I�ݾ'�ݒ׈��%�r�`�T�<A'��yF`鴪��lŶ �g�[�<�g�'Q΍��A����"�Z�<a�	���ji:�lL�B"����BR�<��,�kZd�FNH�5�[GI�<q�h�
f}K'�7.����ƊB�<�]�C�� 0�kݱh9f]څ'YF�<)�x?<,k"�P�5��Q�!�}�<�2�H�'��)��Z1x�����_�<�cEċTBQ�lR-fu5�@�_\�<y���?f�N��ɚ�;
�!��T�<�gH	�4�^8;���"=+�X)V��R�<�P@G5;c�I�E
�%~���Qb��h�<���N� �� �Ŋ!h�,1�o�<a���?����%�G�a'�Hp Sm�<�ÅFG�,�#��D�CnTՊ�,�f�<y���B����eL@�JH����G�<�E sx<��5A�	4����D�O�<!�/,-$���
�#H<=��lGW�<	P�O%8�9Ο�#��R"M�Q�<���0ftq32,�?>�I#�JN�<��b�uׄ(pV��@��U��j�H�<1e/�_gp�E�hi�#�E�<��#�������^��ഈ�}�<a1��Q����{+d����M{�<I6�ȤW�\�x��O5���c�s�<�s
��v��1���2*Ѱ��I�<��b��K��:���+	a���"
[E�<��j�+:�Ma�.βW~줚�g�<��KܤE?<y0V�L�_��T
GIZ�<�&F���5-^=��8�L�A�<)o
�q���eOe)"P�N�k�C�	Hc(��"�#2q�p�ңr��C�I�Hz!SF���@�u�7�P�GۢC�	����5�� d�)��B�4E�iS���M�ָ3!�0��B�ɘq>��M$Q��;��[�u�lB�ɪ@�����aHQ�U1aO�k�.B��%FyP�F��`�v�Sv�L�>��C�I:lKpU� $]3+J���-׳-u�C�I	V!�1�*��l�(��3��n��C�	�Mdq���2{����b���B�I�]18��7`^9�d��Ə}��C�ɀ#�,��J�vo� ��L��7h�C�Ɏ4^�@�WJ̝X�fL�c_!nC�I=��0�q�E9iTi��۠@A�B�I�`[F%����o'��*p�B�)� ,Qs��$[�X[0E�(h�Yi"O��rˊ1�{^͸Q���¼�ȓYZ��/�� ǲ�0vNA?�J��ȓi��H��'g�& ��ٻ�D�ȓA����яĘt �U�Uc�:Z$����:T�а��޾?Ղ+���6W��TZ���C!PS4iR�^�����ȓVad Ⳮ�	%���5�˾Cc���ȓz�F��`��
\�oǠงȓ!���0k׷b������݁eB��ȓ�d@է�VĜ���λN�Pq�ȓ)5�s��*j�Tېƚ:jD�t��C�IA�0zf��rU�L�rZ�|�ȓXy��!�;B2j��S%�?Tie��&RTQ�fKn��Qg�7O_}��%�>�C(Z(�XuL�
v{ZX�ȓK�|� ��1n�0�iC�LV��ȓz�;���pϖ��D�a�ȓ?��y�s�"q>"�yv�KZ,9��@т=!�@�������q็ȓZ?�!�uǀJ��X��&^p3�ȓ5�}�� a�Ń�Ij0��MR6��%ČSlH�� j��i��|Y@,Eft-�aQ6�>}�ȓmɤ���c�'��=�q<�<�ȓ�9[�(�+� 2�	1
d����83慈E��7B�m�d�22�����5ΰ� ��A�P#
O7� ���$��<Z�Wk�b�@0�Y�6k�܄�F�P�
~:�I##�(Yq���ȓm����f��m�Ht��ƌ�@�2������g�ַ!p���ǥP�:�(-��BRj��$\�7��9�MY�LK,��v�d�SwmH�s0Ґ�v��aR$��N�"�a'm��7-Z`�A��?DzB�ɤTy��I���->��y�lA�/n�B�I�nK���G��:U�La���]<C�	�{N���K�?#(<)�萧w9�B�ɑ9 X���Ǝ0��a���Bj�B�	�d�F�@�o�l��%`b��B�I�a:r�c�k�+��-(P,�f8�B䉼=�����x#���fԶW��B�	7L`�M���W+T�xᨳ+�j��B�ɹ`��$�U�ۓH�)6!G+f�ZB䉽g2lY���"�"Q��㊈3�HB�I#L�hP�#��2�ElH:T�NB�$mERI��-	j2�����Ĺ<�LB�ɗ�~��`(Z���0N�6��`�'�L��G
��t���u��tX�'ހP��H�[����@��h�lm�'���wÉQ�i��?_���[�'-Ly����n�|0��@��5
	�'e�5�R0P�T��"�25�2��'�l
�_<#���n91��l��'���&�
<F��V+=�8,{�' �|*t���S��-s��� fƴ���'�N��6��l�a�&m�3t�jl�
�'}<)T��;a��{�Z�Z�pI��'�,��m���V���e�j�'`�x�  �$��a���
[�.��'�Vu���I�b�H�BQ�_	Z*a��'<���t�Z�A��2!
����'�(�cثp�"xPcS��Ԑ��'�v4#C+禙ز�AK�A��� Bm��@�=��ةV�P�Z�����"O&�"���a�|<�@ͷA����"ONA��NH>�y$c�p3F��f"O��'��!�B�����wD�z#"O� �@U,
>�33�O���0"O��j���H�ް�a`F(y���"O�����@�p�*	���>��т"O��ۇH58t��@3w����"O�+%�п4o���2O�0�\�Z�"ON�zwG��w����-�.H�쨋�"O6	���
k��5���Z$QB��"ON�#��	2K׌ ���L��|���"Ou���B'{ƪ �M<3��R"Oz�K��
l��a�G�K�"O�����]�^�)��#'��q"O��q�͛�Px#PG��Y]"�G"O,�Q�N�'je���.1��g"O��8�p:��ڲLt�チϸs!���@E��e�?-JB�f'o�!�$��k�!8ݩd��Z�\�!�D�-XO,5r���Y0�y�@�l�!򤞹k25���Х`ݐm9��"B�!��4+�8h�&^�*�0f���!�J(H����Ą�G��M!F9U�!�dW�i��,�7mB�Z➽��-�9�!�D��h���E�N�8Φ���ݙ#�!�$��"��9���'V�ʴ�޹v�!�d�%>�r�P5cB�J8���u!���~�8�6¬r���� �� e!�d�q#��� �B�W3rh�7�>M!�Ϗ��P�!�'6mf`U tK!��F�j���uC�����	5S,!�(,V2q��_
>���_!򤌸)��ݪ���]^�p���a�!�䎚:����\P\�vlb�!��/Dh$�mߗCx��Ta�4�!�K4��-xp�L�0(�|qQ��)e�!�ӆ��PD�߽�{W��	H�!�D�3'L�́��ɝ
K��De�!��ոMXdmi  � 0���@�L �j�!���zݔ��#�ʻB�xX5,��7_!�$_ |Ʈ]��J�;�N� ɍ�!�Dt������z��!'m�3�!�䂆G� �������#�%�9X�!�$w���Qnͤ�6���%�&�!��dp�1��!�&x��F8,�!�$�c�.��V݀v���&��V5!�W�e�.1H`h�	���Є̃I !�$ޗKR�`�J��w�N�K'!�l!򤜷5��ꤋ� �j%���C�D"!��@K�@p��VL�A���I�,!�$Ҫ�f��
�g?j�h�7�!��C˼����B�m����\�E�!��� pV��x3k��"U��^.$�!�Ĝ�V�)5o�\E:�C�Ѻ�!�$Q)��5{A#y2��
�S5!�$=] �	��-K!�	���!�Or����	�I��%B�`#|�!�ă�k*:L�"J�`�x��`�c�!�$V�r͢���)^"�Bm��Y��!�Dʔ���x4I�SR�\���ēy�!�d��9�q��Ą�t2�-���U�P�!�D�,6��Ұ흽6u�2Ύ�h�!�ET�T+@�� �*�LN u!�� �(��F� r�`�\��-��"O��!�@��$���Yؚa86"O>8�b�6D0� /���@p"O��9�(�m��8���M�!����"O�m���ӻs,�5�5�y��3�	���+%��<u�)�&�$���)pDj� @�7qO ��9Jb4�և�X�.���4u` �O�t���1Yf�K4�	wY�����ĦpR�Y4B�8��Hɡ��@*$��_:�9q��/uf���)�M��-���I2%����O�nZ�(�O�P��+J 5N|hPBj����E�a	�O����V�{}��hj@���d��ۤ��p>�w�i��6�f�8૱	� 9��ѫWb�4N�$�a�
�M�fV�p��	qy�O��4�x����D��d�#�9t�7L=�¬/{=,<���)z��ڂ#ܨ��O��;-�`�����9��� ۓw]P�lZ�FM�5h��=A��ncC\��I�<"k�t�|��sj��S�׮r>Yk�J�d>�o:}h����ٴ�?����il� AwJ�%����-�.���'tBT�t��	<rL�Wb��DSD�3=�#=9�4Hq�֟|�U?���I��I�eA��N:H�Q�������'{04�lZJX��@��ƂLy����-սs�����b�&����$P��A����/��H�'L1#<�Æԯ-�8�e���t�Rt�!�ܷL�Q���I(e��E*5N=)����O!�fO�d��'B>�q�3�a�&��kâq"��OJY�0��O4dlڰ'N��<�����d-+�T0�� ���HQTBѴQ�Q�P���6@��m���xiv��,uq�M�t�i�7 �����X�����$�����Q��G3��1���ox���	��P�ȱ�ٷ)ab���oMƨۗݙ+�`X�h�2n�
Š'�� J瑟@����+T�V�Ru�5+�"���a��2����LX��c�'�+��h�ūN�)'`�h��Iڦ���E�E%��5��j�jy��oӪO����O�O���h�(��k��h��آ={"	��OF��d�9^^�X��/�1T�\X���y9���	��M���?�C�i�BL�q%l�z�d�<��89_f8�a�]|��MҖ�oRT�l�ɷ Gy�1�ђI�tBG�ܯC�x��A4��a�צ`��B�AF?���i��	�C��A��]*~z܅�c��7O��;XjV���̇]��DR��?%��@��cJ�OrHi`�'-��nӐ���~B1�ֆj��h�eJ�O̬TZCN:���4�"=)1$-,%n�r��93f\�v+	z8�d�شM��i��2,ߨ[F�u/��(\���'aLĚ�jy�N�D�<�O �']�aJ&LQ>��,R H���L�.Р�ru���es|PJrCϹD`KY3�q����w����t�I!0�MV�;� ���4z�6���(9�hI:`aW=cOl��6�	:'���|��5�Bp��J�澔ˁ킒��`mZ	�����O }��r��i�ZU�eIܛv�0-���ĀME@�'�b�'��P�z��N�XLX�H����~�Q�ߴJ(���|2�OD�N"<�ik�OR;;�A��!��9�$�&����	K� ��   ?   Ĵ���	��Z�:ti�-���3��H��R�
O�ظ2�x�I[#��y�4g�Բ �I�n-s�E�_�]	p7m�䦕��4E�� ��q�	x8�Ļ��My�֠�B��H(�Qy��7U�#<Q�
~ӨP(&m�r��xp@DB4F��r5X�T�$�����1?�E���/��7�f}2*,�1��l�?)��0��0L־�iP��uy�`�OvԚ6F� ��9O��@qJ��0~
�rt�
[bZ���(��L�@���'�,��$�ȄyQ#��!Ӹ'=�TΓ�|�YՌQ�����fn��hJ�$�<�ቭ!�'���#1���{�L:�I�h$�'�Ex��|�'�!�f�N	^PH�$$��}��-��&#<���>��I˟R��X�H>C���w�Y�D���O(��{��]�Jr؉[�B��K1�=S�,�MSV�1���"<���	��pˀ�8���(��[�HI�>q�	)?n��B�9Bw��2b^�H�����<�fȕ'5��Fx"��N��|� �%�L��t��'	��F'|�1 �?�@�"<	(�O�e(����.��L8��Ev�����$Z��O�D�O<q�	�W�؜1�O�"
�j$�wL]?y�3(o&�O����*�1	�D���N`!GK5F���l~.��>(��4w��	�/^5� �O�h�q�סe�8��F.[e�0�X����M b�\c�0�'�ǁG�'�b�S�������$�C�2��ۨO�����d[3�OL���LR&����f��0��:F"OL�y��  �~�s��A�X�"Oz���P
��)�#�;(_�P�"O2��*Z��z�1!�.Q�H@"O����Ic����B	5�jS�>D���/����+-d=�@=<O^"<����.(y��-�9��Q�G�u�<�eA�<�p��範�1ZX{A	�z�<��a֋���3��(�d�J�b�<���ȃ ��q�bC�*(����o�g�<�5�fe6I�3�P"#�Qe�a�<)��ɶ,D\
�g��bA$_R�<1b ^<�~xqP�؃o\x�2'D�d�<����,�p�J�	_4���A`�<i��Vp��8�5%7NN��U�^�<�p�%i��wIBYɒ�QT �]�<qա�T�)rU��?�t���h�A�<Y`�Y�.��|�@YH:�%1�JX�<�b���h�f�;A��D	��8�EH�<�I� +2�yC�''Zbu�J     �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   �	  �  -  �  '  %/  i5  �;  B  IH  �N  �T  '[  ma  �g  �m  3t  uz  �   `� u�	����Zv)C�'ll\�0"Kz+⟈mZ�p|�57���DB���H1�ѯ&q�5��7�$�b�ی>��+�FRH XY�f��%e$���;F�FiB�'>Հ,y�'mx�a snQ�)�8=s���(-��(:0Lݧ||<Z���I<���@�'�A����4���蟺�d	�
`
�c땘,�z���0�	Z�DΐzRf��	��<��@*��ߴ+��9���?1��?a�n�>Pc�(�[\>�j��¢;����?�
�;���q*O��ğ*K�����O\�ě�a�n�AU��8C�"��%S��v�D�O��'�b,	!���C�?ٚ'9�t-K1Nz�Q�m0\�����ؗ/��2OP�Z'i��P�2���UI֥��Q��̓��'�P�2�#L�	?� �[$��)��}���/� ��O\��O���O���O�˧�y��ېj@�@SS��/m:�A�c��?���i�R6MSȟ�n�˟X�ڴpr��md�lo�Lce'������3�U1�X���J۾�HO���k6�'x S�����0�&/���v��o��@ؖ˞�x`���ڴfۛ�{��I���CwM�
P0����W�k��f`H ̂ �fyK�4c$z���� '�YP���,S�h7�5��aP�d��4l���M�V�N�0�rw�<8��1��!z]�}`pA��G^~��u�i��6��צZ���A:���v%�	Xh���M-�4�@�D����G�#`���pKJ�H����ώ�M#&�i�>6-^�q%��φD����fo��XJУӂYO\(�g�A&H"qo�����1ʉ/m���d�c5�m9U�ٟ��?�C�. �R��$�¾eu�`a'ǁ*Su���$�
����n�8�m�?���� W$�2�8�	0|�8xC#Z|���K'�5�ؽ��t2:9��(٫A�#f
�T�ȓ&�� 눓��#!�ӣMB$B剄�t��+�Xy�p@ѯ
sVB�	���'��Cf��yүY�3:B�	 
�,"
(�J0q
2"h�=Y�g]T�O�d��q�KiP����\�"2�R�'��jT"J"{Ȯ!rP�X2�X���'��:�� �ĥ�WH���
i��']�0+qo� Ub�@�7�������'ق����[z�+B	Z�wA.l�
�'5<%���hS�I���8l'4��#R��Gx��)W&��4@�T�9�%H�K�{�C��05��e%�� �\�%Iרz48B�I�c(@�ȋ~��Pi�㔣p� B��o�^��f���b�+��b��C��,9ej�j��+_%"BR�1p�C�3Z�ֈ9��0m��:�H3M��˓/=J̇��-O�����)e-ь�)"C�%��I0�F�%��̙cm��C�Il��ӷ��2���	v� *o,*B��������Q���h�fѴZB�%"�ޘ�R.#�bro͏�����9H8�n�۟\�	�)p�E���9�nek$�V�T��I������V��`�I��Lj���ƟP�'��N�zΠ� '�
1Ϝ�2�F7�ax2!Z�ː��X�CQp���~�pgN�P��rF	V3{ f����;8s<��O:�o���ء�+��s�$\�Sp��U`Sy2�i�R��)�=,�J�h������L19&JE����'MP�Q�m5��a���D�O���B R5$��"�&V�J�ã�'��I�L��u��ӟ�'��'K�$F�L*���]3�*M1Q�z0�	+.�A���;�l��9���p���M��)�@��.�)§m�ȵ��.�
J���U��j�I�'�����?K~j���h^�Q>6%(%	�9@�bI�K����?�	ӓ*�\Ĺ�Hϵ6�N�Q U-��D�9ڧHՎ��wȾ�p�C��>f�	����?��g�'P��F!�����B���<Y�'�(+�&k�|�ǃ�^KؔC�'&��@��Y�D����DK��MLM��'�T2@��9�V�kW�����@�'�,d21-�3< I��#~�r�'H\��H__t�R7қG��ܛ4�Ĳ�yB�'aH%Bg/��q�6����T/���A���x˚�Cw ����!o�`�2q���Mp�m��'p(���(c��Ш��~�q� �?�@�'��AB�'�(Dô�D<��0��'@�s&�1
W�49�A�7˔�N>�U�i	�'1���<�I�;q�6�c.�d��y��@R���\������	6$ $j�ݳ^� �)�-��f�,�� �I(�산 4^l��)W'.*���*0�"�flr��o�����?w`�*��-�FYJ�f�'M��, �����O:�u�'V2��XY�@%�JH"qO?��M���%���O���D�ilĺp�
>e�����۳�xR��O�u"���Y�.D�G�<ɼ�A�'��I6fך0�ڴ�?�����2��R,)�7�����(��kρ1��'#�Dh�:�p�%B�k��T>��O��̓�*K�.Q3T�ߍZ�����O��3�.��ڴy��A�@���}�El��aqЕz�b	NPx���M~�.Œ�?	��h�@�Ĝ�i����r��!��"J,B�	6b1,��4�ȡ	_����!r��?I���1D��`�@V�bc�z�j�-ZC�$l�ڟ��'Y6��pa�����Ox��<Ycl �����e��|y�"݌�F��"	�;�"QX5��&D q�*�>�I�o�	�$L@@h������9���E*H�2�a@sc,�6p�)��>�u���q�O�L�v��p��
�T�(L�bR�'{66��O�����O~b>˓�?�EG�*D�40fe�:d"�ec����8ړ�O̸)"o� p��x��3���{В�$oZ͟��I��M��������)��#�T@ce6ţs
7\�X=�4�	Ŧ���� �Ioyb^>�ϧ�^���%B�?i��c�,(]�0��A(�5������R�쁪V�����O���t�iY7��"B��<��D�W���D�RN��#���;R'l�6N��Ipޣ<��ݍY�
��b�("y�h;��O�UL9�I��	�4�?I,O��D�<A̟$�AU�͗��Rr��;qM�K!�|R�'� 2��̍1�4!���&{Z�����'��6M�O�b>���>){0�	/�(X�g���5'@��cb]�P�C�	�u��%f׎Xp���e���C�I-���ac�Yr�8����B�Y�&l�p��j��:0E�[R�B�I8
�Xy��U�;�z��'.�"�nB��;g�<T�ʹ�~a�f
�<�,�=I!U�O:Ԍ�P.��z�O��n���''�9��ҚE��@�EP�X���
�'��ty���	OS���f���M�
�'T�e@���G��!K�����4�
�'~D,J(/L�V+#a/\TX
�'v�H@`��`PE��?R�^�{�{��Dx��)�.���c'C�b�YҰ�ƓSTjC��%N�VH�3Μ�-�*�#�MD��.C�I�x|��`�U���E��>]�B�I�$n��ӷ�ˈe����`� >$B䉜3p�l�'+�%.�ΰj�@�� B�Ɏ,<�'�jh�őp�P&F>�o�T\��I&<�~��"�ŷ���%+�F�hB�*D}Иd���} �!�'jȖi�,B��v�ي��Y�X>~qK��E(�0C�ɲ��X��N�&n@ kH<,,C��
U�N�p��c�,������$�d
�$�6���`�K�(���*R�Ūe!򄇉v@ة�	M�o��I�V�M�{�!�����ʴ�[�ER�P�%[�ZB!�)pL}z5AQ�.�k�e�%!��RT/˗'����%_1E,!�� ;��K��C��Պ�$8�ў�P�/1�'i�PR3�����B��Vd����N��h#�c��M�le�q��\A��h�42�ԯ?�����jР�ȓu�Z�?PvN����479��@��x��8h!j��&`<QOẍ́�t���D��`����'*H�	 ^վ#<E���N��9�S@W�t�bEkuᕯ**!��+V�p�o�6�P�
ӡ��M	!��ؚ/j,�8 ��Z��XQ�V��Py�&�S�\@ё'��X�JiFؾ�ybI��S>)X�O�6I&��y�ə�]�����+�\UP݋������o��|"葬�"U��ŷ�eҤ����y
� ����,�nM��ʟ�v~h �"Oܝ�눢��£��t_:
�"O� ���4h,jO�DZ4|S"O�Cg�4�V�����cS�p2��'����'��AR��
�~Yj�a�L����'�4kr��q�Z�;�l�6Z�5@	�'���1I�'H�`�6m�T���B�'X$�$l�b�Y�#�Jr��#�'NF�ph~m��5+X]~�X
�'�`��엣G�}�ŅM=���ʉ��؉~gQ?=Hb,�d�J��"�A&d�,|xB)#D�ԣ+Y�rBi��!=3���@��!D�� u�V��@��2�da�W;D���W�6x۾���O�a��0+5D�xA5�ǄU���Bb���t��2D�܃�n�gl���ȑ�vU�0D��O���a�)����B�Ɓt��ѳ ��V��	�'=r�1�n�Вqy[v��#�F�<T�� H"�sw�H�mg�$�qO�A�<� �ep�T� 	Ѵ"�ZQ����{�<I5eН=�*���K�3���AK�z�<ٶ��
d�xh"e����"��OyR�W+�p>���WC�����^�l��z
d�<�!m�;Z~舡�Q�\,�"�^�<�v�0vo���f&[V΄�,O�<ɵ�;'�	)�
ƊV��h2S	�N�<��
�吠c� ��>d�B�Bx��Q筺����^�b��Ȓ�)^� ��!D�tr����O*4H	���m�Iæ� D�D�fl|_�Yk��� ��XR� =D��Q��4Pn���I��r�`ມ�/D��Ӫ֡@f���8�Z(���?D�L C�j��-�`gD=m0��k;��>mG��Y
�T��q[5Mj�zGHߖ�y��H4p�N�~<��c���y�@�O�n}2�B�,q��M�W�G�y��$"� �5"ޚ{U�1�B�(�yRĝ�6x��;U�G�x�>�@S	D��y�m\�}�B���_w���i�%ΐ�?! ��c��������Ŭi:6�� �Z�+�U��;D�\ÃF\G��<HD�9�؜�5�:D��B��^�r����KW*m@n�H"�7D�Ęu-Я����
Z/+�`A�g�4D���Ԯ o���i7�W�'�B��)4D�x���ۍnp��.
��"e�v�<9ƍE8���u��+
� 9k1�
*f�H��dg,D��6-�'Dv�4C΃�)"��C�.D�lZ�J 0�Q��_6F�L�PD-D���d�+N>d��蒱V�ȸ�N+D��@VgW�}]��9tH�\�l��F-)�O�3��OX	ad�8`�>�k�d��?����"O�j��.��!��c�/<r��"O��Q��4Bk��J�f�B�"O:����Σn��,�'I� �<%�r"O�,"�i��s"b!a@A�Rh�"O#p��A�r��r�2.^�xT�8<��~�$+T;J. ���)�~3܀���e�<��.қC�� ˳&����/�b�<����3���:��+G���[�$Rc�<�Ђ�2r,���4��le�W�<	T���&��6�W ]Ö��|�<Rl���P@�ϋ�@�P����@��*�S�Oʪl��oٜ$� ɜ�X[�4��"O�x��!�����)uX�SW����"O� ,I�d���Hsjȉt��8�"O�����ȇo�8�Qa��#6�ɑ"Oxh�e΅�a���	􊕙`��5"O8�X�"L-�����e��=��X����(�O"A��ÃN�0y�T�S�~l}��"O����U�;\A%�F<m��4Q�"O�9�`A�z���ǩG�D��"O�$Ȕ��K�RHh��z~D��"O�Y�ԫHW�|xU��΀�a��'1~��'�i��6^w�H8&�ֶ)��i!�'	�p#�E22V>�8�k'�����'��QG��O����ⅉ-��h)�' �<�nI�	a:YR`A6!X�j�'�N�1��r��ԯ����
�'�lL�t�B�k�^��ceF�"�҉��X�d�Q?�
rO�(�Q���α'����D$D��PB�&hL�zG�A9�>�2P� D�l�a���%��ISID@�B��?D� Jգ�9L�-i��)Ya�b8D���M��]���In��3��4D�L��%�>��z0O����O@��)�x^���^��X��荃�^U"�'�l��O�IYڐ{T�+Qެ�
�'Be��$��l�xȁ���?:�ܵ8	�'������N�BM<�X
�/���	�'����bN����h��H	<�}��'�y���ՂW�$ŘdD�6`|,H/O�$i��'���窎�"��k'��%,�}X�'?lt�B�'[G>�KbjT'�`��'c��)DNO�{N6AB���	�-��'�A	�˂�8�l��E���}!T�p�'�ܬ�W΃'�I����p ���������HE��
5�@�K�1h��ȓ��})��ѫ �B�h��L-q�����h��iծ"�X����E��y�ȓkߪ���#aB�Y�.^K�t��_�Y��D/[��H5��3;�E��DA���`H��Y��#-(�&�D{�쎯Ш��0B��M���X{���	�ňa"O��Ru��"�n�����,�>t�1"O��(��6=�(��Î���h�g"O\�w-ӱ-��{�b�"u���{�"O�͸u�2NhjUX��T�5��%�A"O�Y�%� V&"5K��߄$���'�'��������>��J��Z(,x(�S�f�4���ȓ=A���p�ʩN��T#�D	�i�ȓL쎁�2#�3.<�����YG���ȓ7�͋���ҨQ�NZ?588܅ȓ	i8�hg�S�&r�8A3��/b�D�ȓ��U��*X�#�X��#��S�`�'�p�
�>���+�뉂/������X5zd}��J>d�tϜ�S��H��R�U��4}h��`���0����Gʘv��T��rnd����U �p�q��0옅ȓn�����&��k:���eI#ȭ����r�6�ɲ(��Ɉ!��|�f ��R\���מX�̼��@�)=`�;��L�G@!���
��ٲê7�hPdeX�B7!�$�fJd���$8�:�i�c/f�!�_��E��j&;�aF�L�!�DK(I����̅�+>�BЁS�:ў+�%>�'W
��#B�B4 2�h#�ʆ?r�̈́ȓyun�* N^�)���rw"�ԄȓZmb���")��h�6!������S�? ��o�-6�%Z�͔+�X��"O$���F.©�FK�7&ۊmY$"O �aS��G�႖�{Ǝ�t�'��p���S�q��)t�O�a̜�y��Z��z���P����
 8(�y���ͩ���ȓ#ҒR!Ҟ1��i�@�nS�t��q) 5�ል�*��D���E��H�ȓ+�D4���'�8��Rk�-d�v���g�����3�T1HR���V��'1`�
�8�r����@e�bICS��"k��Q�ȓ��Aq6E�q`pQ��[.����i/�Y� �<l���R�י
|�ȓ;-2���'�k����Hx������j������4a[N�a��QAx�h�&��XqW*�G��m+b�ԡP����Ў=D�Ԉ7˄!09x�Ȥe�*|J�31�:D�$����	���C �A}*X1�e9D�$���/;|�Qү�k��d���2D�<*�{��a�9M� ;��5D��AnǴ����Gf�3a�2�4��yD��+����7��E��)I�y�k��P����tcʚ)ZlA*�.$�y�h
8�� �A/|ک�&E��yDY<l؂�kς!��t�&N��yҫ�}2��j�f-/2<�c�=�yѐj�(8a�S�Թ�J�?Qb������R!�Z�)�����"4�|r:D�أ��W3I���26	ɓ�|���4D���!Zd���,��>d>@ �3D� � J(�4�P�*�8o  �6L;D�ph!mu�6@� ��th<���/Mp���)L��C��yR�����O� �Ϩ����O��`��ԮF����ʊ5+l@ັ��<����?�cujFm\�;�qKG�n�y��O�2�I'F��mI�IBL*��@���}Ԁ�1Z/�ik�ꀐ��$����j"8z��0X|�!���R�&Gy�R��?����On �1����o1h�8��\pz �,O���d��d��") y4Tmr1Q�2q�}��<1�B�.Ǣ��D��5�D�[��\y/� #��'j�I{���'k�BͲK�U< ��	� PV�-��.(�XP��J��K��x�j�}���!^�
`��D�Cd�X����<a�)N9"�4 G�Ƽ	52Ё�E9h���c"8�JH�!�<W0օ��(��dF�I���$�O��S�V~�gO)"�� ��p��y0�`�>�y"R'5
� ���kji`����hO��F���э�tz�+�+ִ���ܱ_��'�R�+�����'���'5��O^��Y�H*-h�L 0W���$�Яs=\��G�}�J�&��j�Z���
+���D�4+G���`*�׺u��E	������A-;�ΥH M�@X��#�?%�Ɨ�ysh�6��I�i �qP�av�8�R��'������?����r��:���-d�$H�7KH���FL2D��	�鋊H���+Iغ�#�O@UGz�O�Q�|�ՈY�k���wa�u�\$WD��mY�;3	J�踤����H���?1�IΟLΧE6�\`S �8&��,��"�:���ĦG�k�PR1,�+D�I��4H�"?9��O�"�2���:��\j��`!a6)�h�N=j�A>���� 	f�ʽEx��_��?�%%Eq�P�0ð1*Z��� �?���:�hx��k�v@���>E�ȓCOHA��+N����c��U��'�7��O�ʓd�Չ��h��1�����&��(u#��� �i��	�?IńO�?����?Æ,`#$��@➆=����|����?`ܝ�d��Py�SPE�~�'gŹ�3$�L8�#�iK":y�钮�Ow�d��k����pQD��O���(��1]��㲨�/��D�c*ɪ!�˓�0?a�	�~{:��5D����elSx�<�*O��1ŋ
J���t��7B
^����4J���,����� !V.��9��`��P1�Ix%�-D���%V�E�d0H�ڕ�ne��$)D��9�JB�J�4Mrb հuI��<D�� >�xf�:���1%o��rl�M�"ORYR�»B}���-& ���"O�萱(�*Bt��#��r�����Q��O<�}����Bs,C��3ӡ�6�(ąȓp=���.��8�a�1
Ե}�Y�� ��!�ł�:XRL�īƭ;��0�ȓJo2(2�������$�#g����ȓ^���5��;_UB$`A�V���s����GQl���D�r���Ƀ3>p����&L����ō�:`����Ɣ26!�$�����c� +l� �c��?%!�Ď�*�M�D@[3����C뚈R!��?5)~P觌�K��%J3
�n!�D��'B��J&�p18 r�[џ�����M�I>"��=�|�[7`�{�p����X[~b�'�"�'R���aؕM���!I�����j#�����J5�=4�<؀�sz>�X��I�fƚ1��0i��x HK:.��M�ڀ�a��ŋ�Ѝ
��˃A�x��2�I-���d�O���Oh�S5���;�T�۾	a�A�r�P�D�Oh˓���	>?q���L��"� ���,3 ��c��|l���d�u싮Qo�E�f�[7�ʴb"�꟨�4�?Y���?�.O&�d�OX�5L�Չ�iMt�r(��)�(@���'+Q��F{� G
W����e�5d�V����D'��'���K<�g-�O:�'	���qE��i=��2�OW���d�'�z�	"�ӧ�9O�@����$I
Y�'p����t Pb��Op�,�&��OV,$?�H�E�<U�܈��ꅣ:v���5M���Ɋ�~��s�L��M�M�V�K�a(�`ABM�rn&�'t�';:q�J���>�B�`��!�8df_�mt�,�?Q�@�x���U��?9pK�$wҁB�M�bxr�q4gV��r�"}b�3}R*����ə�Mcs��#\�b|)t�Y��`���ĝcyR��9���ȟ�PA�v���f��* �����z?a5(I�T>�I4�����֟���'B�|��i`�:eo؍� �\{�u�޼�'���D�T
�B�B��GL	{O�1�p"��?9�L�����!?��y2��~��?J�(�a"D\��䙈Gヹ�?��m �O���f�J�pt �Ie)ʿ�Tcw"O� G��9_�Y;�A�31�x��xRP�0$��Sٟ,��9S>h��o��n�I���#��X�O��O8�=�OR�Aqo��CΨ��Ȁ�P�؍}�)�	��~l[ЄW�z.�z�_+!��ش���*�3����7�+\u!�Dc��� IX��h$��*�=!���yAb�1k��� Bgk�!�D9;\���(ʇU���goi�!��0�����B�ks��`&X�!��3n��p�P�R7Xtp� �i
!�$Q�'Ʋe
��K�9�:pz�
ʔ�!��/l)X5#�O�:m�=Є�ūE�!�$K
A2�V2I~�x{�"M$Vs!�dO�������@S
����O`!��Ao,U )Œ&A�pQr�
 %d�O,Q�$�J����	"]��y�E�KR�P� ,F�h1�1�!/���7DU6�W�Ly�a��C�t���"�M�DY24p$;��4(4)x=椨ԤA��o�D�NhUÀ�o���BD�O�& ^y��o�X!$������s���AG�u���Q��F�	 .���C/ �D��&��'Y�#<Yϓ 0�d3S �"O. �"��!�ȓJ�d�A�ʃqk�}��J� %�Q��Y�Q�rI�dn����B�\��@��<���a�N��S�.�����M#���ȓ �&�0k֦���C3���0�����_@Y���	�2܊$�	>j����	��sXn�
���d1��b���6�[�r��b��;�de�ȓ+��31�����6�t]$p��rX5S��|�$B#��*ʢ,�ȓ	leX*��f"u��S�"����@�2i]�=ҵ�4�ʹRFp��S�? R�)�D�."~��RfƘ�N@�D"O�0p���wK<3GG\Q�b� 6"Op �#Q�=��L8U�D�{��|��"Oܬ��V�4����Cx%`"Op���*zX>��B�%<ʼA�f"OQP���@��<;#���z���hD"OV]�C��$3���ϖ'�<ɪ�"O8x	%�Ւ9��T�%��P�v"O@���Ub��En�2X
��"O���a)V�C\����j�>CR]��"O������9���)�<\*�"O���wE��U���R�G�' ���"OhU��.J7?�F��򋝟uR"O���(�}�H���F�Np)JB"O��)gf�0L�yp���%�Z��@"OdY�t���+�)x��\	"O�m��D��l`|�k#h�.�Va T"O�@Ѝ�{e�0R"hؑI2�̀�"O�$���C�V�)�MP�2�R*6"O�ݲ.[��t��
>7�
�s�"O~��mX�r���WO��D��"O��QV�{� u��JعWmz�5"Op��^2s�J��J�RUjl�"O�!��� �"��sc˄Y����"Ov��%�C��||z�D޼;B 1X!"O��0X����# O<�A6"O��%�:x�!��eΐ\1�"O���R�B3�� fA0�E��"O�h����>���B�
��*����"O��#M�9,ԕ��)G'}� ��"O�лэU�gj���A	���"S"O2��ݧh�V #� �2o��Q"O�)�TK�]�$�O�-/�>�Xc"O���O08���z - �Iߠ)�"O!��0Y����Nk�B�r�"O�M*��Ӫ�jPY�#¤��E"O�t�mշ �r�8��+"����P"O�L��F�{%�=lc*��Q"O�%�.@z�����1{v]RT"O��!��0�b�ģ�,Z��"O�S���RԠA�FÃ�S4��8�"O������36
���"�<mмI�"O�	kUă.Q��TCS�Í��"O� "�F->�����/.g�~�iF"O�D���Q�a*v���ӛav��"O�ä���y�,
��?U��"O��.\�,���-@T kRkɅ�y����U�ܨ����h����y�DŁ HK��+jJ\Ј]��y�d�2��	xԇ�&�\0" �2�y�χ�k�`@��"R�'rN�@�9�y2GƫJ��ĉI����O���yrb�I�f���ӊ�v�	%C��ygE�td&\[BB��}�����y��}��E��*� � �bE���y�5Ѻ��ī|6���Q�yR��-��b�mtԞ��Ѭ��yb�A�\���D��r}�+� C�y�e�5�J)ЖAęc��yK��N+�y�� <XЅ�«U�DQʷ%��y�#��;\�ьȋGdm�G,���y2�W"<ـ��@�7L�p`�Z��y� R�"�I�'
=6��)�#��yb�$o��8�����3�Z�hf�4�y
� ���a�E!��#BE�2N˘�2"Or}��(V��^��ġ�'(��x0�"O��x�o�2��
�J��>�c�"O�ɡ�	��\Q�*� 	Ϛ��"O���N̈́`t^��lѰK�`�	""O��@V��hچ��b�F

 �v"O�̀��ݍ'�	��
m����"O֜hG�ЙT1P�1�B�?��Ȃ "Ov�cэF#A�j��t�K;\�Np�#"O�yqt��0F�2��_�K�����"O~4��+�i��u�0����H��"O�ȷ�T]I���q��l�]XG"O�(�#��|q>\{������"O��(Gg�cTt-a%N޴N�^ْ�"O̐:$O�P%��m�Uh&�b"O�`�T`�s���U�X){b8Y�"O(��E�W+(��L� PThQE"O��qB�I�>}j�˶�j;j���"O��A�(�w�Z�X��	R2��`�"Ov<����!X��=KGL��p0&`b"O��r*E#d/�����G,P�Yj�"OK#m�����C�?�^�"O>�$�H?аt���&�1
�"O�H&���t!(�b��S0%-;S"O����&��Q�ɣ#4���"OLApщ�����6��� �P"O�+��=JWF�1�e�	>Feڧ"O�4�4���?KP���?$郖"On�YUm���l�$b��d+6�s"O��3��Uv!y��H5�5(�"O�=4K�h�����!R�W����"O����#�3j��b��0j	;e"O Z4���D51��ƕ^cfm�"OZ2sn�pFD�:�O�CEJp�"O��{�n
�\��܊�gܭ]).��"O,�3�+�q��Arc��	u��A "O�4	 A)����!jņX����!"OjS$h�6A��K$i�6l�"}��"O m�nB:=�8h�P�h��$r�"OȘ�Ƨ��sy��P�փ>�L<s�"O�>;���bn(=�b�A�"O��`�CK�oH8�(c��k����*O����`ؿL��r E�T�[�'ֲYѐ���2l˂g�PڒQ�'�FQJ�)��䀡a���3/X��
�'fZqh��h�"�!�
(b�<�I
�'nd�Z�f�"�����ϰMK>͚	�'V�p��\(�t�ǌ³?VD�A�'�E!�֓X:
�@7�W7��`[
�'Ω��.U�u��Y��z��
�'���Q��/=�@���^�b�t���'W$� �dI�;�l8R!�0O���3�'w��eG!T�e�򍊗PFν�
�'f���f� AD��ѫ�H�F��'������\�%���H&ԁ�
�'�R0�L"FwV� ���r����'Ȗ�A�܂8�����lа���'ȶ�y"/�wġ2eˎ/4Z��'��[ATU�"�i%F�0��}
�'ܔi[a	E3+�"K��(�z��'� �j7`]�,�N �đ��z�;
�'���b���&��@0�� �$���'�8E E��l���J5D�	{���p�'��tf�K�3MF����lf}���� ����	���@q���3�(l2�"O(QIըW$r��8�D�	f��
`"O��A�іxI��� �<�\h��"O00Q�70A�}+�$N/(`Y�"O+d@�e�V!,��\q ��.�y2+@=b��!���""�
�b��yɜ8;��0��!������Z��yB`�뎤��E�K
�R(�0�y�l��Mo8Q["�D����a��yB@�#�D@��7x̠�搕�y�h6��$Z"�^�y���A�ņ3�yR@�(-p���Q�n�xqi'X�y�ؾ+��h�����3(N)�y�ܝBpf�j '�H�u����y��+Y�J�@��6"��b�Ά�y"ƌ�!&����9to�������yr`�D�ȓ4� �g#&�{A�G��y�I�_`݁�GAg,,<BBj�$�y� �#gY��I���X�"@wa�y釻J8T���%#��P���y2�ћf�.�*scM#<id@���y�� k�
��$\ANlz.��yb,O�.���D��UP2(�OC��y��
�p����� A3Q�����Ͷ�yB��n�T���!��5h�8b�]��y�$v}�s�� ����a��;�yr�^?*��55g^?����0�[��y��R�t?���d� �RXd �y�d߭K�T�g)9_��J6����y��6>#��b�G"u)��;����y¯\&G��	��)��$�U�Ǩ�>�y�D�5)��cҧ��r5ƌ�� �yC��dN�a��S�oN	���y"l7'&a� B��hh:�.��yr�N�@>�r��
&@�s$�F��y���9��,;�"H� ƨ�+� �y��@�OI�4�������u����y��:7�n�V�	┽�A�(�y���
��L���L��d	��y��Y@�qQi_�J�>`����y�F	:��c/�%U������8�y��ǆY%$����µO����%�y©��66x�k�D��������y��M:*/H�q� �F�����f	��yR�~*A���9�R`:��3�y�
W��H8�LΏ!p\v����yBF���h���z3T=�%�[�y"�Dh��𢠉q�0�T'��y�G�[�1H�V�d�"XCi+�y]5_�渑�	�f&L9ٔ#t!�$�q�x�WD��e��eqq�ڊBq!��j$��A��7ux8Ԉ�
��6f!�d/v�������,rR=R� F�'f!��G�$M���፹t�����ԜML!�_�w��z��Y ��94�z9!�'G7�Ո�*�F?hѤ.I8/!�6T��B�02'�]2�F2& qO�P'0T�������6J�8��|"�ֈQv9{'�A),�mh��yr���Ko*�y�� r�B����W��y��M�O���l�":o��U$B��yB$��>Qԑ:�E�&*T2x�Ȕ��y�h]�orhQ����R�\���!��y�
U�	�"L�B��T�*\��yb��- ��8خ
�fI��/��y
� ���6�I�)���c��ϙ}0RDJr"O�)�	�;��!��D^p��"Ol��瓣<� ua̵�J �"O�XQ�g@�hl
����y�L%��"O���b%�9qw$L��+�>� "O�����؇q���{��:8��"O����W�M��I�bG,d��K�"O�U[a�*6an����D8DP"�"O~��E*؄+>0��[Ve��!�"O���jV?x�՛���+
� ��"Oƙ3���E�>H�Ħ�<ǐ�!s"O����F
N�ԳC���1��s�"O�e8�jG�.|1�w+��n��$�4"O�Ջ5��=��ɞH�@d@Q"Oh8R�/ż`���7��.Z2��q"O��[E#L�@
ژ��_2��h��"O�h_b�8{���i9�"Ozܨň�)C��5�Ġ_�m	�hs�"O�D��/]�a��Qs�I%R�0}��"O���@��$�RF���@["O*	�,s4�����èi�½��"OL�"���,�p��0E[���+�"O��q�AP"����Q��,E�"OFˣjT��}c��Q�97e��"O�e�`��m�v�BT�̡(+$�kP"O꩘T��,y�PȔ8��5�"O� ��`��F�YC�׷q�t� "O�|�-�8���H��E� �:Mx�"Or<"Q(R�^�RmA��̄s8 ��"O�����ɑ�예 ��O��"O�d���7[�t[d	�:HA�1P""OrM�J�)V���$h����(˴"O̬g'�D � ���[s*��E"O��
e.lDj���ݒ[b� Br"Od����PԀ�����, E@�w"O���'� �u��胀
*����"O@�$D	-]"�B��A��.�"OTx9v,�:O�L���+G��"O��B��6Fl�P#�O��,���"Ox�ю�P�XՉ� �!P�yc�"O"�
����%-ӖH��T����	�y��N���Y6
X@�
=��̉�PyRHT� -<�3Sn�O��!p��e�<R��*a�=RC�ڙ?�Ʃ�b�J�<�w���.�T�����.�>�&&�D�<�$��T���qjP���Sg�I�<�k	J�����?�Ҭ��o�<i����LДcɾ�[�'�n�<�$���,�$	;�Y�'�S�<�flL�T\���� M�n��-To�<�E��d���×#ZԐB���l�<�r�%pPF��g-O��~����Us�<�S K&{�>��$ѓ;��ۢ�M�<������"�I����#�e�E�<�cN<
Kʽ�e��/B��D`�B�<����h�n�Ze-G� hT���y�<�kM�@�&�J3	�-�֦Np�<9��7w�n������ZW�ɑχc�<����,0�a0���hRpԲ�Kh�<�� O
��Pum ",���S���b�<I�%�"SX%���=a�����h�<��ԗ� 1�kŵ� �N�E�!��%95��j�(X�N]�����$�!���8%��A�dÕaun��t���!�� ��A��*8����J�U�"O�,H����r!L�ل{�s�"O0D3r��:�"�ó�E'���zc"O@�"��B�T�8e�'�ł���'"Oh �3*P�=Sl �bj��X�����"O����N�.�ts&�
<�H!"O�݂U���F��M2�(u0�T��"O:]���B	\��.ѨB�0�D"OƩ�1g�(ֈ��n��}��!z�"On�S�`_�q8��r '\�'����"O��S�s�"m��/�8�>8��"O��¢�H�}~��s��^R}��"Ox�p��M<&p�ؠ��ٕoB��Zd"OԹ�$iNJ�"Ҫ���E[�"O�J�J۔P0n��ǬY�T����$"O��x"
 � ĸҥIA�.�a1w"O�E�G�*u��XpH�7����"OX�H3h�nвI�O� �"f"O��h�K� E0�L�ٴTP�"O08��Z0��	r�@4Y�ܔ��"Ox�s/�B�.�!j�|�J� �"O�aP�Z$Hf	Aȋ�v�Kt"O|� ����M�`=�q�֝ ʆ��"ORq���ɭ0�F�ѓE�e$�TPv"O5B��!���fD8p�� �"ON0� O�N���.ǽ&4T� �"O��5@��~�X�
�D.�#�"Ol�P���6,3և�(,���C�"O`,����9G�sG�h����"O��`F��s�
���e�-���"O. Y� X;�����R,#�"O����3w���X��F�Y�xK"O��0"��[QN0;f�^
U��]�"O�)$��~x���D�ޚS$�T��'p��+7��W(�Q�H+6�^���'!(\"�a�V���㍴.$nU��'����D�
+R�� �g����y2�'��$j NT�����QA]m���[�'O�X
�KR�4b�9ڰS�69��@�'L��L[<"F�K���=f.��!�'Y�`:C�K�\��H�@W!Q�� �'�|����1�N�����FԈ1a�'Z��r�F�9��10g�U=58
�i�'���y�oO=)�.q���\�*���x�'�m���s��LP���*RBI�
�'�~C��4tJ}0�ܾ$��Y
�'�8�r�L�3$�T����>�D��'�np�[Yf:�"#��H\�R�'���b���:tĉ���B�8�>y�	�'m�2mR"s�(���bZ 2Ƙ��'�D!0+\�ځ����+��P�'��� i�?$�|����Y�� �	�'�\(
�O[���CʳW���z�':��u�#X`��3�� �	�'}��`g�00�����)�\l��'����e�O�7X(��/��&�<�K�'@#�$ѦZ$D�&�����p�<�PE�$h�|�@�ȚzZ&�5��H�<�ul@�_�Ƙ����*6l�R��G�<AAM<E�q�D&�$J�3�CW�<q�b[z.!B�uqd�˅h�<�iH����sA�;��h��˃l�<�A_�U窜Q�CFhJn�P�/�B�<�d�?q��=�&�P*&�^U�RhQ^�<� �,���'E%<P�FK�2�=1�"O1@��R�c���s��@ψ��&"Oj��e)T�QV*�2iȷN1�!�"Ot���h�^���
I�"#.��ST"Oh���O\!yD�! �"}��m�V"OLi��
�bF��!�:[��D��"O��(q�X'h�hl��l�2o�&��"O�Dh�ꕢ�0l8��"�.�p�"O@�:G�ڌ^gtq{G��aϺ�s"O���TƑgX<�J��V�_3n��g"O\�"v�A0k�f�����.���"O"�A�りTE���+	z´�2"ON�!�H\;l���B� ր���3w"O�1�bF��e�<�yQ瀣9����"O�p:`Έ%�pS�]���*�"OvA�F��L�r@��(��	8�"O4Y�ʖ�O�xѓ`0;���1"O�� ԍA��D�d<J�Nx�"Oz(�E��Z�P����J�r"O��墈�
��B��06��ڡ"O�(�մ�H�yF����,�"O����1��L� n��r}�8��"O�qx��[%���Y��(JA�=D��¡o�7�I�+B�Eh�<�#�0D�HZ懊.���Ǖ
=$��l=D�(y%�E�x��lU�F��U��?D�� @*��W��y!�$_�t�cN;D��z��6��h�����H�a�:D���!�0PQ�`O�Q�:��Ć4D�СP� �|]��)�k�B��%3D���E��@O��{��G�"��X��2D� k8tز1$đH��@�1D������)M���m',kڌ0��3D�|q�n�?!�蠢ҴD��2�'0D�T1&"K�'��\{��%\����1D���A�_*u�a�.O��m	��#D�@�E�~Bz�X�O�=��xѣ4D�X�����H1.f,�5n\�=蚌���Z����;V�f�R��=:�
D�ȓAX�|{�T�a]t��`(��4F���ȓm��9ɕ}0mj���F$B��ȓtAn|�e��v���SQ�U�¸�ȓ@��XQČD73�xHk��7I�Xl�ȓX4r�;�e	e���@1f.���v�,(W�ю&Y�x&o�05��ȓ��8zbH f�lD����(3�I�ȓl��h�MH!ft����*VF��ȓ\d��#D�y��ӓ+Z%�:(�ȓ}�t�D����}�a#�5/�A��3���9��9�: o)�4$�汄ȓv��؆jʖ"�����a���ȓay�Y�
_�{G�A@6�	)kf��ȓV "aԉW$��'�6�v��ȓb7�P�吹�� 蓪��]R�Ȅ�NV�� +E=���i�C�'q��q��d�e�K�]`��ې�ˠD��ć�_GLգ��
\��|��S�/���z֪e�`(�lhx�f/Ɨ&*��ȓW�^	j��2Z$��g�J�V81��P �A��aȏ;�� ���$��ȓs�la#��714�q�!
��d�=qԍ�v���a`1m>��S�I�v��,M
|6ܝ�rC��;��C䉡@�h�Srb� .U��W�N�s��C䉠{^��`���~>qH��MtU�C�)� D�A���&j<����H2E��"O�Y(�l�!�B4#U:m:�	s"OFHu'�X�zM pk�<0��@�"O�\��E�.tY*Yq��<[��Pc"O0e�l��|i�!�Ĉ�0=*�h�"O�"����셄�g��H��=^�!�d�r��ے���;�&U��&�s�!��Z>|
e�`.H�5�J�0�凩!�œ.0��쉺]�be�b$�fY!�d˾R�2��ӎ8?�V����>,o!�$
�)��T���U��-���	$ZU!��\
yi�M DQȥ���\�!��@�C�����MY�,!e�
��!��0�����l�F��#���{�!�ϪI$(d� mD�x�`q��K� �!�ĉ*�}B��>W\Y����0,�!�D��Hwň��%BZ\�d�i�!�?#@p��G��(Ḷ�#Z!�d_K��9d�E
^�lI��E8-�!���% �����L�fE)˽
�!�$� ���
w/o���[�x�!��05�2Ap�E1+�̂�Ոw!�DW�.��t���S�6ǲ���>a!�$��Ԩ�IueX(��U�
շd�!�$�z*��V��
�k�?GY�� �'���v
V�w|l1�&Csc��{�'A^<�4��x,1s���_EB@��'���ӭ��y ����: ����
�'4p��%$�5J� �UoN�t�8]k
�'��9��� ����+B��N 2�'��!!�Ð�慨�᎐y�``��'���L�60���C����'w�PC�M�,���eiU����'����G�^'1z@���N��*�'0F�QvEE�Op�9vF��-W�(��'�0T�6�G�"��E�ΦTr^��'!$�A�O��r�#àFƂ�y�'c:X*Q�%<���ɒ�˷@
�<��'���rO�{�V���kC4;��	�'�����ŋ�6��r�K�[�z��	�'�K�(+�Zyq��	�x�,�gQ�<aԀ�7	��$[��yG�PO�<1����	�� �;4z4���Mv�<�O.i���re*O�?N<�`�n�<)��G:
D5&=��9�Pl�<	W�̌_�d$����5�^�q�g�<qu't���!�	�O� l�f�	=�!�ZP]>�sA!Q(~20�c��!�$>x.�;�I�|h�=�s��cA!���3n��ʠ�MM 9iDT�j	!�$I/T���t'�a=XK ��!�D��1Q��R�mF�P� 9aQǜ}�!�$ٽx��������r�+��b�!���2d�D�&R��� �Z�!�$��@�e����w�a3�MT�d�!�31C��3�h�,�I��,�!�Ďy���pQ��;���t�Ѩ�!�Ą?B�h +b*T�X��D��!�Ě�j�<�����#�|��\	�!�	>X�(0j�	�*��q�`�=#c!�D� д1;������C.l7!�D=I�Rђ�׫I�[�CP�MT!��Ϩ/v�P�F�5if�y�f;!�D�/����R7��Q�NG�Z�!�� �1!W�0��j��߮`�~L�f"O��'IX4}��M(Ǧ���̡"O���r�Zy�h�҅��`�$(;�"O���&#5/�\���e6$E�#"O�`�t/��F��s�ɐO�~�H0"O��{��ٶN%@vd��К "O�T��	ɔw�X�"�B@��l��"Ov��0)�((~q��!So4AJ"OvP��)O�ಯ��8�X"O蠪�HS �����m�6t�����"O��6�Ӧ0�dm�VL�fvD"4"OVP�t�ƷN5�	���΍aO�x��"O�E�'g@
f�P�D	!	4b���"O���ƃ��n���B���7a` "O�X�mM`���iG�y
���"O00���/����b���/�1i#"O�ࠧaHPH*Pʆ#7����$"OT����<2����\3F�00"O��NK�7a��1H[���͹�"O�Q	�(P�WT D��[7>|��"OH�P�e\�n�*l��a^6h�pY�c"OP�`���VQ�<P�'{*�s�"ORI��(����R�e��Ȅ �"O�-xa���]!6�`�E�d�zl��"O�V̙"<D��$�w�4䲥"O��9%O�7���`J�"'�X�@"O��b��E+�nH	gh�ZaXf"O�֭�*,��#���`���0�"OJ(	R"�iL��SE˪6vq�$"O:�yf���H�)!���#DEbs"O�p"cWX_�$:�C��ޘ�"OJ�c� ԧc�����- �4-["Or8%��E\r-��	U����w"O^<�bX�^���
��E��"O�Й0�(�Kԍ$�v9�&��yr���j�r1�׀I�"`	&���y���6w9�6�@wN��	0�ybgל?#�xaCjV+l�D	���y�F�i(���	8g	DD���<�y�ɳ}�RI���u�������y��
	�Pl�w�B\&BɊ�	ܬ�yª
UR��E�S�
���$��y��̓(t�=��ā4�d�D�ޱ�y� �E`:�jT�('܌��O��y�Z�4��IB�l��H2C�N��y+݄]��� Ym�ک���Q���!�S�O
���o����K 'Մ͚�'��l��lM�0������h��m��'����ߵ��P�"C@�~�<i��ïS
t�x��E����~�<�烅$;����ŗ�U��2wo�E�<A1,#q�RE�e�؁t�شJ�MN~�<�5�G�en@;q+�>	9X!�m}�<�C��(i�qWo�7u�u�R	Vz�<q�o�1L:����˵H���A�t�<YQ�۳e7��D	_1{yF �@ m�<��!�"#6Q�G׈(��M�ao�i�<�l�t�.ɠo߆d�(`�d�Nz�<���
��&��Kn�跉�}�<��/TOnQ"T�q��BBR#�!�$�@K�ak�˓�]�ȱ�@̰T�!��2_9^ ;a�F<h[LЉ���'>�"��L�+ɲ1��囱a��p)�'E��y2�D�.2�(���Q%3�P���� 4��H��}��{R!>��l�V"O�-�P�D�[u��C1b*���{�"O�1�M�v� т�g�+;�� �V"O$	 ��aڂ����=Ђ B�"O�Ģ�
".�8m+����)�b\��"O@�Ԧ���E�+ݭzD�@�"O�ݡ5K�<E�P����2:qa7"O�`�u+�(����u	X�f�Ա�"O�A�ՄU@��(]���S�"O���S�D�F�9b�'��Z�*E"O��)���&~��bB�� �T�#2"O̴�j��241Jq恷<�0И"O�)�@@�>��@����@�\)c�"O�� �O�{�p���c�z��j4"O���&�4LmӆB�*8j�i��"Or����݃"�P����gĨ@!"O^����o�0�e�Yv�����"O�e`��-fWb%1G/�7_��"T"Ot��%*��qS�9�#�Id� R�"OR��H�8�8�a���M�f���"O�	��)#��\���|�|"d"O���B�,a�x��؁,��u�"Oa:wL�Ȑ����Ĵ�.�y���d�T�oH��#�y��\~D����*b�:ĭ#�y��E�z5v@��MW���WkA �y�	Φ�؉yQo��}�$�foS=�y�]�&E���� �@s$����y���u���"��}��I�)���y玄H0�Zv�Y-�|�3�yrc�'j781xEI׺b���H N�y��X�9+4�欝.a<
d��٣�y�����l1!�T�] B٩��[��y���kB�x�1��!`,��L���yR�c  �cT苠����y�G�25��s�I� ���4�H��y�(��<���{�Gճ���0b����y�_�}_ح�q�� ��L�К�y,�6|�Xz��R�x �����J��y�۲J;��[��]�^�Q�i��y�o�O��D�S�C7u;L�0�y��U�������;qBx��Ś*�y2+N��u��n��I�Ԁ�PybG ���Ɛ+'���5&�\�<���
O��
� ��7Z�lH�JU�<q2o�?9�`�" "5�d�Q��N�<)�&	�)랔���ܹ:�a�`Ht�<飡�/4����6jI%��n�<1�C~|���1tn�Q)Td�<�!�T nE��!ѻP��t��T�<Q�F�t�8������d�5�f�<)7�B��&FazR ���v�<��E�A�����=F�4h���x�<�u�d0�g���-^'^�C�I����f@;$D�M��b�>C�I�qy����H%�m���Oz��C�I���@�G?�����xC�ɶt��di��[�c�P�Z2oã �ZC�ɐ{�QÊӚ5b����B�@[rC�I���h����t��3�A+U^,C�	(-V�[P�6��͡�d��VVC�I�l\:���E=5�����1.G2C�I?V���Ɓ~D>�0�E�X�C�	�j۬|x#aN�M\2!��o	,� C�)� ��s�a=Dh��H3W�(�"O�T"Ĉ$�21j�<H;V�r�"O���c/�<�l��"i�48��"OPQ W+�%xSHY�⊋<A��� "OnȐ�(O2FL���cڋC����u"O hC��OGZ�=B���p��)"O��I�L3h���P��Y�[�{E"Ox�;p�ѣ
��4&,��&N�b"O�(c@��*2:Q)��ƿ|�qɇ"Ot��/[ }_~"�)�3=��qZ"O��K��)�([�Mq����"O�D���$38�`�'6�j��S"O���5�Q'H�h��5�]�5h>-K"O�Hc��>nZ��ʳ�X�g"�3"OLP��)WII��,[�,[{"O~L���_�,u�A��]B��s"O�%�fFD�J��h��a�'K��@A"O�1���jzhM�����T��"O��G�Mo|�ya�*C�J��i�"OB�{�LX���:4�����[�"O ����L/$tE���t���(�"O�@r�D�.��І͌�;k�I�""O���W
��!~)[�[<RS���"O���K#W�, ��	�a5�pj"O-����>T���t)�$\"����"O8����˩V,* Ѝ�yA$� �"O���i@-{��D��+	�8D�Pzv"O��Ɗ�c������]3t@xK"O,Zrn�\���$� z?H�Z�"O�ۣ�ː"���$�G53�2 B%"O�}�v�D/h�+��ߠ3.;!"O�R��MlP�f�!>�m�e"O8� q��)���8p��(Q�؈q�"O�����.3GP0���`����"O�a!�	:5ܰ�PᑻZ�t"OB�)t�vbƜ�B@Ѥ���j2"O�� "�1�H�e��Z{�i�"OԀ2���m���y���"O�Z�NA�2�$�x��Ͼ=&d �"Oh9Bc��m.؈�'Gu@|!p3"O�(�Iw�Hi���a*p(��A6D�kC�Ժd6�#�Ή	^��Ł�'D�4�Gk�'����B�<���2D��q��׌uv� �'ϔ.�M�3D���2 �[��������
1D�C�%�,ZP{�E�z!�`Q�,D�ԪP�O�2��3AL�!�X9��+D���˗�W�`!���H�B��@�+D�$	�/ơa�аRug�'�t�Q(D����>/�� ��`xh�l0D� �G@Lg�� r^�x��1Ao1D�����Y���Z�!lr��p�/D���R#J�?*|dHv
� C2� �B/D�D��E�7�P �e�4j��u:�+/D���S�K5W�4�ZR�� ���6�(D�Q���f_n�e/~F%��h&D����ޣmz�5 ��� �Ҙq1I:D���i[�)y��$E_�K��X
!<D��8 �L>�~�3V Hf�|��#'D���æ��:v�[�!ƄswD�6%T�:�#ܔO�E9Ң���� �"Oʤ��%��&jXpR'P*�8IKc"O<=��/Z�B8�H���S�&uB ӧ"O�8��%k��)&$D�xX4Q0"O� � څ"�\�����ᆺٞ0s�"O���b��(��w�0f�e��"OtIBf�RVH�P&��OO��"O6!9�ObIF@[���B⦁�y�Ⱥ��Xid��>H��0�A�]��y���T�����
�n�6|�� ��yr��!3W��j��Z�]����yb鋮uX��j�BZ�g6!�P��+�y�K�Yu�5QU�A�s���0 
��y��I�.|���E�D4c��A�E2�y2��41x����̸\�z�S�'�y�怭0�~��g���AHN�1����y"��7i��ITlڅ:�`��3$���yr,�n�l{�&�4ڪa����y�Ā
(��9ya�P�0�9�u�'�y�ۗ:��;F�V�3 (P�+E:�y�Y���RnY�*fl����y�V?')
A���@�D\Q��I���yR -b�X��K;�JUX K�y�+�MO��jr���$�/��y��;g��8���J�MP��F*�yҧ�RۄAY�G-H����+�/�yB���:=���q��8�Ń��y�耀>�1�'LǠpe��hX�y�$@|�sFh��ѓA��yg�`���ZKJ]O�����y�i�4D*:u��)�"M�v�j���7�y�E�)<�TmbNܵ.ɾ4���5�yr 5Π�q�nJ�#��Q�Py"a3�N�i�#�mn� ��J�<GI�* 5�y��F�p�����C�<1�U�����'�H�aʕw�<�e���}M�����A$Pʑ��Cq�<Q��ץ^�L5�'a�<���l�<Ѵ�G�K���Z��N�s�2�cgc�<I�G�p�d���.=N�#��t�<)t�	?PL ���(�<`�D�Es�<Y�E@�x�^	�UKҌ�`�B��E�<�S�J	B��Cg�
6��	����B�<1��P���"d+nt2a�]|�<��I���؈�Oۦ:���A�|�<�� W\���#Ǌסg����E��v�<aÁT�0z�� P
q�81Ӥq�<1�dF
|p��p*Ŕq�n,Y�a�w�<Q�)��(t�WeO�jw�)�g�\�<�t,�
p|҉���D�4Z�U��Z�<��C
�tl���ě9	`���QW�<9�&%Qm��Xn�x���S�<)�)�6j&�*���zP����N�<	��R� H��ӫpA�uXeęS�<���4a�ebE%	���ˆ�Q�<�#��*) �k�g^&=����.�F�<u� �Qp���c� S�:���C@�<���ru�yY�Ƒ�@�K�&u�C�	 6�k�L����i�C�O�C䉔q���!�Fͭa7�,�OދHC�I�uV���˲hd��
H<>�,C�
|�A��Tpb��Eż�@C���!�G�>q f�(�p�jB�	�R�`dBC�	�O�nX��.�v˜C�<�n)*S.3-���	@��^?PB�I3=uR���E��hn:����S��C䉨$��Y�4@X�� z�"G2B�|�.%�C�C&l���Z��N���C�)� �䢓EQ?���26gM�HH�� "O���dƆ|_�y�Te
;_1n|!q"O�WK/q��Ǝp�l QJr�<)��:t�c��L�.�D$�DD�<�Ս�;	�~,R�Ɲ	k��K�g�[�<q�Oٲ3�$HI�!BD;����<7$�)*��-��Y�+�<�2�KA�<!��Z$*�k�>l�b�9P,R@�<�MA�~n;s�f|B�C�IWx�<!�G)+a������1AѶU�K�t�<����z�Le� .)qU^�2��Cu�<�a˓ 
j���`m����_{�<�c�27�P�����0s���BI�q�<�Q���J[,��aŝ�uΖ�[��l�<�6�L��,m0w��X�VYyF�~�<9$KAO jPhPoЦ��Dq�P�<9ݼ1��c�� Y<�ts�#C�<9�hӹF�����&HN�)&��u�<�3k�R#���ߟv��M{#B@g�<��O�eB����]&aYT�RU��f�<���(}F�r��C&	�8`���z�<IS��08&tb�e�EM��ɧCN`�<q�m��Yk��z��@}��8JU�_�<�+��6r��"�T�����]�<q���#�'��3�<�T�HW�<Qf�R�@}X���nF�@൐�`MU�<��I�;G�� �J3a��P��H�f�<	��=1]LԠpׯU�,p罞!�䕫P��hC(ٜ%��ɰ��)�!�D�W=��R�@_�QT��XU�)�!�dG��¦������Q�	�!�_�|P\�BD�C���@�)ʲ)�!��^8�i!@ f΁"¥	c!�$
�� �A�ŏlX�Yp��,#!���0=`���&͝;S.m�Dd��I!�� k���kP�"�r����>.�!�$V
ž��dn0>\���!�)V�!�D�,)�hHT�Ϧd@��jbY R�!�t�~H�c+��2v�jf��}�!��A�T��)U�B�*��9H�����!��Y"Kt�ר�+u����ϙ�yn��$��<s���=DpZӆ-]:�y2��^8�u��W?%���q�]��y�
-��r���"v*$h��ɛ�y2Ň�|�RL $����� Y��yBm��8p襑sl��h�����I�y�g[<���Sk�>deh��B��y2OH�X�: �U��%[���(�y�Ʌ��t�۲)�*Z��0;�#Ʊ�y��O1I �IơFM1� ��߯�yB��<����$�Da����y�T=��y{�Ǘ�D�BF��y"�5 ����� 	t��83�I��yb�� �N�.��	����"�ڳ�y��+����c�$q>~z��X9�y#N�]zQB*jC$��'
7�y'O.
�#�
�c�=��	7�y�2�t����X��wg���y"���	,@uR���N�HL�qE]!�y"��~v�� f�R�oh(	�h�$�y�o�u��H'
2� �	�'�0�y�@�o���K��0yb��(B%ަ�y��X4J��d픤({�!1�K�y" K�dy��seҞU�n-ÓO!�y
� lQ��݊�ʨ�v�֠@��m�"O������'�P%�%DD�o!����"O�Ź�8MG�$��"V;<@�"Of�r�䒫�l�e��G;0ɑ"O~Pj�%iwP��@��(� ��I��P]����i����AsV�Ұ.�<`y1�[>������O�h[����S�huiŤG@`˳� >���JJ"���0g-JFײ!:sD��HOdk&�X�L>$�'9Y��9H����T:��G��G���*W�3X�4A�%AޤK��̓ti�O��$������F�oN�i�Z����b���4+0A���!�i>�$���'���xV�Q�0�zN��I8�@�Û&/fӠ6�	�U�|��-Y�t�d ��FS�P`ݴ'���"3R�ܖ'���O�'�'���z21iC�\>EB�ʁ�ɑGC�ć�&VM�3�X6,�J�i���Ͽ{��Ko���$�L�;����l�ʦ�E� C�����x������w~A�t@�4{�1�k�L�dK�(ɢ̈*%� 1 �	s��L	��?A��in6��O�#~n�-
G�eQ�������#��| ��ß��'ayb����ȴ��[?�	�%E�HO�7���'�(�O.�rhQ�F2��*E�ʘ]�HQr'A�<�Co�7(k�v�'̈�{C���@�*S��@K� �D �(0	P����X�F�2k̊��ψ�O ti�i������;,ޖt��N_�� 0P�+KLV��q�D�!���ڦ���g�ɽg������7a~���T>s��k�(+
!H�aݛfI�t�,O��ķ>1g��v���To���%��A�h�<!�  2DÔ�^�~�Ǡ�,#�� ��a���oZ_�	�����<A�����0Q)��?��BcωG#���E�_���<I�GpDX�� �h�)J<1�|��CÛ#�  `pN�C�H: ꋝ[R�"?�%&��Aʖ�#D �d�Xxap��;M�m�c��3r�~�A�,I<gd��ѦF�Fx�!�?�۴Px0�#�����Y�T�X8�jPlD��͟\�	[�IF�S1�~��P�I�A����$G���IE؟Ԓ,A�.T��[Æ�*,a��r�A��?�Ҵi���'B7-B��mZ�t���[b�Q
i�t�5���q��a��B�B��?y���
�L���:c>�Tb�)�#%�擩X:����,R7H<��EOr!�#=hX�{�
�FR2/JV��s����u�'��-�U��.-Ԁ�b�se��	!l]p�d�O���	E�����T��V%S�	�d�7�H�eά�D6�i>�Fzr�8��Q�ʕ_ �8W����p>y��i��7�wӆH�ьW�O��6�F�D�����Oi�7����	Qyʟ�O%Q�&��M���4d>�5aTk4 ��caH9j�����P
q���x����W蔻Mv6y@�E�o� ��k���M3�O�=�tH�c��OC��{S���@��̻��e�����X�Uƌ@��H	�f��x��˦;���ON��_y�����V��?�8�I��+Md8����~"�'�azR�O`{�䎖%Wj'<):Ф�M�Q�4*�4(���|��O���ʿYP�t��Z3vJ�(�LT� ��4'��퉏e~p   �   9   Ĵ���	��Z�:tID:,���3��H��R�
O�ظ2�x�I[#��C�4e��B��.�=H�n�,��x�$�#f?V6͂���H�4;p�1��\�I�$U
E9�`[*P��2A
��l�tD�UE/�7�T#<)�&i�Z%��MX�J���$[���DX���'e �jm�,6?i��K) ��6Mp}"��t�Lc��&q�N�3�jAg� ��
ry�.�OB�6d����9On��$J�)Q����Qa�dL"D�#
(6 ̋v�H���D�==�������'���D$�q��Ȫ�`����H(��%����3##�'(����Ð�> ub$��T�M��'��Exr`X^�'��E.��!���Y�P����(N.#<���>ѧ*�4e@>a����Ty�F.r��)�O�ڊ{@�Y�V-;��ΠZ�<K��F�Ms3�-}n�"<��/�G�ld"sf�|e�Z0�E9Z�p�>�Vn)�n�4�t�xEY�(۵#H��U%��0�� �'(��Fxbn��nfR�� 7{x��K��Y�0վ�a�:$"2#<���Ox�$��q�E���6[�ٱ���OB�8I<Yf�;t5���Q�I^��p��ZS?Q8�\�OR�I0K��p�"�Q�Љ�ޢ4�.���h~r��97�]��4*��ɏ1qࡉ��OT�qakHn��SӨ��
,MɁ���H��܄N�Q�����>%f߷&.T���	 ���3ǄI}R��j�'ѪGxr�H�s�NS;2F�� �%�y�n�J�  �O���Q��U"�GUy�Ne�
�OȔi�)��8�L�)�A�2�"�����Y��M�@����nD
V������)��3� ��w�?.��E�d���V�>ŉ&͚0�?A��:���<�'�?���?9 '�!1r`hlA:���`�O6�?i���ċ�	����۟ ��̟P�O� ��F���ӈ���t}��OJ��']p7����O<�O76��U��v�>e"i�%cLY�c�aA��4��(�� �̒O����>A�#��19�B)(3��OX���O����O1��ʓY��O�=�0��E�F�;!&��em)C���*�_�H��4��'-&��M� �z!��C�	����yZ����a��od��Y�a�|Ӿ�|#�틆I����O�Zc���p��@x�`�:By
�h�'~�Iß����	����IV���3e�4�I�#���@�syB6-ջZ!    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �   C   Ĵ���	��Z�Zviʗ&���3��H�I�
O�ظ2�x�I[#�<��4d�v�V��$�s�ի-h�K�GЃi^7-ƦR�4WU��!��U��) ��|�t�G�,�B�Bc"�3���uH4�,��"<�hӐ ��g�
8��b2�Yo�p��X�`���gxN�Ѣ�*?�W L0
7m
P}R,l��)s�R�9��\�S#Y%B���k\6��aqB�X�i�JC�x�+��,�k�
�tj���@-Y�x�eӋ��F�� �'��5�����'r�[%C�^:�nڠ"S��PM�p�Z�Y�ǁO�(�O�����$����u+��
��$ӬqU��-�Pp��"<���>�]B-�S%ۻ[/�,���К�M��I�)�����Z��20���3j{AM�3�8�� K4}��e�'���=�LB[|��L�-,��A' �⦵��I����!m��o7����R�ԅ1�Q�1b�0y$�	7&p���m�j����ؿW��@�GJL�T��˓��"<)� �	�f�z���@<i 4���	��i��ɮ52���E�'��Г'&թ]
9r�ږ!����yRi�'�J�$�T�7;%f�;�j��T]�aX�����2S�ɄZ��'�f�ɱ0�\P�+x��f��O6���~~B5xt�l��4��	S4�x2�O�T0B��@<L֘aI�ߧp�ڑ��Y�T������c�X��Q� `�'ApE� \E/�|� ��[�X��O�)���䃼�OHt�c`A�M�����E	'Ӕ�S�'�@ �����d�5�?�!\���ɬ��ˣ��&�F%�P�l�L�������/Q�
�B�{yԠ��ĳ?��'�de����;;ب8@�J4�|��'�I� �I�������0��w�4��e����倗>�Bh��J-
6��B����O��$)���O�]mz�IBɆF�
�{��̧L���Ċ�����z�)�S)G����b�$��ԜTDi�G�x��@���h��IE�В��$+�ĩ<����?!��1-����� E9D�	�7���?��?A����$���2U�C۟��	�hh2��^��p��0c�*a�n�D��3P�	ޟ��	p�)� (���̔�4Bx����$�5�g�����ƤXw�QbV�W� Xs���O �(wNҊr_�AQ�٤�r�t��O����O���O��}���<�F�@�kͫn'�J��3p�y�����֠Q    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �   F   Ĵ���	��Z �t��8-���3��H��R�
O�ظ2�x�I[#��q�4�?iU/�+SM�	�pMW�0�h<@P�\���j�6Xoک�yb�$6��[EBhR e���B!N�v�9R��Gu�p�i�vu�o�/�z)���&pF��'�DA�.I�$�*O0|B�99#61X��9��ϥ�̘2���5f̴ �PBP<Z@_�L͓Ooք��Jʻ�ē%ha0P8y�l�3��y�D|�4�%^�態wH�<)�k�����&�����nu���_��YX!�+)
�˲%S�?4`g�5��L�OH��O>	�/�o��z�&Qg@�:�V�<J!i �"<q4m�fWd�G�Nz�<�#�����̻��I�y��əR����5e�9J��,Ӑ-�ۄ�'k0Fx�a�Y�)��	0&Q	t�3(_�,lnڭ:��X���I6kH)2�����FG	��Ȥ���/�I2� K����P�L�L�XɆKǺ2��5`%��<�e�$�R�4KԄ��_��lb�l��P�������D���a�	%}��G�9wH|�,I^�ܬ������'%�PGx2�Dd≋wD�{�Ȗ|.5�q��	�EI��D�xrn��� CIJ�G�n����N=��(��o�O��'De�aߌ�M����9��Ҕ~+�ŉ�}��Fi�F�Ƀ���.�剄��I�1��L>���'�xb��<=�`/ݤ3*�������N��O��1�����
@o��d�x���R/!�$��#� �  ��O����<�O��c �ۜ^Fe�0��b��Pa�zӮ��g.�S�1O>�	�n,�E�Ր
thaäj�!pt��Pٴ�?���y�FGh)�O����PR��T��ŃKզ�Y�&I!lO�$�OB�dv<��s�CW�X�"z��O$H���o���`I\�ē�?������f	<#9�gcH�F���AQe�o}��U"��'v��'t^�LRC�){��U�Vn8�eA�Z�(�J<Y��?�N>Q���?�ebD�&�z����B6���
r�z��<���?����?)�O�ܠ0�Oތ��FƋKL�PQ.J*#��ݴ�?i���?�M>a��?At�J�C]B�l��Z'b�ru'[�f@R��/��|ꓥ?���?/On@B��J�D�'+bU��Oތ�8��.L�HD[RdӢ���O0�H��7�I��������`J 3��b�h6��Op�d�O�����D�O���rG^i��	�C� 9��;��LN�'sb�'	���b��ʘ���ͣS��Ԛ�lT��!0$ &#�f�'��g�/=��'�r�'���'yZcn�93p��+7����Š
I�dߴ�?��4����Vj�S�g�? �HD�P2զ�)�,X�3��a�i.Jls�zӴ�D�ON�����T'��/z��e"��
8�>��b�3d��(�4'$)[���Ϙ'pb��Q�
�#�ݏFmʉ#F�N-Za�6M�O����Oh%`Bk�<�.���d�����`R�hM27�۠a~8���2��'�حb�	.�i�Ov��OLR)F��`�J�4{����ئ����S�R)�N<����?�N>��~�Z��M�z������Q�c��\�'"���y��'��'��I�����OI-r��(�Tnν]XX+��ē�?	����?��*<>�IT.Y^�h�T�P��Ȑ����I̓�?a���?�-O�yRB��|�e��9��x�g�J�{]\��du�I͟�$�`�	͟�hp �>Q0��6�����P�=x(@��b�r}��'�B�'z��|�b��L|�s%�1c*�ɉgvNAPէW՛v�'u�'b�'".�s�}B�>�!Qr�N( X�$@V�A��M����?-O2훐aYM����(��3aMǋUTn�����D�)J<���?	��S�'e�i��a��)��K�C�*pCfEZ�d˛&\�| !���MC�\?E���?��OQ� Ą�?���ۥ
}��ib�'F ���I�E�������ø��q�<Q��&��0"�6��O~�d�OT�I�[�e�
�AO!-��Dk�*��(þi�Q��d$�Sɟ����(&EpKG`اI��Y3��N��M���?��7���&���O�����p�I)5����t��W��c���BK?��������r��ҳM��Ha��M�)@�ՃqDE��Ms�]o�� U���'�bP���i���G�-l�����h��/H��Ia�����t�Ġ<��?�����$^*1�L���"[�Pɰ�m��9�0 B�_}2Z���ISy"�'�R�'�� �H"a�@�B��^=�uȅJ?���?9���?����V���l�'z�6���N�4�^�У��$V�&5ldy��'��I����ӟ�B�v�d���`*�b���l�Y;�*¥����O����O,�Gw^=xER?y�I���	�
�.�*� \譢�M��M����D�O��D�O�$Q�?O^�D��x�dM��2��
�&,'�5�lt���$�O��=��a�P?����H��1W6 ;MJT)v��>+�p"�Ox���O*��ʃFD��'��?�"��T0t����3��yh��S)g�2�1��+�i��'���O]�Ӻ3�#h$L:�I��δ�!�ɦ���ğ��u�q� ��Zy�I�381 �th�J�~t M�.`�m� ]7��O�$�OR���a}2P� �!���h��*��C%U��u�ڑ�M��<�����$-�Sߟ(���H�!dȟ�P�x�hʙ�M{���?��f�=�wP�ؕ'�R�O�I��*�55��2�*�%�@�i4P�P0&n��'�?����?��
#)
ܕ�����JܝH�6�'�hBo�>�,O���<����Q���Tx�gE�r�AI�x}�E��y_���	ߟ�%?�B��>UKpS��K�:�JH@�ꐃ^��	H�O�˓�?�(O��d�O���K�>m9	¿��p!�R3p��z�<O&�D�O2�D�O��D"��a���x�®B�3�$�(&�7rQ�J�e��M���?���䓕?�-O-���iL��P����o8�!
�4��L
�O���O4�D�<�aiF�C����Ps��T1��2���7�V0X'���M#��?q���';qO��(!�&��]��U)�ZLX��i�2�'|r�'ª��q\>�'��T-�7
���D��#㤕 5�P�.O��D�<!��Ko��u�+��A�5#b�ܰ*Vnύ�M����?Ap����?��?������?��/F����^UZ�q��(.#�o����I�"U�#<q��4k3pUqF!L_��H��S��?����,��s���0=	�2�Fm3��V�"���[�<��`�5?���ԭ
�.3Y��[�0k�	S� L
Aɂ�J���.I�թre�?+9�t�U��2t�2Q^�$C�����U01�`)��DV=��՘&�>LpU�����ZLuq��X�2P@�P:%�0��a'Q!ܠ5X�� *d �#���[4:��g���Px6�Ĕnv��k�
�?���?i��Z��.�O��D|>��A(V�S[��	ďRI��\���N�8C�	I���P��͘�-A�k>����D���N�� �D�e0�� ��ph�/T�.NH@���Φ�#��9-$!4�E���@J<y6hFW�¨넅R0��[2�G7J�(H�	��TE{2���M��A�14Ԕ���bM/'!�֟pt�-;���<<���Ȅ�p1O4!�'��	D=�aB�O �]�2mb�0��+l�$1�V5^`�$�O( qi�OH�z>�I���9'�ڝ03�خ�~��'�2�Ѣ�"o^ � "O�p<I&��}��� ��K��Ӆ!/�k׃�}�����a5H �x��]��?�����d�am l��/�;M��&T�	�1O���DR�
n��0��F/�r���9�!���!۲�
Q Р�0k��~a"��̔'�~����>�����	��U����Q�KG�-�샞q�ƼP d��X<���O�`��)d�AI��ͅ0�?�O*�S�4mj��#��#�!��o��G��'�
7	Ҋ8�i��  7A�>)����'`�n���՟5H��d�)}b���?���h���� ���R �\x��נJ�<(�G"O�9rǃ(l%�1�դ�,��P�'�#=i��Ɉ!�Ȁb��x�0/��W�����@�I<M��T*aŎ����	韄�i��F�c�N=b-���@E�_t$�A�^�L���@�b>�O6�@��*2�$�E�a��e��tc�+�O6��Ɇ�и��a�H)���D�A�,Igɣr�������$ʒG��O�ў8���?np�⠅�l�ZCe=D�7e��(�jm#D$�.��kpM??!��)
/O&! #�ǰT��<�1�D�9.8��K\>����	�Oh��O��D�к���?��Oz�Iᇏہ;Zd���̆�]�D� ����x�k�&ɠ�x�E�)8������*F��@	�'Ψ��vC�3H��Dާ���@��!�?��o1t}B�N^M8��r��	o��)�ȓc��TKQ��p��(���X�dS�`�<I@�DP��l��t�I2Y=L)z�J֓x`>�kƪ	#"z`���<�`����	�|Bq�����'����^��YK�O��1��$O��� �Ĉ3m���0e*T~�1���Y:�x�C���?�N>��X�C��t�!��?D�����J�<���O'	���
�o�\�z\@b*�_<y�i�x<YӣI�_X8!B�P�"�,[�yB��&�듓?A+�������O�����0-q��;1�[I�=1�	�O,�d�*$W"����S
#�:\:�f��$UJ�O���*���Ɉ}�.��v��;F,�'����+[@x����٘*�>�PBI?�/2�X  ���U ,�LG�<kD�'�F0p���?1����OJy8$�D)7��$�p���F}����"O$�ڷfܫy��E�D䄽d2	S��'�"=��ɝ"i�)S����>\�V�M�.���'��'�H��)N�'K���y��N���8�cd�+ag �*�C7.1O�%K��'�(d`d&�/&�v!�eGZ�xM�{�� ���<����;&�p��)�="6�P� �.��'1�P��S�g�nM6T+&ܠD�!�kֵhC�I�9r@���F7w�Q:�+L���ߑ�"|"u�T�Rr*�c�I��u��c���72�+@��5�I��p�	ݟ��_w�r�'��	:*��:V&�#����1Ό@!����Onu[�/�B�6�{t�~���e�NM���'~$�G�֨E����#��Q�� �r�@�?1�Z΍�wE�C
z�3��D��ȓ`ߤ���v�9��ZB
"�I���'t�ŋ�m���O�<��	�5�L�5�F�3E(�%��O���� �|���O������'�W�+JXy:���2'�4�A�/��x�E���'[jE�w�ϭ���� #L����<�Z�	D�ɷM�x�It�˵{��HK!\�M�~B�I�( 8Z5�V�3YPc�x%�B���M3��A��0�⦭4 xٓ3��P̓UZ�h�#�iM��'��,s��0�ɯ,�|��6dI7N?V`Sb�w�^��	ן4���<���D�!+�@���*u,��P�o�a:2�Ex��A��uIJ!�ߎ{|�Id���ɾ��<�)��&.#x�[��� _,Ż��Z�;a�C�I	
��ȡ�����2U0!M������r�'�Ѱ�+U�4}�<�u듾w��J��i�B�'��n�[Hؠ��'d�'��w��!!3��:��Ų���E�<Q��i� OP-�P���_M�S=*�1��'Yl��RP�?���U)�I&�����B��	��ȇ�j�T��DU�����X�,)	ׁ�?�`y����'��"�i���'^��C��d�'_��'"��'t�T ��|@$"��F䰔btO� �4ƍ�EFe����r(�8T��p1��d^}rX���	@�t�CΙ^��q;5!̐\I�D0��şD����L�I��u��'\r�'B֙(�0f�pxD�63e��cT�z!�DD+W�,H�t`�]e,+㎗�(�4��F�y'�ؖ��h؞��5� "l���5�ٯnx�X�Q$L�R���d�O&�&���Iɟ,�?��_�K�
M��&�Hwh�`�$�]�'?H����0I"r��#�pd�%Q�c�6wfx�O|\m�Ɵ�'��*�ê>��[Q�5B��D��l�@���Z�,�i��?��b��?������n� ;B��#��h���#V�6g2��S+<�,��K�<����9%������)?� ��D��:�p�	�D�6z���b�1�@x��'�0����Uś�>)�N��$��Y��҇w6�=�� r̓�?1�S�? ���CƘ*
�D��jͩ4�Y3FOulڮXq&��$߮6D��RE,E3A���IG̓�MG�,O������v"N<A �D%�$�P"O�e�ņ(yL�����15���"OZ�r�$��a8�b���x���1"O^��s��PH���	��dF��2t"O،���^e\4\@R�ѩT1�t�"Oԙ˵B)s"&c6-��':H@�"OV`��S�eX h�Ǭ\Cx$z!"O�<b�E��3��\4��$�@"O�s'/�b|	��j՘||ȕB"OT�"�ч�$z	Ɯz�)c�"O�T�G.�k'd`Sw�;<�v�t"O�Rrc+C=P��Wf�)��u"O�a�'j ������I�6��"O�أ��, ���)]ְ�a�"O0X�H�)�(0"�b��X�.�+1"O* �H�.0�%�Uo�"P֬��"O�,�S		 d��W�ϮX�"O���0$�7/`�}r���"� �a"O�]��C�$<�1��D f�2��T"O4�$f ;S���9��o͊�"O�Qu@�)W�$�̟\M��T"O6(��mE5Q�d@���_�7O��!c"Op�m�%K�(P��W(B�y�w"Op�ǁO:䒼�"�B�����"O����ȏ,v(1��O+/�nXk"O���d�V4V����wLJ�#�Lec�"O�`���%P�� IE���X�"O�5ۂH�.m&A�e��4+�8Yɦ"O]�&���u:�ad�V�z��Qv"OhIg΍�M�:a��]'f�D�D"Od��+�K���%��
K��2"O�� v�
+/Jؘ���٢g���0b"O�p�/A��MJ􉍢~��̱�"O��Rg��
�p�@E��#'�n�$"O���� ��Xh������+y�]��"O��#�D�'��S�PE�x�a��8XD;B���t�/�g~��ԗ�tqr���6G��v@W�yB[�&4�&c��ID2�9�. �wL�e��aCn:f���)�����^�*�@Ra�L{bͅ�	b�J 鰈\�9���ɣO��]R�E�d�zi���)K��C��/�(ؤ��G���",o�zc��ӄ".k�j� �#�'TޖHB��)��M��Q�S2���a¢�ys�Plpeh��A�`g��R�,ۚ3�q�'��@3��0�^�Z�<�7�*$�j2D���[�3��+0��YN:!��͹zr�x� ��;�����$Z9򜃗�/vȉCr�4:=az�Ȅ?���s��y��C7L� �K�^P i����y�&N`�p}	�jL�fr�-!��'�v%2%-#Ed��A��IK�N@�1%,�.����C��x!��˨[D��EI2޺ЊD��<�����D\��'zq�#|�'��9Qe��c�J�����y �i�'j���ŝrb�����Ml8s#�"�N�i�F�0>I�!I�}�4�E�8x��D�T��И"l�	됩�Ek��p�i˝hٮP��`H�M8]:�(D�����&�R�Ӂ��	�LXj�*��
�\x*e�˃.#~�Ă	>R���j��c���X�o_P�<A�b�74�� !0�U�/
����J�<iF ��V=� R��$!}�t#Ch[�<��NѨN�كa���5��h�L�<!�,�0?�`(��D!cT\y!��GR�<)#� <�j��D��Y�a��L�<�tE�>,�5�A��!�di�'ɌK�<� \=K�?l��ّ�X�����"O�aХ�N�Sp�%�I"p���Ƀ"O8aևI�[~��#��>���q�"O�]�g
^�����w��A�Q"O��{dj�:��P��>�j�C�"O�pf�-|!�,�3�_�����"O=�p�^8M�R��f	�	�|�R"O(ě���m^���V��4 �����"O�M�2�	q��Y�b'�"ai��� "Ozܚ���8�0��֏�!gNr"OdT�Ջ6ɞ�Z��!6(:|zW"O|8����"��;p4�U"O`5!��S%`�@Han�Ct��0"Ob�Z�GX���1G(z����{�!��%A�����#cK���n��%q!�Y$��X9Ff��:8�����\W!��ƞ:��1��ȝS(n��P'� ':!�ğ�#>2����ǜ#
���f��O)!�D�-0�fH�Dʅ�;Vnd��,!�_(���q���>eCr@	ep!�d�M��ˡkI��D����� ��<����'pB$��!O�P�2�b���8CF�
�FL��I�=ƪ��aًD'����Ҝn�z����&0��' ̪����z�)����w�ъ���^���J��I���p0!�I5x��q��2Vt�O��2�4�)�.�ꎾ R @T�])��'�=@!�)�'v��CQBʀ8��TQ�Q�7\T�!�C�T��'�D�G�,O\��go�7���BEQ�Ig�D�C�O��A�O�צ����M&�p<���ԤJ���a�M+�ʄq�(�y+^l�p��=Q��#?��&�B���qbB%<~,}�ʂ<�l�UN�.,$t�c�3�D�l�$u�g��`,,��C��m�ԟtȠ���?�@9�Y�!��y�D剥Ld��3��;�`y4�� fe ء Kc �-����#ȎbR�]��e3
�|O\��S��cH��S	il�)b	S,X y�̉6[D<����G��M��	$g��)��@�`�ɽ{骰ZS*-Č8��I^����u%�� EĘ�[�`֝5fw�EyR�]yh���A�&�2�5�B"����ƈ��pq(�(��\>�`J<�T�A96}�Ŭ
�\z�)�#Ư^Kv�:�����	����|�pݨ1l�s�#<��.!F)bAS@��d�!&�\�Ed�Ȱ)�c^�+��f��O$��Sd�+pL��i����V�6d@�D�I?��O�>��-υN�����W�:��,)p+G�T�X�u��?jq>T���iP�>E;bA��U�+6!J�eF�Q�'��0�%H�M�Bs��q��ϻS�MЗ@њE۬ԱF���Q{�!�y�4�Ko���10�w���S�v���ω1A��lq�G
U+ 4���'z��d�6Wop�R1��"٫&d�?c�@��'�3>�t8qNў,.�#`)�|tr���A��͉b�_9�RO���t�7Jz9l̘��jM�L@�O
����֬)�:���L�$Ty�#<�*�6.+�����][����-�|P>���!
Ypu�� 
��O����QTܨ��ڇ�:�"@Y�擛>��P(�	̒E�7Óc��p$��Df��RTjA�4��D���I1��DnV�s�-��_2y�L���Ѡ.dft;s�"A���)�S�yW%<����A�T���e����5�*B�}���	���a�X��;��99���d>yf�т��Оs���_w��D{���1�Ä@[;Q�e�M��t����'�z��/ڲjB������	F�9	���.y�x@*��#�z�\�)�p���r1�Ys�X�����*}=S)�f瘸r5-���1�R��1A�b�	��%����ZF�R�3�\��J?����6 ��`�bS5q����u�#�ts�MCҀ�2"&uS'h:���45��KSi%k⎐�R�5N�PM W��TUP� �oe�PD��O�Ă`&N�"(�a�2N��VІ}���OZ4�ʔuJ<�¶��%�0|!L����1V�k$&q !Ц�Y�#ɅX���f��� ���I,R��x���SQ�!r��^1��b�(�������K�¨�ם~r��3Wx�R��C2E�I �h�\z��Gn\!� 4��ǋd��p�cEBæ(y�M�3
��5pw�ÜZ��Db��C����^����*Ҹp���� 7d�d���2qhNt���S	c��E4������Rg��*���(�NŊ&�^+2	UV]� �D���R+ԭkt��Q?�V�>����m�fś�������#��w�<Q��/+��X�㜘�>�xd�ͦ���m�{���5��U��y���T��&M��3U� ��=1��	!8&j��D�g($@;@��KT�R2C���Ԙ�F24�� ��Z������W��8Hz�Ѓ��_�X��@c� �Q>=I��Ҹ$����*"��J�+0D��� , �U��ev1��a ��>���'�Ȑ�q�D�i@Ο��|���.o���x �'P
8l����@��,���,{�0�P���B��"ѡD1*3t��w
RQ7��=E���s����W�9���1f��E���G}�`���nً�dD�zdQ¡Gcr�kea���~��9b�8��4V�x8��IMƖ1PK�u@��	�j@:Hr6�)�)r�K	�qH�牪s�q����.Che� �ə\�.B�I	U��@sgπ`� ��F�/>��'� a�aA�Wl�k!j�X�S��mC�\s����ګZs"l�$�3�p?�aLK�	�b�X�R0i�:C�Մ-G��Zc���a8<%��0�)���ґL�>?S��:tj�,S��5!���ͳ�%�n��VV͑�I2'J�zA̀5K��'����əSN8�kF�Id}8D���I5X;�mbC�"�)ڧ~:�8�߷,n��˘%u̸Y�ȓ
�\zu�G��P�C�"W'�ႇ	@>���	�E�Z���G�hND�+a��
�'^�������"�R���+�,q�� ;�'fv�b�$]�h����e�y���dF"X) 
R���'�lQ!ІCZ,r�*�1!���}KS� � �4 (`Cb$9�'��%�0ɧ=ɧh�<��%�*����W�U�l��"OƩ�l3�И:���Vu��>q�]9 3���
�Ƕ)�G�Zj�F��0���y�@���2T�L<�&ܑ=b���L��^�Jĩ��L��=��)k0Hɵ�߈xЮ�	��L�M-�mG}2��X��ȇ�	T�Sឱ���ɫi,��mH5V�!�$��2��W�XF��cs	)Y�^���r�x�rrG���S�O���� P)p�z�C�k	K�f��'�&�@s�O;F�F)���.G����L<���r)),O��Sv��(*(��	 �$4���U"O@�ʃ��S2���(�ho�t�f"Oș���ۋ"dVPr��� ~�P�"O�Q)4�[�p�A���Z�$5�"O,0�)"<q|�*r�� 9�D"OV�� _��P��BEy"O<�iea�F�8x���-?��k�"O 90�
�(O\x@��D�Hks"O�虷�K�?�|�/E�b�0D��"Oz�:�a�$���{���T��t�Q"OjxP�Ł�a@�c�1y_��0�"O���C�Ι0���p�ၑ==	�"Ox\��AT�tQ́@7�7i6���"O�)�RKD�SK=Q�	
��p�"Oި��k�2"G�p�vZ:u�f]�"O�m�F�ܙn�@[���,��Qd"O�0,]��Em�)���Ӣ.D�D�r(C�D}��ɘ8QG�e"B��o1n�{�)��]������00*B�I�/�Rq�X!_��mawɞ0k�C�	8����W�������G	S\~C�ɻ9���Q�aG�Q�%�6G�$�<B�ɒb<�� à5�Vye�8B�	�Js�M'�ef��`-�' HB��wD�p%��6 c\���C�	�4ìLja�M5z���/ �L�C�3i �� *݄8��q�Q��0��C�	��q!Dȟ�
v��H��r�rB�	M�h�Ǎr⒬���)T�B�	�^�:�J���Qt4�#�R�|B�I�^7��teY�]�b\�Nsj�C��kP�@@,R yh8C��:]_zC�=)L���I�0AyX4��*ޫ�NC�)� ���@�ܑ��â#6�2�`�"Oj8�d��R페@6��dXB�"O�M�`E0�l@�J�d� "O���4
�:ʌ��AN�'�Q�"O�����7k6��ʇ��x��q"O��3� �GS�U)�oCYy�TrU"O��b�-2]�	�0�7re�s"Op�j"$��<�F�R��13T|��"O�<�Q���4V�P���P���"O0H��Ih@�rb�>oN����"OL��.�= ��t
�730�}�"Oj�[���{wx���0D
L�2"OzqC��/:�(਱�7` ��"O�XG��-�<5 FB�%gc��ks"O�4%"�?
�$��!�ULX��"O�Œp"��xPRC��1o9����"O���u	ҙE��a��
�9.\�f"O��(�[�NKV1�Ώ�62�[�"O�Lb�a� _;R�{W/�g�HĪ�"O>l��Y"el@�$�&aʮ(�S"O"d9N��0�*���㟴���Q"O4$s�;N��ɻgCރQr��A"O�1� |$Lu�g��;3``S"O��!r�3HVl�J$]���i�"O�񀐍X�kz��n�!�,��"O��N�3�Ġc�]�ov�s�"O>�!��B#㦉����-/B�e#S"O(Bnۛr/�c�a�1.��"O�S��רk��	�2.���0"O��2Vc�!f,�ŪH�&|�)[�"O�q��۠%
ƀR�A��L2���"O��cj>-��3� ףN��k�"On����0�-��i�4)�"O����� M�L�M�2H����"O^ ��΀�����	
!&^J!�"OH,1Ѯ���F@`�EP�)�Z#"Oܤ�U�\�O(��Ņ�&hj�kD"O�Y�M���t{���!:hx��"O�� �␎K\ �f�Z*&�N�S"O��J�,�?�4q��A����8"Ohqc�S�^���`W?d�$"O�x�����O� ١���]���"O�HeB])�6題|M2�)E"O��
U���<3�`:
�+/(4�D"O�|�weǼ9r)����A|r���"O�U�fo��
���c+�o����"O2���mUy&��R� :q���3�"O�pp�#r���E�9,戣�"O��	4͏�1/$�Q�HסW��A7"OH�x2G�RF�zH��kn٪�"OJ\�7*��&�6<���!#�t��""O�$3�OF�{Q8������t�H�is"Od���k�
vX��6/D�v��Tk""O�x�P�?kҶ��d$�7�tYt"O P歃�t�X"�?+�R��"O��[RM��"Y��$�ɉ*�p"O���x�۔)�w`�]5"O$�KqOP&<
�B��	DXq;�"OJ��U�rpNp�I��<�m8�"O� ���A��� �1ba���[�y�䂁)�.�8�&��Y(�� ���$�y���CT�rD'��
}�qG3�yR�
I�s�
�|���¥H�y��	:"/�,�$C���@ƢG�y
� ��C��ĸ,���0(E1
`41 "Ox�C��:%j<m2���;$�
W"O�XC	���9p
DZ�h�t"O���Nz��]2B)�q
��s"O�3�j�SԾt��g�D��9;G"O���!0ڨ�{�EƂGڒu��"O�%���Q*[���n*݂�#5"Of�p�?�4�A���>�P��f"O�a�` �BJ<Ժ��2�K�*�yrc�]��@�!�CLO5�N5�yn�NKF���)W2i�jW��?�yB)�3���a5��3"���Q��L��y2��6Ks��agH��T� �)�y��%S4 ��BhpՈ
�yB&K��`�V�G~�Eߨ�y���Ju���/ܧS^��Y�.�y"�����������g	֊�ybۖ(cda����:s������y��, vy٣gŴ�BD��cS��y2@�D���m�Z�+w$���yr&�(<�HؕF]?R� )7-��y�o����i���B�6@�*&I��(O6����_�^��F�S
��s�jG3G!��REIv S,�>5͐�P6ʕ�9!�č?E�|�WjW��vD�b/�� *铨�>!f�_*��-�čD/K�8��U��C���!�����A�l ؜��)K'-��eK��:D�4�qṀ;A���`�
�s�<]���3�Vb�D���l�(q	 E�${�,����y��˫B8��5��<"��r!��y���>8��W�7ޚɃC��=�y��4��`P��߅'p%Ȃ�� �y�, 
SÌ! �I2�� ��yb%�����*���(2k٫�y��Tl1�A��}� ���G_7�y��΋*-��Y�HEGX��Ј�yl��k��X!�!��:�^�!@Ԑ�y≓7X2`��7�`��JI�yr���}�Q����e�:	��<�yH;z�< ђK���|�ae΃�y�j�����"HL�����1B�=E���X�RD�����L��X���z*ȇ�[�8[W�E��V��g��\ 0�ȓ[!6JB[�iq�ԣP-ˣk�:̈́ȓ/���gZ�V�p��a�H}6B�	=}�͙���p[��a�bB]B���>�H>9P#�' 乹!�3*^h�r��f�<ф�ٹ3��=��M���|��O�L�<��/Ϡ:�rp�peY�
�� �H�<Y��B�pM�uPHL�Z��M�`��\�<��2�e�!j1:0��&�>Ii!�Ğ<	�.�P$O�6,0��C��0Z!�$��8Q��A�'��M��vH!�RQ� �P�ƛ`�����FWU!�Da��oӷaq��&.��*J�Q"E"O&�Z�	X�_X80��N�*6�,�"O�͉������M �h�T����"O�U�T�S8v"�H��C�S��33"OD�����;|n(�!�'V�(�u�$"O�T¤�ŜH�H��a����!�"OdC���kǠ٪S��
��s"O�b%G��|t���i�l�B"O(�`(`-�QѕaP�:#�1""Or��p��*��u��Y�u&���"O� �YE*�2�X�*F�Hl�*��"O(�
��ªS4`B劇��1J "O�Q�'���ޘ���ʫ[���2�"O*���	&7��E2�q�� D�4��)ͧ0Aj�zgG���͋�1D���U㐶�
}��R"O�es�@.D�8���E�G>b-�%ύ=ahA+B0D���e�Դ`�h��P�0{I�{�	0D�h���[ ��ZƆr�fQ��#D�d����FB<�1���w�2e��C'�􈟸%�2�<�� ��,wi�Q8'"O�!K�\O�u�AB�T���"O88���=a i�b]�zQ��G"O����_���0@ŒjJrTk�"O���0K�����$��+���'"O(}k�L%3���h��ք2�"O
����̔Ȁ�Ѷf"K���8G"O6��g��U]� �F��HjV1i"O��g@w�(���GT����x�"O�Tb�hV;.�����+f�Z�q�"O*��7K� ���N��C$"OB��P�@:k,Ը��Ԝoh����"O�\6&#T��TP�x�ܠAe"O�%caE8XY��4n6e�2��D"O����aFA@|�7#:� � �"O:`�C�
@�R�ʢ�
5Ӡ�:��'$qOZ���n]�]�U���64�0��"O�P��L>M6�8b�P����C""O�49w)���Y�p"����!"O
i�dH��z Z�Z� �6� ���"OШ���:�@����B�C����"Ob́��QgZ]Ҵ��� ��"O�xCMڧ`�@x(��B:W}(ɊS"Orp�<v1ΌK��P�ko�U��"O�0�h��G�̳��(ø��"Oj��$��e��)��̺e��A�w"O���SL��#�m�d�\=���8�"O~Q�%���d�%�Sd�0��W"O9���=+D1�r�Y=7o���b"O��ࣄ�5	�0��	~��aU"Oֽ3 ���z��#<����"O�đ��ξL���j ǖ�S��8�"O�سU�lܠmHw 
���b�"O�0��i�I�n�7ŀ}���I�"OԴ�5�5�`0�aD�S"��2"O�,; :IP���+Qr�*O�����7'h!#�W�l:���'����ȷ_��Ih�MI&b�b�Q�'�Rl�t��,N�PA���D�nՋ�'��h�I��8���0�N�?����'���%��@�d�W��H�Ȭa
�'�X�:��߄����C�4>��x	�'l>�P#�V�6�q�S):�Д��'���s���M��a�@�~]~H��'�����e\Z 2��'*A�h��';,h�#��;�6�zЊމJU�� �'���ۦ���lȉ'�F2H_�4��'`m����{�M���Z8:��Q�'��lZբ�U+HcD�(:����'���D���M��!˳㉯�����'�ڽ��b��&LZ�k	�b��'�>�i4E\�Zid�P�Ǖ����
�'M���ł 2%��� _.,��'[���r	�3ߴtA얬\�t���� �5�HW37G�y� ��<AF"On�	$K*.n�S`n���<���"O��+��ƺ����#@���"O�tS4@҄R����֢Ąe����"O�xĎL�wb���2GշM���`"O���a-�#"��-HC��J�b�R�"O�%;�&֜!��Tsw	ʃO��3"OL�b�^�5�ٲ�(Q��T�(1"OR ��Wh�) M׏@�
d*A"OxM	�HK��Yu���F�(�"OJ��
(i�̬�G�U&`7
b�"ON�9���
@4*�%����"O���%���"�(X�Y�k"OF�aA�V�n�jx�G�+,����"Oޠ�W��3$�� ��;@�
1 "OJ�VÂ=Ft��Rb��cj�:D"Ox��7�^�"�q#M1�t�f"O��CdX�O
j�A�{ (3u"OP@�S��*�|���oJ�VQ�!S"Of<���F��f�a�]�/;�( "Oz����V�[Wz�ϝ�:����"O�P"�ͷ~��	K�`�!Yb��"OnDR"o��$�m
���8���"O^I��Ь}⁮;�X""O�Y��J&n��ٵ�ɭaj��"O��)dj�1/(F�8q؂�,"�"Oi�t�O$�<u�կ]�T��Q�f"O0 (����U�(�� E	R����g"O���֪a��!j�i��	{T%��"O�F��)���A��Ra^���"O�8����-o���B"
D�^U"OT�TM�,&�(�LU�љw"OP�pu+�4R�T�S�A'C- R"O��� ��7c|qk&�R�b/��"O@XY�,�!g��1\�9��I'�yROL�F51�ÞZ��i�#�ݛ�yR��+eT@9"�`��4 �m��y�AW�M�f�`��:<Pá޷�y�#��<kX�)�D�.)�>���]7�y��X�+i���@�'&�`B��J��y��ɨI@�-����dv�� W�yrE_ ,!�Aa�HO���x[�e��y���Qd`4P����ea��y�9�� �g�6���b���yҢԸ_���,ٴ4*��LK��yB��_��x���TqB��O���yR���X�A�dҵA� g���yR��%)|r�1���n "i�����y�a �v*�PdD3Z,������y�lٕ;���j���"�
=�wB�3�y2ÙN���+E�0�\&��	�yb���K��H��FT	*!^-Pf���y�*ӻ2��p�/ε@�Ɂr'_�y2#�^��@{��@�pQp���y¬�6�(g��x-`Ur����y"�I2����DtA�Da� X��y"�K�
��͸g��j8a����y���mJD���'d��E�cd�<�y��
�~��q#T�U� ��ӯ[��y�B��_�ހ!S�$;�0��#`\��ymBQe,$���U 4��a �����y���X(�\�����(�,mB'o���yR�,a��]s���v�['��:�yBj�(V/�%0У�K�t�y
� *	)F��(d��p�A��J�@D{r"O4��j�8YC������c!��"O"��� �%�Ȫ��Z��q"O|5���h� ��#c&�a�"O��0��� `?J� "�ѷx�s%"O����_�@h��0W��N��\
V"O�<���Dtj�`Ɓ��Ai�"O�܁q'�.:p�a����~�ցk%"O����ܲ)01L�'y�p�Q"O�p�RKV`��9CP�Çn^|�R�"OF0�7#zmZ�,M���a�"O�Պ3��"�6�q��O�I�1z�"Or0xe�W9.�����xÈ��"OI���?I��4Ӵ	E3O����1"O�=҅
�2�"v�V�OuR`s$"O:1�n�T6ʘ���c,܈�"Ot��a�O�>�Vaj��WbO^�� "Oʌ� a���,��%W�����y��G'O���G�)o�}�!�D�y献Ae9IW�Ϸx��@rE��y�,ֿ+pT�p���p>��1�S7�y'�#/��rDjR�?j�������yR�ޒa�؅�H�!�L�����yRBM�Yh��{囂�z�B*�5�yR��(7����Q�g�~ J ��y"-�C|ؑK6m�P�ے&ت�yB���Kh��iH|�t�P���y��U�Ҙ�e�oG|4R����y2�D�K�T�r`��c̘�&)N��yBG��?�"M!'�כ[1X��e(��yR�_�f������M|6I#����y"솽H�	Q��J�7L6�Sa�\;�y"·8	uhذ0��\L��˻�y��فsL�1��G�O�ԁH��ũ�yr����;�ܝE|������yrϟ�wI���"�!(?P9��
=�y�+G	W^qѢ�P>�x��L^��y���9�,�[���+Y��l�R�'�yR�*E��y �h���h��]��y���>t��	��%�D�kO�y�Bۃ%2�a�-�6x�f�a���y�fA�YSȕ���r>�|Б�ݽ�yRO�FL����P�=>�A����y2�](Y���jA-�>@�i�G��ybJ�&���Q�֫=�F�'��y��D9%���x'���.�dAF�)�y�+�9e&��(�.��e����yr�6����hT9O�`W�е�y�
�>=�60����)%0Ijv	Q$�y"� Gת	Z�c�(v�I��g���y�F�)���@j"J,�{*Q��yҨ՗S)�=���6h�.�y�@��A���Aa1�����y��+f����.��4T��g_��Py���"E��SG��
��Ɏq�<�6f�%(��"Ň�0V��U��V�<9�[
#?�a�� �-$8֑ pHy�<�1Ϛ�1�-Vv'p��E�8D�L�U,��r6|iqa�ҁX�Z<��j*D�B%�C'-����"�	u�	�4'$D�X!���<	 p*���2Y��D��>D���G-��Q��U<ڸ� �:D�X�#�E�|��su�s�LP��9D�kwA!#�9"�ʰ7S�@��9D�� �xs��N�48b��p]`<:t��"O:��e��0��P�S�FJ�"O��Y���3]���E�3Z��j"Of y���&�t�A�?NC�@s��'��$K*&>a��`s���&�)r�!���(5!IX�����Ы@��O:�=���T��,I>	�1p��	��,j4"OD���@5$��<��ƀa�v4��"O���b̛����xbeܻ(3��c`"O�@q�Y�;�J�`Dװ�d �"O��)U%@9�ԊAC�9I��	�"OR �f� 5����:C�AA�"O��RӏG�z0(`�I<:0�	�@Q�h����i����/O�&�
\9�mC"9�C�ɧ\
�Mic	M� 0q�v̀Q�C�ɬxZ<�c�f���z����B�	!D�MYP`_>#&-����'I%��O���!LO��Y��}�<L���x�� 9�"O�tq�M3�.�:F͖�"����"O�� ����L�4H
0g7J��|2�'�I���:X	���5�^D^�Y�'o,x���:!��UJEj�����'���ۀ@9(5�
�BF���y�O�M���p��%��F����'�az�U����`ݟr4�-Y���yR���-R��7i�<B�`˟�y/�<Y��J�%
+a���aN-�y�L$}]�X $u��Rh��yB�	?C���G5O	�<��&�Py2�^(�����$zH �6�_t�<y�_�XUn	ib�����p�.�r�� �ɹdt���`�JpA�i��"J� ��jF��{DOY�G�����k�,ȆȓD��@�@�!�<��G�T�5`��ȓW�aÄ\�h�l��gkM�l��=��^Yʕ0��5�$A
1��^?��ȓP�@�f���wHdb5�%>���Dm�HW�˛UeL�"Å %5�� ��W4.�c��W�<�.$	�&��U�$i�ȓA�u��������AK�+ ��'��D{��Tcd��	��\1�.�t����y�J��`��6Pp�հ�y��R�e1HHc���-�,lY`-�y��K�#}�!d��<<�a4m��y"��+ ���!p����=ғb�	�y��B�g �Bq��'c$���X$�y�U	H�,i��Fºc!T�jC��<A�����P���Lد$!�8���3LoV�OL�=�}2�-ʬ~D�R�� Kl�$�I��<��E�\_`%�'l,���D�<�W�ZJ�����#CyT�zd|�<Y��O'c� R�lãf�\\��Ba�<	�͚Y�Pӣ"*e�tC���G��4�<�D"��Xʬ�S�R�$����	A��T���OP�Tz���"K�-��!�%��q����5�b�� DD1��i7MR�E]:\�R"O�����_�!N(@f�PQ�t�R�"OH�QB�6zϔE�#i[�d�"O�а!�yM�p��փo��8��"O�+�6'Hā��"O{��C"O��a��5Zr�M����ٸ)��"O.�(TeW?���'�4��1��Io>���2$�f�V%K=kZ�ukSG7D����G�$.��sɈ!sU�e��:D�� �]��	�e��b�@ǻs���:�"OF�ʧ�ٿf�x��V�	
f�"ݠ%"O�Qi�H�@���)!���2�L��џ|��'[�h E�=G~��*� �BT��'�&PcD*�wB�I����w0��ڎ��7�X��j�_�6�I�!R�5~@P�A"O��	�`�4%?t1"�n	r�L1�p"O�U��D]�e���&C # �����"O�%;�`O??&ı�g��`M�I�B"O^���ʇ��KS�\%��id"O���Ai�z�8s�d��\�"O��@�
)U��
*@���t��U�O!ʵZ�`QR�n���!�� �.O���7f�^*�C����T�1 �f�!��B]+��Krt�ݪE�!�d �t���@ /��!���I� �!�d6��8�]�3�@#�K�XG!�D�M/�u9d�V�O��!��Y#�!��-v�$u$'I��E�5	O%n��'�ўb?�X�b�M�>L��"ִxV��g\����I3I� ;�9o,#V�pfC�+&WȠ0��PL R�r&�8
�C�ɉ^!h�P�M ADؠ�BP�C��B�ɬ%n�9���>2X�q�N	"RB�I�1�Z̢��H�mlTC�
�&\ B�	�_$P u��>`H rDG��bB�ɂV��q�2�F"6���"�)��C�ɰ �j@�	�	7��YHr�9$�`B�	!S��6����&A�p�@�m�2�=��'@����l�zL9�E�B;`���FR�����@-F�tٱ4�V<�܆�wv��WJ�4�����̺Z��0�ȓW��TJ�		�JSd��R�R���ȓgE�x�dX a��-��P8$��=�ȓ~���aea�������1^��ȓQ'$�kҨ0(rd�ThZ����ȓ����1������Ŧ��ȇ�B+�1ah s�b�H�`ӭPJb��?��,��q��B!N�@x�ç/Q���ȓX���I�2���X�&Zeȇ�;9��R�C�@�Tp��g�b��|�"�)D�J�)^,q)����`B䉗nY�8i�+ɋ7�
a�C�{�|C��/kG*�� h�B���:nZ@C�	=*���4iy ��	PHӍk �O���D<�z�9�+\�-A��q�(�ў���	�z��ar�ǄS~���smJ�\�8C�	h\ Ku(W�L�H�����.�C䉘N����[�[y,�HrK��r�C䉲W�ٕ���u1@d1�(� x�B�I�`�CV�V�6X� �7D�D�zB�ɇ��-+��?bM� �Xq@`5j���'��`o�<�4�rŤ���ۈB�)�df�Me@��c�'"������'��'+��'9
�0:`�D=���!>!��V�g`0#���-�,��F�9-]!�$�*@�nUa�fX#͌�x�&�%!�D�7������1`���d <!�d4e�4�R+ʕP�1�6���)!�d�
ir�����˙&BdMS���)K�'bў�>��N�z�`4�2"�x):��A�Ic�O�"H��K�	70����CF���'rN��a*FS���؆dX�'��U�g�A&Z�x��7c�<������ �X�so�sd�)%@$i8�X��'����0����#ԉv��x�u�X�]�!򤋞y��A6J�)�P!`�C�1em!��Y���#c�_�TH��o�<�5O�����=,�Z��v�xq�"O���@V�J/��1+�>�TB!"O,�!�
π|�.� Ӓd�X���"O��ʤ뜬UT���cE�N�`I���'�1O��qBӯ(�՚XY&����ៀ�'�ɧ��N�"�
��H���w
��/��-<D��١� ?�����f�	�G�44����C^�"o� �'�R� 3��b�<�#]�����_Y��RP��Z�<9��1J.�q��"��C!z�#a�*D�|����7 9���b��40���1eg)��䓹?�ʟ������P���@&�f1���S�XG{��i�U�Ddc�T�j�D�b����*D!�D�4��JcG�..i� ��34!��D�� aAʖ�(V�K�CB�9�!�DQ� F�$�c
�5
6��S�@6O�!��V�]�����Ʋ7�I1��#!��P`a��+N
tVոC@U��O(�=ͧ�y2����%�T��v�`C�>�y�F7X�Y"E�K�$��!�n��yR�@�~.���WGK3;�X�+�l��y�jte�)PBfV(=b�8���y򩆻X�|5c���D��A�����y�/��.Y,YX��֍;��Qe��y�*V�w 4(y��I:,�`�����䓫hOq��i�ݰX��e��4M���J�"O*i��;��u8oH���T�"Od巤Q�@� vhbY1���y�*Y�� J�P�A�ZX��gX�yB����.P��$��9�d����y"�_T��qjB�9D�0�cT��1�y��Y�`
Z0�/�Xi�Ç���?a���S�q|��� q�ȴ�Ӫ �ގ&�Ԇ�+�ruӢ�_�"���D5
�C䉺)#ެ)���k��Y���fǔB�IV5P��A�Q���l�O��.�lB䉎u�2YH�H��QO��ye �r@B䉣xك�i�"������(qu(B䉃0�z�� �,n�	��\�p^�C�	*�#"'M#���\Y���$�O�����/^Ǽ����Ӹ	7� �L��'�a|R��	ejH !Ő�n�L	�Wl�=�y��S(��ժ�!�h�i����y
�lƎ<�bC��K�bQ�v��,�y�!A�CJ��%�X
lc�eI
�y���c�X���/B�܁�ؙ�yR�	(g�[g�.@��:�/\��y�-R.K�,h����<KF���y�*�Og�����-J�q�&l�y�D�(;��ȃ��Tp�!��H��y�˞%�bH(�`��`B�І��yRn�2Ud�s'�'�Xd���G�y�f��F=5�
߯/D��6Jլ�y§ 3	$v�!�G�)�,щᇇ�y�*�w:]0gG	� ��Õk���䓓0>1sJLL�v�[ �H�5Z�|JG�WC�<y��B�6PJcn�[���1�o�t�<��d�a@j]�C
H:usNHie��n�<���K{[ެАM��=x�t����g�<�@.�$�|kB�[P/�`ąN�<� n�Y��)#W��B0�Έ52��j�"O����FO��8b��D��h!U����	��:�BGm�@̘9��C��B�.-D��mL��0�b�'Z�bB䉪(pHt�C+��,��b�/q�B�I�JlhUXg#H4x�h��L�=!ĢB�	���%�C%]��e3�/	��B�IV�,H��aܖ8c$lK�ύ<BB�	zd0Д�Վwd��'�=��O ��č	^L9ka��=T�ft���	U�!���n�2,�@�ߵ;��H���u'!��ܡe���u(I� ��Qo!�3:4m"fm�̨�n�)�!�	-4��=a��s��ô$n!�� 	�<rB�@�:�\q�3+�!�D���ӀfT�j5�P�PI��[�!�dӪ ۴�"7�E�! �=�u��	�!��C�lq��A�
e*��� +�!��Ty-�A�M_f�b�c+�5"�!�䆞>h$��ʛ=��b���S�!�/ڎ�r)�&4{h�[���3��O���$
�Np0�a�@�"�E�D�!���J�P�K�zjT�JS<
!�$�Y�U� Ύ�+WĻɍ1H!�0��}`U�Y'tFRp'��-�!�$o�1�'�ەB�r��匮f
I��R�jT����3'�<t��S�eǮ4��0ղ��Ei�.P�d�0l�� t2I�ȓ�b-����	"��f*F�O.XՇȓ
n�}��C�n�D�QL�ȓ>��4�K�b'��3D$!5���V�.�� ^:O�x�Uc�:����8[n����0{DN���0mb�Ԇ�:��h� W�.�,+rH�ȓ�Rl�L�H^���E��������IC4!
�,q�Θ�	��ȓl�z`��%�S�m�Fn�#�nهȓ)����jtN|=�aUV�4u�ȓS��q��!��JP��@)ev��ȓ��h��K�����j˧=��цȓbr�e�f�C�g0 �F�P#]k�U��m)X���;QpR�xª�E�q�ȓD�M�V,�C���4m�'�bx�ȓ(�.��͐�Sd�u�I�F�*-�ȓR{�t�sa�V�����"�h��iԒ`[����h�!Jǁ�G�����G=B���,�y_������Qz����>i��LFS|���+��_��m��,��A���C�/�QG)��@����t�������`iH>'!�9��ʞ��툤�/D�H�6��*�<EH0�����UA'�-D�P1�HJ(Y$Q���D����CQD,D��B�� �`�X$��KD�w�iJ��*D�,J�#H.���J��Td�Q�s)D��"Ro��A�6kxȪ1R`&�O�����UѲ@�C�me�yhp/Z�Z�d4ړ��OD-jb��L�H��+�,%�*��"O `���&�N���B!Y�m	�"OД`�(�<z�zh�ǡ�zS�"O�1�$Ŋ&�1� V�8t"OʝJ��CJ��Ю&<�B�Z�"O�۰aw�ꔘ��	���-I"O@�
!n�4ͺ���ܘ�:M�#�'��'
ў�Oļ�)ŀ����M�S
�b��� �#sH�1�H]�w�#�9�B"OT0f��J����ܡe�""O���7	�� �  ��)��q"O��׃@55�QǮ��Y��Y8�"O|-C���";Ă�����R���'���ߡ��9����,J/N5���7]�|��)�d�T���8�	_�1�ޓ�y"㑼^.@pB��L���� #����'9ў�Oufm���\�͋��UU��
�'TJU0��ޒ{����.��U#X��
�'{:�� BC�!��KS
?v2�
�'ܤ����g��� 4X�/{�� 
�'k4\���1�x�dAǶ[���Í�'0ax���d2��x��I�Z�#H��yB,�P�P�ޜEX���a*Ѫ���hOq����w��i!p�YÖm[�"O��2Ĕ*���0q!���8
�"O|}���*{G��Q�{�xY�2"O@�	�@�<\`*0H��k���H�"O�	Ѓ*
���RAG�[��md�'�ў"~�1EƼ}��є$�#9�z�yG�	���=يy��.<C�D�k
�C���2tό2�y�X�*�ȥMT�)�6��>�y��Ģe�>Չ�& !��,x�����y��9L�J�� �Y1����y�(�����F�X=JB�A5�y��*[�!��y$�����?����S�v{ٻ�f�)Wa$�A@[�j@2�ȓH�������<��	��M�.�=��W�l��Bb�7�V��I�*x촄� �2\��枎8_b�����L����ȓ#��49���?�`��\Y�^ԇ�.1�0� �T+�2%�0`�T���	��)�a��͜P�A�X��8�?��.\�y��K�0�q�ë�o"  �ȓrR��c�� 9�HP%�`e���rz��1#DVzt�!ůs��Y�ȓ���jS`�i �`$)���F��+�\�#bK�(R@h��F)�X�ȓt�H��9&Ʃc4G��cptȆ�|y�Ԛ�L�8'h�SӅK%%`
y$���'��>��4:�N)Z�����c�O<��B�ɌY&ب���� �.��-F�B���x�r�`�+���:�lZ2hfB�	�,	�l;� _!=��`3e��U�C��:Ԯ���M�Pv�D�fA��ftC��<2�b=S�7����a �~\C��^a�����܂��[B�a{ C�I�od���"�!xt����H�HB䉵<��mIsg%+X�v�m(� D{J?���	��S�:\�U.MX,���H D��QFL�6Up�i7�xX�=�5�1D��ca�U6E!��aپ��A1D�@���y(���0%( ��q5�0D�P�Si�>Q2�j֋UlxQ��d�<�H>�
�'L��h��P�[Ȁ��Օkv�A��x�N�Q�o�Ojv!ڠ*�_N�?���~:d։%l�`��+T�"�ӥ��d�<�s$L�L�h�'�&aT� i�^�<)��M�#����gG�Ei`X�D�N�<)�nG'f�(� Cl��[%\r�'�@�<YR%���C��:���A5F�ПhE{��IY1K!��X��"em4����H��8B�I�N���AE��u�8��%�G}6^�HE{J?� ñk�<S6h`�GFd�1�"O�С�lL?U���b!�&W3�@�D"O6!�w�є^�4�Bd�W l�I�"O��5�K�%�T�$�ڷD��b�"O�����R�a���_2G�^5��$�OF����-�=*5��*J�`ҡi�=r�b0O�EY��х9��ě2ٜ9�`��"O��jj�	2f�;bwD�B�"O�,q��
?�8mP K/Xh��1"O`�Zf�D��ur��4FI0��C"OzH��'m�P���P�YLxh�"O�$볈J�~�v\7h�.,�͑f�|�Im~�e
�`��T�c �8�xU�p����xB��V�zh�B�SV��훳 N�7I!�d(J����!Z�c�t%.d����"O8��@S�p0�Q��H�Q���"O�x3qH�55=\�S�m�4�|]��"Ou�$ͯ��eyb�d�l�1"O&�4�		1�~}�NN��\6�'w�'!�)�L~'��0��ɥ�@�
&�	� F��y"�ߧIIZ���0f� aˆ�y�����Q�S)(萣�;�y�+ЍG�*-q�l�R�XM���M��yb��:T
5�$�C�0������y�)֔P���e'G�,�Ѷ�W�y�V;�h��7D+`�|����D,�O�Y��fQ5<ײ,s&%ОO�V$�0"O�0�_�g��\��M<h��`�"O.��D�,�l��"J@���$��|2��5h6az�CPԆ��Aa�]�9����y�E��`q`�Yi�)�D��Q$��y���9I^��r��3�Hz� X<�y�*�>-���E��9�>���Ɲ��y�E~}�Cě�3�.C F��yN��.^b��}D^Pq����y"�\&(mQ��1w<uI/��?����D�<a����5e�Ԩ��-�PSE��!�T({��b�̻~��ј�,��!򄛑F�9t-�##MT����!��K��er�(��a�б�rO[�e�!��-)XP�0��E)�ʍ�r.�<C!��
	Z=�� ޠA5��hӔ^���M��4���̰>A�����"�,�P/#D���G �Y�c������ #D�8��`�&>-����e̮>�p��$D�,a��(���y��ԣ$�D��&%D�@{�F@2Bh}	�n�3�M�QE=D�h��J�?p8������ "�%H'�?4� �2oI:o���h��'H~٪���H�'ya|��ߊ&wf��Ӂ�$q���Co��y�g��R��H� @��i���*��3�y���sfz� ���a����(C �y�%6g����Oٖ[ ԼRbJܦ�ybM���B�jG���V+�I�Q��yR�߮+�,�"L�G��:��Ż�yRkOi��0���̀Ft��i��+�y�̓�%+ڬ
����f�iY7H��yRnKd� �3F��¡�f.���y��h�.]��u3p=�jψ�y"��E�%s�L�n'�!+�
�yr	�8��܃!�	:��p&��y�j��-n�����V�8z�x�	�y�_L*��҈�5�@�Z���1��$%�O��d�-8�Ĭ8&�6"U��9�"O� dDzI|�|h��\	5���b�"O(QI��!&�e�FG�7f�<rb"O��C.�%3z� �GJ{�=�""O��+����_�ZV�]$U̸�p��S>���A�; 8�a�G9�d�G�5�O��uP8��`¯>�j@�SiH.W��D+�������9L��U��"�6�a�8D��r��0����w��U�t�"��4D��6��.��Y�c�B���$ D��:�ڲPM�؊`c	
,ތ�uh8D��aө�#9Y�4l��]��)�Aj�<���#}*�(�(\�w숵0w�^h�<��U��} �ϝ>2F���f�IX���OҐ�`�E�b<��'$'9fm����dЬ'?�u���H��>��'V�^>�IJ��\�'%W)x��&ޠV�@`�J2D� y@,ʄ(�PbdJ�ޤ}�A�+D�X{욇37�t���_H�\PGf>D�����W� ��ز���;cƸW�8D�L"S͆-[: "�J�Z����7B�OT�=E�dC��'�$�U)�kj(�Lg�!��"gҜH���̆&Wb�
H�*�!��:Zn�I��O$%�\���� �!�DV:wJn9ڰ0 ��$b@�~�!�D	�'Z��a�ă%Ŏر���pzўL���+q�6h	���A��+�H,ZO�B�	�\Ppəu��7p��e�:R����$�S�O��`��N�<JƸ�!E�M�7�C��Wl�x��l�@�j4	��{���ȓc��1��Ȁ�!�Zy��*�;>��ȓXġ#���l*%J��j�����^~�s�@��y��m��-N6L���ȓ`���cI8\0��p�Ҷ%L*��ȓ2��`͝ 0u��:F�I�&Z4E{2�'�$z$H�1J"@�jE7)t$�����y�C�gH��OE�|X
R����D3�Ov��
ܡq��K�/V�e86"Ot1���ЎW-0�0W�WI�lB�"O�хJ�/.��6G�&b6`���IE>)��3@T\RA�ֳs�l����3D�0K�%ʍW�8W�S�q{�$	�
�<���Ӣ�^�#����5���h.B��D0?���؏x��\�%�7d�v08�kRAy��'�����2dI�&�١+#:1 	�'����)���͠v�L�o��!��'3VhxC*�m+��;eoʋZ����
�'1r���n��eQe\�=%V��
�'j��Y�T�;�p�PR!��O�%����hO?�p�.��V�rVJ�
�}�a�Hx�<I�̌A���Ǌ ��`ht&i�<���.m&�a��+��/�%ȷ��d�<1�(�
5"2�P���QCRd�2�K�<��ήr~h�"�T�]���#KI�<95��b;��C"��Z���І��]�<��B5c�N�хi.�\�e�@y�)�'M989���K�p�j�R&EXC4�ɇȓhfh�gg����ӈ>����_x�<9��ͷ+�V8�CL`�~ YŎ�u�<Ѱ*o��Qr+'|�<�`��BX�<�%�()d�&.81Zd��H�J�<Y��5]�D1KF2v�()B�L�<�	�*�5�a�	��9d[J�<!���
�	+�.��L�0��HyB�'��c��x�0)�@=�(���� |a*BO݆�\��ր541�"O�8�gL�	�����.����"O�c�� -�V�QɄ�.����R�'T�	n�)�=qBΆ�?ST �񄁟��*�	�l�<�P�\��`�A�8��H3�g�<�Q-O�d�>����ـ 0h����b�	I��`P	�x|M�n��!�tp	$D���4E �b;�=愁�;&�K��"D�8+& %r(X�_�B��SaE6D��
��X�d��v+�gG��P�A�<��2��m�Ba?8jh@ C�KL�|ՇȓS�j��g퓃f'*��؏n��݅�i�`�6",(��˧hY��r)&�0�'��>��*V	�!��B^�^�е0�k �e*2B�I 6�Y�� �̮i�d����yBȌ�d�B�&�dT�@Y����y"��ow��mG�X$��;�G���>a�O� Di�=zԠ,c�ȅ�^:��[ "Opܰ7-�7�����b�h�%ZG�|r�'�az"� �Ӡ$���(4І`_+�䓑?��D1?A�f�D�16bPcy e�wM^�<���Z+�� ��?i���@�`�<�eo6u }B�"�����@�OV�<��/�vb��Yr"Q<b�HŰ" Sx���'�dK�P�8 ӆ��$ڨ]1���hO?�	�.���P�S�W�h4�}�bdU\�'�ax��ޜ\��x�M!-�t(��ǜ�䓉��3�SJP���Oʠ�JW G
1)�b�<!o��4{���M�M�^�q�[g�<�A䜬1�)�ɓGݠ%H2( J�<1�/F�
�p���ʔz�(У�͆D��x�<�S���@	��"]�uk�˟p��[�S�4�'��	A$��$�T�K����CY�1�LB�Ʌq�8�����~���e���L�B䉅%��@y�k G��Z��<\�C�ɪfÆ]QT�&<?��s/ӫahC�Q�v�;�e.V����!�mVC�I�qcl��@���C��1�N�'(cLC��7��`�H�8}�W�̲C�ɏq�xИ��ԁR� Ŋ�x���2�S�O<����ތf���ZW蚶gq�d"OV=�U�V ����Z�nWU��"OD��:��yq�KE�8�H��"OB�(�cB
FJH�3%��o��T�S�'��Ez�٢F��ly�:�jY	a�L<��'H~ɩ��I L�h��dĒ�^�-(�'����	��7=YYtcί |dK+O����S�L�@�����P��OC��P �h*D� -��OUd�YUN)3.�ܹEm#D��%�]�m p���*@�.m��.D�0+vN�)���ˇ�4h��P��84��	�>Xr�ҐG
�Z.�t�Y�<�"��:X16H�ON�_������K�u���O�\"ыD�YI���C��b]	�'��"�N�K�R|�Th���8X��d(ړ�y�NY'_�"]����q�h�8�h0�y"J�+e���:� J~dp���ֲ�yB"۶"��HA� �p� �"����>�)Ozd��G��e�-�ʖ��C�=D���!J]
tT�T`��att�" �ON��!�)�'	�R�`q���t�T
E���Ѐ�'k"Y��o�$���)�l����$%��.���k�X	J&"p[��Z�O|�<�炂�56�����ڜZK��Y�B
u�<� ���	�&l�2YB�U\�2�"O���cD�2)i6����&gJԨ"O6|�F�x���P�M-N�6C�"O2����
���⠁�bp�X�6"O�DȤg���Ȋ���;G`��7�|��)�ӄ'�PU�ˍmd��˷�H>�(B��,yθ�ɖ C�L���ʀG�/R�B��7�Z,�� ]!�켺�H0��C�I�	�Rp��NT�|�h	c�:]r�C�I%\��y�"~�8�@�dv��B�ɡ_ hA4��`�J��QHS��B�ɶIT��/�o�>5� B v�<B�	�Hd��l��mx8�IF@´B�,k4���� (=�T��,Q�0C�	�AB���T┦#$4,2�nY8#�0C�I�_�}��"Z$7"�ZtN�e�C�I.8;�k�)L�)�K �n��C�ɅLX���7�[�G�|y��ž|�!�䙴z���2o��߶��vD_�m!�M�;��(Q�/:���_ �!�Dֻ�R���
[ͼ%R����!��ȓY	20��@>0^"���,�#F�!�ײ�x�B�8cpvh�lTG�!�D � �"f�~*��j�!�d@�`��BT�З#FP�2)�(�!���MP�����LKx�`��!�!�NJ�0����$�n�i#���`!�X�<9�h$�˶��R�˚��!�ĕ��45RI�Gޢ`q�
�&�!�$�X�8ڒo`+��*
9B�!�H�o��
�eC3(��HY��!��������+^*�!2���-s!�Dډu�Q1���4%K�N��!��u丼�$�ؐo�h��C�xm!򤈪N�j쫇��2~>�j�@�8�!�ό~~%��ס-f�e�P%�=@�!�d�(S/���T�XIv։�q	p�!�PA���5�,V^�-�d(�.Z�!��G��P�t�L�JK�5H�5<�!���d�w�}W�TA�aX
u�!��,���
�#F/g@�Q:6�_G!�$W��"��A-��s���;G�!�*���(7熃,r�<QnR:�!�WY�����N�8h|\գ7�>YG!��	Ħ��@�[���+���Y!�$��!
`4RS!��[B�����X�!��u,��jǽM���"f팅#�!�d	^6�<�a�@�`�;s�(+�!��
+Μ�"�_-8V����	�(�!�$C7*XZ�e��-	p	�эݡk|!�$��@��j
�,;0-Jti!�M�x���փ$|���=|!�dB�4�t�@)�He��&Z�6�!��֭\hT�%���Y�-Q�nʩ5�!�$ϳ]
�Z�з�.���U�!�D�;ef�����$8d J05+!�D�+��}1� �'II��CB�o�!�D��<٪ �E� 2\H��n�iD!�d@3��I�^j�]"���Z@!�`3�H#0�؎�̢�FK
yhB�I�&e��
�.�H��K�ƅt�~B��C�f�G,q�à
DX[�B�,8{*P�R$��M0�e�r+xB�	�z�$�A�K�F�}��e['EVB�)� N���H�:��h������"O��)�-���6�Hg��	n��T�P"O�9A�HN
�u3��ݬD¤	b""OTA�@��-hb:���K�X����B"O��qG��:�R�h��b��	�R"O0�`C�؛*��1�8V�,�W"O<\� d����B$��zF��a�"O�]�f��S�l�9�A-Hu95"O��褢�.�(���F�Li�"OBura']4���=��M��"O�f,X�6�Blr��P�G�|-��"O lYW��4� ��|Ժ�ѧ"O4����o62�Sd���M t"O�5����5�@�)qi���~|�D"OL}A�n�EHƅ2E�F.*��u�"O8$�Ƥ�-���ɶg5C� ��"O$�82'�.L x@iB ��Q�"O���g���BUʂ(ƅ_����"O��RKe�`乲�Lgj��z�"ON�����2X��+�	E<Upp�"O�q��`��}�tW�qq�ѹ"O&I{����_��-��G͠jEb�	�"O����I!~�1w�V
�"P"O����,�5�Fn�]E"O��q��>i�*�X�o:]:n�K�"O���2�ڤ+�}y�i�*R�*�"O�� P��e�(�JG4�@=��"O�S��̰ Fh*R'^<E���E"O�}�ǯ�}�fb&a� ���2"O$�9�kR�0�Z��Q�_M�X�@U"O�4��/7GT=����`}(�c�"O�(��o�A��M%KӶ�y�"O��'�� ���Gɱ%s���"O½ࢊB�/�`F^�I�.�!�"O:���AڢP 9:�NC/6���@c"O�0�ͅ�-��(	�-�U%��1�"O���5.�H1�����QD"O ��EK?=�&Uj#�G|���Sa"O�� $8E̪����4�9�"O8�)u㊕y��ࣰ�I��.�D"O8]@�݌Oa�ͪ���A�>�K�"O*����L�?��1&K�q���`�"OR�@�Ӳ+�0)`s]�!�"O*؃֚S�U���?I�$�s%"O���7 D)9"�|زe��|�&ك"O��bC$T.XQ ��&d���}�6"O��b�e�2wn~lxg"5z�t�h�"OIs��A(%��Q5�N3o��c"OX�AS���r�lXC�NX&H6"OF0D��-�����O����T"O@���a�lo&(�����x��&"O6h�H;���tm�R����"O�Ɇ(ӳ>���DmUf�~���"O��FC݆L�ݘՉ�K:(��"O*�3��H�*j�Z�Iӿq�D��"O�4�5�ʖ\.*I)p�ٰ��L�"OL�їG�F;�Z���\8��"Oԁ����$�<��HF!t�1W"O�1�"R eR8���۠I4���"OB)��ʨ[�0��Nߞn���qP"Oα#��
|���3�-ܢa�XrP"O¼��kP,�-��ٖ!h�BR"Odts!�R���,Ʌ�� ��i""Ot���>j�^���U��)��"O� ��hǄG�`	⣣��Q\�{@"OT��K:����@�ĳ/C��"5"O:��i��"ul�ː��+p B�"O0���K���1Unȭ4i��"O�K&&��+���آ8 -��Xs"O(����A
9{Z�B�@�r yI�"Oh�[�Z[Bp!a(�?C-4!�"OzI�!��8��+3.˱:�H�S`"O"-	��.�* ��N�n�2�"O��E��?��T�SȀ�,�`"O��qCg�-���`�F�VL�"O0ui`�T��d�J���+�☰"O|�	E��"H�:P��'
?k��9��"O0��! �,bx���f�>�9�P"O��:sOQ���$V"s�D�"O�)*�$_�2 $yQC.����"O�	�v)؆r6��C�R�u�X��"O^��S�β%p�:Go
)$w�s!"OF����:@��1�R��]ї"O*7�8(l���En֋oΝ &�#D�4��gΨH��� �T%>< �Y��#D�8a&F�7d�D�4+��'���5�4D���#*�#qo���H�3@��x�3D�̹�)7<�`,�h64�|aiw�1D���I� %���ĤslAS��/D�\��(̄I��I#�n�wN����-D�4	���c'�#aFB�f�$���,D��Qr�M)�F�7f߸$;�X��+D��GJ�"%ZDx�E$��rA�Љ�e(D���SF�D".ɰ�D�l܊5��� D��O>,�ƝXC��:�x���*D��pCLS�hz%��I�mV<ͣE�<D������	��b�/�4}��<D��37ɂ�HT�� T:��%���8D����׍Y\�m��hΚ8��9P%h8D��s�(��A��p��Acg6D�d��
�����5&��5
:D���w�͙��I�a	��t�U�E�;D��@ԫ->���7'�qb�IZ�%'D��CǏھ!�(i��ɢ/�}:/&D�\��ꕝI_(�*�j��#@VB䉏D���rFK�$��90ϔ�+�B�	�J���� `�	'P�4j��H�C�I%K~��F��:d��G�Y3�B�	'X���m*A��j�|C�I�#q$UZb�W�}&�1	�&��<ZC�	�ob2Px�خv�5���E`�C�I�E.p�yV��&_h��Y��B��4C�I�@�j��\�FN���_�r3C�I�ަ��7�Zl�t�Ŝ1F��B�	�\X6|`��N$Z�dز ��K�B�.h�4:��Z�{�zl�E�[���B�V졻�O 4�HT�b��N��B䉔�@0����7M�:t�w�V�MڄB䉬��f!�Be�?y)L�Aq*O�͚O�!�qisD|���"O��Pa�Q�����U.ظj�A��"O� �� �/EҰ�%C߄J�!�!"OJ��(ٕSR�5ءaF��h�"OVY�b�ϡ}�n���@�$��(�"O�%�Ң��\��p�!7Q�<��r"Ot�h�ܥA�H���;q �8�D"Ohĩ$"�3��!�C����'�qO��/C&"�X�rI��1��A("O�  �(���m����2���`��'�L��'�b�٥(�A�����C5�=Y�'�9�5O.���H�9�|*��d'�S�Dʓ�]\&d����A��h���y�#S��9�TZp�� �T�/q�<���O�(�-Oe������n�H���I ����!�[3Q9�Ţ0�׌�b��Y�hc
�1�2�4��=[��2@�)+y����Ñ��'}}�'|��#H$T]��S����z���H�'�&-�\��؋&q�Ɓ��OTY��O(�	j�Ӻ;�O��36+�3I�h�b戅�3_l�[�'��U�s���hy�!x2œ!F������'�ґ|"P����ʑ!G0|�D
U�SaRh�cVh�<���E3'�$){��&~��x�b�Za�<� �&�,����׼cK\Ը��Z[�<��Ƃj7�T2���yl� �,�Y�<i�E¥BP��Q��8I����eY�<)"�ҰV�2u���\</�B���S�<aL�%����9i��;ui�P�<�f�dl�Q�v�̭8�:a�$!�$�	O�$aA���T����)��k�!�DK`I� o]�h�V�2!�!��˲=�R��Gtԅ�s�\�j/D8��hO?M��9N�$�H�BѧMڢ��U�#D�p	�Ƕj�� �φk��$�!b7D�D
�gH-�y$���G2����*D��e$Եv0V���@C�sh�ʷI)D��Ĥ[�3��(�fj�L�d$�s%%D�p�  ��sž���6M�b�r��5D�H�s�*�`*��b  �))4D��ҐD؟+|���ߞ=�
 Ò�p�E{�����pB� E�:�Ą%-!�D}���c�ϥ9��y��IݪW!��(h��d�3�&��&��N!�d�6jB>�$�&j���0���n�!���g
�51���,�rf��X�!� ���ۦ�L(x(ٛ �ΏC�!�Ԕ|�i�筇h�����,^�	s��0<�I_ʺ1Pd%	�@
��$k�<�% �/\ph�3G�H�U�0R�e
릑���/�T�d�J��N�Ť=cBiF#C�ZP��6�q��VP��G&էg�D�'��~�#w��IF��^~�p��Y��d5�S�O,�A�BG n�&��B�L�a��Ep�'��+�ߓ<6�|	����T5����>Y��	��t|p��PdY>Ti�V*�	F�!�&�>,��gڟ�Kѣ:��p�ݴ���1���O�@A#��a� !��Ȋ2�nM�'F$ы���1�����gH-0A�xS�'�д��	
��uA�`ԛ'�LJN>����~��tR	�0,U(H����ȕ�y;<\�� �K�j����RKD��R��<a�O�ܣϓp��@gٖ���9��$Yݴ��=t��ifjݝ_"�-H�	�yr�Gx"�'���X���1���ׂ!H��4���d>��UeC-Iش8O^3	�(�0Pa6}b�'SP�zg��G���ж�M�C�f�9��?	��:1�ѡp��5ͺ�Q�g��k�!�_�z���j�$�@`�4p6�N�+�ٟ�'��;�Oq�
$z�H�]��dCr$P�M��=A�"O����♎>��<k&�0,��,;"��3LO��x�
�+I}H�Sdl�(%l�q��"OL�l@�Q�dЧ�U�`ܩ�g]���I�G��ʁ���fL(�Jː*��C�)� vh���ùl�����Yk��	tX��Y��[7D(�(&m-YV8��.��1�O�� -a��� qo�; V)0! $�\�f�E�^��p��Q�H�Kc&�z��D�?�e$څ|^x�K#��2�4ъ��L�<�#�U;]l��@E�,Z�D4Z��dΓ�M�O>E���d���B��H�&�2���J��'�H��?�͟��J8jYP�dj2
M��֞~���'��&�'���3k�u�q
�͉���a��>�e*�>�N|n�?'v�,Sp�)!�U�ƍ��l����ēMj�H���؀"N@@(�nLE���Ml��u�=q��T?��r��.�
|�&g�g7�A�:�c6�I��P�p�圜`��xT����84�x��)�S�9�ؙb���-�`���	��b@>O���۴�ا�O���t��0e�`�+�23+�y�O����5**PK����Z8�D~�Gx2-�'�?��w���d�ЀII�58�Bʇ:��ȓ�6�8����+�@D���T�����p��>	��3�f�r��AM�Q9D$����
���ȓj�Z�q3�
�;fE�p��_	�@��O���G�*�(Hb�/Z��O��@u�u!(�21��/����Pe3D�L�� ʗs��yu	��P"��#0D����P��8p`j��a��� /D�dY���Zc��` �]&t���XAM+��6�SܧVJq13��};�B��5A\Xԇ�A�&	��d
��J�ふ�(�Gzr��d�O-��i"���x��2�@83�4��'2F1÷Q�h�x��B�G��4ճ
�':*��'��,}z�;�A]�t�މ�	�'��U�T-S�$�z��T�6Mq��'�p��K;3�Vp�қ@�^5��'����%�ʢb*�<�D�)@�f�8�'ˮ��D��i�z923 �iD�Q�O���$߉j�X���l��&�.�Ԡ,�y$��asCnJ57��Yc!��~R�)�'n:T�b�J"�� S�ɫb�BL��ID�k����D�Eh	�eXe�$(\(�ȓF���c�<A7X��`�Y�"�����hO���`I�/ԨxS��������T��DR���'�(��`�پJ��5#�;6 8��'� �C�Tٜ}:E�92.`x�'�*��1ڬW߆0����[�s�'��,	�)��p�왻������0>�N>!WG!�H�3��	W�F�zg��<�'�Ă�-��؆C�8��S�Oq}g?��(�9$P�-4��R�S/0�����"OP����L�o�D�������'��<�	�O�8{��H�cG���Fįw���/LO"�`�ׄJ�[����&�@px�� ��>1��-�b��$'��3��C�&T�J����8b�H���$(=��ښm�TXb"O���QMX)?�`�6nC�U�ݐ���d�ڃ��D�$@q�%Ŏ8`�Ҍ�S�<�6`�F�8A�_�$H�-�t��<Q���6{�Ѣ��
2R~xx6NO'��c��D{����P"a<8���?�$������y¯�+a�� V���r�|�"&���y��/qGF��'X:w���!gk�%�y҂�q~���T�E^F8;�N[�yr  ���3�IF�T��X٦ ���y�!H��#*�Gk�A��V�yr+45P��"@L�.D201)5g��y�̖�r��a����>%"T(J�7�y
� ���#�uZT�ħߡQ�����"Ox]9�D��b�C�ĝ-F���""O�Ȉ�,���1���N4Xa6"O���dl?��(d�9�1H!"Ot�S�Q�:��eH1�P�U���"O��y!(A�4����0�-\�r��"O�����k��P��B��zG"O^�S KF�Uw��KDIQ�?� Y"O���G0�[Ղ^��ڰp1"O:��ЯJ�j�`�Ȅ� :��՛�"O2e*@�B�\ܰK<�fl�S"O�]��!W�/�0��-ʭ0��<�"OACU�^m�Hs$���1���"O���U
Ĳ+H$A!�ю� "O�e�"���DIpӬ��VÎ��u"O�]��'�:F�nX)�+P�nI�"O$r���j��݊�)|����"O����:��H�$�)cy� '"O�b��E/4%̽�6I5p
�"O���Dbϧtd\*���5@���"OB�K���?A4ؐtȮh*�At"O�$��˩Gz&�j���v� "O.%ఊ��l�\���j!�i'"O
�§�˘24v,�hF�r�us�"OD`�
�z�`�f�C�~�xV"O���'f�.�0hӲ�&O����"O��6���e� R�-=��B0�J�<��
H:`�h�@�pN���G�MC�<��@N�?C�$�I� 3Zt�v�XZ�<�#D�>?~��*�o�1��bX̓`��s��;M
���=w�t�<)U�S "B���^�xTx�Z
Q�<����G���-�#
U���T��O�<Qテ&ݺ�`��5����f�@�<a����Ҍ��Ѵvʍ���@�<� ��&�{Ӈ� <�āp�<���Y�B5���׳*V�e�3-�v�<�v���p攕P�Ƃ�wvL�ѩ�K�<13 �/m"&P��NZn�! fN�<id���Ԥ�>p6�Q�VR�<A��9 �:��\�2�����K�R�<�t�Z� �����y�6u�4�QM�<�C��T��K��K���{S%�f�<�d��P�R���Ki081[P�Vg�<��E(\��}�D��tJ<3���D�<����$$ �X�B��r �A�<��N$(��SpC�P�� �`�Yj�<�
ߣ(Y�@��@�
�y�g@e�<A���VTllá���r�J�a�+�a�<�剓>;W����Ȟq�l@��"D��3����$�3��pVp���!'D��3`ڕN��r��Ȉ	�Ppq �%D��W"Ҭ	�n<����TB�r��%D�Hy�o��#ΚQbpmF��v��M/D��"�%K!Q�TZCÙl�^ҁ�0D���Ug�m��� A+{B"�.D���Ɠ	2m���9o~	�I/D��F�V�H	���� 	Ap;F�-D�$��+D�g1|�q����&�[��*D��������Ul�#m7ܬ!��*D�[TQ/X����.߳2��J��(D����혋u�8ys4�V��`�A2D�0$b��+]�a��h�H��ԛC�0D����(=7�yc���7IJL��0D��`��w#�1�u��.P��D�,D�� ����C�%8tY����L^�iv"O��C��Q���� ��_�`�( "O�)٤�&S:�q�`�4	���"OR䠳�!�Ψ*D�*���H°iv0#�'��	rC_�cd�rǋ�\�Lu�(���2a7?�s,[�xAXݑ�GК~Dp�+��Vz�<�!!Ö9:�<��	v �+��X�
��9�c,��A&�M5.��TrA�;u�=�"O�TQ��]H3��b�!�I�"81�䈗V�qO��#��Y���DNݫ}��"�$�)ۨah�M2D��ۆ�M8l�fbt�+l^�X�>lȨ��6�O���*� __�D3SiR�m���'��H�da�A~��G�<z�Z��O�tP�'�Q���x��-��!��l��	��a+�+f��Z�x�FV�cU�O�On��b,I.A0v�v�T�# �9#
˓]�n�S�.���|"�  !(�b�P��R��'!�$]-���@n��1�a�F��%���VhZ�[6qO�����"GƷp�`<J��m�PE�V"O�(�b��Ey��FI;d�%"�,�	��-)��L<�Q�H5>��k֮�$�f4(7��vH<9"-?ԨhI��M,Uba��E�9ɖ܃0�*�O>��d�_U�`	���R$���Q�'�D�*�K�M�I �j��aD<1U!�$�!XhDC�	�2�\u`a̞��l��
�&��O�`��J?�)�(R\�6��[�M����P+B�	6Zժ�L��A򋝷V�B�I�^�F�ߺh���5↔r��C�I����b�S��";}�C�7s!L咒(d���N�(�C�IKe0�KV��0c8t8׃�G��C�	8��{@A�� ��@���C�5kh�Iq�
6�8Y�	,A�JC�bX�{'D��q��ATIG�#-.C��ol:8P&l�j����BB�I�n����ٱ��	��ЂS.bB�7�P\[�J�1y��ce �׊C�	�H�]0�Q�9!H1�Ԃ�Yo`C�	�.�o�;FR\mKB��e)RC�	<�h�aԈ̕e�\�8dmA�(C�	�7�\̺r��t>���� ��B�I�9a���ҥѤ|�{b�"'�B�IC�b1�FG�-OX�������4�⣓�5��?M{a�`y�,�7��5�|]��"D�Db�(����Fه"x��`_��ؠ0�|rO?�g}2g+4J�D��?K񌽠'�,�y�]�)��񨧭YA��L�fD�ڽ���yܐm ��N��0=ɳM.^��e�Ee�"~}�|�0�Fpy�-��T�����|ZwV^5�wO�`��ͮ5�4�i���+ ����'�҃0�P�'��t(�"E�k��+�/��h�!���01V ��%����X��T�8'�b�qq�]�<&�=A<��v��S�	��/F�9/a|Х|3�Q!'^�_Z�)�E�]{
	ӧ�Z�t��Ј �T&UP��2~_��a��JXT��e�~�B�x"E9z�r�3gۿeI2�6��э,��ں��<I3ޱ�'�^�&��i���	�@�	?q�&iʠ$S�R2TԠ`-F�s7�$@*�K����<)��3c�D�%/ "D2���	�0��%&n�5[�*1B�d�Z����3a�l��/�!&N&�ɵi5��%s�?����u�ˢS8V�(�*��u|R��Y��(2�7u
��T,��t�D�Zӫ�u�RLXs� /L��1��E�6���׈�4r��,͐r�L�3ًs�@\`s� /q���2��G���4bU��#x����D�~��@N�|�BE����JJ,���jg��qPR���v�m��D�;��0��"H\r'Ϛ&KL.����	�g����ٓ�I�a�ҹ�N�*V���8$FX%�c��9&�:n��zg9�L����?E�D�Q�e{HQ���_�,�#�$\2�y#6g��:ޕ�%o�?F�|�UcX�cw\M��A^� �sԛxr�'��lذ%�"k�n��&�J�Z J@2 �]�1���:k�<��'��L�e� h�j��<+�n�1��Af ��VH��Ni�b�	Yol�(4��o���)�$ΐ��,3L�"ׁg��,�PC[�_���2��)ql0&H	�7�����*,1B�B�A�g��,l6� |��FQ
>ԙ�'�Qf�P�=]�6y��]x��@R�^�^�:m����؀ �	Sd>�6	�B%B�h�|t�B ��1D���h2-^0doZ�[蓦ɾ5z}
&�
�o�\��0� �?qX#V;M
R�4.
	p1�� ��!�r��fl�Ojf�j�'��nEr���n_>GAP�I���)ts���D�y�ըH+0/2�
�n� ���.?DF^��'1.h
�m	2*�W,�/.�LM���Q��0�B����铄5$|"�k�W.*Xh�#�!_d�5	W��	���Ae�1*)���]�s ���o���k� �6��j���%���'�Zh���]��)�'�)�^�n�;,�=nG��AS�V3{]���G�-��	�d��k�(a��pE����i�&}��含mV��OI/|�d�4F2a�� B�0}r	��f�Ʊ[�D�}����o��1�8�P��vܬE0wBΩ��yK1�	�5(4�����rڤM�~J�G[�X�`0
��S�G;�Z4�̌@p���%� G�.�P�C� D����Ox����<���&��ƍ�9�z	�Ѩ��[�������+ݹB�:&`[*t嘨��g�-U�ԍC� ��f	��"���-��J��'�X��w�@-V}�%��5ΆP�'`%(p
ʌ/%��Y�>Ap�T�XZD1LI�P�H���L��\1��y�G���(��2k�I�b���5���E�S��~	���Qي��c��1���A��ӱ��bL-a�¥f9f�R�9~��>`�gّtVdk7H?7*�x*��/ʓS��80g'X�|Zt{���o	n�r�@#@�}��,��G�"��L��.�
0
t�WoO�z�D�𙟜��F_�xE3Ŝ�ed��"�)h�=Y�n��PWƑP.O?��Ӓ=�1{�!K�?Ḅ�gMZ:)a�#_��8�s��}�d�5��U0@��a�C��6 ��)�J�>���X�\� �l!�	�]�(���9T��z��0az�pV�H5X�|�`g�-��(3�'W�Y�b��3b���a϶~/5�U�Z$6�����V�zt`����8�� ��׭dl�ȰgG�|��&��p�N��T���x�@A$Vu�<YW�-F��IP�I���@
u�j��R0e�,AQ)xO�pl�����y���Z�:��+�(�DA�����y".�Sa,���
�UG�������j䜰	e&+R��`h���a�Ƀ��T��E��f.����&�?h�bxc�6A��~�2K��pA���q�"R��X6�,�B+�u�<r�UZ
a{�<20&Yڔ-�+h���ܩ��O♡ai��n�B@����x�ZIZa��������
�$�g:H)�"O�=��(�"��s��nz� Z�<��bL�2�Y��`�mCr1����G=ꌺ`�B$*L,���C7JrB��*@*z�(�a&��UJ��@=0�b ��A�.O����Y��xgOٽ:�,؛a��� �:�Z��%D���$M
��s��?��0� a�qՔm�@�=����,`�vKƶjWh!��Ľq:���C�4���@lڗH̙���ne�<uK&eJjB��/$�2��& \�̌L��M��-Lc�h��K�G����@���4x���_5���A!�z��C�I%^ <d�͌7
�Ip g�%+�R]�%��&k�ΒOP�}�j<�c�lΩ�8`A�DN:oq@����Li�f�U.,*�q��;G�*�ȓ"�(@�@)-�̵H�FF2|jnu�ȓ � qU�
M��w�W� ����ȓ���Z`�zAZ,���1>�\��O�T qO,�}��l���*cx^��]�TI>�ȓx�%9��8�J�#�O�<+��n�%�
`�B�i8�P��D�a���-��A	��25b6\O�ac���}�F���'��b���1$�������Y8���'A��9��_�x�噲��َ�!�{"LɀhM�8J�MA�O� �`��;Uz�2 *�� �'�����Jҷ)]�F�ζ!����e8�*i�J�����<P��̆KT%^,B� ���i�<��NI�kw,�8򌒠c?~�  j�X�'S�&�"��(��(�&�ްDA0� `V���A�RM�Z �E��y���in�9`�W?R~��0��N��yU�?�.J��L-��K����'����Ņ<�b�E���!���(�/�F�Z-�pjS6�y2� K�n}�a�Ō0Qh�{Gǉ�rL��OV7���b�Q>�|�����b����;Q��хȓ~�����kd�P��1'�Z�mZ�bҚ�K�!�L8��b%�\�i� i�BJߎ�S ,|O"�ԭ������=ZsV��`�ζJ�	��}k!�d�5^1��Ǉ�q�M� *K"o!�� �8"��U+�RQ��r�n�3"O��� �5�TXJ%�M.0�8bC"O&�A3e�S^J	*�͕�-���S"O��FG�|�3%0�*�ѥ"O6� �j�!�`�wn��@�@"O0�z�o�;�] ��� i����"OJ�X�lO�/J8T��� ��L�T"O�dK`(^K�t}��Ͼ4��,��"O�Q��S�Fs��9��5�V�а"OT	�����ĈF��0�d�"O:U��_Nj-���y�4���"O&���N�M��V䍐C��-j�"O��JW�Gk2�9FYAR6��S"O*D��5p��	�@Kj(��"O��z�ƀ>"B�����"*TC1"O*x�
*D4�i��3"�|<��"O�a7���x�ɑ*Dd�:�*!"O�-(�k�&(���Y��w��l��"O�l�f��&(C℀7G�&�\)� "O|\h�#�b��� ,�|+&"O ��2,�7!S���
��8|�1"O���`�1-^޸J��d����"O��� ߁N��E���>��Ԓ�"Ob��c��CN^YH坫Y@�i�"O��@"�c��l�Cˏ�G��\��"O�Lv*K<){��Y���8�����"OL]�]�n5
��掹1����"O�ܢ�4�b�H���!G�����"O��H����>�NE���7BK�؀�"Oh�Q�.���d�aOF)S�m(�"O^)bU�N WVX�2��	onµ{�"O$9�7�O�J�}f�8]f	i�"O�ap�cL�5��H7gԓH�B�H�"O�%#�H�>L��Q�2)P��|�{"O*�9�+�~�ڐ+R�Nº��R"O�pF)f�ȸ�/�@�|��"O��3�R1+#1S�v�K�"O�U1pBD�FW�d���N�bx�|s�"OK���=�ѠD�ie���"O��h��O���H�U@^@����"O�dH�`ћr��lbA�N=v�\�Q�"O:�r.W�����H�;�J��"O�D���i�@�cMW�>���Q#"Oƨh� ��~:­��L�>�4��"O�Vdݫ)%��j�?V|�S�"OR�q���G��H��
zf"Ovq3"��	�,�+bi��ڂ"O������7>|�*&���`�"O�9�5�`a�	9\�:��iW� !�ě�B�f��eG��.���v���#-!���)��@�C$Y�ڕ���7!��H�����>d"YC�o͚C1!�$��6]H���JW#F���ڝc\!�@�GU>x�qo��k]>p(��!�ą+,|<�b��:Ui��+�N5)�!�䄔��ɡ`�V=,��-ΚE�!���4w�xCV���b�LqslƎ&�!���}5�����t����Gh�!�$ܷ\�Б�tȄHF�D����`!���Mt k�A�H7���u�!�D�n��ʓ)�<@֕c�c�: �!�� �2	��)F�i�*��0���!򤍴�Yy�N^�^�H�[��Ȩy�!�$V3*0��b��D&�E2�(�6nS!�� ��!��-�.� ��ڂ\K�"O�(��	�V��2	��d�s"On�� ��|����3��6~����"O\d��i�N�hr�$d����"OԹ�>�� s�D�0S��"Ov,(ԧS+eu��j"�W	�0���"O��#S��Y��$�#A+5��#�"O��	Fa��X�ZY�'"O���r�"O�x@�Ì�;�T8��8Eyv)�a"OT���Ɔ:-)�n��;f�4�"O��ycj�9	���.�����"O4�+�C�y%چF�X�.�:F"O�p�r��|碥��o�7�$���"O�H0P�Z<�#X�4��䁡"O�Ly�Díw�n�����6��M�"O ���Y�S:�l�˾���"On�1���� QJČ)(�^�p!"O�H(��2" tԘԬ��+��\�"O6<Q��¸�u�2��%�>�"O}[�a@2z��P��	�/K�*��"O�m����g�X�4�
"{��IZ�"O胣�ѦO��5`�ۖ>�<Y�"OX��pR�e����	��LUc"O�9�#�X�%j��G�3�N��r"O
q	E�G�A���# P & �"O����➖@B�q	���
	���"Ov�3��F9�~,�A&�
�i��"O�`:�[�,c��S�/L�u�T��"O�L)�E����Ϙ��{4"O��G.�)^����qM�:\��"O�5�vFF��0��NR$��"O�IPӌلPUً�ʄ"!���"OJ��6%��M�|��B�_���Z3"OT8��Mdܰ��s�ǲ-s2�R�"O��˛/@��ї�_�
KDd
�"O(|4��0�G�U4;�X�g�<1g�"S�H2˂7�l�pl\�<��ŝE��3��KM�T�
���f�<1���dk��g>1kr\�u�FH�<��
De�t��";�b����p�<ADf�5QVLK��`� ��͟r�<1����z	jE�PH�$��Ēw�<Ib�Q���X�&%��+�F�h�e�<��G3q�h�pD:$�^L��-x�<�7��!_�$�U+I*[����⇂u�<��l�ր���ռl�d�f��l�L�h�ō9�'| ���<�TiAN�',!^��Z�a�U�%��1�	\f�v}Ұ+�^�OtuF��O�q��o4;pp)`����jr"O��z��Q/*��ڴ�K�%�V�&�ɨ&���Т��L���K�'�0���>Ro���V�D̴.OJ��f�9N`�O�ۙk���L�c�:	��\*2����FH��X��QЫ��dP��d
��Hg�ղy�c�\;y�$�"%�}�Ƈ�:r��e�"��&�+r�Z�my��Cg�x�}X�-9x��e�C"��`Ä-9�O9x�G�&m�20�f��p@B��*X� r@$�Āԗt� QI�$�O���JB�DI	BiaWJsEF�O!�O�𱳩� |���ǇZ?Z�Z��R���#�SD�$I�O���hM8��P@��9zNu�5f� {MA��h�7(���'��&Xo�=�$�DX�4�F�^3:���C��Rj��
n��)��-�g1�hI�AƐyШ��^29��IV���W~8���k���¥�X�D�<!�BB�j�j!I/]k���ȗ��IqƇ�2�@��v+G��t)�N�btVCp��)k�`h�����Yq�1 �T���F�
�k��Ұ u�˹k�HR�.ٕz�����'H�9�r��7�V��j�&(�ja�!R�Rd��#b:vH���t6=��Tf�23���Ľ?��R�Y~�U�UP�}P����,*s@^���'�� ��FB�R�Za�Wq8R���O��:v��($�]�U��?64ɱ��јoӠ���Q]Ǭ�S3�-3����� ��9�NU%:�"�3����$,~%��*L��L}�S��0*�z���9�����$>�6�s�BA���N*6{P�+"+�'�VD�`��(�I��酊'�(q���zǼ��ثD��ث��E�6���w��?h���
�H=;�^tP�I�zŲ��FX�D�����)4���R���c�Z]t��;0�o	�x�퉹x����lC��9jDHEdH1py�m����9-i��s�F�WL�<S�޶t�Â6O��x�*��X,P��WM8�۰-�{Հ4�?	P/Z$ ,�P��i���̘c�	��E�
�f�L�1r�"���~B @7Xa| ��k�U�hᠯ�V� �3!�2A���������0p%J �9��S�O=�x��	�uZ�BS&ػc�Ų��ƃ~tlPJǰij�cW�\�ZU���� 	��h`@�$�d�����d,�	6f4Yu�F}�	28�!�i5�|X�'���X���6>6�p��"d�r�	��p>ch]�'�0�I�m�iR�h2�S�?:,t��Y"Ym�Q��}���n�U�M	���[$e��1xx�H�뇻{��k��I�D�9�%�5~p��~Z�)@�Q0��-.s7����gګ�1�E҉}ڼ�槈��䓄9�ƕ9`��v������7p>A��,]�:01J�y���'��fL�A��@�D��gΜM��'�کC4O�&B�Uc�L2�Keg��JC";��˗�Vp�:2|z�!�W�0P�}�@) ��"��y�f	Y�hL=e��[sM,`��I6|O5����.�|!a'm�A���c��> ��lXՠR�&�R�\���M����GB#��O�2�a�&7z��p�D�X��q��$�$�&�1bf5y��b?�0�ժe�9�Ӫj�:�e��z�L �0 �lj�G}���iY���� �),�p�*��y�f��
)\	���2A��M� �S��?q���֩���"�N}�aO�Z�$��F<J��v��0<9���&��&GڄLtL�*�DR}�GƱ;�,p�#�i�'M�=iaA��7��Q�Ϸ!,ԃun�*���(c@�y�����/�3����gEi=I)v�д{��0�3+
l�'}\����g�E��H�<����'%#� �H[%r�0�C�^��P������mڇm��I��@�1��t�o�0D���������
]��F�d@D� ݶi�6�A�-�H]+�Mг�y�L�a��� /�h]��)��w�
���'<�����W�]�N�PO?��>�F獏'�4Ec��;+{��2 %�]��LY#��49 I�#I����{@,�*���Z �Ѕ8��(��ڽ�*ń�	2�6�i��:0��"�b{d"?��i�"Y.ؑ�_<< �S#�ٺ#u
��?�v�]��\����P�<�b��N�*ĺ�k���BiOy���6R��#�#
&R0���|�OӴ+g��0Y-�ɲr!+@�xc�<�S�^)Q(�k� �>�2��ݨ=Y���<db�u�Q>�X�.� 	o�.�@�EQ4�p�ȓVݔ%��e�=4��@��#Ŷ�0h��ٳhW��#ꋅi<a{��;CL\Ѵ�W9<��a"֤�9�p=�u��9t��)�.п�MCu
�����(^�l�lK��p�<��
*^0i�C�74*\Kb�Pl�WŚLD+S*�z�}�����r�L��W�e���"Rf�<�c��q�r��3Kψ0�F�`� A ?4�x	goN�	`��~�ւ2�-Z���
+�F�7�y"5{ �u!Ӹe߼���O=�y��Ԟ=�T�pf@�f���)� �0�y�	Ԕl�`8p�;_Q�墁��y)S�,��іo?R��`���;~�6���?�I��~"o��|nmK�愂���BW�y"��H4�t/�7@�9�ɉ��M[#�Ad��Y�)m����F�%8�!��q��=��	Oy������!~��ی����S�	Y �{G��O�!�-z-� �m4<,V�N�9�qO�gQCld�{����QN�����
mk��V�&!�d���`*$a�f�(�[0�:zS2��Qa�'@�u�|�'7�rt��-�\�K�Ϙ��C
�'N�LY����{t<��=n(�(��VQ�5��ǁ2�0>Q����,��A�%G_	e���W��Q����'����I�S4ON|���@�\hqa�/ѯl�J��"O*|g�>�"���A�6s�d�w�$�8F�l���!�9����:�	��,x�®^φA�G#!D��+EL@���P�:0~��#��8Q�
L�J>}b�x����Y�)����a�ԝR>�y&�ÓV�!�� �Y"�F)a�t(�w�;i��iE&� u�$��|"��"u���F'�H��A˒��=�d*Xu�.��t��g 
��9��!�4I����ȓ�(}���s"r۳KN/T����8b`��o5hY*����]9�݇ȓv
U� ˠ/'�����s\���Ny�غ�Gܪz���;e�<RU^��t�BDQ���""~��`C�' cN���x3�\IB�
�u�n|���c�|���9�j� �❍v)\��H���ȓ,��]�p��7�l�� �F	�ȓ|��h�ML:=D��Å�j� �� ���r��z�J�@P�
W����D���� �	q"���վY�bD��S{Jx��,�Q�h�G���ȓ5P���j�*mzI�	�"mqn�ȓ2�1q��߶?�P\S��"z�dI�ȓL���Q�R�waɲ��X�EGh��ȓ�4���ѓz :�b�bT�^��_�t4�b%ATb�E���,4*�X���F���R �x��ce�,���Y�'���xT�ΚS��5�A�(�
�'��J�V3_G
��
ݦ2�� 	�'���蔣�jd��� -��+�'����qf��T�B" �/ ��	�'��X�B�3}g�9*������
�'�d}����i�<�Ï�;e`�Q
�'zq�r�Yj��8aF��zʌ	�'��Q�A �E>fa��EN�D��'�����L�\����ň>��9��'�<�y7Jʹ
ă�҆ �a	�']�`�פܛo.��УK*��3	�'|p��9�n �S,��w<�0�'�A���&[��3dS�����'o�AhG����\jqkW�p_d���'�8�)�扎p���PNޫsh49"�'�p���le�� �a�l�@Z�'?���+c`8ya!�0}�lLَy��O�z�rp��ϋ�<�A�fR���'Z��Q�|,�i !�7r��Y�'��ᢢJ.j�<��R	p����'zh��e�G��\=*R�����'�D���#p�+��J�4ƐH�'�dEz���Ta�Tb���g	F��'*�s҉[�a����v��'t�*);�'��Z׬��m�b���ɲ_�$<i�'�����;u@��"1e�Q�4���'H��BP�{�$+��V
Ji�MH�'�D	 'P� ��!�劆��x��'��"=E�@C�4f�0��>�
t!���gg6�Bs�Ocy¥�6#�����-KE|�ʣ�އ13L�X���{�xݺDT���q
�
�����O�8�ZF�?Q2��K〉\�����'I���1��M.���]U>�YR��	3�ݹ&�K�%ņ90���%��� ÝkC�|��)�q��b:`�8�d�m�����^�~m�%(�#�CJ��h�����������,k��Y!֬ɉ,
�T`��>�R�X�=�����/,r�9���4NҪa��'��	�h��Q�6,�)���5����g�I!B���t�:qp��+~W�*��<�)�'h��mA�6v�6Q�$mR�z�J��ȓW��@��3"�d\��������ȓ��0lɂp�V���ٍ �5�ȓN>�ٛ�
R�
,+�hJ�(5GzR�'�tӥ��?� �E	[�yg��'v ��`J�	�.����Hz��xp�'� 4a�f�4��`(�A�'r�ٹ�'�lKd���#6����HПǪ�	��� r��l�`"�Ѓ�{$�h�"Op<���=J6�0��"k
��R�"OL�4�Ű �l��'�#h
�uRP"O��b�ր �hb��خf����"O��btJŊFX$��C��f���H�"OVec� ߒP��P[��)E��D4"O���D	JMA��K�
�R��8"O�	���GT4:u��F}ϊ���"O8��@#�&�VI����&dv"O��
��'�貴�D�+�P���"Oh\9�jCb��5��G#<::���"OZ �c�]�0Q��fi� " -	u"O�	A'f�$-{E�ԑX�A"O$� Fē:�A��Q�`��Չ"OL�c�A�T̀� ��.;��۔"O�u���� ��4�0C{X}��"OS�&*^�P��"Ɓ.Xx�"O浑B`�2_�,�+���Ie4���"O�R��k%�ͱ��P';O�p��"O |�jIx���A>=��W"O:��t��8YÜ<i�l�+U>P���"Ox`�ע��ę�+P�x89�"OV
Q#�x�������"O �D��i���ҷ+�1`~���"OlmS��1}�� ��.p�dV"Ox�����"$����(��6i�d�#"O���&��;@�ذ��GIPf ���"O����@�6I���#���dW�@["O�@�Fd��K^�!��D�3cT||zG"O�x�u ��pz�!�<���R"Oƕ҇bU�~s��"� �O�N�y�"O"������i�/�d�	p"O�h��B|�H��%�HQJ�A"O@u˶j�>�N���7�b8a�"O.�B�&�yV�b#Êh5���"Ox͒���z���*tC�-���S"O `{!���^dꑄ�=>��"O�����#���$cEp.Ƭ�7"OM�È�2p��ⓣ�r�
"O��3��ri�+w�M��D1	�"O�e���P\�V���O�C�蜒b"O=���ڑ�����@]�� �"OF�b�4��������HՑ2"O�!P&"t�$spE>P�|4s�"O�x��iI7[]r�٣������U�!D�t� &?K�{`b\�R$��u�2D���0g�\����Y�k%���2"2D�����4�(d��'V
o�Ыa..D���f��3�-i��8������)D����C�)��mYↅ�.1bQ 'D���&��^ncf��:~if�0��0D�PQj��=�Ed_#f�D�I �.D�\�@E��WGd�w ��oO���+D��R�/N;/[>I��YQ0+D���a���7�ѝ��rPL�Z�<9І�j�����/ra���}�<�ckS=�K���d���fN���C�ə D��:��;MaPE�aI�8��C�	�^s�Sm�(J:Ł�-E�M�C�ɬ&�� ��U3E�R@#�	�D$�C���֐�pmW 2Ft3%��$��B�	%Nm�šd������F�T!�B䉃}��@��Ή|��cP��]L"C�I=3jd�򷫆t�����k�6x1(C�)� ��	�*!�j n+zy�@"Oj��s!� p�5��ְ�T%�Q"O�81파E6b)q�9(�4�kQ"O�-��.ΆZ&LT�}��U�g"O��� '�wj�²����8F"Oք�6�.�*��؜��(C"OԐq�6�yF)zZEС"O��x���!L��J��Z���p"O���p��=&f Adb�w���f"OL���A?:0ha;�c��i{�)�Q"O ��oX�]��<�C��:9�Hy�P"O�|���	O�8�c߾n���yw"O�遥��C�.T�g�Ό>�xf"O`�H�B
39x���H��t��"OX���-�68��B];H^�"O�x�pgC!n�V 	�CʰTiI"O�] GㄚJ����U��i��"O�$��\�c������)���4"O�Qy�!�'I� U���Y]�t`2"O+Í�;C��Dg6����"O
���M�9�,ܐ𭀻�|Hx "O���cD8)¤*���\�T��"O��±j�%b1<�{�j��Mf2��"O�	��i�2gbtY�L�Fk3"O��a�ތ{	�������H�8��b"O��x3+�Rw�L��Z�s~�YX&"O(�seMٖ �B�BaB� %��a��"OR=����,1�K��ŘVX- �"O8T�ՎK%Ny�5��䄨p9<=Z�"O
��ꅰAD4�z��S�+
pa"On(�S�:L����!	8��� 7"O�@�
ɽ7���x���Yf�k"O��藠
6�T��6Ep �"O4�󳮜�JIĸ�w,�+]-&!1�"O�\���\4J_�W�^�#]ó"OB����>/WN�9�,��&x2#A1D�|Js�Îo\`�˗�8a�TX��-D�t��	����d��`��1Z�+D��'N�RA�YАg��T� ˵)*D����T�2��礃�l�����(D��)V�3}�l$��hC x��`E(D����A��r�3�\�#� p��(D�����Q�i�>�k���:�zq)5n%D���1��n���
d�9$���-D�JW������-�H��(���-D����b��y�6᳖��h�hP1�O?D�$)1��2	�zLZcE�!�|Š5(?D����P�e,|��!R�d�zq��=D�t����*q̰c�
�%]��y��<D�|���45����������:D��7A��II�����[$����9D�8;���68u����3:�k5g)D�Y ��t�ְ�¬�<fQ��0�:D�|ɡ��.�t�$M��/���#D��xujɈN4ܫ��[�d��4�R� D�T;e���,c��)���cP�>D��Z�-T� �T�#3XP0�!D�8ٱ�W	�Չr`V�uzu1��1D�xB�F����U�CZ`�Q��3D��r��ڗ>;ne�fL՘GU�YZp�6D��C'O_N� �̔���M0u�0D��;��E*n��Z®ђ���@<D��Y�)���H,P�Q���w.8D����%AB��⨎<ƀ�b�;D�� �̳<����/<0V�\�"OV�$�#�p��͟�NFJ�{"O����{!^�[nY,eǖ�Ce"O��ᢍ0t_���Ae���#u"O��f��
ٞؒ��Uhc^C�"O�]�i�/`��"�HX�,q�m�P"O($�iH�E��y@���>7P��""O�!B#H�W7֍k�aUH�8Qa"O����K4>�
y:��\>���g"O�0q�	{�d�"����+xx�"O�!����jk>y�㘌}�:��"OȘR��tL�"�a��~�쳥"O�Y���[dd�j�a�!=��H�"O�8�6� �S��z���!"��q�"O\q��*�8<[�C�Tv�!!"O�	2�
;��A��c����"O r��.6r���,�>���Z""Oq37�@"zw�}@�j�p�b�S�"O���� �9�.��(��޽��"O�8�2�UWu�`��L�(7٬�j�"O�Y���E�0���O6�^� �"O>��3�M"}�N$��m����"O,)D���xAd���ǂ��"Op���E��W�L�ci��U�p��"ObD�aL�L�z���U F�y�"O�q�K^=pO<���ܲ.��W"O,)Ss�P<_�,Da�7+BM��"O�����4/�:;�տ<�0��A"O�ܺf$OT�S��Y��|�"OX�3*X!�V��EV9,���"Oz|��K�b�� D��X�A��"Ojt��3׶��AB��w"Oz���	T��pA��r� �"OHX� �ʭ6hJp�r���@��:Q"O�]�1�d��u"jv�y�"O��)!�^�q�t�����A"O�(�"D!z��i��C�6��Sa"O��ӇF�#qp��C�̿@�Z�iq"Oΐ@�DT-V���s���4)��̐�"O�M�c�R�?q�(4"��0�(	��"O��R�aĨ&,�X�A��<<����C"O��P��I�m<�[B틏7���T"O�Ԁ�F	�xW:3���[�䨦"O� b�h�1]�|H�l��)t��$"O� 2�'x8�Br����'o�j�<�nKTj1�A'۸'dD@�W�A�<9���:m�e�B��t?�,2Rf�A�<�W�Ʃ-��YIQ
�Z&�av�}�<�!�IgM����ĎC��KVgv�<QuLC<��,p�49�-�r��z�<Q� �"d�B �R`��#*T�<�`�J�rb�D�"�M���j`��_�<y�fQ��DE��F�<$�fLҤ$�^�<)�F�>���1'��Y[xE*��V�<���ڤ����Y�NY�����N�<1��N�m�4A`FO�)3���I'�q�<a�ID35 ��VKJ"����D�b�<�	Ծu<d�b`�K�l-���^�<�C矚]�TQѥMΉpv*��e,�~�<�a��,}�,����̉!��2�)�{�<�cR%/��a�"�ڼQ�0P� .Tx�<�6EU��~<��f���ybH�I�<��D�$H�H�r�®~th�G�]�<qA�Z�&-!헬 �̱� J[�<� x��K1M�!J��9Gnm�"O�Tۤf��!�̸@�<��b��>D����9Mf������x��C�d*D���u�   ��   �    b  |  �)  B3  �9  =@  �F  �L  S  FY  �_  �e  l  jr  �x  -  �  ȋ  �  ]�  ��  �  %�  f�  ��  9�  ��  ��  ��  u�  ��  *�  n�  ��  B�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�VO&}��a4/zY;�#m�����#D�D1���'�01Vo^w:,�U�!D��1G�;(�x���n�$X�6@?D�P�$�Õ�ha�v�C�y �a=D�t�+�p��xj�N9N|�C�<D�:�K�<M�N<ca��*�Ĥ8��9D���������%� .�7Ẕ��<D�L�p-��h�u W$�[Ri<D�������e��E��V).�&9D�T*� -5��dKq�߾{|��聥*D�\�t��J�9��D,~|qR�&D����O�RtN�I0�6S�L�jUC&D���f�a�R 	!�j�T���$D�d8�FD�p��a���t�L�b��&D�|��揺-����e�˳I$Z��A�7D� �Q��,YX\�;5M߾[~X}��5D�p2'����(��R�,�^)#��2D��"�V��V��7-V,�^�QEF#D�(!�c@�x��V#�FP�-&D�\:�英B>��aι�m��#D� ���9SO�ؠE�l��В�'D��x��̎j=*���?�J�A&D��Z%��.}> Jr`�89wQ��N>D��TBԖoƾp�1���HIF	!D��-�$[� ��T���p`��1D�d����S�����K�,t���h%�/D���Cn<5TP��޽2�x����-D��[#.1S���g]�?�d�Q��,D�,��'i�踰�E391`�֢/D�@�OH=�)��ƀ�M��4�,D��8V"J�Rxv&� +�4U��*O6�E��#Y���d�Ѯ8�*�HS"O�H��E�<X�b��hF�U"O�cQ�0��s�;-�q	�"O�P���,�.�8qe��N�% �"O��HE*UR�����]U�T#�"O���HIi:�֧�\���"O��[����d�@��2�"��"O�kҎ��.����o�-|�Q!�'�B��P��B_�TQ j��G�II�'<VEZ&��9/<Փw�׳*`��I�'ސ�������Щ� /���
�')�9�#�W�cp
��
тTx�'.ıRV�A�Ws��id�D�o%8���'�΀UBDE7�³j�����'�@	�W&ŬI���K���-!س
�'qPȻ�+Ӽ	��E��
.�R�
�'(�D飦�"�`5 W:�U�	��� �<(Ĥ�
N��Y��KUR��ۣ"OvtSqJݲ>,8�&��w�2|i�"O��S��^�@�
�5/ɬk���2"O�X	A� ]1앪1���
1�(��"Ỏ�F�>�`y��-��He�'@�'2�'R�'���'��'N�
 �A"t��I��޵R�0�{��'���'B�'���'���'��'��������)�/��{jP{Q�'�'���'�b�'�r�'��'�Qid&Ǹ Ub4�^�l'邑�'y��'�"�'���'Cb�'-2�'w�td(ګ6���I'Kx��G�'�R�'���'���'~��'A��'��%�B/�K�lX�5�!?�.8*��'�R�'�2�'���'�R�'�B�'�V�A���mО);�,ӎz��Ybt�'��'���'�'���'���'��Q��L1�tT�����.̋W�'�"�'��'2�'���'���'�N�Y�D�%�.A9 ��k\T���'���'	��'�B�''B�'ab�'���4��%%%�!	vMIx�J|��'���'�2�'���'3�'�B�'���X5 Y��N�3ӭ�`3x�҆�'<B�'�b�'���'���'9"�'2�p��f�_��Y{��JZ,����'rB�'���'r�'���'P2�'|�Ju�ݤi!����늏"µ ��'x��'�r�'X��'�b�j�����OtUP�GN)J|�!r�Q9���`&$Ey��'��)�3?Y��i`� �*�Ɣ`�@�,kx�С������O��<�'��A��`:�#M�Ι��l,[��'G�����ia�	�|RC�O��'J��}�f�<ܴh��FԤk����<����$,ڧ �ԝ��@^iۺ9�F��!\r����iH@��y�i�O�.�rP(�{fb��Xz�X���O������O�	U}����b��F7O|*ĩ�3"�L��D�Ew
�H�9O"扔�?Yt� ��|:��k)����� t��(c'w٢��p�X�'d�'�v7-ږL?1Oq� cH�GԸ��`�2r�|���0�	wy2�'*b>O��\"&!�2,[p?��S� W)�+ ?a��Q���NY̧Q���N�?A��W}~P�&Lܼ3��Jb#����ĺ<A�S��y��!�9c6O�3qm2��b(�y2!r�Ft�4��h��D��|2�IU80=x�h��\�* �	���<���?��-)ݴ���i>�0��U��u�3��O�E�5������K�=���<�'�?a��?���?Q��ۧJ(<�pwc�"s�h�ivD�;��٦�RM��|�I柈'?u���0Q 4��@A(�)t"�:*~D�'�7��ᦵϓ�H�����eZ�8S��@��jx����6Q�d��X�����ç&���I�Gĉ'.HʓPL�y���Ig>�ˇ��n4�{��?)���?Q��|2-O�mo�0T����ɽr]��6������部��;b��������?�+O��m��M��Ee栙�J� OӠ�Q$��B�n��+�M��'@��km=\b��I%�ӽDfk��-2T�PTm�-h�����l��j��d�O|���O���O��!�S�A��0�Pȏ�w�@��C�*0Τ��I���	��M��F��|Z���?qH>���~�6T{�Hξ'�\l`�R{��'�R������Ni�v��싧�R�(wL\K�E��;�ޑp ���(<���'K$&�0����'���'�	SE�7Z�(Y�F�*l�Ea�'tB_���4h�������?A����]�75\\�bh�n��T�FM��e��	P~��'��f�:�T>U��g 8y`ezB�� 6[�ѣ�]�&5��(��'�P��|���OH�L>!��N4
`���U�@�9�!eL(�?����?����?�|2-O��o��HH4m�qϚ��`�8�^:���PaFyb�'��OZ��?q#��xy�B 0�T�c
"�?���i" �ڀ�i]�	�L�P{q�O��/b@' RnPb���K�ϓ��$�O���O���O����|����5c���V���m�(�����ϛ&*��V���'3�����'��w�l1��g��H��I3I	� ���'���:��)V!ch�6�e�����	�7`޴JeE��N,x��{�M�US��DQ�Iny�Ob��j�� 1իS�Q�����0W��'�B�'���/�MS����?Y���?�폦z䒘���M<:=����mߨ��'A�IݟT�	���L�b`�
)p[�IC
C�]�'�|3��\,���[����ٟ�[��'��y2Ԍ���$��s�T|��'���'��'��>��	3fA$X���B&�ң/��h�ɣ�M� ������O���k�a��Չ;�m��g�s>�	ޟ�ɤ�M�+آ�M��O �i�B�RG(U���jA#	<r�����.2�P�O���|z���?���?I�U�X�a�V�h鶸�Q�Y7D�\�j)O��n/\ɸ-��˟���u�˟�ңˋ1�HP�E��iW�I�"�KyB�v��Do����S�'�^}��c�Pp�3��/� <�靤);��'Z �z�ES��L4�|�U�xc e��Il�9b��M��|��%n�����i�6��O6�4�.�ep�6��/-�BX��2%V� 4�v`O�$f�'��OV�?��47��O�|�̜`gBC��^�y��!�sW�i0�$�OH|��b���������� ���4b�.v>:ak%"ScZd0�$2O4���O`�D�O��D�Oh�?a����P)���%N�1	�����Ɵ�	�hڴ�j��'�?����;&9 â	"���S��3{������x2�'v�O>�I��i+�����w�R/r��C�YQ�z��B�_}�R�K{�IUy�O��'tK?J�镊¥`����u���'��I��M�Q���d�O��'V���ua�`t�:�I�?i��u�'[�ğ��I���S�4I��Ӱ�k�'�%�6HKr�"g�ԩ������O� �?u)1�$ˊ}���3V���;�%�f ���'mB�'y��OH���Móh!tTL�F)�J���#!H�|�NZ/O��%�	fy��p��#pUc�:��U �80�V-iv�����Z۴�ة��4����9����'��S/Ns�PC߉Ch \ �@��6��}yb�'��'�b�' �S>j�C�"�\,��*.���xY,<�nZ�^$��꟤��b�'�?�;PX)�ɏ��5#�
��7�i>67�g��֧�OTlP��i����o
���KKd'�Q#��\���A�����!�B�O���|���yȤ���F�N�⭹��S&4�v�����?y��?�*O�eo�S�Ԍ�	֟��I!#,e���@��
�2p�P�s#��?q�O(��f�J$��1�A�!vÔ=K�T(��08d9?Q�B)=�~��t��E�'0�j�$��?��ٴ�FĈ�=mpR��M��?����?q���?i��i�ONbf�� !���z$P Lp,rR`�O<@m�>[����Ο���F�Ӽ���Q��lU��m@�Mحz���<�r�iҺ7mæ�	s���e�'�`Ye�B�?a*"�ʿ#h*5#��:<vuځ�A�T#�'�i>�	���	۟<�ɷz��A�@�?V�ش�5!|�N��'��7-�'@��$�O���>�i�OX]b� r_���e��B?�9��<A���?YƜx����5w!�͡�nH"%FA+��ۼ"��ɒR+���]�QEջ��9�ԓO˓8�8�@�W rE�RVog,�����?���?���|�)O��nڧE�\���2� �d  �P[#�Ӝ�$��	��8�?�O���d��pl�%I�Р��И|�l4�f�E�Bl$9UJϦi�'
�$R�?Q�}���P�H�s�ҖJRz1q#�_SwP���?����?Y��?����Of�p����YNVHq��J2e)�Zٟ��Iџڴ`��D3+O��� �DѶ�D*W�ߣ:�QQ�HH%he'�8�����!H���mZ[~�h[�����李p�f`�Ug^�>���Z��̟�'�|�X���՟����D�D�G�=,��c"T/4B�43v����l�	by2�r�A���O�$�O��'j�z�xw�]-y���MY)�T��'i��M�g�i��O��H�eꎎO�bAx��!,�}�t�=�ʴ�4�-?ͧt$���P���*xU#�-

�V�H�KR�؍k��?y��?A�S�'��Fަ�p�[�}��Ѣ�7]@�D��9���<��p����O�űG�55�J���D4`�B�ODQoi��m�s~������Sc��H34���ǐ�Y�Tѩf�ȦG��D�<Y��?���?����?�˟�hE�V��.����̫x=���AbӨ��#��<���䧎?1�Ӽ�A�-"���֌I,A�=�tO	��?!�eω����'��$��o�F<O�;� �%+]���3�6X�~��b0O�\2ЅY��?���'��<ͧ�?�`.��Q	�5�� ���(H%��?�?�cυ��?����?a��LZ�.I . ���O��i��|��ޑx��9YW��DY����D8?���Mk`�x��@7����B�R�nX������y��'�*u�V'D�=�8݊�O��I��?�]
��_�M���&gV��)i� �'m��'���ǟ�H��5l�v1蠏J%h]�< u@�̟<[�4n�U�,OH�9�i�Ia���Vq���yZİA冡��lZ%�M��i�@���i��O�s'�+�j�LĒi��E%�	�Ԗ8z�T�2�|�V��S��`��ݟ4�	ϟ(3��K7GIFqA]�Z������}y���*���O��$�O�����dD[��	K�#G �����Y�dp��?y�4cSɧ�'q\}����i*P�0�J��N'0 B���1��'�N�BT�ş�!#�|Y�@3�]�t�Q�D'C.PZd�F��I�� �I��Dybil�:	XVc�O$Ͱqi�
e-T�0ʔw�\�`�O�$4�	f~"�'Ǜ�)f���U��ou@���C�"o�P%Ǝ�H�7-5?Y�`;<Et�i;���iʐ)I�.�j��w)F_�h��z�`��� ��ퟌ�IڟH���b�#�P�#�̅���
�3�?A��?1�i�رi�O)R�'%�'c�A��̆9�PHRX�rU6Oj�2��ֿ�\��\ǖ�n�w~�7KKv���R1U^t(j��I6J�f�C���ꟴS��|�W���$�	ҟ(��WrS���!+D�.�� t����p�I@y��z��z���O���Or�',e�AHЍav�0�!M/H��'X剞�M��iE�D ���_����n�͎I�gA��)��/7������ˁr�i>��՟4�0�|�i�i�,QH݃xK��W"]6w���'�2�'e��tU�Bߴ
>�M0o�I匁3#�J��Dkt���?���?���V�����0#�7x��%�5e`�x�	1�M��ʞ��M;�O����<��J?� �%@Ü�?�|��+	��X��6O���?��?����?�����I�,�$d;��a�F`���NRx�o��)z���ɟ��	I�ɟ��i�����)T��ҁg�V�����(�	��Şk�i��4�yr	]�e�:9q$��C�b	��\%�y⮓GrLD�ɑ��'v�i>-�I�3R 	jgꝧN� 2�S�^�b���p�	�P�'�|7݅/g>�$�O��3O�d<�!E����w�N��?��O���d���&�,2��J�]��`��9j��dj(?�"�S;I��c�i�g�'A´���'�?	�T/,���Ƿa�&]J%V�?����?	��?��I�O����X�h`򂎎��\@�e�Oftm��I\ܕ'�b�4�|%;3�.f��E���2�::"�Oj��x��mZ�'��ul�O~rL�L		���q�ViX�B@���yG�Hnm"D�|W��͟ �	۟��I�l�@�4,U2L�3#O�w��0� �WyҠe�b�����O��$�O4�������>�<�� N&A�ؕ�4��*\�ʓ�?a�h����O1�F^�~�*�84'?%�5�s�N)"��1�OL�� �?IB6�d�<s�PI@�pp�Z�y�������?����?q���?ͧ���ň��؟dZ��qn�Y7.�*�¸s��柌��[����զ�a޴I�����'LN=��h_�
�ҕp�B�=1�y�u�iL��.
-�@S�Oq���N�:�F�sE��t=�V���<m�D�O��D�O��D�O�'���~K
9�(�\��X�%}���I��	 �M�G�|Z��?AL>!)�t���,��X�U 8F��'�z7�����o;�lo~(R�3.v��f�LfO�|rRg��~B�6��)h���`��'t��͟�]NR��?A�Rp��mU������˥,]���%�H���?��B�@z�����ɔ����<]�Z�ZѬ�g�l��O�1�b�	ǟt����d��ğ�Jٴ\1&$	(���$˩d���'M� @�h�&�{u��t�]")��(ԓ�(��EW����B�'zU�gi�e�ێdɎR�#�1�?q��?���?i4GŧDǌ5X��?��2����j�)"����&�@S!R�T���O���3���զ���	^���I�!��[�O=���"���Bk�˟�Jߴ
�� ߴ�y�'��9��Ǡ:M ��O ����ܼ?Θ����i�"O���%!W%=,�A+x���B"O����a�#Czhk�����%xR���l�t!��h�MQw*]�1��q�@c�)W#*�+7��c��Ÿ��� ���d���h03@AT�2l��#�m�x��q�@	4 l���0�N�)����8�s�BS�.T�\�0o�l��Zt�C�2�㕮X�"�p�[�6r�C�-%�5�v��)�2��%-�#lC�T��CK�'B�ҍˢdY�",v�`dB�0��	�4�߽:f�����Q|^d��I�-^�m#g^�6&U �fG�PF�P�0j�qIB��ee����u�%e��N��ץ����ގ�J��	��&P�'�Fn��) l[�Nz�\j�ΉJ��ɀ�}��I2D�8��^�qO\����چ5٦�{5D��B5ʍ�R��[��U�)�S�,-D���p��*�D]S3B.
p��iFA+D��$��\M�9ѐ&Ւz��hQ�*D�DĬ�1IǞp஖�9�yQ�-3D�X�������X�!n�3%�8Z�
-D��Q��D�	w�H�K��� "%?D���V�H+DA�`��M�l��.>D��*� _/i�E��&H�5o�(��<D����k9[�i�c�ӹ55&<���?D�����&d�:�*�HR��-!r�!D����,B�HHY�M?9�έ[BJ:T���D��P��h���^02���PU"O"��@I�|f,���܊330@"O���'!,~�Z�dG�[2$p1"O %c�bY�[��$����/>�:!�b"O�ѱd�0i���uR�c��t`@"O���
S5�2d��m���c�"Of�)�,�/|x��`ކQ���p"O���s���d�xdE^.w����"O~Y�c$C�EPj���@E�>`(pB�"O��#F��>��}�7 ^S^���u"O���ۃ}�	hQ�߉g��I�'���q��EV^,��L
3�
��'YƘ��	�f�J�C���3��99�'���ao�5K��j5��1��};
�'� $��c�m� ʁHȗx��\�	�'bB�8��=�����4:G��	��� ��h��HN.��#�<Zd��5"O�x��%��2�Y���4_WT��w"Oh0�!U�H>��gGD�ei��H`"O|�A�lS1'�"�
�H-ޑ�"O���*�vq��Q���:�x�f"O��(��8J�q�$��@(�x@�"OTԋ��Y$O�\T?~�x4`c"Oȋ���F�a��k߶y��3�"O�٨7As����
�F�*Ò"O�E�¢�:P��;JI+*�n�Ђ"OX\Xo� c*lT	C� v T�X"O��DN�E"RX�@mZ=.���2"Ob<a�υ� z�1Į�8�:�'"O:M�@,�J�ӂ���̠��"O�Xi�F��B�l!6�E�1���e"OZ5�2� v�8�B#2z����"O�[�
�Ky.���C�5*�,R�"O���!a��Z�u��	6B"ObEzClʩf�T8RLJ�$]�5"O8�z�F� j���re-͉4�ƥ0"O���k�M؂x�5�K�Z��!�"O�dA�MEL[�M�"���zz���"O�x7�߭ �ƱY�i��9`��`"ORx*p�BLl��
��k���b4"O�mbw�5�>d[���9�N�Y&"O�$���^�l#K��8�i�Q"O����G�e�Iа���u�Z �"O4x���[��ؠ��L��,a´"OΙ��Id�P���;O)`=�"O�=�f��R����	O�V�
��"O�]j�G֊<�X��-"����"O"����0|(@ F\"䠀%"OI�ѥ�8\p9!vcܦJ6��s�"O�)�K�%J�RL�B�,nX��"O��â����'O�Jx8f"D���`�3��H�G*̫q�(���>D�����G"[S�q�`$ʾ,E@q2B;D��c� n�
�C#��31���P�D8D���#M���܋�B�U����N!D��a�)f�����L5Z�e��!D�|��.B%<��S�ꈬx�0���=D��Se��#"�mCq�2�V�68D��2�(A	O{�|����;c����C)D�1���`X�ܙ�b��Hж�z!�4D�L�LF����3eE<i�ޝ��.D��!�A>F5��I�-W�{��)C+D��97��=	�N�(ᓛQ�D�҈6D��P��M�o�lBfH]�A��
�5D�haT�M�?�6��3`��7p ���3D��X	�"�f̣���:Y�څ;�n3D�h`ۼYqd��2(Ŭv�Z���TJ�<A���.
-��Y�H1$5Vy��l�O�<�'�q�^�AU�ޭDÀ��ML�<�MA�

t��&9�1���H�<��ꇧÈ� �*K%���#�
i�<Q��M3��*v��4{z1�Q�]f�<Q�m�t�� 5�����P� �^Y�<�wJ�2hX�"�Tk�d%�T-^V�<����J4�A�7��3aD�ٺ$�y�<9���`�ly1���� �
��u�<C��qt�SuU> d�X�PLk�<���9M���[�|�P�Q��_q�<��	�rÌ1��6z���Q��EU�<IǦێ^�&�X6!�-���p��O�<� T�JB'X�+^��dQ�,I�@r�"O.MA�L�E�0h�� IH8Ĵi"O> ;�k�<7s �S�E
�C$- �"O�ёG�>{��a�v�Ȋ�*ܛ0"O��ڰ�8w��qa��[6CےA�w"O�]p�"[�_Yl�2�bH
^��"O��1�ϨGR$��@�E�)�����"O���"�txF�Q+ݍx���"O�ԛ��^_�jƇ��J00r@"O` !�:obzyr� е+D)��"O��#�-A+dA���nF
W�-��"O���W���qF����mh| �"O��x%OQ,;��m�AI�P�j�"OLI���}P1B��\�2E��)"O�e#����vp ���� V)�es"O�$��%�%v���Iط}z�X�"O\�i1g��&l�����^�@ȁ"Ox�B���b��Q[�w�b5:�*O��(�@&�j`J�rKx��'z9�G
�*���yg(�;�9��'��mIc˚ |�\�f���5�؊�'���P��L.��G�<����ȓh>��J�фG� ,�7-<�<�ȓC�Z�@���'?� �q־T��ȓ}U8AW�4�J}�2�S7$�2d�ȓx	���_��D�����H��؅ȓ\wvQ���ϰ�6(��'<[�N,�ȓI� S�����9@d���ɇ�^�,�3/�;B�,�Ӥh 
sHR�ȓL�� H���4f`X07ꑃlA^��ȓvn���� �gȄ�f�ת���D$����L�_�`)�B�t��%�ȓ9O�����ߠi�����Z�K�Ĭ��~�nժ�Ő�DY2��ğ1w��ȓv��Ps�!�ɺ�/	!�|��E��j%�΋{�j�``��G@Q�?�@3,O�pr���U(C~�ҽ�On�+�B�'
��'�	�R�%1�d��B�tB��+Ho���h���ܨ�G<3����$�$���<��BOf
ze���q!�X�<i6dW�L�̐�MO,K���i��TL�I)j��?�}����^�<]c���bDnA�҉�F�<AQ��3Q2$aH"��$.��g�[�A�|�q���2W ��v���x�"_7C����Ɠ 2� [��ͬaP���ώ�b�Tma$��e����ܪ-���sA�F�e�4�EN3Ű<��ν�J&�(:��2t+�M@HL:m��-D��{c��5_��pc�v�����7�x,�4A�{����C�z����Ls��Z4)Ö�y"�-��d9�K+f��X"l4��' 	�9OVQ��̘*h<l�x�ҀzBO�0�F䓦/����BC�$~���4G��h��C���0�Aǎs������9h-8U�剾}'
��=�ͪ>F����K�*n� Ӕ�j�<)�'�����&�;p����Q�I� j0�}��D�]����Z�p�2��fdɍ�yR��l亡I�#c���P����'��U03�3O��s�̈́^�5(��H���rO�q�O��`�2�~�����a�2�pu��~��8HFM�`�ej��\�b������>PqO>��qK��А%
��8;%���y��"c����S��Д�й�yү�v&!�s��97IB���C1�y�,Ҡ}�P���ɩ6K���OL��y
� <���V������4��KC"OB�bاjiX�pA��cP�� �"O �2%B�5r��1���AG�g"O�eiv@�6�ptr��ܼ55l%��"O�!��/�$l�� ړ$Zu�"O,�Br��9gL7��-hv[�"O� `͙�I��5gX�nHJ�!�"OZ�i�   �l �eO�%���"O���DGۂn:2���$H�V	��"O���o���D�n�"O�,a�[=p՜�����"H��"OR�� �Ɏ�J�(v��cҤ��u"O��� ���H�i�����"Ot��V�s!�MbvkU��Xб"OV|� ��!O��e��D�/_Ў<y6"O*%���Tff��W$;�J9$"Ol)ҕ@C)WM(1QS"	�+��{""O���T��$$ \��?�<��q"O|�36/�w�T���*s��R4"O�
�DV����1��ܘ!��)�"O* @A��-N�&���@�4AiR�3�"O.�
/����oB�b7�4Ya"OD1� ,�&OXi+�O��d̰و%"O�5���#+�r�;�Q�t�<�3�"O6H�及,Y#Bݲf����+#"O6�[�%�7Z
$#��
=;�i��"O��x�`�8@֐�1�M�/����"O�uj�/�SGl��e��>fp"O�]R��"fCꙑ�dݫz�:��4"OIHB�ޝ7v~���T{211�"OJ�{#��=����Ꮽ/�H��"O��8f��p0ѣOC�*���Y"ObtH�-V��y��ْ>�:��A"O0l�Î
 ǌ�:TÂ\��X�"O�����
��
_)tX�Cϛ��yr�3�%�6㟎W�8TSoV��y��O(c|�[a)S<xk`����6�yb�
-?��!5��s��u*a-G��y2f� bQ��G�L�p?��p��!�yb�	�@��i�P5p.�H��,��y��R<}(����7n�(��+���y�.N�=<e�wC�z�n!��ق�y��5�0i�@�qז4��!�y��V5jf$!5�S�\.�PgW+�y"`\�o@X	!�Y���!���]��yJ�>��MhT�Չ0��u*��<�y��\!����4.��)�� ��ϛ�y"@I�W��q�bַ�^������y��Ж	�f����R ӄ�L��yr�K%���@B�l�T��G<�yr��<< |���b ��.H��O�y����푅K%f8���eլ�yO��n��(b��>uU��c2�M&�ybeD ;h���� 8mJ��$&��y����V;�lC#KZ!d.��3���y������!	�0,-��Ϟ�yBH͌=bT�)�F"���v��(�y�Lنi�uB���/W�m!����y���X���#$G*f��`V�y��3=�}h���(�jZ��4�y$�*�v��B�I5�VL���@��yR��"a�x������)���1-���y2M�
N� `�o�+*r����J��yGQ�G<Z�J��Z8��0���y
� ����O!o��ia*̜0��]�"OJ��A⒞Yx��B	ʿf�<�"OT,�卐.6��=���Qhd�3�"O�J7O� _�\z��ƭSMV-9 "O��b 1 �z��'c�r�J�"O�X�ǫ�|��MRv�],	�\,i0"O�	�׉%�Vx�7���">lġ"O�a�dF1CP<� !��"~���"O"��F�"�.d��۵f���0"OHd�w� |G����Ȝ�^��,*"OB�A�C_��\-١�Fo�^l��"O4���046bU�7�C�%چ��Q"O(Y�q�H �д`#GL�r�F�V"ON ჈H�h�6H]�.�Z��"O�D��d��>ˤ�ё;�&�q�"ON̨3"�5BP�av썥�\��"O
�Ђ��s�i�Z0y��h�4"O�0�ШyQf��#t���"O*}2��K�i��()�
�^Ҕ��"O$�ʄ
h�����ϲ4Il[�"O� �C�>,]bt
�#Z0ٰ"O��k��$5����k��a6���"Oة�����c�Ԕ�𫕺&=ʵ�""OT,�Q��0���n6�щ�"O\��4�ȼHQ~)�@bҜc6()�"O�����D�*�BG>;
�+r"Oj`���v�x1i�ҰB$(�;`"O�1p����j8"5��87�e�"O~���Ži@������:/��a"OV{DO	W�b�F�8or�`�"ON�c˓N��ūs�F�
x��"O�Q3R��3n��č�x���"O��u �&n�����E�و1��"O
�#�L�D�R9�o�3���h�"O��C��I!Yl\���Ң!��\(�"O<w��o+Hy��R�
�^t
b"O8�Q0��+6칀\.�1�*O��*��X|�-�@F�;N�{�'p�eXd�Ҏs�!���1�� J
�'J������|���Ө<�V�	�'r�x�cG�X�� #���0�h���'jtA��P!�"	�Um�"��e��':���ញ$X����lU2���;	�',|��7�M�5b$8���'��-A���V�U�� �6kJ����'�eNN9YV�AEB���,��'�ֹ���|!���b-޲�i�'vص3%�hǤ���6h{�l��'m����숩 p��QŌ�3dF��	�'��� c�J�i����>`�f��
�''�R3AC�� i�@�+� ���'5� h�GHP��E�N�v�l��
�'��A�&eά"4�Q�9�D��
�'�V �$�
�V����/�&aP
�'E���K�t&�X�ҍ�>!v���'f���N�A�B9��'M�2�[�':�u�v��/r~������?HX���'v���		�A��4��[ NeJ1��'���p�܆Հ�)�i�G�0!j�'{\�I�O�<bߪ�ۇf�1G�!��'�8d��J��4>��W�8�R�'��<qG� jˀ�PE�L>Q5j\�
�'@�	�t !g� ���D�#af9�	�'�.e�S�Yhֺ���(��Q��H
��� (܀w���H�ք+8�`U�"O��3H��8HI���g��+r"O��p�SgC�EQ���}~����"Ot9� �݊!9@��ra��\$��a"O"�c�J1���P��3@tlJ�"O�	����0dj����20�Ձ"O��IR�Z<xB��o����c"O4�#D�0V(��㊤M�h���"OҨӂ�U]�F��b��b�~�(�"OdT��!�b�R���[��\@�"O��4Cbp�3'��2?{���ȓ���2�)ȩB�FX93(��-Hz���t����F�0m
��8e�@�n�6���h9����i����u�uS-r��ȓ2�8���Aĉ%r�h��8d��.@�ه��Z�ҁrQES�K�Ḋȓݰ�*�	N�O��0��0_�`��ȓ��u�w��'l9����* ���$�ȓE�=�@��>^��b�ɰ��`��OD}`�I�O��Q��%?�|�ȓj�-Ζ)�vɠ&
34�H��3��Ti���6=��b�`ės}�̅�Nk�����I���		Ɛv���I� 1)���+q��r�A���Ą�L�n��F�!+,��� P�Ȇ�q�Ȉ��CŀXƐ�g6+�̘�ȓDF��:�4g�U�1H�0,6�ɆȓK�4#��:VI��wCҮ7r���f$�]j��-�n�R$�R�d��͇ȓT\m��8~d��BT�H�0�ȓZ-�	�Bj�/C�X'+Ř`���ȓ��}�P�!Nr�J���6�v��ȓUl�����4^Ȣ���K܆�ɇȓ�m�ᮇ�<�6h�%�+Ha�|���6��j��Dٞ��7��d�4$��5:� aPV?@�a�C�
$O:�ȆȓD� %p�&X�6NZ�0C�;Q�Zp��4�fܫoܲd=��l�
m��U#�'�hd�!bN9Q1��<���',lD�p�U9p���qR��zȉ�'t�q���V�����P�{�z�9�'>�#%�R�5�xā��={�����'ي�bTD�c�=���r�\q�'�R�����-)�P�)�唝t,
���'����F�]80�6�s
��e><Q`�'Z�!��_(`i
���eA5]x���'�N���U�(G�P�B��[���

�'n��u�^8&8��eT�h���'� $�q�����o8f�X�'��X��Q8x�~[�.h�PQ��'"`Y�N��v;K��U�غ�B�j�<iq(0x�R��&�z7@���_l�<�g�����tꏀdօ�D�WP�<ipa�?z�z�*�댹�8XB�V�<Y�씘4ĭ"���5a�8
� ZU�<�'�H/Y����ώ.%�b���O�<A�D2�����OձQ��M��B�<�q̄�FMbq�w�\�����FG�<���(\��@�J���9U�ߖ%!�$ūf��@M�%g��B�c݇>�!�$���Uc��M5~6��R�e�3t�!�C�Mz�$���ͽ(�\�+���!�D�m2l�;ԆM;Ant��©�?!�X<<�d����֏kc�8ȕ�^+�!�� ��VFL!�؄i��L�}Yv��"O�\Cr
���ɂ�DYH�����"O�@�$������&C>#�0<��'�x�3t�_�5?�II��T�]Z ���'�A9�^7���Ջ��j`q�'ΘYS� _�(y�#���x�6@�'6�bt��9X�2(�L�i���
�'f�m��h�>��BC_�3j��;�'�l�;p�<Rj�Dx���C<���'g~@�T���s�$�:��<��89	�'������|z��V
a`�%8�'yPh��L,tmNɻB�L1�J���'� �h6�4���2)C�3�8!��'F�a9�ҟE�x�VJG��iI�',J�$傴L+q��J�,D8���'*N�n	��!�\!��C��0��'�i�J�-��}�^�O�0j�'�% W�V0W˦���
ǐM�p��'����%e:��d��Lpr���'����-/�@	���R�KU����'�� ��FS��i�R�D�q��'&c�!�)U&��g�/@̙֔�'�
%kԏ֦/a�Y��6���2�'��Aԧ$g}@�8�ߤ;F���'.X�� ȝKkf�3�C��$��'��(�蔤!���C� �#F@}k	�'�J��+I I��\µJ�7;�����'�Ω�0B-0t�����<�HU)�'���;㋕�¨��M\̩[§���yreߎc�P�k��L�<
�ؼ�ya/x�|9 �nޖ<�D�0��ǯ�yr�4�V͘�)�$?H`��y�]8$`.�8�fΠ_U��[��>�y�%�qh����0FHeivɞ�y2B+���խ�7���� _��y2aL�U"p�c���+Ln�ڣ��y2��D��(�[�*��M����y�k�G; 4�a(��(k<��C
,�y�%��~X��0��j����QJ�yR�@�`���3vc�j�:��I���yB�ؔ>[� �A牝Z>�������y�(P��@��CR�X�D@����y����J���s$� �X�ẻ��y��Vq�$��B�6u����dë�yr]�����OJ�W���/���y�	��r?p<e��%(���M��y��yK�@:g�Y���}�a%�-�yR�-$y �$����q�&
��y"��i�rh��j��A2y+���5�ymF9d��*Dr�vYs�#O�y�h��[��� �V'l�D�ٴ�ӑ�yc�oT�yXE��%j�,��D����y��@�_4Hp�L�c/0K�j�	�y�� �%`�jA[t>T�����y��� �F�bs�P7B����bgʗ�y�*�[)* �Kʆ�3gj�/�!�d݄Rh~��0w$�Y��Z�!�Ă >�cb�W6kl�X�P�Y�!�D�/�\	�R��-`�y:deC�P�!�$�*}�$��%� uu$��I5P�!�$S1jd>� w�Y��P�"�ڧ�!�d�"a� ӣ��7�2B���!��N!�#$ �t}��St���q�!��[?�>}��e��(zD����:cT!�� �c��A�k�dUp�I��A��A"OT�Kҗc+&�Õ�=-լ���"ODLـ`��0܄��g�H%nFlB"O.���ܓGH�0��pZ���"O�� �t�5sS��H����"OL�ٰ*F� ��Es����)�t�"OV��M
�a`6�)¬C�l��I""O0��a�m���J��?ݶ��""O�Z���Ű7����4�NZ{!�D׾#�=)��e>� ӊ�Dg!�ĝ	_f�����D��E��^�J�!�dT1<�-z�.@A'�ȶf�!�D��1�Z��Z� pK���3�!��`,����!,|ZfO?5�!�D�7���.tX���v&�)I�"O�ث��K�.�q!s�H�( �;�"Oū�h	8�5K�!P���q"Op,��̚�{
���Ə&x�Bqy%"O�h2B�5�E`B"���bi�"O¬�s��(�������{�"O*�s�P5D�����:m��4�q"O`!;�ʑ�h{��s�� 9�"O
���H!}I �wc�$F+!��
~��<f:����W�g�!���8D����#REYԂ�8�!�d�*!��|�J�Yg>2�S	dU!�D_�"�@�b�I4Y2Ĕ�"�L0!�D̗ �	���ۃ^�,�ۗ�҇i!�D��IzaF+K�e;��^�N!�d�iR��SdE�lhnqoA�pV!��4A�fH)E�4?^4���9_C!�DQ3x�:`�iE��˒��+a�!�Ā�zz��ü3[.��PV�ԊZn!��خ!���J�<5lD����>h!�$F$�21Q��$G���ڳlÏd!�$ �9K� � P2A���R6
�!�D�,T�T(���í���C�-	�N�!�ݹi.T�W�y�NP��l��.�!��B�x,(�KL)�hE�S�X4Q!��7f1�E����q'<�@�^*6R!�81$Z5�Ṗ0~�b Y#>L!�d<_x�˖,�9m�U��6F�!�$��)g�E�Q��<hj�A�� �!�$F2<���dH,��d��7-!!�D�_�m�P'Ӱp���aa��!�$JW�Q�s'�����%R�!򄉿~��`��F�2"�R ��!�ݒ42�T�@W����c��LM!�V�:$(`*]9&z@����:L!��G
>7(1r0�Ѩ����H7:<!�Ƽ��� 1�H8�bV��""!�䓁b(���'g��G���H��"!�G'
�<h��̇�ް����M�j�!��#j>� �B/ۃ}FYٖ�_�j�!��ɴ;X�G��<Ci��h%�^�6�!�3n(�b��ΨUJp IWG��Py"␽T��t*ŋ�$=*�&ߋ�y��H��L�ڤ�Ϥ^�(��T �yb˓+k�Ւw��'�n��N��y���u:���w��`Hb�R��y� @3�
\�CL�3Yv�〉̦�yRC�'D��A;����ـ`�L��y���#VZQ�is�p��W!�$�T1�T��oT`r���e��!�� Ȉ��㇈Q0Ҽ@�K�*
D�t��"O�X��*�&�d|����8)��kw"OJ��ϑk A�˘�=�9�"O^�u��3�RH��i�(9Mb�r"O|�y"1q����/W�?��"T"O�����}�n���58 61j�"OV5�I��k�*M`���.�kc"O���`��F�b%��.�:hp��
@"O�M�'	-"��+f��7CzF��7"O~�"��96�G�oj�%��"OH%��n�fM���(NP@�S"O�i��֓~�u�U�^�Oh�|� "Oz()da��-��X��Ң5`\��"O
��E �f���ц����"Ov�#��PPd��SJ��zS�"O�����X���1z�ƈ�zIB"O���$Ⱦ{v���v�Z�L�2"O>�Q���5�6�'��e��"O � �һb�t@�1�V\��"O������r�j����HR*��"O��i3HX�_����b��jE�isU"O�<��R�ʚA�`�!)�䙆"O�H������Z�����I�"O4	�P�� qč*#�I��ɢ�y҈��<H���$Tgn�!�M6�yN;DCҠ�R�W�A���)1I4�y�
�e$�	���7��L� Hͤ�y�d˫~2�i6��,)�`� )��y���Y�:%�2��P�`�PG��y��ٜfP3�ܹIp�㖌U>�y�_�*�"���B��"N߰\�`P��Y_�(r��Ƚ^_h�MO�"1�ȓe��[���Q}^D3����Q��ȓs�bܑ#MKed<��V�$`���[��`�v풓S�н"+Êc~@4�ȓ?���w�O>5R b�
.��ȓdf0� ��#���W	+���4�������g��"�"�\ �ȓ]�����!�?V���˃k�.��������k�	;�%Q�AS�Sb܄ȓZ\�ɸ��[�l$�MH�B!:�R��ȓCSإZ�!�~xݳ�B6T���ȓ_�1'��009IR_�2��Ʌȓc�����O����w:-��x��p�H5p���V���`	�Q@��e E�V`#|Qa�K��ȓLIF�#R�[
m�0�@����݇�@�PK�������
uG��q�"��ȓk?�Y��-ź�>)�s�F�[PZ���m��4��
�5k�,�a�L�[���C�"�y�W�R�y��N�d��<��BN�%�'m L�f$*4��%e��ل�k�4\CWa�7�A��%O$.M4y��RW�XxS煵c�I�!gK!H�T�ȓM)�\�CL�N}�4��Xr`��	�"�7.J	.<H�GY�U�8���&�}+����bQ�IC� ہ\�H���jO�seܲ�XE�vi�8�^1�ȓ1j�Z���x7h����1������� �@�H	*#�	�2
D(j����p�� !�*HKn(s�J=W2�<�ȓ=��H���H�dph95��?J+
y��d� 4�S�7߈Aɗ�;�z��ȓ%�T
����lP��V�j�����S�?  :!�E�<x���*�3��Y"�"Ot��"�������c�'
] �2�"O�@�O�8<xUC��;T��F"O�)x�N
`�a���8͑�"O�ѓ3�>I*��[��5��< !"O�ݫ����eބ\kE��/,HA[�"O���OV�s; 5�FI���\�"Od�QA
�e��gF(9r$"O���Jۮ/�(Pr�'_�mB ��"O|MpDE�l��f�!N�#"O�i���W�kr�Y����>��I[%"Or%Z�,2cx��W�Dzeᘍ�y�@�:l3�d�U�F� �"��T�]��y"��"� EHĉ�8v[U��䝳�y�ʈ*��J�I?l�2��bQ����hO���<�ňٯ����I�2W��q
�@�<	"%�:#Z�ԲD�ê,W
`*c�<	!ܦ?�6 ˶�L*PL0LCԈK�<�a�-�6��6��Sþ�`��p�<	nR�<��9�E��v&�P֤_o�<A�� ;�JA:��.-���Gk�<yf�!����-dN֬)��e�<�4�x� �B�U�~��E�Id�<��Ā�g#R	4 ��h��y!lZJ�<ɶR�7{HT1�J�o88���D�<�&E�b�\<y��PH��D���<�䄝�d��=��ɋ�v�� �#O}�<Y�D��d(�YU��1���p�KFA�<�2gΜ(X�@���-)�!r��F�<��R�0��@�#�'W
yX��VB�<!`
;^�x�� V��Ś��e�<���0i��gʃi��Ē�*�l�<�e��WtݑCL�d:Fb�e�<)fj�,A.5��mF�W��t��b�<a�ɥ[811��=�"<+���^�<�5� &�\kQ@H�A(Nqp�D�<q^zH�bv#̵U���ó�F�2B��"K��1�f�9rc�$Tč�VOTC�?����/Z������%���Yh<y�ՐnP�up"�^�gDu����\�<�G%HC�l���N�a�F�@���^�<I� ��1=��q�鏇_'Np����Z�<��Ӊ{�fC���w��y�f�\�<i@�@"b8����ʆP-nU�cE[�<)���w�@a��*�7�N̉�.�T�<�".�9�pU���{��Q�͎U�<qv�^�@�h]As�.�l�h�L�<��"%&C�eL�V��h1�I$D��1w쐏`t�-��A];)�8�Ej%D��"W��Vmr(� D�&*�̑�o#D���`�ϴMF���$U?zθG�?D�4�1�8e(��[@AD{�8���;D�Hz5(H�)=���B��*v(3�,/D������	9Rs��O�{TH�Ņ!D�,�E�BH���/Μ=T�*"D�(`2 ����)Fi�q����M*D��!�m��6�j�G
�
C ]xV(�O.�C��zC"�l���K��	EQ~e�ȓ]���JR��?>R ��Im �ȓ0�)9�jϡ%�2	� ՅFܔ�������ö1��yҔ
X>S�����s��D���ŧV�,�KE��^��}��-��DaōN}*�KЬ�i���ȓrU��3�M�p+��#�I�tm䀆�S�? ��
�!$�n�
���1C`0Qw"O�(����9�>ѫP���[a��(v"Or���.}��tZ!J<ZHr���"O�S�J������$�?#\�H�"O�����p3�4`��v'n��c"O�Up$LF4��<h �_�;3����"On��c���	�`�A���i+�d�'>b��;\� �!��{�a�D�O�h�p��ȓ2�2�����,�n`���=a����{k����!��Dm�%��Y�Av݇ȓ.��Q�v.��Js��Bƒ���ȓfe�,�`ΘB_ XZdd��ˢ���1��m����3 �0r�66�� �ȓ=��!�D�<� ЂAU�T;$���П�'��D��'d����+��q,a+��=�$���'F���n�+�*1qF�e3�I��'�c�Y�$61�D�LX ����']���T�_��*�E���y2�]F��ȓ��A�@AD`���yR��
3�f��1���$�lt��jS��y�CK/_�@�ʃW'0������G)�yB���R�Խ��-P%&��e�2ꈼ�y��)G��|(&៫%=��3�Q��y�!ħ#�BL:G��I�Ԥ�Ƙ7�y�˛�h��C.I<<9��
�
�y"�,m�fYId$�l�X�C�ݓ�y��O�f���)%j��Q��J�y�C&g2�y`��<75� I����y«�D��pS��!L̍��+��yÓ=Ҧ�CB� .� �ή�y��7P����ՆpR t�GG��y"��	�]�������OP2�y�!�h1��ţ��p���ǋ�5�yN��[� CG��sz5	��y���6�V����@('��91�]�y�$$�j�;1+r�ub5��<�y�b
��5z�&Jm99��\��y©æZ�J�[�Z�d�\y1��ُ�y⧓�N��9��e��I���qD()�y�'ҹz�V�z#k�42V��9%Ɛ�yb�7�؍���5\\XQĢL��y�.��/*@hJ�l�9M�
��yR`��5t��I�3=�t���U�y�O�d��z�I�ľ};f�\2�y���7EI�����M�P*�yb`܆]`�BjW�Ύě"�J��y"�� 7���a� �5���9�y2/���q�T��<Y/.-VDɜ�yb�׫�J�̭Se�R婕#�y�E�<y&2	� 'U�L�X����yB���_��Ys�G��Qc���y2b]�g�T�K���9�)顯٥�yr����AQC��CXVa�A���y"a���XܓD�?��2��yb��S�8���ܷ'�rT����y�*ِa���qh��"��4�vk@)�y�LN7����DW�(6�*�y�چzt[7��:9�Y!&`� �y�,_(z���9��
.�p�P����y�M\�u��{Ƣ�)�����y"ņ���Ԓ�iŐkO�=���L��yBi��|�h�%%^�e������]�y2��wH9K�c_ /��1j���y2��|`�pR�71P��� ����y
� ��;���X���&K΋@��p�"O��)QO�t	�yz�iG>|�LqR"Ob���ɞ(o�ұ��(�$�j "OF��f���t$��Ǔ�F�:�I2"O2�K�f�WR����R�&���!�"O��:Aā�!v�3d�	E�.Ԩ#�'I��'��
���7f�B�1�I��`H�'nH��@^�t��5T
�53��a��'�v��5:H���ş(l4�!�'�8Az��Ț)^�5�2m��T-��s�'�ʝ0%*�}�6����/@O0���'\���c�q�S�M��4�L��'�^�Ɖ�-6= T	��1������?Y
�D�|Ys�Z�W@��q�n^�H���A,�pC#�J?*d�hG�O���ȓl��Bv�4�>�����~@����ް�RQ�P6l��'J�??���ȓ|L��x�&��<�9� �ɀv�x��ȓ:�(`2��ʦ	�.a9�e�>��ȓq�p���)��V��h��޾NIH��ȓĒ0 ��T�B� a�5ϲn���!��}iqiŰm�J�KP�E.��Q��,�p��gV�
�D��2O��;�4��-�:���C���������^��ȓad�X���_�v�kP�`x*��ȓJ$6u���\�$�nHo\���L��'H��q�.#A 2���|�N ��'{�<b��8��y�Wg�80�B�	?+�$�h�#�� ��a
±��C�I�}��I�d�R/bW�������DC�I�0:\35�!rx���
ܾ,i@C��.�q�AaH4�,"ai�1�^B�ɯs`�	(�I�s� ���Nػ~.rB�	�j��@���͐��t�󇙵q�|B�I+MX CG���,Hr!�p�U>B�I-��r+��P/�x4	�:��B�	-+8��𢎐D����>)P�B�I��!��%|r�
��B�f�RC�6`��hS`	�$U�� ӪG=�C�Y�h����
�u�bD;p�ۃa�&B�=yf�@rrƞ�gBjLc����JC�0l�a�&9?NdJUI�/) �C�	�A��X��FI�
r��xR��M�C����س�(E_3l���ܱr��C䉂 �X��7/P��� A��C�I4Q���fe�y�&���C�Z�C�	�Y1RA�7c�+pMX�w�ܗA�@C䉰F��EY`@��4Y��nЩ[��C�I�3֧?̶=p�
OxX�C�	�.�h;E�z���H�ΰ��C�	-yj�(GΓa�\s�96ؠC�I0&� X��  ��K���w��B�I�d��BF�ȸV�0�M5(	�B䉵!��i��K؃ ��Ti�h�c֦B��1[��d���&Ln<[t�Z��B���zi����p��e�'%�d3VB�I��NQ�cW�-g�-q%ġ+��B�I9kŒe!
1*¥YQ��N]�C�	�0�Vq�"�Z���\ ��3=v�C�I�B�,�*!��$��K�W�B�I�&(�4[��G"��଀8n�ȒO��=�}���2��ǌH�f��0��HV�<!��M�O5�<P��)�4�ub�O�<���1;x^P��f$�<�!`��K�<� X���a�4e���vG�,gČ�"OJ9����w��<��GM�\6V�i�"O>����R���i��ۮ|I1�g"O�%���$�:��6�̋;4���_��G{����Z����iF �����f�!�$ܦ@�v=Bum1>ɮ4hݽ<!��� Hz= ��V�TP�!��*�!�N6z�}�iG�^���u�O/)!�d]"O�I�Ѩ�s� ��/ԋ!���SX� �F/
���U�!��Y� hip'�����H ��'�ў�>�3�E�"$
���-Xd���5�?D�\'MS� ��'K�G���G�2D��S!/t�1" �n���E�;D�TR��?U"�y��^�#M$�I�N4D�����P�V�X�o�I��kq�$D� ����4G<i��J�
XSZ����,D�l8�AY�d=pay���5i������*D�H���ܒP倩�"i	��P��N=D� a!�/2d<�Y�ܼl���J�6D�D����%@���+�hL���(D�t"� H�L��&ưW�Z��w%D�(ð�:w��y��O}>!�#"D�X�H,v�"�2o��5e��6�-D���ħD./߮�B6�Q�&�ٷH,D���1"ޑn|�+ Đk��[�+-|O$�D2?�b�"8�|7$�Kεч
O�<a��=h��*�MռZ&^�!�$�M�<a�F��x{�h"c�:E!�g�D�<�E(?��i��H m���a4bY�<)��,Ly���
}
�d��T�<٣'�b�P�r�BYKF�"��_Q�<q��I��J�jZ�7Ϣ�"�I�O�')�Od�)��\�\�@|S��E�0����ȓr�j��/��G���jU�&x� �ȓb
�����[i���Bv'N�Q5,��<?>� �4p	�Թ�'�t�5��u��=@��ڦk2x% R�V�8)����`2�A���EvX�cU���\��v\t���HfN���M"AZ�'���Id��DUg����]�w�U=��a�5D���E��cYB�Q�+�M]�Iq+2D����)y85b��ԔW�֤��5D�H��EB�W78URD�l�b����4D�@;�,ԝfblQ˱� c,@�rA8D��*��V<��K#�ޘO�n�0 �<����
fT���ա�R�ҙ�Cغ[�<�=)Óa!8E�i�/� {�#��D��w��A`)b�"c��R����ȓ2�Xly��#�r��������y�BT�1I^�G�,��1�ֽː��ȓ{U@�W�EZ$u��F�h��!A�����R�;��4M.�F{���<��3XG�tq`��0{���3�^�<كG�i	Tݒ��U�:@m(�CW�<�G/����a��,ew�H&l�O�<A��įo��Z�����ț�A�<A�xK�@��C:�P�3��r�<q#BY�1�C7�ۄl3��"Gl�<������t<��O�>\�q�l쟠G{��ɞ	~�h����B\���E�F���C䉟I{^%���T�*����oD�k����0?�p`��itT��m
.fQ��h�<`"\+~�p�) o§LYJ�g�<� PM#��5�؀!�O���8G"O|��*	i����%%B��Xg"O�9�ת�C�pը�*�+><br"O�˓�ǅ4�F 3��yq��{'"O�|(��
0z�<D���Ӕ']l���"Or
�+���z��ǋ��W�<�""O����	�\jD%_�@D�p"OHrt.\2_J|�ˑ�py��4"O�Hyq�Z�*<���#��L~�#g"O& ���	Z� Ѩ$h -�R"O�<[���P�FP����H��1��"O�yQtbA�C��`���=[�Z2"Oe!îӊy20����̱<PBRS"O��+�ur\�ZCMK�a�U[�"O2���Ef�٢�J�`qQt"O�X��
-=d�%zw*�)&�xQ1�"O<ا&B�VP�Ǣޕ#�:�{p"O� �b-�<�$�r����:%"OdE��BV3Kh�h��a	������"OĀK4(U��@��&E�W��x��"O�y�Q��/kUD�	��G�#�4��"Ov�eFj�<���ގK�$| b"O�E�b�X�i�:r�i�{P��"O�9���R,WVl b�B]4^a��Ie"O\,rGQ�(�f�xᄖ8]�a"O�f�1J� ���Bi�F铷#�<��nnD0&NО,�DЧJ���|Ş<ó������a�-��ԅ�'}t!@�)�����gP){H}��V)��S��5P�+u�6 �`�ȓ�؉�g��zT`S""T)F�(��p�B���H�6
��*�bG)M]ƹ�ȓPSd
e�1^|��NĥVN �����!g��.�D�9D����8p�ȓw����M�"z�h`�P�]�!���NI�lSqA�8��If�в4!�D�����[�I6AVV��E�ӳ�!��1Z�*e��g���1�9�!��qÜ�ۢ!/�\����Y!�d�A�L�R@/Q�.%��	�m�!��V��:�"��w�lв��;�!���r�����ϴ�,�c��Z,�!�d!⺰;�L ���T	�M�!�DN*؜H�e�6>�@ȚVl��]I!�$G.$(@)v��79�Jy�#�BPQ�2�)�dk�B���#��W9O���C"B]!�y2����ɐ�Ј���Xt��{Ј��SH�UT��cf�愇ȓN�������M�X�d��0��D��P�H�Q2�	�u)���g�����8h>�aCM �p��ӡ[�$4��u.A����tw��(���7��?ɉ��~�ч�Kq,��$��4Ct�jՁ�D�< ��=:@i��+�0b���g�<� �]��2l"��_��P��u�g�<y�b܄K �P'�?O�1���b�<��"G�7]:i��:r|��J��QT�<	ã�9��T§B��Rx�����V�<I$/� v5�X�^�1��y��NQV�����n~�  Ӝ!V��'`��,�q͛��y����Tb@$���Đh��� ����y�bŨN���LȨ[�n0I��M�yb��VN ����҈E:�y�m���������"m�t�٥�y
� bȻ5!O��hԋ�g��E��|�F"ON�K��K�2�yr�Ha=08�e�F�����J~"��FҢp@�M�>�L� 
���yʛ ��1�°I��b��y��m�@-��.M6Hlԡ7Ő�y���t�ƀR�%�%=\�ؑ�W��yb�%�-R��Ҕ4Ѿ!�ai�=�y�AY;vI��S�cW���1���y¦�7	���#c�(<@`�/�y�͇^���
"���_��p�gL��yr(y�F��0h(�� @�б�y�����0�+Q����n��yRJ��yf�`�����H�� )6"ƺ�y��kۆ�Rq�į>(�pJE"��y�!�*K�l��./��tp�ŧ�y2DL s���Q(�<��݃����y��D�Wm�QI��`��M0@�N��yRM��;�(�3%_�S<�����I?�y©�.$��B��M>�:A�1�y"m@�n^D��K?3����k��yr�R M���Af@	�U��X�Cͅ��y2.ӊuΈ0D�I�EF&	肤α�y"��/I�t���U�1��ZK�+�yr��$�Dm�)"�� Ӧ�؊?!�D%�e�� ��5z�P$ 
w�!��:WC��95a����b����!���EPh��Ӫ?�l �BH_+b�!�$_��4�Ⲋ�1��|�'ȣ)v!�d�)%��ջ�(�z��"��#Ov!���
��R�Ԇv� ��C�X�^S!�$C"h�x��ԦD�2�(�2��� !��J�q�th�F$�c�<�4
M�L!�Dҟ~AZm�L��
"V0��ȟ5b !�d��h�e����)Q�hH�ö7�!�ĕU˄䒤�ΦJ'|����In!��]�Io�X J�V�j�F1g!��U-D���
�9A&�+EPȹ�"O���C�Z a0��A��#|;�.���"�O�5���Шj�z���DW�Z�J�s"OL�r�Ӌ5�Ή�2Õ#}���@a"O蹲兙�ok:�R%dH,IX՛�"OV\�i��8[x���m˫26��J�"O|r�h^.PM���K��e��E1�"O�T���!�|����͢#ll �`"O�X�!�� ���K'�@�4�X�i�"OJ��L� _�6�����3j9��)""O6��Ũ�.m�R\x�kG�*�0"O�d�G�����C"%N�cr"O´*2j��IQ��Ӗ*g*�J�"O�S뛈.% *Sp`s�"O�)궉�m�l�T��+YN��{�"O�#��P�H�H%
7H^5��Y0"O>i�F@�b�����@�*r=`p"O���q�X�Ty��R̶6�8���"OZ�hƤ����Ƀ+��yZy�w"O
����["�C�ަ.u"��"O���e%`�I#�F�q�#d"O������v��QVF! Y��[W"O<D��R���B%��<Gj4��"O�
g�v���qoG�4aH���"O�M�u�G_W�\��+I�Z�d\��"O��4o�;R�e�jJ��(�"OB43�b^&�X�
�fF�j�±b�"O�Y(ՊW�j�Hb���R�~�2a"O� ��c�ď�(��W�LĀ�"O�lk$�^T4`B]���l`�"O0��ހL:B �V�e~�k�"O�x
���^F���5�ާ>� 9Ar"OX���R�B��"U�@�X#hiH "O���q�_�5u���gcWs� x�"O��x"��X�9p�":R���""OF�9g�'�@kUŢE�\rgO�m
�U�q����N[�� �	9�!�$8��(c%1x!���i��u�!�D�c�L9C�Lb~�XXqIA)2!�D�U���gE�.Ey�,`r��-C!�Ę�v沘�l��?b��i6j�$.�!�$�$�fxR$�V+-�<��0��/U�!�D�5T���*���	���L����
=,�^����.Z�H�9��E�lE~C��2 	(����7�PP�PJ�7�hC�I��R�Y&-TWhѱ�O �O8C�IN��93�ߎe�6db]g'"C�IΠ|����a&,��Hk�B��81��}"`�K�b��l�g
"
A C�I�sIPhʠl����v�4B�Ƀ\��DБ�F*�Rl�'(D	Q�B�9g��=��T#VU:��%�C䉟s����� 6+P��^Q���	�'�Da�t
Ÿ8~�t�%M��Gv�`
�'&0����+(P4��Q&T�P�'��Q�Dj�-%���J��ũ#f�T��'���@�bQ*l��-֓RA
���'��A�TNJ14 ����@V��-
�'ӆ�餦L�wL��Q��*Lk�U�	�'��u�W�S�:�Kq���IuT �'��(��tf�BKΞ<5f�(�'LȅHDE�.L������7]��B�'�����E�h�p2�1$"�	�'È塑���� �v�$\+�'3�C&(ď ͠�8��B�!$X��'a^43����u�����W ���p�'n���!���M��oT?��'k8�2�� ���X�+� �ɩ�'��|�ѫ�%�dH���	<aJ�y�'3��p������!v�@�D"���'���u��>A�}R�#�%�h�<i�_8���Aƌ�1nҒX�FLN^�<�b�JJpz��TI�91�)�X�<�%*�mR~�XW�B�x3r�(��NT�<1&���
<�v"$eĚ���n\M�<Y �T�<1��ag�["9�8b���E�<���� ���:jX���JI�<)ABnt&zp�� �%�o�<!�G��1"�L{��LS�N�tʐj�<a��5\�$h'D���Л�%c�<�u9�z��R��= ���y���[�<A���$'b����P�x>B`9�Yl�<����<c R@S��-B���@��I]�<����n��<���Z�=!����S@�<�p�σ ���1��+����\{�<�$f[�b��,A�#λ;�*��v$Ax~re���0>Y�K��`�����4�^,�P�Z�<�S���.x���ڂ�h� K
V�<a^ɠ� �-*�p`8�gUR�&=�ȓb0��ReKߊ5H��A �$��ȓX�d&b�%n���1��A��$��Vs��;CJ�}���e!6r��S�? DT����D�v�� Qv	($�|�'�֥Ǎ[<��;hR.���9�'��0dg��r�
�Bч�9d�x��'�r�&�ݒNr��b�L5E�q�'��ۡ �8x�F=!0�n�j	�'�v�C�\GW�H�ܳ��
�'�$�;����%�J�+��,��E�	�'�l�W ��	�ō
՘}�	�'�>A�ɏ$8��m�  )�|��'4 -���^�?�V9[�G�3��<��'��h��X'�`[1�_�G�N ��'��ih �Ą-����@ �@�����'�^m@Xh	G��)Sd1Ӄ��y��&>n��SgDF���eFP��y2�*e��&O��Be�X�����y�C�$2xa�"P(;���w"0�y��i�<e��<7�9��+��y¤O<b��$�3�؎?hcg�֦�yr�� �.1��Gl��h)��y YH{�D �-�J�t��yR��o�,=3Qj��4EV�j ��yrb��
�($(��Y�&���y� ���yb���xID3��E	Rm��y� 8] �Y����2�4���́!�y�i��X����)���
��yBA�z�T�*(8����F�Z:�y�Î�,�h��߭-n~�`�*	��y��>gv�2�������6�y�,jA����!H�hѭ�y2`A:!�jꆦJ9r pS�J�yb"�s�8�E�U9����RLH��yg�	�	KW	J88r���y�E�Dv�P#�}�.�x�bK��y�j�&4�fi�U��3y��r�m���y�Y��QRĎth<q
s���y"�؊ -�pk�,C�oe��QŮ+�y҇C8_|,paǭ�np�����y�M&D�0��DkB���R"�ybG�x�X���^�e�D(���y�*Y7*
���� {��B!���y2&חK�HL�֯h-l|�kQ��yB�04�Uɋ�c�@h�'ſ�y�g�7r���E+?Y����邬�y2��%]�-�Ɖ��x�D�S��y�	�=	�v�^�jp�
�S��yH���U�	&�<L�f���yB&�d���c�gB%y���y�̎O�b�����mJM�V+[��yr���M�*(h��H�8{ ����K4�y�L	#�����>-4�r���yrn��o~���N��y����f��yBȃ�H5 � �PrԨź���yr�ٹ!2Ȱ��_�e�B�v���y2�	<�6�C�@
�
��)+V�ė�y��(_�r��6d�����s`�N8�y��]A)x�*2ɐ��ǅ�y� ��+Ȃ���΂vl�d��'�y��G�3�uB��2_�����(�y#���aң��-;�t1��+�yr$�Z^}�G��P��\)P��y�mB�4���ؑ{N�P�C��y"GզW�X5�3�ìb�dLpN���y�H��@>��v��]d6�7�W�yB!��|V�u0%�\�9����y
� 6urH�p��8cg*ߘ�H�A"O����LѓM��a��3O��I�"Oh�kQNص/؈p4%�]>F�A@"O<qS'�ԭ%���:U�͂!=l� "O��)"��N�	��u�H�""Ox�YM�2U����W��2�a`"O��ȟtt (
S� ;�:yZ�"O���v��Y��1����u�L��7"O��Z�$|ԙ�o��~#�]+w"Oy*�(�2�L���c��~,��"O6�����.�ؑ���	���1�"Od�ِ�/w��)cb�J77�~��"O��(�A�(+�� BŮ��6tr�"O\u�u�Y)^�R� 3.ɮ~ָ
"ON���!B�b����wLX�=�M2D��� �A���B�V 4Z He##D�Pi��t2����g 6�R�/#D�l�5��8zR���AI-D^��"#D���5�3D���YwaF�`�B|`�&D�h�Dֽd�"	S���rB�� E�'D������&T�8�#��7p֬�6�!D�|Y�%�8��X�c�vqtY�1�$D��+�$�H�^`GX!L������?D�@R�gO�Ͱ�BJ6?��eQ��>D���ckk�Fׇ�pn�@CO��yR��v%�e�R��@��4J�o�yrIQ�j5��(�ȋ��8������y򅛨c$M�u��z�x� ���y��<y��F�V���f&%�y�Ϥ�I�(���!�!��y"����`ǧ �"��߀-?!�DV�MX|H�%A�9Ft��d,�=:/!�DO,
1�Y!�F�OG��23��"!�ǁ"��ኴP��KBbA!�D�'b{L}��X#`��ݢ�˙�Xa����b���J������Blߵ�y�������̴X��U�Ⱦ�y��L���,��%@37�3�I��y�%K8.ɑ��&-�P��埞�y2�(}q�C)�Q��X��y��T�6�D���eܙ"�(��FN��y�m�F �m��a^���%�Љ�y���Lڑ9�
��4.N$1����y��P? ������\�E�wN�y��.���[��ǲ���q��3�y�c�[P�E�Q��y���4���y�Xo.p��%F?�ࡹ�E 
�yҏW�}���Pd��l��%*�M@�y��D�=8�� �ߐ_?�PC�٣�y��ѐ}@���o�7n�"]3����y¨]�uj��Ύ�=mnihݵ�y��E�J���I��Y�:آ(��A��yRL�Q�Ӎ��>a� ����y2EԺ�,T�V�� {D #�_5�y�MI�A��R�kWL鱣���yB� (�Ĉ�닂3��}h�&�yoD	8$qB� L,��aa�� �y�bʂ:H$�+�c����ph��y"�>;����Pꅦb.�	G,�5�y"�Ix����6�M�q�F�N��yR$Y*����1�S�F
y:��/�y��9���qō&l�(=�%���y�aTt�+R��f�JXFcQ>�y�n\:_���2/�\wH-9tNÀ�y
� B�A����,��A���L�v4@pv"O0�8%4-$~̂��<<���"O����M�-߰�Y�7S:��"O���V�6CF��i�m�4�I�"O�����[5LƐ�Wcʔ@)I��"O��� �H!|��Tb���a��"Opq[5H�2c_��q����SΙQ"O�哧(��Q�|���@\�=PF\0v"Oj}I�
T�v��٣!fJ2-�AB"O��A�ה�n�C��U��`�"OPq�ʙ�L�)sd�(&{ U��"Od��0�,mJ��[�b�:���#�"O�uh��7F��S�/W<�r�X�"O �)����;���w�>�Tyic"O���E^? ��Y�.�g|z3�"OV%@A�T.!�����1~cN8��"O�)P����<�WO/V&��E"O`! �bP�2�iFC4ZC�{�"Ob�ÖfY�/�$p�@���>�`��"Or5x�K��t�=��K�BU��sT"O>���iK9�.yYa�������"O5�fK�\���T�T?>�V��%"O <��,Z!@�Dx���V=4��}��"O"A�Q�AzJE�� N�R�Ę��"Ox1��]�;�|�������4�� "O��I��g��x��ݰ_��=�"O����;]�AH�#ތ|5�"O�i����%\�̩C c� �
"O�H5I��
d$Ԉ�h�E�"O*�aa�^�����ao�?�l�"O��* S�X�p$��x�"O���a�J�$�.%�jL0�`)�0"O�!؂@1Z�`(�D��r���� "O�q����!��)�'�^���"O��3�P�H�r���HK����"O��
tʀ)Hh�b����4�d�z#"O���`?,�A�"��n;�9q�"O��Kf�9��Y�&�Hd��"O4@*3��@f�(8rf�9$<1�"Oʨ��"�A�fhɖO-:&(��"O�����/K]�qc���6�1��"O-2dܵd|�5�îF���A"O�Y�"����qbb�H��- #"O 4؂hL�s�µ{$���qt|�"O<���cOa'4��10T�ia�"O��у��|���g��t;9�"O�H��_ %�ph(�eL�&/����"O`PQ�]�+t,�H@�L11ɼ$C�"O�@��30��*a�EL��z0"O���e����hȉ�d�-����"O�`�K+ H ǄR+08����"O�u"���W��p���?5�MBb"O��z��8Id@��p�_�h����"O�dC�N�%k܎p�S&͡*d<���"On�˞�a2���o߬((�)�"Ox#s% }�� 	��N+e4�hr�"O(;��
#.R�Q
<N�`��"O*�"`��G~l�!�����P�"O��b��+�𸻴j_4�ؼ�"O@@�����L�+���84M��v"O�m�#ц[ʑ����&����T"O���Pa��`{�M�����('"O<<CR�Oto���bB�'����"O���I�F~�A�&� :'[����"O� >�C®w��h ��/,Cƌ# "O�k�f@�k9����F c$4!��"O(�I�C�I-b,S�O=$�H�"O�rD�a��U��q��i2"O^������L�9��'��� @"OZ�����mr���T�x��I�"O!�eL++��<���f�abr"O@!A��I�+���"^,�:QR"Ol�sEN8z(�ș�.��C"O��@�Z  ���z��8J�R�"O:}�5��59�`�ő�P5Q�"Oԉ9����Y,��D�*jp�	"O��X���=�(Myu�R�Z�6�yB"O`: �@���\D-�Q�*<�"O�T,�,Rp��߈K�v,h�"O��ӭ�0L��jʨF���V"O\A�RZ����,�&��lҔ"O��*H�:`��!G�~�J�bu"O�E�W�F�W���7�y�"O8=�"lݨ` ǭZ�^��8��"O�}�bfJ�y׺�HmG�h�t�؆"O�$Ja\�P̜�)qO�>����"O��[b��t~�Q�ɓ3k�����"Oȡ�nӃt��YU	ƪA}��*�"O��ǒ4�u�P�Ґ5�b�""O t�Vŀ4J������U} �Ҁ"O�a;�`U1T��q�BT(|��4"OnQ��N��Z��'�D�E]()�g"O��AW?!��/����	�'JZA��D��U�g�X�kL����'0� ��AIf���Jg�]��'��$���_6^t"0�b�O1gt��'���2AǕT�a�g̯2����'�>XZcZ�Z �J�	��i��'�ڑZ0֝q��4���F 00�D��'��x:U�~ՠ`G�QE�Y	�' ���cǾt}Ҡ�W�8����'x���_�A���r�H�d�j
�'��; `�?>����a�HWvL 
�'/�h�F�Y�5!n$kae�Dx�)�'jt���$�%e��Aa�Z98K2 z�'����+�DٷK�1m�1@�'"Z�ږ��$r���G��=,҄b�'���)�dtÃ�b�ذ���:D���C��5�U D�هM�h�7D���F�2Ű�� 7���H �3D��q&d�3m���b���IȐ��0D����d�$�@�#7e��(c\9٦�-D�L3�җ;�#�ɋ�>%�*D��b,>��I[g.�{d�`rpc5D�Py�˙s�fU��哢)k����@7D���2J��J���MB��i�m4D��C4��J �]ذ�(O�ܐ34�4D� �"�!T^��� ܠe%0D���pcH	2��m�$+�5׋.D�D�FK�2H�P����$]��F*D��ڦa�����׏3�xu��%D���p!N�^�L�A2-�p�d'(D��80�ܐs�tP3�@S�S`�4�%D������
��Qz aV�roj,�FD.D�P�sʈ,[ru#�/U�w�x�Q!,D�j��
�I�8ȩ��:d�/D�;�-P��p�ʄO![�1:�l1D��f�O
>��ICѦҨZ^t�9 i0D�� T��gOI5��
���J���"O68@WY�;G�-���I9�va�"O2��$(�x�V�ҦhD�JP�=0C"O�<`�ټE�Z�*���O��`yU"O�j-Yrx$��dL�E��ݻ1"O��!��y-3U%KA�N���"OLM�fɏ �x5���e. �r"O���:!�Y�F w&P8#"OP�Y��X�S�]�O�!c�P�"OV�k�b�x8ғ�ٙM�es�"O�\ӑ�\f��9��L�'I���u"O�qp�0@� ��%M�V	H�	e"Ox���u�\���Ƒ#��"O��3���'��IVňM&:#�"O�\���A�{� ��B�"i �"O��	��B#?*n��P
X7 R�c"O�t3!M�.�����e^���"O
՚w�� FD�e�ܖ�:5ҧ"O�@ӑN��4b
XBRKC'��(�R"OB��a��lhD4bᚄN�v���"Olz�`˷s�z�[E�]|��2�"O<5���?���	�9]�ӥ"O"|�dl�!+}��za�C�!�����"O��K�eҥ)d���Lc�"Y�u"O m���ޑ �6�{ׅZ+r�0��"O�`8#�  ��9��L�&Ҷ�"O~��J�6�"T�#�P���Y�"O�YG��
^�����E�lU "OT���gղ6{r0��b���¸��"O�]�S�+
Xd��KC$x����"Of�HU��:^����G�M[rq�"O� ��u��@��L�	���D"Oxe�#k�2},4@Ѝ��f+��J@"OP���jН2�����B+
�`"O�0b��Iz�؊�;�e��"O^(��$æ!�g�Q/]���g"O�<XUf�0Y`D�p� R�4)�r"O��qE�#��Lٲ����R"O�9y��N6>E����(@+u���
�"O�]�Ԃ�TU�$:�}��(�t�3D�����M���Y'i8�xY�`2D�8Xd�2��]��Y)?�~�3�4D���'n��i:pI�K="�b��$D���jA�!L�	%�R.O"��2i$D�tˀ�Q�*-�R������ D��HA���%ې��%U('!v�{4�>D�`��hM�lS���z'dmr'H"D�X����~5t�q'�
�*a{�'6D���0͔h�T(@f��n���'D�|�qf�13�\�#��'� i��9D�4�Boӥ,<�t�O<�P���7D����7WVvmQ���,S�X!Qp 5D���-K@`�&�'LZ0���g2D��rl��-o\���@J�3-���.D�L��ٽM~`PÆMI?��H�
-D��y��AP�B�Ѵ��x��(�3� D�$V�* �L˷�E�W���d+D�,�q�@��5��,z���*OZٚ�ꗬI�$i�F��=���Y�"O��A�i	��2�*Ҥb@���"Oj��Pd΋c���,&���'f�\��oY�p�♑��G�*`)c	�'���h�2ZV�h����6lh�j	�'�bUb�ֺ�2���LJ�|ʬd���� @(*A��
���I��ބ[ٖmC"O��)��ʥ}�0����C�Ԉ��"O�)�VG�4IJy���vҾ<�S"O� @�)e�J���#[�E`��K!"O�XʧBP�.y����I^�rs|!!�"O��( �p��5�4OS'©�"O������*~H��'X�쀀�S"O�������S�F	����(}f%��"OZ8��ª���jg�G5=�|���"O1"TG�n���yF+��^�PA��"Ov�1����
Ba� 7\�Z�"O�\��Wn�<��E
�z<��E"O����H�Vs���Y�1�hf"O~p�e�]+_w�h��唟|)�E��"O�dBU;�-;'��>?ò���"O~�W���6��L�@�R�5"O$x;�m�;}N��kX�pR���"O�i��ۥm%�؃���-GKJU�q"O�i�r�ߒ1V$\ g�{,�Q�	�'��')Ԣh� ���X��ح�	�'�8��Ꟊg�dс2�V�_
F)q	�'3.5�H�7[�������U�<��'�ƹSpR�M�n����2S1`!��'$U"w��?@��A޼M3Ե��'��i�#&_-Z@��Ȑ,E��0	�'}�D�AD���d�P�X�tez��'
t�*��57`��`�]�e8�')�L
Ѩ�*_�`�7)��
����'~�Ac��*B������7�����'��l*�g�7E� `�7@ /:D��'�@̉�Ǎ�Q.�Ap-��v����'w���FD��\r�`10�ۄi��I�'�^`3��Vצh��/Z{B�2�'F���O`R��g�U�����'*�sa ���lX*��"dx��'0���F	�s���	�_� R�B�'ɖip���b���@�B�
���'���A�ԱMpbmJ�&�	@"5��' �Aq& D=�F��ѳ7�J5�	�'�� 閏]�]Y��"�Q.�&�{�'�0�/���2�@=R���A�'-*���X��L�y¢��
�'�Fmi�X.q }3v�U�j�dP�
�'ξ r J�<�ځY�7t��*
�'�X(A1 ш)&�C��:��4�'��l9�m �"%>-)�mЏe2��'\8�Xq�#%9�Bc�<s�'ꎘ�'݄/D�9!��X�P�0�'�B�c2 ��W��@�N�B��h�',�A���2 ����#PKX�x�'o��J� {:I
"mV"E�B�	�'�d�c� Ea�(����5���1
�'�
�O�ii ��b葤,"�x�
�'���%�Z�L��c�!��	�'����;lnyHb��(yL}��'`rX����ʸ����.�Ԛ�'Y�8j�0A����']޲�j�'����Ǽ0���'O�d�
�'ټU[��\�G�$E�?���3
�'�N�x�MO	A
�`r���IRZ�Q
�'��lX�I?T�n���1����'��鋴���Fl�\)�c��n� �'xFm*�b֨^���C�H�4Td��'^x��@�+
!�DR�h�x�
��� (�6�C7~�4j��N�`�q4"Opd���h�|(*bcZ�t��#6"Of����c�|! "̑�.���"OU�6���8f��@�\=�\��"O���RGISn2|{嫋�&��T9�"OhL[�*��%��A��i�7k|��Q"O�UJ��o��鑪��7�V�C"O�M�VFF?g���3H��%+V��F"O�9֥�8(�����	�%��Q"ORT���<k<"PAa0��h�C"O>`q�g�K�����@��G�<e"O�iDf�&+���1�NȶL���X�"O6m��c�����d�:
�� #g"O�9�`kD	,ۂ�(����QUt��"O�b�P)(��a�1-F�VD(9I�"O&|qpd�6*r�(��757�!��"O,;6$�5_��6��"&긛G"O�UѴDΘ,�"�9g,��5
�Xч"O�<�4��>/���&����L0�"O��a�ꕷХK�@�<-�����"OT �e�.޼�#���'p�}�"Oα!�j��/�a��EI4V^���"Oi9�Iڞ� EQC�S)&}D�'���I�H�嘧��>�0G��G�bP��y`�|��h*D��`Z-�P�z��[:$̲��5ˤ>���
��-y��'A��,�!<�6��%k�,�F5"� �<�*�HܑD*��H7J��b��dPP#Ҡ5M"���"�Oh<�U�*N�:��(�"8=bt����]�'���#KȲW�m*5�1��F�T-A孂�q���ҧ`��bu�B�I%:b�X@#�!�5���P�:�X�C���P8��Z�mQY��,�g?��̤z)JH:ǁ�Hb��u� \�<��BQ9FWl��
���\�7��ݟ�{$%ւ/����} h��D�1�4k�fL=_����t�N�y�F�=^������
�H\5� �[�H"�| �C��$r΅��D

�Ś�'�v���S�N?xE�C#Mܲt�L<���F�,�}і)�\�BL��)���O�ơ�uK�x�V!��A�?�U��' :`�e�(�H�Pǭ��"�l�j``�'[-"��A�Ռv�v}�����O���'����&T�{���"f �@jԌS�'��Ď۝qu I����V�6IgΪw��!'�R�mq�M�
�wp褆��2id�Z� ���!��a[Xz�?�s�]��HX� �mov]�a,[�;�c��w�
U�%�<iSl5J��x(<Q��^}J\;��-.�՘ �yb�Џg��l��C�w�B��#���P���P5�q3�� U���pc���y"���.1 �8��НqL��i7nՑf��<�£tb�1�d	r�N)N~
��[�$0z�Ĭ���ZL�^��c�54Qa�FJ!c��y2�.��E��i@�AZ5x8�
�mK�%�"DoX��q	g��r��x�j��9i"\����
I�}��A���O���|w$��g�{.�r
�"::�m9��N@.��b�&�t��c\V(<���@��[�h�;_n����{?�%�By����7a��ɫb�\��K�韓^n��;�E��F~�P����!�Np&H��s&�U��#l�G��y�b�:h��#@Ś	5��h	��~��`
4h�e��18��d��pe�H4m�,��	1I}�����������ؗt�0��A�:�R���\-��I��g��g9��ǓN�0��u�	3 P�i5��Ul��E}r�]�{��\�V��} u��K� �(�/R�~��a�4��?	/h�4�`� C�	�H��Y�Ǌ�mҔ�{��L�H����?T�L�fl�(Kh�iz��Y��[%�I��OAb�Ҫ�i��5�<� i
�'$T����Ȳ��1�0-"~����;jy�0��H]2׶	�G�ˍ��S�g�e'�,��(�^ћ3g��Ih�0�O��	��O!$p��� �*"IdI�EC�qz�x���ʪ	���5CY>��'�)G��� �R5�Ѥj�X�b���9��u)V+j�*EK��*����eG�U�n�KQoD%s(���e�a�<��M7���[ �ǧ�ȃR�Py��!�^B@�
 1CxMy��M��(���6'�>w�z]�WBO��("O� R���#$Jh�
�(�~�� f�ŁK��Ɋ{���IAL2�3�I.s\��c�)C5)V��� X3[�~C�ɹ.�d49���#Lu�q����#�H��	ƓBJ9��Z>���L80p�`�$D��.�Z��ȓh���pr*�	}��)��6l�%�ȓ@z���hSos2��&a�f\��&"�|���_+o?@ ���
����ȓ2Rz'���T�L��
�� u(��ȓ/h�YV�c�Dp���SNh�ȓC�<�i�J�N�� e�
;]0�ȓQR��� YqR����U
�n���`��-c$��j���ځI�$�ȓ<�)��GInހM:p-E�Q�ޅ��M<�0��J W��	jdbYH�L���KqD<y�+	�'V���5��v{楇ȓr!4��dB-���GC@�����8��&ɤ91�!�e`B�&E�I�ȓh>��PN�9�ht���z!B5�ȓ.'<�cJ�2��5!7k�9��!��O$������]��<���O�A�,Y��	%R�Vǉ�g^��3bJ�	�a�ȓ^N�UJg��[�d����('jT�ȓ � =��bE [#:X �o�?>��d�ȓe,~D0���&~�@��f@�K����:-� �,�g�}�P$'> ��Ge��BROSF�\�p�S<3\\��}�s�5E���S��'�E��j̬���1Rz��s`X����AA쌉!���>�ȤcJ��)ޅ�ȓJ�����N
�2B:����%��ȓ{nlM�b�� %���*���8`9t�ȓ9۴u�E��$�����9,����"�'���!琴q���2~޸M�ȓTl���VJ�"G����'nI|�f5��|�P��a��w��ԋ�,]Bn����?�L��	��
gL�^�P�
�� D�|H�i^� Və�}�@��w�?D�����[����xEO@�y*�!�vO'D�x0��W9$�t�!F)��Z��!#�/%D�l(GjXR��0Xi�-��-j�a#D���2���D3VM�n��I�&d4D�����R�0L攡��*3�i�*2D�La�mJ��{eg��xָ�9��.D��jդE�������'=���.-D�dȥ��VD��u.��R���N>D���G�3<��xp��E-?䖸i��?D��c�aݷ]��R,��(��5��*O�(#���:TӶ��@ ��_�P3E"OȠ��Ҥv���r��I&��h�"OV�K1�56J���E�� �"Od��s���Q���ԋH�u�-��"O�<�-\!Prz|X�
Ƙym���"Or�H�B���L���D�4��0��"O���`�)������3�<�2s"O���F�5�*���8L� �0"O��Ѝ�l� �e��$ ���"�"O��Ӥ�]�.-*�+
|m��i�"O�1�s��q�t�آI��^m��`�"O���Z .π��P�Ո%�$A["O ��6
IjwN +�S�`�dA"O�^
���% �c�	�&!�y⣝�a-:��a+���,<ju�B��y���-@t���+R�b@J4�D�y���v�\�����0I� $��
��I�" ��*,O� �@�dN�-<n�E1sƇ��~�`6�'<�Ų2�R9W����M�XuY�O�>#h�I\<���%z�p衧O�M���[Z�'i(�v	�%^r��sA�v�� X*�Q�c��R���$�}s�B�I^l0sF�0A�" �>^W�7��g͠)(vH�[hM����}��M��,K	��u��'Z�~\cA�Rx�<��X�$�l��IW�>�
��Z�҈��M�~m�3M��rG����HOJ� �;��˰̓d���pS�'_�Ւb�4C��H��I����0��jX��)ɯp���I@�NL���Z��t����L�c���C'% �uQ
�jc�P�q���Cq�a���=�hM`�c�Zl$��wC˭��L�ȓ5� ����+�����CٶQ���RqK�{��b0�>	4�q+UJ�-�h����:��%/�4-�ZɗL\# �!�dA�M�<:VEĿ`G�Q�b�P}��t`�aPH�C�D�,�VxCU7�Ԣ=��[zYkcɂ�0ĉ��^��ǁ�=��<�6K��r��Q�r/�l�� "��F�xp��4.��M���a.6)9�
��k�@y��[�53n"<A��,�H@2���!W���JK7��6�`@�&���
O%!�Ĉ>q1�eA5�NB�k"j�����3GC[Q��`���#������(��s �� D�r��F��?����c��t�<��ꂑɨ�CP�ġ���S��.]�&���9�\4r�L��0���'�hO$�y�$�+`�N�i��-b����V�'�lˤ��7^��B�[:/j��0��
R<�ST������[
��}+)s
(h��L��kѳ�(O1�P��(w 8��ѻ D�˟�c�:6,
"P�0x�MG"O���3H�7�^dI��37��I��	�>�,DJ��D� �:,C�Y�>Q?�$�0|T B�.4Ρ�Ȝ�|!���B���F��$1T�G�X�R��rhD����#dL=St_?#=���x�4�3�4�`��gqX���	ϯ`^
��7�T#Q\X	�d�z�:�Aц�(QF�("��U����`^jT�h�N
'�>H�7k'��(���fܠC��)��
4P��1�)D��J�t!� }��)���) �ti��ID�]��ΡNH �K��)�'M0,C�<d�BC�M�:����.��(��	WJt�"�n�3b��t%��*�Nճb�ay2h��T��?2�J�"S��w�!��6<hZ+�<rTLzr��'?�M�ȓ(�8!8�B*W����4��!Q���ȓw�"$��	�����N1艄ȓ)�\� ���/"���y�EO<UF������T`O_�pmAQga�z��ȓ��h3GI|�u9e��>F
��ȓAtJ��3����q�"-�>�ri��hĐ)��ۙ6h�qqC91#D��ȓT}� �����"��?�����8g���?�Q�u��-ȅ�_s� �q2I�Ԫ�'u���A�"��'R�*�F�`奐�������6H�fX������j���J˺"U�]�#�X��E-��'���ȓ ��ћ5l΀$�B!�œ�B(�ȓkS h(�%:LHIF/ϋ%�$�����*S,E̕���	O����|�̬2��B��(�z��E?OLr��XUTq�BHG�w��%�I��f�Ʉ�%8j���i�FH����qG\Ň�IO��2�+�lնuT�W��*���zEtla�i�*;�ꙛ����o׮���!�ʝqS%@�BFf}s��v���Q�Z��'�F-򖝚@�V;h�̇ȓ5�f�i�"L�i#C3d��ȓnR�x��ܠ��!�60U�L���J2����	Jqr���eصHN�H��u��}Kcc�#0�Q�V��
/� ��S�? L�� /��Дpp
Ax��Q�"O��i�nΘE
D���85�52"O��@q�N;�@����G��'"O
$��J�"�d�T�}1"O�0r0��4��)څ*ښ�ر0�"O��C��+����vN�p/�%i�"O�\+�W�	�֬��ښ~�@AB"OMR&�ǁj�P�zB�۱oh�z"On1��%2z�p�{�cܩZ#j�p�"O"apu"ז@�6�+���3 ���"OdX�4�%&\b�(� �s�
�Y�'�y�$�9 &t����.%t�`��'f�}Af+V�z��7�ȅ�t�1�'�{� g��\��	�(&���'��d�A��P4�bd`!�,K�'8�աrc@�^��4�^*�hPx�'��< o��Nv�@���
� "�e��'?d�s׌��:`ī"J�F���'@����א Wx�6�ɬr����'h��l�2 B��D�]�dVĝ��'A�$�@'�<-�T`� �ޡ^�ua	�'�x �%��"|DꐅɜJ!.)J�'�j�['�]
#o�q1�A�ek	�' l�!���E��|��n�A�����'�L�i����p�(�굣��0���x�'@dᅞ:CED	��H�y
��	�'Cx]`��YF�;g�M�4�C��V<�)��E{�S�O�Z���'�� ; �2���!@"ObEQ$;)wةP�'��.	t�R�@��΅�=}2xYӓ&UKG-*��	4f��N�\��I$�0�Be`��E�BD�a(�^��8���t��!�6n$4��臅@� `F���.�;2�As%N1�i��1��� O̜8��I��lAr�f��>0>�`�>b�!�H*�D�`��9ghX�n��0φ��@NE��ڸ�F�y��ʧ	L�dI$x#t%?`ȉ�U7D��ٓ�E>Y^�p"'I0�r���A�O^軕%��"y�(���G�[�x��ЄB�̒�.K���� �+��<��ϖ.J���RB�ڨe�i4� ϒq"�2)b墠g�
l���G~T��N��|��zCÂzh'�<���+ :�VhN	P���
�/�cܧz��ؓ�B�v{��!��0��#6�HID_�:��ғÔ	o�c�AM���CG�)>?N��v/�aܧ��OL��QvD �B�^V�9��~LT"BL�:�F$���,m�e����!����� \6B���k��=���񤌀Et��$��la���Dmџl��Ȓ\J`�m�-N�A�@P�����뉔a�XD�7,[)pAB}i��>��j2��*�J��\�S�4Âè<!��w�X���lʌ&���a�)Q��%�}���0[,e�T�R����HFg�<�@�C�1p�D�Ve�*x�P`p��"pq�'��o^t��g�I�+*�$?��'�)}���)r\��{c�1ra*��t����?�⁒P�&QR D��D�����oޡW}�X�� S�OJ$3��I	��12�G�4�p<�g"�v�� ����h-�9+�x�''�XQ�K�H�b}�&�4�l���L*��E��ȮXk�,C����4�Ro?�,��Y�E�Z�����y�1�bO��(j�B� ��T��l��|�ȣ��S*V�@��e�=	���Y{6FX�Ē�y�i�"��[B�¯cbfQ����X]S�+;"�>�26�WH%�,�I?Q������IY,Lmڶʂ�MV8 W�B�6��䐵Vv�X�ưW�\S@�׻xD��'j�0|/p0/a�H4K:)��#u8O��[Ѫh���7O�\�ȗ�	����ض�P;�~=AQ�	y⼀�JL�Vm�x���?�V񃔍Ǩ&�Hb�'�H����@�be8X��S#h���'�S���k3��z�ԄR-Zٛ�@ް0��>uL�=5��m@G現`:V�	�l#D�|t�ŔB��り��Y�6X2�D�VP��9-��I��	� (&�O]Vŋ��xR��-\Ozl2��o*(-�� ���p?	���D�biCD�4��`R��}Z���lδ`I�$
cA�%�rU��eQkx�� |��ց�X�@1���������60d�tj�S(���휆6:�h� ��}�bGE^�VL(0dh��yRB�L
����샘f�ԡ#'�����g�5�2GV����l�n�Q>u�qk��a��̰�K�D���Zs�.D�t�`�ƃ2�t�7Jɰu�t;�O5j�`8�H�6�^�g̓=��0��16���-_NHx��RM�u�PF��B����Qi��F��"�ݗg�1"��'QP���ׯgޚ@C��qn0��'��H�w���Z�!c�� �rM��'�ĳfC��8#����Bi:�]2�'BL�ͪ���RgI�m	Vp��'L������,D�H�`�Tp��dJ�<�Y`4\0�iӺn�V�Ff�M�<DV��hmx�e�9���ᓁ�J�<�0쓃m庄�t��:m`��z���}�<a i�?Z�� ���>/�)Z�b�<Q�k�"9�y"�Y54h{ׄ�]�<��ɃF�P����6�dR��G�<A��޵s~�|z�nG��u�p$��<I��-����� ���a��~�<�`1פ�aV�0���Z}�<q�c�(�^�c��ܼ*�(0��@W�<�Ƭڷ��)2Ǚ?�>�+��Y�<�Fϕ�Od��"S�@�Q�[b �U�<��n^ �6T��%Úg��![���t�<�tiU1I9�Hc�` �YT6}[��Ty�<A��@��L� )�f8	��@y�<���95�Y��l��I۾�_�<�!��RI��b�6�"�A��A�<����P���Co�h��t�Sa�{�<�G�+`�n��J��:p��ąv�<פӎ.��@f�^��`�w%�u�<�6�˰5
���ғseT��Ev�<Q�K�D�<�,
Yv�=4�Yp�<�Uo����Q$Ǥm�ko�<��'I�y�0��l���jW�^f�<Q�N�h�����B/�Z DOW^�<�#\�x�R�� +khũ�Om�<�e�A'xDBB���&��eqM�<�ɗ�\Le1 뙢]��)g�\�<�k)1ZG�xcx4�T�TY�<����6N���c
*��	��A�P�<a�!��QS� ��e)Bˑ�M�<�3D�l��2w�K�G���փO�<Y�$�	9�nI؃�_�d:A	�K�<9�L� g��@BHW<��ҕ��L�<��nK<W$�Q
	�X`�
��a�<1�ۢaj�[6�8g���2u�
]�<�
����6Y�#�&^B�<aǡM��&��l�0B���K2̀v�<i��B�[))p%`�]��{d��q�<A�+�3
�hi�qaܰ�.5µ#l�<yL��&����A �,i�H5m�i�<���(�}�M��7fACV��L�<�uF�7f�������iI:�
')FM�<�BD�h���#0+�+N�`��GR�<�U��)$� �	�S��D�W�p�<QR��6~|����mZ�;]@�H�Fo�<ѣ园^�r�2EM�pӈ���^h�<R�T�LX�d(��W~6U�H]�<ّ,�.>�xhaL�Ɉ�a�X�<��N��Nx�􋀻lwL�+�aWc�<��dEQ]�s
�(�1��p�<yw�ą}�n��ġ'9��dK�q�<� �=Ѐ�èk��=����`D9�b"O�䋤-�k+Jp��\)�xzf"O����ƶ6������ʼB��C"O���&	�.!.����oӤ	a�"O��pJ]�9���A֭��0���5"OB����il��!4�(�p�h�"O��քI�Il@�dK�_� ,�"O� "�e��J�'.�F�� "O$�&�)= ƀ��b�.3�P��Q"O��Va҇/���r�<�n���"O<�h1���~�
,H )[��Y��"O�Q�v͐�5����B�5�4�(#"OB���{�l��Aʡz�<Hv"O��	����Ĩu���:�$lS�"O�!y�&��o�HaH#6@�0�"�"OR0��0����Vr��R"Ov�QW�%<E�Ad�xB�hG"Oi�{�H�A���6�Vؐq"O�9�'�L�%�@yPm�<f��u{t"OD��*� 3�F�x6M��\Xd)��"O�{&�^*[�d㠌�HF�D"ON�s��\7%Sh|�V���nl�0r"O\e	�؃6���j�G�$F{����"O(�"Ø w���rS� c�\X�1"O@�y�֫+���/�_䔂�"O ���/@�Q�	S �C(}D�"O(�'�=H���#d�5nWz ��"O��K�a߻Z����]=��	�"OLQ('2��3Ck��Def�r0"Ol ��[�.�bJ]�jf �'"O�t� ���a��ɛY�t��T"OP��G�98��,znM?k�ڱ�"OuH�h��sMұj��3"O~q	��Hu`�6���zDJ4"Ozၔ���u$�@pqiD�i@���"Oj�i�'p8D=���B?���d"O�A"YC �* Ǆ�<��$��"O��27��^�i ��\����"O���?!��L�$�K@�4Ҧ"O�H���/5}���wm3e1��C�"Ox�Q��
C=��C�L�n����U"OV����>y9���PACqy<�#"O`��"�D3���O��S��h�"OT��5��)�]HA��K�<�"O�d�E��j���4'^���R"O�d��B�:CA���o�/Xbe/x!��K�>�X�v�
tr�"T#:1�!�_�/�a����?Aȱ0QBG�0�!�$^�fk|�9�昣]�`�c!a!!��l�2�@�]�(�H��Aʠ�!�O1������Z���r��-F�!���<�W��6��s2N�>�!�1S��-���@7%�R����Z0sx!�D�*ޮl�� Q!x�0�P��k!�DY)E8�-��������<|!��߾uZQ1�LK��9���!�D�F�� BF�M�p�ڦ�Y�"�!��J#"Y��\�J��AOS
|�!���R%⌂��t�l�z�/�� !��>.��ۤ��1yL�S��; !�S�h@�쌉^{�9��.��,R!��}"l���M�Z\�A��My�!�$N�؈�c��+k�
�L��+�!�DSJ��Z2���Z��@+M�8!�� ��[ +L;8��۷�	b�� ��"Oҙ)�l34Ȣ��b��&P�g"O��P�%�L24ы�W ��"OD���/
�+�r�y�MˈET詓"ODE��mG�=�.�n_�7�"O��9���O���H&�D���t��"O^x�a0w��l�&(\<���h"O����ZtT������7T�\P`"O�Ա��CX|��H�;;�X�*"O�|A�D�Nl{� eFܺB"O0)�T�$X"��{�/��1��)�"O�,� 	�8򔫴�Wg96�|��)�Ӵk/L@�Έ%ݚ���Ś!i�B�Y�z�Z'�S���4��珍<�RB䉥J�`�hg�>R2�����y$B䉡>lܴ�u�_-�<���O�	�NB� 
�r0��!MV��1Lƌ�B�I�D�P��;���@fI�f"O 1��G��E`� B= @ի2"OH|b�C	r�liU5߸�ȶ"O\ �Ƥ(LL��C��0Ό�b"O����^J����ՆZ���)D"Of���^#Y�lLR N��9j�4��"O��X���=6,�i�Q�ٙ)�T-H�"O(Qс�ڨ�Fmp�8pl��V�	��� �"AT�n�N�#�.f
����������	�N�;$҉��..)H:�XA�x���\S�O���5��V�[(�9�o�,89x�V��J�If��|�>�u��?���E ͶV��2��Zᦅ��7�S�O�F�0���
&��y��،uD5��)���x�!h6E��'ʜ]��Q4�ϑ�y"�d�$���jIc"MϤ~�}��,��s��_6	bdKǠ�q�8��OGP���߻~��	�FG<Y�
�ȓEs5c���!?,���gLL�%��%�ȓ�(���_*Kb���f_a�~��ʓ2m��f��@kX�i1�.e��C�=hMJX���A�88�c�|C�I)u5GZ2�c��r� C�	�j� b��J�u^��v�(,��B���d`�EH��4	�C�<0� B�I�ikB�`�æ~1�ak�6N�B䉢*��Cs�p]ا�ژ��B䉋�V8�,�n-*��ֆV*B�ɮ~BtX`f�Ĺ8��:���W"B�@����t/M����&�W;~N�C�ɺ�[�K�+B�Ⱥ0)�Eq�C䉛HZhɳ"J�	�=�H!w�RB䉘[𹱷cŮ9�t�#B���ZC�ɝ������9~�(��/?PkB�ɔjl��
�f��	���Õ��'nJ�C��$":	��(R��A���C䉯V�e �� ��#5�4?B��)5x�I��K%bݴ�3��J�B�Ir/�@(AG�Abr*:O��B�	#(�m�P�U��!�t*ː<|�B�I�l�� qR\�)��mk��v~B�I�m*��u�U�o!^��r��=�BB�I�jU�ds��I�-�~W�v*�	�'��E�Ū��i'R)۵��Zh�
�'.(s�Ӑg��I
�o
��|�1
�'R���.Y��Rh������	�'�2l1��(ڥA���԰Q
�'���H�ˇ/>瘈 %FE;t���@
��� �H���re<	٣hMe �Q��"O�$��$ �yBm�HӃQ�tTq&"O�H9&c�#$$q{���j��7"O
(��L[,���c��� [Hh��F"O�<���%T5� �@L3E0t!�"O6�)S�E�==^�����%!?F�:�"O�8d(^/;��u/��}	���""OX)؅�sĞ��v.�?dKz�x�"O�XU(�b`P3.��J��5"O$<�Q F��]Ґ�������"O�,�5�ߔ�&���*RQ�*���"O��C����	�mq4�Ì}\����"O*�PE	��q �Y"4���&r�#d"OR5a���Y��D;�(OJj"OdH�Q��P�d��!.�髆"O�%X�ԟ@����a�(Z����"O���GcI<$P�+g	�n���"O.��5��jѪ<󐈐>�z�s�"O��#F�;��Q�Q290��I�"O҅��̓G���ʁ���F�z��d"OzD*�hU7'�2P ���<���9�"O���$甥muʐ�V��f�����"O���@aԉ��;�'2s��{�"O�(�$o��cV@3�JW�� �"O�86j_�)��iw����@��"O @���ӽQ9�%)1�Ñ-�x}R7"O����\�B�V����R.J���#"O��B�H	d4�+�Á=W��@90"O"��b'W�)�=����*�c�"O�@! ��
8  �eBI�Kt� ��"O�`Zc�L1�n�p�
��8$�E"OⰨc*[�i A�0J\��i�!"OZ��@B�(3DA;2�}"<��"O��Yq�%h	C�A��Hܢ=��"O�����Oj3v 2�@��K�6;�"O������g���B��<X�6�i"O��`�	�?��
֧ol�MXB"Oܜc�휧0�P(�cGM�syi�c"Ot;�ᚵWU`D�f�>�f���"OL�cF��p���_�-Ӳ5�c"O^���"]� �	�� �,�s�"O��`�$��wi\"��6J��@%"O�1{�EA�55%EV'F��"O�	s�+�/U%zU�"�H#W��Ѱ"Ox�X��H"���"�C�4)�"O�@��ɒ����3ŉ�?���#�"O.iAa��[w%Y6h�2w���*"O�Y��
�z�|z�AS*T&H��"O(h@��8>�CV!�?8��!Z�"Od�z���C]�t8�	P�0�r��F"O��C����2��T	\8}"�!s"O��*�Zmޝ��Ʈ��PR"O�SQ+�^��=��>���J�"O��1��! �1�Ƨ>�6�
�"OX\�J������Ƽk~B-	�"O(�*a�OȖ%@�cĴEi&��f"O�\�� �-ɦ�`p��;Ng�C�"O,�V�N(}inQ�u�U/-K@�X�"O�CM]/Z�J��o[8.�$2"OvI�Q%��U?�l�W/JF ��"OnyHP�R�x�kƺ ?(�˷"O2��G+Y�T�\C7��;,�]�"O$R��*x��{JZ
't0��"O����G��Pr�p���cH�I�"O� v ��F����a4�[=m����"On��1��6:�����"-�y&"OĈ�R09�tP&�=0��Y�"O�	)q�F�D�6�@�f�X��"O����(R�h��$�>1�y8�"O��i ���x:nM�ctUkA"O��a�g��b��d�$c]����&"OL����W��$�TBO�[c���"O!�R�N�&QBR!�<���d"O�#�
2]����� U�t
��H4"Ov`��F��I�t�s5 ؼܙhW"Oj�TO��<�bd�� �4�(0Z"Oޡ{�NT5馤���_2C��#�"O̽9FƱrQ �s�73,��y�"O��OJ�� ����аaC���Q"O�8{A e���еaݪe'�8�"Oh`(�BZ�qGU%��>�]r�"O(p�Gě�f=@��P�a�"O�)0�F�p��%blO.@jrģ`"O.E1���8�X��Eןe%"O"%�mӇ8.�:���F�0I"O��q�F�%n(�����r�H�٧"O��&OP5=Iθ	Fc]� �q�Q"OT=�CFl�9��a� -���`�"O8�s�CV���5?H���"Ox�IƟ2i�,�c�A�5.�Yjt"O	�ĭM�h	X���K�=y�"OfQ�a�,*���ɧW���Ӡ"O蕸�傳<�h���=.�5��"O�%����5 �N�=�BeB@"Oz�9aո;]�d W��'��TC�"O i0t���R�lBS&͝R��p��"O6)���_6Z`v��SjQ����ç"Od�y�m[�u�uz�
N�^�N�� "OH�K�G������"��IW`� �"O�4�Hܫ	�0�V�9I�@X"O((	W�)X0�L�� B�� "OB�@�Y'e�5�5"J3D'�}�D"O4قR逭h�Ȕ�&��f�b���"OB��gb����uP%�����!"Ort�'�
�.M�9�Aʃ.��JS"OH|A�o�Q!��K����~m�7"O�-����6P��`W�U��j�"Oz
!J��ؐ��.�J��"O�i�p��|jH�)U�X&6q��"O\�b#�
nq�w��;YCrH��"OV�@j:Gj�h5!��>���"O$�ʶ��V�$;$�h\��"ON�xU��:sT��g ю6_@��S"O�1�V��8�xI���O��(b"OzPZ��H�u� 	k �|���T"Oj��*M*���s�jڼ=#~��"O�x7��nt���&Mm�X�"OTp�Ej>oR8��'�k[v���"O@�� �G�����iQ3�:� "O���F�J/i����/,9��؈a"O9���+5�L��}�ZUkQ"O ��nTM��:1�;^_����"OZ!9G�M����b3�/N�"�9�"O�9��,H2+�Z�R�L�uMX�;"O�u@E�֝aSb<�r땬C>B|�a"OhQ
�g��u��,@C&e%ʠ"O���DaH��2Ɵ� �l��"O�@�� �[	��"�d�uѼ�U"O� �� �ސX��P��:�Z��2"ON� �L��X A�\!�"OXh��I�z��\z7��>B���JV"O����)4;�R�n�34����"O��I��P<jZ�Y"nY[²���"O�!�C�	l��=3c�J�#Ȝh��"O���D<f��*�kVf�@�""O`ɹ�'�;a����"Et���"O�l��%C%V^n����8Uy�$*�"O���:m�N�p�ʉ4Ds Qc"Od�x�L֩Z�2�Ǝ��5s@�l"O(-�n@�o\@3ȕiF�@�"Oh�3��^�	�Ua�m�U$$��"Ol� jD�� ��j�g�`��"Ox�8�G
�\�N��l�9vu�lb�"OJ��.��d
`�#����S�rp��"O��tGX���Ѩ�*!	v"O�-�l��N�b���Fy�q�"O6�ѱ!T17lD@A�Q�a�̩b"O"��J�-6�.��ĭt3\r"O��aI\��qGT �!8"OȘjMW�D,�0���=t�Պ�"OR�i�+a��X�@���>�~��A"O�!S�d����Q�g�����g"O~��áҧo	�E�T���L�y"O&ъq֏�¤H3f�(\�@���"ONX��R�T��恘H����"O�\b��0�� ��\���	�"Or1�Ud�9<��1i���G�<��"O����,%RP�BᇔRؒ���"O�(QEBrvR�K��D�*L�"On����Ў;3M�%�:�╉r"O"�s�' ��DŅ�
��x�"O���r���v>�{��G>]��)��"O q����(��9zT#� ���j�"O�k��ΏA}�X�C�'l���07"Oȸ�   ��   �  @  �  �  �)  5  c@  vK  �V  hb  4m  �s  ~  ��  �  3�  y�  ��  �  N�  ��  �  ��  
�  p�  ��  �  N�  ��  ��  ��  X�  ��  �  c � 0# �* �0 !7 e= m=  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- ��!\tu�[�輑��O���$G3&9�IUB�:��ab[93�a}��>�@V�X����Jƍ2l�t�<Y�F�@4*-I��P>|۶��#(�G�<q燏+/�3r+��DGt�R��{�<����^H@��ߵp��	C(w�<�6��.h�$Yg�Z�b���
�g�<Y��0r�t�)e�U�nڙ3fF�c�<�R	�P6H��	N#{Bf[F�S�<)vD9Ja̽1���W�}��UL�<�Z��-���!������EZJ�O�`FzJ|�A�]2�nd��M�� 5�eBz�<��J=(������i[�A)P
EA�<�D����$��/�S���)�~�<1��6r&�0�pC[�l��J�{�<ٓ��9R��@�bɛ�ds�Q3C��\�<ISO߸0�P���E�
֢D��GX�<i
X'&k|��񪀅������W�<�B�'5�p����3*h��K�K�<ɁhP�^V|��B�bخ=J7�EI�<�Q��N�����6F:$:�m[D�<)�c��ZqC�2Ao�!B�aS�<i���<�,��C��+߶QXv�z�<a@n	�/��2�M�T����u�<9�ʓ�JJ9�0���2�h�J�cA}�<��W�{ڂ�����U�z��#u�<�w���A��(2-�N^�x�e�j�<�Cf��Why����w��h��Fh�<Y�mD��ȀY!a��Y։�b�<��`�b+b�;��Ԍ���Śy�<�U�ߝٖIhG�Ol4&hyP�j�<��ں ��J�bȈ})�P��i�<��T<��QӇ���x��!�Y�<����I�J(�a��8v\��g�X�<��Ϣlk����#�!�ų"F�Q�<�M��2y�HS�B;V!��IMB�<�A#U�~�ˆ%H�,1�%�%fg�<	��	���={s� =T�X��a�<��N9`5��:F�}�X����Z�<�(�l6����W��D�"��	Z�<)+,��qhq�kj��B7B�T�<I�5r8a`���0^�"�ăT�<Y��Ę3NxH�%��$Df�2c�W�< 䁳	�~iX���A"�8�fQS�<Y���X0���nU�z� gFP�<aҀ�V�ȹ�@o�.�@��s�<��*ɕ�&��!%�p!3 l�<���O")�H�b�̳}_M�q�j�<A͈(�P3�bK�S�-���^�<�3KA�x���:�`A,���P��b�<Q�#��6w�i�
@i� �rA��"O2(��K00n$q��W	|=h�"O�iKvKW7�� uLR�w�s4"OP���j޷����C+�<[Z���"ORh���r�0}�
�0Y�v"O� �fC�oW���D���d�"OF5z��P�e�F���Ν&�4�h�"O2����F/��C�)�R����"O��y�E�5Ai8r�_�N�S�"OA�GP�=$N�Q�gFP�A�"O��J��׌T��0�Â_B�ɩu"O�C��ߛNӔ�ۑE �l0� 0�"O�Qp@�&)Y��At��F$�ab�"O�@#�Ճ4[�ո0͇�[,�@�"O�2S"�c%���v�;�p2�"O�,sҨP�V��q��ꐸ+ �3�"O��`�Ҝ<���X6*�V��J%"O�0�a�T�y�4uB�
�)!�ڦ"ON��Q�R����"�[�1.њ�"O�h�evAޜ�`n��*,8��"O�,*��޾?:���g�[�H;��1"Oȸ�#���1`L]�(�ɩ"OکAS$�:��0D��L ؅"O�a���2�����[�`�h8ѡ"OЙ87A-������C�E�bTzW"O@�Z�J]�I�N� 1)T��"OҬ�����tR��PN�@���"O�0(���'�8�RK��(���"O2��"c����ʇ!;����"O�Ŋ嫞��4ГC(��Fu����"O�A�â6����G�Ca$ �E"O���ge��x�6F�&D�"OzѠ�fT;n	6��#gW9$*n}�1"O��0P�J�ܩ�3�V&.��R"O�呶C�Cܜ����.	�H��"O@��W�޼*�`-��S�|��"O�a[u��!#����7��B�t�t"O~-��D�#~6�Ғ��?+B��"O(�h�4:���*~p<�"O(C�OJc����VǘDd6�� "O��	Ϋw�ne8 fR	<O๸�"O\�q��p�T�q'
dKP��"OD�	`m[��r@S	K&<J08{�"O�-�%i/#��a$��Ct4�!"O��2V%F -&tt�$N��C"O�x����
#���4��=�$"O���*�y`���3(����"O<�`Ƥ͓~�ڱ��$_ִ���"O���"V�>L0ƕo`�k�"Oz��L�g>TXR�� `r,�e"O>�1��T�c����(ҤY?b���"O�@S"�
;)��Ic�Q�6�{#"OP�ɓ�J.%��9�c�n��4"O�5#�® 2�`�@e6�%aS"O��k���?�A�-@|.�`B�"OX�Ju&�z2�Y(+Ŋ6���"O�1��f��d�w	�eo�#"O�H��$UM�xVF%�-�7%o�<QՠϜE�`��-߀Ȼ��V�<�3��#}u}���:��y��ARm�<	6�_��ac��,F�q��i�<$�I� BHÖ!L[�1��+�^�<�@��
;B�c��� $�EnCf�<��I�� H*T�&�ھN x�t�Aa�<�'���1�e�R�W9�B�8DI�<��.ΈHh��f�3B�fthgnI�<!�Z7ƕ�B
,k�4�³�k�<)�	ޅ(��-�᠎�L�"�*��Og�<�AҰ=����1#ϫtf��pS��f�<� &�{t�^�<jV�k$�
M$�(�"O�ٻ@��!F6�`�	�0�i$"Ol0��U�]�xQт��k�4� "O�� ��& +���_�D���"O6���ɽI�(}jƌǆs6�/�?A���?����?i���?A���?q��?1�Ǻ �EHQ�[W���P���?1��?����?y���?���?���?A!��`��:#��K]�U$E'�?���?a��?Y���?9���?I��?	�M�6"������U��I��J���?����?����?1��?Q��?����?�B�*60�q��W 4�@@{�A��?����?���?q��?���?)���?���UE{<y�T���h�H7ȑ �?���?Q���?9��?���?A��?�����h��I���%iQ��[vj��?���?I��?���?I��?	���?��L��Pv���P�%R���hU��?A��?���?1���?	���?����?11�B#(��t�T�ψ'��Q@���8�?y���?����?	��?a���?��?	%-�E:li���!-(�rs�@#�?����?����?I���?A��?!��?��EM��H��
0]~(��"� �?)��?	��?��?Y��?���?Y��A8>��xC'�^���lC��*�?���?����?���?����?��?i��yv  �-C�j��@v��?i���?q���?���?�5���'7�ٯz�0�C���#F���Zf�߽(#���?.O1�����M�P��k�����E&G��1�KCc�2��'��7-(�i>�ោ�f������Ћ_�����Kȟ��	�/��mZD~b3�(��Su���*K�>`4,�"<aXس�2A1OZ�$�<����Xnm[�̑�:M��!'�V43O�elڙJ�c���:���y��l��A�$G��5���� ܾU���'g�d�>�|� L��M�'lLDB�BQ�f�,�Sl�&KP���' ��؟l��i>��ɫNAȔ��E9�HLS!�!u���	Iy"�|�`�jX�V�(�D��M �v�e@�ۧ$���(��OZ�D�O��e}2G9���
D�1[�h�V�Ӑ��$�O ��Vn�'!�1� ����!���d޽6lq�$�K�sh���fm�:e�˓��D�O?�I`�F���*��P�׃�͢�I��M��X~�cyӐ��(���@:+G? �X�'���'���˥V����ϧ)W�$`[��5�q-ՊZK�H.�X����a�	ey�O{��'���'�2�Ѿ���c4�V+(]`)sei�Z��I��M륇�+���O������H;Y�����섋,Ơ���'����'�2�'*ɧ�O(������&(ؖ����%y�䌣an�z��E�Y�d����L{�IGv�|y򇑣qw@� զR6ݐh��
�qUR�'Ur�'��O[�I3�M��ɉ��?�ϖYl,��hY�H��A�*�?� �i��O
d�'�b��y笕�r"�ܔ9D��e��F�S��i��I�mLi{�O��&?!��4L_�3b�8s��Q[�*�h~��I�$�	��d������	u��u�l��ɦE7�$�q����'�b�'
7-3#��˓L<��|r��%?|,k�
ߣXܶt���h5�'\����� )뛶���]3?}j�#�1{J)K��4�N9�����8���|�V�l�I韴�	ܟ���[(��rBD�n�8*5�
����oyB�|Ӹ@y�m�Ot���O
�';�NhӴF9ix��`��;9�H��'� ��?����S�T��;U@�*�L1&6�Ay�������#2(�$83�O�i(�?!f�&�=J��#�S�X�P��N�	4����OL�d�O���i�<d�i���� R�(|���7��.e2*�X0,����'��o�n⟸��O���j4b�`��r����4j��@� �d�O&uxc�gӒ�Ӻ��,��4j�<a�@�yR9fl��m����<�/ON�d�O���O����ON�'VKF��秜�8ت���Wd�0���iH�z"W���k���h�����Q#�N��L"���(w����戝�?����S�'X�.���4�~"<��C aM�h�4��!V�<�#�̾����?����<9�S��O����C�	��Da�a��G�y��'u�⓫YQbU�<A�4�*4����?����^�S��X�$:���'���?q(O��D�Ot˓�?���ǈ=<P��C,��u����<9�(KX��1B� ;�TA�'Q�4C�ៀ���'�$ش�R%#4�1�RL`��Z�'Y�	��$�� �.�(� �>Oj�iC�'wv6-T�*$���O�8o\�Ӽ;���&> LY��$�eSv#�<i���?Q�E۰X��4����e�V��.agR�Xz�ҩK?i� �ʢ�����$�O �d�O��D�O��ě{�)���N/
��,K�)�Tw��'��&놝O���'����'��5�B��=%��m�fjʤ	��YGY�(��ğ\$�b>�3�,�!{:�&�u�|]���O3�Y�.?�4��g.�d��䓂�d_�JU�%�Ѓ�A����FH �`���O��$�Oj��FE� 5� ˓U�6U��DbD�%���e��]X,i��OƂ@'��}�&�$�<1����I�����˟�	�'���]�A��$�����k���l��<��g�({�/��'����� �T��`P�c6���@�JQ |� <O�D�O��$�O��d�Of�?aq��j�J�3r.ލ'�(!�f��֟��I��0h�4B��|̧�?�״i�'����呟JJ�4Q
��Y�ȫ5�|�'��OBB|��i���"!�.,3���Q��P�p	��:�(s���1p��"���<�'�?���?�� ��K`�
:P��F�?�����$��	��/ Ο,�Iޟd�OE�!D��RS0L�??E�Y�O8��'��'ɧ�I_�R�����@;K�*Qg� ��5���?ܚ��t��<ͧNA����9��Z�b��M\6{���vI3� 5s��?i��?)�S�'�����2�Ȏ%��a�CD
�|���2��؛�� �'�7M7�	�����O��a�h�
�����!m��)�
�O^��Սj#67�>?i�H56��	:��n�UI���A�)+�P��
&�y�T���	ɟ\��ٟ���ԟДO�����f�D6�k-7��۷b��9q���On���O���j���ަ睜�R���C�<L\A�v�E�R��I�Ia�S�'!V��a�4�yR�JE�Wο?]�Y�$�r!F�	i����'MY%�ԗ'W��'�(��0,V$@����O�_v���'���'�"W�\��4F�`���?Q�|!| ��[}6�Kv*��<|$ʏ��>����'m��Ȥ-B�<s0�Ɇ��K_ҥR�O�`��m�;�"�c�$����?I��O:@�"o+�n��1�O�y`ʣ	�O8�D�O����OT�}��B[����iO7�	[c���r�A��uߛF�Y�a��%�Ms��w��@��N��,x��/:vL �'.��'�"n ��Ɵ�X:���������$h�h�r��a$��M���'�ĕ����'HR�'��'.$e��J=,�@ rV�O�LE<��Q�۴6��a
��?1��䧎?Y��#M��Y�&O�I:��@f莠Ld��ҟL��r�)��0e����`*I�L��1����y b��'�|$�B��(���|�R����O;X�$���LZ�	��Ze��<�����I����wyb(j���d��O=2�(R�x�|M�A��'K*�hG7OIl�m��N����T�	� 2⒍Y�ry�B�0�^��׏׼" �m�t~��^2^
����yܧ��s��L0l���U��x����<����?9��?����?Ɍ��ۙ!;��k��N�~d�*�%��S���'��~ӆ�ad:�|��Yߦ%�	ǎ�:L[6Ek'�_f��6&.�I� �'��S5�i����p��L0�)n����>���m��d��ɚ+��'�	�`�I����IC�*�·J\s�=)&,
1�>������'F@6�PG.���O��į|�Ջ��%�8irճ�8yd�}~�A�>y���?IJ>�O�
�+��Щ %f���*�� $LIH ���R����`�i���|�����&��WfS#����oŔk���G���P���t���b>�'�r7m�P�q�U�*��B�F;oK6�9נ�O^�����?9�[����&M"����荟LE����*	�X߈�'���V�i#�	;J�����O����'�2�r��Q*i（(�gյ,N���'��ߟl����|���$�IA�4Ϛ�2d�!82lQ�b4mzp�ӁA�(7��F��D�O��>���O*Unz��T� 9(I�����A6�&%��,����{�)�S�t�pqn��<qA��}�Xa�"�+a(H`���@�<�Ч�n+
��\�	vy"�'4� F��ݬ�	E��
����'���'N�S�P�4%�L�j���?� �,��рۑ"\4L���V�Р1��k�>����?�L>�ըB�6��=�r���<h��O~2�=<�*�ˉ��O1>��	 *�r(�/=�^�yu+`�ƽ@P�&���'���'�2����i��OOf����b[�{�5��ޟX�޴HXhC.Oʘn�U�Ӽۗ��
p�		g!W���0&���<����?a�(��c�4���U�4����O�tyF�:��h�C���|�S���	ԟ�������@�T&�=a�d	�BU[f>�â�CHy2f�O���P�' ��'S�O#b��06�ؠ�ӧ].D�ɐ ˭=����?q������:�x`@�	QMx����~Ǧ���GA��I3�-���'m&�4�'�&h�&V, t��µw�8����'02�'Mr����R�ܩڴV�@���,Ϡ����t�x;��"1���ϓe���$[F}r�'��5���H)��i��[���i�6};6�X�yɛ�����T��7y8�h�P��ߵ` ͉1W����w�!_(��K��a��Iٟ��	�4�I���0���2��2E�,p͔]�&Y��?����?���i4����Q� ��4��&O��{Ǜ�<�&%�����+J>��?�'���ٴ���ɓy�� �q,�<x����錸5�`�Yf�L�~��|V��Sܟ��ݟ�`&[!#୰cD�-K��s��ßL��Fy��}�xD��-�O<�D�O�˧i�0��u�БNT� �e�H��'���?����S�Ԇ0L,@hR �?�",jU��Mo�A�d�ƿ^P���O���?AW6��T�2&8q�!g�6��t�r� �D����O��D�O���<�4�i/$`p3iE-h��y�I�(.j�ĳ5�7��	��M�bI�>�@궈���%m��B��]�J���?i�g��M��O��%o������� P<97K�5dLƩ��],���F7O�ʓ�?����?���?������̕��P�@T��z4B׏��Y�Tl����	Ο��IX��Ο�i���S�A�-"��X�DK*0���6��?!����%߹u��f4OҝJ5!@�bK���ůT&k����4O Ě�$,�?��&#�D�<���?)2��5s���F������?I��?y����d�զ��Uň�d�I!��Ԙ�Py�c��9� ��&#�Q�2�������In�	M"�F��'��Mꂪ��."�`Ov�s�� �M�Ð��%�l?)�;�@�ҊH+��e˥c\37<&t����?a��?Q���h���$�^�3�(н�b�3�ԭJ�������Xퟐ����M���wGF$�$��?X�a�g�+9ǜ���'2�_��8�OƦ��'x�a�ӌ�?1��$0A�D����A G#�0 ��ُ�'!����|�	�8��ߟ���?sW�AS���?>i���C�'N��'�|6�N�����O��?���O8*$F�8�2]a���%K&q�CCa}��'��O1��[�	'����ٚkڮU@��:�P�h�D�<�V�=kX��A�����<y6��3"l7��R��V������O��D�O����TQ�@[�4S�|��D`��ǝ*�Z��)�8m)|�� *�f�DJH}r�'���'Х��G�� x���k��u��1�n[&{�����'F@�t�Q>�]b���r���)<ѺL�7���	쟠��ݟL�	ğ���`�Sݟ��3����B�:%�D�����՟$�	ɟxC�4b4Z����?A��?).O)r�&�uO�����1�D�O��d�Ojq��u�:�I��8R��#5̥��FʁxAT���ӂ4�nI8�O��O&ʓ�?	���?9��q���ѤBwq+��Z�>�4}��M���8��syR�k��M�է�O����O2ʧ	9�5�˘z3bG�U�`�'����?����S���s<��e\�Ԍd	�N<Y�.�17��Y9�֖������:�DW}[�V枋VZRH�"aU�t�!��Ԧ���F
>e�^d{�@ʛf�.\��$Gh���I���1�4��'c�듸?�f�`����D7|D(U�M��?�d�T� ܴ��D؆GX�
�O�剺r��!¦H=B�0��4��	Qy�'\"�'rR�'"W>]a&�� ����r� :%��x�#Y�M[Q�X����O������	��]!W�*��FB���̊�V�~���y�?�|RgDł�M��'�TC��r=�=(0H�)و̢�'a��)gC����|rS�D����xS�$J(!#�A ߂C�D����� �I�����ey"`�b�0�/�O ���O�@��H__=��k"oR(A41pA�(�	���D�O��d3�d��{>��3���Q�p`�-j{�	!����)R�E�|��O����	�}�� 9&�ۭEDpPiBDڀ,H���ן���ҟl��l�O�RӺHe�T�%6j¸�R�J���e�<��U-�<97�i_�O󮈔84UJ�9����g�>��D�Oj��Od�JdӤ�4�~�a��?�	Ç��#�{�D�E}��Z��Zy���y�/v<X�i�-���Ͳu������) �ğ��	̟d�J�&�"I ���!gĉn)l
��ʓ}d�	�t��@�)��b�>��cD�&�"Q'ݥ��ȫ�F��a�.O,u�d���~��|b^�pd�C�;����"��7�ժ�jA˟\�����	��iy2�e�H�Z�`�Onh%�<60���	��#�v��V��OV�o���\��	؟��	͟�`���Oמ��b� � <JG��!!.�5mZI~�(�w?<�'��'��S�P��2���j�$>�d���N�<!��?����?y���?���dj��Ա�i�9�B��r��):��� ߴ���O�P7�8�dR�~"̩��꟭
k�Y�&3~�6�O��$�O�U�Z�ܴ��DR�i"pM�H�#!��hA�&����E�4�~"�|r[��ԟ��	�\i��R=�N�$*����y5j�۟��qy¥}�\źQ��O����O��'#]�CD�Z��t�؛$Ft�'5ꓔ?1���S��)_�q�J�r&�@ZlR �W�<��7lW�J	���O�I�.�?��-��*,RH�P�Q*�]څns�����Of���O���<y��izz�*f%��P���Q�P/fnh�'/�&bT��"�M#���>��Znx���z���� W�B�����?1�
;�M��O��Cf$#��M?�q5�����3�հ'"tPv�`�ԕ'���'g"�'�R�' ��L���K��Q�# 1������Y�޴6�<1
��?)����?�E��y��T�p�����1��H��^"�B��)I�$T�7Ml��:W�
�9�ha3��	9oJ�Q��h`�����4"��Yg�ty��'�r!�2-����@��(&;Vh�y*��'7��'����M�r��?����?I2��F��-I��H�H���B��7��'`��?I�B�"���s���]�8ö�%��9� ��I�x���(0��K����Q5T2|�ve�1P��$*˖7J���O��$�O���7ڧ�?�g�Ϡ��D��*��/�R�����?6�i�Ԛ�U��kܴ���yǢV�D�a�J�;t���pI���y��'f��'���5�i[�I�m�>`���O[b� ����03���$Ǚd��b0�>���<ͧ�?���?���?��I�|5�(z1K�ص��Z���B��Y�������I���$?��	�%�X� "��6e�3n�]���O0�$�O��O1��{'�{�v�`�� �P���q$Iݮ��A�Ǚ�4��K�8]r��N�Iyy⍝�|@�8Q�J,2�l����ʈa�B�'���':�OW�=�M�©�0�?i�MR#'�ܐ��KȚ|S
4�I �<�R�i��O�x�'9��'�bd�vv��	��E:bA1��E�&jp9v�i+����HIP�O~�d%?�]IV�t(��!JLX�F�?���	ǟ\�Iɟ���ן<��m�'�Z�aԋӮ*Ҥ쀅+�,��4a��?���A���h�	&(�ɑ�MSL>�q��,��A�����Z������䓚?���|�t�ȥ�M��O���|P J�4+�H��� ,c�б��O � I>�)OB���O����O&�ʃ*��,6�����=d��5���^CWpd2�l�<i��i��<H��Ox�'��t�w� =那��6�`y�OZq��Ә'5B]���IП�$��� +4k�*�f���H%Mr�X"���B�fEѲ�"H�0p�'��t� �P�|2�7:V^�pvA�0}���qUne��Iݟ�I���)�Sdy�Hm�$d��nٔ3� �%/C�LU����/o��d�O mk�	M��埴+B�M�Y���r��G�-� �q�)Z[y�H�:9����0���
(6�T	RNy"ş� `��0S-C�*3T���3�y2V���	̟���П���ğ��Ou����eU�C<=�Ū$�B=���wӘ��c��OX���O蒟Z�D���]!x�1��n�zܒ��3%ǲt����	۟$$�b>%�����)̓b:>dÉ�eB �A$��8�Γ1�8a�@����&�|�'���'y�P�	�*���҂��VB<��'���'��V�D۴j;�m����?a�{@��B ��&Bʩґ��^�ᡏ�ʽ>����?�I>�ԩ��(Ǵ��I�sQ�+��O~R��x��h 5K_)��O��x��++�bΖ�\����_.X�Sg�źZ����?����?���h���D��Hh��_�b����`�I�U42�D	Ԧ��2��_y`cӒ����qA���-�:1��\ )<�	�'#�T)s�i��I)ȍ��O�!�oX\�|�I@M�>
`��"�B@�^y�'12�'*��'P��05��Y �� )
��0)��.�	
�?y�o�埠�	�@$?�I�npt��C�DHxs�m@d@��O���O��O1�PY�0��;n���S&/��	(A���,y�7��kyL@j��u�����dN�p�[G�����"ƊT��d�Ob���O&�4�"�N�v
�*pR��$~� C�^������r�q�f��!�O����O��R�p�|�a�!R=C����T�^�77ؕ�D�h���zM����C<�'ȿ{M��K�	�i��T���(���<����?I���?y��?��D�7;���t�Ϗ9� ���-0i���'rOhӨ� 4=�|��ݦ�'�|pP^�A���zF���>D�A;�-�E��@�i>a������'D�g��~<X�0���l���qg�U)0�����	S{�'��i>�����(��%y"$M!d�	&�\��3�O涘�	П��'F�7�σ���$�O����|RS*�1x��2�X�*ȈTҧK�T~Be�>���?�O>�O���&���&!�Ď7r΄���=l"`�d�����t#��� ���|�e'�CE��b�fe�
H�'���'a���\����4H��� &g�5�*�h@jR�C����ƍЋ�?I�
���� i}��'~�iJ!͜D����2a�&�9��'�����l3��,�q���k��Y��)�g`��c���2O���?����?	��?q�����V�� �@P��M�ұ�4�Y*V�mm�l(�������l�'o�X�];������.v;tES'��&�dE��Ο�&�b>=��#���a�1�64�r��V�%3�+W,$(͓)�L�!�N��d%�������'G|�p�H��� �`�T�)���'8�'�W�(�4<#������?9�j^j�&��m�6���ۺj�n��r�>����?�L>AE��6'�68)�@�H�ZDs4j~~r�<zh�"oTI��Oll���I��g�@e�p)����^^ykR8r,�'H��'%���ߟ �d��$V��T��.Mzh�;#���XX�4jp&�����?Ѷ�i�O����$$�&ųAު KA�\�0g�D�OR˓H}b<�ش���
��� �'�V��%7x�ꍑ�,�N
��;�E<��<���?I��?����?���J���򦜬]���(�ED���DL˦��䫄џ��I̟p�r��.Qb4��%)����A6nk�������E�)�S/@��yh%�ƛYh�Ŗ�pu�8:�Η�}�'��mr�z?qK>	,O�i(�K�� =a%�E9{3�@آ��Ov���O���O�	�<�q�i���XD�'������3�`I�#�U)b����'/�6�7�I��D�OD�4�� a쀩\,�XFf� �� ����7�/?�B�6)>F�iV�䧣��f�*}��)���s9\�+4h��<���?���?I��?����H!L�8���:�wbW�S�R�'2�p�N*e:�������U'���ꃷFy�H�Vm��ͫ��P[�	ԟ��i>-�JԦ�'d��� �4�p� 2l0����B�$��	3�~��|BT���ҟ��	ޟ����6?Ƅ�$^-3o��ە,D㟜�IXy,Ӛ�Q��O��$�O�˧BQV�h�h_�B�N���K�;d��'����?)����S����>�ؙ�2�^rֶ���E��X��S�2 �q�O�iM�?)��:�d���pd8T�&E���ak�5�����O`�D�O��	�<	Ǵi� G �4sf���
2S��X*�E	�pB�'�6�8������O���#v��3w�['t� 0B�i�O����'7{�6m>?A���7���>�R��� ��m�"AÌTr6,���q��'2r�'nR�'��'��Srw�Ԫ�k��4
t�3���v��1ݴ~I8��?�����'�?e��y7�Z�Mx�P���з���5#��'�ɧ�O8H���i�$��aR:̛p.09��5��ČzQ�ü)����'/�'��˟���1K� ��G�Ld�sg�T�Z��I�d�I�0�'�:7-��d�OD�d�8�h���#�}l U���㟨�O(�$�O|�OnE��ď1nB���aլu]0�H'����7.CW;bx�1!�S�W?���x�*��^�@��f�'g�J�x�Dݟ����|�	Ɵ|D���'V�"Ǎ�/"��G�S�><ۣ�'��7���]�����O��o�y�Ӽ�Ӈ�:af�lx��8K�h��F�<���?��*/8��ߴ���R&z=�U��O�j���Ҟ1��	X6��`� �p�|R���IП��IğD�I䟤h7+ �P�1q%������`S^y��lӔ̂�l�O���O쒟�$�A��ZG�!i������� �F��'���'ɧ�Ob�X��
�?��7�@��+�f��K7�V��<���T�>���IE�_y�C'c�р�Oٿ:��#eD�x�R�'�r�'W�Oq�I;�M��
<�y¢�f9����=`�l%���d=�d�̦y�?	�S� ������ɡ|�f�r��4p��Y)��8�.��覕�'਺0	_g�L~"�;̘��7o�/$a�0a���̓�?���?Y���?	����O���i��ͳLCp��c�C����'���'	r6�I���i�O��lZ@����)q�[�tK��9Z:[��$���Iڟ��VR�oe~�C��i��\s�Fs�d���&b��H+�	�t?�I>�,Ov���O���O�0(�H��68�?��lYF��OF�ħ<ђ�i���K�'8��'b�Ӥ/+�5� ğ?�z��%O# P�6t�I˟��IQ�)baoݠeT�e�1bM���iц���RZ#b���4.ǟ�ұ�|��N&�Eis��+�]��I*H��'��'���$^�\��41����V�������+�6,���e�V��Ą��?��[�����@��M����R�zץ¢AE���I�|C�m�ͦ��u�
��t��pyR
�!A�2�A�0T.�ر�떚�y"^�����p�������Ɵ�O~zd�P9a�^�I�:aK�̜�SD�6-֕)&j�D�O���/�9O��oz�1j�Ň�>�L����Ϻ־e �,�H�I[�)�ӠL�
Qn��<����*�B��A��R٨�˅�<���Q��>�	e��Ny�O�"i݀O���D-˫G۔+`I�>?�r�'���'��I7�Mc�h�#�?���?1�'RVi�%S��7�)Bh����'W��?Q���j��4J��J�SUD%0�l�q�'��XJ R;>��}����!R��T�Q�'�H�a��K�9�BnA�n!a�'���P�Zd�>�3r%��Ș���',,7�vG����O$Yo�K�Ӽ�5fǘ��!���?�ll(����<a��?���K0i��4����";b)��O;��	�,�8�<g�O�4XA�%�|BY���I��|��쟴�	՟���B�;5���ŊZ *?��x�G�wy�-~Ӣ��C&�O����O������_�|��p!�P��s��5�'i���	���@Aw�H�k�u���-h���#�v�ʓ|��]$��O��2J>9,OW'N �H����S!t��*���O��D�O���O�i�<�u�iD��R0�'�d���)C��N�{fb��WE ۜ'�$6�8�	�����O
���Ovi�iu/΁��K�0{dDe�Z�Ң�iE�	��E����5�	��\!Z��	�|���7��4e{�eZ5O����O����O�$�O��?]���t: ��֘)E��ԟ��	�0 �4)�ͧ�?Ѧ�i�'�BQ�P��C�>����
e���ѝ|�'��OPX(�V�i���PT*0���Z�
���k��Y=�f�xX�<���'��'��o�D�dQ��8PD���Ef�'$��Gx"'}���!VI�OD���O�ʧ5�-0� ��xa.O&ms8T�'��?Y���S�T�� [ƹ�DMV�ozT�$[��Ή�&
�\Gdݨ%S��Ӟ)sң�^�ɿN��3�l��dLq��Bz
B�I��M�c&_X��1��'��s.�Xp�#7�Q����?�W�i��OԹ�'��L]�u���`"��!7��e�tB�+f	��'B�X�i��iݭab��?M��V��9��ٯ8X�Y��L�Yx�x��x��'r�{��ƴ#*p�ЍS�,̞u�� ^�[��6m�75����O��?�ӆ�M�;H�b�r�&���qh�E�7|����?�I>�|����M#���  jCd����1@�T��<O���s*M��?�a,�D�<+On�ȄJ�:($i��	e�ѡ��'HP7�0V����Ov��@"HH�� ̹o�Ny�nڳ��#�O�$�OJ�Oz8�V,�vހ�RU,Sw��UH���٥�X$^� �mZ���B���3�F%8^�
"�>�beC�I�Z2����I��X�ШP;JB�4
d��&M�|�Ȑ!�0�2�d�L�vj4�sWL	�2e��iU�Y�a	�!�.�x��k��y�45���3.�~�:���+}�"�p�R	�����6#H���$�B8rE0�B�#R�f���ǎ�Z�r�C�U0\m�E�� 4���I"*s��CU+/t8�cS�պ�����/�eR�7(Y"};�Î ,�0[�R!;\h,#�D�,5Rt�I) .������	K�y F-�+]�佁6���y�	�h���`�Oʓ�?�H>��<�<q ����� ��Ï_c�$�'���Y4�|��'��'��<@3�x�$�� I�L�-�Q��c��4H�A�'�֟�'�h���<)�m��%�DAk���q�Ѓ�jq�b���	ПP�	TyB�ڙV���E�dS��#�$�$ÚB0�7-�<�����?��|����'�iJ�̏�v�6�W�@�st��O����Oh���<�'"��t��؟lJ� ɲU%��BDe 7pf�sƊ� �MS�����?Y��[-���{�ōwl�a3K�" �a�����M#��?Q,O�%f{����e�i��4��)����q*��-�l��*�e�:O��$�OFL�r�1�	|�7��#)g,�!3.0��hjb�V�U�'�n��&)s��$�O.�$���h֧5��B?1�1�#��J|�	�2Y�M����?qV& ��'�q��P�4a�L��򉌦A�JL�ҷi����.b�����O����|���Մ:�,�!��4)�����@�W��am�Y�z��?���D�'���ȟ�R&BYQC�ІVm�1esӘ�D�O
�����m�''�	�t���l�2u���V?`��&�K~�Rd�>Y$�Hs��?���?�5�ɲ7Z�H
'���)��j� Q����'���i#n�>9-O��$�<1��〃	� `�K[�����ݵ}���+=b�M>����?�����4�h���يa���.5�0���}}BV� ��W��$�ɉ'���{!F>y,��c��ͶBjA�������'�B�'��Z��Q�.���bO-��R�dS#p�� ��'��M�-O�d5�D�O�$�
<�r�IX"%��DV=���c`��MU���?����?�*O"�Ъ�s��'#�� J?l4H݋�`�0d�n��Dy���"��O�d-,���j~�$�Q��4B@ȲdDq�(�$�O�ʓg���0��4�'�\c�6�A>*�lAҴG��VhȊH<�,Ob�$�O�����X�2b�9ߊ�����G�P�i�iW�I?}Inx�޴d`�ܟ�������_���p�##��X�s����F=��R�(�	ȟ��I|RH~n�8�zQU�S,��P�kK�M5�7MH3|��xn�����͟(������|R�j�:t�CL
�r�5�5�#`��v�'R��'�ɧ�9O��ĝ�''�E�C�g���b��90.�m����؟0;�%Ɵ���|b��~�ǦZ}�<�4�o���(p�%�M����]p�3?���~� �a/¤#��9H`*��� �MK�� EH|�(O2H�O@�Ob�D�S.#Р8�ګK����FS�
(h>b���Ayr�'4�eW�Ö+��Ju�8y��!P6l�1q��Iߟ4��`��?�'�x;]ʒ�	qΒ�b`-�u��Φ��Rn;�	�L�'��AQ:k�����"EٶL�5<���ԋJT+���'�����OTʓ+�d%nM��#�U�d�L��fY�a�.O���<��E�� �,���D�xh�HH�E���@2-գ{J�lZ_���?�+Ot|�Œx�oT�X^(Rt曱���x��ƌ�MK����O6Q!%��|���?����6�D�1q��
WT3D�$�B�I��'�ts���~�#� �3�( ;�&��J���_���ɫ7�a������	ڟ�SvyZw�2�yë]4A��1�K�(/����4�?�)O��B�)�I�#r�܀��
ȷ-��	�^휠ny0�=��ٟ�Iӟ���cyʟ��:o��R���YE�w �в�Bg}����O>����6�6q��I�<w�us�͞��M���?���O�)O�]��36��`�ŸY{�,I����~��Dx"�-�I�OH�$�O<�"%���PH%�Y�r�S�$說��5A�&�0�O���?9)O���Ƭ��f	�L�"F�=0�v[� ��e���'���'BV�X�bƴ2�&Ps�!ȉ!�Ҁ󵀙�Dd�0�OXʓ�?�)OZ�$�O��Dܵ$��(��a���Bt����2`�F��d<O&�d�O����O6�D�<��埫e!��G�a�XVDL�L�@T�MR����\����Yy��'���'G5!�O%�2IF�"0�dM4	���IA�i\b�'���'(�		,�����F���X   Ó#V�Ԍ��!ϥY����$�ia�[����矀��@-b�	�t�����c0+��+���C��ТoB�anZߟ���pyr��w����?1����3o
@�l�恘)�L�s_	++��ПH��؟�C7Gd�(�	ԟ��IU$E���XC���L6�	�5d�æM�'*D��Q h�
��O��D���	էu�ч+�,��c���]̀$c!���M����?���S�'q�� �11)3e"�y��+::���i��Ph6#d�2���O���'t�I�I�2l���5� 5i��ھ� kٴ-ž������O���R�mR�C'o^)��a
�i��D6��O����O�l� #]H}"_����~?�R�#S=hU��͡
yt��.����Imy����yʟ��$�O��,�X��5JՂU�8� ��^3�6M�O�����T}�S�H��oy��5�A
3ي���՘&j�֛�{��m[
��'�R�'�R�'��	J�,P�NϰPJ`bB��a����B�����<����$�O.�$�O����Y�o���S�H-��:�`Ք$A�D�<��?�L~J�Â!P��E�:�:�H`.[(
�q1�����W�\�IOy��'�b�'��Ș't,!yb�#@���V�PE���p�s�B�d�O��D�OL�Uՠ}C4[?��i���#ɃD�<�r���oU�2����Ķ<���?��UK�M��?�'W4�p��26T�'�P�\���@ڴ�?����D�74�� �O��'b�4j�$ �z0{����M�8Rr
ւh� 듍?���?Y ��<�H>��Os�����UUԁsl�̢���4��$�l�ڟ���͟��S������ ���Nt.L*��_4^ ��zºi���'���'LX��<1���5a�83d�Y~2| g��M�B�EQ`���'��'���e�>�(O�	3�`��w�ȡ����2~��P����њa�q���I`y��)�O�X��I ]G
��GfD/(��ZD����Iß��	��j��O
ʓ�?!�'����*ӕe�N�E+DU7ĩKڴ�?���?1�@L�<�OB�'�2O�!8�.����?57i�v/M�S�(7-�OB ��b}�Y� �	wy���5v+��H�G���7���oN;Q��I�5f���?���?����;B�r��ǩ�5@T��¢gw����+�x}V����ty�'���'���g��H;88�S��mN>X�Uٕ�y�S����ş��INy�/QY���(H��R���o&ؙpBi�3(�^7M�<9����d�Ot���O�AAS0O�-*i�	w�j�1��L�Hz`ަ���ß���ǟ��'�m��Ȩ~�<'4�CH��4e�"J�5?���@�i:Q����Ɵ���"@�<��ޟ`�wy��0�- �L�b,
�k��)m�䟐��IyB�[4�u��^��Oh�i،Ҭ�CAb�(��2���F��'�R�'	2؍�y2�'�R�'��I�>�Fx��&d$hY�����LQ��W�h!��ڜ�M����?���Z�_��}��G�#��e�Ţ�ш`Z��k�����O�ĉ�0O��O^�>I*�
ڇ|
|�٤dB�);�}��o�z���U劣�	̟0�I�?U�Ov�J�"p��\�ux'�Z4��X�i�d�P�O|���O�b�[�d�kg膙9m:�J �ʘ7%L6-�O���O�	��[I}bX����s?A��Y(0�TX��]7+��#$Ǧ%'��Pjc���?a��?q��'I�APE�S�u"���`�0!���'z$�b6!�>I+O6��<A���U��sd�qe�Zc�4�ҭ�y}2Ϋ�y"�'�r�'2�'c剫H�p���m�H �{�
�1Ra�-נ����<����Oj�d�O�}�$��3!�fs��_O���b��%����O���O8�$�Onʓ ��\ �7�x��a��)f
r-ô��'Z4�(��i>�I����'?��'��k��yr�N�q?�͠p#��,P�+E�r�7��O����O��$�<��
y��Ɵ��*l����
�B)�z�B��#��7��O���?9��?�E��<aI��Qf,�_�X���F�����#{�����O��\O�,s!\?��	럠���`��!��ԜU���Y��tp����O��D�O���ƅ[��	\y�ҟ�P��=.�)r	�*���źi��	�/�fK�4A���ޟ����dD ��1�d���`�<.���'�bZ��y��|r��K�nq��LўXv�t�P�	y|�F�ۿN_�7��O6���O���s����4�0Mˈk�i����,e�Ty�����M{���<�M>����'f|+ �#N�<HŊ�f&�X�f�o�T���OP��/O���%����ӟ��j1�CF����\�S�Ï&0@o�Y��E���)z���?��0�D����ުXCҌ��B�;A�֌$�i9�kQq�Pb�`��~�i�y�1M�Vth7?��-rR��>ɷa=���?���?I-Ov)�Ŏ8.�`iS�ʉK����S� u^�'���	�|&���I�,ir�*�Y�t,���[�l�&s͊���Dy��'���'�I�1���)�O��� J7%:uK0�BRp��O<���䓰?��P;@���'��9���P+�qiw�?�D,9�O��D�O��D�<��f0Z�OO�tR�	��5�B����n#��r��m����0��O����:��O�yq��<[�z�I��4Ui[��i��'(剁8��KH|Z���ƪo&�`�#�P�ƕ@�Q�g�'�"�'�t���'�'����/���sJ����E$
��R��U�X�
ڎ�M�Q?����?�O���\�b|�5�f�OF� �5�i�B�'��X�'��'�q�N�;1ĎB��%�c섕Z�v�ְiq��с�tӔ���O��$蟠��>1~	hU2���0��<�5io��lF�i��O��?a�ɩ�fu���K)k6*��$ s��$�۴�?!���?��X�X{�O�����HGB�"o}h5� '�
C�Q�l�J�O
hV�Y�ݟ��Ix� ��!�.#��{S�|�P�� �i��&�|��O���O�OkP7������?�P1��g�	Z�$�IIy��'1�'$�H1j�j���FP�	���^�^9���Ї���'V�|��'Wr��$I��� �ǹ�JҴ��#���'��	����I���'�>YK1�`>W�EWn�!��W�a����ɴ����O`��<���Ob����}O����"S�
�r�x�b�D��k�@�'#��'BV����%ϻ�ħ@(�D�P��0]��!F�M�V��it��|2�'u�n*(�b�>id�I�6m`���>�x�w����	��ܔ'`�Q;�a-�	�O�����8Y`�ؼ�\���M�8:f&������1n�ß'���'	��K'$D�p�\�T$�P��m�uy"�3"�6M	\�T�'j�T�.?A�\�E�R!k]�I
�0#�Vͦ��I��\8��c��&���}�'P�w�)0�+�u�D�Rf�Ȧ� ��ݜ�M����?���ڤ�x�O�:�W��%S_����LS�-��Y��a�>������O 2���V��%ځ��� ��M;�%(�6��O����O�����S}�T�D��p?���Q�H��9c���i��b#O���5&�x���q��?I���?yT�e��`�LH� *<`��	�!.뛶�'�T��+�>�*O
�D�<����phQl
��YN��I������v}2.�	�y��'/"�'�B�'l�Ɏc�t�3��oX
d+ ��#<�Ԅ!vk���$�<�����O�$�O�)ۖ��-�~d �W�L�Q� �s1Opʓ�?���?�)O�P@�L�|2�eC,)��KbH�1X�)"#�@ЦM�'s�_�H�	���	�ob�ɅX��Z���q"l��'�E(T����ڴ�?����?q���d��$��O�k�Bv�1ED�92 �����=ϔ6��O�ʓ�?q��?�D��<.��<
���u��5"�d���g��Ҧa�I����'�T��d�~���?��'?L��6.=���2��@����uS����韠��%p�Iޟ��'���ZY0�O��!�|�vA>0�6[�D��� �M���?	����wW���:f�jQ���S2|O����8*6��Op��D]=���Ol���O\�IEΎ�3Фr�	��*�"Qٴt?��qB�i���'���O�����K*fL����)n�b��gM�����gg��O����O��`��J]�d�e�1*wdL�5�>Y�t7M�O����O��86+Fn}U���H?��
��MjF�ȑ���Ct����l�����IHy��'�yJ?aч��S~�ș!Tf�dI�d�D���L,�y�i��u��|����1O����P��p=�(z��aCD���owʉb���:��;���$jY��3��#L�"I�W����W[4Y|�h"����.�RU���2FX�r���z��G�7Est��'��i�@a��P�S��uDF�vG����E $��pD�=Q[L��g%�?35�q��0`�<��L,u�R�T�K�L�����<b�'��#��'9�6��TG��"f2�˂eͭ<
@�,�r(��`W>���g˞17�܀E~B-3�.i �&�k�N�A�A���*EfG�h��P�G�!	$<��w�'cp����?(O�x�Á[�!�d�y�Aϟ��9�/|O�q���[Ĝ�q��ѣE~�u��O.�oڝ~i�q�t�QfD�[��x���IQy��9�ꓰ?�+�>�yb��OL-s�Js��k�@^A�`e����Oh�d+!~69`��ۯzr��z�O�Sl�dj�f��Ȩ�nJ�)0�	������� ='�8b�k`��3��IQ9M�^$µ�\3����ꜭ�e;2��I���F���'��ǧ%J�:��M��M1N���'u@`�!�C��ґK#��J	���
Ó㑞�9�lP6:*�Ҧ�I�g;VH)�蚘��$�O��D�"Q�X�1(�Ol���Od�4�2$�ɯ:�|���kt�*�΋kZxˀ�ޟ\8�a��E�0b>�OЌ�'#�{/t���Cy,�Ҡ�@!lzxe�dd�Ο�I���4:Zq��'Q�(`$���Ʉ/��1�6�' �I�<^n�4�b�=) "Y%���Q���|4�\iq�<)rkJ�1��,G�|��!z@�&q���'���NnЂ��T�D&
\���(�*��Ԁ5�l���O���O�ɯ��?9���ď�!�,1����L�D!R4k��Z���SA�H�,����Y8r��yB�!s<�h��i����D���N�[��!�^��τ1x��y�aރf�f���ڻ^8����Q�O�J4k���?a���1�	'�d5z �̾)�<�k�a��L�vC�I�q���kwBL>,@�
v�
&-hXc� �Oʓy�ұ�[���	/D`�ROR�Rvh��#�/;�Bu�	d���ڟ��I�|j��<.�(� @�3��䃑_s�a%�ܥ����N����xc�9F��h�bӨ](��ɜg~fHt�ׄ,�r�P$��e���%_4��'��	�bI�	x��W�d�R�ƀ�-%xb�܆m�.1VZ;B���I۪�4B�I�M����8Xk� �ե�U>�Ʈ�<I���+wH8�@���� -S�L�B�)� ���T��sOt�pf�\g��r"O^�A�ē1?fX@VE�rP�u�"OHDZCM�7&#N�@�I?�&�)!"Of��A�M$alހ�bm�>{°u�D"OzH�C��}8�5#�"Wָ%9�"O�A�e�<�ؠw�]�.K�"Ob<�`).2ة`1�,,(��s"O�lJ��T�O��"��[y ���"OfD�@��k��"S&���N�S4"O.h��垼4Mz���
�#�^�V"O�M��O(t�5*Y��J�)@"O�%{Q�=�}���ȇ�T"O(0���+A�ذbݔ:%�!��'�XM�4 W�l��	0Ý�-|!�D� ��� Q�;�t`{�B
�!�䘶�ʍ8��F=R"(A���!�d׃*̐���%k��C�	S8P-!�$V�F�%�pG[�!���`�͋_!�� ��ڗ�+E�L��V(�!��Ӛ��d����6��2 M«4	!�$��J� �'�ѦU�v���ɨP"!�$\'z��t)��L�֬M�#ǌ�!�T$)�dl�s��h'ЈZ蜶�!�$�;�� �")^m|h���00!�d-^eX��c���w����G&!�d�&2���r��T�v�#P!�䄽"Tjp�Q`RX��e��fH��!��;i�h+�.T	{�Jy��$� O)!���~PCb� A�
���!4(!�d!&���#̇7�VIVc3]!�D��.	Ȃ �.,�P}���É�!��4�t����J�"�+�!C/�!����d���� @��s��l��J&$}!�dۀD����� �)�����W�!��:N�NUA��D&	�������!�Č���cr�Χ%�(l��fʾ�!��*8���,Tв���q��'>e��ϯr�lL�&h	�UYn1��'.:�Q�N/vN����0QԾp��'a�(��A>4������Q���'vȉ��	Wz�����UN�a�'���1����(��o[���x[�'��p��s�t�Jc�w�vM��'�jU����v�ntW>s�����'kp��(�\zv�
b��p�R�'� �Q��6�Q�D#��!��}#�''.m��BA?v�r�#dʖ,�)
�'~V�2X��R��<&�J���N�<��% g�yy�-��\�����EM�<�R�"Ba:�0���dШi��p�<q��7k��y��,Jw�p�3�s�<�f�H��� {�B%�` �%�p�<�Ck�r���StOҽ +:x�Ҭ�n≄;�Vu��I	?
��3�\�k~ȐK��T )i��Uɦ�kT�ׯBsT�p���f��G��]D�(�4O5$��E�`��gj\�Ww&|� �0ʓN��Aʉ4_q`���� &��w�=������O��yR�vЦP�i�_J�94�ް�<�ce�`�a�D��~���'C��� 	����G�/zt �'<v��HL9J�n����BxPj�O�P�q�U�:�U _ 
�axB�̱V2���L�WZ�AN
�p>9pO&y���2w�E=r�Zx�A�[7d�^) �%��R���!��5�dR�2lߎ���GC�r!3� ғP�2�@	�/G�l�~Bх�M�H(�$�$\$J��@*�~�<� ��d]�7�t�ъYA������'��x�CG�Q-ɧ���T����:�����MN��2���� D�P9�Ep9"���W�^]i`�:?�%Nj/��$�k��M�"�/d`$�DX�+�a~"��5�\!���
�Hb�j_�;\���@�y�/�>�.�+
Х8"����̅&ֈO�ġ�o�%9�B �O�p���O
6M(�K�����a@�>��)�'����A�.�Ł� �'j(��'���e�@<h�by��9��E��L�S����Lݚ��uRW��3�yboICw�W��+&	����"/B�Y���$�,��Vi��ZZ(P�*4Fx��~�)�rc�,g�I��ϧ�0?	��C7����2M�1'�p}����dpc��oSDq&� �|�����c��O�L����M�
���4\~�a��_�\̪���];�^w_�ܒ$'�>g6�@b'�"s�@Ā�'�����}HD�4��19O��!�'�.=�T�U����L�82�	�
uXd�}���D�y�����<�Zl�@�	u8�x+1�'�~���{���ё�Yz#��Ã����8��#
=�?�3*|���͟0)�{b�\���B狔�7�4�@����(O�	*��]@�>x42F&�'&D�����Ji�*̷Hi�xfJ��o]�e�T�6-���D�(v�4��nӔM^a��#Yd9��gL1�'�d�fo](k6L����nQ~i3�'v����/<�r�X�@k��Q"O�L�tV�GM�|��aC�!�1���'�`t{��ݷy�6E6H+��M����.�a�c�0=����NB��iQs(D� k������i7 Q�>�| �U&�/���'	�����r!�����=I�R �$�JLJ:s��,����Ax�,���ޡ$� �%˜�px��2e�w��kG�2�xi�h�f�{C�<\O�ZAe�dH>tC"-M'q�vԨW�I�+VQ��	�O]���b��U7O�t��B8����N)*�z%�e�)D��i1B9.�<@¨8�(�SjfӦ@*��вG���O�0E�J̺��O�kl��� ���v%R3s"	�9:!���16� �I�(�'1�BX�_O<>aG�|?a�Кx�yୟR5�A<�ɠ�>5�f�B�%�,���oI)r�J���ϲd����̇W�P�� ̓<��i 3��:4.�xQE�MP<��GE�&r�����I>0)�V�ݒ5������ "U�Q� P��Y?~�0(�R�Ͳu ���ņ�>! ��@�P�3r��7=�,IǤH��y��[19�⒫�=G]4hʦ�´nۺ���@ n9��q�M��,�*M�*Oq��.�2�tA�c ��S�k@.`!�d��v��������8m5�R�2v��jU��cЈ[RH���'1�<h#">�Ɍ7�|����!zU�Ii�镣Mv���$��F^8�`�Ȭ��mp����ȹiK��Z���"�"d	��茝��,���p=I���GN�����75��B$}�H�E��f�-x0��ـ;^ԥ!�O�ě���>[rU�u+�,l\�u 8D�h1A��v��E�ACKNg1��6�thi�L&X��e�p� 3��)���+5��<nW:��Bs��M��M�e�<	Ǥǳa�M[�B�2dE�a��O�0�z=r��ԟ�
�:��5�OK^��=�Cj�x����]l��ȣm�U����2��>ؘ��c[ ��PB��
l�21l��h��$��.e��p��'R�L� �1�"��3��5
�P�'�jqP�:O>�HU�P/5��M褡'u&"��7�xR�A�m1�1���V�R���=P1!��U?�֩R`E����L�G���M�\���c�
E�=��$<�'V<�蟈Iڠ1�]�ä�A�2�c�=b������'�����5x�`YR�BW�V���{2K�-C��:�x�l��&)�q" *\�(ׂA���'y�QJg"J j�`�V�99<!r����X/��p)�0L���ܼ\����4��Aʇ\�qo�m�V#3�$H��<���N�V8� �솵r/�\C�$E",vN��G	 {�yhq�4��%�d�q?	r�J�W���@�*6�y�<�pXR�E&:[V�ʷ�N�z��7"O`��p�ӇB����.�J2�L����;5k>V��T��b��?9��S�3F�a�Yy��IS�3)�dIrjK4
��T�pa��w�8A��o�,]����.P*��)^r1�R��R��S�M+0!�p��!ӊ܀U"H��k.�4N�<�a��IQ�hl����K�A;F(܄qM��!bڈF/r�9Bo�FXm[Dj��L��M�?ݩ1�C�w���[�'�k&HpАB6D�((��ߍhL��9 ��N�|9j抲R\~܋���c�`���� .(*���m�'P���؜T���T *�Va���u�!�d�|(ma����.�P(�sa2]F�l���4Y�):E���B��pݽ�Ge|��O� ,�PCI]��$��r.T8���!�'g ��(RQ��SEeDW��]k��Z�0%���Ƶs�`ʕ����T�'��}�f%<($��Lµ<�.�ʊ��%3��l���R4�QJԯ)�	�DY��	�A7XXp�1&,j!�$5k�ܤX� Ώ7�ZݨPdU1m�B�U��b�zW�ŭJ��)�'R3�@p�/����J��	��<��'],����1�(T����]�ݳ�'��0�a�֧"ꙙ�L�U�E �'�D89$�<h�9:����\D|�z�'�^`X�!��U܍0!%��Ws��y�'j�䡒�KԘ�"�-��M{t��'��A�W���JT��q��O�N�*5�	�'D8�0���=B�zN�W���'U޸��k�+=S�!�r�(4��Q�'�	�KRo�"����i�ܥ#�'.��A��YI�qCbgC[��Ćʓ;[�E��FU&;��( �@�/M���ȓ>n�����<p���@׭t��u��N���	���
R��&g\���>��MX�Λj��j�b�<���ȓ$�z�a���N���%)ʺ���[U�\hr)��'� 4�DC#B�m���̓��B#h"���p�4@-I�ȓ]�9��W	�V��M$-��Y�ȓ�Lܩ�D��6e굙�d�� �\��ȓ&XArvˎ�g�N��PN�:Rn4��R�iBV�\��p!
Z�3�(\�ȓ[��xV%(�^��@��i��ȓ �28�CS+8V`1�VH��pX��r��Œ�B�42	t
Z&&��m�ȓ���Y������@qHI�ȓFR�BA޵N �YVK�De4��ȓt���3���>B�����2^r̆ȓ$�!H$�Щ38����ԥzz�݄�",���$�6O(��_	u���ȓ;����1mI�7�N��#ņ^r��ȓOy��j"cct�뀃<Ų��ȓ1�rIH�¥0�9���\��ȓm	>k����@��� �Q>E0��I���!��7hX���ʬ��)������8E�����(&����3a��AE[��TY@�N�:�,9�ȓl�� �T��i�J]�e͛�w�Dd�ȓa-�4�e�R质�uCĆ,���YZ�Dµy�H���2]h܅ȓ$��[�㖓KU2$���Y�*��U(���Y�15F̲`+9/����Y�n���,=˸1�'k�@����ȓl�d�
+%4���Òg�<���((�X�%u6�{��"Y �ȓa\�a��v�$�J$�q�N��ȓp�03*h���
�G�T"���	�ع�,H
!Bt�2#M��<y��ȓXM�k�
��E�.���ٻ6w�D��@yNܪ �:�] �"�1�6]��<ՂmcD%VVh5eG+7���ȓDi�e"f,T�;������+R<���S-��bKDi�P$�-�I�ȓ�Vl�2�Eh*����^� �"�������Xo�����*A���ȓT0#rɈ	th0�����~�� �T�(f�Őn_̐��M�Ub���+25b#O��)���l����P��3}��5l�>,j0{��A���S�? lM(��N2x��e*p���h?�0��"O2����>2�D�A��3h����"O�H��M�@��C[3k��"S"O��J𪍤N��[�k�����"O@5j���9a|�(�d�O=.w�I�p"O0���*�HԘ:�ǭy�����"O�\׮]���ړ��z���"Oz���1Fb�X�U����mS�"O �1E��9J`9��,W$���� "O� ��	5�l�S�X�ۢ`�&"O�\�c֌
���F+�W��4Re"Oy�&�����s�H��DU3�"O�C�
�=XU�����F���D��"OH�����!H��W�Lj�y�"O��
��<�^�h6d\FE�m!�"O^�� �8
�`���-טܚ"O�g��=+� X��(ձ-Yb�j�"OF\ b�?>|Z�h��\�"O<�@��ķAT�c��Y�*�"d"O��$+g*�ݩ4i�j�\Q3�"O.t{�+	��n�sR�BZ�0a�"O���F��9�ҕ���@ v̑(G"O@eȷ�Ԛl�a��ŗ�v]|��"OZ�����#J�e0��ݟYodtC�"O�����*S�)#��;JY2�"O�����[��caT}*|2�"O��PsH�uZli7!Ȩ(v��"Ox���4<{zM�W�Ѐy�t�b�"O�5i`ri�@ _>	��"O䵋��_�K�$p�Ã9�>d�"O����L�n�k��O�F���zA"O�Q��Яw�Z�"�xlpu�C"OD�PE�_V�A�OͿiZ*���"O��K�!�:UB��sCP�(�"O:	���L���W�Q�z��+�"O<I�G��}hR����Tr�M��"O��Ðh�F��@]�8
l�!"O���d�<kwN�Q%ٺe�@T��"O����P�)��p�Ođx�x�"O�d[�[0Bf����2\�!"O��j�i��)�\R��X+X��XQ�"O
��r��u^@��#N$r��u�"O���-$Z5Z9+7쎚2�P�a"O��bF���v��`��}�� ��"Ox�GEߔ^��%�v�'\��"O�k��8dbefѮ7��P"O4+Ԋ%q���s�LE��U"O����.T��������F�!� ���gcǦX�R��AK"9�!�Ղ9c~���	�pt&�A���!�Ā7r
.0����@���wb\�!�D8iz1Y�#� >vV���.���!�d
��\p��7.�ᔎ\t!�>4N��Gl��v�B%�p��l�!��T�ĸ� �2V�$AH$�Ϟ<�!�F�H���ReOC������J>XQ!��cn��Tk��BthQh>!�d:4m�ݪ0��;J�\�Źs!�w�``$�-;�qr�틦l�!�]���@2���x(�bҮ�!��Զ���Sb�*M3҃�
�!�^7
���4錎 �,LA��L!�dG�w��xU�/UU�����qD!�$Vx�P��fBG�	���..!�� b��F+Ѡ@���%e����P"O.���T/� U�$R0��E�2"O��	&��>AP��u��;4͘�`"O�L��E��igԩ��fF�"��U�"O��#E'����(����ՓC"O0��6.M��)�$nC�{d�YBa"OH"��G���[�M�?B'���"OaySc�'I�T�{�G&
�̙C"O2�k���
}.v0�c��h �mz�"O`�Z'ɉS.\[��ڃu��A�"O��q�`����*�`�Y� ��"O~Aru��N;$��Da��`��Yjv"O�BD� ~ ��p�`[�"YS�"O@���U[�aB3�Βh�E8�"Oܙ�P��9�*<�ሯf| ,G"O�0�CbZ-T?`y�@C�| M[�"O`y�t�A=I��ro������"OH�Z���5�.��0�.Iy�"O.Q��,�fХ#�&-C9�1�"O�8)/�Z'��BQ&�
aQ��s�"O0�рK���$`:B�ÎdD�\["O��Ks�џ	H�(��#*�4��"O���)N���,rp���u�5aG�)4��I7�U�M�P(@�9]_�!(d�7D�|��Ǖ#LR�iB,ɛkq��(4D�0[� 
+ � ��;C!R��4D�8�bn߶�p��a�n�����2D���CF���0ը�*J
�IA�5D���q��	*=�ѥ�V�g��Y���'D��(��47�>�i3����=�B�%D�\
r������F�b͈�� 6��;�S�'	8�J�	��&Y���ӥL�m<n=�ȓ���`'k� �2��I�f�������ɔ��$xDaD��)%yD|��A�h���@`y�I��'I�wJ&���n1�Uzގ!r �E@�t𢩇ȓ�P�`1+Ȳ#���`�N��b��ȓp�����[9QM��C���h�\̆ȓ>���ʀ�.�����A�X����ȓw�T�#�JȉOH�*�2#n��=q�\��b�
�Q
�b��N�Eϰ-��4j��k�2d�
 �t`�'ƴ���Jw�a%R0H��Ǯ�T��e*�UD�2&d4	���w�]�ȓA
u�WK܍y�����)�$�ȓv�bh�c̗4�D���K"���w�8��p�%W!=p~���љl!� ��@ؤ@$a0��@�[\�ȓe2!�T��	qyx`#�)[5��ȓ<� (�1,�,T�i��ID�86u�ȓ}0s��Ӧc���ڰn��E��ȓ�Je�%I�]�tdh�Ŝ����ȓgNV�����R��T ��ט �"5�ȓ�`�i4h
_��MȐ����X��G���b�oLj��ց~� H�ȓ�6�Rg�9�8�4��2�2m��_4a#�	K�r�t��?>�V��ȓ_��8Hk�7%�,\eF8}d�M��Kw������lh6&7L��H�ȓh@l@�Y�wŲ�C��͍a^b��ȓy�� �咒�"���2�B���7��ݺQ*N�D_ju`%C7��݅�4���	��ɚ/D�� &�ۻs'����q}�pQ�Rh�|P�we� �Ԅ�S�? ��"�]>q�E�R�͗.�� Y�"OR�3�\��zb�>ZQR-ڳ"O����ߩ]̾|���;FԀ���"O�����E��qBN�?5�=�ѽi����#�B��0G��r<%(�D֭Jf!�Ą+>��!��(q������M�!��.Z*�)t�C�U|�d �7;�!�DE��8lXD�\������)�!�g��q��e:�A�GԈ"�!��ɒf�x([u��3Y��a�f�(Q�!�D
;���ˡ���ri�D36!�$�:Q
\X�(\��$�kr��z!�$���ÄƐ~�,; �!w!�d�}؈�҂�H)^���GAG�\�!�D�T(�������-0�b�-�!�DL�&`h�R�����\����'�!�䆇1�\�p���6��Hy��� G�!�D��}�lP���z�&q�S�"�!�d]�8�ѐDA9(ʢg'
5F!�D ?�L��5K�83�ąU!��^���	�G���RI�	S�T;!�d	H�jI���])pS4�!�++!�D�+c (!�W��!.Pi�-T/m!�j1�i�T.ȍ.��Kڈ1�B䉿�P�Y��
v�Z�[��X��(B䉮.겝��J�� "F�AT,�juJC�	4/��UU/�!v�N4��g��@&>C�� .txHz3-�3+* lcQ��,o=�C䉫G]^T��
  ��R�oҙ=�C�I�hx�JR�l���Q�	L�B䉅��Lh@��_K|@0�&�{-�B�	 A�����:&Fd�V
�]��B䉐�&HC�F� (}.���φ(8YzB�ɺ4sN�Ɇ
�h��a�,D�4 LB�I�4�������$�}z��D\C��$s�J� �	�~ձK���C�I�^��
�oێ.-\Y�����B�/{���i5��0�r8 ��@/+QC䉨@�$q�nWV��%�� "�BB�	1�R��̪o�j	��jZ&B�6s�l|z��	�lm���P$*J>B�I3������%�6�:�f�,�<B�	�;L����	P�Lg&�H�Z-e0B�	)�6E���]deVQ�0'X�M?�C�/W�ѸWi� 0�bͱ��ֱg�B䉩=����s�X,e�\�+��W��C�I�G�<����BW�E�E�ϧv[�C�ɝj�!�`�O�n�H��L�E��C�	."7\�Q2$U� ��0
�x�C�1�ڐ	dVi}��*P鈴Z�C�I�*�����0�T��Ì9_<�B�	JŬ�����!�1���rB�Ʌk�\Q����C'�9����2B䉉;�L��[�T2t��ni��C䉗L�Z�1�g��*�2��G+�# c�C�I<F7аhCdӸo 2�P��F,�C�I�fB�]˵�N5V�p#Da��1�B�ɷL�pp;��\�cҐ��A�&r�hB�8(�,	C3Gp���p�G8	�<B�	=v�9�N�7X`��CjK>&b|C�	�����E��HZF0����T�B�	�z4 �\>�����G�rB�	� ���r��8c�΁ F�PnB�ɏ�L*�	�7@���q �DvC�)� &�C�1.8���-��_s�i2v"O��P��%-���q���Խ�%"Od�fޏI�f���%�x��1%"O:\�`�T��č0�eO�L�LJs"O�e*��P-����$�,9����"O`-���X5<ĸ`��V�i��aS�"O�Ds��ނj��B���?�:C"O\4	P��L��Ǥ�5fޮ�@"OR�V$�*l�&(b�5d���2"OD�9f�Ծ>�����`�3����"O�����R��,s eC.YR�R""O���Ʃ).��m���ЎW�<:Q"OB<�Ƈ_�y�2�8$���FU>��"Ovh[�lK�\���U�洱J$"O�@2u��<����Q��N�4D�0"O�jP��&;�(9�Ǖ�0�*���"O�IB�?���Ѥ��}��M�"O��AO�-4���C=Z��"O��1oA�U|�˵aK1a� -"O2����%v��i��U ��}�"O�,EF�Yh}��cP�r�K�"O$p�Ō���-��b�2��'"O@�'閮k�&�ѳ+�蝃�"O�Y�5����𢚯x�>p��"O���$g�T�5�� e�"Oԅ3"& ��"�i��;��"O� I�-W���P�HG���"On ��o�h���5I��T��"O�i���9_7� Q�C�х��c�!�D[�Llꅂ� <�!���ތH�!�dĕu��L	��� B�HX`F��*�!��?�LT���P_:Z��1,�U�!��ک���@�dΰ�T��L�!�$1
����E���m�`�R?�!��ֳ#�ʍzs�U�Rj�a�kA�Y�!�$ѨD�d�"B������S��2�!���'�l8�3���_�M*�I[27'!��u:��3�Ήh�.�P�'A�~!��6r%j� ˆ��$��w��co!��K���A!+Y!�� Se�'_!�D
�$>�a�4�E�x���C�B!��,̬9�E2c�N��B�MZ!���7	5
�ز���̤qAV!�dH&�nL�+�0u��	�%Ʉq�!�䒃q�,���C�XD�� s���1�!��LYp���B9P8إ0�"&x!���	(����%aU44(��A����!�D	4jg�D����-����`IM�!��bD�'JJ�Ԭ�k�!�D�V����0l*C�����@V	
�!�E����c	Ҽ:�F�j'Ϝ9+�!�$��[;05;!ܸR�>�bU�ڇ�!�͵^��2�!˫-��j� �7�!��ϐ#���9eE	6X���(�!��Z�\��7m�<"gB�+��Q�d!�W�@�N��`F�X� ա3�YD�!��B'$��v��&[�� ��F��;Y!�dĔf}V�8��U�O���pf֙|K!�$Ȩ7#Z��o	�9��St�y5!�D�(}�%��\|�&IYg�<@�!�$`��eaW����u�a?8�!�D��2{��Պ��� �e��N�!��:EX�Bs�&"�0AAB,nk!��U�
��sQ�X?m�$Mku��+_c!�� � p��a-j`��JiXd��"O�ܡ���4Xdz� Q�<W���Q"O$����^v�%�$���+9�iA�"OH��1�G�q_�c�ᆽ80���"O,9S� �@dTi�/þ9�lA�7"OB=Yb��=E�x�b:qH@��"O���3C61�(��f�F�t-ܬ��"O��*�L�O����@29&��[�"O2TSuo�@��hFM;�@P"O�`�eƃm_B�F�a�H"�"O��xrM*���Z #U�h��Ä"O�Cf�@3��H�V"ɛX�j4j�"O>ܚ$[�T�!�LS��X3"O�xàE�N�y����o�ܱ�"O6@¥�h܅ʒN׍#F:�{"O�(:���'uh0�m�,[��s"OB�;U�M�^mc�L �pmr�sU"Of{�@�t4�ѡ����q��	��"O���`�+e� ���!}��*�"O"٣��y�d5�3��.I�A�"O�!����QڈHC��0�h��"O���s�R�S�⁠��5a��0"Oű5a�-b��pC���9Ϩ�+"O:��&�>&���#ghQ 8���
�"O�xRe��p�M:��J�D�m��"O<0 Ǣ�]?������"_��}qT"Ot��dZ
��b�IL�D����%"O2�s�!ЀP��dp��Y��"O����ż�����qw�\�"O(�e@�eR��B�]xs����"OȨ3P�-���(���9 s<=B "O�ܻR���qD  ٳ��Q�pm{�"O0��D�R2��Q��0]��	�"ȎR7�F���hD=J�Pˡ"O�AӶ*M{�� ��� �R"�"O^�UM#,��,�ф�U�Ը��"O�(�@5I�0��Y%E�� �s"O�����  {l,����}{� ��"O��YTR
p�*1s�	xk|�+�"O
(.�mI1��$�E`�c�/2!���t��#	M�1�dU D�Ϧ�!�d^�w2��p��:J�
d���b!�	6A��H��3VFN-j�@��4}!�DV� �l��1%Η-a$����-y!�'r��#$��T����6@!�D]0cV%A1S�j�*i��/�>)!��-]3zy�#�Q��e���͂sA!�ĕ%���jԏF6n��;S��B�!�D6��(�.[�GTH���:zq!�_�~f���*G�:��I�#Δue!��%^����#i�B2r�(w!D]!�ě>B���!�$"=fqC�(�!�dH��A�!��2*F��dG\�k�!�d�p�������6)�he{� �!��U�5Q'g�K�n�!c���Y!��(��L�P"ۼL�.��g�3%!���<h��{w���a�v��хČ6`!�D�3Z��]��T�j�^�K$�ק^!���4���/	i��{ 捥VG!�+���;�76|c��F�**!�DS}�~-[�FߧA0R���J/�!��a�$
� 3L�2���(]�!�$�/��j�O"p��xu�NQ!�_6	�L�G��Qc�ቖ!�� ѳ�L7G��+�'�$!2�"Od@�q�O�v��'��
�x4�"O6���
�)͜8�S �5XO8�t"O��kcXP�;��� Dp��t"O���NA.����dO9v�j���"Oh	�t)W� ��%�S�б5"OZ*b�]5��"�#Ы+��!p"O���W��TE��0Aɏf�nEʦ"Oj(!�O�`�XU�W��5:~0
�"O"�{b�7NIP�Yp�H�D|��S�"O�1Mı>�L��兇5w�PIE"O\H�uM6(��4"4���dy
Q1"ON|�+R,~�r���)ƒ�"Ob�S��6��u���ȩ%�i�3"O,y���Bw`��S�Jڗ��D��"O��0'%F�9 ��i��*�S�"O�X�S�@�����>K{F8Ig"Or��A� ߰�h���!_�"�"O�Y[0I)�$X�%�R��H
"O\(���|��C��]�bP��"OBi
�����M!3�]�����D"O��@�2�܌�ď��S����"O��K�n������s"O��e�C$KP �4,�o�h�8��'�1O-i���5<�:��PR�ĸk�"O(�9$LZ
uB�ɰ���8��]�"O(�����+�nك�H

�ha�"O�8RB�9��I)�hӠ(�̈��"O�SBȂ<uD��Fƌs�,t��"O>h�poG�j��ڡ�{��)i1"OT���
�4PgE�4�g�uG��!�䊡Q%��djS�4閹J0-�k�!�Z�]ԉ��-��
��U���IK�!�$W�H�X��"�	z����,Qi�!�DƠ1]�m�BH�-&�����
]�4�!�U�)}X��E��D���5�)	V!�ɓ+�P94J� ��9ń��yX!��; ĞH1�Ҝq1�T�b���!�Z�>ȩh!B�7+�r���թu>!�D^�%#���[�I��"b
�S�!�D!�H��g�T.n���ă�!�D^�u�ڡ�ϱkkJT$#�(�!� J���C�虧e���iPK\�z~!�J*��,a���2#�jT�vJ�+�!�Ï!���`�Q�~�2�Ro��a�!�*�t��㮁�u��e��K�7!�d�Kfx@(_�<��ui�$R!�J�{C��(��	�B�uraǕ�-!!��6,�\a�%Ҽ+�{���2z�!�ϭ�NɑA�	\o|yۀ���:���9O�U�����@�c%_f{�"O����iа�iͧf=��0�"O��x��Z+V|IT"�*����S"O���Z��tMj�a�6a�"O4����4X RiK ��P\)d"O������ ���ufօ`!"O\Eҥ�W2�\�"��.;RJe"O~�ak՝mX�aA�Ϸk4�H�"O��*F-��*��Rf���n�D�8�S�Ԭ�9R�N��AK��|�.%F�!��O3s�,A��+�
f2�cφ5-!�˜E4�Y)F��m=Vt����J@!�Ȭ-�`E*f'Mv!��╠M0.<���4� �!eca��ؒe5�p
��� PTa�nM��dz�(ڄ��E"O��� ي��ɪ�h>u˰���	S>��5ާ8*h�I��P���r�.D�X���%H�x� +��ThRY���*D����昉7o2�K�Eŋw�(D��(��Y9.�6�7����I#�;D� ʰ�Z�!�K�3%^D���7D��C�ǻ��<�F�W;x��lg'�<)
�--����gŕ�佂�`�j�ؙ��HA�!�I^���IU՞
w�ȓ?��$KA��<K�9��)O��v�ȓF���P*�f�h\hceN1沈��8G��8ug^� |�t�1e@1t펉���z0�dM�L���q�L�J����:�8�Ą=W���&b����R�� ��'�X�	"+� t^���9�=�n��F��Q�Ƅ�ȓI�^�,IC0�A�)ϴ�ȓc ��R�KW�4Xa-Wfzф�M�(��.��j��x�ԅ^�C�"���"����V�WZ)���D>u9䘄Ɠ
����%��$�(m@��?��}a�'$4H�[�]�1��WR_R��'V�p��B:=�P�w
����w�4D��0��� "���V�3����h0D�ę�E�9v���I+}����+D�Ļ%��"4 ���@�-]2щ�(D�$��$_:����m�0A{Eo)D��Z�V�^d`��hWq���&�$D�����k�x8s�9��P"L#D���#F�H!R���l�"��a+ǈ�O:B��'g6 ����6(}��ٶ�Ðc B��u����ÄI���9 �ď�$B��#C��tK�e׿b����z@<C�	�A8ƕs6�Q�Zb݊7��#��?a��	K� 
 ��iֽE�����
�Ij�yB�^4�|�t��"A��P�[�w7�B�ɜa���!��Y�L �>A�C䉼_�
)���ρ:Ĩ��K��>�B�	�%��+Ҩʤ]�l� q��KD�C�ɳn$��)Ql]�5�P�)�B*͈C���,u��g_���-��w�fC䉖C;���@1��A1�@bC
�=i��hOi�G�R��^(���ɲ0��	(D�<Ki�9-rt����,��-"D�T�H8.��5*���0C_�x�u.<D��i�Bю5Ɩ]*�a�1-x�c�/D�\���Ϸcb��oS1���j�,D����#�%����R�V����7 .D��r���YW�KdĐӖ��S��<!��Z�P��
5l� � 3�'�D|��"����f��w�r�!e,Ȥ.^̆�Ccع��n��Q&�М[J�'��e��*؟W���"M#f9��k,����R�F�Z{�nR�k�v���T�V�ID�O-'��l!5m��n@E��j>�ЄX)���c��['6��:3�*D�L"��a�v@9"�	�%�(D��#�׋Q0Q�&֬�N�kF�%D��x���2o�PRe��4�D���8D���ՌVQ7*�v�K`'� �:C�Ibj�DK��ԕ71j������'��C�I�?��dJ�
N��d�S��1	$�B�	�%WJ�:P�\�Gd$��L�^B�)� �i�G�*hJl�c!�R�%6v��4�'�D�)y�2���h
�5|Eap"ܸ	!�$�^�~�� �"�v�Հ�;#�!��tɴ4�e��l��T�v�!��(!�j����b8�r��@H!�$RCߜ�P��H*~��o)A!��,4��!�ȋ��h�����1J��}R���u��d��b�E6l�h4*/�O��HΊ1{bU'�TX�,��Q��x�ȓ1B��v�=I���s�c4H�@�ȓ&&�Hg���L��V�ϋ��̄ȓp`rPk�@��]�� B�I
 ����ȓU"�bvg�=t��В��u6<����~��b�C:蛖�J�&5��ϟx�<a�J��-/���6�D��k�k�G�	͟���I�'��Is�&�z\��U�܁X<��i�'nl!�f�S?H~>�PS��K{��'>U["��$f��*��+�&��'����6	�Z�HC�*!Rd�xj�'��i�&
ނ:��8�@��'^�����R5-�{�'B:H=�@i�'Z��`MS}0qh��R�Θ��'܀�[�lY4[o)΁�>��r�'y��Ϩtgk��
�9�&�c�'@~�K�쟐M!�pS�$�i ���'i 4�1�_�W-LL�TIX"/o�}X�'?R���D�9���S��(1$�R�'L��)S"�SQ HYЄM�jP�4@N>�����E�O �D���ѣ[��u��ԭ$!��+`\�_蹳C/��V��"Op��W� �>�p�p`΄�G�B���"O�e�P�.|x�ӫ�$���� "O
Li�-I�k0�=h��.U0xa�c"Oڤ���7Y��\� ��%��cp"O�����!�b�E̛;?���b���|>-�p�U�e�¥X��[�f�����%3D��YV,�oG��;t�������#1D��H�ѫ
P�� Uf]/>��0p�0D��I��B.������$f���ub/D��yt��s��H"!��`�r���&,D��YCC�i���cDF*o�:|s�%4��D+��ƅA���z�񃅋�L�<9 �R�8~��6�E"�m(���F�<�aB��;z0�Вi�k��)����W�<q"�( � %a�6�:�+�LBT�<��c��I����=H��d��VM�<�P�G9Ze���"h@��95$�p�<��H�~�T����!d굹��Wmy2�)ʧz�ذj"�a���W�3-ޝ��h�0�r'�/y�T1!�I���QOJ����� TY/�?y�e�ȓ��0�b.�\��-^�"��(��o}����/K�6�������*E�ȓ{Vb� ߠ<���vl߷
P����uJ(bc�P�r� �����4EG��ȓ>:��R"ei�v�g�J1b�I��g����\5a�E�#�F�xv��r�p��N#D�@�B,�I�$��-p���M-D�XJ���a�Z��b U�y��)7D�t+��	�'�=���u��] �&6D��G�+Hʐ��pJ҇T�R��/D������8�P!�UO�C{����'D�$��Z�"iZ�H�k�?I��a��(D�h$�4a�҅�D��C��:!3D�� $m�
��
P2D�`�S#
i��RE"Oz] B)R�BCEܐ f�c"OJ�c��qx�kO�;�'r4O�!1a�Ըmw�	��S,%A�d E�|��)��Y3�e�t�,.���&K�2�C�Z��y��NCSA��Z0���G�C�	�:��}�p��۲4��燿b��B�Ɍy]��0�\�c�Ji��ЮT�B�I!9�`h��i� tF��܆B�	?�r���	1$̛eo�7S�B�	�tV��r9�\0PcPY��O��d[0xi������
-��Ql�	$<!�����x �Ƃ5���@f�Z)!�P�l;����\-r������ͻG�!�䙪D��0�$2�ʈ�&�Q0i�!��I+���C�3�K�\��!��?OH<h���46��u�:-�!�#v�� QrNI�5+t���-�7�'	ў�>���	_�k.QZ�k�9L�u��#D���S�ӋB]����ăv)�i�D/"D��a�@��:����W�'펹wf D���ũ
(	"|h�3�~u*� D��s��G�b� Nߐa� �Z�j D�`ʴ�:Ҁv-��.��eI��>D���2�D5S��(R��>'�1s�d?D�02�*s~d�w��%�֥cա8D��Kt�M&�f`�#�#B�])�� D����S�S` �P�π(�d�#�1D��d:�J1�B�H	���1D�|�S��8����L)lr�r��<D���PC�s2 ����yE�@�9<O�"<9��,n� L9S�ۢ�H�Ad*�n�<�&�4��z���*"�6��FGhyRX�H�鉭E�L�9�;8�D�����)�\C�I�E�Z����O7Ś���$KFC�ɱ?�X��t�\�X��yC�J�C�ɲy� <��Ȁ
�P�@�d�)C�ɷp�0�!�7R#(�"O�c�:C�I9a���B2��+G����6H-t�"�D"�S�OUd�aQ�@�G�4�wo� J@��8��'��d�����#�,=�\Q�!� 5j!��0[�$ C�><����!k[�2!򤁱~T)i�oN:I.��z2cL�E!�dU�`F�) ��4#��S5��!�$W�m��d2���)W���נ@�z��y��'�'��I��
��A`ԎÖ~
���D>�Qϊ*{��5*�!��k٠Ii�D#ړ�0|�̥�Ě�ϑqu ���A�<��	j6$� �ɋ]I��Dx�<	B-AI�!�1E��#�ƘF�Or�<A#�#��q��.R:EZ�T*��Kq�<��OC
9Ǯ�5�J]�֝��kQp�<�u��eR0�C҂n6�X�o
H�<���İM ���N�!����tKDy��'��@a�ݥ����.fVu�
�'�0�Q�+���n�fFb�r	�'��K��n����8ތ�C�'��;�^1(*����6�F���'����қ 7�x��� #@h�4����y�'�R4�Q+]80y��Z#��9��=1�y2mX�A��P�
$X�APR�P��hOd����gބۡ��`\"�*�j�OP���.FX�I���yCӇ�=�!�Ez�`��䤅EB��F�B�!�� "t��]
:I���-G-E�d�1t"O�TeD�b>,��럴}��t��"O�́��> ���Soz�9���r�O�:�6m0D�X�A���S���	�'���d���.!ҝi�)�0v�88	�'�|�K�&2�ȳ��1mf���'}|ZECL{Ќ	��cá;�@Y�
�'��%����L�:�m��	7|�X
�'���XĤ�/�6�)B�ȝ����.��)�醨 ��1:�
 �xV�1O�Uz(�;Ȑ"�呎g	pl�%,�O��=E��n��.���I�n+��e O�O�!��?^t`(R𧁤�iy@��-�!�'+��-��Ț�U����4�!�D_=׮4k@n�)��s'��!�Dڡl�$830dڛ?撽sa��8{�!�DK���� ��X�ɍ�V��{2�$+^@I��N�A����VK�(��'�a|2	�� ��1�I �Y�Ț�"��y"�p<�#㏢I(�A�[��y�j��nٸ拙�@ZDP{1�
��yr�ےCd���%̃kA��Х��y�M�a�rW�_�F��F���<��ڶt0��+Ԇ�z��h"��N>0@�}�����'�N2@�X���N?-:4�A(1�O��m�����/�#H��{��?*}%�$��I�"����P�1Nd�C�ʜ:�B�	,�
b�,ψ-"f�b�&�<,�B�	��.�"_�foV�D�X��B�ɎA�(Q���[;�Ms��{��C�	�����GO�gspm�ciJ�����0?)�$�/Epᓅ��("���F�i�<����56�{���6>Zᨢ�Wa�<Q���{�.�3���N�����P_�<qs>.�C�����B��C�	5e�4űR�E8jq<@�TB�B�	�
2BU1@$xxт�_�B�I2 ��mSpG�~��ib�:`�LB�I�d/&��Ɗ#Z@�Dc�%7.LB�	�8�� hpJ�2Eb�b���?;\B�ɿ_��gŔ9DX�2%3�"B�:*-������-M�������V<�C�	$&�:����-w�r�A3���C��W����&�b�X@��R��C�INCZ� ���4,���B�2B�ɶH����+܆ت7_�[�2C�	�Z��m��A�u/��$CP9Aq���4�����
�~7��r��:l+�x�f%D��{��F�\0�%�],$����$D� �wL��an��X3�W/2��YQ.>D��h`j޶{���s����/�<@BQ�?D���bi�"��S��9`�D����ID����?Puz��?*;�j1�G�Cg��D7�S�O�|�Kc(׶a�ơc��D
9���§"O���G��@�J�M�b�c�"O�P2�N�O6�+ˏ�e��D��"O��Є�;f`h)����)D��,#�"O��C���	� (1{{�]�2"O����* 4�Y'@��#p�Ġu"O�("ŉʙvr��ea��U
\�"O�٪�#S1��QQvJ�l�M�"O*��%,	D��}P�	Y-:iNM��"O�- MU�U��H1���=��<��"On�����>�`R��C޴�@@"O� ���`2�8[���.���'"O��J�.@*����&�XI�|��'�R��~��Ͳ_���rRd	S���Zf$�Y�<�S�pi� �����zǒ�
�^�<�&�A�S���P���;��i���<���1�sb��8�.�)CLL~�<!�f��`dh��X'7��Ac	�z�<pE� yA�f�M'U�eQ�Cy�'��s�'�f��nު��T�f#_�=����	b�'?L�Bۜ!W�̨h�)��K�'_�Г�	�/�nm����wo� ��'���Ev���@�׭nXN��'�^���GL�l��X�&iG�{gD<

�'��X�!H���x��>kvU�	�'_��PC֢�t�yר�^�\0 �'NzI�U�SE{������c���j2"O�|��!���� �lܔ?v�p�2T���':az�EǠ
6>Dە��,j5ҰM���y��A̎< �c�O`%r���?����2�f `��O�p���v���
b<����L��`+���؆`����q�1��F�Q�v�����	�*���q�~`�2%�_����Z�F��ȓ�9y�b�4fa��Y��ȗ �4���M�����n�)S�sK�a�J�xT�e��S� A�K9v��4�j��7��7�j1pe��r:>)��?��ӃNܞCb�ɫ�����y�ȓ�5FC��m�X<S1��$"=��s�h�������T����J���ǆ ���ĥ�n(Z�n+�P�ȓXj.�ð��V����m��@h��I�n����~ڸ�Qf��2b��܇ȓX�����lMb�;�Ѣb8!�ȓ8܄ѐ�݀Q���"B9D@�ȓn�ځ��c�_������BMlM���HӅ�Y,y"�A�gP���ȓ	���B �_-�0��ueBĚŅ�w ��([,4��X�����ȓkDb�9�o��{L�(�J�h
0��0�dB�d)N���ʴHQ�ԅ�"�\X��oN�Aqaĸx�ڙ�ȓ��W*A]��v(��V�ȓH�:A�p�4]�����b��&�4��K�`h�u+Ez�d@x���h8ɕ''ў�|�0��!q2����-��Q�d�<��H��	0������(!N�H�� ^\�<Ѧ�5,^��҆��gh�Á��V�<i���c���3u�GWAb�rg��Q�<��l���DZŎD=D�^YZ��I�<�W�}nH�Ƈܽli.��7�C�<9��EN�d3�k�6]���� g�<��^�2y�-
%k��=�đk���Y�<���,�<��M2a��B�d}�<I�E�8h$�E1ui�P�w��C�<����v�("���'��`���|�<����S���ƬȤl~��QE�Q�<YC�8�<Xs��V	=���.�y�<��&;m��+�0gZ��8Cb�t�<���ƛg�V���ɴY�X����L�<9ª�+���sR0 ��w�A�<i��M�h�����($0�0(�%�T�<��Mڋu�:$nșCa��J��yb�'c��XX�f�,5���
����y
� �p�dE�xmA2��I�~�́�"O���/8~�V�c�D�=���i�"O��
�`D�'|f8y��*�\!:�"OJu�ɭZ;5���D3;��V"O�H���R:z�<�P��F8��"O���! ��!�k�Dף�zhi�"Of�Cr��x�[�i��0q�@:�"OdA�pgQ0���ꇿ�$��"O����fJQ�eI��+Y��#�"O���E@F6M�<,��+s��M�"O|��� ��L��&�2�P0+`"O�t+VKW(%k�8i�c�P��X�"O`��e`���LS�e�� p"OȀ[U☛BM�q�*A	
&@��2"O�pP0�^�?[މX���i�i�@"O���Ó�X��鱡�P�5I�p�"Of�"�ό-�B�pW�?u/� !p"O`$#&��+0��5���%-��Hs"OTš$�0CA�F\ ��B�@z!��_�l^�-�p�
R�ϏkۄP#q"Ob��#�
�p���ά8�J�ɷ"O�����j�xD��A��li�"OV�x%�Z�)�S�ϝ7�I�E"O�#TE��Q!x�󷄛1Y̎�p#"O<��¡ 8���B�5\� (��"O��)�&�H�4c�-Ҡʵ"O�<��+
(乛���t�X���"O~Zr�<=�:�i��Y-4}�Px�"O�tzÀx���3�e��'ydI��"O8
�n�'/�I0E�3mq�!Д"O��tHC�!����D�UKR���"OT�řQT`)����R+��B"O(��0"	�\�0���F4��iQ3"O��n�)E��"a싼����"O�z %j��5�V�Rx�X�9�"OfYj�k�6�z���;ll@�B�"O� p��`i6�� /��T��"Ov|���ιk~2�C�n�60���U"Oɨe$�+t>N�ĪA�,<Q�"O�Mi�@`��Hs狺v�P %"OZE�@��3ج����bk�]�q"O���'`��m��¤f�3h��ɶ"O�p
A�����e�y���"O��J� �i���6�Gwf ˢ"O4�	�Ó9����$��"b�`��"O ʷ�Ӆ\I:}ca[b�8` "O�81�I$p]qW��>� ��1"O�52�G�=Hf1��Pw���"O�	�b��0�V���Ά�&��H�E"O>��H� Z`dj@/(�N�:F"O g	�G'�4��ɛ/�TE��"OD���cLݚyS&@�Z� b"O����e�y!�yReC0A͂8a"O���4�S�cC,` �ĝ;��1;v"O��w 
�`��Q�E�F��A"O�0�&#I�c@DT!G�%]ʀ�4"O�]X���L���/E�\��|��"O�	�Î�1"��H��ϠAb�8Q��g�l��KH�*�&��'�Zq|Cl2D�t3��Z/��a2mX�Axb��"D� 1,	�1��Y�4��4�����A=D�������q�F��OU����:D�d˃�z�X���ǖDW�m*�8D�Ԋq�ޝX���P��Ц,Op-�M1D�� ��3��K|9Љ�S��q�Q�|��)��+hJ�`#��A�1p4*U!�C�	�9٤�Avb�k��p�b�#75rC�Ƀq� �BD�[�R"���wo�4�C�Ʉl�>Hj5�ŀt
l����Q�6��C�ɕ_R��K��.oZ9#hA��B��0�`�QA@�>U�c�Ϋ_8�B��f��-��C .D#�p���!{�RB�I�e-2ݨ�h]�hi��a�	�*�>B�	�I�ص@�ɌsY��AR�D�Y?�B��.'x�灟AEp�5�߉!ߺB��b`dKb�RT�I{�	ܿO�tC�	�d�p��q��(M�n�� ��I�HC䉫0���c��ӝ^�Х�=J�$C�I)~+:����qk� )�̀��̣=��'
H���6eÑQTr�xg�:\&"��z���iPIM�Q���&9`a�5��p�.�I�`V7,�����׌IBܝ�ȓ{2DI顭�v�\�rM|�H�ȓ^��)��h��V5 H9ff�??輅ȓ�ZQ�.�#y+рI=&I�Մȓ��e����z�����D�Y'R�D{��O�()�vI�8-b<�����F5؄H	�'z`L�����A�����?��1��'�R)��L>$�T9(�hUfT^��'�8["�80�����hI���'}�yR���J4.�)�! �cĶI��'��X[AHāG�)R!ʋ�Z=&��'�nxQ�-.Y�܈;`kF*�c�'2R�؅+�3���j�%� $~&!��'��3���2&�.ԁA�o�8Q	�':�[QBW��l)�����|�%��'.B����j}�$�#��:|��<�'������M$�,�4mUs{�3
�'��L�&8N�|p��"���	�'�d|Ӑ�ҺQ�4(u���rea�'�q	4�\/2�&m�t�`^���'`�#�L���.�kG�`cz�
�'R�%csϒ��Q@�n�TiH���'��`30%Kv�CuA6L���'�2�7
9b�W�Y���a��'DH�R��V6O4��f���v���'���wFB"%L2}@`+xL\�A�'�l PU���$Y��Ҽnxx4X
�'�~�٠CДK�@{�F:9G�\�	�'�ӗ��	˶UC�g� �DL�	�'�D���]#:�x���z��	�'��L�f[
do�\�ǋ���"O��ԩ�ۈ����µ�"O0�"��$d�NY����~VT��"O���WG�5�h ��F�}+@��"O�]���	���G��"q��0V"O�P�H�Cc�\rsJ��y�"O ��!�x��Bc	#5�%ӂ"O�(�CTOg$�D,_]	��R�"O��F���$5�s�����5{�"O���`)�.��0��J�t�4���[���'�azR�גD!8@��.�8>LH�b�yB��5�Ȭ���x��;��,�y�N���D�@9�N��Q��y�V�9�^�"���)�p�K��yR��.0��8R��������]��y�o̪tk�܉��In,u���y�L��}�4�y�h�$
w.�h�+^��y
� 0a�H�L�;�Ϟ7��#�"O,�Z��B��4�
�)�?���&"ON�5��u�ed�*0��IF"O�r7�3?��m�E�%{|�.�yҮ۵>�u3N�&R�����y"��X �D*ĥ��X}86���y��اI �Pŭ���4P��y���3#���I�[�&���J�0�y�̆�+�pl"ǆ�O��1�aԘ�y�Ȝ(�0cʑP���D��-�y"
v��24�"7�Rm��ˉ4�y������
&`M�B�D<�-�9�y�j�> V�H�C�4s��3�t�<A��7N!�|;� ͛M�^IAF�s�<����v�$�@��0� @!q�m�<�'���@)~�c`и B�и�$�i�<	v@1T �̳e+��~&)B��Zf�<ٲ#P�T��3
�2�@�G�<` �/��xh1�J. �N��4o�]�<����#y��:�L��Viq�&\\�<�'�@o�2]�m�*Z&Q6��b�<s�Z)�d I1�N�N0æ�@\�<���L�18=�0�^�b����d"�|�<iA��'��l��͈�/����"�{�<1��VY3V�:���#U�m���S�<aiN)/v#T�Ef�ɉ �It�<�O@z�j0Ȁ�C:��%�@o�<���S=E*�(��1+D�s�Ig�<�g	�>�Փ$��
�ʵÇO�G�<�� T:3�Nɲ��S�l�:L�jj�<����W&@`B��S�.Ŵ�:���b�<!7KN�uq�8������� �I�<!W���U�YI�M�� ���$n�<�R,�oh�a��.d7��ᆩ�k�<��"<	��h�NV!X;Hu��ŜA�<Y�mZ�v��r�F�[���(4/�s�<Y�dH��8<U�|��$a�n�<���1�m�2�I+b��q�C�<	d���xㄢ�%�e �"��<a�h�'.�*pZ�(�O\�y�Gy�<٣D�4��ف�آw>�52�Zq�<Q�MW]-���$K�v�Yq̂E�<�KݗSઈ��Vc�9a�k[A�<1�Eçx4�S�J͒}��0E�<���)u���i�cʘ�����X�<IW�޶q�\�tnǘ9��p+`OP�<�r��%#^r�d�Z�o�li�d�J�<YQ(ΤUv�;�.�d�5�6��E�<qu��3�*LPO�zb�	C3JCY�<��C��6�gZ|�T��X�<a��<�������T��蒇�m�<9�k�hm4! f�dֲD8Ĭ_�<)X$�E����H|�s�H]�<�"�W��B�iE�c���6�X�<�d�ݦR��m�0�	J1��
W�<��I�D�by#&����`�g�y�<)E�еq�B��qf�#2<��{�fs�<����rp�B�7���CpˎW�<�b��i�BY�@�r�c��Gn�<IcJҾ 1T��@�G�Zl�rʒi�<a #�\]t�0��TĐ�T��c�<�+ǣn3� �%��e��YE�Nb�<�ũ�!(��
`)�+tG��"b�`�<A��0�dT�I(50Jmbӯ_�<� ���f��'7��Q(�G�~*}�"O&��摆%�}p��I*@�Y��"O8\���rj���L̈J�N,{�"O�`�#�H�^�P +̧i���Q6"O�u{��bh*x�U,r�X�"Or��qd� A��G�K�����"O��Rϙs��!qAQ�y�Pr�"O��х)�((��5c#Y���Zg"O�H{%j�7)�2h@	'U�8(�"O���;CX	C�b:6U ���"O8	���]>�0t��O(S���"O����kܕ:�&�h`"�1(oe��"Ol�gc��#ͣ��ݕ@X�ԑ�"O�4�$��`�42!���cP ��a"OnqQ�g�>t��QI��a?�q�"O<�
t���Y"�˄G�&&/8��"O����X�O������E�u��*"O�uV'ƹz^R<�نPX`jc"OK��/ t)�4I^�)�7�G�y���m�#a�'wˊ}��W:�yr�*�rl����v`b�hC�W��yR��l:�q׬�(yad����y�-6T�ӱ��!I�H:�.��y�c����+Q�n��@pLͬ�y2j��Qn�y�a�/2�6d!���=�yr�­UhLJG���&��0h��yro�y����+�2�f�#��F�y���C��z������aG���y�j�$�^�R�Ņ�;wPy����y�H��-Ր���Ə,+vH`dA��y���=�Ը���"H|�3�aS��y����l�wM�o;��Agܚ�y`D,��0��V�nA��#�'�y�� !�fq���U�Ń6Ǘ��y��жmZ�HM�U���6����y���;`�2���&3Fa��3сһ�y⍆�^�a�w���.��Q
���y2H�'Wr%��8zZ�y���y�/\�y� 0���N��y"f����(E�:t�5��L�y�a�Q����+�h�^��h˽�yr+�vu�$���g�<9B���
�y"�M�w�I�d��<0O�$AR!ϸ�y�m�`��Ѧ`� `��ґcW��y¡O(G�,!Ċ�-]��{2l1�y�P[��@E��j��1 E�;�yr��$3�<�RV�z�"�i\{�<�N��F��J�b�?'�D@Hԉ�o�<����gd.5�͑�@�	��
�A�<�'ΚQ���PǴ53gc\6RպB� 	F!� '�S���+\s��C�	�2	B�pSj�9Z%ʈ�q��!6� B�	�>�� WI�42�\jA�]��C�I�x�f\07�L�C� ��!�C�J��	1�#�8������C�6IL
q���di̬$�_�$��C��>v��A��ﮜ��pXC�	������(�O�}�a���6C�	�q�[ሚ���piA �+2C䉦G	H(P��[�g=��x��W�N C䉋j��B��H�a��Y�F�Ӊ?y4C�	,���[3�3�D�n��%~ C�$Cs��E�L����h1&��c�B�ɪ}#^p�,�O_���GE�e��� 0Ds&m�����J��6L娕at"O��!0
��̈�P ��"�"O�5�g�vCd 00`�H��ѳ"O\(�mT�',v0(S$B�v�d��"O�����ݶ3��:W��EEnB2"OB$v�T"&�h	��F*}%  a�"O���
.(��|��̀�tԁA"OZ̹������ N +�Թd"O�����Ħv䖸�Cm�}C��"OF�+�@�	
_t��+�Y2���"O2��Bf��J��Ij�)�B�"OyKPыk�-ҕJR�i$j'"O6IDG�5�6��V�I�[��r"O��pDN�9A�vq��j<��
R"O�d�P���O%3�^�Rr"O<4�v��Ix��&��g��RG"OT�kw�V�p��`$fQ�^�(q��"OV����d�t��d�
�+ڶ��v"O>�����2��(Bf���Ix3"O���C��Yh�� �'�35a�y;"OP��@��*U>L)�&ï/�@�h�"O�IPd����U:Vȗ�E��S"O�U��b�+[�~� 2(C�=���Ƞ"OtE�^
���ƞF���"OցAS�C�suͧ_�lu"Oʰ���
pIDX��N�۸��"O8|�̘"$����Zv��$"O �2,G�l��u�}W,��6"O��#
T�.�m� (��2��11�"O��[����$�y ��D;7/<["O:�B	�)?-U��D�0ŀ�"O����g�?\�u��Jجw.B���"O*	:�c�'3�,Je*ނ �t�B"O��ۡ�7t�����n��5h��!E"O��x�l�,�T)�W�1FkB�Z�"Ob�5F���p��'��HL�Y�"OM��F�Y~%�Ї�(YE�ɥ"ON���a�yr�}#��]'����"OH=��Nъ|���Ɔ7�<ٛ�"O��䝝@�6��?F�Biq!"O��Z��݊
% ȋ #x��lr�"O�-	�g�;Z�aq�E�u5���C"O���$�#	�P I�KXh)Ԝi1"OZ�c!�?M}���7HY�@H�s�"O<q`�g	o�f���ƖKR�-9�"O��f���4���Q��z6 l�r"O9	Qj�*��P���%/��Ҵ"Od)Z�҉#5P(ufM=n:0|@�"Of<�E녱!j�E:dFY#F�3�"O��Ʈ�w��J�%�� \��"Ox8�ܛY���K1N߈���"O��Iҳ�f����օX�Z%��"O2�Z4�9<А�4'Y�S�rM�f"O���i�;֔u�R2,�BIȱ"Oh�#P�<��	h6	�0�0�R"Op�;�e%,4�w��	|s\���"O4=Zs�#	jܜXS6
Q�)�2"O�A�C�X7K��/,uD���Q"O���Q3,�|�*7�QF: �a"O������qc��ݙe����"O�W��'y��¤�\��a�Y�8��	/��T�Z;N���â��2n���$??��.�6k8vQ�a!������t�P�<�/D;awڍ0@U�I��x	3$P�<� ��C�����0�A��/Y_2�h�"O$���钮e�\��oB(R[�j@"OH��%�C`�|k�-�9d��\�"O�2�S�8or�HQ*&���!"O�(���wIJ��Χ'�,U���'	�IŞ� �	;{5�pZ�-}�4��F𘭳!��3|m�F���B��/�A���Gg"��[A�<8�+D��;����"�r%:��O&y~���(D��	#A��&%��Z��N����2D�����G���a���L�i9��$��æM�6�<���F��*�P��
�ز�V�<I���˸M8�m��g�Qa�ʌɦ����c1�݈!���V�Ȗrm�E��]�f��B(�y��q�%�^�̇ȓ+w\�c�ŝ�k�xhB�Ő�Z��?���)���(>2=���^����!d̅�yb높 �b]�#" Mp-rT̊�HO��$��-a�3�BT��a�х�'5�!�@���87�9J�$U���D�s���?�S�O]��0&�O�}�����#H�a���$)�|*���B͗po�x�xm��'��}���*L�.|�E$A;& �h)ЅC'�~B�)�'i>F4��ڛ��e�%P�`��Մȓ}�VU" ��)��}��L_5oz��)]d�"sOP�,;�({gl�4b�J���pLL\*����41�!�҅1<&�����#u��+�F�5�Jݺc���-��B��f�4@���;4B! 1�ěp��B�	~�L���-̌*�z�"��B�I �Ѕ�4�"|X�	�+��B�ɂq" h9�l�i�0s��_�&ynB�ɘh�j�����iy�b���`B��4>괠�bC�4,y4�� .�,&M"b����	�S:��`��j��Z�FX?+B�I�^���#��$�'�J բB�̦��(].��]��C��5�T��*���Dz�ԟ��d+}b	ʓ^t�tmػm��J���y��7a�|��͌����$r��`<�3�)�S'!"ڕ���$�0�y(ӮE!����ծ�?��4N�r�Hs �bP���y�V��'���O��S�L<1�쁸aӨl��m�8�!��M�my�>A�������Ӏ:��)�E%�9BN0hq�X��}���%JɞG"J��Ц�^E�`2�`3O.6�5�pl1���N4�� Ц��lƄD~��ӥ%
�C��9D[� 	�Q�@�O�=�}�s�gS|(�Bm	�0��h�nXA���hO�@��ȁ����2�!Z�����'�ў"|U`׈�
킶'A�O$�j�~�'�ax�lߢ]����`��<��H����'��{s��qȶO�ZdP���-�0<)/+ʓ=��t�v�S0~���C���|b�?�y���O`x�9�a �!>8<,0v��*c�!�$�.`��	�#�SE"�:���M�'.O��<	�� �N���K(��A������x�gX������l�@��=�MCO<q�6������[��8(A  4�>��ȓm�f��M�k����N̮���g>�)���#�Id�+y,@=�ȓV�2�7s���J"�ܤ�x�%��E{��d��kA8PBӿ	���ԅJ���'�ў�Og�ۄA� �$��1�B9 �O����S�L<��f	/J�ūPFEf�r��aJ�P�<�M���mq�E�ax�@���f�<� Ѓ��\v�d��@��='�*Ȉ��	\�����O��&۫kk�@��V�8��d�U"O���š��8��F'Pq��E:S"Ol��&��q��˓e�
��T�R"Oj��q]-1����������z1"Or1[s+�m��d��.Mtp��"O�l�祏.vE�Ya�-6\���9O�����O�܈�m$>
��Q�U6;PX�Y��'��'�|�#�#�� "U�ɒq�$��'fY˓�G�]�be�4�(iO@���'��c�bTfԶ�jMPW����'cX�(�g��o[��Ja)��"&�P��)��<)q��,#݆h���X��b�ej�<1T�R'8� m�"_�@+��Gh�<���NCj��1��;K\x+$�:�(OT�G��O�P�F�]<l}}��G�e��i�V"O��7�T�H�y:��'p�^�3;O����ɳ+3ޥ��T5Ii2�����,Tv��DG=�y�?O��o/��h��@�.<m��"O$�m��YH��¬A�@���"O�y��)Pq������͔5��J�"OXp�T@^�C�F��AՇj�<�y'"OR�i��U�/:.`ȑ@V?����O��J⍌�V_Դi��W0��r��c�	t� 
-��<�R�rgΕx5�m�<<O�"<�Dתr{JA�/��Z�[��L�<9 ��v`�A$��X�)�	 A����<��{����C��WM�(y8����6�yB�V(%�0��[�	��� $�y2˛�S�0|��0^�UH5�V��y"+�5@1P�)�Ĝ t����څ�y��[3Xl�YP�Z�le"F�^��y���sJB`�2����%��!�yR'
�N�ă�38[����L��yrP�>�4�ڀ/آ1����#�K�yrM��4B��x�� �%8
x+cM��y�̅�+�l%:d����  �mJ��y�,Ϫ$��8kĉ�e�]�*Ո�ybb��.��}S��(oT�ۖR��y��i3(U ��4V�<y��!��y�ꎳt@�;�`�"u�u�/�y���_3|���M@�f	�]�ӡ��y�.˰+�r����'w�p�� ���'��z��G�l[��т��9!�����j'�Px�Y6��uC ��
>�^����+���|�sN0KIK*��e��G}2�@0�h�ddC��FKx%�Q�Q0=S�"O��g�9
��ȃ#.7۴�BT� ���铕9�.����)�@|(YNw,C䉀6!E���	t����
yF:C�ɴ_E~li�'�3oA^"�E҄UF.C�	;2�<�p�O�
��$N�-��B䉌J����m�5R>���(��B�&`��`�jA�B1zP�ʳXfB�	#9��U+X�%.�عG�ǵf�C䉵L��H���X5��84-��E��C�ɼ�9��bP*n��%E��x�C�	9)���� =^~6�K�."ێC䉷�-�b예HvĻ�*ݰCLrC�I3s��ܣ��T�e� 36%�$adC����`W��X}5���!spB��-���C�;̀�d/O�)�tB��@Q�M90H$��iZcμo�C��|�Qp,��v���Ӕ��9�RB�)� �!B0��)�ё*��3F�M#�"Ob�!%�RX�7L4,����"O�ER`��e�d�l �&p�9�"O q�w �L8�<�W���jڹ+"O*�)G��t-ŉ ̦@�h�	7"O�0b��N�q�fK#@���"O� 9CD�E��bÆD���h�s"O����ɢB�Je� f��q�`<�"Ot,�`.�����J�,��B�"O�����'�|�CC�t���1�"O���g��u�@`�F"�����"O��R蓻`'ָ�� �;�V�k"O�TA'lH��v�bRO�*���"O4��u-�9�anǴ���"O��"��YAk	��MU&C��lP�"O�B��G�ClT������-��"O�M(����� ��,'i�1��"O��
4��9Z�!w��R_��:�"Oy@���*3*�,�H����
3�!�d�5,-�x���9������Į�!�$O�;Yč��O��"%�4�X�?l!�D�GO�0�S��p#5�ǀo@!�$U�^�!�K��BP���"i?!�$?���AP��:!����eDI#!�^	Zt�sD��	T��a���7!�Ѐ#�aql��3����7�!�@a�6$���P��D���\�u�1O�x��	r�8iV��!p��P�ɠ��}��hR&Gԕ06���!�d[�l�	Z%�s0dmr�O�l�!��%;Kܴ!���.��`�B���Jg!�d��% �xK�A�y|<�b���.Z6!�$�L���ᅐ�V�05ȐD�=I%!�$�!g&����"ԛB�b�C���	P!�D�/%c8�GҒ��g��t!�DKd��h*t%څ������ !��N�>0���.�h�R �C�i�!�܏��`���N���ի�n�!��H$��,�`%W���ɟ�!��+n^�yDh�>��������m!�DW#-�p(�2��CV�M��+�/
!�䌪uDҀ S�L�Q�VA���E�!��
2����6"��C���acG�/h�!�d[pe�dgB�#�`<�d��c>!�dU���bR����uS���zr!��)�Ɯ��A��|�	��"�&6�!��N��p)BCmF�=�>-vAPE�!�$J�9���H�ʊ�Q0�����j�!�$�^�B}��)�$uq���(3�!�ǽ�h���+LMjpIbn�.[�!��:7$�ݑc+�p%�;F-�25c!���w^@��q� 5伹�ce\!�D@�?��ɒ1`E�L��rP��6A!�=2��bDK��,2��"��cn!�d��d0��`sY7_����⃈_!򤉴JږII���X�4/�U�!�$I�Y7d���Y-��چn��CJ!���#t�P��AB`�E��
�L!�� �ynqy�O�4��䓆�L�!�Ċ�":��c�b�^k�-�@�@.9�!�dL�J�B!��o�p���_8w~!��߷U���Pff�.P���AN�go!�B��Ne��.�8er�-᪝9�!�
�>��ȱ�)%	�Z�i��ܡm�!�d����U
�
��G��=Z����!�� <!��g�H���Z4�v�$�S�"O\�A
Ӣvl�AJ6�_:Ba aQ�"O�Y�/<8�&�3`�;z���"O|��bZ��J�#%��,���"O~TqDiPvz�yd/��o�X��d"O̭Ya%�?,5zQ�-DxU���p"OIq�f��\�`�d�Pf��x�"OrA@��;(�^�	���d%v5 �"O��)��B2u,\�����7,j��"OVHQe
3<���@����b�"ON}{�,y8X�3�����A*�"O�	ʤ��&�`@�S��p�)��"Or9	c,�2{{h4��aQZ=Pr"O���ą#&M	a@E =J}�'"O4EK�/´%�� !��-�ek "O��Hq`��UK�,87Kl�8h�"O�I�甁C�bXk#��w�B��"O����mE��s	�MNls�"O@���
UX�k�W]͎�B"O��!��Q==E<�����m��XR@"Oh%���oN�Yi@��'�8\"O��p��M.jVLH1φ�?�,�W"Ox[R
I�E��(��_��v�8G"O�E�� (��Y8B�KR@��E"O�@;b��K6��A���JRApR"O,���� 3u8���V��L��"Op�E��#4�����PP
u�2"O|�QB�	F��e1RL>F�y7"O��!&O��	�U�S�Xj6%��"O��sۥ4kh��5" Y~,J�"Ox�r���g�&9[�@��L�L��"Op�he��W8I�/�/jֶ]�
�K[����Ծ:���zc��G���"�B� R�廣Oϭ6Tl�r�E~v(2��7�"=z�B�;�0E|��ϏG#z��F�%E�v@� GX:U��f6^,�0��h��1B�O�<i�FX�;����H�60zP ������2Ƕ���â\Z�o�O�� �CI>a��`�RE��a���"O���U�u�@�cX�e���&\2L�H]zG��e5���NA9}j�y�'ښ�8C��0"6�IӒM��d<<!
�a2Ab-0���Z!�
7R�N��O�*��	���@C�ā�0>�ҮE�eF�<Ç�!^	 �s(�A�'��;���#���҆�V�D� �P0���u'�y|z�'JNH�"O��wo�4b�:��V�ͲI!����'��Qs�.B�k	���MB��W��=]h�Iu,	bp��5�]��0  �v!�8���� �
@k>TB��n�͡�	؍J��yt��g��	T���ьJ]��-�GH�8�"��;�: ��e�A�T��eI�1\�}�rjƙpq���[��E9�E8�O�@S�CԮ~9 �ۧڣ>/4����	�4� �hu������
Oe*��s����둀G�2i� 2{BB�ɿ$�|��`�
1�e�%΅�
�����-��p�Ȑ�\�V���P?���|D�F�ߵ	�|��䐯�b���$D��2 C)SY��H� ��&��0 ��@}�$ƃr��U$A)\:�?�#��1U��E�4�Z�j�FCPx� �6�9.| 3c���o7R�+��1nD���1�L���,z!r�̔j2�,I@��-/8��E{"�˂[�B	c L�'
������.8U`PBl%�l�ȓ1�0ɰ4��n�p��J�M����	�I䘼�&/�&o��S�O2��Qb�
w%���"*�	�"O��y���#H�L��;�}�AQ����"T0d|� ;��'Hv�����>r^��І\Mנl;�Mժt���h?nY�o�0k%\��@&K��=����4�r�� +�P���	&����bP�N��I���d� �x Ś(�t%Ѵ!R��\ܰZ?Q��KJ��EXfH�>gu�����HC�<�@I�ID�dڃLĂr܊qi�t~�'و�Ӣ*��j����Mx��@`�۱��� ��K7�ʦ8�RM
���#T:<Ѳ�'n0Z�C,i���S���1�����`�?-Ƅ��ea�Z!^[#��^���0�V�z��L�@�"@�p��J�F3����)������I��

ab���ķ��!c�T�$U~Y����p�R��bn�4�T�r�7�O� ��@Ep�p��F����c#G �I!ė�u�H�h�}2�ӑ^'��z55<r�I�44�SΖ��]��d2C�	9iQl�H�Ǎ7�@�a�il����6��Vx��0�LV�D�6�X���	�2�0�b�-�|�B ��Q��<!t��t��h Rq��T�ĉ�.G ����
��ΘsAh�>PdYP��S;4�c���N�O.�G��q-���o���V��"�z}��#�<u����<��C�=v�����k�d���W�ħ6'���k�m��;2��L�bdpQbYj�x���K>�OvA#e��k�qc�D_��"d��Vl�H0qƝ�bA�%�5�)@�S�pڈAgĖ!9���8b���$��:B�p<zbN� '��C䉀rߴ9�dDY�^��bH�HS�0��[�AP�����.����ԅ���SZ	�C�ʒ�:����`�����J������"�R��|h���LA~Q���*"�4����"et���F��:�J7MB�/Ed1J�|�.�S��Q�3}B��-{ :%q �=x4�e0�L���'5�u�L�(���������W��DO��#�&i���6�F>e��p�i�?�ti��	�R�|T�d�R� #HQ����=�zIjU��'�u"b�
V��)�O3��R�#+\y�g$O��$�4/�5{�i�Jt���G�@�Op!�d�]���7�:h���G$��pv���ߐ}꼍�VȢD �0qN���G���B��?%9��ġQ�$Z!	P�WIv�Z �2\ORD"D(����������BH���㨅.L}�6`P�~�'Hm�f�P�����D�hrZ`���4i�������MkqO�DK�N'6Hd�S�'o���@���
Mf��͍+����'�-��yP�$֑�0?)�D/Qc����N<M���"�p%F�"E�Y}�����d�O0,E��O�z���ɜ��� @9-��5"OX� B.O�oE ���nɩ �H,1e�iA��Q�H>_�9U ׉$��xa�UXՂ�u�9�$LM?��=Y��]#M����CܾT����Z�e�D�[GLC(R<�x;��>$�X�Ҏ7'al��ag�q�3" ]Q����ZwϾ1s�Y�i�BNP8db���Ŏ?@�(B��#�̰�fG��P���:��П.�"��L;hwf<�{���L)et0�H#!Q�T|�d����OTC�I7R[������Tưd�ֈ
�JC�I�$�rP�!&THٳ�[�x�*C�	l��̰����n;�UB@O5�C�ɺ
F�	b���u��٨ h<&C��ld4��@ق4����0KC�	'
�V�x@.̓.�j�#AJ�*\4C�I�q2� ����16�3(4�"B�0G4����?�D�Ct�Q�l#�C�"}�B���e[3P�4`��*S&N�C�	1��TpB*�')��걍ͤCU�C䉳:�B ��C��iS1�
��C��&mH��p�;5��H���Y �C�ɰq�(���*��Z� �7<w3�C���||��B�i|t�)��3)��B�	5G䬠Q�P�R`�d:C�	�I�F�3���0A�:-[�&�|?�B�]����n�	@�5l5n��B�Tn��ӌ,F���smݩb�`B�	�y���BI�
D��'G�i�\B�&Fˈ{1o�)�pds��׳(��C�ɝ/���R�'��6:$Z�)� x�C䉎w�I*�\����"D
@�	}�C�I�4����P Z�[�U�s&��7�C��%e��9�����D�:cƛ�Yf&C�	w����O_��Q*��+C�I*=X<����) �<�`˗�B���jPR�'p�=a$U�3ޢC�	;^��Q�FZ�1[���§~[|C�� 
��M�	�!�MC�F��A8C�I#Ǩ���/P's�ywo�/f�C�)� �h��I�4��ah��Px!�"O�� r�M �zM15�\�`B̵j�"O�����+��d頨�6N@��"O�q����$8 ��T&
�� u��"O�̈�NN�1����F�T�|��""O����KX�wN6���&�%E�:�zC"Ox���+T��\���J, ��l��"O��,�_Āa��ٲm���� "Ov�sgŌe�����C[�+X�y�"O�����W��r��sO�	�"O>�{���/D�z��B�� W tuH!"O⥘�nP�T��uMI�4}���"O>U���=k��تt�̺s0:P�"O��Cg���EV�J��ǳq>�}��"OY�s���T���C��1D���"O�p�&I��k�h�c��֊-f�S"O�  ��E�L��>ax�5�@"ObIygcN�8�J͠��*	x�xr%"O`,bé��d?@� [!p���p"O�d�@/*=��t���Rz&�y�"Orc N�w�����Z
E��a3�"O>��e�:^Kp�CW��.���r"OVi�OޓG�nܚ��ǡT)��Q"O�d;�
ŻE^�3��K:Ƹ�"Op$o^.%���e��1R,��W"O�TCUV�o�|�b�f�8�$�1"O"��&Ѭ_��<zw�=}���"OƑA���L�qq7���p�"��"O� Y�	�"���B�F�L�t��"O�M[�gЪ^�Z�f)["=2`M�B"O�b�SA�ly%��R��"O2u)CGD! �=����u�"O,���5��܈��ƴ�P"Oބ�5#;|F�Gb��U�t���"O��:E/҃��("��I#}�*��t"O>9a�Dȱ;+����ʖW�2��"Oޡ[�-�?tP� �N����1�"O�1�b�]�&Y f�)pu�y�"O����#B�#F%����"O�X�mH�^]Hx�Q&ц%�©� "O�p`'��G
�9���#-��1j"O.P����E���˂�,bT�(�"O�)�Q	�7��Ѐv�M4APt"O�ȵhG+4���!�6L9�Ƀ�"O����aW�L��a%�^�N���2"O҄�Ph��o��&.Œ.��t�"O�,�`E��9Q����� D�L�g"O�a$k����Ҡ�0��)Z�"O�%`�+Np��eԯL5� ��D"Or�:��X':���@���+6�2Tq�"O�Lp���!.p�yыM0
è<`"O����C�~��S �U(0���"O
��!���n�0Dꦦ@nɳq"O0�jԤ�%m�`�B i�@�� "OV��A+K	Z�-[��}�����"O����+,j��o�"vD H4"O(mk���}�A����o(�ڇ"O�8�Q@�&m����lZ�$$��r"O��+��(iO�t��C�|r"գ�"O~�@өJ�\�F-H#KD\�B"O�9�pe�?D�M�0̜�"���+"O­I`��^7������W�L��a"O���6D2)�Vtp&��"o�T�r4"O,<�����d�Ū�w��"O� ٫��2x@	����y�Pڦ"O���ģM�!�p�a��Ľ��(�B"O��bw�H.��R��Lu�p�"O)�U+��DL(�Y�%���"O$�dF�%\o��O��M.,|��"O�l�� ��V��B�#|�T�"OXb�`��������2O�pp�p"O�E��]L�u��Ϥ �,�S�"O�L %�����u���(1s�"O��r�Փ(�ޭ��,�D����q"Ot��Q"1�J�"���У"O�W�K�Dt��!,rr�*u"O�dF�Y!���a	�l�lH�G"O$��W�%5��|��HS��|�"O~�@�͖ �6YG���^n���"O���*]�R2 ra��[�"O���KK�*9��bг,��}��"O:���A�)0�DO��,|S4"OR!���;!fP3B��d�X��3"O������o�#�A�O,� "O�q��](]�����913��R�"O�	zG�����q �7])���q"O�k Mԁg�H	��� ~L��"O �0�A�~N��1$Où~P���"O�Q�C�s��l�"`�5GL�"O~jF�ܸ+z��瀕?�X��"OX�Y�H�:]���Qg�5)��p"O�z��l	Z����1���"O.���O�g@�I�8��\;�"O��kF��v�Hi��L>l�*h�S"O��x�-��l�,*�lӦC��iѥ"Ozt&?!��l�� !�� "Oz��#�T)��]  ~V�"Odt�v���`pt�U�yK⭩@�
E�<�ӈK@:�m:+݇e֘)e)B�<��@�%sk6x""(�KX���&�y���YT�$�D��Ew���G`�U)�x�5��K��iAT��hX������"_���a�^.A�,
`!?�t��Ez�KԶ 3�ū���G.��=Uސ钗5��\-j@�$"Oh�7=�|���@�	Ft�k��'N�e��.G�Y����;E�d���q��0��'ɠ� %��V�2(��t1���׀T :W�B&ؖaWB����
y@�E�"a��uY�e�~�4�G�H������H�1B�,C`<����@j$x4iT�02$�0�"��B�-�P��͚���ʠA.�O� ��네XB�EӅ!1uD����ɿ7Gd�B�iu�jQŢMT� �ϧ}�����O�+����o�k�a��w�Yh�#��TGjQ��½�}lB��!�J-��)ޡ���� gE�O��V�)M�Ε��Kc�j�*�"O�0�p#U�D�*�b�8j�>y T��1=B�hT���F%���v�G���A�'0čc�<p�#ǤK�nV�m�	�oS�E���]:
x� iGM �aK��O�?�T�a!%�xx�d��6�0>1���3[�H5�N�T(^l!B�JJ�'+��9',�$�T�곤U^�X��O�&�d�i����fj��.���'�:��v�Gj�nhsF&G(0���s�jbt��k�dc|�*c��>V�8�~��*�45Ė�Z�DB6Pjr�F��yR�!1`�b�ķK��=p�;^4��3:!�u"e� B�������վ.�ɻ��٨���Sd�RF�}r�ՉWJ@ݻ"�˹=\;%�Y�2��P�Yq����R.D<�D�֜%~~��g.����O�W�']6�����qJ��~j2 D,�� �D�.Z�hׂ�M�<��ɛ.�T#�����h��Jȟ�� H6%4��>E��f�NKJ���ؘff��	�B	�B�!���h�:8��C��vIa���!	���' ܊��L�U�ay�hWe���Hu �f� ȚQeN��>�q�Ή]�x-x� �	�� ;X��Aa��U���g��{���'Yr�H�
�"��� �F(�x ����Z��t$�A��(��|�4��x��!�ʄj#�hPL�a�<�v�8�*�q5�D�jM�tN�X?	v�8$(\CbFs��`3����gy�t� �ۢ
6e� ͳ_?!�
.��s)T9D����&Ğ�:�X�R/
P��<}"�?�'�j�G ��5�!@��ܡJ�'/��*��_�<�����b̞S��q5%ά'��%���_X����,��S��E2��L$i�@�P�+<O�Q
ga�"c�TڨO����ޗL"8�sjO�	6،�e"O�̩�Ú*��5����U�R�H��|�`öP�J���H\�O�̴X�Q	a}v�K�嗋���B
�'�"�A��.^}0�����+@�ՠi����'������>i�	.�tP𮘃54�a`-Lh<1�g�D����� ��к���
~��yT+�>;���$�/&�,�J�(�ɀ���x�y�� ,����LSS}B ޗE��J�D��w�r�"��۩�yR�^>p~�T���ƙe	8IBf	ܘ��d6a"��]<��#
@J�>q�d@�����D���*v��<�2�1<��ٓ�?4Ѫ#
�+D��>���2����I�{q��˘Vԙ��
T�
�B�ɘ�h���.p�[$*?��q`������J!�'~����ȚRO�Y�-W�X�
�
�SK�	gmV�[��u�:�3��-���Zv�ԭ3�>X�ȓ_��tx��<,�x���(%|��	%��ɠ�Ƥ�������}('��$���dal���	�'�i�4DD(M��eA�2<�$�Pa��KB�'�4ˈ�@� �4[�v���o��n�xX��<D��C���0Z��5a�H�"t�A0���d���E):�OTI7/Og>�K���%xV���Q"O�q1ߴm���rU�=O`�P�"O<�B����[��tx�ď�A7� �'"OL}�#��<L���DL��:&"O��(�	]��u�UbQ���"O���g/��a�H�(bBƛز��W"O�ua���(�t�Q%�lɂ���"O�98��N�N��2����E"O��Y�m��u��CD��8+����"O�Y�B�.C��A@��x<�a"On!B!�yV�;G�[�
;4E�%"O0�R���|fԀ!�A=~""�d"O�1B#�*�K�c\)|B�s�"O�%�!E�<o@��`�-c��r"Ot�T瑔>����O/A�!"O��ţ^_���T�@�~,��"O��zt �?{d�P5G�'��5y�"O�8hI�,�F��c�ȥ���W"OH-���]�"v�p2���V�D���"OV��!�O�axcbƙ?1��"O�`��-9xi�'�De��ش"O̐!��V�=�؈a��0��P��"O������~��V!K|w�St"O�rC� <F��+��@�j2�9W"OL�s���:��(�磟02�n<�"O\���F� y���AɾE���9�"O��b-(O��I��Kv2��"O��ҳ��
=�\aƍї j�5"Oh�K7��p!��b�S�:"�Qu"O���*ǧ~�D��%��j���)"OZ�q��Τ*}�1k�"��pX�r�"O<`hP��%:��QS�Í\o���"O�4�NטZ�@׍ڰ@�Y�q"O���E)Q�
l���3NH$�B"O�s'MC�}��H!N	N9088U"O� ���M��j@Z����X
�mKS"Oh��k�>�i�������G"Ol`�tE�j��M
7��K�y#w"OV�ЗlP�7j�s�!�/�~q�"O:��� X�؝je�؜>mz<�!�$�i�l$r$����ZX-��"O�Q�k�46�&�`�ኲ`�|K&"O�	�$��0�H�d͊:h(�9��"O� ?=-Э�1ʓ�k	:�E"O:�C4(fHw��21��k�"O��	E���R�K%�0�r��"O�1�r�M?&I��;��G�(�t��"O�Q�i�M���DO� �qt"O��Q���\LA�N�-Hbd%�e"O��9�
�4@�꽃�L�X�謲"O\��A�Y�bhȥ��(2��4"Oh�`�c�;A^�;fHQBhx�K�"O��hb�$vc�:H�Dt�xQ"O�Tȅ5��T���� )D*�"Obd�Q萴I�dsf�<dD��7"O��#�ջQes���m�"�cp"O�< HTuX���R,r�QqQ"Or����)\�Y���F t���"OT�S��]��T��B	<OpMڑ"OZt��7/�D�!E ��xGҼ�2"O��P��
Qj��� ��v&q�"O6��l�!�~l����8��@�"O(Y1o4JXD�IGB�<粩Zf"O�8�7Vmڭ�3a��B��\[�"O�Y�Q%�a$iA�`Éx��$�@"O�0Z�	M�/�ĉ0,��֙��"O�m0Ђ�"6�DȪ5B��e�x��"O�l�k׋VH��a5��a4�=�d"O6���8�Z�AM�K�"(�"O\k���B���GM�F��`s�H�A
���/�2dd�Y� {�1O`��eCS'x������H	����"Opp�k�-�+��h���"OD�k �Ͽ]�(h��D˫=�ٳP"O����o�<!Ѳė�/���Q"O&�{���vܪ<k��h'�`��o�?W�^b��G�E��?Ea�aA��R�X$�4PA�����'@
��,?�萻��һL��Y�ȼlϬIIw�|/�<lήc��)��)ߴ	vde9b�'�B����N�#��'Q��e�O&:،(�OQ>����
&�`���sV�jI�O��h�*p?h4�!G�<E�4�]�IKT� �[_�`u�c�\�S2�ѓ�dU ���-OL�����^$���kŏP^aJ�������Ub�*��ɞLh\�ᓩ@� A�/.7[֠�+�
x(�T-�<Q�j�.4+���ç<����E!�"J�Rd)"H�!+;�\�'�U���A�]�q�*�'�M���LQ�좐�B�!�
L�@JZ�<z���
(, ���d?E�TOQ?}1��&��61]<�D��&D����I1n3�i���O��iJL~[wF�'�ƭ9w��+0hY��@;��-QK�sf|Q���mq���
�r>��I�*�Lh��G?ܞ\y�.x�>1ACe 	���`�+n��ᓫ(%���p�W0:}���4f����BB��~1	S�4��O�:Cf�?��Pr�iQ������ 3e4��'1>IU�Ϙ��Ӟ<� t�(�)=���"��\ �O���d�o��I� ��r��n
�!�d�)�^�k�%�14mpy6@^_!�䎲>n`(�"F�P�"��7�!�DO�O���xc:*��H���	v!�d�!X�b���/���Ν�%�!��.�p��,�hm�c����T�!��"Ґy��B�VX5�S�o�!��H�7�v��7�B>W.~���#X �!��z��x��2{��i�bT��!�� B��Λ�3�Ԕ��/�5 !><b�"O���O���L;toȴe��;�"O�$ٴ.��?���ʲ7
v�*F"O� 0�I��8�C�@��p��"O�@��E����z��T��"O�=��G�{�h#Ǎ��к�"Or�;��
� ݊�[ G�1E�F�J�"O|�����^�@����l��0�D"O�Is��!wzQ2��In	��"ON�R���YTa�u@�?u*�x0"O ���O<s�>��i�":�$�"OB����ۀԖ���.;"��:�"O���&�!�*�B�Îol�X2p"OY��Z����unյ#},�K�"ON������~�F�{d�E�Ua>�"6"Ope�#�V�d��F�ڰF���p�"OZ����A�A�e��͕0���s�"O�� d�/��|R�
*�D!�"O�*ףK	t�<\���Y/i��ٙ�"Oڜ�U�F/RI����b�R�R�"O��@f��:��8)Č�
B��"OD9RA\�L�Ҭ_�@�p��#"O�X�D��J튴rtfy�
��"Od5jv.ŋI4 ��lx���"O�u�E�*�8����,p18"O�9�1գ�n%�ğI\EA"O����y���mU�Q1"d��"OV���'�lӐ`�j�7C��G"O��@�Θ�s�X� ���Q��`J$"O5��1�k��ϒA�L��"O,����"'�4�0	�M��J"O2�5
��Q�tHP
&�*���"ON���[7�:��bI�!)�R"O��A&Ӗ3]���'ih���"O(��U�F�M��{��,+R�\!"O�Pyc�^	�T����o0����"O ��&� �7a̫�(�Lv��2e"O��§$DF��1BBN�JF6��"OL� piQ�~���c��**���"O L��łw�m�P�V�7 4(�"O�y�7`��&�nMcu��C$x��"O����D�w[ �;��1'�hZ�"O�;�\�6:���ҁB��v}��"O�\��.�lRQ��@�jV��"O�Ԧ�]�\U��OV��a&"OF�d��>8�JD��n��*,xe"O�����4^d,h�fF��0��G"O\0�I��(y�d%�'9�4a�"O�,�S�3Hv-s�|�@��D"O��e�!� T�oL�F�5�"O�Yc���kn��8�處3�`ĂW"O+7�V�9���R��V�y}VX��"O�p�`g�;s��#F�$ڪ�;!"O�h���޻78ʈ��D�Y!>i)�"O�=S@�j��R�K9-P�b"O�R�k_�y�����g�L �"O�M��"-�j�xa�O?h묀��"O��kV���`98U��%	B����"O~�)'һ|ߞ$k��\�I����"O��Z���1�Fyz"���а�"O2��$�*SM�bF+����8�"OXɃB"T�_�0� [��&���"O������t����F�Ґ�"O!x�藌o1�I��dY�Vg0(��"O� f���d�6�|��L˽P�(I&"Oư���D�$��=AEK]�%�<��"OIP�,�8|�2�M�4o2\pH"O ڶn�>5��ʠ��a�4""O.����Vpj�"��o��y"O~����@-s�(|"AO��]�|8�"O����� tll�"�Nm�4Y��"O�Pc2���g��9W�T�]M���"O�%
@A��TR�oAMH�M��"Oa8��+0V�M�L��[�"O�4[eI�s���C�\AM�y�"Ohi� Z� �H��v�7�Q:�"O �L�$\�n(��#C�ؙ�"Oj��,SOl��s��MA"u�"O�|�%�鶈�F��d��"OL������(R�/�#RP�[�"O��ӅYO�%� �+LE,u�"OX��QŇ4(��){��2 "OL)`B��:Q��R%T9-�	�"OBl�ӊֱ��A�O^�v�!�"O���A��"'��	�%I ���B"OA&��N]^%����2c�D�6"O
�0�Z�q3l��&E��"O�9�$M��4�"E!��U�
�(�G"O�e1R��dz�T獞S!l�S�"Of� B2?�x��U�7�r�"O$%06O��Ss���F��n�t1�"Oj�o&=�i�edT�.�X��"O���2K�Q]�)��
�
�~0�"Ov��q���!YY�&E�P"OL�D���7HH�U�U��|Cf"O6�h@���pR��sAᶌ�B"O�9��ٹdڂЉ�O?Iޞ�Q�"O�U2E�Pf|�20��B�P9�"O���g��t�HER��ǰ�*�z%"Oj=K"���P�b�	��8�R��"O$!���[+�8��U.U|���"O��] �;���Y���a"OZ}�a\�u)v����֛���r"Ov("���wI%!�N*`����!"O���c�
=���-M���"O����:�1�1Cv"O~P��)Uմ�;SA��w�n�Z"O���+��H��	�����"OB�:$F>o�L�xdB�Tw1�"O��G�Z)><���	ca�d�"OFqC�Y���1�-A�R�u�V"O��"2s�(��lҞ7�s"Or���\�>25J���1�y"O:Pڑ ڞ��I����/*<r'"O��*e�Ф
��[R�۬ )8��"O-q�
�FJ`��r̂"P�@�"O����ORF����ʗ�)�"�ڡ"O���M�	]Y���e_��j�"O��s@�Nz���'H�R��ICS"O֬h2㜅y՘鋣�$>|�q�0"O�h�mұ>�(͢�
��Yj e��"ODH��R$�����H?]ٰW"O.a����B"��ct��#L䵘�"O������,%�]z7d��(��t�"Ox�R1h�*,��s�؅,�p���"O�Z�B�k]l)1�+�/�Xܣ"O�`�g���M��ʔ��jv�"O��cH�F"��b6iR�hd$a�1"O� Q	A>l2�ٙ��۔c5^AH`"O���� ���V��u���7"O�a�f\�`�6US���E�
���"OƠ�$�ќ%�2�����(� ��"OTȣ�CJs�Ÿ��.~�҄"O�d�l��J#�-��ā���m)�"O.p��J�5�0!h�Ɲ�[� !��"OM�0KL�~p)#eBB�Z�)&"O���*K�Q3$�n�<c���R"OfA��?"��1�˙�5���b&"OHm�3�ÿ^��s�M\|���f"O� ;�CT&~��k�Vr�M�"O&y���%-�4�[��	�`���kd"O�t��K��l	�#`�;�*)�"O���%�<�:�y�NL*r���Rr"O���e��}�c��X�����"O��[�N��*j��2Rl��N��"O�`d�� 3�F�@�T�-o�m� "O��	!k�3�����]�	_~��"O6xk� �*���7f︨��"OJPj�,8$��y��I�Lv�q�"O"傥%�D	�� ��� �"�"O( �dR�$�`ݚT�"O�ne�t"O"�2+�5P�)����>��0"O�U1q��E���S�f�|J�1Ѕ"O��c���A�Ȅ!��5/�2�"Oj �%��P�bH+��Ŋ>��	�0"O���1���<d�:sD�8h�&��"Or4jW	)#J25k!�y���a"O& `2A�
�l�t��<r��"O�貒&�?_�u1�l% 0x�"On� #�Z�m\���J����"O45�C�َY*r�Ѳn��\��"OI���E^Z��AH� ��b"O��J��Z�GT9��r"�HG"O4�H@�	>��H���? #l���"O@��󦘽=&&-��@ӽ~	�)G"O�<I�f+d0���A�\��dc�"O���,X�W�\jw�F� ��"Ov�8���T�p�F*�\�<Y�w"Oԁɢ�P#~�D�f��
�x�"OR�3a7��������_�fK"O�ׂ�z�`q��fQc�h�2f"O�`y�N�yM����#��!���"O��0�I�7���1 �5l�aS"O�2�!�x��\��@Q�""O����D�
S�8ȖFy����"O� V#.(A#@P�Z���"O���!�Q5�ؑ� �@"u�~��s"O�ͫ!��vfL���C��Zp"Ovd!M"D��I���Pft
���"O����
�u�*��K�os��(V"O�b�"�~��,K'I�� ��Z�"O`��I+w�8��qh˲E�� �"O��� C>׶�q�^�)���"O2D�B�^%)�T)z1�Ψ7���{�"O,����'�>�:v낓6�&���"O`��1#^Τ����
��˒"OhYQ���N�F�*���K�F\��"Of���Z."l�a�J�%8U�t"O��ZB�߮|L�����%Ej8���"O�Qʲ��>B�"̸R�-NO��C"O�WJ������NJG�1!�"O�i���s��0;k38,�"O���:    B+�>O�l�d�4�<II"聁�y��Wg�\�*s+ϵ%�x��f�%�y�%V��]@���b|J�� �yBa��nOHL�1']�c������/�y�c�:`q
%O��!���Y�K �y��ý��bC`�Vu>$���ؘ�y��Dz9pC�Z��Ub ��!�y�DЖ���+��U���0�����y���88 A�ŬM����gU�y�I65-��,�����pw���y2 �Gx� �C�������L�y
� Z`���H��
������"O��G�4:�i��E�8y�Б��"O��Ð�VDp��KP�{7�i�C"O$e�e�ѣ~}&-��C�H�hД�'
`�@�@��#0!�J��񠂄��S��#�/��n�ډ��$0�IʐlZ�w����W�4&`�<��A>1.thR$�h��q�D͑ P[�ea�rҦH��"O�4⃇2M��(��NV*j5�V-��"9v��[N?Yq�7������b�&O�Te��[�ω|�B��4
���5��4_�����K�D��a�0�	_�*e�U�^�(�a{jB�h�R�I���f��5k��*��<Y���`���/�&�"<�v�>K����3�ϯc�̩a�O��y�i_?3F:�,	e�D��Ñ���d�l�CC����3DС"��V+C@ӾpN5;��/Dg�)�"OvD�рӎ"P�}cK�3Y���F� �xr�&2�@=��`ُ.���aO�� �ِ}!�$�v\&O��̅�{�2(p�O	���0���]�(`��� ��@*��]za�5�",OP�K�`�����䗼+�p����'���W�(�~��P��a�E:0��8���#	�iI�4FO�dH<IŃ�	a��3�F݈��M�3�Nɠ�EZV;���Ɗ�hⱟ0�@W'�	��)�Ul!V'u�"O�X�jĉfҨ4�TkU���]q�5@�L�8�K�M�\m��6Q>˓��� `�'UuT݂��N+��ȓQl⴫*Q3h�$$�a��$@,x�'ϨY�0,�Uh���ɦ�l�ã��9B]�W�׈6U~���W4Spq@j�%M���b�%2$���/I�HU��'l��Y�%�(�a���J%�������16��0 0�/��;k9 �P�F6q��!�G��:B�I9=jh9�`d�S��tQ�O|F6�I"a7��ӸF��� eʃH
M{�
�f�,B�	%H���1hD�*'�ƣG�c4؜�΂�0=A�,�$����uL �8DN>�O�08$���G���Wg�k��h��kҾD ��X���xb&4�I��]�C9t�*A	�hO���B�Hc^h`��4lF�B;Pa�R��U@@B��y¤�7+����̙1��݋#�?a�BX�Dش!�=}���+Y/�X���ō*�Τ�����BC�	�I�\�E���ʴ��CYD�r7z ��F������A�&PB"㎧p"Ҩ��,տ>����dW3V������ 
q^�+��P�d�H%�"�Q J��4�@�%$����Ȓ�/t|�ZA�F�M,��˃&5ʓ=l^��g��*|p�J��l���<2�%������J���y�"%X��xR��ѐi�+�	�%)�-fuy��N�i��)�� $��Z*\����=:"���+D�x�O��g���DQ�9�ڵ
��4#��D�!�����0<O��W)"h�`�F%5�b� ��'��<�A�ݙx��]����a\إׂ_А��\N�<�V�R�=<��ÈA�~�"�FK�'b����Ӽ94�F���>^��4�VP �x��&�yr.��q�x{�f��2�v`�(�S�@3�NJ6$h��!K�"~��
6P�|Z�C�����!D
�d9C�Ig���y�ڵS�D݃Wf,�P��{��;$���I�b�����L�V����&�����&����4B��l�3!ݮΦ	�D�[: P���ȓ�2{���!�%)�ąSqj�C�i���S:�E %��,9P��;$�:D��#�OX�#(U��,1��T�0�=D�h@J��G0�Y@�C�AqF��� ;D��*`��;Հh`��hY|]H�,;D�H�eV)e�\S�۔"Yp��,D�@�c��^�(1���s> P�E�'D��A`�G���o���M���&D� T�B>����8mb��ؤ�'D��J5�A7kT�CĸK�����o%D�� .@@Ku��% K'����"O60�̜�zȎ��B1d�����"O\ 0�C� 1��s�#�%Ir����"OX
E@I�e˘U"�ūk҈��"O�8A��R.h�����䁙nI�3a"ODL���L�~j�ղ��� ����"O��A뒭U�̘b��3����"O^��c�2q�B�+uA:h>䴒�"O���e��7���@�GG�m"��Y�"Oq��̾�Dp�&�Sh�ʰ"O*(� ��
R�L(�Cf܊.Ph�g"Ov��W��8��ĸd&J0!�<h��"O��
 �=�8Q�'�*�uS�"O���!��5O�����X@�"OF좒�F�e��z#MC�"�TX�1"O^%Bϓ1�4�k4��iI�=��"O!�C(�y��8�#'2U��"OP|�4L΂g�V !7*̵i.���W"O�ͣ���2�v�c�Iņ'�hk�"O��Y(Ԋ+�*M�����w��Ճ�"O���@ٷF����Ў£l���O�<��H;O&�JF�65�6����J�<�BڈZ��=)dO ���eB�<��m�0����������(�g�<a�i�,� A��6��� !
U�<�Q-�0�L���9Y�ՂAEi�<���H<^ $�dL�=�j��Veh�<	���;A�h��m�9A)�P���h�<�S�$8�@PQ��LC�r%�c�<��kH�T4��<"J`R��Wq�<i���=(�*�� �,���W[�<9��āS~�dsE�	�_X ��e�|�<�W�H���Aō	�bAJ���~�<��ꃓS�#Ɵ�݂i�qh�\�<ɔ�x����ŞN�F	�2�Y�<aţ��,���FeC"-�\͹IR�<��ct�h�p�� �n�!f��S�<1f��y�P��6W�5kaO�u�<���ȸl����LZ9����Zs�<Irψ*�4���8]2,;��K�<� �ۏ�F�b��A�����G]@�<y���XA $#'d�t���`�!ZH�<2'�Mfv3 �����b
G�<9���~&Ƭx�@ĚKe�Y!�O�|�<i׫R;{h��r��E$|E�el�r�<!6!�b�p�q�%J���8r	@j�<�4+�>B:���c/juX�kGb�<�W&6,$64�jR$��1����Z�<�aß�LtS2)P4�\����DC䉺S�Z�	�/��r�S, ~C�)v��t���H
u��p�g�Թ1�JC�Ɉ)+�!�+ݚ*z�C�k�+{t:C�	�lk� 3�6�Z0A��ØE�B��)^J ���u�Ɯ��@_;E�(B�I�oڜ��4�Q�kY�t8$� �+�C䉩?ؐ Q��?�I#*ҫ19�B�ɟoI\��g�3d��҆Aл!6pB�I�[�D�D @Z�&�{�&57�VB�	PL~���:n�Q�]�,B�	�u�Y��J�&�,LqB���C�	�>.�Q'U�Y"ɰu)¾J�C�Ƀ&蘴P��*������"T
�C�I��ek��A�S����tk
�k�����B```���6vӔLPe̌ZN�+�K҂= �[R�Ϲ!�!�� ��Q	ʝ��=i�̄5+�:Q""OX�Y���E�������g��Y��"O�Hq��Φ]L�H9��њ*���b�"O��(��ɜ@����͵(d�M 6"O2���+*��hH�ATvh�E"O���qZ('����fH2{7n%�"O�b��G1D��LhƌE/L���"O ��!�K�/�2iX�*�%x��iU"O�@E��iV�ǉT>[hU��"O6I��v�~�Е(��pO���"O(���NO��(�Th��D��"O�����K�xfSGG�q˞�!B"ODX�`��� &Y�v��q`5�'��0pn��eL�R�*E��,;���F� r�Ì�x��i�Ɩ�b�4��g�O z^w���
B�iΙ)�*}CB�L�vf9�ǉ�b�䘑2���$���d����5/�p��F85�tԠ��Q�W��]���>�QaU#d�P��I��f�x�b0u?�y�7*B�X��'�|��2O~�"�}��b�bLQ�CA�u��РCCP�'H8�)�b�N�S�O�`�X�nD1�h�{�����+�O������![�1��K v&�Zbɖ�ѲC䉃D�z�a'�#���B�.'��C�I�AX��A�˕)T��ys�IG�Y!TC�ɎY�$�Rb�_8�$Bse_8�"C䉬5�0���	�7E�L�u�҅|�B�	'%:Թ�7MF�!��H�є��B�24�:��2��A��x���,��B䉘�3��ÖTz���<YU^C䉡6��`�cM�*	������
�HC�	�y�`4JTȈ5ch�s�G}�C�	29��I�ǂT������fM
�C�I������ �:�\����*B^�C䉿GS|���L��ߊ�M(nC�8d� ���K�V�8!��ڞB�I�d����%�%t,�q�6;�C�l�D��"��U��a�䊙@y�C�ɩ~f�����7��Q�h�8\��C�I:S$|�e�s8tyz��ǘC�ɕY2�S��
�
�p����!�fC�	[�޸�,k�,��h i`4C�0m2���w�X�82�`?C�	�{�^X��낁	E�0-�7i�B�ɂP��Ŋn���I,"��B�&QP�i�O�#�T����
I'B�	�t�Xǆ��;�4lZ�oZ')C�ɤ:(���wA�Lf(�R��=@.�B�	� P���aD$,\2¦�50�B�I}���iBgҷ�!JfB�	�"���F�4m%��o@b�C�	%<|�1ua��P��гF��+�
C�Ʉ~f� ���[�d��Qa��\i�B�ə"���Qō�F��T�K�;@�B�<g<\bU���d=3�����B�I%bѤ����I�i�be���-4��B�	�z��t����b�:�I�I�i�^B�	*`t�P�S��&q�Q	C�Q,�C�ɜ	�~�xP��7i*J�A�^C䉏	"�� ���cT��U"C��"M��L����-����d��;;C�	;u{��фF0'b�����Z�C�I#�t��p�ۜ2X�X��N�5
�B��;q��u:U'�>^�NA@���:%�NB�!>�@�����@8���"nT��ZB�Ir��1�"׬_0�` �Jթya�C�)� ���PSJb�c�4��A"OT�i��l������L/ d��"O$Xc�[(2(H��K�u����"O���d .TǪճ�E!vH���"O�)[W��o���A��'
=:E�2"O|�j�&^.;��u30�e$�e�"O �NI!��r n�:E#�1{�"Oҍ�PÂ,'�B��}ȨaG"O4]9��$���#�L-���"O�\��[�D��,�/s��<��"Ol�a�K����(X�r������yBg�]D88�
J4���$-۠�yҡ͚"W��;�OB�7~�q�y�aGj��.��5���y2x�LA�H�X��T���yB&��� 4��A)��o!��	$@hЬ�Z'��;�� MV!�d�%-ΐ���X��Q��}�!� pGr� `��9n�
H1�DT�7!�S�S��Q�M�ʭJ�nF/QD!��΂Jq*�P�i�q{�!�.ZhU!�$<DBTT�pl�,J�n�bE�^.!��A5AҖ�k��N�X��-*�!��h!��K�P��q棎�V�"]: �/!���H��i�c�:h��RL�}�!�X	C �@�*^�px9�iݷ@[!�D�gcH4��FN,�%��)N!��
X��U�_*d_�h�ta�.�!�D�!�~����ͅi}�uI6� C1!��ǘ�
��f�P b}��X� ɗ/"!�2jShq�'ӓ	h��+��2I!��\'U��4�S�z��Q�τKf!��@�}C~���Ú��.�BC.��0A!�R��n�p !�?�D��f�-Q?!򄖟W��0��o'�*Pc�)��S�!򄁞?��p2�a�<�� �O�!�D�:����5E���"�S��Ww!�	%� ��H�Y�Fi�#�x�!�DیB�F�����W�X�7LCaS!�Jh���B�� Z��!���>8!�D��nŖ�3A�mb\!H�y$!�d
�7��5��#YcT~����@!�
�S� �Ж ��X�<���E�d!�4T��$3B��#��
E\/c�!��[ U����CN!L����Q6�!�dŖO� �S�ݲO⎤ �Ϋ�!�$�$l�P�����
pnh �̆�!��h�
E�����h���UIQ;t�!���{���1���g.ҙ��A�`!��̌3Z�|��B7�D���a�&G!�ȔM-�eGτRvh�<!��P�Zx� AABϮM7���P��.;!�$6_CF="�%b��P�4&!�M�Ԅ
�nJ$K���3�KV�vb!�ټbL%���[�|���*i !�Dk�V�<b��0 j���!�d�#C�T�%W	���si�$}!�׋v�h(�Q�ϼ}�����!��Z.�� ���_�᪔%��e�!�䇳0
��h�k�7y�S�bU�NS!򄞎l�y2gb
2Ba:�AQ� ���dQ1��c�lط09`��PBۻ�y�I
m�$�9�G�/����l\��yR˃6"���d�0�ցK&DK!�y
� �؃D`ٗo��� �ć�2�<XRv"O���$jIg��	��F>\��f"O�`�J�a"lx���9;ԅ4"OP��+*B�j��(��AT���"O$�f޻P64<;�G�jBXia�"O��!���8v�9���м%Anx��"O"�r/!@ X�-53F���"O�)R-�W���b޸X�bi4"O�y��9�(����^MR�A�"O:��g�y?� ���K�!J
���"O�) P,έR�D����8l�
�"O�s��ۼVR`���E/>D��"O�+����"�V���O-�nyi�"O2�D��65_�9��ӹb�Ą�U"O�X��Ė0|����A��q��"O�����(W�L�K��M6 ��Y�"O��r�勲";�q�\64�|k�"Oؙ@�hZ"W���cP�"h��E�"O����Ԃfs~e�$&\�{g~�a�"O^��b��?{�ziS兗:H��˗"O���g�^�e���p ��*��w"O.���!�<���#4,��m �ab"O�Aװ�ȑ�0ʫ[^�xe"Ob��ΐ `��Zg�B/+��p�"O��`��Fo���(�,)h�sU"OV��ŀ	R�$�c�3<XX��"O�q8G�F�7��1��G	H��"O��#r�E�1�N�A����]�d"O�0�l͎^Zh��!�ѤR۾|a�"O*!�!,�6O=������L۸m��"O<H�% � D�H��Γ�
ìhsC"Ofŉ5�M�I���m�2|�:��""Or��5�2&�m�@-B��-�"O|D*F�C9^&Q���Z�~��e"O�5Y��ɉ>�XPS�+ר@W���V"O�\����3�l��e
�$g@�i 2"O���V�®:�D�3�ȇ�i����"O�y�%G�#|ea&mN��� c"O�Yc)W�j)	E� %a�&�)�"O�(Y��?��9 u�����,��"OX!�U�2w��H��V
^fB!��1ik��̀�wJ6Mcߢ�!�D�%{�JQs�%��B�@�T"C�A�!�$U+�8��4n�q��D�O�L�!��0_CȄQ�ȘF�������%�!�D��|8 �*E��JEҒ̆��!�dM {=<Ó�>Tmn�3*��8�!򄍇,���ÂE��,��*3gUJ!��E�"`ak�h�30�x��@�0d�!���>}����دa�N���	�z!�dߴwĔ��S�w��0!B�ja!�*	~$M�#�ۡ��;�*W!�$�P(cE��eѬ5��I�6J!�$�;C�.U�5���d� !4bR�#�!����+��ř8�!؃�߃a�!�4��t�EN���|b��۬,�!��F���I���p��UqO� c�!�^w����t�\	2H��R�R t!��Z;\�� G' N^�`@�V�<;!��&nڐ��ڷy\:a�"��-!��=Ғd��G��M������?'!�$@�Su� K3�Q56hV��r�K5�!�ÏA1�ܺp��%G��u�+-7!�L�X���1!AP<R�r��G�Rg�!�� ��I@"ٜcLxA�D�?�պ�"O��3c��^4�ū"A>:�PȀ"Or�I#���T������^�)�p"O���B��9&"���ӎ:j%��"O�tVG�S,�9��/��H� "OH��f Y�j|"�Q�)I41��a"O �.�wƴzv��^���"O�p�3��7!STE��31d���"O�ͣe.&�zp�S� :�!"OF��7$��i�Ⱥ�M��B�8x�"O>��v�Bt��p��.�,�%"O��G��#/R&�S#�W�ƸX�"O8x:3#��8$�H���<a��,��"O��X�!˽#s|4��׿xR,��"O��ѡFJԑ�"C�1����G"Oz0�D�)r3�@3���X��|��"O�A��+�b���)�>5q��""O�[An߀�
��Ǜi�b�"O�}�G�[�G��|�. 9�r���"O�8Xwϑ�_<P�s�G�ʂ�
�"Op�"4iI �4u"U��v��c�"Ot�#��N�=QL�k�	��H%C&"Op�p� �,����gS�;J��#%"Ox��Tl�a��}�Q,-VӦ��"O�\���W�-B�k�>�6Ix "OH���B��R+���lP�\�2�Б"O� 3�֥^���vK� ���"OP݃ad�z�q���۫o�$��"O��a�   ��     G  �  �  �)  )5  t@  �K  �V  #b  Tm  �x  ��  p�  �  �  x�  �  ^�  �  )�  l�  ��  �  ��  ��  \�  ��  �  l�  ��  M � � p V �% z- �6 �= WD �M U �[ :b xh xj  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+��6\�
�<4�d5h��'�B�'���'	�'/�'�B�'�TP�`��!a�dYq$RB�x( �'���'\r�'5��'w�'H��'��MC%���g<���]�0�AF�'-�'��'#��'
b�'���'#~H�DJ:%�^yc�[�U쬐��'_��'���'���'��'�B�'Q
�rՀA47�(Ӵ$�=>/n���'r��'0��'Mr�'A��'%�'|��A�)M\Ȱs���a8|���'��'���'���'[�'2�'ł�
��;��=GBJ�i����'�B�'b�'���'�"�'	R�'��i1�n�?�L�'�.<�f����'��'	��'�R�'�B�'�r�'�@�`�B �~�6��ǁ�U�Y��'�B�'���'�r�'O��'2�'��`�B��WGd0��%|��<��'6��'+2�'62�'Qb�'���'8���F&/s��A(4B�1�%��'[�'��'���'�R�'�"�'U��`"c�P�P8� �Ńw�8���'���'���'(2�'$��'�2bM�%ָ0q0M0@�X&-έ,���'\��'���'���'�B6M�O>�dͳ_�`u9���4^�}r�AV8�'��Y�b>�z���瘝 C��rs��i�99�E��^� �O��oW��|��?�Q�952�b��d̔��&*�?1��MO��y�4��Dm>�������sXT�0�
L�VeF�˂�̕(�c����Uy��S�:��MB��v]G�\f�[ش0�M�<����Kw���?�m3Q�D��	��F!�X�$�Of�	`}��ʀ,r�F<O��(�_�S��kejC3&�	Ie5O��I:�?	a�;��|R�-�`�P��O�]F!: �y�,͓��� �$�զmp-1扉��Zj�{3. ��.H62uj��?aV��	�t�S�Fٴ(��A
���N4���������O\q���%9�1�\u���9����̨aSJy��[k��(ɵ��=v�ʓ���O?牟uhq�:)�J�ƥ�m8�扉�MC��i~R(d�N���,غ�$?Z~e��'ש/d>���H�	���QiT٦�'��K�?��@�V8]�|��F��mK^�SE·@%�'O�i>M��������$��7"�0������={4,�>Y�\�'r46�=G�����O\�D)���OP,s4�5ز�r���1���vdZr}��'B�|���� >-��N	(p����ÞE9���V�S0������^H���e�ړOZ�Z1�|�d�$����@�B|B�S��?���?y��|z,Of�oڑjv���I�.��6�$;ް�������x����M�J�>Y��?9�=?��+Ӭ ���p���Za�穈)�Mk�O˄����z����wYNcC꛳�p�ͥ6I de���I���I�0����
��7!%�0V�D�7	��?����?���i�H��ȟ��n�e�ɘUl���h���Z	���S�4�%����ß�(P`Ymn~"f�[���Ca�h���z�ֶ�N�ȐJI~?	N>A-O�I�O��D�O��ɖ�C"�,e3r���a��م��O���<a7�i4�aC�'���'��ӟY ��`��jx�q��߼^���z���̟��IN�)*f��_1��!�	/A��5x�[�3a�	�dd��:B��R.O��?q�j0�d͹Z�����Ǌ3�HLږ�ޅG*��$�O�$�O����<���i�+��|u��&�)��j�����������ڴ��'P���?ѢGG�e�v�����
!;�%E�?��m��5Pڴ��D��J$`�c��d�A�v8��;>I��4����y�Z� �	���I�����0�O2|�`���,��
G�)��	��d�LE����OV���Ot��T�$�����%n���: d~pٱ�T�,�*]�I���'�b>5qu�צ�MČ��L��tJf�8g�Ȼ[��͓
�d�۷��O���M>�/O���O���f�d�U$Y<�TQ�Y��<��ʟ���FyR|�t\��"�O<�D�O�Pz冁=i��M	f�1F
�h��J(�	&����Of�XBt�џ|yɵJE�dj���	6?�����.�T�#gS)��',���S��?a�/�;rڭ��#� =�@�vo'�?���?���?Q��	�O���1oni��(Ͷ`y4�{�A�O(�o�3Q�������4���y�g8wY���(G;���u�̗�y��'��'���ـ�i���"l�~�1�՟��w!�$T4,1�wU�+����!�d�<�'�?1��?����?��@�wJ��Ĉr2Y2�A�*���٦��$�����������gKCr�ZA����!ud�9"�&�����柨��Q�)�S�7H��f�Z#O3$@��BГg	2�ߦ	+.O�<Knֹ�~|R[��H$��	���X�`�<3@H�#��ş,�	؟X�����@y�NiӖAS��ODu��j̀)�h1�ţ	�Q}$qa�*�O6lZo�0�I�H�'�`ÈݾT<�pP�A�%iL�ժd!J)	ߛƛ�4�6�R e��/]�S��� �ez"fB�.���A]!;��+G9O$���O��D�O��d�O��?YȔkĘ�hǯS����R��ğ���ȟ���44^R%Χ�?���i��'�����J� $I�(t<���y"�'��I�F]0@mZd~�+�������H[,yb�O�`����ʟ�$�|R[�L�I���I�(Jde��2a�@�tÆ�;�ִ�ů[���	Qyrmr�j�� ��O��D�O�˧9�D����j�� �L~\���'.��?����S��DȜQ�,c3AͤK� ��EɁnK��Տ�5F�d�O�i]��?�$�0�Dψqԥ�+�����o�=gq��$�O:���O ���<�iz�JP!½!Fl)�w�;e��u�!��:r�' J6M;�ɶ��D�O�)0r����aQ�-l X9����O��DP��F6�&?��F�kGP�I:�dlL�|e�TK�v�bP�`,�yrV�`�I埘�	͟���⟘�O��$k��H]D��!c׳1��tk���ɫ<�����'�?	A��y�e\=2e�;�:����!�Џ9R�'�ɧ�O����R�if�� >��rEd��G�H��w ��]��DZ(MD��[�� �O���|��#���� �ʃLV��+�%N>��!A��?����?y(O��o�0w�1�	��ɨMY��(ٛyІ� �m^8cn��?�@\�X��˟�$�D(a���w5h�ħ��j��u'5?�gIJ�%���4ޘOHD��?��B���y"�&=w�萇�,�?I��?���?�����O|�SiE������/}U�e ��O0$mZ2���'��6-"�i�!��C�2!��m�ì*������f����~yB�Q������I�(��C�T%Fd�����]>�0�
E ��U'�4�'���'���'�'S������}$��.�R��T��ٴA�r�����?���'�?��j
24A������;o"�:�#����؟\�IY�)�Ӎu>�9��A$x�A(q�8xFE�2��3G4��'��E,ݟ4�@�|R\����F
	Ab�iTI�AF-X��]ݟ���ğ���֟�Lyr�u�vɨҮ�O���¦�P��L��&y�ҙ�S��OTdm\��h[�IΟ��	�����D�~�+2�M�%U�T	���.SR�\�+���RE���>��*ix����Ҝ]}�<S�%�.F�F��t���P�I��p��K�'s:h=�7�7y���.[-<����?��Hƛ� ɔC��I�M�L>)�BD�C�eK��U?h?�xRa�T��?Q)O6@s�r���+(��C�:]�����Vz6*XZU!��<F���@��䓾���O����O���"cfm �N\v'�𑑥Iw�b��O�˓;Y��!ޢ�R�'W�T>)�W�3e�Ĺ;��<; xH��� ?�PZ������ '��'Q���0��^���3HĿ9���eJ�;�f��˝j~�O(��	9Ua�'c��f�L(s�`���K>��V�'w�'���O��I��M;�o�`S6�a1��<k�.$�����[��u���?	��i�O���'�OP�^�>�����( Y�P(�!W^��'�LS`�i����~m�S�O\�:����E�E,� �f!=JCv	����O��$�O����O2��|R��_&&n���+�(oS��Sq�I
H���eC2w\��'!2���'�j7=�f��t"D!Ml�=c�����%s�a�O�b>�2���=�mDT�uM�w�ڑ���[�zA�1Ox]#@�\.�?�n:���<���?����%�=p�
A�K! )+Pf��?����?i����$A¦�Q2��@��ҟ����8�J�QQ�I�JD��(�"AK�g������h�eW���IŹ%�
��1IS��sK�$	��0�M�&��DKw?���:�I��#�;z���` * ��r��?y���?����h����7(�<`�2
�� (zѲ&�IJ�d�Q�$E�D�ɔ�M#��w'��C�*��]K7�̢u�X�+�'�B�'��)��]F�v���]�u�\��3)( 2�ƹd�%q&�[�5��Q���|rU�,��ϟ��	ğ$�	ßD@�Λ� Y�� E�3VDz����Qy"q�Q���O��$�O^����ɫ�����@�gO�ѡ4׽. f��'G��'�ɧ�OM:e8v�^ M��tX��0��pß�k%����X����q�D?��<q&J�u�N�+�K�"z��=��G��?���?���?�'��DQ�Y3�����q is"��E lA�!D�| 4������C}B�'YB�'��, A	M�@���"Ք���(����f���g��,%�4�	��R�e��,��%���Un��LI�6O,���Ot�D�Oz���O��?�Q�F�	�J����#�v�e@�ڟ�������4�&��'�?��i��'b��y���}����װ	����y��'�	�^�t�n�c~2���z]b�e�d3�U+_�)���Xh�~I�I�dz�'���ޟ���ȟ|��N:0{@BȌ-��� +�=7�M���x�'a�6m� �$�Ol���|"V&N�[�n��d*�4o��5KV~���>��?�M>�OxJ�(�*�����O/W�:B���!\��i����|�a`��l$��Aa��s���
,�ld�%%�͟��IП����b>��'M6��7S������Q�0EWS��\9uͽ<1`�i��O�Q�'�� �I���8�͔28f�Yg��G�b�'�҄��i��iݱ9��T�?�Y�W�� r�����=n2�q�E��rޞP(t7Ojʓ�?����?)��?Y����iC�^�����,�{FrEr�ߒuBtm��U�	����G���H����`&�=CDV(m��g��?����Ş��Y��4�yB�A�>#���Wd�)�j����T�yb��|U�a�	�xD�'Q�Iџl�IU���Z�$ɌD��/� S�,�	�����ǟ�'��7M�BG8��O�d�Wtڀ ��%<ޝ��lY�h( ���O�$�O֓O�Hsg�̡��E12	�S�,�瑟�ba:0��LXo!擿0��oAП|P�B�/�t "�iP>�l���ß������	PE���'����f'�#k� ���c�HȠ%�'M
7͚
1^~���O�oS�Ӽ3��$��h0�K[҉�����<I���?���J5�u{�4���Ӗn"�d���S��%�ִdI�8��,��o�`��,��<ͧ�?q��?	��?م��� Ƃ����g��5L@5��D���Ґ���	ӟ�����%�@����qc|�0N
6|��ǟ�	y�)�*�<  +�/�(Њe����Pyq�K����ٗ'dN�Cń���"��|�T�x�F�J�&��a�2,б���C �U䟔��ϟ �I���S@y"�b��)�J�O�d9$e^�z@�yzV^({[e��7O�o�w�|��	ğ��'sd�BC� �.�yF&,d����і8��v�����R��TH y����mۄn̻-l�;��_?8
���bp������Iğ0�������2K��ݢ0A���/q�KZ#�i�	˟�	5�Mk@��|j��9ț��|RG\�(	}i�< �����l�Vq�'L���4�����V����&J:mB���P��0�L�C�eԊa&(��v�'�
'������'v��'�R�ӣ�=��5��Q�q d�'��\��:�4I���I/O����|2ワ$.J0���T��j� ^~��>i������F��|���|�2�I��V�h��@uҦ���ƾ<�'���������zhP6o�=y�R��#'�2ߤX���?1���?��S�'����H$�O�2��]!�R��1p̕���D�	՟�s�4��'X��?��@�UV�����#V���Ղ�?I�e�R��4����T��K���/O�m)q�͏�hJw �k8�T�#9O�ʓ�?���?����?�����O>�\�8C�� CU$��C��m��\f
h�	ş��	]�Sşd0�����,V�̼��V)������Ζ��?�����Ş)�"�ڴ�y����Y�I�r�c�ݣ��]
�y �.�$U�I?��'���퟼�I�pDXxPFg�(Į��I_3�Q��֟��Iџ|�'a�7-�ր��O0��ŰX�� "&G��P�،W�-&�\�쨭O �D�OܒO=ke�0fpQ�Ѩ��e�ЪR���ԧQ4f�Vl,��'`�l���<����.bv��I��$:N&����R��<��۟���̟�G���'f���ҍW�:���E0���C��'�p7MW�|;���O:�oZm�Ӽs@�Y$I��;c#ڿ2XrxɇD�<����?i�����4����^�%��O���AVE,��*����![<(�ӛ|�P��ٟ���ϟ�I��+�'�L�L��%x�=��b�jy�f��$m�OZ�d�O���\��ތt�v��6`H�-��D�%�4cW��'���)�>�zDsW`�ek�|8#��p�l�i5�I�uV˓d^�����O�AO>�)Ox�xQ��)x�z)Kg@b8�}9GC�O����OZ�$�O�I�<��i�~q���'
d��O�_�d�8V#ʠq0���'�6�<��9����O"�$�Oά3�C �L$؃F����3��@q�6� ?qc��9�D��V��߭���&RZ�C�%ߟB�|��4�u�h�I��I����I����#BǎV����@�˽R��1$ߪ�?A��?���ikD	S�O�r�j�>�O��w&S�>W�aa�Ɔ(^�rD) ���O^�4��a��o���el���B]&/�T�H�/�8�:�0ӥ\"3/��	X�	Xy�'K��'Z�'K�q�Q!t+�8+PJt��Q :#b�'��ɪ�M�ׂ�8��d�O&�'���)U_���	��X@��'�2��?��ʟu����n4����	#X��(��Q�+{�}Hq��* ��|�ׁ�O`�HJ>�t�K�{��ːg������?a���?���?�|2+OR-mZ��`!8��#Dt�Ŧ5UhdQ2*�4��
�M��ͪ>��NR⊙�'�<��3Ӟ�P`����?I�b�=�Ms�O���nK���L?�HB"B�'�^�2�V=aȌ�"�l��'���'{�'&��'�哜3~�9��!�8��aB�I�D�� Y�4S�����?������<Q���yW�^�
3�%� �N�k@���w2��)A)��7M��ɥ���!	���-Y	/Ű���#{����3
�[_�	sy��'E�FO�,+��6�ψ]��Q6�N�8>"�'�R�'Q�	��M�W��.�?���?af�W'�֬�4& �A|�i����'#���?�����za6E��H@&ڊ	ѦD0x($�'+��Ԅ�;�x���D�џP�R�',5�TI��@��U��Ȯ0������'���'B�'�>��$XL�RoРʀY�F,]+]�@�	��M��K0�?q�x4���4�x�P��C�R��6���W���>O|�$�<Q"��Mc�O(����Й�z�� tqh�
� }��#b웋�l�9um>�$�<���?Y���?���?)2�	/͈	��Ƙ1O��7`���d���]�1��}yR�'b�OfR�ƎMAdTS�"֩:�Z�"��0H~j��?����DC�xY�%�%�C�8�6���;�(�94B�P:��$�@8���'	B�%�4�'-�
ƨ��jƁ!돴y�P��'���'�����T\���4u��LB��`=��`�#�h T)��)=��̓}<����O}��'22�'��yB�ה"E�Tї!͡�����������R2�¶w��!�I������@��b����+��<.n<�R3O����Ol�D�O~���ON�?3'��8�0���7.�f:�N��I����۴b?\m̧�?)0�i��'2Jt2A��id�̸ �Z7ze.a��|�'%�O�n�ʇ�i�Ɍ�L �dL�{>�b C�I��9�u��L��0��<�'�?	��?1 g6\&�Mq�mJN�����_��?I����DĦŠ�![cy��'W�*xr�A�Ⴡ.R��[`�%IPX� �	ş���d�)rE'���('	(�9c-VtFX�"��L�� +O�	8�?A#%������A��	�dL���4H�d�Od��O���)�<�d�ixV�f�"jA�%�K�F��-	Í�l"��'��6�:������O���KՎ
X�P!JU�rj��:��OP���<|��7�/?��'X�X)��wj*˓)%`SF�]�� po�	�M����O��d�OJ�D�O����|�W��o^����1�"�ض��b���lŞ|�b�'�b��t�' �6=��\���G�z���6 �h<�(���O|�b>%�DEئy�_���9`f�l(�#����0�f�0��&�O��J>�(O����O�@A/ j��,I��/*��д�Ot���OX���<��i���z��'���'��q�@F4��x*��� 
�,!��$�S}�'��|b��\�XT�g 
h��LJ�`ĉ���@.�b���oш\1�t����\����%l� ���Y�N�XDГ��70�����O���O��:���b��	V\Y�H��P�(����?)P�'�^����?1��i�O�.�6���&g��p�DJ9���Or�D�O�]�mӨ�4� 1Bn����l�v&Q��E�B�����%H�����4�����OH���O��D�c�6�yC&51��E[��]!P.˓	���g?�"�'����'+H�jү��t���5'رz� �ʹ>����?�K>�|�T)�
{�Z1��+Z53������n4p���Tf~���j��I�L�'�剆@�6)¥��;��iF���:pJ!���L�	̟��i>y�'
�7-��8�<������������"�/�`0�$�a�?QbX���I����I'`°!rCI�,�SU/ʍC�Px[@#�¦��'5�B�HX�?�E����w����gF��\���ȃ�(�H�`�'x��'���'���'��1�.\%���k�����&9�?���?���i&�Y+�O��Kw�$�OfP#ʘ+]�fHX�lĎk�Z�hcm7�d�O��ԟ�@"u�i���� ^D]kg�؀t�@�sRl��=Tl2$F7vR��~�	vy�Ox��'���Աٖ�jb*�F�ԑ��2�'���"�M�M��?���?�-���3�N)��y ���u iS矟x�O`���O�O�SKz"��Ҡ�5���ԁ�0T�M��"%�:��*?ͧJ����E�\��h�\餽�@X����s��?����?y�Ş��$��?�(boJ��Bԑ$�Ӭ���h��� }�F�d�_}�'�,�A���e�]� M�[�����T��r�mզ��'�TQ��?��^�XȤIK���H4ꂬQ!�h1�w���'��']r�'p2�'k�S0qh��\ vl����Ss_��޴"yV�+���?����O��7=�b�s����|Ԭ�[& W�h�J4Ѧ+�OX�b>%�g��覽�?��02#HI�
�K�$ޡ0�θΓ3�����@�O�BI>�)OR�$�O@��pF-]&9ۇOۭq�0s�/�OJ�D�O����<���i�v�ɗ�'Y��'����lϯ3r������1���"���HV}��'��O��	���G<��C6e�H6�h���@��oJ;d������k��8e������
�E
c�at��yW�La��U�h�	ӟp��ݟ�G�T�'���'��6EhaCu��:�D���'H7�O�J���D�Oؕm�P�Ӽ��Dޏ|�B�ʠ\'*Z��O�<����?���HΙ��4��DJ�~,T�{�'|?�A���04p����bTe9��<�'�?Y���?)���?���/'�����-UW����������,A`r�'B2�)6$��T��L�$O��r�.F�BA�h�'���'5ɧ�O8H�sՃ#�U25���(�v����(ؙ�O��V���?�3E �d�<9%с>�"�j�)8L!; kG�?���?���?�'��d̦)[f�C��h�aE��j9b4c�1u��E�o�Ɵ�ش��'�6��?����?Ƀ�[�>����YSM�ҊZ>�JA(�4���K+B�$�����O}��۸V�l�R
ռ5Xt�E&���y��'���'U��'�b���$L� q牕^ ���ҁ.�,�d�O@�ĕꦝ�a}>I���MSM>�PG�&o�����L��Ji-k삵�䓪?i��|ƥ�0�M[�O6ԑ�� �U�憎i �'���b�;`���?�6 "�D�<ͧ�?����?91(
?.qM�w��<?ऺAa�&�?�����Φ��ǡ�Ey"�'4� ��A��%�\Y�f�)��[I����8�	`�)r�"*J�~�HX�VeA�f+��ڰO9h�����@�џ��|�e�+A�H�vg� �a�H1NyR�'Tb�'��^����4z��\K�eR#He�<�4�3I����/���?���6������l}��'��-sq�Ƥ?[�h3fCR;VC�!fU�������'�h��e��?�c�P�ہk�5|��t;wA���M/t�P�'�"�'�R�'�b�'���w��|����	N��h��TX޴QJyj��?�����?	D��yGEK!;*r�h���&JZ�B#)ŀx���'ɧ�O;Hӱi��I,eABuh�%�"�Z�z��JL��T�&[|< �'�'=�	ǟ�	�ı��k�,:$X�P`
u��	ٟT��ß��'^,6��-ʓ�?a0"L S�<"&e�	-%���E�H���'@���?!���_c���'cת����j�
�@��Pi'b�5P�&Un��'`�F����b+S�6�"�oJ>��7��x�	矈�	�hG�t�'¤�	B��W� ����(h����'?�7�\�<���Or@o�O�Ӽ�e�L5^�0�Ǥ� &�� I�N��<���?q�HL�� �4���I>@z�3�Of�䒁�I�PJ��s�P+���Q��|"T�������	۟x�	��4�&Β.r	j����%_�:�Aw	�Py��j��Bǁ�O��$�O@�?1UF�*m�D��kJ�v7�:#g.��D�O�7���6��1���<DC%(���n�v�d��O��<'���'L��� &,��"^�~�8�3$�'j��'o�����W�T�޴x5Jz�� �0�Q·'a��駡M�10P���N⛦��x}��'���'+8#�ȅN0���BG!o��K���������Q�,�����	����:��e������g'��ȕ6O���O6���O��d�O��?�j@d�I�H�Z�v�� �l����IٴBz��'�?I�i�'8����B���x{wa����@ɢ�|r�'��O�:�葶i��I=hR��=��qs`�ޜ�L��ȥ���2���<���?1��?��&�O���y@*<A�l�'(P��?�������f`���������O��$��=*n<�e
wzD��O���'x��'cɧ�	���Ł��%3�F�U�L'(�2XA ���Xb#���S�(bF�H���
�����J�jx�bS���)�I��(�	П��)�Gy�aӼ�8�#�'v�n-a&!�A��9����#>���OlTm�t��fW����4k@CőXau���˲"�mh��M�<�I�r�.tm�t~�$VF��4�J�)�	b�0��C�Z|&���T5LR�d�<����?Y���?���?�-��y��KR�zq��y���;Z�hT�tm�ܦ��BNԟ@�IΟp'?M�ɳ�Mϻ`V̀p��P�O�!�"�Ҏcf�
��?�L>�|��F�M۝'�0U* G�CF|+'�^�'�A�'r�1%��{"�|rU�L�I�Q$fUh��Ŋt�W�'f��CGZٟ���$�	wy��V���k�<I�[0��F�@���*V���a ���>����?�J>i2��8[e>���;��q��~f�5w��aǓ��O���	uL�f�8Ĭy�
 	i)�Xyf�ܩr/�'���'A���۟�@���n�D���\5�=0���͟`�ߴ@�U���?	��i�O��(j��u�܏J��H�A w��O��$�O��)��s�0�4��t�ǥ?�Aq��-=�5�� u��N�Ay��'Zr�'+b�'RFʄ(���2��.��xP���@*�ɐ�M�u/�:�?q���?�K~z�2W���ԅ1x�l!�֜>�z�TU���	���%�b>=�`K���2,[�2���9��,7���Ka�)?�s�Z\oB��������D@&%�P�X��eDD 2r�٥ �<�$�O����O�4�l������f �I�����Bvʟ"\xF��H�B�x�J㟼:�O����O8�č-"h�����-�4��O$rr����u���=}0��s���4�>���~b$����n�:P�T�C0pOt�I�����˟��	؟8�	i��)\S勑�wP�F�-0��j��?!�vH�f�H����'6�<��'\ ��q� 0P$���1O��D�OX���}r�6����< N�2���&
��ݛF晫�,�!�G^/BN҉�o�Iny��'���'���T�;�T@փ�?7�6UIa�$:���'�	�M;⍄�?���?�+� ���+ۮ#�� i� s�hy����R�O���O��O���	ȚᚂN�1'� s��^�6 ����uS���b+?�'���Ė��`��� ��,G.pI��̺*�b!����?a��?a�S�'��d_�)rAmE�~�i�D.J�-�p\kC��T�Tt�'�6�;�	�����O�1@��F�\j]�`dƷ7&��QU.�On�d��
4Z7m&?��qBU���2&�L9dp�)�8��5���>��ϓ���O��D�O��D�O8��|�P 1m��E�.WB����N�9)�& �5m��'�R������;A�Tĩd>R٢��
E�9�I���&�b>e#1m
�u�S�? �iso�>*�l����>�Q��;O���G��?��<�$�<�O����CND|k#��n�����o����162�'��O�/�.�Ir�T�d�`S����s��O�|�'Cr�'f�'�p�1�6@RL`��� =|�5R�O����Z?Ŏ\;�C9�Iؿ�?i�c�O��˕
7�l;Tk�4�$�5"OH|��n:r7H��
²&`}	U	�O�o�s�VU���|�ڴ���y�j��o h�5N:���cf)I�y��'SB�'�F��i�I�5��	B�ԟLA'��gbP)��P�,��QJ��=��<q���>+>��Y�m�4y֌�KC�ɽ�M��O��?����?!���VU��D&V�q2�A�D��l��?�����ŞC��e�Qf�rY$K$�V0#����M��Z���,X$-��<��<�hC?� Tc�`��+�l�Fd�~��IٴW�$�3��7#�q2f�K�
!^T���
{~D�c�D���d�Q}R�'6��'�@�b�j�q�v��Ӊ�=�,��n,�v���� F�2��T@�j�S��M2�K��T��k��
�X;���Ro�|��I�?;���Ճ��O�xh0�	2,����ߟ��I��M��W\���s�@�Of�8s� �D�1w֕s����)&��O �4��kPCh�D�"Na�G�)ZD�kD��F�%2g�My��	q�	fyR�dl20���٩P�����͡C��XYݴi��q���?����򉎏!<|�[f�M�@��	�P�	����O(��7��?���/�3��+����]��L;h��y5BԦa (O�)Y��~Ҕ|��N�`i�m�t��1y���:��Np��'<��'���\����4	
X����X.���e�<��Ч�¼�?���{\�����W}��'{������'=���(�$8���ѷ�'���F''�V��4��M�6��)�<ya���\��dE��sw��g��<�-O��d�O���O
�D�O�˧(?t�:!�(} �S`M�G|[3�i�$t
��'d2�'T�O`B'`��.ͣ0:����\إ�S��2��$�OT�O1�f���ad�x�ɴMd����&yC�Q���X!��	*M/�|�w�O��O���?Y�6�څpLM�^0�IC�`ߴ$X�Y��?���?a+O�o�8hӦU��۟��*[L~�-�����aVcë	[�?�Q�$��ʟ�%�X���W�Qk��[4�W)L��P�P�/?�h�j��y�ݴ5�O�0-���?��o۬ 1 �k"��+O�@��1nW��?Y��?����?���i�O�a�%��״�xf)�>?3�(�$"�OP\m�2g�.���ܟx��4���yg
ٵ��9�#A�?T�K4mO)�y�'���'��ً�i0�	U��ڟ^�YeJ
�Rs�@Ȱ�9T�>����,�d�<9���?���?���?y4�֌A�E���P�~�@0sM�����٦u+���꟔����%?��ɹ"*];3 �^�|�J��آ2� p8�O��D�O�O1��ax����v�!��_Ҩ�ha��	f��7��\yR%D[�L ������8q�sV�śp�����ڊRɠ��O�D�O��4�8�4��o�'d���3�f�$��*�h|J����]�b$fӎ����O�$�O��d_�H����jM�'�ܑ��j�8.������j�x�y�8�z���?�$?��ݹZ����w$W4���'X d�蟈�	�8������	@���]Q� \jD`��1e�H���?������������'C 6-'� �Mk���j3Y��=0��R�A��O"���O��ܴ$��6�:?	@d�<B�IB�Y8L��ݨ� hѣ���$���'82�'��'0h)��گY9�a��/�D!(��'��P�lٴUb�����?�����$�fmQ!)YB�����f�4a@�����d�O��$6��?i:PI�8e����#�!�fH���Ŧ�d(�����1r.O��|~�&�4"��Y��1�O�+�2x�ѩ#��Bٴ7��ܺE��o2���`�
5���;#��-�?���f�6��C}r�'SLeK�A��|�-I��	���"2�'���{@�v��|�d�fO���<�G-� .p�`�M� ���0F�<	*O�����`�QH4�N�p� FE��S~�o�/I������|�	c��t$��w� %��E�O��L�6n� elݹ��'��|�����ʛ&2Or$q#�
W���I���(S`�[�2Oꨠ���?�2%?���<�/O�Tg@�� \l����x��B��'�7�Ğv���$�O���5:ة�p�O�p���r@���qY��<��OX���O��O�0*��H�,�d��Z�T�&u�s����/�,x�l���R��Iџh�3l�=*�H��^+�|A07$$D�Soԋd�jѓf	�vBE�E�p(�4~2�()��?��i�O�n�1�(p�A�Y�$���OOl^��O���O�(9Dw�J�H��s��?��d΀�.������t��m
BGn�y��'���'�"�'��9�xsF�òE�޸�� )w�3�MCcaԭ�?����?�O~���W�4zr-љy*~��V��y���\���	ğ$$�b>e#�L0� �!��B�l{����Js�����
2K8�I��>9�S�'�p�$�4�'��e)C�߼:}�����I�B��5�'jb�'i����TU�LQ�4!A"њ��f��r��'�ZHI$eL�6��b��L˛��DLr}��'��'+��ڱ�WQ�D13L�1���J��6�����JT�ޏ0��)#�	��T�fH�h�KF��e�E�4Ov���OT���O,���O��?�b�#��n��@�X
2��0)��� ���H@�4"%@�O8.6m"���"lnX�x���]����%��_o:�O��$�O�ɗ�	�7�5?���B�2�G)��C�ҵB�B��I �T���8'�D�'��'W��'�29�BEӿX��! k̶
֦����'�^���۴*yj]�(O|���|����7o�p�˷i�Żc@�p~RE�>���?aK>�O����&ݳ/B���c+w�0Ex�K�_�^i�úi����|"�ʻ��$�������5p�R#�Pw¡�Vݟ��	����Iڟb>ŕ'
06-��*����$Ȱ`�dr#K��F��r���O������?Y�Y���FiP=�#BZ-x:}(��T�$�r��Iß�bY���'���*�O
)O��2�	�a�6Ts��w��hv9O���?���?���?����	K�rm�����q��L�^��s$&k����O�O����O�����D����q8�e ��ԥ��e��n���IޟL&�b>��II¦�͓!�45���!%Fh��D�H`1ϓAX�r$�O�$XH>�*O�I�O�9갌�Jr��TI�+��+A��O�$�O�ı<��i(t��'���'�&{�EQ�n�6���fu8f�_l}��'oR�|")� zW�X҅ɍ=^ ��ߤ��D�zd�SU/U�L�1�@�{��I�&�d� �Ę�O��c�ö�}	��D�Ot���O�D'�'�?�4nW�j�L�5��� AX7�S��?)g�il��R��	ߴ���ygj�:�:�ze��,n��[� �y��'��ɯx�
|lX~�I
���S�:��-Q�*�Rb����A�������|�Q��������ϟ �	� ��fR1g$l���tjNd��Kuy.k�@t�g��O����O����D�3�xdi���Q*j�2H�'����s���p�
�Dn�D��?k� �!N�e�0ʓ*��!p#��O���J>A+O�E�� �(��|�ǛoJ��L�O����O���O�	�<9&�i(��PV�'J�,s��_=؞᳣
U0y��X��'��7M:����D�O��MTbY�畧t�M(W�R�J��@y'ʇ��M[�O(����R�)4������,[?�\����0���3O��d�O�d�O*�d�OZ�?U3�Ϛwm��Y�LK�M;(���D�����ݟ�ݴU����'�?9��i�'��������҂�!z/:���y��'��I�"_D�l�P~R �YM�\ �9�,QR��r����ğ���|rT�(�Iԟ ��؟���	S��e��L=�ي���� �	ay¨g�p�#P��O���O|�'oo�A��OBK�f�%N��:K��'m���?�ʟՁ&�ΓNS����B�� ��QsBܤ:�z;���|"S�O����H���x����V�`�3H�"�D��5�%��H���!�l�@C��Wwf�)��B*��z�M���К���?;�j�Jg�7ze�jF�q�d�ٓ'HM�l���*�HO���ιm5�ș�$�%B�8�2>�l(�!��ȷ(�*y�(��ɋ�B85��S5)H���P��!}����'�!�ƅ2�#�99����(�'BP(�r�H��r�(�bWΓ�C�
��ET#a�\)���)x��Tʋ�n
���u��B��}K4(�w��%;�n�	#3<$���#����3��4*���'�����&�d����x��� L��,P�kR9���bb�Μ]��&�h�	ן\��By�bh��	w>�P�ř�I �O	�K�^l�-uӾʓ�?M>��?����~�K��&�̳��ŀsJ2�����d�Oj���O2ʓ9y��XG^?u�ɝ&�P�����b5�zGD+/5T����$�P����\��LaܓtlpZ�ᇔi� �LF�2�lП��I@y�ꇞ6�>맂?)��b�	[=��� 'C���`dH9�'7B�'^Z�Z��$�?u��
��@g�H怟
jż�zU�`�X�_�rU�ѵit��'f��O������Q�a��s��� �c��9��������X����OW�Y��FN4��	�4_��} �i&��[��s�r�D�O�韄p�'���);��W��":2.ܐ��Y,�\���4^��y�����O�k��F64:��8��τ`0� X즵�I՟<͓� ��O�ʓ�?Y�'p���f�1]L��q�GYA�$�ܴ��u�`L>���?���f�P��}COX�gu���̦I���)ЯO���?II>�1 �`q��cW� aXcCO��bh�'<�����' �	���	����'0�y��cLT�Ȕq@`C�<���r� U���꓀�$�O��O���O��P����T�~9����~~�թ��WTᲒO��$�O��ķ<����*2�L!h���hC�R���:��R�\͛V]���	a�	۟���;~�v����K0R�@&ղB�����b �<��O���O��Ĺ<Y�#I�����*˯r$�5�#�QG�%2���M���䓆?��pD�>�U`b@�1e�&R��	������1�Iʟȗ'�@"0a'�i�O����lࣵ�ԑx���f��O(�@Pu�x�]������$?�i�� ֡��g�8Fg��aD.�
DHmCu�i��.�V\:�4Z����8����DF�i�xպCj^'��L(��ԑ%n�&]�4���qK|jJ~nځ/����OёZ��1�	�	6�GQ�$nΟt��Ɵ��S,���|z�O?2�n|��R�)0'M�jۛv�'�2�'�ɧ�9O���˭7�,�[�m@���T�l�g���m���	џl:������|����~2��:?�F0 gD�2~P|Q��V�M3������3?����~rm>,��e���=tG�`�tR��M���0mdx�/O�e�O �O�aa�mʹM�(��!,�n�HP��+�D≑m"�b����]y�'ӄlHƅ�gvh���Ԉ'�
���d]���	C���?i�'Q����#�=�����  �H�2u�ݴiʊ��<9������O@0���?�j��i|�mz�DH1 5/m����'y���Oʓ;m�HnZ�7�4��'�σ2�~��3�@h1H��?���?�)O�KA�O��5E+a�5\��p�EE�E���h��p�^�D1��<�'�?)L?��p��G���X��
�t�!&hm�`���O���&ex����'��\cβh���f�E
� (a(��M<�,O����O���������������X�Ļ� �>���4������?!��?��'���T%	���b̚8Rpx"eS��i R\�|8��$�S�S=^u
qY���+B~x�Q���NI7�X=*�lZҟ��	ҟ��s�O�N�C�ne�&�J�@x�a��Jw���m������\%���<��Ytq��Y�6��q
�����s�i��'!�.68��O��f�OT��T)L`�, �)?}Pտi)��|b��~��?���?��%���AC���Q0_/����'�7+�d�i>	��v�B#��Ӄ��<�R�ӂ�G� ��-�O<�����?q/O���G����!lS#|�B��c� ?-$�S��<���?����'��䖨S4�+DF	1cE85�Bɚ+����U��$�O���O�t,གG8�ڐA���d�2���C�8X�Υ��V�$�����&� ���4�'#^�9u�Ī>��#&G�c�u��j*�D�O^��?Ѣ�[����O����Q.2���u$@�xĤ�bA�Ϧ%�?����ğ3�'�A�r�X6U�dDP! �N�H�9�4�?�,O&�d��$ɢʧ�?������ph�lxvA��&����}�>�'�H�	wy��O��R]�t�� ub`��GI;\����H��&����������?��u���*6�<�� )W�K;������MS���dR;Y��Af�G�9�Pt{u	Y�i�*��'�iz|l�ky���D�O��D� '��2CD=:�l¬]M �
��Ik��K�4�?���?�I>��y�'���F�*�L ��)�-,>��
�d����O>���I@�$�����K��0q��Q@����%�4��ulZџ8&�먟��O����O�0)����Kp�)X.B&{9yǬB��9�	YM���L<�'�?�O>i�E�s"��	��ѫX����bs��'�BW����П�I]ybE��M�$H2֦Y��T�Pw(�<K�>1�� "���OT��!��<�;f�2%�C�/4�����M�P��8nZ�$�'W�'��\����/�����%P�1j\�QA�)?����؜�M�(O��$�<���?1�~�$��
c���c�-K�Hv�؂{IZ}��V���I����I]y���!ꧾ?��#%Yg"����b�����CK�]}�6�'m�Iޟ�����\�хg�ĕ'���1ƕ-Pu�A�T�Q�hR�Y7aӄ��O��m!��X�Z?1�Iڟ���Wy�)�L	:Ĕ��$��$z�O����O"��άw`�IYy�؟T�ӡDțm��q�j]�F|�Ʒi;�	��h���4�?���?��'	�i�]؇H�*������Q�8�5Lp����Ov��B8O�	��y"�i��|' �t�Ӧ^����E@f��Ac1�6��O����O@�)�]}�U�;Q�B	�� ��'�����G��Mc����<�H>1����'oL\#�Kюwq���Ƌ2!R���b�<�$�O��DT)=��\�'q����|��e(�kS=mLl�� ��sO,XlZ��d�'�$�����O��d�O�e���K�B����F ��f�`�æq�ɡP�
@�O���?(O���Ɗ
wjF�<\����X�<p{�Y���f�Ė'�b�'Y�O�f�;Ajԙo���.E�Tƨ�����*\@����O�ʓ�?9���?�FJ߄�bX� ℗�| ��f~�]��?���?!���?�(OT���D�|"t,�8"O�x�r�'�*H�F����	�'IbP��IП �I�Nƈ�	�qFE�!���'J4�b �-��1�O����O0���<�f��2R�S��@�1��
�yनܷ3/F��2ŉ�M�����D�OF���Ox��W:OB���Y`,,e$E�G��1�J2��h�:���O�ʓYmH(A�V?��	����5�����'˾iΈ�HQfF�Z�ڮO����Oh�X0)��D�|Z�����l�74��=C�V�caH�s��J��M�.Oȸ�QbB�������8�	�?�s�O��7���@D��A��L�ui���'RI
<�yҞ|��� ^� ���i�r��_�V����7-�O����O��i�}U����J���ӄ��:� ℎ��MSсD�<�I>q��4�'Nn� R��s N2n=��Y8i��i�iNB�'T"��1U����d�O��	&lz����ǵ"�E�t6�-��F�W&�?�����p��}���ᑫ�
	I2���ao�ҟ�j`�[��ē�?�������/�T�pc(OL�qrƊ�}}"o��yrX�(�	�%?��V*Ɣ|8���8&窰�W@όl�`�BH<I��?�M>A���?i���$����	ĳ.>Ȣ%ԫ)�V�H����$�O����O(�=޹�u=��$h FO�e�D� ��K���xb�'
�'r�'��`��'	���R�U?6�z��¨+T.QP�#�>���?�����Xȸ&>�r%/�?�PiCM���֢���M������?��'x�j�{RB�.:�P��q^�F"��VF���M��?.OviY3F�]��ٟ���*:�:�����c���@�L�c�̛I<���?Q���?	M>��OER�0(�s+V�!�%,Ġ��4��d��/Hh%mz�Os2�OL����2!�][�*Xۀ̎1�Fdo�����	4$��	I�	Eܧo�����/^�{K��Rԋ�?�o�n���pٴ�?)���?A��j-�O��J�%�	�8q�)WnX�3R ����"@��$� ����3'�ё��'@,,T�D�0F�L�3�i��'�B��\� O<���O>�	$� Ab6 �2M$��)֭��6M7��G6aF��%>!��ڟL�I.H�z��0-�����S�{���Rڴ�?��d� D[�O��$3���°*�Né4ʽ�]�m�:���R��s$��h�'���'��O`�'C�@�޴�O�G���p��|�rc����v�џ��ɸ4,R����oA��V��)�,��1�����'^"�'��V�������4���N�C��1��DX���d�OJ� �D�OH��9|���ʍcų�%��tmb����])N�LH�'?��'�rR�D��M��ħG�h��0e�1KS,]� f�i[W���	�h��TF
�o��X50Q��I�f߉0|��%��u|���'kV���"��'�?a�'8Q�\25)��@1��:�Ė�l��!&���	ʟ�ASg~�&����
�8Eے�>Qv� �̀�`0mZgyr�� 0� 6�S���'/�de ?���R `������"��,��IΦY�	�����"Z����OIX\h�OJy�����m{�`��4P�JM��i��'�O/�O2�$B�|c�-,L�H9�̲m��dlZ+���?���$�'�P3��01hr��Ɨ'uV�`� S�'i2�'�l%h`g �4�8�'��=8��:px�hA��<���ߴ��'���f��O.���oml�.�tdH��c]"yt\o���J`����|���A����`hY��\#6�X/b4�'rY� ��ȟ���ey2@S�H����b�ԗuX����X�lk:`��#-���O���Oʓ�?Y�U�%����8S�`��e�V��t3 �[d��?����?9-O�p��]�|:� ˟dp����ř<<l�M�U��A�'�b]�D�	����	.Uc�����b��8���g�63� ��'���'�Q��R%���)�O��Z���)>�6Tb�M�t�Q;1h�Ц��	Byr�'z��'H��'�哱SrR�	�˜9��	3r���c;�| �4�?9����5�:��O���'E�T&�/S����#C�	"ՅA
zwl��?��?Q ��<�+Oj���?q�p�C{ݬ	�N3<�
$+z��ʓ#;
�f�i���'�r�O:��Ӻ��� ux1����>2�{�ئ�I{tw������"��Gv�� �,m\��a��H��6�4�f�lڟ����Ӳ����<q�$����f��:I�t���ȡP�O��y�'�F���?y�	� ]�����Ɏ�5ڲ�3�'E�'ӛ��'?��'v���r�>�)O.�����H0#��{���6��$�8r��x�v�$�O���˴P�?���ҟ����d�B ��-��O��	�&&�Y�|�ߴ�?d�5=���Ny2�'i�Ο�����8׆Ӽ1��	1�$d���: �����Ot���OJ��t���o�S p��������af�U��	gyr�'��I矐��՟\�E��
?���٨_-|`���Q*)Γ��d�O����O����OdȪ7i�OV��@�˄��
W�Ўn�f�xR��Φa�	�����H�I����'����۴t�� �̱~Īer���UF��'[��';"R����X�ħl�����=xԥp3�Ť%,"-A�iR2�'o�OIy���
)FpI�.J h��tBX�z��6�'e�'�B(U+R��'"�'�����`).T�Ǣ Vp�X2�"D|$O��D�<��NA��u׺q����Ea��Z�$g�� L��v�'�Bl��"�'���'��D�'�Zc;R��ǲ�d0�4�B?p��Sܴ�?Q.O|��)�)�

�a{Ŭ��|���o�*-�6�Ȩl �7��O����O��	s�i>���A��z{�=��͝Bc䰫r؛�Mۧ�'��'���y��'����$�:L�F���̥UH���1�o����<��	���d�<����~�a�i��W�^ Zb�m�9B"#<ɰ��T�'�B�'}��ⷡ�46-������P���o�4�DQ خ��>Y�����sB5_q���c@�,�N�1��W}"���'"B�'mbZ�hr
� �u���?�� �[�iǼ d���O��D#�D�O��Y�31 EC��5�je����s|f�`���O���O*�@0����2���bg��7\R�A�ɨC�f%��x��'��'n��'ۘy��O�m;Ԣ+�<�r%�K3&��Q��Y�\���T�I�����|�H��Iӟ@�ɠ�͉5G�%K	6dc3�C�Q�q��4�?1L>�������$6�'u(�c���q��qy¯Ly�j-�ߴ�?y�����,��&>��	�?�c�mߤ�%b,�6/}�aW$%�M��2b�5��.��i)�ȸ�i�3Ċ����܏pI�1ٴ�?���j������?���?)�����;�l�!|H\mEa=7ڞ$��i��_�D*�&�S��J��\A��b�� ���*l7�<8��pm���Iʟ����ē�?!�ԩi��ƍ"���lɃ���"	�O>�I�4ϸQqs�E�%{�	c�k��A��8�ݴ�?����?�����O�������6��l�����\�dT xA�7�ɲ�b���I������>�Ą�v��g�Yx��̍�zL��4�?yD�"wl�O���?���&�(�A΋	�Ε�K�k��hvS����<�I�����X�']�ՍW4�F��t�����x��	]%~c���M���� ��0W\�pa*�zpd���k8ҩY��=�I�"�"�	r��i�����d�UP����A�.��0���Ӎ)�(�S%� Q�x,���ۖk�C�3fM�%Ǥ愉�B��#$��$(�	����ؐ˯68��-ƐX��x����rP(��L��,E�҈[�HHҮ�H��+pJQ�%� 1�V̍����i7�A�8���9Q�g���	Q��|�\8�'*H�?�Y%�8�dL��v��t��oE\Y-
����&`Jh�S���
hq���Za�-KQ
����R�[\��CR��'-�i[##�="�I��T�*B�vj*�̉��C�p�4lA��?K��[�>Yp�M�5��´��!&�`���4 k��m���<d�ҝb��J
%NL���Q8��#�$�OD�}���M���cb��xTK�,2Ĭp��g��S���a��B�@�0*K����I��HO���@;8A�x��j�;,�Sg.}��'f���@�d���'A��'��w,����*�%�g�� S� �+��&Htp�Cd�O�����ߥ21��'Z���#+ �!�,8k
ޱ�N�;SG��� Q�+�O@�j�	Y�����RD���
�a߀��CC�Uz������dF/��O�ўpp�"!�h1a..,ތ��%D�T���W.��L�	�}�m	0�!?a��)*Or�Q��ٖ	�:�p��1��x藯�9!!��Z��O0��Oz��������?��O�ZT������ �Ĉ�he�؉��~��B�ɜp"N���Hۦ0r�M�(`2$C��¹(�,�&��8�Xj4j؞����-ê�&��(r�X+��)�`���Op�=�"݁ ;�a`�,ٞ6�̚�Z=�yb�^���Ek�aKZ=���"J�*Θ'�j��������lZꟌ��t��p4�-D�<�2 j�2Q���<y������	�|J�e����&�|���U<,8���=9E^tC��#O�Mѣ��.1����2hT����k��xB@F��?�I>Ae���uc!��V^Ę �Ν4�!��d�������z	�h0�=\�!����m�CG�<9���hD�3����B.扟{�ع��4�?1���i�59Qr�5"#&DFIܯy���C��F8^�2�'�JA��'(1O�3?���	�{��L�⥉�/+D�s��Qg�$�;��?eó望Hz ���KpM1�	-}R5�?�y��$�-Z���з'�ft|��Dg���y2CÊL��k�\?a2IX�] �0<Q��	kw�Hæj��<��Q��YO��ڴ�?q���?��(B/"Q }���?��y�;E�&)�g�bE��C�/.B��l1�	�g���U�|e��ò�AzDs�cѨ�qO,���'M����2���3q�ž' (P�$ſ'��L>�7�B?�N���Q�`Q��@�)�~�<��f��^6�e8AȪ/(�A���x~��=�S�O(.Ѱg˃�^�ŁTi�FJ���l�=V�0���'���'���s���I����'B������ۇR�jy�u�;�h��na<�Rm�X$"X�q���F�����A�A����[ "ljkE�6?c"+�
�$9_.>��!�O�8f�\��ֱn�6 d�	s�)D�\��mߗb��I�v���f��('��9��'L���T�l��D�O�l�P쒊xR��4GڏAF` ��O�	�2s��$�O��S(��;��q�����G��ʕ���?��x2gr�d��Q#`)��l�U��UHvA��p<���B�`&�� xE�я�]E���oRZ(p�s�"Op��6��s�hP[���$E�4��O�nZ��q��S0�Urd�&%^^c��*2���Ms��?�˟��z��'ʬm���f���)&hO<J�	�'��kW�T���T>��H���#/l�P+�j>(�)�OV���)�ӈ�<�;��A�P�(���F�.��'��Q��ۘ��O>��2ˇ4K��e�t�E=�X��'r�eq`��6{���\75�u�Ó$葞�F�E/��X ��P&̙��C�)�M���?���o�D Ed���?y��?y�����a�@�����`���I��'V�9�ϓX-��!ܾІ�E��<5Z��=�PNYGx�Q�-��L�%��M*Ya�FHQR̓]q�)�3�d��T��h�T1Q�r]�4��;�!��U%_d4��r��X����&ɍi~�ɢ�HO>��4	�/g	��0��W$Ѣ���h�
�B�o�̟8�I� ̓�u��'��<�.�K�K"M��xs mUYR�X'fɯ[�!��9{&@9�M��b�ܳ�@s^%ON)�MOy�blTҎm�
f�п���'�xa�&J��V)���Yz!C	�''��R-�,@��cA�2%d��{�y�H9�	�~�~$Zڴ�?��v��b�&{�RLh�J�;�b8���y���?������=�?9O>�voǁI�����N?;�6���	F8��A�,�I������^�bz��zBB���d�2x���|H�Ġ�@H�r�`Q��Y��y%w�q�!�(}8�5AB!F4�x2bj�@���\$C+�<�$;r�`q�dŤev�n�����Y�Tj�%�?9P��( ��c&�9%l0 G���?�>&�)r������p	&e�	\.8�*&}�h2�7}�X+�O�L�����A1���=!T�l��>�"DSΟd�<�j7c�=G��#�ʓ�dnY��aW^�<�.�"����8 �qWDR�������iO��``�)L@�ʲ씂N���'���'��qѢ��'���'�r��y�G:cHH�WM]�nލ���6-޲$�c�o�}����qC����|���>i$�|��B�=7a�S�[%�rm���=b��p��-�d�P��L>��`D	�D�J�F�@X~����E��?!�O����|����@�N�||ʡ�Bi}���юd!��B0^	$)���=qplL9��ST����HO��sy�R�L|���㇌Aўa1"W�m�|q��GO�;��'mr>O��ݟ�I�|�7�#j�F���Y�e9��9  ńY������I��['/��q�*=p͎�}�"���Wf<ag/�)}zp�5�Fs��`
�A~�\�	t����qj�by�d��4*�0� D�`��2=,�AQ�R!ODX�sѪ(扞��'~�j�|�����OR)�0�D"o����t�=�]� ��Oj�I4�x���O瓳X�`��7�d�z�a��L<� ��啟��x�-����'Xfe����cHy6�F7{�4��Ǔ4��%�	J�I�}�� ��/�����i���62S�C䉽.���A���"Ĭ��#Z�DL�C�I�M{����@N~ seĨ>��3^m�%[�p#�iD�'K�ә�����}�,G��:^�� �d��.E����O���f��Ob��g~�Mʕ'~֐:���;9��K�����@J#<����UK&���E/1���[�CO�DÊ^f2���� |F��Y���)��/��KX!�� 4�򕆖�m�����-W9DaxR)�S����QC���Gв|�0!5�i�B�'��Ĺ���A�'���'���w�c0!/͠4�sOM����󤅊/z�y� �;ovR$2��͐:�� rG̴��'/N���3�l�I�W:
����
O���J�y�I
�?�}&�\�w��iq��z�j�tI�X��4D���$�q��@va�[��-�� ?y��)§*� �`���p����23�ak������?���y¾�6���O��SB,ȍ��ZZ[Ѝ��XYP�<020��a#�R?q
�:EL�z�l��F��6��C��> q���6 �F�Q&�@%�ū���O���� p�����z�xq�6�^��J��"O��bω�	>j����(w�p� ��UW�U�4�iŽi�R�'�)*K7}�������J�
���'��$�$���'=��,K�R�|���AK��тY#\����fZ��p<qt�IR����!��m��c�`	`�DY��\��	�g��d!���)�ب0j�?23��qpF�r�!��\��͚Bl�xzdk#ţW!�$��Q#��C2�SQ�G�B`g�%扴rQ�h
۴�?!�����L8���K7^�h��7vl�	]��b�'K�� �'�1O�3?!�ώ����'�A�YŘr��t��?Yc�ߥi�A��ߒX�(����3}�N׿�?!�y���g�$IV�"6�C2u�|��3g�4�y��ϼs�n\QQ$&p��Pe���0<�鉡`�>0��"1��2'Æ,G"�ڴ�?Y��?�-� CF|0��?����y�;2�����6E<��"E�H*LԘ�y2)E��<Q��8��afl	�HӸ���$O`�J�Ԅ��qD$`�ѫ�� �[bA�� �4�<a"A�џ�>�O6=��۬Y�qa�J]b=��"O���֎��c܌|H&@�5�Ը2�������5`/���7o[;zy����iT~h�9��ԉ|����۟����<�[w�R�'L�	�4e�ZIɰ�R�]z�#v)ךZ��J�O����ؑ]P`Q�NܴU 6�[�G�4!�Dؐ]>@����D<%�,y�.�*�L�à�'/��%U&BB!��n�'�<=ؠG���y"�2��p���!�F� d���'|�b��P*���M[���?!�`�)�+��D�6`��
h�9�?a�'ϢU2���?��OUX�
����3_Ҵ`�2&�V0Jt��g�>l��	�g�P� 	a��iִ��t �\��3�;O�I�2�'��'��	[ҧO58�NX���L�z܆|!�'����3JL'5�8��ڃ(p����'7-ȓ	�QcLB+~��X`	Mx1O����K�)������O���Y�k86��� A�e �0B�#)"���?�vĂ�?y�y*��ɵS&���@KE��jq	�|y�'�������S�b
0�G�TO�;H׷)��'�����o�S��ᰄ�F���
Y��AUq7���d�<l�ċ� �-i7��?l�%��'�HO�W�m����nL;	D�����Ц���ҟL�Iw��)R��ϟX���������B`���/�=
P�ن=�n��E�l�ݶ9�牀?b(�v�9��ݐ��!]�x�ԒAM<<O��{4B��crm���d1��.�I�����|R�� ��hx'CU{T,�$��?�y�a�M����	��P�F%k4�ݵ����}���Xa���_<�����b�4e�׊H3�ѐ���OF���O���캣���?��O7�}a��	�0�R�3'"��k����x�����b�@���Lit�7J��	x
�'���zgI�yl�h �ڏ[�r$�aݢ�?��3�LL[�`�]��H�g$M��m��P��a� ��ZHB���Ϝ�Ѥ��<q���I2n�ȟ����2yF=
�i@|�@���μGRY���<���������|2Q�M���'�S6E� I��9�mC�AH��$@-O����$^.g܀�#�
���I��e.�xr�̎�?�N>�үN_,�tSq��9.��)�A��l�<!%�@�c���6A�(�s��c<�ֺiJ��1n@B�r�o����юy���7-�O��$%��HП�ڂ]H������5ipxf%���	�}����IG�S��Oި1Q�U�1�~(�1��Fȋ��Q��ɔ'��?ŻDl��=��;�ET#��{��*}����?�y��d��6A��� �4>�����y�l]'eHN1q��[�;�L ʧI��0<���I �n�[d�X�Xް���ݭI�:�4�?I���?��ߓ@�,�:���?a���y��oa���u�	����̜�<�����y�(����<鳦��|������ϘO�TbծEFܓ,!�!��	�����T�3S� �S�	��<��	ǟ�>�OT��GoR:#SlRc�94�*�(e"O� rxSb0W�$�A]�s� L�ѓ�T����Ӥ)=�m��+��sW�J�4�Tz�^�����I��h�I�<]w�2�'��	ٛMFT��֤_�>aD��gϟ�p�8�H!O���fP�cN.��M�7u� a
P�!��P�c���CE�ѲzV�m(6�ІwK�H�7�'����H�:/X�'G<�R=�5\��yb$,�n�0�����,�1�K��'n`c��+�e��M����?�@D�.Z.��h�SQ�\iسa���?!��J��p��?əOh.t�������0�B}�♒wvD�#�����W&yXRH=�D�8����];g�xR�ÒOv�x��$�?Q���?���n��}x�`�.Fk@�G%�6L�.O��<�)�',=�,�Y��i�PgZ$���S�E��.�#q��z�H�	�y�Y�`TDA��M����?A-���Ygf�O�)!A'"�@�6�� |�����Or�/V�P��8�|�'	Ȅ�V��ň�L�ʞ��M�J�"5�S��=�c#E�f>"0�!N?y�P�OrT
 �'�1O񟰵�a�<.k�|� N�LM��R"O8��eƟ����9����?�����'�#=��Ԥ\�x�Pf#	E����p�e�<Q�
Ͽ&�j��hS��A�JH[�<IE�Y7]'�<�#ꕄ{���'��@�<1��vA��8�>e�D���DJy�<����� ,�����(F�4Ɣu�<� [�q쎝�0ǚ'��y�q�<)��عkp���hYi�N��v
�D�<Q�LY�< ,9#��#D�-<�TB�ɷL�^=��%�%)-��FIZ�Xz6B䉁~x�j7%?G�$ W�ԙ_�FB�Q�^�R#�w۴Y��a��Q�
B�'Qz� ��"p�ppɲfVOgB�	���ɱP�6�A��^"��C�	D6�[q��^�f�G$���C䉿�[��I�*��x2c�&m�C�Ɋ>r���0_��c�̜o��C�I�Y3h���n�,Z/�	*�I�H�C�ɝf����R)θ|VZti���p2dC�ɱ_hk%b��r(�2��{�8C�	,$�Έ�@�)r|\����1�jB䉵v��dѕDE	0u,9hua�y:B�M1d<i���9E�����Do@�B䉍7�Pi&�;B�ۤ��l!�B�I�TS VXMI�q.Hd�vB�	C88�@#��v�	�#��1t(8B�	�-�� �Ӧ��\��S1c�:"B䉽:pR���U]�(��A�1��B��4���'�]�~`�pBiϋ-^C�4�D���6!��$���7y!�ȳ'�a���}I:�`�@4i\��^��x�ؕ�ܗS�%�q�R0�y�\� �H8SiD����`!��yB�܇dq@��U̙��E��Ȁ�y�D?I0 1n�&H���Y����y�Ѥ ��5� 圳/�ډP�����ybcS�줬�ӫ�7TA�²K��y��i.�'�<)Fx�F��y�l��H~b�Q��|�Dl��@B��y�7D��	A�S5|\�qA��0�y�g�3=�4c�O#z���1�H˶�y�m.O �jamW�"�J|l�y�
M� �|��¯�'��l@�P;�y�kE&(R��V
jqzҡ��y�ʖ��e��A=[S4���L��y���/L�d8��3VD������y2��5s9�P�E(FTp���9�y
� �9�C�*��Zg�,w��y#�"Ox*��0`*��ꢀڧZ��( �"O�8�'L�Qp�0x �ʊ_�b�Y1"OvEa�n��i������N�9g��1R"O��q�ħc����o��za�%"O։��}
h4SnR=`gR�a"O��*��rK��� ��J�kK��"O��a*R���Ap� �L`�z�"O��(���]�t���O, O<)��"O5�S��)�P�2&IȞ��q�"Ol@kU��(Am�F�ʍcr	�%"O�x@g�� �A6�Wh�*� T"O �Y�
F2��4'˔@*y���'D�GIʭ_r�� �q~�qb�!3D��j�Ŏ�`�dX�+F
b&xI�1M%D�l9��1\���c����l8v9�-7D��`�mR�\?<�,��^��5�4D��)�� �<E�xᤌ���N�C&1D�\2ri�3?b���ηzb�d�e0D�L��C�:���u�J)Mr
m�r�:�OM����?5ԭ�c��O�� #�8Dw�@�D�hh<1%�C��,���*�2ՔA��Lm�'�\i���/<`��~�boU����#2ᕒ:��t��	�c�<��MW1Z���b�ؔV��j�J�۟4�EhQ�)��m��>E�TLM�c����qo�3H���J��O�!�&pU& ��B[��\�QI6���	ieJ,3�F&@ay"ɪo]9"+�crT{��tڀ��V�<§,l���$���'��4�iHB��ɺ=
�'���he�@��Lt��ўm�L̓RnHQ�%�1�u��O���&ΐ}�Y�U�'��Jߓ\ͮYb�L�>I�D��/g�a(���*f*eR$%�<��f�������8�7�۬����cdK:���!��dQ�<L�E��HϴBx�J��H�^(������$�Ǌd������k���T�'K�ɡ'-�H���Qj�	&P�50�~�1O�Z�OR��p�Y\%�b�IB�a�>Ȣq��2f��T���K,�졄�����u��KW�r��B�A4�(!�\Y��pMA
';*5@��2uJZ����9/���>�� a�3s�Yp1-QR`��K�!\OLl��<�剫U��pooK�,[��� 8o&�YCg171F��hѢu�n��n"�Ӓ/�4�&U�5CS$J���i!B�{�dL�=��!ԿA:6�E��N̈́JjFi�kN�U;,a[[a C��|�Fh�gV�5��`X%�6PD�Ї�	�>L�hH(� ~�<�s1�� g�q�[?1O��{�O�R �7� /7���!� �z1"��JRв��ƚz���e�m��i�U4Bt���Q8|�8Z��-AY[�#U�3���ɝ�U J�B���5��U�2�H
�\��RT�c�;/h�5��{ ��ʰ�Cr���������P��V����ְ;U���΢ʈt�g��?���U)t�^�[PH�?�����кCb/}B��4�z����t8y e��9��'��q�7�	O �3��;l�򴙇��z|�0��`@]�E��-_�9�j�����X����IAJ]ax"�#�T�5![�P z���N�qb�|��Xr^�3�BU ������' Α�'�+c��|��gl�4^��$ �ak�}��o��t��$1\OU1C��2"�P�Vnʇtp8�`�@@5s��a6�/e�}J�cQX$��)^��S���:u�=��T1JY(�#���2�Ґ�9p��IV��!w��c�P5Q&}e����>271O��� ��xr DQ�q�S����7-�!u�e�W鋰/	0Qa���J����56)��3%Ձ,*�awK�CG6���FV�d= ���;67��r�l��dTH����䖁c�hc�x�ׅ��f����)�h'�ɢ## ���9�̩�!�]��l�'dй�f��kZ��J�*�9m]���A�;P��I�Q��I��I�0$�2�d�obT59�h�:!+FDG
	SϦ��"NE�C���j4�|Z�%xmRpbgoG�C�,5� ߁T>�H�'�����9b$�3S�˙w�8|�c��01Y"N��?y��5|��(�	���T����q�?�*����]��@�� �yl9�O*��%k�."]�\8!��A���h���-`6� �MߧW��p�ϭvY���޴̪ɻtJ"�?����c�YDu*9��(ԕ[ن�	?{Nj����-!��pD��?Zz�B�)=:x���N�Vt�)���
�? �������UxH(0J��״
�̌����3<��ɏ)���[�E''�ʰh%�P�̧U�P0�}>� L�C�V�R��A�E�`���jP"O~���̎$�zRo��-pk�m���JǛ�guf�؆���n��b�?�	����0��+c�Λ�f���H2L�!��3p�l�k�G2Ҝ�ƯI�$�zU�.�]06!;�+ݙ*|��K6�O&��1	��Obd�'�?Ţai ��?��P��'��(*[#I\ �k�`��� ���WMb����e~ ���o�%�~2M�*�Ї�IѼ��$"z�(��\���'���U�F9Jd�&*����V8���*j>)2�o�z�G��)x�8g�ͻ�y�ř�6�ƀ�va�+%Z��Qj� Jڜ�h'b�,����p�b�VY����w�!�M��Nm����I�,e�
�:�'�=�"�D�]n����Y(�l���3h�N�Y��n��{򄂄7T��bg��TB�C�Ź�0=�7M�-j!�RTg���o�~A���$�:���R/k_�C�*?�X��#�8=�@�`�4\fb�@�h��f��G��>ki���m��r���2�$0�0B�Ɇ;�d�s)�2H�*}���)J:�l�'DV�ēt�G��O�Ђ��Y`HBv�I���4"OhШ�M�Q��a�$]�E��H���:��5��'/�M��Hڶ	�L��y���דC���pI<���Jج��f��o�%dH!��$oT� "�F���43ƀ==4!�]�V������ j��pO�f!��ՈUFR�Z�I#�̉b��Q&~�!�˰kV�ȡj'I�&�x�#س5�!򄋥R���pc��!� %z��Q�a�!�d��VdA�ƤD�[���c�A !�!�5V��4{�ՎF�
�P�S+&p!�$O���Ի$�;�������!�@$8pp�;pl�cb�џf�!�F���=��G�ye�9��QX�!�dţL2����>X�t��ֳv�!��4�t��B4`���צ�7q!�D�?Q��R�Ѐo�L@�FSw�!򄃓:�d1FE��������9|�!�X���0�G�+����ˀ�@�!����Xh�G�BȞ�2��O!�D�7L\�x��*_+���h�+Y?D!�d���0	���Q���x�+]�~�!��#"�*�ছw���ۂ�[��!�8�I��̺,Ąx��� �{2!�$�PR<��e�G�z$q0*+*!򄃔�������z�ڥHN8�!�d�0h_�,e��̨!gm�%Jm!�D�	$��y2a"t���͈�PQ��{�E����*�5��s�8�+"�T3F����e"O�)���%�
Aٓ���E�*���8}�W���O,A���B���ˮ%�fuH��ݮ
A
xz��ފ)H��}Bu���ظ�8�I8q�4�[��'@X<ibGװ/R�s�o��Z�dĊ��đ"~d-H>ɉ���S�H:r�̓!`TZ��X*>�@��=Yi���Dmt$�����'���g~��I /�0���.O}}rc�22b��'�8�&�Щ�.i����[y�L��4OsNa�g��<ɰV�u3ʝ�F�0r���B%c�<tI�|�`"��!{x�+�I�}mp�r������N�pe�[� �.IH�#�[���"O��RE����U����C΀����/aX����|r�����xn0��5b��4���03	"D�H)�m�;{q�!���d�J�3 ~���' $b��dģ`�8���bX�b�
@�a�!�䀣0�� ��S>S&� ��V=3�!�\0@$t�Cu��{q$���]-!�ވB��Q��ʴb^z)Vo·�!�]2[�QɡH���l쨃��,`�!�U�
ib�����@���R��"!�� b]8��ͦ>�0��ML�HŃr"O�QbtKԫC����nS�n�@kS"O��Zϋ`�I�U��
0}Ba�"O�8֦�)<�ȱթ�2��<��"O��jb�*p��``�i4rh�+ "O�EB�,3�(8�&�P0V]0�)R"O Q�aDC�,�#��;V�VY��"O�d�`O�^Eܜ�����p��r"O,�@e+N-t�:-��Q,S���f"OYH��7TM(���m��U����"O��j%"$+ɞ �w�I#8��U�C*O|!ʠe]�4d�Q.��>�|��
�'뼶NF3H��l�%F�aq��a
�'�f8he,��OdV�%���&�	�
�'?rL�r�4o�<H�)���8 C�'k�U�tAI�`�ʭ��#_���'�>4�rb��;��|�ר�0a�'4�	�cO�X2t��'E?�, (�'��pw��q�J���BH`�'Ov��(K/i�i:e䘿�<T��'�\�H�T`L	  �
#��@�'�R�Pd���hS��v��{{~���'�$3�ǂ1	H�0��m��Q�'R	�cϗ���S��a��H�
�'���!�E�H Q��KJ ��'p����Fb�9`B��x�D���'�N��n� /� t)`��#��Q�'�����'u�UyT��0@i
�' ��ufQ���Q0�b�6'���'E�e`��A�ud\�T+��T����'"��cRMS�8��_p�u���y҆R�[�^`s�.�r`�%JKL��y��+@�nU���i.nq��/@��y�$R&}�^���\�Z�ؔ�.�y׉Q�^�p��4R��D�y���H��H� 蓫g�Y����y2�W�\B���.�p���.Q&�y"��8׶l����s#ԥ�y�G,T����\�@�@R� 2�yÛ@^j�+�9���AA)�y�E
.����V �� y^=h�� �y���`�(�Yf���,�nT�ʃ%�yrk
r�
���[\��x�4��g�<��o���7�V'z�� ��r�<�@��=7�䔠�i&A��� ��\r�<Q�(N!o��"@��#Yxy���G�<PCO�O�\�9F$��paȀN�<YpK(��Xc�D34�S��	R�<A��V'.�2`��K�?`�N��flI�<)��-e��T���A�B�8��bF�<�@��S��	�G,q���a�F�<��)J��xBiے\*� �D�<9V$^�k$ҽ����M���v`ZD�<�@H�o���ʏM�F0y�o�}�<�0�зP����jÉ,
�	���^�<r�D�(}��F&{l�h�+^�<1w��L9>�Z�&O�R_�� �C_W�<�T	�|��I�P�������G�S�<alT�g����v��12���4��N�<��˄(Tz��zF��.�ݠ�a�c�<�BNI#a�V�q �� &v���X�<��/۲E��F�/#��3�d�}�<�D��z�@Y
�n�>����VF}�<�u㜱6��(��\�(](�� �A�<� ���!͈;ntK��]60.��07"O�Z�Ȗ�E�vyz�蟹s��q"O�1�v�&�$9���q,���"OJ�%@��.���`צ^�%����Q"O���Ε�9Q� 	v��r��;4�Ip����Mm�H5h
5kLЙ�*�!�Ĝ<?BV�"�O.p�Y���¢C	!�j��(��=Y�E{�鉹0�!�d�G�a����{nV$���˪vA!�D�~��J�㗯S^2h�(K�g,!�$Ϙ��5��S�&{�8�(�z !�܆X�Z�釂��7d0]��	�Q&!���-
�)9�	�*E��3&�%!�$�7Th6a@��$:�*feE24`!�F�)C yS'��l���C�->F!��RI.أs�ZRG�M�B�8T!��0r�r 9G�?b)&�IeO"�!�$_�-ްy�&ԒP��I)��ߣ �!�DVv��(u���Z`�R`��q�!�$�mkh��@�^2OxJ�z֌mq!���!Vv|-9 �A�%p��"!.$�!��J�� � ��I�@�tLh7�X<	�!�D�A8��X� N�s��	vh�?�!��߻W:,�Ճ�|`�@��
#j!�$̡E��u�!O>��d��8`!�$�p��1s� H�`㨎^_!�dʺ@��Չ�C֗I�h�p��JI!���7X:$����׌�T烄N%!�ʁ1$��ŕ2|�d�y�l�4&!�V0���H¬6�tqp��5w!��ϒ6ª���4C� y� �]�lm!�䏥iPR��k��ZD;��>e!��\�{���+��q�V0�dςgY�䓠>ma~r�qt���sM�.Nx��q�Y��0> �"}blD�9�F���X�B���:�N��y2%�p�X[�l!6C(�H�`:�O�C��O��볫�LOj���Ž>���'/��	>E;0�I(c�V=��%PT���>�b�|�mȢɦQ��*P�ȓ#����UeYva6����8�X��	$��?��"�#M𢽒�B��%�Q�ii��t�c E�N?���'Z���E��DD8�(�o�� >z���'�����SES��B�u�iÌ{�'��zc����X���G|�q{4a�b�i�"O�y�"ʋWd`� ��,Rڌ�C�n�'�"}�'ʰ�y��G/c���IWÇ��a	�'�6�с���K�d0��KЬq�
�'N:9�TE�9Ħպ!n��,��'IdѪ9�p<���+V�a�'�Hl���N�O���� U:A׸8��'�"�[v�S+M&M{2$B4?.� �'���X��Ѹ;Ni�QA�C��)��'@�᫑CE3�n���ڌ@���	�'>H�;��ɪu�\˃i=��h�	�'���b��.������/0h�1@	�'�p������^�
�5(ښY��'�Hy0�A�v�0Y�UA/z��ؙ
�'�A
�+̵�F�r%��!1X�k
�'��:��Xq�����)e3
�'�ڨ��LΒ+����X�Y1fP��'*���E�M�mt♂��#z�t��'�� ��%N.2>�����u?,�h�'<���7����rH%|2���'��	��L".Yf5��B�l��M���� F��5����V��O'� �"OV*E�;*�n���*g�����'#�$E�����Н[Ө�$��g!�D9|�e�Fm��+�d�hPMӨ1n!�M�mZ�*���;�B���Лe�!��y�h�եֻW�4��/�@!�䝧OGЁ 1��5e�@��@F�!��Eb<�l	�,,�0ϙ��!򤐳6��U@�5�"��=}�!�Ă7�FE�v ��?����k�:}!���hz�q���:}[�	��m!��,m�X��܊'e�iO�=e!��7��Z��n&p�+���5e!�F?;�dUX�� D'nE�-�!��D�F �Y1o�	D�(��*D��!�Cv̘�b��nd>��6
��!��~F]��I�`d*qr��1b!��*.����&[�uD��XE�ɗZ*!�d�9`ޤ�AO�;I?�0@F�1y!��ǈ4��XP@�>��Ԉ���=�!�D�O��Q��G�}��Q�!�V�qJ�����b*T!!Ȯ �!�D�.Y��e���[.��ұ�\�L�!�To�5;G$Q�H�0��*�{�!�Ǎ1g긁�[f����2$!�7dH �B��8.��֍�
�Py�B�p��@�m�t�P '�։�yr"K>� tRe
�)t �0�*��y��"Tք�2`�t�9�5���yҩ�#k��	��Ǳh����u�[��yb�V:���8%hB�5hH��샜�y",U�@d����u�Y+�L�y����H��G�~����yRЭil�@��	z{BU�`�ߧ�y�@ߢZ\��H���>2�py�����yr�S�&�l9w�7G�@S���yr�D�w�%	��=�VV�.1|���.�jĤ	�r=*�Q5�U2L��ȓJ�:��J�_|��sp��/H�&ՄȓL+��w���.�@���.e�,��T谨�,T�A�8B�h�3!���ȓ
��#�3<�l�br��:<�ȓ'��}2��݈zL&��O�in�D�ȓpi��kEP�x���&�Զ0�0\�ȓ!k���e"_�q�8Ë�0z�P��ȓV?�B�.J5_� �"t�4}C�U��Q �̩te��A��=b�a�
- H�ȓ|��aPK�Vg��	7�mת���;���� \�\U�I�΅�-[p��I<����h"�e����>�\�ȓ8~Q�ì0�����
�3=�2���9������68,a�,w0�����S ���9��I 7gӦNĄ��	a�'��E��C��&I�W��n�^���'����1@�����6(O�X�v�
�'9�t����&a�*Mt�H��BК����)S��u���ʝU}��ȓ+���萞M�|��%�Ix��P��Ѩl��ɛNy�`�C��T��]��F��{�bȪn�b���ϨyVń���-Y�)��iR.\�H�4�ȓD`-��].^���h4�5�☇�_���1��VU�F��?[�|��-�p�f^ e>�h�V,u�x��S�? ��B���?@m7���.OH�4"O���vHW�3�z�E/�046R��`"Ou2S� Z���Boөk,����"O�Q�F�'S��)Qm�m&Xq�"On�J �%W�1C��9Xt��"O����Ƙ�<��5z�a��N@���"O�x�(|�n�J�%HIM�"O� �a��8s�r #CCBE�'��lZB,V�!�Z@�#�Z� �zŃ�'l �� ���R!�E,^�J���
�'���	��ϒ0�&[�dǷ
'R)q
�'�fd�đ�UƼD�2�A� h�$�	�'���1`�2eٚ��V={K	�'ӎ4�E�@ȝ�@���v� �'٘���C��[�^�{@/%�r�[�'z���U`ڥ�
�'�Z�wp��'!�L�c@�.�p����j$�X
�'1���P.˓x���U��P���X	�'��k�F��c�V8��Em̤��'+\�а�M�7
h�:b���9Id,�
�'zh�R��4a��ĭ�2���
�'���Ye�Z(fnd=�D+��y����'@�˗d5o8�L��6�:�'��ir��/
ظ��L	e�B�"�'˰�"���R)�Hՠ*����'�
�<F 4�� cY�MJ:x	�'qt��g�Uq ���.|���	�'��AQ0���'��'�I�#�!�	�'�N��,G!�@��k,-o����'�D�0&^>f�Ա���Dl�A�'�*	�$ :LO
4S@�+�����'���a!��n�1���������'�ʰ��E��u�O�� �'�j����B� ٠�&-5
��D��'�����$�lq��":
!�'���ԏ��K9�����<-h�<P�'6l�R��>��6V17�\)a�'3����m�
w0Xi���/%�z���'i�͑t�
 �f4�C�#m���'2r�2�F�j�i���<n�Zi�'&�iX7H��T�#dE�<"�8�'΂��5I5nr�`c'�3:P���'zF)���޻{���S��4k���'R~�Vi��w�T$��`�:��J�'3<������;�`���B�d��'�,��@$J3ex���=B5�'����U/H9���B�a����'�l(��۔BoJ�x��#c���'vN���g_m0������.0=��3�'��<������P#�ַ!k�"�'��i��nO:`���`eN,�9�'J�)��ĺBE��ևծM݂�r�'v��"b�	>ML��u��L�f�p�'�v��&/O�&P���� PK2~��
�'�6�2�Ad �SCS<���'�r�腮�.8Z)��@��g�V�x�'�l���_�|f032��!dM��I�'qd�Y+[�S�l��B��
V�"��'jX=[�:w��|	��Y<UFV��	�'���v�A�N�3J�M�n3	�'���'Te
.` �o��{�nU�'ʲ5s���h1^�����\�3
�'�l�B#Ӵ<�<]X�kX�~#f��	�'�vLPSl�	Mު	�ʔ�qI�}���� ��ʢ ׂ�^a�7$ܶw�D���"O^ԁe`�*��,�1���w��P&"O�)aEĤ*�D9L\�`Ǣ�x�"O���$CP�gnbTy 놎g⚌�V"O~�AAa���Y*����sl`��"O�T0��2d�m�b(~d�$��"OHE�#�ޘj���S�o��IR�"O��v�ŌO�Z(�Mǭ?RL "OD嘦�H_.��b׫�82J2��s"O�ۣυ_JZ ��N���]�q"O
x0$	�)!ʮ�۔������q�"O��r�]��!���\�(�ִ�r"O�dQ��3b. �4%�z)�B"O|�ˤ&T�Ȩ�v�&�j!"O~���>kwB5��E�=%�ur�"O��C��*d6� �
(�m �"O��3���m���n6�#"O�Q�Ƞm���#�H7w����"O*�ҧGK�F�P�hF^�#H����"O:�S�,��? L��$ʉ4"FJ��t"OJU"LӼ�r����-k6�B2"O,�����T�^11��[4>!V�"Onh`Av]x<�AF͘c�� �"O���''��)J��$EǳlYD[ "O����+��w�($x���(�@<�u*O�5S�M"��!�ܝ5�,��'�2��v� �<g^��b�9k��Y�'`��y�S	����,�@(�'��`�W"�	4RH�1�+X�:��2�'t!����x�QV�Z�@a*�	�'��`�p���wB(�إ���@$��i�'^ӅBo�����Ƙ9��4��'��,Am�<�8�Q��[�@.�
�'�:�S�g�`�j�kq�� 2���'���b�I�/`�`���E�;dp�@�'Mxۢ�ım��Sa�G~�x�(	�'3dy���¬>���n��jvv���'�D��L�U���A'��d�tȳ	�'�1`�fW�N�Б�w-B�q����'�V�]�R����&H�A���@	�']�d��&]�Hx���׃
�GfdX�'�����d���(��GyVԘ�'d�\���/B�4Ӵ>�ji8�'��H��oT$�����?_��ч�\8�,
�c�;����5�����ȓ ��{Ԏ	�&�`����*��@�ȓ_l���gت3���� hަ(xD��h.M�A#'�X'�(v ������]�a#E
Ht�y3�&7h$��5�R1so�9�0�#$�_$I�	��0D�Ր�ѝ#c�Ļ�I�@` ��ȓ]~�I�ꛐ�L" Ћe8��s��CT��5u<��W뇄9G��ȓ�L�C�3b���*�a�>Z�4�ȓId���"˩gI�Z���:6�U�ȓ
	@}Q�%� ���r��:4T�l��<���g*D�ĥ)`���0fv�ȓ53�������d~�� ^[�<�AH����Y�hߩhQ�DӁ B�<	h�&\��U��]�s�����{�<1�Կ|
��"�*k�X�h��r�<$bW9cɜL �ѝEzL�C#Jo�<��MH5�4[��B0=4�В��j�<�$ŀ���$ �W#��x���h�<� ��0��ۑl1���i�up@�r"O��;w����}2�>�8��S"O�t��i���0�B� ܱ"OR�cw�JA�4���8�P�I�"O���aM�$�Q�aB�/����""O� @틦���#n-_�H黡"Od��(��P����-ɤ;I��$"OD����
`Ҿ��JD���|	�"O@� ��S�~4y��M���ɔ"Oڕ��/V���a%��"OP�AO�PPdY#��)g`�(�"O�yZ�I� ��`[��6hT��C"O<9�Q`�#�nu���='�i�"O���f��NЬ 3��Y�z�z�"@"OF�"���DśЉ�;��a�d"O`�X��]�$d:�I��#�d�x�"O"��Oؕ0T�10�͈�S��m��"O�|:r'��]� 1�'��~q���u"O�ݰ�� Z�6��6N	�`Y�Xr"OJPT	�6@���[�VK^s�"O��EBT��UZ#B�|&�$�"O�T��� 9�N���D�4)'"O�$�! �?8�\�y��@;Y'f!�C��F�O$|H)��>N��lx �����	�'���X7��A������Ǝ��	�'�"P� &W�8X�hI3 g�J	�'Z�ui��: �L���"~YD�ʓq�H��-S69�q!C�&}`ȼ��v�y� dW�Iњ@����(7\e�ȓz�hQ�g�`�J)�
0un�ȓc���A0���p�պEϮ=��͆�	2��wF��!��4��.>���ȓA�.��v�YT��A��z�ŌG�<�#�A&:�xIǞ�b��e�D�<�%��P�~�%���0�J��Ɵ��'aɧ��dJ��u
��@Ws����  �!�dȯi�x !-)`*E�c`D?V�!�d-������L�d�¬q6j��Q!�D�K/���,ͧD��`'�
l!!��*%BEY�C3Z�&m�� :!�G�.�&�w�э#&��:��Ͷ2!�d�E��%��P*M��b[�~ў�D�I��4��pr���<�#��k�'�a|B�ςs\dU��D�;w�h��(��y�ɟ?j�t 'f�k�t|rp�@�yB��|��|� �ʓRg�d0����y��R&�0@��Έ�?�1h�,�yD�G��<Z3@���:��ÄQ���=1�yR^]^ �
�nE�Z�`M ƦѼ��'�ў�Oi�ԑ�)�,�`qzE�[�T��a�r�)��È�[!ZM�s�Kd�,������0>)SÒ�^<1��D�vP�͌J�<�h�Ysj�z�5'<b��0*n�<��͋�����'|�����<���m��C�IT�)Np%8�ɋwh<Y�ڸ`���b4L@68)�F���y"�X�Pe�a�2��.3 ųꙄ�y*
	$�.�	!��Q֜A��Ƚ��'�az�JT={�
�ׇ�7���+�Δ�ybа�8����.��4x��˴�PyR���t��ĔJA"��%AR�<�ӊ\�>�(�G
�> =a��M�<�u�V��Px�p�I����`TGy�i>��<�掝�h�@���M5�LRp'�{�<� ^��r�Ap���R�7f�Q�]�8E{��)���}���Ϟa��L�c���!�# P�(�&�@�z����O!�ęw��;%d�5$k`�{��Ǻ?C!�d(��{A������N
H!��$ �x�sC�:�´�Vh�9!�UVo�����N����1�!�d�*J�:�c��זwu*L�c��2�!��N#� ��%��O����ue�N�!�DҐA��;%	��[R(3�Ꞿk�!�$�H�<�����;1�]`�&)�!��X�^Te��%�O<�M���ѕ!!��J�tt�Gτ~��|�qG	@!�$�g;�I[э�}P�}�U�1�!�8`蜥k�j̦]0(@!��f�!�D۠?3`�d��J,)�g��'Pt!�d�O�n��]��r�#�.�=`!��K�"��+ŬU�vCGd#T�
�';"�$�%�|�DYf�H�'���#%>�� �&M���x�'��걪������+ֿ9�����'
��!K>O�@��C�.#� ����xB��Qج�#Ѩ��Hql�0���y��
�ܼ(�N'QAV�Iu��yR�ߛKM���#���>���+�쇆�y2J�%~Un�@��A�^s�l�r�:��>��O(�s0�S6dD�a ��RE���""O$y��9;,qI��9=p��c�'�!��7lV�]zB����|��1��_u�Ii��(�0�c�))�`3u�M h�E��"O4��mA��lT��߯%:�a�"O�1���즙�en� c@���@"O�((��P9 ��@����q%"O|�Dɕ�F>�k���%{(�B7"O�%���-q�
���j�	h�}Q�"O��s�)^-cEv���α]�t��"Od ����(8t�Z�ϒA_R|�t"OP0#'-e%ZчLܢ[W��e"Oz��t��#3q��)S-E2�"OFa�7-�<U��4)��?8t,�V�	h>�1h��0;��1sD���� �d6�S�''��v�Iq�Ա��}�朇ȓw�X��R�ǐ5J<\���{��!��)@�)���oݰ򡅿A�.(�ȓp@@����T ���#e��A�ȓ}�2����h�*iK��Y�~_�ȇȓ1��d����7k�[�}�,X��7v$`u"��6W� ��'��_�<r�'���Á�T3�����Mp����'���0w�Hp��K��If���'�0��_�AH����ǗJm�܋�'�L���fA1��x��P� �Y��'��1s��;!��j��>���i�'H�-��ā<EP�X�Ïb�J�'�4���'�-jݸ�9� (x��4"�'ϪI"b�����4a���w��٫�'l�~�)�' 	:�%Ǩ�[tE5n� ԛ�'r��XeM�̸,�6������'EָP��R?N$���ku�l�Z�"O�]@�l��sͼU���
���rD"Oؼ����[~"�Q )L�g�Ne��"O�4��M��A��I��>5�!�"O^ �Q�]:5w�tqṽ�;�v8�S"O���&b]Q�V�j�A�M� sS�|��)�3� ��	C�C�L��%pF%��I���!"OF��ЧEI��1�~�>���"O�%�*����]ѵ�Р��D��"Om�ԏ�b�8�c�#� up\8�"Ofq2r䎌vN(<��`�<�"��B�'��:��uBD�#�L T;n��$�7�O��h�tC�f:Z�0b/Ɯņ�_V�U!$�Q������E�mL�d��w���h�B�������
�EbQ��C͜1�H��j�9g(��J�P"O��Y#
A:J̄��@�fi�W"O�y@D@�U�p�rA�&N�X�T�'B�'6+��S�v�X�ZW��3s�Nȱ��'$���tŁ��R',��e$�9z�!�DVO+pɋ�,�G؊�ycNY�F!�$/uD���G�"t���LIk�!�)V� ��&��!�z��jG�X�!�dĽ%�h��&��)S�vY�"H5,�!�O,D�u�`��2l��Ő� Q/:�џ4E�T�;j1�)�G��t�~�ʧe����?q�'	2e�"�A@�aK�gA�z��Y
�'=l(���`���Q����ֵ�	�'�@I5b�&JP&��d�q���Q�'�*��4�ݹ�~���f^�y���'�8\�1l�?W�4��I[
\!���'xz�Q�@_� �RC�� W�؉��'~Ř��^�ǳ�$kA/�^�<Q��V��H��G�	��jS��^�<a�gͨL��!����fT�02��W�<����!`:�%��M�61GRm�C�CW�<I'��|�8A�e'�5q3F��h�Q�<�U$@�L �ݩ�)ʳ/�	ۃNX�<�b �+N��ш�i��2�W�<��):N(��� B.t�܉�&��Ux��GxD'�P��Gɘ<P���*œ��yB�4h�%���D�K��|�S!5�y�b�Bg�PJc��C?�`aC�Z�y���#$��U�޹h�̡	��×�y��H�jF
�j�́�l��  d���y�i[��ꜱ��._�t�"J ��xB�9HP���z�||9��I{��t���ᧂ���r'p�йZc,D���GN�$:9%O�(V	�Ã�+D���p��:`6,�Q�T�� `g)D�Њ�g
a��������k<D�H:���=t�P���^1&��9D����L�u�:t`$�Ȳ\P�Q��K8|OLb���/��/�"�R)P=��H&K4|Ob�ф���G��$��ďoU���O2��k����եB�fwB�R�ˍ6X�
�JfH1D�𪶌^?5u���!k�
��c�/D���rC}��P�f/<����S�.D��а��o=�FjKh΢qKn-D�8�N1.�!���Y�l�(,D��
���Z�4���"x[Bz��)D��i���&�4,��M܏�� ��"D���C�$@�-�W!ږ?��� �,D�)`���Ɖf��po�!�=D���b�Y�F���R�&"Zd�1��(D��z0a��r�[��S�C.�sŦ&D��A1�{��5��E�&E�����"D�XOQ��tCf���H6�	�'�"D������Q��ͦe9Do�A���0=�t��1)>�i��Ԫ�]k�@�z�<� 6y�p�	).~U{�@-)��Y�"Ot}!e�Vj80��N��D�q�|��)[*X�`�dc�$I!FO�yL0B�	�4����V}�<�Վ�	�jC䉻5�	PRM�5V��������C�$9Č���s���T�53)dC�}-��d���`���6C�-�*��͉42�4�4CE�m�`C�	k�����ho�r�ñEH>��D&|��87��[5�5�T��8����ȓ>������r"�8+��GM��=��V]����3�t��pB�,'����&�>MsӬW.A���֥1�����r4��@��R��A�Hx���q��8��>�2��#��l��+6A��x�^�a5�γC3�`Gb�sbd�KE �}�P���*�DC�<1�PY�U�;|JH]�f.��7C�I#<�`�rȚ?�KA�F�*���"O"�ٲ�ײh��xCq��A[�!�"O*����*ɨh���\:Wl��"O�� ���mI�[5׀WF��x�"O�8���WL���K(=rDJ"O ]��˓�#�d����
�g1��J��'�ў"~�e�$2E^}�Ҁ�<�@�1A�P(�y"�O�K��PZwÓ9�����j\/�yB΀� $]��%�=^-Ԕ��)�y���wB&P�B��(�8Y�uƒ%�y�8h�h���P�W�QbE��y�W%QB	��(]I��!#��"�y�2���)�b7@�PX��L��yrL��L���ⱋ>iv��h�E�&�y�U$ܜ�yv�-��&�<��?ɘ'n�i��ዪc>�K7� Or,��'Z��x#l��B�>��n�~2}��'j2 B�d�-uh|*�a�!���'����D�F�m�hG����B�' ����OǪ�v#�<�"�B�'�T�g�Y�/����O� b]�'���(0n�x�Q"E��ma~�k���2�^$��h�#4�8�L�J�j��r"O�#����䩐j��y���S$"O�,C	�J�����E�����'"O��rv�V��p@'�s�l*4V��E{��T�U$+L��I�5h��,Ɛ E{�O���͙.
t;6��{�2��
�'��y-�$0��x`蘰}��	�'��!F�b�&��P��>nvRih�b�'���	�ƙ�X���WJJ���'!D���g�L�ZLa�%�J��I�'j��s��&%��es6�� >�|���hO?��D�:S �0��_�Bٞf��ȓ,p� CB�ɠ��,^.��ȓ@R̭X@DխG�`+�&�ktbmD{�Ot��)v.N&��V�W�u����'ء8��g�8�f�b�#cΐW�<QM��ai�,RW,L%���{�<��`L�i�R`;"gʎV���0t�<�S���B�c	1h�\9�#Fpx�4�'v �7I�0o�,�P�v,I!��k�<12���w�(�ӏU�F�D�
��o���ϓ�dH��~����Lզw�h��ȓCO����Ó:D=y�ʣ|'f,�ȓNr,�q��_��X ���
J�!��S�? �EVOX�0���b ��uv��R"O�X���0��D P��"]�5"O%��͛$#z}�S��9~��%"O�D�Ee�'`Pњ3(	�5u,<'"O��IGm��$�"�� �y	��2�"O��<mTY	1�x��
�"Ob9�D�*^^���c�0�eʂ"O�}���uu̐���C��S�"O�q���ۦF׸e�D��T6\�e�|��)�ME}� חd\��X@�I5�|C�ɔ$��)���:b�!+���p7�C䉟~T��W�.^����n2?��C�� dd��F�K.^d�P֮V��P��F�"�"W�
���(�s�ñs����	/��Y ,�n�x����T�ȓo�H�����N>�͙r�\�(L�i'�|����A�k@"ؚ�9��:��C�!E@|[c��b^h�{�ˋ�Q�x��d'�*�ԋ�*�X]g/�w����0�8H�sd�^�Pb� `�艆ȓ���sj��a����fOH!�ȓq��5���ƧyV�����2a�.���+f��h���R���/!��ȓg�2=�w \*����*8��t�ȓ#��H4 ؗ@֨qQcX�"��-�ȓ#�Ԑ�&iV�{�^�i�M�1q�؆����"JCv�Ε��c�V;^\�ȓ�	y�k��[ޤٹ���,�ȓl4R��GI��8{�E�-ED:��ȓ]m\�Y�J�B����F��ȓf���ԧ�H%�=)Q��M�2��ȓ=�40H�)�/�D!١挌Z�d1�ȓubX�-�!��Ȑ�TT�$م�#�mi�o.lhx�����m}�H�ȓM�^aG���3���xf`���&��ȓ\��bI9�t�b�č86䁇ȓkMܱ1bF٬.w� CJ:JM�e���v�yI�<Od��1�]�	�8��f�P�Hg%� 11��&˖�C�,��ȓR2j̑�l+b<đsHZ|�̆�<�z��#�()���`����1�ȓ<2�H��'�q��e��8p���!`"���(C ��� 8_H�r�)�$ã\ �LZ���L�ـk��yB�ޑm�� �cn��+��	�Њ ��yRfɣ:�*$��B�'V����-�y�C\?g(Pu2b��wȲ\��ϖ��?�'xJ�a��Ht`�!Kȍݴ�@�'����E�8P�E2��ˏ� Y��'}���A�E��`Q�(�:����'��M��I�2n?����[U^U�
�'i�:%��*�de�6(�3�E��'a��Ϗ�?t���vj� �2-��'��M���?^>\;Ueݵ��b�'M8�^!^�FU�'�z�f��'�|�`wEG-8�^�W��w02�B�'h�{��;	窭�d�l�ⴃ�'�.U��̌O�(��˘�4.�	
ϓ�O����N�bÔ��E%�>P����"O�H�5O�x��*4���VGHԃb�	R>yp���-0��f�1�<K��#D�Љ�c̚PM���c�@�p0|<��"D��Q���H�6��k�z6B���-D���D偡icb�� /)I�}���+��w���3� \��Sd�,�0��OW�|~"@��"O�����7��EH㨏�Pq�#�"O�	� J�����%�].Sa���'���C	(c��������B�;D��)��!*�d�q���t?��w*OX$���"Np�6�Y�\�q�`"O�0�� +���!�O�Ty��c�"O���V �o3u�7��Dy�Dr�*O(]A��9dj҂�	6���
�'��0"%�[=Νx�1;Y0�2�'���Y����k-8M��Mŷ<a���'�8�x�m�<��D�l�5�@\�ʓWT��@�x���Gƒ���]�ȓh�����&=�ru/�<t��ȓs���s��fh���>�i��QA�AY7.����E�â]�m=.Ԅ�/�kD(E�?��a��e�/��-��s�e`�ƞ��j���j�-i��ȓB��S"!	�,�����G�>?o~���09°�1t�6,���ضu�V��ȓ�v�*"�L�E�ZEɷ�]����ȓE��� �%��O&4��E$@0�����M�Ly�m	�	�
)�`��s̀��"4��2 [��t��1͍�b��ȓKĵb���qA��ѤkUF���W+��x�*
$ު��ݞVw�A��@�LQ�$�
8Cԍ�Y}���"O���J�V��	��
(2^�q@"O�󡭝+}>h�VN�>�H���"Op�!��N �@���,Y",��11�"O,e{�&�X#���JڵS�T�a1�'��Ih�r���#W�����8��C�	�"�����"tk>����K/��C�
7,�Y�R�-�
�Xf^�E�rC�I5l�(��J;�5��'^C�	5s���`�
[~eȂC˖PBC��.]��i���%}�H�	u�DMZ\B�8-*&�P�*�^�0��^^��=�'sZN�@
J9xeBL`��C6N����Qw(4���یGB���2NO��찆ȓs��0s-Y�8�� ��dG4N�ч�J�4��D\ ~8�g����-�ȓ$�밀�^p2��Ѓ���ȓNZڼ�@iܢ~�����]^�5��!뾍j']�-��{cS�*5��G�0�EB�(���ҶM�/7ՀT��Mk����/��;Kɹ$�� {��І�}=�����0Z�K�>����/C�$9s�^���Qᡄ�<UOf`��ph`�`�Ğa�yQ#�Y�� �'kB�X�d�$&���[�`H�j^���'�){�	�RBBa�nޅg���x�'+��B)ˤO�LТ���a+z	�'S:|  %á=�Z�A�W�V`�P�'�Fy�ӝ>��M� ���"O��B��b�:h"N�-�B�z "O`4q��q*�u  gƯ)�Y��"O�ca�L�g��0�֣J�.k�"O^���E8~��Cf �N�4�G"OR�ٱ/B�H<5zQg�8UJ�)�"Of�!�9<�|�:#�٘D�)؂"O��z����ٲ�A>�X��"O�mcl�{x�R��ع`�p*3"O�T�gղF�pm;�O�<�p��',!�� ���s�הq�Za)7�vT� C2"O �H�(/��%�F �|,3�"O��" 
d�K��O�b�����"O@`�q�%CsZ!6c��it�x!�"O
�����-<�QD�?XevtR�"O�M� c�!H6N��V
�7S:��T��D{��iý@���$$�0BH�ԃK�<W!���-���A�'6>?.����B�!�V4������$19L�|�!�D�	�8�v���+۲H ֪�+c�!��ܲ�jfF� s�@�����}!�΅* ��+Ti�â��@.x!��V�[��Q�pWk�%[!�Dׄ	�N}-���SN=&ۼa
�'�y��O�/
S�֬��	�'���G����@ҋ�Bl�
	�'O�\
4n�=0�iP�@�Uc�'���BÌ$�|T��(��0|`P��'ƺ8���;BP8�bT�#f:qP�'29�F�$[��:ٙf�B��
�'�ʤ�&#Շo@�� ZJ���
�'�L ���
��m��-NZ���9
�'����D.Ո(����� )��ib	�'na*4�3���s��kD��r�'Nذ�I�f�܁��KYOi��']\%2ҵj�*�{�)� �=��'5li��
�Z6����ޏA���q�'����Q$�,D2��'n�.��ݓ���/�z�!��@)P����1`�0�1�"O�A�%��<߼ ��@�W��$��"OX�9�݉Ϙ
я�7 �n��4"O��������z��`�"O8����6_<\�b�@پ���"O�,1`���*t�xt�C�`�!�"O0Y���=$��A�V#W�*��Ֆ|�P����K�
|2'MW�E�0sfJר84bʓ�0?) �5u��brj�3��8j�B	I�<�t���5��0�b�/9E䔰%�	L�<�*L�w�А��i��IX�V"\E�<�$N]�l��q��+O�
����^@�<���Q�d�:l˜}l숓&@�s��UyB�ONx`E؉W�Ȥ@��2hI�qsN>q
�'o(�0!�`*}��\�V/�I�'�a~bM�'�����A
-A楒En��hO"����\0���wo�� M�����$�!�䁔k��8[P��6)E(@���U6�!��0v�"���|>Z�� �{}Ȇ������/�fgإ�#�A+?
`I�ȓ<o@��b�u��@a��]#<:�t%���I�xV���iI�ZD� ��S>~B�ɯF�t0@D��7v�����N�g�>B䉼E�-A׍b�q���
��<B��e\`�s�˶a��Ҁb�7d�B�I�<7��Y�aX���Q�Z�C�	�X8��ӡC�\���6B��"��C�I_���%�B�de�[s�ԗZ�C�	OCL�B%W�(��R2M�,C��;@�X� ��i���[�-R�p��C�	�& `��指]Fe;Ŭ�[]hC�	W[�԰բ��+��k�B�)"�B䉀D�x`fϗ!�� ��=��C�q��I��Q-Pΰ����v\�B�	-[yx-�3��/>�e���ڤPoJB�	�a�,�M[♃U�Y�#$�Ox��� ��遊�
?���[�H"Τ�1��'�ў"~BC6,����O)��M���ͦ�y2-Q�b޸����M)X�@�Z�M��y���1qs`<��M��S@B�b!�\�y�%��lɀ �Ս�"I���ѧ�ݥ�y2Cw>X��썊Bڼ����
�yR�]�W�*���䎭?��Hg�=�?��R�ӫvhT��v̺@���y���3Y��i��	u�'r&0X@HJ�g�t8q���g�*5��'}*U���)S�%K�D߷^����
�'"�-�2�\O��p��N�O�=1
�'��Qm���	Q�B�K��8�*O:�=E�@ǫn�\�� Ƈ_���+����'�az"N@1�,�p3C���p����yR�D�M�:�I�3p�v@��y"D�;L��J��Q�}�h���ۙ�y򂌅nRą�t4	4m��y�E��5��y�+�:[*
��3����y���a� ���F�L���G�y�*�9\����!���ad���y��&�T@�(��/��ۢ-����?Q�'E�����^��!A��S6�����'���@�N�_7����a%� ���'�@�j�1U=�����>g��
�'�4A�Dg�G�1G�H�
d�b
�'P��SfI	!�&u�Q"��O_�T�	�'pe#1gV��)�G��Hr�9)	�'J����H�y���<����'	>B&(0 *�<�AC�)HFa�'ạ9�¤8v�|Ia�J3/�%S�'�-g �2���P�*��O���'2jl��W�$���g5���8�'
b��N6	���ǁ��*�z���'��9��H�-f8ef,X�8�lh�' b1��L.�����ҵ,%t��
�'���ӱ��,�r()R��+8<�J>���E�d#E�_�h�F��EG��'�T�d.�t�eE%c~�26��.��(D����霴x %A9���f$'D�����OK���G�
)�p	�c�#D���ӡ�J�Wb˂u,%��"D���3�#X�rɑ5)�LQ�p��4�O��!�bS�=� ��E"�/y�9��IX~"&�`�\@p.[&H&I	�y�hR)l����"�	-$+^�����$�y(ߙ��X[�*T#{� ��iB��y�b�>U\!�A�ɟ��4IDǆ��yBB8��m�u�@&uh�A
$���y�L�
� �y2�܉lք�bۭ��<A��$A�a��蓨�8��ke$J!>!��7IZD��%�)P��1tID!�D4u۾Q�mX)�,�Ѩ�;!�_!��[����UB�m?H�!�$ҥ@M���M�{��%/{�!�d�4Ra^@��m��(�ȡ�S���}!��L1g2�Qf��bN��3�+ܭ(�!��L(CG��#@�D�o�< &+W9�!���D�S�θ2��h�J�2;�!�
�Qf\!��^b���C#ǉ�!�DӘ-��%��*.] �{�oN�]!���B@���'�N$;�r���7*!�D��F�pb�	�g�*���B80�!�$*抉`�����|B�K,�{R�|B���qY�]"9�F��3��{+ўd��3� ��3�/X,Fuv���h�.�t��"O���q�
v^����cꎬ�C"O��J�� E��Y��Z� px�"O�Ik'ŏ�b�����1&�ҭ2"O�pg"�'a:8�b���1}�´��"O�9h�N�8g�^�i$�Һ��CB�'�ў"~Zw����љ@�	&7Yz�хi5�y��Oo��4c�:*h�m�&�7�y2%®��`J�<5Kޑsԭ���yBd�h��%t���x8�3/��y��v���P���V�H�B����y�8$����甪P0$�`�	 ��=��y�+�+?z:��+��BԾ91ѧ��y2�F'h�� ����<�[��(��>��Ob��H�oRrњ`"J�����g"O"e��c�x��c�5w��a"O޹��j��.<07�N�"��-x�"O"�%��h xb�0l�n�A�"O�L�3�0s��Q{V�l���i�`�'�a��D��)���%Úma���t"ʜ�yr�S:��Q�wo�k��"��I��yR�BM���f
�]�&�`'��y�� ��� �^�L���������y$�5GRD@��E�Da�UE��y2�P2~�d���Ӓ7�vY�E�Q��y��"��J����(,#��)�䓣hOq�%�����A�2Q`�1;�5��U����	1\N��p��M!5t�y٧ǐ'qQBB�	�[ZVq���иr�ʈ ֎NPJB�	Wޑ0DҬ6ޒD�G��[��B�	�e(ģ�N�������?<B�B�ɣQ$����b͟l��$Sw�I>VՊB䉸F_$��bY%Iu������u2tB�ɪ>}��eh�/;Uz���j��j�`�O��D?�6���k�L�e�c!��_+gT�� ���8?<���I�!��/�${ �K�_�Hp�q�!���)ٕ#r*(X�j�((v��t"O`p
!"�J&J ����&��+�"O�xp2��cF^�bOb���Y�\��՟h�?�}2e`��3ݰeK�M.�}Qa!�k�IZ�����y�[� X�70�S3E�4�y�H;i�H����.8*�}�@ �yR%�:6�r�[3ň(+�"r@���y�/� b*��̌�.l�����yҬ'`tV�L�-#�hGNL9�y"�!>����.E�2Dn`3G�1r!�$�c�	j�Y�6G�d��ΣB�!�P��wa�xQE�*"k}!�\4=�h�C�ܱv?ZXӂ�8l!�D�r,�"&�;n"��	_!�d�{H�$�R�>TxQ� 'oW!�dX������.1[~d��n7h!�$�*k�2<�7�U��x���ӭ%Q!�Q!6C�QD��M������}2!��:l�d�'��5r@��2�V!���)q0��4dǎpj�9r���-n!�$��O銙���|O����oR w�!�DF�d�N���ק2����j�!�d�+1\�Q�T��n�Q���.w]!�d�9HA0�(@e@�R����哪pX!���ò����H�MH:dϻ"�!�$ѭ*���a%����a����?�!��
�{^XiS�@
���r#7Xp!�� �=��N�^	���Tm�8�,��"OPmp�&Gxh��b%�Y���J�"O�mK�@܅w)f\ s�I�t�j��"O읠��71m&��G�88{\9hs"O��`m��f;؀k��( \l
"O(HA�-F�Y$\ᖪU1`AvBt"O�`q��#�`3ǈ^ x���jS"O>�KROРd��/�b}Z6G@�.!�:A�,�Ɉ81�O�f�!��:��0q�"�7d�	ǀC�	�*����M��05�-hC�I�^F���e�
f��ꔅٻSS�C�I�^������)�����G�f\lC�	�9Q����u�Y�� [�@C�ɰy�!�+-^���S4nR�e�C�	�ZՊ���#��戱��*eƴC��C�"�g_=T��zR�_��NB��n�PE!�G[�n�z����JB�ɠU:8)Ȁ"��Z����2,D.��B�ɐU��	H����s��d�4덐�C��a`����H.N���HBC��,K�2�F�U8`h���R�C�b#�(�̗�s�䁑�mѽw�0C䉛�� �7������� �z��B�v�1wB��6�X��� S5ŪB�	>M*���p��M� ���i�%j��B�:!?̂�ęA�,u��Ǌ�C�ɰy,�5*6hËB0m ���PI�B�I��!���U���%P�O�:��B�27�Da��#�[�d�h0mP�z}�B��+K�����[�R�rP���8 �B����4EFF��LYӇ
4%�B�ɿZ(���B*����ƥq�rB�	�s�~��& ܟ2AFu���^�M�fB�1"�d1z��ޓ0ze��.��B��/@������"x���W�f�B�q*��bլ�<|�9k%�2so�C�I�/��;�)U,v�Ѫ���_<�C�I�bd�r��*uS��B'_�NC�I=UD�c�)Z37���7�ޅ�ZB�I�#���jTI�=��T�e`[=،B䉧a�����E�detܲ�i�$�bB�I;�m�Peӌh�  ���E�6B�I6���A��1G���C�ʸJ�TC�I#a(h��u�R�}�>D��ǅ[�fC�ɨ)�H$�":�����!�C�	�"iԭ�&�7c�N'_���C��&x�^A4�͔y���@Ϣ~/zC䉖5��tK7��	��M"PB�B�,R���5 Gu �<�'��(V;0B䉀:��#�ZFy���Y�kg B��6 耀�CƇ.� �@�ڷe�B�I ^�D����)^#��hV�� {�B�	#�t �$̈�+j�HR$�6U3B�	�Cn�y�LO
GR���N�>=2FB�	�U�)`e ��\�a�P�^�u��B�I�u 2��^��x�Z�̝� ��B䉁fR�lq郴��YE��Q��B�Ɋ
1�̊�i�����Q�`[�C�	� �z��mG�Y����i%2��B�ɟ����A����,�$	5|�B�	�e�����FϤĹf(_�{g�B� N���Q@������ uEBB�I �.��&O�%����2�� 9�
B�)� ���ϭ�Pಯ[�B$�5"O�ɲP�+wp�<ږA����yK�"O4���E�2r�	I ���dC��'"O��9�'^'��ˀn�:{^�]re"O��	��M"Y�m�
�4\嶵k�"O�a'!R�l�0 B���mZ$"O4��)֊^��9�(Vl���"O��zS��u�X�ѣ�M�A�T�:�"O<�s�hR*)���Æ��!'D,`"O��0�O�*�uq����uf�� "O>�lZ/*<� V���"�"Ol���jM�T �P1�V�$"Oڭۢ˚�z�0�H�nI0�V�8�"O�$ r��sҒ�ِn�_r��3"O|X�A�(G�����^�����y�gCCr&U�ҥ̑o"`�����y"�L&(S^��R���fPJ�����0�y" Ġq����Ae�\3f�8q����y"fT7`�¤@�L[_��7�^��yh�
�`׍.�����N��y����(ÂH�fr���2|��mh�'Ƥ	P%L	<݌���]"r[����'a����f� Z&����dP�pdx��'�jA��A�錙��$uB����'M6���Ə�@0Q�� �#�t��'� @�.�5�}J�GɐN�ؽ�
�'L>A��U;BBtbp���v	49
�'��
!�ӧn ~Dl
�'�@�ڣ-��>�������z�= 	�'��a��
"y�蕊Я˥B�pdS�'��`���O�q���&���&F��'.$����M� � �G�$D"���'����	9�J�y�m�	��"�'TDy���O�!�OU����'����cĝ:C��LHG����	�'�0���ߍX�ɩ�k�r?jP��'N"�'U�.<�Ыk�	;�4���'��2���E��dbR,� .��1)�'Z�i�`�RF>��­ �'\bA*�'����f �d���q�\�����'�tB&ńwf�ʢ����2�'^VDX��݌Z�l����2�*�`	�'Dę��ᖎ��1!�Up�ݪ�'�L���C�X8�&l�Hi�	�',*%�g��1���sI?8�<1Q�'�6�*���%/�y��ʯ<��Q�
�'<t�$�� J���<�.P�
�'Z� B�63��*��vV�S�'�t@���H6aF�}ؑ��=�����'ΖhÖ�ڠu��-r���@)�'��(�@�Âp"�J���f���'���ʝ�'��{�:6�0M2�'S��*���`�"�blT?,����'Q��zU�U�7���8��0s�I;�'ޮ}�Ǆ�>l����ʯ'>a�
�'y� b���2A�Vp�v.L#Cf��'��)��@iI`�-���Q�'����D����"�B�X���`	�'�4�2�H^��;AeW�O)����'�N�#❦\��1���Z<$I#�'|NI�IX�]z��b�(Gt6�1�'c�t����By�LjA�M�=�|T�'��iڢN@� (���Ȓ3���Y�'��X1Ǩ����	�A���D��
��� ����aY05C�f���x4"O����w^B�+Pa�&  ��"Ob���
W�@��A�� }��)r�"O�`�%LUgE(��G�ӆ>��� "O��3��G��"\kE�&E��4��"O����Ȳw�P�����\�@(�%"O>�Yjނdg\@q���4}��!٦"OZ��/�9@��X����t"O��i]R������=���"E"O�H
��3*�̙p%�#U� Hx"OT|h�,�� �X	���Cɀ��\��F{���-ph��U&�!��T��2-�!�DV^u2�1#H�>�L0p�@@#�!���s�&�;f��f�L�%/�{�!���x� (��H�o�����Nĭ!���q�$9}J|�':@4�g@�������p�(��'�J ɒ�8O��t��G��c�6���4���A��@��!�?�xh3�LJ�",jL:D�,�A�Yʈ��an%d����c6D��C"��o:����Z,)�ps��>D�X1�؍cW(�"�Y;O ����0D�����][NT��m@hh�Ь�<�
��v�p��Z?�$�;��S>\qJ�G���h�6az���(C �[�H^5;�~C��4c,��%4��l��!�?5]R��ē���S�,fչ�#8 v@��`��m"C���q�CH�9a>*�s�b�@�DB�	?u` jE6_1
���C&�.B�'Z�D�T���m��щ��BdT0����h�t�>%?�"ǍA�>�ҽؐiZ�{+D�U�<�O��'v
�W�� <p����J6-�d���'�Pt��/`n�8���E5�L\���d8�'~����'�
G�	@Rc)�|��ȓ_�1��7n�4��IF�A��܆�,�©����~L�%z�`_G䍆ȓ��ȑ"��p
���c♄ȓb�e�p*�%&��f�Gd&0�ȓol�ͱ��J
t� j�KϹ���c��?,Oڬ���X�!8aU(A8vԴ�b�"O�,`"*�,�2�b! �1h�!�K�_�<�Q�Q�=OL|S�+]h�ў|��ӄ�zt��e�	fГ�DʀC䉱8'��+��F��*@BF�r�T��?�{R�	�'7�ppRN=�0<�0��%	BC� {Q�x8��g�܍�DZ�L���n�a}��G5{x*�B�#��X���<�K�ؖ'Z8�˶��(��TO����c�@��y2ʉ�������@�  ��(ިO0"�d@�0��0��"Kr��p���e�<�Q.ؐ\{��b�"Xs��h��W�<�bJ�()X0(q0,�4��X�SR�<y��	�V�f��J�T�Q�C�v�<i�ȗ5$��!�e�!�0%��aSo�<yt�ٮ�v���X�q�J�:b.�l�<��� � ��I�i�����h�N�<i���,2r]�tC߷5Ah�����t�<�����L�2���_ͼ�%fKX}"�)�'4Z����*���
�f�!,	����[t0�z�鉌0[de2�ě�r�u�=Yۓ{=\Z�j�"j@�3�ĕ�)���M���R:I�#�	ǧn�q"/�~�<�����B��N`H,��@�$0�Շ�K�`�Ѱ�)kp���m�.*3Ь��	\�'�8$���J�^(���
X�j%8�O�-�O� A@��!@�*P�RDȥO
�43O���J�S�Ov،�Q8��#5�6v%����'����B�7$�$����v=*�(OJ��$HQ�b>�@�ݣ!*���`�8ud��<�O�`�'W@����/YV	)%�	2���;��yy��'}x ��Z+.}9�`�x��Y�¼i[���O���H��)��u�׫�w@��z�'$�$����5$�1Ȧ"�@�"@�,�(O?�$�/�Ɂ
H�
{fY����?!���g0ڨ1�@<i8��Cʻ)���=O�i��&?�"ƣL��U"O~�@����EM�5)"�M��9�$�O���o�g?I�.ǲgB�������T��8���9�y���2Ҋ�`0(G�NZ �	7`#��$�<�H>���ɬl�d�y�G�KBPDsc�r�C�	r�e�EǗ�l� ����
ѧ�ē�p>�'�
SK�d�Q�P�C�ƞu8��$��'njI��d�%�f�I�^e{`�m�<yT'�(Qgx�"'+2Ƹ<����h�'� �F�4���3�h���`�N x�E(���yrÀ8�L�z���8S���m,�y��Va�T|�Ѡ'Q
���u����y�kX�/��i�̑#NA%��6��D.�OX�VZ<f�. ������P��'��	� ?>�B�+	d8��`�⎧�rC�	#Zb�ѳ�B�9(�����F�0"=���T?=s�B<Q����(}���P��"��F���'*JV]�U�#m�ƅx����( �H���F{r䐋`�Ё�'��=6+��ɥ
��HO��$�MSmX3E\�_�q�U �#,�!��hT+�H��{p�pwOX$��hD�ԩ+}!��zU�	 �b�ZG�S2�yr�B�PV6��c[(�Vl��A�y�l� %D��#ӌ8"X���O��ybJR�$
�9,�&���V����%�O� �\�O�h$3D�L�
i*�Hc"O���Ξ�G5 �����,t_x���"O�D��͝<]f�R�o�>1�R��"O�%���A�m12o��`08a�'Y��OLԨTM̕kJ��!N__��@�"O���'bD$s�tS��D�(f�s"O �r%�53��1ɖ�H)f$��"O�)b�	� |�`�P�u`��X�"O��{�$�
H�b��a�à2?v%Ӈ"O���	��gi�ۅő�mB�8���s����j�E�4�D�CR��sC�m!��M�oj�b�rY� pW⇤�!�Z$��Ձ߭@���p@ԡ~�a}ҕ>�E(�I�
�(�o^�h�s����?�/O����(l�x��/16�d�r��:]�!�DWPC.��#-h(��֪N�D&!�$�v���ۃ��\�"]�	��IhX��&
Y&�P<� ��j\���e+!D��Q�O@jA�pF#>-R�{�h)D�sugM8�lR�˄;&�h�H$4��C#�,U�����S�p�lC�h
E�<�¥�B n���$�>A�5#Cc�~x�TExB-\&U�͎�&*�,Z!����y�V�c�MX�Q5j��mS��y�� 8�9b�\�,? =�����xr�ii�i���߻>��mc��I1&X�6Y������'�v�>�w�ۉP�	�B�гP�@����'LO��#zyr��L�19�`*`@U�:!�'t����	�?��xJ�ܳ$��,S ���D{J~� �����{���W�ΌN��H��"O��p��� ��A�-�TyV�R��	}�'��ɳD��5@5H!Q�dis �N;�B�	�g�V	B������,�%h�B��rI�]#��N1)/X4�+�.d�B�w8�Y	�A�e�L,��F�X"C�ɉT/��Z�M�E,��j��"<q?�S���Y�IP���gR!P����T"���yR�F;/v|`�Z�_�*��7�=�y��)�	z�����X�Q�U[b[0��ȓK69!p�"��!�s��M��%��R����R��$�^�� �*a~�W�P���7
�xth�l+d`�c$D�L���:B��h�G��2��5S�$0��{���';wҥ:U
S	\zp0�"�:��ȓ6��4`�d֜\[��-��'����J������p}��;� O�"��w���1eU$f%4�Cר�J<���ȓ1p�D�5���+��%;:�B&"OI�e*
(7���$υW&��#�"O�8"S�&��р�0A����u�6D�X8��%U��PR7��I���S	5D�,r�J>"*  e���礜o3D��u�B�t]�,ID
<#*f cqa,D���WN6����U��/T@F$y�+,D�<d��)V���*uC��u��ɦe(D�`Z�I�
&@��5�m޵+�h'D��
T�R�_��)#C��3������$D����H�0uziƃ^_��Q�3�$D�Da�*I �H�2f�F�{�~m�B%"D��xE��C��qD�@C���Q�:D�����	B�|3v�
���Y��8D�c����%j��҄:h�A�$6D���� ��(QhU�w 5E�� �5D�����X��NF�`iz���'D�ԛ�&�6d���9���j+ qj J8D����F�agJ�ԫ�]���Ja)8D�����Wak���I��7D��sv�L�y�| �_#Dt�"�M6D�|�ԍ�0*�v��ě�Ql���63D���%̞ R���vE�9a�@���1D���w�� k�`��f@W*3��,�'1D�Ȫ1/J!�q�2�Ӡ}w����3D�PqQ��$S���x�+�-Zo�0c�,7D�����<V�Pi0��d<�dF #D��(��]�!��3��x:Jx !D���w��8�LR��9����<~�`�p
��]�#
 LOt��6MB/t2���I�� 	Z�BT"O��* ��2 �ɴo`x�"OEp-P�R��@�l{^���"Of�J�-ѽ�Z�CT[�[�i��"O��b("��Jc�_&P+qkP"O�Ջ��V3_�c���z3"O�`�n�o��U��d�7��8`"O�p{��@'H��́hy�؉"O����(>$���ϐ�F�$ڑ"O�i��W):�3�O\�1�6���"Ol�C��"K�q�7nJ�
���"O�ɐ��U�2QP���D�$��6"ObP�gL�u���3NBxvv0�a"O��c65"��Ȋ�PTy��"O�0V,$A���Q��=^^nĲC"O*M�匯Q��Y'�VATq��"O����X�b�jhQ@$�,X�l��"O� ~�ۥ`ƘF��a��	4$`��E"O�؃�?zt�t�6�D0@�"O�4��R�a�2!8�T�}�@�R"O�D��H� ����S�C��$q"O┐���i���K��Ǔ/ߠ��#"O�J3"�3Bhl��Rn��n�"p�"O��p�O�Y��ã �>&�Źp"O4�r��Xy-�I��6;�P�"On �e�N7k^e{`ΡO'xXK"O��DB��:�Pggø0K��S�"OB��r��H H;�L�+�J�"ON�� -"אm�b����*U��"O�@2W��gT)3PԳH_�}	�"Or��D��5�J`�5
�+f9"`�"O|��p�ɒA�<�P�V�W<lX�"O,�	]���l�1�s&��p"O$%�(S�k�ҹ�MZ�ic�0�"Opm��Y\�;��S7o�h(�"O����A����"G)�)~y���"O.Uڶ�m.�����g��E"O.����Z�k��X�2F�N�h��"O��`��3�d����Η9�b4c�"O�U�0*K��\8Q�dI�A�,���"O>��F�*kDڱ � �:YxhM�V"O��iạ̇̄
�"���ܴfh��a�"O^U���%4�ᆛ�[Z�Rt"O���&�g$� s���R�$�{"O>5�&&} hu��L,2�j�`'"O�����X��U���G����$"O\X�6�zW�-�R�P[�"%�b"O��C�M��1O,�
�I y���S�"O��EFN�$��&FPT�x��T"Of����M/��c��0�H�Q�"Ox�4nƧc�¸�C��8�l��@"O��� �U�"�@$����B�:1"O���n&F�h�h�>v�朲�"Oܙa��9z�0$�g�X*�	@"O4E	��L#�6aY��T:Eʶ"O���KȨ[Ѩ��3��m\��v"O�xh$�'K�(�+f�R���"O,��a��F����(9<��0"O�m�S�
-Me� #2#(��U"O��
�ER�x @�Ԗ�7퉠�@q���S��!D�](x*Z5���/+��B�	5md�%	bn;���i��P�f�!�`̡��0}���'�`X2,B�\-��J��[��U�'�
�+�n�<d�@\Y�f֛d�*�+�"�B�[��ĔWm`�YV�",O-���m��H[�.������'*m�ECW~� r�CĚh��x�ǐ�y���O��TԠ��
O�ة��˽E�qy���8����T�dD�)�2yGη,�8��-�S�sx�I��:A��[��6=HB�	��r�U��]j�SFH�,u{�q�G]��ðֹd��Z�'���v�M~n���&�ѿ]>1���^�,��UKw�Sz�<!�ތs�Z��4�)ADp`����:R���0w�J��Z��7Il�oڽ℩�)S]ܓ"�P�pT��%|�@:c!�,nz����I�c*��F��8��=YB�"��s�`P�h)� *|�5��a�WL88Eo#�����tJ��j��H8O8W�1OJ4:B��S�
 g� �Z�J�����#�D,�9`���	WqFLI#�@�XD�0��<�!�F=Z�&����Qe���a��{�n��u��+m��IՆOcf�JG>\�2��!�?��3�t���$Y�CC�PeeK�~P���-2D����(4~Æ)*���)\���a��(��t�g�##��I�t�ő�5zɐZ`b/�I�bPf�"3n�\�n�HE�����L�<t��!#�'d�+��]��8���N�3n
�y�"��*�b�����`C&љA#��	ӓP�X��&�	U7Vu���[
��'�j��DA��v�A�
v΀s�J�+O:�T�P� PH�u�	����reV�!s�4"O�D���K�o�$��sN�
az&1[��H'Z#�Ę	��=��8����g�X���n��d�b}(-k�1�l�́{�А�!�x R��'��t�Q�R��E�oάn�>��掟��]`E��+����6�n���ѡ�i�A� �^�_�qO�������u�!V8s���J��n�'��-��/��]�؉��j��<�����	̞�\�(�IBL��ٻ)�7&���i��'� �n=�p=11��0w�(M���C�b5�d"�BlyM�
є��ɪ�\䫕�\�H�vh��O����@kĽ^��j�v�N���L�$�IS"ON�s�;i:�V�Ѵ8����#T=3p�K�fӍb�Y�S�ً_>D�o"u�p��[�����/�yG,,���A1+��Hn�h�Ǣ���?� �	)cj!�N���@}���ӑ
%��(�旰��#q�7J):�@�j� �P��3�Ji���|��2��!9B�S+E�n9;'ϐ��O�ز�ȼL��Ŭ\�=@�u�P�̝u���{!)�-59q	f%�2;���H4b���ʲ(����Ĕp�Q��N��bc�`@eO��2��(Z�����Q85$\}��IL#��"I�*$�x�㑰J.�tfH�N�t���wh<���0df��x�.ǌO>��

F�'�Zu�& Ԝc��D{?�`�+)�	�sCv(����+q9@T�B(�.$!���}���R(R�O]H�'K'_L�7��(�:-Ä�d�p��<AǤ�n_H����j��]�M�d�<���]8.@���N{�0y��:@
���%���R��M���<c�� 5����4,�UZ�4����v���1)��-A<�!M�30�l�JQkB�g�N���b=�"��64�|�R.Hl���!���%�x%��,�I�x�ɩ��wF�xC�-��M��Ii萺G����@�8O��B�	�r|�5�˘t	�|Ȇ"M����J�A=]��G�B�$���(��I5 ���	�aO�IJv�Ih��C䉺o��6f´-ٖ�
C�
�$�����J��ji>|�2��1��z���)��)�E�Ȁf$DX�p�H��p=) ��\> SrLܢ�M;Wl�>��PFF)x;�	�V��v�<9![�ݨ!r�(Ӡ|�:�Ӷq�N�����l�i0|G����6~��ڂ%�8��[�ٶ�y2I����q�I�(n�^�iG���x9�!�]$���'�>�I,�����N�_�t�q��{�C�_�L�'���~YhP׬Y����D.y��|A�K��=�d�k����ɐ��do���0>� �^�^$��*dJ`�¾kM(�r�GZɖ%��Z���$!V4K � � ��N�QDy�	�[� �F�t��#`�L+S!^�FN���ȹ�y"O˿|@1��9H��xiq���y�E�E(n�j\��m���y�嘗bW��*㋃�Mf
�k�)��y������c�E�,�H���f֭�yBm��K��|�`('5V��h� �y��̀~2VD1��?#�@r�]����'C�r��K1B�4 ��m��L>�S,թN�$�IV|=)g!g<�s���;tP(�U�yB\�*�◂E�"p�C�G �R��D�.p-v!PϓEn衔�e��(��\�E��U��ԣv5�CƁ�j�!��U�^|ظЂC�
�]�w�^H<����?���(�OL�f�\��3l�Dy�#�>5�E2Q&O�a��A��5q=��~zDM�5 ]& cI'k��P���G�<��*���Lx&H�#e�2��C�����0nχa��-Rvi�
:h�h&?1zV�x�Ѫl�X�wfP�%��j ����?ك�Q���=�ɸ�NɩN��<A��$R�Zh�@l��螀���A��@���~e@9yD`-q�V*��U�^ >�?���W���;�(M<T�t��4 ޛS�M9�
�p6i��k�6{����&�1$�̋b���:�[��BqЉ��<��]&o���.�,_��x�G`½��c?�$�D�$����%CL޵��.4D��yw�S�+6$�	��W�Pc��$-�tA4]��Bs~t�+U&��CԌ��~�#M<Y%�L�X�� *1�SQ�б:Q+�m<QhB{.�J'�������9oC&�
�g(vw�p1JM�#L���m���
�EÒ����@���IIz4���_qD�
ۮ=�4��!R�A}��� ��U�ޑ10"Oȍ��B" /�L	�eQ3f.)�"O.@0�Ϙ��bd[U#I�li�@�E"O� f����׆1��+�W�U�c5"O�Q[6l�"#�a�n��C\t�rw�'Y��ˁ����ɵz�$����}˲��d�	�6C�ɴ3��r����S�*=@�)O$L`�b�8P���Ne�\+��S)p��a`P�_7�ҁB�&�BB��=�6����
t7���b*:d�K`�S=���e��!��L����������ا,�\@���/4���U�U�)�B�zo�uN�^L��1"�)�6a��D���f�$~dڠ��̓&_���M�}n�L�%Z��	�>��1/W�؂$�vO(h�B�Ie�*pZī��8p�O:J邏O�,HG!�9L༽i�"�f���Q��R< ��t!Z�+�Xm��g+R�jQ���B�|`Ȉ���v�T��B��'< D��>�gϟ+e�Q9B�N_��� �`h<a5$���<�+���,8���@�-TG^)�Ў���T��
�{4��s�ٯD��H�AɅ�z�牯E��T�w�	��~�ΓGk
�B3�0\��д���S�"Oȵ�#AY�t� �A*(�R�	���**�X�!� ����
ܩ��Bjx��ɀQc��
�'�Tx�fW?i��!�	X�fv.t��oDr�O,|��Y�4#7�Ͷeݾ4�5��&9:��!D�\�'�H|@��)��'8���C:D����|m�Z��ț �����9D��(�@/`�z%k��P�yP�0�E D��#f+O�?��ip�ѳ2 (D�V�!D��ÕJ�*�8����"�H��+?D���B*�1dn���C�ub�y�6�=D���`F4[d��Pc�
���p�<D�$�F�R!Z,ڥ�4�F=1,RPZ7,)D����-�N�� ��!T��3�	'D��bSK�n��  ��<K���$D�<���:A�J<(�ȑ)_`����m1T�P�t�"�d��F� Z���"OΩp$B�(g����x���"O�XqeN9]5�Eq C������"O@�8U�(q[xm�_9(�� #"O�$[�B�7?��01v$W@��Piv"O���f��	9kzy���O�x��"Od��#��a`Ri�b�;N��uqW"OH��#dJ$u̰S�R
�
9h�"O��!�R�q�,x���La�� �`"O����ę%Ot �d^�E��U�W"OV��$�4�r���Y�BK׌6�!��,�4*V*�*U�Z�Re�+�!�dk����D٩�6liG�A�h!�d��L����q���h�pp*�"λg�!�$ķLt�P����{��5 �=	�!�D\�tnB�A�:L3��ZN��!�D�5q�Z���ݯ 5���EN�R�!�䋺	̠XJU�J�d2�y����b�!򄍼G&yZEN֥B2D�o�e!�D�s�y�*�/w���YA���h)!��ΌX����ŏ�LA�]�U��!D���g�Ɩ7���^�t�2��U/z!�dߝCK��i�)�<�hm�č��!��v�1�$g/U�̐U%V�|�!�d�2dCD@���	,e\rhr�KA+�!�DC�J�J��ɪ[Db�2S
E	�!�d��9����V�JHr��c��]�!����Hf�$.I������+�!�V�b��R���\"Hx��iJ�k!�$��rY�QI0/���(C/H!�,sπ�)�@E(M������,n!�B]}�E���xZ�Y)���b�!�� &qS��̸��� $�<Ŏq�s"O=phρc}bU��A3m,m��"O �f�&*�}��)Bl�1�"O 1��LT`�t�5l�J4�%"O�x�*P�X��]"�b��I�Ř�"O0��b�X�eX�9c�Z
�lt��"O"���Ŭ&��B��T��9��"Ot��7.�p��X�I
~pp\Y"O"Y���ʒv�(��!� q��q"Or�J e�3z7��V��Ujx�j"O:��4.��a��<�b�ŭ0���"O���L�A�$S��CV�!a"O�AbZ-PX82W�S�J�ؼF"O�2p��n̻�
�1�| �"O\�9aꎩd�`����
��)"OX��ɏ�{M�ZA��;���P�"O�`�f�LC�1�Y�}�^%
1"O���lD�؄��!W2"���`"O$�'�P�q�$Q���R�ĩw"O0��fK�NՖ��f��@��JT"O��BA*O4��#l���d�;�"O�8"HQ(_�: B��P6r���E"O�)�h�)Z�@L���(+�Z�"OZ�����sp���T�����X�"O�I�'K�@�F�[rc\7[�Ԡ�"O���p�I2�@)$�.`���U"O��QD�I!T}��^�$�:鳣"O���qjS�:0��6�Z�\����"OL032-�!
DiA���6�\��#"O<�k�b��K���0� 'SO����"O��� 9�z!2a 
�67j@3P"O�1��o0~RS	�c�|��"O`-��锫4(.Ջ`g�*M�$�"O��91!�=~�������N�f��"O��@�׏	���*S�+���T"O�%�c��U��QP!AؠV��\@�"Or���*��w�	�$"4�"O���Y����RNE {��"O�{FK�i����®��:��#F"O��Ro�]���� �
3�H"O���L���P(���56�f	�"O"]Ck�%�L1y��)$�2�ل"O<�v ��\\���9��S"O����h;��9(�L2���[�"Ozy@�h��j�D�`���9g"O�@��*��$8�A(�.�m�H��#"O�B7斩Io8��-��s،b�"O��:v�_�T�ġ����+�n�sG"O����*���A2P�^-��"O��)���2<�hsD`Đ9�L�[T"O����=`wp����B$w��Y�d"OX-�CL�7#���A�X#.ǒm�"Ov��d�����2��/#��q"OLdJ꒳d϶d��F�5���6"O�к&+h��;��D0&�.p%"O���UΏ�j>��_�ɱ�ՔN�ў<���9>k�>���!Po������;����*1D��6�۴*�����C�6��ɸ�Jkӄy�eXz��O?7�����EK<!%��Y�{(!�,k�V�)�%�8
x��3$ӧD����).g�i�O�0=y��]-^w�Xq�Y>u�}k���G8��Q���6� [w+������V��9�fhS�K(q�!�D��BH�a�a.E"V��q�$�ΑR��a8����V �'E@��f!d`�'?��;q`����H�b="��]7G#�Մ�S�? ��ɠkSt���h"ǔ�k���ɳc��*ag
�&uD��O�`���B;Ubf ��y�m�qwQ#���40w������p<id��"����cקlGvh��L f[�)H�	C̾��ǨW<S�J��:rI4(6��D�azb.ű
�J\+&�*�E+����dP1Q�S��>�܍h��҈i��i�<y1��_)�(��P zЌtd �d��C�ɓd��H�����D�B8�b��i]d)��&`Baq�J#/��d��Fg��P����@�	�-5�21GV�@5���t��V��/��"�35M2�xgf'&��\"��V�
o�v�S��gi2)	�K����\�H��,k�i)�={�vm2����,��͑�Q�qp��?��)и$ڪ$���G�AO��I�/ީ\�V�H����o/@��^;���-O��h E��z��z��Gd�|y��V�Z�|���)��XvTqR�=E�<!�`�8[��'M���TH�G���[q�5 x:��Q�B6@)����'+bL*�I2'òA@�/�,.a܅J��%q�J=KR��������F�*.n6��fL�םJ}��e��c���\��p��o��:���˧�>�O��S4�7~z����cO8e�gɱ�X���0�a�� |�}ax��Sn���'���)�CH1�|��$��d�`p
���T�#�> �e��gH���id�^w����U��&�3tn294x��O2%�𯙢u��u�	�dm�:�`U l)dL��	��0�n��'�Vذp��L`ɧ� G� OfL��G�̣^*�0ZC��6tP�b�Y�Fw|��O��`��D��pA��h�8�@�d�4}y�HGl�8��O�1��hC�|JeȐ:�
HįI�O�:`C�r�<	�� �q�f\���U�ܰrMτS� l!���l;�A�'��XD�,O�( �Vm>���l_�-���5"O
}�rO���\�%�we���P�+�4����N')VZ�H�!<O\�	�f
�B�x��π'�P����'���c 	�.-�Y#��P�A�\���EF�:^�����w�:q�',�qS�jӞ Ȉ�UI�/&����{Fגz�u��Z�T��I���G�	%�p�'��_{�t!G[��y2��!������:%�=�7,+D�T�q�
X8[�¡[�'[R=F�,O��1�@,2��N]�yE:���"OhոF�
d�kt�+p>t��֍9gD�6gкC�ڱ
דS��(�T��w�t��S���&\O@�J1G^+��E�!
w��1��:0Fp {V���]~Dp�"O�D��@����Q�=��d�Bvu��	S�Ox�>e���]_�}2g���S���2D�6D�������TSA'� J�QRD��(w�1�J4��	o��~�éI�rY�%��0G01�g\��y2�T�r� i�I��c`r�@Ff�
�?qG�e�
�&'lO��9����B�:��w抱x���AD�'V���N#C�Bb�A����+�!d�������yR YjrJl!���$������(OȘqp`٘ꈟ��që8,�B��$遃�N���"O��bg_ċR������A`"O�E��̙��Uk����GLԩS�"O 	ʒ� ��������f�xR�"O��kN[� �F�[ōҟ;�}�`"O*A�wgQr3*�A���?t��m�"O�4P��  u�(u��'I�} 7o�to�pG
"Q�:|�
Qq�q��'W|P�G�&"&��2�N�4��'Vx@�$,�>F�Q�#�G�/�.x�$N��X���K� $=Sz$�H�&O��yB��c�(49q�K��2)2�k����O�e�� ,{l��hP/+|M�Qf�yP�L4O��xh�v��/02��'N����]C:4��Fа;k���.OT�P�D�����J��#��-+W�ő��O������!LB��F�ī3���;D��+����E�p�@�N[�<�y�hX�4�<b�2⾵����(�������K<A"͔7qS��)$��n��4��&�g��tjR��4\�!��@ʲR�45Z�Ě) �� ��X�0R rB��*��'�\1t�Еw�ҥ��(��U��J�����@]�*7jO�FXE
��H�7]����-}�z�����!h��pc�ɼ�xB�O��@#�-o���p큄��D�-�$��RC�����91������D-t0�գ�F+5_�0
2�y�(�0k����a�..��)����>G�<��m͝�b��"�x���KL~��<��,t>�;�郳`=&,�2.|5���[n��1�Jn͌X`��Q-\�$�A�Y�A��ȆL�6X�����<� r�!2��*sf��`���l1&�'9�ĉ��Jl�����]b�H���ޠ������ѢmT*,%%ZK�<Y�d`�]����	.Ļ�#�@�<!�2��a�iB���	`��W}�<e3ghB!Z�GK�]� Ly�<�o̍~����N/%0P�I�������	nD�'q�)Y�%=v������1pt	��'X�Ā�L�5	�(�V�J)t��`��yB�J�v��t�ƥL�O��y�/�f�Q3J�S����'�L��O�<��My� ��s�$��4�\��%�+O�ջ�2�3}�B�cd,Ōqr4�'�����x��vtP��ՎL.4w �sunV:Q\$!*�G��[���bS�'���q� �V�8�Q#��a`0\XϓS�𑣇�gj>HH�'�,�rf�]:&�*�;�mQ�^�a�'r>�!�)U>!�J�������zJ>��������ӈ��%��!'~��p��ڕu>*��F"Oؙ8��5|#~� O�� H�@���U4DA�R�(1TBD�g�d��|���C��XMf�R� �s%��D�!�蕁��H�uKd�ҰD*A<l�P��]���i�&�O���w�O�P2��B�?��@"��'Q6��c��<��T2�3O�Y�`�1Z$�a�D� s�+�"O�����\b�0��OǱ6f
���<��ݾY�HG����Pt���T�׾s7ƕ��]�y�D�Z�4"�@��^'\}B/[�$bN��e�!�ۭ�(��ɪN�㢋_(��Bq
�i#�C�	�T��a2�*΢F���BmS�[�TB�ɗo��QVb׺Bz�CҬR�'�8B䉒_{�]PT�L�!�ܴ��ǍG��C�|&��y��Y�vD� S���C� AA�T�� �= .�z�H�e*tC�I#%���k�1W�Ӌ�60NC��3�"��ř���!��2{C��%+�eʱ�C7X`&$�^Y�B�	����W�@�i� t����(C�B�	��	
�ǘ:m��������B�	�˾�90j�	i��i �"R;"�B��	&}X\��?<��@B����B�	N�t�n�/b�Q���i��ȓr�hl�e�B"G�R8��l���ɇȓ{N����*O�ab���Ԅ�ȓ3A`���:����L-����9B|9�&�D9���g�I;�*���Z�ĐסZt��O[���ª���%��oȀ���/��x��^ՠ���K��
Q�U	@]���ȓ��C$�_�!�L�A�#4�D��!��(wi	�Y�΀Y���xɸ(�ȓ-�
]�T �	���Vڹ|fZ��ȓ)*DB��G
.M�5�̶;�b��ȓh����O;4��D�$0z\��ޢ��`���c�Zq�a͙�GX���p��ud.�UE�99��XY��}�� ����c!$(��9Q���ȓhL��c�4�R}�!�_8�Ze�ȓ?)JE��θ:Um�:놀�cB�����S�M(Tڸ���Ɍ���K�E=[�O=o�C�6���h�Io�6���')+/�C�I�aVv̘0cǁ@~uZQ��0M7zC�+/
Hl�TN�����صJabC�	�.�����ͤW�R����{�B�	#r`��Kd�_�e��D�&I��:��C�U�%�[�.4Ա��L%xuC�]��7�
l�A�VY�t�Ny��'�L}y�����{�B[�'T� P��Q��0�v�OE���JE�H�%�>P�zb����� ��Y�F�Vst<�w����7��]?���>��4E�=�0|Z�E�XG������=-,��Ɯ�-�ˈ_�T����%2���)§��dŇ�Q��e�!�[�"(`���3RW~��6c��p0�b9���Yi>%���,F`Ԍ�$�;(���sF�M���jf��Y@�f'ő]}�,&>�}é�00�|��b�
�nh �8%�ڗ0���Y������,k^a�4��;DNXb,Ѣ�J̀��3w��	"E ����M�g��S�'��PQUh=)d&\�0��Y��m�Bz�M)#��)��O�3}�*P���q�[��f5#w�Z.�?	������"~e&٣#�܌�U��l���ɀPg�92
�'g
\��"�
���}j�*7H��y"�U��()0)��"�0�$E��y�ǈ�%���� �@�f� "B��y���t�hibB��:�n�b�l��y�o\�S�� �d`��Z�Ζ��y��I&O�QC�T�PD!�W$�yriP�Rkp�#PO�GoȤP�^��y�ŎW6�ÆE8c꩘s���y���|E"�'f�����yRȃ9(jf���K�ؕ����ybl�,����2I�-�jY��c�Py�'�-j�$=ۗMQ�o�$qz�@�<��ҸJ��]kfJ�>C��Љ�T�<���owv�X'f��#�pٖ�P�<AR�+/��v�[�'H��Z�Q�<)���0Lʹ%��eW�U�P*6D�N�<Qu�Cc%n�I7%��-=r9�nFa�<��X�2�-�S�%��)j��Q`�<�ы�R���(Q�CL�	ԃ�Y�<�2J��i��t$��
Oi�511��U�<�$ �%J�l�v�	���*�]�<�a@�@����+:�L�0'*�d�<Q���7F�P]৹B9�e�Ŋ1f�B�	�ag<}�%�]����#�D�I|�B�	/j��#c6Yu6� ��0�B�8�Lܛ�$G���������O̒B䉣;�b|�s�@�q�tt�E�A>h��B�I7D�\��#�J�^� ��C<.��B�I1d,��@�V�MvL8�uc��.{�B��.8$�� ���En(���$Ҁ��C�I*"Z��@i�}{"�X�AN#�C䉜JyȀ��h��RS8x����\�B�ɖ	����2p�e� 	3?�C�I Ӧm����iNܭk�%�	-��C䉓� �`�Iȹ��v �C��"T���`O�<�����[^M�C䉔D}�i��\<"�XH�vB[1��C�I9I`����J�g[�x�)!:�C��2��L#�`]�MB͡��
r��C�I�Y2+F��^�8SAF�)V:��'m�A�NE	�x��h�H��H��'f�����L�8�	cCP�E�.5C�'��q�����eF� 0R�:*_z���')�h�!�J
93����n� c���'���0m�m��y�@�V���y�'���KehO�3朹��F:; 9A�'���T�K8*FXD�҆,v���'���eW�H���bC邷T��3
�'+rx�"�)�����T ���r�'4�2���l�(I+6�ߍ_����'U��Y�a[:!@�+YT����'���3�@^��k����`A	�'�6�����O|�t��;�1��'-�ɠ/�%8�yP�nW�;�<���'�cSD�w��\%ޔ0e������ �͊A@�T�ƨ8CBT$67�`�"O�s���)R�j�� оa")
0"OL-��5 �J��N�
=��JC"O��b��%p�����"#�Qp"OA��GK�0�ݐ���zl�"O�hr$�<0i�U�H<["�X�"Oڌ��J1�0B��$ZP��"O<i�	@�>T�e�(at���y盇jLt���� ��h
0���y�N�d��pY� SG�v:gA )�y��q�J陲�
�2�^�����y"g��^���˘�W�)P���yb�¦���A���N]>��A�م�y�(B3��,*���>*��A��y"�_ a`��{�DI=V�����Q��y�J��3L�0�BY�`��a˜�y�ճ!\�(����2G��yB�Ϳ�y������,)dh�1֨�sRÝ�y��	 �%a�@H�, h\Af�0�y���M��P��	�8$�����y�aD�E�f�80BB�6j��K
�y�&�7hܤ ��e����pxW� 	�yR`�,��4���+
0��e�_��y2�ˊ~"V<����U���9E�(�y"/�$H��R�U� �����y�P�46�PAifI�L�0@E�ȓV����G��d�f��m��p\�!�Ũ�en�*b��?[E&9��uV���g�(@��rS��N�<�ȓ	P��"�]&F��-���֤z�D	�ȓDHp,	�  �s!�i��FHyz�8�ȓs)�t*�%��$K��Xc���G<��VkF�H"�`%����ȓl~,i��n�
�b�4�ˆ>;)�ȓ�&Yq�#�lA�@H+�$�&��ȓ	U\s1(�IQ �+�·{��}��goJ!��`@�F�I��Ǳ'"�B剐g�"i{dO�iִt1a�& æB�I\@H�4 ��,�XhrS.7�B�	�6#b��NA�f�P1萴.>�B��R���*��Ƞ$�7D�]f�B�	<���V�DY;���ӛw�xB�@�(�&ַkՂ��A P/Y�lB�əQX$K�cT?$���-��B�I�e�jl�W�W�#����V�T�t}�B�	�g���ꔧB;�Ї�*��B�I=etba{2c�Y�"�q hR���B�I.Z$��zv��$/��6�.<�C�ɯL�D�4�C�j�5*���DA`	�'�$l)�nȶK�E#�! tdY�	�'��\8��ɟG�f��Kt��	�'}�5z�'�*k N���N�2�
 �	�'�,=�OD�#��VP�SdP��	�'~����aI���f��R궜"
�'`ZEN[��^uL�2-��'�0��b[�n)L̐%���>�h�z�'+������8�H50��<XD��'����A��-u���/## *@Z�'����e��:ԭ�+��$�t�>D��{6�D-��|�cmũs���Bb:D��yP�Uv��@�"�ƎiP��+D���͇c�V]R�K�$VXF|�2�*D�T��A�gT!q��_�~�:�	s$D���	S86�f�afd�&pM�2c/D�� �|h��<8����KS�u�:�1 "OjMs���\cd,���!?��Q "O���Ѧ[�r���T)��|pg"O���BZ�(�PZ��84�@"Oܠʷ"$j��5ڒ��ܐ��"O�8q�Ɂ3d��x�����Iq"Ol�Æ�� @�$,A�w�$�"O\�I���9�p4��J( �6�;`"Or�y�Gˍ{�$x����H�N-9�"O���3A�,
��)A&:	��p5"OV�3JR�H`����G�Ľ,�y�JZ�6P���̵L�>��%��yB
]cqj�"s��Z���eH�B�<sZ$4�̍��ʝ�K���P"O��Q�_�Q�p�EW���� �"O֝����?C�j������@H�!"O:\�'��.�����->@k�"O���Y	]@�H0q�!z��8`�"Ol� D��!)hu l[f
@Q"ObIRp��f���hw	��Q����"O�E!&Y%��9R��>�d�@4"Oplsѧ	�. t���g��?Ƣ�ò"O��q��v�21��֊9MD���"O&)0�5 f!⤣�0L�Mj�"O���4�� ��0h���J6����"O4����ΦJa����[=)>��"O���A�ݜh��$�#�ۛ/	H-�S"O�yS�
Bn~<5����sd��d"Ox���
M����t�IM6���"O��Iec[��\���IK>����"O��`R�G�<��L�G��;���a"Of�×�P2-p]��H@{{�m�'"O��0�-ޝtЄ�ѡ��_hƐ
�"O���J�+�r�bN���)J�"O(�ÏS�^|���&�e���q"ONYЁ��h���֎��
J��"Op�K��F=cpL�Tl�h]R� �"OȘb��{5,1�M͍/3���'IN��s�N2lP����M�:��#	�'��h5��9H��y��<W�Pa�'_��9�/�0�t��<��
�'����"Ӗa�,hK��[�C>:�3
�'�(�#D+Y�]���0>� x!
�'��8�"�<i4&��I�i#�@	�']d�P@E�m(����R�L��'�j��QC��w����A�*M��S�'+"��p�-E%��+Q�U�5�:��'g��a7F��g8Erqك:T�%�'`��jw�
#P�&๠��.k�'�0�H��	�*�n��#�VeY�'�JYZ�F�tX�H
����t �'y~l{�'�39;�a��P�V\r��	�'�� ��*~���*THĄl^��'\n$r0kĩ\����X,"H`�'���3����N1M�*x��7D��;Ƌƙ�zIj��Ǩ#M�ݳ#�6D�\04(�8��-�A���<���t�9D�Сg�meX9�Jc��,�ӭ��y ��cb
�#K�<��� P$�y�K����"��EJԙ�r�Ҷ�y�b@�[�v� �I@�B8 �����y�GΫ\���"F�H Ȭs�I��y"iX�b��d�����>���.ʛ�yR"ԝe��	���E�����C��y
� ������d�p�'��1R��x�"Of���+�A3PY A퓭_��7"O,���	E�j�$H�E%�5/.5��"O��d��q���Pd��#E aP"Oj���Ӏ. �4�w�7'��a�"OJ}��BM��p����P�_�q��"O��T-�EY ��<z�<�U"O 3�c� ^|�Agk&KΪL�"O����@+2\IF�@�k��u:�"O�%�w'
:����2
v��l{�"O�-��Y0�S�Jh�`"O����GT"^�P�2Í�3A����b"O��{�g��:�&�y��ʦ����*O�y��JG���b/G'H�Q�'�ܠ6g�F�b��%X1Z���'g^�
K.'�*�`ܘ=���K�'�f�bI|�<���Թk� !�'������s��İ�E�^gB�*
�'����f�d�"0amY����	�'�bպ�KU��B�X2���V�Fl�
�'�jx�  ���   �  C  �  �  �*  w6  *B  �M  iY  e  q  K|  3�  �  �  �  �  ]�  ��  �  ]�  ��  ��  ��  �  O�  ��  V�  ��  J�  � � , � h �! '( ;2 	9 L? [G �M wT �Z �` �c  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+q��62\���<4�d5h��'�B�'���'	�'/�'�B�'��x�.Z ?܎Yf��0d�tx��'��'���'�"�'��'���'�nY�5��B��0��g��ծ�pW�'l��'C�'���'���'���'b��i���8��}��dK�� �C�'1��'W��'�B�'���'���'?�%�����غs�9
lk��'A��'l��'B�'��' "�'O���ek�92�lu���D�+��'�"�'\�'���'��'B�'�n$Q&菷U�~�
�"��]x#�'���'��'u��'�r�'���'� �H�N$!��y;�Ã+K�f�0�'���'$��'dR�'���'���'�Fx-Q@�蒠�6/X��o
�?���?i��?Y���?Y��?���?�Po�^}��� �	\V�p�'F��?��?���?Q���?���?!���?auj+2��!� :D�|Hʗ��!�?	���?���?y��?���?���?y��ь�����/�&8CTtꖢH��?����?Y��?����6��O����O��DB(Hc���$��[��$�E/U��b���O����OX���Ov���O�!lZڟ��	�P��H���L�!�"��~�-O���<�|�'��7m�?3�p�)2N�&g]��*ϓ�Zφu����,�ݴ�����'�"nlr�q%�E)-`�����:�r�'hr��iw���|bA�O��)�t u=#�h���	W4+���<�����4ڧk���j���=3�6[��
b�,Z'�ie�,��yb�i�ڦ�ݛ,���d�!&�;$,A�;�R��	ΟDΓ���	�^46m`�t�E`�p��%]���2��t�P�p 2Mm�����'.�8bG�C�8 z��;1I�(R�'E�O�I�M;�˛C�Fmv��'֏el�C��:6\ui����>����?�'<�ɯF�*Iɇ��<Yެ��Zn��?���><�ޠ�|��+�Oܠ��l��|���B�`([ LK�2O�0�.O��?E��'Lt��ӯT�L����L�6LI��y,|��,𘟌�ݴ������V,ws��c!�ΗM�k��� �y2�'�r�'o��b�iD���|2'�O��!���N����!�6)����Gb��My�O��'.B�'���_�v� 1��k�/2��GM!n��I��M��aɐ�?���?�M~�<�t�*phR/�J���ӋU�>\�`_�x��4��6J9��	?K��S�%��"�L�;��C$$fx� ��= ��:'h0DrA"ŕ���<��*�I�rd�,�d�>F#�����fM�Iן��	����i>U�'�v6ّ��$��c�b����ѳp��h��Ъ%����Z̦)�?ѕS�T�޴c����n��b�bR?#�V@Zc��&r�^x�f(�6)h�7m+?Q�)��
���)���s�=�f"�|�Pn��hR�鷢�K��ן���ʟ��I����|����B】2`�M��O+ �&�3���?y�Z�F���~%���MsI>��_#L�x��Lՙn~=j6b6
��'K�6��ɦ�/a���mZs~�!P�FO����	$����A��TǄ�U%�ݟ�@Y��4��4� ���O��R�'X`��Y��X��C,�M>��$�O˓�����,*2�'��P>5�n�|Ot$�rd(y�8����9?1sU�`�I̦]�O>�O��ucr��X��3b��)G�D���&u�@(��P;�����{S��Oα�+O�T�4�Q� ������W�K�~���O>�D�O���	�<�T�i%��d�Q^S�D�"B�^H����M��'D26-+�Ɋ���g��,aG�֏%dݫ��ɮ|	�{�FҦ���4xɰh�ٴ��dhVѓ����S�?P���e
�g�Q;3��p����۴���O�D�O����O���|R�ݻsA�\S�@BE%�kB
�vK<k���ʟ $?��ɓ�MϻD��tH��(I'����S�f�I��'����$���tET?ԛ�=O*D`��͖7NF�k�>���S5O�h��$:�?1ᣩ<A��i��i>9��>G���JeF�}꘡R0�S������,����'��7�í3�`���Ot�DS�7���v�6 �Ed��?2~$����Ol�n��Ms$�x�/&|��Y�
�r��H�:���'{����FQZ
�O�T��#3��dQ0�?��G�	�dTc���*d����'�̫�?����?)��?Ɏ���O�mY�ڥ�p�z"����8��Ԍ�O�Mo�p�p��矠��4���y���c���׉wTP�[3���y�EoӘ�n��M��f ��Mk�O��³Fş�s��.�R���Z�y:�$�N�,˓O�f]��S͟�������|��#� ~l,���Բ#Z����Eyrco�N0�&$�O$��O���d�?!>��'G!�Uh$!J(��'� 7�Y릭�L<�|��F��'�2YC�%ۆ�"��͚���ȁh_~�׼5=��I&>I�I9�M�)O���,M00Ҝ3���#MdT	b�O��D�O��$�O�ɪ<���i�j	q�'wZŲ�$�W�n�jqh�,�rl�`�'7�6�3�	����D��͹ٴ<����7���8��G�Z�XT�"�z�. ��i��\�Xp`OD�n �iq�)�D�~�� ��c��PZ9V|��*A9bT�0�0?O
���Oh�d�O��D�O.���Y�� K`��b�X]� �C��Z�Vr��$�O����}	�ln>��������Wy¬L�zr��TOاW��Yd�\>��6m�<iC�i��7=���A�q�
�de��KG�P�A�p�R�ߌ/�h�1 gؑe� %
�+���?���s����uڟ>���O��8B��� ���3v�se�\(6v��d�O�˓&%Z����d�Oxm��?=i��Z��]Nm@�d�$	o���OH*�t�X����ūݴ��O�̄1��!G��BJ�_xP"�̝C}Du��A���D�ٺ/�6�T��?��Ӽ˕�S�\BI���e8X��Ȕ��?a��?I���?ͧ�?�����Pצc�j�����*�B2TV��d�6������ܟ<����]�<z�4%�@-�"�7B5z�C�L�7)��!R��i�P6MA�$7�.?Q���7S6v�i2���N>�HD���j�2�A��յl��6�<���?���?A��?!*��e�(/
����
~�4���[Ǧ��!��JL^Y�	Ɵ���/���i>i�i�%��([;ь����%"�Z��@U��MU�i�z7��<�|���1�M�'_"�"�oQ�k`x�IV��e���<��h�5!���_��������4�'�T��d��?�%��!#�D ���'�r�'rY�X�ش/��Q��?��N.\:�cڎx�a�%�,c��	�OL��?a.O��lZ�Mŵi��	�@��h�e�)5A�KuL��V�>?�抩�9���	W~�jmݕx��'U�4�I�x�P�`&S*�l�CQiշ#;�����P�	񟈗��)�O���O0TҴ�����c͌R��%AQ�O �l?Q8|��	����	ş�����w�~�Ɇ�oj6e� �ԒR�:���'�j6M��3ݴN�ߴ��D��.�@yJ��6x�d��e�V,��f� i4���E�O:�ĄҦ����t�'��'��'R ��*k{�U:��""�����V�Y�4!�(��(Ȼ�?Y����"��.��E?<^jla�*�J��<2ѩA�y}���'ɾ6M��	X�43��>Qr��P`�Ւ���fR~���,r�H�(?I2�K"Z��������'�8Ȋb��gh}Ү�5�*Hڥ�'���'������_���4|t��*�dZf�
1M��i�h-�v����x]H�/ۛ��$�ty"�'��fk�J!���	"��=S�#G�uw���K(m��7*?�"D\�C���+�$ehݙ��2ar�}pc��>%XȘw�Yj�D�ǟ���ڟ����Ii�'�\��(��|�T.@�7�҄p���?q��R����_��D�'JB7�5��ݽ\�����a��`����Qמ0��'�<��4h��O�.�
2�i�d�5��KeoǉBe�l�F�I�.�rŐ�I-N��TK�h�
�'�\��'��'c�'gd1R��6C���%��Iה��@�'��_��s�4.z-��?Y����)]9��	��+���"jIo�������O�7�Q_�|�Ƭ5Vh]q&:ȼ,���9n�U�ЀV�'r����d��`�U�|�
C� V����O��ج�vb�1�I͟��	៴�)�iy2�k�� ;���P, hq��ԦO����LK��I��M���j�>)ƷiR��1#��#"i*��U�L����!/|�R�mZ4-�n�L~��̶"D(<��n�)P6Z��Q��W�c�Dڴ%X�J*��<���?!���?����?!/����F�`��� A�Yl�.GB�7��x��D�O~��/�9O��nz���`S:L�3�!�#Po��P���MK±i�NO1�d9B��t���ɢ!,�z4(��ZJ*XӲ�����ɩG�@]�%�'�x%�L����'w�x�t��x?>��w��$h��!�f�'=��'�Y�X�4q�����?���Y��r��œ9XVM�RÌ�a�������<Q��?�I<q���)�2���E��ZuiANA~��J�咑��W��OP���	�W��L��x#�RQ�H5�.���#C�^��'���'����QEP�^���!ݥ;�b�! ܟ�ڴh�
��,O(oZL�Ӽ����_�H��ȌK:)�7��<�׾i����`���Ѧ@~� �H�(hWn�2��`DE��I�E(��i�x��d*������ON���O����O��D��/�� �Ac�$��I����wJ6ʓG�&N�"��ԟ�&?a�	�x�~��Q�O'�:��0c߻G���ʯO")m�*�?aL<�|j�l�6���� ��^�N���,<i SȈ����Z�� ���)�<�OʓV����9d����R�F�n���(��?I���?���|�+O�DovCF��	u�Q������$jɜp��	,�Mۉ��<����?��44� ���E[3v�X�;���&���M�M;�O�8"��?�r֌4���� �[���<!)����G]�p� ��s?OL���O��$�Ob���O��?{�HZ�Q,�C� H�H�&/�py�'��7M
�5���M�M>9⁓�
���C�y�RG�#�'g 6�Vܟ��S�H�R7M#?	⁍E�b��p�S�my>��
�`k�d����OՑL>�,O&�D�O����Op1�d�V�ߐ�S�!h��{w��O\�$�<1��ib� ���'o��'s�S�/7DX #��#����]�hF�$�I&�M���' �����O��``��<�F���ȓt��	e(	
���Sb��m��	�?�3�'��a&�pr§��u�x���D�\�|(#�#�����ğ4���b>!�'�6�Š����a��B�@��#��Ox��̦��?��S� �ٴv;���S��*,�C�ľcȬғ�iM2�E�(��5O���O�A}�t ����)� �p��ǳ?�����ϖE�79O|ʓ�?1���?����?����)G�|��S�XL"��R7v1
tl��?b�t�I˟��L�'|՛�we�P�� [l_v�I��B�0��RR�o�ioԟ<���OAli�p�i��D��f ���'����U��y��ě�z{�e���{�O���|���!�y�E(Ѻ^т�)�M�P$�İ��?����?1/O�oX"ެ�I����	��vT �F13k��*<p���?��^��	�4Rg���'��43�hLQ��//1�\H�E�!�\^N��M�Q2p��|����OB����+ E�C��w�֑�w�
P�����?��?���h����س7��8�.�G��H�2/�����¦Ey�Ĉ��d����M���w��9;��F�$ᢱ����,����'l6-��M�I+�t�mZK~b�H�,����ӵC���e!F7�ҹAĊ/4�'�|�Z��Sן ����D�	֟ �4��?@�ʅГ�N/}�l��[_y��g�Jmj� �O����O\����$ҋ�,٠�@�*o6�[U���s2���'�T7m�����ɿ�H��Mj�햣0 �C�O�TW�C�C�u+r8£��$+B��?�F�c�Oyb���v@�c ��,���AI�1	3r�'���'��Oe��MC����<�׾A�RUB���}�������y�,t�@㟀J�O�oڋ�M�Ǿi�d�'\�İzׇ����c�ƖZ��&���[ª�5Q������f�p�f�:��1�Um�#$�f?O����O���O����Oz�?�h�!V)=�P�g�B�(F�����$��6�MÕ�z~�feӸ�O:5S4��N|pU���ڒO�@qw�s≕�M����&��(�&��hj�MR">Z��s%�(�\�2p�_ 6���(b�'X�m$�Д��4�'��'���Gg��K��@�%`�mTh��v�'a_���۴S����'2U>�He݆	[@�)WU�P�H��!�8?	�^�4��4*��A"�?�s�A0|���QW�2{،ht��09�,8��>u���|"a��O�1JN>Q�	���	7�X�iv�B��ܼ�?Y��?���?�|/O�(n�0Y� ��R��V��(�I��	��y��-���<�I��M�����>��i[�E0��'_��9�h[�/�M`���O7���06-5?�rȂ�z��I݀��3@9>qRbH�,��H)���2n��<��?����?���?�*�"]��	~�!��_t���������� ��Ο0�Iԟ@&?=�I��M�;:� B��?g\1Be��W���MC0�'���O�И���i$�D�Vq��K���3R("�7�ǐ/o��0��([�v��O�ʓ�?���~�ViA�^Na�"���<E�Qy���?q���?I*O�qm�4�2��	ҟ�	y�.���G	,`;�H�+L�<�?	�S�(��4hR�x�Q
'J$�����҈�3e�<���JA�у��ؐ~8ғ�����y8@�$Ƙ`�ʍH���ud��E!8
���O��$�O��D �'�?���)��rgĔ y~��HF���?A�i�LX`_�|�޴���yW��0'VF����
�fV1=OR��; ����O�6��H��7�<?9�fG�1JL���uf`h叞�EO\���H+�,EM>�,OD���Op���O�$�OW�:К�b��Htl⨚ŤJ9������jd�����ߟ(&?���0rh�
��ݠ�&T �m�0C��b�O��lZ�?�H<�|z2��G��\�0��*8�����'w6U��H���$�3~��ȡ��'=<�O��x�D��� v��|�Ы?n��H����?a���?���|�(O�~(@��F�'$r��V���kfᐟx?�u�'�p7�7�� ���F�}���M�!B�sG�]���F���R ӭ �bŉ۴��J��H�h�'o�v��|��N�~x�h�FO47�6̻FFW/L�D�OD���O���OD��)�S,�I���#�l��TfL�����џ�����M�fS�D�i��O%1F�<A�\���"_�C� �R��/�M�����D���}ћV��0J҅�x��i#��ʠstQ10Έ�K�����'c�&�������'b�'a�8J���.���㐻kpsv,Tk�$�fT�\9�4��@1�OG�'c���wt=Ӧ��9$՚�{堚�v&���'krW�؀ܴ)��]�l�O$��˒�OH����.�)+��ذ��/�,��4�Z�iq���GZ���S�i�b�_{�ɂ0�By ɟ�|��I0$��.Y?���	ԟd��ݟ��)�Nyr�d�D���K�yD }�^-������bΰ�H��6��_my��i�n���啂#���'�ȂF�Ĺ�Hf�Ȱnڕ~Z��m��<��,��!����>4�-OpM{w՜A%�1`A�٠�e��>OX��?����?���?������Z�4�Ha!��);0�d@S���um� ]�-�	D���?9�O	���yW�74�bܓ|�f� �G�`��7�矀�'~�O,���OjPz��ik�dʢ��1�#�ܿK�� $Ɔi���Eb����Hr�O���?��^Ą��rf�Y���1�O�S�p�b��?��?�/O��lڊLGp0������I/��BU�SW���h��ًa?V�?�\�DaݴJ��x�hI)zB|ɲ$D>;o���č��yR�'r!�#..`@�\1\����S�2�T�l���]�r�������a�^�i%Tܟ��	�����՟(D���'��x�Ó 5# �A�8/JA���'�7��r�J�l�f�4��4a�BX=E`D���X�0����O*6MO����ش,Op�4�y�'�4D d�?�Q	� t5�A�9)bR�;p��`>���<����?9���?!���?�SɅ�Ls$4:ъˡCC
��G����dC�����ߟ���䟄$?�I$4hp	p⨗�e2�#�n�#w?���O�`lZ��?iO<�'���'N�Ct�S���!v-���[7禈r/O�dX��U>�?9"�4�D�<Y�Y�(�@i eꝔF��}�!߲�?Y��?����?�'���T���: F�㟼QP*��%��HA���Q�r�۟�ڴ��'���}�����O6M��w�X�(�,_<u>X�CM�R:Ќ��mv���	՟0CE,��Yly�Om��;)�D�	�9H�A���y��'9r�'���'>B��1]n�����0�R���jXd/p��?�Ķi�Dq�O�" i�*�O�����`ܴ�æ������!x�I��M˒�i��4��Rz�f<O$��ظS��)�DZ�5�uh&�X>$}�d2s��?��@4�d�<���?)��?�v� �X����U�ߦx� rH�?�������(T���ϟ�Oo�䣁Ş��V ��΃�P<��O��''T6�QߦA�O<�On�����0���1��w.n���(� x�&��4�` �?,|�O�ɗC\0+��왶�;�N�� e�O��d�O���O1�xʓ]?��Х����2�'W�^p�F�(ܜiP�X�P:ٴ��'�^�N̛��mZ`8� �@6ȝ�U�ףI��7��˦qz���}�'^:Ga��?����d�s�J3�:��׭��zR�8O���?I��?���?�������~�Z ��%q�iB �V�lںs��y���`�Ie�S��I���k5�h��P�7�1R澡Y����&R��s��%�b>���D¦��9+�+��I� �B7MwK�,�@�%�P��O��yO>�(O���O8}p�jD�_�z�`KȔR\���(�Ol��O��D�<QP�ih�`�EU����+�
u��_�_��Q ��I.`<��?��\�t�ڴ"����8��0�D�±ŏ�Z𶕨�FF'���'.���wl��,D�b>��'N���	�$)j��צt|�e�(ɲ&������������z�O�R!I�.&�xZ�(E�r�z���׶(�!f�>ĀD��O��DOЦi�?�;FBIb��6!�x;d�@�����Oj7m�)n�R6'?	T�^�	�����HVX���հb��ÔC0&���N>�,O����O$�d�O����Ot8�7*�x˒�	��|r�ϭ<y��i`�Ԃ�U�\��V�S۟Ƞ`ɐ82n�B�zn���IK��d Ӧي����|�����P	_�Y����2�"u
�d�7 ���N���Г}_�p�c<>�O��L����3��ʇa0�������?����?���|�.O
qm�)N�vp�ɝc�rQ:��܊F���DHDʨ��	��M���<����?!�4+�J�jA�����p��� V121cǫ�*�M˞'
�)FfH����9l��?I��W,\��iG)~���T�Q�>��şl�	��<��˟���|�'Q'��H�ܩN�.pУ�O�O��D3���?���">�6��:����'��7�(��[�"b��zc��28@�AvN1,��$���4zƛ��O��ca�i���O��%&
a�j�k�䙫x|�r�ǆ�C��H���N�O�ʓ�?��?��G�VM񑊘=�T�+���!�~����?q)O�oQ2���˟8��P�Da��K�h�GGP�r�P�X��F���d�b}�f�����Q�)���K�@쪙�������n/X��$>���+O�ɇ��?Ao&���T�X��'�3��$��&ԌFz�d�OX�$�O��<�$�i��!B��Z_<8�@�h�'gS�T�r�'%07m(����DB�Eې`�,]�IK��^�T8��\��Mۅ�iB� �v�i���/\��-S��O2�)�Δ��
L�7%�ش�΃}��mϓ��D�O����O��d�O\�ĸ|Z凁�Y��#qŅ�?��A:�d�K:���|&��'7��O��ޟ��i�qYCJN9:xx�Z�3YF��?�۴�?a�O�O�4����i~�J�U=���Fj�� ��l	����Ro�\����t�O���|���C������ :`n��,�r>�#��?���?9(O\�m�0j
�	����Ɍ\�7+�X�+����І�N��$
���M �iG0O&�����?>��tj%�;��xC7O���I�lP:���H�0����?�r��'o�I�I�cJ�EQ��(89�����*$�����ܟ�I�4��k�O��l��@�㎨{l����R7l��l��xA�O��D�ʦ��?�;��U0��_>a� ��� �:����?!ߴM	�v

������xJ������+v�٩�&R<$�Rɔ9D=<Y$�(����'���'��'���`
�k���Ń] L�|a�[�\1�4h��x��?Y�����<�(�>����N�/y$P�dI�V��	��M���i��O1�����AI���{F/��x!S@�4`BU����"� �/n")BP��|yҋΧ8����@��� � �D�
0�R�'�r�' �O��Ɏ�M��![�?��牦6"G��+=�:�l���?���i��O8�'�D7�P�U��4߬���_�&�`T��GW\��qZ��MK�'���J�?1�E�S���d��Z���4�``��C�<`&�4
$ӻ{�$�O����Of��V���'���\������@�p�Bod�I`�������M���A~� k�T�Ol)�Q
���(�H�EG�p0`��R�	0�M�ױ��tΉ~ɛv���R҆4� zXb� �zy��:����5�\@�d��%�?ٗ'9��<�'�?���?Qwj	��aPa��(p5X)`��%�?�������)�%��̟������OMJ��]��u�Q�j)�UJ�Odp�'��7����l&��'j��qA2��2y܈Y��	z|�ē�"[&��J���4��t)�"픓O��@��a�H������x�%����O����O ���O1�8ʓ|z�&-�-�, Jĝ�88F@�יyB<D���'A�ee�&���ODtl�%s���7�9�h`��*�{gh�+��M��Ύ�M��O���K���ɩ<)���-tN,��5��w�}ps	��<a/Of���O|���OJ�$�O��'#��iP���,Kv�p3oMI��ѓ�if�ђ%�'m��'D��yҏ|��Ζ� 2l+	^�iP����C�4,umZ�?�O<�|R�):�MK�'Z�m�¯��FF���G!��O `��'�
�k�%Y۟�K`�|�U���ܟ�D٪q��r�� ���*�g����쟤��hy��t��X���OH�d�O�)v��
-��=:�M�?�m��&;�����Ė˦�Y����O���ԅV["@�&��<Ge&H�'�D@&�B�m:��g���g�՟L���'��ӆ�W@ubus�׵h���Bg�'���'Mb�'��>��e��D��a�)�"�C:=�m�	��MSf�2������?ͻ�˥@�*�8u���)C�ځϓ|	�FA�O�7
K�\7M(?���)L���i:���@�h
�?W6�r6ǆ Kk��K>Q.O����O����ON���O�T�@<��,h��=|��q��f�<9�iDƅ�D�'@��'p�OAR̲Ek��԰1�Ĉ�'�'4z��?��6��O(O1��A�S" �VKf ��!�a��d�aH�,bn��n�<���!$���U8����DC%G�����K�8��#�P�)N����O��D�Ol�4������)��'�/�%&<i�쵢���T�	�0
����@}BgyӒ\����1�ZB
�h��<(�~p��JǄP��o~�E��`��+�O�W ��YX�#�/[P���R��ɿ�y��'���'�r�'���F7x=S���:�)���>T�˓�?��i!~���O���k�p�O�)�!B��>��I�ꂆ�H:`$\B��ǟ ��ffKo��s
�� ��A<Z�� 3Hy��ҥ��
M�6�$ל����D�O��$�O���H0Q  �2���OeTHB �L�T����O��,��V�ڎ R�Iȟ��O�|2�Fތ[Ќ�zB�^)Q���1�O~9�'ո7���'��'u�;Ƈ��c�r�@�УL��%c�0<V�|��#��4��@���\��O�8���I�8"I����q� ����O��d�O���O1�f�&
�V��&{���p��
�-$�����$	���'ODy��㟼�O�En��d�4�cC6j�n�jV��f�@Q���M{#G� �M��O1�Ș��
B�<Q��>d<B�;s�5����<Y.O
��OD��O����Oʧpf�q�d�ƷcՂ�[�D�/myN��&�i����F�'n�'��OlR+n��ΌG�"��SW
c�t�ԋF9�mZ��M���x��$B֬G���4Op��Kވ_�|	h6שy�Pa�d=O� ��T �?�w+5��<�'�?1�e��3O :���*~>��
�
=�?Y���?�������¦}�5E�����IџHj�'�#I�Ґ`uIՃ�.��d��e�
��I䟼nځ�� �~�d��6����K,p@��'i 8���]A\6����d��Ο���'bR&a�5�*-�w�N�>�P0a��':��'���'-�>��k5ʔ���YO���Ȕ� 4����$�M�Sm���?���ޛ��4���`-���Ց�,�:4���4Or�nZ�M˄�i�ؑ�!�i|�	't��-���O��y�/�s@$Y)	˼X�q�q�\�	|y�O�'���'_��)0�B�H0HB�њ�˔*5���/�MK�,���?I���?AL~��b�i��� !,�"���i�xy�[���428��� �4�|����\�f��?K^n��k�$�$�jiq6T��D��\�e��/�b��m�Zy2-S���IX0/F�3�d�	sj:���'���'��O��	<�MK@%Ή�?ae�4j#(�� [l}�vj�<���i��O���' �6�To��yXB,�k�1]���f		b����	����'"�i�F���?�Zf����w?�`�ή�R�S`M�$޵�'��'�r�'jR�'����*�G�A���;��Q�dV������O�d�Ov�n�6u�p�O���'��I�u�Zh	�|�����J��~�BO<!@�i,V6��^e0�y�R�I���Z��+~&��Q�*����F!H�YJ4�b��'�~�'�Ȗ'���'���'9����Ö8Xn&���4��:��''�S�̨ٴ~�D����?Y����3l�^��<2���X�JW�� �����Uj�����|���<�h\`T!�X22��>~�X��I�;q;������sy�O�ȵ�	���''�qs��F�PJ��4���p��'�2�'�b���O����M3�LM�0v�ms�A�*J`�)r�C:K��1++O`m�S��/J����M����j�A���/Z��TA�I�b��6.c�J����n���I��L���N���
pybg֥"L�k���^u���q��ybR����۟���ϟ��I۟��O�1����x(����H���4Ix���� �O<�d�OT��:������9Eq`��#DI�)��L�׉P�d�T�������|J�'��֬�+�M㘧� ��	t�E$��h���$*zHY�;OPDG��?��=�$�<a���?�ǔ�&��A�H�.����.O�?����?y���dH��%h��W۟���������P+U���k����� Ȗ�Z��7��I�Mk�iP�V�9�mľi@<�%���P�J���m����^D���A�� ����C�O�;�XF\̡��J1 1Ȩ�6�F`�[���?����?����h�n�DU�\D5s�d-@v@\+�F���䦑s�3?)ֶii�O�.<���3b�P:Kj���ЯJ�W��$B���Sߴu,��'_�gT�61O��$�!��`8���,�G�H2�u!QK4�~����2���<�'�?����?1��?��S�k+���r$�*��cw���D���[�}������|%?�+a�����d�78�ti���^�'S.O��v��($��i����I�A�6��fg���c��O��A�/� l��	?U��9��'��u$�0�'%�ૄ+ٴģ��e�����'���'B���X�� �46�Q���T����"�'T�b�Ұh�/`�TA�$��$K}�%q� }��Ħ�;�"�J��9BUQr�ɴ�S����n�^~&�N�D���.h1�G��.��E�Q�M=�|�h�A�yb�'�B�'&"�'�2�	@-Z����%Ѻ�K�o�?1n���O������$�m>��&�MK>����κ�Ҍ�
�{��O��xx%����4���m|��ڴ��:��`kө<���aa.�� �։���:�?�c2�D�<����?���?���I6r}J'�ԳL�8�H߁�?�����d�-�Ӈ՟x�	˟4�O?
���끰����`M��O��':7���4$��'l��M�g/X9���j��Sr�
i��I�*Jv`�կO���4��<��9X�Op�J��H8d!��rO��G��O���OL��O1� ���*H._B ���l�%�>��h��U���T�h��4��'�>��CX1�H�ڦ-���5�ԍ�6�i�L7M�p7M$?�g�2٨��#��D�=�p�8U���M�`$#��y�Z����˟���ퟔ���H�O�L��g*\�;�*�c㠍0����N|�<�eg�O���O����d�ݦ�]�f��q�ȇ:
J
5���\�@|�شJ�&�"���R��7�b��8��Br0�$��y"��Q(j�t(�C� I��`�Vy�O:� �"��q`ę�`��,�\1�'���'}�Z���ܴp�������?���N�Y�ꌻ;z�p���N�66&�q�"��>YӺi7�6-�j≹{�X��7�җS|���1�� $������9u.^�"~А
�B+?��$F������?����,�R�01��q��I<�?����?	��?Ɉ�)�O�u�b��	ʦp��>\�L:7`�O�mڒ~�x���ٟP��4���~�g��<�d��p4^��#���<Y�i��6��O�dKw-`Ӭ�u4r��i�����jʑI�P�
��g��TP��^9����4�h�D�O��d�O���=Ub\�"�d��R"�{W�8%'˓�����j��'%R���'��=�3
�.C^�B�Q	Z.h���O�>鲺iD��6��	ɡN�mr��ˊ*��СÚ�k�D��!�&M�,�h�N`�pA�O	�J>�(O�L��m�J�����	i@50�A�<���?���|j(O��m��6v6@���v��&���)�N�
@�)M��� �M���F�>�6�i"��e�ƀK���'�4�0��p\P���
�Ga�7�&?aE��=��)'�䧰����N�*i�s��:O��K�#��<����?)��?A���󉚢-��Q��"[�����Caڠ�D�O��YȦ5�!o{>��Ƀ�MN>�&N�:U
��s�B�h>�!��ڵlb�'�x6m��)�<eL7�!?�&_�U6����;󔴣Zat�0Ζ (���O�	@y��'LB�'�ꏶ
m��sG��l�.�{�M>�R�'b�	-�M��A����O˧#��%�5���7
�,AE��8�O%mڷ�?O<�OD�Qh�$G�.8|�D*~�1j��Fi�����i>��6�'_|%�L��O�xĞ����C�M���p��ҟL�	ȟ��I��b>��'o�6-V�6z���k��g6 �q�<C������O����̦��?Y�S��Xߴ�ؐeM(�.U2��S<=Ƭ���'S��J�{4�6��ؙ2.TG��$)Ly�B ?Q�0)%N>BަA�f��y"U�|�	ӟ���ܟ�����ȕO���!�M�(����x�D��w���˷��O���OT�����PԦ睊k�(�[��K�{�0Y2���GU�(��4K��֩>��i+3�27-�|�u�-r(�����U�%�P�K1ni��"7+�	KB�{�	Iy�O�"�;T�6�X��`f|e����/��'�b�'��ɹ�M��E��?���?�GJ^�q^ ��ԫ,�d��A����'W��a�fgjӢ&�C��Q�df�*�(*�e�A�6?9U
(n*dk���G�'c)j����?�r�T���!�l��h����3�Q;�?1���?a���?!����Onu�V��-I��R+ �vIΙI@��O��o��h	�'�*7;�iޡ���V$��Pp��?>��Cp� b�4}��o�Ȫ�g�Z�"}}h��柪RV��k��q�`��ш��`��h9��<ͧ�?!���?)��?i���5H�T[�.��f�4�������ha��ߟD�	؟�'?�� v�R���
,\bIM�5�ΰ!�O`�lڅ�M���x��T��� 
���R�vV�	��1�@�f��u!�I?�b��d�'�BP&���'���Fl��.]p��τ7� tQ�'�2�'�����4^��۴K�-��m�D	�OJ%�Ԣ���!k��̓����DJ|}Bs�Ʃmڴ�M3������j2Î4��¡e��J<�t�ߴ����x>������OB��]�2��JI�70Z ���$�y�'�r�'C��'+b����
�p��'K�'eF�"B n�@�d�O����ۦ�P�Iyb�p�>�O�Pc�Ɨ�D��Bd[9`,Y���u�ɞ�M����2�K�-�Ms�O�P㲦G1n�L`� 9#6�*�^"iNS��RQ��OF��?���?y��Z]$�4�P�"�l�Hg�S%0bh���?�*O`�mZ%�'��P>y�m�yb6�C&"xBx�3?�G\��c�4��xʟ�5�� O�֌��L/����� $�x�M֨b`P��|j�"�O��	K>)ԋ��H��D24���9��C7�?A���?���?�|:(Or�oy�y���8p'� �H�vK�QS'	�柀�	9�Mˍ���>��i��lWF�����@!�4Bv`lӠ�o��]��Lo��<��1����� �X*Oh�1�HX�gŒ����*��<O�˓�?9��?i���?�����1b�9�E��� �5�S/1�@n�=K'j��	⟨��g�s�8c�����$�?u���MB; �t��s��L��!�O�O�����A�>�P7Ma����g�$F���m���gp�8J2nD�Lf��r�ILy��'�"�Ε��5�e� �9�t9�߮I�r�'R�'U�ɾ�M�񡌜�?���?��_&���;f,��S���'E,�v��v��O"O~�(�V�x�D-�� ՈR̂ةE<O��$� dtx2���Pn�˓�j�!�Oj���fH��P�ݶ"�v�����T~Q���?����?����'�?����?�)�(�����b�8!��D�vmQ�?!��iږ��'���'l�]�l�i�咅�Y4z@T,�!�X�=��$���I��M[g�i򩎹d�F��؃��%���$z��#U�G�6�Zae��\�ZD&�h����'���'�Z֛&�D="I��q���+"%Ѣ}S���Mv��?���?	I~Γe���
А5�T� %A@t��#E^�L�Iğ�%���"�zR��z2�H
l��C��A5	S �;Ю> �ʓ�4Mِ�O�d+J>�(Ox�0��	+J�Y2�D�:?�<qr��Op���O ���O�I�<��i�^�1��'Z�$h�ib)c��Ǻ�#�
�=���Ʀ��?�4Q��i�4:�B�i�T�ʇ�@�8��8�l�-.z�i��6s�������������/g�S��Փdlׅ*G����$C�0���P�x�X������	ߟ�	՟��F��<D�X,��^�':-3éΑ�?Q���?�3�i��1r]�dKݴ��I�8�+H��4�[�(X�%)����x�"q�V���D��czӄ�K�(���,��9s��`��}������4�|�D
������Or�d�OR��	�\hP*�^�j`(8��ƭt����O����E�.s��';�S>uS����/:�j-"�Ȇ�:s�I%��������S��lA�z��a��?	��9D�A�0�V �
R?2����u^���J���k�	�,{&RD
R�pbe�t(�+)���I��I۟`�)��Wy¤c� �32	��bG���������$;�����O�!oZ]�W��	��M�K�q6!R�V�gϦ�ڶl��2�i��h`ֲi�I�9����O�xM�'Z���h� /ТeI�dZ���Z�'��	ӟ���ڟ\�I��H��s�����ݞ)�F�+���U�^�avNq�H�R"5O��$�O��������<�jI3�P*�� ����-|](A��4ye�&*&����<o��6�g�X2sg����bfhK�Q8�zF%q��� ��f�r��j�I`y�O���&(=b�/�ɚ!C0C*J�b�'�r�'w�
�M�W���<����?�K�<�Y�C��'��Kd�����'��L��dӊ�'�$��G�|�[u�B'\r��`${�H���U,ĲD�X�	I����t��O��A�s��E&4f���8���^<H���?���?���h����%wfha�j�+n�!!`B[������Ǧ#��`�ɯ�M{��w����U��
DZ싓*��P�Db�'5l7��˦Y�ڴ�:-�۴�yB�'���x���?��e��5�\H��Y�2W�`�w#�9r��'S�i>=��˟��Iʟ4�	;I��� ��|��/��!�ݗ'
�6�90�l�d�O���'�I�O�ܣw�(E�����ފO�4��vE�}2�m�j��Ik�i>��S�?Q# E��Aqa��^�tX�@W"m���h�iFy!J<]��}���Q�'��g���ihګ>�vU��ڀ0��	П��	ߟx�i>y�'@f7MF�?ST��]��\����M�e:i��LYD��Dʦ��?)R����4u�ijX��׃H�<6�2�nƔq�.(�"��8]ڛ6��8���
U��T&�_����SEM�
���k�f���W�c���I����I矘�	ß��r/��qs������L�P�Ӏ�V�?!��?��i� ���O���h�J�Ov���o��* ���n�q�e�X�ɋ�M�w��jVN���M��Oz�1���"v$��bF�5��D�,M�~�(���"f��O ��?Y��?��1g��)���R�H��55B(����?�-O�lڭ?a����@��X����k�2l;��M�\I�k��U���d�Y}�Ju�8���F�)� *�Ӆ��b����9j�H|;h=%h,ى6[�w�|��|b��O��O>���Nv��3c�ԣ-�%�'CP��?	��?��?�|�+O��m�(4��o̶|S@�I�(Z�r!I�h�џh�Ƀ�MC�&�>AѴi�0���üvŰU{��V�[=� �d��O86-	���6�#?9�a@�mކ�)׭��d��w�>�Ard
r���q�Q�J��<9���?����?a��?.�
�s��0J�:s��$��Zs(Gߦ�z�A�矰���� $?�����M�;iD
e��T�+d�P�7�H�n���c�i"�7�Y�)� "L��l�<�� ��p���f�g�����N�<A�iD�FkH�Dʫ����4�@����9�����_;���H���H���O����O�˓52��Cߠ���'/֋R�b!
�-�v���K㬊��OBu�'[d7��ڟ|%�pj�D�>��a䛌/�Q�1?���ַR\��a����']Z��$���?�QiH!+�)B���Ӟ�S����?i���?q���?��9���8#C$
�����\)_����M�O�Po�����I��Tr�4���yW/I%�G�#��a�P넩�y�&x�ȥm��Xʓ�Ʀ��'��9�p��?1Q�&�X+�H�7#@�x�)�
Q�Ii�'��i>u��ɟd�	�x��u`l�%"S'�zj� �C3�9�'Y6��6���D�O���.�i�ODk#�����T��on�aKvmLv}"*o�l�n��Ɏ���53+�!�D�b8@q��ayH� ��̡8�ɶ���a�'<p�$��'�^��!���Y�v�7R�"�'y2�'����S��Cٴ`)���sW�-��*
�o@X�yQL?�P�2�u��6���jyB�'˛��'b��ach�!aM´�T�?���:�"I 8i����l�� �h~���9�@\k�����T���9o���T2O���O��$�O����Ox�?�1�T>y��*�������� ޟ���ß��۴v̧�?���i��'����A��<#%$��Ѵ������'���+�Mc������՛ƙ�Lr�\{��Rg�!n��%���2c��y���'l&�|�����'���'^�!RuJ:Y�H tR1�䉺��'��^�@�ݴ=�֭
��?9���$5�Cp�tf��eٖv�ɣ��dM֦уܴ�?qt�铝7J�`��F�gy\�AP�E9n`4�ɳ1&!�!�6��擦cJ�l�k��(�e�0^��R��cY�H��ߟ�����)�cy��m��PK��D�^W�<��+�/	�2-�C�-e�L�D�O<�nd��8��I��M�t�ʟ5�̹`/Ч*��QAA�	:�F�'�Xɡt�i~�Ir�^8�w�O��,��s��]�R��`4i�B�!̓���Oz���O����OX��|�qMͅ>�:�7��jP�������V��x��'����'��6=�
���CӦ+�p���	k���g��ʦ��ܴ�?�)O1��a[��v���$g�����r� O�6B�?N�9���'�$l'�<�����',R	3�F�Fܫ2��@SS)ޟ���֟��	ay��m�6�D��O
��O�D2r�#G\�8�3�����ۗ�+�	����O7M�O:ʓs(���A,M36z󌐩t�
5�'�f4�OMjq:���-�̟:e�'���@��J?@���vN��:.>	��'K��'���'��>��	q�>D���,���Y�Ϙ_cq�	��MÑ#�1�?�����4��)�w*Z�V�>9zao~<[C�O���q�h�ҕg�86�!?������ܩ�p`�)]�9��}Cwj֜'�ҡ I>I/O�	�OJ���O2���O��sY�l���Cϼ%Zl��FA�<�պi:&��B�';��'�����	�,�`�# �UJ.� $�Aky�'ᛆ�'�)��_�t911f�OI�Z�����HVb\:>L�q�'$fQZ��D����|�^�T���M�x�$PY�.�+d�R�)ϛҟH�	ß��Iȟ��Syq�����O���HP�=��a��8R1˔,�O�unZ}�I��ɣ�MKҼi�b�ѦB��M��JoF&a���#bՆ���i��	d��Q`��O
q��N��@T��37���=t���b��e���OZ���O��d�O���*�ӤO�<!��8	�Բ�ᗼ$E���P�	 �M1��|R��x���|B�4@m��3%":�z�p��$�V���ٴ3f��O�d�i��I 3���c�D�2gF�s/9bd�R��?p�g�~�Iuy�O�"�'��P
o���6�^�)؀�������'��ɜ�M�ANɷ�?����?a*�X�i%N�u粸�aUq�HM ����0�O�El�M+��江(Hk�dP�p�n�f�� 3�&�6/��ML2�p�	�f��i>��Af[=��I�7!8A���.D�a1~�ؖ@֦^����E��d�5��`�w=݊�Z
ui���.��TX�-����o�8�%�R7B�G�� �E� �UBmБ��O�8`DHI!_��$rs�Z�FHVQ��E*e2e�nO�� S撶b �A��U;Ԯ��C]:q��R>M�2�kD4E,%A����&
���ڥX�< P�N�'�0���&��jdM?^�c��B	ܯL��D�Ђ��X��3&�?)�8	;W�E�-�&�#Ff��s�*,�d	�y���"�>�-O�$.���O�d�#M�8�"�۹{'Ĭc���k����#���O��d�O��+�b���7������̡V����6 G�7�<#��i��	֟�$���I֟ 2�q?-،Rh\*�� �a�O�>��'��'��Q�,F�����I�O�[Ս_e�Tj�Ǉ��D��EƌǦ��IX��ٟ��ɉ����=� $}�"�m�]���N<E���iN�'��I5<�
����d�O����(8@�U�E*�W�Z {��]�a(U%���	��@xЇ@v����$���Z+0,K2��(]A6}�fC��M{/O�Eۦ�D�)����(���?��Ok�/��	SJ�p��M�AG���'Q"�Ŵ�O.�>����Rt.��S�n� ʙ8Yh6m��A��m럘�	֟��Ӓ��d�<QU�.L�^���\�u]�3��3�&���L���d3��Οt{d
/G����6��q���M���?���Ie��9�_��'B�O0��iQ9��U�E�Y3�BE�i�����O�P�Q+}�П�������hT��X�r竇�h6�hb�直�M��(�H�"]�\�'�V�X�i���'��$S!����K�:�$��%�>�H�$���?)���?�/O�qʱ�� d�@�>_J�8��CP�Qz�|�'������%������dz�'ì?������u���c��'M��&�T�����oy��'vv&�Ӷ-��z�M
Di�'*Mഐ4�a��˓�?qK>���?�����~�ݵnAШ��jǖw�顳K.��D�O��d�Or�A�h蘥R?����n�Y�4��O?�	��A4�� ;ش�?IJ>I��?�6���?yQ��e}R��{&v�rP�ƱjW@1������M���?1.O``D}��<�s��8�`Č	Kc㗭q^�p��
9��<��A#�?IO~B�O�
����'g��x��
B�DQ�4����Q$n���s��Ia~�(�d��ae��N���C����M++O>�3���O��%>�Oc��Шs�Z,;r��,o���M�G��f*e��7��O���q����}�i>����3B~L��ɺ:���j��Mk���?���S��'R�ЍZR,��ѢӼgɞ�����)�x6�OX�dy� 
&��O�i>i��G?�&&�#rDH�f���h�y�̦���H�I�������Mۢ�Q�4�Ơ��F�o���㇞ɦ!�ɼe��Ŕ'�L�'��'�*x�@�-b)�xƧΖ"�;`�"�d�"R�1O����<9�n�45y���<���SR�E)̀���O��d(�	ԟ��Z3T�"R
���P�Rǔ�[�qlZ�%��b�`��Yy��'vR�KU؟�-s�L޽#n��	�ʊN�&k��iB�' �O��$�<� ͦ�[$閅l��;�c�L2�p2�2�d�O�ʓ�?q&��9��)�O�2�#X���=Z`H����{�k�ݦ�?�����w�'$����$�~t�&��3coI��4�?q(O��D<?
ʧ�?)����}E��)7�@�N��b%�/"���&���]y���O�L O�61�"��8M�L��J�/P���Y�� A �M;Y?Y��?�A�Ot�u�ՕM��ix�E
��``W�i��	�,�ɱ��'��禡���W�j{J�"��	�o¬�Q��oӚIaFM�ɦ������?i)I<ͧF��M���?�L�f�&`���i�i��'��|ʟ��O��Hƒ>#� :��1[��-�w��O����O"牉W���&����p�}�蠃��^�WO"$h�Ⴡ6� 9n�ן�'��r����O���O��q&B<`X��x��������A���T��"�>1.O��d�<9���'̙���\r톏9�4����Ht}ҡ�y��'Er�'r�'�剉9:B�#��!Vx5�1��y�f��������<������Oj�$�Of�Xcn��J�D�Y��6��t�I�W���O��D�O��d�OJ˓9T��)e8�깂COB%���b�T;D‌A�ix�Οl�'yR�';BHD�y��ޅZ64ʆ�nު���'��b�H7m�OB�$�O��d�<�cA7����֘;'C��@2�Z�Kf~�jݮ �d7M�O���?���?ib��<	-O�e�f����-��B&^��y��c�y����O"ʓ@���a�P?i����D�=f�TG:<Z,��"Z&����O��$�OЙr";O���<9�O[<5yP�%P�d��iتT�lZ�4��D�|°�n����I埨��������;gC�)}�r��V�D�i���''P$0�'�\��<i���bA�T��S�/܃]i���ȓ��M#'I��i�v�'�r�'l��O�>�/O����J/|T sf��1	t�#��֦��Ю`�T&�X���&��I���0?������T`8���i�R�'��˝GlR����O��	�	h�������Z�E�'�6m�O�ʓ5OZ��S���'p"�'hLrrN�d��4��,����AD~ӌ���eThh�'��	㟜�'�Zc����|�*Q�ä7%���+�O� (!?O�˓�?9��?�.O<U���Y��!��L��������>�����?���Ә��'&j��@#Zv*�A��<i*O��D�Oh���<��I�@2�ɑ<O�|L���/% `< ���]0�'+R�|��'*bN�/��ɗ'M�p����#C~ 0ke@�>���?�����$��q�$>1Q"��j����6f��$ѓ��Յ�M�����?���0�^h�{��I�f�3L����B#�M3��?q.O"0��D^B������4�"�j�$��W[L��sO<���?!�h��<�K>a�O��䋑�D�Tm}��F;G�)��4��DH764n�����Ot�i�c~I�0U�uX��Jw���S'�M��?1&���<�L>���  ��bc������q-�L����v�i� ݛf,r�.�$�O����|H&�t���������<N�(IvL�1���޴O6$�Γ����O�R��G��� P�[�u_��9 m]�7��6m�O��d�OTt���CX�ן,��C?�Ղ͞?;8�(�a^4L*Be�e+���%�Dۓcr��'�?!���?i��ZQ� �N2m�8��C��'��'|��J&8��O:�d&���ܴ� m �p�f��+��H ��BP�$�1aa�L�'��'""Y�02�cɉ�th:�,!N����Ou�|��}��'��'v��'=h������B�P��RŐ+ ��}��(��y"\����8��py�`
e4�S8=���'�^�8X
�j�f[�_�^듻?������?���N:���EP�,@3 ��I8���֥�7�( 7\�T�I����xy���$~7����F��5Y����ܖR����L�ᦹ�Iv��ꟼ��hˌ�	t���!"f��he�Xz��S+1g�V�'�rP��
�����'�?!�'*f��R��5O���w�ԆLI�L�T�|�I��`�I�g#���f�	GB�	�&�ře"���,�w&HΦ5�'oPY��y����O�r�Ou��2{�u��	�F�` 0G$����lZ��0�	�Z����~�ILܧ8$���c�ݏ)�0��'-Τg�Ԑoڑ[3�9��4�?����?y�'[?�O��0Wo��6�>�x��*��`��O��q5�YG���OzrA8�H�"s��:I���Z4�`7��O,��O�lq�"�l쓊?A�'(���H�{�-��X��쭪�4��t@��S���'���'��l�sIж<�yv$�����
��k�,��� �~��>������c�0I�< ����֜:'NR|}⮝'R��V�������[y҉IAd��H��W��stkT.)<�� �Iן�'���	ן�!��EL���RȊ�{d|��wE� �H�	my��'S2�'���;F|�O������~;}�pz�M�Oj��3ړ�?!�)T��?��aĬ yj��1
"^�� p,��GV��'
�'$�X��a&���'!y�M�rnY-AT�\�oH�I�Z1kӾiўp�ɐK����	韰�PW5�e�J�fջ�Ф^��4oZ� ��lyR��=+c����k�٣sR��@���ƅIc!Z�O��d	)�L��'�T?!����n�0A8�N�t����FhӐ���O�P����O��d�O��������Okl	+/^D�S�L	H��h�`	�(���'}Bm%�O&�>iH���:[0��d�-L7�KB̝"�K B�s��cG� �|N�i-�
��]qǀO�DP�qpKV(hF*i��*�Ua��
pI�I�T%Y� ��T;R�Z\��@�ץ��By��j��H�9I��!$�	dq�I�&^�<���{��_<�H`�%\�~�������X14�P�<@�����$#�@�T�3�� B'Y�j��!)s��DdA��	���e���A��hI�(C��\��A9Cж`����?���?����d�O�擓R���#���W�<2�D��o ��Y�B�5"ā��;U"؅�FG����O������H�@�"�$<ߠ�;�j�y�lKcL� L�����9�衱!����x�U����Գ��\�������y��d�OL�=)��DkB�Z4�S(r��qQ6n�(�yR!�;oܖ�Y�H\�R���q���'꓆�LJ��'!r─h��:��I� qC6b��'zB�'p����'3�1�����ڱY���+$�݄'t�7��3x��G��[t0�i
@�x�C�g$�Q��h@7qN� ��i����.��6�|y���3E��u��CnD�	��'D�{�P?z� p���ߦ?�z�y��'W.�3�:V���8Տ9��ě�'��7��^dJ�i7��f�����ޒ\e�<�B�y��	�0�OH
=)��'2x��AL�,�����;(�rЈ"�'}���$a���C��G�`J3��O��n����D������Qل���c���	�0�`�(�gJ�5 ��Q$Yq�O.f\G��7b�,�%�1!��́J�<A�K�Or��#ڧ�?�q���n*�ې��U��,��%�ȓ�{�ő-��Pr��11��	�HO�ștBʸD����1�ȭ6�,�Ĉ���e�I���	��Z��G�֟��Iɟ����}�a+х+,ze���Qul��W�(���ɑV��ӠM�+�<b>�OJ�RPLk���
qA���4�L�7�����O�HIC�3����N�8��6v��0$�O�QF��yR.O��?�}&������(�FuS&�ާa�8���9D��Cwo(s��d��!�)AX�:D�*?1��)§m�vdAP&\�=��ݣ���'a�V�H���2����?	���yB����d�O�"4�,�"���w�4FОx~���Bb�)"��z�͝�w
�q��	�-P���SHIu����W�s������B4	�J�P���-�i�牵�"Uh��
�cj��Ə���9� �O����O����b*��M���4��d#/T�iu�sФ��]� ��i �"+���D�<)���"?��'g���R=a�@{q��sFɄ�%�r<O����'�"?�܁s"�'{ɧ� �加��E���RE
V�����')�Q:�Bj�_��d��C���4����p<��Iݟt%���M�6@݄�ġ߹ U"�R�G!D����/�=7�DH�B��4^��Dy��#�@iش��-A@��8��MrvLӗR�$�<����QS�f�'-�?U���O� �CٚqY �aH��pV4�B���OT��.��d#�|�'�Ȥ"�T����)�#&)[�M�����+�S��t@�y�EV1X�Y���;�bħOl����'Q1O�\Њ3L�3[Z$3#&�.�13@"O@ӥDa��u��$�!5�$=���'�,#=���W(@�8�AD�(�
S��I\���'�'��RQI�.Z��'T�?O'n���x	P#��*\�i(�G�\�1OP�I��'�t���A�z>�$!R�Ɲ5��x�{���<�f�ųUb8�It�;�&��V͙$�'�.���S�g�u5����΅��J��QE��'V�B�	(�i#d(�4 �<HJs1�����"|jC��L� ��cs�A�� B�ci��;�?A���?��'6�.�O��$c>���˕8L�Lj�JZ���@ �
��pB�	 ~�k5�X�ɻ@O�$i�e;��K5&B\�<�g�6�*���$:*��#�O�H"A�V5�-�B8�}K"O��EK�9b�iS�P,?�$���$�S�S8���i��'�0ˢ�E3�D�V&^�i�氱��'���9lnB�'���TsW�|��Isw�ad��\@�Qf�W��p<�E �D�X%j9B6�P�Q"����G�#j���	�AaN�D(�d¡p����Y2e��Hó*E��!�Ĕ8P�le����F���r
R�:!�$KǦ�f���hM���퓚{12};�g1�əv{�e3۴�?y���	��E�B"V�	�p �L�Nip}���f.��'�@����'O1O�3?A��7�Б wk�$@����E��V�=���?iy�%HNc��S����Yc�b'}�'\#�?�y����	<d���Q傁kcx9Z���y"��,�P�Ν�n����[��0<�F�4N�rAXS��[��5
�� f��P�ش�?i��?�Ѫin����?i���y��7iL�)��9�PaHU�	o��dp�y"��<���gy�B
]7?�L�����<�`���5~I��O�a�@�$
���<� ���>�OR�a��!���'(�K�<�6"O�=h��/B9,�r`F>!�Z����i����*1�4ڣ�BjXK%C�o �Z#�͌<B*�I����	�,�_w
B�'^�)ǐWTE�W$�k���C�_�N��FO����_=yed(ҳA��]�\-2�*�a�!��=y;������z箙&��>G\x���'�"�|��'�B���-y�>4�6��F��AK��P�J!�P�66�]�c�Tb��݁�Ζz�1O4 �'���4,�RqHش�?1�\v�$��F@v ���w��5q��a����yrjA��?A����ԢMD����Z�N�<�uB¼I�/X����h�d��	.�}P��
�H��f�Ɉ���L<Q�J ��E�r�x`K��'�L������a�[]�n0[Ө�� N<(��_-�]�c%�.6��
d)ѩ9+���� қ�]�W��<��@�b�$�jD^���'A=�'.nӎ�D�O�;v�	�9��q@���v���FQ[_��I���џP�<����<i8l$���خ$����Ѭ 5�~&����E�;Pg�d�t�*�F�2iR��ΐb���R�k�+0��Oz٣��'1O��`�	 )R��M1����4���"O��x&�Y/WV$�KV��R��E�P�9��|�!�I�~�@�#u�'HС"V�S<<~L��4�?���?Pm��
zT�J��?A��y�;W��y���0��c�$��j�y�y�����<iG. 09�/@2hs-�/�U��N���	9QPxeS�������3*�!o���<�s*����>�O8,�HJ�c,ؘxRlͭV�hp02"O��e�ݒV"�P����xp�r������ᓘ����'=����ꞼOk TB4���}�	՟P�I�<\w���'���#\��S�J�P�j���H
�mGJh@�O&q� ԍr���C�a0C��-&ܨ��1��R��j����b��q��g����f��5�O$��ա�9Ybq�6 �m�vQ
 "O��7��n����AR�s�(�*�u�O��Xs�i��'�yȦ(� ��L�w 	B\����'��d	x��'���F��!�&��fg�i86|�`q1s:Z����O�a�jS��'��A 臶����"o3���N�Y��i�k�(m�u2f)�p<�c���$��WJ�Q���ѧ�Qa^��ǡ(D���(�!2�ޝ�È-N>����2�P޴)m0lH �r$��8�
��^��<��ţ.���'-2�?��V"�Od�Ӏ/�P�\da���k�H��� �O��ć�'j���4�|�'�~�b�&]r�-(�
W�8�~�K�D"�9�S��=.������?��㶅_]���O����'�1O�xC��$zB*q��n	29_��"O�8���E�1R~�Ň�
O�웶�'�"=1�Ê�0@IWD�Y��tQ)�'p��6�'���'P�a���+9?B�'���y�f��qΉy��L�7�"�s��?^	�'��\z!�$glџ(`Մ��"�)���TsDS�m"[r�^�(D�qAA�B��>1��AV���$�`֘qn!u��E��%�Lfum�
�M�g�8u��8T�������h�&E2,_0��%�N�BJ�{b��OT��ʜuqʍ�vh�1�4���فy��I��M�%�i��+n����|�-���
p�\�
4F1�m
�xs$\3��-Xp�jG��O����O��ۺ���?1�Oqjܠ��	��u2eh�b�J�`��ܿ�BKaEW�a�Ԥ	��IT8�hr��� tR���/	�
�qǭ�l��p#!���=9�̀C��x���
a�Bْ6�BXդs���	�?�5�i�Z7M0�I���OC@��&������� �bLK�'�X�i�.V�P��YpC�(%�B̒�y���>A�yҙ�Į��$���}����o���y��T�t[ȼ�� �4|
�<Q��N$�y����f�N��kZ@R����)�yr����++��?)�a�t)�.�yR̟"��m��Dؐ4n��4Mď�y���<ߢ5�FK74��-`�����y"�"w~f�{������C�O)�y"�,��I�S���^V)��_��yңܿ7>�%h�T5m����W�7�y"(UZ{tX@�ۖk������y�����u�\$d%�4j�)՝�yBNr���3�Y�s ��0����y҆ʹ0A�:eHȶpFf���y��tE��x�A��	�Q����y��+w�`�q��c����� �y��e�y����`�~����:�yr��)�DY3�I�VȔ�Ӡ͛:�y�c�w8��g�L$oͩ���yBo]	��2񨃻s�&�j���y-q���B !6��l�7�ԏ�yB�D�
���5��@�Q.�yb��;Dj$a�cK. �,�ъע�y�eT7LK@0�͘�u`�䀴����yrGτ1и@k�o�.u��������y�٠r���O��g�@�E�L��y�63X�x"0jk�NX�U*�y�A�_j���w��!��ʈ��yB㕋9�6 ��_#j<T��u���yB7l�.���n�>h	,����:�y�
͖}<vu��8����
I�y��� �VT3�]�6��z��ߏJR)R���3�g?��	ή0d��k��0~���# �H�<	��.ԱUaK w���Çϟ��a�@_a}�	������~g�٩�j���=��������_���l��-6Uذ� b�쐅ȓC�脲O�^�#"�D5s��0�?��N�"��#�a�1� �"��x�aّ�Y�<� >��ܪ_�DY���b��1��BXh؍�=����O�Y#�j�64��B�%>:��)�"O�a��/�8i�&'U-��&�'2N�Q��tX��j`�����sm��d��|�B>�O��T^d�Iюļ.M�Aᔊ��""O��ǋ�=S��PP%��K�l	R"O<y����
4%���D��U���J�"Oj��q�J���APE\�Z����A"ON�	�͂�a�<�B�
k�L9�"O���e�#՘��̅2�z��u"O�� �%D�uL�؁��#:�0�8�"O�Z�O<�D���)f�(�"O�4(� ۺ:�V]`�`֦}�y�5"OH|�bb@��h�B��\��)ð"O�5�ro��a8���O�GU|P��"O� �t��L�D��L�/Q�e�"O�x���P��Tk��]f��	i�'TƐ����<-n���[��`"
�'ւU�'fT�9 �����:
���
�'�*��O[����3���L	�'�&iY��������x���'\��JG�@���n�4l2���'>�ld��O8=J#N��c��	�'��7hǊZ�(�i2�;
��4 
�'0X�,\�^6$�s�hP
���k�'?�Ey�@W��ʘr�G��Z��X�
�'s���w�P��æ,�$�*42�'k`�
�4J����ԓ{=`�(�'j�1���-:4>�%�مj2�`�	�'OhXb0�I�pM�K�A��dP0	�'Ȅ4��"ހ�f@4��._����'���zp�;ET!U�C�V�b1�
�'gN�j$��$(��[Ĩ��N���S
�'����1S�<uDm`��HB���'ʺ���îs�t��w�M�58�Y��'[�\�
��V��
��^�v�K�'��Q�*Y�%�В��S8�����'�X�9 �I�K-�M�Q���	�@�X	�'&ܘ��ZO܀�XPb�|��qB�'z��fH�	޶����%w�Z��'c��9�k	>�<h�ፁ�"EDh��'	nx!5`��Z�PA��,�AxA�'� ���K�LY��J�t��'��}�4� ��h�Cw�+hn@��'V�c.�	��`�d&^��]��}�$��আ#���lA��nC�	�wx���2D�g��_�C�/̆؈���9��!�ujO> H�C��-Ė�1c��{�U��&ۢ01�$[��7�����_�ΰ>��ԎN'�u���טS���!��G�Tz�$A�ּ��	���L�C�l�"�e��KFvИ���uN��b���/�)�����I����'WF�) K�6��'�(�'mٮ�pU��>�&��Ȑ��ܩ��!�>a�L۴ݘ\��bQ�L�~�QR��Y��	��D
t#/�3�Ix����9��N4@��ɷDC��x�_1hFP� �;���ʲBJ#s�Xy�aX
�#*=�OL�&ēp�� H��T�I�\)p�')���DA� �JlfJ�>���G�<��ݠCfNj�j!-BA�<I�E�/)��
�g�*y�+D�F~���\�kֈ[1��"�&K-��ɑ+[#05j����E�<鴏�L�9چm͞W"!���J�H��P����	�| �c>c��qC�Zd�a�+R'5��4B�%<��1Åی@����`R�F��3�)~��HT^n0�)�tB*�UC��8�9Iҡ*r�H�ቪZ����H�
�@�#�O� ���Q�@�j�=��c̾�&0 �"O�����
(I��]�Kk`LRq��p�@Kй����$♲�ȟ�	�"G�
�VJZI�" � "O4��&lY��Ы���q����u@R�hʆ��'� �Õ/����Ϙ'O�u���Y� H-9j�KHf8��'G�U�q�ʩW��@"�!��M"��V$���:E���
,���$���eIGj��%G|�˄A�=B:ax�-J8V#�yb+_$R��4 LrU-^�r���G�	�j�ȓ:_*a���;���I���U���J�JΕ�Wp��ӭ:�*$�ȓ>��Eh'�&��`��HU�9�Z��ȓT��8 Q��#!����ũͦ$
�}�'����M�6$S��3�eq�(�5B��a��O�b����"O�0ۣ�
ڰ� �� 7p2i���}Z��	%h_���A���g�A�A�
�9�� �]���ɟ<�X�'��=MqFU[��A�n�0��@�fL����oE�E^��a���p=�֌��w�@l˂)�?���CL��	7�,�fbӚ����-� ��&�ֲA\�Aȑ� )I�I3n�3R�ؖ$� ��|
	�'؄tj��ůMG�I��CJ�z�B�MI妵���	S~iKPGJ�u*��PZ���DZ�~�R�Q�w���X��ɈQ�(��Aʩy�����'��A��$�V�t`ܞl���8�!:Prz`��a�mGF��	�w�!�&�u�g¡1��$8���<)�
(sW̩�G≃*�Y�To�`x����∁.��ɀ"���&�<�$T��F�NN���FZ�Oz�8��DR�
��[f�Ϳ{�$$���c�'���
"�۷HTxf=�\kH>9�À5�|�'_RQ"U�=H˞��t�YoU1�-ь	?e ւZ�Ae����_%�̛�+ �OTXS'�7U�jt`"�
�]×O�7��z�	:�FuT���AM�z�	�źi����w�(�����;ɂ�2�q� ]��'}��cC�FA��3��^���eT2�Āj�#�� ���O��#�C4�d�����ɍ3�L=�1퍃E>6����ݛ~���䌁A6&���O�x%*�7]���SCJ�S�P�xQo���?�։S�X�$�9#�w5�I{!"�W�';ณ' C�]��Yш��P8BN>IQ��{�@�&;r��?֠s�`,2�� �E1�nPK��\��|���JQ>�^���'�򨑕(�!~��q�e;LE�g..?��6xBf�Ȁ�E.Ur�d;�cX�y"l��l��Γ	4H#@l��;}� �p��!�*J��u �"�$���E�۹no����EG5R�Ia�e�>yG�l�*�1�D��r�����͙%hf�H3�ѧ*�Rg�;���]�H|��ص�ݍw�.y����}��6��3X;�����/��GǾx��T*�ͨo&�CM7n���Z�, O��
$d-\���'J{�*��b��XCR��l�R�2
��".�9*r�:�O&��A��ڐ�D�8L)r�	w�>!Q�^0R����ğ\z��L�<%?Y���v�	�e��B�>8�"n#D�����>=t�J�lޅ� lNh���ɳw�xݴp����~b���K���4�r �c�! �"�?$�x���Ŵ3��y��ì_� ��BE�^M9�����y���q�4��㉄<�R�pA��>.���D@(�O�����)�$)ߒT�����mQ�Q�n�����J��:$��ScRL��b��A�0����+�	p��X�N�Q����DS0]���{�۶>��ҥ�'4�H�Ѓ���V!Yw��3$���K2*�
5|���Zi�Pa�.�V"X�9!)T����{^2x�<�S�%��S�� X���\z�<����7�A���$km��;�Őu�&oe���?�}��Ԝ=�������Z�����x�<�̍�p� �SE�a�6IH�h�6�@	�{�^5�s�LX���I������Ɠ"�朙�I�]�=�A	�#MW`�H�oϛ�x�~���H�T�_��`w�'��<	��U�ۘ'q�yZ�(@t{X�2ue�_���#�'Ή�sd�3;��#P�V� M>��#Q�����O��2�Õ�hI���dQ�ɸ�'�HHBK���(O�=H|R�r��K�axr��0w"��)��_�Vg�41��Y��yF�,y~E�F`K�`�>�pVȂ5it���'�2��F�R��D�5LO!b���[��� ~i0�٬3�p1"��5#�\yA"O��R[�3�5���S��Hj"OȰʳ	�=s��sc��{�s�"O�<k�b�����$.$����"O2�0D��0V���%W1m�%B�"O~�2A":8Hђ 5NB�@"O�%+@� � �Hc�"�2���s�"O�)#R�ڇ��A(c��77ED1�"O�� ����&���Z���>5`H� "O��#g�گ4q���<o�h8"Oh�CR �uV�y�ڧ\���A"O��XI ���ՠ�7x�v] �"O� �"3f��8рދ_�؀��"O�}��h�xU�PpQ��%YÖQ�"O��(�D>[¤�a�4�(��#"O�=9���7�,كF�Y��P��"O�5;�g�:DH��en.L�:�"O�;g(ü{|0Y�U��,70�5"O"=���? ��c���_4�К�"Oހ!@L�x�:݃��kA���ȓ%�d��I>8���� >�|��ȓj���p� A�b�\��c�J2����*��"�Ӧtց�j�JkB��0��Pp�_�-���b򇙌h�ZL�ȓ?�Ƽ�F���(��ځ�4M ��ȓ}:�TDIܓYG6�W��c}�̅ȓH��HeM�M�l��ȓ2��ٚC��@�i�4옅+�d��7J�\j����򨪴擺m��C�	!y�bqP ��(I��xa3c�mhtC�'.NHP�E�Η2�V��ga�$�C�;Õu��:c�p�-�4�J���'�\�6f��Z-~�"�*���I�'�<9���"V�X\cGCD'��đ�'Z��`n�b����ʍ�lc��
�'y@Q��ٵ;��Z���i��Ur
�'xZ��6"�?�����%`�����'i$4{��;D�h0
�,K=��Z	�' �� �iI�Wj>lS+ʺH�`y2	�'�80q��L�4�(<	׮ծ���	�'��hsO�[�� �-F�Y�l��'��UUhQ1W1<q���4t��"�'�x����4q$��đ#tB���'��`��C��)�L�g�J�nVu�
�'�j�ғ"C�A�4��C�
b���9
�'��]*�D�(Cfl���F��YB	�'����5#\	�������=��'D�x��^�QD�U��<�
�'�9SV� ��3t.�<t����	�'���#eı>���F��gX&��	�'��p�0%GWCL�!�팉h�,���'�@ē�+:n��%� Ƹ�b�J�'���i�f��<'0,�D	����	�'��X�.�-Y"ܽ�3�!,Y�	�'RDP0%�X ;�6���%8%�6�	�'����P.؎oj�`R�bH�"`K�'�%�ф���\�� �F��t��'�=+P��h$��b�)|E�q�'d<ɥF�f:U�5�ʅ
��!�
�'<������5��6w�K
�'2t�%�5w�2�M�}��y	�'b��v�0I��!��|d�l�	�'6�}z��X1l�.5j �S�f�4��'�(��G?s�$���L8KP5���� ��H�%C0m��UI� U_����"OH�h��ۍ^a ���,�bh�"O��:�gS�{	Ĝ�a�_�+�1"OD)��A�=Mcr�c�i͉"ɴj�"Oj1��nɸ*ݘ ���YZ�8<&"O��=@D9��I�7�H]ٴ"O�a�e, �gv(!���#C��� 0"OF�{�/�>Ø5)�ɞ+����$"OČ�!J]�S���"ń���"O0��F�� �2���s�x�zr"O,đ��.��AAAW;1����7"O����^L�`L�s��(`�"Op�J�k�B	w�x]�a�Q�n'!򤕀<-��жm��5����r���5!��%
Y(y�� H�d�F��.��'w�KBV��p6nɂq⨠
�'2P��pq1S��l�C�'jzG/S�7���c�6g��t��'B������ X��Ǥa6m0�'�R���9d�3�� h�օ��'�^]CB+ٿ=~�s)�,� t��'�졺��?~� |:C'T xRt���'��p�0u�xI)sDƟ^����'��	I2�@e<�d�r��*[�4i��'����'�+*��̊Rf�� I�Z�'9h̡�셒Lg:EӴ��FMs�' cG!/	�H8���<#V����'7`��M�T)�8��O�6-�Q��'�ڼhT���0�P�DȞ;֍ӷ"O<�t��0#�&Ŋ��M;�4�p"O��֎�,]�uS�J�A��"O挹���l�΀��nVd@z��"Ol����y:�MB��FL�"O��`� ��~x�Yp*�^���"O"�;�ٴ*pڙ�w��{°!)�"O��2c'S4L�� rU�"`��ѧ"O�����<�� �޾\�61��"O�	���Q�������8>��9"O���j�VlH`V�O;*L@誇"O�`�!C)r�S�J�(��IT"O��!�_`� ɗ��J�Z�"O�$c M��l06k(��y��"O�)��%�<&����c-�:��5"O�C��
C��dL@Q�`��"O��&�X?��#ҥZ�v!(�"Ov�U-Ԅ,�x!J���>(j$|��"OzY�"BH�A����-aT �t"O8�&�P�8����ˏ:Q�=�"O�� "	Ӧ!���q��R=I��"O���qN�����L*=
��"OtH�'�,#��9�')p�8T"O�I�FL�L|�[wH	}�����"O&�:Cۥs�+���i��@��"OX��ՌJ�N�v����ё�2� v"O���$�=���{!�˪^�P��%"O�����N�/g��bTDڂl��m1`"Ovi��(�2f���[`Iʯ�ha��"O�P��L��N����ޕM>�P��"Of����tB6%�q�LT@� �"OQ���/ x�����:=����"O4�E
U%5V�e��`�;�$��"O�u�g��L9$��pnފ ��$��"O���6Mכ@��r2Hvs<UB�"On���§q�ĭxlד%X�ʢ"O� $�3�i�>7G���E_�\M�T;"O��0���"`1��d��2~�j�"O2����"`�t�h D�y(�La�"O�9�>g29P�a���A:Q"O(@�Q�X>s>������*6���	�"Op�����)�$��ە=�Ȁ�"O�26'] ]�zT�#\{J���"OB�H����a�#E(4Fѥ"Ov��c- 0l��1$�.��2�"O dh�o��?�聶��A�`�×"O*İ��"/*ё�Y�E��X��H-�S��y�O������W7f�d�'9�yjĈ'ټm�f^-4Z\l�4/�y�#NT��y8`�L+;�t:����yR��;|M��ӡ��Cg���\�y�]�I0%I�`b�X��J��y�`Hm��Y+U�
2���u�F�yb�>b.��p�@|r��`� ���y��N�g��x���v6���k��y�I�a����G�@�Ĥ�Uf���y"�)_@�-PË��m�f��V����M��4丧�Ol����O�q\��r�`?=�*���'��[�i�u�t�K��ݣ�
P���/qs(���O� YD�)N��i� U`|��K�"Od�SQ߭0P�� �.2q\��X</���X8�����)����W���.q���M)lO��JM>IӮ�u>���"@�a�v(9��M�<m���X�"I�*V�6!�f
@ܓ��FxJ~r�b�;z3�)��"�{��8{ͅz�<Iu"�++}е�צW8e���rǏv�<��KI�:�N�¡˃5�F��y�<��I�Kyty*Q�,eL���s�<Q��O�Fk�̣3��P�2͹2�T�<�f.ߔ{{�ݲ�2=���a*�S�<1��1�DC��
^}P���j��hO�O����dI.7�@���JŒ�t"
�'^��Qg 
��֜`�6wd�k�')��!

�~����"�ҟ[����'�z�#�R�R�n	XG�ܷr� ��'d���v�Žs�Y��B���9 �'�|�����f� Y�!��!��'���`c ^fk�h�X,��'��ܫ�E+M��QbL8jI��K�'�v$a��(�M��-��]�f�ѯ($��Se[4\�*�P<-���uc-D��0���C����t��\D1"��&D�L��h�$���6�]M�� 11�*D���b+C	
�,�Ӯ�Q��؀J.D���D�1�~�+1i J$1	@�/D�A�����P�cU *D��G�i�`�@�*�!�:�K��(��<�C͖;y�B���ǌ*���CagNF�<qE%
I"P$���	��[�DK|�<!!�
}0H��Cӂ(EP�{�MHt�<�B�
S�rr d�&N��!��j�<��� �6��rE�98n �
�c�<���8F:�0b�������h��@c�<qc�N�7)"�B#�F�}.�����`�<!�+ݳl`�*��՗|W��8u�P_�<�)�%/��8�k�8_���2�b�^�<�a�  \�"��H4`)��:%)I\�<�D�C�a���f�vB0:�!I`�<)�EP�o�h�
7o���j���u�<�7�\C�����Q�sb��n�<� &1xQH��_��ᗍʯ��Ļ�"O�iC�A4	�������m��@�"O�][Gaڤ((X�J:-�<�3"OL �Re�j1��B@�Q8^�̨
�"O�Q�����Py��
"�\�˦"O���$�-aP�S#L'�p�4"O�dR���Eb�$�ʏN�Lpp�"O��1ド���	��D6ZȁU"O(ura���hS�����n-T�y5"O<�5���4x�L�p���O)d��"Or����F�<F�+&�O���"O\�wI�&�(��Ѣӯ8�Hi""O�
�ܹVE���c����#"O��t`�@�$L�#�Er<���&"O2�(d�$c}�C�F'p,��c"O�1��'M)	{84c3k��l�@�"O�uH�o�,_*m�/�xvh��"OV����\~< p-L6rf�M(�"O���1�3�tA�ʍ��l[�"O 	�֍á޲	S ɛ�w��<�&"O�,RclP�M����N L����"O�����zG�5y��G����Q�"Ol�Y����|�&�zU�F7 �r"O��ٓ�:'�y@N�frY{�"O��I���r"��`����K	��k3"O�TS���G��)��Ú���""O(Tb��|���j
�x�`"O���\C���`��m��h�p"O)ǃ��F��1���m�"OP�z��ŕQ8 j��@�[ȥ�"O�Ȧ�������#ÌB�xɶ"O�0����=|ހ�r�`�z&�a�"O�-i�˛�Ľ�D��(��r�"O��؂�P���h�E��
��؂"O�᪥č�wS�=0���:)�
TXa"Oޡ�W�W�q
F�R$�)�(�h%"OA�3O��KN�����`C�xsG"O�e��/N�@��@���f.�;S"O�q���2j�t]j�	 �=�"OPM£�Q�\��3�&�<��d"OR	K��,��Xa��?(W$Ii!"O&u�!f�<Z���nI�l\B� �"O�$Ca%�u7� �G.��]�4��w"O���K	(t��ҍ�h�D&"O[���$����mB��ey�"Or�`���?8 �س-ǭR��X��"O��1�菮9���уm/U|��s�"Oސ	��[2��ό#Վ��U"Of4�T�3�U�̋8$�yC"O��b�)B�Q4�~�`"O
��0(+MBe�1O�'��x��"O,]{�cC�O�0�SD�"o��XW"O���!H�- C����̀�94"O���,���+�f��(Z�"OF�Q��Ȝw�(A��iZ;�Z�"O���&�<j�lbj�����"O�h����gq�Iu�	.i�	u*O��*���%�D��AΦAR��'�H`�GꚺM�@��nX�7u� h�'�"�PPFF!mH�t�3]�Y2�'�iPcQ$R�bM�
 T��i��'$�(�'��e�$q#�b4$�9�'�,-����<�$�3��N�L
4�b�'�FP�7�Ō'����ま<��ܚ��� ��ͯ~��(s��*n����"O��kFb- ��B BT�YR+�"O"���6�xq�`N	MR ��6"O$A	��2�"��2.��Oj0�Rp"O4��3J?7�2!�d�J�A\�$Rd"O"�Vg����|�`�$X�\�"O�4�6�̬&t��y���n೤"OjȠ�g��<&8�g�D�h�ठE"O�p� �݂I�Ƹ�FF�����"O4@ ,Ķ~N�P��"�+�^��G"O��@�kQ!Gf��a˜TZfq��"O�}��N< �X[4뛟I,R�"O6�yD.�=�}���I񀔩��9D��aGC�kxb�K�m�`L�v�4D� 藃Қ�А�f@�w$D1�g4D��"��|�Q%fI�򀝈�!���kG� �'��&�p񕠇��!򤁝%��m�s*��R��9A�n�!��_-Z8���� O�N�9v���.�!�DP�"mF �D���/��df�ٙ!��4V�#��ԠSE�t{7 C�T!�I���A�c��7)�A�'
�"O=!�D'GKz�J� ܉.Z�p&�2.]!�$W�O���Y��
D��W��<O!�D���)@�ƫ X�ȷj�"_!�d�:$kf�
'I�W�J�+��%\!��
9G��#�BM��rE1�h��Q!�8c)����n���U��"k!�F�v�L!���*$RȺ�&<f�!��,�*WM�#]	|�`d��']�!�$��Y,z���.ׂ !�]�%��!���?��0DA�f�ڵ�V�%z\!���3��Y�eo](�T��텥Q!�D��#���G(=�6h�dK ]!�ե��`#�/G�8�~HP���"&`!�$Ksj���#��@M��/��ea!�DY�$��+�A��N���B���d^!�D��[3N�*��5b��L�T-�2*�!�$.����%f�!�U0O�!����C��s��Q4OeܕP���Sj!��D9�4��S*P�xu������`O!���.oYP��B��q���sa�mD!�$\��BaD��	Vu^��w��/!�!���#��e��wfn��J��t"!�dڨ�h�s�^� ��8�A��4w!�DCs��F���S͂Tz�M'�!�d�'z/f����Q�
	;E�$Z�!�$P'I��ZU��LpG<G�!�dI$
i� H��
��$�A3@�>!���Ac���g�.��W�	c�!�Ke���BF�H9W��1z����Xl!��W���,��;!������v{!�䈪d3` ��m�jn|XdM"}A!�D�+^^$<3�@�"m]�Y��N�~�!��DG?Y���]�#$�m�FdY$k!��Ҋ��PB��_<7�8���'1�!�$�V�X�ҭ��u�y�@���Kv!�d����e��?" �0q���E!���e%�-1u�|�������%D�!�$IP�M0��(�n��#��wx!�D�'h�2�`���LѼ-R���nk!�d���űg��_�dm&fۀbP!��T�&a�vi�i��	���*o!���H�� �C����ud�*j!�� *����S vB�9K'�[�)�H�W"Oh��܆�섢�H�/#����C"O(�p�gҠ_;��G8���:E"O
%�ժ�1K�myae\0dàɉ�"O q2�\>�~T�A�И/�����"ON�pr��:x��p�_�^���"Oa�sNC�)�R�A�@�7+zT�Z�"O�L��I-�Ҝ��̋�;i8!��"Ol�����UQ�0+!�1d�~�r�"Om:B�R�]��{$D<M�Ƶ)�"O��2	�
<�X#'�W9q�U��"OH��j��bx���w)�@8"O��2�&żs�Y9sς&o>}Ha"O���o�v���ط�@5f��)w"O⤯���8M���ؒQc�`h�"O8EeC��e��a��[!YQ�)�"O��چ*%�B�@%�_�6촜'"O��5��$�BܱuJI9N�>ؘ�"O����&�8qj<�/�1 ƺ	0�"O�Hk�`�T����Ө5аh� "OP���oY�*=�$o�)]�u�"O�=���Y,����QF����"O��.�I�1fh���A^y�!�[��` yvhͦ9X$�3Q �@�!���B@�b��><ZL���3�!��
��Xq�6�TN����b/A�%�!��G_ (*� ��-�VIۆk߽Q�!��D}�ȱ���78wQ�Ф^8D�!�$Q�������6�`�b#�!�$� +����(��t ����!��[�iETz�BW�*��q �Z8RU!�$J2NA~�1%���߄�XĭW�ct!�D�)���P#,���0�Nټp!�d��8b�}I`��8��&LPv8!���/��������u&@T��4!��C�,Ѡɏ)�
���O�~!��
�,,������tB׉՛!�D�%�$ố������k�!�D��/�T� 4��s��C(�5D!��1d�8�R-ŭ1�bE�ʵD-!�J<>����$!q�j8C��z+!��BG���S �V0Q2��Ro!�䉝v�Z!{*�jdŪ�@�aV��䎃ft\T:�/�`"��3l՛6�0B�ɚ\�j�*b� >�4�1��X�+IB�	!o*8Q�a�A����`��8"�B�	'8�L�y2D�
{I��(F��N��C�	�	Lt�S-�@�q�LC+}�C�:P���
�M�xw��I��2_�C��0{��C�	�:]�L�񯔢WE�C�I�[��U�sf϶5�ڐ��&z56�O���� $F4=9��?<�B�fצ.�!��"@��L�L,(<"х^�g�!�Ĕ�W�Lq3��A	��
�'�!�䖉Ә��G�T`��d�Jf!�_k`pxS
����
��<M!�DU�^�28�.�!�4�J�I�=!�dE�f�N��s�+���z�"M={�!�՘O���� cOF�c��R��!�$���X�I� )�$�
��!�!�Dvwr,�jR'=��i��Oǀ9�!��V�H� �	M�dݺ!)A��/�!�$Ͷd��	B+�,(�t�[���F�'�a|!["� �9(8d����ą��y
� &Dԇ�&{69B�ZR38�E"OԄ�tN�������cY5K��a��"O��:�ə7_���%B� ��T��"OB�(��ׅB�X5�t�����*�"O�B��	����L���R�"O�C�I��|���ŕ+|��'��'"��>y�'AF��XJꔒ>�Ahg&�S�II���OiL�a(�)ry���q�̊q�<a
�'ɶ죓�J� ���RG	e�Z�C
�'�v�Bcʙ�g��q���.�:
�'�07 �r_�qCE�/O�Z���'�`�4�ϩk�nI��֑J�ʤJ�'�Z}��A�9~&N0��
�Y�6q��'�T�h���l��zsHՓdQ8�H>�������Oߨ�ە�ȀV�
�Ӈ�d��a��'/J��7�'D>^�[��R-]ђ�C�'
B�q�F`+I�f.)e�2!P�'k�����*|�8���g�^
���'�!yƩ���e�P��9�''�X��1(0��G�Y��t8�'>z�%)� 1�l�{�d=R�}�������O���>�IP�|��`���-0�hȱ�K7D�����3��`e͹����7�4D�pI��?7dZU�d#
c����M'D��'c��6�t�k����~�~�Df#D��:�%�~��01�7>�j'N"D�ؚ�R9,�¬����8�`Xs�2D�DB�׿�n�d`Q?.�tLs�1D�t8&�[J�xh�,:-P�ؚ/$D���0e�=Jit����7qW �8d-D����
!Kti/�!X�l��+D��cC���&I�ϊ	>���'+D��c�N�Nt�"��]�
���&D�<ЗU7+�j R�D�$�8��#D�8a��99ئ���]�s
넌�ON�$#�)�'62�����o�f`�wdȫ9�����'n���2�-�D��ǎ��~� ���'Vn� a-�;O���2D�
��#�'����y%R�r�����V�<�fb�G'�L�R�M�|N�P�F��G�<�AdJH�̙+D��VD�XJlI@��\�<I�iȵ�L]��kА+�t2t����x��W�S�O�bV��"A���
�i1 �����"O��	���0�d|�E� �j�Q�"O`���`�o���r��ݢ,H��8�"O�劰c�vP�i�Vn��S.P�u"O��S0M��Z����,*D�"O8}q��V$�4O��^	��'�"�����#\hJ��\)r��y�I�O<�D�OR�d�<+O�c��`Ԇǉn�h���_8@ �Y��#D�<�E*G�<�NLP�Q�
Rsc"D� ��L�,�9%h��ʼ��!"D� [�C��uQ~@	�
։.��l2�!D�xʄO�1Y�T��R^Nuz�M,D�|13�Z+u	���i��xDb��(|O���yrO
�YLν�A&i��H�C�W9���hOq����J^ �q����8>�|P"O�q0ƄԬ���d��ĩ�S"OY�&l$:����+����"O�xDD�v�6 ¤�P(��I��"O��)􄑶�����ډ|L�q��"O.IY���,E��6f�'�"0�"(��0|�Ao�8w;��bC㖁[�ɳ�*�q�<��O0&�04����'�o�<� �Q@�۠W�t��ӑ{��%@ "O�ĳ�$�`�|�w�5zj�id"O!ؑ���"�.hJH�v��tA�"O�h�gI��
V1�*�=і%�c"O$�Ʉʜ�u�\�*��m������/�S��_]sʨҠl���r-�B��%!�$�;H&���F!%�8�Q�
�u9!�D�u�R���E	z������L5d�!���! R�Qag��]�L�)]U�!���?,��J�N�-\����F�!�d¦g�T@1�"��:	�mE8$�!�C�.��ᣄ�=^5�6l҃�ў���y��Pyb�ښo�]� lS'�d�O��O8�}��+�J� 5/�)f�h�"g^&�昄�#�L-�d�Or���@�	ͼ�F���U�����ꕊ���/X�n���b�G�<!��P�O��fک	a����C�<�SA��4- �����p!��@E�E�<!��^�Q��SW��@Ul�A�<I��B<h���J���	ȁ�T����'gɧ�i/�	�O�N���)\�B��L+4G[WC�ɪi¨�Bj/t��J�MZ47��B�	?V��c,[����S5a�1KvB�I�;{=� �
S����A��:B�	qPN�G�hHl�e�[kPC�I�� �AG��Nbdz1a�Z6"��$q�$�q�	?j�D�V)(�j9�d�/��4�O���À�?���
��8�AV��G{��)��=֠�R(�?!:L @͞�}��O.��"r���:�`�:H��)a�!�d�M@|�N�+�8r�:R�!�D��H��M��@K�+n�ȊtÔ1�!򤑢D1�l��߂$Z���D�חơ��%���Ac��1~`��n�u�����*�H��%�ިi�x�Č�x�C䉱W�T��s��8~�jV�5y�C䉀;��� ��!Nf���Ob�*C䉡W��%���H�h7ܣ�Eݡ��B�	������_��L]�]�C��h�	�[(6�ty��V%m��C�I8S�ʉ�	G�5�����%^�qhJ��ȓ
K1��L&V�*�"��#\�h��X���xc˨Hd\��WQ��eRdp!L��	�wKHm�U��Z�j8a�PJ� ԡ���~L�-�ȓqj:���N�52�	��ۊ#ǘ��{�yb�� �xX�b� I��o����<�Fꇾm���% �.y���	Q"D�|���V�o��x���].���1b!D��I��JO���!N� �&�f>D��*��	�\���G�g�JQC#)D�P�b�ē�0Lq�"�!�Z|�eL&D��o^�n������� ���/�I�<��aϙj�nH��ƷP�ΤzԪ�D�'Ra��"�RF�$1tL^o�J[�����O�#~BC���@VlĻ炆�'�T����{�<��L�3ytr2VO@!��e�b�<qw��`pԈ���	�ø�Sp��g�<iVo�#\�&��v"L���a�<A%�=OL��@��ŗ2��0�t�^�<���7�&� `MDHY�e��Y�<р��  ܡ��K���V��V�	ٟ���C>A���)]�2b�W`�ajq�3D������0
�p�mI&g�j�Y�L'D�� ���#F� ���S��ؚ�B=R�"O�T��	֒@x9S�g9%�Ty��"Ov�*q�
22|�8�`L4nl�=�"O8�4 M9J䔥j�]�x�8%)"O�i@G]�{�:u�[�O����"Oƴ 䀏��D�H -0i30"OU^'Q
���ǧ�+�n���"OPt��	@49�:U�L� &����"OV�y�cQ>jl�hRR�@ ����"O�9I�E�#�8-����k� �+�"Ol�˙ f{�Q�gL�h���!"O�9����K�<� -A�����"O���ք�,_@08��B��<�1"O�p{��B�]�@���dJ��9G"O��q���#���E��^@ax$"O��Qp��� ��,�u�ɺO>{"O�����]�)���"Fܐy��
�"O2�A�D`�J���"G��X��"O�Ĳ��zĘ}��o��1U(y�"O�=�G�B;ZOR��p��6vG8�82"O�P+5�Q�!OHUJv씓{0 ts�"O�����n�y�R�ǜJ5�G"O�]�ԠM�u#�ċ >R���p"O�MKנ]�/ٚ�hq�@�s=��"O S�@���(	��ܷMʀ!��"O�Lz��&s$�DC1�\�w�&���"O2��P'X#�����<U�6��D"O��[Q��u�f����ͮ<�I��"OD��AO��X�.�1 4p�@à"O`2%�V���DY�9�����"O�{R$ %���C�*.�5C�"O�(Z�gC�Hu֍�ա�:X��`��"O8�Vd�/�����m\i�,�W"OVt1�[T�VQ�*@�k��
R"Oɐ��Tl��JV��`�@�ñ"OZ�b��ٳ�L�yCҷ>t�:�"O�z��̈́S�j@!�>54Q�"O�!H�]0��K��0n��њ5"OܐY�����B�OX�k�ry�"Ovͣ�@ ���œ����"m��a"O��
�����LH��ˣ*W&�(S"O�`��܃L��Ĺ`eǦTV����"O���k�.&����$0����"O���qE��w�x���`�U���;D"O���H��DҠ��ψ�c���a"O\H!�<<p���ytmQP"O~�(r!P��åM�E��u�"ODi�v!�y(r8�u.^��xr4"O~�!D�?|h�v��=0���"O�YÀ$�*p`r���b���:͢�"O A�
�
�f�C���" � �h"Otܺ6��:L�+d"�Q�,�"O�s�^�G��=�V��[��ͱS"Oh��䏁 U��1�`�3�D5r�"Of=ѠU:8,t ��/Z��6�a'"O��1�AQ rP� r%���g?�4�"O>8bql�(j��;��X�p��i��"O� Jd�̼S^�X���{�Ɣ�"OL$"�C)%)J�B�l�b����"O�U�V*	�*=R�ڴFS����w�OS| T�
87�P�C ? 6٣���y��.-��� �!lv�81HN�y���:�Z���P�I����)���)�OX!Ȇb��
�%[E患1]H`�"O� �`��$��eJ���GI���yv"O^�i֋	H�`�s�(�`a�"O�ufGUxl�tS;d)"�Qd"O�Dc�� �c�D����s�@��"O���� �?�b@@Gű�JdR�T�����l;�҃2�x�
�f��D�O�˓�0=Q�پ/ �L�΁$R������}�<�S�.}�<8ptΝk�Q!F�|�<��#�8A��a�� 6-���Aiz�<�`$ڎ)�P�p`�%����O�u�<�#���Y\�X��`Z$��aQ���wh<�UO�u(��@BޓQ��-Ё,��?9.O��d_�lì��u��%J ��'I�K��'a|B	�,�f���*���r�'�-�y$_�T�A��Ą ;����¡�yrP.1`��h�*ht8� ��yB�T�?x)x�P?�Da@��y"3sJ�@�ꘜ~`��X�$,�y���-�D�QiR9+	�$�U�� ��$"�Ox@�sb��
�b���5����U"Oȧa޴Y�h8$ �m�����"O�ͫ��� �p�+��ʂ�2 "�"O�\K��E.[� pV��/]���Y"O�*�1�| ����w�;Q"O��Zr�\58��D���["O�Tr k�0���d#�P*���D��r��W�D ��dY^Ȩ6lW�<@��	���y"�?/���G�5"�0�v��3�y�'�pN	鐌C�&i�ƌR��yr���h���}9�3��y��JpI��Bi������y��N�˂m�Cڀ��q�1�yr��W�L,s�F*!x��pjS���'@ў���<U-҆F�ЫVa΄���*ZI�<Qu�ہ��N%m�r�{�f�n�<q���i�f�ŖXJ�-��g�<��×�@N�ۢ���9����a�<�`g�Dv�}�ݐw�I�ƌr��G���O��:1)ǉGK��CѢ]O�(��'i�,
�[��	���0�DBJ>���?����O�+'Jl�*DM� �l	�y�,	��Ӑh�7{P�aW�D��y�ɜ��Ʃ��k5B��q��*�yB�i�bY�uk� q��Z%��y�� �P���ŏe���0
�y��H���	��Z �tH@���y��"'	(A�!ْT� X!�D���d�Ox�=�|��X�aA���
\�S/歙 ��y��[$���J�XO�B�7�6�y"���id���I\�5�G�ѽ�y¥Bd4��pK�E��Ɂǉ���y� �6+�f%�s`��<�*����y⤔�q�@�:7N�5D����]��䓖?���d/d���!'���P �&
��yBJH0�f��f��CWi��!�y�W*M9�a��dƼ9O�}��ȝ��y��[���#J�+�@�`�(�y���S!����R�/�>��n��yb�؎t2�q�M�.��Xib+���?��'j�x9c��n\<t�R�V�P��	�',ք��h��Hn�{"��T	t-�'$��+��O
q�NLQb��/L>J�k�'��t��cY7|���P2�H�R��I�'_t�������za�۶I`l�
��� |hpu�MQ���+
[�B���O��A��
�v���mu�J�)D�l������}xg�S����)*(D�h�����r�^`h�H�=�Sc2�����H�-J8���`��m� �D"OF4B"έiӨ�Jr �2V���"Odc�4
����c�ɑe;l��S"O�t���[�=
��x/�'$��ag"O��I���)������l��r�'�!�D�D����$˸j�(����l�!��8d<�  ��E	�-ۆ�Ώ+>�W�l�<A��@�O6e�UbSj � Z�aSo�z	�'���SQ 
�c�|�!�ށ;��Q;	�'cBEJ�	��|8q��£1#���'r6�1�]% ���	�Ro@� �'\�����yY�i�AĜ�^IT�.O���ě���U)��D.�9RU�J�7*!�d���0t�b��6U��� ���Q���|2�'���'����+ϾjO����I
gT�x��V�s�!�DY�-x\�h�{M�IiE�K?D�!�ă]L���G���fV��
+K�!�ňx�D��@�/DV��p�ʆ�!�N�
X���mF�O�4�x�4>p!�Y�?T6���iC'{Ji#tEF!;[!�$��O9�����7M�������!�dH�u��tphыn��ʵ[��'�ў��<Y�ęݚ\+PLːq8�HтD�R�<Ń�-:�!Kg'D#�i�!b�e�<)���ez���Ӭ��' b!��'�K�<���r�)5犊;�,��DB�F�<yr���U��4JE)�^��E	Wx�<i�=a�y��a��V��c��L�<�u 
V����7)�/� Ȑ�!d��hO�'Q�pB�PixR��jɅ�%��ܚ6�(�h�)��I�̇ȓZ-�ip�7p��E�>/C*(�ȓ���.L�o�����H�d��ȓeR�1�͉/N)IWf�7��9��h<w�Dl�FT�F���H�$��X�<��NĲ)���u��l�WeT��hO�}���i�Ò(7>
�����(�Մ����4K�*O�]:!E���Q��N��i!3�V��8�{fjͿz���bs��$ݚi�f�W���_��Ą�$l��cb��fՠ�HFMV�@0����M���١��&b���� �Z�-Ɩ �ȓ�)�H�-q<q���ɔ��?Y��0|Z⛫K�C�`@66Խ�hVJ�<��	AR�ƴb�L�)0�.�j\�H�ȓ�&maሓz���g��̇ȓ`�`�B��z����$^ �ć�D	:\ui�O�$��I" ֬��l�p��&H 7�"$��d]�z^��ȓ[�&���9mT�Q�j�0 *e���D�r�W�-�J];��24=�h���JH#���.XG:-+���Ht<�ȓg��ly�F7(���!�ARօ��=v��ב"P�$ �/Ԡ]�F̈́�RF��@������ �Y3NEv�d9��3�U)d�H�KԩJ')�����*+D� ��$����I��SԠ��0�'D�Pj0��_���k&oRz9�؈`	 D�ԃ� �j��ӵ��;��t�C�	 �����*ε��/$z��C�)� l��gՠN�fYH���R�UP^���	v��Vn_!{T��G�]�h�Z�$;D������)�B��`��Ӥf<D�(�`H�	$4�1d!� /��,�B�9D�@��MǲVb!�r�O�u�<ZP#$D���DÃ&o��,�6�?+��܃5h!D���q��,&���QTa�0/�,i�� D�lh��ˣX�!�ɟ�,����1k�<q��$-4I:��/�!�b��S�	>`�0`��B<�'�� ���	 �6(���{���F�<��̝g,�ъ���x�@�k�.\�<�L�3`�l4�p"�3[n`[�IZW�<�gδ1����B_LR���,H�<��F�k|J��f)L�p��EC�<��;�}�U��L���kv/[gx���'et%��f�$�L��"Fԋpb�)[�'r8`�(՗�x-�2�К��� �'X�)SD�2�Z�*� h,Y�'hD�ń�	p4�(�U���d�'nf�x��<���!w��~ٶ��'Z�p[�h�3N��uZ�͗*y��)�'2�8���0I"��
�/C�Z!�
�'�H����# ��IHj�	*�ܹ	�'s���pcY�gV�8b�It��I�
�'����nY1GT"3	�%�0̙�'<n��B܇ϸђeM?~�q�'��x��"'.�����ԃ;^���'����S��F�� Y� i���
�'�
̸$%�NB��C���d�,�
�'��VB�2x�[�h@�h����	�'�p�tąD_(�)C	�6wX0�'V�d��BN�rM�AbT�G6�;��O�x��&@22�dT�T�:It��"O�Y�Fو�~mK�B�LNP��"O��$Ȱd�V�S��N�8��"O��'ڥP|.�ZGI�|68@�"O<�˦`_8'�!3�'0l.�E��Op�XĝcC� �$/A�j�0�ˀ�<D�H�fn�:O,#1ɀ�c^:�z��<D��7�&�9C&b@�Q�$	�ǌ<D�ܣcˏ%{=<]�!K�%��Ѧ;D�0���2X� �b�<3�AE=D�3(I6^��	���(^��� =D���$!]�k��qC,��k�|L��9D���5�p|�s�öd1F�9�),D�h��͙)g/��Ȧ���Dr�@�58D�T���c9hI�K��1��i���8D�`�w��/Iz`*S�P�&�~��F:D�h;1�@���
v�M%CT��#�<D���c* q|�xRF�E��� F�O���O���<�O�"���Q慵z/���I�'x:��!D�А�	<<p$�O�4��p�!D��B�Hm��% t�#��#�B>D�dl	���q��-_!?Ej\ئ�:D��낭ޞQ�`��D[����B�=D��r.R�8
�xa��.n�H���/D�Xi%)N��!S�P>d_�y���O���O`�O�3�	$r$�sD��
xN9qr�� ��B�?u�f��G&��/�*a!i����B�ɄMے�b%$8��Y�1L�C�	;G���Թ2�|)Q�!ǖC�IJ��X��Ķb�Ј8&� "6�B�	�D�P�:Nf�ɦ��
�$B��8T'�(�ELw7x�: ��8!$ʓ�?�����S�π �2�NA$tP�h>}B�|�)�b�f����J��l)ˆ ��wy0C�.5�T˂�
/4L2Q�T&	"F"�B�	i|���֟j��p W"M�=C�ɰi���di2fH��3Eŏ/8K0C�I�uH��C�E�c��)E+ C�	%3V���k�]u\"�)�, C�I�
Vq{��O�`�B|0d�3���O �=�}�	Fk�e����R�{ch	N�<���ޟ=�@����Z�>��aj^�<��!��Hp W~�v=���X�<�IǠU���V�Բ3X�:���I�<��-f^���3��D������D�<���z���ѵc�O��Q���e�<!�B�{�tY`�@�cB��!6G�c�<��'E#K�z$�vdԭQɶ�*r�^T�<�r��j'`�v�S�@��bAƜX��n���OAd�� o�B��S�n��\b�
�'�����A�2%���P��4i�N�z	�'�Z�Ru�lf!���)A��Y
�'V�Q�&#á/�01@�@��8�Vq��',XL�C����	V�в7� M>����I0wL�� U�N�
�Ą�å]&+�!�Ӄ M�\@ �ʵ]�b���	X�	�!��A��$/) ���[�!�F�:_t1
$�KO�AzGV�!�D�h@�(a%ċF7b���eW|�!�Ɠr��P���܆u�4��ھX�!��x���D��N��D�h ���	P��(����3��%Pta)V���|Vy0B"OTd���p(��jӈÈq���{�"O E�_4.Y*}���S�S֛~�<ٓ�;n��1�Z�+�&�b�<Id�+m�Ti`�+%���%*�T�<q4�W�������5�2}���	V�<f'�Zqx@ PB�SD�d����N�<y�l�.a?h����$���J�<�q-ԣ�<�b�I�tH
my��J�<�ѫS Ijlq���\��pk�F�<a6f�?Kh:��r��>^0Xa ��l�<���_�
�t�P�W&$!!3��<��B Y��<���<5^�\"'@���lG{��ԑ�x��O�KlB�ku!ۿ|�LE�3�8D���Fc�V��`�K��O{&��sO:D�YF#7ypD��@��&h��+Շ$D�X���Q/FE��F�/1�$�v�#D�� ��^�ϐ����	k���ie	#D�(S���-A�=�j��fJ���B,D�(�kF�E�t�pf8M���0F�O��D<�i>�DxBe_�dޘxP���R%�(�AQ6�y���<�=J#n�P�|�R&�)�y"	L�()V�����Q�"�_��yR��>�l�f�A�w�8!ׁ.�y"G��x���h�-L�zO�[d,�y��\�)��(x'#pg�}��L��yrb��hq6P�c�g��͚�	��$9�S����lp��W� ��yCB�e@p�0��$D����b͋h˾�	����g2Ae�$D�`��H� @��h�I�T���hև$D�Q3�>I�$�R��<'>��'�#D��0dH��Cj�5�r������7B6D�HV.��hĴ�"%f�e�<���&D�h"�ԣ#�e��ҕR�Q+�-�O�=ͧ�O�m����H�r)[��H�6��1a"O� �R�%D�*�Dɱ�D0�>up���Ɵ�D�d)�*V,@9�R��D�� B�Ý�y�`\XK����5l����&V(�yB
�$�5id�������D��y�g�1����'`5�@�4	��y��"=��*"$��[�^5��ӆ�y�IN�V5���'`�(n���i���y��U]6�����"Vn(�镏��O
���O�b>�b�ψe��td�@:�Hi	O)D��P�ԵWp�e�J_�`�8�!��3D� �����.�2�Պ[�E���rm,D�P�r#�=>`��Q�m�Eܸ��J,D�b��YJF���ϗ X�r��&6<OZ#<y�Rf�H�⯒(l�p�F Dj�<�"�īWN�!"�H� TP��X��f�<�m�:zN$,�E�YO>\uKr��c�<	�È�=T8���ƗiZ:���a�<	�	��D���7�ߏG������G�<�-������v��a����F~�<i�Cߟ(���F�%w�!#�@�G�'�1OV����#�z܊�(�`	�pJ"O��%�=bl�� ��t!�̃�"O�)A�O�
k+P	y4/�".�,1�"O��: $���H,R�CD:�|���"O�9�Db��c匄9�(��'�DP�G"Ot)ffE>G� �ӤgN�0J a�"O&D��)bV࠘�Ɩ	6AS�"O�q� .�4�EB^�1�2"O@����0-���
0��K�<�"O���b4^J�<3uH\�+6�l2Q"O �АB��Od9+��4��"OV%x��Ҩ:�,�&g�
l� I�"O����kJ�8��f.T���P"O�,�7�B�#��a�!�� |BV$q �'*��R�nF�f���a@�:�d��&D��HbLM�A�\$)$��S͎ [vf/D���'��/(�p���Od����.D�@�q�ŬUA�i���L	�v� �.D�T��G�&��:�eJ�4��{�+*D�HCQĄm��Q茴:��ܒ�*O"H��,ąV�0H�Q�2�X"O�%� �����fI���"O ẗ�OײhC�e�l�DX�1"Od��A�L�X8��s�S���k "O�8s�G�SՄqa�cL�XE�"OhI�4� B�0��B$T�6�!�"O
	��NH�N�y{��C#:�<\+�"Od$���tEV��/"�R%p�"O B�_J�x!��I��:"O��
3	ډ7&@����-�ni2`"OT�GlV;\��)���@�:=�R"O�,�� �l�Q��p�Pc"OD����U�j.V���k�?r4��"O�4����  Ѱv��f�W"Oz�ό8�T\�D�+GL�z6"O:(�rثm� �x�&�r7vh
�"ON-�QAϖ*9�p��%��KQ
��"O$)2�Z�-W���*�<s18��"O��"P��'b��1�''�N!>���"Oz�b�½F'�Y�#G�;9���$"O�T�����?;,�Xg&�)_6��u"OvPx�&�,�6�A�� -,wB�"O�����ւ
�T eP:5WzQɣ"Ot媃I
V�x�	�*���"O� ���dm�x��@3cU�~zFm�"O�( ���?
����"a]�Kv�ç"O�m�L#
��` j=Ҍ��"O��8̊2��#�/0=��"OIpg��آX0T(_�S*p�+�"OP�{!���"z�E��>"��V"Ol�+��ɎWD8�.>k�E�B"OB9h#��	t�՛��LR5���"O����nɼ*�rp�"�AZ"O.ɰ��V�k�4R�*L\(�٨�"O2PY �U�C��D���&"x��"O�z����6�cB�L�!
�"O�9��d
�Ȁ5F� &���)�"O��"VɎ�K�.�Ӥ�$����2"O�P��&S��$Hj�V����D"O	 D��M�]�T��L�
y�r"O�Xc�K��c6<c�n	!*%�B�"O�@�C
�s����Q+g����7"O������x	�aY')I ��!�"O��+M;H�4��6n����"O"�IˀK��Ie��^,R�"ON�d�4D옽�"��q�P�jF"Or�-F۞�YŦ�� ��y�"O ��^/aa�5�gе��eQD"ON�2� ��C-�pЁvsZ�P"Oz{el\�Ai�����a��)p6"O����6̨\��Z�#�d�Jq"O�P��J�=r�d�`�ꀡSy�H�"O���S��63��P�J��Py�4��"O��X��ɰm�<���Y�$rri�"O��2�,4G?�t�4�L�_���$"O USv'�W�J0��Y"�Ȅ�G"O�S�	�	 \�h���_����"O�m&NF2⪐ѥ�ߟY��[�"O��r7�I�)�.M���/;����`"Ovr��&��l)4�Z����"O�!���Os`�
�$H�r� "O��1A���X}�f�S!mHĻ%"O��tLB�'�~�S3��=T��"OxԁM�Ơ����jɪF���y�E���(�A�	.�X��gO�y��H	w*� �ۡ�Rh�v�]��yb*YR��ш]��:� ���yr��=.��s��P!�L`2Fm��y"��'#� l 1��u!ȵ	V<�y���(|)�! ��n��2�G��y2[�(|�����T�~��4c��ە�y��ѝX����{�Ԡ��C#�y�ܧEF��C F� �6�j�k��y���tSҘ��KM�	1bi�,��y�$�Yh�|���Ơގ�BTD֍�y��Ȋ$p,��G�C���dA(�y���Z2z�@J�?����� �yB���
% ȱ9x���n�,�yB(�"3e*9`F�Ҳf*6r�$�
�'��j�f�g*�Z�G�N�d�;
�'4��P*ڊp�v�+��<J֑
�'9蘁fh�	V��	c���A��

�';�P��+g�*��=:�*�'�re��
��y�U�T��F�x�'��(P�ʁ)�v!�P%�o�����'$�)�#`� .����A��Vi�t�'����$�]GR�p��;�^1c�'2�S�c	�T9��@S�S�
L����� H�eP�$X��@�:��"O^�:���J$R�dZ�I�\��"O������~*�:���T�ѥ"O��#bp���ă:u⮨[�"O�e��������c� �x�"O����ʽpM`H������|t�U"O|}�oϿ*��T�AN��IR��7"O�4j:f�P��@7Ny�u"O�$��Ɔ(�HX+�$��v$°!�"O��(���+���&�G�v�Q��"O�-`u%F7;6�X�$�E19��"O��`�g[`������l��M�D"O��r��I3m���ӅC(cO��!D"O��2���+u �+��ֿ�2Ds�"O���-�&u/�p��ԏH�l
"O��A�*M�j��s��5D䠻�"Oʅ�g+'�J��)�a���v"O }�F\'B+�Ś���#$~ެ;""O6�[�)��59<lk�%.nl(J�"O�-��m%Y�2 ��zU�� R�<���c���*r�8evP�NU�<I�aȍ��B�rkb��@��,n!�Xi�����!l�hIDI�al!�$I�@���X�l�ee��y_!�d��N4:'Nt�d�ԙ U!򤚧/�-�d�F79**4�3���=!�ў!g����o����'x-!�$Nj��Dcf�:e���2bԲRp!��|S��
f#��y��1	��ш�!��?c,M�������Nҷ �!�dP� ᚄ�5�[�A�>{�K;D!�d���|����L��t�l�0!�d��tn����x(r�+wJ��u�!�ů\
�̀@�S�+���I���i�!�D��u^�	ʥ��+(��X�>�!��&12hy�8r�
������!�d�(Hv�C��9�FP���pw!�D iY.���KW4Y�d{E��hr!��J-��h�i�*u�+r�[�)�!��(^2E˥)]�	���8����!��(�$
��X#2��X�d�T�B�!�$��4���
^ $l0C�7|a!�d�����Qi�s|���"S�}C!�	@��ȳ!��F���u�ؗ�!�d�c�@�S�N�x�ZL)�h05�!�6&L8,kQ�ȝ|��U	w)��h�!�D޼l�6p:c�'t*MJ�jX�]�!��]""7�����<>b6ذ�҈d�!�$V��:��$���˕,]:H�!��˔y�mi���FYn8aUe�Qv!�$�3|�~����{W����d9@!�]�6=���כC@�H�d�2!���0��AL�m��Q��͞�!��[)+��0P�d�2�9�6O'�!�$\�r\�wc�)2u���`_,�!�D��eL�D�b�\�'q���ñ+�!�$ .6z�֨]�s�b�(R�3M�!��@��qǄ?-��F��7k!򤟚}�@tj!EOr�pe�	V!�d�l,��%쐁u(�K'W�N!�D�1i�^�'�9p��Yh�.d!���<�~%�� Z�F�I� Gɕ7Y!�ĕ�N�&����^�]���k=i�!�Ā+�p4y�b�;S����[,6!�� P�Y'mT�(i�A4�z�J�"O0�A���	N*��R��U��x�R"O~(M[*�<1���q�(-R�"On���t!���cf	`�4i��"O`$	'HT#����֡w���r"O
dzA�J�^�,x1��i��"O0ȓ完>"�JP�*��Es"OB���I#V^�(i��sG�� �"O��St$�P�F����2a,f+1"O���b�N�V��(xq�ϊf%~4�F"O�	��L"&NJ(�O4��{6"OX8��FK�6��9���+�P8�"O|i��ª.=`4�F�;�$��#"OLI{�H�����̕ �$��"O�|$�S"~5*=	�`:�Ġ��"O��Ӏ�
<�tM����(��"O���B>#.�=��#�1�:��"O�}h%�ȍ5L<"C��3
�>��"O@���N[�b�x��#B�rހ����'8�O�-h�-��iP�p�q�M�H��|:a?O����	 90f����0@+V�[�@n���Lb�	�`,��ʈ�aC���5.� .�FB�ɴ@}�,[�	^,sp
4�m� |��B�	�<�pX@����?��!k�oI�-��B�:+"�Ђ�F1&��A�afB�]w(C�ɏpV��[E�HA�0�����j*�B�	�k���A@˞�P#�۴_�0��ʓ�0?A���=��A�E_��S�b�n�<��T���r���7�H�@��f�<!�E4v�,����'��ᒄ��e?����$ɧB�h[�蓧(���� ֱB�!�D��00zehT)�!7�h��*��,��"=��9Oٚr(�l���#6h��*>	�"O��f �f@չC�ԃ�
<"O\qR�@��L�ڷ`�:q��Is���	:�~,z�Z�ؑ�k�<�!�$��L�`�e�	�1�ށ{�*��!�տR0SU��<f�F�P�K�!��Ŭt<��T"B� �Q�D�0�!���V�����k�3St�ur7J4z>!�$בO<-���2Y����Ѫ�2
,���Os������/ 14&�2��C�"�p��āʡ�yrlH�Z�0H�Q
�H����`���-�Oɒ�e�(<=�p���$
0�t"O�d'�v`�8�f��$��ʗ"O`,Q�M� ŀŢ�11� �5O@� ��Ʌhry+�N�xR�ݐ&(5D>LB�	�?(���c�~�9�([��C�ɐtlI�Q@�$4�������"EsB��.XT<U2�'��9�j�P���eb(B䉆#͠�ݜ��˅��}F�܇�I*!�h�S	�L�x�
����C��+ �$�@����>�1!�e�7հC䉔��	��
<iv�P:g	���2B�I�<.��d���z�+�]��➜F{J~*��S53N��3���HP��+NT�<��JШ\:�L� G��>�pI�1B�L�'_ay"O�$���P�U�P�N��M��ԟ0"<��fX�=px��䆥f�6��-�G�<fj�xjZ�csڜS�|����E}�]�4G{J|�r6��z��s=�h�r@Zz�'�?iW
	�hԔk1.M9cZ�	�:��W����.K�*y!�f@�S-87��<\��hOQ>]�F�ݹ ���*۝A��X��3D�� ���0�ӵ��h*��vc�]��"OA���\�.��� ��F���"O�@����5\?J,�2�]�&E �b"O���B㍏=N,y� �.Y�XXS�'kqO�0�˖�v
+7��Tb�	ޟ�E�ī�*���	paQ	��y �����y�u�䒐�ε8��Dk?�y2�{�-����o�%Y��M���$�)�>��M��[��̹f�L�U�6I�$oGUx���'
�%8��Z�"�|󗨃+Yy~Y��'D���d��, ��H��1W�@I�	�'��(�%�v#>�Sqf�<@�y���hO���U��bH4�cϏ0hV�{�"O�[�"|�rd�� TK�B�"O`��-N�~�E0�y1!w"O�(�Uh�;-i�D�aW�wwt��'��e��a��@�:�)12m�=������?�w&�)�N��T|0��YT��P8��Ez"��Xy�{ѯ�8*��c�!&�0<q���U�dG���fcH!u*�a ��E�>z��hO���f�6;��*���i`"O��+u�[�T̮��m�.M�� "O
d(�����Q�U�P42��S"O��J7$��J�$�9H�w~���"Or�S�aʌ
;��	F���7����"Oh\��Ç/5240��!�17��×"ODx��эM}J��AI�έ�"O~��uM�\����4��MXq"OP����8 �&�8��� '�8�"O��q2�Q� (���ֵX$\�A1�;\O$�(pa^�f&���G��*'������v�<	��������:�����v�<yt�	(bsL!p&�'{�V�[��o�dF{�N#	��Pգ�9B?�8���Y ��'Zў��<+h�^�����u&�	�5"O�M�QM]�n��)I�L7^#^@�v"O����'	�x�"6�ߥ;�d�K�y~��'R�ギۣ.��$�i�\հ�'��}p@��44ޅu�T%	m�<�'�^I���1�5�kW�S��y
�'��mc!�ˮ$JX�`k�
?y�{	�'��A�#�PdE�)�U������'�^qScB-$�.����ƴ:��H<����!���J�
j����fi��u��^O�H�� Y��H��D�nnB�ɉ6��iG'r�0A�f撕&��܄ȓG����M/��]���Զ~���ȓ6�,�pqE��0���6G����'��Ey��	Ρ!*���խM�L�2�k�<�O�%C/�s_��*�KKuBʝ��dk�0�=9�5�d�-p��Q�ŚnL���ÇH��d?�O �3 ��&���OB4kV�1��O�����7 �!��W��dE��C��O�!�$:M��-#���pӖ�a&�(�!��ߖA�B��w�ɢ<������f�a{����5V8Qx�F�f����Sx�!�d�Xk AX��� ��HK��I��O�=%>��4nǡoÜ�S g�9_���p��)D�<����Q��`�B��B��%D��3!,O�~�d�kM/b�-�gB$D��+�ѹCd4���P�a�t,��'}b�)��"u�|�[ �J�[��Ī�5}9)�����O�I��Z�����L=b��\��"O  ʷ m�$���`��E�>=j�"O� �Г�T�Y���[�J6z� �"O:$�u�/[Ƣ��+[�J�"O���`��.o�6���k�I��qR�"Ol�8��~��y�!��4���ʔ"O E�w��eL� �g�r2�"O�CbBN�M\R O�6if�=y�"O��&ÞH �@�2BrB� w"Oּ�SbԮK��P$%	�WZ���'��$��PAH�jԮ�i�d0�����	p}���S�JH~��G�\�p(j��P/G�n��"?Q��	�L��-�d�;k,2I�f�{X!�D)h=x!�.Z��|��]�!��q��(�4��g+�
K���R�3u>iD"O��@�K�=s�ۀ%�����d7�O03�K�)�����ΥxK6\��'�L�����`��`�BI� a��1�/1D�XA`(�06�4�agF8?�TI��3D�� b-�����3t'E.`��	P�&1D���hЪ�i �$|����$�,D���r��X�b�Ӄ��Y@� D��{elBTp���.u����3|O�c�d�A�H;�(Q��?b��*�l,D�x:r��s�:�Ɂꓝ\�t�#�=D���N�V������S�!�8��:D�|�s.C�	Ϧ���O����
%h$D�|�Uj����O��$�O#D���P�E��,bEm��X���(&�<D��93N�,]�g��d|b"�:D�<I&�J�WX4��%~D�s��8D�t����#�`"�O�n��Ak�,#D��C�K�c����bd߈\��%���4D�\0��%u��=b%�G,��c��2D�ċ"�ɻ\�X�uG�;,|�2f;D� 0Ag6��q�d焠(C$�"O:D��'��Z�e=V���Տ4D���4�K���)Sn�=��i�N1D�l�%O�?jV�O\���Q
f%1D��y�=�z����� ��g2D��#��LO��sw�W1	^(�a �0D�XIed��m:��R�{��Ab2D����'X�
���a�;v�d�(�.D��1�e�>l��2͵r�����,D�����li�����"2��,.tbC�	*�M��M��V:Bi � ��>C��c2ʵh�.�*LXޭ�tM�N�C�I�9�"����M���)�7�ܬ��B�I5J�K���6$��ڢN�u#�B�	n��}3&�P-Fe�PX`�؝��C�	1S�}u�_<q�}B$K.3��C䉃a�����g
)�e��ܜw{B�	c�Z�bTИ8�j0�#�)��C�	(hՊTA�&ۛ4��U7:��C�I�N�^%�2+�G��P+r/� hB�I5+��q�sMH,9�u�IӁI�BB�	�]�AK�*פ{R�CE�L����:&�Z�F
�nn�B��ƿq7�8���@5m2ȈrěJ�!�dԖh>,����,+/n�� iAc�!�bK6Mf�4]�A�P�!�$[&7���¤W9k��%�c�GQ|!�$W�+�X<�g�R�*g���W>Z�'����/9�i��䌆_�Fh+�'�NdP��҉q��-�a���U�z��	�'WT�Q�xlܠ�Т�}6�E��'��xfh�!��`�E�ԘC(u@��� ��
f9�
����͝Q�%Y�"OV�eoɯ
��u�Q��}Ӽ���"OV}A�B�I���K�oO����"O���A�]�|K
U��(U j��=�5"O�)@��v���G��x�"Oz��pbY���Tŀ$pi`"O� ��^,S� [ ��![st���"O�<���sy�X@p�
3p���W"OҼ3b�|����,L
�,��"O�]�^�0�h�C_�e#^��G� �y�H(���#��U$ĄK d���yR��<�� g�	7�j�d�ҩ�yR�AN�"X��L<y�|B�M���y�LC~	�m�V�I�"���`$���y�����	���58,X ����y��-��iج
�4��4hY7�yB*՗}Y��A�3R�𓭔�y��EP�P)i$�M�5�h)�b����y��V�4m��d��9z{����K$�y�I��
�(��-b���yc�5�y�&V�	�p��1j� Y�́�7�yr�ƤR֖!ۧ��?S]�xd"J�y��KF|(��G�_;E��OO�yR/�,��#��I�B���x��ˋ�y�gW+�h���YF���A�ʤ�y"��*m�V1ʧ�*�������yb)M�z��V
Kx�zw,	��y2$��e�d���`��E������9�y"b4j��4�蕶KR�TQꂢ�y�f�!U����ŧۡi*0x�hA�y!¿V� abY�{f�( $��y�C�:�� B ��{�t���	��y��X<�v�2+�%Z���Ar�-�yBG�6iX0ȶ���[e��&A��y" �*�����CRTjZfɇ��y�+w�$2�+�K�����y�		�x�Ȝ��CƚA� ]��^:�yRrW�0����=G�@���Z��y"�Wa��92��A�?Ǣ��R��y"
�2<�*T�2��5˲��y�
�6n��r�֯_�h�yr-�y��
^���/R��C��Q��y��Ԫv*�D '�E9v�����y2#�9Pv��dR�O�$���*��y�k�(�q�V w�MЁ ��y�V�aQv��a(�/=�`+mȢ�yҫn0��〆X>8�8�-
��y��G6HT�3��TIV�ҠBJ#�y��ȵ�q�e&ז+2p�V�y��Z�=F�����;�� � a��y��#>��PCAk�]q��z�GD��y�K^�vxbD��ń�#*���N,�ybď�a��)�e�9nP��2'��y�DF�~��r+��d��8�j@��yr�E�D
���ń�"���!I)�y2��*X�<��k�_w�@����y"�ն{tpB�P���Y�,Q��yFG��J\KC��!@[.���Kޢ�y�nW7v�0�+�N�!G����F���yb�����"���~��"���y�bC5ݞ�+2�^&N04��ڄ�y���!U����W$��N��̩!��)�y�D�22xp�5�Y6qk���n��yB���1��N�i��ޒ�p=����s�)��h�� ���%I"�Nz���<4�0�I"O���#L�؈�Q�+���
������*��c<��}���	����Ξ�yW�@a�F�<9�(�z)иKd+	��~ �
 �����ͺE��� =.^�?�'[����.o�ђ�e�Ƣe��'W�a�eΖH<؈1&�W�*�����bV�D�d�g�p݄�I�!�,�H��(��Bv��m��󄁩��"�m�k�aB蒠Ts�a�a
�4�JaQ��47��B�	%,���0`�k�~8��#%��Oz  pG� #�l��K�2e��uC�/c ^T8�C=ٰ��$�j�<Iwf���Hh�����5�*]�5��rk�(��E�j>�\HC�R5Z~���O�h�gFӓb�L��Z;n��O��HVgn� ���,e���E��9:������p��ܯ^�|��Č �عqt-�o4`(�����1�牵!�͸���'I��R��D.�έ�'[q[�0�)�	ɂyؗO0x���ݾ$��4��J�Ș%�$O�ܸu�C&���B+�C�X���d�T,��<�W˟U�44��1��q��YX�8P�g��E�h �H�U�!�EEM�7z2�F���7��4����<n���8����|m!�X�I�|7m��q�-p�\sU�I�?<�	r�P.rgay���,s�<�����X�HP9��>��и/���Ԛ-S-BP(�$ڦL��.��yLC�I|$<�����<��K���K�D���CZ�'�Dd`��	'Dx�Z(A��T"Hˤp���:�3��'��U٢��i��5oE�v�rsl(����]��	�z��s��p�h<���x���'LU�2�O��qY+����O�ƽS5�P+��Ȑ�"�9ˊI��O$ձqI�q ���D�8��$M��f��sR�;ʌ�(Ac܋��OJF�0���6ݑ5OH�7	T��"�(70@ߧ7�B��+4a���V[b�:�>p� j�&�*m���!���K��'o����KZa�<ҧ�T�>�f��qK�	��xh�N	���<�V�/�7�Q;$#L��t��6��$ X(#z)��� !r�He�K��C��RRG�#��)�'<�8ȳլ�U2��d%]�l$}�K>�T���m&y��=Y�RhHCL�˘O�"�j7�[��BD%��0��êO���G��-]���'�IzdE�j��1&��(@a��P$FRN|��۝Ae4����O�vXYpJy�0!����ʺ���$�?��"i#=n!�$I�����$�;x�y��V����9H����oQ6.�s5AȚ�����zy".UƼ۰�Ԩ-�j�S���K�(�ʤ�B��t�
R�Omp�0�)rvjV�5qĔ��+��G��d�0#`�``�(
��ɝ_��Q��I�**� �b۪fI��j�`P�K-B�25	�	y]F(�f�4V˘Ћ����̈�tIG ��p��4��J�'�~�ȸUʴ����<�E	ѝ;�`��B�q���߷]���!C_�3�<`�ߐ?�u�}��/��ɚԨN+X� %c-��V�����/`JpC䉂ztb0�͙�rat�P�t�J9�GGցA݌Ma@�F@�A'˔�p=(��8}���#�P�.�Z�*�[ :#
���GͶ%a{RD�tR���v��">Q!k�BM�����Z�����02,Ԍ�P�ڜb"�'e\�)�A6��Ol�2M^��49��⌅z�=����@gʼ�a�I�~'ZP�dB�1�O�r�""O��s�`	��f�B�
�[�OV��W�P�5yj��d�.`� ��E�����'ҔG�����&�9�F�8��|z*Ay��Ϥ(�DE�ݴ/�%��F�>(�Ha�@ jTDĆȓ?t°A`��+oi�P*��_3d�s'�cV��6��D�y�&к���(F��(�P>0w$�
5dʍ�a{�N�P��l�`ղT�p-�׊��6d��0I�p��V�� ������'U�D�e$�m�(uK�?	Ŧ��,O����O ���2|1�Z*BFтM|ʥ,Ρ
�~Q�mG�l`$��-fX�@�G���N���D�B+_2F�~�p���)r �@���D�>��#�떎t��:'B��h��d�9o �L�Sd!o�`�rW�ˀ(���Hɔ��E�>��f�ԁm<����G�x~�ӧ)̟�Ao�r�� �<���D�mX�D4�`T�[��"cי�M��I�"���M &��/1B��!!��=v���a��&d��3��:,/�Jt����
���4mD��L����[�A�8O��p��Y��![4!��O�nih3�K	w��|�!�/3tU��Zh��v��O�B�Dϑ]S68`V�[�aゔY�'L��C�g'��O?5�'&\l*��� �z�fl�G�'z�Ѣ�3� ��i��J>�(4�t�̹M���rq�>a6�s�b��d�- S�-`��� ,�*%�!�d�%=DZ��R�]�T�Ib�H�>�!�#LǼ�(ǆ��;�t�&H3i@!�$��}�8�b'K�P]���Gj!�$�80��(��ܙ]��%��c�*1T�'��5����i��@1��D�z�d��"�4I!��_�p<���Ֆk
M�'���U7���1�+����c��u��mL/&�\܋g�C	[���ēfڬ �6�C�}4�M�NG�/J��v�˲l�8��d� FEfᄢv�x]�#Cېayb,�B��&�,�2�`�n8�G�
&�!dI?D��鳠Ȫ_�1"&�W�4 ��k1�$��Q&|r�{��D��5q�dIvLX_ሑ��J]���O�Tc!g*�'#�r%Ò�8$̍�Lݰo�� �{��6G�zb?Oj�"e�>8z��2�@�M͚��7O$���G.���h�� �����U�P��U�E�&��D2�˲hLC�ɿd�0t9��ۈf�
���T�q�t�ʢ9�M$\OT��u� 3-,���NB
+y^`!�'+�<r��+"pl�Q���]�M��Ҷ,#^���'����-%�V���?-�4	�����0{߀Ġ��)�p���T �7}}�Y�Ú!D!�D�'�̽x��И.2v��eT�DI�
T� ���{���P"|���Ӈ ׁ�xB�C��@l!�䐳d�N�H�&.�|�P�1)P�M_.H�
�xd�ia"��J��ؕi�3��U��8���r��N�Y>����&��xɄȓSˀ����U�%V~8Z��Q����ȓb�A� ٱ�4�$oM�"F1�ȓ#�tʦ�U���z����yr��7L6J��1��M���	G���yB�Ü%����窞(Ct ᵢ��y�'�2�����I[�9�,�kE
כ�y�k3G�ܰ#��2�*�%���yb��h��Q)ɡH�eQ�4�y"�ئA:&�Z��� (��|���G��y�λ_GH�H�*ɖ&2��b�^��y���y�2�B&H�#fE4�eӱ�y�i֣D��� �b;������y2���х���7b��z����yj���ȓW������7Sl����H%�&M�ȓ%>��Ȱ�#H�\P3� 1�!�ȓX�V$�doɭ�8sWE��b$����(�Q�/��:��>~�H�ȓ_�*���c��]�L�bGU9Oj���7>��'���`h�lZ�LKz!,���/��4&Րj}�D���� �����x�A��.]@>�B��\�
�ȓ_;����x�E�a���6����/jB䐴MʂA)*1§hǤ_�Tt��K��أ�jP�V�"QX5��.xԨ��z0P2�ՓW��Ux��[�� ȅ�l�p\��JS�C&N �Q �܅ȓM�I����/��'��V�b��S�\� �(�
=A�xBR͚���x��h�x�A�dٙeX4��C1}���S]�f`���A#u&�(tֺ�ȓY�x��jU=*׺��Fb�(To�h�ȓ���1��Z�R�k#�M�`�,Ň��*�9��4`���"����P'����c44�P#�_��@z�*/}S�!�ȓ!�P4sd�Ȓ��%�É3AzU��E8�(��	!t�@T#d�z���ȓHEj��'J^�#�B��UE�?�ń�S�? vE@!n�^��-���+��lS�"O�P���C0P�)xeL�M���"O��ѧJ�#D����²+9�\#"O���v�"2t�P�b�2,>qh�"O��B�o�UX�Xg���WN��"O�k��M�`deXS��:��Е"O��,E/X�����gX���{�"O
���!{֩b3�"yƅ��"O���k�<;8j�0�c�I�ك�"OX��&)�:���q◆\�Ɂ"O84	��9��ܩ��\}�U�7"O&��cJE�W��)E�6IT�1Q'"O���Ơ��<<��J�4 O�"O�lA���~3l� �KV�1,�|�"O���z���!	C,#���
D"O���;0�X"����є"O8�0��8$�} ��^	'��	�b"O�PA�K--�4I9���/�84I"O&,Bwo�r	<@xb�/`�4*O\�C�ٷX�4�J��� {�ޕ��'z"! ��#����P�T`'ر��'��#�j�y=�ب4��0XF΀��'�bB��:����#�T+��]*�'V�L�5��!A���j�#n�9��'>Z���I1C�,�[!�j��<r�'�p����+|�*<���>P�|��'֌ ���)X���%D&D@T��'�9�V� 3��s 'V#'��
�']pq�@j�����2Z6-��'�:��v���b�@-�fk��)T��B�'�0��d�4��y��͍;Qƪ���'��m��)@w%x�`^'N�	�'�n बؾ?,q�����݀I	�'��방"�&ɲG����z	�'r�D�'A�;�L��@����	�'�=��c_"D>2,��/�\���'����,��u10�)􏃕_���'�n�
��W5MV�e�C�C�T��L(	�'� [WŞ�UMH@�S)\*v�S
�'Ln�v#. ���&�.r��z
�'슱[�MT�G�5��n���bi��'kB4b`�#$�\ �PJ�P�'4 ���VT��m1Vm ���'R��g*LZeTE�����A��'�",�Q"��X�[*K�V�D��'L�,h��ɮZX������
O�!�'�D!�l��� ?�A��'��a+�� IaL�ZM�6��' FlcD��!��1Q��D�9����'Xx�Qġ�*����@@��3Q
��'[2���ًRb�|؇�U�{1ZU��'����&�2S.
=�F�ο	����'Kx	�W�!W(���"C	���
�'游�u��-R[NP�U&�U�Z�	�'�)0ugY,�ܡ`�52FZY�	�'=�1PġD}�d�V#��.�E	�'倭1Q�1-��T[���Vx$��'_���S�$Ԇ���� xj�5:�'�sq��d`Ip�!��Ȫ�'��!��"R>Ei)0���.N����'��Hu.�"@�� '���@I�'8��`�����W�EM�C�'T�z�D�e�X�9L�&O�fm��'���+J	 ���hňMnA���� fC� M�RA� �tջ���"O*٠��{�8 Z��e� � �"O����;�����C�0}A"O*���D�#T��MQ��@��y@g�'RС00�<h�]Γ!��x�1� �f�\�@� H8NI��Ͷ���L� g�Fs�9g_v��<	S���eZ~�ـ�˸�h��H�rm"X�"C��L���"O�+�f��r`�D�t�ܰX�lep�Q�Ah�UWfd?�F�����	)FĹ��*���$����bC�	8`�ٚp&ߩ;��%P"!�3#� �"�m�m��J�'a{B(�80��q3��5�>h�u���<!�I�7�&@����1���C��
4�q�L�p�T �u���y�'^�-�����#����MH��"����'�i{t�����==񟪀@�OӌD�b!�B�4�Z���"O�����/̼@B��	8�.��A�>SR0��"
'!����O����&��ņTc0c�bT9|�tهƓ8j�8���R�(<
2o�'b#�k�ƈ�8��ayE�á%�2\vB1,O$��LD�&����h8�-f�/��<��eL
k?�5!-q�x)S&�YSI������*d;��3�i�d��C�ɛ)ϖ����W� (���	:�c�8�dS4>���R�X�-QrAQ���(G�j�X��+LRYH��D�yb"���U��;SL�S4&Z�P$�Q�a_�21�c��O����Y�|aӍ�*3lR}:�C,&M�L4K0D�(!dF��"���ju# LN�X,�<�&kՏbL	�"-,O�ؓ�K��K�Θ� �\���`%�'���PU�K<*�&%H��G�Y����_��R!BH<�2�d��5���6�6�x&�G�'�E0Ɯ-8���҇+8�d�h���|'�\@"Oʱ{a�K�vLA�غu�j��O�T:�#�����h���c0�eݘ���߁cc�؀"Oj\�i3[j�u��-O"[������R @���	������	�0z����̯�����L/��Ma�H��2�H
�#$=hU��
��ٳ	�'���0�I�;%�-���$�FIZ��$��&"�R)N��O�U�ː8G�c ��$�b�'C�J��YSP���P�ʩ9r͓eߒ=P�eʘ�ҧ���]$n8 ��Cq�A.xP���)<D���SB
�vM��n
����0�>a�-�4q_.�����EX����*#4e����ڶR�ȥI�B9�OH}��c~��2��-}��e�fg
�m5d�Ƌ�:h]C�	�޺�a���~��BD-��~~b�<����Ԯ�1G ���O{�؈���k�
�5�[,^�����'a��Q�!�_sT�T�<" �&��F:��g�R�B�S��?��
�kl��2eF'EP�lX���i�<�Q �tl�Q����A �40&�c?qso.
%:Q��qx�d�D6v�(	YP+��_��	9f'2�Ozaʇd��N�y1�Sd�5�w�]/5&� r���y��K�F�2��`�ӗw^���.ڼ�(O��+E�ʹC�>�È��R߰ՒD��8���,�C�!�$û��b׈ޫ-�aa�	�:2�+AiQ�u��ʒ�>E���8מ�B�T+T��D2��I/���ȓ$�0e�!n@G��0�P �8	�2��'&(�$����zr�F<��%���ϬC��-��M����>���
Un6M��A.��Sm�I�T)�*¶P�!��QKeĭ!�0��O�FL��'����M�o&��;���?�Y��'���� 97����0��
�'>�!4*�5F���biRd�����'x�qi6��`�$���O�Jm���'w|�[sӘJ/\�w��<��	�'�<�P�U�=�� i�36"�z	�'�ZpP$��1EP�@ՂW�~����'*<`��_
�0NC�m����'��t��`�- 2B�(1���oÐ!I��� D�31d�U�H�t�3�Zx�"O	��c
l��b�C�%��)R"OX����%��;�cPR�΄�"O�5q��L+~.`!pAEN��3W"O�dxDdأ ��h�A\�b�ĲT"O�d@�3L� xh���4����"O���F��B�ԂQM�+U9H���"OpI0ף��î`/A�P��-	�y"撟/��(f'Wbk������$�y��\.%]�%+T�]�I�Ej؃�y�],=נ���J��P
bYô!A0�y«��\,N}(S�D1B�bq�k#�y�oN�\@�f.�'NN������y�Lâ|^���f�3D��0���.�y򇝐?���(ҭ�?�t��ɂ�y�>')�4�F����K�ƙ��y"�ȒKI��xu&�I���l[��ybN��}jt��e ��B��8;wGD��y�Ӫyx��&T82`�l�y"�T qY� �)$-,��E%J�y��K�:���V�$Լ���!-�yr��?!��+�fD�
K�ؘe����y���n�݊��ăxق����3�yR#�	I9��)A��n��_/�y��<���.@�ʺ-!v���y��߄Q��� UZ���M��y���i�ȭ� ��G��5	E���y��h�|���g��8��෨��y2�V�p�ڑ�d˔� >D!����y�O�C��s�	�i`�ۖ���y����q_��R!I�!n%���h��yB�H�B�����"b��h�R��y2��3>�ȹ!�l�u锑k3�܇�y$��)z�q�"�O92"Ή�b��yB
BQ�=SE*ǔY�&hPRB ��y�F�}׊�pwf��V����&ㆴ�y��Q�4�� ���D���Z�o�3�yb�T4�y�DU�L䘀��'�	�y2,I�-�Pċ���?�lh� ��yҏ� g��P�$`������y���wT<�Ǩ[�}vɺ�eA��y� T�$[�	ԗ	7���Hߗ�y��T�Wl޴Zj@�YFZA�E�A��y� u�h ���Z�c�FD��3�y����������^��ˣ���y����Ȅ�,�� X�9C���yReE�JHb,�1��q�����K��yBJ�;N<`E�q�*zcEʓ㙶�y�Jק$Ǵ���ڂp�8 � �y�!��+_�P�hpY`F�y���R�3� ^�AI�x�7�.�yR`A,s?>@�0��6l�H�i�-��yR��F���,V�o�F蜆�y��Ɣ�i!C�(B�r��W��y�k� BRC�``���"+N��y"@�)8H�򲅘�nT�k��P*�y�cN3��=ʂ��q�D�%�T��y�$�\�����	�*>V�9%E<�yBb�v������bt�s%�C��yRGɁJ��`�߾d��(at$��y2%��D�t��A�_����8�y�1;8ԙ��oG�Vi��P.���y�EIP�.�P2l�8u�$b�\4�0=a�d�=Jp��[�(EܼjqnȒmkmjƮЀ����_�<� �,zƃ��!$�!A�Ƌu�Rܺ$"Obm!Ǌ-7�H$�ΗW�t2c"Oƙ���<�h�ul&~*�	R"Oj��a�v�t�_�:�	�S"O����Ct�$��J�!�2��#"O��0�!J�s���!�I��p"O��bg�T
܈�CU)���$�IV"O�Z��K�[��H�T(砱��"O
��[!(C���GK�W@lI��"O\P�VN� 1Fr!�)K)>,�5#2"O�@T�
�;_�Ƞ��,����"OS�U�]���W
�#�2W"O�@G���rP�Y���<�&�(��'y�ov��#�N[��|k�*�>bT@�v'Y�1�y��	 2gh>E3���2����[C�${�����	78���'>�ю��oO'fg2�� �ua ���g�|��pjfá�y&�-~|$������tM�oB�%�B �e7flZ�醓A�vM��O�,�!C��O6���S;'�a��E=l�6�J1��p[��,�e���
Q�
�ӂ�O~��H0/��ۖ�Ue8	�ڴQ�����r�Py+O�?M����`:�9��h�(N�HՉ�4z�=	��ڃ{��IO�3}�O ���m�?]�.�[V�%<�$ �ڴ��"~n����)V�Ixb�Y�bP�vtB䉤h�\���'b!h̹"FʲW�dB�I��� aˆ�m0��p	ǅ][LB䉸^g��8f �A�e��X�B�B�ɏA;��3�&�?hV��g�T��B䉸��q%�;o����7-�$u�C�ɰ
q\(Z�V1kq��B�N�K�C��R���g�NGJ@	%E��B��=s2�a��0
��"�9���d�0E\��J�uK���A�P/!�$]}Y��1щ{8�x@��֒r,!�DB�~�|���&E�,���nZ�e�!�$',��XyFȝ�1�CI�3U!��"g&�jA�֟@x�6��"�!���>x���[@�{Q�y�`C�W�!�4�"�UgE�[GV!QP�O�!�=K�����ӑ�
��p��~�!�d]=2@[�#� #��=k@�GB�!�$� |�>��/������&  s!��%
Ĺ��͂�p�z�J��C�!�C,dM���TKA23ؔ5�bCE�!�$+�����X��YDb��!�d�_�tc������%1!
e�!���~����ıB��壳���!�d�64z|jQA�bk$�YC�Ӌ9���B'Q�hP7O:2r*!r����y��܊1䶜��E[>zP�*�]�y2$�>@���wB�mO�ـ�$Ĭ�yrGX()\�Ճ��űX�D�³a��y��ӎF���yՀ*J��G�!�d��Xy��a[ ��[V�\	!�Ė�n�~!{B	�p�b�î$!�DE<L�P��ȝ!d�|D�1@.N�!�%k$�$Śx�t��;�!��W&k�^|;��P	R�ToV�g�!��˔] ��·K�X��Ō:�!��73��\����/�ީ��AU�`�!�$\)bd��0��T��#oYZK!�4 ��u*�&_�r��l�����U�!��B�7��2:� }@e��8vx!��C�ql�m*H�rc�Qc*C�w���߳Lx*=Ȑ��pF�C䉋w+6m8��D'vh̼jPd�5� C�)� �X��$�"n��4�b�1D����"OBy���N���z�aF0C32��"O4��&hҹ2�n8� ?w���5"OL�CW��n���k�H]�~e֍"O�I�&��� �v�ʜ>�\��"Ov��*��������`q S"Ox�0�7lA����1H��"O��Z��?jHa��nB�w20XK�"O20�c_�i��`Rl<>%ve�F"O@-PF�ԯ$�2�2�֤
#"�83"O8�� ��M�<�)D	M"-
�Ͳ"OR��u%A���80�G�-�ވ�"O��2eD�r�>T����-Aߌtx"OpU�n�4;E̬ڀ�X�!�܍��"O&� f1:�b�2%L	-�|�C�"Ol���,�2�*Q�����d��"O���������Re�ċq��M�s"O*�0�LY�X�(@e�`u�I�"O`�cׅ܍�}�s��q�=��"O�����V��>���B�l,D��"O��獊+{P�Ӧ�>i��*B"O(���4`�������n�Y�"OH�Sd�yL	����:���"OVb�H֪r��43���}߼x#"Oy�bM�@�p�"Z�X�v	�"O��Z� ��}J������.���2"O6T9a'��|.�jA/V'Eb�=�2"On����&sn�rX��&�*8!��i� I`6���0¦�B�%W!�$M%h1Jq�@>��`dU3Z7!�ā�d�{� '��5����P!�ҍ:�rPK#n�@"diAR�2�!��,�fQ`r��z�����ӏ]�!�$��i>0!3��������b�<]�!�d�>>�P�q�g	�a�P�YToc�!�lm@䀃 ��.W�Ԋ'A̚S�!�d]+"�H*X�:6R�JB�pd!�DXH�t0!�c#څˠ ��Rg!��p��f�v}0t�5�E�,\!����D����.\�N�{���B�!�@T(N����w�Xġ�-�<x!��_�h�X����P�3	.)M!��V��-�w�
0$=dXa���W"!��Ұ=c�� W�Ǻ%�J���",!��B&n�F]w��+�p!܃j!��ܢ:`Zq�C)�<P:�S��ԞY�!�0�nq	����HO���S R#�!�ē�R�4����Fi(�zV��2'�!�[�<e�h2�N�EOj3��!��<+ v�{8���
��Ql!�
a�ص�B"�T��5���ɞ&W!�2}:`�IqL�({���P�J�q7!�ޝ*#`L�whM,A�P��Ş}�!򤏒b����AS�d���r�!���&���R"��M)��X6B!�&+z�Z%$Cb������/!�$F/&|�}��yD�q�֥�j3!򤛞Bp��+E�z�]�^d)!�d�9ij�
Ad2l�
vI�X!�ě�TV�ݹQ��,�$\+�!�i!���I�64s��W�w�n�JC� )!�d��8E@0��~x�ٲ�+D�(�!��(-B|@�!��%��8s*V�A�!�߷[��@��p�8��L�!�� ĳ�EG� Z�����Pz��"OMr���0�,�r瀗EJ�<"Ob��RB��q�$�Y�/LP2DH"O����O��p #�oϏc��{ "O&0���ܟm]��ڶ��V�Xqʁ"O�Ӧ��~�F� �'^�v�G"O�Ԡ1-P�������q�>��"O��+e���maZ�Q呰J�Ti��"O-¡��i�}�vF��5�<��V"On�@aU�9���ӄY n��v"O�R�(�Sx� ��i�S�>Ԙ1"O��wOt���P�iqv(($"O2�j2)Y%H2q�);v� "	�'GT\�ԭ�&�Yt� /4��3�'����a'G<t�q�c���0&�Y�'��r���'��"	2Y�X��'��5��I�5�땟�(���'{r�jӆ�,b�j�) �N�|�F�
�'c2�;�/]��&ɀ�![��:��	�'��ZC	!K?�����61$U1	�'����C�7����N��~�\�	�'v�(���D8�kw	\o�H��'� H��g�^X��+ס�i�"Ȑ�'-B%	S�j62R�e̷w�~!r�'p&���M�?n��DY%%�~�
�'~|2��$E(�d���4��9�
�'����L�HV��C�D�'�����'�~���M�������('�Ɛ��'H�]�D�hrT��5*���'4�A��@rꀕ�Ԅ��>�Ԙ1
�'l6<Ұ�
v�Y{�;Z|��	�'�&;p�V��T*��.��s	�'
-���1=F�J�NG�~4MQ�'��L�#n�Y����k�^@(�'���"�C.J�Y���b����'�^T#ҩ�����놁�b�aq�'J�`�W��W9f����T5B�
�'rYE ^���G_�LE���'���C	K8_���)���Ah���'�������[�td��儙8��I�'$p��)�i�N�P!��Q`���'��3��T�V��mZeƝ0rx�h�'�*�i��̮""rŹ�ꙟ ���'�V<��W+�����b	r�'�̛b��]v>�(��S��PMh�'d, qnٺP*�'��&�6q��'8Ԉ����O
���v�X�d����'S��W�W*u�X�z����.u��'|��K���1k�H-z^nl��'{Q�ơ%!6�ȹ�쌮n��y��',J�1v����AQ�X�P�'Q����$5V��S��񈉹�'�hh�CLB1z}���S���+�'9f$b�4G$���Hx,s
�'Ø�[s��r`�����*��1��'�L��N�z^��A0,�Ԝ,��'�<z�.Q?ꉢw-M�!����'9�K�LW;c�%��A
���0�'�h)9�X/)�>	³Ëa"h��'�\�'�T"C;�D�2	�U	��	�'��H��[/ Ѱ񚵈�:R����'���2�̰:B����	¯A��y"����&�24F#���&�y2ǎ=;2Aq�6z|9���y
� �}�����Q���̵s�%a�"OV�k�F	�B�ZP!�Tx0"O���/���2	R�e4"3���"O�xy�Hޘ�d�F��`$�r&"O��
��a�W$
(�(` "OrY���Ln��)�@�[�:��m{�"Ot���J&���#���R����"O���w*�6��,����, 
��"OL��a��� ���[�
�-��"O�AaR�D@�ࠧI�[ҭZ�"O�A$%,z�՛�e��I�"O$]��o
v��3����6���T"O�(�PdՈ�4��e��o�8i�"O�k�S"	�
	5�H�"��Mx`"O�A��ɂ��e� \+][n��"O��N�0^�����nBVa��"Op��ᤏ�<T�F& �I/��2�"OPpQ櫃�O X�6�
/)b��"Ob�"� G�x�t��&��j��p�"OޔA����eV�򲥖�N(�"O,��v��;�P05� <�N��"Oh q�kO
L��T�W=o�T�"O�4q���9N�[���B"Of8��g�����âҨs��=B�"O�}PcMȾ2aP��٨Z
���"O`؂'"�5m9��� ��� ]X�"O^<���*��!��/R:<�ic"O��)D�1RT��ƠR�0r"OHD�   ��   �  ?  �  �  �)  5  L@  UK  jV  b  dm  �x  ��  ��  ̏  ��  �  ?�  ��  ϯ  �  ��  !�  ��  ��  �  �  ��  ]�  ��  ��  9�  � �	  W �! ( e/ b8 �> <E |K �Q /R  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+!��6*\�c�<4�d5h��'�B�'���'	�'/�'�B�'���U�W9��m��Ʊz�0�b��'���'�2�'��'�b�'�r�'���k��.Kªa��͎ 5���Ha�' ��'���'�R�'���'���'����
F	�>]�&ΏfEP$�b�'�b�'��'�B�'�B�'O��'�$��zm@|XpjC�6�D�'��'���'v��'�'��'�"1�)ֽⲵpa����j5�'���'���'t"�'��'��'�%؇�Δ*��� A�B4%
0��'�R�'��'o"�'�"�'/"�'�f}�b���Xs���]��X��'iR�'���'���'��'W"�'g�=��'��"��	�Jw���'���'j"���d�'5r�'}��'��u�1� (iL�\r6e �t|:\���'�'H��'J��'ZR�'vr�':h(uC�=��)��G-P�����'��'u��'}��'���'u�'�;+�'HhufUmzn��`�'���'|��'���'��'p��'�J���R�h�����*|h�p�'���'��'���'h2�h�x��O��"�q�R��t�T�)����G$�|y�'��)�3?E�i)�ZT��}G��E�ɢf��<G�)�'�63�i>�IΟP��fL��,2�j�>LX]�� ՟�����Z�]E���Tn����O6�,�3�=��)DK�I�T�J�yR�'��D�Ob^�'(P�,Þx���BxHl8c}Ӥa��d,���M�;(��j�L�'���	�"� w�8�����?њ'.�)�S'���o�<�C];�NŊ4��6L��g�G�<��'�*����hO�i�O,���=pUl���*П��ik 0O����F��f��֘'p�Y��n	�G�PSuj�p�̒��\}��'Q";O���\�s�(�����ڢG�_c&�'��\��H�����VßL�v�'8�	��b�8�tKS�ćc$��K�S��'%��9O��"��8Q�D|
��N�5�`Ab@5O��n�/Dz���V�4������ňY��L��j�0�1 4O����On��;�6�=?ٝOx���?_$��)S�Y�;� �E�]/_�z��M>�-O�I�O����O^�$�OАqU���R����G 9?E����<a5�i���!B�'x�'��Oy��Ql>^p�1(�%O�!��H�AZ��?y����Ş(�@C�.YX�!#�gʼ�p�MK�_��8S�{��d6���<tg�?^:u�"I@  � ��TI���?A���?����?�'��d���\��
�O�|��F̵`�f��p�B�!�\�u;OYo�N�7��Iݟ��	ԟl���w��m�t*�8~��1���
&�Umx~�DX?c�p�nܧR�B�=������_���S���<���?���?a���?9��4�
5?�I��H�����cR�'��`Ө]��3�����]'���W��s/�$iA�v_��Pm@N�	����i>�I��զm�u��+�,4�!O�;�y
l�/<��@�'��<%���'N��'���'��9�@�|�.�k�n�9��	�D�'8R[����4z2����?���I�caPA/�8@qI1��}��I�����O4��1��?9���x�P�i�7��Y�Ѭ�,���s'&��]*?ͧv�������Hxt��B��p,�qٳG�����?���?��S�'��DϦ=�T
Qw���#:�U��^�3W4�KtU�Xߴ��'6�듛?I$&���	'�X�2r̹P���?����� ڴ���.z���'����iJ�pt+�/R����Ӊ�����IyR�'�'�'bS>Y��	-v��R��%[��S`	��Mc�Ǝ��?����?�J~�p{��w%� �6�Y?D�L���
�\��p�V�'��|���h�>D��<O���'/� �;���L� |�"6O�a��m;�~�|�X���Ʉ�	�`�rB�^�4�ԟh�	П@��Wy��o�@��b�O����O�(v�U]@�Hs&���R�!�!�I�����OB��%��p���a�W�qt��rUl�"*�ɯ��a2��5Nvb>�ir�'Dv��I<~�Q���m�Œ��N_��H�i�mޟ���͟�F�T�'U��1�\4F��8�N�Bo�]Ғ�'XD7��>:��˓ZZ��4�$�/U�t�0�0��ֲ(x��r5OR��O~�$��tP6�=?�t���i	?(��I��E�Du��%M+�D�J>�*O���O���O��d�O���f��W@�f�֔a�������<�G�i��l���'���'��O��nD�.]ԺC�&�rȰu���Dꓸ?i����S�'PTz�)��0)��q��_}�00�-�@�M�'�0a��[� �6�|�X�H�߱wb�9�EB� l���Yğ��	ן��I���`y�h��M��,�O��2GcK��>�Ƀ�ޕv\>�p$��M���i�O���'���'[�Y�kۈ����[8�`�F� #�|׿i��I#�<�c��Ojq���� �58��1pt�!��ӌ"�(K�0Oz�D�O���O��$�O��?mK�������Q� �4@I'�������(�4D�Ҕ�'�?i2�i7�'gV\�S�Q��<�#��Bx��|Z�M��|�Ah]&�MS�O̬ȁ�5hrN�hEbO�@z6�i�/ЂB'`U��'z�'��i>��I���I
jf�Q��Ǉ'���"�@]
t�v��Iԟ�'{X7-�����D�Od��|���)> &��7�U���St"�u~�A�>Q���?�K>�O'�z�!\�BL�E�(f��Ѐf����P�i��i>�*�O��O���f�0lT����-�^��#��Oj���OP�$�O1��˓B��&�W0+b��"`�eА
����'/vӢ�D��O����Aݚ��7�L.Yπ�[0��'h����O0��7M6?��W���� ��˓KJ��sb�:-kLLs�(S	N�,\͓����OZ�D�O����O<�$�|J���I9(:��t��t �Аm|���VB���'H����'��6=���$N&-��!Ā^1 ����OT��1��0\7-~�$r�bLRp���ǄE�!6R��mn�` c��|H��?�d�<����?��n�����$	B��yP���?y��?������1����矤��ϟ�SE!F��郁�E<�CKS��7y�	�����X�	7`(8]��eƾ]��)&+� ,n�|��K���TX4��|Ⱜ�O ����"JJ}gn���މ�	ԘW%b��?��?1���h�������p���{j��� $���D�ڦYp�kMRy�gӶ��1[F{�Β�DP��!���|���џ8��ޟ�P���q�'x��#�%�?1i�_'l��@F�++x������'}�i>��I̟��I���ɔBѮ]��xH��ǜJ)>�'h7�$>����O���(���OJ�[�C\0>pM:�(ç3�;�X{}��'��O1�4$:�)G�x=�I"M�J�Hš��Ar
�ZԈ�<!���@���Q�������P��U�71��QAAH�9V^�$�O6�D�O��4���h7��J݃+l2�\"��f�F-Y�0����yb��a�O�5�'v��'!���W�bX��
�Q�Dh���9H�b��ֺi��I;{� i���O�'?1�];ɲu���ފv��U�DD��v���	�D�	џ��	ܟ���N�'X�D�Q�ON�qڡ�2,Ǭ����?Q�����W#����'��6-!�dY�?d��rE��`L1Ӆ�;��O����O��9Iz7�??Q�&
+F�xæÙ�z���#gi�>	�Q�r����'�d���$�'��'u�a��1@�=i�kWqh�Y��'��U�� ܴ9F����?����򉗠�n\���"+��*���.6�������Ox�d&��?5R����q��q鐥�J�`�1u��#UkD9�i�S���|:bn�O��I>��� (eˑ�^����+5#H8�?)���?1��?�|�(O$`m�Sν)��Y"�&�H�^j�Gsl��'i�6� �I"���O��'hCMmL)j��]�.�>,i�h�O&���z˸7M7?�ІV�T�\�>�b�͹Be��R��v9���e���'r�'���'���'D�ylЀ��I�be!��=�@��4l�2����?�����<y���yWΉ'y@�^�D�����*�E��'tɧ�Oʎ�鷹i �F�(���N��	���P�BԊU��Ā(1���� ,F�O��|��K��r����OҼ1Jý^t�b���?i���?I-O��oZ�:����럜�ɗt�^�
ΔI�N�3�- c�6u�?�w\����|�*���V�����-r�Oخ����' R[4��:w$P�	���������	Q�'<�B��?C��zT(�'��+��'�2�'���'�>��	�B\�����E�cT�Zgc��O��Q�ɍ�M˶�� �?9�<��V�4�
yԩ��[M��Ke��|pB�2O:���O����nKb7�1?AƠO7�����z�@�0磓dRT�¡Hۤo�<�'�Ė'�R�']��'���'C�x��!�3�rA��!ͭ`���#EQ����4
�K,O(�d>�S*ZH��{vdR�b�̄�TXE�H%��O2�$�O��O1�le�P+�{CB(���[|�^l�"��JsH7M*?q��%�,�	H�IRyRnمk���{�۠Xe*E���X �b�'�2�'A�O��I��Mː�K �?�9_n��q����O:�y"�k�⟈��O��d�O���0L���Ə�%�I`$�4�Rh������|Ҵ|[L�?&?e��PԺ	��)=-�,��a��.1������ ����I���Io�'Xa�9ic�	�U!L��h��*@���?1�� ϛ� Z�����'K@6�)���Tb�)2.�5:�XjՎ�3^Bz�O����O��Рv��6m%?��y�Q4��7v@���D��6?2(�qfÙ�?1$#��<���?����?y�%Ӻ�(��	�Ij�<@WB��?����DWئqĥ�vy��'��S���|��#�<D TQ���� �F�	�����$�IW�)��+���z5�źB�:��*[{�`� �K�L�k.O�)�?a��0��2+)���ˮ��1�倎���d�O����OL��)�<1Ÿi�r�3���,O5��R"�zc,գ�gǭs��I2�MC��"�>���XV��nZ2n2�a񲬇�]Z����?��Ś�M��O���ٌ��I?� Τ[�#�6_�L	"��[B)�YR>O���?i��?Y���?����i�S��0@�l�JK"���!��Bmp���ş4���s���������_?0�`�FV9J4$(5�3�?����S�'~�&]�ܴ�y�/�	��=Sr�pČm�b�y�L�>%:q�IQ,�'�i>�I�Sްaa�N')~��$˒��N9��ԟ(��ΟȔ'�6M]��p��O��dҀPLl��#m���(�:AN�=3�*�ȹ�O��d�O8�OX�v�W~\L��/D�?t������@�_�� :Ta%��>��aE� ���K	���^�iw�%H�L�ޟ�I�d��ΟPE���'l\�%.�7i�A�wA�o��u�'��6�י\�&�F���4�p4�Q�Q�x�𮔌*լXX9O���<AG� 0�M#�OH�S���Q�P�N��e�t.�����:�F��,՞�O���?����?i��?��n�&X5jC  "�@�����Ad��S,O$�mZ7>lf��⟬��Q��=���X 1����˦"l,ڤQ���W�S�'/�x� 7��
V4�d8�"-���aᖙn�d� /O�����?���5�$�<�d-T�� [�a�o�����?q���?q���?ͧ���U����Z�g��5��)���L =%�s"�ៈR�4��'B���?I���?�PD�Uf�SW*|���E�l����4��d�#�t��'��OU��VB �y�H�7q��k��J�y�'���'�R�'9b�)	~[�����@�'��c�2$��D�O�F��m���DRyrw�t�O��oH:OH��أ��_^Q5k0���O��4����{���Eu����.W
}�j}P�S�6���k�%?�t��J��^y�O_��'IBBŭ~B�����h)���T�B9R�'�I��M�����?1���?q,�f����Q�8�j<�儮	L8���Ts�O�d&�)��L	]�e��V<Atr���Ꮵ;�� !uA�4Z�d�S.O�iU��?�n0�$U|�F��U���V��X� �F�5, ��O*���O����<��i@|� �&�7O-D(�T�X�1��ckm��'�J7- �I����O��s��Lls�ȐEH(�(�r�@�<��Մ�MS�O�q7'	������<	�M��2�VyIp����#)�<1+O�d�O��D�Ot�d�O��'=�.p��(�Y+�m���8e�h)B��'�}����?1�����<QA��y7�۝f�C�'�'���@��3
�b�'~ɧ�O�P���i��3a����(6�d�H�_���9�d�'I�'�	ҟD�I5lz�%C'2�&���Hz���ϟ��IԟD�'l�6��c�����O����5P��7&�jQ�%e� jn⟌�O��Oz�O�i�a�4P+��`�N/�xi����r��X�ld�r3�SX��S��p��O_7<�|� 	%����ٟ������	ğ�E��w����\8R:���#�*j�ȀS�'8D7M�?x�d�O�o�L�Ӽ����>���B$L�B�U�����<����?i�:�dm�ܴ����~�:p*�O7�8+�DԹ��DR ���ǖM��Gy�Or�'K��'cM�^�TܷB�P����I���M�W�4�?���?aJ~
��G=:��Dæ\���e�-n�L�{�S�d��Οx'�b>���d&3��pK�m��ݠda�Llu3��IByR��k�~�,8J>A+O 	Ӷ�,z�.��A�8h�Tl����O
�D�O~���O�	�<iw�i��t�W�'o�����J(R�BE �IG:PLX)��'0�6M3�	4����OX���O6t��"�X_T�XC$T������}s��4����~�p��O��O�bM6T2���
^]B�1T�ަ�yR�'�B�']�'MR�I	(pX��1*U#:%HѠ@MT�E�����OD��ܦICM>��I�M�O>��`�">L�
v�B	$I���e�9���?���|ꢄ�,�M��O61�5�ך�b��i�;	B��i���(J�b���'��'��i>5�Iџ����d�iW�3n(��3�Q������֟��'7�6��а���O��Ĭ|�3AW�8�b��㝸L�Չ�%AW~2,�>����?�K>�Og�<�p�Ϲtᆵs�iڕ-��4;bfN�6 ���i��i>m�0�O6�Ox�6 �b٠���Ⱥ9><�0��O@���Op���O1���7��6�˲�RB!���f�:4;��N�'N@��'cr�cӰ�\�O���9�pQC 8��	�3Y�'����OB��jp��F�Py`.�S�mp�T��P0	l�e�)�;X���Ey��'�b�'X"�'��[>9w�ޞ}��$�	�WX����ل�M�#�?���?A��t�j��.D��U�������@4k���O��O1�~ȣ�z��I�6?�QP��N�'�P�bK�y�B�Ie���rB�O��O|��|���g�dI�/�`������0QD\
���?q���?y)O.�n��$���˟4��e��2S��S^]��G�>����?i�W�`�	ڟ|&�B��?�{�!N���l9?a��E�9`~U�i�v̧>av�$�6�?Q��n4�iѧ�T�v�b=�scߧ�?9���?���?���9�5 q�R��\`���	}�H���O�EmZ1�4��':6�8�iޕ���%�d��j�[f&�y������p�ɆO��o�u~�)Y���� ~�V�Y�l+h�
��J�W�N����7��<�'�?��?���?q�!^@�(i��݆>������XͦM9��؟l���x&?i�I��`,�wɎ�l��z��X�-<��Ol���O�O1�@Ղ��ϔZ���(#�ސ:��mZ�	�)�b6M8?�����`:���\��qy�,ӽb��[��]a0���)���'���'i�O.�I��M�DJۊ�?iPK�+��Icȝ�9 �(B�c��?�U�ia�O���'���'����,"PD�#m��l�`ɓ0b�����in��$O���P�O[�h&?��ݞ,6$�ɂ5VDL���92��	��IП �Iڟ��	Z�'JՊ���G\�k���	�I�0٘����?���{+��e ����M�O>AB��-B�,x�	�
d�!B�:���?���|�s���Mk�O�(u�K7]�TE�7O];'Ĩp��`7nۖp����֓O���|z��?���k��z$�C�~QX�rp��&��8���?�-O<��	 �l�D�O�$�|�����k_�e#f��TjLq~��>����?iH>�O�d`ĩ_�y���U UP�: �4�AFH�= �(\���4���S����O0���HK�q(jxHc��_������O��D�Oh�D�O1�P�e�FdD(+C���ӂDF��P$��5L���',"``�`⟈�O���.L�r��p�ܹ%�x8	V�ҌyQ�$�O
p�m���wdYg)�S#hZ4�+�����مL>a��xyr�'�2�'�b�'>b[>Q��T`U,�X@��:D1�WΘ��M��/ť��$�O8�?�����uG_�j.Z�Ar��������?����ŞS��={ߴ�y"�W�y�ū �C:]]��Q����y��Ъ
C<��	��'F����ɽ"�>��g��� ��N
4�����	ޟ��'�p7M�y�����O����NAL���>�\|��a3
"J�lh�OL��<�I�k�~�)d��(C�Ԥ�A��`C*�Q�4�a����g���N~��O���sV��ϋ�5��M�Ҧ�vz�ai��?���?9��h�������@�$�b��b'���nm�Ŧ�قK�ByRFn�L�权 ��B�,C8��h�G�~Ԟ�Iܟ���ʟ���֦e�u'B����
�Q"����i��l����-�E&�`�'���'�'W��'���ծ��sW*�0����zEn�s�Z��޴_ ��*O��$*�i�O<��Kt�������zv�X}�'@��|���DE(@.��G�B��,��G[4h��c	5�MS�Z�8ڢE��O��<�d�<�E��IL L�s`�<q�ꀄ��?9���?����?ͧ��D�֦�Q��ܟPȰ��/.�d�2�܈A�,��e�L��4��'����?Y��?&��l9&�*2�On��A����6�y�4����z�����̸O�����\z���-�*Z"�]Á���y��'���'�2�'Or���iVJ�jE�4�ȴ��$�	�����O2��Gʦ��u>�����M�I>I&�V}��,�P)%!��xdB�����?��|�!H\�M+�O���Ԥͅ4�ݹ�Oގ�����]�XP�'��'b�i>��I՟L�I9T3��
Aɛ�	q������d��hyR~ӠECsM�OD���O˧,v�a�hN�OU��9��E��<�'���?����S��F~rq��쓜&J�ږ��;<�`<�w' h��ƕ��t�d"�D	4@����+�88��:1C,h6�$�O���O ��<�@�ilU�U,7n�N���)�@%Cbᙳ]�"�'�875�ɑ����O�H����3��;�B�=3��L�#�O�d�`�6m0?14	� ��>�"��32���W�k��l��x�P�'���'��'���'��Do�]C����P%{��,2�bQa޴uq$Ĉ/Ov��!�	�O��mz�!K��zQ����� >p�9�ʟ���}�)��ry:�l�<IAi��n>jU ��R:���r�K�<��cS���IU��Cy�O2�Z�cv@�I(^���E��O���'�r�'4�ɏ�M#T/�?���?��W8H�49�1@�+Hj�:bh����'���?������G�^���lZ+4{�T�'���EA^3�F`)�)�6�~"�'������Y�a�$��<P� ����'�R�'
��'��>��� �%���$	�|i�Lϻ����	�MS ���dX��m�?ͻ��ͻ���L'�1I�Y�y
0�͓�?����?�q^��M�O�|���܂��7���DJhyad��>A6mVő�`���O<��|R���?���?��x0�u�-z��mJNV[
�١(OL5oZ#����Iğ��	�ğ�둪�\G�9�d Q0z�\y���J ����O��b>rc��b��ѱ��̢,�P�qB/E�n�*FHOyR�GI�]�I iu�'���,X���f&^ɚl�bFe����Iٟ�I՟X�i>��'46�qzn����JQ*n	�Gj�%C-Hq���I��?qEY�T�	ny�
�
��SfY(�p�@��#��|�@�ik�	6�lli��Ok��$?M�]�CN����A�%rb��ìSFWV�I�t�IΟ��	����	\�'�v:F�N���f�#cx(��?���%��,��I�MsH>��NǿC�$�(��ߌ'c��[b(���䓇?Y��|�qo �M�O(���� .�e���0$�)��M� ˓��~2�|�Y��S�x����0�6\�	1�d�׫��b����oR�����py��c�Z����O��D�O^�'VK�L��#ɗ%�1 ��O�y�'����?a����S�ꀄ��kצ�% �hg�X� ���Q��؂T��Ӟwk2cK@�	&+�43�ʿ9Άв���!�<��䟈�I��P�)�ky�LbӔ8Zh�(q��r�Ε8K|d3�@C���˓LV�V�$�U}��'�ҡ�� Bk���үE�0�t�g�'>��K0������!�Пp��t�~��cW	D� ��8R.�<9���<I,OJ�$�O(���O��d�O�˧h�aT�_@o:=�b�Y� ����i�lݢ"�']��'��y.r���2|���YS�F
}�pФm��0�����Of�O1�Ĕ(W(w�N�	�7H��2�M3�,�@�n<n�n牛!S� 9��'�v�'�$�����'TṈ'�۝W����t [\J5���'�B�'2T�P��4��a���?����h�����^=�VZ%S��0�bD�>i���?�N>�4�ü+$`A�C
Ib(�УIt~��� <�u�4����O�a�I`�⥙�%o����y��K�]�h���?!��?����h���D�P��p�ɹT[=����g�.�d���VM��|����Mӏ�w�84�aRGD��InEdhb�'�r�'�Rm?7����֝nQ`t��?�d$(Vg�2�=��#��Qr8��a�|�S�\��ϟt��ݟD�	�����BũBh������lD��h�Py"��hQQ0j�O��d�O擟������m��G��	X);G���"�:�'Z��'�ɧ�O4��K�J��~¸�A�%�k��!���ϛ�N�<�eE !'���p��Sy�H�D���2-�b5@1������'���'��O��I�M�`���?���� S���D%��-��O��<Q¾i|�OT��'�R�'���A(%��gE�Hc��45C�ɳ0�i���<p��|h@�ONq����1p@�C��gy��Y~a�$�O<�$�O����O��.�0{9Ƹ9�@ �^�.�Q�~�Ꟗ�?a��?Q�i6��\���ݴ��^�����!��h]�4h%]20�d��M>i��?ͧW"m��4���פa~F\9sŊ�c�&����%V�}(����?iM"���<ͧ�?y��?�BL�>���F~�Y�0ϐ�?��������[��ş���ϟx�Oں@9�@",��Y�Bَ)��1�O� �'���'�ɧ��R���a���:l>�X�iO5#.E	R�8O�*�sї��S�q�B��G��p5��pd&�r��3'��R���ܟ�I����)��gy��tӘ��#�l8Lp���!"����U��e>&� ����a}��'Rd�&ʚ$ c�톭t�<'�'v�G_3�����Ё���	��ě~B�e����]|`��p���<�)Ot�$�O2���O����O
�'x���e�=�H�x�+�Lxj�Ÿi��M���'�R�'���y�'o�󮋓vU`l�,t��fjȰrW�u�	���$�b>e�g�@�9ϓ|�| �/I'J�<��Xy	���o��t��H�O�ŘO>�,O��O�L#��6�xxi\	|��l Ӏ�O���O��$�<�0�i0p��]�\��pz���;��d�>Kq��?�pY���	|��f*����Cv=��,�� �'�4z��E�Y8�P��t�ڟ ���'��9�N�,HEԄ�RO��&*�7�?���?1���?���I�O~�u��Fe�:î�!db\3uM�O��mZ�\���	̟|�4���ygO" �-ڥ�E�AŰ���ә�y�'
r�'M�(��iU�i��Я�?9 2��=�T�
�ņm�(�.H�h��'k���	ߟ�����	Dj��E��,(ĉ/tVE�'"�6��/p�p�d�O��d/�9OН���'W����"� W�by%
�I}B�'�2�|����W ���+E!G��0Ɂ)�<BNHl��	�剦$�e1��'B\�&�h�'��Qp�cϳ"�H`�j�4#\�S�'U��'�B���Q�h��4"�,���>��t��k�,4�be����� ��������o}��'L�wL�A(2N��-Kƅ�X�!��qd�"�������M�j�i �I��|4검�;\vĐp0-���
�9O�����sK* �1�P&̈́�x�E	8.T��?�P�iʶ��˟�`nD�I�����	1*P�PD#�4IV�L'����ԟ�\k�$mZN~ZwK�Xk�oÊx[б�gABm��
����]I�pyB��T5Ȍ�Oȉ[n� �\�h(��j�4H�� +Ot���|ZF�_�(E���T��0�jP1R ^^~��>1���?�J>�O �U*��"nqT C��Q��r# ڳ2/ޡS@��8,�i>�h��'�%�$Se�6�T��%h�����@�`-�lrߴ/��q�e�X�<e���S)�Lx�^���Ă�M�?��X�<�I����ɔk��B􎸑�̋�[ �%��ٟ���j�Ǧ=�'g2�[#�|2.O��ӣ�Yr�`���~�ڨ��=O���=a��#K|S@'ՙ�i}֩��t��A�<�����O��7=��#Xl���"6�&�x�j%��OB��?��i݆t��7md�� �%o�x/�m[a����taKE3O ��b���~2�|\�ȗ'��pP�M�A<�7M�V7.��Ók+��ꑳ~�����p��-�@<97c�(p�*�c��H��������Ih�I��k���*��%B dY.n�j� Ur�����#�M#%�����P?Y��PT�9E�W�p�6��D�נM�8��^" řsLQK������}�����f�#��	��M��w=@-b���/Bj��	�!�7*��i��'M��'���0|I�֓�`�
�l��iغ"�����'/t���g$O��Oʓ��O Io��%�Q�B/�?"C�����޴<�B��(O���=���~ͺg�	}�$d+��c0�K�O��$�O��O1��$9�OBH�N8�Gd���d��Jt�6��[y��4��D�����D��
��� ��_�bԻƫ������O����Oz�4���>��I�2�OW.a���G�lH�,Lv"��b�~�h��O��$�O@���4Muƥq�c��z���0ՠ�@�LE��r�V�S,������J~��nL���D�3�Q��@ҥvV�ϓ�?����?���?����O�z4�vh�RGjU�%ӈE]xX��'���'�7-�U��˓S����|��C &�p���$da�Q�&Zc�'�����b{����֝�C�`�Y`��0�\��F�N�KuM�۟��|]����ӟ��	�� �Ɨ/�Pa��ɆW�4��&(֟���pyrr�@�`uC�O��d�OZ�'�r �o�p�VS�僣sQ���'&듣?����S�$��f�����P��(1�D'9 l�j�b��x�P���T���0�B
A�I&��7�Q� �����&������`���\�)�gy2n�0��@Jh8����`�bf��"����O��o�B�����ǟzGF�)
� �bO���a��J����I�n �l�P~ZwP�X0��O��̔'[Vi��+ՄdN5"QO��2��b�'��	��8��џ��Iޟ��Is��ႌ?{Bt1��A�v�z ���`[L�6mR������O��D#���OXlz�e�MY�o��X:�H��xؙ�&UƟ��	e�)�S
X��0l�<a0��=@yB����VE<`Q��I�<�gϰr�N�������D�OX�
�q���s��2�(UXE%s���d�O����Od˓|/��lk��	ߟ��IZ)*
�)YF�ۈC���B�	ʟ��O��D�OT�O��h�n�lnP���m{"��*���%Z0���#w�ƥ$?eKW�O��dެLs�1�e�52$<�2�
�T���$�O���O��d:��K���1q�T������	Y�`�S)Ʉ�?�E�ia`��a�'t��i�`�O�9�(A�%�Ի'N\<�Pe1`�`h��6OL���O���C3ph�7m.?AG�"[x��)Me���u
E�l���9@�`�ڽ'�ԕ'��'�R�'y��'I 0�!9G��K2-�5�.�/��B����%b|y�'M�Oc����A�@u�#��)��8�bɊ4{���?����S�'_�����G�&+�������:|�̠B.���MS�Q����`��r��*��<�铰�P�� ����s���?���?����?ͧ�����Ec@��ܟ01K�{39 $��2fo̊c���I�M�H>i�H��Iܟ���ӟ��4H���q
�(��j��XHq���x�8�lz~B!EN�2�S�|��O�gf��!��d��'�6(�fX ����y��'_��'B�'���)��* �ݽn;� (��ԚP/���?���i��r�O��~�(�O���銋4��E��.�)#��+���O�4���:��J�.�eꥨ�b��ș�j�
|k��̟0U����n�Ijy��'�2�'��mQ���1s�Ez�1�N�,T���'���/�M[������O��'JuV�b�ʎ>涔�en��h֘�Γ�?iu^�D�	��'���J��7�ٱ/۠q�Uz�,�� �L#v�޴��i>A���Od�OjY�� �!=�l0ja�$:��A��O4���On���O1�.ʓs��&,����uAŦqf��� �ޅ��t`1^�4�ڴ��'m���?�"��x@t��5f�4^�⸉�^�?���5���ٴ��
!p���į۠<���$��.\U�'J��'��	՟d����\�I���IZ�d��.��c��1Q�@s��3$�t6�ڿZ�˓�?9����s��n >�����Ϳ�B@5eYY���OΒO1���{�"iӐ扣�<ŹT�I�~������	3��	�K��4���Ob�O���|B��FP���u�L@�Q�UEj�-P���?Y���?Q.O*�m�2'"x�'fB�h�h0휱z]:��ѯI�t>�'V�>Y���?�J>ia#�<g=�����7>l�����r~b��o%� ��i�ʒ�n�a�',Ҏ߯'5��G�Y&f�h�#�c�R�'���'���s�}�@�G11wn13�U�7Cʜ	�M�ԟh2�4Y������?qt�i��'f�w�p�V�F��r�"`U�$�<8��'U��' � D�fe�����݊$�8$���m2H8���tc@`�q,[���@۰�|B\���	̟��	����ԟ�`�K.���u�$�0ЕGxyb!Ә�� �<����'�?��+0�0t���c��[�R������Ij�)�(4�� ��[¤;TA|��z�Ҵ�zӺ��'�lЊ���g?!K>i+O�Q3NK-j���C�\.$���E�Oz�$�Op�d�O�<Q�iS����'(����P��ણ)5����"�'7�!�$�O��':��'+R��.@�$�w�Y�O�A�p>>Zʩ��i��I9p������O��}$?����.����B)u��ʂ�"�,�Iݟ4�I����I�t�	y��a HPgn�Wv���1Ȇ�/�e:���?�4Ǜ���.���'~�6�,����l̘��F��A����)E`�O����O���/)ݴ6-7?��A��	�c���2�)K?' X@+V$^�?9
*�D�<����?q��?�K>`�\z�c�n!����G���?1����Φ�X��xy�'���=��U�v� k� q�LP8{) �ǟ��O��d�O8�O���jt��ِ. ������B�Q7�|�F#_@S�m���4�l��'(�'����T P��0�Dě,~�Y�b�'���'!��Oc�ɬ�Mk��d���4��G�
���H��*�h��?���i�ɧ�4h�>���_1�|:��P5�xG�ǣl������?�����M��O�D�����Y��@�+�9E�����`��w���i�d���'�'h��'/��'*哶v�,��':�2����  06 J�4	�a���?q���䧆?���y���8����%�C� ���G�u���'^ɧ�O����i��$�>$�X<�u��xk\�`��?���ŃqW����S�O���?����t�2Z�|�G+��xD�d���?���?-O�l�
;�
����x�ɂ چ������/����)Է:���?�AW�4��ޟ�%�8z)�(8y>}qGʕp;<l٦m7?�↔G_F��4U��O������?aF��8+��Q�E�E<I�P��,�?	��?)��?ٌ���Oʽ�Ƙ �\���	*���R)�OȜl��1���I�pݴ���y�h	�/�kF�$[x���,M��y"�'���',$� �iN�	^�ndC�ҟT�cT��l@�a�?4�~�Y�l,�d�<��?����?1��?1G��<]���`�\h�`o�K�`�'S6M��{�����Ol�d!���O���Bg�P�q���f��8���UK}"�'�b�|������p0�d�Q�P[���}���D�iw�d�P�b��7�<�Q�5_J�:��%e5���s �f�Xi����[�F��&ȷ
B�e���0($�P���2y�,���W-J��	�@��o��|9���"#%zu���Z�,T�rc�K�A���B����?yS�?�&E�t�&��	��ͼ%�8y��Q�D�%��=>x԰#h�*BO( cS�T�[�r�C��;�>�B7+A��[���'
۠o�4~7��"ХY�o>Đ)e�оH���"�8|��T�!�	�X� ��f\<�D
�y-�8ãE�k�2�Cáʌu�p��BRӦ�(�NߤhgM�#F����&�_?�M�,O�*�D�O���91���X4de���6��.��K�� �I�'`��'�☟�8���]���'���$@R�L�v���i��	ҥ/b���>�d�O�D~Y @��(P�L�$E��D�ս+����ߴ�?q����ݪPH��'�?���TnW��b0q�J�
V���BL]K�'-��'�R` �'�'��)�qk`mse���vy�*e9�&������e������I�?�ۭOk�
N��L�ǧ�8�N��f%��B!���'��� �O��>�%�}Z�<�㣁8V�Ċ���O@�ه�j�8�D�O�����T�'W�I�7�`��㌌נSu�J�<�*�Yߴ_��P����I�O�E)�CK��s�jɾ.��������Iӟ(�ɾ5�`�O���?!�':L�1
�%�e�\:-��4��mN�������'�R�'a���2��(b��T}%�|ڄ�x�^��˟w�b��'��	��H$��X�,� 01�/�ؔ����9��R��4�<����?����(/_�j�c�P�1����tL��rI�>�(O���6�D�O���ƺ*8V)Q�c@5O&�����(y�4-��5���OJ��O�Y�D�A�OT���%P�)x�1B�L�P`�@�ݴ����O��O����O�s�P������4;�؂4(��`�^	Ⓣ�>Y���?����$ȴHk��'�?�`�W�k����Q(6A�p��or�f�'��'�r�'��8�����{����[�M�Ět�Yf��&�'C���@��B^���'���O:��(P`Є`&���0*4s�.ݛ �4�D�O��Μw4⟌��A&(:�M�K��q�_f�X�l�D~e~���'��'|�䮯>��~��@�勍�vC��ض]+A�}lZ՟��	0.���?Q����(0�d웳o���F����?��h��M���?y��6W���'���#���8�|0A��Hq঍mӈ8V#1�	n�'�?	�h�wj���ƃ�wn]A�NK�!	���'���'�,Y��J!�4��������)�-��!E�!a��A7k�`��%��V��'B�'K�)E7S\!���! � �G��{�H6-�O�Y��[�i>��z�W�ĕA'�ī ����	(ҎQ�H<������O���O@ʓV�,}�"��v�tM0&�� u"ܓ�I��_!�'�"�'��'��i�=�����r�Xe�%���T+o����<A��?����D�����ͧ|z��F�=:tX��>uz��'2��'�'3�i>M�	$ �T̀�E�g�l��f�:�J�C�O����O����<	0K	��O1��  5Ps�\�4\1�o�Y��v�i*�V���Ity�O��~jT���aQ�}�R!�=cR��!�Q�	���'��#ǎ&�	�Op���Z�j�"�!c�́�$%Z9KK\u�g�x�Y���I���'?�i�y�~�J	�!O�;3Sr�i*l��FD����i����?��'<9�ɋ/
����@3�lH�R�**��7ͥ<I���?�����ܴ��M�H� f�����v�n��(����şt���H��yʟ�M Q ���}����-}e�4��Vq}2�
�O>)#��Y�=�Yb��
�N~�q%���MK�������S��>!�C%]�ess
��{^TX�7�W�]�����D�'�DJ8��%b NR�3���{VC%ț�'�DCcV�@A��Z�d(�I���T:�eU*/Vݡ l����+��Q�'��'bW������ !����&�]v���8I�l�{I<1��?AO>9(O�U�QUkQJ��/eE�r�Ol���' �',�]�x�I�(�t�'S���0'��PH�ٳ�^8hG��m����Iy���?!/Ohʲ�i!�1�r��PpF�󏏲w%�J<	����O�+!
�|���_v�Z.K�bd���ơX3\�Y�i
�O��d�<1�^�	�!y�ty�� Z&t�ٴ�5Y��7��O���?�!�����O�����kLV%�^�
F����!J��'�Q��z�*�ӺS&���7#�d���J���Ћ�c}R�'���Y��'�b�'Z��O�i�%��A#4��s0m��C@�a�n�:���<�e�l���'DUt�cG%ŇtS��7ݽXA��o�<O�����4�?I��?�������C�<���õb���=�q�<�
7�O��O,�O�s�X��=::�!������e��$,t��ܴ�?I���?�R̮b������'���5���Ip$ĢB��ժrbE�z���'�'���<9��?y�����2�L�+/����R�r}����i�b-#K�O���O���?9�쇇a)�<K���&I��q�Ոׁ7�'��Y���I�����fy��1wv��Eo�#%�pX�N6�Qz��>i)O����<a��?��� jelϯO򜀕fˠ5x<9xWl��<�,O����O����<ы؃����q��Y3��S�
l8��_$i���^��	My��'jr�'����'�9�A�^'ZOb���"�Z@�U�R�c�����Od�d�Oh�?t�y(�V?��i��*�&�*P����W�9ä�A#�`��d�<���?i�'��a̓��Ɏ9<�`NxCK�TШ�Xdd{�0���Oj˓��0��Q?��I��|�S
��86���ZFl��aV�g��p�O>�D�O��T�L�Ĳ<����d�]�,�(5�6�Z#S=*Z¬��M�)O��9Ca	Ҧ���͟0���?�Z�O�V� �PX#��ǖW|~��UÓw���'"����y��'B�	kܧ,x<��'0]��Wӌc�ڜnZ�����4�?���?)�'G��	fyB���^�2�2�dӦ��|��úki 7��9���O|���OSr+��f"���Ʀ��K�Hz�`4G�6�O��D�OD�P�(_}�V���z?1���1.�Px;RCˠ`h�
�]ئ��IJy�GD�yʟ����O���ױFJ]p�d �.^%s�,� Pz�n�,��`�����<Q����Ok��P���"3OP RH����5��I%x���	���	柈�	ʟ��'�З)^30��F�&��q���M9%8 S��'[rU��I��h��o���'Ɋ� !�z�%��ZW"a��A8?Y���?	��?9,O��; 	V�|����,(��h��1E�2��B ��y�'a�X�|�	ޟ���,Qi@�I�YP�T�bɕ��O��E��4�?���?i��� &�^��OXZc,-Ё�ޘL$�!��/&}$i�4�?�+O2�d�O����)����O��	/��EJ���6E<P92i 7`G�7��O����<���]��S͟@���?�{]�_���A��Pb�I!`fQ�����O<�d�Ox��=O���<q�O���[AJCr���S)-{�P�r�4��V�b(��o�����	۟��S&����TU���W"�@��fG�1J\����iQ�'1R�'��ޟ�}�(�H����d͖^���葩����L���M����?�����V��'	����Չx�\h�1�$���g�r�j�AV>O�$�<I����'�\M���,)��b�I���\�3SEt��$�O>�d�:VgZ��')����I��Z��˘
>%�rk�6S�enZڟ|�'Y�=阧���O��d�O��ZC�٩��dR7`R�o�H�D
P�5�In��Q�O��?�+O��ƮX�㠜�b�r�k�d+W�����i"rI�yr�'y��'�2�'�剝*4�ɓ2��O��!
�*/O�"���E����'J��|��'Kb���6�'3�]�B��^��k��'v�I쟀���ܕ'��U���i>	�&f@�'֜�ƙ;A(�4��d%�$�Or�OL��O��7O�c��',N�!6�[,��P��C}"�'���'����ؐM|�ǝ~"��Ip'�c��X+#��*���'�';��'��hip�'f�ILʽ3�nF-in��5�=2Dmm����	by�
��&�������꽛Rg� d�p��Ue�$��U#�N�I�L�	���IV�	@zc/��OP0PXA�ʊQ�Q$��˦�'[�(K��z�8��O2�O���S�? Vp�0�T
`�5	u��"̄x �i�'����'`�'�q���
4+J #p��ф��#7�`M�v�i�<� hnӄ���O��������>14k�F�z}��,�!V+p(�rFR�nf�v� ��y��|��i�OT%�陛y���cF���x����Hئ��џ`�ɚc]iK<���?Y�'(H��8!Q8����#"�`�0�4��l�"��a��4�'��' Rp��V����c��V�x�#��w�8��ҩ}<�%�d����<$��آ}�� �A\����V�R������ ����O��d�OBʓQu����摰LȌ��=gf��$E��bm�O���:�d�O��d�5MjR9+&��
�� nb*4�f5���O���O�ʓy�����4��`��I��R�k�B�W�N��EV���	C�'��������#qͤx �L���朷P��݂�OP�$�O$�Ķ<1vl�<q8�O���Ʃ
�u��=`TF�$p =���gӺ�=�.O\��.}���[���������j�$^��M��?����?AS������O|���B"�0�z�0��ڐ{�z��qH�a�����'P~�C���TX8��J�Vl�B<'9�|�g�i�剦/���ٴq�����Ӑ���P, \����\��C�b��'G����D������yxvu�ÎҦI<P���M��.�?1���������O�V�qZPΘ�H�|�[����x� ��rQ��D �S�'�?YQn� 7�n�����:x�$�c�Ø���f�'<2�'�6}ZU�?�$�OJ������ED�P ���N	T�j#<�	.F��b�`���h�Ia�$mhq-�?�*��Q�7f��;�4�?�c��c3�'r�'�ɧ56"B�$���f��7�-"/Q3����~1O��d�O��D�<#BNs8H��e��uI.�"��.4�V���$�O�O
��O��0O�8,d�� d� j���0GΟ{�1O�d�O �d�<!!�M|�)��[<����K��UB� HkR
ps�'���|��'��l����H .�t��GD����jj)3��I�I����'č	v!2��i�������,�j<b�(J���En�p$� �I쟰!=��98B���'�Y�cg98�`7-�O���<�b��h"�Orr�O(Bܚ"�^�u�\t0�e��/��B3���O\�dC6��'\Ō�Sb[�0Ԁ�@P�+~8�'�2�V2���'M�'{�4[��ݔ�H�KW�&fk�I"�J��D:T7��O��)e��ExJ|�A�")=x%�v,�؇G��=ƪ��M����?����r��x2�'��҂��9g�| h�X+qa>�O6�DW��H��f�ȫ:t�'��4"�oZ��	y��F��' �W���h��\�� C@��J�0g�'5��'�B�p"<ت��yD�u		?$�:�o�ɟ�$b��ē�?A�����[��AkRh53oI�	X@8�y}	M��'r�'
�I��*��R\����5V���'�+>�ؖ'��'�b�|�'���H2t�a1�LD>��u��?e�6lь��$�O*���O��Z���f6��AX��J%��u�aC�,\�e�$\�����(%������G��>Aր�]���V�O8�V�z"lu}�'Z��'z�	�HUO|B�Q?zA5{�����4����BɛV�'��'�B�'�P�3�}�A�u����Ќ`�r	��&�MS��?�)Oԥ!� z���'F"�O�0��h^��i��P��,�>����?���^��4Γ�?�,O����n*r�q�ʕ@��q�0�ŀs�7m�<�5�3,�V�' ��'����>��:����AS�$�6P��NB+�F�oZҟd�	�B�B��,�'q��-�V$�F�\3���~h2ͰG�i� D��|�t���O��D🬑�'��ɸ"	�1���F�(��*�vtt��4&&͓�?�*O�?���1;�H]�`�	&����s�˛'�|)�4�?����?9"���Sf�	Uyb�'��d��
>�K���g*5���'L�f�'��	�i�)����?��
�!1GS� >@�˕��\ ��i%��\��p����O���?�14}�aJD@,3�MӲLʡt�q�'�f��'P��9zx�%�`�R��F�O�|�b#
�Lu���&�J�6�BXI�'eVaq&M� Rf��/&���$[f�ܤq1�@"`�dՈ���Wv~5�v ֒6;�p �'��_|f�v��3O;
����6R�9X��E>o��mS�"݄cV�`"��k�4R���-sC�f�_��,��&�(�(�a$�	9t]�[4��)Gj�)��H.���g�M6k�^YSB#X���\Pw�D#A6&�*W�E��Rhq�C�y3f*\�<�=+@�',B�'�b)i�V����1�d� 6y����R2'�Ťj�R��姐�w����'MY�'��Ax��,]����!ݺ@ʛ�I޵��-�$����٘��K�&у�l������O���-��`���^�fp�ɓ@���`�
�l��`� �,7�t�h��Z�WK�U!6M:�O�A%�$I�L�-W����@�19%��$�x�̀&k����D�Oʧmh�����?I�r̸$��,}�}�@�6cnmp'��]M�ʥ>uVĒB���%��Ot����8>�h�s��k/�G�:XU����a�/�e�Mǟ"~�)� �d
P�|,�U"V�E�*��+�%�'e����O>�S�K�U�n��v�̀8��d1šC�8�ZC�	�~e"���D�G�\h�U��yH#<a�)E�ݼ2+�Y��ƒ�CS� �?Q��X� ��U1�?Q���?����.�Ot�d�"@~\t�ʠ$� ̂A�Ό ����<؝����T����	|D컵쓄4��]�ҁ�����9R���W��B���W��I�G�,"9�oA�=�2��>�dm��ܟ<E{�T�t1a�P�*�� �F�	Z�`�$D��f#�׀C��,��!
V���HO�SvyRE� F�6�I�TRl �k�� ��z�N�����OX�D�O�e���O<��y>��i�=M�BJ�%*T���:GG��S���mV+�h%#6�Vux���FJ�0:���"���W*r@��,��tC�W�R��t6��Mx�h[��O����(ݴ�*0.�!��1�� �)�Z�=q����{ؘË��\�=iW�H�!��KԎp2#�B�}L���!����X}�\��{%�\���d�O<˧@�6�"�Hɶ9�B`j@!Q㎐��M��?���?�5$DtڄN�$��0���)եt:���!�m��ɑ�b�0Q�ؘB�C>�l�v��[�RU$>��pR����Ā�!�\q��#�h�0,����8�ꀀZ��dzt���W�)�D"�O���֦�%�>��Ai\�D	$�9U�'LObى�h 09PyAʗ8;�<��t7O��;!F�����	՟��OP�}E�'�'���Q7jK�rņ-k����p ��DC�B�T>#<���I�y����
�Ew���ᣘ	KM@������O��B`�ݧp �y�E��rt:�`_,���D;�)��Tj�OӉ_Ԕ���U�#N�1� ;D��T
T9�� �3n�6�p�d.o����'H�y��lݨ{f��q�����?�3BU�l&��`��?���?	a���4�4pp�	.)6�<�' ]�I#H�%�O���"�'! q���/	�<{�͇w�TH�'_��i�_�=bt��2��ցאp�h�@`����u��H8D��B�q+���;+��=@��5D����m��`�X��f��eӷ�HO>q	�����MkFţ\:|����; �9T��?���?9��?���8��?ɝOX�\���?�d��;]�v���t�Y��E��L0�|	���ÀGp�T��.�	��	��SY�|"����?�����h*���=+�6��̓~��ȓR(���C F�"���`��g/�ȓ<��=��AJ�%�\S5�(�:��7�O���M٦����<�O��u�4��b���5D�5 ��&�*J�"�'#rn�
K��T>��!葭&v0�Ň3��s'�=ʓTm)G��Ē�n?�I�����˶Ē�(O"�p��'3�>{����y�V=P�.�����./D���CL O#��
'�3z�[��?�OFE'� �c��!�� ���$�@�k�'|��ʔÕ��M����?	+����C�O���Ot9
��@>iP��S+�=� ��MU2w���$5�|Fx��e\r��'���SG�*^�&���)�矨�ǤŦ
C���lC�&�Ԝ�gψ�zHZ|�	i�S��?�ҤFL��8�!��x�n�z��N�<٥�/#|���MgZ��B B�'\�#=�O����"�7]q�Lk!G4>��C��'"hBL����'���'�2w�-�i�Y'PpΥ�U�:p��L��d���)�O�Y��֦i�h#)۰lL欣�O���'�����(!���A��:l:�'L	a����=� �tbY�T�ҥX2��ӣ�B�<4G5>�0��qkb����?���"|�4��'A��)��y p����k6,� �n�2�'.��'x���'^�4������'�r˧R���dH	{PIE�ݠ�p>�#��uyb��c����e��({��.jrȅ�I�X�h�d�O�]��S�d݆A�����=��y�#<���O���<�)z���9T���7���_E�Lh��@�<٦h�r�H[�L��[�F�#�<��W� �'5��K���@���O�'_�����U��Ƙzw�X*ed�12�W:�?����?�6�� �?��y*�^P[��N3Pl��ζS7J�)��	%#���j[�%�.$���!9z:L�Ҋ�W�'�0x���h�� �Ux��C<��KG�$	���	�"O�@Z�.�����h ��`qd�'<�O{����glV�Ԥփb�B�p�"O��1�N�QU<M�t)�#�tA�"O��p�&���={�;U��|p�"O�����C
���מV��$`0"O�hrb�&(��mQ$��i�D�`�"O$�bb� �6�dx��i$���"Od)�"M�-�P�I��5�P���"Oj�)�FH8W�v�l��^��!�"OT���Ha��dfZ�8lv���"O���+��lk�8(�"C	o^�,�V"O�l{�*F�3��/�!5B�tXT"Oz�r�(��f8�d�(P��!�"Of����\+@�L���$S�yPQJV"O��%G�X�<�b.��mU�'"O�9�,�#k-�� Kd��%"O^�[�)g1�� �MX(>BB��&"O��ҒHL0)���X��ڃ,�TXr�"O�,�d霞K�rP��&۷t�ژ�P"O� �/ó<����}��!�Q"O"���Ƨ6�������.���3Q"O��S��Y,����Ɲ:'��)�"O��x��6yΥ vK�?���X$"O$�t*�1Q�j;'wt�"O�k�؂=�T��#�J�C"Ol�	� ͥb)B�I�ҭ{���Xt"O��`�RO4@ѻu`\�2��"O�賡%Ѻ@���Y��P�Ы"Oة3p Ҭ}�>\`�g�(/e�!��"O�%#���:xI�8�R�Ѭu�ܥx2"O��vDJ�t몵P��R<"�~�[�"OD�À�XD��=�6�
J�����"O��:��[��Z����B�|��t"`"O��)�Ǟ��4ͨ�㉡1���Y3"O�L���V���BA������"O
L�6�%.�I��ʐJ�|hYU"O0p�g��Av��(�,Qـ ce"O��1�(ګ<�l@:�N*����&"Oh$��܎C�n��3-��<w:�A"OQç�3=�T	�0F����Qr"O��y��ׯ*gZ�q�,D??~fi�"O yb�	f�@���sSĽ�U"OX.@�G>�0r�cاjMP$h�T��(B����=Q���9��!��j�$*���c�Acx����@!�?���Y�}ڝy��4!j*`����\�<���_��8��gR:
����V
�n�'� ȲS�^��h�&ݨ�A�T'���m,1O
=�4"O@%��IOP��ʬui0i�v	T D6��t4�)�矌{�`�7u9�Q�R<3��0�h0D���wɸSS����
�>w � �VM������R����ۺ-#�p�υ}�l����H�4%�|R&[�'�´��^�(]X����0���Fm��j;�Q�ȓSGL���`�xܑ�U��$$@Dy�B�WO\������&m�c��R|��rh.�!�RJ�)�w��>}�M) �/(��a`%$� ~b�"~�ɾxX0�a��B�P����"&�C䉩_-��x�-�#v �,��d�A�˓l�ȡ3�'��-s��.4H;7��{��I9t�H:��݆�I>���*��u���l��D�j�DN@�fF}R�˚��>u�s��N�t%���DN���0a+��T���J�Q>9��'�W_�}r2�?�}�������Q�S�O�u�塀�-丰�'dĈi
HtäJP5^X�
9��)�矜�jW�G*��i�"p@��e'$}R
D60a{
� �up�f��+9��j�+%�z��0�O�}�`� %P{L	����Ά}�*6M5g����\��	��Z�P��|R&Yo�R)��͘�1+R��*�0P���a7N,=��F}2"D�m��>��qbV�[�+W�K$rm|���."�Y�2ܡ�bW�_�#|��!��6��j�@��& �V��C}�W�O�>�s��Ǭ=8�@���O�6��@83�n�#�PP�ӧ��r
��Fv�Y�n
�mm��j�����yf��~Mly�GD/�XY��!����<*2�8���x��liffT�D�a�D�3�Fq�d�3D�8��T?h>J�h-�#<�� [�C�I>?���sF���2�<�Ѥ\(_nB��?YX�Ӯ˾yO�y���Ȁ��B�	3t��Bi�"�H<CFJ��S�rB䉠"�p��Ҙ�2O�&ZB�I-��`i�Q(]�� e�*B�	O�HY!�eI��u��盵Y� B��(i��q(����
�P�C(Ŀ>|�C�T�vQ��%�*��4h�)��C��"W�d��[�&�c���q�$��"O��'�1:}d(qV
O+Ҏd"O�9k$J�|`��
�����"ON���0M�\����"�ZT�"Or��ɍR�����/~�La �"O����h�.+ظ��L�;>x�� �"OlxU�^�����! 5��!w"O�L�m�$����E�-,��9q�"O���*R���T"$&��G|�h�0"OtIP�C�J3Ly���U�ra�"O�Tc ����aC�1N��)�s"O��A�O�`@���3����"On]@p�
@
���F��aj�"O���E
8E*����n?%�B"O�hK�(r\
իH7Pe�a��"ONc#aL&	�@]D�Q/FMYr"OΤ��]r(E*�)Q�?J83'"O����dŎ8��x;���F�b�"O@0'�WIs����O	;���I�"O(�9���_/$�i`���c�"O�-�� �bK؄"���07TK%"O�0�bA^�<�h�<��ɥ"O4��#J�D�>E�Df��.a��X�"Ofu���O�A�:�Ҵ$�x_^x�s"O,��W�Pq�LH�䣙�`��U�"Obuh&K��J*����] ;{�p�"O�r!OQ�-t5Sgڗ\�x�4"OFY�@�]�t���˺u��zd"O�4�4L�IV�Z�/_<�����"O��I� ��R�*�;P�O�3���HS"O���� �3��X����{��\	@"O�P��J�L��9�Ta��1��h2��
��Mk&�kPd5�3����zAR)C"*T�d�e٠�$i���DP�$M(��a�$�"�kǆJ-�:��S���.�� 
�+#�HZ����9�z=�fk�37q��㉁?���u욯a���(|B8E"I� #�4UBa�=NB@B�IN���XC�TO�.i�D�$���'��}��.jA�ه�S2Y��	Yg�eY2l��0��<�
�P��ǅP0P��a�J+MP�����_O��6R�������Ӻ�C�OLAb&F987%��%5r�`d
O0Ӱ�4YY�Ց�nį��Z�� ,Ja��Z��l�Z@���J?��b������D���f�	 0 s��'�I-RPҌ��J%2�����2	Ϫ7Z�U�"`J�Hޥ��)�禡�p� Kpp��fި��6$9D���"A��@;
�2C�=���""�>�W��}�|0�k7<O������/�,��B�;�D��Q�'�&�;ӯJ�u�� (�R�&d�1"5셒�:��:4�H�
5N�"Y�@A?,4I��C1�J�eH���*Q�?������1�$�ޭx�� 
ф-D�D����H��ʒj�.~&l�j�zx����/1���`K�"~nZJ��aZ!�D�p6�|@�(��$�FC䉪?=VH���;>(�����-�T�]]^��ȝ�ސ��䛹/Z��唧+�~�rP��=.a}⬄���]p�I�x'���cOҧ+�� z�cO�O�,�Ɠ:��U�EC�3q�2C��App�Gz��G�=���'�H��}@����0+�y:b)�3/F���ȓz��ڄ!�2��z��[�8`o��9[���Sj�O�S��MKf�X:^�	Z�!ՆS��I8�!�]�<qH�2IFR1���?!4@���cy�̗
d�~���'J�D�Ռ�~0��F"J��!�
�'�v�2%��Xǒ�HA��;q�,
�'q`�A߅�Y����	�R�2
�'3�U3+P�S�yrc�Ŕ2���
�'q|�@P�����T�3m"=�n�	�'���� T�:@�*��<*�"	�'9ܵ�!�ļg�v�3�&F/p�0!	�'��Y�W��'>E�9ٕ���ti���'��mq�D��.�԰5�� k����'��A�.�� �*���+�'�J��0+H>_��9��Q( �@���'ݤP�vm�]߲�b.P8z\l!�	�'dx�c�.H�E����$g��	�'�Ra���O�a�j /UbL��'���ѡ�Z�'�.��4��=RE�yדOd"m��>��MD8Z��A%(�"z�`!z��y�<1g�͔h�J9����|]�1�� qܓ*Ȉ|�Ѐ9���N��S0\F�	�N10]@r"O�dЖ��Zh�M����h� ���+Ji�qO�P���Y�|��������	fF��צ*D�����ݒ7��ؑ�Nvt��$ǚX�9�>�OHq�fI�i�L����:���J��'���A��6?�L�q�Tę��ͷZ� s�EF{�<!���Id��p#ɴ�<񖪑u�<Q��+RHD���lp�(�q�<AbM�52xLa�ӄ6˰lPrdLr�<�֌�69w޵���8"t@XF�AX�<��,$(e�ɋw�?T���1'R�<!#�o���k%��>6�f<BT�t�<q�@N�wT&� �cD�h�
̙7�x�<y��G�qV���58!���"s�<��F�UW.48㏎�xB���Ys�<Q&�߉-��B0|F �P��f�<ɰ��:g^��G�ԭ}ڈ�h�f�<���ʌk�(��H_	  3�a�h�<qe�V/�Ƞ!3���5�Nպ�+MO�<�oӳ�x=����0B��$�Q��c�<9���=A�L#R�Y'���e�\�<YG	�v� ��V�ev�#��FP�<ɦk՛� M��Ì�@�!��f�<�UL�)��J� 8]b}{���}�<)�7 �@��ըM�鸡�M�|�<1�K�,c����hm�X��`u�<I�'_"8���#˕,m�!����r�<yT(�0
�x�
�'0�̠A�^o�<y��A�jv��>
��(_n�<qՂF�D�0�H[�!yԮ�h�<�0R� �2�0"��T�M�Z�<I <s�j�8E�	q�`=
HS�<A�ݱ]�
aZ)��D:�X�fWO�<���R^�'��X�b�a�r�<� v�iǮ٩����/R��J:�"O܅�s.ܱ?;�@gOВ<d���#"O��3�̽9Sj�(�뚡
Z8=QG"O�ڵ$�=����<0����a"O<��
�	R����qH)��"O��B�:K,��ʥ��%o�iSW"O�4���.\	����dax1��"O8H@5@[�p=���^�	W\�8�"O����3Y��9�ω	q�]ZS"O*��_!��j�iوx�\<h�"OZ��a�0U{�l#�(A��rM�q"O:��	���TB���.[��` �'I2L�g޶,&4q#��v7p�:�'�J�h�l�.x\���%u�<�
�'H�N[�c� hQb�JB�x�b�'s�@%�;j*���Ý9Kx8li�'T�id�<�(Y���5-Ȅ��'�
(�����@7�SQ*\�,mMr�'Zyӳʆ���T�u�Q��~�A�'x��SFȵt�Liť�.E}����'/ 8��%;����[	I��-�'��QJ6�<[+ś�B1H(Ni�'�z�d�b��@2��uY	�'��0F�܂X�ʵ�	�'�	�'�\m�5у/�H�t��2(�ȁq�'�@�3�ۃG/x)��f=��?D�,{0��k6lh��F	�(���1�@0D�l��@_$S�05��jZ�B�"bI-D��C�-���C���5�t�K)D��xA&�"_N��Z�R�`�:t
r�<D�c�@�Ny�F.��)A
��V� D�
6�ƃswvt���L%e��A+�:D�t8'$M!:��"g���V,��6D�;�E�#{ ��WJŎ6G�4D�L LɳZB����-�1c)�=	�*2D��0�OA�R'�"��f
�i�`,3D�<;#�lV�8��K���q�/&D���b+M�H�����El��d.)D�d ���r���B.��,Pq���%�OR�����K����.�8o
���M�<��ެ�pEC߹ ��x*`,_R�<�5�H�g�Z,ɠ�ٛod�邑��b�<���A�:I���>-�9��kC[�<) ��-��˶]O*,HR-N�<�db�br�X��F�9(��W(�M�<I�ܻh�L�q4F
�]rD����L�<A���MÜ�
6
� ��B�JE�<q�؍o����cnE�\6z+0Ō{�<ѷ�۽T��
�瓵M�[�/���JѰђq�F���*ǲ�B��ȓH��2d���Ht8�JIK%Q�N0��FȄ���h��>�D��@EQ�nQ8$�ȓO���;��>�P��&�_08��ȓC�ӄJۄoÔĢ�N#�����Q�d�e�W�V}�XR��B�G��9�ȓ��3�CԍM�vd�p��z|�ȓg����OP�@�Z��7HQ�TޢY���� �q�� e��ц^�X:���ȓ��$�q虴5�zhC��ͣ$��e�ȓZ��"�+��3(l���ͦC�pH�ȓD����JR!WV���o�	.4t�ȓ/8F�ۆ	��QBF͇��؅�I��~"c@< ��.O������y҃�̪) � �:��` (Z�¨O��D�� ��WF��X�D�L�N����e"O>�Җߨy��\�|9��OD`Ez��)Z-T�V(�!�ĿAE�j%N,!�D�/�`f��u�X���@1@�3��|�gZ;�.M�*�|3\��*�yrKX�hk@���F�s��X"�.�y���l���'��=Q`���n��y��Sn�f��G��22;t��G�G�<�I�(�v��M�1Q���r�<��gU;^�Y�t��Q�X!��Oz�<���R�B��,:��M7+�~uN�<!vJ��Rt�Y��h)�ԍ��\L�<�d�Q�;����W##��R7�G�<Q��a*�E��i�
� 3F �D�<�%-��lRA�G���{��um�C�<12�U�y�a��;�X�ږH^t�<Y��1}�7IQ����#Yo�<�5�i�F�)u�B�
�F[v�<�F�'��2 �	.L��&�Y�<AEI�)UD�;�hQ�v�I��J�S�<�� >Wb	�B�ѕ5Epu�vF�x�<q9�89���`K^5��l	x�<���v��@�o�`��XkUc
v�<���è#VD$��كw�~|��j�t�<�6�ԥkz��ׇC�*s�
f��q�<��8%�b�F�ĔdRZvaFF�K���O�����X2"f@{B�̌G5&��'xBq��i�!߄1��ɉ�pȤ�
�'֠SH��W�BhѓEN�lb��
�'�;B�#	���Y G�a2�Ta
�'-ԸQ*�@��|��$!X�|�	�'�����L�Q�� �.^7^�vy��'|�[`l��5�d��oJ�"�Խ�'�*�Z��R)�܀YC�� �����'�,�i�)�)
�"i�7!8Z��' p��V�G���0 ��\���'ͺ���ˍ�}��`b0_�h����'ֆAd�E�@ގL1����h8�'H$E:%J�.�2�:FB �Q��1��'l�����Y*���yi\A:�'��(+d��&f�%�kw>�z
�'���Ye51������>^�܈�	�'b�����2�s�U�rhC	�'��ԋ�"ҢE����򯎣��1	�'^����K;���2���{�(�J�'F��V�S�^�����D�,�
�' ���RL�=Yzހi���=W�P��'����҄8�֭�6*ˌ �4�K�'�<5�'��<N*X�B�P�r���'?6��Qw�YC3�ʍ`$$��
�' 6Eh� dxș�U�ϊ��ݻ
�'4H�:��Q86>��CR(��s��a�	�'��}��g�/N�jUK�K�}Z�K	�'풉�K��^l���D=v�v�C�'�J��QӸIk�M3t���p���'[4��g �
i74��sn�#tw)
�'��L�gphfK� ����'$�EZu�K8(�+�"���'�%�穆��
]1����te��'O��ϕ�|ʪlգ�Fٚ�I	�'�h���GW��-���	�H ��	�'".���,��N��USA��#&ț	�'�z���2o�੗	}ܖ�	�'nj�{�F��K��Q�7�^���	��� �����D�s�|���Տ�* ��"O�J�[1Q��Iv�͠Yw�i�"O|� ��>���h��y��S"OI�����9c.	��X&2����"O ���e��!���R�n�@Y"O�ta����L����j� �X "O�1kT�S?p�T�*�ߗ?�D��p"O�,p����Uz�
a���!��"Orlq���j�剋�M�t<��"Ori����#�\qI�H2�K"O�	㓍F'�����: X1�"Oj��w���&p0W'əb؜c�"O�����L.�4�GGǴ%`�yxu"OzM��IS�-s�[A'>G�a�1O���$�� �T�vtV(�U�^��!���K���B�b� ���h�:h�!�Ď
�#���g�"�AC�#�!�*�u�)R5� �C��Ƙ6�1Oܣ=�|�ף��+��B��ť~dz�����K�<I4�EV�����\��h	��E�<AcU�&�q�M
���VJ�!�dԔz��q!�9 mڙ���Or!��N�0���Zu�׍v��!��'x�!�d̕}��sTj�w����Db�!���)>6�x���%�uB�� `���)�O��QD!�3/�R�YD���C���G"O��A9D�)C����U�w"OB�)���S��)=�,�D"O
+EM�!E4l5��>��,Bg"O�)�@�� $���ƃO��	JG"O )�D
ԏ2J��B�fݲ����$"O��A �+F8�)QHJ�=}����"O�ԋ���S� �R#��
3���"OԐ�DG[�&�6<����nq�T"O���ӏa��p5:�W"O�\s����y�d�ۣ|'���"O���I�T��RGFمy �%"O�3��ۣ��52DE�������"Of�R��.�AdéS���"O:ԃ$%Q&y�Q"c���� �4"O��9Wi�e�,��p��Zm���"O��b�aO.>f�ԑ7"�3h	��"O����/Һ?(��0c/S�kJޅC�"O��#�>�$K#�\�I��
e"O�z�@��Q��x#!��_�"̠�"OFa�l��0���`i�.foV��p"O��9F���� �o.8�"O�lR !�.C@��E�G�y �:�"O�x�')�>9�@�͵z�6�7"O&�J��=2�Q��� `����"O>���D�&!!0m���4"O����6�HXVL��|p "O&�ۄl�eb��qk�=9z0蓢"O��`!@�Z��� �J��O
5� "O ��B�A�(�Y�ܸ&��X��"O�a�8����BB� ��A�"O �����&҆�������"!"O����+�(��Ո� Y�
�&�a�"O���@�D�{UhT1�o�	l8���"O�|{ť۝d�p�XBoE�T7�\��"O~�Bύ5V��uXp-̇B���(�"O�J�X��p3��2EPh�9#"O*���K� k���±�
LF",�%"OvH EA�y1�|�2�Y���Daw"O� Փ �E2|eb*4�)6�`͒�"O�!RlD��i e$�0rQ�"O��@cP�D�R�q�Yu�p���"O��X��ıg�5(A�)��"OV0kp�ٞ7d�I��j���b3"O,u��n̍:c��C1@ʅg�t�1�"Ot��,��'�,{�,����u��"O�1��+͸N���S�%U�
�(h	 "O28���ܙe�,��[�q8��Iu"O$Ѻv,
*E�B`b7"�H%`���"O��ؓbؚn��X"�W�N�b ��"O�T�ӡڤ,xX
W�ӘI�l�A"O���է�=ںh����y����R"O�I�3�J�^�$�����܌:�"O�y��"
;�*���������"O�qBw��n�NQid����P5"O����S�Qĝ$Ɯ
M���P"O��k�O�dT�X�A�`X�u"OvѲ�@�+��Y�w��>gԡ�5"O��i��nJ�hڗ#�-flA"O謈�C�*U=������Rn��"OHZ$)ݦx�Ra�cA�bvh3�"O�A�G��	tv�Ipd�|r��b"O(]��&��{Bt�����PH�䈔"O�}����
3�/P<4!S6"O�)��_M�ؑ4녧=�p�"O
����0e��	�"@N�i�`�E"Ov�3�I�=�nP�.̇@��"Of�kT�_f>�1�,Ⱦ#׬�Bd"O��)4-J�y;(t��?#�]#"O��$�L��;tl��b|M[�"OB)x¥¼Bl@�
�y`,U�"O:��G���a�.e0�̀�|S9Z�"OL�ñC�����['خ�N�[�"Od�y&j�^)� �v�ߓ-}ȵ9�"O��١���*�las���9�QQ�"O��S�g�)�Dr-4zͲ���"O�	�F8i0i�U
ͅ��x�"O���0fԶ��Z�/�ߴ��"O
���L���8���ͻ"�b��b"O,���K�r ,ٛƭ;C�$��2"O}�3��(�l�m�y�"O��x��	ll���WK\xPX�0"O"5ʆO��,;��"nH$)#D"Op��K�:^D�=k!���|ڤ��"O8�c�,�#zx��תԂ`����!"O>�X �5_�ftRf
K$S<"Љ�"O�	�bB��FU2�46Q�G"O<���Ý*7�a���3y���2"OX��ȏ9RkL�3��CZ�$��"O�Q*��A�k���6�S�{�m2�"OH��W�
"&�:��14����"Odd蠀�/&��b��E�%��1��'���3�ݝagH��FܓU���9�'m��j��^&�2ջ��$Y�k�'涰�H��_{J@�aD^%p����'a�����{�X<{�eI�uM5	�'�>��G4B�\���5|�؃�'��])T�]xHp1�б_�����')^���MW�@�ܥ3@i
D���J�'v(��ċR)�|҇�&?�n�1�'��m�-*��7��jc�"�'}�0PC��>TqF�0p�W�e�0A��'5� ��Q�j��I0Sf_5aq�Л��� �h���}��Q-0�̄�q"O|�y¤�	I粅��d��N�e"Or����¡#R�����	��"OF43�aS�^�P �G:7J���"O��cN)�p�B�FUW�8��"O�d�и	�,\�P
,E`@��"O���v-��f�[��_���"O��)tKI+mD$qrW�	�8��@Ӵ"Oxy�)�5qL�a��Nmr.� �"O(��wN-������� y����"O�!3B�';�R�@�Ax����'"O��:�G��QA ,W+x�,���"O���AO:X:�T�)G,�Q�"OvP0��3{Z���\I�U�6"Ob��PD۟�x�L	y�n-��"O���/E2�2�kW�G�*4Z�"Of͚ )Q:-�E[�
��o�X��"OJy�l\��^�ӫ8�0��"O�����|�7nv�`1��~�V��ȓnM>�Bw&>n�sKɄ}��E�ȓ8!�  ¿?����n��7��y��%�(:v���o��| -
	8��لȓuUPT�'  �-8X�����C��ȓrJZ8�3E��
�A�^�����ȓm ��;��Ā�4�T$��JHA�ȓ(D� �����4��13 H�>�V)��W�zPH�>h? mP�e�q2�}�ȓa�x�CG�-+����"`�=Z!z��ȓ	�h��G�`��	�1lE�k9�}��[�R�N�I\���u	%r9T��ȓ^��4'�.L�C�̠c�Դ��%5v��� �Ƹ.1���K4�8D� bFbK5o�E��(�C��tS��:D�h3&T�i ]#��P�qJx��u�5D�P��L��H�Ҕ�ҹ���P�`0D��u��^_>|;1�Koh,�R��"D�(��έq:+��:!fj��#K"D���f�ea�)�#M\���'�$B�I�V@�|�w�ȍ\��b�_���B�ɉ:�c鐑d��e馅��hB�o<��LX$X�� $ݎAd0B�	:rsV84��b�L� ���[�B�I�<Z�H�J'8�-҇*��K��B�ɮGnFTX6����1�BF��\
jC�F
δQCo�:`.����ُA<C�I8U��O���I����`C�Iv3�|b�˲?�����B����B��A`���f�,=����_�n�Pg"O�+Є�7���� �ma�@c"O�e�w���&Ru1��
2�����"O`���͎�@1��r���B1���v"O�q;w,��I�2�0��R37�Hy"Or��0.	�G.�&�^�T�@�"O�:0jC#4N���l^�ߘ�X�"O`XG,��I�m9�	׬�\��G"O>��g�?�:�QI\�pҜ!�""O*��ʹ6��}���S����"O��r#�
�aܾ�Ir	���p�"O��+���V*n|0�mп9��X�4"Ox�0���?�2�+�$;p PD"O���3	Ö<R=k�h@�.,.��"O�4�r�388x覈��""O��ƃJ'Un|��
��@f"O�`i�J�
.��|��!�k�X	��"O� ��Љ1r�L�j)G���E"O΀�+@�#���瘭clBMQ�"O
Հ�J��0����h�9m]�A2��}>�$ �<٬�X�F�������O�=E�@��Ij��I$J£:��ъ`e�?(!�D]��ܜ{�
E�%�D���@�/b�|��'kD} �!����0�Ă�+�jh[	�'^2����B�\��-��@Y�'��pZ�`��f����
� ޱ��'5��!d\�D�x�x�k��z:��'�\��F��	W�`Ca�8EP�z
�'��A�S^jqp��8�C	���y��ږ,ɤ�0We��$��a�
D���>1�O��+��0`K���dͻ6E
L��"O�h`�C_��PlʠEҌu(8,�"O�M���T1%� :PN�".�8`"O� yԅ1R�d���L[�l�N�jW"O,��閅B�8�t��j�Б�"O �,�u�dl!0��9\i�<��"O���GE�qy�9t�(��+v"OV���A]UU���IG�P̀=�����@��,�5[p�EC�Yn ��q�>D��C�4:Jd�X��9R�[ !0D���āW�n�HY�'��[����"D�,X�	Q�*��q�E�Pj�<#2�<y
�(x,��!EZ(Z�x�E/�c_����=�䁢�c�}��0n�.7��?q�b!̱[3�
�{�����/!wq" ��b����S��u�.�aGb�\'tE�ȓ;I�$�ׂ̦vc���R.M�/�8���(���2A$��3!b�A�Y*��]����$�7~J�����O�~Նȓ+zR�S�]8i\<Pc7�ǧ��ȓ[)��g�R�cZ|�"��"o˺����Je2�΁�do萲%A̟jt�l�'�a~2��+���̅�x��C�ާ�yR�m8��\u��D�yr쒶� (c� � �X�c�-�6�yr��D�
��A?��#�R:�yr����1	'O-�  � �ǂ�y�c����3�W�#d|u��nA��>1�O�X���ױ>N�%����ٺ�'mў"~B1��.|�P�A�+����寐�yIF0fGv�"�
����еJ���y�mەv`!�MڤvoP�xU��y��ނ�:�y@�P8��eB�6�y�$M�Qy��q
Լ~�FXE���yR����@��cU1g�əW��?щ��S�j^�3�� ~/�!+vC��%�=�ȓݚ�H�(P�R��
S��;
GtĆȓZ ���^n�Err)�;*�.؅�F�R�*s-ۜVex����K"=���g~b$\;�i�ILlY� �?q���T�$�kjʝ#�����F�{f�مȓ
���(�l����� ��U�h�Hv�׮,�ѓ!�F�^�����W�����5�V�oX�a��$8
�'n�)3FL�ލw��'��}�	�'2��p1�U��8$�Ɂ2�$	�'7z��$�}4m��nK�|-�͢K>����'u1O�`�vLߑ:N�J5�R�K�*�(��	`�Ow�l���<�d�Rگs加 ���!���*� د3\Pe�֓�� {�"O$�RvhB/�!:�B��pv��""O� �yó`�!����b�*p��;A"O�M��^bƠd����9T��廦"O��P��v/d� �0^�j�:�"O�2��
WXJ�i��G�k��uYC��~�OP�H3���:B���h�Lދa���D�vFp��9� \�sP�q!�T�H�mcG"־-������Ca!�D�#$x�&D�4�j�����!�$CPI�r�S4[n�kc+0W�!��;i�V�0T�wS.di� i��{��חaI�l�T��zZ`���'(�'Ca|2BӍ
�6�h����B�O��yҭ�0.���ffD�c���`u
H��hO"��D�! ���@��M"!n� di�6
!�dK9'�x�2�%�,	>��iZ^!� "eVy��T�_���0f�1F�}�,�'���p�ApI�!P���)��0<5gF0]�p����C�kx0��D��hO�?`b��)��K����+�'wgH@��/6��S&ǜw�{3B
�6��ݗ'Qa~�\ j�6�I�^�njD$ָ�y�O��j*�1���޹(�H�I7�F��yrlј,+�p���q'�P�F�T��y���7s��Au�/p�ҹ*ǅ�hO���ıs)�U��(L �AbFn��8��O��=���ḇ�B�+�<�aaC�62w��U"O��+��L>_����/�^���P"O�8���OV��	�v�O&n^��� "O��J%(�8}�=� �G�tR`�[�"O���*[?D���J�1.�b6"O��1�V��P�#J�	M�"	�"OT6� �V|����E�L916l�<	I>�N~���`�=4�xA���C���@$-��y���(��a��P�Kצ\�&@�,�y�o�(�i2��z����ȂN1D���##	�_�`	qK�@G���6T��Kv #L��UJ�A��pJv"OpJ�k��c�^��g-+_��� �"O�x����O�r�*���I��"O2�[䭗�F� y�C-f�nm0�|�'��L25� %��$� �9)�t(s�'B(E"�jѿ-#�5x��j �Q�'>�@yBI�t�*$A'K��_�$��''��j���<���F-ۯI%0���'��U@��4��ږdH&p�*1�*O��7�)ʧ	�.��7�]�#\q�D
\ƦX��p�j<����Q�x3���+s<��ȓ�J%���߳
n����� v4�ȓP�P��GL#u>h馠O�P�.���B� Q(헾~��`2���p��ȓ|�)��� d/e �n/wF�@�ȓs*asa��+�p�G�/D<��'�ў�|
��K�(T\9Yb�8f[r1q�FAd�<a�H�$h�@��qJQ	#ۦ� rBDW�<)��L�
��L�"	��
�SO�<��iPl� �����d��Iyb��P�<q��(J8�X�j���e2f˘M�<!�f��m�p��bL�>c~�s���K�<Y#�ދ�Z�b���\l����ly��'52�|��ˢ8���8�+S��7�O�U�!�dļ��\)���du���XA��'Eў�>�r�$Q� mn�ʣ�W{+�<��/ړ�0|�c.ђ.����υP����^�<QWI�:� �T���j���Q���Y�<� ^��v�
C��SDɌ<�x�h2�'�󤟊wj0	�E:�@%HD�d[!�N>y��!ȭ(�t�HɊj!�Dťq��٢&��;4:\2	T�E>ў���S!��U.�Y?�����<����hO�镽H��}�`�V�|���@�`ՂH�!��%2,��ƭ��O�xS�NZ��!��I4��rM�<P�D d
8�!�D ��(�B���z������!���fa��c`@��Z�NW��!���)<tp�1� ��~�B�c��Z4%!��P>騰�M��z�OW�	o!�dս2�@�QF�
��z�섾ZO!��?�HL��'uF�� +$,@!���(��t,[/s������7mI!�d4Vn�$��8Qflu�f	V�*�!��$%/��A헧!X�����I�	r��Z����䜬=Kl�96%�)vv���]]!�Ą�7O(QF�_�G@@,sM0i!�$�T�\	��^�+�����X��!�D
�m��h��aZ�:�ǘO!�$��;�`:�,�}b�Z0TJ!�d����x"��c�|ԚD$���!�Dݿw"F\�B+l��#dcK)^�!�dY0r2��AS���,�`B�K�1�!����8��%�.��=Q�Ã*!�$ط#�RDKQ�H�j�"��։۞v"!򄌍wb��Q���ikj=�sH�.�!������	FG�U��E8��y��'1O@���5���h��V�H��"O�I�"�F-]��=��L�vq��I!"O�A[�	' �L��J��^1��"OTE�B_�Y'�P���@�d̾1��"O���1G�8K;�љ7��){ƞaY1"Ob�Jg�W4���	���/��yE"OD���-Y({�Pg���h��8�"O�-�v��L���l�%4���@"O6�bV��]j�W��?6�
��V"Oა��v^B�:���cq(�ʳ"O���'� ��G�<X�@��"O������e�������4��p"O�P���[AҨxd��a��,�R"O]I KW��Ѫ�F�Jӈ�P�"O��3�`�^�csş�nҖHs�"O�����p�x-SFą�.m�-�%"Oj$�V
G:㎙�D_3GZ� F�$!LO��ʄ)ϪG:�03��1�؀ZF"O�|�s���"��'I	Lx�$aB"O�dp�É%�h�!!��Hh2"Ov�H'��] �Jr��7�.���"O��[�jI�4U�`���Ñ�ܥڗ"O�%8e G�ahf��` �Y�����'��d�o����I��8�q���.�!�dN-A�p��%PS�h��]�w�!�I6Jh������t2��Jc��z�!�$ã3����S��81��r�"�3!�Ş}��agO2R���܀E!�dcF�pN��qα���I#v!�D��_�n����n{иEf�~�!��v�h� ���/jx�HT!�d�2c��\�vfX�w��[scC�g#!�$N�t\�A��Ib�^�HB�	:`
~�k�LAE���c�#*;2B䉺pz�5Z� �#4\�؉�� �C�)�  [Ώ4^��C���J��"Oֈ���DJ�d0����`�E"O����P�qAG��Uޮ�z�"OT�5oL� ��9ՀPTrfX�C"OlezB.��PJ�+�j�p~�x!"Or�r�F�?W�V�Y�E�<`�"OU��*C6"<Aك��)��j�"O�IҠ,0?j @	&LX�SV!Q�"O��u
�
sn��נFU
2�1�"O z�E��1�,�m�=C��"O��S�����Y��K������"O�Iӯ���|٩V
�(^��p�"Oz,ڣ�H$�X���4���KF"ODȁ�@�YqH� N�h��"O���I̦'�xTz����4��"Ox��A�Q�B:T��`Gi���T"O��0A��.�\d+ n��KXL<��"O0iZ��A��Bˍ^]�K"O���:v� �x�K���HY�q"OXX���/e�iB���:�dГ"O��f(\5вt �&D3)�H��"OdD���_f�8'�2%T �"OYP!�.f�*��@�(eIt"O��A��S7:���UN�Զ	�*Ov����*$ylp��
G�X60Q�'l��Q$'ܲ5�Nɶh���v��'��+'O��i�}񘘋�'ZโT䎧X��+b]�EV\��'@� ��.@���� ��Kzt}�'h����пC���)��2E>��	�'�VY�Ťܟf��iWO����U:	�'̐�×�γy:��ʶʒL��'�>�c�i@�4����`��d� ��'���)�ό�j.�(3���0D9I�'�:�*2ʃ/0;��%�
�
�'��H厙���E�2(�.X3�u;�'���򌞷M�d��$�U��'�abBgLb�~��D�:�2x��'�lq���s.��Q�J`�z�8�'�x�*��(� �DfJ�OF���':�p`d!�1���Z�}�J��'�����ۥ:~�,9�!�,x����'��1�1 ɳD�t�E�٩q	�:�'ڎ+�䞨	�9��R3
����';�0�R�T�Q6�ȥ"(^ ��'�J�5(�J]R�)%T�'����';�c[�IQ�Ł+�($+
�'W�i�C(�2?F���À۹՛	�'h���HܪG��(i�D�4��a��'c:��`@1v�8��6L� wL4���'u�A��L�"����i�H��d.�#9lT2���x�$����0(K���ȓ*��x�%�1L���q�ß7z��;��x�Ǯ,FP�# <�-���\DBDE�5p |� ��J����ȓ^�ޘ����Q�Y����c@ m���.u �jtφP����CGu��Y�(�i�J�#zHp�U8e��T�ȓ�܅���H�k��X��36.X�ȓM���2cD��V@��BB�P(�E�ȓ]�� �cp bR`O�2K�m�ȓ~�$�B`�l��U��)�F�ܠ�ȓ9�j���
��>�!�E#���ȓ|���"�HE~
er��G�\0�Ć�S�? Z��<_����ƇI\�$�7"O��#�h^,��&��;?��"O��g�\�	oh�de�
X�B\)�"O�;*J�:��H��ź`F`�C""O`���#� � @��c6>F|�u"O����NĶ<w�<S`l��'$M*b"O�]h�d�N�^e1��«pjh}A�"OL����38���d�=K�ʰ�3"O
��t��Xo��6�Y7o��p�"O$���L1V��1��L��E���f"O��0b��&)�,q��ů|T�"On�ñH��7U�%�V(B1|��8�"OX��DD� �"5�b�Q��
aI�"O�T�EҶ^ج�Y��J�z� 5A�"Ol�C�_w��C�	�8����"O�-�Ө�.��y��R�A�d�x�"O@|��*Y�qmjaA��Ntv!�'"O��kuK�%
"|)�)M�"b<�z�"O�YCt��"6zX��"�ظ�f�J&"O2�qe�͇��qL�2�T��"O�quj�4HXz�am�06j��K�"O(��Bf�uӠ���+�OY�[D"Ot�q��.D'T!���Ã_P�P�"Or�HE�"u�����C��&6���"OI��!�4pJ��k�U�5N���"O�yx��^0�*��'��6"ORXx�h¶(��5�iW�'Z̀�"OL=ҴF�)%)6	ဃ�M�2�s"O.�f�L��@4�`(��16OZ����L�������]���i'D�L��F��hG�����ϕuTU[��'D�t��o�,i��L�ju:��1D��`��g�-w �j���-D��x#N�%z�M�Q	�d���C�e+D���׭��D�p�R�T�W��XzT�,D�x�r$M��D��үG [�D�Y"�5�O�I 0vƨ�Ɲ�,!BȖ	�*˓�?Q	�1�`	�KL&^1\���`����,�ެArE \�T�!%��)�`\��1V�� &���*�ёSJN*[(�|�ȓj"���	C#Y���u��g ��CG��J��A�B��Q�K��ȓ9�~�e²	�u� ��	vp��S���A)�C��u������!��Y�Pe�,�Hp�V�C�nN�Նȓz��@{�^2AS�`s��!]�2�ȓ��m䌜 	ՠ��1�3Q	jȅȓ!�8���k#�����O�:,����p|��I���@Q�m!�o���4��ȓT�
�
��_�0���G�,Z�T�ȓ	;�0p��W(�\p���/Y�r4�ȓ2q*D��,ɝLF-8�l3V��ȓL��h�����}[��[ǣD��X!��d)���a���Z{�c�@�+�:���"8�K�"oJ����^�t����  L=��'s�e[\i��d�""Oj�1��Lc̽YP4S�:A� �|�)�ӆ"�;�&Tx�B�{FFm��B�49F:��Qf�=�����h�C�ɨ��-+��V&CwBpʗ-%G�C䉫X�H	���/m|ر���ֱ�C�	 H�l ec�9A��u �!�C��8�  �"�.n4���ˆ 6C�I47Β�5��-�,d5$M/ Y0C�)� p���z��$b����7P����"OPKtO�%�\Р��G��H�`"OPR���)�zQ3��.]¼�"O&e
V��X��DB���M��]�B"O�0��@�^�!��i113�	q"O�i 5e�*o�6i�"�P�j�H<��"O��AK�*g>����r�f�c�"O�l�7�r������'q>�P0"O���7D��R*hy(R 	&E2�Ps�"O8������Ud��
��ɶ> Э`W"On�%��T��"D��m�T�"O�8��ėo��4��R/^$`"O�tF�N�N��^43I��c��'�R�'w�dǱO��<��Է/��$��cK!���2����^<>�j�2�"F&��h��D�֦N�z%@P$�5�\�bvn;D�`���l������?`�3�:D�x#�	�$j#�Ȥ*[�P"T�6D���Rg�$}���8�'��~��5y�"D�h��x^ݛ��=-t���* |O���yR�H�F)���lD/Y�\��'�y�@��,@(\��>N������8���0>aP0h�t<����%"Nusq�WK�<	'��LnQ
�iΧP?4�c�IS�<�����Ҽk� �'�pc���O�<	ć̐A}Fx��͑]V����)�b�<I7��W���	RDGh�F�r�]��D��ݟ�Nh`��)S���m�C� )�m�ȓ(�(�N	�4��T� �$�֭�ȓxp�a�FD�e����S,��=񈬅ȓ�,,�'@,o�:���a�#����"-�yIQgO�-~���1d$S���m;�@���S�N!xL�w��1��a���� �K2V;K�5J�p-	T .D�X8Ą��l���#cO19���2S D��1�\�I�@���L��q��K=D�|s	��=n�0����2����W ;D��آ%^
�­���QD���p.D�(a��A8(���ѸX@t5b	*D����S	-k����O/GGX�E�:D�@{G"�!}K
5����kEDe�D�9D����(
B��)KV�v�"F�4D����\ג`I,W�@�a5�p�!��Z�@BVAI���(q'���{r!�'F���#�0*ʵꇍ�s8!��NR�\�Cw�K$T$�A�4�B<{�!�D�nµ9fe3<`�ÅH�!�� \���/Z�)r�IƝtw!�����i3�\>X�~� C	\�S!���)Vtvh�E�7l�~��2	��Py����KC�*�5*�(�[��E.�y�n^2q�*���dF�M���L��y�3LD��Xx��r�E��yBn]0xP��3��x�Ը��\�y��I�1��X`��J[(Щ��D��yr/�<JՆe�n˯Y��X���
����<Y���~��ar�JB癰�`�Ȱ��_�<�#@�lP>�c�&�-u�A�3/EZ�<Y")�]��P��M'G�B�[�PS�<�1G�2S�AC$��3BiC�%�h�<���`��f�T��kŋhh<ѱ�N�mc���Bξ�t����H��x�hY��^Mk���/3���&��(8Q!� 6#��4�9:�E��=A�!�� ��'��9`�bVu�2` �"OL=�pē&shB��t��a�b���"O>U ���*U"B��'�"�b"ON��GČ�>{#�Ph��'i�
U���lJ6A�_5����!]�مƓGȊ������V8*���H$�"��'��Q��o
�c�*tS&E"o�+�Y�<��=I��!1�˩EXn��P��U�<��"	�4	xnG&Rޢ���+�U�<��������,��s���T�<��	U�D(<qm�$+�T)@��j���Q��J��,"ڝboĒ:X*ɇ�i��T�)7��KpDՏV�|�Gr��8C�py��]�7�	h�J��fu��O�����fL<��N6jhx�A���y¯�$%J�I4���d\PAhq�Α�y&��Xp%n��I�(	[�.��y��%`6�=U��D�D㇫��yb���T��"Êj<���OϦ�yR�?�h���L@�]�,-x����y�.rP���Ѥ*'� !�?����"㖴��+ �X"��ŽyOzu�ȓ/�ʃ ���0 �;b��8�ȓl��;��ϘT�t���k��c�
��ȓ�0I���rԪᲠ��8����ȓ;E$X
Ŋ�mS0���i8�'� F{��4Kq����LT�0�Ö�U��y�l�K��0�.��L�1&a��ybD�	����6o�<�h�I�����y2��r����7�����L�y��
_)|�Q�>�� ��D\��y�G����  ]�g��늎�yR W2�ͻq
[ 1���<-�!�ߖ|v����R�<��$@;I��y��	,��÷	�$[;*S&!����C�	�]t�M�G4�@x���G(C�I<|�l�#����-����CƄKP�B�ɮ8���Dl��.Mtm�Bh��]{PB�I�U�Q� ��ua�K��W)<B�	��ftɁىY�ڙ���vc&��ȓP?jT��)��P� +$ȥ�ȓ`DqAC==���vG��T+��ȓFp`a᠁��W���G���~�ju�ȓl	�H�$~n�k��ډl�|q�����٤���tE��	��1\5��0�x����ʩgs&�R@�U��x�����B�I�g��jG%N�w2����D2����mHpl5��b��(�Q��"OdIR�ν_d�P��CR���B��'��"��b̛�&�gw|0���>L^!�D�L�zl��9xj"ٹ�(�8c!�K2�f�sbf�"YE��fǴW!���C^\��UK@ra��E&7�!�d\Gľh�AɄ�o&$���<�!�$�0`R|��J�y�DY���-�!�dάY��-PԀ+�q�7H@%�IM��8�5��X
M��9��$Ӥ"D���ф�%U*v$�K�0��8�G"D��Cab�OPM�#JG6�z�!�n=D�p�T?-iJ���._�R豆<D��q�	ɾa%��xq"�=aCFYc��;��z��̋#�%K�lHdÄ�p�F�8ړ�0|"�g*^$y�dʈQr 3�ALC�<�ƯA��8+��S���\ �.f�<� �ٲ����P��0T��"OJ���$��GfY�Z��\�"ORt��y�Ӈ� D����1"O>Ȩ�Y9	A��
AaT(B���r"O*}�aa��C�F0���G�bD
E"Of���&
hl]�p/��~��V�\����KY�U����@����FN����?1��	���ZV�.#���[���5!�Ć�[��0#Eo��-��Q�/M	3!�$ͷY�3G��k�m2Q蝖V5!���A��<	�nʩW��(7��&B�{b�dW�;����0EQ Q��P��eѸ&!�¦�8��&�e3VuXi�k�̟Ї�j�L���)9渺�/�
)���$��G{�����7V��e!��0CR1��	�+�y���j�D!�����5 �p�I��y�@��,���T�vL�h���[��yU�j�
��[�]J��7J����<���$�3�R0*�V?��yBF͈.!Y!�R#>f���vG��k��E�QK� �!���h4Y��`1" ��#��3���)�'4��e"�;bp��:F"�73@����'ل`+�M@�LJ� �fI$T�I��';HY;֍�&E�Hp2B��j��}�'�
�ذEۖ�D$��xA�$��'?�@�W�T4��Q�S�)r��'w��ElK�~�v4���/&1���'tH�Ā�0�PBuj���#n�<�d�R��ZAb�/�W4
5��g�<�SS�Sb$Mq�&��v���B�g�<a委'tl}��F�� �+6�Ed�<���Q�"�(M�aɽ2�ԴۂMSf�<)gi�&~]��!7�Q2<op�CgE�e��v���O�F-�m"j+ؤ�Š�li�eS	�'Ӑ�Pw	>#�4��t�X�b)l��	�'5��1���3�N�!�&`�`��'c��'t)4=[�,���i
�'a��7�R�	ř2Ǚ8it&�s	�'�h�ңm@'H�L�B2��b���Z	�':\�퉨^���{�g�T8.��(O6�=E���m��9y � �`��̹���yB��5NQ	�+P�	@���)ژ�hO������`B�d��*���'�a�!�D�$X�$
�`R�鸬���ؗ Y!�$[ W�rX9��"؞��ⅎ�!�D�)T۬�Rƅ�,;[���b��Y�!�$��R��i�CΘ5PR:�0�O#J�!�.P�@+Y��$�w� .a3�'�a|��M!ٖ�A��f������ �?�)Or��D��
�x���Ֆ/Ch�I���d�!��ݵV?|��!O
/#>�s�3 �!�Z)��M�#M F�WEڦ(�!�ċ�=�N��G�V Q�_]f!�$��"����ʎ'
pb7��1B+�O�=��x �������9�	��F���(D�XQg	ٜ����C
\�ia�8D��{��g��8��y� 1��"6D�0r M�$*����'�0�(@�3D��I1痈�p�&I
� !$�?D����E�x��Eh�8\���%0D�8���J �@@rg��#�, �.D���Id��@{���2֬��"9D��[��.z�,�f����V��O�C�əs�h�v�_�2϶`�	�S�<C�)� �����Y�N�h��Z�l4�PQR"O1�N�)+��f�ëwu��(v"O�r�Q,gq�4rvb�C���"O�<���7!��ԛp"�~�-��"O:���/
�D�t����Thi��Z�"O����@�8L������P;c�zH*�"O�����b�Ex4�	�P�V1�F"Oh�9�m��^h�p��2	��-s�"Oܨ�@�:�Ơ"-�t�aC"O�	q�̝�7�&�ځ�f�^-Ȃ"O(�)#l
T�80�Y�C��
7O���� թP��s��-_D�z�H&D�쁓O�r>Rlb5��<E��p��#D���
 7@��9�vI�:6�`��"D���$�M]H� �$��-\����?D���ЛO�t���J���9!�=D�<9 ��Tz~i)�C+#���4n<D�H; �	&����m�09�E3�k:ړ�0|��/�0�<��%5�NղD�z�<	fӄ!`q�eaU��Z��t�<�Q�A��h�W��E�(����s�<�'C�%azLB�LBd�JKq�<��ߋO�LԚ�f��
��$��ME�<��C�T0|����$6��	���C�<�3/��:DJ�h
�.1��F��A�<YRm�>3!�![G	�,ߜ��PB�<a�Sz���so��E4��"�B�h�<y�G(3Z��
�"nU$�b�<����~�$��G��m�b�a�^�<Y��X�c&r��E�Y*ɲeOM[�<�p/�2 MF�P�g��6HR���*�Z�<��ד
yH���D
�2*`�ѲCZ�<	p�B(u�f �2$ 9�f���bUq�<�ÍO2D�� ��7Ń�A�i�<�g@�)�`���)�2+ت��e�<Y��C�|B����V�(�dAH�<�ǃ��xz�l�2b�|1@/�i�<)$�6�rQ��T�`�NH�v#��<�%�ė	����$AA &2����o~�<���G	%X`,JE�'(x�@H�FU�<!U��9
�<��!CEH����_y�<����d+��)p��T  9����q�<�H���Fa�H�r����
Mk�<	#) G�I��Ȁ%=�ɐ��b�<��� 25�`�3 ����H[�<�e��]P~t�ԫ���9�l�<���)\!V�0�*��c<��h��n�<� ѭL>H�j&a޼?�.<p% U�<)S�@ Sr@Mѣ�H	f�34�R�<Ɇ`̢&Dt%1B`�j�H�+P,�O�<a�B&��J!��x����NS�<�`bO؜�sm_�ZTT%�'t�<9P��z���a7�T��9�D�s�<��ʋ���T�@_=Wex���q�<Y
��Z��%
�;;�m���n�<1NQ�wR0��#�33��!�BD�<��K�;~�r\(	3ń_�,f|��M�؄��"T�n���D�CZ�Ʌȓ"�D���G��0�%��a�VԄȓn���"��
0��`�Um�x4��5����H*
!�U��2𦹅ȓcPXM�Ƀ�*��C�>]/p�ȓ=���jbhZ0UL��bB�I��NL��.Y,�/)�M��H�/a�}-!��  ����D�i캀�uJ�I����T"OY@�"�#T�@ô.V�J���{D"O|H�`�.i��,Nw��}p"Oxh���\�S� �J�" �"1"Od)4��TO��2l��U�ؠ�"OhV�2(T�2aG��e!\!��VC�<!c�6v��4ف畱CF�$�o|�<��#�5��Bc�0C��
%h_x�<�C�(@�\�łP��V(�SIUu�<96DS�5Rp��iO>4�vHe�v�<�Ǫ�T<����=`��Eep�<i�kţ'��C��ɱJ��dAg��o�<���9 2(�)�� -r`H��i�<�˜�
�Bm��Ɠ{�d��
�i�<)թ��DJ�d36�ȕ$��m:S�~�<�)Wh ����I;~��A7�Xw�<�W��hbf�4Q�d@�f�<�R7j�2�*�4o 2%ۦ�t�<s��%��䑣�\�VohXJ�	Cr�<�%�" /܁"�� �^�:U�o�<qa떼���Z`M�r����	�@�<	��@(�$�"KR�� `�E�<I��.H~.t�ҏ]E`�@B$FC�<1C��*Xt�Z�`T m:�L0�t�<I���o������:s���k���F�<�Ʃ٘3�ԃ� �a�p��4 �Y�<!�AV�7l�z�/FOy��!��K�<I�+�
=v��"���*����Jc�<�sL<q�-��M�@B�!�ō�F�<�։Å[�]�`��!EDl���<9G�[/��t�M�8b�T
�A�<��iڻeF>E
 @OZ,�y�%X�<9 Ϙ
GD�P���1�8����~�<�W���&�2L��IR��OA�<�t��3\�xXg7J4����Q@�<AR+�p�x5���/�PAa�C��9VL�ْlЪ^��P0@@(��B�	� v+a���`������B�	�H�&t���:�\EK&+нt{�B�	>H�`�*���liF�%�#BZ,C�ɑ8�P��@a��)gԉ��K>
{�B�	�e��FI��-5��b���.D�B�I�k�B]K��'�D,S��@�=bJC�I<e��J�G��r�TyV�^�6C�I4	�8�Y�Eb,E ����`8.C�ɏnȢ�MVi���ի�<z�B�	&<3�	�D�A�4q���f�%I,C䉓<����.B��8j��D�p��C䉕!y(@�D�\m�A��!$�C��S�@�R��W��5�s�J��C�<!e����iA�F�t���.U^�$C�	�z� 5���=fYF 5�6��B�I�_>-2���4�$�Ძ��d7�B��5[��i[@�&O�����O��B�/I��Ae�U�T���C�pm�B�ɼw�q/�!��4��V�bJC�-^��ar`$>j��p�<�C�	,��1�rjΌ���)S�[ �C䉊`��i��Nw������}�dB�	X�� P��Վ0?�@�aDPY�.B䉾P@D�0��C=����ϐ8H�B�ɯb��P�cB�C��ݸG��})8C�I-H#pk!K�e-x���ɒ])�B��-�(�ӆ�H29~��#�'ƒ{޶B�)� �DML�2L��4��F�ZQ�"O�\c��CM��Y��M�@�(�!�"O���`ūN�qǔ�Y�d���"OYh��'g������Q�ZR�"O���n gs"ґ	��Q�B"O����. r��b���n%��"OvAc�a�'�Zu�)R�8����u"O�`9Շ�;o'","1��f����"O��r1k�*.���R�]�2����"O��ef�)�)��,]�P}�"O�%��F?�j]�*fM�"O��ʣ��x�ԅ��E�<|'�%�C"O"�yr�:3�ssD�K�
�"OB䋡
,�r��Ud�d3f9��"O��
�`��6ͺ��%�_:��"Ovkf�]�^Q�@�O�,�8��"O �S�$B�5�ڜ�.�U^I%"O����'��e��� !��!��S2"O����]�v�^xZ�Ʌ��<���"O��*@G�D:�z�F�TC8�x "Oj����/l:l@��-��B1"O��`s%@w:v��-\+2�c"Or +��b�h��T� �p�"OV�S�#W.6&`2��!wk�!��"O֡!W��3����&GA
�õ"O ,I6��]O�bV�b8R�Y�"Oz������,(!!�%E6`�X�"O�[�I�	�v �Ra�m�`u��"OZ��6`�GZ6j�̔Ȑ�"OУa�ܰB��Q�N��t0D�,�amF�0��Y�a�\R9�s3�3D��	Kq�\[�o�� �U+V 1D��[ǦԄzb�@G���+��c�#D������-U��H�`�}���UJ=D��A3�
�K�Tao�#��� �@1D����JQ!68��k�N�Cz�(Iҍ/D���3FH�f��2�OB����C9D�p2�f	"��lC��d@�LH1�7D���3╳h�`�GI�=	�x�i��6T��@�ם��	j$aC-'@T!�"O�I��'�<G
�9' �8Or�T	u"Ob݈ŭ8Bj.����V,xw�Di�"O}�e�C�xia��_d�H�a "OfI1�''rg�p��1{2m��"O�U�"fW�Y���ANN�]��P��"O�	�H�7,|��"�+Ⱥ��X�6"O��j�гesDy�)���d��"O���B	H7 ,p36�̇kqX�0"OP9`��M91���M:j�x��$"OX�@u��V6>%�FAԮW�Ј�ȓe�C6$�	�0�� $  ���`�l�'舾X":ɳ��	�|��q��M���1���J�8�	Ȝ:��ȓ ���jAl�F<�.�&2N9�ȓe�>��I�!��9�A/�����s�`<���ƬF��tj >P�2�O��=�"�h�5Zu()b��I4�셃g.GU�<�J�ITT��'�#��a#�g�T�<����Z����	��rQp�����QX�$Ey�&�@1��ޫYH J�m��y��߸g_�!�ł*NQ>5�w�N�����hO��~D0g�O�+∢�#5�Θ��'ֱOD\����t�ֱ�B��ۜ�@&"O��q��6fF�d:�#O�V]�"O� ����LN$Y}�4��
�-6N�ˣ�i��d��:�aB���g�.�y�A�>t��D=�$�<��'Ή'ܛ��S�*�VD
t��(����`	ϵ�yrn��:��XU(z�bHX`�2�p<���$��0Ex���O�K�P�@\(A�a~*p?9��CԔ���Z�S&*1I��^{�<Ql�� y^�0���&+r[�5�t�<Y"�=B��D�B���pX���x�<afI67	�U{�*��� ��d �. �`r����OZmrc�U�5�YqTƕ�U
�i��"OL�@l�R��!��G�j�� J�O>ꓧ�=A�A�Ha
� pdM�%H��^z�|�@	6` �	`ܼ��G�_lP�*e�6+����脴u*|�փ�(+��d�� *D�(�A
�*�:�a�G�<{��)Ԋh�֣=E�ܴ	�#3��/�4H�!�O�p����hO��6�$o���JPlH�/FF����a�0��e"OԨ��J5� a:%��;��t���d!�S�'x�$�H��=Љ�����E'2���II?q�GXy<"4F��{hh���J��0=�5E՗s�1���J�Q�R�2�MJ�'n"�}���%?�*�a�T�x
��zbJ��6(����^����b���T��L�r �6C��R�'w�D$/�*MZ5�D#�pj��
��C�I�f����-ż ���T�	pؾ�'5a}(ۙ8�@qy��ԅr��Q�&��-�y2�K�~��h�G
�9=v-�f����y�*�����j�%2kP����\,�y��\=D�t�d+^tlR'����ynа&&(rm
�?qH�[���7�y"K��u9�5r+�01��,x%�A��ynQ�96|��eT�]�0Hj�R�y""W��XDi�nR�JCDe�D�� �y�E�/E�����o�"Fj��1���y�C�����S��l�)�A���x��|f�����~�(y�F�a�tB�I3.��q�S��;��U	�rf�B�M�ё�ۃ4Ï��#��B䉦V,@A�e����*Q!�h��gN2�IZ�&&y���Śjd��ȓ|\j�zUc�� ��ÂM/J^!��i�Ty�&$��XR\k�LIh)8T�� ��xۣ��)+ph�3�))[P�ȓU���J�ى��0�g�#v���ȓK,��sQ"A�r��)񁘞.{���<��ƥG�Fw�������X��>1�a�ڔ|!aCY�E�����u�{0�RD�A#XP�=�ȓ�J��F�+�0m���F�q�L��ȓ��$�����$�F���5�4�ȓ&[@{�@�d�Fa�m��O�@��U��8�6`�0Lo�� �%_�,*�`�ȓ*B��e�\������G�n��̄ȓ�$A���[ 	)2���J�>���ȓy�hl����2T�Eha�_�G1���N_`T!�A
!L�> �]9R��؆ȓ#�b c�*M�'�L�cHQ�_[��ȓ"��)ɇE|�P5��'Pr1�ȓLP�lx�h �Tm�`Z�j\�+�n�ȓe��D�!�)�A�%bC0$8���]2T�0eF Q[f���O�iC��ȓ[��1#�O�+�,����ap��ȓ|%�#o��@7��OP�ؚy�ȓ+z��Ą�#t����I^�s����S�? �t+���<�p�p%��B:� �"O���f�Z�f��Q2���;Y��K�"OR �7�O.
�"��(؆a�~܀"O�Ej�`�l��D�ֆž j�"OH�X%NR�)j�̛�c�d�#"O��AF���^��+�aTp(�"O�L�F��4J^T��K@�c=܉B#"O�@�gMǖq�R	N$
+:a:"O�,R&- 4s�;�(�$&�M�V"Ozɱ5�\�#��X:5I�b�<���8LOfaj�gZ��Ⴂ���s�x\�"O`�SF!�p1�8��c����D"O��S�L�TW� M��%�@u{��'n�tS��(x�lmI��X� ���I�&D���T�.nn�"�)�8D��=�v):<O�#<9T�H�^Xa�u� �_���ZRn�[�<q���f�,2@˕�!F�	S��FX���0=� #Jc�R�e��R�<ݹ��S�<�F�_�8���W��*ߞ�Y磘ԟ ���s4r\��&�'E�5��WF���XW���f�� <���Ģ�*v),��t"O ̹�A��$&�a��#f}X��e�'lQ��cN�gvT����&x��$9`n!D�(�t��;�L-"#^�}�05Z��?D�l0Ъ�9I�
�w,������"D�@3�"��+�:��
Z>Fz��2'�+D��RǢЌ|v	�v k��R�#D�x	ύ(m��ԛǥƘ\r���"D��S'	�4,f�9TLƹu��%҇sӜz�)��)c�!��:A�þwG6����4D��*Rk��	֒ܪ����9��+�<�`�'���H�

��|]�f�]��~2&�Jb���#X q�� ��>a@�7�,}�i���=�T�'����`�S�0��j�Ö�b�]��'Ѫ��C�Ұ}�U��ݨRR���'�����añ�����F���������'
Ni�7 ���D�R��qO*��d�Ct
ر�"�1ώA�����5�a|�|B��9�KRTc�9:�J]�yB�9	Af4K�3H��ag����$�<����?�G�"'!�IG$P ��S��8D����� ?%��Cp'��y�HxK7D� b©�-݂=3�ˣY8�r!/7��G}��OP�?�X2A�:B,��S'���_�j]y A��0��I�*m���'�~����p�� D�꓁�'�Ӷ~�qO��@��M���j��j�\�$"OH@:����fE���7j
�K�<@a2�'�	f�S�O�.�h �.{+�`���>;�i�6�'Hў�0Q�@�}j��J�Ĝ1��0ɗ�s��Il��O�Ƀ���:��hƟ)��Y��'a�V��t��k\���
"�O>�8�9�B�OC�I&;CI��	Pu<H�c.�8��<�����'�6ţEڳ/�آ���!c5F!�ȓ_���X�&��EO�M2(M5��Iw��'��T?����TR�
�F	�6�d���@�eE!��P=�"uAt'(;�>�	�i�)�?��S���DAd���e�ȘQ�JE���[��!��r.)X��8��m�b&ٛ>�!��8#lq�Q�@.Q�8�ITlD�|�Q� D{*��$�0!�1b�RQ�`	E�F}pT"O�t����&�μ"k��*��E"W��I����r��>2�tH'�N�T]�ų�E��yz��(u��&z�`D�utp|�ȓ]�툓�0���b�.L��S�? ���O�F%�1��`�MRv��"O���%	�'1T\�+�/�� r �q"OPtz�k�w�tA��%?��yv"Oԫ��<>�m#�ݯ:r`�"OšAj�U�~�c�A )tQ04"Oj�
C.���T��/�	%̡�"O���ąoN�Q��X��r"O�=C5gp`����,G��(f"O�a�mѻVc���Ƥ�;#˲p*�*O�(!`KJ(Ь�ȑk�3�i��'b����G�"H<�!��ԃ5����'���K�V��!q*B�-yl�H�'r��A��^�0ODK /�#��ĉ�'�P�!�j�:T��nT�	2v�@�'��я���UlȢnn
]p
�'���aꛖw���g-?k��5I
�';8�"Ӆ>�vQW�V6��'��7�_"��m�1!�z���S�'\��r&�#d�X�PM�o� ���'��i����*StR��ܨ��'!R����M;(Zթ��D
��aQ�'U�e�S���E[*I˦"��}<�y�'_Nl����8��YK� _+(@.�
�'|Tĸ��*�\��ۥh���
�'�$|ktG�)4�@ذD�O�c��� �'Ć�tM�VJr�AA�آ_0n!z�'�,#�
�$9`H|����Q"P4c
�'$�ĸW��_��eP`�%z�hi	�'b2]CQMO�X�Q�G�ƿ~���C�'h�k���>�b�s'��/wL
Ȱ�'ؐ��&�@M8�H�lж���'`,y$d��v�*]���ʩ׎(���Ĕ8|�* bS+];gf��-�sV��d�*j�T��4��w�Q���N��y"�S�vF�y����6kf��y��D�b����J��D�`�@�y8i!j�r�,�:@vH����Й�ycD}����⋻FG��7)I�yr�I�q��i��V�GN�2׬��y��|�
1�Ǭ�2.�%��a��y"	9}H�b!L�j4�Y�����y�:*6�2���48Z�������y��� ��x�H�.`7D���Ԛ�yИ^����t��4��́B��yBh��X�L����/�p������yr�٩o� 0Yщ�Lި���ø�yү��F�])FI��D���Z�j�y�ፁI��p	�N��<2���'�I��yR��:�jH;�OG7[	"��s�I�y���;WvLԳ!uHLs���6�!�$�1%n���K�ر�$�%6�!�䊽(��'gE8�Fp����,�!�^Zd I��pn�\��H�e�!�D� `?�ݒp �,!YNx ��Z�e!���-V��ȉ�J��@�a��q�!���rxv��V ">����R� �!�D�h��*���&}�q�ͣq!�d!(�Vd*�D�N���B���a�!�$�5R����#&�U�d=� o�!򤋡:&�uwnX�Z�
,�����>�!���n&�.֢b�`H5�)�!�d /l|���"a|��r�L�'F!���W���+��� ��`��Z�< !��e;��gł�5bz<�'��m�!�d�a�ڝ��c��gf�)O�!�� ��pAnM�]�d�H�]�hzZa�"O��r�B�=��i��>}��3d"O"��P��?��u���H�hU��"O���¥�CN��#cì*����G����7u�����
=K(���l�,oO���u(��=�!�J1 ��%�g#� ���z��_#.f� +�
R�	#/bQ>˓�:��rbP"(m��	D��':2�!�ȓiJ����/g.0)�h���İp�j�0�Z��"�O�͛���T�� �Bճ�T�t�'�V�X�a�����-}�eGE0:�l,J&��A��ȓ9��S�"w�Ԉ���\�(��<���@	Z�0��C�:���ma��ѼQĨ]�/�u�H��ȓ2)����� _��Z�k\�-6�Jc��i�''Ppb��t��̔�',2�p@H�\Y�F�9D�d3<�kD�`�褘�!ڶ1'� �c�1DV�|�M�{K �y�BRf�Tv����0=aq��q�M�(��e�	�+���e�2j�"��Uo�9�fC�!N���rc�ӃH���B��Q�Tc��+���W�@ʔ���H�f�Җ�I4ƞ�X����!�j��"O��HA�T��hH�@Y�:�z%H�K�,N\s�,�~�����I9#ԈmA� V56�V�)B��81�C�ɣF�b� �S�C��q��8vyB9z��֙,���������E���6��C��=Mm�m�뉹n����R��CI� V>Z4v��"䶙��X�E�!��JM��|q���e��+��O�ek�!ʩ->,�s��%ʧAT�����2
M����K�E���ȓ0P�<��j= �H}sp&�^�$SeL1.�~�;b�4}��9Or!� ڞ\q�)r쟃F$�b�"Ov���2���!��V162Ƞ�4O8�`MMW�`�	�d.�g�ŊM����ǁO89��I�=pd��	A3��us�5]V�" ��H	���gl<D���2���1��Ȁ"�����U���=�_�б�b)-�H�м2�؋D4���Fk��}	W"O*-���3EXEP .��H�`�yt�iszs�(Ck�S��M�A�ٴ��yr�8&w���G|�<�u���|��,)6&\���Ug�z�<Aӫ���������Q±[��v�<�J��U��5aWË�w�L����m�<�G �(C�T�puˏ�J�0:�a_j�<ib�� b����ǅ��00��ȓ��y�+�?M����,���A��!����af�-��@p,M?nXB%�ȓo\v��� iw|4�& M\��ȓ?,T|�x�ӄ��'����}�j���1�
�pE�=E"���ȓ/s$�Ӏ�)~�kCȏ-Q��Յȓ|��t�w�;w,��1*K�L�,���:�5�`��R���A��,�lu��REvh{Q�L�C$!;� .xy��.¸)�À�5' z�R^�l��MFi�<��(W#.IJ�e΁,��lrv��}�<q�x���zdY�$�d�2)�~�<	�!��}� ��B�3��h��i�u�<���\��ƍ�/s��}S��q�<�����!
�i��+��7�Hi��"O�C�K�����a�%�� �ر��"OH�8B%
��UC&c��a[N0��"O��� �7|^�9c���%``}�#"OM�&=ِ 7
W�}p8R"O­����X}\� �Q�p@����"Ojq1 )K�[r8(��/�$9��C�"O�d�Y>6Z$9ӯ��"$�t�2"O�p��9pQ
��[0{"%��"O�5K��)y��t����G$ �%"O� &X��O�y��Mxգݶt����"O���p���@�?9��H �"Oxd`��܎t���逇Y���X7"O��"0��������2��Pc�"O����cN�fR��O�p�f�[�"O��	�o1�X�MƤF@�u�dP��j!H��a{�ÿ)Z(K��f\�I��
�9�p>A��U䦵��OJ-i�-��h2L�ef��C�	-k�a��V�IS�ݙg`��<�&�k3��6M1O$�{Ǎ7O{`��e���OsĘ��=M ����UӈY���ǔt�>��.�S
��0�.�+��	^=
7\��P���Y���(!�b�%�g}�LޮPl<���M&4��h3	����ٜi<����9��)�'HF�@(bjڰICȈ:$��5M:�n��	ADY+V�ȘR�h���)C8�����ݧNu:,)�!T���rA�k�D�(@���/��Od�B�"eǮd0R*uw�,*��	t�Ș"�ϡTlC4�O"°>1ֈ��B��E�f"Z)�p{!LN�3�hD�f�ٶm#��Md�Ÿ�M�h�Rhku��l,�c>!��Q�W�,�a��eiB�� 9�I�l���䘏8���f]9�C�&��s������	��75 �9�:C��-AA��1�>��'���k��Q�Cw|1��G�)q�O&	�C�;I5Ĝ O�"}:ցʫUD%���;G�`�fP�c����e� Ҁ�+ġ�k�3���$mz9�I֤q~�tva��f��'������Cg���Y���I[w:+� &h
b��լ��T�����X�2�^�
�֭^Ψ����Y�t%[���H�E����=P�v�H-v� ��)OB��!�X"`����
�v�0�A/4�	Y$ ~�A6$��Y@�)���X�6�џ�YԦ�
*b�|����mvP+��!~�����1X�* �F�$%�"�g���G�dQ� ����+hS0� ��?Q12�Zd�%?IaF�`�"|J���e�tY# nWx,j טT>��a�l��nU�G�ãux�A��dS�
�tap7�:W�PGF�:NV�$�@E��RG:3X�y����~2����8'ĵ��R�H\: �S��2,t���)�2;1@��m�D���?��N�?r�J���$#dp�3V唖*��gQ.�bY2��cVJ]�"	�z�j�M�!ax�E�׼k$�ĕ\cʌ8v䞿'�(�PT�Fx��@� E5BH�c,��"�ͻKq�h��gVqr!�&ӛ,�Ь�$�φyzby0w�Wd"��r΍{�'<<���
1[(|��e_��b���D � 8�����@�w#��[�擊:�(�c|���䜢�7M�gq�Yғa�b���sD�!O|̉6�\�;�R嚰�V�U�XX�·�i���냮T�l|�8È�S�hС[?IHs�ǫn	&�j��N5X�u�Ä:;J �p�P�g�^���iW(<1�CQ6 �v�S� � o,,�j�NY>F4
U[�HG�'�<���-S����Q��x�s��Ol��b������fe�Bw�e1'gRb��{b'pu(9q6(����b��߀I2`�@r�e��IG'.a�1��#�'��D�:;kt�@��':D4��y�ɍtH�e�g�|9X�XP����'	���R����$��[;2�b���*��)A/`L쫧o/�d�OY�t�"�$��x�4�J��f؞$�$�F.N64�z�e�)L�*��
�KxrԂģ*^��$H�O�j=���.O40�R�'� ��Jv����Y�
��ߣpޤuJ�E!D��r�F@"g��g˝G������Uh
���ۂ{���'�� �1�M��x���Ѷe\R� @�*�bޠ)���LV������8��P ���B�>$qԀ�
]J*�l!^f�pP&~}rIĒG�`�c� 1S�	
`��/�HO���ߴe�R��5��	q����r���RV:�	>j�x�X%�.��%��hDI�
"86��/9G���A����cю��>)`/�t7VК����̊E��%���Ay�E,8�� 왅]\ҽ(@�q;N�ʈy��h�ɒq&��؛U�J�ل�z��b3�ҋ���� 60գ��imfUj�!۠pμ�ObAR!��vĲ�0����y�σ���Y!si�mfx�;'iB�p>�1����� ���8��)��Z������ُr�6�'�d��CGư�>qB`��<⑞Ī��T�6���Y� J)P�z���k/O0���-�#RH�\}r�*�
��#܀�j�m�����<�h@�2$[�\��	���?�4$����s�Q���tNL�'�24�h
A?Y���Y첨O>���$�I�F�g����M�M�LC�	�j��H�u')fn,̩w�N�<�x�;@%[3��=��S�O:J�r�kK���*#m�d��'�f��Bb%�D�:�/�d���IK>1�oJe����d
V2D�$I �<�I�	�XW!�Ӝ)R��CǤ	bb�a?�$k�<a`���J����$���Ĕ`@��k�<���K��!JE��
�P$��JNo�<� �#Rϟ�!��8��E#u;�u�T"O�P	�ϯ"��=�d�N�����`"O�ڔ��=G&�5��n�d�pUK#"O�UK�g�rيA!BM �{��u! "O�� �]�0J�͛͆�dG$��c"O$=�Gd�!"5�	��O�lN��KA"O���b�~�Z�*�GV.��"O*��4��$&"V�rH�>ga��"O�aa"#����)r%ޅ|�`2"O����Q�E����W�Ҽ!��"O��Ϟ�	��p��.�Z�˳"O���e܍9�F�KE��rzB� �"OJI)��@p����OadDp�"O���+Z'E��+�2nL�
"O�P3s�׊pU��K�FK�5��"Ot)� eV	GjԌ����#FM$�P"O�l��ϔ�jX3�ʌr��U"O�1�1A���Q�Ӄ/���8C"O <���L�/��E�R�ٲeW�,�7"O<豄d&�\{gܽh%��d"O�ܘ�d�2�>	I5l�)L��"OHɶJH ��8�F7D�0�Ȳ"O���QQ�"1�,Q�*�8<)\��@"O�h3�CTz3YH#�ĩ�!�$ �9�d!�j\�r.țz�!�d.R����w*���p�4)�!� �P�p�^�WX,Bs���r�!�d�5r� س��[;TxsE�#+~!�$H�V4�XQ���s�}�`Η*m�!�Ӿ���AM]���C��5�!�b`R�P5��MN� ���_�!�d�	\<ç�W�*��h�!�4!򤂛l��P��͔r�浰��H�h�!��t*�y��FH
3����1R�!�$�w8�h)�M�	>Fd�C"�"2!�DP�L(d����qvD�@L�8 !��_XE!��78��Ik*�1]�!�Z9s�A!��^�0�A��<�!�D�I�x�V$�'s�d@{�h�*P!��ʳ��-�'��{؀ݙb��]k!��U���Ĺ$]U�L`1�Ǡz!�d�-N�*����ڔ$'j���e�3GZ!�d� `�0P�����1�\#J:!�\�<��8�M�#��!�!�	�J!�d�?�^L�7H��:J��S���)�Py".M08�a���Y5�T9�2�@-�y��%p��gM� �`��E��yR@Ѽ}�hB��2z+B��'���y�¬G�0�1+�"B�d���M��yB�ւn�n���иBR���W�C�y�	�?o���T��+0i����'��y�&d� m`6D\1�YK����y�.ݝ+��h��Q4z�����C��yBh���Yq�QD��p����y2ۦ����G�=�V���ߓ�yB�N(�Qٲ���#��M1����yr
�`j������W��Ŋ���y��?E��uV��>EӮ��#䜓�y���5eՊ��7AE:��C���ybe������,�#�6Q*3�̦�y�)�*QӢ<d�Q-h�L��"���y�+I�Z�Z q!��c`�g�-�y2l_�S����ރd�]�1���y�#ɖ<�&��Je,Fl�q��y
� �q�z+�]�)�0!I���W"O`q�aЋ\��\���!^��`�u"O ��+�AP|z4��q��k�"O01�+O�6���xe�֏�Ұ��"O����A�$j�NPa��=>�����"O�ukA;$�"�: �*`*6�k`"O��i��×C6>�Y0
�. �Q�"Ot�1�+H�P�p�� �cRa5���U@ۉ��:xǖ��"g����QYwϒ�!�d"P�j�pw�BRd�@I�n�5��5*��FN�I�4�Q>˓u������7�X��D�5)����ȓ6������V�AtbӯD���`#��&��'K%�O�UjCE�y���rE� ���1U�'�@m���ÂV�����7DT�t'��K���@�[�J����9ӆU9"�$iˈ�x�Б>�T�<iBBP�8�L%�c-8�GԤ�)�Ю[N�	SV�R{P}��(�^�2��
;%��I�R`(!�RjT� ��'��L��|[	��iǰ�&cG9NK��b(D�$���S !E���.�7I\9��Ȃm�(5p���L��|©٬^�	�SL�� �pp��0=9�,[T��� ��?��'��.&����?%��<��CAC�<�4#�^ ���A�K�����e̓J��ٛ�l�M6���B��q�2�1���;@l�`� C�ɸ%P� `�k�_S���R$�pSP���́5����%�O���3?`� �[��̢�h��LI��0�~�<��H1	� 4��^�4��ŽQ.�[��E��)�u.\OLq� ���'�PT��a�h��Q"�'�`�� ��`h� 	�� ����w�4+*���OŎ��9�ȓY��T��I�sm`�
lV���>1�B�j9~�c�E�&�(���&��UY0�1&�k�����"Oa�����D)��"��m!�P�*�-�q����)��<��陶&�Z=0�қY�;�"r�<����6�F����f�F��a��<y��+A<YF)$\O4�81U>a��eR5�� +��m���'M�e�/�L����(u��� � 2y�ģD���y�L���跨�%�dKt	��(O��WB��"}ƭK�Ȕ��҉]�.��8¤�y�<�R��$��!�ˍm'�d�Φ��@#qO?7�a��Њ���-1ni�0�JE�!���*�6�<�xM	�$�4�B�ȓ ��%:j����T��L�ȓ�p� �O�n�8+N�dD�ل�$��9����&7�B��!n��e�ȓ!
������\#��%�>���+g�pK��qpx�d�J>}p���k����3d*�xCȚ;4���j^H{�4l�a��e��m�����"P�'���e�ư[.����d|pCC�,���ѲI�G^D���,�(��� [ x� Ĺ�٤H�dԄȓ����"Q�#�������;�ȓg�8
 UZs�"/W	1X�ȓmCּ�c��&�\��#�N�3��ȓh@\�Q��3����E\�_` �ȓ/h�i���u�4��&j���ȓ|�Q���8}%���m�Yc|E��2H�Y
eL�]�0�`��V��m��#��]�#Ԑvm	��1:Ɓ��*�H�cQI��G�t�[���%Ңp���8���K��o���s�m�"*vbԆ�!8�B����H9w�Vm�:����P!S�گ:��4%�$F��ȓx���k��_(:�H����gl���h��
M;\@�ժU�xC�)� �a�a�ԑF�j��/дSp���p"Or��AY�05��5�1fr(�"OV�Aηr��K�(`�d�w"OTE��cʈC10�@i₡�"O楙!H�<� Q���U3Wt�|Z"O�bp!�� "[%�X=Q�R�i1"O�����h
F��c'ھ/W�C�"O8�d"Su��d�֧�a5����"O�%�+[�\^��UC�7C"`)�"O|dQ��F0�Hl�DƬ5��,+�"O��ڧo�:~�H�H�dW;�c"O���􎗗RV~��!�OJ7D@:O�ɪ��s�*0��N��'��K����8�'�d��C�A�bT�H�j]SM�Ē�����Ht�qu!�S�EX�\!�f[�"�5a��Ҧ`�B�l(�x ؓ~-��%N��z�a�Sq��3r@ӧH��\��N�e�9�m��:ْ%R�"O�u@��?����u�D���I�8}�k�6��q�@=����O!Up�	��pAh�B��D 7;a����Z8*�n�%7R����ӡj�r��o��W�U���*�x�
Ƌߜ�2a;�DY2�&"?A�c�2X��t��I;�i� e����H�A��Xq�I�M!����rJ
�'N�����5��	�RUD���.��S�Oᠠ�R��b��P�T�"m����'�~iAV
^�3=�]��
>�ti�ǜ>�V�Oy2z�⠟��}�f�4ޔbSᖖ$���iqd����?92�MoJ���ㇻj;@5#�XW!�h��	�u�̼HT+�/;����ݹc�j�E�bQ,V�����0y�%�p��$=�:ԫffE�
m!�$^�6u�A���\/�����gN_2�ɹ_>>����$�Ԙh �Z7g�`J�CL*u*B�I>hF��&�����DMG=���4Xbr���-�$k��0���H_�OHh�)ג$.ҵp�\߈��'p�`5L��LM�H��LKC>�G��Tǀ]�ĤK V�$�tD�����IY��06��jұ�v�P�0� ����2����ʇr6 (��e{��25+Lx��d��a<�ip�g:�O�H��Q�H���*���Wj�Mt�I�'��T3�&&z��T{�iUϧ<����:KK���`k\�.5��ȓF����D@:HX�/�y,��i��ɫ-O�#@��)�:��"ΟC���F����P�ɦØ�P����L����ȓ����­��)B`�Q�Q�J�+٨��RD<-%�����|��-�Z�'��	��a�=:?\�� 윹+9�<���ā��CN18��!�T��-���vK�HNڑ�$R,$}�ŸK�+j����'�f)�#n�U�'g$=����w$Ts K�/��q�ҥ��;D�`:4���`�����U(��4�",fg�&.�SE�BC�A�!Bcs��@�"�O�ě��r�Vm�t��I�Lk��l7�QqW�'L ����5e��Ћ���s�RyΓL�Hk&?�0-zs�Z�*D�"h�Ȭٓ"O<Qr%@Rr����KP02�f��V��{ �W|����k0?i��
��p�cסcl*�
�m��PxLGq����$e�/@Nr�	�0|O"�:D��F�E@��F���ʇ�")�,:4,�5�B� !��e�ܽ1Q(��J�Gz�o=�:u�Ɋ�<�$$�Ŵ��'�l�ض^~�i���L~�Y�S�kg�e�'�Џ.�̴�@��!<�2ey�����2)M�t���-o�� ��̞��Ё�a	ɧ-&��I���]s�����h��B�-n��� Lv���
�M��a�˘p R��2D���5	�Y��)�'�V dgV<4D_��M�1��B�R�z��|+عG�L�*��M�b���ϻG,hh�ŧ���Դb�CC�xLv���'�9��Q
��pᖭ�I�b�ȣB�r�8S�>����h	"� F��-ڸ=K���I�\��0!�" ����A�
P�ax򍇈
�y47OP��t��+�xUY���K���룎۾{���JWw-��t�'�v#&h��g���sc~8� K�41ǆ^B��D�`�xC�+)��O� ���.��csh^�w�L�+�'��TqW�"~������ѦWX,���O�G��?|�4�O�>m�S��%v���0䞺uhX�r3`>D����6N����i�=-{R��#�>�DZ=,yV���S�? ���td�N���֢��!��B"O�p�BH�=_���� B���E31"O"��b�<rF�i����
�D�"O�| ��%N�h	��( ��0���"OP�飢	�(�0&�9� ��"O�m#g�m�Vdx��O0B� `B"O~U�E� �)����S'�"]�"O��
�Śbz�a*$K�b���iW"O�i�e��mL�8��U,}��j�"O���&!.Ȱ�@'E� ot���"O	��"�4I� �:��=<`��"O��)�ȗ9f�V8Q�B]�=�T"O��� )&(*�a��FV��t"O:�{��ϣEצd񂯉hO}ȗ"O ���P2_Ȑ|�R�s-,qC�"O��pd��&�rp�gM�'Er��"O�}˕�[�=�&���D�"O��璏8^�e�(S�IÖ"O*�����L��Q��҉Y��,9�"O`�&��0F΀+#BH%���d"O�5�k�;5�:<q2�+� %�`"O֝�g,�3����Oژ���R"O�u�T����d��Q�ɠ	Ep�;�"O�4��ɓvƪ ��h�3|q"c"O�%Q��"f�ɻ��W�|����"Ob��V�����bT�"����2"O���&��1C���rW L��k�"O|��� *1�4����)��a)D"O�H jÈ��x �тY�t��"ORA�Ҷy�Z ��Q�M�L���"Ot1�r���2�Z1�_��	JW"Ox�J$dA�V>Z���m�D�FD�"O����Z$ۤ�붎Ѿz`Ƚ�U"O5��*,#.݊$k׮W��;�"ON��*B
ɨ���ʟ	a-��)�"O���&%�9�*�w�J�(a�\Y"Oz �`G�[f@�iQeXF�hs4"O�l�B��l^�0��Y�{N�,3@"OZ��1���g�8�;�`υ����5OD5Fj�?D�`�Gl�"IPD����I*F��EX1�!�ȁp�
֔YBvB�.|E�G�	�p��:�h�/tB�I&/��e��'����D���P%H2B�	6mg�RA%��4� HR9<C�	$I�V$ö�M+qT@p9Wd��6u�C��'sAN-Ccm��i��eX%Y�H/�C�:Y ���MS�Q�/�:~�,B�	�;��l"DȣK���̉�n�"B�I�f�Bd�1�:M����LȤ.��B��MnV)걫T��( 4$Ȃl��B��2u�pH$mB*k�0e��fC�I�9��]���O�l^���gO�,�ZC�	�iX��ѳ��"��B�gèJ�TC�	���i�a�;6�a����k�^B�	�Kn�`x�JL�{�j!�v��6m�(��D�v}�-@"[�LAj��?]>�x���*�ē�xz�D5�)�ӣb&�V�^�t4���@E#o���j�H����?�)�'+�腘�k�pS��ză�	I�doZ=�|I���S4���u�_���rÌ�R7^A��H�P��0|�(�nJ�h�Ȁ�YIV H�cB���'���@��>a�M�r�#�N�x�Ju)3�aܓ�hO�O�J��R����0�lCY6&��'���ŀIl�0CS%ƣW�̙��'o}q����\�܀@_�Q���+�'��4;�L}��B��U�H�pk��� F����'� ����!~U.|��"O�ب�	hP��uʆ�AS�9�P"OX4R���HSN�b)��%>����"Ol۴f��o���b�͚C1.m�v"Oh�
r/��Q�<Ӆ�� 1�Y[3"O��)1eK7y��"Ѕ+xJ,�"O82� O�_HLRË�9�U�"O�93
�<c�hu�F˓��52p"Ob���ݎk�A�@�1�h�ra"Oz�	�l��~����Ȩy)F��"OFT;��\�9@^	�d�/<'0�*�"O�MHR�X�5���D�8�����"O����*�İ�E��)�TY�g"O�a����e`��e"��%��"O��������<�g���Vt\�CD"O,*!,[1^�āj��j�P�v"ONE��i��\LE�tB�2�h�P�"O�U��h��s�Н���� ��� �"O��3��"*Kb @�+ܔ9� �"O���_0��+֧�V6]y�"O�=	d�2[N��#��Q��2"O�Ճ���7u�e@�*ό]F���"O<|��(��?�|%r7�Ĝ;_��;�"O�L@wHZ��~9q1"��W<-pp"O�x ǭ�-R���׀S�U.<h1"O��&OK94��RD�٠>�ᙠ"O~��pbX� b���n�L3�"OF��d�ȍ��!#?!)��"O� ��ۘ�xhTl�O�B�"O�SgCG�Y�u*�[8d��"O@ B�恤s ܽ�`����"O��z�D	zO<c�`03D�� "O�}xaMɉ;/D��;I*�ɛ"Odт�I��7���Z�R��t��"O�
�n߂b�ȓO#6�|�"Ol�ag2X�<��!��/�6��"O��Cd����� ��#{R�)�"O�|��ӪRP1f�����c�"O�\Q6�Σpє��rʁ��"O�聦A�0U�=��hZ	g��;�"O�рPg&0��1�����z�02"O�уS�3^ S�#�	J��%��"O�A���*6�<aա���,���"O��F�Ks�y�e.�1�u�g"O�ٻ�_�6�T��,
�*�D���"OP���|t�E�s�J�J���1"O�̺�����t���!7��K "O���L��;���AB;��q"O�(��Ҥ2;�Xڠ _�
9 ��"O�僵��eF�UiV�U�yb`i�"O��)Si:1�T�kwd�w���"O�5��G*3���2T$�u��"Oh���ϷG ���D�-i:��"ODI��RSl�͠RdY+��i�"OFU�t%_� q	EA2��(Җ"O�@B�ꈓ2!�(�ԍ�x��B`"O,���) &�{�Lυ2�2$�b"O��#ǩW9	}p	�`�#oH�s"OVԁ�D��h��B�";�Y�"OH̳Th�"n�zP�#N��Rx��"OT��옓~�u�%��  �@9�"Ofpp¦��	W��&쀀)Y����"O��3�ǚ*h;h|B)�>9��b"O>��6��z�h�@i�8m;8h�"O� �]�H��N�1����#�D�6"O�pX��M�I�,��"��$y���"O�,X$�4@��yS�V-`h9��"O��mG��`Y8#
���U�6"O���Ei� ��� q��6DF"O�r���'�8���@&S�6��"O�1�f��J��xBdE�d�����"O�qT��-d;���cK~�H��yr���-���oJ�m���UG�yr�	�4W^�J��\� ��UC��K�yBF�7^X��SMP�gxbb�D�y�kM�XA�h��_�(gj 1�AX��y�&��Q�e=o�\��]��y�b�&Y�&iU��7Zq�H"G�	�y�"Ռ#DV�+�M�O�*eC��߫�y2��S��ӄ��M�x<���y��4��Y@�͎GU��D
�yZ�={%��,U"dS	��̈́��،���G>~i�iqw� #��ȓ?�t8�ʊ��I��
�n��ȓGC�9����)K��H� Ո�Z��ȓʆ�
�*�MU��������"a�ȓR���P)�,cl��!^0�����T� �����h�h��t�ȓ���a�ȋ{���a��..D�p���V�xܡ�IЬK��:s&+D����� �do�M{��M�BP��@�*D��ɰ��V�؀`�+����<�;D�x��];\�.��p�+ ��uct*.D�P��$oa��G-.���BW���B�ɊpY�,��
�b�"�CfG����B�I�-�\(���">-�Iɣ����B�:Z����6�@>���0�����B�I�b����/T�^��{�-I:^��B�I�N
�)�',�V���31��5�B�ɳ_6��oʮ`�%A ΏGlB�	lᶱ�4,����aK��d�B䉔Z%)�#�b�U�$A�9#�B�	{rE�L�}r|	�SO�!"$TC�ɢc�Шgʙ94�r
R�E�	?hC�	�&I�1j�*r��d�։i$�0��"Oؠ�"b�)BO�L�կ��9�ɑ"O��JD�tb�jA���<�r�R�"O�aR�O��8���*s����	Xd"Oh�	�N�h�*���9��4�#"Oh�""8���s���(C��h�"O�����Q�,y�@��Mx7"O�Y��X302Lx)�,��}^�U"OV�2��p�-q�a�Y���6"On!���W�[v\Zq"ݱ`l�d"O�3� �45��}��U�XR��"O<�1����p��9�f��7"Oz�R6@�t�(h�v��$V�����"O$��0O#���i�G�2ֲP @"ODt�h�"�p�B�`����Q"O�5��$�Wt�@�$��>P3�ሔ"O?H�J9��nU( ԥ�"�0b!�<H��B*30j�%���#w[!��3wABu�F7 ^
: &/P:!���lx���q�0RY�L�����J�!��Q�ap��@���9G:���S�J)�!�D]	2��˟�T)>M�EGy�!��+|��e*��H"���õd!�	&�8�Ȣ��#n(��1@ªX|!�� ���� ,@�4�2� ���0��"Odl8�o� ��=xU�	�*�`��"O�͠ ��q2��e��tS�"Oġ��+�mC���8�,��r"OZl:BŶa���FN�Nr1c"OV)�3`I,� ����B�3"OR�Ǆ�$a�}����)�v,�"O�Ya�Š�\�5Q�m�f1J�"Ol��JЯ;B�B	��J�d"O"��ǎ3
�1)!��P���W"OD��RU����&}�b�"Or�QA�S<��ً��R�i����W"Oθؗ닥yv� Q��T��Z�"O��훷9�b �(́�@���"O��x��G<�y�CҸs�H�"Od��6	G�?��	s��7�N�80"O\E�P�U�ܰu��*�̰�"Oa*��s����-��:�ND�G"O6d�"��)i�hLj�5,*Q"O�tb��/�&���".+���*�"O���Cީ[��TX���5U2
D"O����e�^��9���?!Nh��"O��XƉ��/�R%"N�aCR�:w"OXE[�hC$'�j���o%��a"O����M�;O������1v4�%"O\�@�f��F`ȕSt�9K�H�v"O Q��b��Q1υ,re+&�y"�I�V����ٿd�ƹY�*M��y�BsԬA�LV a[J��eV��yr� U�|�'��
Uvr��-���y2�%j �����BL)j�8Q&N��y�� A�ݛ3	�xמ���I��y⫘2}��	ׯ�;�Ҝ��N%�yb�A&mn �8��K8��}��DJ6�yB,�M�� �%� *?�|X�oE��y2��&0M�)g�C81��<�g��yr'�:���6K�<;RfF�y���4�01���ȴ����Z+�y���ovvmI�hE/ ,��!�
�y")Q?j�v@�a�L
�;sAɃ�y2MË0�1b�
�C@�h����y�M� 6��e8bo1+�*hL��y��(%��Y�V��3G�9"Aũ�yB��1�G�1q��ɔ�O�y����5x`ba�]�Q=���C�y" y�Lh�¡�Y�8l5���y�jQ�j\��F)�@������yB-�)x��5X��2J��h�`���y����b��G�=;]�5����=�y�f�Y%�mȷ�BL�C2��y2����AqE �zx��!�'�y�`V�w������0p��ڲ�!�y��8-�hh@�
62�����&�y��ȋ :��W�M3��
l��y�@���u9��H�-��|����PybM�� �*5"��F�S%�K�<�'�o�!x.Ec$2�k��m�<�7�¼mNj����	pF��ףG@�<)r���5����U� #���-V�<Y�Ǝ��n�C�cW� B�EK�O�<A��O�1�p�KVҞ	9�N�<)$��$� ���#�� Fa�e�<Q4�T�׌�x�)�vct�p�a�<�`-2�����^eD���_d�<� ��J�B>F# �K��]�1�l��!"O�e�֢Q �����Na����*O���dF6R	JQ"��T�R}�
�'R��K��λ)�j�H6E��N�T�'a�$�   ��{m�NHW�<!����SH�eIvcE'y�D�#�$SF�<sB�|��5���	�[��_�<q�A��]B5a�U���H���W�<��$�{���C � ����a)JM�<�q���ugR��DK/�lh�!�R�<�U��	J�V|�@��:>�Z�H�n�P�<�7�Ć_�j�90`�����N�<��C;J6�*��gV�����J�<��K����~|�D�e��jE��_����jѥi��i���r
 ��ȓZ��0!T�˔"t��h���?� ��!cvD��K:��ݠ�A�)B�ȓ
.l!7j�(a:��Tc��<�J��Z̰q�d�F�\���߀_�0��F��� �G�^d󤍘��y��^Vp��ē?[�e3���?4�r�ȓqiD(��1>�h��4 D4eXXɄ�+I<��!��/�:%ئQ`*L�b$Rmd���J�jɄ�	-0���W�g� �[e�	�{_lB�	r�@�j��ԕ+}�i�Ǝ�n>�C�	�/3.ب���?
Sz�1vFz��C��*N%��0a�"P�}PD�>f��C�ɬ@:X���+f�P���/x�C�	����z�ɛ�<�+d)�5w�`C�2� �7&�i�����5!tB�	� rc�N/0����ǘV�>�I���V�<d��aݝ��+,�
.� H"A�' f���� W%X�H�BI ��҃\Z�hI~��� ��hA�J<�(b���(�J�2e�YI?	G)P�u��AiE�֩�0|:�!�0 9I���I\"�:��ܦa�F@�'�R��#�Z6�)�'������k����F��<b���勄)���� �:l֝�3�����0�Ov:e��I޽"��0Z3��$I��q��n���#b�N�ѓɗ<�O�q�FD���ۿ`lDL؆��T���sB?���'cRmxf��I>�	ӋF��lR.����N_~���q7�[\>���&=�-�alƜ:�d��b��4��N�c2��y6�|ʟ�=�Н����>�(�+�%�����x :l���өnQ<Q E�K(g	CK��<>d���S����u��4�d�S/��U[*�A@(A�TͰ�h�"O��҂��]U��(a���]!���"O$�K4��W=n�n��(M��"O2�Jbn�!~bMn�T�5	�#D� C���5���\�-�x�rO!D�$Îͭo���� �Ja$u�>D��Ap�×t��c�ժb�VU0#'D��0�˟��b]���T�9�KU�9D���ӈ��:�|�"-��py�Q3��6D��;qG�2	�&�{1�OzY�1��?D�h鷀�&lɊ%��hٲ��i��B>D�(�vg��s��Y���Y�={�%Q6�<D����KߞCv8�Tʘ9PҌi2��&D�<����"h�A�ŬE�(I;t�/D�P���
	nrm�qG��aJ���"1D��C�
�*K*50��O_H�	fn-D� qV�̙F�4IS��zW�$��c8D�$K�g�y�<tC��?�U`S 5D�Xb��U/=�2<�k-l�@v�1D���B"�^�*MK�-�p��M1D��3���J߆�:�Ĉ %����J;D��;��#G�(�8�C,39�
��7D� ���޲ys<�"�莔 t4D��8#�ߠU��9����f^f[�=D�<(���a��!�!��P�V���7D����>(Қ|�Ԥ[$luT�Ť2D����!W�B���A�W>{$�#�+D� 4DĉG}ޕkǎ�,L���AG"/D��K ��4{�(P��E�ot 08gE,D�̣��m5�v�B�k���xg�(D�d�d�@*/M�<q���$FB�+b�&D��h��	]"5����0LS�!��($D��i��M2L�>}a���|���t�!D��+�J�n]K�M�bM�VE-D�(+��	[��k�ǝTD�5�tN-D�L��E9�;`�*K�)х D�H"��U�$����#��A�yI?D����@�OK�ЙgEٛ8���`WH<D�\:��:LDK����R�����@?D����$B�Y�jK� �Az��RD<D�t�EW��8pd��ހ�ra@:D��*���sX���ЂP~��	e7D�h#oS�V�D�f�	�S�dC䉴"��1Y�R$	`M@�A�x)�C�!/�@xy!gDtX*��Q�yR�C�I��@h��#<n,�۵�C�30�C�^U��x�ʏ�(��ӧ�?f�~C�I��^�3�\�#���h^F�|C�	v�j(P7�� X.ڬ�A�o>C�I�Bf"�q�I a�L
f��"� C�ɂ6����F#2�����T��C��2c#����jU&��WB԰|��B�?s��)�ˉ����ʀC�I)
�H1��=+� �%΄[�@B�ɝPl��:���.P�zt����z�8B�)� ��s�d�?h�LH���/CZ���`"O��[&]mʠX6́=3R�4��"OB��+ �y��q�P%WM^81q"O4�J�JR�s����1+�$yG,��"O`���ҷt�0����4���@"O|�$M3�T1�*N H��`+�"O�)à�	:E������ɫ[���b#"ONA�"˘n8�uZA�T��EP1"O\a�
N��Y��LZ V�޸�k�<�ĕ��P	��Z�b�I�OQ�<ihR4b��8t�0_q0P1s �E�<��#�u�"<#C�σ�L�A�B�<q��
[�V�j�V�W縰I�G�<q�h O�}�'e��f�f2%��l�<�$����1n��W�I3d�^�<����Qo^����8�%k�B�<i��ܩih����ĒurQ!�&H�<9f�G*-�Z�5�Z2�DAw@i�<) ��-��8��n�&�H�-@y�<��D�[(�!�χ^`֨h�/^r�<��G�
��5*�6l@���g�<�R+d�0�"Z�P�pᥣLK�<�MG&����Q�Ll�<	��	��	�W,I�W�>uʠ�B�<A�z�6��СP�@�N��łt�<��֦E�n���lH2Jvd��L�o�<��+�?v������E�Z�1��g�j�<	�F��Bm�])rͮrht��#�d�<Y'�9R�l}!���~�TM��_�<� z��`kQ$8��Y�]	!�].uw0��'���T��)'��g7!�Z�e�����+:����\3#�!�$^'f$X	�GE%P�ǎ��!���E�ҙ����G4౧�R&t!���w8
�'��Nd�H�W��hK!�gĴ���3AcRY�fFN@!�D�<X�`����a�naad��Z!�d��,k�|KV,(5��
P���9A!�DX�!y�m�D��*�!�b�*!� <|�J��>�Љ�+ۖF�!����tmc�c]<O��4YPK� 	�!��i��	�KB?�j�Q�	��#"!�DA�.��`��~�R��5�Mr!�Q)O���A�E�/��U����A�!�d4cMp�!o�3���-�<�!��C܀hK���<�|��"�\!�T�7/��7!	�v��1d�J� \!����8�JՒc�4U)�$}7!��Ɓc����°-d����*I�F3!�$�=7i����f�;[���	���*'!����~��3CE�u�hء&	��j�!�d�� O�ڶ��g���ѨN �!�D�B���t�_��|��]�!��:z�TA@6%.I5v@p��"#�!�$�)4�c���}v,=��F�^�!���8K�쫲խwuԽ"���&	�!��	���+ 	�gk�tR4!A�]�!�H�^)��ÒA�4?L����Ə�!�� P�Q�Ԡ�($>���`��Et!�$W)q� �����|tO@�SR!��RBX�q"��>rh�y ��N�k!��u��Q�'!B�?��	�B�ԧ1!��>:�"18B��P�JA���_�7f!�$W���)灇�J�9YQ��;!k!�� �4��'V Ēl�E�I�Ҏ�s�"O ��g�E���p(@]>1�hL#�"OT���k�5=���e�M/4<��5"O�*�6�z!��N�K(�XP"O�e[�ǂ�X�lɲ@$+vQ��"O�ȩ7�%�ҍ��E*>���"ON��_?�<���.��U�"O����B:l� 9��`S�n�zD�@"OFA��H�*���3��_�>��6"O����g�X��'�7q�8�@"OJ�� ^�I�$���_2P�����"O~�#	��^�P�F�r���C�"O,|G�ǂ{LYh���8b$H�"O��j��%�txq�տ%���"O��3�B�2f��(cD�[!&��v"O�K��h|
y DSy�-�"O������2j߸�����&n� 0��"Of �g�͙;�c���.Pz�鑇"O�I�%�3� ����`ي�3�"OtQC���	�|I�������ؑ�"O�E���
 }�`y����z�¨�W"OVpbqo�2\ʨYg� n���s"O6y!�!�.#A��c�#](8�����"O�}O<��h���C�kuZ��"O|bq�U?��}�����\N4�F"O�}�Ң�\�l)D�
����"O0�+҄V�QJ1�2d�(VQ`��"On՛�"aڲd�����(��"O�!�tl��]'qk��C�=�> ��"O09e@��k���{�B��\�h���"O8$ʐC�V��他��48�>5��"O�=P��o�.Q���5+��+A"O��w&�%͒ {��K�'4��"OV[�[�0Sd�pV�l̉�"O,���!TN����V4��r"O��ч'��[������R�ij��C"OjAi�*Gs���'Hï^�4�S�"O>a�� ��!a�W�3��4CE�T��y�HX'2�DY�Bђ)��u�s�'�y�,�b��}PV#K^
�Hd��y��܏l�1�P�L�>==��$X6�y�h��J��u��E]d�Ձ��y�	��Ai�u���>>7�i�����y�Īe�DR���/?e�qQ�bK5�yB��TG�� R
O;z��2dJ��yrF�5�M�ɑ�U6��c�y�΃�-$�xc�KB�x�h}��)��yBd F���w�G1#��j�JW��yb慖J׸��v@"#��}�ń�y"��_�<h�$�ϨC<p�˄�ǖ�y�9k�0��i�V�Ʉ�]�y��,��]	�
�Z� A����yrfԐw�܍@�C�VKHU��':�yb�g�6��0�șK�KB���y�
�O(a�!-٤���M��yr@�_4��s���t�)�r��y�\��,��rd�1jG���솨�yN�9wh�ʅ	�f/nh[����y�� �-xc���6�fL�a��y"g@�x~��@�@��| v�"�F�yb�̉�x����h�"��3퍻�yR����>`ˤ���Iط�y���(b��]�#�V<G^ISA���y�"!��,I��I�t�2��C\��y
� �:`,W=:�rHC�,A+*�ȍb"Oح�q)٬yU2��pMV�����"O ]�G�ŤkΒQʗ�'�q��"On���à_W0\����k��8he"O� r�@36��7����D���"OJ�SE�O.����A�W"Z�f�"O��EPQ��-!!!ގ,͎���"O>��"Ǚ�q(Xp��@' ����"OJd��e�<(���O
1A�c�"O��s/�7b���3�`P�U3��#�"Oֈ��R#T��P`�7L̰��"O��@"#��x�@$�&6�@��"O�e��M{<�Ҕ�-x�4"Op�J�
��팑 �A�=Sb�aYr"O�L��B�K�R�I7A��a�(Yc"O��d#ݍv�@��`
A@^6���"O��JL	xix��0^���"O@d�˞�-F((���UZ°�5"O�<��c�H�xEH���0D�pK�"O�Y��D�H&L� (ǰu@>h��"O�\��   �<� E5_�xH3�ǀ>�yB/B='�BtŇ�I�8���+�����ʎd�fA�a'��O �c���4:x���@) �F� S"{��E���Ț�~"⇙��GxR�\�~��u�mL+ R�i��R�	NVi�W�w�̼F}2��ti&��ĕ'{4ҍ̪�x�!��F�'�V�0Ê�z��a�-c[�O��:�슎2E�����D�'h�d�(�2w�N����90��+�8;vY���B��"E��c@��ħx@)�V@,@'�Q�_�ES���l��RԂNv��ӧ����`���2r��K$�����F(^
"�$#�Mѻ I�	;�k�j��OC�!{��LR}r`H�Z�Z�i1��\�E*�+���DƱ4/���4�װ��O� 2)�u�Y�k�H�L ���>9 G!�#���4�DS�"��� ���'pr0.B94�\�ȁ��y�gn�%@��)R��o|���!�v��A*�M�7�H�q`�jxf�zƄ �G�r��E�T������	�7���8���C�JJT��i	"2�<����T�LY��''�ܴ�`��Ua&y�p��(D:Bȍ�(�OJ�*�/̓S�LTjB 1�4=�	�'p��p�D؛z*g��$7	.q����4I����gR"t�Ls����'q�l"3��>	A*GѼL����^�:�x��R��$�O��
�L��׈�|�ܱ�u�X&��� Dy�<�G�]Z�yjA, 	������R�{ �d�Q	�m��ɚ�H#O8�#����HU�|���%E���1iD�l�>I���G${0(L���ԼtLP�f�3�O�PF��7qW�,;��� �␘r�>QV"ӕ@>��	Q��)��|��J�d%4c>�W#˓b�pmX��3G�l���9D� ���\�-8F%0N�,R~�b4J�h��=��T��	h��~2$V�nø	�̡f����Ɉ��y��O,[:��LI_:��uـ�?��#ќ(ǌ���c,lO2����Q�y�\h����W��@�%�'Є(U�
�\�8�n�<��I�ƙr.�W�P�{�TB�ɤo���h(0��@g���0⟘�CBǀO��-���ӾCr*)�w�[1+���p1�"O��Bc���9��qC�1I�*L�F-0\����]��"�g?���".2P3�c�/*s��r�Vo�<�Q�K�\�M;P��%^*r�F�`�	�Y�Q B�$_+a{�?w�j�
"d�z �0P���0>	��r8n  ��\��YA��8d��3͝-rc(��ȓI��u*��ީ_����J�}�B�Ey"iԟH��qF��GQJ�@)G������!��y��5
q�4�e��H�ƛ��yb+ߣs���:$�PX�r�a��y2��R�r��GC���¢���'AZlq�N}����+�f��<B�K��B��Ih6�9�����.*#*R�)�	2żI���[7�h��r�`��� ��T��H�*a�LM�I�6���	1S�.ђ�-V14��O): �F+�*R�J]8�E �W 9��')�઀�8/���5i��K ~�/O��ҶbU�d�"��M��|�A%8AnTt�	٩��`��u��\�ae�8H�"�����%0��35���&���>�7��7ET !�1�\Lx�JΎ���+��b��F~�_�Rw|T�土��Ė=E�ތ: ��YR-Y��Idid*�)Qa"���Qs�(z�.�V�I�X�j���5���� f�:ʓPv� ��1 S���pYC�4ttf\zOU�$Z(��"O�(�-?h��ٗ	7D���0�Q�`�V�^=%���GC�F�iȿ@�	"�Ϧ>1��έ3��<xv�5,�@ +GM~��i㏉�=��4��iJ�+0���Ԯ�s�����Ȓ*����v�����_uF�"?q���%-UH�B0d�p@H��g��X�'�"D��eU)Dܕ)'���<Ha�Z�H����_g��CS�S�*�����@���C�
P\B�[c66�*)�.���:����9��ן�p%�K/"±1p�i�5��ĳ�g?l^jH�E���:�.,;�O�̓��ԃ�_ {�h  cZ�'��Qh�"�O����0��bO��"�t�<�l;�#ۊ"��`���IZ!wL�YH��b)��D�g	k��-�6a�ڟ6���S^�,��坾{d᱃��*� ���xQ��S���9�����C�fQ6���d��nH�`r�ǃr���pu ��	D�����T�^�)�����d��n#V�%E�t����#@~��;C��Jm�X�t�&�~%*��'}�h)�I�88��f
�E������QDP62X�E���!<Y�$�d�rNe[c�^�$ϔ�;&��0rV�Z~����ՆH�0؅�	�$�� �wKp\��2�τ;d/�"�B�y�H��刯D�R�;��d �IٷԚr^�SF����'u,�aS*}���F�$:D��J�'n@92#/ν����'�ޤ��"�/�j-Z@��'����G�*��bP�V"����ѻiq������{��(��ŊH�z�Ӈ�L�w���/.1��(0����M��9|���JW�]~�9cc� #)Y�}8���;��t��K13~ �
� ��M4M��x�0�!x�i�f����"|�Y�枀q�(�֪��s��9�G
i��%S���*!e���^��pL�S�B�I%R��\@�¤i�~���KT�'nX��I��6�(L��O�}�NR��ey"��fd��su/��X�����\���U�PbP�y���1q}�x
�͓:8-rał���'(pxJĂ
*�ax��5f��8�ӁN�ﲵ����>�y�!��[����@{��Ԋ��yr��X�|��w�.MgN9`�O��y��8 �Tʔ�E� ]($��y"l�=]U0����9=�bipW���y�F-0��|1�h��7�R5��P��yRi�M�����"�����Ί�?y�dЌl����|;��7�ϸfnޑ2�C�%�a{ͺpF�h���O��e
8%90���N6p[���p"O�\��_871��!PNІ@�1���DÌ"�]��E����jM�)B�K� ɐB�J5)���"O8�j'b�6X���yV @���cсҭs(p��>q�b#�gy��ް4@�� �G�dkr�Iqꝣ�y2�D�Mzt5B�@�%�� ��kK�{J0��V r�hA
�iktȪ�x/��P�#Ϲx����Io4�а�n߼t��$�(�>��U�_�"!^�Q�K_1�!򄓲=$ұ�2�\�o�Rm�����qO��x�LT�r���1��i�"(����5tPYw��'s�!�dX�%!ԩ��k�$h�`�DL׭[��-
�B�(��Z�D�|�'Y$A���ҏ޾p����#f��m)�'�ʤA��'Z��0+$'�SL�|1ň�
�a��i�3�0>y��܀�PKV�s)nx���A؞�z3���Mpx�tG|�ѥX�/�h���!7mr��ȓqP�]���b�1 Da�,M�?��âh�"B6��	N4p!�@�LOD]0%�Fz�<q�&�LV�ԑ�P�1G�\���u�<a2�D;^k���)ݺ>l�)�g�Wv�<�U���B����DZ�l���(�s�<�ǩkIz �q�Z!�ӕ�Na�<!�Ő�~�hb3d��"���2@	j�<QP!��`�49j���9B�lDZ���L�<� h �"@�!�����٫Z�hʅ"O4i �I@�]���8����"O:���	 ?~1���2D��w?ʉ`W"O$� W�7�<���7^�Je�u"O4���jЀ[Jlp�sɳ+b #�"Ob�r��	�=���K�/����t"O�%��RHu0�@�%%Ȁ�J"O���($'�1Y����^���"O��(x�p����E;!h�\��OSb�<�F�
�7�@�1n����G�<ٖ�$
���ퟙl׆(6��f�<q��T=/�bL�b�	�F�ܻ�CS^�<)G�R2�!D�)
%£a�`�<��R<#C���Ac^�v��1j�X�<�PO�!e�*S���d���b�R�<�4��-��UPtd�R`�i���N�<��kL/:L\�`�?�0��RXF�<��ǋ�{�"��%K�!w�T�1��v�<����"�^����B"�m�u�ȓ��:�� ��i��"�$ǖ��E�dt��E1�n��S+P>f%��R��-��Ȍ)A��hjP%�sFf`��$��@�đ�\��	r"�ڦFa�0��t�ܼ�S%�8�c�!���ȓ�v|B�. <�r��23�z�E|��5����Z���Xd2���H��M���>D����.�9T�B��.3��!��Njϸ��CĔ{-�B�?ئU��ӷZ��u1�m�#�DC�3kT���I�PL�qC����b%(C�	3T$�%���)���N���B�	�W>�<!Hm;�%ʝA��B��^�h� E�R�J���F�_�B�	��Jx�B���PH�N�B�əx���sM]������,+�R˓m1B�<E��-��(1̕��\�"�"Y�ڱ�?��<�S�OQ���m\�z H���M.�bܨ`��O����8,�B"|�A����s�NTNU�|�qe���%�x�aE_s>��0`ݑ��y�'��><BS�2����<8JC�2��La��?�) �øo�$ ""O8�æ;�Q7��L�:�:�"O8v�׏xꄋG��rN� A"O"��l\�zu �H׀�1�fB�IP8�L���<�Rn� x��)��#D�TGQ�X��)��+ܳ	�����N=D���-�[��@cj�3i�J����/D��KdD�0o�1�W����(�҄�.D��Hhҁ^�8�G��6<s�Ɔ9D�̙���ɪD���5It.LBBi7D�l��-] 5`to�(*�A��0D�<떫�7������}��Iza.D��SC�:�ԥ�0@F�Z+�)���(D�,��"�S~�]���+n0X�%D���wm�'`kp%8�KC��4���!D����.��b�����B�	�����*D�@:E��^캀�u%�=iL���E'D��́k�4y�\���+d�#D��;�C"H��	1�� ��q�M=D����k�Z�~Ţ"c�3D��	I��>D��A��C �U��#�7{��
@7D����mʕ)�N�b�MC8��I#�`:D��0aG� {I��+q�_1E�E�6D�������g�"I"�J�+:e3�o3D���D�Q4� ���ئ�*A�`2D��U�^�"�\���<h�)('c*D�� �H8Ə��Ib���Wg0`��%�"O�\9D�9B��8�f̅U��T*"O��c�ė�>��6�w���Ҳ"O�����7��9K�㏇c�H�S"O"ux Ă!o|h`��"ĵ$��1#"O�E�r�� g
$#T�%�DI!�"O,���0�@�
 ��M;�"O��X'ʈ)VѦ�yb�Bى�"O����KN�fj,\�qd	��:�Z"O�1��@�=+j��@d]�8k2"O�DÁn� g<��9�CU0MB
!Iw"O���b\�*l> x��L+g9rᰰ"O@�;�-��/`6,�QkC�9�@��"O�m��kZ
G�00�0��-J00�"O��Zv�͉1������]f"O"A`���4Ǹ�Ү�9�l��u"Oԇ1</��O.X��"O��2ȕh�`K��X�ڰ��"O~ �@I�Y�4	RQǹ*0FthQ"O<�������Q� 1����"O�u�We��*���H�G�5^����"O>-Z�k�<�� ��W�R�4�w"O���5��P�Hj0��'x�`�f"OLh��T Ev0�#G:1W��y�"ODћ®�C�xMx�r̹�"O�}�,�,����\X�Q1"O�-��̭i5�-*[e�B��%�P_�<���$2jb�W	
��āR�.D�8C6���Q�4�A1��1XE�(ȃ�9D�8��M[�T�$�VC�Z[��p�b8D��w(�`8�e�S�8>�AH��4D��R��Ș�ȁ�`*"
�U��G-D����nB�S|<�0�
U�3��r +*D�pP1�	`��5)6����m)P�-D���⋗G0ĺ��`�F!D����"�� �2Q!�M�|�l�C�#D�{�5�H��&��QZ&K/D�t���׍_�2�Ac���V|���+D�p�VMֹ:y�A��	PC�%q5'6D�,K �T�Z�Tq����0	�f�5D��+#G�'��)SJ�.&���4D�D(��D�>��|arI 9I1�H.D���֩w��+V�ܰ�$d`�'2D�4Y��G�[�ڼ�P��c��
&#0D�����7�&%! �m��iۖb,D�D+ ��b���@*րBB�;�i,D�!� �=~�������g�(D��P �� $�A�K��,־��B�;D�Гd䙦St�(��&L��&D� "�ʓ�!@�����%o�"�B�"D�H��� M��q��^/TG�S��?D�t�ǭ�@Ȳ����+:��}%>D��s0!�I->d�ق)���I��&D��y׍����S�� =*�� w�$D�� G�#��1�ф���K>D���u!�B���iROLp%��M<D�x�!�ϩR�橒�)�dx|��n>D��.��yRZ�@��$K� Y�f'D���T̛�Ū����>�:�0D����A���l# I��T�C�� D�
��־,K�T�	�91QB�<D�,��B��I�g�.!?��!"i8D��悀]c�ݫ��?��lI��7D�\xU(ĭO�D�+��<��w�7D�� z�ďx�!9�ǂ�x�PdA"O�P���6�R Jcg��0��a�"O�U1��ٓ��X��fY��"O^��� wN��,� @m��#t"Op�e ��5l
��+�^���"Or���H0Z[��R��Z2(��3t"O�Ms���0�jݹe� �n؜�#�"O.�����9<ExvF؎o��TH�"O�8ĩ�u��[�DM�i��� #"O�ɛ�-ˊ!�r�۪)��`1"O�bt�A�1Kڹ���ʓ%�����"O]҂�+U`�l����)��3%"Oȡ@��7b�$`s"�P[D��i6"OTI1R���T��B�|���"O���c��>��9���5�`��"On�f�[����I�
�hX@��"O�� H�-� ��6)��dB:��6"OF��`��2Hv�a#��=B��iZ"O�`#6�ߚQ�����oº:����"O�er���05��x��+9�ޝYA"OhW.�IF���-�4v%���e"O��+VJ]�_/"M���$Q�"O�XHQi��*KXQ��H
R���t"O����w��E��[)��=�"O6a�F���ZU��'C1� ���"Ov"�"�!}�e�  �$�tl�"O�x,�t+��ǂZIfT[8�!�ҏ7��#Ԭ�>A�!��ͯ<�!�܇p����iS".� ��ׅ�!�:5!b ���]�4��c�%��'$Բ��ʲX����I	�Xvl��
�'��9�+P����:M����'ҕ��C2���K"2�T���'����A�936�	���*�6,��'�|ʃ)N2��J�ɖ"rfy�'堘Y���G���g������'c��ǭŀd8aq抉��
�Z�'���;2a�a
y�5/��T�.9�
�'
p�a�L!6��{��F#��
�'�h�s�ыc1x��� ,�B��	�'(rdRE���������S�I
�'|�}8҈�-+�ڤ�'S�!��@�	�'`�
#���a��<��Dq,Q�	�'�bm����Pm���p��'),J���'P�q�fhI=�� � ]�|��'�]�'�	�V���١d���i*�'��H����)'@�i�.m��I�'%¨cP#�(6�>[(��w����'k���M6+,����ѷh�uB�'�12��ϛ2������ڤ�	�'V�q�.�af-�D����~���'-��4LZ�s-:� ǌ)�0���'{6�rqF� 0�!�D��9)� �@
�'M��R��,V��m��a�<�t�C	�'\���-O Zۄ�H4LG#
��@��'�4ʰ��^�i�3.�}H���'04X�5.�	R�nx�g�V)*׎	��'ʀ�J$
D�
n��(�`M�%�-�	�'�PR'�â[L�����ž!~�s�'�%��!�+">euMA�&"}h�'�H�ʵ�/)vؙCSw~pz�'�F4��݄,{���e�DL��'�ViqT5�6H���U�6����'�dB�-���5
!'섥���� p����+U���D^k����F"O�0G�`+dU��DZ;Z�D�b�"O<�Xd�8Mf�,�֣�v��p��"O���kL`J�|9��Qu��B"O��QЄơu���Y��`� ���"ON�����N���b&�X�~<X�"OT���I��
�����j��!!�"OE����\X�$YT��;c�6R�"O�]"��C�<uk�3:�d���"Op(;�����"1 �*F_��U��"OL���C�?#>F��bÝ�0ĭJe"O���O�(q��1��"%����"O�GN��ˬ��� 0n�v�0�"O8�*
ɍ>$���pB�^����"OJ��bA�*Ǌ�Y�.�!gѦ�8�"OL��3���D��	�Ѭ��z����"O~0G-�
Z_z�k7�'c��L��"O½p�f
�|n�&Ǌ(6����"O���� ,~�1B�%�%Kl~�"ONISc�ǌ'�\I2�T�,el�Q3"O�d���I���q�6Ώ�e����q"O�(;&�+F�L��+�r���c"O�����B%_��(�Ӓ9Z�ȣ"OTLK姕�X@l<1p�]�$Q��hB"O=ZR)�H-љ& 6ך0�B"O�E{��B<�y�% ��q9�"O��+�̗�T���oP�a1�"O��"�/#�2$�#j�<,cH�j0"O��Y�Ē�s���e	S�6���CD"O:,��-�f;8����=:*	�"OԴh�L(aӲ���fK+Y�p "O��Ҕ�7\Ř!SP�ұA:4�zu"Of�qTeY3\ވȀ5��0yΰ@+�"O��c�)WC��iJ�$Ū[����"OԄ��*�"�����#џ'�"X*�"Of��fe� �=Ec��#��p`�"O$Q@C��)=���\�)�V��t"O^��� L}�6��T�O�?���
�"O���M� Cl�c�"߭�<5�4"O��j ҫA��,���سkX�Xن"O�|yq(��"��}ȵ��?c��}��"OZT��ʘ{F�$��^��`�"O�̣э(��m�t�D�T�j\��"O�,�F�$��h2E�!V���"O�����?�P����']�`�ʗ"O�����F�a���B��@b�i
�"O }���?�Q)�I�C��!�"Of�@�"��~�6���I�F���0�"O�p�S/)8�6)9ba_�hNyJT"O�p;5j�+[� !)S`H���"Of��6&��D�qi<bE^� �"O�T�F�� +����H��Lx�"O�sB1S���0&V�%�B=I�"OF�2r	�2�V@a��Ϲ{��ದ"OB��A 
  ��   �  C  �  �  �*  _6  %B  �M  iY  'e  �p  @|  %�   �  ؗ  ۞  �  _�  ��  �  _�  ��  ��  ��  �  K�  ��  R�  ��  D�  � �  � Y �! ( 2 �8 +? <G �M \T �Z �` �c  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+q��62\���<4�d5h��'�B�'���'	�'/�'�B�'��x�.Z ?܎Yf��0d�tx��'��'���'�"�'��'���'�nY�5��B��0��g��ծ�pW�'l��'C�'���'���'���'b��i���8��}��dK�� �C�'1��'W��'�B�'���'���'?�%�����غs�9
lk��'A��'l��'B�'��' "�'O���ek�92�lu���D�+��'�"�'\�'���'��'B�'�n$Q&菷U�~�
�"��]x#�'���'��'u��'�r�'���'� �H�N$!��y;�Ã+K�f�0�'���'$��'dR�'���'���'�Fx-Q@�蒠�6/X��o
�?���?i��?Y���?Y��?���?�Po�^}��� �	\V�p�'F��?��?���?Q���?���?!���?auj+2��!� :D�|Hʗ��!�?	���?���?y��?���?���?y��ь�����/�&8CTtꖢH��?����?Y��?����6��O����O��DB(Hc���$��[��$�E/U��b���O����OX���Ov���O�!lZڟ��	�P��H���L�!�"��~�-O���<�|�iӸT���_�6HF�Z��
/��A( �C-)l�	9�M����y��'�����"қy����g2-m��Z��'9�훑u*�f���̧ca���~�6DI�o�P�YfJ�z�����ND��?�*O��}2'�X.xȝ�����\����X�jƛ��!��'���nz�]8�"D�O���3CmX1'�̻%��՟����<a�O1�i��u����9o���3B��\;�슰�"����<���':$F{�O����>��&_*�xk��Y��y�S�t$�0�4�4T�<��f�5KQ.z��N����	��A���'8��?y��y�Y�ЫIX�cHp�s`䆵]�>L�p�6?1�T�q0�j�'T�����?�ѐpI�Q�Z�$s.qR�����D�<y�S��yB@�#�B�a4�Iy�Ą �y��l�ƽP3���b�4����T!�#^��rd���k�f!z�$�yB�'�2�'߸r��i����|��O�x!*�m�E]Z����gA�4HTb�IBy�O1��'��'��ݥk�, D���-��H�銙r�ɽ�M��"�?����?N~��JGX��7h�|l��q�V!{CҠ T��2ش?1��(��i� ��B��;.��q��ѭng^��$,��[>�w���~����:3��ɓl���S$��	-Ix��P)L�9=(T�I韬�IܟD�i>��'B�6-�<>���F�H���#��,ƚ@(V"�%����ɦm�?y!R�4�ش�&�}� � J"l2`sg 3ܼ;�n8f��6.?Y󎟺�*��#���}��]	%�� ����6�� 	0F��I�������h�	ڟl�IH��eq�i�@ۺ,o�	��*B�S�A��?���q�6-1��I��MCO>�T�������4�)�x(I��-N��'L�7-�Ӧ��b�x�on~��I�@;נ�'m*:�B�MO؜�� ���P�VQ�,i۴��4�`���O$��>N���fo	4˖LQ���h�����O �����V�'�r�'@RS>���D��1���]O��q�1?�7S�(�IƦ�RL>�O`C⇒TjZ�iQCǩ}��@���-6�<	ꇠU���d��֩�O�Ġ)O�ѐ�y����e�dDIW��W�,���O��d�O��)�<�u�i��	cŇ�F�RI�%�>����	�����?Yw�i��O�D�'K����DMfu���J.�}Q1E�W`\6�즭r6�\Ӧ��'@`�o^�?U������K�)��$�sH��%��	Ϧ��'2�'3��'��'���?.�ҘieȎ���s��G�1��4,��)/O��?���O�!nz�m�珄2j2����/\�`�Hq��?۴4ɧ�'�(�4�y2�9!�1��,��V|�5���y!�9�4U�I�\��	�M�.O�	�OBaj��V�=@����́�CF�ya5F�O^�d�O*���<��i����f�'��'���:g+ƣX!H"F��G{����dU}b�f��l��ē1���Y�ala�&V�@�������Q~�o��p�`�@�-��D�ںc6��Oxi�@[����㗬�D�l[U�py����?����?����h��^����1�x�ؐD��t������M�G��ϟ��	��M��w�n���;#�]�����DQ�'�6m���Q`ݴm�(�ݴ��$�zJ��'V�x5�F�%_�pW�K�a���1S��<�ҹi^�i>���Ɵ�I䟀�I�j���C���i���"�Ȗ�rTT�'�.7�M�e�r��O���1�9OT�a�.v��($DA�[������D}r�q��l�=��S�'m��|ad�Y5͠�!�ɒ�ZH�"�冤u��%�'�$�*�I̟4K�Q���ش��DD�E������@��l���N�8�8�$�O��d�O��4���<_����	w b�?�^�p�Q�������8�y$u���{�O��o��MKղi��}B�*�'�^P�`��cҬQ��ƛ1O�����L�#(�k�ղCN�OcP�=� d!�%Ȋ��2�� ��N�l@��?O��$�O`���O���OH����Ӊh�Xh@֊�i�QȐ��~���D�O���Ԧ�#�*�ݟ���ܟ�'���"*P1H%����(_0,p5H��K��M#.Oj�mZ3�M�'�@�ܴ����Z�`ٳ�ϙ3Z��G��y�j��qER=�?i���O���M�����'"�'��I�wa!C�f|��X+W�^����'vRX��Z�42Q�����?�������\e� �LM�I�Ҡ1��������?A�O��$l�Z8oZB�'Bq����H�lRs�� ؘa���v�8�W��a~��a�=���'o��Iğ杘}8� ���A�>�@�bЯ^�+��q�	���$�i>IQ-^A	�4�'Q~7͖;h6�q�ƨE�c�phUF�41tc�<�����?�(O�9mZ|�jT[��88r��4�Xyp8���4mɛ(ġzě���|K�-U�9>���~�qi�7H�%�A�ީr4*P(��K"��Y�����4���,����d�O`X�X%�,Yz�vO�,`�ĩ6m�����>_(���O��i��'M4˓�?ͻ:��dcF� �PX���x�+��iAj6��Ȧ)���O�x#��i���k���vm�4���	4��O��č0b�q�LSJʓ1Û�P���ޟj��O/R�L�C'�*`r6�xT	���Iϟ��	AyR|�L�o�O�d�O:��"
�0��5�ti�40T.�O�ʓ�?	�P�D��4Tϛf�rӀ�z0���paA;Br�\
 .	8@R��'���Ta[,
����Oͭ��n�$���?�0%Qg	x4�Sj�^y~Рw�N��?���?����?��	��\�ɹ�ztIc,�/X�0 �aE�b��ɘ�M3Ca_�?����?q����4��/U�`@փ�	~�i ��\���Ʀ1*ٴC؛�
մM������v!�<��t���Y�B(��wa6K�BR:�0�A��� �	��M++O�I�OP���O���O��)\���@I���TdC��<q��iA2���B�b�'����p;��'��M�%^�
�S���	=.9�g�RH�U��vHr�Rhm��H�B��l^O�Lhx��ͽUl.�&,�+ ^8u8���|PSmؼV�)�Iy"am��� kj@2�B�;f �\���ƨJ�d����?���?��|�/O>t�I2p���=^̱���H�U��rB�}�Ĉ�!�?��Z���I����4Q��BD Iz<��TiUjF���l�?�MK�O�m��P���J?e�Xw�IGp�x�FI�&*nxӢ�C��yr�'�2�'���'���Ӆ6Wؑѧ���MF��;�O�cP��d�O��릙��)�qyB�o��O���R���Vƪ���"�~�p�X�i�I�MÕ����眒N��&3OF� ��H)'Ģ(Q����Zl~�)���S�,���IZ��P���.}��Ryr�'R�'jb@Q�w�
�;��^�z'z�`���i%2�'[���M�6 ��<���?)(� ��vF6���G�0}iVH�7����+O ��e�v`'��'Kly�G�B�"��C����,�ʰD�k�(L�"��~�O��q��<~�'a�-³"�l	��C�ҹ\���$�'��'�R���O���Ms�āY ����9Q�*�:�L%�ƌ�'7M0��*���S�Ar ��"2�å���`�!
5b��M��i芁�Q�i���v0u�%�O��'#� AQ .e�\(P�mYmB�͓��d�O��d�O���O���|2��Ʒu\�$�5h�?0G�Ź񧜜j�����y"�'>"���'��6=�"Xq�W�$'�!S�]�_�U�D&J���͒O1����!q���I�s0���ą�Π�2+�:1N��ɿ�H���'�¬'�蔧���'�2������r�\0��4���'�R�'�"]�d�޴X+Y����?����5h�a˭b|`9��ƻ�C��<���?�M<)ck�?<x,�'�^ 8��:���k~RN�p���&c[0Y-�Oj���I5Yd"	2m 4��Bk@��d�#�i�K�"�'�r�'���(
7�M;z���s�[�6U��JQ��\�ݴL�$����?�q�i��O�N��3%Ba�Ei${�E�Ȉ^~�$������M��m�M��O�I����S���QŐ���ԕOp�ac���C�z�O���?	���?����?��Rqa��P�*�1���H2�),O&�o����T�����j�s�Q�	�=}�p�R��pk�����N=����Ԧ�*���ŞK�\+BMïzm�Xfo��U�������-O�u�P��?�0�>���<AF�Ϩu��7�<q�|9��j��?!���?Q��?�'��$���	ccm��dƇՐu80���;UlX��럐�4��'Jʓ�?1���M���W?N82.R��2�(p�	�#ڀհ�4��d�!_,������������� c���%Ɂh��,	�Ɓ�'��'��''��'h�P���Qd�(8�!t�a�R��O���O� o�u���|.�� ��4��$��hN�u°�й+��O\o�
�?�(��lZs~b.�� 7^8XsIA"�Ju�e�՘~��"Ɵ�!b�|�R�\���T�	̟p�`��^ٞq2��W4_���x��ޟ��Ioy�`y�\`�B��Op�D�Oz�'`�z����)+����ذ\���'�Z�l�*�O$O����`<I��ц{�$x���h��8G��<)���G
�7z�z������O�U�K>�c2#�JG`�7Rp� .���?!���?���?�|:)O�Hn�?af�	1���_خ$��C�!H���vCV[y�F~�
�d��Oao�m�h�
�D�x�n�1�
�J�.$�޴�?q!�_��Mc�'�"*D�}��y�-��� �I�ƿE4�ݪ��*cB�!0Obʓ�?a��?����?Q�����-��\�sH�'���7%����oڢz*��'a��)�¦睙V�$릆_V3"����F����{�4"ߛf�'��)�әY�Dm��<)@ON~�N�%A�D�{���<ɧ(֭@X�dW?����4����җH��M�#�I(t�VE0o�%;���D�O���O�˓\����/f�"�'��@g%��"�؆W�:��fO�V�?	�S��ڴ=����' ��*_Jt������"SBߴy���-(N��@o�#W����|�q��O��S��?�J�C���qH ��%��¶T����?q���?9��h���dZ��~�������� vI.���@�qړ%VSy2�m���]�YO�y�7��~z
q�'O�	����M�ǿiJ�OG��v��<q����de�\�FI��g�����ae��]F�T&�������'���'Z��'L�0jpjўVf�-�Y�Ԛ���ݦ�S�J؟����%?�ɬV'.ْ�Ә���4�[vd�X�O�l��Ms���>���,�N�Z(8�C��P�T,�¡\.MZ��d/&?q�E�O�*��]������F�
|Ke�#n#�l��L�v� ���O���O��4�,ʓ!��)��y2�E#��uhZ� �5
��y�i~�㟨��O��m��M�Ӳi>ΐ�����"_d �'T$m����	xț���h�� �3,���i��^�����t��K�톰^�Z���>O����O��d�O��d�Oj�?9)"lY�N4�M],&H,�W}��	�BشJj���'}�6M0�ā<\��D8`@��w�4��59�
�'�h�4՛�OX����i��Iy���'���v��䇙�f�-b�Qq���{�	Ey�O'��'�Nޑc���</94��ҡ9���'9���M;�G�q~�')�S�>s��9��N�Cpj�+E�U�c���t��I��M��iqLO��#O��I��
�P��SF�ԋ];�p0��(;����#?ͧGwV��ԇ��>��ñ���)G�yЂ�҉O�"�H��?1���?Y�S�'����?Miڈu����F��8��r��
�˓d����$�l}�Ns�j@z+�r�9r�L�dߞ�֥�䟸lZ8eܘ�l�p~R�E&9��ӱo��	n�#BJ@�|} `�[ -���py��'�R�'���'("[>A#g�S�L+���|ɤ�'!��M��&K��?���?YJ~�'盞w������:d*�jV;^�� �{�����e�)擉G��m�<����h���!*�Z�&��ˇ�<���̀�L���+�䓔�d�O��d1(�b��1B"���I�?�2���O��D�Oʓ["��C�V��'�bF_9 ���K��L��X��Сx`�O~�'-�7͍� %�pz��Ead��Bϫ$)*���8?2F�\�� �	�6��Q���䏶�?)��2U�� ⭝�|Ip���Ջ�?���?Q���?�����O�4�&��+[�%S4�Պ2r$ԃ�!�O��oچ҄���ğh[�4���y�Β�:�Nh� ҆ڤ|c�Ō+�y��dӄL�	Ԧٸca�ڦ��'ޠ\aSdL�?u��*���и���	���aD#i��'��I����	ޟt��ܟH�ii���?�v9�נ�6]~����<A��ie����')r�'��O+b�'q�,q!1��}�Z�0)��-6b�	�v��O�O1����m!a��*��<&>p�2�	~@j6Ϲ<����+m��Dؼ�����٣s~���C��W�|؉�n¾(���$�O��D�O��4��ʓ2��*Fd�2�i�p��L�#uRl)�#��y"�wӐ��­O��n��?��4w<@��:��XS ��B���P"�M�Mc�O��⅜�:�'����T��6F��������d��0O��D�O`���Ox���O��?�@�G�#F� J�{QыS؟L�Iϟp�ݴN��u�O�7m#�D�PDn�#@�;{( ��G�`6t%���4T��O��0���ig��-!;��؆h��O;T��A����D(`�@l�CK�IIy�O���'	d�xov,��f����k��K2�'"剣�MK���?	���?�-�z�s�C�+\�!�,�~خ�U���q�O.nZ��?�L<ͧ�J�2=��3%*���BT&��\� "��06Q�Ѳ-Of�i��?�F�?��U�+V	 !@�c��+@��]S
���OT��OH���<��irjB�$�h4h���B"���A!I ���'��7�$�	���i�.D�3��'l��"&'̬lv�z�aŦ�ܴl�Q�4�yr�'�81c#���?5��[�S%�V#T��%�
�DM�P�Ghc�d�'q��'�B�'���'Y�,�@q�� LLq ���X��c�,ţaD�O����O��ɶ|Γ�?�;.gH�	������6�K�p�z��0�i��$�>	��|�����S럹�M��'q� ��˷�P�Y�ł�j���'M��(�͕ڟx�v�|�]�X��֟�� &�I��t�ȼK�j!n�����Iß`��tyb�z�ZP��O����Od���hͼ��IR���"t����&��2��d���e�����-�Z���K�~}<� � �w����?i��͌�\C���d��n�C��>��Dmc�4ڣO�!t���E���@�$�O����O��d+ڧ�?��JU$OT��X1�ȘY&,a���?y�i�,	s�'mB�u�Z����d<��*ñ(`��0.�!UVf�Iަ5�ڴ�6�Mʛ�2O��$��	�0���L2�  ���Q)C��P"�����J)�D�<Y���?Q���?���?��DÙzАPcR:F 楫�+���$Wݦq+f]ܟ�����8&?���.rkd���Bр3�l�B4-��sb�(�O��m���?!O<ͧ�b�'4!
-	Pf�scr��6I^>^D��㨏Ge~�q-Ot����?Y��<���<�R���sބ;gJ��_1�	�pi���?����?I��?�'��DSݦ!�be��<q&m��S�)%%J�k�~�kW�z�4�ٴ��'�j�rԛ���O�7ԗ�x�€ͣ-?H��b� a��g�eӨ������"C��,;��YIyr�O�G ܶ@��������Y8�fO��yR�'�2�'{��'�R�)-0zx)��ʬW! 噃iQ-)�Z���O���VϦ]�sas>��ɹ�M�M>��ǓK����2O\�A�bߩ|��'�6mX˦)��i�.o�<A����=��
�}ڨ:AhϺ>(��Q���+@���H!������O��$�O �DЩ�"t(��{mtزF��E�r�D�O��n��̄@��'1B^>� �R�P]^QL'i�XԐ'�$?!�]�T�ߴcf��l4�?m0�
�I�Zh�v�	6X�xa��s2 ,� E
l}���|�T��O�HIH>�,њ`��k �^�7$�Ay�'Ɂ�?Y���?	���?�|�+O�,n��C���#D/۫v���`A�/M��1�Ϟy��c�n㟬ɨOlZUl$���G�
2-Z|�Rh��uΕ@ݴכ�k<$̛v����N��3*���~z��S�Z��]����2�v	���<�-O����Of�D�O��$�O�ʧ��ko�t!��<K�%3��i�~����'��'2�Obb|��n 9���7��<K�9�)��J�ƕo��Mkx��T�SAU�8O*1�S�[@i"w!Nx�*7O��ؐf���?��g*��<�'�?���ɣA�Va�5�F@�� �?���?������Ҧ����_yr�'W��$��A�~���`+=�89�����f}"�aӲ�l��ē����"�A�]� �,��T9J��'&��r��_<r�`����џ�`��'���Y��,0�&t�V�VPƤ��7�'��'���'��>����gl�$X1�H�g��1���cƥ�	��M+���:�?	�)ɛ��4�F�R�H�A�@�<_��s�3O��lZ>�?9�4Lf��ٴ����D_����'?�<���Ʊk`�rgG�N��ru�*�ĩ<����?!���?����?Q����C��!&y�O
��d�Ʀ�"g���t��ß<'?�I�p��i�[L�$�!��rK�u�O��nZ��?1O<ͧ����I���ւLZ���#� >m� +b�$�@]�.O��Q�엉�?�u3�d�<9r�Kh���'#��g���JgCK��?9��?y��?�'���Y����П�D���zD�a�¤�7��V#����ߴ��'����?���M���u�XKgKB�P�t���`F�,�۴�yR�'/,�b��?�
Z������E�F�еPZ���R�Z��Q�ѭ~�X�	ğ(����	����J��'K����0m�<&�h��
��?���?�ôi�I��O��z���O&��U���$�H�*��E[.���n�k��;�M�g�i%�+�^��f<O~��B+#Eƕ1��]0TBmP]ufy�b.��?qE!*���<����?)���?`jO�#b|�J��9��y�3�?�����S���Wߟ|�Iޟ��ON��Wj�
�@����������O��'o�7�U���$��'g��qd��/w���G��%K�@ց�U v�N���4�b@���0��O�$��L��" :�*A(��\$��O����Of���O1�.�9M�)]�%�Ri�u损|�R|�#胺z���R��'e��e�㟨J�O
�m�$3��A�NǖB�=�2�`��YPڴ0���LУu�Ɩ��Q4G�C ���~B�AֆQ��xS��k�˒��<���?����?���?����?1�⚐3��N#�,� �@B+ir\���-՚t�y�����?���?��i��'�2^��N�K?�K�CM�Z3<\1��H�?��426�U"��Y��y*���d�-S��7mk� ��k�q#ݨԩD�J{�a|��W�PK�"��@�	Ey�OG�dܯ)�:ap�$9 ��ji��'k��'*�I��M;����<I��?��lť"�HK�ܞO��bT	���'<��BǛ�Hh�x8%�����,��x��@�02�H�?<�'m�B�5�JT��,�7��埲���h�
��Φ@��8
�zP.lA��Y-Ӣ��O����O���*ڧ�?Y�ẺeJ���͝�(r�Ip�,�?��iw���&�'��k����]
^q�I��@�0�d�2/�J"��ğ�m��M�d��MK�O�A� �%��SMU%\	��+�7�:��*^UWV�O<��|B���?���?a�I�*Պ ̅�3�b��Ǭޥ{=|=�-O��n�&�,��I�h�	X�s���yp�(Ku��d��P������D��aY�4np���O�Ji�'�L�`Q�5�*>΄� �#+ ��*�O�	CE����?AU(;��<�SF�5�0�!)�'�j(Au�;�?I��?A��?�'��d��ө�ޟp�ZV�lk��lұ�cC6�<��^����?9�]��pٴmۛfAj�pɡ�ÖC�^|��&2�M!��
Y�~7|�X�	�	�d��3�O������;:N&h����*��� ��C=9�DUΓ�?����?����?�����O�
812�N�G��y!��H��O����I`d,?	�i!�'�̭�d挺DdH{X{3dPK������,��Fm��)X�k�7m"?�d�g�? �������<� � �@��v��;��?��- �$�<�'�?����?�%�+#Z���򂀾E��0��͜ �?a�����!���ڟ�	��t�OT�����Z�d�p��ϟ1W�T@�O���'��6�Z�%��R�����d\�9�b,;F������.W����ĵ��4��D����̓O�d�'D؉��!sN���U&�O��d�O����O1��ʓÛ�Ǆ�-ޔ ��B�]�fRbG#���Ң�'(2�v���L��O�o�:|x����i�3)��t1*C�En(���M����M+�OpX@������<!��׎mEl��!6g������<�.O��D�O~���O����O��')�H!�.�
�y)`	
�xn&s�i�R�QA�'��'Y�Om��'-V%2���aO�帠ϟ�N���o�"�?9H<�|:�!?�MS�'H���F'׺@Ä�W�v@ !��'m����l��k��|�\� �	˟ ��ፊ}".�9S!�n\�(H�F�֟�	؟���Ey�wӀ���G�O&��OR���ND�F�.5��� "x�#�%�I(��DP��H��ē�&i��h�TȊ�JS�e����'��� 5M��oȹѳ��������#�'���1O	h�T��牌�S;�j��'���'��'��>��r\��Qb�5�ι@B�Қ7yB����M����9�?Q�&㛆�4�vU��E�b�dę׃:,�r:O4=m��?Y�4Ns�4�ش��D�:,����w]p��a��WD�|�"�-���S/.���<���?A��?����?ys��>:!�[G�8)vb���O�6��_ͦ	�E�My��'��O^2B�)Oxpn�bd�� "b�h�h�#��F�O`O1�t���k���uz�/�>R^2�ܮ`!�����<I�J~����:����d2h�t�P���#m�b��������O����O��4���#w��А'��^�^:����!8{������ry�jcӰ�p�Ovho���?��44���"c[�[��	�����$;&@��M+�OX�˗��$�z��?����
*�e�B��.�5av��V;O����O����On���O&�?��b��z��h���sG��ٟ@��ɟd�۴l+"��'�?ᴶi[�'H|{p!��1�pj�H�$�9+��!���O���O��Ԋ�i���/���͘==�X<���Q�hTr(�߼�����䓙���O>�$�O���r�+.�e�1���e��ǟ��I~yr#i��
E��O���Oʧi��8@��'��i1.��T�d�'��d�6k�OO�S"e�މR1m�4t9���r���m�n<R�] ���AׂX}y�O��Ib��'�B@����"�٢��~���v�'R�'�����O��ɼ�M@FXOA���$�R=$�nU���Y<u���,O�oZD��!�����MKe��5��P��\5C�JM��o�Rb�i�2d ײiO�IK���%�O��|�'�ީaOS�X�|����U�&��K�'���8�I�`�����Ic����rX$9DI�B $���T#�6��+�.���O�d"���Or�mzޅ�B��/@�|Q��Қ^n� �N �M�յiW�O1��,K�Cp���IZ2����K��48tL�<Z��.>D���p�'ʹ�'�������'�2	�3n��M���LR�if�'\"�'lbV��!�4qL��z��?i��r�}�rhU�r�����oڃ	��`�2
�<!��M˱�x�%H\�b!O��w� c�ֽ��䞤2-�p;deK�~#1��|��{#��$ǸP�v��ƕ4^�4��A�žN�(�d�O�D�O �$"ڧ�?)4�>j3@Qb7%\\(ma��?w�i������'#R�l����'X<x� ����w�h�0*�H4Z�I��M��i� 6�W�`6$?�G�h�f��	�ѩ�B�
�+��٩%���I>1)O�i�Od��O���O�P����;OO�r�ܪ
��A�	�<ҾiHĸ���O���.�9OZ����Խ>I�5���Ӱk*�Б���X}R�y��o���|"����Ƥ� Lv����2Ԓ���T�n���a!V[~�]��y�ɮ6"�'���R�nlI���f�:ADGB�_��H�	ş$�I��i>�':�7�hf����%y��g�N��a󪚀h�������i�?9�_�h2ڴJB�i*�`�j˖ Wb�1(մM3�	tK��b�֑��`�(��	5��$�G��߁�c�'%��0��u4aC�ko�|����������I�T�����+�,,�����:bHQ�`g��?����?qb�i�dY�˟�8l�џ��'��I� ϕ�b$���B�A��ъ �8�dĦ9ߴ�����MK�'#Bʘ?��h������
�8� 8�P�Jϟ8z�|R�|����Ο���GN= m`G�[d�C��<��Syb�dӴ��1g�<����i��S����eP�5���8.@�Ɍ�������������|���?��(�4�$�a�ʷx��qa�-P	4ƶ�Ѧ�����D�� k�	?D�O�)�0�U�?������Y5Uh�H!q�O��$�O���O1���a�V��>W����e�\�9C���Fm��z%�'YR'pӚ�;�OZohن�YuI�]��@M�n�1��4%��6�'n��f?O�D�3J�����b��w����� �:0O6�1V�ٴ�r�ϓ����O|���O��d�O����|��2DJ⬒��ښ7�dJ��6A���U��'bR���'�r7=�8	�bO�9r�$LD�w\�<�p�[�	*����|��'�JQ���M۞�� �Y[tfT�CɈh5인Y����;OJ��l7�?9�*2�D�<���?�D�^4%�Q�e+K2t:��H(�?���?!����d���I�f���X��� � ��D%:'��H�)���`�2�	+�MKS�i�S���B��99=��0(�G;�Yi��p�x���𨳐Cи%2�bV��Oxdj�L���BWƎ&�t\㥍C�=������?����?���h�>�$U7{��80 �ZbĜȠ�K44�@�ČҦ%���8?ɰ�in�O�.
�4I8�AvA�.����*^�?�ܦ�!�4;e��-J-%�V5O���I+�����'3I�h�C޶sp��)A W�u���ʷ*���<�'�?����?����?	P/IY�!���@$���[4C����$Dߦ���c|�`���X$?�	���J�ٸ|V�au''1�3��D�O^7��X�韼�	���-S��)p(���Ɯ6���͜oؾ��P��d��&�9��FN�IQyre��G9
̃4��halLq7�WlR�'T��'��O�I�M#F�ƫ�?7%�g��`3��]�wʂ�@��?��i�O���'��7m���Dm�^V���Q�D@s��őp����	
9t�7�%?��%���I��ҘϿ��-�i�m����Us�BV
��<����?���?Y��?)�����[1vAٲ�@y�fԈƥ��$HB�'��n� R�4�l�dM���&�t�T�����"G����u���A'��!��O�O��k�0^�f��d���֘5#�$9PNL0�zEp��� G���q��'�� &��'���'4b�'�(\�A∂8���,g����'�P�Tbܴ2ޞ��(O�ĵ|��$�E��}z�
A��N�8i�~�!�>90�iښ�3�?�"`N�y�TlP�9����(n�tx���H�>喧�t@I����|bn�{`dS�NL�7�rh)!�W�c���'�R�'c��4]�T�ߴl�$�����>DTh(@7e�:�|��taʪ��dJզ��?7U����4)d���+��0ًCJʳ*ઉ�U�i�x7�_�U7m:?��K���>�	+�Ԡ����Q��t��udX��y�]����֟������I����O�P8���U�Z[ވi��[��C�mӬ��G�O��$�O�����DH���݃@N6p�pE@�W����e���$���4>���5��	ɓ}��7�s� �S$n�XmHB.�7�6I�p�P�ƁU %��i�D�@y�O/X�)����O ?F>�x4o�1<�R�'���'�剩�Mk2���?a���?���� ��Y��\o>�Ec��H���'��� ���gӬ�$�؁�/��Y��H[q�<E0@It� ���l(hK+�|������O(���D��3w,V?6����/[�BՒ���?����?a���h��ė&%w�M��<t_�RV�[�C�\�d���=���KUy�sӌ��]�ecέXcK��W~p11�@�a�b���M��iS2Q8~�����X1Q��0`���眠a�J]�ri�2�>@����5WuF&�P����'52�'�R�'�Q�4��t쀰u���q[؉X]���ٴ�f�����?�����'�?�D��
|��+Rk��Y���C��"�I��M���'����O�� �e*�l@�e�i࢜HfKZ6��B�_���r-�*j�
l�	jyb*CV{��kU�×[���T�X�y�����\��̟�[yBxӞ9� O�OjP6L܏���8 ��er��>O��l�S��t?�	�M���'�L�=_p�;F�Ĺr"A�1G�	l��0!�i�����e{U�O�&?	���K85�F�L	[ڎ��@�=��	ß�������Iʟl���Oc�\;�mI�$f�I��J%W�0��s�'���'� 6�xp��kț��|�b��۪lb�O�!vP����*2+O,�l�*�?��7���n�W~�b��a�R	�CKZ�!ĩ��PRTq�G�ӟt0$�|�W��	��	؟�3��՜`=`����0qS�I����Ify�Ge��0����O4�$�O��'J(�X
�V:�L�!�3k�u�'��Si�FE�O�O�S�C��T�탚wq�yQ�ǂ�rw"�8����z�ǘEy�Ok>��Ic_�'�|(V`�q�V�%��0
!n��'��',b�O:�0�M�瀋�Tb��U*"�(9�p��7��P��?���i�O�p�'��7m���Qk״o�B��f�<���O�7���6M#?�2/U-Q֠�隁���x�ɻ% �@�N��`�<f8�D�<1��?��?���?A/����I��bܩ)d(طG���!]��D�C���	՟l'?�ɻ�MϻV�x�Ԃ�'��H�!oT�R�d�h��i�^6��|�)�l��m��<I�h�
\C@�^��&)��<Iq��5	��$��䓈�4�����L8Lx8E Y1,�Ęh�T�/K����O��D�Ov˓Z�F�H�zA��'Cǂ�i��p6��,s�h��$b��s�O$U�'��6m�ۦ1�M<��̥k�܄p`��Dd�DOZA~� .zE�}�t����O_�a���1�Nų\�]���i�x��[����'��'�2����J�n��L�p	9���43�`�Q�^��4ufr�.O<nZK�Ӽ��T���*���+c� ���<A6�i��6͙����&�DĦu�'ˤAB�A�?�
b�K#��y[����R� P� $� 1�'��i>�����T�	ן���;�vQ��$E	jpH���� >��ȗ' 7�G�V]�d�O>��$�9O���⥖�aD0p�B��it��`��[}"�aӴlm����S�'O�L�� <i�5H����|+%@Y�<�ZH
�)�Y��ɳ ��݈d�'�>�%�Д'p*@;��({>j�H�՚8BE$�'A�'�b���U�|K�4}  ��8,��@g��a��I�!��:~��͓)0���d�M}�ijӪ�m�M�%���+�(�0��ݸSJ1���k޴��DN�P\P���øO�wNqe�X+F)�Ir� ��a��yB�'�R�'0�'O2�IͬW��$�6e��:h�NZ!Y`���O����Yr/l>e��6�MsI>��DY� �!��G��ZE�\�{H�'�r7m��I�	;Z7-3?��DʄLR��w���I��'��� ���O0�J>(O����O����O�}�V�X7d��l�r�Z .Ŭ�2s��O���<)��i۴D"��'D��'���U/ݜu���хL�M�a��I=�M��'�������0Q�a�cA�O�B������D	�E��(%�5[d)�<�'x����%��Kt�����=NZ�l�H�r������?���?��Ş���֦�pDС&iQ6Ĝ�tTb���훲b�'�7�=�I���DE�EA2쏕�`y�3&��\�6�Se�=�M��ir刖�i��$�O�h����ڴI�<�Vl��]�B��&��3E�iZ����<�-O���O����O����Of�'&W��X%� ������X�h��3�i/.dKB�'���'M�O�@u��΋�'|��t.U�n��a#����,�|�l��?�H<�'���'H��H��4�y"f��Hs��@H�w����f��yRG������k%�'��	ɟ8���/xv ��J�=L��@�Y*]���	ٟ`��ş̖'Wv6����&�D�OP���1t!x��������P$`�>����O4,l��?�O<q�FK)[���h0J�2v?t���D��<���4)� Z�9NL�3/Op�)��?�q��O���s� �Q*Ď3e��;�Oz���O8��Oꓟ�ä	U���ښg��Pb�]�k&�R�o�)^ˈ���uDMğ����	gy��y��Z�q��K���4Z�
�
�*��y���^�n���)�ܦ��'�
��H��?�"ލ"�t(�7+Z��Ha����.a!�'��i>��័�������"'�ܱz@NM*LaN(ТJ+^�@�'��7���:TR���ON��5���O,\��\4z�D�3�^�&S��T�Tty"�'|J~�`�A�M���%�;\@1������ݣB+����d�3;����O�˓d ����:g��TI����d�VLY��?����?���|�,O0�o�32s����6|؀��g\�C�5�ca �Xǆl��6�M��F�>i��i�d�D�v�s�g�e���P+�+ڐ��ь�ze�7�2?a�BW3Q������ܿ���WD��Ř���.p�ȓ`�N�<I���?���?1���?!���@��p����0�K	[Q2ؓ"�,R�'�B�k���@�5�H�d֦�%����d�8P��ӿHy�q�5��ē���k�O��d"E����w(h�̌`6�(hEN��sg��f쪶�'� �'��'���'K��'�H��f��x�T��3�W�
}q�'�B]��
�46�nm���?A����Q�D��pb�� ��i�#��I�����������S�dj�)7�p̉��Ƿ3װa�R�A�`���pc�R0N|@��Y��S#H>�m�u�	���F4]v�(���]K~��I՟L������)�sy2-m���)��ÿD�Ix�� 8�uW��>�2�^���x}B�u�����:��E����F-`�S���ܟPm5K��oZL~2�
�KĨA�Ӡx�ɟ����S&X��Z1BŘ[X��	`y2�'}��'���'�"U> 2
ڴN���k̆692��E��M;F![�<����?)H~�9t��w�0�+��`�M�b,��<��mc�2�n���S�'D�ta(�4�y�_3�T`��KT܅Cp#��yb�K�&ZQ��;6�'�i>��	`�`�x�d��6�X#
޴+٨�����Iß��'9�7-�-]����O��䑗Q���A�ml�ja�ԍo'�P��O�m���M��xb��M0N�"eѡ/��1i�Չ�y"�'eM��8kZ���O���?�?9���O(����
�o|�Q��R�e�l32h�O<�$�O���O��}���+t�}�@�2s8th�d]�� ��#�> r�'��6$�iލ�$� D�Ȁ[���L�P
e�r��P�4@ɛ�os���P0�vӺ�	�$�$�&Q��$�Pv��A�?46����R'��%� �����'���'�R�'� �+f�m���h���BX`�!]���ݴ(z����?i����'�?i4[=T���:��%7����-����ɹ�Ms%�'߉����O���X��pi1*ȣ5�ɹ���8:$���B�	��剳"��0V�'\b�&��'�"�pR����7�.����'qR�'������V���޴%O�;�bך��VJ�&�҅�`�Y$��3��7��v��[i}bCh�&��	��MS�F}���{!m��0�lEb��ɢ1l|�n�x~r�Y&�X��ӻ��O�+�d"��ցBa՛#�^�fL��Ot��O����O�� ���d<�7̒M"nY0�f�P�� ��	�M�`���|J��}��V�|���@��a:W�ǗK�����M��O�l��?�SO�v1l�b~ҋ�=@@0�"�ͽ~i�T�����'>d���蟌��|�U����ʟ���ޟHx��_�j�2,,��2��ɣ���ß`�	dyr�^��Џ�O,�$�O��'i۾�B�C�2��$�@ܯ#���'Ք�l'�&��OzO�3� 2��!Ĵn����\;5����㓊W��A�C/;�P��|�s$�O� O>��j��%�r��.۱S���R'g���?���?����?�|:,OԤoZ�$��*�Z|>�i�nݱn�D���HßD�I�&�#�R��>�u�ih�p�3ǜ"�ly��m��$m��O�7��>g�6'#?�SN�k���C������D�k~�b�[�m��$�<q��?���?I���?�,���*<+pb]�@f�_,�<P�Gɦ�s!�쟼�Iџ$?�����M�;4��8ɇ�̫\x�h	�lށ�N�Av�iYT7-�^�)��\���oZ�<qρ����҄�:5s^�l��<Q��X�/Nf��T��䓭�4�6���.B�li�#ض<��+1��8�~���O��D�O,�?����q��	�Z/�E:6�
�i"�Є��`��[��	
�M� �'G�' ��h�L�:F�*D�&#�$7:j���O�U���8M�ո-�I�?$�On�
[v��F�D
h��I��S>B���'���'�B�s�a�qB�y��8�h��D@ -<�ݴi�)s,OP�lZB�Ӽ�g֊*��TY��۱@L�庇�<�f�i��7��O��	�o�n�EL�᪶��T���/߼�i2N�� �bЁֆ����4��$�O$��O��$��fyi�����6?6%At^�vp�N�6��7;���'����'�R���U*B�
-�Ә9���>�v�i�<7M�O��F�t T�=w��X�K�{��E��9Q$�Ä*؉��$
&fr�D��w>�O����$R�S�9X��V(C=o�����?����?���|b)O�o�f����	1`J
�tŔ����0�R�a.批�M��b��<���M[�Tc�<af�]�X@ʭ�gJ�"�l�/��M�O��@�����w�X��eHBl`иJ�E�,�2�'���'��'���'%����n�����f�=.��x���O�D�OBplڌC���':V7$�$V�\�ED
� ��բ��k�|��<��i��7=�ȹy�`h�*�Zi\8��L�0�0�Ҫ� �JIh�!��(ɸ�$�1����4�0��O��
5*
}ɕB�("u���ǏÐ@�j�$�O�ʓǊ�?9��?�(�H|s���[7��R"r�ȤJb�����O��n��M��4����0S$�*zO�2t�Dh����e:D��z ��O[�i>)���'���$���Sl�}`��r�iʲ'TXP����㟰�	埰��ğb>��'�~6�_	o��q��۠n%���`��>(R�Ʃ<�ǳi��O���'o7�V"#��,q�)�;	���-�,�Gq������B~6-#?��ۦ1��	%���)`�t�3�K���r�*�y�\���џ����� ��ȟДO�� ���=H��Ē�o�7�
) �gӀ�)�O��$�O���$��睥=�h�̀<�Xa��m��� ���4?���'�)擰d��m�<��H�:����mA,'��s�kY�<��Cۯ��������4����_��ʇ,�X� � v��S6D�$�O����O��=��VIƹK��@I@$��@��3a͂�8E&�h��VU��C�����lZǟ�'�P��йv��5j�h޹�LS�O e�����+��Qf�G��?�f��O(�1�a�0,�t|��̢a`�B���O,�d�Oj�$�O��}���L!hA� U"iWܵ��AI=q:��I�^I2���$�ɦ��?�;4H��0�F�k�Vѩ���ʰ��O���pӴ��KY�7M&?�i�;y� �)�^ ���d�؄R��aw"�!K�p�M>i/O�I�O��D�O��d�O\A��a�9���V�U0_z�}�W�<�ҿiOƠ�3_�,��X��
�h�pl��4̸M���`�T���P�4��ߦ=��m~J~*A�;�^�9��\����07K�(�t]��ˆ_~2n�0s<���?��'r剅��R�!Y l�^�J!;��%����d�	���i>��'��6���{�(�D��){���	�{��Y��D]7!���ۦ%�?�V�\��4ܛV�'�\�jT�2
��薭 ]���RG�{�����`��#�V���9�p��lI�R��E#P�2D����3O��$�O����O��D�OP�?��'�Y!^�r4x`��hq����Iǟ� �4�x@-Oz%l�I�R?�1�F
 -�nmBG+��Icy�G}Ә(lz>1��LA����'OH� ��th3���:e^��KՎ�	��x��0s��'��i>��ퟔ�	�8�YOK�=*R䀠�U
���IڟЕ'�6�!7����OR���|���7I`,v�*����C�w~'�>���iV�7��O��~���!34P�����ą��N���l����;��������';��2�gۥ
"XH�T��M�'�Y�w��ZQLӋy
�}"'.�g���ئثш�ye�1^�>��TL�E��[��|Rn��|
���̅धB���O�J��HQLhpc�ҝ�J�KǄĸXBޤ)@ə/�A06!\��}k�gK��ĉ��ci�H`"��߲Ljn���̒Hn�q�

;h�&��g`D ?�:�����6}T�q(���1�^��,�E�ݳ���(� �#nW*+���)�I�!RC�9�GA���QCA��5l�� 4�O�@Y��:D�7Z$��ZC��>�*OJ��0���OH����^�>-��Z� ;d��W#8XÀ�3���O\��O�ʓg֬��W=��tKw�{ �S�@O�Zഅ�D�i����X&�\�����TCQg?�!M4vhT	��F�$sQB@n}��'�b�'剶3ذ�y���M�O<8�:R�S3�*��+��j�nZǟ�&��	ǟ�#l�d�S�? l	�m:�J��K��I��R�iF��'�剥SO��Ү�����O���O�y^�\�G
�9�Lm��٢G*Z\&���I�j�OCS����)�	!��[D��:�M��e�3�M3)OV��H�ܦ���ȟ����?���Ok��p�1�BL�^�pQ(������'��h�4�O|�>�ǉ	�(;���#H#i2r|ЍqӸ���������͟p�	�?y!�OfʓVLK�-yޤy!F�4\I�e�MS��Y�?&mYT~2�	�O�l��)JLv�E�F��lňQ����ϟ����	  ��Otʓ�?�'@�P`�蕍	^r��[�pm"'��̦��f*?	�/��w2�O���'�R�Ō�z�{ū:(��$Z�ꚯ/7V6M�O�}� ��^}"S�4��Iy�Լ�Ī�,�R$b���h*�Q���G}���,n�'���'wBY�4q�G���<4�J�"�$�s�.5�$X��O�ʓ�?�I>I��?	Fb�7S��a���>4�Q��e O��
M>q��?������ ���'+�0����w�*0H-�S�ao�@yB�'��'�R�'N���O$]�R�ǭ�l����߃ 98e��U�$��ԟ���Oy���3X�>�'�?�R)J�Nɚ�x���&,�"�+�`�	M:���'l�'���'�h���'��1®O�ˀn_�/n��!�9j���i.��'��	6f��[O|B�����@H7'
�L�LA��ӛ<�N8$���'��M���'|�O$���1%��BA����[�D�-Y$�6V���g]�M�DR?����?eK�O&!1d��	k`)�bN�ըE�տiG�ɩ(��5�����'�򩶟T�̍c�`q�gC�`�N��s�l,
g�̦Y�I����?!�I<�'gnRy�@&U�Xi����J�B �J��i��'1B�|ʟ�d�O��Y�I'��1B�]�ū���ܦ���\��

��K<�'�?a�'�Ƞ!!���z��2q�V8��P#۴�?�N>�GV?���iZ8�����VH�QC@(a �O�zc��<�*O����ȍ_����cF�.�Hd���3 ��<�����O�����$FF�	�aӀ;Ǆ|k��NBظ˓�?����'Ur�OJ��)�B�4��p�ƚ&�`��i��+�y��'��	ǟtBv�_h�UA�(Y8M�QG�5"��wn�Φ���⟌�?Y���P1$�&�A1�,�2���k������	���?�*O���B�N�'�?Q���Tc�`*F�Aq�1"6J�)s�����O��>��%��b-7LQ��W��fu��j����<���`XJE�.���d�O�����U�3G� �������-�h}@�x��'[�	!F5�#<��!q���d���!�h�j��Û'JH�l�]y�,��7��6m�O�T�'u�4�-?�/��b��X���S���d)�ɦ��'�B�':L�������=���򋛕k�IC���M�	^�ZR���'�B�'9��%*�4���a�$�/0ǀ82p��6)z�HEA���۟`�	o�)Γ�?��+
r������6P�����bś��'x�'襃��8�4���ĥ�,��OF���$��悰v@�ԛ�yӦ��4��s��'W2�'a�OƟ{q%C�'W  ,�a�@���7�O�iۖ �D}�[����|y���5f�і~��A���Ɠ�yؤ����DA�r�$�O��D�O&���O0ʓE�"5P�ă��H+�`O
5��p��d)I�Icyb�'A�	㟬��ݟ���*�5-<M���(�
��f��k �I����	����	ßP�'�x��@�e>���d��O�j��E��8s�51)bӌʓ�?!(O��$�O��d�^�ȼrd �p�ՒKc����1.B�}m�̟P����|�Iry�E31���?�1Ul&e列(
0���b��-pb�l�����'�'�"���yrP�00G���1�~d梇�US���O&�	��'[�����~B��?Y�'#cj�����U�� ���N�`0R����П����0"���'���S�6�4���*�!$2�1�nM%\��V���r���M{��?�����^��ݖJ�.�9�f�<R�Nh��J[9+�@7�O������:OP���yb��U	��T���>iN�8v��0����
OX6��O����O����K}r\���J��1۶�2L��*(!�d��;�M�b��<yK>)��T�'���ru�M�]��e;�Ȗ:�-��zӢ�D�O<�D�]�2P�'���ڟ(��z��p���>��N)^do����'t�j�����O��D�O�`�KS"&��DG�<Mpp!eF����ɈP���K�O���?I/O������e�����ȿv�L��d]��Rh���'5��'��^�@�Y?��p{���q"�M��d]_�,�*�.�I%� �	�8"�,V�l�ѢₜO�����%׭
���myR�'���'��	 )p}��O�,�ZPhX��y�e)K�`�ؑ�N<�����?�����(*��Z���勤K��k�]�i�^��[���	Οp�	oy��E'{�$�.xIU�QPg��AT!ġ`�9�weW榹�IQ���)D~��=! �
+`R��c%�f�΀0�)��)��ş �'�:I���#�i�O8��ExXA�Ċh�4��ϯ
k�D'�p�Iޟ �%fm��$� ��!|�H�ʈ5�����Л������'m�,�dv�@��OT��O�`�Z�H��Z�7%�$�oռp���lZԟP�ɳ*���s�IU�g�? �Ų��2�0�yF$N2W�r��5�i�xJV�s�����Ob�d�t&�����,�L����S� B��f���ݴ @���䓘�O@R  �?4���%�A0�6HYU�T%#�r6��O��D�O�vĎN����P��Y?� C��~���2�J'~�)$��ʦ]&�<��t���?����?����"?����1*�M�T�@τP&���'��]�4�0���O��D.��Ƭa�jL$p0�����q6Rt��Q� ˅�h���'^��'^��*6�  ��p�E��f'��q���%���}�'��'v�'a�� wX)�V-ٙTha���yW�\��韸�	\y�B��=Y����}�E%ЇZ���:DV�l6t듨?A�����?I��ZSZh���K�{3�N�zj<h8�Ǌt�$�A�[���Iџ�IZyҌ�������#�)o��𑳰
%o�$A�n�ןX$���ןP�D&l��O*P�ǁ1~��8WDۖOth�K�i�r�'���@O�]�H|����z�AB���u)r�X�\[5�w�R8/��	џ��I��h3��x� %�|�� հI+ ̀�G�~��ƒ,��nZvy�ǩ0\Z6-Z`�t�'��D�%?�5	��c8E�Q.�}���VE٦�I�4�6�]���'�@�}D,{0
݀c@[�*"4��Ԧ�0�*F	�M#��?�����v��8�HY��*ƞ�^u��j�>q��=m�)x:��?)����'𬉀eC�&]선�o��{�����i�����O��d��Y;�5�>���~�,�X��=Z��g��BL��M;N>�qE��<�Ok2�'�R,V�y��X�U*n�R�	�Z<7��O����Am��?N>��Lv��aC�
�-N�bP�S8:�i�'���c�'��ܟ�Iϟ`�'MVe;"��l�p�B�S�_�N�@��O%#:�b����J����	�=���3��H9IĂtc�	ӋO�9q�������'��'�r^�*������*Ԝ!�8Ɉ�H��Rs�/�5��d�Oأ=i��?�z�"�)C S�N�aH(@�a�\�c��p�P�iaR�''2�'��	� H+H|SH�#
� ����z���4B�f����`��H�ş��	Z?��e˛caj�3�E�/i|m9���ɦ��	����'����2�-���O0���$�%�D�Qr�hQ�g�<+.̒��$�O��sM�O�O��
z.����o<X��!���@d7��O����C�<���OH���OZ���<��O���D�T�_��0�T��-Kn�nZ�������""<����J�<���Re���$��<`2C |4xHj,7h�t�ѬB$������Od�+�Ɔ+�A)�U�i8�-W"O`X��"�GvN��ү�>,� �c�:w:��5;xI�zSt����5i��1���6Ś	p��&3&a߃�*��wD�2(3��ґ�\�#!.m!/Нp[�|#r��"����Sa�	�z��F�<4�}�[�7	~�H��Տw �8�p�hF.y�%�٢si^Z��uG@���O����O�8���?�����X�
(���f�1L��ѻ"��/\��s�G48�=��R�u����8�QJQk��^�+Q�dZ�I
F�4�R�u�t)��?E�*	���Z�M*�̚K�'��Y�lY�e��ɡ�ǃ���Lۻ�?����hOL���4
�xp�ph	�tK��Q7$ D�����2xe,t$5E��a3W�<�Ɋ���<Q3E�����p���TH��a���ڴ�_��ɀU���쟄�'0{��!V�T�*� M���߳�M���Bk�j��q��R��D��d�6"\Э��Ϋ~k�-�a�<�б'H-^����Ϟ�5�����'�bxa��?�+O�4�ІE�	�!���0��h2��$#|O��� �R�2t�Y3$�*
sDi��ORPn��Z��;�m�=H�Nh���J3<ư�I~yr'.5����?9-��؂���O���ɛ>H��+2�`��mKT��O^��(ǲ�q��S�T��i�C(�'�򩁹���`�E4������@OX1��+9�9����H�0��V�Ǯc�l���	\�0��}�>qG����j�O��"�tN���ED��Jz���(O��y"��]�$((�ݯA&6(�C$���0<)�鉥/:��I7�����6�س��A�޴�?���?����5Kؚ���?����y�;$-��q&n�bQ�u8�˅q���3�D��W�d�|AD*�aZR�g�;����(��lC�%��FT�R�T7[���	i�0���|r�� g��+V@-�#0<\d����"08��L>B�^@��"�A8$��	i�<	���P�@���ޭh�� ��e~n4�S�ORbY0���:�ֱi��Z�g��p���|o��c�'�2�'��xݩ�	�ϧY	ucC��/Z͆�K`�G���9� �, ��A��n�#4�^XHϓ)�x�He��*`�H�JΎ�\��T&��b�.3���2d�> R�a�.UR� %�US�b������������?9��tc� ��m U�1P��h'���y��Ř"�TT���t�@�S����'�x����F)l�l��4�ɾ&�u3�e�R����f�0eS�a�I�<�����$�	�|
$�ʟ�'�� 0A�"HS�}8��[([0(��';��،JO�~�l��ʃ45�E��e��p<�.��<$�t���4���C#���<ލ�6�8D���"��1���Q��"MU|�X��6�dcݴf�1��$�2&�d�C\�z��1�<1Ƥ��y�f�'�?U����O^tQ�$�5�8u�Fo���� ��O����&Y����.�|�',���3a�1>'|9wj��V�>�
J�$��h8�S�'l?T�8�([Bp+f)�{�ŤO���'�1O�>l���]�BD�2u`3(���"OJ0����N<�����`���A�'��"=�fD�g�D�z��23��T��� nǛF�',"�'��x8�-XR�R�'�>O��	�_�X�c��2A,<C�L�-
81O��"��'t)r��]Vl{��N4P�0YX�{����<!�-M5@La�a�21*�%S��;��'-�%s�S�g��?q�lbfl�	n��C7e�$��C�I ��S�(4Y��*�@:�#<?y��)§?�����W*]��mA�ō�x���,�-&������?����y��`���Od��!�5b��B.��/��'�� ԭ0�(W�\�-1R]�%��`�,�ƇN,e*C���/1�1d#S�.y�q�,��J�NI���O��$̮mj�C#�7�F-�R�5g�!� -1_ƈA��J�V� a�e�Zc�1O���>A�۸<���' ��O�2�5��׫M�^Ar�؃l�b?O~`�$�'��:�0�Ұ�'��'F��1 CH�jp�� P��Z*Ǔ*�H�?Q�����e�So��1��}X
�i8�����O��O*ESsL��dfl]¶Kں-()�g"O�u�`�kLι#�+I|(�OJ�nZ7KB�D"�`�
L��Q��Xc��b+�3�M���?y˟8�cu�'N�� ��Ҳ6�zKDᇴjQ�SD�'2I_�rp�T>��tH�V��͑�$�-�re�OH9�`�)�S�l0��2��.J���x��V�8�d�'�(�������O+dm��������RN�f�	�'n�H��I�9��@��IЬQ�ÓG���|�7��b�ܣq�ԅ�͒@eZ&�MK��?���sl��� �?����?阧�#G��8Lxd� ���Lv8�k`ژ�'1�Jϓ+nX�{����o��@��#�Cr8Y�=���xx�(3gG�#d*%B ?��H�#�z̓<���)�3�$J�ue �`�@�0d�����
�*9!�$'=xT��Jp� �3G�͔R��I��HO>�D�H�`��0�c���8`�.V��,VOΟ��ȟ����uG�'L"4��YSa����ޑjC�x�F�D l%!����4P�!w�K�ah�P�u.�	h�ܫ3O�!W���`d1��I
%Ȉ�7���'��'���'��O���W,ʥ��Tn�s�2�H�"OliJsHC?lX��l w�j�4��_}X�����M���?��c�iG�Mc��U+PDA��j���?�'���
��?��O t�BŊF�'6Y
1�|X�e"!#
6���![f�*Ԛ7�Ky8��K�K�[iF��1�Ї��L��d
�tJ��`E�tj���
��x��H(�?�J>�ň�Tm�A8ֈ��~K���LX�<��=ge4G�ń8�`�B�LOQ<qw�i�� a��7�Jqn��JwT�y�gގtqV6m�Ob�D.j��ğ��������!zU��&X��Y��ٟX�	&t�R\��X�S��O
l(PE�-(�f����ݎ=q���!�>3�������V>`r"~���
UBY�P�����/�o�D\4:r��ɑ+@L�kA��nw�}�= �!��kz��t��\ъQ��k�� ��=ͧM���tA	���	��.;*�>�ZwHؖ�M;��?Q�&�����?A��?ᚧ��pdA�)�ř��"7�$���#��'�֔��HW�#Ƥ�mc�e3@#_�L�=��&�vx�� ��,�F��g*X&.�x�å��I̓-�x��)�3�?�$`��9B���
�*E�%�!���_#�����PXf��v�-C�����HO>I��U�a0����+#�����PA��+v�ʟ�������u7�'��>��5�dI�
�>�q`���H�B��1�Ĉc.!������ �@���
<�@���E$[=.)+'�\��*ߊF�T���b�$bȉ�6��A���d0�O�U{��S9Kf���@��̬Q5"OH)(�gG5T��b�����C��d^z�2�x����i��'��dPäј�d�X!aU?�F���'\�ֱr�'��I�-�j�Zp�Y�Ɋ9bw�fӜ�P�#��s�8���VD��q�'�-�q`���~|`f(J%D�cؕp;l ��!���үZ��p<�A�ǟ�$�PZF8l�5YQn�?z�*D���G��������9J}C�)�l9�4'||���L�x�΁��Ń��U�<A�k�D�V�'b�?	�P��OD�ZУ$Dah�@��:ֶ�Z��O��D�Qa\�D+�|�'�"�;W��,�p@�1yX&�;M����:�S��`L��6@>N�T0��P9�2��O�	� �'
1O��r��u��-*�"��I��X��"O��#�*P�		����#>��(��'~"=aL��r�Yq��Y�v� ��)W0@�&�',b�'��aYD%�(Y.2�'����yg(
${���(�5{�������z��'�vP�EM׻C�џ�_(��']�+�qӣ8:C����"���3�#9�Ջ`�!�	.�E8�7O&��4뀇I�l�s0�X}Z ZG%�ش�?Y�C�?���,O��U�r�(��&ɯ&��4x�[=��!�O��%��0}�����Z(����t��Pkܴ|��v�'��6��O�˧��i���d����Y� y��WK���?�؄K�C�O����O��NȺs���?��O"К񊓟t��`m�U��x�cY>,��aH�	�:z�y�.Ek8�4�t�:3�@��5@��oP\�bC�B�!K�8lo�U��c�2B�x�LA�3��� �I<V:Ua���21�����b�F�k���p���$-	�9��<K�#ѱw��L����y���	;�n��(O j� �e���'N��Ә'�O^NH��L��Z�pB�W_����'��U��ʖk����ĕ�'dfL��'ȽJ�HKl���b�$!���'P�;�M�� ڜIUKNN��b�'����D�xς��T�MA�x��'��"&��S�ȝ��e��D�j���'̖�#�JZ����kvkR�5�@�'.v��sI��d�m�Ba�:@��8C�'��uj�b;��S��D����'\e�����
��iѨ�;��S�'�)q@/Z�K�6!�׈R4� 9�']l]��������f� %��<��'d�����üG�� 	E������3�';b���� 
)�)��^	����'��1:!)Z�x4�d�d�i�`�
�'� ����G��!�f�V���'�"��v��N���[��X�'�.�WLD��Q	
ARd����'#��eL�9����V�	9D��}�'�|M��NZ�\�Va ��܍>b	�'��`��F���$S�M'����'v��0�F�t�V�9n"j�t��'�P�Z!A@��=�W�Q:��Y��'�Ș��Ôn�h��M�5�"Y1�'�-Kc��(R�.X(�,�=&p�`
�'����{�p�'�J���	�'c082ՋԦk�J���cQ?�Q	�'�BD��Eʀ���
.b(��'vra8��A�$��ri�'���'������-C��a$�p�h98
�'L�;#����Ypf��vla��ռ7z�Oj�}�'ui�u��H��9�qL]54^zM�ȓd|p}�fE[�d��S��2E���ɵo^�E
�'<� ��S �����\;�	X	�_�l�5#�>	��I�8;��ED�1s��(2��Rn�<i�	��nE�����c��!oh��?(�mBU�2�'Gq��0# Ag?8
''ܚ�]��S�? �:�
cUN�	&F�P��$C��ͣW����=���O6��EΏ0$� �`o�wn���"Oƈ�d�Y�Z�	`�ǨA<�����O\�1w����>1ufUiJ���tbWHņ��7m@l��l�'�8u�s���o��!��lJD��'�X�t�4b
FX�t$�7jEnt�	�'���5�� #��JQ�@i��e@�'��ᇄO	 t�H`�dU<D��'w���A� �D�ˋ��2���'�6b��E >d�H*���.�v��'F8M��A׏(��d\��ht�	�'" 0�Ǚy��q�bo��[�rġ	�'�Hz���+O��8��@��X�<Y	�'���	�K'h��P�*��Z�ޅ(�'�v��4
M3)�V8�pė�N \��'�t�"���u��#�,9�y�'A�V�O�W
@Dk���)6>����'���x�J
!)��1�EH6i c�'i M���$_��H���^��\��'Di�U��b������1!j�m��'L�(adAHE�a)Tn��*|���'2� $F?Jׄ���B�f���'�� �e�&E�Q�E#�nX��'Fɢ��SU��H��I%��=�
�'d����%v�@`ÑD:s
�'�V �G&��GR܈z���(z���(
�'�20a���(PP�0ɳ��i{���	�'�b���H% 4�k�O�h�ʁ	�'1� �O� �����D�\����'�l4AkV
D�r%���X�Y$�A�
�'�� fh��t�~e�7.�$CX6AP
�'V���'m@�b���b��18G`ܠ	�'��Ij3@�����3�A�1�ĭ		�'@ě��Q��1�ƅȼ*�����''��PW/�3D2�MI�E��Ęi�'<�a����@��y���xmr=��'�  *Q)L9���u%��Gj� S�'�H1�p��p�$$�p�Y@���*�'ݺ9Jㆄ�r���
aDU	a�][�'�� �E�M�VZT��U�2�2	�'X��Qj�D�l��
A�IH&)�	�'ޤ<@����k�`H0��"@D�a�	�'���[i�8���W��9Z|��'�.X�q�H�zF,L��`�7DU�	�'9��A�ƍ!6ʥ��4[ �0��'Jb�r2�A�W���`ǃ[�R���'%R�9�nĩg4�a�IوB���'i���Pj�.p����Ǐ��}"�C�I�&�(�`���r�)��Ɣ�;	�8
`�br���矰۰>!��O"�a�ΉP��oQq�XR1�	9{x^d��$*��DV���`n� ����.�'"�!�$3m���vНP�ZTM��]�	�?�5���_�D#���ەo�"Ё���6?RFd"B'9\!�d^�z�0t,�;N�[��X�5��u ��B}���̺�����yb��J�$��7�OtҨh����x��N��m�AfԙS5H0�ag7r�c�,�lV�yՃ%�O��&�L?{�`���p���+��'n��k0B� ����>��+�;����3�E?�v�	�$_x�<	Q�� 	:UP3�S��P@1��t~"f�|?����bm)�#bs��T���S�!s
�q�'�Bp�<���}��`�Mߊ^z �����.Z����Q�Ԓ�H�
/fc>c�X�0kr�F0�qg��x���E9�x��kB�w����#bƍA�@��c��z)f�:g�(=*v�X�o�9�KQ4�H,���ּC�9���Z�z�I�b6��X�O� �̲wN�)�x5����+��EK0"O�q;Rd�#}�����$���`*@t~�ލ"� ���U�lԨ#��J�K%�xKŤM4pl��G�e�<y'2�2% ‗�#�@Z O�y 3 \�<a��� |Ҹc>c���Q �Y5�X�j�j����;����%@���B�Q�����A�^��` �>�:[�`���bc8 0�y�s���-��H��	���!�Q̚�?�dM��O�0����+zU��P
L�D��h"O\|Ӳ���X�lI�%I�E(>�s�"O�����9N��
�d�Ȁ"OyʴI�)Yp^��n�)R�9
3"O2T
�E�5��1�L��Y3�i�P��j�L��r\̙�B�8�0|�gF�#sR@����J~���,Eh�<IVhD�Dq0�`G��>t2Ĳ	]�E�K�']v��-��((:��O&M*A�3hP����Bɠbm.Y�u�'V�2��&��	۰���N��Ur ��c�>X0x�a�M�����(��y2r)�,�8��қ��'$�x@�ә�Mc)H/�������u�x]y���!bY��2�͆Qb��:@�D8f����rN$D��`�����횤�?2i�,������f�K�=ST��*�%�����H��(t�1AI%>��QD��߼ G��<\���.Ɂ
�BP��`h<1�k�������؞h�`����.6@�WハY��͈DޮA~���pk���ٯ;�"P��c��/d*�I42��FHJ�=��-����v"��DK�9���'<O�D#E�I=R�ѹE�ݒ�VT@���\\�"���?�^,jwa\7 ��]���Pr�.">a3$�a��d��g��^�\ ��aO`�Z�L �'a�<єR�=��p���]AX�D��/(*�[��
ZcT��d��;j��򆪂��a~"�]a
*�u��.2:0颇Y"��E�' :��ƨ�,�	p�M��JpB\����N̪�!V�i�`0TiC"F0h����C�̤ԡ��=� �{����	�Uφ(��̓5�7����Upl����9�0������	��<	�nE-O�^�JG7 ј���QPx��X�JF5$��ɺ:p"�:�I�!tL��@��:Kw�C#J�X�G˜�m�J��pO�d���9��dV�+< �K��,̴�X�a�$��'Ĥ�a�f~�)�(Y�h�� �)����s�-EW��cD@L'���C�f�$��Pp������dX��Ԕ����7Mn�s�k.k����'��)���8�)��q>���ٍ2�n-��wޱ�dƅ�p�up�ST���%9D�L[��G���f��m�$�#�k��Q���4h�?,�m��^D��6�����-Rz��'ɠ%3$	��H��@���x��'I�$1p�/`
� ��ګ>�����e�%]����*Bl���� �Y�q�?����LF�{�l�C%O�B|�u��	Y�����,
��O�C�"�A5�
/~�����x��!B9è��ɑH=��Bq�Ɇ3��(3��Lp4�OְSbK�B`h�9���N9�t����fi���ؽ�-��A0T��'y>����Oy����I�7Cb��p��S��?�c@�;
�y3 �^n�'�����T
�Ж	�XG��N2�!�Yo|
����M?5V��D��v��$�¯��.��dհ)�$(h�z����e�L9�p�c�ͯ2��h&��#,�S����|����!&Fe~d�`b.�K��ТF�{H<H�\?�5 �'�1o���@�ĞV�� ����'���<a�j�MK�Jg��*��x��hh<�eK��}��}[�#	/�! ��V�E��h��'@�C�D��Iז��U�	�&�jϓM߆���y���&�~�O3P:5���"�y"(*�X�� �_K�1��씩��[C�����doW�m��\:��$	��}Yu�	�y�ѓd�YC�#=V�-�lU�Z����'*�*dZDL���/ޠL��E�	�'�Fe`7.,{v$��Ȃ�,���$bUr�!���?&�d����*���hN��y���"1O"-� OK�)B�� !H�t(���"O�r�)�-���j��^�`��0�|2�_�h�Oq�,�&�0��]��L�
q�B�"O>���9�BbTkœtfF����͊U_0��DA'�h���)>\���!��Z&#��BF�
�,��eH�üEr�O�����3ye�����ɛ0�*I��"O� �2�$��E��4�w�+)���1"O�ɲ�g�>o�$3g�
��2�"OL]� e�bO�#��-h��L
�"OBI5ĽAZ�3!�Шa�&t�"O8�X� +&��t�0d�6w̜�I�"O���gYl�����ϜN����""O�ԡ��Τ!n�!�)O�!�"�6"O�i1+�	cp��E�K�kI�T)�"OlD+M�ll��gG6,r���"O����f�gR��^�8$B��V"O(��읮u+8�2BbX�r�"O�d[B(�-~�F�˶ �U�"!��"O���&�'k��y�a���:���w"OP���\�sen�����r�ʥhV"O�	��΄�"{��S�<:rF�c"OhURnx&P�*��xx��u"OL�de"&��6�W�/�����"O\���?�zL�#���kЀ�U"Or�����	r����+h�=`q"O�H��m��	&ݠ��J�$�� "O<(�Cţ\큡�ǸB9v�U"O6�A
��7�*m�Tj��Q)4�y�"Otha�}T꤀#(L�Pɀ"O$��P�^�+K�2�ȡ�FKZp�<�a��"6�����B)i^K7@�P�<Ydf Ti�D�!Q�	����J�<�t.�\<���(�\g���5OF~�<�"��S9��*����9fT��v�<��揟V�D!D�D�:���2#B�p�<���@<1��2E_8
�d��.j�<q���25�4�w�µO�vㆨ`�<y��1��	�2(�/9
����F�<����ic4�3�ǧV,Ա�Y�<����N�R�Q@Aj �z��p�<A��?h��"#!N�<���BB�o�<9b������sf�5u�J%��o�<A�d�-�T��"&.|�m�@#�i�<i�)��+	VM˰��9�ё�	�q�<���T�x���jN���`�l�<��
�-=�tur!��=(��A��<q��D\�0-���]�`I�s�<��Ɗ�.Gf���G�6+D��*
v�<�1��� �h�p�A�:ƾ!�"HMr�<���	(�u�rYl��(���X�<YG��-#�x���#�z���"�p�<�4�U�_,��8 ���8��Ee�<�s⇫c%ju!��@�ƸM���c�<aa��N�I��lX�W:>�`�Kb�<1�k�8ՐH��݆+��8yr�O_�<!b�3O��\�gNV��<���aC�<	rJ��	��i�g�
�xqJ�����f�<ɕ�_�H��R��T �i�<�%l��b��L2��D�&� pG-�i�<��Δ=M�@��K NbNa��"�h�<Y�Er��Do���1)c��e�<��6D�d�kE{o��U,h�<�2�Ҋ[?8p%��E� ����j�<i'���m}l��cOɊ%��5
n�<i�˝�7��\���TY��d�g�<Ym�$]P�d�7��2zD�#U���<���ʚi ���%��jK��B�hC�<����^��(@#kY�;Ĝ�ʢ��z�<����p{B�j6�����TM�|�<��`����S� �R�A�*B`�<�  �b�Mм?�>=q��;[C���b"O�Y�N��N���!�+<b� �"OP�Ч�Oz���C˃H}6A��"O�y�Jܖa���A��_��d"O��z�Ȗy�)��ڲ(�����"ON��#XwA��⑦��U��-�yR�ɖE�����`Dք��F���yR�
"jd呇.T�g��Lه�)�y�;��IÍ��b�3'��2�y%��1j�Y��Х]&��Q`��y����_���4��s#�=�����y���"1�a��ǔj{�Y��f�y�D�s���R@=cφ�jG���y�GP�-��5劈[6N\4���y�`�rOm3F�Wdl=�V���y2HF�-|-�׊��^��D�f�B�y�S6�����ݟC���a��y�� vۼ�P7n��9����e�̱�y��Q�z�K�E�(c}�d僗3�yrA����/D��ڬ)���yr(��^<� �Ѝ^�*�v�3�y�=hڐ=��˂��TP�l���yK�7�c������$j	,�y�@��^�^�7���`����e��y�*�S���S�F�i�b��㥑��y���7>�S�kקh�lL�-� �y��"�.�Igj��UF�}!g@��y���X���!3�ոD?d\r����y��a��`J��׏8K���R��y��61 rPk��@/�thZU
^�yB���F-2)����U�Y+"�I>�y�@V�yK��Zc�����yr�ߌZ0		S��;Tp��C^��y��� ��`z�Z�b�]�ф��ybc��&ݸ��D-#���Ѷ��y"I�>	:�P��L�� $����I��y��#
	�A���tf[Gf��y2�B>�D	6��HfԪ�'Ο�yr,.\H��"���("b��b�	���yҫA�F�d�W' �d0�(1��'�y"��v�Cg�WC��`�
��yb$: ���1��Lh��i��Ê�y��I�B��(ִ0~�#�I��yR,�;FX��e�Z�� �ũ"�y"GL�'�,h�!-�) ��"uK��yb��$8g�
hJ��#�'�y�c�Hf�����)1��c�?�y���8v
 ̉�.W''�6#҈[��yB��- ��bF_5vǼFq��j	�'J�r��I�L��
J7�|]��'|duK�+a*2�#�|�:tb�'~JySfEbˢ�8���p�=r�'m�h+qBΖU|�(80'ͱQkL%0�')�p�WFR�hyq�*J'J�u"�'B��pjׂp2�@
W 4\IA�'��)�2D�Iy��C�*���	�'��|r�H�#���`-��)^��	�'��͹t�0H Dk'/�+�$(�'9<���i���蘘�0��"O>q�q��#p���dg��y�͹5"O*h�F�?r<b1  <5��"O��፱]Hp�#e��0T2�"O��tjޗF��aqSD�i�|�`s"OP�FG�5hr�5�ѥ!Z���"O� ��j!'�`
"u���I��5"OָsƊ��_��L����5!X]kw"Oz�0t��\��<�'��W��a�"O�1)&�D\�����&l���"O��3SdȰ4�Z������"O��bfQ\2p�_��hME"O�M�)2����(�l Z�"OhnFOI��v������&�(D���7	Z�h���3�	F��yBd�'D�SW�@//��Q�ӡ�*1��T%'D�P�f COn1A�/���M�q��z�����d^
N.�q����D��8c�J�H�!�-���e��@z�8賩M�#!���'
�#��Fw�	�VZ�!�d�<29ny�Td��0��ZQGT�N�!�d�4yT�`1����ش���4/�!�ªt:��*�K��&����d�9$�!�I�*j��r�bC<%&�!ƈ��p�!�$L�m�苗&ߝx�P�gۛM!�d�E��)��� ���+L(!���wy$����ƚ�:(����6�'��F�iDqOq�RH���7d�y�.U6l`1b"Op��H�Ep|x��,�w��%����IܓQ��I���L��2����[u,�xSG�<?�����-D� ӷ�F���a����΀@��/}����p>�o�:l0\tsp�M:m�,�%�^U؞x�T�|r�_�OA�6m���A�*	��y��f� b0��e&	�ò��'fb�q���� PL�48`!S�Hr�P�3)�y��2�9	$GD�8�2����yL���@;� ތzK�i�R���y�ԃ���"N�	<Pa���yrɏ�j�\��G��$�p�劷�y���|�]P�W�(�8)J���y�D��s��[欖�n�8������'ў�Ԉ��W�kEB	sF߁f��!�F"O�#��]q�ԥA�DH�B�1�"Ox�A�fȨ#�p��7����5	��>D�DC B�Fd�A��-*rD� >D��4&�� �У�lp�C�;D�����ƓZ���R!�4jz&��B�'D�tѓ�K#k�=�%���2����!�$D��)`E�J��`;�FP�:b�!D�@p��O�`�n��$E*`5(	y�� ��xR�ҭk��A��J��Ïם�yҏ͛%FsQ�ߕ���%Y��y"�ցpQd��U{1l��B˴�y��J�1��'��6z��0�K� �y⦁)C�����,m�\�ڠ�ܟ�y�Q�n���h����ś�CB��y��
�lbt*r��<�|�x',F�O\���ߺ��t�0zph�'��!�$�9&�1�$�*�42�/Dy�!�$�'S:�D�qď0��Iv��G�!�HuW�}(����Y�P�C��V�!�ć\�`���a)� ��0R�!�ErR��b�̚0y�� $��(�!�Qi�0�M�C�2��W�O�i}!��7���1�摀+�T� A�G'L}!��b� H�AqUVŢ&��Q!�_��H`@g�z�n�6��
�!��p�jD[�( �T�Hq`v�^�G0!�^�m�0pӀ̀�wqLA�Ц�t!�$0\�H�$oP4'^�S��4 R!�� N� ��"��	�&֘<��!"OP�!@��$c`0�#f�a�tȢp"Oԅp��$9�$"�k�Z��`"O������x�n�Rg�-]�V���"O<�*W�_=j��xGNs+�[�"O\�0�E�7� g䏿Y�� �"O���H�'� u���7 e.-�%"O���3��O��yУ�&a��i�"Oz"�C�.zf���%�"O�5�S��K�Z�&A�t4�I4"OL�3�#��h�����cU;%����"O<H1-��@ԞC
���a	�"O��g ��q����n�����"O��[@郐7x°�@���~q(�"O&P+��F��(�J�G	fy�T"Ot�� -S����ޜ9���K�"O@�0�"-�<�rWL�	y�a�"O�ĳ�L<�*3k�E��Ԫ�"O�:���;���S�i�>�@�J�"Op�R�k��"D��"��#�ȼit"O�ܚWL��8�D��5@��U��}q�"OP@��`'2wv$�`�T/�Ta�"O�i��˘k>V�r���f*v(@ "O�\��"�!r�T��m̸M"�y�"O��@���7nk�5�6-�LB�S"Oz5`E]Z�{5�D�D����"O�j��O�8����,/j�Xp��"OZ����������<s�"OF�(ga]t�.��>*fʐd"O<|Z'm��e_.��&,�?c�K$"O4�ڡl�#_�e�W�TxJa3g"O�
f�Z+h��x8%���fq."�"O�Š�&9M���I3`�t�"OT\�O���������!"O�|��!��+2���"�zѪE"O�4�&R�z8�P�p���h�~���"O��A��%hvk'���f�8�
�"O:��D��9��<Aa"%Y+��Qa"O\�)�����Q��V΄��"O�Pe�4�|���l��yQ^݃@"Oj-[���9���i�[?Z�k�"O�!��H�VдG���v@��C"Ob���Er���)�^�-��ٙ�"O$M��R���Lڗ(�ҭA4"OP���HG�Q���P�Fo���"Oة�kĈj��=�4�˃��	�"O@�C`Η� �|�Ѫ����E"O���N)h�>]QFl�B"m�W"O.`� ��#c<�P´ ֙{	&�A�"O$���S%�����_/#�Ruy�"Oƨ!�Ȕ 7S(-ѓ]Ty��"O�9�ϗ�V�X� �m���P��%"Odp*�@I�p���Э�+}*YP�"OH��a�:?-\1Q��HQ���f"O��x��FGz����e���R"O0���ׯj6$�	����>!�L�"OJe�k:��(#��A��# "Oμ���JI���BL��Z��ԃ&"Oj4��۸Bt�3�	!C���"OZy!����~5�3�ٌm�r"O8�0�Y�-l(e�b�G3\r���"Oni� �?@*,��B��6g@r�"O@02���iup#�ѢWK0MS�"O�횔#��sr����I�5>4�"O� ڰ�@XT�0�aJ�i��87"O0�A���A��*D�-=���"O�-��mY�dU�8´/Փy�(�+�"O���%Ė]�X����,a�* 9S"OZ�@Bn�1��l@���UBX�S0"O�Y�  Q�fw��p��U4��"O0�
�Ð�uT�P0�,ƍN#|5p"OvUk���
	_�t�aˉ:g\H*�"OLX�p�����q��1j��1"On���@�|%r�it\ ZP��e"O⤙�MK��A���Z�0C��"OB���H#S��Q�c�}%=�q"O�T[��>�
d
�M���X�"O�ГQ�
iox	�� a��5�s"O����'.���z�j�7�pL�g"O�0�$�C�KFZ �� ��b"O�%᫔�7�.\z0K�r�x�Z�"O�Y��D�*�����o,����"O@Q�5�B7�T�O m��@v"O�q1��	x���Z@hďg ��"O�%u�2Dᩤ�����܁�"OPHQ'��	?`�t�wFJ�2h�lBr"O���$�ȭ<��r�R�F�DӶ"O��(D�X&U,�Q񆝌)6R}��"O0ma��D���ah��}.���"O�鹁��K��ӡ�5d��P"O�l9p���IA4�34���u��K�"On�SƋ�k����T$6�$Q��"O��p-��/�l����# ��<:�"O4�8���,XZn�(�\�Y3"OZ):�H,�ƭ�-�[��aAd"O� ����H�i��i�8��"O�� BF4?$�����l<� "O*���F���A3'��=i��ӳ"Or�iWdE�S\���TeE*J��+�"O0�1�㛋���X����b�L|3 "O�蚱���su����߲R�z��@"O�PVM�;2�l5!F�C,_��A�"ON Q��.}��2 ��R�� �"O��Q	�n������w�0`"O��&��:&�ӷBS)N�l �"O� cE���Dl�!��N�%��"O��7G �r)�e����ne"�	"OЌa�����r�
7`�:@"O�{�̃g����L�$2AC"O��ᡔ�6��A���lH��"OdT2�b�
##�A����$7�%Q�"O�8P�E7 �@�D!��,�ؘ��"O&�q� ПOư2�I��3�"O6D&�t����'H�=����"O��Yvۂ`��D3����~�V��#"Oؠ U&_�Y9�颰*�
�~���"O��0��*�P9�c�цz��rG"OH$�S�1?�ڔ�'B.N�T"O��8�ܘe�n9�Da�P���8�"O���Qb<yH�9��"ў����"O�Ɂ�I,9�UA ��3!5 ���"O �J'���e'�|zU��;l��˂"O�wn@>QL�q�pA��g����"O~H�%��!(���u`���T35"OޜkB�̀���:��P���ա!��Y2Vd
Pe-y�T�Y�"�c�!���D�J�c�A�J�6��S��+?�!�d�i�2���h�W���w G�"u!�� n|c�)Ä,K��гgL��"Oޱb6��	Z�x̹7'@.@��{`"Op�
��ͦ}-FI��ߊ�#"OL���{J�H��4h��0ڥ"O ���!=�:� �����2d"ON�!E�� ����4��&0��<��"O�!R�C�>٪l��H�l��  %"OV1C�ꅯT��� h8kB��A"O�@���RJMJWFA!(N(�+�"O,q"6	Ҍ<�	uE^�m?�d��"O��zB���*)v9��s�`�"O(�sK�p�"�Gi�/��,u"O��ض&΁J��Q3�-£\�$"OV�:�)t
p`׋� �@8E"O�ps�f�9
fHx�)��{O��"O8!q���88��p�Ё�.)�"O�!BԪ�*A�E�T�b�b�hf"O��5F�)vER#3	�,O�d�"OL@&�4gX܂�MЧQ�zL`�"O<� �枇0F�"�nO�C��۷"O<�:��C�[۞P0-ʼ$+�ŀ�"O<�؃&�)(�baa�,�$	��d�t"O�u@���j�8,U-��v��u[ "O�9�bBA�v�#���@�����"O�0kD�5?W.�d$˨9���"O�Ś�+V(\yP�H��*���yr &%2ܭ����:9�f=j�lL0�yr&ފV&��!m�,2zP,��+^�y�F��%�����#<,	K2n��yO�.\gRP#�V?;����6��5�y���.�2@���1. �X��y2H�`��ң"4*Q�Ř ͪ�y"i�nq����^�K4@Y��ڴ�y�g��u���Pc+[1I ����d�=�y"	=f��I�⣄2F���(N��y��@��ruS��W� F��"ħ��y�`Oɨ�Sw�~I�xp Y��y��#�
ĨTŀ1x�ؑ"���y��W'�}r�΁k�:K1����yB� �`��1��\�f/��W�ħ�y"ˆk�<�j7��d�p	٧o�*�y���0=b@
ŎZ0Z�X��A��y"�#p�1QRhQ�d��2W�T���xB&�29DՈT��\`j$�W�+kr!�aGh�+����s�j$�Zu!�Ě6�J���"�7<D��K��F�!�$� q����k�	 ThZ�`X�!�ɤ}Jٴ	G0)� ڧM�<�!�dL�x�Q��$�10 rx�DbX�-�!�N(~P����10:�IP ^�Bu!����
�Aveޒ^������v�'a|�ˌKu,�ӡg�:.��Ff�.�y�+�"F��lxd��52�,��j�yb��Z���6��2�
#���y�2t1�B�"l���ɢHЅ�y�C��AZ�a�W���Z���\��y�k�9A	�]�e��P0�*���yB%	z�9S _�
5��!V��y����yhZ!�A�����ȍ�y"�]"D���i�7rY�� ��y�)�����)ED3z�H!c	ط�y�
����/�� b���IP��y���$:�t��X�"��<A�F��䓑0>C��F�jy�ԡ�a� �Ȱ�=T�� ��B@5��xK����^#����"O���dj��Eh�=�e�# �91�"O&庀�C�f�xA�QJ��%��T"O����O��F�iY1JG1�L�V"O\Ո����̱A�h	+$��ӓ"O� vd��8\�hH�/�����'.�'����>��"�?�|=�ݚ�rQ*�#y�	A���OP����ИP:`���	5u�T,��'P�+u'�e@�� ��gh�'d�y;0E �?��y/�����'c���A�=>���Ūjyr�'�$$���\9i�$�*:v���' zM��e�Q;�E`$i	�b�'�L��T�ȗ#�҉�S�µ��M>9������O
�L�E�=zB�<@R��}!�8�	�'�j����::p�1���sʐ	�'E���CE�iv���.��d��d��'R*(�1�9��e�'@V11Мx2�'P��[�NΒ2A�4�	@�*��]��'�ZM���X/�$x�H%���	�'ܽ�ao�$[���M���08����O���>�B�Bũ\�`�� �&p�2����3D� ����	�~�P��1lQ���b&D�8���4i���F�p���A$D�ȩ��Տ�0t���N]��G� D��[$�&%�r��6�M���4D����I��.A��V<N<�P�1D���b'
+�~�:a#ׯVt���2D���3`��f* ��t�Ҫ"��3�+;D���A�S	U��IF��6J��@��5D���+�<����a�ݜH���H`H D��s���Y%���B`�y�$,ِ�>D�DSfA�N/�y3E� V<���%0D�@+f�@J��k"DèQ)9*C@:D��㡭��!32�0ӫ�%Cep�O�O|�d:�)�:�|l葤���"���D�>�"���'�u�A �Y��8��Y72�9R�'����#H�+@��Q �w���'!��á��<����'B�g|r���'�8���
켄���o�H��'�|���6���/��j���xߓʘ'(�P3�`�6�)��Kƴa�(I����?q�����"�����PSii�/�? �C�o�BE���^�� �)�!�D@�v���C� Ҹ������]�!�� v��d��'GcɌ�{�ʃ6�!�$�N�.��!f�*TW`�Isk�7D�!�DL����z�GG�j8�)Kªܔy�{2�'��	������	��NnT�i�L�\����O`���O�˓��D%�I:A&�e�t��5,u���!3-�B�	;U�`)��D�W�.11���l�B�I�f��'�>b~��:d�L	C��C�I�������:u�j�QŜ�b4bB�IP°tEV;D�0�`ږ��B�IDnLQl�� �&��_�
��D�<Y�'�|��#�s�[e�ZF�KK>����)X�^��u�`#��k��p���I�!�D���Ԝ9�&�&��ҷ�ʘ�!��<Y�Y�%�R�:Z$g*[�!�d	l疱�	���Y��ɝ.+7!�D��度H�"��`����R:!�Z&-h��1�X%m� �	�G�>d�ў���S�)6$s�g=�F�37��S��B�	'j����*C1C&A[�⊊y.�B�)� z�b劘4�h�h� �NRr,*B"O�����$�2ag��@;f	�'"O�k��%Co�q5f�_.�Is�"O��˧ޒ&l���Z)Lp�6"OaY���,2ҵr`��d��jB�.�S���xH�P@��?ڔB�Zf�!�DW�8U7ώ�p�� �!�[-3u5ɐ
�8
A�Ġ�9-!�wӬ�e���:�A��g�!��q�}�W���.��0$N�E�!�D��I��!�IȨ4���#�+�!�� ,�ej���:M������
Zўȅ�ӛTb �f�Ŭqz���V���Oj�O �}��@2l�rؙbU�b�*P!xɇȓA��!��%^_|�y1_�j�쭇� ,^�sGAϑ@i���$�ڕD�<�ȓzI���"o�>X�"mH�<D�ȓF-}����)J��UKr�QpNq�ȓ1�p-��ʭT�޵�� iB�ȓ����A+��B(.p��W�^����	hyB�|ʟ0b�0��bݹ@�&�)%1K��e���7D��@EŧU��h��hA�u=��e�+D�<G 
���HBO�*� ��2%*D�d@bY�5"��+W��8��E5D�D�����5��G�+I�6T8��4D��Z�BA��T	�A�P/ZL00A'�OD�	W�.����4nY`��74|r�O�����.�-�V �8������'9*�IX��(�0��v� ��6��3���X�|i#���2LOB�[��'ra��x��{�˘�y�!��<N3�d�a(�p�	H�!�$׼X�xؓ3�^�P�*�h�"s�!�d��YΒLI�,I�s�:���E ġ��%SH�O�7�(5BcҚw��T��	��2��O��X�<0TH��C�I�s�xXa�"��J��B磒z��C�	�m��$xnԻ`�n���� \LC�	���!J�DǙ-jV�����C䉪t���	��]^|  ��6�$B�I�?�E+jN�M]F�@D����C�ɥq�Vm��Ė�q��%���Y�t���7^D��U΀3 ��ÒA]�'�BB�I�f�l���H���	�"ɩ9��C�	1c���)t�:Y�p� L��C�ɓsKD�� �nt^!��3ϚC�ɳD9~ �'ȗ�Q�p*D�;w�rC�;�P��P�*�.�P-޲�l�1�S�O�F�S�R�X��a����f�¥!2"OZ��2)�,T����B�jX:�"O:����$;!�L2�'
�l�� ��"Ov��6�	�G��(�$�crh�3F"O飦��2,���%^5�Iq"O�<�v���>�8�Sbԙ �@u��"O�B���r�ś���te�Q�	Q>!
M4e�]� �N�h����q�<�����4]��KY!y0ei��@�=2��"OLp�a.=6P�����&� �&"Ole�]�4G�R���R!D,ч"O�lp%�H-(�t�H4e

J��"O�ܑg��-.�D�B:i�(��"OP����x��A$�>�J 2�"O�h���3v���V�4,�}J��|r�'�
�'J`��vb�0h�����ˮ""�����xL���^���`�a��+W����S�? ���Ǎ:���#@A�l}^I�"OjH�g��#a�xP�%(Q�-�XT�4"O(��w�8��1[��	nU�i�"O����D�!Ih�HH֠O��т"O���C��&~#�4ɡ/�nE����"O�bi�1Mq�ђeD�n�D "O D�T��>���D��0*a"O��{���^2,8q,O.~��I�"O���'�B�o�.4�"��4*�|QB"OHX	�k�8W �X�!�ޒ��ٻ�"O���4ˊ�sw����W�h�2p"O�Y�ao�w��VI(��.I�
B�=M����g���F1����(d4&C�	�_�F���"
8�8}��M�6f{C䉱��|�D�N(�L��1g�1��B�I,��ꉢJ&�B�e[�J�B�8��+�O��l�6���N�5�"C�0�����V�tS�G��l�C�Ʉ�d��0�K�R��W��]�B�I
`Ä@1gł�c�ҥ��hM�B��3U\:A�"�R� ��͇r�B�	23_z5aК�!���ƩM�B�	�>7��t �u2�-Q���F�$C�I�N���P!IҾK^����c$j�C䉮\H~,K�-T�_��A�)o�B�	�F�f��dE�j��h�rG]�w��C�	�R
�E�0��6�@Z�j�#��C��oMМ�@�S^�8�J�U��C�ɓm7��b�۴[ .1��	����C�		{]F��A�(�&�:���"qЀB�ɒ$ē��@ ܰ��G�F]�\B�I4?CFl�&E� �v��DkF'(�B��}hx�3�ڋ<'j����ś3��C�	�I6|h��8x6T8e�'b�BB�	�ELj�;��׊w�\��
�DW0B�	�}<�0t,��1K�i��`A9Hy�C�Ir"f%�`�Y�j����@x��C�,N�L�!��.Wӎ��e��B�Ɏ�����F���%kW�83C�	�k ����e���;�хn��B䉙,|l-�1G�?��ś�ЮIm.C䉲DU,��g�ۙ}��,�*��B��B�	av@��Έ��J��F�q�|B䉆q���*ƬÀz�.�����Q�C�:P����A��
���
'��^�C�	�Q�������
�eF��'HC�)$��	�W$�6?��樀�<C�I�t5�"w����"��D�!9�>C���|�GE]�+�Y#ĥ�2!VC�I0�\H��G�r��Dr�^#S��B�� [k6�AIY��H��ۗGݸB�$Z�^p!D��2@���3��]5��	�'��"���>�H�!��A�W3�D	�'4��b҈��:H���դ�� ��p�'Z�US���&0��R�*S�Kn���'d(%H�-K�bwR4�+C�Ɣ�Y�')�@r�[ =$B���*� �H��'� a)�R?��i�G@�,1���'y���鞽;U8E1���S����'ײyX����h4ps͎�Y&�c��$2�	or�7C%XL�9qS�ƫRt&�����<AD�)r�8R�ތt+�)��"M|�<a�/�<(��pC M�z���l
yy��'0Y�ы[4F
؍i���[�-���� P���M�>�e��2(�`%�#"O�aI�#S�-=��$��!T��P�U"O0�j�kJ[(4���gy�8�"Ob��,��\ٔJ�1l~��p@"O<)�צ
�N9�)��C�xq��_�H����4 ��������i�e�����O���0=�Ǭ=� 1cZ�X܈�b�M�<A�'�b4u�6���P1A"�E�<��%�8v�� G��d�L��jx�<)�%�f%����(w\��E�Kv�<1�&Z�p�����a't���@�Pzh<�v��}(Q��@[�X+��Xv�=�?�)O6����4ʘ� �F�wcp\V���'3a|rR�[n��������/��y�#��B��]9�OA� �1p#�y2%�� /��2�	�nx�y��d�7�y�k�+c��ҦǼc"���Ō��y�	GI��a�W�N�\P֣4�yJk���@Ϧ5�뢇_,���2�Oft� �H5�I��ENt9�!�!"O�R�f�yA� �dc�$b,;T"OdI�B��_��l bT�(Ʃ�&"O��@܊[ɸ���@�3U�b�3�"O�RB��:E�q�#��X�6q�"O`,3&�,8_J$�Ə�AЬ@q�"O*(P���.-> Tk�ώ,q�\TR���|�Im�ďI9~[<]�B��G�����+W�y�'�3��\����DiȀ�+�yY�THtA�"Kb�Ũd���y�o�W��ɚ4�Y/S�޸y��Z�y���
gH��e���L�0 Q�U0�yr�^/:;�)�Al0V�H��̶�y�K��`�P�x=$�|��ФI���'Fў���<ɠO�;*H�@ɝ�%���wJ�D�<9�%T�P�����5u����UA�<�F�˕x���ŨԆE+��c��|�<!��59��T���?��A�b&�r�<y7 ����C��}��PZq�	d���OO*�0T�O�M$�	��Ϳ\/B5S
�'V@8kU�^�L����R]�a�I>A���?a����O��P�Y0x��������*!D���"�<{[�ઁ#����:D��QU��-%��|:c$��F"�B�,D��3oDI���C�	j��њ�)D�TI4$ҹ0������̱1\Խ���%D�DĂ˳@�[��+�X�˧!#D�軀@�-%L���%�	>|�L��<9��hO1���Z��ªRɨ�c<��e<D�p��I]��0���˰= 	��;D�{ ��;�$�e�J'L��AP�'6D�|�"b�Ls� b�H
7gܢ]b��0D��CM݁V��h�d�/j~y�v�/D�$
� 2Ei1"D�r��5iԌ.���O>㟄�<�w�\5>����JŇ$�RQZ!��D�<A���D�QņT�MÒ�і�~�<��#�����mS5G��a	a�^x�<e��/iҥ���JN"݊c$w�<iQ�Cp���'x�>��r �<Iã�=oi�0������hk�П<���n���Q@�E�r�y�D�z�̄ȓ4�=*�A�,k��!%@.xX�ȓ�(���0]5rgE�%K\����x�1��Gܗ���⦐�Q��ȓ�]!�F]������̦|_ą�S�? (h�%�N�B'Bu�q�ՊZ��("�O�������`���y�1yw+D�X��ي2'��0E䋨~��`�I'D�xq�F^<GT� R�l�S���I%�&����T�AT��0s�0(2Wm�6if�2"O�`����kDD�d�8)���*�"Or�{ӄّD����V�J���R"O�\��nº<��y�ARCP�D"O���a��CB�( %d���'�!��	_���AI8,��Lȴ
�/\!�S:�	��ǌ�c`(ʥPџ�$�$�O�p�тG�|^����K�K3��	�'v�I�,\ 8��4+W�+z�	�'��-��Ί�4(���F��'`��'q��z���_-D��W"�(�'��x�D%��D�b�+t��,O����4� ��0�P�N����@0��<�	�<���ÉdbL�`&i�7���%�H{��^y��'5�O:�9��1�gKZ+L "��K#"J0�"O�x��)� i��	r�p:@"OJ|Rh8��Z ,��\�Vų�"O�񥞵I˦�10ꆗe��5P�"Or
b��V��(2ъ�ͪ!D���3��`����M7:�e�f�=D���&�]�I���D+�'&��3��<D�� "K�|4�`��9�Z8�)'�D*���'�[ÅY�@�X�	��6�c	�'RPD����c�f���Oɫ2[bXk�'H�p�T��	�c���+�Q��'_I D��"#���B���v���'�����AN ۬���㑬Q�	��'%�C�� F��C�-ޤ�
��'��i�҂�<=�����]4�[���)�4aI����|͂p��M����ȓ6��9B0�L=K������;����4�P�%�;��DҲ�Q�|ڂ���:tb,q�+WB z��ΘJ1������0�p�آ7�*,zA�U�<���H<�Ac�9�.��pɀ��x�[�l�i�<�W��%^r:��3�d��`C��hO�'�R%��:a��BpmQ4l���ȓj�ryӊP ^��J!�N�Oޤ�ȓcd�*���n��8���Uv(��#���(��Ԍ5���RU+��ȓCT�� BW�V=|�(� _Z.�H�ȓUʰ� d-
�8����M L!���F�8�@�]�MY�Oͳ2��0�?a��0|�򨗑|.ƀA�I0 ��Fx�<iqՆqRUȷ�M�t0�EZ�<Y�ۤ}J�s��{bB� 5�]�<��N=/-r0B��΄\s&Xc��\�<їHF)2�6db�&قJ?�4`l�m�<y0bD8ZD��'琪9/.�8V�A�<�U�H�0r�*� �T3�0��<��BC6��0*F�]�;`(�ð��P�<�J�5+��Sb�'��l��V�<!2`�:V��Y�hU	M����JS�<�D��0x�@������T���1��c�<�p� W�D%z��6 4}�$����T=�=+m�*p�|�@�&����7[ʭ�7��>&t�C
�rnŇ�%E\hC@/v���d}䔇�Q\d%P�����};���i��,�ȓ`�L�f�!R��I�byvm��S�? �=R����S�X<�^0��P����h��k�#$��
o�;@8��g�;D����P�c׬]K�a��T҆\(�,'D�<�.�*;}�E3G*�@���"#D���G�^.C j-���V����"D��*��K`��q��B@*���.D��h�� ��5��Ĝa�H C�+D�db�b�;[B8õ��DVe���<I���1A��ܨwI�ж\�_�&�Ԑ��o<���[�#jtX�e&+�,t	֥�o�<�F�E>ex��I��:���(5�Dm�<�ሿڈ8�FF�ul��D�JM�<16�@,�(Ыǉ�ܡXT�V_�<yg۵$4���F!�x�dm��C	A�<���ɸu:>\���QI��E�{x�(�'6Z�rb��h�2�;�aW� �J���'� Ph'��
4,�؃��t1�U��'Qh��Q[	-�
\����t����'���p``��jTC�(�f��'.(�rG�H��8�a�����:�'���Y�OǊT�D��(<5�3�'�v,#DMG{!)��vF�c�'V	�� �$	NE��oP�{{����'�0 F���*H����	ok��I�'�X�` T��vH(�'�`L�k�'Z6e��,{��L�M� Q�(p��'d�ibE)ׂK��6
�-N��@�'!��1"�h��MeI�E+��	�'Ì�7��
 �B�)�(�=�� �'*}z�n��}��ف�쌇 ���
�'�p�����5��/�#B����'VH�9P�ۓTs|��H����5Qϓ�O�����ŤuL���b�G�@YZ�P�"Ov�c&��]B�i�P�E�(T�"Oh)��3-���ZP��PH��+�"OiphB�m*i��\44��S"O��z�[�I@e�g�9Q�>0�A"O޴3v*��US���D^� ��\�"O�,�ш,X���%2���"O�d��[$$!����+ڀKij�"Op���*��),�",�F��!��e�
����]�<��bL�~!�ęf�F���
K�����Cq!�׋E�B�P���5 i�(���k7!���4[Ek�F	:Ă�1n��h/!��1A¨1&�PP�X��+�)4$!�DAS� �kek��`L��s��U�@!�$Vˤ�� �7��A"��B4!�Ę f�,ZՀU)K��d:�Eݕj%!��&� P9'ٮ[�����I��R�'���'@�)����O�n�����m_�1����5N̜{!��?"X�KR.��p0I-bq!�D	�;9L�Q�m�	t��e�ӻ|g!�$�$���-�*	R�Ұ�N�i�!�D��6�<��W!�43��y�F��b�!�$�5P��m���)��U�!�d&H�8b�N��U��ֺ�B�'v�|ʟqO�c��&�4��
�66��"O�r�ڛK��)���A3f%X�"O6i�ƈQ�kٚ�@�jA�u����D"O�-#2B��s�zE��j�P����0"O����M%E6L�p4cڱU���cT"O�a{2�%+��ܳC�:8���;R"OX�$M��Z�@��&���kи����O\��;��3� Px��jċN�	�ƭ5���j��d�O����P-���RQf[�##����  !���'&Gt� ��N�g�N�I࡙91Q!���n��k�UQҀ�!F�.=!򄔖_��� &΀�4x�)B Ɓp%!�D#y���J�c��g"�5;R�@xw!�dK#��ܹ���1���F��-�!�$�1�r��� :��4i���}��'�ў�>���j��O�fa�A�D�ze�v�7D��A�`nHD�g,I<xRI�2J)D�$`�F�(N]�"�̉Q����9D�衴mZ�f�KB$�m?��۴�6D����V�en�b�)4�b��v,4D�`Zrm�@&\!A�F���Rf2D�h�Q�t���Q�6o<���(.D�P+Wi�%T��*���|�Y&�.D����$*N\�b��=P��c /��9�S�'����L�B���d�BJ�-�ȓzeBEɊ�-A��M��L���c�*P �e��[��C�<��y�ȓz��u�����4~�GF!Rq����3fI���(�*�z"!+3�'� F{��d		����M\�W�L�p�a��y�@ȗk�y���:�z|�6�V��yB�4�
���1>��i�&n�-�y�h���߶4�v�c�'
�yR,ݸf��;��+B\�LBl� �yB�I@����,m��٣��yC�'�zY�v�}U>��d�۷��d<�S�O<6x��!3�����W=5t��
�'+�%YU�W��I�Nҕ%����'@D��1'�1�X��KȚNz,1�'4\��a�ШW�IS�UNd�E��'��x���	4�<Sr/�	u2��'�\�BG�1"��!n�YW���
��-���L
���B��ZQ�(#
�'f���K�/u�m�>h��q��'�(-cA��P���`ӀL&3+"��'�PM�Vg�.v��Z��L�;-��
�'��E+�'�0XBڔ[%*81���	�'T)r�K���'�/e��|�	�'�1u��-y��\hb�W��}Y��hO1�J�O�JY���y��(���&J�P��'�&@��"�O#u �,P+�<��ȓP�@U��G�1s��P��)^�����Ųs�ܿ,���0�>
��ȓu�))�$�<�h`��%1��ȓ|��B�
O�Mw(������>��ȓ?�hsj�����Q�-�2c���ן��?ͧ�O����΄�5�2��&I�����"O"@:C�5]��� k�.�'"OL���n�j5�L="� �2"Ob�8�
�2B�
3鄲Au����"O�PցT�c�L)sp'^�v��"O�	���M N����&F[H�t"OH��_�H��x�R���*U��Q�PF{ʟ��'^2%�ujF�[�F�NF.cj�$��.H: @�_~T���$5����#�I���b��u�&n�
3h؇ȓ!�l1s�[��)�@M�5Kj9�ȓ>���A��/r�(�%
2HGP|��1�q+W�3ͮ��o�YQ�}�ȓs3���F#J<O@U��*Ѵff��	k�����	6;\���+M^��a`��]|��B�)� �4�uH��%����`�u�b�����\F��ŧP��a�#�ư%���у�y�f%x6�i�Pjшڌ���`���y2��+a�\+R��e��;aJ���y哻<o��H���[��qkw���yBGB*g�TDr@�ø N��/Ǌ�y����/��P�AC�lBl"���y�,�1#�H�y棖"��`wF7��O��D�O`b>�ദ͔C)��+��+����"c:D��ce��%%�
��A\�!�~-1Ɓ"D�t���awh���]�:۾���3D�H�G㞝=5�� a$Q�<jƁ� &D��X���ӥ��';xZ}c��jXRx� Fx�k��I.������/=��R����y"�D)
t`�C �/�x��S��y�d״?p���,<�k�)���yr$�O;	�g� �fQ�N��y�ǺV��ɻ�0c_��f�@!�yҏ������(�A8DA��yr�_�w�ZԳEN=����D���䓗hOnc���T�Â� X��D8v>N����&D���3��Ti��8��	&��sc0D�ĘT'�o���u���P���2D� B!��.je��Bu��2����L-D� J�\�^�Αpa)W�I �R*,D�D#�س5�\l�Ħӌ�� Tg)D�p��c�1�l��CD��O��  ��2D�Р��_3M@p��Hb�P�k�g1D� p�j��!����҂�!E�<	�q�0D��H�f�
D�Y����ʲ�/D��xk_�XQb�3�y���.D��{AbƂD&��0�%����L-D�����Lh��D�0 ��&"��yD� D�p�BON�=���D��<:?T�`�o><O�#<)��6 �s���&H`|#�GPr�<�a��Z��	6�Ј�d�"��i�<A!ں7��mi�hW�Fm��GO^�<� �ܡG�h���f��qA$F~�<����p�e�X�H"�Ls�<!G�L
[=<l1u�R�H�ʼQ���c�<���M�8�ш�B��q���_�<���׍H�1&'H�[�Q�^p�<I�hK<&NP
rY�#��@A�h�<�㌖D&�P�󥁐c�`=ɴ.e�<���&����d��,�� �g�<� ۵"[���P�?(��R��[g�<A(y��:��I�@��*
�_�<�2Bb�bPۓLܑ/�L�Z!��]�<1b/�4�A�(��h�y���U�<7*�%���:F�_'o^�uKh�<��!������`�<� �D�c�<1t��X�^@ےdO�N�Aʄ��`�<�&��9nb��ee�(
u�@���Qx�<���Q�JS� ��!8�Z�ˉs�<�hD�2��G��(V�1���k�<�𬑰d���@b�((�g�i�<�; NI5���7b��T�i�<�ƨ_�����N�.�\�@sIEb�<����cNt�BC(-4��9�(Dx�<q1�. g�$2K�p�9a��i�<���
{�QGŗ��%i���c�<)� �;ˀ���\�A��x�A��D�<aw�ôx
��ȿ:"tI���j�<��C��D��C�/�2+���I���i�<� �A�T�����y��A �ih,��"O���eF��D��A���҂M|	��"O����o��EJ� ���ݺ1IV1pc"O��3��\4f*��1�ޢ^9,�P"O�	8�,�W$���4�@1��2�"O�ب��YЄqF�6*�k"OС)E M��x(�҅R<=%��	�"OB�h�O��F���bЄ7
����"O��P��3�:8ڇa�;um�%"O��B�ӌ)���JژS�Ȭ�C"Oz<�`S?�v��$�:g����"O�3�uZ��Ԉ� |�ܜJ�"O>�+�mU?B~1�!�
;S�� `"Oz��"9�੢�Y9"�.aQ"O�	CW4;z$+E<�2�$"O�K`i�PVP��i ����"OT�-T,Πhp���ck��"O�ę'�ة}�`��'֪&BR�"�"O�MH�%�#0`N��'��U4��"�"O�=��e�0b6��s0��Pn|k�"O\�3�H�,p��1���|���b"O� 	p�9!�U�A��n�1�#"O��q��:�`}�BH
G�Hm[�"O���r퐠|���%�C��r�T"O"�u+�.�J�����p(i"O�0"�h�@*e 7_��T�6"O��
P�}V�,Ke/L�9.�Р"O4$�eŧ0�CrMR*���"OF��1E�'Jv��Elڒ+�ځ��"O�q� ��� ��B�Ѣ"O:�&��3l����-�D�t��"OjIۗ�F2�ZYy��
r����"Ob@r-\���ѻ&C�3\o�`�"O�h7�Z�]�J�-��rr �"O�f�Y.2�,���z^� `!"O֬(�>n1�a����^:�X�#"O�ݘ!Q+�tx"�̠SV�:U"O��C@
��=����ba[3'��mZ�"O�A+fm�U���H5�	�-j6A��"Op�&aɝ0d4���4.�U�r"O�Ű�%غ>�".O�I��u(�"O���w��/�6 �Q�9w�
 ��*O`��3�W)@�0S��X�PZ:��
�'Tb)a� N�Fd0Y�HX)���
�'UJQз�ц�~�i�D�T�z��
�'�Y�0H1=S�i��+�K��L�
�'攴*#��r���('�N���
�'�9 �\.���W�Mn\XT�
�'�&�5�M� 8�) E�a�D�
�')^����\�I�@%Q$dL6R*~1�	�'P�ͲwU�����#.�;	�'#2��e�9.x�(�9���	�'�F�0�`K�M;F�ѱ!�n߮�X�'����B�5GuTb��O$gт�Z�' IcZ�#���dc�-9�'�"����T�D�6��(��c�i�'Y��z3 [�b��ŉt(E&��9	�'�hK48��AX�b ,(�ʨ��'���r����X�Ė&GZ���'+85HqdK�/�lJ��|4, �'��aQ"F�AshO�Y�T ��'i�5(�T(M5&�����h��	�'} H�#k��6cdXt�H�^
�q�'e� ��N(�F�ۃ$V
�!���� >i�`�\�l����#t�D"O�,R�N�Y�*%AEߺ""�HE"O�|Q� 5L"Ա0d��;Ȁ��"O윛1�/K$h��O]d����"Oz �tE����Pt΂-M��c�"Oq� ��W��A�t�Xw��aC"O�]9��u��B��3b"Hi�"O63 ]�2�Y�Q��<�~�
'"O6"��%gƼUp�C��je|0�E"O�Iۃ`�6��1�#>\y�� �"O��!p'S<
�����D��T)`"O�Y�Ch��~A["aҹ$���P3"O���Z>^r��!�4�|p�"Od�h��U�w5��r��}�+ع�y��\)]q��b�fԉ.:�A��U��ybL�73��,��Q��E�c�U#�y2�X�%�<��s蕂N�B�	�O0�yR�Ʃ9�I����Kx�q�+��yr���>M�du�A�@����`�A�y����E�5p�B_��d	ޢ�y��S�<�<�:���'1�И�ϙ�y��+P�.��$n��{,���Ğ�y�I"z�	���F����ND,�y�$Dv�Zg[F��i�tK̪�y��-�j1��W8>L��{As�<�G�l20��qi��3�D��k�<�5dL"� �RAڞ:��� �a�<�ć۝k���fi�����_�<�`눦6��r��_�~N�H#D��Y��71�lZf(Ӌ$�����4D����Q�s�d��?C9B���*O�QJwc �!�c� G;(�D� �"O���d�@��I3�̾{p1K�"O�I�a�0
>��sfG�(n:�"O&�� 晈;6��I�KL� n��C"OPѳ���<iiFYe�ϮvX�"O���C
�B\��)�i�~KR���"O��V.�4�&�[3�L+A�T*c"O`Up6��A!�\2��.F5�Zt"O2%`�cP)[d�4�G���C��t��"O��2�fڃh�r�2���"O�QKr�  \$tI�Yvp��"O��k�K�?�m���ށN��G"OFa��j�����K\	 b� �"O����n�;4�<q�D�[��Y�"O����,%F���h("���"O��mK�y��;�H�mP� �"O:�)u��A��]h��KY>��#"OLQpV�zF b�c�Y'����"O��ZĆN9g<ti�)�>���"O�!%@�d|��tǗ%p�F�jp"O��ӓ
S>�Ĩ{���OI0� �"OH	@2דW�(X�����$�D�"O�*���qf�����;$�JT"O��C͆4�z����B(
�P�v"O� ���F�jR�''޿5����"O|ȋ�i׹<��&,E.3���9�*O B7D��%x ��v>>l��'�,+��
�\�,1q�m��={�B�	�"έXU��7DP���FaİY�B�	-S�4���|al� ��5��B�Id2V�ӡ�"�D�jvME�)�B�I#8>^d��_3g����#N�ND�C�ɢ*�|�Xu����L���!�lB�)� ���Ў\��FT1�J�Kv���u"Ol5z�G�]8 �Ӣ�	z|�!P"O��J]#!��:��4d�`ˠ"O�]h�ȡw\, �C
�(XBd%�"O\���CK�o�Ƶ��#X�� I�3"Ox�s �ĒR��(ҁ�7�2��e"O�����<���Y'_�Ntl��""O�P�C/	�<��H�Q:jD��3A"O�) �hCP���)pU�4�f"OP��1e�F:��C�<B��K�"Oݠ1�Ȓy�^�J�h�� ��b"O���g� ,�\��նSB���"O��҅�͗(�"�I�&�a�b�c"O�@�c)����A��)$�uP"O*��!ω��Б�`�t8,q+D"O�HrB���4�*pz�U�M�)�"Op\q��(������%7@la�"OTu�#��<WH��A�&�C�"O�H�P��,"I(=�&�Gnm` �5\O<c��� F\ΔDH��)ls#t�����-M�Y8�h�'<E�=a�" �n ��	��ē)�tT�X7�L����22��+�"Oz����Xj��ʂ���D%*1�%"O�k©w���3$�����i�"O���Ř�(�s@_�n�PH�"O&a�Ƣʄ(��� R"�>I$)w"O��I�$[?&2�����.=J`�!]�L���{�dIy�,�;+$���$?@�B�IxI�D�$ܳ�B1r�n2��B��0�`Yz�K�P
ŚW΄;'���e����'p���>(��Y
�h�����'� a����-�,�sx�xCA�	T��y����"7'�2Y����I
�yb���\l5-�1�<�R�M�y���4^��``UVL�@��D�O��=�Omh1��ށ	�B��┑t�՘	�'(�0�OE6J�|!3��o���'�8j�J�Z��`�ҋ/m��	�'	�ݳn���r�g\.g�H��'��<bF��;;�yB,�����
�'�~hz��M9)����tL�<k���4�6�<E��4��X�q���ap��w�^6�b���V��Ṳ��tw�ɩ� 	�,�� �'w�~����'�ġP�D�*�� �ti1�yd��LlT�W��%3��S#m��yrf�%�P��O�
���ɓ�y��d'O2И�Ӣ5 ��c(�YHhY�U"O�삄J =\��jw��8��"O4!��폝'�t���?q)U"O��:�	� %�$MX�E��7"�p��"O�bq��Jh�-��O"b�1��8lOvIf$�1ی��R��0_�>�:�"Oq�7l]�r����(ԓ�l��"O�+ql�8b5��\�	k�lST"O�0X���� �ah�@�&n�Pg�$)�S�S�H��$�'�Y�u�L���d��-w�B��%7=D�ic$��|`VѩǢ̤V�$�<�˓;���aI�!k�����O�X~��mZr�����ɾJe�̻׉��L_t�M�*T!�B�I�i��'��:o�N9Q��'R������&�S�/&7��Y��M�t� &��c�^�?����đS��%.�0U��HdAS=U�OȢ=���+��F�F���9�,��;��:�P�@G{��Ʉ�n�}���\���੗)W�!!�� *�is�C 2v�a�C����H��"O&ݡ��1j��u����Q,����"O���'ݘ!㢝!��ĳ&~�0�"O��ą��&19��P�ep�ِ�'QqO��b7�#*{�I5�����I�� F��-~�<쓶�?2�̴Q`+Ă�y�˄�}Bh�; ��U�E(nN0�y�DM���}*��TS�B��m�:��d/�>ɕ(ȉ#PdH v�w�t��!Rmx���'6�Q#$m�5'x���ȗ|��
�'�n�9�̏���g�S<�-`�'���bN0N��V$���
AÓ�hO�Y��I?ߔ����L�N��P��"O�8%��	f!j�x�)Zm�J�t"OHI��� bJ��b.�,�x=�w�<)��3^z�<�jI�>�h�d�@X���O���6���*�O���0"�O���V0^�. �&���RDKe����x��I+G�R$�ǃ��rf��Pօ�
f�����?ړ3�"| d��X�*\��O�W�D8�O��=��Q�Y��Se]�wL���im�<@ѕ<�&��/2za��)XQ�<4i[���Ț����X�J֢�P�<�ǆ0&�<X6��9��%όF�<�4%֫_�
�Xm��\5�YK�Ɨf�<��Áx�:�$�خk�d�@�DDg�<	G��r��غ�o�d���h$C�d�<��MP�u�r	�e�"0��KS�Md�<E������9i[�|@�U!H�i�<�e$3d�pu���Y?܌�l�_��p=��l�"P,RW-��@�����P"m|!��-2ަ��@M�\f*M�7*ڿf>!�$�4��!!d�YO
��'G�u�ax��ɩRW$tIv�)/\�P�0Vc��E{J|Z�N]7
U�Q��Lt����g�<ɥ��q�!�����l�z�&a�<�g傆(�ĘB�Ol�p�S~��a8�X�0�����1��_F9xfl5D�)���J����!)�L�]�&D��C2*,F4��f�� �,"�M%D��s@�?��ئ��\���)��!D���B�Ȅ`�>���<����� ?D���A&��F��`3a[�L�D�(7-1�$=�O8e)v
�Y�T��I�A��@�b"OL(⧏D�t���i!Ņ�oG�rE"OͨG M�T�uX�L5���"O��Iӳ$f�Re��aD��"O���$��5�]���SF�ⓞ�����)�'P@|+��[,Xz��"�H�n�$`�IQ<��Z�J�{�v�Oq̓�yR��˽�����N���qP�ոj5����߰?QK�o������B�jQ����'�ў�'g,8lZSC��h���EA	Â	��z�r1�f(_ɀ��0�C� �]��aB2�b�_?t-Ճ^� (����Nܓ�2�s�	 <4�"�R�H54��ȓ,C�8�C]2p��!� M�wh� �>������Ĺ%���%���v1�e�T4�y2, �u0Z��e��2pt��'�Z��y"NM�b�)��n�c[�RP���yRo�!πAC�BQ�\2�=���۬��z���O�X�;�a\90צH1��?v�PA wI.�S��y��OR�(��o��o࠱� Pp�<��	]�^�̐;�Ȑ��oZ2�y
� @��Я�`7d��2�E�]��`�"Of
�
�v]��i��?�"���"O�t$��?�D��"�]�2p�t"O���EJT���e�B�<���"O�� �h��N�����/_2-�"O�i���,�N�@K�8�X3�"OJ�(�(��Ea�t�G͇8��B�"OV�P��E�a�H�`D�R��D@4�'B�$MYM��
���P
T=��GQ��	C}��� ܮ8�*	(k܅)d�
�"��#?����9�bq9Bh��z�n�JP矋D�!�DW�a�j���B|m��X���Ik��(��᳴�}�`i�7a�N�T<ɴ"O٫���$5`�̢7K�e&q�V�$4|O���qIS�z8�$M��1J�ٻ�O�\jf�֥����Ι+�\y�V+�q�<���	W��]�0��?I���@CBw�<1�HĘ=�µCY;4��d����q�<郩�2nO�q�G�m�:�C7̖Q�<�snHb!�G�F�I�f�L�<Q% 4<����%�\8e�^�p�f�]�� �<��B�#�l����� aωZ�<�
*q��5��D):}&��S�<�c �.O�B��i��;�Az���S�<)&���v���c&C�Y�V��M�<��d l��C��W�_k��j`q�<)d�FA��ɰ`�:,�"B �j�<�`iR�Y#b�[���q\z���Bg�<Qd�N�t��U�l��B���|�<��E�843vE8&HS�dx,(�@�|�<�#,\m��M�
=k�
Sb�<��͊6��Lx7�L���z���s�<���ܓ����h�6k�P�eK�e�<�W.V�0" /]�ءRTa�<�Ũ�:@$���,�$py��F_�<�,�%-�@�c�%ӥgth���_�<)"N����X�~�]�%�@c�<ɱ	�^ �h:G��,�������a�<�`o�{֤x4��e�a��_�<�&'�t~�u@`�sJ|�� ]�<i�ٕrv(���0O������V�<	q�J�4�����FF|�����[�<Qɯf�ze���Ϣ}��!OO^�<Q&�ӎ"�٨�Ϟ� 6�y��[�<qc5x���E w��E&WV�<���4&�AAԧ�Rf��$.�I�<���G�.fV���'�sB��Y� JC�<�B���J��	�F?\�03���@�<�V�Y*w-�q0�f�^)z]��IF�<��@*n# <q�%I9c�.����@�<!a�V7Bbl�t��7\{r��PGD~�<�����ؔD^�c�Ґ��"�r�<���.Y�Z@�$�A��h��Y�<�'A��v��t�R�������E~�<���Y#)���'��[�6d�ՀB`���� C.s������A�A��$U�/y�tEo�vD|,�%c0D��pTm
�%�!O 	�U�L;D�`!q��L��=��n�l���Շ4D���7M@�!㢼qc�7d��H�p�5D�h 3F�+\�%�Pʗ&@��t��a1D�(Y�nK�@�\���KI��m�6�,D��Y�A0F�B�G*`��m�b�!D��� .�]_�x�GG:R�����!D�����j�Z��@�ŦMg�M���"D�� <�%Ă&9��@S��PR�,T"Ol�'�ɂK_�p���f�X��"O@��f�.i�-u���t�[�"Ou�'��1zB7��>7-5ch<D�p�d�Z���P��F)x���4� D�X�w`ZJ�6�{��P�eh!���?D���I]�2Gb����<P�"g�?D��h�ň�G*��k��H�<)���=D�LrV
�;�j��3J�-~�8Y� �,D�h�6��G��x��ɉ
�5�tC+D��J�;�D i��ҿ7��H���,D������ �l��A�ʔ�DN-D�����E�@!�{���`9D�`�!��f���K(1KxT��4D� �7A>z�dx��:`:���*0D���ׁ���qr��@�PP�E��1D�`�L�
��d�/R�C�`�@#D�|aE�T6[U��y�cѨR�FoH_�<!�N�-�R�8�K��6�ȉ��_�<�p���	U�t�TMԩkI�qh�b�<�c��2lݾ-�E̓�os.i�b!FX�<AEڸC(b<R�٪]��ђ��O�<I�
@�b��\�%ګ%E$��E�<�%�ٯ����WbZ�r���KR`�h�<�	[n�<x�e��lT�i�0� k�<����I�fA�5��G�p��b�<Y'�J
Y|���RA���A�\�<!E쟒K���7R9�N�j��C[�<y�n�%Hm0@�Ζh�T��g�Q�<����SJ��p �N�n���*L�<aŇ;M���Vf��L~�u!�L�e�<����t���U�J�DMPSa�]�<�u�����'�J��z1��[|�<����I�De��0x���Bn�P�<���[�	�f�t�W�5b��S�<Q���7QVh3���$.�H,2ap�<��ƪ
K`�r�N'4�F�$�l�<�q�\>O7����TV�Ԭa6�Ak�<�ЅՎ
f ��̢lv΄�QO�f�<a� +>�P��L�X��H2�T�<y&�=8��rO/tA@�W�<�r�#Z[\ոf����-�UI[L�<���=t������;Р��L�q�<�v.C���Bd+Ĕo����g�F�<����1O���)J�Q2�A��F�<1�^��miA�R�r��q�`h�t�<��ˎ�F(��.��A@�����~�<)GBZp����=�^=���u�<c�
_E�ń�tХ;�%D�<�φ8wV������  �>����F�<�Ŭ˨J}��R����"i�ت }�<���&M����gE����b%�z�<𯈆D��rl��Z��*礝r�<�׎^#1cFT��K:;a��za+�i�<�CN���Bd�� Wm5��f�<��H�V��cA
ʊ{6�4l��<���U#	φ�@�(��i-d",z�<��H�:I�=��	4�pxA0!J}�<��k��CZ1#ӏ�dp^�#�$Xx�<���$wɰ���I�1e~�\�b��s�<ِ%ҁ$�R�b�造h�l�$-�@�<��I^�2U�܃�a��K�6ɂ��B�<��ˑ(�Jrf��lS�0��Ww�<Q���L��i!(H.F+8�3!�y����Q
O�H �T>O� ,		�/�|�����D<4[���"O��x����Z0�%�a�ϑV3J�2#�O�T6@�s���E��}z�E3�I(�%�;#ԡ�#�Q�<�2�ξt.��{૜�Jh ) ec�5-���s�b[���d����?�'R�1jdM�6j]Ju07�\�y�p9�'�"���ȕG)�y���MC���F�B�JĔt94%�2D��	(S�Q �>d���bZ�;d���Dſu|��q�[�=n�$�eO�WtI e���n=�ĨţgC:C�	�k�`�uÆ�z�f����
��Ob���L ������A7[3h|�偠.��3���'f4�Lpg�Y�<��錸zZ0�W+۴'��ƍ�?�ڸ{a��2{��Y�`"Q+h����O��A�O��9U��=Kk��1BOLT��L,x��q$��8a�� ��*S�ƠY���B�*�CV��ٰ<�#)�{�����:WK��U(ax��A Y�TL��%h":�F\	C��?3�b��T��eC����1�':T;�㊗[�*�s�Ȋ\z�њ�y��^���@÷U0�P���"��~ b��ܫq�~���C޺;0B�W�V�����,EA.%�rCګH�P`�*��f��2�#�?��!�gy"�U:���qw�L>E��aY3%�)�y�� z(��iB�a����"/�4��V�
}��"
��ٰ<1e�D�#J 0s��H�;��"��Cx��r/�P@�Au$I�6촥���K-���"��V?UF����B��D�E��w��̣���),�}�(��J�p����O��x�2@P�m���J�)J$Q�(%�˓[�>%)��3�dת��r⩃25pj�c�H�I���N����{��	E G��q̓�6a"��6���dw�'n�lHэ�C�S�R6��5M��:�1h�HI�}�t��'ptK�L��i��y"�!��X`�]�{�ҤF�O�rFqO��G�x�6�K
�rEn�9���9�h���A i�VI�f�Zh�B�	�:i�]��ʊ�L��h�b^��5^���<�u�^��<� �$�S�zǰ���"E!7�|��֬��R*z��Ai����ٻ���Ho�}�iB�}��	�u+��m�Z `���C�x���O?�Y��^0F�q�g��0`���gb�Y~�X!`ò5j�O�2I��G����9�����ǕdZ�@jV���D��?�p��G�2 Gay�/�$褐#f�h��QC-��2���Aq�Ί�?���N7�ȼK~n4i��)ǆ^30+�E8�Iٙo�Y(��hE�vL��c�~��؅a��(2��ܔ������ǣI0��4� ��U���)��O�S-���ˌ}T��S��-��"ж��)G IU@ �&����O����ƁM1i�☙4b�����q �o�����h� hl��ȱхW�.Hjp�� ��)�����eB�-�t]A���r⬐����>y�kJ�%޴C�������=ڧ34��r����`��Ƞ�C^o:%���h)C%ć���|���j�0�q��,'<{��D�Kޡ��t�H��P�ñk\��<���'+ܤp�	�4�li���լ^dar�G��9eC�v�����Z:S��<�����������a����L^�@�!�j\�<u�	N��8��	� ��S��Q-�΄Ӥ'̺)���K�,(ҨO���	L:Hqژ�h۾a����+qݑ:���	K)�J�(ɘ|z����)�r����-&��ҧ���a�D�GiպO���g�:�~2���Ť� )s�!0�Pa2|��IV�-���DK�@u�=�r��([�I$[�z�㬙U��8�CA��#e"��Z`��B��y1 `(�N�1R%
͓��N*�T�O����+�P1��4c�lk1�2V�\=��B�#?��܄�ɫ'3�e�#��/T�3Rl
�X�%�t�*{ر�0�D9&̶8�% R؞|��϶9��D��Ń�U��C@�%��x�#6S*�)���<qXt�Xwh��r��&�*@+��5c�h��'��"���"x�&I� aHf|�ҫO�s'�J�Kp�V�U� �[w��]�p�	ٮ5�\����k
�l����	�a}2�ö$)��o�=���)n���zSn�O� ����"�ژ�vH��5�Ju�t1��$��äi!�&sL"��P*V7x������Ybѱ�����u�h�j0)^	�f���^�)��Eak���``L&�O����f͏Ln���a�+��пi�Ԁ�!)qܓ|l��Ф��;[|��������7�MA+���k!��8	�!�D�%d�����
v紁�1�)Y�	�]t@���܌k�@���Rr?�����[���{�H6'�U3F�25������fm,8�U�'�����S�dW�S˃Yg�Y�\Np�J��Uf^5����ݪ9��`M���懬�, F{"(A6k?�  ��5dW�?�Ą��@�	@\�q(�_Bt1���m(�E;� c�d�@#�@�9mʥ�ȓ;���n�=�H �b���͇ȓ}�i�2`_"lP%Sǋ�"��a�ȓC��h ��IWR�qm����E�aR�ܢ/rm+$e��ni�c�d3d
r�S�'O�dx�2
�9'刵��'3b����J�J���[$4��fb�2'tԄ��{�Y�9mHc?O�KcZԩ��9�T1�DO��Bb%̡e����H��Wy.�3g�!]� �	�����E�D\� ���2P�^��	0��T9��|�Tz��	i�(�<q����/۱�yB+֑at:���۾Y�:�f����|��YhW�"�)�Ӥ)��48���x�,�ԯ�=M�L�>�b����H�Z9P6IvC�2�\v��;��5�	�9��A��L<)j�%K��Z�,��>��=;���<�4AZ-Fʖ㞢}���ìb�.L��؏a��x�r)J
?y6�:�'����F�.R��t�`�/�����O(q������=1A*L"lD@Ae+&��X
6 <�O$C�.LPa,�z���t]�a�� =��`S"Oȁ�"��$=;���
��A�T�Q�ɹ3[2����S�8���㖫D0Q�&�S4 $��B�	&>��I�:8}� ^`p��&D�k���Ӫu�tDb��wo�0���VB䉂H�ԔyDM@p!�T��)�%e�'�D����'>��A�΁�V��]�/��9�'U�LK�ح�P �!ȣF ��'W"��"*�<���Z)DR�'$|��F-Y4|���J� ,B��
�'M���iE 8UL��)�-����
�']�n�|@�pF���.���A
�'�@Uĕ��0\8E�@�	�'���f�
 Yֵ�'j��`̈́	�	�'�(���HѢ8��E��ɘ6gˊ��	�'�V��A��/m��}`@��+X���'�~aV(O�#���T�"&tL{
�'�R	�a��&x6��P�T�Od,�@	�'c�azcW�$ڌc$?g���'�%�bnZ2Q���!��УF%���'pl���&KDi����Z�M��-��'\��% �F�j����,1`j���'���h�ꅀM6���@�A21
�'�*���I\�zP��x`����'hh�	Ѷ&q��fO5m$��'Z��L���T7��~p���'g8���Z�k��H�N�I=|PK�'���q�VNi�� �\�K/���'!Y�˲XFI�u�+���0�'���2�g4<�����7R�����'���K���X�9��Vx��	�';�S�O��!��$��E��D�p��'\����%�HQAD�:iĽ��'4^�*�f�%��`�d@=��c�'�h�2fʓ<s@8ԃ&`B�*zb�0�'|�xx�m[�`�Fe&$@�}�
�'�J,"4	��T������zH�	�'�L�"�,&A�M��>��`	�'� y���S9,x�J �S*|�n�#	�'�4Y�.ۂ/[CG
� �jݸ�'��=�_�@��ܓՌ[)�T���'#b �1�L�����(}�X�+�'U���"��b�AH!H%p�ɻ	�'�J��C.��	�ZB̕7���'�u�d�(qR����
�?�jL���� P4Y���z� ��*�4�c"OX���Q|�@�q�gOF\�"O����'(4�P��
Dn���"O��Q��k' <蝥x(˖"O���0h�;A�rQcPjS�f"�q"Oh�M 0��4;qIü�f��"O�U!�FA�����x�(���"O�;�E������p�P<Ye"O�i.E1��"`��i��(�W)��yb(V�"�Q�p%��eG�P��*�y�#F>]O|�X$��k��daY�y"��o*�q�����q�	$�y�G�:����H\8�jЁF)���y���9S���@ @D��yˉ9=��Hj�A�u���h�� 
�yb,G}m�|����m�y+�j���y�DQ 	�:�+� ���@�2+�?�yR���+��9)e�Ɋ*�Ѳ��8�y���L@��$��_�������y"�� N>x,&�81�� �y� �R����&h*��r%�6�ybM��a�z�	�,���
�M�0�y���001��j �ɩ�Ht��^!�y�)�.L��7n���qvY�z!��� ��&hI�Dr1@���ڵ"OD �uDJ��n�rF��D9TX�"OfIA��G�n����@�9]B�5h�"Odi �%�_f�5���6I 9ht"O���S�	V�`���[9���"O�`�����l�z=���;4jjM��"O�D�q�� ����'�Q:���"O4���FصM{��V��Z
<�"O,�abHKs���`#fA3^D�9"O4����|
§�?}T�|:!"OX5붍��*� S��φ1��	�"O��a'L�V�8��wb�
#
��T"O��0�ٲj�����U�_ê�y""O��y����/����"��g���"O��.�in� ����2CNԣb"O��Ґ��c�H�Je(G� ��"O.�8���! ���*�g߀2�"лa"O���1��9{��i�R��jsL�x"O0�)Ba�w�l�X�+;hL��"O�В'��=w
A���!N�q"O|�yB U�Q�µ���ОJ�=�0"O(�{�ѓ�乢� K�0:�� �"O8Ȫ�.�01��ba@]�u=� R"O�4�۪,K�l ��Q�8<)�"O@���=xTD�R��W:,�h�"On�z��<h\^�iꁧ_�`�"O�� ��)2�@��>	�$kD"O�q����?_�����G�BZ!	"O��rU	,��@y6ӳw���Q�"O�}��b�+o<��oè>���	�"O4�z�BO�-L��ò��1(U*m��"O`%���%k&�fI	2�l���"O�HJ���l4�2aȃ��bIzR"O�TC��0yQ�z�
��-�t#�"Od��r�ћ~xd�G��*d� Y�$"Oָ*`'��vY@�E�m�
��"O�x d�\)��$�"����2"O��Y��AE���n�B��5h�"On���a�Q~z��5f�Z��<�q"OX�
 |*B�B��[�(�nq"O� 
�����a_Z�I'
I:O����"O�I'��Q�D(�tlF�{����"O�D8�j�*��
_ �qR�"OJ0�R*ܶr��H9���&	�J= v�'S
<��	��S��Γo� L 5�ز ��U���O����ȓ;�
���_�4/�ݢG����<�gٕ􆕒)@.�h��U�P	S�=G�aaI�,���"OTp
B�I�y� ��&�2��¨Ŧ#c�(��Ar?q��ė����	�(�"� � �?��s�)�5Y��B�ɄR�Z����w���k�n�T$q	���/e�h�)w�Y�4�a{�d�$g"p���`���B�ʋ��<a�c��f��<ʂK	 N2@ )ԪB�L��,2��Yq됷�yb"�A�~e��� y���S����!|�̻�#��)� )DIW� ]��ș��+��\���(`V�mӣ"O
ذuFG�48�@YV�D�(�6.�^kld�Cϕv4d1I�+��j��� *�xEI��84�U����S���Ɠ���4o>1�D�rD��:kʽ�u\E���C�
�(B~^���<,Oғo�VfU�3�;^v��A0�'WbA�C�U:]q���"8��x�oū?�<��Ff
!Ap@���	gH<�%(X�s2��V�HI'D�9'	R_̓I%L�w�\��U��g�o������!;H��d�Ň�m`7"O������N���D<��l����N���i!Ď�HCz����8�Q>˓?��$0v���� C�7R�R؆ȓL�.��u���v� �Ȏ,#9�	�'VR����	 ?����I�6�2}bT�4�
�{�O������d	*��hS��=�%s5B�AP�w�D�M�а��'"��Oǝ}Qf�7�T�YK`���������*�S?Ct4�0���d���1�̕�X(�B�IA��Z`cP)2��a¦a�95�����N�����ӵw���@�@D�I&
Bz�C��.70��ʴ8d5��P5��ix�BV�!��<�Ԥr��q��'X��a*U�HFx�d:-��KJ&(��ؒ?\0��	7]��-���)�!�@/hjX�Ɂ!"Vq9���x�ў0"�ۅFpR@�iD;$��
R+�v�-�P��Py-ߔS,{���u{�����?Ya%³q�pa�g.}��)�-�D��4fѪ}�	X�a��NB�	K¾hj��ˎ0ӄ�1q.�Q4*�7]|��欏�v����I&0�q���[�dy�c��Kr���)mL�Q�� p�T�
��?@|nA�%!ԸI��5$��Y%kJ�z�����X���,%ʓM�^�	�+�O�v� ��cCk�65���ϥA�Ʃ`��A�yb��j
e��J��-�&��w!]�a ǢV,�P�Tk�<E��{��2@�O>i�~:cV�#�:E�ȓ��)�d�
V�;��P�`b��%�0x��];�� ��	4S��|I6Ū�z�s'냝'8����-|��h�->-�C5e9z��4���V#����'`�q��H
`�ҹk�7J��d��gh�Y�F�H��ЁȖ�R3�:���aÕ�
�bU"On��bEX����F ��P���,S�<���_h�S��?�d�
��d��n�q� ��$�EE�<���D"02�[zZ���/L�2�f���+P��p=��N;��h4H�!8���I4�^}x��Y��=+ ��I��3���sPk�-m�DۇFC��yҍ�My2�x�M�-y���#ϔ��y��,�e�w@
��HSJ �y��N1\�RѲ�+�� rU;���y2o��{%IQ��ĉ#Y(�
���y2���m���Ƒ'��r6�A(�yb�ͪ��Ii�CN�*hF��y���!26����:�^���_��yҏ�7V�0���"<>�����yNA
E�p9[GE���X��Ѭ�y��fyj������������y
� x�:��UEBXS(��%f�A[C"O�i���0t����
7�9��"O,�9w��a~��1���7.��S"O����E�kA��02���hj���"OF�yC�O��@����i2 �b"O��)�$ӿ8�Lh��)Τ�v8)'"O�pQ��>P��-P���v� ]r�"O���5��{R���(�*�Г"O
iE��1��L=(n� ��"O��'c	"����E�(S�`"OZ� �ɥa�금�Z'8��aH�"O�!����8�p
׃R�G�B(��"O������<#צQA���x�|e! "O�ux�oߍ�.=�t
@�҅1�"O���ѦC>b2���I� ���+0"Od9��M�faSëQ3AvP�U"O�Y�7��M�P��ɗ!cHFفG"O�mz�IZ�hab��'H,���"O������?xP�;�$�~0X�V"Oh�+5��& ��=iƪ�;��!�"O�Q�L�&S�H ��pC�-"OP���1 8a�TM�DVqa'"O~����Œ�@!��˺2;^���"O*\!���(l�h��6D�]F~
r"Ox�'�3�ƌ�a�϶?$zDi�"OХ�!B��@$#���ΩH�"O�ЂvC���#f��2R��Ա�"O�z��K�g Ir���0���"OH�c� �$F�FE+�\<`�Px��"O ��&��'��dT T���ӣ"O"�K�#������C
�0x��)�"O����ō?!��z�L�v��iʰ"O� �)w��p2s�F���,��"O`,AtJ�s�fX�e�؎D���"O�Q��'���R�J`�q�"O����Ĕu�B����' ��xQ"O���eD�M��|r�$_W�S�"Oj|e�CT��L�0ZQ�83"OF!�R��ba�=���Ӛ=율�w"O01�a�Ϟ�Q���X�-�2�k�"O�-jpف/�����L��&AD 0!"O^�PE�(,j��Eʑ�qZ�cS"O�	���m ;���gJ�p"O�l�j��76�#�ǌ�^����"OƈQ�KG�8�Rw� z����D"O���͌=���)�Rh��"OjtY`푠Fb�i��<Mn�!�"O6�B���Ij�	C:R_��3u"O b���-���a�BXP�"O�h(����'` ���W3�x��"O�a8�D�N4�<����5N.��"O��0��
�/�0��-M�7
Rl;�"O��;����]�H�갫ʿI�ԌA�"OHH��D��=@y�ə�`��9q�"O��#2�$H^i���#ZZ����"O�l7K̝L�3�DTF���A"O��3&a�4�&I��$��9����5"O%ۖ(��kF:�7�Y՘��"OPU�t���d!�,ϔC����"OV�G¨x&�z뎶k�`PH�"OxTr�<x���z��Q<A~r��G"O:�e� �jlj�Ɗ�S�b$	G"OD����r�R(��dҎG��A�'&�y0�X�r��y�����o�~�E���)T��5 ��� j�P0�Q/*�t��E����k�"OPm�^�F�����ʰ�Qˑ"O*�ki�Eپ�ա�4ug"O�ze��0B:� �t�g0��"O�k'hU,�*H�e��O*�1 "OX�5̃�+bl�aB�A�p%�He"OH,���Wa۳O�4*vX��"O*;��D<_ |`֭Y/��E�"O�ضd�+\��c��Z���9��"O֭���ƈm*,�d��7�nt��"O�I�r�Y�-��H�#,�Ӫ,	1"OP����S^H�)C*C�G̲ ��"O@�D Aff�Z�������S�'5�Q-�2��ԃN�Ʊ���O>�����3]N9��y����c�=�Į�а)c���%(|%1� ����I�KQʧv������t.B�%�7N9\fX��hW!� 0Xa��y�@ƥ<�t!������ �EŊ�pP!D�|���S�D�$�dS�O��\+k�̫��Oy�3�"���= p�T1w|��˩O�� 5�A+����s�N>ݢ�.O,c�<�(!���6����c�e���u�ا$��[�ƴ<E��?i�B���L�aN��H$!�1j;P��FĈX�Fy��>%>O�ΞuC��г���6Ԍtb���1
��N(�S��Ms��ߤUO�m�����wG��s��S�<�AG�"���Pa]�jl5�D�<��� %3�hda�6hn(4����|�<a�� N�m:�K�6�D\�$JQv�<���%<8;��4�ș$er�<P��	^�r� C�UB�B�z��j�<�#�7Gu
�\�OB��r�L�g�<y KO�b��U1�K� X��Ȃ�d�<	G�~�ܸ@,_�} ���GCb�<�a/�z0R�6
��h"� �V�i�<i��i�tA;d��Rt�B�g�<�p �?:�J��%u��"�·I�<�����$R���<�� pS'C�<d�WlQ�q�%��&�т�F�<���2w��$+ch�	H��0U�n�<�&�"�,���I�0D���-�m�<�v �%7�e�DX�<�(�M�<y�36>�`��*��4��$��gT�<1/@�q��p�L
>��Z�
R�<��l"��P��
��0���O�<f�65r���3��X�d�<�`4m�D�iZ�7�nl�V`�Y�<Y��_;X�r�b�_�M����!z�<	FQ������C11&�3��t�<Q�H�Ft�,ц�� \���c��W�<�ĵxq(�k5�N#v��[r��T�<��� ��D	C�8v�����PM�<�蔋@ Bi�v��2��0��`�F�<�p��,�����eN�z�
�]�<�DnTO- <�Tg����%�n�<�1�%@T��u@ϟX�B�4D�t�<��dƥ(����jݗk6Iba�YG�<�/_5�LtٔFUV�Vh�u/�h�<q�JL�[�4��bgNw9*H�r�f�<��"�pPx�#��6|Z��f�<y�$`ɧG�	TdX#Fm��&GC�	�H���a��"|,��u�V�!h�B�N��i����7�H-X�BT`��B�	�Jڙ��)�>{z<*��\�b�B�	���y;��ώ���p�؆h2B�r�ȔC @�G������V�8C�I����5�@B��X`#/�C�&��Yy�ќ!���j�nZ�6B�)� ��A�+� ,�tz���*��e�2"O�= �j�*y/^1zSB��,�Iu"O$���$T��yGǪ7��iR1"O�lJE�8fY��E�A��x�"O*�S�h�0r���#�-ն\���2�"O�eYW����[�@�谹�"O���p҅j%�Ask��r"~=�"Op�4D�-Z�ri)#��)=��(q"O�e�b�6�4H�P��JW"O~t�p�J�`:�G[?)���7"O���%�[l�3 HT��n\#�"O�[օ<$0�p�#)�(w���F"O�{bNݤX�*] T�V"v�5a�"Oƭ���ˎ~h�Q!!��Ш�s�"O�у�'�@O��� ƌ�Q�p¡"O$�@ ��4�p�i�d�C'P���"O��䛥!�,�!D�f�,݁�"O.���A�C1VB�)6%��"O��҂C�37h���߬R5F4�6�4D�8��
W�=#Dmk�A=pr���4�4D�\��b�?lv�g��A��R�=D��8���)Y� ��- YVe�O;D�d�w�Y�ІP2��*`��Jg�%D�h!�(I�4d�C��J5j�sB9D��;�J��N!`�*0*�F�!�4D�$��-�0 q���"͆2U�X<2��2D��A�Ǌ�P�Ӧ�Ĝ9�U�2D�t
���I� ��;jZ©2D���ਆ�U�cW'_K��px�H1D�xK��1t�a���Z�g��d�U�-D���VG�#/+Y��(�f�t���',D�`��!"�X�o�o��3s�(D��!�Ԏg�	�i߆\��H��#D�*�j�:56x�9#��/G��!2� D����鈂S���:�J��>TP?D��0u�@�s���h�@�8J�4��n'D���P�2p�,�$�ɍ(�ihw	&D�\R"-^�9����,�/w��y��0D�<��BH68��5E��+l�6�,D��(��D8�����
[A�A`�$)D�|J�m�$TZԃ0�M`�h���*D�@!2H� tT��ҁo�3-
P�p��<D��C�ȅR�D��@�$�^��=D��Cf��>0`���oVI�,��ă9D���R�zH�ݘ�bV:,Z
H�$#D���#�P�5���I�f�yC"� D�� ��-�xYÒ�)V+����?D� ��.D2L>~0�	�t��lI��=D��$����)Ӕ%A��!��.D��@	a쐍�щ̙Ld��Ʌ/+D����bW�76���I^E~�9��)D�L��i�v�4j�3�B�3sl<D���pKI�[ $ݱ�(Zi� 0�Q�-D�L�bܳ�Px�B�`B�6�,D�[#��?\F��Y��ܣ@��i��/D���mӖH��I����qW���q";D�P��.AU�L���Q�g:r�ҳ#7D��@v#�z�f�"���!�@@�'4D��Pb��� 닚Ah�8�d=D�Pi1���1�j΀L~��@�5D�4bd�|��b'�f��V�(D�|�v��p(�K��@�~��x���$D�� U �h�0x��k������>D�,�œ�>�X��T�]�Z�:�k'D�� �4�FfW�Gb�q�P�6�~�"O���A%r" �Io�ȭ��"O@�@����Y����`IݷL�Fl��"O�x:���5V��xi�!�FP��0c"O��tB��{VcG�
?Q:��B�"O� U�X�I^Aڑ/���}[�"O��S�M�WR����m��
�If"O����b��R$��7�TG"OJ-r ��X���㨛�>I�C"O������'g�$H`j�:]�P ��"O�9�`��0��d� *��\"�"OF}{�`D�KF��B(ˊb��`9#"O�����V, �����l���ea�"Ot��taXiN���D�|��"O^��Q��6�:1�m��P��`�c"O��BvF007�$д��S���a*O�̰D��_(��A�ř��� �'�t�x�Fʛ��4#.E�NH!�
�'1�Q�%I�b3�/L*2�vT�	�';����3:�q#EL�5��!��'[���԰\�<�+�C�1�����'됴c�䛖?v��5D1q�hk
�'E�@'�CK�8��^2%>�{	�'����,
�REQ�,ϣ�LX+	�'%ҬSA���!�R�Bf����H�	�'�R����:CFe#V��LE��'�z5�u��3\*����I5���x�'\���M��)4�����4` ��'N<��K��K�Y E/�+_�͒�'	���WZ�H�d�^%Ge�@�']�6$/Z4�KWc׿�((��' ��H�J.!H���FH��>h��'4��m� ���~"�9�'��t�DC�{�&�p��D��j	�'ǀ5#�/��hph(��L-*���'`p���j�>����ޠ�0�*	�'����"Y %z3�ㆁ����'Sp����"E�8��0F\�x?*lK�']�m!���RT��w��#B��'5n|�d�2N� ��1�H��p�'��ũ�C�lX��Q
�k�'�Q�#� u,`A���(p Z5��'	
�!��G�$#��)�'��j���
�'Kr*��N�̘0�p>��y	�'��D`Ӏ�l0\���m�����'Ry
Ug�F�؛F���j��49
�'�B��%*��M�8��fZ�2� �	�'H����V�r��ȣ��^!+�.�8	�'W2В"Ǔ�X��@��(&xpɫ�'���8p�׀W�b; ω�����'����q�P����Ȓ�S<�		�' �U��A\+�1�7".Z!�5��'��a$̒I�b�����GQDu8�'8I�G�k�Je�d*[�T �Q"�'���0�ꋘ\E�l�S&�G;��!�'���S�	�/�1Y�
ӥD|xd��'.d���,ڮ/�I��g9Rܲ	�'�R���>L�� 3+Z7*)i	�'r�B�hUJЙb�ʏUz�Pp�'3l�`��	ht|���N�G��	�'��p1��D�!(�QJكE9�e��'
4�©�9"��,X�'��]��'�6P�H��
"��@��%����'�hp�ŲP��� ,�
������ P �b�A8�=���� O���@"O����W&�x���~B(H�"Of� f��hz@���凈9�ݛe"O�q!����`R�IQ�5'�I�4"OHـ�/@�vIͻ��L!)��)A"O�Eh0��=����%g��a��]�a"O���Z�F����%FT;�j�K�"O	��(0�ڴ�_���"O��j��mir�c�C͗����"O�xB�`""���50��A"O�M�Řb{�y�é#m�T�"O>�� Y,l�VA�6�[�s�$�"O.-�� �p="�"Ҩ߶[�^	�r"OJ`S��% ue\Ӧ}��"Ovi�	�a� qYE�Fˈ0�""O
E�P��ti{u��.s���d"O�)�"�G
LҌ<��$ٲd�z|��"O���u� ����s$[�3�mf"Ohi��.�54�j��B�.0��؃"O��V/U�i�Btb�K�B(0Xy"O�PE'�;E��`���85#rp(D"Ob4{QJ	9||�E�΀���p"O�1 ����؄L��B3v��`�"O(��F��H�J����$\���""OZ ����,�,<s�ш�2�Q�"O���"�=V��I6���f9"��"O�)��n�fv�R榘�.Y3"Or�b��@l&e����2��K!"O@�ҕ   ��     Z  �  �  A*  �5  �A  RM  �X  �d  p  s{  �  �  �  ��  *�  ��  ��  �  Q�  ��  ��  !�  e�  ��  d�  ��  m � > � n  �& - f3 9: �@ JG �Q L[ �a �j �s �z -� m� m�  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R��'��:�aɤ,��`vcء|�~Id�=D��Q��ˌE��z%O/Fs�mQ�7��)�S�'XM0�UhR: t�3��UU\`1�ȓ���q���*T <Ia�?c�ؠ��3�� �W���TCԺ����d7�-{G�0R�
Ը��̳c����N
��
����J��8�2qz�=��wYu���'R��r����e�4݅�u?��+Qœ�M@\
1�W�1�؅�h�eI�*�~UZD�����ą�T���Q�dD������(m��ȓ	��Rr+���<�Aj3\�Q��I�}Ru��4y�v��`E��2�b��ȓ2�,a양^�d� �N>Bņ�Q����$�Go 4� ��@>j�ȓZ�X��%G�,�Xd��غ"t�5��W# Ct`�A���X#��rg�-�ȓnV�yC�U���x6k�[K*��ȓQ^@d�p����sVl݁oVr���b2X�3SMD�=f8a!���t�ȓ0����I�<�XXC�
�Q;���ȓ�"��w��7+�dȘu�ȷ���ȓ;Ҧ ��B��IT��(��D�꽅ȓ9قu1�f�y_t ���7v��P�~- Q&�Y�F4���-wq�(��@֚,@�ϔ.���V�`'p܇�l;��GD8!�,�w-J*�هȓ5��S5!O�tk���f�<z6�ȓ~t�i1C�M)><)��EJM��{�R} �L�j
�*3ѢM%r�ȓ"��\��o_�4�WbD(l��@����<��;-o��P��&>�����C �3�^�A� ۤO��X���ts�*R)G 0�pHb:�H��?y
ӓA��Pq�*K<T��@e.�'�r5�ƓydI��C� uj���� �A���'7�	P!H�a�������far���'?(��]0:|��F��6��
�'"2���a܋,��aCN��
lL�	�'�҆�;V1�@&� |��TP�'0���"#�"�d��e���'xv%;	�'��$�߸s-V�!K�I�����'i�}�# )�j̓��_�@2< ��'��p`��
(两j��0=l��'Z��)�� �K��{S�L�@�u��'�J�#��D3.��i���ՋlG�
�'�x��&d�0:Ȗq�f&I�a�fԳ�'�\1Z�M���h #L�	a�9a
�'����'�<�,��#��I�*(h	�'�X��7gNa]r(Kr��F^���'-����;�t��*ԑ6Y0���'���t䖓e����FD�y��X�'È�r��4f�� Yu�
~�Hq��'�$3`�W��б�1b����C�<�AW�Zo�h�5˞1M�xS��z�<����6 x�y�� <�|���d~�<��"J w��@Z?&�HP뇦^z�<�0!%B/���� ��X�'��n�<�DD��c����-�{���1�E�<����;-i���g��n&�pT��H�<)f�<ؠ�h�s���sb\F�<!ң)]ݬ1A�m�$gn��P ��f�<� L0�i�3:���b1o��O��郢"O�A��M��]��8�-k�l�v"Ort��
D8g�\T��̜�f?���"O|��V$�9m���a��%
6�ɱ"O�Ī��$$���2���D�l��"O��)�ce<H=b$ٲ+�� �"O����Ο�t+���%�5}ò�ڗ"O��4��M��A�#J��t���(0"O����*ٗcJ��p��d���s"O
�5����6�h8Wo���"O��A�&Jt�H*�%�"j8	��"Of�->5���Th�hC""O��w/�p L��g�
M�$� "O>�`U��c����g̈7�v|x"OƜ�� :�)�k��E���"O$��0��<,��H=�� R""OX ���9^�H\h`Ȝ4��xIP"O���!�Y5�`��D	�6��V"Oй���X"	"m��AI���"OV��Z�SA�!�Bs��"OМ(�F�����*<���x�"OΩ�X�ޙ�4gW*���Id$PU�<�V�O�~�	�d(	�3Ѱ�Ɂ k�<vCʚQ��ݛyu�#Ak�i�<���<&�8a���yf!0���@�<yG�t���b
�S��U�<V�['g�Ȝ
 ��Z̐��FT�<�Rɝ<Gt$�#͈[Wꭢw�v�<��G%)�޽�5�ϊj��ⱍ	v�<y��0E����i�{��pZ��s�<Q�W {�j��B��y�>(aFU�<��Ɩ�5�"D!������ÊW�<YGF�y{��0���8�ɡ�i�<YU��%"
Й B<!db�hD�e�<���;1A��ӑ�ɸ�@ݓ�JI�<!��Z2q�@�D�$I���p�<���
�T'�ٓ�Î,B똙��N�i�<�	A�sP��Sũd4����y�<! �v����L'��5���O�<q����BB���j�v�"a�K�<��#À:�Z`��dݙR
RIȕH�<�e���#��8� ,��`q6��A�<Y"ݧS�i{v
�D.t�B�NA�<!2��>$R8�'Qx���
��W�<IB�֏}�j9�X?f���JB�Q�<��ȏ%ҭ���O�d,�Xc�r�<�e˔.ta�'��!HvZ	��S�<QP�_�K�B-�W!ٝcD�y��GL�<�7���v'ĝ�%�ΩGwRB�	Pd"Lq�J�H���k"�� :��D�[Ԝ�yP�8v�T��:x�!�$�'9]�a qHС84]㷯G�	�!��[��� �fK�56Ͳ���H�!�$�����P������p��܇r}!��50cX ��!�=;	��ZUM�g!�D�%!Z�u�����)ԭ��>�!�D� w#&4��ȯ�t��D��!�$��]���ȵF�? ��ٺE@S<!�d��Qj�%�E��(f� اF��X!��	O��C�A�]i��q�H�<�Wg"��u�ͅg:�T��g�o�<qGO�1�؃D
߷2�=���j�<�b�l�N�L4`B�Uç(�f�<��Ά�!�������8XN� mH�<� �s���Z|Ä�R?T���"Od�ڳhL�,n��֮	&V�&<pW"OX��@�3�����n�,T�Bw"O���w,K�]�P@Q�,жx�2�PG"O^�B��D�L}�,>����s�'���'��'�R�'���'���'��Y�̊b��D"a��?�@a#�'���'��'��'��'���'�F����)�� 	�!�3r,|��2�'�b�'"��'Dr�'���'&��'� x*4m�<$��B�i3�'���'4B�'t��'2��'���'=��I���B��q	�-����M)1�'1��'���'tB�'���'���'?r�
c�KX�<��k��:��M�'�'���'��'E��'���'���'����g�6m��@��եO�A[E�'��'`��'�"�'[��'��'I�0�� �w;T�S�+��I)���'b�'���'�B�'-��'#b�'�m� \<~=3�
;��c�'/�'U��'W��'���'���'!f��HU�1��}��c_:�~���'���'!B�'W��'���'���'�ˆFQ��Y��L@�8�n!�e�'W�'���'�"�'���'���'Y6���NL-+�V�z�ɑ���#��'���'���'+�'�"�'�b�'�\sD�&d�c�\�e�l��'+2�'���'7�'���|Ӕ���Oҹ��ܽ�6	iT�S]!b< ��Ky2�'h�)�3?Q�iTе���z��,�d,����,�C����d����?��<���}��i�
�b��\���یJ�4�����?9��Ѫ�M��O6�.��N?����\ ��Ȩ��͞3�p�+Ql<�ޟ��'4�>�-F0�l홗M�rXP٘��Z��M�&�m���Oc�7=�\�{��͝Z���O��8�2&��OX�d~��ԧ�O��D�T�i�󤙑D�D�y�,W��y����v���e��z�g)�=�'�?�A,îu@�,k�^%l�p�`����<Q/O��O\�mZ#7�(c�����	��[���z��h�n�����ݟ���<y�O��`0��$�Ȕ;��Mol�}Z�����	�J�z$���(�J����ߟ|9�
 OD��4@��Z�&�Wy_���)��<	d��Y�0|+F��=$��xpr��<��i��X��O�-m�}��|��kĿ�ޘ��-p� I��+��<����?���A2f���4��$>���'�hacG
�u# ���۠"�]�D�6��|�*O���H�.��Eu��YR+BT]*Mᄞ�48ڴ(u�q�<A��d��s�]�D��:L��(�K%A����?���yr�&zs�T
� �y� x ��R��$Z�BQ�������U&���?i�o*}�gy�� �&�Ƞb�1V��/�1+"\�\�'*�'S|6-V6c�Z�:���#�ڇg�D����6s^���U�?��<��?)��L;�b��Jr�=�Ƅ�)��y��_��M[�O��$�����)g�����h)<a�6��7�TP��i�D�IFyRQ�"~��n�?b�� w��" ,�	�S"f̓�ƣ����$�¦$������q����2�)�@��0�O�<�O��D�O��ΓL�66�9?a�� �G��~�P!�VǞ#R�訉@�Ox��4����?qTa��:��Ab�/�h<n|�WA��<�K>�u�i�ꀺ�y2_>ia���b�"MbC��\F~�D�"?1V�����|ϓ��O�� 	B	L,C�T,�f`E8I2�1��'@LPJ�M����4��������O����I!H$�q��;"�R\�5l�O��Of���O1������H�+�N���6�LT9դ�
i�`���'��keӜ⟠3�O�0mڣ!tz�x�N��Br �i5���,Z�Rڴ�?�iS�M��O^<��� ��H?)8&!_� U���q��2���bs�Ȗ'zb�'G��'/"�'��Ӏt�>$��ň&h8x֙��fґ�Md��?A��?YH~Z��Y���w[���gg�*N����2J��tM� ��|�,�l�w�)��]e��l��<yW�^�J۔$���ƇU�u����<��-�"mv��W7�䓂�4����
2�\a��d
�d�d�i'j�e�6���O:�$�O0˓l*��
���'���kx�i!�$K]QST@LS��O���'2h7F��q%��J��]�u�``QkP�L���1�h'?��DY |��*`��]�'d���D���?�!�&E*8"���$��9r���?���?Y��?�����O��RT�=Ft>��d-[�Abfh���OoځT�u��̟`�4���y�OFW�"�S������92EƠ�yB�b�V�n���y��㦍�'��(B���?q��ڿ`	h��f�*	[3х��e*�'\�i>���ϟ��IßH���}�$�r��u�$�j�N�j����'�7�
:n��O`�d+�I�O(�`�ǹ}�L!�@+�R��J�Q}b�i��mJ�)�&��Q�P?������K�H�%��`A'!9?�ta4;����D2����dX�dx��>6��\�4jZ�f��$�O���O �4��ʓ��F�
�� �p� t�E��z�̘ �I��yb�aӲ��O��m���M�d�i/��jfnș;�Z�A�8���vMWL����O���#�H?o1�����{�v�N�� ���AL�Fy`ek��תRdnH2O���O����O0�d�O��?icFkK�M�ѡe�,���{�\����	ޟ�P�4'V��'�?	��i(�'�0\c��>Zv$jU���x� Ȓfn#����	��|:���M�O�ax��Cb�\]�`*غd�֭��ǔzRt@�� �O ʓ�?����?���./�e��\��	2�G�6{�H�p��?i/Od�o��3Y������(���?=��5��T���@"Y6�T�bT�0|P�n��I�M�ӱi�lO�Ӊ.��E���n��x��'g�6��B�ؒ5p���&M�Gy�O]����2_�'10r'��;84`�̆.cՌTy��'aB�'�b���O��I��M��T�)*�]��ӗC1�8�R�RLPxP���?�ƳiW�O��'ئ6��;�t@{�� N_X5r��E�Q:ʱo���M[���M;�OjL��d�����<��e����LϺ}�|5�r���yBZ�\�	ߟ���L�	��P�Oז@�F��$|
h)2k��N���07)o�6Ԩ���O`���O��I�|��^w��wG�h��֙	D��@�9H�P�sd�Oh7��q�)�	��4�07mg��XW�[�rh�Ss@J�i�^t�v!q��*w�<7��G�	~y��'��
dڹ�p�*����p O.Aj��'���'T�ɚ�MctF��?���?I�B�TZ4 ���	�i� ��s���?AM>I�]����4
���3�$O�T���d�����X8V{�	w��cb��p�l�$?�C��'�l��I,,Q$Hi )H��3���RMX0�I��0�	�d��x�O�"�*e1��q�ǚ�-�
 #o��n"�y�Tx*���O��������J�i���4��+y�5j�f�\F�<`����L�I���ݴi��uڴ����./Z"���'��X�/>2,�wC�{���.9�D�<A��?���?����?a�.($R iB��xT�������Iڦ��/��h�	џ($?a�	�J6���� ��L��Pb��)�Pd��OH�l��Ms�x���h��gPAcdC�$���#q-(��<)1U� �	�H��J3�'Ђ %���'��L��l��F�\���iə��\��'�B�'�����t_����4d/���,.��z4��{Dy����w�V��k����d�h}RE|�^qo��M3��;[ϊ�e�ڿ�Q�X��9QR���-�'�bͲ�O�?q1r����wk*�1�)=C����gD����'�r�'/��'?�'Z��T!���7B5�Ű�*�f1ۖ��<i��͠�a��d�'� 6M#���s��p���r����.��M�=$���ݴ@���Ok���b�i��$@��)6\���h�fU�q���#�l�:Q�I�f/����?q��?���d�H#͒��2�S5W�1 Ql�O��$�<��iKFD:�'*"�'�哣>[�I��ªTQn�ze���	L����ş�m���S��)#F�F���	��w�bbƇ��x��Qj���7� ��_��:>�"O�o�I�B�|��򁀓B'�0����:H ��I����؟��)�My��v�l	�U���|, w�U�5=�a��J�N˓z����Tm}b�h���jM���,Ð��8N�1���ix�4g5��4���Ó��<��'4�˓Y��{0K�;I����@́\m 8ϓ���O
���Ov�d�OP���|��;6N<�R�F<�����-+��-/gC��'�����'��7=ﰤ1���4�����Tް}Ғ
�ڦ���4;f���O�~0���i�����F�z �ƸO&��rT��<��ĩq@����K�2�OP��?Y��V>xx��ѫ
2�x��'%������?	��?�(O�nZ=dD��ǟ��	�'�D%����bZ�yǊ��x�̸�?��_�$��4����=�$�2��0IQ �J�L�#A�m���9��zF
(�~�&?]Z��'�~���y�b� �g�����N�6R�la��؟<��런��^�O.Ҁ`2:�ڒ�M:�u�0�ιO��e��s��O"�KҦ��?ͻ5_�,a�GZS~�+%A��.��A�F��F�j�ZElZ�ƴ�o�A~�*��C"-��%*	Ô�\,n	�7Aí[
��AS�|�Q�P�I�L��ȟ|�	۟8X��'K����Y�^���H�VyR�iӠ����O��D�O�����C�p��MȲC�?�fy����=*��'�ұi�O�O��WC�!e`t)tJ�;^:�Q��Ί��|�RR��(�eI9'b�
Y�IUyr�[Ol�ԣ���8��a��+��'�R�'��OW�I4�M[2i��?��l	&y���ǋ�9?fq�R���<Y�i��O�M�'3v6mB�uQ�4h,u
��8u���a�A�:�(��re2�Ms�O�<bD
�
1N5�������c�ɀ19��#�EJ��E0�2O����O���Oj���O2�?�a�m��}6���Я�:X��az�kZy2�'�7*����M{M>�������J4i�y�*���J��>����M�Ӻ����T�P�����oԓ�`1���ͦ8���d�?�d�a�'5�h'�D�'�"�'M��'D	!���b��F�i��'�2^�4�ݴ��I-Oh���|�S��1��� Wi��~
����SM~�>���i0�6mh�i>�ӗ=O6�Kt�Z�麼qPI�$�8��sEC=/�d	X �Ky��O�<�I:n�'���1d�c�(��{b�q��'B�'xB���O)�	�M��fW�+��d:B>1Ș0�5,$$@�����?�Q�i��O� �'�N6͛�+`�A��]�FȒ���ҤnZ��MS"�@��M��'^`C�j�(���|��)� Rh``�2m��hs�+?:ī�7O�˓�?��?���?a����3X��� ���Yc��SaC�d�o�8{<t�Iޟ��I]��ޟ�j���˄��2z(N%x�`ݫ]l�T�L�F�eӎ9$�b>-�p�¦�͓�Q�G�Y�:w�͢R♱{����zԪS3'�O��M>Y+On���O$ z�d�8'/�5��
M�ZTr���O��D�O��$�<��iB�{��'3ﬀ��&׾/�j ����v^B�za�dkyb�':�6��O^� 蜁#��]�C�T��H�ol�H͓i��xTL�mTI��·�?���T=+�KZպ�p�'&��p��Z�x0ZQ2�ז?`<���'���'�r�'~�>��I2L@ʉ#7�,:VŹ�bV���	�	)�M�M�*�?9�N��f�4�m;�mP,S��c�_/�$�Z>O�n�MK'�i�p�Ȧ�i��˼ ���\�%C�m�w�RTc�L����{D���y�����>�]�<�	ß@����������Ic�c��Da���H{H����TyR�ӔBW:O��d�O����d�{ؙ0
@�+Y��r3��CŌ��'�J6M��$�b>�� �K�a��IJ�k�^8�cI;+v���6+����`녱*����&[κK4�>ɔ�<�'��Xx�51���r6.�^���'���'��O��I�M��`�<Ʌ�-$���tO�5hv�D����<���i��O�ė'sR�i��-ϙ,f2�2aհV�D48am��(��Y;��i�I�Z�����Og�'y"���8 㝱np�dd�9�ԡ>O����O��d�OJ���O6�?�G�T:zNR`9��0jt��)�-7?���F�a����¦&���@,�?JHL�cI�m��I�v	�j��M�Ľ���'V�v�v���� 	ߣ3�t��$N���|�*��W�>4J�2�'�T��'��6M�<ͧ�?���?��&�1@��)(���
s�x�D���?�������m�#�x� �����O�%�w�@|�J�f�/c4>�h�O�̖'�i�1O�S�g5�x��k�N6 �d�V	4���xf��@���*?	����@�'V�Ӽ+���()#El�@�F��V�W��?1��?���?�|�-O��n��j`�[B��qo@�;
_�U�n��(&?٥�i��O��'Ǜ�D�0U�m�%�Wt�q��;PI�6��O�d`4�xӆ�,��z����OXѪu�U�+���S����	Ν ��u�"��?���?��?I���)�Pܨ�qD\�Z�r�B��%t��m�"~���ΟX�Ij�s�(�������[�U5ڥ���эmb��C�B "J�i]1O�O�D���i��$�e�(X�pa
(0^�R��ܗ4���ƕ ����y�˓	V��W�����r�ԣ{�H��G�\iĈ$�՟��	���	ry��xӰ�`���|�I)P}t1�Mǭb�d�i��
1A�4��?��X�����%�8@��۸,Gd�7c���L�d=?�!j���i~�a~��ۆ�'HL=�ɨu98�+5�q��W2]>�hR$�O����O.�D�O�}�)��H*N�l�)�q`�?Q'2��@қFe܆��� ��?�;Wy��G�ъ{S��9��(3,-�`�v�j�X�D��U�z6�=?YK1>2<�iY(~!�0�&fS�����!P��/O�ImZ^y�O#�'H��'�R-�=��}�0��%�챐�OԚ+���5�M���<����oZe�s�D�§_�B~T'��D�.���������j�4��Ş&
V���ĕ;AqP�K��8(q��:k�Ph�'���x��D����`W�@B�4��U?q9� ���;'� 2F/ޛ*���d�O0�d�O��4�`ʓ'���(��l�R�ُ��%�"������Ѝ�+D����⟬��O�mZ�M¼i8:]a񆐐TJ�H:0��X�hEٿ>��F��pѳ��	N_�d���1��׾8��	�P�N�N���8Oz���O����O����O��?]��>� �ಯ��?� ͒EnNş��Iȟ4hڴMl^�ͧ�?��i�'{U� ��04j�	S��1EN�q(�1�Ǧ����|�5�Fβ"�%?��(�Zd�@�JXa��I�&�x�A�O,Q(H>Q-O��O�d�Oځ�Ĩ^$:2xT�CE��O>B�i�A�OX��<)��iJ�tk��'"b�''�2h4��uM�`����"'��3��|��i56M����M<�'�z�㝪@w�TP���jT���@�8?���t�ߔ^6��'u�����<2Q�|��P� �@��6Z�`�ゥG�"�'r�'x��T^�x��4z���sa�z�M��Ԙ>�q�u�S�?��-����G}�t�$|��Z��c�Z�k �p���J,'��.f�A��i�"�ܟP��&��h����+?Y3��:Rr����HY]Ŵ-)&�A�<	-Ov��O����O����O��' xl���D�r��A����X!��iG$�hp�'���'񟮸nz�킒�]:A��c�߄D����6�MK�i��O�I����逼+��6l�X
�f��,���!"� GX&��U%o���K�"j�dB�	\y�O�R�ڜl8��K��92�h��h��f52�'���'����M�'�U��?I���?iEi��9�ݑr�\�R!^���'0�o��6�m��U'�lq��5_�� B MƑ	��g�o����.ldP��]z�d��zB��O,���Ae���AJM�&��P��ղv�8�����?����?����h�����P)vT���*? NH�*4���d����S#Dɟ �I��M���w����-�'�^	 N�3E�h�@�'z���eӤ�l�pA��mZ�<�q3�(:W��X�� ��1�)��sA�EZp%�/���<�'�?���?!���?!e� ��0Zf@�n�vA���H����ͦ�K/��d��ϟ4'?a�ɱ��@R��ۺ7ۈ4CgO�(JIҨOV�mZ�M��x�O��T�O"�Bʇ1ʐ�2� β`y� =a8|8x�O�e!��D�?��b9�$�<y��$G�
���_�E�:\P$ ��?9��?����?�'����e�&�V˟!㮐S.L��)VY����џ�Y�4��'>L�L��Jgӆ�mZ��B�$jߜ!(&����E�m�f�faK٦�Γ�?��mΌ*����~~"�O�) c��d�5��mRx9�.�y��'9b�'���'�r�	�52�F0Xč�ZBgbߨ+q����OX��m��n>��I�MKK>QQK(T�$���W�����H2$�'�D7M¦e�-9��l��<��%��9�a�f�8�H%M�jE\	#�%����䓌�4���$�OD��P��T��Lε1U���$��Yw"�$�O�ʓ0�����Vb�'��R>A"�*9�x"b�H"�FI�ѩ(?Y�T�H�ٴaI��j.�?ŉ�"�Ձ�ֿ;y�dIԢ�ubU�g�o�l���O��?��/�d�#��S
Z�D+�%���-9.��O��d�O`��<y'�im6��LF	bFH���@�4l��j���>�r�'R�6�>����x�����S9�&�;���Z�,�H���eٴ=�����4���g��{������_̜ ��
4(�xdH�ʖ�bb"�Iay��'���'�b�'%BZ>���ȗ�Gr�+d�
������Q��MS	��?a���?9I~j�9���w��Pf�E��P���5e��i���a���nZ>��Ş&�plZش�yR��|sR9�T+P����yr'��J���OybQ�������'�FtY�M }�) �S����r�'���'�"]����4g�4Xx-O��DO!V�n	�b$[�6.�A3k�WA��X��On mZ��M��x���U۔,�~����(����Y�������E0
/1�����/�ʢw��,�`B£(�ĝ��)@�L%4���O��D�O��,�)�Sf�9�*��2b-	�}K�M��ly���U��OFn,O���՟T��I��֟�<s=&M��Ń<����Ǯ+�l���Mw�iO�7���F��6�{���ɟ`Dx���O7&���
_�P�Daz���?�,���z�Ay�Ogb�'b�'��A4b_�m�G�E5*�����e�.��	��M�$k���d�O���d�Ҡ�k��� 6 ��ч��;+�9�'d6�˦	ϓ�H�~�(�K"�:9�B��(�y��C�~(��`㝟��t��v�B�g�JylY>u�L8�cH��=iw�1��'�B�'��O��	$�M�`���<aS��k����5�W`�����A��<QĹi��O�E�'�±igH7͕�
�P���;��@���#��퉳t�F�	̟�p�ݠ8�T�=?���տCЏ;n����B�/���1C�<����?����?���?Y��4��� �	���E0d�%�C	A��'u2p�t s3����E���%�8���2\��!�"$x��	��'�����f�j�p�	%"p�7�s���"_�Y�j��>�j���l�:��i0�M�`����M�	By�O�2�'b$vD�8��(��j�a	��'`"U�(�޴_8�+OL���|2���N!fX��
�'���:7�[~�F�>9�i��6��H�)r �=IAF,�0���G���^�R�B�!��1?�'/���$����rj��'�n�,��Ռ�-y����?!��?��Ş���Φx���y�'�Īb�F�"'�lJ�{ț��DTq}BO{�h��(ݝ >�F@։0�&9 cJ榉�۴R7����4�����
?R�H�'����Gb��,�:=�|rA�?f0��Xy��'���'&��'��^>�:�.A�p#dܸ$%ʟ��a$fź�M+d���?����?I�'��9Olnz���H�8�����+��ł3��!�?q�4YZɧ�R���ش�y�#��.��zP ��X����u�P�y���#%�	�_�'&��Ɵ��I�)sDh����+T����w�Y��՟x�r�̟��'�6D�Y�Nʓ�?��I�:��Z��ל+P�*� Ķ�?�+O���By��'��� %��%����U�)1>�8�	̜h����OJ���#ʵ����f����j4����g�0�9�QaƦ���H�����������	̟�G�t�'�`���gX�G@IC��Iq2���%�'>�7��5.)���O��lO�Ӽ�R	Q3T��)�E��o7�Ik2���<A��ie�6�ͦ�������'�ht����?j�h�Dg`�k��5�҈`��'���h�Iꟼ��՟��I�OZ�OW�|��p
�b�p�')�7܈9*�D�O��$-�9Ox\����:X�d&	"i�/�F}��b�Rl���S�'0�����*K8t"��O�Z�ph��I����'��e�M�ޟda��|B]��b2��=ir�P��?QI�i��F�����Iߟ�����Shy�r�.81��O>I���·o!����[9�|�����OXHl�r��<�I��M�C�i�&7��:"�`�hfd�;�Z�q��?�@٥�c����� Z 쁬uL���(?a�'Կ�Q��[q��a��[$)�pz�*�<���?����?���?q��mJ-q��� m)>�jp�E/)���'�R�`�U�15�X��ۦ�&���`k��N$�3̚�+��E�����%V�^<��O��	"s�i���)�� Ԅy�YO|�����3:p"��I�?��d>�$�<����?����?���mKp��fI$�pl��?����J��%b���|y"�'��	d����ߝ6�N�rgJԮ4<��`���M�'�i}�O�ӹ5˨�bEN�P@��+�ݑI���[3�k��x���ny�OC��	��'�t,�@��*h���9�LN�|$l���'��'�R�O���4�MK���:[��P�@�]��ǌD�(�T|�+O�@m���]�I��MK���+��K �R?�b�W���t[�F�cӶ�i��yӖ�)��Sa��|�-O�m�ʺ`h�)Rb�fr�Yp�1O���?���?����?	�����gG���1�!(�zSe�I搨lZ$ �d-��ğ��	@�s������k�E���J�g>���KF�V�vjѵi�
6��D�)�Ӳk�XqlZ�<YqR�e��Q@���y�h|c�N��<i����dǷ�䓔��O ��ѽ%މ�`�k�X�k��M�`V&���OH���O��@��F�Y��'�rm)G *�s�VW�����_'-��O��'�(7FئU9N<فHP8*.�(��Wd���CJ~2��8w��@,2w�OR����2:ES�r�8L���.�����(~�'n��'nR�՟ 
��
�&h���S��@�P}�ST�P��4Ul�y�'�X6�;�i�q(�A&6��xU�ہO�>M�$s��z�4_����s�:pQv�uӀ���y��K��4�N
�%V� U`�+=D(L�Tg�#����4���$�O����O���֣E���
 b��/��:AE��8��˓C���%��yr�'�R���'&�q8p�I�Qz�\s�خ!*D02G�>�շiq�7E�)擘`ZB )A�^�ZX�a�BR����H�a��v�!�Q��O���M>a(O�U6L'0AT"� �D��!�O����O����O�<��i��5��'�4 "g/U5@�,�#��Hr�B�'�H7m2�ɿ��P˦�c�4{���R�$&��BV��(��#M���3�i���B�6���OJq���NL�j��a�)�
ˤJ Nݵ ���O����O����O���'��_"��+��"����H��I���Ɍ�M�2c]~�"d�t�O�9
%����!p1��|~I����c�	��M����D��Is�撟�sT/��l&�@biZ8m���Jw�_�9���^�M�4<�d�<ͧ�?i��?��^"�j`��Дh(E�T�P�?I��������:Dl�(��ǟ\�OFLŰ���6 c�B;V0�!��O�X�'��7��A(H<�O�J�kt�P��ÕI��a%m/S�J�b���	>`��O�	5�?��3�d](^��8�j\Ėc��Q  ����O��$�OH��<y5�i� ���\u��b�gRVʠ �G�y��'"<7� �ɝ�����}�G�Ǜ]�Dd84��kOjM8��'�M[��inR���i���]YD0��O[�\����.Ց[V�p򁠗�2_"H͓����O���Ot���O<���|򖠏7o��d#KT!bNz�"�i�)M;��E lFr�'(���d�'q*7=�<e��dd=\т�)C3��l+�������4U����O( B��i �;j=��42k�XQ���5���1�$��/�^�O���|j�HM�T�t��4LA8�a�
 3��i���?����?A*O��n�NW�<�Iӟ���w���F��U3�	�E��4�}�?Y�Q���޴��v8�C�D$�@�-�`�`9��N��I36}`%�A��*�b>E���'�t��'>%�<��8�N�fCJ$��(�	㟸�I���	w�O�Bg�1{S&�q�Y]�����1}!d�dm������ߴ���yG�˦8��$�ӇD�S��U�F�Q�~"�''�FN|�����{�x�q�PK�(�(���]�Yq�9�D�^�GSv�r'����4�����O��$�O��dO�18��c���8G�y�&ʙ�u7~ʓ=ћ�+	��y��'�����F�$�;#j�&B���tm��
z�ɩ�M#�i��O����Z�Ӆax�b掍����gc�6l4����.+�	�m�j���'RV�%�ԕ'�����:���e�7l84���'�2�'����^�<��4'
�T���Y`=��4hS�"{S|d̓+{���D�]}��n�,AmZ�M���^@�c�A?5}�`r�J�Z��X ش��$�� �������O�G�Y�Q�f0�0��� K%`����y�'U��':R�'�"�IKD
x�LL�<Υ��� |��$�O��D���YX�f5?��i�rQ�D
t �ZZ�!:�C��Y��Y��D�&��M����o�H��Hl�l6�e�����@S�lk!�.HrR�QU��?}�M0�<��'UZ�}y�O,�'���A��6��%��hO��(��'�RX�D��4B8�Γ�?)�����Kn JN�/Q�Ԅ� ��I	������4�����O�����C�+%8�s"b������A�K�v�Q��������H�8��pF�Ox�3���Nr��A!�7J)F�E�O���O��$�O1�l�|r�&��O�>��FC�~B�p$MC1��E��O<�mZt��%q���Mc�e�3V���c��*/��i��N:Y���j�
��d�r�|�	۟��B`�C�dd.?���ʧPl��'�ě.lHi��<9-O���O��D�O��$�O�ʧOV8p&'J�Uܢ����ݎ�Nڦ�i��C�'b�'���y�Ev���dopy�	�HS��qU�(#JX��I����I>���?}���N��n��<� �<����N�ܨh��q�!rp2O�H��Ȋ�?awa?�d�<�'�?	�?2j*Lh@�N!t�x�c!c��?���?�����֦ys�0?�������F'S<�,i��ݿ2����C�>�e�i^7��n�I"Z�����s1�!kEÌ�I�v�I� 1W&�4 ���>?9��1��Ĝ=�?9���%�� z!A��ް�4�V�?���?	��?���i�O�1Ov,���ƌ��Y��`xr��O��mZF��A��f�4�0��ě4O�,�����B���s�8O�Loګ�MCd�iG���i���Od���<��D�1%��qB��.�l�"u�^֖�O`��|
��?a���?��aܔ@�f�x<}�4�9�X�/O�(mZ�S�������D�s�DR��ťP�ó���U�ָj�����@ަIPݴRL�����O���aڍ<�.� '��#�*���Ξ(4c�!�����$�={i������O��{"H����Q�i{*-�m[(�DmY��?9��?!��|Z.OԌo�Y1��	3!$R����*4�B&H9D*~�ɮ�MS�⎷>��ie7��Цq˥�32fV"��-L���;��
$�$l�Y~��\�*�p��SZ�'��Ѿb���G�N�Y��u���<!���?9��?y���?���d�/IR���p�JQ���'�?�yR�'��g���iӑ���ڴ��1���
��.b�
�N^!�"�@�xl}�`eoz>��� ��!�'d⍊���1t�;�P 8b��ïJŎ����3m�'��i>�����\��Y2|:��VNu�DC��r4`���T�'�7�����O��d�|brG�Ԉ��
Nyxq��LD~Bʶ>q��i��6M�F�)rc�/�p��%DՂE���)2
Ϳ56l��P8B@��4B�៨2��| j�C�F5�VLC4/��#��',B�'���4Z� �ٴ݂]�墕�.8*��Å�iO2��L�U~�fӬ�PکO�%oj����i��d����i��'2�P�޴9=���vl�f����L�2d��$�~BB��!�Ľ���T�6�~,��Ǝ�<(O����O����O��$�O˧7l��Ȓ$I�4���9�h	�'+,mX�i�~��V��	Z�'&��w��Y��CR�,)�=b��R�>�Ν� H|�4@n�
��S��".AӦq�B(0���!��!�(aj���Po�R@��O�yL>Y(O���OB`��`�v�xC�Ŏ
D�4��O����Op�D�<�Ĳi��I��S����c�(�:�iY�r�l�h�hG:^�I�?�R��ڴ"���3OT�0�ldqn�;y��|zww�L�'������#�����ԁ\؟P��'W�A����2�@c�N����r��'r�'�2�'�>A��+3�T�Ц�Y�T�̌3%��`(����M+�n���d�ڦ��?ͻ���� C��]mXZ��@�0"]ϓl1���m�0n��R�vs��F�b�a�O�|���)B)�h� ��/O�0 �!�Q�ny�O���'���'i:㢒:'�\ <��ŀ��<1B�i���ؤ]�d��C�SƟ(g×�\�.��w	L���P"E�P���������4H����O��X�$���7$Rh�UH+5���굪�L��y�O�MC���?Q �$���<���_
q����;PgF�Z$�'�B�'Z"����Y�x��4wb�)��:���a�/��@I咥c��0������~}Fj�Έn��M3#���]��A���G6%'(�	�G�;���۴���Ԟ$Z����'��Oe�@�{	��ud�Z�8W��j"��	��������П��IB�'�X!�gA���mzF�Ö}�r ���?9�FV��a��$ �I�M[L>Q C�u�jd�3#S L�2� &-32�'x�7����
Ux�ns~� FN��̑�,))W��Is/��O@����ݟ��b�|�_���� �I��x:�莰��(C��X�.�Ґ�G�����ay�eӊ��f�O�D�O~�'n�8�P��K�D5����%�=i}V��'�p�|�ƣqӄx&��'!'����h��b.��%5�`8r��0@����Wk~�O*�(�	�VU�'︈����2�y�
S�&� 8���'�"�'�b���O���*�M2튚M�x���!#z�����w�����?�p�i��O��'���D0{� �X�N�L:��m#`H�7M����A�ɚ����'��Z����?����-�3 ,L�X@ɀ*5��h�<O�˓�?����?���?�����)ߩ��U���^0�s���xhzUn��K�,��ǟ�	|�SǟdZ�����΃�x;�L�� Q��c5���(�)g��9$�b>���^ߦ�̓�h僧	1~�(@�!m��9͓z����ӧ�O��N>�+O�	�OrUy�D�=$�.��u	�+t���O��d�O��Ġ<�T�i�P����'��'��\���Ң�2���퟊A�Dh���k}��r��`n���ēF����7%�92:�1��jm5�'vdjca����� ��$��'�8hASȝ�WB����@���̓�'�b�']��'��>��	���
Km�N��gC���=�ɳ�M���)�?m~�"�o�q�Ӽ�A,�1��	���,@!��#���<A��ia�7�Ȧq�����-�'�FP��&��?2��������ڊW�����m�=h��'��i>�����d������3B����V8W�nux��ۋ/]�ɔ'�87�U�!�X���O��D<���O>��� �&Mf4�����Hђ�M�y}��x�^�m+��S�'
�<8� �!OK�.��!/ɱ
�<�+W�T���	�c��P'�'#~m%��'*��27%w���&��e~�dy��'+��'�R��dW���ܴJ 8J�����@ΑmL�|`C$�N��&�$KB}�f��o�M3e�
�P���^�<�Xz�J6��iߴ��DI�Qp~UI�'��O�_�DH��Ķ8��ݸFJ�wl���?����?a��?Y����O�Fu�q�Ы�p/�
߲� Y������M�����|���6�|���xc�%�"�S8ym!�NADJ�O�$a��i.t�6�(?Ap�W�6-zl��FM�s"�8��G���B�O�1O>�+O�i�O���O�����Lh:-���HB�����O&���<9b�i��s�'���' 哉v|&��̈́�a�c���[)��O�����M3��i��O�S��.Ls��A%-�D��
Ԓ:p炜(���p'?�'7R ����jn�B���^���(��"y�@����?����?)�S�'��D
֦���A�
)��1����GW�xa G-vTf���ݟ�ܴ��'.�J�V�C20��r�(0N���iȧh�86-�զaj&J��m̓�?�a��J�8�ɖU~"G�QwHK�F�{��,ñ
���y2W�����`��ԟ�I���Oo:��FI�J�"�b�Љ2p���e�QE��O����OȒ����L��睾xIDiw˚�2*�[�,U�4P�����M#B�|�����'@�#�4�y��cn��qI?��˃Nۖ�yR�����	�<��'��	韴�	*?�l��f,:v6�rP��	>cn���ş��I���'S 7�����D�O����
%�lM��1b���邞,�����OlHn��M�x���`7:P���\0�#)���y"��5�J�	�� 	�I2?!�'��D���?�ֈS��:M�v)�fm���FG�?���?9��?�����O��Ia�9�fY�C-��xY��ҷ��O6yl�`��Ea�6�'ɧy�LX�U^�,��:s뀗"�|)�'5Z6m^ۦ�2�4A�v݊�4��d�D���'%	����w�U	ReO5K=`yB��0���<ͧ�?���?����?�6!�6&�.q �%Jp�$�%c���\ۦH@x�H�Iџ�&?�ɊP2F���c�a�hQC!�q���a�Oto���M[%�x��T+�}�*8�dV!d�|�� N:V�إ�B�����^�t��g͚�Ox˓X��Lqq��/�H}���I$�Ό����?����?!��|:(O&5oP�D�	^s�A�A�Zܹ`G�]?扽�Mc�2J�>�P�iqr7mH���B��$��Yyf�ƹvX �#/��3`&�m�i~R�)|����p�'��6�K8,+�!�G
�XH�a�C��<���?����?y���?A����F�\b��*�̢@�"N����O�oڒ3(�zd���|��M�Q<(z���7�����	�>H��O��oڿ�M�' ��#ڴ��d��v*
���Я�X(���_lD�ȕ��?ё�%��<ͧ�?)���?��hѮ�. !�
����p�ئ�?�����H馥ʄAw�\��͟�Ou����"�M��t�����,0��O
��'��i% �O�S�K�Ĵb�hTҞ�P�d06���m%i�X\C�M0?ͧ_Ӱ�D� ��+,�y@�η�-yԉh��+��?����?��S�'��d�ǦI{�A�8y�� � �H(�88J��<���~����A}�Mo�@Tx�6k0h�#�E�1�<��"�Ŧ�ش+<R	q�4��dXjjl��'��S�s`�l��Ê�S��->Lɜ'��	ş �	̟8�I˟��N�4̓�K��퉑1*�Ȉ�Q�X6mi]��O��:�9O�-mz��+GC9r�
��	&���Ѷ����M+b�i� O1��sr�s���	��N�8��_�F4I��]�[�z�I�-�)���'�!'�0���t�'���� ��LѤ��d��<2��'r��'	R]���ڴa�m��?��f]����]�&�����ͫ%�%*�"�>���i�B7-�F�I1+Ŏ�x	� ��� C���2������"�_�z!*��$?��'7���	�?	$C�y�I��bφT�V䚐`͎�?���?Y���?����O��!2gFDU*��HE����S��Ov�o�2A�6�M����4�.���޵#d�C�鏭}�&<O,Uo���Mr�i�ܐE�i��D�O��ze��Ҥ-,:v��!��Ztɠq&Bt�P�D�<�-O�	�O����OL�D�O�t(�/� ;Q��@b�p3��<Q@�i&���'X�'L��a5�y��'D�A�G)Ȇnl���2y��V��/Pt�jٴ	���Z���O*�t�ҶtY�`��*���89��Ɣ�r����Ӌ�%���)w�j���L�Z�$�<�-On��@��^@��!��,��X����O�$�O��U�"�H��<9ƾi ��w�vt�'�G�,���hʞY�a�'*6��O���|�GQ�4��4Ư�Ig�Ez�"��eQ<0�H�UQ�|�rh�
WX6�c�4�	�O��t�OĢ�b��l�v��! B<#�]u�܇y4xU��?i���?����?�����?�F矪#��5;%�@<(F`@�%^K~��'�6M1,��O|oE��[W�M.|�����!܈�aI>	�4d/�v�O~���q�i����Oʴ`.ԫt%��K��%��C��K+sS�
�3!R�O��|z���?1�O�а@w�|�L��3BT(��@���?I.O��oڳv�Z��'y��O���K��]�|��c�6h�m���R�yb�'Qz����n�z�$��S�?� t�2,Ә��X ���3�Ը AeG�ªLp���'��	�?��`�'@�E%��[�H��2Ң`X�����	������	ȟ`��֟b>ŕ'�26�ϼ"���
@	�E�d��C��!w݄��������4��'�z�Q���T���o/c\|��0��,>6-Pզ�#�f�u�'��@��M�?���\$����$P�T`�����<��0O$˓�?���?���?i����I�p���K�
��.-&��m�<hmMg^��ş��	T�ş�K����pn$-szp(�Kӄ7.�dΙ=��i�~�O�O�`�
��i���Z>tY@A)a���.���+����W�I��
!��O���?!�Hi})]�f	���M;��,���X�	��x��]y"Mt� ��6O��d�O�0���>E��%� p�(�`,�	����ڦ}��4{�'���G�_جq١H�<<�t}9�O�YC�C�8:it肢�iߟ|Q��'���y(�8#~!�1	@zV��86�'���'�2�'��>��I�ch�1
rN�S�>����ܕZ��e�ɲ�M����?�� ʛ��4�l���_X̚� ?F14��23O��l3�M�ҿi��ɪӽiq�I�~0b���OJxX�w]>"xĀkC
��$��2��E��Uy�O�b�'C��'�	D� z(�
�E1j���]�w��	1�MK��>�?I��?1L~B��t.��&I*wD��r�	9�JU��W���4[���`4���N�@[���U�mª�A���9=6@����V�	$8�z 2 �'�0�&��'��-��MH�l��+
��5^�t�I���i>m�'�6�S�V���d~���j@�l>ru�B̘=�����M�?�W[�d��4ab��b�R)D��5�L%
bI�"��Z)P3��6m4?���V�[K��/��߁��nǟ0lp%I�mB^F��r����֟��ԟ��I۟x��概�}@�L�A۶"��8DЦ�?���?i��i�:%�̟plZ@�	�7�5��G}���KtĊ�GU2��H<	��i7=�n9�%gv�(�T鋀��=2�<�1�*L��g �>���#�䓇�4����O6�ē�u�^c��Y�9p��"
��t��d�O��
䛖g(L���'mrU>�R��,n�L�s�!R�:}�g&?1"W���ߴcțF�;�?�"��/&:I���p{�Yp�FW�!����e�S�N����|�c��O�՛H>��9v�8 �A7���2�[��?����?���?�|R(O$�m��_c 18sgL�TW��J@%T��|��#�CyR�`Ӯ��J(O��$�1h�%S��B��d�'���f6 ��]k�`Pܦ��'�IQeg��?M����0`�7�1kPEڲI�\��3O*˓�?����?!���?����	�U�-�ըŮK|��`S��XHn�n!�	ßH��Z�s�8������k��tNR�fm�k9�I҃���Ҵiɮ�O�O���i��Ę)y>x� t��*��4 C�Մ%�d�h������5�\�O���|���a�vXq�� 3����CdX�)� ���?	���?�(O6(lZY���	ş4�Ɍ�,@�E�?���s�HO�|H���?�F_��K۴j~���1�M� ?���$v��!�R�F���9Hz��ڱ����c>}�1�'����ɫ6I��آ 
<D���Q@��`����	ߟ���؟��Iz�O��M]�#fnH�DOA=2jY(�bCx���`Әp0S��$:�4���y�jl�|�Gw}�X
Ã�y҄gӂ�l���M�Ä��M��O�L���Q����-�.~���E��p��J� �O���|���?!��?��ux��`1��'BM��k҆P-}B�J-O��mZ�Y�h��I럀��c��̚���2�Z}Y��K"���3�K�9���O�1�4���OOl!bv��!X3hT�2�߳ Rm)"�X.
3:I��O�:W$ձ�?1�O&���<A��ǧT�qP��ӣLD����W5�?����?9���?ͧ��d�ߦ��V������$yK��@�ᑆ�O"t�����Mۉ�I�>�Ǻii6mX���٥�\�[�rh9��ςF�	�H�����n]~b�SYktI�|�'��;��by&x
VbJ�J5H #Q�<)��?���?��?!���kQ�cZe���
���J �
)k���'F2/i��,zw=�>����'�C����mtB]H��Z(��������t���w��)�3j��7*?���"�,Kbk�^0R���h�i�2
�O>��O>�*O�	�O(���O��7�ʓ,�|�Hv�ιg"�� �c�O4��<�U�i+H���'���'��j_z%i0G�:*U!"a@�e�P�x�I��M�f�iMO�0TަL�3�M+�l�i1�
�*C%f�DT�h1qj/?ͧ>���d֞��"����C�E� -�%�2E�? �<7�'?�'Mr���O�I �M#U(S+/+���N�	�-#�!\b[�����?	b�i-�O(l�'�6�����i����n=�M���%.w�	oZ�M�'��M��O����@ޕ�"H?	�gMMɒr�W�-��O?u���<A��?��?���?�*��Q�g.p&u�6�%5]2`��զM)��A� �Iş &?%�	��Mϻ	�*��Ӄ��R�1�A��>n4�&�i�~6-g�)���eo�<Qs�� ^ �0c�
��M*h̔�<��3z���$������4���$S�'�$�X�'	x����ݕH�r�d�O����O�˓{��H7�y��'�"j����(�>~�Bezc#H&H��O�0�'?�6���1M<� @��^�ty*�OB�-j��@�����X��<y1!1�ӏX��!��B�D�d~���^_An-�W%N��x��Ɵ������F���'�� Bs��8yt��ᦝ�[x�8���'{l6�Z:�I$�M���w�̭���H�h�ԫ]L*fc�'�7�Cͦ�b�4wp�ڴ��$���J�'�$!{���3�2y�&Eѥ6|	rn2���<�'�?1��?���?�c�'*��q*�o
�P�����(�9��$�ubWmm���Iן�$?牟z*�8rNJ����sȗ�S8ڬ��OZ�lZ<�M�f�x�����@��N8�1��1^HV��P����JI�¨z��r�O��Y,F���`Z?F�r�8���z�,1��?����?���|*O�}o�"���I�7��z̱7`$@CSF�H�I;�M[���>I�i7m�ʦ����3O���+ާ� U!W�1?d��l�R~2�\[�t�����O��ʀ40���V*b���(��Γ�?����?)��?����O�䠈&R�;.LS�KI�Om�	��'e"�'��6�H����O�l�~�I�M�� ɓ/��+�i��\@*u�L<��i<t7=�J4ʤo��.���IS�ǱK+*�����+��eh�P69�l�$���䓻�4�f���O����t�f�A-Z9n��q��O�)�j�D�O6��V"�(E���'��W>��Q. @�����8T��Yp2f)?y�S��z�4*?�F 0�?�I$�
 (f`	�.�C��A����D.�}��©0����|: �O��H>��(�@%S�h��v�޼���S
�?q��?����?�|Z.O�m�*^����UǁWS���'�B(f�LP��>?��i��OZ��'�V7�
K |ܓbm��)Ӗ�1vɥ�>�lZ�MS&��e}���'2���m��?%���� ��L�v ���ؿC
`���4OV��?���?A���?9����d��UFT��!!T/Y;um��7*����� ��p�s�p�������}ˎ�)��4T�~*�-���i>�O�O2��F([��y��DK��٥LW5�t��Ë��y�aL
]�vu�	8?9�'��i>%�I*�����i�z"��t�7T�D��I�x����'�L7�θO���O���99��5�w&[�R���Y<�����$�V}�i�r0m��ēzt��Ќ55\��i�)�/{(�<�'m�,ړ�P,[�R@��$�P�|��'��2F(FND�]�.�`_R����'�b�'��W�"|r�\R��&��>4JhJ/�9��N �/@����IԦe�?ͻw ��0w)�5��)�(�&�X��?y�4w�����"=�h+�O�5��º���"ȫx�"��u�[=
gN���.�OB��|���?���?��*a���ۥZ���)�� 8���+O�}o#CJ��ݟ���m�s�@�r����,��^Z�e�@�L���O|7M�D�)�	��i��P��2֐�ЅkK`<zЙ�f���	�,�zT���'0'�@�'�<U�1d�>����˗��Z��'�'F��'�����TW� cܴ,�������aj�؜"̱���{m��K�zݛ��$t}b'g�n�mZ��MS��A#dB�b�	WkZHU�D�`k&!�~Ҫ��R�Smܧ׿c7�Dh@��ʴNث&RjT*1���<���?���?���?	��4k�0h#N�OґPs��1ck�b�"�'�|�L�R�?��ܴ��K8X�ru!^0���C��>�$���x�fs�\Dnz>!ÖI��crh�I8 ���B�:N��d��N�/�0��W�A3D*$�dL�����4�����Ox�DL�[d`q�ɍ?E�D�#�)���d�O��u��Ɓ�����O{�̺���96*�����>>Q8��O�`�'�:6m[Ѧ�HI<�O������K���V#6��(H&�O�(2K��P���4�d`B��^�h�O�t�Íe���wŃ=@L�kRO�o�7����������d	�
-
Mð@˟h����MS�2F�>���i�p���hCV�R�B\�/�Vx��dj��l�$`Ĵ�J"?Y7`K40�f������R�(�㉃�#h���S$R�$h��<	ߓ�p�Ip-�&z|*����@	��i�B�t�'���'/�@lz�����5|�Ѹ5n�8Q��ɻ�����M���i6hO1��P{si�-\���^ي &c�o����R�D_4�d0e3Ѱ�+�֒O ���K	01��q�� jx�y�P��;�ax�i���ђ'�O|��Oh5�a�O�D��Q�q�L�cMt����7�ɻ�����ݲ޴2��'�i�s��g¢9��_��e`�O�E3R��0��1�?�iʱ�?���Ofy9�/J�\o>��Ӧ	(��C$"O��CL��4���>#��LzR��O8�l��f�^1�	ԟ���4���y�
T���Xz��߫G4LzG���yr�n�R�o���M��OT�R�)�'0J<rwFZ�?	:���d�:����?$D�bgl��5�'"�	͟@�����	����ɨ(����)�+Tڈ�:��7w��'�47�6���Ol�D5�9O�`��ޜNēkR�p�8`�3�Au}"h~�&�lڅ��S�'hH@I�ل�D��d])m#�����_�y�'�F$�%�ߟ4�|BW�0r�i�w���g+Q(S�zu�0.埈��ğ��	ݟ�Ryҏr� ��3O��@qc�U�Dݓ�� �g�4��8O%nZh�m��ɡ�M�i�T6� ���`)֊r3|lcUD@�h��J�g��:�x�(痟*Ջ���i����Bd���_kt��(U��H56O��$�O����O����OF�?�s�H]�p��2���-R�b��3�k������4Il�q�'�7m>�$Z�~�X�CTC$=���@a�<3��%��	����7LhEң��X���� M�x�D�q�V���9m�6,P�'��4$�4���4�'���'��R��=�	�ֽz4� S�'�R�Aݴbb|�ϓ�?�����)��C`��d`�t؄𣜰F������T𦥫޴]㉧��Ws<t��lڗB���GB �p����U�f�y���!����y�-\��b�T�Q����"Dur8����`�	���)�Siy�nc��#!޶-���v�@28���ܺ+�	�Mˈ� �>!��i\dQC�k�5?t�(��������M���i~��٣�����D��AF�(�����"!� "ԠW8B���C�Ҥ~�0�cyB�'���'���'��[>-�À1rb�憎d�5�Q�ӓ�MsE'��<���?yH~�:��w���dGر W)+�O��$�@!��p�lo���S�'nV��
��<YQ���lz�a2H�^��I�b�<�W�V���������4�f��ٔpD���Xw����o%?�����O����OJ�@�6fE��yB�'��,�vk`]��o��o|���a� �[��O�)�'�d7�OȦݩJ<i��I���n�0�bhs��x~�Oݵa�Ua�%�טO*�u�ɵW�B�?;�L�N�?]^�� �]�X22�'��'v��Sٟ$I�H��BL�D� �J�3.�;�Sџ��ݴx�Ty���?�@�i��O�.R	�rY	�+Ĩ+B1�"�5�$�Ԧ;�4�?asAA$d�'��(P��W�?iPT�ȼR/᩵Lژ-P�9eK$��'�i>������	ޟ��I�#���C@Cy�4�&B-6��'-h7��)�ʓ�?	K~���[6��R$�^n�Ph�v�l�`��S��ߴ:C��=Op"}2%�¼D�:T2q�-u˴�@�B>j@p��t�v~���6|���Il'�'�剂A.U�ȚO�b�("%�[��I�I韈�	۟��i>1�'(�6m�A���֍&�Yؔ,�#J..xY��_	d8n�d�Ʀ��?qdQ���ڴ&��'X��P�� ������NC�0��yʕɗ�/.���O\œ�K͖����k��ǏN�k~����-�MX�p��du�P�Iߟl�����П���(]�iq�9tO�.X�1��!�%����O�l�u,���X��4��$�T����8�uJ��G�r�':�I��M�����N0>r0��O�H2���%q�J�J����LU&߿R��(�� ��O���|���?Q�wN(�6�-^b��%��J�%9��?�,O��m�)^�0�'n�R>�x�HF&P�L��KV�(�r��)?1`W�tX�4Lj��9O�b?�i�@��FذI^'$�h2Aɚf�6j�/��~��|����O6��L>Q�\G�؋)N���T��DP:�?!���?����?�|�+O�m6M�.%��J�'$p�$�p�<v��Bs���x�	��MӏR��>�жi)��wo�#yK
e �X��l���j���dϻ9^��@���[!d^A��ԓ~*��N�15fᲷ��2=� ��uf��<+O��D�O^���O����O>�'P;�M���&��'Ů	�����M��hI&��D�OF��t�d
���5Z�� f�=A|�KB���ѸݴgÛ�7O��S�'߸%*���<�@�Y2�bb��U4ҵ����<a`��?*�$X�����4�����3J���C`�� b�c��P(_�����OR�$�O^�p^���� k�	��H1�Fњ_q	p�B��$��Y�T��T��!���*�Mְi��$�>���R�x��L�2��0/T�2!�Jp~�e�aN���cXƘOz��IF�/��e)�1��n�_.x;3d��?���'���'��S����j=�D��EJ�3+bBUNݟ�@ڴb�n,�')*6$�i�)�c��<>����b�C�8E��,n����4���p�8�e&�K����C�:��C�O��UzU.�1����J�f���e�	]y�O-"�'(�'�Dˁm��+��/zl��X���1u�:�M#p%��<���?yM~Γn�4�j�)<}�")1C�D��At[�h8ܴb2�&�;���9��0��n�2R5�-�`L�o�<_$�4�e��ܘ�y��˔V�Wy���@th�G�I ������ѹ?���'A��'��O/�	&�M˗���<A��5N^���C��Q��0����<6�ix�O*y�'�X7-����ٴA����J�f���(T�L��p�0!PM�'�h��' H�?��}J��}��i���+���Ъ˝`̎͓�?����?����?q����O�B�uGH��a䀍2
� �O����צ����(?qd�iJ�'T(���B�Y�8 C��'@vp4`%�$J֦����|:�m�#C$�'Tx����sk���M՚W!�H��ȏ7u�Y�	2z��'t�i>��	��I�<�$��� ݩ@�&��pHI\3��������'7m�"e��˓�?*�DY�3 '+�d�R'ׅraP��4���ٯO�m���M3�'�����ƈP$��Qb��(^�0�H@��\)�!l�i>ur��'
�H&�4X7�ӵ&�ƨHS�	�O��Zc��Ɵ�Iϟ��	��b>ɗ'I�7�&9¶T�s�Y+�l��#Ϭr���y2,�O������?��Z��i�t�? ��6)��@%R��E10'�S�JΦ��ɲ?��(F-?y��	�M�n�	)�d@��!�И����"��
�y_�0�	��H����|����x�O�������?k�@��5X̤�U��M{T$�����O�������̦�]�Y���Ig��AeBEb$�;z|���4r�F3O�S�'?@FPV���<Q'f��\=�2��M�$}�o��<��O�5��D׷����4�z����LP��;��4��a�1��\����OP���Oh�pɛ��ڹs�R�'G"��2W��i��:�����"'�>�G�is�7�Lr�	"!�>8��IV�H�1s͂5	���c�T%�F�
zj� N~���Ot�H�H�e;��	�LZ*Q��Mp9�����?Q��?���h�&���*���@ş6r��I��G��$�D�yj������ɒ�Ms��w��Y�7 �'�����;�^:�'��6���u��4
t��Ϛl~��;�V �S�X��h�X�x|�3CO�5�h,�&�|rS�������	ٟ�	ğzd��

��9�p,� !Ӥ@9�Lry��d�4��2e�O����O����$�9U|�Hd���i\ؙ���UJh��'�@7�ɦ�J<�|"զ�%�, [�H���Ъ�oU!%�ȑs�.C���d�Q���k����O��-$h��Hֻ7���tE&�<���?!���?���|"/O�mZT�e�	.?ft���-D8�!ËR0#/��	��M���<1��Mӕ�i��Hy�)��&gx�te�@�����嗺O� I �O�]g)����d%�i���!R�Ȥ�А����k�f���7O����O����OB�d�OH�?ii���<��HI�vi�p!��Vy2�'��7��%3l��O��lZg�5� �R��5&a΀BjD"Z���͓�� Ѧ����|B�M�xM¨�'rր�oD9s�M���Z(���K�$�N��ɞ��'��i>A�I��T��,;�I�N�9�:l� ����I�l�'<6M�*�˓�?q*������^6�:�AA\�������8�O��l��M�'���
���#�2k�		s樻B�A	w����ˇ�%��i>U��'c�)'��M_�fy����gٴH���$�I�����ҟb>Ֆ'��6�K�]�pPK�̝#���Y���.l!x\ޱ�$�OF�m�N�{n��r����Ɔ��w�`4)����M���Vy:e�A_~��a��u�H�)���(r�D�%���Ҡ�ݾ���<����?a��?I���?-��aJ
;>����jG���ȕʦɐ�DAGy��'��O�Ra����R���R�`ͩ�6Y��C!5x@dnڋ�Mk�'�)�Ӎ{��*��f��u֣T�-����pl��m�JE�>+���V�I~y�O�l�]�HU�E�G0��рO�>���'��'��	.�M�!�#���O�@CR�*U~�{G���̀�K.�	���J��p�4�y�S�\�p,դ(X�ݫ�%��0%|hb��=?�WA��y�� ^ḩw|�Yv'T6pfdu3&"Q�;��q`P��N� ��>uJU��
�&�ࠇ�6mV\�!V�/ք� ���8 |����(Af���� T�q������O����e��&>"�b��ܲ,q�Q��(UԺq�|�W#UU��)�M�v�IQ!b�eK- +$������xł+V�Ou��s���?xQ��
T+v�J�[�@;s��Y@��6��@�L �vi�Ðké?^�}�eR�l��V%>�^LZ"��&J�a�eN�bA���NH�	 �C�c�d��EԠ{�B]kD
L�i�HE�i��L;kuNO����O̒Ok��m�*(�'	O�K�����׷���'t˞'Y�	㟀���`��ʟlA��hPYZ�ǜ�F�x��+�9l��'���'mҖ|��'lb��?���ٍ6T� $hȮOK�Ja�(!2n��?A���?����?�QÀ��?%d�*8,�s�a�;,o Mӂ	ϭsћ�'K��'J�'J��'D8�����M��d��s3LP�4V�3`ȸi'Gt}�'���'8"�'�|U"[>���5E���h�M�pt�Ү��yߴ�?�L>q��?���$�%���f�M_H\��ǎ��Q')x��D�O����O��م��O��$�O.����L��u$�!�&Tp���v>�+��i�I��$�ɘ֢��!�~JDf�.VƘ@#�߾N�*��t�E�	��؟��m�����qy��O��i�q�B�[ ��hh��6��qӊ�D�ON��V�|�1O���L���'��$a�]o���ij�l���'���'@��O-2�'��Ӻl~f�[��
 ���=B#���ܴ�:%ȴ.�{�S�OCBmU00f�`�RO*�iO\%e�"7��O@�d�Or�P�l�d��?Q�'����ƃ�!5P���B@�%ڔ̀�}�ǁ�Ԙ'F��'"�"c&8(�Ɣ8Ga�H�U	X7M�OZݹ�(X}RQ����b�i�Q!�GƲػ���/�
|��>�%��/���?���?�,Ox,굊�4?JV S��ݿ~p�c��(t��D�'��˟�%����˟@����^{@I{��X$Ew�a��� Fh��%���	џT��ty��A��)��B\�	0�]�O8k���}n��'��'M�'��'���[��Oj�2��N�&�ꗮ��7!��z�V���	�����Sy�̀1P��'�?	2N��H�7��.��E	�J�9`N���'��'���'��ycF�'!�Bp���X	Ir )f�x��@�Ц)�	���'�$A���~*���?��'h��R���p�J5Y��$;��i���x��'w�d�KU�O��������d��n�#�kU�
�|6�<� �W97����'���'��dj�>�q�? \I�h�$H��	��L�W����$�i��'��Л���7����hց�%[l��4@�no�7m[�G��}lZݟ��۟l����D�<ф�F�lbY��7��i�����RÛƯ��s��O��?U���?"L\����"Lh�A�ִ��4�?y��?ivm��R���Ry��'����j�`)�fbK14�Nus��^�#��O4$K$)(��O|���O����Ɵ5������a̺�*�A�ߦ��Ʉ:%B�J�O���?�L>�1O̘�!<ܬp)s��*U���'U�Az�yB�'gR�'-�	qBBԛu���ZE��/�|:�KvD����<���䓟?���Z���R���o(�}���&�ڜзK�4���?��?�.O���aB�|���^��x�_�k��8r��͗'B�|b�'~r쒘��	Jm�TAR���F�� j4�US��	ޟD������'(!�S��~��Jm���$҂}ڜ=! �ߡ'�xqe�i:��|��';�؇'�>F�Y�u�©X���������צ�I����'U�*aB>��O����F<��B�8��Y�[ N��̙��x�]���I�p%?�i���M��}0t	K����i!����EӲ˓hPHㄼiC��'�?I�':��I�?BUj7cұ�`šԭZ���7ͧ<����?�����ܴ;ܨ��4(S*En�Ԁ:Nn�o���Pݴ�?���?��'n����dM�;�Rh���u�h�q �"_��7-�O���O�O�s�L���� !��� 5ڴ�Y�e�=���"�4�?����?qC�޷)牧���'P����H@��
Tpr����(���'I�I#@�<�(���I�p��c�~��sl�U�HA�n��9��ao�꟬���
Ty2�~R��K��2���c��L��!;��O͜�9s� ���v��?�)O�����D��щ�:f=z�0ŀש?�N̂ao�<9��?1�R�'g�cԤB��܃�D8eJ�B�&�?"0n�b�����'hBR�h�	/'؊���x�`0�*�Iʲ�Q`��[�<Un�ʟ$�	f��?����8)�����! 1��H}vAZ�eK7 d�H���>����?	����{Jna%>�q�Lѩo�����N�)�hU1!�1�M;������$Q�{C
��/��f��@���)D�{��h��Mc��?A(O0IR�`YN�ɟ �s�as��Z�~���3!�"*p��k{Ӻ��?Y�"������'��1��ys��]��5���ׂ{W��d�<���Z�&U>����?�[�O�L3С�&	���N�5�n4���i剁&aT��&�ħ���ݺ���n�H��K�)x֍x�!c�~�I���O�D�O����S����m��\3E��?Q�@���͸M�,6-Y2��l������"SC܂x���J�2=>\�Ƌ]��M����?Q�����b�x�OO"�O�Ղ5bO�<6�93��> yq�i��W���w%����9O��D�O��$��XA�fn 
��S�%"�oZ�l�'����|�����Ӻ[q圼	 �*��
�m���sr��n}��J(s{�U���	��IWy�ÄB�tM�B��^�@�a�7c
�(�"7�$�OD��O*��?�М!��Ν�d�����-=�v���/�+�?�)O���O˓�?A��C���d�(j���H�f�1`Z\]	�lԻ�M����?9���'���D0�@ܴrjn ����$�0�r#�4b��i'�x�Iryb�'��y�Y>���$�,��ci�H"X,N�.�>�a޴��'fb�'*�aA�����[~�`�eF�/~�P5��@[p�Xo�ݟt�Ijy�K �?�����$�kl��s��z7@�R
��ucT��'���!R�n-�	q�SGj`d,n�X@�@8ѣ�ZR}��'4��x��'��'PB�Oj�i�=�!�/~b��㯊7�Y��@fӆ���O��i هT�1O���A#j�}	j^�9�R�pָi�j�aTBu���D�O���⟚�&���00�S�L�!>����P��гܴZ��|K��?�*O����I?U^~� 5�� `��pqm�Q!l��4�?���?y������?9�O< @���0.p�C�D
���(�#\~̓0�����O��	:_:<��n	�\�.H�Wm�h7m�O�9���<YE[?��?����1O`q�E��^�! �/X�L��	�lr���>?��?I����dצ0i�ŒBF��T��l	�O\?K�9���l���� ��C�xy�n
�/*֌�Ɓ��M]j�Xen�aL� �b�'7�	����ҟؔ'>�DF�k>�H�X�B0��2��+yY@��>����?�H>�)O4� 0E�O�S���&*Yh�Y���=T�e�@[M}R�'B�'��	;Q-���O|r�	ڪv:5�.�%�~��Q��*11���'��'c�I�2�4���D�I	�5��A!A��@|kq&>oЛ��'~�Q� ���=�ħ�?���a��!X�@Q�o�a]&DtDp�hyB�?�Ҙ��ٟ��y%e�+/�2䙵K�T����i�剚7��l�ܴ0���ן��Ӭ��䀚~)��ׯΌ1�H��jW���Ɵ��QfO�Ot|&>�%?7�$i1"y2��7�����	�	���CʲO�7M�O��D�O�i�b}bU����o�\���+���;�����_��M�$J�<�+O.��"����e���R��m�Oǵ6�|�#F�0�M����?���wp��R�l�'���O� ���B��B)H��@G�~��S�iXBX��K��}���?����?�BA�>@����^'|�T�B�
F9��'M6����>�)OX�d�<���kR��)��Z2oڷO�
�!%UO}R�����OJ�d�O0���<9�%D�{�|᥌]z���'-ɰ5x�]�Ԕ'i�Q������8k^����j\bQ�"�	�AC�|��e���I՟(������Ly�L�.)wn�S2��8e�O�X�1c'�)��7�<1����$�O���O��72O�)�B,���Bc��
!j��4!����ПP������'��ɸD�~B��`(٘v��(:��+B�D��9`Ӻi�2T�$�I۟��I�u\�c���*W4�@v��f��{�I�����'��\�FD������O���|!����;Y�\��e���L��I�@}��'�r�'�Ұ��'��'��^�>�^�`r��L��2c��h�i|�I�a�2��4�?����?	��!c�i�1��\�v<EPl�LyƕP�~Ӕ���Oޝr�?OZ���y"�	�g	�R 
3$�J�:�/ˤ]�vBM+Q�6��O��D�O.��G@}rT��K�c�7z���wH�#nP9����M��Z�<�K>����'���x!.�RPv����Hc�@2'd�N�d�O:�dW�4���'P���h�2Y�$�k�1�YY§�5E�H}l�ݟ�'1Ș˜��	�O�D�?�h����z�<�1b�3CN�4	Fe����6���'j�	ß �'kZc���O˻%����T�'��,b�O���$=O��$�O&�D�O��$�<��l�m �u���.��tSp)ˤn�$�1R�X�'�S�\������=��Qp�F<|,�̑G��+@��P!��q���IܟP�	ڟL��yb!�
2���{���1>Ȱ%0碔5�t�ٴ���Ob��?����?I���<�w@?
zZ��(8ထ���׬w!���'��'<�^��Kq,&����O�(�Ө	7ZJBT�V �5)жj[<�6��Od��?Q���?q�.Z�<�J�Dʃ��[�T)�,ؖQ���s�~�"��O�˓b���Q]?)�	�t�6k0��k�j�91������*B�zD�O���OT���/f�D�OD������kCt�8AFè'��cjQ��M�+O�<���m̟���ϟ��ӣ����4M�.��80��͓1�j��q�iT"�'T��'<���<���$���v@p���a�x�9-O��M�HC.%���'kB�'3�$��>+O��k�&A�:��hʅ�N��A-oܛvn� �yR�|����O�DRdNW����c)zK��-��޴�?����?ѥ��&��Idy��'^�ğb�����/��k��Ŏ#ǱO����$�O���O�i�ׯ�w���w�8C�l��%�զ��I3H�� �O���?)O���Ƥ���8 >� #�MA�P��Z����>?���?i��?-O�����ū�B�ãǖ�W��B҆,EY���'��Iן�'���'\2�ϊY�Ń��5��T3%�#�4��'4�	֟d����Ԕ'��Y8� s>�' SD%� ��/'� ����p�ʓ�?�-O���O`���s��A&1���s�ӓ<�)���P�R�m�㟘�Iߟ(�	Jy�ňz���'�?y4"��8E�7h]]�E
�bL����'��	��d��۟���f���f?�҆2Ml$ b�t�:�Ĩ��M��Ɵȕ'��5`C`�~���?��'~�t��7�L�G�t|�r�D�z0kQ\�8��֟ ���|3,��ĥ?��a�b*�8AT�����p��mxӎ�FV�hX��i���'+��OӶ�Ӻc�dF*P��E�!���`�������Hp*d�D'���}�w×5�H�����)��7����c� �M����?I����7W�L�' ��i��)%��%o����7�p�t��>O�O��?)��*2(�R��Ũ3�K6%��M2���4�?Y��?х��Gz��hy��'��I�(�Z�S���&��Q*� ��IQ��'���*u]�)����?��OK����ń�|����h��p��ڴ�?1��J(���syr�'C��֘���� U�U�O�.�E��Γ�?���?����?.O~����?5�44�C�]*5���i��W@���'��ڟ��'���'kҠ��07VUcb��+�P�Ӓ��
T'#�	ǟD�Iɟ��O)���0����2�q(�*�Xi�q�xB�'�'7R�'ih���'#t������3� n��ّ��>q��?i����dAt6$>u���3O�1�����l��D��M����䓾?���C*D+���I,[ԕsO�Ie0�
aI.M&�7-�O����<AhA�Y�Og2�OK�E9���{||8��J�
0~�@m%�D�Ob�D�',Mr��/���?ͣRO�9_����썁hKP���mb��˓f @[��i�&��?i��9(�Ɇ;:���H�*$@���Or�6m�O��	�6��5��$�	;���1gR�MCP�KA�U6��1�xAnZ��	՟�����'������@��<Ǩ[�ʐ�r������O�O<�?�	  �ʕ!��:򎝂�	��8p�4�?i��?�ӥQ{��O*�伟(�%ˉN�P��W��4Ug�@�6�c�`�O�ݚM�G��ğ��Iʟ�rBC������ɞTn`p�����M���3���s��x��'�|Zc�2E���8��u�B�>	h��O�8���ORʓ�?���?A)Obd��$4C�k���{;�p� �D�IbL�>9��䓮?1��b�� ��C�Ɋ&4�¸+#�Y	T��4k�<q+O(���O���<�c��:��i�m�މX��)_�pz�h����|��O���x�I(i�@�	�e�8{A$Z�Xh��7�Щ����O��D�O��<�w�I�#��O�^ ��!oM�LU-.,�rb,f����+���O����-$����#}�@�PȌ�C@M<f,�T�0g���M;���?�/O�t�2�h�埔��P�NL�RL"`�&�"'�X?�8H<���?A���<iL>	�O�mPu���j��0�%B�L2���4�?Y�������?�(O��)�<���.�Jw��_ш[��R:8�o�ş4�	=r���h��8�)�CДs�T��hE� �T	"�72J�z�n���(��ȟ��S��$�|��89�n��T�#���d���sԛ��43U�O��i*���O�Ȃť:��m��`��
�hqC��������I9N`l@�'��� �v�d�#�JÜP�8�����c�2)����K����&>M�I<�ɬ|�0E��ɒe��{�� 7�P�4�?�����?�o�����'�@����j��t��N�J�P�EJֳ��DԊ61O@���OJ���<YCD)�������N�q�Jр6ײ���x��'�'��	�4�I�G�br�	:������"#H�I��b<�I��(�Iry��'z��Q��d@��	��NB���m٬FY��B�i��ş�&�p�'���+u�I��Ms��
4]u4q:3�Z8+�A�l�~}�'�BY�X��Id�~�MY=y�:�	�	#B�1��ǃ�M������׻o���5�x�jE�$c�,O�$&X����į�M�������O(��R�?������j���2%���HF1[�G̥�I<i.O�sӇK�K1O�STݪj��#x�V��cɴ6��O��D	�<;J���O������?��:�n%�P�Y����QAW�f��Um��4�ɾ4,�"<!��/�'�mb��?]���P���	�M�An7�?Y��?y����,OP�'Q����.m�ժ�8q��ictl���?�Sݟ؂Ǎ)
F<T�õ#�j�gù�M����?��h�h�.O�ܟ�3z�8�u�^���I�&g̙`~dm�T�$\To��%?�9�@SnpH��i[.��w�
���<Q�l�#Rpe:
�'�Zx�ա�$+ �}@c�[����:דU�T��n (m��1ɗ��TXni���TXf�!ѩMO(0 �c��p<$������Q�  tV�h��Č�`0�`R���t8Db�P�:��d�V�]'C-����`F)�re�iJx��d�
�f^�"a�U�[` �I�0sLD˕�J8(,��l�q������&n��Y�	����c����,���|z��U�h����l�:Y��a�a@Ly��=����ㄈH��?������	�Y�i$���>I!�͉>����@F��<B��)��i�&#�>dԉ�N �9Rޕ���D�'���؅���!J�ѩ=����yr�'� ��b	��O��XK�52�z���'�6Mȥ����tEQ-a3j���$�0��D�<)�I��"���֟�O�Y�&�'�q�n/2c�|��x�Z�'�2g<%�d�FK�A������O�@��d&1J0�!�(Є[�8�ر��I4>kd� 柨s�X�����_�O׈aP$��;W� "g�����T�J��YD��Oz��<�'�?��`H�+� �-�cwɂ�}���ȓh��R�.�%4B�( �ױ%w ���I��HO��H'$�<i,���+*J��	{dDIk}�'>�B_�`Q��'��'9�w�"ȣdL��0�4�a�B�m0�1�莴l�x�C��O�hx�e���1��'�Bm"���0��H�)vΊH6�خd(}��E�O��tJE�����LR�!�&�E0Y �'��|g�S�����-��O�ў�R�/YD9����-L����8D��L��?�\��)��{P��g�;?y��)�-O� ��.е��(Jq*3L9�P�JQe��(����O��O4���պc���?A�O%Jik����Db�"z�L���Dې�x2'ʜ�]i���g���*�f�!A9�]Ru"�3j:����15��#�!�=bFa{���;���M�m�:�c��U^2�����?y��$=��%NNz=*@+�	L���X(_��@B�I�a�JMK�lM0���Ѧ�]$0�c�h*�O@�	>z�TZ��	6xݢqZF� LY�E���a��M�	㟠)@�������|ڴaT 5�ܹ��G^V��u��4r������u��c�&�)�H���0l�#Un���+#M�)�� ��#��=�4��4\�DQ��+O��
��'�bR����I<H�@�23��M�+,��b�4�Z@��n�.b����)�_xB�I�M�`�W(+6�$C&G��)L$)����<y����_�*�y3#�7Gg���*�I�&B��8���A��-�rHS��f�C�I-��x
C��%K�f:��L���C�
`7~�;��GL:��A�)�!�� *�CQ��?_�H��c��l�$"O�(iVi\hX��K�$�2��"O&�)vk�"��l���&"���(s"O�����[��a��d�Ҥ�ʕ"O>tKFh_X�𴣵�J&4-ۃ"O\]�P#Y�4�N�H@�� �rh�"O� i�dϭ.�,�(�X0��(��"O�pX�N�(��Ȳ�Ş�P� A�"O�`���Lޘ`��]'e�4�H"O�@�Bb�j��XtI��8�|5Y�"O:]C��m�����e�(|R"O�P��50�s^�� $@1"O���f�R�5�>��C悲X	r�j"OF�c�k�Z��P���+h�i2"O"�ⵆ1h�
r3��L��KE"O`t�ԌJ93�ԓ�팚#LE�"OT�!�i�-0��)�W
�+_��"O8�0�l �J1����S�"O0[#�X%4�^�!����1E�hs"Ot-�K�:Y�4�kc�U�fX�"O��w��14���ztF+_(��G"OT�`���U������U�9@�%��"O.e�0�2Ρ��C��\��Ĉ�"O��p�#F1��Al�I�HX�e"O�0�ۈ�Z\9R���*B��ʄ"O�`P4#S�hV­��OC�M��].�y�
�8x`��/Mv˶jքX7�yr�J�a~B���Xm5�<��l�-�y҆\�(�B8%HY��Xǁ\�yrH\�E`|y��2�����J�y"��Y=X�g+���Q!f����yb�Jj:t���U���]��y�	�lm�-c&�ڧI��T �-��y�˓2Yf���E���q��y�)Y�td�@�Q��=-��{��V<�y���9D��Q�%���\���	Q��y��ޤz�u` 䊀r�DKp���y2���~��T�%j˞��T#��y��I�l��Պ�Z��1o=�yB(^v�z<�sG
�t.}�U`9�y"�۸F��IE���(�r�el��y��A�~��s�J�/(��tB5���y戅�<�sB�,�<�T���y"���>����f�r�����p<����&�qO���t���"���+�%}g4H�B"O�-)$˝;�&ip2kW+~ZP ��^����ٌ-�b��|�䫝vgF�j����t��<�@�Ju�<1�kY�-ತ�l F$E�q�dY/FY@�J"� N8��#fȿR�����ń�HR�7�O���q��`�9�LbH�3PH�KT�є��'(ڄ�0?A$�¢? ����nOX޹	���x�'cȠ�� ;�:����7����O�Q[��1q3rڦ�L�
�f�'n-4���d�.Z؁�0J�	y��h@W
�O9⦍8O#t���&�&4%���g}����o}5C�i��o�*���I4� ���@��X Q�+>?�y
Sʛ�SZ1 �%Reʰ�'JN8j�P?7��/%�J��
t��F��r㯁�(�b4���=�O2�j-͛nX��oъs�fx�Ul�]�>��Jڼj{�:�g��?ّ�C{.�����R^���ME�HMiԮ��OQ�L[��	��^���E6XHLkЦ��S"ku!��%�f)�Ӎ#)50$�
�'B��ЗM;d�� �\0e��X !��)=Y��A��Q�Nr�Q�e�%P����#&́�&3��Dg���
'ʓk�`4c��S ź�;2�Z�J��D��
'l���V��Y�	X"@��c�����&^$
*�%b�(�V"'*�m+�&���|�Z�� o-�c�b>�K!�T_;��ç@K���3S���77�����CŴ�85FPs�zw+�H��:P��� @��7��p��h�J�v1��p��O֠+w%Fq}��	P��̱�M�k�����M,���#��yHV�V�M��y %�>��8��捅`�x嚌��*E5���}�0���O�H,�Fj�1?��m�0f�r 0�a �\H�2��זw���OX�p&�ƴ�ywɕ��.i2���d��fR�b�b�<i�/�'S2Q?a� �=jLl���n7��&Y�@ܡJ>���	P�3[��kC�˭F�r��w����艀G�m�V$ X��N��(�>�~r�I�%����C�Dԫ�J�2W�b%t�U'�N�{�@U�~-�-q� F �Z�s�╾Dթ��D�7=��HA��:z�du�#�";��DNV���'�]s�+	�p\,��SDF�{bz ��'�����X 75��Z�i��?�X��#`/М%0�C��O�Ⱥӎ�}?a�MO�Tu$�z���0�Q���Z?�'�g�j�	ρ:i��c�E_��?y���P8����|�M��m��V�BL�3�MP�'��$ATM+���)��ؐ<��8��܆r�����!�;�����Nm)U�	��	�'^^F�݉m%�@C�w�*�K��O%un���I��4������@&�t�>E�T�F�))�d�T� ���s�j� 'Q��Pd�X$
T*�p�� �I�e�D`�'
L��&嗧 �>��uH��z�����'�,%�t�7���dT���q@��:��ӣȄ�)~ ّq�\!T\ա��y�*�+��=YإQ�e�'ԨOX�G�?��R(����Y+z���!ky�ɓ4b0�K�<28�@��VW�6�^>f>`��>��`�ת)�2�1��	-n�<���	�aiV#*��a�)��I�1|8��4@��0�I��}T�ÏÚ
��X�C�g~B��k����(UX]i�"ٿ[D��H�~K���7�BV��]�E!
O�"e�[�n�Xs)�l�頔��p<�DXm�,�0v�vl���Y���Pa	)�q A✈eBB�#E��v���煐�J�$�X�	��	#C����$��C��=���A8#��5 v�ɖ�1Od4C��Фp ��8G��H��1Ο�X�(�.���D	�]L�Z� "@�`C�ɸN�| ��
�	F-�`�d�\�7���r�"m �c�J�FΕz�!��l �W
)�'>���gHK�X>���Ta 	̄��"Od��ň۰q�}Aq�\�90M��E�:L8M�%pN�+��$����O�.b�(qe���[�$�s��BZ�h�{��5LOR��c-�tx�x�F�;Vܐ��D�<aj�v��DΈ��h�-���]������T� i�����V�(��)�8~�qO���m�ezJUH�U���O�Z�K�=;��rޠ�Dt�U�*�!�1x��a/ܚ�Ĩ�v�]�V��I�q�r�1�>���O[�h�¢��$�L�k̘֭G�P�0�'��j\!B��aQsN��*�MH�yrF��n��l

�ؾ ��-�6Eg8]a2˞�z����RP�EQ�v|�Y�&�x刀Sv[�����O��cf�T���s"�h�V��㉻i�B$
��ĉ�r�����E��|t��bFO8�!��5����U�՘K�=@ '�\��'�,d; @/�)�ӠF� �n�>$~8h�5+έu�fC�C2�` @Q�M������Lj^C�I/C2�5J5��|�ـ��;�FC��%
�����CH�C��Ⱥ7�	�h3(C��4K����CE���թB6k�B�	2O������Z�<�h��3u��B�	$;�����8��1
���&i��C�	<n�.�YRlܳ-����u�ڳ^��C�ɬI/�Q�	7���{2`*+APB�Il���D���(�,�x��
G B�	0c�%ʲػ>�h�0��-:C�IzpM�%*k]T���GP3>� C�ɛX�t��s�Ѻb�.�ハ�VC�	4`���L r�ԙ������<C�	�z�T�]�i)�E��c��B�	?|�F�:b��+�Ϟ�c�C䉝nCr�㬐�xx�t�W�6͚B�I�c5"X��B�v%
��ՂR�|�$�F8tz��' ��	j�����#v<	�hIh�q�aƁ�y�O�
0�ꔡd,�#i�R�١�ԓ�y��|�L��둈.D���虨��'9S���?-�?)Sbэ[;t3"�3���P�4D�L`Ȓ����Iv���K�'ǟ�y2rbx��]��~Ҡ�)c��&LI�:��`�����~��5eB���� �HC�	�LbT��DhG�2u���'�����F�)L�Q��k��_�~�ĮH���e(�*  Lߪ=�Hi��DꁯZ��	2y�撟����'D 48q���	�t�$��r6�ʊ�dB�(L0D�OQ�2+�R��:�6ͰC	�'Y��j3��)!&8��k�?�0YҝϘ��i����)"s��>|����ځk��H�� �ا�:t��7�ۃo��� �?W��N+%w\��f��=!�Q��t�1g;qa���'Ϣ���B�=�ȩ�$�;q�8��xX����O����U������J�9����9[��B��O��+D�f��$�r�S s9ᚰm^�fHD@(�M0)?���>�(�Tr�I
�T����D�f�δEy�M,�D�~
SN�^��0#�l�R`Zaht��4�Dm��I1&�vM`��D����F�R�bXh1I��
��P���	l�8���T>y(�I����p����?UR&��;P���ar����0z�C䉆s\�����ݒ6%��C��L���	.熔i���Hl��6N�;*�D�9O1�j@w�تf��i �P,G"<���'�T<�p[�<��-YB>9�0��;5@�%��kΜ?т���8��h���E��O*0�O%u�Xpc����5�yI�剕Pa:Cs�S�g������ɂ��L��U:v��T�)��A��(�����ئ*Ɏ|���t����M����ا�	��d0�`@@A����e���
7��y��
<�\�ȕ"Of��D�S����[Ѧ�@�� p��'L(�Ȁ+ɾm:9Ad�
 3�v����yJ?��Վg���P��?3��)ά>%N�8ӓx�|ÔgW]?���,�^�(��<~�*�΍�2P<��6U��ϓV�̨�g�'�D�wi-f@�*gA�?�4@Ӎr�l�(�����ޙZ����S�<Ҡ%BV$�u����(]�:Mp#>٧B�@��� K��ȅj@��&�*��8S�L�J0�ˉX�b���O�m�Ն&u�����
D8`��aH1����4> �=�l���$� h0ܹY�f˜ �]Kf�ߔ!��Ü�g��IR߷`n�mY�*�"�����禥"��!QO�� W�ʊ/�NUA��S�%jL���ˈ+�^u$�OҼ�&#Q�3�X����+�(l��"O�T�� ܗ(�ĕ���Fz�!��	;l�x�a ���0g�-a`���@����ȓCHh���J�pLБE�	�����9
�閯�:jL 	 ��:�4��z�6��� ��{Ծ�x����E`��Ql�Tp��ǫ�(�x��C�1��|�ȓ��I�� �FS�8�<!����"E�	+��O��B�ܝ�yr�T59}n@��쌥z�D4crAB��y�	��0�`c��fD��*���y���1���l��cS�Q���	�y�痤2S��q6i~8����I��y"K86�)��J܅�d���@�y�DIS^������q�@�K�#��y���!��(��C[/oՒšAf ��y�� *wx9�t�H1d�*�q��6�y��_�n��&E�D=�����,�y"D �*0��P���<Ř=� �Ī�yB�K�~D
uL�41N�P��y"�Xy���� T8_�r��)�y��Δf�L0�k�8Vb4p*w,��y�.�(>^ֹ��Ԉ�5"aU��y�ϱ=���-�0E�rͱ0c���y���np���O���mI��&�y�BA!~�|��#��u��Y�yBm=WJ�U'�(���a=�yRcH�b��Q���N�6%$��y� N�I��ٰS,A�^�v�H���y"ϙ��ޅѲfW�V�RA�7ؖ�y��Bs���	[�B���l?�y�,�0�
$Ђʄ�ZT�����y��1?Vl��އ��кCX�yR��a��Y+��	�v���ԇ�yb$� pޚ�J�	��n�S�L���y
� И��(� -�=Kw��:\�X�"O��Ó��7���Rb��O�>hs2"O>-�"ͿM�D��� �`�;�"O�ɠOѻ3~9!c��-L��m�0"O�LKA�� x�x�!o��agd�H"O29�ׅ^�0R�"A�՚d`|��"O�E�'eܢY�:�Ag-��qs򤰤"O.�1nZ�9Ij�:���H�"O4@u��$Ed�	*�e�x�v,�d"Op�a��qB�2�ᑹ��5�a"O4�L�?��a� �9T��B"O�UX�F��v�V��Woۃ{V ���"O����W�N�{3�]
E#F9��"O:�zTK�B1Z�c�ylr�"O\� #ɋ�'pm�DE��1���S�"O�xX�ˌ�}0�]C��Նv�(�u"O�����?��H@�B[��-�f"O�T1ԏ�	uM������4�a�"Of�S�]�-���*%�0*��Q�"O�uy�l��E��E/^�4u"��"O�}3u�_"Vd��#$\C]���"O�M8b�Zo�q)ǎ�62=T��"OܙB�+8����ц{"�\*�"O\��)�&.�]�1hڏe"U�v"O�Iv-O�U��=��D��s��2�"O�Iz���
�H<pt�̓\ Љr�"O��p�G���A�鐴�"OP�A�A��m_
�y&�V��X!Q"O�4��F&�щ���>p���@4"OFи���rĒ%o�#b�>�B"OL�7�g����W��� [3"Ox��T��h�Cv�ϝX����"O�\���!�e�GD`�)�"O�P�̇,B�ʳǓ�v��Y��"O�4!%��e��6'ާ%�����"OX�34EWT�A�HȚ+�؁�G"O��QW�C:Vp��F���"�!6"O��0Ѫ_�H��w�9k��2w"OrL�P�	�бs'���\0^ثU"OJ��Q�\�{�<�҂Kߡ)�8��e"O48��V�7X )��i�@Sf�A��|�)�ӎBL�s�3@�@"G�Vb���ȓ�z��a��yĮ�>$�ȓ]�03a��U��ᓧi�d���ab>�R�e�V�a`�JЁ���� R�y�ǚrxXY��G�~�q��w|��7X:�*@&�D���]��
!|�`lA=%Cf5@Fmɍ���-fH}`g��" 8�C���w>N��b6�1�����-�5@�&N)���ȓp��]�a�Ɋ/j"	0��КE�ԆȓKn�����Ϧ͓�/�=�ȓsG|��Q
5o���YV�Je�t ��X�x�0vƋR��S7�8&�\���@)<���$�� ��5�J��.܅ȓG�PȚx6�S��v9*E��6�&��Ř�#�$A�Q�.$�d`��&�<!�V�̨��x(��=�)��;������#ai��hQ
�R�섇ȓY "H�'抓�&�v釾Y�r�ȓx��;�/���]��ʓ.n�1��-���@篖�s~J�)OӧQ�ɇȓjE5�3n�p�!��M�����(YM�D&�г��Qn���S�? ���KJ�@�r��g͒O8\KF"Ob����D%: �Q��,��t�8�S�"O ���U��6�q�,Rp���1"O�Xˆ���`�q�+?RZXX��"O"�i�GH�HHS2�5(A�!"O�� 4"�;(n2��_
4�j=pr"O��鱄E��3G�_�X�,�zA"O~�+��^�O�n:�G˛W�4�`�"O�y��Gϱ6\<�5LGH����"OJ�C���
�41�H�6<��Q�"O��yC��zO�x��
9T��"Ox��M��I7�}ˑ'����r��'K�<[��T����O�� �b�(*D��ke��+�m�̉J��jD*D���&��"���(?K��!S��)D��2T�\�=Z`�c^Q���4D�h*E�1<I��E��S��k�N5�$7�S����څ�	OEz4���ݿ�N��ȓ;�6�R�X�驁6)� U�ȓADN1h���;,���A#$�/vq��ȓV��u��(ֈ{�H}���P��!�� 6\�s�A�b򔵰��rC�ɠ+���V�MGl���ї`��C�I�6�}��%��Ik��N� ��C�IBdZ8�ë�%t� ���E��C䉔+B�#�\9!D�*Ʀ�\>�B�I�VXT(����\{lHg�C�_g�B�	6�J<#Q�W�y�J	2@����B�I�Bu��8tF�[\<����&8ŘB�I�f���b@�"9���
ςw�lB�I�z+ؤ��/�!���uN�qb�B��4Z-P<+�Aˊ	��/Me�B�	$�4YI�1 
��G��X<�C�"g����ʋ�w��������;ͲC��g�lH�S�s��\�&��l��C�I�X]�x�Ek��"��HL%6^tB�I�'	2q�c�w��D B@�\�jB��$����&ś'4��F�8�FB�'_"Z1����0-9*k�L[�<\�B�	o��p%&�\�x����<�pB䉫&�򈚦��-}p��7�� ZU:B�I�K�j�U�H$=v�	G��P�fB�	<��!�	B��.��f֥\��C�	�;�BTs�&���j4!bHڇi��C��2\�PD�dB2���چ�W~�4B�I?^�,�P�ޅSG�H3�٫WMTC�#^
I�C&�'st��4
��S80C�� v� PY@�ݠK(���C��,WP=���N�_�eS4��U��B�Ɏ⬉7���zC2���Y�",�B�	�3	�p+f+�(j��(#�[�|�B�	OTp
@Z�ax���j�AF!�dB=~0P��.G:&g��J	_�n6!�D�Y���Β򍒶JR��b�'��$��D!B� ��2���A4�'a�M�d�ߍ1c �Y�G��9!�T��'k��1`L=e>:����՞���P�
���h^8q�:X�ը�`���(,�\��	�
v��u,�>��ȓ6�b�Ӏ�\�z_0 w,H&�LD�ȓ$	��w%I-1�ɳ
�s2l��p�E��l�6��I��iY�6��<�ȓ���z���5n�Y���P�[�"�ȓ040��G�?Įi ! �&8 씇�S�? �cp�Թ{\t�8#B�C�H���"O��K�A
=)�ԐK�I�e�M�0"Of	FO1�4P��FL=c~�h�"O��(S`��,���S� �Q"OTqJF(�&`LR,���ʻ@;�x�"Oh�� �C�<��eMK�?􉐦"O����`�}4���N��a�����'ޱO�xRE�@a�92'�
��]�"O��ZRDY��*�3�4L��"O�a�R��5`�(��P� ��Ad"O"�!�$�(����p��[�"Oj�!&���r�xع�]*@�
lA"O^@��ˈh(���\����"OZy��h�b���3�M�Ht�"O`Z�̈)FKr���ިJ�Z�"O�Đ` �	?���ʕ�_�ZB���V"O�@0�M��LI�p,�W!�%��"O8��&���0�Y�f��~�Q�"O������W����$˃�+ȉ�"O�U����>��)�	ӈq�H��"O��IfNG)��1����|�N�*�"OJ-�a�J�uax��a��Xˊ���"O�9	�*�z�t�M���"Or��s�M��D7�����!"Oܭ��A
j\�m'�ϽAϾ!��"O24�F��*M���85��h��"Ob=!ī�6�	�	��N��[�"O<t��kZ:����D���1d"O��k���)���SǕ>�d�ȓgǒ�@�Ϗ"i�@a%g(^~���%(1�����l
��I�>��I��LZl�CsO�.7n���
4�"e��}ה�Y�-�l�b�A��Z�R����ȓ3��tYKؖ4�9@�C�����=�$���F�64�Ā�<�8��ȓr�22��Q�u�(ib&�-Bq
%��?��ȓ��[jh�b��wY�ȓ�d�!	6��k�͊(C\���VU`%�bA�S�����&
�Nq��y��)hG�ՑC m��]!c�",��w�z�֏K?SY��J5"�^�V��ȓ?}�E(3F�*��������B�]��b(& r��<Q�S�ث,:�����ׂ;�j�PA��8N|��iǍ�F�<�%f�9���w�ϝf���@'c�y�<	�9Z:��6��O
�5� �x�<�"��d��P�a�7T��@A��K]�<i�IT#İ�2�L�8]p���W�<iuf���<�ңjW�Z��� ��~�<a!����ѥ�#P8D�"2�S@�<Q��=l �e��/�(=���z�<�CB&1{Q�#%�5ߞ��`��_�<�V�A0�D�(c��c����1 FX�<�6�Y2-�{�d�7d�	Vʏ~�<1>��K�	�1eA*�q �y�<���O(��@�a�(W��|a�$u�<ч��+LQv$����xyyU�m�<�4'��0Ip,��x7q J�g�<94dĚD4���Q��>L)
0�V%�h�<�bN��W_��h6�O?6�PX�jIN�<�2���Q�v�c���#w֐���FH�<)��#�6p����+�\����Y�<���1. `y�C�RNh�o�A*!��ҬLVhy��c+d`�-*���G!�� ��@�$�8��1��)Ԥ�8�"O|�i�k̆J���C#V�'�bH��"OB����4���`� 	�S��!"O.l
�G�o���("J]!%� �"O��KD�q�!2��[�]ĐHw"O�L�U �2�=��a�I��Ԙv"O^c`l�$t'Z{��H��X�S"OF�b�h߶B$`���΍4Q���A"O�����I�5z0��RN�1oO���"O��r��O8w��ȃ��/G�tj�"Or|��C� D���2L�pԜ�b�"O���s�ԲS��|BQA��yK�"Oژ�f��n���@�?U;z��"O��@�E��Wb2��v%ÂA*�X��"O�#�iT�Sn��#E�\=�p��"O�UX��/0�0��QDTa\Z�ؕ"O0�y4���,�h�mMt�b�W"Oȼ�"K�2��Th�6A6T��"OP����/G3����,��H��"O|����r�赪�(c��	�"O� `� B5|�L�Y�&Έb��K�"O���DǨ����^���)w"OH,���74FJ�vj��X5PP�U"O8����a�z�c��-)�k�"ORĳv��
o��Ѡ!��wF��"OJ9����
��3
��o����3"ODd���):�pD�6I��`�t��"OrA��T0	*�����2$�H9e"O0�!#C�eDx9�aKƟ]�e�e"O�Aࣄ q�|�&j�	>Ve��"O� �l�|���8���{���c"O����#)��C�S��m"P"OJ���4�0kp���tE"O¹Ir�<l8$�	�̈�k�I�g"O88�V����i��E2D<��"O���w��K>%�7�i�UJ�"OMPԆ*�t����2zzLa�"O�zGr�^)�GA�c� "O�qj'��`�&i[R�[ib|e{S"O��򕦟Q��Ѣ�_$k�j��"ON�*S��|5l��RÚ#(��r"OF]�̍�ƢuS�T�c����"OJ���"+p�2'HU�{�0"O�!�̞�0	"T٠��j �!9�"O�eA���.�����'
�u�. �'"O6�hf�)t�
�u�F"{)ND��'���#a��C7���$��	��|�'��\�D��n���
I��|{���'��(��&Bur ȵ)ʇ~M搀�'Rĉ����?h4���v��3�'Q���s����E�0Aq�f1�
�'b8!Pb� �M;�X�`+�7}G��'7긒�GF���UiM#-ehq	�'k�����62M���Ef�+G*�0
�'���u熺T�2��`�K�(�@A��'=�!��Iˋs��e�2�'j	�'�m�U�e� �9%����'.(`�4�Ɔ ���I����,v)��';�!��פ;��X����6,|��'� �����,g`85#M�����'��򫘅+��i�c�:�dj�'�� Bfa܋L�z8�v��,�u"�'�D8HuK�VPZ�rV�δwݨh0�'��y��7BFDP���<vޮ,
��� >� $�"���'HB#�V�2�"OKg�$V=�� �-C�1�2��4"O�0AC�[<�)�%b_�a�����"ON��U���5�P��qQ*�""O���AJN*,�@a�r���e����"Od)b��uN�� �PZ��"Obm��.��vD|��.E�	@6IPP"O���#�H�^-�<r��_$*=h"O�(�F��_E�a�"�6I���"O�5��J֬(S-{Q�:* ��"O��0��]5:[(��M$G=�1�1"OĤ2��:Z���@|���e"O4X�Câ6���K��ȳ7~��Ӑ"O��XCݺ��0���N�Vc�q�b"O܁ �`�{�e���[�2b�1��"O���Cƽ	�f�"��2t^̻r"O�X��[$��a�F����6"O�iKń��Q���s�$��]��I�s"O"��+ >��3�$V�$�w"OVyم�I�M���
� ]����� "O\��F�: ^H�1Q�Z�fh �"O"��#q���t�[����×"Ofx���H�j�y0 %7Re����"O�i�nަ0o�p�i��4Q�C"O����E�&�u�G�C9Da��"O04�PL�I�Y�0��1A؁c`"O�)P�&��A	�e.F��P"O.�H� S760��ǲ\'�
"O��(U.S'��� P�<!�"O�84 �N��9��h^�9�"O@x� ��2%>-�����&��"O�0�C��60�$9S��~��г"O
P�h��0� H�!��$"""O�1��¯]��'�.��y�"O`�� e�-$�2�)WdL��4Ia�"OZ���GUC��puB����A"O����W(\ΌA�
�S��da"O� �O�Eď�l70� ���"O�h�dMS.�b�z���zy�5�"O8�mš-�ȩB@K����mʳ"O&�۷"�5'h,��
�1�f�p"O���'�o�&JDǒ�8̰�q�"O PJf� 8�:EO5OrA#@"O�5"��q1�x�ţ��Teڄ��"O�HB�Ǆ1)-���1-[�-L8Ԙq"O6s�O�=S�	�7��-8|l�"O�zGi�j�D���*7�y��"O8�Ѵ��J�6�vǘ��Ի�"O�
3/�8s��J���p�V�a�"O�1Q�k.6k�LJ�Ƽ+�6t�b"O0���+'!bej��޼3�dT*�"Ol�1W�ɨ~R�<�GT$Z� ��D"O^��Ǝ]�)��i��������W"Ov��ue/^xb֦\!����"O.I$�����J�ʹPq� k�"O���CɃ4��q���o�ޤ�f"O~	��\	i?<���p���B"O�e�?�4��͖ �<���"Ol�C�����8RbG�_%�!��"O��Z�:=�L�9���7���"O(	�5>�j�A3͙#<T�ԩ&"O���D[6a�*%�"X�SbX��"O��t��2D�l��`B�[0����"Onl�e�I0.A����II6#�\C�"O� \Hz�`U�k�`���2���"O^�h�P���4��M�d�Dp�"O��, �i��T9�Z�<D����"Ov��wIF:�L
��S	2B�F"Ojt����	Wc��P4�0��:�"O���"C�w��#�Öw�N�%"O4�[��۬��=P@#�0F9җ"OX����=�D��#��f X)�"O~�q��Af4
	�s��?Pd��#"Ox��C�_l��c�.�''
�����c>e�d���x�d`�.�\ytЁM:D���&iԒ`σ
Ǿ�� S�y�!�d�2!x�r��/ �d`Ѯ��0��'�a|�d3Lcҡ���7��-��BU�y�ImD�II�Ϝ>y��p�c�.�y��ӈ/�<`q�C��T0c1.��yr��2W6l�[���)�l������y�WR^Q���2?2�B˔��yr�M2S:��"��	�
� 3aN(�y�A�l�*�S�,��eO(҆� ���0>9`P %;@m���6��̨u��d�<) �
�N�JUDH�7���v�_�<�� {ʦ\r!��4;�\��d�<����~4x �Y�Fo�3�Jx��'5��H��ғ/-� Y0Yȥ�	�'z��T����^2z�ɋ���$3�O���M�;&�H#��c���5�����2BtXz�a˭;d���#�O!�$_�d����$
?'Pʑ�5gɼ�!�D�Du��٥�U�~�N06�ΰ$�!�dZ�:e&����2L_�� '��x�{��'��I�m�j�j��ȧ�b${e$I�3iPB�I�~�v1Hb�0"Z�9s��6�0B�IO`	Bqn!/<"0�C�G�d\�D1��]�O��2H���ږ�];�i�g⍭o!�D54�f��w�þF�R0H�6�!���#��x@���r$�Z�/�!�d�8���z�k�&a�xݙYaصϓ�?����d�#p�:�/�SN��EQ2 ~!�J�T�Jͨ��W�\�t��f�`	!��]�E��!SmA�v0dQ�-�!�dt�N	��3s�@�k�A�!�Σ~R�rvi�&D���8g��*�!�A�\���(��W�pؓю_Z�!�Ęqk
�p�f�v��Y�e��<�!�*_���"k��U��]`��܄?�!�$PS����6A�����	�M�!��ͳ"�E˃� �+V�5"@�!��$w�~����VVP�a��&}!���5�ȴcE��:r.V,q� �%k!���[���J#�Z1'-�5�ǜ53p!��Ćc�=�D�?�<A�"�	6d�{�Q���L�HP�c.o��ܑ���
=_�8�ȓ�
�6$+t�h�ӧ�օd�nh�ȓ��u1����k) d�S�Ţѩ2D���r�� �4�BQe�l ��l$D� �4�5$1L{�7-ʀL 5�<D����E*wd�4�p��I:D�t��-K T3 �R� E�af�
��$D� �T(�D�6M���B�d�^�pp#D� ���׈a�=��K6�]�(3D�tH��"$
r�� \����>D� j�`^-&)��́y̤��b�<D��
iٿ:�F��4&^@�>Y���;D�� h��34*����l�?4�^I8�"O�5����%Ǡ�pq%H#_Z!�"O~P�RB�Cq���qĄ�pL$A�C"Odz�c��p)q�Ӛ-$� �"O�1c�B��w~��uaFPp"O����&��x&x#F� �,��S"O`y�!m�
W��C�g"E�I�"O���U'WqN1� Y>GW�ű�"O��qCɄy��(ha���y��ڵ"O@5�G�1�MH�	�f�򈢲"O�ͱ҆ɭTa�X��gŊ`UL���"OJ������څF�)X*�Qg"O|��t-IW؎�b�D\ L���j"O�`� A������"�u�:i��"O���eA?��6e�/F�v`q�"O�(w��X>@b��D�d{ � �"Ou�4�)G�5�,�$
���"O��)�� ?<Ĥ�	�#c����"O����$ɇDf ���hڍ 0��{ "O�	3k�k��q�h��g @��"Ol���!
|
���d�R�̭qQ�����!V�v@{U���6�����a�4C�	<<��� A͟d���%�V�C�	�7/A�F��B`�)H�
VӲB�	�}sԁj��\	�Qʑ�� ���`�@�xdʊ$��C��F�-���D�:���h\�A{e�W"�P�ȓYuƩ+A[D�^i��)�I��4%�ԇ��%;��0a�N�V��}�5���Q�bB�I$i�P��W Z�p{Ul\�J�b�?����ӫ��yg'������-�'��{b�$dd|P�F�(-��9�!G�_���IN��8��eT&sgbd-40�`��ѭcUB�	.1W(�!'t�e�VI�"S����<?	s��v���0�e�6XR�W^y��'{f�KV�t�\}[��ѱF��UK�'P���C��!ub��JA+ �+G�hA�'�����6����%_(�,��
��O�d��G�1�b��5�ށvk�U��S����	�6�R�A�-�W���ɤ�ť8[,B䉡n�b���1�l<���&cf��$$?Y�n�Rnj}��/ņK�DpQ���t�<��W&H��u�d�(��uSFk�<ѡ���SԌ�T醋z��5QFg�hx�dExO�5�C��D���sD��hOjʓ�O´2�˃Q{6`q��T�5=h�_�Ȕ'waz"& �O-Z��U��B����[��y"�U�7u t��nC|���C3�Ԗ��?	�'
�$#������})��D38���'�.y(cʁ�X�����8'��p�'c��ٓֳL��d��fD�1���3��?a�y�(��*���+B/ۂx�ިsCɀ��O�#~��gL�>̌Q�;t���s�z��M�̺�Z�28Z�l�M!b�q��/D�8P��]	��L�ǫE����#D������~�0���	�-E�i0��"D�4Yъ�]&�1Wfć`AXDF!D�TAu�Ѝd��	��h��^N6e�č4D� �@��6}?*��H�/�K$ �O��0D{�O"���'���Y�s+�5 HA3L>�	�A�X�Z�F8x�b��d�ȅȓ*��i�,5���hw����\����bXA�o[�JD tP��Ғf ��t�$D��X&E[�2?x�C$�ó�*\�d7D�� .Ys"��>!��abbŝK�p���"O�,�Q��_�z�s@j��Q$"O��+ �:@h�J�,[:z�,��d�Ir�O��A� �A��D��"L� �'w*e	���%�ջ�� �\Æ��'(T��q�?��� �S��Y�'��]���T��แbN��a��'),�c�DATG�D1�	Ħ7�`%��')���-].+f�@��.j(���d>�"���j���E�&�\!p2�X� "O�f.À[㐄ɰ�� t�n=y�"O<���<�� ����]; ɓ"O����!�B�(�����	7��zc"O.P���a��)1gP�g|�(6"O�Us��L#_:�Y2 ��f����"O��qH�x���B/C�K��'"!�D�t
#��2{���LZ!�R�|���AZ���A,�5!�^�V4҈Ȕ�B)�du��+*(!�� 2������u�Fi����.w!��z�N���'ߗo�~�3P��?�!��+m��}��E�g�Vz��Y�S�!���\��(3(:��%XԈR�zl!��$L$		�!���9��B�Q8!��
@B��E�Α	f�h��Ļ+W!��Q�F��ƊL9fW=9p�H�	!��El^\���W?bTr���`ǀ^[!��,�L�s�]=0���#;�!�D��J�tp�Q�ď�a����A�!��N�����J�^v�U#�L�n�џlF�$E �b����V�B3Pzx��cҪ�hO���i�!E��c�C*XF�����!��>8�P�ф,�0.���N�h'���'�����Ą
�F�h�ů5W�e�e�'�!�d��=����4K� .T"��L�q6!�$U'Xꚜ3`��;="���u���x�!�@/Z�쀆����8"ś�z�@��?��|���4'�J�sT��P�
_�����D<�'Z�8#��N� ��-	�b<ܘ�ȓ}�]䂅!�d��U�����	�<	���#o�Eɦ#����Sp�� ���j	fL��ؾ�2`�p-]�DjBP��Rw0%�1�A)(�L�I3*�2xb$���;J�ɡ2�������GV�
�Iu��˟D�?������R4�P�gC�aYU�`��ԟ(F�tIG�--���̊�4jx���E���?����%*���%F8���Sh�3M�����r��B,KN�Y�,�b�> +��؇���VY�2�F
$�U�����?B���9�L��%�]�{L���aZ�b�M����<����32;�E����l�vI���ny��'j��b�	^���f�\x{��$�O�"~���#�~��򪁌_{�$��
�i�<qvė�A4��ab�Dq�c!��c�<���'`��/q�~��2��t�<Ag�W�)�H����'\VQ�S�g�<Y2�1C$"'N&�����c�<1FA|fh$:p���",<��'�]y2�'�B�K��q|��X���*A�Q	���5����re�:Pc��L���{<a`A��I�H�YV+[���9g�N�<�P�]Bn!�p  ;c_�@1jQH�<�FZ%*��݀���9mМ�V�F~�<)1ȝ��x����5hǤ��V�Yv�<� D�԰Z���@ �0"J!��"O��q� ��vt�z�F��Z��=�F��ȟpE��	�.g����5�Q3���҃�]��y+'t��X�!�J�e#�E���y�����k�醦H�����Hٱ�y��^-Q0`M#��J$BFI[����y�ϖK000Abȥ3s�8s	��y��Ǻ��!5�T#$*�aз���yҌ�$`l�BP��!���J6�)�%��g���Lȕ<!���]x��P��V_���U+��0	!��\�nqf鲒�^7RE���J�$y�!��:����g�a3]!�)pq8�'��l�+\�P@j����>��z�'ޞ�k�8`ٺĢ``-] e����'�ў ϓg�v<����w��mۣd>TK�=��e��˓'\/w8���۶7��ԇ�T��)S��5I|��P�.,(���iXN�(�A�v�:q��l�Z��ȓ������(�i��\({P@4��>=��+7K���C#
JZ=�ȓ<���;���a��tufB����ȓ �M�6H�9�h �d�۝9�.؄ȓ��E6Z�J!R��G��4ȄȓYv.�3Fŉ@�:�����	r�q$��	V���(C]�k�L����!"�L�&�"D��eʆ;Re�,P`�
��x*UL"D���*�������@ e�'B$D�l�d�atR1��ìd"��C"D� �*�:��c��*r�@��ì D������im��+�BC�_\(�7�$D�#$�'o�l��C%U�d9��$�$�O�����hb���!�#O�dY�� a�!�@��Bp)�"$WP����_�M!�d�t�2�鷢]�y��B����r�!�dȡ3��a3H���d�ɦC�!�E�gh��]�Nm0��@�:�!���YNq(t,ۗ����*?;5!��uG�bW>_��p��^5/!�ď�vM���a/ T�8 �7=_!��	�b_��1��A��dd� \l�!�ߺ_v�����C�X���=q!��]�[��z1/֧'���h�/�R^!򄒝l0�ĉ��ؒ$�NP�p$Yq+�}��q���p�f�SG��#!N�B4��OZ�D��'􌘛wTFɄ��퐜"�n���'�Z�(�A��,�����I�z���r�'�ax�
C�z7 P$k�>y���PH���y��.���-_�o0�#��%�y�k�1����I:�@�@7�ʋ�y�6��<��ڌ68�5h�K�7�y��ɚ8ؖ�s7���/0�b�G�#�?yI>�������IG��\��	32�x0P'j�-cfC䉟jev����Y.&F��0�\6��C�ɍI�F��&aX�wx�) ��]� B䉉\��i��f@�HB-+�B�	B�.|�I!r(<�:�&�F�xB�	 e��x���/+����,ݤm�NB�	�B��lQ���="��������B�ɋ1Z����?r�D;����B�	�.'�,{�L�5U����ϙZ�2�$��I6>���R3/�!��s��
/<U.B�I�X:*�xSEӎs@��`jԯ2�B�ɖr����aE�;�X��$��B�)� �� ���&  ������Z�T��4��p>�9�k�1�PC�%R�N%���5D��Em?&|	`D\ryء+4D����IN�Bt��3[zi�u�O�=E��$���xI�Q�¹q2��#s�ЛS�!�dԅk(,"�A��$+~�S� A'w�!�Кg^��D�:��I{���
�'���Rj�q���[���YvZP���D8�K� ��g��=U$��FiJ�~r%�I|�����	P(�|�v��.e�#ס��^��B�	:R��t�XQ(E�R�6TLC�I�5i<¥mW��<�[R�ћ6݂C䉀g7�1i����	I6� ���}xTC�	�p��3�G�Y9�abc Դ>�nC�	�r���j��x�ވ9�͵)�T���7b^ze�Ch>	Ñ���ee�L�����*4L��T�Zf��2z[�5�ȓ\*4�j�-��:���f�(P�J�ȓo�*H�C�܂ ����Æ�PAL���x�$ۆ���]r����Jb�,�ȓT�!Iœ�a3|<��IEML�ȓz�T|*Q��� �r4�A�݋a��5�ȓ,n(�v�4D��`��ET �dI�ȓr.0�'�Ή'�������{b���ȓ9r�� В<\�l�POg[T�ȓ�RɈE�^~��[�-�=�n��ȓq	�z�A^���k�)]F�(]�ȓ_?��$d܆S� IG^Id�ȓ�: Xw(�fu�Y*A�6yڽ��Ie�'"�]�`�_fn9�t�G5h��E��'�N8����4�D9�LD#*�V���'�X��W P�Ҹ��V�4HJ
�'�Y#̨~�Pw�G���y���g����E
0� J��y��M�2L��㥡�?��p%���y��6*t���珖n*���߰�y2�^�!<Ȍ�K��e<8Q8����y)MEl����)\��]�դ�y`�U�U�1J0R
Ta_?�yB��CLf�B!�ĆX�\s�H���yb�_�x�4� ��:s�������y«�;�l�x�C!2_���允�yr铭=8�e锨ִ<�����&��y�&(��\��I�;pA؁��8��'az�CT�}�@�8�(��]@�1�-O#�ynHA�a��/D4����6�A2�y��ρy���%)�ҵ�����yr,�nl&���gp�XFh���yR�&h���[g�N�an��ӫ�y
х]���H�χ�f.�i��ʖ�y2(ýu��*��i��i#sdձ��'Paz	)p�P�Ɲe�hL��n
��y"F���Lr `�3a��
QD�y�0�����욵p���8`��:�yr+�2�4��j=d��P��ڣ�y2�!	T����"ѰaO�u�&(B��yroSz�x��!�/"`b�a�mG+�y2GC,N�di��˕�����$H"�y�@&�HAa��HPfh��P#J��y�� 5,/~<q1��PR�Щ�)�(�y��I �<I�P��K]��r��Q��y"�Y��R�׫6L��p���X(�y�Gԫm�rcHҲq��{%F!�y���(}���R�\�J H@-�y
� �-��`��ijz)�eQ�w.��"Op-{����+�P ��)m�H S""O��y�ݫhX�04�����"OZ�20�ےWBj]㖪����'"O�+1,ƞmũYh8 \��"OpYkP�9W����� ��ۅ"OB�K�� �C�9!���)�B�(v"Ol:E�<7�X [&�"����D>LO��P��ރm^�Y���  ��M��"O��q�]��θS+�&Φ��'"O��"�
L��2��5G��4rf"OV� ��i������
)u�� �"O�5ImC<��R�f(8	e"OU���(i�B����9�DQ�U"O�I��l��/a�t�EK��E�Ґ��"O�Q#�LQS�Z`�j����A��'�r>O~�1C�ھ`��9�	޷/�<@H#"O����1o��A�t��m�����"O ��F�R5-��=� � e��#�"O�/Y�(s��9�-��qQ��"O
5Q⧄�$ߠ�� O�<�yQ"OT��RDҦ#��EH��������"O$j�i_�3,�a���6!��щ��'�85���[�"��,�/=49�'r�a�lG�rf2�h�=w:��	�'��t�4M��V���ZSCO**&�PC�'�h㶁��W.Tq�&�r	�8��'uP�	�@�#24�� ǽn(�L��'�rMѥ�*�I�W���T+�'6H4�R�R�y:Z�;)�� ��#� �^�e2��_{�a����+��B�I2!�h#�Ə4P�޸`��k�FB�Ɇ ���fe��j|�sө�?�DB�I�U���R�ڒA.�q�&'֌)q>B�	�-�`$�!C&4�����!
��B䉦B�>�C�!]�>0�H�E�*xI�B�	:��8�ǔ-X.j�ǪF5�C�/ �KE�͆s�D8�!�)[�B�	�����$��"��VB�=z:�B�ɐ_�Zը�� ,F�$ �럂<=�C��>\��]�"��4�#TE�7:#�C䉨#���yc!Z;�`p��ƁY�tC�I�z�2���j@�c}��rG�P3
�
B䉵�����ŘGM\���&�f|���?	���?��'6�~�Y�F  0� �ЙB��4��u�j�QgG~�!���e�4��*��HZvd̸<��W��� ~L�ȓ[����"H���Qyɛ2T�n���C����֐��Ip���K��7rĈ�U�8D�,��ȭ[����fZ M{�(���#D�t�H)1ժBfY�H�n�#�&#���Ov��>�+C�+	y��E��<X�{�� D�\x7"�>`Y |(�$ �G�&h��	*D���DoS6b���;&ȈR� �D(D�4���~��8c���@�r&�%D��[V���Ki�Q��Ņ����D�8D� ��֘L~^!a	�c2����,D��t͖�-p�P�C�jhd�0h.����G����		�䘑��"D�<��1"όUl!�$Ru����$�-s������
b!�ʵm���K5B�Q�Z��w�+Q!�$�mi,$)!��nQ� ��:<!��0I0�@&��08 Ud�<V�!�=�<�L��I�P���P�!�� &J��J�)Bth�(Q�9X�3��'��T6eX�H4\��"�N+
��-���;D��)!����I����5Q/�X�c�8D���A
4`�-X�O��JКq�8D�p�B?]v�ZF2j�P��ѧ"��O���J㮀$R�]�q�Q��H$�+D�Xr!�3�&�c�õ/��p�F�)D���MW�lB�4x��Dh^"Ppv "D�����
#xyF��D;V,Ru�u&>D��0�ֱe�fIXsf��	�Xĸ+)D��g$���,iQ�0u\�I��(D�XPWM�j�FM�a�v_(�ҁ�$D��a�jJ�L�e`� J�H����<��	vBH�#\8��fdӄԤ���I�<Qb�ҵ�7-�h��! %�hO����Xn�0 5��%���C"��]K!�ā'����o͈@�l��F˙�-�!�$��.v��JC�S0�
e�'�]�5!��˹t�m�р#:uhwH�j!�D\�%j(���h̦"@$h�jQ"z8�O���)���Q@nd�2�˰�� h�j�`a"O�Dx ��JP���Õ7�Qi��'��0��IT�|-�R�'`Y��r��<�M�B�Õ��I@T�`����d��b�h��Ť�
Y^�� ��WфĆ��ß��bk֌9;tir��9��IA���ȗ'Tў�>�a��H�s7��Qo�_��<s"�<������(��IX��2oT����O: 0y�"O��Ŭ�!O0x�����1v���"O�y�$'�
�ƥ�DF �t2���F"OᘱD^A�N�Y���9�ȼz"O�D��lY�	�FD��7g�8d�c�'��$�IOH+ѡ�0X�����/ln�X��D{��4CF> 9��*'��p�e�J��hOp��	@�i0��!�f�)4*A�� _�:2�O`��<ђ����}����"OR0�	,QR���D��ȥ	3"O&1AB@Y�^@�A�F
+���@"O­z��խb��x1�ehM���'[�,Si��\�.I�b��x@VB@Ht"�|��'�O�v馭h��P�+~��¢o�x"ą�g�'  U[��Hb����}����r�'KP=3�� ;:���ʶ]'����D ��M�%끕Bj��c�*8�|t:U"O���:*��+�eH�G��%�2"Oܬ��̙�=�Ptb7�� �:hI�"O��j�/6�
�B!
H�dU�ɳ���q>Y"�U��0��1dP&Wǐd ��3D��RQ�R'}�F�!��M���c�`2D����X�eJ��Wɇ�7�~�@P�,D� 0Fm�s�X�u�
;P�p�6D�`K�iL�,�>QkI��)�@�B"�4D� �G��H��[0� K*��3D���BB���0 �0lƻD��q!>D�Ԉ5n�)I4&��!�0�����!D���'�k����5M�! V��<Y�~�&\���ǈg��I��q��y҈�z�\�����9*�X��ҋ�y2B@"��]jN*~�6m�:�yR�8r�j���G�f���h���y������ ����cb)�y���c-���DQ(tV�ac�hH(�hO.�𤒘>���4�,>+*d�ux!�$(�*����ܷD :����)8�!�� 3�i �0CeQTֽ�$"O�}i@�_w�<�Ӆ�w :M�"O.�S'�����Ƅ5��E��"O�Qf��F��MS�����8p"O:D#UN�#;�����D�4b4���@"O6��N7t�����ӡ]��6"OR�I&�-V����/�&dA�"O�S@��O�����8�>-�q"O6=jDG���B�]04pYj"O���BG�	�x�qpb"B�p�"O�c��ۙrch�@p�J@j���"O��x1�s�"h�r��,�ʓ[�LF{��Y$J�𸗃 ����9C	ȴU��D�O(���O����O">Y���hS��(&� �����e�<i!�C
�֖��R�Q��[�C䉛[O�|Kr��m�
�rS�:�C�	<o���-���xIì��<~���Ofp��醤HYҭ�r)&]�`�HӦ7D��bX��ue�/k6\X$n�O���OB�O?9se闕h�Ro�S�tБ��l�	����	��x�	P�'�Ѱ �W�V��&n����'v�R�
�1V��2��'q�v���'��)��#��إI�h�q�l��'"D�F
�c�%��+)R�`�p�'�6���Q�?64(X��E�X��
�'VL���E�=�ba"D�o�l��)Oh�=E�T���S)ĉ+q�;l0���VdW!&fb�'��'er�'4��sW A2g�h]R�lQ���1G�:��0|2r��.=Y�97H�a��9�c�q�<	�_Y�=���G#E��l�FEJm�<)r`��5CBHRa��!-8y��N�<�O�7{��Չ2�U�F�P���R�<�wX�猉\ĺ 2*�w�<A�E�Jc�9���	3����%B�W�<�KN�[��U��1U�<��*�[�<�bhZc��J.	�1[�:娇Y�<�SfX�Oe^! ��XN�܀J�Q�<��ʟ��l���ݽCMzp��_�<��%�p �r�'�<�>�7�t�'�a����=,�&	jd.#t�F�a��O2�=�}�3�H2�A�o�l�l#l�d�<�fO�)[Q)3(u�S�#]f�<!��H+v�T���Me$��3�j�<1�KG�����K7�<�Pb�f�<QR+�� �4���G�;�����e�<!��&]\��B��9Zx�3P�X�<����GV���$&��8��+�^P�<�$m jb�+B4P�-���ҟ����S�Ft�R�b!"�;�A�Cyp8�ȓ2��w�8;V��Qʂ�s
���itfq�E�?7t�$M��X��E�ȓDD�!�͆`���� B:4> m�ȓRSЍ��X1Sq~ #`D �pلȓ1�����䈧vB��j6 W�F����ȓu�.�R�H͍����#�V!x�
̇�b��L���W^U���O�m��L�ȓ$8�Qqn +5uX@�fe�_��A�ȓȪe+��MH�psc�Ԭv�ц�Rh
��e%��	Jn��@�{����ȓjIn`�	P6 �� ��\,Z9��xl���Mݛ|� ؚ^礥�ȓa��H��νfYh����m� ����R�L^��<uq���/F]�-Ro5D���D#��u;���*S���!ڐ/5D�� �D���H�,=�����d��Ä"O�0'L�? 咬�ק��x�� &"Oh����ɳg��'g��N �� �ICyr�'1�������2��`d%��_�R�2�"Or�
c$6GY���CϾ-~pyJ�"O��@'Xኔj�$Y�:� "Of5��ȔP���㊞.���[�"O����.Y(P^p����I�T�p�"OD�A��Ú�p�P%e�����"O���k��Su���`�Ȝ	<�9��'�X1HU�H2N���dDR�O&D�(�P��li0 �@2w!JP��A#D�9�J�]�(1��*OP�c�+ D���fLG�s��R���(�j%�C�<D�h�A��Je�Kd�:_��"�:D�0�G& ـ�3�n�),Qz����9D�p��!@&�j��&v���d�8D���&�!6,y�����o���8��6D�|z�eܽf:�M�b��f����=��0<�!Oy�9P���b��-��!�b�<1�_�^A�8��6�zd*@�9T����i׀2���/MFt\Ly2�?D�T��+v��˰���Drq0D�h!V�J����1G�|����.D���D"|~�-S�gݚ%�l��5h7D�8����hۖ-��d� [`EА�9D�dx橘�H˾𠔥��M�� �u 8D���V���0 ��%f[�<��5D�Dx�L�/N8�k��ڦ5c|�"� D�����ƹf��U�Ø�1t�*ӄ9D���H�Ǝ��i�� l����$D��K�c"Oj���$��h��=D���c'Z�"�⦭ΌeJ0�B�.D���0�z)6�`�͎' ܋3�-D� �U���V�����(7������0D���ڇ1���%�&G
��:0�-D� V�m��F��-y�|S��,D�4��F�'I2f\�p��.㘼�3M-D��0k��H%zH�4��N^`�i"g7D��9SfU⢵���J�s�R��5D������C�0��S!H�K�b�i#�7D��)�%�#/:~P��M[�r� @�w�5D�;��ҋI���J?Z����5D��3.^�gE�8��g$f�42D�\��D��TX1dZ::�H�h�,D�tQuh�3,����Q���I\28�UL5D�$s�䞙I&�A�g%ĨX�l�@s3D���WɎ7{P��sK��l�P�*0D�$`%i�����S��� X90�m-D� ��J7|�f0��
]�TY0Մ0D��(5KH+p�0e�@�Y#Z�"틗c/D�ث4��]_����K�e_�P��!D�T�J�-�N���ʥvT�Q�`2D��Ţe��C�%�@*���b 0D�`�5�R?@$��Fk�:� 苵D+D���7$^�9Ũ�"�'	&>�^]���>D� ʀ��Z!�a
jF�`�@-xO>D�p�L�;X���=lZ½2C:D���U%ˠ7I����MS��jw�7D��2"�*���3#�3�jA�Ê7D���0A��`� G�M���6D�4s���6)��I�Z�؊s!D����JΚlؒD6�t�Q��2D���ؓo��)�RA���j���1D�� D��sE�#p�0p7���Q��y�U"O�p	���9�qaօ9s,Aq'"O�93��-����q�07� �"c"Oآ���hD)�,�5`�.�c�"Od�jTIg�'�Z
px;�Ñ#�y�@Ȫ.Yܵ!��2��5�SD&�ybB" ��G'6.z6])#�2�y�"�H��.�6��3f��yB�J�oS@|��g�J@���y��B{�&��_��tx����y��Mm\�r�J;lm�)Q�y�D��d�5K��e)T��_~j�ȓ?h�H�A� Բ���E�ڨI�ȓ+��<�3'ڴ�(�qe-̫Hr���ZK��@�-G�z��3g
$)Id���_C�H��X1�P� t���[:.m�ȓ1̌17)��4�E��ǋ2`�bX��4�<h�@�L�y���"���؇ȓk|1�cj�Ĭ!�,��	掅�ȓD�t�c��4hX&,i��v��ȓX�$ô�O�'�"� �쀲Dך��ȓ��0�É��J�%)U�;aP��ȓE\�m[�k"�MP���MZ�E�ȓ+F��)�#�"�k���f�:|��V7l�u�خOg�-�0�-�t��5��4	R$8RY�G�Υ;�����Y���ǋ]3� ��NN�@9衆ȓ�Бv� p��5��a��V�%�ȓd��)�Q��&��h-�}ԅ�:5h���K�Yܐ����N��ͅ�6�h��]4�=x_c~Esw"Oᱡ̅�B��iqV`�iOH)s#"O����L�b9����8B\�"O�T��l�T���&/]�g'���q"O\(����V��d�V�W�Ƶy�"O�`��BO���1wo^=z�����"O,-��&�+6�*�@\�3֖�CA"O܌�#�ތER��1O�I�bL�F"O8!c�	�!���s� � ��%y�"O�M��)�o�|���\����#"O��Q�4hx��	�$�A�"Oz4J#kj��͠#�B�%�q��"O�y�_5vbX�SIN,(�@���"O,��b���Dn (�P�ۤ�~hBp"O���v�4�R�Ӆ�z��pr�"Or�0
X��'� �Μ�"O�yS��7 ��@���3F�\!`f"Oh���9�$q�[�l!�C"O���%�C���;A��'݄���"OT���f7Aw�M��B�g��b�"Oތ���^ .��|��	�w�P��$"O��{7c�x&B�c
�	>�P"O.p�t@�M�Řņ��4�<��"Ol0�S!�����r��
T�4"O@S�qO�����[��E��"OL��w,_�#�F���	x��B"OZ��!�S+&e	lˎE��`��"O�I+�B��y�EY�j�,!L�`"Or�ر�ΰ<z^Iŧˠ8{
�B"O(�ɦ��-:D�:���(H�t!�"O��iF-ŉp�da��g_����"O�l�e�]�Sq��+cG8%T�d"O������/!0$�G�^9���C"Or���'D�3��r%��=�D@b"O� ��22e�!V��Q�R5}J��"O��r�n̽A]�M�&�}X���g"O�xC*.�$�x��&[Tz9#�"OXp� K��+E �Jç� �"O,Bw���{^|`�רQ�6d�!�""Oʕ2T(W63�q��$��3/X�0"Od��!V�Z�Z�Edr��"ORq(@��w��m��DQ�5���9C"OT�Y�5���8�� ��a�"O�D��q&��Պ�GkJ]*"O�A�a �B�>�TC8�i��"O<��� P!T�\H�EB��NӴ��"O�A�C�Z�N���Z�ȵb"�A3"O�T�5�S�H4���C*	@��G"Oi
�j[���9CQ���s�j]��"O���qh�����(6�I�"O.�;d��!~n��
`.	�o��<G"O�Ƀ�E�o� �9��G=!��$��"OT�Rk��P.�У{�RVp�<9P�ӷ1%�;��޵}�Mi�%p�<��l�:8�x�;+�}��Q��T�<q2/��]Tj5 �"ϯ%X�)�N�<�3�ǚ*�=P�(m�>�A�kFH�<��e�9���`�K�f�2�o�M�<���.R�uJ𬟝!hl�j�~�<��?��T0�͘i�|����e�<A��7vg���r�W�yV9CEn	]�<ɥ��Tf�A��^�=���"A
�M�<�����@ƃӘ/,ѱ��G�<)BEMQ\�y2�-"j��!!IG�<�g���C��K�HM7q(�(���E�<Q�*-	)�D)3 �>m:2ؐ��El�<ya�**"ʙ	C��X���<ɗȼl :���g$����hc�<��J%|W\9��Y�:�㔃_[�<y�BR�S�9���B�:hKQ��[�<q�gT4~4 P
�ˇ�}��ف��M�<��D�5D� d"�F�X��SA�<!���5\��"A	�Qv��g�|�<Y�/ʆT�p�K���,��u#1D@�<	G.Ŧ
ά(
���H�.ia�<Y#� 3���r�V� �[+g��[�<y�c9,��ͨ�LG4�R�����[�<i�i̩5R So��&��Tx!B��<I��� ���	�U�rtDig�<�go8y^lIɷ��,w ����H�<A5`�C6~h��#�$+WJ�#K�I�<��.�qP�iw!�	#����%�Zl�<Y%+U�@3*x�`ɱ'�@�<����� �PJ�	��p��q��Mu�<�7HF�R-R�p������V�<1/��*�Ұs�C�n�<=�eZmy���v��J>��	=q����G/�<e����<�S�G���$�j�cۜ�S�(f�����H�8�I�bC x3���t�G���	��p>�Co��A7�� ���2T� �Ơ�R�d.�S��	�>ᷩ!/���񌅓ښ܈�-N�<i5G�, �"E��zed�qV�#Ⓚ�\��%�.��x3� 
��`W"O��bEe[.�Qj�+��L�P"O�E2`�,U��%���Q:H"D[`"O�Dӊ��9�� )wF� "O|�g��K��D�Pb+�u�'�	_8�(ӱ�͸ �l�:T�K�`��;�7D�� �q��k�U;w��(��u��iQў�E���A�a���Ĺ"=��AD�����>���<I���Dz[t���nJlB#c�F�<�rG��9q8!�CC
�#&h�� ����P�=a�Û����'S��	��:@�'*
MBلȓN�l��/֧

v���]AJu�d�'��O��|?L<i��yi<���D6�v�#3K_�<e'�h&�1�&���u˂��~�<��!���zg �,%����#φ}�<�%ɜP�F��C`']!�x����t?���'$��t ����K$�X#V`<	��(`��� ��de��#��"\}��8�>��G�Q�� �to�:zP)Fz�'(����[�g<:��ա24�	8�'gdq���Z ev�W��7�%��4��$1�Op�p��0t��h۱(?Pz5�|�|��'�.���fS��&lC$��Ĉ���1<Or�bpG ��>9
1���cE��y�On4׭�	��3�¬Bv��H$ˏ��>��'�	J1K8d��b+��SLD9�S��Py�F�o��U�P��*YxZeX`��\�<�N\�~�JC�޺Q���{5�X�<!��/��e��
N�Nj�X1�i["fў"~�I�j����k�A��f^�a8J���>��@���.����f	rf���0=	N����<^����T�r�
R�7�O�O�Đ%�C3�l���	�={N�;d�I|���i�*!.��`Β#$��Y�&$Ä1�!�d٪>I���Ćl��cG�ў<��ӭa�̫���L�@�õX }�,C䉖!�05�b��2"��(�Ⴠ�UIC�	%J�����hN�\�".˱3��b�L��	��![Q	rn��:�Ȭz��B�ɹ|��+��� ��{������O���?�L~�+�^@���^�fyp�qt ��]�(m���t�O���F�ΏHQ"�#��ۯD�p|��{"����<іƑ��:	>R%P)h�&t����?��A�j��\�AH9	:n��q��x�&R�{6�g�Pe��1h'O���yB-��l�F"§Hk��v�Y��y���
����CE^�U�����T"�(O"�'���d'P|�9QD Y�BdR53} !�d\ql�+�*
6�zQ�7���!�D�?pj���D�%!ފ�#�,I�n�!��?dQɃ���!H�Ȳ
<$/!�D����ꧨ�c(�!�^2OA!�DS�K�$d-�M�y @W/q9��x��8�PJ,+>��6mB�~�(MC";LO��O���Ϭ4��	�Ko���U�2�!���:�L+��D�Mm©U�L�9���3���(%��B��^Eʀ%WoB�8e"ON���O�mNq$��4��+�U�D��'��}h��h���	b�@#�4����N�J��\P���m8",#g��`�V
O����X�J�pT#�*|c�����'�������(P�@c�ġU��@�/1D���*��Q�b'B�My��i�L1D��P4	�wD�݊�C�,/ܼ�C�/D����'Vg (]Y��E2e&���V�,D�x�V!E�H ��A�4���&D� �B�ƨ4�D��K�9H��Ѫ%D���Kр/iv	#ݶj4QY8D���SjG8'H����/ip.=��N4D��	�ǝ(������A�X��(p�L2D�� ����^�`]�v`�<EZ�@��"O��c��I�G��0ȳ��pH�� "O�<�4Ξ�K'4Q�#��]H�)W"Or�i���v��Yu Ǜ	�cg"OFcE!Z=D��ѪQ��=@����'��	V��R�^N�<p�ʚ/��">����,@�ΩÓ�F�6*���� 1%!򤖶y����j�� �З��I�5�S�OJ�U�!+Y	t8\X�' WX��'���4�۳(4bIx6�
x&����'��d�,/KP �5`C0t
�(�'f��k��^E��#�I�4�]���D9�S��I?S�53a"�;\�&]@�㉤�ynI+S� ڳ���jq�a(c!�9���p>!��� /��ZQ�(gT,hǇ1�D5�S�D��O����<�-�fN�I ��8b"OT�2���(Ue�/z8 ��x��$IJ�'�0y3��	��q��߄5u(�')��`�&���P�I+l~��ˌ�;�	V�4MQ�g-,��愙��T�v���yb�6_(�)�����А�H�?�y򋈝f��h �K���ݨe��1�~r�|r[���ʧ#�t!�枹v�0[�͆�npB�ÌK��������#7ޅS&EY�_�`��FLE�p��L��?�"5��"�L��&S�[�� 5Fw��B�	6w�JL
7N��J�����l�=���q\L�q%˞Vg��'ʛ0�ў,G�T�i%��s���a0b�:�뇯I��c�'�4݁cm^��m]`�%C#>]<���2�S��"�# GTQ{E�" ���؃J��y��Y�R��v��%a���� +�5I�v�=qF�i�����C*Q��@��XӬ�V�<I�L�dS@ SUgR*�2]Pր�m�<�ざ)M�<,vL�����a�<����9�4���$8��3.QX�<Y�^7f�였"���	�2�i�<�!C/]�*R�J���H�`}�<)S��>Q� �B�����u@2Hֻ�hO?�I?	>��g*r/�|r1�C�	35�� P�Ž.g�@��^+Pp��P����d�����eN�3}�ak�(��0|��E8I�c�FH�p�F�H�'=�xr�4>�$�JF��5gjmYN��yr)żo� �V�ʥ����A��(O���$�M
,h!�,L2=�7�ޙ3�!�D�>a��hh���9����C-P�!�}���h�Έ-Ҟ��˳z�ay��	,k�A�HZ�PeK���9��"?�q�?�'�X,1&�@�9o�����ڞg�l��3�t%�W��M8��R�;���'��'U�?��WN	L�8����ǻ<�|{&�"D���-X�I�.�� F�[`h�
�%D��� �"���N� Vu[5k%D���t!<;�0g�׺r.�IG�6D��Zud�,gd��k�?n��$�*D�(�ʟ�����)�4d�v�z�C)D�@xOT�\���GK�c�R`j�m%D��4ł�R��`Cg��CNPz�-)D������S�|��ՃS$��ׄ,D�H�bA�f�T@`өT�<(��+D��gO�	�a1�㍣��q�6-D����!~��3��Ԯp�a5D��P��ŉR;�b�C@���%�5D�����gX���6"č'��QCH?D�� .�A�狒d�| �D!ɌP]\�"O��j��%

�u�� �@?rq�f"ODp�M�/"��w�H(78�@�"O�x���58�n�IE�ۄ(0� d"Oޘ C��P��Qǁ5;�U��"O:M�u��\�Psd�E�jH
E�f"O�D*��J5AT�]�׮�f@�q�"O��r�)Ƕe�y@Ӯ�,c6���7"O�\"Trf塡���1!J(J�"O�`�2��0�Y�P,�+T����"O�M�c���*
�u�$�ƈ��"Ofp�fj��D�fa�IH����[!"OF�ҷ�ē�pxPM��Iz���a"O���_9�"��#H8+�.r�BC�<!T�W��|�;`�8_��Щ���t�<)gE]�p��QׁU�t�h�7��l�<i���#Fʨ���'d����o�<�t���f��q��%I:\��)�k�<���34=�� �^�Z���i�<��\ ?�j�8W��:
��Б(�e�<���D%9�|��0E+�� �$[b�<�ԀB7Ɛ3C��&gJ��#a�Ra�<i��޲~T����ޥ0�\�3GOw�<���Q�j���d�D�L����F	p�C�ԋ��3O" ��F X�KyP��<��%�on��r���Ҩ3r�RG�<�"ڮT�Dd�O�B�
���g�H�<���ԫ���c�R�D�Qe�Nm�<��/(<買�*vf��7�j�<�qW=�NpR�h�!u� dV�e�<y���+
�l��-��=o��І�Ay�<Y��٭JA�Xx��4H `2'�^�<�W��mZfL�`ԬH���#�MM�<�A��h�������{��-�AK|�<I�F��&�t�%#�5'T�4k�JQ�<��G\%2[J��S$�6��!�$h�z�<�pSr����R��4��A�l�<	�+ѶtU^12��ߋV�(����Ov�<Aԩ�pv��R��A��b�����q�<���J���\R�M'<:`y�@,�h�<1���G�2X�6���9�D�sq/�i�<)q��d>�M���4X��K��M�<!U�'>Ѩ����ȖAEhȥh�I�<9t�Y]vԑ��_	V �+�H�<A�m��
E��&I�:i�1�eB@�<9ń_4v`�U-��;��[��@�<� R5B6=���1,�j	p�A�<q���U9��u��h^�0� {�<	4��# NPQr�,d�� �l�<1��&<""�E{!ŏ
3��-�ȓ!m,+U��yW$����Y-8�؆ȓ[��iI�/X�O�M�Ŋ��!z ��ȓZ�&���b�v�Jy��ʚ�U����ȓ17B����ȟ��Ia�F�!���ȓ,Φhx2A�'�%JBOQu^؅ȓ88<K���<�)a����ȓ?�Z(�G�����!���]TX9�ȓ?WXa�)T�#���&�LN@|P�ȓ B�L@#gͣ5�=[$��I�6�ȓMc�K�&(1�j@�#���P���u��+��H��ԑ{������6e8�9/l�9!���3.�(ąȓDo�� o�'�i�C�I���ȓa�ڙ��A�w,hDP� �#�܉�ȓ5�5+�M�5`ʈӱ 1bhh��S�? ���iE�;g@�a�m�,= L� �H�p+1��� !���1%�*o��H��G�[��B䉏��U3���"ؠk'ł�,�찠���P^,�O��}��a����*N)S������	[��Ą�3T�A+;�JAz�$�`���l�q$|�1���J��{��I%od&x�!o��D�"�;�%U��=)��tl��:�!�O\��ri�
|
)��|b��U"O 0J��φ����Fŏed�92��٘8M�dX0H�/�h��A�gj�
�)��
ϔz�\$�1"Ojћ����[�b  �ި$� �����>\^�e�U�&}��?�g}B�:,fb4��.��=�p����(�y�FH^������.����Q����M��+0&@�e2|O�|�3��'��X�D_�!$|qF�'����E$D� �b����Љ�KD�X�dq5C@b_�C�ɠa��£m�|�@҅�@�++���7�0@�.�G�D�J�V�.��k2��'H��y�!V� "�pq��e��x�0�Y�y�m�5�* �K�B�>���ߛ��'>�$��&Qv�O�ވ��͕W�n��HN�.h���
�'C����HʾzgP
se���b�J���O��:��Y�|q�K�l���a�mN�(�lp!"#D��;ׅU�8w�<�e*9�2�I�&�rXT�G��Z��|�%ˡ-�FE�T+L�-K�b�ć��0=�Uf zj������,�8_�����˅��c�<D�ԫ��l�4�4ˉ<:�E�S�=�	�8�uɓ�<8+Q?ycC�ނT�(U�%L�`�J��=D�ۅ��9��hhpgF
8P�(f�T3ZD|��a�>�,k�����/dFD3�j:WK
�JE�S�%�!���z�zTc�G�1N!��.�8E��-F6p�~��1�3!��O�.�y>p��i<l��<���8Z�޴x�GI���r�'�ٺ��K�'�Р Q�ÏL����J�.��@��:j]� "ػdH��=!l݌0'�D�5I&>(��I���0s�L�?�0��������G'��,F~���`6�	
.Aj�� W�aK�>)A�@T�H@���艒6���
�A�\XU�td����0As��Oj��Ǫ0IHS�	�'t	H5�҆;��5�R���;�X�g*�cZE��ڢ(G��<��OA���Co%}b��7hBd`Ã�7	���$��,�vć5;4HA��K�uC��Aq�A�iAlp�フ5��O�8`��fC� a�K^�pW*��$F�$RVd�g��IY��xY��ș'�v��nK�z��0$���-pQ���"&*���NƋE�8�iN���`HJ�BR���'H\X��K�����5���a%G.�Z5�ЬB�iMT]z��h����,��.6�(Lc&-Al�<^��B��6؀��Զ�upb	�83D$�j�h��8�K��ğ/O��pR�'d�Tҥ�QF�% 4�����]�T��Y��n�'}���Y��J�X��u+Ŏ\��`�J�'<����ڟ.�B�F?[Z����$�0�@�G�z1�í-M��O�2ǚ�۸��S($2P��>^�n�
@A��J���Gݒ[��Ė�����_r�%��!
<[�|�Z���\��`�!L��u�W�R%8���II�u���`B�q$��?K��]j2�ć�0�� l<�Ð@�CW�ejrї.�� j2������0=Q�bǶ[�T��"�,{�#1+I�b@�@�>,J��2G����D��
�]�
@ã��.y�Ak��-�)���6eX����j���*�U�ay��ˀr:��&��)v�ߢhک�喾Y"5�`�� [s/Ё7�\�2+_
,�����26��SZ�\x�t$��y�`��y�nQ�,p��0F���i^���H,�)����"
��!�>5���E])%ђ��hAK��ӑ�ߝB[܍�mȨ:���d�=>���@�)+�=��n�ֵ��C�~�N�T`�q���M�s�E�"vnu�R9P��w:�"�ժlba�ܹk����&�#)eR���F�5������Y[�uH3/��p@}(��_�,��y��1��*ψp�"��A��4��&_����p�(��Iͧ
@m�t���1g���PH)ι�ȓn�j�R�bR5����$ߍs��<����,Q)JE	%�M�F��P��a�S�Z����.�>y%	_�g@\��sG�"K�6L���[���ae�߹&T���g�=^_�A���$-fxqraT8w��ەE�yl�h�%��4x�i�Oh��+s�ޤz��觋&�i8�aBO���1ZT��u����i�uӱ'�~��*�*"�T��fj1�O����O3K,��� �Q�P����\:� #�ЙR���A�t�y&	ä@��$?%*��T�m�I�٨R�L!F�#D���d�2]� H9��	J���� �^�Os1˵N�#[J���-��	��c>���.?�d#*\u�a�Q�('�b��U��P(<�D��vht��ԈV9b�^���)N�nZuq��G�I�n�3��5�O�ez��#Xh��&��1h,���'Yl�,��&�r}
� a�ӳ&�d�	��6V���B�O�=+��0>Y��6��A6�٤oY��v�,I�C;扷-i�#���w���2H���r�Ai���5D�p
pb¯&��"�G_<D��i*3�3�I:L`
`�d ��^�>�" DJ��P���+�h���#D��X�J�w�)-��P�6��]�z4	,9Ҝh�O��}�M|��:4+:�����ț�<켼��	�"������C���h�H'_��xS�"-��O�@�e
w؞8SA��;!ℨ�p�+-�4d�� �I4]
�
�E]~R/Um�0
5`ʺ��D�(�F�B2OӾ "ɫ�@��<�sLX�Y��)F��?�@�Z4=��{�N]y"��l��,Cf��V�i��@3U���կ�f(h�L�8�!�d,hD��"T
H���P�>1��F���bU��ڤ��̃�Ę�-��$i�ᚌN�ȹv�FN��z��~����'S'b��I߫|�|Ԛb�K�&�jh��P��?�Wo�,*���C�&lO4�PG	!а�@d(��cu�pR���09�@I!ĻX�L�l���1�Bɱ��b�x�(P���G��%���"1�B�I%��H�	/#v�;B��r��}2)�r���
�C#p�g	����@�I�/"t���9H��!VYZ$s#לOH�:@��&ta|R�Հ� ���'f$݉v"�:W
ݛ2�� �3�Ҟn%b�ɳ�Q�,�A!pK�.3f ͹�b��?_c���!�(y�֘�g�͸
*����/�	�V���ɡ�P���ԚrZ((�-��>�i���(~�A�e�L0����L�W�d��BR2`�$�'��ы�O�_q`��!)_i99��j��@�UGf���cђ<����1�U�^ul�ȁi�o6���|��YW� '� ����C2l?�����*D����N+�\mcm��A��I�"��L�n��B�U�5��0t���B%��T��)�D]bÍ������w0��c��L�@$Թr�M"��'FH�{��''Z�l�Hcb$I��N�D�j�c��?� ��Ħ��C�� 4��28�ȣ��?-���`���͉�	AY"@����#7����?i���:#�C��<��M�V���,N�P�h�`�U+$t�0Fl4U�q2G	@'H�"b���=q���	+p�(�J��a8�� z\��V� ��	���!B
�\)���,����GG���2�<��6��-T�&|�f�E�<Y��Ю+�l�I�.MA(�1�BG?i&#U)K�|i*")O��60k��g0V��D�&����V��qa��&|���"r���s:Ĭ��I�bh��a&�3֦� pG�s� .
<�{ulu��ҁrC��'�Zs��P��G�(:�:@�7X�X�s�l0ʓ�@��'�Q��!)E&�Z��4b�"'�u��Sf&x�e�q�<%%��H���0�)P�e\R�(2�6D���7� i#�Ч�řZ�XPie�5D�L��i�*Ұ����S���5g3D���'.��Ua:	RIè�@���2D�(
Ң@�8�P@��)5NdٗI*D��$��7$8<�s�]�4����%�O\��(�H��l�^�aؒ�u��
�'�ڵ�BB�:mٰ�ςB������/b<��I+S���A,�.�>�醤ڔr�C�I<+�py���:*X���Y�RZ����<�A�򍍍y��{>��������4Y��(��D��Ҍ~�[�cZ��S�&a� 
 �˙
�hx�O�&5x	�Am?}��3I`4�R"Z~��1�J�6�$��#��Z�=3׌=ʓr��!�A�*�	9d��x��ST����F#^��0�;�P2V�(�h�OأeA�[5D-��"�[D�G�A >Q���䀟.B�ʁ��������ee�9I}^��&�ǻ@EF|��"OvBB!�T��y����7G>Ax��Oڭ�	�ک)J��s�aZ$1��`�S-,,� ��o�z�L����'M�q�o��<)p�#-(%+4c͹�D�����C�$ƛp1Z�8�)���0<��'����"#�=R��)�#K�Q�'8�[��d�!�^ �D
�s����D�-�n��e��.���3�'�XQP3���ݣ�[<�dx����C�"����>�Ӛ
��z�jM%p�^�Aw!�87D:B��!'��b-ܷr$:���A�@��p�Ι���?�)ʧ9��A�Ғ"*E���*��9D�c��>6 ̓ �`gN4���7D��rTǘ4vE�P��/_;�6`y�I3D����HO���-#+ݢ\e�T�q;D�� 
S)��
�B�L�2)z ��"O�A��F�q�� ���3)"(�"O̠1c I�DO:l�� -x�v�Y�"O��  ��:u�񯃂i��=�"O
�6NF)y:Ĩ{�#I?5b�h3"O�@��D��v�E g �z i"O�}���?.�V��!+���"O$5K�e�[Jt0���o�9�3"O�0[�IDD�h��#.&����"O�\���WX��i�F�H1���{�"OҜyv �5R�RYu.�{�ZQ��"O i�C�n~0,�n�)b��͸�"O�dB�Ɋ"�lݡ��8%U@�"O���$'A��/aCf���"O"�q�NUH�x��c�۲h�F`8�"O��$"�R��m��m׫=��I�"O��qB�#<�LdK�f�>v���"O �A�"�~�c]����"O�� oO+J��ґ�D&QӘ5�C"O��Yw�5O�X����;n�$ha�"O0�qdԺo]�u�0�v��"O�Yʴ�N�m��i!g�;�X�A@"O�` S��I��8���N�%��ź�"O0�+�����;�!@P� IE"O��sG&=��[�S�V�@|)�"O \Y�#�=OX�Iģ�cߢ��"O�9#���y���Q�a����"O�� u�/���vb��v���q�"OZ��ƛ�LVFQ��H)�*�B"O\�����8:�B���� O`>��3"O�u��B�~�td+@-PW��I�"O�5�B�Ç3�>�� lH�(]p�Q"O(� �+R%heB�%��9c����"On�aF�K�Pj@x�TJ�3�lͣ�"O���l�=>�у�����"OX�ۣ��"��Ā��B�z�%"O0��*b�`��<�C"O�Qr�e?F�Ddq�"�����j�"O��ǣV�/��G��f�4@��"O ,Ȁ�C?{���S�\.o�"�"O�16#dY��E��;��qB�"O�t!T@Z�m�8!{�g�kQf��"O�z��!IzZp ���_���u"O(]���ޣT��B��_5mE@@#�"O. y��Q���5��cU"OnX$D�~��XB���]g2�ڰ"O�mDC#%�H�hGLȗE����"O�ē@-�0X���& �<:ѐhЦ"O�`��#Gk�y"u&͖Rd��p"O��0D�\��pQq�K�!J�p�'�,]y�M��g��AB��(0�v�j	�'d2՘�H��ؒҳ:Q���'��=i�n�)Z�°�Ր6f��'�V�c��2MƖ�i@K1]���{�'f�����`�d��d��gͲ�
�'����%��>��ᛓ�\�H�\	�''r��50C<iz�
��FV��;�'BV�Ӈ� 3���b���h���
�'��y�G�T�*��!�P�Ģe��9`�'� ��A�8K��؀G��P�:�'j�Չ�A�I�l��Gh���`��'��X�r�Q4>�ы�f��A3��)�''8hqA%ßj�D�1��˙���)�'p������h$k'�������
��� J����_K���QM�m��(+�"O������%5И�1K�%'��X�"O*Y;�CÐh?����������"O��U�&)L
0��p���"OA�nцv��\�bZ�(���d���>����!P�%M$(�6�ވb�B�	�?��������R�ޭ]Z�����H,r)4�O��}�WF̓���>�Vx�6��m2|p��/}�Y(�BŔ~��*�K@����m�	@��b��"XG�{<	0�b6b�Ry��ZG�����=� j�1]�v�����O��Q�(-�VQ�BH�|k�5�W"Ohr#�#�T]�EGH�f��{��$�,=����L5�h�X���iN2m�TX0 �N��kU"ON��a�1� { iE����d�ş1��I3�(}b)$�g}�̆/kި�vh�!�����F԰�yb�!.tJ�Ќ̚y���M;��AD�J=�a�9|O�ܛ�HVP�4� SH��v���g�'f U��N�"R��(�ɮ	� 9��!V��a@�Y>��B�I�o��Ā���+Mʨ��w�⟐�.B۴�E��c;"���8p)S� \N��DHT#�yb���C���P�1Q<�D3�B��y�H�%p��tDo؃z�AT����'zݰD�Hb�Of@��ޢ������PѠ
�'�.��T�P$~�W�ʅg�x�5NH�ȒOpٍ�Y�(��.�!����A�����23B D��чI�B�,�T��5~j�!��^x��
:@�|r��=O*~M���t�͙5��0=�DW8d���*2��t���4IΎ]��+]�Y;6�:D�`�b��-et����"fUyJ6手%re�
ׇ.�Q?]"s(@�*� P�v
	)Gp�uY`k4D��eO�1v�����JzX,K��ճX��08C�>I�]i�����Zm��	�-�dMZ)I�n[&8�!���f��YJ�	ʙ;P�c�M:,��P�I��b���i���#l�i�fh2Om~�SG��?/�x������?�����'�qY�c�O�'�vТAM��:�����.9�qxG��'>(X6)C:Z�AExR�*Xx`ˠ.5N�,R>q�����O�\궈e����6cקb�~���y��g�f���I@e�O�U��*ɃM�n�ơQ��h1#oЄn��$�dmX���0�M��
)��ټ�q��>�ċA#�/M"�����,͌ȳA-}���6���I%d(�	����Z"m�P��6\� U`S�v��5`S�	pyӅJ�,�9'�A���' y�KSwL����ǶWq���A�]�:�A��o�'>R�6�Ͻ'�$x����)��*G���
��ѵ&�<�V��bO��w����@ �X�� 03��Ͷ��dK�k˼!��?��L0wD�-gU�O���E,�ݎEC��1~�}��nI�]Ĥx9Xw^�4Zq���D���A�$�X�H�}"Ɇ;W&�|E�4FH��p��0N�'30��2A�.$f��zю<�Q
S��-!~�2���-�t�>)�;B�%)uO��yQ�4E`�,c�BB�	�+x���ˑ���k�&ޱw�&��Ҁ���$)P�Cc�k�-�|��`�J���'�R�wgM���UCGg�|2�l�ߓtv��W�H7�\�+�K<da4.�*�DU!�I�}�P�+��"g���a{B F�BN�z�f
�i�xx���O�4P�- �H�2�Z��`�@Ѡ��
�I����xqхԟ�rH����4+!��� {lV��P�-�����Ǣ\s���&E�
W*t�"(Q�9�~(��M zmQ>���R���Bc��:Pw�y���6y!�dX�0��A���2Z�H):�.X	U
�m�O��b�@ܲ���qO�:�:DǄ�
�O�:^6�q���'��jǮ�;zB�O1u�@���'_�R9�ӇDo؟#��U�!��9s��&g�:��4�W���gM����­�g��!2�z#A��'�)�g"O]���F�,�|����C�2'��q%Y���k�	iހ>E��m�VO���Ee��}��]����y"�+ڸ��J��l���+�d�'34���@�S �ϸ'>*�IG��	8 Qp�$�0(?�%"��< �qs^*,O�-�ǁ� x�rd�ۊ���K��?���d�Xa�%�+yH���'� �BH-�X�'��R�f^�/B`(�k� iQ�9D�� ��*�E��^���3��B	-��	��>�G��X��?q��e�h�d��T��/ ��  $%D��!��JN��@J�7���B��$D��x3��nT�P"�m� /��zs�&D�Q��l�q�v�?;0��&,��dSG̓��a|��ؠ�A&���,��.ר�0>�FIL.r�N��8��� �L
_��Ȱ�%/�J���{>d�0�C�G���'�"�e�?Y��#�rИA'ҧ{N�Mr���j�r�ZW��X��ȓ�f��U�0|��0bݞ�nIJ�kG�ZO��g�>����O ���ߤQ(x�JR�!y\Hq�'$4$���t}�i\�,��d���R�[ �a�B���?ٲ�(4̓U�:lO�a@V�A%*���
խAK
y���DP�@��<�g $?a�
V�#�$ui��`ݹH��A�mM����F'Y>� �/#D���%I��	s�ĐX��A�^�I�$��<q!�'��;	2�針�yW��d<̲ KI?Rq���R�y�x�\Eh��)'����`J%h����Մ@Rƈb*O,����)RY	�}B�����O�(��ċ0�p=AVA�L�j,�r��-�Mk�IpZYb�@ʟ]��H�m�����PgU�e
���u�'Ab���]�y����ڝȍ{�JH>z�P�ZbK\�zG�	.UC��C7b�?��� ��`�Bݑr���ವ�j7D���#k��~�P�%m%p��D�;����͐��?�vB�L���C��~�@%ȹ?q�?�h��ï��N�lL��莌l�>9#�'v`t��i�	�r�̖
w���c����0�s�Qq��\�Pg[>;�ly
��
�=FU8w�̗	�Ń[��O�����D
FL���Phh�� �k�q�'�S	�?�Ņ��&�0�&\4}q4�����N4�<чK�.T4D@`θ�b}��c�{���RۓA��-����H�vL�1?�m:$�] Tq�@a00O��3a��D��B�
�`��ʲ8�y2d��b�e�]�b��ӓ�N�^�~�[g"O걸hJ�~�mk� gc]��*�=�q���<h��TC�&���э�n#��v�A���w�F��2�2yG��x6��j��H��'�м��ȉ:\L�o�� ��D`4�ˉa��%i%�Q"3:R�k@J�A-��X��X�U61
��?9:��Er�G5(%�@�Y�f=
�����#MQz �?i����rxrB��<�@G'+: �ai�<�Ly�sFů/���ba�`��+�O��>kL̚2�Q?��=ѷ-��y��Y��m���yZ���>�� �	�k����y�s��d�iۀ�D v��s��_�c��^���'%ѝr4�x���F�<a�ED�D���(��;`)bV��B?ᶇ�k���a��2B,�B�U�oy\��&h���*l#t7m�� ��r ɇW��I�L4��¨@��D��\�>9�ݰ6�(c:(x���Z�¡��#�My�������ɜO��;�	�%�����!܀H�H�<���D�N�"~J�� �c>����/<iT����\�d

8+�#I��	�"m|�q�+U���5�ʎf?^B䉰-��=���MK�@���3�*B�Iu�<�QwƠ����2Ʌie:B�ɇI\~�*��D MUV��䃝V�C�	�	h���/@a����8dP�C�	�~{��:�Љ>>ѹ��^�4�p��$��y��!2H�7V,�A�#E-f��z�fI���xb �� 8� K�"��p
���O&�XW���[8�>ݸ��V�72�{#;2xl�P�%D���Go^��;U�T�ND�������׬(yg��f�>E�4�@/U-�Z7fR4L��F �y��U*
.�*�۟QZ���2"���=��CUe�)F�axl"!��	���_�N�Ā�h��p?	 �ײ����2�ݡ��HŊU#u.rPQA��/�C�	.g���2CA��r4p����Z혢>aVLʼ/<,bpj'擢:UR���(�KdYՆ�W$�C�I*s
�r5�2V�c�e�b]��	+C����h޲/��S�O%��;��ܹI�P5��@�	�:̈́�Hq4�"FNW� ��yǈ�;��x�O&�sΐ	r�q�
�HV�����2X�&)�Q���$H�4��I�ƈx�JO�6/�����&=�	�C&�C��)�@��E�+��A�Ęx� ����O��Y� ��0��>1���#+�8�kج8�My�l"D��P�ܙ;�h�V�D���DK3o�<9���4➢|� `�@�EI�M
���2��joL�B�"On���&0zT�8�)*+�q�"O~�j�ރ.�8 �0��O���Y�"O���a@ݬpz�y"��Y�%p!"O�-���1_ʕȲi�HI�` "O�1@��]�T��iD=un؀�"O��知&�B�+2���LG�((�"O���w%R�r]0���ۄS醰�"O�ѣ(��3e�y6�����"Ona�`��f�\9ԧ��h�As"O�	��
[P��7��(�r�6"Ox��
3�(��d_"�2���"OR�+2�в."�X1G"�L8f��w"O�I#�]�=�8c5KB3A.X��"O�Pg����Ѡ�+݄(�d��"O��$�X�~0��ϓ�9�t9�"Op@���+��"R��#�T;"O	�� rA��+�O�ru4,[�"O� #C�K�M����1+U$`o���'�y����l�h�����**ze��'������>Z�A�L�2 ���'edlp#'Ѩ" �X��b�$����'�|�ؗHǺ�r�������'�<h��ߕg@"4jr�B�ﴼ �''y+c۽Qa���|[z,R
�'{,1' F�}����o6c��x	�'pU���*�����C�P����	�'�b�� �>�����,G�J����	�'�d�rU�I�G��xH�a��T�X�:	�'p�]�j��j��T�qE�{*���'`*����	T��A�W(֨p�����'|�r'�#� ��fZ�>vh���yR��9yv���!F�'x|�Ir�Ë��'�|]����!d�X!Эܟ��B�'6�@���
�L1W�OO2xy�'�:M�ՅT%��t��G�{|�
�'�r�p��]q�(V%\�!(  �L���'B�*ç��q��-N@�����s<���qm����DV�z[e����0|JGA�>z]���OԐ7x�U��E2t�$��o�F	q��%{�X ��ӷi��i��I�`�$�P�T��74 L�5a��`���
w>y㇩Gl���BBN�8���jϧ0|�r�f�(&p�?O��𩉑R�J0卍�pF��U	�|�!����S����'at@��'K�B�kU#Źq>�1JB��,⾈�T�=V4P�Y�y�'M1�,�r�I�$$Lp�kB~���>��L��&���ç1�Zi�c�-�e:E�S�s��'�N C��T�OH�A�OQ>A9 E7��I"lQm�DHT��Ovt�L�$���N�"~ґ� Hl�bt�Ӫ:�n4��� �~�@V#{��O�>)p��͞	N �̏�SŜ���"0D��U
��W��DJdk&o|Z�0�),D���a��s88��,� 2�T���,��9�O΍Jt#�uX48#�Or�(Y"Oh1� ǒ�c����P��`<�\C�"O��!ѧ8�r� [$)��"O�,Y��#��0x�.��)�c"O�yؖ�V����I6/͙X�P4;c"O�qy���$	��1z�oU�$}�9p�"OD���(4�QA� s�慲%"OI"I�b�6գ�FA�2Y$T�""O���R� ?�i9��UL0@�"O��9j��(@�\3�钾�Vh"�"O���J�=@�@�*��H��!;�"O"���,:�H#�ְ~:��"O��كa�/]���k\�T�I�c"O@��#Ƨe��+$G�l)7"O�dÖ2R���
�K;*�\4�0"O� ��h�f�	w��5*,���SQ"O��ТmV���� �4+N���'��`�U˘!�HEK�*��V�0��'b*�QC�ؓI��J �]99���+	�'f�qI1/Ūo�^d��'��*��H�'dr���˃2�v�QG��� p���	�'�,�{���~M�V ͉�hH	�'�Ԡ"��_�6=����^�p��'����.�2��qa�R���b�'r�-Õ떖���a�gT�{�x
�'����a(:�ШA)�!E5�h�'����AJ�%\����B�x��'�2�qB�D81���W� .��i�
�'�8R7`��|:ta���B'6��
�'�.�KNw�Υ��R����	�'_�MeO^��
��4�Љl͈	�'=8��'�s�,,��jû	1��	�'S��1��S4P r�h4�H���E�<ya+ʯF�xؑ �Y�	 ��A�<�!�̋|h�"	K�vl9֌�a�<A�cѪD B��t�<X#�	S�<���
^2$e!f��SA��)$i�R�<A$b�1}�p�Y$��=k��	ɐ�
K�<�7���R��$��=B<���jn�<q�틧W��+��F�����֣�j�<ys�z�(���4�]�Cg�<���U�uHb��F@��T �)�Yz�<a S��j=�T`E&jBz��&)Zy�<Ia��LU�U�A	r2yy�B@~�<����,�t,Y1倠Ip4ab��`�<�#K�r<9�4#�����x��B�<��m�!d��%�����-�<�@���A�<�d2&���Rd֋P��Ի`�KB�<A��T 0�L��'� ��$�E&�A�<!E� �C$,JJ�Z�XԈ.s�<�D�$��<cS��(G���!O�k�<�s�;�R,���X��P;'Jq�<yaEЧ!'� Q�៮#4F�q݌�y�f��dln��ۡU�>%�5G��y��8(��"�(H��@�� ��y��IԔH���/���4��.�y��O3{���b��V����œ��yB(�4M��T�-�Q�$&��y���y� X�4�	
Of���I�1�yB' $p�qqv� �FĐ��$����y�BK�u��!���&D�r��4�G��yrL	�%A	��Ά��<ei#d��y�-�Ȕ�A^)1g�c�@T:�y2oIB�e�E��&��(�;�yr��??�:�`�G��ʝ�t�6�y��A<,��(w�ψaݸ	r�Ǘ��y�+F���u�^RൃƬ�y�Í2�H�!�ō�X��e��U��y�Ƈ��t���M�N��i���;�yҥ^(>���6�ƩE���2��ʙ�y�ˋ�.mx�a@�=� �`�M�y�HN/Q�܍򔫛5��!���y��Ȃ ���R��۪.Vr�J!H>�y��ެ_Gt��`�'tܹY�X#�y2A_�g����-W��P���_��y�Cϭw�DӞO�x��$.�y�/�4�P�1�/M�6�уSJ��y�%�f���S@�5�~�p㮁
�y��+lk�}�@�1x���G%�y
� lԣ�f�(I�AӥDG	=I��y�"O<�*у�I�RՀ"Wg�B<�"OmѤ%�c���� �$�,�q"O��dd�!u]T��� S�" �sE"O��؆�j<P:��CF�:�R2"Oqg��-����S;)5�1
�"Ox�B���A()���>C�lj"O}	0dHi/vY�m�73X���"O�)b7㊄��y�D��i"O2L#2B��`j�KWP��e:'*Or�7T	A��)r���B��\��'g�������d�$9d&���'�.i��B�2�H��[�5%�8��'�p$ٖ��Sw��k�名.�*�Z�'dH �I�-J��ٴ�hh��'��xX�,�6x{U&�r�d �'�����Fڷ"ۮ���d�'xj$��'�j�0!�Y�`����	K"oݲ|��'�hpQ4g��x��9z�g�b�H���'��(e'��5�N�P�T�٫�'-�!���< �z�����)N�j�0�'��a�I��_�n��G�څ�حr�'v��Ko_*'��h��(� cz��[
�'�ެ[��؛b�J�	@�l�:��
�'��3��J�H!�D��f�p9��--��e�I�b���y�M��k��Y�ȓ/���(Y3V�҉�@ �1l��Ʉȓj��7�]�L^FX��*-l�<���	�zse�sO�m��F��@H\��*�#0N���@� �) 2L��ȓ=H��)�㚏i
�1�k+��X�ȓI@��b�X�m2�J�A$f��ȓ(V��j��BO7�a�i��;G���W�>4zՏ�yt����B ]��	�ȓ|�Ja�4�R�a����U*�L��{U�9�B�S�EH
,�ք�"|��Q��\�n�a%���G3Ry��g�(��ȓi��D:`+�{�t�!@+���B����ii�N>�x谤�>h]�B�>� �!�,�0~w��9t���?z.B�Ƀe"ةQ!cG+\�h�g�&d�2B�	!Fn�2����ZI����^�"B�I� ��S�o�'q{�=sqnԧ6ưC�I)O���2�F�(d�����P�S�xC�	��k��[8��dZ֥�$0vC�
"٠Ĺ!�9���Kf�ק-:C�ɍ
C(�xbh��{^T�3�c�RsC�<!��8���9o�D��U�Q @�C�I�Hb�@���)d���j�	>��B�2^T�}�o�	�ƫD��zB�I�9���+�+��7�ޘQ�� -{n�C�I�#nĔaT�޲���2Ѝ��F��C䉢&�ta�D�\���]--JB�4��	3F�=J��$)��M�C��%P!�\���}$��H�$��(��C�I�}Ռћ,��!Q|�C�?msJB�ɑ6����29�PX��	KR*B䉑<UT�ի��9�(S��L�0<�C�	f���3��<Ϛ1�.�C�I�-�x��qbߖM����Dd�lIa"ODcg��%z�(�����AO��y�#�5f�u�� Z +�U�2
��yfӪ�����FK�x�x�81���y�#�9<fT�H�G.wZ=kʖ2�y
� 㕥̯[�D�ьPb�I"O�� ��^�_1�[�( 6��:1"OҜ27B
u̓���=)�@��"OhT4o��>\l%i���o�
��T"O"�&�\�<�DHA��4���q�"O����c���p���%=�ֈ��"O��'�m��tǅ�4XH�"O�pѪ�>0�5�QF̝Vx.P�3"O�x;vC�<��D�0w@��f"Oȸ(Mɤ!Rb�Q�FŉE<	�"O�u@����dAhkP��x�"Oh�{�b���X ��BI����"O����Cp��X����'H8V)	"O�)���!� ����l1��SU"O %)C�-n��PE> &�y�"O8l���^ l��� �h�*��Ђ�"O�i3t�>I���1��*,�J	�'�+1iZ/A
� �æp���`�'��@��dӧ>=`�ʧ+X�~ɣ�'ن5����;�)T#�Y��'� ���U��=�@!���� �'}��k�G�20�BS�Ł^�*�'��� �ei���3���	z�s�'�E���<n.�҅��6{:=��#܂D���.i�@��
�)&@@��ȓ^��q�e��f�4���@st��ȓB9���S#��`�:��J�KJh-��Az�����0���d� �ȓ=��@����<H�獁�P� T������������V!WN;f݄ȓ\T�2� v�x :$D��1��,��,�*���t���Uͭ}-���vx��U�M�5����	U�g����ȓ,3��.�99G���$�x�� ş@�<9EA���pXV�*Q2XW`~�<9 j�;�b�3Θ��x�[�c�t�<�'��:=f�*�%F0uY.�C��F�<�*�)<��Q��-
4�8xD�B�<I�hU
[�\@�AY�f2hPi�dK@�<��~� ����W�
��rϋ@�<aR�ԿjT��Cև}ºm)A�He�<�c�¦*Y�����i��)��,j�<�0�
pHr� �/@��4+^�<�+Q'|�\ 0�I�D:z�+��V�<�q�X�]�d$�J��HP�#Ff
V�<�6�jo����M��k��Z�<ᶋޫ��)�N�'q��D{�j�z�<Ƅ�F�@A)%_%4[�#���x�<�b�Ό	�T׏��Z8�t-Xw�<9�M��1Y,jᔄ�Rp�<!f�8^���J��	 �����Vl�<Y��AS���Ǧck��M�d�<y�#�N:���-´e��y[���U�<�P��Jv0@C"��	E�%3w˒O�<���C#�T9�6S�h��)�ĥMH�<�V��p�lxW�5�t$��F�<Iu�6�(��"B�'���c�[�<�e��o�&\)v�� ��}I��	Z�<!�_�Nj��V�
�"�e��&V�<1���H�Z@A�Z�.�B�O�<���ս8]��ȕ@S�Kᄄ{��M�<i�    �